BZh91AY&SY<a�i�x_�`q����� ����bF~��         �%R�B�=�R�m�UEE*�liA�P�JI"%J
Em��$UU��T�T-�("�I��T#f��
 h�r�����H�A*Ui�֩H�M2�B�%"$��R�6� њ�60	��R(
�
V�l/ c�H$�Nj�*��U� j��7F�!(%hUV��HU � QTB�AQ(��E*���P�ĤJ&��� �JUI*@��    +��@���I-e����n�+'X��T(ɕ
��Q����m�gNTV�&Em�&������%IT��/   ��J +�j*�R����
d�(U�.�T��R�*�5� ']8(�T��� tP�wj�����QG��J	Y�  �d� ):�p�*���� wJ�4�qT4ҁu]û�wI� �.�R
)E�Ӏ (\.�A^�ڔL�E"%mR�Q)<   �� �87v����wl �-�x	:5��� ��+���P���.���w��]��z ]�d(�B�H%Uc�  �<��U�i� �]�*�S�,
R���:�E���v�ziTs:�m��Z��ҩHg��@ sU��ʩ*I%UJ�IJ��   ��R����
��e!�B�Jƴ�Z�i* l�Z�PZSh�`�J�{nm��Mm���J�U� R!R��$��  @.� ��4
�` -��( U (��hц�6�P�0� �6!UR�����B%R�� 7��0�Z� �@(ڬ �0 4Ƙ
 ZB� 1� � -4 HP��*�I)   �s �  �@��1��Ҍ 46�� *�h&0 0 4L� �v5i�
))���    jh� ULh l � ��(h�L X0P�`(PF� =�   R  	*�L�)Rd�ɀ �2d�b)�IJJ�&�0ɐM4�L���I�@)��F�1A�A�6�d�*jR�Q�� 	�4�Sވ�S�<�4`�� A�%$�"�����O��@�4z�����鏔�S�\��|�e|�[���y�q/��w��>�#�����z��(�*���z�������� A?�D@U� W �&���U?`��t�DDG} P_�T��"��������?�`?͗�0d8�1�^0a8����fa�/N0d8�q�0�x�q��'3��8��^0�x��0q��a�'8��8��N2q��<`�8��8��N2q���d�'x��a�'x��^2q���c�x��N0q���a�x�̜d�'8��N0�x��x��0q��`��8��N2q��<`�x�1�N2q���a���8���2q���a�x�g�9���d�'8��0Lq��a�x��2q��l��L��2q��<d�be�8��0q���g7s'8��0q���d�9�2f2q���d�'8���<g2q��a�'8��0q�10�0񓌜`�x��^�a�x��0q���3�&N2q��<`�8��x�8��N2q���d�n0�^0񓌜d�x�<rq���d�x��^2q���8Øx��C�<dI�N2+�x�/Q������2#�xȯA� <e�
q���(<d�"�N2��FaC��q�^0#�$� �^0��x��F`^2��xʧQ� <eG���2F`���2��@x��"<`����0#�DxD��`�*q�s
q��'P�
<`G��N0��x��D8�e� �N2#�@xʇ�<dS�(q����aS�(�N2��8ȧT�(�a�D�<a � �(<d�"�s*�LȏA�
�dG�(�N2#�@x��8�.e���2��E8ʏ� <d\aG0��@x�/�(<eS� �1�U���0#�@xʧ�*�`G�*q�̠�ȏ��aS���^0+�@&U��
�` �(<e�(�T8�$ʩ�2�q�^0��P0q�&x¯U�(�a�*D8��<eW�*�C���a�"aC����(dW� d� �S2��Qʡ�DN2 �G�`S0@3*Q8�!�P0�q�3*a�'2��'0�`x�q���2e�/2f2�0d8�q��fN2f0񗌼a�x��̼e̼d�/0d�e̜e�x��2���x�񗌇8�0�<`8�q���0e�!�C��e��0�a8�q��!�I���N2�2L<`8�M���`8��^0e��x�q���4��2񇌼e�'	��q��N0`8��q��x�q��q�e���2f ��M?=�����������_��]tQ���c��If�(�ʺCa��SX-V�K񈕕�/]6鉛D�s#�x�n�*\�x��HC��-X0eVQ�7�I�e�ej�j�)u�`0֖N��M�N5k�ծ�V�2P��-��m��5nV��#qF�vo"
�\6�d���Y$"Y�z��-�z6��I��{�WC=&�$aHݤ$�22�̸����:�2X�Gf�m��K�*|ѳ*����[%lv�[7���p����SwI.��vȽj�3���HR�QB�R�͖!��(��#�E��u0іe�ɶ��kO4�b�;X4�9�^cSK6E�v[�\���P^F�Q!5�q��� F�Lࢡ۽�;)�m�y�4��ddu�[���ݭ�S�e�o�jڔ��v6Ml8�X�3=pY�Ȃ����ˇJ#�����暲sET��ɥUSwp�)Mvh��u+��JĶEj�6�j�C�"2���N�D�i��49Y�P�>Ų��B�-���Y*iZ���Y����gtW:zP�D���V��q�0�
���<©p&Ɯ���W���K��e5��z76�m,���[�v-�+�ҚURT�ɖd@���F����ԗn%�17-h�&�a��:4l4i=�ͻb̧I5Y�f��qR�X+l��,�Yo������*^�n��0r�8읡�][/B@�=�U	A��rm۲�LY���NVwT�K�ֵV!mXiH��J�f�T���<;���I�2���L��/6�RŧY�e�ͭ��BHB��Sɯ�,��&��6�	jBΊ�d(�@�fJ$l����PEO��`��Ɋct�!�]^���G)�O�YG+d�d7j�U�T�ԍ�(2��\!JZ�"f�9�Ӻ �*�e<���tFPO,�W��Ƴ3Ue�M�Y6�޵z�u��o$7�
�E��f�"]�'��&3w�=������(�a%dr�ٳ��ݹ[s/@f�tl�8@����S,Vh�.��p�sa8"�Cj%l�����'�W$C�v��@��5������l6J���I�]/[��4��!�)�H�n���SJi���i�;�iJ���o1ǉ�!�ͬ�I��I(ˉ�jC{�b��)�Wgc�Q�,��.���	Q�Y[���%�a28�z�c�n�j����֓�n4�[,�w�֭y�'`�U]Q�2"Sr�IUJF6��^�*ڥ��$�
'@�Rk��ӌ*4�ܸ[z� ��^��rͭ0]ʸB�[��3.�x���T�+�@j��hڂH �Jڌ��@s/r�,�wt�o,q�,�MV̅�SGX�z�(m9�U���Æ�JH(n�YF&Hw.�����5A,�Ɍe* BP��tU2*�D^��l�PX�2����i䱻�kl�BӕB�V��p])��U��̘�q�l:���2Bf�w{-ubf3s���S1���%@��kPm��P�J�ݖcV���\+c*��S�b9%�
543�K۰ovh˨U�h<1'+r�1�rdђ��"GY[n0s1�X��\�0�.��^73m�$�A��7�4��]L��
aIyd<s�MVj�n�1�Ь�h;M�
�ff�Y+�n0⒫j���*�iԽ;W�ujV�ES��-����nff��P���bM�d^uS#6�ވN�g�l�7V����ְM悉��"H$���ִ)&���5M{� 1�ӕy���4�Yp�䘣O�͹�'+)좂�������y���&V���n�K�王X�A�m�w�&�z����ի+1k���0l�iL��;/l�I	fV�T�8��N���l\�H�F���Oo����W�*5�.�C�
j�te䦶�w��f�U(D6;��Ia�'O&nӪ
T�:��t��ӑ���#�1^�Ĝ�p���KЂ`aUڔ,��[P���X��lR��Y	 ��mT�^
��K]Ӹ.�E�4Q�9��A$�U��uO]����0F�-	�o&i�����Xh#t��P!����b�(�cb�T0:���y�^�8º�q]&Α�3�%�8�n2�"�1"�%��j�ʢ�a�RVI��ű�;��]Y���N�5ƚ�5Z܊d�,&�EK.�U[���j޺���T�^�"7n�F�Q��/X+j�����������%�U�a�j��˰E��p�8��4�7k'��۪n�:v�F��bb�(�be��\�T&��)���Qse��Ha�+FV���M���?
Ĳ�X,�i@%'��Ҵ�{x�ɯu�@���\�Z���Ef�𥲎n+��>:։���O/X��n���7�����1�'vj�ں�����i�jf�Pt��c �&�
����,Ӫ��7��vXcp*&n�vƄ���P��Aʴ�˂ �ݱ�DM5����F)�SՍ=�9!��t�+���ea�*�-�C2����&e�ʶ�H�VfP��Kv�j�n���J��:��b~�é�2d�7�s(�`!��:�*έ.X]��*�	 Ż�j���7��X�K�9�iȋ��A.�C���+�� �t�٬��;),őٹ���8��Td��$��Ժ�^a'V�*�G28�Y��r�kuc�2�cn�s��	gq�.���B��T5O(�ܣ.�h#�p&2�uw�����9�Eb��;�'Vo.<.�U�tǡ�U�uc�+�Դ��6�uQ�M�w#a-��jm��r�go,�B��3eՊM�a������UYY�R��ٮ̸`��ha*����yFM׷���g����n���i5e[s�i�*��C��6%��^;%�1��L�[B"��GI�3�X2����Ke���G�Wִ�茖��#��1�Xݧ%�66+�9uG�0։���Hi�2��N4ܻ"�v�N3��U]��b�a:ޭ��I&��(��8��s3E�	����$��%��׵h�{e�5���!���I����3QwL7��ܥ4IG̱���j
�ӭ�=�Xa�j�/l��!�R�{��@wF�#0J�M��^M8�1
cN	���AQ�mV��N���,��l�M\�[�j�@�X��B��f�"��4u��eV���fQ�t=��5M�嚔ޗjGreK-����/Y)X�QcP����jOaA�p�P�S&�+@f��}`-��(�.��һ`7�Z�G3P�ʹ�E7cs^�m���)�b��.:K-��2Ƒ���
�6���4Y���*n�w*��q�3E�ûu��J#+V�+*�ے�"&���/4l �;q<U�ļ"D���N����J����e@�ݴX�{
�ً\t�f��N�:����'	�y/!��`��p�4�^�b^��mLf�Gv@��f�x���F���G��ɂ�EM�qϧ�/M�շ���v^���θ�7�v����B�M�Յ���Y[��p�T�W&Z�9k!N�K&�)�Jhi���Qfn<�Z�������I7UU��W~�ŦM\���V�+l��A���p}��4��=`�0��PCM�Uf�@�{�:��>,��5.C�,��(��bV�nT�dj�� ��j�� �묀M�t\;�ՍW��_"F�_PvU���R ��J��'�=��K��Ҳ�ݽ,�*��R�R&�P7gA�H�OD��tò��������Q��pm�-^2���n7 ���%%H[�y!	��md�e��lR��{dA��lf�!X��
�J�*l�+���>a��9�h��V�,BL����A�&��bX��*��%�B�Ld-�]͌��U�-�{t�v
���W��&��@*2��H����<��E��<�+sMn��V�m9�iC�p��ze�-3��y&�v�ch�r����#��36�z���*2��#�NVd<�Һf�)z�@�1&�Dv���z*͕�n&%h8���ܭYXB�T�c��FEt/ƌa˧�͡��U-T��̠���e�QX�J���1�f���ݎ� &�Th㫭�����"��^K��7���6�يџ<��5h��gB�4*���Y3]�td8��̻x���v1�yy.��kp�54�r᭸�ѹU3#��]�O
	�BF�c��Vl��2��j�ElѬբU��X���+.Ç&Y�*)�C��'�7̘�k�������h�&7S�Y��l��vA�x�d��h��	۸�CA���]�w�
�*-��қ����!�n�E��Ӭ��ӈ/Z�,^��<��'#�6�6�m�ެy�Lu�[O�H�0\Ǘ���f햴�/U�窬�̼� t�V�r)���0�ڽv��]3���N��$L�sS4և̥�d7�J٭̆�N��f�N�L��X�Y ��<���J���Rˎm�1��^=�l�խk7B�����ݹ�r�i`�B��4n=rP���ÒћiG��J�]�@�.;��[d� G�Io+-<��]Šd#K
��r�J�Kt�E&��%'UAc�G�,YyCK�f�:B;L�l̥hJ�D݁��v�"M=�q�8��Խ�t�C76PklU��ݑ�J�h66��xl*щ̏�a�/f�j=��3�(�:�U���C �B �E�e�zN֙�	h"��a�l�7�R�������/
+�f�f�M#�Mz�۴�iܫ��W�V�7P�^Ǔ�I�FZg
D���xI��ܺ�PY�)��Ue6�R����Zc8�c9u��nk:K�SUY��}hl̀�yL���yYe+n�!�����ts��s#4-�f���f��^�nb96��`@��*c�AF1G(�;���+�'�yA���̥�&F0�w"�A�;���,��b
��	�v3A�L6uD��ʡl�@�Jﮅ�/X0�	W�1���vEI�0�	�y-�9C-K�h�Ԕ���̨5�*�|h�!ZN�x*kYBD��tiF�۳��ķ;�,��G��P�m�kR�QYW�Bu��@j"�G\N۹wyz��Y��Q���֒���I��5���E�e�;Q�
��V����5ּ�E�u
�7C��
�Q�vA�.�����iՑ�"V�;���d|mN�gCޗ�i��RN��cr<x��Q`��a!�[��2��1OQ�C���{:���c)�3S��+k�L�{�r�ZHq�l�mI�7�P�ԬhR����ށ�W�*�e7(QT�YR����!�d�C�r�T��[�4�!�<�j��/Q�-�X���ݨ*��W�N���6Tx_>,et"���а#H�Ժ���'f�xv�Cvt9zq`�[FMP,�薾em��k�˴5�)&���i����6Yy%�v[-f�+r�j\�R��J�b�+([y�2��z��f�	����iMM�y�U�e�ZIl��Z�i/)W�W��:$J�]����7��I��&�	CV2v;��	�sw�R)�'�R֭^,��6��B��%�N��zf�f@s�[�n�q�V�[&�C,�y��U;�T����F��SB��̶XJ�v���5�ٴ+�_��H��AG{#�c>��j�;ʖ���.�ȱ���Sf��˳�	��C%�B���L�kF8��n�x9���Cv�*�a�V(n�����)i��R���;���]̣�yz V�X(���l,�Y���d<���nr�:j�Y��;�:
�NV���6�����;�V��Y�� 0��x��V)d�و�h�xpj�͗ ��ꥩ��І��Dͫ6�O[�X��6���7`0� *wb�SۨLA\��ő���M#	y���[R�'Z�p )�)D/n��7*��=Pc׷-���h:C����(f�qȞ���[�%ɩ[մ^��,�$��ѻ�04A�T�Y������ ҩ\�E=�)���H���3-(���+P���v�w��^
M�
^��i�䫿�n(˩��b�N�߁6�k)�^�7ڕ�d������#NE	��q!Z#H,��jɢ�Z�'*Cl�b��#b�2V�7fk��V�j���V[�%�
P.�;���R(�(�q��cGQ�[M7�08�X;J'��(�>�Ь�o�`3==΁s��r�`�(��i�VxrмVoA��gT;���꽫䶓�-X	�)D��=��p*��@�c/�b^��aC���h�++]_����q'�G���U�D��ݏ`�����Y���x��H�\��M[���#p�����q°��5��eiٚ��B��m�!ټ8�Ea���������88.�fE�2�'XY�W		99r�2��TVB��,�Hv��'͢���\<Gqw����3^�O�ġ���xc
&h�Lz&0��2�kOcA��e����FШ\v��Y,�;DǢ�x�x0h�M�e��M�=EQ�we��0�]�b��M��]sMa|& �;	�bgN�(Vc69	X�QzNi�he�f�iQ=8H�<��`�ͻ@��������%���VR:�ɉ��:��ҢFr0%�f�Țf�\U��3�bgNG�@�6�n�e]f ]0B&��nn���⸰�3J��"���q��|�;y�=�N�#�0}���0��p)�wC��)�-
��n;�n���^	A}�W��&M�u��LG�W)�����4K:$�q�1��ۋ�V3��<��+��bV1|XZ�D�١Aq:���h��nQ-����s�p�p���f������Nؐ��s%���'0�.'Y�*=�by%�8X`R+�]��GTgC�J�-e���Q2�X�n�DurTՃ��G��H��X[
$�q7�0@Pi:pmE C�B�A������O�&t��< �A���������>'Ϣ#��e1��f,��?6�G߃��"*�����N�h��rz��ww��w��|W�q��H�ÙW�����1�m����U��pd�{���5}.��`����ԋ����[*Z3�u��:j^Y��]�N�A���,�"��Ϧ���2��6��wxα�WV����ʰ�G�x�`���;�oi�x&�;�-t�F�ol�O��╗ ���ɀj,qi��]esۍ������ކL��
V1Wh��f�uQ�3r$(k�+�zC0h�+Y��/���7�ӑ�k�̹&�x:�-�]�t5���B��vZ���u�\2ȩV��g��-�+�kAͲ�m���ռ���	-��j�yթy��s,�J_7�}{d
`3k�1>�ف�v΃2��3�M+ko��{|�uGNX���v+��SJ���T� ٙ7u�V�v0���7�U��\9�KA�pZz��s��vҺ��V��;�i�����y����ll�����I닫QR��w��-N�-2��QЛ��t��%u�
����E�0�	Fc�j�bڰ�U�Ô�y�����]^V�J�� [�^��o�F6k��̼!�IRp��e�N����{PDQ)�He-��u>��<X;����Ǳ��\�/��f�z`<�1�^�"�kj-ޚ-+�^�~�+�q�]��.�u"5��5V��i���I']���A�i��:;���lqb�*���IwV'n���1>1�(����
��w|)���mblt; �;��rvw�u���k�l���Ɲ:t�&�.�
F�nJ��K��}-�:�l�y�.�Z�"N�Ů�{K�y���0���їJVh�e�NQ��\�M�Z��u�oxT�4c��;��>8�r�t��ͮ���m,>΢��u���[�l��x�4�L�&'[�ݞ��M[�8�����c�*o$wc�F�r�(Q��UG%y�Y������w��F���wb���D:;}B��|5�r���h5�֣�^��Y��ewnp
q}�sP����=�f�.ۮ�
I���nm�U5���!֏c���d?[R��-��ʦ9w��%�ж�+{����4�b��N��9l�hmң[8Mtj���!HZw�������չ� ]��P��3�r��fN���﷑�+�:*�t�#Ç
Fʳdn��[�iB"����͢w�ֶ�5�e"���Fo�k"�ܘ��L՟q�ҰQ����1+�I9ZN�[�B�p*�)�B���`�7����i����:�hB��T�{�|�q$�[�w\��s��5Y儿�+��wS��&�a���*�E���,*�=�����Nt�<���$�m[g;{&ޓc�,M57zm����ǰ����z7�����:�d��~�e����<�iv]�i��>��*P�У�t�Nnc�:؂�������*�#�S����r�C�E��1n
_�1,�[-�w��1��X9y^�[p[챇�o�oG���/�;�\�D�-�WG�+��e�6sSa���o]���J<�ӬS�N���v��W�U{��N�:��L�3H�Ȫ�"'˻��\���N�=�w�9�n�ڰ? ��1r��7��i�4Ԥ	kUx�䨕YG���g�va,�T�ֹR��7o;�og"۴��"�Si�:9U�ۺ�W9$��"w��Vs�Y��	X�8���̔%��\��ۭ��;�̚s�f�V��}֨���{p��c����we�:��Fwn� �+w��Wq�r�t�U���̭�6N��AF��4qt鮒6;4i�(Q�45vt��80��!G:�wh�z;F�7ww%����o2��,p��=��7��Us���o|��vX�Qxv�_�%�m��\&N=*P#M��*��GKM�{=�l�+A�r�ͨ�6�Rڬ�z1����L�n%+�8����&q6�8o�Y���n��Ѫ1��8�[
>����DŹ-�[X�\4ݍ�d�A��i���-�9ƞEu)w:���%�s#�]���S��C�ڥ�k�{,���t��z�,��s	W��1�UR��nF�u�X��y>�I�`�aܶud����������A�C�k���Gl�ybJ���6�{6���몇:^�j��ӕ��t�q[(i�k��Qlv,����[T]v"�xo 9�hҗ��#��`oe��rㅛ?-��3�aWv�ݻ��]CZj�l�^�en��Y�8����5�V�t�t���}]>�;���}awZ!���G��n������R2�ZJ�2�*�ׇf���B%������~���:U��L���Ξ����Y�y6��"�)�����o�u�	y5����6�w��b߶�j�%��v�P�WNݱ�K��/��d�X�2�b����-EQ��Jvr��}'P��mg&`�;)Z\�P�q����n�ܮ�>�{o3�n��ݶ��(42䬮xMu�8�b���ʀ����rݮ����t������F����X*���deήMu
U��_w�,�I���嫾�k9m�Qa��S�e�wRu��:\�Z�h���(ygJֱ�͖�sc���X�*2ȉٺbTnl�&��6���ֻp"!�ϩ�b��3�����G�!�
4��Y�^��KL%VE�,eӮ��W���^�ML^f�g<�i��\�I��0�O���-;2�QV�w�銖z�"��:�<�A��j�wk�
�b�[��y�ݼ�>ɚiy�Bol��;gT��{:񫢆>��Ȇ�����*K�c�{�k���5�s�L+�VȘ%�8*[����.�$*�!���0Q;}�7v|���VY�������]\��m�٥mu;sh�u�<�E��φ�I��& ّ��#�g��:�iFV��L%d��v�<P�C�lQv/Z��k�Փ�g5�so!Yn���N�f\;M��B���F�9۹���̲�|�i����|�F�Q͹�ݳ�Av�:n%�	����]��y��ۅa�]%�dN�&���z#����nU����ͼ��E٩f�ݰe�,'��Gu[�j�ß��N�z���k߭K���u����S�c��G���.��0����7-v��gN}�|��X���L�<�*��.�蟍��t�g�s滶C�jB��+�e�4�8ݪY��Q�R���Ν^�0eZIF"	^�hTv^�� ɻ�R6 �nA��Е(�q|�Ă����'gvѡ��JΥ�U&,R_jgu�-���m��ܩWG3o�Jָ����5�K�t��hmY��C9b�L����!�u�b�,R�#�r�q"ic�7�(]x&;�7j�E�Lz�%
� Tvs6.����+�dxV&��ʎ��\UB�k4���z`݄]�2�d�i+na�8�5�o,�;!Wi�6dZ�
��GU�s ��t	;���ٕ�t'쬶lb�&�Ԍa�<un��9����w2qخ۶���H��)�Iٗu�)c�JmG��᣹��%�qU�_ZM��+&"jl�6)���ok��gU�9W��e�+]Z�L�A*B��'T�z��ӻM7�>�Z�/�����R����+�+Ŧyճ F��Wj�lZ\θI�F�ɶ�A�]����{�.�}gi���tm��-��؅������	��$;����W`�f�U"y;rC��=�7jD�u,,����IV]VK��6�g�ENً�7����^𪒑��QK���1���o!Ff�5[��]WF`j�r[��:X�}-�����Uq�MҼs��Z*YpYө�x
Ÿ�Q5g��$\�wH����r�ؕpe0۵�2��`�Oq�Z�j�F��YtܜU�R�L!���f�n�C㙩v�Jv�r���U _�ׂ�웹��j�1�i�CT�B�*�@�/�7�{6��P�S�/��]F;���Wp�&�e�@���9Ώ��׻c����'���e�:y����&oev/-gIy��Z!��rm���kˆ-�zh�y,��[�Aq�y�ۻ��혭U팫�`3p�-9��"b8���ԗCFp�a�U�LU�&�ӰJ��%:�Ȉަ�vu&���Na9��N{������Bd!�,�Z��ݯk��@�U��Ѳ��h�TW=#73�e��pt����m��7���D�ҹ�$��
������&u����u��}�)�{y��0�#�WH0�#����T������j��b��gvv�gY��1��+E��d�������ξ��0X_9r�{��Mw$GVle�{n]eN�Zͺ�ᷚiF��Ag���s��"��ZV���أg)�s��98f���n=|�,���3ƴweݱ�,,�SnsW��#�RWu�:��15�A�]��*��̤�0���X�C9�r�)��j_�B�S)V��rXr�UU�k㻸Tvs^��I³�����^i��}��B�6AN� �g������\D��m�\��Zށ�Ǽ��xʆ��Q7x���][��ۡ��f6zS���K��.Q3�y�J��=�������6�iǣ2�5g�#�I�F�dܵwj�'VNޘ緙���-��1eLS c�T�G�8�Qp�3���х��ɝ�����S#�b�%c
¬�z��h�Q1Z���a��!����N��k�|4��&�9�9��/� ���:K�R�����T5�VRW}J���fѻ\Nݮ�,�H^aJ>�ܠ��)k�܌
�{�2��[��uF���v������	ٲ���F����ɯn�B�	���˝�N�Dq��5Qx�f[.����Rw��E����y�9N�H"���N%����)�a�����+C;�P�d]b4&n�㉁1a����"��xq�x*zubx��-���v�6.��m�j��(rWH! ]�ul��1{ɧ�}�T�7n�b ��L��a��ca���-���qgn�Fݐν�J�mE�Tmܴ:��6ʢIm�����H�W
<#�=۴sNp�׾ª��9���Zج�n��@�-�pw��e�5�r�OEwCc��2�P����zK�X���X~�L�x�ͼ�+��5<�oP�ꭉ�V˺���*׶�ٯ��{r���n)�ɇ��i4@\"�h�.F��@5�U�T��-��n
7��Ѻk�3�f4�<�+0�4L"�Y�s��n�4��B:*u�W^ro�]��K-F�4Fk/��a�3��M��Z�w�mDs���Mg^t�}���]�}�j�"�yL��93B�ܗ%mi�fC58�7V�i��ڹI�ɶz�������Σ5�E�iY�ϱ��V�����]܎Cbf[�ձQ�x<=E�#�c��p�����4���_3����i�=P�ya\٘�ՉW�Ro�V�9b�f�o*0'efs����aG���s3%�bW�]�����jЧ�����"�f�M�u��Ic}|��f��|2��FQ/�y��O�����u���w�\��]ezz{�W�;�g9�t��샦!���}�g�!�U?�$�W��-M��Ҍ��f��{��H�Xrj��=y�*h�Ü}�(�(e��5�U؈��yYf�nVs�ٲ�����X�V�*R�^��K5ab���s�{m�q��1��u��s�ַtwu'��}|6'��m�s��T�ut�΅C�l}g3�!fk�9�orug;�'7���ºY��ߑ]�T�z���o��S�M6��(Ѵ$��X�]r��j&�ih^d׭j.9��N�K5��J԰�=􇺞eeZ��.h뜎�1�{��J�ֶ����cY���;R�����/i� �	�>�)3�H=B���sF���0��ݮ[�����D�-�Zir���r�����9]��S�r��:l&�M�1�ο�xU�J�ǋ/�cuV�	��ZT�#ƪ�C1�u��T.m�4�
���n�2�l�� p�X#���ⱝ&���5��Z3�)"��Zuy�v%㝶{������zưb�<5�֘��z�s�f݂��'3>vU�8oB�d��N[�ů�.�:AY�	}�H���{qⓗV�%H�K�&ݱ�O>�}��҇'�zgB`��1�	Z�(gtF�lo6�	�祭V���'3��)���|I�B�e���uuN�&K�o��T��>��#�����v��2V��o+�wwU'*�^�p��9{�q���;�_�~��	ߙ��ё� ~�~¼��%}@|���rB���x$=I�G�	�=����hO����>�}B�=��(�-������G�~@{�����>d��<�H��H~��_x7<������|�y)�C�.���{�=J�p$R��~qWט�y#��+��
�_䟧��W��|ۑ���<���Q�g�_����
!�=�����{���Q�/vp�F<��k0�Em�:o��l�K��W����^+�2��m:��Tofe�)�k�+��I�+)?
��Aeʮ���Fo78vޕt
��RC�3j���J�����v�s��PHr�E�1��	_Q��%�wd#kKr<��;�s���E���Wyx(G̎v�wV7�4�P����}6����kW#A���ύpb:�.��QBe�[��\Op��uv�D��P�����>�V����	�\i���ݮ��let��x��WZ��3��6&���ޥV���]G[2nG�_B��e����ۧ��;5ד�-�wكe8
�;���dӁ�A��;aŽ�N��a�lTX{�U��ub�I���ut�� ����k�̲,t���4��*}%�+l���ؼu�hn�!�Gg���T��y����ө�vnY����>���ʤ�i_�	wTVhU����*!��b�_u�֣Q��;�[�I\&qu`ܻ�|�-.�	[���[�]|ݨ��8�:)��N)�+[���r*N��ݣ��2��J��h�L}eb��z�i�z�͗��e��;:�L�OD���Q�1�v��]D1q!w�	�����m���UmՈ��x�����D����1)L9��G���������{����z�}>�O�������z��ׯ^�~��z��ׯ_�^��ׯ^�z�z��ǯ^�z���ׯ_O^�z���ׯ^���z�^�z�������ׯ^���z��ׯ^�z�z���z��ׯ_�^�ׯ^�z������ׯ^�z���z�_�|z��ׯ����ׯ_�z�����z��ׯ^�^�sׯ^�|~�_�������׽��w�����|�[�Z���ECn�c�u2}�$;G�����I�ٖ5�&S]@�=�����7�T��Z�(u�tk��A��c;X^�R�K+��u���|sP�&��N[!�CѬ���qn^�gBk&��^�am
×�,m�v�5�k�&�&����ω������`B���tgu��n0;=3����6]q�.vL��\�VZ�i�F�p�XR�.����R�`���P�Z���=X��p��f�op���3%vN-���.P���Q��B�9ToB*��0��<cb�R����f*uξ|�s]�$��3f�x�}��gVcf�>euQ[n���^�J��;J�58-��ח�d�RR��˘gK�Н7vsnb�f�m�p�'��n�8+۠�^l�n��o�I�K��	��6l�q�[�]P�n�[͂j�\�GnF�y�H�]ٓl�Jnb&�c���y��p�3L�Y�)��K��z#kU���	Kk�c��Z$�p�h�WzNʋ���{.���J	�0����/zgu7�dt9;l�.<IwN��s�N�g9Wk�Ee�i�w
�=.4���8�m,Z�G_\�1p�z������d��N]�/�>��.�F��r�d���s�1�*J�w4���T�'\���]���*S��p��T��`��8S�/K��,��x�"F��}�����x�~�z������}=~>=z��ǯ^�z�����=z����ׯף�ׯ^�z����=z��ׯ^��sׯ^�z����׏^�z����ׯ_�z�����=z��ׯ��^�|z��ׯ�^�z����ׯ�z����ׯ\��ׯ^�~=�z��ׯ��^��g�^�z�����sׯ^�z��ׯ_oG�^�z�w����{}��o�����{����}�����VN+vJ}�]T�{bv'u�GO�ι�R�'R���F\�{
:��b��w���h�d��ԝ��,%�)���w��Uvm��w��sjOE�΢�7��T�0�\x;X��6�[ʐ -N��op�HYԵl�zj\�V7��4�Z���v\��i��p�:m���(�W'>�Q�u�uՑ�)��ջA	�8���sV�
m�l���	�vE����V %d��Z�n�2����+!�ؐ�����e9B��Ҽe�=P���7&�G*��rھT�IY(򮍞e0kX�QX��
ڝT��������0M��R��;�i�J���L�WK�!�)�Nۓk�e��xp5^VabG��	�2�\X�y�f����v���3���s�û
5�V��eQ4*�b�:9�6����Y髰��TW	Ȥ�sТ{�Z¥p��G]�1�[O�w�1����.��ٶ�>B\�_=C�e$r��K�Wd��O��%�R�Y���+_#�]�ז�	���m���!$�çbsmV�+w��tQ���!)�2ODL�톥����Ğws��9ݚ��#A�֠�kj���!\T���'@��G�>��V]Йao_���ڕ٫2�j�@�O$�z��YNfC�O�����~�_Oׯ������ׯ�z��ׯ^�޽z��ׯ^�}=z���ׯ^�z��ׯ_o^�ׯ^�z������ׯ^�~�g�G�^�z��ׯ׬��ׯ^�z=z��ׯ^�~�|sׯ^�}�z�z��^�z����ׯ^=z��ׯ��^�|z�랽z��ׯ_�=z��ǯ^�z���z����ׯ^�=z��^�~?Y��~���������ׯ]�߾w��<��ŻP�/hD�ڈ�6E���*N�)YB��t�1	�B�ףo2�f�f9u��oA]�c�����������vj���2fm�6�\�;rr�:l�Ԥ=��'	�]���]}����9��$�D�7{f���$B��ҺV�MwF�Fj]��c%r�@��V+3%���$H�u��L:����U�X��	�x̖Z���oҥ�&!9���3�{��_I���)�7�Aũ�-����e�񍱋8���qsF]طj�$4�R�Kp��0j�of�tKUf��Z����nl�Eeo��N*�E����G6��GC7R��Va�w�D򩦲�Wkd�B�.��ytZ5S���V��V�>�:�w^�53�t�sX�q�c��󴰹˖Hè�z^W���wm��<���q�}+���`��e8��z��l�S���N��/+��6���)���$z��e�]�s����v���̾z�pML寇;�9e�z�A�u�][۸2�C�,���MΦ���W;5�/���jǂ�jy�yM�}w{*����v��#�	�����GQ鼗S5V�7I��W]6�c��]��*fZ�� ���^=�:�IP�_>����n��1z5�L6.�Ȁ]��9۬��ު=k1�����dK�CҬ���p����X쫒������;K����^�Q��njK����@}Ɲ�%:7��#ti����+�(2]e��Ri��Z�*.�"R屻ޮ {bd`ٮUY�:�=���=ҥV��ב�}KJSR��b"+��_h;ۏ�+��A�]�s�bW23��]T����MŜ� ����/�J��;k�ɬ��/�����wI���M奃5u��=۳�^���wdo���}Q��r�سy+�c��0X�ѓr6Y�/'�Ю�9��q����mp'�W;���y�m��,b_]�z�$�:6�2��Ֆt�g����qaW�is�y�P��ޖ7Iަ���O�8E���\���8\涭��Ǝ��{N��c�sF�OO �\�����z�c������|2N���UW��-�l���l9h�W:p9lwv@ [l��s�^���'V�+9�R�c@�����끽x����V�J�u��t]��e��e8��Z�&tclb�������
��?x]B�P��J��U���,rwb*9\6�����ZЫ���#����C3�`�f�mT���ܒ�5�A��ޕu`d�B+E��t�\�>��V�xC�&f=�����_2�]N���wXח�e�tb��E�kȑ��1�x���Ů9T�{�oc&mf˵v�Bľ�[ֵ5�žӘt��nd$(n�WG�F�*�=�;��b�z�v#-�:��P�;5�r�
���]�9�Mf
R݀���2.�@k���mʹ�L�\�,�gRf���b��	�dn���ޫC��`�6�3B�#�NoV�{4��]����U<7v=�g[��Nn��gRK���F�?n�p}��?��㫗�K@�E��
=BՃݻ��#��t��Gi���($ni����F�J�U3"Ե�v��x�$�1i��/l��]\�<����Ӗ��ӻc���w�Yե�H��m�ޖY$g0�;�nbi����������u��#��ױN�ږ}��9g3;�S�6! f��k:��8�<�f�*۝m����d�#ɠ��9}����EI��۴�WC�s&Ѷ�߻�es���+ae�mʻ��PxďK�I/z�Ӭ�����׆n���s�	�GsǨX��q�da�U��,��]�ׁDL9ٱ[�'nU!�*�����d����}��v��Ӓ媽�HH��l4��\6��#�� wn���ck:d�)�G:�f�1��Y~���b��]j�ma!v#�ࣅq]������UU�i%N�]Q���D�pm+�@E�0�9�Qw�� ���
�geC�Z��Pi��c���+�N�W
��s
s6�j��=	�u���2�U��I��rw�
Ð�3���3k)c�[�_V�k^�qQ�5ۗ|� ��9N�ma���#zm��j��L˧]���B�9��ں�Bu����b��p��3���0L�3N����g�%�uv���Z�+�v��\7�-�@�.�#o&˭���k�=��ؒ���*o=7�H;�b��f����hvr���A\-7�);�8���.��Ý.�x@���9�v�mՆ#㛻����xC
j/�3i�r���*��[�-����U���(9O*U���!Z4�bƨ��׎Pu��ۖ@�4iĦk��=ٰ�#h��*�unռCgP�{q��otG�l�����]w8��i��z����(SF�J=}c5��K�1N��^V��e1�	u[��脙˝��j���0��[[� 8�M
�4�)��Iz�L/1��YR ��JЊ�,�r��Rv^����e�r�Ulέ��^��*�X�1�%:�@��۹��М�K^�4�K��W8�(i"�e�r��Ӑ�c�"de��M�b�Ԯ~+�
ӎ� �9�Y[�a�U�*s\��o��f�:Ŕ��L�C_k���w���?yO=��������31)y�L�Gh��z� UOZ�t�����\��E�ǘ�]֓�w#�al���YYu�����ule,�j��`9�f�����r�K�X]��)W�������;�i��H��&΁����²Z��ڙ�זx�D��yo,r폷s+t]T��|Zld�<f��Z0���9�քaػ��ӳ���V�������l��ø����[��F�U��
˩��9���K���nѳ'[�o�8Q����5Yz��`�����d7��¥i�%����+*��H�m�*��<��ޅq辢�@�TT[�p�B{��1��%������ >���/rj:�е��,8Gft��U��زӖ�h�*��Ι��%wp�仃��yU���{,ڍ��iWf�C.��H�7%��K�j��/�b�R�w�7JiJ�����O+Mot훩D�f� �����r��2�p���<�
|��čutŹR_uSZ��pEԳøѺ�*�L-�W!1���,�B��2b�d�C,d{�q��SI;�p����3C���	E��G.״+%?("��\]e+�Ǯw(/� Qk�Cz�I��_]:Ь`>z��&a�׶�f�7����wyR��nv��fAǕe�s,��겑.�5��n(;��v���BW6�up��+��:$;%���8gJ�|��ݽ��O�J+��+�]�M�uAט�򛍊�y��i�y-�8.���g/ju�����83:�ۇ|Lf-&E���r2V�u�QF+�/8��>�㛗KGq�<F=�[�n�q�7Y�	µ6o:�[�R5R������we�����u��3]��y��K��s���D�G魖��4�/^��}b��,�	�����-kF�c��l� s�߮�̙�!�:!�UЅ<ݞ�t���:Y���n����L�Q���Dʧ�~�iz5Q�wAܗP�2Pv��5[�����H���ru��\wB�ք��Hɇ �C�e.��U�\;�P��TA��d|�:vkN�F�D8�((�+���$�ǵ-QQ���i�
h<M��W���~e�ِ�������ʩ�t��o(6�o+i[�E�IH9T�U�s9D��t�A�ƭ tu�j��L��YAs���;U`�k�;��[��f�¬g��2�=A��C,��+(p�t�J��Ķ�fI�Y�7^�A�7��4s_0�=N�;ϫ�)G��k�N�3E4OA��B�5�Q��k�]t`��L�[�w˯J�nl�b����ϫQI�5��z�o��p�FdU;J��H��K��oE7FŅ�X���1��Y�L/e
%X∙.�d	P�Ӄ$2�N��"l�ZH�!w:X%�m�Fq��Tk��E�-\]zGگV�]!:x<h��ۺ�]������xX����vVd��Ǳ�:AR ���zҥ��i	��5��6/���n��8la�^ܢ��û�5��%ni�t�V����%n^�.}Q[ݶ�;���p�,��ί_>�'b��r�s�2���ワˮ�8��ĦͫYƤ;w]�6)�{j�Q���U��<�I��3�r)�n.{�㽉������\]#M/MH��'��V���� �1*5��Fp��oz���]IH�	0�7�Ӕ��3j\WJd۴*�I�g	����q�G�Hw��Q��C)������ξ��WB��ù�\�ɹHL�&b69
9�9R}����j+��n�x��;��ۙx�,a0�����,���
�vYܑL�r�Hgp��M�������Ù�̭N�㥹y~X��ny�v��	��c��O��6���(֙e����{{��q��Y�4�[��<��uUV��] �w(���ع*�Q��79��9�nk�Fe(��Q\o0�1��X4�=���\:��ZW��~�'����V�{f���Yr�x�����Z���lw�F�*e�g3 i1vt�Et�,�ɳ�U���+x���He^ԺCtǼ/�5���(ii��ma���%|��F����1V���zZ�4�.��k�������y�y���pç���qGV�2i��I��8K�M �Z6I���nB��Ӆ�c ��܆4���ED�,��4�n��LH1���a�i���R)#$0Ċh�8��dCP�ʈ�<X���$@��!s���0�$�PLRIQ!� b0Pe �-4R�i�S��	L�O6�L�L Z"&Xi&)��MBG�/9<i�w@�Q1����	y�"��aD�Cy�Qm���0	��ԣU!H����a�E�
!�a�E��kֿ����F�Fk�Cj�!�mJ0���V�v�PԲ��,��՜�b��	� !%{��m�].��>��7:�f��V�L����1���,�����i�}U�Z�����w�̳Z�˕�]�Bx�OfZ����ꃩ�o2gVd�F���p��`(�R�"�B���:A�v=60��
��;�rT�iu-<0�a���ʮ�ީ{���K&5~F�U�H�hw���;��2�	��p9��I���-c)S�f��*+��jigB�':�e;l��⵽��x��L���Y��Y�}��)BU8�z��v���\��X��L�B8݇�vUm-�58�'I�v��//'�Kγ{Z%	՗6Ȳ�ܨ8���n��{	��ˏ�s�,8iRTE�}�Y���U���f�;cq�{^q!�p(�Iu�\�=yo�֒!��;�A���ې���������̾�]���::�G[���T�ąy]�n�H��Պ���Wp)����2S��۹�96�5�e�d.�06;��ε�'�8}����ø�;�ui$J&�V�u�wV|�D��gS��ڔN��v���+C�媗�E�����YDM�Z
��v��&IŌp,��ALkͥ#��q�O0��*!!RH1	T��2�2�A�-Yl
M� cA��H�������'
F��0�L�F8d0a��(�4RT�l��l��W�DdM�ĤM�$1��B\a2"�y�KiH�i�L�@�e�E@De�c��~eO#	(����P�"�7䁅�~N8R"K�UA�1�I��$H���Q��&F[!!9$&�I"�L�p������2S�䔘�N$m���J~!D���2���p�IN&��a4dHȜ �8�%�1��0��!�!�ϓ��l�#E�J`��I8"����4�"�P�"@��M��&"�L�L@���e�
��RB2c$��O��H|�/�Fc��> �U@X)�yH�r�c%4[FHDL4cF&B	�c�0XJ#��Ѝ�0B�$�$A�� 5&�*<K� �6��&a�+�� ��,E�bf���kM�IZ��4:S��h�`�0珏���������=z���۱m��PS�F6M�kAMF\�)�sr��NX�s�<�b(�I��j5��s�ǯ_�ǯY��{��*�6)� [�İk�ܩ��,T�,Q�a(��*���9���~�8s�/O�p����~>>?O���~�����~bOל5�SE���&���x^N�8諘(=��rK͔�cͺ{�W9�`�1��ǘ�3�|ysv����q#FN��"Ǘ�U�cͷ�@�V�p�W
4����������#G�8�Q�qD�H�nd[^FW�\������^��<ǅ�T�F 1���l�1P�f��kX�nn\�J��Ǜ�N�'Ta#F��mnFw-�y��y�s���p.X�p�l7���0���?s����\��.X�;b�A�y��A�Z�ܞV)5�9͒|�4���9�#��F9������Ip9��8�i����8��p9͹Ø�9Y�\��y��jOZ�Ɲs���61��l\���a���p���'r��3n\��sVܽy�
"��n5q���fy#��� ۄ����ሴhլ��ۙ��^p�g�<�N�lr�9�<��95��.Ac�4��^y�\�#my��\�)��M<������ʪ�\����yiJ#xn1��/��;�x�:�G�܃�$���щ(/���y�=xy*��#�"�����Z!�
A�@LC)(Y��1�[�s>sy�9�o
ܹ����K�ޓf�_J�3��'��B��A"F�V��3������M�Ր���'1]=� �5N���H2m2BD��(�B$!2 �,�!�z0�^FZLD�>��`�ZD�!p([$¢F X�CP�,5d�Io�q%l�bsG� ��T�Ct1��m�~$1d Aj��f��¬f�P�'�O-e�U�~����ܡq��r ��"dǳ���U�_z?O?���y����铰n���M���_��]��gЙ����n���E��m�x��#�$Ȼ�G��|@V��ؠ(���9���g@���3�y�}�1^^XKصt�^��{����9�����V�zj�wCj��^U��Q׻t`;3����1�j�cؼ���Wx��!s����u]�?oz��*��^�V{�r��c{U���:t��k�: ,��c5���f�����q��Vck"�{��Lc�D	���h���{z(��@�q��ɏ�:�b��.ͽ��̿zN=����
�*���}��\w���v�w����<�v/Qm�K�\*�%zq���|}]^y{�Di��}d��֙�k�L�aK�|��xo�|�=ӱ4JU�Xt���^ׯy�t����WH᎚{�+��l�bu���c�$�U�o������N�Wv���f��G�:�{��2�A~�����6�5Jm�։��F��j�v��5�#�?���rI�6ws������k���E�����?5����-�۬ n�=���{4�rW78WvU��_@q�����} X�Z盙��M�_dJI��!���t*��=]�f����ЧG���]������l�ܴ��H��3+�ٍ��7���\p�����l�3�h���KCΝ���*�6�s3��=��b�-�����t�C�q���h�ׂ{W_��z'^�E_u����0�}�>���3^�0��Cй����&�~y��; .�)��~�V�Zj���sS�����.�y�egsY�^+F7fi����]��z�����L߉7U�qG�m{�����B��<�bH_y������vI��nG��M��1���i��rd��d�=��{;<9Ws�ڜ�hg��w��������r�j�H�����#�G�S��� ݆.o7�w������)���oL&���nº�
�:�nT�����a^�>��n u��u�ت�D�> �>++D�;���ԕ�]�.�פu�c���x���}I_3�w�f^�o�y�{p�Fu���}L;a��d���\;{�ύ�5
��g�I���޼S��4�gfލխZ����Jw6��,}�>����Ƅ�
�>���/�(?5"A����v8�����XY'��T�W�I�=;��(�4��罐ȣ�{��9�+;�/Uen���v���nd�fDob�ţ��&8��sÿ;@Y
m��_�����on|)��O��/+��Ϣ��F�%�xj6+�ߨd.�����7y���;��\~�U���ހw%�p�p��J�� >��>�w������U���O�t��rxs9��A����>�U�kuc88Bm�|��C=J��j��T���8����7$��T�G&n�A��l&�|�˹���<UBm���^�T�.0)�}������W�z�z��ܚ"���Y�xa��V��T�܅N�N��Ʊ6�lU��-�d9g�m�tlɹ��sP�t��A�~[�va�x�*�<Y��.T�`����]/���`j:�x��J��	3מ����=�����K���,I]�3�R��B���-�0�ʋ+\{��f�]�-���E:8FO����˵��$������~f�S�81�i(�o�n����$����	��=�2qżH��F�ϯ��c�~峺�m��t��б+�_C�8�����<��|��E^kw�YW<x���C��\��S~���=������*����]�N����|7��F�o�*�M������r߇W��.���^�LONᾑ��-}�_L�����}�G�M6�5X��w�Ω6�{u��{�,��P��ۭo}�~'_���>��_y|${���=��g�
nM���Y`{7��&��SW�f����:ە�l��c�ϼ����n�)��"�?���5�x�k��{���{��)�?y�}]�졂��nf1��3��w��"��Ͻ�O5W�Z=/{�����q!~U�cAY�t�Z��F����wA�w2�H�]uWV�W-QFX�n��	'n���ωU��o�oc3b�]u�����c��wh��Z�e˾s�>��}]����)-Nt��S��>ʞF_sͨ��3Z��]���! :�U_Fj�?"B/t����|3Ԏ�D�2
�!�ߓ~qz���D�w�u��Yg?��*wG������J�UwN_�W`d!�.+��ҭ*z��]��)�:�ƸTwb�_����֩�����h9�ʐs���o�ןq��W��>��z*��nj���SL��=����xwt��Z����]X��X��~����g��^2_C�U���2���9�7}�A|{��Ԝ�ï��ݶh��Ʃ�������͉k"�ž�p �v^����<K����rA㕛w�5C99��𼞠����#�x�g�Țw���S���;kݒv�تזf�b:�`�ro��fj����Xn��f�{DOuO��ݲ���,c/��"��j^���b�`e݋ﻸ����.��TU�!�>+h{�uo+)�{��a���`-�+�|C;�0�έ�>�y��Ի٦`2��]y����
]��K�7��Bu��A�d�;v��7v�vT���{�[5�l/��{x���%|<�1t�˷��[#Y*f*���<}�*�2��r|
|.�ZKj�]uE.M$!�)}�j](��+��;u�ϲ<;äzֻ�gegT�0�L8i�u�U�!^*л��H�ϵ��X瓔�H$��2:gd7�DL�A���U�l��{�~�"�@��}�����Ӈ���7���C~�'���֕��o0��9��K`��Z{d<@2�6f0=۴};h�{�.����g�B���cGW1<�����/e�����v�O �Lk��YĄ�0woz�����ݘ�����$����9~�� W�m�
��Kz�r��d�~����霚�><n}]�s�����˲�1~��r��ߍm`; �~�TL	�a����My�mΑ��9�7Pj�;?[���:m�޴F�U��bP���Ū���m쑽�k=�����T�kq3�<��]I�٦z���鵚�O�!�eN��Ru=]��l}@g� ���I]�S����0?{mM���9�q��l�]p1#��z�1�5G��"�[W�@���6�{N�n�Mgd $��ѽ�P�u�7f=U�����D����A�����Q�ˎNR��܂AA�}��m����7T�5���=��'e)��wmh�5޼�\��}���}_`s�NǙ�lhz3c>��T_m�[����ve{3�>/��kS������D�h=@q��'2����ܫ'>�+Dӵ�h�f4����}@u"��S'>y�Խ�K~�$}�N�i�i�k�¦F�^W�!��:4[��@�23�ǤlO�	��ۃ8A�����<e�T����]�L���wr���_��<�S�z�-���ӏ�k����"�+i��Ͻ�z�=�����[V�+_�Dpا1��h���^��@b��=���4����V�elޞ9��EE�Na�3g#���h^�X��/A����UO�{������͋�\���Ko��wv��hzv�?q݊�̻� �9(���c��-��s��&5��1u�'��0fֆ�_I]�l�^�g�:L3�=�:z�;�+�j�iw�*���p�)�ڰ���v�����L\h[_ᕵKNW'�L]�i�j�1g��C35i�N��=w'M�]�S�H����a�QM�I�z7���[ӹ/����n�eѽ�˔#����
O�3a3��0���^f�xzjgov��{������H�Y�b�9:��:-���W7ڦ�F��d]��h���*݊<+���K�/}"��_Yi�dD�W����������`�� 
=�vqǼÜc����y*���5;���<zi��쩸�_Kj*�w��}�n|4q���cʳ�q{��\��E�N��39~f���-O^���Nþ�_�lU�k����\�`�Xô���w��cB>����]r-��mrӄ�x{$��,vC]�:s�宦�qF�a��<�ށO�u���'h�iy�}�ϡ�s�J�5Q����I��B��7��gj��z�L�����������Jj��Qfl�:w�9�����Y-�Pc����z������Oa����=��P�����H��4�iC��ٹo��7g�=]��NMl��m[�=�g&U�R��.�m'ZN�T�+��#iZ�7�1u��vE���6	i�R�I&4e�o5��0*�we��U��+��Z윲68T�rv>WY��L��^�C�U&z��03q�b%����vD�_}�����`B�#w�r�\�v �
�0R��	4��6�E���A��F_#�z��K�}�y_x �����Y��joVWyl��J�>�����3���#�{�f%�3ǣ,p�B��л/�P}��x�\����=B@׬��9E���}">�g����LQu� |9�/���z�h\��K�3����->���|�������=�ϧNޜ=�Ɗ�d�8�m-l0���Rz`�6uϳz��.�q�����'��&^�욶��_�?x�M��~�(V�.�b�'��5O��L�6i����>n��{��3ä1�l[���.���6��q{���Y������;�G���6x�k��;i`>���vN+��z��)��VU�̮���T�>t��*z���s�r��k�#��C_c��]���3�y��5V��/�� �	���U|��9$��Ǘ�3��<a�Gٜ��z����4��7�\��P[����{ec���h�N�"RT����#!�,d*m���&ut~ֱ�_ԥ�c^�|��-��WT÷!�Guͽ����4��ELsFBS�ٗ�.��(�̄�Ȧ��#qr<D�ī�CU@���fv,ͱ����'-q��;]�=�4��Þ�:y�����û�{�&3����IVh�Od�P�9���-tǞ��5��4�ȝ�8z��s�M��XR��B����z���E������+�O5��^7wc�v�n�&�@+����"��o���<�Tsƺ>�-�i��&�_�\wCwM��9���{�󆧈�/vRү%_Ҧ�'�{�w/O�y߁92��	������OK�?)B#^� ��Ow\x�]�g��k��w�M�}�[������7�;+{h/���դ-Yҷ��|���WN��)���c�
#kg �����A���[�=�=�f������\��s�^�Eڷ�{�0��VPH��ѫ{�}������ks���W6�������b���xx�.�}�2K�`��珥���7��.f��l�V�hР�.�:&�Y�Qt-֝�h���B�]�a�b�����
����S]��@�Q�WYӪ��͙�{�#�t,�s����}nuqZǽF�Ь/|,u�=ܕ�W[��6S��S�;<��I��nI�d���y�}B���k2eu�1OS�U׽YZ�\%����Z��b��ve�Wj�=�R�8˫��̽�v���}}zb�N����U�b�m[7�"w|޷��A}�כ3Q���x�������P�XuC�Xa��:��	nƥ�	����w�Y��U[ȫ�|�ٶ��8�����u�2�]݀m�7ʡ�����g
S�+1���9�� ��}��M�-�M��(l/T��Xs��)/�,���B�����B\NuջC��J�:ub8k�^�j�dΉ(nC�D��5�l,�'&�۸9i�2Wf{j�yG�z�&K�$�N�V�Ɣ!��1��E�=O`H���ֺ�Y�7�B��՚��l޸�B�JC�雷+K��ӗnч���`9�T5b-̗�s4�-��f(vQ�|{35��uQ�������3������gy`�4����"��������F�fj��4���ǏV1	��V�W��������\���s'B��j�u| ^�����W�##�1
hZ�Z��@��P>"�{�"���]h�1X�D�G~��J����g$cd�]-a���+�ri�7���vEU���p�ֽ���V�P��*'�7sl��E͊�L�q���t�]�]C��R�,�j�|oH	��v<�r��ʪ�qWU��غǋ���c`�ÅIYh�UO��2r��N7S
��C{pw*��g[��:=�
�`��L�J��]�5�zn!�w���f�\�M�BKQ��m�)11�pE�t���u����q;p�ۄ��0S�V�K�T0-<9�i��guf�E���q�g���Yvc-t̴�`���˳�F¶��mf�t<�fU��6i;XIqK�=�k�i̗���4K  Y��RB�D��{\�̙���<�ut�w��3+��a�8N�C�
���9�+�;�;$.y7��jя�!�#��U��-ʍ�'a9�uz��@8��YԮ��l-Ǎ��y��~y��|t���B9�w#�^��S
��˴+�egQ�����^���nJ�qu7���[m��
��FL{אn8�CN�2Vm�]-���u�ۿhƻ���;kw�B�Ʀ� gQ��������kWffԷ۰�kB��r�oT�[}a��Jͤ���ҝ��ͮ��֔A+��up�},��w-�W�����j䏻6�X"I�f$$�|H�b��:kCG�h�9����j6�����U<����U�:�g�����������~������~�"��*�)*�c��1EUlV�*��*+N*�j�N�A�J彾3�3����}>>>>?�����f~�h�[�M�E{<��/+FִSF�	��ƫTUIl�p����Ϗ���~>�����9�O��ڂ-��Tm��LN6�Vƶ��6�X�ּ?y�y���h(���gV��TW�Đs��8�Lxl�؍c���S��?m��c��)�j5�Z�j"48���95s��L�h �$�#��&*���.Qr3�P˗v��)1Uy�LQ�cՒ�QQ�F��y�^UPy��>΋��tDαkya���i��gLm���\Ƶ6�to�ܪZmf
����b������b��&#�cU�[h�F���c���r0kPVض�RZ6�5������V�n�7	�*�m�TU����E�N�
���"�6��Śsv9r�)�[�8�
(��cLEkA�v؂�)ă�Ix�I>�7/u��ϱ�ع�2�	��l���6#�]^]�`���^�7Kh����G�m�M��MΣ����2C,3�9z�y﷿��۞`�4���6�<��ַ�	�Y������;�`���uzFw-2oo�|sy���՟.�
�nr�C!5s�3�[ �f�C�n��������8��6\=7@:xv�d�j�.���^�I��Ʀ�d�N3���`}�;�4^�'���;��#2�mq�al����YIa��ZW�����~D/������П��1EZ��u�Ͱ�	Oy��f�i��Z[��_۱J�~�@ma�ަ[����'c"̀b�Ic��5��[����D]	����'�]�@<tK͈{T@�~�^J81j��dڲ ���YE��N;�H�0�Ƚy�3��\���N.���":cqѯ�G��xc�Fϵ��oE+� ��ʢ���M�%VK�w���6�/[�����<��:i�����J-������[9�v˯A��js�4tI��S�I����&��[I��|W�bxI!�{���ޒ�F��+g͞0���zf���v�Q������d�n�T:�w]͂�f���E�� �T�f�; ��/��}K���"�i��WtF_}%���E�U�&�xy�L޼i��KD����I5���W���y�;o(=�ʴ������չXb4-pCU�4�y՟L՛W��W��Z|���+�ߕd��l���v+��ý�VKn�9l3f�2:�U�S:��E�+4��v��]�ӽ3߇����9�����1���v�m��xLwo@����`���dS�߬
�����\�5�\s�×���d�C�u���}xb	���<z�x`/�fy���ύ�@I�oSW��\��!��������{�����~�@��(�}G������l�����?g��v=,�I�`0�S��#�K	���ޔp^~�?x9���-({������`
�^cL��͐
q�H�E��RkZA1M�w-F=n����Mʙf�!vf�|^��3�.��y1j��uC#|���h~ۯ�|LsxeA�.2bέ̋��6��׃������~	y�-G�F�h
�8/��!>�x��Cvy�;8}K_~IZj���s7�5Y�gBqـ���s-vW +�K~����~A�O��D���d+�HN�ݫ*��򽿺�q��p�2���zZ���v~�6ކU��~q�}�y_�-���FS��,�����z���oz6��`�@@&�bP4
ܝe�&�6h㞡Lk֮��# [�4�C㚃#�!�H�:��OZ�'�913=e���1��N�b�¹ռ�fmɀ�z9�o�mxV�F��2w]��������¢ٷnMWN��:����R�M���65:.ٖ?)�;���(�ے�-�>3��B�IE�Z>�n���۪=���D���D�� ���g�p$1ΟN6�x��Db�Z���U�c���rp�2U�Ev	�'o]�b�ɻeֽ�T��ܶ�>�x����J�AB�n��V~�/𱤊5p�d6~,ƌr8���i$��@8��*r�\��^~Pdgڀ��~:�Ι7��<�������S���oSDF�/
�tl7=� ��v�@.�c�퇯M�3�O�LY��N �;��淈M��m�>\�2��Lo,��͡�����J�ZU��'���}���𢣙�C�pm��h���s{c��܍ѳ�����z�c[�ܙ厾��g�{���56b �_�-��g�`�R�oB\���^�<���R�YUt��v�w(xL�~hIIa�`n/��Je�� sjP�å�]̒.aa������d�/�� fq���g�¨Y�.(Y�@s�\� k��j �����6�p��\t�1�3�u�����jb1��fy1��tz��ݘ߄\���oP����q�����u�uڶ�nc����Ws�xl��(�
1�`�?s���TS)����ԫ�/�@�o=�1�qۏ������i@v-��'�Q���Z�r ����x�E�aQ��@��}n>?�O������7�;V}̯�=7�v�g5�� w[��z@V���� ��b���6���@t��;8^���P�,5�oC7u�U=�K,�k퓳{���n��T#�i=g����̪#E=Ť���D�#����ܣw1�fԫ<M:�0�ȷ��䢫������M�c��o�G7�ۓ���Н��nm�Xଉ���)�P��QNŴ��b����2�oX������a�nj�[w���#�Ks!����z|4����hO��S��wT�	g�T"=��,"eN���[�9T�zsv�Mm��u!�)CU:N�� ]�F�r~ks sm���b��1���t����-�S��^&a���o�S�ź����x!g T�[x��8Qw>ێ���Fy�hq/Sz*��n�����s���dP V$~�7����;`}�D8�(@��S
��2`"@&BeIexV:�J��qS�s
��^ >7��/n^iw�f��߼�c_�ĵ��8*nG�@0����p"��X[-P:�>lnohQ�{�ny�׫��=�~ˡU�e&�����Y���5��s�u�	���y�(�[�EBi�*]�>ύ_g� 7	>>$��������s{�D�k���,�m��
z������4��D�\�츎Ӷ;��GGt{���ǂ������d�1T�݃��P�/��~�����2d��ٔ��iS�3s��� ���G�Jl���;؍w�,F�a���@�Zʎm�%+e.��:�p��ˈK�u�R�)��ޏ	%��i9l�����gl�M���|��Uqp�2����w�J��x4�0~��}gh��9�Ԇ���M��-o\�Ȃ��)�����Ç�9����a?ZGT�o���J����]��r`�A�7j���o�b�5�r�+��`��9�\���*A��Uٗʶ�go[��1�@�W���)�������x��=��0�1Gޚzjd���1q��s��w��� ���R����W�N+�l||��UYy:��ǅ�꧆��B  �Pe`�3`	����"����@E�&�/-�>����:1󟧳#k����^����[�:S����5��<cZ}f|�H��� ��X	{o�à?�&@�s^���W�2�*�� mxcμ�~`W�o,�cа'?aרN~}����'y"@�ψ߿D�����n5�>����r<��>F�nN0
���扈�[O�`����z8�\��a�0�Y#e�!c�Z/�ϐ|�
p�L����b�;60����8�M��H�)H\q������No���{�}_�+?��o� ߧ��0,���拫�`'x˲.p�9�Ԛ'4�wE3����e�6���Y����E�=�+��h�>�x�j�=+�茀}�nd��s�p���j9�3/et6���0�D�����oo�PF1�$�p3��Õ>�Z��4�h�z:���4,�f�(�Tu���[�r%��d�f�>��f��:(�)�����0��-~���WL�Δ�e轛V.��nq���z��0O�[S�$�ǽ�$�B6SV,���b���Us����+�C�0р��s���������vrT�f���S"�L��O\��ke囦��#":fAxV�i��^L�qΝ��G.5A�}����� �۴��ڃ}���<>j݁��~�����=��O����(%9�v����>���Yb�P���md�lJ:���<��6���wjn�`o��;�h�K�N�x�T/M��ݽFw��"�$�{2j�d3��sN=+�1��9��̟s� c5�jħX
��H�b]�8�c\�F�S�6ADD�]8�A��] �;�W���~�(�n���|��q��:���0�n�osR�?��+$��~%�*�]?5�a�.�����,?��=hNEfq��Km����᜚n.�d�&�k��Bd�t�Js>�hE67����� ;���:�1����zpf�b�z����tn����_)ޭQ�2���_�7�~��}[�ߧ��͡�[<��S&��1F�h��O���w�~j��I�)aʅ{�8�="۬�ʓZ�LL��h:�)җe,(Q�Zx����'rc_$O���� H*}��{ﺰ���P�2'z<i�q����k���Ӗ�n��o�%Ϫ�r/�E��ȝ��� ����h�,�|��������uU]��l
ٶ\3 �w���ZOn,5�T���]��Sλ7��a�d�U�Kk�-t�e<A�W�������}Y7o�o��
��ݾ|�s�+�w�1n.��9�iU\�2𻹬\�#	���Y�P�x��/gA�?��#����#�{t�)�2�L���-_��,�H���`��� ��P�L�J��x���l�����$�9�gO@��駁��DB�a~��nOc<Ҳ�y�'3��ʭ���1�I�;"��\�t��U�n1P�;=>}QAK����>�k�Ä�=���!�p��Mv�c �<:oe�+ ��E�l��D����|Fm�OL>9��f�Od4q�ST�\����	B"����F���dcu
�0��cIe
�ӌ%��/�5�]x�M��fZ��F�Zv(3�l��G��:���
y��ӯ	��ٰ��ߎ������-�.~|�I�r��=R��\���c%�,�vF�-�Qm>��.(�Tc&�07`�l���X���6�S����T��j	qa��U�y���~�li��c=	�d,�f��V\��v�6���:�w�=~�ޛe���t���`��b�T�q���
�[��k�~��un�5��'�_bA�C����E�g���"�?���E�?6%�u�'��-������� tg\��k�K��λZ��z`k.|h/^�FG c���S�7�m�h�:9�QM�]�����\B~*���۫��0eM��j#��~���n��~��<�M<K�Jh�OWum�_��*��7Q���U�?z4)�N뒡*�"{��&�\��f�̮����wzoz&+�w��.��
|�|,����9F�ԚE���"���f��ܐսN<�װ�O��X���x������A�����&�7�1ʹ&!8�DA�R���&ŧ���zc��ZRX\�=G���2���8\�F���d�bg�L�1���3����]m��0K�_��!x�����Uʔ��h��guߨq���.�̿x���@J��&���>5��d�
1�lLd9��Ւ�H�Y1p�\qr����ș���������vׇFD�60�3'�u����Rz3Fn¨}G�ٟ~�i䅯,��*��A��r���� ܳ��Ȗ�s@dy�"S)�d_U���|�D{pf�K��lq ]ô��Z����$X���4�6Ξ�F�����/���K��3~�pmB ��
�y����*z_��!:\���g���0�ux�s�m�:��`��V�·swL��O��F����M�/>��"���)�Y�SEg�6�J���35�db�W۝��g?�K^D��MOr�����1w�f���C�`��?/�z��8.����n#���55�"Ym�����XU�b��O =�2��;ݼ�C5������4������m�V����{�SlA�L�S���i�ٌon��-7����	�h���1�*| ����<GNǏ4UvN�W��<�t����1Y�8q���I=��p1+����	[%S"�l�%-�V�)���0��F�+����9�:KZ*Z�,�tG1ϒ�e�}�m�TS��`u�:��p�jEУ��i��g[,S����	�wC;dH�^�P:h�a�#t��SM��0i�l��\M����8��.v�L�0ֱ�G.]��鶜sm�0�CT�q�c������'�ġ[�V�!��u�Ź�;� ̑�WA��=1��%Ck�;)��S�^aG�R�׶�> �-�z�7d��Ж���܋��.�A�W�����<����?�>��`����L�ͩ�Kg�η@�r�e-~{G��Ɯ��+P���B�Щ��Y�׻̶�/R�Wƽ:J�/2��^}��������)-�25�U��5q�`3�T�H�`���1�zXfi�4����K�l�E��G�<�n��]��;�H�݈6�]��i��=��{�!���3[�wf�*"�*}f�L��w�nE����^�t_S��� �) 6��c�����l�6�N������lŦ��,��ݒ�P��/<3d��!\����f�ٕ�ݳCm�m��Aawx���˺t�&|>��%U����"��q'vF�$(��G������x��S��h�`���=&U�K�
�dI��r�����Eqc\��r;$�ǝ��c��'c��P�-m��\�tݻxx�!�]R�vF���{G�������K���a������C�'�!R�4����ǡ�%� �9�w������OO�`l�4z���y�݉KK_V��3ʳ��
�?;���~�*�N�<���V��E�	���E0�R/4�{�v�[�u�ڋ��c�8`�|��d��֙L��
�K0AvT0�#}4۾c�g���"� KVm��@Uq�MpswX���@�P"�%[�?,m�	mSm��^;���ݩ+��^�W�٠$�C};̪���G �a�ۂ��gk�XgXߨ�L����F������%X�׺j̘�Wz�56��֢�<�#�i��5K���4�&�q�Qu�7[B� �P9�U�I�&��8�qJXE\䷞�c� 3������O��6W��V�
���b�=]$�b��pɘ���m��ۃ0οjhkO������;hދ�FTc����Zm�Wt;@��mq�0��moV�����VƠ���!��F�61�����5ݼ�-��Hꗅ��P�չ�.��u��f�CÒ�KO��{���2jK��~���>��dI"�����a�~����qzIЬ1A�f_gD\e��y�}��|ڛݹ�9<�V�蝣���h�Y����3t����+�r��c[��`u�f��_F���UU�ܼ�v��Q�.���9���U�CUF�ɺ�D+r���ǩѩ���k>ǖ�^}z����x��D<�/c��n��\)��yk2�	m�;OQ.$.�j�{#q���p�>�"�Wp�Rz�u�{u��睃���:Ƽ�/	Ǜn��U'c�(�yޛ���z��,l�6�آ�����X�x9�t�3�ϴoC�����:�7B��Y�U�fu���,�{7e�� K�
��#�^�AB��Z�V`e��wӳNqP��ע���������Z��E_�`WsE�������R�������<jc�D�FyB����\ic�4�ц����%���/[=��T�I�@u��h,�c:��=��T����ko����5��������Qb�ޜ��}Ճ��n�o�����&��eT�X���i�v%%Ĵ���3���1.<��,�*�g;��T2Ur1�Skj鞧��c��X.�mE�!���x����U�h��&*Y��f�7:�a��ޭ]ਫ਼���͈��DmWD�� :���u�5f�\�aM7@&F�Ox`G۳�ы�+����(�����}���%���ի��d=�Ӫ�rSӈť��2��Ӭ�Aنa��V=�b��H7�;DKOM���x�����ʺ���Wn+*�K`�.%.��"�t���I�P �Ecb�Q�ڮ��
y;�X$��E�b�n��9��]�K�=����R@���
R`��UP�1o�P� �m �T��g�r�(1G+z��Oj�leY��\B����c���	��3�w��Ͱ�C8�]�lS�{'d�
2k3Zs2�CUO���Z�h����Z��/D����s��Bb5v��As�>6�؉�2��6�]"ډղ�6e��6q���p�V��u��)|^ku+z�Awڗq�G^9���,�V�'�_�c��Jݬ���d#�\Ͱ]qS��E�$����Y'��6���w
Vi��Ϋ{��z��*�R��Z�������E6F������8�f4������ҧ}�8j��4�l��򾅩��B7ǝ�Z>l����Ur�1>3=�,3��Y��fl���g(��R�c}�U����fo���Z�F ���US�t���j��Ų�h��_;�g�����;.�J��}�i����r��٘�IT«�vZqv<Uhz�P���m�j�}Pk=o�k
����h�{[Zᶴ֞f��x�XN���ˊY�,��!OY�o����yÕllo�m�+��ܹ;���Y�@�ϝ�ZOW&+��`��;��� mr�d�G�үo]�A3mC�)���k�^�+��bp��ѽ��,�$��8����%ۅ�n�R��Ad�{\-.�B�QL���t�A>"!�����mW1��k5kEz�?xnj-b��������c��g<g����������?_�g�bj��2E1-[;[gD[5%SDA�����d�"���;V�ZZ-�4�3�<s����}>>>>=�_�g�*��ű�9���5s1U��s�bѧDTc8����ϜEM�}3���>�O�����||~���3�_�ݢ���t�mQ6�ECF�DSlX��Cl�|g�|�&�d�j61AQ��;nX�*Z��kSi-��b�1�����jO�f�j����0EAr܋f������:��Z֛gA��Zr킱�E��UWͯ6��c%AAM+0TIQj�:��Pp���k��EE#MV����Ql��m�[lUCF٬E�m��ccb���`�֐�rnq8�P\j4h��p�M[-����^4TQO	��#mڙ�����Y6�D`Q�
;B6�l��&���KP��@ˑ�HB� �F#1#=E5�W��gp��x[9X�޷w���ܩj'J�V,����SX��jt?t���vW-ר�η\*5�tn�V�X�m��f��$�6ш��nF�M@�a�� �0L0�$j!�Aю(���"���`)�D�1�Z~N(D��*(k�����煯� �C"0� �dP�J�׭lk����DC�ߏ�"����I�ϛ~n$��D(IM���׋��R�1干��[z���+��^ׄ��>�K�f�0�����v]r �;L��=и�f"̚�4y���C�1�<ƙ����E8�
��:�0:Us>�
�f��{�]��ܾ�S�*���A��X�_�.퀸�uo�p<���i��t�
ރo��w���Ͼ5�>�3�ұ�5��D��0u5����*/��ٿ"z�y�vla�Z���URΫQ���� ��$Xb�`sΝ���}:�5��f��H�踶��]:ɥ]�G����!��-�fYq���ͯC��f�tG)�u]mP��:0�8�ܒEu���:��g�u/V�ڮ�)�.���L��#҃?0��`.=#UK�ϑ�w��1ڜ�F���K���" �����OL r�o^��C���k$M�]X�{g6��Q�`ɓ�V��i��$Wҗ��g�a�
�^�o��n�;�(��iׄ�SP���r_=[�U�cFQk����9=Z�L�\�����}�N��#ݾ.z׶�(��4|�>x��6迳X�����n�Υ���6�LwgZ�蠇�U����t񗈘�����H����"��z//w�FK���ĒUŏ�w�����Q4��k:G�@�7(ge�JJ'5��Z 8P���9go47Ę�%V�]d�i���v	5n�xx��}N] �a�D�J�I� � �0 OE�:h¬������&�ؼz����\=5��Kg��@�Y�fvI�F@!����Hi0ژ��E�yyA�zҕ/G�T��TSg?%�Vr�ߍM�EB�@��"�����_�a�w0����߶�x�Љ�Ӯ���ΐ�S��\��l^\��XP�ך���"2+�ttU�Z�;�D��ⴊB1���L��FD��qqƔ�(�ds�g�bzmm-��̚G��nD�wa�5G2��.$Dt��nZ4*��O�?͋��r�/�����|5�:m�f�0A�LY�V��� �翕H���?[�ˁ%�[�b��xj�)�����)�h�x�#�ъ�(45��[Az/�p��Z���a0��f��sL������
 zK�sv�˙:�N+�a5��o�MH���G�Q ���[B3jy}��uW�3s��'�:F�C�Z�b�fam��~U��{_I��c��J{S(��o��}�s-f�By�u����B��u�J,���%�e�6c�}l~��A�$��4��Y�"};ޮ>���8���g��kxw��YX3i��i���-�)��7�iJ.�{�l��<�Y�jA��8��q{�+>ۆ�!���8��ܵ�c�Ac+��b�K�US�Ԃ��Yq(`�Ո}&W*@�ݭ�޸�͝Z�'b���5���� {�#�a�S$�*��^������筽��ߗ�f�ǄF���)��w��AlB��B������¡!3>�-s��&WU���$�cS�Ǘp�%t�$k�Y�6�%�Y���ߓ߰Tk�ƔC� � �7%a {�T�P��+�3E�:��I����IvQ�6l�ߥ�i��X���S���Ѷ���N�%���fs�嬨��S�+�ԛ�@��~[����˟��@w���}/|dB�=�>�H���Fm�[���quJ�r!0��]�T�|D�T[n+�`\�����5�v\(i�}S��˴iN�ځ1��C�[#S�}~�.��m���u��m��m�<�^p�c%�Iĺ�cաCc)[.�D�W4��E{T��6x�͚�O��)�n�k{x���jW�xT
���咨ٹA�*�z���gd����S�u(��z�D���r.�|��^���M�q��@6���75�s�F���\�ߧ��)�WN�e�-H�Vh�*��4��M�<r5s�_���Ӑ�(hT�f�f�ׁ���g��1�Κ��þ;�r̆1#FTû���a�o)�s�����#[߉�;�^ȕ��w�S�:,����S,k&�D!���w���^���irS��Z�i(��G{��+�5X���9���P��;;U�Rpk����Ҡ0�]&�|���é�Я�2��2�BJT�߻���w��?��>���?]g7�gt����u^��Lü̼L�_���*���8z�g�z��ڨ@�!�I�Ŝ�ڣK�"��_li�9=�tz�}��:}������lt������继��4��v�q�Xn��oa%��^c���n��1��|��t���o5w�Z�&I{�Y����� M�Z㫟�z�v(�k�xf�\;H���p���a̟X�9Cl7o����`5����>]/s�n��,}������C�KL�L�Qo� ����v{�=�ݴm���eA�ᔃTU�a��5s���B�
��3�~��~�_*�K~(>G�;�&�����}-��l;�{O�81�����'�&P�蘖�]�%���zw��"%��i��*FO6lJ뗽Zѹ��9Er�(����F�j̄� r%�e�W]�b�!dۼ4�5�r��I�"���1OM�Ŭ ��Hw�w�Utj�ށ�9�c��&\�ؤ����oOl���ohLQ�|�ۺ�vAt;��>����	K��߃)��8�+����G�ӴB�����fe��k8�����V�1�Hٔ+�T0}Y��xQF]�~��˽�������Q�����?k@�{��N�i��*���z�T鹚��#˓8�*��ůS��t&F��s��i�r��F4;}��������w�O�`D�DHe��H'��v�-�1�\�_~?~����0���$�$���p�c
%<�Z(�Q'�
���L�D[�}�����J�_��'ڸ�h����T���xܛ��-o�w���{90�E[�Ҭ��WA�g�t�� 撚|���,����ad|uK�;1��Oĉ��t�JEz�n��u�kǒ�i����b�F5)�֑������f��.2U�yY�kk�%;M �O"�	j/��/�S&�����s>�hE6k㻳5��n!Zi�oH�K��R���xh.���'��:�³ת���̝gO^9�����t}W�5���f<?���#��_R;N���b��,�6@he���I�Ǥ���#sa'v�vGF�O��W|{�5%~�����t�N@_J�w^�lz�8e��.<�Fb��#NH��"떪�]*E� ��d��Gc�e���W�r�9�� �R��[�|�C�R.�9�vc7�l8k-ڶ:�s��b����͒2�DKm1�-;�S�t�7=3�^/.�h<h�DL��e�v_��u}Ðj�P�NG󈪗lb\b�,����
��*ft��D�zwDj�J[��#�n�f�_oN��[eMSt��6&���?�Bx~9l26o#�	�j��T%��IY�k�g;��Gܕ�d��s��'�	 ��?�Y�?�w�SRC7�>ީ���\����A�����:��ޅo]�]������x�� 0��p���@�E=5�g��\G�*=Kո��w�P��5��ՆD��w|Fm�nh��tn�k�oj�,�i˗bc�)��@�%��j��J��~��!�9[ڕ�4��<M⟊���6�F��^WN���|�^mS��|���0�ʾ]q�������?�]ƹ���]rJ��tUR<�r�|ff}��q��]��'א�Oލ���r\&,�Jq�B�,Ɯ0iW�]y:F����3�M��.=�^$y��a����q-�dd���,�m���-�v�tM��(2@f�y�����S.~ħ�*�X�+y�\Q+5�>��lϝ��. �>��|t��*w��L$��N�/0�ƶ�k�P��ٻ�T���n[���wj:"팗@<@��8��No<��y�������U�
0YstkZG��m��_������?{�6��<n��F��ބ��\{�Z�ޯj�.*�˧���8fU{sw74��ɚ1�)2XH:�34m�&f���Ń4��/Bf5=	ye1���Zn5����M�Y�&0���2�[��f=�Cܺ�@�ԡ�F��f�+YֵW�G��)�y}ҳ:�`�H9��#��}�f��sm؝�d�f�N��N�5���m|�w@I'Z+����*B�\\)Qx������O����ϗ����=�ZC�e!S�:�@��9gQ��W�2_"��j�M�֑ߝ����M	�,.� ���'�T���O����cU��^L��ͧUH���(֗;<�y�N�3͐�&d"�@fҠh�k��v_rɅs����������Dm|D³��xs��p���/�����iL��ܳy�u��b���G�w�^��ǟb�/5d��5뤜F�/�c�=4۳fd~mܶ�#�QL�x�N�&��~��ӳ�N��m�0��6܄���^S�.��-��>k�\edc۹ێX�瑄�fޚ���3�f��xM˩��{KH)�t��4:�;T�9_�4��d�z������ЕS0��η
�NTV����f�M	\�ȫ�6��^	����1_�6�d�Ί!�'�w��B��K&Y�)om5�4̽̂�4ُ�f�6��	�obK2��ۧ�ю̹ٮ��魙f����6�F
[Bj�cMJ�z.*ݑ�9టoL�Z��-s�)����L�3M]���x��^�t�M�Dr���+�ň~�ȑ�;s�t���ۨ%V�Ad�l0U�"E���\J�G=�E���J���tE�b.����W��Ԗ7��mm�u���a�;(�P��IG��4&/Y�G�#�!`�Y�qލK�nz&�aNɀ�ӗ!\˽_=����=l�=yt<�E# ����[�Z���շY���� ?���<{�2�aV�
��T��x,Y��
j�4���j�{h��v���&�p��d�y��R��q� =x�R}f�)s�\�9��t���e�2 ���5�����7��k�c<���G_W0�� ���Ы��Y�i����iv����L�]�$���`����`Ln)��gO~I.�!�W܅�>>Ϳ�����g��1����K;�T�,��M*ˉ
"3�L�r��P"ЩC`3f�CC��>�]��l�W�$���2�ɪ9M �]5r3��]>f�gX��v�_Cv�mUHj-�X�Q��A�!Ľk�q��ث��b��+�oO^�_s
�	u��t�;�?��SvtwZ��	��;�<>Aa C��@.}��1����ckW����ƠZ��Y�xlP���ߺtNW���|�D�2����&�q�Q�}��^���CJ�DS?]���w]粈Ưm�"��&og�(G�˗��E��f|�|�-�g��c+����3#ʳ�gb�1}I�i��j�Cof�JƠ�{T'�]�T�Ċ���Z��;\��A�瑲1��iW<c��9n�
��P�&]v��a9goF�w�!��B�}�u� �loj�FA�������ԫ�OM�;�{�j��<��S,
�YE֫��Y�d����e����a��-t.�wjg'������<�BGEРa�SJ���0>�x�D2�l��N�x%	�2!$EF�DC�\8�[uOR�3�	�`g�}},^iL���Mzi���j"��zw��!�Fo�^i�F���%z.E3{�S#ܸI�S�d Ũ�zi�nRڦ�KhU�n�Ѵ��-�B��P��7	`F��'|l��e�HPE-����ބ˞���N��{Y�7�]�7��:����vV�pμr�S�|���Ȧ��ޗi���)F0��;�WD�Z�gp�����\���W7b�Xni�7���v=R=���O��2}��O3Hΐ�1z��C����7?sfi� ���7��"��#<������y�p{a��sԹ���-Zd�2�[y����#���'΂0��τ���K �X��F�rFÌ��K��֐�dl�޽)�W�U��n���\/���H��-@��WF��*��2d�\�ϣքQ�X�?^*�M����淎UU��%4�2?E���I�]'���^�*`v�s�dkbz9��g��Y�sU�-���5�v��MO��fkr�1�`43���)ƣ2=���m�N,��P�q�=骹h?�8q1-�B����a�u�ڣ�@���2�6��]*�L2�l�Wk[t����s���F,��Z�Q5��6q�Ő��;�	{z���o���X��o%m�6M8/��&;��u]u��(%ًmw�����xx��p"��U�?y�������ur���N�0o:+���t�D�o�b�p�c����́����&�f����ӽj���+r[��/D��З�D�����j? ���0~?ve~>a&$đ����S�mhIO�mH���}������1m����ǃ�sK�Ȋ\.T-,������!�M�(`���]`?���2�k�ś_�ޖf���O�u]��W0ΐD��[Tv�m�U΀U�._r�EV���<>u��X��PEzX6�)נr�ws����!߮�:�q]`��B=AF|B^do�D%~ڊgQM,�!S���:��p��x�9'\�ڴ�(e��R~�����2-7��f�]�O����Z/*��6U���8}�TD��:V�ϛ,GN.kέ�O{�^�������+��za��x`jˉNY�F��̯��G<lVy&vb��zdߔ-O�Vu�Ǡ�2�)���k/͋4�;�N:m��`e^vLV�l���@A����콶es�x����s�O�Y����b,C�� �xxì9�Z��0����&��ɭ�s�;k^�)����ު�`���ﻯ^ej�P�k��"Q�.�1Ӵ'��xo���]+�������H 1٬�\�F�x��Ż0h\jdt�O�P���ْ)�ޒ��|���uz�sv�[��R��eu!��;�f�P��[�WLԤ��E�p�r�v(����޾u2-�eA�t�o��?���]:_N�:��B9���C�P�2u��i�t��TG#+,��_<�+s�q��=;X*e��w�E1��K�d��T����J�A�/������ɹ��;[�V��ʴ>0_u�ҙ���e��u(���h.NC#�w�)ҋ\:*�����b��Q�ʲ{`����Mu'1��]E����wSR���m�Jw[C�ί�N�S]1t�(Q���2��Ff��i8$�7Q:�a�uwU�s#[Df�#-���O
�Ȍ۫۩�/�H�.v���N��nU�燯��l��/J��AWՙ���L�������p���E�t:�&WN��,�X0�6Z��6%I��f���V�"��œ�J��:*�w%���)z��G@�Z��Zȡ�E�S��34�9���j5vy�kN�_���SY70�#1*F��Cm9�Q��M�^Ε�'u1uX�_%����A8;ҏ·
����"��ŲH�V7��&�C�v���З�Z%�S��S�A�7�����zto&��<����|w�%�c�f�Vy"�+�!���Ҿ	O����ڸ�HͱX�L'7��+u��T�6���s�\����D�|���o{z����QW��ڮ����]#���z����Y�xA�a��h�5nT}�Eg��oq�6�޵Ǩf�R���Md֭WSswi�;,�J�=�}a#ʑT�.�C.�M�2_W:��G����ɱ��UgY7&eN̶�M*�Ow�E]��UʓV��'}�e�[��v�7�H��7*������r<._j�ɋ�[7kn�Y��K�+jHg�bBvv:
PL�Gn��9��^9wx�<�t��qL}�r�1"C�qr��䡶�ܗü]ʺ�u�$�z�V�f�s��7�G�G3O1ñ�b=:�ʢ8�[E�C������b����v����Y�����o�)�����RsKr�[Y-3�(�ڹ
/u�{���4�S��&f���8$�9I;��o�kǥs�մ����$*��⥄o(mv��Ŕ��S'XF<���sM�t���. �Ϯ�-���������&�XF�ǯ����y��E2a��9��x�
<�����Wv��G4�,�c���fi�B��Kfw�!b���4j��w��/.v6�����Їl�IAc}��ւ�=NnV��iJ<�UE	��<}9��?o������9��n�vJhy���p��M4Z3D6�D�U�>�\�kMEE}3Ǐ�}��������}?G����o�ܸE%Q[�X���
m�,Q6ڳR{$�EULV�1��珏�������}��O���9���]��TF�E;��j��Ü*�(����W��*(�"b��$-�(�=j�)娊6�`��UG#�����55y�__IETW �l5O0b"6(�E͆nX��EA�؈���������3�r� ���nY�gURLQUmmQG,D�UDMr4QU�*`媝h�`�55U��ZuG-[�4�x�^lS5MQT���d��q��αUD��TE]�A�km��DDUQ�ų���sbv�Q���U� ����5��{�������WW�E�N�2��UӮ��F���O�}dV���q�5�o;�N8U�ru���Qٲ��U�U|'��a���a� s{��\W��m7���g�B_�2OX嬘�{f��+�S���ĺy����%͞�_"�\�jE��K���^iמ 'g-����|hO�ё"��iO0��y�J�����n�z��n���d�[&�� 1�D�f�]�û�~�T{"ѡU�S��m��s5���V�M�r|t�7�
��kTks3f���<���>��LƧ��DB��)�j����s���ل�gw�o8`�����,0�2I`�S���dcw����m�}����\<h��s^��Wi�NMk�P�]ŗ�F4��qCz��PY��ҳ�B��.�����c�n��	���3!���d,	��z���a����aԅ��u�弅�I����w��~���D-�G�\���*g/��I�|��[���qm��sӫ�n��H�9�L��?5�a��+�&<�� T��� p(�}y�ف�9�z�%�\f81e�ݚ�4��e*��T�raf�s#��r����ͻ��n���öx��驞��.9�j)���K�O�f-+�_T�d��1:���S�E�)���ڔ�)���+�s+�n�e�Oo�1
��c�Ko.��6��Ģ3��Ol��d�7W雓x�/q`j]F5JG��۽T��;����"�]�g,]�_b����� ��<@����!�B� ��J���5-�,E�����֝�>	�\K�v('�q5?*_<4�Ä��Oɐ��m�,��7a�۝�ס�1�@�
}�4���,^�Ȗ[~J����e���Omw���@6�{U�R�I ��/[s�(�&�2)�����@]s���+���J�y۞���Eec
E��u�n-�18���k��z0��1T�v�~�D�c'vj.�%�a@R��Um�Pa�0h�UsZ���IX�LS\:��{�ύ4c���e8M��!�T�q^�3���m/I�a��D����y�5���)��Jǖ�P��5~x�t��9�PZg����n�j��t5��{O����$��1�@(�e��27�Q���_��+}!�-pp	�D�wM��[:��Ln��vݓ���KO�L����RQ��� �S���#+�3f����l�V�N`�fN����ڣ�	p']446��Κj̴y��Z��4�q�iZ�?���ci6�����w��|3o�J��~&F�:��Qq>�Ά*�kC���e�zz����^U@���V��4���=?�Wr���lr�[��Bj�΅���^��j_\��A�Ry���G���s��K�F,�ѐg<��J��{3;�#���)+����;2��_����k��˾ӍVd9��|Y��Ts��}�]q�3����t
C �2CF xG���G3�3"~1�ί�}���v-��(�d)$Pq5�AqF�d���S�ҦCM�"��1i�>�Q�vc�Z��/���
7^���db����١3�%~�'{G�9���@�g�L�G��(�����'�~����B�FK�a�d���81�N�M����5�33�(7)	��
E��O����_<5�T&�ܹV#UA��m�K��U�n�>�A<���i�Y��5K0L��<�O�͈��:���a��*��􈕽w���I�SP��"ص��W�;w�^�\�m�^��Mk�Ȇ��b���ȵA?6�uN��=������Ȗs^��O)X��1n7ɰ��l+$L5�}�{�F6k]E��4o[��x�H��Vn� UD�>������zt/�V=�t�\
Y�n��Z��\d�e%�]WH�b�韺�B���gc��[L"}o��J�a���t�Ǻ�����U8���˻��5��i��&�eu��ɦ�9\�zc�!��|ӅO��2s�#�����1�EnuM(3$��k��c�b)>7����`Ϭ��v��b���A���, 7٧�[u��nD6�2+m��Bf����9��;��Pw���q��Mf��K�v���J��h�ܱ���2�m̙���Z.��]�xQT�9��D��� {h}j<�A��g�����z�n���T-�� <?�����Aa��-*-(x֣��R��L[��ɦ�K��7�W9,�Ka�񬄎دC��]�C�d󴫹ڲ�>ը��s�*^/^�1�L���3�N!��3���2n(�ds�gփ�e���0c���R��Qw�T4��LO��������7��<�j�z���͑� e_>'�`�.֘�-��O��Я����L�<��]�qd~ՀZ�s�f?�.,����u�x_&{��l��t�S�d�;�`���́���y�)���ǒKvd����Ǖ���2�1=!-2��0��4s��C��f�^LG����~���{��Oɹ��p�q�a�[/=_��D�;�����ts����*`�9�gO��mZ���Тԇ����9���B���	&'��C�C�D]�'�/L���X��݋��w�*`k�gO��=�3iܟ10��wFB/6���lŚv��X��0� hq�-x������ڵN�3n�|7}Q�~����-,�c"�R����{��Cí1��E�d�Π�����������C�WUH�(q�Ӈ.��2�Kw��r�z&H�Zހ�Gv�1�q��>㣳��C��Gv����X�lݔ���=�ڋ%�q:��}��ܾ�	���7�9]L�c�B&�k�d���9���������#�y�U��C�a�4�a�+B����������6���;܂�_:�.����P���`��z��+섓?|�P��n��ά�4��^��p��'�Ǟ��'��-��Eۊ��N��=˴4Sz�[;qq���j�x��<�Yu^Di��R���)��lt��)�<G�m�#�V/�ٙB��qb�X�$�lU����rT������[ !��HA��h�Re�l�'�q�eϽ�� 9cl�Ȉ~����u�����E�}�������Y��Dy�c��Y2F�LH���_|6*Sm��mG�7P���u�^wD����1�0b��;��[a�m�рg���04^G�6����/�M5Q�@�#�q7�6�m����� [k�wal��1���k�������-��Pp�fL�g�����wcL>J�p��t�����1),�F���"����屢�>��6�=��̛֘U���O5���C0�c����&F�����L�h��t۴z��L2�y���鑯,�b�#�N���Z�q�g�����/�39r�v$�%��w2�s[�d��{�9�#���U`H=�s6@��WpYMo�哖j=z�4�5����O�P:l��Gޫ|gbO�۬I���q�/�zّK�w;5[���<�7d����&L']�p�a3"��}߾�����{����?��dRDp���+��������}���߿	�o�L�XEOG��d$���Q�u��c�3O*�h	���)�ū5ݕ��gr��Oj#�b�D(��������v���4���C3s�����v{��J2�7f�:ṏ͠��h�O�g~�W�]�Sg��`�[�o�e\aذ5���vc�cY�Xl���K��6C�ЃiBf��p��DE���^Y� ՗@���/}�}�pZ�l�a�\N\����NA���y{/D��&Bm�L{(>:�x�/5��a0�B��h�{缰��2����4 �((�W�k^���>��.m�>/%:��K2כ0ܧ��vmO�E��s+��G&���;�cO��=ҀZ=kd��F��e�䪙s�yc�eslZ�I;%�v��]�[;*��uߪ�xD��r�z���FF�\���U)���۶�ru�03;��tJ,޴�eDͥ��!f@~��M�>��?�P�>7��L�p��� �{�~Nbn�����g ��(�O�h�6ג�?2��z�"��~��L������3��[�]_/����vY�T��>a=���K��9cG5�[��Cap+D�*��Z��,U�t/����9�{��\b|�g�쫿*y��c r���ޮ�V�s1�Ȼ1_l,^���R�S�:\���ʨ��HY#�x��r9��3߮���?��o���tP���@������Ø�[�����~����d�$�Q8���\A�v`������ٖ��Ŕ"�U��Ds-d�v?�Q��[]�ѐ:|ָ5/ê��)�s��*�3g���CV�T�)fY�
;���%���/M�hL���͛ <fF<1e�U��")��A��]	y.������D��P�*�u�U��5O�δ�j�b>�ag|��ʟ��`šy�E��H$o�|�w��g?X���1��#%�ޟSMvȸ�
sl��u-ۜ��\�/"�Y�ڸ;c�wf�m�a"�BB�0�61�-j�����y�8�\��hO�s��_;6F/�ǧ1a���b��L�g�o��$i}��X�y-��0�8K�S]�ٍ�T����00���G��8n�r輻�H����X�	���,)t�C{��f3�o��-x�ҟ��v��M
Fm�
����g����\�����O;���ؾe5W���C%Si��1@��*�Rqz}M��ꄫ��2x�e3��AvT0�1o��.��(����Vu�yV�K�|f�k�r)�j|P ja+��2`)dKse�-�S6�mv�VX[�mB��j}ݞ��P��Ӱ��1x���sUh�/��-VؚR�d%1z歪�	3���i�������	u��$�����yǆ	�2�r\�����Q�gwv�S�n��u̸~���|�w�Uz&�X��������<@�!�CH��0+y����������璅��3n����C55P7��.*���-��9�c�ބ˝�{d���zm���G�lU�%�r�M�E��`K%��^͇�T"=����!)o�7�|��wKwTq���e�/�C)v�AD�t{c���>[B�*�kr��|c�,��0�0`���?[wdC��M�&�3"�3@���;0(�x�R}ҤcpVn��ߍ�;��F0k�*0�#���ñp����Ծ������'��y@�oT�~�x�[Z�7C?FIP��D�˛�-��$q/X����@K�q��'�}���4s�u�	�X�d�8�	�L�w6�WU�k0��;��б���M4�s}��rA��="A2o=��t^X�U�v(�]Ο����$��|o���zP�<�/���7����#!���@i���ˊF(c�y4��!�4ܠ�e+]�3���Z�$
�g�>T�֒b���v�ݛ!(��A��O�:��maV���r��ڴ�tMd"��_H�s/��Pf��sB@~z���vo�P�0v�]c
��N��`Rn�+1�hJV$gb�^������<>JU�5�T�x���+��E�k:ŵ6�mcU�S�&��T�(UnJ�O��t��){!���6�23p��g3����f6���:��6�Io+�)u��3�ag<��������JeHd� ���� �`��J�v����l�\3[)�>�1���ˑ�7́����;�����>�yx�P;*hi��-m�yC����$���;?r�|�(e��(}�ͯ@qlǕ�b����
�y7Wfޓ�җ}@(�Y�1P������!'�/��涺q�0˴
�,a�#6̲�7o��V�u�֥�q����Ŋ�1��#�T����8O4���o�k=��+B!���E8����tG��w�B�}��Z|(��q5SE���6�X疩�tt=,�;Lov��u��5y<kSVdk.u�)���3�|�q�p��v�wdu���6��k�n����7g�^%S��	:f�9=�wj�2$wJ�ۀk�,�Ю��,ΡA+����yaO-��!t����B�B.y�<�p ��y�1Aנ�3���S.~!@��5C+��+��~�Y=*�?�E����*/����'������V���:$�(o��_w��A|1R���z�i�b�o2Si���1���֪	~��v��CK��#,������q���3 �}1�
��ٲi�����V��5�3�?OKS�d���V�&���]\��:/���wx�wN�ф��j�wW�ڬ]͝�I��ϸtzj��6����f-5��Uj��7�z3{�sHu�O��w��5{�=}���`}0������Lu-��=�X|��2,{��/�G��Ra������� m��u�~��Ѝ��XX�Uԝ��窙BP�5�9O��Ɏ`q�1���Px��0����z�����%����g��/]�%��;*���/P[�d�Xg� ���5#[���6��k��b�a�;�g�d`�\�\�L���R��
��֪曚}
1����қ,�-ގ����3�܉�ۦQ)�J���i����n��t��D��۰p�*֮��A����٦���j�i�Q5+�����
P�8^/�7��tb�3���߁�-�İ^So{ê��y;����Y�GfV�Qŭ�Dxpފ`�6Ξ�a�ٝ����D:JzW��b��S�&�_�ٵ��s��!����-P�gA�D
�7�i�ꈋ9�������lW���4ܝn�RAj^1Lz��N��/$�Ll��X��^Bڇ��zw��ȇ�����q�&̞���y��l���xc�������'�Ѹ����[�N��*4���O.��x���[kD���kf`:){�p�tzn��͛���ɰIX/e=*Ѣ�m#c ��'[��l�vK�U�^�=j��t�f�R����r�����\���/(�P�ɒR�5���b"ld�ם�o4š��:��3�T��\��2@�u�;�ȡ����T�.B���o"z7p��$=����r�a1˶"�-n�G;��,]U��I����\�]�|1����͝A�r.H���ە�k�&��P�J���af+4��U��,���he���-�ΰ-űe���8~����8�v�C�D����Ǚ|�7�gmL��ßcb��luM��GG�h��jbͮN�����k�î�`�S�8��T����eGnb1�ٶ&�ۂ�ҹﷺ���Γc�����m��)�ڬ-)5&S%�ܨ��We��PvU�Ʈ�I�m>>(M|�x�l��:eA�I�yŒ�N�/��[ғ_vc��N�Ϫ��XȦ!]���7�^
Wģo(c�/.�v�ϟ��ܥ#CE7^J��z7�-	�����[��h���T��b�XZm���"!�{$\sZD,�a^�!�]Q��.���V�.h@�NH���A�\"ѹn��ˢ�B�Q'�fLOS���]1�m��v{�L�o��P���Yޞޣ�̏o%�&6���NT(nIP�p�萱��t�D��E�C����f˲9�i:�m��iDK�)���oE��71�`��*B��!�vIyճp���)i�wUŒ�L)҆1����Å�T�Z[��'ˮ����9���:�7�1VƉOb���֩�|Ǝ���}Ѡ�oq���@˵+J�ݭ���3&��Z�K]�й��V�6"�춍�{b2)+��0WP�f��.�v��<��|5���J:�ȇ\d�Ŗ�J���h �+�Es8t��l3YiX;���8�j�2&�s�#�쫱�S��J�S�iI5u�5:��l�k��A��h�3���ʻ<�c,Z�<���wM=:�Yx5���U��z�Ċ�u��䂲��_+t��-R���B�����H�):.-ݐZ��-7����S�[x5�W�e^+Qq�{&;�ь�3����]xT��73���R�U��+�ɴ����oB(p��#f��%ۡ���t�@m_QB��]��Ʈ(o�j�-i�_Ua���t���K�6(a�j]m� %�8'�q�̕��Fy�4S].C�5k犩��dH��L�9�2;v%T�Ex��G��;�qۼo#.�뺈�x�����vլ�1�h����,Jj��8�fSʕ�%��.gC��;��e{o+� �W�z��U��^��QOQ'��J�j��U�4�7��ME+���Ft5�2��sA�*\��:\�9Y4��9WroW�t*l7�K=5����6���S�A�i>$�x�>!��cwi����<��G�E0TDηͨ��u^?�<x��x���~>�o���?��s��?�&)���Z�-cZ"i��9������h�(�
�7��9�������~>�o���?��s��cT��Üə�0"(�I�&j���AƱQ^����������~>�o���?��s������4�QZ�D�E�_w9��9<i��DSL_m�j�*����b ���J�Y�	�����b 
���ELQRO6��"��m'�i*(�����"���6"&�=6� �b��*if��1LQM4�Q�j &
�Q���t_mDTU�TQ�����Fb����������M5$QD�SUUCD�E'�]E���LA|B��Ӫ��m������cK͊)}X����U@U4R�LQT1PL%4�B#�+JL�
!�����D*"�)(^�≣$���Z�Ry�! da�}/y7�2Eҵ�[`4��+y���n�BzI�̮���bŧ�v�OLU3n�_WK5�Ju���x�r��h;2H�.�&"[.�B��P@��$�%(ZE2cA�[)6`A�dĚ@$�/͖����"�0�
�&2�QDʁ��<a��D��������B#��T�"N�x��>,&R}z����.U�snB�慎�X�$S>E��v��-�[nL�R� K_�K9D�ف�״���@���<�l�oL�[�*�\��)�[�ܳ��]l���]!�*T��z���k��_ o�d��?r��$����U
�����&e�8�6�0�9jmW?�����U�C������U`�C,�
�K��Bm�p?���A��x�Uj�.���o�����3�=2}ck�������FO�����7��S���s��n�5Y}iUVA�*|���y��U��!>U���[b��n�����I氟��'��6�7�#��u��R�R�z"%��O57��k�&��5��};��0��Pf`�|m^*��n~Y��d�,$A��B^L��^[ZDgM5{&����:�>z"��7OKoIm�2�/:�q�_��1flTi�iC`=�������Z���qwʷ���ڬ5�x8� �u����v�!�C��!��+Ѽj���Z�;cû6C,&�Raz��|1H�l�e���r��YX۴���b��K�l��Nb����v��z� ��j�D�EEx-��ix�j���.�~�����{�4:�@���y[���\���G$lע�6Q���s��>�M)�}0�S��_;��
u�gn��*��z�\�׶t�iv��W���W�r�-V���d��=^}=�����ի��da�����0�w´�����$Ǿ��6�$M�	*m8cP��]��������%��t�
�d�}�S�z&)�_�	�hp�}#�z�o b�[O����ԯC>vmU���b�S7eP9�P�p�
g�Z�5��E0]^3���b�^�M�nr|���,�`��d4F�2aRY��љ����Ws�Zkѻ�L/u��(V���6�ɬ#p��C
��r��fcZ'hU�w�s&�`_�y�+�>,W�W'�+���m^��t�k�q�[�q@��9)�{d��Uò��h���r�m�����ֻX*��K3�����Da"Z�.�P���0���LM��/)e[j�+�� ��q��G���v�i/�y����O��b]�4��	�_TO�����Z� r1~1�78��f�mx�r��Str6f�2Ul.b챂4��,�&�xb�+�]�޾R'z�s��w�[:5��Gl,�ٚ"�v���$;��4��#����<1n:2D�ȵZ@���}r�[�`�+6���ɫ�xv�ȫݳ���¬�K�a�kw�L�{U�yS+���"�yw��>�ʭ5d����6O����6��~��ϭqe��l����ƪ)X>�6�)���VRV}놈ѭ�:k��f=�+��f�D�1Ã��w���}�0�R�J�����w��c>φ��L��~|�c.�ȧ����� 4�����o3��+��0�벓׈��[>�Jy��a��:��b1�`4 �S�{�.Q�^zw�f6�[�
���|:g��e�0y�ol�eg�>T�� ��r�66��`m.�5�1曲Y/v:J�U�3�np�=1DW>�CZ݆���WD���+�f����\�r'D��߿sE|_1��<.N�_=�W�	��R	w��O�W�Xv�?��?I��n��lf���ߐ�`�KW���t�)z��>cWck���s�Z݁��Бn;=�^Q~�!C[�/�&,���G3X3��O9k��g��{_��*~�}�����������?A׿*��qmW7#j��[ X��|N�T�(�e�	bo2ֆ�R�K]q�fo�jZB_TM~>�?���7u��x��;�t��<���~~ʹu�O��3�y!6�pKϺ��4>ۉ�ѣ��U��5��/VC�l�۳3uM��L[QЮQ�I�FTN����M�Ȥ�xW��Z��qj""�I��i���u�l��V��s�$C��/0���F�6/2����U�3�f1�N�/To��u�d��N4�L���T9��Ur�^��Lw+.�mw�C]��^�Q��+�j=��y��6�j.�{���;v=�.D)f������
����vw;�����#�� ��<0�7����xo:ؔ�=��k��L��3����:�!ݝ�̓L�~�j�"lbX3^���Р�ɇ�9�w��S+��X&'nֳU,w	��`@¤j�G}{��CH܀��5ϬGU ⢀n��ٍ�c�b�i�	y�ޖg���1�	����y��5�Ֆ�yn���鯌��)��T�����;<G�t�;9��N��3~O�B� qej�W�1;�|z�"�~�E)��CLI��5Qn�8�W�*�rs�y,5l,�%�g�v�mͲ��c3�^������yw��e�e���s��aG֑T+Fk�i��Y���?>����'��sM~D�A���|x�y�]���V��<�2���ze���Cu����m�k�`�h�"۴��a���6���cm����'�K�\��˟0/�����?|�D�/,}��/_O�,~|U�?0����bf�o�_����>F�����h�k��	^~U�a��H���i�؁l}��#�|:�7��?+�G�.�Bٜi�Ơ�r��i�ώ]���
,�"r
z�3�8����.��e����7�,��������I�l�+�;�V�ȱ o2Q���u?L�|�$��7e���z���Νv�fb��Q��'��k��u����A|_[[;���n�׊W�7�V�T6v��N��v��ۦ���Zi0�Ӝ���>a���{=���5��\����z��~�ɀ�KŢ����~Q"@�Am�a�6yY}f/M�r,JSlI�gO\cz�I��R��F���)��U{�t��5�i���p��R�k��YC�&��!߄�- ����IL��Qƍ�.m�4n}�G��D��Y�F��G#.��58�4ƴϠm�)��2iI�_U�3�����E�^��Ю�'���b����f�YMŰFx�woE�g�ˏsX1~Um{�X�nD���J����,Y����tG4[AՒ�\���.����
7���q��B���5>"�����ǻ�eT\qU�×�Z�O(���ut�-i,^�a`��:�����u-z�-l��Ra�ɨ�C&��k�څ�x=�AeJm��`{��r1��8�O�[��qR�m'����!6�@Mq��鵳!s�U��M6����q^�3���T�Ƃ����c�)p͇�WSG�LB}fD�J'u;1���۫�q��D���.$Y%����B�u�y��^UI0�����m�I�s�F��.�E�������v�w��)�Z��������*C��#�5뭞j�B��si�r�}�Z#/{�����������^�e�z��9YD�.Lm��5�Ǖ�³�s�����w?nu����ݺއ��b�9����j"˚�3W��.o�v�=��E�H��r�s��>�+�s-p�|G]@3�vr}������G}C;z3�&d�;�����C42�{��~��������Y��/*���QN_C�g8r�G�7[�^�y.�ʚq�o�Țj��L�k�<�lc"3��I�?h�~��X�з}��㡒O��)����o����~� V�OX����ó�3�C(,�$(�����&��/:2�(�<r�� ����
zG���%~T>L�<S!�^e���9���CP��Yl�~��ob�|\.�y�Iْ���{{$m��H-�;��T�qA�����ƚ�r[4�vYZ�^�|rf0ȗ�Bj-��Nd�5ۻnr��A���Y���Z��@��U��L\����7�ġ�1��^��+�b~QkU�k���M_�D��gѶ�,^�R�ĵ���w&�ѷ��<e�Z�CO����Gz�'���{�׭�7#�At�>�覱9�$�-r�W�����ۤX�{C�j���m
�]$�s�����>B�@Mk`t��*��oy�o�$�:J:\�z$I�	k�%9�v��;^;����������T
�-es�Zgc�+s4n�$�����6- ��@���ZnMl�ۼ��t�鹻7���/w��'�$	�G�f�yu��%�X=�����]�Ld+�����6����*�`J�NY[O_z�u�z0^�z�w����x��G��#��c���J4R�������*xM+Z���l�/(,�a�^�s@���g�B�ү�?����Dj�0zv/���ԆhħZ� r1f"��犡��ԍ�nE������ꃽ�Ξ�  �� x�� ��5K���z���i�Y�K?����<�Cr�wW�+O:�������Aa�.rA�x<�ɸ�H�2�U?�J��\�����
��Dy}���b��lJ��nI}���~TDK]ls��{��F0r�o>/%�{��.���R�֛(ξ�8�~��2��d.a'����=��M��Td5�����b1�`0.��7��ofd� ��Ziu�	H�Pޙ.2��j��2(I�b^Y��v�wf����m�>4t�����s]�if��� ��=�U�����CZ_NP��6�~l�f��.)�Ŀ:,!�_�fg5��Y�/3�jp�"2z��.����>����^A084���-�.��u@g�Vk�	��,��<��^Li~Y����_J"y�g�X�U4s�r����px�2�"���9ci%=�V�p5¹���.��ޮ�zw��#6�8%8���Ȝ3/z��}�\�~�ҷ%�6bZ��B���ٺOwL�g�S����/��}�H�C"�.�]�JZ&������%�)3����t+�p]!�|�:,չ/:�P����7�(�FN$��T�V���t|;���9����ʹb݂ ���3-
5N7=��Dj��q�[b!�8��z�b��u尃mx"Z�ڧb�ͻך������^:�n��"�U�s��[��˵��{������	e��t�;�m����P��m%�*=����_�80:�ͫ
�_~I����9s.z��R-��uk�jj܄�<x���~#7hjQv���r����޸gU�1|���e�GMk��/�}��O�r�J1�k�Ha�2��>D��lֽ��w#��K%��T�&�:5���!F,�C=��}��f"B��5���X�M>��{��\��9��&z�&Bjiz�v�Bb��_���������_WW� `�a0]{�{/����v�b971ٖ�u�	���p�6}����і���V��"���ꐛ�ּ�*�S�&+VwK�\�'IĎ7	z��JYcc�Y��kQZ�ha,���F߇���v��*d埯���6���*<������8������sӮ�-,����:�ó��
f��}u�3�ߌ��ܠ���H�\�+�5^��0�{p^�u�c����]�tT�n��rA�N����\�e_S�~�a�.ę��Ԇ3�~�<�86v�B�%�eJ��qt5&��%g\c�bӛ5�ԏ�.�m�C��b��.���� sG�}������Ͼ}�����!�(?<>����D��O�gwRO�R�1�ɞi9�!&�m�~a���M������j���޼%P����4U�R	���頻.mk������Z�l�a<
f&יAa>����꺖M F&�A�Ia\cZ�q�l�ӛVgE�5�I�a�⮭T�v��!���C��) g���Y³���oղ5g�~δ�D:�Qy�.���?����bɞ�,ơ������q��#:�L.�u8�'k�Sߥ���f��9;{AM�.���I�i���v�-��"Y�f�6xų��wװ6"Z&��<�R���k�(ju܆r�upXj�܇�onAcAA�����4�Ѻv��h<Kb����9D�<���,���r��Z�卄��|!4�&Bm��+��y����G�މ�W��9x����噭����[�a-I�+��4yGyU��ܱs��)��@��fP��^�.&�%�LD`�.� NS�ȷf%ٮݚm��S�4R��5�����D�63��\�5�7ط��6�c��ym���O�P*2�ƊN���1"��e�����l�n2��E��j�m�R\�hE��9��/-Z��d|x`ʀ��N�:a�Wr�ev�?��<�vU�i繸�G�}��}�	r���i���}�`wb�Ƌ��h#Y|u3��S8�&Y\�VNw^Ȧ����M-���ݖ��S ;8������0.<�����W*rWc��Q:���Ǯ��i�|�m��ͶC�ŵHg������!6��:�iU-����ЋR�$d<��a]�,t)���I��ԡ[����R��
�Q�^�q/N;�3b�˵�ՒK�)�`�;���|����ryu�X��t��[�^L�Ǧ˥ƚu�-ή��d
g����;�m��dKO�ֿ���8Z���㱞�f�ײl�}�����x��ѽ(����f�m�^K����F�wa1��煙Fy]@1F<�j��SHW�C��8��pq ���'y����ԙ㟞�S�8������ĈDs�uoV���f�4G}��]����U�@���;�)q������$;�1a>��`T�^���)����M��n&�טJa�����^���fh���Ýݲ�8́8v�ꀲM�����:��K�?F3W�>����;c�3��$�$�7�0,9�t=�-��l��T�,A^���-��qF�CN8�f1l���O=�w���&�yA���Y�����;�Z�q��ش�"��;��5KnX�3d,�ќO�m�
 L
��]���Mq�6b�*c�Z�z���IZM�PLņ@k[��r�Is��;B�",��ذ)܆�2ƙz4��ul���!뮷]Y�P�|m
�ٷ>�M�&�8nq��Y��ն!Du���/��6�r��h�m"�-�k3b-���o��v��_^�{s�2��ы-��6Wb�����ڽ���2Z'!�vwvH�3�Q��кL�Jyj5�Mn���k&�θz���$��"]�9ΕWM�ѹnGzY�&�IV���`'��톱����\�ij�t���C����� _YC���	�����М�kl�A��༐A�N�kJ3*�66�!b��بT:�SBﺳx��簓��Nvl�����3�N9>���WE�׸)���Yܦ���P��a;�k�PP����r���Pu;����Ь�b�c6_9���^3��͗D삸s�)F�H���9P�Ƶ6�r�82�; )���er8������J����u9:��lof��>�k%�64;�R[���8�gGÚ�����]&�q��Ȇpž��|�ǳ�4���}q�CN����φQ��ʝw�7m��mN�la��b��4��f��ڻE�I5e՚���R��+�����Y[e��))�k+��k�B�/]^����"�ZlY�XɌr-�	�2��1B1]!y�lp�sŔR\n�D�a =�DR���$�Lv3����R�����K��˱�^j��>���*^:����5�J��.Q�/���T�[�[�9c'i�5.i�u�6�s]�5B�ϭTQ)�+u'Y/{e��!ڻ7xMq+�Ufw9�B�-8sN��q�&�5k#)��?fTP-=]}�i+X0�OH��6Q�W#|����/�ۅ�	����noN7{2czT�xV�-���]-�4X�ޥ�c[�uP�{	ҸI��C|]tr��c�f��U�����L}�w�V��YR�Q��]�[�2�>��ʝN�b8^u�����T I;T��t��8�ENrҷ��P��#��z���x2qx�B�9�-�zL�1��������VЫ�D�Ee���p<� ��ȽM��IOq�T^/��&v��m�aX��M�U�5��fj�{'gfwTin�%��mg]v�4�xs��_tI�k�V}��"��"Ay�}XÖ��N��woC��_a����(���{��ޤ5D���s�kb��N�S{X�C�	�E6��Uͭ�Rp��Ġ���ci3T C[Bh,�X�C�/��W5fm5E��>�/���*���Yo$��6 ��B_%LY����Nӡ;s�9��)�����ji
*�����10U��۶��bB���*��������~�?�O�������?�ߚ�ъH���X���h�j���4QIr�E4{}?����}��ϧ����}?�������D�SU3��~�B�����&"����oO������~>�o�����翂����g��T ��DQG#DDUk5RUDkTRQ�D4UDUU1RQE	3T�l�h��Z�A�
	*�7)(�����3��[#RAU���.4U�N�DPQ%�b4:����@L�D�*��)��l`�B(���"" 平PP�P�\ƒ���������(���!���|�6��yÎ�PP[h��.R�E͚O��j��j(*�h�b""�h�������z�|��G}�����H��]��TU��0�J�^ђehN��:��Wĕg��ƺb���ʱ��f]����ϧ��y�������bj�[���O�%?U(h���韵�1�w�
�3{��i���L��#&ֵ� ��`K��[K�'�{hr�Z�.E�&7����=������M��9>�UQe��e����M76��kЖP��],�@�������A,9�?����y
�}�b��'g#����7C���{[�_�k�rU���-����ηCG��R���.����k調�4[쿇����%�z����� <I�tڈZ�/M���r9[Ob6<�U���Y[|���5n��9S��d�W�����V��9�^��C�F�pr���nϸ& 3(��w�ɲ(]R���z'�'\����li�ɦ���E�*:as� �yj�ڥu����],��n7b��bG��{c��I$�Zx�#��7�]�E����Ֆ�KO��w�z8F����6y�9e�-l��Rw΍��}Њl��w!�4Q�'Уy�Oz(�O�廨�nҫ-E���'�b.&P���B�u�=���3�qޟס�_!��?�Y�NZǶ��!D�~���}\����p���J��<8k۸�IHjL�Z#��Y�Os��]T�y)Sl�љy_;(0�q�͏�
���̔���ʈ�����G�j�v����HAj����u&�ji����o���*���jv`���!��{�ÊU�D�H4L|^�Ȼ����N2��1���5ZĽ3�,���;�`R����+;��1���=��4Qp����������W�ͽߋ��3E�͉~~����;\��3>M�ĳ� ������l��YF�@X�|Z&�g���}Cm�0�q�a���&�.�RҖu^o<T�I�������(�W��Zé��#��|S��p^|�NN������{A�~�Q]�˙��e�3H�t��u���0~P��9l`k�~���*�(лc�}�����V�z*M�0�@&l疸Q������v�QN���ă0��=��H���qLݡ���6 S��V��zz�t���ox�2�6�%�+-uk
j[`K��v3ʖ���6�e�I�i��Wl�!�h�l����D�VG'�[�𚚽�	�=��'��-���V�͹vt�����]]U�ӷѭ�ڋi��dŚ�M�j��+���0$g�����H�1<oH�U��s��o��榙�����ud���1Aנ�3��mQT�/�'���yF���s]���%��2�*Y�8z���-]�.�r�u�pX��������Lp���\���X����'v��d�}����u�u��z�~U0H�hNv}}������=��#�t�J�QU�p�V�9u�$K۹�e�Y����HLŧ��?���>{
�E¢�~��k~grT�D`j(��0`&��UQ0�>�ػ����{��X뎹�>U����?j���a�����sP�Zᒍ���� �N��T�ҋ�-���
9�<�;�N�^mL���u����@S�U��LI��&D��%��mW0(�x��3�'[kW�v׀�1�F7_u7PFD�vC�v�[�yAl7�3��*����ЄhSz�T���G�q=���q�䤰���=Z��tQ1��3ڋ=���F�=0f��I��ᡓ�sz�)�'��XUF=z�x5I45�oTʈ.�ŧ�ʇ2�nK�l�Z<}���|�@���\��_,6>�xV�����u�:w�UT��%�zD�6Dך��0M|�|�M}����ʢ?,"z�۫�1�|��	����ח9�s��a�a�)�=ƨ�?\����3ϲ��#"&T温�)�:��0�s�uv׸���Pz�'��<��"��;2u?6Z���|{����{�Y}�Y_*�F�D��m�7�N�:��Z�?T��
j/�2\��M��[瑄k�y���n<#t�Yxt^z���{+�Z�M���-3h{ו1����L&�2�BlH�v���
Z�qGXR�Z|��[dx���it��ʪWV�m�3H���&�S�slo^b��9y��O'	.�OoD�ٕ:��Bs���XR��2Lר������?�y�����	+��m�����S�E��dhZ�^ D&�7!4�)�0�u��	6�C��q��b��h�'�I�՘I3[�҈fW�7�s�_�TUm�ؿ�e�kM�,C����-wU>���H�ֻc#G���~!�mX���4R����Z.����.�6b�T˞�j�n�srኋ�W��⃸�P-��,}���ӭҤ���ܤ�ř�搯$��19���
������ٶ�mku�b�!�h�m&�.���t��9J�w����(�<ɧ��!��es�s_�E'ƿ��c�Z��@���/��V�QH���m�]�X��2�]����=�kzgl��<���Ў*IrG2�s#u�%�ث/��55v"��.�/��6�����	�d�n��m��D��]%��O��G7b���
_e��馋�X�P�
�`3b����yu2&qz��t�/ާ�SMX�6f��vYَau�{�6g��i��G�\��cc[�(��*�㟔��]Y�;t2o)Vyf�ǿ���U�$5�I�����W��VՃP;��䅅-���w+.��wdyoeP�7�{Va)Wwu5ί쿮�S&��9����&n��&T�=�FF;��;rV��Q݊7[6�̒�l-_��݋p�X�:���|�0��{x�w"����y�/������k��S���;���"�8���dy�XL>#οF��ݯ�������S���b�����lj���q�@�Y�V.�߬]���1.���M�M��t������2�LVC��d��NP�n�[h�"ĕ6\W�ܺy��|_G�$��7�o_I����
�L�s<=�+�sn�K��p�� ĘfϜ�J#PO��O;ի��5�2�jdM;m���I&����~48s`~o�+�ʔb���zaT����2��b�R:9�b2�W3�̵���آm蜖D����|bW�`j�����QQ�����R�H�y���s���]����Ŭ�2l�ʦ�	m�P�[x�|��>6cMȐ̸�f�`ذ��r{��f�b�04F���7�2統I��H�|���=�S����zt�z��xU]�����ְ�жc�m��R�a9�z���kߊ��ߖм��
���W~�������B���&�Fk���>g��ϧΡ��\h���
�j��F,�'ͰUfû"�
+El]��Ƭ[sVё]l[n��&��x��]�����"����x��WUC��s6Y�gm���$����6����յ:�Zꂫf��]�����s{��Ep��a ��g�"ařO��:峉�'[nK��n�W��q߈y�7���ǚj$�3R�8��������r@� �i�e�W{kg���z�L�_�ͺD��s�s��Z�GlP��g�|a�1���� WǿVA9K��`�����7��֪�ik�x�p���ג��Mh�,�3��Se�w���c	�y�^K��Z(�n�~"ղ�Y�\�o#[�9���3�~�^�5K����ZXM��,�)!ߒ�>�>=��il(�/c�y��B��qu�hc_t��Z|L[�l.����ިԤM���G<D��� r��߿~�fP%�1��+�`+͗�6�.^ѝ�r�ɼ�g��Z��"sJi��2��|���d�uڟf���u�1���qLN�T��o[WK�Q�ȗ�,2jq��-���ƙ�x� ����}�a<7��}�M)����K�;����7�g8^]�c�\DK4���I3m�e��^捇�yg=T<�& ��z�ص��Z���_{�7�,�ZF]�E�k(r]	��_-F;��6�'��/q��i)P�S'�����sKEr�7�X��g�ޑ_c6��K3�>kje��[�W��86o��J3Uj�ѭ�a��N�	0�1)[�S\���é)ݕ�S!����]^\=���բ���]f�Shi�/Je���9'�ٚ���|<��Ű��W;������)�Im�!�Ă$���1���AOL#z3r3]s��t�I]
�����O�-�� gK^[H�<�/s�6i���gV�g�L ��q�ΚZ��2/�tV?^-��1*�q��C�wȚ�����ۼ'`uݻ���zh;���'	�2�S��6 ���-%>�R!���x�d-z�n��wHu�fP���1�[㸖��8�[e�#[#CG��f��]�\���onx[���j|�?%�Oz7�:����]F��"���1m*��k�y�2��M�8�Mü�@33y��on��":*5א����O�n/�*Sm�h�Z��$B�hi�\�ì	xM���E�͝�e�i�E�<�="l�P�������y�X!j)�� ��01�+Ss����K;6t��PԄ�Xq""~��煣B�G�;.����a),$b:��b��D�ؼX���kgo��*�60?d�����[�,���������������q��
~|�tS�����n�KL�B�b�1�s�m3灬���G_�@���}�?��}����v��KBFV2�c"�.���/��&L��XJ����1��Od�?d}��]�=�{�f�fy�t��!+��9b�^��V�����Z���Ù2^݁Hs�挳إ�G�/L�N�ղ�+�Ū���v*�.�h М��A�����z2M��F3��&x����`���GS}������g�X(z��{�f�5B+�u������GH-����T'1��I�+��bw
XQX�%��FDL����$u�������q��K�1p���3#��X~��C��`��:+�dv~$���rę�;�ik-����?%�����zG&=�nei�<�a5�H����ϑ�vL�N	׶�O�+o�>�Ezӷ�l�}jip���j����DBi �	����Tj�G���?�^۫������þ���j���;�[11M~��\q�s�h
�V�/ֱ#b�]����6���� ;���ȗ�2��IfX�r�xy�ڞa�ݚ���y� ;Z�}/e��T�OۄNih�y+�����c��E6�YY�q`�͘�>酑a�q�`De�ZƯ%�>�"��LR��.����z��%R����U�_�������
W�V��Kn��e&�ƅ«	������	��� �����"�F�3m����#�I�ְ��fX7�&Ǿ���{�3� �q�*~xMO:��_�<�'�e6���oU>�.&T'Z;�]y��'bm:=���'0��QSPι&h�xuowk�<���E�k�Gu�oh�'���'���Mi'py��f���j��X'zs����7ȢU�]� ���1	��_ś^��_�ԫ���FDH�Kۚ������;]����}�{����s��oo���m%�g�~�?TO�������꿠���6�y��[��X���*�^�!qT���\�� ������k����}��=��s>��\�aJ�g�9=y���f�ԁ�g2(י��5�ĵ��`�ۂ c@}���%���^�G��L�Y��xV}¶l"AȒ�F��~\�"1�$������b�Ӽ�����y��C;Ǳ��a����ئn��\��/H�E�<��}�E�llj��qz��QU{ux[�]@�ls����K7Ǫ+��-8���S\h�R��%���'r��t��h�$X�iU��ޚ�7�T�U>��u��j���1�B\c��)�9h��-�d{���z��Ƴ������'�q+o�a�w�Z��V�o(|;��.$��0���]��P��S�荔g�UӕO��|b��Q~������L��
�`.�]�'�żD�ӽ���2����h
�+���2.�ȏ��C%`/̘:�Lc�V��-v'�R7�a@�R�p�:n�i���S��wW�?�:1~x5d�K�Xd�%X��y��>D"O����V=����`�)�y��G��ut.VL��h�(*��%k���z���2�*�F��6���k���*�Ϭ���{,�I~C��1����6`EpmضD�ɷxm`�� �mr܌Ի�i��w6l��S(�,�[�;�ͼ����V������<�a|�S��硑��GZ2�n��)�������x�JT�D�>��k��=������;�W�%Syl`ҥ1[k|�����gb��M.H<ST��Hק�!��@ߧ�_��m[�X��≠ο��,�b�zO�Ѷ4�g�̼����d��eDFw3�X��O��Y�x�G�;�5����{sU5+0�Lb̲/���tlt�I�r��~����0���s+�]�ƲD�Vm��v�iz�B+R�߲��j+��+�5��"������3kHXE?��u�m}����v��5-��]Z�S��P'Ts���t�l��^�5�5j�E{B8�-'��N�ʾ�h ��11Z����5Q�g� TW��<�4ȝ�)�^`�5��L���i�1l�ڧ!�a?��5�n^��-t�6�	 M2��0/�A<��]^��A�P�T�ȝ�4���da���Q�;�FbL��'ME�������ɖ�o�V^���'ҷݺn�;�H��Pg:��k+�L�x�X��U;Ӻ�M͠��%�7�I�Nn���ۨ���J.��nB��IX�+4��`�ҭ&w!�*2�7�X:���s�&��z��ꇞdБ���О{�f�w���3 9�:՞�fVKӄ����͇5H��2��*����Wu*o��H�3���f!t�ʴ��r���U*05�+�Y���\������*ۥ]�ͦsZu�m��{�l�]n������d�mL��#]\Yʓ��Z�j�4q޺<��v��x���
O:d�]؆EٰE�w�1�Z��݊���<޶nb�����o6jjdɢ�|NZ�+�2u\�x�=%^$
tS��j�L����3o	=;�eJڡ|�CS)+��z�iܭ�j��N/�n?0���wCκ6������w!�-R���K�L�Ө��vx��[�yw���ʉ�)�ЯB��o����.쫹�d��.�{��d��CD86�:��"L�m�(X��őևvh͍ڳ�֗Z� 5�����k=4f"��ͫ���oba��ó�4vR�NeN= �[�+�Ujr��c�f�Z�#�յ�������Fk7 �j��1��\fP�+B�ƒ�Ǟb��9<�ۏ+u�;h���;�n�+�d�a�^����9ر��Ca�z�@�:�Ę��87w!��8��"��v�ʾ�TV;�NoY��1��톭�Ĭ�ԗ���Ė�����.��:��l���'[��+w6K��G������Y�@�����&䌅�ٱu����NT�!��n�2u7x��R������Ӱ�e'0��3�A�n��2�����g��M�X,b\�7ơy}Lj�.�#+��7�2�����1�T���"ۤ�]g]_i��j��v�H���������8��$9^s��(�9�- �4���a��;����]�<�]S�<H�%�:)`j���Y,�;�>���cuǊ����3eh�8o{�]7h�uD=����:iԨuւ!@�dR�TǙo����Z�A�Ոqe]�}ĺ�*��Qsc�_c�z�������.��,<��:���-�`���k��A�j��Ҽ��"�gk�..�L��wk�j{٢s���A$3L�炖�ג#8�i< y����q>���00�]L�C�ܢc�M�Z�l��XY��ݖ��v��h�K;�ϪoC�egX�-�"�,M80К�E�+{#_�	p��D���1��[ǎ�-J�������EsS3P����� �]�K`��.�r.�����:x��g��qjs�T��$�|A��`bvQ���l�IG�5T��EGl�DP����������}>�O�����3��䭰EP�~��R�CE�yǄ�[`������RD�޾<|}?����������?���|{��h����g�M4�5L@�D�D��͂*")>>=g�����������z�?��ؒ���f�����*���n&�sf��T�4�;s��(���∊+g[8�H�h�c�r�.F��ә�-%�\�&�UU� 4L�3EPڊ
&NF����DLD�Q4P\��p�P�D�T�UM���"�c�E5�Q�11Q�RU%DL�TV��*��hj�����$�)��nZy���T�IE$W�h�)�:�)��"
6}G �����sm[�0�k�BCa�2"*y'���r(J-��%m�c�����ɩu�np�Z��N�]��u�ĕOE�y8%��q��ں���xE����w�ܕ�H��I�ؒ5�<S��,��M��A�0��e�LFP���Qa�j��b�N ���0�#�DYDS�6�
H`�

")�Ԑ���2�5^$���Ϳ�Sе$���8Tl�i���v���j�D��0u0�0���|���f�����d��_P�҄��I��4P�\�b�t��	�-A�[:z�<��g֧�I�BP�K"��X��}�_}�߃j9��d����!�k�Lֻ�vL�t��u���j��<��ّ1�S�q�X���'`gz�&^�D8�J����aP�Ϭs�	?<Ȗ���Q�w����9a�g"h��Fv�z?!*#���{��O��v��!�9��w�|&�.oV0�G�^]Ɩ���W.������mZ�!�� ����薨�%?n@!�Kn?1��I��1m�gHlt"�"�WlS�U.1��&��Ph���6��Ā��U)�M�"z�U��U��ͦ��3*��+�v�{���U�9�B���H� ��a�}4��&�����`3v���Ic�R��4��mX��3���<�������ȦZ�R=����jo"9�K۽��e���s�j������۝�FY$W�F�Ja��kq{񊕯k�9� +}K�t(xq���ȇnT����k����0vZ�cw�o�ٿ"��L�H�6/����w.ܽ݋$��8�.J�L�X����k%�e�H�no_R�e�Jb�tQ���wi�A��fv�_Vr��=-��e��z������K��}��O�����x��������0�1���s��ϼ�z�����cߏF��'�֐_���ͼ��K��@� �������8�
�ب�E�B�i�.*�˧��q���5�oK�/����Z.vB�C�N}�d(_̐J��P5�)?+|}c7S8l�Z#B��0�fǥ4M�Gmi��w4�Jh��7
���}��`iI��`�L���Y�##wM�aݬ霚ԑW>'�����ɵpq�̴Y�
�Ƒr�f��\��h[�x��m��{lq����v�ݖ�~�ʛV�������E��~�/���g����J]��]���Kkh���4c�q�wPb��˙����O��M��a�M�1H�:�f�m;9f����x��j��da�x����f;���'D(�w����g��N��17��Ǿ̦��^��e��|��
�����E_G��`�h%�e���B�螽b(��^c��&֪ɾ�]0�Rz�&�9;崸�V���P�jd�d^�l�M��<,��J�Y��wWp`݅E�.x�t]��j^vF%$�%�m�N�T��80��we={.�u��3Td��j�=�w8}�ׂ�[^+;hKv� �Ƞ� j��r��3iĪ3�:�Ͷgr&��r�ag%8���7h����@P�b'���C	�y�h�5.��y ��R0�����K��%{�[ѯ�gU���Ҟ������K�uc�v��_s_����s��j��IWb��ܡ�k���ʭ}�/2����7�֠K��A�JޮE�W*e�r�vc���7v�����<������Z���B\lT_��퇽v�p�긹l�k�b�x�&��]�޶(Rr0�l���e�q؇K&w]R�}^�r�x�4˽���'��{�p�mRM�-q��6��|��
Oʅž̙{�䟯g�s;ÿ&hw峢���]���<E�e۹��N6H����37�BWKw U�ŕq���^��'������a���KP�
�o���p�S��C�����V�K�ʹM�/>v�ˤ"7QՀ�T���7V:P�毆��W�Dz����3#{�o�
rf���ٸ�W=f?`5C����§��][��^�<��ɼz��w�e3��5���k����N�y�;[8k��*�[�����q��#��+����׼��Lɝ!�5�,x�k/��<S{�z���rw���=߷�B���nXK�]cy[z�w�������Y@��e,�W�����FDM��w6uEs�����V�nv�42�g��1R۩�<�>`�j3T����M�'3���s،����G)�err�VL�n�D���lP�������㏘�Mג�+�U{��꼓�|U��e�3䭚�X����4]�G�U�����ݣ�°z��8�ct�i��ȃ�v	����鷨E�"_wbs��ؾ+E���܊���w-��UwV���V�uuet�y�������Ӟ�Q]�7�ل�r��&�Vic#H�7�s�����)��<�gS6��������H����7�O�y��n��ޅ�ҹ�3�{�f8��W"�	ߕG1!��2ǰwUeƎ^��V�vA�Q���+IZ����vT���x��Y���/v
%��-���W�� ��^��`W�e.�ʼ�D�WQ���N)%o}�p������>"��-F$�H��������/��'$D��q��#m��!#3��^H�B]��Ϥ��������dr�&�u��`2��/:��S�"����liv6pƌ:�����ov螀q�'}�sU�4��_6f��᱘�~'���*�_��k1�,�fv)nw�2�A�(�?�K,�W# bѦ�ټm��%%,nXnݬ���3���h���7Pm��=6��;D�
�5�z��*�R�X��j��ח��C3�C�sz��U�ڧϢ˿��+/7��k�q����;!*E�{0�τ��T!u2���ښ6��|y�N�摐ѽ+���]�DM+�v��<�O>\�O��ޫlv�@�k-�m�
��eΝ�Ħ���Rˠ�K����]:͉7����3�)+7�T�[�����z��Z[���l�@j�k*]?�
rT
�tu[������F��vE�k����k�Y�lY�\س�
�Mk�&,���)���pZ�Qj��Vv֙ݡu��=0̞�M��s�?��������3�}0W+:u7\���4��X꼹�^��a���	���zb씸H��
ofM� s��z��)u,<�.5���:a�4�9����Z���2z�Y�k�G�mN�t-O�SM��H��#EQ8�7�=YAM�)���5!��2[�B}~����%�/�+���Stc�@���V�����{�3lKW�ڎ�w��M��s�=��D���~1�{-�V�<l��廒'B�m�j�V^�5*n�ʦtj��p�#��D$�9�Ht��-VQ(۞��{lco1�����[����/��:����f��'�-���ׯ-O�ݴrm��E4��
͓{�-�\_�y	C;ʴrm�%�����>
<�}Ԋ��p��m3�@��Ď�γ�s���^�M��o4K0`�aũ�'{��.�n��j���ܭ�%�#A'�q�G����6ϴ�q��G�l訦6� .�8�ݳ������"�w)�z3�5楶����$����|hn�/o������O(�ؠ���앮���^x��ޡ1�՛��+l����B?���r������朥�#l������qÎ��G���Y�n�}�~�h�EыXki�,N��6ޫ�#OF(c�������ʼ�w�yk��(�W��U�/�H=�ෝ�k��6�kQvٜwq���ȁI��M�<�[iv]�'���-��g8�_1H�Fbl�_=S8�Ӟ3h��
�l�ʄ�@:[��P�u�*k��gR29��w�uJ�|��|��n��q��ş�1l�f��'S<l�{��r�sR����W
_�����iv�1v]�XC@�{�x�m��r�p�Y�,ɥ��4Ľ<�]鸭��!݃:ST�a@#ѽ�ބ�BR��Vq�["��36��W-�L�F��[;u����x8
�VY6{1�I1VO��n��٥qN�noT�o^����˄�\d����_u��ծw�sʵev�-1
Ozc#���u�%�q���kS�{%�Ȏ������\�b�(���ܱ�ϽU�I������U�{�6�.����cb�S ��,?�Ӹ��R��g=�@8���{�]'�'h3U��F�U�ǎ�-����ս^8�X܃aܼ �� �����k�^��m���gR��	9]K�-���a�f�fw��6���*c7*3�b��x�����d?_u�뷇Ƽ��f�r\R�����.D��a(�gp�՗��b+��x��Q=8Rl1��b9�c�7p���f}7��/u��*rw��0�ǿVHm�z��|���Ҭ��c�# er������d�
�;��ўv_k��M����΢C���6*��e�	�b�L|..�̰׆���I���:Zf:�}� .�;٥u�������C����#�T0a�v�� �p��o1v+�%ؔ��V7���Ժg: �0o����ue�Y��ƞP�ɨ=ú�y;js+I�x�eS5�L�bg�j4�'��a�s�j��y�OÄ���/z �0����u(�<�� =8b���I,�/^>���P�}�R.�<�{�&JW=IdϖS<M�]R���aó�| fi��=��j�����^rXn�YU�ƾFU�����T��(��L�l�� ������l"��O��������.f�Z��c\�1�&UmH�0��a+s(����S��3�R3"�δ��!s%n��]��ѷw�	}Т�\��]���CM�a�/'*�]]҅�v�� ����4��ĕ�/�������w�����ȢM�9�5I�h))���B�P��d����@~�w^1\`Q7ј��,��uY��ק�i�Tk��i"����^v��P�5�<��e�%��vE���f��M]�v��-�Z���oU�����Kf�7����p�6Z��~���N�������X���䄎Hs��L��s.]P7S
�e`&�{#��hf����P;�җռ��	��_;�_�kr����4��E7��`�S�+��Z�����m��]���)]�=�N��{����wdEs32�66Sv�%]��n,�>1��|6�+��O$�q���~$ݝ�V�8��®��qh�Q�W	�a=љZ�mV;��rREe&�u���!AO�db5ঌ�T��0Ì2N�}p��Fq=C%�a��6L]��?NdW�uM��3�j<���@9[��C�͆�^U���N}�/�f�5�����0fS�0�{]>	���,Mr��8^����o{���}�����v�i}Wy�SPs훝�ti�&�<I�GqW�S�-����Q���G�TpN7���:�,Vm���^�.T��"��f}�?������o"ʡ �2���HѼZ����i���\�w�>��uw>Se���X2w��jƧF��⼷d��-���6���@m-R-S�L��)\�pO&��3'�x�6�?I�zȫ��i�%�:m�n�=���C%���ȨϏ�UCr��:۬��Fi���V{t�7���ײ�f�Yhm���؛�����Q{.����a=W9���~������Ul��/d��*^��.���+�+g	W��;�Ǯt�E�����&f&�J�J�%oyY͠f�����Q9�=�A��G^�4�шF��R-9-�9Ĵ�����[�Y���n��'U.��9G��i����ܱ�]�7�o��$�]�WrW�=�t̜=��}k7�E�z�"'��8y��,��`;����h���>>w��U޽�������yI.4(H��f�v��g�A�����E�#6�,��+��5^���϶��������kU�{��WgV6��˪��iͬ��� ��pP�l50��d��hcH��8�{���Pg���#5��2��V�9����|_�nƨi��Z�O�=S�Z7.v����}&@US˺�nWX���,1^}m�sOj����tog-����ek�d�D�S�:��h�EOƃ;����ki�`���͚�6��i$�rɌ����q��]u){MӸ�f���w��N;�ږ�|La��,���Z̬&�wˮRz{5(���y#�8T���y�w1 ���2���\��9�}!z
g2��b�l�Ǥ�����387��y��0ܡl�E�(��ݴ��2�K*�<�U���Az_B��9:c���O:��j���ݭ��_fm��'���*��E�|
�3��C���Xݛ��-��ٝgce��|�lv޳�`�*��`�N��Yb�뺵�`�x>�F��"���2��Eg$e�ՏYB�����	�"��C��}��uN�z3�Ԥ�3[���Nb��9KK�AR��'R�3�y�fQ��v��)/�&�o���[i��k�Af���rl�wd����4�b�4?
��f2{����k3��lM�A��5*G�oq�B�L�b�
���ρl��Զ[���/4I}��M����9s��+��T���T��"cm�+��Q`��V]��X��j��*�����1'	�{�os���=��9�I1�]L�����/+dj"�;^=�Sc����.��L��ɺ㭫xe֦u�5�y��͍[	푊+9tm��^�Z�s(�z�ȅ���-��b{�M�5t���"�B�*��0�1)���N���Z5]�:P�P�kLȞH:fM��:�tv��,�̼A�f^Ý�I7�����J�%��^3�u��ˊ%o1&wm]���\��gg��״(�]Un�&m\�p�Ƒu,V����:i���b�b	
.�V���^
�]M�f��$�R��8o'9��'(v��/j�$No2��p�K"c��b��/c�ѹ�Z�4U�M*�X\���QN�| �z���s1�Ï~�Si���$�QͶ���.�W
��Zb�el��7��㘱V� ���E��t��{E�2����P����`4�����4���d�a�B�q�.c/���3�KyՔ����僦Z
���S�A����M��ƺ
0v��#R���n[޷�ۦ�2�j|�)s�ǁ�-R�"ZXӦ𣕉n��{���P<�=���p(�����K8�9�]�A�w2;ۑX��W`Q���U���ia�:��'��	�8{78_ٙ##I�m�}�����\b-�5(7���
�1���Q�E�v�}4��<8��/�L�;y�S�*T_y����r�
(�h/��4�HQQ%��3�������?�o��G����g�i/��b�rWs9��8�&�"��O������|||||}������N�G�.�3�&��Rj��y�O�����*�#O1L�m�x�g��������������=�llh+�M�6#Z��SD��//-�Usc:i��TEPRDUMU��O��E͆���	
�d������X%��ӧ��\�LS�A�D�'d��Y�4b��9���I��������
��(����4o\���5Q͒�֢*��ي*��klN���71ې^��5��h6�Q@�y9:L[��ۜ4�m�'��Đ>�K�jno^�rط���#��홙�u�nA۷� �,�Kɭ�����.��S�����T;WJ�vn������ ��n�x��=_���N߇��-��i���Й����3Zk+Ts�:g&�H=�s\��$�{��>އ�š�'}n�.���Q�[���Iy����f��5#�[Ȃ���[���'3�n2�ꦣ�Ǐs���(��j��|��]�7�f�Tu��G�Ͱ�L#𽸶�D�OD3��L�i`����D^�=63���'H��l������^K��]�Qj��5�<d��0�LM������bQ@�E�M>�����[�q��[�޽���}I���U�cz�
VeX|����W��F����W���ĺ���9H㥴��)w 7���]XYt��+�q�4�]X�b:�6�fhR�P��K2�-�z},�ýA��vE)ӂ���U0�Iy��ַ�#�0�4
��foUR��^E�t����y��B�}D��'��{��(]'L0���&`�u�\�n�8��&ƕl���-���Iի$��1W'���O�$u*#O� ��WX�{�}!�mu����-r��vY�}6�e�Tĕ�8o�����Y�����bG�㷝,A�j�6��ds}w��|<��v��6�æ.C�Ug��R:����)�U}q�f�ڭ~�9�9�gi�䮝��w��-����Ժ��zy�Z�W�`��By���|�6���r�@�����͈�����φ��S����]����4JL*kv���,�� �vPrw(� �8|���E�~�4�7�mU��onۑ�ڬ8��/?�{�A8=�{��.��]ʬ:o8�"�bl����d9ie�p*�:��|o?3:����{�} U��-�-RN�i�w�!�$��q/�mD�m.���y�N!}7= >,��O���۞���O,̈́�cDF�4�Q';x*2�^��sѐܥP ٻ8&�,�+�o�����(�1qw��Q=::C-v��7�)ćR[��8Uz�0�{�=��������������D�v��4�]�c�@k���-��������X���I<�_{�Зs�Cٹ�K��\��J�˽n�޺R����[���*o�4u�-���s�	Ϸ�2���.�;ݻ�:Wt�孝7N�(�k�NI|@��fi�/0�Ӝ97�U���Ƞ�n�E�ۗe�r;R�ǣs��v�����O�I���B�M���h��e���bBaBR�F��L$DGИ�I0V0�I6דe g�{�ӷ�m{�\�l��S���|�i��A�;Jr�ۦ��힋��kʮ3rY'ȡ�LT��J6���o�?�����/�k�:��n��M�9�r�*�v�W�xJW����/o�K�@g�*��$E�˔�&�d��!Ǳ���2v;+R��*nz��'Q�V��i����>=m��e��b���"VT� ∆w%��ec��gZ^^��]���f�l�7� �к�+(:�/��l&��5�\�m1]d[���Ͳ�����O#��ezق4�`KC�yT�`h�)���7���1XSv�F�9m��8.�E{��]����W�~�} �.�
����Ր?��2:�2*Κ�I� ��l?(�gcn��K�C�Ƭ�E�;ѩF����z�/��U�e �����Z�f4@�s���@�]r
s2��z7mv�����P7
Uoz��ON3:	���6.��xڭ������U���֢Ӵ�����C�0[�	N��9���8�%����}b��2�+=���\i�˖��^��d��I~�td�}1�U����d�';�NU��"h֓]�/�;ؠ8�m-�*��w��~���z�X�ھ��mZE�7^�W>3FB�8���ŸnN��3�C�F��T+7E�k���=��D�6A�n���;ǁP����Upڛh5��Wo�E���|���h$Tq�Z��f�ܯ�x���	 �@�e��Р��֏2��Y�;��+SE��ɉ�P�]#-���\�N�7Z��5�#Y�6�Sh-3��Z�^��\�k�[a�T��S0&o�!Z[~���U,�Lf����w灑�Y���K��ڔ;�6%�M3�<��EI��lMp��̫x!�� �.�Al��Y[���7l���Hk����r�ǌ���C�rb��pO5��@l��8���x�$+��Up�lb�������͡�����*fM�((ot���7�e�����BQ�|�ᵰ�6���A���.��{={�q:i{	��B�!������Qu��P�tv.�4��}+S��F���c�����Ď��鄘��L}i�Sec�g�T��d=���:[���H��|�ޭ��
e�8���J��g6�տ<��[O��:O��U�o �l�����J����򲼷qh9FCR*+�nl�����ɇd��>�:�[�=ҵ_���;OٳC}��H���t�;FM�IZ�h���i�9�Y��y��ѝ\e]��x�~��λ�v�P!���j�D�![#�l�o��!�T�ꚬ'"���ꇹ�D�i��Y��U��1m�}Z[R�/}�)UU` Sʛ�t���3��6�6�[��ks^=�Ka���C�b��c�C�\���i�nXY���ׯ�h��ʌ���h�w-d��4,���&~��3��}������T(��vq�nZ�����n����������Z`3آ\�&��.��*<��=��{��9�j���ݻ���4����� i�p�3^rfMJ�-{K[��%�ߞ<du�A�U���3̛��Xd9~���vn���O��v�ԕ��u��)��B����V�ӑ��Y����c�Ux0�n���5�DT{�����l6K�2#�d
�Gza��o�^f�c��cgQ�nM.ǀ���e��{�nT����\�4·iC�2�c�u3ݟ���o�#�o���Z��%w'�m����U^��њj�;_\K�Q�����e��=��c�{�,�Uz��b�2}��R��7�����2ȋb�S������]�3R.���n#��֎I)Y��_,撥�eSޏL�I���1��/�^����]�� ��Zc���5.�k��U�ۡ�m��k�|ĉ[!%}JK�=�e��g���	�F�_4)�J�'u4I����e��mܹ ���g}�e��B_�}�����*;/��6��;02�)���U^����PK��YHM�l����e<q�|�t�����m�1UOz��ez�N��)�+}��i�(��`v��K�ޙ��~���w[��ogD2��K_ac����;j��O�Yq����e��I����ض�WG�q�&n���ꏐŨ�o:#Վ�m�2��]ܻIL�����<�Y繙��ҍwj���ë���f������$K	k�u����·A�2y�dPH����,a	6�G�w2>����k�~�K�]��b���_�d��
Z 5w��n�1������h���:�v߽\��C󻷚:�k(\�9p��!��������EV��`�Xњ�n-��-묌��,R��`0IW`�+�^2��*ˢu�_���}���D�H��j%��|U��畺���KP7�+Z��6כ�Ws��QT�a�h(��$�M��{F���-eS�*�@���o���mv5ic3!�UЕ��e�O��q�rVW���K%�r&�<X�48�Wv�6�=��9 �9Mo���J���T�%� ��U4Y����N����5r3P�Ɛ�-�G`��4��l�@b�j}u_�
�gp#���8ː= ��ݟ0�ʻ7Kkܯ"N�O��k��� �0:LEU�̇��L�og�Ηz6�]Ҕ���9��c9�v�UIHI�r����3/`(s�������;BLM��h}�/�b��wo47��+!a<��a{��t�Z�6Ύ�o��u��>ن^J��u �'9�%뵲Ų��ۇz]�4�I��:�l��|�'f�u8�;�ί6���fS�u�V�^�	�Kv9�P�!/(P*�����O4�u ��F�?�' uT�����f��U�xv�~�>�آ�k��
�J�Uw�w�� �M�iUɹ�r�fsV�� �5v���AF����-W]���*������n����Z����-t�D�#0J�<�O�v��h�D�du�dF���j�g��ykZ�Ɵ����4���8U�\I�E�j!�a�M���OV^�SD;����a��K`і2�`8���e� 9�rfV�0�bZ���۔��u:���*��͖�ܮ���"�':GI����g#y�M)7�X1��L��� �m�3G�*Z���g�����N���K(kmy�rj���l�M����d�)���88�>`����v��Wy�7|v[�ו:�=@Ҹ���d��_ƥۡ�C�����^t�V
��s���hl�"��$JN=�{�.�{��ዸ��],V�3�-���egL^Et���܅�v��]�C��;��Uj)��[
��NM6;^c��F��؎���P�+|rD?��x��y~=��%�����Ww~&�+�ǚ�=���QQ��^h:�l�E�^�Ӝ-o�q���ǡm���gvw�z9l�^2�k�W��kpN#*��r׾5�6��n�H�K(���b�^�����j�̵�9Q�\Bk�\m��N��l6.!���E��~=�.h��N�m��ހ1��B�wjUV�����x��Tn��5��>jp!Rʎ�i��-�� 7��%���n�7WqwvM�L�w//M;+��3����9>�[Րc�HϚ���j��E��5�ɻ�*n��֜�{�;>� ���F:;NSd�;��6��g��n����8���y���8n��Zg���=��m�rD4�nr7���y�=~J�V�-;�2@�̝�GX1�K��?j�W<=��ՉjW��1��I��6��NlG�\A��g�/2P�o�V�^+!锆�˦_2C0�)����Z�9�Y���¦��q�����:+	+��O���Gr����g])Z�Q�^����8�-;]�d���O�����8��b�\A�^sc+ٹn��y�����|25?L�Tʚ����r0p�i�^R;$���df>���۝+���ߖr���י}ߧ+��3,�%��}��<�D�"��b�.����i��v�il�󳎷AC��ms6(vJe�M���KD3� ���y'��Xs;j�R�A��f�سO�:�vB��(T-�h<�n������'�U���p�w�?���,S�/=�m���2S<���vܪY�E�nok����E�E(���^�)�@ϸ�J��֫��m�a��m��_��'����7x����nA/K�~ N����*�XȨ�\��ݏ �Q�.��]�g�/l�wXԳgMKߑ]{a@�|Gg^9+R�����m���vMj���w{��M�4�ʢ�kx�ޟ?�+����+�t4�ڭ=��(Z�˩CF'L�Ϲ�b�B�OQ��vG%���n#w��M�>�Cr��eANl�E�J��j6	��=�N���e���-�(s�[�p	9�m^S��0a�Q���,;/�bUV�mɻwK���ٔuJ|C�{�g<b��ԡ��LuUR��ŽJg0��\$S+K��Yw���"Q�+]��WW�����D�e�a�Պ����
(S^�O9/Z]�i����4ՉhR:޷�GR�@�ɥ�;.U��/+!�#�s�e��j�b�]���X���ʄ���%fW`�̜�(�ݾ��6 6�y�����-��g-qz��g8�r6��t�W�ѯwP��R�}:����$��5�ڹ<����ɬ��<�TvsQy�l'�9&�D[0�FT�ۋ���;Bg+BC���Ds�4�gs�U��7�%�jB_"e�ܚ����z7�udƧs�Q.�!vS]�ufND���C�u8�i��{t��a���c={�˨�t<p�/w�L�ynF]�֮�ky;���
�wc0�y+(�3��4��Y�5�|�\�'�.��FE��Cp����wT�tE�#�KF��v*S�*렃��:kڛ+�ԣ��%<MK����7P�q�Pc7v�L��XV�=�k'fY/�j{�J�a/o
�ݐ�S�\P ���o&ju̗7Wet�
�}k*���1ۘ����0���0�Kt����8�VS�l�p��ꌤp)�;�3,Ƃ&���&�A6�D!���DR�Jnq����,��]�զa�`��0P�OMO��P^)C�g+����r��^�B�Փ�T��87�cU��j�t�e3J	$!���.W �=��JB�Ae�zZ�˩3U�ϗD�&�sSCSK�R'2�y+��o��X[e^��0lwD5rB�AH�9��.I��cjgM�~�ә�ƪ��v42��)�{C �F7�E��-��b�ᮽc���7hm���*����m���*Ë���nq�V4Z]�x� �B̍C��fd9;,�)I���m�\�j}˵Εb���hν��1�Zj��r�P�����9����,�'�S�6�������x�)���${��(]��fBl�3��
��_���:�Is��v+^�;�}��x�A1�l���JX�hO��z��9#]��T6������+����g[�|uC6��LX��dב]_*Wa��Jx��2ӥg�47����L�C���sq=�{d;Oxr\�z��c4��0��Y]�!���<S��Z���IY�V��kf�f�h6{��F�BAU�2���7��3�[x��Ɛɲ:�7kz�D�b�l�)��k�Kl쩻{��!�xc��,����1��1W�z��t~9-rh�����i�U�>Z"i��h�&y�c��l�������������������U7����9:9�p7,<�Z�����UST&�ޞ?Y����>>>>>?�����g�c�4?Kɪ�sj����N��A�)ѱ��<�AW���<|}?�Ϗ�������?����l6γR���㍇��*�A��X*�	��+U�;�y�W������A�UN�DSQI[Y��k�nq�6�P\�9��9�M����\\�9cd�h����:5Z��-�ZZ��Zh"lgC@h���h�l[<�F���q��Ɲ%����m��mZ]�U[p�-y�E���A�6���r.gN�jɨ���劎Z�RF�l�)Ř��<�-.���DT��ݹ?B���6�Q�z�Ⴔ�S��76�Dnssm�Z����c�h��\�O�>d�B��*� �����%��0��i��ҕa �)$E��R�O�HɈj`��b��gz�l��t�����cܝ�����M�Z&C�fE>:0۰�WX�wj ���CBN�e��C�o���M�:n�'�h�A0%%�e
��U�/��F�@�b(��	i��bx�HM��
�bPMB!��&����e���� ��f���\e	S̐�l��
0���ȉ�{�0�(*u�%�P~�>��:�!,@ف'
H��FT2/"܅S#��@���n;��%|��sբɗ[0F��<g��gj�Q�"^�-$�o�R}I�V�q��v/�}���3��j^2ʅ�1���L��ٲ+RuIww��>���M�/�g\�vI���Y�a�m�33K^��|�*�W�s��\ͫ�t �W��M9^��^�a7!��y�NmT�'͈�omMv��`�!��@��2k�Qj���R罛��p�09�����Ŭ�6�p������{�n��?u�W�:'�Hezm�5F�8��ê��r*��Ht��T/7j�9�Nd�;tj;�E��|k�m�;n`��@k�BYw=�{N�;x���a�?��Dzb����l*�C�x+�U�@�N�bg�|ަ�W׾��̻�Dc7%�rbn������_��6��-�S�m��v!L;5�;��70F�� W�0�~���2�Wfː���V#��sz�{��s���n[�����K��
�_9�[oKj�ތot���iq�U:�B����F@G-�E��Ub���0,�������j��)�����nɟ=*��T�pfd����8�W�\�$"�4weF��&�!�h��L�2�3�3ʤd5�ʍvj�7kz��z��_�Zgg��E5eۙ7xAت�3�a7s����u%���t��J������l���άգ����a�>m�<r�ܭ�gב^;u!��r�-E3�ыݔ"w.�C/P�7y�^d����[�^�U2,�*��`N�4z����3ڌ���6v0��T�*<�+��[�9�]a�/�A�u�TPמz��g2r��>�+X�Snd�������[�g��H��jf�zk�"��� �n+���9f��_6�l�$�G��~q���# N�Y��-9W��6�{���s��ɶ��u(i��j��f�	��#1ڍd��)�	2������[��X�f�0fw�:w��X�a��]�@��@��S{rg��ź�a��&="ؘ,��x�hۣX(>c��df�n�Ͱ���ԞpF��xZ�ia�d��$�T��g�V0tR�f���k��x4C5��,!��:��g,N�u�S�[\�j�8��p����_:k��籸zJ�W�i'/'>Xv=j	�-^V���������i9�y ��x�q���4u���p��aӨ.��rz����LX�<����x�b�F���t�zCr�T�]�;�n6��w���U�4�Ǣ�x�ً͵b����wq^3A)���T�^w>�m1�r���:C�ǚ�ZV"k��w�e�l��.CS�5���d���t�ng��TH��k�~����/߶����e�����:bga%vVun��[�wBV1��NO��� wW� ���i���ܹ�&����͛	7<���c7&�j֭7�Z̔��[)�e��6�d=T?O��P;��z�]��c�;��K
+x����~��ʶ&��ǣ.�)K���;qj�Ց�z�e���ɫ�m�TzV�~@rÝ��,�f{2��h�~�-N!wk�]��D�g%;�x�/+/����w�s��R�V���R��;�7O�6��n;��z7��ݻ�{:2wVo�^-��M���)䝴���^��nž"ω� �e~p
�}t�w9Mc����gs�*T�z�᥻�Vك�a��mI�O�u�.����;{Y�|���:4�1�ސ=���t6��t2ʍ[��Q�~�:]L�tY����y�d��K�^w+���g���,�m�;��齞�wP����"x�i蘊��������������c��Yi��+dp͇�o4�Zo�����ID\��EZ�2ƨ>őZ�_���k�Q���pk�w��6���?ٿ�M/ 3���1��g����
ԁs����|���=����ȋv������ZSN)���.��W��e�>b�Q_�U��mN}R�߆:��Zʍ��D��L֖45�̇Y�bei��EV��g��3^���t[�B�/�����vECw�1�]�.�\5wL$�&�U�+���̚'��:�f�{1Z��خ-�6GK[C�ki��ag�e0�Q9,���^~���ΗWh�
�NlH+��V�qy����O��54�*��.�ߪ��U���Q�i�����K�}��h�K���l�Q�!p%O�;R��k��tۣO#���s�d������Wv�G�9m�2Զ��b�k����i�M=|m�̃b}�9�K�G� ��-C�'��}����#�u<��x.m ߉K�`������|Nb!����1y6��2",��`���ޘ��S���꾄�����nP�uu���B�g<�͋R�a�,��o�����2�q��`��w!�]���jn#��L\�M<D�$	�y��sW%������׎�$۸('��4���>չ���N�l�&�'�f���(XY:�_sOP}�Oj���;�s'�5w9�t�y6�ڒ�Ф����w�-�J�H�gc[�E]w<Tm!�4�A=�}zK��R}�A�;(Y�G8��n�e�����{��v�ڶ��ٽДD��:�d�ͽ\S�J��w���9b��O�͖q^{�͉Ӻ��\r�W�(:����fv {�ī ��eC�I96'-�]c�r�]rg��v��L@h����ܽ-	5���mMɀ�r[9]{{n�5�1O�6D3e���u5�M&� ��l�R{=p��wd��~�>����43�I6>�DWn�C/�zW���^�{�k5�昣	�dk��Q�<���P�ոWJ��Z���f"����Ow7�{/_�'*�B+gv���7����=���31D�3,�*��ЙP@Oہ�7{ĸ�U�5({�36�&�&3'ڙE�����:CY��W�3���x�&��M�:2�R��ƈ��FG��^�R5�"�x�@�+�^2<��P�)CS��y�:��u�6�
�v|��b�����S�P�6���f����es�R&'vo+�s��ǚ�
^�!s5K����b�C#�t���8E��;��J\�h&�ᜃ+�{@=��g��ח�:j%.��C�J�'9�/�B(�	��'�C�UL]�������5M�ޙ\�����b}�ֻz����8p�6�/���K2�%m U��k����9R�Bz����+����/4�;�1�XR��r�A�Z�[�;�-o�)�޵��;�a���n��v���8�9-����y]��]YC����'n��GNܳ�]X��Ҝ�]��{"  ��3���/��*���U��Q�5�7��C%��,������i���E�T;5,�JF�P7S���s)��)J�՘6�[F��w��ؗ']gA�N%X���u�/��:�0�fDZ����Z�HD�H�e�:�$��.�vn�w#MV-a�3��{��͢\�gI�82�;v��1x-���3S�2!�L.3q�%3W��^������{[��dFD��~ �X_��W�3}���:����� u���M�W��<�{�蘌�v���M�D���@8Ւ76ǯ�6�����(���s;��u�'�����=S����/��L�4��Á�;ih�1�*����t�7:�By���~�~���U�q��ӎd����y��Cwf�w�*�.e�Ƙ���&��#�]�N����3Ƅ�Q<���n[���!N��V]�[�����
�bo�{U4��e{8#�ȠEMGE�����Z䈸��}�Z�qK0a�@�*��]�Ygd���w�m��{0<����}���'Y��ڏy߆�4�:�N��L�yx��u��>F���������ps�k�� �*�����-���wE�����ݙ�B�e�3oO�g.��N/���ZCv��7t�Y�&��h����{:�=�� c�tY]�*���wW_�>�) �YtΉy��99��Ƽʲ��r1-�b%�.P�I�8���.pz)�n�����W};�.!�۽Cp�g�oo�#-#����bUScN�Jo
�dO��Z4�:\���5�ڋ𛞲�T�A��k�k���J��Z���ʮ,b����0��ֱ���;À�5�A�����w ����v�F#г7IF�{��c�nU��j�̝&���z��S��#����G�&�:�z�E���:ձ*ձwF3;�{� ��v�?8�X�����h�J��cf�Pq�|b������9�J~�t��d��8|�������*���'�q���g	~"�z��S>�&Ev2�N�H��l��s����ٶ0���!�;�ԾŻ����XJ����i�1��7�A�oNʂ��j�a�q���ŪZ�`lz�]��*�ㆼ�xΓ���c�w��2w5�մ@j ��a� ba���Vf��Y�y^m��$�fx[Xϛ��j'@�����w��x�ml����(p�	l�gSY�+�w8��mu�2�ճ�.�uTY�� �t���S��.L�tx<jܵ���A�p��(�6�.�2U�7�Ѯ��
�Q7�1����lֱ 8�a����c�u4�Z��RvD$�ɂ$q H^�H����<t ṟ����eώ�/BeM���ƍ2��K�/uVʽ���t�ƓM>Y�>ᾩwk;"�56\�S=Tf���涋*-�v���GAf}��($���>j�V�iԍ�ΐ��R��{�l)]ٳ�wA��5KM]Z
hqZe����ʟ<)c�k�g�N���������S5����U�ޔ�����e��]tY�TI�v��{Ml���q� ��jz�8ux�ՌJ+��΄�ġ Ԇ�t�P������\�n�x�l�x�d3ϙ�6�䷳��4�}An�v�۬j��+sZݔ\�f�X��*3UP��s�� 5�M��i&�`'�6�J��&0jӳ3E�w3]����׾���������`	|����VDm=K���J��vK�y�T,%��粨���m�U�ZY�٬��)<Y�o&r7��h?I�����:��_J�eYZ�A��=����i�e1�ܙ����U�cJiK@���x�F.c�=�E��x��/W�=�_Y����K��k{Z�oZ��!�D��� �ar\k�<l������a1����Y�?V�)�K�Lu'���[���-Ӗ��&�:n\uwV��T�9�������.���Y靀�f[
��e�5�[%{�vZ�kwA����֓[��Ϡ�����_2T=ca��GVl�Ыk�k�:bc={-�A��� �����3�@��ȻI��WN�6if��=����[�]y��ƀD��ʠ����e��O��v�l�E���m$�t�)��s�3����"����6|��G���Z��	�����yI���9�av6�Ϳ<^�bQv�7	�P��YT�|i��^TMN[�U�P:m��qx�aU���������f�Ay��	��غ���}����w.�S:-{/C<��{����R�IU�U2������.���ϻ�-���eP-i6�wj}>x�+[� �CK՗��1���"u����1i;[}aŠ�� L�ѱDf�W�vP�\z6�I�z��o�Gŉwg)#�X���K��r���z�@ۀ�A�6���V˜ef�eG����Bo��(��h�u����;�ou��$��f��m>���y��էku*0�,1vsDfkt���ń�ݸ;��T���6��LmX�,��q��ڂ�+x���Ω�ۛP�f����B��`}�T�gE��F�l;Z)SƳwj`�wZ5��4�q��PR|�)Ѷl�ǹ�<R��e�ĂJ�龩E��I�o�X�/*�>tl
�+����s�p�p����4+p˒�f�j6����koaw��-�3A��.����-��K9I���'���0�	]^_Y��RX�`y݂E�O-�q�:��G*b�����۬\�ܖJAۚ�C_ljd�IK ��G3�f5ټ��C5'TB������7M�%]՚��jZ�)����	�̎�e�΁��'!�t�.o�����օS1����	��p��Ku�28�A����;�-��Y�ĉ �{o9u��ސ�L��t��[��x�t%k��7(N�5m�'�q�<������[��k8���58�ɘ-�f5g������9�3	�8�4�����|�Í�-��U�*"&��nц7��ҙC�������ޅmvG���j�m%��IiH%�d���s#x$Y�%��a/$��@��g�l��WWM�t G�cϏQ+{��܏�]�8�F��7��jꢻ�C7QW�o2R�.�n�֟i�2
[ɍ�"��7V�&V�h�zܻ6��/��;ts�i��Lq<pb՛��q3���ï���kk�Y�
H�T���:�oQV�Vr�f'Rb�u�ګȯ0�VQb	����s9��`[�p��;�(���f(aΡy�q���-2�b�ɫ�ww�VSc���FZ��90���÷U��o^�o��8�dY����J�[��oc;��y��@Af��z�-����JU�k��a�p���y[kA;�(jOv6����w���gh�tťƐ��\���T�3/Rӡ�'GI�t����a�Oa�i������%��-aS�YNj <U^1s*J��.�%��⮨�e��EU��f(N-d�X�Nk�7Xρ�J�i��rݣw���YeX��]\�s��3&�:�>W���uh��<����Dt�۹i��tgi��c�&q��Z�q"���`Z��=�巩Jwx��c�NBN�����V훮������μ��[���V��nޣ��[|8�͵^��g-m���e>k�;B���X����lX6<&vm�U9-|��Vc���Q��m��񧬮մZA�O�^ �b���my�M����
ƪƫ���Er�h����	�Dmf��N��������>>>>>?��\����ݷ=^\���k���1�h1Qb�QIh�űՂ�������7��W5��!~~�������������z�������Tb5DA�b��G,�#S��ր�cZ���"b&��~~�O����������s?��߻�Uͩ���)Ŋ,lF��!AZ���ڒ��uV�k�F�^�1�ܱ���l[QQV����(�l��7��>�<����X�:>8�5���;G��X�gUA��[ih��V��j��rͷ9�:4^o|�䔵�bJ���ː"�"ш���{�*���l��4h4���N�cMh��F�Zq���h��ܬh(1&�S�ѣT��4ꭚţ�妍�UG-�ch����69�������V�km�,^\A�V�b+mF�kUX���]z�^c�L/-F�c���1�����H��($�K�㵛��{nvN��s)�Zڗԙ��e��ۮn�ru�(;��\	۝��އs5	��d���*q;�w�0;8��W�B��G4�{�s����3����+꤭����N�t30ex�%�U��)�WD�A5FfGY��t%���r�M���e��ؙk�gI�<��ȸ���z�����	�օp�S����,���b���:i<��'�z"Z���m6Ϣ�Y��T��]�5�v�{�����z�c��C��vh���3	������S���7�4%�L.3�q��Oow��!P�]������D�KV�̳��²{���aoLAF�����y�����#7[�T�u�M�� OAƬ�f�|���G���APbU�\��|�Hw%zvy��=�g�o�w�];����q���AӪ!>�}uM��T>�핥[�r���&��ڿm_oS�%��s�~�D��	��������"��^ش���u^���^����	����#c�-E�@���R��mZJu��W�c�Ɯ�F��d+�u�@~�.���qݍ:�-���ʼ�\�P�S�f���pV���L��e��,�_�������n)�մ:�ȟ��go���I�&�L��~Pٲ뵧�@_LM�.�/{z��(�1w�}��OW<�H�A��-�᩵H���S]us{ �9���l��xy>.&:�D<�������y�yw��r�hJ�<��Hu��*�=��A�":S_Sl���Q4�p���\z�4(*ј���U@-�[Ď�^��ofc��ǧ�z	-U�񣦡竍^ǥ��bG���n𫺠e��nۨ��c7R�	WM���1���@���p�ێ�k��J\�ػ�Գ0��]+�o���ޢGYe������@�>+�FR;L�����t�M��<��o"�����i��=V٭L�/�d��-8�-8�1�}9v�7X;�6Vev�4u�ǻh��^�Z��7<<�e	����)ye�0x��d��[�<�]�L�q���Q��n t�1s`|+��_��e��?s8c��7Z�ɫp������<��ҵ�5ҁ�@T�u�*oCN�㕓��wU�YQ�Wվ5��X��2iU+S���}� �.ol�Oa�ă��G�^��fWF��[Գz"�ơ`�=Kbq���ƃ���]�Q���%P����6BZ�o�~���;ݩ��d�1�T-�<�0�٘8`|oJ��[��@q���Չ�+g�3`>ܜ���ɞ��L�]�2k����#�����"��5m3���9�S��dH���ߴ�v��h"���~���.T:��b3�d�����
�>���I��.��zA���a��9�̈
�zE��z�yz�a�r5m����Gd�r��4d7Ph��v_��B���+pd򚛼���Jk@9]n�R	2W�ppxs�d=����)�m��Wt�*n$�A�:�7A�拷y�u�S9�p��vY���.-S6�u{-�C�%���#5�\=G����[T}L���Oq[D����F�����om�(���Ť����;>�twJ{���Wֲ��	�]���fv�Pjo3OF�ȉ����u�l��UrU�O�oJ�~27�-��O�-_m���8��ג�!Sr����v�-}��g�7V74˲�H�YG��!�0�`NXOi��e�^=��ǉ&ݛ��qr��*��[�與>���Rm�����p������[�B��z'����wS9{����|�6{j��U{��1�> {��w3p4r��zm�)_<��K�M\�������T2r��[�:�����`���E�*�]���Sa������,d04�����N�滼rjR�-���ޮw�jJ픕�Ƙ37V�� 2�أ�[�R�H5��|6-�q��:��%r��	�� ��y�� fc9G�;I��n>i�s����U�^�Ld
1Vl��N��VȺ�m�qO�����\���?��<f ���ζtV%sZ���]�����?��N�3~#2��U���|��׏�ƻ �����,���2.Sa˝|��J�߼��k0�D^��/��v�@����>�c��C3=�{#���Zf����5����j��I���@h'��ɟ7Hc;��{-�r-�1*2�F�W}��x~z^�����37���i����6����nK��3LD�e��{��S.�?�D�:��O%m�ٶOm[
�0����	��f!U���\�FnWv���u8>~��������7�b��S8.�t{sN�:Pk��nc�V�\:r��Լ+��|ٷ\<����_Ulo�z�΂���C>����z����U��H�s���*U�X�7QB�j�[�����"��%�S�9u"�`J9"��"�@�w2���^q˸�ʬ�;��	�x��u4�0g�)o\�WS�.T
aL��^�:	�&>�K�%eV��Yd�7�.|� f�N�C]�ux��7+��lb9�δ>�� �k4�1y�w�;�x�q�\�[q;]�ʲ��33Z[�V��e�(�`pQl�������J=x��L��"/)g�7BY`���q�^��u[�ݭOA�=J�{*�oB��t�])t��,�y�n�z��v+��{�t5�w]SD�@%y.�� ��CM:�-��Fl��b�l4f�@��r�sw����nYt�l��9��}��L�]~&���'l~N3�w�5"c�w�X~QhVt���!��*a��dOo�v�~�d�A^V�#Y�p���.7�����FW1��<w�}f�j`��w��O^*�������6��'�fm��V��5r㫧X6z��㨻\�C�w�76)"2�N��f�5(�:x�����c��{�7��jJF3UT�[@��}�M��/����k��n�;�%�*Z�T�F����i��t�cم]oi��͒��4��Ã�0��Ϗ���
�w��Ye�b��RqD�u�[%��`R]8�i��5;�r�2�CsL�TK���SW�Y#�����؁ʅuݣ;f��m�f��ċcw���(ъ�;�Q5:9S޻aA���ǡY�D�]2oi��~���j����N��$P���M��E�LMuPg����*��c�j;*⽜2<7��Ռ��i��͹�@S>�E��*D����n�Q�=g�[�/ǯNmYnl�ն�-���2�4���׻C��l���T���e�K8ev$��J5�Y����2�j�����°�4]cGأj�z��V g_�6�R޵9]3�ܣ�%��e#d%�X޾Bb��ci��K������B����\�U��ɏk�����Z��R�N�*�#��hӔ�1�PRئF��ә�?�8x�><�4�����&��P���\nYm쫨̶�	�X�N��])��-X~s_嶗Q�� <���<�u�s��J1���r2ɞ�& �/����[���Chg���d8�-�������U3d�3w4�J2�t���Z��3V��-[�xyff��줩&���ʙ�ȦF��oA|�H.��e�bݽD�<�������Lj��Ʉ�7+;��!E4��;���|WqOn��V`#\6��g[��3�f�8.mq����'avU�Tm���Ֆ��G�}�7'�ɹב�W�ٱσ�	��c���6X����*�qֹ�p�����וQ����㺨���\2M��3W�'=>�ui�5��g�M��Wnݩ��q�&;��qU��&_ِ���N�:N�
�X���T���U?'Pw_��T9�U:����݃{lN�7ƃk5���db!a����j��d_-� ���Kȳ��[M�$�C���>d*=.�솰g�'��)�#E�u�x��F�k�3})�e��WI,�6f��N��y� =k�m�u1k��f.���R^�2� q�<o�I������87��3y�c����B^Џ��-\Omۥp>̷�	���s�S�5�kW>Z �YsCp�;ග�4J��f�3 <���~ �;��+�gi(�XD� lZ�,�e�CY�\�7/����ڎ��ܯ�ii�g��!)�G<��Q]�mr�����> �jÎ��Ǽf�N��F�R���j�T�w���w&�_+�7q�>�D�+/~��5�e�NU�\��rR��qb6���B-��f�stas�|L��fnG���z��f���-6%��g)�s��]��c^^N�����ZT��ܕ�Y���\�1'��5�2��e8m�!t��gvx�	�R��hһX�v<�K�vG�W�g�i�m��͙Y�ts5�@�l�
?@���2y�>\�-�;~|��*�Y��+Z;+;����3n�K\b�D��J͝��%~��Y�/YL�"��Lf�<&2l�D��'��y�foG���^Tr�v
�k�o�U���Y+\�ϭӡ�3C��G�~���:�^�=HK�c�.�`6(�X�㑫�xh�J4I�r����]y�6 �뿮��(=��9���cI�7CIH�v.�2�K���N��C�ѱe�,s�\�@[��_�5��p^�(V���p9�YOIi"{�y�m�!)�:���n[oL��3�Zz^����Yc��{f8d�!�|;��,��ʬ�h�#;~�o�,��x�/�hۼ�I�� ��z_�e�CvÎ1񡪎]�b�Qҵ��D%���xnda��6�s^$H�FX�'b�4�z ���| ]Ҁ 8n����*����r�g����jB(d�bGm'��lɸ��ĸC�/K��V�>ѕ�>��k��P��19SU��Kb�xS�1�U�ϛ�6-f�<���t�[�&�㥬�ӆ*e��?V�b�S���,�ck���^��uʎe���=�Kcx.ɟ�x�ˤ5�5�-�z��ۗ��c:J�l��e{��p��*��̪� �V�`S-��0�~�{#/tՎZ_���9C̛Tt7BK
]�A�X��B %[�/��W���
\���9����d㌫��`@� Ը��˫�bGx>l�u;VA)Wv��(������ύ���d�/$	\D��X��)G��ۼ���K�Y4@������ڃM�^�#�;�k�xS-��{}2�{y�A2�;s�����l�Ѐެ�ǋ6��c����r|F�x_	�VCgr�畻bJ��S���}���9�g����>3I�P����;x��tӺ�ժ���Z�n���U���In��������������Aw�^S��vZ뎋��RSF�5�0z���TF�s��Oq3�#����HM��f���[�"
.�}��@Ӿ�L�.6O��W���fXtx�VM�c���u�yZ�Ϣtŭ[k\�h�#��-���WcK��<�cI��;��=�y/�t�J�]�2�,p�c�q�f�J�7\6���kyf�Cn�h>B�����K��cq!���ddq�D��L���tO���8j�x?�6*U�*�ҽ4櫡�(�+~�m:���]�7��c�7 :𰇦Ǯi]8���"���FN��X�j.9Ϲ����1�w��U������~~_��}A�x" 
��*����O�����?��������c�N��y��Cz���<D!���B!�!B�HA�%BQ6D��2)!�)�*H@�0���� B�B���!�T� �(!
��@!�=�������@>B��	P�!	D�@!T�!D̈dPBU �$PB �!PB �!PB �$PB �T�@!	T�@!A�@!� !	�@ BE � @BQ � @B � BQ �! B �$s��@!	a�$�HBP!��$8��HB9��@��$C�"C@�$!
4�$�H@$1"�y�B!C ��B!0ʄ�B	H�4�l�dR�BQ!T�%�b hdB�HB?����pz�=���� QV�PI�DB*�~�����<��g
���Ͽ[��O�]����r$�~�l�n>O� 
��������UE��X U� �����a�<�S�3:�@{v�|-�q�'JT6�C�K���C���6+��E@Y �D!%dB�U��H@��I`BB)D�I� %B RA �$% �H`FQ!%BVE �! �IQ!P��IY�%@�HYD�$V%P�RX��IX��J$�I%B���D�� �
h�(�T�! �@ �P�D�J��"L(R!!L�A �H�@��2�B��, I ����!��K"H�� BB�2!"@0	!B2	��1a�O�����H�����Ң�
c�7����/��� /��x
휨��l���f�)h��'`K�+X9����(" �x����?<�4� �
���*���a��?� A�0��H(�� %ӽ$?�!�hZ��XO>$�41C��8�x�*������" ��AT��vߨ9t�Bʷp�@���!QȈ����� U������C��MK\M@D�St����.]pB|�@����0|�̙�C�?������N�_�UQE�1����QE�����{6���PVI��K�4.��:�` �������f���)DTEE
�JIP@�*U%D*���TJE��*��)I*QJ��@D�UUJ�IR ��QI)Q$B�*JJ*T�T�BRW�D�PQ *�QE*PR��EHU(PT���
UH$�)R"�%5�bRJPP���UER(E(� �$)R"*P(�DR�EJOl�H��A)!T�J�"�� �
U�T
��  ��@�(k3@}j�fm�݁�J��4Е�5Z
���m*�E�ki�E���0֍��(Ym�Ma��d*�C5"RR�!(�T����� 6�P�C��B�Χ ��P�@(ܦ 
(P�T����)@�a�&I���P�[	�cI*����M�
�VԦz�B�KXh�T%)"T�JUkC�  �h�Y)�3RՁ�j�������Ԣ�iR�K�4m%54e���`����YShi� �9�U%e��0��%�QPH��MAJ[   �v�5Vk1�UP,�T�T�j$UP�J�F�H:�Z�5Y�%*Z���4fEI*��J�	U ��   ':B�Vj0��b�V�eJ�Vj�[U�bjh��l�J�*���X�E5H�j4 ڂ�T�*
�IR�G   ��EJ"�4UZ 3S *�����	M(HSiKUR@�����IM^ƅvJ��K`�ʪ��U%	T*R��T��   �P
լ1� 6L �`�  �  ڪc@ 3@(��  �V4P -K  5*�֪TT�U�
�%#� 3�
 5��  l�  �  �� ��Bh
���Ь� �cX  
�� ձ�F̤$�B(�R�  #�  \�  -�  f  ��2�  �� �L  �hSS[B� UPT*���UB"J��  W  j`45L  ɚ  ��  L�  �� 4�  6U` �UX  ���R�  E=�	)*�L@ hES���C&@�O��(�  G���0  	4��UP� �Ãs�����˛=H�3hI�����i����N~���k�g�_�7~g��9$BI�gן�$�I<���HHI$BI��H����B�0��I	������n�����O�?����f��w�=3),e��Ly�-�`F�9b��Hi���H�ӵ//B�F��U���҅5C0L�V���v���'�-�u(5���3[X^�(Q��o\��w1A00�ܧ�c�W�+�<ChStM(MD����L!gVLaL;E50�&en�N���v䈭׃~�w�N�#u@q�F��3W�oV^��9.�F���V�&V6��)��7N̫�!���[�.���6(�F5�V 
ݛ�#�.e�-�ɫ�b��8I{ E
�i�G��kv�UmmZ�ofZ��z-i���&���K7���6e(n�f�S/#fE�co)dP�MM�;
` ݦV���X��U2�F��Bm̑a��Fc"m[MNkSh�>��u1ٻ��	�q�h��t����j���tR�2嶅ǘͭ�q�*�Y�Z���S�b{�.H��a�*X8�x5F�䵵u�H�r��S6��Yn�56���nֵIHT�W���v���\�J���v	�B�w�w�Պ�b��`K�]��X�$��n[ӂ�e��lM;�q�Y	Rj6<5�y�7��F�{0�+&`V�,�R�ǚ�<Dԟ'��V��.f�Q��1@�,R;p�lݺ��c�t���f�{fī�,M%fk����P�E�F�	5+�UȢ�;Q�d�yn=*=�5�b�,���5���!��G@�vDŒi��<�	{q�j�]�i�v�T��)�l�V�V�͛�{H�Luj��{�^�N�Q���r&��(I'w	U{�ɚA�T��Ym�4kvů��
�ļ��]��f`�d�#x�C[s'yMRզ���,76�*1ݍ;�GY����k+(�n�v�I�V��U�D���nֶ�)X.lͣ7Hw��Pꍔ]�:
�-�����y׼j(uXCJ.� _
R %�I�-b�8V�b�v�B�ICw�����,��!F$���,7�ɠ��E!%�Z�E�YD�e�@F�>�]9,f�h��N�U�`N�QN^8��Z���	����4C�`@��ִ˱�%�HH�ܡEmǫ^Ӹ�Y�Ye}�,���h��4�1�L^=qd�fmXɳ0���ƾ�!N�-Z���<4.��f���-}w�o׎�i8�n�Kq���q����3vʌ�c���k;��j2�7h!�SGE��h�����]��toػS Q\�	ې#�ݬ�~��l���c�VęEd�j�P(��-�-y�6��r��уiLœP��,�B�i:�2%���P4.�B�kn�Y*��VJ��/(*�xƬ��]�lm�*���yLR� R1-5�8%n�O!�q��Y,h��Ui����^��lZS���^0�Yկ)8�ǧ%�ua�W�$-K�6eiS��iB�!�SE��5�P�so^�N�Or�%i�M:����u�[L�gLSt][˭���l�x�ܤ�q@�Xo�QelDh�MA�!3%ʻ�7Mn+O0��I�FǍ�ד$�me�Di�Ģ�	���s^�!�ݙ�eX+n�֬�.�Q����D����5qR�7Y������|�mn��lJ	�V��nR��ڎ@J�\�ݡ�7N����K�%��9�F��XWI��<�t\�7 �I^2��1���$�L^Zr	 �i�˴k ud&���f��Q��'urDq�ے�f��2��t��"���S�qHU�#n�
eU�X����I���fF�!�ꈶ�5Wm�4�:@����}A�Y;YI<B;�AoY�M'Pyr%5�a�S]�t��;cF�V4��V1�^ �LI="���M�bF�dt4e�4�͠i�u��e���BE���WL�Z0���A�Y�,2�w�^b[���Ԓ�� M[���Yx�3R��E��y#"�93E
@�M8iۑތy��4�,D�Bŵ�+n���Lm'�>yZ��҇
�i���u^��R��4��Zb�
��z]�����2�ͳ@
���^n�B]�`�ih&%O4fФj|�R�D7Q'�J��n^6��P=����`[�j]'�3�tU�N�P7�th�K{I�)����5�q
��c%���2�2ܷ�Hn�Ɓ�����[7Y?3h]�R��Gp�XgU��Y�Vԇ4QJd{JR���I��.�: 5��[JD����V�՜4qB�%��6�T��D	)�]i�M�(*�aA�6	��؛�/2���k�+ںp���`��*�Ֆ7L�*f�-$�Xe摗t��G(<
26�;���h��bY��N�0f�-���J�2̢N&��#�.�&�FZ�Ө����Ǘ���'>P�d&��:���nb��{A�@�{N�/(̬�w��siQ�n�Q�\�{9c��^9!6��Ø�
Vj���֩�����7e�b��UI�K���[�D���,i�U�S�5�K*@�D�dS%\Tg�Z+&�oh�l0+L�H��qY�Ј�iU�U�T�����К���0����]�",��$(U����b7�F$d,�Ǐ&4Y;�s]�Gb�ڍ�le�R��U�A)�-J��t'P�+U�n(f�F�x��x���{�ݕ�5Q�Q�f
1�jV��f*50�OnF�Ձl��ymfi{N�28b���wSSm6s���RN�B��d�7(Ӯo��(ѮH��F�^�h4��0�"�W@�]$��h����liǡ�.V�a�*�S�N�c&�4��˰�Ke�@��X.j%kɟܭ�!&���RSI�SL$r�bYf3/䥊[6;bG!OoFӎ=�q���Cc�}��u�ع",5t��81Rh�Q�Dm�p�X2��Q�����Yuom�7ji�i%�)h����N�R��l�2Ŋ&�h�E�6��״�)S�;,�rڬTUe7�u-�����g �Pg%�M�{t��a���չ�D��BUتtMқk�%���[����8��M����Y����4�n��ä�շ�n����"��ˇd9I1��X�U��jjWo@�FZ��{�z��Af�iaȰ�C$n�``�`b���H�����h#6��r�.�8>�$fP�FX�m�l�������/��p���^1�#���2}Z1�ït�&<l����&*+n��^6�D��k.e�CC�$�ʍ�m)�#FmY�i:CbN�i創��ڙ�%�hܤr�>�q3�(���\�,���.ee��^j���)-��)�
�B6���Rcw�,aT��a��eL��I�v��`�-f��u�&���4b��pi���;6��(!���2�P�H͒��xp;�����L�yx�l�f`��R�v�M�M�o$��\�]F�I+[;T@ѷ7KT���P��1�ǡUڧj�gFD�s.`jb��v�Һ)%B�1|�З���XĦƬ�NYJ�]',b�afb���SqD,*�K4���e5�x����ٺ��	�6aV2�һ�S���R�+Xaj#n\̗9 ����C��9@�U�[�挅�-<j5��Ƞ3�-ոo+C�2�c1<�Sf�O�,`�NnZb��1n=7�B�^�U�,���/j݃��R:���m�5y�9Pmʆ�nm:2����S$��56��/,깖i�����;��:&� �h��B���Rx/6��n��(-���v�B���h1����md�dm����Y5��VV9YX�)�ؐ�6��%�5�]�i� )K�m��P3a:�R	*�W�p3��	�c. �u��oԡ�7Bj�L�e�#F��U����F���>T,^&VOM=:!wI�}�=�Q�Q�aXt5���dEJ�gCz2���"Z�C7��.#�^���Ws�Y��שR\�N�1�)�b�+��
��܎Aa}�F�m�Ӑ�%dǭ��e
zi�v�R�^��Q�{R�J�i��1E?������b���6�+Z@����g5^!�:�,�W��SRm�5�rԺ�w�����
F���\�!pb�����y%3n��X�G-q�vki�	Jƹ�m�	,O�Ź���9��#��,h��䥻�MKBaRR�n�5�GJQ��Bq�рٛ�2��ʺ�WSQTѰ�nԡL�p�p
Ai���5�Fl�M%&�h[�d����������%ӂ����([�x�~�6𡗺u�q��\��:rkFe�)��im�Zܚr�I!�V��J�u��t���͂f�C-f6.ė5�oi�B�M*�*͖yV��c�Z���YnQYr!o���Ն����Xq�E[� �z�Iܥ@j�Ӳ|�Ո���0�l1�Kt�oHU��IKFihi�*��82��X���{� 7\�Z��,@Kz� VD�l5�ZQ# ��Z�o�h]m��*�mŠ�������=Z1�L����>K�uykő��(�R��Q�"\,$���zN\���2N�����j�m�k[X�Ƭ#��{��V�U��SMh�g�ZF�t<,�
mZd�XE����f@���ȷb�X�HQ:WdFӻzv�b ���Gw+3mض��R{�^&�j��g]8���Ƿhܘw���x�AL�Z�O ;0\�Af��v��إ��V�Z�.�R���.!ő/����tL��x(���D3l;r��V`�1YMӴ�7A]�hN���h��2Aj�����h��CH[Ec����1cbOD��aE��%�QlYk65uw��S��&���Z;+�N]�(��@���K6T�KI���r�&Nm�I��р�Pm�wg��3CTj@�3�K4R�Z		D�:y�W�P`(RJ��@�զ��W*���2��%i�ZX�ۀ*��F�����
�X���!�{mFʓ/�3ɱP�p,Շ.�5V�T�I6�;��ne;#I�J��zf�wVQ����ưM���͵k5�R����kU�h���ф��Y�q�q|����åK�n�S�X.Mn�K9E֍r�)��	\���'+djޟ�]�8ѽLVLf&�$��v��M"�@M<��1f`��Y ��q��ۦhT2	����Z�%���y$Un�?��N�+�[Hw�e�v@�'B�:��mc����wV$�h����Ğ���Y5�F j����Q���0l�%2E�ʛZ�e�	�LiZ$�&�^�L�)���NaKK�1�'�l�W�k�e-R�ZI�J0m\�qϮ ��*�-ܔpw���Z��K��݇H�y�Q�ĄHi�In�l �C����ɣo�,`*�v!2��tՀ+4f���d-����IL��s0<d�+.]7�A��Q�
�C)���hi|����`��U�5f:��l�U��5� .eKf��"Q���u�[g�D�4�����md�k*�%�1]��ȫ�Y�Il��&�5N8��Q��Yz�J��J�6���K{hw�73w(�ȍ�U[Jм��!hQ�^��z��Y�k�&��`:EO��X��x�A�f�Fl��"��E�4ڧ�M�t�Ui�w2 ��5���2�	u�k����2eԛGm�Z�d�Y��6�T !����qփ-	/�ͬ���k �x���J�$Y��n�X��-���R��Dʼ�%NU���V3t, x��[ɴ�톊���dS9��#�Gh�tJ�Y�h�!�D&-��YV�J)<��7r�m�-k%j��ӑ��V(x1����R�,B�ຌ���Yt,�i��	��A%zqT�kH_�'D�mi fѺ�h9J�ߊd��Z�P�ô�ՀA��b<R;Oу.�é�pVU��jE@�s P�0emY��X Į��U�1V,���l�����\�ݥqZ�'[CU�v��l��
S�F*�Z��K��r\9�7A:ʓ��rD^���+i�`�UvNȎb;�J��n��
9��f�P��$H
zoc�Dnn��5�n��ȹh�u�g�`��4ռX�V��m�j��P*Wzi���jAJlY���le\��a��`*gJ�%,�/Q;�>�ѫ��0��n�tS��W�Wn�*����Z�aV6�m���h��X��W�Y�ۺ�3�$���q3���ڦ	�R��53�̖	x���d�^o#E���↱nPTF�Vܔ��4ʳ�
�ci���U�ķ��`�K��Z�v� J��"Jוj���6��n@f&f���bAҐT�<�wv>��	�sS�i�3��#�`�IcB��k��v��VP ��R��v%�J����K����,�����>` @�;h�:�V�e,���*�˷��@Z
�E�KW�$4���:֓-LuрmkR�[6�Y�LZU�MS��/+^8� ŰM�)9k/.���8�����f�� ,ZĘr�[33(�C1�"E�g!fn�`�m��B�J�Kd�x7EC2ֽsŦ�#�/T(� ��3hV��!��I�ܢ����;va�f�������W�t�R�^�E�Չ7.)��FԴ�4M�����5D.��eލ�8(	L�x�X�4��i�On</h���.�
�`�D6�O-[�s ǚK��k����Fj�W���2e[E���S)RlP�۷v�ӏ��R��[�w&ࢾ�n���iG31�W�1�X4l�[�샶oD�((����R���4��Rt� 쑄b�-�P�o%֥��:(�x۔��$d�� �֪���F���a��՚��l:8���j����v�<)�ӡBC skU]�I��s^_��R2����Zcp�0�/nYr[�Xn��n�ƻ�����C��.�r��N������?a�J�5�U��sf���e�<r�a� �*�Լ�EC�8�s��h��.wWnPl�:���j�3��Ydhr���wR�ʙ!�}խ�{1ѕ֧=C��ˡ������<)��Jj�����%�-��a|��d�/��/�u���$Y�w��v��|R쮐���e�d���^��f�^V2�#���̻=�`�%w:�V#lMt�N��������C>f!v�=��!/�8;.aL��2�t����E$q�	�ed�ZN��9l󷫷O�`�0��}n�P�$�j�Y�]��E�hI�j�A��^���%i����ʟ,s���=�Tt!����+��u��n�qt�g�b�ʫ�b&h����Z)�j��C{��i-��B��m&�wĂ�z멷��m_V�������:��p��\��u����7��yՙ�(H.�Xd`��Xe#!����7uS�.�e��o6ʥ]�-�H�7 ��z�î=�)U�r���wp�Y�5S� �n�1r-f�{���ݕ6mJ�>v84�Na�t]cέ\SE�i��+�p��B��r����v��V0�os��Bi��3�.W[�)��f�D�����H7Ýάv���+���sxk�!8�x���΅W	��'|��s��K��Q�<2��^���s�w[�Z#�9�V��" 
6^��]�bݢ���K�.������jZ���8Fm$z��G0�14
:sZ�fa��^���{6��pw{��G,�a����*l=���T���vٷ��s+���y����j�;d��S�^��3�W��Ӌ/�: �da׷彖f�I�:�
MU��ռ7jt5���olۗ���ՍV�9B�������y���]�V�����0]�'{:�<=g�B���\nJ�F�b� �LYS_S J{x�N����ug|����u���6��"G]�t��꿻z����Ʊ%������Oz�Q ]��OF�Z�Nko��Lx�gg[��Ax1Tc�A9��GW����Wω�^����:��MB�C���ۖ+���L�4���1�2؋h�Dm=}�-ݷ���]��������tt+k�,Lj��@K��*�]��orF͍�4�a�x!�f�����q�^&C}�"��H��[)pܾ`�E��u�um�����R)���ZP<wM�+�� K��O^�h}cFk5�)EV.�t�6#���r4�L����b�F��/����J�y�Wy��.^���OS+�per�2�wwt����d�R�	9��]e�Gj�m�X��j����sL˧�)>&I��sL	�e-ӻt�4�krf����{�sT�ż����������8��ON�p9owRIR��5�hL,��K�p��.���ލ��9 �ڧmp��un����j\�K���}�~z��F8�3��a����wG���U� x�x봥C*m�qeR�0@����ʰ���Ѭ�ۡ�s��݆�k�4nru�.�s5���Z�л&_K��F��B�H���zMG.��r�ʵn$�u�q�l�'Y[��Z9z9-]�yv��6y-�k�ռo.����.T�{���Ӓ�}�RJ�=Y���3Gg�W^��M��
��nM-�A��T���*INاf�Qǻ�Q��nt���j3J�A��٘��ʦS.��]�
�Ȥ����;g��8�x.fP�$Y��	�N�����엦���)&��������p!v�ԯ�F�
�g���p���;�z����H5s {���XB1�У���;5�;��_R�Lb��Ƈ`����[9yF�\���0������I8�8��M��̙F��@x3f��q�Y�0XIgբ����t��2�2�����uW^�Uu�l��r�ҫ���p܇�o�o4���*��� �;Y)Ju�V�7._�Q7R���ux_����$�cj
���pu��M��U��2���b-�� �}�oms���R�_F�N���]S�
�F����X�ʡ�`,ҽ	P�Vr����ѝ:��ޔ�ս6���垕x5Wy��ʸp7;���x��s�囊���m�b�	�fv=�K���Qݖ��>.�y����ZΝt��O-D󍋏�S,o2�Y�Ue�wcu��{�����Xyt����ӭ�
0���m��vYs;pG�f�K6��b�;���D�M�ہ0xR'l�3{D�o�*]�`�&�P%�u�5WP��^�-���/����ī��5���g�1Y@�9C06��>=Ô��A.�#�M���(7Y]K	�D*� ˃8$"��K����A>�s����Mf0%����|�c`����<��eɴ�f�I���*���W)s���!�9A��<�������9�b��N�8i���Z=޹����	�?QYzSq۩�ev�w���͝�j�mL�)��]�.�����,�8��|Q4��[�ܮ�&V6��B�P�ml$�B�Ű9\%ѳ��LY���0=�$4�WE�Hv���)�^��](��MVq�Ӛ���[3���J;r��h:��.����Q5׫Y@��>N�	۫n�\�O�%���/U;iL(_��B�h}�--���bSF�nw\��^Q����T�K$p�9��[�`pKwA�nQ�,mV��C�[.��٨��k'[�S�MlțSC�z0��M(�k�=,���j[K��t���{�I��r�5/��e�Zq�T�ו�W�7X�X`��YI
K�>�M���,ӝz��\C+�$l=#�ە��7[P�z0T�4��U���"�kjDh��+�Է�[��v�K�Ռ�q]�-Hy[*��s��W��ĺ+��^H��s�}IR��wce3�L�rм	B�Eۤw���F2�ⵉl���(Q��iGO�c��a�LH����O;����T�Dյ�b�:s���s�OnR�c�]=;�7Xu���nv�-'�-<��ř�S��S��72�"�kN�;T��}���:W�;t_e�hR��}�*�u+"D,�=Go�3�:�^R���,��q��c��`b�T�n��"������\�0k�͔S�(a�T�h��w���\���������=�â	˘�'��c �ΕgF�]G�g%qW��̅� ��n�7Wׇ<�GH^��wH�D1�s6�%8^��k���v�!��e�\v�6���B�ڻi޽�9V�usJp	Ǆ{����n��wt(>�qβu��s����O��OF��U�i"i�8��޼iH�]Z���*��qi6�:�3f_wQ`��8:��7����*�T�&���'��r�/ql�������Cr�i{ݷ���z���ɭ��7VV�(a�1mNz�b�S������;RM��Egsa�Yۗ}	��;�S��;�����2p-��8�;�t�r�oRvM'ۏ3�0.F�3Ivb8z������Ү�9r�]��B����=�zXӺ�/��5�B�r;Gc��0�@�t�1v�MI��R�Q�1=�Y�:��	;M�ᷯ-��ܝv^�Rk�}�q�u)Y&\�}t�����ntZu��o��X��j�;�Jgi��l�Z����Ö�w}��t��%��F�{;c����)�}���S�A�<,�*�-�k&�\_�,�G�9�n��x�S{���R��+u	YH�Yp3��ۑF��h4N������;��U��V��wq�{մ��d����}��:�w� ��^7�Uς%������A&K�e%ʵt(f���5G��M&q������7�o�+�*u*_p���϶�m*m.�0>y�.����r����^�� P&�o�[�W��w8�S�
fu�H���7*򔧃6;V/��ؖ�f�]�)м�0Ru������u�m<���6'g{��=�t�El�sm���_p�5+jW�Q�9��C�;�I���+�Q��������$���,1�N�z�˷gj�:e.�dvko`� m ?������j�]x�&ԫj�\�*�e�x`MB�-��h_6]����He.��oL��h�
��ks����3epޫ��g��hs�jYr��n�"�+h�z�v��&� �r�*%� �_h�]NF���w+�v��9m��H�Jͅ�q�-�GJ˃�n�h?[��΅:o���ZM��+%m��lӫ�A��4!|��A'qR���s���I��禝L�{o�m�:��:��ρ�\�W2i���s-��9f�Ҟf�9=/=R�[���evmw ;�7���!�9�*�3 Xե�r�N]�VR�b�J�i��H�u��7��/E��o��!Pnp��{�N�c���i;���cAg5�:�F�d����#�n��q����<A�8������ =5s�CM�P+t0'u���Y��HWx�vZ9N��[ҵ�D3Z떐r��Ot����h�ր���t�����l��ۂC�r�
�Kub.S��X��=�n�j��1;�n"o���x����`w�	eə3{:�]d�.[:.w#5����5��H�i����[���yC;o��:���[O���U{��y��V�߽�����/.[]��PL��=�y�۷G,��0�+V�V�7��b��T��6eq��}��:<���z�����o�fe5L=Q.�����`+wh���$��C�@�8��JŦ��'���Y��U�<��7����e��tx 5E��ʒ�ZW�+�*r�ovO��Э��|z���Yyr<�n�_d¬���s�.�ZUո���kG ��*��Ύ��-3)���[2��cT!M�!�{�:�:|�����^T"S}���
I�++&m������}�*"��5���G�oN�q���@UޱI�U).�V�Q��zx[/�'B���o��XR�-���6)ngU�"5f���4�g)��.5��C#���9�ĕ��/{H���T�ti�殭�E�w�+V�n��@l�N`t�F�L]�o��z�4��2���ƹ�'ݷu:͗��ju��]Ob���m&�c�-�+������^V�d�>q��GS�ݡ+�F��mZ�r� nk3�cƯ����Tȫd\3d��f��EAox��gw
��Gw7����*WoT���5h�������z��@��3g78P�-uX�,Sl��K���u��<ؚ��f�<,c�c���k�۰>OU��9y\�Ɓ6��L��݈�a���O�:���S?��.��i��׹4�]ܘn�}�[��U�-u���G��o���i�*�@���:tܘ;�B��� r�΀s��E�R���+\��i[D�}\�lh���\I�	��X)��֝��T�Q�`	��_c��<�����K�/s�Ǔ��t���%���t�Cx�q�ӻb���2��mLX���nm(��jԡ;�θ5�FT�z�t�M�7 8>������Z-�O]̆��SS@N�c�1d��o��q��>{9�e�i��������c�9]��i��[�֒�ײ�����MԎ��5;Vq�K��%b�����o&� {p[L�&st޼����t;�*ed��jWR�j:�Y��ӵl�:�y���}��3򧜀���8�RWN�o=#�4靨R}��3a�y��J�	'��u$��NNH)w����wAyPasj:t��K^E���6 ��޺��Wj1f�ej�b�
����_Iz,��I��GG�Ӽ��Z�»����IG6"�C\�0٩��۾q�4�*��{Ԉ�R
�����=P�ݧ6��l(�w>�b[��#F4��w��ҧ5�ݪ�)�&5�{`c@�Y6n���3W$� <�Ʈ�vqaө4s�'gn�.�r�RV>�vVV�X���k@#�D��j��r�?f�II>�]�vvf�y�KdnI%ݰ҂�	�qR�]3��N�'_]�j��5O)P7����g�q嚩��2��ahiH��āsnQ,hr�<����/r�ę� �)B�������\��t̊q����g���]��\�6��Ȗ�%wևf��y>�J7n��+�_آ6�3���y�vZ�y��L������$��H�����3X�7c��]*�+�a��]h��(E�5�ߊ'(��b�c�aQ��\e.��zrS.��9�+8��F��P-ج���ө�݃-�Uu��;AȔ二@f���\��EJ��b����S�)��F�q�e#[&.�3m7P�d���ں��lk���P�Z���]�L�cj��˄��=�&g�d��n�Ƕ�g���r�R�	�;�8iа�f�VX���z�M��,�0n�B�
����s%�)k1��ظ+Z f�_2�2T�eǶ��y]��#+9#ܫ��o����{\��^��������u�@IC�@u�,�yU�Mt�[I���Fd��G�,y3r�LR%�y˂ɺ���4��M�F�8ru�y7�ڐ�v$�����M�y��Ʃ��9r�4�A�P:�л�L�}�UĨ�K�Gm�ow3�\�ݩE;�"G%C�ʾ����U�b�9�E+�d��v�|�ڛړ�@����Oo�tF�E��e��֭���$s��@������2G�p C��;��m�$I��������]YGiYǩ��c#x����a�P�9w,f<���<��tm3׵��*������@ⲓ��'!�U���q���z���r�!�-.��\��kjs�T��.�
��]��d�y�r�}�*oY\:�[��V厚�;�)�{J�>)dI�P���U΍�~�ێ�]V)�F��	m�&��z:��cWq�[��;
�� �J%rN|-*Y9NR0�m��5�(QaL���
o�U���c
Lg.Vz8.�#v,��Ґsyw��k���yĹ�q���BBI$$?��!$�ߧ^�yw���>y�����y�7��
�O�h>��������sD��u=�3/q�����\GSE�4��ޮ�s�u���S��G)�E�V�+�F�Nψ�p�Z �n$:�+3{\�(us�yP��v��B�wQeT���-�]��9�q_]0Yu�٥��A��֌8R�	T�[�k����)p��[ѳk^%Yi1f ��vt�� �
�Bm���� V���4�䫷+7�;�D��.>Ȑы>�q��Ee�H3(�o@�Ҽ#xRݥ+)/����,�K$�������c8�����~���yս:�r��+�u'^#��Uk�X�CP\b�N��1ZI����+i��y�6
���#0�j��� ,�B���Y=B��jn]����hZ�w����JvJ{RKޭ�MK��V�뜢��o�lV8� f�XR��a�p�P.U�����L���-V��[�Qj���xU�8�.263(��6�� �Re���y�RPD�W)�]�ֺ3J�Kg�6��ji�8՘���S��W� ���N��U�|{[ӈ���O\�������ʦM'Ϧ��5��l|���[e�l=�u��.�jC�vڌ�7���њ$B�mQun����]'�����F�FUwE�e��(�]ڑ"�m^�n;��}�%"4R�ҍ>�U�9����I��գF��<^�֬T���&���%����&!�3n���{�.��S^�Dd����Թ޶Z;�E]�:��X*3or��p;�(��c��P�6�;C��"R������ ��q�%�(mk�eX�v����G��lm�O�_so94^<�Me��E@�v��n8�V�ح��,����n�Weq�5�Ŭ�ɹ)����'V4*�{���^��e�J�!�X���2![�'�[�!Q
k�p�Uc2��_rg6>���Àe6�g*웆Q���/��P�
�۝y�&����I
J�p�gP���EV� Ҿ�q�u���k����鹠#�$���w]9ܮ&�Ó��0����FU_ͬj��.��U`�{Y�6�r$�e6���UvJ�MR�z5�*�wV\����gd' 7Ͷ$��]o%�k��w��U����ɧ�,�HWZy��]�8��XB�QT�*�X���1�t�K�����Į���]N�G,���񮃳*VbӷA��1y���̧e���\d��Bo�ѻ,�_fQ�tB���0j�@0����GQ�j��v��T������튞o6���٘�7�c�W'JJ=u�N,#S��FB����Սvr�Z}�1�'d�\hs�#L���u��k.]m�ӄ�HF+\+�G�.���)����*����,�:��e����Į]���1H0q����>�c��O�_���T2���5gmf��p<�<oN����"vAd�q`q�a<b������k�n&�3)���j�:�(�\Gn�|ҵ�W��������q�R���3V���e5�4�겺��O��:n��~���wUk$$�K5��;y].�]u��:�(6��3T0t�k��6���B;ڽyK9	"�cb�
����C �1�)%��er#�캼Nj�2�ۜ@NuƱ>�熻�ջ�G|�8Y��1�k�.�[-C�陯�{��mu�9�I�K��w���>P�\uv�&�i��͢��t]��`$빎�ɑh�6����&*��h�Hˏ�V�boSD�����!'orn�������zpuqJ������,s�C�RQ
��A��CEq�b�^LھN�"�n�F�lP*��H�����t��Q����V�Q#[��R��믱�p7�7Јݣƺ��ՙ�.����V��Kjb%�^1�3&D�f��k�Q�ʩ��{]�K�A�hdS����QR�/#��)&�Ù�ޓVu��k���b^�Ru�%q�O]k�V{3!i���X@�c�k��ԫ��Y+tj�p	d�Dl�R��ćbETJ&yO�b-.es�UN�)R����w@>xJwHQ�a"A��5�b0�����5叭�̑��AI�s�Ԇ��9��Qئ�B�K����oH�x.���d��e����{*�o�q���EmZKR��}-e�9�3[��dfW!br�x�2�Cm�<h��wJ����fg�J`�=J��<'�(SgL3�ޞ�T-�s�J��ǹwԆ����'v�(V��x�oR�{j�o�v�
��F��u
��/u0�M|�f^��5�����ڲQ\�q8]E�v̹v��b�왛A4�=PʾLi�:#��3��,�q��қ	kW"�Q
�u��c�h�M�
)x��55��w
Z"�|B�r��f�r�zo���B�`vk̝���;�ȝ-�c��x�8mwN��'1����wH�r��d�-U�8���Հ�6;��iA��qtSw�-����Y�y=2�e��pJ�>h�B¹�.�1r3��T�cE�B��'��@�!��A3�.o^��9���J��L��MMGt��5�S��2�$jwWV[�q��g �%��g^] ��d"Mh2�D�瓫k�_+�R��,+N8{�m�� @(.n�]�kE�s�*�7�5��1��f]���y��^qpHqE|�;�N�g�A%�y\�A���Q"T���N��kV��c^,w
�@���	;�fZp�X�=H�uu�^A;m�X��i����v�rd�aQMPYc�vûxyD9bV�gV�U�_=	�(���ˉ��pb���iZ][/���QR����h��΢��r%�Hf%���Ga�5�,O�m��s&v�RxvuCm��!W%=sX˥c��KD��XE-�N��x+^]����*���b;��띱9ea %h��F��w	q�3u�=HC��(�[N�r ����s����.��kۮ��\/{o5.6VH������)�+Ô򰬕��[Vs��
"�WGs�M2���Y��;%К�AAF��].��E@)��%��F�"5u�IL>՝�z�(.��`R�"�]��9��mv*Uo#dk��9�e���3S����X���=e_S�1�M�Ŗ+��F}gNL[ӁIw9)�˽U�
���i��l �u�����a\�N��/�����D��zP��׬P���-�i����k���^m��i��-��Z���涥%|fj���:�,����2 ����:�n��pc�k�����ڱ���M�/�������fV����}�vs�C#�R�X���c0՚kN�r]*Y�/n9�ו+�-�^t�D�˻f�D����ʶ���,p6�˫����;�d�b�P[4cΫ�Tf�f��J����e�U��ެX���ꋔotXz��=�6�c�EЈn`�!���f:�v�B� �i��eZ��َ�.}u�hU�u�[��]�R2�T2p��-M{%��
���[��0�g�.���3s���ܢ���Ǔ[�c���'.r����ݴ{���mw�Xl�vv�ak�{Żl�\���:�S:�X�;\�d�@Z�}��:yw���g�:�!άc,�zKL�w���'������b&�(n+�͜/��*W*���j�9�c��t��r���:c%�Z�>�����^wR7�F�YpN��8S5��+���*��Y�����&�$��*���N1jb8ì�����Kz��euf�Hm����E_-�E���˙@��i���Ζ���Ec��Ne��'���> S�6�`�ɣw`O�m���.�h:Z�j�GgT�w3@i62�5����ꊏ	yۺ�a��Gx�T;Iٕ�EQg"i��f�r,�2\�B�ؼ}L����C�-�-��*���v�n�]�*լyf2`�i�.�-�ٹ�^p��uȾܵ���ф���%m�v(K7�
�5��G�N�\r���΢�a�7NU��oN8�(�*L��ntO!����w���:��˦�`�ٷ��;cf���٣KK�wR����0�67- ^�G�Ň�ɒ�%�GP�Ӹv7wy�gK[[�+Ygf� um�`j;�3�psz�3�jM�J�1�d����x45i�{]�3���C)���fd���/�kaJ�G�3���i���t�K�!��_c�v�j�a��2�p냀�	 �Y,�K6|��[�9�n$:����I�J� QHWf	�;&�A��c��u�oaz���R�7)e��6Ӛu�% ZL�6�Sɂc�+t�c"�IU�o��nZ�qs��R�L�:�цzI�*�_I����V*���r�Y�i��W����ʳ�`������3���9��
dE�W)�v[��i��PE�����p�m0w���t�>��[92�@%i��nm�W�)�po+W�-5}[k{����n��Ԗ�a�	��󱬭��e�~u˷����+�MQ�ζ4 쓍>����B������C}Ca�l�r�S$�!�A�֢0ҫyACׄc|�e�[�\�,��DB��%�ǹ;�Y�t�!�|����i����V��\�� Xe���äXp�:�d��o?��.-��)��(3����d��a[���>f���WX�>$ڕ�|%��(��U ��̧��u�f��+�N��n% �K�Ց�M��H�f�(Vބ�b�kN+<�-Ǚ��������q�Sb�]>��ɜ2ъ��b�/���(.��:is�t�GV6����H�x���*�RF�\��;�q��i1��e�pU���ڝm��Z>�*&	}�B]�;��Yv�4z��Û�[�6td����(�i�F���-��v=c�"��Ce���"G�!vuA�)α��Y#wrk
��������r�U�c���[k�
IwZ�z�e;��@oL�$/x�]%�36e�Puo(xYk[�*�9�w��t�ss��e
->�E�$���Ec�i��wb���6AB��am]�G�>1/Sx�m��YO[�V!��Q�Zl���S3�X(f����pC�(��V�,\�U�&�i�s�����E�Yʅ��d���ʮ�/�b��,u��&���g�-�XK2����ι�2�d�;����2��8dL;)���;1���C5�w%�g� [V�V�Wo���i<��Hp�7��f��,�M��ɳ)��ZV��bw��K2h��ǵ�k�!��p��D�w��(��[���k���s�Պu�%*���N�-+mwH4��ӓt��������V3�:v���q�y�|ZU�����Q��}\�C/�J������Zb������F�1�46��h-b����[��4ʭ$�Ti�eu��ç#�t�s'{���+*\���j �9��C��l���\�[՟<y�mwE,YRĜ���@])�y��)faD�@�#��p��lҼ��#����Rд�{j��e҃�����2����Mj��忱�At��|ۻ(�7KO.�B5/%�tx��WI3MgG�y�@�%��	vj0gr�t�H�.�����Fz�f�=qJ��@3t�xMb;>W.�������=�$��N�i��嶇}#qt-R��y�W6P鵝���g4�WW�GS��c�`'�t]b��	+�T$�.��:BAq�x��3k2���o2�|q7\$y�/�s�*˕�X7U�:�+�0��^̫F;��&<�����0��]L�kY���>;�al
Y{lJɈ�L���U�'����&/�Gt�� ��0*U��ݔ�֞��yd��/i&]t�;%	��K��s�8��(9N��nZ�;��V��N�P{����a�qF��n
f�[T�VKD�G�W�ڳW���TUc���t��t��U��.�j]*�Ԝ�M*���;�v���K1G���we��!;+���f�Z�X2b�z��y�rV�R:�+�[��hK=��5sl&�jn�p7��0�[���n.�TQ`')�frH9d9�ySH�zbMl���hm��� �kKnn��;�K8�R��F\��H�AlP�Xۨ�ueӗ��dJ��!7�b�����4벸�z�^�G�v�l��i�䝴�E-����zv�)ڗF�δi���d�uqb�B���0�rk������nn�н�5ڷgo�w�7m�U&�9��B��F[�׻��p^��_-�33V��*�%K��w�(cP+�U�������)3�dxr�u��`�qbeל�����#9���t]��ȋ���CK̫9�ΛԶd�����=�B�z,۾�Ⱦ�`�`��&I���]@�Q,m'n��/�`iU�2.��V1�]����,+f�l�g.;'5htL�6!���RF�|���d�z�k�|7yذ(�r� �]Q��pB��鮙(=�%�����o=д˥� `Ht�ӏMkfA��n�!�vAlCkc�ml�����k���;�9�t=K{P�����_u�@�'1������Kn�t\g�3{�*��+Z쥘�kDp�7R!.�'�f�2!VhV����g�4T����
�+���f�V{5�L�p��$"�N^ݓ��{R��7K��fFSԥY��p�1X���8�ȫ*�R�n���M.LVm\�q�2��I����4���w���빶͊USV�2�H��.�E�貕���]�qc:�|�������V��(=P���}Ǎ�G��x��6��3�ˮ��g_�Ԩ��A|9U�L]Ք6Pm���Ga-�fŕ��n�]����:uꋎ��
�qz3)&	�vޙ��GU-4��R�خ�oG9V�,�~�oZ�Wrp��}��0Ia�:��g�
ˣ֩[]C�ܾ����Ջc%�%[��| <w�nݒ^�g:WW���s�bشY1ޒF�+��ܻ���	V�:�kh��{w�����H��`W9�����uo|�r�}��;ktp0�G�t���6�2�e
�¤����K;D׹�ػ�%��c-G�+Ot�$2�n�A�SdIF�L�N�Z5k� �	'W 6pg7���ru�)����s{��k���/Ѱ�D��㕔�`5��iPQtr4T��fg>|ʴP�)��Q$^ue�,ӱ���h�l�8�����P�!q�%(
��,AB�nv���ǆRT���8���f����z,v�%fs��w��o
���%Ŵ��#t�����-�ܕ����y�r��.)�!c���E��c�I?�x��#���V+��Ve+�횮�f�g^-��>]]�t���h"��S[B�i��s��緮�/w��Kq$q�6cw���X��ZT��"�8u��]�֞��[Lwq�q[G�qօ�y�5Υwճk���":�|h^�TS5���;s��N��1�;Z\6�m��}��$�Zk��tZ�aɛ��y��R�K5v���=�)�ܪ�r�����+�K�!A�;٩m��:뒊���ҥ�<�ǘqwK�4!���JZ������!B�p��C�n�y-Yڱc�_]O���>&LuǱ;VX���}"� �o:�g)i���tk(��x�ÊJ�fBax�Dwַ8�RZ��X!�����Z_1%�Z��+x.o�3!_]Wӹ�4�y���3�<�Z�ł�X�cm��Ŭ1�*����LIR�ҥ�F��X�r��e+!�єLKh�m�c�l*�������mJ�m���ʂ�m��*�H)mU3GR��jc�ʩm�lزVFڂ�m��ʡP�V�c�J��18R�`,L��LjĹ�̒���K(VJ$kUP�X�m���ER����T���X"AH�jf\@��[b	�����ԕ(�KijX"
TYST�@�Q!�c�ZbU�Y�b6ֱ�q�Ab�b���������DeT��+PE� ����e
b�6�,�زh#�E�m�cI\q�Lr8���E��*2��++JYEj��B���C�iZ�Q���=��a&��'fn+�ݽ�U���Q�Ή^���d�r�L���9'�Քk:-�Lwh`���0k<���}�T�1���bGc��T����q��<Z���-֊��+�pxPhɧ�3�㽹�k��	�8F�
Z�@&��j[#��#�����Zj��u�9��+��� 2.j�V�(˪58^�%�؍
��][��e�������CL�Ps9)�l�����螞+�ow>Ϛ�,�F(�Ӿ�򍖏�+;Z1_�:�f�pD	�	_<ު՘JBD8�(�@gu��9�ک靓<�m���Q�����KO1�^)��M�R����գ�oǄ�XV]��A�H�_N��`juî5W�)��z��[�|0d^Y�`\2�o���g<��]Cb����`��hxS��@TG����Wӹ�w�e�h�� �妾��yR��D�ѧ�(�����1���\����/m�5�{W�Vf�j�a�'Q��m�.#zO�<(w�m�����~5�2+��*Z�S�u�3�9fvdc�	��n��Eٍ���Tx�ױ���]�
�P�H��s|ժ������	<����-fVw�-��y��a���k(]Զ��K�~�S��|��,�3<���=$AZ�aŧ�ݏ�=j�p&E�E���>����i��[�wbq��zrY4U�ZZ =hV���<'\�SN9�SE�̉V!�ybLZ��;c@r^2�u]�:"g��y3û�}=+��(g��r��5�~���B7J�E����U=�����-��&b�IT *v����`���ڿ���9�� ���ydA�s���Sy��M_\-�'��p7&H�Z�d���T.���B:��vJ<$![7�;\VcP�zRd��M¿��F(Djɪ�_���)܁?1=�P��U��}(N��Me�o[�~�s�U�9�^�"��tE#!I΋(X��ĩ�9"d�I75=L��<�+LF���f88���'br@�ՁO.�@�Tiȣ�O��G�m����)2��v��9�X�(�\�V`���|��L/�_{L�r�=(t`:�G�y���h��n�q/����զ�p΋��j��T�o0����ޚ%�)b�T$�5���Vtؽ�꼈s��%�zn��\��Yyy��+�[-W���僀
��xxJԯ�O�ʼN{�7�#9����z-��-�,�Īt�ó����ɌS;7��f���C*�uT�iںr���q��F[Ŝѣ|z�S ��Z%r�v(H>���
�7dFoE
gv��Dn6�`��%��)�H�l�.P,�tY[(S�۸˵�AҗwYCK���tBh�͓��:q��͆�E�탍g.{vj�Á2$8���	�X�XXG�G��ђ�U�R���@���r^<ήPE�q������í�kC��l������{��U<lz�6������)\��X������o�{fJr���`�DFY��x����vV�a���������K�h��:�vIJ�T�����%2S���+�,ͱ�����V黥K����p�%�*	��2���g����4�g�j%�̈,.5��TcyR���&��ӑUT��M�&�1��Gi�qV�T�@�0��̡�6�8�,k�/L_���p�+�7�6�)����GaF�Ȕ.a8�E\�1n'�bR�/�2�Dm}�c-��ςU��Na�f3ҷ+ѥ�f��xvc��$ �]Bd���@Jh�`3~���h�/ѵ	���M�]]�i�Y�ݼ�
�˞�-)5z'D[�rJ��h��(oƐ}��W�lMH]D�Uoe�Y\_��0�"W[�3#���N���� \(0����u�=%�����2_=��1���8��\B��p}��V�0��K1����Ó5��tm\���Ѷ��#6)Ef�E�� ,.|ҁқc5��I�Y���j�d
i0N� �d��%[ ��j�u�c�M|��ܱU�jkWE�m��w��ӕ��7Krvv\D�&>ʹ��r*
�:���@�MJX�[�vn���1Z�+,����Pʎ��Tr�x��n����z����`����Н�]��=�z��\wAt�x�Ҏ�-e���yb.��
�u���k���Sj�|��1��{;�5�-ܽ�&��	( ���e����zsrawћO���&RY���q�򭒺e���nrl�<�!:�k�٨^�T1������_��9[7��3�'�TįZ��w`�v%���E�I��@|�t�����CyG�$��P=CE�o��LV�Qp��Iv���]��H�Qq�#zn:���� �=.��)��_CW�"�;�.!7D�;�e��xL��c�A'��D �t�8.2f�� b��o���b��%���ѷU�ȸױ����=S�v����yU��J�5�%|eZ^ҫ2V���ncFK�F)�(!�ӻ��.�?��<3�}�>Q7�����κQ#���C��Y_W�Pxr2�9�O�o75�Q��X�h�:�cE�δ2 ������@.��`OԪ"h�R�ąǰ��c��5��>�H�����gq�i�/L.(�(13�]�:��g�(㻦�]�[����%��ԡ��b�]��
��9�ߨt�:�t��|6]N䨭Fޓ9cS!<7n��� K���] &>̷�]	y��=Fo0I��9�hSBs-R�F�j(]����8v�%�ڳ��s�*�9P�;�iB�Li�Eh B�آ�E�J��)����D��~L�oP�r窃�~��<�g8U�ƈ���W�:(g�1)4:�]��O�r>/ݶ�e�f$����:�k�Eg��{\T�0F�r�t\�h���s f�+w�������f�H��:�WˈQ}�!��DhVX=mހ����N��'�'�4&
� ���]9� =5lLM.��qa�ۈD�o1L\B}V�X;��5��N�۪���@p�X�Z�r5ᷔW�-�ds�y�/a�:*C6U����Z15�h��+�7����v*�����f?
�>x[���q��s��ͼ ��jޠ��摢L�ӣi<��q��s�:o��<(ٸ��f�KF/����L�N����H����(،���=�5]e�_�τ¦m��d1F���0U<��o��]�4��,�?P�.�E}g��cᯱH�e0xR To=�s�o����A��'�z��FҹI��G�:��*�h*��V2�dv�����z%�h׽��r�2���0��^�`vS�/6!C������|�0��z��]�U���^�z]����gYW�f|���Z�pˉ��u����żj�h,�ū�DX�AB*�~)�����GA�3PF��Z�)�(�8�*��1g'S�!�8|�Ƈ�?�������^?|>�O�����R��u��}~�,}7��/<u[<-�I����o�y)l粱*�꺱��%7D��vs"#�O��ϥ��5���ȅ�
��R`]L���V��\��u�΁v���xk �ˈmU�҃���ew1�b�1�۝e�F��ED�2�7���f�f�J?�i���xxJ�J��z�����3�o���U��c�[Q*��-<ҷ�ݳ1}�uvԩ����]<����"���jK>�:��#yn�8-=fT��$\;:���t[�4��/���f���U!
�t���*W�Q����nP��m^U����<�ɽBqb����A�s�+�ሊ_
�ؖ!�?Y�{�O�}Ṋ�X��`79���K����:�����Ub�Ϥ�Nh:"�C,Q�?��g &s
��LoP�댦���\�su:6L�͟�}P��sh�9��o.ɂUj�;M�Q�<��fVK�tq]DQH@��������
�ɹb���
�
Șr�S�h��Gv�'nE�PA`{c8�lP��-%Q�C���r�U xN�N^F��/�롛�gw~F���E����P;M��J��B�}�j��R|~���`�n��i=U�Wq�p.]�j:�2��Q�kT��WcI�ũ�vp���S��s��>[��zǣ�/#�4�F�z���F���LT�hlq�NFe��������(l!�6�֦,8U$2��'�{��V�{q�@>+p�^*a鯵N�5����Kj�,�cID�����4wHLS����N��������5�9:�3���|�=�}�@/]E	�	�ORxl�ڮM��P�-��"��2tƗ v��ʎ�䯰�[2�2Z��)��^Eb�9�=J�����<��9�ۊ��Ɗk(��k��	�<#����J�p�w}W�ݏ�9�`ǹR��qߔ��=�	��l{�>��:�)]H��Ă��8�af�y�BWz�TD�L�K����"qKg��5O��{g����T��q��+Է݁i�;ޭK�S�+C����9�1Qja%}��!q�,`z^�NX�w�l���3ؽ]N�d�|a�o�e�U[q|�-��[�׋�=n�i�Z���g�3�uw���<(��ǁ�|�����jǟm�!QN�ـ�Z��S�)|��ǵvU*�(qbM�u���E��>nu�v�!}e�o���w%+��X��!�%���W֧	�q���)w$^S5���;V�2�iC83$N�Prt��9�ΝoE�m���P�ۂ.#�i����r�D�2{��W<��ڄ��[%��Q����0�:�9*ޜʿ�-�H�́	��pU�닆�B�$$o���$ ���W��;��i;ۮ�T�@+;���W3������ӓ�^<�+�J���u�
�['����.Wa^ob��a-�� u�+�wA�9��Q,DkuPZɧD��'��%]�.YsKE&��)�3�QD��-������ATX�>����7G�ǵ]#P	���g`�R*O�t���Wx��c�n쁯��{%�'�h�¼��|,<�?��x\��%t¬�}[��ɜ��sT6�� $G��2�nA�M���
�ͦ*4Պ*����:��D���+�y	�!�]��o�0�hnfÅrh��g�aYߤ��A�\�l���v�{6����ڲN	%�s?E�뇈�2���}��7t�_@��u�eb�-d4�7�b]�r�k�uun����������U�K�:�\���� �"~j@�'M9����VA"�Zf;���a�*�u���e��^Z�/v킼�o�V+��30V��^a�+}�!+6�̬��4�

�����˒�!�5;���P�É��LE�:��e����G6��&����Tdd��O�Z�I�g(����a
�����=�4�K�������kz,C�����:R�0�,׆��|M1XMv�tlJ�e�
�Y2�����|�8l�T�7hMҾ�ܢ�7�=F�sG~7ꜯe�]+w����gՋ�Qn9���v}'Fu�R*��;�n���y��1���cR{lW���\�<��l�5TQ�j���v�''��fzpe;��`�ok�޳T��f���6�Ȟ��F)���[�U"����Yn5A����>��1Qe�`\�wq�p����
��b��%0R5�[�9�A�K�u��5r�k0V�$-��i�#ƼڬT�������]�zy_�.*�v�]��7��[͍wk�+qL����7��R4t;6J�`��;��ŝ�"�����!a�+��b��N��o��*QfU*�_$�m���բ���a��b����
�U�>��V���ݟ\+%Q��~����'�E}�9�G:�x���j�S9 뽁�w,��n�#�~�`j;[��eH��
�G
w�g���֕Ij`]s�u������Wu���1ڕ���m�>��h�0d�E�j����w'��h��gu��rt���tTo�d*��Wu�����d9|�a�!K��{�wX�p��[��Wv�����+
�L3t^���:�d_f�VE�V�Th� F6��ah���r�TD1Μ����1.��ӿG��]��9�/r�xO+`�}O8q����Tr���Lb�QS�۪�����O�k>G�j�4��y�33;�d�[��7�Sz���L���׫�N� ���1��t���y4%�GT�C.�r�3����7��f�d���D�BwO'!��O
D
�{l��F�t#'8>:�|*��t�MdJ��8���J���I�!���a�+ny�5�	�P�e��w�g6�l�[�����{Up����*�v�}�mq�^x0�C�ϭ��3�YP7�]��8�o�+(v���n�Ց�Z�B� �ı���CE��\. 8:<��v��:�7>]3���9y\��*Ɠ��c��4:��^�g�z*��K�W7Ώ�{��\�V;5/�����.�kS���>��Uβ���:�ο��l�82�=��MO�Q����k���40��aC�*7p�� �"�.ja +�2��6���8#i�C��ug�k�e]�������P@���2�ѳa��`}!z�{a�ҳ��ە��=)VG`ɽd�X$��Gp�Nr�r�.�[I�ѕ�v5�Z{�{~Y�NM�glG�©}��ʂ���d���w�.����}�
�I�cP��.�f�+@��6i��2�fӻ�LY�n���n�$�"�3 �PU� S ��ꂵL}{&��R֭mwb�FNTĵq[�\{s@���F�梱�x��c�0n��M$nT�Q�9��a�bY�ݘ�]��kY���$ڍ��7o�zipxHXd���'���U֪1�f%|)S��+U����A�י�w�+�e
IT�]1�ݮ�Zr��KB܁i�Z�i
���n��-b�kv��rnq㗥+�*l��-��镌	ǱPq�7�M7ڰnJVm��{��1�_W%Ƀ�CY�RE�%��w
��{!ۻ����wj��MO+S��2��h*V��$^R�o��b �@�:�������
���#@]��p�f3l}����Y��ț۬��.j� ��8h�]GY�Eޟp������-�49��$���.y�����)x���p�����8u�z6k���,QӤD��0�]b�9���j_K�O��Q����jc�W��T�8��:����ό4���+����˷�ڷqb�[W�e��yf.�q���/l{�l�+�Ww`&�9�ў��R��p�$�mfl��ǿ@Nd�k���"��L�wb�/^%��w��![��r��B�o�ִ�5�J돮����{:����gbq�<��z��9��;6�d�{pVoԾ�u��*�w�>�H|���b���r�EnBۻA�7��ٹY}W�]���d|�K�*�eG��
P(႟��*�Z�N���T�*'���bI]q<G$)S�xQ!r��a�m��zj�܋�t�AN=J��wNWeu�@�5J��u�ai4�X(ǃ+������fK�j>�k,C"y-�n�c8m�VN6{�0�0,V�n����6�%s;'��tڕʡ�TU��>;�E�QbÛ�TV��+�VU0��72���v�V�Ǔq�jw%����㋩R\�7��A['GW+�|�M��2�*
�U�dD�U�J���N%��{��z��#���ş{={�=��Y�w�J���$�8��8�z�x���Nͷm�q�ip��w1����,[݂�C�݊�U졣[�n�բ:���j$&�����RJ���u�O �쥻�<�ya��kUj�% �)�����Gv*��}l
=��p�+������v��%'3\�y�y{|5�#Q<��\Mۼy���,���Q�M��1�[<�i��L'v��	@b��-��ʩ��Q6��7��e4���1gT� �E8_v�nڝ���.�^���b�ģ�*Al�IT����,�2���֝#k2�������>}��5���	w�U��$Ҏ9w&��|l�W�ީ[���v��X�����z�"��VG��WEZ�{���{�=�}�q���T���j5��LB�fYۉlb��*b0Jر�-Q(�Q�
5� �-���FTEkTX�\h��\�+Z�F�X+-�%�XZ�X�*�Z��U�e+X��E����Ŋ�F��i�+J
*��D���I��Ƞ�D�ek(�0�����*"�
�T���+��ke�
����"�����Q+KJV���h6�"�&e��+#mT�Qc���E��T��Eb��(�)mKj6ٍV*�DT#�Ycb�ƋmR����1�h4KDF�b��"(,��1YZ*����DV)�r,E�D��:G��ݜV�aK��pm�(u��e=�{8� >��t!�R�,�ͬV��XC�s�m�İ��"s^pp����� ��L�S\ԕ�H*��2DI׌ě����'���%`|�f��u��=��C�*u=�����ۥg�*������1}���fL�6�����V��ܿG�"8D1 ��?`
�/{�q��i��wz�]>$|��Ld���-`/�ON��~a�l
���M��=LIP����zß��
��+�����k~��<~﻾�bi�(t��6��?$�K۴�O�Tǉ;۴��Y*��x�b�.d+�X�gg;�hbL~`_3"ɉ�*~aU��ǈg��>���鿱���I�y����8DX�,bOS�ǹ�@�>I��y��:��
��i�4��V��u�hLCn�c���'��%egϓ��ɾ�ɥf$�+>ʡRW��&r��H%D}����k��/�����f�z#���}�vئ�<qX��'�4�a�1���d�:���yf�1 �����lĂ���P'_��xk�O�P�x^���J��;�γhb|�Sj|t$�d鑾9�9D�"8��)�wT�H/�z�Olڳԕ�l�XI_ɦLECė�P��I��&��4g���/�>��
�� �ÿd�J�U&���Հ���5���o훉=������z�|���
��܊4Ì�1���|���?'��H*�����<OĂ��� ���1��C��O�T�Hc�ì/���=@�:�O>�M�ۮ��$D�ڼH�#[����b/�@ ���N���ٶJ�~��%f������5�8�y��m
Î$�����>I돓������&$�'�P��C���hJ�_������寷w�k�X��G�G�]���%};ܛI�+���<`x�=J���w�1���Xy��%d��h�ᤕ
񓉏���C��=a���Ag���l��[|��+^��j���f��G��@�q���偏��{���|��+&��>k=gP�����siP�
��=�~CĂ�3������l���mI_���=���Cԗ���&$��#�c��'���u���V4㬣bhav�@����mV
83������KY��AY���V[wu����Xi��o�QI��]u�9�]�w����U��o�i��mиѡ]��/��C'Γ䦴�y	�^�x]�Buw�{�Z�i��o��:�5�b<���w��9{�~`bC��kT�:H/��&%d����1 �a��揓�0� x}�6��u18����>֠,�f!����Ad�{�&����06s���Ag��1}�����km��y��g��I��+��� z�nÉ'�݆$��~\H|��q��{�p���|�!�>d�=g��2C��K��Y�R���u�LM������;�4�~f�*AzwܑM$��a+�'��xn͠x���[�O��1 ��,:�!�J��ğ!^'Xp��<��䘁���d�Y�%g}�bx}�	���M0�ɀySJiR��z�hW�N��?l��B�������i���>����4ʒ�$'�骤hST�q�T�o��g�3�'��4�Xq���:��m>�������y��Ԕ�s�} ��+~�LC�+�zçy���.ý�d6��Vy3�jM��!�|������ΐ73�i�2T��]�`bAt�e8�La��q��(i�a��G��=���_{2�������D} }B#��`H(k����x�����v�0�,���<��SI=B��;�d� �I�l4��R|���4�W�|2�&!����&��J����?t��i�
�����K��?}C�Dz�'�_������!��C��q4�Y�ְ�ԝB�7��?%I�*}�8��b<���C�J���ɦ|�&$��VbIY��7��7���殷�f��~�ob��?!_���{Cba��iO��Y+X?2m�{l�N!_�k�0�x�Yԙۧ�M��H/ٟh��>�c1�b�|�{ʾ�@"#����q3UY������y�����|C�m@�S����8Ρ��{Xi ��5�5�&!�[ϐ��j�$���ɤ:����z[$<C_���B��
�s�:ɿ/X�C;�$�+�t�����ư��������9�����8�R�{�b�R߾ޡ�i<a��{�	�>C��8����H,�����J�SF�:�!�ia�,1��Az�!��6��T��w?sG�d�Ag��[������\�_?��"���= ��n�TS4M�B���c�Z�ܽ�r+s�媎�to�r��^�����v��r�i����;4ve��7��%�gV�hH�������,��srs�W^��
�j���&��K�_[z8�;������*O=��V��'s]�P�J��u1�<�ed�k�a5l�f+�XI�/,��ٗO�
�X~q<�����i�>{a��N�Y7��VOn���uS�JB����x������;� �0�N��=}a�R���4�3�Ԙ����d�*��K���6��z�z�߽�*mT�E*,�k6��w��
q��&� )>B��g�:�}`T>D�͙����oy���Q�~�k���%�O�,!���P�#����,�����C�)��m �I�>�N��u@�{�@�i���}� Ă�w��4�������CR]���q%}KOu����|������>������m`)8�g̗W�>'Y2�=z�NRc>d�Xk��h�R
�s���u4��ǝ�i!�c�̜M�m�~�Sĕ ��/u�zs�����~�v�wߒVT<OP�t��&�%Ag�_&�%I�x��}dĂ���ҽ@���!��}����6��T:���~������{�5�'��g�{��O�?|/iz�wmlW�V������*a����i>LH)�_sԕğ!X^�b�m*OϺ�I������b�s�i���Ԙ��l1���ϐ���I�*O����}����������ό��^KY܎��
��@�,>eg�vw��
~d��fՀ��
����J�0*�>扶�o�i�-�6�~�b{�IX���f��<�C��������g�"&�̈́��x�{�Ny�$!�s�B � �t�0�§�I���x�Xb��{7�6�Ԩ~I_>ߺ8��AC���bmX
O�w���]ߐ<�6��++�:OM�1�2T��g�} o��a���uZ���8}�M0�0*C������?'��'�i�4��*��*��*��g��膚 �]���O:�%�C2b�Led���܇P�����刯���ri_��+=P��J���S�������� ���Ws�$��
ϙ_X���a�ğ'ɉ���)>v��T���Ud�+N�>Ci����4m�a�
:�����^�V5�#�pp��Q=a:��RYj9�%�LUt��N0	��3Je�l�`b�pU`�U�Y���-�s�\E��;]�#�5+̌N�|�Nv$�)>�:sԹ�嘒wzs�}Q����Q��ַ��9�G����U�mÁ,|��u�)pY��G��<�q��f���&2�VN2�<Nꆒi
���T����9CԘ�e��� }��`�1�GU�_�!�yO,���Ϝ��kn��t�ګ&�C�͛�� �h�Е�R� hts�Wˈ�t�V���r+{��-lkGb�#��Mu�q�2��ʘ���%��@x]y[���ZF���eW��Z{�zs�6��W��6�_)�Ss���iW�E}��O2<�F���k��a���Ҩjj�MQ�.	��L:����m���򀊀��1����ȃt�h�a{�э�=�'��5�y�o}�Ӣ}��f���9X�����oTUi�V�e�����FY��V_t9\%���p�HM8��O��Ʒ��>P�s�QJ���oj�e��G�N�����Eg@�����L1�e�B�	�Q�X�GBc��y�0�Ԛ����M�/������_m��6]�w��U��g�R��������e _�? )��FJ�^0¥Bg�W~����2����ī��tG���WL������j����0�뉩��ܶ��;jJ���5��:�_fO�Gf\�5��No�U �j��JΏ-O4�k�ٔ���X����&زK��)�==8N�[�ub�]V�4\�dmj�%��1��m�"�"3@�b����wJ��2ڏ���ޮ.I��Za�4eCr퓌�����Pܡ���Q�z���2 �_�Z��-Gsn�.��E8ٔ~�1ܦ�MpK/�r�\w�)�'PY돞��a�f�jw>�/��T���,}�L׸���(a<)���L���9�,<*{���������p2�D��]���f� T�pU=[��
�~V8i]_v(��{�+��;JNlԋz�� �+��C
�����F�.T�U"�|��b�zm��GX8^έe(Y���F���ı��:�b�:sp�IF>�r�+��AN��ܢ��0�EL=��N��q:�ϰ7�j0���֨J���S�1΋(Y��TNLÛɶ�7��>��n�]G@<���^�&�������E�ϥ������H���9I$i��ȕ�=��vq�$L؜��_l��
��N�b�g��DJ���Ԁo6���s�sZ�b�8�&9k6O�Uᒩ7[r�X��#_|��}��ޚ%�)b��A�ր��9w]0����|Z���TdK�\�G�9�y,�k����;��V�`�[y@Ө'�(�MsC���Hk�,o_�	��Mx�]]��:�J4tM�N��ۚ�r�ԛ;~J�s{Ƿ��A���}t��Ss{���:��d��˦b��'8��3W*����ʟ�.�"��=��Դx������KU�9�YJ�x+�v<1��V#��X���b2��~GeW��@�u~�x�K�i�Ku�~�󪖬:�)��o�L�#z�\�*�6�x��JW�Y4 zkJ����,]��0W:��h�]�V,�K�rb<�`������$���O&z�©@�U�Q���Qγ�]}��n����0���FD�� Ƌ�x�o@۝�#����t��2��[���Z�.�k�������yC�E�}{�GW�~��a͝,\*C�۰z�f��D���K�VBUC�z�?\gKg�����LIv]�G�s��7Z�[�|~�2���|�|�x�p���Z�tuj^*��=�Ê�(�P$Ԯ0�ܱ֪� �S7B�ܩ�[O� �ҕl�)C��X����
z_�n�Ww<�����dl�1��	�e��<]Ù��X�m�R<\_NUUWl+w��Bn��ª9�0�w�_Wܝ$s�rj6�Nt��/*$+$$l��tƞ;&���]�ѱH�Ô_C����[e���]�v
���&���h�j��i�4�˔�pUJ�PM�U���	`���m�\a}إ�LO-Z�ܹ�(#��Z�9���-� .V2t4oyM�ň�֛��}r����I�V�봤�HO\�#ݢ���;�#�P��m��Z=�������d�5�P����n�2��X�˷e�����ɎZ�j�N��������U��R�C G�ƈL�.�"]+sM�=-��]R�����f�Fn_{��5���^GL�K&6)mD��1K���CD1j�9�e�kd��S��j��<����0�����fe��[yZO�NrN!���7��1�[��9Wl��+�b焋�Z�1B�MP�����@��0�*e��3a��ɅћNI���i��)	����&y�u����=��_ C8�T7U���e7	��K
��t�;����@{q5k��;�޳��`ƞ��i�;��B�di���O�U�-z W�[t/����'7�hЃ|��\�֊�l(n����d�q�����u|��e�U	u��z�J���r���Q�$��z@�뉄.��C1�P�R-�om�,�zc�ΘX1a�9]��Js&O�����(�p�����ʤ��g��_�� +������P����~�'��'���,iTi��"V���Kie<eVX��-w}b%��2��]��y�������}�1R�7B4���I�	e�գ9ܱ�)�P�>̗h�ǿ N�D���7|0���]L��s� v �=�2�PA�O9�b���V�ys���;�Y�kU7>��b��E=�\;!u
Sq&,#�_A��P��ۧS=]YY�:|�m�R�W�����9L�e:c�w����Ek�c��v-fg�7z$3h�xWL���PMD8۝G�Ć�}�j�T�����М�	M���W�@R/|���r�Rɷ�ը`=�|����:�Gq�g���8=+��#�鱂0Kj���v��p�]t��r`]Tla������fGT�3�s���p�1���������/��C��ûy|��`$��:kE%*L+�`���í.F���x��W��S^#Û�)��[v��		���HQ� ��UU���-���SB��^a����.j潿lG�o�ε��w���o^SB ���5��*&a�3�nHh�w���}6����2\i�=�>�b��yܞV|�� FGl�1�wN�k"n��AZ"��
	�5�A��@���qr��d�&M}�ʅ|��fCj*t�5U���I�{ MF �w�����:�	�\�ڎG��{���X���Sw�������W���ˤ���KV|�u�u#Hu�U�t9ގ,d�`l��^��
�
4�.�_�7Z
+I��3*�m� �]ӵe�F�ToU[AX�8+��9FfQ6��{Fp�P�:?H��F3�W8�gA���@Toc�a�O��ɞ�o�7a�iRA��2��}9�*������k�H�t��u|�(�\:2o�}�>�|��	�f�֭�Dkۯ�7bl>�;�D�v�k��;b-�Y� �M���r�g&�\�h���:�z���������]��:w)+uFxu�>"_t>�G_W%q�wrn��GIh���c+S�K�f9�0�nP�o���%ذt�<}�c\v��19����q�:~��,r7�h+�%���mPeq؎sP�1u	��e�������{폪f�C꥘�(�I����E�P�x>�_*�2����;�2���c�.����	zf�T\���j����?Ck�ۀ3\ �=[��������|��gαT����hN\2�op>����,���A���O͛�\��T�)o i
��imt�w����f.��S���LH��v��'�{$`��L����WX�x��UoZ=L��E�z���F��Q�qC��-`��n�j�5�u�Heu�T�R=��4���YO)![���K|4��j�gv[�sBLŘ�����lΆe��L�0���*S�HX59��cZq^^Y���:JJ��<!�D�-o]c�au������mw�O_���w�Tߥ�l�p�f5�}ZdCv��wDRsA��P��AG
ͬ%d�[�Q�80|�M�2Ͳ�%�2G�b��
�n\�	iy@u�ydT<���)�u��T-B�n���@&{�=�r!P�~_����+�aTg+x�6	��R�>{l���YM��9�4�{C����&Sj�\M׮[��/E�<�|-�mY(_�Hs we��C7�V��[�1:��~�p�TG(�\����}�r�-��zkT�3_L œ0(�ؾԺ9�U�7��nPRz��`.�F���!��c��/��KV%��eЅ�8�{�v�u/� M�E�a�����,]��,w8��(���䡚���K3Ϳn��WP�U=\�X,U.�W�ڬ
��3���W��t�[ʍ\��/J.�v9w���L}9r~l��_�����"�T}��k̯Z-������Y��P�u�NI>O��㾞-i�J��V��]�>^�`��n�SE8���26�u6~���hꈄ�{���-v���zK�Em[�}s���Wr������"(����Yʉ�Yָ6wY��({m�p��-�sl��ӳo�96$�L��+8�§w3���1{+�V��lP�����'E�S{�mKv��b�T�L��wc���\��
��^F�7/���V�/�������uւ��CΎ����ec�ٽ�WxԼ�_<��:��?	x�H'���Z�Ϻ9�:N0YD]�b���:��}֖T@��=v���G�h�l�^�Y5Y�c\T��'3V���S��f�cyۄoKYv7��]�����e���� ��;�g���e��9kAu��[Jr�ev��.K3��C��gï�v������Et�)�-<�:�Os!�=@ 4T="�K����zރah����n&���e��7�Qc���Xo�a��V	�s�;��3�j܊��� �t����tG/i��]W�1v���K\�սB��d��x�U���tV���wjtm�T~�#�)�0�i��]���t���*��E��#m!��NϊX�=e_!�-�a���Y2ʱ�;Y���+���	�c8ՙ��Ci�c��D=9V�xA�d<��&Ky&WHJ�"�k�A|�ŋ�S=�1\��%��.)$�pr�l*CY{!�PY6���$Ś+�a=:��*��*队LE'b�t�,)ϐ|j�i�P��k��/r�>���ɦ�U�hr�Q=3rC0#�����VK�g����=�7��C�bHvq�� ؒE5�*����2�ࣦ�KZ�7����
� �]!|w]+����u��lW֎»�E�J�Dj�/.f�+�5Z虍]j˺C#�F���$̣�#��G۽���h�fdڇn�mwR�wu��a�X�F���g�Q_|������]x��l	�un�h=r���&m�
H�c)�� fэ�v�岜L�]�%i���l!��7:]j8˄�~YOo6�����7Lޚ77(�R���ڴm=�Y��n�����ݮ!��=s��4퓱pB}%+�h�#zE� խ��n[o�Ji�Q5L�V(���*�+�ܛ���m1�y �YY�sw�b8o7y�JmX4Af_<��Mo#��Q��6wRmWlÑc��0=Y�Rf4��9`Q���Am�f%�Pol�^ǿw`[#�;ڵ���逨 9cd�p�sEY�K��Φ�s&Ր��d�31��R�Rt�9��6+�#��7��t,Hw@5�b*W�o��y�]�Le�'l1Z�;��n����a+��O�X
���z��|xl5n��m-{a��fw[�j�U]gU�%h9d#�77�қ��)�#A�9P�� [k\y���w�Z���AV����Z�2,D�D��\�k�tɻ��1��ʀ��7W�I#�u��voN��к�q�n��C.���]��j����	�����=ɋ���Gq���s��F�'�ʛ�a�MV�WAM�[����y�����������[׻о�DP�b��Ĩ�F[lV��V+QU�"����bA�6UU��TX1m��[֢�R�,H�(�kD���J�����ԣ��1Um--*���%aJ�Z�lY�QEU����"���2�#Q������m���PA�*R��b�TAA��F��5�k�G(����
6�1,X*8�ѱDDZ��iX�(�eb6�b5�UZ�iXV��cm�U��R�)RS�e�DcZ5
�������DkEF1����[r���m��DEJTlX�
�хB�(UF.Zh���QD�J�Zд��Q�ъ�1kAAm�T�j"�P���2�
�hV%j�ۙ�KJ�Z����Z�+P����Uj �"#6�K�1F�AEkK�o�Y�y�=��5�cȇb��w�Q����0�U&ŝ��u�Gb�=���,�Ⱦ<���,�ӵ(!�lnu�L{�_�U}UU�}�=��ՠG��A<Us�"�����p��,�Ձ1S�����̡�>�XP/3�>����Fg�WU��[��2(��Uބ P�nD��1�'�)H�"��M�ޣ@�I*b�v��϶��ok�J��x�X��}hp�YP���U�H	MAs�#~��}��S��g(�� ��g�6��__m|9:H�nH�f��V	�_���t����0?kY��V+>o���Z��;����JF,C��K�W�P����1�zM����SLf��[I���3(x��۱]~�P�咈�S`�����Ѓ�]rÞ�0���w�u��HP6�5}�}ɷX�^���8������_Z��K���|��rC*:a�`P/�8\67n$�m���E��>��1`uCw�Oԩ��r)�i�Q�d�xOʟ����'��Dw�^�c��h����1B�} 7p�ݍ����4Q���3a��Ʉ�_L9X	�v�h��*��ب�B�����ʥ1�k���C>J�Y� ��7TÅrh�߽e�����W��o���݊�w;��1I�V:^���?n`��,�(҈R:b������b֓z��e�f��4jT�+��v���0��r����յ�tm�qL�-Yݦ�mjx��;��n�y�.��� <�\�zE��ʌ�G�}�mM��|��0Bۛg''�y�'DE�S�j�kYC,5�uW���Ӽv�9q5�bV�}ݨ{Z8�M1R�	�oEޯ�b����3�Ui�N���_����ydBЫ�Ģ䐓�o�³"��p�}܀�'�7)W�vxO�ʘ_ /�9o��u��g_n���+zw���5q�\;>o������%��1b9�]��U�~@W5����y�̪~��}�!�z{j[U��l�=������(�A�bS�*�d�y���)�^��00��۟oϳ�n��vE:cE�z�����Y J
P�^)T��[Ǣ���]�Ҧ|��"~��s��Ą�F��W�KN���<��Ӧ7��R�3�{0��nVǝ �*�]K�\�h��81���ikUw�"�ۤ7 U�f���@�7��S^8�	���ώ�*�#b[��p��.�P꽯�|P|x�vVӏ�֫�������H���F"��&��8,؊�F(�͒��\�����#��<����x�2�Aw�7[.�Z��r=�Uvwț]X:��B̾�I/�Q�w���xM�s�4l�y�o�kUb�je���9�@q��Imū�>�nզk��Q:EX�B}��z��.6��ccM�@ty ��%Z�.󒲶�ﾈ�#��}e9NZ�F�ݞ��x��m\�@�S̖�I�E.����VM»��Nk�uUTH�qcLG4)������/)�#� nW�p��耟%\7%��̋�^���OG��/�gB���R
��y�����mu�)�@�T���Uݎ��d�&�aN�5�.Z��*Rꩋ�w�_f��4��8��5U��P��L�us��J��s���̓��:Gt�Q��%�<��k:�R{��1�΅D���LT��;��{�;=R=7���b���ۃ�2��ʄ*,�(\@�8q �@dhGi���3cq]k�|�Y����Ν��>A������7K�Y�K�Ab���!�k����JU�wZחws}5݈������;Mֈ}S�����+��7�u�ONE2�]�p��`��IF^����a���!���s�N@�n_��.6�)�Q�kv�C��v�K��<���x�`�L�۸w�L�����7�h vv�Όw1���i���K���h��*`W�\X�Kx㛋w�/�2�[�_n��ť�SP:�_>�Ϙ&硁��e:�w�Γ�18XG���YqΆVkbM��ȰV9w��wW�3��q�:ȡt��hu���^�-��UfA�U���ؿc���F��?�W�}��=���&:���~[@S%\�a&���E�<%ZZ=)�O�P=��4��r.�9�&ř�o�-Ir0�(�^�FB1��S�9�{�b�|�o�<<)x��x=�%�Q���"��n���n`�n�C{
��|���@{�R,��a�329��ƨ�y�M���p��$\/�<$Xu^z���W]t�HU_juOS
�J��@ٽmg��[�6]�s`��|�V�B��P��A�n��n�RG9,����E��p�|���1�9�C����|
�s�V����J���32o��W��\����X&un� y�ߴ��{����P㒔|)�9���F)zwC*P0��T��as��V�\ν�P�'�!'z�t�E�ڭ)7]r�X�|1���k��L�w	6�󌚁���iF83"��v��%���!Ww�>�h��JQ����t�U�.���&�G��R�z���]�L`q�6NfY�8��n�0	�5Ğ${.��ry�Ơ��u�H_��m��^�KM4)�.WŎ���%za������nִ&�["7B�$��{�3�-�lf�Is��}��]�;��Fv�����|�b�6�Cn��X��}�����h0�YrD\�K���,Q`V�QOU.�U�U}UV�~~��OC�q�vn � @�X����C�bx�kv�6p`�rt�}��%�oNX\��Q=B�e�U�;!5N�^K�����@ʎ�`TE�1�)����R��1�TdcՖ��Uۡu��)"3�z�����ZY�Y�Y����奈R��9f3��6�{��v����}��;��-���f�ٖ5��*�q��|Vt��]M�����=�Mj�Y
2��<�)�]1���������R�����iW�K���y�x��we�W:F�8�q�(`�}��C/J��@��17B��J����@2��19W75{PA��^g��YS��mK4���wZ/�u���WS_(~/m�ԝȊ����:3�q��5r���ڄ�G��_W'Id�S|kE�R�.U��C��w���6���@�������Ș.W��!��Ƿ8�!����4B�NMtwbߋ��]��WpT{���\���-&��0YS�b� �9u�y�[���d�P���[�*Tn��S�+���r�;,P��Z����E��Ը���]g3N���x�)�B�@��h�kF1��
)�x���3ÓG�A�oB�,!��wj,��d	����b��U�<eQS�[�,��Q�2�Z���yY��uD�{?U}�}UU��I����l�~��UΧ����� J�aw��/�5�iU>�H:�^�xG7[w�e���qަ�!3�jJ��&,��蘥L��USӶ����[�~_?+G���]Z��(醦�����`�N�1�H�� �
��A6 ��b�X��3a����/;ݜ�+��q�Md��)]������C�S<��,,8W&�G�D��1��k����r����^Vy;[7���������<]5̀��a���jU~�S>�� ˸w_W���<}W�V���+~-xW8�;7�c�‟�]�TGwS�((9{��.ۙq�O6?�����J�
G�Y���![���2��{*�p��<'�!�_ /�4=�bd�)Yo�=Í$��[��/�����3.*�g8Q�J�0<(�GX��P�xBoƚg���%����0+���r;zs\�q��.���N���"+�+�F׏�M�Ey�c��J/{���ī|��̗8*������m9L�dS�4_ʳ�F|�Ԉ뇴/� TtR�1v�{����r���-c�:.k|�����8���9m�V�X�ݐSw�4�*�ݾ!v��k�s�]b��ix��e�ꃝtܬX����L�_\�V�$��ŝ�/gP:�P��N��]�8Ys�c;9�����6�m�G7�rֳ����M�����}�PY�w96��`L_���Q�r�Ą�jڅq���0�qa��Sv�X&9����,e4�(��RU�)ƥ`E�*@YuR4�@d\�h�;�=��=T�v���+mS2��G<���
�C��x^*]�Q�[�$ ��vW��Y�6�߻�l�S`���1ti��\̹F�U���[.w�=<:̣?B�N�v@�٨0t%uJ�Q:�@t�`�NB���l�1�vG�j׳i�.%�1�vt��@W�2�b'���r&@zk��1�+C�����)횵�+&8f^��#�,l'�l��e1�G 	��2��*f�P�L_�ԅ�ٖ�`�w<uR���ݔB��['C���'z@�_rw6m�@4r^P) i��g���n�<X��q�ǂ�S%Է�:��S�\0��?����
1�ڊ�TZ�8A���߆OV�NZ���-�YD�����q_�9,u��(�~�^
�E�w�*��{P�=Li������Τ����b��6���C~��Ɇ���L!A�C�`�8�~�"�躻F>�Ӹ2wJ����']�؇)�b�&r��a�5x�T-С���_l�L裖���_����8���;�`\�N��WmX�x��Lt��jf!�+i�=�mǗ����ɛ���Ob���4�م�U�g�K�N����f㲪EYYM����O\��Wz�������,�[{sw�{ゴ�N��`l9��>A��Xv%{�=�u��r|�����]LN�ʵs�������ZoQa 1W�H���m���D&��P�zkꄰV��u�OHY��u
��6�/l�B}N��1�k�����2�S�M��k����Ԁ�xu��9� �Ɛ�{=76R�������
Ȫ�/z�lFL�����ީ���^��L�:�c���eZ��b�gy���5��z���v0��
$�'�f���ڴ�zg?��\�[�0�wj63��='!E�n/i���/��\+'�O������/�a &"�y�[(E�.�vi�X��w�7�<$8��\8/�_�`a�j����������@{�R,��ň6�\J�{��C��3/\F�5_]F�*S��ġ��"��)�P�9�X6J1B#�M�L�n���s���H2���[;����N^���a����V|�"b)�P����ޤ��ԬWP唣�E�������V:ج�$2Glő�=�����uz��#\�Q���x�P*i�.}�g�7���fͭb���8z�u)]�M�ԙ��Eg�R�>ޒ�2�|��H����&7���B�SWy["�)ʻ�U�Z_M��G����;]���X�})Iw�JٮWR�S�#��>����E�`� z/�
`�.>��"�"�?v)zw>�P�=@­�o.`h�1TH��X�8���s֮�Y�q��t����^g���ht��쨼1�c�+�ۋ]/~���j�q��ZM�6GLT&�3LXw� �����>G�siG�����KU�?-ѳ�m��&�m�[��.A�����=μ����<!���dG�>CM��]f���В�5���^�r�3���Q������� X�XĪ���P�<d�l�c9ĝ0�� ۮr��2�ô#h�x��[��ֹ��U<r����`h�q�9��&!��ȶ:I�p��V�;O��/J��]+��6E���g�gh�Ɩc�S�hS������'=�	�"r�r���&5��;��e7�H��v�7�o�T�Q+�-/i�$^����N�����Fl��Ƣ�:zT�Te�k���#`��"�j�	��e&y��2���oV
ksg���=�;W����c>��C�cn]�TpL#܉S��!m�?T	�n�ۅ!��/d��-/��X��&��)���\q�@,Nz�gA�oy�����ӽ�=��̙ךui�[�xF�΍���?�]�>�z�e^�9Z�����wd���n�.K��L���mb� �����<��ɫ��U�x7�U�U}U^�5���.
���+��U�
׵
����^�ϚVG�0�}d��!̀��Ih=w����q�w&��Ǒ�j岷f*/����N�9��5z'[�|
�ܮ��S43z�;X��W]�T��Fx�G|r4����j|+���V����8����u�,9z��(>�ieȝx	EkrȦ���cLB`�Е�U��0Ō*{\@��և1�4����=��	��M�1
����Y4�P=�5R��^&�S�t��^�s皊�YX�X|�85�O�S��)b��h��T}�����-W^U[�~w-\�ǵuX��4����莚��*7�S����|UP�r	��Ӣ�I,v[/����9�����mxr.�C��rkL`��;�t����������.�eTL�9�|+Gb���������9c�j"�;���Ї��i�;��.��@i��Ypn�-���:)���;�ھˈ����&�1�4[V�\��]����+O��V��5I�݃Ae@q��:�A�V�$c`�tY�Ĵ�wT��Z�4֛o�w���_]C�\s%^F��ˬ��9W,)km�f(�.�W�'X�����2ŽUu�r�[���S+T�
�`�,h�7�-����kR�rJ;��u�� ĭ�q�e_v��N��*��L���|��l����J.� ���R`+�8�S�̂0����4t�𡰄��˛Nm�MnQwK6��t9�����6�G�Eݴ(<	�}V�V������Z:k]�i^����V�wÎP��E '�V��P�G����]�o����Y;��<�U��.�K�8\��&t�f����h������>Q#�v��N��N�ݖ7id�65�N7t�;)kږ�gbѵ!ٴ4r���Oy(�ykr�h�ȭ1�ÌZ��:����1H�P�>J��4�kW}���Kz��^���!YwI/���#r)���Op/�3����6�Ҳ�V�7�nx	BWSA�I�zԶmd7r(R���)`�*4Qy��7MV���9V�]��F�^��|���m�)O�M�Ô!�޽xȆW����>�Ơi�U��2���+t�."n�Ӻ�\x�Z��r��
��F�B��ˮ�#�����[�9�1n7��ݴ��n�J��	��b����*s�����B�7�6�:���+k�v�a;D7ө>� ��Vu�ځ�
]�b�;�ޛɦb���`4��4u��s�?��Sx_-�6� �u�قʥ��ߞuY��pW_c��.*�gb:*��* ��ܫU��;������2^�%r����gRx\{����,3BaN�'���t��l�dǄ-���*Ĳʈ_7I�iuМ�n�v����z��{�ۥ��M�w���%Et������B!��Mo�hW.�EK��YO��׃-����4Ozz�mFJ^N�OÙ0��t[438Z��`+�l]�j�����ui�ɠ��k.���;�p�ͻ�r;Me��C��yI�,��7�����ǝ�B��:fT��9��jۣaq]H�r��T����7���],�U�Q�i��wB�1U�F M[�!���y�<zƑR>�\[7��n��;��MlSV�����b��������[�]W����=Z]eKIe��Q�9K2Q'�x^n��S)�Dk!X���E�8l�К�Tzc����W���e�i'6.)�ː�g��r��v���9�H���jSe�/p�q�X��fmtO+ruw��Ω�Di.��}L�܉��hN��9N��KGT�\0��uq��`Q)Þ@�F� ����a�ٸbK*��jh���
 �S!�׭���=O4V<����ל�R���I�������6�^Ssw;M<(oL�بt��uD$n�vmYY��?~Ȩ��Kb�1�.R�3�ĭV#R�*ڱJVU-Ys.�ƴA�����$U�!P�X��(���X�ke�X�EVRʌF,�eQKBŌ�V��(���PQb��PZ2R�Xʔ���cZ�5PQ��X�U��kJ��F#EQF#X��,̙��jQYR�b*���,F1DE"�Ŵ̰���(�QQQ�h�F0f%EUKq�E��A��F6��!�+mVTm����Qb���((���E*��ъ��ڨ&P�#�P��TUUQV(*"$ADb���H�ĭRA���ff`�TF�QQ
��"�Q���1�*1�*��R��UA�����%F(��(5��"**#1b*V�dU *F1�R���R�T$��b��b���6�-
��Akb(-J4UF1�Pe���Qe[R*ZX��Bڭ	�F�.�o�n��C]����!m�n5��<�ꓨ>m�ZfwuL�]��]�+������������+���}�DG�R��9U.�.o�P?�*�m�Ցya���b\��0�ٜ([1#qH�P�y8���M��ۊ֜����ϭ�*.��ܡ�m���(��3Zn>�1�:�aY�E9N�_fR���J���!=�eƧoND9�mV�]��+u�e�ҷxo��jQfwY�t��R߫ݱ�O���%�����O"��C�L�dT��ᰖ�+n?��vxe���E��9�ߨ������&{yu�C�_���V�KN���=	���t;w��LbZ�=�<U��r��׮�����D���Mk�x�b)���Z��{��󵷼���fʳsJ6����t,�<9�`\��v���b^䁪�t�X���37[y�[ѳ�:E2�w�05P#�&���d�e+��X��'��/ZyUoJ�Z�'zBy�գ�&+���ҿB���߼��}���I��"W\�0��p�3�\u|��Ҧc{`�quơO�w^��-�]������˶RV��'pAJs�6��񣚩\�MW�\�U�%��}ZK4�%�QA��T�a���������A��Pj��p�ʗ�;b$e`݁;�1� ���c�)�]SO@�)}�ts�XWu�����i�t�+�S�&���b�v-��At_�ﾏ�蛞�ߴ�N���ht�Wa�x��
����
�&i�7�^D�-�ɾZ_:o�k��*��]���9�����
��/�X�ڏ�@,l���Q>���w��5W�w��p�џ���)v�^z��eR�X˧��^��S�gvT
W��訴����=;}cN�T[Aq>}>+v�"�����o����kN�^��J*;�8|���s&�oTW�[w�Ҩ.&�]\Ǡ{�	6s2��$�c����#\d�(��X�e��n��)o+���N1 _e���#\zFr;�ǳs�QqV(�_iyQ��O�ϝ��v���֫L�Tn\��hW\1�f��qPkZ�8�>]��ַ��ky��%2�Q��iӎS�U}��kY�T�W$nj�D�>UW;�V��9�Nn�R��������?�M��Af�a�@�g6�guel��'#�m�	V=��5}t�\�H}�hź��#��T�R���P����"�,�N��2s� �H
w��0>�]1�
�O0�f��uܣa�M��@u#����8!��`͍)�va$��$�{�/{��,��y|$<ݤ�s�y��]���I�o�R���DD}�C���Zksl���*�\��u��ѓ�sg�T�a��t<��:`MnG^��i��pk$8�]���uT����V�dӤj�*�5`l�*�{ڽ[���X��gֻ���D���[���n�Y�c�Un��:�^M��=/vds��(v����s�O�d�Z�>��2�+���;�/�ä�d
[�6�50K"�ʜ�X~�BR�r7�reAo�M,�2Wd�'�a\��q�s45N�K��Ě�cT-��<�b`�<s�����(��1r�z:�����P穥Փ}C2�7h�޸{AW�ۯ�p�ʛv�3�p�њ�Q�S��V�t�z�ڼD)��g9r�y����v���aX�p:���;8����5��ɜ6�,�P)Nc~}CT>��j�>����+P([��|���C��8R�l�<��)�{��^�Բ�.���^v������3�b����A+I����Svf	�`tם:��ҙ؉؀+y���r�&f������cI��]�V���2�� ���ٞ�݃��
{-w;��U��g�{��Z<��1�o��Fv�)Z}�D}�����m��+3�ɡ�����=EC�g����^�Ի~e�F�7�=�mVJHSf�%m����Ya �ƗU��,�/� ܂E�/llu]T�M)��n�z�b��G!���Y���m
���7zUfj������k�:br4���
���[�J'���2���[/X릕.���>W+��z��+��Cݸz���w���a��L����J�R��s��F/��/O{��6G���7�I�|�Ihr,\�U:�s�Ҫ+&\ݗ��9�`���_OK�>��hs���{;��Tl�u�˘���p�__�J�S��]�-�c9�WBk����h0��;Î�<��u���T�P�)��٤Y�ru�Y?S%nL���j�A��2����목�����>����W�FR�x�6,���C�r���qX��
ٹf��$R��Ǹ���jH�T���9�����E|�К��6�S\����T�p�Ğ���]v�x5��l��'F���^\�\$�*�Go+������e�J��;��(�4h�c��B$���پ�;�]��Q�Z��51#�Z�r�>������o�^���½��c7:k�y?oPU��j���CYg%l&�OJg�n�(2O0sR�;Cm85�Qy�Qx��,ުK��]C�i��`v�Gt�T����ɊA?�lo��rލ�U۫7ؼj����]8�k<�C��)�{jQ�ZV�ʦ�n��cr��ʃ����'1E��QN�]�_Z�cGn{��)��6mz8�Z��6��^j����j���~�9Go��|�٤��O�����#��;��TWܱ��7���ۍxy=����+��˙Ρ�X�p�J�,.	�q��D_G*Ҳ���=OqSݪ���ע�s��~�w��h�^,K�]ⵀ��sPb)�Qg��ϣT��)�j�X��`�ee�9uj�Ms���a�삙J��N�\S�%:�Z�4��P�8Oe��V����@)��+����P��P����Q5���.����s�N/%5vUm���c�.�m�oj�`�����	�����Cz�K��������A�ӅMy��VR:D�w}�f�{\G��\�uF��rV��#�T�ɗ��)S M��R�K�܈�{3v]�ٷyo�t U�;���b��,ݓ!���c��]�Q��������U}��=�7(���5�ݶ��-�k�Q��Ж��'�5}<q�V^��7B����̚p�OS}��oFLE:Fep��Օ=9�R�_,j�WX�w�t끛�a)��TV��wCy
��r�+�k����Z��U��nr+��bqe�Y���5ݡBX��^!�d5�P�)1WJU�UvcD[}�]E.0��'��TZ~�ËhW1�ATrf�����UeU�oc*Ukn]%7E8�u	J��+pR=E.>a��X�]�ᾊ������ΰ���P����a=
���[/�C�җi^o��k��nt�U�aT��p���6C��q��]b�@�p\vTWQoUt��1�Y�T�K�Jx��1��[3��<�J�gH{��K9^�m�v�!�t���ib�g�[g+ �)�t�Q}Վ-�k��Q���7�P�����9���.��:!1B��CI̋ w���c��x+VSN��L��$�8�}�����B�uέ�z������{׻�`ۧ�Q��gWlt�� :�*���xmur�tqE�lP��7�8�b7�a]�au��`s���b�HCo(��S 0I���۬��">����Nv��8��۰��1s��=�Qʾ͊�o���Z�;땘i�|�)�a M*����0%E,f.+Z�����W�T}����ݔ�����i^JZ�m�9����{��H���o�?���}\D�������5���r��Ǻ�Ʌuz�Gf�a݇*�Q��O�{zϖ��>�j�׫;�ſq]׊��=?7M��)`���<rk�wA�����P�=�j���ON���[��}��7�|7r��3�N��ջ[��l�V�F>��!lB�<l%�pe�bs[���ným�-Ϛ�q�Gs&Z�A!0P��bR	}��'��V���,j���0�_}*zS�_�]2�v;yn�)v�<�p��|�11�u�ie}<Իm:��fA�n�Q�(��x�������k��V���W��yӞ�/nB��T���6v��_3����{^6D��o)0*)]�M_\h0�7��Qf�׵~k���A�Q-Z��[Ϲd���J|ځ\��_g��b,*�=�B��uy����w�\3��i�r��Mt��	�ܾۨ"d�M����/�<mt�yƦ�ѻ�I�H��N ��p�)8. ��/�Oi�W���	����Ȯֳv�ՠ�F71���ˤ����v���
�끵����ys&21���������.�+���ڧ�*�o�g^��}���;^Лwvr_B5�w�Q�죊�.s�-�j�^�Բ.����ek{fe���1�)d�}"�j�{��G��k8���׏Q�n��N��=�%�֞�*��\�x��ȭ����.mW%}�y+�<L�UD.�����qu�#.��f����<s�B=��ko.�ێ��)�ɶ㺡lJ�������uαx��r��hY<靯G�>�V�J�_���d;z�ҝ��V�7�QR��[WV��ø���6�N����%uF��_]���O;iͧP�+d7[������(m�1ξ��-��S.i������4�k��]g+�&�;k/1�L������E�$G���mn k�i�}J]�/VL��F�
פ�$�`�������7�c)���F����#Z�u]a�[�٥�Su@X��hS�&u�{���.eN�q�p�9�5m����E(���ﾯ���*��.�2�G]b���*�`J�rʉ=&z}<J�E�ŧ!��>��w=z�Ns�M���v&!\��a��*x��.��nciA�o\�z��%$
ݵ��P���o!W��D�f',�����o9�b�5]=e�k&\b��U�o �&�o�\����L��e�ں5}���fN$�����:��i����ǎj5d�oPU���=�a\Q���B��*�L-�eԮ��S�D�ȼ�W��,b�=���k�O-���SԭP�������[s5��W���.���f�ט����^�toS}�7*,�}-�F�8o��>���q�ʚ��_k���P��t|�j�ū�{	���֫�4�(r�ӞaU�/�WO?K��*��@Y��S��"�"��9���3�ʍ�����Y��9ؓ$�=�1Ⱦ�U<]�6���?!7�J��J��<� ��:|�3��>���Fc��{�|�{���d�E#
�U�V���d��R��s1�3kr:�B ����݇��wR.nY!Ds��B�.w��˲�Ԛ�ijL�u�cj�W���c nڭ	1��jAuA#����|�9tD�����g�ﾏ��ܖ�u� /GueE��QʣJ��Symp}��zYP�i�g�j�	�yV��{�R�M��_�S���w�>x�/���	��-�m)
E_hu7��r��>tL�*R�u-�TWBۉ�?N�M>K
}�h]vk�Ď5P�U�i�L�%K��Y��i�v,��;0R����s4&.�������_G'{ӓ��-qٝF7-��*�%_���\�ԣ@W���sS��g��Qt��e�Sk���&)�(�t�|�jSo�4`��\�[VpZc���Y����PV�p�����_[�0�T
M��w�#�c�"i81�H_�+s!����c��K���)3EtuT.y�۹p������`�6�D�T.�.��u�m[�U�f����Ԯ^�N/�qzy�O*�ǮQ<��M�}�me}y��ޙŀ�o���i-+�Y��l}������G��Y�yVm������Ė�[4�����>�ut����If�<�[��/Pt�;����
>e�K�$�ũ�wPՅ��s&%ٚo���q��W*���<y�����Ej��ZY4ղ�P��F�vd�/�q�Fq�
ك��zû�ZÛ�ߊyi�=AXQ\�5
�Y9�%�r��	_bh�gJ��v=0�^��<mc�����.^��D��u]��WY�O�-Pr��kI@kvR�|����fB-H��M]8��	�f�\}Y���v�_:A�� ^e��79�����LAK��)I��1��٣���uD�M�ۏ:'��E��zp�ST�g���!m�h�����
���8��LX㗔�q��}d:�b՘N�����=6��ܤ�Y�υ;��hur'v\I{h촺�"�3#�p����c��q��Vu��u���c�`E���5E���0���9z@�#�d�Vв��o G��r++m\��6�Ļ�J����ӑ�̘���<ࡳ�q�(Y�q�J뤪�ħ؋��w�%��ww��E�l�`�Xz�@�zD����r�w}cJ\��w9��.�\��Ƥ:�ù��' ��I�(s�;��r�p ���I���5�s%ǳ�����WR-D$�]|�.uv1�=��8�sc<k�<Is���\J���u&3.]�����PY\j�jD��,5��ֳ7��@.��M�oәC�9c��Çe�*u��a4c)�V���L�F{G��y·t��)���5�S{j:5daPV��ڌPehv9kmov]{ɎΦ��|�Э;�\�֋�C�W3gTJ	��������RM�@d8>�\ ��I���#Z�1ɑ�z�jJJV~w;#�DC��� �w!����vnB�s�*nE���w`L��ƃ�;!k;���J����	����Ԉ'���)�@2���w;wV;�m/���뢶����vb��*��!�x����iPD�-����?ؠ�N�r`��E����CB'�㾶�f.rd%q�]aQt�W:2��:���G�,�Wv��k>]SYdлb���/��R��ǩt7��#�4:��#��w;db�z��"��A��2��գeb�@c�Y�-.�tÐŜ�+o���W
��ZzS���iy]F_]7W[3�b��G�Vq��Ƭ
j� �Ew�!�7���n�����,T�uu���(��Q�[����!&��p8Eu�Υ\�5vhJk1��ݟ~Q�u�x��T�-/}f��o��U�Z��I��Й"/w�E"�)�vj�[ŉ��� ����L�og-(��70�n�˼�{��Ⱦ�p�17x�K�AgfV�X�;�9�'��5��=��u)����Џ�hlu�մ.k��4�x�펖�N�6��0��z������ި�P:�����ó/0�1�ND�e]��i���eJF�XpK�lnD')N��ov�V!���W�X��
 �X��*�m*�Պ!���R#Z�KRֱAe�F�,�Z��)\� (����T���[b�ĶQ+m�B�DX�YRTETDb�1QHڢ�\l�ɑ��,[j�EEX�b$PZ�E�V#X�*0E@X*(�E&6�R���ʐ����ik��F0GUEF+c�����1�IEFҪ��1*�R&3�-�R҂��V+�(�ʵ*(�,UA�Q�s
�QƊĬ���EЪ(6�P""���KD���XV��T�+m`"�eTEb��2�
�U
�k*�(�UEB��E��P\���PX���EAX�l+cB��mm���PP1+"Ȫ*$UZ¤E�ʪ"���.R�īQc#-��m��2�qV
���Q(��Fe�m�D��UD+b"�V
�-mX"*"�-|w�|���R���������
�`��@*spLr�'.������7q[��uh�Z"m�L�/!|��^ *�䰬��>������ɾ$^���l���=Q=q㯠.u��r�!��K���e�fE�33��y����̃�Z�q����ʚ��ek��P\vQ�|/X�{S+i�5�
��5�2��X��9���
ٽRx��zp�^|����ܭ��L���֧��C�V�|=�N.=1�����z��}Y�}0��tߧ��M�ӻ^���\�y���7�J�ι��Uq�]��F��<Ov�aL�\\�_%\Ry�$u��}!��W9�C�\}5+Z�����ڥon���d�#��.�#3b\������ܤ�!Mo\'���ؕ_i�j�D����Z�FMȞ�iq�r�qm�F����{���k��L-L9��m�A�Q�*�h��9�ed>�joM<TzWrA�/���:���#D���o!�K|��}��x�y�&�Hg����.���E>�n�:{�~|us��E�����g��U��c9��E�홛�WN�wN_n�����N�8wT8+�2�b&�*%���֒��0:�+�Q[o '��ޛ՚l�>�s��v���+�=n��r�]vP���O�If�PU�N���E}{���w�"�������<��B�[�S7�s���;�O��.˸��/J�Z�@o4.cf�6x��؍b�񫯑F'�k�>�%k��.��|��?QD����M�jI!7w]��wZ��:*�C�!}nx�i�{0��5�>�ؽZ�r�����ћ�����Ct[�5�:�c��}bVm�#[u}�:����.ծZf�ļ���ސ�T�ڇ�M�
��p:����O�����ۍ�S{d�'��u�j5h8�r�jze�6��2�|�g5и�jܭ�+�]@�����XtE'Cʈ8��}y9Q�騍Pb���S�-�;hؘ�5X���l�9��շ�z��kj�������G��Z����,���7|;�����M��&A�1io�cO�^��R����\�"��9���B���]��n���T���2f{�
�z��{��o<���g�\޻ҏ���^�k�o}�iH�2�4^n'��|r���.�$�p�3z��+mѲ�������6ҹ1�2q��j#r�f���l����E�_6�v�];�,�W(پ�xd�ת���[{�5�ˬ�α��o�꾭��h�3Ea��a6���{a�x˥߾����\�hlU8��^G�����7]��oq��J�n5���]W$U���;q:��ָט�;�:Е�E���/�ƫUSˌs�{|�c��pn^x��	ƶ�oT�y��
���7��Z����\d�׫��%�n=ۇ�yr绣�[�܅�< ��q�����YRvJ\*-5��kqri@��[ϒU�2��Vwt髀�ʰ��n�-��&����^�nzS��]�T�fM8;�֓�nb�Cʞ�5�+Ȟ%k�h���ETsoU���%P�ȼY�����:��U�[�*��WH]�ad]�JL�%v�xq+E	�W�Q��a����S��=��,�p��g���L��Μ�r�
��U�؆V<s[�j7�*�yTۇ�M��v�e�v>�T�vM�W���ܑ���<��X�'�T��g'7��bΔ�+4�\�VEK2�+�$�֕�wd��L�U�j���X�S��qX��� ��Og͸��b:&p=��1��M%GC�p�<쓰ιC�<�n�����#L�pձJ�Ӎ�w~{��p�W�F��}zN��V��WY}�o�G�B�{��q�v
�.�V���+�O����ט��r�xP�GX�Y;٭ܲ�ǲ�Xp��{�z�8�~�[�����ܢ�b�������s��7_�n�5ێ�U'?K_O9����V��r���g��'''��DF�sF���U�1֗�������}\�+<��J���h{}�$5�ڻ�@���dQ������*�8�-�-
�57�S��{����F���S�������EaBy�ؗPU��bu��<�>}�hN��ҾAuG#�|�V����	�����<���o�Pgz&)�W��j�l#���UQ˼��j��ݴ��)�㨬�P��Bۉ5%(���jyOF$jyRޕ�n�N-n���n5e'�j� ���e��.>�z��ݶ�^^g���Y�.��}5����p�pOE�S�j�=(X�O���zN�NzJ�-G&"����w�?w%��ڼ~�����Egqȗ�����|�h�Sv�^U��C���Fgp#��ae��Bt�J�E�r^J�n�
Z13��M9V�%�wo#zr��H�9����:��><�1��4�������J��r�M��X�F%vf\�u�ۀ󂶡LE9��k7DU$�a�up.�I�ѫY��\%n^�,+�a�}N���2&񛧰��s��.F8Yq?+�1G���R�a���f1cۀ�zB�O��A�rㅕ�<;��V�	�o5�k���c��=7C���zm����X�|��{Xh#jf�j�v�>�W��F�v��6 ��i�օ�ZL����zNC��/�k>H)�.c5D�ԝj���:��V���C|}[}���q>��]���Ǡ������Q]*;��P�{w8��<ʾ49�L){դz�~��Kf�W�9�k����\d�7W���Kx��v/���N�Fu���=I���r/�7�+��oqG*�/+��Ν6f4;�QEI���eC�������M��}����n'E��|�o!����Y���O*��(N�C����»Jٳ��kњ�;��$x�G�P��qy"�=���<�����Q�̾сl��{�f�)0��)�;{i}������<�*\�
�e��Zc(]%�BYlh�v�+3s��߾����s�M�7�=����>܆�~S݉�{�as=;�N�͢�T �~~h�Ǫ�����/N5z�hN��{��oiM��[q	�T��:wt���ME�n�둏#�����]7˜!]^l�=-�{���R�Ұ�#�i�3o���aE��s��&���;�t�^�P�u7����2�+O�v�C]R�Vq{�T}����	���w��ꢵ��}��	X�]~�^�V9�+����"�bUʘ�����c�fB��÷F����q��.6�&������W�؟�˘�f�YV���${���ݒ���K븓]O�Q�ӸCЪ�Q1Μ�9���7���jrf����Q{�����:�#7�+�w�H�P�1�u�N�!�Zd����%>7�Q9i�h���sߟ;T��8��տR���{���u�۔̺@�zVִ�}*U��[���D%�G��Dl�̛�,���Tocř�@D���9	�OƢy2�F�*bNgV�����FE�P�ͩ�ݖtG[I0l���,��W�ꓐ�ޭ��4��h�7��˓-c�(���l�����/]
9�+ﾠ��ig���Az��*;(㺋x�/'1<;��[��U�7&��Xj�Rd��0�zYʝV��W-��P���^ߟR�>Ra���2wc��L=��Оo|�:j1���r��P�՜s㋶�^4�W�z�[J���a�ʝˇ�
����V�#�#<�(�v�r�k<O�bS�b�����:�9�Bv�DI��9�>����G�ޣ]m���Ĭ��ќ�q9:[�[Į<�G�ٴ+=&�����LN�_V��K|��T"�.���vF��Ӷzj��-5��
��b�%(�|��J�z�����7^��U��5����D���P
�W���ᄨ5nMIK�}i���t�[������j��(���l>q�{�v�G/�";`�밹�w*a:�c�sW�s�x��z�����_�<#�_�n�-�t�GZ�;AŜ5ldº����j�X�M(ǷsN�_f��/�ľر�R���֕�-���ڲ�&{����S�{Cu���-t�}����Pٽ�l�H�g_F͌�b�)
�|8)�n���;�eEγb{r��3��.�ţ���8�0Td�������Ե��85�~ٗ��)��al�����i�;�WP�11�w]g67\kg^d�u{�y7O}�@�m]�n�W���O����{e\u7q,��7�ڎ4�!6�Ө���Ǣz���xf#9��d�[����o��D�ةBy��Ē�J�+c.'���7_m}yi�W�.V2�{'�K�� w�#E�oMI��n�:�������K/����m彼��^�(LF��丝��t5�ɼ���j���}�y�-ؼ�r�����+�:/���׽�W��)�R�z�O?KS�o��3e{��G��}�77`!G��#q<�
l���-T_mc�x�^��T�w���f�>=N��4�<F�,���fxrW�5Q��!{K�UVWڛˇ�����f�R�a>�����f����nW��)s��Fʤ�j��/���UF��F���f6cf�
�]�bI+���j����:Ȼ�g�l{��MA"��֬�Fmo�b<��X��&o��S|�efhm�V�����Ncp4~Ҹ�6�%4z�a���;���y#д�s	��ʽ�mD��.b�M���]������N����oi��j�·O�us?f����};��;�_'���綂N�1.��(�'VL�R�����7��i�ì��
z 5n$��J*�bl_)�V�o=�,ތ�ɹq�LR�ͤ��n�ѓ�tݎ�*��	T����ˆ{啸�(�ө�5rx��c��i1Z|�K�m9R�wf`>���%�1�LH�y�M����p���PZ�:����y\Z�����pl�*�Ĥۃ&�Jܼ	�XW=�:I���=��݂��&�8<������Z���������,�a���qc�
�3=�f.x�j���g��.P�ʸuTO:y0��G{��~>b��(��c}���z��W�vAB��r���>N'�r��[��U��g���8���1�w�c�{dWs����A�Pc���RT=Gk������I�"te��<�>=ޜR<����GEX�B�vQE�И��@�âl�A����X4�78L�nI'P�w��&Lܚ�=��Y:�P"Z̾��m�8����Ö�Zw��c\L�Wg&.��Q`|�b�29Cn�l���n a����A���{��~gk�϶��[K�c_P�P�9���|�k���P6��s{���
uxa���9��+B�B��u/?QMuf�^s��4��/re�|���|�������m����~�8qv����F<�m�^�7:���d:�sa��B�Ow�ieC]��0$����֪�,�����I�5�o�����K��������3�*;��������'O�&�^�� T���S����72�U��z�V����{��Lj���4-����>i�4�E\[@^<��܏H�<�n'�\Ew%8���*⻱C������E���,�o^��4V`Gm�u({q&� ���;���]ܬ����I�f��M@c���V�-�"H��J�K"%?ԏ��]��w��պ��z��7o3�j��䖄�]���\'��aYS�5_���ח�c����}eqW´�&c��&`N�����PfsI�[4��k��yI�.Kmc�϶⭒��:��gmJ�v��FnigG���ٛx1��y�+3]oW\��U9>H��4����E9�mm+��-$F�F���r��HHXp��cL�\2��]� �ٱ����đ#���Z���3'R�޷�1�wOꬊ�+��>��X��F�cs�כ��gT��1�4�i]�bN]���`��ko3Q�ZOT�ES��� ]
�kMgvc�%g6
�֎}η�d�����m]`���R@>;)���[g7�	����[�i�A(bBITk@4	��:�WSpޣ�����\�P��EO����4���\��a7(�؋q[�K=��S���[q/\z���w1R,�v��ᓛ��EA�p#S7J�]>����UǦw��pܘ�U��9�E�ӎ�u'k���+��݃s�J��B�}���5���wmQ�,�zʢ�J���]6X�6��]ONl�
9q�P���pY�55�;l0l��r&�b�NB\�CgK�ۇ���2� 񄀠w*�J7K���
_ev���Z,gX�W�n(.�*;|ަ�˦�8�=�����d��Ӷ��,���{3#]�L�bfZ���,:u�>�0jO�F�Ј]�Ԩ��N�([��V�n��������`�8��f��b�hۥ����]׶hv<߸X(%.
��������s:o�N�s�C^Az�Sr��ܒV$��j�o9.x������� �K�XɪJk���w-s�X�󔉷�,t!��K}��p�R*�$�_s�h�e��墝(q�݊�1շ�33b6��o��Y��.5)vMc�t�N�-4�!%t���;p8[{w����ڻ�v79�s
F�1�,WN�e���Lr�'�^�K�K�:��w��O��<8�H�fT�ڰ�Ĥ�團[r3{���T���?�a�
[�[��J�$Mʺn¾=8�Gm����u�v;u�N+ob>YY�y��H3s�f�]t�z�v�����7��7+e�`��IoU�}#���Ҝ��x�M�6��� qkʋ �m���>���ym![c��p9ҝ���󆘵ts��qh�P�mZ�����M[�-M�Wάӂome[Mhu]�J��%�ڊ�d���؂����)�u��`oyj;���G8�u��F�l�ȋ�sN�̮�\��D��3o`�����s�����9u}6���l��_F��^���ص'5�/3Y�8�5)s<�6`P$6^�Ǒ�k]V�G��+H}�#�&��$<���N�ʚ������uޫ�]&�)��w:�P�7%�+Y\��e�&m�|e[E���tk�%��(cE����i���.m�}Dq��{׹A�����>]��0em ���GP��[w�eJV{/��X��޻DK͖/>�P��P!��Х��+Т�QPƫ+R��Q1*����QUUE�[j""��Zʂ"��[H�Dk`�XT�mb�UE+U*�1QX1H*�B�QbŬ�"ʅEkA��b�aiUB���X(DdQeam(�"��Q�EU��,��ee�k.Z0X�E�3)V*�֠��U�X���(�EDU"(bV,ưEҊ9e"����,Ʋ*ŊE��$b�
�XF1Db��"��PU\J�X��b��q�B�m11$�lTF(�QAb��Qb��U�PU���
�U������`����X�#�`���PR ���P+
��1%f	1PQ*�DQa"���QH�DU�Q_�����!n�P�f�z�칦Kz_@%�n:��)�����JnƮg&�v���7��(�W���3&<��4���Z�]g~����1��S;���欴��L��_GSv"a[1=!v\YV�i�ك6��]�UMvkɚxl���ہ�1�A�'N�P��*��Q<����Gt����oL��Y���y�v.�%�߱�w���y���n�- N��\\�&�Zy�l!S�8���ʋ�U�j5h3��+�k������9o�w�ng&)Z��w�OR�Uc�Oo=�Uã�-����*�������m^Չ�|��+��m���Lu�<��7���ڞ�k~������4���^��ɺ���2v�5���Ve�k�LS���]Q����?q��QPv���y]�\�9�o��OiT��T�i�������mo�߽���&�%}Ƈ����d���tC*(��)��YVsl>]V�-�D>MnG��3����۟�i�	�]�iUc���,�g-�MA�w�Y�VW;�kBw���v;{Yax=��p/O5I' ��w7o���9��M��Ƚ�O`��,𒢕�Jo/��vv�"7�w���ʛlr+u� +Qf��AŦ��g�wZy���]��n�!:nn�D�3C�6����!��-��X������^�{������#�7|�.e��R��}1��
Һ�MA�J&)�W+������L�NH�ћ�r�#4��7�y���au��9T�mĚ�)p��5����h�kg[���������OE�:J�;r�\#�TI�ϨbG"�m���19O�oK�R'9���^�_-|ٽ	��٫C���Uś]G�Oc���X�;8,8}}��ކ�]��+c���_[�0��pPr�l]b����
	��5�1H[�_c{��W;��ML�P�|[�\�W��=�E�=����ȹvټX��xg�X�Փ�AR�hv�,��lW'����ʊ��8�0�'�9SqR�n��˝��U�����i��"}n����Y�Ѽ�-n=��Vۃ��t�w��y~�=�;��Qy8 Q�K�Q:�QS���}�Vl��d��+]8��#�ne�Ѯ�Aq�G�L���ڌd�&��B7�Np��X�4]��|�qb�cU*�,�Z��W��o"U����͚�C��%u�)C.�6�.,B!A�rr�,���U����QN��`u�����(��ou��^�Vs��7�:bu�Ok9q��A�Y�Z��"�Q��o�=��l��U|��19?;���iu.ߟP�z��<�����O����ɴ;�B�윚|����փ'��r�.�<�ulymՐ����r��6��Mp$z�?z���^��_3B%p�q�3x�����o�g3=��ڥ�n%�ܝv�k.��S���ϒ�K#`��
�:�jV�Qg�E���J�y-F�����qUWN1r��oj�e�º�Ī)Bۚ��O�����U�4����6ʚ�����nm���{Jm��<�p�t,#z\��-<W�ϝ,���{i�����M�c���:�ҽq۷FKt�u9]a.J�.7�f\��o���S���7���~]3[�ސ�z��ܘ�H��u<�j^W�Wv�)��i��G<���Z� .̰�n���ގ؞q!�"^^j��}|�uF����b~W*b��uk��[�p̸
���c�~�}/1
FǛ�Y��7/7���:����(�����vA,`�8�Ĵm�:ް�)2_1w��
B8�wΧ uvTJͲyܶ�����is2��3�8���&<è�멑dޝݱ`�pJ.Qx� ��(Yܮ��J��\	��D����ø*��Wǡv٥������3��ˇ����R3k�&��-Ũ���S��n�\p�*�<�뿍>�6��1^n�O���U.̌�%��3�woHY�������*5��/�ܭ@�k�|��z�7�,�N"�V�j;�������?5c��L\�Q8E� z;j�p�0)3��;���^NTbzkT�Q]�>Ghwer������so�/`�/�ɳ��A��Ҩ.;�SO髨��OԱ����܂D<gn�[k`��57����[S����+l��Wg/�^ڥ�:������&gMn�m`�����x��D;�n�k�_,����:�&��kKo I����5�v4�SG[���m�>��t�|��}Q"z�ZDo
X��Vw�w���U��P����w��iO.��i����.0P���^t։���]��j��3�[oM��q��T��Pr�N�ݦ�6*T����i��ʄYʥ轱8e��۔��.�]��Z�/{�^�K��Cr�Vb}��}�ubt;kyҽ͛O��]!S�VA�Ng��]�+��x�|�<�:���9�_���Ό���B�De�'L��-EI�Ⱥgճ�o�t�^�}�v���+�(倫�pgO;�CR�W&�t�=<�˦���ޓ����;+0��˶if�f+���C'�t�'.T`K�rͬ���j�"~���:g�����;�t��2m�ܞ|�N�͚�1?&��%��Z�Mn�.��jJn筆Z
����˞k��_S�I�.㛡��=��/�#y;�(yo)k:���̧��fthq�y9ݙ���PU�;��C����<���x�+��e�=�������6Оڻ�}�c9�כ��[]G];ZJ����⥕sD��;��,��Ux��h9��u����JM����}�{_�U�D�Cp����\w���TV-]�5��^����Ҭ{ӊ-�;_c�5�ʎp7*�����qM��C��#���X���K�h��$ި%a�B�EX�F�+��x��c��^�Tz{Ǔ,�@'�$��3.�.���ʵ����u=�GE���$�N� \坚�� N��N�v,WPލ�XFc[�
<��ƁT���{���*uc���i�4}�����_��W�+�<��kRGK*�������w�mz)���߻�w"�~�8���؂����5s�{��9��E:��Kʍ�]�S�n�65��Y�%tj+�i6k
�/�Yj��#������2=:�4����[��!��S݌��%��{oB�Hg?�İ�#�PgZ��ʢ��z�hN�1�G1�l��p�K�z��[�SٽV����q(%6j%(���^gM~|>�[���0�{�����4n�]Q��-�ov0�B�L�Qm`�Vl��[���fF��iOSQ�W&�C�޶����FLS���eVJ�F�#��5v�t�洨>{(�����]5���|��K�z1T[����5��UNM������t����}���D���ƇM�Û�[nÔxhR�]^!�w5�EY&H�M bV��b{����4�_}�^�$Źڅ*�K�tnh6*�.�;���iU���..{������s�W�G��b})V[}]j�ևR��lc%���-]*뭶�mnX�hIڡ�!�1I�ϸb�y��n��j����|F`���c���)�nR���թ����ʵ5�����LQs��m���6�!y�;5��T�i]�E����m�ov	�n\O��LQ��YQx�<�{5��N��k6�)yg��.c�OB@���@�S��9˕;R�o�O*�\W�\�onIAŗ��Q�n{۫�ٷm�oT�nq�V+��+�>{pw�_^/vu6��O����  �WN���}�I�%Z�:Wm��j��p3�}&�S-��r�ѧl�q8�j�ݸ�P�z����?$��{<҆͞��׺,�Chz�Ϫ����:���p��>{��1.�TtR���h|��8�����Y���+��Y}J��qʾҲ���t�D��PS˙�.���s1��-�}����lJ
�퉨5�U�V0�35�x�*R�i�7��寓ݔ�|��yPZ�"uDN���@"��G�(���PB�����:"����7��۱�V�=�[Tt=p'����Q����-��Oj�me��S'-�8@A��Y�b+���*���TscaĒs�K��܋��ϧכSbpZ�9X�p����8E�����j�0oxeͮ�F�\�5����s�t%Ŷ��ԯV=b�@iVĚ�?�걆�7*]������c�8���:�m+����}��P6�kB��{5�s���*�����JH[��C]=�t������'�,a��Eew7���Za��=;�Շ��Z��.̄�;uW�kp��|�IV7n�Z�s��s{�]B(��W��>%nd'w�Y.���)�7�v�7e�<������l��n�Ә߄������n�=��@����s3S|�m�؝�p�����*��U���~���:��N](;�R%O��#j/}٦c1�{�F��mA�jq��X�Z��ۆ�i.�ɖQ���P_͝��xz=��
�uO��|��I���C��0ܔn��j�cM��uI�a �`*l�z��r��Q�u(��x�yb�7-�<u77ϫ�Zc�Q���eT�4=Eo�q!M���}�����F��`6�
e+͇[m���m��os�ǌ��.^���K�i��˩�,Xo�[�f���7|�u'3�䤩w�88o��Ӝ���4�Cº�l1��̦�R��3������y�B�iY��}L�==^&z����Q��y�^�0����#�\5Y�(���!w�5ѓn.�;Q�"2��wlt<Ow>w�Pݭ}c�f�
�f*_��8��Ci<��������ڳܯOOх�p�}��W�U��w���B	�V�2�{d[�u��m���=��Ɯ�7��&W/�J�{OL��:��>\���j�S0��5U�J��J'��joLE<\wDb��0Q����2zz�5ۗ@HO.�XVZ��	CP��ߊ\-s�O�c�����my�VI��eL%u��qf]#Iʗ	W�9a�pe�$%ۻ��s����?�5�/[�Z;���n�b�b~����i���k��3v����m��+�\���m�&o�9���=���*�!�i�C*o4.Rg�5J��ud�y���z�����j�u���,���[օ[C��ffj�ɫ޼��v�\���6c�IJ�S��⾎;�%��xz���C�*�-����)�I
v�`L3���]��n��`�ft���;b�n.b�>Z�:u.��9���E9��t4�*�8��P��{�x��:FǶ�!�3/��R}2�v&k5��	�:��qL�]]�̺[��u��	�۷������i�U���9o:7�*�6�7��ˎ��/K�ۂq̜jm{�ro�ё�EtS�Z��]�Ը�}k�jf絧����rjf���㰬V�[�e|q][ŵEbߗy��h{A�0R�x��Г̛�ŕ���q���K^�t+!'tW=��)4_+�뒱%^�~{�y؁8J1j�����Oz�gN;;���⯴]l&.y�Yv�归� ��/t���y�ǖ�Muf�^^_w��B�?1�W����v����	\�j�qTY|�,ߵ7����q�֕��y'.6�6V����@�R�����j&aD�UyTY\�R��;�*�w�t�\��-�J���þ;P�9\@ж�8�
l�J)�VV�g9���s���+��r��2i�͸�K���y��a�����a*�5nMIJ3�j��eN�θ&R�Ow�xyJ���s�P�mV�8�F53�M�������j�ݮF���o(v7-��gl��i��+��:�s��%�zJ'�r� �W�m��wR}G�ǧc�0x��c[N��Yۖ��N���z�����R�<�nh��8��ې�%V��Ki��s*M܎|�:r�]t�]u �e�9�&�=v�O���똕���'W��̌�|л�ڬZ��z�r�H\�Zݫ��U���fy�[��f��E�V𗥺��ʽGK�Iս�{�����{�S�qcrޞ��tkn&�WQ��)11��E�p�v�;��<��Ry݆�`��z�T��0��ٛ����ۚ��P��x�F:��Ŝ�4!;SVs̝c��q�����D��n1��zT�y*���v�o-*�ӳ�ʤN��%�9.oV�R�V{�$'
K7�x��:��|Eg5-Ab7��߻k=� �
�L���V�l���9w)ksw����\�Qy��3+��֮��v�뾸N��5�7�R�xu)�uֹ 4L�K��[�C^�$Dc������YL�aVAF�����Aě�;6�5�����܃�r4>�'��"U�=7��8m�d��Y�wҝ�0�]A̪Q�*3O��^���	����&�������+p,���<�	*dp�{Nve��m!�ݝV�Y<�������ǩ]��췒��g`��-"�K^����7��Ȗ	��V����燗p��u-�.����Xb.ۧ�8�s6>,�dO`��	�M�:�wx{�����İ~7�������O9��+���q��n����i�b�� s���V|:��ն(�}1�]�-:MK��u�ʚz2w+Q�@�9\���2�V��=A�C��v�����/�;���x��s�k��%��z,��V垜��s:����h�:�aWGp8�_�ͻ�������'x�u�b��
缤1G�w�.�R���� ǄK����%��F�|��[�m+��W����u��\a��_E7 �1(L�n�(�d r^7���Y��f���S �}sz��]̇�HQ����PjS�3X���὚d,u!�ē�X�]a���=�)9r�e5�8��
]�,�S�1��f�6n���P��+
��-�M���[�8�Pa�Ҹ��cnhF�-J�R�u)�Y]��]}��Z��h�ʡ��Hۜ6:���#�\Q�)�2����ܾf���S�����m��)���Xo��SPǘ{���;r��lŵ����-Զ�$󻻯,����1E��n�l
��*�LY���&Y��,U��[{Y,C�Z�|�Xg�����˻���Z�v��Vww���94]�˚Y��ږ�V� GZ�v���0{{��ϕ	ڶ���`5�?��(}Q-�H�j�b���������k���M)`	چueu���^o�b�����B.
vqu�_1n����\껝|،K��^o��9A�:���4�
������1��x��H7���<�e��o�í��
������B� #D}AX(�1��*�Ȍ��RDAT���V��+F"��E���**���V,�+H�0U��X1F)�*M7T+R"E��TP
�
,X*�UdY��X,DX*����Y���:�1�
��T�PY,`��X�1���(�EF
d`��DdDU*VFکd4�AB.Zi�b*�V(FЬ`�j(*��B#j]P�(�U"�b��b֊��H�Ab,Cłԣ�TX���TEՕQAE�)b°���*AALIDb*��2��`QE�(�kH��11Ȭ"+�2��
(��UdX�XUA`�YX��m�M1cl���UQ�hň�Q`�*�j����"��QcE����[X�*�F�*(�R�X�V�aR��E��(�R*��`�.�:���__Kнԣ|xff
���nH3�q��Qb_ϩe�0,��jÆÄ���QIڥ:��0*����챩g�u��937�����p�X�Rx.T�@T��
���{v�u9sn��S����Y5k��>���U|V��o8+z1U�
ʞrfu�V�:�J:��(+����Yave�N~��cWR�cZ��NYrZ�C��=a�!�[�'�!vY��L[�Q��­�����L7X�v͙��x�z��ElbpU¤�%]9��϶�������X�g-w]}�Jɥ�fh!ז��"�k��I���m�[Μ�����#|��mQ^t�����V��.�A��A���v���[�5��aX��+�����d�T��t��*��[�Ґ���nNg v1A�����N8���]�[�+��r����"����\�1q\�˫�u���F(�GTOe(�x�j�s'�����a����}��n���	�%~g�(�~�9�]��v�R�c�h���Ξ�w\��Rw��paڵ{�"4²�K[X�7�=Z��L�0�� �,l_h�y!~Řpӿ�uZE-�"�f����i���������{n��� �-J���#���]�R�|�`CU�L!�C��V�@���v���ܴ^�t�G��.�vn�������I�3O��䯙J��8��my�T���H������U����t��Ou�M��X�9�+��;�lJ����1Z�}g�E�H�Ͱ�_U���Μ��.��-�i�ok�5�6�.��(.���tN�O�Y^����i�%�w�x~��j����:7�z����J�N��eK0�\S���c�9T��o�:A�K�R.��L�QjS.�6�W����Hz;�+�{�����ǅ�9�Gw�Y�����ˋ���@�L��J�, 4}k�j�/��?JG��\���Yni�x��-�]��m�<B���F|嚇q$��� 7�qJhQ}^�G3�ơwT56�h{s����x��{0�s����� �3�dSʧD/I�a|`�eD5DM9�;� ��Z_���Sy媧ˋ�g�Ǳ#P�����x�}&����z�1�ȇ_)��t�^z��tU:��0�l�y�`>�2=�<�g����T{a:���Ǽ�yND���R/]z���7>G��TO��\��#�/rz1�E%.��0�ꕺR��{x�X��*A�z��}��S���NQ��E[	y&~~�8B���y�:Wr���2�נ2�]*ھ6��7��y(�X��ԳS���D�
��!�42�����Ib�{я�B�����Q�t���=Qʬ�.#���{�'�C2Ϯ ?m� 5��1��>���gB��ϡ��g��댭��ͯq��O5�����29�q�'�ׄ$=Z�n��K8�dW�Hݱ,{�z$���#�;P��{�l���zo��-S�/oeƱ]0f�t��.�]�{��5w�H�|��r.<����QD�;;,e�V�+��,��nf�lb���|�N{`?bVE�V��o�q��y⸫�i���z}�����2�kKH����ӋM��n�s�7OA�U1�{�����B���S���Oq��z��w�ֳ�	H��n����.�`H
^dm-��eH��9Xt\dΣd�E��2i�3��#��#q�\n|��>0��3�6�u�t�WGZ߂���U�<���
�� 9��2�e��ua��~���}Ǳ��:�̪��cկtz�'b��>U
��|��'"	@=����4�V�x�ن�����IhU=�/�$��on3�݌���f�Q*���eK/#L��ϥ�2.�[���DmCE�W�bj`ȩ�BsşD�\�ˁsT˫��-��=�y��ց���C���������\���g+x��i�ղ�j���k	�hY�*ޞڜKv)��u�-$�9c�t�z�6Nְ�U�����N�\|WS�xXwL���2���V�yYd�ݣ��|�*���,�Q�Y!�ߨ2�w�tW��w"�~��Hl����"˟q��k�W���B��Mw���%ȭ+�����P�%����8�r=�]�ȧ�N��'��(=�⨇A�@��f�3ΖMQzOq�8<zV��|1/R_O�_��_�TD�V���q�&�D��-�*���to&dzl�M�{n2�11MV���Ln��X���H��F�u�T�D�(DתҼHA^<g$+�	��4��������\�}���Z^�WO����bڪ�ֽ�1Q�nMf�������D��A�P�Q��W��3c�o7j�׸���}��=Z�YVהo��X�k)&DUJ�h��T���g���L��|Q�w�J9s�i��c/=Z���w�?W/�0R������}�~�~�y�����N����ݸ����:m�O�����1�Cݽ��W�+<��M�=�
��s��޹���6�W=�y����:�^f�9�����s�.<�Wq���r�(�}廫sV�Q�җ���_d֔0�g���:�{o:��*�o������؊��K��<E��t�G��}4"�Y��-�.�a���s/cr�K�7���r��/��oQR�.X՜��&z7Fcb;�rU�w�A�t/hm_�v9K�-�i��,=���H{;W1��	��Ku�����[w�U��XjChn�
:����:1WY����1:��Ӧ;0Jd��Oz�=����:��L�'��!�������ܝ��j=�����J�tK�9e��"���T��*p79�ME�?Wz��L�FL��r9�C�Y���y�@��?u�����e�F�l�^�	�+c�{=���LӔl
n�d\�9f4 �AbpTv*���bͲث>�|����|��Zm������ȫ�Ul� &z��o"�E��!�;Q��y^�O@�)��Y��/�C���m���*�r=�tߩ�>��4�l��m'�u�U�R���L{�/UHڙL�8}+�4�%��pw<�x��r�� ��E�r�Ew�X3�=y����^µީ>��BW�������D�>�a؂Z;�%�#�|٦_��x��Q�]�>����q�|��=̂+甦�Z�^G�d���bb)�m��{���Q�¼/T��=6�7��oه��XCӀ��{.j��>���lf���Vɨ����_a��=�׋�Hg��V�z����G{ީ���<�D��Ϡ<�/W��ȹ��"n|76p{��\�aV?T�Ғ��MR]ff���6��52[��q!��ZX�ų�P�4E�[��u���&�
�[���/��vA{eM_�A)뷷�sS���=�\+38���5:V@(P�$\��*āD����3��đ7�71U�T\b����^�R,����Χ������g�2�}�������$�J�6�(��ފ�7���G�r�}��/ND~����/���U~�W��kk�}��?)�*�2tV��T�f��`%^��߹�� g�T�O�&�:�ߙR���بo>��4�J9P_A��3�&��Ō�8v5���`LE��d^����=B'zl�d�FV����F�`���+E�'��;w����+jzz�k�5�T���`_en%;Y�7ƥ���s��%\�y�ý�PP�h�����iS�Qc+�;�&wӃ�>3�+���v�_G�����[ӑ���߽Q�k���}墐Y�
v]``���&�����}�����X}��P{%՜��51�g|�9�qu�9��R;�q�V�5��g����n%����$p��I��������S���as����L��U~��-�=]��Oy�X]R�vU[�7�%L�V�s�>��P��S>d
�R�]gѴ­�_�y���'��D>�5۔킣�7��7�ܽ�PW'd��t}�j=i��7����R+Ҭ�����j����I�E@��1k��,bD72~��H�:�H=�R �� �WbW.�5�oy۔����i]�RI
:Xy��9ǯ��p�;[��M�n���]�P"��N�	��"f
���˫�nbG�el{Z�.�{�L�ʝ��,�'���p�R��pg/�Ru�Ԕ���:2���9Y*/��E�W���@�>s{7�)�E�{��ϾƖP�T*nNL&kՄm���}�t�ѿ��W��z w��"�U:"���>,Y���4�／��"�����%����'p�w�*=o����IQ/(~�X���E��<��������V�u�S����e�����"��Q��*#9`�y�U����K{�����EѲ.�����vix9�݅�r���V���C��:���Ud�q�z���t'���9���١1�5#��{�,r���^ �^@���Ԥ{>��ו�a�f׸�Gzx�`����'v|A�"��O�+�vo���{]5�?��Q'!90�����^mV�ǭ�<��Z��.�����t�s�vo��.U���%�ݻt.#��Z/����>�3I���V�+���K�>���ߞ�\rլ֟���=�`T[��U����9.��g�{|�=�;Mǔ�*e���:���]�NouvA��^�2�1{��|d{o���߶��q�d��{�ye{��}��zQAo�EWXJӉ�Gt��>�u-����i�]ݺ `U�h�U��]Q7��B�,�Y7����6��F��t�\C�R�	Z�Y<��rԺ�;A�ݖ�99�0.�t���{&.?_wV����v�΄ky��k%s��MQ�l��+�+��fm�}s�X�ɝ��/":d*��>N��m�񯟯C�V�Q�<�o}	��+��/G5~9&�sqU�LT� U�S7�,/gS����^��=�}Ǹ{���W����%��T(��՗���8=q��+�l�`>ȉ��܁��x�ن��mC����r��b''=���Q���u�,wz<���z�.��eo���>��9FE��e��{s�صcݷQq䷞)I+ݹ�M�f��\�֑���#��{�����.��\i!��<��#������;ӣͨ��Pg�G|��3e�Q�P�__�G��(�{�x�EM�s.H�'̘���i�^��ۡO{=@Ǵr�Ui5���2���3��)�+��e/L�D�r���ྈ��^�=�:�����WAyQ�B_�dD�C��)�MV��|7{�,eo+�X����P��(ږ���^�����c��?@˸�fi�-50�c+tø�WI����|0.V)���έR�y���ę���}�����x�y@TB�IG=3෌����ݨw�m{����>����-[����U��p�I��a9�%E����Yw�ԬOM�qde	�;+����pc��tفÇ(ж5��Tڼ�4��
����fRw���ﾍ�V�Y�0�m��ƺٶi�Z�h>��W��/ �CopՋG��
aO���A��ҹ�\{�xw%��,~q#��;��x���t���S��U���QˏU��,^�C�c�W��^���~[�KR�Џ�7Łj�Ǔ3� 8�u<n7ے���!�+�����J+��{R�_�zy��^����]���i�����א+�U���.�[�G�TM}�W<`��G��2n�����o�o��>�}#�!�����O�,�fy����*�x �*�m��u�w�у�W��%R��� *){�ʖc�����c�w�3��L�'�R�~�i����[��G,���r��Whh�G�i��S�͆羚�k�p��n2e���3�\�����I�q[;]���_W��GB�Wᐧ(���P� �`>���`Su�s.$ӏNe�9�[�ڑ��Mᐸ�م�.�9�G�q�t�7��=~�YR��@l��� �{#�g3<��Ϸ�k�c�g�+ ��/K	F�_���1莝��u��~�[�x=����{��}xGE�0���c��B���2��+�3���W���;��ǽ���q#���=�6��x��5޼�����:s�A�ֈ�k�E���Q-����w��:5���a#q6��gmi��g�m�(ɺ�%�P[�������L���Cb^Е*�s��V���fU֩:+�����l��6�r�6i-�Ґ�)����P�!-��o�LLS���%���X�)�>�����A�I��5{��Z�WU����ր��u>�����sĀ��_���>��z_�v@�xg'G�f�U{s�֏oPo���H���@{�� /z��y~��W���͆76Hu��9�g�����;��L�;��G(���q����\B�m�/z��:�p{��@Wϧ�]]�x$s��Ӿ�l���C݌�ݼ��]�/�o�mp�,i��>�噐�檧��qS�����{ <�f���C/L�	�_�þ�>zn���r�}���Ry;�ד����|�m0)+�G�Bu��ҹ��ڱO�.�W���;X[TV&Y�n��$Z9�;Q츌�qb�6kM�7�,
SL�����>�=�T���_��ۺ1�лo�q��Z.!��s�Hë"*���ه���7�}$xebX��A�ں�f»�E��|���Ut?Z9Co�M��n�gn'Ԇ�9�2�]ü��Mg��zr{�w�Z=�>03���~�{
�K�]��⽎�WyPE[��sa�*�7�Ͻ$z�3�z΃�M�0}�<��*<o�qV�ɹO7��	�R��@���pЫ���eN���aɰ5H䣀S<_N���b������=���F��\x�gn���B�TY��p��0��nʳ{�!�G�*ŭ#]G)Ħk��6�:�q"��C+�W�K��3w!����扫b�O5�E7�2'��X���f8�W
͓8<��u��q��füG�bV�5��ڦ���|���#�rs���ǯ=��(VN�AX�h�U��ww�«@m����0s�CW��}sS՛�$�h�ڢRHu%LO�+۾ٚ_\	z�Ȓ�T�Jj�V�(��4Ԭ�v5ge�6o�������nojc{��Ve��ۦQ��P(���ꂢ���^]������"���d�����JH�K�;��w�y3@�7ٴ�d��$87�!G�˙�<��Ց�tL8o�ޜ �5����⩭ݾZ��i�gs�o8��Y��@�E��Ξ����t�u���-=9�@s�lu��	ʱ�#\�=��I��4�˼��qtde���K�G�{�U�=�B�#���c�)��9�f���A��8�����p�ts`�x��[}K�dݾ��,������s��42��s�;��F�<:�=��'8�\�\�@Y��věj��ꣷ�c�;��M�g]j��&Dt짤��;MK��1�aݣc�5�h���Mo{
��Nw��R��������սW���Q�
ʝ�,ݴp�F��e
O� F��7�u��+�+F%ޕ��v��@�7������d9��� �Y�s��G��+��k->��gS���e�/�xa/8U�u�N�HT8�Ң�L�8���Y�����ȱ��+w�
�d�R�+E��
T�K�T�b��sf��:�pp������jSQ�2�vL�&�{��;WK+i=��t n�3�^��G2�օ�8�f�����R�0���^�w�>ͧ�uk�sց֯�p����	�cRt[���e���ۗ0�`1�yy����bEl�0[��1,��N�t�>�t�v��jƅ�ѽ}���c�
q��~]��o!ipʻyE�Y]��S��B]f�p*$�Z��۠�Tz��g���w ����9��1�`���V�Y����dN;v�G-�6R�ڮ����$2Z�ɹ�ҕ�M&f3���k��u�u7���^��(eִԴ_�Cy���J��7N0e�م���
��ڮ���j��e��tݝu�>�zhq��Lt�|�Xn	ݙ(o~Ɂ���,���'jn�[(�u���ӣ[:�H���ï��X\]��bc�6���Nn�\��Q�.����Se80u<�X���*�yƟ�7���E�n뫵j��ع-n�WM.����,�.�^�)6J�5|�5TQ�H��TƂ1b�X#"��$�UUm&8e*H�V��`��cb��,R
"��Ȩ���@QQ�����eT�VID`��Ȩ�b��Q`�X���"ł0Ri� PX�Z��DAC�-+�Y*#UF5������T�@Q�5i�"������,*c���XERk,1���VKh��(�S5I�Rj�"��PETAEձH�Ɍ�ATFTb0b���Q�U���*����#�QU`9`k)����1��0X��X
��T�SVHTc+RAT��V�&���E����YP)�KJA�|}B��PM]���G<���{�4�Lt�F��v�)��mmIp�h��q�u:��	�]ۑK�8�<��5;uj�ܺoP���1�ɔ��9��9�x��L���W��V��
G�Z��?@��������J�x	^��b�̊�H�q�({T�5�q����q��9��7�=q��/xY�����'��y�s��Ee����S���U"�l��jW����Z���~r�z��ב�'����?R͆�x�臗�g�^:�z �j	��UHB�z�%��ͨj�����(ɉ������)e��#��mx�0u��ȸ����8�|�{7Jh��;�wk�]�졽�Z�wdy���~���?r��0rXW���]7�yNH�^��Ř>_%DK���=ٝ#�����n���0(9�G<
Gt��K��w�}8Ϥ�r���p���B�!��U:�<J�:rY�	��!�IN��致G��i�_o��;c+�V.s驏{U)�I������y��O6F��M��qn����G�NT-ͬ�'ä�Ѯt��=Q��b���Ǽ�Nʠ��������[��}�X�˃��;,�*#ށ+Ǫ|�d�G�'p��ͯq��O5L �z�2�?uQ�D۪h1�\Tzp��ב���Ï�)�Gt��`��,}�;Ց����-�%GM�7%�kw���h��3Y|I���>�<m�Z��^hFl�m͠;`�fj���3��.�������t���/�n�uʤ�����ؗ9�� {/��0q�����w�����z#��'�����^Rމ<p�B9�;P��a�L�Z_�H���Σ���Z�$O��gX���O���v�з��{&x�D���'K���	iY���k(|��W��|��ЊT�p3~�vZu�=[��#q��7�s�ὣǁ�N��of^�߰�6�Hx�{dx��Y�}�:�.#}!9�2=��}�<���41���p��l�YX��4�T�M5��y��}��UX<��:���>E�L�Qg��c�#޹��[�0��e7[/w΁��^�Y�x�{��T�˜E�UXSȁQ~������S���S�h�7_^55�95X���)=�g=����H1)����T���욋�?StE�^.�6��S]��OC�3�ʲ�7G+�v������Y+޿_��,��!���`{�A[�UuI�k�W��H亣���3��c�ԑ�z���}�p(�_�G�r|�d�ٸ0[;bo1�TB2�j2�{^n�!Ed�ә�ϼj��}^�7���#
���*U: ��� �U(h����æ�ߎ� <�cSՇ�_)LV�Z�{R��Z�\Q���؊��LL��җ�{ė���'�x�2�¬.�n��ۚ;o��7A�]���C4��va\}$Tz�8�%+����9��ǈn=��u��{
.����ȫv�Ĕ���"���L�)�tdJӸ�[��Ƿ��;����>��?>�y�ň��\$�A�B�s$
���u���1?SU�n5χt/~�Ud�i����(>����w�z��Eo���K�Ǫ�������#�un#+tü�t�����:�4t�	?M;���pg5�������3�z@<�H~7�lu%���^�͏i��v��m{��Q�vVd�Z��ǻ�V�����GTw�~̶1������ު��w&���J9�����/47c`�E��wq��^c=j��A��G��Ƕ��)���ʉ��5�����z��[ :3oo�ﺝ�,�>����ɭ.��b�޹�,��� TZ�o���~�G�E)�T{�uhIO6:t��
��Bs�=�)��R0�Ȫc0Ζ7���r�=T=�L1K����ݡ�*k3�ҋ���<;b��c7�n'����UG��ъ�'Y�g�<���j�A�Z�y�s=S���o����uv����RP�7.p7&b���C6'�&=����`���,�Σ���މ��@�b�2���.Nݪ���F1�t	U�x����&��p;����T��fƄ�����β�0-r���.�(��Ψ��g#���aj�;+67Mqk齽��"�ָ�H�����ė�I
h-tms�[�r�;�m��+�~�~�W�숿_��ìV�d*��_��X��M����T��
�}]3yeI�a���z�e4^F�#�醣����<wO��/՞����e����Y=2�|]owu�y�m�K�UH��t�����>͖D_V�'�l�}���x��~�P�G�i�f��j]Я�60��|`����ex�!��x|9�Wq�P����E�3�p�+�W��gu��b���]�yNn@b|͘(=��LM>�i�%����R�����Ol�N|�Nz�*ӆi�]{t��0V7��=�w*!�znª-OdL���_���O�hޗ�ݭP8��xz6��w*�v�4�/��Ц/�t׍���vAU�o�`��@��W��h1��C�.3��}SW�З��L�i\U���\�Tz��͛�y�D���rz�Ԧ�e�ӦΘ$'�6�>�@�A�֏^N��l�&MF�=س2|�T�b�\N�~�V�`yF�>��^�7�GX���<}��ǲ'���ͭâp�?���uz�s��@�=4g��_�q9�#j��z.�'e�+�G� ��lQ�����f`w�0xin�B�����(�v�b�̀s
�ժ�\�N�h�S�p�ڝñN�]�u��|��t��s��.R�s[ʏ�r�>�ϵ<t�]a�:C]��DbX�C푛I��'M��4Լ�y-��=�������<��/�Q�@�_Smm� _��:��C�u��ߺz�����Sq�Å���Z/�Ew�Hë>��xrva����:��G��2������<s�h}�@Rsl�{޾�)�4��ݢ�dO�F�9X�UP�FCؿNW�&g���n��ҩ�2�{��|6����#�S�k��������RQWh
WV
�����]]-����yR�5����td���3!����r#ޗ��?�fͥ�np�o�xy8KhV׶5HB|�)�}�U�1SȊ��������~}T����aQ���s���f�xA��\�~��+�F;�}'��P�UH��e�E�^.���aT_�G��y��;���h/�k��Lߚ�5z�q��g���!�_�=����J�, 4}j6������=ٯ#�+x窍�D�+l�)��PLW����f��2O��{7��|_W��mb>���/{����x���@��5��q/��9�\
Ͻ�����dSʧDZ�,����i���0��Ws�N�b��yI���T��#[�j>����Y�U�t���ƭ;��)9{TP?b�]׳��
��Z��]ZG8_D&��A�����O.�5I�۽[P����e,����+��W=�]OuS��v�T�1��c�Z�3pC�=���r�V;�c	xj������>��}$�$�<�ꨉ���z'�{ԧf������e�n���D*��i�Q����^����'^�����C�r\�{�9�/�ޛ����8�R{BQ�����Qw�V��Ky����=�tܦ=�)�X��C�kLx�Y��.�~��4q���^����E��߷?p��m~���+�=��%��[L-�i]�5Oۈ-ҠR�h��UG�\���"��!qމ<r�}A;0�߶a�L�KT�����㚪����l�>�W 's��Ns�_���n=۷B�=���mJ<��њN�.������ك�^��h�QX��k�n#O��O@͎�`W֝o�W�Q�|��)��y$v��#�N��Ƥ�=,w�޴�1���\���ώ�?_����Ǐq߼{�}�7qگ��x}ً{}���O�����p�UX��x�q�:��^�9i�3�?:�=1J|w���syg��:�<�F��g�W��������ES%�e�DUXSȁ~)���a{":��^>�����~ݙ~�Bb�'�pu��I���n[�v����{H���c��+�^�Jwc�=wV�}e5R�d��`�9v�i+g�|�}��v�Fe�^�8���ȏs�������D5�	}M�D��f�0h����W+���Q�U��{xJ��߬��������>���ME�����*>�+��Ǜ�k�(t��O]��{C�=�н�q�e#n���F�����VD�,��!��>��r���ۛΪ3�˘��$Vz���{j<�}}��REG�!g�
�:����Eƒ;�E0a\z+��ESYހc��z*dLA�l��i�/ƻ���j�&��ģ{�4��e��\�B��W&����U�z��|3�0P�ʢ%�����V����ܽh{>�R�La�R�Ϧe�z�j��{B�\�2��{��M* \B�>G�L<ܯ�mg�w�amR�P���N�~��oV��UΧ����@�ߊ�@��K��UW����3K[�K��Tǘ���U�_��}yC�Ҵs�8{��!q�UO�Ǽ�,����9�y@/A(����p4=�sv��a�򯙏e���yNݬ�,�\L�j5	�_�6���g:a#��\*�6j;�%��	K�
*���}�5��/dp~�mhW���q�3�o�V_�=���x���}��7۷~��ң�ⅺ���z��7ޠ�]�<�+m��J��{�Z�[�$�\��9��Й���Ή�7qh7d�sE̩ܚzNPQb�����V�WٚƱ��b�����빍h��Y��In���b�X.�\�X�}�U�:\�mL&O�JY��z0����&��\�ܮ\D�nu�t���yfYr����@J���Ef��垺�q�F�o�XF��+�_��������jW��$Y�^����pʿE���x�{�1~B�u��n�<>�,�g��{Q��:�{Pav�����s��5u>�{�}Z;��Cz;�r�_�tSg"}:����j1]1q�:��L�'��Ywp�K�]�\o�h~��zw�י틟S�� �������-I��j8	��û�;1y|��h�8{�G�3���<�w��^ӑ����z�4(u���9E�Ͻ��r�{;���@�+�I�{��2=�{�.\2+���$o[����>�{�Ǣee�*2��5w3���::03��PdUH��`d\��}��¨��?Sfw�W3��6>1����^��Ӌ���; �z��q�>.�q�:���ly���TF΅R�Y��>�0hq�ߗ�������L�_�M�`�r�B��n��H�����8KGw��{'�C~���k�dꔅ����M#���޽�{2�y^��j��=�L���E�LO����x3�x]Gz��ut�2i"�iA����ʖ��'�aή���l�V�t�����ˀ��b�Vb�%N;����αab���n��9�{/9�yAo=OY�<U�2'�'E;'6��[j���5�4�=�͍��4PG��W]S�8��Y�/&o�>�)��>t��X ^���\� �O��3a�̬�E��Gn{��[�1\)���B�RkOitn#��Q��C��sf��@y�uX=��K�^����8��`���.;^�g>���&��f֎ì�l��gC��wP����zc<�N�ze�X��EeɅ�ki��w4�Y�~�iϽS�Ȟ�ï't��tV���?���`%^��߹�� .�Ag||=�	5�V��+�.}�Պ��9�=���ۈ��ye{��Zo\���`p��g�~K(�������Yѩm�3�wò=��"��+E���O�a�3��L>��u���;��מQ+o}�f�����F�������:���z�+��C�{����g��=E����UBk�z_]9^�dע����p(�Ic��~ӑ�⺽Q�T��~��V|�����깼2"[�ˬ՛�w��8����������sB�����>�~/�{'�o�Uj�}�b�@�����)B�uaӅ-�%�D�@>��2��s�X�P�j�q�Z:25ǫ��ɰ�:��xϦj�,��{�/���-�r5�;OW@80����� �Vݹ�U�̛�2���8��"4�_F~e��=�k�WB�j���U�3Ǯ�l�c*:���Κ�w%;|:����eY��?;�X�d)o:+ncy��;Ç4�WV��VR�ۙK8�"�@�3ﺳn@yS���)ٸ>t���E���^sXP�V�8��G��fl%N�G���T��G��i����O���=�n=�����d�W�a��x}
Vfo0��"��ݹq7���B��z�9����~�#_�܁q�7���@�qJhyV��KӋ&{���b�Pg=Z@�9���0��Mg���{H�ՠq�DK��Dw���a��Iܴc��}
��9q/ymI�X^��[+N��� ;:��G���w�A��>�]�����2��o�5�}��;�%��D{��^=�7Lm�=_\�2+�s�=�e���b�۟m�\{��
�1�l�?	��/X���<��\�F�nZ+'*�en�q���k\�3Q�Ǫ9U��=N{%Zښ��q����o:���ho�<��@*�Ǫ|�d�G��+tøO@g�1��͡)�]�^KX�����<�b����/핥�/z�H�bP����L�:va�߳�P��+{J`G[�Ff�r��	�K>�y���`	�V��/V���%�n���V�����>�3L��ă�E�Nf��{�r=�!G�Ę豜~����{��}]�{)"��Ȁ8��M��v>/E�s�Q]�����"�0���q1ӷ2.t��_TMwm;w11�|��Ҵ��,K�^�j�|D�Ve<�: �Ӕ�뫮DB�S*��]��s���.P��@���t�:����7�k���Z�`5�Ż��F���7���oU�e�H�ϱp�-�D9��
L��F���B�q��k�z�^گz���m�gQՔ��8$5�=h��t�Ij�<���#)K	�Ҕ7& ��?�wq7�5b&����M$���,�r�P���o�z�H�3��u.�u��T�
��'u2]�ݘ!Z�p�;n�J����r�(֦����3�TB�`���՜��i�V�ड़R����1��-��7;W�K�- f�gC3� �$��}E��RY�[�DQ!�;)�]gU�N�	�sﶵEmb܂W^_q����g3�t��H$�U����!u����c�[��z��i&�O�Y5p �n����k9��פ�U ���
i�G����7
4�����<S@*ЪUf�6�n�s��� �L��Gm�s�t_Z���6S�5h��G]���C�$Bb�+���:�|fst�BLf��m�A-�3q��ԭ�a�,0���w��E�wb�˛�yo&q7V,��������p�O^�����َ. �
l�F�Q���hs�8iRy݊�;B>��ӊ����ʋ��W��Ϋ@��}�p51����K}B>�a�!X�Y��{[Uf�v\B������:�@�]��@�{�M˕�r��u��"�^��qr�.�З �)�6v��{����ǳGM1�)vJE<|M�]e�Y�]Ձ�[Z���W:k�֛E�w�>���&r��l=�tP|�]�6z*�y��M����xn�᠝�+���AEU��WR�@�N��̊��΁U�]��*�\�wF�b�-Z̾��7��X0ghK�-�p}���dͣ�V�����j����Nût݆���3���w��:_5��G̳�m��WrMQi�9pQ�+�^�Z��z ����W"�:����H�	����m�q���mf�cr�'�qb�hf�����Uk��e]e<��f�	Azr�k%�����֝ԭ��_WV�t��)g:��(�ٰ�/U�ZހZ}ݕ���|Ùl��/�c�����v[�Τ�i 6^�g;Bδ����<���[�4��[5}��L�W�6�F�̳����"��\�����#�O��1YQ�\��Mز��6���A��a���,�xDN�V�r��/����ng*��+1K�����*t���Z�^�GC�k���8�����)�q�XKl�Z��Uf0�U��J�R,��V(���F�c P�@3�YTc$U�J�EB� �1HcU�Ab�[h(��c%E�PX�(ʅ`,X��QZZ����"�"Ȉ�cX��AH(#XUH)����A`�E�R�E��P̪"AH��"AH�PIY+ U����HV,���	P* �4�V��
�V*�@c$Y
�Z�dR�BV
�,Jʘ�P�Vc
�Z�d*�"EF*�kX,��(�,̠b9IDaU�0��AaXT���l1%I3%p���Apd�Kk"�PD
�QIQn<�Gr<w�4�C|�	b���Ⱥ敘���o�$et4�6��0��s�Y�Ӝ�5R��(p݇�iV&��ʌ�*��I`O��\+�%���>��7��6���k������ͦ�:�|�)׹I��蓮���tK�f��p�2�kO�#&w��Bsq�G�㟳��{i����=��J_��k{��S�(*�(�QJ�лl�߶t��K��VEU�7=����:��ϑy�L�Q�|υ�� ��̩�U�3*�ox��$w����q�c���ʏ�+�t]��&�su\�O"_�3q�,/=86�z<'/�۹��ѯj<=�l�z=��N�K��YH1�p;�ϟ���˖쉨�M�A��-���^��Զ�p轢׺��Qi���'I�q>��dh�z�~ee�/c�CsP}(zz1C�;�UV=δ�r��	;>�����p�^(��h�t��~��}�HG������C�Ϩ���V�z.;���\`����������S"`�\\��W�P�'��x�7ģo�Y{	�Z�M����hI^ z�l�*ٳ�ٔNE9�Ҵ�|�ԇ���W��C�:k8<%�g���طV��R��K��?fA�y5� Z�-ɺ���W����h���û�����{�&|֝�ҏ�`�]{H�ʠ�tq��Ǝ7?9�{EW`��������y��%W�߁V�~��Ս� �tW���V1��s���bKN�,:���Y���f�^F���s�l�u��]s�̦�@��!�lUi���AN�x��z	_f��XCՊ��t�+m�z�(�Ӿ�xz5*�p���)"��u���UW�웨{��aߧd��t�ձ{���P��fJuIMG�M׾�V��b�.>j�|n=�@yauC<C�z	�j=U� ͏i��"�;M�C�.77��wѾ���o�>�f���5�e�cUS�/�� x�{�����IG0K8��]����-��l�}<2�ա��;[7���3q%��^��39���:z7۷]@�BW\Ϧ���Yͥ
j12ϖ�'�J��lN�q�ZU�O�i��#}<�-y�W����1>�>�>���u��fa�g�o�*��s�.�]�"'�0�Ϫ��3������r�������w��=\��}`o�^G�p/z�Bw����)��>��VET{}���u�}�⏞tSj|�^.�Yg�#W�HC������:�=����u������PW�����s�9ɨ�vK��h�Ve�U��?�3���G�8K�sʇp:����'�u��������NQe���>�E����T��c�@�@�>�`Su>�I�϶h4{�0��]$u��TG�_�Vz�<_��pS}m]�a��It��q����N�sq��؇0L�ЂN�Û��ц�kq���cϧGo?J�S�w�[1Ɋ�(�l��ybl� �ŖC³�p�aU׌ʝ��΅�q��C���j醎�7��Wr��;e�݀!2��Ѹ���>继����F^�KR�d�,��:s������ �d�ϥ��G�6XU�|��c�kx����o��hW�G7�����>�+�\��1-���U!T��XC+��ς����wډ�^>�rgR��%�S��ǚ�e�G�H�y��"��9�Y�|��(=��LLS������핚i���/F�j{f}�}��1�-U�||
�z����%�������	�������^n��W�7��>�<�v@�xy1>ʯ���ϋ� +�����_���U�}p\<%��^����z�[d���I��i��P�!��9��� �ne�_����{P�a=
�iyI��\֏qț��ͭ�����X�3ZX�r��y�T�b��8����<����W��1}�9qZ��}e7��?�=S�ǲz�ø}g���?���%~���y�uͧ&7�sy�77����t��B_I��	�>�����<��qc4�� o��
�-���ʰ�{jo��֐=��ޝ����ݢ�y����>��T�;;�V�5}@~��Y<S�CĠ��!6�:а�8���"�t/'�+�e��J6c$�vԙ:V�7�۹#%�u�Vq�s7,F�����t��-�or���s@v;���+�g+�R�U��/��;�C�xm�_2"� �"mks���:�h<�7 k��A���@Rs~>������S�C�Ǟ���n�co��!�K�Omg�4拓�ܫ`U�d?|��:�gT�ap72��?_��_��\w��w�<��(�A��zj�ʿmJ�ޔ������^}U`M�w�)�a>^��9��)w�;��{�{%��f��b�6s����W�U�VQW�X�J��W1SȊ��"�����W���-��ء��uԌn�",�t��ݟ.�qs~��@YR�vk�vG�����E��2��J�u�L/f\���گ���7(�X|�o'lw�%��Ӻk�z�q�g���!�_�=����^�f�V�1�6�s8�v�W
��M�*�*��>/ԑ����/>�Y+����?W�����7���k}����~sY����yA�Du<8KGv{ǗuC�}~���R����dF�`��N��x��ѣe�c��^3>4lz_y�����8�=��
�_���~>��D����e�|�2}��GJ+��^ ��IuD4w>�����ZdV��ρc+��^�g�ܭ��J������r�r9��a:r����+�Y4��6�H�E>{��'v��I5#���֡�R��j����k�j>M�f�v\~۽���-�k��n�v	ǥ�ÁͲf��T�����.�n>3�7���{&_:�)Ź���Yam-��JV�Zi���᧻�Ж���.����5>��C��V���K���z��QTz&���}9P��+t�>'�g%�h����O#�X8�8�ˉ�m��PwR5���i�D�A���z���DOT{�2�L<����{2��>;A����Y���gѵ�	����T���S���U	��
B��D�9s����</=މ��Y^����n��p�@��g�[U�Bgg���/�aW�<G�>��{�v{�܂+v%O�&tK�����D���r�z2Z����7�|}j;]�Q�o�Vǽq�ߞ+���dvǷ��G��Bڢ��̒�D��eSQ�Z]��;��\��͎~�{U��o���_��=��:��R�p׹�X���E��/'�V��x�q3��>E�鐓��R��7E�����QU��c�kt���W�۫W��s��,�s��Ϫ�	��@��JdA����}>Գl�!g��h�q��^�@�9o��9�B�����ǲ=#�5\�ɨ�g�m,��ǤҊ�.��x�̪ɇ��_����"���=��4T{���Ȃ�����Cs[�f7Vd�����s
cNv{�]�2�#��Uٱ0����S:�4�)6��:�* ��5<��k͏P�-����n�D����}��m�ѤN�����@5���{���'���S�T[���֓�Ef�k�!v�R��cE,f�Q�p��FE�郱��}�Pѫ�w�����Σ�������C�z�:�v��P� ��7H�}
����@g�}����l���_W�TNq(��3�Oo�ΰ'��>(���e�S�DlU"f)�x�Ϗ�i�����C�l��Wm�c�Z~T�� �����G�t~W}쫪 _Al���u�+���U�u�ۼJc+���}j�,o�#~�������������ND��=c�p	�^��Uyɺ��;�Qw(���{ݫ��{�'�{������6���{���T3�e_C�(��W���p��.${t��@V�{kf|�3�Q�ͯq���&kj�|�e�cUS�/}L7��U��Q��<1���x�-��^�&<h�F��'K��G�2v�oK��������ܪY��^5���o�qy�}���:o�����NJvX�ɭ*���7�o���6�k��Z����{qLe��SQ�����
��>��U�o���ty��>��VU1�����}ig�+<��k����Tc�vo	B>z�_U�ޛ]��"��N��_Z���c�Ղ�-��&g\3�.S7��Ȝ��άtU�Zy�LߐhvޫC���p9��qr9���<}�[e�U��:FL�ʣ����VM�b��;�T�����us ��`4�J
μ���Z��=Φ��C��' �
|}�}�\5�w����)��O�t��UÊ��ם1�P���u��<�nc#���p7�w?W��s�#�~��YhhϽ���}Lܹ�ܹO�����ç#rP��%���z2g�x�<�v9״��W�[=�8[�LZ���V���H���ͺ�=��R<+�]����.�Ey�
��'/6h4n+�� 9H�9=�O���Z���F�c#{��	V�W�QG�d{��$S�L
��<��#e�Wա��l��19������Η��������騿_�Dez���y�RL����>
z6K�%zz�+}~��3=c=�2�G�����t���\Q�sp����`���1?S���Y��3΍�`m����U�G7�tuz{���K�p���=��� ���
�4x���Zj`�������z��7���v@�xj3���d/:�>t��R *~��z�����������'�1�͆6�h��U�t{O����	��z���΀�9.��Ys�f������E�5ل��a�e-��+�kGe�5��J�2+�ϮFqjlfe�c\���R�5mր��
�J�O"wڮ�.���8�i��>E��M]w`��ݘxvn�U�IPI�;���@q�V˛�n�Ҩ����]�O�i��O�J���u���Dic��2Cn�0��
F^f@�>n��;�5��gНW
���ٯ�zC/O�?�uOW��w�2tV��s���Ύ�"�4.��k��ˁJ�;����9S~��e1ހw	�q��<���qc4��jW4+�1�}����5�x�Up�d�������{/ÆG��|2!��s�Rʨxw�Qs�R�s}<j��
�CY.���H뎩y���N��5���\y��;�i�{R�Oj^��
7nT��q[��'�qS�<2��p�&w�x}3}2��s�_����Q��'�yૣҶvU6�VN�!=ah^MX�h0W}U�M����)�\dϗ�9�|]{O�_�q����
����N�;�TZT`Y٭��7�>+� K%�k��&��|�Jj�����O'��˽>�6=���Gc�>�q�Q�
��{�tj� ���-�-��,�������6��^ϓ[�g�/�f֎�y�މ\{#�Do�^���f�!��<کo�	���c4���=$Lҭ�L��zİ���u��Z����Ew���ݦ��Q����Œ��N˻�c����)]1+��?��SdNvO���7
�,��P�ޱiSB��4Q����gJ�G��ݝ ��Ȑ�پH��gVc;���K�;@�S�YJg���	�Vf�y\�:_�#����{��8\g�ף#��P�	����ٰ���};�2��>R�ElУ�O�qa���a�K���������g��Nb�0b�S����o���TG�͢�����5DM9�;�����ǳʫ��ų�3�'��ث��B�������]��.h�@�;�M���=Ea��\�`,er�p�}�+�B���E�����]�L{��C�O���tB�ר�9����n���O��J��j.�<�K?:� \�G��Z�`�vՓ�p��=��y�=5sA��w����>.��\FV�Y��ʓ�
�G�E�/�J�O���0gѴ�	[������rz�ު+�!q��.}AT�K�+X�U*����{�z3j��i~=7L1j݀��<B���G�s#~����v���Y�yY�U�.?b
�=X��*:��g��.j�2�V3-�f��1of2��Y]��|���n+ѽ�>7�Dw�~ǀ���o�O��ig�S<�yM(~���g����~�����c6s'եR�c��+�K�O�����P��YLn�K)b]H��R�R�u�Nƻ{��"<��H�pW�z��I�b�v��
���Rw0r���yv�c�fn�o\��+s%1*{5$5T���Z�;%��V�kP��u�m�/$ٱ!����q|_Oq�������{:Kg"^ւ�����,oѓ:���>E��i�8��=��n� ��⇼���{)�Z����۟^�eD��\�U�5<�`^���������3�iO٣�T�w�������w�O��?W�9�A�S��vC�Y�.X�MĆH�9��BM�ٔ^ϑu�Pѯ�=�>E�g6v�;��&���ʔ}����G�k'0t(B�ܟA���(Ⱥ��������4j�����sސ�3��::j�}5ďz��sc��)Yc�=��}cd�3p`�;u2'�.}��Ng�/Ư��������D����q����99���+�߮���uN��xO�o��T��s�:2�i������X��ܯ'.<��}c�*�������
�����<��-P��d�Cܟ�m�)��Z��͔o�<�����^
�ۏ��d�\?Mx��X�����=��x�}U^Ed�C܏fQu��7bf�ս��H�z�I�+K����Q��1qUO���:�>.�g��|�Q��#H�.�E��kk�s *�0��[�XZfL�W��Y[�ٮZF]:3��]X�S��2����������P�d{�%��uwz��x.�񥱻�s7��\�.!��ﻩU�5����/ub��+I��
�U����zM徚��n�Q�)�ذ�dK�sz��KVb�o`x��-*j��F��a��A���������sVM	:� ��gm�v�v�A`��ci�����,h��[\��jĤ�ܫW�C��U>�-��F��]�%���KA�#�-BWB�Gke$f�Wܶ
��`}��R�Ջ����i�((�u���u( f�Bm)SH�ba�Ѥ.촓��dRM�d�DZr���-���C1�����58��X����]P�u�G2�pEf!�I�S��i�̎�f+wWb}��څ1�)��*�� 9���Kl���L:�ӷaҚ׬S���M�U�k���u�������6˧��yu]ύ�AK][�V/����l4:��؆��`���V�v'hK�ՄU�B��xv���׳O.���L�`��KQO r黴�A4�6k��,:��Yٽtm%�+�El���WRV�KF���u�+�tuuˠ0X�ćp�h��`�Fk[��7$��P���ٶ��!��s��(�����	4br�RU��\5kC���ۮȒե���|����Ʋu��ڧ�T˔{�k�`�
��X]>�d����G��2��$mfjUS3tC8�h޾�Ѫ�����E�eu�{����qb��s�����ȟV��F��UJ�%ɗ[Jm��@}ƍ�WҢ<6��W}j�^Cϯ{�s�u>�S��m�h|;��Y<ԺX�iY�1�H5ē����Cb��wZt��iϻICԯ��^K҆ݰ'1Ba	��]h�_'�N�Zk,v'�#W�����
��7 pX�Lm!/�������mw@�u�W\)�1t̺c@9Ʀ�����X�m�&����.�*�t�ŵ�}�C,c�.q�����P������L`�/���Nԗ�q�9�+5۬"\�>a�.�nS�w�m�a"َ�I����l�����Ve�ӡ��gw-��\Z��ا������Չ�sxv�Qa7�h��n hفu4��ۺ�E�>f"�K���y��s`��jKH�Ю(;�7��=;n���Ƣbc�^!��k�����#��l�
"E�_}-���QH���v	�\��ņ��ʇ_[�f_wW:�f���5MZ�tV���&h��WD�c��$J��/���R�찐߂�_�l!� �J��\������Wt�@fy�.�7(�*q��*���E͊�H�3��[�.�$r����!��K����ݑ/���o!����9�o9�%�s�� ��;j�H�ˢ$Ʀp��)�R��[�G*���^\��ǡ�h�)��]�ܳ̄zr}0^4�D{C�:Io!���ߗh���#����d�k����*ҧRx`��`2�;kx�@b+�H�*���(c%HVLf2�+s2��Bf-���DU�-�	U�Y
8�ĮF�(���%�ԋ
�U�	Ym.`VbTPPYX(��eAd�d.Uĕ�0�#m�b�Z��"�#lC�Ub�[#��8ե
�`V�J�!��+V���IZ��*����V�¸��LLJ�QX�Z��PZ�Ȱ�1��Dae�I����jF�+�(
�-��ˈ��.#��b��X�Q
�B,��G\�`��-B��(��r�E�R���h���JPF*�iE#l.\`�8���m�b�r�`� �b�Ykj-aRօ��\���f1LLT��FE
�2V*���q�*"�lZ�
�G�~��k�������� g[�juv��w��sҧkk2���^ R�Sw�ѻ�o�hް�T�je,q�F*W�[��X*J�z������7j:�6��/��ڇ�V��xo��O�҆3�޻�lDޚ[�J0�V�9�g2m1�|w"g�s������鿴�,	���bs]����>�1Wn���_�������Q)�>nI��}؝�2�&����7��鿸�6�O����{�4�$��8���P=�I��:���c>z'��e.��2�kK3�)�am�x���{�Ӗ�e��bp� ��7=�`J}�����y\7^T�=�M����=��H��Mk�l��U���J�m��y}�('��!�������:�=�_�`s�S;�J
��}bԮ~Q]����/w\�B�@4O�� ��+���z2e����9��J�ko����b�Ş�o�{x����C���^�����6�7p*���϶h4yyTJ�t�����\f��s>Qrwzv��׹��ϓ�YC>��~/A�<��*�]D�`W�,yf�
�/�C�WS�����܏`�ApWUH���1��>�I�~�P���Qc6b[6`���*�*�^+Ar�s5�`��w;QK��蘪Y��p�²�NiI��S%�+z�k����2��w�VAOc[%�"��Kg��n��b��|: LMi�]s�P�+�ĭ���� C�I�P]\��U�p�N<t`KB����>�`'����ɬ�9��:�O�g�����/�Qs{d���p`l<f�X�3<��H�y�2K��Ʒ`�WLlN��i��	aҞ��K�C��)}�^��=�W�+�p.Qjz�����/�;3�=���g�O}�bb�Vѽ)��0��/
�~U~8}����3�Q�+ ��[K���Ua�\)�R�H����̈́6���!���N���{��Q��C���͛���q����)�sR�ټ�����c=m��~��>w�;Mҋ������Ux��X�3��lr��om�vE�*�y�=���T��ꉝ>��z�Y���C/NG��}�� ��)c�`�?g���i�O�j�̛�h]�!��Nz�_�����}�ڱO�Goz����v�j\e{��WT(6/b�sn����Y�r��`O֪�㗶�ztoG�o��V��=�s��:�G�O>z����y��V���Uꇎz�F�@�q�#�lv�s���Q�����1�墐u���s�[5�=�S�<T���G�خ�ד;�>����e������o��J��{1���Wq�%oWvF��XZ�<������O{)Fcg�ї�m
��X�ӳ5tz���O�(�@g��v`NC*fu[��J�:@�9�E�uݝi�����xG.��3�.K%���KN̫���P��y�.��9�˺Q֚R>��]�AS�;�FraG݀lR�!ےY��X+"�����p�&S���g�Ӝ惽�w�3n�ı�}i�M��Ż=���´�>�R�ˈknY~�Y_Kt�������E\�.2eTe�(�?�
�˔�W�w�;�i�Ό�G���?O��:�\z̳�❛>t슩Kd����>����ԧrp年W��a���:b�}B��?I��~�����{��=LȜ�jI�����:���8KE��5S�Xr�I���/>�u�����E��zn�� �yg������y�ˉn1>3r 2}�tШ/���%���&�G$�|�_���G�X P{ݚ#��Ǯ�wL�����Ҿ�����J��s�w �p��/	�t?+�Ev�t�ә��^�X./�'��@;~��]z��UD4xԱ���=Qr�ȭ{^���n7e�ܚqѭM��84��}�;s����ˁ���ù��F���"��<�����t��g��{1���,�<���>��O�d�s��~tO����,�+�V�O�쉛_��,�~�W`=��ג��EG-ҡM�t��G�V'K�taB�!v�d:emA/��I�Ba�]�:�k�
�����1v���ؐ��{2d�E+�0�v�2�L���q4�f�ӻ&a�2�GW:\��橩u,����9�.T�c ��Υ����hđ��^�{]���3��	_�����
=���2�	B��*x�-b��[��g��ES��g����q����Zn4�Ǧ��m[�/�[�<����̪�i�V�~�;�[a��(D��=�j|x���Ӳ�_�[p�2|�oK}7S�s�&):�W��Qk;�{`]�[��W�L��;�Okx����ʴ�LeFMiw�;��\���K�2��R���U����d������l��Oq���w�[e{:Kg>������~��0�dW�g��w�n�+��z�����$?oMy��9��e{��ի��~��
��.��6���� �����9��븭�������7�('�u<,_K����	�����u�����~��
��ûl���N��}`_����@TZ�˭�h���;�]$s[���գE{��🶫F�1��me�ӓT�����q��7��9FE��ݠo얏�#j5}����9�HG��ȣ��|�o��ܯZp�d�Cж��\7T��CeA�����D�>����26_�E�T:��N\�xz�>~�7�0	6�ڑԢoi�� ��Z0��Z!a��#��sѓ`JQ��z��O����oh{|�+�Ws�w�����$[�ɝχt°�'r��5�̌��-�;X9M���NM����"(�ܒ���*��i��o��f�&���.9|�T����fAS��s��Of�`��N��|͘(=��D�S��џJӵ&�k���!�s{u��|�l�{���ԇ~��L_��^��O� W�fA��y^�Gʄ�t��͈��0z��J��+��w�M<7�Gѽ(wd@�2��Y>	����t�K��=w R��m�U�z�3r���\�{l��TV:��F?|�tÿ���kO����|�[�O�ǔ��YuC<r
� ��Mk̙�>���c�lЏ/�:��6=��3v�כ^�q��3�Ż��mUO����0x����¿K]��;��+|���(ٿz$��d��~��c.=8���Ǻf�~Ź�=��܆�1�w�e�MW�59�>Օ��p{M�O�P��v��ɭ*���7�F�_�3���ެ�]�f�9��^ٛ����{�u���/ӼW����G�y����}#��c*2kKR��U쩡��|�\���|ԁ���=� �\��}�낿��=����
l����%GTys�������ۑ�,�T��dΣd�	�T�:㟯�s�s�#�~��Yhh���R����;1�7�Y�STVh�aL^ʟ>s��7G�tpDy3'[�3:�egn�.�{��k�:+h����_Ae��.��yc��/8vI�B��ԥ���!Φ����@��l��W�3{3{��&j���4i�,�b^�����!��F��ˆ���Ը/�\��s�ޜ���T=��)��&X^9	=���^���+r�lpU��7�)����T�(R�B���� �.��Ei��Q~���!��;�P����S�Wݤx��+/<x}�>�:�_�AYR��@l��@>Ϫ�]}.���G�X]E�
;��Y[�������xƩ�|��x�3�g�=�%�����`������&W���I�L�?Ur��{��\,��Ҵ��}}\�.���~�E�}�#���̂K��ȿ��ڿu��[Y9.�n�Ͷ����,���r��|���\��g ���/G� w�pD�e�����}mb�x��A	��5��11O�hޟx�A�g~��^���r ���.� �Nl�=�Q�On��w��pD� }ج�Q.�[�lxm���ղj4�>�q�/���T�9/�y��O=�D��}>�އ��@T>�K�5>	�����6�;�����ɭ,{(W���mC�Law�
�3�d�]���STL���U���M߈ea�x�D�~q�Z=,w�zl�ᘔ>�د��v\SN�[+�(�K)�5������a7�ޅ����0j�ۑ�w"WM�܇Z mf�I������ދ���y^���]�{���mp��h��
l��k!��b4U:vLZ����]n�����ll}��,�A�P_>��Y�mhM��s���R���V*���:b��
\H�sbv��^�s�y���pЏ���kM�k�5�u0&-U���߀��p�vW�n	��wKu �UϦEHg��=��~�$�[�ߖ���l ��@�}R<6���������N��;6�
^��}{[o��s��D#��2��"UhҦC����d��o�>����6㟯�r#�/�s�ڝ����7����"�XP=ϡ-W�"�(�}B���X*f�Ⱦ���S��R��sA�ci�Y�I�ohq|����}�2��{h��Lf��YY�)��[�dUXy�>E�S�F�O�ٳ3����f�^�~���������}����ע
��uƸ~�~��i�&�����Jɟ�R��HY+��mx*��Z<���ǽ�Fw�~���+=7#L����^���v��ރ8޸'�T�=�< y^L>v�"�K�6s�9@���*/֮F�۱���v�o@��S>��RW����n)M
/��p���~<���K�����X�9�9u�C/���n��uCD<,��I���œ�������D����·(<��k����/uZn`f��)�T�����V�w.��IF(*����;���ާ���m@j�r�t�ZEd�Ԟ�N�������tOok��R/�S�����nY*�i��b����j����i܀_��ٴ�*=v�s��J9�й��v��#k��S�̟"�~��O��uD4{>��6��G�.V��wǣ��?e��(�^�s��ݶ*:������{·����R^�I�*"�|�g�urw�>I�v1����F�M�=zj��&Nq�g�mpU��b���{##��r�~�WՐGzVs�>G�ݚ5" 7�f����D�9�V�y���<��L1	_����q�'��#c�!s�G�(�G�<����q�=F<l��3�&�F.�y�8w�/Ǧ�������9�.<��R;�����]��>�Z�V�dʿX�ݭ��x�r����\em¿�Ԭ�i`o���gc�*n{���V;�����;��rv������+�F�=Wq�۞7��O�p2Ŭ�����L\k���/-�7�,�z��O�-��@�ʟ�q�:�y�^G��E=�D�NuW7=�Ƕ�i�R�b2�v�r��{�Ϝ�x����-���^G�=��6����������ES7���'�C����P]Ca̻�g�YAV-��Mew5�]�����4�>�O��J.�06�����I�`�R5��%�.��U(Z`��V�V:��+��
\�3g��6Ur=�ˮs�^9�Xa�x��l��-���S������i	}��;���=N���wP�M�2,���ZNmaQ{k�*�<��9x@���7�>�O/ף܌��?����*�b�^����A]!}�������ݨ1=
�7g�>,���1^tZ���6��Q~چ����\O�w����n;D׹{�{w2����u��+���Ҩ��2<���P��2.��@�h��Pѫ�w/֑Ȭbvj�~Ɏ����Q>^B^5���_�Fzg�]�2Hlق����D�s�>���26_�{���i�A�ײ�M�ODVO�==֙���%�p����S��	�"%QN{�G+˩����{ǔU:Ӟ�teF��c��ʯL\A���`/z��MU=��뉺�ւ3U��Xr)�cS~�G�Lz!���z�q�|3��,'�||�{�%����+�����&x�R�Ǘ�{p�DM�=���0�t��>�����Q��14���<�+����r;�gkJ��>��2��`��c�>���a�0i7��T���_�)�?�����j�|F����0z�U�<}��$��et���g���z����e��NW9]7_�I���� �@O��C�˸���Ǵ�	R�U+����lډ��]���E^DUkF��kop�Ẳ���r.�=A����Ѣ���x��"�o�+�IT���MǥR����%Q�t���ǚ���7��wώ��r�@Tx���%I4�wd���(�ȝ�q=Ú/�y+D�S�:k���:�+ە^����O���;Le�UhW��ZI���>hS����SZG�S�G�ڏk�j��x����-Wq��<b��Wqȉ�:���y����ʥ����`P^�C�e��o���H��v� T,U�>��p��}��;}��Ž�M�L>(��w�c����v�>\J������3�7�L�'ʤ1��~Ӭ����:�e����p3skg���O\��}B�7>��}5�]�xee���㋯i����_<W���
�|�Wn�;P�z��ζ3�9Gǳ�z��p]0L�)��g��[47��YH��tH����:6|�7�G��;�#��iջ��=�(�4��>t숪�u.�X�>��[��/d���]S������mh��=�[f3��*�}��S�T�>�IcLȁ���o��i��z���nTO��q���f�
�x>��x����ϧ΍^��7�Nn;��{�y�}�F���[���o��6L8��KNA-�0��t�r��
���������}DD}�}��@ @?�I�RI���!$�H����@�$�����d�!	'��H���@�$��$�I?���� B�}$�I,�!$�I BO�BI� B�PBO�BI� B�I$BI�!$���e5�mnO�BE�!�?���}����W�7�����B�A"�J������*�	R@K糑R)*R��UT)IEE[d���� ��:P�JQJJ��%T($�E!EQJ-�B^� �:���*ֶaE�0!kj��5"�� �ʢ���V��T���gB�S���T�8�Q{[Z�4��5m� ��T��2l�����bT�63f՚�)T�[*ZT��� �qCn��[��$�;tձ��4n�B�2�n�r��tʠ"����pkV��t,:�n�v��˲�n��*�v�.ËGe�,t%���ۮ��R$������kj��uӭ��6��5Ѣܺ�g]j���+�������j$9�P��.�j3fE��hU�QQ��!��B"
DةP�n�%�̂��J��R�Bd�m*�֫K%*U@\ .%93Yf�Ѣ�
Q[kf�kZASY�Uc@�����S�M�D(U)��M��6�E��y�    0dʔ��M 4i��d��$�JP�0 &`	��0	����L&i��S�A)T�       "PBh�&SL�5'�����a46�R	OI �$Q�104!��&�dɄaקN����+lz����/]�lVj�� ���U���h#`@�PA���Pj,�O��?�?���k������  4�@"5H�# ���8����q{�g����n̊  �_��	�1��H�P���f�!&��ߓ�I�1�Z����r��g�5&�+5��.k;(b��[��]��DB�ְPY���&�L.�[YP�h�c�S�:�륗��`��vn[�SS�ʵIīZڔ2��&���EKP�O&j[A�Z/*�
��ABvf��fa4���y����,�Ҋ�ӧzp��`
��{r�9�mX{�i�U. `�*6��8��6�[�{��I,Q�4�3{�)��*ɉ��
\S���uz��B-YJ�Ph�R���t�ț��^��--@aJ�ˢqD(2Q��3qF�R4��^�N�E,	�7]ݦXU�7���ib-��"*������h�E��Ӯ�k[�o��3r�hhr[��f�Λ5�%#K��z�7v�)���Y�@��e�VM���4�q	���z�hb@�$��*e�Z-�[�f��7����2�b�b۽���d)�Mi��:ºz�͚R�f�/-��(/kd�G�Ͷ��,�é�ͬV�T^Ƕ
���FJ�u�BQCfU�(|�Λp+�ι<5��l��IM�t5�.�K��"1�i&��̄�śn���l���,5����{�BLYw�B��#�e�m�[�G.������'�\aA.Y�hoc�Fm:�ģ�6ہ�*I������Ե��"Y�r<(щERzm�I,�X��kqL47d�,S�D�@NX�Z�!�I��W�ٵ�I�#5���2��-�;a�視Vm�lHn��T�`Z�F4�0ژH+M�X�n��x��J?R��P���&�h�i%����zPI�1�K��F7pb�X���]�MZ�ԔeVax��,B�%֪ñ���=�������]n&g��p��)%j"l�&�n�0=8)�l��Y�XH���RT�SA,h�DT���K�X��u�c�yK_Ѭ�Y��sR�fʼ�v�͛��SWBg�T�,:�$5�������.��2 ��9��^UԲ�/���X�o͖�W���L"�/"���ٮ�b�i�inڶ�
�Ȝ�H��a�Yn9x2QE��8��@��̓�Q���k)L����V:�cݎ&2���TW�X�RO��ÈS�A��yY��)�yx�jL`��m�Ʀԩ���-�aLd�j�B��`Z��FYa����&em(w^X4Ø��0J�1�E9��㺻�+#�+�6��)&�{i]@��ViY�helgX�y�I`�� �������VԬ����V,�VCҮ�$���V,4��(�����-�j�.��F�-���6���,T��s֘�#8����(TZ�⨾�͗򭹦H,PJ���h۽4�mإ�-"�%�2P��$�DTQ��Y�P;[�v@�2��c^b�d���%�.�hu�͔6 ,��w^^��R6�<4	�V4R�������I�R�YM��Wkb۵�|���ċ� � v����l����ނK�`�����[i��@�捥�6:ͱ��F�<;����A��
�7�6�GlSv�JH$*���t��5A�X�FV<�f�z�lڧ{i���P���mC��"Y��u.��Qm����ƣ�6�٬@��0�!,����S-�'�tV�Wp M�ʺ����!��h;J�"�zθIrB�
�Pn�Kqe�>ʭN���K��l8��4��Gr|���]^@
�{�Ѕ�[B9)���������VZ��ϖ�Su�q1TU�5ȋ���S�LиI*)�m۳r�ߝ93�[��-���Ki���)7/F�+pj� ��A��� �Qh!/	���!!lf�&��4.֋CX��)哘JaD)وY��PCo�!��S�6��%�&�xofVlJ\�V��;��d�4�=��Ek�w
��D�E/�i�+6�C� �:��N�;�֕��i���o^vG��f�n`U"��:I,cM�(-��jPͷ2=Lan���V) "Y0�Y��l���)�nւ�k5z6�A��I�v�O�7pfǙTP��u� u�yx����CH��Te����jD�p��f��i�S`W.93xN���\i�J㵂��&��H��f\6Y��V�Z��en��!.MeR	ŷB��`�mC����ѥF+����$�S�J�Ґ֌R\����PeZ1'wvͺ�U�i����Y��X[l�ƶ�:$��ǆ+��W��e鼦������"JTmX��w����k\����Snh�cP�j=̧�LO-�����`Vm��t�zt���Q�V�ڭJ{�P�mPV���@S��.R�&�8��W�[V2�݀��뻔�y)n-��_Cn�4���h�*X�v�"�T��Y��2�X�U*�u(|*���5�F���
�6�;�A��z�[q���R��q]�hQ����VF��
)��3�W��THY����a�4]�ݸ���΋�,R�)G�&eی��G�u1�iY�w�VᎲ|]i*�*�l(��ݫ�!�D���0�,OE��*�����蹳d[��@2��Oc�j@�䅇�/hH���Kf��GmԹd��Q�k��0p�'�Vs�0�W6��1�rk�ٸ#Cv��F���i9W�2�,K��OE0d�c2� f5�7e�"S��b�Qҭ��𱸆}+mC)"�R�/m�s`	b�tQ�R�ŋ�Sd�
�i��H�ś)����Ů��{Z�1Tf��J$:N�X�N�f�!��&�-@��"�Tbk�d5nJ��N��#A���C��֫��Up5h=��
�ili�1=P��U]ٔ4K1�a������oa�H����䘰h���ɬ��������{�^P��kE�cT�jUt�Y�Ir��n���}���������N&���W�T��ş�F	_�g��m~~��}���1�OS�SGT�I1�&��V�7@g�r�Ӗ��y�ݑ��v�-�[���d�����e�o��tR��qp���"�Mg-���r��|tC�����ծ[ٍI3`�-�ӓz�#�O�VjV�u��)]Џ��4��Ѯ����֤�U������mn����MTQpV�6��`S�i���)7�M֗r^L�E���Y�;��i|�m'ڥ+i};;�(����[ouћՔ����8��w[u������ﱾGU���:m���΢��.^��Y����ϳt7���{.�s�Fv��5}��],ۀ;!tc'9�����o�"���쾣3�8hM��Ѭ�v�S�v�x�UטO8S�&w����:gk\r��:{0ҷ�T�B;yU��-�c[.���&'�q��w�꼋��c��A��{������G�S�w���O�!�)�+����{���u��ٸ��X�̉G��g}��6��/K�s3��� u�(,�3���6�f���5"����a�Y:��m8i&��ڌ�ie��EV!�ݔ�O�R��\U�Xˣx� �&ͩ+�i��`7��V�*��C[��,���z��vIM:�܅U��c]���G3O���A빴�X�cN�`Ք��ޜ�X�ժ���EN5��f�e�����lC�D��i���Wg�,�<oU�	��E>����V�݇TP+y>�lE(Vc묊�L�&xv1���ȫ=`9Hu|�䀔q��r� ��IM쉴"�m�u���鬾�\�@PT�B��H��pP�5lJ�)�J�N떚���i�F�q���`e��W������V���[
j�jb���qr�er�0,�o,�'�$H+z!��-xg��LB�[�Ԝ9<M�oy�r+�,ɽW�M	�k9Rb��l�c�ẵN��ڌ�ˮ
S�c)pʵ"�b�9n��V�n��7FJX��"w��;��6.T픣�z��97{�݊��9����J���gXK[��7W�����Qu��;�؎���o���� 3n��A�4�[)	wP�{s�؃q39d����N�\�j�pE�+�j�F�f9�h�4�&p�I3v�L���F��=He饧F�&��D��t+N�N��.8]���9m{�f긻�R
����"�z�O9���6 ���� ����aN��Sh䢎%8ɜ����j��G��Mܔ�*:�f���BP�M��ѝl.H�^���8Ep����}Q?����t�Z9N�V���BZ��W3e��7z��-�p�a7�C�*�]�_e�k
�蠡"�Ʀ�v"��V��X
�s�*�t��ӭfn�Y�`!��`�j��s���u/#����ћ�����z�R#z�ͫ��1fS�v��%Ꮺ=Krp����Ne�]7pŚ 끊�m7�Р_}5P�ܯX`0F�L�oc��/��U�'E��e#�\/�|�(�]g�|��"�V��:n�u�G�Ӽp��`���T�i��[���l�mAK�3.+YՏ
�`k�k��;aY�u��N��[h>Y&����t����S����@.H[��vnͲ���}K��v9����uw5�8�9k^�ZZ�rq���Zvfm��%Mk)Wb�W�Y��ΎK���N�����r�r�[2���Eq���qS��ճi�̄VYuh�790���U�2(`�b�fՒ6���T�h51V�즻�i0�9z�1������h��Y�g���ثj2��:�t�_d�-ccG�_0��M�;iN��+���+VӐ,(`�����vѧ�����t6�MD�uk��>:5�f�5�*5�!W�������Yb��z2�]z�@!;ItЕ�H�%bn��;�sk�Tڱ\/P��"wt;��͹�(�f�Lr�5���lG�U>���G�u����;1�P7�qWX�F���]̃z�>!bםR^.�S	R�y�9�n�4&,��YxY��X�Tj���e��wu�4��!��|�	u|�x0���#>..4TW<������l�r�q0����Drά��["���^�Q��^�0]v݌).+����!Z�v \ӵ��F��>oB��	(�Z��b�rV��\.�dJ�dt��5�q1
���t.d+Fܖl�75Nސ�Ǘ�PY��@u4ee��ǀ��ڵ�Iy�TB��6\����B��V�P9��%�(�G�n��z����Vl"V歶��O�7�۱�Oى�A��Psd\��c7�K�����\*>����U#�k���`0nҡַ��1v�3&��]iJn���VS���I���J��s�VĬX�ᰩǓd����=r�Ό[��N[�<V�Ј��`�U�yCKrO�H¹I���sÓwR�L�<s(����]�;x����C�Zd�M�յ��3�7�um�w� �q.l�W������B�r���s:*�Su�c�F,�RԨ���i�Iک@Ж՗���+��ϥ�ȳ��������0�R@���/�����j��ηv�|�˶gp�1J�E4�f-�4��9��V4�B87nm�����^�t'y���5���1*u-K�*COb�ξAP{�3����w���^��B�8��zb�/L�J�ݬv�ۡ�)T.'HC�.�4�pi��h�I��չz�B��'wT�Jm���I$��IM��ޒy��gu6��I$��IM����$��RI)�қ}���I%7Ҭ[��T�y.���t�ô�*fw�_nvMM�t��R>��AY|�$��d�PH�A$�Q���Fʼ�2j�c������sS��u�𸡫�6gi����Ѣ��DH�vίjLkoN�.�σ�N��8r�
(3d��\\QQ�^���L�������>�:;��=[���b�-�դ�ľ�-��ų�j����t�=\�__H������vk��Vrct�ǡ�F��L&]lI�T�·�q���N���n�u�k(�e�m[�}ѽ�N�mv�b^��Z�'P��=���K_MrvH1MvuI���Ϲ���4�I�Ը�]������`\��]\	�4���l;�3x�����J(觬�tBs��8�P�qUZ��:򲑻�Z���YO�1ʤ�.��ڙd�SN���ֲ@�bbɑ����C�]�g,�v䌭��n%\!@���v��B�O
��PڭF��h����C{m���pl��=5���S���ZM�=�I��w���mJu����h4^�:1�O!1uqn�5��8>��x>[(!9Z�G�40)���������]
�N�݃rk�o��e���ͣ��Y�M%G��'�}v%J�>9q>6uSw{R#:��F�J�ݪ=�pwCg���)��oA���B�h<��_jً9�b����r[��F�A��fa��֒�H��DkΈa�.�b����o.2�^�b^�
]<1���I �)Rp�����{�6F��?s5���0Nu��I|͊��,�[�i6F�Ɩ�gV�A�q����)n��E�E5��� �i5)h�8p��CHb���)f�ꂙ��V�/[i�a�wE�"͕A�j
�����M9r��E�R�jb������{������J)ԝGɺ�j
XI���}����Ȧs��_5j�J��ʳ������B�Db�,�����Eg ��b�]c��O�E������t� D�:��E��v��IV�|oN���=��o5����؆����$�41I}�x���hCT8�8[U7`YjT8-�.��n�EHm-y�'�Qɣ	tY���wH�^���]�1%\�T�e��HH��4	���4�+)�\�J��:^�wur�]p����%t�9�P<k�Ruj�nMacǎ�t�_
TT�u�j��Ҙ�1�u����&�g&vV�����vAR�[z�M�t��"�E���^E�P�����W����W��%od�UÍ.��EiU�Yט1H�oһ:\1vFE���vs��i։��t
w�ҕ��)�ځ�K��R��X�&q]��
]�%}�vp�A;z`Ӷ�E�,dT���R�^uw���h�:c�u��E3���ᙳ:>m���[��`6�-׏���X��0[c�����#�CK;!�t�64�{׼��7���j�����X���Dc@L����쬁5e��63n��R��1�>3�U0�+L�X(�.����-�2GT�@�ʬ�vJ�f��tܢ�����"��-�����b�n$r��i�)m��q�sB̪Xgc�`�n�A[9ۄbSR���}2S��c��xΙy*g;paB��9�����_!�D[�Z���4ڛVK��2w����:�Kov�#��^V�)`��jr�y��ioE\;��q��/�h�����V�d$�ǂ��/*#-�۵u��]�[KV�d��eTdHgݠlR�A+�uʱ�A���4C+�p[�ѳX��(�f��!���Sn9���;�{Ǌ����ܲmFW`��L����>��*!��T�,>�9��k%'1n������ͭ�N�[t&\7r� ���2�Eq�Ξ�c�Ugv�+#pҧ���z���{�����u[��o&��j��[��"U���x믜f㇫y��]����'p�Nr������	Jo"��uJ\6�j�-c,�b�Ө�X4s.�d��2�,�+5�Ǳ�H\�w�E����)��WW�:	����Y(ǔ�ݓm��'[���+�_P	��v�D7�rV�x��m�eB�]HOb�x��
���l(3� �9�ιm�C(s�d�x_��:��f�g�j띅���W>.
�CrQG�v\��G���u��Q�M^S݋�
�yWdqH|����I�vSHQԨ����w^	�:��N���3D��=u�j|_g7kk9�S<��S�.li����O3�9�*^+˚��^��k��I���p���L��KDn���cz�=#�CS?p���$��t!!�"^�b�����3n���dj��[J�]���B�t�m��.�ҩ�V䲳��V�g(0�b�<f�;�ҧ�rJy�#�	���޲z�>O��2�r\�]���7��fgVP}�'��P��KN=ݢ����oI;C�'R�S��襌���ŊT�9�w�������D��\X��T�*�Abmu!oY�{�tu�r����c[{��Cn�֬sM�1R+X� X�;K�Ci�փ��{��8U��������R�)n��O.�[L;����)��(�2�eXI�u��ƍt�U�t��\��\$�nc�P��%\�fK�p��MM8�.�E묏t�����.-�<����Il�y����Q�����6�0�3ۅ���J3g@�r�C�4ct�V���|fS�`gn"��#Pi�j��Ķit	wjU�H}X���;Iު�y�8FrU�Z��E�R���ڛ6% �pH���"��� �p�*7���הRtxP%���h�'�Yٯ�c��T���쾢����|B��Y��ѱ�1�B���P�}@�Y�}���˺|�ͭ�t��u�f������_7L'-�i�bC�U���`����3%.���_TZQ5zC4ji{PFڗ��u�c���R"��cQ��Gs���އ��hc�bwZIt�9��˫D9wς�Q����@��t�&�ꈛ�}uuܒ}��M�z:oG���[����sYXW@��A:��vh
d"�Œ�I��a�|x]s�dO뗴�Ʀ/�Z򷜇�"H�|��ա֥ѭ�h'o���>��W	�~9�C7Ji5"2��U� 5�dSf���Ӳ&Vs��a�䗫������x�f� #�M R@Eu��1V�
6;�؅��n�\��qҐ;�V'Z��,���*ȇ.���lۤ���H"Q�B�xU�ɘ.ڰ������=7A'�ompyP��]��we.��gq"�y@��b�����������l�Z�ͳ�������; {����P:���5�����VX������H���G�,BL�x��L�:�Y�m4��*}C/�Ċ6uv�f��̹XZ-�N�EJ�r�p#׻V-+�}q�蔊Q(�9m�r���ZĹ`�1j�(!�LϔH7IҌ��U%��-F4�ܦ�H�H��ċNd��ZC9�tcd��)ij���H4���TU��*%��h��%�Ʃ��Ɓ$I P��8���i%�F�p��ҭ����#�5i��[DKhQB7qJ�B�]��
*�%G�4ܨ���[0H��hX�H-E-��mL��	�r�ܕA��%2�ib��d�XƖ+C���n�R$��&���)PQ�ƅA�%�KV��B�F��������]���-����Y��������圣`�!�L��]�Ъ���/��܌�W�w�J0h��t���r8p9mv[����t���qMf�MY-,�^LwH�[-������!��('FϦ\���O�"_a�E�����W�%�<��%�?l�r��&ա��AGwF�Y��:�H�(KG�h.53X�F�&r�'�x�K����a~��������=�-����Nɮg��NMr�5�4mb�.�|����`�Ǐi��i-#�Ĩ�P��J�=����N��X���ܽW�4�4�*�k"�lhq�Q���cN��V!Qvw3%m���$9��a��@d2�.�J��xc����E��C;�rQ|:霎�zkV�8?p�Ɗ�Q�c)md������8��ǐ��L�bՓ�����r{�]P�M�n6}�pf�{KcBS�Ä�ԧY{�����l�
��5L+w�M�s��B�#/������PR_gW>(�����0m�iW$-@S��x��;��R��KPp�g��jꆬwmf�����" ���Q��t���f"�u�AvXז���^v��ZA���1��-��$�Sg�˺����w��5|w�4��Y? ���<W�1>}��}�	v8 ��Q�匣s���D���35�;y�G�ưQ5;ZF�Rky�ރg��۱W�ZR�g��z(b�Lx`˿=%sKj�3Ѵ���WO:��3�|o`2�ڼ�z��[U!��� �'/T�c��fQ�4��ņ��<\靚Y}�aC�B�Ꙕ�]lP�پx�O�u�����Ԍ_"�H������U��������f	>���wwOC�r��Cp���F��J���K�-�^����aü��nn�U�ec�u�f�Ҩ�%ZVol��T�\I��=K�{ݡ{k���ڝ�6�jKg��^}j�nj�@�,��[w՜>�8qx��3���iǈX_��9��s@����k'%6K�����'g�e�����q>�^�?q�8	����Pe�<��f�H���I�U��8��;Z]d�	���;\�E��=+V�kYn�R},�5���T�u2x�mw[��F+|
*�4hW-E�7#,��˾)O;GnU���";��&#:.t���9K�GAb�v����<�q؄hz#��B̹���r�Vy�wl(:�q:�0-�Na��&�:����'�P���\�/y��|z�V�װ:ЕW`���1N3�Z�W�X>WWc���y�7�1�Xڗ��t��⎹p62E�C�&��J��[��0u�65�gn�Y	���,)�:4H��+꼼�x��)Y���2�'�;ruY����p)f�P��(����t����xs&����ϹG�t{��̝|z-=ZT[�����S}��;I��..Pvs#8�f�ڒ�{,�l��YD2Ʌчv+���z��X����/F	���/{�N��=@�'k�"V�K������ۻ�R���r��BO2��kB;�P��!<7�/�:�ݞo��A����o3����kr���k�'��;� '����+��.lM�u3���uƠ���ᴭ�n%�)Mŉ�e�nl�zcVC
���7�eF��Tp��p����)4�Mv�����q�!Ur���e�c��V77�%����:<2q�F�W� Y#<����Q����H;�[l��f^)��f���t�U���]��Z�q;�ꁾ����h�nІa�&�jG��>��YC��7�(H,MYd?W��/"��,mvf�v$�{F������0E4^{��kÃٽ�=�A���D�ؚ�9;��9�����)��(�{RgXf��R�6�^�A�{��-w�5l���������VL�Y��q���
�y�j���7^:�ؽ�W��B.�rg��h�/���'5&��o�
�}t*�X|�w2B\MϽ�)\LP�7��c�HPh�j.�LT2WS\"b����l�':�[�vw,W�]HsB��c�G����*\��}�ׯ;�(�S�Q�.ӝ1��aiS�v�.���y�����D��u�ʊ1u��
���E
b���7������̳��j�W]Y=�g���𔙖A۾f�kٔOyʉ�] �SU�ч���Uz_�����k^l�(eN��\��k� �E 3���B�mk�v0	{����Xz���<�����7i�������G�����}��~}}��k�v�_m�ی����0:�o��M]�bmf�茽9x�w`�����El<:��Y�S=������N��G�ڽ"XI���e�>	1&�v��q!�ǳo�K$`�s����e�"t�5rU,��b#+>�v���Ѷ�bDvWrۅ8�p�r�hv	L��{��j��z����V�H��{��r��ۇM5'U�&��+����5nV����hˀj��>u���ؑgE�\떮8ou	�]���-�
�Q�ISF�/k:�Fivg`���u-�y�	(m,۶2��FeZ��N̨����-I��q�U9[�j2;�ν]LR�_�|���h�N?|ղ#Q�o��U<�qP����-\y��)���%�Y�SE0����JTr�u��m��3�)ϔ5f;LK�X�K*X�&RPe!�E6��D]��+U�jͪ�b�mJ	6�'W$h�c�����ݩ��8�(+%�Vҁ����(�tVbVr��р7@�e*u��8���bQ
�Ŋ��B��%�/�J�IC%t��c�R�6p�T1]��E����*�X�4(�u%��l���c�Gw�V9A5D!yJF.ڣx���X�@�a�ƶ�Zd��{��~y�3�< 7��-�-����[m-g�h�*�a����hu*6�%Ճ!v�d�1�Q�T�Ү�T��w+f��q�"�e,#n���^�f"��0��E�0�,�؄�Im�.�Yye��K�IVE�.1�[M��-�VBU�+i$X�H�X�&(��� ��wwcp��+!%ȱ�R�0�%����*�).T.UI	#%F0m[.$dEX�i��j\
Z�R����%���H�X:�E�P�F�R�*����ߜǇ_��Gk�t���V�OjTk����º�s)U�I[p��V�U��(�@�r�H�,�8_z���ۏ�ᱼY;[�*x]�}q�	V'��z�$�;c�g>zK�K63��W�0�H<˶���3��u��u�41;;{{�6q��|ool���U�4���dc�^��;H��4�3h=�#¥Y�("c���;����¦�u��:�/��ݺ ��A�PY����80�:.��Jz�9��������?V���r��f�Օ����YFv���sk�,�����G\f̬NN�?��������-��i��}���Im�����R�Y&�J���I~Y׻����t~!K&�yV�U�yc���^:��-g[a�N���o�Mvy�6v-Y�Q�b=Ū����"^��uLca<YM�}o�h#��{�V���U�Ob{;kaܩô6��Gb𒍞f0��L�m����D��Q�P���?W��e���G������_6NEf`�-ǽ�9tן�f�[���_s���XH�Z���uJ-f@(0�K)�h����D��S����˦�]�377��uR�{����㡑�����|Z�j����Ҝڊ��#�j���Y�I)9�\쾓@u��������^rR9��/.�w+ō4t�[[��q0cU����#i^���W�Ճ	fm��8��&m�z��r%s�V�$�����g�9��C�qoM)�}��L�"��0r.���	:���x�8�8�-��F�L��Z�I�,�V^^��ߜ�ؗ������Ui+�6�q�A�� �V�h!����|P�D��uDKE�pSW0qD\A�֠j. 6�)����L�Ǯ��Yh��m��&��v�ﱏw~��D��Y77�'�[�
�E�ļC1V��E� 7�6��k�a���>���*��UQ�A��j���ZAs�M@��Q��*gp<�q��o'>��Kw��F����'�E+ő0� @��j�!KEM^1�y�j��('Э�q�ZPm�GeƎ#�E��1PL��Q�P���7�����F�ҫ-#UG=5G�v�cz)�]�R��G0Q�s :��3�/;���v��Te -(��11\�|֡��,�� �^�j�Hu��UM_��{��\��Ti-�Ai�A���މƩj�7)@�Ty(6Ѭ}���ԙ��X(f뢨��=�|���>Q�}�*�_B]nEt�dJ��.k
�:Q�Δ1.G����ǽ�G�L{Ѡ�h(=p�|���>N�S�G���֤�;��QiZJ�J7cTT���P�Aq����U�^j�vQXj��3��Y��o�C�A�J4�Kh8�y(8��KA�Ҫ��Bګj����U^�_ �~�s��5����|Uu�S:�FZ(�:���x5E6���P�M�^	X�*4R����}x��ʪ<5XJZJ�x���	�s"�53�bh����m(�Q�JJ��5�{p���!�8���8�f V#�G������ꪶ��*o�\�;Wjnj�ߌ�M� 'C1�K�Kž(�j(R"�_�"j�/�[mAK�kS6���lh^ q�QS0�C0]A��\҂�DLB�h�D��R��m�g���[�*��eW��(��m5�j
�,���E�� ��ߵ��~��YJ�U�GR��q��QME� m1}UR�PD]��^#�'���k��%�M�lS�|�dZ?��K�Ch6��[�1L��������˄�������W���xwZ�ٮ��yw�=�n�^������^V�]�D��S1�}PCP9A4y:�)U��m0����g��VZ�h5#�`��c�/ 1h�
\䣭Z}(�W��U�XvU�E���	{{��y��zPu��ƫW� �P���СK��E���\j�:N|e�E�u�w�����CPZD�%��z#X��R���+m�7�ﵰ�Pi�� b�6���Q���%P�F��h���W�����}�0�P�6���)�h�	�MAK��U�Q��"�s�6s��6^��#T|�tj�J�A�>L��ZPm5A��Z:��B��AdC�)x�V.�یݬ�SIY@-�8�)�p+L�TO@�WZ+�J��Q���UV��UG�x���c_w��m(�y ��U�������
��*��C�U��W��Ag2��w�L��C�M<�|����o��1+�寮��v	ʂ�&j|s�w��+��w���u9�]\}΃E( ����W �_��F'��Cf����~%aU|T��ҿ?fN7RE�v𘜯+�y4l��n[�\Y�}�v OO\�`J���g�t�s�\c�+_.n�۷�榽5�I���g��wqxc2�u�g��6`MJT�c�/����^��3F�|�1ٸ�F:1�}&�C��Yv����n��@���hC��4�_�O�c�HU�(Kܕ}N�"���םq(Z̝H����u]����o/�kp�rC�{�*񤲫���r��={�
�/d~�{�/'N�~���8�t=>���!��mkW��~��g	k[��Q�а�<34�9�,���
��Y�&V����#w�$�ox�"Fl��Y��QmxDl�a;)�+Ю�A�W�/�xVp�tښ�L�i�M�	�jB*��v�`EԻ��f�S���ڀ�&,�BH�r2�id#/�w3H��ĕ�p�}��X��I�u f�m�ȏz#Ԗ&������E���{R���gkT�x����R�w���qD��;͛�N�'`�כ������=�`A;�V%fP
m�N=�ό�2#�����J�[�Or������l̩���x +�pg^�}��K�;�8k���G����d.�*綻��=�Գ��I��Q�G]dyzp'V���f����:����ǰu�AtW!�:������Uv�2pC6\�]�rఓb�r�J�i��1��D{ގ�z���[u���{���ߥ����)��mG:��������aώE�=Qw�͗�ٓ��W2�����Zr��M�bm�ۺ"�Et*���VC'��9����l��u�/�wA�1�؆!�x.��Ԧ*���3���a�v����q����Ռ
HzI�5��g�:a�=ѽ����N���k@�3<0���h���ҫ����k���>	����K�r��
M�N��)���䒐�3#�X���ۂq�V��8�v��Ac�v�qT��4�d:���W.K�Eꮒ�8�X�N����ˆ�W#}����I��*�D5j��U�����)���x5��dR!r����hR���R�e]�Pv�v�.Ep�&�s��%���跒�T����mQ�.�"y.[�7,:z:b��%:ڶ���t�b�{c9٪N�,&�v��Q�os��mv���4�Q�����%wH�_tڐ���m��JZ{f`5�X��+�� C����QֳK��*C�ĪE��L��EV(�T�X�,
g�'K
YV��7���9/�B��x1��]ZwW.��ZMd��*�#��B`Ѽl���.�Z�8��9D#iDJ4��V>v�[�L+*O�W
��[&.�T�h���[��[9�˱��YS"�-+FdʸQU2�FH��M��0���E9���jVE0��&| D�� H�Ma�2VZd��;����\�aa��"�B��)_^]�dӦ�LV_�G+
���9��T�]$Jf��GL�$�e���N�F��b&b9!H�.�(��R�4*���F�hE>�mI(�Ji�DQJD�LH��D��6\҈�"�#���V�J���X�$"�()��*Љ���ܢ+�(��X��)V�P�PU%���P�J��F �a��������4��B@P��(�%VZ��*D�+J�D��QR�3"�%ah��svID4F��TQJ�@_y������=Ӎ�wC��ɒ�=�j6[;����G���wa��ΓU����Č)Q�}\g��h��B�~>�)]���F�g��j�G����-��5>TU�}�B{w���6R�Lm'Z^ر0�^5ų���7�`B��^ë�sWp�3����7��H��{�&p�&�ĤC��U�ꌃ5�3zYfV��K�{b.Î���b�=�� �ꫬ��jJ�Kd̅6/:�a	ұe��M{2�&7�;���!�:����Eo%��wd�e$�=���7�z�]�5�1�|kFت�]u4��5��zvr��풅$)PԮ�3�w:��IH]h^��z�'�W�c�����ź_�=.���Ȓ=�K+*�=L>��w����:�!@hT�������{7�No6%r�Ie�p,/@��%�!#^�e����L{�Im��K6��oy��!/8�i u.ݹU��_�Ǖ;���!�]�sa��c.���{�6��]V����@�A
�Zj��V��~�7����o[_��
���?�خI#�h�gj�L�������{���³�Q���1@�=]���Vd��!C�2��Fk�	�ڬ^����z
��%u��N���<�zd���b��ϵ�r�>N���g�!��>�\�Pw�b�q��5횫�V�Xv�oUs$u�ȸ�{�U�ᡬ}�:34=p[�ݚy�uCN�=�  WӬ�n�����m;�jlU��ף�e�G���ż��DDz=�bk����p8���ڙE�`�!�|N�-������[n��\��i�-�xA�8�^�v�`�f�|د6����	%+
Ş87Mv4E�j���<2䲛��EG�Ό�E񑆡�z�ʀ�u����ї�n��q�����k�u�]�Bd�^�B�'3w��Inl�'q漩k�UO�`:�M���k0n�r�.�����Rv[��x��BxGR˘��"�4�,$b\��DDz"�f��~���L�6#�4���\����ӏ���i�:]�uy���)���=6\%ʺV�N��Љ>�漢~��A�n�sid�]'�@9�\��o�>�
�(Z��Oj[#���rc�xf��{��øE��J_�74|k9b�RH)�м�3������>M�/�&�A=��Ppfʔ�v�+��G���I�4�̫d`���v�-�`�8p���y�W�n���x&��侈��z7���ޔ3"�0Oh��h�폲����CH�ܣ:�:����QI�u�잕����m�gF�:�ߧ��ɿ@�(r 
�{���ҽ��fLֹ�TmXGL��y�mw&�:K������4n`ƍ�|-P�=��yȪB�M�|�!��]���^���I�Ox��"f�SMh���noX���fV����:;�����f��>�5^��v�A�	��c+[�5U�fc���7z,�[-�����;��\����{�fn�o0��z�������z.�n�rz+��\�{]�k�*�!'���s.(�E�W|��d'�m����ͅ[����˭�=��F*#Sj�m�53�ޤ��B����TV��Ŝ���Z_�ӯ.rEz����'Hh��2m͈�f�P����a�QÝH��F>�6-�Zʋ'C��l���Ǫ�g�	��K��wT��f1[=��]m�>�x0m�i3: 	 �!N�����3���(Q�}��4f��.ۥڇt��|>%r��G/��lU���4��C���=��-�ݓ�GWɓ��F.�#�5�Bdu��N���Y�	�#�`B�Zg�=�Ǖ��Ð#�[�<�uÙ^�`���T�FsC^8v�6qSN5]YC��Xu�^�N�f��[��2v�5��ԉ���\'s)��g�CM��0����p%��6$��T�b�y�0�88�un2X���,���+�Y��}ԞL8�=2������G����5�.�rTg��F�6{j�F'<纍`�@�%���cO�о��y�\�Ւ�K��W��^oZ�t����$�`Y�M\���t �ha`���{^�s*v׭�0�9��wCf;!�%"^��(�t��B@$H[A>� ���i�;1j�c&$����I������"p��:黶T˺�h.�e#��G�`d��46f���Y���@��S댑��`�a�%![$�5���꯾�����	/�~e�uJl�U�_����t�1X�
:���>�Ff�c5�����9J��B�A�� ,���'�]���wym�rU�r���iv��q;LZ�֛+�� �G�"p�I�퓒��&�C�w/c���=�D�Z�����iTHї�e�7lj��\'���R�av�D~�6s�*�R�Z�_�
;�����U,���w�:�f<Wy�뵛��4�Uv���JhAq�\;h��uIZ~�\zRv�\��{�w�����d��k��H���r���fR���[F�m����[�t5��Җo�w�d��(�e�c����Ք���W����#��un��.�4��a��%AO�$�A�=G{��J`�;k4��ا�Fc�m�e��a����!c� ��T�2m��>��ˮS�f �⺝-��0%!1��"�d(0-(�V�(��x8������7����ӐX�κ�E/6Ą�Sz���Y�X�I��e�d+�A7`&%�2%N�]c���������Nc&�K��Db͊4"�>p���	�5�+
�mV��G��W���U�uن���@��'���[�y��j�V�=���wO a���+*Zv�^��8P(d�$]���JcX/&(q�j���
(RƲ�ej8�nI�B���Wd�Z��j�]�m��M��N��M>��H��ْ	P#B�i���)bF�U�j�KD�ڙb�"�ӈ�������E�``���Z.P�Ȉ�UmF�F@�2F��dT �D�Qj��J�Dj�Ai0�L6�lH���DiTPQ"JT2����rIQU�r�Т��7��H�Cj�ږ����F$	�Z\�T�
�Bґ��`E.ED̫�����U���U��W��':������p1���~���,a/׾�f���{J��Gs�A^��␪�k���c�b��9+�z��s\M��~�z� ��7+It'u�ʜ{o�� -�뱺�Xm�ͧ����croy+�:Qث�q1V+���
���]Cv5�X9����X�W���
����j�pS����W>�FN�Lm׶na@�0�ʾE�C22P�b�_��B���-��"^\�{~��[j��X�"YTM5aCE���;Mw����gF���I�q���΅m���KJ��^����ӕ�|ē�׎�J������w�W�"�ݜ�/�OE����8j���*�{���,���'�Κ��ɹ�ӷ��k�������%1^[�>�AqѢ��Y���}2k���MyQ@
�~5�kF��j�p�F��:���ǉ��Lx!��k���Ы�~��k��Ǣ�W��V�̓E
�l}@X�N�
���W���fL;s�hk5���G4���/���@n{�����L�n�ǍZ���b�e�������R����xhܫ�@h\k��1b�KS/-�%ZM`B��SMR�VR6�R�
������pAYBU��4��Ұ֎F�Ѻ��y�pD�Ύ�iw�2�����n�Eu�|Fw}���bor�p��ZWcX�&�x녊Gc�w2�84P�V�b8**�.c2�y�O2<]fe����pf"��Zd�0�Lc6�짏7�������aebX^4�]Y�����ӧ�y�5����q�
Vk����H(t{MA �Z��g�vj��Ҡ��SϞ�·O���g��%�w��b�`�pX��(��֕���l��F׭ܮ�OqLWy4йO5��w��\�ܾ�:�y!�M�15�]x��ў�xo|�y��Z_C���ァ?u�B0!�yՅ��j�ټ�5b��xz��l�]-��])7ysLɕnr&�I,�9]ѹ���d^��=�-(��7�}������c�9c����%l�{�u�gW��1Լ�O��T]���U`�PT�ݧ�Z����8��Ӵ�:����� m�[�W����Q��p����b9W���*}u��'�3�~ɍ�|�&�����������lk7��Y�C���H_�`w�L��W�ι�ޡ9M��Yjz�wͅ��\��B\�
�1��n��j���ꁭ�sC����j��P��tTS�]�Y��U�{g��c�0h��P��>�58��w��Ν�EڱPW���x��b�"�R���� �����p��~�q�u9q���y\���h���)�칣�Y��S������s�ϻ�6��R���[L�V����>_
 CB�����q�[��|tk��T���I�t��u^!ЅF�јt~��EMą��U,�㡎�s��n	g�7M�����hѨ��..�7ܟ9�w--�X��+Z���7E���zǽý�4ڥC��S�^(��ע;Ƶ=�gϻin��`����M�iȚ���.`��R�GP�4�n It�	�@5�(���S��������KP\����:�:��n��(}��V��r���]��K,v���B�M�a�X�+7ˣ�y,yh;�,�aI��U�ƙ��7�io)ܞTG1P�d�}��M�ɋ�Q�kG[Y��ɺ.В$��o��h�ҞZ� �� o�ǻ�=|��GC.m4�g��LP��k
 ����@u}�*�7e�գ���xk���J_���Y�&����b*�
tN���a����E1��5�V>b��+E@�q�4e��>v�{�]S[����u�rI���m�����ӹ�@�8`�~�c�ޭה����{�l�o	5�u�\�*��F�p�֫gG� ŋ	��̓|�Zm�qy�s߷�_������4��&Pȗ.a;��!��L����%��UA�r�ׂ���y�ӱg�0ʔO	PQ=��^�̣-�M�X�u����ｓ�C{^���ߐ���5y���[�EB�,S�����{���.g�@{Ʀ�+��s�ܻ֫�c�"�4��
Vh
�������M��i��VЁ+D
��'eB��[:4*�Z4v]���n�X�~�Q|��^*o��Y��u��ح �+(p"�g�PR��CD��8�o+w���+E!(R?f +i27;72��h�U-��pf��`c�g���}�5��ϡ�L��Poz�4J�*٭Wn\��8�|E����Qj��� T3��e��V�Y����\�=튥n�r������(������>��xI+�{�DG�AZ�:�ꏾ�>S�nSD�A<�ǜ�ǵ�+�SsVwܵ0�74����e�5�{Z�82ǃ���ѭ�5Ⴗ����DV-I�n��ѐ�F�5c �̏�׫�/ፎ��{��ǆe�G�!��y0l�|�f��4��.����c績��Q�Эv���S�&y]S>��.5c��եR�<<�1�{��H�my0��_�k�7&�2�oɇK9zG0:Ɏ��\8h���"(����s��z�����j��c�k4�b��AP��
�֯�:�PQ��wF۾wӫ�N�����/J��6���sN�=ώ_mN�f����v�v�#9/��@v�v�e��Vсa�ë�n���R��7���r�1����2�F�a�^�աY��g�Q0wd�/)�� 1��6�S������{�`l׬ئ+�|>��Jz%/��{��X�Bt��Y�Z�M�̡nK������'N�d�u��,v�ӏ=�-[n��W�Y�=���5<��}����$A�j�������i�	��\��8vu�q��④q�5���ƌ©����k�M.����sx��ǂi�VX�v�u���]m��B�?��E^�-��K����B���6����r��`��W�̄��a� <4Z�S�^r���� r_9��b}������!��F�v&&b����8���S�n"�r�u�&r\_��EU{or�pv�Oŏ<_g�gFx�]��(�a_S���ڨ>�¯�Uh�,L5��1Z+Z����3뗴�όMLt��=pE�Wg����B�)7�k�Ǵ�^}�j#d
s|��S�#*2�*b��X�HhО+�g�@��T��Ȗ��5c��@�Ƭ[��\6w\���b�M��DV�c�����^���K�J+֩�L�7�F�T��k�y���&��D�o�0�,8M�)	�^8,��,�՗�^����U�K)4�]�er�
�Q�PNXW��5+��o_-�)m]�%��tPS-��Bg�p�ߛdˡ]Jޘ��a9c��y�g��q�=3�cm�Ff�E�q1q���GR��w�p�R=���ZZ	4t+_n=c8��gv��T��wuH��Nܧ6��][+�v*Z�U�멥�*�[ۻ�*�䳐�)a;^�
�����ػt��3W��F��H'/ow�������%-�4�8w�:m�.ʴ�y��@��˗��f���Ȥ����P���i�h;%E�u�K���0CZk��0�ͪ�*[jm�)p�1��=j��mf흏i�T�n./,�o�y�[�bx���P]����U���i��3�(�S{�����E��ԏj�o:�U��X�<���~�uf ���^��;/&���I-�Nov
�!�3q�*�q����s������E>6e.{����4aZmf�:��<��m"�d�T(Yf6D��"G��ܷ�!V�}0u���	�ES�l�vS��J�T�;{����u��mCS��WP8ȫ��Ĺ$�K�$�H�'u�����u�H��"F�Ȩ-��"Ԅ%*t��Yib��cU]�\�R4C9�s"�%�ZJq0���c�\ �-���X���m�p�s�
�Q"�j(�RJ���*4�H1%ʥ�F�g&LHʌ���v\���9�lV���b�m˻s�V1aarF��r+wp�0�P����G��_S9+�Wl��G(ngo%����[�C}�1�^T���~�tɯ��kGR����PX��t�d!�^��$2vq�x��wW������o	&�b�>�,[?xrw�8�6���^&�u��09g%��'/L��mGJ3���\ɉ� �y�|��Kپ\�����@w�f�7&R�yQ#�eڪ''T�"T��TǛN����r��Ӟ��gP��W��a(x�V|5��^�n���G�׽do���wR�12��+��u�ߦ��=��*+� B
u�Lp"��Xk¬p��=F���>\�d'�=�}�������>^���e�}�ι��@K�r�/8��F���żS��������׽��`ɫ�f��-��'ԇɚr�P
�GNWVՇ��81ꪱc�R�z� |�0��5����u ����Adn���c�
�4F��Y1�X��"eyJ�u��f��n�QO9oq�3|��87�g�߽�5ǿv����0�ӎ��y�lo��1�u�z������e�ܮ9ܮ�q4^�%�z��l��n��������{G�ë�4o.�:w�(�N�&����H4_a�����ζ��9���}�P���(*��V��T=�+G�V�3�N(��y�^[\E�ͺ�AENX�Q��\��G�,�{˃��8�8s;����w�UT;�s��	���}N��x�hK�uf�̄`�z�u��r�dL����H�_%�]�]��<�7�Ze�:�h���U!"�B��^�l��ݲ����شh�5u��b�S`A���P��vO��խ@1�֜�L<��V	x���ə�pAa���Dp(��vW\�HPb��9��=]@P��z&�m/5�s�.��_��N���CX���x*�L>P��a@�޵Dks����ZpR�@!�m�X��k��/a���:�ۿ���)+[�P����{7ҽn�u=�Ȇd-H6��X�=-!�-v�o���C�&\�Sҕ+!8=�OQ�9��PV{~��}<�1���=!�cֵ�=k�COL�7/�Ʉ�w	����T
�<�h�b�h�S���[��p��(U
l�B�/�Y�
�1�׻~�	_��2j�j2��bu�uލګ�P��j���Y��:�7	dA�Ug������6	��mr�*z�[U;;��^yQ|�=�|j}����b�%���jVWK��^�Q)��^�+D8D5�Z���("�q�{���`�ǂ�D���m�t��᣽�|4�}�c\�}XM�w��M6�M��#�N��t���F�*Y�Vb�qb��v�|=u�q<��mn�\���M�8�F����	؞j7;���}_zo��cs����:L��:�s.���?%���׶���=�,_'>�}>[7�\R��BY�X_�ϲ
��h�������xA�?,/O���=��>���K�`�*}���o����{�tkކo{���E�ʂa�p��T�ga+��&�8g3�~w�7�g�<�3ͻH��f暿]�4�W�Ht�3ڲ��\,v�MOr�*P��b`z�\����Y�L:�^=M��v�.A���1���Z�K%�>6=B�##�b�9y�] ���T�{����_
~(
H�<>�4o*U��>@h\i��D�{���ʻ\6��n���'f���'v�ڥ���ÎR�z���wh�6�r�ݒ#%}�kR��DxR|�D�ʕ+�h�a
׋�d
�5xՋFb��?�Pe��X���Z�g�)ի��cZoɕ|�Gۤ��3
Zˋ5X����*`Ȑ?L��.!�2�x�h�A�^む�2��xՍ>$}��ge�bǬ�Q�8pf"�e\Ø�'q ױ��{9v�.eѼYn��V:\��8w����KkC�)�~�\ϰ�[�V+�|o5R8=�g���T�@	��va���8���Y��8)a�>��Y�
��o�n�p���cEd��@Q"������ݾ[i"�����u�+�,��K��JM��7jFq�+��jXG#�ǀ����r�|ƎBb3������Q�����m*�C^����ߓ�n��+��0Z�{����7+K�^���hޚ�󼹓ٰu|Ɖe8ʼT��
#C�X;5�Y�n�׶8��>��SO����q������%dW�D��b\���i�`>Q�_ny�9ȷ���2���{y�;8�L�]�����C8����R�wfc&+&8Ӝ�jԑQ(`A��){��{��1[�cC�`�x�
��.5�P]�������>���]	�Z�WN���cV�,H�|w���y�������y�U��]��dn�#�򻝬u����ΙwL�*�ck��1"����䵭��MG�3#�H������TêF��E�V�?����t,V+�f�_܎��1��*/-p�Y��_,��'Woٱ�nAf��۴�s�<��0�L8y�������`�y�eX�&������ڟ�̝�T��`"��{U�׏��pޜ=��4}!���ES4�p����g��;�m���G�˩BޠLO7�y��19�����Hnq����^���M�io&}��+)����,H�gt�T�T��9�0)�ᑵ�7w���Z��붙0�{����o^e�Qز��đ�b�%�������O\=x�H����UF��Ө�����r$O|o�
�7=.b�ya����+��:Y���q^���f��@���*	�Z�}��j;��*��X�\�w.���W�^�W
{]G�J�[��Jϩz�j��t�/��ٺ��	����K�����
@R� ��f�^p�2�;"*��~#�	�k��5i�D͛&���n�ڙ���X���n5ci�HZ;�e��xV�]C���R�j����xK��;[^�X��_�WP�����Dօ֩rT߽ޛ�^�}�V����Ĕ��{�m"y��i���sy��1�Njb��
�h^p�~䬗���l�3�������13/�&�<{�ô�n�mt��r�E��$����&�>f�/�?iI*^�Z�6>�,!��o\����35~}��M�';���g�ޞ�_y�>���d�?b�u�ԍ�s�6̻�O��LL�K� _��M׹V�XKXׯ=)�U�	��:�e�"�^*�����V�Gm���>�bY�� �ְwr7gE��V9�Pd(PBǇ� �	C%�\ϬS�U�c�b�(x^���4���,���x���� ���mV
��P���v�छzG
� T�(4UKjǅFpg��E}�v3��ǌr#ʦIV�tz��R�����}2�f��"�T�O>�A�s�M rp�Q ;���zE4Uv���wM��j1��e�n���@����f���L8��<P���l[��7t�/��ۧz��X�2@gR�ԼҲ�+�\\�cTRmjYa`�5g3�n��Χ��y�u�]>C����c�$x�Y�c�̺�pX(<��W#�A}Lf�]ND��,3�&�ξ�;h���]�;���\�G-�ܮ�pCZ���2K��6���\ԧ �[Z*3re�{\�b�N+9���6��*�Qa	go���l�B��َ��lԡ���ń�2ӫ�
.dF�s+/KHS�g`�٤�*�ئ�֝<�i��#��b�Ď;�����Q���:��T���rJ�����d��
&��KĬ�BUEWf�57���ɝ%�rUO6-�Jl�uT�,�:)Yj��O�4��ˈLn堝��i����N%�]'�p��z�K�@�fO�;�T`m�C�Fb��1u��ΒFؿ(��3tK��֦��Rޚ	�ԍ�,N�-�Y�-�#��;���N)��
�hM���a��Af�ף��)��E�u������%3����;�it���jq��˼��wvr����t��Iנ��*�Um��_®��*4���uҴ�m�̋lj�S-K�Y�I*�Y*
-\���6�)���Jj2��Ds#T��4��EZ$r��,j�+0���P��U4�2wX-GR82�6J.JnpiK��n�"��2�EZZ�J�����h��\�EQS)z�?�f���>������ԶV1�v~��R���]�K�o@��&�˓>�Mx�Fg*:D��).�������NÖz� f��{�!�%�Ŝ���o�����%�Ovw���-u�f٨F#Wd�|lX"����V��u�@�*i��эfg��s���;C�l�!�o�<��Xw�h�/��q�{�
"�W�⾽T���� ゲ���W�����׆�Bŵ�.OKt����I�q�;����g�5�*�2�}3��SʼyT��m"x�ۗ��L����L� ������7��VvV<'��U���U�ئM7�"�_Z�[�ּ�v�`����Ո&,������u-}	�ՙ�s�\��г�.�S�Jo�"�y�K�S� �8)���kE��L6~����r���-h��,�������ZP�q"�N����[���fWS���۱�i��3U)��}}���M�N��|��2�ny;ɷy��{��n�]ڥ^J��X�  ��,�0fx��e��4Փ���o�h�+��ǆ�)㷎f��1�C��m�ZƬ��i�E<��^�/�����a�e,r�.����>v��ƟN�ADz�ݧ֍�0ߌ���,��uù�r$O�N��2�b]ny��N�u�&����_vu^�2���s�up#�|}��7��(]\��K���Mfsً�YEWq5�׍5�B�	.�#�a��u��ѴJA�DAR��!�0�T�"k�g�QSdZ>�irӚL�����P����DS'� �.cw���=�Z�z�]��m�7y�a�={�E@�׍j������+ƳML�ˉL�.oU/j*��i��t��f�{:���>I���}|��׌A|ˁ䜑s�3"	�7�ؘ��B�9�)��|��7:��I��x��f3�כ0��]^���1���m�#��@z�����FP��c����ٱ(AV<=�g�ڕt8pNՈ+n�:�aO*�V>BηOS��F�������*�n��-��Y��񮙋��´s�$
�@��L��؝�<*�0n�� �q3+��·�*ǫ5R�O?��=m�7�=����m��&2-��B��ם��jB&�ҘR���ȓ0+���V� d��+��y�]y� ������t�Z��a����{$�C�'_[<����!��ﲴ�c�7O�㡊" <���@u�~:j�W�<�cֽ�[��R8�ϥz{��	�׾�#�W�����Yf�ao��p��\;�+2�Z�u\�[���<5K�(XC�%�+(P9=��Z�݊�,T�hnKꓣ�x�L�{x���t�4vc�19�p�ֻSU����-�Q{H��cL�Ԓ��J������GƄ�O£�gl��X����8 ��Vk�*�ゕP���0��3�_9�L2�*�֚c�iѸ~���>b�B�a���&�^5��(��w]u�^���k�m��#Wv�|����f��c��[�`�g�e���ƍ�D?�����Э�H0� ����HX�F���5u5V}P+���������� �r��22��T��_d�^�WP����G��i�b"e䆻<����<q۲�<�s��}�c�1�\z������W�񩵷fc#źUp"u;сLȱ�;h�)K����nj]wus�jӘ�8]�;;zt�w�XĹ}�w^6�{�g�W�l����b���
��{S7�vCC�=z�T�EP��
����5�RC��;������ht�:��r�L��:J�6���T#Y)Q�)�.�P����G/7إ0� ���b����N��f�T���lnC��#1b����+���wI����qk\N}%/V*��Z>��5D0f�L{���96w�_���q�N�I<��ۯC���Z��e��T�V�^�^&���SuYm�7�|�-�F�%�6/����U���T�͛���G���Y�u�w��D�N�	�*�ԫ�9����gP�����.{���5�Y��6��Ⱦgr�sK��m��E����V&�m<�ǈ��^�!��#�w�����]�m���u�k1N���ɔ��J�I����s.N���QPs�0�:��z��ͷIi����i�B�#�[��%�z[cª	e
`�����w�Cf4|�Ie����}X+�u�4+��|*�C-R,���_֍f���:
�,�@X�(���w�|����؀�j��Э8�ʸV=�0l�j�y`T�g�Ee�j�=����h��f���E�(���Z;�ǆ��Π�\�Qo��>[���y����*��!���m���IV۽�ܧJ�4�I&�;f0Yؽ��R?z_2���z�Ɋ�����<6��F�_�佷�A|kt�/j��n�c8���+ �:5��z�2A�0�xV�L	�\XY���{�[�JU�;9����v�̚��BnHvn��x�|�=ȧ��ʆ�?%X�1�b���8��m+�y�@�]V���~����(x|5�e�"��}�˷�]�@�E�Xٖ��f�mh��2:�Y��J�^�ƫB㢴|��]P�F�E��"[ԁ<k�
�~'H��U�آ><m5~��s�U�E�1ƺ{�i�t��uҦIUn�	�Kwy#�����^��f��wn�1�K�$��\L��ι؆���u�Y�s��=��_g/m�b�~\831}~�*�l��̙��g���_M���V�>�)F��6>���V�r���D�j��@`���M1\�O�����
�*�p*�X@���>��BlS�+w-�'f1����sf���G
�v�E���Eo�ϡ� o�������}�X�50�4@�s�Q.]mh�%�3��*]+�l�2k�wl�	o���b��/S.s�:x�I��wY��O:����
ݛ�҈G�%��^H��7�����>�!c�s�.�억]�4b6/��z+i;�\��k��I��(�0-r�24�7J� f�I/��+X���}߉�s��h��S���RuR�mJ%tV'\�U�7��(���	����.ᶭ^���C:���U�W��Iu��>�]%3e��\U$�O�l^�87��8��+&�kkp�a��p*
t3=*��or9��\9�A���^�TKWn+�\i�.���MK��&:!��7��A�OP�F1/r"�LQ���4���0z������o
͡[O�YX���	����))����^'��sv9^8+�VK��;��������z��p�]�Y��fc��W<m�<�=�����ꊲ<N��#W�a����u�{�Y���获U���;+m�.eM�����y�b�\�ɷ3OX�a���qݡ2�&�ެGq�RKo[6�h|>�f�`B[�po+��
�\3�q���h��h���YY+^�W�����q�g��+�<�_[��9�[}$N�����Q4��+.u\�=�o:wȣo�n�s��r�`":�:n��˷��G^���1Ք�VT)]&	��B�����b�َ�D��3.Q(�]\�U�3ੳR���Y�\6�-٩�H�����hT&�ʄ���&�� j��*�X�m��T�xhd��"V�@*���8@�X�CM*���Uc!����!�N�"�
t�S"T*�"��u�����;N�'������Q����+^X��v�4o�q���[������,;��"��.�S���eܕ��q0�2�����4��t�H���-ke�ƅ2��V��WWX�n`_��-X�F�ղg����եE-#rTj.�-����&d)R�ai���rj���֥]�UMH\$�3	�4ңKF�ZĀ�D��	JI.Yt�%�P�V�-"8L�ѹb��H�
A�/Uw)t��f
��D��}g.l^�s�R�C���fجVzCZ�̡c&���,X�G� #�H�\��kt�Z����M������|ĥî�9(>�?L��w梺��\i�\I�����>��m�� �+w�(D�1㰮��^S�U���U��w6M۠�}.g�Sy�B:���4��7�,�G����i��E�]xͫ��\�3� �v;֪u�L�F������w�4���wj}t���5�j.=j;oRj�t3�Rnm�b2�3:���e��ZpR�y�cK��^2���_,~���?~8���cr�Ӄ�{�2��pU؅%v�ܤ5�/k(v3�.��&'�׹����/��t�NdtL
��U�����ހ��^p5�g��V%�VL���>�O�t�Q����a)�-2��5�J:�7�cQ%;;5�9޲��J��/�j��CU�X�5Xd��VĹ�f�,1�8��
}��e޶X�0ͩ��&��;�@��/��pq��+_)���g��M��;V��Tc��q�ݔ���:��`U,��(@76Mb��	���3˅.�e�UQ{��v���Q.�w ��sB�(�(t;Q�E3Q܆��͢�����z/e�T��o7�)7��$���.x�#uz]��`6� *^U����#�s���+��A�aH�{uz��NI2�u�шQ��U��{<{�=���a�;Ia{u;��B������];r&�xG,���6��,���3K��p��C^�d�U�ێp[��w~��;�w��9�#o�1����=���U�%����B��-T{�5���K�TZ��������(z/^3�6���2���������΃X��n�����O�]Ҿ��6��ߛ��c%b>�X$k�����]`Ǡ���I���/('[s2E�;��e*���v���
4���YY��qR��)d7�<�����+�X8�i��v`��ND�[[�!��j��ү��[��ox#|�b<���V�\|~�z�4�,���õ�����>$���޵���OC7v����n�i���C���1�d�GL��1��(�7�w[�'�IC�(���w_1tw�=4�X��rj�5}���ZS��E�����S�H�=�GdG@O���6������θ��n	t��'��tG���i�y���u9`e��A���AR:m�M����d�����ֶ��u\]��*�l^��7��,$bE}�IKZ��X��m�(�����<s�'F ����m�\�&��^/#�T�S��av�ۨ��-c���{�jr�_Y�rG6�B��=ѧ� �+�Hw7g�M��.n�^�p��k��5���z�ȟx��Ʃ#�:��"���+��-�ލm�;�Ձ~e��C�9�-vaN[��+nL5�6v� �1�1��G��"}��&�!\�*^�o�W-�ფ`b���سi�ǈM��w~�ku/bq�~ϫ����	YQ���.�S�kf�Y'{����v�L��ך�1�k]�NE^T���mRt�Bu��z�RݦF����Ne[j�Ou����0T��w��dL� N"fP6�Q�Ǟ)�#��&�>�p*짜��7��XF�,B*�q�Th��^�˗�+��#��p�ޝ����_	��
�Oj\�0_ej6�{'Y�	�����E���D�ؚ�9;��]���3~?5�9�^M�E\��f���%�o��T�l�����N|z����ԗn�Sa�.�&�`�~#0οR��;dw[3+�m�f��vk^^����k�;��8�!i���̽�Ks��a��/�CbV�yZ|	-���	���^����g����9��s� y�Gx�(��R}�x�]ʸ2��7G8�e��۶����6��y���Yk��K�o�$z;2�K��
E��c߅n\�����3�[|�U� ��LF1�}S��SJo�f�X��t��P;p�sT��ܬi���z�V�j:�%'���@Ź�t���W�!'C)�v,��ܷ�k{ڒG��y������ػ<�����M�}Ftav��������YQ�6��`�݁��3'�!n�@��'���7X��D�0wCJ���Q^k"���OkEmZ���F˩�:�WwP�d��aP�ԍ�*�Ἳ��o4wѼ�҅��{����#�=�C٣	ݥ��D5����U��B��s��.͚���_>y��!���x`jVu�Rm�Վ�Z�ȅ7��x�e��eE�=h�Ś��gޛK�B�Ig˦��ݴ�.I��ʿ.(N�zC)o���6�c�A���=��gO,-����Ll
�k��|2'z�f�y�!������LAԴ$,f5G�͠�Y`I�GC9��Y����]��خƪb��<������Qԡ7((�����Ū$̤��
��Q�9K�eC��>�x��ܝ(S�,wX����cД�ɟiV�+Y�i���\6�8۔O�R�ц�W�� �
B�aB���^RG�V���
�&��Wؗe���:����-؜� �c:����nZ	Q�i��j���@��dĂ��V�n�cf|[�����m D3 ����T�ʏ�]!%��
11J�|dG)���vg�e0�`h�ԍͬb�,�������_��)][��(7�\I��qVQ?�L�[�A�M��<(���Ѻ��C.�g� ��fG�b�o/Bc.�]5�h�{��h�*�Ц��?*�QHeZ��[&Z�?`��-�Ua�Lp�������-O���X���B��u�`f�^L˄�Q�u�:u���Z	bgVZ�m8e�.�0�x��w�P�5�}x�tE�u�<ß�`2+Ŗ�,�@I�
�RU��+S!/2�ň�-'v�cF)��6LÉU�Z ?��lB�:�=t�Yi�_Ƭ�"qQ ����Ը�Y�x>�!�-$���H-%ʶ��j��[l��B�Z)j�"��w(s+Ma�QDD�",K���Њ�T�A- � [�2�����QE��j�B�Wf1wB�m�h��K�$IJ��(���F]ݶ�DR\�X�i
�4*�"�x�y��C9��Y��8�VoQ5�"�{�)�q._�zI�������)����鲕�9��i弛�p�V?^��}wW��2���&6�D�;r=��zh5�N�uz�ɹ�|M-��|- 6Ǝ�ǊƦRX�ށ�,i_,��*���g���w�KJ�81/gu�o��S2�_]+�=~�S�y��dk�0�d�r��3Ҟ�G�R>���{'����[��u�8m�H�8�F�Lg�7��ȧ>��#yd'Vs��!���N����/�y��K��[6Eל{:M�	��?ՊK��	"ɇ�z3V��/w����{oݪ��Fa)��6YƘ튟=���z:���tG&�
�'��U䒠ܚ���ݮT;�j0LOG+�n/OyN�����V���+�k�\q��Mr���$���'.|�a>ofL��o��d�v����\s�#ї+�E��6�̖��y�[M+!�}�잧&��Ͷ��[���hv�L0��;_e_5֖3{�L�ش�I/��V�C^�}��P<�/���ڍVn25�O#7�Z{ً�&=� X�a��-z�d���k���%�%W}��p9�f��w��=�@��P��(�U�9����5WT烔ͦvڱyƯGn]��E�_Py�ݖƈN�X����՟:�)c�MfXs/mS��L�B��ej� C�N�׳��Ȑ��q{ w�<��n�q6�`yB�@u�v��92�Ì�ҳ+�{�Ԟ��쟫#��.�{���}\���:@�T��ܮS��>{�c�au�^����u����(&�Y��Y���;����u�5�/l�|Y�q�F����'�0�ʋ�cHۤ~���Ѕy�7���V��׎*�;p��zOn�	�y'vb���C|t��9�Tu6�ҍh��	K�J��D�=M#��e���=��_Vf|���U��m��������#�Q�&F�K��j�f��ߑ��V�X>����%q�
U�0�j�.饌�5(r��g�c��1���c\6;��n��9���ۙ�����Y,���bj�
�Y[��پ�6C��qf����6��{��!b�P�6gB3/��"��Px5�3cl��<2�}�S�+Er�����шKj��|���'1�;7�YC,�Ƹt�x6��J˺q>c2Z���m'A���V���U�0�A����_z"$�kC�W+#DQ��qt�"�z�ׄ��@#V),m@9���Ξ�{�-{|�wBQb��������ڬ�����*��p��\��}m���᪁0��L=�8=�a�����U��k�m�5(�鷱ݣ]��8� ���t�42+/�*�v���!�X���l¦��Hd͊���.�1#gA�;�>ʛO���]�&V�򱡜:q��u9�f���j�J��w9/������������쐹�kk����7�W�����6Gږ�Np]	��d�2VEX΢R��P��<���|h\���^�n��n�}����B������ۘ�Eq��,��K\k-[��]���S&��`������yE�:�`]�w�����O=�_��U���;�0C��y�>��|�ɕ;5�Zg�B�1�c�̅m�w�����Ժh���s<���6t�ܕwдB�Μ�f*�N2g(��+%`�q<�T�T��AV�_,b��raI�%�UԿ!��Џ������|M���3un9n��{ޑ�_T�y(+Jx#{/7V�Ύn�vU��]�u�1��Ӽvj�n����W����ޫ�0���Aka�]ۍ٩��z�W91��}��s�%W�����L;G%ԧ�o�T���Gў��']�&w�(Xe �M󗫸���K�<��YE��m�tA��.�L�t��%3*e�L\ 5��3F�u�S�-J��X�N���t���,�젬�xD!;��5رf�|*��Dিcp�'�b�j*o��R�4��7�J�
|�T����� 9|y�Oy��B�dEޛ��W���u��j*&\���6=����]�$���L�2�Ucc��Ƹ�Fwu��C�S��Ǳv�o$��������n��
�{<Ƭ���0�e��>�Q]�=3�nF:':��|Î���rXL�-v��\�T��,�b�<$������W����fI�������p�y��M�J$.�U.'�6�_�e��v�B������5�oKlb:ַA�����3�y�.��ie���� �T%D�i\�x[��/$wZ
{�C��^
��X�R�2�Lh�$C,�T�Oh�ͽ�L�=��h���;C�����y^>���f�=�s�rЦEf���7 �ʖ��|�v�v7ٓ!6%3D�nm�����9t�ń_X�ݜێm}��"T�2�oX� ��6�󗫺�Qs)'�vVQ�jum��8D����:��x�D=� ��[�yx+w��띴�z�*tV!X�]J���Ɉ��Vn�38eK��0�T��!ńIW$%�+f�s�t72�fփL�܁JʘX��.��jt��[�`]\辊�N/a�7�Ra�5�4��ԙc^N�WYQ�\$��kb;w�åޠэ�u��^��P�;2DQk�l�I�B�h��+��6m�@�X��s;RK�Zlŋ���Bl���(�j��I�+i*h�7��(Ѧ
�/��YO)�av�X�(��FYn�+��p6h8mS�O*8�R`��dQܔ����&	����cÎ�rfV]d7>h����o��`�&��S����#(5�)۹ِ ���%�s*4�X
'>���'n�+WE��(<DĘ��h�a��"�w@e���M��[����F�oz���(��X� ��R"�BBb��]�]ɫ��.
�-�7wp��1ZhUAYR��vTnJ�h�����QL�\��@V���cM��Zҍ*�%��-*D5vԤċի�[kZ`-%�*
�V*��ܑnE�n��BSx���E�HDZK�*��h܈���%��*�+lZ�ʊ�k6KX�(ҺHiŒ����i��
%ZД�[Wa-���H�Y���f�J?��k�qg	:������bK:�׻)%�����!��GǾ��^��r�Ջ�ղ7���++��7�L_E���[TR�Py����g3��t4�X|����3E��[���G���r_�K�Ǥ�[���c-`����y¤vQNEڨ�Sݝ���i�d���z=��A���k�4��G�&�S�Z�y
��"�mb-�����e�Z���V�N�Ǻ_w<i�@�j���S��M_.��%�7�7����W�yr,ή�b�e�!L=��JGjih����O�~�Z{�A�<'�^�DG)���[�P������*Dwݭ�K7X��U�{y��8 i��a��Q�+!�z�<�w�W�m{���ݒ_�E&A�.7��0����MK��574�O?_';��[ɇ��yn�V*����o����f2������}��%x��wB�f�LN+����]�cS����^q+����w�Y��Z�݂����l{9k���Nh��WT�suN=�_�Zs�f1�x2���QQYsoy��j��<Ф<�qo�:�Pa59�
����zuo�eފUh9��T�+��@����p��4�6��$��#`L3D��j�,�k/�㖽����+��>�@�CY>�
��EY8�=���<Ad���z��	�VdIL6 �]`;22*+/�#����9��Lv.���D���X�߶�S�)dr��;W��L繆wcZ\����
�sfaoZ!V�k
�m�F:�������cՆ��ێ��\V�5�.�nf��
Y�:� �@.]�0#�Ge�G�x����Lmv�Պ���oC�u�l?Wv�,�����Y�L$��e�W�c;��n�7����`X����Ȟ�mf�Uƙw��i7`Z,X�����o��bxS��r81���s��{]��I�`��ϫTNkx�8h��VC�K���Q�y�Ze��`�=]�����W��7���y�V/�����b���%Mb!�e�Nǒ8�����3u�ˡ��*5iZ��;XUys���� �oa�Ih�c�O8�qrϽiN���L��(�e% �9�o�m��]V��'A�r�k�����[�@̥Vf���������a��"����j6��e�zg��cϸ� �W0�-�m�����1�aS�FqK�ۘ# ��"�LL�: "��ڝ��[p8��][i���.����c��n&�ς�/JS*����K�s�b�q���2H�Q����U���pϦ7�?
I��\JU���k`�Ei�	�TI���w�^��7�9�vk�s���]%�t�!��}�R�ޮ�����e�ۭP`������5E
��ݝ��Dҕ�Tf:n���f̗sZОp��FGR��R��_g%uz�}�a�3�q;c��*�9@Lً��uh3�L�O�v��S'�<��R�G<����6��7n�W՛a��'K8���r��	dW�5�Q!ϟ�0л���2-Iy����WԺ�!���h�t��t"a��G�t<Ƀ��w��^���i7�#x����>ہ5PTP��.G;�3�g�ݮ�#z����ί(Rἆ�͚ش�8�)��c�.&�j�V0dk��HYn�+�|ۇ�ڔ�O1�!�;@-Fh�]��`�&#:swmOb�y�5�Pb�n���T���ᗾtJ�gP���oB9�q7.b�� y��}�qc\��w��&Za�m�٭�±��Z)�
ͺ\�*����iN�R[t-�4�������C�P@�7X�!7uMB�D�9��b�J`�#٦�����(^V����'�&;Uc�P�b��b�L��i�w��f�.��Gxw8�/�(��P��a�S��f ��u���Ov�U��J"�7;{���{и�A������?L�O���r"��2��_�Y|�sW���8}�4���DD�+/(]���=2�RwkJ�6>��x��j1�5�����K�n$��֘������K���bX{�f�]����ᯮ4�|�
աJ���UJ��xk��7q׵B�Ws�RX�\�u��@���b�C��[����v5������֍'�[���F�Ef�l���%����"�4C["�4N��oOVϝ$V@һ�׷�����[(P�J��X��A3q�T<6�Gf�2�`�n�;��9�ي��sX�U9X����
~��ڬ@�ny�7�"kK���UƐ�[��m^2I�T�K�u���ީR� O(v��3�&=}�xs{Yʕ6̩��D��5�Eq��#0!���D��^ɋy.�Ʋ�v�����0bf�YiMŌ�(Ⱥۻ�F�s|�掅kk���`�AJ��U'
��]����Si�GiR*�u�����Cn6u�[���Xڙ�{]��6�Yە�����q?*}Ck-E���vQ�.�������
�( ��yJh�B�MrEK����]�5�wNbpܡ>�RS���4)�|t��Gr>q)5\�=�/3�,�׭��D��]�l ��q쬓LZ(:�w�P�F-����T��:^��̬������hn��"�v�����r�dNU����](k�R�+M�-;�&e���������g��BEt���fA{��<t%�a<�r^��&l{e2T�����9P�n-.��w1v���NvM�M��9Q���5��\3m�@�K�c-U�o�Z�(r�]!&%ԉG�^w��ڳёo��.�,��0s#���%8w57(��C~b���W+oD�ٖw��	j���$�i��E�/��7�Sۨ���.5E�N;F��9�R���!c�a��@��y�-��0��b��u���h�u��OrɈJ�%QX6�����s5U��$�H�RK�qܷ�k����~4���[�����Zܔ"��QE�ʉA`��wwp�/����-�Zc�	X�hZU�p��K��d�AċR�
ҫ!5%-p��cPs"["EU�UAUVJA1	H�r��4�"��$�h��+�p*
��$��\��G0�����ղ�)k3qq �B���f.���4��(9�R�"��S-EJF�����)m�mT�Ar�R��V�I(��+NX\��*����̕�B�RH���)��ю�g~Ĺ��8k��l�Q��^N�*V�}��ճ���Eߙ�n�«�E���=lm�W�<��_9 ��Qɉ/�b�vOA���*X!�(p��nq���9.xj@}6��E��խi��V8�3ĩ7���a9��GUoc��Q"=�t�;:�vli2M��	�������mg�o����2�a�Y�X�nR�ȓq��>��������b¨��C��l�I떣#i˕�Ȧ�g]=�j�Z�҂����]��ד..\���]Z��^X"��pFy[y�:Aq�����9����̩o2���86)���@|P��n�03c��Ģ�C�&뫉�b.�;j�Y}�A��J��uI���J�\�9���D�]�ԝL �%�,�����I�����u�{8�W��^��>��<�^z%�;�6(�L���N�n�o�¾�M���k%μ�!�0�{3rc��s�3��ѹ������{.Ҏٮ��yq��^s���w.�$=�w���n'������l\!g�q�y�~JQ��i��m6����ZТp�x���I���,'�� pT�ؕ燐��~����ܐXڤ�~q�?Y�>|�Q��V.��t�Yz���XḉVl�D�j�Ř���"��ᚨ��fy��m��KK�g�d��!x�҅�8^�I�n�,�0���h�o��Cx�࡛�`u�^ܩ��)��8���rN.�xh7~錓�T�>�-T��o��dT:�0w�Ll�NME�c�%�0�:�5��t�}�r�٦#�n��M�.<zKml�E�{�)'���J`�s��C�ڨS��0�Ⱦ�oK� 귷1���!ٰWhqș��s5�t�����^[ s�e�.bY��9�˭�XG��9��]=2�<.�5�6��S��z+Yɯ���Z���'gv�Y]/�u���^���:�a���[XL����OQ�#�ݾOko��{Cj�q�U�QݬLT27�5��W�l��'$0a�1W0:�wW'��w*�E�yW�NZ�y������.'ͺ�r�Yg����b��I�c�F.�Ǝie�B}uV�Hbu����Dj��8�\<��k)�U�W�]{SMb����y6m�d��Q��ⓞ}��ө���Ƀ'1X�Y}���)�F�b��Ȼ�{��tJ����,�}�D[]�]�*�����fj\]�s&la����������O�*�ۤh,�ҧ�&��y��;�1��r�>��f�k۔�"/8���N�XVȻ�|N����a-��}<���_g�������[���&����Om����L�:e��S����}}]q}�`���!g�k�=\�N��r�m>��."��:��1+j�����NlX��rW/40�ģ�i"4�
*1��Q2]UîIu>K8��@�/�EȘ��O�x�_v�֠��Q{���x�S5�ȎZK��tlgu���E;�]n�&��|;S���r~u�J{���~j6��p��EHA��p�����l쑷��g���nze���ՍNHy#t�v��	2����=������f�*��.����7����}�Ӡ{�㷽V�l]�S����t=�ݞ�~�Z�������,wI���n�ɳ|�eG6�&7U��l��%<�Z�e�}��>!Op�4�x'�'zX��\�<pK/��zZ9�mD��O�!7v���Y�D�Y9V�J��߲;A
{zx���0�wX;%j���
��1n� '�XU�A4�'���F�ݿ����q/�#,-u�\X��\䃍H�u%&jΔ���$��'�1h>0��)�W�G�J�1n7-t�X�<����g�e�qi`K�
�OA�(W1���a�Lk�K�����^^6�M����-�2��Z��=],4kKۉo�>����z.�ti��D�M<����Y�knGVd�s�c<6c%.qY�~L� �Ba��z3o<�vͬ���.��N��k܃�ʾIv۬�3��̕؏=Y�E��;�7�{�O<׾n��b+zj6ə����%� ��}[4�����|�U\�@��P*n;Ԓ�V7
�ȵ*)\n O����x4vb�u���S���&�������MĚ�u�2�]6��a˼���!@����K;��Wi�J��y��ƪ-iߥũ{H�����	�L���^�|_�{N��>D��II$�I=�J
  �P���}�䣰��}!&���)����p�4��̓�`Όy6�U@(A�KT��Ֆ(��аs	��Q�_�Q�]��zܝeb"�A��ͧY۫����k]<n�)\��bT�X��ud��h�g妦6�Mz�\�q�w7�l�(�����q�+z��  d}J(?�Aª��dJ-O����N�p����O���*���;�Sл���@�<=�:���i���x�H<\k�45��RcC���I�|�^�ZKX)O*�߳�����ɩ��u}�a�W̃��L@A�^o��ڝn|+��6}ҡQ�i$SW)~t�-+_��s!�]9���h�' b;�z'V��inO�� �(w������@�Kls��n[��x���?mf}�?�]�
  �ɣ�U�jsǂ�����L��a�iWu�r�ƞ��f=^O�%Ӫ���zh=���Cy��;4D�y3]��X���a��7uRC�R��Oi�0���Q����R�(���^�h��>.��
p\~�� �J�!?hթ;(�4<�ADa��H/i���݊�LV���C�2!wt��hF�)D�%�[U
�YQf���{n���r"����`����tO��r���S�3s�?��J�y���+Q�3�'S�}|x��$O�>���J��y/��"��z߰�:���JP��_�I�"  �~�y3MO��Cn����7N���Na���L]2G�(}��*�U��87��������b?_��'����T˶�Կ?'��|{��᷈g��%y���D=�
�Ϩ��v�C=��n����|��p�H����X/�a؃�>/��:9��梀��=��v$�`=~�ݘh�"�}*�ַ0��H�!�(/��H������H�
	t>`