BZh91AY&SYK��֤߀`q���"� ����b?�� �`0FfE!�bP�Q#mYdPd���F��PM������U��RV�AlSmi�R(�(����#,E�{�v֔kaa�hє���Z��Z[I���e��J�UZͭ�M"�
�-����;M0�f�%6д��m�c[U��lɭ����[m��f�5m�����{-�U��ų)#m*YZЖm�d����XBFm���cl�l�Fړf���m�2���6jV�m-�F)�������[f����$�Ԉ��  �j�n�m����1u�5�F��[����:tݫ\���wuˬ&�A�t��v�f��GT�����ͶصJ��Q����   s��gwul�S�z=���P�Sw�=v�*�Ç��U�*V��g��B�&�[�7U.�ڤ�ޏw�ZԡVr��J����/w�J�]��(�T�{f���l�36�e��M�6�͛�   ;��P�V̰��y{d�(�{�s˽�	T��{w��;,���^��
��^�缯ov���Lq�{��F���-��5%(�����{Y�*Vxn�]d:{{h�M���[6��!����   Ǿ*T�	�C��Z4�7���R������7<��ܪ�v��ݽU.�׏Wm4������u��s�i^�U'j�l�*oyW�J��,���m5��	M)�V��k>   X��[u�U*�-�b�vv�ܩ���H�sÏU
������[ov蔮���R�֭m�{�y�V��T���W��*�B����x
�ki[�g����&�q=l5K-���kLҕ�  �|)XU*w_W�������e�ԭ����u��m%w������L�<ʥ*������K��A=�<��J.{g�����Zׁ�R+MR��{V���U���kARV�Y�   �}�b�������c.�S��w�'e5H޽N��\�j�;��*�ޙ��7[nƩ*�5�BQu��.�$6��J�z��WZ�҇��� =©�RD�UVKJ�m��   G��֛���վ�m{� k��76Ͱ�Ž��kW���;�+� m{{g�U���{[�n�4�e�L�,P��3�  ��۲����7z l��N�UcL�uG ��{�;��n��(WC�F
=ݽ𮺢���*����l�USUL�6�����S�  ���Q�P�t법�;��7�7=��:מ��� ��-��л��z�.�����U7�M�CZ�{��P
��   S eJT�L	� �0L A��{F��))C�`&�@444i�EO�2U* �    �)*��    S�UR�   &R�#��Ѝ&OJ<���A�C�����?��Y�������ݤ�P�Y�d���d��Y�!�c7_M��������z�r�g�  ��f�c`�i��lm����cm��?������������d?�*�����6�,��;c��lccm������{cc��6߫86��� {ds������1��v6�y1�����Lm�;cz�0�������&�z��d�d =d6޲coY1��6Y��v��oY�m�&�z��Y1�� ���|�m�=� `���1�������c`޲0��m�d1�Y ���Y�6�� `���z�66Y�6��L`��q��@���L��q����cz��=���86���z��oY0���0zɰ��oY����7��c�L|�����^��u����W�r�r�Ĵ����!��&����m�T�ަ!v�	���=���U2�5f�R�R�(j�/s-��;��c��ԈI����;9o3y�
r�"�X���"*�k#Uy-�,ZبG������ ���#�G]��s����:�н{��K�аł�8Ù���LoEb-�`q�5SB\�7(�L�q ��������]���^mҽ ���e��Ency,%�E�գx����L�YZ�+��)e�;G6��cuv��km���IzSSʖsKT�8�6��f�c��P���Û-�f�����'�Aɲ�1��Ѡ]�44�������&�@ ��2����ۢ�ױ�)I�,:ġ�ˠ�L� z7_�@��J�Y�2J�`D�MR� z�^Cn7&�A7�I��%ۉ�n�I0�h�ܘ�ui��۹#�ƛ���5c��� HѠ)Q����9�*��5�٤S��J���-����}�3y�MM=*�(����fQ�i\���$;F��Q���acI&��T.��%�y�Iuqk)$�u�!`RE:��l�w<���ȳ2����x��hqj�W����ڧS+	���g��4m6Z�S�m�3A�(*i���]��zC�Be]0��2��I�j����ŖiG�)b�v�Żw(bb�^m��(nJ�a��8�kX�g&�s,2VdF�T�z��H0�r��Mk���]���@����(�̽}�
c��Ѷ�g|,0�9e��v���wE�r��\���%:�mH�$h]00����!��ݭc�6��lMf���Ik j�(���ʈ��(��m��̔㬖LM���2�ҳ�h��6��ܨ��P�,�� ��*Ƃ�6[5t��M�-mc�n�n�ӭ�#6(�T�:ʀ�EX�Z-��!��\���ڸ���v ��-*�l	�ҕ�oJ�`�4+V�,ײ�=�3�`Vb��`�ݛ��������Vh�f�J��Hw#i�:���lݏ5�-*�^�!�� �x��um�#2�72���2a�wiLʹ �[�Low�`���i�a#.��5A���1mʲ�[���f��I�H�<h����Y�Ùu�K�5b	d���6�u��goC!��kn���ٗlT���ͤq�`����]�S� �S�E%�6���m�w�B `'�խ�4��D��v�f����H�&u���Xw9�/�3�%��U	Yu�\�2i��[x�Rܴ��VH���}�Eic^)*��u6�m�e���@M"��n�HP�'Ʈ�&L�i��漲���b��2�;�<�e6����E�WI�����f��ڑ������n��I)Q�ӕ6
'BD��ܛ��Az�%�%4���kT6��t�F�髊#CV�=7z0)�vM�k�Q�����l�:,��YΙ7+kV��]	�T�9�
�U޻ѹ���m6�J�#9ZV,z���]m=����~j�&���1�RK����<�r�V:�V��`�d��h�3�;K�L�+�ʧ���ivi=xwE�B���a��[ƵX�+ve6�k����
����:�ngRW*��O�I��9yePс�+�k%���Ƽ=��b8����7 �T*=��ш�SqeM?�AڭC^��j��nK0�Y���MܣF5��e!5��qm�`4�a�2=�˸F��=�r1gu�ݬ[n�f��Q6���eD������{TM�լ:�-lښ%<��֌�W?mK�TQҫ+rY��vF�z�P�8f+ͧ�?AX�$�w+&lgd<�G1�+@���7(Rt�u�&۾�\��'�֊�v%�zm�����V3��-$qmi��ٳ�E��n�K{���`�4�12D�fE+Xx=�)�){{���M�i4a�YK+c�c���m�.�-*L7S߻O],�	b�he�V0kx�Z�qf�b���㿢ɍQx�;E��a�HyW���Y�p�b�ChoM�Z��o!*R
����
�c5Q2:�U4%�~�Z<�W�h|3��F��v�*-�L-N�4�Ѷ&e��F<�3%�����`"cֶaإ��y��Е�+��W�am]��HU$�e�3��Q	@��8.��l�
I�&m#f�6"��ٻ{e�Tn����2��l2�{��C��c�Ň�nV�GPa���7o�\U4awW����B��f���J�bv��v�KFA5��pi��t,���RyBK�)�A'I���� $R(1X�m�zR���[����T�˳r��X�����[�z���Xi��J3�1[�V輗O+r����g,呀e;B#����db�A^�����&� M�)��*m��8��\*���dr�*f�V�W�X���f�֋��r�?���5�ض�S�,n���l�w�ʢ�q����e֨s1��'u�<p�,1��`�[�U�f�W5fM���%�R�Nn�8�Mmԫ�5R�"�CX�ܼB�����i��X;�8Һ6)�*�&f7�:[�M9y.,:Qj]#��f�o.����De��(3U�8*{�Yע�+sh$�v������\׸�M���2�[���R�����c"&��/�����[��b��;or�2�(�U�eRWX*Q1k�3
*�r� ֚;�ǎn�&a֫���Ek�QH�AG����uy� ����YUv���Hb�Xƒl�&LQ���A#cl^�X�iYx#-=n�V�v�eB���l�l��VQͫ��}k"�����1�Сw#�9���V{k3n�	hꂬ`yWQ��۠v�U)D(Sb�-�^�n�9YCa;���I6���S\�.:tdː�*�e��u�4T"h~vN�ء����d��ы-��D�R������*Th�!9	o`� /��ӹF���l�#&�%x)47�m�Fh��4o"k��?��ʸ��a�S��.�jF*[{�x4�^4�i$)x�ZS�,���e1��b�# ��2-��7m�S[���1Z��=���գbO���*��LD��c!Լ.���#�7�t��d�q]�7,$Х6�ȡkK��ej�tv�6�vJ��b�c�5�u`� 7L��&f��$�9�]���m�wX2��c�i�X�t�7�E���%�ͮ�o��W�ݒ�]C�d�1fRv��'o,�CX��N��֔���ۧ�#W��n=o[N'[�f�Ym�\W�� ���w-��e�H�c`��zmTbq�[����.]X���DᳱىVq�Ή8-��Z֩H��ݺY�A�ތ�*"蓘ڻF���f㊝c�opl"֧��Q�vU�o`Ԗ��XR��Sjc-���uB��54#�.�Ӕ����i�e�j�V���VAON���!;B�<5.��Q��C),i�kD8ͣ��z�D4�.  R�^��iT��b9F�@�-�͕0E6�	���+b�F�T�YuY�5�#��LXxBDz���<PU[�[\Z�oR��bֽ6�C5K�59�\ ���=ll��b�A��2+����4P�8qۂ�'b�ݳ�Gj�SJ�xk(�'T�eL�Gt�x�b9S�13u`ծ��4��U�̄��4��NLte�J0�e�2B}������c2�Ѻ/6Q��f�㬉6�g���\YM����J���=w
&����jJu�KpK)�W7m��欂��N�^,#Dqڸ�$&�6�;���&��g$HVkS�61��<�'e��-R�f�A��p\Ƣa��%����Y���-�V�"�=6n�h[d�*�u.l*�а�]���J�Tx�ʭ��n=� ssـ\�&�5SN1X���	K�H9�[y���*�'@i�z�B���/e�Q���WlC �N�3r�3�&ᨪ��@LV����Y5�TPN�ׅl)j:���`�Нa��7�V͓��p�X]�ZLV*��!����/ ��Զ��40�ي6C�+j����t���Xw\+#�4�x���d�-�i�*GV�l5��;zv�F�sp`N�f�����^^�Sۚu�#��Si�{�z
[�-�wF�S�r,����v��br�h�k)ĝ4�U&Zkf�mZEZ�p�I������x6����d�PŶ75�e�0u֪�,��7	6r�j�͹W6����j��%��h��[���u�CP�l��&eQۥ�D����D!z�nA��'�{0�m��܄�5zk��+��2[{���旗��=i]җs��*9j6��# VV�lX��:�h+m����ܶ���[����ǲ݊�Q�I���oX�vT��u
U5Hӊ����e0����}�2�;2��9�K�&�Ʀ�R!f�B�މ��Ò<�Bnaq*�,�e�4�a�,b���׺�v�"���ͤ�O���@�������@�e���g$�i�lhQ�s%f�HM
 1T���Q�ǵ����S!�Í�S�Ӊv<��ش������^#k1e�eJ�`*�1��$L�H��f+�VF����z^�)����G^F��6][�Ab�R��(^l�Puy��]Y����U'6�)g�:3(0`:��p�Y@�)�c������[ٯn^šd��1u"u�nnn��(����M�\R�{#(�sh��Dӷ�H�"!0nި]�y�	�%a6���t��#ۊV�x��-��bo^��ڶ��C�7��	V�ۏ�v�yY�H����O�*T sz�kΞ�Y":�(�]7���@��ҩ�F�"�2
��G��@tKQBX�V���?���F�9�E��Kp���PZdSF��5a�F< ��,�L����ǹX�n`^J{*!ԕ�dz�o6Ҧ�-o�l�2:�4;��/6Q"��U��mXl��J�	Lt�z�#y6#w�ۚX�mY����+J«u�4��m��c`�ed3p�=�Vʌ��&�ଅ��*1AhMۍ�jh��S�7ʕ!�z1fV���Y���gRy}f���<~�]A��z�e�kn���F^�hR�y��c�.U�R����q�F��(lӌ�Ŭj�$��zݒʼ�YLx`�[��ޛ��d�B�n�&�Y2Dҍ���bٔi��o6���a��e`��_�P�����9t�뭥�� X����w ��&� m��{��T6�۵�]gR����ɻP(��&��^V�EMO(l�,��JZ�h��
�����A��z�g`��nZ��SB��T+%�	�%"ݛ�HE`<�6�j[�7�@Y��OF��BIQJ�K(�c�:G!�3)c����x'�RY5�T�r��P���{flFP�H��5Z�%2���횘��X�^ǫu�h]����,��JR�7������
�)���s�Q|U*V��U��8�Hî,������P��Y�T�ã��0�3�u�� �tiM6�����B�V��2�F�hVh�"�¦+c����M셡��Q-�ڲ�m*]c��K�׍�Ֆ�'l³v�R�0)%��X��JZ�ۛ�e]�:�bR���9Y�͊�PVj�ib�fa���m�U�/�1ư����[�Df��I�!�ia*���d� pn~,]1I�t0=TH�MIiY�4�b��jc\ȱ�,0ŗ0AI5��4D�4㤣�i
)7MmkW�Ǒ(�=�ۻ��7�7��a���p:��4R� �B��M�i,��6����
�1����Kde�Yy�%G4��%ne'hVFws�`E+_������RiP��U��֖ڋt����G{{Q���xv�ьa��]�`B]E��-	��[L������3b�7o\�nV~�S��0*����Y�����2��Y	 ��u3�RZ�-�3+)j�c2,)���I�r�Ӹ��� i��1�F�-�Ưk0^�锅]`h�kP4�/6�
fbJ�k��Mi�y.8A�u,�n���l��BlY�
�BG�nYNݬ����K�L��U��|�T�6���[�j������L�%���gv�B6	k@5%�dײ�ThS���)�f�b[YX]�D��%{ *ڡGښ�,�l.lb��s[�Cr:�m����x���QLܵ��@�����: ��)S@��8�]�Y1��f�}�������
e�U�P��Ѫ�]H�[b��t5���M�������S	L�%�c0%j^`��k�5i��C�{��#�m���\�������N������*ye��J2�20�0�{���mnp;�˷~� �%ݛG:!�K2����	+*�M��0���/?J�.�<�M���/r��Vrh/n�̽�@��V֛݂�[��y�5HI����$eh���!X�k���_J�V���$جзr-���j���2�5�Lవ=�2^�J���[��ҙ�ܧd!�#m�kq�*�j�c�B��.m�q��(h�%�Յ�ݕrV��1������=t2�XV�%��3;PR�=�6x��F��YW׀F)(p�Ա[�<^�F�m���B�ь�j��[���OgpY|��Q}�}�Z����;�R{���JV^`Qǎ\�W��m"�ze�:�֊T�K�2�']���`�R欥0#�1h��Wsvri$�v�����i3��#�tb=}��~��(���[W�aǭ���ׇ/'�un��6��d�S0�{�b@�ne�r�Jf��X�e��E�*���jƇ.U�y1��nLeRyd�Å3R����^�H+{.�m��S
��x R��ǈHs��I33i;��̻#f�Kgx�G+�;�%eo_ӲcPm��v)үXM�c�Y\uô�C��T��������<ߠ��`�Ҽ+�0=�f�g�w����h)��R�n��.}6ڦv �杒*m�g%�NQ�/{	�8"Ԑ���f��v�՘�V��h�:y�7�z\�J��r�]6���?"�AA@��өV��|h^d��U�q��^�}T�������EC���� j}y�V �9o�N(�o(���W��*=2�ޣ%�ד*V���!��}��_>USq�6�\!�r[���(���T��3��K|y]Seeo+�r�Jf7[��y���R�M�5ʚ|+2��z]ˈ��m'G�����ACڱ�o:��]*�������E(홢�!�:3t�Ͳ��7�ޥW�i\�$��;;t�*�B��v���%�!��J�f<��ݲ2
ֶ�����s�x�V@��v��zn�a��|��dtQ6țr�P�w��\pM�E��5΃�2�r�P�Jd�M�2��}ϩe˦%7e��nG�376��{!j�>�x3��9J�t	���#����LrT�� �ENElB�[K��-�[�n�=-J���$ݝf�t��Ќb�婭.�j���ֵ;�>P�w�ŝ}{#W��VojR�7F(QEI�wZ�3����Mg*�m�.C�D^Q��8��S��C���@=�ٖ��[�o-�Ǎ�ۜrV ��L#e���3�n��A�bU�[�C���Z��U�4�{H�;����!�7B�B!ң��N�'vS]��5�����9����C���,���k��Mi����]0b��O�i�ݩq���)�;G�T� �ʾJ�#
(Y��T��.��o5,!��ɝH%�r���HHt��W6�����L�ע�m�N��A�R�7n=�0k$a�w��i-7M��ҝ���L�%E<�X�<k_MQ�:w��+^o�3AuMz���jX�5���E�����tY�/y�v�s{��S�ҵ���a��I�Wtifpӗ]Ͱ��pk��H������X�Yb�%���Z^�mMT;v�kaZ��9��U�����.�vK�ɺ�:Л;6�h�2Uו�],���M�`akX��Mb�q��K#��]�{7�k�Xr�5*�H�\��d��i�$�]��y���Ĝ1�HY;bp�hg�c��GjI[Cc�JwD��V�ø�;��o�H�-�)��5�����t�y4(S�h�>K7��`L9,�v�Y�8z��X;8�e@̬u)^r�LB�=&,�\3��j6n�`�'s�%�rV���@���ĪH_p�ث�����_Wm0�:�`�i�W�T�:Y��N��ƵP8�,K��O�\�6%�ek�l�����s	�X �-ևY�����i�A���&���u�������+ ��,�b�]sF�M-�Eئ#ݗZVv卙��z�r2ns1�;�Nfuv��#"ڿ���ߣ㵭�0j0�ϋ{έ<���%Y��o^��U��-Y ͈v��=���5V���=� <�]����q�Io]k�;N6!�z��31�d�U�����M��������V�t)�rG��<Y�M�R�t�U��`"{9���3h _u ����"��IWGE`��4��g ��zn��&�j]o]���v�@0!����-�٣��i]u� �^���B�3����S��:�H^𧜱>٢���r]��Xe��E�2omnIW�,S�Bʥ§�ۀ!�Y��k2���5�.��O0u+�%a�enc7{�F$�je������A]���D���%�3�.��\���ue	��VV�ǖt=Imrf�쁅���ȝ����әl�㳨u��'���k/�;�S��'�����X��ND���v��l1���u�YG:)����+�n4�64b�<�N�{\iJ�xR�Ps�'r�k[�$����n���i�r��Y�Rwr2l7΍v�Ś�F���Q�b��r�U��F��S�&"'8�&vs&��4�뺱�E3����b�j�v�y�POm����˭k9zM3�]vܔG�8\Jb�.� �S��G��$n�e*�¦/��c�r�����²��tj�Z���(�o��yڦ�=�x@�+�hAPo�ɛ�c�iH�_kTҲ�5Ԑ��^�o�b�a]h'fZ����]urƇ4Сk��+X����Hط2b��T.�\�a^�ގ�>%���/N�yiR��o2o2a�O� �x!������Y�|`V�E<߬K|,s�u�y�����wv.��n��})�Ĩ�l���=���f��]�`�l�%Ps�� �JV�.��s����y�͇�CaƇ]�޳�����V���)�װ��ܯ�3R�.f��#�9�q<dL�uQ��l/�2����rARcW��7�����)�7]A[��LH����'X�û^�S�\���R�EЌҏ�)��_MC{+�ֵ�&Ξ��fm��	z�7��#���5s�D@���' ����v]�<��֧�ř�L��:���n[���ّn� g�
x�3es�Rx����⭇��h,�V$���YqWϯ�����udӧ����۝�Tt�w*��r��Q��.����LUz��Ec�7v��ý�0��-����^�7����J;�s��GP.�8�����G�e֚�굫z<��?EC7���ʥ'A]������9�Ij�PtδhVH�aQ@��ݵ՜tiD7� ��	���-�Mئ]|;���Vr� �4�st�/Q�\7+9��<���E:�}ʝjVθn�[#������ �4���G����WtO���:���]�L`��i���wM���&E_�:P�E��Tx��Ȇ�yZ0��y2�`AL���(�!�3&�z1qq.T�tIt��Z�"l�p�Ko	��^̬��T��N@[g�ȷ��)sF�Y�M�[Z��x��uQ�/J�v��&�vr�e	*9sfF+*�GsUovp�-��gm���cX��@�م�@!���޾�f�ѓ�7�s�)T���.۟�2��P�9uZ��&c�X3�\���&<�Wy�гBb�̓�B��j�!�Wl�N�i��2q�%W�;�VQ�KvTc�"���)Eش�]@�}[À����:j�3 ��X��09�L8���~MLWQ�:l���F�\'oN_n�ギ�fLfqZ
l���eDR.]ؕ�Cj��v��D���tje��͢�/Kѱ��Ñ����|��xR'O<:�o��d�*��6f�MJ}t�2ُ�mZ�}qڡXr�ûv�4�j�Fɒ'�gU����jV*`�y�F_X�tf=u��7�l�ZN���2�S���C5�������R	dS����x�3d�X0��/� �ۗ�G*`�F�uX��]8S5�����]�Y�����!�r��i�/\/X�1�0��D�W+��,�<^vmѺ�/�7y>�b�%%�|�BX�%��	X)��՘�M�7�\�J��ݴi�\�=u�;��,̥����v�õ��Ą2"�9��WۺQ(�	��E����o�-�o��t���7	��fc��B����Y�'m�.�HP��a�C[���XY�[�[��z�K��(보��y=���������kc}�2خ,�I�#�L���*�[�9��|q$y�~�U ���[�6�^�V<��v�K�Wav��m��6�6"�)����p��ۺ|����������x"�5��f�}#[6Y�YBD%�r��\܎v��m�^��󱮲;uų�ȨY�;f��'CS�i|��+�Ħ�j�<'�Pp\�Fm�\�k�&����Gs�m��S��혮��8Fq.+L�} �}��݃$7�&p�0nJ��ޭ��Z����V�rKSY��-�Yd�-r�b�lnk��yvu7�.�U3�/�T����)���m��r��x�e'��Q��w���^�N�h�, ȫwA�3-Q�KX�38�d����9RM]�!�oP0�f:&����S:�*���F���w��8�V����n������Ք‑��WVZ�aͽ�Q ��*E]{�N����Z�(?N�zT���F�p��e��f���E%|Mp.�3u�v��ٔ�pF�R�5���\s^ՉK6�y����-�n����?����B�fr���eY�7^��]��-WS ��w��Ne��`+��%�y���O>W[DZ�B�N�x����z+'{��u�WK ?&����[��ĳy	��iQ��ga��̺]F���1@�B��1e�͕;{)T������*�]�Sq���CV��#�U��<���n9ӥiP�ʴ���H�ᵟ����e˘o�	Į��U>H����x�BN�Ҿef���%y��.�nGo[��K�ܓWL;�`ێ[��	W�F�*��f]�"�x�$L�7;2h�� ��7$9�i]��
hw�k$��p[E��%�q9�"wF�c�(�hx�����na�%�N뛛�Φw;����\M֫�=\�]�^붠Vecy)"5��K]JX����J��g�U�5P���j>�SEa4�7Q�DM6AW
'��&e��m����F$f�R����:�`���X�KZ�N��D�`0�&%κ�'O_���S�7w{��q��MW%��16�۸sf��)�K�u��U4-�Ph�����LL�\�f.B\j=��ɳw�}l���le���y+�oo0Vj^���
ن���+���Q_V�m�����;�b����<Ѻ���YdX���\�Ǿ���Nn]���Pz�u�DzN�p�yl�ȭ�KGׇ�At����dg:`�: [��;�-��P޼\�m5)wmVz��	֎)%�z���}�˥��V��P��2]�.����$���Nw�[Bl�c�
&����a�UGE�\�CV5IV 8q��{.96�e\4�u^��ni1�k�we�䲶)�f��hfM�m^������F�:���m�w:�@9�ޗ;�'��J�J]L@[�t�ӧ+�ܬ��:�u�5����a�zV����U�H��cw���|¾7�j�R]O�bw����(E��h�)��h{�	ٷ�7\��R�U\��J��K�c�qn�8�(�d�*��I���<"���d�\�:��;d���npZ���{�
\Z�)]Y���6\ږΐ��-l{l�����P�Gu:Uˎ�+w'W����Gp������e����YO�K�ނ`��a�]t(%A��w#/��U�3���p<��Ӗ_u�mt��g�$��M�N0[Vd��K;[�H�:�.��[�uhj�p]S_2K��+��!�)���*Y�7��*�H 핐N��gw{lju�)��ŧ
s�ƪCŚ��u�f����mF��ZZ�,p�r��@��}M cT�T�V��4w+Y��wٙ�$۫q��-��\(��p&���x�N����9�J��%}%;*��d�?Ǒ��Q��١���(����+A��V|E-�D�1�6u�r/����&�WgL���Q�33``H��7��8E�+/6��(��J�(,���2�㔋A_yj�!��y��El�}Sw1���\Mt�]le���)��HG��ٰᖯb�� w-U��*A|�+��"�hڛ�0y��SGQ[�ܦv��U�+���4�H^�e�J�#J.�(K�4%ձ�(�]�F��RT��8]C�%�Y�9��[�0]^���0��뮌�P�4��Õ4�n�S6�F7�����Xb}��Op�]]%���͗,G���u5֦_��)�N�.r�Wa��wL^�t��:ne܉��V42��Q��T�
B7y�=bIWS9�9�LnD	Ԛ�M֫��\h7,K ]ۙrk�NPݣ��we0�k��j�L��72� ���`nZ�-�8ٚ/Y�;���sy�[����J3�ĩ�+ege癏�ۺ�9a����V�w�	��#"x;�oq�1�6�yn���hѐ�e�x��VS�wη�=&��pM�Y���J����1�o)퐦��;@M����Y�qR�IF�+lֺ���}����*cEr�#�[n�F��wB �1;74�>����0`L��@k��Obi�m�8-�{
$�f~Q�*RdV�*f�0e���į#Ƭ5�{f�����(�q3e)Ѯ��]+����=y�@�Umm��|��Ajs�,UH�lJ��V���um����ڕ�!��
�-��&�H9�"�z7גցL���T5�8�Y}2���m��]�!�V�\XH�k�C�o7���c��8ܧO�P��ȃ\4�.�.��@))=�Gm�t��XFh!�r�2�@ڑw�<k8Y(�u�	㯯�Y8+��#q�ro��Qhzx]b����ږ�%S��&j»^�/���w��&�@1�D�Os]�����){B��,�^��'*���R�\E9�WW*j����p ��$��k/���iSO��;#�;9+ܡ:�ns��b�:v�\A<��zWjЊ�|��*ay�=ٴ�Q�i�/Ei=��\\,�S��N��{���/�^`ls3�-��������4
9z�v��2gGh+��f���;���oF�-��1,��y�VB�exzP����Z�"5���Ý�CQ'�N�k:�X���v��$���"���LJ��ɱbU���م��
��f�4@�J�9�`ʇ��вxq�B�]��Q�C�u�+������¥�)ʢ�%���{��=u~�d7����K`��e#=s6�YGh�J�����Kd��]b��}�^�k���˿��wU�\L*����\�m�+(S�d=�I��o���]�\k+[��c�Zj�ˏn�)�1킰ŏ�Ԋn��뛯��T2��[�8F넒.��zܐ,i����m�wo����JF� �7M�y4S��[[��� ��Q�ja�Pd�.�'����P$h6��5�)(��Mh9-������w�}<��{��_��_W��l�z���{������ߟ2�_��Na����+f���&�M#p�ţ.I}���Wa���*v��&��b�sƷN�٩�����vS�G���Olyi����JNP�b��b�����B��erN��n���^���8�\��b��,�T��t	wV��+�#�׃Zj��F'���&PX���{��a_WwW�+�6"��QHf�C76�+�yx:�g��`���޺ew�]N�^����n�i�����(p��Zeulڭ�}�,U�Q��}�\P_��#S��בt�B�V�K�y*�O�"��/D��0XS#�*�t�kk8G��UǷm��t8�����kAܗ����iX���N�}}��m5,�F���������c. ,�ڤ]��&F+E=�v�j�.�ZU:糩U���(!��0��r�2H��a�rG���0H7�f �Yф鍫T�n�� �]�m�r��s�ډ�Q���{p;%�޴�a�y��0o��b���+�A�����m�g��V�e�ݳ��-��YT��uy�M|��@Td4�F;՜)Mw{w2��ۋ(etyJ���^��Bzh;�%��K�I.�!���Vj�`X$�?7�)7:�\���|��fItq��9�,���J���W�R�ic��Lފ+��&,c�@[�{{�kib���-'L,�n�o7���mu��6�T3F����&���KN����ll[vx冮漅��wO(�:���2
��P[ṵ�D�s���h�ɭR���{t��t�ս�^��I�Zr�0�ȑ��AD9�;;��vN)+��o�����.���kd�8J�����].���MUę�}w�JR����c�`�8>��}|ҵ��1*�WNoU�#H�o3A�2��t��\����9�ǲ��h��qiѹ���o�&��&������.��Û��cj�p�Z]�c�ۨn�.�{�X�J	WX�1��_k�i�#���d����&CV���� �lR9�n(owJP���#�����mu�|*��p0(#�Fpƒ�M�6���FV�7,�"�Z;����2.�Twn�������q�b��ᇹ�u�;M�xX��3Dt���(�k
���^�u!V�Rs�'�1/1�g(�.�6���@AH���w:��]�tɅłJ�����Z�q ��:+o6��!���Q���J*�/�Mpyٽ���2�Ѷ�;tCF�|ƽ|�9m"փKGuDow>{�lwN�>ȳ��\YD���a�vsS{�*�,�"�Ww�������7��<��.�fm�`d!��Ru���p�����ؙ�۳I�d��}���rM��Y}}�0A��{���C�kb*XT���O�53f�&�7xD3��P�#���a�/P�����d��Xt�:�>�)�nd�{ǩ���m��O�@�ń薂����%Sr�?��>�G�>�Tڝ���n��ޮb!$�{	�81l��W�F��x�ʁ@���S'V��HF*&YV��PҺT*�r��J0�2P�Tƪ���Ʌs�|j&�/���RN���td3�^RF�;�#y}�c���
Rމ��7���u+Uj�&�GL�a�����uhu������=k�)M�WL]���UհK��2��q���*�P�0=�Z�"�|W,c��,;Ζ��kkK�mDo'8�L����L4_�����2�0�Z���S����ck�������I��^��� h%��dt���*rE���4.Ч
��0a��iź��X�bљk3��1Fp��E�NO@-�w���9Rs���oDt�'��NM�r��X�a�wc�J�0�p�NkVj�:Xc�T��f�xD�@���giGz供��bhFi�R���b].7�q"�NF��V��yIf�!6��`mM{��܃3�,����bC�A�1�;U�ʚ���Ѐ���@�k� �e^�;�c�
��h�V��6_�c�uq�֦�om�;d��<��r�
}�YWQ"��Uݺ�48��������!ƶ�nS���ƍ3�#O<�C]�S��s�R��&^�Bf�{�A-y��cm\b�ӣ2������msBc.�+��6���o~x����Z�`����"���"�40�m��]�gF!����n]�K��䜫�Z���;�ܶ��2���S��:x|H�o67κ庵�I�vu��+���e�M���������)��u��᏷)
�W���H�{#���v�#*�!�R�7˴�Q���wpf�3�EfÊ�9�4�J��ژ��+	R�ˣA�]�ܹ���u���n��2�LUxE[�<����\=-�nM���g�ڨ�8;�3��^]�s��I�f�g^R���Ŷ�a+�Ĩ�3����Y��̜�gb�6Nl!W�թ� ��a�l�Cl4�[F*�e`���J#i�6gd���i�*���'�EQ��e��%l7J��[�������nV�
��vF9h����e_g��}��ȏ�^�㭵�����!
�:�됫�kؗp��^2�!u,ut�r��bxC�삔�X�X�����f��:<,���%�5qM5�`��3�������P۷��:f���Οp�3dݭͅ��
p��L��^���c��C�Y݆Z�k�3|fq��j){�u�%�m�w\0�d4�q��l�KTŗ��u@���qp�{y<%9GaK��0�~]�ҭ���r�8L�iRM�r��t�q������mY��6�9��qɝ�a}a�5��[��l{N�ʾ#-��iA�P���(
�t�C�)M(���4������x���R#�i�'��^�Ff�p`GtC��]��rh.I��*�f�xxv�����ܾ�V����<�2_4�n��]����m�.�ho$j��M��'z���9A�J��e��j��qɗM������V6y]�-J�v�1l��7�����ꂧ,T�8���s:F�GV�S]s%h�2f��"��l`J���7��$<:�P�*�U�N�����qt�Wo%�GrD89��p�mC�:��b��򘡱
)]Z���ڊe�4�G(hν���ݒ�%&-�}ZJ�-pC``S"�����X�
��u�5!g�VH
�[A82�ܬЭf�|ʅgb0��XƊ�y.w9�NwV���� .D�Q:�kQ;��ͫx�ɣ&R���P�_��c3�tY��n�`\#{���堬з�9�Z����p�v`��o�m�\��z�]�Q�QL���E��jw"��j��A2�y��*����i3����9z�zC���9�.��׹Ի!��+��J׉H d�'IQ��Zq 
Jݏ:��ǧbE�̲c֍�F%�A��E�N�Z���pM4?^�����I��F�k�'Y���U����AЍ/���թ�ť�ޚ�ں�K�U�T}w��[[r�AM���wf
�ɡ��!\�:��6�c����\F�ӛW�z�q/U�
[1i2nPj.�Q5�N�K�'83���BVɗ���G;R4�w�}�x7f��o\�[��m�V)m��*��,]��Z�2����SB����S����v�]�K�)锞�#^��D	L8��C5ğU�3K�`�P�MU���q�^�k�Y����ϡyv�����VB\P��ZF ���G�鎃�q���,��,>P.�V�1\��1K�sF��{%>q\=D����Ø.F-���x[s�;ia�6����0�$�)-�*�h��k���4��-���S���٨��7���Z�e�Vh�,�/a��C�_=���t�,ɝV.;��wD��=w�I.]6���9޹�'����lE�7M�� $�ح�����+atv���X�e�&6Ů�}cӞ��5��;2mu]�LL�Ԧp�Mrݠ�k�:��cZ��w9-�����S�w���g/�Isub�Z9;]���ʱȋ��c��S�t)��ފ�z��ȶ���Y(:�N ��;��{�V�a����!Q�)�[Z��OcK�����m�!��¹kⰰK�{��wgU�� Go)�+��i�t�X5ߺ��D�F�ۭW�qJ�C��]b�r�w��O�K�r��c��$3W�On���u�5����1:I�\�M�Ke��'5Vn������"��ʡ;�A;K	�1;�,�̱��9�ആ�t�z��QO��dOһ��z6��ͷ+�l9B�gn3�Y�{�;�V�v�Ԣ��fm�U��Jv�5��n�a�Zc��V��ed�\�=��A�3�Jm�9K�浵����;p�+"�@v4O\C���[8�lAxb�@v�	��ma��֩؏V9��x�x�k���u�ѤV��è��,���a١�Y���T��E��}]Ih9�g�VU���p.���-l�h�ږ*/��!(�ݨV䔺w\�fZ��\)Ӏ�͒�;g6��$�	��Z�n��;���7��mvN����K�m�QvO�f^B�t]X�+�������y���:�r�6���4�[s�U1�\�ط��U�}���9��5�#�vj�p;�h���xZ4�Q�hH'6�+��,���6�A��o ��e̮�u���݆(�We�9��Z�xd��Ǫ�%�����5�ه)����7��u��:���v�phAI,'����kzɘ*�u��f��
p�	�-��b_�N�����Z\�KeI}*$�u�`���-�{kEg[O��$(��M�{�R����n^�qT�y�'t!,"���I�y�vE���-ɽ�x�⾌@V��5 ��c�{ǔ�R�7��Wr<�H"8�*�mn��J:����b��r�M[��m�	��i��2��)wu�(F��xlګ�HBp�+*og\L�JQ��rwW,�xT Hs���ldA��6��5�O��Z�ޢ�~�m
jGW>�W'(0f�e;g.gXo%;u4,|�aq;��Q�,x�u:��T���$뵈`E����ՓS����Pu����H��w s^��k�wPEf�593G�i��"���
�;��f�wy\U
6�70���Q��oe]�-b׏u��B�0Q�T<�i�JOZ�tp�����r�}�e����q�����/��z�ہt�A��%�\��}*]�Huf�j�3���f�i��frI���a. S.�{9�y��b�vs5Zj�P���̻o:�v��_�;�Q�F���m����7�ו/k���hAz(�-&qWq��o��d�����9�8! ��V՜���}֤�A�)����w0�7�a=Ѫ�T�P����y�ߢ�I�4��k �OT�v�
]�a�T�=u5�2��'p-�k4z/����>}�XU�	b-��'AG�
�|��5�:.[�-!��n��L���>!W�����4V��!�;<��nrN_d�L�b�_V��Aٓfj���������/#���iPW���sy_v����t��t6�f�s@��B��0-���4,8�=�G4��3.֡Ĉ'X�JL;��sEm����˰�������e`�浬)��G�T5��9��	����X��%@�9ӆ�A��,V(xk�m�꺺�@f�H�lHtB-��'dɽ�\P�&(B���MJ��ړ,��}�yV�M��l7KXj-T���j;�)�t�m����T�R�G�'^Lpf,ã�B1���JBY�/7�m�֎���WT��6	��:�`=O,�l��܋������~��z��m�L	h�ػ�j�u��4�0�v��ηR>��P7�+C0�s��A��֖&�]$s4�B���I�&wk�X�͈,n�Ks^In=��Νm]d�Q:\�!nI�{FW,j>�Fke��YV�v�W���v��.���QS��$�<"na�.��P4�re���FmӗC��B{a�.�.�]��)BѢyR����u]au8���5oV�	;3V;um��f�Qۀ��.Sw���.]ry�=e�v�5���F��5팈n��)H1[�BI�έR�n�)�����%�{���S��d��:闢�'ca�m�S��<�o��*�#�++c�%J�4b(����8�{)1YVf�x����K�..�n�d;�(��v�y��������EC[���IQyyx�x��u0�����W��w����3�d�öb�Z���i�.��[������D�""�+5"����+r��Zt"��&W
Q6p�;@=�&:��b��;$��_m�8�f������\��6����+*�]C�2�\���gw4�M���uӴ�*��}��nu�@4�2)�kkh�Xl�9oj�V��ҩ�8�]�ԟu��aђ��Ic�9]�Tu������o��	�>b����2�i��ޠ�������R��T�v͊���[]l[����WV��zL���rmJ2>�,j�v62�ڲ�Ӗ��Р-��9Y͝c<A�X�^
�6�\�т�f���J<�|%f�7j�M)]3y����,�8�k5�TW��t7[�H��%U����L]<�&��3и�3���[8���G]��V���	>��I�4[�Z��V�J��!B˜��;B.SeglT�$�j�����"�`c�:J��e��ˠ��n�DVq����S�'fc�s�n�Ƿ{ܝ��,��1r�\_^,<�;�w��#���V�T0��vf�ZM;��hNA��u�3�����T���̳r�LN����:ә¶�c�t7Z��ڶ��y��)�|.��\�$o�Nӕ�ā`�ػ1ul�q�<�I�����6/���u"��+�Һ�]�3 �v�x |�<�v���|ɶ��*p���-s܍ӓ//�q�͑��h�ǌ�0�y>Owy�u)8��2�]�,�Z��mw�9N{n�Z5�[1�����^�\�9��;��/�m����>�/������������ѿ���7����%{���V��}���N0�oԢX�qT�b�խ���"�h喾m��m'��뾊WIoX�Z�{c�Fn��xq�Mt�3ujX��S]���Y����^FG'�Qҭ��w�S���j�@��vV�EZf�eZMh�����b��T�Ko�ep�4s�08Y6:�q*Źu�s\�WLַ��5�',�K��zH���/��񙭨�2=�i�zhn��K�*<S����3�L��E9|��;t'��g+�Rd�
Q�:�W,��X!!�r�ZD�Go>�K������M�3s�\J���Mw�,aPM}��Ep�y�]E
R�
f/�*fs��̮�{�;H���A�0l�{��:����7��N� ٮ]V��9#ڔ�k/%��b���p�5R?(��W͡����saWc�L�X�/E>��ˍ+M�N�M[��"��� �h�S�j��m��!��RŞ��4ȼ�k�]ܥJj;'���+��	l�+@R��fr㙠ö�İ��<�I3҆v�֙!�7��6�� �m�37����Gt~�ެtQ��Y�;��jҢ����I�9�n�]��"�,�r	#{��e�*���Y�܊\�<���q�hO6K�:eA/ήY&> ��2����)Q�յؔD7ov2�d9��^>銮���;���x�]ueP�:=�<�硷��N����r>R�BaPhETW8:`EAAd<Nz��d�V�I���W�'C�Z��U�f�2$̥B��:�QU\Ir��	�TQDUu��ZZv�)\"/��D$�J�D���㊑+@��F���]I�^#üN4üT�x�#�*)u�r+��	��*(��Ծ$��r���Ǖ:��\Q2
9&�,�"�"�������O+�rx�lrNQHa�ei]#���9WG\�0�����&TPp��˔]�K�$`�t��y��%�9�{5L��wq�bt:�z����"8�V��g����yb|+�J�P�DdRO.ʺ�|O:E�1C�D��Ȉ�(�1d�R#�%ȍ2Z$�Ң*��atY�����r���J�ʨI*黮G:I`QS�Q
�*:R Z��R:�"���Ǔ+�_K�ܝ���f��w�ή�=/�m�z�Y�X9���F�M�b$��9bup���`�����:��C/�ne��T�#y�ϪI]�Vv��]��ej���u��w{�U�����罶բ}]���m)5~����/u��BUWX�7}�ڀ��:o�vĔ�~��D�nzF���vO�r��ǫ��Y�{Vm]s��2_�n{���}[��|�I��qk�.۷_���{,'��T�\7V��x��+��}�ߩ�9����=�����m���}� *��3�����e�����|�{�{�7��l;�	�Aך��3�7r�3Z/ҳ_+�4E
�h��d�^N�w$��Bʷ�lL��څ:`�<Sp�{�X��e.���eP�<�k�ON��h���� >���k�O��f���R��ϼ�^wӴ&2���zM�;����"�s���V(��(�3\�(����k�k1{s,L�oޏ����u��[�@����_i� t�E-8��#���Sڙ|�ez˻խ��%o�U��V��;��C����"��.=�\-�鋝^��{3|�7��w�U�˺u�w�I��g�8o)�ڭr�)՜���Iȸ�Y]{�Lk�P�|�G1'qә(�ɧ3�=}ki��W���ʵ鵔�o�o����sp$��n�/F=�lvm_��%ͩ��R���3�HU�`]{�j����Z�q��dE�癉[Jz�R�ފ��f�n�B�����<�7%�������ݺ��f�dow�N�H/�t�d���c#a�}c�?A=��m������!������qH��M�X��v�C�^d^|�G�� }������S�Wկh�7ߊhe�����O��gX�����. �S�N��3A���`ټ!��`����̋��Rܛ��n�����dӜ�9�Y�f�v�BSo:)�%��z#�=)��u�
�s��O��G�֕΄x�n��ۋ}�{Od�S�L�^Y�{~�<j��b�W㶦�5�ֳ���>��l7\������~O��#���������x��r�Rp�1���4���wY/��B�m�+�4u��Ka�ud����h@4����c�\x�mm΍�J5q�&�ָ�-%�yX(��r�e V�g��ڸ��2[�\J�bU�[��p=��)�S���/h�j�ã5;�3SXl�U�\�G�t���zL�9�`'�]�f���٧����>b��~������.��z��=��]�0=��LΒd����zZ;�Kլy�=!^M�.�{�~�~g�XE��K���B�^^Z�Y��az�F���9ޑ1��3���}������\D^�ʏ���,��C��b��^8鬥�ڨ���.�����[��^����Bz�e�ǫ��㌹�+;Rkد�)���v�ez>��m{g�7+g��p����1�5��Cw����g��[�kAl���ļ���ПL��;/g�;I����~�r���Ͻ^��ճV�関��s}b��s��������P.nW�6�t�TRN�~�'foVOu�yuL�+=sp@�9�>}bߖ_-����YC�U=K�=no�c[3n�e�M�<��%�����~�L���L���õY��U��WyBٗ�y`]e�:�ˌ� �8"z�p��D'�;t#d�'ke?r�:��6��2��N_4nc��{�lǷ*+�����x��{�Q���PDM( �u�y�3�c�J��)�
���.��w�`yM�Mv5���m�+63͝�"�6�u���k[<�"��*��lΏc������~���_�̕�lN����Y�����{�7���o��;�X�{���x��{�NW�\ٗ{,v�뛍p=,���e�����-��0�79��t3�Ɯ���Vk&@�o�m3�hI��I�-/6w1�@�"�K��;���yuOzC]��^���yuپ��zXΓ�{׎��I{4]H���r*x���Df����$��̉f���5��]�O)L����a���;ݱ��{���K}��4���O�/����1�t��rg��Π�������.�#��{��j��m}���W�C�[3�M���Gi1�'w�{�n���M�;��b��N�T~y� �N�<�>Ӻ�����{ϧ�>l��^vmϜ_Wch贚���i�Rī�zoٓ�5�2����Ö\�_X<� �䞶�fE�10��0١�ѽsgm#�5���Z�Lۼwx�}��9�I,c4\͵/�i����`�o��ۥ,�rſ��,�����,y{��5�(G����ޮ��4AΙ�>� ����F�c���h�sn��&oE�&�Z�Sa�oM���b�"2u�G�]g���\��/�I���<��i�s1{�2�p�ڶ�ܽ�Ԙrz�N��
C�f.��勶���y'Z��G�+u/u�z��{½�����W��T��ꆯ�ց7�]g��ޞ-�<��m0��Oٞq�/K��k�m#���j�Ƅ��F�a�<d{�sO44�M�P���߫{���v�^$��QHA�E�=�[N�Y���]�?���2Qc�Ϗ��6e���.��������g��}�{���=���x�~�;v�����ݟ_�#�m����}��F���A�9'h��r+A����m���x��eNw�V{{	U���]t]�0���&ԙ�%�w��n[�V�ix�Vkq���z9��+p_�d��K^�ߺP���ݧ>ػ����̶Sp�i��0w���5��}�^����TûT֝y�6�h~��b��Ʋr�ǛJn�&*4��iH;r��tx�۬WOq�f�ܹoND0[
�K�wɋ�jvK���-�IM�r���Y��D���}����ҳ��cA*�I�/��\^ӏ4	�ؤ2���:���z�G�z�*G�^��}Y�͓y��e�nrѱ�|Na�RO�:�����>m{����\����j��H�)�P=<d>�6[ǽ�T���}��L�<�k�OK���*;��S�Hs���>Z����6��Ϧ2Y��b|o���OgEd3E�/�ww��;(^���g�}ל_Vc����?/y�ŏ%��%��f�R{��So����qO���[���7��k��4=A�=�3m�w���Į�м�K�7�1�ٻ����2�!W�t���(��j��}ѫ�c�b�� �U���G.K��U���m\5j�P�������'B�)tV�v����_l����S�'[����,G-!��϶"p&I�e�oZW�c�gZ*U��,�ھ���(X�[�{Բ�.g��r�w��?h�{���}[�#���QX�Kޔ�i�.�p���9�o��C�e�Ȭ�ݡM�F��46 Uk��w�=��e��"8&AZq�'8��������!G�<�&T;&����RV0(½� ���Y�l�[9N�0s��Hɀc���N��j{Ij@�)r�/[�]����rB{��ʀ���9L�j�v�N�s����{g�C�xw�����}����a2�\bX�zXY�G9��DX�{ݎOvr�y"W��u�TT9�.bOL�Z������ݓ�������d���z�Mχ��Wx>�g1!H��(���Jw�����L�y�1���q�����t�8������j�=����^ԯz(�5+2Qo�A���KL���oގ种xo��cݵ�'77g�ě�-`���$�v�vV���C����K�U3�X�37��2_	��$�ˈ���;���0I�xj��K(8p7���06s�܂�L��i7kqt�'��u��^?{�=��,�5Wk�w�;1z��/�n4���܇��Mq���=��v�����尿�+��f��Zq�f����<z��q<�&��˓Ѷ;�x�m�3�	��{X5��^��O���a�2�i��$t^(a��`��؍ngaU���ɧwW´n� tؙu� 3���f�n������o�'��r.���5���]��r�o�
y����)\�:!��="y��j�ػ�>�L��B�.�z0r�1��Q躯��hT�̻k�sO�q�u�}YK�ĦьW���^��^�E����5q�[��.��}����+,�P�J���ܩ<�)��կ��}�+��~N���E�1x�&-nLy)m�SZ��:���	~J�w`IK��C���S���H�����{�R�]̅�Ϯ�k<@*sŞ�Q:��m�s��c�Ӵh��ū�ߩ�R�9�$��4�i��_H�bZ'��s��Q]<�����jiQ��1�v��Z��n��T������~߄
`�i�8�/��Hn���f�nu�}�u�N׼���"�Or&���P㮭7z�,���^_�/��~�����Hj�{˧�!��z���7�9/"������NQ7�"��n�P�g3���?�i;@6���hև�r���{bJ_y6n2�S��x�3�U�����=�%7���q䧡�(�[4z V-��M�{Ք�`����޹��d�ҝ�s�Af.���n��ٲ�Y��l=�x.���a���<���#�Ǌ[	v9;����M���v��#�:k�����Ol�8��f��Wʅf�.����u��������z �W�����c�@޴~־�!��g?�ѡ�N�Q��"�t��1T,��]�=�Gn�ȫ[R��~N� ��j?n9Ց=��{��3�5���jO{�&<|�s�7�ͽ�|����G/T:�V��}{B�{U��ȟhs>�$��E�;>�n��j��r����Bt�bx�Pع�_s�HW��^U�`�^�������K��A�yTG�k��Yy��[5q���RC�R��N��uR�����R��K�	��DM����p�W���������C�Z�u��'�ҕ��X.-S�ƶ��EQ����Fi/�H��r2}�X�4 7���^ы*�*�~~�U�[���)���}���*?t�2���OR��ȼn���"rP�C��׻7��ZHg�GuEj-�i{ںz�%yo�O�K�zm�%�yk�7��'�������"r�E�V�#��`�Xٍ���:��᧋G �-�x˒^���T��Q��&�ŷ��ݞ�j�[��e�V�}�H��c�	��a%�/w�䛐
w�J��V��.��+Ehb͎C�+Ul�ql�<jQ����ξ�{E�w�ĩ>�̎����^w3��wOT[^�p׏Y�o��c<���N-AK1�6������Ja>S���,�]�7��<�M���Uo'GQ'6n��c5 U�̀�Ms싕:ϻ�o]�~�A���y8��V����c���k$���q#�a��?̻�7�wC��ڊ��jI�,�}I����OCy��6�������x�����Ծ��}=�m�����u�v<���3�h5<��n'��m/u����&o,+)�;�gȽ�@���g��Ճ�L��FY����c�e��� ����t�E֝m���z$�c#����0Ѭ�;����>���ߟ��:1<<��,.�hj�S�az�ޭʞ�囓�%-�ʫ^�YO���䆺ݙ�:x>r[9��<};��צ;[Sw*CW6��`W~���:��������yU+w�~DKf��3�����ٕ}��_e9�S:i��ho�7��ٔ�m63�y�]��T��,�겦�`�|�o�乭aWw���}�)L�Pj���̞z�Vs���V�&BW�aˎ*����Uԕ6U[���Ll�Di:
��:���T�mN+H�;�rf>&]�5���eLv�$�9�*LFuR{j�J���1��:Nޗk!������\�'A!;)�ؚ�M�;4�^�F4��l9�5Ռ�Y�x֜s��k��g'a[�D��Ӵ!��|Ԕu�&������LN��Yxk�*��֍�NU��M��ݪu%4���GF�����5�I��Cs���=�����;7��-��O�7��v��>Ԑ��#�`��t�R�*�r�� ��7�:"'1L�M=p5�$��5�8�.G\7l�<3���m��0N�Cssbμ�� rQP����O���w\L���D;�(�j�	��A1-���Q<��:�6���U�]:Ár��� [�w5np��<��k�j��9tVT��yKu���&z� ��Ln��EӎNtZF~#4lҺ	HIJk��u�2��N�{u�NՐ�H���g[Y���b�qfp��f��"����v!.Ʊ��e����lUE`�T� �p�ه�OaE��Jb�K����*I�3t äJ%��o.n��J����o\�x�)���`�8�i����+Y
ԫM�3�n�d�J�n���&�z�0vM��m��}��M���6���E:D���p-h>����ޓ˛�<��Z�IP�Vn��cڃPX��}Wl$]�xiά����wKU۳-[�g�)�����Έ6�דp�������m�������*Lw��v*Zf�eh�!IvT���4 �Bd�GN�í��=�r�PM#��I�U1���[و��]J�}�-�C����VoCd�ͫS�-�t��[�M�=��SV�j���r�B�?3F��)���!����R��YfoWd,l3�]i��p��S��jSs56�)�f��c�#�M˱ E�3+]e��,i]cnq��TY��*�vQYz�wʷ7�7\� Sj��b�Z�U}˦}�ǏM�]����D�Fe�S�^�n�ft�xV0z�۳i���N��T�hl=�q+�Q����u���f^�Ꚙ��p���OG��aR4NZC��tb��u)���͜����bTt�SmE����[��en����wBr�D�ّ�/�C��o3�����u3PvЮ����Wqt�qΙ:��u��ܥ+�ǽt��Qo�nU��+AX��f��=��8��ǈ;��]��\�;�t�e���瀶`�����Tȥ�k�)�,ۓ�%�pu�PŹ�7^w.���/�BǍ�։W�u��sO�w�Kk���3�f�j��`�y�]xn��շ	�\%T"�-��WVv��7�.����е��wA�Y��O��)̦xȰ�y�H� `�(<<x��^mu~��!�jJ%�HW��* �:U�Z'���
�ͅw�k���g"+��1
�EN�z����+B<�v���$�Iwp�=J�GU��Α�*��zR�S��sP<3� E�L���S�U��tO<�"��d�E�E�E�w�P�> �S�j�a�����9QB{�9˷eEEF�(^���6��

	4��.԰��QQ\t��t��u:��Fc�q&�W���΅ǺԬ�xꮋ*�����.:!�̅J�
�#�*N�EZ�,XT�W��O��|�價e]G;�P_�e�a�ɥ��\�)<I�^H:-�0�/��'6�x�\��)�Y*G���u��E����TEaU��Ur�Zqj˓���y'��.I,���^D%p�AW����p�Պ�VI�9Jн��!J���*G;��\=3�D&UTG)���έI;"e'L%d�y%D�H�H^Ks����A{�Ts�!�wVD<+2B"  �@F�����rG��4��;zQ���I�̠U+eԳa#)�!�f�gD�%m�����'U�93sD ,z���=�ʧ�r�N�)��H��_�#\�E���S'���Ȅoj�=׆���|L��)Nfάy�Ђ����������Ԓ�v7��mBF	�Si���:}1fzeY|��5��C�	x���P�A��sS7z�'1}��NUA���H�}�X9_>�E��D8ـ^B�I�/�fi]1�"�����8��œ�-0�-E�.��ݓ�\�>�k�|�����xٺy���vau�֌�X�{�Z��(��(��/r��]�\�]z2i�˩<�ʺi������_�B��'�-07����ĖsCɓ���c���P���܀�J����	��2j�l�b7SHc=�����m蘤���["�(7�v
��֯fB.��-��EWO�ѥNO�ocvo1{�,.{e��06�t�\�C�t�x����B��V0֠	��r(pPd�9m%���;���/�
�"Dn�a�k+�w:L�ϊ2�[�r�A�SY�T9޺��jv[�8�^�T\!�MІ�n��	ZĨz�J�t�PY���FF^���/�`��+�o�{G�P���j��PZ�A��nlhĄ���`�6�9J�*N����D��;i*���Yx��n�ת����zU�	<}�q��r��E͔`K26�,<�$��Km']��iB�Ϸ*�9ْ���:V$y9��RkdA���RC������i���0h�d���B*So�;�=B�bJ *��!=��V�*Z�b�O<��T-�2Y���؈�v�.�-�5�����Z�v�(W�}_d1Q�㢝/��e��a��A8��
b�Nod��t6Q�v4�L6����kg֧�)�Wڎ��4��h��jG��|�(�J�MI�FN�>��ye.3Ln�'��'�lF���r0)���Pu@*����	3_r �wi��{��ϧ}{���C&��̤X^��BB~��7g�oz��yi��<v;�JK��i8���W'=7��ݾ��5�(��+0���m0��B�R4&y�I8{{v��ش��Gr[;k:qY�br)%N����)�@��akc�j��R�_(�U�s�H��n�v�}��؛m..0Pz7.�c�U+R�J�����d�~�*uϡ:���s���}B�''��6�(�_�Et�[���w�'6P��q�nA�:d��ȓ��W�}
�V��Gރ�E{����ɣ��+1$��Yu؅�ǟVe�0����z���\W,�<�X�|D��	-��L�V8?y�n|&e�u�gY���0*n)E�'J�N,����L��v[g�E�_�:�=�(���E
�W
�je�se��[�a�h`�)��U�.��b��ǵšB����_T�/�[�o=���n�N1{_��"��m��B���;��P䚡��H��ê�'����/;�k<;2������U���9��quY��z�t;m���������\��5���j!��7?={^̓�2��S⚃%vm����8�VC�Y�:����]�m�5�q�*D���r��_O���r�LV+@�6o\zm�c��s�u��S<���8��U���&o�7�i�*DY�L�T%p;��5����qC���lT�C��f�=�1�S	�tȯ�Գ�[��_ZٍY�x�kL%a^O�P��Bg{*��wC�~�艩b[�A{��C	>8hˊ9j���d�Y�3�M�>+�PBɦ%�W��L�}�,��󖥩LF9j����=ݜhV]9Cl�\<�u��7�=5RJ�>����e�ߝ�N�G��(YH�XeςS�p%���h�����璓�}~�L7�⠫�$���s�Rg��Xc�YX��D�
�-�
~9�@Xos�,�u:�ˣ؇Y�v/a����jj{o��[U��UO[�(��NrD��DH���(��H�e���8����dCw��J�s��#�O^о�;�=��B�^�^�$�}p-c^��yo*�LV�y���9�EN��Ә^pt���_p�m��,�6f���rՌ(��5��$�âLW�0�Ki޽��O�;8R�r�wHr��s��_(�@n�f��9��=�3lDd: f��bFq^��Ꙡ��RtIX��G� 62���ؼU�]3B��]e�ML�B�|ۇ.�y�N����m{����Q�QMh0�:r#T'j6�U�wa�_u5�a��v����Y�O2�z���=�˅M�5���V�R�TH���Q��mW�ۈimN���Z�.v%R��^5[��O�w{} ѕ�R�+j{̙XUt+�U��.����؆x��'�/(�1��u�U$�K��G˜�Є6�����}�v��s���]�X�)Z�oZ��5��zH���XW�*�����+K�Wh�.ՉM�u�ݵ#�����k{T'vfs6u��L��L�`��2�t��\�B��e�0�T^L
��WFޔn�����®�J͞/={[�z�Ԇ�9!Ў4KלħL;�T�wg�85��~�ү���L(��k}�-N�M�GNZ'�wb5;c)������7!�vq�.,Ғ��E'�\���J��%@0φ��?i����gyE���������{�{j�1��g臟g�)Jz��kM.���h��yA�sbs���8�<��<�Y�W�k��.c�P���Z^L:�]�j�Rru��N>{��Lv��n�׊�I��
����_�Z|����e�YB�GGP������Ճ"Bl��z4�κ��ܷ�,�I�L})ݣD�yȣ*)S��U�#���JR�g����=Q��է	5�`�WF�q*4��o�L��y��l�5&|�l(����tC��G/6�m��Tw2��43���	�(X8�?ʄ���	Rp��ͯ�<�X��W��b��WN/?�9fm����UY���;]<��KzB�r*�u_'~n$x�b�ݭ���n��d��vU}�c�EH��*����rR�@x#��A:!q�Ӊl��*a�W���6�Yɍ˗�VyPy�R1�=��.�F���UW/^.�v��4q"���e�@}�Wۛ�����39��J�(nA9��ݻl���J=_5���ċ�s悳˷�kȚ��6�C�0֬0��(���Pf\$�jq�f�{�wsn廌;aPCd��.-9	�&cfn,�r��	�[ ����7��x��E}�t�8*�����t}��WXԦ���en�����m_5}����}|�_{�po5oڡJ�qd��a�T��"�d�)��!�ъȻ��Y��d]uUvꎴ��@��$���Sm�-�k�j������'����JmoG�2�׎�|�Κ�Q����	����B�6{�{w4����]c���a����%�aV����k�IKv��9q	C��J�;FJ��M���y)��E�yK_8�{ɠ����ԫv1Q�-��|A��Aa}�q�̶C���L�B�Ȯ���õ��|d��ʗv�pYzo��X��8�LROU��k�H�t9ϭ{Ü��U��*N.���jˑ5q	mj�}�&%y����9��A���,-r����櫖��B��K'kfY}�9�55ɤݹ+;j�#r	N�1�_�$bȜd��KY�Q����dn�\|��L��d��nXIh*��T���/�P�t��r�����S�Ky�_quV}C�|'�l���ʥ��o�U�Z�3p�Χ������̊: �t;�zz�jJ>+�^��2qa|{֩q�g��/��׵y���Oov<���l���z.SJ{�FK-�3�AJW�IK-i!���7^��t�.7�n��K��qe�(��L6��憀����}�5��d++�?aو�t�;Go��g�}؆Fb,��06ac�y�O`��N7<���lb4�UW*n,�_w-MF����è�����4I&+�"y�7t!��d}� gk�ܮ7%1��ފ��I�ٕu��61DЋ����[��5��i��F�(������ͬh�W�ę��7���fa�vk��ը���V$S�(*�Z��^��7����-Rj�e�WC�:|��c�d���f���4�M%;�N����(����ZM��Q��t���E+u��MU�2��Y�5s��v�rY.�]e�ْ,r�0�?�1O{v��3��]��5����jb���C��x�B��"T��&&<u��	��]F�$�LL�����8���d{J��O��l�PT��}	����c�ꛞkn;�n�]x�5mo\�n���n��Sr�C���>�0�z�P�mdKe{T۸<����|sB#֍�_�q�95�ގ��{�-�W	� k�Ǭ����4�X��p�?Er~�c��rߦ!Hq��lR�.��*}7���3�.|�_�ҜJT�5�u8w�Fĳg��/W�E'�[�/c�s���"�OB�k�"1M8����"}p��1��w�Y��s(H��s1T1mK1�)�O^$jt¼�h~�1â�</ub�^=̡���+e��Xg��D�9G�4%p/h\�6�A>��N$Q�57}����w�2�u�s2���Ly���*ꡆL�Lu��e�y���t˞��n�K������]զɚ��|����<�v���3	�{򊔝g���k����N)�R��$u�*/��D��B�0�Z �o�yOъ$V2a����ޮ�/���EY�E>H�>y�����p���T9��2P����z���7if���O?]���\�y^��A=-�~�W��(v�����=Iflժ��dg���r�&��@a�q�o�ʷ*����u]��Ё��R�en�G&����6��OX���u.����8�r!�V�&��w{3Ue�K5}	4���a��
��7��aR��PY�	�s��T�p�����p�E]����@�A��=:�;͟84C9`��S��3��E2�vWYo_�:�e� tdt���ͫ��VԮr�P�م�_Lɲ�tYMv�
���|7�( �& >��nU�c`Ң��_Td�qOk~Y��r�9����wV����x�����Nr�G'�"g&�T���j}f��t�a��G���[Gh�x�!���o@�g�S4��Ru��ш@ud|V"Q/y��,踺b$���]����=��a�;���m� X��U�h��MV�,N2�n'z��V9qU��se�'mMp�L>��Bj,�_��l$�k�=	��p9CX�7�|�^��=���3Ɣǜ�Ӹ�pCɄ|�\�MjTl�X%4�=^;�̟�����!��,��)=(1�[�/Ow�1����l��_����0���|�O#]��W�}Y5���*����E��x�3Ա6���Mϋ�U������U勿bڈy��PJ�RH�W��U����6�۲^|�7):�H���4��(�˓�{�Ҩ+ֳ�P>h�zQ���i��@۬��NRB��7zii�h\nG��m�v�"�/s}�!�;+�o��'X�,�Ю�`d&+�
r��V`��Y�\�����T9�P.�}����F��`�:'��[]�͸o^�~��P�S-�US"�<��n��8�AQ:�9��ӣ���~��7o�.g��19��&����cA�{!LoS��%���MܢZ�W'o�zm�^�q6�gm����7�f�<����fJ:jxBn�d�ay=ƑqniQO�.m?7�5��冦��Ί����a�����*>sa��8������f?I���Do�U�ӹ/���w"��ūz�o/sn�ɤ8M.��05F��z�AZFDC9�r�[�+6�u$��B�:�%�:�[���cca�{�-���=(� N�B���d ����TP��.g��ݣ�*�Urk�7�wpa/��p�)��t�-W��A5Z�Z�ؗ`�Ĉ���`=6�/S̠fL>��D*�rz�4�Ӭw������g�1�}��!gLO��.:�qt���"�z��w_zj6˼�1uv�
��P�9��b8�Fv��ɥܓ��
s4��@�
�|�x���=�\n����('��(Y�~���R���NwfS_(/���=�3�7���8y�(��~G�7�tqԩ���gt�<;S�_Y�b]�{���7؇`7[����Ѿ����e ֹ��*T5�2�=Q�*��.+Q`�����uM�$�y�c�Qr$#�k�ddr�q\�]n���W_v��	}�(���Y�w���J3�����//=���_��C�U��0h���;�B���V�dٳ�Ԑ���B���NA�<�b4v񫌓�w�K��l�=�k�����U=.�*��Z��/t�SZU׽����:���?�ܤ럥֬Y:�c9�������5J�;�C�J#�U;�z��>r�[�	d�u�2�k	u�-s�wHg\nB�z4�r�1c�q,Yy��9����c��G�/`�y_<��T�k��Xv�u��խ�`ۻed���s��p�b���9��6��^�U���:f�k5��!�0h���ݵ8�|��)/�Qʸ�v�Α�8|�.�H�x������2���&��n�s��^d�al�����Xg�#�O�A�O��3G��Yڽؕ�p��+^(�쭯_��5vו���q��ƺS�r7v��A�͐�aZ=^�W��r�Bm+.p�f؞��Pkݾ��L��\��_^�TdY��y�=ꁩ(+�!=��/�	���ަ���s,���m��}�.�x�M]�h�٨M	��{c�B!9+��H�Z���xP��������xVK�k,|���ڝ�ֆ�K��f��J[2��(��{�X�z��R����F�%�;nҷ��Y1��6j�7��㇗FM�km^�֑g�oMö	��!PU����#+�1�5;�<����Z�@�ZM��G��`�u�]�s������)�����y?:�rPtЧ ov+���f�K	�4c>�0^�j]M�k��\�5�+tVu\�ђ���_ԍ�t�����r����0��[V�!R_i�6o� cα�s�s#3){o;MRͶ(h��;�ŗtS)Ȥ��'�֛Ws�Z'�Z��"	Rdu�wE���cg� �6����;��%��h*+-C�Ʈ,���5+U|ip�m�f�Q�2�S�/�7u�i�ָJ����A��$���Ν��*�.mv@��^T:��i���Ѻh�t��yI�Y��4[2���jೊ�lk���`�q�6PD���kIh�y:*��P�C0%*Pj����:��D1�����yԚ��[CQ���8����LĽ��Gw*�k��A����&¢:q�m�u+���iLjq�<�Á�t�E�Mh�";�3�M8"FS�C(;�gsz���P�̓�c�7P޾�jj���evJ�k�ߒ���;�u�j9�P��P��T�C�pNη�����J�|6��:� %��x��	ܖ���T`��m.� b� �)J�u�������s�sZ]u۸�~"Bg2��f�L�������Q�4eN����u)�,��c{e1����=Oi��G�Z5��~�f)�7fJ�r���ցe�`l��X�E��2���*�,�8�/e�%��u�R�j��xSw����:�V6K�e�9�wz�[9�s�T��Θ���ѴVꖠ�;'Ln�Uu<!4y����AE��Q��X�X�eo1+�a�8.*���g��v�3��h��.W]]���CK0w-��}����蠻\1YT�k�*�׆�K�<�:X�$u���S�����HnF�z��S#r�u�o;�T/[�u��U��u=b�e;�[���������1��]v%˰��Ыx�yW�l\�|o9s�pۇ�]���ܝX��o�i�.��ȗ[ċƤƵ�Z�h6�!�2VAq݁�nƤ�nޑ�ɻz�Ϟ�G9ZS�)�����R�=�u�[�7�w(����l���#D�a�U��d�:�N�Zl>y��!�rڗ��vQ�Xd�����9i4�% ݇L�8g	]�i���R�Y`ZE<g�:G��E�]i֬��>�+�z��5ۛ��ҹ����]`q�y}�S<�UrΓ3�˽(v��hĆ��'#{��i9k����¦j뾺�t��<�RK�]3�J����V�b(T{�%����doʝ�C�a��R������h1�n1{]�A�F��fiSm2���lG�aʶ��3S�t�P��H��;�����=�4��K��b��PLˌ���,�^4����&���|j#Q켹^�V��Q��}8����j��������"��P|(��p��k(���L!0�|`�L��AS{����p���/R.V���(�R�Yft�(�39p�D� � ���#�k\��r8�H���(�"�,&QA�+p���[�;�AԂ�QA�J�ʊs�|�K��¨)%�3��NE�T��"���9g� $��g7S�s�z�S�8r#ՔQE\���D�!�C�j��=hy���x���r*����/�#�U�ؕ9'+�fJ�R�n�GT�)R9:^�z!ȣ2�\��+��TEWg"]��\��C���G#�˺�Dk�.S��M�u�r.�!O<��:.���D;���
�3]Ҏp*��*TIj%:�$;�x�U*��(��X��$��eU!ǉ*
���(%9��QȪ��Z���;�դ�#! �9�냩���a�-e��.����q��_^�J'	�R��J�̫̅f��:�&�lӾ��bّ/M����1�&�D�UO�%����<��4.�*���y�=Z���1<���	����F���9��8�u���X5T��[AI�*�5;;�7ܺq���P�8���
��۬ػ$�E�coU]�$�e �O�p��ഌX��2���7'���~�����+<�ђ='	a�\���C�	�{3M
[�+�j����@8���#2=����:ܢp�v�}Z�q=t�2ͮ��;����r�r��g;��$�3���|�<}4�SؠN+G�G��8D��Q֠Cj*R¢�qg*��}�[o�3!{��L2�HqEBf�E�ٳ�]AS�}	����_L{�xi�1�q%X�r����}�,Eu��YQi�5���gMA������w��W�\�K�T'�?ΰg}�s�o�s;5���a���T"6�n�o5�6·T�{aP�l�~Ų'(#X�M�~��oq���jByP�]�rV�}!lJUN9�"�)����L�'jZ��4�p�ZU1�������쎈�.�U����v�����0���}����j� �g�G���𪸾4�T�LgZr�9�.��|��;D����(�N�k�ʌ�3{�6�e�g=(�zsX�ĺپ��@>f��������׌�˯E15
��x�G+�k�N�kYC�;Ml]a�OvM��9�d������K�JW���Vs޺D�@�u��S��=�v��&3&��|�#>D�V��t3�]�J��bB����Ls�j��m����֘u��u�w}{D���4i�����1��*}����b�c�p��`�~q��~�	� �s�_N��B���:�-�o���wT��50����Qn��c��Z��+�n���uK���o��K��09�z��=���߰��:��H�>�-�]:Dۃ���n�l�RUc�����it�$$�>�.��5�a1ڏt�6.�T��nϸ�|�/�%�%ݛ�}窮7�OWrõ��T�\$�˵\�:�+ⴂa8�U3�{=>.���ޟY$�3��妕]S��{�f6{r�=��wG�󪣦�Řk�{��'!�����m>�{�ϔ}���9�u�-e����a�5���}z5RZ�xJ=���B8���DH�����\�I�Z�ۺ������!����~��b��H�+��L�f�����g�4"=���ىR�T��v𹫲!	��B��[^���C1?,��.^q���0,g��`��3��y��E2ׂ�0�5���&��~#p�ع�>*9�}��}s��Ø �k��6�e@��^�ַ�5�]�}ݛ�Wp���m����>���+F�� �u�o-[/x�艺��8y�2M����76�X��ê�3�̓l���3e�ko��72��s�Eۏ��=Vvx�n�����D��}ap�T
��9��X�f[��\&X7�k'��~-���"��ͫs��\Z�����لo(8�8R���z㚶�U��ܪ���!	�˫$R��k�Ie�b�V�W�:xg�җY�	.��B�����4���|��N߸\�a�S^#��.*��u����ׅ�����O^ܳ��~�[��T|�ũ]�je���)��|f�W�,m���̬�"At9 ��,4��Tǜ�]6ڲ��g�)�����1���k�8���'�ǜW��檱;&�׬t�����1)��U)��*��~��&m��������Onzp���ýQ���`�3r��X�;_\v�@[�/P;.w���R~k�������i�eN��n:r�U�'�d5�._0KZwQŲ={qL7��#�N��'�M��cS]2��9��째�@�OYZ��Z�� f)C�:��� 	�g7�T�̷<h�}ҟzV����ݐֱ��GE%ܶ3��x�1r����0�;!K���L��2�`�Z�˳�ӯ]1��;j:�⥷�t��&�"�?jS�sY_b�s��m_� �gi��۝�u�X�9X�.`�R��Cb�9�}.`�7�;{6L�)8h���:.������ʽ�]Zd�۽Kgk�w�K�n����P�՞yN`½UU'w	�Lv�ʏ����F��JT[�t���?JVt��7(������>[��[�Ǫ�V\;n�8��۪NQk9Y���ٴ��ɫ�K���V;�(>���}^��j!�\��lV�G�Ǣ���ָ���mMql&2�'����JѠg�9_+��i>�c�5�/�9S3�u �����PM�=`̻�0�
��͈2�I4�}��;u���FA�d��f�-�~־hPC��8z�G�����1�|P_�͟�kv{��U����:��ޫ�Q;��q���9M�"̇�R�~�kL�������+]�̖��?�����t�x��ξ����1F���0��(,�ʨ���YN�|�-�'���z1�ʑ}d�d�s{y>oLm�1&��Gj��������,�PY��Uo'W���A�\W���͘�3Ӫ��^�d(vq��Ӟ����C���j�<z&):���I���TU�<a�;|�f�}�n�37��w�����#�@���%��nQʸ�_di�|��s֛U�u}�A1)F�:纞����xHʵ6���M,�T����@�n�8;�%���%o�[���w3�����tH"Э]
!�����:𖣴��r�"���`�&Ľ��G+�}Q]^Z�ť�$X��3���Y��|�7�郵ɝ%������ԎW[��;�7��|���&�4��.�	V0f�?LZ��d}uEE������Zʻ�&s���E�%t��P��ǩn���NA�(�.w<M�Ab�bUІ4�_SDZ_J�����韼��|:O:sQ]�2�)�3-a]�B)��a3,�\��ǹ�n�o��{�R@�h'�:�F�˞t�tvĜ��T�8��&�*K��R$���\��M)�0Yctz�yw�ю��>��������F�fo��,\��]�S�=t�d��r5�����&k����?��\ٗ�X��]�3[�g'y�j^JIf㊟��xԡ��fZ�ޑ�;c��	n Z�
	��g����n�����Ne1�,��t�	\|VjFU���9��>�Gy`��%�I��szng��C�FD�ٙz�ȳ:�FK�5W.Q��zu@�P�`FG�T��=�6���~��Sؐ�I�_��׎F��Bg_�r5'_r�jT5�6:�l.��j�����@�qdlXj�j�-�fVI�~����n�������s�"ɐ9����\����'���8�u�5���sR��P�MLV�����R��	��`��̕veC(���&Ft�X���溹�VkJh�v{Fz�D��������a=.�5/�n����]�^��6+휬��Lعԓl�Zz�����S�UU��nt�i�P��ޛ��B^�ŵ��_r���t0|Ș�n:�>��>IH�Р��b�RǏ"�-�9G��">��*�E��ۀ\zɊa��c�0�(z"����P��WBԴڗP��1�_m��i��F�}����T_���Ɏ�/�Ȭ��뎉M�~&.}�4��sbhI�2!��(;��3\��y
/����߹b8�G�ѝ�6jSa	�ˉ�3ΰ�8.����a�W=�zb㲫��ϩG��}o�֝��3���gn�܆�V�1�k�R��x���Wl�=c�!�Ln�μ�e'Y��Ly�
�l�f�l����d�����.�2����^|����n��B���jZ��R�K#uK<Շ,����(��	�0��-�+B����.:_�fn����K�:��7��~��$ٞ���Q��`~�#g\sK˱�����>�`�1Z*H��LF-53�xVO�7�B���q����%����
�V����V�}�P]j�M��p��T9w�( �8�Q쨢�흮#�"36M�kmx�]���m'7����5���Br K�ٙ\&b��>���)���PsT|�t�ኗl
�7Zѣ��x�%r��5���X㞋�9���ixU�ۯK�7��Gk�Qo���e^�S*�y�i�*�+R�o6���-�Blqt���=o��ڳ�45%�>�{�7^��v������R� ��|����k"��ހ��D�H�7�h��P�JJ�K�#������� o=Ry6Gr�+>ޭ9
��x��	G��	�H�E��cq�~�1����Ţ���9G�#lE��έ5�D·Ô�o@�y̲z����+e+ϻu��j��;���㝗u�^jR"D�⦲Q~녫�q4����\���5�,s�d��vs���q���t{(�+S��Q� 6Aa0����p�wO1$̴6�0���P�j����8�A��%Iv�8C��H)��A	v�M�+��"㼮P�V�h����-�^Dv�ʰ���|a��#�ߨU�c�"��b����?���&"5��U���j��5d<�zvo/�eS��\���nKZ�$�ו������[ʈ^6���g�+� %E�ݘ�\�*;͕�yݯl����H���'���X��*��s�]6�Ae�0���`W��E'4v�j��e^��f��(�!���k����m��嫢Zl,���ؕ[myd�~o<5��9%�n���hn�1`40ә���������w`u=$�W'��a�z���K�?88;@;3Gn݆9�	�����7:�U��/9w?u���Â��U�vn�\�J[R��+q]X���Ez�����oQ��в}�,#٧8�J��{�w^���y;�KL�����M���4�;h3m�����S�k����*v
���	{�������~������.0�\|����k	�8���Y��?w�n��m@�K�U������6�/�q�̶���m���x�]Ȥ� `�S�:���&"�𩓃Y~Ȯ�E��n:�k��Z��^��+q��}�u�'����;@tg��
Fw`*�{�ͤ�ؙhc#*�v����I�zhhb�.��6t���9��ϙ��UkW�k�z�l�Q� 9;g2\!��tX����C��p�Z���j���������>�g�g�>������w,���WL�U�%O��E߸��A�
�"�W�m]õ��9�+qҡϨg�n.ܴ\^�U�z����JK���N���2Th�d�\lJ�3 ��ݦ`�oiά�6�q]c;��f,����k8@�{��ATw�5Z�,2�s�^׆��6MF1�ݡ�畍�2����tR��r#Z/��t�V��r�J"����PUޔ�꤯��"E%6�Z���%��Q+���[�:���d�U�y�� <e�_��o�+<�	�2r�칥3V.����ǲJk��Rqk�ӹ$��16��.�Nj�=;�3g'���j�-�L0��Ա��Q@�Q)S����+��Aq�� �p�V�9��k�H/���;sh��{��z�Hx���2��������8�a���VT�(�r��΢O�c�DHyQ5R^�㮼�Dsda������H�"�����sRwD�{�2j"Y6ߒڦ��[Zת.ҞEdR��51N�P�[�}���;+�2D�*�W>�^��_���)��ꖵ�H�s]F2�ɏy{�۽���u��5�t�[�Ɂ{�F�(��p�2��B.7��ik�T��d��^:�{��m����S�|��Xni�1ꋕ�vG�tQdH���t����&2�����]�k/0V��v��tڷ��r�Q�e��H<��k(l������:�C�C�\�ס���J��u�YƋmJ>{7��|���}���le��T��eae=���Y�0���Y�1J}Y��.1զ%N-�}R%��r)�݆L��M)�d��g�hE;�tZH��+Up1o���b�xD;�G0{~/�K�r^������EQ­0�ڞ�Ǟ�5ʹ*E�<�Um-�س�֞
��a,��,�ˊ��%����<hu�3���F�1oib�kz�
��[�}�N��5t��t������#ߦֹ}}6���]���Ȯ��'��~ۦض��������uf��c��^�s�8��.I��[�(�Q��3�������
9ՒR�� L�9�#��4�7�N��d�p&J�g��x{��q����Ft?|��n��_K�t�M���Ԍ�s��'��#���;]�/Q�-u��g�p}tb�c;J�nx�󙦅��V��,�P(N1�_HL�j�D���� =��������rY��4ϐ㆙��x��L3Xl*��tx��j�����@��Ļ�q���I����=e��O�oз���N��P�L�R��?7ꂤk�Bz�8���H��<Lǹ�G��c���]zT�T%U�G/�C|;�R�&����H�����'���ʋ[�����$n��E��Β���>k������U�.�y
⋮���L�kv�S{�M�YQ�B��m֑F��bJE�^>����[�W�9���ú!C6o�;��i���]��o'���l�n�Et�s�rEe�����,1��kE��M���q8�w�y�tvN�?�~�Ζ��2o��S�A��N��O�7������~��+`V��e~���O��}�r�X������4��A�^�;���$���1�8T�eY�{F�f*��3�����OOo����W�����7����Kѹ�-W	nb�$�W<�����OO
:���4��C�-��p:�5���.>j�:oVYyV{�hY����O���ws`����+�%9N|H�ݮ�Z`Ł�m>���u����V��v59w���2îI�o�e���e;��kvф�k��f�}o6�-�t��$�/�DV<vy�s�9;f����ڹ��b�t^V��SwP[��%3M��Y�O��msژe��B't�7�aJwQs�R��M�M\S����z��ud�;j�Ӏ7�r��$�V8p��~��]W�=
��<)�|��k3�rafU��1��C��b�r�f�ܢ�}c&I�u��^��l��;�;��w�l���4���b��-�>aq/uRfj�F�B�ȶn�A���.��{t����si��M �J���9A����K��u�6�&����<bʋ].6:fm��R�Z}v`���J��gu���s�gc#�%lZ[�0j��[ P�Ђ��:�]�nң[�-`�����gu��i�Je�����AS��)��B�����;nwp~�a	M�bl��:N{0(EJ�o�sT4�Ǝ��GS���l�Ȟ���k��ZD����*ٳ�L���_;�P8��Z=%����dۮ�D%g`�}����!LD�d���;�n+���nGCM�G����D�y�9�Џӳ����"��7W�� J>flzQ������N=�l�/+E��Nun˘���K�$�l��,l��iV��I��
������O�p��z@�	V_u��+����+U,MӘ�?F�r�4���n�ps2��W$���y���As��z�N��w�X��t�Zv��NE�tV�Sby�tl�n �Q���]�ڔ���Y1���mӗ�J�:�D�����{�]�F)�a%E	��Y$�,R���d�5ͬ0��7��R�W�ֽ�Gq�H&�h,m�>B�OQ�㽰;�,"��t�\�)�<�`
�݆��N�э�|��Է�â-���p<s�Ti��o$�J��tݚɋR�U�=���FC��E���pWJ��yKS���`�xM���5������>��4Ǯ�LR�m(Ӯ���k�g��c*G�5`�nv�(u�pϚz`��K�yL}Fe� 8���y�g��wR�}�u8�Y;��4uK�s"%W`�e��Wy��M���{G�J�I�q�*����>]N���6��H��w�MY"sme9Ѯ+bv�`��ZM7:o&q^]:`|�5�k���x���[ź��qV���m����YSk�\���14�He
�7�F�Mݍf��.曍+(d�#^�Wt�	��ٴ ��O�J����ڬB��FSܚ���)�;0u�7\��C`ծ%�[�����/<��ݺw�f�:�DS4@CƉ xj���<�9EL���D=�r
#��K�'I��,�*�� �&E"�J�� �Id��W*��4�.r<�WP�¢93�)̢r�
9AUWV�3�\"/LJ�Q˔^�	�K�g ����p��B�s���9}���Q�'*+��DUȂ�)�ģ�T�=Y��M.Uuyй�u�DQE�B
���"�9�*�F�
�v�$"*(�dG5�hX\ֶE%QTs�e�p����Q\����좻DU&QE�D�,�YG9vT�N<�I�Ɇ���K�ʂ(!(�dUr���r����6s��9Ȋ�����t�*��"�&T�"���)Ԉ��˦AE�/rS��P]�`E���}��|||�^�;����%9�9���������N�F)e0�Y��E@5�* ��s1�ý7i.�|Ԡ�b��h�K�&�$��v������ �,oI�7�����%��׭O)|�)�_y����ML3١l����	�`�JOZ��<��Y�I����Е�0�U��� m�"��q`S�(���V��k�]r��9��yVz"]�n��[��Qh?�1���w�晘I̿�;8زT�q���Xjf�9�;S�5�9�J7�e��$�q�[N��Aޕ>:A%��s1�w�(����LV#{��G\D�o-+U��j1��[�*��Q�C�Y���zB�	(G@Q���{�z��B2�,�y7B����R�Kv��4��yB���cZߌ�>>��4xJ=���B8�v���.<�j����G��ޡ
rN=K�>����Cq֚��V�C�V�L�Ω�]�)8r#�z#9K���^��ipU.b#�E��"F��7s�{��:�fC����<�C� xc�A�Զ=��~��Mｏ65[���Z����r@7�� W��p�`�ƇwU45�L���i��*Ŋ�ś#.u��Fr!�{�D�{��M^�!\��x�2�ߌ�?�f�]�������J��-�Y�As��+I�����->�ΚL��uׯ��_� �V�s!���n.�ego;9
0ԋ����Sޕ;`˲�c�5���ɑ�f����]��&��|z9|r-͠��D�gm�#�1v2SxU�L����wɄ����g�U� ����Ӽu���8�֏�eP>NpU˫��~�t�}�#�d��� �W[=f���+0Ъ/m#�Wn�����e�i��,_�l�.����U�œ�o��U����zj�y���/Nbr����� �7�@�tI`LBe�L����Օ6����Wp�xu�uGOTn��y�A�L�l�0.z݂@|��+T�9�Eu,�4nZ�%�+���>����2_�g>����^���J��Y����f�)
wz�!ຝs^�ҳ(�HsU�q�e��������;����_K��T��ޯ���b!�5;��ǷUKztb���We�A��[-\�k^#�>��n*�YZ�r�T�0O�=C�Ti���M�(N��g3=�zhnLj[ʋ[_jU,���[l�F�1��v���HP0�U�;�^49DN,�M�s�j���T�����,�f�5�TS���eZ�3T�U�Ů�vG��xI����;�U���)�uA-_/j�mH�;>k,wO�eW�f���_�m°}Ŏ��1��~ϋ�7����
�c�dthu*���[�����CJ��g�na��-��4}���.�G�LB�-,]�T7���h��=t)�Q��5[���o8*���<uS]�*��?�<yU�2�:�u�KԪn_tQ���CW�m�Y�����$fC۔�M�'gi��N�m���}����Zl�ngK������3[���fН0��`P����ݲ��ī'ȹ
!'~�68*~��c/�	<7��>�a��h-����F�ܞ�0}/�ƀ�TWm˶�=I��E��-'�L�w9�鍥���G���3�`xX�>h%�)��)a���rW�A����j,��-��%j�Q78��pUc�J�1�3T��hN�����8��|�)_��T�:
����"���8��n�j��.��R��К�u���`��O�;��d�k�W3��fxԭ��JS��(�zǇ�&�V��j�8�[#���R5=dԃ��+\�t4�\K&��M�
�ּ��+G~�_+�g��]��h���E�0K���m�0mݳ&Sy ��I�%�9׵�I��˔G�X����e�fv⨎4�n}f��?�Mu`��~5��~~dn���y�?)E�♸eP�/�"v�n�⌹�]���ZrsǕ��6�ZI�2�ǲ?��t���K�|u��vN_1O
o� u��śv��s҆vXR�k���8��a�����6H��sd\P��:C\��7�K_��bG&�w����;hmI�lm�ٸ��Q��[N�zG�^Ė������^YW���m�u;`$w�����[�j}I6;]7,]���Q�-fܮjq�R�zƞ�`�zp|�B��[�x���Tr����z����xx_vq67�[f���ۛ�����e��\���F/�ѭ�;p�������0���f�K��"�N�fnh+Ԙ�+�9S�����m��{}=*����)���[����ywˬ㑪��@��՗z#�nk4�I$�$.a��1���8�#�M%Ja�-�hOB�Ϟ��ɵ�_T��;R}�����������c(��X�U�	kEt\=x��f����y̓M�IW*yE�EL�ޛ�b�RK��T�,%ƼȄ��$N@*�# \<jS�չ?ck�(&��Ft�]����5�³|�AQ']�(,5DJqo�%j�	g`P"�Eb��yo�?�Qw[��k30

۱6̘�t�<I�w��J@�|����.��j���@�]]6�y'w�x����w�D/NO0���Ixf��ّ(��c(VkBI8��&~n���:|FZc%�=��;(���Y
i�>l���rJzڋ��1d�B7U�/j`�S�n8A�6/�2w_�NT�͑Y�"O�눡w��8u��!�]2l�&��b�^ꕯxaP�9���s�mﮱ��
ۡd#��?����v��یu_����z�)�1z��Ԥ콝]���:L�ml��q�j9�V��;ee��[���������}M�t6��i�RX̽Q�gUl���v�Y�#[ح�R2�g?�ѫ���r��z�9�t�r��sK������s�������Pg����Y�_$���?;ê���/�<D�c�>~+����;C���a'��>,��|T\�cS!�w9ה��v�����qw�[P�@��/hǏѝ�6hJ�P�ȉY�܎���:�yFvFc�f;�l���&�_�̢��O�7����3(m�YW�ع}w���_!��_�#��q=Wx��Ժ�2C�b�]:^fO�Eշ�}����&o&;&�r멈f��_q�yf��O�Btg
#��g�P������P��2;�暘��r0ތ�P6�A��-��u�r���:,�R�E+.�C;B`3���S�F�8��_Oj�_�ioK��fG{]����xsrȶ���刨	&�;@LF-53��G�gqL�/&�������h��N�\^�1έGs��T�q�T?>��!���_ ��j�3�{��GLs�Q�}ۻP��t�M��#�����I�s0t����5_r �J�q���(ެ��A��voj۪�nƝT���{r�ܲ�֮��f��cއ�}z5RZ���Q�ܐ��>��Χ9N�n��
D�u���_d	�h5��ތ'�r�i3���E������%y�6��H�Ne�~���7~׋ͱC3����W��gr�l��Zfڑڂ�[�m�K�8�5J57�c�K͊�8��
H{���^y�O�� 6�Z$��K��DH���ᘾ��m���f%��~�^�=�T��ylD�5)�k)��(�Rב%Z�`��%��&�y��t78���P��\�r��A�v{���˔/��R���;��(gEX���q���H��`��H�|��Sط~Z<|I�hi=t�,Sf��nv{r��X�A���7X��
u���0��nK�1m�������٩J�)�-n��܍zRڇT���HJh�jBm�UЬ{������4��v(��/��|���w�d>��˽�z�C%����o\U��ɛ�bT2}>[4��-�oiUt+-����icIC��C��ǻ	Wz�J˵_J�+$��6��������
�c��.����R^����[���{౭ྻ�Lf��F"�ئa#��G����A-r���ħL,����L�&ɀY�gm��c+Qs��%=��T�>5��d4E��9�8jtC;_\v�@^�O�s���6����N^훙W�i�\���4�p�f�.AR��
��~1	�:N-�D��{߲~�.'����-�5�*��P߷3�/8XsϽ��L2\��$wl�岶�6��m�⾼ҢIftx�1Ƹ��ht�.��H�4X�y.��6)m��<:�q/��J80'��.X�]��LK:���7^�KS.������Zn��:���|�?b����k��E0v�=� ������d��%K{���C�V��Gr}j���Օ��$��$��uJ� ���+�Z��y_�ۚˬ7Y�4��V]SP�[@8�KQ�(s�:�.��.Q����!@�n��їf�מ�Ww�E�⧓4%IÑ�4ouε���Cξ&���U����=�f��\כ��y��,�G� Q���
K�ʄ���P�M^���u?*$ύ�՞���N�t���9kw���1��)3CB8�D�|z8����+�/��8��|��̸_*dݘ�s�CE���5s��f5�"k�A���^�;"����wnP�q�����4��k�r��r�s��<~�E�Ndz�p�p��z+�KjW,0���r
��3.
yFt��O\rZ���{�2��i���^�9�U�w���X9_҈�<��������P�^���_yo��^��=����E�O^W>ܿdM���aU~��-D�<KT9�h߱�"*Q췑�� �D
~�u׺2OZUiy?�r<����O��wnļW���3�c�&�9t�6��������S��; ����}��(��e�F�:k�ӈ���y���c=��4=�e�4q�g��޵�:	�}�}��rs��h��*ژ�@s�hr�j5&��Wg8�s��A�"�V���pe�o!ާJw��}��ﾯxx�a�:Lgf;�M��p��x[�]�¹M�0mݳ&ɼM@�烏@����g��]��@14�C��T�U0�En+ʏ?E�߯!Rt">C:)/n	̸U��%�]�>��=������6mtg?Np��:*-985P����5�������� ��$T����#����W¤�[~�Y���K1�U�"���k �EEE�p%@��X��\��`i�����=�]靹L�\�C��̬�9������I�1N��!��Z������a�#��_�O�<���D�N�o�W�߿�.����R�_�ԉ�ӊ���0a��&��z9� �|��n*!��L�3J��g1z� ]%X�$q�h'��P�yA�O�
U�v�{��rrȿ|�
i��Ƿ�`�N�^*mҡ��=��Msv��?��߻ ��J�W5����l�P�͞}�6��+�+��m�ӗn�\n"ې���Ϊ�W�ł��A�a"lԉ��!�9{����i�E�U=�Y9+�H{x�)�)ݤ��۽x�L6��'�ĮT�T(�"R�B�U��sa˲��p��۞�+i ��j��i��P}�'r��g0���<�r�}�^6u/c�P\Wƕ�N��K�=�07���1Tx�'A��%@���F�m��e1s��el��$P�:#. ޞ5��|�gl�˱���u��ʜ�yY�<?<���F��fIn�#3�/��״7i�X��H$λ���aw�e��Ρ�])��)g:�.i��Z���x;!�	�j0!zT�L[��#���ؤwV�C8�qP|bɐۿI]/���ۘϪ����C�/�Z���"�@��d��%�\[#�#�T�9a0�
�h�ՓZ:0)]��缓|ƹ�Jw�"��G�/�}t�%=�r��ySl(n�Z�y5��/r�e6eI]�Ct&�+Vy��X�|D���R6��b����}��q�R��!\n+���y��q����Sc_�Be�~[���wX��7�*��*M�;#M��m�ԞR�$���v=S���szJj�y�4#g�Z���M�yW�X6�[�
�ho+����y`T{��;;5g�DNYѻ/�C.ђh�2�yJ/a��N�tM�.uG����N�Ƶ]+��Zyu�o4)��ea�*QdB��T�uY��^�*
��L$���_��ΤW5E�K��k���b��v{����b	���Y��Qv�G��^1�F�R+o��|ōf
���>��E\n�ne��R�*�7�sc���k�:�^���{i��}U�]�{�18v�96s��3)��ļ=���ڝy�+Q���fI�[i���.y��5b������Kq�;6
z���F�o7Z�Ԛ[�
%�"{����V�%��o�`����{�����2�p���2��~���K<�y��P|V刨!d�q�hLF-53�N@��ٲq�tFz���Z!
Y�Z�y��W�n�~�7�P�=+W�(#ⴂa8�E���P�]�fg��
�v��E2�t��x����Rc �),�A�Q�_s�0�ȃ�P8��hn�4��jYkV�|���l�H�l7�M�hi�e��^����s>�����Ļ�}�,է��J.�k6�F�`���P�"zm��Z�',E���Zy!|�C�Wo@�}�<��E�����n-����AK�lIX��>�nP��
W%=��%��n��Jw.眽Z��j���\�v�X��F����SW��
����V�}�mOE?n�|3�=���a��]y�\_5����_x�|�j/�wG��H��ui#_���F��I�������?̾��`�=��n��蚶ݎ5Mm���iHL�t+ƬiX��꤬���{����|�b�<��!�=!�5H�ʿ�t)�%C'D#�l�l�{$f��Jۘt<+������`3�� �a��-�u�k�L�B�EqI�n�4�	�.����o�B�7����ʺ��3���F�*ɻ�F8�TFԻ�έ��ZnE,�����ض�.�$Q{�]e��@�jR�I�Ҡ�S�:_���z5�O[�o��y�-���ua֦*�7�=�Ԕ�u����"WL��tn]t�R�d�7L�C}X۽�9δj�	����(���ewgu_v�,sؕpWh�Dv�^	Ѱa���%e[��D*���$9�=�DӆPy�vE��U��o7WV�
bv�-����wf�
�{Z��mY
+��x��4��6ݚ�����xULt_J"Kݡ��֓~���c]h�v/����7{�W���G
ʫ#:YS�)��\Ѳ�)��N�y�Iǹ��m���rb�ʾP�{u8��PV��&�{v��14"�&�q=%.컖4nt�kCy�y��1 <�oa����k4�J:[o�u#W��?���U��R�1���X���Ki`�$�j.*^�����UɅ5��JZ��f;r�f١�[�053�p���J��23z�n�}�5]D��uc����m=���4ᾠ���=��;�э��R�rd��)V�_�1Jm���EG԰q�����%���y0�[����Ȯ֒y�.��0=�U���5OhZY��է6��FL�}��<�Qm��7}���@�M�ʚ�^U�G5�]DL�����_ՃUh�h}����9�4=Ja�7��^��%�HE����3����K�k��E�@c�/0�:�+���-�Ԩȃ�pʰ�|.L��`޹�YάB�ۍ)�V�f��P�K����B�l� ��1�>۽�PYRcM�H��C��w5�nOT֙7�aH��w1��y�3{��ܙ�tj"3C���wlf���w
B9] ��8�lV���Y���j����^\��2�Y��FJ6�t�,��rg�c80e.!C��e�Z:V�X�rԬ��K��Ġ�/J�b46&�On���J4U�N>\ng;wt:�+���pק
Oy-�y)e��s�j�>,��<���vj�8n�1ܗ�5a���e�b���ێ:�k5��dY���[k f���Ru�]dzV�C�#�DE��ZX��L�����^�!]a���'�gX��љ��ἦ�7�Ù�3V����%̀�M�W*�ӕ��ơy֥F��j��ɕ%q ���q�L�C*%r]�S�/��QQ��
��f�=ɇ"��@�TжS"<�ëB�-R�.Y�5�An� ��g�`*����ܣ|=���U+��G����us�z�x}qڰ�˚�FF2��y��nD�<�v�l����J�tGUq�9�EC�]ZO��I˲h��:�Y����}���gy�]��)dVۆ�QA.�*�t�d2��2����:s����Mh�8�g]nJ7 �bn��B��NCW :��Յor��BZc#�C�W<T.���A@��T2��
�9�9	⺕\���3��We2���麰��<��!DG#Kd�Z5�OV�r�O����PEk�R*+��9T�C�.��"��]��W9���*4H�����#�(���R��K;8DU��z!G9E2�T�Y�^t��Ȝ�e	!DW9�Rt.s�DEQJ���M ���x���Z�ҩrvxt��Ȅʂ����Ur&�e��+����r>�
��2e��9s�L�Η
���&UEʪ귰�:Q&s�E2ΒZQQ˔���$]�P|e9)XJ�j \((����*��gN"�'W0�&Dp� �#�O)y�9����S2�w�QB��RIPP\�I�%E|�AAv<M9@U4��P�#�TAr;�2;I��<���9<t��^��ٸ������muۑj�����@�gL6���\�����[���V��bUa�ҧ,P��3��lKɝ�ZV�M�|����諭���ׄ�`W/R��o��L�ḳݸ!�M��`����|L�dp��E�.�m�MC�M���f��\���u�����X?v[�N�n����U�n�h,�t�{䡦CPi[toV:}�x�I�Z�r�m��u��WU���JT`G9F�hL�����hBױx��lЯ�����n<���p�0 <���-L�zk=�^*V�5��*��yT�@�|�%�菐��>W�TM�fV�k�jYʡ�#��eO'������CYZ�v�H�@B�C�f�A�V�Ebf���GI����X!���dp�jm:�KPYaAO�� ��-CP�v�7Z�\>/@�୍8{��N&(l�'�yWҥ�5*N�٣{�y?g�Ihʵ^f�fu�b��v�8"����5}�h��=h��2A0p�����1�?G@����|L�����[#�:��k�1�+ى���J\t���' ����$8ﰭ�qv��C����YQ�kr���Yv�k�b7��2,c���txD���҂n1��q�,��ZW��2���z2r��7]�7L�ؼJ�1�C�S�X(�����K�rۭ{s���E�ҧ��"|�ͨ�:��b<\�V��c"����vb����j�<$�M�4�
��0K�l4�.���+J�=�i����Win�H;�}�z`�Y�;`�����W��[���<{�G��k��ܭ4��S1��mr,H�>h%�)��)a�����`���s��/Ӕ�H�wӊ�Y���H�5��H��L�Dx��)
@�ꆫU'�r�W���`���Zm��t�SH�u�j=�Crk��W��ʖO����`Za>�v�Ք�/e˗n˷��4����瓕fR�Nڕ�G�Eȣ��̩�f�|��� ũdK&�g5����{�����qL����[�:W5��V���8�P��+�L�z/���H����>�^��7�z$W��k	��v�ӵݱs��]��["�	Sx�ڮ6}y����)�ڄ�.�^ݐ82:2Ҟ8Z��WgfgS4,`�F�4���+\���H�76�s��v=�A�1��M>�����~�9ʉ��_T�8e�V�G����S�C���(�/���@���H�K�:�צ�n��DdF��̇��zbJ��@J�Y�(<r�bQ��8h�J.�<{��:5��Gn�M��Ô�3ʲ���g4�)'�XE	�_J����O��D��(�;�s�	�?��t�}�K0/K�g�p��y�������N�VM�\��ar�ؘ����a��.��zPx�:��^���o�M�H�ex�=1�p9K~��8vΖ�j����yaX�.�TGx�M�Ӿ�:��/�M���/�X7�͑���RҔ�N���s�}E^Ӟ;O)3 ��� <'4�����f:�=�>�E;�@l6;7�"44?�̼��1^����6���8Ȫ8U��T����s`樭"��5���/����qj^&Ĭ�*�\��2�,�L\�+3~1ڮ=5ѡM����K�9Ɔ_�ϼ0�<��C��Tq`���D0�7f��ێ7�����>ه�p�r���rB�z]���J��ë��!s)�?.�#(9�hP]�+�j��Ί���y���O=����k�i�Q��0$&[���#��;g��6�iȽKz(�3����E5C��`�d����gP�>D���U;.�s]'���M5c�7[�'��QF����x4��?>1��x�QO5w����Gd��u��n(�6�H�8��
���U*��.�xu>�/x35��&d[�=��<[�n�Jm��q�����蹈sA�n�B"��m˃oY1LU�Ģ��LV�dt��Y���.�@�y��R}��+m�Պ�!l�^��,ܕ�_HbR�x�nsMԵ���n��ѧ|ش��f�c`.���Ȥ�~;�/R���+nXP݌e46q����{��C���Q[��o&ZsL�ap.���q�^%�l�t�\�?2���}�u�i��Աj:씵�{|�:�hu�4ŗemH��7���ǀv:�-����-�c����=�����0tq�z���)���I�}��ip�i+�B}��r�\����Stj2���������%�N���[�%�g-�4 o�Y5�I��̤��*|��X3_*�n��(��k�N���}�H���eN�z�z�,5�p8o����кe��<S~�T�Boh��N�s�jɽ̭��1�����1�aP���D�C��W�-H8^C�8i0�R����7��F�!g���-����9��(C�0�Ŕ�v
gl	����m���Rع����w��Wn3�����Pz��H���ųѤm�>+r�T|��a�v�G������y�}]!K��^����0�+��ؽ*cɐ�y1������/��cҵP�Aސ��
S��΢�W���7����Ox��E2��-��V7u&r(,�*�w��u�;ə����v��ݣ5���3?#D�	�m��m7Q�|�M���cٞgאT��Ǣm��_]�[���h�(4y��	�H�T������/��|1Ι��Vxj�|V�ux�U��r/�ߏ�I�%��_-����ĕ��`��.o����e:^݃�fd8Q���<Tný��\���%�郰�B��B_�����''�+6�Ҩ���U�jQ�U�X�'��qSnVּ������9}��6���tp�<��8�RV��׹դ�w�Z�i#����y�;4�[���n2g)��em�x ���$�vK�˯�;��lG�	$��!�v�l���"NI���p.��}�X����V��r���=[���v��9�(@O����H���� ���لz@ȓs�\׊�m�X`R�zw}nt{w���MR6ꭺ���6���	MjBm���S��4�#�6� +���<���ٸ1��ͤ���{�∆��7Y�_q���d�gf�u��omybϽ؄��|��;�N;�W�W' Mz,���x.쩬d��7}q�۶��j[�A���H��n�VԂWX¸��@�w�=��'��r�/U�`Ⱦ�
}<�S�0�!�Q˭��|��7����~&i����urf�%��-m0T�kP��� &�T�櫠:���͙u�t�ae�� �N�sV�)�>��i��ŧ�K��T��+ht�a�;{�������l̀�_�1,�ۺn[�NH��9���;���m��YZ��J��6|��ȡd�zS�B�TY�_�e�w���T��]AO��#�$�cЭi��º6[^{�n�ˬ�E��Ƀ���̛[�W�s��T�|�Io�]�1 5�֮G%��T�unjkY�x���ɽQ-8�Eӵ�.��+EI���(s�8L�^��C��d�V<4��6�4-�F�qV�C)X��hΫ�c��g1p���������ᵖwfb�����@|R|�	y�F�I�#'6�|75�3ڸ�S��'c����^u�o۵q�P��ܣ��OO��!H9�	GU�-SR6�hA�{O}��I�ጚyqܨ���睞�:S��O|c|&����IK�}�`���\q/�T�ʆ�M��,˜��ͱV�/u�c%^� �'�b0��	(3MP���$dB7�~�&w<k�1Z�-R�>Uޓ�wr�m��d�of�4|��<���p�b~n|�K�S[��Cp�&d���Ϗ��5��>�0|&�T�Yw�?3ws0tn�b��)��e��C�˧�f�B�/b�$�'z�FIz�iB)?���1��W�^˚�:�)�U�,�))L��U�6��y�%��~�]�]���F�P��+�^�.�э}��;ǂ-$d
e� ��ʺ��U����g�c73�۪���>���L=ʣ��c�&�x�PߖR0K�=/����c��&��6�޲Y梨һ�sFu����ɥ��RsϞ]��["�(��{�9͜�x�u�S�}=	/�?x��龭Ȧ��xt|�:Y^��	7M	X���� |�	e��1^m^�#��+~��ғ���w��w��ϓC���bD5mϸ�]3�{]������K/���9��ƈ�k/�ml��փ-��i���{��YxRKR��{�RI��&�������K�\Xs*���ӓ��^�YX�Z�71�^;ʢ���f���ӏ����nFe�F���ʸL�7:���x�-a�T_�E�ĨzX��XW"ػ-1����#q>�8�1�ѓ��LR�̌��F~��R�M�.���F��۾u�+�q���շ�I���(ig��!��R�/Z�����*�}=~�����=���̻?�V�S����������?�
����IK�ѤO��yA�O�6x�g��O��X�Z�r�Jߨ��=�-r��^�l��ɚ��z� �g�L��I�g�}(m�ES"3�U}{���ܻ==ݑ)׫i�B�a.�e��P�s1��n,�}ȃ��nJ�H�Ν��F�fud�v�֭�Zf�^�j�yX,�^�bBx�w����
f��sbW*�)gMYY݂�ݪܬ��	���@Er�^/�no��]{.�괶�X]�2�CH*�6��(1p��7�x^���?�JW����s�H��k�0Gۙ�0wVw(�2q}��b�֦B���o@��ݘ��Ю�)?��]�`�2 i��:�鋕N��w��>�{ذ+�p]��R��/��4m2q�q:�/�[�2U�w�}++�.��iە�`��n>¹�G�G�I:�u5���:*O`�*���0��]N��2�9�c�mH�����;�<�5WWq�[���ћ�۱��gC���z�����==��~N�z]Q��\����lW��]b��u7��!��^?6U�_e�ʩZ��O�8�]�I��>IH�>�F�+\��~b�UDY�M���ufʞ�9���mxz�����5�VqS��r�x[��楫�wB�\���������z����y���0�[{�崙w��j�*`�P͚�^�g覷�2�����qv5mC	��U$��û����ʗ����٩M�$yq1�y�>��E���O��ț����fe����կ��f��b+�#�V��B���3(TK�j������`m�}���ޘm?����_X~݂�n��\j��㽲�2�(>{v�1J�k��"��}��R��_Z���蠫zY�?p/�M�6�+uh���Jxv�q�W�޷.ШnQ���/ghJ�v��gyW֧Sd�/ó�ɫݸ����m��
�$�Z��<[��>�"�����-E@HY0q�hLF�4��M�e�2m�ܽ=��sJ��Tx��%�3�ԩq�����cu�_)�B��J�]��]#$~�ۭՕ���V3��7���,��ԅB�^M=	�@ͣF�<��-tjj���Bsm�W9i�jZ��&�����N��PA�@�$�W�Y�;l��8�4uh$=�fY{��$�0��jmMIw�Z{H�"�z��]�����O�j�D�|<=��'(���d��`��z�/Bf	Լ�`��M��'U��%'};'=�q�̷6ОvGq*�)�c4���@4���B��ȟ�,>ܹ��t��ˮl��fSޭ9���tn��/��������s�C��xJ9[�MOإ.�VE�Z�/�x���Mt@�+z��)�e��۝�U1S�Y3=���K�%'[V.���>�9�T�O5�`��U����F�9����d�B.�:0���bm�r0H�5x�2jvaZkbJ���q�7�.Һ]�O�ޤ�7nƶ�3�hj���c@�`�bD�9�AX��'f�*����/��y�W���X0��+���:J����P��@Z��ht+ƬiY�4��ʚ��8)�=�[��`>�����%SC���}ƻe՞���E�ol���]�F^(Y�7���6<!�{*!O�V��_%v������+�r8��@F����/&�8�0G?Y�a׵ͽ8���Q�l�+�,(�����}Wz���T�6�h#�Ɍ��r����$�F݉_I��d�r����l�N����D3R�f@F��fV��2�Ii<͉,�����T�I��;vc�*�tٍ�O��\�M�J�$�Ցn�*O��5�m�{4꫓��{2Z��m�L���[�Osm��p��>�������<L�m�?ۯ���������d�rq��=6�/@��A/�Q�@N�gFk�V��>�vN-ӹSn��z���)%�y�*���I���i�n^->�.
B��
����48wu������o?B�ח��o������1"	*�=�D��u#��Tc?^�ˑ>����~O��}����hUjR�H��!��_��W�����^8�Q^*9�l:�-���O�:��2�b޼�{��Mb�y*> �d ����Ό����q�g=�1s1{&��5'���e]�ѹ�&��Ug4�����j� a;���	�|�Z��r��4��1��R�3NJ�5�oN1��T�k��[:����F��>&��Wmr����	��	
0�FJ��$���ƻ2csk�YLڧ��uNp���F4��P�A��T�<
#F��}`���.��P4��:7�kq�~N��B\i�+�z]�_u|�۩#n�q���06�=zӢ�q�tL��詷���8lG�:���&��{2~�[�2���R1�����vҺ�C�������}`>�1>��¸p��ә�1
�Ӹu�B��ua�xU��3�J�p�+,j/ԷA�]�}L�Ⱥ���3X��	�3iv�:�X6n���H�58JL^f�c�	O�1z5K�8�7���v��kJ��r�Z�}2��!hT�ݺ(o'\4'������g>ha��&`�S2_�D�,��Krb%�eU�7Xp�Ig1#����xN���9��L@nQP����T:uf�Y۷� 
��z�6�W&�.
�	+���+^ֈ�` e@8v�6<��yAI�|M�HᣊT�V�*Q7n�9�U�L<\ ������LY)^�۷ʃ^\�Kz�:��qm>$X�&�J|r����VG��u�y�:�+�[֝��w���$�u-mao�y��+���6r5E��B�~�uh�뜪T��"lO���Ѣ�4Q!�5s�ۓy�����6fH�[}(�b0�1V4��2��^ɻ�C:�b|�~:$��Qi����Q׬uU���6��1v0�N���,��.�F,��&���u:`ٙs�_$��V�vb�o3�D-��ǙB�/�4z��`:�v�x�,9�˖��OyV,�V��fe��DzQF��\۳��t'�ǂ*��%e��1p�%b�{��un�bVWNR�� ��ưTŲ�\a.�H���d�sb$hiWA��^k���1;O6��4����rD؛4ժ+S*�䬁>q�v��n�jQD�Ԁ}��dI��7�8�'���Rڂ�2;��d�B��d��)�������=�����r��Xnr�h�;*�;��)5�M��^�۱�!I~5��-��3�WVI|⩙����4��4�ltL����@�g*��pq�d���l2�6��ڮ��>pcph�iA4��^�^,Ge֍����-h�yj�l�<�d2AzifB��L�[�C7��*j�Hr�z2�鸌�$q��N�}*�}7���­)�gZ�G� ��:�}�Wh����莺�@<ȕ�\c�
��`ݻ{�W¡W��C�C�H4�s�VX�(1�*ߡ��ZZYn�䭦�Q�����-�|i�¤W}�m�3x��gK��S�4������"`-����;ޞ��Tģ���m�������(��������so���iJ�un;D�.����۹8t�R�d��H"GM�Θ�C}��:��=���b���8�k���㍗��LKܽ�+6���E-�hҶ�@��/��An�ʛU��l�|ݰKv�����Հ�0�]Dr�[��L��[Bf�6�@Tڎ^Y�P��	C,eti�B�uΓ�n��y��:�]��lT�2�J�׵�f��#%��+��X��8���̖Y��ie,rӮ�B�(�	2�V��&3�v���νŀ0ȗ��=��\�W��#����\�S�|�@+5&���A/�񕸯T���u6��=���%��s����M�J9O���*�� .P��PTE2��AԢ��wR;��p�S�LH�+��4yk�	��	��ů#i��:w�F�Ȟ2@����9AF!Ap͡	|�9ȣ�S�
N�K���Μ>tp�D�4=H�w��O�&\"��5��.��S�E�*�HZ����u(�� �*-aM"�˅AZ$Tr�
�\���P]H)�+�r�QBd����wXD
,�G�x'��(��'��͟�.�.h��
(�&E��si�Nxv�,NȄ�J��2�;ǜs��Qg"�$����@�R�D�'�""�b=�!-R
(̈���*��u��a�*�g�É�=J(���ucr*���2�*�{:p�B��
u�E�����W=���<���w����0y�:CyE\��ύ	�.l����|4t��(:�ࠣ��wS&�]R�o��<+�  ���MP�?��N�]QUzl�.�_��յ��{�s[���v|��q��{H�{<���*�~��|ޥ/O���D�G�"uR^j�]�\�y\	/�R9���~�;O}�cfȢ`��Q�~꼖���żsE���'(7u�"ߞ"���d�.���6UZ�$c�A�,
�|TR*�"�j���̬�h�~��(v��qM6��kx<������Tm����0��d���{�6���܍�M��7fa��cA��n��}/��
�VTZ~X5P�������s��{�X����t�U�X�Db�FcO�2snY�s��}��Yl�TW��|6�K�Y#��r�����M��5}�gy�������*�<��yAf~�j�s׮���"�3�p�h�g�u[2Ǩ]^�j��D�2�o3�w¶BH�����u�z�/)��H�y�R)�u��d�Y���֚��]���J�t2�k��N�]�9?D`1�q�O��yP�:�/
U�g4VC�f��78����7����y�-*��N�j����z���]����hGȋ�N�r-q �<�y(0daK��0@����)��)�������;*M�q9���ڹ��o��a8�4Tљ�Pؒ��#�y�+�^�����:�<`�7�֐�}8�h�-֧*���UΟh�Y:��"�{Mtcb��a��z�=i�s�{�����&�c�yݤlΤ2�}B�z�P[A�֚n,�D0�7�k�,�7
���ey�zm�_�^N5	��l�MV'W����c�%�ҙ��ؗ.d�Í��ӥ6��*ҁ��cW�O�B��2I�ݙ?pwÔ_%C�I�v���f�{q�,ʬ�{;���|_�c�Z��JYԠN)�[�M�z)���sh���1�%n��ͭu"�|��ϱs���x~�5�_����>_qЧ��#����U*�
9n�%,j���F����^=�:ϵ��?p��X9�_�"NN��JGd����Dz��T��f�6�(��K��ۇ�4����u�����0m�� ����=��Vxk�"�[��R6��Y�׺:�ų���볗Cm;���tJU]����u���ĺe�Bؤ�kv��Y�/}��yp.V�T�㗯�M�1g�m��%�g3 �H���-C'��5�ץ'�O�V�ƺ�6��Ǣru��B����g��|��Э�[h%��?h@��^й��N��~]2�g�a��?z��9��[�od����fNB�֚�Ke{�n,��n{�ǅv��֬,����h�gI��Nʉ���u��o"O:.Q��|��5�;��XVA�D��.�ұ�y��=N���z�]RL�I5��mH&p�v���SRU�%�[�9�&�m�ba�t�'�ekQs9�w����uTOs]n��i��5�Wa�*�乃��i,���.����V����٪���PwC���u��G�rz�c�g9_�,�����hd8�	O�~�����S;b`3��ә���,���w�n\Q�}�)����Uv2�r�s}u��!�p|V�p(�!d����A��ei��{���+���bs{s�9ƅQ­S�ލOI�\_�p�i�,A�1�w��%{�aK�;���k'��g��n���f9��e==E�@����^k�g��q��/��>��� z�������@�܄12< ,>ܹ�LtҢ�:��L�\�^Z�+����������UN��!��8ԈG}#"�A-Y�Flӕ�y��d�m[�t�-}�hg(Q#K=�8�c�S4��RmAX�">�7�"_!sY%:�O������Y�8�isn�;:[E�I����#�8�袚ݘX��m����ݯ��XZ�s�/���p��̋ݳ\��ֿc�Z�:�����p���O�*a���k�i2'������*�m`��T�rc�bR��������G�7u!��^��Q!�Go!�v�~��AZ��Jwa~B���Ԑ���|C��\�[�J\J]���� ���U���T#9#�5�o5�]��춞͓vV��۷Q��}U_N��3�L�����g6����40-:ꭒ�{��75�P��jl�%t+U�	⌬���8������;/$pY,}D� ���q��u� ��Y^- wm+��T1~w]�dd�&�٘����ˋsoN����ƻ�x\�zaPŖ�U�iA�֧��;�{$�鵴�:$���t0�3�=�k�q��d���AuS"�
5�ו6���j��~��Z-zY_�6�����A7�n��W���[[v�/��a,��L�Zdxu,���׎Pw�ں�Ǎ�Z��(����{'<�*`�J��jBv��9�v'��EŇ4��a�SZ}��Ӎõ�D�J��|�td҃s�M��SMkp����R"1��OC'5�,g�T7�	���\�%����ōx�Y�r�N�B�^��:z]"��&�-A�!2#�gf�L����q�:���6P*9�\H~�U���]������R���G��'\���!H���T%N�`���2sk���:���7C6|����ݓ8�f�4��0��f5�Y��r���=" a���)�>2���~:<��+�)�/r6�$R�O���� Ͼ��쟥;s�uz�x�D�W�$�[��[�Ђn��{qo]n5r�=��y�CW�}��m���(��N�x�rn%�)�\f���	�������Rf�7[�Mu-u�"��4us���M;���W��3�+ު��צ;��uD|9�
m9�u>�g��duM}?v�JZk�8�DA9�"_@���q�N�;s��j��r'��se�u�@�iȲ�rV��Ϩ`�橚] D�Ԉ�e�n^x��#Y_{v?�"ϰ��\x�)n;��v�;U�v��4{I���o!�6�;��Of��A�PTT�ͫ�nOm���RXJv��NG5B�����h��pפ�42F��N��e;)�{���N\��&��Ze,ݢ��tqT������n9��~O�9-@�aXU�����rM�V��罸b�g�[�+�_�W�Q%|Y3ţ�n�R.�d��R
y�y`�ݽ��U'��ѧ��b�[��e��ɶ�YT�����I�~�E��ܬ�%�����^���,N�]V=�OU-��Y���K���bM�����E'6Ȧ� ��{�
���x�s�>��W�)z<�u[��{-S���{(��,��#�\�C6\�\�5�@�B����a�`�����lO[�J�-���b���D��?O��Z�-&�^�i�J�[����_vҠK��P�dp�%��M��V��j��O`�w:}���6�i1�=��5G4����(#ٜ�3wx����Tϴ3j���?D}<ƹV�8�u֬*�LT2U�7
m��I
ԭ3���[һZ��i��qct�L�}r��:w[T<^K3/�S��Ү���ɸ��UU�ǽ�䏆B���o�_W���P���R�0�)��O�3����ch&�Si�q��I�׋���f\8p���=�RP
�0�Odu	Q��J���R'T��"��7;SZ�G]��\�]��u��jN�(�e��}y����Ť�LF'D�q��T�|�o�9���S����0�� �^�*�yq�����C�+MvB���4#�dDY0�ҫ6�(p��mz���R��.3L�k���6&���l$hcu�F��3:����=��w{\����1��-��3q��.����v�o�28ܖ��-ܘ��f�-�������3/wr+E�C�&1JW��L�V/j��$�P�ͬh����1��^/]�O=�M������{Jd�,k��:��W�∯�����M��lw�ݥ����x��Ѧ���|�S�(9H�8^��^�lœ?�PT���l|qĈS�@^������5�g�y�������v��sՊ�a�y�U
���P�C�m��	7Y�<EO%�|����?e��R��o��뮲h���o;�jBкq��75�s(����P���6|�̓���ԯ?��&�����l��,��N;A���b4�Aq�^�s1L4 �%fWj����{u�j�
��V��/y�K�cL���ʹ�[1<!�;}��gl�>ܸ�Ϯ=d�0��X�΃t-E'�+(V��XE��B���by7஍C��;���e�C������5]���þ�,ٲa2統I���Ҧ��<i��؝������f$v�ɳ�dř�B).L�O1l��E�9�E��"i�(����r}�_�)cԵ��9�wQ��$ �t8X��/8\�m�g��/��<j���3K+gFT��}A<S.~�T�df�_�e����]�_ֈ�����n���3�q{�P��7/���W59�U25�3�s��_Xq��|��	�0��W�'eU��������6ft�G�fϷ��jP��u{_���a�.(��Q�_5D84U��ȢE�Z��H�eƈOB�zV�y�RԽ1��0S���G�8ػ%R�kz�=z�w8�*p���\�9먼ۅ���T
y�Y��-̘K��@�gL�:繘���)�������J�F)�X�����6"YS�\x�dt��^1i����P8�oHC#�mzh��.@�ˣ־�ҠTb�'|�ޫt���<�,��;y������א7\�V$��e�{�Kz�b��u�S��b��~w�^C���ý']�evق�(�,���d��W��~��h����Ol��wC��
�|�6�M�àE���T}99n�ӹ/�P������+���;��i���-�M��Ux��=B� ��0�(O�D�M�E�"r��ޕj#��n!u�Y�NBx_�S#�S{J�CI����|��Rz��]�d2"D����hhh���;�o
��̖�v�oC'��a�;���m� X�����5[0�:"NV�vz:齈Zs^,�dh��I����2j1dn�k*��0}��
~n8CX�7_c�H%�����i��?`}#���x���+?3��=���BP�Y�;c�8|/��b��&�*�V=p:�{���{�Sr��0��B�T��K���>�6��|�s�ݫ�k�SmD�d��a�:e�"L�b�ǍM�u�],�1N���Y�.��j!�yZX�B�R��T�Ѻ��p3�9�l��ڨ��+x�\vU-a�[q �S"� ]6�K.��OW00^C����0n]���L�����;��y
k4���u!��U���9hN�0[uy*�Րq�����u�P]����k���}7~����Q�.pG�����PU�/����y_��r�Λn;��w@PPy�XO^,�<E�f���y9�v�;n���d��{��~��A�X�{��9�����p�ҧ�$�FhX�vLwӄGA;�4�,mx����QG�ޑ:m^���N4���@�ORCx�k��Ԯ)]o�_5��"K�l�KC0	��Kn��~���|@;���lCT�X�b�og�"@%V��b	tqԎׂ��2����I�}o�� a���%~�Wj
�L��L���~�f�Cu&��/_11���vl]{N����=Gs!�w:s������݀���T%N&jT�3�Nmx�M��S]��k��[�a��_R;j��q�G����0�[���ʤ#��tI�m�����pg��wdB�u��sV���g�l�{�FEuE}#��R�_�.��*�"R�[��W\I.u�I��djz�q:]��r0�M+ih��0W�f���(W�R#;�s�5��o>�_�V�o	�2�6�C0fo������NWh��0Ғ�v6�m�BF	�Y.�<�DaM�
��s;���?��?x�`�Zi�3qg��2�ә�0ln�R1_s�M�i�1K&uK�wO#���I�(��綨Ѯ9�0��Zl��ߊg�.��~Ԧ�W���,�m��ʙ�����p�|��L_�o�V~1%u��p{M@�p(����n�z��
�LW�;��oe><.�{���R��jI�^����!QԔ?y���IBU��y�â@��z��h`=y��ֹ$󃥴y��.�S�"�ڏ
�:����ǟ(������;�]���� �SY�`wa�Y)]��k�]
��ͺ�J��O,s�������G�X�i��z�s�o���(r�Z��d�D�m�W]���3��G�/�B^>�{��3��u�o��+�ݾ-l�]ڐm�� Y�^��v����c_O�x��n�����B�w�W6�ZNi�f�mvs��LJ��w��*Y��}<}�g�6(�`C�T��ǜ�M��"�@~�d�/�=!��\�f����IӐ�S͏��TY!�?Lt��LNfm�G�kr�'�G��MfNA����aD�gvM�r.�Kv��WP��q]�hu|%C�R�>(��ڥz�ODMu�5$�����E�������n�?�c�}��ި��I쎡*7U	R����P�ISN�;.oОM;���B�]z���lO�,���B)�+��G�i8�$C���~����#�L]V+���n��t�΅='�*E�0����<����kOb^+��ԼM���TZ抜�^������x�Ԡ��T^s����c�e�K�c,�h?PUU�^n,�gN=�^�O�kf:tfA�ӳL3�witdϞ�(:�4;��hV	{S�I�y<m��*S��>O����{�kT�]�������+ �P�$�piM����]H^-7��c=Z����n���ļ��e�y��W}V%9��P�§3m��Џ�vDި#	�|(Kt{2�"����󺷵�#Om8��ŏ�z3y�i��n�,ض3�S$�r.xfӔ�,w@�p�Թ��:�3��֞Y�����چMT+˟��Y�̩��Qs���T�̳}[4l�{��³+h�=R����´
���:�G�����K�N'	��`�N���XYa��2/��i9�������ܵ�k_��A]X����[� ���=�ܩ�V���f�"n�Y��^)x��z)w�=
�d�&V�P1s��a�sP�5Q�i������B[����vNhui��Wvښ$����J΁��t��A�uz=�W��^k�v�}�5�Yܾ�)�n��9`�����xp���W+�G$���m)����@� ����G������]vf�3���ɫ��S*H�0�wQ��k����}9(k2�7�t�p4Z��`lҽ�]�$pڭj�����2�%�[o����M�mṫ��r�y6m���sl ��C�λj}|R�
=�����ή[��c�#����e�in�%ESO���z�$VXw�l��NRW:�0�㺅O����ij֚����ϱ��� �E��9L��{��gy>3�X�]���PJ|v�[�e3���ͮ��pu4Z�)�[�Z�w����#'K[Oj�e��X[�����G H�{Ko�'̶��wV�,G[��Mm�3���S�J}��N�Z+U�����3�ͻ���әV��}!�]e7;��gs6%�9�
͌:��6ùa^�����9]����ݐ�t�w�z��)�SWn�/x����;����Ħ,���(�w���l��d�!j�Wwqc�`�r��{.l{��[��y^P���#ˏ5Gu�������j�IcHiF]:f�����V:�SԔ������{�����|5s��?���&u�M��=�Wt�&Sh����k
7��[�J��Ik�[XTv3�û�rCz���Snlvtg���r�n�!�aZ���$���i�J�*��x�.Z�;�Z���m�(����Q������t���e�\#������ʷNY;t�J�����ucV�jv��k�`�C�U��,�].4��]�Tܠ�*�
�bթK�ΫޅV�pVvK�H�!�z�a�zwcc]���v#VÜ�ʕ{���O:�c�L���Hr��=���t)R�J����,I�wg���hrRɈ��]���yf�!:T��-%A;"��V�65^�Q��#��s�:嬤�Υ:16�]7��/����ٸ��`�31KXu�C�JkZ��Z1kk�^ʵ-Z�/y���vp����X��[�:��{�K�f^�X�6҂�L���'i�ܣ���Q�7�u�2��ޗ��1CW]u����w7q��P�L}o8y�G"��Ds�BNn�S)(B=�(u"����5J�j�qJ�2*��»�Ι�h�PWĲ���hd^Dr�� �U*E���vI�(�*���D��R���(��TR��R��Ta�,(��&��f�UU��IU9�f���	N�I�+��PQ\�!*�R��J���%ip�*�V���$�I�p�E�X�M(����)�br���͝��$ �]�Hs<j�QE��
���ւ�&�&ʈ��S�)�6r�

�EQp�F	Fa��IHB��X�A�W+Y�G""(�QI(#�	HEʪ*��b	�	��6��B �eAʪ�\C�QP���s��̖�s�m �Zr%h��:r"�,�G#�J��j�������
�J��Up�����>ow�_*�Q��.�]�\� ����4�+.W"��Eb|\�
W�ӕ�E�z��{9��9�}`m�ʌ��8�ϫ�P� O�V-0�v ⏗@F##ګ����n����>�p��~��뼥�	�>�Zs��>�1�I�g��Otx��j���  N)W�"@�8D���ֽ�#�ߨ�7��>����4��֋�|P��8�O��<�QOb�x�7��)�!{������.��H��̬w�3~�H|Y�9om����t��PC*�^�0�}��P������/����������{�)�AlB��2��`ak՘@�T=�>�Ȝ�udQ�Ǖ��N�z����~��q��Ϙ1f�����R�q�H��V�
�_wC-� �)��{�/n�
vb9�/1=�f��mQ.5;PD��^��
Q�;�,���'ˉ���zŰFɢ��6�;z��Y0��w��L�3=��ӋU�ǣ��6��9{Ob-Aw>�q1jO����pm�{#u`�C����3�u��S�(������*}��f�mɛɎ�3�e�<F4�t˞����3�ߥ͜)��}�޺�OԽ|�,�ui�g�󊗋��i���$�Y��t����i���Wd��)����֮���|�$�ta��$�ץ��R��,�qf,"��־��μ�����'�:+-\7�X���,c<�a�����[K�ÈA�����w��%��Yϧn�\f�eeum姉����y����1>r�=mU7ɽ��l֝�^��>x7!��q� i�6��`k��)�,O"��q�ͪ�,�z��H�4V6��[��w�y�%^�{��Bم?5���-^��\ߪ=�����%R�kz�=Z��`������ןp빺�_�A5I�D��d�#��H%��z���E2��-��V7�>�>�b��no�ެ�}�g������ʹw�(�!H!������W�N����A�ɀڨwY�kd�o�]X��Y���J�]U<OP�z���)��C>�^CJ|`n
q>&��m�����ޮ��m�4�2 a�^z&3s�f��II�ؒ�r_g�����{�z t�Ó�)��E~>�e���ख~��˧0�o��ASlQ�gO^0�1]6���;�9v�W���C����dOб���:o����>�e ۖY������e�}�s�������0cl8!����Q&�֨�.�}(i� e��u�)���(Ih�Rh��r�̬������|^~o��4��9Q�.�������#\���^��[����炩[�8h%��}�o�7m츠��X�l��<vy�S5���������{���+�ɷ���(��!^�9,5w��I.�Ǘt�q��R^a�OT�+A'��Y�q�|	y�o�3�O8�eF!_�>�}��|�n���έ�\�R5��q1|Al��U���,^����bOV|�R��T�e]����<ު����.��sop�4��zh��YaS,S����Yu�(��!��y�7>T'�Q�]��ّf���O�Ӿ�,A�t_�Ga�^Ƒ{�酂�Sw`E^7gA�&b���q:��r*ԧ.�y��DD�Ү�,K����tPU�/����o+�kO�{r���Oz,�n����u���z\�о�@�5o�Wﮒ\u�I���Ȗ]�a��LH�	U��� ��UyC�ض$�r�>��ѹ��B��F0/�qB�j��5�*�_��%SmRZ��;�]3(�����ںcv�u�]��K�wd/B�-CP�v�0��;�|\o/}���J��i��tꍚܽ3���/2m�ҧ���-}j�Ƨ���r�W�= D1�[���\��9�]�������Z{'nKK�:Ǥ���sw�N�6Ϣɐ�F��$ܔ��Ў.H��^��p�Gw�vM��]]�!_�1#b�P���]�r:Zr,�W�3���H�.f�:�~��/��g�([ sܠ|�9�︬�V��|=nB��A=�B�4�1d�f��[Ϭ����;׾ˬ릡�v.tV�n��Č`5[pG��7/"/L����$lT�l����|�+gc�=YcJ���o�1=}r��=1Lü���cs����������M�����	�m�C�,����}k�q��8��J9����cz�K�Per��q�TŽ�'�][իx�dlk�A?��J�j���J�+�A�=�8�˛��Yi���I��j�ĩ�y���L\�?6^����,�4�e�cH$�P/�����b���.0�-E���k�7[�X������v�2V�����W/.Pq]��qW��h߆;�D�-Ǣ#L��W
�J�#�"��jNǈ��Q��hܛ�ٕv�g^޹
�7L���t��C�;�v3��=Rߞ"���S䮙��{�����3c���խ���۫ &��_���1I�>�Iͣ�-��V=W��n�6ݙ9�8N�uH��\N�Zv�`�ܩ/���۝"��|���K\����j�g��F]H��#�����޻�x��Mʡ����
�|J�9�EG3@��giy*-~`"��;�p��S���l]l��l>��;~��%���v�(�C��������E�}�חm��9���@��7�]��k̺|R�j;q_gl?�la�o��{�TIAXFLl��B�Ra������X�����C��W�L�.��7�=.�N7�:6�A\\��v��7Ww7R�z����By�<�)d;���U���961�got��N�[�4�����J!p�n�TOtm4-���WT��� ���$cGKJ���$ر󕿁`r�EՍ��NJ��.
vV��d����iNQ�n��ǣքS�WCc�l�hfO�2�x�%v��ٚ�5�G�΍�S.����=��y�O`�0�g�ռ����kMvB������7&�r��i���$J���-Zh�|��9�:˙��p'F�1�#!�B��z��N�N�uen��W�N� �O�|&�N�/�KT�X�wW�߹P-!B;i����~OR���n��B�����pv�.V5JX� �-V/j�	�u��3k=��bPi��������.��X��*�G?K5���MP�)gP
��s�I��E?G��c����+I\��D�Rή��}�w�\6� ㊂̞��E�Υ��䞯�8ϡN)^�q}�EG�Y�S�����V���/M@�n{]}�X��Ph{���Pn9A�7X��)�Р�څk�[٣���ȗoH��g7�w"#�?��e�.�6�n�o"�n���V�peP���h�(��X'���g�����<M������G�߂��G��D��x���z��f��)��t�\�O����w����.J=�ش���#����ѵH٣Yj�F�gC	�K+�%|5�gF�RK��7s��vO#z5x�:B}j�ہE� �4oV����ƚ��QI��f��VEoed��>�x%rΩ���jsp�9:CI�0�u27�5��#
�d�9����5���N�0�/!���oG��N�̡v�ȯ9�Ʈv��X���9Ǭ&֔N�����/����Ǹ��n�č>��z�?}�]f�{[Yߴ tz�@����#�?][wv��	v�z�t|�)�?g�S�+7cnL�Lu���B��Z?���\�M�؟���y:���c���5AP��D��w����_Z�ӔܼB�ƘJ~Y�W��=n���Mך��Т��ӕr��ʾ�:��<���F\U�U�
0Yr��1C[>��l��7S�շX8�E4���5�LB~h�	��T{������Z��͝j��uY!9���G�6m�޽wu��ӚA�=)��A�!@�i���j�3�ب�S���-�ꡓ<�nH+d���mL��=�R�򼪩��О��@���>�
NC"`,>���E��}����vha�z���Q����ˌkƕ��*r:�8�w��հ	�S��DH���JG��QS��YP�%����4��33չ����n�P=�P�,���f��II�ۓF!ud|o�ٞ!_�R�����V��:c��,���u���n]
a��)2��P�yŝgƒ����Z�O3�ii�����^s�&q����D)>[K��.����#�uәc/�K���n����|����sDw���oD�ήh���s)NR=ާ��V�(��o�ä˂���
���\�Lϵ�9�_E�G������z{���9�5J؈��7C�&��E��6	5MB�&P��W�ĉ��%�8������z��� ��ި"F�Lʹ�������@�4�窼w[�6v��f/���fU3�rb&s&n3݆�i���P�^�fEP�QL��n�����ڽ'��@*|+&�[WklϮ���gtv�m���,d8�d��%��*��7�P�����gވ�SH�jO>�#Gb#�S�U��wV-Ȑ]od����2��%Tȹ��m�*m��� P�꡵����j":DRZ�o#v�Zs�B����{o$HY�ګ�<��0.��hf��^uɈ:X�x�On���g11#���#���7����HS�iҢ�<�)?5�tsm�S��n|+k��{%���w.'��<�"�T�4lt٦41N7����	U��:���(jwS羽�7a֭���M��X��J�9���Q�LD3��Bd���Qx�]��}����|a�X�9�7���ƭg$V��NSP'S�a`Fe�p�&����@U��U���6HW8�<�V�7�XeEu�_AW�j������r��;7�9*���O*J�P�m�0���E��]�}+���{a6��q&��š��M_w]�s�v]9����6�%����q�cҎW@'�@P0vB�\o*�^y�unY�j�3*�6U�3�_`�Z�Ӓz��Jy���拳>�|��W�v5�A���@�zB�i)}��a�E�>�*�΍�s)�F�5V����hll�Y�ϻ��zC����r�嫃���']�r^"Ҷ��	��QL�(�[��u7t���C�e�ı�-�(9�io1��{�Zt{"\V��h�.Dp�}t�n�0a�q�B��nA9��L�o�Q��rA������.m���*��*8}N��޹Ƌ��3��t]�X7�2`����9�g�ٻ�P�G>�aRb���f��;�;mb��-�"<m#\_��	�Ҋ������r�^��7��Ć��l����R�W���>k*�ߛ�':�>���mTD{�T���P��>r�[�pgA���9g�KF�b�hT��"�o,w2�n���5��ɶ�wT{��a��9�Pg�qXE
}�y�Z�ݛ����
�g�t��4M��O��7�q��s�����E6PM���|�b���V�˲.2r���<�s�*��
]Ӊ ��k���M���׃�����d=s�u.�T�c�r�����o���XnF\Cu��2���y��1��9y��{֫9��z���Niɴ�c�W��c�N1bP���l��9��R^�v#c-e���b��M���LʼH�~�c�K�9�9��#G*T���J-99��u��X��F{o={�;�u��?!t��`��U�c�;]QQdLs3��Ak+Ѥ׶t�c[�.aQٺ׊i�h��r�Y��&P��@-�����*�P�T��4���Dc�B^������{�����к��M���K�'e��O�\�s��{����l���C먫�(���ξ�ew9�6Z�Ʉ��o��ڕt���"K϶qP����])��������}�b)+��%$r~�`�}VU��.W��v��3��P��_J�OT��{:�{��鑍iMp~7?5�Y�<
��ӱ����ܷ�����Hf����c�q�H�<hO}�"��<��4:�s+�n$h[�htQ�"�[����q��V��*��v(��b:��n8̄�unO��;_�p�<��T��m2�OdwWr�c5=��]�3�gDO z�.[�RΠ�Q�p�##ګ�	�u���\�d2oaR��Go�]�Q�s�=+ږ�&���u&�x���Z����X�.��Ic��P>�h5G�QL@��ܶ������dRل|{i�)�ʧNc�
��	kt᮶ﮱy�+��3�v����϶��Zo]WYHP}сˍ�ę��ε:����T�1AR^��u��z���[��ܲ�L+���U����ލ���hsLb||#��K�3�B��R��j�5V���S���Y�6�s���R����$d�ɽ9Z��=ʝ��������g^�M�Z|��k��id��75�j[XPOH7���l����u��{�sD�y�J2O1�{�]l��ɠ����u]�R�!o��J���m���N�u�Q뛑�p��m�U�)wm�}	�,�mi���Z|׮�Zz�n�����)%�f�*���"}xƆe�)�D�2��e������˩����8�>c	�<���U����O}M�!��'c�/�1��_���lڌ��7
:˴m�D�(������!��s���+h8s���}�݁���D9��%ƽ[���W��sM������JÞ�0_u�11{SJo,���D�`�H�H�ޘ��	=��T)FW�k� ���<�>�o�1m�Jt�}?_����y�E�V64�c]�6jUn�S���tVn���X�*�hE����9�z��,�K�F*�o+.��̘ZL"����J6����=��W>�*ܓ_R����lm����[�e�dq%�����٠$tU�%÷Z�-E��N]�KM�w�7y���y����^WA��5�{�@�n� �.Z���]���m�1U�9M�+���R!v�K������p������P�Ӯ�~��t��|���D�J�nX�F���p���-����	�7p5@ҹY|�������W��]X,�,ŔU���Nm�Y3��4��p�1Pb���T���;�'�aה�o]p�9�pm/��'z��Ӵ��M��\)^��z��i+�J�4E�&Ð�#\!�0GDh���p�WU���È��%�i� �F����^�
vq�u�)�f#�cҠ��=V��<uE��1ɭ�L�x~Q�U��Z�W}٠EL`��T#azA��ugCM1�%k���٬V���W/5�P�ut1L��\Nw<z]��V@��,f���ʹ؃j��`��y�Wo�5���!bOGn��nƢ>Kv�����%����+#�Y�e�٣,�=���72VV������m�ïl&+l�����k�qf��ћ�����Vq��V�	E�e��6�Z�,=d�3U�xҌR����Y�0뻷�����K�/q�J�Sʔs3�j]ni7�e1�b��eT��F�v0I�28�R�j�2RL�-:���!�%*�Ѹ��}�����%�o���{O�3�I�X�����7,�P�Z��ƲD������G���\�]I�j|���
�)�6�-y(�Gl�elz�&b��-�%זS�L_�$+�R��YJP:G>��nU�&!Ť�{�����c�8yS��*��V^��CVis�ZĴ�8�c#����K4f�=��sfs�6������jf�F޶:�V�'k���u2��^�lh�vN���e�'c0�N�xJ��"ˋC=�;<�='���˼p^����Ù+]�~�T��󫕭�&�ײ��z�2{��͕.*�4�ur�$��/�>�r�#�ӎ�׫c	\m�8�K�zm��{�e�)��.��%�E�5�իuGU���fqIfғ�\Ď��%�R����j�#��X%o���wv�]5�'w�H]fL�� u��P]�	�|��
� �a_pi�^dՋJ�W���,O&9���x�M���L�Z�x��x�~�M�w9^M/6���k��[ۉ��$a����e֛�ɻLa1r:p�U��vAE�0-L�V�U��6\��*��,�3����o^Z��P�g-���w'V��QI����/t�V�
��Y�w�q�:.fT�vJUǨ[��XjNL�;���Vj�	}nSqջ�;����#�bJ-Y��-o �:7�h��CO$%b[�d	�%2�Fq���Yws{iKTQwD��i%)QRr�.rfK-}\H*�A�F`UTQS.\�LNDRq	���"�U	TU*3*��S�Eʵ�N�vQEQ�DJm0���I"�9TiId����P���Vi���Q�TAY���r�W"�(�.+J��<1SD�5-���'ˑKR�r9eNw
"*/Q%f�扑��T˅�Z���!KP�(*�"�e��f&U@WP*�A����M��] �������Ep�
L2,D�"�A�BW��j�^��U%A�����TUUbse]��gSb�W(* I,;p�ʩ8�V�	�2��.*\��#I*�B�%�Q	�$�g3
.Q�a�Ur�B(5�R��W�3�sEG���Wm��S����r���*�g�s�Z�� }v�`P�j�D�=�61(�m�Lթ���Eu���ة�w-<s䳧H����{z細[���BCrt��kγ�1���|�d��y�L�������Ԥ@�>(=�g~H������E��L\��Ol��~'i��1ov<�0g���-�!�r;P�R��sً}W;�@�r;5�����'[�6�N�%Z���e#���[]e�d[#ӹ��:t᭘,@5'�F�>��ktmun��JcA?�(_��k�rtB��󹲯2t-��v̼d5�1�H6m_�t�wK�]�=뭭z	c\TV�l���m6���GKb���1U/f�GuNڬ7�32�X��3�����|���9Q���(��q����;�M��dT;�tg1����zѿa�w'>���y����6� �,���Z�����=^/$xm;��#��3��wot�Y��{+�&���|�T$k�J�amd��Z�W��N�ܳ�)��!�f�Km�6Nk�
'r
rʊ=��4|;Nc�*�������_T��k w��?_�N����rt��w�@�]s1)�����9�xwt�j$�{Cn�b�GiՅIW+oK\�����C6$��խǮ�r2�kzjW���3:�ڵ�&�w�FYv�"F��u�k����J�KJSz��q�A��x`٬<�v{�c�gy�"�u,�ҿ>���=>�Pav�:��`4.%�ژ/:]�?N�m��+���z4��;��Y��_����Ng��w�}0΍�4���7q;�ӻ��)��kg��Q�ΘY�<ۘe�K:���a��>G�K�7JRg���U⻖_�_N!m�ɸ�}vÙ�C��4V+-|�Ơ�Ǻ�^�e!2cے���l�=Ȣ�����jc��z����ʊ�</�_��-Vd@����k��n�dݍB�6ə�h1ܒ�3ò�eOѶMi��`'K�{v*P��XUhԶ��)�7��ip����Q���o�[���v��c�q"t���^�6qFx��Ꝇk���f�U��GkE��}V ��	�/� ە �Tm�f��^����|p��XGy����m4D))չ6�WS��q�MÆz�~8)���Q�����"��vnJ�w:��"�&H�e>6]j��#K��4�@��	��<%��2��wtR�X��`���K_W80;,go@3Rz\���t�A�8A��z�=*���;���e�YZ���
R]��*Ԣ�O�^�Y!u�G�*u t�)x�k5>|��$L���v蟻'��Ip�����k�#E�<R Sx���w���d��X���^ ��{��<u=o�G.�@��4;ae_ R�Y�d�Vm��^tlU����y8oH�'��&�^l��m,�
�寔�ӏ�o]+ ��*�vy�I��s������D��5,�M5Ϡ����p6֚�c	e����]+��&������l�f$���g)���E���l3��������H��/v�N��՗-v@b��/+v�]��n���u�|2!����n�%X�{K2�V�ڌRo�����G��]w+nܔ�?P�� 6΅�9��Q��mD���.Ӻ���mDf�mJ�Y3ل�����9P����[�G���!�ޤh��曄Vfł�H�f!�64�{�S��'O1VoN�>��Ъ�U���E�oX�ʻJU�<�II�n4�1L�78@K���у/S����*�4%�h������VRs}�ns��[��<}uy�w���{9�Ǡh�Y��R�7�B�Y�2�7h[��mG�}�:K ���
�T�l�frEM�z��j<�H	�E�{!XG��-���r��w��֮�:�irGk�mg��Wy���^��V�Ve���1�y�#p��:h����3d��C����=]p�'���#]�K ���t��Cv�3� @|��'�~�H\9c�u���8�diQ�p����8@�F[�����e�c�e؍���*�vf�C0�>lz�[��f�g�Ϳ�n�x�6=}��5�;%���Tk�����r�=Ol�@�;16���Ԭ2�h'���9Z��UuT��v�	���y�޽��A�]șj2\y�T��Yb��M�6��K!�)I�n�M���I7���0j>�~���~`k���=c�\�/���U��~vfNѪ�s1��N�약h-��ŷ��٧Ul� �zm� ��D��bhҔ!�^�u3Um�m�t�=g�i��8�M�U��9^E�9���|Z�?&���M��ݏ:�V+�`b+`�����)PJ��|$�1]��w_�k-�;��@��w_s�5D�뽷{��v=o��K��9Ű^d�������qC���ѭ�3.�	N��u!�}-�*�fЬT$=��hy�e1��TXs+�R��BI��3�w�z�5YX�W�A���Ǐƀc	+/'v���+7���z�m��<��R)�y�;>�s<~������r`���䨚EX�yK����[����Bɨ}�ո�=מ:bQ�sR8�,�K������ ��WR�e��̬��Z�cuVc�ffR�B���e�gt>�G���ƫĥ�A�۶�S��힖����ue��u
n�����KG�����>�HF�NfWr��&�O5�̥�j��tb��5G��N��W��q��XbY��vκ�ھ��{�3*��T���9m���fL�Pn��u��s������U�M1�nt0}:�M>NK�Y�F��=���:�~/���$qY���u\�/�I�^�=7<�
>�t�jO	˫�V4on��� '�t��gn��@�C�w^�ŋ���A���޲�U��"&����]�3�(:�����9X��GdX*��X������U���
�爸i�Jvⓩ�s`Fa�Y�"���K��Э�7Uz�T��TD���L�{�M��Ǧc��΃Ӏ\��%Kޭ���;c��I-��x��i�=���|�Q������a���T�ɟGt����R��"0tS3	�n�5�O6>A�v�#R�J�֫i��%m��2W}l�b{�:�b���.�v3��wG]���c:��.R���v�I�qm�*�+w�V�E�2�����eqO7i�e��Gs`�'����t���-��ժ*�9*�T��3{��7Z�,��n����V��y���-�7A*�U.�J��Mc(���qoYqݺ(�MőW1]K=ǟ������P;t�H���V���z�/,�kp��g�Kܖ����-�l�í�G�s{i�VMD�r˳F{�{��*�\B��R[q�y����C^�W��/9�D<�7�*0]x�˧��|�����]�Lе���j�+��-�y7�;w6�6��&j���|޾�؝�1��2�m���-Y@��rj����xA�h��4��]FT�C ^#	��A,���"j��L^�ii!�yY�Xz"�e���9��Sop)����䩭���G
�1Vu��;#�˖倢��[!��98f�}\(�5os�J]][O�*F��ˬ���&VaW�&�R�D�՘���Y�Q��<(B�&W�wVn�!�PD�1��\�ܒ���[@��j�Ͳft�Y�oK��cy�N�͗����^@q��%>��`ý��IZ�����f��L\[\wmzC��$l�W�.�r�LD+2 �T;F�ê"�gǈ�2�7�1���]��u�P����54�GCb��^�16o1��4��&�M⛼�5�+���yć�Q'�d�.�h�N�ò�Ԍ�X7c��EuZ����@E�{�kF�&���RC
���l�S�������B�q[��{�P����C쥗�F�MP����[@���%y\�K�.cw|ΊH9�I�8����#�V����Mq\�g�3�q�y�5��g^=�E��k�wu�;�?`�Yi+ʢ��E�)�Σ�g'���Ak|i�-<��<�7������7�^+}�����fכ\l\O�@�$5�.���P�,�P�
G���+= ���w��^�{]��ܡ#�*V���O������y���=i��B�dҊw�%3pRW� ��ռ���m
�<�"Ywz̦����)4��얊��Qe�T�![�D�^�Q�3A��Q�������nzv _��Rh9�˶�s#� {�|��5�Ojve���u]쨑)^OM�h��Ҹ�z\�m�7����F���/rR[UV�p_c����W"#��ccl��&8�(TU��OHK[[*!� ͝�^��}���U��}�HF��>2=��uli���Y�g��Ŝ`e�*�̬��ɺx���{����hb��þ+���/ذ�K�n���w�ˉ�o�M��3ҕ�2;ڡ�;o4y�
��<��íV(|�+#M6��n�>c��8�1ۍ��:A�� _O�Z���{X;e������g��I�6r�e%R5�I��p��C|k��>q�t?6������#��	��y��MZZ4��������-Bʦ�<�m�f�Οe�����8��۬��<Ty�jbʐ"o������R���Rw��78XgD�u�<*��s�� �p��֔���1�Â���j��ɾ��4:��㡭;��;l��k�I~}�Y�c�����r0>��e�i�������J̇^u=ɲ'�S�	�L]:�Z�G�tކ�ےM�,
��(y��9�AL5�z��������=���w�@���h�����C٥�(��MvjY6��Q���D���x�>v��G����~@d��wW��Jw_{����n�>�q;����9	��Yy#���X�y�*���K]Ǵ�d�M���Zɪ���4���ӛ}9=5�{(�7��|��9S�[�̾:wJR��57\��v�3]�:��6��WɨrFX�F�b�䯂�y@ɼ������!���6�ƣ�&�!��RmWB�:,�H�J@&��V���fE@mM=Ѧٻ��}���	z;C�����5���j*��D����* ��3�ōq�O9�|��-�@:�Jވ}�(����O�)O��orU��r{s	��ˮ��<[��+�}�Kj>ށ��ᴴ2�w^�'a�2��F'�u�7����L\�dU�)v{q)zouZ�y3#��T0c����!ύ�yׯ3%����Ӄ^q��M@V\�Q�T#;��h�{���s:�F��	*��G/i§,�[�Vj����k8�Z�%�Jﰼ�Ӵ��P
39e��a`�rm�R�q�j�����|;8�����i�Hv�b��U�ˣ�4fʴ��;cbu�J�r��[<�xI�n:��[�7H��Z�V]XT��M�W��8T 4�Ǣ��[b���n�m%�x�	��
krl�������p�0m�i����	��X=�wF�f' S�Y���\;{[�M缧��J�[^~?�CqT�~ڠт�|+bl�n-5���I����&�`��Y/q4l�U1�Xb�F.".V۴i�S��g�:z�f�Gu*���ت�A��л15{�v�b�6.��9R� ����˿��J��=fE�w��Z��O ��*�7+;M�h���Mi���gw:��Amyv���$K�-yV؋n�t��}vfߺ��p�Eie{�!!�d<R�A�8�&R�U"s�7 �TK�T�`�g.�s���Ws������#�i��]�A�{Zu.�7A*�*]ަ���=�)=��m>M\�w9̽_+��A�m���u�n��>��x���}y�3bޢ�^�ѷ�����e1�.N��C\3w����U;ʦ����iԼ�
$d�5crNP��=�[��\	&{�T��>K7���iglV��I��b�{Ky�w�Ϩ`c/IE�u�M�\� v��8���LRJ1�GTW�0j����T��ښ��#E��i�kzSz@�����B��@���B�T8�����!�g8^��dtw��R�v�7��%���6c��t�b�s��ngKo� �t>�$��9���GD�>��^ՙl���l��-��N�\2�8�I�mJӴ��5�M�m��s7��f��6q�P�s"`ue�qS����[�4�V�9gZyЃCU�,{�K ����&��/��X��\P��������vjT�ܒQ�����$�Hk�O�?�:�����x�Ϛכ�ig	LW{�[�Y�'K�'|)7w�6] 4�	�pVA�2�O.fb��\ҷS!Jෲ�*0G��#y���Q�0Y��Wi��W�n�WYz��ga@�m��X��m�=�7,d���J�Pg[��"�c�]u3���p��Q�N�N;��nv��kߢ�#�"y8qG&aߌ=\ƃ�pki����j��a��s�׬ţi��!gN�f�l�owYIv���[o1:�í`���ͬt�(�����c�S���Y��y��0�y�:�)`���1�uGu�P������-Ѱc�i�P{ؕ-�n���8g�<$3��Y�|��
��xڌ�y�*m��Z�M�]����c�&2�7{ͪB��Xc���&}i,�~	m�T8x)�v�v�ظ�)��"���!Ne�{wO.�4smX��5��N�h��Vz�`5��ِ�xv���m�c�!Z#�S?���Y�:��/qf������m���蒟tw��NM|7�V�2o"^�p���H���5q(Wv��Gr��)�3(�/p�g��\�cr�#��5�fR��jc���vp�V�C��Ժ�R�֒�6NqQ��}v�u�ޮʋ.� �9G*d��J�F��R8+N��2v;���}v:L!�òU�Mc�;#��ytq�x���}T5m���P��&*�S�ܛ�E��˻b����]��t0:�rlW��Noš��#K��QX6�R��ʗ.��]�l!�8����BR'��L��r8�yz�*t��/�l�+s�I)y:��,&�S{Hqcᖪ��)�y�:�IO�m��������ԍ4+�b&�:	#e�ݭ��^Œ�G�ʸjӔ��6��J*��i{����}o��qP��G��%�)��MZW�Ν�B@���wP�����K��6��2�j@�q��4N��ښ��"��Vȟ9�AQ*i�нE�o���~5r��o{|����{�)4c�w��bŲqD�U�<`ڂ�h�<���iSp�`�/o5�S�n��^WjU�F�I�B�4��!cN�J��<����.�-��u�v��$��!�+��@ �U��Tt�EJ�[��^��E� OqdW.ʻ.�;�EUU2Ô�gE����H
���BuR�����f�)
��G)Q �NRQQ3Zd+��*�C(�;H�H��E�(`����ʂ*�����i�bHq*iE�D��
���5	�iP�C�Ȯ�-B�M�rʌ���";�T����Ң:Yl�*�B"��TYIe�*�9�B�N"��� �R�Re]2H,�*ȥ"D�#K���$�b�+��0,VF�*��f.����P�%R#$����]D*:r�T��"�����,�Pe(�4�%*I��S8�A�6h�bIZQV�p�8r��Ң�(��>�N�1j�v�ǱTl��	�;���1���������n�K�U-�ގ@�����Lrk���-�lu�ov����#�u��@1���]������گǻd$��B&t�3||��)�K|y�;߭d��p��)�V)��t&�?5����s|�mv����ZfOg�KN� �]�c�˼�U�q5U�a���5�Lq�����`�����?k;�əs�هzkۗ�{Ȱf�,�s;��w�Q�{���$��jcG[D.���*��M�co7������W����_F����~'�ڽg��#��2{�]wNn�a���H��;ڣ�1�dF�a�v��CWA�+Q؄F��iF{��r!����u�=ۺ$lN��hD+�S�/�Ϡ�]�d��ںr�yOY�%�2��wK6�k�o_1�G4r �M.i��6)x�� B)e���p4eu�=w����Fw����>�A�̲B�v�ʝOKb��"�1�v�ڋ�<+-�Jk�&������('�G���q���N+r�������b|`&�fF�m˲���NѭB��u�8�����u�;�q�3�7���v<��fmd�.j�'Ie\{*=�8-W�q�[Һ�.�,E��p��C�	�h�e�eN2d(�gZ��I�.J��^-���>��C;��&����hy�2W����$����|�$S�_�*��Ǉ��T��YW{7���iM�o��e��AtMr/�	�Zm�Q�La����z2n����檽�*�+�.��<-Ԁ[�e�D$6}|�kO���2i4,�eq�'�L��el��w	����7kh�ȟ܌T}�������w�:�l�ɽ��ͼx]�l�p�Ty8l��f�vM����a��U���
.7{ �n��şFS�˴�Q#��˗�����:춆FB��h;݈��ë��>��B�^��j?�	��B�Wq�ʌα���zY{�׳ٍ��;R�f��矆�q��fgc�j�r+l���D�^#:��?7��l�����������#����y�F��C%s�ܽʝ/��j\��͹��,Udf��7��(����3��|��11a�~���^���v|PBR	� bw��0{d��>�գJ��������������0�AlƦ�$
��ޙ��Z2K�4Ia0�3�"b�o:!ط�S;iԼq)b����G!1m*��Q�mp�c��pWV�]��Q�E��v��s�a[6�Ƴ������3��)LK����ݑ���i2]f.M��ǖҚS�4��l,2��8{¡*~��]7{�-�QJr6=ZV�v�Lҥ"_�I�p�������T띰����P�����8OK�`�s�|"l��]^݆��-�$7��Ub%7cd߮��-ژ�w�{�+U5�LZOԳ�t��yyHɎ�}��:v3�>�GxL�Ĳ٣�i�:Zԇ7��f�_���O_��[4Q��Ӑ��5�*��'<gp���i�U�X�,�@k�k��Z�)׶5��a����!���t�_���*�ee U�W�㩼e��zm��r����g'4���`j�Kۡ���?B�Ў_������$r������:��q�'����\��Υy>� Ɏo������$e�$o��IY��kK�+���rOxoL���O�#�#��W���PYv�䴚EZyZ�_<�DzD_�sz�Ñ pp
����n��,_ry�+3vD�������&j��dIj//�嵗w)ΫfM�8r�el��������dӈ`X��.rY�U�54%�2!'�D�S+mT�-oVF9ə�I*�ffn�u�By�Kml��H�;>�\wc����a�~�����qj���;���f$%ɞ��9#��n�|^l�Y�s��x�8�y� w�Թo8���y�����&�;�/�a�B���z�=��޳�;��]C�鎭�;��53DL��yY:���=���k�3��d* ��ۺ�)�o{���K��n��##3�����\��[�z(����}�[5m7�Y�r~ݽ�I��W0�؞!Z�aܙ��o+8���g4:B�M��x�m�KT��,{���r�����[�"pS�Qv�fQ6�z��Jc(@��`��I-��,FoZc,�vK��G;Y2"ґf�ۋl�C�z1�g���V�e���F��C�<�\��hi���|��SY�M31w���VUpl�;�n���S!�{��n���)m�o�v�)����Y���ߴ��ܹ�N"v�6H�Z.�Ŏ2..�7�qv=崗�ո�Dm�xL}�Ԥ˸^qx����o~��`�:'�Y&�:�{=�xI���Q9�����X�fQޜ̽�Kز��:�����^�z���[�:�)s�k��l����z,�%ڽ�[�������e�a���s�F�hP&�wB� �׼�Nׯ���,��j��e>>�<�ٺ9gi�Ʀ�G̫��k�d<R�O�Ɓ2�������tF�fq�N�ے���?~~��O�d�5��d?��ͩv��%h��X�75n-�@�7���Mg_^�MGr���m~7��<;��e�7�V5��N-傳/3c'M��uZ��IgW�!��0�l��m��WaNM
W�Y]�ձ�RE�u>�F�˂~� ��±��G{w�N_?r�ʂ�������̝���hL(��5Q���qt*�ܱ�v��<��S2ԡ^X�ș��NVR[G'7��:Ŭvσ�Q[�C�j���\M0	���M����Rʪؽɾa���}w�u��[��ܪ`u��M�8s�,�ݍ��g�﮺������Vt�5�fQ4g��a�?�"7�Xf������ԙ�/�{V5q���ǎ��k��Aj[��L��o���4�Yb�p*�b��oCy��
�`�������V�2��ӗƑ�@�����5ʥF�V�@P�u�դ�};vT��׉��Ġ{+zE.�)%�:-h��ə���t6�u�
T������W�8$(�-�H�l�q�ȼz��I��pb��kݪ��]�&L���;�uε�`�d.�� ەڌ��[�+?A�ċӓ�R���j�?%���oF�$⧟���~{�u�~&�,��C�GlOv��ۇ�>jU1�dD�V��6O��A= P�	T�*e����S��o�*�ʻ���k\;���g�w��y�Qˢ�&��l+�_!ʖJڞ�J���֫���a��~�Ly̜u��������Y7�?�}��}^zGfkȌ^�]�m���'ex�ɦ*�$^2�kM5��3�,�9J"F������zns^|4�ɴ
��c
��yf^�&�$���)�Uwg�˺�pӍ",���iǤ7%Ĵ,�+�Y��A�w[i���Ђ��L��OÄ<M�|َH�;|����F�=�rz��nE��֧&���+S^���"���-�Y�.6|10*�f��!�YB�G�ۭ��ew��,���j�����nn��*����Gps�
m@�\�U&�Ӛ�D��yt�[.�}�r�G	�!�3[��Ԣ}$��s�u��C������56���딦��I�|����V�t�&�޹��z�����ۤ�µ���3� Է=6>������m|��_h��>�o��q���u�Λ�Ed�u3QBJ|�QS�k�t־�N'�c��Sl���t��Q�p�JȽ��r����'M��d��:�f�9\u��[��v[�=#~�E�4���ԫ�/u7N���]n�띾�3Gui���R�]i��G[AM)�dvK������+\i�qUٻ�c��輹��N��>�� ��զaj�,@�W��3�6��'32Kۭ�{��S�֢2܁�t����|�$u��-c�]�k�[f�)I}���������>'���?�}T*]���Mw)y�@�4m4�f���u�4A
��l�Ɲ�͹�b�|�%eѩ�����[z������w[noh��"���79ZmUX�,����@�b���?��e���˛ImN�ޠf��(�d-�ƫ7J��e��N�a�;��Y�{wC䣱u��\��wZOdV6ei�*�J�=��7W�:w��Ԯ��f뚶qk㧍D��v�Q���/���H��0��.��{wkm78��ȿ	��?~���B-eex���n��Hk��ھ�֥�� �m�hZwi�[w2�Co�c?9�n�r��M�z�]�W+ȡsv�R"�lT5���y��Z�Ց��͒��~��|��La%~���+c����C�<6�~�w�e�2���;������=R?��"Ͷ�%��E+���,�������3���i�v�6�K�tí~\w��<�D�Fah!�6{CM�S�>�ܵQ�JY���o�w.Ă�dB͑ϩ;>����[s�]{�kr!J��ߨ�ڷ�{�wmg��M�}� �a�K��O�3٭W���vd�^u	���D�Y���k����+!P>�����73ԝ�ڲ6��hZ����IX�~��Þ;W�;��<a9����e�|RSW��sɛ�Q������e���{Ǐ݇w��>�:ߗv4�����
e��i��Q.����]Ե��Q�ЍyV{���n��@���p��jd���,�\x�C��
�i�+bߊ�|8�����p�IvgfF�}ډs��G�'�z��������i�H[��EJW&'�mCSgl����n���*��>.�NV"���Դlj	�c]h�}�m��/ B�"���ѽ��ǦT��i��󯩧Wcq�:F��&�#l���/k&}T��7�Ȇc2�ܦ.s�MoF�F�7��rJ8$��E��m�@�N�l��
.:��x�س|��)N��v�|�0�nd��b�5r��
���E�~���O/_`��<�Cyz6�����S���:�.�R�78hwB�����N�y~g��p�@�g�Ct������]�*o,����P&��F�0�PJJ�<��=��L����$T���d���W|��3-�i�c�����5K��f饯c��4�q}�˛�Ii�N&�p��+�� �[;�9M�#���<4j�"W*��X(�}�Ö�O�lO������ւNuA&[������ݛ�����vOEe���ٙ����f���~:9�
���8V?�3X 2�ѳт:��H�E�}�*��eX��~��M������%%�#�3�ҊY�4�~�<��޿p�!��,��Xټ([��Q����;-mG�j�ot̨���V��Q�����U�U�Q�Satt�V|{�[��u�G���ӵ���R�s�I+��
<c�SK^B˦��>����~c[hSf�SWPꃲ��:���G��T7�o���g1fϵk{��f'�>.����3'KSի���zZ�:j6O>7�A۶P���@�� m���Hc���>D�6Pȸ�VF(�6-N�D�ό��6��i�쉟F��T���bP�m��zWk9���fߗq��Y#c9MD��\dٸ�O�-p[�w�O�qn��a��U��pK�Љ�����0@*��z���nB�xc�u��[�|��ȋ�x�s�w�v_��5��#Iey���)�+'�<�
Y��]�76Ȭ��E���ʽ�Ρ�I�('����r,�k�i�K����]��#��'�6|���e�`�[뉏n%�/P+�ac5[|K��iw�ǣ��W�Aȹ��MP
mR�<Ɣ�����mo �>�/g����Vg5p~��Ԩ�2���(;��Ju�ܮ�bYVq@���΂�RgL�m4�	�z�5����`�՝���b� ]2�w�b�B�M��k��4�ɯMy�:#�� �MVZ��;�&�H/�
=�7����'Zx)�Df˔7�R�&�X�kf�g(��-�8ū���7�N{���b�!`&D`l�h��j��МP�y�·Uv���S�r��u���l��JQv�`�g��R��xR�d�G���2��[��֥\Mf-�:�ٮ�y��-D+Y��O����C]��Sg�n��8��]�ti�K]
�k���]7���S��\)��V|'t�H�֪\]p�N��"��+'�����+�fV�%�%f��N�![EgȷV��Z�GE�Qjr���q·;��y`GI�vv����t�
����3f6�
��5)-�M��(
�wy�j �j��(�x��J:{`ŵ�R�
���NO���Sz��i�;�p q�ƦD�I��#l>�J�������p�ӥ�^�Շ+�-�Y�h��h�2 )�Ä�������]5XA�:��镺��[�R��w���y��<���ve{�Ԩ�ky��}�خnSE:԰"A˳M���I�)w`W!��Ҹ�R�p�w��ƚ4Ʈ9�ʽ7���i�yu�����<�8P�]qwS�יԠ�h��v�������h{�J}��ý9۲��Ȱ@E=���s�j�t���s3��̂Z�]ep@`l��{En��MC9�
�<�5�"��A[�����M��=��3�U�MA�b��Ը	ʔ��b��1���a��;�Zw�OM��H��L<x�~ݬ�Z�\�]�����kk3���n�wN�c��oy�J���N���}2�M�|G�ͩ���_FUeabr�w�p�]��"_`�g(3��P�4Z�F`�@3D�3�M(�o����J��飽�01Fu"�v�<��V����x�������n��ƴZV_}��I�v��8gbW1�����ݡwB�.��� �x��,�4�xK���_w]i�)-����l؎�K���NK�eM[�Np���Âf���%�EӫEݔ�k�rl�<�����vٛ20����>�'BIOo-lGb����*x�����k��k�p�[��c�ipT�8�:�I3��x���խt9M���6�Jd��J��&�����
�jΔQy�\F�s��`��1���Wlʖ����\{���D��<(���7vm6�k&�/" ��4���iuRXkQ�l�z9���P���dg,�)�tT9�eC�^�a��Շd��y<�F�u�N�A# S!�3�F����ȶR��df����vNص]�f�ߝ0%�ؠ51B��^��s�ɧ �nW �9W�M��}�5��W8c��}S�	.[Ҭ���g�uq48=��� ���(�G��ah��$�ʃ�PZ�*��%Vh�ʪ�Ŕf�*���E\�d����RR(�3A?[ X��N{������;.\��$�NP��,�EJ.r�A!�B�"�Q�DQ�Pf���9���G��/;=/*��9��uqN��L��iG˞Z�R^'����i�I�U�kΞn{��˸�:\sVP�&JJmJ����qۦ�,�Bc�N"���E.�T��T���efʊ�o;�\�LXE�<q
"q^Z�	*D��G"H�9ʜ��"�AEE
Ш-J��i�Ⱥ$\���*��9TY�YI�-$Q�NQ\#�'*����5�QM%���{(&E	�@̵+�B|t���I�jRy�g���\�Ls"��,�R8�+)�:��C�~$�E���R�7�����kf)F�s��G��S`4�bw��9uץN�e&xc���Z�I���Ψ��B�ڗS��T+0��R[����v��;���Tg
��V�g�_M5�,
hO��9�Sv�d��9uv�4��eĐ]u���5tZ���;�'�U6�DF���,��y�Q��:�y���������'��edyWVTu(�X��l��m��x�L��z��S�*o��s9P�\K$Q�~ܛ����d�<��5�y�"�����<�9>�<��aq�q���	�7I���q�_\5�W^u��ֳ]A�3����M����~9��[�Q�'��4�T���ј�������T�ԟ��֎7��M�{z<���~�P�&����D�&ī�&.H��w,�Vlb<��JV�{ڣ�1�o4�݋�oٜ�Z�K�Μ�IX�q::��4:�)�,h1ួE]gQ���6�m4������P��|@�@]bѮ�I��/|���r�I��L^`U��y�a���XCC���ņFf)x���b�^�{*/z�a1YI9�@3a��{��f텅پӸ��m���QX����w۫\@�d)�zØ��ᑁ���z��8{_E
��y-�]޼������Ӧ��)7V�ۇ��jVϣ�)�P���S�N����/�0ffa~źJ!,�I���S�����x�cL�w��y��Sf����Ϟ6Y���+�.VwQb�mtp8���;����eL�42s���EFO�[7)z0�X�*Z��&���e�/ڞ�/�f>�ܥ�l�����UɭW�X��=�5~��'\�^����g|�пP�؛���7��TJ�7iUOY��Cv�&�hY����}��{Hu�`�fz�>��^~�49���+�Y*��X<e�t�[�tw�" �5�Hl����n!�����Hߙ����3����|j��V�T���Bȗ/������v�h*(!Ho<�M�˴�Kv6ࣀ�f˺���ii��>��'�k��u��#���wY8�8V{ �ee�5d��s��E���s��L<�:��Qe���ώ�?��yV�����/}JT�>�2V��7+�f�y�ȕ�[]�Kv�Y}�F��*Z������j�����x�8��̈�����Ao���e�TsT�U�Hꄤ����+��q��՜�7���7!�D��Z���v6�c�DWƂy�S���N�g�K���F�nr�Ť���-�JO�>9�տ��~T�Q�+�#���a5�[8�શ����c�e�jRĿ_ﯗ�3߀�)�X�/}hNgg��[M{�.;��di��oU���Z�6�nT��u�a���8�:�7Z�UÚ�0�9ѷ��l��̣��h&_�ȹ`ή���z�|ݍg���LUhW�r��=�v��}�[p� C����C�=�����߉��ZLgt�y���t�bM(�)��m�{���Q��Pi�LhjR�y��Wv�9]����{�1\��DE��o����z�ͷn�`���N�VK�4��B�ۊ���2r�R��7C��IM�L/&iR�Uj+�����ٴ��k�A� ]Mq�~dT��7�7�J��ql��ŦP�Ζ�t.���yýn}b6�<ʎP�M�-���-�&Rׂa�����TGk�c=�k -�|w��1�jJ�羫g�2	�>N}�Fl�u��d��X�-��{B��b�*9~A����Zʷ��0\�3e'/�r��u����+�(��-��3]t�d�\8_5:d\o&�n��ƶ��]���Z�yx�=���4����&i]/Se2�1�m�v�q*[�7���n*�o
��ah���^f�W??z�f�z��̝���O�[(�9��$�2v��~��~#{�{G.4^N+.�Ig:.w������κ�O�*.��5�6D`�pk�^�(rW)N���}��OK��;7.����x�Ŧ/7c.�0k}"9�y���@mL��}:ʄWr���8cuVm�C�C�i��"�;M��A�?��\f#R�۽��;��a����ߵ<��	����W)�[}�'��x7�$g��f�k�����LB�V�wKe�z��16}`�d��������q�]���\,Eԉ��������]95'7��=:��ؚ
JC�rv�s�og�-Z�B�cb�M�n��d�j4�j������9��E�䢿1��'䇭�ޡ���ILy�M� ���<�]���Lތ}��0�v���
�k\'v1L%pk��<g�O��(D(
c��M�F{F���^Kir��%Vl%�>�w7���+���ԣ��+P+�l��@����x�LjQ^���)]�`���B%�5iv�"�k�+:��9v�3�^�f)�0Ɨ�d����'��E{���H�f�gr��
�Uo�Y��nO02R�eO�n�{s:F�Tq���֓G����
1t�w��N�:VW}��Ow���D*��U/]K'�����K8�QqY�xO��"�����C[w9���R�)S�jdE�2�̵Mr���0��jM�D�"{,um����i'h��qVRW�o/D�If�O[���o��q9̨b3�T��ט�Y`��^�W>7kk��Iݪ�p��fB��Z#s�D�>c)B�C��3R��rI_��ݰV*��8+a���|MY�h��u����F��]|��ˇt�7��r
���`Mz�p��n]�T��<�m'$[�!�L.6���힌�A�7;J9�����oF�MF�#ě�-
l�����y0�i���2;�Qֲ�X2)!�m���;��V�w8];�q�.�Z�6#W|:���N�y�P�gsޠ���Œ;����#���ƕz٦� (˸����bLe>�9W��Of��_Ts���#͎����k�z�Ym����G['�z�iY�����s.iO�G ��T�Z�[b=�3v���?j�t}Kv�q��u��@�oC�p��봵�f��6d���[r�j�J���,��E�B��+c=�P�.�K̐ⰼ��;���[�s�a�ז���e:��>��׎%�=@�aV,z�Ӿy�sY8M��Z���c��H*}b�^�{H'�&�����"�of�Q��q���1S��C���Vf&�V���*����R�4�l^�q�~��vX ��X��;���M�^6 k0ҟD�Uxeb�Y����v��=W�z�:���{x^��ِ�O t5�s���=�/p�p��ό�uU����~������P/Hڪ�;Ɨ��+�e�d�G�����<_[ï��� �Z��)���+,iKh,��,̐
^��X��pn��N�4^�w^?No4n�4R�FQ���6C�����Ў_��M���{��O6�C���?��i[���X����`���מ��&���P^����:�� �t*_�D�U�y�2{���O��{�7�J'���Ԗ:�te�ޏ�tU�g.T��9L�m]f�5�p��*]��9ƝJ]�b{��/�����g�6�B���s�
��)�߄�V�{�Z�#>c�ᵸ�rѣ�A*H���4��g6�����znKr8.�i�Yv���
hU�DNU�kU��ć:zهn����B� �䕤�X�z)ጕ��s-�ȩ"�����٭R�o�����s������y�R��B�S*��n�mR=�ϳ;$;�l%�xM�)(u��3s��h���w�[�73�o�����-y(/)�o;�؅S���V%ϖ�@k"�#:"�l�w��=�ngF�
Q�t��J�m�r��r�v��N[[���Еâ�3�ۦ���Mp٘�2��-������0�����p�{���;�FQ5c���Ӆ�����U�%R�4 �k���x��DYV/f��(��W�[q�G%��G���$i#�&�#l�ݲ��;�Ԩ?XId��D��p@˔ޑ��O�"B�j����w_T.����4��W�a9
wv�B����ۛEn���\r:��{��D�-�?!��c�E���,|������#�;��-��P��v^�Mv#/N�]%\��lp�u�d��5�o�l�fZۂ��ѱ�wn�;�d���/f̇��LP)E�W�E�?�^���i�=�H�$�Tdf>�������ɿr�L� ^l����=�W�>�^�y�'۷�ow��e����<���\����]��+��Ӳ_f�I�n/�q��散w+�m��UMԲ��d�NR�^}�3w5+{!��C�/�ӛs�;���G��g�@�ȟz˩$+�ju���Y�I���\_�f��Hn��*ʥ܊���n7A�����8�P��L��"(���1[@�(�\Kd�#��W� ��{�KAԯ}�[�S���+š����kg3�<���*#O[�G�V�����{j��D�������$�ɀ}�0��C͡1���-vO�ʅEwZ���L�e����Ȋ �,gڛ���@u�DO(�3��������4������3��6��8ջR�j��[%�8aޡAjk<I�h���m��u�Wt9���[vP���Nt�S�����e�E��O�p�����ŷ���aW��E��n%o5�U}Ukq^�H2�Wop��S�s%�&\P��f���/2̩��8��s5#\��߯!m��0y��a�we6�#����ps����tq=��{n-���}GXό��6�{]���wO���+���upfߧ��G$�H�����;W?j%>��Q�Q&[�2�l6sL��V�6�Xx��ٻ�]f1z��\��L{p�����:I0JCe�V7mY��<y�E��QM~
[�)��=�we��ĉ(��̰%F:N�ˢ�3����dñ�Os�6<�Ԫ}�DV^����F�A8;.�οz"�Ў������g[49;#M2���������s�&柋T�tMµ���7w���呼G*Y+h��Te�w�L�C]���_�ל��r(Qw�@�L��C����u��]���@U���*�*�l��6�u��F׫Z{�����n�8ɭ�n��1���D�4jVf�ͅ�N�l�fr�7���� �ɺ�W)1L))��Sg��-Շ,������v���%tv�ӡe�Գ%jf�1jJő�򧙩��f��Y���b�̧�#LN���ku�!��|y�Jz�E����˅�t�=&�����_tVV�O4��-MF�k�������|ܒ6^N���"a�i�����Xh��T\Y�u(�o�e:[0F��P��3�����zuN�a��^�
W����d����Y�/)�g;.�\g��`m�%I�1�;?e��ō���� ���|�����Z�#���}b<�6D.Ɉ(�������j�X�5vt����@gA+qs(����]�Z�{X7g������2�W<���[���}
��*q=֯A<��-��zR�3��'wO�y����;Y�Zi��5k�}�r�W����U�즟nޚ��Y'fUl�nٲ6l�`�H��B{}�v/��u�������Kt��`��yr�S0Ԟ�!�[�vӾ}p�^!Y�|�tl�.|(H|�h竆۟�'�RR��[���<�H%�Ghal,�C���U�� |�~��~����|��clm��lm��|������N�l���q�=��t�c{;ld�`�`;� �C` `{{�& �`��0aŜm�ww��xm�����0mgcm��m����91��v�l��m��m��g&�l�m��m�[� ��n�v��Zm��9  s���v�l�a�m�s��g8�l�cm�� Cm�� �l�6�9�m�� �m��m���l�cm�� 9��v�l�6�9�m���l����m��m����9��g;m�s���Cm��m�rlm���p9���6�p!���[�!���{�_��9 �aq��P� �o��}Y����������?��?��� ������r?_���?s'����~����6߸?w����L66߷��cl��3~���3�������?�}��`�X�cm�_�o�=��&���1��0��>^~?�~!�[��0`��6  &@�@����ll�����!� ~v�6ŀ����m�p&0� &ɶ ��B߇���N?�����L �e2�m���0/��}�o�
?����`~'��}f1��ۃ���;��g�w����?�-��=�~���}x1����vُ���>lm���@��o���d���1���������cm�����<A�<��n�?�/�포�{;��8 �6��?f���g����6�p|a@��=�@��q���hhP8��� �4clm������6��}�}~�����.>�|}�����?i��_0�|�����|}��1�����������~A������������ٰ��}�B�{x`1�����|��m��X>���d�MeB�[Qf�A@��̟\�����P�(D��
�����UB���0R�Cf	)-�%����֒��D�IR��R��H�D� (���R�R�U*��JR���P�$" KF�:�R��U4�YT���ZD�P��(�U��mP�%R�+�UH)	
�QUW�*QH��PR$�I
EUBP�H��� ��J��J�)H�HkE*(�B� �E%U$Ph�R�%UP�|   U�)Jm� �h5)c��l�Y�(i@6�6�@jD��e�U�`�)4�@�-�	hZ�n-�&����p{�R �HD��J��   ���}��鮅bE�MҤ�Olm�D$[�WxQ!T�B�RG��z�2[j��0�"� ���T[-cV�cZ
)��1��Vm��^�խCA�m�h��-JP (�$U
x  �{N��Қ���KΒ�`fMTҀ�5���Rb��������`��J�v�5@�_fT��am�h���T*���THI)J^��   a��`b`�-�-��m�6L5[*e(0"�հlL�(4իU-�mA����Y�օZ���ح��j������A*UJ'�  gU(5����hb��F�{�� Ci� #P*�q�qS46� 5�w2T��*D��ҡ*T��|  <PH��m� Q5�RB����Z�DkZ�TT�����k#SQ���4����� ��UJ*%UU*���%�  t�-�"�Q�Z�*e 6�cU ��Z��Q���6�Jl0PP��b����ps�J%�I�T�턅@�4�$�`�  ���UBE\��JR�J΍Ȁ�]���wvjI)�Yѫ�)D��B�Up&�Q˅�Q]�:��U�҆�AI.�ƪ �"B�T&�%�  �R�(�y�Lpm��a��$�E�.)(�T�Q�T
��rGp�Im����S9s����1�� �֝�n�"�r *���%QR����   {�)(�8�H$W���R�v��SZP���;�P�bX�RJJ�����Mv��-�eO���I�49�gT�(�O 2��#5 E=�	)*Pa2 US�h�T�z@ �JT�  !��� �Q  h �)PLUI� hf��x���ߏ*���l��nם�����a��`,}�\�b��J�v/��_U}�j�}���`��ɱ�m���0l����cm���g`����� =�xxx����h#�쏓f!���4[�|���H�S6�%�^��M� 0|R�j������4�BTZ�m�U�Y6��k*S��acL� �y)ҭ�N%���Lj�UgPOL� &u�ͬ�I�t�	[�eϲkw���E�*�j�+�;��D�7I��b*f�D�vrQiͽXdH��U&�	��%H/h4�Q��ذ�I]�]��yj�\�MSr�Z-ڣ�� �[O4�a�ʌLH����cm�ы˚����F,� ��^�s@��2���F�J6�t7p���L����7H^�*RB�Mf�keoM7y�wb���х�r3��.Í�gsKU��ܠ%�����R��WP��R��XǫNK�V�1�لEM��Zl�b�U��iu���JčӨJ��z(�7���հ��T�����:��V�P��TkVRԅ�K]Ll`ŭl
4���pVM��Ip^&`+)������N�A0�֥������]���%D&�!�5��s[�nc�{-�y�ٵ6�K6�%��yI���j��Zt �)���KʹU���d��������x�PQݡ�P;���ٓS�ckh-F��O���jVB�FYlR�MW4^`ee4NK�����j�SӃ4>@�(��)����#�f�L�ڐܽ��ҭCi�� �c���x23����d:�c.�] �,m;řCE4x[̼�V�-&���wZs2�ƥIJ�ɹ��b$E��?�JPX�d
Ƌ{�֤f �˚�N�x�W(��̓{� ͙���(K"���i�r��yw�un06��B�iM�H��5*��Μ���������+uWR��3F�{����<��*�[���@8MZ�r��N͋Ux�;���u����ِ��rQ�8��[Y
��w���S3�"� 8c�+���{�ѡK*�HP���%h��]�Vn�P�)��d)fX�@^l{�gE�ĪBK����iI�i������cLۭ�0ŗ0�H8��`���f�t��U�VK��A�씪;j�5lb��ƨ
�p�J:6=�R��'CMxm�m8uK@�aZ��	C7�W����V�VI���P9b-ܬ�����ɪ�����;��2`�VU�!N�h36�T4a�.��YV�PR�u�ŷ�aF3�����a�5u��fW`�L�k��1ݎG���5-��S�K*3��Xջ71(s���i�������V�J�ݓ6�h�[�k�7�E1[�Sv)�vV��a��]݆p��L��"T�w6U�S0L�^�i����	Y�V�V�@�xkP�!�hC+r��툫~�!֢���0j��H�$�r��kM#{Q��#:�+pkW�z���%��m������E���W��+�t���v�/ ��\z���eh���0��Z�����5�/)�u��\�����e˖��q�r�2��K�|�(7v�cx��[��1Mq�� ϝ�CAf˅)��(4���y�i�·K�V.�sY�̒��9j�'W�Ӹ����.���2=&QGw�M�
�Vf�`���2];�5��K�՚v��Tq3�l�X�NdW��wi�+;�a�4YΑJA�JШِi�4+�
�xB��с�en�[�.��e�u�S8c��Hr��U b����:�H��mѴ�7Z�ܹ�mF����F�E�ZWA,M�z)`x���"��0YOᛶ��JS��4ֳB�TW���(Qֵ�WB�nݚ���K0@-yZťPM����)S]��c*��dt�h��+��*
����:e�	�^�Mcf��u����m�u8�WK.�
N;�*[э:j<wtsfP-+��򃧐XͨD�*��<��[Q:x� �Cj��y�l&����2"R��p&[����E0j-O"B�,�#(Jq�\�&���ڔ1cįD�iCO�p�eܶ YQei�,#7M� V�[�ʳrE	:��)����%���QW{��,1XVJ��{[�ik��G
�zI��Kx�ƫV&S�1:MKZ�ca�#�R��՚����ȟ.��~�]j8kcjӑ�&,�Mx,vm���
��J���'lBl�l�P,m����Ȗm,��kf8u3U���Md�LWVLSCzH.�qe�ƍv �6-�B��t��#5&�sxĭ�������ͭ�I�¤��xfIlmݽ��x��5o�Z�V�����U4CPӵ��d(�:�m^�m�0�n��W��]�بh�%�0� cm�����z�� �l�:$��C&��Z�����(aD��B��`i.�a��՗����͵P�սYf��C�,�X�;�@з�1��%	X���(^�X�����^bf��1'�)w���6�`��Fb�:m�[ �-�����L�9���j�p�;' �kȩʖ��+U���ҕ%&-Z�C�v؃-�*����12�h$v��3/u;8XճX0����R�*�;N���W��6�2a�j����!di��z����~ŀL�0ҩ--e��ӷE�)��6dW����J����H��ve�{P���;
@��n�e�E�'v��0X�5V��㬒U�M�MZu"�ZN�)���Y��MEBR:�ְ�� �iet���ŏf���{qM��Don�t$d�yb��#ʚ&��Ae�S�r��vF��f�a��	�fZG�mXq[jc����G�A�,���ަ$xQܭr�\z�T[Q�.U���#�uVeGVMktK���1�[��E ��zV]�2U�i�W�X�fcߜ&�
�$.d���ћ`ې�!���:�^���^��0��v֦cV�Y�c3r5�CjЖ��N�«CSiZx�bF�]���6PdV��Sfcd�(5�+LT�.pʺ/ς����;�Exf�c3Z��$���I�w5)�4,��4n*%)6�ۭ����شꉲ&H�����̄�r0�0T�0�81e;���m�bଭ�F���,�@��a8k5N���{�2K�re�&��Ua:b�����pk2��7�=X�PH����J�lۥ�e�7���|UnĴb���/1��4+� ��)�a�ő�$�����7N���%���AF��>I9��J�&-��0'kS��wKjѬ�MD5(�bI�6n�ދ�%;*n	F��"�+ݭd�(=xp"�<�������ZZ��6�B�te�{r�Z6�M�"�E�J#��fn-U�)]$�� ��[Y	u��oҕ�8[�P$5TY�l�P��nɍ��1{����d�v���Z*��j��[�����c�xi�4�dWa$��0,�oiML�x�<�2=��;�.����6حvP������:"d��;?-e|��5�𜍜:slD��\��ƅ�K�i�IX��uǪ�<l�}�'�P���i*��>[H��kT�73U�ԣI����  �װG��k`�mR��Ŏ8tjtp)R��ˡE�A�Ku;�4�*M�-�v1�	t8"j*�ݬM�zR�5�A�X׶��T��%���a�Vk�L��j�	�Y��$1�t��{&�ˎ���!@�~ͫ�\��ʶ�4��Wr�n�j��f�p#JֆQe'[c�t�Ot����Ww�͂�N�h݊�L�`[	1A����Fe@��U�[���rb�͙�*��⛈��
���1�t/a51��ۤ	7PnժD��3h��ɡR�E�	�l�v��6��HB݊��B�(�E歽
����1V�޻���d����]�Su�3@�[���-k~dd"�=&��)WF��S��I�
�:�J��	˛��KY.�6:-����*�R�yF��`���2�Hk�iӰv5K��ce�aL��42
�f**�V��mj��Z��5�Q�t�csl����7-R�ժ�Txr�{`��P�n�RT�f����Xx�[�.�,a��������:8����u�3���
��ź�*J�0�r�8^����^������a��n=ڐ1���e:�*��׷"00��	���c�5�i�
�:�A�O�Pf�,��H(�H�r�Tu�D���_C��7R���%ӵ �LK%5�6��z ;t�+���/R��ǶBi�˒��C/Du�5V��R=D5w���cgt#��	��*���js�dٴ)�p���H�M�� 0�;�m�<���I��3n�Y��1�t�ԥ�V��^+3	3�@:@�z�ط���W�t��N�)j��2�J��C.A`F�݀kjU�,wVP�R�N5E���n���Y��Q�L^毎
��{��D��)��-�s7R;O*�Ef��f<�u�޽fMm(��L�VF�෯^�gA�S�U����6���aT)�+�u�ӎ��������Ib�t*����,ִ��9V�]�)b8�$T�!v�W�Y㲮�E�1�2�'3e��\1���ϛ�Z�1ͻ�VN+��wshS�͇n�7Aa�a�����p�'�r�J�,K�S1QwL
Mk���-6l�oQ��"�73b
Wc�7�2�E�axx̩�Y���.�2�:�Qa�e�V��i�i�tO�;�[o!&�"�n��Z��@\��M�5IZ�&�x�5�[�B5��f���J�`�u��VTj@3DX�� :x�t�*�V�ݢ��j��4-��JG/�Xc�F��y��F�ِl3�'G1;�]9�v����:���֚�YM<A�q��9���"�mڹO1����S��Sy{�����]]0Jt0Ӎm��ANa��^YS���'ZE�F��}�1��-���*�MnF-C�-C%e�:�+FSBx��FMf�Pӻ�.�Rɻr�2�$j%b�k7L:IIBM�HI��f�,� ^��q!��Y(��0n(�Ƥ�Y�w��-�G.�̺��ͱ �v�Z�@���]�kpv����)�Xt֗`l�����0PUb9�ȷA47���0����(�Y�f\��
	�	����Z��Z�&|p��%ⒷAۋ(��}���<�ʩܩziU�U-kc�B��[,�h�j�J��՘�ټ��4�Ƣ���^��%<b�*+q�7���m��jZV�MM����tkrA�ƂO�"��`�{H�0�w��"�X�ґ������!���eK�v���\Q��c����Z�2 �4,�G]k�,l����m�Nee@�m��E9��&���[��al���Cr��P�ĥ�,IGVB�����4Gv(�4u뿘,
����J��YA�9VV�͙X:W��+U�dg^]���i���;m�k7N�꠱bU���b��0�`�0�ŌEu7-J	t��M��_Y��G�Q���5J���3	�%b/e�#���7���*֔6��n@�`��{�<y6b�N��ϙF�3Vb��w*��[�*�7���e���o�+N���7�$�u3�T���w�u���(��\q�:�庰,�ѸU�b�f;T#�l2i��i,�,�g,S��Mܧ��o4��
�jYw� �>�,
��ݔ�m3Q�Sњ&�B�e@2�h��t���P�Jޓ�N��b��2�R�0Ps,6���&;��/Q�y"�{�Mq��ۉ�۩��3�Xke��Ey��'h[�jr���2A0��\d��6�+ak�Ot՝�252C�kQE�c�4��#F0p�E�ҩ��,��MN����
ȓV��dV dJ�;ON)�7�-e�%N���$������P�V���CZ��iZ(�m�6�LLnб0�v<X�H�g�t�p��u8u*�t��4˩��C�#�M!20%d�4HNYuU7*-j��^�Sv�q�;V�
G�i9�2���+e՛��֬f�eӸ�խ�����3pN�A���۴
���h(f��� �gG̅�F+b�� ��$Uts��vTԐ�q���.�ǒ?���SF��B��j�wDj*֢�ͽyP��a$Ee��Dg��;-�m�y|i­�&�.(嫣n[�����;Tm���nkޢ�Z��dYwD�z��N0���k���_+�1�R�۵N¼�RV��n�<eHXUm��A��.܇L��0������Mƚ	e���>6��zU��Jj��8��T �,=7����DR2�]���Ǻ�����,�6I5�ub���&���e�כbb���t��q���9Q��M��âXx��m7��D��C�)���7�*Z.�`�^BFՕb�U�-�*�)�H�[��;�$z�e���T).�u�oƌ�9]9M�6�(�@�Zq���W�4V�A�:ڎ4�ō"��U�Zt���fTc`��8�r�Ҩ�
Z�j��'s\v�(�,{�jK�W#Vv[s\e!��ZЌl�2X'�yf���L8� �M�R��;����z�ɣMq�ںNƭpfKg.���������&��ؘ�k �`TV�{�,P�Ck-R�[On�݅MX(��0��*8DL�%uceN�ȬK���A�8f�A�{��zrM%2;���X�L�*5�Q̳C��'�+5�v����n"Ἥp÷��C7eժU�G�[��7�#� Ɂ��@�:~�Zs�V��6R�K�1�u�Q�l��RT�������w��Z�t�wY���AJ��b�d��%���!�2J�R�
����y�F6���ݗW������f��gd�*��8�����%6�ŗE٦�f^e�mf�D�]�?wo)x�Wjw;�gE��`��v^d;I��Y��-i��#�ҹS��{�FJ��:�tÜ�x��ϴ�fto+��6V�Q�:4�*n�Ԡ0���IW_:m.��u��������T�z;vc��Ekm�8J��L#�a:��sf�Ù\�J�O@7$][�M���a3�Sڛ�E��pp{V/,g7�)�`ue��|���ٹ>ޠa��ξN=V��qPV!Mk�s���Ր�-`828�AC*�&����1���r��; �8�)h��Rq�tA�/1����s���r�"�(�<l�+FAO�2H%^�G��r�S"�3��(WVY�3Z��)��|S�;�/a/���h*�H���1�gK��ز�u��WK\W֬��)�̇3�T��=ٷ���c�X�Z�{��ς�l��Hxo0��D�{���w��f�*[y�9��6�[�vR�"�$�{K�)��'#}�q���Ў�r�L�k����;=��swL���Vҟ>�����"og
��A`�qWE�̭嫻lR��Lܽz�J�&�QV��o�21��-A���^x����`U��{bY��I�9�֗+r���w��+��p"�����[��^X��If�ߡ�쏚]�X�oY��V���K�eljt��x�[��n1ǳr��A:����h�m傭��j�un�<ɨu�W�{����70b}�sTL���bt3w����m�����2�p
��129���>����uխ������+/�ݫ�К�o/�HN��m���k2��?u6�:3��v�(VѱhB;�N$ ��b��ݢ�_7v3�l3a������Ҳ�Ԣl+ܠ��4�)>����U}%r=x��S��=�h���;�ǡK�c��Mfr\�(V'Ϩ[���{5EC@t\�1�fr��p�"�j�ƈb�9,�k؎%�ܛ/_�>�o�X�I�ղ7:��Ҭt�@k���X�O�_*�Bxe>�ųkF#�V�`q�F�q����A���E��i��+�ՙ���w�9���PJ\��Z�aiwc�I�9���LGWS]A�7�u�r�!�����8���Z+��r ���>ױ�GD&��W�F��iÎT�N��8%)򾽩#�u�^�+n�}E�r�XUbn<�F�f�T����+v�`Rbv��41����s�rIS^H�WD�`BfU��Jj�齂k���|)�.�[ύV��:�qU9��
��X5����i�
��$vIy��b��f�4B ��1��"=Je�l�!
6���sj����v"��ӷx&Q��;�`U� ���7�7zu��i���d���B7���/�7�����Ԉ�(�з��c-�.��4��h%`�Y
	U��C\ky��Z��*7Qb⵪Qw�J��\��H'֚0%����U��w&���ٺ�59�%��y�˲�@���qj���꺆޷ɑ�6ק��B�Z�cxW$�VV�E���;݋�{˖I���|���:ufmje^Y������K�!X���:�A��
=>YP;t�]mu�a<�or���ы5��q�m[\N��.�Wt���Ç�N�}fVZaw���KdH�YÆ��%ݧ��.+�*R|�fY�0�-`bS�s�F�x9���Jb��|����5Usl3�/h��ӣ�\��[�hJdsxG��+]/H��O욗&gTڄ�Ñu���_0�D^l�/�/u��V�S純a�Ǉ9��Ò����!��Fv�n�=��h�@���Ǽx����Sp6iY�Z7q���i�U��B�osV��i�N�u�}���ESx���E�Ly�%3p]��Y\���,�`�QB�5gaMh��
��c��V*y-?���W��/�P��Xz����KCxA���Br���K�gc��=�MM�t���>�2�}��rF(�Q��X�l�5SCC1�' �z�3�gU-z����O�S|����=sF�A�g�w3��n����Duh���Q��Rnh��/�M ��Z��y)�[BJ��6�ڽ�֠��kS�nc��vor4����k��'�9�l��m�&]EY��TdY�M�X�sLS0��k��y��b����s�.3�)���2��w�)r�r4��Z���Ի�h�i�8��{ܔ�r�n^UtS����;���Y3RG���Idf:�0N�����^Qաd�)]�e�{2�>��k.bOV��)��P
��0���;]�#���E�!+��+R��XxfgHKF���c���(]u�s/���}p;u$���6�b{D��Dm����>�4���2�P��u�Q�K{��
KjUǝ������5�X>���!&�I�1+xL٠u���Y�փ*��t�K�⼼X!��\�/�J�F��v;�U[�.|�[�e��4�6�W07�W1�<��^g�� �ђ�[�H�aU��i�x����%ۡ��Z]�����+���+�1����6��*���MpP��s~h��-�;�����^�����h�{�wĪ��P���ą7��U#+�U�e	��s�$�����{�,�]:�.Ȫy���.�nup�/U`Xxvu���<�]�g�/�ll!ڜ�me9J<����_����ݘ�8Y�C��̉u���i��� y��X�a��Sf^��ދb^��[�1\�n���1��W�]�wgbEb�k\��`�M��z� I!�kV�]r�Ep�z���	�-K&ٜGN�&��Wj@7��r�Zx����Ͱ
qU�ʙ#�}�M�/V&�R\���{;�'��m��z6��ʘl��Tٮ��T��?{�@ڧ�>؃M-{gaP��:�t�:O.�Lt�h]s.͜��a��RK��i���m���\���S�p�ɸ�EƷ3�N����+�Q *�x�H ����v���!ƳRG01������u��(t�̥�3YB�4���vLI3G��=Υ��M���қ��ԘEu�w3ҧv@4�B�Mvf���Mݧ)}(`=�^#��b��b��5�v����ф�Ƀ�����k��8l	:���a�����ع�!/4hV���q��F7w��他��ȣV�n�:���󉄀���m�\�
��9+a���9ݰ�Mw�8���N�q��	�8K5��k��#6ۋ��ۈ�|� �ѻ��V�1�gD���T�`ǜ���o>+�k�%�����D��,ȺWT�P[g)`d�ŝ����Y{z�̗��U�>ۋ}<|+]!��N�3f�ɊH$�f�ΑC-vʡz`�Go�?�ێJ`H5�7,��;T���S�r��7 |\�ب�h�����Ƀ#+�5+OP[��8rbX[��J�)%��o_w,z���t�-dލe�:�U��[��E�,�+zܐ,��yTRVd��d,y	�I��b�v�����n��I �= ��6dݾ�[����5ԕ����灶��ᕁ^�իS'��dR\�Jcxe=��ժa�y�{5�}t�Tz��h�]]�  �;��cv�_l撙n�52�5hmة2���hb���\㓊=�):��������PKi��9M˹5ӝ�v� �α��GY׫jd�t���.6⮨��s��j�ܸJ�h�	��_MSVD��fg>X�])|15}c7l^��u.��dyǵ�.�L6�����V�vY��X���|�ۙ�4���N괰1>��f7��@�}��a}���	�������ո]��B9�صn�$1�y�J��ڼ}oaX�t�K��\A+�K1[dZo��r���Zx���[�9O����/*5Eu\I�Y��P�����b��G��P�D�E�d|�'/5갞c�Y�3�O��	83�q閱�Z��:K}%^�����1�Jr���/8dM�\+,�Ŗ�3�Ym�sk���fe9)������0��l��Ӝ��o&�0�j��l펊Ed��ܡռ:�d-�37yp���M	&r�=h�6UG�.����%5���)�.ڊ��v嫥&��UE���g�k2sٚcب_%R���J�>�㯳j������e r�D��-�B�;��{y�5�c,-ɦ� D�ȭ����Z�ΆZ�K����c��]��t�+��;�mEZ�X�r�o�=[�֮ë�+��+�-�|���|{ӯL�{y�.����� ��!����K=�CO��%2O^&W]9N=�Fu�U����L���;\�h�2�G����E�-����J�p&u�Ŋ�]���O_7�D��yWxj�sHk���ר,7ty�k2��ﻀ�RS{���k���뮂ęq�y�0�@�f9
��¦p�_61���Ν;鍘�n��9�<�ц1O�^ �<���ҕc�hQ�o	C/RN��J:��K���:�X'm!�\]�=6q�������,��ъ�M��a�H�k@�[�)2���:f�U��V�v�^^t�'tJ���U�4&a�=n@�௥5��u�m^�t�L�	���=�ՙM[2�=�j�nb��V�����An�,�����%����Dm�X_/���kU�p�&�R`r�5�t�ڃITޗ;HP�]�m��(���̧�e;+���c�����l���8+���(y�ru�~j&�.�ݱǟe�:�Hq�<�\���r����8v�B���s���	��t�}���<�7�(�-����A�TS4a�ﭶT�I��SZ�G��^��g]^�����%�ݯ���y��IBd+����X���ݵ��-����s�k�P����Q
��B�67g?>ª�NF�n��;72���o:s�<%���(`GR}�c�|V��vs5o���EQ�<rj������d�%Njv�;����k�1T����o�pc)���gz�%�es��K#�+��r����b��g����QE�a�eA����r�V�U���6~YáI��8��ˇ^�P���r��Xe�r�}]�iggM�#���j�����5m`iV��ӧ`Ɋ��^m.�94'V����Rt�F����OB���
�RfL�}���r���I{;�"�k����7�h�eh�9�P*gkT��e'�$�&����C����i�k��Ů}w|&���de�2Z���L�05W���Kn!|^��=�8���&���6�=R�]Bi쬰�Fs�i�v&��O�ʍ�3s{K�������7�#�5;+���g(
ĥ,���{-�s�bhU�1�5��8p���ۛ@X낓v􊶟Wr��O4��J��P���ę�Z����i��=���Θ��E݇+xg �+��<�n�v��yA�&��F�'2ܨi@���̳�*�D��u-� �&l��YX�_#��*U��n�xg�b���
�������p�����|o��`ym��0-��)� ���1���3��M��.�Tb�::[�5����Z�I�ƀG~�ت4�S�hWe���� o��i��?p=ٙj�p���^���zA}�3��Q���V/-���x41�Y��}rg4����[ �4f���W5��h�X�<x��z��|j�Q|iuf>y���_t�s�)�r��M���W����_u�)���N�뼶eC8��U����X!ͪQx�AWA��<)Ά��7tO�K����=��S�6��O+��|D���F���̨l���*���{��4[A���3E�Ŕ���I�f�∔�٘2���Գi��<C|��0�k�*`�wد��B�r��@�mV��3C�nCG�H_U�Ǜh[i���_.cb��]��U������r�7��!��J䳚�&Ι�hM����_G�\e�鞝�題K���i{0򅹐�e���N��fv
�Z�Ā/3|�V�*k6��c����c~̀��3*Ү/�ve��cr��
'!e��:��oV	�Ҧ��]�{�G�s�陕;7{;K��qT�u ���Sq��d�����E���QQ4�^̭{V:��}o��)v�ݭ���D.`����+�p}1=�Sx�z����R�=��5)�A����`��wh}�6�r����TN�]u�a�C�o�H}�N�}��m��! ܆�;P��M�� ��ƫu��}jK�%�嶕,��&��>�ǲ�\�y�Bj�W@�ѻr'v�U�P�����<ʧ�!ٟl˶ˋ#��� v��,�	����2�c	Z�E�Ȭ�:��g�^*v��)�l v�䦭�|֜��4�:�\��h�b
�<�,ջ] NO�z��� ��/ɹ�c2�.��퐻�	�gQ�X��i;P��Nȿ�:�;:��oS3�Q�Op[V��F�,�[_=Ϋ����l��,���9j]Lh�Ҿ|���Ն�5Ǔ�Ցک�`.#�us;;�f�b����j�rK`.�L�X�9�t�m�3J�R�y�u��M��W���pV
ي���.�ZtX|]��ӋK�k�*���p�j!�J�WM��-�3^ȭ�v���]B��jN�i}s��tq\>t;::��Y(����	>���p�=S#�$Ub��:�5��;vbi�S9	Ƥ�}�O^�e�����f��@�[yuq�c����p�`�>?���ӱ�M=�!�Im�1���E������y����w�;;B�8� $p���|8R롅%˺Ή
y�7]��ќ[���t�)V�̚E2w�Ԗ��m�+3M>�Ҧ�gZ��:�T<Q���Ӣ&�k���`�������Y�̷ʺVu66+Vqv��WB�b�Nİaxr���Fd��=rl�G,�����P�JYηy��>��&�B���3N��;�	�ۂ���)�=�P��b<����=[2��S�⺝Y=@�e1˖N�d�.���F<�;w��PpS��\i�_S]Xln��4..ҶN��������W����>������vp��n��3-E����U�cGV���S7��u�JT�n�	ε�.�pA��yX������@f���[trP�����X�!ty"�C{D:��5z��s1�g��`�G�}R�Ԯ@�K����yb��Hn�)R����ǸɱV-Ч�h!���\���:�U���Ɋ�=�����)Ы
�厩�dL���J�sZnJ�ȱb���L��Pw�8V�����,Eͅ���!yB��4:v�z��+ޭ�b�0�v��W$�)�ԡ���(�
�wӞ7[qMJeon�x����0��oc]ꛦ��Ȏ�!=�}��	�6L�E:��۟R�ur9ך��8.L�X�6�}C�b�Xώ|-���jmN��n_h���'Yv]gJ׬؋���K��Zu�K�lJAj�"xk%;������M�^h��8����YO/X׷$np�-�F�9��>�%
�*�Kd!��v������R�yݢ8��X����Z��.ɪ+��E�l��r7�;��:[Yƣ�~���YɣЮw%��V�*K��ȥci��`e��.�}j�e��Zl�_�^�X���X��q��iP�ݫ{����V��s؟vf���f�o�A�k�ר�P��%2"j_�!��������D�N�B��p��n���ԭ�:�֪��}�Òq�PhM�X��'�L�ș�c�G�*�\rBe���� nKu����Y;mo�!T+�⺟ͣ�]5Ec:nk��.��j$A�SAw�
j��&�+z���x �����ܷ�[kD���%d�"�h���f�Τ�{{�d�4��O���6s7;���Z��n��2DjY�T�^�Wv�g��p���RǗ1Ggd$<��MݦT{0pV5��tU��Δ�>
;`�f�у��k�븣�6q��u�K���&G@���ۖ!�\��cb",]�K� N��a�B��[˹W7E+c�{�ty��uB�k.�lRc*h5j�ݼI�ɺ�ҕnL�4.9�[8/V��h�a����f	���[_#��v�Ggh�w|���.�@��6m�"�݁v=%v#� b�(d����@�(�&	��be敐�v�&3�r��۰�Yi�{���wmb�+�
RԮ���I�*�h�<Փ���ˤ�9j����p��X.�e�٦��e��*d��k`�p��z���P<��1%vj��r"��{��j�9�)WAԮ��l���߻rA
fE|1��<R��%��#B���LcL,����yl�)&8uI��7n3A�mK]a��{EuaC�7k�\��Z��'�[���g6���о�N�Ae9Q���NN�c'EH��t �j�{�oz ���ީ�)�o��r�O*.v)m�N�b�
�]gK����Y��l 3�v�:ͪ�
�6Q{��n�+Uܷ)�fp�:�].�-�N�:�t
]mn����k�������H��\���]:n�0t���.�x���椝�Y�s���ݷ`dF�F�2f�w�t��i�����J�]KUz���̭q`�W������T��w�	�}n����;��B.��ͣ��
6��WJ�<����m�mi�ބ��8��QUdéP�2�-�uܠ��o��m9�jr�N�8L3$�C:�H��'��ȣgod0���H�N�uٷ�����A̻�ݔ8̦�=����wۄ���xm�w�D��v��9�ʌ�׈���b�m��)vUй:�#�����w��	�y�]���KAօy������/��	&e�*ը��|]���L���l��|c6>+�?���0]K�}�E��m����zNH�<�]��MC9��&������,��˳�!;1�uw=���|�O��.�dǌ�=Z�^� �|���O{��,�9�i�i�<�ej8:j�;}[1:�/�h���I�fk�ރ�m�P���XY�)�>]�;o�5���D��	㽎r��j�K���8B����'P\Vm���|�^7��9������,1���5%_bڹ�<�1}�
c�R�p�)X�8���S����� �h���yq'����hfK�ɼ�[OiA��� ^�N���z,�;�V��K5��(����|�oen�va�j����;��N�U�dS��\�E���q憛DEN}�1O,�eה�M1N���v��^�z��c��P���Vȫǒ^m�QEXY��l�dZ��5K	M��-�:��)Y��ZơRc��S+��S���ۏ0m<�nt�.�n)�a_T�5s�@t�����g\��=V,� l��v`_n����)��i��b�^�Yq\�H�������E��R�nc�m3d�\��/��[&D��-=O��S	z't͜�ڕ�;{^jG�-}t7(^�]	�1�z�0r���m�jŲ�����hu��ljQ�HՅvq��Z
�R���U��ӗi��;��ηA��v�\@wv��RKkT�v��x�z���9����x	(Z�(nz��(�^'j�y������3c�W�9] �VF��o��wz]�kW�q�N�4��QG�Az��b�v�f�����l�J�٢NsO.;�gR%k#)�I��m;�$㺈�]���\�1!D�TeW!]�Rt�t�ǳ�A^��mc�!8fՋs:M�Щ�	*F��7i�\�4ĥ�K���e��H�ʴ��Xu�΢��+b������VWev��b��/No:�zSMk�l��TS�asR�h�֞x��R|���_c��3|�p퍃r��k>�\;4�����Z<!A�"�u��[#�#A��+�HE�;W!��C)�Ej�oZ�<�Y��mem��7T�-��1���4+�;�n���c6�]�,"F�E��X�K8�40L"�c���_#H�|��{�q��.Vn�������ʩ�g��2��ȫ��Y�q�S�Z�ZKh��v��8Ұ\�*�x��w�bvL�%8�ާ\Gj���ȶmd������i-��!�'J�Mv�ނ��:9:���/��_^�����9Yw����|;J�S�������*��]��,�F U�
6��ˇ����6�V+]7;�SѝX�� lM�^�0�Ԩ�ײ������ɽ�r��*8U��U�M�����}�oxM�;}m��}��V�X��v��уgB�g���}9cHh�B��o��.�[��X�f�v=�����0�ꄪ�%��Z�h�k��2���:��N5� �̷\"�__24�П_2F�[@�97z!Lu�dm;����|�͇�4՘{Ŧ���	l��AQ=@.��<�i�(l���4]݃���1��aƸA�vK�8+�MZ��-�ZnU�.�q������V��_d��\L�ZH|��eKUԘs�r�C����P���i�I>���|�m�y�*t*��[{����p��b���`�ڲ��$�˒9yR`o��Ү���]˰bD�J�H�\��M�&�x�&�=�3V�\u��V.Qd������[������G\s���<�Ү�hS�	�+3�8��ei���X�aBK�K8��p��v�gf<���
������gK�1u�ےЦhL��l�M�����ƕ���R-�;6,��	*�v��]��7�ҽ(��Xk���յϫ( �	z�W�A�ku� ��ܬʜh��E;ƶ﷩F
b��m�-g(2�H��b�'R=}ܱ#[3o����~ժ+�#��,��`���������0r�G��o%��X�nY��j����]��f*��d�q�1G���Knpa.+I�Vs�ܾ4�ʈ�>Z�	�
�0�Ǫ�[�j%h��h�Ł�*��B*˝wBei��ʟ��4�˾�(i����B�g)��5���Υ�ۥF��l�`4�5�Χ�5�z��V(']Ӄ.H{�g`�.�L[�"�%�Z�U��ɦ�ufw=���9,��B��]��7���4Alu9����f]u��`���5�L���['pn�K/�.⼨:���R]Ȳ�x�Ճ��f��v,6�ͻ�mD(i<��8a�\����L��v��}��Z�j�{��+h�n�����,#s�ɛ+]�Aᠴ{I3W��&�rΛf��R�p=���%: 1�x{.�9u�k��(�m�dg!]n����Q����&3����6�okf㷉e���ʉ-��_;-���x�8"v7h`t���t�x�5��T��T��r��͇��֡�3,��Xlm��ht��[�O���գL��m><Va�;��hF���;� �ۋ��P���`ެ��V��FoA��I���N#���Ǻ.獛�Q���f,��ja���\v�G�U��F���B�6�J���F�p��)]����728�:ڹ��ky�K�xx�+ZwuJ���q�I=�Zo:@���>����	޷j[���N�
�,&]������#��/�:��`Q�Ir�ޝ����v�"��{��	� 8�8��]��`iz��E�6X�S����w���s	m�E�=��R���ȼ���׷k1�vۥ}�4�6�<�ۊ2)�=�˄ed��R8�9��ʴ�Lr7.�HZ�SL9��WV��z��������+�l���I[��|��R�jĳJ;G�SC��h��w�n������*�d���V�9�|s#��q����@�խq�7�K�����Z�%�o]��f�D'S�u]1Z��m������h��R�x܆�aM�q�|�Z��M�U����:W�
�
�}��Ut����b7F��fJ� �*<�T�x�H�n`�g8�I�٫мHK7��0K·!9�\	��:W���j�̅�U���f���%���7��X"��jlK2�qY�s5�ͮc^�6��tV�	�3�B��+��K���)�p�1��Q��`*�%V�Jas烷�3�Ẕ�GhBJ5�x�O�Qw7�ۙ��C��sw�cϹ^�B��E`��� �5su�/kM��ֳ*��͵s0Y2��EZa��j]5A�Xo�p��8n��8j	��ٵĎ�q2����ʃR.��店�]��퓻�6�v��ui�ʋv�9�ij�c�I�m��c�v�S�*@�]�j6$VA&�U@n�WRb���֕] ү��\�t�wk';�egOi�:�R
(ra�t��(p����V�0hk�nѴ�]:u���U���DF�(fJ�SJ�OV�f���p��S743�Ļj�(����ֶu���ʛ�O�R��
�v�M�s�lWE8V��Օ-pf�Ir�V5#�;[s�`,#,�8+r�8a��b⧬�_Ĩzk�]�n� ��yiਜ਼AXh�k���=.�;:,�O(]�v.u��-��R��r=��f��GX�{�/)�3�m�����R��;���w��9��V�GnV)γ����I}B��f�S�0b��튄l-�;`�ŉQ�|�皓�3F�Ǎ�цS�y�U��;\(=D��y���x�tJ�(��,*�V1�\�4�
�w�@7��so�} ��*�yJ�V�gIPCYf�n�����QN��T:��og�r��X�Q�["U	 Ri���܋�P�	��R�����ȧ1N�)��X��0����K����Xl�wU���g{l_'�e�a�W�Ք�;:8(�e�yeQ `"TQ��J!�٣���]�BT���G��r:�:���)��+���3��*7�+Ed�fJ�9�'N�2�T)��n�V�4�YAY]jU��E�o����ݻ�tgfĤ;�ְ��]�Ix'�׳N^�y�ϚO'��6�)��b��^]J��t��0%�:&p�
Ht�8ﰲ��l�'X�5��ͺQ�x銻�g%Kb�жVS���V(%`�P)ݑ�+tύv�B��W���J�`gd���I����;/����v��5.��N��t�"�2ii���2�L؀��V�-��ә��wWG`^�Ӌ�m�^3�tn���;t�"]4U�G^�4K�+3s��F�sSrԎ�����UH6j�N�t�u<�U�q\\{[�ҥ��ۗԲ;�Ν����j�K�}@T�1!A�ѡ���j�<�Y��ݪ=k)�v�F�C��P���l=�$�7q
���(U�rr�kR�,���mɖܽ�b�d����ҌTBQ�u5�
9��O�0pI�9Mn�R#��)����|g��C+m�λ�ϯ*����u
�-�FN�*K��P�]W8ek[Zsn��#+�ƇH)��m�㔻/bY��Y�
m���p�Q�/��嶹�~�-�'��K/�	�t؆����9�K�Q�ہS�Ԩp�N�%X��[���v�j���*Y����t��LV[㺆Mh�j!�1!\�{��v
့�]6����ʽ�o-��9�a�����u90��{�YXGf�n�8�>|�n�ɽ���м�Es�|\�+{�.�VL���c��﷾U<�G��Ǖ�ܤ7i��o��"uK�ٜ��J�H!\�4:�2��'*Ø�D#ec�ͼ�`�R�aR�/����am��f�N5ݣF�&�+�� x��:ݘVÆ>2�]�]p��X�L���EA1�T���d��:�v�c���6]hGY�]�l�Pov���1ش�\Z��X�em�X���䵠��[�]��M{.rۭ��n�%�z��Iu����3r�4�λ��6	b�R���LuaDu�A,���%@�S[ݔ�b܍���+v"6��E}����[ܱ/�w�.V�ׁ���5���bCz�s7����js�B�(���5f�z����ю�1��ty�Ѣf��kZm`,j��G�ٚ�]x�u�]0���X�C�dP�������IW����ٗ]�V�7]�vdܦ�tD ��[��񯪾�����U?mL�HRi8op����x�X���T�4���$.k�g�Z�zޚ����f�N�(%����E�k����u!���hS`���lWN�����7�L�Ux��6���*ni{v9eS҄C�^�q���&W.�Ӝ.���_�,�2:z�������]cP�qn��0y:�2��ѯPC��x�	�J��Q��R��V��l2��>&���!^팎�m,C)Rx�/GK-����N�6�ڹ#�V�����:�8���՘��Ϗ6�w|m��H6E7N�cŮ���Q�-���@Pz3Cw�vQ���c�y����-�v�5;,r��.+�ѵ��dA�����ڨP"1�l�Yݛ����adr�u-j.��Z�l��R^@U�.�e�V�xE�ԍN�j4vq��U�B�<�����j;,�C��>��v��ޮ*�3�;��;��C�0bֹqݡ�NuS]L�w�ҕ�Ҙ�ó���P�ϊ�R��y�p�b7\K������w#;���E�m^&��A�\^������݄���9p�O�j6��>��fN�Γ����X|i>CV!؈���T��k��;r�-�7E�Uv�0�$}�K,]u7�bCU�d������tt)n���g+�S��
���My��s˶�q��
��{��8_:�u�o6�U�e�a��u��8'<���[j���fn�s��ٜ����|z�����$�A{"W"�S�$\����"93̼�"�J+Y"��E*:$�(��D ��9\�&s�q��QjGr)u9E��TU�΅(Т)�M���L�QATG�Q	�����y�	�;���!GJ�(�AFEС̢�29Q��P��az�^�8+�G�*:�p�*�TU�2s�����YAEDX��ЋZ
�"�0&���ܰ���KwptS�p���{+Ԋ��wD=X`�����ۘ�/\Ni�!� ��w=s�Yҹ
I�W.V{���+ծYWQeEHC��9�qd��"�s�DAT�u3��ӮwB�Dd�Y*]�ҫ���b�u����V��^�E$�3R��nw'Q�ȏ1�f[�	Ӝ��Vl��9^��TEA��*�-���̮��R�Q%0��Ȋ�Q�"��Q�t���z��N�]+�BPE���	�n���ڎol)�����qS�ݸ/M����Y��iP���tn�@�P���f�X���nѲ�Ǜ��J�}l%X̿�-f�m.Y�!_��=�� ]�c�y]r;�WN�����{V'e�$�M�c漈�q^�y���� s�̲*� I�7�ϐ�����u�k�WG<�S���:駝ދ�%ߐnw����W�d�ޠ7O(��d���;`��p�R������*U�Y�sȽu��h��Rl�����~��+��?*+�BPU�#pt�u�Ф�X�B����hwd[	&T�5+����i��@O��� �Lh����{�b��m�(�^F
���7E�;O���b�48�9Ǉ�b5��״����<� tBu�o����`����+y��g��~�VT�mh���g�k�pB�[��~���;���'L��1l��;���z���p`���I2��W��� :�x�K��'�t�=#D��N����ۦ�t�}�yؚ�51#��w��~NX�{�x��@ s�T���v�0��3U��qfTL�R1I�c��[��p��R;&4W��1��=Zi,@W�\��|���UA��o���Y��ʑ�q�hua�Q�Uw�(�Ua6�l�<�t\��G{��btp�o�=��V�u�(��X�S,u�6#��ʮĮIĖ˼;:'�ٕe��ʄ9Ctu�sxoF�����>1�1�2i�-a���=s��c���٨+=fc���G; 8�j��U#n7��-;�Cr��B5n}~�B6�D�4v@�q�N5������K1T��&�es���DJ�Z(_�j�z�{�� d�o!��6�z�`^(�n�(F晬����#��2���:Xp������Yq�E.�i�ҁn@c��ʘrںz�rxU�f@q�0*Bx�$k�����9��y��m+��U	�8/+;7aV�ߓ�՟O�M�u�����28�Z�R\4S�����4c;�@�[B1j�Z��n�	�hi�yTp�d��\�����d��ƀҊ�ò�|)�<��Tkl�	��-�	�v⚾��]<��Y�X(eAt:�����n|�ګ���I�(��Dh{U��U~5sGHy2:��V�28c���j c:LW��p�Y,\!N��7U"+�m��ɰE{X����OD�:�r�:��[��U�ߦ�HW�� �u�W�p��R���%�u$CK4�4����NY�/�Ì�{����Ng@�=�@��ߊm}w��N]ޣL�o��!� p+���3{&��쓓�uWa$���B�VL
��=�Ҙ+�{hIx/���O(�q
�ߤf\)�y[�4�
H��Jz��t�`̀��X|�ۥ[�7Sx4��6��lԄ���3j1���R�uigl;���b�k�98��Uͺ���p�Q.��U������-s�\(��tj�t*�1C�N�Y{C����^�Oeڽ��Y�u�����g���U/��v�j��DZ�n/j^���10=�AG�j!א��׷͈Ѯ��Q�FzOQi�����\����Q�1�z������ �ױ�L�����騆�_ƽ�>۩�;���r��'�g��^N~c��t�^�y��{�/Ʋmm��g�D�9�X\j{�2���g�81OaNf~;�#I5�jw��n��V䃁�a�ʨO���zX�x�Wl�<�� ��lÚ�Ej��Ʃ��X鄈ِ"3�D� �J���<�܅\<�{q���c���f�
fL<��k�\�+��=��^�h�����!���W�%���A�6̙����oJ���`ܸ|�f�P(.�����{GǎY�TF�@��qR����
�e
Z� �t�s{����W9��]n����)ˡ�dC� J�J&�&�ʞߎ�u�rm��['S��h�|��T�p�hʈI��U9��Nf�Z���H@|�N��G��`��V��Ԯe�
���q�^{*M ^�j�1v���K�]��\0��f��+����5�]��f��:�YW+��͗�c���z$��ɣz�nM�.ۜk�У��ɛ� ��p�+<o��r���S����,@V�v�ۧ�Ẅ��Ĉ���;�v���p�s {-�YU�1���W;��ꍑ6��� �õ!Z���<�κ����vS�L\B2!
�mP�L���9�\�g;	Bh�P���'�T���͎f���
�i�� ��&i��BmƆY�;s=��cs+��K:ϸT'�qKd���Z'%��e#^�c�ŋ*�p��\u7:u�=���{)uENR�������Z�'<ܝ46�|�ɳ�œ!��9Hd��o���s��6�~�|zfY�8���9NN�`vD9�"|�o���p�bȼ�c4�G3IB'ivFh��*�]o`�4tY1��@w�X��L@>1�W:6Ἶ���F#�F���=�u�\H���a#^E����^Emߕ�F�b��ih�p�r�y�����Yڨb���'�i��5J��A��t����-���Jj�p5�������kE%gvy�-��d�=�;�v~��8_+dVN@-e`一�ׅmC�z}�[b
|�C���,ּ�-ju.����Uv�P'rڎ�Z�3^���G���g'������@.3_PI՗�:^�K����������%���f��"�q��t8-�(�o�{6�/7�%ȗ��ͬ@B$���ܫS	fQx����o��4�����%H���[�U�%z�J�9��.9��<틣�+B�����a�\(n�Y����궥g��t�����;H�{�*L�i�	�(B�*O��蘟$
������9x�+;�=�nK'�����[L'��!��C{\T湀5�e�D���3w&�H����^b�oZ��VWC�
U�ߐ?T���Ń絫����Њ
������	�j�^�����B�!��D�=�\�M[�][F���Bco&+E�}V�7XG1\�Nm:ݦ���[g �(��dW�� Lcx!�yDu��;�+����hު����[2n���&�1�/˒!<�f��Rf��.�c��fD�Y\+��c��o�uQ_������ñ��q��:�,�0a��:5+��j`���SXe{�%z��l��@l.��4ͮ��I�}����J�_צ��؂��p)�p0'���1�K*8Cd��͚~Ol�`���u��f_+��I�(�QQ!9uU�����8j;]:XP��O
�b��s�*�r֣�Q�U`�q�Xu*/H4)�C]�ߟ����]F796]��]���<�B���Q��)�����<`�'�
6��2U���GZ��侚�w��-v��T�����M��Ij��n��N�9*<E�Tq���8_D�@�U�S�y��T)NНUo�"T�%<�b���>�/M�K��7�X�~V�}�p:����N��o�O����*յ��6�nd�!�ehB�B�=E��,gG�����[Ho	��Sb�K��Z�>�iU�{XC�c���+��W�ߛ=�n���h*'�����}3Һ�
�o��TU_E�;�AEi��dN�Ҽ������ң^�pbQ��W�'��<�WxT]�����6���XW<-�+w\fd%ʼ��h��C!�m��j�߸P�#6J��v+U�˾�̮hn��U�j	���΅�DLB�Z(_�&��;q�r0�7n�W!pj��H'�%w�����Wa�z�ӎ�I�޳N����c�����h��S��� Ay���*��Õѐ�sJ��@`c+fC�^.�P<+��w�0;��Ļ���%�늞S+w����c����R͚XG]�}���:�j!r\����m	
�ƂLgxH`H����:�W�S�ssGQq}��P�T1e�"�rw��d1 q�3O�#-�#/��=�`��I�C��.�n��oXɘ%�QĚ�H�ى��-PW}����U%oY�p;猶k�U�^��ڭ�F��=RӾA-m�W�revv�p[�eu-��5����m��Z���L��\#�t;�e�<���ֺ�v!o����f��z/�D^&QB��u�ngĢ��%��8��W˅0>'���^̶6�
��J�����ύ��x\�5Q=��$Ɔ7P!�оE��4ñq�����^�ʌ
���^΂*;���,t!L6�Do<�8W$.|bF���jG�3��/q��!\�W���\^T �%��d��n`��s�EbNMVRIv��7�bC��^l�:�=+�/M�J�W���>���7��{����ࢻW��3�+m�o��F����(?��b6i��xʤ��,{R|��p�<�^�O�cˈ{x)yiRx�G|e�y8|�P.{>w+ӶS�yX�툋�)r�C�ty�N�m@sz��&u0L����l�㪽��.v����\v��M�_�e6"�w�XpOf[/�(��z�����G(ܲ�=�ۮ"z�������j�;��6+�eC}e��g������{�;�^1���rj�@���w �9ndS��,������,`w37&��h���6��[{��_����B�Ȃb5�L �J���<�܈��0���Ȁ�B�eں	��Ό:��aCW7ƥ�M�`�/�N����r-xh�e����4���`Y��P��^J�HH��x{ǀ�oe��p��y�=���� 6p��vF̗����Vf��>�͡���[h�K�Dk�1�|o�y%�&w���y��n4�-;���GH Q�v@C�/K�O�G�����]pQ����	�R͎�^}βcߐy 뻮�ꞥaΛ�4F�s˾Txs��TT�0N��Ы�]p�{�H\`�:�i#~���U�ҙ�.cDp�7#
�yd"T�NɍS�c+�w�"��Obfg1���+uh���!�K���9�s��f���n�JY(���M�i^c��;�{��VI��>���ݨ�~sC�sL��59b×"��9��ݝX��٠�\���"n�u�V��[��[�HC��L`��R	Mc�7c3\���{-�H��bp�.�"�{� ����0��)��O<�b�Ѕ�w��c6��\���;Ӊ�n��@�3C�uT��D���n����p�}��p��Y"����V�n��/�����<��R��)�;��]0�<Je��g_����,��Q�Q9Ha��"[�ڼp�qlM��6&˅�C��F�c�5�1�h�8�w��\U��'LW2���T3]�����v�J��A�۾� hp�ϻ�FgL����b�$E�������FWa��꺔��,rj�=�כw�ak�+��K��e�����n����7\�.Q���qd�)+:�\�l}f���2����:����X��'gD���՟ /�ݾ�6�:i���$P�=��m�mT��YN7���F�F�tJ�q&,F�L�f�QB��_Emߕ�
�e��k�kunT:��V��Ňa�����`���۪�KK�|;�O�4�π�Q��zV7]�)w�|�>WF��R��{�	1��T��XЧ��F�[
@���5��B��#,�(>0�LY[���r$��ܙ���p�c�L'M�cp�c�)�?Oi:�+B���Oс~�]��r�:.�2��]_�+�Q��+<4m$�#�O3��C�s����Gt��T"V��T�����[Y���pNiXr
�b�m0����9�G��{\T�]�d؈��"H��`�]�s[���8`�'H��:�L�cq��v�ceM>(w���-{�u�3o�������=�b@vU</���fn��ݺ��=���s�Y��G�)ӂp�I6�7w7�VE�'$@���^��:������2#��3�lU�=�8r�i�>�]3{r��D۱�����Xޫ�vp9��b��C'���vl#pq��g�W<��{DU���"��&�9Ҹ��lgap<i��F��ۇ���CN2�,Q0ɚ�nRa�.{�}��f1�F��V��WgD����<�/dʇ��p�5 4mӻ����<Q=��o�:�y^K���C�ͨɘ7�x��<��e���3P�Xv�fzᩂ��3�����Q�q`�B���1c1���9��L��c0�E�
���]�Ѐ���1���p�j�p�<�P�!���}{A�������q{<Ԭ��.$�Q9P�Y�(Fg<{U����MI�[L@�y�ѳ��f��R�(�iۧ��\�C��X��HV_(�������;�(�u:>�btɖy�Vf��ݸ����S�f�F� 3#G>��[XUq�p@�ٝh<5�_����n���;�8G+'[Ǯ�M��SF����'�[�a�����s�4\>�\;6@�0Jߪ�z�8M���0yb�|7�y�*�D`w��nh>�XXo��e#�&4T#\c/ڪ=��bv@�b�C���<TY���ù���'/���A�YU!�X��"���u�㌽5
�߮�`�K��ǖէ�_v&�=���M>@^�oYQ5�Ip�gk"���'��>�Q�6< ���ZHEn?S�j(KŚ>��:��i�Q,��5�J��Sq���C�k��gw\�O���SR�A��i!��ZT:���U��2�=�SQop�jL�e�H0��ҳ	�U�@�̔�P�r�����	9V�e��7+;+�&�LR�\��P�k���u_0��5�g�����o�F�������]k���b��N+f�b�E�q5e��aq�J��Y��o�Q��[�� X�2�c�.��m˙(7rF�۽�˾�.�PړsV]���' -�L.ǔ�;f�c@wXv�m�@^�5t%n6;*.�,�j�6�*R��k�n���تˣQjt�����=h)��ބ�b�&��mL5������-�(�Q})={؛��V,����N�t�}�}��f�������)�\n��-�xUF���J�X���J�.Ύ�ڎut�r���T���f�s���k,"����u��w�o�#��;w/\n���3rF%�L�P����ƹ<���f��5�;HI�:`��k�B�OZ�KF��;Ps۰����	�M���K�)�׃��������&��%-Dp����:�z�ҭ&[ɩ���"�䱊�f��-�iB�7�wE�x����Ebߵ����On���V�^�5�+TF��n�39T6q�]˹^Ҹ7Fa�49�Eب�L��|��x���V�b;�^Ro\[�#���W��U|�u�u;QPu�o�^R㒮�n�*��n�l�j����J��O$2�-ts���u;鲂�柒`�7η8���]nތo[��;�0�v�e�I���v���q���c��B�
,S�۠=ż�����r�;������z����Ӻ��$��\��{��h0w6�"��ͤ���]�樷�쬛�K\��|��'s\78nWZ�I [ǥ�K�f�N��I;���di�2�\w����wfoD%71Z9fӓ���ǯ��GQ�f�\HP�7I�#toLO4�ޘ0���A�)�*n���u��j�V-�1h n����a��֗�**r�P[+�X&�-wkY�#J2��E�O�u6�A�FH�mrW`�ԝ�j��z��,�6���$}%��
$���y}D;n���Ϡ_X��ښ�lAqf���A;۰��,.V�������ޕ�=�ݴU0wx��v٧��ҸjAZ�YK�� �݆m�ˋ�L���l���֩�����5��ұ$v�1w����`�"��y,��]��E5��I$��ٳF��ۻF��!��X���,L���6����]�\�4�(���ޚ���R�m�/��7`%�H���Ɔ��n�މ�q�	ƱGS<v��$7��>q�[4��x�=Y�����dnK���鶵B�{;@�F��R�4��-�M!	�8�n��Vݜ�r�ό�T�̺�U���ͼ7A����J��w��Q���nG@��}���@@;�C޻�¸������C#������ҟ�g��h��t�h��,������=�Щ�z�����DUQTfy;��Ћ���-wR���r;)0��%9#�N�F�e�j�����r�L4��t=jmZ���g���H�$��E�y��8��.�'Vs�4��Ü�u�܍�9AAs̸E�e]�������\Bu
s"�us��V�+�)�]U�U늻����S(,�]�����.8I	��T�H���TK���p��V�r�4]�w!�y� ��(�GsLs*�Q�E"�'@�we�s�r*]�\5�UUs��<�t2�Ow�9�A �v���8��D*�^l�wJ�G#�8y���\ʢ�/X�D�HE{�8�!#X���q�3�ːf^IQU*�AN�]YBy$AQ]�
֕ȦEQ�T�Q���::��NH\��S�U73�̨��Y����f����z�T��EDr�Fu�����M�T:��QJ�z�Hi;��Dd�D��Ki�&u]���w��[(l�Л�_v� ���)�XR�ʊ�ż�����{�Xor��֞<���v;qs�z��?
�1a��Z��@wue�-�=d6d�SOK���S�8��G�7�w�¨�"o��s�����ÂC�}O^c˾8�_=�)�hr��q�*I�~��<���}�ޕ�HO�e�a�na��; v�;�z*�!�t
��̝�چ<5��X`��<���a�`N��y�����xv����ן)���c�}t��$���S�s��x|�'y�}C�<���iɽ�;�G�Dp�؇3b= �x�{V���]S�>ū�,��P1y�[�<Hd���_����߻�yM����M������	Ӵ����^ 򛐜y�|v<?|[|Os�܁�'㴏�v]�7�/��n��%p.;�����Ϸh��ߞ�����r�j�Vj�SxS;k`�x��w���ߺ)�\~O��ߐ��<}�����=>s�����<�N��������!��C��]&���x��a~��|�X�zv��$]��Ǽ�5k���t�}u�|��_X#�*�Ǖ������P��8��?��ݷ�?&��=n����]��߱��n|��a�Q�&��GT{�ż`
� ��q��'˝�܇'�=������������Mցز���uG�@��#�~�P�_h'�ݼ����>����i�Oܟ�����k��,ro�O�o������!�5������>��~��xM��S}��߀�7�E����FZ�Z���r��=#�"G���!'���9G����}w!�����)�S~O>�{Ohra~���< ����!�����s�^,����q}�~���@�~BO[���\yϼ�P��s�W��Խ�������<;ux3 ���s����a�`����\���}C�A���N9C�&���?��]�7��^�~��®�=�'���I�A����?�z/� ���x�6��/#8R6�e7n޽�ha�lo`�Ae���7�#�֓�I���ۏ�?�r�����Ǎ�w�iǟ��<';{y]�������s�x��<!�4�On<G�������57��+�P�C��Y�O*ٛ&��;�����<��C�������99����N��'�����U�|߾����_(z?x����4��|�'�94�On�������O'��v� �����mj�tP4�=5@��atK�V�9=}�WY���Hm�U��ζ�29��n��6���Ѷ@w#o)�xq!�1[�|>��U�
�=�69ۧZv�R}\6���{�Os��+���9���gZ�K^�]O�n#��q P�3:�@�u��F��e���xvo ��a ��a}<��~v��˥w��ߐ�S{�zaM������<��&Ø{X;a� ��`5��y+��
a���Vk�O�s�Υ�q ���7"w������GT�̹G�0�x�0�A��Cˏi�������o�=o��m��z��Í�<��>�|M���������ާ��7�7�\�o{���umcNKUW���V�j�󷹀vˏ�����,
2�v����<����;N���o��n8�9={��>������HzL/����|����ɹ�^Ϝs��w�i�+ŀ������������st��Ol=Lnoy{ڪ�_�X	a��}v�>Ǆ��������ܛ�AɄM��NW}v��''����|q��|=��|w�;�o�����L.>8�������fM	�u�-�ԇXa����rZ�}����s�J��ӏ��;)����8�N)�� Xa�)T�	a����;��>"�������$��o������>���O8�;��!=h���Yf��?_�5`o�4���7����C-��Xx3+f=�ސ��P�o����Ă����{��<&���}~��뷤��'��<$�&��(������x},���,FD��=�#�3
w��
���Q펷�R�|>����30�0ϽM�iAdxP����~����<�yB���o������?�M�	=�p��r_G���c�$������q�𛐿�p�vx����xDr�*&B���B�t��<��}O.<z��r�?�����w�i��x�}C�}v�y������Mm�#��aM��{Xz����<���<G�CzG����{Z]��X�j��F:�k�3V3�U�=������=�!��㓓�����r;׋�S�����>F�90��ߐ��ʻ�i�C��������~���X����~���1&������y�8��:~a�o�M�=�W1���`�qwV�������a�o/�f,a�̜}I9���{��P�Nq�=x�'���|w�~x?��L)�Տ����xC�{�c��$����= ~I=��P)�{��ɀ-�!���`<��}G�c{g��gd����u�7���!�{_��T��w�k/�iK�Kh�Ś�\Tӱ
W}���Y:Q���f�+�ܥm�Zb��ѻsly(_*x�Z.bt��!�{y��k-k��v_:]κ�5�J�'v.{��0��]E������������� ��-�[��o�����=&�?$�;�m�N�>G�<u��r��&���m�=^N	�?<��p'�yL.��=��|���v��nWo�&�G�~}���|mdKC��]�M	�C��[`�\[[x��'�����~���O~>q&w�k����&���G�Ğ��M�'��]�3�8��7�$������3s Z���&�� �×us.�aڭ��ï���
lozx�o �x����}����	����xW!�z�Ǘ�;�ɽ�v��}C���'{߿x1����9<�޼�
����~1�9hrĿX�9P���`?$����+WQu�\�:��U�z�/Y׽L=`|OǸ<y����}^���{ps�|���ޒ@ɡ������M�֬uY�o�J���ɼ����'���<!���?|���yL.�����nC��LRsZ��/jʽ؛����x�����ŷz� ������$ޓǨ�_nܛ���xW��u��8�O��?�ߟ��=&�>>�����"��|����������g�\o	��8}�-M؍�9)nZ�ܽv��jo Xl~�>�x����raO^�i��o�`��Wo)&�}������w�����>��;߾<������C��yC�aW}B���ora}{��������}v�!�]|e�b�y����v�
�f���[ӽ��ϜS~BO�޼|�*�SzB|��{�_��������<;s�}v�F��O���aW'�?�����!�(|O�s����z�zL.���w�>8,��M3�SL��Bb:�!�0�¨�����&�����\r�XT�X �x�t�oz�{��Y�ǿ'�p)��}�����|@�xC�4������s��Hx�]�S~`3F�`��:�jnY8�襹��X{�Soo�"���`�)S�7��&~E?;���P���ǁTߝ!���w����Ă����y@��o[��xN~;ro��(�Nҿ'�'��EA�9,k�GÔ��[]� �����	�	�߷G���;H�M����X�����r�w��:����?>�}O�ɇ����S}|���Oa�����q��������v��T�W�RU�Z�c~�W갼֠�gNt��׋>�8�:���IjJzm>P�U���vFo3_@!6U�Z�Ѱm7�8��NI�f�r�ͬ�)zY=��\)1���h��,�'ϪL}[˸��5�j�_;'zZU!+��/���rK��`�(��'W�����||���~<YC�aW|O(w���]�O���i����S�.ߙޚ�=,<�Û�-Q�fo �=-�P���~N~�$�~�ɼ?��xq���cˡ�1�}؃�QX(z�Y�����Kj����I�]�{�}gxw�i��m�'�9�S��&|w��=G���!Ʌ�A��O�zC��|��x~���+�����< $��������]�7���/�a�[�3")��nk�qg7^�ӹ�k ��ox��C1�L0�oN>>�����]��y(?:W|v�	ě�'8����xg��?�����'�������ސ��P�J��=������_�$�������s)���#�k_b���`[�G�L{;rf���'���>�}BI~~����yC�H{>��<<�"������m�<�xW���zOh�9���D����;{�!XahS4���'�e����=�=�D{��OЕF<+��N�~��C�a}�������ܞ�r���.ӧ~~����>�c��
���߃wF�97���Nv�{q�RE��'���&����~�����;搜��Y�:�����������<��#X��9������4�s����c���{}��aWoA����|��.���K`�c�G�0��.�����=��w��Bq'�=�#�;�50H���K�5���c�*��}�x@����/���ɾ��=^���N<���}C˿;]�����!�5[x>��O��aw�k���;ʦ�������nOi�<����c������l�$);�~�=�g�!_X�+�|��	����s�x��M����x���0�\I�����n@���{BO�nC��}CÉį�>�|�o�N$<�o��ߓ��O��{O�� x����3o�^^��2���(D"����+�`��q^�Uz��^L*�[d� ��]nυj�Z��df�:�������%��Z;�	�j���w�mQ8 @u������n���h�~7Ykty�zts=+��kt�G��e�³��1�=�:׊3[��-Q4��	�>��!;�t,��RC�vfWcf`���߀��1M<�B�3�{gIͬ�:fl|��Y�oS�T=8)jƬU�+�Z:�s3('W7qHd=�^�CՁ�kݞ��|�0��{��(h�}�x�l� 8Ȫ@A�̗QHGۗm�Yv�7*)�Έ�Kf7�Xx��L�vLh�k�eƪ��^H���[�-&�����=�@��3�Q�Rw'�Q*�;�������r\q����;�X�P��-�t��X�	���Pv@�qN�q9�̮ޮ*�h��U��q=�M��/��1�o{�Ը �J����n�?�C�7�ӣ�}fɭ��%}r� uN� 'g{7^�ܳ�}Y��*��F	Aq��..�¼�Wq_=L2��9��9p���m�K�ؽ�Piq��s	��.���w���t@�)G���"��A�f��쥦�N�*^���pF����-㠍�o��͢����:��$י���L���iT���Pe�b2(,�Yݣ9(�fIB��ն�l#,m��bcyK51�g͒�@q�$�|�pt�5v�@ƱD�+����u�j���t/�����%��r�y�R=�//��h8Ժ���ծx��W��]$e��ĕ.Y��A׌��?z.>Z�uxV��ïNS��[}������:���"��2>%�[;��H-�RԾ�ml�fn�墛����z����+Q�+KE@�#�I�St�/-�2s�t�*��'Nww^�r�o���2�?x-��9םz�0�ɘxv#\�3WP����&ĄD���i❾�=V�=F���ʐ7��{��k�΁���rzo�k��u���I�[N\����~��N� ��M�s�C��pp�3zdTBRd٫'��J�����`��-
��UX��͜���7�{����N�7�tc;�S�����H`��{Q�bR�`����r8YJ�v�N<�G��sZV�`���e���S=�xX�-گ=�:J9�Vw�$\�t*�}X�'Z�����`����p�u��y��]ҍ�{�����pJ���.)y�q��V^*Q�CV¦�Q�d!�骤��NAw�]�ySE�����Q���3ˬ�e���Z�+��z����8X0r���4蚬�\ 4���,�5X��~�����>�3yHu"�'�[�c<wi���0O�������!K�L@H�*G\O6��U9}s��x8CRé�\h_t��K��܁[�U�����䨍��R�ù+��C�sԵ��8�z����g�Z�Dp�������j�ktt`��N��*��I"���e	D�j�fQ�s|�7)�>�!U�Ђ�^����h�Kn�l���t�f���K�=ϛ���������ݙ`�Ć���\	k;d�42Tm���Ib/kc6�G�\�b�0��26[/��p�Y�Q���+!�0�T�Olù����1jO���T���>%S�^&�>�WƲ�I���[��'s7�#�����$ʎ�ǅ�h08}�A��;�ߎx
�]Q"�U1ݾJm���%'V��o0SNy���{��dgIXL���'A������]s�}L䛲�:�0sNh��23ZÈa���G5@>F� X�5��(n\���n�,�zw�;;�O	��L��q�c�� ?{^�1��K(ߧG�n���YG·�(v��B�L�:�|M���Ʀr��oq�U��3e��sڦ"b�;`'8��=�m����-��R��s]�	���^'�(HN]h�ɡ�X�7��s��,v��#�ub<���TR���ԕ������1��^�Yh��T��*��C��1_�<�٪��**|b�,m�Ԩ�Ѫs -׫G7/7�~K/�5�Q��%#~�4�L�u*�q9����:�k|�MnCV��%��Z&���f�辶g'�g�fw�$Uû۸�o0R<��sk���.Y�v��+vՒt�o�wr���p?f��t������>1�S{+�Q��ɊG�R�/v�U�h����CT�&��(;p��������v5���=�~��Cq��9T��z�\;#dOI%&}��9֎;Q+b���W��Y����$��Yxn1�3z?��������@-`g��z�{�uf戋��+
�V�z�������'�=:l�i��B:!���{c��.�]턅���n:6&���Z�`�)]
;< W���\-�:�*C�_�;H�8�l���]0׌�곀Յm>��:�~�P\!�ϻ>ٻwsì�S]���W�9�G�y<T�wx�X�l��#����˷=��uY��p
��sۤLe��)�FPw=9]�,S�{�G}���ո�LU�4�o�����
_�v$1�ו��5�2ez�z�!]^x�$#c�0���#f8C���ᾫg �@GC� 5��!��"�5��+����۴(�P�j��o���2[ͦˣ��`��a�rxp絪��&�}Q�I�e��L�t��6��05f跺��7��:�|��#4p=&M{�Pi�߷�Lx>��;��<��d6b�.
;k�243���Q"��ǅ�M���a���[\.��k���W��cyW/Ǩ�K7�J���s	��h !�Z�����7!o�7{���h����.��-��1���@`��>�³Ui���鲺���c]��c���z,�7����������`��zf<|��L����bǟ�Xb��?��� +ڭ�1�&��j�OB!�a��]���˃�}�2.�
q[�E��>��`�Q9P���'v��S�P��]�W{77��<%(��	:�K�V�ϐ}��[af�Y�%���\�y��:�����Q�����lB^9�{�h���_7�O���d�g%։~�\O�g@}7ʐ�ק���o�q����˩�������$���>�any׷Ms�4\C�ǳ�"L ��:�1=�)D�n�]����*9�m!\i��D�V@(</��{��1q��j�{�9)�Y�C,ؿF���=�� J F�L�&�S���ޅ�R�N��KGC!��zr�B�QW��R�ׯB���َ��U��'��C��<��䰈�[�.j���႐��R���J[S1Sǆ"F8t����} 癗�kvh��� *_��f�v27��js�<K#�h�����"��!ʙ�1� ���$g��A��~�R��`��֪ۻ�Sthn��{Rо��,k;2�������]����S�]%-D�z�c��L�~���^��PE��o�)���7C�:�.�o���W ���s�K��[������sn���]Iֲk��v\jPw���˺��mVP�:
���舫�Wv)	�}�v�O�.I\_虄�A�<n��
sѐ��j2�ᢟƏ�)s+�_l��љ�C�9�9��e��v��&+��1~.q'"VPp�Y&����e�ճx�Z\�Ob�;�*.J5<"����vv��w����^K��L1秢R��
/s[���w�۳�ėQ/ɍ�j�u�Fs,m�CA���Ud��10���ݡ���O����˯|�ߺ�pX�Oב������Ӊ
�+�%�v4� I�&m��ۻ���j:�h̙��-JuC��D�Z+���[2���v� izo�l��t�J�N�����r��iR��Ĳ���0���f�ȥ�ɳ@p~;T�p�A��&W\��B���u��v���"��\��钼,N9���>�Ǻk�=n�:؈�"����F���w\�o(S �(c��a�ɝs\�{��r5;`��^��M�t��Y�3N��(�T;�,C�x�r�TU��}䭬Ե�V}��^�o�>��9�N,�2m7�4�{�M�7"5�r�*шf�|F�-۷[r-�]}�X�m�ksj�rk�+u�[43iU��$Ҥ����q�L���7Z���ԕ�kr�c�}��u��p_C�d�#[ܧ2�����*Rܭ븴�vb07��]�Z���c�Hx��'��n�v���5����d�M�8��k#{�p� vi���luM�Ҭ��'��ů�"��]���}�RZIH�[���:MYbL��nT���-o5�	�%
�Yo�5I/叩a�'v�Bx%���]�N�n�m1J�u���u���o8�� ��Yκ�i2�ț�vq��c�P�7�wK��մ�@^f
�k�%�S�\�|u�N��H�7]iW\����^��4�'أ4��#%�F�Q�,���eķee>q�y��J��;�9mKo��k���<�a�P�w8�E����f}�8���+.'n,g,_]���¹�/n�/�����L�������E�ťb�6�	.�,�G�&�ŏ��k�{� �j��N�DGx���̻FC����w����yq�H�Ð.�}Z��xJ��*08iW�Gz�9�����j�$��ǫcy��]�͎�+�y�$���H�O�Qcn%Z�����pê���K�s�v��hSE��]�����jN��V̨��2^�d֐��i4=J�/�g�z����ˣqZ�;>��<�\�YY��9g�%qm:c�8U�6i����)��g6^�}�ᢸ*�gf0��W���{Ya$[�؍�Kt��d9�%f�e�6�����ޑ}�祆������u�͡KNl�P�1]��u/��vYњr�,�F�������m���R��N���������r�QD�F�^:\#J=�ʭ�`<�"��Dݣ%$ő�9���ЂТ	'�U�����h֧]��+3^K�N��΍)J����*�T[x
mmDs��(��TV���M���*n�)�<�����e3/"ݛ
eH^�J�Vn��f	n�BN��鐂��m�r�N��AY[܂'F(�.�ۜݎQ3Z�AP��d��-E�)�^;�`�8� P��J9b��Qu+Q�^e0��.�TX�Aj��J�Y�a�|')�M�ɮT2e.�M�V��GVJ��@������֪"��9��W+{&b�������Z�ݒ��.�cH;Q�*�D�`Eԯkr�\��9�/Cx�
PV��ك��r�3I˾N���2��o&Q��;�W1�P ��yZ�5�ږWc/&d<#��9���o��n��f���4��ٴ��mk�Y�I�
�Ъf������d�H�%!�&ʻ|��uѡ����N�\�y���q�\�v����m�NF�ޤ����O76��	4��9ԣ�4_gCD_V_4A�M�`�&��t����M�[��ȓx6� b�+[p;N�Nv.��ڰ�۰8�	>w��)�;{J��8���RF� ��*�&��w�t�f���Ђ �J��z;�t��@��Y�����e�=wN:�����

��UK��㛺�-�I��Bه�\�+�4ȥRH�B�"��WD������D{�r��̥���\<��]3+"�]k�s�Ё�rE*��JqrE:l�"�E����*�@�Q�P�p���<�r����^�zx��r��B�U�G�*E�FQ7Dn&&A:�^g#�SP֗�"���N�YUuH�U\�����GM�E��s��=S�U�p��t����p�P�Ī	A�u�(�"wp*�Ȫ�G5�p�I"��"��w\�WC�=k=��D�Ѝ�I��NE�Y���n�K��r<�u��e!F�	�w'<T�Ip�wv�!	�
�Pi ��/�TE mٮ�`�՜淸�51j�ĮcJ�!��11�N��\e
Mڹ���/C�-������������^��#�j����Ĺ����xU漤g�>?R�R�ʊ��N�d�a��,���z�.�Ou�ʭ�Ö�V�a�wRF3̱��90h�`�Y>�9�*��J� iw=&{2����e ��*�]IQ/EY����V��<�������E7uM̎;@n��xp���$�Z�����m��{�p��}�Q���Tr�i������p��E9�#�y�l��7;�1��Ӿ������(�z�~�ͽn��L�1�8[r0��<��N�N]��w��8sZ�r�8K�mD��u��"iL1����9)�z����1p�p:��Z��Nk��N�粳2,[�\YU����.'Ĵ{OE��&2�TH�R���F$E��H1S'�,�J��Y��T��0���]�Ҕu�k,��<�v�W�G��}G�io�;��mа�`�2�W�����s��� -�� !��ls7����qٕ	��\�;'�5�
.���E���a��g����[wp�\�;�~�a�Ixu�����1�m��p�"eo<�U��
�.����mQ����i�Z��-J"���
T{ntWh��x���WB+���ѽ��E;E����YCL��.�y�$[��Z���XY����C��S��{�v_G]������Z�wh�E��:ػ���S�#�����9Cyu��=�6���ޫ��k/i�zM�LD�S�wX��/ٻ^�k(�}Sn�aq^������J�$Ċ��{�oʶ���\�U��o��/��uECɴt�븽�T�&�\͆�SԵH���w	��@�5X���-}��ZU�� 3��}���@h���e���\g���`�S��q}�G��o3Ɵ�B�1������>��]�-1�3�U�Ɲ}����&��V�絺�5Ա�
����ò6D�פ���Mz'\�m�cA�;�d��ÕuP��-��ƹxo�1��Е_F6���� ��V�L��^����:Ţ�����J1�>���֦(5	}�t����;M�9B*Ӷ0ܔ{��|�g����y�ZR��p "l�HpzP�e�w��Q
xh�����+S̽>��ɹ�jR��u�U��V�.���|Q��zR��&��N��<��v&���4�5���Ƨkwz��,��L��n�3ҭ�T��:���T�|���:�L�cr�}��UӞ��7D�
.���A�0N��L�4�Y�KB��b�w�4c��%�,�&��θt~����������W:�sl�B�q̺�]L�Z�ި{�з�2r#+�-Δ�ɅfҘ���B����^Vb�G_t�C���<���w?�3w:��-�S����Ub,k�@�u�*�����p��V�$�g��O���OV+�w���/3����|����L`��ئ-��gtu�,���Y�NH�&ޣ>C{�Y����.�|r���"�^�'�w:a� *�sa�v�;M�;����Xt�
ܙ��/3���4��"�5��y8��f�)?����zG����{[Xd7�p����i%�USm�k��{�d0�����H�M3k�����+U{1S���o!������e)&�T0ڴ��m��G��8�t�����90�YzP�'v��S�QO�Mޝ��\���WI�(@�C�ܟ!���7d��ڗ�w�خs�!�R[g�w&�핾���K
��~N#Ι,E3���TCW\4d>�^�'��L��f�x7��7�YLtG���Oϟ�L*�&G3aI��.��0���.,!c^�=��F;�+��9]/s����Q�H4�T����q��1P�a3q)Շ����S:;��\kLgz��!J�%�7��Z�u�p�wm�{tpT�����r���[����ѧ�	F�7bf���p�6�����s8#����O��SwY�Č�d$F4<�#��3G?]Ԩ��|7R������d�>6��k���e�seΔvv�x
���Dz&��N;���XZ�s��9�F+6�C�����ȆwN�D� �Mi���Q�}[����`�~���ǐ��2Ʉ8���N��"��Cr�p
Y�[��*0��\�y�3|�WmӸ@R9����p����Z'��TK�/�St\��/��>�i&^vTq�!
��G!�@��l��OL��
��b!#�3m!�_J4�]]eJ��%�G��6��y�Ҩ�3��yZd7z ��tB%OI�L��*����״X���p!C�.��N�<���,)1>�ҸcγRoˤ�7�I&�w�:�l0�vZe+�$�3��#"/��Pc��}ګY�e����ʈJ����n|����B)&,VNU��y9���D�=g}&433�2��\��kN���y:�P���9sW�4���[���*a�=wB���� �`�����NϞ��W����砻����
�v��Co��"�p1qΪWI�9�6[��!��`!��΁�{\�^������n�2I���=Q��ϢM��wk͙�����|	���\4عeOv�w�a:���yA����*`��u��%�T!�i�n>0__�]��ᔞ�����ǃT��m��;�xi�4��{\z��a-S���t�̡��ވ�G�����<�N�!Vs���;ր%�MBs�j��>��B�����0�X{;,*�-J�V.�v�P�#�-�D���yT�Om�4���Vx6��pj����ѓ/*k�vvF�0�W.����7F��R�`�H���ҭ,��HE�u�J]�YL��qΙػ�����y8�G�k��NZ 7F�A���� �������G_�]1�g�>��3�ڊ���df-����AC&E��Y��1�D>=5T�����ɼ0���+��:�Dp@)�{�S��٘lz����_	\a�e�*U��RMx��u0�R�%��\�q8�+e���T����9�>���ۇ�	�!x�X��v�n��5%�;���E��_�ۮAC�ݒ|�v��{�����>�R��7 G#���r��S0Gu�]g������'���R�/R�ᮢ�^��7{�i�\�B��2��a�TUI�}�v�4�u��T�Q,�F�s�J��=%>U�b}�ϰ�
�3�ӆ��o��4uq�9^����u��Oq9Sp���x�ov��p@tZ��X����{2mo^{��e�`�f�,��p���(cW_%�/Ƀ���o9�����WKB����љ�j�ι��P��������5|��G+έ����
7����\!�_UU}@�%��cZvxN���ɈT����x��A��;�#�Vt�˕o�GU�}o�YA����OO<��M�
ؑ8�Utn�ܑx9�=<��$�/bn�u�n��"/���u���ٸ��lz{z�����o��n�1hȄR�S�a�&� ��#���.|T����+�	5��NE�?V6z�.�j��ӛ�6ε%���T;(���-��=�
"�Oi/c�����T��j�4�����L橈��N�	֢���騁�����Q2�8���Ԋ�R5.�já�E������u���A�\<2��q�k�s��]u^�t~�`j��	N��6j���O� ]�H�l�WYώjf�ez���ƺy����{�g��� 8�t��;�p�_��d<jU�]�R5cJ���g��_H���p��N�ϟ��%;y�S�^~��<��#�z����G�W�y��t�����vU���4���j�2S���Ì�1��1�����F�̮@-S�����{=��wI�ZVdU:��3w���&
;�W�G}b����� Z]O�ɼ��ު佝��o��{���ׄ���&��YQ�OyI�Ǹe�AQ��4�6�h����;��VVm���C/i��{�H��KPt�BT'�z=��F�p\�d㉐%Oޣ�kf��̤bA�ڄ�N[#L1�y�!�t��m
;�RT�	+7'�H��dy�x�BE��[$uB�&�v���p�3����V����Z��~����~���,�T��Mk.���b�^uX�;ׯ䉢�c9�z��c�=5�5���xv{�:5�Ј0�'@�R=s�Q1�t<0�J>��v�ݷa����FY�KuÂ����n�x� ��#�I+O_�d��0eT2�2]Oe�n�#g��UE��p��}7"�	��P�ճ�S�#�
G 
�e�P��|a��*&2W3�=[�{FsP��?{2�uj�MwJ���s*<��Z��6ڠ9���JQ�D:�ƛ����e83�4U<5�Ky���F�):�\=+����`#�����ͳ�#�e;[�UZ��u�xPϑ�4ͮ�j������~Ń��~��{9"��oh,���V�w�UCݓ���
�5�t��p���m[�a��e�s�]�Y�j�;��-5�2��8^� JR�}��x�F��gr��ljǽ��ź>���>�r�<6�r!o<��Mz&�A�4
o��9ˬ�u��r$i�te@��T�sת֣N�OA�؝^��q�V���������$E�@tѽ������3��BS��`�Of�[sl��������y��S����X����{h@�s�+�z�!�e�bm��e#�}�|��6+��Ć�n��a�u(��6c �k���s�M���G;�殸h}�}T��C�^ݯ(������o�zw~���.��3�%Q�I�ҟL0��w��{�x�����f�w�ާz�p���*�	��p�jىe�9��aa��2��y1�'7X��V��9��-�΃8�o!�e��K� �k7�o'��fCiד��h��)m�O#۳����h�'����V��sF�*N��7��N�x�C��<��]dEk�|/�k�:�t�7U��d�~>���j����lwI	dUu�<됬��$<#X��Gp�/'`�b�+mG��\p���qog����:S"�J5`��b*�t�+ ��m<���K���5�+���qV��3~s���(�H�vzL{N8��Y��L�u5�wv� !�G���p�F�L�n��k}P�f�r{Ҳ��EmJ��ӼT�9�ֺs�䛣sx7���;�d�ܵn6ȭ6�����x�v-�һ�I�K�x�测���3��Sx��S=ݽY�H�g 2&R	tahl=��<Z�1`��]�\i�R�WLDc��k�r�����}�ͣ}:[�!� d�+&��H[���}����E�0�ڕ���rmuWm����es}%)�N؇��@{%W��b5��7]��X��^����\<��g%U�s���]�5'C�!LW��������!�g��1Ӓ�?��5��{ؼ�y"o��O����ܬ�Th�D�)<�AQ���W>�rt���@�c��4{�y�u�2as3s����1���Z=9�lQ�4�&�9�ĵ0l�7�BD�'!�}1y�R�Qt�_T��:���X�\����U=�و�ms�6�Jv�b)��� �����l�d�t�$7��a��y�B�x� ����suR5ϯa'l���<U�u;[]"np�Eƺ-��n��y@r7�*��8;��y^5���
�k����7xՅ]���t��7\SGt���OuF[{e�\d�1�N���f�b�r�} 65A}������ev�W��������+�\CrƩ���F6��RF�0�Q��ܷ�S]}zdRd{�������nu��X�D WHc�*��`u#O-7;g�Y0̼j��K9��K��F��{��U�I�3��'{��ur
�ʋ�������w�.���!f��=Bs���˻��i(9@��J�|��.������������ϛ2r��!W!Q���N���|w5�#���b�IG�Ҩ��ڧ��ZV��(�Q�!��(+��]pQ��>E�q�n@�G�T����¤M�I��O�-�1� Zٹ��W�bD�/�\C�����,ks�v�7\ƈ�58Z�ɉ�-���Y��S��F�q��C%�D���sˮ&��,qr��F4e%��n2�@���Ħ����7u�r*�6�,�v���B�OQ%qWu�d��.��ڥ��0we�o;9��{�J5�3{�v-���
�\�Ҥ57&88f �Uo����>�:�o0�J����Խ\GZ@��۪.#�}lh�V)��dBڠb��a8 	�rx���=C�^��?���=�ok�e��ޘ����3p�e���K(�=���l-���t�v�vj�}�:���b[�w�TK���)�-��Ʋ�{��m;@g*�Q-���\���ʠw�5Yo1[带�g��(�Y1��2�r��ɡW,V�T9�Dj�:��1ڐ�uۡim��J�j�b��rP�{Ǚ���Z���J��O ���x!R�k/hmo5�v5��s��Z�2�^ q�K���a�{����mb����X)�������N]���.�#����9���[c��p��wO���ts�5�n��u���S�{S��-�i��u�ϰVmw%o%a��eѣck�h�lEV��Ak���5���rX&j�z�۫J��t�[��#+f5U�+��/@U�rX���;N����u�v���^F�9W.��;�_A�:�R �l��8�95�cO2��:f��K�t</�*����&��N�h�}o�M�[�������ś�e���l�)�7��46&��;�n>�GS��cU蘦��Z�����e�iچ�q�K�רL���:'cÛ��\z={3����,�V��R4���Wۏ9p�"w�*��J��[z�[�����IYk��WU��a�uL6A�c�������妷����9�cmn���јvaB*��r�̧�s5�p+��{�������+&�%E�$:��u��d}��������_iϵ凛����/����b��W�j`�z���}�D�n�p������R̿���Q�(�[�����4�:fe��U�[���۰� ��w��9�DWq,i���0v�X���v 
��Bf�\�IJ��_b���c#�<Ȏ
ĉGY�r�땱bXS�ÉV=�N�rW@�c���;4�����)N��kVG���f'�ڂ�eKA�;�*Q9�՘�@��W��-�L�9#�a�P������H���dU�!�W�%c�Ť��$ns4�b���Ʉ�1�\:���j뮿g�kq����Va��v��zݗ��Z�ޑץK����T����{��{੪�/�����5Øt �xE1dU.�J����G�)1��ad��\V�B]���fk����9mL-�v��]�Pus�8S�\���wC�j� ���ku��]���r�]Z�ܖ�D)��ekknė�{��\{f�|�J::���}1�T*"Ax��|Ȼ6�ʹ�ٗ�$�O5[hS�����ďu5��# W|X.Gy�Gf�s���doFp)�ˮ�r����ﶜ5�f��ZK�Mr
�sr�gD����gM��&l�-��4�����.���tLA�a�-^Ҽ����v�\�W�k�u�n�Xl�53^���D$J�1\��\�-mZw��B�X�Vt�;�Z9�V���M45)�]R�[9��d$L67�I3Bv4��U��P �8��������\Ht�X�Q�C:��u;pe ��&b�5��z1�%�w{X�+n�%\G<	4�i��j�ԛ��j�l�f�]���wt����FU��kGs��&��#ԍ��rp�<�Lª�J`FI�i%ȋ]qVH�w!3qI=:�[��N9�)BH�B��
�Q��\t��=�G
Ԑ�GQ�s�e���BL�V��B�����zDH���nQ����$Yd�.�ҋ,�J�)jt�O9��"�%(M΁9U�����i(�;�r�UY긷t\��+�Y�*J	j%�--ɉG���!�l���W4��!T�GP�(҈08���+�q9f{��e�iFQd"i��Y����&V$auk(�D��,R2S2"�KPBR�����#�,��,E��N�8NHEDA)a]R�`U
,������TB$��%L ���ؔE%RWP�F�YʣAQ+,���u�5IVfe��%�$F�ul�#O1ʠ�
�>��ˎ���(�-=앪^��,����dCo���q'�+�ٴ��{X3]�nq⩍�����_s=G��}����K4��ߕ�o���l�׷�]K��xi�i�G�{eR�D��3TF �R��v�0��wr��ZB���T�Q�ً�C[�����]��g���*���xn�O�#'lS�j��Λl=��L[�KW�(������B�鎵W~�m��O��S��r�:˔�y����:ۮ�c���۸L�Jj�c�����c]JR���ӔDk{w]3L����^�q�`b������Vy~S�T5��6��hO����%�^����.��#�}��$4��hTy���˅����tuB�&�)<H���_U�$�ܮ\^٥��A=��ٌp���I�~0w���򚞣D�=�#Wym0���Q؞�x�ގ͢��io���r<-=�*s\�.�lDJ(��Zx��{t���:X�9�'l(n۴������Ύ~�JO��B*#���X���3.0C�a+O\�M���\y���UK#È����0��!{����e��� ;b�d&H�JTX�ˈb�g9Ӫ_�ƽ���~>�}���g��.�
��'5���]!��ҳ��[FWWH����M���_u��4*)ûs���,]�ɮMwK�����#�.���V_uj(5��b �*�ut�uwd���p��Kifb���o�:�unr��mP����6^�C+W��V]E;z+�kZ�3��������m��Ɲ~�+�>�גF��5���9�h�X����ٶ���u�^
�q8hP{�5>��M`���+,��
uE�yY�gra35҃�'���j`��0U�f!�ŇUw�c��r���Mr�-���F����:��q^���,���u�)��/��/+zuOD�V��K�]�(2ϹhB�O^F�*�ʄ,=(t@�8\T��wc��7AԞ�{NGM�5�mpP���P��pgz#�^�W��TW��U���*��ߨN��Uw���er���$ZϪ�� g�\�u�H��b���s��	�!�7��kf�\�)W��l����S�K�K�Q�w�1�����Ȑ��jN���s����
���4Ğ�Yw�K�Ł	���@�$��v���p��rل��'x+ ���7)������x�~|���n�Z�R��Բ� k� ���|����?��C�������2ǎJҒ8k�[��mj�SfÍ#���^�>�=>�V�+�d�\ˣ��ߙtMp�]C�=�����&KB��2�3)���u�KZ�SmZ�,^r+�s���@� -bx���|�Lѷ҂��2ռ��k�^!��i5�����٭��z{�e��z���Q������io��Iu�eb	�os%���UW�W�Wv̓�Ɍ�1��v�P֛�8�����;�Ge��O:I���3��h�����w���$�x
w��hI\�K������7��� `��L��)F��!˻��-����]�n1��b.*�԰����#^a��+�T&l���V�:�S�"��s}��u���֣���q2�^0x1��*wdl�L��'p�BLW���b��\���0ԣ���q��o3�z��/ƀҊ�ò�|)�<��F���s�x�����X��{�NC��WB9ï$~���Sy��7~UgPp�5�Γu�-Վqxb5|p��S��k�M3���TWW���ٮ#���׻��s�Qk��J�g�b�0Cj�.NJ
j�'d(�=S�H��T��ʆ ���/�UJ�8� ن�(H��W�\�7q2��}��B����{�M�77����W�{�b���iL>3qً♽2))�Y��/���Ww�֥@0W�6P;.��\�v�و�o˝��2W�Gu�����Ba��c}��
ڇ��Դ�[[��&R4��n>���S���l.��ʺ[H�:V�C�����t�=��;��a�]<�X����6;0��I�u�i����.�7W;����qm�Mm���s�VE��}�ot�:���U��}_P�;s��ۜ�wN�c�"C�r�CGC�8U��s�Q]{.��/R#YiI�Zo�]�GpP��_�4үW���A[��P�7�*��Ã�_y\V�pO�$֗w�7]r��"��O#�MSG]��vb�7�Y���"����H���b�*���;��;-,&��ރ���j��O���n�V���Y��@U.�h�׊�Ë�
{j$ �]VV��t{����uc���:n��RQ�\��O:�,��drC�1��~%�S���h�/.�(��W�9H� CF���`�Z"�b���{���oy{vD4��3�J�f�*_�:�om&n�qW:8��ɗ����]�i��>��U�}�GˑH�j�o��n�:��t|��Da #|�tֵ[�4���0�L2��̱�ݐ)K$	�+�����\�bb�TH��;��|0R3����φ�v��Ɛ�bDX�Iճ��IA�0�������B���0-vneo%sS�g�q�U�=>��;�B��������`�vVz��<·F�h7o�b�a��Ɨ0�ڎ0�n�^�tف���`�+�j�b���!���}�Rs�f��ܸ4F�76���0���I�������&���%sv��u�:��Ď��ԣ���6{�����b�Eg]������!S*�H\q�<j�|��ء~ ��$���D�d�m���7 MetOz�1�l�f���C��Q�����ë��H�C/4�j{[v�,8����Kì�F�#���J���\?rV��E)t�Ns�&�kz�ʹӈ<�w�s����E7��H_A�)^߮Z�[֌dЎ����v��Qco�<�Ҩ��;R��H`�t���W{d�ܸ֚��i��xW�*�N�	iW��r�O�U�������כ�c�J� �R�ū�
������F2�H���Q3	�[z���U+S��k67�+J����Q������P��c�]��x+�dl���e���Ǽ�m1����5�>��@Y�e-���Jj�p5��5�F59cB��C��U^�*�������g@�2�SE{2y�$gI�Ä�����d�8� G]R��7��A^���tb:vhG��Oр�(�ю�F�)�]@��yQQ�p;pC��=�iBN�����ۉ=��Z��=Q |v�X�u��9O}�zA7����=L][�
��������Q"���CG���A}��kx���g8�'a��ms�],.�T�l3���[�^r�N��m�u֮��|z
�=�1_�"=�z$����c]�2��}�&s�X�P�Q%I� w`�(��4O3�B0�'�d^7@����<{b�xX�>�u��:��hz$'���V�����r��U��F&���A�6��33E�}3�cr��H���J�E�xP=mހ�����J�����./��2�\�����O�h߻���j4EGrb�d&���Cr:�� 7ށ��I�9(^���ndW�Ύ�{{�`��|(�[C>v��\>ǁ�+����h�����f��j�h�T.�sS��ՍVetט�$��Q=��D�7�y^U8�(i����'���o���]��[%��J̥��Ko0�]3	�<���L �עJ�
E�]s��Tf*`ӵx�l�f�+�:��`8���c9�Gh�/.hWC[gL\s�nLpÓdYzPN�w�U]�JU��H���#_�P�5$^��bzU`���x��,�)��6�n�Ǚ*xY�7N[�`{�������`k����(�ų���|"���2h�v&���z�o�rRZk���.�9d(+�j�Q5
֮[Fn�*�PQ\�Z��}�޾E�7��8� ��|�O�x4끾J_
 ���=.��Y��G�<��i����8����M���aR�Q�=k;1I�|n�w��ʬ�aN���DG��ѵ���oGq��%�ϔ�|=|��T���lo�����\���;X�ˎɘ=�^c�c��i'��,�*'�����&y�eZ�-0��N�8+9�^��������[S*��-�Ɗf��_�Tz�@Z_��Ip
���2֎뭴<6=D��z����|�r��Q?��;{��g�\s���K/DH���U*@ޗYj��� aI���,A���8�O��dC�:(kM_�\Oq܂�0ݼ��_g�������Q����t��m���n
��M�/�eK�yJNF���v�{�CM[g���J�"��N�[U]��s��v�����2�fވ��/���B5�*!��*�T&l���� @܀��%����j����=j����E�%  �Ǉ���9��S=�b��oИ�L7�N�E�U����l3���OV��u��u퀝͓�fL-=(�S��G?�m��nvO�+�ת��f��ܔf��7I��Rб]�7��3���ϗF���:8��>F�y���A�Qxb'ۑz�g����m�:�m�R�.��ec�Ӗm3�f3��؃6F��[�	����̮wM��*�T ւ�]�+ꓙ��oBęB3�8�94�i<Q�hE�!կ"6S9ҀKoB�T��@�}��G�O3��K���Ӏ���QB�C�!TW�U"+�W���A���+�ߧk�nQg�Be����3o g���5�끛��`	JXbU{�]���T/��L ��a���#�=�.m�0��G��+���g����l^L`��L��S X�Q-<�C��vle����T�%un���)�x��w{~���Y�qg����?)�I�\���vɱ��ݎ<;[�Ӻ�]u��m����c�OܬV��l؋��������K<�c�¡�?��6z���>'ٹ孴3�Ev=&�à�!���W�Y�>n�Ń�M�
*���W�W<�' uM�v_m5aM�n��(����j�:�^�3�J!���p�����hS�U�W�G�8@��hbɱ5����K-��-�cg���B.U��C���2�����o���&8 }�H��<�ܝ�>���Ed�p�Â�e�45S^@���5Unn��ú�QG#\��Y�H�=r���yu�F��O���9���jvb[����=Y"�V�n�$�{�c�҉Tn=ǭ>ca5�r�\��?C�	۳F�{)�Ir� 	W�V�%��]���f�t]_v��K� D�f�`�*�n��j��n��Y+i���iD��U:�B&ۀN�����o�{����������QP'�2�;��Xw9��J����.˾����9|�+T�5��쨻�k�y�oў�Wr~7.�9˩��s��JH��3{�j�j�s�����7�u7b%1����xVJ�� O%����}𖓈[�%��:�5'u�C�]��r�YffAE��lu����Ӓ�,O٘�-i��Z��{^N��rCj#S���P�ve_�˳j�Am�� ��-���E/i^i��*N���O�{���U�5S`們� :NWG"�q�
��~Me���;������^/��r���M���gB��{;���\���{{-X��mo��mą�ض>��3n�m����p��T���-�|-���{cep̯�Oi����N]�j�-�=x{z�-�&};a]�_�y�Ž�x��nJ&��m�s��o��Q��9ۖ�j���%g��:������(��JEgX<%�Zy�5��}�����]c�E����7|�X���ᇣ�g�^#R6��M�c8(�9��+
����:�N�����b�:vZJ}����2�=��Ws��W��O��������:���#~���̓��'�A�Yp���j����D�~������20�C�emc�Y��R����zvD�8��m'e>p���t��]4st2�~�q����8=1#]J>����9m�p�:�������_k�O��;�S0{�F덧M����wB��s!.i�����ݩoai�����N�1g�I��Q��쒲b;�J��}a�×c��lsB�\n�P޷Wuuy��^8�n�yz*ޣ���.��̫��T���`q/;-�[������z_D�u�y
�ؘLps#սwi�\���;�0������{rku>�2��O��
�J;k���w_cz��G �x0��5�~��k����:y:�����O�EF�~v,p��\���ܝ���n���O!�Ek�4���z�Ţv;��{��F�[��X�:g�]�|�����wf�^Q� ��+��uԞ]jS��ʄ�����s���y���6ѷZ�q�އ��T�k���I���l6��6N�Ŋ�Z���m$ ��_U�p������WQv�J,��"wBv�0�,W˥�
���&�k9�LwgH�^m��C��<�)���f��0�Od�ݜ�fFM��V;w�Up�e�ø��.�i�':�urL��Mɝ[,e�;���aF���)���9�7�xVqnX��}$x(rn�Y|n�w}1pY;_	;�ǿq�����m��ē�-k��R���5 ��6uu9t;�{�V5��o
P��Z���B�������ۜQ[@��;1T����=j���ʤ2��帯�R�펮�%�+��d�����s{�'wɢ��p��;���Xo3z�Q�6��K����z�'%�-�u1P�B꒻������qJ�G;�0,�W��F�K�V��9at;��LE
���)֞�!�Ȭ�6���VpY�t����TyJ��w���j0%�V����Y]R�8�3;�����5OZu�^js�H�S8�3t�T�� ��+q�<Z���F��ܵJJ��3KB�S`�U���;o0_a�W���	�����9Fs�ݜq#�9��>�Z�S�D��|�3=
�ټv�- ��gၴU��Br��Wx4s�m@�d]�l\�u��oo<+:+���e
@�Qe(�u9�J`_6�=�h��j��J��yy�!�f��6��h���K��m̮<��U�ǫ%�H��#��h*%'�~��j��Bn���Z�Kʾ{����N��l���f��z��5`��-����}�A]��Z����o eʗ�:��Z�oE��/U�u]��&��n����K�{�V=�̥�R�;���܍E/�2\C� ���q�+�0�	�no��ճb���5U�Sd��)��4X�֡vQ��N�Ŀ���.�|�N|N,���_V���X�����W�E^��$7�o>�hp-�:��ݭV�.�r�qM��Xj:�k;��<0FŞ-Ė��#xT�d m�z2��J ��%��g!����-X+[�5��p�+�e^�U�.I���eږ�<M+6����6kOz����h
3��#tF����.<7q#�ښ�+���`��I�$-M9�5<M��8�}YJ��r�(֧;/�bʧ��	������su�٨�;u� EX7����䓦J*�����z��N[�*r��W�3�l�7[��]K��C�Ѧ2�Uge��a[���8buԫk�Y�lP��ǺCzZ��S�-�qЫ�
�a�oc��i4Kxu��I�Ս��O!����`S�:�u)��Sr�b��X�ǘ�����ܣ|��(����F�WWrժ���5���\{ck��Ns�I}�����#k#�[1ڣ��e�Aq�.	��d��Ii\���J�2�'I�}�q�m,�갋Y�����t�[/���6��P ,� �i`�BQ��j�mf�AȢ�T�4�(�®�l��D�B�"«0K,�L�J�UZT�X��I dU��U�I&qD�"H�I�M2D�L����E��i,��YG)u�ꑤhi�Ed��bmL6R��D��4$*��2�R"��IX��MG!"��.�I,#E@�:K�JT����*B�PJJ��$I@�2%D��da��dY*R�Si�J��\��3Ii��e�!$�X%��Z�e+U�TH��Yy9�%2��J X�d��QR-*�`�$�J�V�C3��(�eS*��ABK542��P�**��D���b\4BB�V�,��W4����b�eJ��r(.d����RH��,�B΅fr+�
��2U�Ȉ�	
�,2N%���:%WMZF(���U 	!>D�F��*�w����p\+�f�_ wh�;J��λ]\ �nv��5(S�Z�No��m�r�}�X뫕��ʻ�]��+��d�?������aի��;�b��ݒ��U=~w.�.�MuC�л�R�+�s��}�����t���0K͆�]���C&�Mz���mm�B�/���^[�"�xV.��/f�-Q���M�lZx�5��z��]�u����-�̡�+3rW=N"r����8���{��t�s[����d��u���ƴrj��~�(��-�J�8��NO+��Yp�{~z��\�%�W���/_/{�94�w��1�7�P�=�j%EkY|�B�N�O,đ)L-Wڎ5r⥮ڙ�q���O�֫�XUr�/L��=k�3�Nݨ�u�I�S/:�yR��/���5�B�Coj<���酵
���/	��#�k�7�wݡ��s����ID'���ה�B����k
N��f�����ݡl�	8�����kGr��R�����X����6�!�
w.�G�d�huZ��k���ۧ��n7/�2`nV�j���*G�ʺ�q���ݳ2B_Cp��VIos)�ӹ�O��w<�c�'�� =�n̴�BOwJs�R�n�[���>5,��/tz	�p7���2^,m$T���s�����꯾���7�M�԰����	�Et�@Z��.��)�h���w��f�Q�7p]X	^��~˴c ��	�Ep��yS��Gq&2%`��H��4_N�s���q��	�og�-�[
�Gj��J�t�]ݢ�(��M�mS��5&'��n�y�����ם�.oײ�n��w���g�����y�j6��̎k�8���'}p��-��ѢfK�?ͯ݋Ӽ0�ތ�u9�z����r�V���Ϛ�j���\�us]�+މ?x1�,}y9^����8�TظO�C&�%Hp�2z>�9��խ����}k�P�cx���ORϏ{�y���r�cOz/D>�o[~��N�IioÍ���ώ.��g杷���Ѣ���Me���':��.�}�?������6�:�խME�MJ|��D�7]�y���E��@/4��]��Q����VZ�W|64����N}�Q�Ҭ��Q�����5i]�.�i�(�9�|�<��u�7�R�L��M�G�F˕���44�"�f�s��/2��Hs��`X�*�����y����U�3��}g�\�5���!�ڈJ�k�{��<q�6��Ğ�[-]<�x�Q�~��}�d��>w[�zm��=��Ơ7�"/g�d�X��t^�9�Ip[���>�\*/�˅��[�|So#_�4�K���
�͞)*7�y�r�s�Y�s;�H�	p�Z�壥_t��:���4�n�x#ޝ�l[�C���4��Q���%<t'����5:vf�M"rۍ���8쳜���<�n�B(𢷨�9��bV�}��B� ,��bu>k/1���o�Þ�q�f�]�7B11�|V�A�]Z���WS�B�!f�����}�;NE��;�j\��e����ti��no���!<5����i�Ǯn��Qt���NZ����l�Q��cd�ά��;�#@{��{y��^b�ǵ�����m�=�5%p�=WG�A^�Ny'�hCg0��9zz5w\�ss@R��󝚻��g.�����ndֲE1��r�:�YW�z7�J����nS쩼�����BU�G� 垫NY|n�P�']���:E�e�]���K2�m��3U��+o��S�����������M\]��]�h�h��%��zq�E����r��o9F���a�x�⳥N;P�V\��U���!֞VOy�^�7(�����lz��k:��њK��J�I���&�<�����>����^�Ҿ�GY�>�,p;�g&vCSa���q�mFtc�ζ�7��e�o���d�H7hZ�`�����,y�[X�:T"%�og׵��8��W!�sb���Z��D)��R�n�uG9���l�-��O�fw��u���ܺ��|�ky}�6���ܱ�)s����>1�uܠh�d�k��e&+��T,��	>e�#+�7:�N��>�]��m9��P]P#�|oTK�	p�Չ�=����kqU:���l���)�u_�i_�kU�n1s�P����U�p֌$��f�\l�����oZx�����
����O@���͟}��	�x�~P�Evۜآ�)��!� 2��X��c�W�NW)�Z�������#�v�5a��YkO�r�t:�w=�u�X�t/F)�j�=y��*mL�4� i����\c��3+?J��V�U�:�(J��֊V��h�������j����/b��b_+��3�|�]p�+lc	7
iث�q��Vok�s�F
��cvk��{�Q��r{ɍ�o����mF��w5-���z���Ύ���&ޯR��`�xf"�W9��S��F]M@�:�ͥ��O^Ч�BY�7R�������R��y>�Ҋ7��.�x5��Z
�$����Wr�7��}p��B�;��d[=���o�%�5;)�g!5��)Km_!��}�t��=�nQ]���-I]R�֞��b��gu^Nv����&�6���b}}5�զ���eZ>��s�3�J�/3���ss���Q��s��)�p��\s�3Z���yS����b�}�w�N+�Mţ���'����~œ�}����IC۴j����I"�=��y����?Cq�TzJ�*V�Q|�B�LUe�O3j�Ry�5�7{��*-+7��D�������5�Y�X��^�`��̸�ĺ��4�B���r��]��N�w6a�����/:�T5G՝���c#�9�si��3.�2d�3s{yP؛�D[�ǽB�r�1>��Ç8��}�G�
ұ�%���_��k��{�5`]�;Nƺ�'y���Z���.��VJ�َ#&��|㚾zm�oiM7q��ۅ
f loTv=Fu�k�Ec��b��Z�G+{;4�\wm�Cj�C�V���N˫���F� �˙	��\��8�'�M慎-�3Q1�amo)R�_<�kB��s1	O]߂���鴥�NL�|���7Oe-5=#�rE�axd�F��[�q�=�2�UR� ��������)V
�	�*�ɞ��:�݁0��0V�l)��ò���U�n��6T�iU����=���I�mCނ�)��^����eVJ�|��9of��s��ps8��w�:�%eߗN&���R�<��*��z��K�F�Wv�wѥD�s���W�j3_z�R��%h���ۙpk��k.�=�)��c���ӓ]8������� �S3AW{��#'M��8V�,�U�5\9u�ֻ=T����/
�j�M�\Ow/o�tF�|8B/S��[tt5�u,��t:F�z�T��OWN�,c�1�ǝ7n�t�IN�Os\�Y��}_Dy���Ovꎋ�p;���*�[�Q��u><�Sb���7�t�1N6�sT�5'�zj�y��"�:���]Kƺz�^��o<_���`WĽޓݳ����[��lO*8����+ܓ�����.]�V�^��O�먾o-�|��w�Qv;����4��>/��l>�'Mo��Ʊl���ֽ��}���)���x^A���j6��ͬ�C�^f�!��.%A��+��W�Ra>k�y�ȇ��7}�U{ʵ*��Q�NuZ[I�b�952j�pbR�|��-*޻�	�~��^tm7t�a���4m^\,��7_�wHiT����
�b绒q� c�����������w���9Faz�o:0��L'Ձv^Hك�l݅�8;�'�{#*o��ٴ<������n1W�؉Hp{ �:�Ǟ��7Ҧe��Egџ��Q��4�h���[k�D ��0^:�[|9����էU�K�����J��G�'ww�Z��v�"7�;���ni�]ó�a��hq���
���i��X�u���>��)h;�u�KoX��w��;1  C����b�2��C����l��9��)��t��&���8V��-d+��c�[��'��,�z���Gb~�"Z��Ow��	�ʄ�;C낭׃���r�6�:���U��߾�z簪���!'��l�-�l�+�>]��i��[U�Jj2�m�������W�j3W^�M��Hv�+33�Y��mg'�{v�p�ʥ0�]~�,��u_[�7���:w33�;P�p�3k�Z�)T8��q|�q�n�y�^�7*죊�.s���]+��L�g�{ޥ��|����G���?C3j��{����w�s#4�3����yS������g�q����b��>ԯw�v�=������y<�:O>)�z;��F��d��B�����5�m�Mn;}��y5(Wr�X��Pħz7^A���J��֢�.������Ʒ����]�	��,k��Nf��	[L��֞�2cC��2'�8�|r����	�Xz�h9�����e�ٷ!ս��r�룧{kV�Y������Zc�
�t��z�[�j]����=޳n���vv��Ũ�er�UuJ��n����ݭ��$�:vw!������E/;{��r$�wѶ���S}r����u(�L_%��D��H�ۀt>��o=Mf��[��e[�fS�Au����[{��&zn�Wkau�fp�i&���~�4�+��P��FW�ͼ虛������G��\�����?w�ᒽ'q�y�\8J�T+���idM¾�%�UmR��y���������8'��]p�ô;����i&�6�q˝��9�������Y�f)�+rksSKF��a��L�����T��hd�#��Ʈ\%f��xf;V�I�5����}��1*Ԇ���������p��:�
�%vz�^3��Ɂ�1{F�d��W.x:wpK��_;�q�M����N��ױ�au�'�w����ҍ���w��'+1�5������U�?u�yᗶ�#%����K]{�U��&2��܏.�d\ا5uS����Ύ�b��.��$���*�/i]�d��&ܵ�$�^�����,���9��r�<�Ѯ �+Y��{5^�J�9��"��m2S��;��0)X��b�M�[H���5:V����1xx{���/k�Nh��l���	����}��z���	�B���>ΝyS�t,���;h/ۡ�T�b%���*�{C��]K���#��V��Jp�V���=<%N��\߉������'��_%%���ʰ%<tz���O^��;OѺ����M,��7�l�j%A��j�/�����B���]`������cWͦ���)�ɸ�����#]J����ɋލ|K�X�NcӻA��z���w	󡯲և�ی���h[J��Ț��r�VE��m�kcq@���#5
���h�of���Ƹ���8Ɉn���'�6�m����\��]�p��sИ��-0�%W���|sZ�r�p[/���t�6mO%�mxp�W��+�6fZ�vf_�JU�w����۾�{�T��MS�u�<�^�v'ȣި0����sH���U�M�^,�C���̬�"��6�1dkDf[:�[��U9b�4[�ṇɜ�d�����s����Mf�wY�����M��^������>2ֻ�����ϱ3��K����d�!c�D؛[ls4T�u��>ӎYƯ��Zo�g_:�)��(sWk|�'9[�|H��`�*��[*�k5 d'X�#�[ˡ�D��$v��,zkj�)֩Ƥe4�uͣv��:,\�n��V��q���e��aʸ%!��w(���Fv�ڳ1�9O�*8nS�H�����8�(�w:C7���*$RY�Mmjٱ�8}w��u����jۦ+F��Ҿ˱ORբ�z(vh��G��ୖk��y�}ھ��b��蘟xnߧ`
�lm�4�n�Rj��bC�`����L��ky7��Ua��C�r��g�$+yΙ����8�Coܕ+��e���z�_L���ڜi֔�vQ�
̑�9Jj��!iE�ռ�s\9ۻW5���� �k�:�w\�9Sr�۫��#�f�sy���tk����B�Y�5����wCW��P�tT^��/�1#�f�U�-��x���l����A��֣Y��k��Ԟ	􊶭̘��{���ʧa�68��1�xoٓ7Ix)<�Z6����Ӭ��͝Ž\�Ĵ������Xh[�@��&��X)m���J�\�ݎVЮkl���k2ɪ��1�3��T��9��qdm�|�p��wW����)�\p�xn�+"��e�vS]E�]�v��h��,��6fk�2� !��t�T���T�ifت!s��ôn�%�.����]$�Ua�R��'��2�R)Y$����suc��:� )������Ԗ�l�/�л]\>C^鷄u�}�*]��45> 2N9P�)A��T�k�&�k�-���a�)�źl-̡��c�g ;�*E2ј3(��f'&�Q4{+�Ln����,��Ds=IU��1��p}(rX(��%c������Qp͏��MsS�.fgP4���`l��Sca��<��S���o��V�f��!Ap�4��xsfnu�a4>ul��h�s^Y�Q��.�5kth����-\�魕
]�os-���{�k���W��U�-gtZ�ٵ�\��i�Cmc�߃�BV,\o@ƹ��}}N�,i��G-3cB5�"����c`?�6]�8z�FVu�Ȅ��RW����H.�]0t]����13�P�Sma�� �s#�,�G%p�j�*���N+��̮���5����l�:��DgbT� ��BL�w���ׁ��\UC�&�o8GDb��jd:�9��j�'�����]��sf�=�{��|�n
�+4&��"�vX�[�@���Xy�T�ͅ�ϲ$]e�cgN�z)��Ϭ����������L�fg>�yu�G
�<d��S�7'6:�c3��;.�+�h�6e��Sl��;�i<��0�c��EL����%�v����n�����]��G�o�F��|<?3�i�R$��֤Tet��T�GT*&iYf���$"̍3mT��4�BTH����Qi�p�M2�*$��$&��t�)Ye�Q�:(&jJ��Ē��*�
.jbj�Ь�TJ�LPB"���l�U%�s��"�Z	d���TRr�0���NY뗙� ��2��"L.j�
�SEJ�֜�����US�-
�4�3:uB����-2���(�&�J'1H̠�"�,�EJ���S���r����B�ӥ�����3&Qt��Y�TPC�\���i3�u��3b�`FR�R���M�fUUe�r�QL��C�⦳50�
��2���"�*�q3��Ce���=w���|�(WF2t���ś���\w�����h����ζ�m+�%eoJ��JR�[�xu�s{)�k�vŷI�ܗ��}��v�+e9g77�����6�������	�V�[^�wI;�Z���zj18192��m���ʆRLU6��U]ϧ[7���.�+���j`��"���o=�uoL�-QܝBtG9
�G{��]@\o�������k�<��W�%Qy����xf��A���]%�>�vƹL�u�&��ט����Ŷ��A}���޼���O�s��M���zE���ײ2}�F#}�~n�W�SMx���[C��v�1�M��|����q�Rlv��]�W	�ݼ�]r��k�����7�e犱��z��p���`gB�IJZn��~:�m&�<O��K�����hq����|����*?^�f���O>:�X�kr5��=I�:���^�e�&��)9��W�x�<���b��*YI��Ʒ|�.ۈm�)V���[�/�V,yJ�=]��7z����$tj���QC|��/d�6��V`~�]zau�jݵM;�i@Z�Uά�̰]�ޠ����u-w<j��c�-���۸��E��?����{d�^	<��6�-95d�tu:{K���� ^ت7Uh��WV��,
k�z=�̀��q�\)����:c����TlJ\*/9��Ο+z�M*��g3x'�
N�q���9N��������2�^���p���P�s�լ��OuL��d]i�r�c��S�i{��L%>����]��+��p��rB�[�n���ס�CcE���Y�9�C0b[ٹ�|fs��N�.owܤ��=N�<L�Q�݈�LpO"����zf��.S��	Z���d׻S�A�.v6���ך��
x-t�Ù�7s��9��j4���ѥ���oLǯ�I�BtG9�]ͅ�JOu9�{)�N�Vjy��w�j�s[Cg��]�@�3��c>�ޟ_b�2�]n��r�j8�_���p�n6a�uX���e�k* 㺿��P�Z�qg,�u�5���Ët�Zx�4/|�y��kj����6{h���OgLk�i]���"P�ð�l(�����(�����Ӕ�Vv(E���\�Y�Ȕ�΍�a��ŵy�`�!��9����7[R� �-sY�"^n�%��e,�����6*ws��ȕ��J�;{R��.k�n�?����K�Pķu�p�77�4K�E��5�Lʂ���In�6CY����殺o��z��������oF��<��Х��\:{�լN�vM����I~?n����Ru�q9vs�,㣎1\.u��M�x�ny^�7}��� E�yhb\�Lu�)�m��!�=����z|�g��_?rߏ�y�w��5�~�Ӟ�?wM-��|��5�Iq�z`��Q*�QQ|�B�N���2t]Tv�z���K������v���.j��v5ԩI��I����m���Ft���K��:ﻝ��y��ۍg9���B�}!��pxd�"k���I�#;���v�k�-��W�4�J�5�r�c���I\
G� Gs`S��U@��CY<�WL��'}3�݇�ִ�[�]m>A�F�*�`�U�S���r���<�Y�pڈ1�b���/
��	����;�x�H�����i��m�\�N��7�뗕C��[����;��91�\�X���f_m�g
ʫ�V���C�x �l�6:�
Z;Î�y�{Lf�չ-�;��HѼ�=�m<�3vr�T�H4�^'���G�1��B�W;��À��]ˍ7K&�I�n�Nná�^V�?gg��y�V����V���c��{���^���c����y�F�˚x:]1Y9�l�ݣ��UCNZ��a`�u׊�F�T^b�1��d�A�m�s�ǒ�..�����;�pԕ���D7��+Z�]A]�7�*��Gg3�9��=I&P*��^mՕJշ��4:ֽ��k`�S��26���L��r�Yc<-��c���[�}Oל�b�6.!<\̮�UʁӖ?civ�4��KJR�PT��ٓ[3��V�\�n3y�����q��r;��gB���=�S���V���~m�Oa����>��H�
��E�M��r� �S��m�ks��k����;����*�ZP��W*Y��;���5��[�������t1��m6����w���pv}�^2s��B��X��u���2�Z��'�-�i�j��]��F[�6ƹ�=7R������������9�����Y1�d�I��:9�f%1�n�дfp:�b�Y�!tf}��U�s�Ϲ݇�Qۗ�c�2W{�I�̫�.Վͭ��p�e)��v^=����Ш�!�\z�.��%�er�@I\��ĭ���[�]����g?&g��w�~�q}S�#�
��X�w%��কÍyQ�6$f=S=�ɵk�ΫP�%��S��	d��>��\�֎�}�J_tuݛ CwWy�ڥ�S�72-ӤjG�s�	W]߂�ˎ)��|��
���}��SYv\F:M�;�\7
}N���z
��Ep��st��`�� V��;��g3/[����_@x��*�����0V�x��.�ƔX������V,���M�\�?'A�LSơ��wg���IR��=ݸ�u�x7Ճ�
�^b�Zg1h������u�B�m�r��aZ�ʹ�r�ݼ|�;�#@~��ʃ��-l^=����vr���<�Du�fS�-��;�z����#��R�~�oЯ��϶��[�GހҞ����h͞C_���̝��Q�K5�k<���%��]�=<��G�W�ڍT���X-@�0�[��Jo��K�/J2 ��J��0�B� ^EOV���=X��{b��R�xp��s��v�
K����j�}���] 8����$�y�	Yntp���v2�'CxQ$�*8mR��+ ��O����yZM�0�:����K�Z«��')��r���^j�i����PU��D�9���L�^Kܼ�Z|��z�愞�]m�ب����+�n�o�`��4�������W��0We������NW+�:�\k.P��7��=�D�X�e�U)�n���v|{�Ԩ��2��N�S�p5<�zo@:�E_<��}�$w�������O۝B��^��-Э�1+���p�[Ѧ\�r��Jm�]�u#]֠�ʳq��L�̹��N]`xEO}'��h6��Dd{E�t�;^O���n��8��S�b�>��%1�.*�HȺ�Q�i�:r��.˿=N�%5�p�G7�-ؘEo|�G��3�0��O|��Zo=8�����r��6�S=�!�st"s��+�o"l�~�@F;�^]�>���>�E�}؋��^$��jf�a�'�&9�٧q-X��¯)�N.�+���+{:��[�ߛV�s��Ϙ�/g+��n�&k�g�f�,���&-\�s�rb=y؜�[ӅwtjĎ���j����{�qc=Ћ8��Hyk�@J��]�o'�+7-f:n�K��e7�����X?k���(o����-��)YS=�`�Φ6��hh����)M��y�R�����q��������ĩ7��`k���@V1Ք9�=�.�+�S�a}s�YƋ�|�^�;˵|��7R�V.���e�k(㺋���������[o��j16T�%;)����9A�T�o,|D�ʏ&`�z�z�ڡ�Y�;�9�~�y�:1�W��Q�;�}9�����M���o�ݧ��^[�zƉ�v���(��ew+K�ͭ	�{�UE|�3}W��[關ؾn���-.`�����ﹼ�ύ���S�&�߇{��3�Q��'@�Y������̇&�B��=͞d�dK{Z��ov@�+��J�:�U�Ui01����0�
5�X�J�j;r߃���k\Rr��z$vj���]DJ>���<��@Gc�[����.�s��On�v�?7��4��ܷؼ曾6����ތ�7.�封O�����`��ǰ[..��F�zLTB5h
<.{)�Mw��Z��&c�=D��9�wSX���س+B!�s�
��
��[��p���w���n>޾[.<�v87G;.�f���ZF�����԰]���~�g6���
��-���ϸǛ�M+��'�72�R�Gr���Q�3���ve��Uܽ҄-q]3>���-j��Rή�������q�kb�;lf�y՗ͼ+�!�5��\Jח�E��{�x,�`�ZGr��5�`�H����ܦ8����[�[��b;��lU�7)�<�!8�U��=�*㩻|��0^�[W����Ԣ�7uf彥ԧ����������o��5)��LrtV���@��ra`�k����bϣ3��}�k��IݻjJ��淔�+���p�:�R�E�� ɞ���V���N ��-՛����^����խ)��ør��qΞ��|��./B��xq�E�U�ͭ��׮'��ظ��p�,�˨��o�<<���z�e��Hfo5k~���}j8�~>{�u.==�T&��N����h.J*���N�;���SB���<��u_d�Y�����"��W�m�N�V-�spl@�����2�Kʬ�� �ބ��� ��xqi`���5�$Ffk�az4�vJ��OL�+����d1����C�Fy��H~�ǿyˇnC��<�3x���2x�Xf�����n�ݔ��+���ש�/;��K5�댃�W�Q�{�'dXj�j�I�ۧy�Ki;��8Ư�Mv;z����^.��A�J�
-ͬ򮝽>�>����C��3ݵ�K�ɩ�k-��mf��m,�9;Ǣ�Ґs/Z�d�,rp��65d��	p���;�|�׻�������l���/{�]E�&�*9�Sv)���	J�y*�v�O���/J���%�.����rͫ�p38ue�5Ǌ��A����0����31�[Y���H%�\�y���MyΧ~4sw�؄����&�_j�M��%�!��׹{��Z:_�s���nRa��M��\p� |��}ѷ��!���\��˹ڞꋉ�ﷰϻV�A�'C*b�P���uP
�R��t7��ByIG;�r��~��,8D�ZY�N\w6��8Wrqޥ0Ҽbe��CB�����	3	�o
R���U�����n��q�ɨ�rwr��\��.�h��ذ!�ڶ��b%�z����,珍��e�6t/8�výx�U�O�]]�XJ2�K�թ˩X�b��6��[�1��M_rwQhW>Nt��H��Ǭ��vG�����z��2�
x�̯=O���}YUݾ�����!6�pD7˫;�q��5�����[b�+z�/'*;S�w:Nbn�]��)T8���cxи�\��v����S�Wg:i�����	����h{��W�x�(��&�<����u5}4��u���V4�	�,s�/y>�~��
/Ohn��sb���rW��ި��kx��}��g(Bxe�z+S�i��+��T� cYm����w�����構;UJ\r�����Q*N�|�-�i�c[�p3�[�[i��ݶd��j_+�B�2k�J�K�sV��3z1�ȩ�|��oU�%{lw%~���d�M�
��;�$�6�����r���8��,�63 �H-^tg8c�ڂ�H�<���w��Q�q"���\Uv�4��f�7o)I��YWX�����8�z7Je[:�ouw"�)+�[�P�p=_s�^S��y���L�r��W�.`"���@26��7��r�X�N_����]��l����K��+(氳��DՉ��ݒ�S�})�}�9����cr�;d�����v�,��������s��S2��	�^vϓYZ���IWI^o^,*P��e,��M�� ]��O>"�T��%��H�O:��Z.�nb�z�ʳ��y-�7��;N%�E��cVMb���8�^x�C��'�X4�:3�Cir�m�������m�˛��ϥ/g@N�7�Ev|36���q_r�f����􌏈��+I�A�,�Ҧ�e��m���s���Բڽ�#�j����,cEf�"�\�ʕ?�ś/+(TvrΘ��k>#�3�6�װ���z2εse��Jn$�k�T���M�];�-mL6㭽噲������H�CL1�^�u�7r�4Scn�->\s�+��]X��k
	�ѡ��.��iN�x��;�Xu̮S����0�3�T���b���pU���}����Y��E���p����*N���*�����f��w%B��۬U�;�t�+6�xջ����g9ge���81�s˃)j�fe��,:��S�忈��p�t3�o�\]��wph��(f�M�˜Ͷ`#�'�g;��ԩ�VtwөWl�i��;+Nr���se���,�g�p�(�1�E��Ta�Av5:�uVڔ�}y= �$gΝ������6�����:m�2��6���a��b�l1��Um���Dsw4o}V�Q*�����������K* 4NF��Z�T*l���T�=]%�En��xCꂓ�������`)I*��1�n���k�����2��(��>�+$�;ⲵa�B+ZY�YI��^c=-V�T�)Ge6��F�jf��V\r����i����[��i~-T��<e�ѥ~��-X�
>I��k*hռXsa+�[����/�r���ϩ�Y�W|3m�!�#b��-Vt�4;�8!�S�m\ ��j�6n��ڗg�8���m7ӽ���Ib�*�oeTr��M��ˬ����O��p�[2%JWB볖T$�n�����"�v;Lɝ�b�q��q�.�9��\��_>�YYh$/����G6��|$����
�ݸ̃���.�]%*�sE�e�NIr��:M�89,�d�\����T�����³�#�ﲔ����Lm!������iS}��ý��W|1]�2��y��D��϶��Wu�M�K[-h��%W�v�;��	�di�u���!I^o}�C�!�J�.Ų�ƲTrv�sI�{|:��^k�/o�R!�-�6r����<�k����jʺ�>�x��N�U��u��*��A�x5��(�Vf]�t�EӰ��hGeD�ĔB��aM:U����)#
4.S)���r�DY���ZT��ʤD���q"T�]����3	,�B����b3�e$��B*����b��H�E�+Q#i�#*�"�H��DsPZEVp���
���)V��B,ʒУ6�TE�N�.��T����$*̊e�]2�"9���%�\�����aj�	dV�J�b�2�[B���E��U�(f	$�IU�H�1(��
hUQʢ��(�����)"��Qz�:�/w(�n��ʧ8��;����E|(}DP&�	�޼$i��%̜�!J�����uk�.��M_C�9Duu�Ֆ��ն����$^]��hX��^&�L�ԣ�o)}�#��]��M+��ݧ��6��m_�d�:F�G�w:0�H����[��w�)o1ӻe�>뱽�}��<Jh�Nýq�+t1x��7)��qH���:{	�FQ���b�k��חŭ�Gr��]nR��ቚ/���(Ri&���q�	�z��ڋ`�.ٸ�Ov��ʆ$��p�b�6�p��r��m��q-Tx:yk�4��3���Ůo�=�3gN�}O*<���b�Bߚ��CYj]�O���+r��;�UoBL��>*Vq���(��f�;��X�K�p�l�wN
��%�Z���f.�GD����W^_�!.���OF=Jz�Kp�������Ϋw�Q�nP�)�(�����T����;f����]��{z��B�[^}}"߯�✗��}��{���*�_����*�8��V��+���.�n6f͍5�m��c~�p��bKڴ����:ʧ����q�p��X:F��!�Ҷ�OZ��N���o|�.�������3Yl)����#X���8���z��7i����NhhvHw�����s��������T��E�z���'>���|��T��8[=�&���o~����D.�8���Vo�=d�k�^^y���}����Sr��_���q�z|Wq�Pb'Z��䫓�c���C�ǘ�y�:7u8�_��]���B��7�iA�9�'�h=������q�ԕ�y�{|S����5�K=�m�յ���q��܉�)B7]VboqfSln���zdf�Qi��Z9_l�M+����2����2o,��c�=]�7�Et���p;����j=P�t7z���ZuB��{���|�nH�yV���y��ek�]w�4����J䍓��m$�{kf���:�<�Q�&8a[��SV�m��>�;^%���~7;��i��tp������O![�&8L��-�^O[��i�T�a.�oM��������6��5/B�'�뢵����aq�=37�HKu ���5�r�rUǏ7���2�R�k{��dç*A�����,�G�V��S��jV�׾9�ό��h���Pg(�B��X��q��&�u�SշåmJ��bǻ��nE���h
]b+�G�.���0�޹�5����ۿ:U+�';�K��Z:�+jҹ(���1�}B�z��k��}ד�����䩻khc�X�q�1|߹�?%�Q��G��o�q�>}�NP�Q�#�R��h��5��i^UjƆ���筳^��'f;F�|�g������ԹQ/N�\�s7�;�{�':�����S�{�'U�o�Mţ����Ⱦ�U��s0���{Hf3� ��c��k�'����=�Ÿ=�����L���<d��}�N�������8�����t��	ˋ}kͦ���go:�n+�-I�c�쑳5��WwQѫIp\Z��������(��O��)��[��U9Pё������Ζ�˅0��9#z�\��U�X�w+{54����GeWNSI۔��`�=�Ʉ��T�U�:Z�}�����Gzu֔n�����5�v��%���k�\"C������^�a܂�nVY\ Ǧ�|u�h%b�Io1�Z�q�B����˭L���u؇���3����o���u.�RY�7jg+[|wn�E��u6����T�H.�n����}�o^�;�ǚ��n�9WW>�P<�,�N��y���E��`�U���yysr�a�5.c谧x��ی��J:�x<���o!U��<(��	�V�0���˳z�`�[nowܨI����������B�v4-J�̌y����Qe	Z�/����>�ׯ�t��F�Q	�4��x��7�c#|&�7؝�����u�U�*��s����:�
#�ɳ�t�\Ƒm��%8��W��	��:� �ʃ��/1U�ڌ���^����\���&�s�F���t����n�m��ml�G�[�W��o]p�5��ݘ����^wE�lo���ᡓ��y�l������YVFf�:J��?T�<����z�?�z��s޳�T�U˶�����p]�p=}��r�W[�;�)�&�ns��:�|�뭸I�O�U��vMH�M��_�U�To��}�b-�5�M�]��1.}�uN�N�YF�8�6�؊�r�-Ω�J�]�-�-�b��38Y5���Au_Ky�q��A�D%���
[S'����z�'�Z�m�]7V>�,8quu]ъd %/e��sy�D����9GZ����{G�iQu�TY��nU���ci��VQ�W&��5Z�I���Bq�{���u\�����r]s��N{�l�Cڳ"!߆ys�=� ��I����B����F7*�.�]�;�͎TC�}��9k��&_{����8�n���7�J�.Q�1'�gr�"�����6}�s8ɛC�'�Qw/R����&�u'�C������\>���4��`>Wpe�v��)���7�\8Jb��pU r�Mn�v�Xu,p�5��6�{Pa9�%k���P��I��s��<L�D��~y%��W-����b0��Kk���]�^����r�uTh�9K=�SS7�;�<�a=jT�7>|�C@Z��ڼΨ��b/��q���)���s6i��M���M�5|�򾞸o�_�ߊ]ي��O=:�����V���&f\�CiWl9bəܯ{6�I���5��M��VǦ�39MA����]� �>�a�V�»fNs�n���q���������u����#ˬ�=��
�k����yQ]���f���V���]��,j�f�X�9��ee�un�r���;������n�S������^������+��Cߐ���ժR=�o�)=xg�OJ̼OM��jx�[C%���5�0�U@�s�3���T�y�JQ����Z���mNTv��y�k
l9X��юWX�_Z=�ӯ����[گKhq�9ą��8��V��߱63�kxV,��h]��~�f0�E�e���+�nF8������g�ʮQV�r�2���Gic���r�j{q�C[����ˆ�w\d��kҠ��Q'6�tr�����m\�L���q������jyx�.t��.|��BePt��w)!���m[�@�v9�v\���[_R�<���_s�p�n1��t�z8�H�6�aV�����\��#�
��_�pU���Ҩ���,%�,��YB�W�l����;Gn!����F����Ձs�Z�ĥ��j�v���+E'��h+I����uģ0�>fup<P��q���l�t�/b ѻ�P���T����mm-x��>�cY��Ƿ*��ʴ�ዎ����]a+u������]�3�*Ik&���N��k%�j����}�����ޱ�{�Wf��I3-��]����%m�*{e���j�$~��f�S�}�:��STu�l%��UMC�9���n��&8L�Pal�S�&�Sy-��x������q�r�cil�]	�WQ��	�c��{���Sc$�1��N�X=�f4j�d`����V���k����+�t5�r� U�6fφ�e^~I�̝����w�&��h�	s�rw��O�RW\>��ܻ�u�A�� V�f'a�))�u�N��E����ߵBR�rZЯ{���CC��I;�lv9�V�V2������]d��h(w�ϊT}O~/�Gt�f��w�;%��ץ�������mCim>���]��}�.��n�W%�p�ɼ��'z�"56+�M��M�*�^�]�ʅcf'�7�>�����ӊ<�'Κ�|�>5�'�}�i7��5��k���>��q�x�k�*�ڹݽ髁��8��5��Y�@��~/�/d��aY\ǭl��h�:U~��^���<j�n}��z�5'�Z�+�3�WdQ�ދ����=ܪb+���,:��};]Ka����3^�r���ƚ���t.��r��/���P���}[�Q|�-��r��[�5���WW�*����:���k����L���w��IB�.���p9�z���+9+F�OSG��{4��aj�tloT��	p��n��{=ȏ.�{�,}x��>6������v{^�9n�3��[�R<ls밹އ�j���|ojY����	q[�5�/���
�d��#�B��� �A�]ˤ��k���ܻۨz�;iu9���p��w�s� ����j��K����j�Eԧwǽ�63�"���W�c�n�͕q����.n���S�㷣jMrɒpZ�;��O���v�}���\�m�bfP���>.@�zb��7{���ض2��\6�uE����9�*�'[��]�<��Դ����۞��=}B�g�5��,b5��̠���]�W���c�ͱ�r���Z��b��A���'i+����]q/v�S�T,�>�3����Ì�'+}r�^��2��iN��d�X+�v��G<PE�����]@�3�\��pHGd���u}o�.K[�Ê�U��{&�N*��wt�j� �.>.��|�+�ݙ��,�uC��w��W�8����X3X�lZ��T9�qbU�N��p�<@sԵEu'��޸��l\'��������r�6�UC��Ӻ��E�H|�-9��"�-5�6�b�Z��v�����5��U4n�2,Cb�Xuɾ�ÄȺ�Ѿ�i�v��g7Гb�'ګ3l'�C�u�L<��T�I���v;���Ҩֿv��Ʊl�oR��N���a��,w�y�W�4�z�{;���Ϋ����Q��N���R}4[���CR����gRˈp�+ͭ��w���P�Fƺ�R�Az*2H��3]��F�3���o]�ҿc�ێ/a�n��O���d�5�����q�C�"�L�[�ߖ�[�gasJ�;�X�̺G�"u9_.�֓���!k��}P��s~�}<�.�98e/�]"�Z*�nN��ˋYX��y{Þ��4�J��l�j���!�()�]����,�0%��"Β!��#y}c��GhD��Y10���C\���l̅��i
x�7�J�l�@;���9�H˾�*X6�<a��=u,���5��m�ĺ`�\ӗ�f�I�Ϯ�!��:K�2�[��
4ԎĳU�X�/���'蒸�����]"bi�}�t�Lw8����'���.�]H�:��Td��u��,qE�^Ȋf�[%��$όa߸��<��4��;b��G3}�[EXa��ծ����	�#�>�����?:���������I������F9KW醴�eB���F\�l��pP�;M�a4�3'��(�۸� d�4��_���nnP��om#���|�ͼ��̞��n:m.�X��@J��\���N��p�U2>�rl￑������ڿ�`��S���E���.x_��Z]�N��~�u�3���Q������߭��u�-YBu}*�ܞ+si�g;c�h�`��:�.{���&���:�)<Y��f�����"�%����3�̯��d,Ο�o�g)��c��?C�*}�a����J�[��+1����}>�$c�N;^�Xl��-j}��°���E|?��/�!��v��q�R���y�̠V̎�o�(��EL����)f�V����Z�y�&FPX��׭?#�~U-ի�Y��W J�,r3qR�^����70ok!�[���^��R��<=�_V��Z�wu��U�fP�>�d]9K[l7	���*T~�8��a�� �m�d.u	;�F^t�v[4wV��_N��s��)-K�u;��ǪN�OXu��7o6�~\�H�z4c%�a4��Q��Zu^�p[���i?G�,���GA<8���Ɖ�H�]\>�1o�wJ��ԙEv�}����`WfTL�&gT�Hdv��}�J�2�=�3�l���ńyP�Cz��6t�2�kXgV�{u<�u)��+-���[}��jSz�=���D�\e'V�;��r�Y�1Z���ބ\W�C�����F��Lv���V����V�(�/���l�잒1�ޮ��V��*S�OMi�>�dS�w�*,��RUw�����./'_Aj-��,Y��������^<�e"1�+�A`͚��{����I����e��w>��TM��0|/0n�ka�[]Gǘ�b�/���ثWm����ї\���u�)� �5e�$�RBU]�{�6qb��ݑKd�fttD�P��yW�Gp;�ֹ���bU��L.����M8|�*d�U��u�J���n6t�B!��6��]�w��; E4�7DV����e9���CX���f�3�qÓ�Z�U�M��՛���ǺW�٩N��Pf+TR$�k:j��q��,V>���W��M�|�Ǘ��v�9��9H^�@��\�i��dU ��r��]��k)p�]P\o������e	T�3i�း>ˬə���\�vΛ��:�U%��[�&R�q��6Kʜb�E�%�6$I�O �1Vz�x�ى�d>�U�޳̧ܫf5���)�/�2Ofj�뗘�������ߺv��4�6�.5uf�� �D��L��۽vy�[���2��kaV�랾@wb��]$moZͥa��N�QV{3���㫊��Є�{���X�Vqw�+Yz�7ko2��&';������C�6�v��Z�@��Sr�������A����g��gS�Y��r���u��q�{)�Ɋ��嘵VJ�x��2u�2�&#��@h��6�ǅ*�z�y8R�B�b/Uep������"�Y�ޠ^��R�YG�B�f�w��'yƴ����"5^틕o:���%��i[�+J{��x3bio�9���6*!Ykg2���ݧI-�\-r��p����D]�_wM��*U�y���9H�����>�x�ri;��C9���yEn�i���O��/bw�7�)�++������;!�}��&��<�oI��xK��{-TS�0��O0/�1N���;z��x�<P�sj:ǯg\Df�X��mH%��3���r�:��h��]&s��0�t.`�ckW@�f�s�\������+9�2�����aAi�Kt8��C�4G7Uí�����T�$��!"����}�p�PN�&s�9�B� �2"����X�h]̗Y�AÔ����M�t�UJ���˧J**�̕.I��ԕ%�U�e���UVF�$'(.Q)��<�I(�s��E$Rd�m*��s"��P'J괒�.	4��&G*��U*
�̏J�9IĊ���SS�%�ܪ�:fs�I$h'bI��S��T�8��J������h�f#9�L��4�GI��E^E
��aM25dQ�R�EX�d$\�5 3�b�XT�ÕbR���(��,��$�6�pU�I8���q3�X�eʹp�8(�U9��QR;Q�UE	#�8Xl��4"�T*R����r��I��;O6n轙}Ъ�^�����)�f�=�'s�+���I.��3aﱫ`r�V���LB���n;姝5�6��T�Y�r;�!�`!���Q�6�Ca띎m�� *�ZgX��Ŗ�-����'�[)�y(|��۩
῭�)�����R�V���
%HS��q�@���n�����0&QC��5�= s���W�l�o���!Sz��t����9U�,�}�9��Z��U�P�e��+<��t	��W԰������<����s��{��L=�~���őt��p�^�s�jY��)�5�4������ƭ	��S��H���.6,>%JVd�|��6L��c �zi6��e)L��J��Nt�ߛ4�6@���J�6r��a��ve3�q�N7\E,�u�+�a�'~�#y4�%�(׏΀��@]��d��?$��b%�GE\�'�j���/�h�W/L��ϯ�5��M���U�B2�U��\����dag3.6�B�șe�Z��Ps�rC�&��-����9�fgN��~e��M3I��(�UO�n��Gd�7�������� *����i�p9H��<.#6kM���ζ ������A������Lc<�ȩkeJ���ή-\ᕊ�ui�$���U�c�u[(bx�ԩw�}��������;]�5S�]0)dVt�]� ��ȁ����i�c������S��7�h�t�ia�W�Y�u�����r}:j�3;tUvb��f�;:G���pc}���Z�7��ͭ�I�8ra������i\����L��6�tC��>�5[3,���SJ,�������t`��t�����QQr9"�
��j�y����v�:���5��ޙW�Q2����n��g#�Q�%.p�*��HA���q���(�D�6*w�t�\F�s��w:���'�Vi�r��ۓ�t.~��,*޼ߝ�Q���`��T����~�����T��*��j���]�~
�a�sWM/�̗��\���Z��7����lL�Q�}uL	��G�sJe�ڬ_����馁n�Y�eg���̽]v��v�0��5_��������k���&���D�a_����덡�*&��}����ug�>��M��
�7�E}���T�`���Cgb�Т�����CU��4���"�X[�}�o[��F��ґ^?}����|'E]:�jeIv�q0Xsx3$�ǌ鳽vsp�ߐʻ��S1�۷�k�E.���QEN�(�}����)̹(�<q��잻*��,��I������J�F�s�զ��mM�xe:�;l���Q-�U��3/ΕQGi�s�ŋz*n����s�y�̊�t=��3�(�g�,�V:de
ӂf��sFs����7��V*�t��W5���S;�Dw]��O-�ԧqG�%,w�r��R�ӣ:\,9|_,ϳ�4����W?'y�[7@��pY�bWJ��7��%�IDÔ�50�r�%��;%s�s�Ϣ�d�o�4.��#������Ӊ�nN��j��;��]E&'��D���SnV�"�NA���/ܞd�"���3bQ�S�_m�֒�Y2Q�J�{�3t���NxԻ�e�7Q������*y�9�W�k#.��N���]W8�Д�MAtC��^[ �%S0Һ���N��Ͷe���b4u�j'Z`*ډŮ�]b�
^���#�!7k��L�'�R&����_J���WmQ�P�H�7_<M��1���u.�!Cru�E��:�->{P֞�j�l�|�1�q\s
G0��dF��1�x�k�	���5c\��ߎ�;�3�Ǧ8�_���4�w�f�[��l�!�Kgs�3�[z����uv}�����vq���v7������K=�]6v��M���G�i�o��nl}�I+1B�Bl��3�m^J�H�ݟ^��Sq5	�W�7�p�B�!�י����@���n�;5����S��������Jb�u�S��\.�ZS}_P�#��m�ý]����cv����7oN	ˑ��V����j��{��]\ُy��;�/gt#�|)��ws�P�X��8���)�W;�D��jP��b�'6X�FZ��d@i�+Y��_}�ձY
�3��!��@:}7M����{g���ɿ�/����`�eUf+b�-�O]���Y!PnQ�jӲ;��h=�%*SP2�Ϙ�n�᪔K''��帐��_R�g�7����c���V��Чt�r<��ف*z�T��~�1���	����LL'Q��?�=��q�,}��p��[�^�>�zP�CK��c��VkМ�͚�*�h	�Ɠ.{ˇ�cI#��)�N�g��?3á�G+>{��p���yg�M��O���e����D���a��?k����X�:%V���9��)�dW?t��ld7%�"����+�V/��Ey9<MDL��_��c�r�!��_><�}��b�Z�ܡ4��`�*�(g�Z�	t3-<��L{S�4~���/Z���V�~��d�������OM�km��a.P�̤%�v'r�I��/��>�(�9i�����=�_�T���?9?���~���Zo5��g5Sҩ35��u� ��Qۮ�`�e�$3�f;��h�4�mp�a]�İ~�h��t-^W{/)�:�8ւR߹�,�ٳ�(�<��է�h.�f��HWK|�wڒ�q\t�mY{`u	:��=�F��kT���\��y9"�2�@j�����Ӱ��z�"r��w+kLK�
���	1�9��hg�{�F�kf�?�`_T�]��C��6R%�Zf'۳�sQ��i�^��P�ï�!���h닅�wMė��3��K3��@�' �W�oڗMN�)�F�M��������}�Z3墐��)IY�آ����̰�S��7"��[N��mu�oieU�C: gb��������Y*د��%Q O�F~���:om��ۺ��+n��)���hן��Tb�f��;���XdtN�5k�ys�Q�;U
����Ib����:~�� c��B}J_��J�{u!\4��+%B�q^A>ٟW(�+ky����M�uܮ��ڨ,�*�gK+�Pv@�u_Q�%���s�{�}d'��P�7�1y?��2歾��-���WN�)ҸC�l�+�!'R8� Q�h�UvBn��H�ay�)�hU�Cᆮ��Ҋ��=AP3^����R�0/��*�d�ZO��*:u��f~�#�n씐����3�]ӭJ6%T��t%6�� R�-��0��L�<قfy�
1����A�
ܺ�{�u�����/Z#��oR��z�>�"k:6��UCqD�r�n�>*��e�l��vbG3;'w;|��!�.�Z�F�[s�97�]���K:��_-YH;�l�",�Wz�1\�����N^U�/��U�Pl�pl�fk;�ФYzS���W���9�r�����(�]�O:�f���$�"t潶K�)z��1#w�C;r1͓W�z_��n'������\��F\J]���2�������~ō�Op։+��˕�d<�m�tzM2s�}�$V�s*Sɤj���q>�/Hw��\�,��u�qf��0z������ten�3L���u�5~��`m��B�GdI�*��mz�7���̸�&�t�eL�4�u�[N'9o!�i�n:M�R�>����(2;���ڸ;�5�݈^N�4xVu*D��8VE6��Ȇۦzl�h�w�)�,f�D�O�&�f��o�pp]#��<-z�:L���kO^�S#*�J&U�#��_\$o�<W��Q^��!i�a����q�٩b��A���u{:�,'\�lF���-uܥa���aMvpj���g�6��V���HƢ%J�Ds3�_�W����~e/�e�5�#m^��_55�W�8/�5���̶m̥<VD䋡���V��,جDs3�|��7�76��G�9��J=q˲u��u��1V~�V��p�q��v��ҬW���;*�<�����
���]1���
���{�/���&�)&r��_\p�����c8z�<p>A���*����Lrr<�eCE��q=|k�˚]u��rۖk��B���l���.
2��j�o�w	h�?��9��S��v9���M}Fr��+�����LDe5;�{�#x(��֠~�>�2���[G)R�+���bۯ��wn�>�xnW���)�����%{��N�nȉ�B��@%��x��%OK��yrU����GS����ӛi�F>^�C�j!���46�>k�#!rJ��Q��ϑ�'L���E*��{�B��{�3��+7�9�J;퓄��߽1(}V���=�Guf��_�4���l��9;�&:L���^j��md�%"��`9�:ja��Wı|���G9�c3��\�	��=e���^�U'̵�s%�)eᙰϯ+��ԐE�bV�L>��0�g��kw��"��C�b��ƽ���V����壚WD2�C�H�s,��z�@��MHw�˟���ӎ")��o5�\
ĉ��ӿS?D�L�Φ �Cw������/��$_�U#_I�]��8K�wm9�ox}HK�����k����W읭��.��Nh�L�+�R&�'�:M*�,��ݶt�DL�K�u�Fԓ���J�B�@�t�Ѡ%ƚ�{O�}����qwB��S����F�}�G9������n��nz�v��El	�]��]�KBc�+ݍ����D�)�k��sn��B�V}�\��4X�*V���h�Qlj�����y,T�G�oR��Y�D֊b����ǿX��C̾U���T~��vx]���%�b�u�ߞ��K6P�R��<��:��7ˡ����FR�IO�/�򵿩~�-pQ��lg�P�d֖.2g~;.Pj'�����0����� ��w��m�����;+�_���;�Q��%"C�6�b/��/�3������6�2*TDAU�aDNkb�2�x��Xoغ9~��P9MV�e,�f�v|xr���<fFl�Z�=���އ}�ey}�N��6��B�A��
�ءY�6^�����*c�NQg��f�����G|��iE۸�sQY�s�3>����=vⰠ:�HT9Gq�N��V��(P�A�<v��Ҥ�iQd"�7�'��3Bf�(霹��\����a|wQ
��Yp��H���q�iٯ�f���KC�m�.�#��@a�x~4ts�J��z���/%=��{��P�u��wc����3G�տw����N}������
r�"nK�&&�Li!�����Q͙c�cY�%�K�I���R�J�hk�,t��~��i�g'����a W��P5��_��τ�������1�8T�U��a	��r�'���{�Kx����)�5ш���]����,L2]	�w}�>��%��D=��������w���-��-�����T���A���,���2�@�{f���;,dԆj/n=����f�pΖ��b�{k[J�M8܋����d��S&�������52�}fl1�}�I�n���][so�C���^̎s��
�]ΰ�)hM#TA�;2ý27\cڜ��1htMkg
oC�[�.:��I���UŲ�}oVy���~F@J�B�=3�M�Z��.�&.�n��kjOk��%��~,�XΉ��f�~蜭�Y��oe�}_[ '���῾o����zf��)\�"��+2�DO�\�#S��V�6��b�,�q�Mi�΀�U�8����1)M�1�a\dC�նF��qȴ�KmK풇J�lP�!��*}�a�������_���KS��Y�⊒����� �ܮ�m�?����õy�����8d|�Rd�=%�=2���y�+̎����v�|2�;E�lvΡs25�22�����폲�\:x���Eg�@�H��f���}W��|�r���g�T�&����<��ɎD�.��)��Y�O�dmZ����J�Dʥ�����;�E���OH�~��M�ٸ{u!7�!�q�)�p���d(����beܼ�rd�g�JF/�T������*���C/�mN[-޾�2N���2��wV-�l��w������7do��+MM9uZ�k{���v�.��S3r.`x6nT�w-EMKJ�'e� �Ў�1�.�c��9,N�����o���.�7Mlԩ�D�^F���q�p9_���D�Q7�~gr!��r�,r	|���gV���w)����_[�@R3�	O�10�]*1PW԰�-�����T�Y���������/�]lP�������H��X�}r@�� (�O�ٵ��8���&U�qz���/��7�%��s��-�M\���ױds� >��>ID�L����^R�i�1
���m��{��H�{*~��L�v;��M$�e+��i=.͹�I3JY�(�������L�^�Z�<�6M\��˴ΌP���ЛkT���ur�V�}v
�=�	��s�e^Wk�N:�S�0�z��簩y�m�{��'G�w\�5�[\?��|+���U�2^#Y���/����4-e��uS�,n�4D�g�2��6�xT]�i�[ř��@�Z�߉w��;K��R��^���}��Ȗ�C����C"	�Q��ٹ-���F@��;�+��j�b �ȉ�9�ӱjx�k�^!{<���]*Q49=�ҝh����t-���k$�ۉ�3�5���ѧO��A����5�-��Q��x.'Q�7.t�)��}kz��q1kP��-R���9Y�ԇ�9�X��*�d�O��3��ɘ'4��]kr���W����Ӽ�����۱����ם�@9|	��v�Q=�\��*F�e�8���!��״^�9S�R�No�ú��s˭�BQ�7}b�wW�!����T,���)��wT�Θ���y�gǹ���q�2C\ �ِj��e(�r�l����2/;6��A�r��ԍFyIP��3WX�nd�^S˼����H�1f�S-%�S1=|1�o�cͣ�������u'�bO�c1%w�970V��!��2�>�
�"Ð�+�,�_f>G;��`���*f�����b��t��n����;sjIdn�u������Eӫ�&XT�d<����M��v���(��]xR� �)��H��k����n5p��F������|�m����7�w��W8��.�7w|�KɆ�Sֱw�gZ:���V�_|7+��oY���
`Y��f���uz��B�j��j2��Ov�k2	YEBZ�����z�G1�n������.>�o3v���t��1��U&c	���ܗ*^�L}Nڽ|�+���V��bV*w,�����,���_`V�v�j��8`�����O�J��a��w�NmIv�t������(T�f]HH��f����aI;�Y��Wo�1�-ά��/�A2[+��Vс ��)<�HoB!��1�K�q�: mi��],-��M��M܁�YS-�]Z�4qu�cjq��3��Z�u�
��`���R�Q�jCZ��q`k r��>)d�GN�`ޮ�(|JE�(딒͜^`�tt��Vw�k�k�$7�;�&c���"�93g� s{��Թ��e�suY�tbJ���u���W!�Wn�F��6V�Yǧ�s��.�E6���IY�sjE;-��{S�	�jP��u�LxI�߇>��ǻ���n��p�Ԝs�pPG�{�]�}ʒ��n�	`&�aso2��R��!���U9��P2�gt�|�FA������F�9i�6ģ8�$��6e����;O8t�X�r��32|4u�;y�V.-����vj�.j�&$�)P���t�n<�00�]�C�Y��Nb|�*H�gGVj������������!��Ӵ>�b��poGW:����L��^jKT��g������,Fۗ��)��S&^��\-�ه�]�a�W}���j�x���]J����֡�sr1�5n�����غ�ݸ$�`F���"G�p��I"�V��Ŧ5ݔ�VJxrC�[�������؍�A2�mG60^FƎ��#�`΂��k������C�grx�^����B��NPUS*�,�*��t�*�;%!$��HŬ��QCT=t��
�KB�B�^��QG�PP����s�ŷ:^��M���t�(���,�@�$�""ri�u
�+
��!3$��E	"��E©P�
���=����sR�T\��rJ��˜�G.�Ȉ.\(**
�Z+�T��E�r�
(
t[]�9t�*�.I��s�'
�̈��.�PNY	�(���2�I�P��
�*��$�j�DU+�rN���Uf�8'Be5٢�z,�fQw!/u�=�"��Q�Y��9z�:Uª2�9t�2��\�GdU^��r���(�J������ �ht�q�-N�rtB�]ܪ�D;��tw]�D��+ԣ�8Z	TT\����**���s���V��}O�v�J�[�+S+��v�����OGS�5{v_GO��WA+�7@%:���L�-*��:�S�=�m�G�����GQ�~o{?U�2;T�ʽR���������g{b�V\=Y2j�L�:���ʾ؝��Z �;8�H*�V�O�V�&r=<���w)Xh,~G��T����u�ޭj�y�М�D�ާ=R1}�Ol��#d	F��@��0&�,^)Me���C�������L�~:ک��^���Q��W\��j�0�	�Q~UL
<���L��R>�oY��x��V{�j�]��Q�oyU2X��r���z&4�[d]{]�8þ3����cx8P��v����b�g�F�J�7�p�ֶ�O�f�t�+֥��<��M@˖��f>˻��C:�s�*L�]���|
��t>�j������<:�dD��;����o��G�OK��9ۤ���d��U��c-A�স��h8��Sm��y�`B�;\��k	ґ�=�'�ϑ���;�T��Y?B��$8N!�شq�ǝY�c�Y��#}�0>U#g�f3+}&�FM���3�κg�N�3l�-Q:L=�e�e:$_�cӘ{	��M{p
�i��R6q��V����?�O�e�u�RY�{_M��-�8�!�K)c��Z���¶��v���oBT7�"���S8D^7t�ה�8�
����T{k�ͧ�87�V/s��y�-���r��]umuw�R�R��
������,���wLJ���}!U�8�ﾾ�ۻ�[c����m�v��o�K{ܝX�[�󝛐>�uEBbx ������ו�ag��Ov&L0�3쟦�ٽ.}�VOД>�T~2�@�Sɰ���Ntԇ~l�ƣB�٦wbz�TC���f�3Eg�|���%�Bn�P�s��9��
K�D�ʭ�]#{1�^��u	�
Z8�:}j�+`(����<��=��[�S&�>�v7�P֢`�k��kMG�~3���?"�K<��_{&����P����9��� _)Le\Wm��m&r����F����@n�ȉ�'�cto�e�H�F��SŞj&��q�:@�S-�2j�4�b��E��+!F�f�\r��07�T�"}TϘKl��"i���;�}xӳ�d�t��#rt����s&X+O�u.���k�tL�\�A�Qc�A�5��@���.��}�)[�u��cw�F��_;�GC��
�s�*�#�o�j9��ϻ	�Ч(��!��Ѳf���7�e򅸡�9L���L���of
-������h�9g}i�)R��G=;@O93g��~�0�7Ϫ�yn�2����yϠ��F�J�]I%�W��u����Rs�,Uj��%�옗�M���{�s�m)R�<�/��å��}H�?]���8�+��V���{@��wa���:�gR����;��j��ꆃ��L��$n��Kv^���t�!��x��3�ՋoWf��(�B��G���L��J�8��4	M�[N#9��U��E�Z��1S��-��tgl]L(��vS*_�k>̂+�Y�,��\�����O��(�3�J��3b�;���˞�ߐ�k��>��]�|������]���>1�;��q�cҙ�ˬ����GZd��D.�iݰ�My4[Or�E�r�؇��(��rx���;�]f9<���>�ݴ�h�J�ݨ���Q���G�����h��R�i%�L�D:\��p�;��z%]�hjޭ	�����<�e5ql��яU�6y�~d�̅������5�#%�)�b*���<w�����ݝ��3��G�?��9%��c������`��GKa�� &�ٿ���ڭ�g'����}s�;�;�}F�w��{M�{�2U�l�,�s�Z�9�οl�vpj���=Ʃe6�Ĵ�����J1�V��CH춁�Ƥ�z�ʈF��8�
��~F�;���M�.�I^Fd����8N��]Qp�.��Q���%�y��;>��1�����"�q�^�[���e���8�9��j$ۉO��H�����kKxC\����Iko6V�N��E;F� �\Y��:��8n����w���':���}*�����&�L��N6HP������hL����m�ФY4��t�����uVێ��j j�;޺���_:d]{�Oa�y�
�cR���Ͼ�(�}�YOI">�Y8�n�|��{d��fx���"�4�vC�'��@6b��a��kʟ�|Les�*��e]}ڬj�'�T���;늦&��������R>���>���b���F}Z�34�R}uљ0]��(f:�!D�Z\���H�"��4Ke��e�x1�ؘ8v��ǥA������팆��l��;������BS���7r��D�h�"��	.Ue�ļm�[Vɽ^����0�6-4��=V���T9j�c �W�d�4�V�����߹d�[��dm'4�֘	��o��r4
��;KﳀdnV
dq1��ԫ_};��D���;�F�Y�3��7���]��œ?���?D��e�/�Y6��;��8|Y{��m���>��������k��\�R�.{�q�6�Fzg6ͽ��7O5R��3��0%����?c�H�K>���"����*x�X����:dś��k:� ε�q�H�	ӫ�*�hyי��7'�#C����,<�x��J�/��t�u2��1�O+;I ΠrX���[�b�����C"�������'���y]q�V��Z���)nN��5O�v>�$בd�݅c��Rv�:d���n�2�ԣ�c�ֳ>[����Ϩhݐ���L�6�Ĳ��pXG�&}�!�a�p5ME�9?iޞ��6�k�] �[���q�Y��SQl̂R�5ys��>[�)�hj]mӉ�n�4�u�Z��2�K	y�+n�,��Z��VJfh��T�����r���"�U3�^ӛ7�A�S���#�f9����f�MS�i�����d������8��R��o\s,�n�Ӱ2ZrJ[��uR3[ςC�P�����HzoϯLq�2�O�.����NLƚ��_��~��ks�1%I���Qu۩)��M3�,W��U�����T����ǖ� �%;��\t����ٰ̃5_nKlWnYO�Y{1B�AK�2�䋠\�#hXw�q�O�9��>iD���fފ��ae��ꌴ1z�usCJ�/��v��}l/��&N�*�~RMx�t�Lk����4��V���XJoN�����1r��V��9i٩�)R�ш��7W'=���^�Q�_��"�wo�j�y�ۥB��<��^f��)�L޾x�4�=_��j]�����)i���I��K��ʬ >��:��'9l]�7��Xl����I���q��}s�r�kJ}bt=�ok7x�eB��Fk��
��v�A�7&�+WZ&�Ə)�҈������vV��>!��WM
��L\ah���
1���
{��[x�ɰS��b������i�5��5E�X����n�Ȇ��F��6ٟn?#)wH������'MD�,�1WpYD�Zu�	��J��eIdJs��{ˇ	�>��{F�1��8��B�����U�^-�ڗn��(zf�t�q��ǜ����?]9'�O��B�갤Tշ�W)�37]��Դ�Uēm+TKJ]�����|�`�h�gƀOaS��QvF���:�wLp�G/��<�ߪOљ<:����3��Q���O��2f�rשΚ��;~ﻰ�5S;w���_�~�s����/Ǯ����2���+$sGt�L����ղ	T�].d���������|y�?/�M�vXˌuYɹ��c�3�X�����(����B�7�V�vUn�_�bwky�]B���L�ro����=�5M<Y��:hm�v��;T3d��(��ɜ=�S�=Ej�[�ַe��ݒ��CZFD��A�7�޿�K5�4ӽ�"�s�o��MN���B(�m��@��	Y\t���c��B���-��������}�R{��}eI�)��{{�c��a卲�G����M��7I}��sS�m��
]��}V�����Qv��l�t]�t����;��u]v��cwSN�����clMT>���_G"Z|��-9����E�YRp��g�3�;D��Ӊ����v�sK�S����<7��ql�r:H�u�VR�Zo��M��3�m^J�M|0�1�G-�nt��ȹ��<!�NT�Mһ"#��l�A�B�B��nW�T͍n�1jz�=�/���wo�Η���?����P��LgQ�����-������ݜ�ڨ0t%c�WnbS�[m��W�!�#E�#�Ȳ�q7����>��Q;�iS:��U����w��_v���Vc���="z_��H �A�&6Sd�ӈ���ە�~]� �]�;�����H�6q�I��ϫ�Ah	�ƴ��ò8�H��Tx�aM�r EN�L^9���-r�ŶHJj�F�U�1I�p%TY�=ɟXǃ�a���&�|����C�۽gz��.�s�k
G2���������Q(�N�	�HD��b�L�Nu�gO���d�ݺ�z:�x��6H������eA�*��-99�t3-5	5N�νW:��R<�(B��������ìS�V�-e�!݃
���ӺK�os�K�[�H��=h�1�х�p3(�VV���V�4+k/i�ʮ뙄l}ڋ
55�Q�$�n�-���<*���Y؊�ڝ�2�J����R4|G�@���k;7,}~ͭ�w6X�2���%UC�{�]?3��R���c*�ib��9�3�Yw�I����^����?o�i��2tV���_�Ζ��uS��wJ�-��j*j��ǽu��w[��6`,�]Rh��ϖd9�7!���Vu�Ԟ,�±��4�~ն�t�0}�օ�k��$J��'R��r#�}�p#e���s�VT@�=���F���*�dn��1�%Й;e=�3Z�]r�%n��Q���N�2����(�&㧤��q�>W�fZ���{B�s��d
ɑ�N��W�`o|�t;�Oa�b~Ee����o*�M�����Ɋ������v(A�z@9�����i�i�Jn�~G_�-?I�$�Ǵ�f�Ϙb1С|���l;d�S��'$N���c�%��;늦&�������ͩ�����2��A�Z�]U�׽�B[��p�U�~P�5��8� �fȈP`�D���1�/o^H��V��*�Y�2q��r��b�dRvj���t~g[uԻ���"�<��U���bF
���X�Y�Z2�IՇ�Z��*;ݝ�SFH��*�]�GH�Y�j�����R�n��.��Ee�Z�k�^���/7sz��T���&�c.nS�t5�1�iu�)bV��:�RY���f�ZZӋ��׹V �(L�)��˰8�{r��?����]��x��\:��9��H��}�p�eM�R�p����{��̧6v��=�L��
����h��R0��{�@���*~c�� <�臹ck>��0d��o�&$��XXd8)�u�:9G3��7��f{y4���!��c
}�x�Y�NV�Rڪ�ͨ^ԒaN� ����x�k�P[c��˴{s��)�yKH�����rEJ����6�J���e��������O�g�{
��#��GdS�N`]�c�ٮ��u��L�r�ȸ�5���W�ҳ����'s��<2���13�s�Q��T]�
�6�̛�}�x�`l|��wg�Z�qCT�f��Z���󖉸�Q_}�b���V���Z9�V���WTٓ�*���/J���٫��;���L� WJ�O|q�+�y/�WT��|+C�zء�0�,�l��eg���U,�G1WY�i�<z9�19D�yd�;�n�����^���2{�)e��^T29m�x��T��4z�s�bvg�;��ľ�����n���7��	�Ђ��Wq�0�,�����L#��j�%�=���Q~`�O;��T�tr�<�T|<6�U����{ַ����i����`!�yG]��VS/7y"�V�ˡ�E�kB6I�
,�VSPU�
?�^]��G�O��҇9����s�4��m�NXg��Zv�����y��"�	��Xs��H���ۘ��|��f�T�>D�1�RІdoj\댩~�9�.�\�#jþ�q�O�9���J'�_��P�X;�����zI�[f�\��J��q)�������}_sUoM�q�
%Q��b��g;�i��7����}O)���(}pQ�������&̱��M�sY�,���P��VWU�)]�U/�L���fF�!q���c낋Ī+�}i��A3�A��Ǹ؍
�{�u>��m�f@k�* b1��;�t�W��6���Un�������o��k��t�����Z�t�9�~��'�eʒ.Ke0��]"f���F)��`�˷
F�d�d����4���b:y��9;�t�e*���&����j!�.
g	�9/ݱk%�c[¶�X�y��D��#��:yCE��m����B`�w�/��蛨|��T�%�*�"���"л�s�~§�[o�KBmN�%��穖M^=m��S�5~�ɕ���vK˶�"4�T�f#^�41g:�v�m3ҭ�]���B�#�[x�a}KM�(���dt\�n�R��9��!�ؽ�,Q"�,Z��Y�
��eu9p|R�w����*�`��X(N�eP嶩�"�����Dv�Un)wR��ؕ�dSpvfV����.���2*��{���;f`�+�/"��v��;w�T��v���.8.�n����]�άoD������ya���O�M�{�n���Xe�%��4�8�� ��8��sL`�aQ�ז1�C��Ss ���1�v�d�l�.�Ƶv�׀�����(
�5����ս:�w>���]��q�4\8�a��P�虑6(��X)�X1塂״�K�S��p�t�b�f��ٿXP1N�[��wS����oWU��,e�8��x���ݜ� #.���ёn$�N�7|(�֔��;	т�`/'1�x��[v=���$�p��Wt�c���6+h��<-�}X�<j�"�͎Q�Э�T�n'2>���oJǯ���Et�cXj5����
���к6��8U�|E��l�u:���c�k�ƌ�TD:@��}{4"�W#m�θ��f�Ep�Յ�&�p�=qDi}ɴQ7g�>��ф�UØ�N�hu�6�#RJfˠyK�\ ?�;�w����Ǻr*�Ķ��͇Q89e�p��u}�D��W��Ҹ��}��\;�����2Eu��]�5���jPu4��p��
Ɓ`,�Ȁ��𽴮[��q=����\�o
���}8V��suѥk4u�Q<��Ց����ޑ�Vl�������:t[��#L�$�y�,�z���E��/vV<�g�C�4����6ۭ!u_-9�2��c8�'_jK6�`�9*�:�����z1��8l���;����IU��6ب�l��6U��jWBȢ�D�:;��jԀ�9���lѺǓ��٫_=����
t��ٙ:@��+8�/�\5�+�&��ѧ#�bt�g7�&_���IS6�����pH��,2���C|�v��_!g!>�_k��{�x������82�<�M�өYUeɼ���6Gܫ�v���Vko��"[հ�u����e�u`��\�"�ъ��+z�kw2�E� Y�u�D�.�h:n�M���]e�r<����ҋ�s�9R=�LYC�`���Oyo�O��I�����Y��]��{or�&�I00iJ��e%K ݢ�N�&�t�)����ϝ��:˙�����c�A_vR�T�Ջ�ڻ�w]��mҬm+��d>�Z��s�}��.�'a��\ۮଔa����cZht�XnM��lF�f���� ���>��:��qq�JT�������2�- �Z)s�$�����;5�e��<�yN��M%���E>���P���*=�j�P���l�bp�U;Ǻ��ٜ��������X�oVo�f������'J�k:���+3�T��}�)�vt�em�c�b�|���b3ǼxUAfe����(����QErՅk):�E�!�@�� NEY9ېTNdQ��A:�Ĩd脒vb�ʪ�!�N�QS�9�n�AK�Q�w*EPj�6U:"l��NʯV��[X�]�"�hZ��F%C�9:�T�C���,�S�+�9�r7wԨvZ"��:Y3��eeE�g����+���I=
s�2$B��p�=0���;���s	֪8y8r
(��"���=��2��rrȭ:.������粨*�"�8����8D�E�W�㫍Ȥ�u� r��S�i.{���L*����tD�I	�y&�=�U:�:��t�wMGt9]��a�U�rīZYY��::�l�I����*�&��*$�G��F�IU�\��*�Aeqɻ��u��D^e����g9��^�8\�YPt��PQD�,�"�s�H�n��ؚg;���Nv݅�Z{r��XX�ֵF7(Xw�&���1I��؜�u�ҷ]f���b�M�Z�Ns���g'�2
X��(�Q����l$sra��k�ϯ���Y#���]�k�
<q�qԪdL�vA��";�2[g4[t2�c�j]�zN�/b>��r�oٲ��g5K������x�ܾQϾY�� �%[:2f���d��j�6d(��O�>��{�j�OvEd&�9ŭ>��ْ�,�0��ܬ�R�7{����jmc���݁��l񋅂wI��e��8Xy3�������k�#���Kqм��f���]|�i
�����)T�bڃ�L��%�I�q��h�uu<Vsή�;S�b�K,w�=^9T!P\��OaYδ� ��l�?������H�̼,<����@�c�l�kB�u��9�����i��O�&G#O�d!����Ƕ��ScOD��2��z�S�3;�K
�����z������|�P��J7��"���fӲ;��ț;�v*����Y��P������C,�* 	���)��Z%{%����BO�n�pT8�};�{~ΥvrR����c�P�3��5������BAt��1�`u�G�Q�xi����G�)��'A���J�O7$���N�w%��zjڸ�o��j��@�O4��y!}u��]"�M1�"Ѩ
�������pD�7���)�s�r��@>�|��o���5|U];pҟ[��B�/��¸Ԙ:ؖ�sV
>˒�iI,�����g�.�צ��e������w�fA�Pؔ@/�0a}�H����d�e��LO���Zd��TQ;��1̤%�Z�lJ4
��;K��}v@�(�|U�E���28����58�g��_*�7�)���tsy4cHKbQ�n�Y�X/,6 K�K3s�,Pj[qo�V�n�F	N��s����>���T[����*�V`r���g)2d%�̴��C7��J̉��̥�U�Jl�$�<NԂ�،�����-�E\&xqͅ�w_�H�UAHKш��p|�n�'�{w월>�uT�_-�����Q��e��I���������?\d�7�u�nNi�¾���~���_Xw_g�
�9���fʉh������,�s�nC��5�h�J0*�Z��?J����3]�#U����I���D�|�_�YhP��+E�`��q%��5�G5��1�����5W��҄�@��2I��Գ�T��,�Mi��
-�<�����h�}l���Sl�U�YK�'4b0a}~��(*�w��;���uA3�<�㱵+z��=�`U��K��1��6�����	 ��MO�K���)>��s.۪�S|)�{�5��Z�{3#dN�.l��_��y��Qۺ����_Wr2���Gi�I�A�����o�[ӫ3�3z�"��#��5FI��n>i��הs�TmF�m��ם-���Ҋ��b��C�}	�Vl�*����T�?��4���)��"y<7-9Ұ�A>��))}S��Q�r�;�v�� >�
����l�(���\U1C��v2Pl�����4���MSY�ڮ����>�R�ё�p�U��D�
��#+���6k�D�Q-������ɞЪ�^��$%e��̒څb�mj	tsH6�f����?T1�Y����$��>��RwuEo�
{�ܘ�
T��H���
�yi�_RG>���7�E_��E��4��s�DR���?]�Z�Y�>�+��^�SB�VB�D���g��IP��

�ls�*l �3����O��e��_�G~�O��`��z-QN{N����=� d�%�(�H4�`�roqea�3�-17-Q�?zw(p��$�3�Rk�0����:��!ׯ�q�ϧ����r�AHR��j�}���>�����&�����5�Y;F\�!�l�����69�����-��.���Y���}laz�u�'�Sf�n�jJ!�Ϋ�eA��h�����a�{��q���h �Zb^i�q����C�$,�^gt��9�@l}��lT�w�z� Ⴈ"��u�[�l�2;�L��[̥�PVWw� ��������K�ݽ�;��ͦ�w�Ց�ť��tq_�aY�<�@°�_j��ˮ���t�]Q�"�	f��8��U7K#�F;��\l�}h�u| ���b�k��V�;^{�̳���zh�٣G�����H}��&��ǅ(�2�}�W��Q��E\E���׽���]*Q<�qát�fVL2��n�ђ�u�,�m�~���p�1b�o%t���������R͔9B&=i�j�+;kb���K�wY�&~t��/!�oY'N��{j�(�g���?5ȍ�A�D��6�j2j�ͪ3*����b��#�l*|� %]1�-����R%����7=�b���og9�!��*�	�,UE҆�ve�9�5�.u��*�Fz'd\RRȍ�a�L9Xu����#b�j'�e�%,�K(�2Շ���iLֺ)��~Ӊ:kމ��8�d9�~�`��}����q�ś4�32/#��GQ�vH:z�@Zܣ�нBv�E��%*Ss�w$��X�-Nl�^u��LZ��wv�2'��� we����E�Uξ����38�i�J`SU����7k/]�K�%�] �_M�`���P���sai���=�}�!]9#�l��;4�Y���$}��/vUl����~5��Sy�fm5czw����w5N�����/z,A�wf�k ab�h>��t���VtLCtY�[�{]�;��É�ni∃7m�����
�h�u.�U�;�Y�8gT)
γA0��$�.��˻Ŋd�{�t���U똦�w�:L��aۉ���D]"f���B?KӧC<��]J�z��<��]5�����m��=P��y��6�J��G��:L9�;/0;&�;${1Z9Xn���J ��۶�����k�Q(��e�����X�o3��w�(��ȕ���/�Koi�7F�z�.�Uώp]�aS^����M)�Q�%�b���+ESc[�*1�0��}��7Z
.y;�uϋ�$j���W���Iy�d�FBUR���㦼�8r�T�g�l���ܵS�7(Rl�4R'L�m�!���S�ty�pг̱�}X����V��f�t�W}�7�{΋':~�&�?{�!����U����{�F�ki�E���lO)�05�#�az/:�q�.69����LU��8��+kdD�˓�Z�;��K��ʦ2�kK	؊�qM����
��p�����;�׎�d����e;���-�ܨ�|%#q%�=1�ֲ~��ئxoM��@ي��T�x��\��G#���ا��΅�/ʡ6ODε�%mH+kꝝ�.���m�ۻ:r�~8"�.����swiΡ��ir="�:)�}���ts�t��9[�����:��������d��1Y�W9�\6�������wX˥�����>��`/{���mwv�[p	\�a�����.�6^��
�=8�1r�J>���>ٹ��&���aL����J;�s�_�s�}�e��㳙��x�	�1�s�ܨjt+�GMq
�:}2�M���L���J-��>p�٩���Zd�|/�;�iR�Ο�����L&s�P��)�Bl2��m�P\�)��Z%{%��܇�B�_i3�cnTH;5�{պ��Zޤ�m���ȵ�)� �l �.wNõu��UٞY���e�W��mϯO}�ÿ��q�s(d}��.s~�5�}�W��H	c�vC��[�Ձģ1=Qy�&):�B�6�,����c���F�MAFģG[��`?����O�O|N�Ϥ�x9E�4u�ځF�,��ݙq�O3��@�t���do&�iKbQ�WC2�.� �)?�R�U�?�+�)�	��>͒�%�{l1כD*��d�/��P��Zk���r�$�l��N&x�]y��'�9������`l�(2��c~*nXW�Z�4���q�K����'�³����ed'�i5��dC�֮؇�>J�B�7e7���/I3�'���6�}~��Zk�]��Oēfz��ێ�ӕx\�sj�t�1Q���iW�}Xp�Dn��!��B��w44]���{Xpet=>j��|�%�d�:�YV�����a�9v�9lb�o96�]�6nu�ˡ�޻����
0�BZ3��p03����?�U�÷X������7�vۗ����
��e]*�3j��b��*%�W�Q��#�3�k�ǳ�^z�c,Fg՗�1]�>͚�k��#U�9����+�q�q��B�����k�t��)��������
���D�M:�7;�����j�_����~)9�������ǎO^/����0��T4}c�<l�i8� �U���q:�wm�>��7!���9�K����|G����;�vo/��̯�3��,W�"�(���%TL�=uL	�סּy)����/��+ZO�-����ܲU�^�t�i��Ca���&����������	���ϩ���Qx.-��nN]��z�e�l[;:ʘ�4��Q�h�a�tJ���׆��;dWU�}�WFOO}�5�U9�-�V��e�R$���R�hi����^�t�z�3\y)TQ�`l��n�DF3� ѺJ�4m�-ܢ.�yF�KG�}PR��62}M��(��E[�r/�~l�Q?/=s�/�ekP���/1H�vnFt�Q�F�=����g�wH����q�v�Y8̱�5�l�������ȼJ�}����ݑ�y��/JTtI������g-��bV�'�<cx���/���zwol�ò�Z]�o�.���̴�W0��"\1nF0j��C-�(J��zY10��˩+d�}rwaw)�ڭ�Ի���ϸ ���+�L�*I,r&WI2�w��wNy̽7���,�ʽ�Kʒ����M�C:�*��L9���S�,��ĳ�a�W�c��!��V��λ�-� R�q��{����	���Hˉ�]�뢡�KuA'[��6�¤<��Qvy�bS���N:��\N>v��R���1[	�r�'�F�K*���w�mX���7��ܗ�V�����}'�kr9�Iמ�ߞ�+�Oz����j����*SW�D?k�`�@	T�CJ�h���K���ߚ.�e6l�E�'|F͸Ro��O��,�G|�f��R��kO] ٍ����D��VOf��M?[/4����0�g�~�Y-f����AǞ������ _)D��4ͫ���mM��sw�J����?o�%p���⸫�ݶx��#t�lتC�ɭ.�g~�3��I�� w`<�)���qCr���j�r=��֚���#�YE�<JF�\�=uL=�cnP9�	4b��ٰ�{}[cݺs	���L�S[�6ԗB�B�#�vEג��5؛�_�>��،���(����{��!�T���|���ֶ��q&�P�b�Oc�
kq�'.	�@��N�e�
Y�/Ej�"ݎܗ�>�k��'ή�fPSoI�W��a�ZJ����5w�ig�]ʹ�f��	%��M��R/6�ae��~�>��:Lվ�z�q�|z�㜦ڳ��;��uˤ�)��._>�7��qg|Fb�����~�@	�?�~¾/sòA�Բ�7(�4-M�j��[�4%-/#�v�G�r�4 �Ȩ��tIngk�E�@�KG��Mdo��?RFL���~��.�k�%�2ĕ�������`�2�����j�T?#�Xmk�3�+MC!� ���:�C���x��'M$�g�ԪK@�~s�Ϝ�q10��De9�n�2��T67����6�n����h/�kR��N:p�V�'zt�Ͳ�,�Ή�a�a����
َU��>��qA��M���_��[�b��o���O�X�Q(�]������H���όLδf�x��W|9�`^Hdt�F9�.�aS]қ}�Z\/�ܳ� }�˻��<f�ȉ�>=sUT�[�5���'��t�s��ڌ���=\�4=����7#�����L�^�D;�N`3�}��]�Wh7s52�4g�5>wM�e���n�K�cϪߑ�o9x�W�}�Ɋ�3��[^�l��S�o��c-=�Y�����t(3����X�?#��up[��jVH���|4�8{71=c!����B�H���<�ϳ@®��݈�����H'1]y�U��n�Xq}���܎�[�b�[S�,�s��]���℠E��F崾U��f[�m��OCٟ)�]�lΔNY�>��{�j�Q�4�Χ���r���OUkw��#bo>��� mW)�3��1��fkdGeA�3i��ܗ��T�H�S�>[��|���kҲ'�*��߰ȸ�f�C�T��:D�+�Zr��%B���/ZD��3)B����.��%��k�UFq�κC	�V�.doi��"�u�üiP�'bm���Z^��{3<����XD)�RPJnj�סּ~�AT-w�/�q���ӛ��ZN>J��V����2�����}��2@���� O�����L�{V%�y����}<�(V	���4coj��
�5���GlǺ'�5rQ��#E������ܖ>g\���~��x\����X�����/��U����dwЩ3��5���ì�,���10�z�Q�@�_���^�.1�z�.y��:~��+B��_C�i��΍X����Y��c��>�z���>5x�j���f![�DI!�vFٯ�n�L�;�#�ɖC��uCw�U�� ����=�����cm����cm�c����l������6m���l�������6���6m��`�1��c���݃`���6m��o�0l�������6m����cm�6��`�1��`�1����
�2��γ�x	>��������>���������>�PT�BS�CmH��TIV�m�M�����mc)(�*��TP���mi�V�j%
Ei��9��iU�6�ڑ�jeL���5Fj�X�m���kUX�ͭ0Al$�Lm��͛2�kk"�ôu���񺽦�im�Y�5�����kV���ͣ,��e�� kZ��Ʌ�V�4�	13��[6�۹��e_9�lձ�a� =���*Zi2�R]�n�h;�!�Πژ�0�UT8���:4�
�%�+�����w� �p	��rU6�`4���s� Ҋ ��@@�X�R�(��s�(( + h P�LD	�M�L���ԥ �  쒐����hcCUM��� m�
�+�km�I��M�*��tR�'NR���W*Dѓ  x	׷-�Ҁ9�vʒ��m��wwHi��ѡ�m�Z\���U@u���5���a�����  �=�N�J�.]ιQ��������ܪ��q���������Wt�F�Q�v�B�;\��u�n���gc-J1V֒���Uc� ��)��j�*���C)��ꫭ+��軻Eъt���WW:SE:����ӌ��j�Q�:����]ij֨��liw  =�׎�&ڵ�P��ΣW@%fse��h�wc7tU:ˢ��4��+�Z�R����4 +ne[3k6f��Z��� 7W�%@��ٸ-J
�n������᫭]�wgNMmM�*����s�9v]w]��T�Sk�݅Y��ґ�P��o  =�oVܦk��N�v�*����ӵ�]erv�v�T+�-��7wn�ۊ7]ю�P�&3�rn"u�itZ�kJu�.�� 1�'�� ��6V��^�q�l�D����t��j��sD�� *��( @ ��&�R�10&�a40�ɠɈ��0�ESP      ��d%R�L 	�  &��"��h�I"a0&�4�#ɣ EM!�A�)�L���6��Q���jy��*
�A��6�S��4��4�oW���n��,c��S��T��[+�2�(��/M������5DS���ʍTT @���Q�
(�������6��~�L�P,"�A	P��$!!�I���#
VK�r�~��*���ʽ�𠐄�vN?�se��q<j��C�P���hР?c�ʇ�âg�/�MYw0aS(�X.�t]�~k��N�Uyv#�Tؙ��Z׎T�X�.�x���v��լ�f��u��n�6�lV䂵��6&�d\th[*���Nl����C"�l
2�d�-kH�z�YǶ@��Xq�V�wN�g��M�Ҫ�n�V�"�J�dܡC6�ٕ4�낵͛g�%�^^I��m!��z��`O�,�k>:5�[y�3u,�v�J��L��i���E�j �_A{���Cl�C�ndx��]�� ǒ%!�r��uV4�unh���hY��:�CMm�pU��a�j��$S$�Em�劌E/V醄�E[�g��u�����t�
kn֨X���Q���Eͳ5�Z�i�b�D0C	zUJ�Z[�j��*ڃ!�v.C����c6�G×0X����,{CF�J
�h��^a�V����Q��m�	�R��JT�`	z.�曭���^"�1)f�1f���z;A����R�࣎�F\��[��d}#2f蕸v��*i���n���qջ�6bVSVM��i�tn��p���Z
`6nj�nfb���B��zٌ=�%L�����U��Am$�:"��M;.-�S��P��a�SQ 3SZ�}��'��}Yt��XWG�Й%�Q5C<E7UM�3]���{[��CIkS��ѥ�i���b��1�ڼ��n��"��,�CF�"�1�(Q۹��xB���Rov�*�$�]�W>m��&�E�S:ʟ�4�w�N�k�%��̑��^��Y.A���L+�D����PQ;���5���І��B齺ukM�2��k9�����k쑙R���36���>3wjBjd��t ���/>��j�%`ܫ�l�-a�I�:j���E�n�u��o^-ŔC��-��פ:y���h����Leڊ�G&���f�*��ZT4��9��
��Kj���@f��n��3C��+]F�^��Л�8M�A�sF1D���y��,�^i�4:�Mh(����v���qneF�� ^!(���Q �F��i�tv�ա�͊�ҧb��Md�#����f�oCWJbY�E�r�A���ի���ek*�ݧCq�L����J�+R��:S/3p�z�����ו��b�G�t�[Ӑ�t!�o��QSQԄ<`�����T���@�؃r�\G� p^��]��'���B�1ܯ�\�_/����^�,U��RH�,��,5�e,8T�
�uZә��3j!A����7��k7wFKȊ,-RQ��昄۱t��{[��[R���b�z�6��yO2eኂ�ƙ�3>�b����װ�:`)���z��U͙qRW���x�V�h��%"R�o,[X�[��2�e��6$��x��E�{#n9SI�ȁ"�Al�M�R���"��^�jF�j�:+t��UM-�ah�6�̽��[�A������z�!XA�GfU�X��g"oc+h�kr�{��oSz�j�� kǙSD��,ܧ([��YQ]�3h@�ixˣ5
��m;5���s5�.�&��^�W��uk][w�2w��ۅC��f+��%U��+J��e�:�����<�i�N0���6�P��I� L�ͬ��f�won�^�w*��{Y����|J]�� YxQE�3v��n*A?�-�n���^�g)X�D�f7�Ħs"9."v�x�����]f0�,�[�-�5g��X]k�vK��2����*�@ϳ(f	���V[�ݦU0���ฃ���uk� �U>X+30�90��R���R6��,��ɪZ�˺�Y-�>��H7Mɦ]��ic�X�XǳV��>�	e��Qi*�{w�|��l����t�4 1���.���HT���Ǻ1JV�v^,�7e�u`Ĵ:��A̳��n���T,姰ۢ�r�$£/mE��6FiL��m����,��C�9�rֈ�՘�$k�'�Ʊ���@��D�U��_j9EY��n�m�m�oK�n'x�Kf��Z+�G�nDhe-�F�ۖ�|mCP'MR��g$5������P����,�#��݀�oZ)Qwb��B�c,+a�I���ڷ����TuPhW�8K�����aErڡ�5S��{��"��0ٺ6�j�
[�V6[�a����mi�J�+,�!����nM!���*�����5P��B�FF�F6�͖�%P��T�u��Е�ěZ��6��:!�1e��|�]:�J�Y�k�q�,��	{R��&��6�a�zCU�4�7-M�&f1p)l�Ս�B�W#ܽ^���K.ڌ۔�][{��;�)1r<{)��{z1��?c�K�w�E�t�ZL�]Dby��t�z!��^R"��ta�.ͫ�jV� �I6�{z�,Z�oN�=KM:J��!�u�P�A*4�MY�J�y+,n���[h��V�l�mk�5�Mf"έl��T�k4�Lڼ��Ie�3hH�� :��K(��r��z��f`
CSlTkZ���1�>��jY)��d��n��H�E��J,��Ow-�4���6f�P*y�L{ZoF����j(1u2��Ic0L��mާ[��9%މ��Z�V�3
�ը��Ij���;��I�l�t�o6ա#
��j���qf���:��OHO�sKQ�v���(ޖ,�[�v%Zc�yV{�*�=v�X�f�i�.�.bZ��A�ƾ������7-Aw&�r�#�Y���l�0�y����A8�)��oa6�V�l=�&�u��/�VE�������0b��r5lKm^�2���T��{0L�
�ѱFU�q��c�,�]�LO�N��鲡Eˍ�w�M�W���#�n��Sx�uJ�%�7�T
�!���wX�GoXi���ϱ&J�5R\�إfk�LS+��KL�u���{W{S#AF��,�[IZ ]�	�%=�J��㙢���쭁��[ҩ��a�r��-/�F���dn��2�0�t.�!b��[+P�A$ju��,���Õdԩ,&*P�a��ݼ���h�C,��L�(���Ș�Q��~�@��ڥ�L����i6���\��2�ll�	�)+��ov�8��s)Ig ��ɰ�iQȄ�5��c#&�y�/S�7��Y�)�O^݊�f�jU6m��,���1�S0�m�,���H�L��V���(�i�����A(Қs�l�i��=1���&2��ְ7B��4��ݡ����-[�T��O�hn�K]VʹFZ͢B1ԀLT�kԞ}wz��/M�,��'��-*�2"D�����Z'^Y��\qf�ű�4e�+!�n��t�iډ;3n���SV���F���X����Ӷ�Vi�S)��e��a���fڵP�S�ڷ�EQa{u{���T��Qܿ�ި�
�k�"�N�i�� �R�d�7SL�&�	�/L���Q]n!��Q�"�\�Kȣ�4LN�7F01�9��%�^��G(ku{R����"[o"�8Zx�ă�+F�B$Zr��cw�v�3`(��;GC����c���ù@�Z{M���ܷ�\��SW�C�(\��q�4��aEn@2�:��N+�e�8vjҺg0Y{t�Be�,%Un�{$W(wݱRE���0��fIK6�G��|F��ڪ@T�X���&`�[�N�IW$����r�t^-ۨ�֓���a���`(�����E�$�TQ{+-��!eE�j�@3���Ռ�^P&&n2b�I�.���-\���Ct��n`n���a�*�:�kJ	9x
H]����֭�ޗz���t���'&�M$��h/6���{v���N*�E!IHI�%Z��8f�t���$(6�v��g���[��2�Uɚ�����'�����7pn�6mem�% �M��z�n=��T�����й�nU�[̎I.��,^�{uk�ݦ��n-�.��u�U�gǮ��*��"�#pDK�CR�%�+�k:�af$�)��!{{(��n��P��Q �0�
�O��:*�kv���F�v�$�L8${�f'Z���-���j������`*A��#���`ԭ��g~�ǶX8*݌M���7�s�۲�:��B;i�NWe�,����@|��.���1'��i�l"hI�]��'�ߘ���dմ%��*K�]�Yyu� �d�4����[{u�%���f����d�y�A���;w�vu0�]�
b��#X�R��F��	XQ�e��XR�iqwz�SI�V����*���x�1.l�F����n��Y��P�M��^:F����65�F�VШ,��r`�Ѩ^�crI��A��ٯY��D���
;H��6�5��3�׺鐖"U��r��^,����"Z+͎���QD��ön�6]�-�S[��M�[��̪'6ʤ�&V0�^�?M���5��:)Փi��Fn����N����N�b�ӛ���Td%$�NPs�XQ�d�Uh����e�1���Hl�Y(/��%�ދ����KH;�t$�(�hְB-A)U����Mʚăa�]��T�*��a9�x�7.`
c�nJ7X�[���Y�MӗR�fV8�l���.^e�PJ�:�Ȍ]���K���g(��w��tLd�$��%v�k�uz���D�5�%,FĢ�ٸeW�[Y+@�cf�4���1���mr�m��)��xaDMіZ�6)��Y&�4 Ue:ssiH��w+�C7nBV�yD!�������I���k*��4F&��l�U�,�M��b�wc�M���XEr�;��hV"۬�l��HܶЎ]�T������y{�ȩ���GA�_2��S�e�$���/ŏr@��z�w)<͘��;�>����4�Uf4i���Ǫ��eX���n�Xc�fչ4\ɲ�5��,��U9[Z�P����Pt:�^/PyC+���|�C
H�z-��o��m1�Z���l��`vm�jh7���|���_u69����)�-j��EB�m�ջpՀ%�H��:$�?_�5�w;�q�z�������������G�t2%=_;T�ɫiCY��͢ok_(�oKZ���c�����ކ�*U2��v��������7Β�0�q��jkgolv������M*�����z��3VK�)=�I.�t9Jg��[=����+uw(�P|{FC������T�yޫ�v�ol�r�,���]h��R���&#�!�Q�<v�:�9�9������
���B=^\a[sѧ� V���'2���z	%2�\Z0$�l�C�]��_���5׆���]E;�K��U(��}���[��ˮ��ގbIl�1��л�����N;W�g+�5���?�`��;I��}uk�ړTb�3O���K}#�r�^�:�ep٠a��(�w|�Vi��:�
n�Y���iخ�=��� �J�v��|i�� W��Ln�9�����\
vnX�-���Rޖ	���dfڗt*܋sFes�t#�!.⮫���֞��5��iqCB��J㛉�!6�
��� ��j\MPC�)�@jx~E��ٖ�໓��F��y�;�{�6�,0�s-.����f�CK�����:!̶��Wv��g�L��V��]���ilӹʬ��d�����\�H���ȯwu.���N��s'�gn�
-��n\;8���2O��n���/��\[���>moLXy;�Ԏgka-�$M�wp�%�Ƣ��\;/�,#zkh<�o��yF���ӫ�1��K�U���(6����۲�]"l�O����Bjz#�� ��f�j�\�B�J������w-�; W	����*����d�rnӎ������
F^���jeZ�)ӑw��%X��=dd����B*E��޶�}B�C/][�r��s��(,����s�I�kN����]H`�r�j���5�l�L��b!�hT�L<J�FD��b���F�)�uo�4�������3B[�;n067�h�>��isy%WO	�w'VkI� j�{��b=�,�%�J5��'��M	�zQ��N���W��\��y1�m<K����ڃ&؄����i=��f��*��G�x�^wn�`y%3ޱp|*YӋ\�|�Tb�S�\��^��q��l�c����Z��PQn�7 ۝]�V�u�h�S��7N�r���å�켩{D��ʸC,5�U�`q��xp�L�u�o��2"$-�YlnԻ��E��F�]�.>��%�n9(�V���6��4r="��m7�#����e�]�F&a#J��R��{c�{N�*�l����c5��v��f�
���&���ix�Z�Ҩ���t^*
�a;���5��x5Y��>�S�^\G6�.�H�ۣd��b�PԖ:��EK�z4�^�ܑ���e� 
ul��^��-v�v��a)�uwŉv_p
o"�(�#�7wF:�SR�u�����(jR-g[a��l�I��Gi�7�W.��	�xG��<L�_^]ЫJ�	G�|$�����kf��mT%ֵ��f!���p+7�z˗@�ma�I�����J˱(7�Ȧ��c �ŲJh�pvǑ�rbbS�7�&�On��0FevX���N��K�4f�)�N�@�%W���j��eR������d��GFSr݇Ժ�$V��:\�mq��#p��%]o,�4G��7.�N�l��- Lx��xL��4ZU���|�����C3��飡��Q�ɭR`���v��Ц�3Z܌<�1\}�GʫY/w��[�_Wu�Oi�ѸEs�9��/M8�-,��
��Lz�*��-52�K:��V��-�N��:�hw�7��NY����;K{�[�ޚzt�SreZ�`����D�x9�\��a��6-d�S��&��8E�y���̳��|�Y���nH�5iÚ�O&-�d�AO��	�kR�2�<5}G��@3�{�݆9|/^]f�Zv���>����|Xnn%$9g�UFv_uu�z��G���v��P����J}�gkM��{;j�4��=Ip��4��4�	oוǳ%��$"�Y�r[��V��:��_9�Nۍ9�+\ @��5�YKt���3v�t�P��M.���ލB��=�%i��#*�6h����}��'"�lY(r�;�&�;^���5ȓ�h���S*�c�c]��mj�Z챵�T"�Cޣsk-B��.�:#k�LO֬1����n���ˑi2	BkLY��l��fia#ڝE�a*�!���rI58e�>RKHN`EN�Zg:��]�7����k��3�W�e^�D�v�-��R�;]�^�^�b�"�2�r��D�M"�r�����R�1ؼ�S�-��;]���N_R��6�f���dmn���E��L��q*�m�d���y���]�V�萠$c��}�y���v��-h��B��-R���7�:1��
�`r�&+j˕��O�e��;q�.�C�oW]���L�1ڽ��k�t-�x��ϙV��y�E��`2=��Xg(&58�t--�2L.r��9��镜�������@���D�m��y�^pu2�z�
3]g\Uy\J���.�8gSc~Atlgs
�Y�mf�{���
�k*�(ES��i[�z��U����p��Ž���z]�}(�_'�f=%�v�� �.*\J�qn��Vˢ�v;��	�|��d����>f�m��*w-�Gkr�8�tܡa|���Z1Aøj`�#��y�٣�}PZ͠���v���r��l,q�X�
&���0�Ww*�h��A��,��`�ڼ� ���;@*�N�ˬ��p�q��R�YF��F;/�c]��8S��k�L����-}׺�d�5�+`��GP� �58[\�-_}i=O�����	��&"�W�.S9��_]��e�r�"�v�x��AqȎ���D�%��V ����}���%��q�&ȧ|$;Mڒ���1���sv\U����Y@���R�ۏ�F�� ��N�?�z|� �0hCF��=��GZ����C�b�<�p�v5\�qdj%[�ۖ�`�M����aKJ>G��5��S��7q,�L��N��gH�:��} ����gc[�!+�}��]t݆��1qޜ`����D:��!Q R�]�$6]:�YJ5�����p�l�˽ka���f`y���v[�w���MސF����8]�-�X#����A�AGg*�ii���;���k��#UAJ=���	�h\k���H��E�Ȯ��c��uc:(Q@�$��g��{t�r���ky�M��aw��;���\+%uO$:%`�E�� G���t�o3XT�W[�`���-w�[;���@Hl�u7d�Z�ipaY7�>����y�_-��ڎ�p�(�V�N4����.��V4g+��ih�]B)��_b%H�LWF��b�P��l�m��&q*��d��ƵR�ա}��C�a�W����_��i=��󮵊x_9�kHwr����t���ZU&7_-[u��Ԏ�@\{��/jl$,��	��l^v������2��tȄ�^'\N�Ql����a��Z���[̵�1H���]V��v��f���˳��&�e\9�9��!
�`�ȝ���Q^�����Nt'o�����l����gj�X��}̷o�y��"P�1>;5A���㴞��`P�duδA�救�4�nK�*�V�:aB����6��s�!<#�7�^��ke�1#C���Q�����ǆXJ���vd�ۺ�Xd�%�t�q���3�ou�QK��&j�wV�u�jۊ��}!xb^+k+03�~~�Op��8�ά��2dR#Y���pm;<�e�`뎂�it<8��x^���E�-��G9��y�N�vurE3a������U�v�F�ٯ-��n�a�
2���;f�m�\�f���ֱ2k���;L.��a;}�U�G\ [T���t�:����O}��)n�/4ʴ8���ϳ����.M�"w��:�-Re�J�K�,�K��-z�x;w�0.C�y���7+*�X�-:��4�f]!Bg4�w2wKb>��e�N���b�m���G}�¶л�|ʢ�u��:�7"���"8[�x�^��7!:���v�Z��]�gq˥A�W6�<N��-��$y�Ep��:�V�]vc�65cB\Si�ӕ��d�������_1�v��1�I��V����#�{4�WFI��+],��]�YY���\�+���Ó���d��]���M���\q��jqX�����FJ	V��9`���m�����+���9]�,W�E�L�*fZ�9�b�O6u�_=��u�,8��dA��eg���ZΜ��c�B�ZN�r���j�m�]��oGRsUۄ��b�qJ��L����a<�%{���0�,sxb�Ko������'*�M���M<�YE���*T�5���;i��Q�{b�m'���0�����B���z+���L��!�eN!&�"/���brd�#&'�5m8�{���v]ltB�Z0`S}B�b����|v�x�5�݈�e<�%��S��Z����^'h݁�aΠ:+��l��"q�9-�qz��F��1ұ�țC(j�Ǜh�Nd����{��$F�ɜ�9ܭ�{�.7�1�{�GҖ���-�eq������r��ߏ`�۬;a+�����O`�WӀ�r֚�Np�rog�cE2�����W�+����J���.V�V���3�W�����ZS,����N��۽��[�r��l�e7(9�S�e��|�x틨��S�ww�+,�C��W�fh���pqdnԁ��8�����v�!`�ni���@ǳ���]���r�T.&�@-8�t��l?���
���H�I���̈́�a�'Z�ݎ�\��b�M����xu��+0`�xo^7+{�H�9b�.�V���S�$���حr>�B�{���̦yQU`���ڒ!�;�m<,�+�t2fo�8�C���gpHP롶�խ�F�1�n	,W �b����]y����e��j��۵�����`P��U������u���^KK���x����]�*�<7k����<��y�ǩn޻�t��µ�;A~Q���hw�DU�o����>�ާ�eYC@���#<b"l\�b/b,T����;�e�M)$�� TDE4Ԑgzo�
�)��@P�=NuDDE:�͛t5l�U��pS,Z���t�a?��+}X���f��T��u�Bn���r�5�Q��镩fTc�!7��6�zbg�[�:����o�9�ۗ�twf�	WDJkvC�f^�OL8-��xzPC�V8��k6��ܫEb؛�n*��]��,��<	a˧��,�_K�y���/:��h�[qdۓf_@y���a��e$ՅVk��ô̥/u��j��Q���T�*�*�ۋr6���,�����-�u2�8�x�c\Ӿ��B�"��u(>[�[!��j��Ib��r�"�܊>7W��"v(��x����d_,
�9+(.;�c=%��I��[��������o���2�q+`�=��\�r�e�
��ABYT�7:�'96�A�bRa���1
�iQ�p�2�N��8o�ܬ��b��cy���H# U�b�74�Pɛ�k�]t.|9Q��J��3��������SF���51��G�n�?�`TgX�[�m��}�g -�Ix1Ύ�IvmuX��4qul�6@��`��I�V�d}lsE��X��}m�T���XY�����́�.iw�Z��NtQ�_c9��r�-��a�]��շH^e恳��]��ו`]��2��a�t{A"���:sb}����57α鷜�n�b&+�Y)Jev�!�u���ݤͨ40���I�MS���Ւ�\E��PTl�������2������3�z���,���ҷiAh��z�Y�[�S�K��]p&���ᛪ<2L�q�Ie=G��9:��%ɮ���_]��Y��-o(Ѧ����UgZuU�ض� p5��L�*)D�K�[�Y����o�s�V�6�c���9�������=��\���Yt�	33-�v���T��u
���J��� �3Q=W/e�.N��HQR��l�u�����h����͔������J�`��od���:��oL���6���&��d���~��y)�)��Go��S�V�Z2����l��P�p��%7�%��[�c��kv�Ău�����1_'F[�P}�o>8n͊3n��y�L�hM@�Ի��]v��;��\�	��\�gOC�/X bՋ
,[�x�S�(�B��p�ޏ(�1@�����������x9_�u�n }S5:�Լ�[�1�S���1�H���,�U�۴iK��lJ���$�a���:�Cv����m�(n���3>�M�Qǰ�x�Q�ǉ���:��3un���&���vkw����&��CR��v%���y�ٖ��
���h�^I�L�z�`�E�uϣ�kysV��*��6Ț"YX嚿�a���N������;���n�����3��BU+���{G�f#\�2�ӄ9A���a�@;��F��I���[@�Y�e6�/_s��õ���ӡ�:��s|�Q���Z7�W��X���C!��n�����.�n�<)�Sq=�ju�ۡE��Ѵc��DV*1�:����{Ҥ7yw�ٴ��eh�YБr�b�}�*z��{���Al3�¨,[O���Nس������M���v�u��4�"�Rnv['+C^Ô�t��{Ϟ@m#���ۃ�֑�v���n@�]T��-�5;�N�5պ��L�$g������ N�eK}3R�b�e�����%�/�0 �I�|l�	ŉ۳�d3O{�u��_sN�P�������Y�m�Xy,�������?��A�N�����|2�ں*�%��RA[�5.���132���8+�EK�A*�qr���-7���Tu��2i<;��QZ�X�,���e�5�a\����9���us��ѭ�MԾ�o��;56>z�p�7^_M�<��C�5�C٪�]1�[�œk�w�܂̈fZ5>Ԡ�.�v�]���9�2���l�Q^�)�2�:қ�-�n'��ZGzVl'+f`�9��n��r<nӔe��ǅ�#��؉��ӵ{YK�vV�"�t�����,�iz�"��"��ԼS���B��)�%�o]f�ا@ݍ�"��Yz���J�����6s��>=�2q���vTȏ
/��E�iZ�gKU�"��4�*���-�a�Z/�K,�U 7{8
[r�*�g�K������AZ�Ya�\�Ŗ/�v�,n���		�P�9\�6P�AԬ,�T�z*ձ���')0���m��d\�u^^1]����b����N�Q��!��`�Ltk��8�.8)VJc���sK�ΥAd'X2S��[.���R1>͈�E�hW�,	�l��]��CE�6�αY��T��j�.�&�`w����+6p�,ٹ\`���IVZ�G.��`�58�V:v���*��h�{k;�c�2�U}ԣ-��Z\�X0v�w\�n�کBgI8�k��.U-�o����be;ゑrb��|j���u��kn�E��1@��1x��z$�Xʹ��`٥r@����I���.�<�X��Y�+z���ۮKK�E�6��U�r�#��ܳ�G�qu��۱���6���=�T���mv��tDRى:��:�ఀ&M�GE�@�ݗs(䎶����3�h�/���|B;����6��@qa��Vn�Ϯ�u��������6o�\���JsᑴX0$̓�����4�	*��AD����������wI�t:e,�4k,���m5n�+5����o�����(M�Bry�^���H�m*�C���;4��q}��+�"��nt$��M�Z�����b&IN47���On��f��')2ћj`�vl=�w5��B��2ڗ��0��&ԥ�z'zX4��fsJ��ڻب$o��rr�T:V(��}�K%M���`�u^�x��.#c��Mm�;˷3h�-5\{�f1ږ�6�v�ly}��&�������Wv�il¶��X(����N�+Z�zXy@0
�վ��o�ǫ10l%I��9�D ��1ܚ�].:�s���#�҅e��/O#%w+����eElZ 3���|E���8?I}h��n;�F����wC�N�G�Ҧ(� ��q�W�������m��Ƕz�Z`�b�lyX����%�����9}�3;[}�!Q��]���ޕx���;.P/����j�6B�`��_;��S�/�3�0t��@��,ȣc��&�9̴WbZ�ӨOc���w�:������6��Q�S,�R�2ܶ����;�Y��Yr�r�`���`��I���G�v��Uft��桎[f�8�n-Ǵ��]��-��x��N"�Z	wCXw&����k�7�p�n�m�'>9�9�#!�Z�4�qJ4U���l]��{e�|u�[@՗53�-t.��W��Ơ��zb�eɖ�W��ł�TKc�ޒ�o`�{��3�6�+N�!i�����G\�W5� �X��n5�ha����q�˳�Pd��qQF�Z�Ml*VK���K�lY$2��O[���X!�`]���]aM(�ՈNO�c4�r�гN�J��Ū��R*��GcJgr�N!wvəi�BU����]@9�L\�u�[�^�e�ݭ���v����N���Č��:k�;���)��@=�.�Lt�͙Q7˻2��`�*�Y�X�4�}dLw��_^R��_J������]�q'�S�N�Wb�U��^e%���jޓ��V�M�ڂVܖ��>v�,�B����К�P�3dJ�M�<��∻bX=K��- ��t�! �e��vA�v=��6&�{�z�ָ:Y����e::�?v����C[*���[]Gu��k�i�2ݦ�)&%�t��&�|�7}��V��9�yf:��]q��޶��^�Jl;r����T��v"iu�.�m��^mK���=��;*�9&0��2��!�R���Թ�[��)�J�}��QZ�ڎ�`���B��3{/e&����]b�o���Q
��Hf�]ܘ�N*�]8G��[����e:m�*��.� �(��&�k�T��.��3��AQ�m�+m5����3Bp��GA��+�'P�� 'XڍJ�k�S���z/%�����f����i
�і{6�'���;�u�Z
(LQU�ʷu�*է��1��c���ڠ-0��c��$=t �zN��3%7ll��zN�ֻ��]Du�w�8���G��2ř��y���%)�Z���UL���]�[Sͅ[�p}�[����V��]c*��^�;�����;��[��bp�w]#ԬKԤ��v�ޣx_h�6���V���Ĝ�ȓ�\*\b��|w��ZY6�AF�����EUͰ]�ʓs*�v����!�l^n���i���-�A�D��\�4���SY���Z�3(3V�������R�X췷m�$�O%�o��l���.�9Xf��9J AG('�����Ʃ���yB��2v�'O3���n3C퇍Xe 4;��*kr�]ܤQ��T<̭����h����!���v���蒵��6u�ge�����^6��ebvN�ܺ�W��7�$l��FO��Iό�S�f[=p�����L��.��Zf�XG�W[�D�QY}&5�M���������`ő���W��a��7���z0r����;O���(�5����z�
2�w0`N�1�c�YXƼY��mN�F
ouf�hR�D�=J��v�c˻�s.�⑸�m������j��������m�>O|i�v3xt �q��-5�H��T*oӉ-�/@ë^̫t��orYC��,�ue,�R�D��*
�Ԩ�d단�Pк�^0��9J�wE89R�����B��N������ʐ�;�VBУ�9����Ph$iT�y��R�S{���;5c�st� �I�IW�������t�J��[�3Bќ��e�����V�xj�&�5A�m7	7�����e��0�b�n��V�'sT�%fYAP�k]&5w6�����W��b�ܕFS�ap�h�c���z%˙�<�7CA.�w�sV��V %VB8ֱ[�]H�ڼ}��zm��<����UӃO	�1�41^ٴ7/�����m�O�ټxڢK��M���;{��AA��v��o�^<���ߜ~��?�L�BAR/��>�~~1=��!�־���?�x���~�0��U�Dk�� �O|�CYw{�R�Q.4�;���n�i�)ژU*%���7&eX���-�mU��8\������x�w>�,��u�fn��5�C\�kv���k�3S��gnV�sP��;�g�4��te�9#�y�]s�O���2r�+2v����4�S���u�\�z��B�
�b���z�r��v�A�=�i"�%	먬8�������Ivll��=�7 Ա����sh����[����9h��F���^
RV�3$�f7.f��=�D�AC:3\�
���$�.��;G�
�0.\�2�AX�goV���l]�Ik*df�}i�"�� *q��g&�jU��d���M�g��#����ھ=hqx&��ஶ�M�F���iN��!B�Yܑu2�mV%RFn7������^����u5#[��u�B�8���Dzn�̨����%e.����Z���u��Bso�SDw$'z��}�%�|+y���w���С͞��Z*�s��o'(�{�J���ݵ�Qs�\5e����=�v�.�,�s�E�����9��Vl�~W���F(f�\�"�ER���+Y�36��R����-E"�P\�PP�̨��
�*cR�q�^,����-�k�:��.�%eL��Z�&Z��GYZ��F�D�*f�V«��Q�UU�[j0����EU��-��2��I�X)(
��Щښ��YR��3+P����֣Z�*��(�"ֱlR(ZYY\ʶ�#!jJ�V����f]F��[h������[-��QPY-6
�EQU`���5�ń4	�?Q�����׎��{��g�ߓ�z�7\s��nn�VoV�H_Hv��qgk��w�D��p4���)����O�o�����H���|���w��;��]���y��q�;�������Z��&l?�j�q�C]�T`x��dr���K�u���Js�:�ڧC9�A�E�]vtc	���lg[��J�����嵗����¹�/
�����1�,�4쪿]�M�I�<3̙6į��3�����y�u	:�RՁ7ʑ��>a���e���k2;��lo	��}��d��#6��ȍU۫1�
c�����sJt�a��#ɮ�L��5u���<��L��M��)��aR��B�{�Y9f���O�y/�㹻��T�q��2��%$O�Y�K���;/#<�YSkr�-k
��d�5�:�+��M@�/z���c�uN-�7�2�!��{����y&&���I�
+�5nWi��w�7�?^C/k@S�#Z�ϼ�S}�O�^�����ƿU�����긇c�[/�LpO=���y1F��n�S���6����W���k�C�vի�i4�6f�9=E�ڢݮh�_h�����ׯ.q��5�y�5�/fы>���������l���Η�~���G�}��'��mf}9��ʗ���'��O���rBjk��6f��[p�
,���[�I06���A�.�e*8���w��q��v�SS햆6�X�)
�j�=~s.���xvD;�3$�˲�r	2o�6�P�z�����:f�ջ�0����vl�}��XZ�O�C�/��i�8;6�[�8Gfb�%5%8]�E#��˘�FC�����`�u�mlR��bn��WI�p�*<�u�r5u�B��*�!7���J�����ݺ��X��ʘ��I�n��ޓ��Z��Yn�fQ�������֢�i޴�W��Si��Qo)mŹ�'����d�4���2����ld�c��|P��f�yy�`��ݰu��ܧ61��캝d���r�+]z�����xK�¶�v�	�z������~�"��yf}��S���Ac7Ev:ѝ��c����¶7�2.�F����vKs�N��!��R���(R=h\��uw���n}�-q�lV5<�M8[V$f�	�Zj������j�o��k�?s#K����\�Oo�{����1]�/�����������܍�P�Ix�����.s�]�-O�m��+��f8~�������7q��(Vj�l)IM���P��:���es�$YM9Y��R\��GT�??�����x��"�з)�$;W�����JjR�66W��MW>�I����n�T�~�w�P��"v)n:S��V��g��և{���fD���t�<�))��VjzJTǟq��	N��ϨFv��h��kKiE�.����bm��h�g���yZx�u�y����+5� �w;n���:���5~�qu��l-e��	���o��-�E��)����T�<ʶl�t����ݻ���j�Ø�9�N`��;B���9��y���7���@=����*��_Vt��{�JԌ�3b*��N����5WIʳ�Cxj�f¨�m�6�Z�����]�3I�Zjggw�{�`9v��LhJ޺+/e��
�6��Ѫ����!�0�Cj9ZfI�< �J*Q�/��e�zz���Q����S��ӻ�x��R��K�([��R;./p�^��UH]oy�����r��zj�dYMKW��Ƭ�Vw{��Kr�ߗV֞�o���y-g� �by���%5��엳ߒM�_44`=��l�=�M'��IM��y�[���G�������g��ܿ����j{��Pz�,���p9�,� ��^ ݈�OzKʝ��CK᝸��&�,1u��;�,1b���Χ��؂�����f�vpx��HU=gb�:�jt�EC8\h�nbPB���܍^ʈ�[Us�C���C$|�V�dG~ӳC3q�)�Q���{1��^��&s��ъڬ��b���颔�rh��X�7��<��x��B&��zv �\�ݣY�:���������^���I�P`j!����D*u�Y�����u�d�Sc��ɏ���C�����Y�F���B���{�/���?k���f7�?e��*���ԪMI��ˋ=��Qy/�ʮ~�g{ҋ�1���_ܶ��9��o��O�;�M�/�z+w�mؓ�1��ǧ�MŰȮ����;�ϟ<�*S���=U�l��2^�҇���X�R�y6��{}�����}��j�f���5_���$'cO^�;�dgx�HZ�#ˣB�t�7g�w;�d<��~Z�&x�����=��g����l��:�tO�`�����Jҭ��ޡʆ7m��B:�g�|O�{��Li{�y�8p�bE�hS�`��[Q��އ�j��
��N̙ճl���S�����p9��b��� ]��[Z`�����6vT��-F��k��L��Laut{A8U�꾠{"�ӛ*��s��%���(a��Y��l=��%�;o�\�j��h��-�[��>-���R�>�6�+�i
[�2�ק�Q�+����g�Р�+5X�e�w��*E�<��c;@��r��Bq�_1^�jk���U~{��s���_ӝ�&��l$]�Z]���MM���1_I�xP�ivGFP��^�Ts�´_�ӣx�3톞k��a�\|P߳)t��K��rJg�q�ϣ5�����2`�k�[Y��d��N�{vc�v};Ƽt����[���=�0�w�-�Űyt8$��qܵ�������AW�Xy�Vh98��ͬ�۴�.���|�ošt�ӽ��WW33��7�wK(�K��z?OT��w!�=(�j�HG1�$����Km��f�)f?E2�{*2��2oe:�n��|��qI'��]*U�����ڦF������,�]d̛�.-��>�PY*�udš������jw#V�=��J����W:�����m0*���g����5v���a�m{�~����P��t��t:T��3�vW_Q}�N(n�����xx�Տ.��i��M�\� ���]������{cg_Ks�1S�t)�x��p��Cۻwy�zwq.2�2����6X�'��J���}���i�vf�nv�����#����m`��k�ob�����Om�*�8��]�J_��{�ە����.:��
�4�-z�a�d�J��l���f�z�AL/~�,���-�}x(l��1�Ca����K٫��A��Q�1�L�9�	cO�<H7zs\Á�F'	��Y�[8m���95{����y'L�|)�ziav;����P����t��蕖|�{����̗�B��Ȋ�+�DiKu��<����rs���̜���~����J���^���)��t�h� �S>�(|�pyM�ϟ�ɓͦN��̙�7�&߷*�A�lb�6wt�{���G����ڽ��?5�ި&z�e����.�F�ɓ9v���RO'��ƀ�U�&�+�d:(����Exѱ����Q��y��@"�g>�����,�g��%"D��eC���&����ۖ�����Sv�>�*Q��ρ|o��3�O���'6c����]_��]��&l?�f��Aoee��.���ʓ%�H.��P����+���TV���m��n�Ԯ���&�a?L��&�m�ɰ-�>�܍:��T�|2Q�NL��P��ˊ8�ay
=�v�bF�$�0��[~�j���!�v�s7�9u�����R�=��KO��<:��,�J�e׊�~7I�"T��#�(ԅy�ϭ��z���7�W�����uس�/�����MG�خ�Bc��D+�ky��$��l��NUq��*_�	C�G�e������;�@��e��M��\��y]�C�C�М�R�������3��<�[���yn�\/2<�Ԫr(���p8u��^>i�u4m-�׿*�B���/�=ɮ�- 둻���8%�6�A���gշru�b��{揂�r���3�����gJ��o�{XuXhu�q/}J��W�~�����X��3�����~٘6�E�>/i� ×�a�k�{�j�'��}���<��/;��lnJ�V���%d�脟k�V�g�Iˤ��W\� m��z�� ͗�Hlڹ�
�@v�f^�Xn���Lnr�H�\dw6���N�J�Ȁ�Ӡ��|������<�U�������m���F�����3�T�N�N_���̶:�E���-��$-�q���]��M�*ƀ��`�F�w��k\��N��8�v�#Eѥ@��ڏ1���	����ɏ� �\��jڥH��MQ��gV�z�7��ٺ^�����Q��8k�+��u������E�X�c%���jv�ҕ�oqCa��N�bYVUgEO��@|��*��wS���dV�.<V�܌��`��j��K����v��7e����Yu���ݎE�����U�۽p�;,Q�+9������Ul��0e;8O,]Z��6l[ou΁L�PubW��F��;b�8�ݞ����1l<%���� v��J�s59W9>���fK困~T�>�&��&��k�N�r!�2�d�n�)�B�;���'~����s�6,{�t?�/�ePN�;6Ŝq�'%Q����d&�Ǒ�p�_a���(� �J�ѻV1�>����ƾ ��/�eԀg[��Y�IIE$�)��ie6լ�N���ZO��H�w�VD*PVR>;M���?	���R�.HA!��b�Q��^�!.��VV����h�]�d�;����-\���Y�mZ���n�Co	��U�[ <:�X{#��'u�-�v�:��6��f��ڊ[��*��E5����t�u�B�]�8k"�Bf�  �b &�R�tWڥn.yt��:�mĨ޾�C.�P!͍U�F[�2�zy֨��p�����lw:�
�I�8���Ud*���P�S*��]}�e��� [5���[n��F:�F���b�滵�1�`f����^���%�Еn�F�|�(�(J�tF��/fYe�|��A&�{��&m����I+��D����Z�v���M"���C=�f��Ey`^40A��O0
=x�5nh����ɧ��P~��h'n�k}���?T�	$�Oߒ�ȥ��"�-J-mj�݊�U�b��b䨠��͈֊�k��֍Mj&A�֤DԮl3\˶+0��ZX�b�XԮE��յV��ж��.�#+m
������$B҆�
*�"���KZ�Pֲfd�q��]�(Ҵ;6��*k���t�X�j;k3pd26�mAA�U�m�f��[ij�U��S����#R�j2�J�T͎��l����jYb�6����m�)*�Z�j��2�U\--([��5Mm�k���-�a2Y�ҥm-P�em�V�h�T���[��\�r���Z�����.�EKi�m-e"l쥹3D���F�*e�*",G7�%�U�mԦXͶ��SS�]�1U����ϼ��~1!z��]��1ek�x>Sń�ݷo�)g��N�o�-;�9Mn�\��_4{n�(9�F�1�1�C/�ޫ�ig����l�1����=ֵ�	"��E��¼��Sf�'�y�rf�}3TƮ6Go���/ʲG�یv���k���c�G��>��{��~���k��:|h[�-��CW�P3�sFu�5S����X�nur�h>�o��N>F����<��e�WS��u�=i��foR\�.t�/�ذ�� �pD����ٴ����:�[��Tp�aR
�t�������K^���Ձ�ZLZb�L��b���Ӿ�V^�k�Q�>+��M��]��
�v��7�'�&�y.�I6�'�MOZ�����H__y��_��z�U��g��@07�����G�B��ܾߵ�
��~�ڦ�"?>s�`�=M�����^�<F�����LmV���i�˩3��̽���'�O����|��y�,�އ�Ӯ���vE�xխUӺ�}W�7ķ���vQ�2\Wq�oO�ٟxJ�v�n�>��M�:T~܎U�GԽ�ϧ����Ζ�U�B�z��jqde�oE�*�}�#=h��4�-�&�$���OW��罞IN��A�b�K�-���)��/,������8݃��W䇓�(�P�/��s�=�CW�왪XԪ_+�������i���]�L�nz�5�߂`x9\1��?��=Ig2�!�}Ѕ=�ۅ��{�]R���Y������Z�,Nf����{�r�^���0y��F7�NÙ���̾�f��9�v6���ӵ(]c��XGN��5�+ʺ������DYە�d<wW��ae������8��	�*:�)҃B&�.le��朓5��O+yoVK��Oy�а-{nPѾ��׏�I'�2��n��a�V6W�x�Ԩ�/����P��>�G���01{�A�Y�V'���!ƭ��<�\Q��<����A�WCy�;n�ǛHul�4��y99��}�FTd�/����]EUes��rsU-�zo��:U��S*q�:u�ƺ��7q(�����[JT�A�v<]���ɀG��	:��{����QugT��8����T�3ܡǲ����;�p��N�������Z�ʪP{*1��Y�)al��l�n宬��J���ӽ�p��#ϱ�p̫�
����qh��}���|x��9��d9���T&�FP\:�ީk4;�4���:vŖ2a:�����ŸN���E#ow-�5��(��c�L7��a��������\��t�[$�D��ڙ3�l�^mkw�i�Z����m�k��;C�z�����{�{I�f����N	�@��}�r:o�x��éV��G�P_5]V+^��6���I�ߞ�*�J��Z�R�敯edl��?y(vn����iX�b���['2h9�)�2��&�L&Y^;�<m�AR��K��G��+1燷%w0|*H��6�;y�q����{7����9�t�*pV\	2}�����@��:c=)v�|��9'���Zf��|09C2x��"������`wC�O�	���P>dև������ROY;`~d<N��t�������Ϸ}	�������	�8C �d�Ԟ"��$Rz�wa�$����䞵����!��!�������"�>��W%���O��ӭv=T��kBƶd+1rޢ�� �ҝ��}�?Z��;b�P3���Xf��u!�~y�蠖��h%�nm:΄*����sY�'Cm	"������?�����	�<Bz��N����rÎx�=Bp~���d�>��O�|�8@�?X}Œfq��=B}�^�o}��ߟw�����]�v��'O|{I\QB|��'L�P���'��=d8�O�p}�'̞���	��N�,',�3����y��|��������V�sa�S�C���~@+��t�=����P���C�9�C�8d����s���RM9����`n~��o�>������~��Y8���pC�>���״'̆�8�z���,��N�,')t�IL�$��,��O�����{�ןz���s���?2N_�Y;Iݰ8?RO�r����hN���@�~�=g�C��7���Xv�?'�b��!�W�Y��A?���C���ڻk�{�<�ǌ�זI��ޓ�d��x�ć�4=`z������t��N�:@�����q��$��? �4 ž���>��Y?*gI?2z�� �}�N�97�N�O������O�=@;N�0���0�~Rv�ԇ�\}�\y��_~��kؒ����}�
?O�?"��,������d��;@�{�C��'�'��<�O�	�$������'�{��y�����~���T��u��I�2P��Y1�Y'�z�'�'%�h$�9��'��<`psI�����l��ަ��׷~���>y�^u�����'L���t8H|�����ξ�Hz�P��,�Ğ֒s����z��'�����|�;��6��NR�*Z�g_�4�ZtMM	�V1'�9�N&�r�7�۸���i)�9�<�G��g�K�=g�Ӂ�J]x�`PDj)ے��3y��hG�4�[�w|uL'Ma��%+9��پyI=C�!�?0/TC�t |�_�3'���Rzɑg|{�
�d�0�N�O�X���O~=܂�왹����ﾲ ��?|,~�	��Ls`,������:B��C�����Xyd=d����q�*J���;�|߳����,N�������);{I8��Ğ��Vrq�	�!�'�X~�P�E���w���L�'�Y�*�3P�߸����q}����y�?w��x��$�[	�9d��}�z�~����'̞̈́#�zH��7��J�~w�^������~�������Y;�C���䙇����i��C~��!;NCXN_�O��7iP��VO {kﴏ���A݁��pW��?_��o�!S�x�����'����C�'z}�ROȡ=@��'L�Y�|���<d�!�<i=@7�q���ι�x�sק���/�!��P�L��|{a;@�8���)��$��	����T>���$��~�����l�YP�!�97�Ϻ߯}�u�}Ϡ��ϸ��I=$��I?0���S���<gI�	���8~Bu��$��<d� �����/v�_�k]��y��È�C�@+'��ad��ps�'�����d��`q��N�>I�:d<`z�yC���L�����q$������}�w�������>�XNR0+'jÝH~I�'���7i=�I�VO�<`w:��C����{d<@�=��ԝ��wN��߉!5*��{/maN[��P��W����ފ��랴�E[��$}Cǹ�R4p1E����A��);2�#1���3��1Ӿ �h9N����\6�Y����䷛|f���p���XOVC�t<d��:�'i&�|��'���XOX_�$��N� �'�8~`{:�� �����z���|��Y'��	�O��=Hv��bO�V$���B,�'̟2u� z��|�$����uϽ_�c�?q�������_߻��>	����@鞧�T��&�!<@���'�9Hx�{�a�(�OY��N�Mo��>�E d����]���$Vm�^_��p}��o1+��C�t��ϙ'��9�d�8�`����,�d��}�	���(���,�[	�}����uϾ{����y�Y:d���I�C��7�	��N��!�!�:`w�����x�4>���OP��އ�=dȦ�^<���_[��.��ϗ�?����~b�U|>�X$���Oq�������x�~ğ08�'�*i�!�,����ĕa��1O�k�>G�������|�P��u�7tXp���[$_�:;������8���CĜu`)��>��q����q��{����aQd���|��'{�@�[�q�*��|��)3�I�М3�N�C�IYǶH_��2��s����o�|������}|���L����*O����_��������|ɘq��
��x����݁�	�pj�9I�� 4�?n{���,�6�������>?�u c'LN�$��y�=g�}��3�2{l�g�i�t��y�VX��7��3�'����߼q}y�;�N- ���(惟���X}]c/�XR:���F�w�B�g1ǪP}0i=ƝA+�i���u�;�m�K^_6�(�˷
��xE����̃�>�@d��[L=������z2�ݟ�W޿��C�I��=�Đ�ğ"��9�t��O���'H'~P��~a��C���?}��?����#��߄���/�??�	�����C���d�2�6��ROz���L? x����'('����0�Rp��w�����>������w����$啇���O_BX~C�!�*Y9���~I��OQI?uƓ�O���I����,����rcʟȒ��?�ȋ?�~��?|?�]�O�Y8<�:gtR�1݇�8d�����z�ϴP�\{���'oL�2yl���w��~��?u簟�t��O퇬���w@���|�$
��x��~Nqd����Oa֤;I�&}���d jԮ�<��Y^��'����$������Z������>g(O�<��������T:��~`�d�"��x��O�~y��o���>{ߗo=���>�i'ho1<I=O̝����� �3���M�<g��N�������݊�O�����Ǜ�t����;��d�"����P9@���?hO��a�|�z��I?01՞�OY�9��C~��'�y��Y3}���߾�{��~	�J�LQH��d��Lk��N퓛d�$���x$��'̇�0sHxΘ�$S���������~��z�ϟ����ߴ=d�&E���+'��I�yb��XJ���N�98��p�~�CwAg,�l4�>g�L��#�9�ُt��̭�Ƭ��ɽW�E���Wd�D\��(V3�y���n.��cgc�l�۫��푊h���R/o��ʓ�vh����;B���%�ڵRC�</�aS�5�I��3'h�:�Ğ��7������$����v��J���@Yw8'l�G���8��x��-����ߎ|��W�Bd8`|wOMՇj�<NC�OQ`y�	�%�?}������N��a�~a=���O?{{�O׾;���%gg]�C}N~Hx���3�x�)=N��� ��=d�Мy�J��&�9=��u����~�ɽaM����73���x����a8g̞�� u�x��N<��8@8�'L�$���������IY���ֲ�d>a�d<=;���Ϟ{�~qߞ��'�W氇�:gHO_ڀ|��>d�0�R�:�d̝�����ORz�g�'H���Y&bw�9��u��w����^q�>~����T��:朰=I������P��7��3�	š:O�K���Ųx��s��'��r~��2}i~x~|~�;����z��'�',<������ߩ�X~��'L���(C!��I�Y�ᓀ�� �'�}$}�#7}���nȳ�|T���ڨuI��O�9��>f����I��B|�i�=�$���>s��q݊C���ä8I8�L�$������������{�����8I�\}ĝ�O�<I��9B|��z�����gO������y��VN;�C�I�+�	7+�����7w�}}��8��`t��,>ԇI>I�=��|��w�{~�@��s|<��̪T^��5�R�c�{��;캆�@9d9Җ��G��u���zd*mCs����b�wl.��IL쥶k^�cݲY��*����nf;wo]���ɭ�4�cE5q6�$���[�s�C�WS��WcŢ'����Ta˭�59駣�Y� �|S#������o�F���x�N���������g�����=G�8*�_*s�U�2�랎����_Z�Yu$��F�q�cU=���ٓ�p��O+}/�Pb	IH)V:��\�1�z:������c���mI:Ё�L���W�!�36�~Q��ku������j�^�CeW�η�ܞ�]
K���"�mJ�a5���X疩$�L�91TD�;y�ܺ�}Ԃ=���C�OzIm2��A�*�Ga��q�ktd���`?�z9�|9W���kZj�!͚�2+��u���mӡ6�Yt�'��v�$��ZǨ+�7�#wQ\�`�s첥��W`��A�֪\��0TȠ�ֽZ���	�����[i���i�c���R�-��o�]�e�Y��+LF���朚����_e�φs��n���ٛ�����ƀ��o�A�;�ϵ��-��$h�Y��j��7
����������/;���a*���&n�(���L�ι�U�/]�1n���7�;/~lVh�/��{�j��ϢqǴT�#�-]��35�c͌^�0�4 �j�]r�ݍ�-�}��h�*!�NY5e��̕)������r�Z��`�+�"��&�0��&;1��nZ�m]���K׽�l���6-Zr�hӕiR�e�S����JH6��t�_�w(G��(z�Eά/�Z�&S�2-��Ii�wKG�[��Z밅�&*�n91[��v�{0�W1��]�	֕1���t�uΦ��0ώu�y��eر�@٩��9��ED�����Y.+��t�Mj��@��y\_�%ܔlz�=�)6���Y�w��1.�4��62զ���N��A�	0�¾.��f7τB��N-�-n�E�+%�!%�R7��r�ܙn�;��@��,H;��w����v�+"����k]�P��T�i�tV�[F�*F�] (��\�.�Y&[g2ଆ�p]ab���E@X4�ڨ67A%�NOk����Av��f�ҤD:��Ƃi�}�v,X�G���:#x�}6�7.�Z@i� B�����јؼ�@&K�5yY@��a��kD��՛9��
���/�;���
ByU��ջU^���F�@��ڀG3�6s���Z�֐����%)uw�!Y���Ѥ���Fq�c ����s�E�}��bn�Y|����dH-WKm���:ΰ�T��o`{�6�+�4G���J�݌S��:8ݳ��U�|1M�N�k4�B�������{�v��-�T&V.k�%ؙS�N<ta�����i�^h};`O]�[�yK;���:�T/5��]����mY�K#�̛*9�I7uo����k�
�R�vc��Z��Sj5*��]+[m��j]J���ZVѕ���Q�E.��ZU��n�M�Lͩ�)TJ��ݦ�%���6����J�TT�ETԮK+JT�Q��p�U�����m�p�m������mS4X�l\ܵ�u�Zʺ�"8d�jS[�˚&EZ�X�[Yb5�j��n�h�cB�Ke,AA�j�u�mZ-��جԢ��b�5[�T�S]��-WZ��Q.�X�]���jʭj.�Kh��cV�9V�ʵ��KKEPE��F����ڣ��YmZ�6�֢ح����lZ�+b+�p��*�""+Z�V+����X�kU��1AP�*9��dU�-�,�A���5��i��ER�kd���KB���uu��(����2����?��z��]ف����qz�\�yKj���z"2$sz�r�
oIa�=��)��O��W�f�[��#�ѯ�.�C��s�8I�����~��JïUe/o���t����7͖�ך�-g�ܟ��'a79�%/S�;��s����+�x{y5*�ޅ�k>�
��Y�����,e1jȱK���{'l���{�Iȍ�\2�A��mY�o��n+ ��+���wy4�b�u�����I�+��(k���*�jf.2<���;��܊�X��G���kCY79=Ԙ���W�IL�/�TvG��k��}��fK����>��R�-��"|5}��hd�򮅼��y�h�Zk�E��(\Hj��_I�U�]71WWq��{��d��8罍8�6��v�
^,Rp�E���h��tQp�u�;��l]�ͮZ�����Ai�t����V�FqJOv������rކ�D3u�J~���}�"�O-'���jR��,�z����:5�Ei�5�=T�挣�!�į��X7�����돱IҞ>ۃj&�1B8m�*�&�}�b�'1k}Ԁ�f�_�$�sS�z�\C���eF|�ڜ`~��y)��o&{��o���jѦ�*�w�ҷ��2d~�����z�b�MMN�gj��cU��d�
D��q�k�mv�S���2>�"��Q�nF/T7��+�#��W`Yg}%�9s�u3��',�J����YrP��6^�0�ɳ�6�v��M�s�佪૮iթ�oiN��3aNoH��ӏ��q�Rk(�y�"*�:�Xw�Iٗ��jy��o�)�d��ekR�E�������M*:�H�r�_C�5݈�u�9tf)�KRd�������]�^���췚�M��u��3��.
��Em�Ͼ��7��8���g��e31�~Y0���*�j#�Ev����:�{zOI�Ѣ�f;�X�>��C[�V�@L���^��$�я�[yC�������5�oݨa[��v��JSS ��
�xy<hT=J��3��\
gU�W�:�y��J�����-3lS����,X��ߍ��觭��:�Э6`�.)	p�1(p��uw�1�=q.�5��R]���
��A�m"����\�ɧo���rtm�oɚ�ʭ�.�cC;��ʑڇ&���w�o�m���z�3hCj�f7�j���\����3�2;��ط�����eclV�\I�%N\#� WBI�dü�/n��V�A���9��,���ޓ�P��]S��S.�J*P!I��m�|_j�[�vkA�S��l�&���fg-3�v'S�k;����}��}�ϓof,�v�[�ܷ�o�k���ۢס&������5%e�<�	�R�n���q��j�3J�!6�q�O�	�.�f�1�]_vK�>Ċ����/�s��$�=�ħ�2u�p���G�˛��Yn�e��I�Xb����e+��*r���ϯVM�W�{$����f�ESg&��P����ΐ�T6*�`����б(�T�����J��H�9fkܫ'|Ͼ�X�8����y_�o�o֬���9I��������ܺ=�_��J��9ح�%�,w7C�_
���r��6���!�+���^�����	w"z��uxTd���(
�ˁ��RQ�Kz=y&Q��m��C庨������A���ծ�(͍�R�o&�T��n����V�J����Q�Ҝ�������9��ծ��i=���>��ꠔ�zx�g��![���F�Uӏ2�x5��Þ�S�_�יջ3�l����Q���7��o.+j]>�CȪ�U��z.����E��2�"h�ٽ�̫���='��'��z�P��B�	�i??4AO�����=���o<ҝt�A��7��S&7�q�ϼ%֞�?k�8�^��;|��`�l��z�ùkY����^
�O75>�r�
�Pz�Nϼ��G�;}�g�)szz7 �~E!��.�[_ct�튆)�wxӣ{v�������N��^1����e:�}��=���fDm{�1���WyB��(�x���A�ږ��WG.o]�v|	 �׷�-�g^U�5��.�<��k�ﻞ�=rw� U*�c�TU���d��x�]w�mM�"N������nZ���d����3l������G?>���%������]�����ub������A6��{ێ�폔��^��������%a�1uߊ[�듥mvľT�g��i�?��
�쮙������CЧ�.�lr]�bɨ��q�4]muYL�W�!������ug���S�� ���P��Up�YBp9�#]��x�z��g�7�u�:!V���>b!^�y�=��,�r`K�̯I�Z�˿Wz�)�*8m�*2U��w�s�/rk��K�f41�uS�()���^)y�~��z4���<����â���<��d�y�������R��z�%,xE�V��u���\��~�W�s��o����ᛌ���<A�p]�Ǔ��x�I��E�϶��g؅�]�z�5�ta��L᮪���qEr�A�\{�2��sw�`h�C5��Ks��-�H��٥����Wb�����_}�W�ڌǖ�*{2��N�}�m�b��
��X���ժ��&v�8t��ၽ9�DmYrV�s^=p�Nغ�����T�^yJ���LF�h��EZy�V#���N^����G��`�p����o)�;��t��zzC(��x��z#�^��Ԫ�ƣ�'�ː҅��~�܄�hp�@�l��ylǾ:��O�fzB��]~^Q��)�j���i��q�]��<Z�*��*��}��g�1�#�0)�AK?:aѻ���*g3f�1٨��el}ϯ���VQ����1N�	�q��#׹�Y�֣�{X�z��`naqlXI�b8m���nR�\�|����z��*Kl�Z�=��!�T�j>�����v��ƞ��f�Ug��c�yYq��⌻3��r���mk�4%���!��sm
qӭӡ���U��g�Y��7�K�=@��1i9G�^�(��|�N������|�r�_ ��P1Ǳ`�U�aV���\]bn���6�榦1�'��o�\j�38>f��g�u�{�F�3�u�4z��Օ#��Ǉ���'�}�*��6���I�+�{z"۩]�0��q�v���k�v���/.Z����1�-��L~�'��y�����{&2�6H��uoD��4TܙLP�V
���g��o�a>���,q:-���.��/�֒!�$��g�J�{��ԷH���zX��12�o���ٽ�î�x����sQ�#�Q��4ҹ]u9z\��Ɛ�շ�^�{�N���w#WP��v�_�x*�f�ć/mN)h��ԭm?o��y+�q�M�WDs�hr%$���:�^�^d�&�z�.�԰�*đ�f-Zcr�$��7�u���}��~I�I�?^��*K�:mfE�k�$D���b�US�պL�=�_�Փ�A���"ǿcˬ򗎘to�T�C5�4�B�������ֻ��R�S�\M���;��(��3�2�TԨ]<�³�-�zo����1��͛�(�'��[d����V��\�ꑯ�PnM�6��H�(��wB���˂�U�/��o,EBڰ&[7�/��Oԥ�c�b�pῚ2�"k冽���c�t}�5Twuy+�S����g!��N?5�ob>f:��8_*�eDs\��Ӆ{Nv(0j���
d��d���a�������y���V���C~~s��r-{�;�~Kβ^Ef�=Oۖt�U(V�h�� ����U�rd���/|�7��ݺ��ܒ�=�Ԡ��1�Yzy^Օ��Z��'oD\Z�T��E���l�\W��9�U_WԷܹ�;�˵��YU_4=c-��oF�Ȳ������#q�긳�(*E�L��e2�P��[]�(tЖ&x����'}I��x�r�W�#Z*�C+D��ެ�;~�8�Hڛ�a�Ԧ*���8�R`���p�ȸk���������e0�g�2~�5��޾�O��+y�8��O1��pU{�J�2�n����Qc5S�g�gB����n���	3��k�^:���5�r]s'y�z�<(:�Ae*���>��9�&fA�ܻ�����h�f�������,/VP���u+BY��F��ʰg����[H�>�D+­��x�~�o�ny�P���PeC� ��t)F[W��Z���Z�w�T��j��oi���]ފ&JO�J`l�����f馘-Y��=Oj9G��^���iDr��7]D�lKܼ��]Ų�����&�T��[p�%���Fi�VQQ�!d��ޯ��GP��� �����[n�R�]�Z��0�arى�[@5R;��5�y�K�1Դ����}�E�Û[����LA��_�����]c����F��.b��8˘r�;ZK���n����曗]Jc�{ܯ9������d�}���W���PY`C���o1��>[����l����te����>��Vu9L"<kJ����І��ۢ�z�J����d6�:|��;M)H1�}�#�~X����2�:Ѕ����	���;e�2V,����x^�+��L��]��@v�fM�e"e�@C'*��c ���5�[#�������p"��g�|�u�]��Ǳ�Ú�酰�]!9�.���R"b�0��Ei�b��ܦ;�7�Z�t+�C�V���{�yIGBN�]'��Sf�C�*ժ܅Eo�2��'����M:����CƏ�#ܒc����i��^��,���g?'�C0QF�n�N*�(K/*F~��"��#(f�"ٞ���$;�� 0��
���� M�	9��q���	n��ǗVbr4G�D��`�sTіU�a�3%�U�P�G4�WnBç����Wk֩��sR��f� :к�2�Ȧ:Ybڬ�R;�+/�"0��Y�[gw���H[�A �8�:�l'��J�V���O{����S�hÎ��`ǣ��L����c��[b�n�tT�Z�L(��ggu��:��7 �6��l(�j-	�uKp  �����[��8e��	�wy�i�)�����/1��G
��z[C�"�x�*-��:���\�%�۵�\��u���^T���h�[W-��Sv��ؗv�s�`����X�[��*,�L䅗da�`.rޜK�r;X�ZL��"Lɤs_��0���̵6�m-i��e
�+jg35sDT
�PW%UZ���MjV��mA\��F�uF�\��*UKj���0bU�*R[\5]m�	R�u�%ԣ�mkkJ�-Ej�PuҬnM�K�,Q�����X��3E+-n�e�s�rmZ��R��*�VX.��Q\[n�QXZҹ�5Z��̸)u5�BܦX�.���i��C#[.��kS#Wn��Me�Z,lH���+�D\�-�Ҭ%k�˩����j����k��Z��b����fM�ְjV �k�"�i�u���hR��ԮV��)nGX��J�Z�ڕ�9��Ubͨ�5u�Km���v���iD�Q�]5(�5.�Mu�4U�b��	[�f�m�*2�ըZ"�#l}J1�C���r�`��n��v�
CL�֦�Nb�[����*�N&]��^}K5�X�'�   �i�&y����W�
�	CX��W*"z��]��A+gw93^�r�U���fD"�;����W�-�v��qԽZ���6��+|��]��{d��w�ϵcS)�G=����z&rgk���ɲ{�'�X�xb��]-�L{q���7�+���ǯ#ceZg=;��%!&���3���O����A�����q�@E����u飼�j��s�wE�s�H�����9�=8�>Z�`��{7�W0i��к�֛�~�5����8P���v�긧<�v�}�V�xE�k/�����)��WP��>�3S�پ���!�>v�ץ�.(�z���rAW3D꽽+p�]aXv���I
c�����1%�=4gN��ٲt%�K��kLCe�Up�]:[�v:��t�����r�N*���t����������-i^�^bGu,������>���Z���y)���{>�Su3O�F��w.��df��ۀ��(�	P���n��PZ��g��ޝW���$9'��=~�v�%�131M<C��'�Otq矋�د:A��ń�7$;h�O�/���9�*}�k�V�h��v�h����ܐ��r�c�Z.��|���k0GB��Ƈ��V�7���#5"�ϧ��q��w��K,�<�[/���[���q�X�X�^�Y�o����Vr&62߼r9\"4�
�f�c��M^���_�^����?�W9���ENɎE��n+}�ڱ���ԏ![zST`��aU_PyQՎ�Q���v�O}0e��Ҙ�{�7�/�V�I�+m.U�7������ �M'���vW�A�"��͏zk�u����f�B�9�=�?L߃9B��%e�b��k�Gz�M��e�����&%��Nǟ�#�2�]C�'+�ȽE��w���3G�N2�D�xۣ[��^U���s����E�[�>�P��ʱ������H�ǳ�6%�\z��to5�C��X��ӵWӅ�
���3a��Rg�\�թ{��M���V1gOV��R��n�~�X�&i�����纣E����S.�Ԇ���B�t�^�nU�,A7ȗ�^�*r9z�H�Ej2�`e��z.���ؖW\FQ�������[Z�쀩[�C�G<��d�έ<]L�YghQ��r�q� ��C"���~��ں�W��2��].69z�"7]���Yܹ(�˳+��¶������mQ�;Nq�1����}�� ��i����ڂ��e��hʸ�����oec�_y&z�<�Z[��{�߱� ̌E��ո�5�n#�����vc���e֭h`��̗�Y�_��*��izg��^lN�y��l�ܥ]&Qn�AK�5���w��S��e��7b=�2�m`����9ڡ~��U����ٳ������0_���ĝXy��PT�3�P��]����x�[;�2�j6]������W���r�,��3V�~�9���TA��ue?ˮ���HEy�SzU��[��2`�u]dx��ug�Ud������Ú"N��z�JO�E����Or^��ѭ�/7�讹��Of��T&�Z�D�S�!����<C�gU�gH�2�.G+M�����O�iچKÒi�:�-뫑U�*,\����ITW��Pv���T6�y�S���_W�W�>����.�����M����)�ǎ�/�\=;��}�MJ&ꚂURJ�xh�]|4�^Z�qZ�|E�7X���ny��=��/������D�!�{���~��+ނ�C`Cͯ�:6#���oe��y�n���y�8��SxP�A����ѕb2}���%A���N�ߌ��)�����;�{��\�H���{w���N�'���2�y���[����M�zq��7�RS;>ɏ>��Q����c�2I��^�ܞ7������^Y[��G����c�}�UF=���%��&j�#�jW���M�����5��U��=�޻�xbt-�cY��z�g��zC�:�:�[b[(�1���@ͣ���ͨ�]��$[(v�X��z�Z����3ͮޭ	�������=�)$�[�"Q�B�����1WU���.���˒�w�����IQ�e�Ͼ����-��������jѨ�f~raw��#w&��s}<!=7<�G�n��M^E�}�j������>�ͧ,oD�tΉ�s�u�.{֙�}�G����S�:$ؽ���@A���t><󕻍�~�[�Py�d�y��sm���0D͇�i�R�������To�6l���׮�]�7C-�h*xЦyފZɐ8����^b����U���X�Jx�(X���-3lSF�?o�H�p�B�wb���V=(#(g�Sr�z�Mx'm�v��e���s/��%�S���y�^�b�Ѯú�a*okq�x�E���^y�v]�Ƈ��?�P�q�V��y��=_����
�}��&ؓ>^���?Oz�c���`��Z;����7x���x9$NܔA��|K���U}�Wՙ�r�������8ʸ�,5��XA�!������!uJ��P��'���;<�Q�����`i������?k�ekg�A�l)�N��h;��z�v�1�4���r���|ňᱛ���dX�,�U�}������M��ӆP�vvZ��d� �g�߾]C�z��5��fz䞓x��T�yLti��)Q�L�o���-k'�����K�y���i�pkw����VG��R��p������^�%�鏽E{��j= �Rb���jӥ�/p-~Q�܀x���jݣ�}�ŭRcWq�`?�=^�3�}��\�3��.�GDp�_f��Z�)Uzp���5�xG9��K�Q��	��eTUu���� loQ>��r1*��w�J��������>| ����Oe[�"y&O�o
���R�:ީ��PkJ��c�0��/Ey��vbf�أ��U���V���R��b��C[S����k����-�dz���&ojn=��О�WÕ��_��^�Cp<�O(lyw���y���N~?���FM��W
տT���ګ��
����-�f�lXݱ��_EŰqޣ�9E�����!���s��[~��}�����FU�M|�׳y�����,vZ��<ƜyV�U�#�K�4����~Æ���Ã��ո=��9~�#�����ֱ4ƨz�i4d[3�Vy���-�3�w6m��]G�ԱZ{ˬ!�/m�!�s��y��5��%����ڜ���$��XC8�|�1��Cۛ�+�o1_gZ����;��� ����%A�*b�m����զ�4;�`ٻ�H���v[����牼[R�e$���Rkբ�V��
�Zԍ�.�w,G:<ǜ���r�UU_P����o~+�|��W�8:�V�3Z%��3���0��mו��3�ޗ]o��
�
��c���ޏE����k	�tzF�1�Ϟ�wMІ/'�� �P�Q�����nݖ)�V��x��ƢN�gƦс�\<K���/��֛�A��գ��ۉ�f�#G���'�D��8��
�R��G`��g^KWǗ���P�oB<�dpc�n����u)Vj੸�#DV)JɥH��CEӖȣ���_�f�|�������Ϫ�&R@<���1c5��в,�YvL�ԽDI�o{3��Ƞ�<%a�����\!�P�;��W��]�5��]{�D�s���2�F�u�u�˰c�"���qܪ��ԫ;�O�j�ż�����i�|\�]���0��G>�:lh���E�lGR��t����9+t������[��[!�)M6�o�4U=<O_a�F���P�����<����=���H{Y(5j���N:��ڳ-6dһ�
އC��s(�?~ > �o�9)��������K�a���H|?8��T��<;wJ~���oKu��S��%(�~�7%��&��"#<k--�^rEBc�/�餂�}��oi����ٞ3>w�}%�Ն�x����R��I{��}��c���3^#Ζ�a��MD#�;��8�p����.L��3���>��gb��G`�H׈�/�J�S�e:oR��rܓ����K*u�Cnч6[86[�>�e*�6�gJ�iW�+x�O(�wQ�OU@|A��S���Ge�<.[3G[:G��ex�mV���)m�穑�aT'ƶ��B�8�Jq�t*|�T=XͰ�ԝF�ό�O}`�[_e��r+h���\��s$��[Z���m�Ӿ�3�����F��MN|[���@p_uL��RQ��+���]c�����}tCU���&�a�
�L\=]}�q����yv���!Gد�uT6ܷ�)ҧ�Bh��Cw��S4e֞!��%��s?>F�S9e��
oZ���٧$V�`��NG��%��O�6�cRѧ�P.�ęC�i�}�g�vZJ��|#�suq��kn�!��慄�
��ݺ!(Z��˗O����H�b��{-�dm�*�=v'\߱σ�p��D�����v�*/�w�R�_tB�w��*Üj��C��y"���=��X
��_k�(5�]�ʓ{e�sk0� ���û!�y�q�Vp�u)GJLD�Ւj�헛��=X-��������_R*�H�R�-���
 8�N&�¹�@QO(�W�ց��̬� B
e
� R�s���n:���nok�!<�25Xom_>.:��|%Y�AE#���(�����+�S�YukUM�RG��
�������l`i�OC�6�'��ӥ�;�7zE�D�Wv^*���O^�oE�W�&j��:ts��*�w��!-t��Y�:��wԋ���C�x���C[V�!s�}�v鎦*Ռ�-WF3�[\k(��s ��_2�*A�'o���C`|��v&u1l*R�l��J��氯 u���)��7pN�е9kV�SS�ު�Y�}N�g�ĻRިT��غ{%4�f����q-�R, .ZZ>y�a�|n�C��j7��cS����C:�G����	,f��t�a�����CE��*%ô�ū�y�C�m,���M�qӴ�\�)���B���ꑄ�ŔZnJ|&tu�:��AR��.Y�4^و���'|�_|�*B�#`�vg�l���|%h�?DL���ޡ`�v�6J�YlP̧,]�&�+��$��Q,�]�����fSO��J{��8����Dc�8�ꖮd��.p��ͭg�KKy�l�k��u<ʴ��[Xu�wps�$_���Sό{Z9m�jճ'j�d<K��0�]]�Q��[��]��\s�����L���-�z$-��?s�O为�ljZ�Y�*�Y�nS"���5�R�P��Za.*Q�#s\U��]p��\��W&tIm*[�A��P���f��1��D��mSl1\��V܉�.�֙pѠ�U�[m�5æ*��ũ���d��Ѷ)��ڸT���fq��ܙ1R�ҙ�in��AqB�ַZm�)���gsu�S+WV�U�˩���1��Ʉ]��l�-1��u����v��E�qu��3]�Q�.�VdMhkqX�E�-n�3F7j9[��t�+m�͍�8��2a֔6���L\\R�Q���m���Z��ت%.�eq��Һ�Jm*�\�g��\&5��S]2"��rcY�T�[D�v�"��mffecm��Z�̅b�SZV�m�-ҙ���A�9���3Gkv�Mu.����5�R����-3MmB��B�Q���n���6�jJ�ܘuZ /�� >$�@��7==�T���3�Wo5g���tw��#��onLʽk��nY�]�!q�7���_}�� 7�ڜr��%��G��`ϲ���e�U�}U��J��#����ӷ�O0��2��"��#��&@��*
�U�X5�!��]K�Oq�=��fTz��*P�<.eӢ���Q�GGQ(�k���$��"H�5��T�u�T.ϼi
�4�~�M�doZ�w�(^�6'�d�H��%ʨ�a���[tE���h�f䱫�
��eYQ<�����+�V%(]�tX�A\ʲ�C%i�L�P�z)�^�C=���`&ڇ�=�\�肑�����g���GJ����b�"`�r=a��9�8,!�8/ǨJ��3h/qW�z�]�������{3\���˫X(�5u��
hb:B�����0�\k�A�p'��f��y���H��>;����QAR3M�,OW���<�~@-z
*�].���]�{0kk�p��}�P���H/-\D�[��ߓޣӂZ'4�����c�7�uh*�b���2��"E����{S�����
�������.ȱe�[�i0�Bu;���.q=���������bPؓ�}���k�|r��Â4r�*<����r�s�����P.�v�1V*Ͻ,v["��������|�2��Id��V��"�r�f��|5��\����*�{|)3\{���>.��H�����ֳ�'��iX�k���𰇄D��0hSU/F�[������<��Z<Qs�L��y���K�k=���|,V�P��/~�Fr�ő�{g��e:B��E�[�m��W�=n�Q�cD<�*t|)����vL�g_H3��q�9��6ݳX�X�o�T<������dW��%�����ծ�@ +(pt{t.�Uk$p���b���3��ng��֯�M�g6���X2��$p�7�h^	�Y*|��c����K�wI��}>��2X�cÀ*�+֐�K��V/\�p��ܪ���@ӯX;�U��x.2L�f�R�C�a:+��7���K�c�ڲ�ww�:
i/����X��:����Y$n��Χ��xI{�V�ҽ���^󫋐8�����S,(�I��s���ﾳ����pe~%
l��c��P[�H���k�5)ʬ=���4���rR�;�~>4B�x\:~g�ݭ7���(r�eI��YT�z�M������gv^8�p�烨1WO�h��m
�O��yOg(�X��M��V���\��}样��౪����WQh�Qս�ɽ���ˣ�hg�|gz��P�S>U:�;F�I���+����z�8��<�,UU�!�%�F�ã��aU	ŭ+Z�(�7Ӯá(x��n���w���� �i�:?h���ש��}��Wp�y)ĵJ(u�.�S��/��"�)�85�87Q�6-㹞&��Z�~Y+=f
���S��'M���E�gD�p���Ϸ�{<�yw�%���*!SN�K4EE�Y�B��vQ0�SP���uՁl��]k��-�;sP&�d}<S��qHx�)�^K�3r��G�O�L`�&]G��J�ke��6J{]�\�k�>=��G.!�\�X��l��'��}_}���iI�v]~X��|`�,S���e�x'���	�B��b�O76E�6��A14JT	�S)�3�Q����O��ĨPl�7Yl�E=��;ȷ���!\)����R��:��.������8k����gM�r���Vcf����D��tM0�t)����6�C�"9��w��t�S.3C �߮�r!u�C����V����(o�fnA������x�8�������,�q��q؞!a��G�Z=,;<Ucw�o��@���=��zg ���~�5�g�߃�E���U����ޥsW)z���,3��\5����
���9�ķ�<gn�}�D���~b��*̪G�H,d�GV,U_K��������s�u<O�gOr~�����=+��E�-��n��YGY��0|���+U��FW��΀;�;(��3F�Ŷ�e {�����Y���,��SS�i�j)�{yfvTl=����õQ�*w&�O��L瓒y{��C۾ƺ�<��7��  
��F�/�~���%������ɮ�eR5):��?�!��{��w����K�;�Wt��xl���V�?:F~_�m��!��ɺ�/��-m��ܝ��C�V�e��k����Sh�Ur(�(�	7�����{�kL�6�C�H���`���T+��a�f��,��d��zy�ݓ=3k!<� ~����б\<��U��K$|sj؏^���D���0q:�D
bU^1��|ņ����d��{�Ū$�]�(��n��`7�*���R��
:���{�gN])�5t���$X��J���a��f��IBeq�#'�L^���ܭ��	�æ�lѹ/����]@]j�Y"��7>K��z��b�Oɧ��;3�J���ʚ(iv�eY��ßJ�Ν+s�!{fż ]��Kh`#zL�菎�������W�k ������֥_m_W!�=n��هv_:&2�sn��H�WoK�zv�g��;F
�c�&��tjc��M�<!i�.6$�<1��_}U�V��^���&�U#�G�ŋ�a��*��MV��K�Z��T����*������z��.}��d�U�e탂T$�׋F�l��9	w�zz�~]��q����Z�|~�gn�
�g�۸Y�UO�CN����b�'�ҏ���b��/O��9u�Z�W*��t2*��n���ٓ��b��]�mZ�Y�X�n��P.��^0�2ڝ�oR�B��<��B[l���1b�_�5Ƭ+��SRlZ��sǧ;ǚS|I��UW�+��^�f��>б�ch2�,�Gp��
$���Dxp�n���M��1h�8Z0Y�������qM�:0��Ln��>^��H|�uU�wEz�[��cEg����i��)5f�7ͺt���(�`�ag��|O���qp�!�a��!�<�iVVa�ė�,)u��Q�����1�5м�M
��P��*@U���U���b��-9�Q�,Hx����+h�癮�9o\�ݣ^+����i5��6�| w�ة��g19�G��;0U�f�"KT�/���s��¸���n5���u�Z+��!��^�����B���V�GF¦�ut�&{�o5�tΘ1\#&�C��,*W��tG:�^m�q]=�g&�e��Jy��v��w��XӒ��Y��Ӥ1b_�){6�_�]1�V�p���z"ȗ�=��e� X�>��hӯEé�pJ�%	��)L���2W8������f�ۭ:w�w�����]�^{�yMxU�;P_�e��K�
�3\\]E�����M^-��߰�/�^�S-���uuT��%3��׊]l�pvd鰪آ��l�K=V��s���z�?.4;��������E�g �J��[����	������t�W(�����@�(p~.���f�ދD����CgxS*�D��y:��Tn���X����Ϯº	؆�-���@e��F ��:h	,ɵ��ͦ����&ՙG#��$Grsv��JeZ�0�l�="��G?>�ꪪ:Z��*U�z�o�p7RٕL���
�'�ڳ,
���0tc�2L�|�l��f=u�>wd����֌�.��5�9����Ζ�C�w}G;�67�歜?O��3q`���"��8�����gw�.2�����=�=��}u�<8�
`��ЪF��Q��D6|�����3��2Z>?k�=X*�%�s�mb�k vn�"���j��{�G���2�.�66��L��n�l�N1A�P�f���|=�wsy9��4e�૨�K�H5X�!=T����T���t��M��ֺ&D=#v�v<J>(?��!WX^LM+? _��VPa�E�z�~�z����J��D�{Q�|�N4����'c9�I��[�~��gz��Zg;�Y�0Ñ�4/r�aþ�#��A�F�`yDJ���g�գ��.�|E�l8M����;.�>�j�m�о��OV����u&e���/G\�)E�����w-T����;�%�c��t"}�6]�\���P�tSp�r~}�U}U�G$s<��������˧l�P�b)�#G�\Y�hvH�(�缾�0pC}<�s���B�c,��a��#/L�
/:Ĺ纬����{hi�´�VI����$zm�k�����H�G�_\kN���&V�Â�CLѯS�↛�a�L�U�Y��]�q�nskl��q�P�ß��J�`�h�J�f���1���%�߶�]OF�Z�Vz��0�z��ۇ�;�=���Sχ�W@�@(&�>W)m����ܬt��x�P���e�ƳHE��d
� SS�-5&oyg|��7B:�ޯ��k���қ�S�M��G�>y�i7��%UK�O]6n������F���t4K�ӓ�:C�T�����oy���!���X<g]�F�|�UJ<,5�4�>�+K7��&�o��lʕ��9�t�`{f��6>�%[�L�^�WU�k��EL���e� [�are�ՇI��jR�ݪ�V�yI�v��:��Ȭȡ���Ϟ��.�ޡ�eo)��~�}�|+�ڹ>��b��G�ѦeW1Pڣ||MA7�Ur�|��ʚ�<��E�q�.�nT$�	vk#�W���|Yˬ��,u�߫�jٚ龑O[CL�fW�x��,��*U(�i��,�kn��޿��R���L���_�?Om���?v�ӎ��ҋ��×	ZY�<v�r}�{"o�u�2�ǳ�E层z�HP��e`(�R�U�ۧ��KJ�$ɡ��^�YCN}�oo|�.!%|2��UqMK�r�3�&K��x�y��N����iѵ��GN:�>�eT�����^��|�y�i�V�.�� �$-q�Z�c�%�il�(nGWH�˱8���ڭ0_,G~u���Q�v���5`S(�QB�t5N�$�k68��c�Y��}�a�w�����z��`ƮƸ�a���s���t�P���<�
]��Z�W2�9hT�*Kl����cu�7K�S���-�nJ�}5�g #���,:D�܈KZKKO��GXS&ꙏ�m1�*B�f.�g[�Yr�ƭx;x둧�a[�1�yXv����<���2&ye�v����~oN��ҧp�8���r�z�;b<�������#�h��E���@��2�{/g�V,�<Xg5�5u��"d�ied�ֶ�"�x��#����](�r�Ĩ|P����oe-���P��R�2��o]��`�)c�����A<�ߞf�r�ȭ&�n�޴b�o�f�Դw��,\�U�����C:��I�e%L���M>�e{�,űs�4����W��^$й3�1zwj֛�P{Athf������v^Q�3�<�9r�]��\;<���i����[@>vc9,RRn�Y�Q�ul�J��x����m�wK*!��Z�:��-��������#�Us��{Plk���CGe����,�Q��;�,{�V����fܛݢźE�v�c��Z�ö��+̈́��%r�"�`T�����0�5�*���[t��$kl��x��$m�U�h�WAguE	��nj����8����4��!�Rs��M;�5z+�����*:�^��v�J��b�ph�<��S��B)_]]�^ۥ�-����^5����u�S.�X4�^8n�`��%h�S{5�I���BcTj�[D_��(���Ga�c8��&�-5�*�O��|�,��t���ע�-)Dq\צAո�q��FlyY:��2S����&j�7LչY���rcN���m������s�;�ohR�.ɬ�w^3 w��}��g+�B�@3ZI����R���Ҹ�Uk/�دE77r�uqs�}�7��-��X�WL��:�s�pǣ+�e�ܝfȊ��Q�ӄ��d�c*��^ܦ�2���Ū]�;�Xh�"�䡦�B����`�a�0*�$�dȋ��]������v1���y�m�5���֖�p���Õ���uyj�!�Z�O-z5.W��9[�Z�N��]�%�q�b��F���PdZ�YB�Mt����[嫎�V�}Y���xy�i�c��k������qܧ*V�[]�u�)�u�Ϝ��%�l�6�p�KJ���u(3�c\T��YZ1+�q��ekL�����5��Dc��֨��Z�T�U�j��Z���q[bZ6l�&Cl�M��kbQ�F�u�[��YW\�Ʀ1���,F�-v��E��fK�R��qp�%��P�.�ƣJfۜ"E5�mU�*]J*���j#��[�Z�`�RW9�U2U��\f��9l�ZVQR��TQ*Z�\�U-e5�@S%QQ��%J`����+
*EZ�[��d�h��M�����**��u�Z&`ܢa*[�+Z�P�R�B���(���TTEU!R�h�ejUJ�m�U�U������iU:[�U~kO~��'kV�	��k�ˋ��kq��s�dY���9m��jc��諭��^�2�U�
�6=}���WP���k�Ȭ��U�k�,�<��"�����A�с\8���1ha��(49���]^����o4��k0b�407�U0Y`����Å�-t�4T_�zd!ڻ�W�j
W7	F�W
4���*�Ҭ6�r`��
�%�Z0��+�y�<�����(髻
��P8:�$�L�)|���}Y��^�S3�L���(x��2�p���.��l�-�n�	�-�,��x��z�p붽sWě=�qT"e�:h��V����ʦ�Cc-���9��A��Yc�$ǯ�T«�g>UlV	��o��/�i#�q��w�{��q�|1��R�
�]��6<s��v�M�XC�'n��L���uF�;y����/��ƈyBh�p���U��
�ev�0�y�3�7��\��zN�h���wl����}��T��J�����.��h�vʹ7u>f���4q�/S�+������	�*JV͉P٨�hr�����]d�H�s��Ȟ�*~}U_}@&np؞ɤ��=�h�Lx?����lR���A�,=�*�m���Ч<���5J��p͖�u��������t�:'n<��n��[�'�k�U"g���hvk�|��c"���t�q��������<���珌�A�qC�a�˲8�;�����f�_oG�a���G�\�����QW+�.��lî�{�Jm�ǝ�g��K���gWy���'o.�^�=�U�xB@5�崴:<L��k�uV��9U��O=���-QFT0y���u�O]3E�ƸRߍ@,t�^�p}��h:�]��軋��:��ʒ���(�
�T!�*B,��wK�)ܹ<�S��<Ycn�_�kE�.����|��ގy���@Q���zİM�q��_z�Չ,c�Xxe�"ި}�.��o"�C�(��q����XI�m���H�*r=j���0��)�m_� ��W�E;�Otל3���4�w�XIH�S'!�[�>��n���.��3�_ȈA���۲!�	�W1t�]!λN�貲0Zpi۱]�23S�r�����mɭ3u^,��Cch�HR/yT��ui��
��N�����`�#RU:���74�(�}��ͬa�����g����r$}��q��O�%˲*Ę�5s�{Ѱ�Ca׽P���t.'Q�x�������m��>�ԋ��u.��Ƙ^՛����L6'\7�_��>�O��yj�]b���UC��FV��1�:d�#k�`߶��tE^�ܛ�� ��ԕ]� ��Kb�T����0�����S=۹������:�ǌb��ׄ�,���,��I�T;+AQ�U��y�LC;�J1G0ͮ��R \���7�����p���}��ؤ4'�rzC=������GN���BtAYF�PTN�𺾴v]����t�-G�n5Xz�tӬ,e�2��)Ѓ����
|�G�B���-U�WG��\)���9�����ʔZ�s�I��i�n�as�7�Vb]v[��������(�Q�������ε�wɢ��ԛ6�����y�=��{��-Y��-�T=p�5xB,ӢD>��J1�p�I�Ƒ^l�Qוxe�p��ʥ��
^����͚���ź�wY,؂��R4Tk�|�}R������P�Ɯ��w^��]є}��7�*�K���w:<<��E$@!�J<�8a2�x��jt�t1�>48�+�dw*�1^��4�[ʊ��C1��×���i�v��8f��on�(�$Z�n�e{ʆ�U٪g̻2!ON\��V�}t0(����}lђ�Tt0ҋ(��"���ivb�7;WF�]^��p�C4�dg�v������]�ɵg~��E�#٤��1rSb������W��d\�0/�A��(|;�ρGMQC~Yo\=�g��4䊏��+�)Q����PX��/�P���3h:��zgh1�X���5����4�ܛZ�=:<���d��mK�|�\y�B��WB���ק֮A��l��q���nկ�>�jx�TM�c���n@e�~�;��]�����`�]ǜ�綹�Is�����+������G��G:���[��Gn��[h�B����o��Ե��Fd�8�d��!�U��֋��n�5EO*����.��%^�{<ܙ��<�U@����a�f���I�Q'��[�x*9��IL��~p*����W�u�m�k}��E��
��Tģ���'y��B����L�UC0W]|e��e�y�}��fL���t���x�'PEl���Cb
�tup�a|�&��H�-4v{v�Ah��{xȠ��{ي�fm��* �:�x�pߩyhl��c_���K"e��w'��Ƌ.}v��wĭ�@嫫ub�*�n�����Eu�m�%9�r7gn��A��GMm��m��4�U�]�ts�W��6�)�$�X���A�����Id0Q��)f뽵Y_xb56g���r\AL=�G��_��d*�K>�	�ɕ���sƇws��z�l�>W�yr�W.Je���5͡�vM`��Tt���K�ݹo/���2�La7�Z۳#}!s����7�9�*��ݖ�Ua�ѱ��72�,��U2�p��8z���%�#�ڭ4a���+Eޗ�ƛ�l��g��J�g��F�r�w�%r����a{L�V�lp,��D��<.��e�����I��O��LF�u���f�(�Jg�2X����U��ٺ�[V����<�LL���;��Áz٬�<��+H��|>�؏�ޞ��g�(Q����Gp��<9�s�L�Rcw�[�bc��Z�In�~�NI2�_��7�Ȱ2�̆�l�uT9$�E�l��bY�|�d�x��z��@��0U	�dq�k�Bd�lj��Ӫ��K���5�\fu�������v��6�u݂h�He�#�pn��ؒ����]a��g����vM��4+��;�L��L��Y��%wd��Zۨ֗�H��u��I�hn�j�
���l��I�����4rw�}����Z��?g�`�ϡ��Q5��N6N+�/�::�3��q�ܩ��:qm���v�D��ա;���..ӹ�6鴷.'�;���y��c��?ʡ�e��+{G��lPX�|�5���ժ���R鿅/�V}�j�\�R���,Ⰶ����0h����*K�!IM�
�^`$;wC]�h�}�\�#�B]:�fֈ��Ο�K�V(���Ι�a�v�
[��==ݛۀ� �!HX� ]��m����t��(�PEX�-�-ZsSH�#p�S,���T6�a�<P�����T���^��	���q��(7K�q�Vd��5�qx.�m}g.Z%��Ùnݺ��O�,K�B��.�j�W�O�r!uG�]gVfbM��(*ȩ����-}/�`w2�P��٦�ؗ�&`�M���'��{�˧���_�v��eC��FS�1��Å�Ɋ�����X������no=O8��d�3��]�9�����zR�hË�8�r�j\/^R��� ����v�I�2��\��T���𥢉rj�z�ծf��fx����5q��n��]ѭU�����is$���I:�#��^��8���]xI����G{-#^"d���@hEӽӝ�6`t���V*D��P��,��ge:��������a3�xf�_��X�`�p�U�/�A��k�I(�?r{�����/��ma���5S#�<�VM�����A	�k򣻛�������T�f�g5�ʇ�+��K��ꅛ]xYE�`���=ꚹ'����.��ls��p}���C�X����W[�������3c�ƣ�a�M�@DkB��R����*�*�����g���4}� ����d�Y�|;���Ih"� 4��,�j1o�+�5?a:Vǀ�"�Xtjxx���x��fQ�s(kV�L��=m��||`*͉D���Yd��vk>�ɵ�a��Σr�#���ťZ�x�&๽�J7��I�m��|�+4�~�����Y|đx
��K|��fao>���Vac̏{U�ǝ�2��X�{��2�F�P1�0��C�+^�ɗ1�'�-�1����M��"n��u�^+�����D��.�ʬDE�%�����f	y����ԋ��r����F�@��ʄaj�՗)�v�:o���k,�IXӞͯ_|g����	~���kJ���Va��w����9����("��������	����ԍ�~�nI�~�,;�׽:��^x���j���#l�6�?�ih���y�}�{H�uH����/�H��Y��k��<;����t�`T(�A�nD1Of;�L����R::[>��}�~<y�>g��E�<$�<�{Ә�hC]C�>�r�u;⏝d���ϻ���N��B�9�F{;��雌j�(�  ����XWP���~XȵyT��}���t��!�7��MS4PT0;J�u���QŢ�x$p?P�����'����=M<_-�7J�v샆�u���CP���(	����y�έ��v8d�S�w�`�:���6��+���%H��]��㐤�,u;A���eJ(��0�w��9^���0e�����m���w떎鯹o�,�x�<x�.S>7u���0��["��V�V7(��#�>��묥�~y��G�S����4S6a�V.�Y�P=(2J,���Uw�*ݥ��o.+�d���W��D!��n��v(0Q.�H�7DI�aId�2o�z��#���`tK�M�d!72�,g���c��ܣ�[�/L�;ǀ�݃�z�̂c�XՉil�(a��
��ӄ1P�T|�ӗ;u�\uc2<G[P�TF�͑�V*��4�h�[��q;���yyr����r��Ucʦ�ߤ�4p��3�ᱵ�7T)��o��1yQ>ME�g��bܲ��A߯K�_�T߂ge������]9U�)���1���y�ɚ4`(�;�ʝR�)����M��%�����\�-���Y��d�mu`Żh_L�C��� L���j���L�d=���}A�U�ԣJ��I���<�i����9�r�T�{���S��w�)T�"�Eڸ�\�a�3����M��Ԗ�x',$o����-}��޳�4�$����q�8�<|F΁p�j3�M��i}t�5ϯ��_Ӻ� ��?ea���Q�kK�cڵp�2IB�S���\��-������TM�j��D #�G�2�v���v���K"Ik�ڡK:I��{^]d���:[jc��H��;�kFWAd�2�u٥;C�^�+�
�="mM�(,��f���f�������)(d�$������T��U݊�=/Tې���s_>=�,VoQ�[��������K�V�������FU��&��1��N�Y����s騝=��T��W+��m&z�\���te���HV���Գ0����$�GW�;�g�:��sy�[�9IM�83[ϑ���{{U�C[Д�.v��nuM}�`U^�h;e�w������X$)Wz�,]�a8L{��}SV������Ϻ1���LJ����Ш���Y ��jb�{q22=�C�H��xp�t��yʶ�8/��	%OU�j�n[N�Պ6�U>uu��#���9���7���w;��j�+��L1�J��	�x�KU�L�"�j�W�Sr�Ղh��d cP%�g)���t�* h��m�����g>�8Y�2��BH�U:��U�Ҿ4:�����LY]POo6�ݘs�R��J�,�+ˎH��4͉��������9���lX���4*��n�:x6�ѷl9���է��42�*�\��b.����l�F���������층s"z�� �!-�6�=�n��c�ob%�7���ز-�zpoh�n�ŷx8��ۙל��Р�E�ӹ�t\6c��+w.�<�@��+�q��/�g2�l<-P�ej��l� Ⱥ+�p57w�,>�n����w���z���G��,��\_��zӍ̮�Jш-2jZ�y��_t���̾]b
������YE��bG'���\�d6�3��n�����S3Z���E�e�V�mP5�5�V��5Z�j�m�Am�ګ���m��,R-j-V��m�J�Z�R���EJ֨����T��,UB�V�j���ZJ�J�QJ������)m�h����lF��V�J�De�T**�+R��--B��,V(�6�[H�1h�R�j��¢Z
�Q*��V�F�RՅX����ҥ�6���mAcl�J��Q-b���D����eaim*�Kkh��B�j5�6�h �Q����Jڅ���EKK*U[e��Q*�V�[XVU�-`X��eb1�jB��h�m"%h�F� �� �DJ1�
�gOZ7�Y�s�Za�b������Q�_w$!�\�k��u�V5�o�)l�ɱn����g7yQ�P�dd���R蛕��*Mq��U�אc��X��4=׳Q�P䖈䭖��,/�f���/v�V�4գ�@��0mؗ�]�Ɨ\�6���=�N�Y���uݭ���Ӹ�p�X5d��t/�@i��Q�f�X���:[���Ӄ��z��w�/ �hd�qP�t;�m}A�_��Z2���G?VW���q�x����Μ���~�V���*�_�u5E��	흝�89���~�]|,A���m=uEV�ޅN�.��Y΢��1�#����Lq	
uB���2��L�1�g=_ICբ�#t��!��cݻ0%�O�z��4�!��@E ���}|�W���E���sX=:k��20XN���n��a���P�"�4�����T�k×r�ג���������D��,Xn�V �ԫ9!�/MC�0s����X9�vm���ݑv�P�e{�i塘�>8�����C��d�����tr�0�E(+�����*Y3[�	�Q-��KҴ_�M�s��������)]�W.#C)?o�d�jP��@H��q��='ޢr�*ȧ�~�����f;�Y(a�#�i���1�y�M.Ny�,����ײ���U0~�P��Z2���4
��J��noZ��qs�ʰ�]�3]�+�����]� ��A`��P��R�h�{�ЬJ���ɨ�՚t���K��G]xs�,�����m�j-�p��ۻIs�·�.�cx��:��;�C�y_71ܽ����=��T�5z?zv�D����c���Dx`�-:��'D�h�V�*�����)V�#��홽lا�1�֠W��0��(O�kr���z����ﮅ8����|o��~n��;���Q�5�s}o��槹�ju�B�`��5��<�^pl�s�S@A�!.��"yQ��և�+b����6l�����.��0�7����;�t�zi*W��i��%1	F-[����u�;TP����f����J�����C����y�s��-އ��
srl�X]͝�"�Գ�������ຌ%|��ւxєlGkE�a�ߦ���B���.��+r�rd4p.�Σ��h"�Pb�����������N�|��`���ӎ�V1P�VD�^�K(䍧};��r�>�>,�4w��N�d��vk"�l?k("]MS����Ӧ���X��Y�00��u���h�R����K��k�ޙ5���uFl�!��_]���̄`��@��:�j�U�+��<;��ně�n���͙�9�L���ʯJ��ȼ�0OP`��(EU-���۵�׮v�▨z�t��ު�݂�KDϼ\0i,!���'��v�d\ �tN��k���u��k��vj贍-�\�z��53Z�=-���U�Y�3�0��t7Io.�T���_V��0��n�ØM�l2S��t렐�:6�Y��NB���H�V^��5��[J�,]ر�;�緎��Q��\����kPʾ�vH|yB{L�ѫ�{ʸ�fw���9��sL��W���g�|�^�g�O�Ƙ��N\&��y���ԭ�4�3Ă��ǁ�~�j�v��(����XY�d)�8U%�L�M������������P�,� *&ib#�+���*��3s=�<�\�H��mx�6X�̺������Ҷ]i����ֈ��ܪz��b�:����Ux�$��>�,��σ�T�jR8��Xg��T������@�̓��#������"��D�]��/�9�ϒ����FN=T�qh|FWG��p�U%QU
E��"M�l׳6׺۬AS3|ԓ�:p�t��7��[#҃66�ժ��
%�5f�˭%�9ljkG����ֈ����lyh|xR�o��Պ���s�U����q�L��UI�^�AX��LcI��ǆi]F$=F�cϗ?IV��B��ыkyj���k��z����\�c����'*C"S-�(Юq���*l�!iV�|��>�� �W���mj��<���ns�:���4��.����N\F�*m�w��-�)T;��#c�gA�N�5A�������w=�rݭ%z��bV��Se�Ǝ������̹DU�5^�N��X�Pu3c:���+��+f}Am���(z����^;Lx��M�ʆ�˷M���9�e�X�U%P̖�����{~+��ʄ�^����sMϖ��D��V�e��P
혎y\;%�	�n��+��&x`�R�91��l���
�lϪ�$�=k�L�%")VTjgy$��}���+�����aU���%A\<O	|���.E�[ޛ�w���V �D�`|tM5�t�&����/��#*�w=����`�u~��w����Z0:�	���FU}��Vb��*��_P�/w��퉿"5���E�yx+8<���4�*��^�D����(�bp��q����M�:���<�v��U\�Q�d���xTs��/s�J�3i�ni}��U*Ƣ[�F�j��ꐉvLˊ�NR����[���3�b՜�u��W�FoanWrm�9M��
G_X�j���P��l�x}����%����.v�0[��l����9�7nٯ;7Bȱc_�� iZ�����r��=�~�w�� ����i�M�A�U����Ꙇ��as�Ǝ�v6���q�Ю�9{�k��b�:E}�,\�co/��"u���%N���&5�y��y�uV6���ZaC]�a]�V%��v�bW�D.��=~})�IK��;n�^0]:�����p�g���"�;�M�x�sQ�?uI�w�ښ{i{�J���e���Z[B����Q��L�;��U[��]>��qZD�鬓<[�G�u�zݙ>ܶϊ���JN���{¬z'�%��ٓ�j>�b_��p1Zl.�$�fAAd�B�����~�&�|������X��D㢩}�:�T�4���%����(���~����Bۆ�;�@��n����/Ӷ���$�S�j�L��ֲ�!����=�Sڝ^�[��>��ϠƌQSkk&n[@��O;.um�_�ir}3�8]����l��ޙe��+�ܜ�x�ac�Ja߾+@�m��0u��+UK��肰��`�^߶o�dU�\]��5�CR��u��g�;P+�8n@��v����ױ�~h�+���2W����/eC�>����̿d&9�N��ܞ6��x�V�+�(�GǸ�UCz%�o��z�V[����1w��"�'J|��f:k��Ut��.�èBm
�C��+)P��ɓ5{���8Ap�W�TԱ�ʨ���W��8 ���3.Ѣ(��|��yU-oE��
:`�'�����!_wXTkV갳A
�v���{1$�k��e
�X��(��Vo���@��It���'p�uJ�i�@:C9�}�T�p�I�g�� vEƍ�r�����9����&,�e{tGz���f䱹����@�keM4��skƕJW�������92�]�Q���N���C�6��jc���r�vKy���|�%�r�]z�%�V(���8�x����7�#t�N��}(r���I{�ķe�=O˅��&���pu�hO�2/-�'�0t���w;c�0�7uG��{+@}�+>�4��+=~*��τ�2wɕ:�g\��e�L��N�p9Zk��<�:5᷊��]]�]��E�r�f-�L��r,��Ŀ��5���g���7I\u�L�2���%9��0/�F��k�G��/�����G����k4}���=m�'�]���(�G� :~U�˺Ư���~7<�..9���am����X�=�`0ׇP�� ��×��U�
�/��{o��w=����<��mm�[[�G��\n���~�Š��n'�]��h����`�|�[��fK�C�V%U�L�]U:��5i�P����w���z���6 ��Q&]�bU�IS"��V�*±�#L�q�������V�t�w=�}��*�U5�{�@-�s;^*NѼ_Nf��L޿gD3�ޒU����C��B�[[�#��v�as�B�C��61���p��N[lE��s0��p�Yח�Z��\��:�*t|�$�?�PD��7ԭK�춗�ׁ������N�!��F	A�&��
sEm�=�p��n��P[tY��p �u�U���VO�e�//L��^��-�j��TmWUX��4|p�C�z{n��C����=|W��^].[�h8p� ����s�
ڇr�4;(����c�x��/|�^���IָA�b�{8��BjR3�X�	\��|h��>�Vw���~��B��N�����W�x-�w]�����_����y�&�|g
�,ḋE՛0�2;�+�^�p�����ml+z�n���\��c�;%
��Ϯ���/���hv}���p��[���@�CZ�H���>�lº�7hԖ�*����Mz4�@vZ3xڢ}F���s
�s�V��.�2dz	-m��a��3Yz�5�#&/�g{j�$b}��3��e����˚XzN��x�	r���'x���қ���� s���iNzv&9nӛ2��r�������,�V=T�>�\�V�۶a
y���e�n9��!��]YG�w�o��p*)TO������cl��l�]�{'9��<H�����x_�StJZգ��)I���Ы�A���pgt��\������t�iT8�÷^0���3�#ƈ/�^��~����6 ��n����u*^e#c%�3�=l�ޯ�Ic���I�5�7���M�%�9F�jݛ�g��vL����Տ���J�g��<�I���D�ag���7�f7�b����"ȳ�=|h�IeӐ{���z�7�n�ܾ=�zšP�7�X�)�X�ԫ8$7F��p�Ů����~{�53�tH�:���ÃkK(h}��Qb\f��z�c�4k;��q�}�y�f}��|?�UwE
l��EÝyA��2��C<	�v֯��Yy��ױ!٠)��zl��V9�ݴ��Vd[�7S���7�@�x���`IEX�'w�+r�W�����Y�+����P�RT�͹Yp���А��vOGRhH,Ļp$��M�$T�OU4z�f�VeRC�pӢe(#�-elv��z�j	�붺�į(�w��B"�5۽��D"�]e�o)-ޡ���S�':�:hY�sY}إ�tk�V��v��U��7N��ٚ�jM�ZҖ�5$,s|�<˺};&��߃�$�lZ����J���'��L
�{C:୮3���q1�&X�y5J�2�B�R�ooFY5v����� ��v��x�k�j76={}c��6P�Մ�p�l�I���/6k"�a�ӿG�o�zOn�ǜ�#�m�����5p�#�n��;u� ���u�ற��lJy�X�ȴ	�(��rS5D�i;Lmu-��&L�֨���{@n�i��o[i�[mwA6������6.v����I`�=�`���T����~tX��m���(��A#mv�Q��:��9�INj�WW!���{]�q��l������Sf��*�jV�V�y�(�&Ŭl*��ܮH	"v#�Fe@[8ݫN�×3�f
wJ:q$�V$�)�W�� 8�>Q�ZE�+.�<�EL�e浤C0cu�e:���Y,��V��Ѻb�t,\l����Q6�R(��ۋ�JY�F��Z��*śh�K.��e���͹�+j��_>Il�?\�F�S*^^�Nڴ��3wg��(ѥ��mP��y�Q��l^H�חtuQX�U0e\��t<f$�i��k V�fV���n�1�=���	�f���p"~Ȱ��z2�˻�n���1K�[W��]�c4��
��wK��ݮ��L��bX5X]�^F�F]�?3eM��1���N>����<��	;�`����C`�tּUw6�v�Y�N؜7�l!^�'cBg=���˦�l�N�r�5�նy	�[�k��dt�
�phjx$�� �ܚ��f�v荶�v��}ڲ���x֍��8�l\�[|$�9�}u����v	$SRlL�5����;|��@|E(���dX(���6�-k,�V���*V�ږ��j4�j֔h�D�P�H���ԵV�+PT�@��B�F�`���+j�[(���h��dP*5�V�kPm(őb�Ԣ��Z�b�B��R�����,V�ZEm��Z%��P��il�U�c-�m�"V	U�Ye�J ����cR�""-J�j��TB�*�Ph0�
��J��-�(��U��
�XU��Ҭ��m���Z�`�+m�R�V�ص[lA��bU�@��1n�jr�%�\�Xy�[��*��ޅ�7�9p��<!�V��9��R���q��$I����ok΢�t^��_��I�6�:�/�h�k��;AQB�����.r�Vt�+�6��	���;$Vu�z.�܃�`�Jż��wo��y�삻�����)`~��e#oV	{��q
�k��R����-�
|���\�
�~��pr��J Pw�6����{	�u�Y/=��QGʸ���W����^���#�D�'DǛˏj���=�Ω(x���ʏ���|x{�h�O�I�<}�`,��f=�}I%��5��3~U�B���8�:'�|����g���m��H��o)Jϊ�C,�; �B��q��0��)�/��g�������W�+�Gv.��6/��tK,1]UD�#GjX�ZtA�ϛ~{���3���a�UR�����\�z1�4r�p1\f]�D;�s�b�B,cX���T�1�綱�k�����e��S2nJ�f���FB��V�+ǻ�(�֛d���W�C����IftAg(^�gu���S �ʕl�]3A�MR\�˛[սe��fʄ���L7�:
P>b�G�0qPtj:�LU5���s_��\�ʠ�t*��6aGA��D���L�-#n�_�����ff/I5=C�J�]fԔ,�f��:�68mY��.3��=����_Ox��'�0}U��K"�_�x/ySum�S��а�|�!���>��ӗV�o*�GhÅ�1P¼)���W�ζE层{�%�[�\�hh:F�>�����M�{+C��Y,i<,g��z��l9Aŭ8�i���'Jt�����(CAg`wZ���W��I���KΞ�L�����Â1h�_������;Ls��8@��Ew݌Ki����y�OR�¡De���൫�Fq�8x��~<_h��X�^��K�L���e2��
P`�������������qͅ��$:oP��;��m<���RA�<��WOݦ��7��5��sU���,�;R1b>=���D��bTk���1����G{�໤�8g�k{N�Y���6Ip��nd������ٲᰬe<���O 0k1��y��^��.xU�=Q��>#�L�XAN��u��0*:�q��A�����'l�M��L���wL�T,�Y�۫4<"�*��e��Zks2���/�w�ޖ`G��֨��j
��9�tx��W
 ӠZH���ۯ7�{۾ry��O��Y�U*��e���P�gMX�f�@�GO��}�'��I��� ��s���a;��_e�
�zA�U����ҋ|`��7N�ж賝���ź�П.�m�h׸T��.�9�̿#b�e%Tt�*�5�,�F͏��2$�]yS6T7�*x�w��������;�x/��-�w+@��Ur����fH�[7ǵ��lYr�~ܱk����=+Ϲ^U6^�/��Ϊɦ�g����A��w���ރ���6���&뮕8�8ZV���G#�`�̱V�M�:']��=��Ʊ����:D܆mQ����][;&k5�/�hI�\��ێS����M�
�Vо�������+-���v��&U5��t�7)�f��>�a}^�'�� �B�>~_ܮUg+�Jf^�Q+�C���x�Md���S�_�WQt������U��l2N�ه�\�3����+v�p�q��2�
R���]�yvG����D�jn5�D#�ץ�uPJv#������R�����-�-�#� ��������F�fTO�����|o|���u^H��2��Ӳ��M�uh�.�-O���S�Pb֭�����[z+gC��3Z���"}�P�V�/�8�p�0�]u�v̊����>�|��z�ud64+ �h��!�4�t*~\)�b����Ъ�n��s����A�]|T���|��B��� = ը���>�L8����^:�sGYq�]�R�&k�oOi5Z̻�{�㻄/(J�y��)�g��t#�Z��7׉��q�+8:/%v�e[D��p��y�mɫg:kL�9)X�6��6e����׀��
J�[7��,P6A����:�>���%E'��[���+���d��b��p���Y�Ѱ�߇g����OSi�����'����Qp��xpmi�	A�y�T�T<��]��}Q�C�������D���3+o�V�C����{/�c������2�1d��#Ǐ�o��3��l>�r��Y�b��0�u�)��X�7��dJw.V:,wr�^��^���ჲ���9��3�U�[�O�;u�*�m8%�/L㲑���{��+M��$�g����N�5��zY"mt5��ʺ���н�©��*UͰ}[R'y��Ux��ld�U�,���Ƿ�B���P��e�]>��^�Q�s�P��n׍J��.�7��*%��p��Z��SN�o�E;�{����8��0zr�ܮk0��:ʊ���Υ�0����]J˻�)���:V��|���\�8�=uq"��}]92j���;(U��f�����V�0��:�sL�nB|k<~�I�&q�����_zX��c�C������J��s4�,�; �B�|{�����B�:�b������3'�|ݪ���Y��T�N|-\8m'�� �c�z��o�[X5��I�^�u깏!���r
�*/K=ٞrL�|h�tH�eφ�,�v��0<4)P����S ʂ��%OG/ʆ��2��B�g�X6YG;���½HY$N�YsC��+"��{���6�����Z"�yRf�/��i�8m8���ڇs=�D���U`�k!V�"��������#��0f�H�$�n���[��)]i�%Ò���~�Ɯ��B�����]��}��f�O�#��:X�pz������J�^}�+%��YJ�Ńg=�^�� �n�	nc��/2\��Z��)>�
%������+w�Gj��m�/%��s��[W���2����%IJX -My����zV�JK�h�w���Rl��ѵ��]r^y�,��n�<a'�F�����<'�yuȽr�5ݥ;���>�!�48�7Դ?����Hn=�x^�2u!�7���?R����,��uǆ��L辙ʇ:P'�[=��g��XκUA�tU(A���r�v��(�K�^{��x�ű�;��=~"�������|k���d��F�̃�<}w��Ow������7�X��0�p5}��K��?���ÍD�G���{���w�{�R;d�<2j��o��Lu�u�_Q�ML>�#���x�!t��\�ý�5���o�8�b�Kɘ�,��@������ֽOy�8�Z|e��X2X�]���=B�T6Y�Wv;�{�W9%L�IKh�:C$�J�1v8����ΐ�Y�dxJ�Ѻ z� �J�8c�3���rUm�3	�0,\B�l��7�|�)e\�]��tm&���'W��=V�	#K��`�/l�1�r^*=Z���;�����nܘ�O�c��E{A�溞(ko��efx�)X�m��G��_n:x��r�<�jd��lTx���n���n�9�~9U�rZ8�=13Z����*���,K�T�!P��Wh^ڈ"P����D��%m"�y��x�����~S�z�Nǥ��K�n[,��w*.�|)�o^�w�Z�v�rf�[R�gV�nX�녉�!%|�}V/��[�ƎE;u�+<���}B������#n���1_����Pʓ>[L�ě5y�k\��Ph�`=��WQb�%��'��
�\�8�ʮu��)h�Os���Ó���L�)+��X�vN�UlV]q� ���U�7�z֬&�*�a���襺�C�]v�r�Ш,uw�We�t�\��כ^�)�G����>R���}�c���5�+��A�:
��h޼��{�s6;Ԗ�|� D����1Z����Z��0�WWO'�S0.D���m$Ѹ4���}��9b[v���]��߶�'�.�c��
�lQ��O���z�L�=��|�J�J�M�M��������"�W��#�PT�pk�pjV)��������}4���#��.Z�v��T*8����4+���֮t<���!�6��#ǜ��Y����%�z]S��4EE�h�W�kC�	u+���;���S��p��I���'��?���.\rҡHX�I�h�0{��TSu�S��Y�V�z���`����7�[0ѿ��l!XC�����;�n]��kTw���X,���3���Ut;���|P~��M�)���=O����:<ҧe�`�ZKLX�+�*Tf�"�ڮY��(�}�\��j!u��R?�LNվ��\�``ؓSm7)�ڛ,i��Y��OQ0���eg���.�?l�}�=C;m��8�^�^�7�	}g�{:�`�m��Ծ7�GޥPp徜��k5�o �X�������_6iFL��-�[^do���|�&�Sk��k���N��s`	mK]��_]�0�#�yK��Zz��B���m�(G�Kǜo|绍����I��}��CҞ�E����H����.�q@�K��l���n�ޥ��䣙����1Y#�m�^!俼{���u>���X�^��L�:��8�]x�W��̖�{�/� �������etU��F�(�ǔ��5�sܷj��UM�t_Z9�3�Jf^.U�b3��!Yr�E�zأ�n��thW�X�0'½�B�<�\Z-�~>��O�������W�xC�|Qf��0I|{��a�� l��8��̓L�_�ϱ��Dz��*3WZ��.��uJF��1�yB��Q���:eu��{m�R�U`�b��yR�~w��4��L����A�ܻF��tH��S7�~�aϝ_y��v�<�|o�5����d�Q຋������x�PC�C�Vo��~�
�[�@�{���p{p0�mKR����[��|*^θI�U���淸6VHX�z��I�:�f?�X��Q�Z�p��nO�S;��+0&vkd��Os6L\��R�ʬ�ٻ.�Ee��\Ե*�M�W�
�@ތ���g@����2���e��bu5ܮ�+���6aպK��SGS�[��x1��`Jty}.	�Dą����겤�4պ�����i����O�I޳W��N�	�"�4x)	���q��@{��7Am8c���vn����0K�]�:��y����#&kc�5�/�E,���W�������ӹϊƷW=��o��g�x�lR��d��*�8 ��m�ݦ���qս�&͋��U�>0��j��r��Ҧ��q�'��N�0!�4m�G������N1�q�ڰJ{�i���z�L_��A�sA����V�'w�V��2�^�r6�����N�c��@,uX�/
u�k����=+�C�h:F�����5��K���f�&�Ӛ�juQFb.�d;�%ы���*se)�o)n�����u\w)����:VPP�N����81�q!��,�c��)fC�e7a�2՜	)Vq,啕F��]Z�5�I�0�G�V��T�N���+.��D&�0wM�٠���"��ٛ��#���KwF��fHlږXf(�� �1��9�a�wn�j�ƸJ���RΎڷ;���`Sgl�ުYۦCe�Z�=�[F�κ�e��7	)P��i$ض�U�N͙;���U�B*�"�7q� ʏ��`rM�;�G����g��xu��{o����	�4{�/k�B�-3L��E�]^ͧ��N�5�t�(b���%Sz�ee�sZ���4�p�bc����#]cN����qv��zI�]>��x�%-��z֝ۑ�3��3��(L��*��s�֦����9���w	�d����H�b�d5+�9j���a�.}�w��_0zD�&u]�ۑ���v�/����nͤ����4*��jQ ��b!D���Q�Te���ڊ)�Z���IX��U*�bUkT��5�V��Ԗ�VZ�ijDb��J��T�h�b�EAQ+[J"TF�QTKj�Fэ-�*ED�YZ�J�b�b��1�ej[,*��[mAJ�(�,��e�b��IU�aX(6��YF�+m*4m�KQE
����+iZ%J����6VQU���
ђڤDU
ʔQ�*�(U��h����TZ�DmlZƍ��B��+*��"��F%�T�ѫm�V��h��RҊ*�h"�	iF�,T$�7{9�<����Z$tV����D�v�W�]��$��Q\�
�H�[��nP�����ޱ2�b�0k������t}���L��6���>�����^�r��b;UY�v4�E�V�*Y�����V��������dǙ�x����S�Z�ugC�	ZY�4�(��0cΟ��yw�v<+՛yN�C]A3Î*�XtA�gL�7��i���^R�R�m�7����v����['\$��-�ߝ��o��ao`wK�d����o?4�>���4.�T5������UhT0�wǶ�%{���l�s���]X���^�e
��(]y�b���r��.����o����)K�=Î�F��h�
eϮ�
�`��ܫ��uR-�~����SR)�w�ꝋڄ)�G�5p�
��b�.r��N���g����y_Jx�w���Y�����24�u�[K�J�h��>����}���Y�-�^D�r0���ת��7��|���5+;S��&fC�xN0�u���B�`���R����.�!�g��6��v��丹L��8���޵��mm�5�:__V�2����D��9L��P���-T�ٳo���M�K�'����s�W�p�8*�F�4Q�]��Rv9]���	�%VCz�����N>�0��t��V��F�3Z0*F�:KB��^1^��:��:�r�����`�X6]�a:����qp��a���C�
�=X����M�]����e�00�M�K��K���ZC�o**���77�}T�O<�[*�ˣWC�d��R6�Ӫ�
�$xekP2X�t�r��Ts;y)�n�D��q�VXB����]̪r^z��r��^.�o�oP$A���~�t�GCM��l������`��R�^�1�a[P�*#B1�Jv��o�k0��ZPh�#�K"���(8u�Py�T���l�����R'ܻ�]��k�~ڣ����xO\0�;�V�� ��V�%+��=�{"�4{��;ŏz��<o��+�U�.��!�;���$�}v�3_yY��e��ꂝ����{������}������;}>���.�b�l�w�pjd���]��u�2���m>�a7�8�l���fկ�-��r���M��b��-��]"U�s��Z�oq�i��u�V��g<�[V�3�5h��G��B��0a���ߌ��ޝ%b�]���pa��G%yP�XΌw��T@\׻<*;�Ə�2�U���~Z9.�wXQz+C>���z�3���vOxK�1��x�.�K�E�5|K�%î��W�=x|pv�m|�)&ǲ�o�M�5��7^5»�OH�iR��$��~>�P�b&ǜ8W�M����I���q�͑\����B�V��iR<btΆ�yp����G���O��є����Nǫ*�]�G:f�f���t)����u9N׬����w:�χ��[�	��`��6ٸn��l�F���A;��I�1����bZ4lg�[˅﬛b�:$W��b;�{I�D�7�h�I��Mlh�S*I|�ϲ��'^��of�v�ő��O����G4�8���kI�}N��Ck�ӫ�!*#6�p�r�W�t�7;Tul2��Y���y Wk�y�^|�w'�I��%�oS7Fl7	\fZ�f�1?.�b��c�W:(�tӇ#��^��RδhN��y%�zj}���~�i89����;G��p.��ʹC
>?f�ذL�&�x]vWJ�.�"��Aɻ���)oh1��ez��w8$�#$��6�L�/k��J���R
*IS۞��o���1(U�#P�J�,F�q�z�K��|x�΁��=z+}��D��"���z#��D��ٯz��z�t���}L�U�^ˋ9���*u*L-�ci�Z<-�p�����Lp���y��-�-��9f��w�����j��EЯb�m:��\:���z)>LO�<Tm��ywAW
���T��Z>�*����<��xߏ�T�|�͚|�������a��a�vA��H��#YT&p�jy�b^���Ι�4I�����4t�Τ�����h�`¯($.1�-\K�<'�[S�<556J���\)v����6�����F�;3��X��d�� \�-Òeu���};��B]ex�|��
�j�x����x�
spf�q��yNDw�@�1R��c���<j�݋��IV<���ӗ�I��h�)��]�D]��`�F��ch�nt�c~��2�J��jf;/�����AaC��ԗ�������ч����UY�D�y�p5�ݷվo�J~�lI��Uw*p:�*�o�k�K�ePUD,~�Gm���6ɖ�3FF}�
�^�D戥�A�'���U5�k�t����O�J��U1�4��\ʳ�>^,pa��D1r���Y�#s��tw�mTW��uz�����u��+��*�D�a n�U��ƹ)�����m�8:�����I[4Ȟ��������;�w��z2�R��ӷٚ�D}�]_��gC���]B��Ur���c$�o4n��ʽ�̅��V!j��,��[�Uo���\7����0+� ��j{o|�q�ϟ%o` v�B����n��aJ��n��d����N<���i��V^���G��������Y-kx����#Cg���{����{�:8?���#t�Tj�Q@�����j�T�J�پ�[�3.5��y�_��Z��疇9h.��R�/�*��ܼU`X7��֋�}��<��yn^Uq�V�A���2��M�3B�F�؆خ�K���\���s����}H�����h��X<�4z�f�n��CP�B}P��mn)�/w)�/��2�qr������GE��o�R�[ภk�wִ�f�=��R2�?x� �B�uY� ���肦���R=ؗ�z$}a߅GL���7�c�y ��
���/j�Zƕ!!kzs��	5<��G %-\�*��pִ���TU��G���3$��WO{�Sǂ�l�b�4G��N�ϣg!��W�h�G@X�}YNT�����fysy�jyg��vΚ,pv����eW��y�YF�����ݭ)?&^�W��<>�k�*�*���KTE�C1VywtP���bH���tH�m�C�U�c�K�I㳺��V��1�!�$�æ9C/QA�(dF����2Ɯ�T6^1[��d����c&Ƴ�,��ǹ>��[�V�0|��KS�mR�b���c�{�y:�3��_n��=�A O�>	~���)���ߝ�5xx�4��D}��y.�Α&�C��U�lM�k��V���!�uf�z�Ɍ-��a�0�'�I�7j��3D�f~#���^V���u��n+�$h�yo�{f�ty;�&kC>�Ƅ���U��٢b"�V��*�ݳy7�����`�����<������ͻ"��-_��G%)Ŏ���D�~�Gގ)���PT��m/|�E�m1�~��6^చ�S}��b^��R�ߪ|+VҔI<�7���LW���Ԫ-��y�K�?��p�@ˇ���dw®��Մ�:�6<�-�< �����#��	�u��H�\�+�i�sw�Ы��Ө:!�+j��.�
�}�hq\��E�8�/��ʂ��Pv$(��l��ֹ+{o^+����iN{�(9&R��CՋ8z��)Ҝ�*Qp"���C�8�ܤqJ�Ӯ92t�zݽ�&u�����r� ��	����:z��#��
cũ��k]׉>�\��4K��5}p����7RP'�Ph�׷�[0��OOZ�y'=ɾΨ�PB�Rܴ�*귁����#|ŋ��Y9�{f�ԣԕ:��Ѻ7��p\eP���d�qm�϶��ƻ%�7q3<9aȦ��3�Tq��:�����gިU���I�8f% ���T�[�6��c�a�%���0���M�bxP��vC�]vWJ�����ף�gcT]��.u�� 1W��V���c�|rK�0?{<n+��d����PL�b��s�뾣�,B�VT���*��F����\l=x%�wǎ����O�sS�^�=��R<pH-e������&���\�(u5[���OÏ�svL:��0��kbE�֘|>#�h�2e��[]���E}��|a*h�v��,���;Ju()Kq��N�&���έ�u��ǝ�p܊��1h�.��VK��X�拒����6�a�VX�]��l�v度�,޻�7�X��[B�?���*�E{�/��V'�=��	�eq�Hє<�Pk����fh�gHY�I���6ru�\E�����Z�?J�'4�KGj}8^���{�?z�̯!z��T,َ��PՇdm�'�)X�%/{wg>q��@U�pnv#�O�>�qdN�F���Ѧ��۟@��"�Y�򺮉��z��{>4�bP���+>�R����UX	Uϒ�*�z���lt��;|�%��A��"�yLhu�`L����a�Ꙏ�����rR��<A�&WR^��>���TW�`��gÃ�(]}�L�i��}&i�ֶ����4��l$�:�Uf��aױw�]�|ռuެ3��,�}l�_{���{���l��K"�ZO��r9g���="g-�.��Q��&,:���~_;��6,��$nc�8!W���˗�7%��1�k���G˄�IZR���̓h�oVV��	\gQH@����n��l�v�*�t��^ʆ ��u�֝j�$��}�z�Hwv��eA�P��K�-K��,�Ȯ�����Ǚ{�V���s5׼`�FJGO����0s�*�J
�
���}�*��e��.Jjc����6t>�o��byþ���56�������2yG^��UV��^�>���^l�;�y��)Ϧ;��;ͨ#u�X͔�_���<.����})6f����||��4R��F��u\2��8�h����%�oL��%���Y]�o�ɴ�����ו�=�0���ԗ���;����v�[��3�ƭ`�+�����8�����4pɘS��-iI��k]�@g�glm�l�ʷ��tl|�ņ��6�gO��ۼ7���:ե��M�X�_o�0�����Ց����Y�R1t﫬��:��x:�#XU�� �SH���G��G���\�O,,�+[.ޡl3kZ�V�Q~�g}^��t<��@@f���F,b0ڎɳV��r�#���q��_r�� ��.IRbv*�s#XTD�vA>^�wԎQN�ڿT�"7C�;"�̧4��73 )>����-!s��J��
�,�'�t�u�lC.vdu�h8��&T�2T��mr����tuؽd��z�R��WB�fH�21�6e*������s
���K��R-�C��\�nՂ���ߧm!MU�oXo����w�;d[!�Pk�g��K��SΧ�S9�o]�G��X�.�N��B�'L�ۣ��S�E���[��ѿg::���{O1t�=
�j"��7�\�b�MkY��3d<��O;6�Ǒ�˻��$�ҡ�biT�W��й�1���э��{OP�-Q��$�`ު�;�,���d,����p�37�����}���T\��/7ծ�׻1�/Q]��q[�1!�WC��P�t3�
��M0�)u<�Y��XO��}뚕�4�W|W����5�e�6�T&K��h i�NRՕ�n�<����۩du����R^���z�wSܛ.�(-N��R��r@LRgV�z�5�F
��7b�پ;vS}�~ٛsxS�V�4�f�X%�PP�	7t����z�;�C�+L��(�b�j.WҸRWq)��j�y[ ��1̗�`WT��|"�Q�+i��7$i�Y5gr���Qܢܒ���p�����Y�Ë�V�m]�<�f���Hu��wB]/�8��vU�@c�J�)�cks���tF��j˼���FSe����e� ������T��E�-T��fv�t���n<nŒpY xl�y�m�3�$Bȸ�!J���I��%�)+����7V�'�dg;k9��G$��	-3��7nf|�Q�ku[=n�R���c���M�Q*�&�¬�d�)n>�v79����Gy�G�%]�ô�3L�������]�dɳc¹V�� >��6[J
���QZ�[E�	Rԭ
Z���ڪ�E��\�У�$\�.f�#����FZ�:�dͥ�[WR�+2��-�%�)u5�,Xf*ն��ZQ�U�X����j)M��a�
�ͪ]jje�X��`VV��٘h��ʆ�j;mln��f+�� d�Ȍ�d�L��ɵ��«R�-�� �eTZԋ2&B�Dd��L���h��b �bֵ��fH��C%a�J�-�R�4j�Ò���ֱv�,���PR�e5�F�ԮUY+�®��wϞx�����魊�rd]�GR�P�E�B��8�gs�X�t�LƉxo9��7[������' ����i�S�V�*Vǌ�uz��:
�M���]��>	�<���^J
�;�N�$>�W��1�*���r�o�5u�I� �$]�o�*�Ԥ���zWG#g���O��K�B8m�*"\�ơJ�?5���S�3{/���Cq���R��q����n��rj)�Y��ߨׅS�����ӽ��M�5���[����.����ں�c��������'��{R�-�����3��o���a�[��>���������r~Ne��m��tv}�|�{\����Y��&��zxDu���o��ƭoG|��}O�CaMji��]2�}粒�u�^�^�5�Py���^�K�^�ǰwh���F�9V�ʇMXb����qLM��Eu���n�:�N��X��֐3l�hH��!ɯ�Y�M0�S�.fkZ�����^Z 4�JWQ3���\��s}�9�Xp������~#D�S��h�Mf{:L�S�Ʋ�{�~���q���!���C��1?���3s��oZ�E�杜�J]t4Nf��!���)�|c�a����<x�Wy�IՂ��|�!��~.�)?s��'����r��C�n����N�2���ao�o�isO܂��BSVsx_F5���,$]Vz����j�r?'fhlW��o#��@;�xZ����N1�<c�s�,�}R�|���,w���ǹ�˼����M�R>v��U"�qM�����2f�
3r�#
*���/ʜ1ـ�<1yn)2�+}׵���Q�.�F���|��-O�:����99���%�i��s�*S�h�gK%Ώ@���)8�y�%-yw)�4�Z%(Cw��!B����a��%:��I<�_�A�����c�#۩�xE��'X=�(朏�f����%��b}��O���#y_��a����x=[�w�J�a��bC��'�	��{�=���љ8aNϟ^���=O�\�cf�Xˑ6{f>^��F�x��ݗ<ӕ���6%��P��p�󱏱B�65���9���k�ȥ�ĝ��ˍՂ�X+�\�ʜ�a��5���\��d���TA�T�ڷ�Y���~�ӊ�E�r�~�Y>=k�Z���9W��j�6���5vK�se�@xbZ&�^�i�E�1u�zK��4A�$�x��۞c�<�һ,�^��E���8@b;T��/d0(�X�~�~:���,r2��KPZ�;,�2��W��1�H9��j�tE�L��x7OÀ�1�VD���$\w`�T�έ���_\IӋ�����BZ�fop�uCn+G�%9ץ�����)_W�e۫�,�x|�Ͷ���MZ��N��A�Rh�n
�gr7�GS��b�J| q"��-.���8�+9�'�#>9���u���P��U��Ãۼ�}�އ+���c���D�<���q�җV㶶m�F�XB.Po���m
����{ynz1����+R��s�I���e�z%�u���[�s�g���:N��#�����m����ʽ���D<�T9���;b���nlx�ʹ��=hg����KfE=���������4�1�r5�)�Qw�l�%J��Vml|e$ۭ��i��Go7gi��sT���ݤ�l������1��2�Lo9�ӴsY|�ܓ�����:�L\�[\�KY,�:�65y:�^�{%I��4o6��b���V^L�~�`��G��Z�� k�ř~���y���}^W������^ε�%�go��h���s�xd>L�N�<���Oγ�Y��O_��#ܢ��k~P:3���*wʯs�a���~�/`�������:*�i�L˵Wx�2I����sv��M�����m��8^��-��������z	�cES�PA�H�6#���������V�D��7.#W�ǛHZth��w]�gأ>�����8˓ޱ�7;���R��4%Ç	�!�^r���e�u�^yyu��n71�e��<�c����=8x��z��*k�{�h���p'��qc#3�1q�B|�'j��Ro��M��֨L3���D��2���uzjݷW�NV� ,i�8��u�y�\�{���N�	&�����s�M}[v5��5���R��S�X�|��Zz�ha���+��w���ư�py�i8Lu��J�����M�x�k� �f����z�?Y\��w������p�u�:.{�d�ɂ�J�
lf�;�����{k��+ۮ�w���I���y�A�2(��ɢ�a�xD��,k��ne����劷ܦ���E�?�CEЎ�˱�zN����z�d�搵�X�/�CI殠Ī���Y����9'x�p߼�򡴜���)ѻ!�����=�3�A��:����L�
��瑁�rZpm]>.ɦLy�]��@�6��Y��-p-�Y�<�K�T�{����o�]�a"��a���'$&�5<�#���$��n �$��=��1B,�&�M��9���;����%>bB+;SD�����ؕ�:���|�N����j��Ś)�ۉxxO��^���6�2)�F0���#Y�;���&����
��q��(^����*FZ�Q��ݺ�S��Gap���y��kt����5*�pG�S�PS�'��^��/_�rg@��Ŋ��Pj�ò{��K���6"��2����|/)�y9�y��ۀV��'cc�k�|��]�ڞp�r��{9(�I�=�u�;2��t��=�2^�&2��s�F)�LI�|�������x�Y�ٸ�I)�1�f�w�){ȵr3WF�\�Z�b�8+y��06]6OYlU��i�d�1�5��m.ެ�Zް�L'���n�[�2Vm��δ�z��Q5��9�qV�_��	�S<����s=�hcwd���8��r^2�RvǨ�>9�^�cD�T�C�(E�˿)�forw����U��sR��cz�̎F�O+}��l�m�!����H{ʩ�	bl����W�<ˎI⣿|i	F�Q��e!ᯫT����P޽W�٪NM�xM�(`�)
V8j,ͷz��`c�=V�l��Ry�<f���cC�Ўb�1z�T�kSyGܥ�Q�9J�^\ʠ¯�����!{����� ���E�N㕵0c�+�{=�s���<��i�(y��П�u�{��� ��-�~���6��~��)t���l�=Q������)������p�R��[�&$��KU����dA���rYtJ�����gɵ�91V�s��D3w�e������6���f-�gn�R^������B<�m�LSW�Q=��g8 3�����bS�`��p8�w3�9G�Qn	e���zw�W�s����(ן�s{�{��J��7�6^V���Tٶ��l69�[H�����!��Ƴ2a�M��5y�����m�0�ă�3�w��<}�$ޒ��.t�S"k=�[^-�����:�~Α���b
��m.7�̚�\�����U����y���|����;�O�vӘ�x'����Z�*�F��oLE�$}WW��n��V���h��?�J����L��:S�'�Q��ᦫ���:�Q�SVN����T�+�2����a�8i�L�FAN�Ny3��H筺�G�V��7T��µO�w�fzz����>�,��/�ܭ�#�j��I�w�A���仕��v��\���٨��+�(��s5(io3���J�����N31Va�2���Lۖ�Y�q��&��qɽ*y��JmH4Sc=�*�t.���˙���=��H��OZ��_;o �B��dp�(r�D��>��E�q*ʃ��꼹���=kb����9cۗ��n�ʘ�8�U������<����X���>�3j��'��pn��K�?eG4D����R��^���NL���z.�����Q��rd�/y��^��QS��]/Wo����ĥ����9זzVovW�)���9�6v\�O� �xjF�o��k<�黹J�MqjE�S���������TXѡ���6����/*u�sVx������"�OJ�|"zrt������?�*%+UUQ��-�!HR$��DE<}�.b������D\<������S���y��R�+�
@�����q��0�B�~�lH���)���P[%�Vq!�ԑDS�@�l���w�xg}���i�)��0��]-n5"� )YTr�\�	�:��ϗ���XPM�9���8�����:��L�W����%�TDE?d��*")��bV�#_������Hۃ�>�$��S���t,�1���DE1��~���D��O#EKv� .��_���Х�3q6�+?�j�=Ժ���	�蘍*s�w� �ә���PA���+�'uO*\�;n ��X=�P�&a��;�&�NP�Ҟ�Kæ����x""��xY�_��m��Wc�>�j���p5>�M`�3M��Q_7�������e��$��ʂ")n�]R@7�ؚ_����~�.VO���4u Hd������_��;H��,���n٥6!п�/���1DSk�@@F8���@|���0P�?�I���C�+� �)`�x�")�~�`�W��,Į�\���2,����7?�K�ʹ��!�� �B7HG���(�"�Bؖr~'�� q�����=j԰O�?�:��^�x4 fS<�X�(�����m���xf�� ��E|�B|���~�8����k5o6�5�m�@|����
��C�_'�\B{Sڡ�7%><6%�"��Q��m���#�3$�s���	�DRWа_�#����� ��v��x44^���"�I}�*P �����o��0������xD{}��2s��i�XA���l�L��H���R��H6�oCS��d�v^x`�TC�l�v��
B�")�0��xG���6�q��Q�^h�HK�v]:��n�	\���J<�K"�H>$�߯b:��?�]��BC^�Ӑ