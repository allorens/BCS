BZh91AY&SY_�`c�G߀pqc���b� ����b(                 `                             iE($����R���J� �Q&��7   �@�3*��td � 4 
X�@�l  X   �
� @  @'� ���Q"��HD�T�
ER�$�
%RU	�*�H��Q%U$!*R�RTR� H%U@HC��T )�@�:$D�*T�%)U����d�-��A��J{�ʐ��R#�vh��N��ѯYP*���TI;�U��3 
 txJ
>�>H�5*��W������P��P;���:<�J;�:������U)�Ͼ���|�Ԕw��� �ͅy��<�J<�>���J>   gХ/����Q!E$D��	ww*�R��˾�́����T}o�{��*�|�_|J��R����g֩�����_}΀��.=�r>>wϨ�>t n���pɥx   ֌z�M>�K\�ɥ��>��
�>>�P��v}=�p�>v�u���z������|�J��d�&V�݁��� ��|�P+�  G w`�V�*��*�(*!D�I![B[�n����J)�;0��zyozR!����� �w�@rhQ�O{: y�⤕�t.�S��   5l{���+�j�P}�s�Z=� �U � 6Ǟ`����(��z@Ns�Ix���q��r����  
=�_m+]n���R*REUUU
�i��l��y��`t�ڀr���`�@2 �`���;��꒩��:3��   *��S` >��]:
�΂U���`A�@e����@��(9 ��=��
  �AJR�x���BJ�"()
+M*�|'���j{9 �Y�B� �r �d�ǘ�t	g���{�=�  J�ꔢ� ���g}�<{�R��y �b�F@j[��V ��`;�<��"��>}    �     ��� ���M� (�� ���)*��A�    ��T�)�       l� J�F       I��U( � �4  B�=Sz�M@ѨѤ�=G��=FF�)��?��߻��������@�iP��Q Q��N��zS���o�zsO>~�AW��L}��x�$AWDT������D�:���?��b��X?��U_��" ����?� PA|����~~~l'���2x�����633����2c8���Ɍv�0cL8�c<c`1���<dƘ1��`�Ox�1�:ld�d�`�Lc�1�d�N�q��`�q�:lg�	�d�`�q���L`�q�<q�q��Ld�ǉ��l�Ɍ8��Ɍ���4���ˌÏ�8Ì�Ɍt�����8���1��Ɍ��c8��8Í�1�L`��c��q�;g1�1��0tÌɌt�0�&0��2�&2�M�2c'l8�.0�.1�0�!�7�'e��\e�Lg�1�N�x�ˌ�Ɍ3��0��1�'1�q���La�N�q��q��:`�g;c���3�c>3���7l��L�8�1��8���1�c8�1�c1�����:c�1�g�0`�1�c�q�c�n��q��<q��q���1��8�1���3�����c3��2c�1��q�g�c1�n��:c�1�c1��1�g�q�`�1�g�8�1��0c��x�ǌ��0c�3��<1�c�g�c�1�g�1�c�cƙ�q�cc�q���q�1��Ln1������3��M�c1��3��8Ǎ��g�q�g�q��xc8�l�8�3���38��1�`�1�c�q�c��3���8ɍ���c�q�g���0cό�8�3��x�1�g�q��1�1�g�1��1�zx�8�1=�c�q�g�:c�q�g�Ƙ�q��q�c�q���8�lc8��c�1��g�q�c�q�c��3��1�c8�3��8�N<1�g�1�c�q�cǏc�q��1�g�g�1�g�g�&�g�1��q���n��z`�1�c�q�c�c8�1���3�c��c���3�c8�3���3����1�c1�g�8����ό��1�ǌcg�q�g�q�ǎ0c�3��8�2c'n<`�`�q�d�q�g����Ì�3�L�c � 8�8¸�8�8���8¸�t�ʸ¸�=�.2�22�21�*c
�q�q�1�q�q�q�1�d\a`\deLaaS�q�q�1�;d`G �dddL``WGW��2���c(� �ȸ�8�8ʝ3����c
��8�8ʸ�8�8�0�<`ed\da`eLd\a8Ș�8¸�>2�2.2.0�2�2�0���d\ae\eae`2&0�00�0�� �(�(� �'l!����*c
c(� ʘ�8�c L���+�#���#��������Ș���8ʝ�0.0.2�0�228�<`���D��T��E�T�A��G��T���A�A�d	�1�q�1�1�q�q�q�1�q�q�≌�����*c
�*�
��0.0�L�c �8�8�22��L+�����#���#�������q�q�q�1�|eaLdeL`a\cReL`adadee`�
c �*� � �ʘ�8�8�8��c
�(��8�8�8�8�2�2&2� �P1�q�q�1�q�1��WS� 1�a\e`�GSWG@� 1�f`G �1�dC@�T�#��c*��2�0.2��L����v�&2���c0���� 0 v¦�c"��&2)���xȘ�'�q�\azd�Aa1�c�0c3�ݳ��=2c.2c=1��3�&3�q�`�q�<`�f�g1�g�	��`�`�g`�g1�񱃌��0�1ۏ:`�\`��1��N�q�`�e��`1��Lblg1�1�d�ǉ�8���3�&0c8ÌɌ��8�1�g1�g1�1��0c�8�F<`�q��1��1�1�8��q�1���a�^�pa�d�\d�a�Ld�g1�lfd�e��1�`�1�1���Ɍ������3���������t�Ɍ��&0cq�`�g<`�Lg�`�`�1��e�`�&�\`�\`�Llfd�`�g<q��q�1�`�aƘ�a�a�{s��$�����y�� ���s�� ͑fcʘ���\�F�fYەrRt�vd��-ɗ��޽w��`�+͙����m6��sM݀�X�+F
�X�Y�V���),��m�U�z��Ud�mlZ�V�T����H�C�n����6��=���h8���*��K�XV��s*t͓�WG&R�(�kt2i�[2겎Vl�K�ݭ���YAn[���n�h!r"�Á_�����h-�na��a���W�ҙ���m�n��IgMMM���TY�l�ń3U��ӧ��V(���L;kEeD`I&�
f�f���� ^�fG)8�ъ�T��"�s4�y9r��d��A]�[�Z֚Z�
+6r�h�d"oi��8��6ڼ�m�̢@&����c�P6M��əGULr�w�{v�ɀA�h�U(��J��uj�]��l�;�ҷYb������n�7^�p���Z������Z2�Xw�61ZT�R˻Tw@�t�k�"��/N�ӥ��^�r�zn�աC2¼��Q�d�Z��"[��WH]M�,	�m�.�F��̽����4�XEj�����v�0�#q=O�vtU!�t�ƌ�֥�5^ӣ{� ʖM^]"��R�2R�)w��u�(�;w,=>@����t&�a��ݹ�j�P� �ЎҡZlB�+���l\�Df�B�m����'P�b�H�j͑�ةC
����{x3%3��:/#^�fTw���W�As-[�͎��q�A����1�mX�ib��KV,(2��>#1�-S�n�ce�a���)ݙ��U�=p�W�Ѭ`���t�D�f�̵�f�{vP�Ue�Z�yQsn�@��)���6T�l��GX6qk5&b�63w̠vJ� ��P�%{g��Q�v���-�������,ʁ	Ai�oN��M� ��5�*yLw)㩔�`X�����S5���iYd���N��Z�҆=��V�ox��A���v�盼����^2e�ՠ]Y�t��t�Ndn�ӷ�s��.��ݭ���
fF$[��m��ҫ'c6ܺ
ڣ���ج:�m�۴�+b!�u�A�1W1��*�`݄]Wb�Ût��S ˶"mD���Sw�5������y/�ț�p���F�ˇЙz�樘4H�yz���7r��P�1-��wv�VE�kX-S���,ل������D��J��w@�Q�PY�啹5뽽9{Y��*xS̥�)i��n�7�s}���'4�VN��°�̦u<��-ֵx^U݈���dC0��
�b��7��z/Z�ц��K�܎���:7^S{���ڗXl�q%r�&�֣��X�xS�����4�˹4�e�%�du\�֌�4�[�t������f�nj��En]*ik�n��V�V�n���kt�v�Kw���=��`U�7[��L�����DI�FUʲQA����v�{�����Wu	;��)f%5/-=X4Ći���
�0]�n��)L��x�f�B�CW����$�����+}�en۸
�c���K4�rX����݆���/6��wkrb�],ݫ��*��l�G�`;zr�6�'O�ê� ���2��]�;r�L�2��lS�
�77S�����J֭��yn0гV�3P3Cy#���"Y�����]n��)ovm�&��+T���,�M[b��/q�V��t�+h�ͺ�xc̪F�@d%��[��Z$�����F��h�;w��w.�؋4����v�-��x6dh�kU��e�[� �9���)ڶ��8�k�/5n�֨8�YiF*Fma�1�V�fy�����w,��{e�n��&�]�f�;�j��K �ѧw�Y�%�F�f7p\�VE�&�uj�і�k���L>�[uy����f�z�f��m�1��-��
�P�Q3 ��H�z�d�i�L6Q��`b�.V�]-����m��kwsw�$�x���R@]椀P7x�i4�ڰ����k5ݝ.�F�^�)�جLl���Q�D=ֆ�;ו��P5���h�YBֵ�i$N�(�b�[����x�u�;�-���/t�Q���dU�����U���,���l���ܕ5�E5tG)�r�m4�ر�Wt�M"��;7S�v�
�70��
�e[�2�S�ym^�CmG��[��wS���a�/i�����l�iC�,����-��r�^�X
y[��w�v$){�0xL��h렪��2�n͊�wgPw,�
�;�-����ȶ�0Nha�0�s"����d�eX�kHƪB6�ǵ,ȱ^oo�^RV-�����7,=m<�Yzá�k4=Aa�"Zn��3�DIY�V��R�5y/R�8FJPQz�K���L� T �]K�Y7wj]�R��&��r{�q<�dz�rٻ�.:������hժ��)Ȳ���%�FM��۩�cJ�苺�j�LQ��&iWf�iU�5����lU��:j�� q�l/hT�6U�{g}��w��v�0��ժ�B�9�Sw�VQ+n�4[ M%˻D��+*`ZFh�Bk���Nh5zE��wxn��m��bT4��f�#�\�Z�<#7)ކ�]�X�"�D�U-�ὂ	��r� R��VU��R��RiG`�z�h7Y�]އ[x�/]٠�:�g)3�m*�
�/^=�v3_���e+�&��b�Crȷ�S��״]؍�ml�[����B�1<���X�5���$x=4m����f63/C�Sy�1mX�S�n�m�sn629��AGgn�N�p�`�����Q�J�
]NTB"�U��O<7�7ݽ�T�׷[�5K.ݺe!t���hjղ���+agqQ�l�Ni��(�m����F��^�m
������A;VNV^@��CY�4�$4�Jՙ��+
��J�
J���z���9C5�d�,�~ ����ݚ�yNk ��ʳ���Փ��Fx��[k��[�S�b
��c�Slc�5�f'��a���aY8W���7��0��G%�Yhfѱ%+��iY�1V�+r�PU�n��T�K/VIz��JG�$�Klf M,-,���y�-��Fܣ���"w&,�w[�ON��/+���+��i0)��0�[�.�J�!g��lR�u3�D�g$�H���w�X� [mR�fKi����ۙ�4Ҋځn�la]���.�f���!Gv�n�u�SF�ыU��%+!&(FCCs]�m�q��l�S�0�։hͫ�Z��-�ޛ�9�W�QЊF��iG(�ֲ�S���n�C8�\��Ufh��P�sq�Zn�{y{Z��-b�Q=�w*3`�u�tdy
�,��I;��ފ�A�%73#̤j�������wy�����M��ȴ�1oA`�Ulfe�C�2��Mc̹Wsi�^7����*�f\��7B���J歑�˃D����#�3�B���`Y�x�^��w%�%$���u��M5r�W	;��Ы5^^aY�N�6�,*KH^]�����ڃK��MfjK+op&Pwq��e$�o�xn�"�&�6pt���k:r��[���	�WmH�ǃm]d��^]+�V]j'V�^��#l�X��Q�4��@��^��*e�X�'�����t5�x�7�XͷM����x.����gu*#RZ+v���͢u]j���NϜb�Ig-�j,���L{�A�⣪���Cw�T��t������� �7���$�ӭ�|2^���N-ӓ�/n~���k,�:�����L\.���9�c� or-��Y��a&�eֶ�UDkO ����)�P�l�p�kP^ZĚ�h��̾�(҉������IJ.��+r�g6�U�[37]'�}����X�(K/N�����ܙZ��i�F��oTn@�'7	^�b��ьtK�hI0mm�k�@�,�BI���dӂ�3�ٴr��8�oI��qi�͙1�6�Z�Զ���7�Z"]�t��E��#Ԋ�v�gJis-��h0��F�q����4Ә�6.�M�.�x��-Z�i"Z�Pۥ�ҡ��ݘ��B�s4�"mc�ɗQ暷u/��-��7kb8mn^��q^����K�.�X���n�*
]\�P�gr�ث����ґ��7zh(��U�3c.1AKÖܢ��`5��͑���"�o#:��+�2�WwQ<�*)j`�T4�(剗�h���4�e�Y���.Е��P��9Iհ��`[٦��I]�%�Z��� -�@B
�x#ۤC��
k72Z�e��O�Q�����u*̧&j��J�ԡJe��f�0��r�C�[�<W1h՘�gjk�XYafT��^�"\����!�2�а�n�R����`�4or򠲳(*Fl��Q�w�n�5������)4�ڃr��ka"e��óL�d���U�)k�<`A�o72 �f�X-����z�e�:/�Ґ���6!O]7f�h�$�*P�֮lX���,5*^�������0:�����nM�U�VF�Yc+3!�.��R�Z����@�n�lѽVe��gn�Z�g�X�	Z�&b.]a܂�la��'i	j%��Cw5=R��e���zo�
-�@'d����oXΦ��
��"T����y���ܱ2
��������K��olBTjf�`@2��6���i����6L�(�񺛌i�Qӓj)in�nf�́ �^��pD�nK�l�ӭ���V��-y��ؘ(mѩ���`�)b��f��ƙW��ȋY�I7o3QԢ�Vz$�a�u���Ǭ����E6������Um*r�Gj�*D�2��mRaT�rޛ��*�X�n��c9q��O#M�Yl�
9w���
�^����f;	��R�u�jMnܬ���]l�5��k�U5��<�˫����ݦ��XjY�n]�J�o'��ɤ�:��Բ� ZL��a��jAr�=�4�<�;�ݗ���l)�I6+Y�lRX�0Vm(�t���t�
�9�[X*��9�[���R�Mx��|p
UM���1X��Z�8�F͘-�h��˻9Zo2�]�4�nƲ<њ�^���a��9B�Y�e�e�`1+d6���U�Fj=�.��k���{�1ڋ"�[4�"Vǘ�+yJ@�nȬrH���F`GN�uҔ5�Ӹ����|���Ct&l��e����E���ه2��x���j�C`��cMz@(��MeM�Y��	R���+[x�� 6=�n�=ݺ��bY���Q"1�H�:}�j���̗d"�e��o7t�׺)P�]Z��O,�\gĊ�~���������*�/���e�d�+M��i8���K�Wk�T��mu��Z:��*A��5gQ��d����'��&i{3>f�0�V���I7��&r��捸�t��{��Q}�`�\�.�����вB9@v*�tLvyxr0�j�������+�8N}Y��-���ژ����'����{
�a,1��l�C8D���O>��w�>�uz���Y�M��Z�a:E�	��'�Ҿ3I(�9��n���~�LK��.�2������^��]Yޜ4@wK�P1^�Q�t���g}�hl�����]6��1ʭ)Eׇc��홇������Q�Z�h5�N�CzE��3y���=@�o ��:Yf��8ȧ����$����Z��v����<��gg0�#�hDl�ԟT�%�@&�尽Fj���I���]~�
R�$�� ��V�P���{�P�=����=���q��S+NYj~����������儞%�^���P�eTOz�l�Z�'�6�U�xM Mвg@
��wKߞ��l�0���R�y��t�2�߉fiH�=b��'��I;�1�gK�b�2��	JY@�e"��H�)S��$<�!�B�tW��p��t$��;
�}�Y���[�ء(�V'�=��w_*��3���c��u�+Й'N�������C��f��~]
�5�m�U�f���e"�zL.�3d�<J�p�������NE:�]�A��*�.Y�R�Q�i r��I)�S�A#5*I'I���a������0��5J��֯�ޔ*�<��h�Ǻ�,Xޑ���x�g~+I'0��4��o��\�����������	�{J�K�1�$�s�U�;vш�'	��"��YZpS������2v���>�Z�t��IAw��:g�F̯����J��8��*v��r�D?a�2�?'���>_�b9���7�d�����+
�X��8�n�O��5�1����G�����Z�E,y3�y']����²>��y���m)Q�/)�`�H++�'˒�Gq��ق��+L����A�,ѿZ:����K�B�*����i�-K?2��J�Y�8�ɰ��КM��~����C�7>�����{6�v� e��|��7���;�`��Q���!I��P�NI&�$��uzC�~d�xQ7���o�����at8���~�w<�PXG�/�8�)���7gI�.�
�$Q��"��E��7;[�_�Oƣy,��ő��Je9R��L�c�l�&�3�I�zK캹w����
�q,oE.�Y\u��KM���%�+8�d|p�����Ax]��h�3v]��a�����Iunb,�)��Qp|(�����6�Ϸ�[��ms_<�yQ_�i��O��]9I_wG�w���
�.�k=:�ʄ�P��c޻��'>:�Ҿ8NPt���&��V*}g�W�n����jYH�ws䒐]����#sI�t� W�T)��L2Ƞ>��}���_yz �X��::�#�e��ģ�$��T���;�L�>�U6�xI��JRKڽY=�<A�)}�i��|��$�J+�=��>�e��,��Lפ��н8M������8����JTJ|���6�W��v��n�VrN�S󳜠Y�oC��q(V)Cd��;q��\��mޙCp�L�Z�'?�~G�+���(�u��]*�O):��g�싌FG�sNi��$��0��Y�9f���I���o��K�">v�0���-��Yh�E����'�,�.�e|����o9}I|O�Pf�\��6M�7�4�k�JAK;�S;�k�8��Fg����_9>�0���8?B3T
Q�PZV�)AhiD) h��P�(EhA)JZAV�F�B�E�J)U)��)T"JE��) 
@�D�EJ �)�P�E�F�Z@Z(A�(@�@�)D�T(JE�h(A)�����
U�F�h�
E�hPi)@) i@V�@�D�((Q
��U�DJF�F�T��U(F�@�;���@~.�a<~�}��@����I��NbX3;XhPD�`Ӊ��� �;N��K�����{����u�h��|�bs���ҁ�}s��&`�i�-:�> 0�;��+V� 3�<����)�lǂw^�P'U�y�:Τ�4�S�!P뗙�ܲCԋ��ZLH�]���	޴�̌�0����!6@lզ� ��54� .Ms�Y�����
���� k��@>d��̒�����I=v�cԞ�7�䓾]{`q8��T�l�'Y��;�|�i��S܆]ARc7�\�dY��`�Oh}�	�q:��c;�}�$<B��$1�Y��Bu�i4��CԚORh���v�|��V���'ݧ��!權u�E�'�'o{�>�w
L�O��0��@�˴��h��vkr����;�:�^����RWy̗$7�)ܙ{	�} �=�ߴ��ٟs�IĞ�d7�2]<�d�N%%�bŻ�a�j^�_�Y��`�����	̘��%��k+w%�'� ����Ӏt�=�����������ϨJ���� bF�g!Ȋ�P��w�L �y�с�� �p�"��A#�Ń�� I���Ú�$���䁛��Y@�˸���w� ���QS���?>�E S��}��?��{���3f��v�������!�R���~߰?ɪ���w8�Z+�5sO<���;�,���屰ձ�Ң܍�S������2�Kf�s�ݝ�n]	+{h^���X囃���2(>m�:ߌ�ֶ�K��VxY;��]Z!�(m�yجѕ�mWÂ� �(��]_�\��NWndU��̎'ʊy��ya�r��\2��s6���a��bYwSoj�^W�na�j���(��������%GR�WO.
а��fSw{�p���Х��ۦ���Q�0a�p��od����zΪW�k6�.
�1�Ę 	L��C<S2	2�Z�Y5ٹ���8��2��詾k�{V��x�ÆMЭ��s����gw]^�����ݷoHҔ�ʺ銊j.�L�BX�)�Q���� *B8q�K3�r��2��ƃg3����x�|^�� ��Cݜ
X)�������^Q��1"��Q�0�	�]�!����YZ��*�2�2�ve�'vӝ�R�P���Xۻ��|6^�:�C�3j�(�� ͬ��wG[\5���S6�қ't��D�p��r�z�er�JK͜���a�VK!E�6�M�D8���<������>����>���n�뮾::�u�\q�����]~:��]u�^�u�]|u�^:뮺��]g]u�]u��G]u�]u�_]g]u��Y�]}u�u�]u�_���������~:뮺���Y�]u�]u���]u�]u��u�]u��]u���]u�_u�^�fu�]u��]u��:뮽:뮺뎏�{�;ތoWU�qW!��J�٩*�r�equ����{}��{�չ�*�vpG���e����2�*��u���/�6�Ϣ����G��op]��1��Lo]wwij�/�}0�S���Һҍ&j�S�U =����T6�������k��J����Y��-�-U࣡Q[���X�Ʃ��8��K�>��e��q�շ<Ǩu���nS�2���r����n>�HE&���z�҃��Ȫ�Ӽ'pc�����g`j����
�MX[p��L�|3yhƒ��Y|gD5�4K�-������k0�S�_.k��u�V5R�=v��{r� ���r�i8un�����7���˼[F�y�zvp�Zi
��.#������~��n�ຈ�:��l��az:)��23=��(�̭��݇.Y�Ɏp�L9���~���c��uw`�5��s��#�:���s��[�h��W�p��\=G^%W%�j�z�c��%�x������"a�c�,��_y��`�5[[������60"7������������}}u�]|u��]|tu���]u�||||u�]}u�u�]u��]u��]u׷]u�_u׎�뮺����]u�]u�]u�]u�]u��]u�]u�����������^�u�]|u�^:뮺��G]u�]u�]tu�]u�\u�^�u�]u��]u�tu�]u��]u�\g]u�^��{���?��^'�%��*fT��A[\*Z®r&��߉�\�]�V�gd�ÈܡY�����
����Bd!�a��a��Z	C1 !U��i��e��s���/��L��m k�� ��R����Ig8F�u� Ȣ�i	w��ǜ�4`���Bxi8}UDUW�Zpݙ�-�1���$d�L��P�uU��;空M5X\��^; �Q��R���j�B��\Z�ӹY:.hC�-i�%@��;����k�K
+t;+M�ꉠ�K�#�����շC���Dm��X{�������!��٦���C��eXu��+MD��]�|-8�(M�QYEYPH��̘}{�V"����� 	2Q�uݰKZ�0���ھ����J����8�.��wY6��Ǡʍ�'Y���A"�T�����^^=���Q�E�V
wU���Qo_3v��_v0�J�b����xo��T��]�ʛ��p����,ր����Yf!�R�q*��f)�:�bF�nSN� ��h�&6J\KF\��@��X���5U�H�v�:s�i�'7�.�n{7%�uU\t�� ���o�OE�7��р!��]�;���W��gN!�������"�C�;����/kzؚ��Pj�Oojr�U5�lOV�X �5V��'o4ר��Fs���lV{U��}^�#�Uh#Qŷ%�xstܾ����R���y
��uņ��߼K� a��g���v�:$�)S�YO���J�Y��8���X�Xʼ����5�����63�64�뮺���]ztu�G��믎>>>>:뮾�:뮺뮿u㮺뮾:뮽�뮽:뮺뎺κ뮺믮�κ뮺믮�κ뮺뮾���������_u�^�u�^�u�]u�]u㮺뮺�tu�]u�]~:��]g]u�]~:�C���뮾:뮽�:뮺�㮻���
���[���N�$��mx�iC�t���z����ۻ�������'��^�_gg�줸eӭ�=:�Vh�x�3uv�+Y�����c���oE��7�ض��=aՔU����y���g^�T����W/�{��P�.��F
�[���W���Ll���U����5U%�-J���uΆټ�ˡǗ%�e1����+�euj�F�2�ͷ�l��qg��;	�U]=������o�+�AƦ��Q>�|n(^Ә�F�R���bF�
�e�+�:�'�OF�X���
#�=���ȩ�[ٕ"2붕�R/*��-t [�)��Z5XW�o�;Uu�i���Z�o��J�дe�5Y2*�QW�/��kE�Ol֊�����O��k��l�f�����C7ݳ��<)N��i@z�o:^���΅�p��<-c��ɓ�j���}Qѥ�b՚b����9�lJͩA�6�����洽�x���w���P\�M��
P�.d�Ԡ�
Q����E����*�xd#�N�*��`�n񚣸���z\�g�ڱaE�L�^�,�s�ṓGs��t�["ŧ�ϒ!�mœ��/��A U�����y\Y�m�9Kk:n��f���g�k��$���N�RW)�C��V��^������2id�������������]u�_�����뮺�뮾>8���뮺��:κ뮺뮺κ뮺뎺�Ӯ�뮾:뮽�뮽:뮺뎺�N�뮺㮺��]u�___�?��~:뮸뮽:뮺�㮺�ۮ��Ӯ�뮸�뮺뮺�뮼u�]u��_^��뮺뎺�ӣ���kkkSkkk;[LLt�D���c`�I��6�rU���v��Ա�_'���n����Rb!����]ë���芹��7�֟(ǷG�d�yy*Z�9,�ڻ(�{�ڃC�rܭ���;~�g�I�KH3%,��ؔ�/m��:�)]Hs�k���xE������ڠ@�S}w��,�3W�`	�Q�丞��s���U�=CMFj̤ۣ&�gf�+s|�e��R��jg�H]B�&��]V���+�.7/���p��gv�ub��.��O3�sls�I�e�o(`�����h��X�yw)7�k ��8 �\�d�^�՚�[����=׎PMx^<��\���I�&=����b�8���M(���t-�ۢV�s�TZ��k7w��3]VWZܕ�MVu�ي�0�޼U�k��Z�����[�x����;@ʞ��ŗI5kn
Cމq�&G,P�`N�9��œ��u��wn�Sy�n,^���v�{R�YJ[s�`OF��[y�a�i�x2V����ݳ�P����4����vmj��C2z+t�q��*<e"��H\�3����3�1�p�#,w���0B�7檢(�鷗է�{T��M]��cٯJ��+�wm;8'��,��(����J�������r�4OL]��������{���OO����:뮺���㮳���믏��oOn�뮸뮼u�]u�_���믎�믯��u�]u�\u�^�u�]{u�]u��]u׷]u�_u�]{u�]}}}}~����]u�_]g]u�]u�]u��]u׷]u�_u׎�뮺����]u��]u�]~0뮼u�]u�믯N�u㮺뭭m����i�4<D;�ӛ�_fVS�r��NDK����e�ق�Jc5��w��+�8�c��З��\�j�5�\�ͱ+F���X��P�UR��Y�̥~��oo��,��}3�f��=z|'D�;�r�w,�{y�c9mv�r�Tm�}�` 5��� R/c$�uW+:3B�u���f��0+�
�˭r�n�
��N���X�Ѽúh�(�p^��-\�RS��-U�i��) u��ev�{������gc'�:���Tg&b��R�� ,���C�g-�s9cn���6-���]�n�j?xa��2�N�v
v��%���OE[�*�S�B�n�H	�v���f���uZ.���[���5ף���$(.
:yT3s��l�.�oO+����BJu\p������{LM�u�8�KV������M�4n`�)B�m]�M�0ݻ��8Nڤ�kv!̪R����U��}&,�u�X�:o�S{Y�b�n2qҾ7��)�Z��ժ:[��:��beo6�J��k�5�ޛ���}�K�n�(,�^���g7���Þ	em�T��;�+r�z6
��l�
�F���K��ɸ�WN�bɡ���������6666�N�뮺��u�u�_||||{u��]u��]u��]u�\u�u�]u�]}tu�]u�]~:�ǧ]u�]q�]u��]u�]q�]zu�]u��]u��������㮺뮾�:뮺뮺��:뮺�:�N�뮽�뮺��뮺�ۮ�믎����Ӯ�믮�:�u�]u��מ�[�4�:�;;�+���8�볹nʻ���i1�_hݕ�Nս#�{9
��;�1���u��uQ�U�R�;��3��B�W�О�wglG9�)�^Ӻ�O=z�FѴho�!w����cN�^ŷ�r�V��">�܁[���W~����˾L��*5�h���[���Q��U/�]u�+%s�,ѮMμ����}�+n�qp�ȩ�glZX猛Cyp�X���T��d�+���l����2�s���w���:Źۄɱ� ���h�u���`Ϳ`v�?XtP�M�ݫ��+���*+�5]�cSq_Q��`ʼ�]`�{�EƳyzrv�nj��UL���t%x�������
�Z�UTٽ�%<Ѭ�oC�6�N�ہ��Sg�=���i,��#r���L�����tmGHSW廼��&�Ð����޳��Ur(s8��.�ڵ4L�;u�nkں0�!�un�3�'],��V�U��f���o&ݳ@�[H�ٓr���\���Z� ��X��h��ec��Ӻ����aδ���*�0���:jnL�-�!z5���A9`1mZT�T5�M����ݾ��(̋g8gaz�nq*���mJ�VGW'v �>!j�9:Ճ��<j#���(-�u���KIc�̰��;W2�W�x�*�g���
���$۵�7�0�Ev��6��f��G�ANU�-��M��Ms��t��T��A�Cx:��tʃqX5�!����+M+ܜޜ��6�aN��I�m�v�ڇ���^��d�k���Z`�W�iT�&	��-M�覚9��í".r�U���Է����:�4䘮��81y�5��6�]gu�ݷ����R�ȳ܆o<�&]�Y���O��yS���,[csu�	Yɫ���d�5ۛ�M�uuu��ճF�"2Щ�ᷓ�T�T7�e�e[{�\�]ټb푫ܼ�BOE���9�8E�������C�X�5y��h���"̰��i�a܋p�X!����ʭ��\�s�sv�eP�hZW+�P�@F3�Ev,0(��{�g�;�� �~s��m��.��&�nO5��f��>Ղ�dGU�gΝn'E�n���ݡ��QF�`�� ]��i�ft�59ʌឲ�goc��))s��n�O3Y�ykn.0R��f�w<\F�i�
ʺ鯦��+��ŏ��SN��tJ��m��
��[3�I~������5�Łyۑ�:�<�{O�]���Z�vu���2��w�f��<������ڴ����j����L�,=����<=��dB���=�һ��pegID����Yv��Ґ�+D�v�:X���X��}���9�j�u��&Z�}��s���Z��vf+v��e�}��(�յd�;qj��v�q��ܶo���`�5n-뙯rA�
��s���ì�Q��le��+)l���4s�{�̭�me�}�e6�M�!C���L�fʴ�{A���04M�^���i��\�`�������7�[k���1�X���6!�@a�m�s/d7��g�������R)4�z��nۮv��n����@�vH1�^������j�z]�;a�I��Æ��p5�7J�\�gK7�0�2rUΪ�쥸�qwi���;4�܅䷗��jg��N����p���X��X�l�xC�t8�!wa�c�9�/V��k���7}���p�]ܲ��[���G2�t�KiVh���a�ͪ#��t't3
W6�8��=r�.kB�{��K���<AV3��ق��m�YW7w޸�_f�=��y��~�u���V/S�Aͣ�3(+.��$U܎ˬ�C/k�R��Sy� S�2���RǄ�~{�F_�k0�}�*���ȱ��޵b�g ^��;��J�Ӹ�q�Z8
̬�ŵ`k���E^��8`��'v�(���t��h�%Y��:5u��#v�Qp�8M��S��]bMG��J��A���;;/9	jαL�sV��Cp�Yn��z
Ⲟ�)�InM �n�����Zy���7@�-��>9��Eͭ�wod=%�[L�`,_U�xbm��q�F��Y}Çm4��fA,�����N�g 7c��s��د�O^u��we^��'TU!�Z<�PH9�-$cWZ�mX�˹�u�%��+P��y�v�Rf�(@�U6��{qs�a'&N#�۱�2Ծ���U-۽ۗ��� kNɬm^#�hxeqPھ�-��sqn��ZA����]e����a� �鶆ĝ�x�ehұ�]`�Yռ�:a����o+���Gg���J�l!Go-�o�B��,�<<���m*`���ϳ�suw���],�J�1���"CfiY
���!�ӬY*F�3��  `�33~�K����������~���p�/����~�	eHP��^%��"Rƥ�����bf\��7yמ��Qft�em�f�*P������g�hb��;�Q����z�3A6�P-��[�|����J @%7[ˈ�n\��Gj�7;CMގ�c�ZY�Cm�����
o/���޽6m����W�vZ�Z�cIn=1�(�����+�,o��`io�=Z:XK����=�}]|��9<F{5���.��ˋ-@"e�n��
��x����]2�4��ѫ��4|�k�w���P��d`o����3����=�l�;$��N<Yi�M]�����!�&)��y-�4��v���so��o�C�6X�3JV3�?^����F*$j���fyu��כh��䵄m m1X��ʫ��YFh;��΁>��_�]�"���
.�l����+��6�I��a�R�)�p,"�Ļe��bՉ4e�.�jj�QY���0��*�+P�G[E�r�]�m�dl�]xI���(�8Lm�ڹ�r]��T�F�tel�0�j�i�!*qT�e��2�-�Ĺ#3p\�%v��2��k���C@4J�μ�X��2�+YQ�
ҹ������]�i�C�/j�"B22�ؙ�Q�R�
�L�3������F���jE��͙�E���wQ��3f� �l$Jk�;@5Wj���VWT��,�!Gqk�Z��Fl۬pM�[�@�"�QY(�)s+�1���f7a-\�]�)r�h�
3L-3�j1�u�n0�q�`C����-�)pB��F���R�l���]�Z킍t�ڎH8p�BV�]fYsVS.��.ф��u&��ʵ�:�)����u\LPS�SF 	�F6T��a�F1��Uv�m�\Q����s�d�!�ƭY��f�-6�!n�d�bhVԹ���b��؂m���K	��֮3Vaf�ep���\Mn����k��Ҥ��%آ�6�6GhY�\��YB^CD9	��Ά�ƹ�-��͖X�GP�"�s�+B����x���SJդ��,�*����hf6�ͭ2(ړ�YWb�̩qE��CL�[��i�K�um%�s2�XX0�ƺm����j�!)%q�֗L�mv�5��V��.��d-�����u�g1���3�[@�+S�4�H엗i��k(B���>6���Wĉ.r0uGb�Hb՚"�j���a�L2�-b��Xb��G������Y�qv����������G����Ѷ����$n�S�l��ҷ��F��u����k��n��
��]�0���m�d��i���e�RT�g,��DV���&h�kF젇j��ils�[�Aщ[4�Ɣ
�.��tɱ���v����%�U�vh�,46�f�lŶ�5�������Fnա�#��2b�2,Ж՜Q��.�X-����Wb��� ۢ���&6Rį# Ѻ�^
�k��b�&5�j�֮l��k�7��:�̮rf-	��,b�Wj6b�8�Mu@2�j�m�DSA���UU��p���K,-A�5�t�YYnB�K�gHJ��V[e�;G0f�K��1Ř�r��2j-\�����F�l�F���  ���3�(�����c3a���c+��l+�����$iZ^t�q�,��������I���&KvtƎ&6�Y�F0����T���7S&�&!<�Υ+#f�i.�v���AҰ�b��K��k��񎻪K%)H/6͝eae)V
�cS&�$-�.�mGd��D&�2��DU�l�B�f���f��E �8Q@��ճEԅ�um.�@V״��(��B�$�{$[Yt͂ܡjY�bv�*�P�T�e�3(�J�f���b����A�2�oP�5��4����������
�<6]f)`�[�m�×u�m1��ި��e�jWm��:��3I����$��cKfe"�mk���J-��Z62��-�6�=k��JRk0J�b�hf �J��j����sw+4�*	��6��{ÛpU"T��L9kZ��ˋ�Vۅ��[�E��6%.�-@�mI��-u%%�[�[1m�j㘍n��GP�$J��電\�����I��a�#'��V틨^3jM�f	�JX�*,tt%YWK+e����6mp`���,�(#�0�/\iuԑ�A��p�L�����V��uXSV�8����s���z�͵�#�D#����riYQP1,ZMJƇbʹ�e�I�E ]�K���ǆ���2G�1��a`c�eԻFƒ��[���f��+�e��5!���GL���M�7lB�`�r����)ka�u�H��&f�F��h�`P�`��e�#���(Iv����,!@j��kZĺ��0fKSM�hd�3LJ�J)eX-���2F�n�@�4^�k�QU%����j(��3V�C."́i�ٕ��m%�gCx����Y+D������W��0�8\X�]����f-JE���1��eIGd�i��؎s,J�.뱗h�[�����@�4���e��B�֑�XP8���5��WeLX���iCd,ƮT-�
��(�]��a��:iP���<���TU3`�2��m]��m�ց[�jF0p�%��*Ա֛J)��:�j���p ��Xĺ�e����W"�!5�,���|rI�1,\jԛ��]����c)n���Xn��Ը�i�X"�m��2P���fU�����i�:�n&�{E����X��9(����ۚh=m)�3j �,�e���uڜm�fYT�2´m�t&�+6�J������T�:���H�����M
$�S-�mfWM]m!��-�b�)�{GZ��X�ʉk�8��b�,%a�]SFSh\k4l��s���zau1��3�.4���6(�Q0�J�[�TkX7s`�[�Ir��m���#�)����p”�,�
�]s��K�%��٥��F�l��\M��W��0��+1m��q����f/,�Q�7^B�J��z�i��*��A���Z	Yit�]�E���:ݬ�@!F䎁
�B�A��*Mm±����Q�`h��K4�l�	0�1��؎��[cvu�jlq���-�2�\��M{C3M�1ݦ�ñ�H���][6�K� ��JT��Q��|��uh8��%�X� 4%�sV�j�ژ��5�:�Wki̦��iT�R� �V�^�vX0ufױY��1�Y`#5�!��e�f V���b��HYs.��:T�(��YJYfґ�K*q-l�@��d1��@D���f��%��F��͓D2�b��o���39Kv��YH#D�R���\�@tH� �-��
YcKS��`�۸����
�&<!q�%���˔v�Óh�$�W%�m���&-�ZS�*��x�Gu�%ؔ�шv�X�����h���A1L�˥e#6������ėuK-��v���Zh��L�b�u��2��gQ�J̲��.�p5�Eq��
�ڶ�X&�6�t�Ű��e5�ɲ5���3u���d�d�N�kWj)I��c.�P�����^N�f�2��`�#�fX A!rl��Cb\�*�h/]�Ń�nv(pqtFۚ΂*ש-Ժ�������bWXK�eͮ[H.[�,Hc�D�C�`����v�W��kk���mڔ�3��;V��=C2�g��R-���-tlI���bX����ms��� �b�e��^!��S���9�063�:�͒Y���-"��P�N�թh9��tе�X�-�ݜa6�s�P1�Y�۫5aS��Q���b�'��!���0e��B�K\q*&�k�fa)"
�W\�.�B)W]4��APhu�u�:��@��P��k"e�M���v�.���"2�+o-X.W$j����׆]�#U�^asvԍ�qF�3�4"�m�2���x��tn�6�-�et��f(Ji��:�үR�]�	-�j������&J�e�sl.Һ��i�p1�ѷ7X:g,�sQ���孚��X]T��j��U%�Q��m��1; �"�7:�W��K��7�kjF1F,XRٶ�ے
vmT��Rb^���,�3$nb�[G��YkAk�F���*�S9��Օnpb�{3W5�0�r���&����UBl6�%ÉPpYf4���j�ȁc�e)�mv��p\�h�=6�l�`���d�e�6���T���0]�m��x6]cTk�ȷ:4�Թ1��[VnR���7d��6���%�رLQ{Q���)u���@m��'�.�f����fm����o^�����kK<T�|o�hO���7�+1��s�:�Z	�u��������M4T͉q�)�k`FP5ŃJ��X�6��:���a6����:�&��ʑ�-iG������yJ�`�1l�#.GB��c'��}[=X`70(��_���F�m�mA��C�5�is���bUJB�D&ŕ��o<��e��Zg&�@Ö��\XA�ф�<h�H�	.jAe�L0v��8V[��i��]1��fU��7 ��)���<M���[��%p�Ǝ�)�O]�A-p���JK]�i�������CеŹXM����%`Mf6In9�f�aR»9unRÖmk��[%R%��D�[q�1�̤��"�^G��xOS��^��
1�͕�sI�n!aS1�(Z'`�M�w��8����pz���m�Ek��7SB�����9�)-� �2�^YX�;cB�GS
u�)[�������x�=t���YMr���=��ζ�W|�ao�
4�c���}�r[=��R���\���6[k�-X77� �)r���mֽI>GOx��{]�`ҫ��4Ͱl�o^G���˅$Qv�h�I�>Fz�>@]l~�Q7�5ۗ:a:�=�|��PP�\�{Knȯ�>�f��X�z'�7��f��g�@l��N�����ڪ2���0QЃ�5V�4*���QX�H��%��S��V"�"�������Q�xu����=���}{{{{{u�κ�[�QDo��f��b�J���5J+J��L��㍵�fB�E���O&F3n?�׷������u��c����:A�9ejTS
�X ���@�WiB%*��z���BE!+SHb�V�5ư���U�[IUu@�Vb����h)$�[t��"*XTb��� `��!]4\JT�Oc1
2KK'M��ZbJ#{<���f�'g�驩����;=�σ���3�U�,����!m�-��[�3�Y��!YX
��cl/�2퐹d.S٫��[�mm����%@mU$��(1�+�[%����9�
-k3�q9IQI�����g����^����ߣ��_�V}m���-�Z��A���ZK[PP�B��#)ji�����	(!׶z�����dz��2�KKe,��J1�S��M���[�j{=�7,g'����jjjjj|Nϧ��?_�0�Up��,�uqn��+]Z)���%%�VLS�[c���Vx4ʖ�K���S!�Q�L��5,f�'�����������O��{�`�Y�`
)�lձTbVѢ�.D�U4�4˺+ێ;��	�+�lJ8"�*9��Њ)zL�)�(ζ�[�]�F��L��*i��1]R����,~Jn�i��T��|�n��YR�Dĵ���-Зl*>��:����#���+��4�cF���F�"+Y_�q/Ϯ ��b}h��c,�y��BN���5q���e�~���^�uh �X��`�n�[!.�=�p��'�3<u��Ԧ|�3�@͆��!�g�`Z�nVRń�Yn�Kq�	�+��m)4׵4��HT����`8[���k.�C�fܐ!fѱIB���&#��˕�c1+mk�.l��"��܋���M4��Ś���f&ݜ5���B�SX���n��i�XQ��l�����6S���#�X�[����k�`�*X jJ�LZ�iM��G+�&�� �S:�&Ԛ�lAqv��/6�Zl�و
ᛶ&��y(�0�#�k��K`ڶU����L���`�h\3$���u*�7�\7f[�i���i)4[��.54M0[���t��wQL,����1�{g�afҋ[��"9�0\[�X�"d��܍��*I�4�� `�03@XZ�f�R00:ι,���K�vƵ!ʤ��d��V˵"�ab�m�ѤJ�C�6�����
�I�tr�6)Z��3It�WJij�A�VQ��%�vv��ZF\���f��o8y��M-Ύ�E�H�[��CkS3Kl4C�L�x+�5��M���h�5�A.a�ikkJ��b����{9�%\�kV�J�����d�֘�!��l��cL�e�9�dB���q�ꃀ�F�뫰�i�]���D�̹�Ƙ�:aAQ4VYp�RĚ�ekxU,M�j�5���`]1�e4�nnq��H���7J趎�ÌK�bWK`�
�.݇H�m)f�4,�e7[M`�ٛmA�8s\)vif�j���J�Үrc	F�Kf�;�-�(��L0�	a���B:0Z�oo���H�̯e^�1
j[��1.��l �6`��aZ�+0�\� ��Hq]�0ŗsZE�#i^�����޶���ն��̍���v�maM4j���m-K�z�ﻻ�O{��v�OF-�KիK=*�hu�5�*-��(�-[0�dD�o^e[Z6XV�������!հo6�YZ,l���F���,
ڲ�HQz�Rĕ�,F��lKm��P:�!V�Ė��c�eIbt!,!H���l%��j֗�䲬���V�,%j<B#}��r�F}V�S6ecjQ�X�hJ���C΋��T<$H���Oxߌ����p.����ۼr�@2W�m�r*O��|i���	�G'����FKW���>8Lw[�}�>��/�HS�y��5�]y��O����zU�Ar�����ԕB���6� ����_[��>�=��6f������΀�a�}*ۑߜ>�5L}������Թ��'�T'�����ߟ��#�.�4U�RX��g��`���z��ѹJtG���ʙ�3�<}8��<��P�E�ǈ��� ��b/-�V�\���Ҥ��
z�L�(H�W����)0�B�]ߵ�1;wV����{�*y6��kRl�)��j;囦!�4��Hi��aWp5��,*Ѫ����V�W�K�]�&_\��x�����5�+.�����4�%��!���þ��u����]��ާ��7mi��}��1O�4ϋs��&�}\;�x�[����L����gb2��i����|�`
@�و	�{B����鍫�>6�\��"pdM�;�������n�@�&�'}�ճ�^�Ƚ�b����3�˴Cy�/�ek�O�ﳺ���+���J�)P���H��:�Y�QRٴn����=�QV�uG^3��N�xl݋^����U��l��u3kosr1�^_j�h4�@���ن��O�qj5]����w{�睫�>^�}��9�u5�Y��Cu�_�~����h�� %g0���58�wϻ,e	[��X��0d 
̺ꊨ�f�W-D��u��v��a�Z�B�-
�j���ϝ+�^ 6�!��fN����7��вɦ_���QYw��e�g�޽R�y�p�	4����w�J���F<5��ok�m����%��k[[�H�������/�t�R�Ed��|�[wv|=hm��Q�����wg~�ϳ׿����l�*jGk�p��]llt�Ԙ���*�,�k���H����f5T��N��]{²�Dz|�{��ڡqB�gi � i$��_y������Q��+����׺�����c��ch���u��4zi��j(&"LJ'[ߝM#П�7��o��[wv|7�jKL����N�Ng��к׀��R�"�e앷�������uez��V����9�w�6�[.�@#9O'���vf��������,s���9�(VdQ���+Bu����	7��|�N��٦י��wK���F������g,�|�v�p�PV�{�����Xf��8��F+Vpl�u�ш�+���z���S�4k��i�e��#ޛ�o����ݗ��0F^eי'��^� 9 HT�&�v�r� �����R/l��ܽ�t=��N��g$>��W�n�p�.�
%Өi����ɰ�^��'���c�je1i^j��ϯ�����uw&{쮵;5��fdS�z��=z��*�x	9��S]˪��-��솗-��s�Z={	�xC"�Qs^8��.�<5ʋ{x>B�M�x\q����H�ۈY��Ybk;v�f��������L^��f����\�	�Uwd�<��  +EU��qɝ5��8��@R22"�3�qִ�����bP�gmH�][0�I2$g;�7+1K)��'7v�E1Cd�J^���sbٞL)P��6�.�ײ�G8�t����jQ� �u[�k[hM��]�p�9��ٲ�]ar��:�K� ��u��;Zb5�E��'&���k���E��k��j�Mt4�B���C�XT��FQ���mZ�ŻH��Yp'k�1�{���z��vҕ9eP(����cm\����P"	A���I��` ���y�S3W>_j7�:�ݤ/��rs�³{׬���B�b�&�6�/��?V��}p����-U��w���f1���������˞�j�l�"����K�����}ݓ��٫}+�1���d^��A,j[�~�0�>u@۸ѷnޏl'��W���T�2�-{�z��(��@{�5RB��g���c)�nG�����]����I�ړ3��TM�I��[���)xSY�\:ׇ����	����<��ڻ��Ghh�F�DQO ��UaZC|�ޮ\�~� 's3�����՞g�Upݿ�N���)z�{%ā)��$ہw:W�'����1{����L���rP3�߾��aj��uɵ�fl{���hެ�X�Sk%�z�c@�����^�S�t@}���:�s[w�����@KG�����/c�	������Sm�F�0��{z�Wݢ����O���8w�nj�k��VfW���O��J�Id� �O�{B��l�;>��K���}�gV|�q?5�5�T���]Ԉ�w�Yl�1Ҫ}jB��,�K�؟-̾\��Q���?v���^���B�@9��wYBG@�iv���P�[n��ݦ��Un�M�f�T��V�w=�<����Vۊ�����}�2:����y����f��Xl��w]�U6{��Ε���U�W�_�r����e�����I~�[�B�3g'PS�	Pu���f�o��|T�[M����X{^��h�¬պ���T�ڗ�j
�P=Chu4��t@� �ϼ�<�gh'�H_y횪3�)��Pߕ��@h�~���*ϟ=�e�R����ω�����Y6b�ߘG-P�t�OM�����UUp4*�ܢ#�^-�W�_�r�G�JgޒH��v�{�c��� �IeG2�ii.�L9*�1!]%H����]�T]L  A����H�`�!��#�K�qK(��72��t��M���C�ٽI9.�)��^��@�8����Ͼe�+�1�^��

�S��zVV�[��/@H����=-�^y��LkY�g���=ެ��b�^��9�)�>�ԯ�xuK�Ȳ�{����M}�����v�+�u�Gcpfz�8k>����nfswN����;YB�fp�"��K��S�S��)炼NS�y����ZH��R6he{ b@Jk�I֠*���0��y�J�0e����:�i��w>����=3�XgvD{ {<�7��#��:w�C����B�z�8��׶�D��]f�X�y�;���Ci/�ϋf���b���ϯ�*\�}�a>���xA]�C[�dй�i�2�jԾ��:k� �CK�G܂:k]u���s�wwB�j5O�jC�|��W����X�������)�Z�ɠ�K	�;Ux��L<��ՈI��UF�t_����Ǟ�ٚ��d;O��C��U4j���S��:m�3�-��oQ��B ���?T��7>���GR��n�pod7��dh���j;к��F��lk�Y�Z0.�]@�ի%��l���������R� �-dz�׭(��:y�����@3���Rf��b�[3HK�$3�f�,�6��M �5�a��С��͈Q��+tlu��=���V��b]i�+yF�sU��Z@�.����(��l���+5�^(�%�Ίͬ�nr�F�����k��H`�4�i��v�.n�Ԅb��GC��P��f��aL����]]wqם1���T.9@�j��3f\*���$�į��w3M��%;M�iJkFѺ�k�b D������+Ig�{/�F�7M��_m�g?�BE���2����@��CL�Z�@������ l�g��vr)�.�ǽ�mz��$����9�?���l��(o��.�1�Hyߛd����B��_g�o^w�&�wū��
�$��i"Q�O^�E`�R�@9�9��8���{>�������2��,��{q�ttH'�F��WRo�>՘�1i"�%ln��^���CT���ǣ��~�f.Ƽ�YA�@�
δR�F������I��7$ٹ�)3�׻�G푦���*���^�������O�S���x�+�Д�Ϳ������dQ>�)�̦�L}�g��t�_=1NI��˻��V���v���B��%+�T�Z�!CF�N�tO�qZ���$�,ŀ�>(d׽�z���x1�*���y�_���{]֊��.�+��;�g�.:�ϫ��Ή���a���/��S�'������ϛ7��;����&��:�MϾܣ�߮�L�^��m�Z[lcߝ>pO�v|��$��˳Ҽ�}�i9��f,[��JMQJ�§�m刧X���V�l��=��[��ƨz�XB����|��Q���|�:��1�k1w�]_ntT����s9o�k~wug܀��~`����.�awE�^V{j.��k0�c�K���D��y]�����OO3�;-.L�L��w�����u�)鱮��N�Lni]\lbܜ�W7}rL�������h�|�\�ܓ(�S�%���d�pw�T�D,�ږ��M�=	��,�Y�iA��o��.�m�76Q�3Y�wt�{TH��`��'y����]^>G8Z�M�uvE��hf���0���#ٴ�i���MVh:�
�4}۰�_M�y)&~��%l��A��+5����t���zk{v�[�P��'%O9�Ee4�Vlfu�/B�]"�J�r�¬Y�<�W^4
��$ե�*|��%�/�wgX���K�Ѳ��ь��]E8N���rn�ܯd�iÂ�A�"��ͳ�J=��+!D��t�h��ܫW�V+$
E:����w\m�G�e�����R�@7{\��9�&�j�l��e����K�����N7�w�ܧ7��w�f�&����`��ً��"L�f�D�h�Z����ʹ���u��K���kf�z��T�ɭ�����k4�d�u�����Y��Ʒ�;F�;�۽ﳁMV�TBl����ٔ��v�d������7��į���L�-͢9h����E��d�����#�r��:]�i��]�0ν�����(�8Ye�'Ƙ�(�\���m�q_]˻̀0�u���g-�~����w�����0�2Ofx�Pb���>���:���NW��yJ�R������*�
��]a|>J���}�Fn�vL@x��zgw\x}Zz�VȨ��onL��DQkQ�*��a^!�
�Z�3#ɓ��f�����{55555>'g������+�*`�T�8��5Q��DdX�Ҧ쵨�c5je�[j�3�S��f�����ooooo���~���΢j=����*-�TbZU"����}j,j�[m��*y<�ω����~?_�ooooo���~�얼&	A��U��ՋEES�i��(#�[[D������79>�O���������}E�V>R�V#�{�S��$X��i��.���NCE��;<�Fp�q��u׷�������~���&�*����-���C"(�Z�-�}k����f��٩���nnjjj|O'������ѳ׹Dպn%C�������˷X[z�J��-g��X�J�LC#�����,QUX*�&�4rب�14�k(��V�R/ j9eF �j��-.�e""ҩEP���b���2؊�U�}�E��������PA����[J���g�=�F$Ք��R0H�L��@׏<��߷��y�o�/�?�L`��0x�C*�8�$ ]!�I��Qv@���Ie5���=��5��=�<;3j ���Cq�;CGuӺ9�tz�c�t�}�~؎t�!^5�C ��{�Nȭ���xB�ޯ{���=�'M�6�v[�2cQN���=[U����\#gQ�^0�f`�� ���{G"c@�kfk�R2h��5��3֔�ý<-0�}�/�v�к5(�s��Ccr�߯���Op���n�Er��=ީ�`é �������9͘.�2&��?]<��30+X����wz�#�q�ڟIp-V�~� � �3F�^�����;�j��O<���{I��
n%Μα�������ܾ����Ͻ@���#�]�.�!���ye�4bP�0�>��퐬3�� 	,�� 媡����]��sS�O1Ʉ0�ϷǅṼx/��	�������)n�l������S�mj������%}��V������F�|.�t��]:�:G�A�p����1`C"1#1#d)!�(1���cy�!��z+�:��������w����{�P�@��n"�V���lg����Cy~CM�XxɹƓq�No�~�m~I��m���{ל�]V4n�Ԋ�Q�[���%&�6����Dw;��D5�`��)�©K����������?8��*�.���4/�&�I�p�,���n�k�r_��
"�Ǚ�-�	��L��E�Wp�����ɑqz�4E�V(^��rF� ����Z
@{C�&�3+B�P4���!���L������{�mG�&j����8.�4S����GÞ���ټ�d�=��B����p����{������	��p�F-�
*W��k�L@L+ϭ�c���Ц,-'"�k �)Ys��3��Y��"����u�|/�w���i�C�̔e�C��{:�yͫE1U\���īv�"&���H�:���_�qs����7w��,Ry�5��j)�D�>��w~�hR���}��ĞP�bF$A�s�Y��}Vh�0ރy7�k�_�:e��!fh�8 u�m�c	�Ӷ5��j�֘��8�`[L"�m�J�%��R���+W�Q��%�:h2���E�)]r��G��4�l9���f���bl���C2���P-�)��[�jv���BT!��͎ʎ���Ў؏lYs�`��ZJ1���3X���l֪X�J�cՍ���_�t�%MU*�Ɣ{K��5�t���V��e9��7߿>���O��xb�����$�Xy��L��v񝢽�'c��C�@���sj|�c���}���o�Ly�{�2�.f���$�Ha����we�I�`X���5��{޸��F���N���@�dµ
8{= �g����Ƌ9�NZ�i;�`��ᑪL-��m�݄��F�_�]O7��(s�0`��F����*.�[���:�z�A�C�>�pCIa��a�k�pZ�n�]�z�׸d�zR��}��J�Ň��R�@r7�RŅ�%�
"�0ph�Bvo^=����+��@�g_�n/����L�:Z�a/�"�%0WA��i|�$G����[Ý#��Y�ˠ���4m��cmJ8�[��E�ٟg߳��Q��m[�o�?{�D��ܡ��D{�L�&�u��_p���`O��Ϋ��u�yоY0��}�����Ü���vJ��:w�� �����U�+n���#B='�߱����v�:�}Y��ӅA:5��z��$m����	+E�{?�/�L%�R[)-��1X�D@ɞ�	���i��ۣ�o�����b�V�r0� U/,��l%�yN���K�A�S4�E�j�L��pu+��+��u����e�#�~G��`�|�9O��s[s0:y�TXo���ݹ����y)" �Z"�	D���A5*/�e�u����x�&Z��1�n�ư�W���Yu��vd����agK1,�8"�6os�^���X���"��ܫ�2v:R�Ae3h
b��L�13U/z7.W���?����������iJ�BV�m�cX��iU%�ff5��X�����Р�5� W���E�j1nb���᪡�7�'��]�g#W���b���珞]ݵ��c��p�_&r�{�?K��F��Q'��3^{�;+>�y �k��<�2w��n様�r�9���u������p)�d=p�������lL��M(�WO�O�ưcv���5�*�����f�]��(j�f�R�tH-�����8*�{QV�指^�n��Є�oB�>f��2&e��	fFd#,e�e��c Cr���]��N��p��������R�I_<���^��x#�]A.�����#@����Iv�`�e����O���]�g#W����'`��`�	W1f}�s�g�̇��ر��IN˫q� �NXH61�@xt�R1��`1�c���}����˚� Xq�3<c�ph�I0UN"l�Vo.�G�xE��5y:s�W�w0
B��1[�շJ1��`�s]�߯��%��zd�� LX�f�M �;S�|��{��t��H6�81�8���9�sCU&g�Y`���,!����\pz�
!N;
hn������9������iaN�`�U&��uy~��4�[�?v�V�G9C?K�(��Jݱ���?<X�`��Vu{�ϗ7>`_�~�����0�a���r�;�.�Iaw�J��vk6u��b��;5j`$Re��v�����͎�@k�mi8��tu��U�Y�k����8e�yN�_��y�|zY�̸׷�(����D��;i:"�;��,�,�`=��w�$��2����X�2��I��b�V1${���{`׷�`���^*�!��e�y�CL�`�M����Iָy���޻��F����O�z��l4��j3���s̼�4��p��hH���x�AQ
�Z6sf�.��E3m�%̳ke}�����EtGvr�����3Ffk��\��XW�c���(<��j�����og>\��CC�:3{��B�$����C>�C����d=��{BM,�@�>������lX[�x� 1(6V�S��矆lz��8��#aT�{���t�`�@<2a�~�D;ɝ�4!�Jw�>��[�7U[���5��t��1fG�!i��`�<��K�%�(s�b_ǇG_�Ӓٵ�A�`
�' kv��������Ȼ�`Obd��pXOo�q][J<J0n�{�rXj�q����ٮ�ۣ����Ie9�^W���3c����&q39v8C
�A��p:�6��k��.�5���S�;��VԾ�p~���ȡgl���΋mk�42}{{]&5�7��j�h����;�t�~��jH���@82����� �I�P/�O�Cw�ղ�Ƭu���#/�<��QИ-.��\m��&rw1ٮj!v�I�
VR��&��R ��yum�!��"W��.`]��cJ���^���o�� \��A&x����q�vҌ��i���6�h�atl����}���e�
�؄šU��M6r����ˈ����b�����%�HKe�FV��$Ɓ�C#�uS���������&2�.0]�Y��Xݮ[A�Jm��C�s�y���
\W�K}���0G~�����aXXX�=>�����<�ny�pv�K6��1����a�EZj8�!m���Dk�6}�M�����Oz��$�'��,1)b1G��*��/�#"���_�� �&�&�P��3U�8�~�I�)��a�=J�y���,����e�@	��k�U�G�����ߴ1)/��{toFC���a�l<��>��\��JMU�5}�b%XM��1���]���L:n�A��X8~����y�N��p10�XV�Ń���؎r�Ј���/y�i�J��r�谂�0�3���J��^c�o��>�9�p��y^�gdd�ט���L �9. v4CK��_�7|�u�Q�f�l�b�6SV%��+�M`+q1�`�:р\�$vO~o^���~��d�8�T�]��������ߟ��p� 5 �[Ǜ �K�2;h,	�L2ń�N�8"�D�o6v=q��{��-jߊ���X�u�/�n��M��<3��W�d���/X ��ׇ�����j�?or�'}g��X}���un����! ��"HD�a�XdĢ��!�8���E�j������z��³;#d>J0}�n�����Ǟw��óvmr�D>�=���-�ѬH�$�ఄZ�=s��"z{/�}�7W�,r��F[�s�b	j�Y Rq0ä蛁��'��0�`�i��8p[���vnb��nmzc�˰�xK�H(p {�I,<����9Ǩ�x�������=����l2<�;���G�_���1�bb�y�>�+{���g������@g��Ȫwi����04[0���Y"ȱ��:x)�t]l��1�k����f��m����|��^��d=ߘ/�P�	�C���Q����y���v���_0@�,1��O.m҃JY�S�pXU&%��,֭^^UH�Ϸ5��u0��L1��x�C�z��G_�Y��&h�ɏ�3U M�"/r[b���o1GP���rɝ�8��,��7�o���訆��@�v&"�;M�nd���3�һ*r�fn����C���o&�����mc�C�E��(�a�Xa^B���bA 3VA�o���|/3�-��(|�`��s��L�h����Ia3{)�w[���fH����b����~m��s�ݸ�f�m�^A1a[&�wLMb�5��8C�^��(�T��a.�űh"�8�F��`<q�ѳ�j�㯗Y��.�@F� �G�av�� � 2E�S}��߾����E,&�C����R�n$�֚����Ԛ�cߨ��qn>�I�����0��N��,.�����|/��s:��������6�8���� rñ�F1a�4O�T���עFi>����>:N�F�@�Zń� �#/���Y3w�-L[��H�హXŅ���~}�O�b��,5�j!A����,f�R�w���ws��"��6|�^3qz�πt���LBf�H,	�I�S; �Xfܩܭ%ޏ0h�X���X�`���������&�A i�O�o�-��1�#5��o!]u=�_4��-�\�/k
�sO�������#�����Q[i�7����Z���
��|��l/Ud���������C!wa�M������˦

��XQay�j����E��g��6��/�����&n��a>L6�u�,�d�f;�^O%��.u����?���s ��K
���LWh�Z5��Xf��?=|���b���G��X~��`�����0����|��7�v|����k.�Y�]܇"7I������G�7�����cm0r6�G�3Fx�s�"`G��¾����|/�e�gH6n�;5RgӁd�vrCI=}��e��v��u�����cT�y6������7|$�<�qus�ID�2Nrͣ�z�&�h#Xx�p@Ӯ�����2�f��7����t���K�B�^�ٻ����{_h{����N�{�dD�~c �dkȤ��ukZ��_����\/�]�:�� I(ש�G�la8v���0`!�bG�8��X��{

�B$Y�a��j�Yݶ6��G�Do8��i�򳽏3]�o)s�@n�[B�n���&�|B�VU��Nf9i�w3�Na����lX^���xV�v1�f�<��J��;�ۂ������6�7h��^�81���<�n��N�B�;��Fl���1eX'�*�[�fp�U�g����f�V0�t�Qf�sW �M�շ�oTd嫘�m;�xo�r�vͻ�v*��Z��e�=�t�gQa0h�c��wj��I\�j��s0>�$��86V&����q����纝� *��0��7�f��}a�&��D���J:��a�4Meɵ�]�x��>:�v�k��t�H)���}S2���l�W�n��w|nc���azgAJ�4�ӹ����'�������(��3�%���N�]��X�U� "u�cT�cG*��ۛ����q�8�W2w\�3��"��^��3L �y��Vv��7�*��Y8����~�wm]��fu�v�ñuv^��wGz�Q���cG���\,��m��e�F���\_7`\=�J�)Q���{�}d�a�w���m��e�_oW��̞},ufE�gbZ�%��p�|�i�GÒ n}k��% Т �|�JC%�s/b z�e
pۡ��9�hE��M�8�ߊ�
3m�+��o�E�ɤ��*�8>���1Q�6X���<Xic��~�R|c��TB��� a[˼&Y�6��8�'�����1�bU�֦[�U)SH\�Ŋ"{J�E���ƣ>�?]g�����믏��oo����~}۹z2����Fz��+�\���ܔ4�5jyar�S����f�����};77777>'����|>�낈�EW��|j�%���vN<;B�3�׮?��>>��]~>>>>>?G����{����1&����b�㏉�L@ѐ����ֆ�e6��(*��}~�������~>>>>>?G���|���}ȥ�D�{Kr�PZؖ�V�rز_l<��O�4?_]u���������[��kx�to}� ��M ���ޚ1j�3�k=�+c�-������/c���o�������u����q��T����r�[n%���*9e� A�S��Ucd����!b+�Ag�FTfYCN����QI�T���ڠ�"+�EeEĮ!�P\am�jQ\��[���8��.�82�"��t�f���
-bʌDb�D�u�1Uwf3n�E�*[C�wK���<J�ӤKeE���ӥ���9sm�H8(j[=�Z��
	�Ë&�̰+M��˯Xl;Y����uA��YI@i����Z��p��CҌ�io�[t�Xukg6�M]-�R�nn3R%ib�]t%�Q	,iٛ�5s���S2�z��E��n�b�V��ԡ���&3%�7QrYm�X��M0�F$h%\�Z�R4]�m��b��%���c��̈́)-E�i.m���.s��\e@�9��b��m#����@�r�cmҵJB�l%f��okL���j6eUD�5[����eԫ��B��ci����6���,v����޲��%�D5HM6��Ñ�GWU�U��j�]1��ڦ��`1������5q�S�l昄֓\hō�fi�uf)�ۜ�i�����K/ ��mDa)�VX�]��efic�#�H=k��\�
��p�ȥ"í��7)���c��i��n��i ��5�`ij�m���F3[�+�9��X�Q��#--��6,��P�:)�Y��̲���e�2R�D�ґ����4��3m2c<M����X���wE%��� ���燗倷$K�Óڲ:+mtk�ɹ����{�V�wX��#Z�0]3�ѺV d�e5���2hf�^H]X�!�LmJlUͤq{	\K`YD�����<��|U���F]�Ѷ%��e�6���iU��Q%!H�t\��J��ڧ--��(�L�ɦ@.G�gC�5�ʍ%�i�%��T�ݛ�
�D�	�jJ4��9�[-y�[&�-�a��VM�m���d��V(9�)&ѓQ&	���1=鵾� �HҕQƪ�n�3qr2�.q��f\�,�Q�cXQm�]e�� �Y�-�F���m�k�`v�C�m��@�v����ֶ��4���bcv��Ռa��i�v)]�jD�#4ڑn�`�����fV;^t�l�P�:\�(WK+����͢�.���k���ƚ�cx�Bk1�^{R�gA�����ZB�_�@��Q�@a �� R��	@�L@���;��o5}���w�裉�lk<�¸��[Y�L�`���չ;������@�
�`�AZ���1f�2�[�.m��&-���/	m&�klN%�ٱ�1{5l5�ʁ*�%i���e��,.���kvV�#�M�lݖ���4 X7�!��aw4�1��7��M�Sf^l�t�cWz8�7��Q��A�stit��H��dw���<���������.�e��q�u�+.�WA���	q
�]�à����P�x�߆���,�Rp �'������g&�h���y�e� F��!�Q-�Ղ
,໇�N�Z2�벉Я� �BB����Y���f���v���	�NF�b%���O�wu�{|q��ǁ��6��۸��=���)�p��鉔���@z[��6;�N��~Ǯ��w~���~����>�:M�gu2u��V��v�C��|�޴�܌i8 �jc���\�s�_���᳓w�$�>C������y&��޵`�����j�+Ĳ�&�� �&���������{�L�O�;^t�L�r4�H5I� � &g�:7���}$�U�{�^�;�\Dl��˱����TB�P�%C�W@��D�3AÒ@��ͅ<�^����`�b�-^�=�|��x]�S3{2���zk�9`G��똄A��K K����(b�g�m�K�`�~}�N�]��m�뽽�.�z����j���܄±�B������};3.���'1z�f�s�!�ְ-i�6��Q�k-���0	�2 C
0���� ��H�Q		)��#��2�}s/�3�龍nM�-e��A�"�ρ%A�8Tw+S''��}��R*�3��%��SB
�g�����K���+�����}gkΗ AmL4�nQj	.n�A �8�0n*w/8Q$a�	kb��3!S���{���|&�̒�N���O�*K��0h��yc�	��C+�����݊�&�������5��g���^�y}�6��G�� ;\8���R�����E:�u�=��:AC�xNf��%�f�Ԑ��X;(�ZL$vO�o�~���q(���f�⎧��o2ƼJ�?s�ȼ�� 5NѾ��[¯��x�BNAryh�����##Z�`ÁT�����@7�;�;�u3o·Ps$C8\��5Vf����7}�;�-m�@,E� �"�*��7l�[#�ӸI��SI�A͖F�;�J@�	z���{^�G%tl��;���[
Ė�����2l�KK<�zHY�RwnD�'���=���
"���u�<�Z�_6��<Ýu�£�U�Ⱑ��NHQ�Ua�'��^�Y��؋�
?H7�8$�'K;=&D�8z�Aqo�f�G�5��A:� ����e��5|���v�tw��pD��R�;֬�������D� *aͷ�Śi�2DF/1�H���a��X�p&'�
�U~��Ow����S  ��y�cB����I�@�{�Q�JK�O<~��}�'��ښatv�fq�%Ԏ�\�,�+fa��M�����߼l�6����=����d ��41�@;dחfF���x�AcN"������L�5������5	"�]��bӌpIB��Y���r��������7`�q�u�^t���; ��PE�RΘ��L�K`��񠃇��(�s�dD��0�/�rh��;<��G�[���O�
��$��%���s�`�9�:���Q��\���������X������j���֪���s�W
<I&��t��Sџ]�VՔm�#����<�N��enǍ�ލ���p�r�}X{H�,a����Z���fm��G�$A!RF#+��Te*SYNҺm*6��8�w�?�0�� �|a	H�#	 �O��K9�o�Yĵ�jɥ�w$���s뺬�R��;yx]���t��Ё�NE�A�$�|NA�ޚ�{�vǰ�ׯ��U�����"��5�a�&p�(��P�~>~D�����A�w�'�^�S��1;�k���|�xp����8��Q���@��d6�3y<I%�7�k�;�20�<I C�X�Ėi��H�ߟd���ZYL�8ɮT�6;�5⭸Y�-���$H�;6G�%�;�-��x���m�7�����oy�D�~�pܣ���Y�Gc��W� i��{�\/���o6�ܥ�⾡�]
�H�<獣e�ao7��_Dq©0ryÁ��$���;s�Q\8U�2\�"O>Q�/�r'�[��~U��w�����E��]��X6�jD�v�j�7=%��>�z�c<I'<����c�,h�8D�n�Z�q�~�{�]e��L�<"f�w\Y5g[s�tR�VV���v�.�B�i�n����}pvg�Wekj�C���S}�CG?�$�$BD!�_eN�¯RR0�
��~�n�kJ'im��ǇƠ���
�B&��tl&)���c0��X�$J\��s.�l+�lx]���YA��͙`�m�y6�k2D��e4�auZ��e�����60:�6+p(�&�:b�L��!�Ua��f��2��Z�T!n��*�F��rZ�3+`��40��s
VMvI�g���l���A��Ͷ5�:�-u��y݇��/��'�і<j����V�΁��1J5�؄�W����x2	?p�8pX���y�L�
�ƒ ��ݬ�ًs�.#G�3G��4bpG��ܒ5H�Aq��d�K��>������� �g@�|���(�*�!���U��A�.��{0H#�C�/��>�DG������{�Ȧ�X�v��k���hy�z;�5�~6�ԵOeg�a����0z�li�d5����$xu=�����9iڋ@�m�>x�̍�t��LX�}�#����=g�\E��<�F��Z"���r$���Dzz��fx�5�����������WwɈ]��.�H�>���,�1��EOyxVp�H_�O���
��T��-#)v�f驅�ɚQc���ZC{�}Z-ģ�~=��{����^s1�N���_������ש�%ې��s�S�	8��Sy!߳5W�B���F�4�K��$aD��^ȿ.ئ�<�����ŷG^Ơ����o��ws��b�s�}�*��OdO'gb�4�8 ���Մ��t�q
�g�C�z�����k����5���5�4�M����wo1K�����s?���Ԑ��	��!�H�s�/�I�Dd}��s�3>�̳�������f\n�C�� �:�ZY�]�Gz��C��j4��tϥ)��]5hu��綥���TV�
��Bp�\��M)��bw��D�̖��k\�1��u��k� (pG�(���E�36}v��g�'j'�iP�&���+��d�#A�1��@3.cfD9��:��IH@�v�UV`�{]�uM	6���&SWW������:\Aʓ�`a��s+� ��w���
���\Dv���Q����c��nV���h��abZ�Shci}O^�߳�=��`���#��c��)@$U8�8�����W~b��.���<�����'��Oȍ9�,O7�|���/|��"�N���vtTް��L��@1�ǧ����z�v�xI�����-:eD>
Ғ��9}��]8t�wC�H@��NԹ#Z�mܷ�4z��M���jBV���=_^�^A�v��(��n��f�����ES�ȘQj�zH̟d�2���u=�u)��@��TN��Y�z߸z����H	��	k�$�'n[yp�B��Y������Y��-T��v�=�Å]�$�(�i�!۞7��rA��A��2�Q&^ظ1�k021y<DU�$��O��Л�j��v��:�s9n&؆7��B��20�b��s��?~����~HO~�>?��������9�Q�2�iSRB�MD��-a0��?y��b��FI ���q�D��B�n5���J�Mf?���VN�:\I� �ӛ���{�5h��n6'9t}�:�r�IQ�4��� ��܁����®���8�1�x� �����f�"n�d{M�i6F�pA@zT�1Gڜ[ �L��rH�U��"�0��w����=F<�	�!�m�����ZrX��CN�4	�-������=�p+���!��fz=�|+'w�s�&�݈x����u�YȪЧ�]a(�����S#�-(=�m�LDs��2�y� K1i������+x̻����w���S��ȧP~�m��H/����`^H�D<��` �Da�~�R B��Cl����R��y�f��fG���X�^H�q
���4��쨃�h.�g���M]�b
�xb��D�U�rH�w�!1j-��+w��hfm�H���~O�֟���]4�1��A�z�j�KaJ�P��m�O����J"��;k��E�K��u41�RZ)8�6�ۢ���Wq��RE��A��$M��>����9̮]r�7Fsfi��Q�|����9��{�3Ȗd�'�@}ջ�>²�}��� �'�N�-�\kssc�u�G �`�0�P�LA;Ƀ�H�v� j�t��㼹�^�c����7�W~d����EyÂ*�r�fM�X���l:~���眻�d����UѸ*��Ex9�)��@�;���0���m� T��A�t��F+ݑR�bM�v�{�|/E�n����1��Y�;:�I�LQ�X{r�_?�~��2:���T�o(��AS{Of^ާ]�CoxtXҮ�`Q2���:+VkFH�(N�Y��X~�oG������޻��#������n�V��ȧQ��Xe^�x0P�`��L���[e*�30�uf���2ݖ]阂hJ)i�EH�.�Tښ9�L��[E8��MF�b�ec+��v)-�sa�WX�p庀FX�bi����]F5J��X7%e�+���mIy��l54٢G\9ш�<���B�٦�h� ����yu���m]Ĉ�zb���؉�lk�=����j����)h�v,��`�j�nϏ�������+�bjmfҖ������;.uv�l"���a)˝��A�U��1��]�~�{��o�����w�5�E���������b%�Z����2')U�.0&�^�Nz�L�"PZ�S�b��=Fn�i�����έcB��^T#�c��ł�>�Ip�2�.CA�!�����p���b3�궉��g��xe��9@L����&v5I�� �l��嘖����	�a	��8V��le����k/�ulF�3�J]� 5��E�g"Jo7��D��P���Mӆ�DA�4��1ro{Ѭ�t�~>����+�9��-Ct%k��D�wU�Rpb'�γk^qw�����I�mc�j�;�$���Х0M���`��>�[��m*M���12��qa���*�ڋo��;մxe��..g_��[���kg592���1?2aE�1GuGg�P`;����s^�J�t�r�Q��%g�B%���h�u��/n`��[z����u�V�鸯����K$̀=tY�n**��Y�=�����E!�`���"�I$�a!��G�����]��9��!߃�Y�yÑ��W����2d�)A$����H"n�g!P,-2�N��t�CՕ�!;9d�]nU��z��爖IjA�q�l�2��DZg0�{H��u�9� ��H9,�dq5"�ݙޟQ�[�t���v�ŵ��^�g7Yz�Yio/Jg=j=i S� c���A��2�*�`f�+Z.V?��<#�ʖ_�.pN�d���Z���DdS�j���v�J��]�iF��PG2���9��iXؘ3e}O~�-���y����$9�u��Y�ZqYF��j��eps�{f�W�<�
I"�>!������N�z��ُ�{�3����)��b56O�3ޝ��.�|�Kc��9jf�\�}��K��ڎ��ԭ�y��0sT�%,�s��Ԭ�@�F`�0{�r���L�E	K�g�/B�	gN%��z��`WZ*u�L֛[ v��w�ǹXh���6��,̤�:33�n��>�zqG��N�t�Y��n:��Z�`}N]�ڥoh|�f�����g;�;��^��v�kw3hee�%ei�ӡ���T���e	�J�4���������U��e:�Mȶ��Ҳ�k�j2Au������n�S�)ӷ]�]��AY�1�lfq�{s=׸�]j�Z��8�jx��`}zq�op��>����}�-a��E�K���p�7�Z˿-A�o��\](~D-�;ﳮ�����e�ͤ�o:5+�ϟ�~��+�n�P�
��ժW�W�3�!�]h&�λܭ�[�v;�ѧ�辬�.�J͹Sn�;N�tP`4Y�Y���U)�CÀ��ܗyC;�T�Wdu]޺$Aϥu������34�i�a�l�YD*�ޝ��������t91��^���@۶�R�~vqYs]�3@ڻn���g�]q�0l�Ǉ��w�ApYٽH֙��	�ȭ���wVN��vJ���Q�n	aa癶�|���d��k3���M�\/��y�aX�5�Ȣ��t��x��<U���$����#μ���"���t�U�n�n��yt!ļo<�>��W���a��v��Z&��.����0[�kg�P�6��0Ų�рL�����A�I�N4��JpǨ�,:��6��땞��*��f��|��I}X?.����rS
���p�sJ��HAھ[���&�bLCѷ냋J����Z�|Lr�L�cj��Z�ҿY���;7>��7<�O��S�sss���u�����&��8�����"����w+��"Ņ���+�����<q��g����}~��������*��lĶ�m֭k��U�@�%�E��\q���l��X�waUQ�Ƿ�=�����׷������>�ϧ>>Q�*e���6k1՗W�6�5h1Em�����rZ��^��O�6M���'�S�ssss�}=�O���.Z�YJ�iw�����gZhi�K�`�+"���Z��ZS[[cy�������ͭ��o��F{V��F�CNaAIR�`%ƊT-�^�eWB��JS�������~�^ߏ���������^�!���9jL*���xMM0]R�*8Z��U���`aS��|2İ)"w4:�<'KS�͸�,ף���C�t:�:Z�lE��E�CI���V=iXj�l+{���BP���2�x��P��C�����r����G�V<k���F��+�%Cܦ�t��(@�)e;���:�3��U�C�M53*�g�~" � d���C��=dC���	��!B<C?/��N�/yR��%�pN��6Ƽ������5���d"1fQ���*Y2m�^&�7i�ª�6nf��W<�oPpa�w-ꂣ��8�OyC���4��th9)�4`�R�F�����~��ȷ�k2d��wz=G�]n���Uc;@I�*��
dT�H��!����ś����gQ�+���L˵t� �4n�E���h�K�߾)'���jq	 ��l�DT�õ�g?����gav)�1^�n�=��;b3�}���D��{ۨ�{˂9���۬=�6�b�Ko ��6.b���x���8bBd3 Q)��p�B�����=�W>�����pȜ�L����<��i�Fm]uǨ�˭�t��̪�F������8�Đ*�3��e/1l�a��Hv$��э����xt�<��!.�$���k��}1��y����׫*=�4y�Pv��@w1�7Ȏ��í���<C��E�SD^���R>zk�P����A�Da��a�RR!^�זxv����ry�|��h����n�iX��x�	��l��О�N�ٱs�ips�z��d�^=2B�Z�mn�|εs�%��;bD�|}��}ˠ��lG.R�.�B`��5��.�@�X��o�o��-r�>���?L�����O<�!yvfy{h�˝� �q��s<_9��z�7��C8E�����S��� �y�Cgp"�d˹$�,h2B�	�c�_{ç=0����+H�XG�L�]�N�xK�`kb#S&W	 U�妽b�&�U;�r�R=<��^���EA��d\��\�ר8x�EQH�s��9�h�<󏗳�J��se&v-E�O^���G�^����Ab1I؏vV��V�/���9l���
)CZ�A�̇`M��y�:����[��9�;HK�t�D�,b�oܩ�7}�Td(.L=�<�jޟj:�����1�q�k�|'m��)��<Z���ײ���F�8�[R�kw����{���Q�?*� �(~C��9V�U)P�~�ˇ^wwҵ#+�,�3T���B)U��+u�8�Ș�r�cYi31h����k�3V�s��4���Ku��"�q���mQ%Ŏ��k�����[��������]m��K&(,.�n�Rh��)t ⩈�b�֗d�*]�鈙���&[�2� �:i�%�:��K[bd#;��2Mƻ8��CJ��-[Xf�Y�i��m�տd��I`��]�顒�r��x�1�HƤ˴Р�]��|�|��[-����Yg�=�-$b���F�nzNd���_q�����z��<H�n<�w���A�zcȐT��rH6CC�/O]��$���gٸ}�G�^��%lG���-�vWiC���>�L�k�v�x�%�>�L��p�h�ER^�����g.{�T��!.H@�>vES��
�0P U�}�^lǷ�z�� "��@�fӍ�5y��1}Ɨ0E�ޠ��wzf,��#%zt9�Nh�|�#!;a04�3'B�r�|�'xb�LB���Y�{h����$��I9b�AS#H��6sIɡ���{".�=��g�6W5t)AHĥ�4�P��0�6�T\r��e�����V�(��B&����������ҍۍY[��q���i	&y7#=��Ռ<��0O�32',��(o���X`z�O�;�glڮʈ�x���
�R���W{a'}>��V�̣bY)�^�=�ޯ��rPz��&m��:���5t���S��Ӊ�'l�tk�{���?�}��0,0�C�/<����0°ȏj4�D�w���ԙ��g�����ǭ�������A�2�1�l�y>}�Y�p5��v�̸�41���Z[X��#1���g�����g�´V�o�\&�p�D��K�����ɹ���`H�k��3�9x5�S��é@��B16�8������vl�"v����%�ٷu��!ٞ�턎��&�J��375f��Y�^i�9,X3�R��*ݰA����ѹ����;��*�W Ɏ��6������N��՗z�MG�DK�e��ͯE�Lg����y�NX�2��~�%�:y6PL�{f* ����ؙ�g=;�Դxλ�쓽z�bo�I��d� �k�� ��1I�z8����~I~�D����4��Q���bf��`����nf[�ϓ������"|����٣S���6�zs}���+r��.*�2��T�s����1�ۂf����#�[X<����w���~:�LD�[�^�����3��%�� Ey9U���u����>���;��3�c�\F,��^��lH!-�=/�bf;���.p���@��J��� ��0&�<o����h:Y-jpN-��j/��vȇ��25�����D�?(�:^�^�z@�ae�z��O~�_*�&�>��>����o��p�1��qN�M��tvB�E��pAo�D:g��j�����
̭��u�� �'���十~�fy�~�Aqf�8ɓ�8��͑����}J�����+��p���d�.Xig�9N��Rm��:�C��\�߻�>N���%9Q��Z�8c��\���5��*m�~~����:ō�~V�F��b�M��@�Nq�18��3*�lOY�>�� F���&�Lt�9qñ�j��Y ��p��<Ď�UOя�	$wp�#֙�7Ue�����[�@3N�ɦ !���]���9�Kmy������Ff;Ya ��W.�gMąu^�ٺ��V������_�8"�3�A˂Rr�|��������	��A���ql� ݧ�Wz�c��I���Lǧ�k(���AFb62��U��fAr96o��� ��ճ�^i+�R�`|��0W_�9��k7�wv��+��>��w���M&�͎��0��$?��˰<�p`H`!�z�)��
��s����������$�	�5OL�I��#����D�6��A��`���k2����j���jL��'D*�L����,z��+ԕ\���3:�٦�
�ҵ��+n�c�vM���Y��c@�������b��`"}���ps���wI�
�����+�q�s�D�W�-��?���3�/�3�s<ˠ�nSb�׎��⍈��c��B ��e\�������|9�Z���,�����o��0k��%"���pA�f�
��B��:	��[C�g^�g���eo$��"mG�����X9WjZ�QpG� fb1g����%��D���8[���wQ�9��`�c�
j�����vQ|�V�>1
�;8y^܈��9e�9_=�8s=��>�I^I���vZ�>�֡-�`��k1�)���2޶������!ܢ������D���l9z 2�f�\�(�\�Ç�CFORk�44� �y�O���6��#RC�H�Q�#	Mu"�_�_���>L�=-�euVف� lh��<��j��3,��a�¼�R�����f&�Xh�%+L�v�v�(�lK�B����9 K!�RVJ�[FQ��g�k�vZS@�lWm��J��2��Qms�kt��2iF\�)���:��vvj�]r6dю�vk�K��̓�.�fԊ%�bZ�lfM3	n�m+7EhR�T�u��=��C%�.������-��5m3ZA�lkD�fصfn3�'�7Ϸ���e���k��
����8@U�1�&n�L���t{��d�$�r��\<��K��a�YG]�p.Nx����C�O7t���Ң<��N��[���*������PpQ��1u�b;t�5���� �Җ �y8�B�9�i�ݭ��X�*Ϲ���}�k#rפ�@�5�8�A��D �
���K�n���}����,G���&�8�,�U[��;���Amx�b�=�Lp9����ɡ�]OҜ��NJ\�L�Hm ����Bոp@�%�.�enEC�6�������_Q�Y�B\,4��N�	.:3>�mM�$W`܋��4K��S���mv��!8.��M��>[=���bYo$�&�C���-���|*��?��t�6z9��[e�P&-ñ��p�m��ǩD�o��}�M�xfl�\k�0���l�A^y_�V�_	�����������wsy>��~Ok��R�cO���̋�|NM%�&�Z��O�0=e" �*JMP��	$r��R0��v4�eU}�}��'|�K� ŧP����Z
n�ݬ s)�6��33g��`��u%Nj��{g<'�����˪����j��BHp8@�/zIW����5|�4%���-&}��brH�OU�����Q΃�0Q+m�@"^�����w���$���w��d	�p�E�1+r����N��ٹj��Y�Mg�8���{��<���-ޙ0Z�����z��1��y��:�� �P��$[�����ZG�R��unX�+���ӣ\�Ҵ����������ڋC2UI�k��������2S���y7�瘸� �|��5b)!C*�CE"�Xßr>�}+�5��N�g�k�M�ޣ�ɉ >!����9�)>��]��V<�҇��q�)$� ��흮{�D�ܲnD�.��4�Y��L�0�/'��:f���ӌ�ҭ��W����?9O�{���;�G��.�=��D��_�"��1�Xa��d�0�u4��~'�}����{��I|Z�9S&0�Oɦ�&�4�CcO$��;�:��@��"�p���o������
�v�������z���Ey���2���) �������E�;&XY�O��5�i��s��G�s��\��I#�p�DU }c���<=F�Ӛ�5`wN�;;(�L�fn��aL ����d`�L͛�s���mZm�҇�����/�D��UHv��SY�����]q���_���;W��oN��\�c����w$QLZ� ��9��C�>!��������W_#�Y�A\��!1<��"�DM��v����m(3��r	�N5-2cv��ډ��;
m��F՚u����sB�`�1v�)�4 ��m�z��E42/�)���	�.���Gem�>���.Qb?��3p�?]����tьWD�q�*Z�O8F�Ɨ�_V��٪�p��Dו��[\�o��;6��5�缶94��oM��*#�7�b@1�@�d'�bL#��L�����^}q���u�#��"'{�<L͏Ps�l�����W{
����)�6B �y��P�E�z��Ί���������Ԫ�q]��Z2�1�ՠ���&Wd���B��m"@��O�yɆ(�S�&��y��MG1;v\��T��s��E�*��+[/���_�R���y�9���>�8��S�,��2�-L����!uU�㣲��_y%�b�;jd�HFM�� �o&�~MI�ߔ0�rq5�J^a�D���r�T����0=z�k4b���!.wb��.A^vi�I%�T���2��+u&"�`5��� v]+�T�\3��G��	+Pq<�'v���/����T@|��
�y((����q$M����;����Nz����}�3�h��״�9ˈ��@�!��}�뚷]��:�u��_�8)k�.�V=�Ja5��v�R�<�8�]�a����w3�Bk����*�oe�e-ڙ�`ч#�V��WKm������fe�S�D���:��Fc�K����Q뽵y�2�Vp�g=e���3n�4Η8fl�aTs(���e�����<��l��/*��Wk���V���d�\:+���Ußz{7����]�VY�����]8��I��yn�7
�\@n�����8�RҲ�-�ꉌ�78_��fƺ-!�c B�۵��ev[�)��Yo3U��Ap�R��Zi;��2&�h�f�����:?w��kvvcb_.����l������T'w\�Ɋ��[x�Y�wڸ�5����s��^��:���[��;����nR�1�Mo��+�,�÷C�=��COHE�"ά�b��բ�2u���^�l��u�n������b��v&G-V�˥Z����}NVoh�Kn���{�ۏm�݀�{tOe��{�5q\{�Gf����=����Sh�MK.�:-�]��imM<{���j�T(���b��ɏ7s5,�n���!CEb%��{t���;;�&���f��Y�˭bo%�ɐ����R�c�o2�RQ�z컥r�f��ҽkif,��Q�p'ŏ��+�L�D�6KhGx�7Ϗ��G��xY繟�����8����{��e��z�2s>���{].ph|��N��)
f��nэ�d�Yt�Ŷ����)��W��^N���^=|9'��v�ED-�-�eT��7��
��[�b+����'�5�]e2(��٩�3sq�N�'�sS�sss�}=�O���u�Ar�%-be��C+f8��\B���c�Ky�h�jv2ϣ77���{75;777>'ӻ�T�o��Me�a��E<CQ/��͇�b�j9{�n!P��q�	f������Ygќ�ű����������̓($
 ���0� �tĴ�b6���z4C�m�Sժ)�"�`UC�̽bX��r�>���g����njvnnn|O�O<o������Ze������9�b6��
P�6�݋���`�R��p���e�FnnN>��_ߏ�������8{WS��:юfc�U\�M+��5������SMt�,T1j����Y�g������|{~>>>?G�ש�(��
��"��\�����.���r��	Iad��KPF�� �ھ�`MkyX�J�0�Y�V�v���,�QJ�j�R����$��pF��1HYb�K(WXb�1-����Ɉ@�vL©RU��Y��4�J�Uݱ��NOy�Yu�M����d�0���<�7���U�gb�p����q~��y��\q�R;͛^)���-�ި�O;]*�E���Ys"�"Yl8Ť�iB���ᰄՎ$�ÓHWbf�����j��j�5�B�͋E�k\4l�]
ᬵ�.��m\��[����t�"�[S��n2��8��ͪ+�����-ٮ���e��7�.�y�-0Pҝ�Ԕ����Z\:if@v�&�G ���e���SDf5�j�t�d���-eu�!K3J�Z�9.����3�\���8�ܺԦ����j�5Cv��i�ٴ�Kc!Z��dii�m#m�ZV Y�ُd�e����v����m�cJ��2��� �Mu�Z5q-W6�MMʰ���!����j�75�l՗X�n-45AQy�qt��vMepKuq����cDغ�]�q���.tR����A[In2��d�m��v:F9]�A�r�˨Y�1-w�5pVl�`-���[j�E��Vg�"D��b�)���Cam���&ڋY��B����b8��mָ�̈́M��n��`�5ڙ4��ˋv��G\V��ꠅ�F���V�.z�Ҕ�Q@�gg:cNx�kJ�v�FRL�lt�F��m�������*9� u��K.��k���%��Ƈ(�WUj��#�yBG����$�Y{8{D�R����ZFm(�5&bJ"ɍ��@v�cŕ�ى��(�,F�![b;Z�iGbĄΕul�̛���Au���
k�����YX�ـ�r�Ɗ:�F��ͫ�cZ�HX�6k�cjJ�ņYn^j���,��r�`���-6�5�Į�G&j�ұ��k67��-���{{���Wi���`�Y�M�2����p��c�,��Xa�3�N��������.�ǣzu���ZU�5���zX{�6i,%Ś���a�I��6�U������%c��]���)ͫ�}�1���tqMQ(�f!�ݺĆ�kZ�M�Q�6��'�q�t��%8�`$A"V��[+���	}{��Е�1����P3ʡ���Wb�Q�-�,��kF��l]�
L��4l�8��e�E
�� 6���jl &�g�B)օ��0�`�$�u;&YM�¹�pm���� �2�sx�3�YaU�8�p���
�e����7��Zf�j[Q�m;��ٝxrE٤M`�`�-�Җ��Fz����?�@�;�m,c���5u��噗`�n�*�=<���Y���1�|�'�K>��(ث��۝��#+=�$�����پ��H@�q�Fm:b�N�$
}�g�Ej�:��:�E[��kP/)��O��Y{N�]���G�$���/1sDd�h1J����t�\/( ���)S�"�5lm�W�7*��V{#_y%����56��Ryeh�<cDn�(9iñ�4�*p����uw����%��B�%Vhy�)������2����񻎣_<���#v��]N[ɏ<�LN .}�����{9�2����Y�S�zcT[�x{׽�C��g�"��p��a@����f���#R��]�J��?�ߧ�߿2�:2{���d"�Z�wj,�9~ョ;c_|��"�{U�@�I�ɑֽx�A1�E�� ��AƲދ��9ۙ��2tt@��΋�������`��Ӹ��ܛyg�m����Y�ދ�&v!"
��u-��q��هQ$|��A�D�)<����%���0`�ޏA��p��������^^v�������S��>)*�9�٧T�[u>2�/h.�3k�oy�E{|���sp��2�\d��A�K�A<�<��b��n��8�7�4�����e�vt�YoL{}�M�ƾ�x�w-��S'c��#�n=�r\�m8P.(��T��DB�z��.2�Yb@׻��_/+Y���\����	M8t�X�g��l>�QP�F ��!ϡ�Dw8�W$h�9�K�z�d��$�'uM�$
�ı���ݩ�6��PX�U(컧������G��w�}x�Y�X�SX_#���%��R��%D�0�00�6`�8�Oo���,L�/	`GRLC�d�^����.>b�P	�r��@h/j3�e����p�=�h�G]�����П}Lzϣ���/(3��i�޸Mlq���%���|��A��pf.�*}����)������w�gVQ��?K��@@]����H:X-�H��f�Y���) ���*�a��������̾�
���E�8pES�I�$�v�����.�
u-��oZI�,��Z�@��)���{�(ۿ�m�Ğ�� ��B#�0	��"#�s9�A���2w�`��}�������H�O{�����:��1ŧa��B��Kwyr��ʵN.���h.�'�+a	��bB�4�im�gC3BCv�Зy����$�W=�k�( � +e�4B ��A��{��U�s/����8�etFM�nBε�n1L�4M�-.�H.Ғ�Wr���3�Ҧ.��iT�ݹ����S;~���㖜�A��8&,-�D�-Qd�,mA�zT�
�cH6й���ؽT�[�n;�Ƕ5��\Ac����(���:�W˅�:�G?���S0�:��\86Bc]�9������9��!.�P6Bb-��R50���{�c:�u�7�o��O�N�"�<�4��73.܊wa-��7r
�[����n)f�oq�;j" ��̤Q��J'�������d#)$J�! ʈa���N����e�~ ���_u4���-�CT�}7��C�0e��˛�������>����DKf��`��B�u��`��uX�9wK\ �l
�WcF�)�jˬŦ֓WR�:��7)x�/g�����*��ȊpᨆM�5���E�mk�nwMe*Gk^��.dL�?����1^M�����N��#{���?�ۉt>>!42������v=ze�HK�d"����Rx�o#ď7^wϟb�~OW��)���2�F�j���[#>}ܫ���Le_A�� A9H>2ñ��Έ�p�����.�������H�	�	�I��2y��x��}-�.��]��r+u�MnB��d>v�#��?JuȪ=�1;�f����&�Lv�k
eNo��{���_i	;>1�8@A��ek,�G�jB�ȅ~Dc��-���;��	Y��Q��F�t����~9�}�_Ε|:����֋��H�x7�f�*/G�a�����a�bC$H�Fm)�R2�G����:��~���C{�w�z��1Ò�8Ŗ;a,6�Z�ҹ���fҔ�W`��u�\+�V̳b#�WB˴Q6�`+)k�Tq��c	GcU��k����t(��X�$ԚcG�v�e���H���	�f�h$s��rOZy1寘6u����F#FK��kHL@�kbɣ6�k�@����l"
"{�~.|M~b�m16s�i�=�_Q�њ�y.�������1�t�tn4W�cQ2;X�gB)uq���ٕM���P~a����1��"�]���A7i��]��N߰����C�W��$��&A����� �h��IoP�����}׸hLi�4����gg=Lv־�%�S�8b0�3��K6��	40���'(6!�)��s���{�'Q�0�z�p�~(qj��˻x�9w�<�4B ֻ4���v5i��9�}Tufo(" k!��I�Ve��V߰��r�q�B������&W�_�Q��9���O��1!2d]4���y=�lL�G��\�ɮ2�ݞ���}�H��A��)
b�T����Y��!��@�6�S)1���uÕ��efm�
�*��8'ƀp��Z!;��
�`�7}��Ǟ��}�%��ky�t�AR7�܍�ʮ�.�Ɠ,pA{�$:
��"39��v���e��k�� �,��X��t]���!'Eʡp襞�����TC�,��e�!�@���|�b�̤bFD-%3
)'��ρޮ i��)�N"v�����?A��1��x��F�:����n����Ē���H@��RiaI���|N���ldLnξ�%���ϩ;�;7I�&�kfA'o��&����cgb�
��W�,C! X�ti���N��iL��d F�z�E�������jN;;x�R��4v�����	b.��l�� �f�j�z��f6�A�����9�	��pE���1�x��h�xmP��ާK��nle�SG�4���]Hi�Dr��a�~�{�/�Z|�Gs��L������%=���%=����&;g_y��Ʊy������@�Ajdk�� ��MFƒ`���w_����V�>m#������u�����0�ߜ;!̱AyÃ,@5���*�-��[��I9wy�T'ҙ��#T�)U��\w�֮����wPڵ ���cc�\bTl��uv꼲�q �Ct�0��Z��L�|Nn��*K��9�%f�.��E���3H;Ă��D=iI��0�J)�}5��Lm�A����i�Pr#sD A�p�_$�P3)�{ۛV���OQ�I�[*��L��d�_���1�:����j�GљW�W�M�L}��S$��� f!�Nc�4DV�����u݃��߻�o=��;HtYp h� W�9s4��ld�%ѫ��!�{NHo�]��5Y����J����,�Rh1�o_>|���C�\vRcLa��F�'Zyλ�~���.s�"_�W7�\�C��E�Ñ���s�Ø�n��^�	�th���U{ �x8�K&ȯ_�_�c�u��\z@�t��"����3�J���>fy�X��6�΂I;�<2�E'iL �"��p��-�d�����m��T���<K��`��3��v����Mzf��0z�*ԐF&�:�'b	�N#6���c���[��b%�.����8;�C�����}c"��7b�fsS��y*�;��0��,�ڸS7�@j�l�3 �9"�خ�Q���
R87�C'��R%�#4���?���o��3�[�������F��q������ � ��2n��=�w����Ird��b���' ��>�N�h#���c���\��-+Cm`�1�v� \�Y�!�q��{�=ϒ�}N���O�fЂ=h5�������js���K<b��"#�W�4��ld}���N���l�e��w#���y�m�p޶�:R�Ʋ�QysN������#�}h���#=+�*33/y8:��mC�l��ۇUKD1�=-�N^t��O\?L{c_y%�Bc�P8��R�,)����\Y�F���Y����5���X�E��~~��9��vAG8&D;i���v�|�X�:����/&�K]9pQx{BXѫNA��ݮ��C2�Y�@8{����1ݘ����.��A���T��& ݸ�}�~�\O��.VB�����4�m���S�<�L6^��U� �I�3���Y��V��c������f�q60������]�s��"	B �����K����k囑�A�қM4�Y��X���(��*(����\%�d\��
cF��F��6����l��"��]��W�VZK� iIH���&�Ylv���\�n��k����"�Yj��vE�[ �D˫ٔ��9SsK�:k���,#�A�Msi�M��,q4�KV��i�]�P��ũ��P���5��2��M��F�������?X})[�Yfq�t����Za��FT��B��X��Ϟϯݤ����e�|;���`�DR�DRd6����~��}�4m)CFn��x��n7�Dbvv@��5H;óA�0�Z(^�6B��P�Vgur|��x˻�d��!�\9>]0��Z!�b�v}c �&b��eM*�9`F2���3��=>λ[}x�~�>��_�E����G��%yy�O"p�$����U��B#Б��gj,������;c_y��������b|�R�����'؞Y
,�)���T�ede<����H�Ă�z�8���{��G=.�s8 �	�\�{c�)�wgb�:�ݍ]��$�S8�%		���#��Pݭ.י��MS�����%�$� ����[)9�($�gWi�2�'��U���߱��C<G���G�����"�ñ����m�F`v��b�޿%N�Q9�Qq'�`��˵-���o���P��@��O���inᗺw;5�����|��jڕ6UX�E��]!#�|��H�KZO����|'y�'_ba��7ݯLvƾ�K�'ҝ�,��W�5�/�t�̓�+\�������AyYE۰�5�7ފ>�/�ϗ7��#^�{���x�L�19�2o�`�.	�NB�̕��!3P�Z���%~���~s���B�p
���=@��r]�}��NyL�dý�iǩ��s,r;�+rMhV�l嶻۶�^7���@z1`uT�ZB�T��{\9>ºxϮ]לz����LR7�2�Z[��K��XƷQ�Y��\����ׇx
"xx�ìDj�K�F	 �T�=����{#�k�A�p���#��Kp�Y�Y�0�Y�%���q�(f;��ϮpǞ������O��[�z���y����A,{cYb�ʡ���P!S���{c�NiDn��U (��L��b�t�^�]�.��z��VeAY�:8��r����{DL�6= ��|U=���V���]�Z
n��f>�6\.�������=���em*A n����K���zy�]5����u�xtv�urr�.�R�C�����:­�k�{�ۺ��h�kq���6���.�o'�{�.�6A��_�.kʗ� c��Wh�3�����fX %��b�����\!'�eGY}��ƷRU�F{8m�7+�����*�v� ��T�UЩ�H#tn��	�ɤ^�a�Vs٤�z�V�F���̙w7i��6�ͺNO�5��s��h���
Y��[��7�3
������9�.Zg�f�6c��PX�.��EJ�=�YHm�����G��h%�̺�k''���H�-��<Ӌ�5�jUƷ1QGd7+b����c:�ɹ9�ne�5	2ž�ہ�[g]�����*�<���mVr;reˡ�:q�H���\"�&������t��+�H�v9fzwXP����al×�鹶+�v�g�	76M�*$���^�d8w2�2S�x����^���� w�[�؄�;n�O��9Hl�4�ܬ�_]}�ځة�����u�tg5�j[��_;�
��+�?��a�臋$���I|X��Ν�޶�&��fPye^��^��7�F��.��s	i	7e0�$W��҅f}�W>��|*��9��RՋ�����Z���2V
ͻ�^����a]�}Q��r����D-ڲ���t<s'�.�����z����z�˂�lЙ�anZ�2֖se#�J^�j�r���L���51kko7�Z�f����x{���={�k̆لL��)=��'�ۆ���$��4l�Z�F�s�g%�}���gg�ٹ��ٹ��>��(�{r���r�\E��l��z%!}�\���&	K�Ŗך�Z���̲��e�}��䳳����������O!�ȧ���Vփl�[m=K�ѥ�dLKێ"��Xj���k[V�,�ϣ77;,��{775;77>'��R/[��ƶ)	��i��g��r���6e�Z�4��%qlѫ�Ĺ���ϦM��x�~�_ߏ�����?�[���QwZhpEwv�cɺf���q�l�ˠg���>�57;,��}775;77>'���ik<qX�Kcs'�9������ӄL>��t�nx�j�޶�}	n<Kb6�R/�)ƅ:0;����F����O"�'=OP� �-�����{JM�y�]�%��B��X[�tn���>	}�(�������;�
Ke�����*��V�*Z�S7�LB��Z��S6*��E��ew�*,6��sF����ZD�#hjw.E��S����lv������pD�0��n"��NL�SR��w�@�v�O_����vNER���	��{~Ҋ��x�!�F�tm�.�񳠃s�΅l;4B��uj�?�	*Lo3�<�X��V�����^��Q{��{�]��u�\$��3
0�T�}+$߉Ӊ�O�Ԁ��3�u�We��\UFf��Bڍ���ܸ���'�7���,�m�^}Ox��� �{����Ɔ�lE��N�s�z{��JX���aOd�I�S<�A�׷&����G!�I�Y|�Ȫ����� �6D���w	��{|�0��$ C�Ѕ=ܽz�Zim`��L��b�QY��Rg�{�';���˼h���u�&;v�&PM��C�ܗ� ����7��}1޿7����FRLC�&B3����==��]��s��x#����l�O�td,�����ϒ��wF|����W��ovj����{�fq��X7p�3�h�o���t��Mw��zr�=�Z�2'	O5_7��!�	�D�i�C7;���/P����=40A7H8 �ۇ)����U���u�\�_�}ԭ��;Ig9aT���\��=�� 0m���H�W�U`ݫbҲR��[�,^B�0b�W[�ϗ�eB�Z�/1�#���:�s��lP*Ӵn_[�`�W��������~ı�!D��ct�>l�F;Ă��M����Τk�C��e;��d��~Y�Gf��I7ԃ>&Lj�l���^Ə/5� �@��Zi��iTB:�]���j�D�m��m`����c(qH@����w�)�#(��Le�I�Ա�&uf����-2b�@U {n�E��{�/x��m����!����8B �8v"��DP��qD]���eȦZ��>��C��?f��$��}I� �L��S�j��n��em�	�&�jݬ��p&�����p��Pى�y;���G���;��a�=�J?��D���D�+
Fi)&2C�^��r֮6������	fcv�`���MQ�^T�kf��Ћ4c.mpdc]ee%5.j��W5��wQ;R..�X��!�;	^�k�K� T���"�k6��9�0MY��i�F" �u��m���C�-��N6�1����	,B���4qu���Q����%�Z�m]�k�/s�3�,3���\�p�����Y����պ��S�\Ыe�5��Wl�6#t$7n4��={8���`Jzn~ �r�T���p�h���8����j�91%O%?I�r=�j�2�Y�@%�Z� ���1��Dy3�[�� U4��g%c[!�t� &����"�?��R�5��t��A;h9`Fc�.h�e�"�]R4X�}.䒄�9�!)S�2ƒg�(�����]C&=={:���zY��Aҗ�%��PAmL�)�,�%���@�@�mo�Pq,�R,`��A���d�{��q�|�3��H@Ջt���'�z�h�ԁ%Pe����p�e��Q�M��m���c��ۛ�����:\nm9$�{d,� ݸ���Ұv�[ͩa(��F�:%+`����M�qD�f�X�ks�}�BO����~q��eC�r*�ڋ'̮�~�����&>���:��M����pSJqNH.	pE ���C��(�	�zE�/���`����7;��o7�g�;)�}NR �(��?���F�;>�2����o{�Sn3���	-��IXR 	��+)L"CP>4B �j�=����]ƭ��8&H�!����ʛQ��q��c��v�%�֛�AK.�2
Sc����1Kq�՝����|���r�rc��D�Unc�F�#��YC#��NPP7Ka>L1�Y��b�p�8�^݌&A���o�n��Ip �ZpD`~�
9�Z�u�1��F�[�
���C��! �t�͑aHW���F�����L��Z���2�s�� �a�+ci�؋L�V�+��we�����C��Iv ]���K�V1cͮK�V3dZ�ͮ�>���o�K6/�e��+��(�E�{@U(v\��Zq]�܇|���r������E��C�ED�ZHCO�Ü!z�a���D�#�Ev���X1�
wv4�?enC�o�i�޶w~-�NA��G��������#H׮����$��Tӌ[��#ZB���u�tM.鿄ߠ�JCh����>�·���h�n���:�p*^�9�yy���A&�8$P=_'� ߍԺ�5��� U��r�n�FFD��2R0�d�Pd��0D ���>����k9��4@BqĆ"�v���K*��蝬⢥���&�$�V�X�Sۙ	�+���Ꮊ��� �w���:�(��5���y���J�����mT�yze���ِ R����u����xhv���~��ӱ�Is�� �ӻ'b�beʭA��<.���uq���q R#6b�a�s��T4��m�Y���g7ﯿO�Z&��Y���ɏ����������뵜%�\U�J��R��Z�G�.ņۍhei�a �:�f(�B�-Y��h��#�Yo��Mҍ�e�Ou˹��G��c�����&VEpqOx��Xؗ�0�p��L��J>!y��,�;ܙ:��:�s���b*Uuþ{G��l�;� �b��dƩ8"��9Qv󰙷P�i]�R7ٕ����s���D"1�ՂH[��{�=�0�D>m��i�S�p�����X����s��ۍ��j9��t��8,Ȟ���3w ����]Ϸ��i��T?���"aB��	-%�!1��nxS���Ϭ����y���I� f����Fy��;��U{pB|����G�l��E��(��1�gZ����ۭ(>w�����1k���m�p�/."��eu�;����	Аt�;P��@FZ�r��Mf8v4�?z�a?{�ulpˍ1����g�}��)���r�I1q��v��x6�4g��׍��Ƙ��p!�w.�]v��ʦ1��Li�
1Â"ᦽ���5]�ͳ�%��S�x0�z3V ���!U4S���M���������E��]��2����&��$�81�5�OYH�sHv�!�	hS���h�m_��{�ulq��Am4m�i~��w���q�ZB��8�A�TM�����H�n�=^�g��a�v��e4B6�
�i��}b0���[�D���(���f������\�;�ޠ�����g�����?b��Z��,)(*���khآ�t�\1��l;��{�sfh���)## ��Ai(R��q�|���O�-��jꆼ�l6)]0��q��6͡6�F]u��,ZR̖<�9�&ss[4ʣS����]S[Cm\��`Z�,�8X�$�+W5tcX�.��h�E�"G�V�fjf��k���zc1�L��fց���rb0MYk�t�9�҅s����3*�k�5!���utڴM:,%�RZcCsJ��#2X�"M���h����O��[��U�nхԱ��f���4�[�J�طv
?@E���vsv���q��!>W~�;:�#�Nj�����#eñ�(�)c<�\F� �1m2�2�Z��wb"#�H�v��8������V��y����t�F�UO��e��Q��R�c�w��� �6J�L��AȼAȲ�"���v#r�^N���a����w���N2��0Ns�L���[R��ά���z)�Pg9a��@-R�{hd����y� X��G�+�1��\J�_R���1�R����-_���� `<S�H��T����x��Z=��A���ձ�Ip ���X�����ɦ�����v�^��Π�N�)�乴mJK�����Թ��e���(�|��Q̽�G�O������Zd"!��G{2���a��g1�q�f��y=��"�7nt��L�I%�ԝcL�:rǩ�O�ֵ�b���[�&t��Yj�&�h�ab
��JM.Xs%;�88����;���6���P'ԼV]b�^�<ǽYkT�>]z��:������1	e�f��������d����pG��ZBoX�D,��=��;�~p��Ap��S,h8"�Hb(�;U�jC��vz��f�n�l�u���Kkw�Sv�Oj(L�^��!l/}҃� ��Þ!S��e�o�%��s���L���S�Nl<�{�O���i�씁P���.��f���D{$�s�2L�`�r�ve7�U
����J���b�c�`ra~�5)YRVU�7R�m���NC�H�
 �P�-V
hn�`�r�j1LXA������p�x�|;����[�Վ�-E6֔�YsMg[C��_�Ⱙ�`�R�mw�'�ތx���3�Ɣ4�^���M��:h�l���{J�5W��r+���!U�e;;{�3C���U��vuvj�H��S��[%��zN�'r��)[�d�1Ϧ�:�}��1X�:G�(T�����O��w��ƿ>���Q���H���=v�w�ك�kO���f~�@CޖzI�z�z���ƹ�ct���wP�hC��ܖئ�7����~���nny�'k�n�����=f���[&�B�[aUSNJ�e����c�Z,M����麭�I��,z�lB�j����;���c���NŦ��[�2%E��:G�llF����U��z��k��s�爼v|Z�RO���z{�����MlO;=Ja���D���~����a����hi����ey�����ǏY��<�E
��HUU`����;sW���z�X���>I���t�u�*��ꎼ�S5`�[��2�H?YH�W6�֙���b��$kN^:�QT�%ՙUuN��~xt���fA�YSW�;��r٪+�h�R��z�w�k�����n��S�#64�/r�b/��	���ǩDJ���<�
V��. L���l�I\ݵ�wUv��M���l��^��;�T���UR��Ϸ���w�g��u�;'a�Z:@�P�n�-֥g%�yýԀ���9&o���p�Sx�S�_�o��7�0�&G*��HUD���|f�6}Uc��}654�o0�L���v��6c�.��:��g��p�m7��ї�g�acU�އ�2{������f ������5W�������.���X�O���P�,����`C3�룵ӱ�"�ʔ~{����+\�yVKfS�ut;{�m����\ì[�z�ٷ���O��ЭZ�w-�cU���h�M�����ü.*��)�k��`��M� �JtyT2�7���[j�V۰�5t�i�.��@ #5y��IM�������K�W�l�9�Lnt'j��w�}ju<�F	�ܩw1M)�w9�V�ԷDخ�"��S����jEˮ�����(��ٺ��r[K��V��N�;|&7]��:��i�b�g�-|f;'����ՋBFu�C�u^1y]Yhv�u�4��d�Z��C��*���\a���^�2P�VQ��[BQ&��]��_v����7�o��:y�K�1)�]�2
�톖��NnVf�V/a|�{�c����Uݣp�3�UK�6�iN��'/o{	��;��1��z��p{�a����ѩޅ�r�y]K���ǹZ�-��{��Ur�H�{��A�ھ�I�|;,ќ�쫬ɡ(p�@sq�wgc�76�ҫ6�T��.��?�=�C�:�F�g ��㭲GV��u[oL�ۙ�M��B����e�0�f�t+{�����bc� �p�0[���V��̻��:����eѻN4=#�pB.�Dۉw.��x�;ؓ��CEX���Ԯ����D%b����N=/!`�3&���R�h���&;��톯����f#/Tyui
�p��u݇^R3mS�����djkè3j��J͚�i�l!�8�P�7��[]ō�� X ��l5�!�h%&l�*P�U�g���'f�e��O���f�����}��O���idH�OgOA� �xHeh/�f%&����Qq�6ҕ�|���Yg��O'�ٓ����������O'�؏�Q5�i���WQELJ�U-]e����� X^�!e��R�?w���q���~�>>=����j��jQ��fV��j�Ī6�f�%������g�$�oqv�օ�*�ѴK�j����e�����>����9=��g��gR�Z*)bY�����RFްMZ���i����i�4�HЉ��z�3*��r���<u�ێ>�?^��ޜ~ω���J{��K�q��T��а�|}Y� K�����zf�e4 ˽kT�V����U����^=�}z~����8��~���{o\O�#m��')����KBXZ�Q��GV��]|K�Ic���톢��CBPP�Y�l�Cy�4��e���U�%����(X�*
�YQV����,G�Qv����E�j��W�e)m-*"9J�<��-kJVڝ��ݣ�U�����km�PkUR�m�
�Q��V�RҭJ� ��4t��s��1Mh&����0�V�i��O4%��k��ZF�$fl�EaL�F\��	����FS��`R:m
h��8�:j�ca��e�B�flFZ&�NC���y�c6�3t�-� �Ƃ�]y�P�Yk�CK@��`in�8e��[���kR���kb��efv)1t�k�ͭ6���3�lz�
�f�3�r���B���](�Nc0�S4t5f��m�ѦZ����Xۀ��i�Y�S�͇�8�J���jgE�Ԏ���@�] �jjh[�Ė:�1D�:mSC5�4 �2�h�+{�Lh�$�T��iG5�aq�ѡAq6pjݠL���*�Q�4�]�vh�l\�v����3fX�h�[oH�Eض��4#��՛`�WB�ciT��V�lf���&�s��ck�2 ���]q�d�E��/�R���ᴶ��`V�t�0�_���l/:k	�n�m˩0��X��
2��`bk��+2�SjHv�����Ga�Q�ر2[�dMrh�g`J*f�Xj����CL�&p��!�li���`5��mV�ja�[Y�(�g3e�e*6��G �2�ư��1�Y�RCku���` leB�Ψʄ�p�ݛ���9��m	+���m�Rm��`��T"��f��5��p���/E#i)�f0:`��L�cML��eEH�k�eq4�٦E��k[t�w	0���b;Bimt6%c��X�YUe�2vқF$-c������YF�riH���KS!�i�`*-��PSWC]v.abű�,ҡ�vĹ�a�r���a�5��Zk�k�8kM��6�)�֑CE�U�B8�st�.�.f"��װG2��e��gf��Ĥ�XM�����{�|�##�n��!�&���J 	�qf<c0����2]��eV�#�k��Fl�t)a��uf.K�,vN�WE%�·Z-�	RP�u�H��Vn�7�"m1�0�e�3���i*K�I:�q���Jėѳb��#�2C2�FR+��\b�����k/���Ҳ�iQp�hW9m�Y�5iFi
ި�TL(�5��
Vc]�NMi5e��F6�0��8�����Jv
��e��L��Q!֒;^��ͩU�f��b�)��䫜eѪ�Y���cD��j��9#A�C&�Y�k�q��
3KiL�w���}\~��;h�e8Æ���h���B�G6�6O�o���}?hA&a��L=N�R�	�*�;�=�scd��f�.!��� ���n�.׽����(��ϕ1��e�o}ё�9{���L+S�WW�i������|H#�=�]�j�j�L��a���W��	����a~Nνi�T�k�I��KWi��j+�<��v{T@���~��|9�Il���Յ���C5�71�L�.�W*��9V���Coy�j7=�NG����&,@����S��x뮮����i'��D�!^
	(#-҃��cv�D��pm≄W[篟 [,
�&���w��9��
���Ћ}�yγ�{)u��#`Đ�YS��J��M�)7`p�c/؀��w�T�J"�Gs�>�}Ζ�wu�Ռ�G�r)�rk�I�1��V���v޻�?[�OR�M��~H�4��k���Kkʮ=��<�7cd���1g
��r��Z��w��A$�����I�����5JFGMO��7�R�{�@��~���I�A�̐��ޤ�����6�R�ƄX���i��X�gjcoӭ^H	򖢃�8�B�,<+���"�S;������Ҹ] '���,�)x�d�ߧg�����|�����~M��4�:�\�	�C���l]��J�R�����샘�� ߟ��nC��Z�ˏfz�����nox�Z�z������u&�&��6⠒m]�=Ի����#�gP�bo|9�s�֘�5Fz�Fz�z�B��i5BHk��[ކv�������]�J������U�f��;o��p�����V��l��u�]Ru\|�f�=O�ܔpR{���/sg��u�@�_���BX�Hb�A�5�7P��:�'��RdŮ*Z!Q�	9�՝�'��*�N*�YUs��s߻m�o|g���g���=L/"�I�R�������MwTn�}R9�x�;��	���Ws[&�[ $yݮ���C�X��E��`ű8x90�(p��P�h���b9ƹ��i�����*ޅ G�^������v~������N��s[�+���i�^�1oT��O�1k�k��x�\���㱽M����F���n� &�*�s���K*i�w�I6���
�&��/�;���#�r����w0�$}oT� E��hNazr|ۯ���ɕ?�������d��Ӗ�{��]#�����c-4�[7�P8�Wa!.���۾�+������,-ϧ��~��৵�+������Sf�)������=�zq�����*EC&�M��n�j7�[���p#��>�d{۪�s�)�v�*��!6�T���/�/DU��B�X�l3�`âM�e��	��@�;bꙘv�eMkT�u�/Nv$E��Ӻ�|O-�UI�U!�^40N�p~sl��Y֌�~�7�eɐ��7�9�D�AЇ�֯�r�����>�O��>Nެ{�>�]��'��;��Y�}����B)P}��&�#F����,EV���$��f��z�#}�o{�c�Ba>UH5R�l˘�{�N��1�i��ӏVꡣ*��s�A%w�ClG�0{@[�
�9h�Q7sdڪݩ���A����k���0����5��j[J��U\i����� ��/p�q�Sܔ�m�+��>a��НFF>��7.�=���W�z/3�]LXC�̷7ٛhBQ ��b�7�d�L.�
X����ju&5��k��5�(�a�b�5�(h�\�M*9��	]t��23)u�KqRF�-w+��m9Fݰ)V��B�f6���e�@��1&�W:�@���A�,e[�,�&�fLB��.�F4�Jr�����S�io-���p����,�LY�����P�G-��J7-���m6
�˒���WM�#��Kv�S���[������?4B��
��԰�T�WCg.R;�9��M���d���_���X����nhg�C�Q}o����������6d�ĝ��BqU!`a ǉv��;�K�P2^�XYg
�e!��T/MVp�t�����:jt�}tqy�Ad3�3ݠ���\C�z�줽WQ�:an���>�U��*�©U&��~�=鈎����琪�}ol�^_�C�t��^�a���k5Fe�6[y�<���$�lPb-��Ux]c��~Eb�GR��Y�4�������T+�si��x{\�_���?PÂm��.�j�h2稈gu�j� K�y�|�o��QKd��C؅R �Q{����]���K�o ��ݤ0�r|(
�g�$�4��{�\w{���T�B��*����`M""���B�Z�iH��x�"�Jx>X*�E��_?qOf��k	�g��f�fA���"a7�t=�K����y|�g��t�*�q��֮;�!d�bɋK�<@3�!�bMv�����V���&0V��ޤ�Q����B�@U;=R��+a\�)dd�HMg��^�zc��r6����n�^��g�}��Ϸ+�@�ʌv���A���]�Z{�e�z�gy�.r��3D&�T�U`S�����n]��������g:��lu�Ʒ�.��5HM4T������R}0�P���[Zn��M��Fb��r7d^��T�kk�f� -�N!5�ֻ����y^Ol��\K@���ҫ������܍��.T��F���Ӭ�$���
�Ɉ��`���v�k���]t�~s;�l��@O�@����e{��^��^P�턅���J"�֌����Ӹ���'n�Q����C�6ub�W$33�6��vs�^U�� �C�����c8Ć��I�dT>t��rM����aP�@�P܃Yܩ��/����Go�u�r�$N�-#16Z�B���X����zc���h|������gjO��P����J<;��5����:��av!BX�c]�Ek5u
 �D�84�C��E"Q���jH"�I��k����ʾ)7�!��dw{6|�ҟ!UyBH�|�3��fyV��ܺ�3Ǒ/��zF�
�2���~*�{��@
%��������Th�/�J�ӥ�z(�"�Ty�*���W�j
6oKi%���u�,ԽD3���!|%+.��˹i:,c8��B�����,t� ݈P��7�Q9s3'1��6ͦ�;��\-B7?���:�����Y u�8�� ���
N���D}�72��5^���H��S��e���ѹ'��B�
��E�Ʀ�"�'���P^yg&�sʪ�z��O�s2o��^�5��?l�w��1m���T"8��s����.y7b�e����2����ܾ��=v���8���I.�i�bBbCl�4�����h�RJܲT�X|�d�V=���X�2c���3��Hb@�t[|H9���D^DEf%>���>Y�����:�x;�3�a	�s>���N��#�ZI8^Q�qc���v�2�-���bЫnP��ϟ�Qj��v<�y�g�M!Uw~��؎���=;z�yV��&.|�	eI�.������U�8��q���;�*W�rG� �&��.��nfMrE�����A���nҪƖq� E�5zgf���ݞ��d�w�|{��/��Qu��~UHCT� ���/Uuz�䅱4}#կR�T!�^���t-|�>�"��y#9�Q3##�(����c�+����A{�^��ml�^fMt2g<��4�U$ƪ�{ݓ�W��e���r��߹d`X:�~���-3�*�y��깛�Ck퓏����8��<k�'�I���(@���/�B=��U!�m�5c5���=�¸�Ќ�5�\u�K�ty�Dx�h�1(���h�f��2�JJ�e�
[��w"��`�U@�Fs{D�+C��΅(���n����cM����Xl$5봮��h���`me�;�V\�5��X���L+��b�;�덜X�d�+*�����-��6n���U��߿Y�ue�H��ZCZ�U��r�]^Y�4�Zm]M���9w0�-���/�ri���N�}����apT�*>%<�����@�]`�����Js_�½ʞ���l�>�l�g�-wu�^���J�p$�;頻Vd��M@U���i���9� �z�2���M�=�M�����8��>;�K��ײ�c왗�n�-ib��G�C�FKn����g���Vǻ�t�;#&%���b�3��g�5�d����ZEڶ�B\+�����*�E\ۂV1t�\(�(��t�bW@rڸ��C������A��A��z56R��	'3Lt�K��2������cܩ��崷�=(SYZ�w`kAN��6z��� ��[P\G]Z6�ڳa��Ԯ�0���ײ=�ͣ��+��ͫ����s�:�>w��i�k��bG�@P�&�,��2#5�fg�?I���f���q����H2�{�&#1ߚ���/lgi�t����_�v'^u�`��c|��U&�AH�����?��M�:�P��NS��u�Uő�P�kL?,鎻�*�y5RH���65l�5�z=m�5LU���Ջ���&�UETm�|�͢�X�6F9(�ɚ��v]����ұ��p+�W'�7�w�,�Hz��a��h�v۶���2�����O<���>�8�fe�M�$��vv��'�P(T
�i�{���(��>M�'{ޜ��t�eO ����z�^���Fn/3�@=�URUU>��o��V�+���������88:}����E�������m��9:���`�]J3�
G�M�ÃMg��:�]�.�0����HiZR�V�-��5�j�����T���Ū�V�+op��=Ce蔀���FyԽ�K�﬋�����<%_0K�����xkٻ
j��2pLt{+s���_]�
���Y4#w�%$�N���Ee���+����bɛue�k^��am�9�(�a��E.�6�>�U��a���.O&o�hZ���p*�X��&56e����'�6���Pb�+i�yI *�L�ZU);�U�ٜ��\w���/�(+������˼ZoF��K��B���w�YU��m���h�-H��TX]#b�Bh>6�ee���Yc���V���[n�va��G.ۼ��'�b1[uznv�6e U��Z�ۼ��M�'�����v�Y�fس��[C&vnV�;����+�2rڕ:K�V�3�ty��*M@z�a�Pd[D	s2���4�m�뫻�Wr�(di��Vr�0^^���[���c�v|snF��{E�������9ٗ���/L�.[�!��f��9v�(��N-a;���fK�Q{���pq�����_=P0Y��9e�xa��
ѳ��9J�5��OJ2)!�Iw狁��M!8��wN��4��h�����(��}�1�^z��]��{��^yx��LԹ�b�`�0���.��X!u����pvL�ǩl�^�r�ރ����(i߷9Hm�h��{L�����q��Z�Ii(�D�Z�f8�:s�a�ۦ��3,8��v�㼻v�dA�aI1:���D%x�M��4��t�
� �C����עՄ��ȷ�\��F�  *E�Uu1�Ϋ��bl�b�,��UPUV*�[R���kV�#l�pq(����*���.2�=�,�Y��������������O=}�KJ�b+hT�g�{ h�-���)�*���+U����:��MK=�jrvy2}5552r}>'��A��)�jX�-(�o�]�R���X̲���Q���3���g����ϧ�SSSSS���>��c=+�����V*�=E���7E��e�"*��m+����%����O������'��}==��W���ƪ�l��܅J,b"����Ee�뉌Ih�&"���%�},�����jji�����~�?=ښ��`��]t_n��e��f
.4b��k���UX��11�����e����O&�����'��}==��E=Jj�#-[-[T�lEQ�#YQD�UD�.YQ[k�殙\�\�*ؑ�G-�*�Z*�%-L�C.8�з̦"���"v�DDuh��j��TST���FشalZ,��Yֱr�eTP�5Z���nC#�_��DTTES�QE�h�(�Ut�1���~*���KZF��+sΔ�g�T�?� �/RI��Rj�m7���!������{��\��lFJNc٧�oh�T����;Z����؎�lo���;}W�S����M4����_d{WX"e��C�T�$a<QN�hs6�\[yfk��f��]M�T������l�� �Ǹ�*+�X�K8�MT�dzy����Q/+�ۛO7�o�G�#���Ho*�T��GJ�G��/�5zװ�ȼ��{�|�>��v�ϙ�{�ȿ��ox����^�L)���H=g����C�=�bn��(�ʊ�m^eOc;�)��h���1�4���\X�U��UT`��*w�9L������l�Q>{���i{�`�Ɉ��M�����g1|8m�Ev�p�W}�Y�����<S�
=W��+�,8<�Y���*v��,;�7�6$P�@�#��~�R�+���3���Y���ʵw���f�w}���:��}�����*�!����ݛo���;�"���8t�M�8Ή���9&lڴ��l.��i���p�^�l̡��z�.����&x�=HY�`��ߌ�mY7u�xR�P_y��	����{t�i����u{۟)����Me���Շ�5���9�I0Kߐ��v�Gk�R{��d�n�|N,�e.���	���Ŧ�\K����/ó.k0�4����.��z�&8�\'�U��x��-��-���OV�*C&g!��7ұ�\��h�wnr�y]ӈ�*�>�y���7"��ъoX7y�9��&�U�|l�c��u[o�r�6&U��!x�q���f{+w�D��<X1!�X�d|���
[�1q�ff�Цj��Ƶ�ٮ�F��,�u�Ǧ��,M�J�I�j&��K�h��j�t�-�"*�@�3J�i{+Kp��:��4�IEm̭z�� �ںL�(��ٌZ�8�*L��������jR�[��j���:�aL�RM�h��".##e�����=�e�h,�ͯ6�]c�������l�S�m���ͷkG#�5҉�p��ۄкZ�a�M^ ����9ST�iT�.�ٻ���t�y�w��s�Ȫp-��6�[�M�]�1"�׏8�� v�����U�>�ɎK�\ 'f���L��6�$�;� e*��|	%mĽ�8��ñ
e��X���ţ����Y�*qz5EGt�u�oCUK=������K5Ϲ�v��B"��{6�R��A�̜�b���&��0���ϻ��[������ó��DUr��x��/�"P��ҁ; ��T�%�AMY�:*P�1�C)M�F�Z��_#��G,�<��:ZukE�X����_����
WsuY�w����ܫ{��z�$��L@����qׅ��/vM�crR�(�A�	�T;��m[
��
H�J&]f�]��WP�j�p岻nBz��$����9�W.���������;���ٻ��:�f�������6c�l�1��i� �{g[�
b7v-�]��Ϸ������ڮ�z�r8�0�N�N�*
���!ʻ��KK4y�q��Y��	xA�ܮ���ws�C���'tz��-zRm�s	D�f{i��e��e���ln�����Y�Z�"�^[�`o.j�{�Fk3�·&�$����W�@�;E1H^Wi]2�79V�eKS38�����l�3<y��SN��&�pZ��o��U��/�Ǘ�2;ל��N��8�޹arm���ᡢ��$L�(�v�f�ES@ʭП�����sN!��W��Lg�W2��$B$��a���E
�gd��G�&<`ڍ�B��,l�x�ߧ}����p.��V��54p�o��#��n�ѥOO��m��b�U¢jQ\�ňbC q�����:W��}G��9��Rkk�	�R�{��>1�:���]WɇrH-����^�Gs�vPvL�^*]TBU�@RI�S�T\�#�Y��u��dg�|b�sN!w��-�+D��*�Pk�����M12�&�i]�eb�����1r5,�O�7�~�Z����&��Ou���Q��W��u�Z󛘑5�#��*�;&��X�ՏoM�~Y�f�ŷw��V-�]�G��c#�vB��!��zu
{�ޱ<I'\�v�i-��y��.����	tz��aޗpƶ��^��T���W_t��Y���2�3���}�o���1���r^ @�<W�Q������v»fB^�x�1hԉ�'�;�Ӟ�8*��BXs���c�[�x,�;�A�G���*OH� �r����LIm"�k5w�J�[� .އ0�>M4�e�Kau�	k�^��.r�on���^K�8p;a [UT
�|]w13ځ0�H�H�8D��u��e��m�Ӕ�H�!҂By�H��� �6����L5;P��S�{&����p[�h�J��
�2P������Zu��y=�|	1�fs��=��n+�K;c8��ǒ�^�ò�	oy{�QjieJ*�=�;���5�s�����9߇��2�eSs[�gy��1&�_���T�y����^�	OG��@MIϳz:�sn��B�^f���|�מ�;ˣz��{I��W��������>4q�����X�Z�ހ�����uE
�qR�Ь[YJ��	\��y73�������h���z`�`����y���[��`~'�OiI`1B�3������㴥�-�6�l]kk���np�X(-�[4
1tk32SY�a�̭�&��.�!-]ECcb$��m]�ع�\���h3LJ5�p:�zʚݕk
�L�Tīu��I����h9Z	��MWn˙e�B�3͙�֚�j\m��n��ٖр��uCKsm��FɈV��J���ƻǘ�����{�g������l"��3��K�� ���f��^ya��t�2*�!DC���r�1����,���[&f;J��ֻ�=�/�����NE�n�O�B�p��&V53�qT�N<n�i�l��5��d��ɯw����p�ް&uD`��Ih�\���0٤��>�\߶�짎�ޜ�o=���pǱ7�Q��($���6�@mgM�-1� U�m��uv�Lv�&/ބ��p�x>�=L� ��Bڐ�4��"�$|Z��q�g���r�m�\�ٚ�xR{=-�)�C�A�	�4z����ˢx�	�[X��	�A���Rr��VDat�� �gW�J�rĨx$�3g����؉}��}��v����\����XiP���&5J��N�6]0�mO~>8��Gߩ,�S�λY�]A��)��sf7f���l��*[�v����G���>���y��M,����^ʚ�	�F9��%K"��Qo>���uv�<�����8�4JƇ�?}��fO��yW�p��Mџ(��^��3[�O|��לL�Ts]�2{���Ϩ��B����nrSĖ2��cڽ��v�����>!�u������,d�p�Z�L���D�k-�]k{׹�=�����458�MUy���U��)�����ߧ�O�Ѯ��!�@Ѫ�j�9E�����M��Е�kH���������1�����r6�{�SkGR�{=���+�o��
�s/ݻx��JC��L���#��w77��g�i�	�{Z�6��4���c/}���3ߦ��d��L���e���T���[��:m)Y�n�O��}î���ש�y�0��VA�5fq�q��$��bj���^^�}T�;�X���eϵ��HL�.�=r
Zj��.Nb�^l����m���Xɚ����"F��F�D��l�P�Ad�!ڪ����;�<Ty��k�n��G;un[S/6�a����:=�{v��D��m������Ѐ5v�l(X��\F�	.a�CPWif��;�e���&�BoS;N���}�_�_��2���N���g�O���Jx�j�.�����w;�=/Yܖ���o3WDu+��={̗7�Rj�r�%���0��O��̏,]������9ܴ� 'm�A�}}��t0�yO!7���m��s2{S�c��?����N�?⮲~z�B�-Η��ؑ��WD����B�f�г��`ò�Ǖ�]k�����'�|������?H"CkZ�:�MJeK*گ���5�Ы7�׳�#��*���1���Tv�p���c?�O��ȏ�
L'|��`����@�Э�pu���ery�~�߿*	oi�� d�@�>@Ku3�H=P���o���n��鋋YZ���/P��|�=	)�A�m(�jT�^���g��n��u[�U�d���	֪~��T{�4H:����4�^k���R�;!V���g�#��S �IQ���f��zv�分��'����|���=��y}6���L�Q��cwm:�5�	{8m���y�1Fgj�1�{2�+����Rij0�`���[V>�vU�o�,;��vm�ڜ��n�x	(Nk��V���z�J���v<6�����wvB��G��:�V��R��2��6k_n[1���r�d�2�0q��2��w{w�w;l��!�o�kI�4��`�Gθ{o�e�n��f����ĝE�K��ھ�S�4���:�Z��Y��_S��Y�m]*�
��;�"���6�3���x]�@6�d���
�>���˜���7���2��J)�Uy�gc���o-v���6��yYte�D�V:	C��|�u�!�C�J\�`{Ԋf��Z$a��xT�.��Ee��9F����n���oui$a���Z���1h�VhűB-�|J]\�z�� K�˫5�6�u(�/r�Z{W�ʾ��h��U}(K�g*TB�N�����T��s3�<�r�Yۙ�h7O��7]�:�w��P����3���
�ؐ������	S�Ux�h	�X鴅fl;�s�H��9�L�}p59m�E��Q=���2��|��j���P��j���"�z�o��}����U�y[��oZّ�ILb�Y�u��'r�rO�]ۍ=��o1�(�Z������w��P��k*kV3#�Xq�idV&�r�0�ɡT�qT���k�}�٘+��G)��jqV���m٭Mf��Z�*���YaT��_��c����f�Y7A�E��R	U�L6㴢5m�I5��G�l:R�Zֻh"e�5�D��A��lDA!im�3�R�?�=�?��������~?��tТ�8�1�%ceE"�D��)}l���b"�aF+�t�NK,�s����������v|O�=�}U��|�USpe��DD]�[Tm�R������1UT���:Ϗ�?_�oooon����ֈ*'��W�UYR�YU1�G�������V�N%����.8�o����~:������~?G���S1Q*��C�څ�,��-���J��X�b*)����^8�Y����ooooo���~��{�V�[B�e��ʈ�MX����T�*&������~�g�Y�����{{{{{u����um�B[�UY2�֊�X.Z(�� �M �ұ�*ow������j��J�ʹaX[\��z�8q���/���*��\��-�,ilU�(���Mk#��"DX�PEQ�]��J��\J
J�5���*�(e�m�wV��b����KKj�~��_P�֛l�0�R[���H����\{/�����f�%�ε.i4S6�j��nĴ��i�=��x�z�[G�-[�C
ڷh��X��	����u2MI}1E�cu�6�
$K])Sl+ͬ�-`���Hmh�4n�F��2!0J6�4.
k	���.p�X��`�e�ȜJ�&�V5Մj�LS,�U5���:��4�^��:j�jJ^��c�K!6���嚕cե�9�������
��x�jd��kZb�n&��Y�ʰ���R��[]l�sf-V�o!7�rki:a��]Vhe�md���,ZX�5SFl���*���h��Ye-S0G�+n�]5��$tĎ�Aв�7@H[�MR�2�K.uTz�.�I��βǨ��lb;WA!9ͬ���k��EWA;k� �SR�h2���5��M��T��μha�]�u�Z ��U%��P�ԫ�1a��0F٦�Y6���rm��@�B��VV^�ti���]k�0ex��	v�vHXn�@̛!��SB0�ƥ�J�ډ\��ԙfѦJYV�Ò�z몹���Y�z��Yku��Xv��B���ٕf��ؚ7Tt��5T�^���m�ma�HX������L�f54"�d��s�nK2�B��hܦ.���]t5���lb���.�3��c��C�Ks,4���v&���=�Q�Z����ԃ<s�1��;]`��׆͢GK��1�j�X�5�s��D,ɉ��0k��f�k]���^+��T��aM��,�1�Uv�b�a2G��՘)K�Ya��s�sY���Ե��7Xf��]�&eZ�\
U2�EF�[���͝ &:����ne�Ү���<��e���Ӭt�.V˥�+�k�B�����9�6&��i�%6�!Eڱv�9ֺ˖ aةvm�w;RCUH���H4��+ج��[e�V2�<7�Pz-%��5-c5Z�Z�D��h���q�6�94�g)s�c���Ec4�s��RYX�\�s�ic[T�j��e�,Q�d֊�B�P�b��B�˴��׈K��v��L��@����)h�#˓J�:R����b)�4K�i#����dsk&Xe��-�78��� m]�ܮ����v�[3�2�&�ح�`E���͕��ݎV܂�3ftZ�)f�p�Z��E�秾���	Lo�%3�&��W`Mb,6�i���`.4�����ʭm�������luP�5��^�p�É��me���	�g��j�/�z ��H
�D��}���u��V��)׽~<��:�H ��X�<̈b����nv�;�w��ܻ���X�L1d�0Y�L/x�m�nߵ�2Gn�����t=>��Q�xk�]���(��϶��&�d�,�)���L���JB�=��|*�wv0y6c�9�����"�����x�l�uC�a�HV-%�����U
]��	�,�thK���~�� 6�w#e	�g�Z����y�n]�u��7�Zfe��y��cThC�cIl�Me.����TL4J���-Ÿ���[�-��wǠ7B)[ƱQ��%��~�ո�ɈjƷ��|��L�z�C�i���dC QfJW3�\fO�c�j79-{=�)��5�U�����P�@W�1�*���^7��g�E�U��ݥ{;��x{v`M�	��rI UKs^Ϝ�1�ח�M�t�{��.�;ߙ�*����~Ў@
��SLñ�-3�-׷�\WH���:רe��G��d8�z�S�ޮ��OW��>I��X�MLt���l�ἈJ����]f�,���Kr�^�-���i%��1�}��n{ү�wc3�V^��l�����# ���o[5z���M�d;}���^�˹�K��0��!��Â��k;y3�B%Je2�Haܨwwy���f՚�V����4��R曼>x�Թ���]�H����UҬ9���N��d�i4e6X�I���C$"X;�<&�^�-y>����.$^܇�Pkb�z�z���g�Uteg��*�kv0Sv��V�u��VK<@$�@�0Z�Ҫ��]w�v)��:�1W{r�s��=	��)K���r;5Tc� ��8~z��GR�� �r���ta��t͆�w;*�u�RSh+7p��wwx�$�m�s����%�>����������]���1�����ωM5T
���I]�v����zm�v�3�jv�����q&�� �-�k@]KQM�\��5�[g՛�u�pޗ���Ψx��rͧ�)���[ξ�]���̏3Am�9E�ʟ{�4�[O���!���}�*�Nة:[�����!��q�� �W��kZ�{6t�=W�yB�5��)�6����6�vv{(vջ!w��ۺQ|j�g�~�{}�{��c��W;��(���V���+��B3M h�1� "�pMT��ҕW[�E�����ߔ��$�l�>d�ҙBN�����r�3�⧍ގ�pM?Xx�����zv[��6� ]�;�����Kͭ�q�U�z�z�w_Tk���u&�� ��/k�%OX�M��p���L ���I��4��z�"��oc)��-ll����&|-TryO<`�^E��9��#�wnT�r\�	�]<��to-]m'�ۛ��5����|����YR4��2�IS�ݕ{�(�
����u�b�Ϝ��-��K�;���t/�r��(�˳�o-3+H�n��ɕ�.���7��ïn����%�x�]\'K�Qk	�t�%�{B�e�M6Q�.�H��ͻe����B�E�ai���e
����tՄ-��QH7�Us�tݴnƉ�Z��{v�뛆[�iSc3Rِ*�,���.W:F0�-s,M�C3(�[�i����6l
v�Ǝr͒���m8ی���TTMi�j�qdlMa�uhL;Fąԡ��V6�6�G��j`�����g�ϡ�Jk0k��#n��W��nҴ�	���N^t��HGZ���m"e��L�۷��Lv��`vS�@�h��ghjt�.�GV���<-��v�zb�#���9ݹS�[M�eD����p���	��M��M2�2 M�ǣ���ɻ���4�ۙ3,����S)���O�_��C@�9�0�x�cI�V�zs�gb�c��q��y���˗�e������Um2&�7`r����9�ۊ����B���˳���IN��]�--+��Kg�yA��C8%��V7�B�5\qRZͦ fX��|��k�]��v�	�+����ȟr��_dl�2<Y���;�GoS&��3�.Uz�st��z����Z����Ҿ��Fc��w'�A�E=ΫW��@[�kj�G]������!�uN���r18;�$3�Pa�[��\��nx�f��v,p�>�
a#��jJu���mٶ �smM үv����R�}�{i�3�#��T���J�Jg�n�4�eH��vC %-���4��썘=�ʟ����Q5F�c��{�l ����b&P��<y���
򼽿�Mt��[�	m�h���EP�w�(l���hEr�d�# �;Ðwu
؉��'�SkR�KX���16A��%�ow���mt�hCR������z��g]�}����Qp�����r�N�) �~b.R�^�F:-����6��6kї�;0{��4�Wjμ�wp�� �|W2�ƫ��}�1�b�:�^�&%/5'���iw���{u���&f�Z�L�;;٩[,��_gݍ�,���PK�Q�$c��zk�gbǛ��U�I*���mU���M��d+�go|gs�om=t�<%���Jay�{'l4�#ކ,���*{n�Q����������\��'fsAjo2��j1�fv}r�����}
Eh���@Q��lY�̑"�t��6�E#I���{�ipw)ᱤ���Y�}M��V］5ճ���׀��G���2��	j���u�'�T�׵M��ý��7i벩��2c�C���8Q	�:�H��ꢐ+i�����a���{�w�������يe��&�;UH\�����yrA}����3	�U^}���O�W-���vJ9�v��tJ����������ց����uw`=̎��Tפ�^[��G'm��\VVL���=<�{��沾��M���C���V��>I�%�#��;��s:��;���fX�@�CZ���C���7�t��=��[�O]�#!
.�.��WF����⎥`�<"���0��"�h��;���S�.��m����b�H�or���C<%��F���V���23��T!� ��d�	.�`T$��Ͼ6��͎����w�udl`���U_��|��߆j�qR��굠늑�j�����I�����Sk���fN�_����@��v��@�@\M���"�QؠP5��!B�\y�nkz�Wm#�,d�j�����&H��-C��͗.�Ze3����H�m�������������Ɉ�M\����3�t��4u;���t��街��h8+[�qɻ*ի��F��!��[>�m��>��`x16 �C�M�҉$p�"��%����?h��3��Ku�`z��]Z昺�M,E�D\R+L�j��
^�]���U̮�D�-mj���n��\%[/�-leXF�ci���ʰB]e��Ͷ!R\.k��.&�kJ��y�Z���b��.l���Ck@�8�96)PК��R�jH����R6Fa�bZ�lɍsΎ��жóf���C,�̥-�l�2мB"�??����H0"�̈́,-&p��ք�1������Q�������YEڦ�p�5;�qT�����غv+��p�� {b�!�v��y�]��$�5������4������M��z���yg2b�c�-T�N�� ��S8t��L�3��/�r���>���z��g�5���%&�|���g�wC�͝mso�w��GlWd�ŭ��՛���Po��*�i��B)ش�}�dzl�,�ʚ͚U�H�4�&a�|��_��|�.�l��hF���`0+-�p��Yna��-�Z���H�&�j�R�����}����`�8�c�=�(��4�yL�E5�ߦ��K�e�cd{aU�)�u�F�vs9FK�SƇו5ڍ:�@\��+kVq=���HV�c�ۉW���T�I:!�4��$3� l!�z�_v����b�SS 5 -�n����d�y��֖���R�X�&��̦���pDu�0�=�w�J����cJ������D��;�)�Ҁ{;c����^d���y�}駬����o��o������u��v����Fe�c �݄���SD���"�]go\d��	k)��%�z��o{�R:�蔋� P�-���l�öн��$���j�랩�F�31t"���॔"3t�'������:�9Hf��um_��vbv]Ú;�/o�@|eQ�m�I�%��LZ}����{ɮ��~��J�ͬ�5cs/%S\-1��Ē�F��E����̠<�>�o�/�F��{x�O2�(v��0X]��ծ,}(.@ zM������[]��+����yX��X8�"�#( 	���hq{��Z�hb�^_t�R����6I��q����k��	�pqA��:����S��ʖ�Y�������\�FB�؇.��+��,�5���YW��!����Y]�m��:Ӽ�a�JZ���ܭ$V1k��<,
q�8E��ɂ���m'5�\;.��Y�r9|���n_+!�&Q��d̲�ڬdl֋�^6r�����E�v����_f=j�=�Ζo	��^�ap>�f>�joI�U�z9!�:(��nWmΨ����jq�y�v�ܚ�.l�7Sb����`�TZ��w\�ّ
[��v�V�c�c\�E�UڈS:�x�θ�LT 	���Q�����+��k���*Ͱ�N��	�Evz鉙%iZtWvQ�GŴk*�������k���2�4y�F�]bю�7�W�����iA�Z�d�`��z�^��:�. �\�
�k��K$��;����㹊��^v���K�gk&tN>AT�)g.�����ٍ��gI��m��q�٦�o��5���ٕqU�֯���a�;� ����r�?>���2��� S�Ivw��tJ�>4l�f+����}>
�l�
���UkoD�oĻ�bI��?�_Y��;� �t�]є����-ꬖs���j���:�&�*�fٷ�9�Ub(��Qr�vg4���R�#;q��׷����_�׌�wIخL�f�QUT��2��#d�ʋ����=����������~?^4�zz��"#�q�+-
}��8��J�-8?\��cP�����ܛ������o���ooooo����ϧ~'��R�
¥E[[Q~n�S��F
� ��C��W��ǜ)��<u�_��oooon���}==d}��V��jT�A2�խX�PPj�b��Z���i���PXǓ�g���8�~������_�׌�t�t����m�)R�[�F1/�T�����f\�Q+H^�^�g���׷�����������t0F#���jX�<��p޵�h�լƅj+��̦�Sm��T�����KKDWM2�Ktݍ��xUQb,W�J��Z�Z�iG(1U�o����)efaP�V"1�b�j*���X#�9JP���e�m**<J�lG7f�2�f
r��Vw=j�	�%����}����|�߻�7��7�-1cdU!2���R�)j�}��3S/��.�U+|ۻ۾�Uو�@2��G�`)�� 2y��C��ݞ��^�#�Y�y���U�X<�y	0�Ja*'x�<��{޿7��D:I)<9g!lKv�U��d�"�!b�S����idC��i$����}�1MH-�}��[�] �w���Ow{<�m�7���S5�Zeu����>+�{�ێ�^�zmWf#��Fӆy�U������9#��Ÿ�g���ce��z�V{��<o�_x�Vm`�BN��v-P�{�ӻ�S��\�ч�&ᄦ�_���ݵђ\�
;T-z�Vd��i	���I��i��f�h�f�.�eat�֫��\��v�[y���{�^�]���xD&�k^�G�
�L��YN��<���<������ֈ�׻ͻ�U���{�4
��Nr�
D�o+�<8��9s��2��d�Y�$i�fS5c�mܞ���}Qn=ie���S�_�nz��}�Y���C��U��Ɵb);�M<�d���@O���y��˼7��2A�r�L��S�\춲�:�t5��g�a��+c�������p�L��!!��T��쮸�ƥ3pL��e7`��\Ŝ
�3������Uf�׮`��R��,�9�A�����CU�|�᣽%�Gk����b�5ң2��T�� ��~P~���'��,*�"��\`�r�Y��7�I�)e�p��%)���ˇcu]��s��%�g�k�8�6��|�M���th�N��n]S J&�F�4��]��if�Pn�B:Z���¶\#ݶ���0��@S.�Hi�)��Y�E�����`VaN���Ci�M�..�[5\����b�,��i).��#q�-�0����m:�^�iI
b��B���ǥ�9�.[a)�,�Mn�R�dƌ�a������f�n!�ǖmd�d�.�Y1�K�t���ʉf�k�C;}����&1F���nqʑR��e�����M�>��R�>��:�_M��\&	��޾���uZ��Dw��X���l�S��$�@�k�k����;V��P�kj�흿o���Vm��^�c�h�6����"� P(l����C8��m����X�z�q��y�]���~���Jlgei��151����k���#���m�U/z'׳�=f;1�iV�	UBIh��UP���^0�^��m��2�3��5Y���,b���yk�;��(M���?2������LV]�I��b��]�*��ǯ]e�
$�]�ޙ$��{��9����rg��b����SXR7n���������s'e����u[/�v��>���:~� ���Z�W[���A��]��!W����$_  , 3�hd������g*z�vbu�)�N�����ˉ}�O�,����8����O�c����f���	l� ����
@�T5>��&a�XeR1����ȁ�v ���xmg?,'��h�}�/��CC�|B�Z�S\�����.�th��=�/��ޜ��1�ėCv���XĦ����	~�y#�*�$��>�x�6�c2BmR�Ŵ̓Y���T��7������{�{���V!�0�u����~�������2��<���?��x���z�J�[jBR�6�kuX=�˶;�o9�a s\ $���s���wC�$�(<�v�/����Ĺy:��S�V��쫰��Ѡ�T�l��zB��������+�y�_�)��~��0�JwO�[���7�� 15H �����VY��Gܘ���D���D�,yL���ם�~S[yX;qky��j���K�i�����-E�}���Z�Jv�es:�#�=x��͍������N�FSE'Ix	��\~T��0�ŗE�XK�e�u��ĺⰋ�z��,�*��<���enG���5�1Պ�wDs��	�-��v�MUS���׈�o�K�&�wf����ʱ��[���;b�4�k�,h���e&|#�2������sx�<�[&ZE��Jd�nllQ�@�E���J�- M 3#��̚�Ո�b�j��}]Fڟ������'`��E�U�j�PR��Wa�NӺ�S���ܻ<����0��X)A��B-4�ۚ�����y��KF�_o��Ml����LX����2��%'�O��{�}���.8�#w[�2��TL�X�"�l޾|��:pI� g!-E�Y��c�6�w$M�$ѻ�n%������8I�1�L����ӕ���M荭�ɪ�X��KOc����i�1�$I0�Ƥl)��U!T���~�����˻���;��mM��@ޗj����]��x�ڕ������w�����O�3���z-��J3��ד��w��>�y�#�ua�Wk�ܾ�'�ub<�KeCIM'���%��<���R�).�R>[�৵ۗ�#����t��A�������_�����K��LR�vLh��k�g�	 �'��޾�z��,��kh�ۓL�tf:�.Ȏ�r�����SKbۊ��ј�� �2��r8�	f�8���k3�̣�X�nR�ۚ�[*V70��]R�n%҄M\�H5c�R�LB\����Y�kZ�H��iV��LQ����7��j�Q�Z�N�-"��m���ٶ	��%!��Nh\�c��J4�j�30윱������a��&����e��t�_�.37a[Dmf����bZ�	50��ߩ��z��m�3�y
��E�|����[��c��<���nx�d�o)�f���	��g�d��M]��;k��{�h���xM�q���ǽ��d��w�$%l������و�ܚ�Ո�[kS���xϲ��@��ЄO?u<�&͗)��7��vr����z�U��ڈ���$�Ե�H�I$.�y ʊ��s#Ngz��eyj�E7Z�i��j�K}˞&�y�$" �%�����:�U�ᙌZ��<@&�N��U@�$5���n�k"�fN�6jxN�'e�su϶9�?D�z�
�>S2�eW{԰���u�t���nn���ge�}u��E�s8���l���{�<�٠W�l�B�jo�;i��U�s��r�s;�of������@P��������M��cr�p��~i�~�Nc���͠m����[����w�����֏�\"�֙�iT.�b�%sd�qbiN�u��uSZ�P�Gg��jxOV)e�Li7,��x�����΅�U��YővL��7Y*r���_�6��{��v�RD�as/RNG!�ē��![c4�1��,�Q�i����0�d�eM��TكZ�\�����KO;���(I�f��{�k���{�'!/',()��d<&��e��g�#��x���ז��E]L�G����2ox�W����*w�xЙ�~e�3�x��S�=a�L̀�v���~����p�b*��g�IBA�!OϬ](M��uoK��=��[.��X��0�2.�CYc�G�\�0���w��ݸ�۩����h��}����ԭ���GP����{�k���z��{��V[>+kk�v��	���=5�>~�o�o)�D��]�޻�8*|}��-����}K�;jGM��ҍ��eðZ8����h�R��~37��I)DE�ON��x��2��U����>�ŏ�aO>�X���ۆ��8��i�A���S|e�b���X�j�^w�}��WR:� cs`����I�X��HO*go<4^�T�"��?��4*?]��	��K����ܵz��

��7ψvNu61�)�5S��a��Ls��^1,���Y����vS�5`�뙦� ��F�,Cn�\��o%�r�㝷Ұs)��]<j�����f3J�)�#�`!������!�����e��bW{�����}��^}]H�\&Cz$~jg�J�����mVmV�_f���Vѩ�f��Q6-YCUf��D���τ��z�	M�|$��Ş^_ދ׾�S�:���1�5�@)�t�r�3�H�<;�|�xߗ����^�y��ر�s{_Є�5(��c��� ��y�����E{`{��R|1J*�E^g+}��\NLY��.�$� �ڈ~�[�1��}�T�nn���ˣ>׈�["߶6�D禚�U��5�v�cUk��%��[���yQ�C@�(�Ic�?�������~����x� ���?���i�W�򢂯?����C�@"08������P��V�A!��H�`R�����f@��`��Hh� L�LJ�$4�0H
M2�0!(����������!(�B G�`��(@� 	 �@��!�8B
�!�@� ��$H
�8��H�! @��J�!�@�  J���
���p�  BT �P!@�U�	P% %U`BUV% �U�X�U�	X�@��	PﾀC�!B!R R!R$$R�aB$B!C�A*! �4�4"�! �!=2��`RB��HB BE9�@�P!
!*!(!��@��@��@�*@�"@�
s�� ��HB�!B%�H��H��HBa	D��<��y��*��R �!0  	 ~��G���?���e�?���h���Kh�o�����t�?����}�?��@_���O�LA����*�����?"@���i�?�?S���AW��~�����Cϡ��ܟ����'���������\��T� �I�I�	�	�
$�I�H d H�D��D"T(P��UZA(�A&"T"D �	�%X� �D%�%B%eBeaY�hA�Dd$F A�bU&P`��I�A�D`!FA�BD`%%RPd!@d%TdRX�Dd A��eHQ���$F	�a$FdiA�Db`	���!A�RRQHA �iA�A�H��f�A�F�`$X�`a!H%F!F�hF�IR�iF	T�`�aRBQ�BA��eHFFF� �d�`�`
XFF�b�� �bA��!T�V@!�d�`�eHFIFB�aI%FIQ�hF�$�aB��Q�Q�d�a�f�%� �`�iF�`�d�fA��f�FX�!	�daZA��A�Dd%  � �P�T)
 �
�PD�D�	*��%EhPD�Di@
Q�
U
"DH�J(Q)����V! &E) �J)Ed��_�p�?�����O�E((@hTT�P�����?����������:�|�<�"
���~��������O�?���?��i��� ���P���^�4�""
��U��?k���" ����!DAW ����8��A|�(P��/����0�>�@jH��?���O�@Dh|J?�o���O��}���	?������ ���O�@DP���;
O�~~����p>'�8�����{���'��� ��dT����ӈ�;�|�������I�W�( ������>v� ����������� ����d�MeD&�|��f�A@��̟\�M|0                                       } p        � 
 
 
        P       P    ��U�*T�B����
D�R�(��
R�QJJ� EP Q)"� URJ$|   F�RUT�����QA��w��j�]) <��Юwr��(����M{� ����ހ�� @�=��{��z��K�E
  �   l }��ي��t�(���%\��gE�h�w�����Ѷ���x�Q�d[o;���R�5�w{m�2�m�  ��  �U! J�@U�IU 
���ynśl�� �� �����y*� v�����JQ�g�@4�`i��=UUYǣl�����S���P ��  ��h(�w P�P��y����Ы0��݀g����M(�C� v�� (P �� ���BJ��@�D�}�̀Qݝ�B�t��S� �F@Ҏ�:n�t��B�plu�T   ��(�� |�l [�
�@҆A��@ݎ�7E��@��!��!��PB� 
�J(Hd�R�%*	"��>})%�b>���:z�'zΕA.�Х3�蔊��*��7��D���U�֔���
�U    =��o���RK0	c����u��Y4B&�";� �EJ� a���w 9O@ Q@���   �В�T��@QB�$�_ ���8��@�v: �uHK�lqP� ;��A�` 㺒T� �@�   �   ������@#��B� ��T �08���!� 1���p m� v �:!����i1��P��T��$�*�@  "~�T���Dd�6J�$�@ h J~�%R�   MBL)RBA�_������_����XI'��/>>br�Ϩ����Ѵ���� �!$�F��BL�$�HHH!	'�@!I?����$�HHx�7����VV+ϝ�=e��qj�J�^[LS�6��x��He�`�y�-+4��(��S37^�Cj|Β�-�H�E�B;�y��FZL�Xv���y�c߈���-^m�*�J�k*�������
��q��˪-L؅*N�<t���؄�4og�Y��'#�2ʧZa�d�*��)Q��%ҹ��e� �MV�5F�Ц%mcʗZ�8_�6�B��u�o±�Yt*��=:/&6�ӳ*��c��T$�u�Y�Z����rZѳ1QQ;�h:��31����ۦ-��xs5��*�Yj����2��,bolDj��y�a�	-�+6<��c��V.G4Qڎ�KW��a1�r͆�5I66�U�Z[�;��Di����VjY���,q��`ۭ����@�M��ڤl�6]���yzv�h�ON���Tũe�0��˼t�^���j��e��F7��4�&ݔ��QZ��{���5�ә�m��z.�[�jnIÍ�3J�.�5��T��#�nEskY����1i�h�7���R�����ئ�Y&�mi:ФSJ�M�A��Kq�))�JwE���aU�F�5��T+���Z�ZuV��5��6��uR"��I:�İb�e�X���Q�SJLr��MG{cl���-U*� u���C�d�?n*�+3/f���nR�Ӣ�8˔YF�ŵt.4�e�����kʹ����vU�y/h�X�=��xooU���Y�N�����ڪ	^L���m�I�j�+U	���kSh�Nk@��L�yN�v^Fȉ��.�^��V$�NǵQ�{�٧f�ǲ��b8���.���9�ּT*���ה����EC�J���lm�l9��b��t�=���5y{M=#9U�qv���N<9`��S#�6��-eK�+.��:�y�pKY�e^�47~,Y�je�+B�m�%��wVUݫ6.�:�먕���ݬ�'T1\��౰���T�,E��3 �Pһ#o1n��(몙k�0������E<�E�q���
ɅL���x��eC.�I,�7���XO11e6u"��h�j�hn�����4���٪G&��E̲��G1c7zE�qͤ\n��ҏc�5gsUP-��mٽV.}/Y����d�p嶱��iCUVa��#e�y�5c6�W�F,�A�tZ�z�Xrձ͂�՚��I�5�+%:������u�vA��%2�^�-kۨ����@�uŋ.q�Tw�m%E-�2wUc�D�ӃP ����*,C��ꕤ�
��V�YG�̧N��A��y���ma�
So��%��I�bzION�Z�X"�ܙ��
����

��A�B�k�W�fY^�y6E@�uԩ��Z��e�:�PnY��w��QDlfC�L����wklH�T���`���t�=�R�W����Ke�
D+�)ī5=��fI���`����̔Nd�u��to]�aGQ�\ɥ�X�1��}�v���mi�z�m���a�W�Zv�̎¹��3�������2��C�z6��O3h��V�X4�JmX�`�N!�Nn�h��I_@kr�p��f,w�����h-��S��iI�/kc�2<j��T��(B�a���N�Jʿ���j�!j�,nm�^nI�Tc8eJ��ܪ���ʁ	qI��.3&�yV1�U�Rr����XsV)��U�M�bۆ�N���6�2�.v��iIY�m���e5���r����YhhVT��wAV��JvVldIt�H�[{����K W���E��n��eXڥ���eV[�Awbnm�[R������bOA�l���Fv�2��oB����^�˛q}sw]a
�ܫtÆ7J��nYŵj�f�E7+�6V��0��1'*)u�j�w-V*M�V�Kհ�K�ڭ��K����جU!M��#c�LSRRdn�0$kj�M3)f<{�:��
i�
�����Y�S*V�M��`��B]L;���1�A9Q�Ɇ�����֐l\1��x��y���BP!��3 ��n��Y��i���3`�jwUb]f,B�9���y��;F�}J�u�ӭG���h-~S����Hؑ����]�F
Z�wv�����df�ti�;�&��U{��ߵ��4�E�;�򶪶�i^"q�hE{Wz�L�B�/\Ʌ�Lr�9{��9l���K��m���Y*�2�)����2�B��Ɏ�8��%&��æ�b�mD�6y%}%�����c�
�T�p�-�r�E�a;`X4m�z)ڶ�ыU���f�K+B�vuj��d���$��{Z�Sڭ�Sbl�걔pV&�x��,�"�v�Z��wF�rf�n�2�-�Z���//41TQl!�f�0*�{�Z�v�Z%���vN;�j�Һ���K�EIX�̋%ͽ^��ed(��Pڥ`�n.���-���2����m��c�͙�;�µm�I�J�Wo^�F-j����.���ߨ�a�p ӌcR3�Kf���S��B�Z���Y�Zy���s0�AZ��M+�70hN����K2��R�u�ݻҋ��^��f���e"��AG�L��%V����te�-S�L��]Pe\�v��$�-�36^���թ\���2-��cV6Cߑ��F��;�k72�jwf�Nk4rR�*x.�+�A7�^y6i��m�����r�9��J ���䪏j��u�vX�uYo��/��fXe��j��C��oS������H�Oǲ�¨T�/NQ���5�X��H����ڋI5eE��z7&㧇߱�lV	3En�%^�Q��VS��U����xU�!B<��YtJ|t96�J�ӄX����K�*�[��lj�,�n�K{K1�q�rCu�&�mG�&�<���&�sJ"�b����-/�C&eX���t��wfJ�vl�:,E0�(1����j�Ø�}�Â<���儨:�,�u�{RT����eD��ԍGiY��4��B�F�uX�K�6lY&�/j�ʢ�`��a4~f,Gr��r�ҫ\²ݠ�-W sNݬ/fh9�b�7X��{tm;��/8WZ�g3n`��o�YEj93lҬ��.�z��ک{%VV��:)*�9�Tpd�f�*�i�ڊ�f���.�u������EG�=�"a��U��;�p�U���8�5��ĦA�*�bi�6,��X���u4��X�X�]��i����T~�k�Ø(쭷�c�b�D�N^��Ɠ�p�&�KZj�R���#q�V3I&��m曘]`�-#x�)@�,�l��:ypb�pQ(�ׄ�a��RW�!^������F䴔[����4�ҧ�*��q�-BkJk&�w��rF.�9�rșm"�4ܻ��yE�ZӬ�r酙�(��꽹�--Wa��q܏Fml�pJy��V۫�Enl�򚮍H�)f�X�T�S�؉Rf�*��wn�<OhI[P�h���PRɓ]�[S֡����j��Ma�*�-+�]���L����a���E)�4�X�J���Y���T�fd�.���B��:��3Q|ATr��cI}#�{Q{�������U:���<�݉d����`��lDU�/>�ckv�dR��4l����-J�F�r��RXQj�#3B����fcN��ʇ(�e��uZ�ȍE4d�ӭ�Z��\�5F�������Qh�Flۆ��-��<C1��6��J���÷���ݩ��s+p���X���g�/fDj$J�����I�{���2�wZk܂^���\���^]Y�2:Re1n�\�v�-9�o
����wUW8j&�"�m�p�:EJ&D�oe�ĖOk��\F�a15������檦��M��ͬǊ��dYU��n�W�f�L��/ �pT�0�ψ�9�4������!&� ��KDhY6�;&f@Yʛ-^Y�B�Y0��e夾����y��2��yeܽ��Y1��#�m|��zn�o&`K�Z
ڼ-)�i�*���V�{�ӳ��y����)���6HUM֑XRy�6�w�蘒׹��J��9�� sdז1���b��z6��An�[*�v���VJ�1OP�7GA۫��B=�0�WzIMWH��\�c2шeXP���Ӕ�K˵���[3p���d���`�pd�n�
��D�R�Ymku%Cx�����J�oRZ/T�TNU]�У�:�5U�¨ڪ��J�lk��1kN�SӢ�Z{��O.��r�!*kƄ�� komܦY��ޭץ�4н�*��z�T6a�X��1`�rɁ��{��5e^R��.���/Q�^6�^C�j� IIV	K�A�bjm�ʠ�
����PR�f@e�%=8���-҉����l	B�1q���*�u��j]��Q*ě�����ahЍ��F^�c��:�(�����۲4�5Z^�auT�&0�̫����l����<*�U�.�n����ٙ�,%Q�y2�!��*�a�f��UKՖ��EZ9��Y��bN[�nѭ�Y����;�j�iA�v�TzU=)��.�V���֬HnT˘Ac\����,;�s	Gq��P]ͺ����R��vܭx�p��7�w�5��
�4a�J����6sd[��˺66���ښ*�	��Y;��*�p"�V˩nU6���x�f�W�,����5K����cX�Y��������6e��&�T�kfuQi�i��/](�#^�eSֆ1�*�[�Ō�m�R�O�zw1�Hm�2Fp�O+t(�W�7�ʦདྷ~؁u��sc+7+&:��uun�@��H^�9u-B�����@�����VEm洰L�sd��uTA�IAe��%�%1�7�S`��W����t�:�SP�,`7-H�BKTO뗺"N�϶�Xܪ:�ܥ"�$�[y�NK?f�6^ڪ���GF��fM�t��@���:,����Hq�{cX�*h�^ڣ��R��i � ��9w/)�n,Lګѳ�]n�uw�,c2�8�9�@�I�ոY7y��4���c.���*�]l�7��:	�.�֍�/+p�YD]��r�%0Q��~�3#GQ5�Jۭ��Ew��9W%lU.��f�b��e�9a	K
{������B��z��˅��0��y+)����pV.��[�ADֱ�� ��۫ ������ͧZ6�9g�@�uV�H���r�V^H^骷x��0\�Z����s>���Tus��eU٪�/ckd��7Kb����~�4r��Kܷ�/V��F4t2���%ؚ}E�S�6Ʀݍ�t
�+
����ϭ+�'4�]UV�O��
�Fԏ�`�����X��2��ѼU��b�u�T��%PU[�����Ap�6���P���m5WKiԻ��B�"	�1�Yv�iT��Gp�W����2��*�dۺ��ì�t�Ұ�6]-{��m�8r�A���o�v̨��kV�Y���u�n�zA������j���{�A7D��tdV��膭����Ш�Ӧ`�l��)���u�dH!ګH�L\�+Rћb�d�w}Ñe���X�Y֪���7v6���t��y�I]#Or�V��A#
rut.�իJ��n��Y9U�ҷ��њ�3�"�%]�n����.�5R-w�6푪]nfY:ԧ\4�;�ꃔ��(�(��*U5�ۺ)�W�&�eH�M(��ySF�$ţC�SX�K
x�`�Un�ݺ�]IC>�F�)�8jP˼�>�^�������֊��+6�Cm(�L�97*!
���kF��T�4'�7,;Mc�F����I+eX�*i��$��omH0��E�Yd�4t�A���=G*��W�7#�n�e�\��3ZW�h^��[�YXq�Yn�dGq]�
�c�sN˗nmh�6��ee�x���*�:��CM��*����3u��o�l۩�U��fh��Z�5��ŗMay��u�j�2f3�r�pUN��Y���ѹ�Ye��K76�B���Q���)(1��x����;�jȲՍm\Ū��ai[�z�5�L[��䘲<�0^m��9�TѪSY�x��/-��J��[���K�z�2�X��n���mK����WU{��i��2��d�j����Mܬu�fh�p˫�g�^�[�N`Z�:_]�c��-1U��ۚ��P�
�5��p典KuY+ia"��u���ۺ�w-��}W3,`�é��P��U,h-ٱ��1Ria�E�p��9NȻ�KM;�܃��8BPR̷���t��fY�4l^���˖,�����:d��lB��]�ux7	oF��Ma��4]��KB]R"�C��^aR����*�N���M��������]6
�Cr�F)3GK���-mhZi��T�����o�
�ڼ�����t3fn��ʪ���rY�{C`ihj���E��F�5*|�Ī6c��Cw2��Y(���dZS��J֦W��2�e��̛UVa��<�oM}3���7�F��.����EҷdK�sr�^cW��)Y�cZ���،2��P���j��*6���f�f͙!Y�Y� ��z퇅�U��qƔ��{ݖ��TRT����Y�ҕ�M�H��RYGm�lXz�ޅ1��*e��Jq����Y6�7Vc3L�ε���fYD�9VF�ZL���6ݛ4~�"�/fʫ�0�Ymz�F�WU(�9���+f
c3r�U���ye�x�k��,ш��]�n�+v�Z6j%b
Cm@uխ�5�el�����X��t�F��#��YAHu㰳!���Q˗�k��ϡf���çqc,nCj�bm�����{u"
n�+kr��k6TX�p-�($���
�������ٔ�l���q5,����<����0�oVjM�ᴃh�G-�!�U��؍T�R��KuM�$�5WLj�����b���f	yG^�Uy�Y�u�[O[�+Gnn�ۍ̋#�{v�Kj�EU�.�+�/Z����KEF:Zt�z�K;�2�nQOq�)���q��.э�1m�'4՝�3qԫI��3V<V����)�N�e*۩-�GlU�UͱwRȎ�����f1����CA�J��z'�l�n�w��BL`"� ��H(B) E  �B�I�d�P �I@��`,��d�H (HAVHE�$Y ) "� ,B,$� �d �$���
 `,!$�ή���*���.�軮�
R�)$�I�	 XHAd,$ �����AI$P�"�B$!$��) Qd$�,� X
�� HI�PYH�	�"�E$�,P���II)! ����,!	! �!H ����
HI XI�I ��@��BBAa	�$RB�HAI$ @�� HH)$
 �)$B��H�!$�BC� B�W������~'���}�*W�t�CH�`�S�Q�r��c۫��#i�w|(L��y���w T�]���X�Zw6u�,�kh�f�]�����.��-�*V;C�gly��2��f�A^����룘��2�ސX��tbŠ���WQy�;����sh�5�oA]�U�B[���7���>�5enȃ���BPך�^�F�{;���C0��ܾ����H��P�f�*��l���v�����h�YQ�^qܝ�^p�51V��5X�u�ƳtV�el�;���0��9�5f�S1��5j���e��;��X����
���볆�-��.[ܱ���tWjN'b���p�͎�A�a��_�*Ӿ�k�i�C:�^�4�e�#�-�QYڅɌRy�+�ٻ�*�����(��w�����m�r�ԣ�@|&�+�Z�ԓ�w�r	M��m���geQ�z���YLV�SQ�9�p�Û�`;�W�j����x^�w�X��1e�v�˾Gp����}W&q�.41;N"��"h�R�h�ї��uҸ]1k&�99�:��c�]^��q]��&�sO�9��rmc+)�='���2�QX�.�l�ݹ2Z��B����m���x�P�x�]Z�r���MsyÓ�sj����X;���S�WqZ��^���Б��>��fg^��ڹ�{��`ѮE�Cp�!���Ǻy����Y�H&����*}��A�9=�����׌ܶ��s��V��,���;�ZT5�l�fx��ͱb��;�Ǧ��A�1^M��+a迏r��˺������t��3eQ��s���e}�FD���S�4�k�z���(�Ǻ��3c�R��;�93�*�mн�N��W�o(P�Z��a�Xɫ�V/̻���+��[�D/������y��+*,�O[`ڼܻu�4y�^��zͻ+x܄ ���m�� �7bvYЋ�s/���U�+S����e��^v�{�;E�QܰwV�iv�J��3
�Z]�[��9��Jb��*j��C6�X��
�U�ۄ�X�����-WYEp�Ü�����LZs8�(Ԗ��a=Jo{��CƑ���0��k���:﬋"�ؿ��OS쪠�޽ါw����㖐[Y���6.P�&��S����	V�3��l^�F�҃.%g)�X��L��r��]ti��S�r���U�ΖY!`̗)έch���e�t�M8���z3����Xɖ�]�]׸�Uu�wx�8��>�)��h�^_F%��7CH5V�<�T�]*�,Q���X�Uu+N�O;rֆ���r�Ȃ�u���}�lX�-���b�(gM��1������wY��N�{�:���͕���'P�.��3]_WM���X��
�o`t��.�ش�޼�yt
�i2����֪��ͱ��������co6��C�ggC�K;�uU��dfS�{��Nяc#*�4�2ne���^e�J�T���������"��*�
�ۮ�Kj�qW�Z�����&bKoRJ�|�U����Υ���쭎t�Ik�qo31���Z���B�f�S�r��,ԍ7t+���K��yC7;��m�m�x{(U�bn`yC�^	�f<BU닱���P�9AQ˽�;�u�1�2B��k�̨.򳖚�����ǒZ��BY����7�Y�M^��j;Z�P�n��]ϮP����kr[n!4'ީ6[~N�'�Ф����ʧU�2�PN�un�b�8*�YW��ʭ��3�p���L�F���̗��KV�of_��������uY�a�β7�G��Ua%�Aw��hUx&�����X�S��ӛ_n���L��U��O ��eMz�^�c�"�p8��;['&��NpM�͹G5퇽f�Qq(�F�{�y|z�V_%$1��P��T�eˬ�4�6x�"�WUt�J�#T��^���"���ԋ�g��c+9�������mfff�ԕ՘9U���[cht����u�m�3sy����}Ev�K�]Ы��F<�Gww���ٛ�Tyw�n0G]^�K{P���/#��+so �"2^�&�>�m�ᕻ۽�*lJM3��㵨�.��۶��]�D���끚JbE��k*��y�������b���f�!*���U�N�$� k[�b�V�k1�j���[�d�x6lia�XH�m���Lˎ�(V���5���܈�#o`���-��5rºC��x�_e�ݺ�t�{Kz�1.\孳�55o	��.�#��s�6���IM�AO6i�xj��[�q|���5���nJu\yS��r[3eevtεf�ŁA��Δ�֖U�?Y[�WE�ոƗ��v��T��=:�����2���[v	�����j�7��q�v*Y�-�r�u��ŉ�&U�w,����-��Ƿ�X&��U�Y`���X+:Ԭ��*���Sſ��Lϒ��ͤ%YڛsvWUԾ��I}�c4��s9f�6�nh�͙}]n82K˘��}STBi�n����ne��W	1T`�Ǯ�`�i��d�G/��;8�r-�����-U4w.�:��$�����Y�Ұl�F�E�b��1�O%�ظp����#T���:��u�)��Wu�گ4;��Zµ6sy��p3�s�ͤ�۱O*�`9$=d?��c �X�vV�[�)�s6� �����&��]�uk01&�nU\F�s�`��P��x\k;A�!��\ڬ�{�ڒn�Vޑ��A�P�Uܭ���Q5O��K꧖��e��R���E�>X$���9U*��Q��r���2�K�rZզ��'���T���ڛ�5N��
��GAG7oI����
!Mt���a�/��*D�U�yw�N��9�(W�oqXۼU&����XH�@l�J��<��ܼ5��{�n��f�����۰Z�q���%G�5�ꥴ�qӒ���&KEv�o5m�V�ݣ[:�P&����!n����{G��΋�'3�EV=�����|�سU,��_&dde�˫�Y���I<2�A�Z��u�+PyW&r��Ah�<]f��ƺ"]-ŁrlF��:����W�VMu�	Fr=�C��W�ئ�5KDV"r�+s*�^Լ��=���q�M$x�uo8��ڷ
��k���GAZ�U�ݵZ�!T�\E^}T��Vm�Y�K�el2rx�m�,�7�4��s(��'�5%�N���L�����Z����;�Vt;�5h��oM�(+]��s�&�mwWr���˜�����)xr��"��}F�P;Csvٻ��k�������ڧ�A�b�84).�X���ɫ���	�6��
�LJþ����j�U���ݩx]�[�t�"ֱa��K'G��p���V��}��Z�E8�]�"T�$5�T�[����� �$�}����N�u�bWz;�+6��}����h����r��ͺ۴^���`̵�BɆ�f��j�ݻ�v���g���%x�7��]=T.$����LC-�6���ۮ�|��}�1_�ʼ��1%LmWb�m�d��e(�DŜ.Lw�q�6�̢-+t�79�`�6T�{3=�5z�qw+oZ	\�}�J��+rl�os�nY���gl�uv]�S7+�GF�Zx9�lل����,���n<a�='v-/�Hˬ���h(M�͂�e��GF�0.�{�nʣ�W�(�j�jt�Y}����� N�m�������ٴd�ky��z�u�K���F11+xBv1���xYG���I]*ћ��̈B�aaԻ��w|�pf�R�ތaV����5�������K�p�:sý/x�vG�wb�:�Y��yD�W
��Cj���@�����}$�I��4�X��Z���0QX1Won�û�w[N���wbPc7MUp�|D�.��Gy�r�m������R듫�U˭�ĭj�P�޵�H\"��������X�;��_U'ovv�gp+S����۹]��;�j�7�[����ڏ�-V��[[����K�����5���CW���NI��mi�v�{�fi��5L�l͵�j6X.�u*ٸ
�����Y;�C�H辱i��Y�hm�iu+EM�Ό�w/�j����b#}ITV��In:�T��2�u��ԫ��x�ɻv,c�t��"Vm���O]}Ǘe��U^n�_m�=�n�����M
gqe탽Ju*���;/1V�ə����nҖ��3B�T(�V���U�T9ǚu��o9Vb�R�ϙ#���E�]�L�ܯ�����F���K�%O���ɷ�5+G�h_c�J�R����37�wޕ�u/{r[9�;u&F�d۪,5)����/F,�8p��ǹ�75m'4�9�s^�!�c������r����]��>c���uf��ل�{�������vr�zu.��٥�͝Y�U��o:�6a�42NΪ�����O�G����H�9]�N3ÃZr�ۖ&�+[S9���yM�w�'I���Q���=K�'�yK)�Nle��̸.�Wպ8�{�N�)��i�CCv4M:��-�N�2c�&]c���CW/ΓR�$d쩅�n_���]:Wԡ<꺕ުө�4��+�f�CkY蕾��,[��9];2(�ǵ�U��{o�j�?c�Ọ4���ZY�1Wx���7(*�\�E��r�R�'�xq�x���s����]j�\��������l���W�:�y��}ֲ�oT��X� ��\�V�y.I�{.�$-�iQI��i�T���2;\�q-wok�{:`�k6�g	�IAx���i*�+���#�����ڷ1�RyZx��z���	�����]�޽�5x�}f��������w<��9��lYj\�Ǵ]�^��g�ڻu����mLǷ#=1���'�1�5or����j���Wq����;���A�;|�ݼZH�T�7E'{2U��[�z��Mu�}	i�6��
�p{�ӗ0�`�Z�d�7���:�vm��'J���e9CEl��p�6�B9����7�pBgN8�n�e)7�ĴmmU[�k*��חt�����<�����h�Z�ǐ�"6l�48������MJ�mP�׸0gY�`��a=�5vL$�on˪4ru�b��{��73�Ֆ�MWkt�ۙ�d___ͪ5�k��k�7���Wʱ��ڕ�1VZNY����_5���Q �_Z�c[�-�C"Jһ5�G
7�l�Ǖu,.�V]f
��V�UdR<uq�8oRSq+�e��	gLR�l�Sm�T	�Aj���K���]p��������u�eAy��=-]:��r^܃��yV�v]V;&(ҵg�-T��x�*��0�YlkoPpu��P���꺇Lu�leU:ɜ�;tq�r��z*	o��S�ٺ�e����cY[w��;ܽ�h�'N媬��Dj[�U4^<�q�n�^@$�ht�gS�&�T���T5�����,̸��:TuD��]ם�v�;�7N�+�a������'/;.�ftx�rk����f1��V���7J��
s6�h�a�Wzl�o�7O��o�*U;{D�;-��)��%�x�U����֨V�OD��^}�0���s-P�&���y�;�,8{Iݝ��l-��v]������Mm"B:�
;p#c��J�x�R��b�Y���.�V���R��U5�c�z���uU��+�����X���TUC�4��o!`��9��s�1m���A���\f]��<��)Z�p�C>�Bˡ��X�Օ�U ��u��0V^�u��*wu�
d�ԺI�i�s���]��İ��!��`�d�mosRu)��۬����ۛ��5�0�����c1l)�9���Y�Z��Ӂ�Wg�b��swNn˝*�\����U]cp/�u�X�_SX��w9��c�u�#Y�u0X�aEZ;��(����y׶�����}��b��ʅ����h�r�q�e�\EIY�zVgMZ��t��-c�*wus�9vet5C<���}5kV�}v��:�eYڣ��V�鸈0P��<�f��Ԫ�
a|�	��5���a�9N|�WEP�u�WU��XV�'�+N��3%7Ǎ��\^[al=��>�|����[���%%_�@���Ss-	�c�����	���'��֏]�F.���m���F��k��x3!o��m�j��J�F�ׇ���u��5*���A>�--��Wn�.}��nQ[qkն6�զޒ5gTܮݷoiUXdq�Zp�ܽ�3��[��!�wBT׫2��U�]%cz���ܬs2�t�y��uu4�݋j.8����U�v�AB=��5��}wUL����r�K�	7zgM	
��uܥ�&@��kF!�yג9�U�KHF��`�]�b�B^:�>ү;I�q���:oQ��vj5WX��z���G�qqcQ���Ꝉֺ��vn���`mr5Z�qZ�E���ݎ������F��dq���i��l��c��Z{���/��]�:ʱT�ݙ���E�_����Eh��e�����ك���٣�.��������һ�\���}ٙW�Ne������+:�W]+O�ږ7��j�vU��s
&�q^G��L7�:����8<]�������C�W�p�G�ȓX��wvQ:�ou��b�ei���]�ꆪ������(�E�U�s��7���	8~5)t��b�(���S4)���y΋U�UX0\+�hu�v�T�fЫ����Cl�{�[�`թԻsnn�8�v^���<�?�gR.�M���(�i�_"tv+v�����y�cw�{�.����f��Y}CzSvl���rͥ*��f27w,r�ɭ�Ւ�=��[�Ō�E�YFd{C����f��&��u�%�����XA�Ñ�.�M*��M%�h-����ν"mid�*7�yx�����jY���˦vV�f˽w�6��"�f���x�*-����W�K��[�*�]�r��սחZz�S�WڇR��s��ĭ����y�1�}���b]6�]����|�P�'{�vv�gVG�	Ė�4Vp<C\F�۩S��p�E+(r4)�n���w_j��� �$� �r��-� ��;A�ׁ5\�=�Ut���vm����<ú9{xn�nC�x��� u5B39#�LZaسkp��-#FU��$3F�%3I�Xd<��ų�6������$��:��w<�F�&��b��˥�x�`�*�u��Ԋ�	�p61��u�⚊�\�ivz԰���]1��Lh풭��ˍ�z��l����5��:�m����[nk<�V�/%V�C���f�kl�B�����8b{��r������Z���'v�u��=���T��nM��`P�庎l[��Md�������^>"�U�ڸ݋m�o�i�t)6!X� m���t�B�c�*1C]�����d���U�d��M뱵��[��yp�6��G[U��q����ikT-N���.5��{@{k����9�M�&�U,n�-	�;�%׹���A�%�j�qH�%ѻ6��e ��Β�u��m�m�X-�<����K�W��Ab	Y��3,�i��@m�Ls�;����s�##��ᮁ��Oi����<�T�Tp��u܌p�qvl�x���j�0fa�Ҿ��ܹ�����%�
���m �M�k*B
�s	�l���7d��
��;�9�:�%V�A1�m���j�����z�h��2I���f���&���G�^"�n�9�M&�ۇ������sɡ��i�M f�cs�QB�\v�dLU$��oO.��5�ٮ3�U��ve1� v(;r6e�Y�#MH�fhJ�Rn������H��b��IY����Y���F�J�&���]IW�M� #u����}��z�;EԦ���ٻ$�: .Ng���\��n��ʴ�9`��][C���j�M�4`��'nz�=zg�n�սD���=�oS�	R�1ūf�S���e��ˣ4n�Y��"��4���%NE�1Bl��M�ڤ���C�k�.�<��3t��8B[Ile�1�T����t`��7m0��s(�.��	��]�Nm0����BZ6d���+Xé
Mc��ba꺐�2�g�q���i�k3�[��a�`��0�T��#*��\�f!6J�4&�FԾxVx���uЂ'n�
Z�6��iu������;��yuqב�'�ȹ���<����i����"�%���{8&J���շm����X"|�Fx �݃<Z���i���v���4z���h��bD�A
�f��3��t(�f�`\�Cldۙ-�>N����J�x4R[�Sj��1Vi�	�F��0���H]�=e�$��Ϸ�]l��;�b!Q�9��<![�3F���V���6&:���ӎKn�(@�l�9v�mʤ���O)m��Z�kr��1������&㮧����>�;g�c-�:;����e��wb��m�u�n�Q�涸S�ﺮ_�����E��ȝv���nH����Pmd;v�q������	�ֻ#��sJQ�Ե1�D���@0-��b�Yq��5n��v�աR�H_n�9��ﵵ��k�Z{u��4�MN�t�\���u՛�aЈ�ݑl���]#�M4��h��F6����Z:���X���xȅ��ɱكGH�0�X�� [��6[s�q�㵘��-��V'J�������pŵ��^�C��[CG[c�����Wmپ^����"t�z<�]u�ǌ��lg��-��
��و/Y���Mmu��,��71J���@��n�W��8��/4�9��Q��;�y���O��c��a���ʏ����ٹ���m�Wh�U�7X�,�,Z_3_��g-�ieܠGCa�qi u�pa�M��]�J�8K���m��ۚX�Cif�
J���a�n�1�N��c�&�tq�ѫ�\n.v�{w�#g�6�����{uV��6z�hsᥝۆcB�`}vlr�s�l��0��lƛZC,��
K�0�kn�0s4��=:�nSm�۞���낎1�ŷ�d+��i�:,�;v���U���ʷ��e#�����S<�d ��[rph�WMM�.�]����JU2[m�d,sv�m�Kz��y6����������c�wd�]�n�5��te��&��4B���s��D`ޢ�ch{`t!��͎�+k�J���-���m�of�����jp��m�^�	���-�t��{=&=��@����,�/lA��J3��u:4
]�i�k��Hfv��8ۀpoec�^�en+@X����.�Lܻn�t�D[@���R�A�.�lr��ĝn5�P���%���6��N�&�(SY`G`��[���۶��sq��;j�ĥ�� 	k������{LNm��G<
\b�{�u��V�5�d3�Q�cp	��.�NviF���1��ٹԺ�8���v�������&�]Fv��ݝ��ǧ��H�miWtv ���96拭vrv�n��a���{س����&�����[vK7Z����k�nj-&��blĔ�� ���㇫�`�X����&kll��3��Q��i��b&��E�6�:���	r�Sȕ�Ϯ�N���<�=�;969R��z�S��c	\�M��B����Su�p��{�Xrvӎ�n�C��#�e��
ho�F�����T��B$�sMj�9��#���W�m���5�� �Y�v�����	#�݄�P/��v��MI��Q�6��l�bXM4I�&�W�n�;gsQ�f�j����n��0�X�c�o6�����/8���ʷ������W|�xH���o\�+`�56�n��M{&����F�0��wE6�m�t�9;\�#�I���2�.���x�h���ͅ6��n�8Su��g��et��꫈{��΁�CW��k���Z�� `�BY�tu;T��a�Z����sRR���:���'��13c���4Y�v����,NZ�'y:��/��bg�[v�zC�`�.�)�8P:h��v��(�gV����Y5Ў��EA����5����H����U��<h��^�.}�\j��.8���nr`�>5u<`a'b^��{F�vѾ#���Y�;��S�.�ڱ�b�l����	s�z��,��z�q��۶����i��#�X�ev�,��H�A��|��M��#�]�`��s@�j��m#���x��7��M�,�^w��F+ۄD�<���ŗt���&��HhQ�歸v�[H<YD�ݞ1q��ɥ��Z�prV�9'��C����i�З1�G8��W�Ku��@�t�cvZn.�����n5	��{�zx�^�k�����CB�hU�hF`dipt�vWbX)1l��&O �ލ�V��3�l���N*맧&T�خh^���6ջ�'t����ݺHz�P�㳍���WLV&��ڇ�Θ�E����֓�cq�2�'c�v��!����hҎm���z�F���l��u�i�F8��3\��aϤ�i
ݺ�y-j9�s���s�;y�Mۏ�_|v���}�5c:��gq]E�qn�yC�6ѭ�M�i���]�Nֵk(��8\�m����A��nմ"]�If���Ԍ&�Δf��#�ƬE��<�0x�d:�do����C�=���{�[\��pt3
�s�bR[��[iCtA�j�ӷo)5�/RXx�\��t�Mn�4�ؠ�\GG��Lll��4r�
����H�ɹ�A�y�=v�8�5�yL�����§FGTgQyQ��o	�������˼\j��](�k���d9*����ŋ>�r,v�/V_=��s���/h�<�i��r�����W<ώ��x��ymUs��4��:^̴m�lR9�-`�7;�ǜ�R�-��#������ޓ�F��ʘ�Ŷ�]�ە�v�8�8��rM�dl��n�N#m�#lg`}Q�f	.�oi�n����Z��`���)��=g�Ջ;��{I[����	���n����MËa�;[o`��u�ۺ���i5u�K[1cK��FС[��`���`Ӻ�$0[P�`Y��(e14u�,���k����b���+q���1,Y�d�ޮ��.������2�I���ѥSм��m�l���Z�cn���8��I̶$]�2�@;*Ц�m��8�Z�i6�IE`Eդq^�Ħ�J�=�;�pj��+؝tݮ5�sݚ�f�jy�7c��<Z�y�@�:U1|�T�9�:BGWm��#
�O-s��fx\n�!G0�B��&5i�ܠ%��*�A�k�bRl�f��ue��ss�;U�F۵:6��J��]�(��~ g��"��g]n���j����ǀ����K���A�7�z9��/f�)�^�"��ּ�j��ѭ�t�]Q���;9$N������Q�`dv��0t�F��7f�mۆ���c5�ڝ�9y�G`��f�܏���C՞rv��xŒ��8_(6	uj9����>ۆ��ݭc��]dx�G���=�o�Q�%q
A�9�Z�L�\Ale� �u�&�v{����+���g�*��OU��7 %�,�d^x���-���s�IaZ6\�cc ���Y�M��2�eQѸ�B�ku�Ӹ^�N��ӫ��#h�װ�Hَn�=��n%�(�E�!��ShM�j6��ٳ�`}�љ�9z��
�C3a�v��e3���-7H��[�v8�&a�28�x��j��`��ݵ�Q�7P��8[�h�qgj���܃�cmZN�8�ae��z̼]�5���2�[.�+�J�ʡUq�$�3���;u�㧌��e���p�۩���u3L�4	۴4 �Ε�K������c:�3���^�=j� ��SӸ���T���Ö��^�kb�2鬥h�q��
u!��XH�XQ0X2�L�k�g�_g!�n���n+��6����v3{U�8�}��m��i������*����]����w�'��B�	��t\	ޱ��)�k[bq�$]�Օ�L�;�� #��2���9�Y��e�ۭ6ǽ���99=�{���i�3$WHM�m��\��"*��2���.N�<�G�a��̽�D9sv�췘��Ş^E��N��HN��[j�E�tf��l����;���n)9�drw��׵��QQȶ�˳��Ȋ;��b
�⬬����;�;)�y�sn��v�\U�y�e�kl^qu�Ue�i�֔NE"oz��w^W�yYݙtOn���&��h�ˑ �2B�7���vdt{��T�j�wv2�8���xY�e�6���Ք6�8�=��!{V�N���Q�E�zt�ӓ����^p{d�dq�XRHU�uWs��U�D��l	�޷v�v����ͪvS��	�ps��������v�V-�Mu6fG���R�dt�0��k�����+ؑ�q�� 6M��p2�BX�K��b�LO���Z4n��ct�F<�����n���M����v���۶�������m�t��܄���1S�����"Ѥ@⽞�pn�����h���q�iq�q��֗ϭC�^LV��:�2�%΍�㶦��YR�9iRa�Usb ��.�S5��m��g"��=v���&n��Ɨ�/dϩ؞�[�s�2��Wh��3��h�Զ���j��۹�Ǳ��y��65cE�]aR� ��Tt"8t�F>�ݎ�&�8�b��`�;WR�G�^��nqڬc�^;:$/	J�B�R��j`��m�4GOr�(x�ý��ySgP�4�جr.z�c{d�xa奮m.�����$cMK�i��P����l����ۯ!�ђl����)������u�]�S{]���c���`{-�4.��d-��q���u��+��zm��r�����t=��\�&қa��,�ΰ��e�]6뭷��ɵӍv�1S>M��8�n����=���t.G+��m&�0�¬���cvƓ����h8��LW&�[g)�6���	������pmՑ���ӫ���b\vC��@��W=8��^�C`��֢8�˞��XJ�F����e!Xf��	;��uk�a4O>^�c�s��\�p6�02���ن�gaD��E�̰F���s�^��=7odEᘪ�B�,A�m-�"K�z�p<�g�ސ2X�g��d�2Uͯ���1��&s�7�G)�sd���ɺ�0q`�F;]
�ѻ\sK�p�>��;E��G'�������*t�'Q�8�u��c]�����ze���9��Ѷ����R����v�=�mB���3���kGh�i�I��cJ�Hj�D%cc�Z�-�clD,�[XF��K��R��X��Dy��Q��e��B���R[e���k���<������@�C��"��Ue��j�oV�E�B�фE�"�Ic
G��!�兴�I/Q�-�K*�BVՅ"�PjѶ�%�Z�����e��5��Z!�*�f�\�6S�|��u����4vp���`�@����p}�����[TA��b�ގ�=�O{sEI>�8��7-�-���7)������Jd�d!_fW�.�����b�ޫ �!O3v:��/I�������s���������w8�]س� ���A�X��A|@�X�Vgl(�έ�r����tY6�}�%IV$C��/�,ة���eUP�������IA�z;4�{//f�+m���֩"E�*+woo�lGſX�$� ��|A�X�d���ܽ=�`@���eouI�������ru#���U�d�wR}�;[�h�+�"Nu��WD]�.�X�h�33M�e�l�P� �l�n�[�Gv������s��@��N�M^ȍ�e��쥤*�s�l
�D?�"�X������aI��2JJ�r�}�.�߶]]��l�*��wB��Tͺܷ>��o����=�$޾��dxv��ִf�vt���U_�Yٰ�����������+v�~�Ub�9bý�g��q���a�����ĒD����e#W���q��2rD�mI�"$�,�*� �G�
}�W/]ON���M��z�}�xX''P I*���N�Y����ܣ����sN�������? �}�M����7_i��{�Ǿ��1�Rs���嘈�����p��,�WM���zŻp�{�W��O���<�����?D��%���0}w�M졏j��T��B��'�.�<uRQl,#
�lgY�ׅ2��`�������,����'K���"V�O+}�{�����h�9Uq�)����H��תA$�g�B2J�2��V��e!5A`��|~�,X�}�<���&�tY6�� a@k2D���6�Cs;��W�d�	/�B� �FIVD��֚��.��o�&���ʹ��3k�2����_E��jD���]g�L�D��N��KV�$ً�>k�a���ɬ���^AjCv����`/�Ŧ��E:j������_{}_XK�/����W�׷��{p�0͂ْŝ���
6�G�{���m��9�㓨_�u���Z�͢4&ՀD}B�� �2J�"Ib���3�>�t4�5g? ���ͯ�d�%Y	k|���m$�P$qV	ö��B�6�ۆ�ۘ�
uK�]�t������R�T��Pz��P� ���$�oZ�������O���!�W�v�a���"��dgh*0�9�<�/N3f��A՗vodլ`8�X8��oTx���|6�s��=d�A�/�������w����v,��}��D����I,Z]i]��pj�Ϲɺ�_ܽ��ͯ	Q%��*�?
"IB����˳w��P�A���g�}rK�{��ګ/}v�����Z��=Yu/�*�{`�S��rY-[�	���F^�S�̻wgn�Z4M�hJϷ���ur[k�nQ��*t4<,`�ݾ?j_ޖ,%}`�QIb��UX�^w z����!��ݵ�
��α��?!|d�D����6�j�ഠD�j��c����_m��&x��$c���}s�'��zGZ�k;҄u߯����r���9�=��{"k~��6�+)i�ՐT�M�Y����rW��|D��$������w!�a~ڲ7������ڪ?cb�o�h�N֩���B@?`.#R�V�P����c�`�P �/�%2	��搈�B�K�{7I�^aUݷ����k��0%Y�%���Cٹ��.��]W~�,_��K�$��-�aw�A�@Wt�f��aD��Ô�{��3��U�A��(�%��$�`�_$�]WJ.�ګ��xfK���ڪ?=b���<�>�U�r��~���X����j��a�Χf���g�(ON��}�c��⑱���:v�[����QMZ��j����շ��>�D�D��eb�}�8�����]H�*�S�c�Qs�Qb�`���a6�g�7#\����fx��g��� m��<��P�e�d���2��#��2`�wԝX9���/�s�3�W��51j��>x�{d����g>�B�џqY��X��n؅��5"n� �]�l�1ļ)-e�:�;=�`K+)�6֛j�4��<SN���kiB8���}�Ϗ�լ�ڤV�#�ipR�t[�M{u��L.�R�*�TQ����@Ҿ"?P�$�!@<�9-��b���wݯ��M�����B#��9x#�s��/9*�ta��pymm?4�wu������~O�]$[6�@;%�I]�3e=���V�3搐o5	�#$� �%����ϩ֧���Q�lӝ�g��}VA�9b��/��Ń$����rߌp�o��� �h7��䷾�5��[}�s~	��,�f-����d��}P��_���IVAK�%<�����)|j�����o�y��k�H�(X2J�AC}��n�����:�_����+m��:!��l�[c{�%;2�5�l3'CQ�6�]j�c�ϳK/������#$���Ňu�;��j���4�w���M��y�wP^��& �2K�IL�D+�F_oD����E�36�kßl���y��{@i�͌�&F'v�h�
-|&��ۛ��L
�]��5�u����������J�c~��z�A��7%�e��^ƛ�������'�/��������Y�z�fc�`�� ����%�&/����b�ެE���o|��+��=\�[6�A#
���d�d~�e���}k��f�P����U�AIb���ﯼv�y���?�`��R����ؗ?B>�АrJ��B�?I/�%{�Yfơ�E��D�\�|�/cM�}�|�ru���2J��X�u�_�(��-�P�6]:�t$�x�n������K�٢Zf0�1u�z�Ҧ�����y��TNs�eW��1g���@Wl�fׁ�C�Ø���1!0C�7��U�H�$�I(_�uqvV��$_�n��7dM����Ҭ۱��w���=����$���1qT��۱�_Y���,%Y�\�C� lHY��r�Ԧ*��K�9�X���P��td�)f�4m�w_{��a�NT(ȹ�d�(+��w�٩���7�X��U�$�q��Q���o��o*�5뾈��#=A_I(XK��K�t�z�z)�^���|G�gw�ֽ�ׯ�4����j'9̓<�dFII]^w/`�~���eo�g���66���|?�U��+�1}$�Ҷ�j��p�\ ���f���� ����)l��|��3R���0��S\���IC&�7��Yz�� ��b��U�	���ѓ�G�9�n���!��>��X��XfP�>"�j�"Ib��/��J���32���0��zp���b�O�"�j�}����{�a@�6K���<ӹ�W ��=�vǜ�`�a�$�$��j���=<Z��lKrsc)���}����K~�|D�Ń$�#=��4�u*�`f����!A�h�;6{'���}�v���P�D#M�ްR�Bw��	����/��|(��;e5i烅>bR�.w	���n���D
:G:�����>�!�/yWY�Ҭ��_	� ~2J�D����ƻ�.�����,%�I^�XO�"9�*fׁ�6Jd�d!Mӿn���u��	dD�Q����qAǶ�F�=9y�Ӯ�5���f�֎i��d?O{��,��P�� �@�+�X����v�-�o1��w��F�۫Cb��<� �9س�%��Ib̒��A��Qco�n��:�-��q��4dݗ���כ��nxX �z��~��+�q���ƴ@������S�$�,�_$�=�v�ѺnWn+'�";�*fׁ��,Y�U�!@�%�%�@ȣ$��Q��AH_�}$���z=7�nv��w}�@�fz�������n�z���/����*�A�X�d���%^�Mn��(����G}=k����<,�� �������'��6�������� ��μ�f�]W֜���2�2�5����2���@Ir�ӎ-�&0��f$;.���Q�{�������k3f�R��VEvVk�x�p�O��<�0�����`GD�l�!l��1������܉��HT^Ĩ�ڳ2r/j5���5���c�Y��Rp��ۧv#�|�;S�����K��<.��gj�0�$�ǳ�ś��mqn`* +ƚW��K2�Av%`U��h�\�uEe��"�4��f��Hj�8y��=D�YY��q'"m��i]Rf:�-��O^��Pݨ�m��_������5��Ƿh��S� u<Yx�Oi���S-g.���D;��a�s��B/��wޕ$M��R�6�=0;|b'5�0{�^"�j'9̘#�r�?&��U��#y�d�zŵ^��ҫ}N���V���RE<BO�b�!9U�Ŧ��Ϝ�b�l�8�$�,%_�x�<Ղ_e�p�����޼���{}@Y��*�J�LCy.�A7}F����zX��A|d��<��]_��,��S6�A#
����Q߽�@;�VA"�K����A�2J�\״���M	�Я-��
���O���o�	�����?`K'�w��جg�)��R��F����F���9��`�D��A����ʦae�}o�����z��=�f��� ����F���||�]�w�3����~e?g��f�S����9��0�*�T#�����������e.�[}�
r�No"��.�v�-U;,���c�v�U��no�ip9�U��F���8^��ڢ���SG\e�~��1���Ｒ���������� ��c�,%:��z��m�złw�B�B2J�K�����vήɮ���c�/9�}�@���oJ~��$�,%Y�}k���!�a�s��oW� �!C&��o����޻�ﷳ�	��?nm�cO������9�3�P����G��/�����c�}S���`������p��t��^��(Y�U��B}:*mT�WN��1R`$
D!*fK���u�IlՊ8a��	[bgK�����1��4�?P�A ��*�Ia���K���{Lϝ��l	!Ln�*C{�S���"A��|d����|D(���z'?[���:�Y��F����}귯7��yCK�BH'O٘�l�f�;��C�x/n�K>���o �9�1����,$�;w�ܻ��o�S��T��e�^�t6��%��]Ϋ�Ƀ��U���j��2uFMm��RR����E#$=�f��Q/Lo���ةJ�j��hE���ɓ�s�U$��>�0��\��r��4xajgm�ʚ]C�^G5�`��#j�V5W(M��u���ըi��9���K3$U���t�`��XW��}f�\�6�z�Z'9���2`�I|����o�=�T#:]�m�����h�)F>�{�Vԧ�j�l9T�P��X������_5h#O���C�V-��g¼G��EG���o����ڰy�Rl]G�1�6-t��j�V��'N�{Y�u��b��>}}W%���t�6�IŪ�>�Lm5���d٭�j{Q���x1�KYN�Un�F2x\���|�i�Bil�A:7\h���p���Pۮ�u��1+����.�2d.뉔��ԏ�����2�t3�fq�&y��_n�7�I��+�7y�o�,�m;��	A����of��'YV�ޡZkX���2��Z���v#}}��v�.y�5N�z�o^Z���z�Ζv�V������j.�Z�(^��0hyV�i:=�1�Ufn3�����K�v:��Z2���b��E�W�X�s�a}ʍh3�K*e�2�&�d�33�H���/�0_$$�Tz+*����*�2:�V����,�uw�[6nE�t^��^]Wdl���}�;�6ѮIYv]��e��S#��3LȖ�9��Jj�\��r�3��;��kr����.�efi �6���,fi��G�*�ϳN͛)m0�'���:֏��(��Qb�T��X)�t�a8%����9�f�E�j��@�d^e�6���l�<��<���y�.m���6"�s�N�-��6�A��׶��m��������f��Y��e����I-ۣ��+�pw��IM���u�{�޷��-�{[:��B�죠�ʴC���(�!<켵�g������$Q�n�l��V���Yy��xڻkQS-E���ym����s��	9�[%^y��C۫)6�]<k"�V\6�̊��J��(�"��fv\�c�I�/
�TVu�qq��ZskN��u�VGeg��������qdQq��e�y׭�Y��qRH^wll����w�ί^�Geeg��w���Ɣv�:�༬ꈸ�N'�r�[n��,��8����g9�j�˓��vt]�4��xû��Kk�O�� �t,��$S%/�����XT�{��Aa�� w��i
H){P) ��l>I �y�����g�����bA����^��R�)��޸bAH(i��i ��������������k���y ��?0���Xw�\1 �
��w�:}|�[�����H,4�W��� ���\1 �����M RAe�������§{܆�
A@�{f$�
Ad�)}P)�k�<~���{���o_s��H,=Ϯ�R����Y�E��ԯ��
Z0�{p�i��
!���${�������_��k��X5�d�F�m\FU�G<��G]s��!۴�ꬬ��˿��A\����
J�So�H)]�p�AH){P) ��n�^��o���Y������w��H�vb~) ��}��{ܓ��@�:$���y$�)}���Q
H,��^�
@�JH,;��j:H)
*��{f$J!I�^k���{�) ��
a��p�i��
�;�4�Xh�f����_���w�����H+��- ��)����
A@�߻��M$�@�Y�9C��翽�
A�B�~�i �`R�r�M�YC%/�!q%$w��i ��
@�{f$�B���~�\|������w�r�B�6k>��ϵ��|��H,=߮�R�P��1 ��Z%z�RAK)�{ۆ3C%$(�{f�) �h-��������G��~�.�є�P?~�f$�IT�D�U��$E��9�~�k3�~����y��;����) ��)~��R���oף7�k>�۪���|�����hة�V��0`Ҧ-���n���q�b�2�W�&�ׁ�2�Mzo�*��Ϯ�)�Ы%��.��|	�w�)�v�I��$J����.%$�l4� �*���bAH)��@����L;��1�	�>6�����5��O���-�N�]��^h Q0�w�A�w�dBq�D�?�@�ݵ��~bMX�$�Ҽ�1�6�m�-� )^wl�u�6��kj�@޿Y�� RAe2S��HX��
?{�$�����H)~��? �ض6\��MM߯;�"{�$����~�W�[�@�嘐R
A~`RAM�S��f�%$��bAa��$�!L;��1 ������~�~�o}��x�AH)��tAH5P�?\4��>�ge��{�=�b�M�|�ա$r$P�O�
B�%$�w!���C
@�{f$��g�g�߽�� �X�x��������P?s���R
Az���� S��f�) �B�l�Aa��_s��*Lz���{6}�^uy�.���H�G� �R�n�R
�~�H,4�^�) ��w��i �#�����@G�����.Ƿ�X�U�m~�O����X}�\1 ��
@��ى �i���H���������k7��=�H,=�?�
B�P��1 ���������8���AN�S��f�) �Hs�l�Aa��$�X��
J��nɡ��P+��H) �`s/��?k﮲sG���=	�_�&/6�ﵙ��w��_{�@�~ݘ���(d��!bJH,(�{��Aa�� w��j!I��)��/�}b������?�H��X�^[3"Z:ľnܪW�vI�Zڱi5Y:���WQ�ރ���n��_ҫ
��5��c������KP�q-�M�	,&�ٳtny���]��zv��q'�<�6��[i�=��Χ�2���	����cj٦`B棙@k6�eƐss�hP��h7<��t8��e��F=�$ec1��JF�����5c��u���)HZB2�[����vi�h��tQ��sm�PF��,�����������YY�ޥ��i�#4�8��Zp��z�e:]R�٣خ)��d?�՝-���̟�t�R*��f$Q
H-Wn$��L;��1�d������H'�����_E{�y�][�$�|�RpϽ��{ǧ��~��x�\1���H(��1 �44�W��肐h�w��i �`R{�1 �i�����RAa���wߨ��2��R��1&�) �S)G�A  2��F����ޛ�����?ڰ�� �*�o���tB�U�I. S��f���W����rm �q��4�XhaI~����
J�S~�p�M2�
w��I���
��YtAH4T;��4�&�X�f3XX�/��}�6��<@�����I��K�@�,II�w��i ��;�ى4�$JKځH��Xw���t�Rsڳϛ��
��bA��RAh�\
H)q�{ݸc42RA@�{f$R���u��^Fyվ�iMG�AH,3��bAH(��}[�+�ƿ[���M$�P.肐X{���R
{�18�I�){P)II��rH,5R{�1%�y_���z�w��H)uP)�^[��?mק��^wG����@q�HUP��1 ��W��
Aa����d���!���$~�n��{:�������֡I,iv��OT��[���IC,è#l��г����t����ጞ����S��H,$�@���l�w��i �����=��J}-��U�$|	~׹G�o��'U�
Aa����i ��?~혓B�R
��RĤ�ý��
CEP�lĂ�H�r<�g�fT~�&\��geИ
��dώ�T�՜���G2�wFa#�`-C�gC������s��t�]"�{=��<jXOԥ{ΦQ;� ���)�����JH(�lĂ��w{������wo�G��Q�G���.��2�
���A`i�������W7�
A�P���$L
@��Y���)���@���X_{܆�0���bMR>���O/�Do�W�;w
�nSK7s��̾m���
Aa�n� �w�Y����W��
Z0�{pĂ�PЇ{�4�XhaS�Eo��w�cޅz� �܉?8����j���G���J�3��3k�0��r�E��cs� ��I.��P�A������"����,r���y�/7�)��w�G��+��	�/��K�U�4.{)R�޼��~��-խc%A�=���ӵ�]�lNy5���i �3\���a_�ߧ����,��~�K$� B�ݍ/K�����7=����/��`�j�C����9VI	�/���������rv�����">#wdM��FޏzwGUn_N�ͯ~#�s�,�*;��B��@�P#/(Y��Y�@�*�"Ibe���םGS�6�Xy�p��Ty7.��L�;���U����t��ԉ�B�M�����6{]ap@�p����^JZ#
�=еk�hvJ�i�L9yR��������nԑ��7�͜�w�� M�U��X��K�$�`�*�!��U~�����nD�o��=Yq�U�*v��o��D�|�	"�|�$��Aw�_X��L@�%}bIb��6�{�����w"i\�;��N�iUK�>�- �F�(Y�U�	�C#hb�5$Ζߥ6�9�f�;Vj�mF�$`��6-��lI�C`eS�ʼ2���×�L��f"R��*��b�V���u�y��s}�o�A+�s�q��H�u?x���X�$� �
k�:�������@@���}/wյ�-��?����IH�^;�Wl=��W�k5CC�b�� A��YIb��_%��_���mQ�:gz��ʿxuV������
 �,%}`�W�I.��o��*��0A8B=:���Ō�V������2�շ�l��"���ꃦ��y��A���Y�-y��weԡ1�!3Ryザ�k���z��r���f�UeH���En`5F�t?����܆��7��ds���Ɠ��9��BUŜ�u�b�#�v�s��|u�ﵿX'��,�x�d���/�y:�N���!s��r���^pQ�Y{f�fJ�ؚE�#�F�YQi�3�~B[翮�|��^�x��j���$���i6�KOޔ�ī�� ��`�<�Ń'�� ��L2J �Z�<»�!�k=Vޔ/U��7}��um�[{Z��~�;T,�ǻ���L8�D���$�!�Ӛ���;�9���[ks�cu�gP�!%}$��� �^��_����,�~RKo�G=��Ww[�^E �/iм�:#V�ՊA� "Ib�2J ��U_�Y|(�:�
Z����,b������=#�}�o�@���w�b��/��X랗z�F�R����^M�`�.��u���8T�9�FS_>�������Z}�޵b��/��/ds=�Ĭ��+n|T;we�s����5~~���%^�F��c�x��uy�#���9�c�/��F����0�q���^�<����˘��0;Z�#z�D΂�e�f��%vAm����MuGEe���		�)�1�,�m0�Lcu�3�T����=cv�����C@/Z2���ئ5k��.�-��Efw5pq]�vh��nɮ�̩Mm�S�ԁ���N�î���U������n.w����?��jb�&�r�0�Ku��PKs���.
55`�S+��Y������:Џ{�0y�^"�h&��o���s�c~�׋Wp��V���(y�^Dy�a��J�9s���܉��4�P#�z��3�@���I�Cn�:� i�G/�%{En@k*�d' G���[�,�a�$�%��P�e����~�z����y�����@ ��$�"~?d}̑ �b���5����
tS��9[_H#����v�k�1�=�G�o�Xxl���HE�r�߽��/9��g9�0g(�q������YQ��n�NM<k=k~
(��fIV����ڮڪ��R���=u�H��i�k��e�oS�d�s�U�y�n!2��r�.�.�E�ކ�r���+�K1m�۵���2Nv���|��9���-�|A�;���ř%Y�!@���uw���K��Z�7N�E�t��2��n�X�A�8;�R�H:R�3H4p*���_��I���݇�{5�ݱ�y�ąz��1Q���� | �ٲ8��~ ��*��;\��=wy�d~����!%)�D�8�yC��HzJ��X�~��$�Q�������8.z�nt���4���,�+�$�3�a�Uޓ^�]��w�V�P��;s۽k��/�:}�o�@���dd�F�u}��b��҅�$��A���W�J�����o�W�P"��Xusz��=n{뎾�����2J����s}��5�|����B��_Q�7��`������zԘw����-���g��}zq���,��IC �y�̟���Ν9V����{Ya�0����Ȑo�A"�K�~2Jp�w�J\�?L���l��۞��^�i}����< ��X#}��LΪSEK�A�~��3ޫ8�Kd���D6/ۘku��5hD�w.⋛�k_��V-�RrFn�����U�h�Hr��k����?oևm�U�T=~s5e$���]<���|>�JC��a�]M�o��� ��BQ%9���9fFr�)~�k��f��zJu���Y� �2K�o��>�eS�u�u�	Q[�m�nU�@"�X�L�������w˽���V!{/6����6ߩ[x�>�W׾��&����R�eVk�fuwT��w/g��s3<��r�B �V�SS6$M	Y�)��2���5I�A"��r$�R
�� u��/={m�}�k�C�,����Ͻ�l�y(}�� ��s�(C��A�+��K~~���hJ��N��}��͝�xH��r�|d���K��(ډ�˜�,؋�s��Dy�aSڱLa���Wh�:6ߩc{D}�����Ń�A|D������YT����t~��,�d��34@��|��;n{���B����(�����v��??��'}�/ކ��R�����qV*X�i��9��|�[:��2Up���$O�gr�N��n)7�{��U����Ӈ�I$��O��^Dy�a�9E�r�#9�a��a����d���
�jy��]��͝�x4��7,I��?H�*c;N4�"!�(�+����1�-ցs/�\֦8����9����<�Y^��l��Y���I(au'��>�*��,o�o�"���[

92�X���%�X�d���!_4̾�7��ՂD�i��V?��f�L�/7�m�}�|,�{�,A��$��8���4�A�X��!~�I(Y�/��J�LJf�:�_�:�nų�㯼F�nW�J`�D+�$�bL3P���ª��CA�HE�U�d�/�=�����ݛS���\���2��_�=U�>�TM�dy�VD���%J�ןmVQE}��n�Ξn7=���X �B�'� d�D���j�,�����,��wd�'sl��%j�}'P���2e�v��3����Ӽ���Z�ss���r��Ρ��ϲ�αP�ݱJ�3c7�������8\)v���*�4�h!��W�WQ=j]�p����a;09|Une�亞��ʍ�o���Vm�᫝s>3��FɪGh���HX[�����䧼���J�
�"��&��Xo+��՜�#�2d�!r; ˻����c��7ؾ=�n���5ݚ�{:vp\��
k�ti�)ي��ԝ7��ʓ.�Z��Eo�VfFz��K���S�c'EU�m�h�J�%Mel���"��W��R�WS���$���}N��C]5�{s�����#��W�.$*m.�A5ԮS\*���}�Q�x���ӇB��|E��␅����q]2y*�vƻ�Gs�U�re㖱(&m��EW>6^.�[��m���6�+v���n���SO&�$�gnX�ż���
ר��t]ͽwW/����n� �4��0ܹ�pqI���S�N���7�U��SV%K�*������#t��skM��v�����xu'r���.��L�΄����:ٮ�|ח���n�N��N���C�IvX7P7�s��P���cϘ8�1u�����e�:t�^���w�ܥV*=ZSwL�sI��&˙�̾o+�u�t�@��e^�#�K/.�f�pc�ک*Cz^��I���w�ڀ�X�vunV��Qƪ��B��#ֻ���'R�S�R1�y8+9�;E�חL˺��5"6R5�Nsm����i���]�o�#u�]�""1wf\t�~5�i��\ۻ�mVW��{׵��;:Ί${��⓻�Ӕ<����mv�rw�ۅ�X�'O{סGG@���k)ʓ�]E�Qŗ����ub��N��ΰ�����Ȝ�
L�����[n9.,ˎ�8�#����IN\��^nA�W��yv%��η�nΰ�*�(��9����s�fY�T�v��v�tG���e�Yu��jȣҰ����x���YfW����8����yv��y"Fue���⴫3�.,��qqI[h��c]ggq8�n���:��tGE�rPw��Q�w��Pw���F�N����+��K���;;��ENM�my�tv]��)�ҕ��0X)?V�}|ˤ�1�-��ƱU��A�t׉���,n#����,5��m�r&0�z$��l��a䳮�8lrW�I#LM���'��U*�06�g����:�;v �씛q�.��M��&J5�	�f5�&cS��
�iN0�õ�f^��'][��ֻ�M#�����dv)�=r�GG���j��dy�5�X��NV�[F7d�n����f*�J.��R4N��#���{K�`�n��M�Z��1=����۵Q�vr��sU�%�e�X=�P���1���ƍ�eG�~��И�W6v������Y���3�lR��㣯6���خs�e��N���
g@��u�Z����W!ssi,b� P�eU�[�ɋr@���\��t��U��`�-��cp��
��P��;��	 e	�g+�N�����8T{sÐ賫�MI�\�ю�K�;Kv�v�����.$#����7�<Ѡ�pu�=`��S��ez�G✐��ƻmɸi���0V��mUe��� ��qk%�eĻh6T���$�+MO�[�R^�=`�(���X�y{|����m���nX��"�8)�c�[�rr�s��5��=�r��:d+�1uTF��5��.��^J��:*�R�Y`���Tar2������[y�5����8�9��B-e��1�:�ښ�ڷ������;F�sH���]#�3�z���u۰����k�O;[5<k
��3��y�*ݢ�ű��z�uenw�ɭ];�y��\ F�,+�eu�g�374P�[@��e��̀�U�\Wx8y4�����`;lT��3
³���	�p�[�@���R�%Y<����[��덭�;F�J�V�1�<E�M������M�Sd��l(/�9K�B���\��u�� ��9�e ����DIk��75.ynv����v���vu�ł]G��2i�Rn��
Ս#�.��mĺ���y3\v�n�U.p�sf�v��m6}N��t���y��ȝpꋂ���-v�,�����ٴ!�n�a���Y[2M�-4-�Κ��6�c�}��]�' �l�lb��t/b�Lu�ġ�[m3�[A��;�f]�\]3[�GSc�����8�&$��v�E���ugw	���E��p\�)��u���4����HC�N͌z��O=Z��+X�qq;g]n����4�֖�X�������2�K����f��m���蹃��[\�p7���չ�f'���,�|��g߿(X?D�?I,_Ֆ}�Ǒ���݋ge�^{���!�s�<��4�b�r��"fO�9���j�\��+5Y�q��u���Nؘ���ݛS������ ���9�=�ꗷ=�١��y�#��ř%_���A~��4�K���ͱ ����<�o�����:A��%`$�`�@�uL�b
�[}\�����g�_����YgϘ�Wު[�l�k�4�En�ɗ~�V�^�7_YQK����(YB��*N�W�Md_��qct]�N�7�h�A�jA��X���I,=�����S���u0���;v�A��{1W9:MѸ�nݚ���ŕ�viSy_awK��!C&��	�nm��j�މ	l�t�M	��nϑ~g��Ќ�9��P��9s����ε�ۊ�;��s�x۬W���b����ok,��z�>r����IK|�SGn���|����2�+���~���[��Y\���@�9���=�YG�������X���(� �w��f,mɟk���\�e�C�ȐM�$!%YI,<'(���F���߳���҆:�o~�����s��3��]��'4�Б
2͂~�~�%�W��d��o��ܽo����`�yвMz�z0hd��B� ��,�%YI,Y�N��o�4t7���Y�F8+��Vǵ:����ܡfIV !�PxK�px���O
���u�kX7��f�,�mp���3ؤ��k���i&�&�`�u���~�/����$�x���1ctK�.���B��Z�b��uX��Y����,Y�U�H�.��,�a�}W��(ɣ ���/[��;_7HH���2=������;���Y�7R�;���9f9U�9�!{+����LA�C��^�T���́1V���BY�a+1m�펅���2�tn�y�9�m�T�]��|��k����O5�BUW�]��| �s� �g��cڝre~ ��|AnX�d�d��$��U�4��hѧ3;�@~��*�"Ib�<���=�������s����v�Ns|j���4X������ւ!�Am�ͧ�n[�"����}�:y�m�s��t<{΅�A>!%}rK�f�F��ŇO���*�%+�����5x򯐗2�)
A�:�l��n��FU��뾏�R��=�"A�љ�$/Iw\N�R��'\y^ ��y���v�%kpC#3�Y�����_�2JV�ڶ�U� -Iۑ>��f����_��7���ͩ �Y���ލ�Q;5ꋛ;�}w�b�-���(d�/�$��=\��ukS���nd�;����7;��C���|<F|d�`�$�/��K����ǃ���j� zK~��$�.��?0}��m\Ǔ�<�|$iD9u��K�ա,Mx�0��$GhWX�J�20��V�h ���VMҽw�V�5���]�ٴ�E�y^^�oc���A��w�mˋ҆[H�J_�Iz������D�М�00G�兘~�R;��sA�WeZ�Y��&u1�ó^����������_I(@l���>{�]�z�_n���j�B�Ў�a��Y1u��im\�n���B�d�a�.�
ߛ�o���@��P�d�dD(fI�f{��V�7;������*��,��U��ş�@�%|p�5>��P��Ú����ʝ/��:j�<�Q�x4���P�dħ4ЖM��ތźE�޺���?L! d�$����j-�j:;�LO�lvN��������|�2K�U�Eս<*��C�],_��u}`�WْcGٞ�앷���c��{�̂hw������[O���x���1�J��*�I,Y�?y��~z���uC�:Go�＜7q������_�Jd}�����EG��3M���Ћn�O[�G�g"��Ϳ�/���;ݞ���׽��iY}.�]oM�"���ƓJ_������� ���D�E-Y.�C��N�l���e��W�8�׫�Fe�q��P#XDz�S��0����JXmq˄r���.u��bN�{F׳�]��H����b8�+`z�����U�K1�,��k��hʦS����&e;h5y�2�;$�l��5N۝�a.KnV^7lۣ�Rh�ȥ�q���ն{��͍>^�F�B�m�N�%Ŏ��~�������ky]e�>�����C+���sY�����A�Qm;s�q.�Y��>�d�#$�����g��b{�;��;��!��|��^,1�+�����_��(�w��l��V���+� ��d�_�>��������`�{΅�>!%Y�;]<ǖ�h�V�?y ���Y�%�?C���N��p��*>ݦ�������uG�� �(c�,%X �D?I3�dۏ^�y�J�cn�0A<~���AK��Y���VS�;;��<s�X#���x8&r�8����,X2J�A��~C�%���*�%{�;��Y���+c�g��>��������/���B2J���P��G=f9G5wr�VԡP7hd����5�jM�kPIu73B�Y���-^]�f\��׹x#��!�js�����i���[��������	z�jƱ��t8�>���)�A"��0�(
��(�9X2w��kzq�j7�z�f���z�yp�H_�-��y����Q�swXw����;:�t���}�4
��wʵ��,ly��m��*v�O��}����Ԃk�\���<ו�5��>@��*� ��zŃ���;��;��X��:��"s�������[�o"�g�=�T6C��{+��>�5�_��B��?I+I,X?D��7�n���&]��W����v/��K+#�=������2�h Q�Fy��j�y!���v�H x�$�`�$�`��+���^4�W8�X7io|�Fָּ���o�?NZ��=b����%��h��I���'���2��%�b���&��5;�r^����t�m�r�Ʊ�����W�4���2<�/�
�p���^�v]��F��;��˶��*� ��U�D�Ń�K�%Yz���%�c�����ȕ��sch�na���)���O�G,Y�T�9F/�(�G^P�'P�0�d�d����A������U֗�)�L�P�*�Շ�W%`ˮ�V��.2�R԰�=ƻ�����qWUy8t �6����-�V'w�}����˵Z�5z.��o���*���|D�ř%|����
��a1
���/풙�����We�m�Wz'綄�,z�Z���D���nX��� �I__�K���{y��u�����Q��5U�ׁ�4���%X �������|I5�_�<و���8�+�g:��_j��Mu�n-h��V*�/$�Ao�,L!%X �$�e�s�7�OV'�vw}~@�-�w7ʾ��[�_����1���9�2<�/�A���{]����{������l������	�#㙋+��0���#�|.�zU��Ń�A|D��W,��M���z�<�yj3���r�k�4��X�$�P"Iv�[^g�������VA�_�o��ފz�=㳻���_W(f�]=گw�w���#��T�؆YI��G�qU�{u�\��Hqu�����OQ�2��т�U�O5�%���\jZ�i��@�|���*?��s�18Ќ�9���U7����b`i�K�dw����[�};�m��O�FIW��%��[ϯ1Tz�\�E)DĨ�2J�~�\u��j�M�RXJQ�b`�̸$��V[����%��zuޖ/��_/����G5��X=�)UG99��1�G����ےŗ�V?
I/��(X!e�i^�붕�r����C~�`�ٗ�ҽZ��s�����*�=,Y�B*�7���r��s��u|�#��Ib�2J�"̼�!�Y��t��׳�ߥ�d]މ���'�:D�U�d��>C6�]���u�fx����2��`���$�b���륃ޒ�Ts����#�w���V泞�_>���xN($��d�,	��%S�ѹG~_G,Y���/gJ�����﬏�+���,_���J>˯e�ۢ��𾵧(Q�pu���*�X�9�n����?�n�Խ��nt$'��!T-Q�6M˦fk�W����*��b!
�4;�}������r�9������k`�Z�e��D���q�'Y���^`�#h���c
k�i �=K��8��0� w���yk,'�.�� �*m��l�j��T��W�# ��\ŗI�P,	[Rd���g)u��U�Bh��ۇOG�l� 8���+K��s�*Y��qN�uۀ�ҝ�1�����Q4+��hٵ���Wp���λ1֮���{c����ƚ�e�ńVf����d�v5�/M8���@�TQ)D�$)�+⪪���r$�b�#
��z��w�տKxȻ�'��TS)m�P����U�d�,�@�%X#�ؒ���������$�k��~V�{�R��rsk������}�G��w_'�=e��n��;�Z1�b�c�y���6�W���w�����<�w��	ƾ���g�_��n���wt���!���_lu����3пW���>�猋���BAD��9{NH�|�N��c7R������f3{�ϼ�׮�����({9�}v���Z��r�k��Ҿ �%
�W���tO�^��w��}m�&e�q�����7�]�j�q�<b��$i�,��k)30�,A�f �)��|Amس����gJ�3���aow�}�*���lFw��#9U{��� ����>���Ei��󱶸<��t�o
����/¦%9,z]i�6�e�FE5��NtqPD�[�C3�#�&<���]O� ��m�8���\w/m��.��dej�HI�#�wg6�z#73�s�j3�
�V����*;ݔ5̫ߔLWyz��7�>�ҩ����$iD(Qm��A3�v(d�ٕ��Z�z�|~��Emذw��+�ҫ��<�w�����0�7��?Z�� 3�TOv��w���H���w���>0A� $Y_Vn��{<��/��N"o����`�� [_Sn��5���CG��i{��bb�R��������p��rI�7t��
�Z�B�R߫@@���c��/�����mʟiܹ�^�j�ւ3W�B�Z�^*�pY�Q�_v�"�hM��w�B�$�\Ym�B4yQwu���}+���;�� ~8�}b�?>��q繜~��޲��=x�u���w��3��{'�ty��6��}E�7s���'�Q��+��,6ʕ&E���<�'�y.�o��G"]���UףK�SS.��q�ז�q���޼�e�+.�42�9⼻����Z��FUaeǔFlBĢ�W�f��v��^@�k���J-����o��#2K�`��Fi�R�^:t(�6jqz�rYv|jdHiP�'ճw���� ]�U��
]��=r�����Ϫ����'E�$r��	y.l����/y_+uC�sf�Q�*�\�H�Z�U,|�4��/��x�K����r�����L=wv��M�ʂޛx*�fՊ�����<wfA���y�DOCBI׶Wue$��T�K�:�wk.��T�vh�R]a��R.�n��x��-^��Yf�nUM��w-s��*Y���-�Go��ڽ]�Z{VZsFgV�Tw^q�;�ٝ5'�D������E^������I����X�&
�[�ia���˼"���M�t��[�q�^J4���0���:��Y�e�
��zU�Fg'ϯ@�:�=��Ԩ1W/ͥ�,k��O�k��Շ������e��7�hF��y0���źqUXR�âfm�w4s��y}�UQ�U��W���k��˵�֫r�:�e��J�t�.KH�ީE	;U^��im;mr�U��
,;:��Ƥ�1�P��\��̜�Wf��I��5n�]]���,�S�Ɩe�����={T��=�ku��Y�6)�{6�;rf��cʓ*T�ԕ���\�ʏ�ܙ�ܬ�5T:��-�t�6�5Y���n�kN�ֳ���}_5�ni�����8⸈�#��{��%ftu���{�ZW�qۢmYGRw@���Q@y�)Nr�."���%@��v�<Ԩ8'����A�絲���ݷc�꒓��8������ԖVv��r��J{u�đtE�Q�t"����^vDw'r��u�f'wOm$+���B���Ml;��mvwM�=++N$���N����Ã���ugYy�\^q��E^g��8����l�9�nq&�����9���
)8�H�a�^�j�ݐKm(�+�l۠�"�+��.̎�+����~[�������KUyl��;�BA� � Amذ~h �U�/5�xW�svŀ~���n�}�o<�U珣���{+��Q���P�li�*��݁@�ۡ`�!|[]�������+�݋3۝�[=+��s��a8���Y���AwC$�*g���ͤ�
��Uѻq͙ �>yħGV�mէ����ڣ�ܺth�9��Q�ͺ߈����g��\|D�Pcc�� ����!E@��?4 � C��k���,���P���s��r�Ҽ���	���@��}���痽42!@���~���F� ���+C��\9��-�.U�M����Q΅��_�
����0���{L~��(ޫ��C5�{͎�}z��&!�,2�4U5�}�&�0�\ӡ������Hܼ˷�f�䞞��=j�,�W=4�{��$GZy��e)�Us&s$,
��*KO������ͯ����%�D���*��؆��}m�z��ݾ��eS���HeD�(�XC9=V��#o�~8.�=n�'>�]UC;�uֺ��s�[��*��)x�U�X^U���lG]݆;f�X�w?d���+�;*�'x������;כ���_�
�VA!��7}B���5e�U�8��c����~>}��|D�P gP���"�#�'�C��,�}����?4�-�G�O,��9!���}^�ʧS�^ ����%
�VA2�!��]~�v�4����� ���/��K~ɚ����V�9��{�	ƨB��	������|D�(�Y�m
-�[����l.t��#7n��z�-����hH?2mW�6�;�ަ�*���z�Y<�+��o7�F��2/>���>���w�0�K&�����J��Q�u{�hw��k"�3;䢅>�92��>}�5z�*���te�b7>�vMp���[��  B���B��ݐ��N��V�ru��N���L�kq��ɞK:�]Kj�nh�gj4 ��''A݂� I�an�(�R��j�F�,f(B�����x.�9�9M������W�g�e����� �lghxx6�f�OpɍC	��y���5�>x"n����ɓ4�,��߿����~�Z��)O��|��O䵛��t�惢��v��j��\���
�њ���n���1����y5��a^[WX�V˘n|�e?DM}e�9�Ȇډ��c���L�ݏ�5w��no���TA��Ń��ٚ�u�\��s����P �;�7^�E��ãE�Yx�m�� �.���o�C*Q�������\��<�񽜄�
�%���j�-�~h/힮�=��孬 �俄?ct(w7�w�/8ʧS�^�e�1�zz��5��~��"�hM�w��c���i��ކ������bt���~�������;�� �����~i|[����{��z��৕�d�h+��	
Ud�于rɈ �։�F[CT�L��<�3��Ϟ��[=����6�=�Lw��N�ogK�Η��8����^���ܾm�m|���\j����m/�2�W��I��Z��
���w]̩�O0^�,�Á/�p߳l8j]��>Y�vCϻmt�@�Y��r�꿀}����ހ5��̇G!�Y�yn�4]����>����9	�n�|�v>m����x�=�~�/�-�s�<5���ͦ�{�ޗi�}��C(x����=����c'tlt������++�{3���f7Z��.�]ڻ�[�ۤ�G�W��y=ǻ�W�S��g�m}"����+r� �۔�戈Q��H(3Bpdlƹ��\��Ij���f:��]qt.޷�~�3��{�sn�~�=��/��"��;��>�:}:�����}�6�m�m�IyA�/�g�:��[�,v���޽�/�|������۽�*�}>�_6�6����iu�}�w���gk��$�g���9{s���pJ��.�Zw���*��KS59pʃ6�/:��F�}aI��|>}W�a��6UnJ�Vw͡"m���������/y��m�ޞ׹6�]�v-�s�=���{2�w��j�& =ͼ��͠�n��wT�{Sk���X����sz�t��n���h6��sڳ�M�V��J�$��tQ���J1��[b�7�����F�'q�۳�6��~?��!�t�_6�}����5��ӹ;vxNU�+�ڟ���ޯ�n�m���߂�4>:��~��y�m���b��;��c@>tl=ih�ϻ�[��{��m��m�m�����%v#�;���ͷ���z��6�m�hO=)�k�a��O�͡��$�S³�&�N͞E��v'w}.5�욜�U?x�E:U���Ҵ��L=1�/o̔��|�ڬ�/kEU/J�	��J��v���q�}�G~A�j�T���u������qw%N�G���ju0�kf��lΧ�S����5����5��W�U�ߏ�� �xKf���J�p\�ݱo[F6ˠV�BݠB�؁4b�,�*������ͷ��yȱ��8'���:V�����
Z;��6��@6�o-z�Q���D���y;D����tE����~�DۼF��4j��~������6�k�޲�*o��~�s���*�����cA�o m�����_����䇳σhc���?y�=��Ҽ=n����Q�[R�v����]�m�ܶ�&�v�B^��9OY�Dә;_zE�6���{�H�W��ex�����Xֵv�S�7�l�]����7>�����^.p�K�t�j��fV1�T��j�n(�yWm�y/<^g������`z��\Q�I��#x�ղ���q*��
�%�7���ɲ��Nf���ګ��X���0�V4��tu�p��6�2�e�<�g6����:"u��8N^+��@x���Y���� 3̗8��5l\�Kz�rkZҦJ�(\�p��������3Ⱦ1�ӭ[�Ĳ2��么��5�=�i-�j�.�E֫j�:u[��,�o�>e����1��I��Ofz�;[P�V*�a.�#j�x㫣k�sg~����ۋ���پw1K1�j~J�6�~5C���e�r�k��C��n�m[g~�h��B�}{�>ֱ��c��lݘ�Ε�r�������ۼϣA믛@63$��5��Y���g9w��Ml����E�|ۯ�M������¯_������� t;��b�c��kʝ6�G�^ڱ`�[�i�_�m|����My?S�Dh���>�΂{���xz� �|_6�Cy�,��%U�y U
FB�Ф����<�h[Jy2�ۘ�0n�f�Bb@��V%V[�}������M��v�3�u�ߔgfN����˻���!��#th6�m�)%Z0�gA�^��{Y8*h���OШTR^��J��W�G��;������n��T�{GO/j��3������>�]�7we�ǣ{��z)�n�돾����3�l{<��������|�����+sF�9��^;���ޙA�m�6���z����ܿ��A�[��o���3Nޞixn��!&�k�XҾ����M���|��p௦��ɞ\�����V'���ﱠ�Pm7��좖Yt��ff��:� ����-������C�D�"`�����&߾w~�w��{���o�d���C�x�N���<��7�`�߆o��t������y��M;�5�c�3��-��sk_oO	��"mҞ�u�gJl�E����P��_6��`��#;���$��ٽ6�F�v/wz�pKN����u;!�V���Vs�_�YC7�k����N����w�_M�́����j��X߶����6�p.����ۡ�k�5�U���}�7�ld�����X�N��2���&�q�������6mP����~�}��>����j璵������"m��������4��	UJ.ԕ�r��\p�팃�Ƭ�w���x�{!��n������u�{9��;���>����gN�`��}�|���_6��MT�sR�Y�7���'���'r�rw/��|�yJ�X��>�t9����z�σ}��S�/`�u���2�j�Z�_xw/�M���~ڢF-��{���C|���&�}�f�S�g�,O������Ҭܵ���f�UOtn�sƲ��e����Ʀ��%�N�@��+-n�Il��O��i���z�r�U�ɫڂ��IA+�6�~ �7��^�6�������1�(E��O�O����X�N�S�h6��o�_v�[��ܺ�T
6�M���[FUwcny�'gq69�0�Ǜ�sdٻ�O�/���_6�ޏ{�ǩ��[�������[��;Zޠ�vۢ�$�pƕԛ�}������������=��G������^�|����m��­���;{r�p�on�����^�+�����S��:<�˞҆���y]�����u���ڬ~o@o��&�VEpe����+�i�۠M�{85~�ȷ`��'����nwl�Ŋvwv��of6�s�[z,#���Z)�n=��f��)��[�"�_㷁-�l�9.�ح�#��W���Ƴ��0�(mk���C6����rf�yl���rP�uX�SӶ���c��,�*�w����-!2���Ff,�9�ݼ�;A���N�/��l��:���܆�ĺ���Y}dq�洍�3rh����f�K���
b0�r��}|:��*�4����%+�+����W���:�J��,��n�<�q�6ݞ}p��y�@��L@�-��j�Sw*<��]R�fL@�96�*V���g��&����C��ve����'�Z�}�h-y�5�k�3�>D�{1�/z�g@����m�3.n�HѻB�n� �B�y���x�+�F4��#"ne��Ğ췌�Hu����f�4똊4공[X�Q���$��*غ�f5���7��j��I1�s���j�sr��Y�u�;SP�K�v�g<��7+��:v�2*uNC���o.�>�H�2n��,�����ի�٥xťU�����iP#wVS��=P���9��2��VEɵ��;噦�"���7�u��ʷ'Jg6/���֝��]W�l�X�*����f��9�nd�ٔ*�v��,<�k��y���Ȍ���
�S��vk��r/+��7+�s��&�+.���#�Ow٦b};*n��Rҭ�*n"�r���ᶥ��ݺWf�&()�%aqw�<�c/�銍��ʺ��!Ō�bTQ��V���3��;4Ք^0鍊�wZ`�u�^gz�L�$�\�n0���o�ǂvq�4�2�b�J��)�z[�؅e9	��6!
�,��=�����.����+/����)q�v_;�"����n��[�2����vA����}�-y��Qvu������ǙQ�����Yם�E|���Ս��⎤�0Σ���/;:�:�+�Y�v�f\dG}��u��i�����u9Q������r^U������DP�����}�>��9�T�֝$�Eyw����ݐ]���Gq��Ug^|�����+��l訳����r;��:2�=����}���k#{��쫸u��)�[�G��]�N:����p��Me����ڇ��z��������U�@�`�8�n[��5��K�<wDb#v�g�S�zP��6�u�.���n)�3Y�e(愪��maR�M���ix͹�h���� 7ir$��[Ep���hk�۳q�igڃ�d<9�¼���GfÉ�[y%���A4RД9��g9�`�Vݭ1��):�gs�\��E�݆�u�-��fa�a��/�Lm#-KE�3�x�R[P���䜸�6��4	�բ�Jq.�627[�^X����a�7R'm8g�k����Cr�%���bv��E��y���w݈�]�편M�۫�ܭj�kEL�K��B�1tۋ�h�jM��8�r�y�2�$H����X���+U���X�E�D���8=���V�l���b��6�$�jk)���ݎ����n��u�5�Y�=X�nw`�^�l<��W^���͹�M6J]&mOU�l����s�Ln�gf�v�a��q�G}��*I]�v��{M��zh���nt�x�в�:1���t#An��u�p\xq��V�qd��4[Y�;=�{pM�6�Y#d�uO�w\5���m�������&aeå^���02��BĩJ��6%������z��<mk�`��:e��WvA�@4��d�z׏%�i2���m6�K��[�1�͔ XYb�$�g��k�®f�'5\&�[�N{/���G:��pB�{T������}�=�9�s���[���%���9���0Kn%�Ř�qc�qp���ZCw[Wř�-I�y�m��i��J��,"�$76m/PT���Y��Ve&��h��HѸ\ٖ'�9�p�c5ӱv�2;ny*I�������ĕ����4��]f�4����+�2���.;C��[�{�k�8�h���n���2��M�k����<ᗒ��=�\�ݩ�B��F������4�kv8��6ڸ�e����]�N&���wui/�X)r������F،��K(]�4�n�`�ˍ5!�طli,HU iT�+FR&��v���ٞŮN�9tHi�8�l���W��+�7��\�H��V]�t��t��,���`�9K��L�kJ0�n��K�S� �ʖ/:�Z����ii�j�e{ �l�#˳�p�:�[�Z�L��x.�A�:�>Ѭ�;p�E|�?��#�T����H�l�Mo�qֶ��&��\وH+�]U�e]�Y/����m�m�9�����ʼ��S����������|tA�$��Uc(���=�;q�{�yW�޽����'�� �bǝ�+�:6���ޝ_|�vo�2wke��\�vt���6��=�M��t$����ޞ*�?J��Ǚ=�f����ܽ���Ҽg���կ��+��ͯ�m�e�y�-Q�`]=/-�h�暬~o@�C�y�m�-z裊R=eU]/��vf�X�T��Q��fA�6�k�F�q���WѦ���;�E��)�:m�{&e�����m|ۯ�@>ɋ���|}pf��	���L��B�M����ܨ*�S����X��`��Q�;ɵ�[�;w)ULGQ��^�qw��j�v�۱�X�'�}V/t���m�}9|�].�s��w�z��w ۠��ȕ��NN��z��ξ�ܾ���۹]L�y_�߭"[���ۡ�����b�;'M�����!���{�y��6�ͦ����]��e��h�&{٬?x�w/<�ɵ�m���~�B����S�+(��V/꺥B�W�#��R�<�3��-��&�f��.�B�LŪ�M/�s�}���wU�����
s������ݚ�3g��x���y{]|�m|ۡ�h�omdZ/������u�Ov,S�t�=Oe7j�4���)2��m�[
�m�y��n�ě��R�q"놺�ĝXt���Mh�،��z�Q8��h���Q�n�uG��m����s��b�vESQU��(��h{��~�x�����y�|'/�_6�Ͻ^}�U>��K�������瑷�4n
s���ߛ��b���W�s�r���k��������A�ӻ��L�����Oq�3�t�}�����k�^��9�H�R����F�T]�ܠy��&��]�S��-�n��k��1���ڃ��_7����z����܏�xwzR����<��f0��y ۠�������AM"v��:�!ױ��xh��1V7�>_H�|so6�hxkM�t�:m|�m�]����d���;�ɮ�;�a����hr�@6�n������y �Oަ�{�+	ݝ��̶�@��R��eM"��ܨ�*Jv2��$G�!�u��#Db������955w���Ifo��<���Y|�g_,�9֏>�-泓GZ�Gw3b��Z��%�~���پ�����A�����oK�|�MlOL�:䭝�=�t�t��쮼Z���.�ۡ��}96�f��\��V�� �� BcJn,RƸ,��F��a_��+�{��&���]��Eݙ�����o�ߑI��D���B��m��7���1	�����_	噣|Ol�ح�}�l�����������mK��P�۠�}NeIc��V����\rV����|�����n���P��ߧN�r��I=�p���|�OG�eޯy��6�6�ͯ�g����-�A͚�5�O�-��V�����ϝ���LS܈��u��N��a��-��n��5Ү�!]|l�I�uf�ݷ�%ej��k�H:��ZԙտE)�p�ʝ��\�W���%h����zY"�8�ۇ��BQюp���I� \����]�#՛xG�]]uu��;˻V�ڱ��uO݁=����N��֚0�C]K4#I.8ӊ�=�;�q�+��ŮZ���`���2M_l��c�z��;��}��-wQ[,I��6'\ڗ���
Yl�$pJ�u�Wf��N.(%�u��6�ݤ�:����]������M�I2�4%�v�'�gr������R��l�0��%F.��}u����f�y�5`w%l����^�R.΂߻q�����6�_6�Ӌ�w�����Wl��gI�ۇ��M��C���o�o���}�T��{C�|���A��v/��=2���������G�;��$M��t#39������2�&׶s/���8ܗ��'�r�$��?K{�;�͠u�mә�K��,�^�/6�w7<;t�\�����(�l�뮓p{�j���	��7�[AB�q��q�M���7O���!F7n��²��/u�����n�mc���������/v�M=��1�$�^�7Sh�|���ih���Jg�%ߊ�ώr�u����h�N�7F� /E�ön�Q؝��S�7p2���u��c"�R��j_+9N�=�w7sU?�~�| Y߀q��ݳ��~��jK�ݏ���"����� ~���>ޔ�vo�5:V��a���~~np�OWN��ۨ}�Sh�ͺϝ�+7�S�+'���.�tkIݚ��H����q�~�����X�Pm��6��SU��CӞuj����c�|�Z��wc��C�x n���ߑC�>��	ߝ5��mjn�6���I�<ڙ��U���u�/gzM���4�?����m����6gw7<#��ӻ|��vy��=����5�Ͷ���_�{�}��{��9Бc6#�f？�䏹x���7�e7y�^u'�V��@6�|���ePPn��*�M:�K�A+�y=���r�wl��y�����ٶ��&��C.���xL��a9�I�Z��AQu�.#��}������}:�w����_H�u�m��8��a���ݠ'5��6�z�]��o�Q1z�h����_o&�}�h6�o�w����'2������q�/�W�ɴd���ס+�D�QP&�4"1]�𯒌
'���m��<��p�oN�w�0k��j�*������ok�s�;��j;�ݍ�JB��|/�;��ͯ�w��^���yX��M+տ}Ӫ�{e�N��1��ϻ|7W��o�:�:�4~m�C�7���ފ�Ot���9p��#U�oJ~��>���eܛM�����DS�b��>�ձ|���=>�y_u��>�~�6�`Q�_�x�޳b���x��/*�&��4z� ��wp�s	�r���mnwkb�+����TiU>E��mgӛ��۫�|���U��#2_,F�P9C���g�f����t�o���p+B�_\��=��*{��s��=@c�.��u��$]�(e�B4G�`$�a�����q�LY5\��k��[�d���Џ;CV�� �|��m�k��<Ͻ��^~G}�}^�\�.X�4��6�6�m�Q����6����O�<W�u�wv�}܃��w��od�F�m��z�m�ͱ;V粗��of{ީ��]ϻ|>z����m�����40�;��|�<'�{�ۇn�[q�V�4z�L?3XvKƠ��5��_6�n�o}y(﮽r��T������{'a�q�s�q��س�k7'h�Ī��U{�,�Kͫ��y���U�]zˁ�a�vj����oԱ�7mR�+6�nU���aڙ}I�;�vОxeTeK��܈@0�!1*ۓ �#���9�%��i9�Z�ٳE��2���c��2���&�Պw6RWC �6Y�#m�z��M�&gy��8�G֎}�������/y|k7۾�~�6��B�ֺ9�g;��#J��'N.�d��k�Q�(�V�+�,+���\��a�t���s=Ci�ݵG/ض�z�yL���\Ma+��|�?�����5����.. 2��s�Ս�3�kcc� �1�.ma��oo��s���m ۡo�w3��xs�s��S�l��Q*W���I�7������Wy�n�s���=3/e��o���w/|7�@w7�
�x��w�{O�=]�y��o2�F�a/пn�{O.��v�}��E�6�|M�V7�v:��gދy|۫}ճ;���<aN}����C�b�� ����m���!��j�١����t�w.��^�J�Eܽ���܃k��O�����_*���F��URJ���H3��qf:\��`�^h�Ηd�lG��=>����W͠C����w�{�e9;��e���m�o�x��=�精��ͺAE{����u�����s��[#%�^�z]�7��l\�=�W�p5��;U0]����Lʦ�L��7h���v$B����t�T��.q�ٺ��|�=�����2��o��_c��v]eg�{.`Y�=:��փn�os���2y},����9��Uq�=��@�>m6��K9ڽ~�{�_tM��?>���{�*����tOH��ӝ�����C�w�m��6��O9�[�b�����r���T��%s���P�������ھ���|�ou|u�:`ܗB�=�Ym�5�l8�C�SB��i�Jh.�:T��|�����o>��0w��P���U1�=�{;��>S����m�ͦ�,��=������@s_c��:�?��T��{��	l���j֊�|�ʱ���(6����~���=����'r�4���E���z�d��Ka[�#���uP�ʯ%��x8/��B�D/3_U/$�Rh;�:�qm�y�]̮\�CB�:�v�ɉe�*���J�XW�6U��t�K�`D��J����5ȝJ��}i[�̙w�}T�͹�܍�l��fk��t.����s�H�ZLD4��F����5�ʥ�v�
���%�B妔ն�S3#������X=��rk+u��tҪQ�e&e�rzF�|�H��۞~']
>��a$|�[Pf_��Pm��̲�t�;�l�o��U��J
X-d�4ҷ�˔W3M^5h��-h�QWUU�L�,�jAa�Jv@ȡ}�����-nV�;�0kk�,�X��9��J����>����׻[��	)o3L:!k�t�\�{:婰�XKѼ�"6�n��D���[���-n[����ʯ���!��F��en}*M�7��7�)6j��{T�.uYz���T[ذ`w��p�Օ�.bǖ�[a��;�UeLV�ok�U��/�7���q�qT3QwjR��ae�[�JZ�j���i8�c��]��w�ڭI�ɦ�[�g�՝��fYe��lGe����Z��,��)����a�7���HO�K���w�*�Wk����ۘ��^eS�������2V�����c]��XI#�	�RD�u��f��hLVǓ+��5f����՛�=Q�;ZOW+�t\���t乤i�<skf��7O�қ����*6�*�C�qK������ڶZ�L�U֊Q\���f�; �q3�t0���l�l�&��*t��O�@���.�i+^�ͮˈR�h-��Z�Aa���y�u��sh��.��^����+��Pu�I�gǵw�[d:f�������^^W�^���g^X\u�o�{����3�<�.^����n�I�5���m�5��RKK�Bem�&*�k�7^)zk҇4�!d�8�k'h��al��m\�=��Ϝ�,�;}��;{���ޙ��\������7�������vwf�g_+������n�����]�|����̢���cJ�V^>���O����_��^�1����f�];���@c��ͦ��j�ے�Ӓ�m}�0{��P���U1�=��T��n����?z�C��m�lD�9Zڻ������k�=�m����t@H�m����:�J�J󼿬Q�$�J]R���ݛd�r��;�\���F�ٲ��f�O1Ѝ��6���'vߺ-�/�v�`K�|�,��8�W�|�m���T|��w\��!�2UO��jU1�=��(w ��y��j���z����m��tϫ�9U^��=샞��w=����A����g�{�{ƺ]+U`=C�|�{���������f��y���1dUr���w��.ҡ6������U�e�ܷ{���^�9-��I��Iw,zO�P��]|�4�*����d�SUW�|���{�_6�m�a�����}�?A*��<��*�3Ǽ7�S���ny��e�B���[�C�Zk.V�*����E��O.2F�A�^�6#N�m�"H$@��E$	���p7m]��q��|����=�7$�y�f�W��|+�v�m|��Ώ*������x��h��������u{��};�٨|���+�F�w<���۠�џ{3x�������Y�7�iT�=�7�S�h�|�pVY�7mMɔ� 6������d���'t�}�����H�� ��ѻ����~9���wr��; �M���M�N�wo�jWͦ�<�+�qg��9��[.�U͏�K\�g�[wݵ�6;���ē�n��
������Z{��, �)z����d[�c��}�3��	l]�m����X��`��w/�X�v3��6z�c�rF���q�Rp���t���dL��r�MŲ-�c�c��sr$�ي��0cc@���(99��Е��]�y���l���	�:p����i�����pn�G'K��Ņ�E��]�u�`��uU��#��d�(�L�� ;"@�k�5a�g��!Cj��:�ٷ<Aū��g��Oű�A�ʙ*%ꥮݧ�V��ِ�U�cGOeB�hQ�5f�������_6��ќWT���������N�~��{�x���OSiN�7;�>~���L{ܓ�g��&�mxT=Fv+�����>ȳ�]����ܭ�V}��koڵk��&��o�5������N�T�&��_ً�}C��ٸ|W�x����������1{���=Cu�k�������[u�}�&�zwyzi�c;�wL��D۠���/�>{��{S��.��\�	kKl�k)l`͋	6���n�,����)X(��J�7K��率��n�=/�:����[�;��|���wJ˕���h6�6�Z:�o�\�W����=cFg�r���9DaD���'jbT���x'Hӡ�+'L��_��ƻ�Ӭ�wyU9���3*_[��]%���#�W�fa�����/�G��Lr�!�mW�8^�[�1��Vh��^�什�����m�m7���yCm/M���.�[p=�;�{����_]�2wDlM���{�5�v��ܖ�׏�s���f �U\�6{r/��x>m�ח���U�r����R��g��ޞ�u1�{��P��_|��=J�îЏܪ�B�$j�HY��-PY�.��GX���!4��SWL#-ؔS��??�ߢ{�����=�<}�o`��w\�ݞ���"j������J���h6�\[�Y�v����=����[����~����Z���_ݩ�_��m��D����/R���j��m�����UX���ż�ڑ�{r�}k1Y�5ieB�� �b�9��wep��.��y��J��(��0c���j͖��7sh��Y��
�_cM��o�jW��O���y|_	;zx���o ��w\�� kp��T�Fټܯ�_6���6�����eƱy�_�{zϻ���=�;����gsxQ/^y�ׯ�'���5�@��"J8,�e7C0�\c0"]�X��kFW;mc���O_���߿~�n���}ޞr�{Õ�1�	�Pl_lA�A�T�^v���L_F�����{|�yܓ���!􍶅z�O��=�_���hߣ(j��~Ｂ��y��{��q=y;����;���m���CQM�m?��֡wz�#T-a���>��߆_�b'��h��]a]�z+9^�Z,D���gJ�PC��qjcr��ًk,��U�է&��չ�jˎ:6���X6�0�v9���C?����G��6��o߂���'���?r�o�אM�;�xH��|��oݺ��h�ۘ�����eu�@�GN�MK8�`��wm�Z):�"��6R�l�տf:����k�ƻ�OTǊk�������N����OW��6�n�mSiK\r��ܳs˩W�}�ί�,������}w��I�I���f~��� �z�>mc�V�������v����N�)n���%'��A�{��DmH���*z�<Q����^%$W�Ҭ����Y��>@	�6��m���H|�ëJ�ڭ؝S��zx>����}���6�m��,��g�������ă�/��7.�K���������ɶ:�{/Ǆ�䐍�{6�O�����;��}wV����W��w<�C	)]rK1�ڗo��.�kN$T.lָ�3&
4�Kei5K-U�6�]���v�kh��qN"ɻ.���9�8l��7.��e���)u�P��A�H�2�LŉŮ4�
ɺl�W0�g�7X���ƕ�jџ3Ҋ�=��������[��M���Q�8t���6��V�˛��b*�7f�tnMS6rݽ��"l�E�-ζ'��W���[�O��j���ؙeik�O.�;#��X7F8�۠�$J$���:�wp۫���o��p������3��!�4ױ�O|�M��	�91wZ����y��WG���w�=��������}m9ܻ�K7+���ͺ��z+'��
�t���������=����t�[v�����m����mOv����/^�	n>��D8������΀�A�n���2S�lgX���z���)��N��^/����l����M'��/�*J��V�2�T�k,S�n��n�b]3��e������ ۯ�C7|���㾞���3&���CҬ+�z��ͺ����{��1�~�U�>2��v�O���]�xpt�P�g#���DWS��WF�;�&�=V��*
��������k��\��C��k���{�e���{��F��{k��x��y ܯ�n�m�����m�X+jSy���tw�v=���Ҿm|���b������ ��u�X4���y5��߇�Tc���M�ϳR� '�����d_��{�{YV-� <�e���d{�����[��~n �������kK��=~	��ݑuh�:�f����v)��16�یS�� � ���?B��ǊH!����fd��u��^����sT{;�5��3]ly)��z�6�ĀFfL����_tЏLs{u}?n����䰺;3�����C�ƽ�H?f�����o�y��i��+���A./�IH�L���2_�ϩ��i��]x;��m��ɢ8�N���Z���vj���7��Q��N�P#�q��d�gv�u݁![�v�W�ۛ�|�O�eݵ��wۆ�$y�S鬷�m_� �[��7fb��Df �����V�f^�>�LN�T���W�<K㙒&[��{{.k�u���	�B��Gr�����OE�v���@��'���3#��\��1ѝ��ac���'����P߫��&��~ 栈�K�fH�_��s�3��z������k�qY����3mrlmY�<��ț��
�� �VU.��{ǹ{籖_��7|�Q�B�zw�G����Me�V��Ȼ��؞��,}ւ7��sDf/��3��~�����m��6��{G����߹��������D���\�����TGs��B� �_I+@ �(Ow�6��yj���T+2�VFg:��X_|� ׹O���#1/��"Nd"'�=�ǩ�tp �9��P �s!v��ol�wU1���|6�����Oj�(���R��6�x��'K����[5a���ʥ',�4�8,=af�W}[�$g-)��;�,o����->����0.|8-�U�:�彆�5�����V2P�� Nf)������Ŋ7�Ә=���	�?O�����v\Ϩe�>ˎ ���BShĪ �+�JY犺U�BB#���<�m<m����d��l�Izz�:���;5]�j�^o�� ��$� �%���}�tvo��az#8 ��X$�cٜ��.P�'/�Ib̋�2* �����p���Y�$�� �������9Ȝ�z6����~m}����E<;�G%�( Ej_c� ~�A3_̑��k���g��/ݛ�/3D{;�k���TA9��f �غpi�{� h�A�RA�AU�vK��Gb�-����&��Hݓ�b��|�n�ّD�s2D�ȼ��6�z��u����
�u������˷�i�w /�!�3�s�����K���:�`b��ݕ�鎙�N�Zjڠ�pס�e;���3���7IV�tV݋$pa�.��̻�]>:�ɪ��a��Ӻ���ʣ�bxm���L�+i7�N<�d��7Y�{U_P⭅B�<R�Nl�rV匲��Qs����m���]ׄ����6�#V[��=xb���-�tx#3�7&���b��ά�"WS+rf!��Qݫ&�Ι�ϒ�*㳦�v�^On��h��mI3ZZROz�.�c�wj(Óu2+��R�3)BmKdu햔4s��cT���<��f�V��n��B���[���c�Ź�F�f�\�ynF�ܡ:c#�_�w���$����uU�[��:�ie�.�����W��*��6�H��v1VB�7y��\�z�l�`�{J�ޗ;1鋋�c�̝7���>�ǻs5eU%Y�m���^���jP���aKk2J�|��+����x��F�ì�ˢ2�-}�(+�EW��b���A�JV�Xs�eowf�ʛ�f����"�l�1��ku�W2����������Y;n#V�ul�p]Kf��.t�1�M�riz�Q�
��03�oZ�Y6���UfYݾ���,�Ys3�geJ�v�#��bY������qN�բf=��X��M7p�::
�j�����fn�MŧY��V�}���ʐ�h��N�*��uV&���Y���Ru�%���ۼb�j�AJ�:�;��br��:�\ۨ~�e��M��f�Vnmgc�{ΙÿR19R�e�ݶX�Ji�c�/ĳ������w��1'cax�e�:�f��C^�/���-��:k�6F��ry|���n�̭�y��ڂ�����;���g�]en��^r��$:��V��#jǵM��`�';���׶:���m�Pvt�����׵y�M��]��zYԇ.��r��8��[��5�.��*=#٨�.�ΐ{�wg$�i�e����,�;�XW���;��׽���oj���)*:�9̸�'�����{o�^�On��/>^��<��l���Bx<T����n�gܷza��3:O�bw��>[o}��[,�}��-�V�cü�w��Y|ʕ��dMy��n
됻5��m85W2�9�<[�拭<vZ�����LG�l񧉴�{@[�Ws@�W7��M]��Mc�K4���s�G.�^ �
���A��z�m�{�厣��������d����b[�s��3fɳ�Պ�
���]����mq�hc��NU�n-�ͯWs������a{m�Ļe�������[]@��wN�Xk]�u�6ew+�&�lc�\-ۆ�c�:�3���td9��K�tƎ+�+V�g�$�� A'e�B;���;Ϭ*��ok�wgl	����KD�3�n&�*0l+�f�u�s��.ƞyS��ؔf���fˉb��"D��BQ�C���l���w@�<��ꍣ���h�w1]G3!s�b�!]���:/Dus�v���6g�z��i�s#�gc�w0cQ�jM��2�"SKKs��р[��D���Kmtl��h}�3C�Ssv�=���Yǉ��8��v��<ݎF��(�6�qmq�Pi6��76�����F ��`W�K��n1��\��L��g��[�wH���ea/-c��hX��6.q	Z�c�R0[Sf�ҧ0��	�Gsu,�;�kv�#�����oi��4XJūv.S"Z�{u��k����]�ݶd:މ�]�r4aL�9���5c��N��Ξ��;rp�n"I�8&�4�w�W�9�۶�vg3���G	��x��mC
.֠:9���J\n��x�ֻW����৭�U�Y����}�.�&覝kI�����01�5�]csŕ<㳩�+S1�ۈV�5ؖn6o\�;��m��b���ƀJ�@�m�P�{<�NolR����nȺd����Nt�pI��j�{W[c��ݺ�+G�kK�h�#�f�[�ݹ��/R��G��[��Z�lb0�V����Λ/Z1֒�]����I�)�f�]��C�����bwSX�ե�^�O&��++��>1��:�tc)��@ː
-��īD��0����!Lspq���!�^wWGP&�5�wnv�j�JZ.���z��[ؐA�q�WU��E_]|WU�=�5���tF0�bYݬn�C��vP�u�17��8磄�1�\:�&�9N/Y	�r��ɖ��lf�`�P�3F�"�,i{YXZ��/f���Q�g2�W�\�<��R��pl��{������U܊��糦��qc�zi�)�.�z�C$Gz��A�]���iڟ�����fd�������Y�P��=���s�p���w�y�/��������&��"ٻ��V�9�\��<_f��m�����-����8�) �3'֜N&6������'�QIb��P �1��1�~~����:kا.���� &�_�RA�"3 Xޏf���D��1+@ ��"�}$��Ͻ�����c�w��߁�_gcߺ�B��|y�=|D��"2W٘���'3���:�<����Ob��X_�� ~5�R���3���͜�ˎ���F�U�Wb�4
7a]��da�6�v�ЌV�Ԛ�^`�1BXCL�*Ks���e�	o�H9�� ��ݫӱ�v�9Ȝ�z6�n��3"�v�������2��R���s=�zE"|���R�7o��u���/{��r�
pך\�m������r��]@ڬL��Ι�����f���ù@����uy���}A}{�H���kڮ9����c���>�DO$H9������&%�SV�~�� � �b�A�t���G-��7�V.k�؛�~�_��kܾ��Fd|���s!���d9�B ��D��@�s!ڽ;�wT<�MݾZ�ۀ:g���M�ƅ}w�/�OGV���(d�`�%
���`uI�>����"f��-{�����U�]�����<� �B?fD��/�M�՛��/��[F�*�ҳ,U���$�su*h�c嚌�CA0܇��}}�[����� s1}���|�|���\�%�/�_#��dsBx_�E����������̟�"�'2!�M���>>�D�	�^��绪z&������ M��9��}lb��^�؂"� N�����#1�f!�O��;�F/��sR�&�ʋ3j'=���9PKP���;�ޡ},!��d�Ӽ���+��{4���X��W�5bꍸ���<���t7˷9ug{}sټ�̃]������@�7��E_A�P"LAH�锶�eoow�d ��?�U��_*��3�Bt��� M����5��u������V�ӡ|w:D�s!	�W��$�,ȹn��-h��ʃ��}�wT<�MݾZ�������$��Y�Z�%��n�z�DB�������vj���c�����X�h��v�5H3u��V �.ڒ�����3$H���e﫣'=��q��}~��D�lw��(���R���ŗ�K	��_�N�M�T��{T�����+�Q��[/�_/�ܤ~ƀ�4�/7����0����բ?�V�9�0yʸ��V;Ɔì�\s �*�G��O=-���`��
 ��(�*�"D�=�g�3l�F�(��b��/�fHT޽�:�99��w�_� ��_���ez_�/�zM����w��$�x��Hg���,M���O�w�}�%��u�C�6���o`��[��[����9�� ��D���  Fdf)����_]c��Mu
�u-��/�ߵO�����34��'����<w�he�LV��y�x�"�ݗ�`P�:�]�n�6�#v��f��{���{�"Nd '2���Ø��O=1���"��A�~��T�N���__�P�D��L���q���똺{����� m��k/�]o���=��q��p?z�H�s#3�{C#*�1@��A�B�!@%X����5~̜��Cf����K-��/� �}8�@�PKdU����}B/Ƀ���x��u"A��ِ�޻�:�v��1���� B�Վ
��bA����A|̀�f)��b�Ɋ�q7hN����"so��o���=��q��qT/�"�H�s! A9�F�r��C���-��>�KK�M�~;2�i��cow��Pg�9tN1�����@�s#ǟ��f�Bm��.���=�Sh����)�?@)�R��+#қ�r�-����v�+D�=�n�3�����]�'����-��W��-���q����F��s��͆�5��!��Xј�eݰ��ça�#�"R�-�/�f�qq�	�6{mF>�m���V�-��ک��X�<Kqc"�X�kj��q����W�o<^l�s�F�\Ŝbj�����7�5� �7M�v����=|�TN�/ҝ�;W� ��㬙$��]�^�#�4�Bmnf�Zֈ�s�����A�_H�B��yhu��t��/D_ �d[��������!_<��P�dT&E�8�g����?�D���8�wq���1�����C��f"���q=3�:k�P$8�@���������32DXс�������=[9�����'��7��Ȩ��PI(F��Wi�x����G�ڠA�!W��6�����Ͳ�E�@��� "d�Yɍ�QB�t	�}����b̊� Ȩ$�`Ȳ��b�E7�Lg�[G]�e���y�kz~쀀 �A�RA�B�C��]!s��L�?b���J9�t��N=WX���������'GtfUV)��7~�����=�,Nrˏ$�^l������fd2w���N�.���x�p �ݿ���2/��,"��F5l�z������y�짃�=^�]����v#��U����k.e-n�ޑa]��q;r�wF~�޲��\��
5b���*�<.j�V3�����������tn�Oge��e����Z�m���w��B�?oz*���,~� �/��D%�"�	�W�ߧ�{�0	s:o=>S��2��f<ᵽ ��~x�3�Fd��1��}Я���Z���g¾?	%��gw��f�[/ ٓ�F��U�"}������	~TD�łd@T�(%�!�>�g��o�P����l!}]��e����{W��3���X�`���o��.��H`Ud+�vI�E5��_4��|au�lЌ�Bk4������T�l~����B �~�?�@����'W��+��y�}���\:���+e��@� �7�O�f@@��'3�?�9R&|���c�'R�m����V/>U9�5��F��U|A�ŀd]`�;J�f����Z���P�"�J�IZAP��^x7V�\���F�(ɱ.�.����ǽeg+f�N5ND����ȼ��r�gl�֫Z�3;��9U�&J���1Wr��[d,�:�*ftx�8��?��g)�_�fbs#��͙�f�2�q��ڑ �B���	�n�S�{�1^�c���$�降�s���>�RA���|��}$� �@H?x��s#b���<o{�?N�)��V��\}��y����ȏa����x��
6i+$$б��F �3\L�F��&3��Zb���Y�C�݃���!Ʋ#\}���9�/_Xޜ�r;��s�s�_ �Mݘ�q����<V#{�����ľ9�"~9��'2>��:ΎP/��/a��=[�Թ�Y�o-�z�[Z��8ug.�Oգ�KA|Gt|�����3�/�ٙ"���36%�[[�_e�ڻ�js�l_���A�,_�E_�TD��%G��[���m�c�@�I���loNm����������RB��f����yO%J̼�r��>ɋ�����D��+�E���ː���n۫E�����l���GVfUQ�	8!$Үn>�]�$�B ��@��BNdr�YetT�+}��n����<��7�'u=pqf/�f!r����Ͽ�>{�薾�"A���3KN1�\��i8��+(e���pm- �]�?��䌲����>�@Df �9�"W�������Qx��>"�n��n|���D������$�`ȅ����2���0��_�z!����ۨ���̟2�Ew���$�@��B5��v�Q�.Hp.�~<�|A�3/��L��{���U^��6eg��y���������f*f@_��AL�헰f�-��I���n �9�"D��땽�0T^>��?z�|B��cz)E3M����x�@�}$��"A��$�3���1�B��f\�ͣ�M�|�h����H��A��٘�ffV���K�<M�s˛��B;m�!�Y�*����i��Z����*��,vY���K����<�r�]�����/�`�YB�n�
�»�jɵ��]0.�26�*�U�J��?��w�}���.#�Z[��S���Piq\�#LrV�R��u�f�����/�����T{n+��l���E۝�8�y�:��w&�lG:�wC.|� r�0������k��Ս�s�Tv��m���`���N��\1�T�.��k�p7n�nSg!q�n.w�~�ٖ3n6���7<k��mch�xЎBi\;G<��1&Ў6��;_� k�,XE��������T�h�o}#}�z}�סu���z	���{בr����9��7�N��R^#5/���Dϲ��9��%9�S��Z�������S2��{�j
6�29� ���9����bz�V��=���>�}sH��fO��]�����`���}RKdT�C��;��c#w$O����d �uǊݸ�q1M���i�D{�n\�2{���M�ߨQP�L���$�$����^���r�+ovL>�W����|A������_H�~2/�i�?OL��]���% �P��#]w4+2Xh1�c�KpgJ�;Z��
fٻ����]%�/�_ވP!�
2J�A1V�z'6�����3�"�7{ڳ#��R�d6��>���,"���*~�-���IT<��xMz��qm"NP�����,���:�Q�����uJʓ誴���[(Տ8ޑ�7����Uv�\�m�\�gaw��H �Bڮzϊ{g���o8o���k  A���\�,��>�j��o��H��RA� Fb_32Eo{r̝Oi����瘝Ӵ�~ֿ|A�ޖ,ȨL���ɑ^����A9S���� ���{{�9�4�_VFy���sܤ}b�Z���=���׍	2 �s#�32D��츁�}�GYa��p�����g�Ί�pW���� ���;٘���B�;Q��]��-20���fH����U�����p�v.�`:sqՔ�����um��?�r��.ԀE�̏�1
�{/���Y�i^>��!ċ1]�ڕ���9�O��T~�QJ�D�Z�%�Ͻ�0��V{z����ߩ�s�T3�����D�xO�a���fED�QIb�̅� s">�z��������Z�Y4h�Y���h�ij�Ӹ���)��N��#n�S[W36�rO2�����q��˴^+���7�&+5���7����iP��XP�U�֦��|j�P�.:��=�2�^Ϟ�wݦ��m�[X\(��նk��&��G�oh��k�������f쀎��9m�n�Xq!���؊�Z�xs����y�,X�R��sw�%fa3:ʻ�ӢC1],k�=ڭ���$Ê��b�9jXe�x8q��XF��1����זH��|x�\�������	�x��LҎ�9æ�cy�U�;C�ľ�zէu/s;v���Ԗ\[��nfS�F�z*V�"á�]v*�Y�/N���	����$�ի� ��
��!W��/2k��yo}�7��-�f�_-Ͱk�r�S��^��q�}T�˹�c
{%���r5��b��R����ǙB���o3���e�o����P�"�����`��%��1
�MG�Y�����W�uR�-��S��^�#�n��ޖ!g
�uAj���w{M�UVX���M<q(�c��r��M�3����������G���'mVwK��V���7l�) S؎�$��;2�u_r',W)Cf��צ�2^-��T]]��!U[,<�Q1�r�܅p�H���E}��Q��3 ���̗.���%�Z�q}��YU�F�S�jw_.ӗ6��UBV_v�E[�[�iDɝ��xs�w���'�v��黹(r���a�qZ����-�.��F�������]XhvV1����aV�a�f�&�V>�I2"e(���̪hj���G��rvw����n��K�;^�z�"�6w}�wҳ�v�V{jH^6�����H���f����Qa��)��[��q��:C��v�Z��벑�r!	mno�����_n�ξYyVYY'N��Ol��(�,6�G}������ƻC����L�HwYh[/�c�9����v�n����h�^Yu���bygY���'{^z����n��S��e|�/��8{h����u�����7e�^۶�����ϝ���{xu����Μ�݅�y��Z�����+��眾������o}�I[BZ�[�)�H�J\���YgkL�m�K�{��3eR2�ˡmZi��f��ûh�7�7��� � ��/� Q�%�M��8xD{'���$<�Df��fd�+0v���%yF������$tվN�2yv�5p� ��@�̑ ��Fb�D<�Ϡn��h��vv(�4��e�K9�/�?�_Kh Fd|ϟ>i���}%�O��mJ��n���~q�������ş@q�&�``3�.��?�������~�'2>G2�����G�ay��;�${�#6Q�㢼帀��F�Wِd}wk  ����Q��=�p#�_�++1��w�+�4�U�	�� �K�����%�0��~��`��d�FIV"Jf{Ԃ�+�x?>����9V�cg���=�~��/�IH��ú��1�9������q� ��Ckm��*���o8o���Md��ҽ����%�D��1�1^�@�=o6���36	5ns'F9'v��K�/���]֒��ZY�hUի�����syH^�Df%�f) � ���#�½꿚�2jޱ��+��Ss�k_~8���Ń"��ȏ~ݸ�/�����K�.@a�v�,��Z��ޤi�c��C���b
LB�Q�j���kA��~ ��^؎�ۯi����q|"��y]mz��;�Ur�­�㙒$�Bs!��un�BTƃ� wa���/�U��o8o���|A�_fb\^�s���9���_Oو���3$R#�voV����{�#4=�s�jo;�h��F��`���"�D��I��*������gJ��J��F?/��kL���c�����${�oq�5W��S���
9���2>C3$H9�4����W{������=�o4o���d �b�b�Fb���ޕp5Y�~�u�I�}�&��r�-�]��}^����(�;�bX7�g�g>ڭ���Jt��E�~ub��I��`E*ႊD(vN<�'²�V�fn��,{:*Yb���G[�a��]����w,�5f��+"aY�<��fT�	�<є��8�-��b�h�V��'=�ךx�zu�f2�Y����tp�!hE�$e�������u����q��v4jN�٬{s!u�r��Wn<B�����k��F��7;scqֺ'C^�;PohwQ�k�����kWc��Ϟ�����X���)1��-�Ir�/��v���n��EH3���>��o��e��1�f%�f!#=��gz�˳Sx��;�g;�i2��"����t|�̄Ff!?��.s2:�bUr��uꟈ�}[�6;6�l]�]F8��_g�H!����k���/��7��_WG��y~��s!|A9�d۪k�mS���r�����ސA���=� s1H��������\�Ƭ>�ѹ�_v��;P_��$t�����b�o]��p��Y�,W�9|��򯈒X	�
$��f%S���vn�F��w�Q�=�3�?�)��� �A|s2F�͎�������o��K��1nH5�F�Qg/�<���	v9�Ѫ�ƉI�&��>�������|��"Nd#�d!��y����c��y�}�#f�毸E�  ̡F?U���%
�L_vYiw_7EF�i5te�}�>�n��,�7�4�o����ּ%�/�x��4r�%���Z������t���B~�~�#��*Q<�_�"Gy��p�/����~m~��5DoJ�/m�'y �=/�x@8��jAz�3�Fb���-��,�[]V.�n�{�g N{��Ch/��A|FfH�s!��}Δč�V��=���H=��?fB�k:�G�]�m�����������yo<�J��*�,/�^� � 3<���?~�A��9�e�>����nG�����������6���ƫ�F��`Ⱦ�$w���7�}~�h���  ��" �O�c��=� ��ˢQ@��/5��7m�.ɐ����ɥ;�����?~� �7 ���X���X�xFr�`qrҜ����Ym�=3���/��	�}�g��������o�O��ݐ�Vm�#�wa�'�y�7��~���#���b>�톜Q�g�Ed'P@�w5}#1�A|~� �ԭW��Q�#7��>i\ZR��fWl��wDou�E�#N��T��7����1�]k~}Ktd�{[�U̛�����Er��y-�s�[����~ƨF��fd#�d FfH���}��w��p<������[Y{��Uٮ������s��K�qng�;�h��O/��H����̄9�"NdGO@�B�txO�ﴏ5��؟y�p�����A��H9�U��t=��-�	��6�W� ̭����X���툎 x��b.4��k��ѵm��?�~��jA����̑=/���9�����q�4�#iF�7��[]v��E�@���* �"�$����QR�y3OEg��w�Au�/��y���X\�N|�) ��#0��>���L�߹E�z�q}��2K�E�@2,��������=�b}��wPhp(�ԂhH!�:p��O����:�D�;R��r5^���8�s��׏o־�Y�;�_D=��e�{{[�J�s�YW�0���}�����\UPJ��e�������ܸ�w���Q=�k���ύ��f�I�����@��6[v%���8�ڐ~n��Km	����py�3�%.)4�Vӭ��Wy~��|�s��A�� �������'��}K�[��L4�+����}��q������Ӫ�$[,�),��a���T�W���=��"����R���[��5��c�<����}�E;�({��ܾ�܉6� ���/�<;�f;�� �=�D�޶W���O�_�q�G��%��2���k��b��_أ���2ǳP���m���ۑ.�gy:
�����ۊۛ��<��s���"@!��������TS[p�"�dH9��n+��t3�}}���<���kZ%�sla�R��D�K�ڒ�� 6��Owδ��=�����ٌ����O�_�pY�%����p��ǠW/V�}��6+�.�ڛF�����Eـ��t��l.l��C�������7Y��<����5��h⺪�R(P"�T.��k3SR �2�,u��lz���6GqS䨞Ss�Ys3�9v��m�B%��\�I�yA�<��Q�ӡ��3r �)_Nu��M�3�a��]6D��\�5�! ==��60mٕ�
�ѯ"�uL�;Xb]yKc�v����*�s
��0���]G�a1t]�z����k-��� ڹ��<�-�GV�t�]�u�v��������k���%�p�x����OFNv�H�oZ\ͥ
3vO������ZwP_��CnD�+=|���n=מ��\�=�舩RNٟ^O*#���3�_�r$��Kp�����P�F/yî�̾k����� �:�c�<���H?�BH�6��vF�cU䁷A���$6АCq�m���w0��r������ϰΌ��s�}����\&� ��Ȑ[j~ �� m����dOT��J������S�܉���λ��]Y�au�>����u{ۚ������{wj[jA���mK�΄�[[�����b���wzA5���A��ڐAm��.%��{=Kߐo�aPi�1gaa�e�͹�(y�욥0Z5�L0���&f L+�	��$�6@n�ŷ"v�����=�s�x��k�V���E����Q[.7��'�RA-�ͺ��h�X��^n�'�f:���|�ڬ��i�xLwk�9�����w6�s�$�G�A���㇏�%W������h�y�W���)����</�wjH?ot�ɾw�t�Vz��]hO�&s����"~!�x���Lz�I�����mȒ�RA-�y	���p�;]�h�ۦ5���g	�C���$4m� ����{Cӄ��5i�]܉��k�m�;~���g}�fz��z�	��
�3K���h�o�Az>mԂ[hH������y��{�"���ںۉ�]��	��g9H �����nE�/߷~�����ۨ����%t�u�2�[��)�SA&�s��dJM�q������,��|>_n����Kp�M�d�up�/�y�'w�w�ٻ�u���Z��� �RA��= ���A]"�]�B��h�Eb|CΑ?u�6g�;���׏�ָ�d"7���ѣ�$&Ӵ���Î#}�$�n�?[AڐA�#���U���O����6v�B
�[`��Now�$�\7{�����"�©I���q� *n�6�&���ZF�5Q�v�6v��k��[����}5��}7�.�'�g9I<rt�6�H����G�mm��Äfd|��ȓ��~ �[��t��|��c�<���	[�Iۑ��}QC�(�mO�7\�!�͵$܉!��&�ܞ�k�=����r�4y��Cxg׏�ֻ�	�����"K}V~�_�p�޾M���T%|�	�S����`�k�PֹC(d��R��&�m���2���H?��H#6����+=u��u���]w]�O��y�{����V��-��ڄ�Fr��n~m� ��욪n=2+�<�R' =YOK>����y�p�j�͠8sA|[k׆���[�6��܀������ w=��;\�,{cv��3����\A� ޹[h���p��k���A�A|v� �ۑ7�����A��X]�W�sܤ������~�i8���J�o��D��݋ks��l���{iwb�#W��۳U2v��"�ʥ)|+�
�rR���,)�Q1�Ep�K�3p/��	����A-�ɷ"Am����� ���o�*ٗX5�C�ᎏ��p�oH �BH<�@����nE�b�{��E�1�� ��X��GVd��λrM\7n�sx�k4�7��n�3(��ƲԐ@��Cq�mȞ��������^>���fq�z��u���g=�1�y�{V'{ܘ#���#�{k֢6N/1�;J~#7P��&�;��}���aw�_|�=�A�"A�G����)Gg������A �B��r$ڐA����7��K����a���y�}�?V��6���n@n�߫Dه�1P#kP�C����6�o�o��7�z��] =q�W��jv�Ɍ/�O�_B��܉����k�ڜ&+e	k|�x��:�kw��O�WU�����$6��_܆>C���;g�*Ǔ� m��H�w�V��-�X�<zZ;�;%L+kF��x�s�oE�t�Ua��.���7��~ܹ>�]D���V�3]ay�5t.�Y��r�l� s^�w;�U�X��uaB`|iR��\��A�>I�*ː.���ւ6S�n�ňaՒ�/�nة�^R{�W�o�m�Y�m^<&���}�U��_ZY�AY^�SS��ڕ�l�n��ޫ7X��;t�gaEk:���J�^([��;f����ce�EPpA�:kڻ���,�k�M�4��[[�oo2�C�o�nFR���vU՛���/��4�7k9V�i�*Or�n�׶�9�S_0R����2���Sw���f�\h����;[Lԥװ�\쮆��B��
�h��K��:Iy���u)fN�[P�'�'^����)�����&�E��*�;:y�G�����nm�qM!�-3-K�<�,�;�#.eV�+F���]�.�캮5��g���ԱvUw
����T��6���`u7C��D.�T��8ݚ��ݿt��#�9a��I��s�d�j!�)��w-q�Lܗ���I�+k�3l4]�7�g�6w�V"���dN�e��#i�Y���Y�ó���n\�7��j���JŞ�"X�T����%��5�����qa�!�0�ɷ�L��VP��.Ka_��h�^��O�F�I2|1��U
QY����w�bx���-����H����>��R�L��:�W][`?bUz�:�U�Í�.�Y.bU5�����z���1�
Rh�|!����ٿާ�����:��=�m�v�1���U	l>�Z�i�0�J-�mX[m�^,��,��, �^���d��LI��yȑיM���l���w���*mi�k,� ���=;/m�i�`��+�;dؐ��å���N�:8��%����׽�k������G$����kM��(��ΰ��-(��2YeB��$���˄��fr�r�¼��'K���(�#�Q#̑Z9�Z��9�M�:��V֜���C1ׅ�n�t.�. �8��^Z���6׵��+3����r=���!RG�n��8DFv����ma��^��eh���JC���G<��n@#�QA�N��H��m��
r#�{Z�;5���m�n�nq;#mۉ#����hm�m��9s��w�-��HF����!I��0[em��J$�.8�Sk���D9�e��/7!�	I����/mC�V+UJ��/w{���ffJ���PF��f��\��[s�X�Gv�mm�eh�-��s=#s��bg�¼e.��6�!��Jp�3�ƞ�%�5�9��n�A�%�Ko1��m��[�`��^�E�CM�����7A��ŬgOn��������)J/��v2tra����8���U�	J.5	ae�#4���A��%��q��j�0[���ݏ�����k�\���1y8���C�:z�f���I�m,-�T����T�M�pŗ�@�y:��i'��u��5����l��aฺ�Yx�\@�g����gOe�Gy�'%��^mR��X�++� l3�7��ܴ�x9ݛ �4n��z8f��1�+-��:���g���M��oQ�X�WO�����D��H���k$4)A,�n]/hŰ��Ņz��9���g�kmȶ�ܦ!#u��뗞'�.��;i隶ٺ�Pz��î��H�	��ck��y7A�Zg���VNnx�ޞ��,��視&ɴj1W��e��E��'c�p�s��v��aG�q�5n����]�"�m�x��Z��ֽ����.��Jx�Q����qꫜq��3���!�ult��d�{[h�=��`�NB��ȑ�y�=v��k�iphj�,��Ҷ��3f�c��0�BX�Z�5\�`mUc�[T�2���Mv+����_R�ݛ���t8=�{M˔ǵ��G�H�f�c�[����7�{өӦj	�n�q���)"q۵�qG'���j��8�j��!q�ݬ��8����B���{^ѝ����)�։bX,(�[�c�N�^���]g��Y��g���㞭�� v��.���I�ی�'9�B��b�kl+aZ���4-��Ltn�7ζ�m�ESn���
��n+���:.�ߛ�A���ں�����R�JuX���e��ɰ�*�P�n�Ԕ��Kr�0S��ܾ��&3�\;��9��'�]E�Q��s.���qF�"E��ׇi�\0z�+�Me��ew��������6W�c\B���g%ۓsWeR61ZS�7D�����-�b�L�ʺ��iE���� �:�h�F6��i�R�.ĵ��lx�իć<�Ʈ݆.G�ݳ���	�ˡacT)B��m)��ɥ�N���=���S��5p��f�Վ�� 5�c{�-�g���u��,�3������o�{+u'ؽZ8�O<ut��b�¿�����e��ѳ��BAm��!.�֏�eүc���H����<X��2�� �r$�� [j@!��.1b��{��cA�}��O�z�N�ޘld�����|~��#q�͵P�;#\N	>P���$���Am[jA�"�w�{�9�=p���=�{�g¼��aw�T3����ȒK��mH#Yң���Z�Q�މ;�$�j�~-����N��|˪�[���5���DM�i?r�M�A� 7H[k���$6f�O-��+�=y�Įs�0ع���\&�>[�D��R?��6D\����U.gA��$)͵:����-���LvD��m{v�l�PTʎ���O��A�A�R!�"�_���L�W���zw�
�x���"�߈=�"A����m���׋��T
��؟vzD%9�p�+���e�a�k�3ܫ8��vD����`�X���ۂn�9�1%Z�'Y
!LG7�:�9r��r�&f�~;�U�~�U}��:�V�U^��=���kBAsA�D{ұL}���WH�sR�"A��?6�OU�kq��7;잌w���\~���q�͵���/���Dx�G�\ ��JA�~� �/�nD�M�o��O�]U߰�ૂ�R].���7�~vWU���"�dH-�'��|Cm	-���g�U�
p�kX%����j����Zy��mI�+�-z׿���r��=�%(cPc���]5	��#a�r��۳Jؕ��6�.G׸�%����m������e��c���]��Db��J��i94;^O�#:П�g)[�Cng��l�hD�,q�/E|smH��Md���]i�7UwX��Er�r�7"A�������wЩ}��?�D܉����n��yR�٣	�cz����9Y>����P�lЛ\�^�1�#0����[#f+�Ԡubż����$����3������e�����$�/:N�����A;m	#�m}-�Ch![4���|/1Gj�.��?�/�����3f^�C��7�t��!�5����~]Zdq����� ���h"�Q�}a0t�>J0?�^ȟ�f�=�މ�qu�_	��O�1��_ۑ��U�6�#NEǽQ�)H��J@�m��a�Z´IeaR�f�f�a�.��be�ˇj�oo�?<���u�͵`�p�[�Nq��������|$���򦳜U��4(s�_�} 6�H!��m�tlm�L��#�>O�Fnp�S�z8���˥��d ;�~m�W�b}�%�|��$�B~ �� �ԂmȪ��M�v=��s���3�wx�Ep@�g9}?crt��܉����C���n��<�$z��p�㨱�����U�yµ��Am�$@���k���"*�ݞ8<��Ǽ�P�W�FC�Qީ�_�Eky`�]W���6pWH��pi�M�r�5��0{Τ�U��Ps
����.a\Ɉ�c������Ch/�jH!�"Hn�zT�>:o�MH���=����v_�M�e/��Dn4$ڟ��ƾ�鶯xډû���u�r�#ۧ�8�Dl��T����	��feI31�4'|$m�f��mI�܊��[�/�����V��+��68l�{�}��Ȓ��6�O��jH'�W�-�Y'U\'�� ��\x2v'�s�UU��Z�A ִ'�9�E�����|�J��;�$쀀;ܾ��nD��_nC��9��%I5ū��M7ה���d A�D�ړ�p���Bj�E_g�sWJ�}���CnD�O�wl�yy��\r��$)�3��ژcH�_/�{��m}e�@��[h��b缼�40����y��Һ�xz�����H&�� ���m�ې�V�����W�'j�� ���.;D���=���Ղ���;�Dk�>��bʛ�T��?{�M�}���u���y�XhSprǶ�LV�r��-5@��B�Ѥ�[ �[��[[��U4[�aQa+.F�ŸH�E�S0�zޣ��	�5\%Еź�!u�%���ɱ���v�`��3��x��yƄJ$6���Ŗ��H5��e�mnVиh�)�8hB�F��]5݋�N�õ���}N<7-/�coooj+�=�^��=t�{]�d���=���۟�uu5bj�R͍�z������t%�Ìb�1��V�@	���6+�-��
�F�ڱ�t���y}Yk��"A��m����?v_����_P٢�{3f"\�*85���U�Ÿ_ۙ������Z����vѵ0�������}sݳ��}�ux]p����/�6�H!����iǣmߗMȟ�<@v�����Ÿ�#]�Ϟ����:�rV+��=uV����ZП�9��ڢm��\�ꆻD�'�h ��G4� 6�K�;Lk�v_��u�. �r����!Q�T������ٰ���A���[A|[iE�m�?,�r$�������}�ux]p��?�)6В_/�͹��r5���$BS0�R�K�8-?ϝ��|�e�c0^�'vp�n��nyX�
������@�?gH��m �&s���
��w�m�)�5j�'=܅��Ƥ�@7A|�S�!tǄ;��jV'l/�m��^�`N��q�"����Ε[�U��op��2U_c�[��� Ε��nQ:X��]ͻz���Je/^�?k��w��G1y駝�K� ƾ���,��t��_"�0O��}{4X ��$[Aڟ�-�q�"��T�O��&z������<�=�H-�m/�hH-��ӷ3hz}3� ~۹w�ŸBX���u�q���|6��hO�B����I�F�w�����C.㾬j�}"Hm @-����I�r�kf����ڑ#h>�k��禞ve .���D�ڐA-��ޘ.tl4����.��b,��b�ؠ|��u�]k�wc(!"B0Tʍ��H&��@��mO�ۑ/'�=�=�Fe�^\*yw��E�:��A�� �?6��ڲŸD;���9�5�/���H?���6-��}Ʋ����} �ք�Ftm,rVp�°{螐+� G��) �ۑ ��|CnEծz�A���eDBE�D�ȭ���c�б�J��G6�*�g:�a�gW�y5"��j�f���oƄ�_�m΍b��O;2�N\ E�_6��~����UC�2."h�͋�<#-�{�~ ��Nd���OtH�wW��]��O�ZӮ�6����ρ����D�ڒ	n�nD����{�9a�9���Ju��s=V������ �9��k�m��n��30�L���z�f�Bci�G4�4�A�3����6�tZz�ۊ�i�32�r�^�����F{���l_܉����Pu=��M<��\G�kTև.�o�i�{"~6�I����RŶ��Eo[��7}�$�jH��/�z��H�wW�օ\'=�A�"Ho��t�l,��=�"A��?��� �ۑ%���-����ϊ������Ng����} �ք�A�ڐCm	!����T�ǪN`����ޑ �Ծ?6�H��j����/*i�fR� �DZ�l���]gMw�S����a�?Lʯ/B�Λ�Z+d�F��'\ҕk¥<���Xp�U&��
n�t{ʕW����*��9� neě˺����?A{6�H �П�!�-����'�%0r�T�~[Ѿ.�ch��'=�H?6�I��m�kݫ%t�3S�5��	��!��VSd�z�[z�s�,�5��[ �k�2b5e�������j� ��L�b�+����z����/��x�x�	kqu@G�T�!�"Hm Am���|zx!E-��4���gl��{�6#S��^T��̥���@�/\��P����GOG����}>hP=�-��-��ۑ��8�o)��W�\x9~����&�p9�S�6�H!������[k�Ӏ�݉nȐwuH ��	�,[%{���g����|$ZБ�.�8Ψ��x����_1��I��m��� 6/I��U�^�%���D��w�qZ��b��O;2�5���_6�[�����E����'����V�e���8�.��n_���2�q�e-O.���a��tӸ�ns�*�a�I�oo*�mo�a�P#!�r��~>�_r��b�4�m.W��(�ɭ��ꨭ;�U��q� �:���X�Q��WH�W8�{s-��f�Zz9�Ӧ�KrX͒�t�����sK8��Cp�'\�nuYS��d����ԉ�q�����ƪ����0��Z*����}�C�k��:�k,��l�K���rz���fb�^+Riu1�5q��.���g���i>�-Ք%Q�u#��6-�\��HKmM�6�k٬�L�J��} ��! �3�E��[r$Z˭�;�Ó�M�~�5�n#�q�y�}��"Hn>m�_ڟ�%�DD�Q�1;1&y�5֤A{L�b�+�ݝ��w�m�Ƶ�'��թ��O[3}r�otgZFRsuH �܉ ����܉��p���o��G��ã=���.��d"�r$���s#����uU�z)
����W�܋��v��^��X�:&�}��?��w&�c.��#�/�����An>M�mz������ѷ��TR�7A[�����[�o��kZA�͵D6�C�򣇸r�g���x&H&��� AH()���Z- Xr��j�,�%C�$��T�^�
�j�3���|d�7�z�Enx�y�v��W���|Dޡ'�� �[��Ƅ�<�E���>�1��7��u�_���5UQ���n��7��]ilI۴�~�+�\�,c��r���9��/�����-�FxP.�}#�dH��ۍ�t��J�9�7�g9I�D�Cn,�+��l���}��9j�O���_~mȒ�RA�����~r�H�=W�3rs�n�V�	�Y�I�h [k�����|b:��y�˟rs��f��6�H��㵕/x������A��G�	o������jH'|�B�m�$76����[g�=�d�1�2dKV���T��J�9�7� ~3���ۑ ����܍��=}dթ0R$��OQհK,n.�O<�Qf؈gL"�ͭd6�g�!xlIJ	B��.kao�O͵dp�S��8+}���rj��Α/]Y��ǰC��4�����r�AmȒ_ Am��M`J��[q�����"�cWn8�ܱ~���� A5��n9���J���F:7'�����]2	�hH �����[r/���τajn
�K�(uZ�<U�S��x���-�FNR:`���}�F(d��]��i�Ca���2��F�nټw|l�$E��olM�q,9N��gr�ժ1J�J�eu��#*���w]E��/Vhgº�ʰ���n}E2}�&i�j�0�a�ݻ�h#���/W*}}���V�����D���ʫ���^���u��\��{�)]m���9%Q��q���B�K]+1��]_�
�S{�`o=�԰¨�X���
�����}Xv}�<][w[�F���û���l�+k�������ؚm!Y0Z*�OV�wF�:;!�T7�M�ܩ�pX�6q�3�a�֨\�����v�wd���mc˙�H^	����{���ш���}v�mԶ�H���5�"�r��ռ�0>���!Q���rL�n��4�b���@��9�slZ�62��yfJ�U�[�nn�}��%�[4���l[���n&v�]\�v�e��fu��K3�n��&'U��w*f�B�oN�<�f�F�IT�;��l/�ҩI�pf
���>�<��D�%�;	+5���^㪣R�O.E�tX-)n��xV<����\QUf�L�zf�՗WWW;GE�b��wfI�����-= �Ч�jO%i�s-_���Ŗ�mi�/����ڿ��D򓻶&c��u�N�G��od�����뮂��[�q�M�F	���%f9I֧7���s]��7N���Sh��ާujV�qU
�v8�G�̒�*�O����՘�m{�y���O��
�^�}}j�}��ycnm>nު�y����9؊�_;�j�R����A/�IY"�B\̭�-������"���׽��,�p˴f�$!:N6������{`��3=��GL�-��۲p!�98��8	!��q���v��r'8��CnȒr{e�fB6Ȝ��鼭�[c��ݝ�DF��'9��4�㤜t���N�6�Gq��A�q{]����	9�k-39�F�'���{Ӗۂ��,��Nvڑ�bAE���h8�Ӥ����i�����	(���aם�����3��m�Ye�C6v89)�.������D���"�.s�{��.(zm�ݽ��8�{�G����\Gw�rOl��F[�3,��HG8tu����@���"\<�9�qy�w��7�z�e��8N�����v�ڲ;�Qi�k���'�9<������%�v��I�^we��Q�%*�)EKe}�oO9ϲ�;.Ռs�o�@��_HmȒ��k��3Ӕ:.=Og8���%�RA-��)�o ���ɻw·8Oխ	�0��N.~��و��5?{6D�H[jH!� 7�3M㳻�C��n��8R���T�U�q�B#q�%���q����}�E�>��`�B��J �DQ�4#��'�ې��y�Υ�.�@� j�
خ��y뀐MsBAv��j��܉��,��LP�v�c�|�&grg����;W*�dz��_/�nD�^5 �[��G�4�n����� ��/c�F�����]��} ��B~ �h mg��i]q�l��r��Gb@�椂r$����ۑ˧�Gay����rv��g��=M�z��!/Z���Kp�m��n(6�2���Fds�[r$T�{�:]���	�� �s�MzGE�+��b:�B�4onk��"n,��/�c:%[��u%�o�|�c�W�t�v������PL6�C<w�ۼ"�^��i.���?���ڄ��RA-���۟�k�9cE��� ǡ����)}{�n��𭾐~5���~������nBw��R�YG��6ݬH��P�������CY�κ���D8��B(�fd�2�'�iꟈ#�dI���:��':e�:9�o�־��8�Ї�����ov!{2D�澟�p�!�"A����@�Ԙ�G,OW�	�1��Ԑ{zD��{��]͌s�nΫӬ��:�f9��O��w�s��[r$�ԐKq~̭��u7�/�/��R��F]]��[} �XП�?sA�_Kn@n�훷��>U;�b�A��Ώ�͹ץ�>�k{��߭�����񬏽�ۯm�x�[����A�����܉��A�U�k�ι�!ж9[���ƥ���6���qΉ��^�!���Cq��[���EA��x�&������tD1�Y���<�{?L�$"��5�y�U*��8M�Yn�7ʖ$��wKv����"����]�&�Yo]Չ͘6�b�a���!�Q��9�m�0J�Y�!�����Y9+u����vծ��^�"p��M�4#�ev�I��ǉ����ƤR��M@��L.E[�]rY�z��O�Q�h;[G�vM���٩H\Zʒ�i !8@��5��Ɲ�Y�l0��c�R۝es���$e�8�CM�`�l�Չ1a5eÈ�V[��=_��H�LZ�BU�2�5օ�kk-����+�5۴V���;�b9;\A��G�v�����p�S��T��싫�|+o��s����s�e$$�+P@����t�ڒ.]k���J�*ށYa|w\��݆����?���t���"ۑ?��g3� �����!�BK�BH!�-����0�u�������̙�-��Ks�k�?�)�r'�Ch/�mȐ[j@"W?>u;۱��2�D��_In#��f`'��˛�z5�	�ZВ.�l�9����K��D��@�[k��C|����_�R'��~�K���签���k!�܉ �Ԁ~n+=�)��1��"&�;b�Q��i�ز2�w��qE�Sv63���k7��U�U���=�,�G��ǽ�̍�����Lԝ~����5�FM�oMK��Q��_^^H�3P_ۑ%����"=8��g޺
���9�m��f�c��2W��v�^���3��J�r�y���Q����]��<����[^De_���}'� ��f~�ά�]��:~�hI��ч,GI�/[�痡W��Fr��� ���_�ȿ<G	���8vS���,g������d/�xАm �W�6�����Uˮ�sh`"��澟�r)u��9;w��k����?2+-"��oX�Ch/��\�-��[��$��{��)�[�����n����nmVU۽���kBAsA��6��˻Jܟ�w���87�A�r��E��h�6���������ƴ�Fٛ�{~2�_�������Hn>M�����ʎ�c=m�]."��z\8쪉/�D���~q�n���m� ��2�%G���Ɵf��c�s�Nt���؆�W/�r�AmȒ��=���y|��ι�ݯ����"~-�$�q�w/o�����3+��W����h��:�^dIR����h��R�3C��ývL�R^���q}xY�˝/3�97]�%�>�}���{���B�>��*��o��MkBA�h [jA�܀�!=��百Ӓ���Ȓ5�ŷ#w5�ά�������R� �B!i���F��o�y��_MI�ۙ����A���mk����ޝ޶3ީ-=�yz�/u؆�_.�I<rt�m�W�"D�C	=�	I� :��V�׍�Z���Ix��֔&�jG*W1��(������t Gg!?�����g�%���u�v�k���BcG�{ֆ�] ��)܉!� ڟ����}�ϮT�[Z#�|w6D���ΧQ��X�m�V/��@��"KmB8^*=���Xc@70��d��	m�m�!�����k�'<r W�*(Nu���u؆�_|�>|��܀�/�n~m���`���&eN��F{$H:�}?��ul�$���u�v�k�ִ$$o\Y1���P��T;:��Ww�������ة�L���SI���M	D�m��_�V��][p�fǍ�rةVDݢu~���j�����3��3zD�_ A���ۑ ��
ܺw�=�;�u��{��;���,y�>���~5�� �r'��R%������Y螁�P# �s�<t�u�i�Xe���x��Y��]�QN���Rk�#u[jHm�k�y����m؆��_!���vWz��]v���Fv�;�������	x�(�B�}�z(�R?��l�P}]��*��o���u	���[k9�W6���:���r$���S��"Hm|�!�#�W��u��Op�/n�K�ǝ�Ֆ�[r$���[��u"�o��}�y	 �?e���Q�-m�7�ެ3U�
oG��RGw�va�2���X��-��#�Ȑ[j~ ���ۑ ����j��CFg�0�y����o��.��Ƈ ku	 �A|[k�m�XQ팍��z����S�,��u,ZN�Y����U:l�c����;cv	��}��O�޴9D0�9�>!�Y�]�f�h�_۔A4M!uF���/]�F�=]��<�"�/]�k3+���ڵ�B0����	|�i�,n�m��N٘���7��\u��LM�;]�7Cr���s�9ݓ���1͐��;�iPg��7��Y�Ny�Y�ǁ��%����ԗaBZ��``;sɝn."�<g(q�6MX����9n�Y�IJ�`�Fi��sڱŬ���7i5p7]a+��{�o�? F\�c�^�+�دg�+Q�gSA��:��;qr"�D+�Y��R#�Ȑm|�!�"{w}�˙>v�VZ�;��'������|�H3��~?7���ʹ$�]=eOޯ9�[ǅ|s֤_9s��]U�5�b|=|����mȐn|�]���������V��	ޏ�nD�[k����z���U�+k�;ʪy�s{��[�I�k�گ�?6�I����TK���mȟ�n>M�m���n��s���_p�ʇG�5z�l)��f������_Oʹ$�_6׭�Z�Dj[�@^r'�����g�z�D���������I�ʹ��/z*Q������L1eHG]m����q+-Wi����)��v�!1�W����B�mO�[��.�zP�>�w��y�szF��y���I���T?܉!������i�l�u�Ό��^V�xU�l�Ң���U�-I��4��Q�� R]�,�L=Kn+$v�~P�Ǳ-�V7ۻ�����k""��;#�/���}z/��5��m�e� �����[r$����p���,��`30�U?H ��$Ck��������O����z��}v����� ��Amȟ�������sV{t��u�.����D�|Ԃ	nޜ�q�C=���W���C�5���rE�V�����R�/�	���@��R!�"~!��4���q��y�x���z/�Ts'����\'�m�[j~ ��پ��[]f���� �`J���RP��Ǎ��=3�=s L�Z�($�m��]nC!�{�Y���� �����܉����w{.��v���/o�9/��+1	n��mȒ�R �V�4{_J����5�H ����[>��kx��z�ṽ ��BH s_6׽�V�@���q����ۑ$c����!��zޑ��8*Ķ�b��ڔ��n����Rx��I���lڼ�s�e9Yڳu���O�[����2M-��0��^��mb,1�m�e����|�܉��-�!�24z�h��:�_U ��S�6�M��q����z�*o�W	�� �s���Y�TL�џ��_�9�m���[���"Am��f��m���1�����3�#k��g�M��hq��$���RA�279zG�1 �B`(R"L�/��k�非7�Fq�q{"%��Ն��f����z���o��/�mȚת��\v����S���^�a���C�B@6ڐA-�!����@U�\����>�$��.hs���]uՅM��w�z�|�B�����M�~|+� x�������=�ps:�,�"�5�sl:��g�M��hq��'�A�E���nD�Ch!����#Z�#�АGr_6��=^|�/�F�'{N�|A���O�֡����'�� ��5���o�S���˼OD�E�2��>���Lҏ����}K�46�:��n�ׇ0�cOݛ�$|-fIR
�%��X{���َ����]�#�	n>m���BA6�-�t�Pz�o=��c���d�ר+oG� ���CnD�@/�m�S�z+�>WJ/��-�O��E�K-�cW���A�[C��3k��e�v;R9Q3;���O}����/~����[R ��U�9R6�g
�z���H>������s��`Fr㯔�Am����mI���:�>�kD�����O���}��8X�m�;\'��m	���{vf�h�y�(�F�O��� ��k�ڠ!�"���V@�eP몎�dۯPV�>@�z�I�'�K��n~m�"�d[���{Q��'nD����p�����N���W�[|7n�<���{N�=�g������@�[jA6�I��Vlh�� 4��zP�q7��o|#E9'lu�	ƾ��}$������������$�� �$���B�T����!I?����`�$��BI��!	'� �$��BI� �$��B�T���@$O섐�� �!$�0BO� �!$�BO� �!$��BN@!I?�b��L��WUk�� � � ���{ϻ ���ï> 4P  
P @   	 
  �       �    �g� #D�P (� �D @�E���JP
Q*��
BI(J �!�� (�)J(""�H�IR"J��
�"�
 (�JHUQ@���T � $�C�  Z����H��^}Ru���G6"�t���3�Y�vDr4p��
�s�*����� n��9H��(� N�S���]��`�� �a��t���W  {���  ެ�B�� z	QJ�)_   ��*UB  ��q��}^��N��W�{�J�ΕU[�V�ǭU��]��Ԯ�Ԫ��T�t.l$��J��(�  q�d:}�t(�U��Svq
�� rky��p�\ 6�=�o0b� ��� �P  ��Ƣ֠L
$)D(E)*%���@Q�3�G@@3�*������;� n�=9 y�IW c�Q݀�P�);�l�J���x����#��]�(� ��@�8�́S���O:� [(���;����Q@|�H��R���B ����G����@��n(��l `q� uGw� x���#�@�P">� 8v z7n�ܩ����z�n`<�	t�`�:��G��tH b�@*�@	�  � T��U(P��3RNN�Ӑ�N�{�����wo{Q��e��S.�]�zW�7;\��=�w�D�@UI�  s��a�/N];Z�����ZӋ��5��\bw���n�msʤ�=�W� �w�x�v4�;��{�    �~�L�R�@       E=�)R�` L 	��`��5R����4�`L��#!��M��Ф����4 4� �)���J2h��hɄ��0�	�DCRF����mLj4�3�����>g�3�}��}�z�P��#��7C�Z�z���D$�G�򍟢 �/���ZBHBI ���R��� @!
D�w���$�����h,?ٮ�M4` !2X/󄄀B����4&�i�H!q���9�O���_������ �*�O�*dɦ�[���^Ð�A��������^^,`�2`����)[�F;8�E]]<��Q��@���w(���u	���J�]���^J�71��h\���+wf�/^ӭ��q�Y8�`.W8[z5n��Z&���tq�F����B�%u��h"�)1��3B�w����WWM 4��`⻺��\FQVm�V�n�m��ia2�5`O~R�;�¦1fY�:�������{p�WH=�N�K��m�2�n�Zsۃ�#L�E<Y`�[G6���N����M�iU��%kݫU��Z�Fk(my4�x+Ul;j�p%{����̩vkq6��Ti�70̰K��l=�*�4Zzv�eS��M�t_�]b��^Pg��^dSn��Ц��M�M�Ch41l��q
W��+��xkK�0	��z��Pka7r�hÒ�ЌnT%�D�[r���B0�n���ӳ�6�ų�G�҆��f˱%��e����1L&]���1K�ch���x/E��&%��ɡ�Ҹ%`Dl"��I��NQ[��ͼrD/r�9���Ge���+˴GCj��\���ګ32�ɠr+&*�f��3m�-K�G#�.��4ڹH2E��F�v��d�k.� �����Zٹ�]�׿�����hX�f���C��cY�X���Z�י��e�,VZ�ؒpV�lK�Z�H��i��f�v�i��-mM�J�IyI����{HRͬ�l�������iY�\5����q�-�4om8j�1�ѬXko+bN��8���Za��6�(6b�&��R:�-gt��Na�`o��,�em����+R��q�u�y4��Z�X6�̼���B��3������M`@E�٣^�QP,�X�m�&1i�ùD�j�`�U�1n��kv�^�I��UHU~/�K��7k�GDc,X�u���R��i��Gw+5R[6Q�h�Rљ�+,1^>ֆy����w��,L�`l�i�tl����}(\ӭ��Av�̲)�Q�C����歖*�jPE�͕��,E8%�>$���%���ԡ��-\��wu�v�T��XZX[O!������N�a�(�+���r�*�h����`�v"��f���2�1���!���7�(�p31��W�`R�Z"�S�f�4!2�V����ԩ�f@n�k�M7���_X���%��1@��tۚ��TPR�jBv�*�pRNS�e���-=R��8Z�U�ܻ�/r[T���lgeP���ۘ)��X���f����̬�L��k5!�0'�+Q��٨� �k2d��f����/ԋU��h�.:e��l쿋�s촨|�� ��V��~�뷎���U[��mB�]l�S��0^h��ױ��N]��O>�9��%g�X��z�*�e2d�o��5�5���b�E�[d�E�=�򈌽%뗒	fǣm-֊u�U�!Kc;MѼc5dQ���U��(f u�F��W�6�[h��u��D�#�wm�*��52�NЁh�l71�gJ܈�u�kTǵ:��晪7��דm����,e�Ւe"a4�Sݹ��
�����ƆPukb���T�.���a��e\I,��	L�N���Y��0��YX��$��on-���H����[��d�gMѺ�kq����n]��7j�`��5Q�u�n�V^�Y+h�V�U���WiM�2	��$��n��u7E��yyn^`̬X]��q���[w��Tͺ$ۡn)/%��hj�6k7I�kCt�g�BnmU"y��n	[q���0�x����ni����д:��wCVq���fe�J�%�'Nf �X�X�K8��j�+I�1}J����e97.�s5U�sI��`6��o(Gְ�s3�z�k,Q������b!ZrCX[��;����d��J��k^)�4����ۋK�Z��í̤��2fŐ]e��ʄD�w�-4�nD�0mZu6�vK�]K.X5&�U� 8@"��؆(��'6��8)�M�B0�ïNʠ�Vfѫa�z����Q���cͱ�yN�65�S�ƛ�Ǘ�7YvA�r:�&��ޫ��u��O̖�<ܽ��:�B\t�V9�ƕ�C�Ǣ,��wx塴Z*��/1ڸm�*̱6VZF���Z�r��]3�(Ҹ��.��J��^�{Ln����k0Zˬ�	��ڦ�4���x��֩����~t�ǛK̃�O��[	��D+���]��a]К7FlTf���l�ѫ)�� V�BB�X�M����Ws/b��a��u�n���!��;�5x�V�l��-S��tD-
s(!OY�Va�&e�u���B�7�����J2��"1�N}��V�ɱ\��֑T�R �]��mѠ#��w�ʲ�p���JU6�)�e�L�G'��d�4ʿ�3i#4�t~��v1��o4��[yj���&�3M᱄�zͤ�c��7F��E/I�F!�jYǀf��Ot�����xX��"�ޜ�������uV(e$����;�Ղ_MB�lt�͋*n\�#M7(<Kkې	Zu��*�3�1�~Tk��j��Գ+mZ�vƀ]DOP���j�){J��]�ٛK�BL�c����X�V� {��$;H��hnF%m��X��,�y�&�{Z�۰in���K�So2�Vw)V���0�(�M�wJ��!�*�Q��KV����V�����;���T�6�a���kU�,,Ɨ���z�:jU�B�i����P��{3�˴UeF#
�)�)�1'Y�Ie8�z՛͙�x-Vn�Ih�T�l�@��+h���q�a� 	�Z��PV�!��T�X��[�eV��Z �c�)��b�w�N(�1[􉫹z~ �n�Yv�!UhI�ik�V�Z��X��Y�f��w%©��2n�����؛O����\�Ȅǚ^-% ��0l<ڱ-P"U�R��rG�Sb(o$VfQئV�G�j��>���+:IN��YV�5f��Y��R�мd��N-C^���:��e��iV�oc����l0a�s�s1� �9n�goՉ&�ǁ��d�(��"��/V�i
x���Y��'	��n�.�m������Sy��S#8�.C372+y�d��Nk���Ɯ�vܮ���xX�t�v@)\U�Z��F^�'w6��ϗŝ�[c�ȡ�V�+^c�]�E'�lA�M�B����&�Y�����Ё
�c�-g�1��Cv�U/�cÄ���_KgXѷ�"��F^؅3��[#>C-�9�n-t󆮘���`bv�t�Fҧ������%��	�ͼ�4«�dn���'uie�;i	k,ڑM�bS�ѳf�q�j��Q�U��U��©R�Z�	f��G�kP�⼠��d#Qf��B�5d�fL�[�`�r�!Orj��^�{z�5_�ۃ�HX�inJ��-�zd����B��Y�]��b�p���L����L�Q�E�@E{B�4�����UדU��"�,��, W��G-�˸@�d́|��.cr�]�An���+-�[���IXڧq�6�Ն�AV�8��j���]�4#KK-Fɕ �Y�BjSfKwqI�NH-mH�7�l�{� #.	2��ʎ/.#P���r������&7[y�������˪��-셅
¦��D�*��ssVe�O3mc��7��U/H����Dn��΍K^��W�6��{yWti�%a� ���)k�J!��n�Y�a���h�X�{b����)a��LӬ:��c���(���`�(8ȵ/Mfn��[[X�-��R�)[�7�V0�x���kF�o����a���-��Dp�+[�(���c�S����HX���R�11Z�G����a�i�y��z��<��'��q��NZ ��r��(�\��֛?X�d��#+n;8��&Z͹��¶2���.�r�e�6���n�3]�A=��2cXq�8i�Nދ�����AGv��@!۷E���WY6��-G6�V��d�k42���X,�y���]�I
�H�яnк�- ���H[�T1��(�yb��wYm^'B�k9[N�6��]0^`2=)���e�9r�5 b8l�j���X�"4��2ٽ�F\ �4�Ǥ�*�:���"�{T��ے�t���a;�i���͛���$)�ܰ�sIW��;��W+.Tso)e�G#N���`�t�3S)�!�m�3e Ż{e�Z�y!;lѫy�2*P�OU�S�ڻ2�:6�������k��E����/�𱛈�YL���VG  ����Ѳ���C/�,-YD�n�2LآqZ � $!SeK�ZH�Y)�{"ՙ�Ь�A�Xr�Y�40�٥`��R��DEn���֩�#�v��eZ�wK;J��u3f��"�n^u��׭R�e Z5m�a��3&���;*9�:�jnb��y�q=�׷CfٸۚK�܌��[�V�є�uj��J��e�o�Y�J�m�U$�OZ��%�Z�t�-��ܪ5��N^�3(AJ,b%�b��={2���.��dNd�u���-�^n9$�9h�*���i�.慱�ZF���X���;��mYIIX���-��E������l�D-+��1o0�.\m�E��M���mV�l��F��4Um�Z݉�B�U�	��(ᦐz���{���^Ô*[�je����͗+����M�����ov"錺�����.�qejeA����
J�JC-V�_Y6���m�7��s^!�o���mڼ��R�R[j�㩘�M�"���e����.����5NCe��ѻ���`��	5m�6��� ۺݗ@�[vn��3uS�b�ܔc�f�r��)2v���EѦʬ2�	�G�f`�B^4��lea��X�oō"%Q��.�ɯY�wSwE*4������7L[��R��2����j��pn�h=!�Պ�H���
7�/N�	���4�/r�f:�kw.�
�EҎV��d��k����ɪ�ʍ�sh�������k��S쫾��\�ت�LnKwI��n�k�h��;�[i����ූqm��5��:�I��l��J�tDثU����4���-{Oljk`��i;�|��&��ڻ��ȴuӚgŊ�I�β��dXc7m7NVfT��	=�:,]\�nꎡ��u�s7�	g�f�	�-�U��.��~|���^:��A�C��^<Bƽn�fX�.H1���!#�EMb���w��}�T�l�Җ�;)���O
8j��@G�y�@�2��{Kv�a����:���:���ܥ���/)Q�ԹR���ƦXd�`DC���e��P���MCCn�jt6�|h�̔�K`v63^d�w�n,�,JX76�m�+�çq*��Õ���-���f��^�d�v�Gk!F��&R�V�9E�+olV3v�Ø��M��l+M��������X��IC����f7�~��Dj�WyX��s6Tہ�75fav����*ƥOaн:С��'m���e�v��W��;�GE�2�.E���Lܴdɏ0A�@s�i^�;̅m�"V��ZL��h��s+w��eZ,a�r�Ŕ �bbI%��aed
:��,��Ǧ�f�Lugq�F4M��K��ER��P�s*�c�)h�z5�TGY�f������]�F��m��S�zR�P˳�h�5t��Bm�/6Z�,̰
�7fUm��2䂎��,�N�j�ܛ���$��%�m`��9yhҤ]M�ub�L��-f�;�&]�UP���ݗE��Q�r(��)�ɷ��Q�0!�0��g�L�;��M�n�.���W>�wbZ��a��;SE�YmVe�
�f�h�H�/*^""���v1`2e�4w���Q�R]�B����Ɛ#ywm�$%;�0k�N`�x�ܗt���b2��vHiL�Nj�
wtm��h�� r�;-�UZ�)���x��n?���\���[lOQ��# ��4���h�HI6	��:����:���뎺��*�;���.�躻�;�*����꣺ꋻ��ꋫ�����軸��ꎫ������㻮;���㫣��躸�������+��뺻�뎫������뫋����;��뢢�����������㫺�.����K��������룺��������������⺻������뢣�닸���.��㪸�������:����:��:���������#��~>?;3�����?}�ڐ���fno`!!_ܡ�"�йH@B���5g�>O�3�>�j�#�5;7����w������}X��Wk��s��K/���'�r�<��n�񾬬��I+��2ޠ!v��[���!i�LI%�d�bv�n��G�a''���aƆ �j���Yj32&(M�v,�~;���^����n6D�O}�!W"�x�#��|��;�u�F�J�0���S*�-��!c��S��=���������;��WW5j(��G���k/�ɤx�)5�t�OJ���!x��6�	=~ղj͎
��*TG�X���YU��ۺ�Eh�q��:)��F�n	��݁��9�}�k{���'J]rc4;6f\K�={��;$�����8ls�Vz��N{IvZ�1��f�b&w]�ا/����n����#�c�Eζ1�Z�U����\�5 �sW�I�u���}\.A�6��	�%�M�[B��ӷ$��Ѭ$��u��+j��\w5�}<T����F|�YĵC��^I�EL2�,-t��vƆ����'��we����w*A�Ήn�j�@8.;��De���5�+ ��A/��!��l�]4pbղ��p:��Ů��]�K5
[ט�bQg<�s��
�>+��s0���3��\�<*����J�c^8�5g�L��#�
p� �����6�%ݗ�ǅ�	�`F�k�r�8neL8��vlYչ����ԏ�/�˧B��B!|V���@�C6�.���8�SܵRK���^��q��Np�3w�v�'�z�(̨��/t$drL�޽�����T���:."]��oE4tvP�EZMN)0�d���RS
�©5�k�[�2�-��溷(���H��KKOU� ����f����޷	�U��j�\z�Eಇ^��Z�T���ۆS�����%{C�FV�<�k�jk\�n����6�&�Pu����+�?ly�;F��];6%�f�Π��X�c%*�i܀-'s�I�rjw�V����y�/�I��&5��`�dAB#���)�C&M��b��fMH��,�)�#.mf>�i�eڍ��MN��!Xf���XYwuqÄ�K�.���EB���h�u��%f����(C8jT��p�$���+�w(��R�shr���Эأb�s�8 �����#��T�3��E[і���7qz���z�e$<n�_���[1�//wj|{wG��ogG�1�ƈ����N���㨛�1:�5�^��3(���ć0f*~b���Z����o+B��i"�1i9��xV���٫U�jj�z��Ø{�AWd�[uȳ���j�&*2X.��7�r`�uxE��T��T�G�^̻.�ݣ��Qg嬲�M�)�u�����Sȣ�s*�]�̅ꇶtt�+�gL�(�C�:�n`�6�fFnؑJ��:2��W���6ȬᖆFH��+/�a�W���edn��!��BIxtd�W�Zl`x���L�ȑs%Մ��=���U{�
��y[�ڻ��ܦ�mc����k�q���f���W���J��7�Ъ�����A���C/|}��Ƕ���\�U���ώ]k73zc�ƶѲ�z�#H���"'A�����p������N�)�^����P��^^��������2�N��d֎�Ul�v<i��jƍ|Uc���I	���G��ivi{kqر��Y��=�VQ�{s-�lכ�1�z$�@Cܛ�)��Gy�<e��6��=�G+�3��(W��y�SJv�t�eսO�U��>ÕݻBƂ���0�3��e5���:Il�T������wq�Ybg��L�
��;�s�����m�wP��Md9Hd���Yf	���ߒ�W��hpa1�O�[�ȥ\��%Ѳn>Y:���i�C���e����H �t�g�^��H٬��cB�T�a���ܘ&�����c5Y��-��+�K5f�=���X�ڔ�޾ĺ��mҕ4��ޡ3���S���?�����FU����ے��vnӹ�^'�[[
���F�a5���Y����kC)Z�O(3�
��fn](�H�r��
�˩�g1n,�q�]����)�]�ǳU���j]���f���Yja�լ�-�:��Qɕ��c�����yP�����F���YD��%��bj�RILu�f-pu�����L:lciKF����!�{̻!b��/��6����XP|�K��3o;vૻU	�Rߎ��]�!���\��V�/0�%�]@eVh�̄8Q] �|���-�!NoM3Q	N�D,:*9�A�&g��<��@�'g�����F�G�%�ڎP��D*���r^���G/+1�J#�\az�[��}ڡMۋ#Ůg����cw�Y�ڝK^��-�lV�U^G�zI�B�l,���c�r6a�}t����QG}e�V��je^�yr��=Ӽ�cf���к�Nk}����@��<�+���a�H���5�.���]��ڪ��"M�h<��Z�Zx�<������ޜ/]� ���UY?E�+{΂�`�TԿxX����ߡ~���0�ե$��v�'v����o)�v�tec�ڑ��|����6�
ug1���n%���1�}�mC#�Y+x����̦���J�3������q�:t�ٯ+z����� � 	��jw��1oƊ8ZzVM.��/-M�Y�,{
!�t�X�\۶=�t�S�,V�f7Z-�tex������^���vÛ�g4y���������\@��1�hnѭP��5`OU����Y��������K�{%e�(T�isH�Z.�y�c$�bh'����!圬���3ޛv�V] ��W���s�vM����sL"�Ɨ����S7���ov�4��8�3�j���
�p;��y�j�;�ڙ�#�,kL�.�x
r��^�{%՗�}�v�A�6#��n�vNhϒ(>|1Dط�K��ً_p���؝^��/)�U�gs0��/t�t�q=�	��n�hfA��9x}0�z�Fj��c��"����X�x`�j�E<{v�Y�i����T�fs�Y�r+� uj,A�ފ-xՍu�f�/k_'����s�^9u�a喥�,��7��r�v������H�6��U�.q�;�4�v�ϣפ��֥��f�f�:6o-U�"�ګ%���Z�e[�;綫\�i��x5cȁ��R*]a[����9[�%�囷Z>�p�6Y�J�hV�V�p�J6˽��v�IK��ly7��w�J�яX�o*�p5k`ėf(U�v�jk(UE}y�J����ew&�ˇ����ŉ`CH�;��'�=Ip�t�:�ǯ�����Ұ���X��d�/@xqn�8 ��wuz��J0�Z��TƂ�iQ!��i��kUu3Qu�j�f^�J�ɜ.��G�፧E1��R�59��¶��t��9F��х�8|��cwY�Y�	K��x�t1rKkP�2���
ͭTp5�/[T�����#�p�-ݽzO�#���hՕ�����hW��la����m�4uf^���/�,ݱW�;oiowVxu������y�_ö�m��ƞv�zuYP�M�QH-]���E��ҥT������V�M��;�Se:��5l�r��bea���3���@k�e �n7+����t�p']���8ѱc�Цh�es,�X�W;	����i�8�wZ��+KK)õ�Պ�!���C���kH����Jxpgwx0@/�n�i�`x>}r��[��X�������v��(�V*mi�d��i)��/+�yY%#veALu�Й�����.�5��Yم�\��]:���ݜr8��k�ɻI��'���#�m��[A��C��r7�I�W�^��I̲��|�bj�؆��6�6���o	m�Wrn�aZw�Ǚ3Ѧ\~m��##�m�|c�fo@�J�{���r��Ⱦ�+V�9,�y�Be��ň
�11��z�ÂgN���)gI�T���dV��ppuz�ys\	u�>�h�\o@��3��f�Z��eQ:�ɍ�,v�d뷠��M��U留Oz
X)�n�t���TY�'f�d�Ġ�AF�M�96�u�^˲��f�c�D-�ϱT;7b
.;�!b�qt�s4g���|E�n��d��A❎���拢/	;D�Qښ�uva�&:{IQ�Z
�uq�;Z��J�f8R�4�75���g+x�&m�3Y��bN�2��9}ie�PN����:v	���g�W;Z�R'3b�=VU��.A�Db�tLٍ�������TMfz�y6-�F�b��F�xm�H�̙3r,�Y��ycl�[��t���z�Ӥ�J���Ȗ����ڕv۷������G(����S�����X;l�� �3��D:�8CǴx���t�z�wZՂm��w��<'���z��I�[)����J�B���quIV�t�R��b�y|�����,A��f\�tl�l�^�W�0�C�Mu�(ԭZ�ӑ,w(W�Da5���fM�%��Ր�nocW���S�]��\��F�ɔ�F���V�՗!Xj�s1A��s7ر���k/5J�]l���x-;���і�W����Vn�ݿV
Z�"��TVzk��񉭤60�u�LsicK��X�otҹ@�Y:���u�v���q�7�2e���vڴI#�A��MF��M�U}�G�myf�f;T^;�چ��G�E��Tzd���+�)Zr�YG:�pS��7B�f������k��E�/�c��C=f��1V6�ʄR�Y��������϶�R�<`VI׮�pV�Ubuׇt�N��!2f:�Lun\����%Z=��nL;�Ir}��x����Y�fM/r�i-6�h��[�w�Cd����S��k.�r`clLP��z�7�Z�1�&��Ng@s]���{�G3�#o~���<�Sp|S��B�k�s]M���%�]u�����ߣ�'��=�O�5y�[c9o.��^r��J�k�4+W}���2���Y�4.���:�8C�h����r���r�B;)Xx;�R��EpYs^t/71�Q��F�����n�Y�{[�q5���S�v!�<��[�@���:1��e��P�,�J����7]{�g��K����VmՋ������p,z7�p䅚eJ��᫽xȍ�0�߶���WN��t�:�Lbq橮��Ū��.D�3^�*J8�n�Ǿ-Ȥo@;ۊ)70��!����O �W�gq̽'
$����}j��2��w�,��Ek鋬kW\q�w��e����{�m��30|7�)�Y-=����-��$]jvkd��Q�%���6�����WM���ɑ���V1�3NJzc���f�c�U�_iA���YZp�aR2�V{C��M=V����z�9E�k8K�E�2�-� wA��v[x�I�Wxem�^K	{S�l�����"Թ�N��	��,�v.,�W5Py�2��u�P!$�� 8�t]+�j��E�Jރ���8� �f�77��#�*Ñ3�������z�m��Hz���ŵ���x	�pem�9NZR�z���\Q�b�V�AA�}A�"�4��6��H'MΩ�T���c�\�gU�7f<��K�d�����n��L�6�NU{�F[�������]�К�0�n:�!�b���˔�� �X���NwGVm�[r�=�3/>Rƒi*��z|.i���w&lxۋ�^b�\�6(�%�~I�=���&�l)��K܋�"���cW��GWC���/S^����F<��+��wxVo"�(q� ��;���6Lr�yk�ґ��x�[rf�d4-��w�x���l�w��e��-�a-��+���x��>�(��Z�!VԈ��dE�_��Ya�e%�fmk��UԐ���P�̪oe�5^�-�/ KRh��em��>H���{vT+���A����Һu˕��G����,P��n�
�.�4�\b�w�vk������h�}o����_���
��R�qҫ�on�p��<К@3��t��ҳes�w��� B6����	u�:ށ{�?�����m��mI��֦�� Ҿuc�.����z٘*����-�*0�j058�5]Jf�ȶ�l��J�ۧJe��������c�x!ω�s�t�s�rkQh΢�p=#���R��Bsۜ�ʡ���u�`�b�j+�ĳ\����#ٗ�����6��]U�|p�f�ճX�@+�y����G�ˡ6�������	#�>��{:�GC���GF��۪����e�7L7C7m�v=>.�b�zp�9 ����77�GvH8�p�5��ŷ����7	��^�%i�뙢�c�`�53����kns��k4�X�m�{<2;tr��0걹8���@x�g��X��n�s簦х�s��Js3)�e�m�C��U�2s��痱��ځ�˸�����;�7|���N�� ��'v鮢ۚ�ۍm59��vy�C8ފ�C����SMWRY�rʎ�2�!��bF�B�W[e�ǵ�����n]s�����sG�^�Az�l���m#���ppQ��qa���ܥ�5@�s�FU�*��������8�Ƒ:�����{�-Ep�9����t+kdH��{\At���&�]mx,����WM�f8�O�
	�nr\�Ya�K	I�3��XY<��O<�N��RI-�s�tm�T��� q��3^ŭ�V��X�SJ��2#c*Yx���n�t�pIuc��]U��� �Wq��x��Q��l�sp�ol;Jc����m�u�Q'�cm���	m=����N���s�F2v�b�W6ʧX���upp��n:β�앙i5��V3��b�ƶZ�F���q֙�.I�����6�����b�s5 ���.L��^� ݛ��ȸ��y���Y\�
�M�5�����˳���>w�a��Ѻjz���pT����C;1��k֬�y��b��ur�Vz�rI����&�a]�#u��F������g��� ��R/���:�׮N�H�.�X����9�5�����	�����"��={]�G�&�����gI�g���mn�a�ϫ�͢�Z0t&b-����[U��\��2�R�@�ZBL�-e�b��%�����g&5��c�O�ь�:$��eXC7[3v��v�*Kת����c�+�M��3�Z�Z�D��7��]����Z����/;�s���]�E�EZ�$�JؐZb�yM��3�^y� �v�]M��{��\�Y6�*{m^¬�E:�R�kT�!�5!�W���h��q���bz�S��x_]������cn{�ፏV�pBU�[ی&ܻ�yű���9Ǉ-�m>u�Up�^.�;��c�Hb��m��u�����k�C�2�a.@x��Y�����n�4S$T6j��,�&�#p��T�X�b6Rl�j�������P�NlO.�<S�F���mɍ/���5�Mc�9	+n����k��j�;��v\lDN�ۄjK��\SKk��wf3u��5j�.
M�LY��0v��A{�H��7��v�QҜv֍sǶ�e;=@�\�� ��ܽ#��-.�z^�p��mgi�ۊ���X��e�Y�-�%��!z�F�)ڱ �_mO�nfۋ8ݮ=X�oAn�y.���)�sO��틥�;d�]�<��m�	�둑��r)d�GP��ʭ�)v����������4�&��\�n�k44�)%Z��3��:@��6����Z�fj=pùn�㵢����Ui#L��meSi�fl6VC'!1���݉V�Y��Y����Zn��k$ݵ=���Z�&�J�]��їJa*�d�.�{s]V9وwnkn.��\����F�*7g�[	���3F.��B6��ƀ�r�=�k����#���L�9�:�X`�Zp�8W�-nN���Tv3�i.�{d�l��aՄ�Q^�x��f&Z�vuG
�KQ[lu#Ka���]	�"m���98��������6�e� ��FiZ��2��$�FX���z
���W(Lm㵵֯f�7�����"�9�:5��=1���S=�{2VD�\��݌I��f��GK,uSB4i4�m%\��}�_��G�� �gk��Fl]��L��sB��s,.Hy�ڷVqۀ�0��m�A�b�h��P�I��:m<MqjGu���i��ܓ�����[��[��6�!�w�a=����Ex��In#&�����sHA�״�s��EQM.�j��ᚶ[s&a�z�)��jj鹴m*��nvm��X���M4�n
mkl9e%��܈���${�=1�Ԃ��ϊ��X�[	�du4kf����K�\��7Fg��Sq���v����n����W�7�{q���jPF{AG8�'knz:v�n��
x{N㢯��Xlh�9nh��D4tlv��5:�����r�ۧ`cX��mOI1�'P;��]�C����=0��5�εF�ƨ8�ԶvoC��q�fݮխu�Nx���%vmu�d��**��8���n8���;����!���O1n�T'g�d�`�>i �{컺�����*�t����l���K�+�#�u�7 ;�a�'�SnU��%�a4�����I���յ�)��]t�K��L��i	�<v��m]�l۹���TR��z�T���ێ4CڶH���fΞ��>�a�Mݓy:�>�n��|�G�m��.�\ݎ���q�D]��xK��Y���{]:�J�*MI��-\R5��^ye��*���2�;/9(W�9�F�ؙ4FC����^�:���Uv:ke�6��.V`�,Q�����h#��,,��ݎ���LZ�t:�x=��x;G�6Fc+��2�
RR�h�kYk��-�V�8[3L���v�G]�+�r�q�9�4�v�F��Z��۰]���]��F���Ł�:��{����R�w �Ϣ�Z�3B%�%��1�m�֝��Yqψ��z:�E�ɞY�D��f-�CXX!��m2}��|W.פ=���l�n��)tX�I�J��=(��V+�Gۮ8,��эup���p�ˌ�j�c�)�{X�K45F4n��cG\��fӎϱ�oWFöR��dRx�d����q�}���}s�{t�aͷH;eql�"F����4��bu�L�ֹ��r���U�f��Ni�eR6<=,Ć��&0i�:M�$�cR��+&\<�5�eZK.BF���[H����Yn-{{:������4�\���n$�N&�X�r���B�%�]	�i/G���vZY�[���p��$���й벱;h��ۧV��V��4�x�
�6K/3b\K���.�Fq>�4c����+V�x��<�<��p�eH�Tl<��uF�����4�l��.���q�,���&[����x�݃��OY���=(bc�ٖ5Y�s���m%5ɶ�ol��B�m��������K�,eK[�Ԋ�f�Ge΂ۘ�W���k��&�p�ՔU��<W,����z�c�i6��<=���ێ'��k�{??h{黎��<뛉l����p�΃�f��j���s5lۉۃq��n��<NN���BXq�0�89���4u��`sq��DB���]{��V9{w�\���9@�!��m���g��ށ��[+U
�.t�{t��Z7<XH��4�kl/���u��({����<�x��Ù��;rė1n-�����k�N��$�8� Z�tv�\��Nw@�7jz�z*�]M �7���m�u�3f��j����9���Nf;tϠ��g6;�χBIncA�Q�H�>Xx�@��&2p��8���=}6�Y����h$�(����5h�]�2#�y��E]&(�r����c��nËu���sgn�XK��7SK��\����iB0,u��1���+���6�t�n�>F����������.5�{V.7��v���u�K��%�e���j�7H�b�:�и�v��V衦�!\܎�)�V*fI��m�(�[K�vZ��n}��7���<n�6�\��j���V��O��;#��,�5窊���`����t�R��ٛ�/�`�au
۫E`�B�i�sT1-L]����/�x٢-s�nÝ�2e�	�}�1����5�.��mu�uֻ#���ۋ�q�@(�k��+���-���}��e̫'7]׭���dMDъ���6ʪmn���/]��j�b�u��]�m�s�V�� X�퐘��7Sa�m2,�6��ecD��W�I�F]-q�ͱQ���0��-�}���,�g�@�ëa�GiM��׼��QdZq�m�i����e���ps���d�[`H�G#7D�G!�l��vd3̶����Z#痕!Et�;N�m�H�&MۧH�te�M��yĜ&i�R[c��!6���^^{�{`�&����3�ֲ�Rʳ;lu�����[�;k��'#�v��a9�ӱĦi�gi�[�a�n��'m���(9�jY���5'9�e�X�,�^��fp6�-����<��f�mi��TnM��n�p�;m��V��m����.��qmm��w�\�E<�{iΗ��k9K7yg�[�ɻ=���l��I�n��;����}���7` ��jgA1�(�^�N �t�g�S�%��\.��QXgJ��4M�{�3�[�B��ց��8�s�7Eۖ��Oq����۪ێpq�㫘xwX=��],�����ʶ1@��茻�)k��
�R:Y�7jA���M[�ѯ�}�S��r<ԆP��p=Fۙ��r��*��ڳ��w&�����O][9�ԊGd�M�L�Y��ങ!T��.�[�Y�������:����]rp3���iK�Z��M!�������Z��s��ZrZ����K��Y�ݜrv�z����j�lp�v�qu���c9��g�YN�⒝����ZeU��R��P����
�����@�u���/<�xv��Xn{	#n�q����Ys�.��v�W�f� V����F��#��Γ�q@��sL�':�#ɵ�P�a�5���S�%�f�葶�W��rg��ܷ=k�N+#p<�=7��N1㎂m��#��4�9�E�qw����<ڎf�m���� X�����4v�%hݜ!�u�N���k���V�S"5b�[{h͈M�T!�chJ�����n4zS8fx ��2��--8獇=̐��x�{�p�<;��y��v[�\��vK�+y�ӟ�]S�@����F�hZЎ��=���L���y5��ם+&���q��[X4�ۇ����)=z�v�����pf�.�!���u��c]Xm-��P��U��#�ٟ;����u㎃u�5ǜ[mA4��e`���gX��vܦ�K�N]���Ŋʁt���`#Q�ѥX��+��zMҒ7��8���.lZB�7U)����]R^k�J�k�-m/1��B��)Vī�ڭ%���U �Xѫ�%�6�@X�Ė�c(Ʋ��`Ij� [����*%�$��:ڪ����R�,,mb�)kP�s*[[W���Yj�ICs�=���!˔�)��ϑ,T�����Ŗ����Qn[3�M����s9�u��>;����G�n��N����o�ƹˇ[�o���Nu�~���a�������E�6�2�w�.oWyVɒ>�!��M�pe��B�u�l6ٮ`�D�N=����JI�n�u�̡�����>�|����������{2O'�g7�
S�|x��}�T�3����l�s}1��3.���;��˓$��g�}6�e��Ͼڬh8�2ի�MѺ��� ՇT&v �SN+�d!�i!WTn�F���e}��(fnżkN�=���܍j�`�53�w���M��Sc�Ƕ���b����V)�2�m1��fK��3t��"���z�ͻFn��;����a�0{}��Z&kxNB�QL�.Cs}�B��rzz�d��P�o��>�����<fϵ��y�l}M�ʃ��X�����/D67��y^D��!��Gn���V�M�7'�J�OQ��]'��,�N��l6�Sg3c� l�����m���U�>���_�~�?}l�o%ɛ�X�J�ѩ5����-n8+�Hw�;�В�[]���ve��onK�����{���p����]�oP�̼���l�D����w��]7��`����wP��]P[�s�Z��6)�x�1�p-<B��
��tDn��i�'u,^�o[ǥLX�q��ܩ��-�:Y%uUzIܞ_`�/U�9uR���VX�%�ح�\���hfWٙ���f��@'	������{s��r�~��P7���eK�<���*�Sm��߹�w�<�}r����u�{�����b�7��}}�>����<;]���5�(m��I0hV�	X՘-ݫ�}��J�鹖c��&�ݻ.��s~����XDF�|�*������������킓��7ܤ>�yw?D+`�����\EMN�lSn�W���>~�AQ���uݙ�̫�zN,.�]}�C2�}��wk�.�38��^�>^���R���'[� ���x��ڟt[oI�w+B���2��#r�f��l�V�=~4�-���2�=�4WxSc��6)�,�fh	�Ӕ�G�/�.���͊n�֪�r�V2U��k`v{N�^ ޞ��Aẘ�BK�Cbm�)���s��_N�Scݹ::�����ko�z�����y�c�!�� �[}��{3b}~ڿw�pޕ����W������V!N�6ߩ%[G�9��!�K�ˤ�C킛̱�W�~+��l+}�]��m�����x��Ŷ���w]%�������M����s�>H厷�����P���7�L���m�_foq���J{�!��owlU=�<�$݀��6v�WiO7�n�A�r����ۼ�eqx�e�	Ʊ�ŷ[u�s��قɻ�le`��'�s1s��C�nL�qFnmeCim��]崬�6��O쾥4�CF^iL�̥�v�G���B,�r6�µ6�9
'�no=m�[Y�j�7pu��8n�ַs����'��n���c��1��z�ȗZ�s��V�cW�tFh���l7���c��9o9wj0g�l8�qX?}�~Ƣ�ci�Eٳ�V�/X6��ʵ�a��5nh^������|����&��K����$�y�:}p�Q�}]����6M�2�s�>�-�Z���)���$���w�7�b��b�ڥ�L�t|�lSx}
�(Ư�n�O����38���e�̠�ړ�X�o_ú�����~sk������7�aRHT4����2�(�̧�J{�#��~�;�zU'����t���U��~;����"�������aR�U�ic��ι��$Xca��f@%�=������<���6*����|��^���u<��Uؕ�m�_6+zg�U8`�et;��*��Ξ�/Ex4�$�K,��
��E�[�p�Y���fE��̲~�:�]�9�����9�����_>w����ޭ�����73{8wz�m5��^����c�o�3��r�Wp���]�'�����Sc��L���O*<;�Sc���ZO���9�}^c���nT����y�a�׷_Fld��>��s�sޭ����V��c��W�}�o"��p�$���㕒��g[����k4m�4�"d٣t}�|�{�{�>����w~;����I��{Hvb��Bh���굄��B1�o}���?�3��y�e7s�����sh�{����7�][�r>�n���X��6]�é��_1qe����H��ɗg%�nkp*z�M���w���ٸ�/oce7�����$���>l}�!����7֮1�\�6>���v+u�~�k_t�����x�فky�c��7�ӻ��c���n�؟��N�~�W���T�2��+��g�˘X�u4!ƍ��n�s���l�Xb���툂=4r�;K�χ͊l{w!�}3����'�x4{��}�'T���6M�+�A���7��L}7c�<7��k����M�Cx9a��1��6*�7�X���sg�O)~βZs3�쯻s,ʦ�.�j��19�p������x������:y�w��Hj�pe��t^*���G�`g�d�'v�)�yj�v׏@�f��,����$Ӥ�5S5ؗ�y���_a���հT���T���M��=a�� �
w��=�-��?5��?Q����M�Q��#� r��f�=�[�dGV���Z�as�ݶ؆�|�ׇO�߱M�&���,~˽;��������O�N���خ�5���2�
��I�k����ݑ�4+cg�xvJ�,�����e}�C2�+3�'���Ԯ�Q��D��I���M��b�vxYط�U,.M���NY��w�y�/��j�͓�g�V����͊��7��#�m�׷�[���z`��羦�l����O|J�<Ǵf�{'�}���=g��j���65FXW|�1��w��л�ׯnvh��߷�oź�lЁ�P;k,^�*9��b�lL�m��V���雖׮�ΰX�F!�!m���!���׃.�5��Vg�Ȏs�.h���*�t�8{����9�y���C�	����#&Kn�bf�J152�v���XYF^{;:@��c'�^��MG��� �;]���F�d�<����Yj����َ�-V��d�;6X�*�J�7D�U�J�t�g�P��fIX4.��� k�������3J=U��M��c̮J�PW{�.t�p}M�^|������^�^����c�h��_6)��iP��V缠�w7ݯ��vG<��AI�lSy��m%}��?�������>� ��6���t�z�������Sb���!�qm�۪89��._Zα)9�ݔmfP�gm7�Ւ}�|>S���j�Srm�ը��\��u�e�r�-��b ��|�}���lT�ź��_���yzk�{�[��Un��y�bn�t����������t�gܲ��F��@^_��l�*(���oi�y���z�^kr�R�%�h��+_:��^��f�I���vb�d������vK��A�a��6^{)���}�c�=Տ�\��}�+�6)��y����Ł[�c��Ve	�[���y�I{��=@beHg�w�
l|���Tؼ&�*��8|M�}z'{��[&����̱�No��z�,'��R��n�ݹ�6�Vy�z����Q�ۣf����ͷ<�^�}���L�F�=J�<5�>�����yM��F�O���{ۻ����H����׼��>���tt���*�s���3�<p�9��i�/A/��B��F9��a
���;~`�G&�}ku�U)��r+�v��fɳ��Aه����G���Ԣ���@j^r=q�����e�r��F9]�ٱ�U�uY�_ 4�O�fTɗ�D�2���q^�|�@����-�6F^zm��%R��f[�c$��c:�I�SV�Y��p%Pm��H�^ڼ�r�D���sb��BE�J�
�3�ǥ����[�\o��T��ރt.����=i��[�NR�m�/��|35��o��MZ�U��$F��ۋ;X�̙y�dϞ{�!�3��~"��W�L��zi��vhz镬i���5�kF��/U��+�j͚��4^�����F@+��Wi��
����b��TOǴmͷ����<��:�4�ʶ��c��4����H�]�<�Q��k���l��U�Z���0�f'��	bl�*��\��,�x\���e<��h�CB��6n��4�Y@�ה
<(;��J=�Z�s1>����_6� �E��{����P�Y,|�wH��o��xy����7vu���י��TҴ���������7�__�5����{n���f<]3�ܬ�[����lZnu�^��o�+p����4��,"0w`f�k�����(�9x ����f�Nh��s3�*4�yMR:;���nvN|x\ՃUu��x��9��_�@wj?�xr8Y�'2��m�X��Ig�{Z�����i�`�kN6�H^�����m�J���m�	;[�:"#�n���^���l�h��Rfi8��q9��{^����n8��:=�K��e�opE-����rY7v�k�9m��:��QyY���H�����{֜��rۚ܄���������=�[w���Y�\��9e�Yԅ	��=���mY�{�f�oy�;� "��E�A�rc`N^g	'O-��М��m9]�'H�'�x؜�cL�ȉr���4�mNjO^�g��'t��{���y��ط��[71�{�*��bU��߻|f���H�O
�~�} �|޵����w{��ܽ����u��'��"��ݷ]�}��6�F,�v-�w�]�ΐ�]�YM�ia���7��~�wχ͏��<�}���^	�3²j�ly���
�Ͷ�yr��@�\�M;�}�3�J�6�L���R���_y�;�>��W�2�e}�m�/�fG��d8䧻��T��c�����u�ko4����ڸ�l�|��{Ͱ�3�ʦ7�vwU�����̯e�����]w��.rk�4�����5n>J��2��u7�`y>�G߻���>�T��W�0=����t�ǫ�:��;�;��+���͜��6﹒jU��6AZ����wv.��;&�@ԫ]@�^���HU�G렬(�����2�=m����}��b�_z9Af����������{�f��}_vP��^�ۈp��=�+�y���*#�kY[��M�nذ�̽��g���U�s��W`�����M��Jd^�t�<Q�ˇ�
lw������}�â����~u��w{��j�
�����6�E.|��<���b=��q�g�>���o$ͫ�I�Q.R

�u0Ph���v[�z��̗��_m�{#�����|V5c�1�������'���[OՈ�,����M4nf���4��u�ݻT�[�����7>�tO(�n�ŝv�[�����"����a�f\`v4��2����s��Iu����[��| �u�YŻn��u�ط��
E�.n/ix"y`B�۱���8�:���k�r>(5�tt�G>:ǒ�����:hߟ�~A�?-eu�+6i��Ժ�&.�yQ#4;FY��+(lM6�Ļ����~����:fdھ᝶*I���vۍ_��`�>l6*�qM0�݈R��&��n�Y�J���g��e[o6U��Wa��m�l|�\�d����ڝ�k��3��*���UM�laQ�[�&[����p�����}.��n]��zǲ������l6�`�ҥ]�g��ӻV�/��v�|��lSh��u���z���;�k`�|ܺ�]��r�R�\�YmҭwZ���z����v3*��f�M#��3ܝ/v�^2*rx�lU7�r�^W�ծ)�^�u��T!�g�w�w�ج�R�|�Y�
�h|�����Yz,[��(��j�V��U�S|�m�w���[�,�VL���A��> �������������+�|۾3�dC㢦��l|����/m��/�����=}�y��7�spQ�B�#�"�Z^��e��^� ^T��A��UP3��~�r=ҟ��� +�McWR4"�3�Ｙ���з�F�{����P4%UUT�
����d�����gmI㝾��� �@��wp
Z��(D�UP�X)oO<$�����z���2X\�;\k��xW���x�Qh۱I�	nT����G��w�$���� Ъ�	K
�@J�U�����S� ;�4#�����l����P�hYP���T 
��!�P
Z�{��Oz�!+�BR�.�T�Տ��zzS���jd<Ъ���{ۏO-�	��-�zJhC*�@UB�
��_��Yg�9c���<#���2,�T���]-��9���_m[Km ^���g]_X��K�Cc�]n�&����Vt�BIk{�[��o��ú�x��bK��R��r�KU%0CMP)�*�%���55�8�`F�B~�D�� K@��+�W�����;̷~@w��� �hE�_'�*}��!лp�3!��U@KB�U@)M��"X*�@�N�����6�� L�׎�O�.�Ʋ��
� ^`j�
SBvPT!-�U �����w�~9�Ӕ'׀Y�0C���+��[]�Mg�:�3��e�B1��*b?:H�	<�;�� ��:��
� ��UB���}��z��9��4#U����햃��[hC�J ��%��U 4T�%Us�}y{�7��&�]�%4!�.�'}Y�s����c� ;�&�4��@)Mf\�
�u|�t�3-���9)�4P�&�P�LT ��U@�^A��3��j��4���:k/<��B ��/4#; �T)�aU	�Z�z�u���u�U�-4!�H���6І0���ܪ�OOw�S�|�x������B>��Ǳ��;�z��
�qg��BȾw�fż6^�Cj�d�9�+�С�X�g+j`���N���s>B�� w�����@PhJ��H"F�U W���k�?�ta�����z����;��~@w��x`W �#.�hUP�!�������?/���¥� �9x@9b����U�Uʱ�Z���Ɨ��:Rݕ���$��:I��'~��+��KU$hT J��c��=1�~3��@_ <Ј���gjY��y �4.�!)aU�m	U@)=�/��ٓ����_������І��_�Uw������j�]���0��,T �{}�R�V:��@��F�0`w!
SB��D�
� ��0�����,A���C��yI���8����y�`W �h˔"ZT-l*�,�F�{����+��B�J ���ET Fv�������Π/�hKY���L���b ��hCs��������*�#BT�4*��l���#3�����{2�ӳ����^��ڀ�І����R��"F
�K@�UP����~��~#$�Me�6�����2��N^Wd
5�4Z]}���NuYc'C��r��<
�PY\��DV����'wwO����|����D����%=��Ց�6�ٹ���Pgv����k��ȝx�u人�'9�{l���M��'k��4�ƛgI���r��c���Y-���H�!s�efiwPVQ����u͎�oX���K͊�EG�UM����ٕ�p='���e��͙l��i\�i�!c�b5%u������I�гWY��(lu[[Yv�B��ݷٮ�b\���t��$��c�UzAЪ�	hCL*�>̾^wu]�|��<��!�/;3n��2y��(D�
� JhT %�U@HІ�U@)�_u�F���u��{!	Jh���z�����9~3��@W <4%��)�3;(� |�y��st�C�ۄ��-�!��B%�UB�P���e�W5�Y[���p�e���h;�#B�PT!-�P#@UB��s���[�&��� �M. ���T '����U�>Ff�j�B��@)�k�"#�ʩ�g��!z ��1�\ %�UB-T��5U(D�UP��;�׷���/�����=,�"�:��� ��坐D�*�BR0���
߻4������YC��F�ڴ"ō�䫃��.�85���뭔,1��l�]����d��/N����)hC=r *��!�*�'�ʮ�������� v�<Ў��3�o���puflhC[�� �4�U�cB����T�{[��VAy����y�� U�m���xP�Xxm�ok��_��T�,�L��{p�1A�y�����*������P���|z �hCL;�	3�|������g��c� ��ˑU ]O��g�E*�,�#B�r����"F
�K6�� ��/�ߧs;��z���"�<���y�`k!
Z���U@4!�*�#@U@HЍr�������z5xnu�*����$hT =�W=�����r޲�ۀ�BA��)����gk���Ў&��0Ch�a U@m�`UB�!�R�*����Uz��B1��j������ȼ�<��@xhC`s�
F�3.P�hUP�!�*�;{��y�_m=iT��3sN9̀ۦ4U`b��2�4��=t��6"u`�S\�#B;p�KUJF�� ��gb��׫��+3�n��eu�����cB���ª�P4!��ku����fF��s�#� HІõ	=�U{�����r޲�ۀ�B�wp�$��,T �r#�����4s�)�*�%�������KB��%%�H>��������:u���	�O��C([�Ʉd�a~���Q�ۭ߫��蚮�w6e�f��?�?��ۯߏ]�H��?S��w�q?�}�|���nl�$���� 	2�@UBؘUBXT�#3O|��� ��a۔"Sy%4
� &s����}Z�\�+3�
� 	�B�Ўw��y޵�� SB]�Z�F�0`U@)hC*���U@�5���/����F0�Bo��fkѽ����� v�<ė� �hC=r�*��`�U ���ʳܞ�p�f�L8p��ٹ������&�CSf��:tP��
�_�$}�y��B��e@"ZT#Bª}��竝�G#3�*ɡ�WL�[�`wpmyR�JhU�Z�UBXT R4P�&yw���0���u��k��A�G2 $��g�;�V��9U���ɡ���)�% U@�伭q��d %�.� V@-�!�J#B��$hC��UW~�t$�h�Ԋg���|��w@;PbKۀR��,T ��U@�T��w��w�|�9�B�І��KB����T &����k��F�31������s:�Qc�y����o`.�gC�S���3��?eR���6*����^�۴l����wĉ�d!���?c����u��k|�Oy�o;�H!���h\�)�a}���Z�
�)��PT {[ߣڌ��� [� \��>#=�{U9U��nɡ���)}�D�
� �hT 9��z�~�{���%�q�fe�ktf̵�M�)��x�V]���e�d���� ]`]� ��(D�*�Z�UBo���u���sܷ� ��y�<��s�&qL �%���B	U ��Z�T!JhD뻼}��r0օ�@І0̄�ٻ����dns3�PM	sp
SB2�@U@����z�A6�_a����І�_`��UB ��hT >ק��߫�׫~�fs��\�Vg��B�B�І_d)�U@4!����U#B4g�<ހ�`&�>ԡ4.� ��6P���r��ף{��q� �@��%�~�[=߲V�{7+�m�b���ų�8�0�Şj>���yI!y޺��e�o�})�{�o�jQ�_�{-,�8w���t��V7�G��ݽ�8Opl�L�������.(KØ&.��%����mN�so� A(Kk7z���)q�� xWA��H�,Vn�\2C�c��}�d{(l�B����s�C̂�{%�uCBzV�h��'}�,�DV��(��s�XQ�D�l�����b�&[� M�����yI����LY�����.�w�.��]�ڗ] oX�wݜ�oT�8^i��f�EzBGnf��oow6ٻ����*�:p�V*�߳n܃HT���UwGN��݀���9����#O�CІ} e%��`�u�픂���%���{�z6�R���S�E�)�k��� Y/w�o��]�]a��)m�Fi>^�l�R��S����\�>�kY�ᶫ4�@(Ɔ��8X#��u�8ۖ8_כ��d�������Ev��i�4��;�:Qc��c0�&�M.ʔs�%֞&�mYr@1��_sՕ��Ԋ�@/Xޚ/mf�Z�7�c��N�yw������@��N�]޺��q�wM�̗�e�O��>o�wQ���DZ7��>7��r�eʣ�2~�׹f������_�Y�8��B�G�Ԥ���"�6ju��Φ����_�[A*�%�wf<�s�T���c�3=+-|S���+w.j�EP�ks��+f~�-o��~N?�$��n�;��Gd��쇚��� ��)e����';{�r��Q壂8��8�-{V��n��^Xpk�4�!���^e��2*#�p$�����$�{v��//;�a��R�k^ZYX6�՜�gy�&���汯:��'Yc.į,�7;+ٽ��1�O1�@Y�(����%�ezG�p���Ѷtrm�ΰ�:��=�s��(�:6���T�ؼ�Ӱ����w�{[(����:L��z'I6�!�Y�r!8]�Yg{d8��wgu��H�N�\M���u�����JQW���yy^FV^e�k��X�q�-��ms{�z9��_����B��ҮC��G���N���w�
���B����d�Dv]�̒ĭi��CG1.���(f�̷V�=�����n:���S�/��v�$nٍ��tK��ŸQ��Gu	��l0�^m2���"�$bu��k��pWgl��s�Ecq^1Y5�Z�e�i@΀��u���d`g�э*f.�5��3Kv������2���`���32l�Y�V�<���3pk��s�������m,�X�l,Ŷ2%�l�O��R�����uxep3�<�<�{��h��b�	���sX*��K5��9��vv.��71�Z-��k���G�#c�Үq7M,ێ�!�6�u��9��;)U7�cst��as�%{ʑ"����cj��]�iDta���!@�˳������%�]�������Z���㫆V<��=`{��x yMr���K��Sv�:�z���ȓ����q� \I�k%!�b=kζ��qv� �����k���:�	-�';یMU�qLf�n�%��e�;l��R��g�8����h�»�6+���Y�x�^ø=\��b�p�j���YI�:���~7�lo��u�n�3�x��T禖p^�k�Sӹ)����m�8�r����\�F�ER��y���s�631m�e������6Ǯ�ύ۴n�c���].�bp0����=��Y�z��nܨa�<i����Aړ�غK`��8ɱ���I��unW��2���n�/�F97��1�cO\}ϥ����h�vۘ�X���Mwg���H��(rb�.-�2���"�܎Mnx��x�#=��8��g�Q�k��$14�����v1r�\�m-��ճj�(�Imo���{��l	��"�dM�p��G�N3�Mc�5v����ƵlNa5���N�;���:`X�н����p�[�[��&I�Քѧ��:߇��po��u��s�n��7�'ph�ꦸ��������Ga�9ൣ�j�q�]q�B��k,�u���;b��0-n��]�9x۞�n��5�v[��y��b8�M��������M]p�5Wh��dL̦XFR�t�]���ݰڮQ�o����{�O~��Ϟ�O�����ޓ�s�]��!�m�W!������6+~��}0q�*��jo�<�=����=��������=�p��e��}]�͓�q���^NH^w޺8���
�۞X��U/����ޝ{���#&��N����yuc����e���ἲ��N��s��v%�|��~�`�����X��ڠ���f��Y� U�rl�4[�;]!�y�ìe��Jj�M������������S�?{�w.���d��^�����{�͆�a���|�;,�xk����$�L"�E�ޡ�7�5W����+��9'1X��.Q�5r�����Y$�H��Y���k�\������Ί���'�Cj���xH�U6)��z�Bߩ���\�{lws�{{Ca�ا�ϞN�N�����T�{fOt~�ܻ�_��>{��"#�+�Uk6>l<̉�#���4`����=:nW��w�������j{v��w��]�X*��Q��'.J����]�Ǝָ�ؘB���b]�׾����=�e	q��w����&w3Ћ�+��̬��fW�����w����:�����s�I2S�۠�ŻW�xggo��|��~�a��r��-����ö����_]f)�*m!f���b��Ѧ�T�U�*�wr]�/}	�w�ʻv��+�j��wY�����k�U}�W�^'�gN�lq���2��̻Y�U���g�T�M�����Hy�^�w?}^�����܎׎����b��T�g]��IM��ů����;��s"y��n�̬���z`�[�w�.���,y6:��w7� �-���S-��t��i�m��޾|�t���̠�M�N��6M�;ㆍx�K���|
��6)�lu_�ӻ1���ό�'5�kޖ5wr���^��s���$/��Tئ�e%�}��3}#�r��6z�
���������n��h�y�ݰ����c��)B�V�ב"n�{�*�i�-��q�e{�ي����m���̈[+�b�7�L3K��^����Ez� ĝT�X�|<}|3�w߾����$_���39�.r�s�0��mj���z�R����^��*���c�l_)q����]t�6�l�F-��Ƹ;]�x�l�k��׆{n,R7f�3~��e��e绝7;�Ss%������T\�̩��|ئ�͊ԯ������}��8�����Ju}��]����<���y�{����w?7�^�H5�����]����M����]�.چT��7l��w�7:\��Ko�_��$1)#6Sb�����F��z��WT�e��ə68��:�̰3/�mՑ�pw1�+*��w~wm���gȗ8����n�ܯr����WL�S+�i�X��\^������%<GG� }�������2d���\6YL����i@�[��6�Ƹ+b�g�����[�i�c�5bd�9��ı� ���ѵ�+DޞSMr/f��XW�ۦ��ј���-�l�4�v���2���/L�q·lv����n%ô���]L6��R����q׀V�.{���c�u�Z���ߡ���Mr�\A^|R	�4�c��:-��YQɸ�����������=��{۝���v�<�{��G�;�WP�ǽBxSb�6>�$�5Y�p�ױ����)����_7Y�W��;�MK�r�ϩ����t�v ����sx��v�����ئ��ۡr��T�n�l��}3�=���s�%Џ^���T�'eÃ�syM�������९wpӟD+wc��u�����e��ٔ>�t-�����y}��ΗC.�ΠJ�.w[��Y{�F�q���.�+Eb�s��:2�̮O�Φ��;za�y͑�3��ئ���ߨgR��
��\��#���N�<fiD�B�{�'�e�S��V������ɫr�{3|��ѿ�������eA�^�y~�X��]���`��ϒ:[�yag�UA�|1��3(f;���o���.�y.��SB�Cb����^vW4Z��z��3,4�b9ΖT����㵯�![~�O�m�6>l6�ы	L�/�A��z�Ӎ{s�����̬�c�6����_��>����W\�Ƶ��cnqN�cs��]
M �Y�Yڥ��Sb��[�wd��=�0T��ɿ.�ξ�̿�(E��a�f����]���t����窎����cCb�&���]�>�)���z/s��q�Lr׫���W/:��֙Y��t��}y�x�q��Rmp���c�����v�]��(�x��<�{�5��s�7\ޯ/7�^��M�����j�k�޸+�//v���͈����'zn�b��|خoQ"�����A��M���6��C��t�|9xs�7�R�&�6����ՙC2�>�,׫��w�庳%�h�Dt����.�a�i���tx��%Uh�y���«�6*�|�c���k7���ϕ͋}��ف�|�l|ث.��Ӡ��{�����价�Sb�h��*=X+to�C��X��o)�X�����(��N|��Ӧx����|�nvZ�w�,��w�e}��ǝʽ�����JU��^�pj�o��L�ɑW1ҕ�3(��Y�6���R����mF�f�+��ξ�ޢ�xE���j���h�5��������TB��a��o�V���˦���;s�ks���F�fW��2�d�Y�燉��+��[qU=�^WMw#i͸T�al��q��-���r����1�8�:��ٷ�:��]�8eW��x6�|�d��&N�ݼ;\�;k;�n�{���yn9���31#�1�]���B`�P|ئ�Ϳ�w]�ɻ�E'��ۻ�vﾦ�}4Sa��b�w�1���]v�㯳)��{�-29�s��Ʈ��I�>�������M�����ٝGh���/5��/m�q��u���|�l�����</���3G��]���h�O�Qg�)�yڤ��?`\)��f�]���j=/�h�
�U��G���;���˒A񬩜�u�Nkh���l��p���@�j-�&R;f��1
1���l*�LCj�Z�.L�/$4Y�k�u��Ƶ����S	��I2<���[�������s�l�ƪNm��,5ƃmG�T��H.QX�^NI�4���%n����q�'��o3�k�I�)�ة�ķi��`�UH�o����~/���ޝ�W�c��zs�B�Gh�-���u����U-�������<c���ww��.S�)��>�y�a?5�}.��{��{�[*9�o��h9n�m��U��S=5}O¤I%���, �y�����*�=���w�����6�Q�<�Y�uT�ɽ{��OM��w�8)�e<~t{���vL�H~�M�����r��>=r#�G6m��h9�v���~�6ٿ~�������V��6���Yn&)8e2&{,+��L^B���]أ�Q����$2
�\#���*η�{�s�N�V�l��[����
JV���Л�wx{#����p�k}��:$	;�\G��k���J^�&�pMq���e�l��y6�{s;�� ���~��o$�l��?I��f�p}[¤�6:?6=f}-����"�I;��z�x�sW%��9�o�i�!�@n�ۺ���^4g�Tw+�/��sίn�]��8�p�HU�B�{���c��~�T��!��v�}�sZ]�mOo���ur윟��I�#WY�l���>��B��]�9�dΧ�k�@Cq��V�R����EQ
»H%b�͵�v�u߷�W�gd�6m�a|ˢ�~�����C ��Խ��u�,���]�]����;+�<q��ߗӫ��.���6&�|�8�RJ������}~4���N=���0��MG��ܞ�6m3�76�L�v�W��~[h�X�V11�ˬ�e���$��+'8�8.���U'\SfH6��K���mG�i�&+9�1�k�A�r�gK̗8n�h�=r�D����ujT�/xa���ޖ#�W��^rY��$ۀ��l�zR�quz��-��2a{C5��)����򷾵.E{��EYŐ��9�//5aA��l/Z1]+����W�(�1vn�bї�f1˱R3d��c���Ăa^�Й=uiRۧZ�����W��VAG�AZ%m�ܢ�Aj]��M���F�HgbI���˗w5��V�w��ʯ�E��Q�yg[|%��t�/ju*�1D�92��6�B��:���������=zMc�g�kg�AD�.�_X�[�@Ō� p�&P�/y��W�6i����+5׳G>���4���ɡ�w[m�E�zZz�f	�0*|��Mo0-$�X�_i���q�W��AU�_kvU��"�<&���byr��;'Z�6�Jx��N����Rv���`⸳�:;�4�,f�ѫ]]b�yv3T���zՇ�u-��s�c��XF?j���HV/e��W/w}��o36�w3h�y�]�<�k�ʓ#"釢cޣV	��9d�]��r�)̛�au���ۚ2ܙ�V�u�[�2��b��V�m�
;;�6�o|�u�2Ū��6�d4�i�b!���^ێ�㳵�<Ȝ�f�3�f���lvk=��8�����.�m��W{b�5i��F�:"譬E��"�=����[��Z(ʳ4�"��W�B\���l�'qrE�k+"�㸎C���H�ّ$����{c��e��m�ڝ�s�Qyv��N^�q�
$�.+��lq�vP%w�d&u�~E)yE�[/2�-����w��8��.c�B\�_my}������{gpwn9-�e&fi9�ێ�ﶊp���8������� ����dRs���zE@-���{�HUu��]��v�y����r�̊�������s�!5=�GCeݮ{q�o�[%��3��b�,|��e��e6>z*HdT�H�|K�`��y�X5��0����~��5�
�%�s�V����k3�͒�kMw-�3m �����b�!T��&����������3�Jnt�n�����.ޱ�Zw�!K{�5$����'�g=��x}ω�}Υ���/f�}��s�ۼs�T֍1�G�n���@��>{J���Ff��V���ۚ{��$�J{��m�F>��ܾ�f��;�(<���o��V�y�st�G]�{��2��ÈS�\Wj�6p�|��kT�RX!��c�8Wu���NC�oS�$�J3�뒲*���UA%H��d4R�����i���w=TX���E�,�x������VQ%v�v�\ll^^�G��	M퍛�������}�O<���},���Yt��s�^f��ok����I$�w�F{�G7Y�r��l��y���?o���w�_��ͷ�tS��۴7hݞ�R�A߹]��Em����jK٭�|��s��}�_n���E��7�ZΠ�ݚ���<tk��i?8�pv����H(�n���dT�I����W���ر���vT��������ICwP�U�#;�A�2����I�������ww|���R�u��9�v�&\�쨷�[6�:���uB�kfejY��I|�>��wwwN���D����`--I4��Pl[�bi����b�.�C]��V3-G�1�i���h�pm6�7�9fh^�T�+[T��S%��b�vyF'8�ˇU���-�b�z���aU��[�1%��'c�5 �ΞM�{x�2o��7��Ug�gs05j6�ݏ]tz뚸S��z�ƫٙ��	��M�~���[.��P���R�]\m%v�<l�7��Y%S�|3� ��h}��/oz2u�r�kw�^s����}�wW�H*H~�l��S��z諾�vZO�9����_n�+��{t��k�욾z>�H�U�̳q��Í7�����<�Ξ���H�I3�h�4V{�V:��^��.d�r����,y�{g|���o�T��}Rn�ݩ>}��߯!촟�s8m:���{�8l�=����($B���v����哴/U���֋2�9V�j|�<��=>��Lt���C��n��7�؟�3���}����O�P_=A#VCt!��m��}��<�4��"�@�^Rx`����/s��~�ov�y�;��n�j��Dz��]9k_N9�����q�U���E���gW�9���;1��.o��~���R �$�uM>�����U��!����k���hg[�V��;0x9&]��9�W�r���[B�t�#�����0��hո� ^ͥ����ߟ�@����}x,�(0{yY�"K�ڰCtf_}��s����|��Lɮ�����R��t�%��Y�~cڼ&���}��X��nɥj������f��j�ZM�h�`�S�44�PK+�Jww:�7����ߜdM��l]��ٯ�j(D��' � 6�Yn�n�G
0��syf��[sG�����G�2�yA���!�҂"��l�WyO��8RA Dā����#��D6�ŷaMq�o�FG�);|F_Z�������5R�����ݵmP���eI��6f_W#"Rv�{Fa�_UW�^k|�.��z�Mt���"s�X-� ��n�m�J�ۏsq��kA+!��\k��2&���������D7t�`�=���������_�B�u�9�i��X��r���2l�cn�lOgX'҂ ƾm�7C�yz��r��Q�W.���â�SL�t��ڗ.!0�Ћu�V.����Ⱦދ��0��۱a�2����ٮ�W�/ex}R� �:Ń:��_6��[��ŏP3�^7ܬD�q��ueۿ8ț��7�X ��&]��c�zrA�(��F��ĉ��Jc��X-� ��9B}�=�9�z�,-����	���"5�m}��!���yGV�k�}yC���݋}��cϺKR=i�q���/<����+�[�Yx<ۼ�&K�#���d�}���{aΘa�: ʽ�"Q˃$9����|++j��܅wrq��)���]�θ���ǹ �V���b�ۮ��Ww�YN@7��mo������:��-������.��L�j����5�q#�Cl1OWW� t�k�`�H��n���s,-����;	:�������VAm ߂�[jȥuYW��� ܁|~��X{�vS��ԑ�M��o)'!e��_��h�{H��:6�m����j�����4�|a�l��޶��ݷ]<~�Ց�A|Ci|[w�u���w�32G.�n������b�n��]�su̴V�������A�5S<�g���em N��F��X�AF�?��Y�isKӡ�#ֵ���q-� �[���뭻��yT�"��������=���[t0=��S`b0$p�}�x��+��9-���,�n��ꪯ����xYd�j�m��-i�˫�L/�ƳNDxmf�7.tAs��9ޯj�rs�XE9�-��s��<H+���Yy��3���!�Wb�,��u[�6��FJ�@*ڭ-��L����r�lݱ��O7�%..�k�Y��۰�k�Ѐ���X�n4z��ǭo`�A� y۞�{QMs�|������ݶ�fk5�s÷m��(����<�,]]]]���^�G�_����m�!��ےs�^o�#"mZtN(A� ��ŷb�źD�|���y�df�F:_��'�ێe�����>�4:�+ڧp� W�/��A�VA���6�ʹ4�?/hÞS��3��n	RG�k�o+��b�-� �[��x,{�]V�5w~�;���_nЀu{��q����2&r�ۛ�ރ�n�����e�@�[�Amؿ�uC/ey�Re�w����)#���͜,}(�h [k�m���\�w�k����E=����m�P�Z��dat�k�bn����nd4fHҺ7d_P�s9X7A�_݋q��1ޜ%9k]qg6�[�����m�<��t�mؿ���#G����QS.�f^Oz�A�㮘��L�o�FoX�^VݯP�є6�v�9�R�H%%�g.�l��nwf�y�S6�!}���:a�_Տf������zFD��x����ז���5o��w�u��Ґ ��Yn�@�[�6���Ʃ{Ҝ�u�}�u��A[Aڲh"_ �={{���&A�A|Ci|[v/��{����'#mk���yH�_�m�wA�Α��D6�X%�~m�m��'W����M��ϵԾ�{wޑ�3� ��`����׻�[OB^Z޺^���4E�#0�����3�v�ń͎4�e�M�h�N+�Bm~�%�_����0�/�%�Azo��A�p��}�!��G¶�p#҂lV?6�o�^�`�w��c|iRc��m|��%����pv�zֺz�\�u��<|ff:��3)=�łc�� ����u�#��T�`��5�]��zu�.]l�O,�~\�[C7n>��!��=����^2��mh1���㭃j�浗[���oGϟ+��n��2&~@��VA� Ch/�nł�"/ݕ=�y�Y�P~�Kd��-�W-��%¦��H����w�mװh3b�Ct������h nEt1]��޻�oqF}8?I��}��W�gX�[�A-�����r��}����%����0z�����.L�i�#-(v�b쟪��A}]{gP@�u�m` ����ȯ�ۗ�#"{�:
G��&/}� �/�nŖ���y��;jl� A]%k�Ƹ|�
�'�"�}C�?6�-���g��飝\���/��!���݃���\I��k�v���d�M���l�,�-�ͼ���u_�����yA|f�Am��ȯ�ۗ�#"{���E�����3疭'��u����mۚ����|wo'c�߳J��ܛ�}���c��z���n�z��#E�$
�Y�V���dא7ݞ�
N��4��KWq,-���ݫ�<�W&F <�(���R�f��H��P����hn�f�z�!�SM���el�c5v�ѶWQ�X7f[���«Kc� An+ ��/�m�m���۳�ٓ]7_m9U��,P�������Y���H��� �@>~��~O�������VA|���9���y�����j����o޲3].a�b�}��wV:�[v,�H�u���	�z��{tFϩp3d�$��7A����=��)�� ��"6%���b�;Ǜi����Mt�p ����
{��5�zVLu�o,� ��G��䒂��xWTo���r���뗾5v��9��������4=�._�s~��b�9�d��s��o���y�H��},Evy��}�o�����VU�mex�-=���YaW	R\z��L��	}V��@��m-����Ф��UtC�!@Xw����E�y�.U��<�f,��8<���\�P�s���R��wHֻ�ݭv��d�t��bHf��*��O��C�i�ڳKc�\��ħ��Ion��Z��j���:èu�V]Ⱦ�a;�[i��@��{Wn�BWuc���;&��	zY7`8%�a7�%ȹ��ț�2.��Y�`v��<%	B�Ǳ5¯�3�/�A��mt��P6�o
)h�:�Ҷ�������`R�!�Ed���:��B�+��}ϰ��rS�WK��'4'��9ȹ��e����s��͎�Ŭ���`�������z�!�eL;�dv[6��O8o*������-�dث��3�]�>�g��Ѹ�
h,j:�F���۔}º��7�fn�[ ��%���H�0���"���S�F��w�Q);I��wIH�0�wWʶ2��|D�8!(ٮ�F@2��J�vs�-�q���^e�v�)�.��I�7�Z�Ɇ��q7v�|Zo�]t[�!�;�Y0ݬ�e����8��˶��'����c���[��IGt�0���E루�����
��~M�l��qG�`=���y�kRy��}�{{YRTE���}��|���m8�wl�^%P�����Kx�"N�Il���n��iQd�hv��m��{���!m2�t%/v�*t�[�ަy�$�j�����V�au��K,ll�7Q�X	�c�F�Y؅�Zt����h�ˋ	
N�^�����ټ�/���x�K�h�K{PR7�R�ζJ�@���e �tw�8ɞL'�ܒ�'�Ѱ�,�[Pj��$)[�W�����g������^�[��:��ޮz5F�,w����y!Ğ��{yyr]����,����.�J�i���F4y������9$K:��eZ^��y�Z�ޗ�e�I�����n��nLљ���y�y^q�hw�_�>��2�d�W���٨���m�y�a.г
Bb!6�e��Z�_@ܜgy'��x��t��[1�R�΢QSM����b; �jgv��7��p�~���>�u���:����w6�М��޻IY�6jaZqJ A�Uc�i��bhD]˄�b�ݦ�^V�3r��L-�KX���A�tG��y��R�9�e%|vB�5��C<����>�m�$eX3�'!�ЅU�$�*:#�Gf퓣V:��[1
�
�G����"B޽��=�ܣo6�k'%Wnum��Î�Q���=\��z#�6��vL77M0O/F�9#V��3��9�f���\8�ڪ�<7��ygX����EKR�,u2��V��T� s\��lFz'/��燏�Hq�l^�{�؂MN���&Z�L���L�u�.��bLZ�����������9�nRYpfۢ[�ֺ�1�<��68w�V8��/m����ŧdI�nuW!��l�3��oZ�`],֮�6��c��C:�b�
�q��yَ������|��k�WH���A��f ���eE��������cqY�![���-�cwZy@�ZMf��8[HRJ�l��ι@qٴ�T�i��e��ԁ3)�K
��1�ź^#*�))�i�s	�8�b����y�@i�3aser�8���l�j�(FA��sn�C��}l���2��WF.���E����j��rD��K�iY���촍I�64b�[6i(���M�c�.���)�.v�@r�g<�-����k�C�Lp��p�\Z�k���3�N����We�X��$�tΗ5����T��u�o56�b݈6�6���쉋��D%�6�����%�ڻ%��N�I�>��G)SgR�i֢�ٙ���&n�B��⹘ԦLn�<xi42m1j��U&���5t���-�El ��HB���ܗ�v��C��8���Y#�mfK�2ґ����s6�Rc�컬[l[�z��ҽ�k�t�펼l@������{:���;�㛢��0�K��L�n�bư��L���|����L�m.�6-��#��Q�����ܸɪ��^ۨ$�Y��v.׫��rRck�� �Uu-�p��X�'�'X~�{�[����3�Y6�6�@�ڰC~7L��s_�b�;Ǜi��&ܚ��}���_X�[�'o�2��,ۤs.�1�D7A�W���x�{ݡm�����M}=�\���=����}Ά��۱e�_zf��ۥ�`�a�_wVAn���y�p����zN��yA&���y{�ok�<;����(�ڰCt����{}9f�Ϯ�ر���O�C6��[���{H�|����uJ��?z�l0������*�xغ���g ��3RH����,�:�: �-�[C�s�ny.Y7_u�/|k��}����0�������Yn�E�_,0�s�r�Y��r��.\�q]���`��	Bk<阳�ڔ��I5���7s\\и��Q��j�չ�[�/����|=|��sk�u ��箌���#��I��yA��-�o�����C/����|�6����-P�r�*���;�en�M�/�?k�[���������Z���܂=�hq{�i�b�ɺ���x�ڌ�]=i;�g����NK���7X �H�B�n��z��S��Af{�J����<�`����E������U�a��J���ݠ��3�p���.��X\%�s���c��-��l:J"�>�W� �A�|�z�_���v��}[����R���jx�۔�<������_ky`�[�2��Ó�me�03����)O[quw�^�����/�P�Ct:��
�w��P����Y�����|u� �tĭ֎��F�ݛ����xKUݷ��s��L$ml���71������Sl;�>��}���|f�z������w���J��ř^4�( A���ma���+�V$��KLDh	<�zи������:�6/mq�����tj��T<S�"	��/��Cu�my�u��5��ꙹ"=�+o^HD�o�X ������������S����(�4���ږ1��e���nƹf� $l*�P"��.�����n� ��T��l���й>y����|�2� �A�Y��D7Aڳ�x5?]S��J_]4>�ƽ�w�׾��8�=`��D��[�qב����C��ʫH����6�-�`��.�S����к\��󌈸 M����� Cu���b�t���L�d�����u` �[��S��l���й>y:� �P_˼*�Q(˴1#��wxP��J����ŗ�1����Mi.�^�w�/���t���f�D+Qk��*ڻ�e��|�}�k�P@����ڰCt!��/�X����ݍ�~�=��-9�^WA���}b�t��Z߫������7TE��0�&-�,�rL�m����6����Z${ә��P@�5��mY�]O8.�7�q����{i��`�4�kK��[��n�����ڹ�\�lC�� ������ʜz'�"�A��-�6=#J�s��w�@��?�����_݊ܿWO/vӾ�}�sb��{H��}7X �_6�X�8l�nj�G��;"���S�9r�s}�P�~�`����*״ƾ͈_ź@�t�-�[���kA�Z����ew^�����;��7_6˫��5>O��O�4_g�(s0�'�
�/�5�I�-<��J�*��Z�1u�;��S�v�!Ṃݾ�7�w�#�?�$��>C���-��mB��Ka�7(�v.h;�f{[mi���)��se�0���9�G.��H��V�;X۳����/+�k��1��#��.&��XT���]e�x�1K���gv�	%p��1گ-�s4�m��r����v�rpb���N4����|:ە��RR�Zj���>>���ax[�^hpc�<n��vW���!�̺ `�iV����������tA|Ch/�mر��K�参s"�W<�tk:���c�c��ź@�݁`�[���3��y��O��+�/�<����C�|�".@�{�� �D6�]Ϗ��wiAn�A�b�t� ���`�x_Ufy���ln�ڭ�is�Je2���c*��T(7����j����#�����m�s���{�X�'2/ep �{K�^b�f33�ލe A=+��t6�-���>�>b� ��|�Ur�uo�dE���V2 �!��m�j�g��$t$��b�u�Xmd�B��=��]��֌`��� ��Zk�6�=\��k���-��z6jp���|�Ǜ=�<R�]]��#6/�6�!��h^�D�]����e�,�_*��O�^AD���>멷}��^N�o/:ҮfdԲ\��L��c�h�Y���Y�<��)3٣G���Ӻߧ��o2/eq���\����9�~K�$��΀A�m� ��v�X9��uMHZ�8ȋ�'}��n�_6�_ź�6i�oP{�Ӯ� ��_R ��u߼�58�$�c�,^P@�J���ޮ�4�j�'PD7AڰA��o����^�%��zŷ��ܮ�Ox'5�mq�����"-�v,ڼw��Q��#�h�5-�J�l�&
�Kl/��u���hI[��c���_6��C�9�#�GK|�".z��[��-}�@wW�6�Yn��K�=�ٵiw��m|��]w�F�NzJ�糾�~9� ��-��a���b�^��A�'�+ ��!��6��ث��\��F�syu��B�<U%^X�J�W����T|~�\�mX�1P�T�Y�v�ʄ�D�َ�,����9���=E�Ҡ��Ճ{_!�X�[� �H�݋��i�"k����v�FsVCt��ڐu>eo�t"�;�VC��w�</4��!R���X�[�A-�۱`�XU�x,[�G�����9U:�'='ޓ���A~ւ����B��5�kl��1����\�7IvG\Eń,���Y\aj왛�Pn�l��m��n���{/w�ɭ{k�
�W�׎W���{�ŗԏ��ͼ�An���~���1Y�tWa��"D���s��2�$t"��}��!�!��l�^�{}��i}HAnŖ�~-�w��W���*��H�W='ޓ��Ne � �mY���wy��� �A|D���;�0�b��k^������M��aPpx����ς�qem�����+6�fi��ϳ�&U^���/<���o�]yW���`�XmS6���Y���5�����6�wzZWpK.�]���\i���0��K_WN�|�ܑЋ�@�wqX ��n��m��gk=�-c�\�m�[�]����.s�i�3U�(-�j�%�_^�2	��S��-� ��%��]w-����w�/*��/u�p5��}����_�@�ڰAv��r�����A|c�/��=-�/o�Z�W�� Fȅ��>y�j�x_[�R#s�X?��M��m}m�TﭜBݹQ�S���r����Ci|~m����{��xE����[�nm��}��]w�hl�-������`�������<��6�n�7Aڰ-��!�麝\^3�M�n'�>���dֽ���_n�~-�̋=��'���V�ή����s*G��$���]���Kt��I�tg+tO��%�ya���**��/�}_��:��
ʶ�qs�I�5��n�p4�]hi�g\b��\���v��u�L:f�,�n�,1۶��v-5�v�.&n�km�3BT�l��9�e"]���E�8u��z�Sp�&^D؍E@ë��5��`�mn�0Nҏij���݉�kaι�QG��0\��=�(童|㋃��
4�fhz��?+/��[����I0o�d�c/���:s�1Gk���G�y������}c+mY�T����O�Rn��!�^��J���4?/�n�n��-������T�b���w�:�����?L�zN��?o �m<9^O��� ��A}��������c��Uj�{e������� ��u��|CnŎ���U���,Gr��,�@J��9�O�Rn�����U�TOW�a����K���X-�?7H�v,�w�+�G ��J���	�Wdk�'�'X'΂��7�_���Cƚ�^���x�4ӹ�+#��9�]�5�*��r�a��3t�������K|��Cm/�mذ'�y�u�npW1�m}g�鷙u��س��E�@���`��E:����ى�����Ⱥ�c�]󥛨wX�+ۍ�];�Wom���p�����u��X�&쾺.��r�Q9u� �$0��__�Dꗕ�T��2k�*��+!����J�s.ř��?+����d[��j�����ʻ#Y2}ru�|�/�ޠ�m}a�~�ʡ���_kh����݋�u社���y=
}uw�}����?T����˔���Kt�Ŷ�y
z=炼��S�'p;�5ؕ�wج��"K�۰o��w��;(�j��bŪ�I؅��w�%��v���eKj1�Zͳ6�?�e�������Yn� �[�/����dk&O�D�o/
���T0�' �mX ����������m�vV���=:��:��w���c�mw���"�b�uY�7�V�YC���v��6����_W�A���"��|���XYa˻��k�۩�ˣ��͋�L{7O4�S��ni4)�_$�W��,�G��י#m�5���^	�O:A>�oH����U�խD������9*д�lj��Νt���+-e]�nƘ�$z/ih��47	1ʢ=�k�/m`"u��Fb�<娍�'8���3GS�܁U�e��r햶����z�eY�a���t�M;cZ칬���H����jK�G	ao[]
kU�wm��2�p��1���+����+9V#Pb�r�F[�������u��<z�U��y/r�ގ^=H3�	-�|Y�xn��wˉ:{�Q[3���ۗg-;��gVQ�T�cF(WW<Q�Q��楎�	�R�*��޹ׇ#�����癿J�W�s����,�9U�B�T\_WY�]����W	ʮ�7�7s ��P��Qp�ޔM����׬/!���H�b����"䱔^P�sd�y�/>;V4��C��3#�h2�I[eqrv�E\�{(t���Ve�mdޫ����V�@�(��Sm�vt;�T���.V��Z�.��'��h�M�Uo���&�q�J�Q������x��R����d�f-�����{	�ޱ�;{�off;��Q�6
~����Oa�o���V��e�'�u�� ��s($+MH"��PE*Np[���"����|��w�������[g�Ϛ%��Kd���Rv�A�`���%�w	���o9N ��MY�kr>���������{L��eZݻ�/�ﾞ>���+e��z�K�ḱ�Ȳ�f�a�����l���b��u�x<¯[n]�Ą���1�a���[bK!ce��^����ݖ4!:��1\ж�Q��,旅�l�sIf�f!t��TBSĞ���x��/�y�ޯ�����^�f�L��;ڳ4�����|�myE>ݯY��Y���o��ņ����8��\��{�w�{��I��^^��65v�\�mꐐ��v�s)\�{���rV7��v�Ej��Ɏ;��{V�՞���X��{�l�M��zL�����G&�!�U8�ՙ�skXR)b�.��=Ef�;������^��|�3o��k�>#=��/��9�z2>R1��:cY�HCh/�nł�}�r���{+��&KvR�.�{۬W.��̟\�p>t�Aj�yO�LVF����mXj�vjXD�k�|�,��;c�[���&��l��u��t��<������}�Ͳ�]��5�]Y���z����0v�`��m��i^��v;� �A�VA��T�T}�Mv%r��R��.w/v��[c��U�Je����)N�%��vri�X4̤A;)u罺�WvlS�>�:�e��"�R��={��eP�t��H����_݆n��ۻ]j�̾SNp���r����� �,�"	n�6��8�sͼ`�P�A���k_`m�s>��"��v%p_Ob��}����,v|R�j䉗���GX���qr{_L���oV��1Xd3��/���Y��������qz��dQ���}������|w���G���B�n����~�x����~�F*��������_�( �mX ��Mg^�Џwծ�PTV���]��R&�-ڜ>vx�h7���]�3}��}����Ѡ���?6�\��<��s�G��+��k�7�__�lYr�n����~-�Dsؗ:�O��uc��V!�	W0��r.l�bU|�ˈ!���V��(��7��ΐ�u"n��X?���Xo�3��H*�=��g�D8uC�-�Ch Ci�S�sj��tA|[v/���14�
�]{k� ��#�[ln����.R �\���An�M��k:<�v=7A�Cƶ'�.l�bW L�/�H�o�|Cn�{)�̀�fS�xo�N4�'-��f�����vX��%��V�ȳ�5t�]~Q�[�|�;�����_�����~1)���5�=i�d�n%�2ۙGHڲ�,��dmj�v����]���'o�s��N!������s4�V>tb��=�lj�Ĕ׌S�v���{O�䮘�w�:��a`5��@��e�����p��u����VE�seG=��R=�eڽu��dL�Ɲt�n1�\EP���b���S��"5&���K��U��1�f�A�(mpr��6�<��,����}���tu��4Usݐ�g�N��Z�3�ӝB|#��Ch�%����\3�����t����Yv�բgV�[�����>5;��ж4y�L���x��ł��-�`���o�����gy���I���W �f+��$@7���[����A}[uU>#B�J_-җ�{5ѭ�ޅ�|�C��A;+ii��.��-�`D� Ck�-�d7@7}Z�o=����w�y�S�uDۯm}��R�vK[���GE^WS�of��6��Wa
��wg�́띣[���i\M�86H��3�����τe�ڰCt�Ja��Z�/c��f�uϣ�uk���$_�v,�@7^�����l��݋ٚ�%wgۇ0�xF���E�z��oL	ٻәbۓv�l�S�k��%xw֫�V!�7�`�����c����C����kV~ޅ��G��J\A�V��QD������۱��n(��:|;�M���M�"�7@7L۱b�gS�c���A�VAm%)��p}j���� L�W���r��L���-�����ز�Ca/}륗����,�|ϖ�	�Aqm�!�~����_W:Q���g�ȋñ�'�M������c��J����x; @��+ �����ʹ.����;�&�{k�|���0�ZA�b����H۱`��/���j�vye����Y�.�7������<'� A���Ȁn��������6��e���_gźD6в�#�u�k7Õ��S۞��w��B����uE����-L�Y1f��/l^�3�x�[�d�.��R������jVŠ�?W��%�=��e�|ϖo�䠾!�������x/1��iD�H���݋�=�;�þ��^�� �v�:Ou׺xz����&:D6�_��_[A [io�p��oA6��ީ�$�.g��=�g�}r �m�m��G�������.�0L8#ubh�	&�l��h��T���*��3j�(}�����ϷC����#rh��������a�.�U�o�0�J��h Ci[j�U��_�G��#u���.��ɽpw�؛u�yHF�b�n���p��F*Dkw`��A��m� �k�_)�>�|$��2��=C���� ��!�����"Ig�pU�A��~�m�jld�ޭ����	�A B��I��ԎR����`���q9�]��LY�[�R�ٹIݒU���Ū�Y�3n���EL�ؽ�Wl�n0Ӽ�f\�<$�ɓþ�t�׻!w�-�d7@7��t�Ϧ@0k�/�{�gz&�{h��6D,�An����z�}{������v\Sk��2m���\���2,�*�!���F՚VP5i^����_6����L�}Ì�s-�ܾ�Y���O(f �r�m����n�ڡY�9z�{i'�䇾����>���5'�Z;⟲���2 �m?��lK)|~���~25di�A|~��{7�uFswV�u�=�ם}�� �/��> ��|�@^�]��f�x��=�}a��3�wqz{�'��O.#tK���q�P���%��` �[�Am����������<����
��;n&���G|��*��WNW͵�6�5�^��젝}��׋[V�����
���[��#=&=��j��]��I�_�j�0z�f�j>���u���ר<�$���^�(
V���1[�N��ÉҨ�e�<��Q��;�9���6ln���,]tlZ8A���c��bu�n̯=�I5��!v��Vh��f<ccZNz�	��ɵ�Ɋ�	@��N�e�:����u��ۤ������y�]�r�h����\Sg��殅�����f��E&��������ʰ�4.���L%&�T�n��aS��V\��\��ٴ3�?|^�F�m�ŷb�ʝ������^u�n;�⬫��a��A����A-���݋� F�Z�~Zj��dj�()I�N����\�r������W��)�z꾿��̤A��H�B�t�#��}u��^1��n�S�^!���m� �����smЖ�$�k-}��Gr_݋]yRs�q�=���θNz��k3��6`��&:@���%��� [h\{�=����P!m5���kS4���	������m�륲���,�	�v���
].v�%ֆܲN]؝Ƃ��/G��'� �A�b�u�-�^f6=�{�����8XU���`S��9���@A��ذ����@��VF^����%p-ɖ���;���mי�ך%��/�o�Ȩz]��Ϥ�m�㥻�t<��"�{%�{��k��#؂��ܱ\����u����G�����{>�ŵk��(x�H��b��A��m��C���嫥{B��=��m9�\𞯽<�g ��h?�t����w:���,�j���~�6�����,~ʿ�h�m?E\�.�A�U��@7�	m��_�X�]�^�-��陖,){u���{=�םq�yH��rł�#�u�g�7��Y�}�blA�&�L�����˧��nHA��j��6� �j�ÛAF��m`!��L����s�z��1�f��oW���������#�t��d"J����?)t�fgql}Gg޼C�yA҂-�v�L���@���6+!�����۰sB�ԝ>�����^�6��~1�7��Mi��S�pt����ZZ��V�TܘvY�������;3����>��S/d�O'��y\&�97_a�H�݁a�����ۺ��s�X ��.�v�Nf�<.p_zb�%R�𭮺��Dh/������7GK����V]�x�7�����ם�����-�d7Cc���ޭ�o6��1s�]��͔"��q�K��L���淋�I$�������>@7��mب�����O&y��!e�zd�xi� ��ŝ��%�_ۻ�A���N�E]4W|sb�A�!)�t�ÝF��e�J��`���o���+D��9XAe|�nŖ�KuQh��ǝӟ�Sn�|��=y�X'ҀA��Ղ��n�
���Ymz�x�j5���6�Tw�|����G^u��� G�����\<o�7Ԫ|!��M���3][/^ଇ��;Ya6�y�w7��� ѫɏ*v�� ��k�+�k���Ae"w7A��m�p+�;���W�[Yn9ٕ�̱ۚ����' �!��n�{ڋ���b�o̸�ܦ��z:D4��^�fˇ&���������]�Z~ݤA��ذ[� �K��n���}L#ם���Rb��;]C> 欆� CimY���2(�?yn �.K������o&z:� �sԁG/��ȯ�u]�P �H���!��_[h(x�ǽ��\�����x����6����Yn��n݉FR ��ř+�[�'�ۡc�ES�����x#��X3ؾ�"� ~-�Ch"[EVC�y�b��׫�l���G^u�����9b�t� �h������X�bکd�I�;nز�!���^�,�0*V�\9ċ���6��Pa�ka�H�^
w�(	��E Ӯ�U�4���HS�޵�v���e��y^��+�f�[[��I،��9W����
w��	���q��r�gݚ��R�z]ں���'Yerv��'�b@`l�1x�rz3{�����E��ݹ�-�w��2%�e�܂\+�ZD�+��r��%���[��v���F>����"��ٕ�a|� �u����nhoc�Ts�ޭM�쬉��ޘ�����E�^��l�8mlRu��,���ܵe4�`������)���x�w�T�d牫�|�Y�=W2fU�ht��VT��&��S%CPD2���zH���ڎ(_s[����rﻵu�%ϔ>�����V�;��<흻�ݘ�M��g�`�k%��g�{Ȥ�9Dᙑ�8h�j�����Cn�U�T�0�!ݥk�T
�L�F�ٴ��n�v�y���/�
��we�#�/u�ޱ�oA���_S��2B�����W�
�@���4�c��5�_kǛo�Y�y[6���j����B�a��Z�� R�˨ɫ�8u�ˉ암�݃R�o�������a+�e�->2�]:����_;%]��c�G��q��79��Me�Aep��{��os�ʓ	� kQs�9pj"X�6bͳ�EǗ���w�_/}��Y=�m������X���R���C��F#Z�9�8��)���[ąke�����3'y���;rٷ�X��䷥��I�P�z�z���RM]��W����k����_/�M�f@���m����ԋ�̐������lyn��1��ZD�m�;k{�W��Y�3	j�۷I ��K6Ӎ�����nv�k7YmU��Ъ0�� (Yj9;s�m6�����͚f�!a�m����{��γVu��;f�u���N��$�Zv���i<�{QDG6ȓ[-�ˎ��i�ͻ��z���y�Jvg&�K:qm0Yѽ�����X�.��l���̆l���ߖ�5��ǟ��<{4�CFӻ�.�
�F�n.�\و֪9�8��x�ۆ�շu�ݱ��b.<vl��sq^�r���iXf�C���ڒ��W%٬��p.��2q�e�g�%�޸܌�4lˇ3R�\�y�xΎ��.��p1e���c����c@��|��n�	㭸tr��9�r�L$��Q��5vt��+�5�A�m0]��Z��z���$�Fvv5���a5����v�T�{w���u�Y���`�Y��F��^h�j]b�F.�e��69�h����\��O.r���ʘ6Z��ʦ��]�z��1��j��l�;p�`��+Dfp.,�Zx�	���n�;TŖ1��W2�u�ٱ:�x���֪NW��mj���Gu4�NM�z���%�s�4��U̘��h�aؔx1��g�ۑ������$iK�����ը;;ir;�ZNk=��H��QR�v�0������b�F]��qv�&�⋎�tvї��1,2k($q2s�)��6�Y�q�����Jq͞��|�g���7ss��*N�m w4sYU�Ƥ�L�0"Z����Y�`��4�!������:��+)� L��
k*u��I�X�f �i�3�g'Z�������pE����F�"�,+��cv��}_ p��=���Z�n�:P���S��'O��2(裙Q���h@2���mI�7d�ln��k�2OӽsX�u��X���҃�f��T�c��lݸ��G�W���հI��I�)[��<��̼�\É�ӎ ���y�G!e�ݸ��T�٘��3i�v��ms��v���m���2'5�u����m���8�3Vh���r/,�t�ng!��K��3X��[,���V�%���9��ڽ������f,mƂݺ{T	{8�����]N�D�u/�'��1�%�
�z���p�f�\�d�c�<<-ō�̃�I��p�\��,a�_=�v'�V�b=�x�vY�ɥ�y��$�`�I�P�q�x��z'@{N�L͘ھ|�o��vLiWAeLM��<�;��;"1h�.��+(����`�A|����A�x��2�q�,zP���=n�]�R���/�ޯ�han�n�Joi���n�L�� Υ'�7Ec�ES���P@��|�W&�[^��<�@������!�`�YvO'ms=ng��u��Ԉ"97XA-�!�b�A7�<�(_�("j���6���ve@m�̱��|�|��_m�w �k�6;[���_�_7@��}�yx��-�{x��s��G�u�� ���mY�'D�ϧ��{�O�V�RiYh��&k�#��N�!FW2ͮJ�]���j���� �!�b�?s�S�5��ֺ���9{�ueX ��b��@7_6���-�@��N�Xg��_���K+h�[���{��9�TԆK���\�.T��>�. �y nީ��W3Vץ鲐x�*S$�޳�8����!i�w{*nFe�:|�}:�l�6mz��Y,Y��A2R ��[��ź~z-	���':�w	S���������m����m!���ڶ� � �|�_݋��۩ǚ����]q�}�ڻ;͛������?k��x,���@��w]`;��T2V^I����%�>@�|�}N@7_y�`m�W��;�{ˀ�7��F`8B󷝤9z��Gzw�s36�љ-��|�}����n�������t�~>��L#ל,(���@��P@��A|Ci[j����D˾s	�����,(����u5��GZ��;�@�#��t15�6�n�zK	n�������k��bW�|ʕ{&ѵ�:��m=9�gշ�ZD�Zj��ѕz�LT���_(7w���Y͝Z�l�Gz^S��*��Zkc�h�^z9�ɰD<��	����A�_݋�_�<=7<_f�}ud�s�`�_"�.��t�c݇��#ם��}�5��e���^�ώ��@ւ!�������ؙ�~��,X[���S��ƦGM��wԁ9b�-����s4��y���C�>�֦(iu�yV��R�i-�bY�td3P��jͪ�V+�+w�m"5�ma6����u��rl>A$�-�g����: �#�/�ͻ�n��K�<�κ�s;�JD\�:�M�q�p�x���`���Ŷ����UQ]wG霂fP@��� ��D6�_6��^6wu�gvc힮�-c��ֺ�״��,�|~n�m�L=����;<�=�X ��1�{�a��d�P~��|���E�8���H��9	��s~{3N�`��Ό���q�[�t��x��CO2L#�r��v��cw�e+Vp����|s�ł�"-�6���>����z���k�k�g	<E�u�{("9�E��[A�G���a�>�h�VZ��u�ج�+Y�\��+�2�A���cm�[�E4�'��o�"�� �n�A�b��d�WD��k��
�|3}����,Y�@7^���� �A�+۱s��;"��!�{9v�D���y���D6;��)���#����X9��'z�M�u��gK���s������Z��is�+�8uA��ڰAmCi�Z%��.���X ����6�]�ٳ�˓�;2:n��n���=���K��H�:�m�����_��ކ�RK�`��	��k���7�5w�瘬�����ŷc����a��G2��������2MX���s������aL�y{�e�`��bN[�6�42��O�^}y|���[e�])/f�:��Wc�v���st=x�(�D�F���כa��,'���#�tX�M�^��.��n��K���&�6ȑl[�[I�f6�����
qj�m.�؎���C��\�:����	�^c��m��3\��csf�Z՘mZfMe�\�Qx�4qsx�б���1�}�|��8hW+z��t�����Ƭ��N�4`Re���\�;�_d���4�"	n�V^=j�g��W�gW����:�3�����Am ߐ?ڰG����:/�v�X�;���;�]��������2:n�~7)�b�t�\�U��g�2��wr{�"͠�m���kמ��~����P7�5w� A���"r�/�mذ[��i/ՙ��_gr�H��8��Vp�.x�y��� 󻺽��Q���{b�A�n�����"eUÞ�����T���~��v1̎��?\��D0�HAn�Ug��$�Β�7�9�;�ݍ�����!�ֲ�j;L�쩈w���	��#�m|��{g]�odjX�C*OZ3�m:Qq�_�/�k���@\����{�N��܌aJ"'l���"�O1�t3}��^�{����-Z�z^�o��i�m�B�_RY�'5��.#~���*��w�@y�Ⱦ�+׍��s�k��*�����t-���*�LB����y���mCu��go,+�v�o8rB�1̒����nW�"t��w��s�n�A;h {��A��ǲ{g_{���%���\���A�pY�ǻ�Yn� ��[w�t����C+/$`��=����hp>t�m�К'{����Ϛ��6V������%�YӀj΍����7f�6��T��ؾa}�U�F��A|~mػ���w�d��p"�����:S+�1�c�A����n� ���X촴��,w+ Ȃ3'�.��Al�K�qy��"uCpٶ�ڨ�u=��t�����{��B�tu��K�Mdu^5N�0voR��Ÿ���Er�4ѐ��l��I^�Bͅw�.��>�j=��EؙU�;�*�nY�������k��*�_�t�E�����A��r�oj�A|�#�_�v,\~΂gs��$Z���ܤF��-�q���M���<� �m���Am[i�=�r�n��� /��waHL�X����`�9 �|�C�u�S�]W���m�e����)4�ú�9�N�d��l�hP61��_<���w���+/g���k��*�Xʞ|=�ܪ���w�E�_7Cm/�j�C잡��1����|�-�Oo�~�j��mf�m�5��;���)����DN�/�"h/�mY�������oC�{�z�e$I,Op@��_[���?���`"��۰mܡ��金��/���-���3ͳ���OW8X?m> y�k;��Xf�� �~:Fz��A].X��R�(��e�g5��G0;#*lG7���S:�
��B+�wa�AvW�i�,q��`��m ~-�`�� Cy�����o��ao_���|/K�"�\n�Cd����^ؽ+�U3@�tF�iu�eE����W*h����nq��Z�D(������)��*�牍]�+��aQ�÷a��=�z��w����6��+��������� A��^���e��p���G�!+3;������*�X?mA��m��_`�܂>K��h�� ۱�}o̮�n�C�>��H�WA�_!�X�� �xۿ�l9���k���b�7�#�/���ue���÷c�y�=�w1|�m{��ł/P_5���-�!���뺱M>.n��տmw{c೧��M"��A��D�k���>m}��S$~c.��h�n�L��+Ɩ<{��;V��C�^�����rJIe�Wr����X���x��Wm��i�0���
Ŗm��./'X�(Ʊ�؋-�:���LG6�8lOO+���w^�6��vK���"��FXb�v�-�:9��������{n�h⮏���~܎�p�ڄ�<�8<s���Л����vq�N���m�`�ny1���^^y.�2�6q�uv�Y�֏<�&��+.&�BK�ef�7[ѧT�q�1��~E���ݮ��Z2�V�gYtѤ��f���Y�n��T�X�	��%���C>!����q�:�xm��"�\CFq�~s�;������"w`�t#s������nh�\j�P]Ypn��oo��hL�	����C}�46��S���g��u��ί�h`-�?7U�_�?5LU�{�t�7�W�X'�A|A��mY6�!���{���Y��7_&݅����{�l?H���	�H�i����1� �R!�b�n� ��-�]U3���lIf�Μ6���bg/�1X�@7�-�y���?_�ߏ�����1�p�!���������P����W8y6�m]ػ7yZA9���_7L@-�9��/:f7�V41�e�$��tn��q}a�t<[jȤ9J���玑�@O_����|��z��_S��S��v򁒮�<2���z���ӯZǃ��4׌>�6�MF��݋�~Ζd�a�F�W�m�#dB�u�[i\n��H��b����"�__͡�;vH��T�8�L�[;�Y"�]������X"J�/�h_źDV����_]ͱ`�H�n�����w�k��+_}`�}��eU�zT��E���!������@��]xt���.�[�g\o��#[+��"�,X-� ���;ҟ/Ȃw�Dݕf�*�P��-ɓC�Q	ݸ6���x)`�H��Bʫ�pOt��<� GJ����hq��rNw��bg|���T���㸟�� ��6�Yn��[�A7�c�)sC"2T>�����Mw4�և적��@�Ի��aoo��Y��OP�w�@��}m��m/�m�χ�O�}��+/�<�YQ��iYL;�}��i9�8��Ĺq��ˤ�ef��:42���6C�:/�e\(U4,��yHf	����� moZy�cG��$�8��M����ƶ��g6-������']!<�)ݏ���n����2\��f1���u�{�i[v�ޣ!l�f�Zl��"�I\�!���1�)Q�MV�D��Dܬ_�vr���X!z�r�l6�)D
�M�g1y�bmڷ3,��$�u5i�g1��fAC
�1U;{�N=��F���&��F��vX&�Z�k�z����ô������t��Xt�ts�	�ڰ����ĺ��&ۡk����Ń��yw�T����z�$�%�u�d�{t������&�9)�d?�-{gQ�c�;��N�% W��ʔ���Dz���4����CU��-�#jN��^~��:˫�~��5ktHh겠�o���v�3�i�`q
�r��8/&S��hO&m �Rы-e�{;76��'��K��Jǧ��9ٯ�����Bv4l�3*�q�¸���-�ϖ����r���XM���]�b����b֧@�DΟ�{��Y��{0U2��Cud?M-]U��%g�SGk~�a��8�p�y�ǰ�\���U�º�,l���o]6�@����oxu�z��wd�p�4(%ӱ_;&қ%���0�[=i�]�  >��r�?���4�+e�{Yq�h˛m�9f��v��g�����眵�oK-��͵�=�K��]m�Ύ^����stX���dNݶ��r�ݶ��i�w�Y�X���e�(�')jKB�8��͍�%) �e$���ڵ�m�(E��S�{�م��۔m�-6�m�춷�ye���Z3���'I�����f��{n�{nY�y�i�!$��k" ��j������󒽛P3�� ��7�v���{{�Y����fnvbme�f�۬�f۽�咆ɫj�m���q��9�h��q�3l���m�h�ē�ù������Y�!gjq-�4�m7	mg��f�r��~�p7�6��ml��n�@l�,�H��n�!�b�6�Jݠ��ު�.PGdV-��,cvN7����}���&�w�^*��P��kC�n���"nł�_�m��{�+g�j���{��\dV����!�ڿ�n��YY׆G�9�[Զ����Z���A�_VG#N�x��u���r`X�Sj��v��~{ߞ:�'�X����6�X��b�$����m9]���'s�3�}���gz� �[�Cm|���"�%��������R�68xe��<�M���d� Cf��wp%*�^y{+ ��,�K�-�H��JsNnww{ݙ%�Ek�{(/�!�m���~B��Nͭ�d�D��݋��tpya�6����n�2mĲn��z�(����,�$�⼓6����+Ƽ$����F��䝆�CQ3z��t�:1^�7&�p΃w��	�-� ��D6�� �Am|�J�̞�7>������<߄����D7_ ۱�Ο�o޾����|a��R[t�n�b���Yodrt��m�U[(]�hU
H�n��Η��`�HAz܋���Ig�q�}�;������FP�;h ������_6Ղ+Ԍ�=����Ge|�wX���΂N,?Fӕ�n�Q�[�I�{MV.ӡ��q.P@�h"�W��=w�/��o��9�)�O�o|����� ���m�`�H�+�Q��;zŞ�D�)�67����FCM>��-�ʺc�\�}������-�d���S�8�F��z�v��18JyN�i����H�����Ku���9W���~��ƍ�&��l����$ij��ֹ�I�Mv��]Gw*xkd�]�6�r����%�>��>��Z_X-D�{!HFV�q������t�KW%s�0�Bz;����vgCn�G�a�z&]y�щ��%ĳ=a˹Rqco'۬������3��l4ں!�֡Yk�Cl�@q�R�ǆ���rr{k�q��=Si�jS9��#n����qV�0�Yq�';c>z8��ֺ�ʅ�cB��V�����~���`趼MnxPi)A�$5E�����-@����C����4�ܠ��-�������6I��ׂ'�*�B��*�;Ԭ�:�w$���ѧw	|[�Bg���U��ݣA�~��Y���_M�2hq�PlA [j�CG|`\�z%D�@�[j������s��T��74w��\m9\A��G,Yn��wb�/o�IA���1������6l�R������}���/k�Z1u��_�ł�#�t���t�6���NV,](�6��_=�2|,��� �6 �mX �����p�R���V�U]�h��v1�7T�ӻnt؛�iK��0�������~��/O�Cu�m؉1�p�1���+��;�{*R��V֑�hX;ԁ��B�n�";u�/;��(�y�wY�ߒ�ߵֺ�>*��)�Wj^�ס�n���Ĭ���{Awr��in�����UG*�>t8�V	���{8E�x"z&������"���گ�^��]ѡ�,i�bS��wq,i��Ӗ��������lc��b���X'�A�-�`�A����j��{3�Ղ���۱�1�p�1���+���� �^7����CNe A:���X%�[A�8{4�4���Ax9�"�<=y}��\A�_۱�����Q��6�Y�����L��\�-�zk�Y�W!j���~s��ϳn�n���t�lo����b���=6�/hBƂ/yY�~��m���;읗�c#�f�f��#:X�PvA�e9��jJ���"o�Yn��/�_3����'�Z��hi�`��]�)�ܫ���������&��c�=ػF�Ю�\ۧ "�U�˯i:���LLo���6sۆ�!\��N��i���$��OD�}������_6в�}�f{�0ʝ��r:�L���Kt��,��x߯�jB}`���}���16���t=�m����dy���^�:��m�z�q=&]�ԕ�����[�%��n�'����Eٻ�m��L\��Y�2�kd�)`��k�F�vI�a�&���-�� � �-����=p9�p���Kz&��v�6{ʱabe}����}��H���@���hz�Z�j���
�s�ܪ�{�Ԅ4���@!�[i�cr���mF��<ڲh Cu�m��g�9�C��}��2L���+�&��M���a��@���9��n�Gn������جCk�s�/1���M��<�	�_+�ޱ��V%۷�PX�C0�\�43�o��l��[Z����r�26p�[x���|���xj��<n2*���C��\�VWe]���%۱e��$5�N>K����߫�{#���X'r�[͵��B�<t=���z}��7ӳvֳ�hk-Qc��=�u�:���9x1��6�E+��_j��Ct�6�ŷ`�r�d�w#RW�޿��0wWۑ�"-�ͼ�Kt�v!��}��VAm\k�%�<މ��qYPD7x�wvw���ľ�XA�D۱e��|[��:�ۂ���n{�w�HCQr� �A|[j�!����v�]'�/1t���A�_݋�s���=RV܍I\~�H�׷��ל}~B���:�6в�#Z�L��^�RT7�h#�Ms����'�ӂ�qYP�/�ͻ2����ޡ�[wZ)7�pb�m�Oq�Z�s���sᰝv�t^����4ӱW2#��N=��c��5侣���l]�'��n�l�6|��b���t��"���Ӌ��'%���m�ѽ=d�Zv���nsa�H:�ײ�͇`�'Íᶄp��[�L �ڮ:���[��M�&wQ��&��O�OC��&9�#^:�ⳙ��+��m.�1�����NX˵�{Cv���ճU�b��K�����.W���ݎzJ��X1p�Ԕe�{m�i� �kR�����gr[�%�^�{��z�}�*B�Z����("�}���~@�ڲ3�|����| #�_M��e>�.R5%p ��Ho�Yn��X��5x�]";��c��!��ma6�B^�-K/ll�8G�܅=���ˈ2 ���۱`�H���\�Պ�U`������	n�����=w����5����ֆ�)��Ϻ�p����ww:LwrH˵s5+e��`W\�8S�T���r� ��,���'�e��5�SJ�*�E,�q�I[H�Ƌ"3 �hbt4��]��ϒ���X@�_6�Ch e���g�f�x&r�����P����7����Yn�����C�H�˽�t)u���1f��n����LȔ闝���5��q�0�p�*/����]'���y���������s���jw���<�E��_��B#�郱���������-�疃��f_�,-�削MRW| ܤ-�����|�ϬAz|&����NA���~mP8��n��&p@��V�nm�.V��F����`�H�t��,�W��4*44�R�q��~W5�3!"^PDh [j� ����{�IA�W��!�46�Yj��;A��%�+s�lS�B��`��������y�ϐ_A|[v.����>�1I�J�/ᛳps7��|?;yY~�n���$_e]�*�L�%��q���^+l���7c��Mɡ߄�sج@�6�v��������R6���-֍��y]�^_��zNɞ���lIi�ϖ�����w�pQ�-�� �C����t"�o!�9�]�s	r��k..��^����EI��/(/��Aڲh"����u.�h��ܠ�q�m�2��ũbd��%p ������箽����@�u�����%��ͯ�j�pz.�o�9|2s��Mɡ߄�_g�X ��"����^~��aPV�}b�ٯ����z�������!+V�$�I����S���kv,�@-׺����{������=R/V�� A�A {b�m��	m� ���{-\�V�!����X���>��L�2������k�[��꧑��/��w`�d��!��Ղm��<�vQ+2��2#7&�~;�	�b�Gu��m-�y˚iV����UJ�b�X�����[�س5��_����w�Wz���� ��XM�h�c4���f-3w�B}Sh`���A]Yz�]�����%��Z։vh�t��%ۯW��VA �m Am� ��=��r��
�˸�	O_oz�=�ϳ�I\?�� �������������0���}�Ɠk�]�X��u��i-�	@+.����5�tE���x�X �P	����n�����7&�~�e���UI���܀ۿ��?7H��\�Q�9�1JDҦR�|����z������y[jg���w�e��"4�V�D6�ŷb�_zx���m�{�����o*:���|���/��|�u�o>�mo�]��Gu|��|n����d��M�=9�b��~�ۣ���0�ݯ�}��u�t�-�[�bx�f��Ԧ�xi����}'+���<s�|'}A~�A�H�B���Z/���h�up��O�N�m�9���,��:+MK܁���]"�@gF�eG��Z�C�w��uùJ�ٜ�����h]6���K�l�`(mF�w�bUH4�h�g0�����VqK9&D8wr�B�-����cZ���*�X�DQ�/zȏ�&
Տ��.&T�]�K�S���<�s��u#���+-e�`WxH���o0�K�8��E��Y�C[s�ݼ�S�ް3:i��Y V���.ԳIGm���B�Y����U�vk���s�����4r�f�}NS��^�9;;|���Y���Dt��G�_{)����7Xɹ�)��m�mi����f��R ��̍�OQ��e)I�P�sWoKȵ5o�X�K��qP� �O2ξ&��c��TV&����6e��<3�%P����V�t�������i�F��ޚ�0�7�� ��=W�wd̋h�X���j6�7���`�ei��]5�A����ZN�4�=�&�C����6�r�2�7׸6����H�QC�G�3)�m�����Q�q��G*ấ8�����R��O��OxmGӰ��!g�6�6X�}�S����Y��q�
�7�B�|�WR���˔JC���(�嵏o���=����n����44^ˡ��9,��\p�l��� ���I��F��6�7��m$�%�cga��l�F���Y�*�2�$��8��c��f�^���Z'cX��;!"�r[A��j�Yd���Y$c����x��X�ZhOmkkj�Kl�	�!���fR�/=Q��3�����{bq�y�r=��Ԋs�G=���FڎL�{v�s��Ĺ�X]��Qz�{u�W���XI���/2Q�p[e��h��ѵ��ٰ;�=�B�Ҵ�m���ox�O&ݘ�5�C-,l��!�A�9)gjI��Z&����Y��y��E)�ۓ�{tۥ���v[�0���f�)�$rt�,^d��ɶ��p��]�m�rY��Շ�aD"t��{�&���ߙ�~�o�L������;���vMƥ��Z/[!�4y��M�q�7s�A7[�^z���v�#mEM(n:�nnǏ+��g���5n��%u��q�c� �fڅ�W[����Q'g��r�����Y�kQ��:�9������m���γ΃�]79Mrs&�n;f�L�8�Mf�]"��ku�ۗ��]5%W���p�Wvѕ�����x9��'����|n��%�7K�B��А�&r��kV�s��c&í�( JZ.��l1��bS@M+�`YB3m�v����/����\q{��F�iu�ǎ4Ft�Ⲁ��\QXb��.��:��ۛ����2�� ��*�x�k�)[-!cl��\�V�i�ns�����kŇ�0��C��ۈ�5�qLu����RV,hbW�\�jm���y��M�uM�0���c5���Y{������\�7f�ۆk\Lf�cq�����Wq�Pۊ㜖�9�.����VM��n�M�4��m�(Py�	�t�KK/��V�u9������x�]]Rv��Kc\��2�[	��Q��8)竁�l�o�8p�e�f.����XMu�XK�,-��[�p�-ƹ�8��N�7cM�^�8{BԆMӷf�TV�uix`-�n���
����LY��9�\�icH:B;8�&�X�8Ճ�9�Y��-�ӄ��6�Ġ4]��1�M�G0`���2�n3[3XZ%��a��,b,#WQ�s [�v�^�}�z�M�	�F�fB���;A�ы�ݙ�(�k���KZx��>�'*6��;3����eЁw �8�%��cj�6���/e��f��:-s5�g�n%f�RѮ+7Cq\ Y�.�7Gq��u�*�h;e�n�ڭ��D�9�o-���7W۳K��ƫ�g��f����r� �[�ۋ��
�٢��A�:ZG����wCk)K�t9���7�N���!�/���I��۲'�`l�k����� �L���f�c�����v7)���玸oBǌ�s���`�V:��f���������l8�G!�kl3�n��X��졻J��MԸsM>��te����z����P}ps�]�&�ʎ���sc|�ܒG܉cTJU24ꠑ�^�wrڂ�HȾ��=8l��~ٜꑾn��
����s��Y$��GȹHwPGv�Gv�[���{��mH�����IO6}o��}A{P_���n���5殰��Aւ#v�[�>��wMWpɷ2��?\�����mW��e{��"FUJ���	ʩ%:��x�yS*��g_���8��4?N=p�xL���x�H��!���%�b���xV9X`
W��T�
KE�av�kX��uЉq�������n�����ݥ� ��A�9��_d��ϭ�]�a��(+O|�hh/�@j��CU �W 7SϤ×���hǕkE��*t!5�B��rD"��~f,�b�M%��q�w���ْQO'q��]�	�K$(�&��=2�g���4�}��wg+�.ę� ���"5��we�u{ ��DgP@��ۨ � #uJ��%.�u��=^����N���3��D����A�_}5j��V�����Ar�e{��v����e�{$�͟[�	�P�S�ZY��F�5�!U���U�UI#*����ssڨAs���Ϋ�u2�Tu�n��Gv���f�j�^E"�RDUe��	V�0�l֔��K�D�B�
�if�]<�#-������ ��<���ۜ6+���g|����u�~sj�ڂ��h/���� ��5u���N�����>ې�ߵw��훛>�C��� ����q�bƪW�v+]	W�H�䒮�YUU�UPeʎ��t�7 �t7h�<��F���3�bi7��vs�Ѥ7���\+�_��g>��oE-�vN�qN���\;GޫP��4~�������{�<�^�XAւ9��uy��S�6+���g A�R"��Wk�}sY�d8�_�uQ#UQ#��U��u�h��.j&�;nv{��7����� N��ڂ;��?n�ex�aN�|;��$�i
��PGB�͎�e�h��l�ud	���R������-���Ϭl�ǟ��ޜd�qW�/�G_R�2��wk^ޫEmX#�A|_R ��H��۴�Ι��ߥ����"����s��\��	���R9�>U��{�Jg�Ưt} �W 5uw ��ݍ�vQ��<�}����{g��w�v��k���
�\�B��A �%��)ޜd�qW�/�G\'�_@�Iy!>�C�[|��"4#֔k׺���Lg�����`����J�@�*�,%�\B�ʝ��oS�围=���5yK��Ms�)�RH�U5RK���zk�9��8mˉ��g A�R��������AP�v�fߏ�$�
�`�Bq���<�Ϟ�]���v7kٲ�Sb�������~ ��}�^��B_�$��K�7����X�2ߍṱ͡���A)|F��H�H�h��}�3.������Bu�2{�W�^/J���������p(��%32ee�,aU$���IsC�����rέ�=�nz'�	��=Hg ��K�7PGv���Y;�����G�"v��r>��]�^{g��w�}A�Jx�At�Z��'v�Ẃ��ө�a�A���4;�as�
���zTu���F�;��?��ט�ٗ�I`�+1b�~�����VW{��k�rhW`�
Ӟ�
>��e���<vvʪ��;��ʿ��ڴ�# �nf��ckP���7:��S����Քq�!��hx,sa̖�lPձ�n�m���Al��P�6�
����&R��.n&e���,�`Ve�@07nͺ�΋�x�rsQ�+��͍��	Il�MՎN��L�u����ZmE��[W*��fM�n�7J�:��S\�߳�����J�a�t̪��a��Qf�ui[J*]���)+���W�{���#_l
��rԇ���˳R�~�5he�>���c��U��R7 7Wr�Oq=��m|�ڞ�q����6g�}o� �"�_nי�}ީ�^�دP� A�A|�K��Vv�G������ao�^+�q��1���#��}����X���P�/�#�HwP_�R�q���jU�W����ȴ��Xkn��=?H>W ��~�?dɿMJF�S���Y�L�#2l�HE���]�#�K��C;)s�po�#\ʻ���ib�ڢ�!����Pֻ'0]v:nQMfc�i����=e��d��\��u:zq�ӂ�t�+�}�߽/����؎|�$y�)��D��I��S!�S��(�I5}��if���K��=z��|��ֆ[�;�TAe��ns]f�!���W�V\�k=�����^�-lv��[���xL���H��|�#w��xy�]��̈/��Dd�ݠ���\yuEWI%�3'���M�rn�ˡ��uQ#*��UI+�6��jdz�B�/�~_n�BON2{���C��q����/5�{\��h��� �t��A}�A.CG��/kݳ-:�g�y�'v_�N��|&rz�@>A��۴+�ѷa{���ϙ.�
`-mv�-uL�lV�v频�۲h��VѰ�>[LKt� �_nׁ�M�v;�u�.B-�Bm����B���#u�Awk�6�ud�5c���������'����Y�q�)�-����DL0|�/��A�} �AO�#9;�o]X�q�q�j3YnWLb�2��^e��xmGp<>͗=��F�1�S���P�q	}E3]�wv��&c�l��8�ȫ���դ>;�F�B~��� WJ�I���䗨}�t_n׾ ��\�K��&\�^��}A	�y�}�ͫ��/�"4��"������ϜM}UCG�ݣ�����Y�}��)k����wh������=|5�{%}�n�,]+MV�52�����fi�7j�M�(�_V�@��q���"�@ߖ�;���N=�Us�yv�́��D��|wP@�@�wi���ϻ�~~�%� �w�uNY]&e�G��'}Aj�r����XUA<�]�>2?UԄ� ���{�}~���>�6d��"̹q�	�R#A�@�wi7PB����(	�4r�[�#�y����ױG��g�ޤ��Z��7��ʥ���K��f���Ք�?i���nӰ�ºn�_�VC��k-���R���݊�1!�_��A����|kqN�)O�*�Ǿ�zv*}3�B=��;���_n���C����G�<Ow��ЫHX�$�ghR�u4r�*�M���5�3l��SM�{��σ,����v�}��;�isȷ.\u�+���^�
�䫨�ƝTK*�F�	e]�;TcY��JD��3��S�<z������z��w���C-}�/��#% A:��A�H��C���p"VW���<�ng��=�8��@����#v�n�(�U�/�c=Y���#9/�ۨ)��wm.{���_p>�D<u���]u�^P�/� �R#uv�_n��ݪپ���P��=��[���弾�:=���%�R�:�8!r�3{x*^���l4�͏[b����)��":{v2\ǢZ�x�{���m��ޣY�A$	�2�����iۻ~!oBlm�C��7�9�Ih;g&���FQ�n$A�R.{p��j����n�8r�\k��N`8��6�q+��1\'�܌�n
:��c��ǮE��)m��s�mOGi�.�L�;4�C�ɓJ�qZ4C=��9��;l<l���GG������w����nI�ih���3jm����������ln���ɑ���v�Ԁ�M��^����2Y��7��/�ѩ�Owy&�=������P�Ϫ��w�1�۴<F�wiWן�,�_IA};�ӻ���Kܹq����F�ݭv��DL���xHӬ��UJ���2��6�������~�=�#�<��K���Ծ#u}�@ͅ4Q��5��������s��wy-s=��U�Q����9[�IR�!�pѺ�������5RN޺�iO�0ԍ{�9��u�����Reʪ����Є��p�|�|�������l��� X2 ^�AjKjXڏ���=� ��s)�P.�������|��S٭:n�fvB��S��U��A����PɹS�<�ydˊ�þX�ؼ��]E�����i��&��w;e��A��U������Ѹ�U��;GZ��N�!����V��Q:����Dڂ;����fj�$oP�/��"�4n�'�w�h�5���ݷ�d��5�����,a�*�6��%�S#�ŷ���P@���9)7h/���E޸;<��v'��7(qT�n�Z>lm�܀�]Hh��kة���}�=ܻ8�;ڭ�dN�����ݥ�5c)�g��رeXUEYT�Z�#E�6���wU��u��1* ��W4�{�e��l��e�x���);:�����̹q��%}��*T���g �u A;���Awh#�ۂ��c>�#mo)����:��Ž��r�z���C��J���R�y��:6�rIO��ˍ�eT��
���ޢ�&����� ����9�֖����]�����z�W5��7+e���b]:�k���uï3��d�B_7R!N,̠Dݳ&��������w�&��:������>��vv���	��J�ȶ^J������iˮ�xim����C�.�|�>{�[�g�X�����Ӡ��$��CЍy�7f��֊�6�.y֌����6����N���퍶�����T�����X��� f�ϰc�M�����<A6��uq��U����'O�jm3;nj�{���-��i��N�ײs�0Nefg>.z�a�ol�x��Z���c��ͬ�� �B;����9��~,����?c����;�^r����T��\֍��.�n�ei<�� {t�;[� +������x������uGo����� ͼ��F j�7ev%ݸ�ٷ����*S.+�ޥ� ʷ��s&���j溫�R!Y��;�Ε�V�5���Є;�0� gs��\�jm�mq�t�Kj��Ձ�j�(��߾(B5�Cjx�c{�X�DԒȬ��7��l�ժb0z�z��E�m3[HnB`��S��4���v
�S����P݆��*�m�=a�S�y-l�dT<ߍ����$�[��������
֞�����C�3YH�p�5ó/ZK��-��F�U��D1�H<)ٻM��6��l����W���r	�i�m�hA���'[�gyۡH�AI�r�',f�X�ɵ�kF�s������n�ٻD��yyk4K,�5����w��E{dfw�m�ݹٸ�^Xm�mYh�L� [b�L�{N�%�w���f�׊�{���x�h�n�ݻ<�JQ�6mVyވ�Ķ�+2h��^�pV�̒r�X2��{֧��"m�������Xے�6���z��Y�8�i�jI痬���A+(�/J�Oc�:&^z��;{�������D�J� Q�5�k@ -kH��i	:�-mm�n��nө�kkvv�M�V�̘��e�v�A�5��w�t&d�6J'�l�1��i��p��&�8M��_K9����*nJ�)|�3������IeT2fej'ԈyA5��u;���ή����\u��K��=IﶧX�o����>�Q���Q���5�K�p-��$��N��8�;�"8 M�����v��qQ�ݍ��u��%P5d�F]�=[���.��]`���n��l8�e�_��,�ϧ>�=�׈ ��z��Gw{S����� ���s
{�@`�}%x��v��� B�K���'�g���<�u���R㯻�}��2/�h{���@�����C��Q���4n@j��}^���g���dK}u������R � �ݯ�ۨ wi5��Y��A_u�;���S�����C7�@��P_��VKB����KiWZ��0�AZM6|^�~���^p�]���X�D�Ov��������WmjY��[�{��
�}+*B�r7U
j��ʭ\:cÊ�jI�vuwa�/v�)sk� ��2 �;�� ��o�f^���Q+hҳV#V-R�1qK6Uԣ���jHG65�i[��e�쌳�� wi�_nK�_g�Y��Q	�5�ʛ����i�t�����H�"5s�u��<_WȽ��v�w��z��Fo M��#��WZݢ:�� �7��`�"F2�IeT�h��5U������~|=Y"�{U�զ>=ƍ\�X�T*��K������ ������ڪ��̗ד�㞆 ��&�H	�=4o}܆��M]�.�$cTH�U$��&os�mx��{Kڻ���]��Fo7�y��k���S�S���nY^�n���%�jM~�F��*#����{P�g�{�y[�,��N��*v��O�QU�d>�3fLUxEa h�����j��St]����v�bx��q�g��7[sri,\kp�y�4�<Q���	�
��[�!]��3�"^��Ѭ��:�*���Z,\f3��4�kc���M��9覹`zr���=8�uu��2ݭ캴t�U��\klC�'�^�.���	8��������r0�X�,˴������WJ&�<5�%�3���*�U��.��_=�3+��A�OJ��:�E��>{y:����$>�����܂YU$��A#^FE�����O���4ܙ�u��>���x	�Rڨ�H�[�_ �����u ���Հwj�O6<1:�[�p.�<%錌�K\��B���AC*����/y���ѾA}�+�7P];����}1K�_p0j�q����z��:�/��j����#���W۴�ȥ����=�$8���O{��=�o�ߩ~�@n�}�CB}zϣ����=˪]���K�P3����+Hs1bЅé��G�,����|c|�l��)ڣlR���[1��� �{j/V�u�q}�%�D���IC*��UVS��3w����^�+��t���[T�g�.�wk�r?����ʗ#�b��r��=��n�n\3��V���7��;������eK�]�e/�?H~�z��yT*�|zc7�-x�"j���;�/��|�PWZ�z�$5�o����L��x7�oԈ v�����_n׏Ʈ�ǲ붟���|�8����Ͱ��
:�Fo7������'�W�+��$���UeT�ʬ�=���Ԉoo�=�ي{e}�e}%��|d&����&U�u�"�^]g��
\����Zb�V%"�E��̅�nw��'���2����xz�Q��f�T]��L��o��Ȱ����Q�y�$g{
j��U1�U��Y3u�t�J����lR���l�hf����E��}�;,%3�U�9�"3&F�"F5U!U�)��L���M�U�w��6��j+g��x̚�<]���Z]6��vd�
w�7i���ݳ�l��k�f��Y��"���~������#��<���?{)%�";���
�^!��꡿n�uw��+�;����n�W\A�����[�y`h_�7 7��R7 ˍ��O�\�~�==�׼Ǩ��9�_��?w�*�Ϛ��φ��y��+�&+���M�,��q�.�;j<���Mc��i��̲���x��<y����C�諂�<����b��j��ʪ�c2����S:��UI*�	˝��SB��̤APGe�ʝ��OG�x7� M��Π7Gw�ؗ+4����|�u"7h wi~;���^�������6䭡�� A�PP�ݤA�� �Y���ұz�e` �D�۴��򞎸�}����ߨL�Kq̹�x��,�D� �de�����-<w�fn�ir}[�2�d:���p,�']Nm�"SBk�����5W[�v�#v�;�+�w��생��&�)�'�|��@���#u��)ʒ��qv��U@�I�@�h_;nݤm7b-{Re��Y��Urٮ�\b�1��}������ywiAݥ����3:���3H���u`��̸m]^C�p�AR�C��J@�c-?`x��������:��>�yv��C�]v�7 �a]���o`K�ҙ��f䕗���GU1�I�eS�W�t�y�ޥ=��o�@�~���{�7k�+��*�^�3e��W�~�
���JByv��-^��7x ~;��|'�{�����|A�A F�@��D�P���6z}Y�o�8'����O)���WUi��G�	W�+�tT9�!A��$U�Ռը�
�K�]��l�'��SN��+D4@���ʝ
�$���џ|��_~}��h����y��i�Va�[[vI��!�df0ۭ M�lk`�4�-�m=��*�]C�\oN��n9Nf�qJ�����0���z��Kp��8ɸt���+s4���� Y����Ԗ٤rnk�!�î4��z�QYM+h�s�6����%�Ƽ��irM�p�c�tm,I��RS-)�b�������tY7�㕱�V٘J��h:9���v��E�q���\��A�۵�7h#�����Lɂx7BA���=�*�Z|�����uwk��ݤFt�u�jx����?nҶ���;^�9dn�@��}"�D����5�I�P[3�Jʅ%T�2�?_�!�jsO ���S}����G�h�]]�>=�����AQ��丙^���[����yi=����Ɂ�7���}�~�E�ߐDM_/��#�HA���!�W u�8����ZeK8��lr�����1��_m��A�wi�S��i��������m�0ꔘ��U�+3u��U[T�+Ű�W�J鼟�������<��瞣��!����|��d�S#�#�}.��ӳ�x+���pUH>�|~�Q��-~�˟�;�,��t�׫zV��/ȬF�oʳ=�@pK+Լ��C�+ep������8�P�fR �A���go%=��o���H_ ��[Y�8�/�}r�=Ծ ��Dn�۵�~ݣ���wvj�=�7��~�q������D�;��T��UL�V\ݽ�2�Y˒Y�$�7P].t��˩VI�2:����!W�:NQ���M�9ԁ���_ N�#uwj��g�V//�A۝U����s�o�&�K�P@�����1�1�Ϟ~��(��6��昻mf�.���]������T�KL�؆}z>�,��/Ϗy��u��՞�#�kޚq������{ԝv���1�D������È��\K�:�J�|��)=s#�?&����ӂd����*�p�W�Q���|d����= �mb�X���G�ё_.&Ï+��Ҡɢ�Wq����[6|/U}ܳ`���� mtV�,J��#8sJ�	�8�]ηw���x�y^�oR\�GzZʥ©�l�t���ĺ^ʝ'�
�#:/o��|)�د�3	�y��=��v��ל�'q�ۓ.G����Y�eY�DЪ�tB��>�d8/t&��ƍ���n����Y��p��p��l6+Ӳp�<Nws���ץ	j�W�ϩ`�U6�}M��<�r�Ob��b�{�=�=�״�7{�꒾�}����.ޯ��u�ݪ)z��5�����o������C���m�<���jt�����|�7��uVN޻�&���`wXޕi���<����w���Cy����T�cTTab�29�W����^.Hk��{\���Il[7�y:�w��en�7M�uiuM�l|ئ��nk�@S�����ȟ��N��j�o�����Ɏr��uW1�݇MՋ�K��]��;'X^���W���Xs�(�̡�elw�/'��&H�<��ky�UV!�Sm�͊W�^�wU|�J[_ISe�����I����vevw�{�Q]��}���m�6��:<�lU��3��#^�Bt~��:
l}M��I!�T�g����Ovt��0�>��ڊ������1����͆�͆���I��������UDU������0�@^s�\��?q��}��/��`�z۫������wW@!�~�B����c|_ȈMF�QQ�d��F��|5��A��$�1 ���/�0$�7D�z �!�l>8_k)B�mBQ���0 B���0����x���G=������/�����O�&�P�H���,��G�I��v�I��M��-V @B��;����~�����B@B�0b�� �/�ք�!)?���~���>���/�p������̇������K�@8>�ށ !
����+��m���� ���F_����������F�G�:�D~3�o���ч��>�7o��W���D�c�?��@@By��ɏ�G� @B���A"OM���F�QM(����e�m/����@�����9�#��Q������@w�
Ѡ�k�/�K���K�?�(?���������B �-�*a9K��.}�����A���5�����%u(���?O��9�~+��>il�/�}��??C������T}'� Bо�N�������?��]�����TA�#���_$��Bӕ� @B��� L���h���	|�Z��C�+(�@#���N󔐀B��-�4���*G��?�,_'I$�B[ [(b_Q��b���{�>L8d!��Ѓk����5-�7�W!�� !b��~��?\����������蘇�/���h���|�>;�> ������D�??���B�}�a#��z_o��y��>�O��_��� �������>o�7��BK������ @B���ß�v��o��g������=GЏ��'�?_��sh��	J ���0���������������?00k����o�~��.JY����~+����͆~__և?(��q3����F/�����H���r>�6��(ؗ���X������Ŀ����_S�K�#�U���$$ �/�_Q���C�8o����ℬh7S�J��vq!���A��@���/|�/��ܑN$=���