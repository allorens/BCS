BZh91AY&SY~<G���߀@q����� ����b@�P   _{�2�(�e-�����eM�U �Ѭ�ڑ��"P-����Р�&�-�"�@�b��M�A�h���TV���Q��KO�@�e�m�Q����U��-��f�ʶ6�eLڶ�j��Skj���
�Z-���mmX��eV����Z���[mm��#l�25�R�5��yڹ������m`�60*l+M�ш�[iek4[[j�H�[�i��Z��B�iP��MA��2�m�*&ћVfjՖhhY�%[f�MnZ��VMml�m_   �}U�X�ڪU��f�V���S��T(wY�u���J�v�q�Wj����4ݙN��:)Aq�
ꕭ_o{m�k`0�6��*YfƢ+�  �>t�h��V�T���5I
�Ș�
Sup�AU��\�((�v;J  9��ά�+���[�4U>��ؕi4-k3C*լ-��m|  _�P��sp�
U8��^�@U���N� 0��=P7���)T9�{�(=�׻ݵAB�{�{��
 �:��� (i�Z����@�h��ٙ� ��z(�w�熇G���U���������>��)[�{� (
w�ϼ�ʅ){���TIJ�[�*��K�gA@�wN��(�hr��Z��l�kZ����mXl� �0{m�S��ҔZ��B��f��Nt)N�Q9���S��)�R���]������h t���Z �\B��wtjE�����B������ 6� �;�j�hP7k� �&��P�vۃ� �j�PD�r:�M+����
;�\)BJ�S�誠���z�5l͌lil6b�m�  nv��@)L�@;�`���Y* 
�ӻ�%(P�U�

`���[�;@
YC���eu� �v�Vͭ���6�����   ]� ��q�@
7.� h�c��47u\ h�  ӎ  L�� �� ] ��i�*�I����JiVYg�  �P�\ 6� ,���wSp (s9� �  v& ��,+Em&( [ף
$�E���Eeb�"��  u� 	�\W@ܗk� Χ  -ڸ�Q� v ۭ\ ��  lS*�U>|   � S eJT�0 d0� Oh���P   hh ���S�@     �O��%RP      �I�&L�&Dz�SѠѐb�OT�~�% M  b  q�9q��ˌ��x���9`�#6�sK�U���l��i�h�)��ɇ3�)�  U�* 
�  "����c���%UTW�T˩� �ÿ
�ڪ�+����Um��+�k��j���ϗN�uB	0�Ճ�
XD�`R���+_Ś��k_�m��5L���{�k������6����Ͷ�-~eosZ�-�3j�-�sZ�-�sZ�-�r��W�j��k�ֽ�k�-�r��+^��k^��[�6׹���k�ֽ͵�kܶ��kܶ��o���[^���m�r��[^���׹��͵�[̪�5�sZ�*��kܵ{��r���W�j�*�7��{�׹�{��sZ�5�r��5��j�ͫܮͷ�j�+^���{�k�ڭ��Z��Z�U�����m��͵���k[�6ַ�V��+Z��j�������^歭�U��6�[ܶ�����ܶ���շ�mk}e�r�k{�[osmk{��o�֫{�m��j�{��or�[ܶ����ͭ��V���k[��ս�U��mmor�m�j�osmk{��_�k��m��[[�֭�ʵ������Z��-m��kU{�Z�U{����[m��j�ܵ��ͭ��+m���U���{��e��ֽ�׹Z�6�sj�+^���Z�ʿY��V�-^���6�sj�5�r�{�osj��{��sm{����{�׹Z�-�r�{�or�Yj�6׹k{��*U�ф8�~�(g��6@��7S0p4�ymZZO�Y��=m���·Ն�;�����q��f���zt��ҖK8E�;LT�2�x  ]ڰ9'N;�f���F�b�m^�+�	�-��Av&�B�2�2���]K}ltiz���]�B+��Ѽ�)Z�{ե����l��]5!��d�O�F��o�Ǣ;���:
��,;iPL^��J���C+�i��nB��aP(���[�wm����d�v{nnΏ�*���,���I�q�Z��dbb̤1���6��]ݼGF4 4�ZQM��J9z��C��qCpub,J9|��^T��fl\��8{��C��G4�����D+3���#�O�ȏ'L�
-��P�7p-���tj�T�8��,��v6ª�F���>���ٸUw���u�cy���T���&�״�)��qq���a#��a��7M�D7���ڂ3�D[�XN!Ϩ�]���i�y�\�λx3l��Cc�^�kA��i"E�J�b�0��)��K/�yD�{z(��T�U�]�!	�qM!k飡ǝ裷h��&*�u�+�f��t��j�J�㼅s���O(;#0��ξ�A�����6ŀ���煩݆\�6�`˩�KA;�[���k}7Y�dΫH�5�$vDu���	����p�ޣ;5n)�[TE�9N�%�R���6��ʩ�[��NV)��]�X�$�����WGY���%�[e�q0wv�7���&,���ZyK4��s5●M�
���\N�ǭ,��9z�L*��4Y���b�J x�Sv��gQ�vV�nh��յ(�+n�fb �z�B�g� n��uɶ҉�݁f�sfQ��d�4�q���e돮隮��a�2�]�n�=n�{l�{м���Y�՜��6�_i�����a �����xW	��9T�8hr+6[�!݄j;��E��^��`��mS/\ �wXZ������*P;&�Hm5���x!��v�D��}ql�7k5�	XL����*L��9Xtjڛ����ɹ�0�E��hv���ĭ=e� ��c��u.U�,��uM2e1$���mkPf�ź8\G&�#�!�y(�2�vS6O����v���i8q�x��r͜�������y7K�$�yuZ�*�Y\|��We�y����'��꬀�ӥ�A�v�8��ٝgZ��y�z���,�l�gԡF�ܴ��gkS�H*k�$��q�+U
Y�r8t}۹a��b(0�Z[���k�@�[�M<$ݣ��4M��\:ےj��o����G�>��9�`�ۄG������dש8�P�3E�R���J��A�ю��"8�Ql�௩�Z�H1�(��A]ug4��.�F�,�Vգq��w7��β�_^����v�I�>]��b}�3Ǽ6��O�b��ڔ{�#{��g7�8Nΐ���yZ���o:c�u��25�X����n���:tn�~ �ou跸 ���ضL�]�1[���E.����1�qb�b�K�b�yA��9Ȉ�6��#of�Q	`,d����5��t�@��[�@��{#ݗu1�7V�#Yӷ�XI}ð�V�9��rn��M��^���`��	�6K&Z]��a�x�ќMӶ�ޤ��Y4�Y�mPy���ڎ)������`}�� �sڊ@��yW�0�Nm��K�f��v�����ɯXݸ8Q��PT�B�"�f�ö�ׁ�ݰͭ�#�LZס]kt(�`���=��ɇwe/gQLL�Z�am̭v���4(�#i��s]:���3���WY,qt}7��p���4��iAN�	bܑ�5V��N^eލD���y�]0���d;�4����ר'��~-�0wL��n9L:IG V^ɇAO뻝Y���A���_v�va�[6��)Oc� �P�W�6����;e�.x`��^$W�U�b��F&�5�3 �ӷ��D�F��nF�snC�j�*�D�Q�&�W���e��_��Xl��j	����s\�e��΋؄%���;C^�t�����S���y���ӽ0W'SL{}X��s2��{�_��aI����6��LpIV)n�aw4hYyR�ZMq�i']�c;�>\-2�ekC�gy�os2-�c�ʛajs��sd�Ι�ܧ��gHv�)7:⸕��/&&�|U���Q3q����rs��z7���E��
�<�Ԧ��e[�r+a��?�`F�D2�\������o������w"�I�MJh�S,f��\4*�����̪ζ�oqS|L?�!��4o2F\��jFQ���bz�1IX�8V�ɗ�2�H:��[��e:)�il��]V�
�0B#�$X*6U�̳]�]� #��Νt����>t=#�C{ �Ƌ�Y�"�ٽW)nZ�BF.]���Xq���-�LU��8k��T�KE:�8E��Fig���ѽ�U�"q.�L�ڱ�И��Uz�	ͺ���(鸥;ǚQe݂��;��M+*�V���؎��v������X46e���X�G�? �s1��T6��ܾ��U��̈́oQ�ې������kƞ��I�fUˑɞ����H�J+2���7�%�h8��z_]�fX�+z5g2�	�n��>�/�-��ك
pS5��#��;$�u�j�e�=�sq�d�j>�,�+��Z��'��7.�L��J5D�D%k)����N�ͪ X�]�5�/n(�+l��!"���*4>�ܺn�r���S;yu�1��)�يl�J�PlDp"�A�=���0�;���jda9��Bh���h�����M�-&�� �+�^�������ǎ�$5.[۴�j�G!-0d�mk4hŉ�����t`9F�fVX"�cP��qٔ�'2�.�@�u)c���oY�ǁ�f�{Jύ:���(��d��qP�q�<�JB�n�:D"'������fj���%��vڥ�flf�8��ds�P��]��1�!�8�{����Cw��fκ[�zl��ƈjX�&嶝vh�����N�̅�ٱ��@Z�1�L�pw�I�vs��f �[�Gv�#u�ǋx5˜�BE��w�p�0m�uf��.$������*�1��/3����4Fv��i屔,�t��L G`��ӆ�<��;��Zޟ-a�P�]n�+��f�|³K��E<�7 �s)�i�gj�Q*���@wt�1��=�QD�7�Z��� 2�`���;��3'�"�$ec�3)��+qو���]]�e�r���{Z!@㡴AҒ�����`�*f�^Ѧ�8��n�1�����;OoKNsbM�s�rI�@Rx�v�����u��h��Qv�su]���8ݏA�K�.�5��Y��1�8]3yn�����z/HV)�y�5H �G}o��K{`]�;rM�u�\�&]�L������sv��M��X�%�i�X��Zsj;nn���qaТɵ����;n°��^�K���ጬk'6���0�!��MY�ۻ�!���lf�[^ �"a�.�.@�,E_kC�Rփ�Xvl�XW;�i�)ƬwbX$�5k�.�Yf�}ϙ=z^�2���7s��eS�T�cB,���l�i�t�Q���]8s0w�k���*И����hNYj�`�c��K��p�Γ�e�{ ����h���-{��c��:u|�����Y�.�Ĺ�Op��E��q֞�q��,f�\�nN5ٺ�\s�W�޵Dv��7�{�@@X2;�e����UtQ�*��U�g�$Ȱ.���-]Ʈ�f�Զ���x��[	�U��J�����D���O]��=��	�7�wI��YI�uq|��tX����dnE�� ܳ,d����8�פ$漱pnj�N�͆	�Ty�O0�Té6�1?H�n]�/�$�+��v�!Z6q�y��U��n�T��a�D��P��i3Ot%��׫��5j�+Pb�c�f��g�]�ˡ�i[򉝨D��%�w	��kM��|$��M�b#@I��@ᗁ�&VE"죑��7l�1S����A����R���]��BCg��F�.�R����Py��a�dQ��3״��-�_9�_���S�ux��������aש�5ig��֯ͺt�H`�ŵ�Wen�	�쫲�z����;yp�cCG������r=R�F�qz�7���V����xP�y�w`����F�L��0&���b���@GN���Ci�UL�,�RٍT1jYZ�sB���10�GT�;�!UV��\����܊eܩ�"����hy���oݺ^ݲ4���1F_��,�GLR���d#�ðkUe�U�r�j��"U$R
���'6�h�83�6�]����jz�svc�C�3h�6�%����`$�c��ඍI��\,/ω���U�����s�k�Qؙ��S�i/��X ��G��4�1��C�b
i��Y�囀V�>��x'l�ݪ��k��퇙�Bԃ�M{�{��:\�7WY���zQ��Kְ��nm�F��t9Օ���r���9.�L�B���vY�<�(���K�s�5j�_v�~継�o�A�P�b�%���i��,k绌�4-G��Ğ�3]���Ep��#�.FflBV9��7"$�{���Jl�,0}m�i�y�bج�G�ЎW*?&��C� �h��'1�M��\�������>����L�Ⲍ\��l�N�L6��NÖ�c) �5YZC*E]]Cc���bR�7u�x��멘���S�֩s��^����ԭ�6d�vE�2%�"٠"�ŗH�6�8&�����Ṽ/���j�����S��<G�.�Ѩ����d�y̷����\O
������{3{��!ʣ]p���6�-�w4&�M��ї�7z?�'�-�jMo%͘��m��<%��8$4=�p����ے"#�m%��iΝ�ӛ�oR��c��\�>t�s6)
��İ����ڙ{�b5�[Z��Y.�z=�U��ڤ��FC�����04��9�ʢa룾�7�M��Ʃ5��nD�wWW<�k�)��2��u�\>�GIZ��w%M�';�-+�!��p�
bѳC�eb�e���
�Qf��ֲ�@p�۳/�a���^JyN��	IejSd��:�Z#gՇ\�Rnl�ʝz���9�w3��G{4��sh.���Xh���
kQn���Z�*�J�B�bs]��VP���g[ۡ)��d�U`o ��*�7�gp[8���g+v<R���ѽ�B9V�MXc���:lKv,�E��.�Y�� Nv=�ÝҪ����{��@����+�����&[�e�	bw<#�?o��u�B���c-;��X�H�6��;Qȩ���+�û��XsDqG)納8@����
�n�ӗ{iCa��#e���%�]��aW����Z�6j�C����ٸ�|�d�����R�ToE�8ꣻ�z��t]�%�"��b��*�w�]��M�]�&n.ѐܜduq4�a��c�UD�`��F��ݽ-	�ѽ�t!wi<��C�����7	�cMVN1��|���ȃ�ژ��qW��:�_ht�9���d/�$�7[��˧fd�p⼭e��&ФG��Q%.י�?4�L3rzÇ�w}y���F�<0<0+��Q�pe�������,WGh�X��w��ݧO�庵f^S+hP�x�y�E�f؆Κ�Y�ܾ�Ә�Tάۈ�G���غ�ر�2�S{{oIz��{�}59r������ψ���k�\�@Q���5�f�Jmލ=��}�(���du��:�nH%����x�0Y�'%@�n��I�1�(N��Z�Ѐ�`�a��o��s�¡s��8vk���D"�"�M�N�!�:2��k.��y�$��G!�jA��Ib��E�[��On�1�KԵ�%����̼��
��!�0֮��ل�,�FMBr�6�1J���j4�����K;��(wX���g��,�?zW��e��V����&޺� �Fj�i��5h�ON��s�����[�� `��LI��)�tzw�V�FOS��壵u�/^(;������s�](]IS&�4hVZ$FJW`����cӗ��luNe6f��'�CA
ov��-+uzF13Pn	͋~}����#�B�Č�c�:Ae�#�k�Z�Hcj�:��]�
-Ilrm�qU��"�CUl����Θ�"��f���&J�u-n-�wKKw^c��Q������;j[e$�HD(���	.FnY՛[�N�������(!���K��n
]�����H�RJ+zd� �.�գ�;/CTY`�sE�Y��Kv��]0��{�홧x
�$L�M]7Zҥ[���F���'�|���.�0��@�.�fv�����$o^(�R���@�͌R��X�0i1�t/2&���6�ݕ26̎[��EB^���2L�hou�����v��iW���l��r=z.#�5F�����J�s����djޗP4H�r� Si��:2|I0���`[O���w�<4�!�n��yi�q���������k�xG�zC��&ٛ��F�4���;M|u���s|m�樧 �f�WG��|��8�w;������˃~�1���xM1����⿉C����1q[�IIr�`�M��)n��;�8<�����Q��Yrq��k�#uCB̕`ǮdZ��r�h�f�4l�kiB���o�q������^�E)c�:��|/E���7����?䚾og��=*��K/������8���	���u5���I)���9�ǋ��Ϗ'�����{����>z�>gW'r)Mڜ�Z�� �T���N���wb�hf��R9Rj�k1�%��@�d� )p�ᇋ��{}�����`]��0KnA��x3uI��tn<�/DOo^t�`�4����Yz�t�V])X���L�W %m`�n�#b.�r,�1zxB�z-���n�Ca쇍B��[1�7������Dcm�7��f �K���W
�؛.[�/�9�������h��'$-�ۤO!����$�@��}K�w���gmY��X8*&�L\O �r�֬jm��(��XbJs�Q�/�W<|�9�k�0E�V������rW#��-�׶L����4�Ȗ��i�I<��ȫXٗ�Z�-Wuo�	3����|L���������V�h���i5�W:vJ�C��n�!���C�;�r���	��9�"�,5���h'BǙG<����2iݱ똫��R�P��VF@p�e���r�szwma&�ú�*ϻ��]�ip�/�4��-�7��#�z&x�ʽ�����xOĊD�m���Qx*���r�'j�X8E|8�3쉚��<X%��.�w�F��X�
��v*���.���6�)˔�VA�T=�X��Q��:դ���e�~�д��1_q�f{�b�Xxk�;�8oU�r�暸�^��{y����Z~A�s|׫��k�Mr[e�q���:��8��F���m����z��"Ϲ��
UP2=�B{��ܐM�!܁�×G��r�M�5����趲�X�〥�̓w�{ �*c1\E4m�
��=/$�:�{�yM�k�	��YV�����ܹ�g���3-M�W"`�Л��Lv�Շ�
�J�Rh��][l��J�9����2Z�vb�W�R˔��`�;[���5�o&���ݱ�6�O�!c%���v�M�*���T�^�7
��𻵏w.���J�v���VޥK���w���Um�sm#�S�{�?L���r0׭�;����=�'�㻝����|v�"쯕�7�U�bZ��G���/��i�O�g�Z�l��D:\u�M8�aAɚ&�H��t����-���k9`ˁ��<�G3{$EJj�����3lV6�sVr'���1d�{��0�1v�ag�-�:��|�5x��˸:ml7��uZQ�y�H��U4�ﴄ�cP�{��� xמVpf�v��8�>��yeÍ��K�d�o��Os�y�����Z����:��n��x �v#9(3���.h�ޮ�B�][��p��x�Y7{;��K��on���f�{���N���J�e�š����tgz����O*��.��YK�/e��:'�x�A��ۈ��WL�,��Ϗ6�h�.fs˥tyD��6���|��hv�#����8�/�oNK��o D�_����D��={�2hW����~g��^<����ȹ[�9�j����X��}b���QLR���C���y��c�.@z!�l/<�#�}��yw%�%.�XcU��xxŬ蚮�����KvI�hd��K��}��nd3��8��p�ܑ8=A�fn�ѷ��tpġf�r�|�KV�u�AR��6@+�᭭�:�Sgx:�{����&��G9OyS�;б��ZM�2��/�ǌ�=��@4^�|�<�{��a�m�c���(�����/yl�I�Ղ��p봇���y���5Gs@�V(�i�����z:f
��(Ж%:zm�V�.�&j$7;K�7<7��q��L���}�����bW$2�C�X2ޑW��P�(Ga��'�)�9��UbӉ/�P<mC�������'w���q��j|�I�m�sfŴ�-��L��t�{���I�xN�tvAv�}}OQ]�{:nn���m���*��w�]�ڱcA�&��S��G([qf�3��p�s�UF�V\ĮW%�w5a%�ys8iR� 9XDb5�N�dЈ�`�h�����?~S��'��t���RO®K��ҫ�\�r-�2���p5���o��NMmlN㻺]cH��,
Ă*�nڣ:�r+�PE�e��^bj��A�&�Q�ڽ̒n̽�U�}ճ/�j���i�����M�_!	�;GJ�nq��m��a
�Y��0=S�}�E��Y�Է����x������=.M�ZEr�5����5���*s�t�t@́Vέ�1M:����w0N��B�@��=�=ϯwm���0l�Q�T+s��L��N��}G>���Ӽ�R��RN>
����1#=��\aB#/e�6���ӁCllV����Y�';��'�Q����c�~[%\��v�89����>��z�#X�`�m��y}+0"k�����(���%�m�kPڃ���<��}�5�{����a֡��Ƣ�0e�#��L�ou>�������t�	8�S(9	lwD�:�B��jJ�:(#v��e�Ͻ��=�:ٵ���h�t�ou"��=}2͚k�E+q�Y����@�{��@e���38:!R�DY/i3��q���`D���@DY���s�n_ �B�����{F<������4��Q���������MpݎsH�}C��t������o�_��LLU��07�H��wJ~�t�b{�7��ۨ�7��mp��5-� +}+Xͻi��+��-1��T}1\|g��cO��U�n{Y{�^���9!}��_4�G_��<�u�u���c�ZT�2:�p����oC���ͼ��A����n$]��Ðb�m���Ν�3��3mՎYìr_YJ�4��J(�]�	RMw,xr�mQj�{���T����m��E���W[tͳ� �.AX�]�Yf�{|�Þ�)�/V=�#��ȩ�$s�o�Yj����y��ۧ�}: |���y���`��wf�u�n��#W�2=T�7ӹ�n�QA�YX�]w��j�t��j�v�!6*���g�̀'���*��������c�塣�r��z�r�P� �6r���^��w��8�s�6������ϴ
|9�H�O%�Lp���sf�3�&�z�vl�6y��p`�[�ub��܊L�[�]����F����@��z$�Ms���k���8�VcgS�1L�E�D���5kK����;��`Ih�EE�ղ��܄\[ƍ��]1&�8���#;3a5��b�� ����æ�/��PSL~���������u��SO�$�aH��W�ȑ���M�� ���P�{I�O1ue&:@�#t�OU�-f�$��U+�Ґ����se�L�(�.p��t����r���t����Zv��T�l���#j�l3h�1Wωum�\���`�S��`��e~�(�������M�X7w���%���3�������)#�g!�[�P�pl �kz��T�����[
qf��=�O$������:��8?6M����Âɫ���4�;��{����m|P�,��&���i6Os�� i��Ki9V�qaf�cN0Z�6ok�%.�K�TK�tm�gVЅ�:�a���AJ�Ѩ�[5k�며J�X��{6��q��=R��ݏ J��뗴��u��j�UiC����O�¸V�y��� i�!��\��M��ܻ�缬=�%���CQ^���i��g{�3�f��`���(�ݜ4U��N��=pI�ʄ f�mU�Y���.q��&�Ԕ�4[x�+��;Ӥ�$�C��X��;I�����$��٪�d�bd}}�������P�vL�M�Z��g��{�v��:3B=����O�.��بizO(7�4��u�+��$��Fyw�����%������5�cb�=�D��ܣͩ����l�{�s���q��^YW�K8�}oo*T<ho_-�o��d��Z�'�i��u;g���ϻ�D��|����&����~����:#�'6~���b;�!l�B�%,��_U�Zi�oU���-����{~c]E
>��;<���8�Z�W����L���:�������)�8�xJ�/�V����	�(�j��o7Y�L�����SZm�`'\���F���3~�
���۩[��K���L�Y�l�Y�|���*h)�{���v4:�8N���{�#	�|bcR�����V=�F:�kb����:J�̰(,GN�r�&�$��v/)�,!�1ڢ��Rl��D�Zq��)�u���c���E�YܫN�pR<�-�Q��{�м������m@m��J��bH�2���z9{ؙ4FD�"�Zo����kb�:yּ�j8_o4l;���c�����:껾��Ag:��s��w73*��b����t*�.r9�m�(G��U��)�m���|ﻝ�zA5�L�[�*W�{*�;��H�s�k�S��D��LU�c\C#���JE�*�ZJm�
bFQ��]b���qK+3n��E�i� ך+x8��&��{���V��-dx��7sAyӂ�x�(�O�L�����/8�:���`
]u}�ڎ-�oN�}W*�X_7w-G��0.]�B9��mQ�v��D�1*H(��X�kzfQ�{��u���������}�&����z�r����2�ݰ��pgjc:��L�y�Hۋ���l](/ov��If��2�ʦ0�W�ï�f��}W�U�iV3�f
��q��y�	r��b��4�L���.�k"������\:F�T�Ǚ��~ue`�n��oq��{|`�1O�������u.8���3%C׏�'F�8��3�c}:Kg��px����Cr�;A-	����kEދuw�<{����s9{D(/.�-Ӥ�����1��E�a��ڵF���k�z#+� &����!��He��K����s�w�q4p�㺯F�V��Kk�����DF���9���\8276�mٵ�x�9��m�lDۛ�3��^�Ƨ��l��M�����5�c��}��*��|/c���q�&;9��e�<���+$��VӅ���9���n�b����)�h2���C���G�&Ĝ�c�i���u�!�kubo%$#�wM�d�/R���_V4����҆1 �:�@&65}臩��üd���x(C';�4Wvs�-n��1�<��&��n���fX��<\t�ӆ�l;�d���ዜ�xUt.q�3�
{Ntk�2J_xkÒ��^A���\�����zcă|oW��Y����<,���o�7^�d��4�WMJ�4�jɨɖRK5��=�d�x/��xrFf��Ɍs�pV��Oc����h�B��Q����SVwli�P�-�zi�G�}�&�sv�ܱ-��AS�d#Cs�ۤWn����=��f*�uJ������f,�55j0�N��o��{��q����wA!�'�'ִq-j	v@�=�cI�\�(*�;�pK���R.-�!�%��
�R���y��m'd۷���������1���L_F���'f�$�h���W�kC���$���L�|Q'yu��K^]�=�85�=��X꼊���U-[y/ ӑ�lu&�A{1�u�6F���U���Tdyp��3~����X��y�Z��iC�3��A�;�]�R=��̗S�fn�tc:�(�>̢�}Ճn���Z��qpD9��׻�w�x&��T���4�F���*:����<?y�w����v~�MzD����wA|�1uq�Zet�.�*�ƃ�e��T͘�9�C��dvc,n,�F�Z�q}��Ն7�.�Ϋ��g��L�R�v���Еվ�� �h�ri�kI�ܗW�Z�!5�"�8�V���m�Nbi2�]��9u$Yd�	�����c�G�ҿ)1RݹdE��u�3&�4K�PڱZc�FK����v]���{33z ��J�q�V���.��J�ٝs7 �7N'u9(�u[[�`=kJ]�]أӖ ����7��J"F��@��3���<|�mu�S�=\���]P�Q�&ck�٥�w��7�y�vv���m���ջ�������9��kU� �j�Z�T��m�N�E�v�܎�Q�%M��m���0WD�]٢�L6��+.��V�ؚ�}�u�������9�����gL9y��'p���� �7o]{�������(�S�I��V}��Ɏ����K�>6ħ��m����Z%����m��9��f�N3r�7���j.=���~���W��-����So�@:�*�#ũl�s�ninU��1��-�g��V�v���f����)�S^3Ok�5�;
md���6��G������g��ʋQo�^��2��.��	���g-�durŻL՞.�`j��[��bB�]�@�uU`��ǰ�Ռ�;�"�QA�yB�j�v�e;'4�e�h7�oCCy�b��R:���^���l*��Ch��w�+O,q<�����V�G��,��)�63u�edۛ�jg5�;sv2U�F�7��7V�5�[R��6���'���Zs%pE�pg:��V
XnC�7JزΎ�u4��5���Z��BS�zU�W76�wx˷jZ\'n�Z����򲰑ʰX��)��W��U�fĿ�r��^�Ѵ�wK��Qaܒ�\S���oBd�P���JfI�k����Śr�SXN��e�{��m�[Y;���&�ֵ��0l��o5�*+o%k��,=^~���x����u�
�;�1�E <[�H�'$�Fe�u�\#�v}�$�^�y��s�py�emc��?���AB�=
�z�$��%Zr)9[E5� �c����N?��=�t�) � �v�F��Q�"H�)JEH ��b������ytN���5�i���"/d�|E1e��e+�9ٝX\Gd�n�G��ʑX�b�B^�EE��q�� �m��F����������ߟ����wڵ�?�!Дn��V�Q�|�Gy�K��Y9�~�o�ͽ΂�
� �M>�NTZ��Ы��J��nQ>��^���Q��d�DN�["��*o_q,[���֖��-*��,9o�e���ue�lPF���1i1{��9N9'��?f�0�t����\�=g�>ި7�삱�z�'�9uKؖ�`�9R�H"�ob�3{]V�d�t�� C�@�9^]��;/uX�.�Ϙ�M9�7�Y�c��U$u\��;	@n�F]E�KC��w��>�V��V=���	��N�gE�ٞH.�%	���5��:�Wh��Ek˥�ܝeRw��%d��分����uu]���i�_���'{\�G��.�Zu�sJ�ō����o;)���Cf��¸�ohsJZq���2�-u�;�u�*�AuCv[�w/h]L1c�K��=��r�t�$�<!��<���K�6��Y�u<��e����Tx��/?y������J�N7�{=��ˎ�`����1v\2��5�]X����D��<����y�1�"=k�D6�9�� ����p&��cMB^uum�\K�*�2���>����	�3d7�?�^^�5���tW�8�4��yy>���W.�mӔ��!陹�2V�XE51��&Q��hi]���˼{�:o�K:�D�Jxu��r�`]� |yH�8�e��Y׼����� =\ƖGGm�e�X���B�f�_jXz��t��M�h�D���9�E~�ܙQ�;ܠ��OK���:��lti�-ԯ�i�H#iu1��1�[�$}�^ݭ����h�=o.�gNf�b;u�ʸ�F�w����l[�q�2��]9MS��'w��ݙ[�:��9ٽ�]C��PV�
��%aJ�v[�+~�3 ���\�G%u�ʁ�k|�U��|-ڛA��Z^f�2�ӶK�ۤ�fm2���,Z�46�K�ed��[�8�ͪ��� bdm�	k���z[w)�ý�t���:�REKn���&�M�,&]�x]o�����3�ǖt�~�������w6QH�Z/��6��y@�ț(q�C�ݷ��Gt%���?e��TEs�{��=o��L��c4<��T �j1�]��Y��[���|��II�����s�����F{;�1�F(��w���3�({�y���#���r���L�\��nC�]^�r=�~[��ѬJH����iYI�P�$Ϟ�/k;s��#=jΘo������g�o���D��?;=�qL�su��x��*�Χ/90�=*��C��\��G���F+�Oű����guXB�,�˩\��h� x�ŷ��������IT����εQ
�yO�>u\�R�@7���>G������M������(|K���z	�h��K�n��=��8ϩ��SWV.v����rC�r������g���-�����A4a�]�s��Z�F�����7e����)}f)��p7�����j/�r�O=AG|�k]��_S1Eݍ��уZ3��\�2$[7;�]�v�H��xv�	�%�r_V&is���֞�b~�R ��=��o��`nI���3;��Kc6��Ν2��:���ӇM���D�]��l��+J�l{��eм]��*�V<��w��Y.��tQt2�7K�|��;-�Q�(�R�����0�2⡎�J�ԮTdR��8�$vޤ�d��)|S"Z2����@�
�]*:֦݃M�v�U�Pbh[����۔�b��ںE�B��xf�s5T3��	\�KD�|;�����x���(�B#�"��0<� <�XC�u>�W�cX�O�wz�P@��z��Ý�H"v�)C�mL�dC�����L)������8�i=}i
� ;�O	*,�;#�d��nL�����ɮ�S�P���c�Q>nvdKr�[g�V&���̃�捍�:`����;�V0Z�1�+T�0�r�$�`����r�̠���*��������mZ����2#$쏫s�g7H�> �虓%�\q����?��=��=�x�;�9�%�wK:P扵p�V&Z�	sJ�՜���j�y93�]�&�.�H�0��6���Cǯ�l����m��X��,,W�OI�N�S�3��F����.�*5���+�r�;f��jq;2�h���ˁ9Eٸ��@���U�
�߽�c���{,��ds�s3ޜ�5���}(���9\g`��ǒ��,�Ik���U=�B6��������]$!�����#�;y��ȕrm�B�7��U�g.���oA�'�4�>�7F䋲{$�b�'���,���c���,ۮ���w�":��_�vS7���A3R�(T��ԳAp³9�	
�Ԡ��5ej(��:���9�p oH-j�yՂi����@].�^�
�kF��K��+0��e�"z<v�ث��L�}OQ�X5J�$��L�=�ܗ�.xߑ�/x"���_:�um�ɹ/]|v��C9�u��ʎt���~B�1x�Va�t�<VW�~�E�4����//�[�l��N���Zӛ�"!����aM�\t�.�Ay[�k����*(��x-'N�$��D}u
�.'�k�K��l��Pɝċ��=��v����n���^8yQ�[�ߺY;gF���cW >}ʾ��1G����xH�96����S�p��ff�+>�ԫЎPK�uj�z?��E��ܪG��^� �X�˷O��|Zu��	uxn���99:��zp˚�*�Vg%��q��%��f�J�_?{[E�=�j}v�9���`�l�_h�Ej��\V�a-�#�o;Y%�����J��5|��VT#�J1�ֿ��כW��l#՘��R֪�W�Ӝ���� ���X���y�k����Jt�~�?�
�c�����t/#��%��uזtw��װ��׌0c��d�+���
�ye�\����R�c����#�ک\�R5�页��`��S� �XM���\N9m�8<��罕I�
�bI���O�����gAy��Q�8�ѫ�[]1T��p���m��g�[}�����fon�Z5[ƭB��>>]u�L�9�6<R��}�3~�(��&hi��b���Ha�����͞��Zw4�H��|��������R���z�8s~�`���S��}෵����6�r�wv�e�YI����T������*���<����]��h�qN܂��=G����{<yY�z�7��y˽��O�vt��2�g<�Ƭ�2&�K5z��	����PޫA�%���L�mX�K7�錝�6�wnT���>�D/�<}uo��	83�1��fs�<VJ`��o�䗎 �)<A����,\=�F`6�@�y*�3��QFܩ�9�B�a=_z������f�}k�s�t��O�j8���\1�7�nf\���
{�[Vʮ�f��iL������A&ޮJm��&-���e�׎���հ��BZ��S�,a�����E.�k��im�p�X�]�X���l�Ҵv�z� �#��>9��o90���Y�w�B^�gL�'�tI�>����+��o��\x1Ưc�KO�������KM�WW,�2�v17׌�|�O2�y�8h`��9X�:u]����g�l[$l�{tM1�Y�Vf5Z)c}�����\j�j�r�c���2d^��C>Z:p�u��v)z��y�r���ۦ�$X�q��k�D�T ��ȍ.�N&�[Y+}�G�����>�S@�+�l�x+�L!�xV\0�uwr3���>���I�I�5Ղ2���7]y��K�l<��z)�`�N��,�k9*Yձ��0r����_ǯy�j.&,jÙvCZM�
p�x�--.�peB���tB˺��9������
:���4���ڝ�X�u�q���l2�{���8i�Z�t��dQ����(c{�pW9�^�g�c+���y�]M�(�xHn�c��1w�=�����4��
�`�űg�	�M����Y���f֔�E�ASr�rw9��ˠx�ɛ�<��3�3U2��Ф{p��ս����᠄.>*n���t�R�wG��#9w����G�o��j��x����k����X���) �(���K�u̥�����z�a�r�^Z3-&�3/�K/{Vm�v'�B[9��� ���*����/A�x��w�[y��[f�;�K/3��շw���50���nw�RwI_LQc��nu��h���of� �J"��̺��v�	��Q-d����g<úpu=�V7�ݻ\�"���dQ�C����8�G�����$;Ռq��I|�/hz���Ptv�Z�ۣv3�e���MŏLo����*y����=�p���-�a^`.��2�78���lA<��\�����Zv#���bm���ۈ.#��W��&��v���9�)E��v�-n�^��[������n:��z�e"���A�06��y1�{Y3�����g�h xi|�P��o�j2���eKE
D�VM��Z�/x"=����b{�����˓=�{'��i��`�*���|�.���}�u�_?gU,�����d�aqE�լ����4X]�[�u4T�S�{��3|&][�f��%k�ɘ-R�M��Y�Iֺ���ja�4��L�7m�.�����u�#8d�˺�r�s���
8ܗ�娹���� SW�ͺ0滤�s;.u�B
]b+3�L�{X9��[���3R �CC3�˾�
�іC�|�e����kڱ}�?�~u;к�?n�`�.E�7�4,h{�
z��{O���r��T��)��:-˼I��+�d6y�sФ�d�o�-��.Χв� a��
�9u�J��eV�P.�w1�z�����&��KE#y�+c9rd�����Mu|	�5��q�Y���/S�&�T�m(;J;�>��"����(�)4�hc�µ�s:���F�4���k�������}���FШ�7_<�U=���]#��_N�(���c!��2�T���ûb���3yQu�HQ�80��J���G��!H^���ꃰ���--Aǆ��<�jW-���:a���ON���X����$�@�znSܘވ���5&��1F���Yu�!�c�^�j�v^�/9�h
3}=������8�^B;�Z�{�8�I��(�F� �H=��XUYi
�{��[��@r���-�� J��:�"�ݗ��v�Wj��O/��1����3��.�z���0��S���,s�>LW���ʎ�$R:��9�d�-�lU�y�w�@��ٚ�'��yq����
Ҵ�Ҿu0닲��L�H����!;�uw(��B�W�Z�����u�J���Q���+H�Fq*��Be��閇&����[�ג1)���Ӳ#Lh�*�U'7D�s7w**]m]�Rf �G�z��L���ݓNe�����0Uq�Xb�w9�﹆M�hܙ�*���OK�&n���pe{�!�.�LL�,�ε^z����"�h�{�@�x�8������]Β�/��\�v(E�b-�:E�\<�Guu[�%�"ݖ&Gӹf�CB;E�n�n9�ie��z��	|"6���Jq����(�o|O�ۃ'd�G�3��9�gk��|��3��;�k���
F,��v�!.��l[��y���E�t�>�˥����E��I{��^����{�3^�2���"�
c'[ծ�W�O]Е�|�����1���{���񆷀
o��a���yA������p=�KG[�ŦE`�8�x���&qG�)�F�4�+�b�_U֪%�E��yYN�V���v\�0�|���FLI}\G:Hҥ��wm;/��.TH�ڌvW�xh�7T1t�R�b��4;��ΰ�UQ@��5�̄�A�j|��N:�US���'2�M��}�{�1n/y����<״SD_���[f����5jt&u��xY"QZ4�4���h�N���7s7�m�|7��Jxߡ��J�x��/ސ���=��c�J����F��-�/+�������ٹ�С��c�=���Nw���2�sw_ż�{&Շ&h�R�6DW���y�:z>��T�;ʻۨv�^<Kɜ�jpW���5������7�nJ���:�D��lϴuM�|>^����n�7~�8�oU���q�zQ;��l�)���w�y��^桭1j���iX�"�!,�j��ص�.K/n>K�s"��@]�+�6ewA�w%9{a�j� y�����D�G��;ؘ��	]uP��i�[Lr$`T48oixŝ%^��J��^��v]���v�{�����}#gm=Z0`�m���ƻm�`���ke>݂�uNsC�����q�V�!�U<����a�pA|����eV��n�2�C�݀��f�S�\桹J,ׄ(d��-)w&�1v� 4{�}.ip��5�O�D�e�5b�n�C�:o	a�]�T�%�ˏ�٤��.��:��ө��d�Z��-�ds��wޙ����=��wX�x-G�j� ��ٸ�^d=�l)�u�Y���ۤH���#R�hS-�x/�יv"�k�m�6;#i�s16��K����6-�L�Ҹ������=.�W���;��͂�.t��p<�1��[�WJ�[5���V���fX%�g��`Ψ��D��Lv��N�&"�B��f=�������ɾ�޾��}�Ɇ�G���_}�5�R�M��{�`f�a�ŭ�;�a	���������nffs��u��!,h{�l�.�7�7�bB����2?��px���������q��׽�P��/e���#j�˓@o1B�e8�"�J'|���:����� ��i�q����4��;�/7���ݻv�۷n�r�������<��p�Je�s���g۟�1�\s�8ޑ�u^�p��ɛXY}7؀�S��3{,���M���U�ʁ�1[ח�BMd�X���ަ�ˉ̎_f���m*}y1��V]V`�x[PQ]��`})T�������)�n�w��}�ay��ʮΔ�w�4��A���/�5���+\�o{A>��|�|1yw���������%d���J��w{h.����WQ�d�{��x��I8���.�Jb�a����ͮ�ߍ��ιI8�y8©�J�Q��F�����[�`EK�.�Jރ�6�O�J���T�ݗ����J�X���Vgc�:`�e��x^�{�F+� ���7swl�ۖ��|�P.P,ڝ���l^VM�c�h�
��w�6�<y�\Y�:i�3�6r.f�bT^���B�fmް� ��Z�F�D�����L��糱˺�Z��p��'���Ƭ�/��/��W�!�owp���S+s�WU���ҧ�M��o>���+���S6ygn�ʸvm�.��׳��{�z�JQ�\���:�9�.��1�{���MDμ���w:��GT��gU���ćd�|�G'M�d��B1�$�c�W'��x7���H�.�(�Pf�@� ��<�5%B5��z��p4�]�T{���73b�ǓZ���̑����q�ź�(.Gy�w���r�L��)2)���]$�>>|��|�|}���h�R$�Fĉ`�E1L2_]��, e&Y�D�K��c1��i4A����I�fI�A%4$Ȥ�"	(����΀]܈)��wU�J��0F4��I�Ja$��S,CfI�t�%"�r�;��"+$Za��]�c$JH�6aI);���A�ݮQ&���"�$�i4F,cQ(�۩�I�@��Di6�,��0$���D �:RY���h�(�$4�Cd� 5*`����ȈI�k&�wW9nRd��AD�Gu]$`��Fa)��i(�A�I�̬�TP�Y"��L�����ߦ��=����vn���#�W�{:�L�|&�1�6{m�:��)�Yn�=]Փ�����Z��uB)��I3+E��}X�nh�Z����v�"�GF	ت�d�8��T�dVm�Ӗ�Es4w}��A�'�$�y�5[�A5=��מ^�a�~R��0:0\�< 
��r;����I��� �����|+�t��j�Uw�tS{�r<��[��o��/zty����1N��_�o*{�������~��� 9;>���| ϫ�9˸����nʒ;{zO�N��Y��7x������]�3�L΅�s���{��v�L�y�7Gh���[d`�0F�G��D���:��n��x]Wgk0ߑ�^žA�N��Ԟ���柼[�w9�E���N��"��s����fN�=tE]N��S8���}�^���=!�k�yso���觭��[yz3�/��_�-q�`=�\�m��;7@�_{r�g�)�����1�KU��M��� ���b�̇���0++�m�&E7���Q��]�e������<��Z�x<�{g*��T�6s�����n̛���*�.t�)����B�z�">����s�q'/�O�vH:�
�-U����v(��b]	�4�_��[�b�ze]
���V���h�}���<�{׸��W��Ik��Q��j�<�Uꂕt��:�r����z�Lh{�� �D���n�Oq"x�4�G`�Ǘ�v�: }�m�7�v��#����"��so9w�4�=�_z����<O�4���xKgeb�&=���g/�2�Vm~�bpe���Oy��2n�I�i�s<���wd��:|��vâ>5|ݢ��l��Lf�7�H2(�4y�$��ˀ�ɰ{ޙ�Rc�~�;��h���;*��$G������Z;^��Og�wjT$F���{�g���^ߞ��u;}�1؛�6:�љd5_m�n_�w	x���<��zA<j�/e��θ�R����g��X���b������W��L�7��'���wdwWHkl�>�Y�p�$lh;�x�W
|~��)�/�mJ�]�w�z��"r�Pw��O����</Y#��T҉Ut��.=��z��2G��ˋg �a��/쵐�?���&�\�����g�HMϬb�#TL���,�I-��?.�[���!�<�p:\mcBh�tLЈ������y��pl���о-����5�t��g�=.w3,�5��E�{����xr ���j��i}�v3���gy��bD��6��-�Y0������>ܺw�J^ʺ�a��������<q:+_�m�6k���;�Gᵱ���1��G^�3�;�h���Z��ԛ�J����pi�K�7����̺�;9]1��bȷ���NįL�y�����jw�9��|{G0�g�3K��ź	�ݴL��@wQ��K�/g�Vu���צJ�w�~�����+\��#QQ�h�D[{{�˲�%-P�RSw�f���=�>Fu6Y��[�S���2���2�#�P�Bo9������u<�]D�viݡx�~�xN�9��2�` t���s::�ۍ>�f�6Y�C�<,�q��O߿Lا�+�Iym�t��םM�W9�C{�>'��k9#R�4�����g������CL������ks�6���C'��'�'��\W���#�ճ�k������gAmf�Vew�8g`������]���hF^iqZ��ɧ�Sņ�▬lr��{�����Q�'i�q�fVM��S\oA�}��Ъ�X��~7Η�M&/$k�9�	���A�v�@٧5mp%��H���u痳R��#��]�U�tZ{X�8����h��<n�n:���œ��J����i�o��=�벨y�PR�֎+y�gI'��!�zx�p�.�7�d5��/���#r2HcO�|� �FJ|G���N�{M?Oe�gaL�����N�1=s�G���ln ���r��7g���ӫ'l5���t�O\X�i�~a���h�HS���������rUu��n=~�=�i�z��kx�nx%��H|��ⲼM-f�R��'�t�[��CCASdu̵�j Ъ�=rE�@9s`l~F��'�o���6�J��$A�y~� �u���=���ެ���Q{q[[�>���x��x���>ڏ���c�xU�z���	N��ٙ��ol9�['��X!5�N��o�'����kMq�����`�xvT���mW3���`��� ��g�g�ፈ?i���쇌�t��-��nIr
���T�U��ޖ9�U��m�*V��0S��(��V�s_(�pJ�Îj��/p�NQ@��Q�/�+2���P4��,��U~	�팃��ӯ������o�g�]�-����fn�1�ֽ�X����@p��柮,��X�U�� �D�&���gsL��+�*q�N��xD�]Pgޣ0w{ƳO�ܬX��t�Қ�G��^�0��4D��#�rg��F�X�I���}�n�|&�v�����G����^�@=w:���sj���g<b~Xkާ͂�GE������@FF��k �}�}7�<����	��%:G9���C����ۑXσj�.@�DV��V�� ��P$���my^�&;���ͩ��ﲣ�pE�䃓�$c�b�p�[Ц{���,�7*\uzW%*���ͽ���ǈ��j�3���N�o�| ޷���<�=��:}J]͹�}^��������k��ɑ|������K���d�G�H���A�W��՜��,��1�#�WPʌ���@��g�e)�-��i��Տ�Z��1n{~��t)��K7��J��l�vy�~�'�ze-�;��4��N��3��kO��e��[}�$ǁC�JϧBs��N�+�ڕ\��i�9���خ����j�y���g�ϼn��=�Kn�n6G�l�;b#`��OSaů�N�>�pGT�4M�tx���&�d��u0�6Mf����]���v�ߌ�mؘ��^��,Md�q�z{�8i��!�ef��j��O�ʾ���k�D�e/���Jr�x���S>4'��e�H<.Pu��U�����i�ٯyO0x��d1�x`=}C$��h�y�j��`��+��ޜ��J���z��O���&EW��{W�|~���t��V4C5�
�cs�KA⠟cpӝ��tz��H�$O"4�G�G���n�GG���4���2܋=��^��>�m�ܺQ�O�ɵ����]�G��=��K*N~��'�]f��Ty���ﱮ�������A�n���m��E�v�{˟5���J|�h����]���uw��q�3���b�4�[ӭ����}z|�����ܰt�{E�"���%�'g��/~O�����Y�j���p����?$�q��MK���{{Px7�l�l*$.�% \�%��جT�{��:Y� �#R�; ��go��Il�u��GO*8��kh;�{�=On�hs�o�x�2��
l=��<�~���:D�exz݇��o8K~��y�u�X���=%�~RVD9z���9��~�Y�0%���\{��8]{������;+�K��Q̉^8����3�	�F�.{��dT�E%�i��-�ߺ��zNU"0��zz���$�<�#ryŖ�M��ykޝ�ws����^�[���)TH�p��#4l�ړWŠWy��:l����}׵��mSźN?�o8x��u�>����y���|�����6��m'�u�������Rv�e�]bV>�w�>�x��h�2d95\_o{/K�������Q͑7����k����~<5p�a�@�����O>��r���)����/�Q���4���v>��^ku~�l���"�g�guVDc�z_f����&��c�����~���ƹ��	����hkX�b�EkԦ�k�Z�wܻ�M�
*;��&�Gph;������e�?aa"��Q�����xD7p[��r��_���73�d��(��K�]�r����*.T��:�5/���Af
����܈v��T�z��8a1Uߪ�q�;��%�7M����r�O��,�����r7�嗞ޕ;�z�[�ʔ}�3����Φ�Y��[�W�̱k\��IYY��NV���yM@#���עjv�y=��j��`e��N��:���/��t�?}�{C�.��,�0fz���p^(�x�]4���zCp��ݒs��
1�N�Om�����bP~���k��ζx��E=�P�$��7�J�/��P�O/s�Uc��VD�>n�l����=�h�1�ه�O���\�\�z��52\q���s5;��k3���|���W�����ez�>V+�]J���)�����=<~�{:a��u{��Q3���'�ӓ�x/�ntF���5=y;}헧����X�s�n�U��v���ݼ�#��y\�����v?��?~Ey�nt"�s�wP�~��+�wpD�ֺ�+iJ}\{B�����X09A�o��۠=�����f�?/R���u�(ʱLd�nsu���e���߄�r{:6V{�b��s�].?q}l<�s���,c�{k�D��R��s�������Na��~��i�^}�t_}��;��?C#EK6W��#���(��'�=4����VW�����/�&*�Q<go��w�Y3�{�X����s�t�� 퍑�WVy� a0���O|d���_W��)�Ĺ��4�އ��~~�[&:���'�Iw�����M+�M_b��j��XE��$��m�}}#���Ua��c"s�F�OY��,����o��!{Ꙋ�`�u��F�q�2.�:�A8������č:�:�ا��D Es_{ٳ�KㆽLk��*䙳�����ެߌ�I��z:�{|Əs��Vp��3�-y��C���ў��Y�������y��^�w_�{�޷�G4BU͵J�`��iGKV��7��d���{�:r�g�� Q�4 ��x�<�x���4u�/+��G�y㐠i����q��y��S���5x����!��h�)���_sN���0pOh�p���.��-�����Yk9v2��.��y�ӌ�e�5��s���4�K�W��Z�V�N\ӝU9�+mY�T�vv[H}j49͙�-]�H�n���J���ծr�z&%{�ǥA����Iwt�d�'��Awm%�oǬVT��Wm`���Vb�M�����]^��Q�7�<���� �w�ٰ���11���!�Q�����dADn�ܮ����Y=_�E�q�Ķ�H������a��\E������]���x��ֿv�^ei�WŦEqאn��=�Kn�q���Ɠ·w�5����]��?v-pM��OL߽��?x���g?gV�yS�(w,9q��콻�����c�;��k�k>4=��G�g�9Jˑײ���~1���>~��pm1��ѥ�g��:�iL��	�O��ʺ�����~)���H����1r8������Æ�h�L�b�Vט�sN���[��yJ?I~A]�^㄁�7$��]#h7F�Н.[8Gsf�Z�r��ݻv�۷n��:UZ������d;����u`G)Z}���%O;n>��ɞ>�⪜����V�!v)	��UM��;3�w(GH�澂�߲(ND��)��]A�`�
���lyr���1G������Ad@����0<RpV�`��X�{9��o���nW'��La)<赈UoXg8)Wkl��������1���t�n�1�^~���g?q�#����{�������ЕŁ{����K˛����-�ڮ�9���r��dE��oL�s�Lo��F�s�<�gUc�����C;���we��ԍ�vn�"�e��L<�in��Eu�	�/�Ս��u�����9X�9B+&SR�c+lu�@�0I�ygT�����*�y���izu:z���ya`,_��9�3T��k�堉.�3���8]l5ە���=m�α�"�o���lm[4w��6H�����:��V���6�u�E��pfa�NT`�a}������^Us�A�׷��~b�Uwx,�<��q:���2��7c�Ŧ�dqɝ��P7�e�{�I�R#�
<<�=M�nk�{ř�2
�h[xu�
������lx����#�WE$�[�	M_o3�׉*������g{����q���F�7m's��jC�+��
��tTOL>��t3%���[UR�DR�)�3ô�u�H2e=2��� �Lm���ʒ���Y���G����O's�{I�tyO���6�|Oz����/{�%ec}��_ ��]uhA*"�e�w5��VU���~�����s��1\ջ��{}�m�'�m�Ւ���vuJ}���p�F���p�ee�	��Q���)��w
�n�����Ջ��Y�Z��9F�7��7���n!,�WAx�8���ו���]�F�|	}�f�`�-��{�N��^�ά��h�ʰs���Kj�n���yõ����e��D�w����3F��(,�ͫ�l�o�n��y�Q�4���݆�iWM<�b����cWA�-TAeϛ���3�۔�{�W���Qe�����BG�6\����y93��Ts����V83�Z���}�H�T�Z�<�����ڏ���{ٰP`|�_y:=���0�ܮ�n�.%�� 7.)W\mE^a��S��ХݠU�v������*��-��$���V��A��+��t��o�����P�ޞǇp���"����U�M�??w�=;&4mۋi������}�<�qI��ږ=7N���ֱ�[y���	�v����΄�'�Ey�>ɝ�	^��I|c��c/�\�-v/�:��6��c:)z�(g|wYJ�ruĩ� Ȩ�ƸGO��� �uulN��5t
�;��\���x��C�Յ���e�n�,�Ɣn���������f�"�:���
:���6���>A�yh}�I��E�_)�I��H��Js�]��;�}�9�zW�h%?�e��&��F K��h�Jcc2@C�λ-!&�!3B  ��(Lc��Hi�v��3�I�,X�ɡHTFG.T�Dbdb2!�I1@FT�$�"@dLc(���w[��bM�ADh�Br�E3I��&��_�&œIbѓ"����H,�IQbИ�6CA%�H�k�ʣI��+�b��8h�wH�F��];wi�+��Rb �n����qX��ѯ�yӻ��\�ƻ��W��x�E�E2cpۧ:�<�xú���]�wx�Ew���s]7-t�;��I
�y����w7�E˦��3���������k�8i�nm��S;�2������t��˜���r��n�w2�D��KI H$~$���x��D��Z��Y��vO>;X�8�<���m�	&�Fuȸ�+��Tj�.�P�����4�\Ay�_\0��
ww^����a�nL[Q��c��ƃ���	�-��$�h�BQꆐ_E��lEC�<3��Fmj��-�o�.�*�q����g|��z����ng��L�}�䮂�����Ng8�:��6P����1\9M<7���
.p~0�~0�)z�Oӻ�Ώ�ͨ�ʂ���팢�r�9��d��&O�~��j����56��W4Kȋ�O3��y�"cz'j�W~���Dt�/H�6�n�s���S]��޲f��ON0�ј��O��<���� �*d$Gf�!�������+TӜK���h�"��b�c\ LK"�SL��o����e|��W����<���<y�&rzۡ�m�-�7S+�l聁_<���	�p�'8�KrH�kk7'��"���=b�PP�E(;+oS��I��*Y���p�0Z,�w��$��S��t����sQز�vJ�yBM:����a�w�ݬ��Aa�C�mN��:m���*]��&�z�1i�g�H%��I(�z�e�T��^r�]�L�%^����� ���(��xr��V'\�u�9V�ل^����D�:L�>�M?o����=��'�V�U�H�&6������f�<�yX����L��Z�O�XK��&%��7�O-��%�xM�6�R�!W:@EkΕ5>���Ss���I�=��Z��3�����`.��%��p�t�_�}��CYM�D����=����b]�i"�1���"~]��W/�OAG�o:����]n���wl��i�&7��,s�R�s��=U	�TF!�� എyXh���T������+۱?�ys�r+Ps)�:��X�˧շ�Q\k�p/�G���qG����o��G��Y���Z��!�z��?>��g�ᆒpo���~)���Qj	�c��������%�<�)�gW�H�ܵ�h�gm	���1��~�����Pn|9�$q��b8˱�a ��HTaOK.a�߳�7�1�������J�e���5��e�Ӎ��6=WFY��l�vo9L�#�zCb��~�\���?K���Zz�)i��D����X
ݟ���s�u�ح`0A��HsV�fK��U���	os���.�!�1���8ʆ@�t��p)��'$����7���h��,eEV�ڧ3��R�jЂ~ka�j<%�y.�g/��ٕk��38A@���d&���Qz;1�?:���a��w�+s��j�-{����
W�TXSPW�7���z}m���~ciaSͽ[w�]ώ��;�=)5���o�H�]q�����p3����Dy���/2i�Q,��Ӥ�wi�"\5�)�&]��u���p��w85�$�C�#@S����+�')�FG��^��7Q���;�==��7J��a�����[���kE���g�&����t%���3p�_Ib��'�b%9��W�TS�a膖�fȓ��n�<F��<�eŴ3�+�>��cH�H8~r`��do��H�J�L�8LS��X#��]&mk֙��B)��dl�|�����~�!?P���q�YT�ν-y���6�gq�\�]ڍ= ��qu�`sN.iz'�� -D=�C�Q�ܨNu�����q_�ͪ�]JZ	��7P��W0��+��\��_��x��؈��&�/��S��nov�ke����=u�����u�ؤ�޿O\�6����E�Z��3j�H��v�4��@�|oy����yj���</�B��<���A�hgz��`%+u��Z�9/L��?��O0�̼�k眼�r�N|B�0��f��ZD���-��,9��R�a?Mc�(v�)Z�U8<� ���ch��l��ʼ���?j<�cC���6����fI��K�N���4c���y�,TRV|gO���QƎb�m����g܅�j�1���$y@��a��V�O������oC����ɀZ$_m�nv���t���2w(+/B�a�P���:��X�&_�ٚ��>�ͷ�]ABc�^�	��v�RC.�|����V��}p��C�'v�釠��!�B�;�Bt�o�-qc�.��(�&n��(�5��6�`Vd2�~��⟝z=��GZ�
V�X+�/���X0��=����9i�P�	������#�l�RM8^��k%Su�+�SQm������z�lZ�f/E\�3槹t�:b���L�=+�L>�W��s�se�R�5�v�?h���B�B;�^V�������!sߎ��,�R����7�#��b\I����2��_ClU,��\S<N�>3�A�3��0����)w���R&�Z2)8Y5�v=3�ˋ��*.'�f�(j�ס�V�^���Ơ�I��!��<�_(��B�[�0�17�s�pYOۋ��R��EP��{3~ո�ʅ�I���}��F�,��!=z�@!�@��B3aNE�~����/�5���E�� �L�躐�ƼQ���������֏H0͒"�h�Sܞ�c5��To���a�����͘����H���Ɔ�S�Q�NY�6��z`��;�p���{~�{����p�Ƥ��8j|$�N��Ut=z�Z~k�J�%ߚ�ך�8:���*��yv�Q};��*��_؈,�t�W�6Qurf�����J�/K#��*�����g���u�-����:�oL�;FB���@�v�M�Q�}��`42�s:���5r�E�f\^z-������J��89}�˓�v�w<���k�7*�jžn#.uv���.����}����l~���^]��26 /}}誕��k�?hl���Sٷ���{�U�rV�]�Df=0���8��`��G�í~���mW=E���6�}˥k��	<>L+�߷"�]�m��zޥ�\�n�htY��s	�yF����;�/z[&�V��y�9�ʢs-ݼ���tm>YS�Ǣf@��f4b�;0�p1���W�55g�׹�ј^uXQ���y;ɩ�2�E���`�zHz�$@�b���b�Aݎ{�k����\?^�xμ�����0�f)��V͗�'c5�gdf��K�t��M	�CI}����~o+3s"9�9MX��o�k:���?g���?4��>U�������i�j��q�J�!����oU�ɗ,+Mrݿ�,�g/�)i�5
���������9��G>^��R䩛��ɼ����vg�s��9����ߒ����~ϣ�f|��O��ROX�����¾��
P6�����2���k������T�'�Cs!�Ms��z3������q���Y^�	�	�}jm����X�͊��+|�U��A�!�(q�d]#��4������Ξi��$�+���aʪ�b�F7S\D��g�v=7E�Wک�w��~�%O�ȋ���wu��U�O۲�8�&����udk���#�ۉ�5M��78gKsuO�A+2�c����2(̧�[�`�ʟ�����{p/}A�������c�}��-�m�fs�hp>���kRB����v�����>8H"�i}�N��x)�%�>Ƽ���Ϸ�o�"��{l���T������݋�H�fƑe�Н���,�7��'q�T��b)9X�"�b�a�Oj�樝[I��~ͮc%E:����l#�!�M�;<�:m���*]�Y����~O�[=� ̗�̨����'�y�Y���W��aH~�C�=���CC�ܬN�G���h�����%5KS����K�lx[d�s|�!���H����k]��˛ƽ="��z&�\u�J��O�{�Dv��^�i�{zJ~h�d��W�����fڸ�'f��O�@\ӫ�g���o���;cQi��];^�O���BՇR�ès�̵��}[`�W5������;B�_#W�K��t(Ez�X
�=	�}}��hGVI��'3LM �y(�ԟ�{0��{��6�͍e��w�	Q_�/�_�5�^�6d�wW�s�ÝBk��v�2�X6+bV��P+�����Ǯ�0�V��^m��6������o���:��l�'�}��������`�'`{7���1gN� 3G�y�����:~b��@'�Ia{8PB�ho���Z�>�����"��]e�DK'p.,(�r[�Րi\�fN����a�8��+��Po9��
b�:�)�6���^��u�An�z�Kfe�]]]�Z���vxh�}�{����]g �
V7\�o���A���DBE�7���?f�I?�<��,"�{�d^�5r����ٕ"ʄ�GGR��᳏'�U0	tj(� Ũ�CPH�*�l���Y,�Ih��6�@(����F�4�s���[�S[Cz����oA	��� ��@�4�V3юoccd�C�p��Y� �M+�k2�+�Z�Dۍ�m0�wi=:ū�&=�A�{Z�g�Ӭ�
�RXKo�d�ź�)�QhG��!��Yv�΄���
Y��S��{ײ��}})�s�d��D�%)��S�o�lK-����]P�����WN���m	�^����:A�����Y�i�]�M*L��}����tXH��w��چ�`��tO�͗�|��1ŀ��0�'����Y7�m�̕lg*�{'�?_t����b��{��"�ع�n��M�fng���p�݈n��B};|5F��}P�=2�������xN]
��u�es�P�Qy*Y.�y<;�Gd><���/8��>���s��Щ��q�K�]|�='(^1�n+x�,(Z��3a[ַ����>�uz.���XyvPV�4���j�{-I� 㴉��c��u����os�=��5Ӏ6�i������t�gv��ӂ�����)�r���:6��#޵��=n��Wf=ك����ۏ52[�Bb��ft݇~&㘕[��L���}UU�U~��wd��	WH�5���1b�5����9��Y�E�P��pOҵ�%�T"�C�����;s)���}�T�{{�5�'��!f"���A��19�=.˨a�a�XR�l'�pv��-��6V3Ɯ}�N�Xf��^]���p���z�	�<F���*Y�u��޹\�"m\�e��:;��0CTO;P*]�^��3�tF1��l��^]���^a�>��q��e�����s�λ�Sw/L��Z44�$=x�4�].��tE��xc��q��v�N�i�Pع�ƅr�Ed�{j/��`��̈́��U�@�UDך}q�髦.7��-q��)�F���_u;��~ �+�0;!�C����%Zqa��U-�y@Z�(,�o�Q�޼��]/k�]s�ш���f=Pꁊg��&Ɛ0L|�#��yl�%s�-�A��M��Bd޺�	�u:ۼZ��z�:z��t%vP��u��=�� b�|�I�&Bo��4�)�v)����q+&�1Z�(Թ�ॱ �'_��LT"�]���Zv��m�J>�`5��e���?��S0g5�����{.���[f*��=�mӈ㞀�YK���R�����&��C�d��o	�=���=־:���Ԉj�G�kq���^��}B�O������2�s�_�G��!C�뵯�i�F�[�t7uV�8�j>����6�k���x{��{�Y�&�U��>r� wL��Ĳ.���Lhi0�&*��~	�{^Uj���śl����_F���XW:�s�Z,�w��0�ʥX��K����,�\��Ԙ�Q�|��-�Ui�����d�G2������,��&�N����PX����۹��ˆ��cv�8^���\(>�`嵧�Dku	٤��Ͱ-XNP� �F^���sO�i1g;,e�x��f�Ɯ~Cq���-N�l�#��<�ԿW�f�U�Qkeb�oT0�֦��tT�8�&w��*.��>W�o����9���a1���~h��Ǎ��^hK=�]d�����=������(�|���qɈ��{$�W�;O0J<�о��W���͛�~$��������Ώ�����ɾ�_��IC�o@�	��-�WXh�q 2�-0Y��v�j��D}���H�3i�N�k��d9 fְR��P�z�M	�=P���WH�[�LQ+��Y�vK����ϭ¸.,׆?��Ք������ui�nf��,
U ����J���i)�N̓�b�qJQ��8��x�.���8�&{}i��u��)ᅣt���«2$��5��ܾf��S����z{d�t�wnTp�0����F�C3s�mԡe��b!tm���5�x�<�\�J-���F��S��ѷې���{�z.�$X�u��q�<�V��j����N���|A�|i��YbT�<���5.J���G�.���W_q�֎N0֠I���@ǫxU�)���a�y�Q.�$���{9�CH���\E�a���n�-��eMV��{�ӌ(�ǯ[ռ�|w �e��`����������X:�[B��<f�2z���A�3��Ĳ����e~��?��%�:'����Nf���t��'���5�,�ׂ�ܥ�Xu����I/��'�)��T�cIMl�q�!��6�M[Y�J#1pw���[j���
��4�6קg�,0�ٔ�$i�I9w�� �"��k9��*i'PV��~]ܱ�����K�����5��;Bl�z����*]���&�p$�s�w��OCQᜲ��RzԚGW��a�?`N'X}C��Ƽ9���+�Q��i�_a��T�B�7�2���[��7#���'�Cʀ�bC���q"Ƽ(����]�4����v��R��c�Q��y�1�%��V�ze'��`�ʨ�
�Y��-ݛd�4�$F`��2p�ˆ�]\�p�Ç>~��{�粒�{�p���A���}��խ�X��-���x�heM��mktW
�X�Av
�Z��h!]օ�3z�S�T�sE��h�^�0gmG����c4=��J(T�b���%�>�&�.q,�bdf��Y�Ȏ���D����j��TFL~�b�q���)�z�����>ry\ቻ��a��>�ārx� ?y�Z4���-Z�4�������'e�"q�U� ��[y��.����t��SK��h]��E�qk�����C��>�C����kw�^2yA����F�;�Ğ����͛�o`Β�SN�Z%>�?�桼 3��˕>�Y;H�R�Y��S�c/:hѯ��{��?_�Vt�����W�9�	���A�z|4q���޺M���t�<xM�Jj��RT{k
c���\2ý���Y�ȃ��4�7CNHQ���5�e��g�
�uG����v�zE�����K�@�6F�̏�f�/3��p��f�WiU�r�N�w{�T+w������Z,=���T3W�Yr�֐������5ӳ5�;x��*��{��7��+ޮ���ߤR*���m��/N4%6UTݱ��#Úy�^A�t���>L��^AD �	*��;�?�o'��0��Zu��[]�aE���N�W�173sд�G�g�ʩ�w �khl��SuNy}�n3����6�����w��{pU�1۠y�P9b���C[ث�ps�MBzL|�ʹ��r�8�
9p!�Q���c���9���i���&�X��H���aѪq�Z4��m��[�����BoH o���{]�2Vݓ�k;/�I��ćuD��$�ӵ^f��4i�/��k�\4�e�v�$��3n��2o��<�j&ء���,ä�^4�R�U6%Z��w����6ݾ�4�z�är�k��q�m�V��X���B1
`�������n��zL�f�|��{x�;�Y���fBC��h��[r�ɻ���wN��]V�n��Mf2(fv��+r��O�S{ӽ�������F�n� p�<�@񂥱�"� �n4�T���k
J�.|��4��抋,Qk9sD˙#r�Ѵ��!*�i�tj�=Ë��wW�8Oݧ	�q�VOv�+��)J���[�YEU�!��,q=�O� ]_q���.���V�l��2����K�w�����@P(�����H�7}���̜f�I9�p��XuZ�`��j�ޱ����^��� �M�=���!�W.��Ό���jUMM�o��"��am�*���FA�����k��WW��P=��o@���i�HU��c��B��3������S!Qd2ξ�I:�/�<9j��ϒ�[q����м�$vӏ諘ܸ;�ޮqf<F�}1P��_e�K�5�_s�we<�W;z��u�Fw9���F��1��Y���ee�6��Rfǽ�����C$ԣ���2��!��L������	��W\;��p�74F�ݨ�	b��Ts�r�Εr代�L;������uwdB���k�;tn(�����wv��+�"�;�^������G.\�gu�1PT�)�t�D$Y ����c&�ѝ�rs�����W9�&���1EQ[�4F�n��Bm�e�\�ͱo���$oq�Z��sE&�&1�AQ��]��ٚ"�c���8A#Rm%���q�c)����h��A�*1�H�J��!b&X1f*6�1���������y�����?;�1N���'��0Lzv͸S�i�31w� 2mZ�fD*wě%`�:��m��fs��p���xO5�j�T����x�~}�3�VJa�ƲǱ˧շ�Q\����!۞j��T��wu��!�k�0e��0Bd�;�,_K��u�&��|.7֓���i��.i�y,��PÚ���h%�������}è
���Bgh�����;Y-�u�9�&��m�F����h�0�m�"{�?jE����hwʹKO�6�� ��o�DL$��m�{�}=o�t�GZ�e�7�D?ٰ��f�/6�5F]���>r���l���$�3H��<?|��L��Wa��{�Uy,��^�AtV�v�A����HjHγ�l�,qL��sӼ׌��Qr��M�Ug.���Ь��=k��Ue;/4�7���]�Z�,k�uc9~��̨�s�������U�gQ�؃5��p<s�^��v�wN�l�\��2׾QIՌJ�+�E�4pkw���>��t�5�3�?�mu[�����\3�ힽ�n��-^��9w��SiA�{���O`�Y��S7է�o���;������b����E�Y�i��/^v�{Rd{)i�v9P��b"*;����Inm���=�`�L܂3�>k;/�n��ީfT������9.
tY�D	B�"6�uBĵj�4�-v)�,�*=�a8�vlr4��+e:0��s��gJ��Om;������������}���>�� �����%�uĠ���6|�1V�"�ׁ\h������td|k�9	�������ن�ys��?h�BX��;H�)��)�E�.9�4����r'���g�Gڳ���5^u��*u��W:�I��=t)^L*��熡j����Ւ�U�C�0�u��-3^�)De�ɪd8�A���0{e>�	�=zz+�ߚMг�$㋾*�
��̦�ְ���>����6_S�WQɯuc�T�9�y��>e0Ƅ�m�2)s�X�'�Z�9/L����/d�ʞ�Y<���w�^V�0B�����|����΢Ú��@���g��	�7-�8Z�w�7�k���9@R�ǜYr���0D����4���S�%��}�Z<����v��N���O�w<�e�����B��"/ʩD��y��g�W�숉���Q�F�˫1oLe�m9�L�h<�H~@A�r�v�l���jBs�Cˬ��x<��4�5!�8�F��{Qx��3`�׳a ��,���\�(My��)�o�*���<W��HQ��h���{ŭ�0s����6��A�������K&{�C�۲��:�R:1�� C<Vq�ʽ�{���;!Y�J�@	k�*��
��S5t/q�W�Df�
�!�5n��U�(��HK� ̌X��S�\���V�){[�r
:��#*���|��1H�|�?\S ��XG�9.$��/bj1���U-�Ar����R̡G�I���O.�5�y��ë3�[Q�j�x/<0G���^��6�sP~"S`��=�-���B�H�<|W���6��`!|�~�/��vz`���i;-Ѧ.X�����t"��f��؇<I~�)�gEH����5�վ;���c�:A�$j&Y�X7���b����f2�g!��DeO��$��d]ybWI`����a>��]���������ݸk6����=�~#�U��B	�a%Y���Rt��T��tS�����NYֻp�%�����fz��CK�[vb���wzzAcXn��N�ʮ��Z�O̓�=�^�DvМTz�p����N�+q.=����yy�kP�5����uch�0-{�(]��˝�N�*��z�kE�����`�f�@-�E���ǵ�8.#�y����]Bl��\�4U5_NcU��,�Ŭ�{w�0%��)ϕE�-=��N�g@A\9��y@���;����z<�o���rmxU?���j�nt\ou���kPӎ���ͥǫ^	�S�y��K�SNe�MY
\��
���U���'H��D���Yl�J��2ƃ�$�u;y�
,%��b�n���Fw�/�5xw	0t�@Z�uD�E,�CP�W�}�}_�  �Q�ܡ#Oy;W?��m�ʔ���u>XF}8�	���,Ľv8`3?����Y�z
������y�E��P����v�Q~�^=$=qh�1^�:οY�X/���rQ��q������{C���\<tY|���gsg)}�	���T3���7�dgn��^T���0���g�\)�>0�~1�)=z{�9��I�Zss��j�K4�������3ZG1��P��ޞwyll<���T)�|a�?�x�T�9P�a�5������5����33a3r�3��1�����؍��}�=[¡�)�08��a�y��O|���鴩�n|�3��u%Q^�"f���ɭ(����`y���[�z��x�
i.�˩*��dv�l.ЙϷ#����5�^~��bY���ebQ��q���L��n{�UM���i:r�|�``Z�.͵/��hAz�N��D�7�E1H�jhѷ��J̩:�f�����L����8����҆m�N�	u���fS����$��S�^�_\�v��&&�,���5��/|�h��]����ț�����;��Q��O��琹��2bW�<�P�����<�,ңZ����8)[wb�P����2!�6. ǣWR�52�Z1k~�f��Ӽ�w�Z���Z��[8Mu4�b��rେ��΢-�2>�^~y��_�B��[�m�ƭl<WVJI説�B+�fQ`��1e�Ͼza�!�"m	���C:m���
�b3�/K�]\�2䃼�L:���)�jM#�#4�'Ǥ?s0h�<�Agd�arHp�w ��"o/?&�o߫�}�r���5��y(�zO��ûP��v0m���wAeM���Z���Ky��[�!;B��t	c�	�k�	>���y�s�UR͕�n��>�`ӗd�g6�祵}��Ν~�����؈� f��L�0�_[�]>���q�|����9\�&c��5za\�N���{��9�Y�Z�������hGP�I86��0E4�Q��c�̜F�Ѽ��V��-i�A!��L��A�`��?�z�M�O��u瑇:���c'�KEWbg���R��؎����B�C�*�-?V�c��04\sO�a'W=8�nz޶uܜ�qoUt�vr�����Lӽ�rSl�W#.|�1��=��*��-�=a@� ���B�:әm���ʶ�t�ϫo6+Z��^L�� Ũ���3���8ʲ���9�������(9�k��;�t�ͳ�,��u8���ի;}E!ᯣ&���@��u��������t7�~�s�q����gG��!�[~�nOUsl�&Qo��v�ee�C���]^{���J^㱫�nk���4�Z�^F��l�ha�g;��h�w��E��_���%[QZ�kZ׿>����E-�������frA\6�����fB~c��r����uk=��|m��i��]C�;f���̍y�����͠����2�1<�5�nL.z��A��r��
1*�5+fs[NXؕ ��鉞����d�Q��uW��47���5�:N�/d��'�ǒ������
�K���m�Os�\�Y�TS��8�Gd[B�Ӎ�>5äH����3Pk8os���ݳO��ۆĿn�vA�,p�a�E���6 ͗�|��� B
<͍0�'홇�s��vf�_2�|�,^�-��]��*Rz�Sl���Ӌ�F���.+�AYZ��o�s��_.�W�h�.u�~�Ԙ�s�Iц�
�fW<5xZ�E��T�49m;	O�� Oc��g��w���/gݯ�K�����!|z~lq�*��\��f���c��­t�����D����']���j�oz�+?Z��+��g�[�`LhOH���q�jéX���V�k1ξ�mZP9�ߵm�2�K�<	�Y��L��k�_��9��e��Xkw��k|�,1�F��b��]�o5��U�|L(��'��q��\�-%֟o������#�$����=�g�|t!�w���6j<��'�b��\���=(�
{E���0�i.�bqcl���WS�z�Vh9O����ׅK�������TUl[lV��U��{��{���UȎ-����#�k �����4=�g�+zz�����w�~[iskkn_�1N�s���P�.�8r�^�0͸��4��c\ŕ����y�c�{��NS2��{�3;�p�m�
�e�6��f�ȲkL�C׊��r�v�tE��tM�1�ʎ�ő���у�o��e� M�X�=���j/��`��̈́��P��roR&D�撚4�w���*V��k�pܫ\��LT���?�\��|;��5Ţz�h��B�:�2����+��w���f?u�6��D�z�8�}sk�΃���[a�s���K�;R��JV}�Nj�k�S>�}�
��FG1�Z4)=���0�=;�X�i�J�?+7��e��
����<}����N/pd�'Z�A�΋<�$-��5B*�؍�ǡ�����	>���a�幵������=�xc��D��^�3):��d]g����4�c��pC�Ls���k��ګ:�]؝���ͮ冗�r���N�f):a|�Qu��LkS�g��Y����[4�T�v��=��e��qxCM��h͝[�l��Wo=��o�����t�|,\^bʠѻ�A���y����ve���&�j��X-[|�;J������7{���B)�����Y�:�x�$��rݸNLn����S��'����X��U_�m��mQZ*�6��� f�f�����0a$�;�u���h*/��8i���{gA���c=�/׾?��{��0���K�%?X�f� �)��$��Ƶ�%�5'��\>���:mh��l�/�zY9�\�����y�+rr�'xor�u�;������z�U�߱�&���~|G��4ں��m\$�d�O�˟�;N6�B7�P�ҵ��A/r��4��f����7p�DqvYE;L��w1e�5p:16>3�z݊nPU&6GS�gӏ@��j=��hņv2`3k��:�O\��U����/��V$�#���L��́���*�܋Ϩ���;	y���Ūq��I�x�a�>,غ��v�8�a;Z���D�}a ���bvl����t��23k)z�	��E<W2g&�mF�췯vT�-~�[���8Lp{�C��?��ʄ�^=���9�i�V�`ֈ3y�T��+�5K^ܺ+��p���z���y43Ht\C��� ��/�J��&���Y�e�Wv׍�S���� ȅ��RGh=f�'�z��C�S�-�ی|�{�&���jx��{O���緦a1��~�����ZǗ<��#�4��Z��j�x�i3&��8�ON�ݧ}E�������%�z�f�L-^N\>x��L����-�'m)T�;f0h�dJ�f���Wh�n��ı$��$i_z���0b8[?���ϳ�0e��mX�Q�j�j�%@`�`���7��xi�c2B�L�\>ڭa�~ڊ��%6��(2kJ%?	]8G�]�0Z�OʭbH}�o��Y��oҹ�M���%�����7�9�"��[W�� ���d_3L������|f٫#-ީͲ��2�s;���l�����Ivl�r�g���&�Iz�%:>Q��"���Lr���f��� �eۗ���{:�1e�Y<�K;7Vӫy� ��f��^��͵;<W�f
�'q�iRN��ɷ�{2z�lݖ׺�ڷ^� �E_�Ú��LYz|�>�� ��Ȅ��gM��껨znxI A�w=���F1���O� e ���4�E����xG�>05��?o�~~���ҙ���MPXr���ۚm��խv1J/�[C�e�%�ޥ�:LK�G�1��y�Ӳ���Է*yG{�kj;B�u��P�+�ߤȦ5յߗ*���#&�UG�ʪY��-ݛI}ǹ,Ryږ�h��L�z��3ᐰ��=��wf���'���8ȥ�u)�S��{�.�Wy,�V�p]#�v�3Wo*!��T!���2��LZa���Nç��":̢�Nf�(��?����#�k@Z�;k��c7�rgssm�ۇ�.�Z�J͟�G?'p�B��k3�͔��\Gv�lm���{G���X�c����d^G��1��E'.p��^p�j+���cf�W�������y���i�"o�� ��d��������k�R��m;lfS6�bX��G3[TZ��h�d�m���f�����%o'ccos!5��Y7^;����OC���~q��׵#Y+���M��F�Y���D�.��j��b�	��tE��y���!��q�ߚ�L$���n��lvÞ�uܩ���Ϣ��3Mi�]��N2^�e�}o�*�-?V�I<bK7��	��5��N��m
�'��\�5�z������CW�3��3gW���{�]��)�r�m��n��;ا�A/>��z`n�(%{QV��n�+�'���s�A=�T	m���w�,�2�fQU��g_��sW�����X�N29��N�l�\��2ױ�):��<��\��dVd��|��R�J�aMK�q�uEë|g�"z�,��;e�p�})�5�<D������[��S�1�E��(���IP�`J��Z�d`�v_����<���z��׌�&�NM�ȱs��;�/��o��wI�ˋ�LU��E���7l�;�0�h�^i�hG8�ǅ�f�&���v{�~BvB�l��˽�����O[�m�t�n4��zk��C�~�O�����x����o�����}�^>#�UOK�ۋ�~ók�π�g�έ���Ǎ�Mז����X��m�]���7��f���(����L�Lƛ���a��o��m�D�^2�9F�qF�͝'[q�#�Ɋ�ͦ�*v�s�]����!r��ܙx�<��y�b5}*&��Ќ�e'-y
��6o�E̋5�;SJ�,YJ�ѝ�Rc�e�qƱuM������E����u�L�7�8ܳ�7;i���"�D>��\	'�ؚoX�5vn�W�8�}�*���VK,���N2�=w'Gn$�='��A����.�@!�ɉzOg�qլ����ͳly�A����r��Y�y�Bs���[��E�9�=p�{�W�˒y���´�����5���e���'R�r�e�E�l��Ժ�UϞڭen.���E�^�\�lz��|��}è�B��6��qh��˺�3w���=����|{��+CPh}*�J̳���*T45�t�fS�f��e��S*�����Uv�c]��l�d�-�M}���P��/&�Z�ϱ_hR�n�Dr�N��4�!���^�;F4��-�j�N(6ZHU�J{��GFjq��K8᪁!�᳹JH�=M7�i+�Ky�;��VHfԖ
:�t�%y?�At�6�G����Ӻ�fz�ec���8$x��(gX4s1����� �9Ѭ��D�XE��Z<���Ó���F�tf�k�<�:m�=��6�=�t����U�=1⢭���#;"H�Fd�!"����9d����@��1�n�4�I��}�{ԧ��Iz�2���2/�I\gh2﷑�4�Jݪ�K��2��n���h�s�/]�/c�J�/�ači��Ұ����'��NJ�?����a��{$]r_QX�A��&���{��,뫦�;��ک�Q[�4�w*γ�ow)�鳶�(�L���է��Fܖ�=�7`����i�ϧf��"��-�4�4eDM����Q��敻�
S�X7f��h��w��)���L�(�;��nz��rSK}#���v�m�`�4�Z���p��//��v�w����>��,Tv�&�69�M;�
��TB�V��YOk��D��7i駎�*[��WݙSy��V>x�&��ɮO�7�^vУۚ���^��qP� �!Xgm�sx���oz�x�t=\=�_s�^J�['#gDt��JCXO�+��х�m�r��N_W8�>�g�1�㭊;x�7}����=��]͋!<&Xі�T��z��\���A���`jG`+m���i�='���7�E���	Cv�0�*zm`g�gejIҫ�EV����՜�@���%pT-�oGf��̵��1p��r�ݼL�8�۸��os��6�뛰h��96���{#�A���ׅ]��p�i�2z{�9�Ə3��{ɓK���s*����c��+(�r�5`YaW]M���8������?�����ߟ~;Ϗ��~*��D�m�f�ilP�уhM�PX�� �DX�F(�QFƨ��(�iF�*dc!(�h��#E��cQI��Y1���(�Q�**1�F��J#2�%EF5A�Tj4���cm�$`�-����F�#DZ5�d�Eb�&ŉ-Bb�h��D�Rh5Eb"ƍЕ�Z+M�+Eb�lE�A�Am��F����>{|�|_��l�r��·9Kn��w��x�����r�e���eo������[f�:ْ�Y�3�%��Ź��������Z5�[�[X�d�b�-�TUڍ�+b����7����3���J��Z�(o�1;���z(��R$�L*��熠-\��eIc\����n�n���q�N��Վ���P��2e�-�"n/�ΠԊ'�d�⤰"�O1��Z�%���2r!��}���(+?�h&5h�%6]y��sL	�zzG6�q�j�J��d���ط�Ee�����k�Ћ�XU
�bټh�j ��s&#���69��,�y�G���?=��^t�Y�Ř�������e��T��{��r��nc�,�j�C���:a�8G{)��-��nn�Գ.s{��hj�L(%����f�z㾪�<��l��5���R�4tK3��7
�T�BP��0�_Tm�19�L��Y44�$=�˥�A��e�b>.�.�\�N<i��S8G)���p�s�!�8{�I�ME��_�a7��ٰ�yj� \����wj�"�s���/v��ői�c��C���ä�b�h���Ʈ���ƥ�B�%#��Bk�)V��٧[��ܨ5�܉�MAW��O�5�����/�#�D.F��2@?����9wdK<{Zvj��j��<�Q����Å�;Z�GG0�7ʚ��g`�P����V|3{����~N�C��g�|�;+��Xa�C/�SG�N]�y��w`�N��}��u;���O����!ߗ�J��ƐN����]�菊�b�ގ��}����}�}�m�֍lm6�R���kF�ljiZƱ��Ŧoy�{���ΫID2������؎k��2*�hR{
�ݔ.���|i����v@�6�8��l�A1mއV70OHW�^�׽��Bb�ħ9�0L�ʡo�i���W��?���vc����H�hA�ݴ��g5������3):��,���tS���:��*`s��������:�'f�#�.z���"UY��>��0�ʥX�ƺ� ����\;6>��Մ˩�g�vB�*�πzb�c\p��BzBc@a�o�i;��YU��,O�,+���}�;NS�.P�׵Iw��\<{�����kH�OP�+��������[�:���\̭Δ1�e�dw9�WC��d����ݰB��0��Z�>��-"Nl���o���V�cd�6���HU���+��\~�d�s�A�P9���q��8.��]Xf��Wn��4�ö���M��Rcl����3�Ǣfy��f4b�;��j4�XF�����p���@��W�ϗṔ�yw���"8��Gi/>�7�+�n�e�'z|�>ڪ��;�[��З��w�z`p�7�s�W��}f�~yrC�d���v\����䲴K�5g����7��wY|�"��Z��0!�孩��;WT\O�gz\(�$���Ɗ�ͧF�t'���K�
�d�Iƞ^���4�6@�x�������ܝI?���_�~�	����ص�M�̴���j�����a�2t�!e>�@V��]�v��x!���\H�Se�v3],�Ǎ��
^�BA�HL˶J�����%���@�ن-���b*��=���!�l__��}[3��)K��9O�^����˳a3J�:Ê�o).��^M���:I��aqf����R�b~K;ԙ�yy�젻v��K��8��K6�;(2���RGh=����V��"��0��mp���(��u��}G�g��L?)��3�����Bl^��&�Ji=���z3����Z��̎5��+�w��8��xhP��2"�d���_��D�.��d���Gw]��:"5K��c�<���������FҸ9��sȜ��>�����%����D�;G
h�j�P*��e=�5gzH>���]I����%��.Q,'�٭�BR͵;<a�`�̧pb:��T���f�]OoG*�ADW9Y��h0�\���LYz���=�A�"mN����ʴ�Ž��ޮj.�t�M�M��Z~Y�R	z�o�u��i�H=!�CF02�G5�_���M1[_���/K�+���tfw�ߜ��3tf�	���YW�V��V/�ː���,�1�^�`���G����k{�yk/)�z����2]a���s[�V�}o{B}L�7Z�����wF����`Չι��9P��cJ�ڢ����#3��x+�^����M�
�"��j�+%cj�_������>��~��
q���e�W�:7�s]��E�H�2�?s��������ga�m��=VVe��3a����;�'�"y�dS2j���e'-~�d�ͫ�B��l�LYR���[z���a����@]�.��,�t�D;k��'�����hZ�:�èfAxN�_.�m�XW�%1�l���n7�_d����b����z�(`ZS �-��B\ay��hd��΢\T��+t���gwZ�>�*aIsH��_�\1|k��A�L���0|�`r9���f���n��Cw_^��Of���Y���.��2�ZI���e��OٚE
j~� ����K1w��c[V.%�*�1O���Vc✝eo�;�ъ��͵�Iv���F]����M�X�I �b��<�q?|k�o�}�s{�l/bj�ʳbq��! �5Æ�&�W$5��=f���6Jtcb�}/��6J��a^Pľ�A��cY�L�HK��U��[��AG����n�q�K-<7����/�Y������*k��	@xy���B9����~5���D �]��Cj�4!��L�c�tE�,՞���V(9Ek��`9�w����u�+���ߎ�M۟���w����w�D�)tv
_���g�ʤ}�RT�ק����.*	L�����x����S�X�1N�k���e>���l������ӰS�l���Ծ����5�Xձi,U�mh��7�2�I�K�.׬&D�Ҩ����0��m}k
ax����&�'��н��=oIw-�m��h�ʶ�ק7��Y�Γ√rR�H�TS����;"�{��|k �D�)~.�)��Y��ы�a��3he��.�eJe�[�:��Ɓ� ͗����}� Iû9�,)�i[ogE̡�NhI����}eS���)=X�6Ⱥ�09�j-#�bu�uewH��r��S3���+`��s!��/ C���@O@\ߤ�
7��
�Y��^�r��PX�jW;�i�����6����%��b��������cǼ�NuΠԊ:�N8��E��Z��̪8:Z�n�T�(��K֮݇�F@y����t�}ni�a1��ͺ3�Y��T��w*�3�E���J�F��g��r^��T"�`�j�;���vB���9�W}a��d�E&����]�{�Í��V��.�ǾP�9DԷ5�0���g�A|<�Ν>In:b��^z�]%`�#��f�tw�ۤa�,	x.�2����fN��4:���7��®BfV��8*	r�Kk��sPq��ʘn�x���z���ܔߺڽ�����z��#����goB�od:oG3�O��AC����kz5폴��pu>� cw]D!]n�}���OK~�J<#�>����L������[
ݷ�[����7��g� �0 �$0�Ofo�u}��������y���ۜd{��U���?'2���p�4�*���1���v���l��"mẇ@f`�>E��̔��5�m`n���t��u�A<��o�f���8أ�1��ԅ�P����oi|k��^�
��1x��S�w���#=��}���L�s��g���+���nK2�+<q+�AW��K���tS��?`����a�/&R>~�L�r�v�g�z��8u�Ak\�&UiP������t�cռ4����
ϟN�)��+Ӿ�]ُ������{>!��kw��ȳ��A�%)�j�U�9�Z��	�(R����3:�\e�����E�{C���u���p/W�|k�4̤�Ĳ.�S�7�&7��.d��P��Ƿ��{�g��c>o���~i	ٲ�Ba��=1�"D�i;Ϭ�'L9L"��TK4b3��N��{�\�\�=H�@y���$�T_�P͍1�tt�}��Q�����⬅��f��Z	��W$�w*�K�����'�7����D�~/�/޲0>O��x~?��i�~���H��r�X��`e�8�  @~<<��/W�x��4V�\��Zy��۹1������w5���ؙ1p=�=e�J}�y�E�G-���C{tA�g:cU���=��F�ڃ���+zo��%ڣ��}�XSF4�U�T!� �vkre+5�i*L��L�1�D�.�Q"X�&르��4.��ܡv$�
�=���5j�w=yd�����#�a��<uTq3�K[���|@N�2۞����%X¹t�{*	{��q̮��s���GH`ӧ.&��D�u��U��7��t$:�>ZV$w0/z���������R����N=3�G�Y��a�0Ǡ�K,��8zt|�~�Qϭ�P��Lx>�MY�ciz]߫6C�Ⱦ�_��IŜvuňL�L��:���u�j�5��+�բ-�P6!۹�܆,0h|.&%M��N�k��h9�6�����n�}	�"�-b^����{�T��^~:({�L���R�v�p��e��!�Za���=�Lf���a��)��!,��i��,y+��R]��:�`�-3�U�Ś�|�4�n}/n�U��sv��[d�7\���&�ӯB�g�<U3u���ezm�d�$9͜OX�o
�
K���wz�sg���=n��G�S��g�j+���%6߹J���4�E��ј�;I��|lt�ݶ����O4oo�$��.����`�`��BA�J�j~���Y�$f�?�Ӓ4�Ͻ?YQ�ܬ�Q��h�9j=U1h=`o������{_�M^�~J���4��ʐ;�n^J0���@��e�]����r:��N�A��TwwK�So^G���Ni��Բ�����dS����._{=wg��ƿ;��<:�;�z���4��lҥ4�f�� ��@ �Z�Jbg�%S�e[�X/l������d3����&�Iz�N���͏F�U>�PY�fn�q�Ws��S?�#I���v��66rS��f�t��sӳ��2��M-�bz��,Y��us��$�m'�\�`n�F�W0�LYv���y�[S�	�s@1�D�	޷.�Sus�+wb�u��2�6a7C�zOȀ�A/Z�H��3L8~��`C�=(�o;Q�Hkp��W+�D��:<���y\���۬Vs�n׆x ,��e�~��'�q�yď��k9������E���B��)��wf��S�+�X�"�׌���0��FM��W>h#Nd�Mum%�QG�����7�]y�_��i�A�A\��./>�m���?>�q�j�Ja����;m�����`q߾��������h�e�q���<�&-0��^�'a��gµ:�֡���m^�4�}�a^I�v׼돏^;�a �re?�p|�lD��=��Aj��Y�u�=���y
l�	�����'��=.Ť��q �/\����`�?�����s�h��6ϡ�뮡=|�\o7h
�<���޼1�-H�msДϦ{�/
�q��u�x�+��♝	�6��P�1�-4���(��/m�{$�PyF�5]��~��A�������>4o�.z����CK�����^/mk2Ȯʽ�r�>���}�q;͐N;��|�"b����6۬�E�f��$�PJq�j�e����<��3�55������t�o�1�`� `���[rx��O`�Z�] ��A��쭒���z��'=GLFgf�R����m
+�ܩ&,s�9��@'}�mAt����	��Z��ck��PgG>r�~�C��լ����/S���ʀ��ϨR�+��Һu�>:�RC�f^���P��9ծ���61*�UԻ'����q����A�n�|��^b��u�p��)}3���E�2��9w��"��E8��aլ#�E��A�4�t�Qf7{`(���h�3rq]�
2l�{,�4�v�*S./1V�Qr��/�\�;�0x�.;��:�3D��d��"�s ��\C ���#�)=r�d]&09�4����fg��v1�6+�>w;܌�m/�%er�+hy�!�z��No�n� L$Qpޅ��J����R�*xMM�{�;/���r�/��(�=�Z�����D�^�'����Mг~s'_� �G�N?~��/7��k��>/�xF�>�����z8:t�L���|���SnU��Zz��MI�n�f��n���t�B���Ф��p�hR��q�PaE��w�>�s�����>ҕN�u6�q��Gr.�]��6G%nۮD�9d�ӽr����������l�Iʘ~��3~
�XHOv[��PX0l-=\x�<�>|�̳{I�kַ��v�[#���ltT�֪9���������~%�k�_��ZJc�e�Z���#!��Τ����R[n��P�9^&���8���g2dK�Ou�j�e�kOLE.���l�۫Rͩ��Dzg��Ey�#Cބ�������}�38ԑQ�y�~��[=��;�p�C�|�_W�m�29�L��쇝0����]�Y�PU8T6ԓ��ُu�>G�Ձ�g�s����	C�O�� �����+Zh�:;���
������g>G	W�d[��r4W�5曌�M���\����������r��ݑ-R�K�w�]�{ysS�_��b�e
6Ty����	���5�L��&Ɵ`�,ʻ{6�S��h8ǦH4��ݝm��-�^�"Se�W�*��vP��Ӻ�5�E=��!S���*#u��E�d5Ġ�^��6���|���!)�g��(,wT-�.� �o_������{}��?���������c�Mf�XN����Ö��n������9yX�t��L�E2=�`�d~��眗bk���إ�p��F�������#�ޙX�e�.���GB��}n�9��������S$˹��PxFT阜=N�8����۷VPʜ΅(HS�E䗘R���W�@z�W�����Z������%���7B�mf�n�=ǋRKO��]�\B6����]�FwClM��t(z���ӵ��2[[8+��ٮ�G�lfM|9��ˎ#Y�i�%���Nr]]���ow&w�]��G�$,�u��(��ѩ)���/�J;�z�Օ��n��&�l��E���_B���^X������}QuH ���rK�5�X��;��v1>b3(�.��s�`|g���q���3�z�j�#�+�)�p;�v��添e��	��#q��e�-_J�ːdG.�]lu�q�U�:X-�jVԼr.��Iغ�J�y��b��w]ȳ7��NƧu/1:��W*�a^k�!{N�6h̯����|z)1fo���6�w���5���ph�v��w_.��m�<�7���d4d���CE�Bm�=�ܨ6PCC��_"|p�� ��W3R[�<֓�_B�2�p]q�}���knU!�a��hdG1�pPw�p����ͥM�U���]3@ؐ�y˒�:šf�}ܤ�i��m#��5�t�	gxǭL��7%dGe��㞮c ��|j�yޭ���zL����\�{i7ǅ�X�0[*���s9L�ӄ�=r�����,�"6N�y���s�T�RUn���c���Js��bb����/�m��w���oZ��%m��~܋"���H͵����-�x{=����'A���pv�]0��sRhv�\�3�8�
\��Λ�ZE����?y��+�,�y>f_H�<�z���li6�F[���O�c�� ��K��zaדr�4���]��\_c������D#P��iRI-�!`3/���|k�3�t��!�%�dr�'[4#6�f�|V��e�_���&Ɯ����:�7@Z3�ܧ�����N��n�*1mʀ�{n�=�
�����+S����Za�����Ukx����B=�.�)˔`V����ly�e��6�Ӂt��@��'g<�{��VF�U��͠�F�C���Kg8{u�s6�)�%P�zi��&d��F[x�K��I��ʢ!7�u�����7-d�(�I���ge6*�O�����s��&��(x�&,I�ң������-���W�b��oL��\k�ܚ�^��9�`{5��>�r^�[�}��/q=-��v�}�'=u(!���v8�}���:�*LB���G��l�tȱ�4�˲b���,#9+;�q����1X;q�+Nm"@�c�GkL���!7I�%�;�#w$�ʌLZmi���T��:��,<�c_;Fܴ�:�E.�'G�< p��+N 0j��#� �NC�(��`2����3�>� ���ũ(�K�Ѥ���ѴF1csp�j+ 拥!!i6�h�h�Xlh-�v��L�Z�ܰ[Is}��nn[�5�uw\�ەs��N뤑b�+.�Tmr�F�E&�R��tAE��	ΣZ.]F��b�5�G5Ԩ����dDF�'w-��[�sQ(�Q�(��L0RZDѲ3n�1�m�ۑ�#lh�j(��!���I���\�h6��o ��}ホ(�
���D��?k�6�e�=�ϵ����Zx伃�t'nR�%g^0WH�ʝ���C7���Vᘸ�ʗW�ꯑS��6{�b�x����x[G����O\�_�e'X^%�t9�����a���a���'�e�{��0N`���̘�����a����18D�Uf��يN�C��dEW@0qe\�Ʈ�#�S���g�#���^4�:�AQ�8g���ٕ��W���z�U�f!;����Mf"�)#���4Z~k�PX֩.���� �����d/������Z�akPw�Q��s�j;y^9S�l5�8��UzY�iT���,�� �8x܀��:M�&��Z�$�[0`���eʝ�m�z�[+���W.��S��.|�:<�vퟦuЇ�+��p8��~=.�C'� �,F�(�����B���[�Ԙ�eO���qɈ��j�C�k��Gks�!w��I�Uņv�`38!@}�����P���d;m�"���zHuA����6]��s�2HwEzV�����s�]�,46
(����t�q��A#�G_�Jl��z��������@��A&a��o�؊�ou�g����2H��Iϛ�F�R��sQ"<����顼�k�$�7�S��<�u�{��OrN�Yv���'H�;A���z,n��mh����r����7u������Pm�e��K*0�5��k���S-�}ur눶4^p�ک���|E��`�-�nMTn�:)5�����4s�9��où]�?%C�}�������4��B��%�<�M���6��Hזx#�Z��p��><�mtk��-��g��}Bi�>��{3m^�J�����,�`Z�:�f�'ƚx\[]�k�چr��w}�؅��9�C��"������^}��"Sm�5���+�(�x�xI��3�q��\��~�_Ui�P�/!���-8D=��VJ�j~���Ⱥ��ñS.E-���:y�c��bUԚ�Du�5���JV���ϓ�'2'�P�xA}	x�cN��Y���m�w�7����r����D�T�b���������_O�2p����'�M����/T5k�?�&�Obw~�l��Al븐;��O��zm<,�t�41W0�%辇�����[!x���a�dڇ���k���������A��t�R|*��&�~OI�5ӊ޷���f�H=�j2�w��\b�D�N��!��!��_B=p�'����L4p�/<�|0v�I�����!:6X2Ȋ�W������Վ�/,�>#��y�C�~4�
�W�2)�&����N[�O+��Y�i��w�晴�s;(;܊[�h�	{�\V���X�m̔؇��'y�E��������z�`+Q�3Q�D���s��$�n̅����f[��3��i�s�N���Lb��+��S�J�K�����)���=��ˣ�{���~NG}�*Y��[�2����@?�v�E�z�s��\�S�N��vg���zf.Q��s��O�l}N���-��t	�d�qO��|QӞY;�Gy/ �k�f{�Y0�'�l�)mjpo���
ZmY.&������-A�s;>��ıs�i'Eэ��Ǣ�[+��6�&�c��sϰ��Mq�.�;�=��hU僔��C`�gWX���]��غ�\ӝU�%��i0u�t[m9����4�:`�nJq�nF�[�Zr��S�Blzʴ�fs�)����\F�'X@|�k/sW>����Al$W�BZ��!�d�檡[O(�
��7>����z��+�ʒ��x�(�zaS7 ���m����I2A�B��l�y_�a��\?yem�_{л�ZE�^�c$���3x�4���M?��i�UZ�e��ػ��`:߹�X�
P���л'����\c<�%�!G��9�m�YͿ� ��<%��g��e�,�/��nwL��)�%)�O�8�}�Ы����dK��Z׉�}�{�`q����Ћ�����zs��WH>J{����[՛l�Gi�~:]/������=��~~�S��*�w��ƃ��_�r_�O�zKia����7�	�����*�Y�0�u�O/����饍(n�KO^B���|ֹ��7Z�pPE���9}�},�4�b�T�)�L�8M��\�2	f�И�=;���F'�fO{���\�Ç��pO�= �������Aʔ��r�d]`c��l�ރTL,�݄"��Cw[j��;73���<���>�!������n��I�Y��K^`J��,j;�����R�����m#�ŤOjX�8sX:nw	���k�Ֆ�='(Y�L�"����}u��	7�ӌA.���G2�����]��� ��~�姠!i�?1����i��mu��{�23GL-�1��r�}~s+u��+\�%锾�GlN�{�96��V}k��8������i�6Z?.��ۛ����:�t`�,9�� �˦��ܡ�r�&���q`dl9`�	f��?�uD�SՇF�����F0���C�u��T��z����m&Y�^���4Nө�-ޞ�y���lm�b��ť^1&��H����ۘ~�wS0�/"�y� ��8i�T	����t�!���]�h�e]o�lg�`L�\>d$�5�m{��װy�`��-���-Y.���qw:��p��]:}a:�bP�e�f%O_iG�}�Y/[6�7����T�^W\��:��i�,_QG�����ZN��{�潑��c��y8��ڍ����b�[�\7u��)ڝ�NI�k�ccZʇfq���c2�:�z�3�0�t	��磕}s����y���֮���w�X1l��P��8�sE�p�\җ��]���ޮf;.��[u�km� �veK2�J�8z����Gծ���m�k}��UJ�z'w-֊%��˲̜^t�����	�G)	�ZT)=�We=�>��xm�l<G75�[[���u��� 4(M<�t>C�3���CM�j�B�Yx��(LEP� nWr'�����q��l�5������/bf~���E���
�&8yP�8EoW�gL���s��r`(��O�<c�,(�qOw0^���A�l��.z�CD�T,�w�������y��K�z���xn�gi�Q�NZ��kÇ�A;65�8Bn�<��jy=b��&2�莽�(��wBʮ��j-?5����j���^N%�����/����dc�ʿ՗�O��N�߽	�ϖ>![7o�=6��a9B�Uz#��XWC��di/N=��ZUd�y]xm�����"�[��ؼ�ý%��	N0�˥k߹A/r��8��,�'���ﴎ�H_H*�Gz�c7��l,�M�QЌ�[2���p&�1�����[�d��p�s-bX2����)=��*ɇ�2��	� g.����P�ܘ�y/�t\���J��]�^�iI��<EҊ����4s���7���׺�:�u�ǜZ�_�}�53ݣſ��/��L������x��U{���ʤ�'�{�gӏ{Z6�L��Vm>Λ�����7!=^v
?O0O ����jj���d�Y��E����Ą��uE�S��0{uz�: �@ݭ��oϡ�uv<:%�<���𸘕6^����Iu�ۗN�>��ݤ���YX�w����x��?{ަg��_��Muc�?��2�r�/�������6�U�mS��j��z/\�ui��L�W�[��J�!\������B�}Ń2��~����>{7~�ӕv���������/\��|�[����n���*����9!�"Ӯ�5��^;C�~ov�\�����삒``B�,W������AUk�j+��Bl��0�5ZSI�g�K�W]�"�x��Vl������*�V�*��xy�s�`��[��2�sS� �\��l��ɫѡU?i��u�M1�*4��Du�5{gOMn�$*$�6T�&
��D"���z���]Ԟ���/ק��Q��˼'$j�Lh$i5��ܞj��\:��?�f�����k�����ŊE
�]�6%��YYF��E'�tSʾ���X��F�v3�YY�<Gw]��7#ƶ.p��E�Wh`�F��翨�ʭ����Z��;�5������,���8�c��:����Ž��!��C��a﹕74	K4��w�B>X8�-�7�0f���(wK0龒�'M*I��Rr�7H�X����*�6�,�����=���)���Ԟ�D���M�ѡ�|3�ڋ߰�v��G(����K��3L7��O��"�滙�5v�H0����`����q"6%�=��n���mk�0�/��]! c{<�j������s�?�	����R/_���~=����:�r����/o��ƻ�)9cS��/��=��V������T�n}���(lw�!����?�X@A�y�mt^�=ϵ�hZd��R]���A����$�����1��]>�2�͠��}�CX.Aun�X����k���!�qz����t2q��sL��0�N��i�{�@�b���Z��w�xg�h�gi�����vd��o�(� "c�������7<�Ρ4��^�.Ť��q �/��y�����nsB�ʡ�7vv!��`qc<>����m���>��4�5�Iv���F]�#F0w�ܲZ6��\�{��K�~�9}����PI>�	bI�#�ql���z{3b���A��A����:6�:�����'�+��.s � �egWYJ�ˮzi��ǔv
l���D����v'�q�3w�ӋEg[� ^�.��������uR}��^NbH��7{k�e��q]�hs���e�`��I�''��޾�/�_Df���t���d�L��m_���y���W��ʒ��2�?�S�Y���.{"�|[YQ��k��'�3y:�_�/���F�sn!�y.�g���^��5Ú�΂�pXs�eG9��1�����P׺�}���K9{�@tA��r�N�J��J�*,)�vN7K�:�q����(�p������
q��s!eRf��xX�^��E�-��$���*�J��[�[�h]�f�x�ׅ�GMi�E��C�[L:!��6cW��C_v�4�2�^b�@����=�t�9=��*-|��h��[N��ᄎ�B�>�A?P��Az`K*���NT��|��TVt��	\�D證7<�2�-!���~g�mA�א!�n�OE'7&�Q���
ܬw�z�J�;��:Gr4��ˮw�J_���{���>�,�=	�~8ts���y����	�u�e�gz�:l��lN㋰8�,(]<�l+�`���g=�O��(x-= !i��/}.ab��fӖ�Mf�p�m�uu�`iT/�Ԭqɺ?���K�W�N��j����_��QQ��;��E��d͏��[sݓl�h2�������r�*+����y��̫L���Z�U����%�k�>R�'m�nP8t��6#�ۋ�#�R�YX��x�*�p���\�uw�F6_\Ϡ4'X�u����(E��ѵ�<�I\�GF5��z��4C'U�Z�o��{�,R��_����M���Ia��~e����N��Է5�1�A�ŕ��8�w[�o̽��]0��p�����omu�B~�}��u��`A1%ڀ�.ݯ�&��ݍ�yF�T�BvU�-�x��`��#^]���@4<����������w৽\�C����7�@��cA�sG=�-�{�mᎸf�`0&|�Yq1�)=�5�^����\����2�T��?m��%�_�:�W!
d\�[�:m1p輳�, Xt�]�E�K��X�y�mҵ�΃sJ��^�qeT�5{ǌ��`� ʂ̡F��p��8�E�T9�6)�ԇz�
��d���т�]�cK/h���q� ���ޘnnr!5���ekU
Or�еј�v�$���.�-̎y�x�}gh���i�q(>W�B�||�jJdY�9���5�^c<d�@]Sy�7�eoK���ze�BUe�m���o���-�$2^	�_M�O�̤�8�6{P�s�6�sG�;W7S����i7�s�8��s	���H0͓��.z��ƽ�H��-n;r^���+z���&�gݘN�v[�/��F库ճ��p�f��1]�k�}��{Uyx]�W�xߖn��'}Q[uh2���`��̊�f���vXo��-���m�:7���I������"���GPɾ�Vuê�^Je�;rU��c�joT��[�;�y��q�E�7E1�]N�^0i���8nvm!�li�r�6��^���C�[�*��zQ���]�B�󨻊�eWC�Zq6�9�(�5�R]��'��찏up�e�O�8S_
�k���z8Be@I��7�3la7"�Ī2�����u�9�����t�lir̩��{��r���x!AB/���h-���*������t��h���Z�T�/~W�t��q�r���B��z�3b��vCC�<�#��6�k���/zm��*�����V���.�o��VloE>���vK1��}�%p�	�y"�g���˫����Џe�R;+��26n��ý��F����I4���W���-��C��t��h|.Yv ����C"��v�27;�?N?w�f�0���C׸�$MC�O�P�������ո9�6He�ob����Jژ�ؼ{Y�C�@��L�����PB�)�(p���H��vT0�^�����!��I�y�������bȾ�*~���L>ﾄ���*'H� ���?������}�w��������|�=��/?k'7h	�Vã����R���v��Uqާa�}ϥ��Z�\�,T0�Wl�V_'.��Qَ%hE6/�����o���jz`��{k�s>zB�hm�mcZq��G����y���x�/�!����U��	���sF�k�פn�)�T�݌��kT*h6yW-�R8%��f�{sحz����I>�J��
t�Gd�e��4>��]���ʍsujVd�`9_j��v-Ld��_>�vI�5�,��N��C6c�5�,#ݯN}��*�c�b�Az��q��|�����5���Խ�L���,�����Γ�c�Nf�#_7$^ܺ��V��圍N��/���[�R~���� ��,����Uz�"V�'�]�k����ͻ�!7�s�7V�Ա�WG���S��r��w��5�s� 4vL����\�F�f������@���y:	��;��2��|���7���r�/i[r�C4r�W���¡�P�Db���d�x���~�8�J87f���=���]��=��1�G��Ļ�K��kNH�kߵl�DJp�[�F1@Jx��b�<`�g
8�+m+d8&}kU#�M�P͠�v�[�0�N� m2��Vn5(��[�{���٫���{`f*(���lP�O��QeE�A�l��S� R��؟�9�Uh����Bf��[�}R�^�f�`��p���h���o\e�W��`�6�Iݵ�/D�hQ�Sh����>���u�x�z�HxX���G}����8xa�U�w]�d㹪J/vu���M���}~�00�f�u���ݤ�m��w�z�͙]�I�J�/��qm�@�y���;�V5�g-o��2��,�z����s��tR��`�;��2v��|�f�!��t��_s��/��u8�iN�kEYX ��+���a�{wE�k�-q2oFna�q|^��v���M���uz�z;r�I��������+�.i��F<�x4�Y�>�K��=J<M�Sxg*�*��qf���_Õ�FXUK%�л������ެ��)d;Ynޓ̱{E6v��tW��GK�a����~{�FA�۞�O��<�_wz8�{�Lc��Z��7l��W	�(Ӑ�yB��;Z�O����Ob8E.���۰�R�:4��^�x�9�e���퀠�(B��v�Ӛ��J�.\��1��g�
D=�Ӷ=镌�����/4h��Z�DM��m�y}��B�$�wW�L�0��\.d(�+ ��{ЅΪAX�ʨ;��ك:�N1�-�M���R���&W��\��{ȕFqytr^��1����x)�֣�s%��x`�=06^�>���$����3�K7��`w�c�+}��ʡ�W�QE��[��9�q�p�f렶Wu���Mh��7@dw��R8�]7,���aoq(:s�c�&��:��ۺʙzv'��.7�:�0��������ۘ٘ ����eͷ5�I����ʹ�d�"�ܷ.鍰!��6܊�RjNV�*�(����+����b�ѱ��.\�7.m#�.DIsn�^Mg�\�Nuʍ����\܋:�ʎ��M���Mrܮ��p�F�]��I���wc[�ݹ��ʹ��Ks�7(�j�w]4i8h9[�N�:jtŹnnj��"����ڮ�ۛ�1�̹�ۻ����oʊ�X���N��(�뫨Ӯ�v���6wQW"5 �Ō���o��I�ye���ي�ѵ���)K�guz��K��KX�W}���������<�^Q{D	�� �. �Q�z4f޷�Lu�?��DW]g�y<����*�`����H�"Sm�R�&�E�U7'2�����:z�c�]8��z��x/V�숐P2@����!�v�"�J�k�٩H��=L����B����E8^"[y�4�£I��3z:���<����A���]�+�^k\)S-EF\���#iNk��~w��?�Nlj�LR2������lz�\�� f��=ܪ����?D<�oX��q�2�3r�ܠ۝�Q���T��1��n�G�nIN'�`/4Հ�aˉR�I,DN������=Dc���n��6Ԟ���S>�M��='�|�A/^�ZGU�YWC���Za�v0�p��_��t���i�s���e�Q-ۜ�Z��e�$k~�A����F�}����#Vb�j�C`��
!�c�!w$Oˋ��
�W&E1�&���k1��%o�3�v�NY.2m�¹�yUK6Pطvm�l0g!��������������8��CZ��-����hik�a��e�~�������m��uv�v^��	�g�濴_\�����v��b�TZ�F/��NE�8;�_�摉����/�0��뿎�:	�md�8�$����/��YIVG�G9������ʣy{�ǣ�yt�B�6!�_sr����uh�Q������/y���n����5Է�ݐ����~���~����Nç��r�Xi'�s4��D�|%!�?W�P�e�~��~Qx\�����5=u]�>��ѱ�10u������ �^�7��w�<}�>hOhw�?!�9��`q>k>��+��;����لP��A	�&:����s��yf����%ڒ�d�N��<�M-�uۺ1p��β?~���P�->���c�I�xCV���\��뼧	�ܿ������wd�@iU��]��:���km����γ׳gc�+��%�ǘ�����TE	 �=��9��Q(;V���\��s��L�Ƅ��vO^YX�K�Y����eEÚ�΂�r���)\�OPrq��`��<콻:��##���C&�5�N�)��,(�vL5����FW�N��q�V5�&���尥��^3]�^�1И��Bd���s�*�IN)�-�<�������x��-\�zB�~��O�6He~��b@�2�#�iRe��&*�t�/�j3�y,�a������Uwu���vl��6��!���NH� �������l��?��kޟ���M���H~]�gF�Kx�i�shF�d�2�>�p8���G�Vr��Jtg�����������m��Xi�������97�$l\"��V�[� Wlܻ��rT�j��#mfs+��ѭ+Ep�r��{}��]�ad͎&�U�{}�-p�~��q�}�rЗȃf�-wb��OE'6$�
7}m%M�z-6y;n˹�E����<5z��/6
�}�lD|RD��k����yW�>"ę�/]�vU=�ڂ�y^9����N8�*K
[�MN0A=�}j� k�Ckrܫ�&�V�Hf�L���A�S[(ʄ�m��VaTc����)k�Qe픿0�v��W=�~1t��+n�W��&��`��6�@~�5;.�hgQa�XR�l2�{���9@���{���.����୯���B��>H��Bp�4Ba����:͇m8r�\.ĜRS�����osw'h�]�.��;=\ŕ���Ly�y"�XE�����fKO`W�P�����h�Gb�)C�Pn]��.�xc^��0��q�3%'�0�N����kp�Fs78�1NYQ�7�Ps�{�}6�%r�My��]6��tS?{D�����=0qB}{���El�=�F5����w)��Ȭ�o�*<����q�^����M=>��(��fݥ�vT�X؟pc=�g������������<7�Ѣ�� �&S��I���#�y��=���s�w�c~�r,���y�6m��d�5��7�a.���[��D��U�T�5r�]��	T�sG�t�c/�i�/yg0�u�����f���b�{�̽�`��r�v-��ږ��fD�����b�)�Wm)�_�S+>�����>��ݟn/�*��.�8t[Iq$>T�HM�x�>��Qb�!2�^%9K���6����9�c���P�л�l�{"����^���Cj���b���D���e��F2�P�t̝Ƹ�;�����7E1�i0�?Er�*���py������~������3qa0�)�x��)us�����E��=��ۋ���f`���M��,+Ts��j�&W>gUI�
�� �3��+'qU�*��E��%�j���A8���N�8�eZ}�WfÙ�c�&��D!�zvh��	3lP�r���˫}��^WC��di�tq������\/uc�@U@qB`���@p�_�b[V�����қa�K�k�PKܾcI{e�/�}��O]�/�R�˒r����
�ØO���h���H�=oE6�0�1�� q��{.\Q�[�Qs�n�O�t�q�3�v��1a�����s��	;�s�}�n}���u˅t#�m���SB����+�q<$�c隼�53�=w�o�pf3A�ߺ5Wo��/�;�;< JNǛ�We�&�"����3�GToQTU��v7�/�US��vۆ���9T�݆�:fI(ʅ^m};�{/�L̼%,�N���g��dV�𫾞����0;���������>�-�����lZ���g�]�����B�[T�l�Z���mJ���b�G�A�skCrC��A&[��_E��
�.�l�>�g��)�\��f����`����T';�~��fnf��d��YA
�%�<�M���Z�L��ԛ��Φ3�)�
yg����A�Ϗ��&=�/fq��.JY��J�,�`Y�{լW����<���TC���|i���%�p8��,9/".=</֮�V�W�o)���
``6Z]��gE�i���[!���=8��z�x/V�(�"Xd��t:�A=øV�4!�q��6{/?��:��`.+�Ĳ/a#4����k�����t�On�$*$�6on�[�����Lk��+��F��K�DJt�D�7�R)��&����O�p�G�����&��r�Q�{Z)3s!K6�o���fٔ�4ʔ���~(7Ny��a��ŗ����թֳ8���ov��� ϜhA�o�]	���Y�mE�
�i�\&��9E�+)�xc����NL\���o[����F��!���`<��v��p�R֋��+�
����i
%=�s�n��Mn:?C�N��3���L�c0>���:U�
�Ŗ-�y�V8�T�M�}�(��Kv�nw�=�
.øc�E�U|�������<�H^m���Х%Ll��}{(��0���|�Ƽk�_��i�9N5vE�'M��]x;������E��ܼq!�M#�^Cψ%��{��~]��N_?1�2��}�Ӎb�il�+w�={ʛJx�k�o6<�~c�NP�i��5��qx.���H�q�c�ŽGg4��/nWr�}a̦^/��G�L������۬t0m���y��l6j�qY�~����>2/Bz�k8�B��RNڇ����B<�Kp	�c�����*�#��V9=��~���<����`���R�`poJ�kz#�ZEϹ�o��QF{����K�X��b_b��S�����D�N�ON6۞��=�6�Z`�mF�\��9:iΎ��!����[cW�?r��հRL`�|ջ?yX�~��f�k=�b��]4���O�ۋ�8Athnj+$����g�oE��dgO#���X03��!��Y����ff�P��b0˜�C�yTU��A?5�� �ncA.�*����� N|>b��~ni�*��V�[���Z���7����~��}�*�r��N��S���>�~��Q�֍ax��S�s�kn����M��Y��8Uuᝤu�;o�{��ه�c���N�k�ZT��l��Fܤhm>ꙛ���HP�kP]y�u:�]8R�?��-�x�{1z�D����!>��v�HޭbϮu��e�|���JD��q��d��S_U)�'�ZJO[s���Jܛ��������M��By#B��~��ū�$�D�6
T-\�)Ś�h����,���H��ܕ����c�!Ƙt���!�x_K1"�˴�M*2�^b��u%Go���KVX�Bm��4�����[�	�  �cO��O�'�^�ʅ�;^L���uMN�z�[2炱�����3m��1��#6�ҹR\W(���}�ܲs���r3���6�-�q�/\�9������\��-\��eIcC�Ӱ�����Ǘ���]�>�?Bh�wb�/��z������xǒ�����1'_%�-�c)]k�A��sۇ�p��c�r��)�Z1���
�Ƒ Ʊ��ͻ��B��Ԭq֟�k�PK�)~a���g�������+~ܽ�{qz�]��	<@��?ĠA�i���e�mxgQaͅ)�]5�|��r�R�����յ��s/����g*V
�A�y��|AKiv~ʄ����۰���6��[5�b���+c���}�m�b��s}��B|t=гoX���.����m�.cfK5y�_�a��K/�T��g�u��4�媉*�{&���@��=��]�o_�����o���t�{�E:��^=w׮x��|ҀI���Ow�������ō������G|�b��+�x2ү���y"�VF��0��)B�epzd��x�z�l4I�L��!�=�7�	�� �w��@:"�W�&�����fЗ�&�gV\�2�
�)�csJ�צ���^�kM�Z��^�J�!^Dך�%�`1p�)���5+��뵥��e�C�ʻG�G�`]hGw+�ń	����Ơ)���A�yfP�`%G�>�[��e\�F?Û���T��Úye���`��!r5��?}bmCǗ��>9��ʀX�Rt��d>�s]�Q۸�����٤
�;�^ǫxi����֜I�&BE�x��|���L��� ��q����wT��]�Hj���B*�����e�'�[�Hql� ���O^��qEA���#f�7�~�����s��Y���=�&�<���'�}h��"!0\�\a���X��ng]E��V�;����]��RtÔ�.��Y����?R�:�
���[����"���O�^�D�ng��zL�c��9b���qw�Q��j-?5����5Iw�'����X�`΅qQ��'ni�[�z1u���ۃ������||����չ���NV�:�:S7��v��,��)"oQ�W�;�S�ϱ-���l�v�����5	��m�����;u��iX��vNY���5$ĮLW"��Y�w{�L�ݯ��C��Ǌ�����ubL���'(Y*L�Y�j���s��{��,8�����ٴ���=8|NW��`��G�8s�ѱ-�D��W	V0�zV���;qB���W_Cp����R���~0z�R!m�xB�tP3@zB8�÷:g�v�|�3l��f�w��������k�{y[�6����fy��B}_��}�	�a1�������kf3q/��5�+$1���������%���`҃��;RQ^Z��u�v2D��Ņخ�U6д�:�ƒx[�p���ƽ��ސ�skCH=��'�!{ќ�E��kt�'���{����(ۊ�����������3�w�g|�C�{��9�ٸi�{ �=)e�/��xH��ƽ1V��v�=>n��u�6��/X:.`za�<��ʟ�*�{&w�Fm�vPe��-��%5��f?uaL�4��z͜OC��׺E;�am^{G3l�=�+b[%��h��Y����{��r�-BҚO~���`y���[�z��xA@����DCߛ�q���w����x��݈�f{�c�I��K����6���F#n<8���e�Z1��]���÷G�������{,&ͭ��A�]f����m����	C�W*�;�9��-�����^k@�}�/n���}��������D�W{\��t��#qN��V�Ք��z6{���%)���r��(�E�$��XTi5�G[�P�t�On� ��7�w�"����5ge��v�֥�0ʽ�_I/])�|"S��SH�kk���ȸt�h�mb��(u�e�cOok�w�`���C1i�Y�m�N����f��4�'�I���9�����b�����|{��gmpoq�����t!�B��&��՝6�^�¥�m�M��Z~\^�J:�!^cny���w�<�	�?O�E�2(֯C��S?Z{N��MɿB�#�T׾���lrxw#Oq����<�w:lw�%ݣcF�A��r��?.�N�\��X7�r�x���Ӧ�ub�r�������jX���>���v�;5�W��?�Z3 f{.�u�6��Z���x�r���V�S�^5�=��O����h/����#��XI�*j����ڼ��k&�)g^���ű>	�~}��B;��K�VhRy���1�g�Hm
4y��U7�̽�n�C�)2�e<5�g� ����χ:D�3Eڇv-�7hջ7F��]8p�ˇ:�"֭�)��Q�z�	%V!o-f��P��S����ہ��r���up/��V?���m��k/���h<s�O9w����Os�]�'�W�^���N��u:��_JWi}����%���l�Ԯ�˳�)j�7��2s��p���!�{�\�$�V����ɒ��f;��Ѓ�:�ݨ�S&���)�_6)�7p�fJ��+�s2ܠ�a����K7�*�2.X���m���fJ�Pa�#߁.�� ;R���*(�G�]���J�>ɿ4x
�9�Gy[��N�X\p]1�4ά�L
��T�eY�-�8�V
���Uua3+�[L㡼v���]�̉vX`��Ec{]���ko��ӳj7ȵ}w}�@/5�㡹{���yz\���n���k't,�޷�+~��A�8=Sf��)����V�뺜�����D�ٍ^b6���5}p!���=�^2-��+p�ɡ�o�{�t�*�'�sy�xl\�Ǻ�-��_.��u�˻��V����eJ�,	�C���� ܡ�bz�TMC,H� =黰2�<w�	x�f����ǈK|I�I�f����]_r�'9�pH�!�3�Y�7ul���rov*A��9��ގ9d��1S�c�r�ݵ��B7�E���'�ތ���u ,[�Q/>'�!j�d@�������I�x�CifL��|Ι���i��,�*��k�嶍�����O]n���\�a��iV�١M��R�ƕ����ϔ���
-���Rժ��6�����ݷ����y[ǧ��H B����o�)�_F1�&�7Y��s��톡��цܽm�h<Ö�f�TޣbL��v��,ڻ�Ӎ.g1���e��f��&��%u�kpX�@����Ý�b	3`��9�ٺ���Q���32��H3n��1�ү/!�k�C�����*��t�ކ�3J��af��$$�gqr�y�u��I}FS܀�<��[y�oJ�h�e 0�w\��
Eo<TOwp<>�A����e�
(�M'W�gur�)��`R�>��'�w /�����b�\ђ8��J+&k��y:���a�(R�/h�YNˬ�D��Ń(/E��[�m�{2�h��:�pIiZ{�t�rPV�}�A�^��m\�p��
P6�t��;� *-���낎�̖�	�i+�X{�r�v�H��Nk�S۶3�̓v�^�b�|�ʆnT���8����Iv��8�q|;��:��к5�Q�d���ԻO=Qq�Ӷ,��kyUnz6O��fғ��A�I	E���"G�T��w�W%�um���J\��Es��-�<��՞�S}�yw��+rI�
�;��~�[�_�[Y�%J6�0w1�o�r\muZ�-qK�h����EU�:��wB�w��w�	Z�z4���a��͙uHa�z����k���e����5E������]l3�5��*��{q�왴K�'-(�*"�eC��� I8�Ld4,�Ϩ�`  ≯u(Blk��r�r�b�\�F�棖���˦��s�u��WK�g5\�s���r6�u�.�Q��k�[��W�m��S�r�X��c�]wk����y��.�"�us�Ch��ܮ�qˑG(��7)��wv�4RX��\��s���#���*�,r�N�;4�QA���;9I��(��]��9��
�9&��ME��+�ѻ�.��9ʒ�sTu�p�"�&79�7wj�wTk��WwQb6'u���' 	��ߜ�R'u�J���v����u۝��զf �C	�KC��#�Py1Q��C{i�Ib��VsN�t�h:��3���W�P�@��8��*ON9]َ����h�;���>���1��q�W�G���k����߽����?~�>��1�!�\�)vo�G��k��{�k��r��հ�4���$�<!�v~���>���e��`�6(�$��y.;�[%��8����VI�j	�|ط�qL��=;�0:O�M�T�T�gn>̠mU�����**��[��	�,�,R��}1���2������9x(7Sk|�:�E�&����z|t<r�p�,{��^%B��TXS.��|����Z�r2+oD>�^j�{Y�#���3]�xI���WBnmwL.�b%9)H����SmG@�\��W+T��r�pP�Iȶ�C��!ƟC�>���[|�6A�lM*L��٭���t�i�h2�Z�Ǎpf��w�xa;�A�C���zA�	dnnYe����,�l��ߑ�G|�y��/|��3�0mt�D�\�=� �k��9�쥵�[z�ҷ6��^�g�*z�V�u�4��Z�E�����p���D�4�}�b ���~�SW��}M����4ˁaߏ�g��}��]'���{��[G[��}�bmL�k�f��˄رP�����jJu��N���nS�E�l�t�/��}�.��=���h�S�$���m;���ǚ{�o�,����fRX�"������s/��3��.^Ώ�m��@�I�LW9�7B̓q�߉TXP��̦�֑<���]��0�ߴN���N��ȽU�C^����L��?2�'�sN��:��:���{*	{e/�. ��uB�8o�f��꠱��;�8`��39� >'4'e�m�,9�aJ��˦�ѹ`ݠٛ昍i����6w'i����W�@����̙��� �oו,�:�7�ێ���c}6j\]�e�3�s�0^���T�v�2� �c�)��{^]� `L��ݡ>0U4�e&�xװ�y�������&��ȴkL�C���ˢ0~��g�N�>�	�b|����}�I}��ճ��>f���4>��'�N*�Gq�א�yj���J�!A^i�)�WL\:�P���2�e]�_v,gC[y����{Q�]c*���(_���fP�c�Q�	��Xu��*��/v'r�h�~wB�l�C�1L�:ll�3�~v�-�d�NԷ79�����έ�
JB�8kvݳ{:z��u+�����|���흠 b�0�2`$$_W�i�y�����'�T���S�w�<<Y��26֬��䮎v��KC���I9�����d�x683-�K��=�U:�Y��g,V���),b:vW�κ��| U<�e�gW�uG/VId5}ݧ\㍌��'[�樆��s/�L��Ձ5]��د2B#���q䇥tE8)l,�q���Њ�v#g1�k�<'��|���2A���"�|�Qx��]���Z_�A%�^�wL��Ĳ.�7E1�
4�P~���5��}*/��G�t3h���3ds3va��qJ{��t'a��٤�>��0�U(��7E1���ۋ�r��k��e�]\�A�<r-�Mo`P�-ً(B9�OH,kУxi;�����='�%�sT�~j�Y��fX��j3b��p��-ê�d0�t ��kJ�O1��u)�k&�Wr��K#��.�5!?�F4?av\�'ŏ�Ԑ�Ne;�
p�7 8�ç�:<���X���j��-l�BU�-ɱ �^��A�j�s_*g�g_��t<�$�/}q�&�Y��-��
a?���4uxǍ�SD����9P5du"����kX�FLm�v��s��u��siܯS�����Lg4pt��-r�N���X��n�E��ۖO�7�;t�}$�_�x�0��4��zA�Ũv���µ��%Ū��v��z�vi��E^���KsgCa�$={�@"I5%�[�|ޕ���;��K����{u�[:���[��g
����Q���,JL�dm��Pǈ�x����yKP~z�w��)d�cb�OJTtX��F��'���<�Dr��[+@�wL۷,a�3/�1\�|Rr��X�9��N�s��=�Ҿ��gv2�_���L��p|a���?���I�OFk���͛�Y�{$�4YA�m��[BJ͑S{5ݜ�E�^j�p�_-.�7��?�?��Z���J��*�{&��;��u�K����x�s����'CrΜ`Z�#��l�|i���"�x��a��O�b�}U�}��;8����7=N^"�uy�%6߉�5Ji=���Fcׅ�[�z�� �d��ajK{�(뉋b�̖��D�u�����Y=\��'�%�{IM2�F�]�Du�5{gO>��rboQ���f��4Mv�#�D�f4%ק�"�K�'S�E'7�R)�������ܞnr:�:��B\���g�[��[/�#�C5���6����-T�"l�w��$�b)9Xt�=9�vE��Fj�~~]ܱ�����v���0�a>�H�!6��l�{<�_
�n�	���.�[��,+���ݨz�;VS֠�B/CQiH�������@G�J>��q�_r���(��,�~�ʦz��˜�[�}&8�!�#X�_|���$:~��ZG�(��!�!{�n��ߣ�6�\W]��/���gn��"
F7\�w�:�k�6��wo9��Gbˣl���$uԬ�vsرם"���L��u>�g-8�C�L��t�J����S/�RH��E�4=F�.����H���t�� <Ҩ`X�|�ާӴ�ʔ���;¨ (��U�;F�v��W��Smt���0���ɷ�\���P����'uk�q��'��3ƨ=d"F�eI����z��z����dR��S���r��q��m/���ݒ�g=T��i��L��;D�L�[S螇O�3��i'1�F����:��=n��^�����ì��z��?Z�����px?��?0�́;#Y+��s�ÝBk��g�nL��O"�Ob$���N����q+C�T9KO�6���`�o��7��?z�⵻pwO���ɷ��݃J&��&2!�wf�f�N�8�7#��ԟ�疟����bO���n��Me�cY۴Ϛ̻������v�A��A�pI��CPHγ�͜eY���=;Ճr&���	MR���ټ��E���v��E0^ۭ��6���L ����	�d	b�N3����N���V���s�^��v��7����`t�.29���:ɨ�\��A�?'��ё%J��d��{�DFe�ZRbvqc\�C����.a��^v�^�7	��ū�$�D�=��:��}���O�t��Uo��e���Ư�C�2��0����l���s�^J�y�JS6�;�>���t��W�9��&����"��r{4w>�m���������b��'1�9�y&���H^��J�y=7�����a�ӥI�΋Tr�&P����o��.�3�����������6g8��ƃ@t�zA�~�D8�2��bo�����]'3+�������'��P�_@+��(��2�v��k���:.f{}��mV@�7���ZD�Gv��vT���)�t�ع�n��������l���ҷ�+["�]��{�U��W:�I��=t)^M�UfW<5xZ�E��RX�-�a>M"_���,�o���ū�r;>��4 ���ܞ��W9�&�Y��N8�%QaB�O1�WZ�|^�>�l��V3e�t٤zF�^��,2:e,�i&1�9�Fq�jéX�?JװT��V1�^�R�������
�/FX�j�a/�(p�^��|�Sb?m���R�c��	�9|�SFԜƫ��ʵ��v��
�nj��^��g2dK���D&#m�&�uq,y�\���Z�i���P2�
�&7�a�÷c�̻H:"��������ľAއ�V����.�+ovTY�v���[�����f���<�l�CׁPi���>:"�WD�����������{��uY�j$j�g��Y ݗ�Q$�z�	���2�,*�kmvo!����Tᵙ�7�鮤�]�H��e�o>�7Og^PR�ޙh�Ӹ�4�������:�� v�p�p̬7�(K7$��k�0
�H���|5]m��w20n���W������T�#���Nrm�o�{�%���J�!�My��)�Qe1S �n��h[3���9B��Da�q".�ؚ�j�ʩlj��!sߎ��,�E�����cQ�{���yy��áfq��q�^���c��៰G���^��&Է5�BlL҈��g�+T��&)��P����L�5����n����4�Py/�1m!8��S!"��Cŏl�*a�v��7���Q�y��x�����	�T.�g1���Ŷ;�am^*�I��������D�����w�Ĳ.��)��Ɠ��_8��r'�Ϭ�zw�x���ꦧ�g����'~���p8/����NS��P���<���̓y����;_!��6C�r��ޑ�A�ל9h3sO�p��S�5"N�4��W���z�����'H�1W-�0@���7���"�;uKϡ���aP��kH�5����u)�m�r��*���gQ۬\Y�~�U��_�F������q�.���zGB9�a������s�Z�W��7d)��V�4
��/���;U�w�T��nqrs-{_��q z���WϢ�"s���N^d���x|J���|����:h)�*+q�8.��B��E��\�f�KW�:��Qm����WrU�9��\;��K�+�A��X*k���r�u�Z2�l/��S�%On�������PKܽ��9���6�E��tØLx>�D���4{w�Si�x���q�i��'j�^�m��I��Q���=�L�1ۆc�ņv2z���㋴�m������u6��c�Cκ/bL9~���7ҋ����!��Z3��@�:"طPwc��X�gǎj��p'�ڵ��#C�q1=6^����KsgC`�ŗ���wzo7_O\d]M�S��������>�ߥ���L�������6;v�6�����i禐~�3���f?vl�^�1tgb�H�%��9����+��s�P�y�e�������^ff��h��F�GZFm�$\өe��XF��y�F�K���v1wl�n��+d��#���%঑�^v�̑sNdU������.7z���z��E+sAn���d
��Q�$�P�Ʃ��u[�ҦF�Ӽ�Y�׵��{�|���_�^69��*�$���?y����~;�H������d(�Y[[d��+z���͸�?Z׮�r	^ܹmuC�)��(l������Z�kY�![;��\��^52�y���x�=K��n��U��e�������[�WOw%��_z���dU�x��bE[�D�ݮ���N����M��cc�yy��\U��<F������ !p�o��7��|
�e4{L��s��"��ޥT�k��+`�}�?~>�{j�X[���P�َ��4/�lӵ��ݷ;wu��rGo#0�V�2�b�^�fq"�@a�^�r7�F��1�e�{�h]|Df�����Ƿr�_y֙���?�݋��!nc�������2�/�+�Y�Y��ۇ�8�f5Q.jsJ]@Z�~���Lי�gw���j$M��R�!�J��׽�X@�^ptȎn���y�\[U�ݝ&�����ՙ�0��"�^cṅ;�Я6�n��pЍe���l��^�o�늧�c����[g��b*����X��p�Y�éXì�B��S�Y�rh�4t�E�ڐ}Xؤ��D��E9��tG�_C�J��(�lx���,����]�f^N�Gl���D�dH�� R�U�ndl��1-����	촬H�hTP�8zPOS�E'ٖh2ڻ��9s��Fݬ#4K��TՕۤ	��ܻ��[�Э���m3ո�R&��$������轕���+����#��
����U��
R���T/��.������x.�ݛ��	od̵�Ӧ�N�F''ka��N�������|�����*τ��ה�պ����3�ٙiF��:6�e�r�	�*�� �{����W7��tpڋ���4��u�"17�ֈ�#����9�WQ��#c	�5���v[2���t���{e�Y�:iԊ�x��w��Z8Ej�b��ڔKE]��0WKngJ:k��[t�́ ��H[�
�RB�ҳ'l�i�ѱ.wu�b�H�H��d�<�=�k�3��^rT��혍O��f��uΡ�1F����)�j��r��ͲzzCkl2�kV�DK��y�������U�c�����_%Ues�*F(��hr�\�oOb�O"�Q�k�l��i!��0;�q�<�O��s�U��ʽk��*�N�ﳦ��n�w�Ϋ�S�泳(�ËF�Om�iW�+��}Y#����}~�g�����}��g�������W5�=A���l�ͺ�m�N���ԥ�5�����-�8�=���ݮ����xfC�6����)�D��/�e�p������/G+\p!����PsG�]=з{�Y�����$2RN���*�t��\.����'8[n�>4�7�^b�(�L���\kظx|�q�rՌ̓x�`�&%QM��ǀ�yo��?y��=�%lWs[���vF��r�N�}/n��-�z55W@��TM(x �<�Y}���z����:���}~��� �[�/]�
��Y}��ȯ�����2��x�1Nm�|� ���
���~�6��>�g����<�o�W�dͬ*����@s�^\Ϧ�F:H����P�uvs;�r�_���R��}c��R���� =�!�A���}^�Z/˲����b��E�Os�,Y�BEt�̵j�N�f�Nddv7�����a=f���v�}�S�,��}�l��,;�k�j�[[r������C��l��Y[�t+MԮɚ/$ۑ�l6�wZo�(kI6\�	e�ф�p��	�Ր��.yV���D�a�m|�1	�كkOOK���Ra�k�˃w�,�$�;��������VG��>2�����<N�	�iF�|���D=׳�ɜ��q#w����Q��jO�)W/��_���;~���mLǈ�ѥU��ށA!������ݹ�Y�9�x��>n\�ԝZ�k��ëQ
���S�3�왂���hK(*m-�]&�vt�����#�xM;��ݾ����t���E����]EI����Z�U����|2���VG+;ڱ{�g�<�����M��M��u��B�x(h��cwڻ� s49�.����t��PY��~�������Nmc�"�y�����m���N^�nT+yU�Z��?I�GEĆ�WV�<d��b�XfG���RWNʍ��XK-����"�r��y�ؚ��0F2v�#Ѱ>}�dX�I�e��s�9��V�oF�;�h��a{]>���?�Y��g�o��܌k���J
,�)��i+�ǈ��e����V^���ٮ���]�զԩa��iȬ$�ُ8�z�,�q���-�L�1iŴ��A��ޭ�[Ɍ�m!v��h;�a�bfs�r�Է��C׫-�TXL^��J�������T��𚶝��(�nK�^f"��7���CN���]sC�\������T�f����J�(ó�������I��:Y�*��خ7ݽb�S�'���q���3�������L��Zv]Z#��s���ps�E�u�=fT90D�_	4JZX�R��7uh���-[s��{t���6f{�vv���y����}�)�@q�y�襖�W'8m��s��A��~#���mMTmi7�bOV�F���`��0��ː��Ӕwg>O������ⅶ�|G�$��H�J\�;���.�q��ፁyۖ�s�d�n��\�r�W:n]�.U��,]�b����b��S�ܢ7#n`6���n�q�\�F���"��W-s�惜ٜ܊	:d�]��k�u nv`�I��M��9�+�t4�hE�:�A���
s��t�I9�L�]��
a�#wU���Ý�`ܮ�p�:qːRc����t�D㺍��%Q �wm˧v�(s�wUԃDN�%5ݻBX�$�wts����s9�f)$�f$i�U�I��\�;��;�]ݴ@Y��7����bLA˒d&Qwn�JfL# ;�뫥	��*2�;�����(�x�")2�O��~8��]<���1�9������I*����w�z���#�s�Ӑ�y���I�0G�-��������=�g4��O�~��mJ�4`����}��<��y@�3�&�����ݬN�ǅ�(��C�����ۓtKE�toj��6��p-�x��K�����;r�C�<�	�;ͱ}|��4���Г��}C�>O���qm�n!t�����;<�B2�U����"3I"JHH��tJ��N{*��N�t�-�4wM�L��c�Uj�D��X���\G#$`=?����jW�G��	�����M{o����`�a��עnz�b�j .��������&Wd{t$9�HzD�����Mi�����:
��~���FGVC1����~��9��o����<�׭(��B�;�"�ȫg@��FW�!�\�֫f7W,Iz��.	ml����s���%*�US�܍�u>�g:�H�[*rس�f�=W*�!ȹ�`���L��:(fzt��?WHk�@g����pS��w������:wr_�'F�oY�{��2F�mV�z�S��wZ�g�ݸ��l���fX��=��~��Pl3�C�o��V4Z�Y�����ÃU���;Ȏ]�K������m]k*tQ,��GS{6�'ܬ�4W�Tǹy{�Vt�U�M�R=5��n�^���KZhOg�p�iT.�WA+IW_���Uߝ������ ��~fPֱo����S�#!�;>��kɳO;%kȣGSi�٢Ga�y;�?f������'�u[
�����7[����)�Iф�*f���m�3w+��o�H���kt���u����0�3띭9I�&���lQO�I~x�������Q5
w:�7�v�����]�q��'���h���I��bZ����8���z�1��b�J���1��2h7G6�M�\�\��M�ԍ�v2+ <u��m���}���z���Ż/���tY��OT\_n���q��I�g�j<F  </��v�t^Y���:��Vo;�w� |[�yp1���/�2Ǘ�h�,���:���ydDVKԵ��}�8Q��V�3G͂j�V�9�t��؀�P�Mz'�{�>�k]�2�1߷w�Me�(&n�;=�Z��帪��s���5	�+�n4�g�M�/x��5C�rX����6pXG{�xL�`�{��T���v�ʙ4R���R����ٓgS�ץ�U�v�Wl�;�}n��\'�,��8WK����|�}���i[$��e�F�x��$u�fڑsN�l��u��ȿd�{
k�N7t�R��[�Y1�=^�!ux�
i5mQ��e�9ʏ[���K��[�F���h�������/Ǵ��[#]�B)+л<n���K�Wޞ��j���w�׊���8����v%p���&u�#~��0�<�Mk�mj��OE<�u�7����@B��	�GXS|
�e42���QϝD�F�in{���d1���\Ml��]����9Sk��~�=�3�Z2����4n���� ��8��컸>'�@��%�y����F���:� ݷ�b�S^�Y�|}S�/{*���6��%�+��A����7��n���%33վ1����/}CEa4�1�#��{J]V���eT3e��[��T*ڣ��ƹ�zD+��ܪw�W��L�w՜��x�_��0C�}V��۔fS��{@��s,�kD������R5��%�quIa���wp{t�8(���݈Rvՠ�+�w{�׹q[gN<]v��=�I5PmZ�&EC��$��w�����.���؍p�E�H�F^���+V��7woi��&[���$���T�j^�7�L�"�p��e���|,�ź햡'U�����ǍX���7��,8a�a���Y���uf���9�bU���b"�q�r�d�3����-�A%Ή7�Nd�t@�}�$ɾ��)���U�)�v���n�w}y�I�5%�O���Yf�/K0i~����-�3&���<L�nƽ��I�]^�����ؐ�;�pEv4��V���LJ���&Ѻ�����6+``�k�V"m1r��� ɵ&��c9o�'&w''{eF!�c,��~�L��p�W1!n#^�]#�t9J&;��/���۱Oݞ��M�243��Q5�%�H�g�ze&��Q�F\Ewm�˭z�g�?S�f�x�).sƨ>Zܣ�G3�^C�-�H,9Si�m��PݢZR#���N��C��\e�v|�Ng1�`�Ǝ�����x�F�WO��q�L[6k%[7�zOƻ�]�_��������8nQ�|�;GI��sm�ױc�er0Q(
��T�9��Y]G�z,�K���L^q�ަ�YXs$;���7�WSr��{�z!��b>�-����1k��\=�V�.�#:ƌ�ߍd�,n���N��#$^�*��w7)V�\m�,\۠���:�7os/S3�z�˴�i����r�L�5=^�J���T���a�Q�1��p���=J��a�@a�ò�^�U�4l�N�ʅ��g{i�64&Xg>MtB����Ļ@��0p7O����`��U�I��Uy�*�stN[�\���z��x�Vq�c����s8#y�͊��,���$k�x֬.]�{m�Q�]7CT\��>�8h�cp-���Md=�:r߻���-�����ן+J��o�LG`��i�3�޳���'WvUuU,B�ԨF^����bt�$��\��JPJ#A���ÕU����zI��D1G���ں��oh���WǕIU�\���wtw���L�k���6������^���Y(j+���K#�3�2�Y�4U�����츺��K�7�c�"��m�r>g)c��SI��i,���x*����wB���
��G��:����#0�=.�m��������]� �2>%�4ga��;&��ڝ�SK���v�OC�5�5���k_3�2l�t1��Hu�H����h��=HS�@�����"�{g6���M}��펺�rJ���P�.��۹�M9�V���V[(g�=l�`<e����XB�����֯`��m��m2�4�l+��bg4�ԓM�������m�G�x��)+/�[=Ǌ���[k�m漝������=���
/�uOg�B�E4gI*�*E_���H��a��v�\���(0�]�q96@d�)�!�pY!�5u�\�R�ȵ:�g�U���Փ�����ۙHrF@�[�`�6�1����9O���ŝ*y�([���Kvg]�;�4s�@'t��4�������{S;��C!������0�����K�R�KJ&c�?L��2�쁾`G:n�0w7�"��u��:�Iqe>��{�h9[!��ҧ( ���u��{�Уl�����������~���n��%>ξ�(A�-��%��{_>p��;�Cu�]��^\<���雍xſ1lI"Rz�������̼E��yP��]2��q�"�[hm����1|��4���1�I=שl<9�c-ӷW�vQrj����1��|̐�:�h�e�]���0�r;t�k�M��� ��2#��/��)��nc�3NlBŒ�zvg�4v6�@���;?�0��x���:��bG���31,���l�m����Yϫu��,����;Ȯ���~��Q���T3N���Ѻ�ȍ�=�qu�H9�yJz)��%����U#&D�����Q����{J�$w$$u��8�"�	l�Lju��(}�X�%;�n�U��7ôW/�7Ck8�Ll� ���4�����d�sNO�i���-��yzΣ7�`�V��j�[��K��@$�P��1���Z�먖Ȋ��$�x}��6����g�"ݕ��"�d�3��;]�fx���޾���|�Ҧ���>�uә��@"��8)�����ЌH�"ETF�j���;��|ټ@m��:��:ُ�o����x����}��1qw��1s`�"��V���Eՠ� ���'FA�Ԡ��4F̦��g���i�>��g��!��ۆt7z{b؍��?/lѿ)�X��� l}y	,���ܮ�Vҧ��Ӏ��;����R��oS
V%զ��!ܦLpK�̺ԙ�+���:~��=���4�<+~=�6���c��:� -�#��[��t����w��amPi�3i�H��%ez6��ƅP~Z��iK��c�a��tF\0k����X�S���aΙ��B9Q.jsJT�Lw��
H��zA��ih]j�"����`g<���S�5��������e]��s���WPt��Vn��s�i���_�޽`�؏F��ǽ�R3��3K�oQuS{�w;ͻ�W��iO���lt3��|	�gU��-�ɮ/�Y��4c��'��S�e�i,3G}�4O�Y�.%��=Lc���0_!�s��#S�z޷-���Gg3I~�ެ_9+*��Y�2����<�5ծ���?e�qi�u����6(bA��M͋Ųu h�J�!���Vp'�X����Yw�d���X�T��.(j��6z�LZ�GaM�9���P�͙Άw��n:�Y�J9��� %9��%j�x�wx�Ń�Y��/\��r�_���D�T�)u>��!-{#fpW��>Wv�Sn���O�G�`�M���qH+7W<���{�5#6-�X�2�� ��vK�Μ @�h	���x{��zov�D�Hϙ�A���1���Z*5���B��6�[
&e�Y����ԿuEn�>�fO�i暀@�("�А�/��q����P�ӵ�g�k7����W��4IHs�z�7*F废vd����ɨ�;]DUQ�7��E�#th�ޏgA'�"�t� �2�:*\�̭��g��g�zU��S�{E/�'Ѻ:�B��z^�+����K{^�Fɿ�L����.EN��X�	�w��'=f��_%T,��oR�h��8ݳBz����*I:E�u��%P��6yO�,��w�ѲU4f�]Wr�7o9k'I�iNMG^|[�f`� �쎦�Ð�l9�R��T3�RI���s�	F���I��<sr�	�j�썾��|�9���E���Ӻ���7i㷚p��0�k��M֨��^�:�w��Q�8�w��f��z��-c9H*6�}����k7l�2_�8+8���uwq�9�}N|o����ɚ���2�Ya�������&O*(U��fQ(^ݭ9��e:G��4�!�]OENRm�:8P98-!�ھ��rNڥ�@�+a�*0������z�we����H<Z;z��@��	�d�-׀��v
�m�>�>�t�-x6�hf�u]��X9^I���;G�,��$HI! r澛`]��*�b�z~�"���g��zJ}W]��xH�=3���C���6ǜHHV׾m���T��O�.�P��]�����uSJ�����x7���_�5O$xWe.����4�vY
�
�~����ٛ趆���ź����1����4��Ҕ�ۺ�sul�l�lk���gwP�5���2��saV�ǶzU��8��B*�C̡��Y5���)R�|/���O��`W�d���+x�IYxElv�<T�6�Xթu�lݦw���O�%�?uy�R�����h�J�(�hI����C.vn��\�bz�S<�j�D��l)��������rhYM��?���������{=��g����x��5���:)����ddാ�\
�1�����/�B�v5�]DG�8[h�||������H�rl�U��`�4� a冚��ȄX�ȕ[[��z${�l5R���m��e�K��~٩����{���0���:M�|8Ǹ%�դ�β��̲Z��3ζ�qgx̓�H��.=��j��%ջ3W{�om��;�@�oL���9��u���?��v&��qm#O,պm�f�<�u���:p��Ч��Ǭ���{���kN�f���B����l64���U՞�!u�o��c`5�n���?���eI_˩1ڏ�{�>ܗW�uȟ.�ۆ �N��{�׸?` ����u�k{DXՑ]� �y[N�#�g^7ԟi]p�6枷�h8�9{}���d�x��/$����vΆt�^�v�ҲN\�}s�؏1��rI��6�N��8p+u�}1�]�ʶu/M��j�P���f�R���/	�߰�ݖ��!è�n�w��Ħ<�r��;�C��_b���Lp[�#ޗ}���%2�c�[ E��a4r�GH�-^�4/�T\P�v����㙲�Da���z8��\��"E�{,e܌]cַx[̆��pa�<w1W�$�tO���L3��׉�{!Q�/�	�����G;�2��3�{�{ս�j�ǚ�Y�7s��X�s�`��4}3��j�n�[�c�Q�rU7o�mB[��w	T郸����<��L�Q��3[��7"�搔�<׆�m�����<���ɣo��I���7]0��C��;q�8Z;'h۽p�C�8%�o��J`����h�Sz<���Rgt�H5BTs�5��jǯ4�M��;� �y�rVj���ױ&�L�;�{�BT �;l[������r����g�Ou���c_{�%�p�Knni$y�E9�ʱ�zU-M��=�L�h���[=��4�\������3�v�^|�q�u�%eck���y.;�U�L���w5����*��ᄓV�`ٖϧ������g^:�Vi��̸9��gO=��p%qT�#X*�����Y�o&�!E<����=~/���5꫙�o�M:��}6�u׆CK�`�c����������&#��K;;��W�
�G�^�ɻz�8q6�VX��V�̊}��C��8d1PS�u)�F9�i֪'���N�v�#F��>��4��e�A}��C��\���Qe�7����޼<��5^M�-S��\��L�<�����}B���=o�����a<��L�,��B�׌G&���|�Ml�ܹ��ʙ��r�ycvl3K�/#{�.������D1�$��W��2��Ws/%��GAc��DW��sgpս��>�#��@�/�O׀{�`;T���;(d�#���,�_��'����'n�!t*ƫ��u;����9����`��&�m�A5I2Sv�BO��%F'�p�R��I�˩��4"R?N�x�J�Y�;�Ȳ&��9̑���&!H��9r��4Y4���j#]�XL0a��ܔ��d� ��(��b��#$h%�v��!�$҈�D\�Bd�
 P��d�ѣB$F�ӬI4"d�)0����02LF4�͛�ш�L� �h0Q��4LJ�qJ2Rs�!`�sqPL�DȂ&$�E($L!���5H�fL��Y�DJ��dD�HH!��	�H$sp�����I��fc�	3)����4��e�����������|���7�E��(�5y��.�puP�n:��B�����ƖB�mI@l�,n��L��]r��,�'cmn�a �ޜ�l������j�����J2���l/������R�x�y�dmY�d�Aa����%�K9��&�O�0}�_��7�I��1O;��^�W�+^�]��;5����~�Ty-���S���I�|7ݙ�i�6f+ȳu��/���m�b��ܑ{Ԩ9[-�n��9D�H;b��L޴� ��S���ճ�Ȥ�8c8#�>ٿF2��Y}�G���I�qn��gz��r�k��U�^Ft���fA���w@�K:�~�ĳ[t�3;�����W˂��3�½=�v1�Ï�����a7^�gC=���UyF��:v��n�N�\�3y	Z�e]-yp���~蠂S8ɵړ4��m��3�Ņ�U�kݝ:M����q�R8ۛjn�F�f[��䵭�r�tE
����»&�;Cx�����R��v��>�7%�"y�S?]�
ڽ�:ySe�˼R�c~+�<�紺��d�uwH�u���]��(���F�z⼫�zN�"��~�����/��7(����)d|\1�P��Gs:D^��`�.w��yu�A��>��[�r8�a��a�u֟<[���\�tk�u�ַ�,6��
���#˵M����P�(�JR��׌b1�C�m@�'z�g�g����ԁV� 	ȩ�EW�G�Fu�4��Q6��ݘpg�vI�\�R�]�u#L.�� >pS���96�Q ����=m�b_�u������=>���<N�^p� 9	���ޞ����޿5=M�.\))\�r��mkgd ;��޶i�����p��T��9}��tN��
��ިꞾQ��^M�f�]ڱ��������*&��Ѿv�'�<����b3���l��F��JT�L]���Tz'��[�~oU��
��n����G8�u�i�^}�ɵ^�ɃٍSM5+�g#n������(8d����Ӿ`���G �gZ����w�}i���n��8Ξ k䤛�A1�h��y�G6��W_�Ҭ��Qwq����ɻ�0�F��Hl��q�Jd�N�4n��y�~�F3'�n�`�9���zVAa�V�O{�-���u�CG��g��'�]/Ն@���o���Cyc'No�mNή=��2�%Y.ƫ�h�Ʋ�t��u�H�{\�-{��Ge5����ʳP$tf�OG	�m3�%��E�c!��j{h\ok]m���x��7�1u�I"�h�Z��n^X����͠u���a7��
r( =ި������xrN�x�J�
�V��Ԛ��:�f���q�5���ng���9�_�������ɋ�=���^9wwfV{X�	f�S�	;�?��X	=q�4潥�6�9��� Yh���s�M�z�5��g�s<��'O�oM&����ٓ�O4�=PE�C�a�}�Q*fȞ�)��^H�E+�I)sƨ>Z�T*�
��QyaYiԲ�e�ܜ�	F!�/A��t"o�"��3�?���tT�R�7:�u�f�p�Ǳ��c#���ä_)VSh�)P�+��mkd�U<���Ǫ������ӻ>��_B8�;r3f����W<�G�����߇�X��l;��ln��tM�|8��c��Zw땝@�5M[�w�g@wb I�"����G��i���չ��5�nw}ǭʓ"�a�����<��d�Y\MXݑN&���b�޿�œ��*.�N�r=���Y��G��3��L���2n�i� ء�9����5�m[���*�3���8`|!L4�R��V-���ɿ�y��*�d��u0}��|Wdgj���Q7.D�˒��爀;o8�ܹ�r��RS�v���n��
9ñ��|HO:��Tf��Wb���7>�)�haH�e�t5E�o3�3zy��ЖR�^j�v��������Z���x��P�mVH��x�_?�8�d�b�t���f�L3��۱��퇱�cڨg�pE�x=�7��Ԭin���� $�����kT3�U�Gn��q�{��c6*1��m ��BZR�W]{��$Fu+��95	�|��m~כ}�X;�5\�y|v���)����e���d���}�Y����f|����8�i���4�vY��?�#�^�m���s[T���Cww�2#8�t4��ZR��Yګ��5m�4��Os���Y��+�y��xc%.�sG.|��.\����ːG�; ��c��5�ة=%Ǒf�2� ���g�=n�zݲOjP�}#�^֪��bQ=�wt��'n;XQ61Ǔp�3FI���{kpar��΍�D9���S.����f���Ύ@F�����'ؤ��=]�M��d
�+���q��۽~�h�2ww
hF�Y�{�)���p +�.#&��G����)-gEdl5����x�Q-y�٤�T�u�n�^k�3�gTy�[��p�&ѝ$�[�J�h�:Su�p�̜,gf�0ݞ�����
tp�>j��&��=1��VxX&]̎�bj��z��/�#QnF�[a��a�ky5�õav�W9OhuGgU�䬽�J1>���	ݐmO����l�s�h��]ݚ�:f�fn6��Gh��q�O�gz��K�Q��m�����d\���8����$(��;��7���P��Ly��ۗ�'\���7��߼���5�
������}�q��2��?�	�c϶d�Y>�/���z�����w�f��B��e�d���x�-������ w@��<+4#q*�@>6�4��|X��%Tz�x�����s���^�X��O���D��C��g���;�}��5{<7u>
5����c��k�8�k<yۗw(A��apN�����P�z�n[��rUr�v�C̴�QN�j�� ���͗'u���d��LC)�Gm�)��&�<���P�o	)� {�`�>�������W�ݱ���w�" �����;�舿v�)R9�WK^\��g����$�^@�H�?=�6�!�μ(9����	�C���A#��K.�"�ON�6�$t���7����� �����*�g.1�;[\�R)GH'm�[��nЎ��z��v2��?H�ÇTz�+�\ .�7g]�B!�`%<��F�kӳ��<��Ֆ��n�S��pt'"��U��z�ǗyX5U�NV��ez7�MYǊ��4*�Ϸt�M�"�:B8-��{��Q��e���g5����R�uƼ�=�Ww��0d�x�o�{��!S�RΖ��+��9"t��2E��-�%5ʗ+e�-kd�ʑ���f���vَ�M�OC��8!�t�y�pԽ�&�ԛ�+���H�x��X�?�<Y9�7���zgӭ�j�bd����*��W����J�t$���v
���۰�Ə\v��,6=r�̡S�ve����k)Y8�� >=���m]��<�u|�ű�,�ֱ��%�\sLk2+��+or�D�81�TlL�(M[����Z;N���k���g��y��,�Be��>U��:����ƍx����)���/Zb՗����w&:w�9!�B���h̀F�8HȎ��J���*�c�������tE�p���t�������!���#E��]�z�<k-b��*f�T���c=��xx���ɻI~ög�A�t3��|
��c\���ػ�݋P465��������2G	�m3ļx�=Lc!���8�&򪵺���uT
P���v��VM��DN�D�F�k��O�.k�a�[�3�j�fp�4�l0ё��5WW�4�@�J�:Җ8���y��m��"rw9���a=��U=B&�W�b�.KA�˝�Gº�ru��wP�ֻ�������p���=b~喋=73Wl꒰1����桴Gs�^��^���̑�Oi���ȳ����� �\�v�MMdS�FG��K2�7�>�~��}SL�e:�
�-ZiWNv��k;.[,-ґ�y%PH�eF;1��Go�7�+�-[�(���K����m���S���.�UW;�c����$�"�.����n^�l1wigc~��W���A}��;8m7T�Y�"�vu�J��4J}�<j�-H��\*�>I'S%=��Po�����l����q|�
�Љ�H���2
�-���A>u\��՚яS]��vXm�t���C��GH�2�)��Z�q�ڈ��z��:�7fڍ&��p�������0���t��f�OP�J���n=L�cgw/[j���j�4weUoiy��C������yk����~�ą�k�䩽~	h���U�=ʭw�[�n�����#{�>`W,r�{q��g�v5썘;�
�U��*�ڲ��W�\vF�St��i�b43�k�)n��v���X�!Ř|l��G��B��>��6ta�3���q����Rn2{��M`�}C$r�l��Ɖ�$qn� �>k���ݍS�&�<;)��d�}�dN;��Z�y����^Y�$��������)����kU�l��3T8�U��O8Yvg���N���T���h�h�y��8H�R0zO�xx�}\0���)Y�P�|�44���^��쒌1]	�:��XΙ�uf�a�`竂t{��prH�&/4;I�-漑�Fi�ٲgj��ㆯ��Z�rx;��nhD.߬|+���V��|΁��Z��k��N��΍v��l�d�-骫���n��}xx���O�-OE<���^A(��ɽ�-�2BWUu����s`���)o
:�YW�v4�Z�)zl(|(F�Χ����h�nZ��	E	�MFD{9e#�L�\���SC��\�v��V|O{	]�����?�G�ڧr��D����t���%�OP��ѵ�����,R^rr�["X�W �2@�Jk���3�RV^���٦��&�`���~���(A�1�Ƅ�|G������N�Sd*)���e�E�����g�����ҀA�A�kv}�í��[}S�v�c5w{�w�ݎ%݆�SX�	uw�U��]y�q���ƽ�'	n&���a}�-c%�F��l�4WEΚn�C��FR5��}ܺ&�'�wd��������۰��&f�)7Q|��ʩU[J�G����دP|��miȨ
�˻͋ !p�n��F
^�E���J�z��N�
x���o��9���;,���ݩ��硃��������� j�Aʹ]ܳ��{)X�������om�����:�zl3�~����Qқ�N�� Q5?�Ȼɺ�9� vt�iΊ�n��O���8@�1��"��1[���{���Y����Y���9���b�r� t�1ܚ8�`�3�2��������ٟ�iVM�g�/��Wkn�1�����hwF`<+5��I�۞~�9���f��}���8�v�}�H�,`�;Q�2�����C:����&:���5.m]��3j�o{�-��M%hH�Z*�Hا9y���|7m�',�F&��b��W��^���:���h�q�fڲ���F�C�Zf���7��s?T��n"e�`W�l=ܪ
�*ɍ�o��$�Q���&�=�w�|pU�w1�~��͚HY̟\ә���QB:�]�E���Ӕl����KP�Uw��
��wv��y�F�z��
�xӑS���dt\�fի��gV�۷n�ջ�V���Čg����=�����]��B�fۜd���]�ф+1[Y&_QE>�:���#7ԏR�ʻ�d�n�>���Z�+����c)eM���/n��[���U�a�S��o�iS���F�+u�8u,�ݑY �ؾZ���r[��hF�vT}�WƝ��F�����<�U����+������`K�>3hsșܗ4q���?h���m��r���զ#Z���}1i�4u͛9a�p/K���^�,��b��/���I�\vw�L�:=t�dK�����kY&^N���z�u\��s�ԩnȆ�%d缹��쾼hؗe�Y]���Sr �:<����1@Q�z�(�j�>���f�;�c�}\[ZJ`ڨ����p�]X�I�WbrZ�]�����m2je�;��r��B�6��fx��f*�=�{��b�x�y|�4���t�����+��<��iO۬Y�{�An=���{�op�ʅh�7����z�w}�;���W���������|'�i����'y����`�x���ׯ����Ֆ�2�H{-�]�c����A:��=j���M�#�i&QK�e�n�%���`��k.詘0�v.�:E�%&����}P�)��k�>הJoZ号��]j`Y�f#p����t=��u���ve=�sP_p��s�כTخ�M� �r�o��cju�v�>��[3k$r:M��C�`����3��k�C&���C]��Ұ%��TH�7O�Yp���P����� �5*[E���ͦ��),�����m@�8>�Z����
�μ��w�{�4��3�������~�x@;sS�K�~}��{["��0�w�s� �Z,p�Mg^s�[�¶Rm�E��t�t�h�K�V>��wٝ���AyG����}�;�������wދ�b����H۩|�����rS�V�Y�	L���۽F�GJ�Ӏ��*MwX���zzvzX�^2����f����Y����V�û}���F�|2�N��_�_\,M ��q&��Һ����kܘ��ǸE�4.
XWW*�� k;�:s�o��.�%v{y��<���l� ġ�r��D6YЕ�wG9N!1��'>�D4�s�N+.���fpn-���WS���YoU���s��ccmO=�!�$"�#,vʷ���q��R���ɓ��^�)N����;e�k����Gb)Y:&����kϘ��t(�k��0O�.>j۾�7��Q�g�zA��^�=���6OR��儑�f�^����K*�tY{�jSP*Źci����1�Y��S�����Ʉ��$�-�Ǆo;�����n�X��DRY��O^q�|���$�m�~:tz��vZ[ՖM�L��ȷ�1�t{�tVf��U�5��3�yu<;F��mM G;u�'�`��5H��W��������?]s���0D���]�L����@M��]܃��\�L0��6f�A2��!bb! ���,��J��F"-&�$J4�RB(4��;��,)i&�#2H�d�L	�$�ȌH��w\��F��JF�Q��i4DD2I�H%4d�
f1���A*L�XE0��i��4BI�IX\�DwWIK�1�b6H� �9�(H�&��2fJd�H��LD%1@�D2҉�,i���Fe�b�DXfLY$�XLlDbM0K��@'����e'��+�:��讑/�e8�B<��<ts<{uӔ�� 3��~p2�ߧ��=�7�R��ҷU��r�L���l��	� �9����I,zo��F�H��ہ�N��K�\H��n�rb���8�����a%̷�F��WG=��^$]*���D3�c���B��v��s��4{{$�\�r�[��{e���ⲝ)���[ݵy��`<�5>���=W�k����Fk�����~͂�v�Z��j�����8�^�Zl��l��xϣgUG���iKj�]���ښ�/Kw�f`���>�`��`Fl&�y�E����R7���>�>N`��Ov�%�m%�Td�7�7_�;!t�b$�u&��⧆קD�;�8sN��=@���ݛ�c���Pc�ӣ��w9�B��ۙ�$��6(�{=����n�g�G	ͧ��s��K�)���s�7��8z�1��� ��}�Gt�"t�$$D:��놎8��z�;�5�2��c�3�~<EޥVY�2w&�hZya�Q5l'U�$�F|��w�Jsi'3og6�v�9׮���m�j��S&�y� ᡨ�n�t
aJ�m�Iz��u��J�2'�� �
�t�-�vbƭ��K;k���T�/d[��k�`֤>gʽWT/Ͼ߾��V��S���ُ�W#3rgU��j���PJ�OP���3s�Y�G��f�֔�~�}�������mI��i=pD��,�qby�p�5�v�n�c�V·�o�r�v�dߗ��9
�#'�����ْ:i�i�=5a�^̛��kw�;�+�du��-�������V^I.��&*�-HܷX��uf���V�e�%c��.Do7���~΄�@�:lg��0����Ctf�4\�v��܌�Ưлp�6����#�`�4�f&�2��\L��T��y�+���nyR�,�������+x.�G#>�S���u��ƨ��~4�/i�t��N|z���ve�(`����6�썒�q����������2x�h;�ۗR}�yPY�eN�����0q�������S���>���X�>G4g�S@����%�Ƿ+���oAi�х��;�v���/^�t7ݔ�C�G��9;c�-қ���h9$W��e��Z��:�`);wK[�c9LAf��,���ዉJV�c��F�No}.vy��&����sm�f�љ�z9#X�*t�Wj���K��{O��T�V�v���XuJ$XF�g^�H����=���U�#@2���pw=�������j�I�q������Ϥtn�k�������/��!)�l�V�$���3��]]�{���A�����:�zpWr���b�
��b9��/,ƚ�f|����x�#���3f�Z$q��8+Z�9�/(5���6����2��sJhƍ�ݵ�r�{}�|r�D֯�!��i��=��4;� ��o3m�x�W�c&�Wْ�T�=�Y=��XPR��]m���\ә�f�[�%w�wuo�⎇"�TN`pw
��*�'ɕU����Q�'��<����Te5����y������9�!_fzN�$(��_8S�΂�P����m�)ߢ�gjF^g�fx���c`M3�
�#2*�D��R[����촄�}���徭^ⳝACw_7���?(?z��};��h��wg�5��>4���U� �^�CӚ{�3^T��3���cVM�M+9}&�g���ÌV�ok\*�ʗצ�9n��C�:�0���z\�Fn����J
f���N-�ۮ�:�}P#U+�Tm�X������Z���_��T 譩�
l�{���"�WFB�Cl���>=7ˌ���,������S��,�2m�M#�]G/�0�ь�e{��_���Ǩ괉�I�Q��a��gNf�Mr[3m�:��'P}�f�m_�X�[U��R�y��6�@4�q���tțH�F�w�؊~*���"6u�M�$�)i[�jTܐ���d�VE��f$��{��dU'��#��<b/�����LV�v��_Mqnjna�N.z�n��99�ܢ���+lGHm��p4/�!&<�e�`�/�z"L���VL;?l������Ou�n��&:N�3�A���u`F<���ܡ��*%�\n��[��^���I�G8{�`�;� d?��>Mh��n3��P)�"/u�c�`�!ծ���]�RDwoIZ�`��;�<�E�1K�c��x����̊=y����C|�޽d����Sݾ���̀��l���o{t�p+R\�-=킴R������굎H��غ�0��8h��FV]l޻\�[,��2���zV�m��+�`82	��=��Sn���h9|�09w=��-��qc�Μ?OP��<��:���h�GY��z�5K��N�b��7@�g���V�M{ʱ*&6F�	���W߹Y׋��HM��^}��%��G��@#�`�]���Vi�&%��8*����f�R�P�d�ުu�m �r)���;]�\��3׸6��:�9y���ץ ���SϷ��i�[ ���u�왫Ղ��㲨�.�#��-�)+�\h6��8��ّ�َg:�z�	l��,�=݁�
�2�:�]��St�Cv8IQR��zֶf�����=^~�\�-�~�I]!>F���n���]^���S"�k�6��36�'jW{��L�AΛ����q�� ��`y�6uW��0n�Q�O�P�3�{3�;zO�n��J<��N��3`��Fc�+��=/����;��]��m/OE�fF����+�o��y�P6{�μa�Y�"��Ut끎���A"k{�E[���'�Ȟ}0_]ܓ��+A����R8;V%�ۭ�.�9�p(Gp/��C��KYS|pn(:�7�Q������2��I ��Oç�����.�4��{ǰt�����7�]s�<D]�3��~��Z�ۭ]����["�=@�Uɻd��;fGPc�%�����ڰ��;3�]x��p��h\�J��t6d�zxV�Q�įD���<FZ�S������j�b4(�-C�2�V���7�D��� $D�q�#���Sq��3x^]g[+o��:m�E�D+��v����9�RS[v�Ų��(�&�Qu�{�U��j��n��s���S�g���}F���	ƞ&�.�'���]��A�jJ]�������W��0�1�c��ܙ�4���FwO9
�rF}DɯA�TfOM<��竇2������F4tZ^�C�Fh�ZDV���RV�4]���s���Sa���s�k���[��z��x��kH9~"�HY|�\c:69�(t��%����W#v��[d{��I_*�#��I~>���{;B�ї���3�XE�ݣ +r�|�^�Ο��U�\2����zÚ+�<�a���c�HQ�Z5�ZJ3�7Ó�ݮ����Z�n�[sroL�:�fv�SN컓�SwL���i��"M�WF���o�tL<�L
�Ow�H��Qr�Di|ah��<(�Me��d^#ۭO�÷*prՇ�gǧ�0�Ly�_��Fl��hט]��M�.���l2�s9Z�;�"�#@���̤��<�|��ok.鹙�fi��.��ڎޫ�#k'3\v\q�w�*�7[����q�����N��nZ���A�0�f1oPƓ%X�VW�V<�=�%����SpN�C}���ng��G��`J�w@{n����
F�e�k���5wFGa��v���6kN����W��a��&q�}^!)��Z��&H����N�F�ū����g��؁�+gU���p�}c�
�z2������vlpr�A�kͥ:;z`��+n\�pT�/���p��,�zH�c6�~�~�K��"�Y��g���O�h�y5�Z��}phwg��;M���`�_߿��_v����<!���^ک�e�9�Z���hʌ����/�C���YrN��۵��a�eW-���;�=�7�aȑ�F��bPH�6K��<7��ݦ���"��R�܃ݙ�zu�P�S����r �OI'�m`|i���1ο���Ϗ}͢�����鬋�)ox��@,�>[�ה�%�f��%�9��'��oNSP�0wG�A�Tdg���ZR�uN;�����*n/tC��Y��:��qîI�Hg��o_.�΂���Q�	H�I���8֞+�=�O!�߳��?>�϶��5@�(���t��[��+�l���e��p���Y��g��z������Z���*@tVН��^s2ճ��Z3���[�����M�@ݞ+���n�"���WO��ǃ
p����zWF�>⪓�'H�Kk:�YM��אz��	>ԛ�x��NRp팢'����I�8/�a��5���B6��g��K9���k��'X3����yO�^�3,�	�*�>��W+eK�J��1-Oru��
疌칈ѻ�E܊�ԝH�p�8یt_ѭ�"��Pr�z@x�j���v��o'}PH����@��ee�Op�=܆��{|
??5�p\�4����o+6��v5\�\��.1�E�4���?]g^<�� |�%�要�M=�t�	H���m����'-��4rEk���ۜ���+����mH�ê�3��Vq� ܴ��l���GT�O��#�!��8���#}�"1�oj�;���0z7;���{�_�>4����Lq�G=�������LR��"uDn�;�mUo}�F�ؾ�$qc �<�Fv)�FC&=-ofi
CWmf��ɢӦ�66���B:ΰ����tDH��i+C�i�]�Ә�ˬ��t��^֍s1�:%����:�2"��N�P����!ևoDw6���,5�k�eVj:�/7)�e싦���(+��a�1~U�d>���Z���I�����8��z�'�ѝ�KA�ˉst@#��]���Cܖ�9�8_@��%�r�%�#a+�BL��s��Hl�
b*҃��7�յ7Npi��c]H��4_:��qRx$U6���\D���=U��ܥG3�Sw5�h���~|��)��i����q�g��uuy�e{��Z���U�|:��b�|��v��ix77�YD����i;�U�[�r�J���=.�Ф5���W��u�ã�� �i(;na��#���(����N�E=R��z��z<��]��'�����Km
ͩjE;reI���t�n�j��r;�ʟ�����9Qt�5ɣ�%49R�~e��������z�=�K�wm4Y*F���8�1:'o��q��{t��w��X���t+����ռ�p��V��,�v��׆����z�	����趸�/"��^��'zE�(
�f�
�`����9���Ƕ��y��v?T���D��|����wU=#X�n����1ȵ�+^�m��۫D:�j9�o�ﬣ�_�p)��	GH;f|:�:ꔽs�Eᐐ/'w�c?�s��k�\���o7E���:��y�=���g����-'^DN���]��Q�0�x[/�h�n��"1�ަOw�X���$�a���G؅{w<VZ��n�C!
-v����^>�Xo��)�}�}�c�}c��	L�i=/���gLɡ��%Z�]�=���RG�  �/P(���}/���"���}u��Y_M�y�5Uu�ٛlʩ��+fV̭�[3[2�,�̭�[3[2�f�f�eTͬ��f�3[2�elͬ�TͶf�f�el�[2�3[3m�[2�f�f�f�el�m�[3m���[2�f�f�elͬ�m���[2�eT�ٚٛl�ٛl�[2�3[2�f�f�eTͶf�eT�[3k2�mvZ�ՙ�2�etֻ-fj�*���ՙ�3[3VeY��-fU�j̵��2�f�ʳ6�5fm[��h��%Ua� `+ Ͷ�3j�ej���S-j�j�LڵM��ڦm�S6�S5�S6ک��S-UL�UWe��3m���Ͷ�2�Tͪ���lͪ��m�f����l�US6�lܮ��f���m�e��2���m�f�m���fm�ٖ�����[m�*����f[m�6�lʪ�m�ٛV����f�ul�י��U2�el�lʩ�ٛY�mݼo5�+fV̭����̭��̭�[77V����fV̭���[3k2�eU�w��*�~����o�mm��kj�[L����z���s����}�>���o���~U8n���5#�;�R�~�i���y�UQ^��<~�������*���@!����aОh_�}C{�Z��+��������@�-�K�s������C�$DpaT@��m�5�m��6�l�����d�U4�m�Ҫ���m����Z����[m�mJ�����f�����U*[m�6�l�[U����kmk|q� �Ogw�*���
"�  ��	���ǳxD�~!@t��~� ���As�Z}��ȮD�T? ���;@�e�MR�'z��+�9���>ix x*���q `���!EA���3�@  �P 	<=) �Q}��2P�@З���̬:�	�@(�����>��UQ^!t��m�<é���΁��6O�h{�  V���<|�UQ]�m`��РD'E��T���e=R�?��4��0��UUTV�h�!��Ή$�/0�]tuL��"���&��APEe����~BHsO�b��L��65�`<�� � ���fO� Ąw�}�J�@UK��UD��J�	D�UJ�A ��B!U���R�E UT�J���)@�ERIU)
��ERl4 �$UI��ڊ�9�
���R�RD���-�����Q(��!*��
��PZʔ*�hJU�T-���!RU�B�����R �E)U}�����H*��T�S��(J��)TP�$�
H�JI
QUQJ
��Ah�R� �<   Їޝt�g:L�vշM]�K :�tը��f�Uݻ�tӻ١jN��V��n핬�S�Y���t� &�Mm�udV��u��krH���I H�!A�  3=z(P���n����zDP�v-��ދ��
�C��aBx�q�j�cݹ׶���]�P;��렭��ݣ�]��픩�n���ڔ��1n�Un��N
��uUR�D%*R�"[W�  	��B�mR�چ��Rښw��v��:]uv����2۷���5�G�۶uήݧr���۩Mvчv�tηA��cZ�Www]����u]��4�r�DJ"%%T���*�  �����ZX]�9N���]�nuR��n�"��m�f�[������P�uå����wu���*ڡ�m�
 �%R��!
B���E� ;UE
�ae(�Q0m����` W���J�,�
%EY�Q@�-5����4X��Mwt���R�*�
���� ��Kf6��R��*j�@�T�i�4�Ŵ�cC U�5(�  ֡E���P�**IBD"�p  ��"Ѣ45Z�cz�t�m]:�*p� %Le5�C1ZԪ�Lt+���5,  *�%�T�h�Q	 �)Ex  �h L�S��԰� tֻV� �� K� ����  ��� (]�p�4vꃡӡܥDm���)J�(��^   {s�  A�B����ڻX t �, t��Fu��:�tt��Q�� � 
в�F�.�U"�(�J�)K�   ���nU�6�  ��Z n��]�t�vl��v U�5�C��Yֻ� \�   �{MR�(� 4dOh�JJ�1 ���)F�4 &�JUO�   � �� $�JI��U$  19urvwg�����n|�b�nb�ڇ�m}yv�&�z%Q�ǖP��<=���{.�uw���m�m�������m��m��kmZ�5�����/��Ϟ��z���K�`��e 3�p��ͺlZ+. n��]ZC(��;@-`� 5eME�z���f]�x�N�i$ۈӻ���mIW&Kzj�V��a��0�؃m��@���u�ާ<��+-O�b��Q3t%4G�%8r=��5�ũ�)xE��n�<`$暘&ݫ4M�^5fl���{�Uh�-�{ yg\g۹k)��Jˤ�K��L�` ��V����:��Ç�������rU�t�I�>�	ږ�댵��w$�n�V���ĶjQ�����A��I�����9u�Q���=�F�8�m�{\-H�^�룷{�:���V���m�/5�-�'��`Z3�StnM�67+1�J��"��'/f����݂�r)����-��J��V�L�)��j*��;���@��w�3F��*qң{��ܶ�̲@�kl���w�jݧ䂄ZIfcvAyUi�P��{�N�f�
W�����jh2Kt�ڹ�,bR�E��/jl��ų)C
TJ^61���kChY��/��X{�V�VK�A�6I�Z��p���U�$�u���Ƣ�}a�Œ��Nj�ԗX���n#H
���v5�	<݆�).�s���C��HnZ�t���`�MՓ��^*��4ԤUG��
�	H�� "6��l�S7i���J�J�����+��2�lm�تX���M�W�n�F^�ha2�ёP�5{�1�ӎ��C�[Iǲ�#2��EU��,F�����"yf4Hݖ����Q������]�����D�0���z�ԫr�n}���e��B�.�v�4� &B��p�,�Um��ǂ�b�v����|&{�­ˌ��s��VVD���Vf�Y��d��aa{m<�D� k*ͻ��5j�0�1~w8�_�M)Ki�t�.�sLfЈҊ��SwJ�S�5�u����݀M4/m�8�fk�ɢ�K2ۖ$��Ҽ@�WQ��
�{@�7�R�a@�۫�1�
־[l���E��w�".j7m�G)h"���˕G61fe^�Ѹ��.)M�+oS �@V]��ֽ	\M8�un�7In+/����D���+ �1صg-�#(�wHT�hV���h�M���n��6K�b�Z?4q#[��ӑnl�#�h�"!b%@`u��)���h��+��ދ( #����d4��iʍ�KJ�I��$4e����A�4
����o4e�2-r��f]��~���UwE�#ݐ��d��R�Y�n���dHR�F^�2�Q�t�W��X��R��q똯�ː����f��D�!t0\ʘ�'R�n�����rVT[W�l�1�P��U��w�oi�.���\�w5|��zMj�p�$&cp�Y[YH
��-��I-���غ)li���e�&�[F����W�(]n�\d��(��5�ŕ����hBC�H�
J�����1��hI�j�MQ�P������cQ���z"/+@B�I��J��L�A�ǎ�:�&�#Vh�!�r�V�ZJq\�:�0�RЛ[�)R���u!htC-�����T��mhU+q�l�F�Gi�j�O&1�2Ҹv���.݂��nLy�L��7xr�m�7��'B�NZ�����T�����B���E`+m�X�c$Y�����M4'vU�f�u���Ua�6�uti+
BK�,�c/3F-�M&o�i�Vj�s/P�0ӵ�h�>��D�Or`Xh[.�tel���zS�$�J���B����`��unhÇJ���{�l�t�`Ȯ��^)�-�4 ��4B��L��:Ka,42��<r��!i=�35ܷ�bE��řn�V7D��f����n[��j�7�f|-^E+,e��)I�REc��򽨎;�@c[��6��[i8ޠ2V�卡����H�����V1�;�n6j*��Q��j�(������nbi!K\�����[������@n!�4f-2�]�m�Bd��H��Y�h^����9��԰Dkֱ[��y0ks�]�%�Wvjm)��!0qP�աz�ci��R˛�ԥX�*�w^��E�40�č���(~5`Y����%�&�x@���w�𴊨_���%�f]���*.�7N��<�- 텻��+w0
5/Ka��S�ː��*��Q���������nZ���JU�V�p��q�`T�wq��wQ�-�f4rB��;���<�w&��0�òmmm���C(��*�Ų$.��1E(ˑ��5��l�n�/-YX�බ�š�LUַ���*dAܬ�WwM�m�7o�P�oU��V�Ȝ��\`YyN��D��S;J��!�&X��V�V��iS%�@K��[�4�rBY���:E�"ʹ`S��+�ڔ�gi���s"��E5l-�7���Շ4�u��F�n$�i���e�EAmV-�\ƙ�j�׊eԶ�AvY�pg��sT�J+Y.���hSOQ3E�I]�J���]-!�1F�P���
9M���Sj�y�X&�T�bFk;GI��1o�;�80�w�b�4h3Ɍjզ����[R-�Z��oJ��B���9,;��� r]⎶��uWnn��ӊ�hz�ɰFἥj�#sQoK��
�����	X�{L��z��㡥&�儶���Z.�Ea[�Y��tF�ס���1:L�j(D%S��eaZ2Յ���P��3��+sv�d�!۸��������d�5��K����P���(���z��3d�ƫ�ēh���Ŕ�F�h�L�ën��f2�o+m�or���SוfQԕ�.�<�!d4r����",��&���t�;*�Ow&V�m*0�`��$�ۡ�H�p�����@9�ㅀ��t.m��qM�yIZ.b8l�y�%@��ƥ����$H���:��.P�U�o2�=�b�R	�����J8L�@\VÈC��Е�e�(��C�ا�.�%�fM�ב�Ah�E���4*��*ЭSW'�朵�ۢ6��Xcj�Pf�ެ�n�¥�m�b��%43��&�/�*]��[1�n�^�-0�!�Ź�;�nS����q��֑�"�;y�r�6P��Z�	���H����r�ȝ(E]��x��3U��Y�9 ��t�6��P����S�sjM,������Q6sO��-������	�w�4�w�h�����*i7�n/J$ �kl� �f�9��j�	f�SV�70�XL��Z��a'��`-���5=uy���Oi�{�AE�,����
r��$ҧh�[&�;�#�F��dCeF�A�3#�Ka,�U��eK5�@�kYD�K43a���Ո�|Ȋ4��V5m����AF*l�gRQ;B�U�j`­a���La�L,&K��r�a������Tmbx�Ԑ;�k%L�V� �2�)L+��!4�.T��O�3,T�լxseӗR�m!1E�,�j"G�pP�����
{f����f`�s[%�B-{���a0��2��r&�����Z�7Yz.ՇN�±�'cY�@���\����ZE@�i�;5���j�kthHa�w&1t>�U����� VVU�2h��{i���
Ǧ�[G5շ{y��(^��o"�w"Xql����o7��l< c&�aݥJ)��e��Iu�a��܍�B�Գ%�o �B�ݖ�f�:����xƳ�d�n�D&�^ݽ
�L��pР�%�J�槗�ˏnLvט��칢BV��C�f�*�ɺ`�'�u���m%ov�XU�u-
��-���6�]�K���J�$��H71}vӛ��M�R�[�f���n<ɮ[x��U�5eE�Z4�l۶&(�Ö��2���+��9j���f�k�e�mH�lHD�
��J�Z�J����I�P\��V(I[�����M�D�X���K�m���Ś��p� �/I̸�mic䈰V)������(�lȆ<D�n���L���ʧ�^��B��ں;��2Z5�9Y"�Ch��j�bo;��-iZ��ܣ�{�mG�&Pk�Ұ�h�7b��.�u �d<n���1ʘ�J�k�[��f�3�iՙ�j�2�oD�[��䩊��n����Օ1Ԡ�d�R�n�͚�x5�mV �j.�t�đ^��1�P���bd�@j;KU-W.M7-�XI��nP�EB8i��Z�X�B�r	(���bk�X�^�l�{��X����8Ʌe��8�諧d�ƨK�$۰ӻ�����{�TKwP�=OĲw�i�]J��L݄T���iml���[��,���W5'�����:�f���@����8]M���Z����V=ƍ���Lu��jm��B��@f�N'u��8F8�`����4��y@��dI�FG��+FX;���.�8&�;�O&
�eIk{osCv��efY�i.+�m�~�@;�����JF��Ɩ�ּV��1�U�nl�\o`��4��*Y�Z���:>��VE�:U��R��u����3(���ח�$������V��(�JÎ����S�3��G)���5�L��N�Ң�Z�@{�;ǷyG��ONZS��Õ�?*�2�4���#
��{�cC%;�s��i\�q-'e;OYШABP��m�����9Ln#�B�Q��im�������4���=��h��`qމ�u�fю|չ�{�EH��mTW.�]a�Q��.�VCB�caORyei[k0;6X�*���++`��GdJ�*��;+Rв�ʻ��X��G���o\�5'�S�i���Z�k)f�I *��
�ʘ�ÊLˋKz����Z�]K"�Z;O�ת���:�IA��U�uR��+$(*$X��)&��*�C�*:2�u�v��S\U��jИ������
d<I��y�U`*�tj�.L��.gѺ��,	�`a[��R�����)�(�1=i���Ct�j���Y3>���4�a,l������i�Xt�o^3�)f�UE�U���� �@�+bh�>�CsL��ɬQ�Q8��<,ef�l��*�(-�v¥�4%1�PR���٤��1�ꗠ�7Ma�ٻe
(܊!K];m�֓�k�];j���X�Z�:$�x����Yܟo*��qU�h3�^�����w�U�S���mf�*E�n�@�B��Ā�փ�dBdp\z�J6��:��g
�{x7UCO���oei�4Ŷ��Y��f����ƥ�1:z�BǄ�2��v�L]XɈ}e3-�6�Fc9���͉��Z2�g@Vnf�bT�!�i��RC��.��I��!�f��[WYO�MDѺ����:�J���6KO����C����	m]�եޝo5MT��,֗��F$��y[�r��w�$�  FC�X���ʦ��{B��̘ �����8�Af�.��Yw�����A�#Vm@��ko3P�p#[����&h�I�����f/��Y�,(������C�Zʸ�;v�7�S�J�27���Nls.�`�(Yn�-M�`0�t�9Q��/F�b��Z��p�;����T��E�HV�7�%��̠�0m^�V��h��$- FE.xP4e,�p)J��[r�0υ�Ywd<�(h� �V�^�T;K0���-*X�kl]hJ74 Ev���:Vei�N�X�t�[KT�p=1kX���V�1bD�yK,SP��"���̫�WYB�yTe1b`��jR�B��)�[�X�Ta�V7Y[M�dG7����uE���H����q-���[[lP��Ѥ�c-Cu�X�J&Һ����sjf�[���V�ZD�gp���}lA��q�[f���)C6��`e*�Ņ�~'0�dt���yz���y�%�3M��;:Z2��w�yl��K@/wwMŕ>4�U`M9t
ܳ��� ���^;�y��;$����L:LX�GY��D�p�9uxend4�)��Uzb��CuU�2�GeM��Ƚr�[wy�!̕(��.�
���:LWi9"-��X �%�M�(enӆ�W�:Kz�ɫ)��lT��3.�El�!lV[Wki�W-�Jb�DvYZl��;e��d;W��!��-@�Mϯ�@h�4�B��홷7hUi��u����8�̥)ui۲��w2���
au�	^�U� 6��f 7���h��T�7���+X�	fXde+��V�ֶe��I�
V�lj�-#e��*�"��om�	O#��c����(�E�X��fB�mՉ��j���J ��e������/�"([g3J���,,�M�cX�Z0�q
K1��٣P�&�52�&�J���.[1=��V-���Z��+^�mS�m�.��%�K� �敖��C[݊�i�	�*[V���ڍ��^�}.L¯e�m�N�w��l*��3�4 �KK�^;_��8.S��?22��	��؉����//j�C������n�а��Mnkb�U���/m���H6qb��H9�����Ko��N�]D	E��0At��n�e�C o�3�H޻���Fn��1�{B��0��A*D��ڡѵ2�9�E6�
N'�*d1��,P����,�3@���c� ����z8��ˢ��Vkr�cR�,����Yګ+u��VTɘض��i�$En�=XUd��멥*x�0�m�9�Ķ������կl-Sv��m�e����B��%�R����-=��|���h'CU�tr�!�yC�6�5�P�T�&�Hӽ�`V`�E���+ZF̂64Q:mm�m��kV�SM����8�E����Q�/vM��(�o �6jU��ie�!rnm.]���^T-#׶����!�0$/u��.���N��C�̎�妕2�\r�l�����iL�7����%�u�x��	�y��R�Å\o�<�I������6���	�tS�dt��Y��4�\]�����w]a$�M;�,p�w����%V��}j�n��mt���c��{��b���B����t���.�17!/�����nl�J�P�C�)��oVf���a���U�-�uqc��ӜٝP��������ޕ���2FK����]�V�^��$�"֧f:�C'Z��#�WG��� �� 1�ʻC�N�P�z:�\����/�č�s����S5�;nma�O�
�2�ԝl��R�ݸѥr�W$(��lJ��k�q�3�v�ǒ|���Ry\�f���m#S��p�K.�t2-<�u�e �B�9�z����YY@�b����J�k3�-**SV:��_kJ�'76⮻�~$:Z�W�z��K����#wCg�V���j��̜��Wa	�y{�%�Ȟʜ��Z���0DZ%���WFp�,��Wf�Ձ���+��jL�����)���rv��4{G����εX�Wg�o�v��r���z���e�N��r����Z$�!�t�]�����ѻ��+�j��0qי֫��q���l���.�D���ͺ{�gY��3ZǙV�& �-BS�h��U�r�u ��c�9�IHޤ�����u��QQ�o��N�їx@�KZ��vN���5�q��y(S���Dr�{��#Lq�QziC���n൘���@'�0ִWP�r��B�W�a����}S�e��f���;�:�;����.�U�0��a5s�ټ��=-k�j�M����*���o]�T�����E�l��DŸ��oC��,U�:��
�j�0k��w��Z,���.ظ�q�ۥh����t�p�-�"U��μij<�]�����*�v�֡Y�Z�Omq���Ρ%*"�M�{29��˴����F���;Qԯy(с�������J��~��b��86;i)�;%u��goR��y�Vw-���n3g/LG��8��q�B�n��g<�U�UclA8k��LЦ�����[��'�h�NV�jW bέ��F�M%��b�Т�]K���GS���ڗ��c�%�{L��mU�o*u�R��Vj{��V�%���)�=�z(�6�uaq�qQ�H"�:r��Ԅ5��s�o�t� ]�	D��-�Wr5����p����5MڭW���s�fc��c���Q�1`7R"��)kN�=q�n�|>���z�=�P�Kc��r�;l�y�ۮf9���Q趥e<��n�q��k���T��0��*a_e��j2un(M�3�ʾ*����W{�����ɽHV�"�
]�V4�#'Ê�(*2����u�s+�ޜI�V,e����������_��������MxV�RY�0_PđEl�z��N���j��4�'��Z�s����۸zcU:;Y�f٨3��p�2�`'ݼuu*Z���e�B��,h-�z��Ӵj��R��32��Y��v6*B��JZP��jٜ��Tӷ��Ĥ�QJ�!k�����a�4WF��=��M���$�X�Ɣ�ٜ��	\���2c܏^O����4ʺ�O�+��SF���5�@������f^Wgu��h�tV����uK�|4W< e���&�*о���a�ӵ�۵t2!׆v��tk��2b�Ҕ_N���|��p����Z����W}Q1Dc�����O��/f�w0�N��.�Hۻh�]B�c�{%!�;�/«_#���Xub�#�và��:��,�L[�͜iI(��l+2�F�ҏ]����W+����}GoXaȵ�c�A�zh������J�Z�/&�Օ�Ԡ;qJ˄�7��.�Ϣ����3�)"3p���N�a<kf���&��ɾp�#&�P��qCsQ�Җ�w%�HW�0���F=�,3���L��74�}��8�#������x7ehإ�Ww[���1���Ѳ�E�ե�U��Х�BYJ�DshPH!W�c���ǽ��M�;ZvgKʁ�ԫ�w(�]�}��Qإ�(p��ܿ����W]�Q�*�c]�f�Q�e,S���d�BA��� �v����RҼr&��ZKG&�l!\]k��rѸ!��r��-��/��UBC8q��Vq�Px��U�(�4��f*��ŷk�����w����g�'\�w��^��*{*^��)��1ݴhy�Tw�&�v���޹�λz�[����4M&T3 ̓5��v+�S���x��P�k�Oq���`��(\�kW8����p��6�e�+7,�6�-;�&F2��V�һ嵝����i��(�u���guR��>qׁ[Ws�[���ݰ��hn]����ύ+�����P�,��m����0A�|��gZ���9��yZ*�:�x�5Y�-2.�\|��ӣ�gL���Z����Li�+�&�yt���r�F��`U|p�&�ޮ+��Y��>͠=s�+�y\͑>���/��ь��]�pbԝz�9�/����O�U��[��6��rT��V$�oR��xwi��^s�|�cWU�	���HBM�>oA��>=�5�ޤ�����"k�n] ��i��#b>���'}�f�e
�>�]z�.�ntޢ��D�Z&�I]��Ҧ�"�BdwNZ�2�kA�LA�Ë;fX���%r�ˆ1������+O%h�U��;�I+�^L��W\��JØy�4[���N�m��{xw3�����_o�9p�y�W�P�-Rk	|d�TKH� S��8���vu�]JI�#���`��t���|1X��)Ҿ�75�	ې�wk�\��d�(_^�2��[�o\�'B�l�R��wH���-�Þ
ҐG�����^���x���A93hh�ND��Mv�{�У���(���˒�Ӓqb}��ļÎ�L��|y�Qʹ��Ȩ�N![��)����r-rF�=��7���d�}�<n��t����í���R,2�㗙Kn�ﳺ�oi�g�`T�s���I�[���ʱJ�ŕ��]M�z��FJyK^R�h9;;pV�0���&���*=}+�j��I��ڽ�t�e̵����X�y��qU�JF�/�8�͖��I�g\��g(��f4sQQi�H�;]���+iJ�9��m��� 1���
z��vn��@�u�V�N�:��+UR��B����r�=�f�1u9!�u�j���e�sfX�Q�(��R���Dm�u�2 ���������wwee�Qm��7;�M��RAW��o�|&�V�9ј|q����e
FҮ	_od4��7��C�W��r��B� �jg1Ý��C*\޶�\w�>�3*�:ĻC�JDM��]���P\�24��)��jܭJ�tFJ�}�6;�����t��X��89b(��C��{2�V
6i�hV,?��a:���^Pg��|&���o���˧\ڠ!Q}�f�L,����ĬI/�8@��[� ���S�z�io�h��Pu��䶶����)wu�b�p�gU�Y�mJ
�ܛa�����6���wN�.I���UJ5#.�y�&��g=-�l�n�
�� g1�'V�2p�MY�U��0���e�|��Tl�w].�,�J���c��	�3&����J�k����;����v)A3!��*+H`g�q�6��:�4K��N��Mv��S)Q�#�.p'۫�%���N�N�-lS]V���|��;���r=�Bl�V e
8l�6r��� c�#����![)���b�Z�C��j˕�a}Cz��_2��0�en�Lb�m��D�4p;���{a����]j]��09��U��d_���P�go��	���m��5���J�CfV�
1Y�j�U�Ր&�M9X{�F-:	5���w�������Mk�W�K���J�Y��Y���`�}5o�]�.*���ȭ=OW ��/�7rLe�BR�yj�X�����	p�
�l�v��;AZ�D��6���S�p�k�]b�}ٳ#�������4s��E�vԁ�uw}�h��;\5IYJ�o{�\ͮ��g�Bfh�I� A�+�J�$ �;�,+��)�6�1�t��Y��<5�o^ Ү�c6���oF孛��Qq��n8qw*Ƹ���EJ�Q���2���W@垡��ZS�3:$�.�����2����)ӣ�$������Nև=���Z���&����۵7(8]k�	W�~��@��T�/�R�|A��R�����x���_!-�)>=ؗ^�)�,���ΧI�
�59|��^gWZ�(�������CO+Gn����z�Ea[C��SM����V�Q\�X`F�$�Mo,^g۠-����~X.��F���|����x#Ӕ����o+K\�f^i��:���J��tpBgwb N���ϲ���Zj�ތ>��r��a�oF��J� C��]�<�w�=��+�@V�I�f���fR�Z*Xˮـ$�Yy��L��k&�f��M��t_v�	,j��W'��(4�l�L�' ��Qcs*ƅ���<@�w.!b�`(5���
����1���QT�Xt"��ڵ�u"��'P�-gG|��w���2�6�1�a����Ko�4<�p�KMu�:t_o6�SE�NN9t�wk#�]�e2�*+�tIѸ�(�m����ǥC>ώ��Q��F�
�]]�|7K��;��t(3-�i7ɑ[�`څ�����\���R��E���2������xS�H��7^��p��!�(�Ι�eX�[EW`�q�, ¹�y�,>�e�6������O��,�n�X2��8ŭ��s1��+y>c��ư�jNRˮ�n:v�6E�(���j�t&Ĳy^'����hb*����
��T� Yt�T��
[�ӃPBV C��bv��s����ӓ��Ff�DI۩���S��5�!P��t�\�v+�uΖy��a���9�KbPZ���`�zr1kB��Y28o\��t��n�F�V��\^�o'W��^���	�o�%�H��f��ʖoS��AjJB.M��*�S��;�:�	tM�N�kw��qQ5�E�s�f)ݶ`��-� I]Q�[Y�o����f��Ӿ�q̫*�o>YMN�5"�јgF�9D��x&����{���T���B:��kq�[u�;��Sa�W��+�{RhХ���d�V˷� 9�A�W���Q�w�	�"�V3R\�շ&���o:�/�L���E�l�J�'�Ѫ"����������yfdqW����p(9�s�N�@Ӹ6qod66B�X�yM� ���]��=�\�tuqt\��"���@��d��u`�pԾ1Ω��.���!x�3j��8�����Nw-�Z��],̬�j�r&+�����x���V�n��>���.����i-��f:�)�՘R��&k�/�3���uՙ�>Elٷ�9�Zt�(>S's�5Ǚ�'uHi�4P�=��N�{��S3�^��{��w+.2F����S�w'��"�g_c�(j�B��0�[�@�;6h(r"��[Y�i1�;�eq��7�D�ؓ��j������e��`����+j�5�s���YsG8�����g_)��y>��f���f��X�Jټ4[�չZ���������{;��i�޿�Vl<>:��l�'<�\���&�4�H1�u�I��#�Q@�3$єNΈ�����0��.� n��<=5�Q��w{[��Fج���T�:�Jdc���o���|��V��.�W,P�z���lr{\�1M��%Q��X�W-�j��F�J���W��d	\��{֜��]��)��s��av�*��n���w��]�r�s6��Ʒ����R���N���QM�呝��H�Żt�|g-wv��sf��5�B/���D�e�ú�)�����FY���Z	N^����k6
��W���!z��+
j4��	����R��/�N��Q����Z��I@)�W���F�/����~:�l�o���a�1.��j<K�9�J�Uj&m#cwr i��s3FB���,Px$��$좒�Q�k�΂�u���nJ�K�f���J7t"�!5&X&����2'�z>�P�ٕ;4��H`J��F���C8�3)�0�h���*��T]:U�k�e��z�w\z���ýhk;�۰�'��(gdó��ʺv��zY|nj�u��g�8�̲W*�y����}P^�ש;�iv*��CYZA�+c����ws	��wGyٷV9�Wa�����۔�j�S������
�m9����Q��i]�t���p��y����p}�4���l�5Ҹ�M���!��*_0�[�Zʇ0�t!'Hhn���ZV�w��y�%l
���E���X��^o�����|��v���1�M8����3���Jy�\�Os��H2��Lt>43���d�<�H����3���XV85����)��8�/.����
%��u��`el�|4nR�vbݒ�� ҳhv!����S�t�9�VM;K�U�m�RBE�Ah���:�(����:��=���x�!P�����W\5�L�u�a�F�@��m����Qu�3)�Ld�~�\e\Ú�E�p1Gf��ġa��_-IB��ꕜ���'no��H�ܫ�m ��7��sf'{�)���- U��ԂV����ye<��N��@��J͉�������ɸ���E��Gu�X'}:���p{�"w�;:'�*�o+�ķL�Nw�oc�o]�b$_d6�*eL��r�K�$76I��󕵕�k\��y`��.�&��y�'�t���gSK�Ün�����m.svpY�r�'�J6��H+������]Ƥ;��}�}~�mkmj���ڵ����������_^}��[�U�<�M][THu}̪���U�Ӈi�ڜ)J���W�*�]�t�6�0���q��j�z���jK��m;����G��<�	�X���κ����}rsD�f�9*J�J�r��א����n�dj�Gf��H�He�d�)�zl>�[�_��_ΐ����n�%I��W�c37h�a\�5��Vo�@ب�M�]��Qm�D2��[�\]E&xRY�%��n��7r]�sa���/$"X��u]�f� �S�аr�Q�j;��#���9cvݷ9�<[���U�Ѵk-��n��V�mJ�(+Ŋ8�AK]	�j�7�Ja�z��v-�ԫԲێ���kq�z�=Y�,T2gS�\�0��֚���mfog�֬Eĵ�����]
�X���F=��Rl����6aX���.�Hk�-'yar�F�F�E릯�(�a�/�ke�K��Q���b��.�ڇ�Si���,�[�G��\t���%����y�^m�]�)�����MػI涰��ᶔ�4$�Bw�6�6�tPNem�W)�i�;Wm(�q��N��P �흆� �E,O�=����]�0\��vƶ���)��I��H�-Q���TV�]cv*�X��}c�aW��X��C:�v���o80��@�$�;^��`���W��2`�;�ʓ�P4nr��"N��0K<ֲ�X�-�8�R�or�(���=���k���ܒ ���D�S- �݁`-��f�ʌ�A��4�<o�<�Z[-9�{�X�ϻ�4��]���z$0���t��|�Dئk�y1��5��ػ����]K��M�6����6̺���p�C�h�p4�}*�-��4n�r��X�	4CV��ߝ*C)'[Yk8���+�n��oEs�I��ԶO$�̨Wҕ�ܑ�z��w:ʫ+C']�q�^��۱�k���G�]��tH����b[x��,��BVc˨�;�&�l�L�]-�ٵ���p	��|�ND�Ÿ�u�P��!J��I���8�xF���r�8+E�q �L�3f�c�Z��e���ɤ�p��ϲ��K�Ν�����6l���u�<D*�.�i�B���@�m.z�ܙ�b��9���v:��Ka�ݼ&�	V�U���\F�]�.Y�>�l�Ѯ�P���
��YW�g`�-������}��Qٝ����/�i෋7+*S��]��kD�����k.�l՚�U��9<B���c��f_�-9����ቓv�'w\5_d�R��(�N̠��P��V[u%�V0[�m�¶7M�A���[̼0��B�T�� X
��ۺ׃���pr���U�c5����)Q8�ػ��8*��9��n���,�; <�'�:=������ ��fޚ+tRrK	�i3�hز"�r+b�F�'��̬������JdP�;:v���(V���dzRܨ����9W��Pk�q���)}�����؁�%E��պ��.���v�"�]��m	{��)I,d��e�������V�gf@�`v���.;z/�*�R]�R֮�?�#��@�S�ӯN��b�#��J�t��4�6�^nE�0���f*�i�C������t2���s�Q|�`�寺��0�����[�;wYh�^��q>%��l�AU�����A�)U�i^f�k9
%�]ו�܀Ą��TҕaMd�x�����wk�}��]�a��P��tM��	�����)�r��'E2�(�p˒Q����]C�h2k�ǸK�X�vm�^�w:�g=���`QX%^�V\cI��&��N㧵��)NWh�RY%u.�؏P9���
��Bu�bP;�BG@�<�2�[L�ۼ�I�ו;sDk�w�ic2�W����m]�W4��Zxmӷ�)Gk{d�n=nqEVw��u�Ғ��F�w�Gׇ��l�Dvc|0�)�8��ge����̵�v�3���D��RG2�蘐g������.��bžV�w>����i��3�jnGtև�0���^��%e��z9*��݉�P�]��oX�B�5
�Ku�g�`�`���O����rm�y͎�&��{ݲ�"�k�弽?6��w�����^^����C��
���CeC��~�]���ݴw�j��Z�5Փ�#�z�Mb��ߊc�3��dy�>v���@�Z�g*���u�������j�X�髶��f���T��ͬuaj�!C.^dKV���ˍ�O�V��˟G�f��E۠�����iB�ljDC�$����Ip�a�]U� �k�P��y���&�����h��!El4\���t�uA�N�@��&�]ne�r�e�p����WGc��o`̹�/���H�]��ѹ̇Z�vHt�|Vt���h7x�	Z�p��BY��b��#�Wc*:�k�%�.X��l��v���:N.�e����PR��X��'M��]y ��%���驪���-:�m��̬��h�/�_fK��NS��	㫛����n��┩,Ȁ���#�O[obx���u),Gz���@�	��4��g�Ø�T���J��h=�mԥ�d@��E<��rdO��x�d�iX���Z�ܖJ�Ԧr�ġ��������A�n��+>��A�2���z�Q�e� ���u`����VA]�
oU,=�v ��ej��8�����ٶ�2��u�ݲ~PRkql4�lls��cCՍE��F��+��`+h�/�< ���e	��P��^#Л�e�̂E'��-�B�F+�!;Sۻ�c�l2.�8E4�!������[ڏ#Ұ�g0U�fR�9U����Ơ�(V�[w���Tťrӊ��1�{3.��ӊ��lQ�a��_G'i����Ve2Uu���2[�-��Mm�9.pԧ�,)�.�
�Z�Z�)�\�P�G���]�J(�v�ԣ��i�S��nS�2�W-�&v��xz��t��^�jg�x�D]�ɺnԑ���IR��]����{��,!��t�"ډ���W9D�ٗ]K���r���|J[wқX�؅nr���z���R�/��M��,2�؅q�Lƺ�u�+���8
���9�x�3l3�J���ou�$�[*m��]�HU��9m'i�!S(������W'u k.]�]��d�I����7V�G�Y�����	h�����.Z�>��zz������^�V�o�U�F�����!9�� RW�"Z���콕���ŖD���LL�M:�Ǐ/�t��޾Bk���[z�.���ҙ�h<�嚵gG��Tc�� t-t����ܸ�_E-\����`v"�,��W��c��s�������򄊎�^�����o9Wkl�<d���K�e��ӎތ���� �o*`���u`�ve��*��;äi�U��+0IS�*�m�[ۂ��5�U��U��<kF�`mq����fj�6V"�L���-���gt엄-��a�ۓ!r���̼ĖN �H30`�-���л ��EW����67Q�X��t1���^ݥ/x�jS]|�f�B�˰���\�"�D��}}�.����OU%�ŕ��[R����n��gd��7:��Sܲ�rڡnϋ����Z��K�w��͂"ћ�`GjJ��23��ޤ�Ps力-�9�(���A�� ����yb��Ϫ����.�Wj����W���A�Ե�i�Bۻ�����\V�H�����@�L%�9�%�t��m��mv�u���ŀ�N��W�v<��\��C��Y���2)R�im���d�T�eJ��x6�.��F���-v��%�swu�R���u3Z�5�����"'�����U���y¬kq��u�2V��'��ooBz	�C� �/�@9��@��J����j�Vƥb�D7G����}�Y�R��\9�"�6h�oWvBՙ�Ԥ2��$���{W�vSs�5����ø#��k�����cc[}t��S՗jh�JQ�+6��vTOE�������躶Z泫��H��޳��Wϖ�T(28pGk/��`��1��eT�lz���֚ػ�ڹ�
Np�Ez�Tz�Z�/��
O#����+z8u�I��v=�C�LW*��΢��jt��hp����w���L�u�g��.�h0�jA.�Q�����|`�n�������_-����{�k��,œ"bP<�h��fS�ۋi�������FMW4-�negV�H���{êt5��P8�#1���Vl毎v�9* �j��W|�i��εKY|�='.�Q����P}]���f�k�8�;.�#��ܩ�wtP7b���� n��K����_].�h<ۏ--V*rR�w��ꩋn�-�x���m��e�.��r��2�`����`����r��1�7-r�(	�G|!�*m�t.�KM[ � �][:�zfjR���$���;x�6���֕
:#�:�k�]�s�x�K5ۈ��0���l'�,�]\���[]�A�6�l�{��wrY��c \���ˏe�u&[�2m0g���KVK�k棽!P�W|6���>؄�k�ܺ�iz�̼#ej��!��iV�/^�&Iv�w�]�Ⱦլ���]����J�V\}d��=��wA�X��f��h\�N��������a�HoZ��ى��h�1�)�g2��U΋�R眩;�a :��綨hcr�e<u�`i�!wY����V+�Y%鱳lR��MD6��J��֊��KZi�4I�%[&����;O���Z����F�t�;�ͷZ��|{�>ǖ}���C�GvP��U�yh6���Ξ�9��λz�E[�D޴��jY�Z~���0�G.��l�:X��ȇ[ǨS�5wP21��I�� ;'YH�A��Бl#z�<����}|�����KQ���k�m6��W*ފ����jL��ʛ��h����+q���g=u��e���քr��v���v닒��&,��%_rs�i[Yt�������h�W]�n������]��}�)�7:�ݪ��M����wtmͱp4����@�ƁG1_1PKn��1)QTX핝L�q_dw�eһ�iZ�K�]@�d��K�L�|)�Yo�-%�V�2�6�I	��p���/�����A���[���˛Q�,�O_}���\�n��L!�D��j�>���vSZ�l�iiAqQ
�-���yO�.��=�z��gqy��4GǇ|b�*���Lӷc�;H�m��s�N�Z�V&�v*NrDQ��nY��D����Kp�<����|���s�
��Ra= F��y���>�qG����oc9�Κa����e��Eݚy�� 4�y���ے�W��9�����Z�&�"���gS8���t�fn�)bw�J�)%�Wr�p��P���2L�.&�@嵆ڤ�:; �d�E�b���<����FF�<��H����<��x�䢄!��f<�}�\.�n �=Q�u���Ă�O�:o�ur�슇m���w�p��<�ݡdʳaM�:���TL�]Zyφ.��0�cyH�w�㎴��SM�,J�#��6T�Ps��3�]�5q,�Q�˭�i�9��hQ^@��ѬfQD��ۙ�ʹ�+�X�V��Z��ڸƖ<�i�k[�y6}P觭>�J���%�B�.�G����@�/6�Y%����&�'���5��uݔЖ_����})�:�ְti�A���뽘��`���z��)�D�����ԣ�n(�.V�v��nŹ�O#���n֦���}#�_a<���m۠K&��NN׏!�o��wKR�����'���;�A���ܬ�����8|IѺ�jf��H�f)��u����0ͬ�݂�4:�b�;ْ9.�bO;N��=�+%`�b32���"��Y�,��ٛuk�KMb���9��_}ֺ��r5�έ6��b��FZ��ѽ`^��hy�)���Vq�ٹp��[%��h⧶�u��i�Z��u�2���ݮ��p"��"�U�u9d���pj@<j�ɭ�l�{)��@p|���cǂ�a�C]�����s��=���@���G��z`Fݬ���]�s��2mi���JT����׃����x{xᙅ�O�m"���u�ۈ�(VleP�[yl�U�|,�³�\��� $������$b�EX�c����Ҁ�-�]���/�c�}�3$P@���-�s�ۘGWԮ�j-;���!�z�V>�u��/��e��,.+s��X��Fu�B[=�ۤ���hoN�%) �z�ř]}����Иh�.�i*0.ߕ��N�=h]���
\�cG"���Mԓ毊��9��[�L���Զ�օ��9��V%;X��92X�x˝���Y�9Q���+]�ʀ!�l�u�6V�kY��M\w�K+FM�h�ٮ,
�͙9�YyT`ցD�;q��t;��$�0l�t��ٰg1@�&��$%�y���Φ���4,7v���ؖ� �{�f�Gj��1Љyz"�l�wg_aH�.��������:�����i�у3���ɹ��#}���o���L��eB�4� 
W�i�Q��p�Յ�`�:y��7Փ�;��dt���f8Ţ��en��
���[F���}h`�<y0�&P��*��ǵ�m�9v�maZ��)r�Kv�U��!�{�4/k*r�"�m�1#���t$�m��嬂X�e��7��z���Dв��{ݜ*cx|�ãm!��>����Om(x�"����[��� ��9�4��S�y���
�׏�)�V��P�҆=���#��L�����
�[D�'h���{{Vo``�zՊͧ�,��A���BT��F�+nneڬ�z錻�BPߛ�
�*�ع���ƺ�*�s%ml�
��I��Q�J�y7�*��/%���+�5��Fݔ+;')���Ǉ��<=�o�3.VF�m�-Rh9n�KC�xog��Q�f։4����vf��to��AS�w�f�}{!�LkO�vV`OMu%�̼�FT�g,�����B�or'+39��u��ѷ��tknօ)s����,99mݧ'B��[�2U#s�\�Z�GÝ^ͽ	����G�ÕλB���N��c39�U����Hqu��o��MJ���X!h,d���]���3R��b'�4��	��$�ͨ{�]"�9�5��/�u��7�K������V%Y��Y:P�h��E���|/������:L�:�7�8�|8*E�uՈM@:�Yӷ}��Y͝\�܈7�p�*�t���7�%�d��7j�������vR��8؊	�����9l�vAݻ�9aw�4[EaS8����Fj��P�sX��ԓ.�V|��XޥZ5i�)kNr�/�_D���,Ȣ�K�ۭ=�[��b��)Hn�^_.����e1uf�Vl()xi)+f���0��^�\���\TN�a)R�+
֎�hC���)�OtO���q�)�X��+vj�^n<\y��ͻN��6ƪʙ.�)����6����[u�B�b�G;v�.=��C`r�� �(7BYaw�'LX�R�
�$�T����gG3�g{%�![�f)�,T�j]���y�uҍ�Y�
(3n�mq�־��]���V=�}��U_B�
@P�i�����H�DE�D�$�D	�Rd���DL�̘�	���dE"a BA	�]����t��iJc)"s�eJa(��Q�@b4D%� VS ����Q,cb�1�$�jd��1&���U��D$l3dFsr�(��X̢�̦AJb"��lL�.�TE3%FL�h�]�H�@��뮢��4�c����ns�(`���R�P�	�3;�-1�t�Q\�d	��D�ҊBds�1�A9�J1�"�%(N뙆�M�E�H؍F�gv�) ��(4nt�E1!,Q"c"&!�I��d�
��p�1DE�Gt�6%$I�X�t��g�����?<����m���S���h$�Zɀ)�$��u;��,E�gk�X��h�5��\*Jǎ�5׳��כ��>�-��<�(����gIT�.�*T{�B�E�r�S��ݩ�8��{k�C�eܰ6�����Y�a���Z����aAa�~�kc�=p�z��1�y�k�X�w{dC���w��L��{ț5�b"�u.���}�笪�zW�W������KgH�����:�x"�9��٩���Nh0�\�#BHT!��4��[I�p�GFS���{�t��Ng��s��wc"�C��;��xA�xkE�3�(�+��`4w)�{E�ctsU�
�5�	f���i��S?Jd�7!Y�t"6j��<�y)D���{��s���"<F|o لciɠ~:��Y��xL[��v�<.c��ѥ������o��k�˘f�Kĕ�f�Oc���z�ҋN5��=�avuxkٗ�U9Ɍ�G�y���OF��	vrT�c���mL���¿��B�Q,p�x �˄B	s����ʚq���R�ᑣ�;o�pڢ_��Ӵ �߉�+N�������~��O��|I�S�Z���Z���g�ՌA�J�d7Cj@�Ag��V��/��ZD���fhO���x#I�������
���+#��Ş�5�U4�jכ$FIe�o��޹�F�)��#>��d�X�0a�㚱٣ة_^tY۞Ywh|�i:�+g�!�ӓ�\:�e9��S�I����9��=�������{�V�v沚G�!�' \�9
��&zzCh���{Ju}�� 4��A�y��ڜs�7e-���s=G�P��@�����T��Y�kG�eԸ���'ǥ�l�"��� �m���$K���߶��N+����f�Tڱ��#hME-,�!!�������&2�0�U�4�$����k5����?[�]�	C���T�\Oʁ�ί�Ǳ�r�G1�o��Lٶ��M�P|�1�[��g@g�o%{Y7�9TɜB�Lc�:��S%��0k�}-j5��kwS�t�U+�]�Z�z0�d���t����tzʇ��4�v���]�wVfL�՚�y�P�)���I��G@�ݧ.Ƒ����_dd.fP����:pܙ1�`�1:1�
���烩��+�_b�n�d�������W������RơX��"���3�ط\�/i냜�}瑡'ڰ��Um�G���Ua����%L��N�z!]C`9�ԓn�6��ԖZ���G����7è���hvh=2��%�*$��^_Q�:�б����������wq�;�Ww���+�`�7;��LP@�G	��%��M0�'�xo�Z��v�]/:�\�$;n�2�k��,��39*]o�}{�ۜ�Tذ:��Ѧ��q.�ʊ� ��	O3����¨��yy��~� ��d��ב���]6}�.ah�|I5������5F���j&J�����2nu}����s,<	�a2��� ��ف�
�#H�3�Z5G5)�JUc�vV��j��D��3�!p���N��z�9��~M\>ϠU��3;7f.(�R�6b�$p���US�CBѨ{&]*s�p��f��a�H�e	[rZj�u̷X뉽�st4��:
h$t�<���Q�������t�e��K:��N�e�d=��ٮ2�q�Q3��sG����:����bʲ�V���o|��:��TFN�Ef��k�?���\�uE��D�9!=m-�*�$	G|%��M΁۷��e�#i5``�M�^����"0�}n���GL9���6�9$8P�uTR������xLS=�D�Q����I���Ը�ҴF��r�D�:j�s�A	�N%�N� x ;�/����p�TIf��e���)��e-
JEC�1Y05�c���
*t�.�q�۸�u�pM�g+���f�R�=�x�ˍS	��'��Y	��Կ<��ٵ�tcz�YP�
�	}���ѝwV��6��	�Vzǯ��ڕ-��w�N�ymg���ݕ�.^!���^�d4�yՉ��oA���J뿔�$���Be�n������i����拥��3j��h`M��!����bBh�9R[����K��Z̰z�!m�7Y,��*.n݆=DV^|�ܺ� l�Pl¿������ɼ�L_ٶ�Τ�Yxe��i�j����jfz�M��q����[�Q֯f�P�*��c�S��ϩ����J�ezz�N,+���Wк�<�X�L02$�!����uf������PK���C�B��dZ�/4v���\e*�ڧ2����t�r0���/M^Nw��0l�½����]��VgY�w��,?}@�:'���G<����-�3n)��C\C��� U���������6�L���g�(��C@W�Q�|@�s{d�u�7c�0�87{9�*�����}wc�%�6ײo�&�t����-�ǻ���n��^̅�Lu�@��
,�����c6��r.��݌�*�������"wHڈ�+MxS��WM�������`Or���T[��Q�.uK�(�H�a��^�f����V�����T�v�
^#=O\��Y�Yc�i{�]i�֑���a��h5�/��Q���j���zіyn� }z��՛�'u�f�]�YHTu�n5�U�`��>���oEi�3�v��S�Y�A�C�ѐ�Lƛn�ܯ'�:���ӭy�{��횴}������fN�#u�l×:�ޮ��;lFz���ف��b����X5�X�͆�������]�F5 X�@�Fn6ч;9i�O�ˋ�(6�1�ZC��QU{-��I����r�z�tF$���&��B���G�^�E�i��V%��K�_�h�C�u�U�׻��9�92B������{�B����X��4��ۨs��aLw˞ۜ��l���4�4tD����^����t����k�UD���^/��,��
��S���v���U9�Gw]â7Xb��Ʉ�ތ|��*�4\��˂Ui�%pׅhF.(Z��ԣ�j+{�2>~��Ҽ�|����z��xP���T<sg�\Ɂ�Nh1Eȱ����R�nDH�H�o])�o���j癮#�*X��TɍƲ�2]Ø�f����7$�J^[�!����e��X�qP=�U��|�ٍs�Y���E1R�3����5g����uI�C�H��4���F�����n^�m�	`��K���͚FK�<����?g��R9�{$�W���*��ȃ]9�'dʲ`�C��1�-�`N�RpY߁=�7�7�4�����o.�$�dd��[K{%EQE���k8
�xz3�7�F;\�+�,ֵ�*��K�(�<4i>�+�8+�V/���0;�y���e�$ۤ�q�׻���f���ٝnΡW�o��Q��܍��8Z;�����MC�~�
B�Z��)Ƞ9)����*%Z��v�Pq��/.1�6"�E�Z��Z8r��k�֗�/�^�//֬��Na~���T!�ՇC	���,�yu�>�]�쑦R�[>*J�����G(��q���<�.+�|�&>���ퟪ[7<����N���?a�P�P:���v3:���{��,�7��@
�d$k�Hx��,��Q��ONDSj��w��s��p���wk5UآA�as���jm��ϫH�చ_-��ثG���:v������6P�vm���Gt�ŕ�.jP`�o�!Cƶ����$O�c�2�.���9/������,��c1��Z̉���9r�V�>�C�������=Ḳ����ۊ0��U
r�w:��;�|���ݫ��m�X �����h�I��U�S6�S�xAݫD��>�x�NW=Yrț�/����8 �CVZJ�ѫݧ]��������My�����vۿXV�Y�_��2��}1k73�8H�ޤ�i��I�����>���N��B��C�]��a�l*<�#/}#�ZL�]��+��S�.]Cy��;v�@}z�IMoGأ����(!�Һܜڅ�q�	&N�o��y�W�
���:XA87R��R�E��7"�/���yJ�u��{X~ݥ.�i.ySێ�����g�����^T���סD�ǫ�+J�S�0
�C���Z��������c��ʱ7	�c�n�n'z����y�g�=��Ѧb}�����Ҁ�c��0{�e����3��-��@�U�0�m�p�B�ܞ�B�.���s�݌"}���ۦ�:�IX߅i���#~=Q����oX�vNL��t�}�/�=:��f:oT5F�ZH4����1݌��]א�.�zv��WuH�k?+�ˑa̰�Zt�Y��� ��ف� �6�M�X����NM��F��puX�G�%�z�эN��k�T�2��������l펕�;n�+�ɝ��My!Hy�I�W ��HO�R��>������C��֬����'�"b�]��@{��n�_LK��QV�'M}��*�*=�	��B��m=1N���I]��}Y���9�4nY�IwJ��<|�r�5�B�+2��{XWש*�3�`�����t$52z:�]��שb64\.�E|���fP����j�qv��3�ô��%����^*V�)ɩV�}�@�:�>���"�M�2�(�U��z�]��M���^:��,�. �ּ$�^��[�eH��]���ֆ�HDj��1�!+���[{����#�H�[ຢ���prBc[KqJ��������Lv��Zy�݇Y��\�I�����t�Pul��*�UT�B'E@��s���ɖ��ޠ��o/y��
�4�Ҭ��7�mN�B=�j69�`�N�5�Ҍf�EC>3Ӎ>;�nDW�y[��p��/���ӯ�k������:����$��� �]Sàs���I����kJ���������fx	����c��=�uע��ݟ�nS���K�	�CF,�ǻ{�f��-����������g�B��x�`��2�c�V��PTUz��gh�n��{9D29t��v\D��U�6~h[Vb���{'�P&�S��K�>+�ס��\��[.�ݕ}����򪈨�j��Ȕ�$�!�����4|Ȍ���ER��T,i�I)y7���>�ΝYmL����%X��L�U��Ne_�9�a0�S����f�9����TVdٜ~[g���s�J��k_8+��r�r� �T����v_p*�"�\5mt�<�U�dx���x��ٝk�)��_=!vq�g�M��sOT1�X6�]��N�����:�}!3%���b;��.���e� 鲝-C��|˙���+��K�/+y]!Jx����A����>���ϴ3�ɷ���:lv8�{J�*�wyD���==�[7���#^�����Y��+_	Y��t$?wR&at�r^��s����T���o���٘��TN��>�R�g%�$�G��	|!��Y��^�E�4`�юĢq:�F�����(F�c3+E�=dd���'^��:G��5�Sw�q�)�`kȬ�o;ꩻ6۸7T�b�-c�Z�D��=ҍH���Q�:�y��D���<ۤ���&L��g�4V0�2%N�0��Od}I�b0��a	#{�U��g���[�i-�q�ܥbۅ�ܖi}Nr���7����D�r��O�yu�S��a��"�
�%���uhw��o6�mģEE;��!<��'e�˺\"��K{�J�/�}�S��V+;뻠��:����y��N?���:����8�;���:]�0�dU�Vd��\��♞۷�(�x��8Ƕټ��O13�b�3��nn^���bG�š�o���t�J,J
�CMe#<�샋&�"^f)νDK�2:
�bꄜ�����d�D<��+��qج�MM=N!�鶉�Yt�r����YCr����\_
Uv���tc���!QSz^3˺}4�%F�B Ց�w;�A�{Rȅ�K�iwk�-s}��<мs'7n���{��X����V>���r	��bW>5�Z�i�Y�E��׏��4��;b��_�ܛGYHԘ�ε\*�x"���.���OS\(�!�F<��ȫ��^�~8V��������ѫg�'/��Ln5��!��á�o|ٹ��;?[X�a�dF)���7�����QU��i�8���0<%��M��(_Nw��C%��f��&Y�{Z��PjǺ��*aq��u���-��~����������]�ɟ���v��eLu���svo}L�uȳV�����xe��U�>�RV���y=�[C��4�U�;:So`3�=�n��M��*�������r��R���e��l�a4�����.i����$�N<����	qUb2kDJrf��o�1,=�)���M�PW"�p1�&\���vn����A�����y��#2�Rb��6>�ZN��ퟨ��NM��i�9����s�P�".*
qq�z�KŊ&���(�������S�#�L����ڿ�]�)�L�?D}�
f{�v���`H�����9����+�K�1*]*t,�j�3���W[Y01Hݐ	���Nk�Bx�7�L�=�j��3)m�k�Z�����c�rb�p�a�YǱwd.t_݊؎�+�_h���t� "�f�����ur;�&G���rĈY��K�{Z�Tt�z�'���d���1�ڮ=)�M�պs�mf7U�)�+����5�uAW˱�a�,M�s��!�����w�U
��Z���L�l�_o�'Q�m"����5}�8r=��mg2oV��^Y�=���5ǫ6���	�e��
�.�g,��^b�����/�诬$�U;�r;��o�o+:�#�;-���P��N��	1���Cj���i��}#7��CX���]�<�9\*W4-��� �i�ؙ����h?���t��Y��t��w;�v�[棶������ݢ{^��%s�堘쇜�fJL,�����*cԜ|[7�#(^3)�Y����yMZ�WH�^���P�
}X.<�w�#�6X7R�Y3�0�;�\� �)t��1��5��T+]	��E��F��_S;�l�#Y�c��-,�Xz��-W�W2P=ˍmh#T;.1]ڕ���دYo�v��ҥ�(Ͷ�At�[������[˳U=*�5��V�m�'�U���oIވ�=�	��T��e�/�BwN;j3Sh+���а7��6X��j�:�T��9�a5�nM�;�UbP����s�]��ޱ҃���I�3�A�Yz�.�"���n�PFL�iҺb@���
Q����n�f<Ω��i����$8�f�6v�:w[�w�G���1XM�m3�)�S޾Yy���,\��;O#쮡���Ac<�跈��m���o�FG�2��m}W�ŦWf.��p��e�]�8��Z��
u5\��[ssz�n=�!n;R6�W�Bs8v�;9�m�,,L�<m�q��y^D�ޢk����u^h�+���ezf�eav����+�fk�V��b�u��RQ˛p�w��9G���t.@�ؙ�5+'��c:��۝ԓܺ�l��{4�H�ws;��lA�)��}���X�<�)�4�
ą�Jkk�>����]�͈��O!��t���Pa>��]y�c���_U����/e�t<�o��tLX:GJ����{bS��W����i&v��O�3��Zn�E���)�*�OB����n��Q���fiN�ή��SW	mn�1�0�g;5���WOr>F����9C�*g5S��:ͳ��?9-��:�8ձݽ���2H��g�]����7y%�Mx�x���]G"�^ۭ��B���|�_7n�#1��.�]\��VT沑�1/�%�M�.���	j㶱�O'm^K]n�Y�`���/�Ɣa�.Eq��;7F����$-fof���x�"f�B��1_s5�t�P�wxVKZ���)�-����`�o���_̖(6$��%���,L�H��H�T�Db�W�k����CD�wt��A�k�`�&e0��H���"f��$�	
� ���pѴj$�ȒDh4���P����J���L�"b#�H@3,hd�@̚�Q��2H�b1�E!(�H@����$E��#2F%��,S��)BX�M�S
K&�رE���$Sѣ����"&Q�I1E��4Rf�2HH3X�"$��`�I%�a)�-h1i �*"E��A�c
Lƌ�4h�(�0��&D�P@P |�:{a��f	ݘ;�uJVߠ{L�`��(���-��I�=�w����d�H�J�oa���M�_�F�b;�y������^���_�ɯ��_�r+��[�7�W�ֹ��+���m��h�C~^��� P�c�I}����Z�������ܫ�����Ϳ���ۦ"k��w�Xq��g)�"�q7�y�����������7-�\������߿����wo������~�v�u��c5�����>ux����:�7�z���������o{�ߕ�/�x�����;�h����	5Wz�2�[J�G
�/����W�������鷍�/�|����y��������ssn��{��r��˛�ί��η�xޕ���ү�4i�N�6�/����u�ס�ת�/�\�l���D<���^YN��ڬ�5[��������|o��������M�_��|�����Š�߿�W��+����=|�}W���o�|���k�����W�<���oj����������7�ŧ����������0"~�}RK�OIk�/b���;Ϸ���ۖ�}����m������V�o׵�+�;�}y��-������[����_����W������������W��^7翾m��Z�����~�^߭�����ֽ�z����~�¾w��o1���w��ڿEͻί���->u�׽�z�ە~������/���+���^
����-�\��ߟ���?�k��n�����o���Z7�����ߝ����߿|����&c��Զ��Ǥ���GTW?_oM�۾u�~/��ץ�ok�}���7��^/�~������G?�����_�ν,}_��S��/�ۼ��_����{[⹹�~_�￟�E�����z���y}���n�.��ԞsZN~؋La�����������ƍ�����ߍ�o�����{k��߻�o���W���[�^7�x�+���u�Ѿ+�x���_�A�=u�^��+���z�|�}W�����LD9�?@��L%8�.���x*�]R���#�@D���������1i�W�u������W��{�ݯm�[s_���^�ݷ��m�~u��ǋ}W�߮��-�xߞu�W�ѿ�bʏLd�71?D-�6xyf}>�����b`�7:g� >�
�
�T�ﵯ����7���}[���/~}�zo�{o>����}�y�h/����{�+�\��������͹���W����m��~[�<m��\ۖ�W>��o�������߿������ZV����	�2P�����U��YwK���6�Gy��,I�uԒ��{~rb#�_�|��c^T'z�X^ʵ��)�����齝�^@z��*�]ޢ qҝ}��C������o�[��@��w�7N+J��;fV
S�N6�u�׮nmq��B������}�=�~~v�����������u�x���~�����o���}�_���yڽ�>����^/���wϾj��Wּ_����꽭��Ǧ�U�W����ޮX�i���{�A��z'���t�_���#�&����b�.����W��yzm��m>���{���� ���E�?{� g���|[�om�h�������/���Q���J+&�����$-W��옊��/�u~+��W+�����[�x�}W7��.k��w�_�徽-�\��z�O��/��ߊ����[_}�����*�]���=m���͹����^���ŗ�������w�O8;s�C�
#���#�Gן�.��\�-�x����o��h�~/��^-���������->u�"Z��zNy��!�}�/y���s���O��������a���ՙU�j�5;X�2~����>�>=~�$�����~��}�����������կKr��_Z��|�\ޛ����zU�u�sn�ǌ�ܴW�|���߭��=^����#O�#�=������˥㝾���������ѿ��_o�����~-����V�|k�m�{y𥳐>����y��_������^�|���ߪ����k׾��x�k�^���<���W�{οzU��ϫ�|	�>�#Փ�����.ͷ�������>�|8�#�>��pG���d[�y�ڼo���+�߿ޫ��F�+�������j���W-�\�ן|�׾��x�}_�y��_��r��/���#�@W�c��}�!�FrR��M��]�/�n��~���Z+�`����>�������6��ޛs�������[����[��-��}�_�u�o�{�����~7��������_W��~+�{�>�oJ�
��]/���a���_bu�߲u�˸����Q�<�y�����s^���+����o�~]��x��������o�no��5�~/��^7��o?|�-�\�m�|�����[���Ͼ����u�ow�>����zL�������
�1���.��>���wu�x�׿�=7��-�������ۼ���zޛ���_����-��k�z��W�Z/�믫z��+ƽ�{�^�ur��������گ����{���_l����'��\�Q�v�G��-�&mB�X�{w��D4�_ig](��B.9v�A����v���YLڵ�G��h�J��Wv��L=�
�:�%��P�0{��Zj jP���SN�fh�[$�Z��2�[�,݅�uaz�H>��\�����U{���ٚǼR���j-�߿}W���~u���z��mʼ�?~�xѽ6�z�z���ƽ5�ShG��C Y�!������"�����o�M�oM��+��ߞ�ކ����1 �Vs��f����k���η�^/���~�6����۽z����o�Kz_���/š�����}����������k��o�n[�}^M�noƽ���o��;o�x~o<�����~^u�^��}~s�D�[��nO��z�QT�����W�~z��|k������lE~��=_�i���뷦������^}~yk������~�_�h/��מ�ߪ�W��>���w�U�x�m�!��Ӳ��Օ+�FO����}�
��� ���z^���[��>��^~��~ߞ�����������:�7���o�����o��U�}���>�x�[w��>�W�}_Z�7z���Z7��_�;~/������ځ�z�ÿ��绅�>#�+����Ll�����}�v�*�������=v�m��U�{�<�6��sQ�+���6���[�~���~7�ܫ��~����F�͹���/��p��}�ޖ���.���H�\����q�D9��"+��⽮x��~����+�ߍ龫ƽ��x5��^��Z|�}W�����m������������[��_������������W�����;����[}^���6�Z�;/*q�yf��_���Q?|��?)�k����[��;o���~E�����z�~+��Z��{�׷��o��o���7Ƽ^5��~yޖ�b/.���W�O��}��$���x��u@�<	��{��B�;��y�z�7���A��&fc��=m���W����w_[x7�^��|�r���ǻ�������+���������?3���o�ݫ��sn����z�����`��|}�I�x﹯{���������}lDT����M��9�����翾��{Z7���z��\����wμ���k��?���V�wW,~���߾������oz�~v��Ž/���y��{�ݢ�\����W�����}��Gvcs�'�f!O�?|&>�s�ѣr����_�ƾ����U�~���~�yo_�k��_��Ͼ��}W������7�~����+���}yW������>��i�[�{����}m�K��_ȞWߤ�9*�;3���@�D,k��Ϋ2:�"�\x����be^c����i��;}��ϝ��NH�r�}�
/�U�J�˵ݘ䀯���h���^�奣0o1�# /S7��u��jp�L\�v����x�]��0��6A��9Mr5�+�W�W���閵@w��3���1�ɟ�P�� �}���u��-�W�]y��^��=��~m�~M��7����U�{o��_޷E������׵���u�_�Ͼ}[��L�����'�|8�|�[��]֖�w�=�*�d���y�c虙�阒"*a�zZz�����x��������o�;E��[ڼZ<�[w޷�x�׿~m��_ͼ�{����_/�������xۗޘ�8<��\����&b�B�����<��"�����4�&ϼ�v�ｍ����/{���ţ{m���������
�/G���%/8C�q|y�����o�_<���_��W���~k��V����ꌘ�%��1��n\oH�׋&$eO*{��Ϋ�g�� ���?z%z[x���}�^76�ʾ}���\����|�׵zo�ܯ��__�7+�����W�ƿ��wx5��W������}k��z_[ҿU�^6����߿��Ͽ�+��mr��^9��?9���S�b+�?��_���������Zu���>��k������������5���o�O����{W-�ߛ��+����\�������m�zo��$�{O��z��2yR��9�^�Ϋ��2��	��g艘�ψ�76���u�{����o�x�������M���ƽ����_�h6�|���W��W�O�~�Z�o�ռ|_��|׵�h�v�T���*���
 
��5�H[�o�����~���W����V�>�$�O���@��^���zo�n[�{��O�o���W�!�@�?}S���ng���ңĻ�0�b��0���`�Nmv�d5�[^3�vꊮW��n'f5�M��3__+LT�L�+���l�W�Z��O�y�@�P�͎�죘�#�����u�����0;��O�D��փs�IyB����_��Z�1��<mC���jD�IZ��r��=mj_mhoyY�b�6��E�z=��9oܰ�Dӂv頲/�Nn�mӝ�����P q��%=~�0�u;ᕃ-�`f�hn��0�i*z� n��f���'Ҹ���O*k,r���q���2B;ά��'.i;��0Gb���y �j�	=���^?�W�|��X�����78��pe�ȍ9yc�lE��c��vs *RbҒ��+y7;P�ٻ�f�j�(VB�U���%�93GR��9԰�f���0��(+�#�r�����w��	���3R�!W+���i:�C�~�lt���{��u::����G�rf[�xZ�U��S�6v��̅H�a!��o�g������?(�{Jv���ڑw�0�U���ι��}��G��(q�@��Vd���ʗ毶��j�X�5ِ�\�Uf�v��XH�"��� ��:L���8���+ۨ�FCێ�>/ua��ڤ����@�)��'���d���ˈlà�����˙���73H�B� �E��b����˶�=ۇ�+R\<���=����F���� �M��y/.��E�8BAd��6Qr݉���mJwԧ�&y�������-u��ϒw|#>}_:�)p��'D?��XPG��Ec,R13�"n���%I�G@�ݥ.Ƒ��=��68���ԇJ���PP��L���Ѩ�z�Y,����t����Qخ��qw�^(����2å��eW�V�.�Tx{ld5=Kh�<�U;�Z��%��z�gU��je4�n�t�&r��F��V�����Ȼ��G�d	�'�Y���T���B}�T����7��F�5L@?����r����%7��ez�]{����oj6Y��*�j��·kxC��3�6�Ś�9�z�ܦ6��~P�����ǎ	W[;g��-���bL̳��T㺆����ض�o��gT�h�O�'��+j�X
�m;����3���ڧ*����I����uC��ݶc��9j���ՊhʍQ�:�8.�dɀ:u�m��Es�6��2�Xs,<	��'n��tCU�g
��Fs�mn:!�	����������~7[v��S��?v�eN`s(h��;�66�{�������}S�"�'6�g�����_���BV�]�vGK��ס��xX^J>�)�dLL�-�o�h�\�8]S��)�T��d�Z��v0���݋JAG9mB��ja�qV�,BI�V�:��뢜W+�6��v!3��c3n�M/�UF8�8���=��	X�s�\�Pշ�ש�r7��k��X?-�?�L�0:Ɇ�@uV�E�s����-n�=u�Ky���S	c�|��{�f�?l�S��i똽]	� �t�T�˸���*���3G.ۀV�M�d�ۖ9n�bY\5��V'�g]#p��C�ݓ��+"��|��'b��/����� ��<���=U�M�vHo���}�}�D$��]���P��������D�6.w�F�}l�N��̰XM\ʄ�$���%��&�<0��RɛZ|�>)S���a�U�����p��]�v���N�M1�;_��F���F�/-.ٛ��SJ1bY4�pWJ�����]�pp��'�%wzFTU�˟��s7����. �[�c��z��b�������g� aκ�_H}n��M鎎yW=�[ˬ��Ĺ������ 8_� �ѡN�o�`�G1�+��}�O:Y|��k���Re��6/6����������`:�LQ`_0��ҡ��z��$:U���g��p��YD迍R`!�UW�\<�Ja��gۆ���՚>dFH��� F]`�[QR�,{�&Y�RZ-�K�ļ����r�ڧ2�A�0y�a�ϋ-��xFmvFTsQ�ﶬt�\����2�e؇��0`V
��+�P+	�h�Q�C�X�c{��3n)�h+���E*��C}����q�k�g�*i�]�������4��o�C�r��p�U��:nm:.j�6,#�}ǉn]�v�Gml�4X]ݍȪ�Vc:m$Q��,�-wA�J�l����ҧA��$q�t����O�崵�:@R�mu��%̙��k;)���y�DlIwU�u(��x������P-�P��]��W����᾵�M�����)�߱����w��tkNKbԖ�~�!�.cun��ij�eH�:��������U��cy���a�j"��o�`�u� {S�wU]m(�Y׮�ەDB�p�rޛ��ڸ7N{��C�ѐ�LƘ��>�|S��[���^����Y���+d%���xV��_f�`=��B��]���G{�U4�@�Cd����^�w�NHP�U�oT-}�b!P��g��s����t���[�8V���^�ld�m��؝W#Y�9�y��jW`�pY(Pj�50�v/#Ow"%�[j�Q��wQ6�'�f�6�}��P����=D�0��bԮ<S;jWa����;E��n�Pwe��Ǖ]�V2��݋o�FȌbe�Bt�uuUGJ�|�A^�P�':nFB�:J;V<�3!����Ԫ6L^����˙�eVF����yw=/*�`C��u�K<�X߻0ѓoɈ9<v}Uk>튲�.:��8dwRc8��|������1Χ��=LL��3=�ř7Ó͇{��㝠������%|�m��QKj���w��x�Q��F��mOqAS�܃�P�ӈ��b�7�K{���g�o�p��0�@�e[�KBU�y�����w���4)-Y�%�O9���34v�֬k�%׾�m-[J��}_}�}�yB��j۝����a��NVJ�XGƇK/8����C�d��1��j��jZ�ڭ�d�;O3�{�i� ��Z/�(�UpUB���q;2���������v�ʛ͂���>���~��w�jv]��n�K�S�����ŵ^��2��=9��]�87��vc�X��M�M�k��:�=.w*�ݦ�p� �'��3�o��Ic�2>ng=�ӱ�������>r���&Qs���t��p$��إ�Z�\��*0=B��i�B�,6��H�Υ��#G�t�o��ˀ(L��=]g:МmoS|��J X@�;�f�~���xߣ?Q�����ΧGk{������o�u�W�1�d���~.�������-LmW5[��t��L���6��km�ta`��P%�"^K�t� ?.�����P:��N�V��<��R2X��G`_U�{������_A��e]����� 6Pr�� [gfm㸢 1�Bt	ߩidMgZ��a����Q�R��ճ�,��
#���{�O)|�Y��w#%�h�+do�V�^��+�t癷��n�R
PT���e������o�i��w��v�W��e��e�Uxz�*oP;pby{�\�1����H*7�h�=���.}fR�wl��Zk��_}}�DW3��_9�xy>�w��I���:���>�\���!3H�B��H����;����W�jk��U�	�&ju�#w�p��}6���YI�E���8vL�G�	Ł+\Ȃ٧��:㤫)8+�kkl���'��]g{e�I2tB���b-ґ��[�׈d�u��ky����y� k�]̳��B��C�Q�d�ZB�i�
�Q����E<���W�{�͍>��]lTS>�so/Ӫ)�+���
�Cdc�AZ���V��U����Q��o޿D��~��x�s�C{\�B����fF=J�|B�`4~2c�OX�-�Ʃ�x��8���P�35|�ʔD6u�-�j�c�뭘�tЁR�Il�K�h���O��)�]��2�J�҉!�Qڧ*e����g�:�u����b���L�E}�_sr��$׉�l%�q��)�0M>���eȿ��a�N�!ۿ�!ci��<X�9����S'�
:]S�A�t
����?��k���������=^\'���to��'e�m�!�M��qL�IbL�5n���&,�ls3V�8�]��j<���z�&Sd��-kw�v6F��޽�tt�(p�Zݙ������E�����W�,W:���՚Q�n��r�u���N�pSVhn��q]��
2�-7 o�ڛYl}ev&ێf_�����g\�:���hu�������O3����&��y�j���t��K�Ⱦ<���Gnflt�wV���E�{�|HF�n��Wk(3���Au$6� H�,\�W-Յ����fE��0)�2�s���ذ1��&mp}Osx��L�V���t뛳s��k'YƁ�.<�����f�oT�苶��e�z�t���.�iPX�I�h�vL4sA��V��r����&(%��ܕ���ӻ]34�,\��mݞFΛ	2�,�����Y}��N��`��</j�r�[�l��9K}�j
x����2)�`;.dk��y���K]Dve�r�,�z�����i�2n��F�̤4���T�6>���t�ĝ�([%��@��RZe��/(���J��4�6��G*`-ۃįE�����Z}9��ק��-�"��WmqRL6�ɶ�m�-[�J��hf+�vy��t
��ݢtH"��^���!��*ie��+V��ڛ�Z�)�x���1-��;k�8Q*�\��&Mt�s�L/���gV�&1W��p#�n��1]��ǙV�۳�V���K���ޚ9$��:��k�^3�1��.�Z�nH�b
�`�p���D��b�ʾ��ū��#���+�����e,���4��~V��5�	E�_E�_f�]z��9�أa�h��b�ں��P�A��r-�K6� �%$^�f����X|cZ䱪c�qX�}++���}�mɠ^�5:]%Z%�|�%2�cn�.��a�At�x^t�(�vN͇8J�Z�V��L�z+E�nZ+�����!��RZ�����1��b�e����#9�^���D��v�,A6���E�8�SZJ���oC������W%����:�h,��Ð����i�\$�TgR��u��	��y%�x �m,�Thƭb6�p��gs*�V65o.��}@P�MjwJ5p02�Hk=u���]��˖gB�o���JP��|!v�����ffB�X+��>*N|�A�Hd�w;;M��Q�[8�N
�e͍`���	x�3�M�t���o������]`O�6j}�}5�Sh��W�R�4�d���%��B$0
y�1�%�Ol<�f�� 𦀭���f����e��6����p(�7!�Z W���Hu��#/;�Hw`�On=�o�:�ut�S���HOoU��9���F�ƶ��;b�2\v�U�z�M=p��lnU�Y�ԕ��UԬ=�p�8������m2��-.d�w����ch���2�(�"B`�&X
���B��I��f� 6�,$Tl�kd�V$�&ai��I��wk���:Z+��H4	�)�]����9�4V �F"�� F����60d��X�J  �TW6��]�2lQddCHRF�1�&L�2��H1���(�� 
4lR,fF�$�g7 �EPb4�!�nH�*K�D@A����&D�	�Er�D�TT�,���#i#E(h��0�,�#d�U��fҜ����*H��lA�"�-.�*Ch�O�ޞy�|�������q���݆��% �`�N@6cܼڰ����˶��B�γ[����avC�Ӛ�h�܆7���������y��0���:�묑�Iί@0F�\�Ȣ�@��!��q���zzz�1[�w4Tʡ1�����o����Ou�Bk����l��κ�>�j*�����M�'uWtCY�S�\��S������+/��g���"f����B�
�p��>s��m�̪id�bUc�`*C�Z�ݚ�x�'�N�:Ɇ��$_����'�UrD��^�pk-���Jˬx��\@�k��Vn�8���ޑϋ#�N���ul�������M�nr��웞w&�X�Hz���|R���qg�9hO���S�΄zG<&���`�x*��t���΃|�:"k�@��ҚXy,�O�Bq�2��(CeN��)�;�[ �M(q��Ѽ��/��.%+Ώ������dcrAwk���)/H�ŹI(�x^�Ϋ+dˉ㔦�%�-u,L�����w.��U�s��ok�Wf\3��z'���Q�}��.��S'�L����UI��Ƣ����}�7�ȱ�6c< ��ez�=�)��`���sS���46no^��3!�:h+�[���^���-�%	��tS�m|�;�ky'F3�^��mk�!�v�{9ձ��7h�Ks{^lS���\���n�^�W8-8�!�l�<�`i=�v��DK�S�ꯪ���t�#f���G�g	��@!�U|ц����3����LL唽�z|ҹ�x��+��f�<&��tO�+�p[\ǹa.e-��I�#-�y\P6t����wgF{a��H����+�v��G@�<%��:Y�q���`���s	�������A�\n�Î��;��m�T�O���*���\&F��]M��]��y�'NV��l�D��q�ޘ.�ԫ���~`vJ�O��U&�l�Dt ���D��Tk��ڵ�㫊z{'�>�lo�U����H�Υ���0;�k#%suNϵ =�7~������ɾ��wX*]z����ڂqj���pU{FD'S1�-���aNP�{�����IY����U��Y4M}I��ƊL)��S��t�}I�b&N��.b�r�[���x�iu�t�y�h�[~(?�#�S����"�jb�s�N�J�.�t����S��v���9��<�éfv��f ���R�b�R`�J���/q>��=^�{�j��u{W.�W7��q���r4x3yG�z��ښ+u����=�9�?v�s��"M乭R�H8��^�R�I��l�ꕖ�����@tr�zV���m�<��Z{����t>�q��a�W+.�˫n��n�cүS�,X瘝Ղ�E����}�}�����"X̡*c:��͢�y.�μ�?\�&`LW��T��)q�m�(�?U���5��^d)�q���\���h�8�˓���muUd�����dx�m���MO$��թxy���R�u.]f|�V���t������oH&�09�>��sa����K���E��q{��H�-Y�4��*ʜ����I���v!�6y��x������ݭR��`��zoP~�0������ճ\9V:|ճ�GG�ˌ�N�Ys�K�s fn;5���+ksuv�.>{��M�0�Qyk�Uƀ��U��i�8��Ms�Y�羅�9��z]oWm�w�|�z|%y�x��G�a�W��P�>�~`ٴ�Ш�R���[��N=
�~�l	�^�<��Fsxx�9�1�0�O��IZS�^�q��_uY��1`wύGP3y�]����ё��//�b/�Qr�wX V����y}X|��)t�ت@�fj[0�:�b�U�����[��K+�t�1Ӓ2��D�;q��ݶ���c.�f�����Y9<3Z��4��5�F�Tz�IR�2�yݿar<�;z�fn3>|s���O�Χ�I�z��ȭ	ӏ<�;:�t�AU���n�K��nFN�W���ڥ�W����b3J���*�M.0%���菾���S��1n�����\�L˜��OW1[!!�B�u��l�D6:rn#��HmQ�uv����v�ح�HД-��V!�m�kT`D�B�E���F���\�t���OL�99&%�U�vs�����.5��ĤWt�jA|�����D�?��i-��g�h�h�vp�wP��cVF�4����ۉ���V� 6Pq.nP��ٛ���%�蟒6��K*�:D&8t73���<5��X㜯�&)1�	tɳ�:s3��E��"U�W��{����.�x�y�Ȇ~��y"�z���_ͪ��c�8�ٙ���\S�R�a�ט���B���,w���U��V�>�_<�czk�wx�+�}�goXs��.�vh=�OX~� ��1]̳���yJ�j�y{k�7�~5A�W�ݥ@�s���,����$�t�e�S�O����xg����Ԯ��QUHl�u�+UT����ݡ�ן=> ����v�Y���N��9	�ګ��=0��ǩ]�*��>��������y~e�3{��K*t7�!�6�'�E�.h<a�X��n�p{��﫞uZ#��&�<�X��� �~���s&�WEi�
�[i^徺��ͱ�]Wi���|�F�2����+x�^��pk��9���˺��7e��iU���/{���W�G˟G��:#c$���3>�I�N@�c�)���}���S�n��Z�\l6l8����m��C�Hø�wdW��DmS�`0�<�0�a����Ln�Z,ϓk�s��s�zJ�w{
^#�0zb$���a,�do�T��0M:���\heȰ�Xx-:l#:�)�dƄ�]gK����8�$<\5Y�G4U�	��|+���?�n��:*a?��<>WM:R��(��K�9�\�w|��^y�痠�^.IaZL��͜Hn�bi�C�N�$5��^�i\p��`���]��Y�,���|��A�~���@�SP:E9���Z�fm���El6nJn?)1���\Sw6��3��i2���\�G�� 4,�z}ׯE$RR��X��3��!�7��������y2���&��92���+Q�z��5�z� qB�?���<�L��p�݉�L\N���>�E�u0��:���%!z�T�Z�}�}w ���A֚U��Z�<!�O}aOh��r�D�u�hD��j���=1_i{e�-6k:W�!�8V�ђ����G��E�z�)���ĺ�f��h�-&wZ�b���L���]�fRD�ִ�zn�s��{X�7D_���<�ưÇ��'�/6+Z����Q�Ư�6wD����d�sos����着����~l=}�b����*�BiV-K/] WJጛ�(� l����%f�T>78����װ�gL��\O7ωJ=����[��y�%!]�c��$U�fod>q���K�官�q����N�<���B�g���� �ѡO��۠`��׊��Oe�L�Bk�ʿe�ǝ�s)Ld���ؼ�V�$K�Um��՘����{&;�m�p�s�,`����U�B]*�G�*"ԁ�m��9�#���ɜCm�u�a��
�*^畮��w��+��ô�e�^�_k�o�ඹ�r���+�
u�]��[�0�����5��\R)�ַ^��)3ڠ�{f͊�^�Ep��XxJ
,�8����o��&>S��|�6<L����_��N�"{�r·��|���ޫ��w�+_	Y��T����w~��5��y��P�ޞ����n�s�qP�/�[��X;9>2�(�%�xB��;&�&&.+��f�.��	³�<�U�"���/s�b6񙕢���N�'�bA9��s��p3z^ֆ:y%�=3�ѥE W��1�r�cO�����jvV��d��G�;+-;�V�b7��w18d5��C��{�p��l=��&L��+��
��VE����òp�j��S�����AH�wQ)�s��Q�ų)����r�g}�UU}�z���8 �"��b�������'x"т�*��	B�N�cL[v'6E�#����%ʃE�y{\�l8W��R�#��.d��a]�¬p�/�^�Ȥ��hr=S�ugk�,l5/��cH��vDjgR[��P���(�c�*���}���K�]n�=��]��@���ˋ|wz)�=���_r�I�Ԯc:AyH@j�50�}�2=��� ����{IN�����_��4y.�ω������"F-J�GmW�ꈪ��}7�cTB��5`}u
v�v���m�Ch��L�����y�nl�/1�X-���F�ӡuը��{a�Y���>J�d���
㓻ы��eVF����yw18S�G������PV�}F/���t��k��9�0�_�v#c�<�a�C�77;h�s��~M���~�F�Lp��z����g��:<Mʽ|_�W���y:�T#w�Jי���Mj�ٹ��4�߭�3�v���{O�vQ��C��y]l������1�>��P�<��Q5roƠ�U0�L�ޱ
�s0��gw$&q�{L�em�Pb�dh����E�K]��sy��Y;]���������) �%Q&N��E��q����#S
��go�l+=��_�{���v�iWJOދ��Ni�~��lr5�`�u�c7h��|o(u�˼�]鸯�6�[�ץ�螠��̥�����`l	�u��sq^oG�Z��*.$��g.�?d�-�:/1��ؑ���P�� V��Y���#G�^\c�lC�Np��|��T�]����vլ��4�B��������þ�P�9TK�����Υ��4|�v���UV�iӜ]|W\�L ���� p���|T»�ҫ������x��	���&P�v3l����gwe�,���+�����Ĝ+��+�r��T��Nȫ��y�+�\U[�h��������{Jw=�_��!Z��{H:����i�!V<8�#�6쒋|NE�K7ЧvF'�&rLrj��l�"��7(��7����#䂼�go
�c&j]kȳ|��(.+�d_]&8�r����Le�$a�M�HjYs3�p�\ʪT*�q�ve<3��w�%+����a?z�����;�Å�CH���\.}_ͣ%e&� o���*7ukk��;Yq�FH>3+��΢
�G���}��7y����W{�Z7�ʇ��CF���}̠wl��'U'�Uӽ�/y~�Pv��S�tEn�)F��1I��՜�+���X9K�]k�6ԉ�K��ں�vU�}}���ɦђ�7��}�}��򄗓g;�w%�R@TY�[~�|Mv���'�څ����Y	;�TՒ�e��շ5>vt�y���x���A��U���U��PUc�z��Y5���������r��d���e��ߔ�EK����Y�t�a�2c��q��#�T�Ȇ:���qJ�\&�ĩ]sY�aH���2���shS�gɞb9�}t��'���+�	�����CՔUe�2�ebQ(���qT��%L�S{�h_�{�ϼ���=��T�X�hT�ϼ��;8):8Gy����x[��R*����O�����Fs�������Ln�qZ�;�RvaF=�+�^���t����>yiQ<9��t��5ʤߖ��2�\@s,<b�g�b+�9�]�=\B������k
:]?"�J¸<oc�۶��㕷��S@mQk�/s����J�Z�?��.s>e)���*؈����ƨ���Z�wY�xZ��V��y	6�jV�E[���L�R�9-]4!}��C��|��A�����r���;~4V�[�e ^Z�YN�e��ЧQJ#�39
JYjݛ�mL܋�{N�C��f\h�|�Q�ŻJ��5Äъ�s�e�*Ǚ���z��:�`�*�r��.Ss-=�w�,p`�<����:kz*^vNaڋ-�ƞ�3l1-#9S#i��{�»��3��y���D�2?t�Z���Sw2�>�&zxb&oa���UU���ո���)���� k���9p2��i����=�5��e!,\�b]��i�ٗ�m MV<~R�o�♸y6�D��e��&������ᓛ=I�����["�:�u��(�<�o�u��ؙ�����az��C
��o�v.U��6�73�5��/ک�&��"N���=�#m̾�
w����]	�X�,�u��.s
/A��ف�Ц{�9�u�3���˿�Zd��˪0�9�s�辨eZ��1� ��m�*.�5��!���VmӘ]�T䨜9Nn9�/����sr4"�Y����1���N�g/�����A�]�=C4¿����Ɍ��:��*D�UW��՘���e켤<*<�c�|�\�fq��d�2Q΃z��Bꎫ��S���Q|���Ja�6�t5t۵�۰�ž�w��S�Q�2P��R�k������8-�cܰ��xQ����xJ��t*/)����Wuo�մ�Xe�g�9���Rb�,��ї���|{W"��pG"�Ҝ=;B�D��h��%�+)Wn�ᎆ���cy!;q�&E��[)��;E��޹5�n���J��vl�@�s�ݙ|��ne-z�V��O�|�T�t�/� oo��b퇡4�[�[x��ʻ�rZ/4F�2E�u�����_J����fjH��4]=�N�U �1Sn��H�a�6
=̛��R<�� 9�1�@�G
e�������xg6Gp�3xem��M��2�c��#
鉕��u����`�������д��;�]��mB-�d+k�]mͧs�Wz�Ud
q�r��^(%t��bH_e�����VB��6�E��&F̗v@u�
�>���07�[f�s����@{z(�D��ݺǢ>�x�5���qմY3���Ӕ���l]��˻����b>v�]vQVY7��J��;2��EX*�T,$w5Үrz��JҨ�Ӄ��2�^�"�%����e�9ǹXc�t:�z�!���^�4�D��cHKi� ��fK��.�\ċp���s{��qp�ܥ�>�\8����f��8K���_�<�Q��ۭ�U֌��2�4�h}�N�ˈ�k[�$΃4�i�5����+2�L��Z�
s0u։��C��^����*�.ov�&��7�>�U�a�42���r�͢ypx�0AV7_;��j��w�u�{��N�\��Z�7[]H��)_ǚ����>7V���f�n՜��֢���d=c�����v�	��W7ϯ��.�Ռ��CB�9���Z��6��_}r�}�2'f!���J�U�[�tıvm����׆�O^��Ɛ��ڈ<�j\��^P=sC��(�q�Mڜ@h�3N9{�6Z�*#t�e1]�dw]K��U����01d�mݮ�xQ�U�3 �!CMe�Ct�9(U�ĕ	#}�͋���u���U����0t
B���8ʫ	[�ƭj.ݽ�9!���)GML���F3f�9�1$�Q�;��s*�.퉓-�ʖt҄�B���3ѓ�"����s��g�h�X\��-��Gl���9\����E����b�r���г�.�=�f$T���)���xҬΔc˨+�(�>��8����s&�I��6֍$�g{T�cA��T`Q�Z&�L��(#8��o�8��r��a��|�c@T��@�Vg7A�g]0�'�]:�'�DCKZ�M�ۛ����!���� ��E��{z�Y�k:Kt,�mN��;�v�0Ñ�哪<b���N�㎭N�w��������]���T��-�m������r�T��ҩ`��PA��9��t�w,�+%��@ܫZ�\�:vMx�j�;|���]�]4;P,X�si����m��^�]��Y��"]�u!G/26��$�y���'7��<��7�!/M���u�2�Ե]������U�2�ED����1��I��b2l��I��E���T��`�؄�`Lh�K%D@���[���$Z6R��r�Q�b1�U�\�	Qcn�X�62m%bH�D1r劊6(���I*H
�ƍ��6᱋X�$h��b���&�2I�������n]#j*��h�lh��K�ܶC[P  UZ��Ӌ�Y�ˬ������y!x0wPc&L��ܛ5%���(�\Ѿˬr��P.;�����Ĥ�Қ[�u4�7��}�W�T�N���W�� �����l��PV����]zm���>�Y�q�:ss8߸�O�N;-P�S�*��[�T���6;>vz_P�s�F�C�.����O#M]Z���Ϋ���l��g�v>f8�����â�1Ʀ�	ې7��i5g,�X�ص$��\۠���r+���&��s|!�)���1r^��$^��K����qK�E��n������g�j�TJv���l�%�R<��^��q�U���7��)ļ7L<��p�w��Aӂƶ��Oz��E�������[Di��2&�#���S�B�==�Rv��}h��t�ֱ#�P��"X�z�e+�'P3Y,T�UA*�,��'�Q��F�}*���5�s�\Q�͢�m��y�����y��̶�a��W��J��1ԀtO*��V�`w�	ߗ{|�"��µu��C�<�V��Kx�R�_���_O���X@y���9@������B�����=��*UP�+F}�P�j�n���6���˞�:s:!����ٰUmzC�ʮ�cCS/E��K�O��Rr�ƶ�jnN���19�6H�3�=OkFY+�7Q���[�/`T�(�K���5]M��Y��k�m���t3���F`ޑ�n5+�C��Ǟn�kh��]�uw(Vw5�tq�uH;,~�����3���g��H�p1*�l��.6��hjUXLV+����v�������+�(f)B��eceuf���Yq��1�B�NI���8�Ǹ���{�k'�ڐ�C���y�|�cWĘ�w�x�����
����5l�*�t�j���:<M��뻿u>��&^s��]R�Ow�uүn>W{MȦ�+~^[�v��Ss���8*�n^�Gh�\e�+w�fv_S5��9'M�%�ج���������F|lN�X_��ؖp���P�nc_�JM���Y��xM�M�l<.c�=.w"��]�jq�r�����js;zu�4�.��V�M���
BQ0�82�f�����p؋e;�.��-��oا�	:Ι�"�����ώ��oP�e��=ˌԋ���X|
��9��� �}�ic��	콕�ǲ���� xY<��®4RC녤����з�K�Û�(�n8c�l��b+��S���?a�P���� ���A�H��o�g�����g��(]L�;�k/�@GG��%]�dj�]�<R�����9�[t�3�Q3N��aw����10-�+�P4��b�pnQ� �8��d�S��I|��2qS:a!�&�F*oI��'%Hw�Vk�u�u���v����}�DGu�{8Zw��=z�����W��K��;��������&��LJ&R3ZsSw���d��5��:��`�F
{Ҍj��\L�MZ���L�5�vf�;���#��d8�+�F�	]����d}�$�.+8�/��r9_�O��I���:	��K.fvm��Ԯ7�$�N�"�{	�Zp�/w�7� X����MO1�g�BO��m�X ������sk���܍:��O����[D٨(�V������LxAΚ�??��O��̪�Q���VŚ��:�4���/5�S�Hv����J��tܩ�ӥ#'U��|X��Y��s�k_��lN�P�x4��l��Mй�m����!f����rd��X.4 7o����0z�߳Ƭ�������u�� �2�:�̘�F�!Lb���"ڣ;�)����S8�yN�2=�/W��Y��
,"�l8���d��U�.fv/���_q���5��s�^��tj��n(fH' ��,�Y�Ɍ޻��^� ��fD
�qj싃�иڧ*���K����qUT=�~i���Щ�]]-cfo^��
�)�D<��l�v��ys��JuϬі�;cv3��Y���ѮlU�V��@m4�sas��kz���Z/���4��;�dL؉t�Д������v���k�Ur:�j(Eu\�1��L:����R�u%s{��;�}_}��1��=�B�~�X���I5�t�5[*�l�j/���ak?+��=����,b�B��s�ݱ ��������CO
ӂ���pP>�����4�Mf�dt9X`��cmf�B�)���?[�eNK�C95p�[1�q��u�\�w|�T��++Ʊ�����n*�r5K1���R4�?�_i���/�z�g�"��+X����{�E��<z�M��U2�N�o!�J��Sw%��s;�F�*��u��-��0�]wT��{�ԺFq0 ��z�y�3��=ٯ��]��ɔ��s����#0�1Cv3�/���/r;��t�֠��6�␡��B@������Vn�=b�w�F}l��8h	��Ǚ���gU���6��.�u�rH>40��o�p��^��Du�)��J
�6��˺u�#�.���B�%<�&��N�	�Vz�T��z4q;�1}�CN�k��*�Z�S��c3χ�1�~��O�w�ٕ.e�t7Ndb��wU#��Ū�l���Ycꂘ��W/F�t�'M�����A	�m���Ժiu��&�A�5igqu
Q�^>1�+\�UY��?
��v�^�ۇ�"��/�l�z�b���	� �`�ތfm�NI��5M����:�u�A��f�T���aB�l͝����><2��}���;q-Zĥ�U���X�u�L.��s�WNv#�.ak�`�rd`Sq��ф��Yb�U�jr�q�z¹�7�,�H\1�c:��}ns�V6~����c�h��z���k���c�����">Z�к��c����>io�U���ձ˒�I�A�ꗽv���s~l=W^"��O`A��%��o��k��,'�v+X��~z7~�_�B�ְ��3��;�(�v�)�fe��^�x8
�>��Gv�G�^�%d����|��;M�=�]��eL&�l�p*�A��i�3P>�Kߖ���a;�O�I~�%��{c<]dDݏ��U������渨s��egWx��f�l��O����ng��|������}�hB?F��F��\���v:��y�d�,��%˴����4厽��9ks��Y8�P��<}*���BAZ�s�1[W��
��bE�/]�2H�"��:ǜ�G]��^�\��S�������
�s�<+�:�_[�k��s�\ϒ�g9+ٓ �C�v�]
x3C���Ծ����=�ǸS�����Ρ�Rj���[�o`�t�df!�j�Q
,L��o'wl�r���R�]�񥳔�YSq��L�Xą�;mU��Yu9�uu�mf7�6�ܣ���k����;�������ڻY�����l&1�FLM�+����=�����B�wژ�l�^�3�/)(��ʞ���GZ�ο��7קWv��@$'R�����=J�ű=B�9*�_���*A=p_`�3�²��.[�D�Q/�}�S�t�u�|fS���C4��P�n�I�x�Z6e�f1Z���ۨS�n�)���ϛFȸ�be�N�·���˨�[)�Xv]oov�[?}MY:���ꍨ6>;��n���%Q�z.alG'w�32ʦ�j�C���D<{{?mݓ.4,�s�\+@���P��:Q�\���'M�����(|~����B�]��u��[]�'�TЯ7�8s�&�?=Lu���~c���F�y|-X�ճ�<L�8,��<bD={��mأ2��vB��K�s�j�w����ӿ[XeW�\�i�n���*o&s<���xs,��`h�^>����{�<��1�;.�\�j�jM.h;�͝�57���rG�3=0�e944��K�����`M���Q��%���G�s�bvd�5�UX�K��N�����;8��넴!�`Ӽm��&�,��B.�:�wWa>�;�O���I����J۫1��t�G��9�)���B���8.gr|Z7���y6�|�4Q��Z�q��OT�Y���?'��E�зN�}UUU��'���ݳ?K��(o(Oc�p�5diZ�ofB��?9wl�B)#�n;6f,���g����_�G��@�iV�N:K�_K�
㬔!�+�9sSY��o��)�l7)_��މ�Y�D\��}����+���ǧ��t� < �+Nx�»�ҫ�����n�,�6�����z�ϲ��_�봆�s����{�����ȑ0�	�Fe�oz�$WCf���8B�c�����K��;���.1������u|A}�&�6��|�3NrW2�(��	p)��\�V�zp�&�7����IM�:a�J G(��SO��;�*$�����j��/��\�o��n1��W�x������a����������(�Y�{�LB筵T)�­y���ީ͌Ny�+�S]Oƪ����E��g�{ydK~[��i�r�@��t��O\�9x�f��\:Q��o7_�:�s,�߭.��K�_J\�Y]�ĺ�{���C��e�9�8��#�ǅ��qӡ{��v��dXJ��Pv�Xr��\/�V���Ia�E5e�ݽU��T�Q��(�y"��W�[�X;5%�����U��O���Us;�b�k�s��e*���
�->Qhu�7�DG�H�p���S�*O�y�ڷ����Ӫ����jx��.��O��0)�9;�nP�Q.���]������N�fyp]��5���2���>n��U�/\�sx����.�F�������[��
+�&/�I��f��K���M\)κ�7��ȝpví�x�H�:Y��j��\.��ܘ�܋�ս�K%j��t71m߫������_�9�5��gP�~�1�D����Y�	�ε�����л.o�'��ݶ8�3���ƚ�c��v�u�G�1<���]�c}-f8Yɧ�G�=\�zT�ח���b�����!�^Ԥ�Zƻ#\g��Z��������gJt΅�+��U�!�����:9��7�-}R�t"�9fIJn�gE����,�Rwk�6	����
L�Lh\�%o[Ӈ�J�޷�7��I��m���>��f�Q�q��*�eϯk��mW���Uyķ�*@�:/��U�
�( �nG��5k��g�>ݘ�e�j��o>��+�-oe�$	�]�6��<��Xd������<X3^Z6
�ov
Å�	ѹφu[P���;c��\�DNf���}�˷���+])���1�
BW�H�;"}F8��ȞL����N�'����/6�w����K��ۗq*�R��S�7�lT{<����zR��j�M�/��o�_��ӚM�>�VEF�&���M�2��Ϋ�8��_z��Kkug.8�f�,p���<&#^	�sʏ՜�/j�!CWȿ��y������Mj����^Ƚ���Kl����U��ȉ�X����k,�ԗ�a���V�O���� ��w3��d֎�j��u�wF8���9�zswőWX'�=�U�M��Wq�ճ��%���ޗ�W�H~���
z�UC�Xq籋���]���R\fL�A��K)���R~o����oUvf¾��la���
�F��K6݌r�|{.�����z����ܘ���\&�\3�l����v`��A���!ăӎx�D�b�L�Eh#^[�.�؃�qOR�j�|�͉\�/��N�j����B�n"L���l�[��̍܍��h�u	�f��B�p���}�y�;��Ǫ�7��mH�hSQ��<1n��	ڋO� f��b���V:�5�U�ߣ�V��x�'�3v���v�Kx7�Ἴp�4���L���}B5aYt�bu�O3,�����@P"W#��XQ�a��);��m�c���LTΘ�%gk�Z�E=�%�b1&]G|�W�9ߴ$�i�T��}��*�$��=�����r���u���)=���:B�	]�t�؀�ɍ	�ϥotV0��[qo/R��8h��;�z�K̔���銄%q���N����l�u�P�m#aB�s��i�{Ӝ���K�T��b�+�bG3zۉ�9�-=�B��n�YOj�7�|��|h��9w���U�&D�C�W5��uԕ�8;�B���������Vw˞��ѥ�&��e��*� �ݥO�CF�]ؗ�z-�DZ3s�mR�~�����;���+Ն��ٍ������P���-ڞ �����M���p�	��o�+��>V�K�2���ܼ�w�HԬ�,cv�^&�&0�s����4�_G�/��k��P�;x�S㖱�x6)��Guz��_uei�Z��S����h��9�Šq �#6�	�UǴ��I��6�Y[�.ƅ�P[���9�f���3iv���)�Z��<�����Ve����[ë;q�IϘ�{�ݹ(g/��c��Z���s��,����rm���*�+c��c {'Z���\�yYiG�Sݣ}m�v�S�]P��0Y�b�S1ؠR�j0��8Em�ݝ��u�Σ{���7j�;H�yr�J.ȷlu���Ɲ� �8�R�W!W���kyt����3b�X\,�\�À��u^U�R�.Ŏ)��7��L�C�����ܦWW����;Î]1$�O�̼��'�**���ԓ��z3t�����Dc�ć�m�a&h�
7w��istվSQ�A!Z�kd�/�R��1zE�۠[��FL�p�V��Xȱ�k�P���I��(�Zw$�x��i�R���;u}�4wZ�����|�ԙ<C��o/��3�r�YX�nL�n���ٺ&r�n����4�+��a!LHV���bjp�>����N�,�wF ƃ.����Wa�P�:�T��j���qm;�F���	�vm�=�	��[��R�_>�o�X��k����r�k�aN�R�e7�.Z)e*��%�J���`j���z�D��M�ů���Cy���`g���+n�S՝���KYi�s�7d���^�������a���v�ǯ��(�A����Wv��Y���x�חy�M�b�x��K�;�Y�ﱵf�C�PW��8.��7��1(����G�V
�BK�(���t��^%z���0�ҁݒ`��f�U���5�����
]X:�a|NEhIK�\�cl�̽��V���kmPV^�FE����),W�ዯ,䚗��@�C:������~/F����Z_'����c�[��7�H�j�2�U�n-�ئ.�V{���ג���V�@�)C��ۙo��iR�ͥ�A���b��4v�\�#rm����)��ڹ[p˽%�Z�N�Y\1t(nH�c`FZ�%e��{r��TM�|�lޏ�^p�`����n�X\�1#�YO-��iMܾ�̀����X�Kjr>hu����^^J�%��]u`�w��vT�X��eΊa͠���)�F�6��֖�
�|��7��+8]�Q}�z+S �*�Aa��8�2�oT�:�zJ����:�����Y��sP�w^Vm��;Z�+��<I��.V�Xҝv�����Y;9��ە��G������ŻVr���͌@�V�y�Q�Me#�xsr㱛�^NC�"o1�$�2(���꽢x����e��7�J�~]&Y
�gJ�����f�Y��ڂ�%<D��]{t�x��P�j��{V���j9�]���k��#X�$ɳ+Ә��Z1A�j���:X����t��5Ҏs�����˳d�[wv�j
�4&�w8�s�3T`�G8R`Ӻ�(M���]�be$[Er�Z6�B�h�J�v�Z��)�,U��4F�w�sr�X��k��sk��p��s�wr�v7(�3���Q�"�ܸ�'
�p������aT���۵�w-r��W"�u��Isz�����k]��kg��t������Ic_R=�,׵�餴��-tR2WZ���q��m��̤��/z��IQ����خ���O�Foﲩ���S��<A�֖��}iv�D��jƩ��z�=jm����-�j�79��L��ig��֕�� ����\��{&�*�d�Zb(8}q�E�Lu$��2�\#ۦ������unFW�����%u{�d��#Y�,шҡ-�K����M�v�:���5O��Q���y��VC���s;A(�W���J���U�o/6�vIv}&�˖L���>� &�k���1&{����@��餞}
�e�kb���"��e�H��H�o_BYj;
��
QS��>��}=�ВGE꼊�B���T�;Ѽ�������9c]��4ſZ��^�eT�L��Ě�h3e����:!K��9�����i\K�[�����ʯ/\G	V��e� ��1����%��NH�ʎ��s�Z�-��ɥ��.Ԧ�,%є��鍬��d��$dɱ4�D���B<ĦFr�}�Z��9�����:�S���]m�25=
%�D9�sh��s��9�e�ލT���v�w@�Ak�j�\n�H�s����`��W���/NS��@��V��\�en����}\;˙�keѢ=����gd|�<Wm^�f)���	���C���
��T�eul\��^@�|������Ã�ͣ�ή#yi��]��x1j�q��F�6����q���d�5�z�֙v�va�3y�U.��v�;���o$������v��tm��?7���f#\�}6���",�Щ���O���x3(�4��w{����j����.���1�s�QYy�V�_���Ò�U^��|��e|�V|q�*��'��Gv�of*�;��I�3|�K��<z��5ӕaŸ;��(���&.�n]�� ev-W����¼�������d�q#x�f��Z����iz�u`W�>�����ؓ�O3:[=��m�%L�u#Q�N�����᫑z$(��>|2ܚ[r���p�\&�[)��;�Gg�L쯟(��1�f�mn*7%uũŸR'um����@����+ی%���%��
�k�H�SEG�[��c����y�it�[m���{�o��@���X�i]�k�����z�WhAW���e>������s�]�o9��5�>n�#w�/Z����ݘz����j���b{��hƦ���e���iM=��hę�s=�!]��={������Orq��?2��I��X�f��1o�*Hv�ѩ�nF�=j+!6Ʋ]��?f�|����!���_Q��uī}�	�ȣ8:h��l�����>���7~��;��c���o9ojw��y:��@2q��f��{���̓��,�HJ���F��`w�L蓪���~���k=P��9VT���:m��.ܸF1R��D�q�G?c���^\�2��|cz6.R�N9-\��7Ə4�&�]���Bo��U�u���Yw^$�����r4�������8�f���6�t��b5�����)R}[[�F���y���9�if�����z~�8���*��w��UOx�L'����z��vu��=�ip>��r�~S����ǇW�R Z7Ʀb�%��Ao(���*s�S�`f�l�W6����e��{jΆ��h<he�6����P�����vW*ds�O[��Գ_P�v�ň;��6�չ*ѩY�=�D����ûCB��|����2�;o�cp^Ґ���y�6;d�Ȥ�1H{Y����eO��ZN�����Ҋ�#���=W���({א���5�[�3\eW58ή��w^�y�d�r7��t*[:j�za\ac�Qz��Q�sϛ��-��ߕ�}{c	R��j�6�F�O�2�h=mGC3��*<\5��\�-d���m�y��Gm�d�1�`Ύ�6+�V�gDͿ�lJW��t���U�o/7��i��٧l�R�퍫ʍ�o�^b3��j�u�.$�W)�P	|��IR�n�S�����5��c�Ic�uλcMg;�V�:s�[&{�}�	I��K�i޴_S{7�yLGT���k(C�v4���q�m���
BUG}�AȀ���j�cH�l�[�,��B�v]��9�ҿ�޵��$�&����aw?�^4��̮"���勺X�����M���Nr桭��]�W�C����U��t��Ƞa�m���^�ǓdB�5���Zij��㾼4��"0��s�+���k���3UX��w�f/&��_�Jv��KM�{�]l[qg;���9Z�j���z��O���Y)����*���=2v����\�P��S����/����\Nn�s�e���&a�c���4娖�ʸ?���m�yz�B��,�����z�≠�<��V-x�hшX�ӝ�
�b�fL�۴Ψ̹4����G��<��~r�N{�z�R�9VX#Ex�%�x˵��>���/e<&9س���]�b�Ꮻ���}֎s��+�kT����ˬ� �J5vj3�;F�}im�}���m��v���-�����ӗ�(�N�U&��=��kf�g��֖�)b�T�m-/�˒����A�����&.)&����ݵ{�b�9�2r�3̾�4��5����Hմ궔._he^��M�C��M�Et�mc	�Gr٥��Qp�m�0zgk�ʤr��4��	R?`k.;N�d���fw�n1Cz�n�=�l���;��3��)����h$�+!�.�P��.��ٷ&��n�6T�b�|�j�-� ��֫�=����О�x��b!���V�e�ĸ�8�D/�z�{i�kk�������KOi����Y�98���qK���t�+叩��`���%wo\4��;b��Z��ں��e������}݄�1�crM�4UK�kn1��o�����=_wϨ(���^�-1DK��s��䧖V5�U�/���9[[�/[s��F$ʮ�����X��6��*��b��;�dB؟oD҆ugD'�&"ۜ.�3]���D��ڔ���9o�V�^U�{GJ��[Ӈ�J�%���y4)��"�ͬx�,>D���;ٔc�X��Ì�#��]K��7�?>S�9s�Q�}F3�Ŭ.rQZ�ֺ���go�:�X�o��Y�<�>K7k}����!�O9?<Ni7�_k�5�z5W�ۑ%������iHct��q/�>OJ��gn�tm��1�1���s����<��UN\� ��7(P��<�[9����8�9Sۅ�9���gO�uS���WS�I>=�Z��rD$�*�\ns4ս�o3�i�*��d'�[Gw,r����	wFQ3Y�w~�kv�kN�m,Ws G���l��X4"*���<H[+���D�VW�W�X2K���U$GF��,AHΛx {(���;ҭm�U��]�����bL��+�r�b�*Z�8T����0����j5yp\D����_��g���0:�"W#WX~�	�d�ߣ�&�z��V���ࢻ�9�)z(��e��f�E�1�R��W�q��1Z���ݡt�,�P�8lj_^�ܖ���동��w�{c	S;Q�DH�cM:�AWi���׳��\���S}����p�Zm��)��;Q�c�L�,Eu��)s�1��Yv^��M�w�]��UdF��\5v��i��-�3ڐ�/�N=�k$�^gG#�d0`D���5�b2�/h�y5�vF��6�qd�1=쭞����X뉻q&r����)l���f|����Cސ�G	t�}2�⬶-�S"���9��BUw�T���n4.y�o�-�������E�_�uq�ɖ�p����I��C�2��i#;"}G�+�jbiL<,�oC걗��J+J�ا|�7�Իr�U�B�)��$s3׻ʡ@ה2"v��`Vo��I�k����YgL5ۀk]D�YzH�5��\�^�WEǼL�x^��h�:��0�u�+�]|�ӛ}�j�h�H�Gn�2�z���Vcwv� lp�{:<�w��Ն.r5 6�K�w�����p㻹ˡ�2�1�����9;��wq�/��{9��}�_|���Bn5ܬ��D�)�u7]'�����w�S��wC^fRy]���8�f�8u�ۉ����8c��HL���Z|.�v5|&c�w��uۨ�Z���ӏ�y�\:��-�T�Z4mC�ή\ӷ�s ��Z�3��.��鵃���{h��������9�̻��n?$��7'L�~+>�����x����4;��!eܛ�ڲ�X1Y��Rn]b����}�l��s�`+����-.*�.'8�/3\����BW���nw�76�{h��<p�ҥ�լGX��T�:�Л|�8$�������VKsвZ�M�u�: ee�<�w�ùc4M
�t9��5��������_�Ἰ�m=��:X��j��w�Ko����d˨�3Ҡ��~�I*U-���^k�����R�Yv��躚+�cr�\$�4}�:��G1�]��;S�������DT9�5��	���p��y�|C���S���e�k7���ѭp����wյ���N��[�h󺵟-7oW(��K�1�fn���<�	�����:�ɍYܮ;�dv;]8U%=}�ꀠD��Ƅ��;��P�r:nWmR�Y��S�T��ܻ}��f�np�B��]�u|��[:1T�������o�㗬����&�3�C��	���:aL�ɤ�k�Y1���`qwk6/�2��s��Sf����C}-K�*ዊEkY�����(d�'���8�zbz� v��]�����/���юi˹n1�:Y�lf	:��^���v��:/>n�U���r�4�-�x[�+���ѫՄ>�
�KY���jzn#)w���.z�<�ћ�Kio?E'k��rX�c)ak'����by���߫�
��8��;��̳Ғ�U��U�J�k�n]�ou.�x�.7����U4g�S����ȩ�i���C���-�1NG
y3O�N�K�<⺴�PNs9GAƚ7+�u��gv�ok�v0m��vn�U���x��F�
���+Sv(���[��Ў��W��<w�1@�o�|�q�;`u�ˁ�#���]g�[[��&����96�|�������D_ER��WO��c=��,��C�:���]8@�;���^��'ݻ$�;��;V�Xޑ���v����:n�0nT2�*��]+��ث��_P݃���h�q����Y��j1Y��BW����������X{vd��=S�J:�=�f��!mo��@�Q#��M:�P��R1�9 Fw,�����m�_#�U�%v�����=\�v�
K�cM$�l�F�(Cڭ��}Bޞ4W7��_c���|��H�I�߽����==uxb�pnD��y��c����w����vk��m�I�2���^@�;S{q���K��87����!�O��iC:�<�qmͽ�P�� ���G�m��~߷����cJ�+Q[Ӈ�J���Y��s��q2�l�Yt��<��
A�2����Ѫ�������u�����qﺢ��qU�-:̽�Ҝ�ԘT��HL����n�	��|��e<S
�Uj�A��P7�f�t�j��!b	ۼ�;C@n�:��n�λ��Sە��B%�P�zm�kB�L���ה+�S�7tl�qe`�����m��q�VC0=c+cgS{F�xh��hEW�wy'/����X��s�m.�I�1�����B��Z�
tj���rǶ�G�	p���yl�z;�����Dqu��w�%6ּ%���a�w_ �Q�W�*p��*�lN���N폠�H/�y�hB�Y�m�g\Ԣ�$=���{�=|�E�*:3�Uv�P�G,W����T�/�3��\�m
�IW�Wmo��tiF�:�����vv�2����)��H���{�?�ꜷ3	Y�s�;-�lR�S[@�V�G(�[Mf�Y��XU�)�E��yb�/�Q[��-�*D���=�N��{4:������wG[�qs�ܧ�Vk�Bw
YW���Q�߻FV�����uf�k2�I���I�+Ԅv�Z%��n�{6Z-�ҹ���h��^��z�ˁЙ��Y:��Tp0�oL�v��]�����m����c:��_+�|�ԅo'�jG����&�=��r��Ir��vO�5�*"s<z��J0���l^��~\�Z�+b�l���c+)LZ���ڢ�BeX4�C�����[.�uF�����eY����4e�?=����ڔn_[S1`�K�mW 5�*mud��oK�Û��7���
�q���������f�k�g�x!�[�}���z��!�P���`�ӘÊ��9�h5r�[���C�W�Ù�r��H������`�o�ȣ����q���.�c��R��r^zv\rCo)�U�.-����<�C��N�]|%���\A��n�LP啺��{��r�#|�^���[�"��ĝ]�t��_%�;_j��oMt���MYF+뜙���^���V�9�ڢ�����\�U�͵,d�X�Vk��ˣ���:*2��J�[�5���$l��ٖ��-�-;K^/mC:�ށ�ޛA8������ǐ���n<��Y�wr�9�U�˵:�D�c�O:C];#ozb���r��wx\��CzPCo�)9�����j����Ksw���qWi�����*��:�r���ͺ�q�e�o��Z�K���9B�7NK%:E_!��^���4r��=+0���V
�V`V�>��|�o3�i���P@��_ �#4���=�[�C��U���,�b��M8�ѕ��ٓ�I@�vD�m+���;z,e`c��Ѳ���ڕ���l��`�أ�������&���[:�j��b�q
�5NE>� SOJ���ÇZ�:XΤ�ۇ���j�tb�'Ք��Lc*3�������j+��\��V'W�"�LO���"7��ޮ��nTw��WQ���V�d%�+���l��pU�D��d�^��G����t8��!f�-Y���]���(�F��m���ff�����*�|� EPW�A�����gv�����;�5]6
6��͝�wtţ5��ܤ�݊�͹pӻ���ns��sb.�.s]�b��c��ܹ�naΫ�4D���9��w!5���5͓�ͣ��J[��r����\���s��[��s��:�\���rŋ�KEs�wwJ�;�5�]ܚ���ˤT]ݻ�b����ݨ�v&w[�.w(�ۚ�msk���wE�wwDU� P
�����j�	������u)Q���+63;���=��vZ��WA�n�&V����^�NrF����Y��}�c%�=��.F�'4��N"UTk"j9N��l2��H�X�yȵ�	E��������kRgmk�F-��?7���f5�P�quz�;�z�̖�_+sx�S�1�l��b��?N�3\�S����9�L�r�n�O7�&I,i�dw�*���g֗����VU)Րq�j���5Tk4w�j���z^e�z�yUN�:��Tz/����+��Y�,�ycUפ���w'�_���Ot��'������߇�k�hj��'vẩ�	N]�^���b�E���I��v�:��w�{c3���������̈́�s4�u��:�EwD������[���o�'� �Dv��T��_>ҏ��YO%���xK�X�/J�
(�GS{z��94��j�0��78����ji������]&#wZFYe��O-�k������+0��J��ûٵ9��k4D�l��))����q�L�T(n=��l|��7��������ޣqS�39�v[>��Y5����94����p��^X��e�V�L�۴�\9�q���m[�z��&[���%�u�ɕQ�.�
D��cG5�o��f�=�;9�d~�a�yY/��F��-9��:B��]�U���:<�7�I�"�@�a��w_we[�2]�N�����7�a�*��&�1; '�}o�-Se���v:������zp�˝M��ߏ�Ư�gݝs��ȱqq�R��&�[�n�U0���Y׵���9f�F9�4~Mƻ�Y��&��5"{FV�K�V(�﯎|:$io���|���0�4V8ta���u�:�r:�j�V"��&x�/>��GΉ�<�����y���#�=q�iD��������s��6������Y�ڴ�~��/��J'�ٚ1�K�jw�nP�����f�ʧ�i��\F���G4,��0�q�@��x��U���V�>�����
*-4�Rns�gW6�v�c9�0�
n���H���[V�s=��%�X)j�Z�i��eξ~�Ut
���GB�N|&]K˝ҡģ˨�]=�\���o8L�(��dw��T���z�oun��`S7I�:��bP��kM	9رrvv4U�M2ٔ��|ʷ�[g9ak���UIǥ����q�d�;ϛ����#ٶ����C
7g	�ͪY���[�h(-��s^5��Wt�>}*�r�Z�����/o�����{S�*���ܛ>���b=�7�cZ����Z�a��7z�ň��pie��ˉ}��6�㗻��g���PP%��	*U-����\.��7=MnP�j�������LE��?*J*z�;���''BHG��7�WzV���O�ｚ;��>��EC�Z�g��S�/�n�['vόNd�J����"V��pJ�޵�Ssn!�
e=�?Tĭ5��5�����Q�N'$�G���/zs�5l��J��.7�wN��c/]k{d�(��8#9F��]��j�y7�[{T�r�c%ࠨ����y[�fJ�����O[������%��'��0�� }J+K��$V���ߧ��5/e�ԕ�W�p4{oB�Y�{k��7Cj�B� .�ӵj[|T}C��l�K��v�⴬Չ�ׄi�^�W��'d��:	3��Zx�B���zX�mVu��Z�VNC[;���#��h��JU���)��[}��b�ԛ3���ӜumƵ&�^	��=�'/���+_> �m���a�IW<�ӷW�go�[���xLj�f5OW�k��)�uSu��<iڋXZ�e[�;n�7�;UO/��k5��9�s�gT�0iN^֣�u6"�[3�x<�S����P�9y�* �N�Rn]cޏ�;����t�R�vC�9w[j�z�?����v<��梲:��g�}S�b�&����&�B�B��zk��쮿e����\`+���Y��BW����]ΰ��^uo��%h�ȇ"�����������k�Q�
={圖������Z�+\F���yq���S�xɞ�3��P%�s;�xk����M�ܞZAX㬆��f��\5�1��~����ۙS�Nk6&w/R� �%������!��w��o�yc]��3m��c��HY	J�!���U���&B�i�}������k�aI�v�zw8P���r�!�7��S$C�yx���M��i����b�D��D-.Gh�']�h��wQl�\-����k�w��d��~��}G�e�Ky���e�Ӱ�c�KS<���t�e��ݧM��-��~s��~b{��.�r�����k��9i�* ΅K\���w�.K�b����9���{�+W9e��wm}����v��zE����,=.yb�c���D���W�v�����ɞ��)�V_>:]a��3�m���c�.)G)ڐ�q�r�qWט��ͺ�x����-�rZas�q�h��bsF!7��D�)ؾ��`�wX�A�`sǩЪ�t�en��է�V�;k\:?[Q:��k�u4�V�	[;�\�X5��c�k��Os�ټ���㿹Sۅ�9��gJ���;]X�j=�\�L�<�0��s��N\Fr�8ӵT�lgB2��ڭ���*�;�E.�̞~�����vu���_�nT;�!�kr�]���9�z����f��3����d,��C�Xq�u�o�ڋ	[�t�<��$�fv2з1v��U�6��ƕd�i��w���i�n�y�kk4���OJPa��e��2�w�lW]O=P!�U���tu-���q.=yd�`Tm���U5�}Ûy�N�ws�E����iq#�p������T[\��	_;!����+���s�7��}p�n���*gk�Φvg9P�]N�ӷx�X���:�s�ek*�7'�p�Zm���{��q�g:1���%��az�ѡ�α�.�l��rWX�ۍp�_��i���}��ܒ^�w�d���u�ݹ3��\�3�9=ݰі��hI�V֌j�7� ��u��|�B���N�Hɕ]��P~��Lh��Z�
Q�����~�@��ú��e�{"��ou�삣�J�BGzĜ���v̈���QH;q��7|m�nt�i��nn��l�_!+�D�Fvavee@�γT�]LpT���Ϣy3zp��E7��]�p�gʔ�)ڗ�r1����c�3i�FS������ev��o-?.r�7ƌG4�n5�D��u�"h���_>ÚW.8;�����[����K;�#|��n$�W,p���A:�b�^���y�;r�>�}v.�NN.�J���9D�0H^&��K#�+[!���_�r_q�w1��i���Ket�q:����@E�+.����N�d�4q��kd�C���w5�|�2K��yP^���\�V��E���C�	���p�z��Y3��[�E��~B�\Vy��)����ϻ��ո�U���G$�n4;�,��?Wd^�N�s>~ �˭eU���#o����Z����q�}��k[�<��v�T���G4/���;��	$���uUN[��{{�C^�%��O�UI�ϙ������Ⱦ�9�lt��&@�L�)K����agn���q�Ɏ|܆�r=��(���1���0�N2փLM�O3u#Y�N�F�	\he\`nLB�kobf��ܕћK+�i��TX;Q�aҙ܈	��93~{�L�x{��Xr��bkϓ5,����Ki��;�"L�Dr��Pb_-��⌴��.��������־6殩�5,���ko�p���©(����}A@����f�g�S2���]�,���:��C}�*�nD'�ۜ0�
�%w��x�'�*y�X�ҜI/��9&e%�h��o@r�ذS���t��V���D���^�|��4����Rβ���ǒ��FN0��y:��܏c��e����m��Ke'p���7��^�LC�̎_�cT�]���i#p�=�3T���p��VooYu#��ħhP*d%7;��ҷ����R�Z�y�a78]1����F�9�,��{����?OH�	���{��{�{˚�����R;r��3�$�l��[�r�1T��6%��ۨ]].����ϔ�����B|	���Zw(�,�����w*�"j9N�HZb]�[�xy�^���
���ܥW�L���#9�0�ã��w�N�Q�z�mi����<����z�1{�W������{oj��&vָtbٜ0��Y�=Q6�
�j���'C�6j��
t�峻��ҝ���sq��k3�2򣝋��ƃ�2p+)��*�G8k��b�	Jn�E[��rR��u����ˠ�K:��s}��m�v�d���bNa�������
d�؋䘺I�.%ow��s�v�9gm,�����t��K�F����if��T%�9�ϖFi���qt�������8$��n,Fc���w��]o��p���g�S��Ţ��l��;CR�����F;��ꈄ���F[��p�]*'�x6���5toOv^�J�=��r��pX�}�gs�|$��g��㱽R�͔��P��Rw5��g��|�ݶ0�S;_u#��uуj��?`N�.����ac�F���G�m����;�S��gh(��_^��bCz�fݥ(P�ѮM��kRyѮ�p���-�#&y͎QS�	k�(cW��H��8�����-:�>�oO�r�D�I���N��^J�����3��Uc�'-ęʎ�:)-����9֞��W��\�%�d���d�]ε^[5Jr���B���%�� s�?i\�"V����sm3��	]S��V�}4b񃛽���ܻRSyb�8Ą��]u.ʛM[�ܕ�k]f�8�^���p��M��n-�
��jBfz�q|,s�:��P�ƞ[W�����]�h�X���7�UW�Ț����{���Ωn�'���X�����.8�&v�k�F-��?7���W=Qw0@��[���2�*@�C�^�BЏ;�.�;(��櫸nN��UoA��V���g|q�T�v3[���\nS�A��%�A������_s�Y�������O_eX2�f��Y�zK����.g9���o	�%�2<t��΁��%�9v���m�{�,r�7j�m<�������8�9S��k�h��y��ݡ��陏n/6�����:���	�V�n=����N�^�?VQG��3�;ʓ6���P6���[4�Ϗ�;:��臷��+aw��߲����nm��6�G~��~�1���C��[�~[T�D��q=X��Pe�=xܾ#�n�s�C�p7<�x�v�\3۬����L蹶�q�X���5���Q&'����q)c�_hnM�ooS)���L�3X��N$�M
AɗP	|Κ�|H[�GS{q��p��f�
�7$�}`�lֽs��w�1���Q��_`�놌���?�J�ލ\�.x/
grk�8Ů�1
�2eTwϥA����q��z�~� ��%�֎e�9˷ۉ�Ɉ����2�;��s)l��Ν!F�2CbgG�1�Հ����K�����<YW�x�[�6��e�)Fmӥ�_!�ZڼW�m��5|y��{������!ے�]��3,؄0zֵ���ǉ��^��VL���w8�0˸M���q�xt�NP����U�vf��� r����$�t�v4�٦&鹪G���|.���w���҅�/��#�Z��R��[�/�|�v�����7Jֻ�7P7mD1^�u�K�ڱ@���3�E���:�x�*yb�Jb%��%��.�b�� m5|��6ne����sF>O#Z)M�Ȏ��+�2X��q�]��W��@Xו�[W.�Z���D�-��ƍ�َ�e ���8�� g��Z;E1FQ$i��rRކ�7�]��f�oVn�wb��(<����\Sټ�G��wu&���B�j+�d��W��e<���6B�\����fǱ�T'��˓,�Z"�Wf�:\uͅ�i���@]i��������s�����fڊ�R[$�d�� q���>����#2:��ҾЃ���dw�V6��J�&��V���rtf�w��IΎ�q�oVJ�?vk�p)���ћe��2��u�bS�v�v��N� ����k�����:u/L����] Id��8�7:�CNU�_^}p��rܫ.�Ҫ,Q+�ug$+������i�]�"7ַ&���n4��)o6.�:Xypf�◶�|]8W�-_8�!�%�)1}�
E�򞢖\�g��ۗ�ScJB�M͸��+�Z��.ʂ�5Pj-sf�gj��s6�Q��,eK��XB@(>y�O`[ܭ��փVy�!DV䖔+����.�����5�ˌ�v�N��\��3��չ��hL�j�'1�G+W\a\��P��W�6���}
�d���5	���:�ז%���hV3�WG�v����Wi�]���NÓ/8i���8���L�瘡�w_�!����nʴ{��pfQ >vA���J6\��=�9*v����*э�V��{��pQU�R�(���x�g�@'��r�3h�oE�V]�H��i��r���˩ǩh|�Ӹw�鹳1��6�����,k��Vb�.`�����3������@�lL����S�)w	*v�9��0s2��{M�^mg�"�����Ze.�lC>��s��� eYMX����'��VkY�1c�/b�E��fs�2��������4F��K��3�����YF�*��sxƻա�%NʩZ�j�6mh�-�j�
ud7����1Ճ�j�:�
�\�RV���S�}LZ��z�]�����UӜn�[ �3M�����|h�l�4�"�ߕN���A:�ǋ[�Y�*�P�J��Аެ�*<Ƿ�lۜ��x�t��\�y�Y�y���e]')!϶jd���(C�`.��l)@F����&V
oU>γ�X̵;�Ot�hk��K�)�]�ȕ�m[Muv�b[|NW=v����������S����[��t�wwGE�ۻ�j쫆N���6.nk���ƹk�LQ!�]ݹ�sF�rƮ�wk����sk��u�$l��b�r�wnj��]݉�W�(�;�����':1!,r�;��g;]ݱr.�\�nb�]+����wt�2���h0�'9�]
�3�h�wt��r�qwi�U�twj�].R�ݑ�;�(��wPD�����\�;Qnb��'wv�˕r7J��r�\፹�5����(�Ỻ�hݥ�ww.]"�n�Hs�"��K4Q�4~�������0g^X�4����軧M�Y�v���.���l{��9%���㦋V�w�B�q�a[�9�~�ŢR��W^Ut�����Ʋ��O�ɥ�i��1	���HJ�4�l�.��۵��������G�ͽ�Z��]����]��:�FQ�?t*q�y�C%@��r�����Y}�o-+���?sNi7�,���d�r�<�p���z��xݼ�1״��[�x�.xgw{qZ�7�
���&�osK�=5�慨�{<�i�ϟ�e�{iA�VN~�y:����\]/8:�r��u=��u�;�~�}Y�e���.����]z�S��S�W^��.���G
���ޔ��y��U7���慟��a��h{�@�J���2�o�t������i�*�ܺų���<��±3J�,y#�{yd�y)���.F����������ϛ���{h�n	訸�0KrE�蔰���b���H�tӣT%zW���!w�n��E����J�l��n����ˉݕ]ynb��W�jY��ʭ��f�l}җ\+��$zhN{ǲ�Ȁ���^	Wx��bJ�8�ýF�T����oYdX��3:Q 5u��uᨊ�H�9
�G)����d⾥',�F���U�C�DK$^��*�"g���w��Nx&<�'�f�7���}F^LP^��,���o/-0�{p�3��g�A�|��i$����1N*�U�o���]�6��<��o/�5��m���I3��>��j\v��4�D�K;�v(�r�
_��'oN��"��o��U�܄�4ŷ8~t�|��w�nb16߅e���5��e�����N�j�f���a4�%޵��$���d���,b��1v��l���ɸ���r"Se�Nr攷��Aj�CיͭR���s�{�c�%�j�Om[��]��j�y7�Xʽ;=ٜ�S��*��~�)<mK�_�KƯ�w�\�N�3.��2�=�s}�TJ�=���i�w�ñ�b޶Ѣ�ä�cRiF�\��=�хF)
�Q[��YCс�%��^�˻�(�Ӌ����g5��3��}x���_�[�����X�{�q�2/%vs�;�
?t���y�%�v��F�9-�t(3qx�}���(܋��i�m��D�Xz�|�����m�of������BD�:.��-9سL��i���K*pt+G^:���ҷ�ɳ�+���峷�����*���k��錼��4z/%�˲<��/P'���ih�����Q泍H���z}��q��}��mB/ϳ˞t���M�/ЕOZ[T8ק*QY^�:���2��LB�[��!����R�!����qxYw��`+��F�kiBVF6sv%˥��f*]��žks�m���o�v���*gg��#���˞lh"�z���V��q���U�����o��e=��ˆ�u�Z�DW���,�����}eq�5����hƤ���[x�i�|��Q�Ae�`����ӻz�9����@��В��]����/�5���S+���@����{T��I��3��wW�'�ɍ�dJ�?F'�-�ٲ�3Ԡg$�9�p]�G/y8]�&"Ӝ0銄%W|�l��=�W=ȕ����9^�Ѿd%��j��#�䆝���`-�,�c^���N��=���:�y�S��gL+T���ɰ��X/\�9��θir��n>�f����M�v�Yr,}Y���9�խ�yf*=+
�Y[�O3����V:�7���j��;(_^��9R\^$�[�w�I�y�\|v�u�0�g��HS�v ��L����y��'��\�M�����R�ԟ�M�
ނ����O3{y����B��@Mы:��7��\��ͣF!bsE7�%Uk"Lژ����#����^*Ǫԛ|f�D��������;*+�q�QM�N+&ƞ�8�u�'��H��}(�&T�v�}�/W���[\�+h�NA��w��.eR��m�G2��;K�-�=�Z\����S�������u9���W^וO8d7����e��ju��8קG��L��ޛ&���)���߾��>3��I�f�Lg����u���5��["�M���/�5L���J49�]���ny�K�������0��ya�(U����s�6��#x�F+TJ0��z�Ἷ�o��S�t�9#&��$mUZ��+���2����V�ȯ��A��eG=�qw�7��֋-)�{yѾI�K�赢`�c ����!+V!��^���:JL�蜰u������M�;qC6�`R0����rs����f�x0�.V�}���!鎮Y�����ڕY��R��%r�Oc��0�4u7�����%���m�d�͕�+nwm�)��W9�����r{��h�?2������.�+Ie�U;[*�7�X�dk���p�HɕQ�>���J[&4sY}��<+Y�f��b����n�O��[�O2z-���
�	U�|�K�g"�Y�[���xċ�ޅD)z1��7�-��M%�����?&�,)��Ou�G먑�[���B�r>Ώ۹ɗ�8ys��o��K�.�\sR�&�՘�˶�U.J�	ۨ]+��yi\��щ���?t����Rj���b�j�ZU�O�/'��u�4:$~[�x[��C���p��\���ŶѼ���㨦�t�-�~B߮*��jқ�HN~x�=hNya���wY���<����8�8U�����V�5��&���Ķ��2�����+���)sXk�J�adVoU�����f>����Ut��������oL�fZ������w�F���W�]B�iU��*��K0*����K)Ĭ_m���G��n�b���VGF���xf�r|�v���e�
�*�&�'w).����KEI����x���������v��Z�6���X��.$�3(j�|���v��r�s��7��GɩoǷ����+��z1���D��ӭ�
��|����}M�=�f�}�e�Ef��]m��p�%Oiu#k)::T%zW��y]]����o!6_V��������^��hkɐ�\�;���k�֯TXy�.�sCՉ��b�ׁ�����5�Onފ��3
:%�
�q^�MX)cn+��Ϭ��~��I��8kn1����F$�W|��+�bm�=����9�o�b
*��S�����_T�����{����.�+��:�^a��m��/�'e��LF��D�i���pJ�]��&2�B�C���i�u���LW	U�WӲ s�?i\�W�V�jb*u�Z� �WES�5�z��P�[��N�p��lݝ�^��y��Q�W��3x2}�P��v�x�)�͡/���y-���j����Ϯ��cJx���B}���/Fg�Ԯo26��{�ܡ9ac��n�=�9�[�D̮Zե�Qu��H&�ԕ��;
Z�'�Z={�5��2�j�OS?_?f�ޏ�w���Y�G^���e��\�G�ӗr�c�a	�龉�K������|����[�^b�|��x�%Əbt~MƵ;�����L^�t��k}�Lׄ�RpT�7��;��VZq\rgmk�F-�/����3�O7�z=٩<��z`4�	��o�[;q���,��k����Or���Q���=5����pg�ZW%]�+P�9q���8ӿ�SS�֐�]���w4��³Z@�K{�d膹��B��"Q;�-����u!��U�t.���rSl�?G>ݵ{W�0�R�%�{1�;��������C��]Z�L:�ԝ�Kr���=����Jgs����:�4������D��2`~��o�ٷ���}p�{5�g��mNm"��{�ڷ�2��ù0��IW��_2蔒�Wۏ��B�}ݮP��1u���x�(ɵ͠qo���ו�Qfo9G�f��^�����b�Km���q�j�!B��=Fu�<s_�ԗ�N�c�	ʳ�NP-�V+�+��;W��(���<��M5GE?o7��6�aO���6����5F�N�b�q7n$�t'���\hI-����JN��5�(Δ��[.ăn�Vնj�܋���S�����KKd��"/��ރ�Oq�kX��%=\Q��텿}����$�6�u#�������Լzz�C���9�
ww�c�z�9���M�z/�MF4�C������.E���ٛ�U�Tsia�&�Q����ME��ì�\�b�C���5�l��U��ܤ��6��.���N��\��T���<�M��B�L^�uJ�Ezn�F�gr�|*zz��đ^~�E�W�{�,î<�����ss�u[������W%�i��� c��97���9�\��W{.q�]����~i~�5u������������o����`(��ktB�V�Dd�wK�O��oӂ���W��rf����v.�F�܍�&����04�"�����L��a8\��d4R��rY"��xe[�s�۾uӨCt_�/���>f�0[�	Ӗ������4�묇b��X!;%����3s{P�8y�����D��]�^n�K�]S/��<�Ӽj�v��d�] �bV�dU���NK{2�e����V�2�-�Y�����n�Q����6�;�v5ns�}��_�/:�;1��vOz��\B�#F�U<z����O��t3�u��iQ��H4D�&�-U&��m�$�8tF$��5�o��]Q��ӓv��@��蚧>��>�]�-�}�^�[>>����zs�]{ò��v3�G^f^ A�/�Z�V?��7������Bz~��|f:��y�b�}�r�}^�7��9�?x.}+f��U�LZ�u�]�m�*�(�n��Tzgʜ�GY(��f�n����{���?7�������5�^ˏ$mL��{���3諨FM80P�gʢ��Ady��������r���nNW��E`����;>������o�ҁ�� ښ<��=<��I�\��M�?+c�۶7όs���{֐��<ᓪ3ޱ;~���T�
�(e���=�U��PTq�f8�Q#�}�}"�RCӺ�r���O�،ο1�3 ��\u��§O��#����g����]0�x��D�p�=h���ϯܬN�ɫ�ſyX����`v� ��(�����b��H/n0�b�e��Ը,h��Y��=um�a%��r���t�br�#��q��M���z�ȠؽG��pG��9am��3V�l�u�w��e]�;Z\��Il���^d�u��ɞ�e�+p��)�;�z_�?G�Ӯ<N��%_��i���]������z��}�I���>u6�7���N���@�u9��33�?]ԃ���D>z�|wF��4��٣�]�o�R��3<�9�#������</��77��Rʼ22_�P��,v9q�>݋�z���v'^�q�{q|�}�x�����a���'��f2��2��.V��g���/�Zs.��/�Q�=�`�=��:�ǝ
��^�ag���o�W�~C�V �'#��D�zO]f��5~���Ӧ]l��P��4��9���#ӌ����9{�;�հ�����)�2��/_w�s?�=u^�@nȃ�
z:�o�A�f|�������k���o*'v-��}�3Vp�9�C}�Ys�2T^��a��
�|+��>>"�ٙo���3��"�`�1PF��:wҸ��	��7NZ���>�ʳ�Wa�10���Eq�}t|A��P~>���,�yށ��v�����h�	��?�����>��Q�������%Q>~�)�h�ņ�1�ŝ��v�ǅ}5�vl���������{md��ҲYDkp:-$��$�k�N�l�=Y[�iN��H8�=����h1wf��A����ڀL��"�an�;gqa�ĺ�5pݨ�c&ĕ ���|�VmbD;��Lb�ڈeoe �;s�=��|�	�V���.-ܥe�}Xb��GF'K�n��똻5�����c[�I3!��&.6xo��9�O)o����o)���,CE�B�1�,ˁ�&���3�ۦ�.���I�nd<�+�ǥT7+:�����f�x'[�.D���u��J$F80���6e�	�ά�y�qo.��8Q�Ңs%�P���ki_`�d��	D�֦A���v<��ӭ��Nn���E��P��bV�}9WMm�s����;1.�������;6r�3{i��뉓Ol�u2��D^R/��f�% X�q��jRUX�#S���b�J��N�y0J�9��nv춀ts��.���Fc���oY���P�q�[�o7�SB�J�^	nS2��c��N���7	?t����oi	��9ڍɜ������,���
�±,� �V�ι�ݔ��u
�Ojw��x��єi�x�RccM+���8���9������u�ȾfV� N��3��)XJ�K� ���,^Ú;�{�GLD,������r���X��f�ز�ѣו��>S6gk�Jzq�,۴u0wJ:��q�Ԃ�9毪ƈz�W��*Ù��X[����(��U��f-��.����{V���}�Pݰ���\�GZ{�3Rƫ��n��q�S:��	�ko�"项�)b�S��&��%!ʸ��BA�����X��D����+N,U�q�)t$�b�����A�;:,�U!Y+���b��%�M�VW_E�s�0W^�U���q��^�{L�M\�����K���������������X�yolRq��	��t����.ĺ�{���4�R�`:0n+�h��0ڌ�)�	�4]Ɨ^D��W�����w��(��1�G��	��֮�Ǔ�CW�>�tB�˩��j��8y��������{a�]�Vnc��困���L¸��i���<�S����?dю�X=��kx͛�zC-1��P���Z�j�R���=��j�$�����G��1AD��7X7̤�e��*W	���xǹ�љQ�5Ō����5@sC=�{�cʻ�u�&��<�䥌�G��m����ha��E�E���A�x0Y���h�3��g���a����?.|{�����;�1ԹP'�����6��֝9co���yX���h�T�Ӡ�,��=�W.'\��4��kz�RJ�d�Ki��N��v���=�@�}`'-�*��]��f�;�s��S4�旋:�[4��6L�y��,�k�1�� �J�:Y���r������϶J:�J��f��v��2]t�/S��F�| �@#᜹����\�+��� ;��'uwGK��p��BN�c!F)I;��1�۹�b#IW8�Has�])�w\62wt��:�#$:\��Qnr.�6K�v��˻��)sn�ݻ�����]۔(�w:�L&�r�g\Q�n�WMw\L����ݹr��#%s�;��7u�v��I��*
锘a�h�
���w9���R��2���w:鑙��R2�A�9���h����r�.�	2�FN���u.]���ݺ��$�k���.˔)s]����IDęu�ܺ�s%�w..\���%4QF��)%��"�2�=�~�{�������Y*��t��p@�Q��%t�fX�%�Zi�b�{9X{�eaPʇ�!@\���y#�l�Xo�t��Y���B�~���)פ�C�Dz�b����>�F�����+�`���!
�y������̞��{[���_���!�p#��.��c�&��S�z��85}�����WwiAOߊ����F,y@�~0QA��7�^C2Ul���Z����nr���V����]{��`͍���`z;}p4Z,�9��!���;���a�{�''#� �@��:���X��z�g������X�Y2~e�QUN��D���j��/��as�[�Yz}G��1�ux�^g�=�O��g}�K92~d�Ԁِ�VO-ܑ=��`���������}�WSclkК�\{>���k��/����Cw=>ʡ�
�xhS6��S����x�ь��%��9�NVO�{FN���NGu=�nB~����z�t��X�����Q�S��w�S�]t�/��.�Ld	��t=ᓱ3�vw>������ۑ��2�O�׆�ԛ�ޭł�ō{���v)vơ���̅Wy�Y��Ԣ��5��9gO L���m��t��G}J�U,Z�ggW�{�ب�FzZԌ̬f.����l�ꛍ��swd� +�v.,����[�|�ꔶ��_,�fӬ������Ј�My��8p���sg1��0��; ���(��[��)ѥz_U���	Br���Q��]4�k��6��_>I?�c�T�<9?���]'=����̱P�O��i�t_ƫ��s�M3��Q]]������\��/�yS^ޡ�P�yy�Ǉ��VPۋ�����^������ޫ���/��#��J%��U�e�r����\{�g��g�gj�pI�I�?ێz�Wk���d�B�w�Q���j���Y���2.te���>�T�{?W�z�ǻ_TS���A�	�U��A�$?|+�5<����*�(��:�ro���ӑ��s���m���*h���񥖜�¯D+��	��
s5!/UM��M���c�>2����~.�Wh:o����d���A�������YF�7A���؁_y��3���ݖc��{3ٚ�<��
�b�x.���ߧ���j�⧀���"v�L
�UAQ�2���MR���w�g�Pv/�k+��_9f���Q�z)1�����=]>���.C��L�ޫ���"� ~�7�M��W�ob�۽Y>SC�}K��o����^��)����~��<��c���c&K�uU!ϼ�}g�wA�;0ok#��I��\NJ�m�r-��F��1�f�'fڭ�I��[+��u�n�[Ё!��bEE-U�zf�V���$�	v+k����a����2�v�Չ��olA8Ԡ���Wd�޲�ӯ���=��P6�l�5�1m���}Kf�i��)~)V���g���/��9��ת=�q$G4�#������^��Vw2��2���w���,���ر`z�*�97h������\5w��!�]��q����՚�/=٫���,׾�|J��Y��Sf���Z%�����I]l�����W�����;6WQ��g�}���w��,��.=�d��������0���S$����c|�kQ<큃ܩ��/|�ӌ��u[��g�vct����(e�r4m�S���w�[7s^�uਗ਼�n�]O�z�:,~�mR��ю�@\+��dCn�,��@ɬ�y��ϼ'مF�BF�����Jp��t����9���گL���H�^/�ӑ�xv;��Y_�}�^�5q�],,����5�X��嘑\�Y>"��2��>�y���&�����N���Ũ�2�:r)����{���Fs uD~ K�|��u���!f�n�\č�"t�4�v���M���k����Ѿ3/����(C4�X�b�@Lh'�bE��[{o<}�ŭA����J ���5�����Bmv9�m߼^�Z��G]LvK.u��&$��֐LR\1թ�L�W":��р+�6��+(5���j�B.:�.���U���Ҝ\�mt\�\9r���y,�0t�Q�V�L f���\����=a� Yo'r�!�x֜���1z��do���y�D�\��}�fjuH�垝�w�%�����3����&=��C�+�E{֐���p~:�ޱ;~��U!���;�T��U��rQ�H��$j�##E{���1\�������m��ο1���-���}e�A�V�iڿ-����FUuQ�:���
�*��zU9��9К�L\C���������ƻ��g\����`g�t�D��(�A��&��"kpA��yu�*���mz��EV�Ji�{3�r'ԍ�k3�K���~�Lɝ~��0;dC�~��0i����/>n���fq��1g�q�E�ϣ'o�����ȷ�3>7������UH�^�d�jf8����:`������f|�����A�y׷	?�C��[������ڬ���*�q���]yt�S�R:3���}9蜭�g�iS�4n����{������&�?��ޏ�;����t���/�+V�@o��x۳�:�e�^1S�[�y�d�g�o���\�Gc���������^���e�VJ*�>c�fY�b��~~�Wl�(�lNد*��4�i�4pN��!����0+E�.ot+�p�6��������(�c��Afl�\��]mr�F�ܵ��=Wc������HӤ����xػb�!�uu=\�`�hl�#�D��W����i�8�֋�<���xf���W��a�f|�"t�d����*s����$P�թ��O���㧐�YS�1�t��5������P�\a��$qu2��5>��Q��W^w���
��}�ޱ7�~�v���ĩ��5��a�����!T<"ć. �d�o�憚��j�T��"=
�Mx[�]������nDo�=�Y���OdU��@H9 h;����#=>�qQ^�i15�3��a��d�^��dx_���7�߸w��=�(o��+���a�x-P����v.�hD�� �\	��)L�	���r���x��O���S�����ީ���OH�5q���{t����F�:�� a@�H��QA��7T��u��O�T����v�5�y�E���^m�ާ�{�/�����TS�(0P�nKǈ��h{��k>��,��f]V^.��e17>�^�L�Ԁ�?:<���E�#��C�o��AL�)�Ƌ���Q=���{Y�v/ݡ^4ƟD/\?��ɍ��W��JG���g��rd�2y��,1��|��?F�+�.��w=Q�Ь�Kee�����v
�2�v֮t�7{/`bta�$�}RS#����0H;e�gA%���ee-B�r�����/�w��E�7�lg_���^�Py�\�N�--Uƥ<w�t��%I�V�3{,�w�����.ˊ9�*��E?I���:�!�	�uǳ�wd[�~ �����&z}�CטMN��F�/gT+q��pt���J�4�l��I]�𸆯nC~����|E��髶6��ٴs1��������`��� �NTyF���^ѳpS<gqs��r}<�}��4��O�z����]-Tdo��+�k�`n�@�^��!�>�pi�����̎����x� J:F_���/�{��O����x����dv�Nz��07lT<�P��:=�?xJ&�aJ1���{���D \̘����t�������T��a��Cv��۪xl���5��'��s3aB�.;����Dz'�/�����>�:~��\{�g�\wg��Rs�(l�/s���o\w�G��L�t���|j,�2\>�y�H�����~�x,���=�W-�TEǷ/G���9��~����?�yu��P���?���1p훓��ӳ��R�K���,*���l�X�zX�}ڮ`�b��AO�E9��$%��t�Y�����&zᛒ�anI1�ې)�k�:�*̺��5|)$�^=��&=���vQ��]�����[����ژ�o��$P�W��J��M�s:d\2ML�ҷv]�96�G6�'E'UҭP�6д����!�5r�d6P�[V3i��9�a�����,�X�V�Jj]�U׽
�7�|��x-��q�ht�M�`��"��q�K����ӳG����!��z3���*���r=X|�k�S�\g�D���4~uAҙ�n��N{UڣN����r=�o�ݖc���Lj~-�՜=��vE�z�f�W�FP
��>>��k�����A��e	��G�o�g�t�ʧ�{���m_�_����|=Y�=��ɔ�9�������L��]UI�
�KҎI��]�f��\*zz����#м�`�܅�X����rJ;��i�g<�s}:cuz� a�r���װA����϶����\�D�ȹ;r�����:3�7��3��j���2:׳f�㽦�����C�����t�y!������[����fϺn}om�}�����+"7ג8\{(�����.6�bFJ��E�=Sݱm�ޜ��nY�-p=���qgҙ'���/:�;1[q����VP����Ѧh��a���L{����^�����'E�\�C@q=�/+�dU/���dG���w�}��w��$��ł���|:�?t�@ف��zg2\.���]'u��?>��]�z�Mq��RG�Y�,j�]_)��;�o<`�塌.�k��>��HP�r
T0��.��{�K���>�ի	��w]ʐĞ.Ԩrw�b,:��u륯�]`�qݽ�������p�K���Z:V��t[^c���%��V��3���=#ƽ�o=u>S3������j�Y+�_�+�\V�����d'Ơ������,�2�ȉ���<}"G{.���C��H���Pֲ�|�z����>�| ��4�Ň3�C���}If�<n]V����w.���G�c�=����E{�s|f_?>Т��U��
 �
�_#��>R�oM{�V{%.�lo�]�/�w�7Mߴb�O�vF�̾�y;l�.�E��ʦgʬ��!�ȯI>6��[�E33�ˑq��}Fu�c��)�x.�::�ޱ;~��w��]��vo�{<���#����D�S���
~wX�B��*VS��#>ο1��ٝ��g%x+���FT7�e~�~�	a���"��h�"��L�ל��ݫ�i�V�ȩ���\H����nfVj�gg���`{%�ȓ�aS��B��v4���!���ȹ�����7�K�I&�8up.�q�3<%ϣ9ݙ�y��
���"zE��D2���,��b?Kd]��OߠX�����2cw����L��دt	p���! �e����U;�𙕔����*�h�W�K��+��~��@l�M�o�J��]��(��u+�ݖ�>�r���V#'Y)Vh���2X�+r3�VGxL2�J�{5�U�I�+`e��U������Н��m{�ӑ�3d[������cnn#���U�����l��/�lx�q�����~���v��Ca*|/��ۅ�'���g�Vo���{,Ρ����_���yϲy̜�nz���P��*�kg�;p���p~#:�ǳ�h�D/z��>�����9튺5��y�z+}�և�%n�Jy|��_�۳��Yk_�J�^�2w<�=9�%�= qݷ�״x��G�����ڍ�vG���Х��"�אsp�M��L���h>�3X��f:>�k��7�e���
�m�nF||}���x;=���`yt
����0��df��^�ٜy�/nB����ݔL�{����������a�����{>�=&!v�!�8m�`F�R���K��Cм��"���L>d�Q���3}S����\{ʯ���6�Q���	�����/؄;o7Ҏ�����fj'�þ�_�ӱn����ܛ���2;�>�F�����}���ld���2v����\}x2$���3)�S���T�+�6�}g�3���{֧g"�[A�%��Q���.P��FhN2����Nc���ph�%�)�P�]Ý�v�Ь!�t�7M�U΀�,��B(-��r{��G��e��̴ŷFk*��̉�1hAv�w��<��LǷ���5�3f��w�.`I� �vf��]�&V�vq���"�"�-�uG��1Emv"=,g�}p6�>�ʆ�N�/��Ǝ%�s��'�gݟZ� ʁ��Fݮ�͜���o}����>�ݥ�����|�a���-$�_�x�t�x�!���_{3˄f�vg����q>/o�ss�NO��8=��D��X��7���U�r*[���i�����,��yS��4�cO�\{����ۆ���~�R=����C���d�aS�Sp�yt��^.��N��w5�3���<�51�7����\{�d���? E���3��2�WVO �cݪϳ��/n�z�u8:{b%VK�KF��I��/��W���>��!�-Ǥ�ݞ���B�Q�?�b~�B�5P~c5���5o]��k�6m[<gqs�λ���ƹ���U5��\0i�K36�{��N��x܎�9$Ƿ�J|-rWr�ߠ��9��zE�g�%���l�F{^�6�z�g��[��>�b���y��gmt��a��T�ݑ�@�0��o��6�>8����v���Y�d�o�R�~��1�����]oC��h��/�c��+|a-�����������k+�
�Tb�PNK5�Ac5樛��񇌊�n�;b�,�tᚻ�]�4���je�f�]��e��Ά��a[NgZ�2�ȩǙc��m�/��5ֳ��D����&�����{q�yN��[��gG|�A9e��ce�y��9"��X�
�S��L��ܗ�r&�к�G,qz�=,PX4�z�q�o�j��^kt�\v4�<,*��R��-�a�S�L7BA��9^
�]�A�юː��+-��AN��PWn��r]e6I=���1��|w��1ҋ��d��buR��@Ӱ'����6�� b�u,���[�RU�;���dc� �4�(�vp���.m@���`�n��Aq�{*�e��Nqފ�',a�����w��{BR�������*��B`��A>��˭̈����ka5H��pVs�Ň����÷~`&�Q�Je r��uPh�{\U������i�[��䙷�W:=y�a�ZDW�zʧ�*�u�K�g:��:�\�����̮��umofL�b¸�{fT]���s�7�e!�M��V_*�%9����ʳUވd:��v�Oj��M�w8���;tĢe��wC[�uҳ7@��&,�;���[Q𗎅8Kפ��Jı1̡t��t�1��l�݈R�WN����g,i��u}�� _j�3sf��[΅��6��0KE���Ǜ ��t�'WweK�����yI,���{���U�u!�%�V�v|� n�fs@�g�e�X��=���&�- ���&8uIU�Ѷ�kk+�������M5;��u���‷ݢ.pd�`zBa,ג�RWf�u�HE�ؔ��q9��ŗt=� G�g]��u�-�r�oN���������ش�R��[`�ҕ�}d��;Bå�P��G�b;��wv8X����R�WP隞���q0hڸ�s���w�Q��Y�s ^;�@�6u����T�:p2KE���������fH��`�gk/
ek+��
�T؜��k�Xm�|(�\ʽ�`�{�����Zyc�V�ϯ�r�d��]�:y�C��<�Os{�ڧ6���vS1�8$.�w+���1Q�b�bz����opý7y�l��9�osy�b�<R�!���&��ik-E{���ϫ-'bo�v�@����Wv$�U0�ݽ���ۍ�;���d��:��]W��:1��;��니֮*�s+z���sU_�5�l�⿳�]B�S���\2�:1#�)���u.��10gk��9��0��Sx������X�r����{oY�gmJ���"��^*�\��VؾO^��]vЮ4�^�
c���,q�9p�4v��W�7�y��:����[E3��A>��˘<�3�kX��(jyr�L��K[�M���$Cν�d�/Z3�wVn�����-��g1%8�c�i��3�o�ψ$EQ4M  %���a�mȩ$�#����D�s���Yw]�2DDӝ�� ANtX)!C�(�����L�\�Jd�И���",F�f$LR)��0%wv)+�a��Df�L�(�$��+��'n�$�2a&�6B"c]܆)���D1���7w#�H$��M$�S$Ѧ�D#�Q��RJ1M
4%Αr�sq��9���D%����gv�e�1�dhD0�� �S"���B���n��f��JG7I9�G6��9HȘ��$9ӻ�́�Y&�#&ic.u�`�����\�`��&�&Di �$ ���$�� ��)�k6�w�Ӹ	�#�ZGϱ�s�LcYmu���^:=��D[-֢�2ŷزa���s4�ٷ0�c�u"��3���٢�d?�~�"����Kc������&���a�ޏZ���e�y�B�K��(�9/h4��й�E� <~�S�5]>�U�Q�y��z���H���h~��g�zgyz5e�����짷ރ�l;x_��8��3R<��4��WuL8v�ɿ���=,G��ScN=U�2\[y��%��+�.2�_��=�*�!��t0��
C��K�S�T۬�v`z�֤Ge���t�1x�S��&}���}�i�~����R0tC,ø����	��1�s-�����G=w�Yק�H��F�lnzY�b�_��_��,S��>C���@�z��K�.�:0�̷T����Ǡ׮0�f8�q#�}E�H�	b�c���)1���'��6=����o޽��>z
^�#�΅����Mkހ��G���p	�^*M�-�ؕO��=�Lm���-���������y��2������=s>���UJ�:�UG��9!��3�l�9����yD2a��z�}���[��Y�F�Q:�T_���(08�T>����S[{9l������4l����q�8/EM�EQ��U%�Z en\쓹�\vde��՘��^n��T��xK�7%ǜ9$�f�L�)3�w�}�����+��v��荬��
u�V%����Q��ܾ�ƵZ�b�� 7SFP�9TԝFŽ�ٮbRlg^N��Np�)�n��ʲ���ѽ�7������#�{6nn;�4�_��T-W�|a����7��;0ܿ{]e�GRt��_���E�����S��}�>o�����3޺���`lNJ��{�C"����W�3��~���\�h3U{��η~�d�k���γ��V����e�>^V:8�Ϧb��k���}?AMg���@\��>���)w%�i���c�/��dz�X�y�%���[��+��87��'������^�����W� ��g�:h:�:�=3�G��.!x�HI�{�踳�ے�g��J���U�W�[�쮊�+%�V%r_l���+Ɉ��r���Q�x�O>{ʦ�rR��}"}�S��{Üzʟv
�Wa��l@�~"���G��}�d"=����^��}ֲ�;��g#}���}?[�pȫ��1 DT8���?����⻫=�P"�?z�c�Ɂ�~�t��B�:���̾�D��%˹����T�hv~Y������� )~F�C?>i���!��2�\�z�g���::�ޱ:�0��;���o�ly�d�R�b�g3�6��t�1�rz��5�yj�Ж���u�R��������a��ʜz*]�Z�+��N_k��T����w�\�our�-���ּ��ؗ\۾�������i֘�8ގ��-�"�hu����>��O��_�����D�ߩ�!����r5}]<����=�m���5f�7��{5~�Y���o�\"X�`�hCj'������¶W�l����ܬN��շ/��V��o��:�y��D1��`<�ȓ�~T���k�A���\e�]G-yד��s��X�5�~D��)�|�ؕ>�$�|�π�xW�w�.�f_���,���G�a�J�
�.��,����y��wL=��>�y�"�{�3�o��stgc���!��>���+8�W��<��v&����pv���jT�g0�����3>*�7�`u�{ۗ#KyH�_9������X�ܪ~����W;[>��Ө��4w���.3�\{����+��o�u��`rG�]�z�V�u�7}}���c��X.�������4l��XF�_��T�V�G��w/L���^��/^fV�H�GY�C������5��`n�¡��&����zo�fg��ty���\!�x�+��_;LT���# �|��Li�]+VT;S�\��)��V1�G~�{X�_�No�P#e+�|�7 �y��Z&�B�����[B�+�!��X�]����)][�v#�� y�{��2�5{Pn�$/��2�
��ۃ���u�,]�;n�toxZ�1G�S]�(����]r���7���|��YkW0#�ǳ������ȏ�љo>�빇��ޱ6���]������ڟO];����0R�7��gY$����׮Ǿ�Zc���#�����<�������ۛ�yVG��OeY�J�Zfm.�y�	v�2��묐���ϑ�_�d�^��vG�ǯ���sw��z�����T�ܻ#�w��=�W�po�*�+��r<(-Hs7*��t�×���޿&��S����������ge����Y�&=�5S���~�~%�w7A�
�G��&��}Bo�^u�Fʏo�#:��s֙Ujrٛ�W7~�Ο�w��-����|�a���(���
���nj�@$�����	��c��O�w���;6����z�q��`[����z�qG�U�q"������6��;ݏ��T*�$s�G����9\{���ɍ��W�-��H�O��g}�K92a��W�1��ժ����h2���$�.;&�1�29S�״Ǘ��ȸ�����3�𹨽\ｴz���Fϔ�4n��T`e9��d�4�l�|}'v��^�6�N����N�7�C��[y��sW�{b`R��	Lz����*f)��A��;�M�j,�Djc��ZW] �5�֓O*���4[�C��R�]����m
��`)�N[�{c5
U/, �S��M�G3���nd��<�ʙù:�۳��z��=�u9/^���
��<19P�Ν�C�2v��vDw>2�̗�2�"����;��'��}���=ީ�R}�r;j�����ݑ�5�!����jÊ���=��<0%x�=~r3�������O���~+�����mt����L��{^Y�3!�2��&5N�މFO�x�x\A�~dh.fLbo�S�;��PϽf5�b�*VB��c:���������Ǉ�b��'Y���Hڅ�]�}t�|�GUz]Əp�?vǲ�����sUW��nr�Y[Q��X鯌����<9fj�]�Y>5��d:��7/���
3�|=���7L�O/o���a�荾��4��W��u�^��>���,�L[�nOl�H�~���3jEoC��\�\x�w#|e��~w�W��� a/�[	�,��fF7�����J���j��s����_���zL����!ގ���#2�;����߅C������!���9��}
��Ъ���F���b�^��8=��s�l�
3�"v�Ĺ��:cΧ�	��D9��5<���f�F������|ؠT���F[���o?;K }��K+Y��.�k�RQ�|���,�5X)�R�����vR��a���r�ֻ�^��Ս6�+oy}P�̻��&�u���]]|l��۪P�6�ѩ�	Y�/����Y�-�u"��>��U8���\����K1�\>Rcm?[b|/��'�Y!6rd@y��)�u�q�)�M�\�Y�������4�햇Ol�~�&6�~�C�y�>��ҙ�@+�i/ؙ���_����W{0�UI��0*�z�Q�w�����\r/��׈��}N:�k8֌��Qќw��g����A���=�c�^�@A�тlM{kog#m�p=��3=*d?�ϋ͟t�a9;-2L��ύ_�^�;;���}���^���j��,�]+��'��g��U�?�}�3��?uא��.v^u�����������F��G�Q���M��U��.ۣ>���⇳�=��4ì�!�j���5S��,�]U{Ru�4j+=�{-O��spTg��էp��N��>*��o�P;=1Q�-�-SM���=����3�Z�m�HXhx����?���׫o�<�]���N���x[�����>�ӆ��:ͪ��������х���^���{ ��gg��ǍH�ڵ
�n��W%��|h��CBw�������Sh,wU�����ՙ�-�&n�} S�t�u�B��a�N��3��u��I��ڒط}g#����(,"�}j�w0�aC;�,�ܫ��Ν�W��@��3m.�v3JťP�⚈sy�tm�͎�}��V��s�W:�"���"��&�hۜ��ᾍ>�7�z<\�C������>�| �.�H`���E��癘Oq|�;=����v��W��.a����Ѿ�����̾�~�>�W]*�� ~A���Cv�g����.+�b|1|i��������)���^����|.3ȉ�T�ព�)�ѥ���5�� �37�'�}/��.8Sa�>7<�;�7^��%��Z?T��<� a?ov���d����<)�@�u�GR��K�z�����_��R�)��B6m%�q�b����s�E��?L��5�ߍk��I�T��j��&�/*3p����.�>�_lp�G�|��a��ʲ�&���>�������T\K�QK�L?MT/\�`���E�QF��C�l���A����'�}�\�ɑ>��+�6�π��zg<����H���v�Þ��B����Z��n=J�U8�?�H�+��p�k�~���fȷ�3>7���g���77��R=����!Ȟ��m��W��6Z6�z�;��{��(J���ۄ��Пx�����::�n�#�ެ̟�w(2BF(��&2,��y�3��-֫6�6��دy]�	O��c�@Ӂ�.f���݁�p�����:�t�wƏQ�4�n��#��v20�>�
Ä�/=Xek�;� �fq��gg��j^Mx�G��Y�YV��Ǣ��㒤�S0 o�$	c{��n�9��v�-S�����_ӵ��N�+/����/��Wϙ��j&'�o�5G{:�=�������\~9��������W��h�{���4��7"53^�ܗ����0�yw_Q���t�yӥt;՟}�I̬��+�nՍ\�ܦ@�v�v��jC�F�q��W�������\���~9���>>��iNh������v�ҹ/�SJ�0��i�7����q�qD��~3>y��s>��X��t���a��dz�O��"����ju�}0�����]�����=Ap?
f�]qt�|Ɇ�x�FF���ۑ����g��O+��9��@9v��){�Qc����E��� 1T�jZ0�:�n�;n����;�߸dw�|�{!��w�s��5i�zX�Gj�]���r.B@��?
s5�xU�×Ʒ�z�T���1%�ѹ>{{�(׵���>�=����N�����x�!��t?()��&��}Bn:�y��&��"LZ4{��|�����\��)�ۜ�{:�=��{���z�h���Q�D�Ax��yVp������Q�j���͵�}[���"��,�&�Kh��j�kF�'+��5��l�#�K�����?d6��Q��[�{x¼���Z��)���e�8���]�W���,v�ن뿡���³5z\�tگ_v[�)o��ଘ^��Yٕeՠ9��Ie�����0~d~������1��|�N��~v�}�@yϫ%�q�x�ϯ�+]W����3�x�Q��	'efm ���=(H�^#!]zv�7���������#����c&W�ÉC����󹛀�?�+�E��:)o��U���xu���>{�=��oi�'�t��)��s�o�^L�۷Yޙ���3���G��)�G���4�l��������4p��ܦܯu�i�ɜ�發�v�%�,���9{׶.8{E`���j�t컈5�7
��;:�fV�wu4`�u+��Nz������#"x��=��q�$���X�s��*�Mf�kC���]�b��TQ�R�F}�=�R75_�gq��L�_1O��	������3�jr�SwpeG")��Y����>>��%T?'E��^f��1��T��Cƣסy�+>Xz_���R��^`����p7�����-
�*ד�fS��=7��Lc��jJ��H��r�����s�C����Z��v�`mfu���t�5^5y����7/#���:��W�f/����:z��'�6�ƽ� =�}Y-�썌�á�3�<b�����胙�7ak�}8���!�FyU�/B���f]-�Zn�~���=���Y��X��^�B��iKSr�$���Ý�0��F��)���])�ŽP��B$�	2�r����L`}���[��Ǽ�����Rs����G$V_��5#�9����d,�Lz�41��x:�����m�(���F/_����9��CSF�U�C�����< G�Nf�%꩞p�ь̜�u���VJ�_��z5ـ��~Γ7M��r<�����:��*F�e�wt(LO���щ�~e�X��Mz��`h	d:�����qW^��3�!��Oq���%�x��P���hߍlTt=��;g�X��I�q�}T��_]�f9�|���~��DVp���+$]z3��Z2f3������9�W��W�FP	����$?WIj�C���T�=�j3����}�sD�'��x��9/s�@��92�uU9�FT/\J9&�w��.���Ⱦ�^*���W�%��3�]�$��{���z��ϥ�����g*\M{�koe#��g��g]�:PWz��3���s����������#�{6no���� �NT>>�*A�ClW���{���h��>�p���+���>������3�Vo�$p��Q��{Nl|o}��̬~ޒ�Α;S�ľ���w��o<� j�� �]���Zjo*i�ɗ����s�1*��J[�(�Q�� �&�������!��;�}۵�:^5��+kDy�.�����+d�������Z�0/Ww#}s���h��	e��`hxOKV�=��M˵@�!ƥ��n�Jxi��[�J7D��^h��qâ�Ǭ���e.�:7g�����
SZRJ0�[AP�i����`�%8A������b1�1���gXNQ�+Ot�5,5����#�X�� s�n�e�K\B��WS�&�ㆶJ�:Ӂ�R�@^Dmje��b�1�V��]]޾������G[toh�*�a�=�#>�x��s���T�YQk�[i�YW) M=3F�C���n*f��C�!�K ����Y:�8aӦ�g[�1t�O)����hNw���.l�,i���S�+��4��s'Wu`}F�Jí>n�G���Ky	@%�j��v_k��:�rD��8/�ȫ�9iV�u���I�UgL��iɷ��V�=sS&���8���׍[
�m��J`�ዣ���J�WkB��.�!�D	k�n�
�˗_��Uw�NJ�%{Յu%vy���6��"]���j5��Y��nB�*&=H�wi|<��_]�5�ǚͧQ I{��������� ��6�1��V2lc6i��V:3��i�e�[2��SXJ�e�#�)�\���=D�`�D�S����f�v N�}�8l:���T������������u�2��}J���5�R� �+�yé�����e�Z9Y|M����B�ΧBP�:�ػv�{+���.��>&��o�soٟ��}M��A��[��{���q*�yT�#�=���]��Y{9��]3�A�b�L�Cf�_^�v�X|R⺗�T������ϴ���5b�A�GՁ=SYg�3z��;��̀F,N�c�(�\���h1Ghf��[�\��aqG���vʶSi���.yX��g>t�Jy�O�j�`տl�����Z�mG����m��,��+U`n͙�.�lt�3v�v�wgU� ���ī<�]�i�q�Wv�vK�ɧ��{�i�ř��4��	k�F��D�a{5iR��h]܃�ic�ό�r.��[�]h�i��G���.�sDt�(Z�!ɋ�pIsʼJ��R� �kf�t���m���>̋J��)�C��V��/56o6D�˘��kM�o�+r�Wv�req�3_�`S�����%Y�e1��3+C6;�j=�y��v����,]��N�p�N�rWM�T�����ĉ_q2:v���r��M���t�ݷlS?-k�Z�����É� Xv:�n;�����N�%V�K0��Xݴ��j
Y�)�Y��v�����Y
M��f��%7N�p��u�!�����Q4�#J_d{�Pi(3��s��_/����~��ϟ���b�!���.�,IHF�F� 9ʈ:0�d�(�P��lm�vl�&����ʹ�De�2cE�	�4�0FĐ$2�0F1��vQ�ȤW:Q�`L
��)�#YIl�&�I�H�F��i)1��� �# H�04�LdHf)AE#!1�FL��d��"DR#f�Xs����Q �b0P�Ta,a0d؊$ĖKܖJ!,�1BDbi�q#F�4؈�a&i@�b)
`BR"H�F-&��PdbT	�DX� �f� �ѐ�]�I�	ws%�0,1�s#$d�0H3�� i�?}_�|���z��X�F aΤ�Ղ�������{ky󍈭����=]M>�RN��O����j�;�"b]}ט_c9���x�`g���TڇV����04dj��g[�N2O��?Tw�8��y�q-�߷���j���t�/�(b#hX*��g	�4�C�j�N/#L���5����=�{y�������w���r�;g���W~GD�-��t��C��i��گL���!�I�o|6�'�R��yH�b)�#>��xs(����U�}a��!�Ď{�|Ecu��ʍ:̝�O,Y����3�.���g��������>��s�G�*���Id&;�w���7�&��>I�j����GՐ�Se٘}�!�^�o��Ṿ3/��ϸg�uҮ&�!Z^�K���8|�&P��P��@
𨸚f�����wp</��!���>u���̾�D�BSH���[��X��y9�X�̿P�3פ{�6|����+�u�ZC>��p,ǫ���]Tj�Ed�N��G���-��ۈT|(��P%~�5�6zE���r5�)�ʂw��4`HN�(��~����7�ݥ w�HY�&lmv�
��[ʌڶW�?D�w�y�NH�9�q���8A��l4+r���7�O���f{�kz�\����<��'�Y��$��8W;��O�)a�%,w�V�0]*�p�;��v-}�W�D3��z�u�x����u,�+��f��%Ũ��DV%wf����j��n�RE¶�9Ηp�� R�ݣ�m������>�/���Ռ��~e�����뉮���R}���T�O��ޙėR#HŴ}��}~N��o�Wfo��|�<+�;�f2g_��A�L��U>��N���dxf1Z��ͺLq����k�~��y�"�������g���r��@!}�lQ֯��;�T��H��Z22{��T�0t���l%O��u����w�x������~�Y��y��#�J�u�sO�	��h��ؕ�^�6�:X=>v����7�O��:�ǳ���p�.��R��N�|�3ݢ7Ur����C��U������^��"v�]�����H�`=��{24VY��^ՕnǮg��d9��/�����#�7=��xFz�)`f!P��y*�I�c��n{�L�gt����Ƒ�o#A��/�R�v�~��|}��Ҝ��l��5���/t�x1*}<7'n�7�G�3��H��i�]�<�G�bo?z�c�}>Y�S��=<�myt��ػ{{Vp!��Tߢ�@W��Q���/����0�h��O��#}q�*%Z�q#�䈹��#��VY����0����fТ��pGc����Cw0�'G���p�!�fn�Ij��0S�)��p���4��Xm�K��F�Pff.����2�Af�1��Dn�분�� \$��`�b48�J[����ٙ��/)vD��c%Nh	r'4ÎlY��m�Շ}~��X0�� ����|j��If��.��G7~�M:༺��VRYnPLy�Kq�\>υ[�\�
�3�E9��K®8Sa�>��vC�c���>�s�1#ns<d��'����ީ���{�n#ı�n�
&e-"j"�}BLy���U�Y�$WG#n����+���SҢ��ng��ө���񁃼|b�1A��!2�L�B�s�v�����Y~����{t��l����;6����������x���=qN�*�O5~�jNv��TbDޏ@T&�q�
��"9\?��ɍ��W�-��H�O��g|�z�K'$��G>�Z	�5�D��뙺�B�p2C�Y&��g
����k�c��yݑ��ɾS����jZ[��U3��1�f|1}m��-q�O�I����ՙ��e�NGq|&�ҭ�ʮ�+����>9y�~��]���z����9~�틈���㇀Fr����|k�6PC�����E�����|��G#���g]��q3���}�+����F��'��5��CvD/,O������X5]��59}/2�����Ҳn�#�ҎF���fv�9���Իl�q- ,���yb���~Y�njO+
қ+���pp�bgN�Y�ܾIs���O���6i{��\+���M:�
T9�6�ԩ)&����V�Oo��|w�UxX��(�5�7#U��;�w�Ͼd����~+���f�u���a�Ͱ�)A�C�/%+�@="�]P��z �{�,���&�u*���g�ƾ��]<�gn�)G�3Ǯ;�D�O��X鯧��/����O l�'�O�%�^�q���\/S��a�Y�g�*�m���C�����Ƥ^G�TŁ�?�6��O����O�E�fC�����u�Gg���)_e���v����FXz3�z��Y�l��!�)��BGNf�y7�u�g�R��6����A嵝^���nM�����z<\�o�����=�*�!��t(x �
s>n���M}վ��u�gT�=T��>�f��_���o�'������3�g�H���0�n��nǧ�.���B[z1z
�LH�@�ɨ‾�^vY�B�5�\P����]{������;�5O�xɺ����\Iy5��B2��Hn�FG
h{w�f9�j3���m���Wj��웩��]s�}�;�e�T������'Trv9��T�}�V4[�IF�;�J��q�Rcp�ѐ�F���J�����Kk�f~/��2�n�8�<��oy�󵻼I�O�&S�.[� �G'2�Qs����]s�otf7{�y�q"� q��[z��|Xj-�c���g���![��8V��pÜ����d�yɵ���u.�@���Y��䫘՞��ɓ��T��"��%��xܶW�ѕ8뙭��>���.�Zȕq�+�"ן��D��^�@t�7�NT>���z;�� M�'�����{'�������'%�~$Ϟ�ύ_��zdu�f��{*�oW�Y�P���]]��*����5�#�|wEº�-J�=7�g^ߧ'�2xρY����/�FB��HM���V��s�mԻz$d����Y��.S�4j�����C$�]V�?^ugNAET��omV��+w=�̿In��\u|U��Rk�g�7��=�-Um�0+~ُb��"4�S[�M��\�=\Fp�|�w�W<�����J���ȗ�����l�t�A�g΂1k��9S�O�o�9�b���ܢ�z=��="�^���q��Ў��Z.���9�"�9�$9^�w4<����iDx�e��<n^}���'=�8����g���H<#ba��%����.=�sQ����Mz.ǅiSu�ϫ!f�p���<���g"7�^���L�~*^���Rb�f�KXk[ђ�,��H�7S�J"	!����}���|��[�uvC�h�t�(bOE�n����g9��]!� ���&��:A�nMP �P�U��� _M��u�����w܌��ɑ�/�9�s����d�E�w�VR�Pj�(�}��S9��[b� ��.2���X��P�e���e���wp</��7��FB�O�vo���27�F�y�[����W�ׄ߰��H�<UL�Th9��Ϥt��{Fw��~W��Hv?Eo@w��9��w�e�A1�i�Y"��F�|���@hGV��a��q��ߥ�!e��&g��C;`>3cLG�����z�t��
��5VCw<D��FH>���vwM�]����7�a�/��bv�W�s��V<3����T\N�,��L�!{'=�g'�GL���y��P� s�G�.���G#���y;���&{��|�½3�ϥ�lɏ���C���M]7R2����ཇ���I�S=�|��G�܋�^�rȬ��C^�����6E���g���gG�=��7�6b�n���\��k���7�U#Ы�##'�'E�؃�.���7���ۅ�'�
��]�v���nΧ���eW�Vp�����Z��Y���b����>����{�ؔ�h��X�0J���꟩�>����{�z�\~9�����p��ց���;[.�a*����cV�mќ����u���J�����J�q.��8�/1��YG�E&�_3ۃ.3p�c��ҟ#�[c������ڞ�ӗ��R����k΃ը�(����V/�@�O�r-h9���<�{8�t���T�htξ=�*E_*��Ι3jp^_%u��z#�s's�#Ӑ�~�H߽g�Y��ϸ�?g�֋A��p*i�z�Qb��LX���啇<�Y�HV����̜N߅NC���>>��vT��y]'��5�]:֧��~;�,j9Vx�s�*;�=}n�<��y=w0�}�%Fz��]������ڟOlu��(8��^|}�������ެ�g��KR0ﮏ�����1p�����{xO��A/��?��O�\�_��Y�?S<�m����O>_�']%�������u��vG����5Q6�����}��\j;��5	a��o�X��3���
�ȹP&|��)��³�6�~�	"�{��Wc�b�u�֯������n��N�D'�����tu����ۏ�;���	��=�;����wg�3�vۇ^�t'Ъ��nǅt��*zTW���@�u�{a��y�\���<̏��(�\+��!�s���^��*�E�]y�,�;|�N�~e��� �>��ǽ�>&�?8=�'tS��y4�R�V�%�@��#I^��/�t�����\y91������������v���������ښu]{o���̗�Rth�x����7 Eu�IL٠E��힡
]�Qϴ8��B�p���]k�=�+I�ەpI)�>�ք�]����[A7�*�%�V2�r�3&��ꢑ|ֽ��f�
5qk�R�����8�7�,�ع/�ws?|1���E>^'C){񇕆���
��ʟ�k�q��ҬǙeG�8�#y��<�w�#��L�1�s|=�@¨aQ�e9��d��KF��I�/���yxΝL�K��l��ym��g���FC�A���#��z��������D�CW���w'ц��Xw�}��Y�b��֊�����u�ϥ:��(}�+���nG\F��&!{`��ةj{�-44�eYS�z�ag�o�5x!Y��i������#��2}|�?Wx'f�dvWOw�"�}52nc���m��*v�J����
�`!����5O�,��\̜M�*Yޡ�Q�k�������5ۼ��M~Ve~S�����Sh����C&�����D���������;^C\1y>>��ܛ�2<�W��	���qݟ{-I���7n��@/���<̇W����>���a�I>s�����>џ?W�G��>�	�(Ք���h����Wڸ���GF��j���7��)i	�wTǡ_�ɸ����������o��ݐ*�!��!����^��uKgn=��V�[��3	턌��ty�m۵d+�Z3�~��,8�{��T�VB-���0�$8.��yt��R�/�v&�#�јq�q��yt����ek��WƸ��6۩֬�PJu�{���+�C&�w���h.1�Y[���&�Q^3>�F���Y������&n����y��~�Ю3�H�l��37f"JlF��Y'��X��A��Ɠ�<Kߗc�c����qC�V�|=��v��zx
(Vg�܁���{��I��������@��z��Sg�\p���~�c���Lm������˖'�g�9�Н������YqeO����G��6�j-w+X�a��I�e���*���룶=�����J�ds���^gA��=՞��&L:�URPc�����rM:�3kמG̀,ߨ��<�T�{�D���WdE�?X"����=�c�^�@g*^ߢ߽��g�1gv@�b�t+Ĉ�w���F�p9�\��w��>o�fm�����zdr���eT��mG���zr���'V+Tk}��
��CW5�#���ߕ׸yjW��ν�Ju^ПxρY�����f��Xf�޺Y���"|���jql�����>���_Ʃ�25S��w��d�k��ə͏�<&�o��c�[~�}^�u���ܛ1���U#j�u'����a��.7X��e}���+K�?SLj��oLT4<�����F�/���|�ּ�``W�ce�A
Km+']CA��J\Z�<�ԕ�Ӆ�
u��!��tV2��Y��ҳ�ͬ�bg	Ds�������h�*.�W�nT�MS�'�b\���W&G��J�_�~���߆z�X�y��P�����l��uNp�WJ��>��j�47���ޗ�Z�W����Nel��GB�~������\oc8��5��0<�S�������v�T������Br}\��ȸ+�|O��Z<}"s��s�������݂����i���ok{�O���";G�2�㬟Y0�;�o.a�����+���3/���hۙ��Y1>Se���ĳ7蛠�A�<~&|�r�����~�>���>uƦ��\Qq`�?�;e�����Lצ^Ρ9�D�w,aT��Q��k�l�E������w�pON�?:��o4��Yq�җ����՞������z��Ǩ�FT�
�(#^"Cu�28S�s�V �8�s����w���{0nu9�S��# {:��Ǫ�@��\��R�V�P��#�x�+��P[���3����m:3�����u�����ۄ��\��������T\N��1G�Nz���N%�����gf�z2��WbgE�]5�s�F��Ĺ�ɩ1��b�Ϊ����[j����[j�����ڵ����ڵ��[j�����խ��-m�[o�um�[o���V���Z�V���j�V���Z�V������m�j�V�ݫmZ�{�m�[o���V������m��kmZ���ڵ�����km�e��km����m��1AY&SY9|{�߀rY��=�ݐ?���aV�����T��}�IJ-�#CB% �[6�"!I���Sπy^��fM�h��,��SU�k��k��Y�TW\��[i��Ei�A΁��x����e�M+l��V�V��hi�+1V�ͤBf��3[-a6͙�^}�4�ۼ�K�
z���%��f&��W.:���Q�\�C]�W&[mS;���Eͭg���1]�)\��m��`Uqt�< �w   ��   v�   X� ��Ӯ�4�r�o����ܴvή��^�whg+�j�T�v�]SN�;�Z���F�fwpJ�]-����P����ґ졙�")�X�%��2�ꃷn����t���c��+�l�sp8��99ŴGx n����0�iѧZWm���V�n�q�I�5�tӡ��ښ]����u�FʒJ��ST۝�������&�x���ֶԵ�7f�n�:��-��5�XC];l�el˻������Cm�A]�ŵt �j�[jk������ {�B�*5��e�E�N�gnt�������k��7)]:r;���0ݕֆT��úݖ�Cq�ɷ6v��x ��7��w+�vΩ��M;�u�J�vԩ֫�յM��P(�6i�C[�C�]��rskG#���x =�%i���kA�ݹ�m���M�m���r�e�gs�ݤ��]�S�Zl:Ӆ��� w{o#WY���.�v���!֚��]���[d]u][��Ͼ J  0J���1�2���a���U � � �  E=�&��T�       ��%IT4�@2�A� %�U=��~�S�m��2 M0A&��4F!��MOSQ�Q����Q�l[$ˡ�Q�3�D�:�3�4�x[�l����?��Q���?쒈 � �����1�i��BX  d�qܟ�������G�p���z	 �  (@�!ʐԐ�0)B 4���n���9 ������?�p  �����,*^����>��?j�K���C�~U�y�(dEW��f�n<�{�#joI�f�U���ęb�R"�X݃�[t�n��ޘ��`���葴g�̰�rQ��錄�S���s$��)G��b���:L�0*̰��D��a�u�$2J��U��32�e(^E�������)�i�7���-�tK(��e���>��C6D2#pZ׆��Ńq�̇6��efZ�2�Z�X��T�O�8�9tod֫q<qm=�Q�"86*k"-X���`�f�̹�nc	<��K�V��`�R�"��V�ɮ2�|���&�Ea@�7E�&��7qV�8	��Ot��ӵ����9/U'V[�B�u���'���]-9A����cE�V��DpZY����6T�~�]Yy[aw%ŷ� ٭=�>�agQ��l��aɟS��M�鐄Ѝ��D2�G+2���3M(��#��<��P1��mҺ%f���0�tuZF��E�t��<�ENowfG!��b�*�քYV���FG�B��G-�x�j� >��}��C���Y�c1������H��֥1��W��݁�eixCq+��2�J�<�Xi�)�X��dي�ܓJw�ͶKiɂ�ë&A���ۮ�o-k�g�O�n)M>��O-�Ø>t`g{a��)�-��)�.�`�ܭj*�ajLZ�͕pX�,D����ߍ��V�fٹ2�m��k��^8�4��z�FĬIx.�,�;Xp˘.�9V�n������;���P������U\,4�̫S:X
�V�LLMt���ܻ�AT�1�2n�(P�b����d�Ll�)�u07h<TM��*�d�N�����;�kr�ͦT�L��-��L�Z'�Gr8�Pwtɚ[�%뤎	Ǡ,�R�d.�E��b+7mݴ�[@�Z��*���nRr)N2^6j��n<W�7v5��^���E�y-&Hܺ1�7C�*gp
�bb�c�$�����T�fb��TZ���r?�G���F��Hm�0P(5� ^�P��" q]3t�L�f2�z�ݣ-Z�6mR	��ոdw۳���Y��e!L8��-��`�lVn�{�,!:±���B����%��i�Bn	U��S+u��%`�d!y-��6�\1Ŵu9�L9�-��E���s.�Y)�S��"�v;͚r+ڌbN��j��%���[�:���y�&���ef��i m�0�㶌՘ea�@�8�f��y+u$�?�1���Ksn��fb��S(P���u�(���H]h�<rm�YDf�cw�y6 U��O������$��8��f�jQ�/lcݹu��E�[U��ȫ��^a%�5f�1��-�T�"n�%'J�cu�T��l�Ú qەz
��b�e�v�J����#$���,#�J���A���ޑ��oX�Q�[�Wx��W%2�U�W�%HX(nh��2�Y�wo���G-�5l���(�=�ֆ@Vm똱�"Ot�"�&U�QT�ۛ�I�xj9���:�恲Vf��,I-#hچ��e��7C��|�:��g��������iq�w�%K�Q뫼u ��	�QK6�3Zp<�5]�=����	Q�L���]�[��� G%�*�o@C*e-{G*��WGi
�s2TA��U�T�om�QM�Akl;�ke,��BM�19�tf�ۊ�iF��'H��C���6� qRf�Z�b^��h7�R��s7*ܼJT(���sa���:���/<���`oҭ�E�%	�i5c�24�u!�����;�6���[N���ce@D����2�
in�u�;�����ƛ�]吆�j�^�:Ͱn�7tP�.T4�\�3�PJ���X��X+T�RT��Sr�͵�)���Ĭ^Ķ���P���$�M4p(���d��˻��c��s+C�ƨKNi2��;aM�`�wE�t��YSMĀe��i�r*D�$ ��C]�ŹX*]2n�ԊN��"f�!e�%�M�3�af����]�Z�
����Q�o䡬�*�eJ�p�U�k ���x�D.<�cX����=/e9�Uɺ&ڻ���z�/�j��̽.����,5*���#ݒ�[��w4H³r�r�a1�Te��{B<&�֣���n�`�[�����h�� y�$�]�p#� �;{��1`e��)(�����lc��7�6c#vӦ`�j�=��+�/M�`@ݭ� �:7�!)�w1[�T6�-H2�	$���x�-G5�cM�pLMEY�fʌ�i����i�	�܅Էc*PM���N*pФ*VX�t�U-oM�G�v�����$��M��6���۠���aT6��am1Re��mYH��(�������D2�B�7f��&vu=G�H�Q��b4U:OC!��b$����&f��#i�YX0FU^� hL�&$���qZ�c��n��0Ȣ���51�J���˗��i+�壶C� �^P�K�ª�* H����G-&`m�ŗy��P��7F=ڼ[�`��VMe_QT���a��)��B|�Dv��u�(T�[u���k�P6hQugtS�R^*
Pܴ(��۰6��Z�7�¨B�ޘ�7�����QP;�AeR�[[QZ���2�]�&�>�iJc�6�Ռ� �+da�vgQN�60V�Ȃ
J�R���v7T&�l(��YR0�(��WV��e�(��7�V�������m1���nJ��X���a$�i�g"4���*.ŝB���E!%n����J
-��̵�����*���;�`Hd����n#(��yX/"{oT�5Lf�NfR�U(�̵���F��ӆ' �c2`�FM����N�c�Ӈ$˖76����jZ@�:��9�L��5$H�ˏM��-f q�;p��k�f�A!V������D�����/c���Je(��KifY�0=�0@��\�2�t�-���B�Ә�R�Y@�D2�d�����Ջ�$���^���j�NE[_,���/�J���X#jT�bf���xk3r�Gmɘt��e��%�� a�-�36�`��D��J���A�'!��F����E�Y�f�8�cz����U#H9K(n�H̔j���w�����ɂ��-�L�XzVc��Q�U�ˬ��J��X�(1�0��c�.+�{f���Y��l��<��q=Б%<Ҁ����7\Q }�����r���W)ǅ3n�du�F�FoY�C�j�ܬx"bTL��6ʺՏM�hS�,j�r��M��[�T��"wCj�.�k�S��-T5F�G(X{��RL�Z�iͳx�J�!���lS�C.y��dx�M�1QV�g��l��6Y����门d;[SYY9�*:1���DkjΣ	c���r��Ք\cMԉ�H*�N[�b�I�sN�Y�:��>D��8�2m�;��L]\�(?��w�M���
���A�Aշ�e̙��]�����l��P̃ mk�i��N�M� M�Wh޺qV�ocN�;S-�F�KS1���t�*�OV ���y�ǍZ�D�$���P7y��eWc��WC��a�Y˖i��ѭ�2ڲS5eb�s0��R�4U�h:p��e��"y�e��V�L͗CWh�_;�����1'�:�MYL���ȬLE⁆n+	�f�,锥��`|��y���E(FNQ�.P�:,:�-:-a���m�M1���̆ڊ�w�׈:����S2�J��h�^�[	�S�r�F8t)�]^��tF�T��AQkZڳ,�Y�E�yR����_����*�ŌNm�&X��N�Q�P�x�b�v����̭����(�X�5u�Y��W2�3�J�%+e"�Yڴr��x㊶���	�C�����P}��Bc�~�݅A#.}�}��w��ʨ}tы*�����h��D3���uL��        p�n�f                                                                                                      UU��]7���Ъ�&��D���9���eӝ(MpkX�D��j�yl��)4�[�]X�����Gj�"�s�bFn��o�] ��rm(%�k���S��k�
M�cL۾�f�&��Ń7u�-*��b����3W��Y���j9��SF��3fˢ�DU�71� �]*7Tp㰲n�nPH�t��LQX��o0�uQ�(�MZ��4���#p|��7�Y�o���픴q�3_J�@����+U��]��,2U��m����r�,�k��|뱝Lv�qγ�IWzM�+�4ޖlZ�ʖ�����[Z�C��$BQ�|�e��!�>���\�,�}�ŷh�;���0so�$����k���y>��gf���:J�Fk�,�#�d�C�"�1ROV�E����/Y��#�il�{��	�0�3��\��m-��y��T��J<��6ލ�X.n�
B��ҫ�Z0�/:��+/z滰xd�{uU+)*ƊH�f�}Ǩ��2>$W�hJsXy2����Kf�a=�r����U�}Ƹ��$�e�f<��A�n�ܱ�/��R2���,�5��7�S�}�xؾV����їm��a ��C��a���B�6�;x�z�k8�+��t
W��$�Vv�kFen�����;	�*fIM�%BM.l�(�ًZZE�Ŕ�[�Qqm��L�_ʎ�+5��P���f�vS����Sl�o�������aWٱ��U�q���V�x������VADj�-�4���ᵜ7��YOYw���F�8����cB�y;��5��P���<ʖ�ء4V��c�ȞȠ��7�M[A��<��qY.P4���_V+W:��U�z]s�	Fa�����i��R�Ǌ�ZK��B����'Bw(GP��Ƙ͛�E���4:��]p�L�%����:��-X+�k��k�����K���z�f�+G+"�lܔ4�ǈKt�u�-����p!9ΰ��]�o;�΍,���"�F��6p"{Uj�x�g=喉6س�[�
n��a��������ٮ��bRy+wq+��q�]i��S\��j5�	ڮݫ[�Z�v�r��y2��)rL�M�V˂ְ�F�g=���{���d�hU;��+�x�ղ��r�}��\�����#���w*��G-_UwT��&�2�`�`�v��@�Т���v6$]�`E<�v]عD�x�E�f4d����wg�r�:��T�j'�+��S(��8.�1��h�<�:��V�����e����; p�͕'��DQ��>ɰ.��m5�qD�$�A&��:��D��u.�jNnP/Ue"��5��5C�=�#1���uh��Ћǘ��#��ލ�LFҋo)eQ��p։no-
�W�o^�f�����DE��n�Nʨb{ ���� ���Z.��ȷ��m���ciqY2J��sQ��[�M�쉭8(�G
8沲���R�Q��&Z�ǫ��r��h�V����F���؏$��:x��zV�sh.�_M����j������\�\��<�+��5�ɬ9��3w]Շ£�\����d�@�|fӺ�㸚�-X�:�LU#�Vs�{�e�и�%VM���M-�WLg=�kxd4��B'Rᵔ���;Y]bgm���Y�%[49��1�p�-Yp�|&u�w"r��|��P`�X�")��O�)����9��쨍����5f3�Z�뵁	1�u�[YmW�K9�JV��,I�J�:��mqB�s�۬� d����1K��G�"���qf�2G�Z�>��Mr'yݚv������	Gq�g3k�ىgލs����D�՝f� _j�8UGό3�X�X"�^��
r�\�ш���s�˱Z�7n�rS���6�n2ũ�g[�n ����I&�
�5�c#GV�Q�X�����YP����>����L���XS�>Z:敖��پ�Q����+�Vwv�גK��n��{([,-�[�t�1���!t+ot��F^ �ꥵ�r�k!;7�7[�R��o�]��owj3���A� M�5����3,�I7շ7��.1���T�'>J8+|�w�1�8�n�Î����1�v,\���*Ce�(]ز8ں+�5�ǫ�w�����鼦����5��:¾���<b�/��}o��B$�ޞ��7�f�/�l�y�ՌR��A�Ts*ب��@a뉪u��W5P��r=vUӦ�EmWa�{ٲ��j�}d،;�ŝY�kL!N��	N���]�T�,Iŭ|{��A_:҄�#�mh��-�݁]_T�Ib�6N�z�a珮������Y;57-�bANK��K�׈:����fH�ı[�x��7��!�7�2 �:sn���7kz��sYǿ`ȵ:����2�,�Df��k	%`/U��z#a�&�U�÷���3	�o��D����q�/A���M�ۖ�2.��)G���#S���̽�� g*BRާu.�DV[������L�+OZ�+\}G*pL�W�/y5cd�]�C�?�e�G[C��T�J���ǎ����Ǆ�}�����wT'�{���=�����[�dMm��K�ܭW��-���9�i@��.��e�*Ӳc�;�k��V�u�����:f��#(*�����f����%����Ʒ��J>m�*4+v���>c�cFT��2�̫�R�E׼j+�}�{F�pM��9�<�6�.��hj����p�5q�O���h�ħ^��y�N��Q��u�j(�0Uar9�Mc�\U�ew�&�O	�Z<˫�پ�w�#S8�f�λ��Z��S�e��"6 �om1��[�U�b켮��\��f<����ǉ>�>���[�#�!�� �.����T۾Tq��=t�ԩ!�թd�i��yٕ�70vY�x��:��)�a�"�8�X��]�k�}մ��Ӊ��ķ��Ït�nV.b�]uZ ����T&]�s�dȄ"�<�iA��w${uF���^h�vN��*�ņ��B��eZ���lq�J�m�`W�&<Z��.�#諴;��+��y<�iv���	ˉ^�I8�+�^�M�׺�5���Vւ��fij�cx���Kg��wْ��4�١цõդH��xK-�����BYK����$��]��i�ԙ��Ρ��y� M�A�vb�I�є��p����1�keJ=����&=����=m���74Z�6��ճէ��� 5Ǆ٣K�
,x�c0>�XX�����2Y7٥��s��ϖ���;�� ����e��Ȅl�Q'���,g3Wݸ�V���c�u	D$�+�Ԉ�>�9�*Vsr��e:g(�ބ�,�b`��zQU���]���C�BJFĠ�1vk���n��K�o}���XK�=Ŧ˰\���g@U��|��Y�]��^Ķ�0����ܖ�A����r�IHAY�e+vc��Q��h�k�n�ݏ[Ɇ)�����!��\H���V�:W�zٍ�&��Mp����2J�|�Q�|Ep�i}g��7,�������bd��+��חK��P������+WH��qIh��r�{��[���#�]�_��J替�c���5!���^��8o�G�[ԞŚ�poI��V�r��ё��
�w�,d�ʾ���j	�wٚ                     5=]���N����d�:�Iőw W�DEESq��3W�                                             �=fn�gM�=9�=U�}a��6�%��\Nv�����������~_����&|��� �5��B @�� ��!�>J�T��$ ��*X����Y䷤4d���Y��yD�3Z��!��c/�\��9X)��C\�/2�h���*�puX�J���x����0�B��n����v|�.tX)Ə��(.�X�+.�вa}H�-�9��;t���X-<)�E���05�m��[V��V{�Aw%�7�Q�p_n�׎�N5��!�ã���U�[��Cmh�K(E�� ��,��Ę���kQ�y�����Y�(/�"^�,��@����C���mQ�E�}�D/������^<���\��.�C���m�^�䲑ي�
u�냻7�oR�**4��TLY��9r�R5��U�^X�6F�u�;f����)s���ϐ���߃"3j�`�ħ>��AVi���Fi��a�2e���f�!M��U�**}�u���6��+�J,^���\��v��C�-n���m�7U��m�� �WpVᛔ�"㤜�<���[��9^Bɉ;�Nϙ��jcЉ(+��X�F���%��W)��֍��k�]��]]�3���#'m�����5��՛a	��TE�)[`�/U�J�PJ��7�B&�I�.��#=�Y�Y�f����e�hXC]۸��2���]b\۬4�3q3t1p�j���2����
��t�Y��ׂ��TU�Gao!�Z���M�f�s��t["��vk�r1q��Rk�I�m�6x�\���>�����cݫ���+�Ǜ�u���������ҡ]�f��������G2���@mޚس1'YZ����n�Ch\�Ѥ��`	X8H8tޡ�{&N�r�XH,�v��*c��Q���իX@�j�̠��rz	�F�ҼV�B��P��R��m^P�C2��2Ȏ�ആEm�nf�ԑS����\�Oܗk]��%zrs�f���SM8�s�i��ѯ�����8cg۹ق�+-R�����ݰ����$n֥�-�{�����ɠ���%�q���`!��5����!/�就H��5t�K��U�n��{V���J���֋B���س;�>]8��
�Z:|��J"��U}�P�E��3���]��-̡�r��ۄ{����#q�yd�ΝA�5��L��^�J�Tg�Q	�����&�<W\�G%���yQϜ��d&p���-.�#|'�=�g ��. �ܗ{9^��M�KF���h'3Ndi�Qn;9jgGx���!Y�)�$A�k���{MLepU|�y�Y4��}��<7~���*L�h+��ޑa�t#���H;4jO����(\S����bS�N�+p���"�R�{��rVY�'1pb�!��9�(B�yd;�i�4 ���8��	(�t!�X_�=t*�P�:�JT��7��SyznF40^20�h�"uMo�~��ed�,�)���de��Bj��lw;��KV�}���T����l-+D\�S�8[���lf�Z��֪�J�3r��;�o��+�%�Ŧ�Y�F �ʇ@/R����:���͜g5�T�� l����mV�x��
ڗs�"Y��r���;���ξ�c"o/ᆧC�y�W�q�
��x��l�
0ӢKT��w��GS镵��T`��b�L����vb�{�1%T�!^�f�A���B��H��I\��eǩmbY ��\r1�hP��� Bp�p� 6qBU��-�{�v�g�L<���{j�r�<"ƕ���:�W]�0�?a��D6jO�Vv�nV��i	H�]^�XѢ�Z�Ep��kJc����ӛPm��u�/D̬x�d8.�ξ���;H[C8;����F�%�i^�U	�έ
�y������-o��2.��$���t��&�DeLЮ8c�녋�P�(�h�9��)r���OH4�>�����l���Fe��s��5�]��A���k#�=�%�+����!]�q�k�9NP��7����#$+�	g�6�U���!3��F^̶��N^�Vr�
��)�1`�� ޷�j��%b��KX6[�^�4$���Y��U}�P�/~��Ge��BV�\-aV�MUڱKs���8�J$�\ﲆ�QɊ��Ս�u��,ϩe�V1Wn��
��p�N���̻�pݤvZ��������t�c��\��B�c�s3r�t��FE�錬���*V�Xh������t�y�Wyu�a�"B[ବ�[J�+F-����V�G�Ӛ�Z��Ƅѵ��ZU8+����Zź�x���3%J��Y8o:�%:�&}bD4b�gq1��Vçg,`J�*W�/)p |�@+7��(��:�e�d�([�N9J��u5�'�:\��Xw�G��!a�|v�0����s���L\����M��!V�N���F��D�m�fՁKκ�ZLF�Vb�>���8������wX|3Z����E���@5�[��F3:���,Jt��śk�Ukm:=����ަa�Ǌ��yp4�>��T$��Z�
�wh��Je���۽F�C��p�7.&�E2�eӑW���r;�f�W��fU��wW]�V�9|�Bg�q^;�������DR�\Qg�fȩʝR��㾫��p�C�|+��7�oP����v!Nn�>�h��m��ք�z��04��x��3K�~�3���I�WF�[��Y%Vs�A!ɥzq��:ѿ�ֽ�9Pݭ�])f.��Ķ������꽌|�-ˢ��,�o��HJ� tQ���V�ֆ�	�;�쬿����9���Jp�9a>�O@��^�tK���"�J�۸J�}[��#�k�9�7ݢ�M��8	�SzN�)m�9YRg>}'Q#n�:u��*�wբ��y���={���H6�1�ʮ�YW|K��(����rhO�7I���� �y�Nf_�f'}ZC:�=�����l�\T�"��u���kv�2y�Z �yZ�v1�뫶c˥��#� ��*�͏���@��*�e��DK�}���C�%�6�o*͢�����aa�w�ވ��3K2���(H0f�E��H�:�
e���e�\Q�٩n�U�bT�NiD���-�s���Y܌�6���v�7� �M��fi�y�2IM�T�5����A�`|Ob�`�_]�ڻ���U���Xxh�.���~H������QZ2E��eo� �N
��۸�BT2T�5�D�p�`}O��=LWIR�.uh��nnG�R׽l��{t�ނ�ac�f�C2�;�mpVn�Q��jkjk�w`͙zM
m�oL��Ŭ�e
�1��/��7r�.�wR�^�V30���{XRj�+J�Ÿ��kaK���u��՚��+T�u1�Y8ZK;�^YtFf�n��&�fօ-��n���I�]�7ӳ�@m!��r�"�4�����m���X�.��t�Y��5��nJp$�Y�'&�j�m�$m�&��&2n��L�[en�^�	���r��V�XOt���3$
`��yqֆoX=�H���f�Hl@r�E�[{;V��P�0���p�K�A���A���>��<C5Al�z������'Lစw���� ��B���N\�Gr�[�`�" �q;q���ӑL��^32�ۛxqj�F���I��j�µ� ��TA�;p�:ꭹի�b�^��/]7,�!YDU_Ug|���^�)}�Y�\�,�P"GC�N��;5�P�:����/j��:�5j�;�l3�!���˲v2�#Z,�Xv��Ĳ��bz�d�RX��۷[DJÃ����s�Nb��Mۙ.�{�=`P�F�+�c<}�K�P.���t����+��o:\�pz�w<���T)�?R^k_|� ��� p������� ���Y(`)gq�����{�        �=�3����Sx�t�8�M���3�BҰqp��׆��*�6)7�@H{�P"����R��E���Y�i�@��=�Ƕ��VK����-�2��T�	���«+2IFd�ղ�')�o��oA�\䒖 ^X�� ɦ���Cb��u�ݎ4-�yz�u�˹uc�.�o4���k��ǿp�W��s��C��d
�绎�l����Ar��
8�p�Ά,���o@u,3s\Q��%^$�ӫ$���2$�'*�w)V�n�=�3v��Jm�ޒ��=An��j�[����N/
�xl��T��g���k4q�ӎ�6"����5te3�>�uq�z�I��.<����]�no-�l�0�qOۺ�]�uz  �� {J�܀�EY����6�)�%1He)A`�,b�"v�" �Y-'�KT��
I0���I"�i
VE��4�HZH-�hB[!�2�B(,�d
@YQB���"E	:��
He
@�VB���b���- �"�3T��V)(�����a�	���]{��RᣛM��+��hTr�qʂ�
Q�y�M�ˆ�v�4�_��?����[��F]��W�r4������k���B��4z<�2��E�J��9�0�\�ˈ��iBC'��w�ي��{{Fv.F��6��K�b��a�p�[���K�ŘɌ!|h�YYW��{��>�'�K>�co�H,1ӕ�H�:ۘ뙛�6��k�!�9őM�F���K8VVߠ��h���	�g3x���z�W�����]��u]��q�=]��B�l�s��R�;�rC܇�ﯣ�ƙ��M�����'���?�㿯Ǖ([�x��C|B�M�]�=<��S�JR��>�rb�&G�<]>�l��6
��E�}�%���'�M8iE[o��J=ug,l�w��zk�z̜��lĢ�X�����ϖ����Op�!c�'�֬GZ��������O6�? �^���z��^���軁�倿3WΟR:��gy�1��1-�~���9q��T
��.��k��d=B{��{o�}Ҷg�5�i����[�<�
*g�ՃqB=�Q�bs�*Ӊ�U�}�9Q�Y�v�Fd��s�_��=�<̯m�5C@n���SJL�Uy7�C�my��U8o��Pv��\�p���_H(V3���꛽�]ަ�"�;>L%�����w��'�fۤ���#�<�9��>�۸��0(��|']������8�"I�ɴ�{�a���=�Ǭ�<��9�/5{e�#7�	�T�xb��_xVJ5����Ko�xE��%����/*��^�(�k7�jb�+j��ѹ%�4�J}��m�+9bx�l~>��G��<��<��ٹ���xa���'���x���^�gp+��v$�lN�m��?"�/d�G�9�Z�C*Yb۠Gu�|& }�)��]�q�зj:�����#��T��a��~R�}{s܎v߭�G�GN4�����v�u#�7��%*{E�Z�7�T��»�O�1���F	�e�<+7Ui��f��q�w�� ��N!2s�Ƿ�u��v�����2���J~˹�՞4ێ)=�FNL,�_$Ϝ�3�$C�e��
{{S�}F2� �����3n>�i�J����V7qn��N{ͭ���6UN�j���2ո�~��i����i+��j9�\���<���x��v.E=KeéT<Z�{��E���J�31&���&��nYL�:je��Oyo�k��?<�'��n�����yJ���n�_������U���MX���ʯ��$~�+��i�@�=�w�g�|0y��"K����8��*�t/�]m�L����!����s��Ay�L�����x����*�z�C���q�6mt���Y�^��5�Z��nI#^�G�n�=�{�����
�$��
4S�~�hק�s�� ��_���3 ��]aa&k������w�.䘼ʹ����x�u���-�����~�����Ƨ�~�@�[a}�5�j�����)~�c����*sǳ(���G܁��n����M:�΃x������<'�<�������]��ܮ��KH��:aC��n���i�%)�l��*2���=��ȣ���6e3gr��\/����]���R�o/��6J�kF	�9TWO$kw��+����w���F��%z�טE_�$��c�2ֱ���u�{����'a�|��i��7��yI�&I�o�)��7�����B�hN��g�s�A�s���|�`'ٻ�a@��3j����2�}ή"����Z�%Z��f�Y�xunH�O�=�K�^����˚���l
�d�jF$�j���	�j�;Ʌ*=
�"�]�<��P�WgT�A��hI��)�����m����RzC�2��O4����L+��W��k�fT�^s�оX\fJ��]�IqNy���)c���a���`Z�Vuo���oڛ~���=Aߩ���˰Z�o���}z�U���Y����ɤP�D�1e�^��l�X,�A�7IbV�r�LF�*�)'9#�Ii���T�n��Z91J�ܔxr���:�3TϮ.����%���/A��T�z����{�lx�¤������򣂓��Y�v��%��<n8����݈$������MM����Z����r'c��� ��v�`;Z����<:G�q^o`��s��������=¼�]UR���HGS���|��u�̈�h��l�Q�^S�Ϗ�a�U��c<�ןZ��v�-jMp�UU�JxM�����E��y�U�]����+bje�rD�U�V�LN^�j�y��VKc��.�'��x����r0�����k�a���@���_��1�Q��%�%�c�y����"�^�}\=��D������h��<�u��ܗ�S|x��c��4�<n��;����Y�ԛfo����kyzx�_bsz�U�ӵH�����(�|�Y<*���]:d�臆���]��c�z���CX'������ʒ�⣼�߽Wތ��z�=5u�~T�뽙6Fb�?�n˳��]no�b����P.=޾���oK
��8�E�s�ygsQִ��'eZ�L�UA`��*��D�*��B��k�����h5e����X� D.����x��ZĪ�,]�����/-���K&��%G���3��[��E�¬���B���;3�G�N."���E���{���*��,�<j)Ks��!8�ō�r^�G^�&U�u2�6l0\�Ho{9D��Яއ�z�b.�^���������WuK~�E^�&��]㧓��v4P�P���OIx��)���n����0乼}�A���P���AI�<l�5;&5�7<�@ ԓ�n�|�\�N�G���TUĽwZdb��59���c"t�z{����k|Ϡٮbs+!p��)DT4�z�	7m����U{����,-��*����Aߌ��{}Rg��N�������]s�n/-�KG�L�C]�ѝ����6�~5��샿p&-_>�Ք���Ku��;��f�CA:�K�j󳠔AgtDml�3�gS�p_]N}����:ȅ�7�Ǫj�Ӎ���÷�m�À5{�������Z�tA5~��U���/��D�6
�h�d}Θ���
��d�Ӳ��sT7q�o�,"mn�fzg��o�ViMO@�AOh�4���F)��0o�u�[�BJ�k �9Oq�y�[W�7=��e�{���tQ*x�q�kdE��]f{*k�I����<�����S���i�q��B�a*ǉ�|�G?�,�͍Xfȫ�[I�����菗�472��y4aJ�	z���(��S�3�T��EV�ybJ|�u�2|�u)��`s�ZW��`�1@�����FE_�+�Z�t-gHeB
+�m|��^}�˝�_t�j�uy�N�o)`$�O1^4h�t7��op��j�Y�E����i����Ч�]���"w��rV��J����^^���1%�֨��U]��+��V��:kh�t��fC%_0�` {��ga�6n)VS���סM]�Z��d]w����}j�3��S#�h�����f17�>�پ�o�<�h0N������6�PԾ���#�n[C��]u�ǹ�����u���
l̓�H�/�B����$�v��0nl{)+�����F������V��4:�<��-g�K�9Z�N�+hsK��S�����k{(�>6ku6�h�u�p�<���|�l�jkҥGe1RB[H�;�0�Ƨv-l���7�|���N�N�D`)w����9���         �뙋�J]�}Ư��fwd��B�O��u^P�ǘ�p�b��;7A�x�)����u��i�#���c�,ŇNrlY5��κ��>Sh����b:��՗�[��QV��%��0�$��섫ެ���Wt�I���F��U�t�r�S�5gY�sF�'tq���4�b�'jv���m=�N>����D��0-��H7�NQ���Ʊ(q��=:��z�iϡj��k)�ϱ��C9r ��'pf��fflc;�4i��5��J�f�xS�t�*4�:���ٰ�Μ�xa��:���nⱷ�L]!ʸ�����:D�yU���]�0c�J�&N[�Q��b�̾�ދ(ƺ���43B�0���  9�y���s�ي��
�̲PȱE �	H���P���C:�*��E��i(fRH�"@X
AT����u�,"�d&���CKBT�+0��,�Jd�,���ҕ*)d�YJ�� (�2a):���B��uR�Ii���2�i!���U"5T�E$QCQI5T9�E7'�Z���`�ץv:��Y�]���D���~q���l^�s��$g��|�8��Z�?\pjy�Y�A]'���w�O�w��d�ޭ(��?��%~��}7����I����i��V�ԭY�]=ssڟ�l�^X���~O��j�e?u}{o���vS;�Y���D�.�}�����:��V/a�Ab��eHAb�*9I�b�ky�e	Y�%�����T��˧z�[�fZ���z����	����R�A�O0�j������mi��_��/J����dyO4���(��+qq�����{�*Oh���,ȿ,y^:��5� ��o:��yݬ��(K�kq��X!5�FӁ]��W&��Py���};��ȗIQU�*��4K� ��Ѵ��.n���e|4��Z�8�kmX��f�£�e�WtWJG�U׈�O���l�O,;E��@m�w�A�Zk�Y�z�=>���*&]���U@�Ւy��\ƇῬ~K>*w�$Х}�^�mܕk��)��1�,g�{�����*�UEWa�>X�v�T蘌u���%t�f��[�����#z9"��Hw�c|�v�_lb��N~���~���|9W*��ea���}o7C�CV���]��}Gѡ�vLGvvz֛M}�7�ȗ%�y��{�_}��?QM2�T����߹�_�u����<��P!�޼�vׯ]�xI�{����v�����7�G�`�3��^���h�h@j���y
yo��n:\:ZC+	\z;�4��oy��;3Nˈ�Ʈ�k� -�B�N͘M���ޚR�����nz��9��}[���r��"��4n��=��	^9~݀�[����%�xl�[�ŕ����:��Vߩ����$�H%Ʀ�|����|����am�1���� �֎r��!I۴^:s�,����﫞�kU�����Һv��Y�������P�~E);G��hQ��{u4(�s��G6NV%|D:ݼy�W��|�����j`�(�#^��8�(��mU���m}�s&�y�Yʍ������i��Q뫠4M�A~���Oc�,E��5c��VC=[[&ae�};����94U�ʽrI��>t  �ȷ�?�/#톢E:�W�խ����y�l��^��f��\Ѫ�P�+̥G���1��k|;��s��֮Uٞ�z��S��Ư�Tv�k<G��]<¡��;�Q蚣�X�(m��s�;)kTi���x��j��鱸(�}�:L_��}���^��'_��{��|�ei�P旟}t ʑd�WA��A6�Y�>�ֵמ.����~���l���0����`z��Ci'7�Y!~b��y<�OXU$�r�λ�����q�y�o���m	��5P2�B`�eP��'X��ϵ0�� d���RN d�@3�:���w���y�&`,8�8�f�Жb�3	�2pf�2�PǴ�.yF�
l2q�['�����3�Ӭ�r��c{ ]��;��䶈�.a>B������Ͻ]��G��tf:�E)a��{��yF�\m����}$�S��07�����[��fKw�I�v��v�=0�O�h�� e:��m	��m�'�&��IhjyP�I�e8��I}�{[l�g{�o~zt���BN�5d�``�֙&�N�m )�$7z��!�OP�`)�&�u��׵�M��W5��g���,�r�m<I:�x�z�/7$4ȡ<C'�!��THq0v��$�Hs��9�s��p���O|��\�I8�&��&Y']$�d��)
��) �T'Tm�m'���t�n��_3�o{�!�hu��=<��2m�d�;G�����>0�� q��O'��O"�m�7�No�s�w�@�`,!��u%�N���x��h8��'���K�I&�0y@q�	ē����߯;���w��פ����)��Uz�D�I6�=�m Y�Y=r�(q$��:�o���b�P�|׾����5�=8II�Bi�D)	�*E �P$��S<�u����!�Z��!��a+͚��~߾{�OKa6���'���e2N!�(���aL��h���Ja8��a��0d�}�{��7�=��]�Δ�q��!��a8���d:ͲC�$��\$�V�S'�Rm����⤇ݎ�wA�o�I��/տ��zi�7!���T֐ѻ��df`��BV����ߣ����cq��UK���*-���;��Z�g2i�X�t�/$��� |%}�T\�9�{�-$�><��!s4 ��u���L�!�
d8��$���x��Ԕ�gTE���5�z��c�*�����6�a6��!�TÔ���	�C%%0��Z�N$6���ԓi'l�KB	�y�/u�ꯛ�|���)�I�ӕ	��)�z���ъXM����[!���<�q�R^���a�Ú�;�>s8׽��2{�nI�N⤧�'�	�LU���Ԑ��z�q'��2�l�(u�=�!�s��W�����g0C�[2z�a�����!�E$�z�i�������!��R@׵&P�!�4g�o�{�kݞ�C��-$��������@�'�Y&L�v�:���i ��z�Y�I�����9ҍw~�^p�a!�MԇP��	�N��*�/Tu�׬&}������y�$�ċ	�[!�[��ޝ���{�w�B�f�$���H3D�2�:�Y�I��F�:���a�� �{�=�=�����y�m)��=�[ꍤ�C�����6�XI��m�Y�uY�!�I%�RM�IX�;�|�<�|�8���	�CR,���C�8�M]Ii'�%�:��!�ڐ�'�P�!�%��'_}���t��;�^��{��X������1�.�c�f��t�g�]x\��p�Ouy╉���֯^�<0�Q�K���9�t���5�z��9�9�s�>~|�$&P�MVu���p�i �Bi�a5u$>Z����E��d�I��ڒ���z� �ē��EoX��Ϻ��w��{$=�e�I���@���T'��&C[�
B^�m
@.{@x�la&}�m�q��ߚ�g�s�uݝd��Cڢ!��$��=Bd�=a8�b�-��I�3<��Ƀ�l:ɴry�{���s�g{�~�S&L7T@�!�B�S����S$5���8�ǵ�K<��C���T�׼���[��j���y���Jd�Ъ��&�Lb�:����C\��%���_�Y&��l!�
Hq�� q��xp�<�k�{�{ �Ow��XK7R,�r���z�m�7D��NM��C�&$��Cg�$+4u��CW޻<޷�7�c�w�l�)�� ���IL!�rS$�W"��(�-�q��!l=H��OP��u�(b��{���~y�d�II��_*��m�<� q��T�� ��Bi���$���Hj��z��O�߼�����5ߍ�6�e$�0�)4�i��C�ja'Y8�d�g��I�M�)'��M�`,!�c�ӽ���k��;����N�	�!�C�R�9ڐ0��N0B��d�ԓ	&|��1D�I'�y�o}j����f�����|��i3#�kp��x	8�lcUȥWQ�!�}n�����C������K8t���:�@��f���d�᥆�?�P�NE�����h,����w�s�����N2�L��]��:��>5P�0��I&�q�l'��&�:�	-�y�>w=�<�g�������ڑ@-��q!��� S��������Hm���4Ì0{F���u���Lb�W��k�|����I-�a���B�P�R�1�$��x�S'��%����T<I�M��T@��]{��s�;�k;�����2M���u��ē��$�9a<Hb�J@,��`b�����tHx��~�5T��}���y��2m�:n�:��q�<@�[��N2`IēL��䇉Cl3TChq��M0�<�J粒�{�w�x�zUC��d1�Y6��Hx�]t�m��I5���q�M�
��B���6� ��N����}כ�	-����3��u �c52wU �0њ���QǨCRx�Bq2b�-�6�+�o��������d)	�"���}�r�Kj�,쨳��iQ�V��FZbv��=J=�S��6�B��u�M�p�|�1d�fnei�<|f	'�����{k|�tg=3�K��ٵ���]]������#߂��N��C�"1��W�v�,�,]��\͓E�A����<�o����I	 X"�@8£s����7���ߨ�*XD��V�x�Y���~�9׬t68�����c]������Ǡ'*e��c�P6zP����E�p��^�D��/m�s��䩻#����ߧ����]�:�g.�X=�9Y�~w|���4���7�l��4�Y=��/�Tr��]ɳ���U�w��ͽ�q�ǚ=S������bz=^���-\���hb�Io��}��E��}<p.:�ͫ��/�����SX**;��������ž��
v)���{��nOL��a�Q���s"�ָZ��~hR]���j�1oc%ˢ��ٸ��Q���e�=�Z�#ML���s�k��9�7�Ą&ВEHH,�Aa ,�� 
@$Y ��H�"�Q`���RL�O�]���y��۴�ӌ;�f<���{��Ҩ����O>�r�X�
�\w�6g�򙏡��;5��}_>1�,I��{.�eä���[9���U�����:}��h�A���J��5�)����OQrq+�:�)�{�h���v�s��D&�r�a�N��bC9���i��o�,ObX���%g�R[�J�;�MxN�g=1w.�
�0w�yu<k+���������z{s^%�n�f�G%E-�?�z���P�K�m|Ϸ1au�\v�nA���q�	�ɱQl������9v\�RG��"����>�YD���Z�M���2&�qAd@��(l���R4��L���Q�U�}
�&�7�|�6��(�d�k�E��̘:��v�gu�k9����͂����[�ٷ���9��6̓��Wiˊ��ӕ�ҲFq�;wP��r R���Uv\د����W:J�PP�%V��������Lks��Q�4�n��>�!�M.��W��J�[M��Hϒǃ #9/�I���j�1�i,{P<Z�ky�{1��vmN���`�hq*M�3����;�`;���W;��`��Ŭ�h����P�5��5�a�(3��-�,M��cҞ��$+Q�Q��]5\U��h��i+ۡ�W`xt_j|�<����*?)���WH��Vp{�Hz�Vm�~�6#��_         t��H�j�0j��M 4��y0��a�뫘	wtSc�e�r�v��TR���Ω}yՆ-�ĦH����ǽ��gsF9P�̣R�=ӥR���U؃�l�&�y͞�SU{I������P}�i�cQp�P+��ӎ����}����3u����`xMv@���(۹|�hJ�/�����!���c.v��Y��:R���/b��+��Ꞌ�²gGn��N��蹂.�caƱ�yhfpk�By��=��(Qv7u��칌<�	�v�\G
��R�wY�������,����Y�e:���uSL��W�����N���7,	�Iau�2�.�=�uKwS��TӪ�͓���Q�Ҹ7}�sj�+�&:�N��� *�� �9�o\��9�+�����*�E'�B�'BؤE@RO�B�C��
II��(&j�i5��AKi�%$\��h�I)�T,��B�H,P����fZ�e�L��J`|&��AdSĒ��`S"���Rc5-"�)3�����W���~��R�%#�=[~���K���t�Oa��t�m�hYu8��:��������w|����-�}�"V7gO߻����?�aC=�aS��M�����'� �t�oC�+3oD�o1Ը�\��|7�ˆ:��b�_4M���F&3��<r�REr����Nu:����p�ᣌξ�Iݑ~�x��B�
�`��,���y��gS���^}#��}�j{8�R?o���i��s6)��*<��7�S�j���W�C���%=w5Ɉ���kw]���-��|��(�kFj������/�≃�H�~La�����Xc���d�+�����½c,������G�E������É�Y���hw�9rQ���F��\㫏�g��|>�N�G��bXW�GG	�y���&{;��~�3;�<���	�O����wvFm����b�1d��,	��z�f.N������,�Z��K�`�0��ojR̼)zI*x!:���L�sK�N�B��CpzL�9=�m��P7���^s�]��~Ԋ���K~��%o�-��)�}�d���m��п������r����gZ��f�=�`�z�x�������~緤�z=�`��q�Ա�h��e>�Ohː�g�)cf����l�x7�s���YZ���g��'�Bۋ͞��t)�������yU� �i��]hy��͑�����#�p���Y�n�I]3�WE��t:׋�i�]�w�!<g���"S�ҏs�o
�]�NN���c����F,QU%��pj�{V�7[y����<٪8��_m�uc��~6b�zk����+�3��֣^o�r<7��5�0�/���ee��%�o���^��<�?d�k��'x�A���ʗ�鹛6�S�>M�C�nOP��[c=��O����|�k.�%x�]y��r]����m�=�)}d��j�b���c����1Ӓ)���%2rU���a���y٫�����z�����;������:����7W�w�#n�Ԝ�I?�>��s�xkjʼ�ϕRť�E���[��^q�}l5(�RUk��ӡ�b�k[G����~�x���K�qq�Om22=q�u��X��9�{r��
�"�s��%^4_�wN�4����X���9��.��8���7�ش�!�h;~����|^.��z,�m�vU�S<i �n7u�M��u�Qʜ�,j��黷�p�$|�G<37�<I}h7Ƀ��̡&f���c�k\�p�D�Zy�5�������?�񀞺�w���ΉA:���Z�(��8z����h��ܻ9�0=N����:Q�s��(�yT�j� :�#3����m�����������V4��2��!�U�'9��m���:��j	G�엚b���)u�nlLݹH�^���ȱ�.��_�̮�SӾ��/�B���b&l�	���M���9�4��Ζȋ��������8��w��ʖ��y�|<�SO���6n�\�1�/	r⓬��؇�U�v�e���,���/$�B��{�^nӷp�;�A��*��2a�2��f֬�":�&-R�Lr�7������1l�W�tԳ͓up��u�~���Y�,�>ma�i�:(y9�(b��/��������K<)�E:���n:�����{���R��T���NUs�;�kI�H������G#����YԷ�1�˔�f$�|�G�Wn?,�y��OLj{ͩ:�K9}�����t�v��������(H&k�f3�'�\\G�=�^UV��������I�1W�G~�m��@ᩣ<�ޤw{ٻ�K^	C�ʮ�����*z˿>ʦ�ZԊ�:�(Ș\cf�):�;WWV�{�Er�ٽ�p����v퐦�� ���������3L[��ا��/���sZ�eUp=���%�ؕ��*�#���f}�g6�y ���vw10�sC�U�3­r��*�o��dӠ�̙<{�]����hi��b��H�a"���Hgb�# �Y �p�4g�o{�͔���~�;Y?���>�^�%�<V��6�^��~llS|g(�7���:�*%&�.��o��9��I���Vϳ�B�S{��}^������5{�F;\�.�)�~���/m���v���|��:6���g��^<�;�e-,d���ѝ��^E�,�xZF�?Bʠ��O}hm��~I�)��Uܓ�ŐB>���c�]���~g3��rm6$0yR${[ˏ����x���z�[��i�7{��q���
À�f?ݤ{�GW{��>�^9^�~Jr�q�76v�֜����6���w\WNt�unE��qW��y���6�[�K���٤�/�����c�̾��h�-���r�,]�sf�Q*���W%{���(XUS�P��a���4�\�ͪ5&�x�[�R�%�y�o��j6�V$2�p�XNl`��b�!����
��GN���+�N��4���f�.����9p6�x��G^��8��jX=㋎��.�ݵ��8�P7�8�f���=�o�ǘ�;����7i6�ŧ�}�k�["�g�f�N������(5�zp}���#�+N�n��Oٚ/���%�t<�}4��\��:q��h^�+0�[��K���V>�-�=�hwB�)���j'R���~��nnI�>6����7߽��0[��*��/y�ֹs��-QB���Po��ܫ�FbV�'<35hBh����ڙC���^�יN�6z�RZ���B8c3���6E���^&N���h�������R��}F�z͘q��វ���io��}����-�˴'с]�q�������f+��{ү:%&Y�&�j+����.��yǋ�Vv=XV����y�j��|���5��ַg4�L�7�1����s/ek�<��.7t���z����<7ۉ`s¶�	=�<B�0׊c��N"u�6�ڕ9����֣ ��5H�l)���~�Д�������;	K�B��3G#�/�+���n�^�?H�
��ˆ����+���1��태�5+}=b��Q�o�N��sԱ����9U�U���qau��>~ur����/MgR����]��f��Ϝ������4[J�T�\/~�{�>������ �^����Z��p����ٚ�l���׈��F��x6Ж!��l�S�[���	�x��U绛Q�Z��=]a2�Z���ߩ��o�|��(+��S9�wmU� n����gK��7N��ST�n¥���]��nիl�p���-��ڠB�iڬ�la�9)
��+��.��u��Q5�!�Ǿ�7�h���)χR��i�����Y$���?+�=�L�}'5� P�)�j�����v� T�Qg:�isx�Vq�Gv�C��e�Ukd�M�6%�,�o�4Ӭ��8�*e�,���AD�{��X�3��3���7C����Q��n��fP�W#Fb:S�����qx"�d�\8�����(��ZVn�a��|"��\Y�nS���(v���Y"�:L٩5�y�/R푶�ZF�g'm̲Bʘ3����*ԅ|y]aoI��Fq�6j6�i�����:gn�vnܸ(*�El��gh�Ɩ9�cH2���4�:��ƘjΫїtѣ�}	ȿy�~x��@        L��Xy��b웍���#SP��s�j��*U��9]^��й6(��gf�
'�u6/M�	���YQ���H3y�*����47smҨ���N�t�K�:lE�cmvk8�V�"��YR0���M9���H7˞v��r5u�H�J���՚⬰�تc*1E��0 '�}hH�����v0LmV��49�
�[1JK�@��UiQ
\���n���MuǡUv��6��u�Q�,�ù��hܠS�RU��L"L��Dw�U�]����+�Cv1���Ԟ�w�l6�q�#�b�}��-��$�9�7�u�"%>�CU@Y��@�,@��Y�M�$���qn`t.��|��0�r!7LS��L4�������6���gr��м���8  o�s|�:|�̯3W�v��Y���D��i���dR�Qt�VQ�,. ��UQeU&�(�+TJ���E��()*�fZF�g i��$Ti�i(�JJ�����]�RRҹJ9���UV�+1T��`�(���PRҒ2��d���J�JDQb��"�D�L�]f�a��RJ�KbMUUU,\#u.����e1dJ�H�F��-/UXj�AEK�*�S����q�v�S7Z�=xiLxʾ��p�,N���k��.H�����\r;\�[5�}�2K(_�:��uu{���H��.ݖ~�&
7lQl"�W�o^��.Wx'WTK�8�H���S�4��uͿ��E!�վ��!Τ�*�1&����+Y�G��wQ�2n���9��1b���繯c��dmE0y{=G�M{��5���\h��^�g^�Sfc�$�op�$5&}���e��*����GD�&V]$r�{�X{oH�f{���7�U��M�� zӵ�spC�<�:���i�����/)f��م�\0g�(mc<)��̎�Რ�,þͭ����5U����;4MYa4�A�3�3��9�Z������M�w��Ɏ���'�����`��ǻa�=
q&8p]�;�f[��S^������a;yR��=��(}$�mK��������nN��q{�7��by4-Ɋ��������0]�k)�.ٹ+��w��~�JK)��>z��u8^x�n��g)��G=Sz�7�/MAtR�f�!fgw�g{��m2D�b��lE,Z�=[cõ�7\Պ�ܩ�M��f�R��j�.� "nޡ{'j��Y7rm�
�N��WwSz��8���+/N(E�~=0'�r2u�s���1�fӕ��Rfъ+{�ژ���t�������3*]��4��ƌo\�N�#f�Rͫ��[-;[t-9��̧bzY�>T�Up����{g%q�.v؋�yK�z"��{W��=��O1m{�&k�퐨�"h2�T�O�;��>�Scqfv/AT7r����<�mi��X7$%���	��]c��Xgv�Y��k.���{�ա	�z���=7<��B�9U�y��O�f�[�!�?o=�^~� dl��Wm�O"8�,iyk���o>=F��z͜������`΀*��Ї�t�����S���a䒵Ι���VH�����Vc�pU�o����9lAd�	�>9*�k�9L�G߀� RH��_���Ҋ��_.�
��"���-/O;�n�Z���^tY�
����S|�һm @�c��n�^�!^���Z�SǏ$���w�n���ĄKDf��q�O��R��G��e���=K-����M���&���P��+�=���҃�6w��5	q��K)��V7U|�NO=�C��R�������h�\"g���!�R�-�6���6��a��Ԕ%t�(�Թ+OZ���ž��ֽZ#1k!-�u��"ά�9�x��]��c���1Y�V9dI�T�CQf�8�􇺒5��ɓ2eX��be���!1[��j�c�f�~����1�W�;�P*��뷻�u�^9pﯫ�&��U�Wa�$��f���ջ:��'�˲�#SeK��z���^�6�6�x�(�~�6w�Q�M<X���ٽ{O[i��P���N��1oW��"dFkj���:�j�#V�r/�Km�k٨�fيc��w;o]�e��{*��Z��놽�qZ����=^7吵�K��y*7�mX���:n�邸��xpӳ���������f�]��8�P�g���kا@#k��j�̯��
Ԫ��:3`�|�5N͍���1�v3�]Z�E�['w1k�����֡G�P���2�E3g+o:\g��G�|>�����9M:�|���4�/w���+���RZӓ��Q���;��z�L�r��Ǥ�k2��j����	cz�MY]SI�J�)0v��2�U�`e������b��B�=��Z\�2��E�T-?^c"��S�����<�	��ē>N-	�Dx��K��#�2��`�I���i���p���T��r��2��|rPڼ�Ҭ�E<˻��������1�Qp�r�j�Yr�RL��Mg�I�\�cc|��ZW�����~f-c%�ݍ�t�*�Tˮ(W$5�^��W`Z4V���oD���1a�.�R�kXZhf�:�v:Ҕ��4
����#?���_��_�J��N1[�9LuB�:\����Ζo0l1I�|�)\3|�ė�v�Lc: 
�%,X<��+��%��\���2���D�Ӛ��$�5Qn(�������>>u3��R��'"����դ:<�7�vj�t*�0*$3�/�0g�xW�7ђ�C+(�{F�2��uaf �:�TlX�ڨ;�^�w���z��+EN����偳Z&� ��:,�����8�2�R�{�Q6�x�`6d���n~~|�k%�Q�$�r�us�ya\1�� ��f^5��.�=U�7�{�<�ym3k��/�t(��4e�d�����\{��]w"86nMC�$�MYu/{�m���	����È����W:5H����}��4��7��DD�p�Ң)��4�������k�k�r߳�� ������3t��
��=g!U��������Zc�|4ץV"x��E���S���jy;Բ�;�#��加���xY0{E{�k��N���ّ�P�V��j�DGD�64*�b����Ow{��>&���C&�q�����c6�*��T���ݭF�H��J�1X<j�/�*�Ufp�Y���:�� �wk�Ъ���]�E��S��j�е�N���ʝ�;]q�]	���
B�4b�����y�0�=���po�xk��`�0(w�בT�o�
Ѩ�{��`��k�%Uo:jݷ��B������;}]���Oeo'�V��R߲:�uf%�'4Yo�-}��ē/cu�˺��� ���̌�;m�Ҩz��/'�/{��yU"4�Q~u͹��t��5ᮉN-���4sq这�t�#T{|�ޛ���G�j"���R
~F���N>í@oȎJwR��Ƥ�W ��m.�@Z4�h�$S�Ue=��ɞ�;Sܐ�*��F�P� ��.xh��ؚ;�2���XTr�(d*j��*LX ��{�Ϋ��W7�(�׵�#�v�_ʺZ"J�|8h� @�l�5 �������}�~T�K�u~T����:B��͞|6q�S�]v$�]N���l��EYζ�!L!Oܫ!�q�`S�$;&i�}*_o�z��j
�� mW��O�	����Z=)�.�0W����9��5�o��x���M�so,un�j<a] ���<��^ዝ��-c_���G����U���&m�e�c釣k��<yy�|(7~66����]���񡢬��Hp��x.�<�YOwfM�ct��5�]�z��*�{F�~#MZ+h����`���N	�*u^�5=n�'�
�t�|Lϋvkr��K�;��������c����,�O"����=�c6�A.�!����a�2�Q����o�pW�`]ui3)����O�1"�tp� 
�Sڧ�e��Q�3}=W�/�OU�]�u�<M]qо4`�壬�S S�,��,o�vl�u*3�U�i��@U��4�kQ�:;�O����{z�	fV8p��x�CEd&�<��FR^S2{z���Z���z�^<8V�i���.����QB:�:i<M��T���c��5�s��˶�e�ne����
�����thj�M����jK�;'c"pY�^s���.i7�̀�C�x�-�*n�cmf�S�쀞�ァ�����m�r	k��֨��@蚁�S-��
��|�8aD�v��.�{7��o^����3�44r|f_b�P�7�F^�7�e�U�pF8�*�-�7|
-� vQh��CƲ��H�
X��ϯeb�A^�uup�U�:�e�g%�{96TJ�Ov�M8ò&���/v��՛��/X���r[2宄+r5�C�e
��(�6�G���8A�۾���`�F�n�]�ͺMh����MA�q^1���ٴ���[�S�����7���U��i����'EժYoǛ���e^���v�[CW�M[S���  �  @  OS_m���VKƸ��c[�g"y��kke�u}|�jc���]��f��h_�Q�ݦ�:�5M��1�א�ك�Sr�!�����榝��]g���.�����p3���t��ۊ�R��N���7K:A܅G��J�Y���r�lu�f�#5�YW&��{�~�b���l'�w涠���3Kݔ�#��L�y�˾Ag�u����k8�q$*�ˆ��G��V��s1�f2�ͻ� o/L�}0&\��B�����\;҈�1S�cxy*��a�;�C�#�7�u����.���˾[�E�r�=Dҽ���S�/l3ұ�FR捴��jIvV�.�(�5�D饫s�Y�5��ư�1���dna<���� *��  ;x ���z���K�Rb�r��*���h\�m���R�n�f.��1n��JB�e��+IL+5�\UB����6[e��)-Ņ�Im⩤c1Y�����]b��m���SXH�1X���(��ӛ,�*��5��)�3T����1XT��*�%��!U@������h�]Ue%&3v�2�UU"����]L1{��L3	S^c�gF���Z���-Ei)�))�KUm--*��P�ʩԤ���9���񦪀�n��}_���풱�x�q���pL�w�-��~�u|#�%�%ֶ���<�5$�=.�wS.ߧ�n�-O=�:�d����#��3�:�m&i�(��]����O"2)
������^�4Pv�F�����ɽ��H�G��U(��Mu�
)����9j��1�D�G=OG��Z��]|���S�Yty|��G�MI��/�'���L,_����G
=�5a �V}v;ƯN�\#���r3��8=��b����
|~-pu8*^����������:X�G����AP-�U�_&�T��-�wE\ �j��&r�ǅ��Y�x��^"×�듽N��&� ɧ�B1A��U�
�3�7y˔9�wz�u·�'��d�� :?��l��䆇K��.��������j\��E<�p�%i�]���� ���|n�Zًd�{|\�*�r2�c��n"E5p��;*��r��ݥr�U����f��vțpcT;����蹀t��,�UJ��޼5;�^D���������Sب��a
�!#��q^��^{�Ү��~�,��2�.��+F�Ѵ+S)9;��Z���
�h�O��ȳbuǇx��`a1���QEᠫ��'�F]ңs%��b��!�V��$�/��k�����r�\@�U��X�2)e2t�f�+-n���ʥ��L<d3�#���C�-ZU*Əۋ�I�>���=��������E���X�a��7�3�l�~�t��\Pz=f����tkiS7�~;=^�ʑ�TVM�Wꇃ&�1[�Z�<M!��e��[�h��+����ꕵ�4O^5�o����IVƙY�U�m٨�3����ȳ؜��t�fry������
�lV�fL�&e���r��v6�����}��O�5�q�tѳ�v�����
����d�}sޥ���<>�V���U*��۪��Z�P<��!(�}�9���8��W`~�@���#jm���^3V!�;���܁�R��-��Jܿ��
�PK��T+l�\���9%Z�<4y��K�Gi�<+Ã�h�%�RU��!�����ߓD;D)�/׌S��x>��i����k�ُ��mzy<H����(|�*�Y氚vH�4����vN����dG��e��5T ���m.uj�?#L!�x�}[t/J�2V���PA�.�Uj��u�OZC��mA�2p�͜���[�#B�-(�qV�PM�YC�#G�yC=~uC2.�ʢc��\鲭��ԩ��QR�5�]��i��sњ񕖢�]�oy$e��n�u��-	r4��ԓ���o~7�����&�u)����$U�+(]��˨��w��X������oƀʜ��X� �4-���m(y>��wM���1]O
7�
�Ck(o���Ô��&�H���߭� p�Y����<0p��]q��'�)ğ@Fm��z����0f�מ�HY@���H��;��uOK���M$]a�)W�N��Ɏ�=�E�4��+$��غI���7{�����Ҽ�n�C�V+qb3)՞.{zt�~�j�f�� 񗊼����ƽ���Suq�hg,��܈}}q�)eM2۶�w�%z_S������9d>|Q�	��o��+��ڹw�۵M&;��ƾo-�7O���o0�^s]ҙ��-��8��>�w�5C��+s��
0���Wo���ա��/h�[�i�U����]P\��?�;�}M�{�
ў9��$`�k�D�F���~�����ӝ[{������������,��T��� ��iV��\��!�wL�	<:����Q�Å` �6h�+.�"������d���Uג��(p��NXu0XU���U�#�y6MW�Pw(���-
�+�:4>v�B~S<s�:�bi#a��>g=-dZ���~vsw�\[%t���jhp� -#����h��QWƕ���˚}툨���jᔹ�n8�T�d��κ��e�����C�c��[o7{i#�ܪ©��� �d��fS^z���$�dnɪ��U�9�u�� �����~�k��o�;�˪�Жw":��=F��차"f�3_W ٬��JYk��E���iu���u����_�B>��f���e�!/�ǚ�->���)�x� x|h�U������"�Yˬߢ�Z�����]��/:Z@���u�+k��j��~��XtIs�ë7I~ ��}Xh�V dӇB��L��Ӷ��}���M��e3U�NF�v�� @��@�~H@��kӞ�Ssf�u�q�Oب�6 ��:4B~_�ڣ=l�˺z0AՎ���}u,y�R���>�`b�M$DR�~�܀��xQ� U�k�n��V�D���Qka�1c��L_�ƌ�.�?m�-��t�UY���C��o����{j4�q�!٨�^�ULGQUdq�/>nwM��괫� ��DT�(�����j�³M8����8�0�t��#�o�������{մǲ���Ǔ*)Mv��2//ޡ}15���c6�s��ĝk�0ߒ�.;� �΀�ӧ0fe'y$o�|9ƚs�_�nX*�������^�K�h񭸼 ���#�ҷ���١���l�u��w�9-���-Wr^֪�r:������
f��Vd@Dt@Əf��gU�j��nwp��wk�M��52��-�l�䩎 ��ǻVw׾�&U��pl���xl�p��cP���e�DYPw��R������T�e�5�t[��{�ה�'W�ؾ9L3֫��� �򬰠
 CS{�K�����&O5�wUx��u����J�L��{2����7����Ы�[���U�G������˃��xW�������y��)wK¬xP4�]г�� h�S7�g�L�y����yY��=��*��j�G�B��\f����U���9�'	S����PΖ1��%�g.J�Jwok	:\g{���-��ﻉj?-_���
˩J�e?�*�k?-2i�h�XQY�}��]^Ӿ>�ƹ}9� �>Oz� �0'�={��N��H�Xk}�
U�Zh�j����|3i{�۬������4�SƴZ(Q�GF��EA6�[:��J�Q�+s��׳�>��Odz(���4	N��E]S��{ڭa�z3T�Q�E+7���k��~4�S��t�h
�u����;X=<�R�
v���AxԐ���.���;<��E�s�+����W�_��h��Y_^V�N�:�{1'���9�x7&AC��.r�8�Z)��h�����SCE�u�i����T!�;>��6,eo�$���(ѺԱ�g�X/-�p��mN��.� ����t,�1Y.7u�����h:��G��u��JnvS��4o+R�ņ�v]V���:$m�t��v�,:�h�uY}RZ�M�[��!�~�:G��1/zG{[ﴛ4K�[�Hh ��e����G��^�=6��}��Οg1����U�j#�0WpW-�x��1X�Ot�v`PU;�dטP��7� U��j��\�]<��UM/a����ʨ(i"�
>ȡ���/����+���n�������Q~u��G���t@>9�i�5����{ӽ�K��|,A~5ٴU`����.�!*�����wp���&�j�4~��5�����>}���&1�����ܪǷ�>��ᑫf��Yr�C��j��ͽ}~={�6�'Exz��dD{E�W�1�O�.kR��[�kR�]����7B]Z/�q.G�cu�98�����uAX7^�أ���z\ܴ��6�hh�d��z��v���u.������I,�o]�����-o9���MH�go��T��|	��V�7��m�z� �Cc!��o��<�:��Q��8�+����x�Ȇ#\S��X�@��օAɏ��
�#ѭ�f����x��?�\�^U���QbB��5���G��A�iըsTY� xS���xh~�+"����-�^�{Ϸwi��1VZ� g��� `���ǅ�b���Y.�b��;�8�u�;(��9��� 2k��F� ˏݻf^㸣�aF�w�k��c�t:ź5T M T�^�u��=��X8<=��p��D1�*���A�|���ˬh^����.��u'i��p�2��Nӫi�Ә���HjAj��燊��_��Y�͘�X*�����������iEO����I���
s#�ZaMX�m�؆ZK`�B��`Ck����5I�j�W�l��e�6�qI���)��kօ���Mh׸�&��!tn���)�agZ�$�4]�%0Λ��5/n���t'��	%�� Ye����1n���;]:E��3:���?e���=�Vh�����'o�G������+�`��D��U\�:��P;vƉS�V�gX{y�O�ţ�w�d��WI�#��j�ŷ��K:1GVd��r�]+Ń��k��^\g�\�h�z����&Í����PFLVÝG�N[�9��ܥ׆^bɠ�R���E2ѷӌcm�^qޛ!��̓f\dxz�NG���ժ[Ǩ�5YL��Wjr��Ec7vs�9	����[���!         O]�C[^5o�kl�|4�#kr�^��m�w��˫��"�P5��p�>���릓�7 ��'1�ͼ��S.r�|G��-��v�!`�[x���E�1�W\�Y��;�3DѨ�L������,>w*P�ݥ�����.7�0¶����515j�5(���v���q|�����5H�Wo�7f<;E�7���f�ՠ��Z���V�����fM �,=�UBBf��^�]��p�&
�.���0������G3�Jx�6Ub�*q�ື)��`j�j�|�i��#+�c��n�s	����;Z�x������a���tC3�)Hrs`��A&�m[벮�{�ȟGEi>2�I�.ZVs�R���B�tngQ�7�I�l�p  ��ݼ�ٟ����Rq�Sb�s+�H��M��*b�w�]���"7T��/	qn�	WE9���-y�q����J*�ZWVSV�X���S�TAe�1E���ZZ����/b�*�X�9�b"�	H��9IL�^�
(�a�Ċ����D�*]������[U�)��T
�Jj1m����噩��c�P�
��U~?�J�5��"��cxe\�h�"��Տ玥�&io�Ǡ:�Js������ �eC����<�l��u^�z�j�Eh����2G�<��͡Pux��U*�D���!Z1U?L7f�k�h��}���Q8 #�����9 �Q<)bULG�>�:]׻�̞�pA�*\@�h��"�Q�Z�^���B2���*��b�g��\q��Lw�����Vx���zl0��5���s5�il��ZWʗ�����Z_M���ӽ�am{M��;��W���C]Z��t>�@Q�Z�Z�����=�8{L`	qg�&���BiW���H�߀���[��/o�J��h��
��B	�����>5��p��gk��~F/�s�x$�KT�V�o�W�E�ɭ\�L�v|�#��L�qx&&�@>����� ���[��x/r�8=y�C&��	�����{Q�z��@��N�-3휟ټ	�+�:[�F|�6��M��ݟX�U0�Z��DO�`��(�]��~��f�ez�M���.b���X*N-��O�X��ӵ���|hJ��.�T~L��������vq�bq�R�X2=V=��w3�ꚴ�����=:�rI3�l6Ly^L<���FQ���U��g�2i��m�x=o&����T��ºNt� ��ĸyڠ%��
��m:��3	v<�μ��4V�� T��ty7�ӻ{�Q�:�:�f���Įt�MXt,n��zߧu<�^1�'�Nd�^��^�F�� &6Mw+�����}�
xF5hӲ�LƸ/W�@N4sʻ�����M�=��v��e��d�r&t��*
w�j�DvޞXe"��!v)��V�Vf�M�ٔ'��.X���I�g7U�1�xKJ����M�"�>��?}U_���X^:C+M�ʵ[.P#�>y�6����է�q�**��@@�|0p5}o�����D׬��@T�YӴ�ww��z ޭU4�x�B���eҷ�*�d�~?*�ޑi���m��N�U�گ;��aP���T6�:kf!YϺE���u,W�JVRCn�aw�	r�q�y��;w��xg�c��&n�C����R T����#�e�K>K({�OԮ�K���;�R�)���8h᧕y�Q���qbC]@vx����:ܷ,�r�����S�����P��,͝�O7PMT�\*Ӣ��'�t��P��p�¶�F\�N؃ꋅXdզ�!�~K9��� ��3Wt��之ҩS�XsF<u�K`o7�F1[ɗ�^j>��M��v������9��ɧ�7"�k. �ڪ�5��ޒ��b�K���ӿ��;;���\TCo�I�W�5�ӎ>0k�觠�=��}�W��Aa��J��Q�eS����X�U�ÎWJL.~�����U�&֐�Z��^
�*��L1�|�kT�'Rhw�Ep�F�D0�|�b��*�7�P���ûy=���M5����F���4Y�k��ʝ���\��w'�q=��vlk����A��λm^	�K�/�^�wN���U�V4y�;�1�P+E�ۯLU��wx���ןD5�)�(�.
��Pm���.ƣ���ŏgI�����4V*��a�8������`��Ou(��lU���^J�, E�a�0vypc�6�����9I\�tcF��_tz�6�b�yn����$:��Z�sn�-d͘�쭝�ћ�P<%	�]�9NopԐ=���f��rI�>���an��l�����
���wxd�F�u��D�q~��b `��7��¯8t|�
� &�Ç:��y�Խ\��a��>����U�� ����
��^N/�US�p*4k9�'��l�<^=e(N�+Grx�;;������v���=Y�jƚ�@�u�gVx[��B�"�A��U*����/�h��0,ݘ8+�۲�ӽմ�d5�|*qf� xRĪ��9/y���`����8<0��+B�B&�VFE*�<�Z��e �5C�w��©��4U�2��Y����8TK��X!���@g���5�x�X�Ʊh!_*�U������2��l��yz��:��9R�n�#�u���tv�Q{Jf�\^�<�Ymͪ ��<�z�7�x�o2�s^�̧�4��>d�=��4��طN����_��v��X�!{�����6���X�xXb�8ޟY��+����PWU��ߕ��6m7L1�����>��S<J�k�*ǅ*,���8��S�j��V�F���6*i�������l�&���Y��<�.���VO;�yl6nN�-j/a���~5�_�����䒈��i?5h	��,���UF��UXf�B���:2��Dv�}�B���*Pu����I�Ur;u)��l97Iʍ�ں�F沌5K��G:�X5�(q�6�B!�5�dLc~�������ˢ��j�m���X�`��@�}w4���Y���j���t�+�s� ׵xDO_�����#Q5��g�2�
)���wWZx�ŏ��%`����X�z�o|��L�iIyZ�q�e��n��y|LOo��Uitd/$�w��E$�;[AW�_���	a�3(b�A�u������y֋���-z�����b���,J�yC B�=XAA����!�o{�k+҃@\����e����>U\ �4Z���_�g��`@z*+CmJ�G������	Ə����KP�=� �*��J��P�ZlvU��},a�C̠�;t���0������q|tX�j���#������xn�*��S�����bT�NH�ڡ(��N4i^x}����R��At�}4e5��u�ڧ�2�C�jv1CQ�龌���Nz����
�aP���W�d+�{s�ƕ�xS�2�=���\��齶w.�<Ls�\�n�^f�>��YZ��+sw�Zg�� �3�=��͍}�]D@R�J�(Wv�,؍E�1B���]N=�9ɭwc�<�X�uP�P��y�گs�ľθ�S4����|QO��~S���v�o��%��h�,�e�jy�|�:#��O�I�x��vkC��j��Wq���`��������M�,:[=���^����+,�IXt�ᡢ}7;db<���2��˥wt��S����*-]kwX�-x�M�S�ziW��|���(Y�T�j��S�ly�'�Ľ���	�AC�RU��g�*dYz~���U6z��>ܹ���N5�ʨ�	���&�t������]_�7�r�~�㢼 �3Q���n�@�oέx�zj��׷M{�(Y� �F�5TD��x4�:����oުg��fǜ\ �^G�+�O*�h����S�n�a�L�c}����Աd��%������r����n�o�fdv̈�/R��p��vI��\Fv�܌�x���fC�m�v"G�:t7�{��r�#na����
�jƈ��Ll��5��̕ᛥ��~��Չ.W���t2�ҡЫ50���,���39I鵑���xA�@�Kh��!�8��t��^t�c�}v��Ԋ�h���yXa�N~\�=/5ν�Q�(z��Bq���&xpU�V,�ѠC��^pm{���:�y��aVҥ<t1C����Ό� ���>��7�m�+p���0��q��_3@�{x�eS��^#�q���.Fc7;c����XN;&�*��	e�=C�ѣ/��TKH�t����D(@��W�
����,�+EK��Z�1/c�=F��#�k�5T�@�_@�h��0,�������51��j̀�\�(=�o�!voBT��wX4j�-�.�m<�"�)dn�ҝO����r��p��$ea$���	��	����J;�Nϼ޺3M�8�t6K���Q.��x�Brf� \)���V�?d��c��(�z:�)�u,�@�i�Ee#AO`��_NݗW�X.�1Z����xp�i�l��q��{ۘl��ih���*	��uC�?b�E�#�TӬ��{�~��\X�X<=���τk4�t}ʕ!��ۙ=��`w��Y�����,���!КU�b��|��H�Z�:M�Z=�Sg���e��pC��k�C`�yUi����_97k��*���K9{��M>R�\.�T4V�>#�5e�wv�:9��N�H�W>�-�\�z�lw��k(�B�}���
 C[�����p���X.��r���KQn��r�|n�.�iޓ�z���^�"Jΰﴌ����1�ʪ�rt�����k��(��K��Ś�À'|"Vq� #���h㴆����,vk�W�u��5Nb�<���33)��L�gK��	�A�z��;�������=���&��%��N#�F�MNwc�l�G/�L%�|��`1%�skOi�E'YLK;No��.?���E)<Rpry.����+�������Q9����Q2Ь�/�9�%�+a�e�̽kqK��b9�(Z,��y�]�� U�D���僓�IΤ��a�k�-��7}F?�=9CJ��%\H�y��x�Ϊ\\��#���q �
r�r�
Pe,pQf���d�͓#�{���uUJ����s���\���J�x)�"��J�n�����w���w�.��s����L��
7U�.�u���U�>ݝݳ���I        ��c�M��t&�S�#�S'77]֭P��[�բ<�]f���.�qҡ��zEޙ:�֋V%�њrug��,R����"z�E$�ݽ�F��Õ���;P��Uϑ��U&��2'V\4����.&�7{�	Nb�����H� ]/:�;��;Y|����jmp�v���X�Է[	���qAt�1'���	�#�T������%���-tRp��w���uK��Y�z:�4�_"
:Vf��w�;��1G|st��f��Ȕ.S{_��6v.�2U��cZ�T��1�Lp�rF�ܬ������㐭-������֭�Aۢ�1���Q���lvWqj�1a�0��⣴� �۴^�1�\�n���hM�gfop7�  �q����%ܣ-AUT���[J-4�Ui-GC��n��T�UQcm
]�T5Fh��a���R�W��T�*�ڪ՗�L���Di�K��uv��JV��U,U�[%�����Ŕ(�B��l�Ab�(��0��V]-Ae4*��P��liUUDb�ն�P1�1�.�H�QT�(���T�10�����% ��1Q�R��!L�2Ѫ)i�"�U
�hR1`�DTEi����UU�y�o��3�g^j�W|�W���A��vt��3�Uqu�F�kcM>�q%��C^���b�Ɗ�I�k����u��'����)�[�'ݾ�=j��X��b��V�H���@�|���˻�:��j�g�V3��E�G�����_�L#<��{㸀��/ƴg�P�]u9҄ =��T�}��M��!z* ��0��"�K�t
��ذ^U
[���7;���5��+:8pr�yQ�@��2�0�*�j�_��5����u�mR_I�-4L���8h�z[�����#�)�D��z�Ʊv]i����~.��"=X�Z�i�{ke�t�x�E��b��WB�q��U�]u�:�t�z�xj��㢸J���@���חc�upZ���	{���6������1��J�)�d>�͉�n�s�B�-:��n^�t�
��f뫉�A���L:��ٕ	�\��/��54㍪��m*4�0p~���䫣�>�V�58ҴZ�]����OwX���u����=F�4e
�x�5KE���F��mt�&(��g���Eg�X�cX5�h��yU�g�����Ѧ�z_���6w�J�&��-ڵu�hؕ�V��F�I�~�u�՝0Et��h��{R��к�yS���I��>�U���V�t��0h�4ћ[��r��}<|����bP2��ы+Ua�GC� � [�{��7�	PeI�w��W��&��A�����p��~xE苒T<���J�5�xX�ϳʺ]G�
�@~����n���xp��F�<���t`ڮ�ן`��g�ҟ�
�Y-��yZeq��
�4hPm��v�c/�l�-*����F���S�\Q�j��f;[�5��ٍutt�*��]�m�<�'4���O�7������*5��T>�h�3�B���_/
�\�ή����}d�t�wǽ�b�C������;{ۉ�u^�8Pv�G @4ɪ�%��"�~=����2�=���1�c��h��za3�~�r�#u�*� ]W�b�c���&�Y�Z��4���5�� �56�ӽ�6t]�Sի�W�X�S'E��*�U2o/)j �0���Y�~���!���xA��'@
�h�U�׎��^��_9���f�u��>g:*��^-U�$�+m٩����g)�4i
�T<�"�W��a� )]�Y�(���^��5ƚ����;�ԡW���Cd��,m{��=�Ĭ(ԃ�}�;�B�b-N��J�K+>�ʥ�ѝ�oKս3e	��D~� $��y/>���	q���V%�h"e����<��WA�\vv��-��1���v>�c�]���뤾f�
���T�Y3���);W���p� pf�_�AK���ʼ�xT�U����O^��2:Ƹ�� �����갴���$d�2vj��T2����EpѢMT����X���:K̏3=��ޤ!�0`�����C��U�?)uD��U��Jz�GP�̖cz'¸j�0ҫ#�q���
��+."�ʸ$�.h ��7-�	�桱��4�a��h�Æi������'N�=Z��W��Z4���LT^-����-_��3�z��v� <~
*�j��Ȧ��(�M�6%��Z�sd�ZV`�WZ@b>�b��+ M9��x�t*�dʝ�=KRkK�"��i����������1λWc[(k�Q��Xt]r[2�d��*�!+'D�Gdp7\�4]&�jm'U�r��ӝ&I��}��lާ���
%L~2�Y�8pL�,W�����S��g��d�k���UhV`�R�<��b����|>��+�w��9�^���Z*���}�<S�W��.,�u�W��wG����� q���(@�<7j�h��Y�2w�,����C~��0:�C�r��vf�+8�Gi���WSؕn�j���Q]���aF�4��+�X5�(�^�@���|(Dy��n��o���������h~zE���uB��w�p�&�b��?Q��L�vHќk�q����r�Π w������0>�,�PSp�]e���=�C�A��B��}ș$D
��PW��7�Y����7ƽ��2���O�sվ�e��pn&�-]���v��"ĝz �7.s�ӗ�͵^񮩙쓺Of�z����к�U"�.�Y��X�w܎��ֻ�w=�8���J��yS��X�E��m�g߷;[ڏWCDW��=\�%�VbI�����i� X@���N��g�~u���fI59��u3��4&�Ӳw~�Zy(e��p�Y���������of���"+�+���<3�U���e:������f.�5�5!�c��Nmh6jW��y{b�(c�O_
�n,�[�fon`"H����.S����d��^�/A^ýh7zФf�vN�}�ua炥�7ş*�Q�.�f�Du��9��Bi��ˆI�]L�{1�	�Y5w� C!��0k�ի7��]h�T�>
�W�҂�P$_�� @�j[�\�l�e^�l�c�B�:*��=9�UZ*�7�� JhUU߽�k6��V��}�k��[�aF0�n�h$il�8��� ��F���<+/N�z*0�B�1_u��<8�K�$i~�܏6��̧v	-��^��-�Po�5�n���3�}�I��&F��G3�LmU��pT;�9V�r����l��R]�r�gvX��o�l410�.�5�|t��M���B���ݭǼ`�CEM&��<"J��5)�f����*�s��z������P9�4T h�i
D�s:G�Cݞ��)\�Z&^x_���z����WS��-z�y�6�1��i�&��U
�
���!��"D�lz�����*@q��U�Q�����ǡ�{dv�eR��?Dh��*�v�6���~�|�|o����:,�V�w�1Hn��涡�I=@V���5�b�k�xa5=
Ɨ*�y��G��Z�y����bW~��(��r�sѶ���������o�y9�(Ў�Τ�G�h�)��y�]xd�̃r�7$0\�����յ��rV���umEpu|/��D��|(�Z5Ĺ�K��V��e}��y��7�U�tW�+~�Ն8:>��w[x�I��C�Wg��v|	�[5{��j�%���*�k<��A_{x�wg�ԼB\Ki����8�^����:��n;����'8�5����|)��tt�7��}���P��*'B4j���g!T9��S��DCKcp+�\6U��3��0,5��D)ȅB��(���<����&������]_�{�c�)e��T��:&��H�\+C�\!r* ���[�����[�J7���R:xu��8��ȍ
�F�>�>s��\����X��,ՁǇ�*_i�(t"k{B<��픞�������^��F̗�jk'Ym���`V���櫙2I�,�͊{��9w��K�[p�z�V�Rܸ�ƚ�e6\�Wvk(6L5�x~2����)� �T�1r���v�w�2AuJ+��r�a�d��w˅!Z'�f�P��Z2z����<�s\<)�,[�Xo�`��~�N*��d'�i�����=�CW5�C3� ܮS&��â��jf�>+�0��@��K���]��9�mp��-PD�i��e�t�ƅqx������<>�<���[��i��EDܿM�UX�i�Y�B-Ţ�U�){Uk�{x8Cf�=ks&�!��0㪧���������5cB��Kn��}X�C<|+�Z�.W҄����w��+�&�aԛd�s�ζ�'���!�g��=�R�����B����K�G�q�rHX��bv�L��s�i�����_'�᝾���,�XܼG.�j=܎#|mQ�vB�)�8(�!%��V��:[�F"I������_�c8㬯�xڪL�g�_^ܳ�P�D�֤�����q�
�h
L�����ts(.5ʪs 7J���Lr�;��j'_.g�\3��j�!�p�j�o�F�:*{Є��z�{�W��
U4-%�ip�>�U�P���r����;R����:��{��J2�Ga��-[�u��z��}ؖ��>s��\��Q�P�ȑ *^!�DR�x`kʞB�������;ջ��*NTUg���\�����6i�~�/�8���n��=��n^��V ��N4i�w�< ��3������-��=��=C�v����ùqS.�������FV����Z7����Ox�p�.��n��*W�b��U
��ӣJ�:�O2��ݢ�TH�i�k�&�t�=Ǚ]Z��,e�#�`J+Oe�]_i9�:�2o3��m�.��:�N�B5p�u%�\d�����޶��^U�H�PI����b�֡�f�� ޸��8�QaX�Dd�1��.�����nTκj��/�)VOn�E����]�A��Wf�t�h,.�:SV��_^�i����(J�vy�Ѹr��\E��qg9�r�n�h҆
�/��TEҲ�-�s o:��,Y<�3����i�{��'����=ѼjAAA�N�����\nL���\"]֖P
����\w�"�^9jp��T�\��]De���r���(ږ6�[n����Y4�V����o ��VL��j�N���ՄA؂���,�;$�k�����e�L��I����w���Sy��         �ms�W<���[M�6F����
�z�F��ljy���/*�-k_.Fv.�J�C	9��r��\%�&�p�x�-��/@�ב9ޕqb;�u�wD �˰���Ɋ����q��(�.I�p<�W5Z�B���7��Z�`!��NSI�.,�c�♇ǩs�8�n�bі����\�밸%�n(F�
�j�f�Hes�V�2��|�r�X���2�M�i��{.iz�"�]^�]0�9*����:�Ň��u�A}Ǹ�*^��u�ѝ���uB��#%��Z�V�f�����&��O��9�/�(���	�����g>�P���4e��έmd�=�lil,�fB�մ�}�����/�N��1�Ki����=#<]���x   v����<�vw"��Y*��)IH�TR��>T�Q�)K�%��B��*�X1e�8qdX59r[ba��))�e�DJ�cZj*��JV%S���
��YH��)Q��$��dDX,(�CL(EG�J��7wH�"��U�(
-U[.餩TWR�*�TV.h�"�*���X��J
�*�0R.*���HJTb�)��X�e2�FA`"�"�,\�t�R�AHSb�0��Xb�1T(�*�^j�\U5ALR)2�EYuRЫ*�"#�-Y#���K��#�E(��(�Z�C
��R�R,�AdY8JF�DE�((�+�]�yޮ����
ݟM���l�p�1̸/B$�*k&��X��.n���$§�v����	O�����ʀ��g���dp7��*m��lҼ�kpm���7b��	�)Wr�8�K�|:�˞�_���u���h�|k��
'��^:<���϶���P��ibC��t��7��4ը�D�(�3.�o�=��O�;���
�L~8����5ڗ���V�:Z�V��I0�`�ר��ϯ�8v���c< �?*Yζ]��:K��ݫ0�
��P� Zrh�#���>�]�c�v�b�hۏf�bT��Â�(�F��O���3�S�����}7�q�@�P;Y��]B,:�- `�P�y�*�JC�+�o���^��C��C���/�.��ׇQ:';"��/K�YO��WT-n���ZRa.���^�*�7���Jn�[�b�ŉ���5i��+���X��\�5�����-͘
�Gn�;nHK�&�}#sgp��Y�B�
4�PV(@����Wt�<�+
ze�}�"���^�v �T�ׁ6Zaٱ��9Qp��O��z��f,�GO9�i��.��6�8���|ȗ��͹JZ��0���@׮;��
C�}��`5%yo�&�Σ�L���v7٫(�eF�������c.����P�Z#��)�74.�k �o1,C�P�8���q��C^{Z�	�0+� j��7wtQ�*��m	fPT��X�z�]��oc��,�d�:L���j�: �j�0w�U�fܳ�5��/N]'�:����Y�/A�Z�$ <`�𥶴*g�G��5������x��U^Q:5q��ht*�h%��2��S�2�0燻�C2m��f�E���7�ʬyH2eta�tA�$��[�OW+al�9�j�m2�a;��
�;w�u��4Vn�ҽrI�8�>n��]��o�M��k�/.������нl��R+���=������+ώx�4F�j� :**�,�����C�,1�|H��:<�SN��N@�iy�)޽���"ǉ��<�7H�Lxxp�&���Z:&b[s��W��I��v���T�gEЯ���ʍY��f�p̋�=ﰏq�K"��YhӾZ+)���W�(|�yy���ϏI �W]� w��a����������Z:
v��zf��U�vX�Y��ᢸ0� ��adׅ^ԝ��9��-�D�S�b5�<+	z���X�E��X.����{{]!ǖ�� �6<,`�nr��d=g���1�k�3�d��ԃ�'mIK�ο<�va�4���ָ�\��u3R�q�奚q=Z�(xv�5gBl͵�Js�Iq�37�=�iE��hoo�򥜒H΃�}D-#����Vt�
^����a�Ւ�+,G$َ���gُ��w`���וY�%3b^?J�&��6����U^�������
�q����Ea�ݫ[�ro<"��%v<���	�\�O,*�dU��V:����
x{C�`�J��~5P��p�FBBK�����{�t����ƴV�ZM]u:�\ѣ-K��m�|ö�h��*���=�G�� 4�x��hF�+D������X2���G1�7T ��S>���KGG�o���J��/M{(�gFɼA���ORB�����´]oR�B 6=o�ո/���Ԓ��{����#�z���,RV!ֈ� K��2E�}qu#�{]�o���|�r�[��X��-��=���؏d>}��3��d��GO��+-�:Q����ֺ�αc5ӈ̒G��>��r8�`��w�� �о\,V�L��Db��l�4j
�>�̧�%��"��[@�3�%��)t;+��W�����^��f�U�k=��Op�j�:�hU�2W������s��s����ۧ_X��e�pa�Q �W��\���i��k���f�n�*T������_.|fQ��N�����4I���㴮��0ץ8��(T�V�&�Wi��Y��������
��JA߫�x�P"�۴B�5�Ec[V�7{�7����*kh*R��J�yhtU�� �^���B^�W����.�x��ԄiV
�=�S��B��·�7��V8�ʘ� ��u�G�-
���Uyծ�~���4ʄ�p��J��[�5��9�Φ�
x�\�>�{p�Q/m�Rg5q�u���l�gs���rಹ�%.8�o8��I�¬yY��(yX�hP��U5a�x���Qޅ��'��w�Y����t4 ��thT4VBhz�+����z1��5�w��PU���	�����׊+G�5 ��7�K�{���M�>S�J�X�_�c�`uR�W  �H.	NXV���{�܀�<��.	�t���IZh�Pxp��F��9�8��=��;^��8*^�G0԰O��i���;��_�v�\��X�p�/Ulh�W\o:�UƩ���De��/*P��;�mwֈ�h�b+�<�K)u@��t6�\{ٜ��+ޟ>���B�G�.��G9pw�Rg�Q:,����!g����>�u�Y_YY��.9t�+b�=l;�mU��Һ��܀��:���c��X��S�9\9IE=b���}�PuiQ��T&.�Փ!�-h�DNs�xu�\D���E��yy#x��Ȯ�Ȣ�#i�#�WW�kʵp_8�;0mV|��E�|)�CW\�`1;Y{��t��>'�҂�������t���`�����οg��ǰ�W��$
>;ŞU���PxxRgG���V�*�a=.����������_1@��\��yz̨.vx���]���,�r��Xo�/.��!X"kEH�xz;��n�}���4�°|���j�U�B��B ˷m)��_{�l�c¬D�:Lر�q��*��z�Xr���dDϴ��7"u^��O���+��j���ÆQ5�@�
�n��˚�{M��V]��On�#�"����=D~�c�9�w��a��@�ҫ"�Q�2�v��T����r�{WR���s�]�7
ШJ��VҾN���������M�uY�#�*G�d��	T4�N^<���A��ޑr(�ot10�W�WY�WgEd5���-�À�/��vYX��(��+����e�ds�k�\�.P�׻��5�z?t?L���Rnfu�噕{�
���k+z�[�U�>��T�U�|�SͿo��ʁ�0��o�����^^���oާ�[��.K`���u����ŷ���<F�K�
WXCu�=�8ߢ�M.��c%��2�^�M{���}�yH�'��
'k����-ƹ�5G��Ԏڵ��$;ͧl't���{o�há�꺨˯���%]�Va���H=��=]�6��r��3���R�4���ߏ�7��z�X�'J�vaϺ�d�Z��qU��=r�	��'���y�߽)�����gE���~�v-�D�/I|��U*��w���'ֆ氈��L���^�0H7H�/r�ڗhnQ��������xy1˕,#۟^�F�;|O�M�90;��P���'i��+��z`�Op��;�8^�����K�Rd�/�/�/��S8J�i��6j�d�d�����y��|��3�{���(Ĭ��Z�{Jo�&�Wd�w�N�4�[G��5Lժ�>+Æ��`����+_#N��6��W��&�S��O��]��U����y���\v�E�C�tUHvb\��2V*��XmtU�Cm��Ӫνu���$������|x��_��6x����.��Ms&��M��Wtܗ�\�Ԉ��.9���Ɔ�)���8�����C�=�Z`.Z/iK���I3ٖ�׏���a�)nU�pn��랞��1�b��������S���*"W�._��dYOCe�T.EL�~��t���!���G��p����������yy�ref�	�D�/��0WqUrTVnjF�ֹ~-(i�s���l��!��j��mS-���c�ϻ��U3O�٣��ou4��.G�� =�M�^<��DW5���4�������u� -v�A�{��׸"=������z�k5�\���ފz�U}���];�j�-���A������.U����tp�3s���PL-��ԇ�����hB�}�'_0l�e���"Y;l]��Q[� ���(�Z�8�W��Q�v�Bn�u��P�X�I��4���g1�k�c)E���˼�rp��l1�-��4S�f�y����)C�p�ʹ!��r��R@���F�������5�k�*B�����uUY��Fmh���Tst���<�u����5�,LF�eZ�]����8*-��;2��@��V-Mt��yu��$;��R7�]��u�D�3r	�;@X�����ιZ3W5hXi�R�ҢW3���G��7���V�N�p�����[�t��S��T3������;@        6&{���*Iݔp�H�[0�pY��}��-�,ұtR!����b������V�j��qh���އ���t�%U���P1�����U���9�l�Wn�uv����4��_*�R��Y[vB�?���D(�֜f�_�s \S�s�Jx�L�_'0�bt���`�nC��xMʘv��}�59f�
\Ό/����wW�3�a��}ȼ��=�V��j$_Q�5*�r5���;�)�xf��1y��Lb�uXfw/j����P��**ᶤ�D��n`7���Vb_ȋ��S�w/�i	�Y���4�3�Q4gY��ek7+I2���wvgS�i��l��/��ՑΎ#�Q֔�m��MV��F	��l��*m=J�bqA0{��.� ��   8e��J�.8�"��qS	,H�AcY2��2�,DwE*�m%(�`�X,�+U
a-��)��Ȍ�S-4�%$�������)�PU��[%�Q��)�E"�e��e!�PX���,��YLF*�`Z�X
T�1K�2���T��$U��e��2e��`*�AVDLUH��1d)y��D`�� �(�X�X7RP�"�-�r�`Ud��}��Zə�{{� c�jZ��ā�hb9D2L�$.��'T��/L�\]?�=�����2	�õ�8(�����k��*��Z�\A�"�ܻ8'��ږ͵���A������
���P��&.���q�7l+:�g���	OcHS���<ק�>}�*%��(`�c�7��S�/�o_B��
��i��Q~�e��^��c=�R'�Wֱ�����sj<�5z{S�?:�:��ޮK3���ׅ� �.z�;+�f/x[0W�wN]�l�r�U�)5�NbG��^b�sږ��j���l�IW�oŕ�w+b���1m��̎b�	��**�]�w^�O�2FL�` ��;Бp��*ZQ̋68�c2M�h�d΂۽}�~�}:?Xo�׋�|����ʎS\�U]��Oٽ5����y�S��b����t��R���U~{��̞R7��߻£۵P���{�%�b#�dF;�����mvڤm�^�@�}C��lgy����^<,��ޱ�Қ�ýK�w�u��{3n�&��Ю��n�Kz�ɍ�%�0��2&�K�!�������Z�1�3y��~L���o~X=�8�Wc���j-xn%0��/�#�13����fx�1�wN�A~��z��z<cG3�R�F[�[y}����Y��nI÷[s�l�)j��󼝺e�grU�'�#�)z�9�#�qXW7D���=���^�ݟ�dM8<��~^�p��VՈ�q/�<uy�y7D�����9&@|�YV���fg��y������ƳR�4l(v�|Y~􆊯/X�Vy<�{�p�c��f;�K9m����jw̥P䧾������!P5���o��Bq���۹�3�k�J�/i~���9�]��� ���br����g2'z�M�P�ʖ^��z�����z|L/&J[Y&zQ�5;������������t��[�Gk�������\�4,F�¥doD޾�D�j�j�m���m��Z��b��_-=D�A�3W���9���Swt�lfK�@��B�u����%�s-ʗIu��͛R)�K3#[��ե��*��|)�4����疢4�ue���E<�r�Y�+��ty�o��nת�'�!��̚����U,S�նu���X�S����|�,��\�m�#'�m�W/I��b�Ԉ���u=ڍ���^�t�\�z*�ds5��K�amZP_{2�W4���u�?6��d
G�	l4,
l,[/���
�#�.����3m���W���
�G��v��*��Ee+��0���_�#�S�N4ۼ��'��y��r��	H$��?��K|�,�_,{�.D3�
٥m�����H��(u/E��J�I����1nw=^���}%Ý*�3�6���]���d����K4fj��=��Xm5Y�a2��P�s���jx��u��隖R���`��S��P��VjX���4
��Vʩ�+1�Xq�Z�et&���ͭϞ�J`�{棷յ�o���S��͆����F����7���"�ս�^k]_U�"l�	+G�|��9��ӡ3��z/:�Y�ٳ8KQ]��g�ߨ\��������a�1�%�N�D�J�~l3�`v��v))t�C)�]��-v�X�fAWŎr��E�Rq�oz��F4�햝�ҽSMG�Z8f%�q��N}��ȇS��4_\�}�9Y�г�ͳ�����Cŭ�ڏ.�C�`�V�������R����T���n[�q��JMƜveI�Q�7"�[�࿪��(}��>�n��R�,qPJ���Arx������ۿy�{nM�wٺ׫MG��n��D�)/���R�o<�ײǧV���C�S ~�=`�*����J���;5��3�T+��^Sl�6�q�f��7C�G�$9^,F,'e5��xK���o���4Xk���he'����5�Ϫ���t����CW�����s���s��k$c�W�4:���z|.G�]Ü�fH���4MWw�0��D���'q��[�B<u댴de9#�,����ڲ�kޅ��`�35*Z�Ҟ���o�6U�y��)��/�V�i��]�.�U��{�j	Q�'�wo_���]s2Ԯ�wB��`+�,�:�$�L���5à�6�)�/�����(ѽ�n�{���ݒ�-8Q��~�\���O�)�����p5{�@ƹÙ��tv�X�|=�=��*Ǹj����5[f����{ǆ�>�k��~�GZͭ=]0<r/A3=���>e�*�`�뷞Z�yq>��y{d����8�5ו��䕰���83�����t����P���\&t'�k+~K�H"��ꋶJuO4��V�䑟�s�ݽ��W=98�8.�7EnNM-e��5��%��bZwF�RX=
�c�9�0�/�f/g���o<ń��ͺ�$>r/L�r`��zZ1�^�Y�_���-y��{��-������~��}d �&z�ø�L^��>�t�ԋ�}��-v/gd8���)�����y�o�^�v5++|5��o�X����n�V)��M�b�����n�a�R{S��Nn�5���ڨ��{S�����F	��NoFF�#e���dw�T��Hʱ��~z��[�7oS��qKy�/�we��N]	(<�=��OC�kv�ʋ��]�F^t�{�T0�}j��zI�Z[�;fN�}�IpNz��%�O)z����{Q�e���X�Oӫ�H�]���!����a��M�J�術zy�[���/��ϕVE|�USR�^������ ��$9t]����ۥY�T��w���-9,�fw���'l}�V�������iy��b)��b�V���y��M��\�R��;���˱�	�B,�OJ���%p��cgg���^�G~�:��u��T�ƭ;J+ǌ8��O/��aQ�o����b/�<:��:f���V��-�a��!v�1SE���u��L����<��W����*���߷<�=n1Pf��e�M|�GovR� �o;%�1���/��й#i�I&�c������q������6'��H2�T��-mq�9�>��Z��_Kt%����\q���c72�m��P��y-�K#�G��a9���Gؤ��Z�G9�`��`WjYdN�^vӳ�O��|j۸����q���<�C�_�l��$�j�{�;6z�|��#��[g�P+c�HwMK|�V�+����k��é���am�uſ�k�)�u��SEÍ��xT��T
Rֱ�1�߇����8�*�T���V�3�ЇR��l���(��/�K��mV��]�oLUoأD*��Vjծ��S^ �b��'�ԁ�Rmh��/m魕��]1s�2ۼ����A������J{-s�2�B/�pޫ��RqDr�DzP�t:(�Pc�㓝1/e�h�����j}&�����F��;�ީg@ȥ]#,�e������i�r����yΰowX13B�	�&�=J�@�+�wok��ޠ�3`e�ǈ��w/J�����G��5��TDS�9�G,JN����4�������976��z�n��%���7\:�M��U˛�2�&\cբڝvh���Ɛ�Y�d���7>雎8�6�S�(������YW��7��P�P&�s��-�j�7r���.���7�%w���%j{T��6��� p       oUtGW1ZfU�w2Q���4WBB�Y�F�Ư�Vui��'���ٜN��Q����%���[��[[���ob�_mp�T�/���]�:9���:[���'~��}�a|�Vo�ei�� �bS�Y��!r�]��-i�D�6��H*���dC$����_Y����l�@��[�5}�.�'�a9��l�%nn�W�v4����!�b��$�D������FS{\a�E�T�e�U�(&L�f��=���ܒ�#6��-g9� ۂwXӎ[��-��uoc�Y�5�^�[}]nԏ,vh$|t*��^6���)����}�x��'��,������:�&cF�-������e�c���s$�Ptf��;��7�b�w��À.�@  y�����L�O�`i�RH�`���|`R�� ���L����Y�Il*�,��uB�aL�d�!L��RR
���*2�-�@-,�����J�dQ@
HZILa)!��aR,�%b�K`mdH�i��Td�`["�P"��,FA`���Ab�IUKB�"�E&j�@X��<������9\�z+���V�l�#�o8���.�7\�\�C�u�|�b����8
�u���@:�Ԁ�]&w�=lO���St!o>U� �NG�ۚ�\�2�Ԩ��b�vSYX�/nK���-��{�$�5���^Nj�;���F�2��.E�MJ�v����g[vD���#7���z��g\[�b[��,]�Z������}���y���xf�ϼ��y�$�#ܸ�W��$�}�eu�1�  ߛ���u�^�S|g)N3W���ʸ}��}�
2��DO{��x�!(b4�n�!��3n�{n��J���=��׾��y!��Q��Y��6�@|��+'5���sV�:���U�%va��AH3C��{�ژ��E��N"jr%I$�3k��	k�����-U�s�@�q~^��z�z
�^��D��v�]z�a֊����-I�v��w��[n���|=�aQo?1Eϯ��ȴނʥ]o�m?c���(��<�Њ�'	C�[

~+g��ivA������\�M���/t���1����? w/m��L�U�sF�w.���ryn����jm�&S�~9����&z*�B.��E�����:1���b�!����yٝ�Mڭ�&9�5�l&����87�9P�k���7yWS��k<��j�����T6�Sr�����/����y�>���)�4AGH�Y��K�vڗԌU�b73k�:<�G�+QLGWr�(��m����x�2̈���Q�t{�cL�U�7��J׫`2�����r�?�d��Չgj��u���� �	ë��%�6��Y�����ܥ1-���3 /ٴ
8( �],�=�=ڦ�����������j��<�t9���M]�~�rx[#����5���*��F��>��J_{Ԇ�'h_$eJ�3���ڐ;*ܘ2��ڵO��ߖ�J��cH:C��)'���{z��UmxepD\v$�4<�8�����x��W��JCfn'^-�r�s�9��v
��ꫯza�0���y�u�ђg򍅪�
�\k��b�et�9�L�"��}�����]j�4����Ay�r�>�����̈́����U`����La`$.�����/F��^�f��Z�{��b�}����(�kѮ�vpNm���\�ze����V�G+�םRn�X�/z;�a�S��k�ڕ�^�Kϊ�2u+�o:��Mk:���;a
���qهJ�fq�b��b���gB���a'�_Z����m��<���8q�ߺ�_dsFF��u�=#>�<{����P�/�s�*��ڧ�u�p�0�=��ZFv1�9���}}~0r��C����s�|E��Ә�q�6l�w�[pT̥����z�r���6�y��e�$y��5,)�S�:���Z�бt\|�x'V��Pw��O�k;�{�-���g�0����󱽵�=�CWj�E��d;��-9�*�n
���{��v�v[����Rb�wM�����v�S���$�/3�W������h+��9��6L��6���Nɫ&���M��_ɔ���F�3���'�ś[�=(��e�̏.(+1w��������S���+6��e9U��B���W4ٲ���>�Vz?_Wrʱ����Y���p9�0���
��no`g���C�dOx��S��P|�P%v��.�<�N\�#�W�]"�rH���&�ֈ�3Ul�m��<J�ֆ8�j�ѵ��%��ɋ�<���<lv�wQ����W�Y���N�Nv�oj��+�د�q_���K���Q�f{�)@|rM��r�E�E~@ا.v!�^�^��ABo�{¼����QX�^y=���A*��9c�u?dG�݄���5�۱���}Ie�>�>P(Q;u����o��_^c���WC��Ĺ�Fmj�G�'aQ�f�rnA���ٕ�̍�bW-��ѣe����lݘFDc�ط+X����(��T��!�yB��iP�ۑf+�p�M_	7�i���N�n����I��))\�d�"e��qI]���p�+s=3����w&/���,8gmez�^U6�T��Y���n�ЖdK���?���h���\訥Rƈ5�T�lՕy8�M
=F���G˫���s�?A4דֳ�E'r�)Z�G��	�����W��Qy�sEbͼ
��t3�rt�HԘ�����J��׫��W3��D3���}��.��oi)��BE�w:s���9ứ�~�,��f��5^f+����g���W̸Y��X�O)]{��Ѻ�#���k/0:R�Z��RU�"��՝ԍ�����Z*�13�ʘ�A�)��{�^^�p��RWj{D�f]if�/$�tg�i���5���_**���)x��?G[��8��J,��څW�����9�г�S9*��{�~�F%B�x����
��J=M�ܬՁX�,zL�u>���6��L(��f�[)}7�f�Zr������~��S�;Z�+0G��k~����^v�_��s�}%���³㵸���ͫ���w�^�k�vM�×{�*�N�����Ks3��{�꾉I���e2���ߪm=����e[գ�gV���d!�wy;Δ�*���9�iԥ�J��p���,�̚�ٙ����a�s�0d��\;V��^^�$m�4�{�3L��lғ}����a
���{�iC����[���95%��r5J�mA&��=y��?7��ڔ�N>-}�Ǜ��{͓��K��Y1�5��P����.p�Ԟ���Qo�E{���V��#��K�i]�\��{�z�VT�C�>���k�j˯4�����Y��n�_�O�Uڶ6�i5�8,_��I΋U �v���%�i�2�]��e�׹���b�T�SIG*��\z	�UL��B�_]����+>VE,���dn!��"o�݆Izxظ���_̝��];�6�卧k��gvS�áz=�A���LEZΝ��HHhǍΌ�J�<��zVǌ��-!n���{��ݗ���3�%����bQ|���BF��gOktr��j�r�Y��]��h��5+�|�~�[�A���lZn�׵�𩋞�y����������譧3H�yq>����%l���={��Cל�;@��֡��Օ�S,�ݮ7�F	��F
'���w�g?O6���6�-��/��I�^�	�^���_�.>�3��J�5�V��i�gG�m��9�"6EU0a��b�U���  @����@ ���Q8  =T?�`��~��aAvj��_ T0꿼>f�gS�Ġd$"B@�		 �$��a B��<^`��y�֢h�TPQ��B�(���3���!�f{P�	�!h  @�ċ�|Bq��Z������C�XXx��"\ԙ2f.}��0C��c~yE���aES��y'�HP��3��y�@  �C���~�t���$� }Ѐ @�0d� ?��$��0���\0`�O��7<�c�s�}�������}���4}��  6�'��a���" {�����C'�~����XJ5����2A��(�l���c��ԑ�_Y�!���<�����~�j]��?咀 l��ؓ<��)o�cB&  !��'݀��V@椩e���XXg�?��0C�j�����~�  @�I�M�%Y��`}g�>f>|��?�!�U���
�&C������&T� �A�5P5��Zn��|��2� ?�*Ft�X~�#G�C����lр����}(�v���ioD�쇱`LȐ�q��ب ��D�5���������~  ��2 �����" ���$ٰ�l,D� (���vB�UHc� 	a�  �!����p��	���>�����	7�l�($>F@?I+ ����X ��\�����6O�_! @�2d�2O d��}��2?N��5t�J��	�H\�Z�?t����'�g&������  @����?����C�   ���I��$���~`�$���>	�!�w�|�"t���̟B���O�G��ֈX��'��>��ɇ�������}�1�?�(   ~��L�G��H�
������Cph  @�?�C_�;��h��=���zO���Y�!���!�؇�.	�ߕ�XK~���������|!����tC�?���������C�g��>Z  ���d����}�d�}���b~����������L(C�ϷU���(?�3$?a�0�  ?��?@�� �??����O�?�}'?Y��!  �������H$�0�}�uI��c��M�|��p?m�MH|��a�	�EI������(��w$S�	��r�