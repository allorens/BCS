BZh91AY&SYT)���ߔpyc����߰����  a
>         @     � w}�    z            ��{�I%�U�+b�ǀ  |��@(BB�
�]��Gº�ݍۧ�G���j�3w��E���^�h�i"[d��cAѩ$:�l�ã����ݗ@ �R������ �, ����)
鄸B"H�DF�L�0r��
�q���4-�B����c��(���
8 q��a��fU+���cv�IU�=:vd]��R�;����Q��{�K֒���]�ǣ����G{�v{�8
W� =%gw(�/m.��e$R�4�$WY�z8�g�A0U ��IUF�q�^�h�m��u;��ފ�����H�A� x�cj ��ֻ�vݴ��+s���f�'��5.����e�]@M�c&����6�J*ֻa�G�����!>��       l�!J$�P� �ITE@@�P    �O��J��cD4b4 @ a�~JJ���LCA�#�db`�	�<�TDSF�@      I�H��h�����C �M*zz4�e4�6Ci�z�(
��LR�H0�!��h���h4h�ɦ����B�-d��KT��:N�$X�seEBa������A7����?(|�U��]AQG��U�����0�����9��!�@pAQ�X�p>Q*��$����(��r(�0� �I$�I$�
|"��!�C��^�����=��_I;��s	r�jQ�q2r��ԇD�a�0M�U4&����7sF�G7%�M�dk�l����:-ԡ&	��jڛ���# ��(�=�!�Ag�(�BhjABh�L8'M3G���Ǐd����aDzU'5ʕ� �Jq�J8'uel��D�8W�&&���6lM�Ғ�t7����F�J0㺕�U!�l���9�S����֦��D�g�N6��}Bs�bo���|�uQR|��ʖC�7��G0��WR�M�p蛸�]�_ȋepM�35'~N�62}�D��J���[0t"pÒ_Ɇ|�)0��_gj%�l�Ojt��I&��ns�$J��Q��}�'j}��j�䣜�Ђ-T�F�55R�	RG����D~���l��m��:jڛ�eN������wQ����Yӣr��jp���l�_$�!uuʩ�����5�'j&Έ�*"X�%8j��!�����TNt��ӢMtGvU����(�0i���f���(ܟ �G{���eN��w�N���N�0�(�}�ɳb7Һ"�,Ј50����QFUN6w����J�gG�0G��C�D�cS�6�J�NԱ83
K�RhLț5؈�
�67���TKY�BY,K&�hÅrpN��.��������7II����\(��G�,n%PtMH�Dı���+�0�m+Ie���M�K8S�~����'�'�#�Sbh��u(Fr���y��G���m)4pNRT�p�N�Yt�ѱ8'��Z�YץP�!2��l撑3�KƢ&=��\�[;�nDؔM5>~d:����nCf��pO�A���5(�5>��U>A�TDв�Ԝ�0J�S�J�S�dçG|��ۈ'V��6oq�q�N�\��'��pG;Q,���pGuQ,J0w ��S[�"9�D�j�p����ԉ�tw,�Ȗ:����M��2	c؈�d�s�PND�cS�D{ �u,Д4�N�&�%P�*"#��0��f��>N�T��H�&�h�[�!��""�:h�H#�*�,�N�+et؛�",�G�r�Bty$ؔA	#�H�?X�"<��5sb	����8"u�I�\�w$Μ֥|�d����тi�&ΜD��Lu*��JNW�+�MJM��rRo8TFI�6C_$���%%�8h�$D؍L:&���|��I��?"p�r��DÜer��P�KɶU�D�1�Iæ�D���WH;��c�]0ٮDI˔�l�E<+5�E&��e|��~�IL��uԤĈ�%t���I��TP��R�6'VU���tN�\��Ad:B���U�tD�J�6#�'M�T�O,����ʦ���M�H��L6�U)줡/'�u*�7ϢpN;��'���~�%��W��檟�ƹڧ{��:�����LuS��Զl��'J�Ã�;Q���T��,�{����J9!Q�A����U�(��e���ꪵ���0�I�TN�H�Ze���+UU��4��뒓��]�ãwT�I�~�����u_"�!��K;Fz�r����x'�}�S�Y��|��֥|�d���}���Љ�͚6&۪��kU��B��pK�jpN�N���&�XY�N�܇�)0���NvW����D���Cȉf5)!l�E?DM��&2N�Ȕ�Rk�r%~�A��O%"?"9�VA�DY҄ǲ�D�+����uܭ����2�蝓B&�ԑ6&�6��D�R��L��zNpԔt�Dӹ[6�R"9,M	����9���Wh~���4e�BΛ�*��R�Ա,y��тs�;ԭGq4��B&������e|�}��醹R���&�1�jNR���eD���U�͎B&X�v�I�:7�M��<��c�hj�|�	� ��$N��H��$F�4W�"Sr�6~��`�pJ8P��	_V�蔉l�IH�q�9EP�47��LN0ٷ�fΉ�Ie��gA��	mT�F�Ԉ��P�*p苕0�bd��58%���Z͝%��JN�Ī:q$��Q):ly ����[¸h�����g^�&�U5�] �ؘQ�C[(Ѧh���BSʮrcɡ(rhJj�ɢ�9PJ(y9��&۪Д�V��N��RWaD(u4&�5U�)j�h�������?6r��˪M�a�e�����f��,N�����'GL��+��4F@ϴA��;ȗ{�z�h��UYb�&QE��0Ll"!���DG&)"��z�P�u�X�r�>����b%,��(�r��Bd��5-줃�'j"<��Dӹ_?]J؎�'Y"%�bk�PDn"w]4c���t�t���/R���W�l~L6�Rt:ܤG>�!ڝ4�W�I�c�V%�䩙*����l���+��K#����l��6h��N���ѳY\b�0Kܮ	ӕ�{$�E}>�%A璜�,�f���B50M�bP��ڈ�"#�|�u�Ȉ�D���A47kU�u!����d���W�9w�-uĕ�69�R���r�b]���%�:�U�'��d�3��:��6��Ʉ艴NT$�&Y����:C,��6"Y�6l�.NQ���ba:l�_&Hh�� �e��>�4i4W��P�ԉ�NyP�8L�7�QZ"h�jh�5Bu��:r�r�ٲ�ԣ�'�Z^	ژ#ܩZ�ц���E�S��X�ɣB�3��Q*J�"�%��T�I&F嶅U!_ 렆�ft6{)�X��?��֙��U��H$\��V~�u�}�2_���o�>��~~���vl���6S��W��n�fO^���<����ن�t�~¿]���f�b06AǏ.^}�2��	�7�����QQ����C$��m�����x�9+��>]����%���=�B�47�B�N׍VV�(v�B�z�%9����{&���0�>t4����Up�����6t�VN�����e}ۼ۽f�gk��8��F��}�hjmm�ǳD�o6����{s�f����\���"�5��N=�r�ק&8sa���x�*�r�=i��T���b�����$h:����kz;�c����m�d�'8��W����l��>¹�)?����r�zִ,/u�N\oL�-��:����g_��ҝ|��|{��ܕ���Vp��cG��yq�=����5��H� z
�f��(�d��ә3x�p�JFȮV3��]�M�	�.*�:���&8~#7���GBy�ק�sӈ{Żr��J�dЂ2]��HH@���$a%����s���^^.��,�)���6w7
��D��:����o�Kb#p�χ����U��Ie}�(�������~���"�8�͕�4u7�o�L;��0�ێ�1�jި�߲�k��޸��>ŚM_%�}/<:af6����C�_I���%������H�!N�t��f���3��.��������RV"��G#c���f�;N\p��u�6p�F���?+Bx���9:����.*q���9�R�
´�)]� �L��d�� [�t�ٹ�l��3O���Jӻ�o�g� w�o1C=�`�"b���{*���xza��%���Nsxx��W��^�]�s�߭��4_f�<|g�d̿�Nj&���D,ř�Js�Q�������`�=��@�H�iT��6��� �V��(�ٯ�/�Q�^?�Xf���i1wV��{{^.kg�۴�I�_��	?���Ğ�Y����q�x��ݥ�@^O}�fV�-�2��ƍ]pd$��z���� qM��/N�Ǵ�h���8z���:�~駽��T�s���S��Y��+7˞C�hg!ar�V�طZ�$f]V�o�(�}9t�bx�y��ɯ��x�����gڽ;�aS��}��"6F���Fզ�K�<�ɲ:~�O��8_=<~�m�␖�4"C�e�������]�K㮙β'��|�%(owz�ڍ|��DG7-��ٯ�$	""��i�!W^rú��>l��V=M�G� U;����W�4��*���)M�`Z��c��V_���%��)�Of�8���$�ˉ7��� -J|S4�=��&��O�d�>�i#ɛ
�"̯��,��&����~l�������ϝ+����?/�?�_q������s��N���L�#G�
y����I>�\�Ӫ�,�!��]Y��/��R��"���we�r�/r��f�:�.H�7��Y�!��>��6n?@�^D�=cǪ�3�Ӳe��"��i���=�)�6���&�7�ִ6�����י>6�Ov70o�Ӈ��֚a���ǎ-?������/]4�$��6�{1�'3.�˘)g�[oN���}�H���L�W�@�-�ݰ���d��1�"j_�fz�Ll�����o=7��M=u�v�*�BOA��h���D��ـ�A]�;6��pd�iw[m���*��gw~?��߽�_�iG���W��b�������̧���\�ς>#��V����'音J�k.C��4:BP4}̩���?����3�M���u*l��N�x�W;���fm�<ҭ,�Bg������4_o��b��;������E��Q&���H��N}=v�"��x���:#��s կa��Uu�G���Ǧ�;<�Ͳ;4�&cE�׽�/<�Nj7}3���6qZ�>9}��VQ��O���a�'$��k�,r��E_���B����cMz`�٧浓�]�3��=�_XyC���m�y��j.�/�D!+��3o�{q���l���6#�]��{���8���/,l�h�Wp�̘fvi߈(��7�_�>GK�c���Mj w8�^+܏K5���L�su�?I���&���bVO�p���c��-{�raӸ��t�$+��_�<oͷ�?My��҉ҡX�?��{�Cע>D��<��FI+�ٮ�~x�hp��;	�%��禔}����<})�7�m&��E""�ތ��Ná���vYk+\wq5�W�K�D�^H`�V�F����z�r�OXZQ���?=�ܠEL�0*�=�N�wt)� ڔg��K��M�x��	d7Ap�r�d�Z�M�		�#E��K��0���M�/�32��^�wQ�93�=?$����al�wL�����I0�?��\z.���Xw)w���%��K%,�8��c����ek�����{���B�g��m]�'[m�,�v`�äϙ��6��w�����P���y��E*8�rf_�U���l;0�+o��7p����=��Μ?���t�q��?i&{���d��<��%���'�in�<���5�qۧr{*?
���6�}2َme�]wT��/��wa"E��]�3�>��y?8J�����؝w&k����N\1�pv0�S}���9�g���������A�LZM�n��²��L~׊i�Ť気	Ӈ�JxV�a����.vBv"�bn�m�~<W����3P��㤼��×^���bf�p�,G��J.�K/x�^�<rs������s�2��V9"N��|�8y�3M;$��F{76�N�m���O>t��魘f�G<��A�S�����sZm~0�<��
�t1p@��>(�����c(�8yM4���ii�/>�ʏ��D�ܟ��^�<@����F��ސ2+�S�4�4���s��:d<X��8O8��$�9釸-���ms\~,�����:�c��&_8t��4��G
�u����2���kֶ�I��������>H|�!^��s�M�:&BG��@�:���m˓�o	�b���б�M�\�Q�������Kej�aQ�m��ѕ����#u�4K�.u��RT���Z���)Y�"�]���$�Q�#	s�;L]������Y�����V�1u�p��_�4�n�ƒ��.Ѳoa�����ͯįi��m�v5�d�:fbT1�%\��1S.Zd�2$	�cB�_�2Đ�_�P���"	�����$�%&�+��hDd٘-ۙ�5p�ç��'�Rg
�t�5⨆f��T��6sܝ��R?vѻD� ��^�+Lie4�P��>u�����7�s���
���<{XN�_����#>m��I�]�5]j��Է:���L$;]�jg�Zv��Xb������\DT�1Vh+��huQ�9�E�]A-EP2!4I�D<�6llw:�f2��c�U��:�D�_�}�G�3�{:�5dslc�7�vL��<��|&�4�D�I�IWR���d�$I�"�@�,���h����cu��»uq���ң�����QW-*ݹ��Jm`mY���0IM�2"��s�8�y��[9ex�}�3]�5�w�_C����t�XMi�sd2aR�^SG�KgELL�}/O@��K�RV%.禼�t]�M~�<��b0�L��cn::�n��#l�>tq�z+�#�z9ηD�b=[�#6�!�)�&Ϥd��@2d�����p�	����l��#b�zcA�Y��bCY637g����d녘���u�AA?4O)߁�Ѷ=m��LOyc��=���eF�Sa��p�}e��e�W,�q�%�p\w��S]L4���p����x��a�b��kхP�)E���Y��2s�Y�x뺡�5�J�|�"b �H��lZ��?4F�Me	It���Ś:�3Hǣe�����%יCcR�M�V=���g�X'���\���	���7?&��1O��7�;̈́��d9�a�n�a;�6i2�x�P����`7p��;�!n��s�êٝ\f��Y�\N��x��ݳ�Qd;gv���N���U=H�b"��ʨMO-8���&��󲭙�c��'֩�u[9Г�j�@6��Аݿ5���ȅF�x+P�������x�;U
����H�;�k��W�~��~���hҪ�WJ��^*�Uz�*�kUqZUn�w�ꪣ�W��UU��U��t��V�U�iU[V�U�y��p>��������+m�UU�UUq�����W\Uګ�W��U^��V���U^�UU�UUTUX���/v��Uڪ�Wj��^.����@>��@�$���	$�[[ͪ�Uz�UWUUQUV֕U�U�UU����x��Wj�t��X�����kJ�����V֕U�]}�j|}'�'�'��'��k����g�Ux��Wj��Umb��"���UUq���ۗwv��*��t��Uڮ�W�UqUUUUU\a��B@X��d!E �(DY2"���94E�$d$��ᇻ����5 ���Cy�t�%Γ3����P�&	�&tC�pM�hNt��BQ�E��(К,��	ba�`�0M�,L�ı,K�8lMDM	�X�P� �$�lD��	�%���(J �	��l�lAK �A�DDLI�QD��؛�N�D����a�BX�&%�f�
,NtN�(D�"lK�YÂ&tC�����[6�ӧ]an�UXJs�o/�v�����~�vn�sl@�MrT�a+�145�-�JVn]��4cq�$���%`�$rߑZ�*X����Y�.����ńĂ��5D�.��$�����.�nf�Z]��9�@���V:Ғ�I�P��*�y��c���im-L��`�s]�k.6����ږe�2��M2����Ez��D~R(�d���j;Y��튭ҷni�n�^�{%������]j��0��e��]v�bV@���DՄ��-�[�4�)�n�XG�\�.���8t��b�{h�Xؙ،�e��+�t�� ��ōuK>v�):�x��ͩB�:��m�	����bБ���&K@��;l���o5�F��:�D�;f�[pJJ�n}��e�Z��c�x� �k��L6���A��6���3K�i4��θ���X��V�BlkVW>��6-��UL�X׍��bi�8�P�!�KAU6cq@�`���TiQ��l-2�����L���K(�IU�($�A* R,����J5�g�[�65ţ&*6i��R�rHZ�$�i=���6��CγX��U,�2�֤���V�k�ٲ&��4��,�� �`���e6B#�	D�(��)U�G���Pe&�?R�7���e+�MkYG�sw�+1��\I���R��)j�1�9���l�7U�ZĿ3��'i�A�"NB� �1�$@��e���h �e�f�-�0s\�sp���Z�g���S�6Im�m�k#�lh���qv5��\�M&Է��%L�U����4��W	���j(6VW�.)G[L�颎��64(�� �%�XM���q�52�(J� �\Q�٘#."��s�5�����:�F����K�5����4	f3��m�M$�p�D(���$�a`䤆  �tD�(�
�é5$����ַ����PCVWmZjٶ#�5=i�6��Nd��b�vfڃŚ��R[��G�S�W|`��h4�I6��-�ax��n~�}���kv��Ժ[W٘�'a�b[����\#r�X[��y��{��Mp3�6mt�uns`�D�1��X�e��CZWY��F�)L�1j�ۚY�4��-TT�DEH�CKw�Y�ݏ5j���cX`��d�'��[��������>�=�{�������O}���}�{���wwwv�{���{����������UU,-��|�<㮺��؉�4a��o_��v�Y�k�wB�S-�6"d�QJ �n�
�2�ۂ��hئv����\v��<�_f���(�9҃6ʺ��.-6���-#1c�� ��B��Ԇ�k�v�S&0;A��:S�p�C;��#���ڃ��PA� %��L��ZVQ����y���q	Wk��fۆ��bksWh��fa�m"���:�&BY��$�ص�.&�Mi�iv�q_F�� � �fvyi����G�Q!����7H��g]���-���k��uE7t^�C��w�P����ӜѱV����)����y���ó�u��C���.�������80�
RtS�	�˝�CM=N�{'F�ag�gY�u�m\�x����<0PJM�!�R@��G|�6ř83�C�
[����?vS�ã��	��L,��4&�0�tM�;�
�*��!���Q��i�Tk:ۇ��'T=�}(��~���jS���&�� �z��n�Mb�|,�C���i�I�K�4��(w�^٢a]���SY��)��PO!d4��'=����{]�8���SL+��Wu��V�Chu�[0�`��Y�6"hMa��߰�mCd��a��s"�U2h��0�Z]t��N��k:�S����C "F���(�������=�6OqC��0�Z�vta�ù�s��hXB(�����3�Y���	����#M>왥e>ah�l+k|˯�0�0��lDК0Æ	Ӝ����=�ᝌɁ0�i�#�}��(�e�n�
�ېڙ������U�GGa���2�ŶR����|J�)R�xk�J9�\�WWU�PÈ��r�O�)�-m�?6ҥ9���l���F0�-SL���%{ˣ�Xmǜu�ĳbhDК0Æ	��wMyBDPТl�م+-�S[1�)!�]��RN�21ԗ��H,�]jPS[n�[�K�k&�1�G����zͱb�
i�L�������{C-Bf�z�o��Y��l���c�J;k�=͹~y�S�N��NN����4(�0f{W�'�)a�E=�t��3g�,8`���e_�`���Ɉ�M,(u�>杝ã�p;���><;0�<0�}��A�N����=�Z��)�BB�U��(ӧcv�7sr�:�L=,=��s��L0�ĳbhDК0Æ��-�M֣����*km�(J��$�óa��Ox�"�����Fv;T��ЇgPO'x�T��9��i:�zI��d�c��(�?{ J(߼��a�%��sK3sNk��L�n�<<����僝K#���SZ��S��d��w"�bKEU����>u�|K4&�M	�8`�:^L�U�����L@��@�g'<Wv�c��w80L)����'$:`'i	���lOx�O{�8�������h{ߝ�����q�-2����r����Ñ��C���o�M�v�
�Y��]�>q�`�t��7�ps��K^��rS�Ȓu/F�)��T|��[[N��	�X�hM�Fp�::�;��j!���h�Hz��ޡ�襦A4�J���M2M��%ǎc�T̶��8%����w),��z[�a<,�b�g��d"�)R��Q�d0ҩ8h��0r�]U��"�mʶ)�C���V>�1U�|�I�05Vô��l<�l0K�	�Bh�'~��b$��e0�!��ˈ(C�&�JH�W���m���hYm�AΚ�����T��ae&t�5�@��5m�C������m�Cx�f�0fa�"q?A������tI��Hɉ�h��\��|�P^��{Og����6s�[�"xw�A}S5��Fi��%C�;ߜV��I9���ZdE};
rX}֘�'pO�s��I�è0�0zQ���J��]�jV�o�L��6��R$-گrL�ϫa�^q�]`�%�B&�ц0N��
#f����7'x�P��|F�v�J�?z6Ծ��}ٽ.R�a�͆��t��!�(l��Hy
y�^�,��
A>	�ֽ^���n��P:�&���m��	���l�2���^s.a�)6S��7Ü�퇲��M�Ħ�����$���3���o\Km:���|���c�?1�^c��|���ˍ��ܞj�<���a����Zx�=s�1��̱����������8�uuח��uż���������q~N<�<�&�_]������e�O/ͼǓ�:�m<�a~e.x�#�y�2�<�y�{��1������O4�[���g�~tM4t�����R�aK�����m��a��/��'�����-?�?'����?#O/o>o3˷�q�'�_^_�_����y�mo1��u<�qo'�///�U�/ͯ��w'�]�������x�Rx�M���0�'�$�d��\�O-m&�-f�a���A�~������=�م\5�T���֗��<�M��o<�-y�v��]�O�G`�8<sr��fS�s>�N�H�a	
a���1��7r�C���}�X���c�]�z;.��5]��ݻ��e������!��u}��ד0�A��=�\Lu�m5��^�9�E�9_;��Z����w�����3�{���뻻����|{����]���g�k�����z�������4x��<xN�<YBhD���N��ڞF��U����}-nZf�806$���B�D&�����aC$���!�M��:aЉ�A��Ķ�E���'l��8!�=�74�#Q�`��00I؈�`��N�I�M?~�W��B�b��D��T`?F���ļ�-5��h��q�(��_RI�`���j������%W�L�Ja(��Y�"�UW�۶2��ҍ�%P�Q�Va'ݦ�ѶQ�@2C)@Q�"2���?�UT���3{l�QhG��b���Ue�y$Z�Ct�~]+�����q��_<���y�]u�m�$��*{�ʫD'����?V ����d;�[
ly�H�J6�����Z����[��~!��,�@�.0��T�O� �)���I�!DD�d
�UcIUY��:��3R�" ?!t�Z��T��z6�DDQ�?	a>�-i�A����I�E1(;j�8M(��D��,�\�K��i~�V_�Xx?��'Qt&��pDL��t$'i�g�2OD>z������Dj�V�uD�wU�>i���:����<�<��ˮ��ͭ���f=l�ev�rV�@�؅"���$¡��O�$c��&��s�R��\��>ұ~Í}!�� E(���!3'Ɇ�Cc�����$��D��N��-|�I?A2�"O�Y&�#Ə���v��O���y��,v�/Da�Ӛ�9�7�g��gp��L�μ��ׇ�ji�d�0�#!(�?$;(����2����{�L�h���dd�B��`�"5B+��r�KW����������'BjL�;�" "�C�E��)�xY�P���}j)�3�'Bd�%d����/V[�c	����%�C,�B#%�d�Lq�.EŃ��ň�E��)�"a�$?P'�$�I�(�I;m�<τy��n����˘mݥ�3]|Dq3*��z$�)QQ�)]@�2�:�U����ݒ�T�K=#e���d��r�S����;q��|���<�<��u��y��Z�)��S1QDD�,�p�H��|2h���d��N�,D�~�2rQ�+��G�V��qO�b�Wī��]}-gWYEm���'�����ȦFNɄ�Xh�E)�N�Ibt�DE%�B�w�n�rJ�J��,��DD'�&�|'���Ns��o�">@�{�|�D!~�i5��\ۍΉ���ɳȇ����x2X��Uv��agR��N#h�CH�S�d4в>�!�"~&�<Hv0ċ$�K'СX~�DD��Us��1x��4�R���"�:���מ~q��x����6�/�
���B���dH$ҏ����ϸ�����2~�("C�>�y����tQ��,O"s~W$�;�V|�C {F	;O�L:��^I0��&�0O���,�<0D��4hp;�C!=MHv0���~2&�����<KJ�\����4�!�£�tU����d@�()����JI*h��0�'b�D@D�)C��$�JO���8~F�q����"0�2'c'���,O9���!����7w3nf
!�t��K	S�S�6	:�t4��N��8d; 'D�2�[%�qp�2�N+~G`p���"	*�S�O2}Mv�>J1��������${�1.n525����t�����2�.�ۯ6�z�ZȰ[�$/V2�ͳ�}�����DD���%N�_�������=I�&@Pdcɲ� !���pDO4���%aH!J:>��E�Z[^i;d�d�d�l
�?� �K �j=�Y X���s#&�P�;�lĤ�S/�.�W)�.��K#��"lm�%*#�n���s�]���5F[�ȱK��n���JG(�7IUZrD����3CuT�w���~�s��Y=�!1%	���C؅�%��#��ѓİI<�{S�C�w"!��`��:Zc"	Y��U4~m֟??<��m:u���2�.�ۯ6��3+��+F3�_�<��)����MJEJ,LNj@�1������hɰ�K�E�g��*A�G�m�mȏ��AW66�����;i�}|�'���*��������W���o���{s�'�e�Q��=��.eT�PBn+�=�^�p��e�w��>PS&�����,���,>���.��G�G�VP�%��~J������� `lOa�Hm'-#�����I,��A�@�C�E8��D����������*S���0��é�(�v$7�[K��������K��;����I~������ )FHT8lUl&0;(�"'��I��������O�nHl@�`@��pC"ȅC�F�H�C �y�OǓ"`pB�s��.[��?w��!�Z���D;#&�؁�P`,��	���1 b~�|��J�"�P�i�������iӯ<��a��u��y�'C���'�}UU�2�<M���)@�2`0�a>#���+������R-g�+㊍8��aG�����X'Ǧt::�7｜ɉlL����"㨽���'�g��,�C�
$<;)�O�pN�n��e:��'T`'��n��S���}F"��f�ڜ���W[�d���7v[���T��mT�h�cGe�oM4n��?6����]T-�Im��7+�h�F��gj6��*w84De&C
z!���as2�>E�j��¼ێ>u�����t��-�e�]u�^m�bU�V��$��T1=9��*�!�I�<)�M<E:�U}�*-ϭ��/*)�Զ�D���/_I�O�[�0a�qm�#�NJu���˘�É�%��D��LȖ��I���t�t¡�G�Y:(w�u~�6�&m.�a�0���'R����P�짓
CH ҟ�Cbp����U��1'��:��Vj2E��5v�R��$7�L�-�G�
x�-S��Θ�1��Zk�϶��g��`����[�i��>�`%�J}�����~~~u��:���y��i�������l2Ւ�[�>�Ub)<�Ԟ~�Z�}.B�pJl�%ؓ'���0���D(�OK���<8x���O�]��f9��M.ls)�x%;)и�J��(�G[t���+��Gꔸ�"�]0�"��j�D"7�ikC����G���G�2���bݬ+(��F�y�ڈ����By-��BO��|��-%��p�e�6Ǫ~������;���9g6�T��c�]4�;��~`e�r��/���~_?1Ǘ�[m�:�y~O���y6��6�L��u�<�Z^�_�]������c̰ǑǛc̯o/����:�����uż����t�8�8�N'�_ɤ���x���yzy~O'�y�8�4�Z��̢�O=r�c̯��b�_��<Ǔ�\�~<�-~ap�Q>���覔U�GO��W�������k����y~e~]�=���<��8ǘZߗ����?/��_����?6�d��y��y������:��Ou-ď>c����9sk���$~u�N�1�����̯Oˉ�y�y�&�_�/�8���\��N�s�a���8�<�yyKO0���F��Z�4�r���<��s���Ҙ��9Fk)86	@6"�>Y�\�u����a,�D!5�٫%˭d'a�IcFbp�	����U��h���������T��c!2�k� �/�i�Ex�*/�y�
.�n��n"�.w��Ŷz"G�:|��B�J�!�Q�A�M��i�"�Uӹ5�'s�!C�[���fb��j.���E��]�w�X��X��u{L0��vo���*�O�=�L���!�����(�l�ϵ)�d��ZB?b�)�[��Ӵ�ko��)1!�o]?aJ6��N�����7Xg
�毚Ma���}X�q�r�������%>�>����%�Ph��\��-c_�$��� B�0J�5jKY1Z���W�.�S��ژ�V�L�P�E3,#�K�Kc&��[lһm�����@ʩ"'��4�
���P��@�.G&�;dn���BZI�GEhL~6" ,��i	E��5�$T�����b�&��m���x�榵[5���'��/�|�]�����*����3.���U_{333/�U}�����}���DN�O(��G�ӣ���~��g{�l���;f\�]��5��e��׈ڄ9f�J�ި�̤5Wm�֎��G�p�K���f���S���Lfjrc$��p��l�Eym�:U�B'c
�1���d�R�+l���u1#Z�Ax���8�.�G��v,������Sk[v��qf�1�{Z���������>m��-�L2Q�$�A���h��∅�x��I`�E�r��X�.z����닶^6gv��}������F=�\$~�		W��O�C����v��Cɧ�)������ɪ�t��=H��cT�0[�߫i�c�\���~>3!�r�������ͯ�Y�1�;r^�F���:�d�r�'�i8u~x�ݺ��~|q0�f��q�i�i��uP��+����ք#n&�BO�lg�|�X-��0��ey4��Ĺ�#Xei����y��t���y�i�]mן5!!�9I��$�D?%.��2��~����p�+��[n��j�9OݓmS��R���~���^0����ޓ��JEFϩ���j��~[�eW���S)�n�n��U?h{�Ni����}T���m��W3u��;wL���zu��6vr�5YGH�*�I+�_�b�U���K�v'a�O;��|2n�N:�����*R�$�]�n�K3_�;FXE�����m:u���4ˮ���v'OXX/�ř[=UT8׽r��s��s3�L8�?1�[a_����e�[�LV�ϩ�kLU��y[���}��Jzi:=��J�_������B�gh����;km=|�������c\^��>=>�+W�$d���k��u���o�w�[���*�WOC�,N�)�'9�p�0�|�*�U�]r�Gs�Z˹>2Ӕ����n��g��VI�mN�N.��|�:�5�~Z��:ۮ���ζӧ_�[�0�L��n����Uu*���0�>⪢O�S�P���i��>%n����Jf�bHI]n�q�0{����}��*�5e�������|�i_����5KC81O�[��M��n���0�ٶDL0���#��VG���=����!�3?v���i��N����8���6(��0�l18^I��;b(��k�ez�Q�[n!�����dC�J#�Lְ���[iq�ǟ�~u��:��y�i�]mן����r�>F5��C�2�=��q��Y�d�P^e����16ȁC·P���~�쁟�	��$����Jl��#��?ŐHt:&R�װI$������j��N����7J!�'F�dk}1F�[��g?S%�3�^�\w.5,ЃKl}���sx`�z9�<[�}η����΍��_!�h=��e��0�+橇�ߩ��6��k`�L+4�/շ����,�ܒ����Kb��'�ق�2rrr,�6O%dV��\���,,d�)���a`�!]�۞O��N�2l���|a�=)����O�������YK�;.5�!��LS�q��Gu�ú�/~�!�)4�8�8���?:�N�y��4ˮ���W�3s�L]�WYi�UTC��.g�NCa٤���̷������r�f��=I6~|u$�a�����8a�M��Oߓ,VS7����4��~���V�F�}U��u��4��-P�~����K\�7xݜ���ي�t}>�a�><�rJuЧ���l<9&���ĵm6���9q^��bw�m��}Jɭ�I&��F[v�e�<�<���~u��:���y��i�[u�ó�-�g.���t���F�B�$���N'3���.���x�3�~�l�dy�_h���+�m��&̲Xj�c�;=:0�?wޞ\���!�_U���r�Bo���c%�|�����P���$�;,S�z�8c�7S�߿Z��{>2��~��p�>�=	���!�����h���׸RRɆ�HynS>�S,�$�d���U�r����8'ϚG8���ζӧ^yo<��4뭺���L[2�*�	�_l�@���AT�Y+ s޳�n*��ra=����fM4�L���0���*x���AP?Qs'�_�#v��A{�8a��:4���SN��tl0(eZ0��sZy��Z�WϪ���X���$���e�d���%����6�1OD��2J[h�F��l¦�k<SMN~W�_�N��M�|���j3g��Ӎ�����kn&�4��<���מ[�0�:�n��/�cD�XX�q�H�Z�R�IiP���tc��SnF�Gmq���D�l�;:�җ�94��&\�Z�.�`%�����o�$�
i�Hn��"q�T��Pk�T_�k%�"+o��UC[�gJ��!s�5�ք�g�/����WżQc�wٕi{��>Ψ�Sh�Ð?��ꕖ_��u�O�L���6���_��_��3Q�5�-�����1[v�i�+��L����9Yw{L+	_����W�|�[gK��ꛒ*�-�m�t�Xi�J����fT��O�Çs8&�x��=��m�6r�qs�"�O��<4��Ӆ���Z�~��+�a�u��\~u��:��y�^a�]mל��K����p��I$C��]�u�unѿ_��r�6۔�KC��cas+e8d�ٽ?;i���d�Һy�����ݷ�p6��?|*�w�&\���N�<vp��������.E�Y��}��.�;d��i�!�roi��q���.D|�m�G�a�zM����S���S��a���Ggq��6�2��������6��~q��__�y���<�&�_��m-��'��<����e�镭����Ǘ寯VdǓ�<Ǐ��y�ǖ�����I�$3���)<B��|�<�y#I���^_������y��O8�̗��b����s��/9�<�Չ��<�y~N0�%O_��Kyq�ؕ�&�2�L�����k��q.��L/�/��y��-�<�y~O>_�]����?/�~L'�n~y�����1��<�:���K=���a0�F(�
�<k$����<�����^_\�ی�m��O��?/���?/���>y���/��u�b]�kZx�yo-xL%��<���˷��[)�}�[߭��?k�M��8m]�@�/�-��;��h�$�(�R���͆\���qC1���-4�M�|�� K��Z�~^a�^����I�.���4�c��LP��Q�G���|sk�?qz{�=�1�s������GcG�w��7�	�Wft�F;��7[�������3333�ފ��333��UW=�����誮{9�s��y���:�<�Nu��/0�ζ��zI$����q*JwV��e�����~�����ZFx�:I���"*V�Ù��Y�o��
A�	j!E�O��:��nng�S����O'����ґ�{�n8�/���6P��Qo�+t�I �Hi�i��|Ur�.ϡ���J�U��sN����b�[[F�=�b��Rc�8��yן�q���:��y�^a��mם�5��H��H�EEEJ�>UU�<)���ݹ����hj6 ���G!��/"ZA����HHTG���b�|�o?T�l⟝m�%}�2���r�o�b��L7Y�,���-�Ed������֫�:��+�H�!�?Ca��<6o��Vxt���V�4��M���(�é�	����y˪}$����[����ʹ��^[�2�<�n����z�1�֤�Ѽ���Ҥg�5s/���"D�?,����R�����T�[F�^&�	yjnRkX)�m�t������P�Ard�~T�O��CS�a��B��$�H /迮~�#��A=80 f�^�������a�/���
���2�%�E��>��a�B���`'����0�Y߱�ݦ�m��I5[��ڧi�������@Q�p\f�=$`�K��r��'k����4�ߒ�Å06�9��|�=Z�B�C�҈x���a�({�-tm�e�q��+_�=�ݴs������g��hb1M��9.�l�X�#��Ӵ�҇�����q���:��y�^a��mןe|��I"Uu�����o��Ι�э~��h�ܟ�l�i�b�3a������S hti�c0U��`�1N5���#mU�i�SY\;<9�;9��;9���co�Z��#����A�"���:��3��i<�3]��m�N6�ŪJ��֩M6��-��~u��iî���e�>=:=>�LO�'�13�UD7�,�F�O��y�?}ܳ<�TY���������2��߷˾V�����W^Z�0o�-�a�.a�\�����D�(ϡiK[�l��w��>�������p�6�%ӂ�W}8{3�.s�,N�p�!��Bps"a����D��P��z�OgGgG�n�/Պ����j��G��Km��8��m8u�~y�^a�mןl�U,�����Z�b5��*x����'�0ᓵggʜ���P���'�]8l����_³؈l?����2��kn?�[q�S�"iyn�m�m��%�h��[8?�u-Y�eV�!�a@�,� ó{[N���Mo�|S��c�p�x�q>K���4���?}�..�j��2�2��˪�Y��F�[N���ߞuלq��p���2�(����+�ā#�(�q&�-��/}�+���ј��F���>�g7oY�jP�զ3)��M�\�nL���շv��*�!�_b�`��-Y�Pg�N�H�0��;I=�AK@�_{E���[�EH�[���($q>���p���`�C��v�4����[C�x�~��d�i���������߮_�~}Q)���ά�w|��cb��>��][�}���0�q�|��?[5^�:��#r��4�Y~����>��D?v����؇;�`#�i*]G�a�a��B���[p�ʻ�������-��G��DI�����5M2�+m��qǛiî��<�̼ӭ��c�]cU>�����#S�UM�p�t~��0�ݬ+M�0ѭ3X��)��v��/nKW4��[?y�պ,�a���w5#�6�il�����2�s�u�.f3��ƙz?�a�z'$���5_�'�W7�%J�u��M>7�5ؓMS�>����}M#-��u��iî���2�/4�n��*��^�H���F��Z�>|sP���"�C���0;�óJ̧"lA�||Q�qJ"���ͯ�����nf`���<2<<��`�qn�ɷI5�>Z"��m�5]ql*0��d���ynI,1}NS�߆�؞��� 'c&)n5��1LS��X��ލ��u��.�Ֆ�4���|��Ky�u�q�m�����2�/:�n��ڻ��Lb����w�}⪢d0�a�ΡN	�����mKkR�S�rW)�s��m��*�`���{�a�֘6�d��3��K�{�\K|aF{��	�;4��'�e<;�.tN�8�-�>��|Z%�~}��&1�Dh�>������i�-������6��ߗ�;g�q<�������<�e�>O'��.mo0��^]y�4�Kyq<O$y~[�y�_�����k��c�����'W�y:���Oa��W����Ex���)<&��L�G�_�_��>c�/���y����������痗�֞b<�<�<�'$��G�_�y�%�����0�ԕ4��-i�<�張����q'�^X_�_��\��%y~O<�=s��ˏ\�?1o���ɏ�w�?4����/�q~i�:��痷���&+$�XO�0��Pʓ�VI�.y�O:ē���&�Ǯy~O2�&�{�̺�������6����q��O'Q���[�G�io\�q�Ct������ˮ��,�R�5x��Y����= w\e�"Eyz���gIǝޡ�!��(��1t����qiޒ��㓳��m�����{��K+���R��{# ��$�H_��%/͛��۹g��p���]���:�RYl&�e" qG��f�_.V�ʄ�����U���X�}bU@�ꊖe�P1!�	������K
��\�G�,�����+`�P�:���m���H!o��S�y_K�L�aې�^�AAP����y?�H0�q㘁4n;��Ls}�����ۋ��U���[$Ai��W� +X_�L���W���I����!'
��_�Y���C��� b:�n&��w�<�im�[h?M�E�ƣaQ���;-��9/%ٗoT�΋0�}3.�����sklw���}�5�а��L�u�?m����]�/��B��T؊6gT��@�`����f��X�V�GQ��C*~�̼���333?Oz*������{ޥU��ffg��R��{333�<p�G����	���<'N�����(�֥`p�ucD�^�f�f�n�ٚm-1,.���Ե,��E�t���!�-5����T�R:�(��)er���4�QbA�^H�74��D�]c�� ��٭N��R̆�,����\�u%�l�D�h�4��>g��|?~8���WGĎ�$Xګ�+4�s),���i���()���ज़`�Ar��E�v��^b�R��k�������U����%��hЅ�#.4�_��I ���Z�O�z�=��20���XZp�]�G3:��c!�?q�եTQ�F�A��Z��Sƾ��/|�1�'�>j�C������yM0�u�5�?[�-r�C��J�Zv{Á��	C�^�dӲ��#�:Ӏs'��yj\�A4�ȷ��MV\�X1hE[��=���0�K6P���{��r��-Ɏp�[f��wf+�əl���~��	씸%��`vv���f^�=�)�_:��|���?6Ӈ]G_�~~0x~��/���c	$\9������'�t�4#���0���������A�y�j㙙i�pD<8t��DAC��a���}0��4�Z��=�q��kh�=Y6�2��2�?��B�(��)�LS�A-�q�>�ϒ���x�RN�ٺ�kZq�����������za��p2�ם��ba��Ɋ|�q����0ݲ�̭��O`�8`"A<x��g���9{���N��E$��_K!�k53<;UTC��iv|���S$B�&WKe�χ�DCm4aH]+��f�N�M2qV�DC�LW�0V�࢚S�����'8_����ؙ[f|������h��Gwxc���-�v�^��,A4�8}cR�_ǩ����u�I�y�en:�8㭴��Qמe�_��>�*�!���/r�m>��`�����Ij�	|D�D�`BdE$��8`߈�����HZ���գϯZ�фj���~['h�8�3HK#�]~yD����eWN�g��uv����-�ٿ3����_6��ĵ���NUF��1U�JKM�ղ2�n6Ï���q��|u�uיy��i��G�H&x�4S�m�9�Dkl�I���AO�Cm�(��O��%q(���X��IJ��!���A@��8�18�ZI�?�6k"�Pn�>�CF��f6!I$�����
v�I8)C�A�����50`Hs z�Q7�)4!�	�{��N0\fH"K���p�C_C�l�&�� �,�i�����!�>���{�V�x	�JKsӘ��8O����!,�nfe���,���}�Ȭ7H�E��W�'6a��a����d��m>����i�Ç`���M9�&�a·��?;s����WM��7.�`�g�gp�򽟘�w��AVv�jآE[�"B&��+��]4�L:�����a�t�`�O<l�:'�S�#p����%�'E�qQ)���"u6�X�Xu��,��I���8S����wN�L�ɌF1)�[0��l�/�� �Ab��!e��Kp4cm	_����.f;8ye�a�ٺ{�տ�����=���q����ʹJ��H��u��ͣ̶ï:�:�O�����/2�����J�bD�F.%y�{UTC'f�aA�����g`��9Ԥ���2��;�Ä���É0?yݫ��e���s5�3yL]��d��a�'7�[Y�<�=�W���]5X�0pʖ�y���v��鶚r�3{)��vn�[T�0����X~A���(��S�"�?q�~q�_���q��|u�u��O�>=:=;3��K�L��s-�������6-�"�o&j�8Շ�\h��ͻ��r�0�/pό<>�t�Z̼�)�&������~�r���6�d/MV�'>��w5~����5�iݬ�FXy�nMU�i�Yd�m����S�..�H�k�n}��]ʗ1�W~u����µ���:��Ɍ�5�����~y�m��]B'��6xN�g�Z�I[�
�oTc]a�����y���8;lS�@jI~Xkˌ�%d�H`P�`�-�(���$����A�� ��v���am�Pk�Y��-$�H :Y�v!�N��B��5Ts	�{F��] �	?ab:�H*��D܆�։R�I9f(6
�����Q��� �E0�T�4��j��2���~e���eS8~䚦+�~�ԯS�2���(y�p��(�a�Q'�2?W�2�.]�C��,W�k�G�}MR�V�柩t�V�R9_�0B�������5�5�v�#1��a��9�Nb��7�zy����i��2N͆t��U�������I3Ʈ$�h�+u��q��q��|u�u��e�[u��n�(��r;�Q'Ŕ�J"�����
4PfJ+|�S�b�ْ�S��[��U���84O�2L�Ml%u�l�z��s�:�\w4�j� @����_��&�(�@��K`d>���Z�J�Jי;=��b(Ku�5��2z�ܓl���4�e��^�o�3L2�4�l���N�x��,D�0L0D�͝�tАM�,І� ���4Ab'K����0,Lı:l��&lѰK�DM���4PP� �$4%� ���P�$� �l�a�d!�A	BQ�h���6�u�XGN�<��-�e�:x���N�tDؘ%�%�bh��0L0�0L,��d��4�S����պ���x��<�EC����'��F��֫���7���O�j���H����y�
��U�ϲc(O�\�O
�����!P�w��!�f�t b�R��S�!���h��w��o1�z0�+�	"Vt�*&*�	f��j��~����U��U��2W��v&�N�R=d*����L�֦!^��L����j4ߵ��B����\,cD����`7*��"��������-�`c
H�����g�33=�z�W2�������*��������iU��ffg��㇏,�a�t�`�M<l����'�5$�"������ӽZ{:)�DMAh����D������e�Uk�I���oF|i�����,���}޿�a�g�h0�Q��.8]v�J��Z&�ӑ1XB���M��/��p�<y+�LW��aQ�Z�i�Ob�Xa��)�aC��ҥjy��E;����ޖ��`�C�?L<Y����`�p�D�&�6xF�&x�~`���#�L�^�I$I� ���k�U��Ŵ�b�A�bX"�=���?7suҎ�n�ѳ�O�sl�q�`0b���e�0��h�)�q�k-??0���?x�+G��k_�^��S��(��Ű��������+��._��F5Z�:0�2d��Q�J�����em�ج��׺�|�>y��m�̈�0�,�`�M<l���=���K�8���h��"�Q#2(C*�Y�6г�\���A���`*�]H�u�g0�eH"�,���I���~���zLv�f��ô8T'#��(?#�Q8���f���={w�C�Mub�2x<楚�Y�2�R��m=�t`u>��R��<����[���>vI��R0�����^�~4� ��Lj[p���yã��f��ҝI$��V�}]2���K��9L�5U\n��l�+Cu�D��ɦ��8�d�BS��m=��t���s��ѹ��p�۹r빬��\_r{=?A֯�uQ�g޴��G���H�|����ǌ0K8X�M	�g��u�TA�VĒI�_SO7OneVms
�Mni�<:�Ʉ���\���ժ�q�5�b�N�����~G�D%<�l��[�~-��Z�w�e��}5����O����=�߻�O.�h�L��~>�F�r#��ˬ�����o�~��r��`��i�k�H��NH����?���혚�t���H��[������8K8["ABx��:'Z�UEQ+.g�@�qUQQta@�������l��o��?��4��߸`���n-����I0�=H�����2�E�"_"�$"	-��-n�0��yN˸k��w�R%H����O!bx'|i&�jXa���=K��ƫ�2Ga�sL0������j����c��6��3��Bp���<&�<&%�,D�&y��u�LһrI$C�uL�X�Xwrֳ#�PC���M2�YΆ�_!��}��s6�\�6�r������øi�N@���s��8���Z���Io�[a�<�:��7M<��|D9�䑕V�����kL:�s����#�8R�?�m�*�~2	�����tt`̰�^i��~e�q�_4뎭�Lx~~��]��q��b!81�m2%?���&N�0��J�Gagv�Te���A�	�
��f��]��<�����Pdh���I �7�IqIs>�64���,�G��{g�l���2��G���]�7�W��<H�wޘp����o8<�����{����P{,�
!�Sɰɑ�M����١�FN�����lQ<2��P�*V�co�9�R���,6��?S�z�|����p���r'�JwI�d�CF�dC>?[v�קw7L��LUEG�}-Ç���=أٳ(ٺ�]�������M��[`���0���	�P��<l𞝖n�hSњ�j�J��lL���;:)����P�g^6�:>��3=��L��4�����e1��2F[�6�.���S�z�2q�1e��Nd�8�4�Y��R�_G�3��5Qط�O�zk�l��cW��M�7N��ꏚ��&��e?Q��h�m8��$*K�I=O�n��v��}�n5Oe��Ym��u��6~��,��%����2����N��(�v�ĒI��GpC�l��>Z[8i�l�2S�2�|���I�+dC��'sM����CӅ&���\�ˉv�bҦ���Â���O��@M�a�M�u��[?C��є0=u��w2n��J��[�1�b������i�KN��D�A�O>��{մ:w	P�����>y�e�qǟ4�P��<l��f:&��z�7_W�UE�0�:z�[ꪢ{���Krzv"?#�h����ϖ�����b��G����;�V%mH�o9Kq�m�h���~Ėu�^��.g"pe3M��DQ�PA=�~c�Zw�>�Mߝ�K�j�_�����ɝo���8r�[�b����VS��MW4���$�g�>Cf�|��im��%S/��ߙy�����M���\t�0DHYÂtN�	�GMQ��ABP�6"X�tИhDN���,N�I�D�Κ8$8"'DЈ��4h�(�� ��:a�6&	dC�A(�&϶6B �A0J(�(DDN�����ӧ^y�a�^y��y�κ�gM	�YbX�%��å��agNN숉�bpN�.:��iӪ��<���<zI�Kɑ�/���h�¬7�ުNi\����RM�O�XBьFӷ�����ff��=�z���}��k���^���*<��n`��ˤZ,^!�Աy͌{Hy��W��̵�.Cq2�%�D��R��3����<�C]7����c���^M�36ʨOV3���D�I�V[��)�϶�6��� ��Nm#m���!آ�%b�V�7Fq-�	%$�Ϟ$��c(�Ӭ������k���:��u��n�)�=R�s����ѻ5Sq�c;e�Ik]���������3^���ѐ��S�G�|PٮX�_�U#�Ӳ;콹Ǌ�������ډ���5�"[��-"�Z�?G	g�qmۜL=T� �'%mz�
�csÍ(A@�tD�J�(�4ZD�8���bR�ziu���:ŷ|{By޻��5U\���!�L�u�)�F,8L
8~I��I��噀�T�gmn��m���zc�Zܕ\��og5���J��b�fg�33����W3=������*��~�����{j����9�i[ͼ��θ��qռ<�� �<<4{�R(����L�2B�ٵX�\u�R�i�X��JarPs�&ɲ���DZd.6
P��H2Le2YEILQ�����sLZ�^Q-��*,%k1S1lCfg/i��[�R��c��MJ��m6�̬�VZVh��m�-�4)Ek�@��h�:i@�f��3����i��]��!T��������XQ	s�8���S���,�M��k��Au0몄�������((�R�.A����I �������P�mP��zZL�x<�n�I���(|��۩q��b�h�c7��B�t�k��w�D<Q��]������k�Ø�N���?a�
~;6�4����S�|#h�7��n�ҵ�?]b�E����8�j�r��8�IP�m)-��D��9��;[��n��ݫaa�|z�<|� �6~:=>��n������������3������-��u�ٕy:���V�-�����'��1��Z�6%����<&,L��F6&�����>����]9ꪢKQ=Kb�䕊[��2C���_�V�/��/�|�ʽl}�ob���[ד���)�<����PC����S�i5M#��j��S9�,��r(B�$�P�E�W� a��w�A�@�07���鐥�X��ifLźr�����5c&+2��ϭ�1��u-�W�p�A
t^�h�����Ǆ�ŉ�P�h�G�q��Ļn��$��hoRb��!n�>9�2�:l��]E�_�~���SE�{�׵�W�N>F���Lq�a���j��l�-Je2èw4L0�2xӱ)=���֞O~IǺ�-Ut��|¸�-��D��]��l6p?D�>>~��a���1���S���|�3
d��-e;�D�O��O3�h��y��y�~y��|뎺Ì8�θ�獼k�����Z����<?y<U:{(������D��?}]-���F��n��O;�쥁�؎�zLt=���GX~�]J�ɺa��R��lR>�����_�3q�p���\�ܰ��ܚ'S�Ѣ&����������M����ic�����ԯ7v�u�pϿW쇰��bi��?U�����]�.��q�\m�y�q�θ�8Ì��>g�|�x��������D�%	�%BJ���u �p��cāe��,�hn8 �$�l���76����b�y���U��u۱b~DX�C����"i�<���t��eS+��T�b�D�oh�W���g=p{�л0�0�	�e�nv�������Oe8y���Y0�;$���Ji����i�HLC�瘥F��H����񧜇� ��*Q;�S��3Ͼ��S�aD觟�p�'|�������Ɨw&7�>/��,<����3�������ea�+�2�/�%3NV�a���~i�כ~y�|��]a�eǜy�1rYB$%$A}�Ub'Pڿ�����D�0øvS�:��nz��5�ۘ����k�>�H�Iyb�H�0�ۣ�}NO{{��p�WC?��m9�^l ON�"&��̟���3�/���֪ܹr������+�����OM��FG
&��3���V�W�]#�h�v�W����Qh�W5*t�r?BzԄ5�\L`��?O�!�Ş0�D�x�,Dц�4�����{N�������M3�VTGͰ�.*-��<�7��;O4�9_���)�~�)��K��"5�L�{�\s.ގ~����`�	Jp�9�Lܿ?��ڹKM����̈������u�6"^�a�<����#�Â&HR���})�g���w��ն�1|��Nȉ�(>��C!�����q�Ќ<��Deo>[o4��~y�|��]aᇆ������I�j����1���z�~��aІ���riN����?�iD�m^�Rط(QNN��@��I �~�j@*E�
��>�m�N�	�WzZlH��`�u���;O�DGޮy*�ީ[y�����w;R7O"9t��5�����6��r[.>�b�|�0]r��6e�0�8�V+��˭8��o�:�ϝ|���p������
��X��1�P�X$��w#g�0�8K��n��0*,m8�e�>���ȵ�Z[�F� ��`�
	��I'�?~�E�ih����.l����~��W�rC��%=#|_Q�?;�a�� ���ۄ�J"S��td�Qϧ��MJ}=�)r�6��������\==�Wsp�C��Y�֛DjS���)�)��~��dq�{c����ᦉ��r��4O��h�����?�+P<�R"�	�����V�X�Is�G�~��;M��̲�-m}Q����r鈆�m�ͺ����<&,K4a��x�ś䒜m��(6(YҪ�A8a������a�T�5N7'��>��X�N�L�;!�/>v�uF����r��n��vz%�)FpNU����Q=����D����^]�Lr�۷r�3�~��@�O{�v��NA��3��J�Ç��2KDik|�<�ҟ7Uh����?<������ї�4������0K��D� �4pД@NA	GЉ�b&�K�y'ȉ�ą��X�'D���lHP����Dw"h�B	���H"i%�pDD��Ӧ�GV��:ʲe�FB�J �%P�"""X��Y#�N����/2��<�o<�N��&	�,�,K�N�P�&,K,K:p���6X��BtN�&�l� �%%�(� �4x��T[�_(�e׳\��Z�M^�'����Y�'���nLDˠ֡x��L.T$�I�s��/~?�z�w�e�6v�(V7���F@�\�I�G�w1�&H��<������4�OĢ?6~����n���)�I���u�)�_�z	�f#�����h���õ�O�sux��f�Y��:�$@}�{Tћ� q#�$�HÆ���W��w����̶����;�K�l��{�������{j��������{j��������{j�������<t���:'��ŉn�Ì8ˏ8��L�$��7w�&2�C�{�������<�}4â�D���4�4v�;L6�ͼ��2A���S�E9��tM�ܮn[��E;,>�ON��4�S������q�w��}�������>��?G�bX'e���p��������3�L���pi��ҟ�7O���DZ+���u��i�y���q�ξu�a�\yǟW'�*ΔC\���U��:��!�S7U��Z8��e�yu�m#<�ߊ{w�x�/0Ez-xv}��g�Z-j[����<��D{0���/=D�=�xtr1��x'�u��U�u�_�<�H��	~O����-��8��i�ٶR���H�b��7L6���ʶ��^<�Z~u���O�0�bX��l��,Ϭy���h"Y=�ȋA��4c0������i��9#)z6NS&����EIFH(BЁ������,�ہRR�
���$��b��ЍT �d��H��MeƦ�ْ9���B�R��H��B��W�3�AƧჅ�a��z'S<���̻Y:;��?6؜8"v.���p����;�Q.�Ji�a��b`�>购_���ϖ�����|�Zeh�E�]i�<n�����o��=|ҹ��V�"����l�us��Ge���O�����Ѷ��o8�ݮ���F��~Î�酝:p�,N�?�ŉb&�4a�Ϗ���1
ª�����Ab��{Ҫ�C�gߡ�9>���i���|����6��b��G~>����20�O���N~�Zz��w�7)�=2f�Z[h��Q\�f$ULa��~���m�p�#��-�ĉ
�E']��v��8K��ø���;�uK3��O��5U�oq�M>���Or�~�(r��)�v�aj�Ͳ���m��\y�u�q�<���vx��y�bՠ������<r��.�t�-��Hg��nc+f�)/�$G*Rӂ'����v�D�a�a���$�Z�m�>:��J�L�L�D$D"	��n��O'gǳ�I؟D:b�4Dg�ܦ�v�r�U�DFݷ���e�3��ߚij��g�*G�u��ؼ�?>��3Z���m�\mםa�ıBh�fx�g���p�$U��D��Qg���Q<'��x��4��cBFcl6�II������/�4O��s�.���)�ݤGU\����c~�E�G*�#�x��c��g8vp��4�/�Ҙv%���zj�v��h�_p�	���������j�G~��4�	ߞm��?0���'��M	��Y�Ő��bn �l@�,Ί����d'�e*ч	�~���@�5�W��%�79+�vj��X�1,'��O��=#����PH@��\�Ƀ�/ACd����:zs>e
$�"���0YNC�3w
��mwכ��j�R}ߵ�V�U����3M�Z3O�un�R���3�n�*��Z4��6O�������~<�pM��&�����z�Oo���g瞬/�!o�0�l���m���1�L��0�?q-�d�3K2��Կ���[8��.X[{������9>��z&�+!��'̢���,y�<�O�'O<X�"hMl��,C���$��玺��y����ci=\�_�����0��t��7Ze�?7R�z�:��_a��>�/�Xz}�	�a�'����p8$�λZ�����BS̤�J0�~q�����z�==��3���~�<�w&��QJ^0�_Nɼ"?o�IY���0�?8���8��o<�>y��2��|��mf�bU��w"�D�_՞øt�5nM<�}�l��JCĢ0"��y��_���=<�d�'�'��(a�_@`�K_�?��RM�90��Ju0qx+�D��L�vx��Jx��VXC�ʬ�5��������/n�n��">�զa�=��D|�îv�K5U���i�a��0���D�g�4&�6ag����H�T�U���P��j��C<!������Y0O�۱�PPA��Jk� �τ~$X���O�/�s�[�B2v~����ه铨�ɦ�$�]4��#O�Y��q���nKz(�I;����p���w�8i�a�g:�^N�C@�5�]=)�R���2�J�4�����e0��i���??<�μ�:��M:ӯ�e�u�aգ��D�Q�4"<��A��Ie�bh�,K�	�	�E����$0D�� �	�(D�8tН���!è��ӧY2FYDd��Q	��B""&	�h� ���g��7�x��ǋ�0Lı,D�+$�0�bt�,��B$8'�Yb&8'������(�%	Bf��d���Q7L}����/5�D!�䂨��L-[���T��4�lr7N��sy)-5�sy�	�i���IKi?vqP��qӒ�3����8Pb9z�u��V!�����+��P�"�J?v�~8��<��3R�M�KkHM�a=��P���#n���,�TcԲ3�fv�����!��u�)Mw�x�X�]��$D+ŸlnT�������s�nF{�2U�Ʋ�(�a'daf`s��ıta��U����N�<%5�zi	?p�*v&0�N�Y&]a2R��%��B�|����&:�\������_V��7�XԽ(���Dn�v�{d�3h����b������.���5.2���[_Q��l/�	�b�3�q[r�6RI;���2-T�P"�i+��w`l%-5Ѯ 7�d�p�#M�a҄�! )=:��(����ы�6Qd�G�¹�h��*m��&tu_����8�e޻�h��o_���^y���˿���{�����v�����-��������{�ww~����㇋<a㧏�,�b&�ц�,��h�Ӟ���e&���a�l��
��m��/����5�F�N8dd��E�blQ�X��0')�[YQ�E��B���X������#X� L7Y���Z	)��eM�3:�`˵���L��]��Z��B�\%�2��:ֱ���ih8v����ZXj��A��E6�Wf��E1tb�Y	�lX2U�3�t�����)������)XGf8��I)L�H�D(���$�� ����I���o��;��U���3��v��u�z�ִeT��Yl3R��u����`_O�;���y���F�?��Dtgm���K;)D��a�xzHJ��RFxhv'�9��EW����-jB9M[4��֎��~����"�g)M'����O�(#��D�ԙ��[)����G�µ�,�w�a؂tS�m*W�tڣ���	�Έ��'�<X��Xq�<��>.UD�؃n�X����NCN��Љ�;����O���Ð�L��`��)Ѵ��ɰ�?}��\-[���t�O���7N��ժ|�3�I'ȫ�1"!��e4[U��dA��p�}��a���_�/)K''�Qs	z��/<a�i2���i��y��xD�g���F0�ǋ5�8Q!R��t������4�4��;�e�k�W�|�]#Ֆ^wU%y��P�����m6���Kzږ�V�ܭ��:��n�i���t�2�-.��5�}�Ix���즩ǝmǖ�=R�!�_*�Xi�Ug$�4�5N6�W][��jN��<&�K<"x��DM	��v||vu�m'l7ޕV"~�7Qt�����R�r�i�7X0���}��aG.q�Yt�
/����ِ�������4Z6��Z]~I8�".���8����m��˓,8�髹�	>&�9�#~l�	D�^�/�4����Ͳ��5�6ˏϟ?8K?Ox��4&�0�g�jr�kEV6�Li���%l�R�ˆ5&e0F�xjCK��VJ¿�K{�
7�m&�Kjr�Wv����@�q2��I$�A����R'�H�K	��a��1�]԰2z���6n)&F�j!1��1��9��j�3)?1>���	�c<:=��u��Za���R�z��~��f��:j~j�~:;��C���*��j��������ӌ��b�2��M�����w����""~�\���Ƃ��lF�1�[g�`��dŉ��66 �~�6�ܛ&�h�0p_e���Z>k�&�It�ut�l8돞q��κ��y�a�|�Ϩ�D�֩�\=�Ub&��YN��&]}U�k��w�~��[|��O'����)ߑgz��L��0�DDd�|�>{��ˎ��ߩm��z'^,�����"9��m󎙣s.9������᳇����:(�C�� �_=���`�6����.��n�MR-�[�`��8�,�Z�5|��]�9i�z�c4�:��n8��Ox��4&�0�g�g�I���Uu�WZ�:UX�L�a��81�4�n��j�y��W�"ҟV�W������o!��>�؝����L��?|`��9��6%h)c�"Xc���k�u�i�e�t��ޓ��F��.��W�i�TLSy��L?l0IؔN�����هpӿr�0D�W�S��ێ���ξ~uן<�ΰza��ó����Y��30��U���a�ѽ�)/�>	&w::��|r(��^�6R�M�\�p~F_fvK����S��}O0�7]?i<4��m���M)�^B�ׅ����l8w�J"'ޢu����`��oy:��ӣ4�6v9`�拴8^�Q2Ca�����Lۦu9��߇��֫�Ϛa�o>q��:��<��4&�0�g�l�%R�{M�W*��H�m�Feq��)Z(I$��6U,�$caʉq,"OG%�m�5�s�p ��pP��!}���_�$�~ ��=ڮ5Y�瘩���<�G�X�5��ͺ=��1s+(d����K�{��|O{m����m��Ӑ���~�����0�0��M4D�g�>9�JѺ�C��tI��b��;ÉȉN��ҶQ�D��xa��'��U���K����h�a�2��,�-.:��5J� G�6�wͫ���oBWꖜ[��e��u���0���hMa���g�u$V"0����	�2xv���,bᄫ�m�i�N7NS/nN0����$�r�4D}Yu�w$irtx!D�.̝�O)DM������(���Z�3'����q;�5���<����y���=d��>����OS��+?2cSr���I����sr��e�n�4�/�~y��2����0L�x:x��f<��e�����n����Xt�p��D�0D�;R"h�,M%�bYĜ0��4P�P����aB%&� ��:hDND�Ή�!� �Aa��͐��~d�	D(DDD�0MA�D���,�㧏	���A!ba�,L�K�&X�,l�8P�D���	gDL,��!��$!�6B� �P�&���o\��k�e}���'��^3b�y�b4�
k6?"<�t�9�/_d�0���� AE����L0ꇍIjJ�>�� � �7���嫣�OK��{�3�	|���-sD�t�+r=	N�CR$Amn
\�j��Әg�"��[�xVu�wW���G���]�����ϟ\M�d��?!�2��V��0#׾����߯����{�n���~���{��www����{��[���������<a��xD��y�a�qן>n���I*!qUW�xs�^�N�C�/E��m3�����Io>�X>F�z�Ԟg�'����QIȣL� D�vtta���Bώ���{9��?�WM��ԝ��{bp�0������4Ӝ\�)��	Ԗ��m�Ӭ4��~L-��uǞq�_<믞y��a�q�y�i���kjI$�O��2Y�|m���A�|C�w0�u�m�[*(�Qӱ:>�m��q���a	ϐa�StI�2s��R��
'�~x��~�:0N]y���v�e���wyf���F	��d�`ø}ϫz;�?p�0��G!�����1�:Ԣ�o�4�#V���;O4�N��<��8xM	�8`�/�Q&sz�i�`R+��Ä���O�Y2���R66c��B��F�_з�D�8�DZ��v�hPI�)��I'�+����~z��o��H5�cd��x����"�Rf*�L'������^�$�w"C�gґ��1�l���S�in#V|��L���&1���Fi�_��8�̣��ӗr�^r}���;W��=��[m��[�e�z���'9eğU��0�g䬪�d�DJm���b�U����(��⤐� F��@�A!N��]�/���M�_�:̶���?2��<�κ��e�u�i������+bZV�Ƃ���U�=R�1KDe�kIm��".��$
�E�ؠ+�X�����R8�=�1w���ݦ�֌a�9��w/��8�0�ilV�{�-�7x���c����v8w��7�P��LbT.�n��/�Zz�S�?�j�;����o?#G�u��_2���?8ۮ����y�a�q��mW+�U�UV"s�
-0�JQ9�\��(㒫5���T���(���c�Uv���vp���>��t�t���i��1�<� I*�Brۆ]�pG�g�fNA</���ż��S��a)[ﾗu���b{��l6r���۳�z�	�s�Q�v4Yg�<"xDK<x��u�i�[y�$�z�w	Sj�n��D�ν1v�ǆ�WA���x��������<���������Ȏa�\b¼���NO�hù�>��n|vv"�=�?bp�&���]��T6�ڑ��~ܑ��5���α]~*��;�����\�+���z����wi2�+���:���0O�Y���4&�0�t��ۭ>NJ�Qu�ĕ�R6��2Z��MM�ڂߡ�S��aE�!�F��8�(j�QD�EA�"!�
�9S��]6��if�֨3qD�$�~ ��E�7�Ԑ�bm���������D	_�0f)-�4�	-b�d��D��noٔ��w���be��3�r��|v}K>y�}V�ͥ�\�T8�>礏;^q�Coo�w��X�ާ�}�*sg!�k{=�����oA�'���E�/��������S���'A�����3r�`��b�ȗm�;��~�td�-S�e�������/6�μ���y�a�q��s���is<���Ij�C��\����㖜�Ua��p���'�f���꒤�\ޯm5g���籺���?c�>5UV�/$ӵ�κ�ޖݕ���ǡ���=�X��A�N���H7�(Q%��F�!	�7�����B��~N��6��hʮ���IQv���c
�c��Zq�/8���:돞y��a�q�m�wAd5��v�U�̉�kK\:���{�`B�؟����?��:s����&h�b;S����)is-q�S-�ǣ�?�C�l?}~NO��C��}S_���m�b����>����%W����~Oϕ�i��#��|�:�<��^u�<�/<��8�N:��Y!R	 
A�!U���q�n�{ZS����Æ��iه�s��[��\(��f�y����%��p����;���p�T��,���?qS��]���?8�u�Y0�̛��L�cU��'�~ԗ�IOU��r�z��7Y&�)16��ȁcT����N��F��
��				J~ok�=�}I��~�XG�m�ňhQFT��%�(Hĸ����`�a9ё�@�X,j�A	HB�	P�����%T!	D!	D9j�U@H�`�DH� ��%T!
��T!��T%��EBQ
��EBRP��!*�EB�����!�T%B�$B2 �"	dA � �"�  �"�����JB���B�JB!)BR��!�P�"��JA�UBR	U��!	U
�B���BR		HT!)�!*���B!Q	HB��!�!�BR��* �ADD���0FDD`���	�$F���� �FD`#����dD�#" �����%��0F2"Ȉ"	"2"Ȉ#H#A �#A"# ���2$#@F��2"DA Ȉ� ��F���� ȉ��#"$D�FA`�#D`#"A� �"2"D`�dDH ���"� ��A"2"Ȉ��D�
$���0DF"�DF	F�1 �"	DA�#D`��FD������ �0b
""0H"0FD`�� ��`���1FD��D`�A �DdH"D`��#D�##""2"ȉ�%�F""DH��D�A`�#DB"#"""A�F�0A��0DF"0D`�"A �Ȉ#F"0D�A�DF�Ȉ��D�#""2"#A"#"A�F��F"	�"0DFDA"DD`$FDDdD��H�D��
�n@��� �D��H�b �� �#A"ĂD`��0D�" �D�AF �D���$��#`�#"2"$��#@FDA#" �`�#a�F�"DdH$F$FDH�"DdH$FDdD�ȉ�H2"�D�Ȉ#" #bIH���"2#�DH$#" #"2�"A�FDA"�D�#H���#��F�Ȉ�H"A� #@FDH��2"DdH$�#� �#"2��#""2$�$�"Ȍ	� ��FD`"ȉ�%�F2"0AFE#
	�$D`���H�XZ��@X@J %)Q)��B�T"!U)
�����!U)!_�J ����H�������xQ���D�D%!��)��*T	Hi�)	P�0@b���� �2!�2 1�HQD#���Z��D%�J�B��,`����D!!)%.)t�BRBUB�Bd���� �A������%B��%!R�!1f �	HE@ȂD`�"�!d�!(�!)BUB�B�]!B�JB��BUB�]!�P�J�!*�J�B�T"�D ���
��D%T"��JB�P�D%T!	P�%!J�TB�P�"��"���D%!�BQH�"! �1�0A �A��h�� �J�A	UBR�T*�����!	HD% �!�D �1A��1�0A" ��J�A)
�J!�B ��C륑
�J�A(�A*R��J�D%T!	HEB�	D"�(�!(�!*���!R�E@�dAAD`�U	HB���T%!��"R�P�P�D%!JB�P��A	HD"���"�T�EBT!A�`�2!� � ��2 �DUB!��T%!JB!R��*	D"�J@����BR	H���"����)!JB*�B�"��!��B��j�f��JB�J�!)�*	H$"	HR���%!J�B�"�)BUB���HD%T% ��BT!UB!*��JB�P���%B������P��!�"	P�J��BR��%!�UBQ���T!	D%T!)����J!J�B�BB����ID �0AȂ �!	P�J�B��HD �BUB!*���B�T"��%T!	HD%TȂ Ȃ1DDD#" �`�DB��!R��%T"�dA��D"2 �$A��2 �"!
�!(���!*��"�IHEBUB��RH�dA`�0A�		HD"�P�T!	P��0A`�DdA��BT"�Q	HJB!)��"��T�	HB��JB�P�B �A�DA�dA#"�D �A#6� �1D 12$BUB��!)�J�D �D �B!R��JB!*��EBR�JB ���D"�D*T"��JA�B!*JB ���"P�T�D���BT!	HTBT"��%B!)�EB!*��%!*PJB�	HB��%B��BT*�A�BR	HB��	����iR��&̛�l%�ZF�Š4�� u0AUA"EPT�@(�%G뢷����ٞ?<����t' �"\O�3 ������9����LB�&�A���`B�7��,��=�)��yG�F�0�=���ۂ������QC�����~_���LCzP�������QG�ӱ^�}Y�A?k��z�D����b���*	Dc@��܏P��X#�NG`��d�H�)K�~`���s4<�{�1����C�D��QF4cƏ�<�B�@,�%l>{Љ�/yB�#�2�"Y�ؙ���q))=ɑ�0�4u�Fhbe�O�����0��Z�	�'�bm�R`�Pq�@ ��k��$���2���TV�AF���-��4����V�Y��R�]`���<.`�v�~��op�5� v�
�D*��B��
*@� Q�+ (+P!RX�{� �W@0us}�;��| G��#�v�vw��4�E�����B>?Ӹ����HEQ����W������E����(��w`��30k��� �#��nb`t���i�}�b=�E���o@?@s
�s����#�t�QG��R4_�j���6+Ǩ�� Ր�$���TF�܂(��H��"�!<1=��(���e��jzF��ங���b����wЂ�7n�r H��MFĒ����u���J�9�nۈ�q��J��)
�1Q�CA.�X�� �b6��`}�H�,A3a%�f'�sUQ�AӢI	�;�P	�Ю=("�<�ޒ��$�ޜ� ��P�@~������u�� bH%�MC��s0��c�N���=!ۨ�� �$��,��P�π����S QE� o?�� ����+�AQ���5��C��P�`�Àq8�7
n7¼J3�@��E#C����p G0���o3`��@�z$���^��R�C xiq,w�;	�ظ8N�� �(�����Eߋ�RJ��q8�ܡ���8Xy`�s�ni�9�i:�HQ�& 툥��P����Bh��� ��?�1Oϔ�L����ݐ�Cq���<C�����<�[.'f8̊����\��Sڒ0�% � 0Sp�_�����H�

�2�