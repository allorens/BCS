BZh91AY&SY�����_�`p���"� ����bF^�    � P     ( �  �      ��@      �@PP    (  ��}��P�R��]j�*V��l4H�JT�a��U+fUUi�4JUJEE[2�B(4d�*T6���D%
٨�ϳ�"
D��@$��TTU(�X��"�m�QQR� ��UUU@�U*�+l	P���U�P�TE*����H�p   n/�Vڱ'�����h8�d-�Hꛥ�fFn�R�
��uCjj�GEi���ڊ�mt4��\��V���r��T���!$%�ԪO   �̕JR�-��^{٭0*��,��5MJY׵g^iV٭��ޔ�wt�Sq�{L�iM1ޫ��hZ���V:�!mmǟ|�UJ�U�6�j�KM���v+U���IPI(�/�  �>U}Uj�u���
W�ٷz��ûv�e�<{�/Y^��V�x_w��m[kjZ|���_m�4ն{��l�[YK{�ޯMkb���{>��)��i���<w^Z�
Y�ީEU"UD��%	R�W�  ����LKm>�;��b�j�}���}�����Q���%�s�cl����ﶶĦ��>･��������ڦ�Z�ϫ�*&ڶ˽+��j^�������j�,�Y���1
H� IRE�&�   65����ͭ�6�����L�Z�����y}�Q�)�m��ԛ)Q%��>��鍖���}�}�+f��_+��OR�Ye�z<��m������V��m��{��{T4��]�}�NcR�$H�%A$"�  ����c*�y<�U��m2�+�u{B�em�7�I�筬�����m]�\u孚ҵ�{�G�qum1{�{��֥4ӂ:�VF���n���U�ծ��DH�%��U@�2��  �W��
�9���v�[vj���k�m�ɕ=�^�E�Jާ�z�͊�*�'q=ڮ�){�7{Z�ٲ�Gy]�z��[�[q���+�� �t�EP�UET��RHEO�  Y��)R�y΂���а��ފ�=z��x�T�w�{�B�Z���z�q�^����E�Q۷U��=׮�+Z��%AT��%)&�J"_   6��kG�+pZ�P�B��+��w���u���({a��.��n��=0kӡw��A��������`�+��U{$�֢��U���  ���s�nw�+m�<M��5���y�{tX����{f���p{���Z�W��k\�n�=j��W�f�U��  �  � ʒ�A��h@4 )�b���`	�10�F@�~JT�� �    �~��� `   A�~@'�� @  � &�D5"�� �CF@�h�OD����?��B��?��^^��#��}��ޣ�{����~w������]럶@ I�@�BH~�$��I 	$����!����$?�B H������Đ �Oq�H�!$I:�??���~���0�Q�?|d��ѐ��HOQ$=�I?|��:����:�"�@<�Ȓy# �=�I�`D!�@�D��<����<�ȓ�!�d�DȀy� �$Q�yC��X�� �0"�`DȐ<��Ȅ>FI�X�<�'��y'�$� FI�`FI�I<�'��<�'�$�0#$�!<�'��y�� �# ��y#$�2O"�d�DȄ<��Ȅ<�F�HF@�!"9FB�`9C��I#$!<�$!�aFI��c �!!"!�BBD�CȒ<� �� !�B<�|��'�! X�@�0�"!�@y"I �2"H@�0�#"'� !c$�y"B�d$"BHyC��$#$�<�������$#! h��<����`HD '���<� O#@�2=F#�$�"BHr$��Ȓ�D�@�0�O#"BI�`I#!yI!�B<� '� � O#!#	Ȓ@" �I!�HFH�!$����3ȀHyȄ<�!�BO"�2�$ч�y�yȐ<�C���y1�y��y���<�C��D$�<�!�2���!��>D���H#'q	�$��!<�!�BF�0��yCȳ���B��z��k�Ŧ���՞����;5���Zm�:�of�ܱmӑ����k_s�r%��=��p��'4d����L����Y�8�b�o�7�!�lkIƦc9WfS���:�$:\��l3�G�*�j�T�{����:N�ӸNc/o`�����Դ��\/`Wz	�:N�n�/U���f��IW��{�P�W"Ƽ��9���s��ܺ���:����b?#���P�;���9�j�у:��k�q�����s����t,v��R��)gt�84��h�ey(�y�uX--*���rla�ou�N����Ѻ6�n��qG��n2���ʭhY39>@a�L����MQ7�OQc�*��3���%�&ay@��'4�3M�G�֩;�(b<�QBT9��]$ƺdТX�=a ��@�6�:
��\���yـ�V-Ki�q���<4�����n�{��sZ.J��z�E�ǆ-�L��	�-8��<���}�yl1[�PV]��u=K��@I�z�<¤�״��H_b,��|.���}���E/�K���+f��w�eҷ��V��dS�&�6m�&_���5�)��A۸	���2��������4�y��v���an��9��6s�e���sz���#��v����\�GÍ�P�ĕ{0ͭ-��r,a͹Q�de�9h�I��t�;���NW؞�;�p���=Z��+�]�p���r�z��l�cRkt��ƞ�j7���թ���`�I�,�veY�Ni��E�cBZ�\��x���.09�$�(5j|w �w�Y�\��x�&�ֹVw%=�k�����(q�����:M�7�B��d�d��TD���өv��$vi�����'!���2+�J��7L�u�.8`�u���H�^''g`5hO7j�� ^��J�����R�;��+�
���Ǫ{�l�a�a�oʬC������l�r�tu�-��R.\�!�·2�`����ΥZ{x8�2.�TP��0�_î��;V\��u4�-}��a��F�&�=�+��<�hYCŤtEvS� ��3m.�*�0
�=n^��^�MM��&'�nl]��owe�t�@[�X�00��<o9��88�}��n������83�6�"��1�e�*���<j��Y�x���aAy8�"{��A4qWzO�-8�>٫t=�ۛ��=���<�I^�l�+��å�ًnۖ��{4s��q��7v'�uK0��%��­�^�oH�Uxb9���ׇ���Ǌ�j��Nӻ�3#���Z��A�א�P�0��^)�k�Ѳ��%����#�TػM3qb9Jq�4�ɶ7���X��H4�и�^o6��8�
�v�Lv��[E]:�y��u��*�K���\�(�r�:pU�p��K�*�Z�^�f��B꡻Z�yH�q�t��DqD~2T��{:-�[N����F�5����7���C:e�:d�;�f�{����b�C*��Ƨ3�Ky����H%e���E�y�7����f���6!c@��nk9VG�vkZ{��

���ui�6�H^�7"�3��ov���:D8�QL�:�����;�sC�W}���������F0��� �w�إ`=L|��vXv�ٔ�Yz�f.ٚ��:�VM����-<䲌���j[zA�;�����^���<��dq+�S���]����[�j�uܼ����Ӝ �MP��Z'$[�{i�c۹�o<�ȴ2���;ZJ��#��-��n��3rNר���ѱJg;�r��L��wF���n������)�S)��9�9��-�zY���W���]u	��C��sg<��}�ؗ�A����s�h�����N0P��;�An�ǈ�p�+��3��ͥȰs�m@���2f٫n����F��n�I�0�5�	����9*�P�k앨��V�ے�\e�S�DkY�]�+y�v���w�RB�g�ڜio�qk�&q����^�l����g�A��Y���+ۃ�.��t�$Xr��5<���X.�v�&n�Eh��t
^Z��pu�{���t��UG.jf��y�E�WY�إ�����{A���t��������3�Dy�x`LHI;�}7�ݕW����=�Z�٠8�^e��|l��a�'�rc挽e�J(�.�;[�8��7���D�8Q��N�{wo�,�`fAڠt�G,�����:���M�B�?���+:�=���~� ®�w,�&yd�zt�F<�b3��\Ξ�,f ���!�Uh�6���ot�u�=�k"L����p�,�˴m�4#�U�)hE�,9.C���*��R�W�Lml	��F����xN���׵vls��K�y���gV�6*��x[\wdDk|鰙��o�5t폯n��#�����}@���[�3��՛F���sS�d�-�t��gtX =ѧjc;v��x�OXX�r'�%�w@��V'����I�m3��L�u�v�Q6��V�g��kSB�HzI��geҗJ�RG�A#g"�ZD\:PtI�%���ݸ�e��007�S�ʹ���r۹w�nL��!�{�nr2s��:����(y&��pv��%������܉����N�(�]�W;�&Kַ*{��7��N�2��@���9���_Q�[���������Ć[����th��JR���t�]�NԷ�.�ۥ����aw{"�#��oM��x�:���	�b�(�/K���./	�]��@h�5������M�mhHu��������56V��n͚����ҡ���pI�$ P�[4r���6�@w]�N\�NC��.�d�m�]��
{
::9���;����pM"7����ku���5;qL�+�u����`�L#��XF���� �����5�<͗v���C��^����Z*��1�X�a�j}��A���{u�ܽ�7�m��t��,Ԓ��t=��gd��Mb��z��8D�wPyфJ���z${`�r����J�S!��	�0��Y�to8������\XnHq[X�ӵ�Z�7ye݁t���e�.oIN���3���SB<3�Re)����n���8���n���b'Cq]��t55H��>1-���r�����N4f�{qn×�&t����H�3�۩b�w�w[4��oНΨ�UnLN�.�����W]�񩕺8Eq����Ҫ,��c��,�7 9�x��"�8���q�KS�3��d�q���w�� ��\��P=��х7�jD3_Y��W�������x���k�s�T>\)�Ikk1��w�w����PM�2�Q4d�{�W�������8NI�E2(��Xxu�����\,�����Z�J8��B,�ҹ����;@e.�=/yr��2n+5��s�S��p��d�c�uγ������2Ķ��X;����U�ڎ^������M���ݳ�)�ڭ��s��w�f��6��ܧ;,�hݽ#�X��n�ؖ3ft��&vn�	[�\ب�
��1�0����SǋA����S{w��7U���A׾�s�:���.>Z9�p�S��#+}�v�v����^3�"0s���Cj]���{؆�*roG4�E-���͕�㈪h�\�h��in�
+���<8����n�Ls���m�'	��e� �7�ܼPT
�wZ3zMf�w�kd������s7"Ϋt�n�=���ӛ.���Pŗ���7�X,)��zy ��ӣ���[�m�%˗{�Yh��FM������r<��t��l�}�Z��gE�i�N��w!�tpL]2�͢���FU�as�g,�c� ��;�dxu�ě�j��x!�	>�o��|�m�jG�;�Rsj�u�U��Ց�;���G��Yǀ���Yr�彋r��R���@ ���H�F�%���V,7���+5�z����h�X/.ʖ��m�\�/���h�L�,�N���c�4��t��ʀٖ1�FN�iѬ1�]Γ&裳zk��6��J[_J�M=aW�d��q|�ś&rH� z֮���$Q��F�p��BE����5d��������ٷc;����^��p.\{x������Q$��V����S���-{��,D�&{���(^�5^�q�Ƌ��nv��E	{�XK���z���&���߮V�T�|(�<����z۪�'��گ5Q����b8�ܺm<f����#�;��jf� �K�n��t�	��q�����"̈T-�kk��3v��:�GD۰���a��;��L�9n9 �r9�jT��/l�N��Xv��,��P�.g�bd[��&�v�:f��t��W�S�]�HN�Zs|�h�uw"�F�Tʴe���t�h;OhÒ�^< ��Ѱ�Q�MߨDg���m��5�/]z"�A4�L�k�j͇;[�o�NK��E�
Ν�7�xY0��ȣ�e">�V�]��,g�n��j�1>{�7n��H^΃^�	2��fn��'qL����V� �`Ki��F�����pTPM��f�ܚ��MHQ���!���W+*/��~�����p���٨r����c�������!��|��I�&n�׈���{���
(&�.�h�7�'"� k {# ��cF�%2Y� ճZ���b����Ʊ�#b���gY5i8��okY��
��#��'K�dw���\	\��v�\����8��fĪ�p��~�A�g#9>�Qڑ%�K���T�#[�n�sq�C���巯N�<=B�5��ͤ�A��ְ��8 Yݷܻ,ky��X@�˫.M�N�nn�ov��X���5�o*C�r;���㻋s���友���>U$,Y,�M����9�m)N�wyT�͍���c�OQe5��]���8��	5E
����K5�;N�I��Zy4�d6�� 	�M݃wonZ�F�G0�>�r���;y	�S� 0M�6x\�u�[�gj�;��l���V�\�E�A誖Ll��FMi�
bۖ�z�4f��'��0�]��Fsrn�ON��ɽz�[fkTGd�I!���zY9˶�e	
�J��E�v������Q�Z��k�Ʊ��&x/���=O��)���H�Ŀo��	� Ίt�.�V1�:�j^2���BsdD��\�K�A-�ЫΥ�N��CPw7����w��@u-��%m/�5�٢ނr�+�>��n�^Y4��]]t�_Z��T(�Jz7A�+��)2v̓p���,Zp�܆Kd��ذe�Dg]��2�y����Z��U��{�G����5��'�C��҃^3'�9����iιF<puy�:ou�L�'M�C��n��s~�ֳ@�	�Z��C��zYN�ғ��9 �Y����$��P|0N�1uz�K����L������=O^�S[Ѭ�۵�7��Y׷��9�6E�uVyw	0�sN�d@��_d�e�������o:Ӈ����{H�K�kg$�Nz��W79kK��p�GJ�5���#*���!�׸M'v˄�WL�u�ݲ��5Q�������Q���v� 4	{r�Dv�/O�pn�8��f^���`R�EA�ǃH�+�FS`�����`���wH�,L�H��$�Vj��o&�F����6�����Q^�_p/B�D�SX�m���W]�˛��2sA=Φ�702��9�+7aP�٫w�<�Ň��.���U�9������)/,٠�6�-=:��Q�Ԧ��:�9�ʄlo(�.�=�ij���8�y�VnŮPl����F��J��&��s��cy�ZQ�&MG \7.���9i�G�D �J���j�r�S#����
%�ywv��=r8�y��ր�6M�g3���Y.��pf�v�B�����ń����JX�q�u�'I�,�ٸmYn5��-�� B4����AJ�陽V��9b��{r��6�ٽ�X��MH��-�3Y�dA�n��cɽt�@@�+i��P4��5p�㺊�\�oFdn��P\�Vcec4�,�b�p�O��E �~X"Ԇ��Sn��6����IFvӫq/h�1�sx'8Q�GD+B�s� \8�o�J�c�H�Ϲa�"�ކ]lk5��/�귻�M�M��-�����n���F��4�1�G܉��#�t8��%q�z�ɠ�9wPf�	��h�����u�t��æX�m{ݺ%Ulˬ�0v���V4k�Ʒl�A��IU��,�1Vre��:��'8c��WHGx=UGh*�bw�b�"��զ-k�/�콦a�yh���D��Pyy��ۂ<:���y$=E�����IVe�\7"tt�{a�^ômcT��[D�'g.Z�$0\�#Ὕ9[p�z����R���9+���ؙ`����.�8oEvh�;����ra��M [xv�9�9�o`λ���Ŷ�鿳}��;@N��q�w��p�)WV�~X��|��ivp��j�Jଊp�ك۰�xv��VH��.hVʐѷW�P�k��rea$�-�hl�w5�EL�]��s\o`�,<%fi|�(�=ۆd,#�gb��0R��9��|x�]���EKYoq��Σ�-tb���Q���i��R�:n��;;V4㨓I�ܯ�=�N�<C!�R��e+��½����H�pu���7'��
1%����"���X��&}�v,�x������ian�n�L�h�\���m��W#a� ��yJ���=��������^�>���I��g���;�����I�::�������6yC�t9�N��2sp��i���8 
��G��"�Q˖��m�����r�Ei�m����C�.�ک�QȚ��-�~b��c�sx	��o����z��V[�v�ck�ⰾ�Z�K����O�����B#Z�ʻ���a�yc�r������義�ܰ�D�\�x{Ccօ*&gF�q�ۜ����&fn����g��B�M����/��;M��`��]{�mpv������Ϥ�T���@oe
w�ս�7����gs�@:;�9��8g?�B�G��%�Nf�p�x���p3���;����Հ�&��k~����Nz���'�=�4x��pt�O����=L9�Dh���t]X�{Ɏ�����"�C)k�$�ы�Z��N�z_m1���):�FE��_����� ���E�7;N1K�>����sDuv�4E�%:M[9��(Q�]���Q�1mV췭˙��2��!C:��Me����e�/間?.ᎎ��b�#,����8�Jԛ*"Fm�D��:��j���$��j�Ĩ��si}B�Č����r�Kw���q�cs_�vX��eZ|0��Zԇg;/3��݃r��e@br�������Y|3Wv�N�2�n�5|hڅ8���b���<O�;�?D�ck��Iݪ�h�MUכ��W]�u���S��(�Ai�lK7\��P�٫�b��o��w`�%p�%y�7קT6�n�wju-;�bd������Z|1ݡ��^ؗBJx̖���,���1>�	Xz鹂��-��S�W���OK��YU���S�Y�8�r�w�M4������d=։����{Rs,!���G�b��Tz���Y�x1�x�X��`}�H�}��ͷ�O��o@&$�^dCúg"x�����¯?[�s��!Z�A�W��z��
KVk弨Υ�0P��ͥPfH�j��1�W�xخAj���4)>d�ț��
O^*�ڟU��ڋ,[M�6�s}ԋFặW x{ƥ�v3���{g�n��cJ�9�'9��᤺�	ǹ3j�=n��X�<G�����ޗ-p�S��Ct��-S"�BBU��q4ե7�;��nR��oz4j)��&�PV�[�pa��f�Q���u�dͼ}�G���f�����}J)�N!��20�zŇ�!��UsL�A�����ҧ���}R~�-Q�Jǀ��j��o�,�J����G�c� ���;[K<b�6�W�ٹ��kX獮��w[����&S��_*�\����m���Ң�����ν��p�}����f�$.R!6��Ιfe�*��G8b��.�%y�"�V�ɴ�)zm�4F�\>d*Up� ��]ٲ��G:P�Z6��u>ti���w^�vd�m��^���_�\��&�� ]%\�����`YE��yBUQ���
u6j��ʬC<nU]���T5C��.���H�xt�i֚���&^�t�?mò�ڶ�lZ,�;B�[L޻(%fa��� ����^����m+�y����E�y�Q��7	Ʉ�|�R|�y�nQ�7r��)�n�7�>����%se)C��/�nۃY�],Yt�#��}�`�@�d�¸.�jP���� YR�9���M<��ʈ��B���ݔ�D[�K���_@��+������A\�0�A��W�~��ef�A�4��f��'�OL��[�n�.b�k�c��7�9A^˥Xdս���!>��؞}�Y��v�����-=N@n��
�_fI�:�;y�0s�@ٷ�\�@cf�k<���< �
z�/�X�s��޾�b�7Y������5%:�Ͱ+v�ؑ�]��B:�$R-�<[��H��5���І\�eҭ�.�x��wo,=6]�����Msw'7����Z�1�}�R�����v.[nun�y�1�R�zM�,�c�t�T����;�������t�M�ކ_p�R�7`�`u�=��۬��m
9�-�.�q�N��B�'N��{���cգ�)��xZ�'*���F�u?�k���`g��j�Ѝ�M��:�x�Ԧo��y�B����Ú��$���l��-^�IE�/"�׫�뇁4�t���7�p�������u��Z/Lΐɒv���HV�qz����>�����<ww|E��Td'�B��ӧu3�-ɳ�X��$���<����טu�#[ٍ�df��2�m�Xv��^�#�z�m���b��t�׈3������l��¨r%}� ��z����l�:;Qg,%��]4\���f�m]��ԭ�qm瀨�"�[�K\���4aYֳ�"0r�7�yƷ��y����Τ�R瞾�\��UxD["��d�tZ�C�},{�kW/��H��$~}pe��������+1W�ּ[Bcq�0WD�s���u5�+U��ŮV��5p07P�,k���B�h�n�E�1�z�7��תt��I{;r�"剨4���kV>5������������Y��v&�oC�֑͕3%����N��e���ɰ�4o*)��kJ�]�WFwl��n��՚PB;�/(��W�+d�Off���-�XMl�$]�������S�:�OJ�*�.�09§X K��`]�x1sZotD,ܜ�I�E�:�t>v��tTB��]�u�S盫ۭs�M�١� ��3f줘%ǘ�b�ٛK,r*����W�葂�^�ͫ��u�[^wH�����BK�+fQ2?�t��O�����_Yq-ݨ5�C��}v{ܭ��=.��j6l���������U�h[Љp�,� ���TLӄG��&���(�E�n�=ng%������:,�6v<wݺUhVX�N��2��`��W����s�b�>/��R��==�_uK'(m�M�Kn�l�0����E�:a��n��|�Pe!���{���a�Z��������~�8��ۚ>9	��n�����t�5��{�#����Z��y�sh��<��w���C[�}]�{�W:<	©b.��I9�|
�E�NZ�<.���o�����1.�b"4A6�G��+�v+��wK@�4!.�͇/y��榚Z9n��}Հ�{�n�j@��sF��05=sA�@ci'`�
t����X��\��pP����H��`�J�o�Y4#���f��<kǓ�����١X���y���cй0t<K0�M�7��,6�'����˞��9C۴�I�b̭
���-Q^�w�8������Ior�-��mK�J���Q��8�y�K��)a��l7��F�"�QVг!8���ӑ����+���&߶��ۏ{3M
RWw�j<�t��F
�%m'}�N���Qe�k���ݯ�3��^�o�}���@�����oSL%p�,q]�u�T���oe@X��ϲ{i�݅�E�g�Ӻ=�>VTGye^&�RR���y[�3 �����e�ڧF���'S�g@���M�s;8a~x}7b��em��ݍ�nM"ȋ��Ǟ*��{!�V	1�7��ΕC�"��]݁
R;�\tҮ��S�5�YV���*�� >�R!�L�7ڲx.gs������=�3Nu��&��o��W�o(�v�{D(��u���>5}ik˷l�X�Yސ����5g��m;��|"�lu���	�Fک���j=2�:.I��{�%2s�(�Ԁ{oTy{���;WF��$2��_��{����8��a��ض��� ڗܺk����L��@�ā�ݩ{+ �t�|`�X�3����J��">>���E�y��ɪ:U���ط 8��<�q���'�t-�B6n�jU;w�0�L%���t��Uw�4&{�:䮝�>�jm����pۗ��J���zB�U�^E}N1�_
�r�!���m���XH�������w���Id~l%��qd�.xz_C�2���Ǵ[�=(IJqa���[�C6��F&�u�Y:��+v�nCԙ�%r��@�y�S#�w����g������fP��wi���Y��Ui=�Yc^�Z���\��O�l��;�{Q�'o��3uÅWM�F@x�1��w�I��{0�B\�]L#@fEiU��]�U��׆
"۷���8�C�	S�s�%�܊�$���_O>�o�!�y�K^w���\�o����]� ��){WS�g%�ݽ��&B�z�Q��-�x\�B�x���iL���0�J��HЁ4����kB��luN>̃��C�bf6GZ,ӗ��s�\�{�j�Q�8AAD�eln���Kf�����9�ǧO�L��w=W��k�=��6�,p�~ʻ���#HQ�ԧi����K�U�e2h��	��쁠5��-����l�,�[e��� Z[�8U���]l���&g[ݝz1���de�rڂ�h���.�ӵeϹX����@��$�f��#�軃sT�G=�J��nh���]dGz(G+0���i+.�� ���nBi���k�xB ���l�=X�f#W����쾎�Q:���ƽz��p&:h�ql��³�-���NV!(س��=O3��h�C�I�y�̾���i��vm�9D�f��h;뽣=T+�-��F�x�y�<��8�#9�H&\��7���Q�n���oe6�B�+�oP�IGl#��8U��U�V��6�J0Ч��J���$է{P�TH+GuHe�-�oK��Y��K�E��{�'w�"��۴E���Ɔl�,/.��1ux�J;N�V�]�k4P��g�Q3M�V1����m�G:"P��k��%�m��7����o������A��q��`'yr~+������YD>μ���9e~�p���M�Sq��V�
���\�gd�`[ܚ�l'��Cy��g.�;�:�>Ít�De�]�����N�9�d7�Ո˵��!���t��ʨV��2�k��*�[+�M�:e�|fS�v"���������n]��x���ǻo���Z� =Q��i��X���0�>y���7��}��^��o7դʗ�4�Aq�)�=�ܦ򴫾ݬZ���;�ӹ�cS����@x���b�֖���ya��ŷ���^�n�\���/��S��Q��[�1 ��޸�ĥ�5��B�!�>�xӜ�I��52\�J��3r�
�"֑]N�!�m��U�r���6����=��Y0��2R��h��8���:�rK�g��1�'yH�j�wwLI��
UueI�T.�6���i��ϧK�#�. �cO{a�o��u�����9��j���{��̮����8�9k�ަR�)fW�bE���ވSl���\N� �{�q�f��h�7���OMn� �p��5.�xYsw�Nt�eo;�Ur��(��\�c�F������~'n��;�ue����V�{��P��r��';�i������F{X����1���/�b��rT��F���
�!�w��"a=��
���DOu��d�u��Ө`��"��i�坎����x���etٍ�u
�pU��n���)eu����W*�]Vkz\�q��f$��_c���G��ҹ6yRP���;5��a��hB��^���ncjA݋���@*���:��b�L>��/�����g���T0eW{��;=4����D��A56A��Ȋr[3//WxΦm_m6y�)IK�����9Ӵ�q�xh��3n�"�ݳ&ڏ)���Б�d+�[����^���'��r�+TntR�\��Dv�'����\���K6�ܮ�(�ُ�S2F�o<��J7+��U=�}U�����bu ��::�.�s�w/�:�ҡ9�ui��B�CIKrc��dyx�P��f)�F��?h�O�\P �ӝ�f9�]���&�/r�{;��zMFv�K���4�4k8Ϝ���k-���fW^ooa%.ƀ�w~�B��?w.��n�#�8�B�����V ���^A���:��vf�#����|��u�']誹ܲݮМ�F�wp���k[�H�S���2r�VGY�T�Gs7Y�5]�-��wc�E�3���W�1�<�7K׊�rs�~�D��f�N;wwʫ:�ָ���{����M�]�@��X�k�p�����m�Hk՞���t�3�n)7oR���;l4,����+���F,_$"�aȳ�*�0�g㗟��up�UW�/���+��L�ǽ�2������R̖_^˗�1>�݊5���M �^�i�n]�5��뙧���5y]9*W6f�7�"G.�gQOr�m�-,�=|��R�?7
|s�Frwػn��c�J{3�N��V�s��OX��oS�����s]K�š�\��0�dĝ7x�(,yP�?A&��\��Ş7nُ�7���-����u1��o-;&�E�@���Y�*�Mv��*�՛�O<���̳ɟsM�8-��iw#:�e�Rv���V��G�U�ִũu*H�3�9({�gi���U�N�S�+��d�G���4����}8�>��f�8�Es� G�+��t���t�'{),�|+3l�}&��l��8E�S���vۜv���L��6h�g�:�5Nȑ�u�͒n�*Jse������:u�ѡ��w�*2�S�+Z�V�rh�jSaL��7���est��Ϻ����f��c�!5��ҟt���k޻�u7V3R�]{�@�R�u�q�qh��di���ǸgSp��9z�OD֩m�%!r��bG%쬫)$���)"�I0�$�w/{���0������<-C�y��/$�h�E�V�Ci�K��Ő�� 4l�� �/�E���H��?�c4\����:}v:�<T�_� ��jtM[Mk�<��f��kW��3]��{bX4|�2*���9�6�$ x��<�������P��� �u��z��'\������	$$$����w�� �������d�� @������o�O���h����w�Z8L�ʩC"� ���i�K�{,=u/��=�d�� �'����1�m�r�Fq�N(���`�vE]Y �(��=��(Gc,�̬7ˆ`���(9wY�3����l��/?+�3�Hy��;�.��̀�Vxm�����
�K���& aU�����U�G��ĭL}F����c7:�+�0�:��\p�2l��M��]�2� b�'<�p$7��Vdm43<�1�q�e�xy��v�T�&ˈho��n+�&(�哊^�[<9ıe���7N�M�}�dː@�IR��_,��T�ҳ�(&�8��6J��:��A�0�;0�{�n,��e�2����+�JO:q��Y)5�4�Jp��(���;�iűf�OiN�\K����uK"}՛�t���?�*ހ`��`o���E��7Z�e(�C/���x�wSۘEG��R���ӷ��4j�̽�u��j���΃kzp�໳�zҥ�����ҝkYu��U��������cU�c�z,��r�fv�/RZ�I7,�	V��X�y�A�N���K����	�����:��s���nx��̤�n���![�I�MЌ=Խ�5�J�0[��i�7�V/e V���ȺX��]W«0]ݠj�<'�Z���� �e��w~k��f`��개�����t���9z�,UC*��w=��t����|������8�os��X���{w��*��`�t�����-y��
&_M�{H���L��3է�V+�US*�^�Pr�ƀ٘�]�UV��6�Nc$�2Egl�;�B-Aeq�f��|kN����gE�qo�S��^���wG"�J�>�
���Mm���F�����r��o�z�y�"���v�ƺ|���g�{���MlP�1�^�,0/F2��oj�֋�IzT}�Q�����'$��ɾۇaŚ3�N�M��HG�Hw]���k�'�Kt�n�;ug��.O6���R�,�*�j�J�Aۄ4�J�q2��m�1#fu�J�X�N����o/��}E�J�����Bɜ8�ޟw�.J��3�E�q��;yҲ�u�uo�.�wˊ؆ufDi���5��8��ɻ{�)xڠ��]&^�}s/�O�{ڴ�X�S��d�Ao�o�`L\s4�2j룫ج�h�Q�]Myɵz�eλ��U{�,/���L� �`M�u$d��ۺ����Ϩj�**|�*��;�خ�*ԃ�c���;�%j����3��E8l�A�^[�Us�4%�"��W��3�l� �~>��;���ǰ����e�\�BS(m֛��aQ�Yր�W���3�k.�5������j�.tX7"��qg����Qh��v�"k�c{#q,&ijY�-��7�� f�9u��q(+Rc�A�T`�7�^��GH��
	-ՏXp��}��:�攧8��vҩ��";ʆ�ӂ�4��5�.�n�:��g���v�W!�AAz�P�s��A���>-�C������(p���w�ùk��R�ū&��9ym�j��C�̞�����r�Ox��-��6�KO7-̪�������js��� ]�3h����a�{I�2�E8�W%����s:�X�1b�x)��{�W+3���d�����/]9/���i�����{V֦P;�Zъ��:�c�ؖ�&�y+�]A�8��V²!���)�}���9�Q10E��r��o>��M!��+��e�;���-I������ý���������ٕ�����!��oJg!Y�et��\�z�k�2��N��B�:��aJSW�n�:n��H��yOr�F�gq��-��Ӆh.��ˌP�#wM�ݫ�ݪT��)�7#u�Z�홡�ߖ%��R�<�S��.�T7�ѲV�͇7@�+�My��\3\yȌ�S�y�{�$�>O:c,���!�k2���ef�����))�)�-Y�{���s��՜�M�i���q)�7S(P��a❸�������0��]�Kf��F.�9ٸgV���i�*u��t�V�_	��67�b�^�:T��%o,��ƦDp=�2F��X�����y|�S�7���U<����z�޳'�f��{�'�J���)���=	fb{����t���s_d}�s���֥�^��?8��t{:���ıBKc-fF�#E�����m!xp՜�V�����I���꣒��Ár���vT�B��ݞ�~�Π���n�&üL�3�f���m��WW�fА�J�����UY�h���'�T��*���6�g^A�T�tL��m��OɺBG�^ �m�Kż��Y:]�4���O����xR�s�wth�c�$���3h��Yu�=��bׁj�cC�M%�{����7�92c�ݮK/����fvV�˱.�Aܱ=H�q�Wb3�N�����]m#+3��{m�[�ڧ��>�oN�.G�i�_{��}���A��zE���3^9�]wd��5�w�"��	3q�u��ӈ%��8`ʻx�c���9X̗O�_9��n�FuNƚզ��*t�d�h�,,:_	
��Vlc`_���x�KŘ4����ʋ]Z���$��h~��i��K4��Y�^
�J��p�a����ކ�x�H<�� S�zl�x!�U���~�y��͏�.D:�� �Z�xy�wy���@��DjJ�^c�.��1��S�||h�UL�3�l},!J��!(j{�EN���9{AJ���f�Q��U�a��f��P3:s���ќ]��ω.�ٖ�V�t�0�c�vtV��L����tHo"n�6Q��(J���q	:�O�w�^ܘzS\��ԥ]R]�6k�0���T��������O�j���]�����w2���;l��J��Q.J����{��Yx�o���)
���v��S5�oveU�]�t8�|L���m��Q�jgh������ac��;P�h굿-;d^".cN�{C�ͯj߂�-L�����1K���둻N�\o��7V(6���%��fv_ԫ���/M����R>&�^T���3.��.Js�4 ���S�d��]XF:4,��;�Ju��;�ø[�͋���-[.���V�{D8�
0���P*�.�1��V<�}n�*���).u���h%��ځ���R�PH��M++W<Փv��j�1Ba���L��]!��V�Y-�VGv���+Yh)�
�:�Z��6���9�[����p�w)�/��鑕��J����dVT��0l}w�H��Ï;����/�\�q�|ft킄;L���;��2��TOuk؅�'�>�<���v��V���F�X��yՙ��7�97SG.u:W�Uq�5���{}��x�Y�ɵ������u��DgM�*�����nqє�7t0ԟv5�j�X�[��U�TKC��L�A/,��nӯ!�78<=���oj�88[�},�BЅ�tk���t��*�.&>�����z��DrZ�bt�ϴt��v�����5����Q`z-����J�LA���'�����4�5-ؗ�I:�� Fu��_L0�ub�#`to�u����O"��͵�.5���W|�%t�v7��s%{�žVM�+�=���^Q��ۂ����WS<1�Q�[ݺ."�>-̀n�E���|�J�4���`
-�I�rz�3�r��S�i�Iܾ�v�e�q��2���FX��ѯԎ��^<��B�fWv����jF�<F��,�����Ł��\�X1{~��g_fy<j�!�����/�_<���c�ӹ�۪�)W��m�n�sJs�����ޕzܥ`�5����:2ͤV^*=Ӹ-B�+�B���#/��2ɂ�bH1w9�-��ȁOp�8s5�'Q�8�{�,��I#�3}ޥ���ŝ`��@��ȹ�t&ؽ*̭j�`s����8�Z9�.I~�ѷ�2-��y[� ��W��{��"�X�r�Ź4`�����Of,��v�ۏ�gU�����!4Y՛{u���\e����"+��k�L�yct�R�}�\��|;�k�o ����F��ohϲF�_.ŏ-kǭ�"�������rɌu�O��Ei"k����f�ا}���_K�O�z����� '�c��{���p<��lR�k�Al,�V]�����I'`,h�4G>��h,��ݾȚ�àR���m�U�n�q���J�=碥�Ij�b��W����Gpc|���6�V�2鮘m�����ݮ˷��ueY�׻�{چ��_R�M�������Ë{��D��ƙNg4u��c� �[�.`�W��破��x��Y��d{�M�e�ښ�.��wQ�kێ����S@$ԫ٩�&W�p�5�&�5m-C;���5�ǒ#�u3V��;�U]��97|J7[��2�}W#0��$��o^ޜ�X�Z N	G/�H�d���r��]�Y�}+@|2�A{o�
ת�\�2q�K5G&��+ݫΡ���8���>��\
;�^x�|�W�$�\��b^��B5�����Z~W��~�`=����s����+=%acQnW��b�ȕ�{Rh��Pt:��%B�S^R��s\	��\�J���ǅwYs;7�oν��cy�7���oM�63X����x,�$Q���A�wo�����-��W��}�'�)rtnGx�回캮��h�~{@(k�K9s�;���Z�`+���G�w]!���s��Y�FI\*��a��޶�!�h��E�*���)<-�43��K=J���Y��+�]yǩy1�|Mj�ci�[o���;:���h��7�!��8��{��=�NC�3Ê������moR ��\YY���15�LX;�ox�wٯ��[b3F1Mc�Md�B�w/��i>�ը��WB�e�O8`m]�ȥ��7/z�V%"�@����l��D��.���ɷN�٪%���]>����|�+���0�����O�Y���|��$W(�#S�`�%pb[`��te�H�l^�#h���5�?@��s�Ih��؈wq���0�{��婪�;�$48�[ژ�wX�n��c���=��N���8] �͛Clܕ���3+UK��N�f�R�R�֜��CN �1���4���]͋N�}%֫�6����&���{�zZQ����$��kV���7��D'��~Y�VvDu���� �"���{�Sb ������)Ív������
�y7VLG7 �K1���E�v�tS��"�96=���^Įە��1}�++�o(}�k��b������]ƥ�.���������B;�RZ��(�/�ݙr�bPp����%�������JR���X�\�Or5`�!o;�7ێU�[xgI����b�v�N�x�ىt��EK�ʾ�+/�@w��w4@z�/���uz�{����Y9֒vЫNIֺ�$����zԜi}a.��4\ՠ\���¦����z��X4g:�X� �:�{�|^F"�f�9^LP1�{��������̱�U�{�u����.���Yl����bW'W�Y�C}�X�qSs������d�����!I. H������6�@{��i�:�fָ�^RM]�i�Y
/L�C�-���~>�/$���X�h�Y��7j��Y�s�z)��1�Ƚ���*ZI�[��{B�b���"�ʲ:��u�p ՙ5Z˔)d�y=��qjDwӈ�Z�]�/8�1�Y��Hd�fj�MJ4�"��i9��^Мr�/(���;h'v(fn���h�%ҫ�)�ñ�[u;t�rmgZ��r��
{[����Z��n��8Gl3�Nb�*�f�bl�Hi
D^��PӘ� ��{�*6>�2_h�\�7�)�瓕�e�>-�hu�7
4:�ڂ�-N
����u���tx�^��x����חq��8n%�g��76tc{X�0.��F��xvn^�g~Ք�E�DD��Z~�4x�C���cϢ�+���[�ήhT�N�p��Ge:�Wa���,�ӣP��l]�ب@��$�tu��P'��3�kB�f8��~��D�ŕ��3�9ۓ�����r�#F�"=�ɹ=�߼{�f�'��FH����(�J`;I!h2�Rs�r��{y�@����w��.5�_7P�ܭVg"^Y�ҍ�Sɀ	�bE��������vEWO�ZQT����撽�,B��{z�=�n��w�L-�^��/	�fvV�]�6^�@7��AMp�&���t!`D��c-|�����e�1,��	\ہ%os֟T�o����wݤu=ۣ��N�|k���˧Ԯ�˛����f�z6q3��F�Rz]����f� �͆��}=`�W_���E��b���;�:'��%�B��!JnV<���t�V�GN'\[s7,���Ά����>�U20u*̄��(c<|�$08D�����UXg����/f�W��"�P*�eĲ���b��6çڏ�x������=_Z1��"�j �����ܧxn�3��c�b;2g����te�܅f�e+f�B�q�f��1.wT�t1P]N*͐7�֮�E���ne�2L��v��ãT�.��
�#G*��YI��ydh`��k�z`;��he!��8x���V6��i��y��K�&`}aM�w\�[�����F��V��=Г�-q����{����s��.�$�;�h�\6��.Rr[�R�E���C'��,�}���3�wD�kU,Jũ7\���$aW4��X�)��{xWl��e5�]t���J�jU�hqE�����6� �C�(�������ݽ}�*��/$:_V��'q��Cum�3���_�����B I�����_�����?	���?9��?9��u99?2~s��,��?^���|��ﮧU�((�Bީ���`�;N����e�����5zMO4�Cܵ�2��vv	1.a�(���<L�N�.+��@R4�-(}�;}i2x���Qܒ�w`gc��eQ�V��)|5��	P���%M�l��@�����t�,�Q�c������r�uD��kGr�Ψ��ƥp�kV/�D�M���=�V�mn���-�Q.h���:!� _�g9�����g� &�&C����oE�8��r1N�.LV�{7/���x�{�Q�!q�ґ~�x[�zT�;�>��d�O�p�|}��~�=��y���,@��c���_ݪ=��;j+��D��u���n+9h��q��Y��=ޮZ���ڧ�������֯n{�+=�������yZ��,��R��(��W�=וj#F���7��	Mm.̛G*Q�4(}|m���dК:7ۇ�� ��Mk��x�w����e�����z��aw7��4���Ի�R:���NӸ�pԮ�ƺ���)ާ�e��/�r��ӷ����㷢��w9�'�%��K�B�k�B���>x�[����g��\�4=��ޣЈ�$��i]��'�ӮC�0ônr]���˘�.����}}]ze��Ĕs]	�ԧ%�CJ9'M(�0`�7�^nY����gP ����raZj"6�����m�Fڕ�˾^km�V,ŰE�mK(˒���Uz�1D�,�QY[iR�+U�։c*��*V����P�V�MV+�Kl:sꛔyXµ����Uzg�ZD��U5m[�\�<M5�E)R�V��J���6QR�h!Z��S�L��`ѕ�JU��^���+Q�[
�o˅EMJ/hP镊"�yeK��c�ڂ�b��J2�s��(�n����kmD��j
�˜ ȜM��QDb���c�QF*��M�".��Kx���f)���ڪ��(�m�!�p����\�"��ͮCR�k*(�,T��56+R�j�S������k���U�l�ZJ""�ͪ�i�UAJ%N�.*,�X�DN�Ǒ84m��r�q�%�kD�V��j2ѵ��Z���-���Dc��2����Z�Z8h)l����\�j��EJ<r�Ussu���(�m���o/5*�
ޙ��6h*��:�YĢd:9������u�α��0�,h�e��8E�m�}������	�[[���'4ʞt��b.��:�����e檄����dm�db~�̿����v)��?�(��l��n�ꘟ�J�K�w�>=�ZRw��x�����9]�H�'j�=O/���֐#��H*e�כ�Dre֖�x"���n��e� ��l
��sTGt��\4�����=T*�M�OGH�v�m�j�/��9��5�t��'�����ٗ ^;��u������q49������>�hT���Lѷ/:Uݚ�4A$�����L���ύ�m4��P����]�蠮,���L;�4{�N\���z2x�g����'6��!@ǎ�O]��yyΆN᪮����Z}2e>��s���O>�֏��Twb���~5��Nۮ�H伟�9T7��LH~�YK���{�h�_����{W�bE����r[ئr{�91���_�%|M�;f/*�`�ܮ�3Ԍ����^~�f7� ��ŘͲ^�դX�X��_��L��go���1�7�íL��h3r�φ�y�7�!(�(����]AeZ�\���������js�odA�J�j��+��+hK�E+�,�$u��[
����.L̹&r��3}��z��5�����\yAn�������Tʤ�k�k)t��}�����'�x�\�=������s՚��.GwPƱ���_� E�K]:���z��X�*OE	Wr6Wn��R�3u��گ�և�p���\��X�Q�B�މ����L,���u�\�}*L��lk�I%��x���h_/�ٶ��w���yLy����	����7�������y��=���u\��i��;��ݼc�ym^qZ����+"����O*}Fo�0m�1��jz�l��|g�8����*�k���*m���*�l�4���*�;Xz�+��j���;��k�SǕ^<�_;�Ov�o��D����4Q���G�=���L}��n5�3�d��g��V�&{�r�m/��;�ql��M�órL�	��/d��H��4V9:Ǣ3�?uW�{�+j9ةh�����s��N�2��q��{ƕ�F'��}h�ԋ��JZ�E���x_�8׽�|{wK:��|�
�Q��}���6��ӳ>u^mf(�٦�;�C~��\�ږ*��_�ynv3�S��[�9e��gCb�!(H�{7�|�����c�P��-�o�,�{lp����n!�]�ێ[Y:�_��t����礿OW�jϏh9��Iڊ�]�d��n��@�d��'��;�F)<�p���q/'��!��jbW�1���$�u�`�mF�>)�kUg]����+Ԧ]7�G���2����O���C촺��<�uk���#�\z2�n�qA���a��n�F,��}ț9��G]�,Zx�=l����8�2�8����5���c��֢�:#�����������m��V�w,��V՞ǟA��ƃ�����kF4���Hows�o3�xT��|�7]W/��U���|m�k(M�Pm�2ԩ��1d�w��׫P�_8ȑ�"w��7��-��Nu�&t�V}�-֦��S{Q�΁7Ѩf��
Ҿ]j
��Q�T��1�/;�ʺ��R{���e+ވ2:�h�|�i��|1Q�:xa��q/h��c�6���]IÑ����XQ�o�ž����GJB�������Jy뛮��W�C��;��\�W�	��tRn0���[�<���	P�KFs�6u?�>ٝĿ�b#ͪ��Zq%9��e.�s��}�չ���e��]���!w3#��㣟���KjL��3�3���n�_�N�X��;�0��'wǹ����o�c����P=M�I+�c�����7uH�5�7YK�ݰ;��`�-�Mj��x�-������^'r���d6��U���Ɓ#'y��:>^bgoz���k�2������4�+}����ȯv�qyJ����h�����I`���XhU(;-����_v�z�<o�d�1:���v�ތދ1���k�do���	絒�ߒ�mt����}��v����z�>��կ�s��Ř���a-Ӏk=��e�_b�m����v^욗E�v�'��='�����-w�]��_��	�U�U�D9���(&�u==��)���wO&=�l��Sk�ͽ�9�Y��W�`��	뷊�@k��Dwd��ޝ�Ö���X�� D����k���H'w�F,�]n�ݳ�ʮf��U�@Ó��h�l��=Z��I�m����`���)y*u��ވ^ۋ�z㹊I��NT����Z̾I�=z�V�%�9O�3�_m6�8;z��Ⱦ�p*��`�Z�@=}��D����΄�e��kO&h�3u�����B�zw���	k"�6��<����\-�q��з{��3}���qz�ő�TB���B[�P�_z��O=�^�+o��R�·K�yM����l���ZR�ҫz����0�TD��ox�l>�2�tv`�]��F���3����*ЭF��vSd9��on�� ��ڵur����;���
�vQ�B���c.;��b�*���u��_4xw��x�3�j��ԯd��-s�j�S+w��x�Z��r�e�z��第�l��v�=���i�W����g�.Cz�?N���}ؖ�r�n�@��3�z�����2�a��U&{����^iu �w�.�si_U\ �VR���3L�9���p���g���Gu�T�[B�d�f%щ���+�{��	��{�B:�'�C
If�d{s��i�q�6�.nm�o�k�=:��ÄC��{��L��2��s0������,�w�ad
�"�(x�j+���y��2�@n�AL���dK��Lt����ݮ�r�$ձRڀ	���F��eW=�o4$�xk��o.��a��m���g���7�o<��yE!^��<�6�eܐI͡�@����|��4��9Qg���sݓ>}�\�k�~5�'�{�2wd�B|�%Л��nfQ�������x᫺�w=�+���7�~�䚸ݝj.NwC� C��p�v;5���������puu`�i�hJ[w�=��Y{��QٿmO�����M���{|�Dv�xޯCi}�����}�.���>~ٮe���RW�M�+�7����.����a��X�>�}�݇�����3�dϹ�
�"���?�ճk��HW�^/<���9}�Q�fŨ�ѻ��C��A%��<�Tw9)��[Aщ�L���{��cz�J�'[3�:!��}�]�j;$��L��:�e���1:���l	ｶ�!�(�sOd9�Q��9d=�#�������wi���Vڼ}�ɟ"�f�6k��GPr�{tٍȫ��b�Z;æw(�\���}[Y����d>�����!�*��mk��鑤ӬS��3�t���N樊�qj]E}tE�m8hգ�:^:�|��;6���|�����R��2�>t;�{H��d򦮴�S&��k�{�O�R���޻��s8Q`�zw�r�7�C�Ǩ�N\=��߽���cٺ�N9)�������'�{'Sg�/o��-[<x��\��mM�(������� 3�βW�]��73^��H�r�M㳛�u�:��-�5u�N�L�=�w��Aޕ��߄�Ze�^R~�������{��w���i�]<���aJw�n��:�� φCCr6��ێ�}{���2^�yX���V5+��yj��]���2��,��n��<�܊-�3��ڟS�ث.h��u&�̓E���쿈�K��.���G�\%}��x��`��,��p<Z���՞&��9�x�'�g���o�����):�j"{۝������}Z�Z�㕷����k�c�<{��n������t�/^k�NALW�K��G\Yojk�s��#%YӑV���s��܅��֘���������QǲS+B7s���v,�As:E�-g{��h�|u��w��X1�����×�(%��s�͝M����p��_a��c}j{ջ�C�)#�c�̝#�NkwU��ʻ�5�'',��̓hE��=��9YC9��W2�p����}w�T�ޮ�.O�3Pz�Xv��i�(�Pd�]�b����|��<��1Q�G�L�Le�UL���۬�}�k�=��+���\�^|���F�=[��	�j����竹
��7*������Vv��߮irS~��[��j��M�ޱ�a��z��r_	�cЀ/�q��+Ӕ}^ͣ��5=ڽ���9�1��V*�xr5B��ӛ��C�}s/u'��hy�5M���]��>\T��w�M;��FOC��VNt��`�@�%��y�	�p�e��~���NX$�P97�t��������u*	TGw]�Vv�Z�8��/���v���'0^Mz���[#raIi��23��}ٱ�j�
��*��=Q��\}0�1/r��'��vݔI�Bt�E�׽J䷡�ߞ�l"�e���p��`���^m�9�LХ��MK3jȎ]�P��ᡋHX F8��Tu�:r��3�V��bz:�ʇn�"����^����oE�t/!�$��O u{N���U�u�$�IlÇ�C2�|�f6�ވ�y�_�<�nz�]�����~�8y��.�X�y�m������	��a�"zG�ry^��J�_P�&\7�N^x�=�=��m�^�j��"�8K��G�>y�^-��7�;6��S�kGU��p;\�����rW�E�Z�~̒]� �.I�����`�z|]Y*y>�d�G�Yվ2�l>+��k/Ҫ�߳�LÞ���nMSe���ZU��짝��h�˝`Pz��S!U~�+A^]F��\��yj/wE1�����	��j���w�}/({��i}�M�3�F��,QR�ƶ��o���Y�����#��Y�dЍ2�c�qZ����S=jrN�f��ύ x_'�J�j����OtR�\Ge�푄V���mނ�kM����se���Ɲ�a������[=��7�x���o��^�.��Vܧ�{b�z��d8u�ꫧ�ŋ�Z+�)]-�����Y$��u1	�(֠�v��D�}���J/:7M3)��n͹�h�����N��V�ir��i�ս9lz�l�a�]��\۠.�yb◔� ~�ag;���b��g��n�ۼq[�(H۽N�'��P&W�zF��#��_=nɻA��<yŻ7�F���ӂ��p҅��f�L��*hn1T�=�xS��3O��"�=t=�.l�Z����m��ތx��i�S��b�E?���J뤮�˽�Z��a]/�ޛ�h�Ϳ@i��~��S���͙�A��wbl}�-+���}�s҇�pkF��ߧ����^Rvj��k2�J{W56z�=���ɔ��+K�<������Lk|�k��"���N;��g�ju��t��vG׈�}u�M��a�g��]��@�����Uz��m����G]����b;5%|M�,L��������U�ݧ���ot�ꞽʤ�?^ܟ)}-��^��C����Ȍ�ogy�,�ӽ������c�&ސ�#}����@3��Ǜ���z�~�w������^#������ L�^�f�su�I�'c.o���� 9���;����r6PKA�	��ӕd5���yZi+��h��&7��^��	�n�k��-�� )�V�1������ڼ���܄�z���g�ů]�CA��K|{@�����C<V3��)w0^�;7��0��v2�WHs����/n��-�t�	-w,�4;�'��ؒ񳆳��V�zl���{��^&2fu*�{*�|1�O? ��� ���~[�]����z�&��Ifi(q��oՑx�q�>�)�N)�e��%�t�N����*W��G��G	h������{*���j|,��Z�pܱ���C�*DR���v�:1��\Y��'<��;j��[�x΁�ʰ�-t����ŕ�'�!���"�gz�鸢A����qh.-�/���n֗4r�|���|N8J�܂SX��·XZ�>;�@mi�v�����p{'��<�����a歱k�.�����w;AoA��TT�:��j[S&t�Ѹ��b�Z�齸|�U��T�Gv�.e�ʽ[Eɀ�6V��}�n\u�k������-���}�ɍ����q��ZB�@�H�.l���f����f�ϵE����p�ܬkd��O��D�)�$gc'o�Q9ҕ�ȁ�j�M���B��~���k��j�ݛ��3׺<갮��w��/^B�j��t�zX�I�z���gU�Bt.�/���*
�Ȓ�y�bS<E�˲�œ����bڶd�9�g�jyy��k]�غv�B�!��j��dc��/�^;��]���=�g�����4�U�q�n*���{8j��w����Lj�KE����vXˤgb}��(��F�^��ʭ�G;��(��'M��_T�΅�p�o��7���Fz�V�<�[m�H�8�i{����u�y�- g�v.۠�֮�v�uo�f�J�4���V�ͱ3v����O�S���wq�����o]#�� ��k��S��|x��k��!�xF'!'$=��(EV��]oc���x����]�.I�v�#���[3˾�'I��YQ�ޓ3#�:&��m,���\��we�d܇Ԋ�<��dy`p���w2۽1����Y�Tn<1>��͠�DK���3u�ׁ��.��Zg�Κje�g�
9�*J_g1�✽D�=��Ƹ(�{�n���%h�u�6E�Vef:���k�!�����M͸Wr%v�@4n��t���s�>dq�x`�+��vST�C"f�N#�
�݌vܱ�#&�G+�pbxG�va�� ���WP�[�x�>Y�$i8�vv�ˇ=4�G�9"��!���s�07��R�y[V���_44�����6z�ƅ䟈�e�J�[,�-�w�l��dr�x@x�x�t�Dy�n�k�ٞcا�qz.KUa�$ꄾ{W���kjz��7$�����74h�P���ģ�R�]��*F	�����E ����ι~��EADS��h�Z�ѵ�YZ�Nӆ��b�n��1�*j[m����h���)ěT�T峊���f���DT�j&����V�X��*Z���ʨ�:�r�""�JڕN:3*^�����#�Z�,Ǧ�iEii[j<K�R��\�L��\Z���N�x�]t�s�%�eJt�����ޞ:7�;x����ėE������Ns<��z���KQ�����5�����%DJ��lٞpS�3hU6��"�i�qV%���[�5ծ�U����[.��r�ǔh���ˑ��M��ef�\!Qu�O1����N2Ķ�YF-��V'�UD�"j\�b�sS��'F2�Z��1�S�S��Èb���Z�Q�G�KW��3��0�֕��u��ˋ�K���[v��\�����Vڶ�.oprh��K8%��)+F�.��L�j��Eyh�9KĢ��u����e�*��꣭L�fa���K�c�{�r�VV��z��]J�+�-�J5qJ��U�i�˓%�h �j**�a�X "0�B��(���Z�ꭾfO���q\9��mj���fJZ��h*S�ܥ8��S��̎|��=Wu��fs��.�Pg#��q5t�꿡�o_�	�d����̍o��Q�w���Sa���!�Q^���6,geG��Ib�����nN���hC��|'�b�~Sd��2������^m�g����Ӈ�����S�ڛb�ҧ�0c��p���N��1F�*?�\;V:��g�
.�e��Cߏ҃m#.��y��uS��r[*�oi����Z��ɿ~�*>�Oʖ�*���`ɬ`kqM{��'�~�.a>���fnnlp��`>�ߋ7:���90�F(��>"��ʾVK=��J�"=u���n��3��N]����N�;9������)�d�z��-����5N7���[���Ч���%�H�%5���+�Y΅5����m�g����x6�;���Ϛ�����l�Sx�`��}l�vS���Vy�BQy�ɣC���+[0��h�~��v:֣XwG�.,Ī\��������,�a�@�������4̈ѩV=n�����
�"c�3�Â��G}Qﷵ������dC�5����m ��*�(�{+���n�Kv]��f���t!��(��Y�?L2�i�z�xTeid:������g�����)Ix�w�7�\(����\X����S�{8o��B.;@��|�<)�Z�6<��r��/=~}e�;�O-�M,z�v0�o��W�,��P��$y�#�0ۤ��՝-�)'ۀ)�a�E'B(�{O�c��C=����w�P!J�S����觻��{WG�j~m�tCs��g����9/��yO��H�~�R)���:C��n:l
�ėe�GLw���v_�G�7C ���ѤH�F�S�!�Fd׻c;p��EZk=�ck��<������{�~'����[<НfǪQy� ���^x�l�ZXY�G���WHg���q�|b�o�z��N
0{:-=�#�rh��k�;V��u���@P���"G;R݅�qS�� vl����3w����/�~e,�;�q���9�9/���VQ;˄^B�\~���OV��P�5�3���������Ɉ�L
��PBFt�W���ی�&>y���һ�}u~}g�w:�:v���{�������<�H\gK'?�,5o�&�<Q��7!}��:fD��%�]0�ӼŚ1��Yg&f�7����u�9Mê��j�E�pk�T÷�3��X��}�uK���3����C������K��5��^�h����(?�Q����C��r��;Ref�{[��o>�Sl*��Ϻ/[՘��UȜFm����w��H��c�xeTs�)\L��\������3ou�n���7je����"�֝�`,��-~W�&�����y��<-���6��sP�zZ@nqԂpX����z���+�|�6Tt�Zܾ��T�Xr
�i ��jӝ
�w\�h�P�.�j��FO�@"?)����#��W ��ߢ����L	�[���W�>8w�/U�'�s}�B��n�S����� X>n���34�9��uF3�`i��Y�?k�@τ��kĹ���F�c�"�`��寑:m��c^�VT��<�-�ϒ����P� �۝{w�q9�#�C���.��c�5��(����#dѹ4����������(�Z��"�xг�6����{��-��ƟC�\P���B�I�̐O��{2���é�t��`��b���Ie�:'��+J�ЉqK3;��X|6}0u�Ѷެ�]]Z�o�	��/"��pɗ,ڮa`�%�/��ό@/������D�#ݭJ��n����.�Ѷ&"ܵ	�%��{�����T�ƭ���#�����-XȰ���vQ�]C��陶G*H`f��L0�)��z�@�@��-�%mJ:*�G5�%o��uM�˚s�q�BX�� ?��0�=�
��!I�dH��HG�\�lhu*����p�����oW,�y�m���׬a��xe��0��0qϑ�Ts��;����T��|>�L��o�}]��6.u����>˗jlau*��E=l<���G;��s��12xI]j2�녌��^=��:���v���u�+O<�[8�L����\�n��+�=���g{�Z#n1�
܊>� w�N��UҬ)}�u��u#n^_�K�� &葙���*��4V��_�~��3�mo'��o�`����N�aLy0q��l�>2��L�JJz�nf�4��N޽UQ ��xË�E���ä�/��Csdq;��d>���������dl�O6�&%ob��¦��E��-ݙhl܂�^�P�m"�'Ժ2S���#�`�Je��v\�_5�^G�*��T\d;T%5"�h���=��Bi��X�UЬr�n������z[68�&%�eD)���!+6O�Q�:����"|Z{�V0;��~�'1Qj�
����sFT7�N���{Uo*!M�Hj�f)J����n�r<2�E(H�3J��k�4��η��S<�p5L���۪��0����J�&�dZ1��8�Y]ؑ7
�U����2(���/`�N�%0�5����x�$�m/g��!ig�F,�/�9�G���μ#���;k!8 ��ݑ�#�y��j�ʂ�;�>�]�^JV���=JC;�o+2��FU^E(s�ú�>�����_�ó���C�[�g��W'Z�%�b���v�h�b���OFuq9]��5�0�����M$�r�p��N�#���XY�'*� Y�	:T�_T� �S�6��\��H.L����Gl�c3o�?J���(�e��-G��P���V�{�z��S꡺�S��B;N��qE��Ꜹ$oN�F�vt�[lq�k��}U�}s�����B<����d�1}�@�I3�T���u�d�������kZ޵�g�7�6��u��>�備?j�3Y_F@_��-�,�>���f�.GF����t��]�h�wO5�/�O��G��5�3bw�27�����w�1{��4�����D$���z��m��h㠦�kW�5P�tǲ��Q�*J��oK�`�<>h������o�֩�Ąשud�ΆT>:�v���^ݥn� �z���x��j��X���7�{r�Դ���=\�>
����7\�%��yX"�dne�7������207d8��3Y;��w>3e8��jR�! 3�J@*�A�q�V1�ɯ0机˸k��moW��,���	Y\ko� �������%����C.|�mť`J*�!f/��T&��dn7��<[+g�QQ3]��GR��|��哩�܁G7��1���2��|�b�U����e��E⩌5-�"�����
��}˾�ja�X,�PY��ʣ��n~æ�k��w "������>��R�Yh��:���=ܻJ�oU�)t��<v;��Z�U�J+�#�\�2E�o�����V�X�.r,od	z��V��˹yg�D�#*Vw�Q��oL�ȯ�=�.S�*�|����u�F|%�<��\{7}pu���xgm�F��uq�YW�6�K��a����ꨏ��>r�Ю_�֑���x*�q��?�8��?:�>����-�E[�����m��%�H`�wp�Aĥw]�:X����ԓ�b�SҎ����������N|����Z~9��/�e[xkdS+�.�z��]Q1C�M�}�I�%�c��ȵ�G vuAG����ކ�k6˅�<�Za�;�Tw4*��c��nLu>�Bv��
!Y��W��3�8?��|S�q醎���
��cu����,���_v�P�0�{�,x��:F�=�������_��9��mVs��*Z{y�����Rȕ*^��JhN����?��&LE�ج�0��0|�C�yo�ER�T��y��ɪ����k�������"�����hO^+z�vf�O݈�?8��0�6 ���S��l�߅���p"uc8l��B\QX��zx��Ley@�J�cRΑ^�^�k׸ņ�猬�U�oo�Ϧ��H��U�FB`9-��]c�x�%�7dqg�w&˷~(�١o-��<H�f"4���(5�~���gIP0�>PB�b�2��w�-�c�nd��y�K�}�b�NQe{lߜL��)Yg���V��6�r/�9�2��z�̽ݛ�������y�s�V�b�-�V����m���=ܧO r����;I�OgZ��Ή|j۬�b�W=kT��TѮ/n�m�A���Ģ�No,�(�r��u+� U]m������C�40h���xx-�x�<tq�[����Gy�pћO���Љ�ҡ�,�s�LLY���W�5(qN���V�z���=��f�O�R�p\ ���w�#������.�x�7�xF�^�=uU�c��X��J1�w�P��y���r$�|�r�sp����5�o�t�ay�7w�Ž3��3nX��SsD�w���L
i�4��(V�~�"�c��O�p͏)�̩z���Y4ѯg]{�}Q�I[X�����tK8lwC/�5-o=��}�F�x��k7�n�o]Y��cn��RKjM�;.�4[z=�A�C�\Q��]���_j��r��3y�J�W�s����q׮�V/^���dod�3�`�	��J���,�l��!���fP2FK0'��5h��&�mo9x�.P��k�y)�M#�6ę̘��t�Da�L�U+��+O�ǽ�ֳM�E0T�ļ^��i����wOa�I.��q���^!P�r$�V�0��Z�z�^����6Ն[P��>4��QB�q�$Q�Z��Y���9�,��|j����OgYԧ�G�q�u��/����j�;ػ`w3����g1�(0�@��j�u�֏U���,ve��a�z��m;�m�� �V���Ì��Jx;g�
\��I����#�\��������X���6,=L=ݫA�+v)84H�i$mQc�ww���� v�4d�s,�3G��,<����xF���O����\�	�E��c݃����*T8��-��y�2Ғ��nu��cd+����ZPJj���t��h�S �	��&cS���S]Y�[�꠽��z2:&�{�5௝�w�mz|�28v��;Q{c�	P�
�dO���4Y��\{#�[2J]�Hv�!v+)ޠߕ�3Ӡ�}/���a��`�@����8x<pG��%c��{��
�F9�{θ�]<_��T+�BA&[�f�)aN㐑�_q�����f7|dm��7�ך�ӛ8ՍGP��2Q���+�G���Csd�5C���W������o�y�j�O��@Ţ#��%ʯR�6's^Z����@���=�h����{@�X'�x��j���#��������б�P�ܺ=:�Q�c��Y�pɗ�%�L75!E~�	�(��]���{"���ڈy�|iР��	F6A����N>Ẽ�>]J��)��OcO��M2���qx���o6�����X�r'1b�&̞�W!��}�hه{�(���'3��򣷉����7�	�)JR�e�ᆥ�NKB���j�Z��sIp"y�:�NQvF
��z��Y�.�ЦbW�=_|b"���Z	>��)��o�"S"W���*�8@��ʁ��rv��|�������=}�8�@��"�zj�s�N�� ~�(�)��q*�E� ��cc*q����!��;�G��r&A��	p���n�%�0�y1�i��"8��_L�t�#R[x����8���ƹz.&ߕM�-%��Gs��T����\��O�3Ցd�)
{=O�Y�TS⋛/��?6ϒ�����8��3��)�AL.�[@����֚�\]C"YO�u\��a;B(qU�ӹ/�����Z	��z�Y��Ψ�AY���ی,׊\��0Q^�=q"!����N��u�f�u*���M/�`ᄻr���C�������Gptw�@�`.�� �x�2��O�*F�Τ�&�TVp��S&aS+%RNw��P+���g[�T;
4sJ0/���b�[�B2�ޜݚ�C�:/E�m~�/d>�g�&`���?=�a�Fi�SИDW��eqӓQQ���Cnl ���69�v�l1���@�iw�Ǩh�h� b(40�CtpX�,sm.���m�ܻO~��>�8�~��Y��+ _m�����qQ�&;���OB~X��#&��K(��V�5Ư�Xú��n��?��E�$���r�N(롵��Q�$(7f@̃Y���fn^*�o	j�qb���G�I1]�G��Q�5Nd3r�c;��R�a{֤�W��m=.��Mr��F�Tw�  *��f�p1B~�w�7�j��t�p?�B�ZPp���\�uu?kNd�4���n�I�`֫�=W]�b*Q;Ԡ+�j��Ik(F� Q�����ꓡ��l��}���ܚJ�]Ӈ��/ ����x�,����6Z�a"��$��5ċ�;�'a[�p#l%e�;�$�'��Y���ۥƯH]Vm��}B��f��<�;m�i��!A���'��o}#]Q-�s/k>�K�D*wk��u���
މ�7��fӬ����*o��AU��ބ1V�9�N^Y��k�z�y�c�������Q�^)�B.���O�t��yd�.D\�f�����Y��+�����]y�1�Ǚ��G���q���u�F��n�l$z�BhLZ�/J5mK����k�F�u�ra��u<���u
��	P�T��@���P���&f
r���ٟ
Uza�5	:����^ٌl�qY`�7;�"�c��en�e��Gy]��ǲf��jWw��x�B%�L	e��Te̺hO�.{g����? �71lF<B�>�g����{<}��W������~#��������_��61�pT���Q�.���"��LS��pbp[���&�v6��kS�+�����&�r�u�JV���B�ZO�������e��E�t����[��!�x4��N0?�H*�I��g3��M݀�s��S��U��
������\�q;���A����eZH�_z�Ɔ"��ԪA�Q�wϖI�����Eݛ�ҁ���G9�w+2��x��q�-��nS�LU{VT�9DY3ѿ_C�x��J��wh�����9�T0p���-��a�bn��YBeFL�h3��z�i��Y��:��3!G��e��r����!��Ո���%�}F��\Y*��oT��ǸsóJȷ- �:����Ŝ�b^�sA厏K��5w�-�����g��T�Uɦ_��\�$�(鋹hU%��-ͪh�>�����v��kQ��ݸ<q�R�?��瘾~7���׆�֗l"N��$Ǟ�f����\Y�@s�YBZ3�*������v�:\.��� �{��4{�֠�zI����e�y(��ݘ�]n軶�w{�n�
�"0���h�?ca���1�۽��lYF��/����[E�؇�T��tv��G�팻���+H���w�5h��4�tֽ?K�<�4����V�{��Db�����7@�ܪ�xա��=8�΀�ι�Viz�M��좙Uu1��&n��2��Wr:Υ�S*vK{Շ�U���\c/R���{k^��zj���b�z�V������û6-\��J�6��)�4��H�Ue(`~�������n��7�����r`�g��
��j�&(�y���7�9��b��F��e�ٗҋ&���A�b"r�6ȩV��Δoz� d�ޱU�-�z���ݼ[}4���o�i�~�3P�S�N���}z�u,�׌c��52R��dH�4[��A�\��b�kZ��	�$Du߁�h{��.� �_<*Ԍ���>V\�O/�L[k�4�ie���Wb�$/8$�v�I9�uc�&���go���=�|��jΠ+�Bisv����خ��|8���礗z��C��w۞��r{�n�a��ZF���a��驋�����(��<s������:y��q^R�o�T��֑��p����
##�{���$�k!�L���X�[�W�}à=^%�%�r�Ks�F�zE�J~�|e�ζ���.�8��Oc@�ˍ���6�p�@���}CӹfY�0������ې���g�^~�M�o�w[�}q��+�n�Yʋ;��Vj�{]r7��ؠ!�u�L�+bԎ0����E�-�g��g:]q��cn%���7ȥ�j�U.Yk��Oe�/�؂=�ܩ� },Q��'mu���=��q)w>M��i:P0w�?*���s!�8z�m^>�s�U��Kr����OUtt�)���J.�79���,Цs2����[��{p7��)�
�4V�73�ݱ��ŹZ�Iir�z��c��i��mVb:6��&�p-<�\I��aW٦o�G8uϰz(����᱈6ʍ�VV'IPDR"��t�yJ�h��-b�fu��V�B�-EADQV�"'f�iQAS�^���~\��b�jX��U+D=���PR�"���Z�X��H��1�eO�2��^^��T(��h�{e�x��E8ъ,�*���h��H��5�Q��5Ȋ�*�QVD�"�Z�mEX"�"*#r�W�T�R��4��/1��yh*���-��[j�R��mX�
������9h���V&�%U��ڢ[UUk)o�*c�T�'V��PV�j(�m�EQQ�*%�j4zt2_**�0̭jEDi�i���TV,�ETEb�(,b��[EA�
���B��/n^�+%E
�����6��T��J�[C��H���j񢣚��52�kTVЫR�Y>j��n�R+�
+F)5��V%k" �ͮ��D3
���K��j����|���[n��{f��i{�-)���@�O��t�B�r��i��)�P�-�W����r��/v�#9�k �
�ث��� ���}ll�]uN00��ļ���~�='��"����l��	��fϢ����?l�m�Y�b�����o�ө�>�=U���🙎�Sg��O��bgS�čjY�#kҪ�􎨂}~�֔�L��݄���({�H�n{�>�K�}��a��c�����^2�rmoxOm>@�T�Ҏ��r}B'й�![&�R����uBp�ؾP>y���s'�OU��d�ڭ�fн}�&����*�'n��%&�	g�
�A��	�`�
���IAOu������nj��
�N*~1�ϽR�{�H�~���&����8���vմ˩�ꇼ].�^���ڽw ���'-z3=�~�����D�o�"��O�j[��������VN���!x��dU}u�2�:�W
H���^���.U����8y�t!��Gy����%�n��b�D1�>��+&�n�??�&�AǚR7e�P͚���cS]���IH�
��	��ա4�k��B�kp����E�~����B��P����_�F�Z�x}�=�,�����槫Mn0�9⭽�hS����ʪvpY]F�Iu�e�x�J���9�B��撳�6��t8�� ���=��Խ�E.��R��ӆ�V�9c:l��Y�:J}������&��h�cq�� [/^=�X�k�@��$��ksVlS9ڨ���~��ވg��(>���0��wv�:+��ςS�M��/^�j�߹ml�ũ
&Ь󕊥x5�7dxv�����9�c(jٔ���F(���)�jM����]�,mϦ�b�.9j�Qf/�ٯ��#�վ��}�7�i�3��R�Gay#�Ɠ3	�rꤲ�
�B�!W��]��/�_4A����H�1U�+jB^-�LĽc�<�j�~�'\P�j��F.F'�-w�}�>�Pҵ{1���x�GD��SHa0j0�I�1*=�vq�Y�V�L|�G�T|�Kƺh��Y��$�ɠw~x|�@C7)��;�P4A\A%��s1�z���U%�|IV4e=U�q	���n��{T��~�j��WşD:�'��*��;ҠG��H���2<s2�i�<�Q��\BS�[���Wf�����FO��gK�1�1� �-�s����\�b�U\�p��?l�������������u(�{�0��Y�0��+W�#�C[�d�[�w9�;�ꌶ��1?9��q��*���żN����H�)M�i�)����0�Jӑsil��NV�HJ&���{���Z�0�Cn=���G�0�D�ҽ�"�{�%
 v�ש��*�M�[r {�ll5��:�;Y鮙�=����
糨��{�	};Fr���e�wpoJ�R��G�3i^\��^*��7��w7Y('�sb���3�������> {��	��r�`���|x��c��g�%���K�wj١�vd١����V�%����]��ف�����oE$�wCB�0�ީD>�G=J$�>j��Ag�:�>��Tx�xC< �3�L�y
��z�^VD$ƛީO�Ê�����������0�1q�=f�|h\xK(��z8E����e���q'���~��v1�D)��i�&�"�#�M^T���(���������Ƞ]p��s
���Tǜ�R3b�Sb'���QPm_����	�G^YIr���*1;(ql��2�a�B9R/`�Jt��U)����c�m���6�Hp����3{�~bJ��	`.�F5J[�d�;�y���g�IN������F\g]�a���ۻ��e����N��rB��Z����L��P����^�W�nO�s�wk�g��n튌=v{=����V�3��W�\0}�:~kD&��kHe����@k���T#^>��T(V�J��c�'<�=��x�znQ���4�==�b=E��#O��YB�� �ɹ?�5�#a:ۨx��Z��*���3�]� \���G��j{��Ɨ_X���&\�]���=C���ݾ>�ۧrC��3���W�]���N@������xdS�����݆6_x�y�E��=�.��c�f�2�F��m~����{���f��޵���R����৶������|z���g	Dor4sJ0�W���{��O++���N�X�L;'�fx���uW�ge�]�7�~qjZ��v�1�of�1co*0s�_{�)���KHq�}�*z3ʆ#���P�bdcsY39�1jF�f���3!��_V�m糅O�#ܑ��u����?[��_y]�/��̘!n��ZTp�ïz$�z�9zbc�v��BB�7��eq�,�	B�ZPq˼eʱ�~����$N_��z����{?%���,�і����Da��U�5\�-vT<7���������h9Ы�$��pTn�ǙR��J�_��2x���b�
����ܡ/ʢZ5����GyEz�;o��t�$���n��oЃ��E�qNX���i��`�V�K9�yTw���	�R��E/�m�-o/d�����ށar��-t@�Ƥ{����z)�σVzm?.�-��o��2NM5cV�.���ܦ���>_s�K	�)��82���$t)E��Ī<�='�p?��Ň�WqJV��!��d�6C�z��JO�ZUƧ'קH=W���S�P�����]�R��e��Zw�u{p�"��La��c��vq91�<c����lV�u�R�I����޺�[\W-k���ι���qGZ1���|���g�=��{7\�pŧ���$�E������vu�L��78C��Ul9�i�=��v
�x?�.C�.ց�ΛQ=�����D���i����ӼH7��矱h�j��U"��;	�Aؕʄ��~���n<S�U!.�H�2�v%����j�rK��ܺ*5�=�i&��A���en�]k�����y�x}���>���H�*����i�ׯY�M	��#%���+g�{��#�"4�MRp�S��>ͨ]}�`�dYz���%�8Ȯ*SAl�B3ד�s��tO݈�?_�o�c��Ti5_��"�<��"2F㊐\3�R�s3^Ǵ��4:ƹ4���dS+�
h��D����8\syq̯yP1���1�����p}g��__ng�;i9�:�sƘ�v��ӛ׍�]��gu�1�a;����,#�ki�	��,�Nj�w&\�lfE6�gE.��}1��x��� ��x�w�q�l!+����⾝RNp0�����_a����a�/=�jl��08/�Ve\�������+����@���>V?}i�����R�Lј�ol�-s��;7�: �d�̃~x�G7FV��2U�J��$�h��o���p�H�T�_=��m��HqՃ�z.C��;6:�a��4��~���䦷��ܤ����}B�0��h�N��d�d�;�o�{�ٽ��}�Ia@�=w߿Q����ǆ�qM@S��f*�z܎ҫ�;���r}β1`�zbL�j����z��ʈ�&ol	��W,
��"�(�����*ږ���Nfj��f������4z�AkR�Y#s�m2<��v
��~_F�L���G�*P3O>Zw��e�V�����^��9o�$6˭��	N6�v%[�/{&m�;j�C�A�Cރx����:پ�&f�L��r��N�J}*<����B���s����Rs�"[0��/�w���*����սy�Xd
2�gE�)���'�X��J}����$��Es�3�J�*к�{姯ۍ���v��z&<��]/���4G�:��~Ɠ
�*��;)��OD�u+T(��B҅��V�V�}{���3��s��F��(G�R	���s߇bypɗZ�a`�%��z'��C2��8k��o*�w�E���ŀ�r�醖�6���O�w�1:T�q�w���x�ɾ~Ⱥ�Vk�#W�r�\R�!��7+UD����	-W+1�z����:|~�j��ŵ��
��S��2)��������zj{��1�0��D�d��w�ti'�!d�{�Vs�5	�~{g�h�?:�H������گ"L,�d��C�f.�#q��F;J�1,.�D��{B9Kꦵ.,�Y��C���j&<����!)�j6�?w߽��� ��w/[�����B��FE,�h��T���-��f�C�:�w�)a�0��R�З�%�������:-miV�9��	�jz���f!�|8�Hu�3��F}�s#oH�,��Έ�n�Ʈ5֩��.!�Z�Ga�`(?@:�ŜQg�`c4�+��T�:��,���p��i]�F�ޓ��"e���ȉ��4(	��Ս�Z��"k6;�r߂^��2<%��
�ĝ%�u{c�5�j|;�5V	NLy0���'d�2'�X�
Qs����̘9�'J�u��7�
ѵ�7/Wu-���*�M��#�kD_�
b�w���Z�2��SS4z�:wgO1`��N'm8��+�m�y����Z�O�(EYQ#��H��&�w΄��l�S��w��o�J�T��%�i�3O�K��)U�c��'��4^�{X~��X�w1~��>U�K1JTl�J��J!�u��V�\<���G�@�אhs�a>�L��d\��m�WXCg���ϯST<��/;�bL��9���A��O���J;SK�X�g�B\�s�b%:aiT���J����N�0�*�=j}5�>@�g*MF�ں(*�^}S{�L������%�Z�Ib�p�/����3��x�l�,7�p��=���`s��K����ݼ¸H������1��i�n�J=�d�[�C�w��ߧ`$T��γ�g��Q��m��;Z�*�;)�G;�Lg����f����7��[���_�B��Џ9GMOMՐGay;�mC��%=��/�23p
��~�)�W��9���}x#��+�$�p-#�Zc���1��qq��U�t�
:��ծ�q �#���jr�1ŝ4;�RQ�4G�=|�g��6�WDjy�t��釚��vp��4���_��=����G.#T��*2���yo5���y~w�k���*K9�Vuw���8��+�;T��E�����gc>���6	X����7꒲�|-V�������qz��	����/����pr~|���T�P]у�B<>��e��:EG:�������
0�3c���S�F���a�'{\\gN�\k���rą��*�G%0�m��~��Q�\��������n�I���»�ݽ[2�6 �H�;�e�њ��1Y8����(?���'�*�U[�=]
�/��b�0���ę���(bI�e��h{҈�-�"���SSʒ��°0!F>��|}��T}�óR6���:��6��&V�%���/��L:UsMZ��(��><j�>�t�Ň4���<��+��̻=-�pl��� W��$H��[OgR�s�튋��=�LL�[pX���Q,b�����\�[M<B�୦ٮ2�����j붚�i>̐�I��=����ϕ�ۍ�`g8�z�sd�EJf�^w4r�eG|�}�2"$*K1P�;�����y�n�q�
��X��F�遚��5 �xK�EM@Z�d�`��m�'����O��ћ�������9�zI��
V�e|��7.6��(���������ˬ[v���:)����y�~����Nʡ���-�RVjO����<��8��r�P��R�C���Ϗ�)~�����=����_���
Eq��Ǫ._�v=Y@;�0�AM>���M-e�F����7+�&�/ιu��
 rQn�m>��H%���P�5"r���=R��^�}��m����.�o��݅B� ǣ�K!�f��O����?Gݮ/����>��$� �k��G��+��5�!W�twV��u%nm1*|���K�b�M]�L�Y�M	�$d�� ����P�đИ%Q��<���ze ��KD=��e���e?�i;�⬰�}���6=�N�����* ��Uz�����-A_0�6�~��`U�'-���V0�O@t�m�Χ�����V�T�p�)�ye\�D��3tpTTd_F���.���<fP���c۫Y}og5��@��_h:zp��3J$dsӾ׼�>���n ���}>�Z㵞��A����Z��	���N��:.�Q��!�Tt%��v�VNY��EΚ��[B��_�祥�u |0Mo�� {�{�m�2�fE����xLv���g���|H��C�ߟ
c��=���b����,' �"����mG�&��7�9ƅ8�0�yJZ�@:���#�|��	�1}2
�+2�;MXF���$�p�L���ϐ��L6���g����	���O֔�����!�ȁ����PB}��@馸�P�D�Ƣ�(���B�����Q~��AR9��|�:��D샰'l��F�>��ԟ�D�?<}�Y�1"�Ǻ�tnG�U�y��x�rt#s[��wq�7���9�%�������Ȥ���ꎴ�I��<X90\)��ql�1+}'�݈�/sB��#k���5�F~���q(�ـ�\��A�ə�˼\ʝ=b3gr��E�t!�>��ؔ�����^ځ9�u�Bּ�#qY}_r0�|�ް�O�߁�xs��*O��x��Cj���">������J|���/^�^P���^���♭�{
��8d�B�l��q���f��y|�@�7#A�4���/a�u`1�n�9��!Y�s��j�L|��H�y�ޏW����z�^�_���<�������������,���X6M�^���\7�n2�X�ٰ2����}��
�<�;������7[�6��=���ן�4�K��]���n� )�.+*�K�iųnP1o�i8�t�F��@�!���'��Ԥ����a�aΣ���N���x�qN�����N��V���;oɣ@�[�>�n��6,(hxPt��:��>� z/hɣ�;#7Ҩ�˚��7�T/4���z�\Ɲe�Y�ٓ�]�.���!T��B�Φ��Ñ�ua�<p�+r��ɠ^_XpK��ݾ������1��Ou�j�A|��;����f\'m�i,oqu�FVf�ӻ��",E�;[��nZ�����0����}}����xpדū��^�F��KHfF��]�wz�Z
՚�CJyKw6l�e	Vصa�:�U@w��X�W۵���r��C��l�M�ƶ����G̲:-�Ozb9a�so�g`��[�q������/-����ѬJ�K����.�=��V��@�S�kٕ�D�/G���|��t������wԶ-��}U|M[��o���![նSY͟<���Y�M>8������͎�-�����	;+��ġ�R�Z�u�R��4�/h4Efӷ�Z�e;��S�$*�Yrb����J���S���Z.�:v<{�"���3q��l���a-���=f�۫��y`aN�M\w�sx[hQ���)񧌹)4Xc����������3�zk��!�0��oM'(�5���y}ǃ��f�/u��eś4ؙ��k�sUh���YkPrw�P��J�HmEj�.��[H��4o��V�n���3�z7{N����x���Ue�Z"Dӡ��G�I���C�m�H�.y+
�N��C �T�msC+SJ��@���ݚW^�F_m�]��e�8�*`��SY�N��N��M�V�B���`���|��^��ʻK�9'x����c������*�e�\���LoV�#49��v�Խ��x�r%�ӱ��w`�D5b�o�dT�����x�jŸ{e�%�b�Ǻ11h��1���cÔ��41y5Iǋ��ہM^i������|,�X��Q��強�����Pv';kvd���v��{s2�C^�{�����9y��;w�oz�,�Hg}x���#D86̓]u���
yNZ}�:�
��/sV� z�|J�R�}�肶a�lR���=�ַ�D�b�m�oXǭ5�zz�5�7Q[bG:\���OІ��TYS]���E$/'m�]��h4xk�o���}�|���r�p�9��u�&���wjA%�q#4��m"�j��o�yc';�N�{vU��{��:�N|X�������r�Eݽq������3*�ou�X�TAEkT�/WԬ%j�e3c+(��30������*�T��42/.3LٕEBڳ5����*�`3y˃���f��('��#"�̬D�bq�T2d�""�\�M���͌��cy�A"�"���°�Z�aZ�m
��XJ�-����h*we�J��3
�R�B�\�"��S�""�T^��3īDDD�Db-a�-�#TQJ�Y
��TQ��ȥ^P�N��JΒ�
��[�e��V<R�Fӷ��E����C�X�(�6�m�^sh��R[m�j�5�}Z�AC�
µbq�Ե�QQTR֒�j(��[VWj(����b%B�����\�i)J,Q�aP�TS��{�����QN�zj �69�"������f�jPꄺш��Qm�E�ז���թx�V"3QE�Pe�V,�Z�Z,��j!ն�U̶�ӏI�C��-m�P(fT*w�ǃ���b^��v���b��t��]�	(a�.߶m��qә'�_f���sO��RSvv�L�uͨ�JB�G��98��rY��a}�Aa$"���P��7� ���ا����!��/�d^�<�=�R����`za�5i��}�Ǜ�hu��nT:W%圮;Lzg���PQ\�O�*C=�CT��T{=F\Y�<¼WO7�g�U[�X��v2���8���*)��	�%w|g�O����^���-�ꊭ�O������ʀ7��s���fi�'����!�=�+�;�WL�yD-k�*(�	���d�<CG���i��j���U�F:���UM�Bx�4�v{
�L�r��!x}�(@��}+�{����wACetKsjF���L渲b����p�C�|'��C��āe�Xa�O�H�����=����/=/4�������wi�������Uz�K9�0�/=;��S����%�nx��%�^Z�����dK[�8Nd�;�B������F���pg�q�cv��g!�V����!���/��L$Y�-p<�P���E���w]�6;a�*pm�Nm^^i��k�����+�9�77DC�h��P��{Ɓ��!DKr;�}�7��y�@%�����w�A$ a���n�����\���6�d<����<��K�/l	jq�l�X1�
�:��(6�3yif{���U�J�
1ۗ����U-�Q�g
�O]�z)�:��}�	�;k�]�2�\��u�|�}��~kG�'~�~�������)$:;�������z��I�G�	��3��D��H��B�ne$_&����|�J1�K���f�L�e�'ʭ22�B�{Z@���0���9���og�@7yb�cʈR�I����f���	߷����!&�d�,�B:$����p%Tȹ��m����aEFd�����<����Bm���}P���/���:3�!M���W�)i�MԳݟ��X�vO�(lp�
�f�m�ˎR�%͜�Z���fc�]��	�	��@o'��^C��4����)v��b������	Ȉ�z��U�:���s��~'B�@��S���K���m~��,dv�otޕ�!_LKj෻����BF�{��]�$w={T[sP+�P��%=C�WDC;�{��E��FWO�"��B��nu��	�d*Ӊ^>��'2��v�@'x���K�A��6��^��ϔ��m:�<(,:*^[�F��P��~��˖�!eyڧ�j���\���j����Z�:�u���`�A�]�~dq�3����j0Y�u������}��*鸁��.$�E�g�lm۞ۼ�$�ś=����.��u�a�"�> �F��j��]��7/���N$��|.��1�/EZ�`�{o�Uq����%�{�<���ՂĻ�9�.wns�z����}[���cD$0��M����g��3ئv��]&)H3Z��CA�w����I�S�D|q`(Y$@�B � )$�,$:9ϯ�|��ϧ����@4�.?��Ɉ'`!�@���vg�7��9FNq5��Hgz	C%���s����ov��~�[��Ԧ�"/f
�'��}_�L_yOՔ��="ن�����3\6��@����S�=�=~��h,��Wp�򔸒�P*�A�q�EF`wn�1��V�>�l^� ��k�*���B��`Yu<�Sܩ-tD��K`Q���μ*Mm��Pv�+�r�ˠ&��vbm�Ѻf�V�8~~����O� ��r"*�[�sy��ra�o�;�ù�H�u�:�&���`{��`u޹��50Y�q'�,qʦ�++Z���d�T9ج�ܩ�C�4ؔ���}r1/JF�����M{i��8�*�i�z��B�O�8}�g��F��SFG�m��G�<_W��I��T���l�uI`�0e�	�g�_%�Ц�r��:��<���t�Z~8Q���ɦ��nL����1��M>r�s��#z7ud��l/2'�Y�{[�X���A��3��@M��E'�Ĩ��m�*�w��ܥf9�>�_@����t7��9�m��2�3�Bd:Y�9@����R��_H2i�l��?=[a�I@v�6P�Az/ ��]�njmm�qq��j��ӒX���q�Y��K!��}���:�T�҄�%�J�'�9�n�}�����|:�u�D�>�	"0, �dD`
<��ϟ/�O�O=w�G���1i��yv�/��57(��G�t7Di�~��'�@�a�"�a�r�4E+�"���OB@y.L��|�H��0e���hN���1>���]�5ÿ=<����Mur.����F�h���`�) �'�B�j�����Ι�8�EfϢ�7����f����n�<�dL>�����
�X�w���b����fn�5rj�/߲���o����3h`���0�X����C\X�Ƽ�<I'$��2��Ƅ���2>����(U.�6���f��e��=���w��1�x���a�3œ�0U|"|���V�x9�0j[��s6uf���KU!f��v}�S��}]���5���SW�Ej�J[�j?h���*��v�WI�b��
�׽F ���ّ(ޮ�C~�'�VN��9���v�i�n��#=��^����0���Y�1B���fQ������!�FD�c*���Oo1��|m�$���(>��v��>r)+��`^Tu��$P����!��}�N�w�����en� �$�en&d����PX�Z��کZ��VZ�emry�����iX,+kn=�l4�-^��aU�z�d��[p����X1��
�Υ�k֖��3��+]��_s{�N���v�P�=J]�f���*��0�]$5�	���92��?�U}���E�P�
@�@��Ydd��~��_:�}]�o�~��TV�G:ïSH�����>'d�~eȟ�ȼ���tJ�w��Ns�븤ZY%˞��g�vyvо�U����{PD�B/����o��W�A�zu�Ŏs��暶�`W��Ղ��~� ��Q|�T�%gl^�Z���9mF�c�a�P��T/]lZˏk��Ҝ��`���J�^�ݡ��&�v:p��L5%s�y)�J��6�����g5����Y�} �	��C�.��P��Ax�qPg5�Fk\7������Z34N���+��5��ɩ(����A�l��%c͘-�0qzu�4�{5�(]�R���S� �4&	�H���V,Q�Zq���1�x"=��8'�8APLX
��ia�0��_��ƅE�uV��n��R��z7�I�~������D�'X��/���BֹZ����菆�q���yP��k���I���g�e�}y�XҺU�{;�89?l��Z�Na�\�pV�����``E�tN�Wm�;�;wj[n�*`���� S]:i�|Lf��c޸�3�ԙ|'�S�PA���y��*1��c���:�F��D�J3���o;5	�4�ػ;�P�nx>h�ߩfN���NW��j,=}����(J�N�Umq�0^�\������:m�����:ے�=�z����O��:$�
ߨ����Ǒ��31�GPl������x|���`�R�P �P��G�)���*NV��]�M���YpC�����f��3��|�@q������g;�Bz�ޗ]:��9��|�؅�ߝ�so�p1�7rD��x�5�Caj�UUO��t�9L<:���Hc\�@�1�0�<RV�����L�R��c^fL�9Ovc���In{����0�0w�0"��d/���D��9���l�=�ބ���p�[��T�wq�c8�*Z�3-��H��^�!6�*�V+� $UcʈS�JҲ��VP�3x�9����\e�^lE!��q��{��g������5������w�.�<��"�%�����>�}U���K�'�Vp���~�����#;�Y{������(�wXA��4e��]9{Q1�I�jS�Ԥ�.`0��:���#��|��{+����4���)��U)��C畉��B�������������lO�`�pM�̌��N��|T��E�a��ؼ6�۸2�2�����y�Q}>��y�z�ؗ�Q�'��}�QkMƑ�]&8G�.���#D@��/2�Ԣ��U��(������uA���vn+!���E����l]�,��T!�C�*U�9.NX+��ynn>P'�
ji��WVɵ�-c�SQ���1�4�g#�yP��{)[�Y�f�Ǘ#;�����J�|�b ���q,	 �(C�����������7�{�OB	S��?s��%�c��'��ǒVr|^��+��`:"ݟky����݅�n��F�*d��=,Ѡ=�Ԛ�(7y�&�y�Gk��P�yuf������*�;|��WC	���_�c͚�{���_��Zs�j���\�S[�*)�ݪ���%B�A�,+�4��Q�T1S]�9�?B׻&}��VzF�����a]m�gj�t�?��&<	�� �����L-��t�|f�:�=������4jO�OM<Q�<7xfL��rrF4^�J`!�<H��(P<� ���	�b��wa�l�V�(]SKtvp1(3(��nۑ �O�������a�)��`+�Pa�5���>���g�ݍ�qWD���G�s.f�sv��s���",��p�uW*K](��tT����L�,|A�s�{�lֳ ~�Z�L�9_uU���4��q�O	Bf/�Ҳ��9HC�T���uD���r��i��'���!?H�2E���M�H���_ö�ǅ�z�F���N+����k"�[�DƔ������{my10�敏؎�n��ld��wS�������Q�{�bL��$=��j%�v��</p��CL"~�k���)�f�N�8��5�`r}����9Y쎱S�����w}�URt��|>d ?xy�{�����=�Ka�Mp�����<4�@��J͇p3>��H�8�cR=\�b���SO�����͌������'i{9�{��m�3x��
��z͇�T=����ܓ�28�G	�B�@s�ѓ�3x�2�7{����5�L�I8�O�Q�f�;*�kP&�%��e׃<c�gSW�2{"��wۊ����2n'���a�o*�v����5����)>�%@ɇX�htʺ�z�y�1�&���cS�nj���\����(h�|��HtoS��X�o�Z81���6��	99
�����B���筑�/^����~��=��[X�}F�4+��&K-���w���18�:��κH���^RI�K #�#D5�e���j$ΝW�B�1R�e��]�=�|f�4h���Z����g�*�����F���	� 	Š�3��\nƔ��4;��4*��`��m�[�n��j�m:c���3��io���q4"@����H����p}d־зմc��ZK^��u�
68��;�n�^&��%����P�/^�R����2bI^�}�oe��=�S��8,��&�[[4�w:��ܕ��|���]d��l`t�^����7S�g��gr)D����ɤ��/��S2=8c�kW+��;V�δp<O=�5�v��1X�Q���P:�,��-��av�N���Y'!���9￼$�fHEdX@A�~ā��;Ki�+��	��I¤����~,�]ɆkR�M@�SBz�K':�=Zz��0/o6Z�����V��<|o'��j�q��?=�,��[���^�-� R+rY�dk���g2�N!Oe�T;�y�D���{�_�� ���1�.��U^܄�׊�J��^-�C�FI��̿od��P�}�t�q��l�g��_R��q$�J��[E�R!߼��2��xWR������CW�]�
r���~'(V�5�)�b��y�}@ÓJ=��)T��]<-5b��2yu6�"�Q%��z.{����v���7�U}�*�/!�1g��3��Ք�j�;b�:�v���d{ ���G�����sP��\��Rm�$k�,B��R����ա�� �dM[�{���.���'��/-�|z�a�Ȱ݆7r��|be'AtS-~ (�B�v3oI����/1؟k�ۀ�M�*O�V>�0�@�3e�?vo���C#_�H�X�R�:�0
̅;�|��3�^a�}�P��ȓ�q�������v5?
��W��G�����ǐ�W��99_O�N���$����\ciĸlZ�e�w���S�Ү�D��������<���'7o���q�7����cH�����*�?�Vx��m{ �g`�S�V�F��B�n:��=����K�[LW:4>|���	"$�D R}z��ׯ<���}eլvG��K-�x�{
������!�!+�4�0蟛]��O�b�$�i޺{x�)_fv�jrGs�������j�DϹ@��M��^y�\i�"���n�귖���S��ɤ��qPģ��x,�h�USkW�Ŵ,���u�x7��֮�[wO���^���r�c���j�i��T[���pK�S��p��|r0��7�n���#MW^�^�	~�GЎ(
�"!�5��ZD�
�n9���~,�>�`c5����H�|Xy�G������'D9�/��	�;�m��I8b���9�x�<]�-��۽ʬ��и6$�A�L��h�]	jz"$��G'�L-n�E�nFZ@����^���KwA}�mOB4.�gd
��/C��A�9K�!��7N���/�
`}l.�*�Q��wC�睙��D����z,�캣g��f$S�Ϩy�
�o�H�Ǖ��%�R�c����kݗ�N�L\�#�ju�̚�j�*��q�d��];8��J͋|WQ�@�y���O�����z�^�_��_O�}_�(�T�<.�]��nl�Z0���X�]u�� \r|����]KJ��+¬��1{��7�X<���p3�5��yP�c�C�9R]�DB�N��Wۚ��h���b������S T���t�����4�vU��i�q%K������G�-F%ϵ�&a����酋���ɭ��V�T���=Z�Ya���7)�A\��`ޚэ��)�_~�y�����c��VFq�ٌL��`C��W��d�R���ì��l����5&����Sb�^Kե88V(���Zðcio�x�Q�H��ձ�s�Ҵui�Ć�}t�����c���]���~��h��>�r�Z�n�l,�5h�K<H3�V��Z��kI� �����:���S�`ǝ�Ξ#|�t{��|�On�Ww�L�}�Ol9�9j�<��zM�~�F��U��)�2n���Νv�x���i���0
*ԗ�j�Rԭ�0κ�����;l��D�������]ճUi�$8�-��j;XK�#V�y�9ϡ�X��2	�uNc#����^�,�.(w���/&a/=�
�{+wl�<��I�ɣg<�ý��Or���u*9� ��j��Lȍx��9;sb9|����Z<���_�����[��#��e;Y*�{O��1�b�>K����,t=ytP��'�s��䣗��yÞ���fV�ɛ6��5t�U˪	G�;���M��ą\��ZX�9�i�$k�����փ��&Q4ث ��Γ��4����~Mg����]W��!�#�ɔ/�!��� h�ŝ��y���f��}s���ڵL�|�������|>�c5	��Z�mCI����ں�ͺQf]�~j�;�������2jL��V����O��k$���V�R��[�zo������ҸǢ��hɴV)���K޾�.�R4���R׮t�C�5f�V��%U�i�yNs(ؾK�L��Ų�������sN�=O�]�q)���{E44Cmor뿥��XU-4�SA�\N�F��工sp����%�cI��!���h.r_���OJ�֍�h�ַ��ۡ�sG�]%��i�LR�x�@M��X�V5�#��P�����.� ��D�]@(�.l�wO(�(�U�st�}:�͈6��8�j�r�q��eěŰ$<�Z�n��~��@�]��ޒ\m
�y�X�:7�
�.9M�g�+��P�r��dE^�3o\��p�u.dp�X�DV����\Lum:�	g�B��^�a�]$d֫�pg�'N.��78#o�^�9vv����U��V4-��=X�hl5Ǽ����-^�՞��û�����i�3l��X�:S0������Tl���B�l��n���;�r!v_��<V��XCX���N�j4��������:[��OHT�>�H��\t�*��e
e55?VJ�qp���]��8A�O�O"��I�`(��MLr�Q��#բ��F0<����+Xĵ��+�Z�-Dr�[l-ec�2Q��5��*r����*,F������u:ō���,[eL�g��*��%W��c�P^�eN�0E�E�kS�PQB��3*L�^�D�i(���q�x�W%��8�X��L��1���j��A]�����ɩEu6�J��8���٩�dQ��DrX�� ��[g`=S+":�Z,X�$ج-P��D3m�QEzj��������oWZqڙ��Mh�ʗ�
̔E��-J��ZǶ�QV
t�2����,L�	*n8DQT��h�q�r��i��Ԣ�t�i�T���/�Qu	Zr�b���;d�q(�¢�2�F�R�EW�ìZ�UZ���yF�U��(���p,a�ms
��)ąQ�`�J��#mg�U�&�T������9j�=��E�H^�J�,{,�t5�פ�|ۻ��,DR5�M�
d� 
��頲�����0�.�o������P=礏B��)���u�Tѽ�0X��6ih k@�ܪD�a{�Nh�Y�Kz�wN�a`����B��kP��� �����#��"��1�" F$�">*w.��إb�g�qY.	�A���=�6
���vrú!2$̱��m�����[Q3�.�2�MF�8�l�E����}H�L����i����W�T���_�(i�5�x�G�7���NEfD�-�Z�Z_��x��^[�Ȍ�wW��J��(���dc��B�<��{coxR�������JO`:�.���m�����@��'f_s�%�^���ub舞��k���e($j���Iz���{�'�t�_~�~�+'�B��BC�S ��rͿ�vO{:�k�DY�=��Ǝ�ku%�87y�b�2�֩v��c��Ry-o9G�T��_�����fY~>�cޫk�S��<�KFR��H�U�;�,3V9��љ��ʂW��p�vd#��}��Ň���~7�����w�w�>�gѰ{�Z#�ݭɕG��p�h<�*g�,#�1�Fi?����fr��W�@c�9�ڪ[�GA���q��[s�k�U�š�̂���\z���4^�E�����d(���0e�x��|�����G��7b��!�����m`P���RXT�ol՛�q��+��%�eQ�e�0��t����ii�+������[��h[���Y6$N�;4Rܲ��81����rLLh��1�z/�}R�B��Sf�a��],`��q�������O~�}��`��E`��#��F�)<��]��y��^�!3nq4��n,���0JSi����T�<�-2��
�Po�l"r��T���I�g�V���/�����&�C"��s��x��4�ujB�S_K��i[mɱͧ]W{��g�<�Y��>׉�\M�O��3����4�'�*L��{%z߲N�0���GE���uAmJBf�G9����2LE�n����T¹n��"Gx��#�N�vC���Ig:n:��:��"cwV��/���j�e�foNd�Įԅ둔":�7N0�q�S�6@N��J��o*b���^�Y��E5���v��u�����R�"���)&�����?f=�q��a�[٭/
�z_��pk�,��S�d�簔ZrWH��,�a�@���:�����q"J��,��v�z���a�h�gN���J1�0�׼U�b*,:�/��a'�v��m\�i=�[}/��u����><��
bT[U+��6�������8�jt�N��m��X=�Ļ�U�"W^^��>��+��s��e !�yNU��<���Y�&\&���ϻ�}2�K�L�)�_W���ɋ�d+م��
������N4Wwn�J4�.h]R����.5�ޮ�����Y�X��G�$����R�g:�F�Һ��ܑ�<����q�!pCRUc��Nhl�u�Y]��=3]�oo��|8}��,��� ���dX�IϞ�����߿4pw￑��L����d%�BZ�E
8�4s����^,)�s�Za����a��{{*�����t
��]z7���&A��`�:��Š��Fߢ̵�&�|����"IT��{�dZ�C[�ʝN4�"ج��:���s/A��ă��H��V�F@q�}�'��홑	�z�۫�n=!���5����9�:���3�s�yO��L5�B';
��!c��w�Y�o��T��ѱz�$:bjrg�lu}��Y�윭8�I�R.�ާ�<���yO�w�Odd���OX0���	�x!����j������Ջ���`�2qH~1�a����5~��]Df���O }Α���g�E��?;}⃳%J����͊���;T�C��Pۯ{3<Z��������R���H��i�z~?Q��)T�gY���E�Y�������Ϣ�^��ʶ�Ȇ��qM�<�m��XE�s�uB/��l�󃩓4&sr�����{]#봛�;1{5�r�z�[�kl{r��Y�]����������eڷ�y� ��5���ff":�U8l���H矕D�'�.)����͓��4`I2��Z�!�R�ԁ����@�X��s�8*��:wtN� +vm��5v��[Zд:��h���78�ա�ք�Ү�6��N��F*�4��q��?@  @A�@P�
"I\��>���H*G�!�~��es��B��¹7�>�J|��+�<��yy#hr�2��K7L{���!sk�c&�ڕ��>���s�|z�@�ll'� ��>$�OaD�I�qE��n~熓�$[�U�=.�������R@u1�b�!}?�=)��i�sσ��m	��yd�a�jS�m;�ͦ��Twz�%[@��IJ�༴"\WD�cn^-G��/Nߊ;�,��(���߹EM��w�d[~����"^�?RZhyj*C	���`�a��/�G��qu�y�K�k�}�������ؾ��C�>�G*y��"^����{~
�x�c��)��>d�z���UQ��gͭ㬱ׯg�ӽ��nK�^��k���,;�f9_�D��N? ���K��;o��i���2�#��i������g�՚��5�=	b|���hLC��߶�xŔ7 ��Dꠟ�D���*�ZD��Վt��ta[�
�Eζ�}\���w.���*O��[.��;�����_b�|�/+�m��F�ۙ�A�>�II�Jgڶ0k��7�VbT��v������2�^!��!�*�f8d��o���SR��q�&S$À!�,G1��g�s�/�5�l�^Ήjq7��,+��aa��7��BR����I�ުΌ�tVi"1�: v9[b��ǿ��ؔ�>̄PP�����й��N�._��`�}�d`���29�4'���� 	m�6Aa"
����I9��*�zV#dx��\D�c?��5���fM�\\#��^��"q�� �?]"���1n���}ύy������wJ>�ġƤ
����L�=�C2��gk����>��CTB�ʒ�野۱2��YB,c>u局4����R�6���j
m�o)d�~�4�l���%ybπ��ew�{;��!׋ۜ U�bB�hy��#s
�3�۝�ǗQ°Uto
s�z�ύ�<�E�@��N����#}r�B�Y��+�A�����&Ep�>�fq/���A*��~&i���Ok��.+i��&"��c�tО�b���=/«�V�#�C���,:�E>y�Q~k�������5��Q�+����"!�95ܩn<�(�Õբm��j{^�R74ܷ����*�;'&a��P�z�������`h�']��-�ӷ�΄L�.����L�g�2vw=^6}�̟ ��ᵧ:��5��	�F����<��'���~����[oU.(��Q���<������ߙ9d��#دt�k���ap�h��U���W��$l�N�k�fL;f�IPGO6ܕgj�Ʈ�H�ښ܁v���hR��`�gk\C���|&K�K�s����~}�r{���X�,�) REO�{�����T�~'��D�࿇��2���,����U�w%E�{���+��D�ө�k�JNm9����Ð���>��/�x�Ҋ�8'�_�fo����]��k�O�kF5��T���Y�ݷ�9�+=�`=ط��2���a�'�1���!F�1�*'��l�����:q���PdR5����z��'�h��x�%0��{%hypA���&�&:���5l�M� �8rc�6=�Z�/��z��G��4�q�a��	�h
��7�����tdkݽi���wWA��]�x�Õc����
.�e	�ޒ�y��H˰Ɛ�Ƞ�j]9ظ���.�Ʈ�0k����W^�{�T>#L10�,qj>뫉�:����vzKSM�'U�i���1��!K��m�ٱ�p��@Ť�Ӫ�Zf�����֢E>�8�MG_8u���;,�7��;��'o�v�<<y��Q��ei��k��E�u�³r�FP��D�8���<�����9���C��m����|�C")���(�}�uf�����#�#��$�q�D`���~5�zT���� ܉���g-&�S\�r�8�V����b��D�a�@V�%������g�A��.:.���'QX�l�ME��V��0��H)���j���S�����.v�wN�!=sU����s/_u�Y�^n�N�6e�7;n0��x|��x3a�f��~J��ρS�$lt��):�=�ܗH���l5���Ǡǲ�>0�(6n깤�Tҏm��6�
}�!�����}�Qk "�è����^�X��*�My�Il&����l%�Т�#P��{�迋�	�"K5�e�����u\nRu�2�@�g�O7<���V��5%�_��j�:���IĔ��%����T�k�{t+�c�'���[�r̴��6��o��Nw[t�ok\�����'_��58�$F8����D?���^�q��Η�zb����ws\������{H��j�͟��s\hG�	�+����KI���ό��WY��?=�پ��^F�Ra���\>��f7T,�y�1��xg��P� k��DPi"����F<p�S|tt��V�+YH~.k#ؤv������-މ�a� ͗b��:9��Zލ5D]�Վ���Z� }��p������'m{Wս鴴�ޏ�A��uvB�~��%i��L��xu ��8�w�
���o�&��AF�'���fd�5n�q@�L���N]l�|��&���"k��;6�;/yMg�r�yM ��d��j�e�7o�	�i�.P�e�� �>ǧp<�x�ݺ{5=(��5�j�m�:`����j��k޴�h�!i�ӽ��޻����0]�u���K�k�w2��lc�XؑP�@�D����}R{���W�Q����J�:G��3ȅdI�]9%=/X�ڮ�t�2�ܺެr\T�yb��Ş�nn>��9O��.�P��T}k��}Jy��UԢ�Vѓ�NO�2�e����Ϥ�۟j���.U[�ko�<�[a���41��)�_Q�9 �Z�}[c}	���.�\/a8�)}�����+���e�)��|����u���׵H��u��s�>�K��Geʞ���i�E�g�Q�2��pů��צ[[����{H�*wr16ʜ�Z��R��+)Ԯ<�����3�V*��_W�#��z7}Ν/Bm?�'˕J�ez��Ᲊ�ה:�/�֡f��D`So�͢��#����3��8>�y�G���Y��A�l��'�95N~��킴-w�Y�^�!���l�+�s��qϬ�%X9QB��1��Y7]�͞�z��B�Ra��S�7����a�a��(������àTv���Ҟ�u=\���k����Tx�f�0*T8��즧�q��_���%�Z��+�dc���wBAg!���*���1o^�gC���Mu��?�΁��1�~���O�Qh�It�\S��/OkH�e�I��Nb�-�&Y�^��U�t�2���S���pz<y|��ˎ�92>�
jӾ�2G�ү)���5�$�l;݌����0����,���?���"" �<���3�������Ȱf�<��3A����:z�z��걸�dPYʗ�7���;�~ѹC��XW�<�m�{�qG��B�C�E�Zs��>�W�D����ܬI��ш�f��$�3>o/�,7Y	i�|X(LC�B)�0�z9Cp��|g�G�EA��oӂN��Nn�<���N]q�^��Tf���������������vϞq��8�ư�2-�/����EW�{Ϋ��7ij}��x��-��z(����h'p�B�P6�/#x���ӷ�D�/��>�ڦ�ܿG2�)�6/"�')ud ��wPGB��g�v��w�u�b}�v�x�>RX�+[Fb���.SCh�"SMzԄ�E]
ǰ�EPǕ�����j5������@x���/㚋��l�O�(�;O�;_��}��<z�M2�kۗ�
g�-K#n���j�ֶ�n
i�=ʈR-bO�|�b&����CG�l�B:;�X���ѱ������̈����լ0"�O���y���VT��B��r��e�
�x����񱓨����ݔ
�2/P��L ���!�`9W�F>�0������L���� KE�7<9��h�^>p𞳨f��)n�\�����q��
l��D�[� _k;HI{�Ie��W����a�l�n,Pp81�}u,M�.��	3���_U%>�n-�Q�i�D�L,y.�M�B��?,���T�gc�P��Wy�l��8�!w�
�2��5�,Qc��*�!�GQ�Ү/�s���G7RR���T!�!<
��R��m)����w�'�����.���}ت��`���*�=�Q�'�@�[����W$�ϳ�?M��S��_&�e_!�W���eL�ю|h絺��!��qǞÅ�7]��Y�<�Ԋ���יS�Jh�p	ΐ�h0�8/��fz|&cǛ4+w�|v���d��	�F^j����ͧZ����c�W��r���>��� pG�G���5H�c�R�F�S�{�W�����s�L*�k�1�l�Y��$�zGa�l��$0���3�P��������q,͙�%�K�(��n3�7����3�1�?.s�y)���>Ĉ��\S\Ǯé�~}���/�?C#s�n�6�^ݠ��vݻ<�d��PB�ʹ|=5P�R�����6�M|�3�����х(7�z&2"i���c��qv��ޒyt��HB���pHO&�=NO'S��u:�N�S��}�}F3���?~����,V���n��Б�=q�=2'Jo=�W��<�G�YR��K���4c�bm��s���8���tg�A�0H���qJ���2��@�i�r���>�40vR�V%��41��VTq��*�oo,��RdC�#mk���#h����_c�͔ՙ,�Ť��;��.����eGcc�[��QMH�o<���rV /�ve������|}�*q�B4�l�<-�Ǹ��]s�����R����D�>�oL�L��ȋ��6s՝P�d�r� �yQ1�38U�D�x+����;�3]�6��d�1�Ǽ�,���� -d�n�{0kdl��n,�Cb�ݤ%�6.�,T�%�-��| ����]�޾x���>3����g�a����3�:3glˢ��7F�e�-Y�k8��\��4�b�3�3���\��I|�xz�7�j�o�;'?>��+f�cսvX�$vr[�.Y�6�����S�J�^e6��q�f�[�u=@�S4�mڠ՚�;Zq"��Y��7%Fa�S;/2�l
U/+Y��ʗҨ��6����-����S��nü6j�N�&G\�wxn���w[6��������y	R�D�wW[(d9�i����S�;en��\C��㹑���Yx*���n��lp����*ҷ5<,�bg`�-y|�t�ypy�oyQ��j�u�g�ǎ�$$�a�ŷ��ǐ��t��5���/�=�̺��#�ް�\�� ��Ù��n�t�@	��N���ܗ�1��+�E�cW���l(: 3p���Y���ZJy����i��.� ���;�;�K�Ƕ����"�Dc��� 5j�	w��ι����nC�50N�U���$��T�}�F�:딉�nx)�6t ��ԍ��=5��r�Ƨ�;=��]��yxw��B`F��Z���cȪX��o�ʋ��vr72�v]�1*�	�+��驽Q�T�s�	%]u�x���hݹ�ny��R�{��yn ��9�v�;�ڶ��F̵��K(h�y�]��G�!����x��w�%�bȭհ��ku[h�MHl��y���E�H�a�#5���*���{K�>57�=�ݓ�*]5@gF�{��R���݂���TlisS�Z�������ǴeW���W����nb�M���8���U����ڛ�`�t��J{�9f�֖�ο:帙�x���a�a��:-$r��,׹�>��4f)�P��v\�#���s�tn㛛��N��3��y�tK��}�B�#l��2Cs���%��Wn��8�$���x�ޣtĀ[s0�<Z�ri��y(<��z�B�s=[��d
��}O���u|����=�q��X6O	�� �Z�D����)>g=b�]Gq���뮲�����{wjM�5�����;�c����(�9!�1����3�Db��Ro��7��
��`��TV�t�x�XEKV�X�trQ���\�
�C�����)�i���8Q�*��Ʌ��8�:�j)z�KM���������/0q�Ȉ�q�P�B�eQE!�VdPQE"�h��X��U��,�v�^ "���u�FE���8tY�	39�Kn�j]`�Ajf-s9�7M�QeKl*TD��kAA�΋8�Y:J�z�E�==n8���QQ�D�8��t�J�Q���P�YP��!�&I{h(q
5��[MB�8��-�������Q�MK�E"�9�ZTiE^|��DµR�Q�ϧ�����[����Q�_��6�cDmk%�4�y�d�m5��fMnM����8EX��o6��I�j�Q��-�����U`��#XU@��R�)U�t*6��k�v�^R�?Af AB!�G��/*h�̰n6�Ck���V�Ԍ�Fb��#�X����v��&��5a��:<�Ź��{���A��2Ց�5����OO4�t����=�����=H�񶸦��U����
��_ynl��_4�:�g�ؔ���ew���jx�>�1T#�G�D�+q"�/6��煯nw�z/L0��"�FFǿA!���4ɷ�̶�K(��ʬ���E>��+7 ���9bc�#�rw��s�F+&��ˡ[c.�@�/
���N���)�{No��՘a�Sy�������;�w5�O��p����p��p���^usQqo
R{J,�,]B��ʶ�+o�ߟ�F�ۣ3��w\���e�p�'!��j94��hQ;�V[�*('���*��hud�jf��?{l�Y^X}�%�<�T>U+��j3��Q������T?'`��wтY�Ĝ5�/�*���O��e�jy$��Bc�s�+Ql��p�����>d��} ��&�J��m�Zܞ�4�nY{�k��V�$����q�O��x��0��;�4Ui��s��S�y׈��w,[�:dm�����?E�7:'��h� ÷�}�B�x�|��U��[�U��.iVd4��Qu:�@x�ז��F�l�,*�sWim�VzP3��w8{,��K;G1�]N#�/����>�.���u]���?_13�3WM�tt���{���v���4w��D]٣6�z����-���v��k�w��f8�����]Շ4�ABn���y�*�c����j:DmJ���3q�� h_��F��|�����J}��_�bu��zGk�Ƃ��m|6㊹&c��<��_)���7 �v����թ�p�P�XP�a��8w��9�d��o��⫉��� �2؅)>22�b�kA��Yx�h�,����o�B�B�~t �C|n����ܡ�w����%e����n�z�z����GoWuR,��dc4�]C<��nWG�TOЧQ�@��r[U���(�VE���fg9�1��RQw77H��%��P�o-�{]"\g�"���=?%�(�Mt��j�3��9m��2�㻋ò�w^�7!Y�د�r�[�kly�
�~�"��4���G�~
��jڋf��6罺Z������蔫���f8��g �_+�S]a�P����y�AW^��xq�J��"�H��%�oF�iƆ��324�S�Z�z��_�a'ԣ��o���Z�nĻ�g��ߦ�ʆ1�����BN|�aR���!�P�4�!��B/�f}��N�)kb�z-��+S؝���b��2��1�U���R���0��P��t�&�5����HnX7un�5���]S>�]�7�8�:�i�[Yt��qI��d�F��lqAA4�CJv;#;o�*ⲗ�o]�v��j�.�Y;��|1�Nh
MNr8u U�p�kS�ӄ�z����	ܜ����U��[^>|�^7�&7b�KF���%a�>�,��6_�f���)�T�^�z�3c���Z�Oqׇ���=��0|t"n5�XAZk�g�`3�S|}Vk��b�}�t@�ջ�D�2�t/"��q�-W0�_���<�������X��c��O;�z�.��i	7v3���A{+K��i��}_=�Ȝ����!�7��x����oPVgL�ȃ�(3�T˦����;T��40�L�>BOBf8���]%�G�ƤeQ���
��;�0s.ņ�򗏠���ï��P:�܄92,@Zo�\�4:�Yf/z��֧m�I ɯ2j/�?>�+��|�.��hzu@��#
��p�+�q��T6c<�+�0ת����E���sPEk?/'�Y����7�\��}>L=)}�_8[�ϧ$ĺ��V�g��$7��Y}U�WÚ�=ʊ���N��Cl����R�`ܢZ�L>%�k�	���%dw��8�s0{ύ<-逄�vdXQ�ksj������*m�5B��p�ja��h.=�g�;�;K{�
�R�Wԩ-�c�]Kg^닯��a5g�� �Hsu2h�G�q44��c�����i��Z�eC�\�J���Os((���53�tS�s�ZtdwR��$������XƇkfWN��ݻ��)y�|",;e�����{��;�iP���{��:h}(q��� ?_ۮ���m@-��K,^��cȭ���J���|�3ݣgDY>H��I���P��y�W���{�(6G�Ot���P���M1҅�c�|f��kj��A��m�^*���[˦���r���H���&���O�Gj�O�:�>o�1PS��W��r{���UL��H�1���a@��0-{b"�]�\W��*e�C�5�9�HWɦ�g[�l9wUɼ΁�H���N�_��-�q�M�^�i�dR7��P�/x"0`v��Yӑ�f���2�(	�݅�<�4���S�5��yq|�����AG�ڍ���5e���96y͵�^��OC�Ȗ2;Cz���T�u�PK���GOB���EX�6����l���z-�)��)jL�I��9cs�M����I�@�qA�����+��8S1��fl���ai���J/�'O�؁��]�93�T�;�G�Ƶ�"H��k��S?r������~��]�u?o�26y9�Q�����2��a������x��޻�fs{'X�1[��,�h� �qU%��Oh�c�	%\��X��F������r�7�l+�Z���ﲺ�ے�]nwjY�oe9&�����\xix���>s.&�)g)چ�<���p�^WϠ�3�zD�`M�1j?}V]nm�s4�FǼ돮4���v�8��?Nt����0�D3hNXT>ၷ��u�$á]��#���|^�8�w��CH�qcjU��F��lT.��?G%0��$E���]�^��vT������^�Lk�lh����e۸��D���Ӈ13	�1݉��5)�;��/"xz����6�j0�2>㹻�w+}�&<��>dE�o�75DպG �U����������%�I͒��a��R���5I��bS^��,�qc�D;�c9M�Z�bnp�h{�_�k�b1��RKC&��,� /9Q�D]	��R�]O��1$��g;:��E�,��)�Ŭ�2k*��Eo��i�qp���pJ����#*#�#V�ۄ|¨8$H���j�]��l;���~��V7��|�\S\���9�Wc�r�����7�M.ل�b��iEh�>ĸ����v�g����"o�Ӥ/�J索Ӓ�Eo�l5�s��疦y쭶.�����p�����Z��Z�P���䨱w�M%�U 1.�y��+P���`tW5�̫��zIaUs��V�Kַ��-fǻ��].� �3���]��|�o���5_LR��̋��j����K�<Y�p������JY͛��o�$���w����'�8BNb���݂�nZ��)�}>�n%y�^[��_US���k���5"�o�/�4F8Pι�K��6��K��c��Pw�S���8�i=��m���� fi&���s�ǼϬ1�l�2�L��w�%�����B�F��o�WPj.��w_������%rZS��FK-Ͻ�}!�Kk�RG��h�^]�T�~^������؈1~f��
����S���w+L;�9�8l��(�j;����\%`!�A�6���m��oƺf�0��\q�ƒ�ƄwF'�����y�#hK���T!x�R >N벇/g�3�U�E�*��p�l�ů��ne/�7e�O�UI3��FO�]���^��wnl�s�f+F�g
��]��x
�B�Ze���O���ۗ��o,'d(�%\�.�f(7w�5{�-��L��v'R���Ѹ���IW���bКTw��}�wnP�[�*2wі�9�������d��1��n�
�sh�cW�<�"^%��L;}⃳8�TY���c.��Fs�&���L�:܎����g�G�k�K�|�m2�M/�lȲ>�3�����.��Y5r���vfՀ/*-��;P-q��U��oh��Yfp�к�� x�¸���I�qg8��N������>���-/
նVF����K��_a��� mx�]��Q&�Po���I�3�~�Un5��iZ�N[�4!MFF菷���oL���ԡ�rSR#;P��Ϡy��,|�m�VF�;��=P�5�9N���|x��S��#S.=C� �������ɍ uGD���w!,�,�n)���B��갍��r�A�G���q~�d'0�}Gg�)�d�P�)x�#�\w�=��4Z�̢�Tywr���R�/ѥL^$��4?��=������L�-e��/�B\�]�l�a��ܡh�f�:�^P8�	�5��wA.������i�����]uO�[S�Eј)Xk�i��6#K���+�[�r�N?a����k\+.��}&K����K.�?*,S�p��	w�"�W�#P��Ӝ�d2%\ᗉD���l�5[��(��=fL��:C�W�eqB����+M�i�;�R��}�w��O|��e�<3ǰT�?Dg�J��fאO�2�S�=�Q�ŊQ]�C�2���قV����\ h@�{L��ǪT�8כ\>��}C���kH#4��L���#Jj�m��{xӎ���Y�*���!@:��ސ��FL�
�7���w��^��Y�=uqW����S�߫rJ�WΖ�4Z֧jJOu�Q{��!�+�i�{����td�h��s�њW��`3��Rٽ��c��w\ĳr�N�v[a[7(��e�nC�;��r���{���v.�z]��7���)������A��T���59KᲷ$ɝ������SQ?��tW.�6�ّ_[c�	V���L��Gi�3�B#�(K��dx����,df��a�k%5Sj�0�螪\�`��.��^�ޗ�|��}����a�*p�@�)��7N��B3�xWEc2si�E��(�݆��z#����P,cs��5C���X��x����n�%|����TU+l��`T�[ȱ�ݝ�2sW��y���dNP}Y)�u+�ć��Y�{c-��7�S�
�Vk��v�Hq���׍�7��,�Z��J�o{.��u�xs=��ݍP�N��<�{Q�R�~�U�2��P�QV��vkū�M��,���س�DN^��c^M.f���Fy�8��o,]�ʈy��kU�,�!*6@��F�9-��;M*�y�S�m-*�"8��E�`LG1�US"�<Q�cb��PE���y�(�:�-G���y�'�ΐ�L��d��[�0�؊�Y��i켧L�-��*����:�rf����d������!�Su>��s��u�����8#�k su��eҮ/�nl�6�ܔ+}m��<3����c�wc�sJ/�C^b���m
!m�S�܊�2��.���}���g��s{P]�Q��ޗʽ3�Uz�\�n7��[��EW�yA�����:�c�T�vLz*��Cu�̬�qԤ�R��m�[��ǎ����;Y��>��ou�$1�n�	?3ǲ@����*_���W-�%�F�U��9�]v(����_"�q;�#4��Mp�L��J�b��a�L2�CIxfԶ1��>����P��u�uw=�D�����6����G5���Y1�:���b7T�x�/��,`c͚��i;��F�*����}w�V��7��u�5��{���"��J0/�P�0���G�yB�9�G�!�~�>p.~�ɨ�/Vٯw?���?h�Y���п���w43��z�B���`\�ud֢$���H�%����#�����]���ȟ�9�ĸEF���=*�꫘���ſ	�ެըL���,8u���yd+@Z��r���\���F��
*0?:�Am��)�~0��o���0�p=I�������c�����̡7��C�����.��yՉv�l��ǳ�\�R�Ι'=%C��L,QA��o�������C��N�JʊӸ�j����'#S[�)�^�M�6Z�a b�Ihd��n˃�6�E?�����$>�_=+�1W��IR�bah��3]{`���U�V��J���C�;+�8g�,=y�Mww'�-K��W[�;}��f�0�ᛍ�\<�#���[����@h���Z��7]YJu��u��֞�&8�f���_��j���!�OY�j,�»�h��*���w*n*���x�F�'����5?��'_��d�Z�,���=�=��Mc��-�>J͏\�㺉�IA�֩���u�C�r���.Q�\7��|��~�kڄ�s|��v��T�༟6�L��:�&��zb.n���w~GM	�I;C#��8��
�!f%R�Č�r��"�B���k�����#�]Vq�\A���b��AV ����!�.9����;P䤵����C��q'f��ss!Ѿ�2�Gh�u{��όF��=`R��BV��,��(�7��	�A�x��k�:��]q;��T��~^���X�m�Q�����kmOdz�Gr�R�z��
�b�s���7C㩜�=Qs(KOq��C*j{H�e��'�XL���d��,����k�b8�zr���BC!~_�(!��̎C��~���.��:dm��0�͏����jTW��lM�Wq��]f������N���Z�\`��75#�{�=��5���P�O5�����3q��%vN�o'�n�G!^ �a"n
�H�����P��o�v��pwkË=K�q��w�D{G����뜜�������O'����g:����n��|�ڷ�����\�כ����hW򵉧7�__1��[�}�v3뾩�_�u4�yٸa�7��Ӻ��aJv�W����i��lV��Y:��R�Z�Ji<��mX�F�����-�O������nwi���B2`�Cg��C�i�P� p�a�7�$�YÆ\�˅��øc�A�ѣ��s�&��t�%9��\��v�еl
��]=0D�w79ݵg!�ѱJ��#�[�a֗�}{��=��:�:�N����T-M�ӋW��xk�cy��Y�/y�Μvs:�whi+�����Y��7*P�u_.��Y#n��y�s�@�X�U�8�{�g��n�V9j���|)I2�ꂞ�ͳ��=�o)��v7�g�`�2)� ����晫��;a�N��o�c�R�~z�򘲎z}��R!k��/��q�_S�}� �"�@q��:��g�Z1��z<)�����>�vkd�9��˔:(5�ڌ�n��.�yW�_n�g�Y�q��u+��336�:�0m��\��vV�hY�IYW+7��S���)*�W����:K��t09:�8-�-ڼx)d}�8�?#:{*�M� �@�AмYsF�o�{�<�Ǜ�=FX}�1/��Ѹ�����W$�uV4]�Wbf5`ћ��M��Y[��[�@6Luuv��Ѧ����2-���\�6h�].��aVH��sc�q���>�eQ�~6@�E/b����1ӯ:��J�h�č.[�)%�x�)ײv+vw�Wq]]@�/8��Y%�L+��[}����Ѹ�:�۵���#:�n�=�C:]+w�M��S�1�)F,������v��H������ӹ�u~}�;jpge�����w��5r��k��[��_,��S1e��7qɆփ�4�Ҧ�S�W��Pz���1�cS˚�]���T�=�tgg����x�}��+��#��zT�h�)��\`w��,���Ɇ�77k�y\�B��=�O|�1�Y������	x)B*�܋��ERSa���ێ����8��H����GC�-˻ݧ��j��f
ud���7Z4�a���Y�ƀ��Mjдm�Hn��|��c�d\-[_kPά������\�C��gx=�;��L�ױ��e�}D�7�y{H�Q����D�]S;M�bT���}��[�Ej����G;�Ŏx:��5��]Y�Fh�`3v��T��ʓ�w�)�����ȩP2���sT�u��i�`5:���.�m��Xʽ������6��6�M��f���n�>Ŷ�z���]�-:߷��tZl7"�5�,�l�ϯ[ށ�<e=�ɣCG��X����ړ�I�^�����P�\xE��	�_��4�.��������+1gL�`��V7q��^��d��X�P�z�:�[�$ �:-��i��\Fd1��wR��
��٣��u^N�mU���2�NM����s��̕YU�ھ�P3L���7"�X�"��(1��ZU���*,M)X1k�ݱ2��EAr(=R�u�m�L�hU���wʩ�axZ���5���X6��uə�+��[k˗+jҲ����5�6����&t�Ѡ,*q�,��l��fa�3[R���m���A�Y��OIӑC��FШkKq��v��.�ېօOZ�T�^������q8�C�A�颲eyiu��[d�S5�b�մ���Q�۪\�8�*-�k^�U0�T��YX���q��n�mX�c+�b�QH���S�n�9{�E�W��E�����#m����YP�̻SU�X�f�]Ap��*�BqܥQAy�-�����bʣ�S��9B�b�+P�����!�t�-�Qb^5���"�آ�[d�J)���Tf�h��r���T(�L:�����|�|���VM��}�x�Z�D=|&�x!��H��C4 ���ԹE�WM]�����R���gD����! z�G�1���a�89�T(��N�ʀݦmcCv}��Z�ɸ�mR)��[���܈���W��f!���%��"�֖Nt���=�T;Ƣ����Ų���<{v����N� g�n1�u?d�n�
�sp�t|u�1�ߠW{}[E>p�ى�;}QzvO)��b��۹V��A�D���p��z�b�D�f�������T�,%{J-��:ԈȌ��3���31Yθ�r'i��kVG����k�Z�=��{�ɦ�y�ò
�_H]�P<�dƞ�!C8hwC-�jZ�{�/f_�f���s]^Z��~�B��!��E����<5�Ĥ����hm۽>+c����ci�6u���:�A���}�^��4+_^P�>��V!n("E���V*��ߤ�f5�]��e�u�&N"s{*�5j��<AN�2h� ��S�g,mɛɊ���R�p�|�W��F�k������6����2�tQy"�z���>uSڞ�ǩ�z��1����"��}��Aׄ��X�5�bf��e��.I}�|�r^V(yr�7�eN�"[r�
lYɜ��!:���V%p�y�,z��,���0�oR��tk�#�vLs"պnu���;�:��� ���!Шˆ9���*u�ԅ�����x)ғMl��j<"ǝ:�M�ǰ�,\��ތƦ����Ug;A&�����L�> �_'�U|hÊ ��
3��^��(4d��@��RQ�M��}�5.����n=��;"��b[^Nn����b6���זGs����vϬ��P�U�����޵W�'�D�ؐ�8$�yOе�P���k����僩A���2�����Tv�ѵk��!�dp��Ax�7��Q�aƺapZ���2�9�֫�:Ξ�b"����B��V`\��n^j��I�mqZW5�s�w��`g�Q�s��!_^
����>��*΂[_�=2�W����N�~XP/�W�	��&�j�_f���t;MsJ.��>ꁫ�f=i���
��3��5��@�T� �0�t���E�k���]s���m�𵁁�j��r��X��ѻR���2�A����VC��`�{��=�MV���+�GBG4�6��VV/R�C�)��=M̛5�g��6�6Ί�Y�.w����}�v���O�9���4�64(�H��51�w�֟�ۯ�c��]p�9����^ͺCG�{ϝ��7�<,�!0��_�|��D�^�r��[cP�[r-FP|��U��tN.ͼ����n��W-���
݌�-��i���Z���mVP�F��.��]S0���z#pS�Wg�ttjq��qW=�ܶ��4����O'����ıώ�7�%yb�r_E�;�z&�dPK����(�hu���|�L\
OO�ٱ�F�O P�SE��Ye��Qmy�Q���^qy0+��N��7��vȪ�:r��L��Y�=��>m����h����i�b%:`��l�����w�##��0��N�a��ت��{fUUN{KW(�Ж#�b���E@q�\S�U���R~ktsg��T��F�99��
�z�����А>�*&�<y;�}h.��o��Cz����W'�>]�<V��T���sg�x�4+b����C���H��2(�,��^��������_g�Lg<��9�~U�n��sș�K��oc>r��|�ԣ��;����wO�H.;ʥN�k�Rt���6E^3W��*u��R�����{�_O��\�D�ޙ�;<��(���8�(�%\�LƬ�^����Dv����)���l����/u�g݌�d�}��.~oK��� 1T��p�N}i��rj��W0@C�l
:1>K�9�r������
�n���q��9�1��B"2�+�?\������~��^U��BF:�HX������ �ʁzs��WxfÜ�])�0a|ۓ�{��5&w3iPk_K.@�� ]�9����������sq�$u
���6�e�!�$���0%d�w��Z���}Bw#k���ɦ���Up�B��cRO�ۉܢ<Gg��-`A�o�<+�
2���3��;CF�l�8-�KH �R�3��L^=U�c������W��d�y	1� ���\[U5}�2��3Y�VlozQ���:�E��]Rh��=��k�3^\�)���j`�K>5�I^��H�'�I�&��Uq6��i��ݱ@<�����Q�|�u۟��fע�i���a��"/�2Mq"���n$W�t����;�7~I�i���(�G��F:�s�o@�s���޹���v'#��Bp�y'&��PFq��ӭ��mTAw2�Զk;dtO�Xފi�ϵ�5�ϨY�*�W�s���8�gJr�+���#�G�ڢ��x˶������<B�\_�J�ρ(��WH��Z�n� �a�jya9qjXc�L�c���aX�� �\G�I�*��"{����"����^�MhfƘܝ�KOMfB�|��h"�H�t!�8����ІW��3�4?����+K"]�P��^�cn5	芽0�j4�L�ܺ:[
���/��2��W�.�]�>���wo,�q� [wG�������u�՞�H�n��,q{sU�֫A�̱��nV6��2�{¾ݴ�b��_t��C9X&��{YcM�3��ހ�Z�I���E�r����z��G�ߍ�4尒}�[�jvAm�v���u����3�+3`g�I�����{��O'`K|7�z9r�S�`ۤǗ��	�s�Y%�A���sa�dc���h��5%�N�47���aS�y<h]��F���S͟�����l++���:w�6��ދM���N�2{��`�'�����J���he���N522-���*� ��D�e]��:X�h�@:��!"r
|���ύHO�c��k��~��Tm�WD��!#��>�_d�bչ�+�D�y͘�Sx�D�aP0��%��˃�ޛ`X繓�����۹"���;�r��]⫒~�����ܳ��Y�R�j�Ѩ"��q�ho��N����Mnn�Q�7���l�QA�]^�/W�BG�2Z��`?z�o�L/:Gӫ�M���qY3xT4����[>�U�31Bj�uަ��@�g��=��j�N��H��e=[�?H�'����q3S�g���Ј�� /J��SdW8x��%��:W�-o�Ȟ��XE� ���X|a��Fү\�ir�0�D$}҈���[�z�� �eW��V�����L�S�S\G������X�fd���{!�(���6�ԑ�MWe��QE�(숺5�J�u�!z�FJ��f�He �K�Wg����f���
�E��m^���ﲒ�z����ʙ֢ͳ��A	O_H�7���ݪ�D�Bk�]b��*��N�E��F�6Om�u�g;�V>1�,����p�$�O�]~��1Y�Ќ�������;�1wk�u炾�P��SLez_��٬ӯ�8M=$��l^�W�6�嵲�bԅhg�+P|���{~��]Q!S��{>�[u^��/��2�x�/�7c�����LW×�R�b/���p���ٌ׍x�nY��§-���'��٦(=a��xԦ��Ԧ]����T��,��^��b�{^<[��2u��BY��|WD�0����C��h�3^����b�_0��)�ts�������A�~���˞�r{H>&,%X���~<�3r��G�;8ػ�qV��oF�V��mG��3[t�].k;R������3�>���HP4A\A @N7�Bֽ�X:s���uSy��ְ�kk�U,�f#un���/Gy`T����ʂ�1ڌ�,'�W�a���}Q%����S�7�=ق��}��j������f�|���S��1��@�0}���5U�ې��+p�Of�}SD3���x�]�"��u(�{�0����|�'��E#�~�A��+qt{��7�Gj����F'ǂsi�a�]��Ѩ6�|�ݡ��Q����(%�?��L
7�}��g_K�׏�n��RP�Z���.m���g-iy䤝���S�z��V�s���]c7O�3���dkj�����B�H�|[]A�����kb�C�}ƣ�
��1o��������
�4a�s����W�fӜ[��w���k��Q��n����@�&��E�65�fL�'�Ù�����ؔ<�h�R�CJ����7P�E�K�ɦxȗ
�^�"P�S� ��2p��JiƼ]綳�΄++elE]Hߍi�eC�딋�$�pM
�ИF=ҀT�O�+54>�3��FV��к���e���k���ٳ�o��X��4�E'�f+%�$
~#���Z�fLJ�[:b����r�X�dq(F��
�t�e�L���M�Rˬa^*.2^Bu�~��Z�ӊ�C/%�p���b��������R|xEG5{Q�C�rz݌��H�/=J���K{,�0X��F��0��/��8;K�~;(��4���E����|a�
�=S��Ö�DB4��T��P��x��6pT=C�c���c�[�f�����7L׹�V3�#�tw)N����e�c%P���61F@�����K�6�[���G�[�Fe���
�'�&���Ebb�ۓGC^��Yb
��p��0��F��}fl������JՋ�۷� ^���/z1��[��Ø>���i����n�z���tƱ�;7m���{�B�.����;˭J��Ӻ��wޣ=��(b�Շ{�6�.���R�% ��%���Z�y���@� ��
��[�����w^�l�u���Cܱ�1Xj�$v��z�+58��ic����:8��7���3��x�n���f�8�F}s�ѽ��ز��ơ}���^����Q����m�<�.�j��43��k_�g�fn�uZ���GvtZln'�Y�oa�2i����^���=c���́
��}فnu���ݛ�É�V�~�E����a�*�
җw�u�5گ3$ߢNF)��6����γ�I!��,����]��8��7�`��B*��}��r˱M�oVu1�y��2�I��n��V�[]���¢�P�}����몈��VMm9:��V�r
��;ʡ�Ҋg]�'){}^����\R��Z#��<S�F�ϋ�̈́�{�8�4w7�t�ק�%`6�ELJ�[��q�&�KQ�yz�]���K:�64[�W{R�J�t��i�;8[��_u����Z	P��&q�8�a��t�ox�K-]N��W�ա��@p���Kj
bEf͸���8d!S�i6���8S�:d�Vs���.`���UN�wvLv���q�cC�T�>��fۂ����Jk!�G�5�����0ח5�'�_���j&�$����,[JP&b��V�D:yl^*��V���g��-�&�G{�u�A6���=�e�oO�´%���N���"��2�K��t�R��������<�����#�3�֮��wT�_�ت��Ms[��q.$�u(Р,il��ͱ�Jz��vE����:n_�!�}{�g�cMSo"�2U��7�֦ع�X�U4a�Y
��̿�ځ�V�1=0��tYdꤳ��&\�L"nmMq���t��ȃƃ��P2Ǝw�\+8,�������B�C�Ua���ٞ��G��V/GQ���z	>z6��*�A{��m����l�dI���;���⹟�E�Ɯ�V�=�v%��,>�V[]T�z�V1�HΜ���C]q�w�#����CZ��ӣu�O�a�w�+�M���?�;��u�������sݝ��Ν��e%��
2ȡ{[ܣ{f���3�Zu�}Ƹ�kt'����R!k�y�3.0c�xqW{¯]�Ȼ�ɹK��u����u�]�>�Kcٙ/;��P)�Z�y*v�.�Sj��fQ���Zy�f�SY6�`W����L��Yx(�^r��Da�������.�[����t�׫3˲
=�	�f��\�TQ;�,��O�ӊl�㕤��8r�����9�P��itªˮ��MK�q�!l;���}��WQN�+e�O��xlD����o7{l���K��l�He�`m�!<]5�*�yasM�^��<�[��r�fD��5-n0��d�ZB��-C"�ЕWz׵�w`=�z�2�I�-�[�J�
�k�2纷�Id���;��� ������s,�{��;�ʷ��ƑW�]�+���I��B�ޤ4�<t��F�܋�w��Ϻ�v�;��j�n���-]⻊�ݶk4��%���Uw�yur�'�=@�X��z}�1zg�)>PY�H �{�|��g������}>�w������,�]N�9�y�|a�5�TNa�#�.i$k޹7r���N�}|��ݔ`�;%kv�=�9D:n�7W�gj�tn��{��/Z#͌ʙ����Že���3x�;���}T�R�RoXu�)o�<}{ ��{�^tuY�mze���A��"�̖�S�,v�/�l5�҃Je�EY�X���[y��1#�,F9-����wf2u��E�X��؟YTo>j�;l)Jn��8���N���� ��D�ƺ����Q;���'k/���-?�AN�]�(0�K�J�To
�;���}��4
�/C
}�7)�W1n<�$����U�(]�^*Q��L���n]KN�p#p�gsx�A���	y }R���V����+Z�oT�o���x�@}�C�
G��;u�&������N����gp2�Mc�������.S�����tL�u}�i�k&�Q���V�ۦU�vo׶�˚�(���|}�G��얐�w�vX|;*��n��־5h���7������R��'��`�'�,<@B�\7VYJ�ݏSFo�Ӌo�c^�.��o?�W�]�����EعXj�o�P�8��{I�D�0d�-�ц�]�kq6��\ ;Ø�V!���6\KΑ�qWe?q���fﮆ窔+�凚���_Ή�yqi�r�"V����Y���$���ب]:�-�HgZ���tn͠az۾3{+S���h�o_���w�+;;�ݨ�m���Ǜ`cܩ�꟝T��Ξ�yU닟�@�������W5s�r+[�(����ZUl�C�P:���mhS�nb�ٗu*^��8�(�����ᮅ�
���s����`���Od�!�!�]"�eJ+(�K^Aw�S�|���a�p����)m�1:T���k�Y��G�Uu��Y�[f�Q47M�� ��(��Rn�h��M+wk(P�}*S5��a9�s��dX��X΂�ϢL��U�=y�?r��pՑg_-1��Ȝ���E!I�3��y��+s�h�1���EJ��Y�G�[�9�� ���O|_�C�Ç�8���g'#5e<��36RER"����<�o(�Z����5�9����	b	�̻S�ۻ-ɴ�����٣

m�ժ�fJ�F�.�R���*��%���E_��l�Z�N ���`W��cI�%i�����R�T��F�Q�}��F�ݮ���{�(�*��V�9n�V��1,'K�	W�A��ʶL�4G�f�
e~�r���{�؏L"�*�>�>����
\XY�h�:��]����{z�n�L�O��ș]����o��\(�oY�R��Vm'�1��.h�3���j�`�+��)k�G	wH�q��oX�:��y�7~Y���^z�κ�ڟ��b �=�{��b�*\��u�n-*�ϾFrq������C�c���ii�����L�!��АIQ��OW;�\���G;�Pk������b���{�Ǿ���J��i�w/V@�Q�k���|�5��)N`۱}�ۓ%C�Um�93�:#��DqTl�*(5[�Tf���ֶ�B��nq���[R�L�9X���,Y�+X(V���N2V[W� ��qfs�m�|N&C�����[E�������/%�d�����qs���� �m�ɑe�
�[�m5�����gZ²����Q��\�(ʛPե�bXɮpd��U*X�J�8󒓃��n)�n`f�j�m����T��53�a���6��ض�U�F�[ak�ɩ^0�8eb���rQg�88��l�ǽ�؊-DZ�Zzg��x�ݕ2Uj[�ڪ�[v�J�dX�dP3���dS0���b��&8�ۜ��Ֆ�J�-�h�ƚ&fuo��%ME����cL���93^�r�9��Qb����"�m��Ѷ�Z��>���J�������*[N%VC5_�5��~p�~�寝��Rd�@͙݊�fX�&��2t���ڲn���Kꆝ��}�B�K����s�8c�\s}�����=m3P����ǎ�6��sρ�o4[�"5T=��I��νa�r6�벻��z�f��v����k��o�t���1����06�+��e�P1>�9��_a��]�6� NSOǑ�Hn�cin,:��=��X7�u^糣�gg�l��s� ��:ݍE��%H�Z���}J�:;p�SW ӯe<ZV.;}�n�n��2|y�@F�eK�S�4�*����k�w�6�x�|�0��5U�d�Fi1�͇�&d;}����}����R>����)Wz�`�jE)�Zc �h�����B��W;2o#EA�K���P�L�������]�<�B��t��]�>Cz[�J�ݞ�=M����$w���I��{_7yU�ҏ���7pU��Sy���㋩K˜�|:��F}�pSY�J���%+U���n�P0�&��n�y�2�`�����1˥&��U:C�ېYozY�*���:��(^en�$K��z yޫ*���.V_wc�ҲH�����n�{w���Zzb��=]R��f���"�l���Z<�1L�+�q���Xޅ}�WM���Cc3��pb϶�;�1z�nZ�>�k~��>�����IObJq}�9�)���U]����Ջ`��Gz��K�����u�_m�6�!q�3֛D�F�I��7�=W��ס�]!���yDh޷���2؎Lhm'�����檞�)�3b�MMΖ=��7
� �3����1z�4��r�p4�s;xԽ]�Q�&$u�	.�eC�hk�ٙ�A�i�om�2��9��|��')�gT���HL�r���^�`��J�z�#�ӓ�E�yGl���w\hG�=��'�P�]k[\��Ş��n߮���Mv�k�=4�����q ������Fy�4��0�i��Vn�v-�{��n=on������^��a�W��7�\;B�E��� �t���`�@�����ب��Vp򥄝�[=H�oQ-����(5�T+�3�<p6�*:|��5��K1��}�05��fL��Oh)J���狻�+}���,�{����$*{�%U2id�{���V<�#-��Au���u�c�n=��|�6��f�JV�-a`䵉P�^���K��fɝX�{w��3�	[����Y�7���L�=ux��G�AC�(�vs�9>Npk�>]���H��W�)[�r�R8b���jb�c�͜¦y��mD���fU�
Xk�6����bOx����ͽZǌ�+�wVqߦk�E��⫩̀*&3���@�Ԭ�U�RI{n����g���']��Ws�ph{�MZ[6<��r������+/R�d��r�^c>ÅO���n�skc��V�V�B����AL
ᔳ�>�h�%�67rkjڌ��Dk�<U�=��1]d�й[<l�ݜ� 9Mr#���|�y�.���xgv�{��:��_T^i�.��ef�[
���Tg���2���ޒ��YH���ɷ���pĮ<���F��6���ϻ%�`h���|={K2T�����ö���e�y�fOM�2�r�[��:ycKd�1�r��w%ď>f:D\t��!�T��f!#^��zf��Z����rο=X�Z;����P̨ڍ
��4��G���oEc�w���-,�ND5�m#[H,�I��v�펫�4Cr��'�3 ���*:{UJ��g�pڃ���^�CzK�őԛ�Y�=��yg��������)\��*ekE����(;��w_ʪ������xfv_��|�8d��Gj5��x���tN���	��q�22Q�a�oA���c�Ձ�?�O��V*3WH��j퉔r�ҡۊ��s�VT��N�v���3����,2C$�e��I��sx4�վ�����z��̀�4ds��]�|��e�N6V	z��1������҉�42[#�Vr��qH^��{�Ď��YO�����uc�j*���S-�4�=�LM*���Ồ��M���$�w?{h�y�����efeS�` �=�}�:�UO��H���ٴ�w���)ye(mY���syI]3Y��^���q`ϧ��#{d����KWً�C���"����á�s���J��[��aÚn�M�}&����r�.�׵�U8F�÷�vK��w]��ǌ��R&�������?������wi�bP�|�GVNp5�q���)�ܘM��H%�#��Q�u��_D:v뛬�7���;�z�0n1��o���p�˨/N��{�nlښ�y��*ኬ�٭�LX�{���Xq��S�F>��Tv��L��.h�|����ᛰ> �4�4�m����4��1��A��Vʳ�A�ǰ�0���x)R�pr�vY�ܓI��uv�Aa�.�/vY�7��q�U����uk)�_ad��Trޱm�U��E���`r<�������'�@�$�'�)s��tf��|�=1�v�J�O�Ў`�{zD-�����큸�T;ͫ��ج����S;�F��`l�=�|ue�#飼3p,�x�7�-p"�'3�\�$>0i�[�q���/+V�*]!�W��Tv�}����ؔ����ZY���F���=�u���>}�TM�H�%��9�Ɩ��a�v2�t�@��򸛮���y06Ջ��;!�����ZI��H/!o}�xԚ��n�tR9^O`�C��Sb�7wZF�:|_�}��+��c����1�S6�'�vzO<CP�O�16n���w/"�I���aUmqY�:�HlDe��0ƥ�P��7��8ME�g�����2r�8��
c��7dzF��U���Rǎ{��y0��Wx�G��L]��\�i.�� �,B�a;��.�ᘧ ��Ipd���#������;��sUs$Z	5���#5�����hy��T-��wr�ڝ5V\�]��Rw3�z�G����ɥ��-S�xl�{�X�V�&٦��؉Yr�UWP޻b9nk�X�!H�����c��P{������w[�.:���!YN��t����Ft��J�%)PY9#�Z��#u��Q�_���-�N3�8e�a#���t���J���~*�R���q����˺���2&,�W1�H\/3���������?{��9�KVft�v��˝��:�Y�����8G������y\����{��B.h]~�)���uǉ�:s�/*��38�����l�^���uN����/2�g�슻݃ijK��	����6n��~}��19��׻��{��6i"8�Fr��Q�62����oύ���x��P��{&�5xי�n�K9��$�|5�<�\5�]!H$�oC�]���d�#�{�N���o��sV ����H�i�7�*�B8�b���m�:�Un��ԥM��ʴ��ݰ��j�yPw_����f�M{�\3\�a����Q���y�J�'��Y����9�Ĥ[?����o3w�ď���B6�>�웅�[��kh���гͮc*`e:�KYD,��1�LK�3������^��Xp]�x�{���Ռ��2�\[���5S㻺%���0(>��N��8#���Ε/D���G�wT�k���l�Ghq�;���\�k�2˹L����{�n�m�ףL�F^Fi@�(�+-�09�r/�yhz�d��˚^�L���g�s�kl����؂��N�:Qki�{�%}�WeL�0���Κ��#�-��«{`\L)e�
�jVQW9A.�T�mE͎���^p�@����bh(e���rS��:��Kj̜��v9=s9��t0ڪ�"㦬4��C�W�6�*��xE4�0S@������[��gEen&hy8_p��������ʬ7Kk��Iݡ�n�5�!lz� y���jv#�C���sCL:�����Z�*R���h�0�.���Z&�^\/����x��ǵP�uJ�E�����Wz�U��,_k�is����u�r�1�;4��㚹fh�r�
��k��&�{�~�I7pg/q�ˏ��$���g;>�߽9�לd�V�P@'h�$+�G`N��m���Y����3N�ܓ�IU��!+2f��cȾ�#zW�i(��t����Cd��X:�nZ�$>M�*.���ј��#`m�T;	��z����	��93
�)��9��E�S���&�D�3	�<��(О}��w�E\�����+�٫T��2=��[3�B�ML�}��LÄ�Q����g��~���e93�w��7|��S�n���]:��g��c�1�G��[8U�w�"b���0���lQFkۙiĺ Nz�l��-���FK�s<0�q��I�2� (�El�>�蛛�38F�=�v/�a���PЪ��ʛLx瘷1W��ܦ�ͅ���y�sjbj�cF�n�zx�H)!�J�j�T)�tO6<����6�v�ħ���ҟD�]x]�fy�Y1>�"2O)��>�OL�\
��vLҝ��~~��{�Y���L
v:D�`ś�e�K�;cdk�Bk;3�P07Is���J�m�'��8�z�O\u`�xo�U�]Y������U��T-�L�k�1O�4i�;X�J�|ޤȩ��ދ��*F.Н䩗��7MKo%N���2�?D}�tT�k�.>>������!�T��jc�T����6sa
rh�e,�n4&:+,���m�q���[�D�c	�7��ؗ���wط6�����u��뺫�>%�1J�Yy(&uB�B�֮v6�L����C�y��뺡�Y��f�g9�)#aml�Ur"��nj�6)��,�PS:/��x��0�q��[Y��볭@rFX�T5mwrY�Q�rj�b�l��&:�:�q#x��ϐaʄ;�X����q����Ż����=�@�ϻ�f;p�Ў��<F��'���fͮQ����i���7ʼ@$�p�u�jIOݡ����/�y���a����������jfh8.վkٻS�4ov�Ld�k�c�b��&�+Z��3`,�/zb5������^�k�a��d�«��v�E�B�xz2w�ǫ�A�wR>j�#ґ�m1Qp�/NE���7����I�#��Ю��N<M���
���`p�;3��˼q �:BgL�%�:Еw���ӓ�{���n���w��ɸf-���@�x��H��n�4�v<���)�νe9	z�t�w��s&�Ύm>�U}U~�qy��.GO�z�rc�����:	�n<׋���\FpΏ%մ��X�Uv�b�$\^k���,���g���Hn=��~x���j�.���;1ˆ�rn��NBx(8n(�3��;u��Kq��n��	���5=v_��b͒\�mD����z� i@�����f+�V�����1qOV2�Mdk��n��\�H�mql�.�h�O�6[>"�Kś����tS��T�[�¼��n��UE=|o�KhqY[~�����Q����Q�"��ғ�_�5�)x����+׺��7�SKeynyel��+���14�>��a�����#F6.47���t߇�v���_c��Km#H���hZ�O	⇘��㳍X2��:X^�'���g ��K�s��~R�n^�R��c�zw���{�{vMo�@���
�+Tns����|�>�7�������}>�w������6��f~���h���
ΪQ�7
���)@}Y=M�]�N�p�ˬc�Ιr9�[�-��-	Z�kz*6q�1��;���]����\�t"�ǳ1��jա �(��� {=�æBzTǝ(K�>�w�� y�03�.լ��FA���D\9dӰ���
�|�ۦs��y��[�4[���٠c�[y�-&���x'�;a��%݀H=tj��za�ݕ�[�9�園5}u��=��Xu�V��B�lLzr���ٿ'N�\3c�F�)"�KSݨ�B{=Gܔ��}Ɛ6���k��뾍-��/�v�=�>��<���ڰv��>�>0K}��~]����ߦ\t^�V��_7-�	��M���>���Z.��:gss�/g{�h�q���G���I�9����B�ke'�!��nI�լ�\�����hvr�, p��7tR8��a�W�`w���]���_H��rc/������;�;�d�̺�g!j��X�
�zo�>��b�´�i}t,Wi�3��9�;M%��*�6��4�R����hB^@��]\�C3�7VG'�ߡ�=�9��Oe�J8E�8dC=����
צ��w�W��@;�k�
3 �<7t����;܂���O�ڰ��x��t�v ��-c;I����ysn瘸��$G.�KYV��	ǯa;P�z���ߝ��PXA�ǲ,A^��n�|���@��VdK���IhYp�����7���X݄� ��V�e��ĵ���NT���Sưp�k��p`����@��<�wFs#Gf\W�'J@�K�W����u��B��;<!^�����y�2���>���6����syc%2�fuKn�J�ݮ�u�n�z�7G?]��b䟴N��_+�ˤ!����&����I!�⳵�����ɭ=� ����ႃڙ��:<�	\�����K�AWM�\NZǔ% �..r�V�C�*��(�6%ݙZ�kM��x�vVC��.b�c�g��v#�Ny^�	���E��h���9��g�3o��T�۬K���<*��ӳ1V�^��war��L���Th��н��Ӹ�!��@`��%��Q�w�ˁ���-ԛ�z����g/{����b�_��Y���̉�I�sP��@��\��u�%>98YˌpA�7��S>ݺ������L.g��������i�G]csd���w�h61�}Oi����+^n����=F^��h�OÇ��������D�u�V̠�S׼�;�
}�mr ,&Z�,�!A:�= jԕ��;=����;���Yh|`����{yM\�z�/�$��m�-��/8�������w�٢7�'g�1�^�~l��4	[����l��Hr���2)ؙ�MYv���H��Xz� r�K�XӍ�J$�����"���U��;l|3�O��2B���RH�d<�N�T�R���ׅJ���m6�K>3kR,��b��x�V׎T�VV�mkF��A�/,8�Ux։R�3W>kʢ[J!X��WP�&�5P��m�iAŵHfe_\ʧ|)3*V-��iY�مF�N�b�EL��VШT�)E���*.Z(V�˸�2�ʅD��#KmV��[(���pƉ`����R���֥T/,���.���t��Vډ�pխ��N�<�%
ʪ%VU�Q��(�˹�r���`[R�5)�(�jn4�:�UQ�lN)[P}�u�,ƣh���#��5KYV��kf�	����.uiF�y��(T�+ӹg5,�Z�m�(�*q*;��G[ѩ�j�ܕL��E���X�F�+Cu�9zN�pz��IU�G�p�)uZfa����Ѳ��E�em)-
�j�f�V��8`�PR�����X�9J*�Z�+����� ��"�y�9�)f����R�ޏ���Ҿ����sj�P�}�ak!���Y��a�k 92Eݹٛ�U�&�D#]��]ϡ}���r&�*4$� � ]�~��m��y�K����k>�Ot���#�x3ّ��-��=�ހ�w�]�Q�ʼz��t��(zr	�љ �}I0.���ϡ���̪Fm�6�j�;��[=���鎀6�go�$u�
��YaC��h^��OC���{��3��oH;4����~�;c7��|��&�����'��čpS@:��{��U�WZ�D2F}f|.V�����r�OVг���j��-�a�j�{y�Z�$�:��v�NI}��Y���[M�scL�0P����w�&��w��-���Br4	�A�ε��S;��t���򌫱1�ې�e�/D���of��4{����v69Q�o�B\��w1gS��ۘ{��Sy�(�����}E���̲R�h�:��>V�'��
�qp�c7k��VᏣ;&&�Ewb�Q��J<F����u<��G�V��æ���^��Up��Da&�-n�TL'4�55W���곚<����;J���h�T}�/:��q9k|�7nP,���ON�GE� ��{r��g--ʗ����1+�sm��rʗ�}-�Dw.eձ�wMf�3��ű�0�Ԗ��x�.�f��v=27}�J�l���]zyEt���%�9�{Br�s��=�^@��n�w)-�M�vzR�]F%󊷽W���J�c֎ұ�z���Gm=�iU���ʷ�f[���\�\2�q�� �[<��ַZ�w}s����n��� �d���+ȟږ̯L�0B�w�Q�V�Ꜻ���ZA�����u��%B�8���KaW^Tg\*����L�i��P�k;xnD�l�{���.�+yHޕ�����S�H�
3�Z�{i"���;�s'�o�D-���om*�vJ�]ǹ�+m�y5'�7������ �e��%Dp�@1�����c�W��-����K��`²[?l���q�+)��������o����|��.~�NJ�:8�z[���9{ΰ�T��wr���dB��M�����>�s`U��}��!�Wi��򫥓B
��$�N�}A�m���-�q f%;k;�N-n$\�;	�hq�$U���c�/	=.��:E��.�Λ�-��Ƹ����bY�Fsr��U�J�^U�)V�q���ﻠ�y�XL�T��QHثz��'X)h��C��u]G�����U����7��떑��j��k�(�C�d�ָ0�t�x�dm�luS؝�P;��B�eꑼu��}���aѓ<�PP�Tvl�+�pdh8���n���K��r�"�<Y���e�x�o��:��JB��[�!�뇖�z{�5�ċ�w:�5<l5�ZV"h����0�2����kv6����C�vK��=�Q��^��=�i�?/���OZ��΢�V[o��ov9���+1��E�#��q���T��C�P�i@�; �A���5!P	OqY�u�T��sM�9Ѷu�-IT_{h�׏X��E�.��Z���dA�Z${��ã�l�/�mnk]�ѲQ�A.���S��m%e�9I���;��Q��d�4��m�&�H�c	W�J�K�e��S���v�W]]K������0����A�&�-�Zq\Y��K����I�#�|Mt�%w��]
�~f��;�n�j�N剫�w���e穋���b�1��~�s!|	���s����������x${2���L�����I���!�3��u�g�a=�I*�'�y;t��B�.;?�_S�9)���~83�W�D���f�c�^�[�M8'K)�my�F����6�zj�$�*�wJ�}�i#0H/z\��{Wǩr�s17�>�����y�/y�1�w��H�il#�l��m��xJ���ӓW�4�6m�H��*��+�sڶ�����s���3�K��3E�����R9��^/c8�Xɀ6�@:w�y� ��W
�F�A��%��n����f=bB�9-�>հ�v�������K1�
�L����M����Dipl
�>���-<#1H�k�7nЎ-���2�M�}��&��9����wZj�(�`���׽�t�-��T�����W��=S{|��+�(�ǭk�����l��&������EQ�~����?�۫P�ު�O����]o��\�=4|u�SM��i�^B�Y��LY~�pK�y�]c'�mOf̖+�5邐�����Z��$$x%��[睮*�2ڗNR	V��W���y>4�!t�J�J���c-؟a7�7 ֎�E�Ǫ�)vV�foa�������v�-��PoMw2�V�����+��5��>��[d����.�C�-ۼ���%E�#�o�
iA�����\ȵn�v�3s4�pC�DqW�׫�4�M*X[_�wJZ�-�z��s�o^N*���֦NH���W�!Foy�k�XAf��[�����h�%���*�
zv��ݓ;�v���;�Z�r�I��*n]��"
hr�vP^�4M�n>���I�lp3Sp��Ut���Iv�IgT"�Cupag�t06!�Iz��h~�ݳ��1�'�����]����ϙ>%_Q��Y*�註���᫸���0�s�b��-���M�<i�F�}���lF�T�-��5�/b�oez�&|{�A�O�L��<��r6�g1s��l��9�n��;K�vj��+,���:��2����7w,�O^�;8��f�/W*���E��:T��s=�����Ȁ��Yn-#�]�>RXw�ˍ�Zd��S�9��<Ӄӳ�|���*t�1����WT�ޮ=�j�6�E�GF�-&ִ��;��9<����Y+bCk;�*��!�	?^P�d�]��!qަR�8�0VC\�e�|��g1l�z��?�AYunSS����t~��pzy�py��^���������i��D����u��"���m���tz���!*R˩�l�+J�n�� x�L����I�J�x�����/#7�O�"��,���G�S���ݙ��@2j��L1��k=t&ȉ���h�~��!E.
��-�Z����L������U`���V3'�ٟU���`ۺ�yۇp^�$��e}[5`��K�M,73��w�LzZ���i��ӊ�)����M��������6��v*�J�ʠU�
�[!��>|ɔ��౥�j�]0�h�����F��r^r��BYa#�G+$��9^D�ڟ6d9My����h��|G	y�x�
�p�X�+6�[
���T`���!��Z1����f��P78�s�tg�/,�v�
�S��\AEi�
6G�����`�ߍ>7Ag6�����LP3Y4f��v�N�j�ܹוkR��`
Q�ʯ��:��-9ɼ �$:�m�SpZ��K �~���M��Y:8�*�p�j`�m����ݎ�ZOw��o�WG�~�{U�T���Of�CF�dڔ�;�wd%��#��Ȏ�w?�U=������n���s��q�6Ҫ�L\%�n�E�8D���^K��^�ݚyTG5���4ϟ�0?���́zDBF��۽5��ì��c�:���u��ޖ��ə�y<J���-�����خ����L�.����Y��ӧ����.���qՔ<��gЧdM���1�y�6(����S77~�ݏl��*]��{���7�]6����ho݌� �f�yE��y �h,��L�"�D���.B��4d�gx�u��а��ϹS����L��R�mV��]���h�0��=n~7ΰc����;���X�12��nz�����"�dS�;���ϓ��k�*"�j��]�7]�L�.=*A�����MN'�g����n�Ɵ����UO����tG���E�e�R�����;ַu��]_I��j��*���l�b�x�Kly���C���KT�n3|�ج�`{z����˪�lsW?I�D7�v3�i)�Th��ܦ;"��Ҷm�B۔f[F��}ܗR���w؛[���6Y��V�`��A��*�B�6$���˻���P��]P\R���-��e3r��ǵ��il�n��%)	��d��*��'�o����J�Yy>J�
�6�E�.��7l�v��z�Cgno7ZA��U�A�R,�����:7��Dǖ�Қ�U���S����EY�mFh�dP`�7�k�H�r�A��ŧǒ4��RwoI]�JWPԙxg5ٹ8��s����*a���#��ł�6o%��H�j�Ok�kӆ��"�b��a ��&Ӕ큷jC�F�-~\m��֞򞌛{i-Y���߹r';�/?t�� �0���zD>�w+�9�:7��;���w�L���K�ɥ�d��I�Nxp΅���/��Y
�:�m�r�&��t��":Fj�w[~H��h�������,*�UL�����(:�[Zk���O�)�bq�t^RTc���&���c0g�L���5=�2t��g�S��]�m�p��Ḷ[�Y{,|2>�Q����c$eÜ��j~�2r5�PS�7�콼��F����:y�΃L����W���5����͍\�Y�w�O�N��Y�tkyC�s�%��M�1Q�Pg�.�hj�ml�t�;u�ځ�on�1.[�ǼZst/��x�RP�E�Kb�g+tC���h��^v��.M�^>?��>og��<s����{�	s
��R,_F��K�R�̍㙋�Ϫ:p���C�Yc�'?��U�5�0���7>�r�D����L����=/>�\��)�"� -�m2��[�`Qd�TJ��"c�*oo3i�x��]S��3���F�
��9�yh�"U5�6�,�ȴ�+w��t4t����c�.�_O�o�$�:��AH���[ֶ�̤A�j}W�6"Y�Vo>��wrA�U�ؖ��^��8:��R��:��W��f����cO[G�Z�z�'׌�Y��Z��8`��.4g&C�wCeF�}Eﻡ�/�!)v.:�uU����3�<�4 �Mj�Zh�k@y������ ^\C��wd�ڷ���ӯ{�xy�3lw���t���4Ӗ�$�~��=
����<�ek��U��x3Fk`���bG8�L&������=Tʉa��Nǐ�W�/[[7�n��e���Hv1�������ײ�m��/۷+�녴H����S	E�z�Q�xz����%O*�����^˭���8�/H�V	���%m��V�Z�fu�1C�G^pNub�㋖�0e���<��ݹ1�f,6��qN�/fu�r>��R-�}���T�h�"��k�P<�C�Z�	���Q�o,c�G��/lGs=��jrKWaF5�Z�36Ŧ}�|�zgp�J��ݴ�Q|�䮮��n����������A̎��2��g��>�I����h=Lc(�h/���j�\��#�d��Ϯ:A�l�� �N�އff�P�/ow*��I�e�k��{2�r����{�`��ϔ�����V���D.q&򫳭��Z'1�n3���J ��y���Xy�HJݠr�M��9�$;<T��zZ�o<h�������U֔ov�RC$% [��:��Q����G!=�$�K_4z������8`TLbK+q�f
�(~�����T��ٻ�w����Ț��r�mR��y��ϗ(�� G����y�}�^�W������y��#�s`?S��l��r��22~ӧ�r��V=���@\c������D�z�,���6��B��we���!:7�fκ܅�m�8SL���J�+�_j���s�X%s��Y4�$�b\qsrG���a�s�PG���n�0��þ��8c˔'x;c����n�ζ�%�=��\�+��M��6S�&�85L�Ŋ	�����ܻ�%)x�������^~����.%GWT���V�\=�x�	�s�@���Ԭ
��݁(����#	��k����voq�w�燏�����W�jVŖ�N�S��-!���o9s�?��Q2����ε�:��۞���j�s��(=���Oq����N�Ԓ6+����p��vl�4õ�¶�˂�f����$*){�(=+���R�@����_��갢�/#�&�!����w�3	�"�"T���s(c��g���N{O �����tvv����\���!��o8��F3�V$r��	}+:��ʝф#t��)zrY�:1"q�g۝��/@a�#�a�ߨ���|+�h{��$�ӗƥ�Ϻ	w�3A�Ƚ�>z����]�JQk�Ƞ��uu8�ۜ���rQX{U}�ы�Д3�\DNgԙ-e���c~���Ļ��{Rlh�\O��Ui ���op�u7���AoAm�]��:��S�s �TuŚz0r�i��=�un]��q=���/RZ���㳴V�7��cuxtf"X�&L�%K��]����w��� �u���}�8n�r�$/�1T�/Yf]�<Bg=sH�6v��5������(PM�Kr��/+wm3�!���Xlhͳ�ʻ�|&���D��0P���L���ݷ\3nj�~��xo.�GU�:
b���q/	����k=�\,�.���f[3w�_�O��^��ؘj��w���pX���Tc (�[s4��]���K�c�=�A�0�4Gz��?ji��dqR��p4��a���E�_h��B�;;I}G�5_���pf0:���H��H���hK)d�|ww/�ު��k�#�w���w����ݕ�Zb�(�������M��^bAy-h���#:��-��Ʒ�NM�h4 �6zV�|�@�������i�7y�am�(A��}40�ө�f�'/�QaN3b�oj���;���yݿ���0�qi��y��bb�F�e�ƫ;Dm\��5F�i�J�u`�� V��34?z���m�"��U;�����vp]R�oq�t��Ӎ=���^�R���p"P�i�A[ǉ��N/W�,剳܎I�b�c�h��V�a�ȎgEQ&`ǻF��2g�u����=�l�nc�q���#8m�bl��H=o:��y�DZ������ۆ��vgv�:Ɏ�[w@�g]D�+^e�f��F��u��}O6� lNQ��E��*u�H��(���wC.�;��C�uG����eTL�]j��Q�-�e�U���l�\�M~%G��S �`���52嶝��%��fmgl�����h��cU�u.��%�Nr�妶k\���m+m��U9͡D�6�����R"�U"#o�*9���RӖ#�Nr�WY��rL�^���Fڭ�:B�e�-�V�v�qEX��U�(�D�����b�J���g)yKKN�u�-��X1rT��V��Z/�ID�
䢶֔mX���8�ȶ6��t�嵕�(-hʊ�kj�J��eU�ST���QX�ب֊�����%��T+u�*���b��k���W��\x�r�Ҋ���[-�iAkEJ�5�Z�A��+Tl��+W��br�]J�[U�b1���l�y�5��]G��J���D���Yy��88R�l��u-mj�EiRT��#��jUDNm�(�T����UZ��iXT�T�i�Q*}��}z�c��^p�v��ӽn+eY��IE歆�ĭ�ps� �����:��c��j�y�Z�|v~�޿<����ͪ���<��nSs�{��oL��ӳ:��ol�X���m��6�Y�ѝT��q�rk��y�E���F�3�0��M͓t���o���fzN��QL��V��}|�&�!M�m��Һ��J��Vm������P���&T����X7T4�k�5�`�Rd����V�&�2��QJ�7or)�P̾|�{o*��1���+u��OH�ȸ�iUve,�}5l-�^��/Lk���V9�5�ڽ����
�sf��k������x�4��[
}�� �y��+�s� ����'Z�g��|����^����]�MKf�s���n��dn��`��3�6�N�-y�o�!��j��9�"!��������\ge�+׎A'���q�hA�%�qηr�K>�S����3?\$�Er�@&�#�n���i�b5���'�P�8��G�_�MW�+�W��'���_/ Ėr��B��]s�}	��8&{�PQ����`"��uB~<	��2�Iw��	��MKpE���`O��t[��'�i��x��H䬾�0��p�١tn�9�:��M���}��,߇�yn�Ik����q���5��V^/���������% ��4ֲjUc�O�j�m
+\v[:��<���\�9�&����<�=-�f�U{ڳ�Qw�k��Xtm{�d��� j�.�X�*Z��GK\<D#=�H��Kt��ԥ�S�_P�=Y�U=GmV*w�l:ܹ�}Y�Z��mF5)���-���6����vjIjV��ª�ٷU��u�M9�7���5ߚ.)%Us�_�Zk�}&�Π�-�y�Q��}�׵�ݳX�v5��8ʥ��ɂ�E��o�Mw$m�t����g � �kj�C��N�Ǉ��To\e%%�Ɏ��hz��o7�Svb��F]��?	y��ѶGi�s��Ez��O���lŮ�=s"�0pʓ;UݝJ�*���q�Q+J��u�� fp-��y�m�`ڶ�(��e�󶆃�M %�_����<f�����v:���x{Ԃ:?V%B�7�z�s��0K��؂G�����XYF��}���1��+wsU[��L���LWY��{� �K�����,���z����c��W���͘��7��yi�8f>ǔ+�r�"%=�rF��W������"�ʵ?�UqI�1�wV_$�N�; p͏�SKe�@�;{ڟ����d\�ߨL���ww,Y���Ӓ7}K��У�y�O�7WD�y[KU��(�h��F�\-uz۫����=�o$���K��ǉd��"�[��`��#\10���!dH�}�e����er��Sۛ��r�e^�G�oQ�Ȉol�B;`�Q<��,\�*�� �Iѳ7c+�P�֛k����Bɤܥ���^Q[���j���s�at��k�R�*�m�v����k��h1��C�G�S��o�r;.<����;�I�&��d�xT퐣|J[@�����j��$L`��S5]�3{"NO`#�l���rO��{�t	P.0���[c�P%A5�6�6�t���9^�r�f���4Ro�wQ*&;	��r����=,2�k�R�����z��/���ً��Y����T{�a��إ����KcF���JK�2��3����L��Nc�5E0�VHkj�8���0�W�nM"gRb)�&�i��|��Ϋ��_d�0,��|W��X���Lw٥΢/9A���F�O��ւ���x<	w�����k�*�&�6i���s�u�v�}w*뛺%��^҂x�vM-�*�B���q<n�]9M�,�z�u�"����vƦ��T�W;n�:9�g�XK�RY����\ޟ;�;ρ�%3�_Q��,���w]J�9C�W)e�׺3$��@Ϩpx#]��>���v�P�WB;��-ݷ3��'����?���wftNr׋=yzk�t�D3��k�|�C�.��F����J��9�<�w2b�7��w�}l2S��&Ijh�{6�o52F`���o�x���Y��w���Z��G�x{g�b�9�?I��anwO�p��'S喅�)�r�ӗ�WC)�onu��E�K@$�hϹ�9���a�3�u�ML�lWm�����(�3���Y��ϧ�y��0k�����T�	�:�;e��������x��j�o���+Kr���뭕�QX����y�[��N��l��viw����h���2�o�.�nk��x�;����}vΊ�2��	6��[���֋�z���0��!٥	���a�K�UpYl� ��V�=��dԫ&?�V���|�7�	��j*w+��"��c7��lS���>�"�����;R�+#�j�;�tgn�\*�8��B�ՉW^�������D�K&Ӽ�kxϮ{0g׭����wS���gSA��N�Y�������j|�,r�(��tv) �NP)em��)K�L��5�5��+��i�;��Z.�N�Y�u��{��.'�����k�U��� �|�ec������n
t6�xt՗��Y����.���#�G+$����$�O����B�U\{^�M�S=�$���������s��P�4%�+�4TQc7Y5YF�f*�WV�V���L�;`�0*u�WrޅǼ�Z9�0�dԢ.v�wk�\v�ΛD�M��s���l�p�ߎ�@�#U)ף�.E_f�M���owv�j��NH�%|@��͑oO���'��赯@Pb�{.�1L1F��RT�U�{�6LU&5�K��\oWb�::հv��L����]�lAxxEc�}��5isl�+���c��A)���u2t�d´��������b�N�X��Wً�9�Q@nM*m�V�#�d�6��q�wK��D5L��Nw\�U���T��g����v�Öl��M����>�h1]�g�k;O2CGd`}�Sy�����f�`i�Y`�X��6�2ݝ�0���A��\��y���Q�"pV�ˁ�:ͤ�=!����M#{N�����8����"�z��d�wkQ"��1�Ԟ!Y�@*�u����a[Ka7��lW�p�^W�^���+<9:���j��w����R_ww�s����t��(t�nZ��X���=��Fk��qbz%̍M�|�Y�����ꩻ<yͩ��;���s<�	͍"��Myu�@�O���s����jS��Q�U�h�������q�^�!D�Z9<jn�v�W�[��v���5���y��o8B�o��5#w�\��Y>�)u{�,���׮�b�F���d��k]?�0�xq��w�0Y��O�d�G,�6�kp{D>k��t��M�M��Yݽ%�͌!�+�Տ��Ĉ���T}���9�!OS� +U�֞�\�Z���X9��S�^��t�Qk�Y��8�8c����d*���:��ղwwi9\�Uq�u���r�j��b�z��T|����5t��/�͂ҸN&c�uQ��3�/w*��Hk|�� B[ \����-C�3�𑋻ۍ���]z���M�6U]�yl�9�f��qޡ�-��m?Yvֶ��͜�ّ��Q�4f*� 
�J�I�����U�\����~�;�}[�AW�8/z�ŵ/3q��+��Ҿ���z�J�*��-��0hl���\@#��ثY�9���.�ƥ��n��)a����x߸=4v{	�T�5���o����R��t��k�����9���V
5����:��V�%>��;|�t,�ye�{>�"��}>�Y�����o}�8���'�����ݢ-]�b�̐�cq;��dg����
͋��Z��՚��p<�7,Ns�����Er�{��{R����v���2/��YX���":;9S���ɒݼ`5�\y��B�Ż4u��i��~Ά{��8���9��@y�|�����I7Z��{&�?s�M?��+[5�S�v�����n� ����yS¼ÞQVa����ۿlT��''#���Bf�Γ�V\6�6[@�V����x6��.�y�磚�F� +�c���Fer�B=�R�Wu�ئ�7:�\�5g�_H·$}�n������Q{wB������f�Hl�ֶ]�i�R6[�lU�n��]�;�h���0�&L�R5�Qd(��'�z�϶��(��B4�6�������lR�mI��]�S@�0B���{�+�Ū�lu�uz�ē�K2��>G��ʹ�����U��m�����z��1�����7S�Nm��'�E��^󼉼.�/7�7�/��z\�u6�zj�t7�������*ң�c�������R|�p�1O|U�-�>v��-U���	�,�����y�rv�]В���ϴ�`��90W����ѴMK�d>��i�e'��N������i�|�%^³�4��5$&�V*�X�Ni>��
�X��!oP���SK���T*K�Ӟ���zכ�/1�fy��ю���<�9�`�;��>��J�wzl�Dk��cZ7/����1H~hvI�:x���(�
������p/=�T�g�^$j��hن#�Guƹ�W0D�'�Zs$P�G�-r��ӨݭQ�15�K��-�?z�;�@��c��o`���2 ��{�v��u"��)�?:�b:���>�=�9��T��*ޗ��u���H߯,��s[]V�0}�z@�_Z00�i�z������<����� �ϸ�s��anw>#���3�f��Ӝ��V�?�&6�ϛ���/e��>s]���6t��2~5{��*�N��w��!�-֓�0�gl�8|�Z
��DR� ���7fn��>��v��x�5��B�fd=�f�'�ry�,W���,��׹X7��GF�q�ہ>����u1F������(&���3�n$�_�k{E�jr�FE��ֻ�>q�D�������;8ֿevo�k���Ã�%��]]�I��B��,�sj]�S.���Ơ�����ٳC*z�U{�p�����͞��ҲE&�8�h�ʠV<U��c�y�y�d�"�e{$�
F�?�í����V>c	$����T��r͔ ��8xfЛiӱra�H�����S)��sC�8$y!���o"�3n^ �����ߗ+ձZ� g�z�X�p�Ti�U|�����*�X��n9���JP��>|&��ngR�L��S6��K����JT��$���5Gxo�)]�wa��h�+40�����X;�k���q�g��|]��{���:I[9����~��f���ʜ�qMӏԣ6�5��l����6硤V��Zr��]�,��O�����˖̅gP�&�>s��θO��e���n�. f��Bk�[f"���r��s��������[��"*����v��/�����5�w���l�6�+W2>U�zo�4�w�Z�eG�9c+����y/S�����$0�G�.=^ƒ�gOb��<�9�D)��7~�	�49�}5�w~Zu�S���{6��K�{��M]�M;�$F��-3��,n�o���{"�Z��(����P��v+��8�1�z,%dա��UW����T(��W���=���.��Vo�W�g��yB \�:�TNhy����G[�hDE��X&El1�a}x�N�����99�}����?����V�~A $��$	!!'�OS�F�2C�Y ��B��N���&�D�H����"$BD�H�	 H�I#$b1 ��a	$ $d����H	�wb!����H 	I$H� $��'t�� �� 0'IIH� ZN� I[  ԛ )+@ 5&� %� &Ԛ H��	H �! 2B ��@�  �� 	H �� VK@!$"B@0�"B $`@�#  H� 	$�!  � "I0 �� ��I"D� ��I"FI$� � $@ 2I$H�I"D� �  H� 0$H�D�H�BD�H���H�	2" 1��d"FI�$H�"D$H���"$d"$BD�H�d�#	2H��D�H����#!!"F@?�ݟڇ}�N�����d��"�BH�������y����?ؿ�����?������_��oܟ����q I'�������	'�=Ą $�?�?Xx!��C�ϩ�����������RÐ/��?������C� ��?0�M��$d 	H� � � I$��2I$D d�H�� F  ȒI"F@ B0 �  �@$` 	$� � F  ��I#$ B$ H2 $I$�$�����$�D�� 1� $	 B��
4�����d� I (EA@ ��=�~���o��
?��� �g��~� $�?u���u�D>��;??��O�����}� $����~�����$ $��! 	$�?��a���!$�/�G�d� �N�@���!C���
����؛�y8� I#�~����?�! 	$��|����}~���?z�?@<�����%	 	$����JB I�������~@4;��C����{��|�|���u! 	$�;�'�|�XP��zC�z����I��!O̜�P�u�H@�����>�O���`~���d�Mf@(����f�A@��̟\��|�}*ROmBB�)
BU�D�T��� J�
�)��$����EIEH$P�H���TH�������))�i��T���R-����%	#�LT�R�*�[jM4[2h�5��)1h�)El�j�F��
R��ͥQ!#O�aH��*T(���H���jUYe(P�*%� �� �+mU��h�Eli*H-��
5�R� �BJHUQPI��m��el�  ܜW���Vi�	]ۍ]�h��l���]gv3T��S�.��ilm�V���v�n�m4�vݪpە�iƻ
�U��Ķ8�]�j���1kM��kbV�H�e$�k<   `�B�
�=ݞ�B�@ �=����Р���u��� P]�y�4���v�(�nvʮ�ܚ�]Gw]ۛv�w\��u��t�jۚi$Λ���u]�V�N��VmPU6�$4�   ���q�U�l��j]ћk�p�-��F�ҳgk]���ʛ�n9'v6շn��K��J��[G-nt���ݧt�F�ݝn���7)n��Ww*t�Y�TT�Z5H-�[^   �e�ݭ���4�꒷f���WT��.�ݦM���R���Z�n)S���Z�ݵ��mβ�mMN�u��\P4(��8ꪶ���ơel�*�UEk��T�  f��O��r����b���:��p�ږq�S��h�i��F�n���(WMi�X(j��Ltt�;��۵)�wT%֦�V�ETmmZ�B�x  �z:wLUGvsU�(-:���r�uP����U]��siQղ����1� 7N��5mF�J��N��[��$6�ص(�J�J��^  e�Y1����6��۔�*���.���e]ӗ4v��r�iP�N�7+l1؍-� ��\ 5@mS  YR�**.�+`ƌB�<  מ� `  wp�  0� � ���  � � �Ӏ  ۶� �m �X6 �;�U*�e)��R�
  ��  n:� �NҬ  �  (M;p: &�p 
��  
\� ��@ 
����@7m6� TM���+CTx  ��t �0  �  uӝ� �� N��c� ��@ u� :�� 4Wn�@t<���)P  E=�	)*D� �U?�4�=  S�A)J@  S�&4�*Q�@#	4�U"  be�f�A���4�i��M��)H`Օ�~R��銽n���,�nL_����I<����$I;��$����IO�H�~�$�	"�BC��Y&I��@R�x1*C+�1� �Y���Hd��;��*F����Y���%6Ñ�(���*ݜI��h�^���jRR˹Yb��9��/%��jM�e�ěܣ��M�Ѽ�,@�ʬA��Ȥ������%��Q7)[Y�Tm�iU�6��ٗ��JJh��w��J1����0��Z�qF<'*f5+�[Z��r��6�iǹ�>��V��6��	Z@�*A!R����/]l�7h�
��
�M�v���TDhOl�^B��f��C/,I�����3�V��gI�2'zű~�5�v�v��cU*I���xU�(���Ƨ�2`f��/^X.�e ٭��̫�􅘛qP�)Lј�E��)��)I�t�WĔ����p֕��6��ޠs0�Շ��V�ۧA�kX�Y2�(�d]�p3�k��j[Y#�2��h�t=i������f�ϳ!�`m݃�6�ہAe�Ɣ6����j��)M65�A�t���c��V]�6�uu�ҵ2���ɠW��	
�b��9��u�*(�Xa�P������z��0�;[��e�E`T&��f$[edbe%��J��GVWz�&� �R���O2�h��Kg>��#�kkf���p�fiE|cɓV�ڀ\t�NP�ӎʡ4��ɍ���$������ja[���`�I�@��$hB�sU�ְs"�`,{��t����T�B�nՕn�6��'��<��������|��̮�F�j\9�tmݺ-0�ѽi�� ��ʍ�[t[�RM��Tx̪e�e��=(&��h(%��%�z�:�N��f�Ʋ��G
�QÇ!%h��j��$T��#��Y����@�ف:�z\{anh��EG�L�M,���cJ�@� T��x3Z���>B����eOp��QB��#,'��4�ݖ>������Çe�պ�+�nۊ�� ��oJ�E-Q��щ��&���C)���?d�p6�EYX@�M�	��miTpJ���y����$�#�S�ǁ�ʕu+F3(@�ڼ�R�)��h=��ne]1�)����,�1�Z���,��ҭOi8\
�޻��L�4UЩB�����p�X�r�0��G�v؎��j�T^�n�Ʀ)��ZA//7X��fQ�J�f�1YR^I/c����F$;x�zʱ5:�M1�j�4���-̔���IˋX�ע�ͭt�ʖ��4U�.ɤs~��`UIo*�[�Z��ȱ��#��i6��,1�-Cxr��pޗhn�rb�!�t�%�[p�F���{���oD��R�-4匍P���꩛x�$C08��w�*nl�eDAeMu%�y�t	n�,Y��w%1Bx�.ɘ�M�t���c�Nniԙ;���`<�fV�h��gq:T^��R���%�fTB�XA�j�[�;�R�e�%I*X���d��t��(�ȖEu��U�%pڳ����@kM<Sou۴ ��PY,cԷ��f��j�2�]5)��7��,�/�sU(�z�e�0�oh{R�C-n���z��Q���艝����,ֻ��[�F�M�I�&�
5�����SY�`ǂ�<ZP8��S�vpf�v����B�U�9iU��nȄ5yJb�sV�LJ<�-��e��Vh�ZpYWx%����c"�	�������ǅ+:�D��	,�b�U7�G>�KI�lA��e3F�"�-��ua��ɬ�&
�1]�n�bj�E�\�Գ5)��f�F�+)F�Kl��t0�Tx��;��r�����9���Z��e=v���Q��E2�MѤR���[��mHCyr�o%�����z/.��b�a=�{H�VZKhcn�t܆��A1��#L�0�7HR��"ˀ���۩,�dj��8�e:�M�̑�HȨ���T�O;P��j��!tl� ���x���������U �0�Z�OsU�1�@�O2񤡫�2a�g7r�͙nbBZ��щ�ˢe$�h�X���y�L�n�yon0�M�T�x�-�L��@
xt1�N6�=Ϯ͚����q_ٕ�a�E�#]<�Yi�sRY�s%9�6=b3`S�@�;�f�A]	���,h˼*���$�6M!���z�}4$0h�wmQ��n���Ի���q��Z�?f,�H"��l�2�����ح�z��N����gö�&,ۧ�������EG i�K9��^nU����J��1�� H��Q�Gg>�N��U��1�p�*�G*l���{4)�2(���
��g��CM1��ʈ�b�ʍe�*WN��j����^mԼ�/$D�Ѵa4� om�CS�z�;�#zf�rd�
U�)��������$Szx���7-mܠ�����a�2�xF��hfe�]�l�;/q@U�\��Fwm��&��X�EErmභD�W���n:vu��v�k��vi62R��@ǮV���{�jV"�+N֩b��-��"��[��&��5�nZ�6���kAlX���%2L�J��n�WuFhSkh��u��	�*:�YeK
��k��J������+6�J�uY���Q�9M����蔯0�v�V52L�
ڬ�*��!���d�u���0ˤ�����u�V�#S[���𢮳,��z�<R�We�IOi8��� &l��)-�1�X)[j1S��Q���V�5���D` -����df��l+��y��-u�"��e+�\�z�^�[e����V��,A�jon�#ڐ�J�k,�e�љ������R�&��wW���3[�mS�%�m� ��7Nեuw�x�����q�ɨ�� =�В�g�e�Kl7������vĶv�$����.�Q�1��%�kQ^���m�*�f�T"��J6�c�/f�M�����<�M�-1ZC���8�Yf�a�R��}D���j(.�O�Ӭ�X�m+B)��H��� Av�ܴ�K
�[N�� ��[3T�Vj6˶ͪ���n��5���&�ZXxo:&c/��n+�m��	z�.�Dl
�h��b8���`��L�+E$�i�i���hs\�&��V�v���1R���[�����K�f�<�����Ϧ�IE���<�5C
��1�Dj��v��m�-�f�j��������1�@�\�X�C[��@�QLC/E�s)�*���]*�wz���eh@�&�x�dP�)��،���kjd�!�^7f��h�a5�j�Pj�l'%櫨���Yz�+;SkmkE"��Ԑ�-�I�V�#�U��y���T�(����Zۭ��FiZ��NQ2��n���̍˔�ٹȵ��Rm(�Gofh"�B�G0�+`\�u��|���M���E邒H��7ou���um])}���V��HG�C05��;iq{�D2k2�~�&Fɸ������u������YMǔ+.��;�P BYЌ����
�wI��\*`��;x�h���W{KZ�M��%m�{��6��̺�퉴ɧv/�o�]W:����;@U� >�(͍܂��Un�Z�U-!{�om+�6��{L�U��w(3�siM]M�j��բ¬�I��-k��t�TJ�LQ�^�>��b��-Gy��2'��FVf�C)^*��)=Á�U���#3c�
#)�
���0Ҥ�t�eMh�w+]�����J�Zf��RI��	�ώ�J oD�j�,Vw�k�˷��yc��U8wQGZl���X)��m�*m��N���m"�!��Da�x�J��2�t�H�,t� 7�t��wLd�y��
[tm�1(hʁ�i��SM���3U7��y�yL+��Ee�)q��6�u���/�HQ<B�[�V`�!��<�N owN%6����(�֝+�z�b6�K��٤ֽ��ek�Ƒe��� ���yjbD�7�b��e�����ݸ&�3��Ѳ��BU��T��̨�0m,��A�*�G-xB�6,N���)(-�!��nN=�,;O�<�KnE1D7���:!�X+�+ݝ�m��{�[ ��1�V����b ʚ�{�131Ҳ�ڭ�t.�@8�Z
�ijur���UM0��T"U�m%�-F��֋�M���f&^d�U5z�XR*�WX�ræ�>��IP�Xl�
����R�vb��h୚o]�gu�
���Bm�-٧�1 ��c\���J�E����MH���-���j��r�ɺ�r�#-�'��SK��y	:	"��{��и�u�i��M5lа]�jcA���=-�Hur���:5��7u�p�t\���+l3ɴe�0\ͣ2b��y[5P;�ZH2Z�`��{e�XͭH;i`&��� �ןm	�ڈG�+��A	��n-x�i���۬�u���P5��IJ�94��L���;����@^����wM�ȗ��S[5l�[�)󙠀�b���
"��0J{Z��$�J��"��8�Թ-���#hBT�a$���g�ۘ��6�ڄ�쨱:5��Vm7��h7Xd��ɷn�B��e�����*8ˠ\p�z���R��J���8v�6T#@�\�P�^ӹd��XGY��ZRVD�@:�R�hѕ��ю�Ҭ_2�����u�"����jlȮ�r�Zn��wv���9R酊�1[c+482��P�M�by.�4�V�r|�f��n�����ޜN�t5ʂ<W��)�l���H)J�,�Z�X/*�8q�mn��D�3i��*��)KmA7`���m��E��!�G�`Fl�4�cY���]��yu�Kmf��賙j�xY�QC.&��m}{���㣫��Ɋ���{��]�F�UyJ��es@�nb[xp�Z��%f+O3��A�ll��B�ci�h��>�B��.��P�v-W��;��E��4r�nZˁ�.�]g6vj
(^ҳWn���f���cb����m;6U8�����ȥ9��&ލ�.�y�ڥqfZA-'�Rgض���Z`�kd��-Z5X��^�����H.8�:�%F7)m].��ˇt�&���%!2�[�Il��ت�v�8+EF�Rue��������1�j�곮����f��a%DwA�s	�1���@V�;NU �,� P7�{��K)a�B�>���P"Lm��I�X%�B��D�����H�g��z]�5�ņғl]�QuJ���] �ƥ�C�Y�$Y8kr��HV�,b� ۺ�������9RQ�0],e�hG�J#%�xE������}���x��:�,M��7aʴ W��s�NlmY0��蚹�a�rBsl3Sk"�{;����I�q]<�޽d��)��uD|���$V5*�rj�BXZ�f��j��,�����W(g%*@�f�2��Z4Ǻ��u��wh��ʢB�(�!���"��^@r��ǻ@AS/4* �y���gM\�,i��L�<��bSj��uŐ/m��6��4u�#F
{��i���h'�� &ަ����BhdY�T�+EAR�aS^�Z��4r�PVm+ssq��H�҅�4��t3!�M�퉭V̈́��kkki̬�m��$
V� �5o�Î����[�c�2`�"ù�(.��E��Z%й/���% �!6(f�MR[�Q��Q�M�Z�^�Rm֥K&%s5�6����8:&��l���c]EN͋jHa +^\����økfR
f���8�˺d����HŜq�(�ձa�Z�i�c����������ʒ�O+�oH�a˦`�t�'�x�Vh��ˢQS
1���V�;��W��K%��%ތ���vPӌ%Hj���`DǶF&������cq,WygLB�P���M��ӹ���7�VSD[�ı�wp�h�E��\��Q�`詯vXݻ��Yra�E�@<Ɲ��	aL��<�;��b[47u�SCrĽ6� xÚ-���	����9���-c�zD�.�l��B.��^�ښ�TU�eIWJ�T��v�5���VK��9�I*�c�]���R&G��Q2��)�3������,��&�Q3.\@�Q��T�f-��E�X�ˎ�śL
�v���� ��LM[�fP�߅�R�����������m	oR�엫�*?@��&�Mt���j�j��Hl&��v��)�H�8m�6��ya�ubV5j�)���-d1j�B�e�{͎�D�8�땬�pPw�%�-u��5�p:�FLJn�v��?Z"�5�gڎ.yWZ�u8���^��a�e	XCQcV�ފ����,O�5�2��QȢ%*��hN����D�R[[�2�e|m��i����UT�Gu�7H�M+��&*�lm��X�nH�&=.G�&4L�lj�%#7
�ۑVֻU���/#���]�Z'p�,b�:'v�!w)���t]n�
}6L{!�*�,�F�6�[�aS�0��1BjJ�;�]d��$�h?`F�{P��T���+�T0���O[�XpcWr�8"�2�$n���nm�ͱ�ܼn��j/;i�Z�2�h������YSFRw�MJ���C6���z��ki]7�L̈��2�*��LU�/D]�7u�x�-m����v����5)	9(�o/51d�DKv��a[[��K��ǻrJ�w(X��)-5*��
�A�)rLm�@ŜI�2���Pmm5BӆV1*��+lkn ,���8�Y��`�@e���
�nD�/�B֪�4�:/r�:��T�Y%�vM��X\u���N��)V:�cn;Up2��JU�˗\A�L��I��V���ӹS�)�o�5ٖu �4pf2�m��I�+j�ꥏEoV�kHL���:	t�����y��X�eL�m�U�K��}f}���O1N��'�N�b��\��=oR��p��կ'qC�� �ʯO<��Jy�]�{֮)g��'u�ޗ�6��+ TzJ�w#�x2�a:���Y5@T��7\s3����J�V�ܶ��O��]90��:���&��m,��)D�ϻ^s{-�}��v����zQ���<�����o"򙛕�.����Z����S�+2�;uʋ��*���pY�h�ފ_Mn,\R�V��սXCn�gS)�O7}gh�7�}[R�kٷ)-�l���%��S{���`��m���\,?�����`stq���ob�U�mů�i�+f7{.T9�ӟp���Ql^�9�w�))�_J�M�W��hN4��ΎË2��[32g�8�/6 V3���5isY���,����~�]ۗ�Ho,AYB�z�	�����Iʋ{<��A��:�\W�{��eev�y{\A��Q�J�}�Y�e^���(��h�D��O�wk���!��͌Qm<-�&쾾kb��QU��N�B�{����N�hLfuk1�����ڴ��J��V^�̡vy<3K_tv���9��e��Wi{�i�0͗Y2r���(S��ݲ�Y�� v��؋d��c���Jgc�s�N�R	�&�Ok]���h�K����I�:Y���.�v�'BO���K�����$~��
����mO�p�P�W���,'qG�����z;���ۏo.�գ[l��h�x6�&@���)Ҿ桖�t�p�h����&�h�ñ��^]��Q�[зw����i1fHբ�}xa�Tﻵ��]��oS�*���B)��r�YR�����EֺOW@�;"'�I���ւ��m__RщwnЦ����l
�۱],b�X�d��+TH��^־�;����X���0vT<��=� ��Z���N�j����f���˘�{(�\jS
pQoQa��?�˂e=��������N^��t�m�ݩa�	B�l��UR����/c�ţ�+�ZJ�zM�ﶒg���u;��wڦ��������W2{p��%�&۶L�������:�%���B5*����au����>��
� M�"�ځ����Ѿ��˃��R2#x��<»��Š�z���.]�݉�̳��"]v�I׊���O`�����"�Q̼��m��,��~论Y}5mL��S�vl�s5r�� �׷�x�C������淬���P�W����'�s�^q�|����݃�o]��e�	�;L��LѠ�"{-���%�6�l�1�!�WJ�J���]���r��co!��9$�5��L����'	��4dIѡs5�,�k������Z]XpW)�λ�G�'�gt�1�j�g�{�uaHWU���u%zup���3J���}��GV��ۮ�\$�>�)(�]�W��no?!��1����{���r
���wQ�l!�Ǹ�e\hbi��(Z6�]����Y�^�;�.+1V�p}M,ϲ|�n.�l%3�+n�!���p��r��!�F��S%'MuV/7jnJ�P3q�x����k��d	��k+��hT���_�>̊X�:����Wy�����c���[�ٻD�.�]�]�Ӳ��Wh
7�>�][6��ԫ��0ި�f�������>[�3�4x�]n]6^�6B�@-�cw����!�չ|���jR%�v�%N���ή�ҵb�3]8$�6�AD��l%�r���^*u�qw�eq˓t㐚u�;WfQ*���w��� �)���EWx�7�@��j4Uɳ��h=L�Ї�.����o���e�� ���W��s��Y10�L"Wh�i�T�h�+���o��<�=h�՚����Uu��ax��x���q,U�����oa<�/�5e���XgČ�f�w�7Ya�� f�떰T�����Ԯ�&'�@�x���U�v#�ȷ)�ך1� �k�EM��	w%�Ѭ38St 62��.�,�e�V�Œ�`������v�]ﱘ�r��͹{\�re^�JZ�a��X��p}[#���B7�jN�̜��6�9��a�v�0a:S{�V I�n��r��S:8!�f,T5d��s
�k�Vv����)n�uϴ7����9	�]X1�l���*�O�t�em�a�`�N�[.~dT�9f�$Nʱ�|�Pi�jN@d��j0���8�΃�QYrp,��[/�yz�V`߳��i��2� R�z�7�;�)֒�,�VӬ}{;��C�@�N�7f�L;&}���Hj��%���ab��{1��7%I �p�S�7��4�[�oZ:����9��E`fk�_6%�P�9��d4)3I,��t@� yt�%9o.���E!!��j�Æf� ��tKM�w�wpG�ц�v�Ncn^����!����Dl��1E=u�or�N�Aft�H�Ӈ�i���Y��.��e4 ?t0f����5u�����D�rEN��㬢%mg]�'�9���gL֯��Ų��T���,٬-���q���&��Ɯ�����[Vyu6$�za5���:�{n�����K3n�ؼ@��	 ���Y��g*(���^������t�T:)^/�^X4D�{}��bȞV(tأ0�n[qG�N�l�/�Ͱ�m�e�ô�V�ђC(֮*�J�sJ�Ÿ�|:����R���&�cO�&�&�b�B��^�Ǌ�#W1ӗ�v��2�����e��U_r@œl�Z=��ʹN�����u[��7�:;��Ls�&#�4�f�桔T{z�=����]H4��Fg�M�)ǁ�F^TwZ~.�'�����(�CA��-]m��ۖ�z�#�D�7�n�:+<e3Na�\�II�pEhW!��1�u��O9.�J�=�]���ea�B�������v|�*Y��iNd�)�MH�;���^)QY�����2e=�9,�(s���xa��0�����$u�Z�m��bԹ�j�$�����N��u�ۈ�R�ֻ=N�7)Wr
��� Obt�*�����ݻ��r�J��B��{xZ�������O,$�5i��ٮO4�R�x�6k��|*��Sg�u���4}�#pV��j�+0Qw|`�UǏ!�d��{�P%�.�`g��=�p9X�t�O��f��b�͗��rL����
8`B�8��n�����fkq䡇C��v[�@�YY��I��r�כ�;5����CH������ʽ�n�vV��<��=�T���.{p��b��\� ��*���_qJIM����٥��R�v=�S�7(�f�΂'Tz^Q3��f#�5,��e�4!�M�ͽ�,1V�ƍv��dP��}�Ų��(c��Gd�ʠ�ƶTI�GJô�46�r��ks{��G���R�2�G��(rP�m�����Cq�b3l#PZ�}�1Һfc��Ь�jFZ�H�����s������.��I�̖U�Uvҭى�e�����T�R�\ft�U��F���@X�kj�	5܃��VSfp�a��k���*�����&ܻ�B�� ���2�Id���۸����.���j��74�c��T;vT�V�H���AH��^�H��2]d����u#�I�pIwۈh���Z�m*c��œ�>���}/m:�3�A%L�s��r����Kc�MJ����Kl5��ۙg"��w��OY	��m��xx���x�U��u�&�ҵ%��n�whR�y���k ��}�ƎeK����SRn�r3�^Pa�T0k:�8�V��?V;'BWᴁ7��b�
�<���>�mýۻ��'f�.KڟZ�rՅ���R� v�`��e��8�N͒�Z�S�,%p �n�'dm�*�w�	6��O�`U��4�׹���.���S����{�h�����[��v������x�l�_-��x�܈d��t�ǒ�n���ƃi��Z �{���chES�^8�Y;ƭ�cǔc_K�[�tXV&��������(g"B�8Sv;٘�m2C|g�ۼ��.ͭ�e�!.��;_&����r�8@7j�+�[�7e&�+X�ҒSFXw]3]�8^�,������{2����q9��ڱ��'o�R�¢����&�*��F�A�Ew!2���i�W7S�Bg����X��"fx���Ɍ��5�eڸFJ�F��+z,�M��A���H	�	M\'nE�^I�A�-``�|�yu��8��&��O_D��>�2N�b�W��Z9����sn����9�{
U�1Cm��$���szt��v�ڒ�v�k]�Srԭ�OfH�սW�\�z�m�b�<��2��dg�-�P�v�B�WuwMd�*�+�n$�Es;FJ�j6�Rż��U����l�#�<��q(�'�:ћ�}ʅ[��You�J�C�c�\_:�F>$�m.��^�G/�!���{ho�{)��W^��a��lh���]�V�V��6"/�X�fF1�3M7����҃�X��ruf�Lqm]���T��xD$j�[�7fE<�ݬv��5�`��YA�Ф�V���FU�Tz7|Un�۬�B\�#1�?]m���,ͣ�Q�9Y��)���p�`���f�1*�93m歆�}/B9gJ�@�9�ST-����hP:9=\��h5�}�;	�ݹ��Ȼ���@"�f��ZF���E��Lp'���I¤$��W�U�å4��;����f*#̎�D�cH��]fXg8�[e_Z]�D�l���n;������4��M�z[�᪤	��y��M,�����g3x����B��V�̩�!#d�G��d]b�a�N�w*�U��Ǔ{u0��<){Y��P�J�C��`���w 	CR�u��:���7IH��K��T<0�G����G�E�"5�K�Q-&��8���v�!x�ǊM7MpUۤ��Hh�9��ũV�7(U�*��9�uu#�^ɍ���:�HWAr��K�5�=��9�v�M\����M���V���v�uV��ö8l_�/X˗ׂ�P�FAwR�{�@pWw۫�;)gpN!�!3S�wTz��RV�f��*놗x��c��s.L]�m��ms|��Td�+�6mo9-�����y�SQ�B�&l®�#H)u�΂�<��U��k�y�՗;̌E)�VY��*��*��ѽ�ګ�F9��^�6���*U�CjݵZ��{���=Sb�t�U��>�q���R�� q��e��Pb����9�Z�ҧ)�ۆ�CV{.��8�Ԇ����ck^f�]�T Jk���������і�[-y/�|���0Y�U��B��[/�:�s&�3iK0w^@�m3�d]0]���<͕{[��} o1ϕoP��;����C��eG�Ώ�l÷��Rk ��V�#*w߮oc�7�s���m��K[��T�(<NM�m�M�;�aYS>�
�=a�rl�L�oZ���Z�[��[�����妒����{r
��蜾���(��;^b��9/��.���I��v�y���p[j�ҪwCxd#O3FWM��lW�9�R툟'��unG��Cg��5�l��Md���9)һ�_u��y��D6Ŭ��k��6�ԙ�Z񫰸_vH���ɂ����
��ڐ＜P�Q[~^�
ӛ��,�%��Zk.˔��s��[5:�h�+k�֣䬽����!�ꗤ*㝑ȱ��kn��  Q��t�eȻ%�nvPǭ�Ǻ�5Z�s��[)l8���.`��*�JV5+�ً�0�Ӥ�4���Ã�1y{����g��f�2]�[EZXj���Hn����0�X�gm2vr(o�YK��l��s��#v}�mL;�Ĭm+A�[u�ڬ��/^&;bMݚР�ѩ*�u�myrpb��c�����_qI]\�׻�Vx[|7*��l	֊ã����^�`U�E���`�褄؎�RU^��n'fs�6r�v�Ʈa��Qk�3b���\@�Q���P�&rھ�d��ߔ�s*;�5����3�p�4�6S=;��mq�6�w�"��!]L�e^i@,rh�����/{Q�{-[:�-��hb��oۢz]ijz�q�j��G}y�ɝ�K��9����{,P�Ց�;nn�U�3��Η�Jj��2��y�b鰣WpWb�?<Y�10'[�oJ[�%��yx���o�Fi�x�# �㱗n��8k�wV=�`0]m6 .Z⺥`�J��3en�)�Wm��Y��Jk<�o\�{w���x",#ם�W%��E�+B�	+/�ǩ�a�6��=�kfv5Ē��P��U(f.=�n�9jՄ��3s:H���3��:V掣(E�ʕݝ����2֢��r���:���Ni`��s�%;Z�=��	3�w������^h�\�=�u�����/����\�ֵٷa�n��i��jdOֺ��}]�Qu��B����J\ox�3���+�L���(�3�Dʷ&��T٨N��L�$臷��"�]�������ˁ�Q�I5�Q��zX�+�f�QSգi-������j,K��6��a�@�Ƿ�id��RvN�����U�BQ�W�i(�t��1���p��b>�,�����m�=qɷRNrC��uzơFP�WB�9���l�7	s3[��ub�����,�:b,��6��'9��K����@VN�z>����s�s�3�n:�]t2�]����*��{�&\��/w�e����J�C��47}jKn�a��2Ly�2l��d�f9V�7|yp���utSs)�8����`%�L�M�)Q�z�0��W�	I!!�@�$�kλ�_h�-�:޹`lƘI��aVg�A2����|w�k���:h�}��u�jҠ�W��gS4�iS4�^Q{s���:�X�<)����a*��˥m�`,���J�fɣMKz wkOf����LX�E˖���[��<��8�M�+��;�!h��c1�,9��K�o�ήP��X�N���V���tu"|5�SY�����He�V��������5
ऀY����5s���U�U��9m�ňzm��@�u���	M:���:�Z��"J�Z[���5̋��A�M�+con�N�pI�֓�o/⫝0�j���U���/jIP���3�Ǻ�q�2��a�s3��2�Q��B���9�'v0���(�e�;y}rjj-\��}|��Y�I.Y\���Roh���uVz/R�"�c�`̺W���Őn�6�`=C�ݹB_����X�GI�����W�c@�N�%���s'+�QV�PH�=��lVҕ�m�>��[|XGm9YW�`s5�K��jV����K�lV��'oaj�&�NӢ1h�8��.��ȶ�%�]h+V�NG�c���ص�Y���1k	ˣW�̃�e�H$���(oKx�۾���ۂ�D^�zf[��ڹ�4k&k�.H�ی�V����U���u�j̈ul@.��;S�ʾ�xd��40��0kw�P�u:Nr�+ �!��)I�ar>k9Д�,q@=I�Y;fX�mN�\aa�YX+p�|KO�)�fڱ���^����r}L�
�l��c�u7���(+�9ع�i�z����#"��qS�فE��6]�Ŧ4��	�����54�����|�sU�PD�j?1ػ��z��E��ݜ���.�Tq����u:U�{���U��݈w.�PO`�wR	+�z%�k��0<���yR,�le+��T^<�S*�۹'b�/��Q�確w�|�-��՛D𘵓0���GK��j�qWHr�.ۚd�*շv�Y�|c��*G�v�AF�C��C�.]r͂@Z��-ך��j0�z4�@԰�&;V�q�z�����[���]���[w%8^"�b��t�%+��
�n�����Z$�I���gm
@:?b���U�I9��mP-�)�����v`9��*�T;�z����؛s]v�,����ڈ�bv�yYO����]V��4(%/ ��sF����p����9c3gQhƲWy�ؖ��U9��3`��}>�ݨ��)��"��Π�Y�Y��Ȉĳ0W(���;z��XE�Re����kx��x�i[�ݚ
�����7,�u�9;�[��Ixl`-�`�ã0A�-�Ů�:<�&�� ��+����Z*	:rP�B��9���Ԣ�	{s�I�oyн��
ƥ�|���lf}�¥V�u.-�u��)0}ԯ#q+7ZW-�Y��y�!���*��E��ܖ�BV���vˆ���Pμ*�G����]�o�ǗL�5jP����WC]�栮���_`�N��c�7��D�`>+��d��3:���V_S�b@nM%%��'֩Wf���E)�ۡAJ�Eɭ��[{j���������w��W��E`� �����]�m�x���(V��JS�h��㏆i�6�c�������T��g����t���5��,�������ݥ}�جU�m*��bN]����oN�@��V�gDkS٭U���I�[Q���YJi�`��v�^�!9��a)�7��v�Z8mB�"�@���g�7R���2�YtcR!�"Ͳ��R�z��ީ���Dd�\m��l��R�r\�3�|�u�.�C�ޱ[��3�C��f�f�ƪ�"�s�5,�D��D���[��Fm���hUs.�wa�.�ڧؔ�)��Q�����s�gV[Ƶ���u�:�����dק��]@�u r������y���97h^�ek�k�M��۱D�K9M5�	�b�,�-pw��7�KS)��e^�n�`�=ʲ�B@,�UI�/>�.������S��/��\�~xŘV�Y%���	��u`�񬩑-nǩ�)jW��JD�9�,SZ�v�J<(\ц��^��
_,o��R�^�U�b��[jN��̬)I��j"+��3w�s��o�be�"I:i�J�����+����̺]��^ۙcj
l����ue۝{��И̼z�6n��-M^ҁ+\�ޞ}ڞt��}R�:�t�}R������s
V�70p��Æ�a:��T�" nA��4�ܜ(��z�a�>�ͻ�X�[���WwQ|Ѡ�5wO2�h�<�a6]+z��o(+r�
����A����7*��|.��;,������Y.f_Ȫ�|oZյñ�S��G]d��b<�hV~,$�#\3����<n�_��OME-�t�`ŋ�����8����	���Z7t���_o]� (3��ܕ]8e�kK��ur���ʾ]�HH�VVCm��ڰ�6���Wuͅ-�+��H��q�ygS�W���{�m�.[&�HFͶ%A�vI�Q����Dkw���L���4�wg�׸B0Ye��p��GQ���9��� �Kq�E�w���~��H�4���Z �3��$k#��aW<P��7��<��Օ��m��uV#lK+���Z�k��\b�1��:TZ���6���շ�GVa�]IV�ŗϝ��7y��4nLgU���syd�P�i�v��[\�Ts$e�!���X�9�׹P�{��x�v��i,La�B��i{&e��C��QҭzU��Ԁ[�C{DH�&�[z�H��0����&�85�Yi>Q�M�v���u�0���6���vI�<�!�p�A�ZU�0��R�y�p� �l���Gb���<n显	V��@<��=ܥw�f�E#�-{Ҭ�֬�'���)��*Ǿz��m`Vz�W�)0���3�r!o,\��2�X2
�v��ƐT\�;�%��������{u�Q^��w��{���s���KuX��`)i�MYM�p\Y�d)mKh�*�O��.�^F�H��7����ec9���� �h�����ɮ4#��y'We�2��4��=Y����gU�r&����*���S���_��}(K����㕱���WY��
ܾ�\w���q�ǟ���F�r�8�N�>[+��n�n����D�gZ��D*���gJ|��q]�M�Ԗ٣٪�ӕ�jG�RK����Mϋ���S$�kM�l����	j�ƕ+VA�&*)�('"C�@m��Z��7s�R0�
\�UӰ~��ǐ�8�8�ܒ�Y�ub2���u��\#�S�;C#�s�
�&�.����'�S/y�fij�%��R���9òc+�i��]֩]W�j�ԩ��:�8']���݊N�I�f$5��dCgM��^��4Dti;��'\|�b���f���7����u�u��!�z.!��{v����l.�2���L #sp�a3tB�r��w�*�(��.�syCkq�]731�6U����خ֏C��\��x4m�]o�憹�i8.������%8ͳL�J��5Y��$2Rӌ�������F���pe�f6U=���<7�4��_G����<h��� >!�՜�������a�\Lε�&�"eʣ�l|:t�h7�J=/+�=n�ˈ��2p�����͉�[���_Pe�����G�m�ƞ2E䡙6�5ږd�[��A�����+À^X�l���	�YO�/]�p�l��}�0��|���v45�猀���a�Ԩ�9�����؈�:�����F�J[�E��4��=�*XB��m�� H��<D���P�T͡4�Uhb8�<:�1�^�-
�ǫC�Ը,�3
�`�b9Qs�- ������{��퀬fT�:rhU���{t���Zf-�sw�"�]\���!����TY.J�q�jvc[�b瑙�y침(>2�R@����ѽH��yu�n��Cl��GN�	�g�27�X��y��z�Sq}�]��}�K�Y���wC]�z<��K73+�P��o���"�t%������#�b�$���7,
��� �E[�������y��o^_�m���y�+�I^TG#:�3Q�nbX{�_l D(�.��p&�S��ѽ��m,��������4cR�>�h���|L�N���{f2)u�NV'�{zٻ��;s�
��۰���ׇ�zۤZ#��k�fE +'mc��{A���w>�iN�pIv��fj}Fe�K7�N�������EVgf	o��N���s9"��v3QZ,c[�5B��X:�u#�Z�p\>�֜R1nj�ųX�
X��v�ṫ�h���&�f$lE6II4�i�ۜ���L]�]>8��U�͙��Ϗ�Uuޤ���]����f����(m��Ȩ�VL���߮K���m��E5���%���xټ�Ǖ#p�ѹ�b%Ot��
}OS��٨n���`h�ڂ��|(�'h����U*��j�t-���p�R&k��4�1��`y��U:	��� ���-�?�R�Xۦ#����V�۝M�7r�i3ol�h8���ƥ�`ͼ/2*(΄���,��(���<�����2A�j�`�W�h����h�6NT�>++&2���#w�5glٖ�.���̩W.7B���i���j�z��I�{�oJDE�p����+}̙:�N�9���NU�#M��9�@��ՂɁ��y�4Ex~�ɘ��J�p������uF��m�6Ђ�H��[V-�i���D���-�#vs
�[p��)Yz�wn��s�^�D�j�-	j�d(�έ������T-�[w��y���N,�K�3y��	��t����һ�&�s���RA��j�>4Ť�!4N��Ree�u���S��ekyu��D�Z��	�ȋ�Q����7�t�V�Y����7FK݊��g���*6'����xb�����f�0)w|:.*�y� �'��e�y�Ю��Ctk�
m�!��&�i�{aYs1��c(9��dM[���5٤TF�"�����(��*��X&�C���A�FXu|i�@�v�T�U�K7�A��|�-�06��̠'r�a���2��/#�.�u�m5!&I/U���<�Z�	�4�yp�oJ�V{JјE���Ƈd�:$qAyy�9�]*�!w$K5��9`��5��7i���F��/@�b�kb�k�Ц+e��4n&��Zc5��Uaa�Nt}g5��GVI�q�O-U2���:5����@4��w�iH̬�u2�q��mJ��j�r�]i����pm���B�ܭ�ںJ��ީ;{^���q��+S�]����a�ٔ�P[ω��â3��X��ʇ+ $�I;7��,iD�t�{��ΝÎ��}{�����M��n���X:g%Ŵ��w�r�T+Y��I4�ˡ�VWt&�y=L�ot����Z���b�����N�kUm��������G4���4;�F�)�Z�v�o�TG)<����+.�Ѷ;<����wge��k��k5(�=Zr���0rή*Ս� �}2�EpH�g[A�p��g�s0#��Wd�������5�G~����k��6$�� �1Rz�*W�j�37l�o��Xc�nr���QVv��v��l�l�~_L�-�je��������x+�W.��z�i��h���s6E�o-/e &�μ��E�s�RU�̥%^)�T�J�w�u{6��|c�BA[>�PThB��,�[�j�^�����) ����3��[O�'�Ȱ�05�nؤ4h��V!�]��%�־��yI0��w�R�^���G��ۧ-v7x�ˡJq��բu6go-�d��q�SY.��6��m�Ȳ�
��$Pf�p���_�.�>r�3G���zh��-���<�ءe⥍�˛X-��<R�y%nh9�vޞ�F�R���.��3h��ESÈ�cW`�t�F`�q̏@�4L2���؊���d�N�ϫ��;��wI��8�٨��Fj"�8��:�_;$C��_�������@�P�N���X�K����</^<���\�qݑ��[N����vب�CP!��G���ҧI`R�(�ni�m�6���t+���ZX����\)����f�{��g���`��*ȶQ���K$�rE�Y���pɛ��9�����F*A����}�f��2��-$���(���wD-Ac��]��,f���J�y�+[��L=�'�Y��r��L)&�����E�7�vcyc镡r-��s�k�޺���ʭ2�˽�܆&�H�O�nv6*����!�8�/K��N�ȏnݗy�<��E^�>=�IՇ�#[�,�VQh�S[�4�7D(sb�,e��[Qn�WX�4Ћt����JU%!���s�1`��R�3w|����J�7y���#�nV���h!���Q�M�KW���P�v2�ƴ�;��RTHS�>���bԼėM���ĭ|Œdo��DepA��Z�5����++�u�ї�인Hu��qz��9
A[��u�h9A�a�xM7@uɣ��
[5f�>��Z9��ݎx�"滗�x3+�Ф���ܶ�����	t�7;��Aa9�+t� >�`u�v���.�q�RܝG�m
f�5g\(���Y::M���OR6��V�� 	>}u=I��ف�KW��B��vF��Ni-��[�G
Mc��.)X>[���6f��{�w�kc,��]MT�)���'qo�E�����']�g-�ȡ�C]�M҃v*.WZ���tе\�l��t��U�1��jf�t�G�7��K4�}R�z��v�{�I=D]�)��6���k\�c�k;Fs�HY]ěn�ѹSx��g�ި��b��@�+�JƠ�~ �\S������eU{���y���Q�:J+gL�k9f㮚;��i�U�T�s���spK*�Qi���L��l[[�Zś�Bj�"5Z�p��2�_*(��jQ��Bx�|>�,_�l�lI��e9�C�v���[�����6�8�
�3t���\Ɔ�A��V�_O�R��Ȼ
�����_3�)4�"౼�]:��eq��C��� �k�(k�l�"���f�*rn`]�6�� &no#�@:�u	}hu��!K{�x�J;��^È>�ujq���Y�q*mI������\�Go�F*�ͧW�"&�_G���%��Y���R�@��㸺�:�T�r	ǳ9m�g�اh�^PX70�t���M+��ȉIML����NU�9|t�X���� �RD�U}:�r<��gm�r�	v	W�MLuE��B��(oR!}{;^�2iFlʗa�,7}-�Ui���G[����5��܈����Ӄ�4ZD�5BkN�έ���XB�Ҍw�6e�{��ë��-��sD63vl�J��1j��zjSv�:���.��Q�7�j)q"
��ᬩ
�i�j�2m,�T��x� �v��=˹M�a��n�"q�KB�;�ڏ�O`�ou<�td]����_-���m94hsw�����\�|��ۛ�ȝǴR�IW]d�Ձ"9��qs�7Gw��ve0�zُ��O�y�dIݥɛ۔Ə� 3Y����iX,U�)�PMR��H�P�2�e(�J�EX�ю��Ʀ�U���(�A�+Z����1-�B��b�6Z��\2�,���4�Ō����,X.��$R(������0�)�nd2ZTU��EbX�QRڃPQCT��RG-a�VE���UM!�)�Z�%J-eX���ULmib�(V��$Qb(0Ak��I�����`��J�c��Y�i[Z(��T�
����Ym�T��.�Pb(�Uj��*�T(-��-m*�����ʕET*�Q+,T�b����`���iA���������Җ�*�R����Y*,�X��.R��(�eJTb�U1�ULj֕��Ab(�HI �| ��q[~X�G#Ŏ� ��:�w��.sJ���]��̴zν��-W�:��0\�7}G��T!^�ةcU :����dx��@ߢ��;����һB���P�Я��p�<���{gf?�n���w4<:\#�H���f�����l��X�a�>f}]ʰ> T��>�w{����ݩu��7����2%ު�^)'�G�L���1�_�������
DQX乨l�5����Ho��}��"�:�m��V/-lw�Z~�$t!�&�G���osǽ��dp��lq7��c���j])�6�֛��y�b�O^F`�k%Őch��A�S��3#%�9�>˵@_2GW��4��揄�g��{e�No��r�C<����2����ި�L�)-�=X��ߍ�W^G��8��\��� �n󽘛��==��2�4�%�gfo��__������k1��:]�"~�#���ss�N֏.�M	�x��2�gl�V4��\F��\p�%�5Yd�aYuP���	�n!�?W<��-�}Wu�wNy%�=l�8M��H�W�c��_��
-�Jԭ9(KW�О�{n�E`̳xy��l\�t����NѢk��P�;f;���d����z�q�ndܞ�ӯv��`ru�x�a^61�Ӥ+�V�37�=��NB�5ϯ5T��u<}|3����gkH`��i\c1hC{Ľ�}wQ 5v����ep�,5�DW)YN��r��Ԗ�[5]����SC$�.����]|c�B�}C�0��ʼ�Ncս�%b���K�2t!s���&+�]�ܞm�H��q&���8�U�PU-]mX�^>X3������,7�YHPS�Z��{�(�/�K4�w�Y�[�r&,��D\�=��O(Ϊ�l��4 'P� $U��V�#� Hn��Ͷ����眄7� _��hlw_��M����"%��äa��i�Ŗ�9f+(�˱\�Nt�ѭIұ&O��Q���w�������$��@i]��R������*!�֜u�S�0�{�g0�A?�9ˀ�D+�V��N�|R��eP%1[CNPuBo���P˵�F^��m��ʄ>�εG���|zGMqߏ3��(�+�g���o������r�7=�q��R��ͪ�	�����+C|-��9aO2�!'5q��kQq'3�{ko,�5˪�� ޺?jb}���%R]�'�z̫����VY�S2p�7��/}9�u��ڞ�s��,���[W�h�r�ZX+xA���z�M��<!�b�&�T��\�v���'b��&��r����09S\��YV�\�)jݍo��tt��������L�)˶r�Z�8��q͗e�q����Y�^��WN���,KO���s.�V�����|���L�{�4'-M�.�s7CO�L⃯r"�؍�d9,
N�^��ѣ���b�S�t-�:��P�կTG{.���=�/���{fJc����vb�`�4z�vz��T!��PN랽E�z�'.pC��a�ː���D��7��~ח\�c�\.P��<�VMH�����w&�yb�(і۸�)��=�Fx^��__���+��_��?Czi��F@���vuN�S�e&��՘����wOC ����a"q�����>��C�u��������,�iSW+8�?K�M�h�|���|�J����9}�:�i��㙘hvk9?Dz�V���tש�yc\��3]%	�P|��iW�5vX��ٟ@��z=Z�j(�rF�G�=��$\7Z#"��vh�OQ�T�(�1�����-Gڇ��mz�m?oe�Ν�78��T��4���َ�I	�	���&R5�ڥ[��zK�w�� �3�������C�rn�w��}S�ŉs�Dswp�t8A!�4��F�B{�9Nw�.��K�yۃ	r�Un
�M*ySF�{���{�wli����1�o.䄮�ֺ7�V�=�1�1l!p�Z0$I�6����w�h-���zt*�!�+�׭���"�Q2�y�3N	�����s�f�\5�B�Xgܸ���j�b��|��7�N涌L)�_'F�Mq�ݰ~{��Z��<7�{���³ւ�|�x�~�7��1}C��T-B9ͮ6vQ|xDȇ�2{�K\�#�q�M��b�i� Oo�x�?�ylM�ڴي߲�1p�ar#�{u[ͼ�Ҕ�z�5�A����6�~[c��T)��^f#^���V�J����s�jn��s�.��o\�17M��%YÀp�.�L_o�P�i�5a�mp��Z��q�LrGd�t��Y���7juQ���3خ�C4PR1���őx�i쿑�^�&6�=��s҆�;f#��q�OV��@�"o�&����.�13q���Ζ���s�HE��f�����왾��C+��WicYR@�E�?-
j`�*ep؆�:p�n��R:��m<��5�h�=���g�}�2��ǟ:� �O6)S=�9\���49xW��QU�Ӗ;��v��B�OW<�j<�>���a9͘Nԡ�x�SDb��|���c#��z�]M�����ɧ@��>i�aMMqX���+s��JFot�`\��\q[��1W�Q�\�N��gʏ��Cf��2� w6�e����oL��e
gjwq	��&rhX�b߈J�^	�WP�]SYOc��Ձ�CG@���X7�8`ѷ�b�]M��C��N�{�P��{�N�q@I`X����ޣAF�&�if�\�f�������R�l�ڰ�zp��ޑ�<��b����n�!���k�.��R��֊�4� ��&WY?.�_�?��4蝕�<�	΂���q��z�+Mmu�{��oX��cg�HX��Z��MB�뇠Ξf�Dq��n��&z��Nzh�kE�,�Vo�'�bA3W���]OI��fV�̕��
{����n�"��p�����L�0�&F?z�!�_����u-����#X�.��#n{ʛ54�'f=͉ꏦcؑ�5S-��n@	�d�E��;_z��^w����-���U�;�;c�Ѥ���{�����`�(_JZ��0��2��3�	\#>J]ֱ����q��W����?.2�W��������`�*�0���*����<��^�[���oj��͙���s�}C����eګ�����5��S�>��ĵY9���S׆.{����&g�I�d?z�[4$��I���޼�S#�v�v��J��K�ȸ�I�la���,��6T&q��LU�%ӐG���9�ȸ�J��uӶ�`d�a%�9�6m�>2����8',C�[&��g4�f��:�ǹ��d9x]llzX�Y.�==�Y}��KR]7�
Χ�Bp��j����_����g-�b��Vט:����{c��p���4��Z.R\,�3�ί���/ G�p�;E-ADr�՜���W��ЏT�]q�o͍�ηf��6� ��xh9��3ҺZ\k�v�zf�Xi�)d�E��r6����r�x0�\0��rP�=%"dh_V��:�s"�TFh2n�=��ޜ����"�]S=ӫ�S���b�ϵGn�؞"ƕ�I�%΀�iάou{N`<޲��ĺ�x�_l"�y`v����_\B0���C7���ט؉YŽ����uH�[�;����W�)L�����<�z�����,ӝ[���Q��k�/r�>g���-�G ��� �:����B�"V�4��V7"����ݻB�(V��j�n��w�:e!��u_����I"�4X1�񤡄aht�Hn�HLn��um�4M�p�pG�h�L��}_wm>ߢ�9�N��b���@i]��\)����j�L$� F<��n�az�q�#�SIJ�f��2ܚf�ux+�<��]�L���1��.�q*3��	pT6���NWes;B���[t��hurkw�"Z�s�)ϝ�	�0mAd�w8g:o��G�u9��Ava)���U'<
���Y�w��{��]��� O�P��p�lU� }������5`�!��J4=Ces����Jk���ݓ+���2���d�h�� �׶�<1
��e=8�6Qn8{�J�\G#��(�(t����"�y��P�Bװ�Y���w�k��V=�iąx��Ŝ���?Iu�\x��ژ��L�d��a?e�˺ɧ�OV�,��-W�:5�D�NJX������V���+2p��`53wlKH�=�벍�
��Bσ��"�؍��xϩZ�r�Y�ig��b�x^���>V{=<�f�|"��qڋ �+F!ݿC��_.����V�ve.VuH�󨝞^�A���2�8Y�t��bu}~�'{��q�Ф�������f�p��Tdm����]w[ݾg 뾫�xkp��n���JQS���|ڧ�L�$����ϗ�C�������m�=ӵ�N�#���΅V���Q/B.{�t��o��_؇�s��Ь;:����^���W���7K�GP�G���Χ�(%j^���x~�=�C�.�̝c�ͳ��FFovaiRQ=�C���p��.��\�0Ｅ~��-���m�w����Ael�F�b��[��i4�
H�ėY�r���1�O�c<A���ܩ�,䝜�(/v����v��r��+7����#ۣfZ��R�ϜY���J\|І���r���@-��Q8k{���E,����bN��Ht��K��\`!6J:BCF����;y��DN���%ibf\VM��o��6�Q2c@�00��Gڃ����Kt���j*����1�b�ü��la}��)}�G%�JQ+44�0��w%>��~��4�mR]�F4��X����8�^κ;k��cÝԦ��M��[��|fU@뭷�%>�조�k�谚O�����2�p����ԝ^��3��'��]�������=��jڥ�ͻ�X5� f��z,i}��f(G=��f�x�R���Z���7�k�glW����$J(�Z�	�=a?�ylM��W���'WBr���:�h���&`ܺ����y�S��t�Q-��6�]`1�T)��6�9>/ �^��F��譤�J6�����U8|n"�;���K�������]���ՇT<4[V�^g��F�9]<�fn:���1x�D⧝Jg�\9�F��w���\kO��+j���]]��ץ����������+�V��1=�u5�M� ���+s�.O� �:���ees�к����䯈�F�����e������G)e�W�K��e�oW��KL��Y�����pPu�p+����d��1��&;�^M�^ETFg,��:���!���M�}7��nk� ���������Ӌ�uYQGM5���2w
ޱ��H"(�HlC��y���U}7����zp�|�:v;\_!����X�^�x�KU�l`oU�����<��ؤ��s�ϔd�Q�Kdz�{��Al������v��L���{I�9����{k�ZD��Ni�������+=���R�/;�X���Y�8�/�<��&-g�@@�����^ǆͳ��U���ZJt���g"5�'�N�L�#�|�|���,9����)?	��䆰�n-�����z���V. �P�V�Ə�\��Oo�vs:��߈�_*�X3�z.N��hX>�����$,
Xz׾Jj�����l9إW11��uQZ1X�nr����ﲣS��>�%����Z�EJ'�s��f*��6����8�{�T!6q�%�ػ}�Z�p�V9��ˎ]�.�0��'pN��j_S ��|W��]#��k���1��<�GW�Z��a��5��n���{9b*���Vid���[շ�T�k�t�F�S�[�4e���� :��K1�|�&�+��<L5�d��&Gf�F�XX]%=�m��xS��~}�irݢ�gĝU"�R�}`��`����N�/xe��ܗjro��_e�K�g7Ɏ6�Yݷ��qn=��[�h��>��O-A{�e�i�~S`	Ϛ���S�ٸ��=��}�������ӆ�[RO���8���R�S�όs��#��a�&1�X�"g��D��R)I#��þf򑼳�k(y٢*��	{��lt���,mu^n����E�[�a��io��I���9M��{�ֶ�m;71C�˵_+�H�p�����o�=�Z�~%���H����+����S�j��6Ծc���s�y�1 _O�c#��@��*������7~1����C{Y�w�'�g^u�l*���?X�w�"~�#9�3v��R잙�ug�l'�BI5���dh�/����k�lFn _Q<4��
�zWXė��y���.{pM��=���>�ve�,�l$-��Sz ��\8�l���#�X���������n�5�@�9S�˺�M3�P�62r�;�=j:��"�䭢���'xs^h�b}GP��zˢk�Ip�gk"���
;�+��i{�|~�}���ok,��������m�X�)-�n�C�HrzԵ�p�_J0w �g�uub[M�*�wǆAWM
���8�٬'}Vj��YԺ���7-f )J��y�{���.�{4��N�k�Mq�B�5[ˈ Xn:2,N�4����e�D�t�j��^/�.]f�|s4b��#d,���T�E��;�A���a0��Nnȫc�|��TW7��ڽ��=���c�v�b�jy]uaM�3oT�npA��.wl���K!"}��Y��9�]�+�dٶ4�&���H6�s��yJV��֣7F��6q��L��	b�Z�fB2��m��6Ҙp�:2U���|����<����(����� ᛴ�f-ڑ��wi��6ɓK��d����w��!BU��'*B�_�+�����7VH��CD��N��8��^�����U����r��soK�aDӽ�ooTv����5j�|���\=�5Q���݋�^=��F�]Kc;�ӤC�ueu��6���̘���Y�m{�tS#�(���]�U�	�y��ל�O>�y�t����7�9�c��H�θ�}�2��:O�t�^Ā��ë�r���	�' 6LS{Mg_*Up�;�V�&��S��!}N�;��(�I�L�n#����½#bCi�:߽�ޓP��ͻ������2��A��sB�N�fl������4�|ىA�%��B����{/˔(u8Yݎ�D��M��|�]G2��c5��\�1�^�<�5L��ηm�i�}7R$�h��*[i�!����t��w���:�%��n���s��\
k�r�W��*�$�7Qٗ��*oP�n��4�˪�d�$74MIӸ��k.�ͩS@VWQ��uܖ�G���U_�g�]�*9e����xAh�K���\pkߞ-.5���$V�J�Jj���u
������;�����Ԑƫ�����c��Z1�����!c�wJN��o�����2J�T5ħ ;Ġ)T\��3���~�u�K�DXS������z�X��<C�KG�� �R���v9�ێ�Gt�u���WW%IQ�y�>���5���=�N緶_}�l�:p7��Ư-^j�PC��J�ڷn�.7�[G��/������7:��XV*q$���&nM}����
��
6M�v���9*wuJX��(��$�%���7*���q3�s�!Y�hD%*��0���U�v	[oy�2�49i�Y�looQw-����������/�e���x������]��5��Xes,��N�g��3@%D/i�ݻ��ԭS�a������ؔ�3x:U�G����j'���lvT�R�Y�����h �s��7�J�O�W�vb��"���kn�)q���M˫�ޣ�h�.��2�k��`4^]I��3ctd��R»/w��׸�X����$�ʷk��\� �.T�:5ؓ�n�sg+i�v+bb��s�A�+31��;���^��}�� �Q�'V�cR�bňȪ-ed�ũM5V`�1ıQ�mPQZ¤)hYm%l�T�kX�R,��TX��B�cDhU�ڍ���j�)�UU(��
�(j�r�+(�V���q�`��)�fE�m
�V(���Ar�6±T�QUA+@X)YQB1�E(*��Q���������ib��DF�ikeU1�XeiEE����PѵUE����"�-J�eJԨ�*����EX�������E%��dDV6���"EX�RҩZ�fZ�Q,`�c�,��2�D�#b�T%-(�ы��B�*
)YX�XUE+(���H��#UP*�KiR*���EDED"ȌAA`20���`��j
���+D+QE�*%J�����F#-�C*�X�-m�Fڀ��UUX�Y*�J[%��QP��-��A��4k�߯�}�yه�kQWnDtnRx:�Mv��}����x�Qg^�t�5��Q���n��Uy��8�7������#�=��3Dj��w����ך���xô��:�>k:H*�ȉ8혓S(c����i4Ϙi1 �S�q�hx�!�T>aS�y������u�3�g�*��Z�z8��i�LC��Y��7�ދ��4s�o3���p��LT��̊NЬ��9ָ��d���P�i�E�J�����(�I��c��|�OL
β�S�g��<���f!�z�.󤂩8�����<Hs=���[�4se�{Ͼ3b:c��wM �����k;N�z�L~I�9���
��U�w�:I�V]�P�z�|�C�՚@�W�J��d�6��O�U`,4����1퓲��K'|���(�d�l�jc�0�1o���8�{���:H*é�z�I�+��u���q1�0�Ϲ�|�2VVm������2q�YR]�c=�t�]����;5{d�iQg=�y�S�8�Ǉ��hEע��S��c�e�v���ty��>0����LCi+�vj�:a����)4��$��Z��8��gz�I��C��3bc���3��Ħ�})(^>}����DA�����LtǵN�� ���vygJ�TS�����4ɉ�*$�j{a�6�x��ތ�遈q%�s��0Ǐi���I��z�T��=�;V�I�,X̭��u�G��k=�������y<�%B��q�&!ީ1���b�f��� �M�S��<OĂ��Ag<�b�C����S!��y*M�XV_}�<@�8�N���0����)������%�V�y�ܳ^���Ͼ*J�����hY�%I�/\ߝI��X=g�fP�&=0�T4��|�OS�^��Af�x���>��AVtwC��O�:�;a�1]!���ҲVT���ׇȚ�;��7�=�|I���!�;މҳ��L|7̝�����}��& x�:�zԘ�x�Xt}{CI��8��Sm
���ǽy�4��W��<���v�Y�;<��Rm�����!����W�vc��vs�`"O���~����y������11������|�'�z�s;H*��*u��������1Y�J��״���'��ް�CHx��ѫ&$�
�%!5�g��^t��|�z���\-��<	<�G+d�ϩ���\��mrӒ��6+��~�S6����ʺS7oX�26�ߡ�@�Ŧ+(�M�=,����j*ۨm�B�At�b�ˬx�R+�]zͳ��1+M��X�B�cÉ?�WΤ�zuN��Wa�!��eoΒϺ�G;J�L�g~��4�Ry�����W9��C���OS����=f!��{��v�Y=��C�1��j� ��䘉	���~יU��p�<��z��:@�%|Nj�񀡝Xx�mua�;�ɶ�:ΒOY�������l���oy��'��ݐ�>ΰ��w1�o��w|n�9�{��n~���EL}><�)�8�AH�2|�ϓI�Vt������k'��1�C�
��]�}�3�;H.ӌ<��G|�Ę���a��k<d���dP�m��tk::���٭������[�����	S����8��v��VL�4�Y�ět�I�(bAz�:��Av������3����+>g��x�T���f���=C���������|zyg�ｆ�zn޺>�'�ٙ��>�y��LZI_S��$�T<I~�;�I8�gy����obO-ea�n�:�c>d�P�1^�a�4�PSi��0�0�f�|�Ì���{��+̙K��3�	?���?2�̏٬!�AB���gHm6�2o�c�
��]���9��O��s���N�t�eM��I�&��i�+
�vOOz�I�J�:;��,�%I����~w�:��z<���>����p<���1��O�Y;f=p<�t��q�;�s'���!�ְ��>�`s. z�'�T��05���6�O9��%d�ߝjtͽ0ۤ���kb$������U	˩����b��/�#�K"��5�I��{��d�Y�%{2�hi>d��w>̑I�+���Nݰ+>I湝;d��A|.oG���'3Hy�L@QI��}�����߾�͛���y��\��w��9�'Hc=a����3hbz�zCI��û5�LC�͡���IY�~d6�!ĕ�>E�$���ްz�*M�^��2u����f�t�Î�$�|��~W�o|}���}>��p|�R��9=δ��*At{̇�S�0�3��M!�>La�vj��$m��<���H)�vf��4�0�����/�:��v�ĩ=B���v�N�q
��Y+#��2�p����N�NU1�f��)��0�Wd��c3WLa�vT��u�9����>�P��>����g`_�M�[�($or��ܬ�6�Ωf�]w'��P�у�J}�K����+x�*��Έ�#2_n�>�=��^����Ry��aXW�l��^tT;IP8��Y1VJ��7�CYd���*&о�;O2��P��N���z�$m���פ���2w���Q�]� �߬b2���^��;߿{uu����s�<|a����4�^$ǌ1<�u��U����Z'Ht�^'��5N��%I����|�víSI6�O�<q�Y��B����N��\{<��=9ל�[듁��N�����8�~���4����`"���n��Ax�ɾa��=M���L�0�2��16_{�z��
��w��i������C����DG��o��Utg�A{�du����6��*���V����K�񁏉�L�:C�>�i�d�P��y�J��U@�|�$�8������Hx��s��|�$t��^?��B�U!_P�����c(W�?�s^��RVT4�C�Y3�J��^=��P6�'i����m
��0Ҽ@��d�°�������x�i*φ�Ξ2TYY+�,6��d���g��ʏ�c��f?���m�G�뫟��{�������t�I�Ă�����I�����1Y;J�ש�4�w@�`�Θbҳ�<æ3N�c�<��IY�:��t� ����C���������213��Pl׭�y���>��5�T�2��s��t��T��>�V��+�������P���&�ɯ��N���m��n��^�
�3T=xΒ�;2�5�h�����<G����������̗�*��u��uﷻ�gHm
�s�T�!�;�v��b��<�xt�Ĩz����ޏ�;I�*f��bt�'��L��W���Cԕ���&�+6�R��T�:T�B�Oz~�gY����n��qiC?�m��*C�����q�'i�O%��6�C;��h����z�����T|s��ԝ�m*O3�&?2bN'v���U�u�CL+
����\�z㐬6d{d��D�11�<L|d����Ğ�}��W���4��P�7��2��*g_o=��m1 �9�J�oI>�OmVNҰ�뙴:H.�;��GHq� m�?=�~�5����eu�i�f��(��ڐ��FS�%��u�pX��ׄ��^ۨ(4�vQ�;��j:�*�Y
�akǂ��m�E�E&eq�MwWq��P��zڋ2�~�f�!vI���)pf�:z�h�#�m�֌�jtok{ �n!�5�fa��;F֭���������X�����4uC^�t� te1�q�>��L|�&�H�q����xN�q
�a�9�NՀ��7���ɴ�l
����i��7M0��sP镒������A>x"��E��@��H�_{�1Yy;�D��t�^'e�\C���S���Ag��tӤ��$GY��
�C�1�̲c�>a����HJ�w�gN�l��hW<>sY~����`�F�DV-yLK���3�K�Ĝ��N��%ea�����i����h8�+>d��s,1&����sVi�
���3�2�$y��>gHz�!�;=��I�T=OS��a�Av �u����]f�y�s���\=jN�;J����<xɉ=��0�*�2tn�'�T���;Ԙ�!�*C��2TYP�,Rq���eҰ�B�N���N���|��L}�1S����u��v��n��W>�l�'�$��~膕�Ԭ�,PĂ�����q;f����o2VVq�&;�皇hv�U��;�.Rb�\��&2f�z�̺@�TY=jt[�%I�*|�w���}ֿ}�㯎u�t�X
O����交:=��W�L�4��@�q���|��������	+�bA��y���1>C�{��:H,�>��:LC�1��1P�*u�+�˶�_��z�����*=����z��+93xM q*�fP`���)�y~:�^V��u�{��wR{-���i��<\F��/ç�3�W�B��5�ڷ^{�XV]���c��S�>��<�X�=��H����JCg3��̼��[���������� �38����NLLb��@��g=�;��.�[�1J���{��v���IU=-F"~�#�'Gc��c��ҫ�M��w7&���CX֨�:��ъ	J�>��k��_{R��[G� 5��[���Z�-�6�տaYL�+1�O��أ`�9�8���+�-��0U�6l�П>��T��절���q�f��S�Eb_Vt�=}�V���8��#ܩ���9������|�`��gN� _�A�M�&��X��w3�����1\-�Bv18�ve�,��p_Q� xF]p8CK.�	FX!_<�;�}ҟ��;`�|�iL��za%�3�������Y9/�Wpr�r���cUa�B���k �sJ��X��� 3gϣ��M��ɵ�1=Ն��J�v���S��|:J�V���3s3�,�R���Ĥn��g|�͓Z=/�ߺ�hA[��L	��/�����wc�E�ȌAq��lY�b6�BB�T���x0��[$V! �xrl����-�bGx�������)�=�uT�
]���!|$i�,t7�,�����ȑ/�����>�%���3����.�� \�/R��E_sY��Ǥe�p�����u�,���<TaJ���6.)Q�f'��S�2�nc�	}w� � L{��c2�/�ҿi|q� �e��펒�f1�hzx���>^}y��%�,
�r���e,e��M�k{(�q7��Tį��I�E_	���&��n�hq� ��V��H���26����]����s����B�4g;�Xta��:v��\���ʛ��r���P�;����*�W{AR�9�t�����
�ɇ�����)�f���[��|62u�m�T������+�'��;|3��?I^�q��6p�W �X��7�b�����*B^�<������k3�f��rzo���ќ����\z����Imi��	�'��\L�yW;�B�Pu����#f���n��*�J�Ud<�
�1{����<ځWt��F�x8����`6q��h���3k]t�>����U��ŵ;E#�rֽCi�qܯ>���c ~�f9�s]�F��9;r�Lw���?�yu��L\�7�͉d���������PK ���M����w-�PU|�j����ɵ�V�h��6��\��;ޭx'�ud_U���Dŭ�O�<��xZʗ�	�>��%��+#t�MI�t3-f߸��P�~�:I��_̦H��
��PZ�S,<?iW�Vڲ�I��=9]�U�օ���s�7/�f�l����!�����Q��(LB�g���	c2f�����[}��t�ǐ��[6��Vc���[��4FE�/���R��l3��d��:K�ޮn��<�'�_��(ĥ��"�w[Խ���B��5�Oz��x����n����j�W6�b��&��j[�UD
괩���C�zV�?7ò��)W���}LQsvLhw���l)+�
4YG6Ex�v.$t�RA�YX#�n��T��م��"#c�͔^8�>
��f��r�IA�or��T4�sw���Ѿg��,/y&�9y�L͇}}H�̯V��1�|���KU��U��>�U`��Þʩ<Y��rt۬��OT���8޾��4.����.kظ��Xw��.N�r�^��n���b������z�T�� ��.�����]%�;)G]������ug�:]nrz�U���͵z��y�]]�g����_	҉�3�G��W�%�еm�ѡ�灤��O}*u��0I[/�\��b�8�p�o�� C���U�{�J��j���\6���*<3�k�7�XcLou��Y�7����Z��v�EA��<�:�A���;_'����j�rI�>t�����O����Ӗi��/<e
܋�ٕ|�yO�\'rP�4v�\ZV{��J����u@�����l�d�±�OZ��|�*���>�x;���������(�V�@�F���O7�V+]tR��ju��HF	1s�Ba�XR@��M����E	ɴL�kJ�n��tMIv�uڪ�GؼGN���{%�'��ڎi%$κ�|�	t��/��z5ʷS��l�J�<tC�*~:}��^��Ɂ;�Jߩ[#��ҵ���� ��4nAf���W��a�A�s{n��Ӓ��۲�uv37%���꯫��u�?k�����Z1w��o���������P�����;�n��kef^��ֹ­��oW�C���b;>�mΟ+��jÔ�ʌ���s��(Ol�|q��7c��S5�^b1�U쭑�'� ��wA�)��3�)-�!t�w���%�՗�5�-�j���LP�K�D'�cGhG"�^�WzD/ի�2��aS������őAv[.cz2��ZݺZy���=l�[�mZ�t���1���s�:S�ઋQ��ޞ�*t��mw�`d��*�#[���䪊�w�s�������aL���n����uZ����;!jeP���Ϙ�<�՞l���P�*me#��n>j�Jz�T3n@��J7{]u��=���s�$g���;Bu�#R���k�m�_p�R�{����^n�{ԚK��}�R�x���$�W�(���^��ƒ`N|�ĸ�4�Gu��c����w̾�R$�����5�*�)h.;�K)�g�9�Jx�X�~oI���]`{n)�,!$v�nf*��w�L�K��Ø}��5u1'��b�y9��P��жuŔ�N$�im^���7I�Fc��Oz؃\����
�l���W:���G;@&>�{>]uq=�\o�<#��)ۥ�Ŝ%��e���Rȧ��x��i*'���̽���U}���\���XA7���g!A[Ӧό��f��������7�c���#'3��l�R*z�p:b�}�ε���1��#O��n�8}���XV]_ +�c���Ȅ���$1kN�a�A#��hʄ��̺��}}e��Y#����R�s�y��l�j�)5�eEi������;��-�ZC�~���:Ƶ_�n[F,t��O�a(��Q����2��bw���Frv�/�T9�u�`߹ҝ������a��8�L�����s�/{Li�۴!�F�L^۳+>�xswL$7�GM�p�p�� �p�IU��w6���*���u�|K�F�t��YwR��3�<)�����a�|6ޙ1���Ud�t�C\v����qN�+d��!Ԩ�-�$�EsÇ{�|�K�~�~��Pݺ~�f��2sqY��Yyps��?.�H�w�"�;X2 ��O،O9��Wc,[9y|�&��,�ݭ�}�P�ﯙ8h�ٮ���,��e $N�Ѡ�WZ����gI�]��p��X�=%4;˼e�MM�D�ҳԦ-��7ڭ�m�+%hE�᭘�Y�W7��n�ʚ��XyK
|v���()c �sf���p�1:һ'B�/6��@pJ�f�P��F���C����p�Ϟ}��|>��+9-e\Z ��J���Ͷ�UG1q������$�u4l�z׃p��
�C$s�j�y�e	\]���U�#yf+�z�	8����Û�\Շ2���x@���1JD��Θ�G\v�YҬ�Y�?U�C���Cm}|����1�cr{�ؾ_v*���uZf�y֮�k���7�~֒��Ļ�4�:���t,�.8�|a�����^K��<�`ޅCj��9�z��ކ���^�r߸�6$M����h.ko�F�x:5��O� �5���ֲ1?=+���g�a��5�y�9�Q{ث��9�^Ji�X�ʫ���}-XT�����(�����6KÎ־�*Y�s佱�:����6]W��DXu�4�'���ӪE�z��Jo���}Q���:}����l�xn�g�f�gb8М��χ].eXkO�[�wvD���5x���Pb�\�o3��v�?��F��G흽#�*��������U
����(F�����V'YM�����F#>վ��noo��� >͹�
��(�v���!7�q��Ċ㺸����dh\�����������t,��=�:�9p���:���'q$
�hp�,5®��j�Z�H;�c�S�s�)�x��s�i���߬BUo�H3Yz�4��;��L>�P;�a�r�lY-�G��ȷ.�����O����u&���VJ9(S�Wf�!\��1Jn=�Q��3����T��!�/5�X��FXQ%�X�ʕ�swz�T|q�/g՝r���0�ub�?�>j�p/U\P���T�3J�TPb�ܬ0X�>�L.�/T�)��v��u������K�Wh��/-|2�]�����u5���3�0���yL�ٴ�ש,���q78�Y��Z��Y���1-.�h�����7B�,���6:�ނln��V�!e�wGp�2G�7�>{/����
�Ծ��	l�9��鶬[��.D�b�w'ZC���}%: 0�4:S���M��Lѵ/6W}S	j�����2e{Z�#�4���S�eV�0!�ᘜֶ�6�aחN��nJRu'��q=+fR��v��Q�U\web��-����.��hN����3�<� ׽�E�>�	��V���J&uu<k�����e��\dո����cΣ�������WP��/4c��d@��B�V�ڐ�V �1�FR�D�j�Z#�<�w"y@�쿐��V>ܔm�O��oŝ���t��7����7JQ�K9VM)͖o�h�C�B�c���8���Ou�%	935>ۦ�C"�ug_^��r��Z�(�m9��҃����M�tʢ;�
�n���4�psn�A�CF�p��-�]�>��� � �;���v��>��٬ܥG�+�؏q�pc�ʲ���O	�ɇ��*���M�,�ڏ㎡S+ׂ`f�N
�E3���M
�snpJ�RVԝճV�s*�^Q˸��Ӂ1Ym����tSY{�����+��ռ�-gt�7M�cҬ�޼�U���b4sw=F��Jwn��jV�c[\��U����{-��˗{d�|�)S��q�`�o�\��t�Íњ(m�T ��V���8���1�9�K�D�i]������k��5 ����@PӵlmԜo�k_�ַ��݊�p�׼4�i��V���?��6��.�7��7&�geZtȠ�����B�[� U�^n�Z���ޤ\%Q�0���Q���f����s�87#�uj�HZ�e�,��u����vLa�beL�{���"X�j��v�W8���,�ٵ?����S�z�Y��	͸a��wm#P���讧�*��M7{;m��&����Lm
��Ihe�c�*,��c���s.�f��{��&�इTysa�d���=���ͪQ�k�(;(Sq��:��
���T]�R���J��7K���Eʦ0k�tEb��]d���˞��3�-;b.ͻ�.�n�욵� ����HȊ2#&�b(�,��(���VҢ�?\i��eE�Z"�F#+l��,�,**ʔDE��P6�-b���Ƥ[J,��iR�%j�
�m�-b��*�E�8�(*Ũ�k��:B�Ęő@��#P���eaE�� ��Ȣ��j�U���X�B����QA��%�,�X嫔XQ#
��-J�l"�%Pƣ[`�6ʣAb*��d*��������E�
��J�"*%A���b � "�(�F"���T�"���B��&�dUX��L�VV�0UX��fQAG-�b�X��UPQEYU�b�P�(�ѩEA��*"�����0���1�+&\r(,-()څj�ذY-�SY
�$TdQ�����3M���UVEER(���j*V��-aR)�DX�*E� �."�jՒ�Ŋ,�U��2,����XV)PD��B��&���W[�v�ve��Q5��un+���b����ڲ�=�U]��'+9b=�b"������5�s�﷯U�~���>���j���wd��{PCY���iڵЪ����K�Z*���<
�UEܱ�g�_UuO7 v�r���K��_.7@J���iyk��H����V-o)��l���C�k{k�H��}������P��v�3:����C�y�(�&G�%��/��84b��Td�#�u,c��{d���n��Ω�h���n��=l�6�Iͷ	�߹�OsU����3��0�j��V^����B����sc�Ў<"h����::��Y�<�uKDC}�wW��#Q>6���G�gz!�:����E����5� �{X�W�g5�O�#�<V#��G�z(������t����9uCW����Om�� ���՜�������\�B`��9PG�N5�x7ڱSs���{�P��)�Y��۷�*��/������M�0��m�q�L�=���
v]�l��RsC�L�Ӑ(�1��
�z�xt�#�.�:g���^.�0���o/Iw�=Ͷ8(����&}e���
p(��{��Zø���[��.�uX�߭]t������,hc�y.�k�M�+�^�U�s&c&��\��F+?$L�ڴ���!��)�X4�R�p����U���h`��(o2�*�ku�ڥغG�\H�k�w}H챐�\���j[�P���������D��t�J���V���w8<<�3}���ǉ�g�����[VX�a��9-��Kyu���ٕIx��z}]WҼ�^�~�p��C����c��Pٶ�m�k���6o�0W|5�Q$ߕ�����:�����"rX����}uv2ujd�A��|���{�Oui���fƢ�n���A�9P;C���{��Lȇf����c��P��S�C�z{)��gZ�j?+?w��q� C#�u�A�P��)��y�97g9L��I�C������:HGez?z_\֘������3���>����);ܬ�%�lϡu��Y��
��p�K�a���wA�)��;e�ۤ��J7]θ�c3vU�(���,d��Vz�.|A�1��i��vu�!�%o+���[Z3�M_�1,g�;b����J4}�%*_rkY|v�*�$�b�(�����3��g2;U�u�..{��ȱ��d��׈�47>!Mj*9�@E��# \#p�.�����㛨�\������'_�d���B?4�ֶ��\���v�Y�H3%�%�vq#J��L�i����lK�",����2�+��[��b��L�}�5~��=�$J�����O����H&�V'��q�xHaz+�j;��U�j^D�ws�U�mR���| �mV^�YӜh�ҳ�%x�}��¥�Y3�<Ϗ�1�5ZD�[��*kgm�7�[�:�=�/>�\:2IMF�$��}e��N�F{��v�Z�5/��h!�n��߀����5����Pc`�/�ǃi
���L:�@U���ڀ�'�uH�tvmZw��tw���d�͚&�ߪ����V���ߖu�����]�ƸR�Z�����y�^��ɍj��~^H�k|�E��CE�H�5tmxzQ����2+돊ut!/w�c��ҳ�H�^����0�s��e�O�W6�kMh��k%֚�o�n�:��xAaYw�
���G�˲F@&���r�i)�����G��n�%j��{.|����N��G�����D+�>ǡy�v3k��O'$}���Z7�3׹���]�1��s=1pѾ���=��:e�\,������|0����p���s-yxƅ�d��#�]�	�G(l�ݗK��K>�m�B��YM���RrrF�l�/�3T�9?-�L�ݙxn�9�2n8����\�-�����n-k����S���[��Ί�Pkʗ�l͋g�9Azcm�x��遷�݃���y����_k�z��1�Z��%�:���g�w���B��h*�t��NX��F\w��������1����v��YJ2�j�D}DGЁ�0�xt&��K�A�$m�/�y�խ0��I�t��ԇ�Ɏ
�#20�n	\U1�^䀘�.�y��epr�������PHC�W��y	��b{���t��U]"�s5c�ǋ{rV��Jk�n@d�N�X��W��&�'���B�[�-_�!���S;iA�d�'���6�4|�_G
><I�筓���Oy�5]�=L�]�i���y���cɡ��7r%��m��Xu�|�����ff�z2G��ᢎ��M����7���Ai�,?8�׬�b���Rq��o#q�.�]S=r����A17\d��̂�	�S�6�1\��դW��Ԇ���w�,�<�=��2s��iظ��'M�q��.��<ぺ�@,#�S�|.��@y�ƨb�a�+�xs�dߗ8g<(��q�g#��w�jW����Y/hl�{NJX�vk0B9P�\k��H��唧��w��j{{�^t�ω=~za�uS�ծ$��(�[֫�9�^Jj�lO-�����k���>��ݛ1*됡V��K��ș�T���kTv�vc}a<Î��a�� �N�B��.��+���lm����#
U���g�/�ݶyN$Ō;S��Kb��P��<�:�xL�5|���Eq��$�$;��&¾=.Z���_W�}UK�i.�>��+W���s�	Bqo*ѦgJ_�LO�ݫ����E.�1����L�=���vN�V�q�h���^�q:w�`��Y������XZE��~�&Q�k:L�F���4�;@yթig1��B']|v9S.FC��h��ì䮺Ĺ0_Y��El'�Ծq��L}s�iQ���}xpD����G���C�����ü:���3���3 [3��׆e_������4���ծ�T%�y���wb&�:�����C}賦���g��}��g��MC�yh���%��FeՁ�|�LE%|�Ua�}H+=;y��E��V��j���o�(��|��Ra�|s,gx�3��8�8��dt��ے��â�ݮ2i�<���;�dY�����n��)պ�Nh����
��V}:�3;��^0����*��
���+/(L�j� J�������w�/�%V+D�y<����t���"J=�Y��f�4M}�i��cթ:�t����.92��"����`~ˠ���W^��*խt�V�tN�dc�k�͉����m��J����z��u%.��b����8\l	o���~���Pn���,���2�f��h�J�����!aL;��ͬ���	�-�^���ܑx7E®EEiW��RJ�B��ժ�C��	��<��U}�W�9�j}g��2؏0AT�n��\�}� �p���y�A���\n��C��1�9,O]ұ�k���Thax�^k�v���O_�\	��5�6*�4n����[C�q� �S��B,��u*l<ײ�	^�5��Dȇ�2{4/�<l�	�R�-(rʣ��0u�1���L��[�H�U��^�3/�o9}�,IU���c�S���d�{c�U.G�f]iO�F�#���J�����)��c�����dQ,��2��ރwp���<����yˏ��5a�8h�����药>5h�f��NW�<8�e_-#;�j���hl��n���</|n�C<!;�p���e�?�{e*�N�	iW��\.���F�r)C�Oڌ�ym�12�y���l�oOsˤ ��E$e|؜�����,��h���u�>���n�⾓1����#]C�7���w��k�o�z�v4���}k��tj�,	���a1�������1�w��~'���G��Y9 ����U�Q6��G�Uv�N�'�5�{�3/ԋ3�����CQ�[� Uo7��kTsE�au����Cn��=XhenV5!;o�Ց��3@�(4¬<�
e+x�Ř��CSJ�Io�E*�8�ʾ�su>�	�e�폙օ�rJu����}_}_W�Dh��g�1R%��KIV��+�-�z1Ej���J����s�2SeH��`9PT;4�S��^������&(A�JZ�	�6rire!ԫ��M^ڐY����%��K��Ɇc�[�� @HXA}�i���9C����W�}�z�oH���Ty�N�����(:�o�� /���C|
E�a���D�6^	��	?H���j�l���k�L�Sow��9MY�sr�wCgfQ�d	��{��	���2�{���[��݊�k+�#�BSz�>��X�a9:��c>�Fx-�	3ǽ~GӚ ��sZ�:�+1_{b* �>���=4�x�]Kdc��sz�,҉�>��RZ�!XQU�תb�����4cF��o�8��?�p��WO����_�_
�>����{V�#�_�w�%Iu����t�x ��G��[���)Kő踧.�%����x�j�
[;�E]�!ȴ�&U:.噲����vhi�lCc˱C�l�T.2GY7Hm.x0EC&�р���t�і]���QW@�l3\�)+4�h�{v�re����Q2�ԴfE���	̶vI���%�Vc�d��'�dA䴙�J ���]���Y��:8�!6����+4�z����ݙ�V�@`�k�O 	�ٶr�evl�N�#u� m^.����`�̒�W��W��Q�l����3K5��˫�l��콥�j��W�����*�����dD�쳛�I7;uvz�7n��ݙ�o�k��<)pm}8˯v�n���ԁh�T�8�z6��%V�l�5rwn�dFh��N'��
�a������k�1�;����z��}o��'���y����v�g�J�=U��%	�v��Xq��X7I���9/�A���'m�����=���렇����2DJ�o5��za.�������5>��s��enm��=��~�ro9n}���W��_M��VuG 3e6�R����t"��V�_ON	N�ȉ�zL���?p5�2FBes�[��x�"'��V���Z�]�Ɖ�7��nrgS���+/;�t4;k��,��uh��
>�dᯏTl��^�(�@ $T�ؚ��{�.������kH`47rU�������ѽ��� R~��5\�yW�[ޝ���V-��� ѾX~_8���+�f+(�T;���U�y)����`m�����ޜ��\�޵:�uɈPueT/��Sk<�#y!�;e�nU앇\��ec�+wIgҰl���֤&����V��As������бe�Y��<YK������\���ш���I�kw�J�p���F��r�v�g�����<��](�)�"9��?*��<w(�0k�y��W�	%������3$}m�׫���U�I'#�+hi��	��g�k��;�{=�Ն��\�k�zP[�a�l�:Qht����L����X:~ǿ{~8��4���L˗uǶ��x�d��QO��a&�><b^�ќ��ΡF�W���Z��+V��g�`��ȷ�B���P��^���FM��)Y��\��U�L�t,��3
�Y��Jz�6�Gc]�����c���ێ즍Ơ�scz�`c�v㿔�>y�۶h|d��ԯ6��uޏ�����^q�F�Zg��0[y��r����9;r�LwwD��f=��~�u�zE��|� 7F�@8m��_ �*����]�x֎��1�[��q�|��V�,g>:
������u�X��|���4�;V��-f�s�!�{'l,�|I	6�5��U��L�������6|�s���~�2���C"2�>#]�W�&.��Q���i[��QF�BE��-˓Y"�/=�.�es"�M�[4]A^3{rW����~��MKW�XUJ
͠�=�X���4�s͏��ǜ32e�c�˭)7N��7z��J�LY��2����}�+rs�/��;]���={�^�=���| �Nn�'y�Q���K��l��g��I�l�ѹ���Izn�AdJU���ሊ�;��3��U��9�uB����u�A}'����'}��1�c�g~xQ��ĹQ���M�B���q��q ��~aq�a���@C�U���/v>�ZO	^̧u-Fws��:�r��T��i�����m��'ц�o���_rfX�#�8B���N�ӌ�(��!�痛�3'kY��⼲7�07��+�[���_�H��?W���6�4.>9���L\r�z��)=2<�Y+��н���(�kDB{*��N5�{��4n����4Ųt���sf���ָ�t;}�_2!��(��<��߁��_{�:h=W{�':�l7Z���z��=���0S�����rG���T�����P�r��J^ؗ��{72�Υ�_�S��1_�
�Oa�5�X����[�5 �k�:��g(�	���[�f��X����o/���5D8a+��b�2����veU��zx�u���m�4\�Ru��0XU#����w��3�AU������;D�Ag.�|��+B㽾 ��Q�k��3t�͍[\j�n_����=ܵ�z�S��JJ�t[�'E�w�[{�ڝ*	�t�X}i��IE2��+��n"Ûn�OZkF+قm�Hh�8o"��S�6�y]FX�w��6��R�vq_j� k�.N�ʙ�.8�K����Wd��V:�m`|Ԉ�v�
U�
���ISw��\���>n(��� ��֦19�뮑��ub��΄���؊9�XR��	OS�)�MŹ�ͦ��Rt��i��_mrW�!�H�g�{���Eh�
ᾴK��AXH�W��X7t�M��U���H��[�������>/�;W��8�04�eC�+�T7cy����3���[u2�S��"�#M*j�[e��(������6K8���3�Z�[���YB0�<^�X���W���BU�]]�\mBv����^��#���ܳwI1E����v����u���6���F�Qy�&�¢�r-â(��1^Z�ܺ1&�c]"W�]wO�ݑ��9�d�i|�R��
Ƈ2��{�ʖ^EY�l�˂���*%�X��k����n��j�B���!��eֳ�z��]��w8CW�d����At�bc�8���V�)�7H�-x㆝��=�4�����&]%[��*��a�{x�!�a>�a�}�6�j�(r��v�T�z��s���!ڸ�W_>�C4w��AZ�q�}��<2gYJ�*���k��e���{I��G1��NϬWުwf�2K���T�z]�u��r�J�J��*V�\
��8P�Ғ+F���f�u�'Ux��)��I��Fu�!ѼI䊮����qp7+�VԮ�t)R��b��b�Q͡>����
5��ޗ�֍����mw$�	6�з�o���m�Y9��ӄB�mi��ó/5��@�6�5��b/B�]�+��Ggt��ͼ�{B�����WyYۥ��fj�	*�	t��3R�`��w%�l�n0�q��3�{0��,�	���F������ƇWYoU]
�:{��b�YY�G�*�m������`��=�p��#&ֽ�w�^ՠ[M�.�h,���{j_MZ�9�f#D�F�q�w�[Ř`�P�m��}z�$�
�k�N�FwS��Ћz�ꡏ��2����g�La�\�c�;O#\#��;ٕ���`��yQ���
�J�:p���2u�c2�@�q�5��S���ru��b��/m_f�p͹��t��
U�I�U�`իT�16k�m͌`�a����*L���]#�븩H�{Z�l5�Y��'�C*S��P�KX��&v�XmT��VrF��;�I�Cͧ�7+�N��ٴ����UA��J�J�¥H��H�J��
Yb0�T��EQkkT�eE'�q��TFE�T
"őH,FEQb�R��5�DD`�f$�,ְ[j2�Y��Q�%@�UX��dP�UE��V��"��E �cX
`���KKA°UDQbŶ�1b�(�J�Qd��XUb��l�X#�Z�1�bŬ�I�*"T�Cc1R(bJ!Y+(��T�J����1�-H�*�(����U���aY+�YhV*�U��"
)Z(�aX,-�ZX�k����H�TF(���T���EX��Am�UR�((,
�Ab0�@UQH�U��"����E��q��Kh�*�R2ڪ��eYZ��-�[,���ر@�LX��� ��d �WB��f�M����~f�`o��Wj�bq2t�ڦ��cgz^�Ը@�Џ^�V;�.��q3��lK��^�9����jή��)H���[��>�,U��x�Dݪ��픫�U��}iW���	��+�Vt΀���2�uE�:�ۘ�����F�t������BٓIBƁ	��C������z��Ҫ�Fu!{�]�e���T;�ﳙ\1���t������ˊ�fA����<b�&��X��B���b��ٗ~�%pei0��m�F��د9�!�O��*[t��N��YƄ�0�ڐg���\�^���FxV���A!#BI񇐃��lÜ���
ݭ�^5���l{�&<����>�!a['7»�iG7n�A�Џ�f�9�a���V\1-��J�j�GP��P�_r�sZH;���E�xc�`UI�V�td��ؗc�5���>�Z��GAo�	��:r����m���������r��:�����27���;�O@�Vjǅz�h�̻� ��G_a�D]�)������uQc�]m/�i����8�	�^�`s�$g�P�'gyR7���A�qQp ů*�ϐ�۪>JgO�T��5��ݎs�[f����7�����y�yt�x��3+ wK&NF��uǩ�43���#(v��]-��,��x�.��7��4��b+&��p�ƻe:���G�E��\ł��UϳGm0����X����V	N�GV�%�&{Rl�z.��RVg�������*Jѐ>^��,�W�-ԶFNX�Va�2��`{|�Ƙ���-��S���_]n�Q:G�����[�/�M���N����?�}�|�p�n�뇽����y��{ˑ$�Q�3�������kv�Y�"��9I�9[���ڕ���"�>)���a��T�?��k`�l]rT�oj4�@��}�g��	������c��.ӵ�;,�5g��Ԓl�=���K�&�b��3���V�ݹr�Y��`�=�w�k�qtLI�B���}XE]���$�^�?o��`�.c�٧�7���zG�{C�L"�(5��x.��0�B���>p����o9����j��8�X��1V�c`�ȇ1�w��%��W�t��K,%���7���!��B��	�ȳ�x��6������Y��gR��J�{\c,F/�e��K��\k7��Z8S�mK-3����\�*9n���4p��k�>��+��6��\
4myS,$%�=s×��s��~]��'w�:�2䄟,:N#b#��x of_]�û�ޞ���\����0_)��*��
���t| ��U��z��Lݕ�o�(A�~PF�z�%=����L:=6hRT:�=r�J��=D\����9B|.OOb�n�5l<���� ]Cd��LИ�ͽ���7�dGev��3'S/#���4>�XJ���Um ��no���Yw�<���N F�/nt,1�St�n�vTHz����Tl��^�G���i���hu����h��3�yt��@ݾ��47r%_�m��Y�w�To�'[30�9$#�%�d�|gN�p��%��P�Z~_8�Ւg+�L�q����C��\�5g4U>����q��{�����ƀӅW�ܪQ��ϐ�_1q�,���P�>�B�sܗv\��ڶ5Emnps�k���p5����?%�rR���ӔP��t,�|q��z:~�Mw�533sf�^Ý�D&$P۩�e�� n�M��f� ��?���ߎ$+�O=��r�O�hڞ)�4|*�dxS^<I�����NkV���|���M�<�론��cz0�'��.2����R��8�w��r0&6�o�B���+��\4ϱ����0���D]�N�(���7:a�x�����)���`�&��te$h��/�T�t�3��06������^�}b\�����gVU��~
�,2���5��Q��A{eMZ�ᚖ�6��=:|�l��՚X9㊯�<O*�ЖVGR�ֱb����D�K�yDu�&�<8'����zB;oAՋ��Ǽ��"">��9�Y�B���r.t��V�=�������1��Y�q���\�3����r[��Se��<5���J_S���t�q�����u~���n���ʥ3�j��U��i7қ���,%i����gv�Z�n*u�`���m������X�ϗް��Gj�UP�O5~�!��m�
�4!��u�����1	:Y�ÿ+9C=��� \�6f��������yx;�����e��46~��za��I{4�w]����P���8�����-�ܗus�W�;2D:���[ ���.0�)+��t�1L�B�Ӌɱ��r� s�19xÍ�x]�G�'�����<�&.�,
{9֘?=lş��y�8��(p�B�~��ᒰT�Pò�\!���2�Z1�U��zJ�ʼ,C�j}��]]�.�v��խS��5W�a\�|�{��yj�1��&B�	���F��4����&ܗ�:��]˪��d��8_��gg:壜���d��ã���|4Ѹ]N��u�܎����X,*fwΜkGo��F\��x-����`im��Y�%�r��Ϧ�"�ujvw�ݮ��/��ok0�L�Nc��2[��'��y^
E�^�kgu��q��g[��\����sH����0��ٜT��W���"�E*W ���{�ӏ��n��M��T�}�u���}_UDm�����.����vWP�0�iɕ��>�k����.�x���Z"x���VBq���s���9�\Roj��0S�Wx.䏭wn煗�Y5�D�U2wonҫJ
�Z��Η��<.R^d����ǥU�x�a��R�j�k��ޭHM����,�.�{�����x��}>�WgGP`��n��>��l>
�_�ޮ{�;�h�A;�˝��އM+���aw�@~�.5���lwe�½��p�'g��^g��,�&�U���96]D�^��퉮��{�Z��k'�xz{#��B0�Hu3uP�
c=�ܴ���-�,\�ʧ��Yw�9Q�#�Ȯ��t�[�:U��$�����/]p����s\Λ�v���oϝ}��2���a1�+h�t9x3�#S�;6���| .�*��n�F���d�+	�l�tT��]��@�7����;ldN�9��ԑYF.��Qχ�	�[�8c��[t�Q"��No��ޣAG4<�臾������{s-d���uf	3�+d��cV�
�GR,�ȧ*xo5.�H��ý�X�u�oz�#�P�b�V#N;�42;4V;R+�A�,^�s��Y�r�X��Z�v�"�u�%u-�(�*�Zy�����{ky^Ͷr^TAṙ.*����|a|�d�@K�JKT���>�w���k��C��eo.����8�� �P ��=�A-嶭F8���Z�uy]��a٤�o�ؾ�Y�L�x��s'{�[��_t��gi�F��q5���e,�F�Y>�Zz�O�ϩrY�_w=է�mY�1,�#�gfQǙ`�Q� .5�>�U�7�l�
'Ըf���^��t���L_�����՚���qI k�Y�_�/hތ�͡�Oz7hP��W�1�dy�x���|��U���2�3D6�e�����\;��˺���>ኊI��nX	�0�ƌ;^����k:���3��w�$]�y���-�Ύ�{�^E�	(���Wp�1�V�L򦦠mC��R���"��u����7S�]���&.e�-��R�T�[^kM��8�����R��Re�R������CRV>qr��
�<��O������v.W�'�:N�����pr���M�|M{�:�f�'��}�­�5�2���}]����o xR�ڜe����v��|,�䲲�����F�a;����cF�c����ڟr$g�����"������tT�\{�*�� ��/�Y׼3�����7+!7[����zrܳ��Ӵ��y�`���/&�H�Ry��8���iukv��n�''3Y��㡥8�cF=�V��"�����着��K����z��3�Ul�tl)W�����'�#Q������;�h[�|�k66��S.�F�~�Z�</��v"Q��:V��3_A�a�B��	�n̹���'�.�i��C�|{)�^�Et�!T&G��gP�={Fwr�瑜.I�#m_V�u6���k���mo��r�F��6�Gw	9c�1Ш(`�Y�X�Pj���/j�����ӎ2�;o���a(�HI`O[.�M�p[��m2~BNMI\d��wy��S	�W��ϔDR����%����A�f��q��|J�L��3��iU���g���ܛi�P^�(:]i3,�6����[�bS�<9iNv�=��d��f	�<]ngIe�Eoh�F9�b�9���{��\���Jx��y����U�N��Yh]����aQ9�4=�E�K���~/�F��6�����j��d*�>K=�.���.��v�grG�*���V�ɘ 
q#���.:�O]�Y�xjF��ȵ2��}Dbwn���C���d��]2�j�7����*mI�	����%������l�����qj�-�g�%W��m-��E���w�kh)�Ȼ������^�x)�ۯdlE��oZ��Lk�n���e� �ӝ{� �xS{��m����&J�d�oE�⊎¢���������l��,L�o��M�T/�bz��ypW#;K���S���nm���H_^��ۚ�Q8^)��E�����CioÍ���8�j�^��q�ک;#{E_ry]���r�%G�)_�S���t�˞�Aܗ�jgP�_�~!w�,�i��Ύ��,,���ҿ�>��}��r��I���A� ��P5}t����U���n7�ϝ>{-���S{q�+�f8��
R�:�.��Z�]��Jo{�[=P�|ʚF>�.1:LFR� ѫGs���>�++�k��u;��es��z��	��t����l\�ܢn����GH]{�=�kjⲍ�)����.؂�V�&P/�
t����:���!hڡ�o���5���[l_�s�z3^�ٕ`���Q��=B���-�aw,��&l��C1�# PH�v��g�,�̄*��BV"6B�#Tg�>���#�#��q�;yW��_%�	V����Į�s��z��.�3q0��G�t�vY�y�le���g�	w��T��δ���/�;��P�}�P�o{��z�L��>0[s|�@yp٘�X鰻/�kn�NkB(
=̙�]�4�7�wd�Q��rN�=P��D��0Ӟ����k$�N�1C�*r�N�aq���=��c�\����%l6����� D��O!xگW�uV�897�e۞���QI_��ڶF�{��~�/���{.�1m��.���eP���M�����k'��;��e�/h���x�����inUI���Ά���1�;I�s��X}����>ū�{���+�r9����ᷴ��\���>�V�Y�w'k�ә*�|k�ܣ4�_[�gzV���p7#�N��n^7����6{u���3�p����={���tZ^��*��-��J��Aɡ��{�rg���7مe%�k7_]:����ۃ�+��GY��T�<KȮVN���h`���kq��Z7h\u��B��i��7b�˙�)���o�w�7�\ k�o㾶+g!�&�A�w���}�s�J��y/n��9�R���s~Y5;����5�����w�qx�R)�5�Q�3É�z����s"��\V���+#�+m3O��Cxq�ݑ�t��=U��o��6\[�*9i�4�)�8-62[�98�d�t�{'}��w��<q�z �V�wyRP!a|��-��]�0f���2i���w��n��uͭ@���]��Z�D�U�w7�ڎ8�f�1��O$dH�w��V۪V
=}�g>�ڭc�p[n��Mt��c�VY������HoyQ9����<����2ga�%,Ζ�K�}l�ʞ-�"�q�K=��񾓨����_�Qz�����u�R�g��=�`렦�7�	�+i���y�nv!����c׿	����֬�Ά�͌���U��v�sA��4�[�Xb�0�_�X�i�a��lZ����W�.V#�eUq�������-20v�[����b������!������XȓCm����Ր���̒ΠP��[�g}+��?���rY��6:m`@�����T��\�܀n�7�+��v[�Gi��Nӷ�	�bĐU�7n�`�cm*����O�ɕ�M多���T�������7`ZrM	����F|3�yj+Y�g
��]������(K&8���ځJ�$��WH��]o����LrbJe\�mDz��\j��Y�Ӧ��;v7�C-�я��V��%��i�ۥ��#��O�tȆ���{*;�)�ܹ���\�%\z �!�ӂq�:S���ݨ���mR�S-rj�f��R�M��m�?3\��E9RW\�e���=ʠ�qWxkˠɚ���I�^��R]�T�K;\S�
��ےJu �^#]7JWv�T6��i�fѸ�މT��ב��-�oB�׹W4�2��n>�v�_u.<�@�	g6��ݫO��f��e^&AĠ�Lm�ҫ�xAW��Υ")�w{�;��p���nSk�fr�j��#�G��i�W��c	�X.my�Qzm#[[��Y�wm������ �%�)��eYQv�0�W��(����.���3w!R�hWB�]Ǹù���Oh`MU��\
{��!mNY���e򶜦���c�v`gm%DK&J匃5T1��J=�.��]p�ju�,���R)���J�gr���������X:\�˽膀m`�a[����\	U�a5�J�[feb2Z��}�r�H��}9�ݾ��iN�P��n�[�)F�<grf��-imv�qm�.A�����Q�f�j̗�I�]��0k�W7�K�NĀX����k���B;��#ը���:��(�%Ȯ�Y��`�š|��f}��=m��\k�������������&([��Ӳ^��~#����e�v���in++4��E�Vs�m�S����ǚ��S�s�����Y�㍕�����<0V�Ȫ�3w�3}�Ui���6�'g'9�G.��Y��S�K"k��հ�0k:�	����wBPr�Y=���Rm˱vq._d��H��psh��;�4<���A��Ք��8����
;�Ѭ+C	�6����]o��	\�`V7�BlF+P�.���g:��� ��*�n�p�W&��v��i1����e݌(ҳ>!J6)=�$�-9z�.}�̷j�{�G7Nݺ��6n&��{$B���NJZ]�{�*3KM:�r���,��+�P>�j��}���LT�Gl��ֹ�o"D-*gMʽz�<���+#��.�&�b�<q��ŽZ���]a�8�՜��Ս��e�%��F�=X��	��!����������gZ}/+��Ǎ�h����BA���� �\=���!��{7��})��hv��e��5t{5S�;�J�+����gI�Ѩ�-gDJ�-���򾡲���O_AƟU���}6M�ЪbS="�+Q���3����_}��zv� ���J���UQ��R,�b�Db"ʃe%cj�
")KXU�)�T��6ر`�Ab�( VU����
��E��P"�P��
��\�"�Q"ʩ
�ʄ����T�`�T(�J�P����`�����ITAVڰ�T�6��T
�01�J�)���R��PX,X��Ģ�A���c[mdE�b�(��W,�b2�-�J�Z�Tm�`�h���X�AaDPeEF(#�E+"��T
��"�F�eJ�
PE
�e��Y2�PRa�mZ¤��*d��y�]}�@:U�0��H�+�C��{�]rڊ���κ�ykcT��]ы��^���*WS��K���I
��������+F��'�av�{R�(^S�8���;C�л�R����+��ٴ�X���p�[�n4��|�����1C�t�AU����:-�����R��Ь�p���
�Fe������*;-9)������4�Ka��z���Zh^���^�v�G՞$&�{���mWM�i>�9й���=��L Tj�#{e�+/ze��8��r��Z�1�qˠj���(z�c��1�L��QԙD����n��V�m�5�=���t��(�k �L��L��܈��gn�W��d��$ϩ��6��͛�2XZpg[��Ƈ�I�2�8[�����iw9�s:-��F85��L�wvD���/F�lf������U�I�;�N4�n��Ԟ�w"���������	�p,#1��ي�G,7Z��(�M���*:(������LD�d���{��}�<�Gm3j����s��������q����+"�ūQ�m��.١��ھ��@Q�,N���FfY��:+ 1bKC����%L�w[�T���y�c�[N��0ud���n���GNH��0�[�qht�F+�yX�C���s �-�ri������ɫ��}�V��P�K��7���r����V����Lƴ1�>n�eWG[<�r����w"x+�W��P���':҄R�����Ҏ�Nu5aV��j"6�Y�V�/�GP�q��f):n쿅��>�؂\���\�Jw��~������^��3�1Oa��o _\ȈM�d�ɥ���2I}Fʸ������z�m�k�Jm@ƍ>��gn{�t�7?�#X�7��+=ۊ�vޭ�_^(��3MX]8�mD5G��nt��;��,�Rb�����6��>�&w�iX�yz�TG�v^��Ad>�'zu�3�V	E�%���.��U��l�u�}w�5�q��nT�ܱ
��&�լ�r�|󸷝���-�'���!{B�����Bc$=�5%��I��_�Nu�w����Ǔ~Bo�ܗ�mgP������mf�;�#���
1�nrΨ��Tj�UO� �U��pp�w������s��HwYÛx՚��<��,�J�.��Wol�Cs�Z�u
��tO�ُZs]�\�w+k(����yK3���\/�)�A�v�v'Y Em8x�8
��z2������c�Y�J�'(�n����1�����[{p�b���>9���kF�����
���-��}�3=�iz�g��v�4rbl����$d.��Ps��t����<�-��^��6�q��۠Ņ�,OU݈j�.UO+;f�S��a���H0e.���x�{��{�)ۿu>��y[�pZ�9/��[4���f�J������]����CÑ�S�΢/"��{����T�����Z��X�U�fj�Qq˶���M-yqN�7TZ�wk*�x�n9>r��|��ypٔC�������30��r�`Uwx��Y��ٛ_ܮr㓶a�g�{+���^�9��	`��������ps:��Q�լ��9\�@��=���Sѯ�'����/|�,~��l����+8��l��N�%��p�gz]���7�A�:4�. ��.,��Ջ��j�4࢒:�˷z�i�� /�$��B��=6�$+�1谺�Q����#�2(��YB?=9-�yt���ܳ���̭6jT~q�C/��׋��((�`��(�VR�CU�'�G��!���M��.c�n��,ɸ��,���|}��V\b������� =�����w�(��b}�V�u�Nv'�����s�C���P���Hњ����t��1���m�nn��f���b#w��\_�F��;�r'�/v�aa֜Vۇ�:�1F;�S�?wsr^��)���q��M�I�s�:���-�_���y����ϋ�qc���#:��%��ۑm�£طzR��v9AP��^i��Ó�`:�.�qN+Z�9"�f9��l�sM-���w�grh�&�S�<2�:��[�=�Z3�N>�4K�����T5T�C��o,�gGf��um�XK��tf��̚}:x��J�\��lû%���Iƥd8�uί�NWܾKtWQyې#�5�0������d�6� �������Kᒇ��yG�������F�n�z�T�h
k?^	�\��V)o��s��2����M��ᔐ�v��]"��v�կ�����ԝـ`\��sz^ܰ�3�Բ�Bkp���Z��:Ǜ(�=��ˌ %��!�P�840��7snL5�?���=Byv(h@>�Jku|O}�;����h����*b�w/����ݨ�p6x���/�-�SKr��1�e�s�	������.�TO,ը�o��X�x��t*c��u����6[�Fk�F��ӭ6� ����5�g���ٖ����iv�q�����t;��P+�w�#�I�v^Q�V���j�h�to�96�wǲ ��*f��'ԯ�aL��Cju����M�W�R�~���D�n��q���4�U��kÎ#���sc��+�ӓ	��<�o��йj�uewtB�)�nv�'70�u�xk��F(�.���JL,[���J:7Y��YΥ����o�>X�L�Xfv��u��VF;�#U��Yn����9��L��J^��c�z�����,-3NXp!Y��gh�S�;��v+�OE(-��3���7�6b��nN�&ѝ�E���vZ�F���ӬQ���SM�6��4`�"�Ҷ�{aR���-��CJ�BSo�62��g(d��j!�Ԗn�A^]��R�޺ι�0H
�H�
��4��/�_W��ߞr�����oai��Ȇ��wa���W�65�oU�:�uf�v����([��TBO���Y�gComU�af�US��m��<�q1��2�=��/s�V�����g�{[�6��}=�b;\m�n�0��N����Y��Ĉ1e�:�����|����'�p�l��X�^��Xe�gp׮��Q��)�sQ]|���ĭf�<��iT�绒k��y�uW���J���2̵"����og	g������]�+�&����U�~�ar�̝�l��8{�6����T"�M��\��6��k��x�PEyT��ennwt\���o91v��Ҍ54'��=���r��U�3S�[��W#h���EGkw������Sq=q	SSbL=���e,�����1ͪ��=�Q�z�Vv��cv��ѩ�8^�S��4�o�9!ͼ����Ϸ[|�#�Ts��X�r��9qd��J��pȭ�5�#��d@�-�1��#`l����.ӱ�;v�/�Y�{�H)�bSb#kw�v���ϓ �7la�����]q�u;��lލ@t��d59<m�Ll�s{^w[N�����z���=���v�6e��l�Vr��q=�P"8ڋ��]$əoPJ'����i�P�Vk�n*��I��̸��b6k:����S��9�?���^�ήk	�񅶫�&��ͪ^A�6��8�ܞ�8��ǘ>Pr,�r�#��8Z��Fϗ777�!���XbͲg��3�J��(Em��זs���o�b2��iZ8a�m�ܶ��T{
x��w�#$U��ܛn���YZ�g�k��|�:|�h��>׋�!��TN������ ~�~w�W��J�-��Aɦ���0�z�z�#e����b!�����af������?�oqt�U���/�Z]<����L�/�pY.n��%���6�P���\��3.!M��Y���V�;j��~|���.�y��������up�s{=�ƫ��1H����Wҙ��n�J�޸��w�vO����|.�yvs=�e��WB�J9q+��9�Ϭ�x�/���H*�]n{���H9�3p��N���^��I����}y���8[ō<$�iTư�z%�{.�J��ܒ���<2Pb��iT�4�W�����r��;��w���za5��,�l#��|�7�]�m�gk���ȫP�+p�i�Vc{�#�ˎW9q����nhJ�SE끸�@!�(��ʣS�%��9���Q�����b2����ܠyΠ������'�vV���"��x���ps�Ƿ�d^'��.9e.a��1��0����X���3h�<d�ߚXCYc����1{C��3���h\�����9�73"��.�q�!�<��g���~��qI��k4ַ�<�M���{�����Nm�[&ݷ��9�L���"/ޤ��.B���W訌ј�Y�1�-N���/��Wq��=^�s�]�׽��TLS�-�>�ܞ�7��]��*bڥ;���F���չK#c�;tz
*�ԩ�א:�x](V�drG嶙�|Ά��F��͋���k�_�:wԅ70]�e�O�`nNj�9h�dG�d۬�Y��0��cjr���B\���0+|z�f-ۋ�!{��`���X�\�fG)\���E\W6&�s�,�b�_3�zL}8]��!�}��R�nM�ʨ����Cn�`onz-=�E^�ij���lk��QI9�K�5���'�sU�5��]2���������[p��3�I�D��ͯ�1&���^��q_������+��u�=�|�F5�j8�*���c�%_L$���0o�eA)='^w2q�8t��D�&��ƨ\s����p�=��L����v �d�o}�1���z�oW��KQ����ɶ�t��ڞ��k(f^���9g�N��c��L?��9��&Ӑ��A���"Q�����d_��j�K�����w?��V�dB�:l5��'���b�]��<���P���.�ؚs}%�h]����*w�&�i�a�Ů��� ��}��Z���{�>
�\��<�eW��O�5�R4����Z�^��b���7��{����ܬ��jEDaQ]Ų�b鞥+��mw�[O�ӂ_<�kp����m��=d&���#2l3� ���V����d�"r$�5�rl�B}8&$�9ZO�V�~�ޛ�n����ΏQ���Ύx�8J��Z����ֺ�[r�(�Q�(��;�f�44��k��2cC������7�N���Ʋ�jp����^sX��^���f��pr��F;�ꊎ�)�7�I��S՝}jrH�F�����J��ଋP����^_�P��p��>{�.�����u�r\���+R@[�_�;�໷__���m����3Բ3(;.9\W��'��e�9�]�\�5-��z�5���^�[���XZ�Ӕ�_
Ε�����b��OP���*���Y/�6�u7���Q��6���+����&ϚI͹�{AZ�پ��jܼ�w�S�qa�t�n6�al����B��7n�[�WГ�u���ذ+��r�%�L:���{�%��q���l�P^e\����q�s�g`��'a�������J��Wv��7���p.��:��m-˗�l��=C:����)�K"I�k:��6��c��J�,R�EA���L�ڝÏ�gc��vy<�ř��Ht��N�Ga*%<�UW������M�q�׾��ni��.���O��tX@7�g�j��c[��H>F]��|B�����R�VV�;�y/��r#�ɭ��g`�65�J����%#2��.�9F�.�[�p�wo5q�C���bT�a����g$,��km�����(n鼪�ݩ�q�kmЦc.�:�4p�s�s�!v��:���H��/t�kc{}t0�icu�0�Ѷ�H�|�U�H�-��u�p$�GXħ�6�gC�΄�]����a��0�F2�VH�7�����I����8ui�t�Qqڍ�)�\�Q]}1�9�Hv��r�U�<�s��]6���(�g��Z�[�h,�e	Xz��v�wW��}���c6�5wuƳ�J�1��iF���L���'�mF9҉
�I$j�u�����^ͣ�ǯ{�Ғ�����u�������Ʃ,�S����.��Ot��X����P ����wE�e�����BM�F0�9����s�bN�fԄ�n�kƞ���v2_���6��ƾt>�G�C�.��P�":x�X<�h��h�Չ)9��p=�At�¤YCZ1_R�F�.�#�9+u��o�]�&�a8:R����i��=(��ʶ�>֫;(k��׵�r����ݸ�a:BX��u��:}��p��k�Y�+���!ڏ*��q���P=�<o���n��F#n(��So�������ź��zew��s���@�����+��/�N��S����u,�;
��knc� ���nRe�tl�2Iopei;v*����v6�|�"�o�7Ԟ��]jΌ�6�ηN�E(HadƑ��ݳ4U^T���{X��wx^�1@g��2�d��]J�9f=��W����u,�֠p�����XzU�6{Hr����H�u�s\�Oj��ʏ�Q�w���0ek�P+Y�d���l���n�q��y��м�ܝ3eM�[����U1�g�գX�b��kO���9�}&X����۳�	��~I�����`�͕22ѫ��JU�e7�����Ϧж�}�]�\�Rmw���>�[����S�=J&N'1�F
@�������c�:���>A�[�;���s\޽5݆aɽnf���8X���y��p1ע�T�ֻB,�����
B��œB�����p��jkX��.�xi�`�`ַ~x�C4^��}y��ť�@p���j���$��ύ�b���3U�mt�5�4�Q�K6�ȟ6��cLX�rݍ��ݼo4b�O���"�=�a&GH�S�i��׊�ٜZR�nW[࡚���e�r+@>�R�����˼��(8+���;�nl�o�.it����[/����˴�WMX(���4oW��lzd"�ޫ�������Ҳ��l0�S����a��XE`!��Z�0��[���Z�-R���!kk*�1�}]�$�:��>p'�wt����r�ٚ���ӱ�����w�߿^���|����*�q!YP�PPU�����L��9F��k(�N%[d�T�@P�Jʢ��dD"�
��f!�B�a��TXi
ԅBc*(�����*�fX��(�� �"B�*!YQX
�-q(L`�R�8�*J1T(�2ت,�$��.�&j�B`�dD��X,5hk$��eKK%Q �-(��i���ő`�hTX$Y���S5���Y+X6��L�ă���B���4�2
A�Z�*�LHfPZ����+�� �K�V��E& ��(�

�Z��XTjE�r¹mI�c �6� ��1�La*-b��
�f&�8�հR�
!�*"@Y1�%aJYYEE�
"AH���� ���wsY��ut�P����l+�������}EK�]5��X�P��ut�F{Hǥ�̇.�:er���&VLG*����z�b��>��s6s�拊LJ��يE�4��s,{�^�ZyCp�k�^��g���զ"ZˎW&�1w	�}(��B��4�_f�״�]��x�#8Vj��B�pw��X�EGj|�^�W�z�q����H��pU�	�Ab`9/��[�X�NjӘ��o�f�#wSy���1�c&
��¬)=���f��Ƭk�l�趂�|�|V-]�6��ȏV���l�1��f.���>*O��:E4��-����ֻQ�6����^���MZ����,8�@~X5An���:i{�ɭ����=W�m�̸��W:�X��uT�#[{v甔ͶWk:��cv05������r"��efƼr_m�OY��G�_GV���5�&��*�tm+G������|���x	/.����]kX�z�T���������|�Ο3����ɽ��[�>yo��~��5k��u��X�08w���O��O�XE���AK�.�ಯ\\����*�<�s�VSn��X��D��H[�O;{���>-�E_9�3��ڬ�)C��3�^*�2]xk�]�1}ԍsg�J��zH�p����dvf&��Zq�j������c���fѯ�Om�uS��(1It�g5��ԋ�aU4��
����Y�̜c]�+�����G|��#c8$��7�2i��~g�X�ˆMZ������N����lw�:�9�$��	�l��Q-�'�%Ns��X�:�^4��C.!�4��R��~�:v+;��S˴֩l�Z�i찖��q��{0�yɭ������_�G^���hP��������9�/�/K��mR��5-s���w�_ϡ��7�1
́syn��;�F��n�e�fK��i�θ/EF,uk��n{/�{:\�@��W��#Z��P�~`�����+N@�g
ӏoVȨ�O&cf�ш�w[��oz�Z�!8��u+�xɿ�>X`5��������t{�k�̵�_'�.&�_t8��f�]9�^��Bx3��؀�."'e0\"���B��n�7e��V+���ʃ;����tu��2�]��gq�V�(g�0��tү���M��[�%�Zzn����ڒ��m�(kL�s��e�i.!�7�:X�Kb�jfkZMh?�i,�}��+e@��}����Nl��/�@T�iؕ�&��u3H��/��zd�vg�����*R��ϩa���V�w�=�K���8���dރ=[o�P����$b�1X��:�Z��<ou^f�{y��==om����j-�xxk�-������֬�W ���f���R�x���ˮ��?*��N��m��vD���/�Z����L�S�LR&.&R��@\�9o9����ڏ�җ�`Π�rq���7�j-?I�K�$6)��7yG8�N�{ɮl�Z�7Sһ����t�I�q��-E���p�3W/wV�����ri��j?c��m#��1	^Fْ\LP�@P�Ǎ^gO�� �US܉�̘���ZB^�wɽR��:�2*@�9�1rsq��#n���=��'W�)k�n�Jm�>�>����kK��ɍ<�A�;��[�3Ŏ�ק�.ܠ��\Ps-���.���cɽR�!v)w1��]���^��»����i���({�֙��AX��<W=]�z
c�G��r��G
a�n�|%�K-D����,>��9��nވ/8�e�F=:"1} U��A�[�x��U7�4_s�x����!t;3_Zs�pd��3�o.^̺*�<��m��G����Qb�^�=�L�6����Оi�a��lZ�9�j�h������;T�(�EDv��K<�U�5��yl�A��L񸀻�\M{9�<��Z�֊�T���V-�:�R=}��7X�x����O[�۩���W}�3(/��]l{��]���Θ�J�q��Q_vZr~OWO<òJ��Υێ��ԯ���o}�������(C���������]�1&�� ���5�eOd=��s~����/ ��n+�'��my�>�Э{*�x�����N�Z��qk���8�V��d��_ӡEkQ�of1M�|���׫��&�����ҹ��|u�M-�P��+�u���:5ϦLާ� ؆c�Tp
���7{T}=�,���3��8�n�M�-��!ouB�*��v7�v*g�y�ܫYC�Ɨ��w4��`Z�?H��B�b�wlUf�$޷p��84�Ԭv�kk'Y{�Q���߱���s����2�ڤS��9�%��.c��I��c7���5���C�v�w���8 M嬗��T}5��y[�h�sVm��ҧ�بD�,q�����g�O��iq��ӆ+7Z���2��������;=@�������oza�Y�)۵��r����d�*juҮ]S�8ҍ�m�r�4��HH��l�� fݍ��=��0Z�t��W;T'*����=(�7
����7h!9֔�]ɖ�~�<���9%��iO]�Cr�';i���0B���R,t�]�֑;x��l�j1��Usn4�9����ɋ�OT5/"ul�Nx��N���R��5<�-�q��Çv ��Fv�|�]�Υ&�s~j߭�b�w��SY^�E��i��=�w'�W{�dVb��m����ژΥ~jR�n�o;���n������-r�t{m�o���rջ�ay}Cv�� Ӂ]�)��]�*�Ǔv_�g������nJ��5�q���ʹ�u�m�$GLn���åu��;�eԚ0nP�nG��-��Il��\y3m=�6q�[O�lQ���<���B�貦�:��뜝I�����)>�ɺD���y&����WF��M��;t�#�����ή=t:����1J�埢!��T���c��퍼Tܻ�;�}�Լ�ߡ������d���^1l�铗>���.4=����ܛ���R�P�-:�u�3ݠ)Z����/5��Υt�oF�㈭��[�dcg.�hT����4����n��$�)��7U�9���#����V�TA;�c+�����<1�;u��J����$�'6���ww�6�f%�B���@�K��G�l�����UU�$.s�LǨ�7Jj�]Q�=���$?U�
���ʫ��ѓ�<��U֑~�`��I�]3UН�_N9�����Tb��R�]$�BZu�M��P-���ݧ���N��Ua�3p�{���o�vT���g\x�۲�sZ-����Շ�]�~��6�5b�}�Xf:�l��cEV>B�F�շ�#���7��z�tY�.�g�9mN�[��0��N9�qxM�:�M�H���g�o:��p#XoB���\%��v-��)M��)w(�埲��2�'xP���(�.�y�VWK�q)�yak���X]u�펜���hv�+�x�����\�v�C��k�\{)\�{:����>2<,��o.���D"eD���6�,���>�>|����?3)��4[��w���JS~��2�r�o�<��n���*����=7�i�4�4����jlI��x�[����Wq�ƭ���CzFAQ�o]�sۏp��
;e|Ѵ~�2o��,?����q�v�K���,��л]m��g��p"���u��+ݿ�Ϋ��y���Ax(3=
u�T���wu�e慗��q����Nz�a�ۍg����W�:�d�w*q���᪸��{xy_R�.xb�w!ssq���ճ:ӊGB���ې���Ŷy�2��3�<=j��Vo���R��W��i�kܒW��<�c����=��ݑ=+ttR�Z���[i�=�aݽo�m.�P-s������������`��@r֌��rq̱��J����e�#C���F1��1}3��Jl"G����k�X��ʸ� ����m�+V��$���^A��jՌCړ��~�c���r����k���ԍ��(�K<�r�ٴ�۝ڽ��\��B|�'u˗9��Vt��3R��O�2��)]4��a��Ι�8�w�4s���W3�Ҁ �����芰zW��O��۽���M̪�l�r\�kq7-�W�a}}8r�T1�(q��D��\n�})���15q�.��t�q�񃆲����E+���a�v�&�/�҃���6�n΃�����Yi�!�m������T��q��3,؋��
n��̷`\��j���=��sp�ѬiR�&K����,��Ț��_�����;��#V��Jp�?��w8��چ��X����\���7&��C��f|�ϣ��F<�Q���%��u*����=� �>��
��U̺ypz<ed۪܃Z�{�g+/�XTTw�5x�u�x��r�4Fʅ�f��։��5K���c7곕���:����NJz�HK��ؼ���ess9��	8厱r8�f�C�H\���.��]1,�9�A�-�o�>��J�[���=��5(�ڏ%//DY&��:G��v37�	�(���wϡr�=�"����k�=��S�yi?0^h6�A��Я�O����S����y93^��)vtDv:�S�M���չ: �^������.�r�"��(�k��)xƽ�MŴ8���ΏZ�#���ە�!�w��)��FHU�Ԟ)���ލx��Ǜ��KZ�r�p{ۖ�vY���<U��~�i����am�����T�nGf.?d�&Z��H�m�i��i���`E-sg�YA�4�:��bo6:�f�ͬ��Y0ѭvǀ'����[�.(��\���T"��9��>��3�R���vq�Qo Ϸ�T�`\8�t`���z�;����L:�^����1��4�e{���x���4k醶Бֶ���۾&Z˯A��G��b�jS(���V�0����¸���(t��p!:��L�����8Pq��5�}���|��i4h��<�p��:n�rWK�<����t�L\{������_`�X��<��\����j��Ƶ�2�[-n,w�!-z�N�:S�bJ��{e���3����R8=6:�/��W*�/i�*��ОX�}�l�f��4/r�Ca�w��}��rq��7���Yʑ]l2��M��uar][խ[|&Ä͆��-���b�Qr�e%��2�L���JCtK��6qg�Z�9���7�]�^��zigF���ZE�<�
9
�����3,���\�g1y��Sp=����a��F��/���B�c���4����^��+��z^���m.�7*�h��էՒ"f��;�^N'F�ϥ�feW>SO+9Q�[C��b7�����X(��m��픾9X`����7=��۸�u�z���9��;̪SHZ��YG1�3��sڻo��x���x~���5��q�놖\g�嵷9��g>���{p�˱݅c�V��H�&j���_�}��[�����,��fᮼޢ��6g����mXZ�����J+z�^�_gF�q��$	�n�[�V72x6�l�.#�������Y_A���_8�M5��s���y7.��;PԮ�ֿ�$�����Rvٞ�����%̓&��9�f��ۮ��^�M�.B���з1� ��/��י;���ڨ\�nv]�D�u�(Lo�ӝx��%4�N��#D���^�m�};�m�Q��]_ج�nY���n�خ�����~*�ѳ;X�B�qK��k�J+a�TH�iW*E�vE�/(�)L����-[��l���|�_G�^��u��=��z����ͼ�-Kz�<r��Vh��̢j%��Tw��f3L�j�p!K[ø�f��е��U�te�źY۽
�r�g��r.�e���  ��f�MԭUz�������e�ˎ�u /��Ƹ,w�Ԭ�r�M�K���+��V��㭐q��p�A"�q�h�Iv��u(�N6V��^V�8���W��*�vf��~YY/�[}�:�73��q=vr���4+�~��o.��жR0�Sxw^��:3��a��-�S�d|�,�׹�]������G:��0F�2��r�d�����w��1S�LΡ�o.e��S�C�͗{H��X�e�<y(�T�=Db�=0D���n/Y]s��u�g�*qȀ��>�+�ɼ��j�X���'KI��,��Y�@��"�"���9S0���Ɛ�y�$��koM#]�%�gm�W���Ue;]s[8�����=s��@!��)OӬf�W`��������ˏ)��n}�3�`M��u��
�y0�d�h�Ey��C$I��c	��s���R�����+��������r���ҕ�.D�,�,قܽH�"��b�'3(�/1�#�(cyQ�so�[s�_���T��:�h�3ͱf��ݳ~@���tK���r����=���mk������
 �u�ޒ���Se�;;Zn�W������UL�;�z%:�獼�1��f�kA�M��^��K�h�
�� ]�S �;�Fdؕ���2Pߦ�u���0v�k���۩3u�x�S�e݊��DnZz+�z)�ז��u_M�YC���w����ީ��&ꋲҰ�� .�$�W<���Ř���ݜN� B�9�2�y�$�2 �BƮ��������	�G&u�u���7y�ϗJ�]��vZFM�yh�U�c�z�4�U�	e%Au>�z����.U�,�Q�0kOM�լH���_�|�`��t��w[\
�J:Yh�1��|ܭ���Od�u����b�\�Ws�����y��{\M��m��';���>�v{6�\Y`]
���%��0��L��)�0��D�@��d��Nh�:�ժ�}��s�RPX�+#u�*�[����o�P��|�3$}�Mh�1���]8�)��ִ���t(W]���u]��!˫��/B=���>=fH� u�	��T���t�U��b�`�j"���7��7�\��tF��� �k�<{�	�j̥���^���6�#�2);�����[�w@��u���f����ds���Dg/bN͒5��JF�a��79�2a��E�܉oE���UMd�[���{���޻^ڕ����;@�"�b����]Z��(���a*�-���9H�1QdQI���5
�k*Klj[B(V�F)R�b�E�¤P�(�:�IU���H�I1��Lk%UY��*E*VE�Z�`��LIYKE���j*�+E�KE��Ř��[�*�V�(�ea+A�Z��Q�L]\L�Q�۪)(Ա1˧j���d�1
�(�H�1RT2�2�-���%��\a�1��X�`�k*E���2�]2� \`�R�T2�t�DAJ�lղ�J̖�%JֺE�a�5�2��+0�0m-J2�[�r�"�EY
�f�kV1�f����IQAq��Ը����SMj����P�

�P�����r��QAV(�5��U��m�H����|/ 홊�FCKD�r�g��7ϐ��e�\�j�s�n�-�iR��u�ﺠG�[��z3��Ӫ���E^jQ��DSش�:��*�k-���e!��W���Ns��8�iVBt��KlB�;t������k�rJ��9&Ug{�'�s���HK�|����AfQ
�tо���{��?:�<*v�9ϑ�D�A�g{��=���x_�E �{�&�n�M�C�L��q�C��.����.DR���O�_ܮr�;l�P�e*a��k���r��{�K��H�8鯗m�
�P����N�󩽈��e��ӏ9�'�a������;`
�P�Qt'}In\�g1x�h36��e�ո%&�+�,�\�%��}�2��j:�����ˁ��ٌ�ϭ}��ͳS	�:V�u��+1v*/m�	�.��q�ϳ��9��w*�3z�7w�t�%{��&�V[5�p]f(/`֨���ٴ�������O6k����Nݝo��,�3Ǯ�P�1H���cb1�ޭnS��d��6���%*��;M�ۋ����w�]V�畓F���:���'�-���9Hpυz�R���;=�׷���1Џ]x��yP{����d1btХg�:�!5����f�e����=�* ����*�{y`/��nl.7�]Q?]��U1EE���./K�&�roÍ��ٝ]�@�)�y�vh�93Ь�x���m�\��o��U�vD���.��Z�9-�bJ-UȜ��W�-����Ԍho4����T~+TO`��q�moZI�W6�u�L��.g+:�'��U4�����g�ۄt7S��d��3;5��L|a#w�����T#�Wɤc\v��2��H�u]Wǽ�c���ֶ�w�k���uG>��̟�&�P=���A��9@�s:[�3n'�sg(c���;6��u�>��J��<���ڞ�f���v�U�L�k��=7���W����]2�t+�o�g5����'w5�����N�m��&z�4���!�Ᲊ[].ŭ��Ԗj[����aQM}`?�뫇�o��Z�.�mC�8U2a�=���Z��&;ڷ5dYb6�O&M��~���rl�{�'.9L(������	�XF*����
6��͙�E'#J��܆��Ӧi�Z����r����#�ìnb������4��(bW�M��nVc��]v���v������-�-����㿠�
Œ;S��K<̈́a7�S��oc,�9]==�.C��&m?��E.ұo˽a�[h���6Z���ƍ���xhMD�t'��N5`ˆ�r�챈�z�>9K~�Լ��;޶�]?��[��M�ꐑ��gt�֪͛����"��"F,���1F%��*��']�E���]U9�������7�f��j���q��d�����w��B�����nG)�w���)��wm�+q��1�+�j��
A%��=]`���Zy���5�߈~�6v�K��-�����w9����-h�U=�M��X�ԛ��D���������z�oS{���Joz�7q��r�w�%_���Û63�2��/�a�����J��ũQؖ�IT�ap�e7���q�ԙV�A�j禞�<�;ŉ��0�~H(��F�C����8�ʕ0��X��9�5%� +hg[�oj������ٸ�:���+�n�I�6+A[�t�\{xH�:�
���ԍ�o>���K3�f�L�R�>�[�y��W4��ѻѦ�<��_5|�N�BkV���,�xI!i�zq�*M���d�q�ڎn�bBJ..W[;:KZ<����ҷh�%wsx�����0ޢ�qU�B���$YD4�Y�f3�RuS�x\Ova���I��'�����5��*��ɞͷt�8NyqQ��u�̸;#��+���=�Mg1o��{��+�(��lCx�jg,����Ns��ݗ�i���z*0��;6Q��b�7n�Ms�=���s8�6ybu8��_����U	��I���=�&��[�ݍ���[���k�{ᮃ�қ��b޹�+��vҋ4`�p��dS���{����Y��jr��>���ͩ�-��P��]��:��wF�4��5��ʯ�Aw��sy9_-+�ͽ��[K�{��.�x��z6}�A�ܲ߫��db������rnS��r-n�y���\T��x�Q���o��Q3.�۹��k����u�g�����]ٯa+�F,U#/��yw�|�h�P��"uk���%�:�r-�]ff)�>4�7�w�7VR(K��F��]qQtYO�������r��Xt�`S;�N��1��aO����i#	Eq����2݄gn���j�#5�e�U��5��A���n�>4)�ܩ指�Ky��YC���}��Z�\���}9qٔ�]^��;�h����ws&��U|�O�D�NF;��]�l�W����z)��K3\8������aS�Çm�������%|F��65�OgeT�i�F�b���m�����s8�;�t'=���2�fէ���Km�3��E�f�T-oFr��%U��]��Nrw�i�s�b=(��(�sL����[2��Oo����u^�7�}#�Z��N�q9�rk�}l���5t�j�}�f����-��5�5��C�ܟ���Y��/�C���P'���ИC������P��}��W�fZs�-��9�oX�`���%Wm�.�-��ܹi���|B6�MD5nܿ�󳘧m�C'k�zjUi����}}�5�N���W��{����a9H��ģ�cQ~����v*e�˺S�N�VH���e[�p�+T�F���֕Awr�
u0iJ6y�C!�$+���}zJ�5x3H�N�ҸM�xUL�J����ح�z���o�ṛѾ��̯��TB[�d�o�K'��Fx�F���x;�:�֊��&P&u�z��>������R�="�2����Uv
�+������.Y��V��Q��=��el�xy������==�c��m�sy���5�����:�Z܄bՂÙ����C^��Ј��|���1��&�72�mnOe�~!{h5��;�:�>�/L�ܞ�Ns>�~�W��w��U��pub�w�A�S_�7�g�>ݫW ���I^�W'�����\B��cY����ѹ@+�}��������~�lvXw	{�K]��0���C��{Bp�|4���.S���<
�cn�����_^�ݣ���ܚE�c*z&/z@��b5���hR�2ٸἫ�1uу#��w��o{����Jv��/���o���#r�N���\�U�������af�`�:<U�K��u�����f��|��Ǿ[
�R-π�5bBff#�@r�m��8��,4b�&��mwwӲe��ǻ��7wD��*0Ucᡎ��nP�5Xc���yj�[yB��K�oNpF:�/�T��L.ہ��}KY2�0�'p֍�]��+��ܺ���q)!oT����3By�'s���W�X���wp|��9�ז�ܿ�s����ɘ#��țN���-���dr�z4��t�8x�\3؝����e̝���d�:ɜ���n��zC��e0���:Ś�'
�F,�ڞ�|�U�&�v��r�J�E��|F������q�2���\H�d�sG�w[f+jO�3#UY����/K~Z��nm-	�ː�0��7�+�Y����+<=������s�0�w�\�<�̼ڜ��m-���G��jk��Ʀ�N�3����y��YO���sf�p�$�0�W��{.�������jC���nynoQ]�.��F��ɻ��{���V�x8�r^�튇���������.�2�#�����8*�$�wyp!�c�����\Dd ����M]��*�ԣ@��;���(��z�44��p��o��m#Y�/����� B<y*�d��06�l��ةW@C�������r��	l�[YX��*9��u�:�`[�e����;Jь��������_{4�=�9�Y�^Ȕ�Kҥ?����F.��]r �L7�q�;����x��=k���/ݚ���W�+�u�I��f7!E+ t�3���9�^�:㐷��^��bg����K���D�xy��r��x��>�_������V̥F"�W2�Jv04=�~�����;we%3.��W���2�O1�讛�af�_��L�����Q������]a�^������=���[��u��q^�����j}��/$��*~��]�=V�&T�x�2��R�=�辭cg��s:߮5���Q�V[�VW�bQ���Ś�M�Q;�|�����בU����8P�?Q�|r�__VP��zU��ɜe�T�uO�XJ�h���2��%���z8R&��mI�<��7�e�G=}B�d��qs�)��N	�������ߧ�]>�}H.��?i3��u���y�0=��^C9^��G�V[ڃ�ڍ~l�wvR�a���[�i�)lы�٭��T�����)���,~�]ǟ��@}�z\�i8����V�7���ss�Zl`.��̔qi��o/�b���eL|�Ug�_f��M��x�pN���x�8Q�,��l.ݸ�q�m�Z+�5�1��k1;	s��N��R�}�Qs�~�4���Q�2`���1ޠ��r�N���\V�o'3��6���W5>����ݪ�gзBc�;�N�}�b�О��P�7N�}�⒞w~�Nm�蔡�V��r}���
jO��R�T�xƧ��c�x�NG���<z��1��ԧ}4��{����S�[nu�.ܫʽLeV�us���;�s��0%�h�]��t��%W�Y���U��&�u��އ��k�ٓ]���.����9U�z��Q�l�?c����z�����;;��'�+���ߧ�z�㞟]�ʹ����Ru�*{�S�x�cu�	���5�<��ލz/���ў
V����s�?�/߼�T0����s��Ç��+fq
�x}���P>��.��Sa��xw�}[6�|}9�[t��-�S)�MNŷ������_�\��R���ĭz�Ws�lF@���5���n�{)���F�R��,/+̤�c3�GWxG���EF��� zx�W1�����sF+��A��
��z�y��u:��6�e[�����1%��q���s����`�~v�3�$�A��PG.̛�P=�mr�Lҩ�JQJ$����jg�@ᕕ�����n;IÀ�b��^�G�&.���x�����Q�����;����R�v�C����.�J]�ա#��D�; ��F��"}�./���**�6����_�dmWN�M)�u�=!�Y�´b)6�f���^�#����>F�7�*FU68�U����W�o�ll�ݮ.�4U��9��G37˙=c���c=N�}���ϽsBs�?X@�J��.x�m¸>��C�Q��-����{�)��6=��^3p�
��3hg�i1����12���;��S��9�<�t�ܹ�p>�9�ڛ��Wk���y�ϗ�è;�xL<��0'�<��j�����Ee���C۽��S���
��)�f2�oF�zGn[�Ig�=>�k*G�U�{�����'�k�_z�
�W�G�������ۃpi�R~��^���������V����Q�%�������9���o��ߢ��:�\+��e�=�w�^�\fz��X���s>";p�Q���ٹ���U���W��v��J�;=��c2��H�6��c*�ե�/*:lOVm=�Z�e��4��O��Ͻ��i�^�vo� �F��+�Nz@g����˵Gߗꁎz�����ޮ}����f��Z�I����ݣ;���bx�6�:z閨ݺ��[Y����|i��V�'[��n�.q��4WS�1;�A��N�J��k4�v�m��YqQ��p�2�w]bu�*wY%�
�d�vS�m�.>��vu��j�0��S�yVEG�)19��s�F�Ҧl�X�ӆ�^&�J̎�0n�)[m�{��9����4���$�W�}���r��Ӻ��ғ�*�P�Ki�.��@��o��L�2���ػ��!Ɗ]�޼���:)��3�y��6��� ��N���(fL�AQ>U�u�s�Zv�͎���B��&6��;[���B�37v�oR+��$���j���yh�����h�em��vm���e���0s6�p�Gl?���)(�esN���,p�тo�d�ƵI�
u�l��m��EƑ&St���v�SyuQWw\�/�vF�ξ���p�bq��]/�aǛ��2�{�\����I��GW]���
�Jⲥ��(ުK�r�7݄P)5��gM�/A{\u�����yv�d	��UZ���0C��=b�y�a,�cX�!csyea	�a���8�.���|&J�Tsc�,2�*�$ࡣr�p�������/�l�u��؁D;�9�)@q�@�����[԰GL6;�헼�q�7�O������ U��!n����ˉ ��.cEJ��PM֙돰�!e�7�^kֻ5���' ֿ�'>%�A�YE���op��UMV�)n^��db����&�0ZS���k0��'2��t��Τq>��μ�Z#�U��:誅2�H�g��n_:-�0r�t�%�网K��,_\�ϒ�I���
�t�]3����M���s&f��4B���eAnm&�w�գB�Ռ}�+�wyG��^4�� osџ-�g�0�g!�)��Q^F���v�DФDO;�W���u��N��U�ѭ�?��X[c�Q�n�]����Xa��,�ȭ�Bu��c;,�i�y�A���*���`�Y�Őv.b#�n�������M�J��k���My9dgj6N-6�9@
T�"J^ugrFwG�s�ߟn��i_o.�<�2 ���W�L�)
;R�B��=i��ב�e�-S��Gr���Vm��8�+�K��U/�;#�G,c��ɮ'�NٲɸZ<���o6�v�QхT�ɩӮ��R�`<��;G�fл6ѵ���"$��)�͵�VL#�@�3��#P��h��Uw�K��㳧27�uj��dV��E���)Z�Z�1		<�K�5\V�$�inQ2<C�N��];W��{�6��$l&
Wt����jxTfJs��b)w�� �xa3`f��`y�q��e�E�\�p&�G�GX�0]3�s��-M��#Zz�,˗+V�9rԻm��^�熍	�ι�y�B��]�aʶo��n�k��J�Mmb���R�Z�5�W3���&[5�J!YSYL(�j�*�k�J˔�-��2��4m�R�2�6����9P����-�"270�)1�lYPXb(��V�3,���Z�5ln���Xi�"�s)�bT+.P�5u��`j��Y�V���eʒ�ʅ���UV\���mRVV��u�ӡ*ј��h�d�LX ���,0j���3Qf:�"E�+]3)[A*JTD��q���`��f��a�a[q�-��Z�0�-eF"ɈVT�*�4ªD[�EƲ���¶ʚ�c+SE\EEZ�n�������LGT�DqXbcc4����,̤.4Q"��je����
�1.R����
E���׉4�Z�0M��QN��"�6�y�����zm.&hս�c��e�i�6M��ү
��bu�fHZ�z��9h��U��A�mWuzr=����^�[�����}�q\s�s#��Ll�r1ߋ_���N���e�}����R��e�>R<�(�C�ў�>=g�=�!�ֈR=�{��<�dǹޫ�P;�xL���=+
�'�/&_�)�P�<���J�F��7|��g��r=2���Q00�C�b. /Z�� ��gѬ¸yi�ֲ����+.�jfɝݞ>�7څ[\=�[jC��鿏����tadH����S+����� hn��>����Ǻ{8=��b}�}��@^E�h4�#�{���9�"f�X�.*����}bdO�N%�����^�U��g��F��ϽU���q��O�G����yS+��eׂ�b*��=��+��w0ұ�|u���ߡu�W���{^���8Lɍ)ߨ��{��:ء��� Uހ�SY~�G���J�������;^K1���.;��?u���������ό?:����?3K9�#kt�N��7�U
���Bu0�2���kn�F^�9^�~�u��nfw����8{����� 2�d��kN'����]�+:�>ܹNI�ݱ�´r�O��\L��7�9�(.�CRv�ksZ�s'b�u�5
/��4�ϤU���o�1���v��B�l��Tv;�t�t�8��X��;��r����tyc�Q=59lK����)����0?N۷���+3����=�. ha��x3�P�mރ��N��wT��O���ؕ�3/J��1�x���{�����E암4i��9�49&��w��oci�ۃ����˯F���\ǧV����7}��a |���5����d���$v��/����[�dƷx�yU��UoT�\�Y]�3��_�?u��H�.=�Fw��f�iQ57=o�Z�ܼz#�����h�0��V�Vi6���l�y���>���5�_�i��o5-8�f�J�ugc��C�Gx�!��/��*1v�j"��v�#n��������߳f�x�ٺ��b�f|����ˆ��N�<)s(�p�:�u`t�x�\9��۴���C�
��� ȿ����hv��tק�7�gf�����C(0�e�`t�to�sa�R0�c�N�]���[�������+���q�ԐP�p�5�+f��|vs�T�z&e�]P���(�1qD��^�����:�3"C��3U��ǵ�k�W��<�z����.݄�����}F���$�L���2Jܥ�ǒ��a���,����K��_���{��G�"kT歼�U_;r3��:�+w�����5�-�{を���}\/�WC�p\�A��cͨ�*�������\c�\��`��D�����IA�U��O�U	Y�D[�cg�h�B���7��{^�j����Q�~��t���O�T��ݰ;'�|�{6���1Axi�q��������=��Ο��I��g��{��5����=U\T��,���{�[2��ԉo�J@�(�>1{��_P��G��OH�W�}[wrW�:����ʡ�핎����f��n}&=^�"Y��ex�ۆ~ͿpC��S�c�6̥��z��7����2;�'��{�L{ˬ;��T�h?VӜ��z�Ĝ��^�:�����9�n����}U����B��d'}���F����j1f�������F�������fwo����W��ӆ2�B1^��u�﫴9����������_p>X�X�����"�/g�17��ŹθG�&���x˷9��9،��Z�g^D5~̞�^��u��A��ȧ���[�y��9j���<�BٓIA�n��_؍��5��^����dF���^��r؛>�]��g�G�W���}~�0�
��~�jV}SJ�(9J�UÙ���a���n}����g}�%�9��u�N(U�ެX���1��(ne�Y�����X6�t�ń92M]�eY�un��Ϫ>M�%no%ԛJ���ֳ�M���oT��giһQ���ݒ=� @�	�%F.B��|��B�2�s���dz�j���J�rż�%#g�i��FG�������}>�V���+s!Hɞ�/�Ù~��t�e�)�����x3���>������fi�~F=�!�lg���7�����Ӂm�$L��c=մ�:��LN݌��\w�{+n��s��b}bU�G��~-���w��.=��u�s5mf|�V�:�����>������sq /�C��:�,�Z���x)ϟ��t;���j���Uu��
_���6~�ۺ!ǲ�Y<��t����_�`mn!N|~��l)N��UΨ�1�}��4=�ﶲ�B�~�)�fጛ���*FU48	��~>���׶6_��祯D�{շub8��׮g}G��6����<=S>�
�fQ~�"l�X@���"����%�W\�Ĥ�&�E�rq~����~��;���kƈ>�!�O	�95@y�X����,�e�)1vkZ�ͣ~gUB��y����V�WO@�p����'���z�P~�Z��{I�g���vS�b��X=++c9g�b�蠿1[nY���񌭛�c]~�[��R>1�j���^��;�݋�ݝ��ۢ�X����
�]���o0���h bp=�/�Z�d�� %v����}��Q�ߋG�l�Lv���	�r�!_�uD�Ɏ�vp��y^[�M�3su�A�t{|rv<� �r5��F��-f���)L��8]97��*���2����������[p��~���m^���w�3����Q����z2��5Y�+iy��N�9Z���k�{&Mn�,�.����2�៳���w3��[o�����F^���#}�� ��c�W��c�
���;�-N���R��#0�{e��7)�����7��n�
���޻�0���g�J߃]|ap/�ϧ9PAʙ�������ϽU"'1[X������=�q���j�9��o�W���>����W���{��x�n5��Y>�3Dz�ɭ�e��fL���]����n���-�M��Ǜ�9��ߘ���:Z3ޯpu}�̘�����/-�ߡ���}�6�yUz� �@d����J��x�ܯyۓщ�7Z�X�ؕ�|�TyhĪg=��G��Q��%��:[�T#���fF���
g�Y���{劄��s�6[�jC��̹�g���t�ǌH�*f�e�eU͇���F�I�pz��5���q�A0�5�G��f,�{���V_HY���s�D��.ݪNWϪ�w�B��&ϯ���f���^9,�V�Q�.%�W��v�']J�guǏe���ŕ���Q��v�t}ø�MiY T��FnTkaR�e�n8P�M�+�_ZRqK��Pe<��ȸZ�'au�j0jK�r��|�-�HKJ�V�����t�ԋ��(OqWlO��X���+���[~����>�{���P߫�s,��`c�!�i���KvV�G!����'=�bU�Z*o}[�؅=	��f�~�P~��ϕdS��?{��*���� }q59�3�ѽ\�dPHq��q�b2�C1������q������,��˓v��)���vzk�7�e�5�'�,�XE�LV�/��6�����*���
n%>U�w�߇\�oXY�F��޹��{	���1[��@�g�3X����_�ד�@b�y=T֌�����1�c��y�36�o��lxsw�%��g��VJ `��[Nr� �q�;~�y��D̸2sў�:�.g=]ν<cW��>��;��x�C̫���i�e	�g7:e7��j�7푵[9ﲯC1U���k�N���gq?H?y��X���َ���̛�uq3r��ǳ;��ѣ ���Y#��~��]������f�)f:�2�E{�g��{��9릯{�GNNf/9(LTa���P�^#�y�Y�lU!P�
��nf�� ~�	�/M��@w�=7}ޣ�ד�s{�SY�_`��<��U�`	���w�p�a�#>��'�IS��c�抆d�zFJˇmP�gVAY5�֡�T��&���1s|��1����ݲ�r�O�`p%|fT�T�C��nu�5��Y���ԗ'qp�K���Z+xA�����QK�c���;�.z��vC�wVL��E\9���@���3Jr��/�h^g��w9��<�#>�R@�ٯOvk3;7�{���q]�&[���n�§���_dئz�����x=�\�?�D?PC�Ϸ�[7�,ܿUz�R&[�Tm�$���1��T硻��\�dH����߁����#�����>�N�s�D��G��};u �Z��pw����衾b��̫Lw�J��r�:߭�/�֏�2=Yo�OǞ<���{XT��Bu~S'�>́G����4�F������;"U9���f}���.���[^�7<�yӹ��J�}�MH���ېb��i���㗺!���.4=�����K���|�O�zw.iKuT�����`zL�p<�~sA1T紊2�n�5:O�iY�r�A����]^_S����Yۅ�p�a�������C�˸�����`V��{�뽷�����Ѻ�3�;�Y;쭽��1�m9����c���h����,���о�ٜ��M{"��Vǥ�
�FvA���3i�$�o�CN@�SE5���Y�E��Q���@/'sl`�գd�1*4���h+��f� �k
�u�6��;mG�+���E	�su���t��x94�
ݰ�����gp�*��	���`��	����2����R�Eu��ۮnD��^Vl̳F��v��� c��:kmN���9��w�b����&}!�QA�1�x�	�kޅ6{<��Ś��:9
�q�Yz��Mn�,�*�%FU�r~ʭ�5��u�5�3���f�zW��"���f<�[|�o���1�T�Dw��s&�\�n�?�mɌ��=�zL&��۠�����󆇚���^�H�����u�O�;�b�;��iJ�#�b����Ù����&�/��q��[=�G����	��ߑ�g_�f��	xߧeC���.��u3J�t�z�1f�{�R��V%9���B�= ���h��9�#�^���s��hw���9��L3�T�:E�^��tuOL��S+��������nC���=6~OűR����T�����\���M�+s_$Q7�[�W=G���>4x[�R���X������`�%n^*S�N��MR��{l�߼N=�'�6�/~�)�Ӥ�It��?H|���^��h���� 47r�>�,���˜y"��5}��T�2GuZ�e�޽�j#=�n_��T��S/���}{aoE
~~>��u�ш*v+j�`����M�V�d�j���DW���ʀ�e[�ٖؼ��]������z	��
s�;�݀��*Z��V�ZykJfά�q��H��4b,�E��:�o	D֜�>į����U)��'�\v����9��_����y{3+�3bu箐 zVl
2��r)��w[�2H�z�,�N{���������)���׍}�s>@3w�ˠ/�� �y����n��cU���:�8r�W��
��ER�����/a4�3·��dǏ���fL�-OJ��z?��[�[����9[7�ƺ�"�p���������␊y�U=}:�|f��r8�����Yfl�zkD�5��3kn�/��ڽ]Lﳭ̅,���SvXH̄��_�;��@?}_������57��쟖Mn�A��Ȼ���/nz��ά�k�K�����;����oG1�����ûW���mN�G{E�1�A1T�UJ�d�ϵX�����q[�&�_�y��e)^\ɍϓ���u?��;�W�yӱ�Af��(硕QQ9mW����f)�N��E�L�q��^�N>6�3�ώM�p��������x�lY�8�����Nϸ�T8߰����ڀ_����M�T���eZ��^���|�T�H�9�U�.��x:�p873���5�.U���*`ծ��h9���s�"O�`9zxv�X����^��h5��������J5��wI�I���|/!�OCݦ��UBah]x�8�w�U�JD;�����|z��p����ҍPY_A�f��Y]fv��щ�5�ka+�P�Y��j����O	�[~�`6�η!��W�}�nn��͊6�-��z�|{;�gMn��z�r�����tc�2�t�ٻV"�/Z�� 4=�z��W���	�]��S�oз��ɧ�Hc�ڐ�|fzO��L����>u��e�eU�ǹ�#w�)c7^3�������U$;�&��{�\_Rk=c<�ԇ�>���|�MC7n��U9|2���.�&}>�=����S�>�}bk�u�7$67F*���~��1ȟ�Uc��One��Uf����yt2{�|@����On+����Sq�|;!�=�s2c�ν���?xͪb�����["�MM�mUWCu^S�&��À�A�F��G/t3��ֳ��W���_����LӇ�h�YT�����u?e\��˩~S4�����^1{�Ϳp1ޮ�^5+��m�qn�/�{ϣ7��{&g��ڱ���u�C�K�����g>{5��AڦƘ��x��oz��6��^WE�=�k������u��Z]�~�a^1:/ݜnO�轔@р9>���8*��q�\3��)�&9y��\7�uvd��àh��l6ܷ���`+�$�O0@;�ȳ-���y-r���A��'�A�=��.�G�v�Yn�04wl�d�z�����ʱ7����2˲�V��.t|7)X)fбJ�mm�>K��z�<H����V�}�6R�yF�9��(�Ȯ�q�31u[,^d��ڻ:e�7���j��c��z7��Z��}C1t�|U���-���V���͆�Zq�;dߝ���J7�<��It�v�Yo�XZB���*R�3��!9®��� 	.��+���������V��4k�z�m���Z��:Y7ʌ�.	k�H��������k��c� :f�!]���a��,j�uh�%�lż�ӂ�9v�4�F���5uK��I jA�%�t�) �6.�IiIؒfv�"�}�o���\�5���өt�V���*����c���/�!d�ŴLoK��y|w�.�_"�+�:���t��dg�*�"�Nʜ�{�)�
;���x-��R�76�I����H�`6�����A�s���`K����u}�vu
.���u�7A�t��1N��mL��Uv��<q�ѻ��9�~��]���1;�_�\ɇ���;�øw�(I�ȹP�Ӈ �1,��Y�����_�/��tI�A�ٳE50vN��=�m�W�wr*�6l��,�I|�/�+3zeGԞ�|�*W ����!ڴ­�d]c���2��_'����qe:�i�J�Evݭ5:m=��f�*�.L)E��ͩ@�'�y]�����X�����|�iX!]�=;��Ʒ:����]�b|V��Wk��o&ndwI����ܢ35�}%*U���^���r�m�R}[I��:lH�����^��i�˔z�]�p_ ���w]�����{}�Q7�D�B�8]�����b7[�K)�ބ@ژF�B�HgKoH����V�巽�;*�E2wCK�|�:�@�ͫ�Swt����|J�̐g٪n�ҁ�+�ם����[A���r�%��aN}�m��:��[ ߏ[��-����lv�)s�.<r�mw%t�u5�#Vlg�%�k@��b��;g�mzXXw^n��\T���v���`4$������N���$-�w*��iV��C��'7q��FL����,���]��W,�ʮ��X�܊	i�4X5\\�^���Ø2���U�i���f������I`�ŝ���i��U�;���"�M	�U!uh��*�0���kX;o�̊��y��V]���u�:�!����s7.^�C��9�{E������wm��FZ��]3w�7'ц��YI�3(�͜���'n�7�Cs���=���Me�9�¾��J��� s(<�++m|�r��建)*(Z[j���DmZ��DER�����1&&�����Z�Z[�b"9W.`���H����
���
ʅL˅iekM\D�Q����YI����ELq1�s3
Ҕ���,3
��D�L5��̔�d��mBۈ�"�(.!PĬY[-A�P�)��-�JʅKeQJe+�\f�)[�RۙG.fd(�-+�1��,K�1e�.%F�V�[��̊�-h[Dk�J��,Dq)hQ+Qq��CTƵձj
[k\�̴-�c��!�kX�!Q��*�E*j[E�ZP�3ӆ[eV��V�(�5�X����upʡU���q�Ld��`ԭ�*X��3�e�ZQU�Kk,���(����U
Ż�lFS�Yv��:J����%���iH�щ���z�]�����g0��(��C�X�o�E�6��P�ڂ��r���s��~1�즍��ν<cW��>}z�^����M\i��i�G����o0O�Ծ���w�K���1v�`�~ʭ�A�w)�Wz��'��=��;����A���0/=Wgۛ4j$�|7�z�?Bzk����d�7nf�w��_�iXD�uR֊�+{�$�W蕄�����A���~�������Up�aQ��s5��!��{w��Np��}vNx���WS��Ͼ�l���)��z��;6�����%�t�=�p�ۤw��xX
���-CUG���ۀ��?,�ȇ�l�MzWdo�������⭰�ȉ�\�-��{2��Wzxt���w��}�Ӟ3�}#A��1a���p�1��f������������Um����3'��dVP�3�*�o��fD�+Fdj��}���
���l xG�S��"`G���k̥5���_xL��P`z(44�QP��@U����z��R�7��g��S��XKxg���ڟ�pzF{�/Լ�J/ِ-��� �Phh���~*ڽ������F�o�SX!p:�/[>3���/�E��mGxE��S��y��,�Y2�B��ȫ����K6hL�;�Z,�ԃ�L�g.���W�gX��%ems�J�X��"���t��8����R�fT4��k�t�\̖��V�A�wU�a}C#�n�>x+V��dҊ!�(^c�ѥk%��%����vX�W3>U�Cf}����� �W�����2�D#������6{M�g�}�l��o���ٸ��ߤ�Wu�a��ϔ���O@y6'�@@�S��+�7w�;�����R�g�Z�������o0�s�;�j�Gz�x\{����Y��ޠ�/lIg�Exg2wv��ۦ<$��S�Nw��em��z}�YA��r�dz���T踏vq�im.(	�K�^�,�ˆu�R:��Jt�m�Õz��ލbs����x�y��m�"�L-���O�����b��c�Cy�~צ�AY5��=�ʩ�ܫ���Uo���s:���Pݭ��B�札�$z�����~�!��{�z^}��HA�2i b��8���Fܟ��X��P���د^�.�y۵�;����\L���#����}~�?;�C��w�ᘊ�\v?|�q4u��m����yV��C�H{:��w�0�������7��R�O�L<�S4���t�7^�f;���ٽx=�,_��W��Ra���C��1�=m��u��|x��g��׳��5،�U��� U�6��eP�i�z�%̵�}�K4arJ4�(�����S�+�]ޕsJ�ZNo�]ʃɢ�������/ut���5"Û!J�<�\�u������so'"Y��P�F.ڛJΜٔ��Б���֣�3+���L�e��:��L��?��~�3��&FS�1��hԳڊ���m�?t��$���I���� wJ�s�٧L{'��s1-�QPݛV,�`t�35ߥ��.kjۇ��&�k���P��϶�u����f#=�n[�$48�T/\@E[�����gf�B�U���x|�[i�����H�S��C����;2��`L��� �64�U2�\MEGA���D�ef�)Ey���c���ݑ�q�?M��*��w3�σ���}�%窐^����s�#F���%1�9'��%YW�/C��*|&f�K��ީ�С����2�ݟC�>�o��
��{[� oxWO���3og�7º6�誸]N|a<̏/UQ�T4=^��b�9T��ej�b��m�=ޅ�yc��߃ёC�b��?�V�񌭛�v���f6��BG��񽯧s�M	y�{�M���|g����3g�u�ޑ�6�cMm�̯pr�ͫ�u����v���䳪�c�5�����ϲg_*�{m�3��x�yaSr~ע�L,��(<J�k�,y^T���%(V�T�H!�V�$�Z�@|L�����WO�deVVm��d�YU��Z6&b������V�S����ټ{R��+n1-c�^�U�,��$�����7�5�7�bs;���p5�]�v�G�ݩ|�B���fOiE|i�+��u����v�_��ec�!x�G�����)Y�Jt�S�[�þ�{w���.����܉�~ʭ�1Y^��W2cq?p���όw����w�����K���ӜkZ�3Y�gd#w�<�3T�zs��߆B�Y�dh��~������}��]!;}���C|v���!��d!�[S<�ۙ����2��=7S�~*}�W���=G�B�ά�����y*&9�Bu���ǺV]1�:�g���X�����븞8�4����8�n�c������˜k�m�uv�����Y�k��_�t�b�X���k���:;9e��t�)�W�\w�=�!rb��!����<��鸃��O�^H�:�U2ص�MI�_�%f��t��X0��D��x{��Z��q^�B^~�3>��y6��ڡqz�?
�[%Q?S�u�Y���4^E���D�xn��J���^��=U���RۙQ��C�w�J���`N����;���"�����x�K�KEMƺ�R�|���z���/z�<�{L��'�`�����l<�
�#�ڼ{�w �HVqv?��b#���Z�c]���˴��T#o6��Mm����yW+�̬�}7�9D�P���ol-}K��ܫWf�q阯:hU��&��}�
()Qv�	�˼�fk'V�P���QF;j�3�b�����;$��8?�Ӈ$�d��Xj{ӊ�+���`�μ�'�oQ�k+p>��OP�u�*�qs���|m�H�.�;�c�\i�:}��0|�uמUϹ���7���,����^����Fm����Cy��Eo��'x�;�ˑ���*fm����y��T2;�3��7%{F������V=�!��\�9��K����R_^�;�X=��1�c��������l_�_Pϟ�'E��^ɏ=�VPѮj����
���q�v�w8�c$�ˎ�W�����:��^> �k����$G�#)Х���vE��O�]����>�>�ar�u.ʫO�ZY�T�{���o��O����/�!{ƨ�̅Y�
�e���.�;�6<�Y���!pG �4�$q�s4k��ʭ~��mK��L�~��/��O
��H��o٠ϣW�����!�#����!f�R|����3_E�!�ÅB3�
�|u__o�ѓލ>�kX�#��;9��44�{�ҳ�K����6%�8f{Ʈ�����٥�+�V������=�q�����1�lg��p���������*�<��-ԛ]<�;'���<_��4�e[�����2�,���Q���tl�yx�=^�;)��v!Ag(ަ�Vs+-m;u��sun[��˨Mt�'�t�y����7��q��Y��Y��3�Oy(�_wQ��G^ϛfՕ'��2ڦ�������Xu�`�w�9��8����@J܌Cؾ���#9��V��lzM{ٞ�=�� (7UU�q]�������D����TO���X�d9Z3>�o��1F��xdz�8=q��W�R���c"�k��K��݄M�.݄ �!�/?��+�u�9�׭p�'��>���6�����~��r��i^�دWL�F3~��1A������"���]z{���B�=�H,]���ԖD��=�@�o�~��}Ք�f|b<	�q�� !�������[�ۭъ�3ޚk��P�h�Y�.�*r�zo��~�L���ٓ�߽Y�I���T���y�ߏ	��N�Q_�3z���I�����͵���U�t��-�NG��0�z�tw��ǜ��+ӗ���ܗ����ѭ��Y��p��h�|�zU�x�ڔ�>��lz���T�t��J{�֮$���+�,��E�9i����
pe9=�zM`��S���Ng�ڞzA�5�����>�	�cdz;������ˮвkt�<Ynr�*�91�[�5������A~>	������vS�!���t ���@ɘ�J'kfu���Vp#�C��a]ty7��`I�.=�H��Q��Cي��$]�e���[�C/{o�B�{U����u�t�)�3.3�5-{�˓H��-,�{���lВ������|�o�;]t���2�����BٓI,��w��rW�3����x2����ŝ{��X>����W�Fc��G���>�OxT����R� C����%wmKv��o�S���ߣf}	q�1^C��0�y\y�_�g��l%�����ʷ2���%F����]!�����g��c��ϦE�>�/hŅ3W�H?e&������<�Ԑ/hxw�^���EQ�v3w�|���$��v�LϘѵ3ʽu84�s�5�	I�=6��������=���#}\U3ϴz��~��<��߬9���**��ڱ`/�X^k�K�K}QN�B��Q��M�)TVg��T�S����:�=��)�|5}QP�pmo��4{��&C;��;<�q�A*ke�=�l)U~Ֆ�,��L��́7/�T��hq��|.���6�1�j��޸����G����r��`�O�T�/;>�s5�Z��p��D��=t�)W�V��Z�QrU�i�m�?|���}���~�>J����k�V;�w3�7q홏�{��]��O�6z��T�� �u� ��ײ7�dÃ�WY�֒��Y�NИ�&Cr־����2��o8����� ���a�'eQ�79C�h)ǹǕ���r���$]:@glǯ��׌���ܗc��
���q+3-wi��@y�JW�r�m��V�U�[�F89���fG����C�/T{��N1�u�u�������b��������4�ߧ���9[7���*��Ο<�&,H���;�j�Z�Ɩz:}��x�l/\��e�����A��Mv�A�������9��������4�%�\ʿ:ҦN�>�	ϣ�M�c��ұ^;/2�vMn�,���q����Pޖ�s�^����k]����|Ds�_��[[��R��==��}�A��F'0cL�f`�qo�[�^Ύ�}c'��q팪�Q����2"���׏�lyS�}u�/{^zg/�[�
1�0{�|m�Ϻ_�ڙ�HS��w隈=��U'^�|m�b�Y�g�=oFG�^�H7푾X:���*�=�Wl���5�����X�\Z���߀T���ef>�����}����=-*������1~(�^�R��K�2��n����F��,� �����~%Ab-,;��{�L�7�{Ǧ��~e�}ފ\;"7�3���#���p��%��6[1v�F��W^�_�*a�*�O���;_�ݬ�J�yK��&ﷇ�A	5�c��93�UaB�t���E^���;y�g4��$��:���L�DE>՗���C�?Ʀ.\�g
�{���lG_��
WZrmd��V����q�����Y�[D�*���N^�v;�}��0� �����g-!�� ��mHy�o��T����g>�W��1"|�ǽ7��~�j��x�h�r����ɇGu�͓�]φ�~��k�W�z��B�x�̳�{�����&4��	6w+nO;�����P��V�nD��G7�0�����6=AmgyFd��{�<�W}��׆���@ `Ty4m���%��T��Ȅ)ΘLɍ�VI�"{�i�f�:0�O����$�|�+ճ�,��μёC�q��p����zz�뭑]ᶅ��Z�z�Ź�n2{�;�γA�~D<��W��ϲ˩�2�9�P��{�Z��zY�r�T���V�CdW�����$Y��y��T3�s=q�7&!{E��j���*۞�?c����z3G���?f��1��uvۙ��߀�?W0�B�d�g]M��쿾��΂fW��:�fx�UA�VWM���F�ݥ2�K��퀰1����]Rodµ���̎���}�Zi�'po��X;)��Zx}*��ʥ,��w�b����C�O!�y\��=�vlb����(��e�h�L�]V��5�&�d͍��ÛS�E���#��fs���E��;Y<��ǝ;�;�-��̓�<����R�����w����sO]�yՃ��Fi���6 91F�%²���e� A���.
�U1<�+`�ɪS�.u�ӄc��d����ӟ~Z�0��Y#�Eۙ�]���V�Vi6���K��)�]Ҷ�5P�,�z7֘��:����^#������lU '�*�s=u�x2|���.���g�=T/��&����#��;9��|;=�����*\��`f;!�; t�{����=�fԍ#���z��������U�hpߟ��#�ǯ�v��k��������Hz��,Nc��gTW���y�H��3�U§ ?Z����{p87���R�<w�?Q��!��j�d�~�������5_P�3�j�pU��^C3��r�o�ϒ1F+�g�-��h�a�������j���B��lM|�۾�9A��/l@[ᓿRѹS�ج0Վ���t/}Ε��\���U�e�U�^���� �hh��ۗ�"����gR�zsvh+׫�9��U)�d��S>��U���+����7՟G�tϏ�9"L?M9^��Q�|�<���:�;rJ�����g�ڡhZ=g揧��f�&!z�0a��ϖ�ϧ>&�ߜ�C6>��P���?~���p�Ec�������98P�	Y���5]�g-]�K�K_f�wX8D�X*r=��&��sy1��s�_u��%խ�'�����'§�W�`Ѵ~P��W-
���N)���-�Y'l�B��
J�Dz�iuN�Z[��6��p�w���*VSX�Γ���]V�nW,��lR��+h�qLv*�*|1���{�ѱY����g �;o�lp���_vNՖ��F�29�^�+t�����*y���ɏSX3AJ;�2J�t-�Z�����2��o��j�7!��Ɩ[b�/�b�Eu��-"D�C8M�E|Fv@���}s�+�!������8�:�1iP�Mj�܁����/',v�h�<Q��nr�����,��L�K�YM,�yX���q�-�֭��].�-��r����i�F�j[d�Etx�N���������v��Yv�sJ�^���L`��528!��W��,�1�7�E�n>��]�j�ޤ�E�Mc�j������p"�ڵ��i��i�|Ga��mnO�--��u�f�8��W�Ky�Eu-
Іwu��k>O{T�!��K-d��`����-��i��n�?�J�<g�i�E�V��z�j������3I����'R��Ai�۩��2��}�յ;[4_a�� �
R]n��l�[���B<Κ#��gn���NG��*��;7�s��omN���T�"|΂`�,ކ�;���*��$�&�&V�u��#��:�"���ܚ�/c4�*m��Χhw,���o��2�[Χ��"���A�xܖ~s4^��)~���J�gM5���-��ـ���N����r.c�;��Ϯ��̢�,t��S��k�BWeY��}�����<n�:&���oju����Nڌ}`�����A,��Pnժ�vX�k;*�4�f���NK�&�}��C�vX�;	*�&�uK�7v0�����w��â]���D^��d�q�՝ 2z�5ج�� ��.Ȟ,s-����'���k��,�H/�96^��[����.*
��gSS�<ul�L9˫\�#�+�*E|����u��Ɇ�\�+)��fn�+�t��ͬ�殀5R��+^��͆I3vIA��B٥Y���/�v�ou�f�3�%�����S2_u�P�z���u�,���n���]f�=�R�]D����:6l-p�i��:K�Va��>�5*�A������:�O��j�u������]��N��w9�He��Yf�ԛ��Lf����� �s��>뾼��Y��ʉسm��&U��8U�;�f�i���:�v�E��j�;Rf;V��cvh�F�YT��ĵ��ףb�`If�o��9݉V��e-���B�E��q}��&��R<��Z�Y s޽�}������u֣�.m7W{!5� �U�W:�f,d��x��ǁC�R�I*�ov`�>��s2[����HrH`u�M�D�%�Z6n:N������z��_jt��m��Ծ�������bb�DE����G5�mj�C1.8�dĵ��(�,���֢��Xhh��+(�j��\�U����ڣh��EUĆYqiecQ��JZLj�LLH8�ZcP)J���*E6Jъ���Z��"9�)��hcb8�ۍ������YP�j"ܮ�sU(�D[lm�%W.a�PT�U-�4�h�F6�@F*R�r���Mj�E�Ֆ�eS�*��L,��6���\qh��`�V)KE�l�*4jV�DQT����Ę�JcY�c#up\˙q��֝".��QXZX�*�Z��[�ben%����J�ܵF�,Dr�2�Z[Eq�̘d* �Ħ0�1�k*Y�U�´���C1*ZUZʫ�
d�(-��m�-(�"[EET��q1DP� |�?#��q��#Y��l���Rw������\ז� ܮݵ���Q�'�{#R�m�Lnׅ��fȏ���Mu-�������M�U�mK}��To��\p|Y���{��߽��c�1��{ۙ�Yg��h�7Y�����Z�Gm5J^���w�VK�5��t9�U�3��ǹ���FS��3��E�������vQ�=q���i�
X����.?�i��k�xeg���U��;�bc\�m�{��/$z!��AH߽�\%q�5�ad��1A��˷9��9߲�|)aQ��}X|u�5�e�zeg�,3����'���5}=�e�ގ��B0�HtPxUC�� ��bw�u��%���g�U�-vdW�:݈�~��G�ߐ��D�~��>�)�+���#S�>��M�{��^��}4k�W3~�nR�e�0�2��p��Fo�������?;(���.Y��M���m;�]։��������fۿH߲�������Y����������tm�����K��Dz�v�[V�ϤL�,uL�?_���t�2���}BR����>�r=��Po���<-�ú�����_1����Y���Xs��5�T2 ^K�=i[���.b����T�̾�7x�#�/#oS̫�5��1��:�� ���������L��E�U�f�>�{ ���O�&��̣�>��1�݇pm���%C����m�tc̾�Z�r
�쥬�O�Շ�Y7{p�ɮךlv�j�u8Bļ��R�6]Ee��ټ���L��gu��E/Ý�=����l��́o�FCCMEB��@@����*����]���\w��w�M9�����>�+>��-�Y��c=�m�����MUb7�#ѕ|g�M�9�����"��X�Hn��.�	�o�����xs��s�[3*��$Lﷱ_������yĳ/��h d��*x�m���w�/6�Xϡ��3p��x��w3�/ݴ��,�F����o���!�@_���{��+���9F3oe�ͿMhs��WS�&I�?8��T&��U]�����_��
��+�����9Y��~�z������9[��6k�k��+����/{2h���[٣�/&}�Ǒ�ϽX���޹�G�,͟{Mh���h44��<9~��=�����>�ۦ����ﻪg|c8�f�Y~�/�O�Q�}<|���:�^�27 �G������=��5q�y+���f�Q��1_~�����g�G>� ��\��_K�,=.s����!�u�`b��52�f�2�q���pz�X��Wp�2�}C�0��d�������?��;��4G���"}[u�~��g�§yۣP�'P�NV�qB1P�am��u���5��G2y*��dLǎ����bfU\�/L4�J�)��4(�W��}�����{�:�+��uST���'k�uܬ�Fyw�vХ�/t6�2�q.c���ܛ�7j0M	i�nueS�W)ʑ�Ng>��0���u�ߺ����Y��;����"��ݚcNG��}�^v�|�y�%q�!�4�϶�i�g�T�z.�z�-���O��
|B�3lW�����Ԯ���}��9��}�=����ǲV]1�)ظS<����@�B���kcٿ-[ÝG���y,�f;|T��yۙ�Ev��z�v���!��_L��彝~��w�xU��t�N��"s+H��$f���H\�~��?m�>���>,����p��d�O�av���dz^Wz"�g�(T��d(��
��/{��A��.�򮐌��fe��lUJa�4�N�K����n�P5J^�����_[�ѹ!�n��UOAo�q������[m�y�LQz�^F��܂���}�4�^
�������nx�zĲ���{~�ȉT�r�6�����i��NO��#��ו���k��0�������GP�b��F3N�9^���:��S=���=7��so��2+��^~�C�W�Y��;��1{f|��H��)�X��V�/D�_x<��B��zһ�ugT�+�\�I?u��$��V��e9��n��[YDA,ѣX��\ȼz�1�c̾OQ��?*Ww��9�PeLc�O��t���;�;&�`�ҖM5(,�iS���o(@p_Z.-)�D��c����]�P����w�Z��8�߳a��аz،�.���W��Y�s3P����Wu�C9x̣���Ь?��8o�H���>�~�(.�ҽ��]�;�W�=�T3�Xh��Q���f�n3�1���2!x���g��x[5~�v����:�����r����8���s��0�ey:���3~��^�{+]5��t_zw�)�cЭc�9�Z��
�V{������X�Y��Q���;���pg9�¹��.�xյ�'�U�]��G�_��#t{�\k����80��Y#��͎�r��_�;��G�{WHpF+�S���wռL��B�1��=������ϟ���v*���{��v�w#|��Ƿy��]���Y$<�p���L?K�!�u{�g}���_��;%K��1�K���~����_��zj��C�3Z*6}��`L=ϟ\<��1�lg��K�g'����n��ʪ+]�][�w%�w��z"D���:�
�ڐc��h{��9��F,?ZA?PC��|N�{��s+v�{������Ǖ۰�D�}F*�UT�@�V�ȍV�3��Ww���&L�5ݳx*�=�.��`̹/F�JzN*�#�mE��t��(i�ؓ*���C�p���6�Lll���5�etR��Ѹ��w�1�;�EVd�n��U���1�"�~�4�N��81�__�A��{�ZΫ��
��;s�ԇ`�:���q�7-I=�z�Ն��C���~��=�i����n�>���QP�pm_[���χ�hڼp�:r��{�{<4��d������}]~�>��z�+ճ+�&5����n��v�h��<=ҹ����]�s�=��s���2L'�>��A����	��� p̏o��%�۬>�W���a��}�<q_P�z=}OI��O�=���>��w>�*�bt��#n�����ux�>[{>;�U��"��n�x�m�����*����7���Ȏ��Z^SY~��ݙ�l������/|�]`>t�T�h1[Np��]���~���U��n��ǳ�X���'�{�+�Wo�[^lh��ﷺ�KzkA�<h5�S�����*�#�W���S��
�)��v���ݮ\.|fws��ｷ�t��z����5������h:��?r��Z�Y�z��S��������^s��=k��#�;\fy���o�	/�� ��N�����Dr����"��Z[+?��4	��5�<��b�A��F�NUoz�/M�y�l�܈���d{�~C�����jru�E�]ʹ�Y�(4B�A+��y�&a�b=]�0���j��Go_I/��8z����WR ���*ˡ��U�;���{�f��X�y����n�.tĒ���PXoS�wf۾�^���5#M������h�%�siWnӭ�T9I�6��7Ȅ}/%��ˬ�r�dͣw[��}�73�UBnuע�:f��f�L3��a�d6|�/���
<����M��W{޽5��l_�������_�2�ٞtbÙ����=�4�~Whz�IFǪ��95ꭓ���U,!���W��� -�a䉖����sa�@�>c_P�s�K�/�(���O��������Q�6<'x�=��'i�����5�F�ex"3#`f9EL>}�o�\o���_�̹�^�AN|������L�9��<�FKC{ꊅ��=@���dz�OaW4�P���{kF�����}��Hzr���w�-�~�ɕ��0&���#�/2<b�N���#��EOV����S9����[�����\=	�kg����;��`w�2�|�j�S��9��Uu�/τ��S ��
3��bQ�m�G�ĭ��;����h�����U	Ǫ{:;w��9������m��X���4�f�Kﲷ¯i�/�����&M��58r����Kz.N9�PU�;��Ǳ����0�*cOշ��~ͽ�`Ь�.�>j���|wD�h�>�u���27�e�g��6���g��m�E{5��'�L��k#\×[`�cx�S:�˕�#n�7ljcJo�t(꣩a��/B�:��<u�S�^�튎����ll�}ş�8�0!;ig)�Ԍ�3S>ƾ��)o���9�$W�3J���}���V��g�޹b��fl����;�]��hhچg6O�mi��$��^q�c��O���1��w�8���e�����@dy�O,*nLk�{%d��F�|9
���bk�v�MȤ���I��i�q�����5��u�~��}��=��ù;R�����g�w�s7n3��ma��}�<4�)��bx��cv�F#�0k�1����3��S�]��u
�<�ue-����%^+�Cc�ֳӑ�n�Y�4�9R8�ۙ=뇹T�z_]?�U��.D�]z�7>����I���U�}���KH�6�i�����S�Ϯ�z��R�'�0Q��uY2�^�������H�'z��}�^�a��^@V�.)ظS<��B�����pa&�k�ң��qp\縉O=}7+�V��Ѿ����dzr�Q�-ѨP�.Ѭb��=����]�p�� !���bU�x�3�O���
Cy�3�p|Q��G��:N+7ys��α���[꩟x\W7��D ���W���6b�{��ϣ՗��yd����?�/e�#O/�l��9��kaO���*l�Y݇�(,�qh6Z�x+���Y��[����I�-�}��d֫U"Q�/nt���e�
�pt/����i�%[�g�n<`�\I�0A&P6���"�k��;/gLUn;/���l�F��U~S2|�����ҡ�^���T>�*�պ��3*��Ʒ�0�*����,�`�I�̖�<��Ѐ:.��ʦUǽ�p]x�hi�nx���.�-7�|;֒�z���n����؟v�v����~�Pa���VE:��lqu���C�Q�h�^�~�H���L�2*|Otߗ��P���Ԋ=j}m١�<���:��Q�Y�-X�5���,��������fW�=z�/Fm��t�;nfv>>�:�}Aw�g���f�{d�w��$�~�9��4s=~;�Xƚێ�c\<ڬ�Wm[���Zπ����������:<H��=��P�Wg�|�od�졣MR�`hrMe��ֈ�s9��ק�ڼ|�{���1��9y��K3߬�WzG�0��fe\_o��������έ<>��~U)g��"z�\�=���M;��t�����o�j�{^G�m��	�Y#���|k���k�𓌌��SW���\9>��ۺ�^�����C'�T�m�z=�����Q�T���
��y��sp.,
:ck���0{��b��W^���R�P}>e��6��]��y�:b �=�]�m��)�\��j�����^��jS"dB��{W��H%1��>�n���R��<�k��̧���\4��(Ě�퐶��[�\�2K���������s�K� ~ݯ/Vm�?���~���E.�~�?R�.HX�g�6X~��"��]����{]3�%���;'�օ��������=�=�z�������^��r>o��]�Ni���WXC�$O�\�-ѿU��nԃ�����LĮ4�O�!��B�ƻ��7ޝ��<���/O�π��L���.�*�n :������!>u�jww���YY{j����r�𣏕Lgު��z��?g���yv� 2�C�EB�V'-�xl�$g��s}�����ǥ*[w̐}ºt�~�Kڥ~�1�v�T<2ew������ �A���u�Z����k�v�H�w���Cyj��T�v}�ΘN�%?Y��S��VDS�������7���Ԏz���4f�Xc�xW�����F��RR��L{G�������ߤ��&��:��0&}9���(�r�<|'���}�4<0�t��F[7n�6�å��t��l���y�������zVV���}�>�C��	��5Dls���+@���ެ�FT���&z�WԜ;���(���Ӻ���;������o۫��N��Ȩ��1ϱ�h�&U���ɴ���`1�a�W�V�~��^T!�
������O��5ٝ�J5�ŀ7�+��!םZ�Nΰf,�o �RX۷J�b�I}ZY�� {z��C��F����}s��:◕��<h/)c�m��Uk�xY��Iׇ�ݕ��gN���%�8��������o<:G�M��ͭ��r
�a�/�~���L�EU�0cdl_�����<2}�^�5��y��ο�_��k�p�.�x�z�����z�ɤ�E.�!��}/Ee�w���b�n����3�z��@�V]�7�+/v����S�����<~W�N��o�D���}pzz��C�~��k�qA�Tb�=3__x�1��-w�C�#Ȏ�h��6���1.�z��<U��;�~2�j���5Lo���+�=�1a�����	��k��o�#��M���T�wrD��Ϛ^�.�	����]2ϧ v�!�2ؿ�T�#�sp4>c-SS(;��ի3��{e�	�|��M��[�*���������\`Aw,A�q��)�CUB�]��������z��ޯK��TъL�;���ǫ>ڬ�^��;�n�,��\}�jږ�����@.!Z*�mhȀ��ÿ���NE:��jG7{3�<&*}��A	'��$I?ā$I?�	 BI`IO؄�!$�`IO�H�~�$�	'��  �!'��$I?�	 BI���$��$I,	 BI܁$I?H@����$I?H@����$I?h@���!$I<!$I?��
�2��lN����������>��������    �    �P�  v�E*�B��%%D�*���Rm��PUJ��%)"�R�$R��P(7w!A����*��U	5A�ԕ
��D6� �J�X�R�,���*�p ꁑ�Ī���{���� 8;�%D�QQT�Iv�J(�8u.̨�(��DGZ%�ȉ�`M
9�TJ���Sl H���l��uf %��.�0�)P���PY���(�tv�����j������Ί� X ��h�H��M4UH)(�([
 p�)T��AT$�Q)lʡITM�E��r �f�%t�*@
J��m�
p .�u�D P4 �ёl R�/� � P ���T�I  @    �x`�)*��� �#&�i��2A2$�4�45OB=F����jg����JU     �4SEOԛ��S�OH��@ ��@ ��!)R0F� ��`�4�sÅ�S��
뎭ָк��	!C�2� D�?�Q����y�*
XЊ��VWo��ş��z?�����$`�A!P4��B���Al��FE/Q3��ϕu�{�3��==��-��
j�x�V�5��S>����E��4Ѓ����~��L������O��5� ��n�ÎN=Ƀ�>=�|�I]q²��f7q��"2�/E��ݏ��fa璍�����c;�z�
��F�}wy��x���i����jr��wM�
�F�掐�ͧ9vK�'���Z����`�8z-���3y�"��AA�[,d�dK�L�:�=6�Ѭ��$��;���H�Aݔu�;���l(b9�Eㄫv\��x��놜���/f� ��"P�Q�z�A��!�N���:P���y�BW��L|�y���z�z�Q�Wq�w�*���|\���:�^=�ܷ.S�;?l+P���
`M]�Lv�07p���vܼ
lA@{ۛ˖؟vˀٯ�,�ܟs`#�1��ӯ[/��_lU䝊���ԜŬ@h׭LgA�oK��D	�,_��
�<���㷻.߈���8Q�H�@ΰ<��۔5����⫷�)�������p���M9�xP���J��Gtb.�Csds����-�7 9Ԝ�g�i`���~ub=���j��*n��[�vK�h"ossy�H�g�f[y���F����j���H��b��#�}�<�사��45�W�dV-�t�k��cP�g%w\��\*Ӂ-tt1��8C�\L�Q�F������Wsw&��2�2mJ��æ7ہ	�.�0�l�tӯI�D؇T:����,�#��N�艢Ӆ����B'S�����=Ɍ������6�輓�JFq�,�Nt�of�`e�%�!Ьߞ���T\�m4p�N�滄ZZY�@�jR�/jܡhN���{������h,����r�
d�/��� l�,k2�&�Y����u���� =�pp!s߸�towќ�1*�ݯ����XV	u���o��X�i�B�l�&t5��Op<��
G���-�����0�`�gM/�:�ܹ9�~��ȓ�^�ݻ�v�V�$�K�SI�(���fU���9sFՇ�<SV��y��	���N:�] ��U
&���!����郣<�LZ�2��V�=�^�`�w �]��֙ӌ���Rɢ:�0��ؗ�w�Z��:gA���:�}w�$��r�r��C��
�@7�}�{�@_^�h\�q�V�Ƀ�5E��7s��݃xh7x�ã!��PQN�x�����繶�'e�9���/��4ږ���a1�
�wbF�}m�c��GV-/����n��&��/�:.�5;���3�4�=���Y���.��{��5��S�.dk�a`����^nw,Ե��q΄jܤs���e[&�ڗ#�0==�uQ�ۅ%�Ҥ�7W0�k���L
�l�N�Z�0���N���vt�X�u��s�p:K�M79[+TG�,d���7t�ͭ=�}��\�ׇ�тLZ8t����3q� %4��&���PK-�d�B)���Z�/�Z4�釓Ox��E��ǁ��H��q7�> v�}Fn�93\�f�1�)so�Z������<:�w|�Nك$����ɞ�xX�tJ����Y���7�&.�\�uF�#�_Z���Ֆ���n(�gh�=���s@�^v6�{��=�g!t�[��S-� �+p[������u����\޴�	�M ���x�M�'7w�M�T�>e�^l�ۈ�s���N|� �f�}�;��9��9��B@sp\"�����}�����l)�8Ah�m��A|�$pm��y˳V����R@�F4��.٣��oa�4��]Pt
pQ����zf����[�cc� 6F�>��X�̷�M#rk!N��/8�7�hg�٨v���.�����YJw$�õ�i�.u�
ᏦN��ޘz�s�@ ���,&H�q�g\���yDeGQ��>`Z�8]kun�h솎cQ�Z�s��v��i�x
`ԧ׃��kv����	����:���0�����'09�ݨ�H�i­ia/�����:;n9���Kz�Ў���tt�	��K�.�c%�(�~w��:����voj�������&�V�UN�6˳6a���Z�ϸ׼��%d�{n�WU��rO�����������Wxa�;�g���++�x`�;�z_a�B'�U�,��ӻ؋�RG���vP��4�lwg2P�����ak���ڥ6�4�.���G<t1󙹝CY����ʪIƭoN����S����c}F��&SI�{.�&@��X+*�v�D���ؘ@���٧�V(	6�ژ*W*���1����]���UYnv����9�x�lh걹�U�jɤ��|�ۋK���+� n��c7R�4>9�b0��eN���n��ʦv�5�k4<7u�09�3o8�ǔq&���Ь�e߻���	�-����{�wϪƭFH0��5�$z��ˬ�¶��W��Q�W�crJm�I(�%m�)��$���m�X��b��Q�J6ےSm�IGI(�nIM��%$�m�%6ۤ�t�����n�Q�J6ےSm�IGI(�nIM��*�ֱtnKSt��o���_=&蠫��򖁒{��]�tu�9��sw,g�����G����:2�b�+*6fq�C� �yj{�!�J0_zޘ�P�H����V���K��Tk�H�`���>+�%G�� w��X��g� !�'���5�7�e��hȆl;�q�9hͥ@�붆f@uN#�w���#�: t�ܠݫp�ڗ_J�n��<X��w���=;������|��F���:�1]���x�h�r���׫:�����s��E��Fl�y�� �{gc�қ��=O<�M�=JC��!�R|�@�������(X�i�9f�r��9v�۾h��T�^mu���s��A�gg������MuY�Pf�g,"�ж>�5ey�y�sh0�x�i��;q���1/\[��a��f���eނ��<���>����Xyb����4w����}��wKE��T���P.�wڤ��ǑgF��l���q^G�R��-=3O��W����q+n�ޛp�MO���9��y�y��X>���7+RG�b�}�0�퍞_�������u~�{!��xk8q��H�Gk����sK'qW0�y��d{rk��޾��v���ȼ��\w}݋�jh�L�n��f���>\ߜ晋���
y\�Ö0�X(��k��P���ct\��yE��غ`�������<\�)�X��cQ��w�
�Ԏ�G
�)�_d�v�#[ҧ]6��� D>/x���
4�V4���������W���W���b��~�9]$"���ʂ�[�1��G���nI7�ب�.İ173oh0!Mr�G�R�D�f�P�I(@%jw&�^L�K�k�n�}�A��87b�y�_��;�s���^CI %hbe�֚7`]�֮vH 8$���7rbxtxx����3�e��"���~Ƽ<ʪ��KYn�X��|%����v����`�r�XҲ֪2=�h<!ض��&��7��
�%�݅���φ	L�8
��&��+�OZ��ض�|�b�.�g"����B�GTG��xF@|̋o���gL]��>I����'8�&NXF��t:=�v&|wlH����3v%�N�1�'��wG�*{^mh��:�JT�2[�ؑ��\#����R���zK�����َ�2��i������H�7�	]�ǡ�%�ƵƩC�<Nz�>#��~�n����ᣁX�b�@��>���3��0wo�"\2�y�.Q�K�/����1��#��$�)�w��~�A�\���3I0G�Z+�"��'Ms�{��z��2��=\��n����)z�i�O>^f,�,Pe�� �@��Ab�d6�� �`'E4�\)bG9N����"Ϋ��)7�߮U�z�g��y���z����%Ԏ��5O���wj�9s�ҁG�QO	�I�	N��M��/�%���_l�nQ了�v�r�e>�'�3�!��,'x�s٫�����6r̡�m���+��2D��nZ���N�gK0�-��T��y��n��N���fru#�T���е�8d�L�[��wFu���x2!�Wn�4��g�]��K��]�)ɇ�9�D��>��NY�e�7u.���$�Ɗ������'��Ф�g� �)�%���T�B�=�$m�SE�iv- f��ā������tX��\7X(�Ner��a��hyA�Y�_a�$!�1����D�N���B�3j�4�RN��tL��G�W]AJ�X�R��j�[��� ��i+��ˈ�-\�=ˮn��L.�~a�K�r��o@�9��	�T��|�4ھ��;-j��Z9@]��K̤�=ļ6�����Ä����f˼6c�.W���x�s�L���x|�qOzO�՝��+/`�u�H��>y��bs?��NX:�(�l�o�����z(����)���2���i��a��^�_�A��R��\h�{Kq�}mԹ��t_uҾ��g����]��Q�3�d�`5�SYƭ�}��$x��`��q��<^@a�tw���l�`)�tGe+���(	L�"&��b�����/g�������/s{9t���U��Cɨ���V��.�\<uc�o��_j*�V�����n�Q��kɛ�cn�%2�Ws�2[S\Ǧ�p��C��H�qs4A˾q
}��٥M=s��V\{7.��Y�}!�כi���F�Vj���2G��\���-�uz�Ϋ���}�ﳩ�t�g
9/N��U�`�kwLM�3l�S��Qb`�o raTA��ky^������j�]THـK��b�M��xwyTv�Uكܐ�#��M���T�1�*6�۶&S�V���_Z���Zִq�_����w������Rr�����vά������� ����Ӯ��U�,OUKx�=��Z�9�6��˾�����>� �n[�:�_�"��I�r�)���v��/q�F�!��$<ː���Ep@P�� �}�w�҅���#�5�.����B���c��мh��ٱ#;y\�V�<�z����$(ƴ�9�����!�l���moq���8o��rn��5��3=��Fo�<�R��O��9Y��]���)�u<:Y��8��7UD���x��7��v���X�_�J$}Պx��+��^���?[�)�~0���{.%�ϳ�Ph���̋VN��o�%H��PGk�~?���]oW'�c����D�i2�unNt9���m*f�K���	�������;h��`F̡zӋ�qof#�:��I�s̨��&p�XK:�x]�l�箖��o���G�W��_,��&m�ߧvo#z0��d��5x��aE�"޳�M�����0��'�4.=�|F�7}���C�Ȳ�[0�۵,֞�:�w�VK�r��V�+Ӕ�Q�nʙ�6����|ϒ\�^�N�w\=���\;��*'��d۞�z�,q>�^�A�<$�/CQ�8���+��wx�������5f��܈�l����	Ѵޗ��ޗ7:U��%,�@�a�k6U���q��B�I̪g9�7���	6�.2tnί�5s�`=�n�W�i���ք�g�C}Ӂ�Tiz����M̗��o�L7r��/�U1*]�^!�&t��f�쐕P�����zg���rY�杨��g�f��{�ͷs�}:4��x�����oj^%�.��k(�����kZ�o�<��޳l�g� u�OY�V�ӵZ�Q��unt����r�}t�]�fk��j^S��9յ>C���7�(�c��>��/WS<'��C�/f�Ҿ#��_L����lW��l�1x�vr+��6xKH��SK5��h���$��l�y���+Xڃ���۹�ү��W(���R���x����֎u������۫\�j/H=�w�� <��SRӛ���w��I
s��=���=�PA��CZ���߬�A�Z��ί{�nx�q�����ᜇm}��;b�����xw�&��a�i�q׳!�-�VƊ�`��	�s҉�H��
,|�2el��̛��͹�1��p�Ȟz�ȱ�Nf]%{��b>�{�w-ͮ��Z��|F�0�B�ՉLY��W�wպ���oN�D�v9s�%􍁷�������vq���;�b�3N�s�d�lWg 3+�9���s���W���`� �t��KJ��$�^{�v�`L�Ζ^�����С��ڮ�}�ޠ���� ��A[�yS"�����^y�v��n=[�����f���ڭXx
k�e��u���8S�Z��Y�)W�zGn9�ȴ��ʗu`���M�����g�yf��yC�uρ}WZހ�^7���Z�BQ�x�XE豈7ޛ���Oh��i{�:�#��%W����h@=ϙDd��Q����7��69{��=�rZ�}��7}�-��]S�Q�Q����B���l�с泱#�ћ	�9Ъ��Ų�����q���U��)�榫p:���h�+۹	����^�á����5^R�ԁ�A�`➭�K\�\��d�;,�d
y�z���.�e��W)XPe��k����y��#&us�O8�v��>�=8x�)_-�M��٩ʀ���|���.Lq�t�5�>��qEzW�jܿjO'�=İ�L��^Ec@���<��%��|s"��}x��x�nh�{n��K��b�_�&{�3�;E8�����ɀ�����s}I���6�8����Ǘ�l�9�h$nMc��p�%l oB@�f�5Jܷ�t�<꾱hh�oGB�l�G:�ܫmr�s���a�r>�1Go���N�`N�kz�Kѯe�CG]��W����Z�G�kA�E��ui��7� �w}2�"Z�B����S�WX��+;��.�Y�ފ�tl�O���\|� G{tp1�B�� Ô��V#Lo­�.v��N*ڷ�&�E>�K+a�u`������<�Θ��6yQ-R�� C��7��Nck����2����Z��t�����1ha_�M�MJ��w��]|��4�\�|w@�lx�Y,��Y��S��kr��{N{ފM�%(-ױ���1毬��!�����w�C�B�Ln>/����o����&*�s	o����r���xB����]��j��[�)}��Զ1�v�wy�žػu h�-U��b� �s+��������@�dSh��팉]v�n���i����b��I��4�����V�t�`o�M��L�o}�6p֯��.:о�ه���|$��%�W���/'���H��/5��;��{B�d�x����㈞J�zO�K��#�")��)8��t�=S菠|;�y�_��IZĕ��]:"`%R+�9J%Y�w���X��e��@[��.���5?��]cs�<z`z�����I:}��.-F����Q��N���ܧtlq}�]��Sǔ,Ð�˥�ٳv�;9���=��lLC��Ժuuܾ؆���ۥf�e�9cfi��T PmtZ�Y��E�ߦh���(�<��}�ɂ]u%�}L�[y�8�hئ����N�Ku2�Y��L����6�sc�j�q;LGk2�s�r�K���c��8�ip��:@��Ӗ#Ț�YpIq���s��뿀��Aʝ#�3b����"��2��ҩ�L)".���!˥)�E"�wr����L��$2��6@2eM���X�>KX+�f6�dH�y1(���
��0q�1r�N4�*j(��G|�4LJv�c�Ws)�:�R�j\P�6��榛�}<�BǤ)KM1�0\�W�̊D6�ir	�c��	˛��b���IJ�79i����2�`��  DE�NF�E_�q���������<����|���\L��Y+�Q�q+��T��l���2U�v��-��ך3^,H�8p����~1����\WJŌ9S3�a!��ܽ�	-3L�A,�f�Ю�qQ8(�	�xүzb�=��	��[��:/hߏKe��x=	+s|[�m���o�?&Cy1����ٟ�	���c{��ɩB���MC?d�^.�&��!P�w��������),�L��\mn��/%&�^�k
Y����V�{�5%����5�\pnU�����S5��l��g�FY|w���c�f�m��Ho��B�fB�)��Z;T��W��n��t/��E^�[>W�[#Ņ������2i�~�IO%��,K��#��z�y2��v�)�w�s�2�Ue�nݹ�@���\��dN�m�b�xE� ���q.�����e@�\����+��%����.���W3f��{Ye-�����H�0f8���R�򋷂��tz��Ƽ�&J��<��d�禂$�W>N^����N�+�|����ߋ+�g��r�;[�k��A�����p�u�z�(���N��"V:x45SX�@�W)�Cm�ˊlzr9�{���g��'|��Щ�1�p�O�=a͑0��9���ޱ��J���u�wm��S|��[V��-
F���ަb�<��h��_��b�i��Y��9�*����9I��ڏ�G���v���9s
��v��22�BR7�6b�p�$�5�uF�F1b���s�'
�
��')p�-�]����(w�>
��b���	�?7�N芶���˹rГ�Gi4�\}"�_qDl�.na����l��j֌���5���J��������{l�^�6/ݚ+���&Ej�b�X}�QVS��ӥ7j����0��+�����53�uL;\�"��2�Ą�e�Әe�W��W�(���s�5
W������j*�f�e*�L�hB���28�j	K�z��1�W@����o\�Ԍ����or�ݫ�sO�Z�8([�Z��[�RÆ�L��G�ۈ�W�';�Ħ���T�k�谾��rv���M�t��ݚ�^��[��F�{O9k&�zMnt*yQ� Ԇq��31q���l�`��S���Ƈz�A5Ә�"w���˞�[�-]�<0��L��.���,V7I�G�3������96n��L��3�w�m��<���N�_M̔�t�k�6�2�����yS����
5.aT6g;�R��!�(��=��xy�W�yz1O�"^Ȅ������4����U�oʅ�p_�S308��OFkV|�R�wf͜��.�M'Y�\^�΂F�*N,�����&ߛ(��ɇ���h��a�~�2d��^�b4��]�D���0�����\e� w)�{Ya������vƱIn7U�꩚����z��C�<B�8�A�"�̣`F�m��i�=EP�3����z����o�5�O�/>W+fS�E	�j�}��ĺ���C������+��g�(�@ޟ��h���^�Sr�b>��n��h:���X��G=�y��|�]��]e��wE*��	g>=X�T��1��b'n�'j#
��n���|]J�vy�����ѭۨ�E�Y�M3��o)QԶ�%��\����-H���$,~&�l��u����@݁'��)V������̭ŕ�13���=��~�J�:k���{	h3إ���7��ٻ3R��f8�����X^|�3k|��+� ��!ѤZ�y��N�V�24�H�5�"U�0�c2��eK=��^o�r#*4Y`7�w�GX�����NJt��2�G!
4vKY��>�t�%�$y#k���?Vu=K0��ko	��k���]rG���n�FN�U/���.�����R��u���%O���؉�%@�6$���*tb��y���<iW��4�j�����6UROj�'㗏�[�k�fN~^N!�ϰ�x����SI��7 Ъ�:��P��]9�[8]�;�[p����}
�6�����5Tb�;��Ct}*)����!�޾Xv���A�ʏ&�e�9�L�jV�sy-ƒcHdu.� �(��
ΐ��x�]O�cC)���	#7�8s;e��q��땹4v��ˌ���J੭�aWP��tc=�x:�l&6'.*A^�٘�>v�%��kA��mgr_KU�l����a���'�xg��sE�c���[��oe~Ņ>s�|~��w��ۥ��y����a�vF�j�v�ԥVߨQ�6�� b�u�U���GW���Vx%�%�*���U�qF�A�W^H	A�1��� &�ǈ����L��7$#wF���6�׶-5|�=�Ԗ�c���ĥR�:�J��&����iƜX�����@6��� �*�dӕS�ͪn��md���U���)�GDmsu����ɊHY��"�I�y�Av���j��
�K��vk�>�P���e�m [.�3n�n��ۢ��%�l��ܪӮe�w^����{g�Kk�A�r���c)r@'L�{2	j��%>���nrU"��4L�4���b�B�.52��L)æ��$᠖���-���4��Z�Ց��&$Eeʹr�.Z.��H@! 	jf�nE㐁X��#T�HU*V���!��h�\���B�P�M&K��Mߥz��,��%�f\�)Q=֪ɥHU����57��ý�!�h��M'1^�oQ�q����L�3��_��y�Y��̏�D��o���s���Q����.�~�@vO~��OU�Ǹ�P��1����k�7�����>���>q���k0��������ۢ���1>�u�i��ƛ׶=������k)^�X�%v�o���-�i���킘����'ަ6~HJ�覵n�?}�.���I��^Ĝ��i� "�g��}ϗRn��0<�B�5�8��0y��a��D�{�T}�~o]]ۇ���E�ߩy�Ѵ�*E�D���6���~�,�ʬ����~�w�������ƴ'�E����<g�W~g���������Ů��
����?�!'�_}�0֊�F�ۻ��O��V�H���ɸ}�2��DE���4k�J��s-
�w΅i��]���*��K#J�5���c� uEY��3��9�3�qbnǆ�Hj�"g��@$��9����B7Rg�ڸ��*l��0e��T��:�׉����r��5�,�0��uD����A�Rv�B
nT�����B��2��=�s��I�u[��o�s�k(q���F��62�{,R�G6�{L�W��j�$���^�ak�3����[� �4Wu������pP���]���d��6*t��� ^pɜbM�roD4؊\N��JD?}J��y��u��{Yy�r.>a�l�(U�'%��	�+(����	����o3ᴂ���9��ǭ�,�H�R�|L�M�ë�g�|-�j��5�sF�A�~�{�լW�W_��!1BXB��B�!*!�9�X�b���	���W�ZG��P�P��4��$5�CP�9�n.�nԃ����(�������\hR���V�*	�T	�f:��(j7�n,�c� �[Qj
B�Z�/�Q�V�C=R`f ^�/'Yp�*n&�ȧN�p�BZB�e���Us9�[o>޶�fufGr����+��`9�-Nz0�fu��y�9�lK9�-nv�I��`8���瞯;DN"�W�/�J���=D35 $��I��1Y�m��/Q� �E/-T�\���\@z�j#h��3�3�=gB��x!�h�D��( �B(K�����X(��Q�$��̪�����1-qSSqj+��1� �*f��Ÿ��㬛T��z�"�����&�l��P��*q11o�� ��~m�9Q�CqR=n�8��#�F�ҥ[6b�-F
�y��^y�i��縵o�D�
^/9�N`n(\�����V�Q
c�!p�Es�]o��oE���A�CNb�� �Y9����udSpL�s���:�&`�&�e�b���(n`���)��D#Z�!%-�Bo����U���1(_AK��	�'4��6��]@�T����h��P�\h�������,w]_���}(����s�Ǳ>Y�.��`�kZ���w�s��p����*k��8����@�@1��]�JbjՁ:��Ak�KAb��j9ެ!���P�D��"3�y�ε�� h�� �q@��4���P���!�������Ơ&4X��5+�b'S��ju��Iq�N��)@�������CQ/ o1D� ���	x6wH�!����f*Mg�߮u�È!�T�S�����J��#�%ANb��؋P��1��u�u�"f�8����S����"�Ix�����
��}ϼ��n���$B��w�D��PC��(q@Uy������J(K�"�v����P�gy��)�$���NalҥuA��o���P�S<�:�=q�3�(H����
s�mP� �!�	�qqC���4�q�3�۞3¥�5�B�4@"��ALa����/n��0S��;���y�WI �Gvd%c�ݺ�-�%��n�2�Bj�BFl����2_�ʖ�	"�VĬ�rt�A{І�fj���q;@������ ��3/�v��``�T�a�(�	i��L�~�vO���2z^������-
�

�v�~;�8��퓔k½��v%�\IAO,�V�8<�p�$M�+b�nI��V�\ⳮR睻��{6v�:ڹ����V��c���G{P����:���]��pq��[��x�~��[��P�y�Zi�}��Io�RYxg+Ii�g*�� �I�������1�DE�j����c>�����D�����.���+�r��\g���W
V�f�5�@|ʳh���ݛۓW�9F`Ѱ����Myŗ�䷔��[#V;��J��+����;\g��W�,��e��q�z3ٓ�\�Ǵ�>�T&
n��L�)�얱��Ț�çZLm���Y}��)�|w�Ѳ�1�nv���SQo�ks�산�����������k7���
���J"�v� ���_��q����6пGJԬW�<���T�{&���N^Q{�:�;�u� �Z=��J]��[򸪾[��Â�*�6O�s��ڹ��̬\R���ߙNc��c�l�����54U�^TdR}Ƕ2��J�L��@���ao
�9LӜ�Y�%�M�΃�����y1?;;Ԕ]��P�ґW�;��y˻���Dt�"=3���	 ) ,�� H! Ȓ�$ !"A�UU��?��υ�fo���C���-'6�ٸ��I?��xͯ��V�� �w%߿3�ȏ�D�n5�t�2`(}����v��{f�������S�]Q�Ot>�&���F�^\s�9�~'����gd�"8��)�Ǚ[&a]L���x�����s?��ԯ�t}��kÖo�fv֐�i�6��͵1�d�)>̴� ���B�P7V�Ro[��ݎ��6�Ea��(%o"��)ګ��ݪ��(:oS����6N/շ�v;��=R��gF���<�ͬ�.���L:�m�)i/���{'��9���avJ�^x�dz\=��]̾�Va���������f��eE���h��1���Ӻ�=��a�i�ՙ�T����H�g��E�?<�D=4/C����55�|�`���ͨ iv��'��p5
�A��u�Hʠ���˓"���M���w0\D�f�劧$�q�a&)��܌lcU��[cp�T�>��!���4�}Z4�V�5]Q�[g�F�2�� �S�6�t<Ь�u����f�WXa��f�!�L͎زLnuc�Qj�^�Q9���+Z[�N��.����yr���5E��ِiŏV�Y�D5�ژ���f�v��6(�MX��h�~�i�щM �(�Mb�\�S��-z+��UGvZ��n��K��_~Ҙ�B@��}R��T�υ" ����=�0�k��p" Dd��H�!���Cm""m1@���s���B�@�1�"ؚV�� �"'Q1D:M[Cb���I&F" D�H&ҩ�N@��]nҔ�LhkV�cLbVH�04�A ����vЁ1�%O����Lg`ꖍ�����0Ҍ+]�Z�ɝ(�fb�D�	�֚V8�4�K8B5Ӽ��q���-o5(J��#9�\�	W|�bܧA�)M�Z�_��DG�,Xs����Y���� ��&�������O�ѵ�9��3��J�j���u�o��7h�&��P��y;�+�[�U�X��)ɉ[�in�5�kK��h�0�N�Ev=�s�;a�˨ޭ���U:�;(�xO��78���c���9�NQ�:n�S�Yqm3�@I��q��K�7�'-^f���*07y7&�_F���0��Y�83�$��ʚ1�%��"=�	6�ج?"�4ě Lw-����l�Ыk�~���sy�!�N.�����X�a�V��ݦ��!�E&���o�N��zO�˱|�����,Ox�WS>�E����}�]�LQ��>x�xZ1zT\4i��{#B-֝� �]t>�T#f�N�ձ���t���B;�5�w�:�5g+k���{f��ŰK�u���q���x�(1������bÌ������X.b�缶�w8em����<����n�zF�\�*d��н��Ũ���E��H��������l�a�`�ˀ�v>-�>��`2,���y�]�C��y+η=$�]�m��?L���IA��P���
.�S:����^g0�8H4�[��Fk�Q�P�wR��Ҭt�' ��T�w�Hrwf#"�؅9��Dz=��ҫ=�_-���ʗ��M�Bs��cMp3��@�I�.NE^�:���M0�j�!\=�u�z���nl*A/���: q��Ó�sd�38/�w
6Ҷ�eA�s���Izp.h�i/Y�;x��H�?{,�E]�({C�!�[Mϒ�Ү����3)��g�ט�Xq��.~Czki9M\�ھ+�l7�Ek�*c��-P�ﻤ�E�[���=���E�S���T��ENd'�mgjQ���0�K�n�n	�GS�=�']�^�9Ʈ<%^��O=9�Z8�a�C6��B�e&���k{#A��}�����ЛE��H�o^_�j�l��:ǥ��<�s@2p(*��}�T\�bQ�aK]���}�W���7��W*��om�=4��+)HF.t9:��Y}�l�`�lι�if�В�6�lP]W��qHoߢ=�$��~�ě��Q���N%�)<~���x����+�6��	]��c�G��X�]\���@*����.��0(��F��b4�O��Ώ��_,�2^*���>'���Me6+���h���*�2ךY͒*'(�YF�;����(Bx*��~�y��bk�)�����F���ԪxmJ����׵�J5��Z�݃D�q�:ua�fB�_W�> l��QzH��D1+� �*���7��RfAIJ��X��"t�RU���ϝ_�������<��|��mh�ь�� 5���]��~�����LQy���j�Н��5@n��y�W>��Z\���X���fGH�N���GYbo�4��N7�wv?~[��tjW��Iz�Z�c��4��	tˮx(Q�(X�P��H6q����:v�_%X��muk��]fs�ۭkl%������{�_}�W�����w�މ,շѓ��R1���7,��|��W5|D!�g��g&#3Jr���{���*�Z*�L#;ڛ���Ո�9��ƟJ��.�6��5K6�/J�5�L�|\���0�ٶ)=�����|�+8/1�7pfO�Y]Z���0~�Laޖ�x5G�(�ꪯ����4W�����2�<Go{����[O����HCzq��2�5/'A !'s|����~�
/��|�W_���tJ*.��J�pG�[B���vN7SƔ%�
Z�«�M�~)���h�b����E�wE�S;�;q<��eb��n���"V�>�x%a?^]�k(�n+��})�Gp;T$80�q�����ۄ���!~�����f|�C������������_^�ꮠ7Fe��vk	S���p�1>��Y!Hg��w��a"�Y[���r<73�{�h�C�hf����}a��4u�3��䏤�nxe�D|}��x�=5Fj��9�d��Oro�hVVѠ VÀ9M�j�y��$�C����|k$�9��+��@�x��������0�����
"7tQ��Ôx�-W�gU�f�/|�\\����W�^u�iܱ�*�8��p\��Hv�@�"�҃N�=w\�"�u�q��)o��J��N|��48� �6��r��\�h�tP�i�L�&2�'%�qj��N��@�z�����<x�Cǲ�A�1��){T�ηr%y��덫nu�"�'�#h����5[F��/v*��ɕX�od�~9w������7˻4Q�T�s*��z����Z�|�ߖA��I$�����	���� ����U�X���X�AJ�����3�Њl��;nݩ�j�����	׮���P��n��D���a;��8�qnъk�j5�.�H��K�5Ly�Qu�s��ǵje�`�D`F�s&V#�i�i�N�S�4w#��� �S�Y5��pJ#z��nͻ�۶�-v�v�۾iNH`��a �S LL�2q��H�<l�a1#[Nj����Z�,#�-�&tK!$9n����84���!�h�n�K��I"�֙-1�#��I�G�`B	�T�3�KF�<`�X �
[B��@B�� �����I������0KD��74ԉ����:)m 6�0m����j�y�B�J�{b]��,FԹu�<�������"�<�&~ч~�x��8���#&`��A�뵒��'�;�a���Mq]�6]��`"�V��1����L>��B���Y���qώ+�	�7-��]�a����f�_:���o����f����g��C�V�T'�7�Ñw�#��|E�XD+3ЯX��]0�M-)L��"U{�rM��"����IOް��m	JGr��D]F�*cT���[V��!����FQ7�K����	]u�~�D{��3w�ο�Kݭ̛�����>�<��X�	k}�+n�\��x��pU�^�Vn��ő�u�=V�D��Xj�\;|s��)��lɞ��ю@U�@ř�=�Eҁ#���HCWn^���M�g�,j�ȸ_� ��tVXz����2(�K�J��c�##����+g-`J�X�Ʒ���dH������������?"����J?Z�d#���Yg�w��:�I|ڣ���4mHkeIQs��A��������˩Kq�.w����Ǭ�����1�����x�/*Ｖ��/;�ЮT�+f�T=�،V`��p�n�`&ʒ�SˢN�t�`BX�f���!.�wN�d��mU^Ÿ���yD��i����_>��L�吧{h8�:���F	YP4����1�E�'O�UW�R ;��5��iu6�n$��O9݊h�)�'Η����p���O⊡�!�u�P
k����2Dt�j*�J������R���&�4+�ۻ��>�Ik��/C�-J83J���!��*JT��Z4T'fC��s��p�Y+�L�p���}9��c�~�':ҽI�ݰ�kT��,:VL�7�°���]�h�ć}��DE��|�7
��*�y�h���Ӆ�����{o�;yq�C�:dF;`�ڼ���5�Q.�J���|B�xU��Ʃ�\�;��C�l^pYۓ�B��X�y�C΋��><���g>�\hj����j�a.|�(T܅���a�q��*�h[O���0?=}��y��^��}����f�Q!��Q�:��j��4)@X����ˇp�]ko+�o�X�,N�=�B�����;H̯��ic�l�v� ��߲�'����w���X�t��2��rn�l�
&�:ª��a(����#�Ҏ��9���=1�Z}�zM�
��_��+�����]�op�5��~}d/��S���M�l^��kڞd�[U{�������ք��0
p�r����n���v(�F�)��#����%~�&���կ�`W��|;u���<-��:�Y��ϸ=m�LT�o�z��oΣ�u�ڝG�'��[Z��z�&����'ל̚\�jL,��$��Sк���44��̆T.��������}�(^ɴ-��[zz7R�����9GSV LVF���e̲�̞�����V�}k<�Q��f4�IBͪ�[^�;ִ�E�=�%-��j�Â��WS~��b�u�[}u�*,W/,̦��]L%�d������i��؇^<X��/x�J	:���2+�,t�An&�˷��ߒJ��{���k΅'KH��1q�l��2���������}���+�3�ό�
���-��eJ���ꎿ9R`�S�d,�+��·�N���ְоʎ^�R�2�W�9�ɏ�$�^
�	�ztX_hZ��y��e�#�&\T�ǳ���R�q5#��]�e.4/��Zi�r�t\ѭ:;�+��{�>//QGV8�5��\q��)d����<$�(A���qwy���8w�f���֜,WmI#t��Ü�{��Ąf���a�nk+o�W%Tї3e��*����㠣���Jne����ߒP���O*�J�}��#����]"�����S�r'\j�e��\k<Fq�Z|�O�yޯj@Mq�*��(G�^1[����}9�+��(Nޑ>z2�#�o�L���ޫ;֙�{vT�,�Y�#�,��n.*�k9�V��k7��2L9.9�S�w"YmoG�81_6dP��]�9�rcP�q�įd��u�4�ы�d����sh�
ļUg)P��\�\�k�5��s���YH�5G
��g��l�9�o%>�I���Ub��O6����=�N_ftu�N�H(Λ��z
S%K��r��Ϣ������.�>�u��EOe4xMM�No-��{�[��Ý~�Hhrf.�ݕAV�-P�g��J~n���mvZR\��g��gݏS��=�b��tE�7�Z��=�V:��p^��^"��(�k�ܩK7���5�ɊNx�����q�TFf��u��z����=.=0'C����ݜ�(�	\mה�I�q>iI���
����w}K�]��ho��G�M���K��ݔU4��'\n�U�|<p�4�
��>wدpU�k� �IO3��.��!�`>�I����p�ת9�=�{�ROJ2��^�[V��G蒢��g�{�]+qnIr�+�l)��v^���n�W1ȉ���Ρ%�YZQ#2�֭�B�Z�*갷*�NC��h��/yy+���=��wx�٘AH��>�=��
̾S\�+������f�j^��,�J��e��<�XYp��8-A1+��m��ziÁ�ê"�'	���>[�պ����n�����n��{�G�枧�e}�|Tl��M�"��|���)f�qh��I$�I,9G\�}W�Ŵ�Th�Y�z�b��B/(˫�����#�x���I���X��= 鳛�2ܙ{8"ц�<�6J�՗]��6��7p���s<r���<.>�Y�$M|]K�ի�A�
�;��D�C;R���|:]!q*u�2���-ÜM�h�8�gdy��H���In�bUa��t��پcS��r���.J,��{�R��m��l��-ݟK5wfB���M�)��y�L[ä�E$-��t�H��'��mH��w��31�P��l�.�͊�b�(c��8͕*\\��.K�/*B(Xa4Ц�O`)ǃ������ 5��.IS�2D��Ӫ��UJd&d do]* �Ne&b'%p��� "[�	�52��� ��cl�J�D�MSN�(JneYR�	����q��P؁����@��,nܑD%�q��hF|��w�!(���B���B���|_>� U�޶-9�O�s�۫�4�yi+����xZ[���Qrb⣾{�R���	����o�\9�db<-�\8/֘��Ԕ��Z�o�ޮ�s�E���L1cM�M�s�3E��D���<����a�ಽ�J�I8�*	�%WZU��;R�F����,�ĈK��X�U`���]�����^��Js�8���Qc�My�Eu�3:�7��|����*�T1WxTf�UC�9�g�U��?~vwn=��鲮�"(�!B���\��������n��D%�^-z�fgI�Ҝ�bu� �E��W8w����>��/�g�	���Ɩ)=����5�<*볊�|z+s�޻��Ε͞�8���q���(�t\��:���wҷ���\~�׊#����'�g}�/���y��ջ=([�,Z+"�ӧ��ݟn����P`��85�q�� �{�uT�~��޳^�x��*q�qƑw��O���uX�1�����ε�җZ�xן�c�N�<zLj\T��q����#Չ�}�ٜ�ߎd���:�EO�*Fo�r�Cp�qe���N�5�%��*���P���ߺ�_#�ED�����p��r���;���:B��U��[�£BK�V�9��|������Z�_��L�%��gȜ�/���<M u_��R�u룸�"�$c �ܜ���F/5u��[����Ú���'�r�xvs7��^n8��{�-�y�2��#��i��Pe;��da��Rnɦ���3K|�x��:3Eέ���(FrX�,~��H�� �=mi��j�G<ů9W�f���t�0�k5Ƣ�_wI���[�Ò���atD_�N �ip^�?!5ѴE�Pk�J���m�ǯy����}�jkиzZ]��˟LqFkb����Zx��g�p�G�OG�Pt[g�Lk�i}^{��҄�hB�U�2z�ӣ�G���Ϲ�d��
Ή`Ў5GI��Lڎ/��5醮��;Wv�U�Ѻ���J�L[M
�cz�==�;�HW��u֖x�<ދao�J�ㄞ����]k��-x=��gw�j�x�/]�����޸��i��������h�g((Z4+6�঳3ު����}����J�Ec	3q�N;O���5��ZN�{���/]�Z3r���$��%�Yc�T����9��J,�D�D��5�ىf}�X�[������5P̷�N~G���W�_�/y�%�ߦ��>j�DI%|��}�+�b��5��1}�\3*4d Ϲ���kT�/��]��L��M�Ja��~��w�
˪����r�]Kk���o��t��t����(��.��O�]������#�����ZD��覓�w;�����|vw�ӧ��]��qHZ%|�q�{{�xҳ����Üp�\+{nowWW���4��Vi�]�b�o�O
+���-m_(أ;uW8(B��~v�ѱ^�������l��j�"������!(����/ _y�(Zh��E�ke�?���u�n��H��HG^p�mj%c\Ƨ����}��'�"��Ŷ�����θ��J�iCe�ND^q|j�o����ᇱ�c��X,�Ո�E���{�f8+%t^"q�o�z;1��s/]�gh�N(�Z�ez|M���V.���]�y]8/LWm�1�Ə^sm��~�?C����4���X�r���*�����{�F��8����-?!�dA������{>��ks�
j5���L��^ )S��,8d��q���Ip���rr�_}�ޮ�/��_�r���â�F��P�K��R�t�)?�a�~��/Z��n{�],h�0��V�ׂ�oE2���x�3=:��%E�S\�ٹF�S7����j�w��!1X�8.�6���m�e緜k�0��X%eu��2|)'�|���������xbY.��\��G3Ԝ{�;=ֹ;>��
H�4��u�k���&���|+����E�kN
�no�5{������[�bi�R�Ҽ�tZ��{%��/a��n��]�}�M��Oh ���xL��/��iR�r��9i�?�U[������h�]�*����Hn���W�m��<8PC�s���A������,y��I�C<gZg��l�"�\Ɣa�M�/y�؟6G8ㆋM4Y�Lq�����t���]pqθ��b繗Z��_/��N8XP����A��s�P��V�:GV�"�¼�<Ec\]�+��7�M����<�/ XC]i��B�J��O��JQ�-8WXh�HTץK^���9�v,�ú�gfI�I��PU�s�-L��`��^b�c���ё�#��n���I�#u�h�Jt����\�H�E��!�z#� n�誈������nLg>���t�(�����G�i�����;�I�X���Q��H��5&!H�Tm�=�j�-md�`[�,���tI�o���79�����V��
�g�8c�/2i�Q�?qw�6s��XU4�Ғ��V�ߦ�êڡo��z.q��5��1�=�Y�^�"<,9ƺ'�V���g��p�Rov��X	t[�mX��p�쮶�7���w�r���V��V.��䣾X���)��� >�-g�',�B���ć&#"z��G ��I��	�-H��&���J�}y+����-�� ���XMak�As�iˈt�.6�&�G*�:%���^#�ғ�aɹ�k
�W&��k{ˤ�1f�;�ԝ�Xp��b��r��f_=�X��.7Bm��Y4�g���,�A����y��^��*0�u�I�r��'���yQŎ1��N8+<-0�}��]��=�R���5MP�
J����8�P��7ݕdM�)P��B�^󥎯d���?d��]#���4����p����qO(]���;�i����ϱ��U��\��-����?}�s�t������[ė�^@{��A�t�yI��̉[�ںZoX�ŎGEC�b�L�-�l����S�o���},_p�܀s{u]��	Kz=������s���8<Y�0?;���#0�ś;ʥ�w��;�7׺kS�KYcAѠɝ�v�9�ÊΨY�ӳ����d4�k�ʺ��s�v���K��[6�?F�G���'�֜�d��)�:�.�f���+*�v��ni�495�&�$�d��Ҝ0鱵sG$}�7�\{�ҒEsj�Z�o�k�mT��������*!
+w���"�,�v\x���؝WÂ�+�=�9�� 0�6���5��兼���V=FH�r�)��s��r�/���Χ#��ו�B>�yvj-���zJ��;V�V��N�0��v�}˭�k����{t��<��Kiv�d����cL�y+�v ���S�3���0c��-�wc7/��(��g�RWo�۩�2�+�B��ż�k0�j�t��wJ+ܴ�ĘrA&E�Ґ���(�Ȍ��anl/�ˣ�u�{n���r��@���u�!����ne�c��Դ[]n$�ƟT��m�0�h N4NX����0��$Nm�[�&��M2���(J��*ɥCe��*�/�h B�;I�Sc쩓F)��MZ��e*��4ږ�)!�%�lcG1"V0�!�L ",����j[��8?�Ӽ��OgM��2F�61�E��C���k����$��������l��.��4��u��5ç�����((\���gW=�qu�˿�k�uִS���V�b�yMs/�x�<,�Y�6�k\F�!�s�f�:U��)Ҟ���j���1�ҍ]-9}�*w�sư�-�Vq�^gO*]�Mߦ�P�WQmxG��w��_���E��iE}��#q��ǽ��U���5x�i�81xTOZ���]9���s�Y��:a'K��������Q���9M�VݮX(���7��C�Q�=3eٷS�.���t�����$�jm���t�*N����m+�Sw��y1������xd�%l��+�q^ju��z/N,,��w��n���
����0]ֵֵﻙ�/D��8BphԻ��0r�y�nWl�����&T9�-����Q8L�:���ӂ�z`���k�
ΑZ�v�<���e-8C�U]�'�l�F-Ƃ��2j�.K��x[/M����ܢo;ʹ��3�p?5|i�Ǽ֣�-W���[��"�ۑ*�~=��zU$�2��P��ذ6�j}���V\��k�5�����B�W�����E�7T㠄���5$[tM�������z������_��"����*��ظE,W]�gw����P���G�t������{�[;)�vAp��7Z�4*N�=�7�O���1���s���-%
���-���;ց/[Ri�NۏLw&W��Kyw�+g��k+3*��7�B���q��oZ���{�k�q�k��ұ�
T�E%F���ofy&QՔ�.eLM��Y1B��Z���t��]8���i8F��A�߼����~> Ȏ���Z�P�%R~� �U޴�������d�1}���K���XP�k5���¥���5������[Ŭ�6-޵�Z�D�~�Rg]����B]Fӌ����饷�:�����ƥ׺vrp^(�%
��t���u�ޣ�Қ��OZ�>|�-`��6��~�iRr�b�a8׎:-8��]�]oD��ꮵ�Ʀ��ʹ��!:��L<q��j,X,4Rڒ����Rg��z����͘[ܬ�Y���P��s+^U�"B$T���t�YG�����j*�x�v{/�QA셂
7*?�q�L�U�B���I4�d=�Xx�Y����S\�e_�eU������82��]og������vb�����B��12�������X*9y*�7�n8�5��Q�Y��*�3E�\�Ǽ�+��]|&�^���oov(�I�-D5֮vxM��Eb�=��Wwj�|�:^����m�R�Яwh�|�=�/,zh�x�.-kJ#��Kg��u���|�����'�o�q"�i<��qd��E���W'Ɩp�í�:-[u3��.#�\|Hq�Wbo��;����C���ĩYۋ+��� Z|���A�u��p�r�rKs�r3S��m~�� {>k�#�.N�,UǄ|+~<����da�/$�艗91�'�.�^�]�9R����L���(�_M��ԙ漅�5��%�%]r/zSNs)J�?
��ŋ�x֋|�JT�*��mw�l�[~3k'6����_��|e�Q�ɗ̳�.���0�炜k�	��ʵ>k�E��M�^��Z������9�-��=q����u�=6��^%å�L,�ή��ي�,S`���Nj{���	^q����N�`�X�"�!��s��u�91�S��:g9}����q������>��G(2�e����ݬy���	2H+Zfy���F	��S�/:�~D��=�,�3�o����Q.����Z�v��QQ==6�a��`���ǨW���җ������=�{s�+�OVihJ�h�S�#��j6��~�]4���`��Q��9�_5���e{��,��=a��aK�nU�~kM������g�;=�����M��r0�C�C�۽�s�2Z����b��*�ʭ�tJiP�|s�i8�̿Z��~~�i[�IQ�ы��n>��l��uLf�/��*�U�x����L;i��"��OZ�T֞��{~�j�E��q�grSE
��2��0Z��":�[0g�W�ѝ5.:r��\��.�a�E�.+Q��L��8*�G̼vaι��O
E��)�����8����\)�jƺ�Oe`�E�}I���o��Ш�*Giǅ]jV����_��&�M�/L�3�%�:iz�(J�׫Լ_�(5�.퓮+�%
�wW�Ŧ��Eu�NN�K�=J&��L)ف�������9+�mAh�Ֆcz7���F��	^9H1�|��'˞a��A�
��T׵P��SR,,_�4�5�u]�o���\B-ЁL��K����5�2k��p�Ɨ�;.���t|j�����'��z.*`O���0'��rsiM>Z���q[S��<q�Ҕ]8��w����5��>v�Ů�K�NZRIC �q��N��ݵ��7���7F�D=��L9��uE�A��t�97���)��k�Qc����P�`�;٦x���b�y�Q�u����(�l��֛��mke����oH^M�|oc��D@��&��q��q���=��ة����f&~�����t)8l�{ٹ�JD���>rO\i�o�q"����iq.)
͙�����ѯMO�|�n��F�<�5�n`��V�;��W[۽�t�����I/�Kǂ�xۙu��ø��Q�](AR�3�;����5Y�K��!Y�](~j�^��ن�ep�kӮV�4��+4J���eݮ�j��֘.SS.�z������\���&��13���ok�K3*,�^�+��$A�*��Gf���߳��۶��ʔ�2��^�=��I�F��0i�L����p�O���d�3!ak���u�\�aCa V��9J;{��s2V�����Fm��v�=mïn�4��9p�˽�,k��!��f�_�Tr�T88e���Y��N��k�a=�i���]y͇@��-���hKq�*�1���C�@���JG\-���/J'mNù��e��j� �nP�6�φ��,v�tu�^F��&iܜ�	$�j�7���6z�-6Zlj�J4m��S��ұ��P5ӕ�>�z�l]ٸ��U�d���(�Kc"�4��J�P�.�)*M%IK,�SV�#_k�`�ӎ���p�m��M�0�,��=� bŰW]#~!�	.��D�Zt:����HC���r9�����ц�J8��\͊��M`��Q(1�&�G0�D-�~?T��M�)yt1n���9vG��䴜������m{�w"����ۻ 6�v�}�a57��a0��Q�"��M�Ԓ0*�P�hAHm;�Uv�B�%@��ԇD緝�da�A9��
�rD˙��(ƨ�MM�u�L��!)�)�ܩM�Ge�Q�f!�3ݚ
����|j�j����N�!�M6���beKnG��H@��o�|�0F��X
��"�����]��ɯ�	��������#��t��3�8�K�����@�5���Ϗ_Д�����	�$1'N<*���Å�-��au��vH�d��2���!�&����;�bh��ڧ��a��5��u��8�D`
��;�]u�.T����ƶcgI��O;Ť�� �V�=�wf0G��{rn���i�:a-�O&0虦����Z�:��b�x�,x�E��0��S���J��j�	���p��Ɓv���u��R�hмh�+^���p�U�����t�\;��q��q�-�arwϗ�w9=Ū��&Z��ށ2+�2ǜS����J�:�p�T՝���]:���p�r X)���o�	���ٓ�U��}�-�r�N"<P�*֭S�5鳶�}+�mvg��\��K%B��+��i}�������|~+�M�ь��w����;�F�1Y�[�o4d���{���:�4k�:ٚ��Y<���ǃ�N�����7R��	�B�h���.�}�v���%y:�|�	=��˽��`�"�fK�X����΄A�A6�fɣ}��g�|[�Kｑ"t��fR�}o����;Eaml��g��=O#v	�6��y�6�D�N�ɭ��~�Ƕ��O@**4�
�=�3�6��5�&G��O�Q��x�!�0'��q�qQ�o.pUZ���FM�~x�O΃uHϮ��܎�ܓ:tQ�r@z�&:�`E�/�q3c��p�W���ݫ5k�O��Ռ��M�9h!��*0���~�z,Xy���kx��σ�QpHsu���Q��uf!����Y���ED\�A������<ʽImg<G�X^���G��(ҵ�םH����:����_�T�T��6�P��ܞ�EX�ŝ��ي���0#�dfK�"b�Z����(��vT�L�Ϟ�dd��Q��wVK\��K1ua���R��R;S�X]�eR�$Q�j�
���{�j��y�����ϙ�*7� ��{ݚ2pזoՕ2��޵~��,/�k�Z��}ֈ��3�eY[;|�a��س��QQ��k��hӛ�,]����6"���ms�t=:1�.Bj�ر�SZX8�� �˧��|��1�N���0s����8]c�^��Y�g��+��/�{S�1A�E�m�#�퀐r�9�/��Z'S�f�1v�pc�=Ć{��M��Įt��},Z�2_tw2'�����~U��߿��yI���d��ӹ!�$��\�9�s![����k{�Gc{պ,5�2�%��W�5�Ǜ香n�n��B.��zxԵ���Mc����÷lPw~����WD3�z��aMt�=�rc;.��o@�U�A�'	�v;'ڊ����s�g�vq5�����`�s3q6��ƇM^n^Vc��k��/��rp*��-Wø�7�U�f?��W��NO���&���.��1h�Q�!���V���n�Z���]�v����*+�S5c:�r�8�-o���G({�s�vQU�r6+SK8����yԽ�v�*%v(�5{��Ok��"��u��x�>)�{H��M��GʷڃR������Vw�c��V[�	��.�6n�������K�$Ͳ|m�֒���mw]#}����Xbpİ��X�[���w�B_u�H孜�Rr����Dwn��kG�H��h�qǫׇy{O�ά�@c�`'�}	\/wsш����y���yQ�6ʕ&��ײF�Į.�z�6��Z�d�3����D�l��2��VvY�M9��ޚ��[��i�r[���6�gmN�-��Kb�f�N�o���W��#�����S�N��V3�ؠSf<�ΟLg�s���p�o��Y ��J�O}�&��B܀�z;��"0�'γan���^�� !��:�CQ��h�a��ytA��2���I�#&{ϝ����[�#`��{�n7�׎xowt��A���~�czp��+;��wE��0�Q��:�w��Ei>?.���B����Z��n<!7�ܞ�lW�v�9�r�g9���sY����Wt�9��s�3�R�69',J*'O�}H��F�<V�������^�üR;q"��Y�W��׺�~ ��F��|DP���5Wjq#��nd:ǅ���.�L�ـR2�<F�}& ޕ�bReF���,����
�N,M!�OO(�w@ei<k��J�+�}����!×�Ρht�e�鸊L"�{�+�|��Y[��;������O<mw����{�j6x�@V�\|�ՙPuwu�F��ѫt���ʳ7jwu�34�7�:���H�F!�&^;�8\��w���o��H�ݼ������{yf��s����L51J}����kO����C��ځ�@	I�E��	4�fξ.vi����\yZ8���d䮺����w3
�bT�.�n�F�kQqvM�N��+[�T}R�C\�>�je�K� �
q�0)]���,�,�G�߽��r'a��l��i����.\ۿ8f锬CF0J�+>[� �i[
M0���pd�@q�@��D�����MТm�f�RY��Ś�И�uD�+d�Gp2�@d���)��Q��TP�F@^*���	Q� Uf�����p���h�����9��3K�W�F�e���w�pk�ǚ����5��n\��^CLت�&�Nðd���ǹ�Y �v���uɥZ�٬[�nݬ�N�N����> Id�c���i��b��?T���\�E7M�M&�㉪�r��ƚ2r�+=IR���H��$B$�h p��2�B��� EH��i�R���	9�ŵ*�N��L��l���ђ�K��r�q�*'�<�"���R�NP 7��ci�&����"�[]�%&AC �K�fH�Ҁ$b��vPCTp#��V(Y�vw��i�F����.�q��$/�UU���0���~��[T���z%z�VuQh֣9wh}�nR���&���d�s̼��.��ֻ��e�O�b�D��9��q�'��V��ȳ���/ٽS�4���n��:��5��5�c�g6'oݔ���%�4u�eA�t�-�9^̍�C����o�_�s�v���(�.�OH�pW��ʾ�t��㸖��V�a�Zл����|�z=r)�џ^3�3�^���2~n�3�Iī������➽�{w`�8޻>�f�W����`��q�(�K�5��jiخ�j�n.��Nqm,Ȍ���]bx�����ۮ��W5��j��Ftly��C����ܸ�\KRꈍ�jtp�Y��u^1 �-��'a�i���O��ͷ��u��>�y�%�8d�1(�ԛ�#���<R����Unw?G��Ԑ�;K�������2������؉w�-��.�r�mfpW�Vz6��xj\X��+��_��e�<���ma+3cbo@)�)�6ޙ�ۜ^���ަ�]�b�"�TQ��{�Og[��qV�u�Cܢ���fD}�n����_
StOM����*w�S>X���'}������5�d~lg�J��-`�u����:�<�Y�d9��7HQ�G�$���Rm��U[�{�i���(� �ܹ��=6C�R8�n�gge�'ƻ2�xu{�R�kx�;&%J�aˬ�UF�5f��������f_��Q�k��̅����;�6�Ԉ{eQ,�ֹ*�!��9<��WQ���y!rn��6&�`.�7C�y<%��
�w�q�9�μ,xc����o�ch��yg[�4m��B��ֻSi��;�1�Y;��َ��Mb�iI��UT� ���k�~����5��zϹ�Eʿ.%yS�%�P�/�!v��j1�yݕ���
��*&b�,ɔ����#��r�~�ǈ���\���Q��kFt�YѬ�U�}�{h�>�5�[<J���(q^��NN'�U�u!|;+VP0���'��-o��z���S��2�a�m���JY9x�QVm�#�Nj��L����n�H�\��f$7�D|[��XG�0VvJ�iЗ|��ݷ��"&8�`b�R�����s<��(�=�7�)�L��QMGٞy	��i�*Ӫ����e���:�ɭ�D�3���)0�Wh\�Q�s�O���s����C2�E$����w]se�\&3f%�\vX*߯��*]����s�'j�E�&�w�$����AJ���Z�&�������U��e��Z�Z6��av�>�"���V���;űI=p�}|o�����A��s޴�-���-��Y���2��vї.�v�����%���u���Yկ6)��du<r��0��c���<��(�hv�k�k!��Og���,�cǀ�p��>ٛ�ܒ�p�1g2���0$벊r-��*
��	�^^�;v��H�T]�t��Y���Z��8��Ǯ�F�`���Pd�G��*U�{ވVC�c�����}�dZs]	8z5��������8��v�n��kcڏ7[E<ܣ��l�����i Ҵ�	�}�6�3�eM�q��,���/7�S�$q�t�0���[������2������4vaf ����VQ�g�KT�d�	����^������`Ŧ�˜���vD���O��l�t	�tt����i���}���pv��U\�a+�V��u�q+��,�Ve<�u��&Y�Z�9�ؓ�g���SQjA�K���K9e�n�lS�]�������K�7ra�����ӯ'^n����f����O��g�������bd=6�p��2��Os�13^r�9b,5���;�����s��ڇPT��b�[�Ś�U �j]}�;���~�7g%zF`���::�����H/�=��/�X�#:s)�X$n�n�3f=��[��B.�]"�a�[Z�[��a#P(���Ǧ��W�Y���X|F�dc�X���5N��0���/WS6nO3�����O�:��ٲ<�����]�t�&���4��)B�]y�4�^l�!Ao�V���"��X�+2�n����Ś�]Y2��Z�T���w<=�V�$#�J���Q��ok*gh����t5��;u�]X��u���m�1�z�<[g}5�L��XVgf�l"��_w���{�~G:��:=8��bo��p��؞Oq3�z����r�f�r�z���c�L�0�h2��6�(83+��f42ὐg�����tW5���V�ќ!����ٚ����[�t�`x�����?e�l��{�Xp�n;��y�j�8Ci�c�YN�&�Y��3��Q���u�Bu��]��RpT�O����/�m��[S/�mnӑ�ڛ�:Q�ʵ��{t��2��ɦ�����F\$��Tܙ�^�G84�5ɖٻ�72����-�k����qn�dm1�\��f�f�~֮,��Ot\�G�`x���z6e��M7se:�Ę�`Jl�h*t�c�)=jP [Uz\tܛ�;RI�(.\�!
Ej)$��-��' 	 .�"��-P���6����� bb��М�M��P����������i�!��nI�T55U�M[A��
ۖ�E��`��eJ+�����*i�Ѐm�*$ ���S �Q!(�RІ� m�.�%0&[l���2�A�	 SP�Ьd�.8�`7m0	�)�t.�.�P�hbbpB`&M$�p	[����h!��Ii" ����!K`M�����KV!ʖCtҔ�;)~}^�;��5�!E���:�JM�{��q�}U����r�����;mۑ�"�Ǚ�_���P��*2a��"F��1��BkR*.��}sq�4�D�T�#q��t�^�A�)�=��]������r�Rv���Y]�l�K}�s-�G<��v
��8y��o��.i����I���T��H���F���:���	�35�Arl�-������&&WA�VL�����e�9w]��}�	I9��M��9b؃��Xp����z�T�b^��w�M��R�&�R��ˬ�܄��nww\�	^�ǑO!�3���������Y^�tsg�<=����?Zª$2�ù�f.�\
��ן.�)�^ Z�V�'γ�/�
x��#i�����+�ݦ;�_�
ڃ�hS�3��.j��˺��2.��v������'������o � �Uj���D�Ot&>Ĉ�h2gᴎ��W�֏-�<|��1e�rpr�7}Np�`�\�Lj	]]Vt�3kM�o��˷���5�4e��/vD�˽�:��>���[�"�,*�Tm\s�a�8R�͜�H}��uy����K&���K���_��:o��U���^�6����ޮWXh��+�(�*"�ɗ2�	3,�q)
�7y˻���b�|��	�#�󽃴_)�zb�,��e���aO�o+r��M��V��ŉ�*)7<t��s��6g��[��ܦ̈́��r�u��M�y���sL�p;�4tx�j�O���wv���`e�=^��7�3Y�ǳ|Fiػ7������\1J�q�j��3�({�{6=���^�g.�V�dc���Zl\u�\])^XE9��K���=߽ؐ�a��]UP���}u������@v��>�4���I"#֜��r�O>��s���c�tu�{�7ǖ�=�<�J�K���Qkk�/^^k�l^F�99e��nr%_>{	ޤ��ǈϋƭt�&�`��x�AA��{�7z�lLg
KJ�QuC19Und'�Gqr����S�9��~�\)x('|��\��Y��+��.�+^�'rm�i���0����q��Ѽ�(�a$��u ���WްN~F�0Ezo���\� �{����ʁni���ee�,��ű�uv���VV�*9��[�%�g�{�w�8���(:�=~gL�M~Q�溏������՗
�=�p���ػʀ)(P�A%�nw���M�=��-G;�=�wd�O^��(�J�h9�c���o^(w*�)�3�^�u�ay�;d�����D�S�o3�fia����D����+�kJ��fǞ+�6�I��v<kMz[p�K�-G�{[�}��V��%�d/�Q�eϻ���Wy��#v�Wnu�(��Y�T��1@o�K��{]��]�)t��;|�e�e��w.��ԫ�C{��Y��\5|d��6����"�>�)�y���%�bi��S���� Y��Z��i����g<������ۑ�V�-�W>^��ƆL�۲�**e=͎I�y��?7�Ѳy��fwZܸ�P/ί޵�Ɣ���t,}��M>�7�MA\Ҏ�kX�p�m@��o<<|����y�K��(ُ_g�`��;����8��������:Smv��9��?�ʇ�����\d'�/3U�=UtOmΤ�K޹�y�]%�b1�p��\dO���K���]H�� �׺�e�G��r��Ou}9۱���}�җmƭ� �6	��s�*�[i��4��^��7ڮMĵ���s61'"����(0�r���>�:�������[O���N��PBn�ˌ/��'��7N��F�����Y���I۷��0$u��9.
��Z�Z�4�˜Me�H%JҶn%6a}i.cpi�Ubs�͔�����>ʪ����<�BJ+�'M�;��]����8Z�a��^�R)�~&�u\��_L���<nJ� vdQې�-��|�6p2f�"Wk}��F����/���(�	ZV�q䴕۵z��1�3���)��sba���P�
��z^B�,t�����Ok&B�lUW>H'��t�_�K�^$^����C�z�P��K��9wX���ۥ��Sg����}N��/��y'����;9ݾlħ��CC}�UO�{�:�K۩Sp �m��u���L�Өu{�OJ����23c%�Yz����)S7:k=�B���y������1�B�B\����ںnn��l$x�J�s�n�ḱ57į��>���b�\�X**�G\�CByy+g\�̇_آ|wn�qf���ǯ��Kg�j���ܠ��2*(�w�Y�T�J9$�I$�U,	ѹdQ�s��Ȓ�� O���.�q�6��OHd��Y�:zϋ
7t,��Ό�X�l3n3zp��)�d²�n���N���g(|Y��ٕ���r[�7~���ID/�����1�ǱL��\��^1�g������=\B��۔"t�WW�yI,*T�, v=JI�sC��v�Q����=f���U�}Qb�W���ZP���s|�I5qt֘�GM90I p��*ki�9��[�:�)JF � �L8�wQ(�Sa��S�2!��i�-4�
�P��hP�@Ou�H�E�˒�R A
Z���D+n V�	�9I�LcL�����T��%7�r�`�D��әlT&$D�) ���fx�D� �B�
f�t�+   ��Y�2 !��)��BMM�˂\X�*�R�,���b�� ��T�ºx(�)��Z��T�!1����Pㆈ�� ���R2�je��J X$�!*o2�w��MQF��z�l<VI�A	�-H���Ţ�����lY�6�����r�FdLƫ<GZZ/���Weq�k��S�ۃ��x��Ř�o6:��y�e�< �D���� �:���,�r5kr8ޫ�j�.qpz��<[{���t��%�{,T�� �������=�r.���v��V��x���1s�j1���؝�V�v�@���Gߗ�~4���!�͏K�1�rI`Eи8�b�ߠ4L���|]FGu�5v
P28[c����y#�XE��/�3�̢�ޣ۸h��P����NQP���&�CUgoV_c�p�$��.Kb��9��9�Gɖ0�bv
�LC�xm�P���~]jՍ �nsU�!L��I�HQ���B\k`+�d�������u8���e��*�j�Om�Â�>� *
��s:��}=�8ՙ�ڀ�ڂ#�1��cs9�,�:~������?�x��ܯз�ɾ�*S耇���O����B���Op4(����s�!-@q&�*���Ri��6�p�����!.n2=<��т��ڦ"���	�.W+^x�����Knϼ]�ْYW�F���OJ�6��+�-���s����5u7�p�|9���l�"H���1o��.7y��{�����b�Ru�m�_o=An�D���}��{ϧ�{����[Y�;cn�XǁU��ů�I=�4h�~m�^N�M�P+�}ۺF?w[����b���f����dr��RJ��ɖ�����+-#�zѰ]�^�f����S�2�~Kt�;܌Y�{n�B�^��bs>%]�/k�n�;�����h��W�w3юo��/Şq�u@�xq�q9ts��pl��{��Ǖ�#����+8�Ol3��_&$���������7#�@ҽKa�b�bK��2�Z.��Ď�b�#����w[W�+��N`��a��m+���Ga�Vz��by	S�&�5�ҥW��޸U��~�~Rn)(��<c�Q��xYQ-��"��!���e,�^j���"���oH�CM��K�b����=�"�/���%X�}�c����7�'�o���dXK�NRBDe�.M2ȋ���N,;������Pϧ��h�1#m���Q����}��,FҞ��vb��Y�,G�����o�Va�h��][i�Mjȝ��XP{=��ݭ,0�E�K�[ͭ���=�od^�E�G=���':�c�~�Ȳ���������7��s�x�9�B���u�g�X}~n���x��e{/����a�u�t��udB��Ĩo9I9X%�ǵ�#F�V�ޡ"C�qg>l��!l}�U<5]g;BI�bX7���85�9�D�ǾK>V,{:$��pYڎ�t�U�{O�sQi�-������`>�&��tLo|ф?�S:uI��+��U��j��������5v���Xq�o�?2����lٽ{�ǻ�yu�X[�<^Q�/�p'�bVfř��r/۾W2��d�ڔݩ�@&�dq�%,�jT���?U. L����q�����K
J�������b<���gp�@M}��yx<��˰U�!�f�y�4�����`~d,|$̹�\��q�'��A�A���pe�#��uar��'ܯ����߆`��=����š�U?�<=��%��afjӔmO;�}��kEw�I�{��<Ժ���k�pT��%ؤ�N��@��ܮZSe+��H�����=������Ƽj�⓯Ey6�/,Ľ`�m�CcD�Q�s���f�;Z�N�8J��;��J�')�pw���kܲ|�*��ЮJ��ҍ4���!wbk�Έ�Z��Xj-�D��ʣa��L�Ǹ�sF�a�=��2b:[�j�/5�yM���~��U>��[Չ�<��e��i�oA�[�p�AL�3�މ���RY�3�vJ�;	��Y��A��7_���N
�kUq�|��<��O�������w���O+%	h�m��ף�F[1nr'Xade˅ŝԫ�YT�(�qw����F��mx�Ŕ���+}�Wݷ�w�g������C�]i\�~Z�=g�Wq��i�bT
+��SfVvC����,N'��a�f�"���g�c�y� �=Đ�I$$�}�T�)iG��)��F���
tޏ�$���Lj�5�v��>}��.bہ��A#����SZ(��4�����/��������apik���F�DS� �ۊ�	�wc�����m��_�[!�yܖ<�6�����&����"�w�Է�q�K�+x���( ��i������@ p��PAO� �S�'��%-�i����΃�?�� �G邏ϵ������}}Ϡ����Q����g�판z�ۏ��aL{2��3����l��Z+_��
�u��q��| |�Lu;��gߖ�z/��"�� �s���j�X!.")��0�� �e��h�X�E�[����y�N�����(�
vr�^�?Zy8�<��~G��t�I��)�`;�d.�1��u~�C*�9�c/v��syG��,&H@�#Se2�'=)�
/��zZ�<�9�S�Ԓ`p�����ϫ��	0�+�?�����u�!�3�{~G���=A;�Y3^/�d_��֜:�!�%�xG�K�*�)�Y���
���H�s�OJ*R�Xo��+����р�N��2wYS!���HF#f�𠟡��(

F.
_#�2��[�Rf�*��g
y!����%Ro�/���`�y���|��DR_�=�~�Rw���<�~�4��)���Pf�SċqTA�����bx��������O�>���K��c����%�
z����x�����=>��I���
R�0�3M���O�����}��x�|A������9Y!�|(�@��{+Ӻ>K���a���?g����i�;�<Lw{���
{}g��ߴ8��In��\�h�ǀ��{�P��C��j8�漴`.-ޘW��xA"� ��`�;|�ǈ/��������w��
{���z@�_�C��ˌ3-.��8��g�k`�w�XC�JWӮ��������)��0�0