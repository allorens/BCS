BZh91AY&SY��^�9߀@q����� ?���bR��         ��R��mm���EI!T[h$(U�61� �E(��m��P ��k�T(E%mk!�l*R*Z(]V�tٵ�3m��b����6�TV�HH�*՛L"٨�KeV��Q�b�mijm$�ml-�cjI�)P�J�ڙlRѠn� ��w�m6�F�X-�Vi���65Vִ��d�&�D�ق���j�Ae����[j� [+4
�)��U(�A�4B	!f�5�Y��f�[���V�j[�@  IӾU@W&������ Q�[S� �d�kZcv�C�WT#vTu6�*��f�GA�Uܮ�t�V�Y�bʤ͠�[4�
�/   �۵5���Q�8�e �e�z*�U�E�=(PN�ox(@#���t�l������J �s{΀�Q֓�^� ���T%AI�k&�f�li��   ����h*��x �z���J��y��� ;U�< ��<�
� ^/;Б� 7���G�U�x{h����z(��m�fl�IVcV��)A+��  n� � ��^�xz$=��T ���y��P
�v{ޞ�*�y��d�r��xh�A����UD�z���( W��^��SJ���T(]�Z�m�̥D*��r�:
 ���z

 �{^�@�z��  ���� ����:  �^oxyR�j
��{=* 
�x��� +� tIGWT�)�ICF��4(�   �� ֛���<�Q%.y�xu@*���{�  ����{C =��=á�F�������
��W� ����� mw�wxwa�WA�T�[$�F��m�kl��  n� �l9΅�`wp�G��v{ƅ �9��]i�{��� z��
P-v� �� 
�/n(�8;mV�2֖͛V�Z�H�   �yP+�Pm�� � g� iwjq�����@Ks8�g����c�� ZUҐ�Mjؖ"SY��Ec�  w�@��\�
�+@���:�.9s��Q��e�@�6�8
 M�'# Kn��� �Rvi�ڳ��"K,��� � S��
�{�n :)�.�Cs� H��
�րиLu��I��ʲvV�]��Jx  �  �j��Lʥ*�0 44�� 5Oh1JJ� h4   h �&B����      T�UMT`      I��2y4�h�@M0$�$j"�4���L�M  ���-L��)K(1lrv�N���k�����Z����/�~C�|����?.���!BI�B@���	$ C��HI?�~��BI�&�������������iNH�@���Y��*�H@����O�C�hd�		'?��_���4I�����$�@����tH�FN��td��ѓ�A�D�: t@��蓣�D�:0: t@����=t`Q����C�!чtd��ѓFN�:2t`tHtI��'FL:0:0: td�����M:$:0: tI�'�N��4d���tHtd��ѓ��tBQ���tHt`tHt`tg����FM tHt`td��d��蓣FN���0N�N�N��FN��#ѓ�D�FD�: tQ��C�!�!��D�Ft`t`t`tHtd������tAt@蓣'FN�:0: t`td蓢�D�����Htd:0:$:2=:(�ш�D�:2td���'FN�D:$��ѓ�:$����:0����'FN��� t@����FN����Q'FD���: z$:0��'FFFC�C���$����'D���N���萁ђ�	� DBф�BD��@���BN�HB@���	!с!р�J�D��F���$� HH������I�N��C�F� �N�:0�:$�8 HtH���� tH�tH���Iђ��!��B tB@�� td�:2�I �� tatB@����ф�$�� ��:$�tI td$:0�:$�:0 ��FC�	!ѐ�$'F@�F�@:2@<:2:!tHHtd$:0�pa'F�FBC�I� 'F��BI�$�2 tI	:! : �� tH x2@�� @�'D tBI�N� :0$: Iс�	F:2@�!:2 �'�$��N� : `�I�$���  :2 x0�:0tBI�!&N�HN���tI ��!'D!:0 脁�C�$��	<рD�!$�âFD�:$���'D��d�蓢N��td蓣'FN�0gD�t@蓢�FD�0�@�ѓ��O�:2t@����&��t@�ѓ�t@�ɂN�:$蓢C��JJ2td蓣'D�: ta�'FN��:$:2td蓢N�:2td�:2td���FN��:$�âD�N�: tIчD�t@�âN��:3FtIѓ���td�ã'D�tI�'D�tetd蓣'Ga������;����N��~[�s�%���(�(˰�i������+J&��-�Ƙͽݖee�
,3	��[,m��^B�h0�^M��ʵ��%�vK]*�mJ�	:��\��mU�M��<7�U
3Fl� ��M=p*�&\GTƭmm�6����K��̡WWKŌ��J�����2lb6R�T��\b���ۘm�Iۨp���dn�xE��#ɬ�VeZ�%K���ikfC-C���&�Y�bI��X�YV`�{��6�Ej����f�e�l%�{MU��?��k�kni�"�f�F�#J����le�eര���(#��-�0�1w���Ļ�v.a�k!֒}�n���Ky�����`�%�{/�a�Ic��)��z��D��#��5��Ce��dI{������&̗l7��6^U�s1z��r�v#W4���˒�Ueea�R�M��IWrdE�ٴ8PN��Y���Ջ��vU���1��t[R��@F!�פI����N���Dم�.G�x���\ʕ�v���4Zm�$]$o��a*�lP[����	ӁeV��Ù�%����C!�yp���OL{x��v�֩R J��� !bG�m�k6��e-�[�f���Dd��ڔe�zf�רY��A����!�^�����s$�)�.�\����X�[����RZZ�!1!�a)�GV):jm)��/7s	vn��R^ �nGz��!�e^��#5�j\{�hS��P�S[/r,Z�4�ã)��0:�v���[��1H�ML�A�%p7md��bg�Aǒj�[Ys6J�`��n���b���P��]@�nM�D��
m3$R7NM	��9�����0�S�[ٖ�3tn��;m�R��
��w�!Ӫ][�E�U3�݂���;�G&�5��d7��Gd���rT#w`WG2՜ǹNd{E�"����{�LE����٤C��^��3l�:Z�/v�qG��7p�ITT7�.�6r�Y4c���Y�#��(n�hOv�Nh�1&v�-�b�5(��nlz�8��5�!هR���М1K��l�+(���F��Y�bd{RYW,�-�5tm�h[���m�F�,���FEF�ȠGQ�oaI��0E삙G��CXMU�"����nإ�u��J��m��F�9H��5�VR���v������̴�����yx̷�C%��%�e�'���/X[zd�j�Y�b��v��t��/˕�M��f![v+cfV�ѻ�aٺ�;j��6�&E��^kmI��m��\%��:�����ԛL]'Ak���du��d�ɉ��ǻ�����Ek�P�k*\۵A��U��5��0�.��ڐ�*YR�t�q�rZPF��phV��\YZ�lͭYCf�潬I���2wv��9�gvŦZ32�{2\�(���{`ފZq������b�I���V1-'�5���ͺ�l�r*"�e��z���Ng��Y�4�5u�5�Y��9z�osf	��)+a��h�K"";.�0���t�y��2^��)��6�@���Ȝ`CRCv�eeC+p��A���bE	NHo"7���h�mV�+'�i�1�j���ҍ����E-��]�v�Pj�M(��Av�ǉ֨F�XC3v4q��jn��W2����T���j��"�FV���)�4\�C��*`��I�xe�@�:cZF�Z/M$ʓF�
D���y�(1Y�@c��#~���x�1�ϱ��e�E��u!����nC�V����X�k�#�1��z�A�(�AT�D�D�QL7��*�HkhJ:s@�=�W�$+4F�͠LP-�;�
;twI���äSq#��R������wyx1 A��̚۹��]��w$&��v(Bh��U�A3��Ii�7�<�������քe��2�˛��VI��;G
��n]�0��0F�8��w����Xm]��nHF���+M
yvl5x��?Q�/$�W���Ѝ�����E�n�1��ݩ�'��P�h ��2m�x$	MI��'!��KT]���
���Ʈ;�Q�kb�x"�/*��x��t�F�oeسڔ�+��]�]YŘ�L���m=Z��v{:݋�oh���[b�Tm^�* ����(�X#2��vl_����+Pl0�["�����y�wJe˵&�O$$1��a�Cy77m�)m��˩���Kum(�ԹO"Z�i5��K�xU�3n�ts3h����ܭ���5������f��YLiD���"��^��ƭ;8�E�47Zԛ�ac�w�������k4��ۖ�\�]:��� �呑�`ȣ�:Hl뻲�͆�m�i;�K���b+��B�bw��<z��v�{H�����U���*X����	��!w��:Me�,����1����Ê
FB�nS3؅H�1�%��$i��_��7
�˒m���Ê���y�@�T{��^mn�T�N��[&��%��e�k�ke��y(��-`$�������p\0U�0yZ�iҷtP��r�bv�b��l7[a�H�BUчuMx^*�Sc2����7Rj���k/z[&�ۛhV�Rj�rn����tɭ��񋳮T��4m9�+�YO������Ԥ�[W���Mk�1+�t_�=9r��X),��rsn��z�=;�!�Wj�dD�j����0�D�a.�7��0�Y{Zu���F6��Z'��6�V�[`�{���6�X��r� �ԟ�^��49Z+!9X�
��h����mI�(Q��Qؘ*+JTˠ&J4�)V1-ԳM0����� djQ�Z�^p��ڔ��z`؍7��v2G)�u�i�$��3�y�R�6,����ǫF�w�Mڻqs�J���>�@br��6p�ΥW�	�n1xo)�Sr`z�QT漥ev��(iT�o#���\���7���U�I�.�Jt� y��m�i%�Ǣ�:k	r�7,XzΊ��4j��SH���G�!� �ll;�H[ycc��W	��H�1^����%�k�l�w��ͬ��\˧6���2ۼ���L�CI�L����݊u�)�B �q=1����9H-ŭ����P�J�X��&E	��t����#Q���j�Rہ
�9�ǎ��Z.���nʤ�X�[�/w����X���N�E�	Y,���Y{���:2���h	���f`�!hTTD��<�n�f��;���#]�5q�(�)���{22��w�Y�q�+a6��5V���F�kN�ʗ������S����@���`J�����m�� ��eG�^��eɧ(���JOƳX7�w*jl���,e[�{�,��?&�^�
=)�/t9,�뭓tw6'vS�е���M���҉�0˔kDĮ�YQ�1�[ՙ�m��a�V9�/.8Ց"�.��m��4�naYXn*G!\�Z���X΂�i�WY�k9h�2%h��Ne'�I9���1\C8�щ�5�52��wq��[`����m��,ֹCc+1�~�X���ڼ%Ǒ���*j�0��rM�i�Ay�KX�'R^�(ܧ�X]*z������6g�����#V��Z�Õ&�x0a�3uDXt�3YA�p��������+�6���G�Ҽ��3^����$��2����%�F�7�.�3V]`�Y(�W�Q��e5�K|i1�eil2�j��76e����h�6�%Ŕ��i�-yn*���w (,52^��b����k�����Z P��2|e8$ɚ����Y{��6ݤ�42��l�a�ڬ����0#��(f,[��D�dz��e�MU~kr9��=.�Mu�+�{Z6*�JTi���oVctkf�2f
 ö:F��W2!R�ԗ25�ic�(����r��ec[�[�_����OL��KX�$�*εES�RZx!�[�o,��ʍ5����K��N��$�X�r[��Z�3̸�QX.��Tr�Lш�F㗥�l�ȝTd�lf1љUe��n�V�� ���<Ou�s"�L˭$j���p�)«du��X��M�R;�
KZ3NgS�f�噬=�z�˖&�{~�C[0�f���	�����[lG[�Iz#Z�I���E1/��a� �2ʴ�S�Fp��Vwn�䳏)�҄�!��j1��V�7]d`-U���v�^7����&��z�ZO��;�]Y�x�(\�
��:��}N�-۬x�`(��Uj�6�)��`���A��#��	�B�;���z�bX����J�r
Ry�r�HwPȖE���g;��O(��w�]�#��k��cr&u��S��k.�i�-�*�4�< �[�:��F��^ev�^�ͩ�z �W�%֬W��L�GW�T5k��0L�-�y���!ֻ��2K�C.��WDj��ic��b�	�D�'FD36KlQ�VN�V�������f���/IFثsh�w�1kboU��.ʳ�� jl�mL1���jJjʪ�r�!��Bq:h�H6�l!Gxv�+��L�d��5�CK�,ؤ��襯*�������YcLˆ�l�-e��2fe�U��dבcW�����l�7�L�M^乳u���e�`&H�U�Q4��oX�7)=�����C4S�v֙d��̣&�mo��A�¥�q���¬�U�����T���d�B+�Ь�2͒�fz�d�˭�9�0�V<��5Cn�0�M�����T3we�c!I�y�����h暶��+2���㮢�����)��I����F,bx�[���M��vm�BJ,n[aSW0bh��G42nj�(��F$�d˩0 /U����ՍAc�S*��(3L]��:&a��A�W�Iz	����D�sc����9W���az�fS���R�f$MS�aY���d��-�2]"7wS����-[�1�ܳ��	���͔M�m��i��a�)�������oU���mL�ku&V73oT�J˓M�YVJsZZō�B{[�e��vɶ��ƅ'z�ձ��x�JҤ�c8Fb�̦޽U�R;6�U�5�bm��~�;���Ɍ+-����uf��&)���bQݍCsi��N��M�yU�bVӁ������ZUV�pK0d��R���ӎ�ŷ�j#�ol�yb��C��BU�P3Z�*�{����v����KXF��&��p��7.I����%*�2lQfm��%;۔,A!�)��A��&s1e�iZ��A5�7��Ci��AyW�;	M�I��6�:�a��ku�j��_#�Gf��-��nӥ���6�D70���rmm���m�N٧�j�D�I0K4"�5=�UXÄ��F��cU�w��n��kI�c^���HY�j�H+F�kl�;��.�2l�H�F6e1{N�!\V̅��;z��5�.�q)��L� O�j�<Vq��h��]�r[�ݷ.Ź]�=��o�wS�5Y8����hS���k+
�rم"�m0iM30�
,�G2Q��=*V����aǔ��ҥ��	r����ٖ]�:�l��8lݣ+���n���`��B������#�6X��,�*ix���K���2��u/��MC�uH髚٣.U�)X��6Η'�,@ٻ�<򍅙���:o@�� �ѷulq��|9�e�Wr679����j�T�&;�֬ˣIkIY�Vr5i�1�4�3��D�Ă1:�7����3C.Ζ;HVGB�lA$�v���\s1�z�a͊6�	�� �aZX�z��H�	�3�@��L�|�QP��,Zp"��D�ޢ�ٔ��o(^��tsr1z��f�c�p{k��b�g��n�V+1(�潨(�Tڛ2+y2��0�;)[ݕ���w,���V�WqR�%�(��K���JȫfR�h1��2Ӕ�ź7Y�������9J�"͉[i	75�ߦ�N�,\^��3��\A7���4���8�l�ˢ%�J�L�*�r	�{.�r��oj77bC͛�V�`Uz�.
�n�=Th�1�30f/՗5ۇ*b�E��ek#x[s,P)e�ٹ%
lf^��M� ��6�4��x���/�����*W�y��%!ʬ-��ZT5��h�FnѤBׄ1�/\�2�n*�at��G4�R[�vh4�ꘋO+@!���d����h�y2q�"����2��2,{q�X��vƦv�Q�@M�w�1�b����uջx�l�a��K{]�Wo�ȧ�E`}�1G�N�a����Zk:(�8Ȇ��T�@,�s�f͵�`�5E�[7Z�M�g������K*V�aQv������ܝ�����5�M���E@��0���e曊P�E���gt4�2;@��V�61a+r�&��f�%�̈�b�1�CG���"-�Æ���m � AW�����R�}&n�A�G���	v4 E�}j��� ��C�p
�� 1��jA��V�`Łw��n�]�@c1�`d�dc�hK.�0V��Ac�2��[5��,�f�х�1j�I'/0�H�h�C�17��1BM�I�e��A^-WY�q��U�㯏�k�ǫ��ƹ�m�5�Ac�P�-{�(�Mk���c*��q��\<K���z��@{Cx�H�������,L��mٺ�R8�8}�9���wUc�E�,z����
Cm#Wm�b�hX���.�7�I��dpT�*D�4wk�g �B�~�����̈<���k���<�0�ю�*����z,`�� �4A��,`z���>W��wfL�8зz�(��Jm9Q��M*m��7pe�@Se����A	 Lp`Z����>Rm�?��o�
rg�����	���@���oc3��7# 掫/z�u��P��,�7v��K.zعu/"y��cWL͂5�6�:(�J��k��E֌�q�M�7�!��Z�9�+ؗ���ݣќ��Nv�z�TQk���J�5�ag�kZ$�z�sM��o)�QM�������W5vc����Δ�t�ÕJ��U�e�YU�R�����.�nA[�K �b�Y8��6�=�y'ZS<D�<��	�Ԝa�7�w7���qU@��,E]T�l�9+�V�s���k���IM�8�Sq�Ʃ�Y$��J]r�������+�P�]xoW:�T�v�Ԉ9)�`�-��v��wע��Eܭ6�HJv��a��+qeK�X2H�%��T����hei�j��]�/(�TN* �pb�99��ղ>�ӛ���H�3���E�i�# �d���ud�������N����ݠl�$�d���`#n�!R_�ِՈ�QF!q�G������"�����o���RӾܕF�wrR�>�;�E�G��{��
�j`̕S�y�f�n�(d�.tM�e@7��4w\Ҋ[�-���nW;�9KB�tr��Y�yݶ�[�� ��]a�4�e�vG��Uw:曉�:B_23Uy�*ނ��ڑ����Q�6���w#�*�6q'e�B<����E�n;,e=[��Y,�,�Y��ж5�����\!÷�*�ս���'���t4��ᛷ1]���u�ڂΙ'c����l�v��H8�6�m���r����l����v��K5/�4��cz�#xﳔ]'
��bj��U�s
`��z�)ν/s �����Д�g�w]K8����&��1�^�*#��n�n� �[�t��5����"\����P��Y٫;wP��PG���3c���ʊPҰ�u5����v"������o����ӷ��z�f�u�s	����duu��͇X%w� ��Z݈��M���NoP�YN']Ms$WpnPSA#�S�"L�O��Qu��u/f�N�p�ାU%�3���79�cr�3�9��4ܙ;.�]�Q��kX�M��I����l�Pv�7F��л��&�P'Wd��-�ׄ��{|�1���/��ru`y����y�'7t%ɮ^�*L��&��u�l��VR9k2�LۏR��ǆjåu� ��ҳ�A�r����QM���"ή��[le�7�X�Ž�Lӗ�ꓩ���ǔ���nQ0Q�s3]�Mͫ
I.��$�Y3k�����6��7x�ܨE��Z5f+2�C�/�XS|�L��+j��<�q�Wz37l;�:̨�1zS��6�����h���XoH�p.y�6t�E�]1~1�u�/b�wɇQ���k��ٙ����b����u�7�r�NG;�6
,5*��:U�l�jZx�N�SH�Mǡs�O�GT ����X���q4���7}��;������&�w&����ݸ��N��ƺ��g�1��ᄻ���,��f�7��ܛ�^�;�1P�TU���KJ�Ū:����K1��U'4�ֹm	+��;!�m���iCA�ۥ���{N��)�� x�	�����ѣjLEJ�ҍ���\(dt�}z!�^M�ʦ~�q��Uf��v�%�Ѣ���܍C�6s!U�f�O�ѧӍ�MIN����n�qmk����� �^���b��6�d3o�G3'P�C�B���m��O��Ǳ��I��f�9N�ּ4�����X��t/@�+)����Y��q���zx��/'������T����^5\[�yC�U�H���❕³��IK����b����	d����*�O�-YcpJ�̬���6O1��"v�x�ҹqDr뮚x��o)�7u�|��o��t��K"�c`�)p�Q��ջ30H�,���Э�D\9*��S�RS�2�ei�"�6gG�"�֦�,�"F�R�[u��{xl֘nܸ�%�u4�{n����s8��1[�v���,K׭�n�]Eͥ㚨�3q�W[�Nk;Q�ʝ��Vkڂc��gYՀ�A�֞���B��rX�6��[��xH+qi�p>�I��|�;�\'l����3&������]�C�6��&L�Y�pbǴ_=�_,���ϸHb��L�\9g�Xs\g:!�����d�~��q�����_[�ٿ'�AP֘W.���0�׵0�'Uٮ܅�ڄ=�����|!���_aO��6	+�[ao�P��oҁP�LM��.��u#M*Kibׂ�t���omU�R�d<-c�ɗ|�֚���o(�����/3뒵vh�m�!ʃ]�]�&Mܙ[���H��+b��9VE�j�ۥ�;r�k�5�*�K��s�*N�S9u�<E�c%�j���y�/n�oZ��9~�g^s��ےܷn��@���Lo�v�ԝ�Nx�s:�I&I������)'^�ѷO2�U���̖�����t�2����u���;^�M���JoG��w���v{�羁�LD��1�e؛��m^t�.#QE}#��X[��n~��(G�	� ��� wu�jI�ِ;e���er������/�uP,�|�,��L�ûu�|���ދ;dX5�kG"�[�_^��*u�c��{�>�i�R�=����F������ރ�\U�h=u�� ��Q���
aK6���1K�D�e�T��B��ݑݢ:����	�9Q��:HJ�a�lŁga�I�6�J���E�T|����m����y�뮆71�洦Q��v��,����J�/-C�؎���y�yf�&����V���iS���y��[���v	��<b8����FI�����*aPT��n�����'
Cr�kpM�c=l_Ye�u�1�i��L�I�q���2��
5i���@�:�
1TYi_P���C6�L�%+ގ`_+�kT��Y���1'�����;iN�G3Vf
�sj��e']�}]� �+��leY����s�$�Y2y�ֻ��em�{8V���9���([z��tU�S�����cu���ے�Ij�E��,�q,��QٳWl�vH�>ܧ`K�%M6������؟R�s��X��U��m�t���oAp[�n��㋂{�w�*S��Av��ZNp�؃��GT��6
�n�]#YR��ufq�J&CVn#a�A�0@e0�U�w7�ڼ��y�W;�*U�в�)�"�z��7x�J�����{���;4�)vkq,Z��o1ᏺ:�(�)ݿ5mkZw����:̛W���R�l3sT����g9�9�YVEݱ{p1��/�;&V�D�wy&n��Zci�̕s/�%�/�
n(�aojA�@i�l� �e�Z!��Ɋ1�/�W7�ĝ��q9�&\V9 �`�������D�6�n��%D��[wS&�T�n!��|��+r۵ԭ�˧1f��2�L���ea�d��N�A�ST���i�]2�5/���^r�(�I|��"�s���S4�N0fe����6������^��lJNt�8��pU��\U؀b�]��@��1uPh�R:õ���t��vv��ĜYx�2��2r$�\}�����/�W�m���9SR��h]2*8��ycsjcŻ0�g���M�W�6��/b�.��n����E';L��t���F�sM���V����+g[}	����hҜ!�c|.99�.��;���Ү[x�#cF���ώ���hNv%z��(�ԙ���VV��ɠ���چ��]g(�i�@�����f\�T�9�V��W*�st&pi.��0<t��N0�؅*«Z<�]�c�dYd=�Rp^
�V��������w�u�Z�l<���ٱ5���h��L���K�5u<W���M�1\�,�r�ɩ%K���~����kJa�7�v�2m&�8��gw*�N�k�׉[䳁�8й u�dw�����͍Ale�S���y�j�ӹک�|n
����:NÌ���:�N$��)K�u�b��2�:��MYǩM{K=c��I����3���	H��2�c�s�s�ʙ{$�]E�L�A�]��E�}P�v1�W��MVX2��=�[Y�qƺru2od�'T�Z��ޤ���f����R��k��+V���9��dn�ϳG!WS�XWfj�n@�E�qSi���˴�u�n�Jrr�]�Mu7�u��w������]�Ze����ٛ�����j!��>7�m�3Z��Řґ�nT��s��W.��Q���p=���)��2�=}x�t�;2������=�ϧ*Vݧ{�
]r�Ro2�3�v��0��M���p�z%�Un;�҈����3ӄ�*�Գ�zT巙���M[��t5�_��\�<�]�!Yv�>`o{���i�o��ɋiԊef���-O�AH��f��k=��U$��.�mڧ.�V�<�k��IQMڭ�sb�S�u�����PO\�04B}o�`��\,w�mm�W6�,����p�9�VhY�wY֫�*}l8*R�l�cl�S�La~w[vT���E�6¼��uy����k�S`H�h���]W&�Ǐ¯�¬��'��t|�oQ���Zj�!�Cr�e)�t���ۂF�}��[��*F&�_W:�X��A��[�L�f֧�:
�),�#���`]T9������5�b�V�u�Ğ�i���c�r��A��p�q�NY�x���%�wV�!��]�ˋ���~ęe<��^,볎��+熞���F��W[�=$�p�}��hruµv�S3��b�M���]�zk(��v�NE�Σ�p����H�p���ƸTb6��vA�b��1{X��r��t�&y��_�ʭ���t-��lM��4��eci�l���R����wgoH[Y�n;��3�3���|[W�싆�{�՜�\�St��VDycq&p0�u7��g���Gn���l1Z2��+��ު�}�qE1�@�Zk�GM�Cضz�ap�6�eD=Ђf�,^�c�oY�ڒ���wۮ��vB+s�	��|(),��tqv���E�����*�h����ѹ���Y���kln���ir�%��by�g@�pQ]�U�R��s��wy����x���*���+N;�C#�h�!�k[!�ӹq`�zxi-�U�7�:]Y�s�Dc�P��k6��hF�>��d��#ʤd�I%��m�;�_-2�l\�(�-(��=5�"o*�r���Y �!�Rh�_{�1��q��	�%`ڴ'��gJ��Z��JČ�3��J�eV�ܔS���iW|Q�[sF�;�㗙U��� ��6k�]�BI���;�Q��/�`ol���T���wLy��`�X�\u���J;1�T��,����8�pW���;�7(��
��[�����`SCw֥<7={��u��U�$��ں%E�ַx��('G�/k�+;P�_.�#�c2N��VC�&����!hW
9]�� w���6��z5�Z�8�`��*j<��w�X<A�rm��дJ�֨�u ��ٲ�N��p�D�~郤����W�,��[j����S�9��Z�=����^���W�Ԭ��&�r��aR]�nCe����\�����ܹ�U�s�H|C߸�"��9�U�����k�GE��S�JAZ�{2��;zIϰ�3D�ss:q9��.8��Ӿ�%�gQ���46h�Ż�A�HZ�u������XU{�z����Lv�=���7*��������W���xS�t[T���/�Y@�a海9�٪K��j�4���*�j|��JV�J�Y���SIgF�Q������f�..O���4���}m
�.��OO��]�5}���|u��|�^A/,�W�[�c�X}����l��WV^������Î������Ψu�
)|B�S�yʹd+kR{Ve�:T�.��
с�G0"�LIoN��J.uϬ]�X��!��@��)��z˗��ñ˾�����L&5�r#�����9N��r!9�zs��z0�{.Wr)�ǤDa4֪Fhʔ����W�����q�N�2�U�Tr{�s�1.�Z�:X�eR�vrs�h�o6��](�0?U�(S��n�ÝX�P���P�!���(�q�'\����%�x��Q��W^�6���6�z��V��Je��XwA'�br��!sS^��Mga�Oa8��ܑފ�C2�WZ�M�T�j�t�V�}.�)��fҎ�Fd�\M!9���
���3�}6pd�:�msA��ّSj�reG�H��1ɲI+L�#�OsL[�$Ī��6�tybJ�V9P�^޺R�T������ڇf��\�m8���E'N���O;o�����C�)ɳ3���\\�;�6�[&�;c�B׷�[(���6ڥ}���ܲ�)�&	�g#�QI�;���Ů��xOv��
�%[ku��Ym�u�+U�Zi��o�w�L�{e_�K]k�1��e��n�$� �.�f�����jn�0������H�*S��,�Qe��UJ�P�Qp�#5H �����a~-�\�oh����a�Z.�q����*���	�Z�z���,\�j�Ga�i"�ӽu��$�&�Q
�
������F�p��!�h-/����5_�XҸs�M���A"�l�6���ۍ����Q)I�P�m�_�����%X_��!S?�Q�a���(�Q�&;��$��Id�08�0����"ӵ*�� ?�D�(d�@�)6L����-�:��Q4	�tb6˰YA�Vj+D+o�2BU��2��,[i��6�V�1\l�|��@%_�$��*�&;$��h�p;%���YB���4�G��l�e �t�jRZZrT�a�-�Y�l/ŠӬ;Xk�Ār	fbR�n�+�sx�Ҹ��ϗ�B@�'����� $���{�������B@�'��O���iћj��l�YȴN��2zU�jX�����3���	�r�иN�V|o.�^Ci�s�w�1���o����%�Ⱥ˒��Htõ��p�t����r����`Վ9:��	{���Ii���b*��8��:�-ó����C{�ژ$�+�l��#s\=O/3D�`lu�P��K5��R��6����j�e��<���h�]����.;Ƴf���uu�@��q�iMAJ�Je:��)l��μD��UZ�o�
K2��X;�W�8§YW<K�d@y{7��d��U��2�!�gY�hq��w�� �'�uv�`��M�ŝ�����q��ւ�t�,E�;��ԑ�Gtrdf��\�0'�ou%��(�nά�QnͲ{��/��sMh��x���&����콫R����p�Cc�SRX�����ˆQD�)��<94�CF�k��ˬyb�i��^�4��uܸ=�.����	Rh�L-�3y�S�P���Uk�Mjۤ��K
�S�n^����L��Vα���;*���^f;���˶Φ�J�4g�R�ı�a�RK����@�+���f3�0uF��v5�0嵵��8��;���{��2���z�i9QVsM�s�v�6�i.���A7��D�]1���B�J�P��i)D@F4��E�3t]����/�i�m1�`aB� � �DA ���(AA1 � � ��(AAP���h��T34K�r�5��>��l�N4ˈ��V.Vg[]	���m�r���hs;���6�Wܖ�9�f���ٹ#���g!J�	��Y�Ypeݹ�Ǉ�s�w�e4.�����ӝiU�C�7k���TSa�#)��Sx�toM O:eN+'#ף9��,e�5�ie<ljg��9�YV���{�̽.s$;ꎣ�3z������n%x��.�*�\����ᕫB��������{ �1�#��6�܍����>��+:�J޶;6i�U8J�$I��JR��1C�nU-��`��:\�Z��iÚ$���gvǺò(gk�w�K����U$��s��f���rVts�B�a3nW!ѷ[�ŋ��{x"]De�ܺ�u��J.��/`�;��J����=���C�m�U���.V�ʔ:m��Xَ�Rw�N[�ȯ��N��u�����U��أ�d��[;����)��B�����v,4�6�\��ܜ�Ǳo`�c)�z��I�{sm w
�S�u���H)q����ݴ&H�Bh��p:��{L�`����Ng^�u�ѼJQk��ot���B�e}�&%���(�f<�~�n����%��9{z��-jQ��Ԛٗ1-�����	�v�X9�ڼ�c)���\.���[���3c0���~�T�n� �A1 � �A�  � �� ��AAA � ���G6!�9�s��fw=�g��S8�ԫ�u�"n]���x��1����x�b�l��w ������-�{D�%]k�V!�Z�Ƚ�i��Ρ�Q�w0dV�{#�H)η�a�5[�.��g(�bW+U4�����:�ö���m*
��H�y.�Z��c�B�������f�@���*�#b(]X��m�C��X�n����q�l�w���rh텶n�Yt�v�Θ�4�Sf���r�1Y��_:���V�m�ŵ��μ�x��lۻ�0kt�FJ�b�bW�U@�b�驳l@.��7�h_P˂���"��]]��@hS���
d�Y�-ˮDixFgq����D#y���[c�V��V����l�k]*:8l�X��96�3r���������j�vs�{s�59�wT��X��ֱZ4f'W�պaΖ:��c��On�eɈ�Zβ���o�c��!U��Z����tU��b��j��^$�Z��]l
F(�RU�3̅^j�+�}i�.��U��$W&'
�|5�G$��j��q��i�)�ɵ��`܍�G� �.�oJ�^���.� )M���|NU�.:�_;6�.a����[u��(�v�ˠ	U��&��	ݘH}0���i�z]�"Y�HN�:j�һ7�!`���b bA@D@A!Ab �8A � � ��AA�E"��5�gX��\N{u��&�w��ҽ�L�O�#��V�{f��V)��[)�Nޅa��!8�Α�5C4]t�ol�:��,�L��E��.ʒ�J��k��u�`�U;%�[!��A9�c-k�f,�-L���3s�Q���:��&N���\yݼ��k7�qXĚ�y��P�Q䂮*M�ͪ8h@վ��S�N�^Ģ��D�V`i���\Y���ᕷ�f��,ꡚ.�P}�$jM�k��)���u�L��VG�a�]���;�&d
�
wi�����@�v�C�ʞ�
RAN�ʕ��+2���M�3nƞ�YF���w�ˎ	L9b�Ի�H�#Y�l�2�{ʵ��E`��K�F�����ţVlvY��Ț�B�;����+"'+������$��G1]�{OB��}�4U�c$��:f�xT4Z�?��j�Z�h���^�
bJ��T�_����q��T�n=s�[����{U,P���喃�Q<�ʻ]��J�;�q!]�(N�ZﺝJzveb�W�F	��1QR�n�"
{��L�.������zoe"%�\* �9��|�[�73:�*���AuB��� \�^)��ar��V4G ���,��^��YE_z��_eg%	��]�|�R.17un�m)Ϯ۵tL�ܥ�mS�jJ޵e��ͼ��C0�A � ���A�,AA� �AAAAAAY|�SΣom�r�#�'<#�ܫF��N��: ����:��:�6�^�B7�uV,2Mッl��4�Ƣ�j���|�Q�8��d��2+���;�(Ԗۀ�&Y���Awu��W�}�2�󧋙�}):r(Wt˔��tl�f�Ҳ�ji��msyz��w�.L��9������5���r���I#T���}�r����8:Έ�Zc���}}�c!�e�ݝ:[vds@@T�{z}�� �y�R�d�[|�YR��YE�m�*<�F�d޲.K[�.�чY�{׋ric�˱$��M��թB���rh����+z7T[�4�=x�f
q���L��>��;���(>��%�Yu�뻲X7TI�.ӫ(��O���+0�,]��f5��U���|���}b��juy>\i�@��MUvF�^a�*ؙua��˽����@w}�4�ٲ�����:�u�I \�t ?T�W\hj��,T��C֩r�z�6��V,��iܓ�]VF�����nw�1�w���X%�K�n�vxs���&T�%e
sc!4z���w�7�-�K�K�0���:�;4N3XRs�|Ļ�Zu�팜ݻ��b�I�ղ��uA�t�1_D�@���lpWie9/U��ը��ީ�gcePvOu�� c��� � � ��AAb�AA� �A � �Ab �^�Xs�k���ku\��H�QLRQ��s��=8�^u}-cH=��8^P2v�U�:+;��H�o0�*˕��-7�,�3 Of[���;��f�,͓֯ڜ�	[�y�m�e�}&8��4-%P%p_0�k���5O8��Vi�4�"�"�L6mL-r|���0�"tD�ۆ��-g�e;5��[ee��?S_*;ք�s��/�DPً�i�h�o�͗ߕ��O.�E0c�8�!�.�r���+Ձ�R�Wfޙ��r��;��V�zw�z�:��F���;3�ҭE�5�Iucm��:ٍ���d9i����t�S*�l{�7x����Njx�P�/�>ѹ�4�[*�lY��g����"���YY�=֜��O^"ފTP�����{u-)ϻ����%��Ic��%�9A;�P"�����q�s�-����7�pe�h��+��l�v�h�Vox�n��RG� ��1�v�伭�W���MoH��e��Iջ�^�݌ҷ@X��wr� ��0P
N�*�#�Gf�pF���u��	1'���R�o~��a����*�1c ��X�k�ۘha[gN��m�(-eT��R��NBNYN1�A���j�K�}-��1�ؤ�{����^K��x�O�UP*19��F�4�G1:9�MN�������-�" �:6t�E����X���X��0AA� " � BD(AA �AA� �Ah� v�}�Z�x���\Le���`yZ�B���^�bn��@���I�0�B1-���[g�.$�8���IG���X�jn�yAs��՝�ӹ���N"5v����:Bó�lڱb�v]ŕY���r����֩����<�t�����yFJEf�.�v��M�|oEU�����]|>��޴P����l[���)%��X���
�g7�v�u�9M�v�W�:
	nB��Vs��sq�vֱ�cy���R~ 3}����]o��<�d]��u�:,���;���ޚ���2�Ae�6�m%�C5m��m���T}ͦ���K�QjZ�����t:�S�ɚ�]�+P�M
���CT| V1���;��n�(�[�1�)�HT�&�l��.�Ē��;w��E��03�(2��wn���vⱹ���E�w2c#�U�1�=|�B ����*�eE���d�״��4�ñ���P=fer�����	�Yv4�ͱ{y�#���w�-���	���T[�lMk	b���[V���A��X7��}��ݸ�p�&F�<cCG}��"p�8���s85�Y��qЦT�P~��^�"�܎����ٵk.:��H����8榅t 
v��Ne�,w&]*Я;�2�}9�P1T:�&>'��;�8.�sI�J0O���^[��qB_L��v�㺺��4 � �0AX� �AB,D � � " � �X� � Cj��=u{��8��:[�q�ѺX�NΫ�;b���1�2
y5&%�"g�j�{0�KÄ��î1e?z�{O:�Deh�;6<�v]�+R)�;!�y����Y<�܂���ayv�\V�
[v0��_YQ���4x���mӟU�����TMU�|M�=�о�w�t����M�Շs�a��t�Rvp�:_X+�5�	qKwMj��f�!j��$�Q�΄Ժ+�Hx�>��1�֫/�b�]j����[	�T�r��k���g[f�e��_c�7qǠM�8*�ćG��I9^�hU{G�>]�X�`h;8	;I��+M�D@ ݖ*�����^鳱�e�%�:KVx�
���ݘ��JS��Op o yd����0��O�'[&峀��� �t�vR�C��V79y��=��
{9�fͼ����3{�:���5�M��%�B��_'���N(1ȵ� D*%Y����X�ʲ�E�݇'(�ՠ3���ޱH��y�޴(w#��2���A]+of�aJᛃc���q��IYy|���1���}�+��q��t�n��[�<�����5�s�����۽�9ά6	{)����gf҈&p�wWol�@'-��x��.o_�y�.��y����^f<ݛ؂yw��.���E6��eg{{��5�z�Nx�R�Җ�R��8P�ز����7|���,��zs#��8TxRg���o2`�n�m��R�.�N�*��Ea��Ab �Ah��ł AAAAAAAA�ߝ#5����*�ۯ]�P�gI|�[�Y�d�y.̷K�+�N�V�]]�V�A�b��B���X6�XgK��eltL���*3V�W���yo�ۉM�[�CpK����#.�3���i{�]��Ζ��Ր�Z��`$���b�� �%��:��4�:P�u0n�����<u6l���FB��tJ!̥���(��3��u�zVin�+M�S�0p��j�q`�"��r��Z��8�{uV��Pg��gl�T��J8>�ZG$,�I&�nv�˵Y1-��'UV�o�&�WLFU�[�9�޷e^�����e�]�_5��Y�璨�װ9�R��Ե�lOK/�b�W���l%��{H�T��;�Sy��C&c��VV)���ja-�դ���מ��'<WR�yb�w[H7Fd�M��$hq�}�!B�B�CY;Q�mY�[��{�M��E�[vb��Քl7�p�ȍ2��Q��'A����k���"�:F�+x)u]2-P��I�*��S�v1�v5��U6���s����`J���1�WȻ�Et�8Q7+���T���I��r���lP���	�l�QŌ�����bg�A��olL��1R�"��WWt���q��M�����J�]����']�$���ҳ��7ԍ����։��VG�_�車<d�����gΨuwf�����s0..�5Z��>7\y4�m7�n>�n�>[5ڄG6�w��]T#��"��+=�j�R>���b���X�ٰ�
�@� �p�|c~j�on]���pk��Ǡ�°T�m�:����u!��-.ͥ���9��v��}-|����&��U��R6T�I{y�ع��n�� ���$dk�j�����A�Zì������TH���9��fQ��)�Hk�Y�uV�~7���#�PZ�����s �J�j��C�h�V?�-�+���v�T�"+feщu��|Ө53;sr�� խ#�U�s|)=jo�x=�.�5}ua��u�:�OZ����9���-˖ �]������2N����L]C�9���xs��ڠ�S#��˥3f唵��V�N$���<{�U���s����Ƚ�{3"��[�1.��x3�<�T��u��m����f��ѭ*,ɂ1�r�R{e򬕼��\�����ĥ����#��ۜA��1ʷ$X�.ٔ*�A�G{�4N�Y��g^:b�˺۳��4�m^��N
ل�����X����z�b�G;Gq�s7r�]����Z<\�Ր��������d��y$�Ԯ�h����Wg׮*�)����|�^�+k/�A5�w)���h��^���\�j5k���$Y'n~콜ܨ�G>���0v6���݇���o�)��9]60Nbe��0R�#�����S:��!}	#-���4����a����2\#o���7�	��R�gcL�cvT�L�v��m�[ǩ�J1\R+�Ӎh��:�G�O��"u�i,2�GNqڭPSor�;�C�(�P4f�������R�����]w2�Z��d����;%J;Ӎ�#N	�7�5ڶ��wmV3�-��/��M�j�9I�m�O��J������q��(e��Jz���
��\�X��c;������+8�(j�,ɠ�b��}UG5�0wjY˚;�{9������̬�Q���G|��+ttT�}�&�z�Z"Q�3�Nvvl��yac�#0�4]��jvF;K[+qw�����P�f���|-�E�Q��N��ͭiѫ%��Q��v�i��iǙ��p���Ֆ]VMgT7]Qw+�o���Ֆ�+�Td�A+g)r�v�e+i��^cwc�cp��������y��Ht׻'+j����5U��s��
����Y�N��� ��Q��� m��ir0݌�!AҾ�@�՛Fa�o�f��O�Fdтe;�nP�*Ȧp[l�7��7zmTzlt&������t���Z{a&z��As�:�G8lnN�ؙ&ۻ{6;�RB(���+N-�MeǏ1�U��m��������rF�EHm	��QwI�d������H�b7�P("A?��u�B#C1��*ym+�c2ؖՔZ��L�)ƣV�*%��QK��­���Ӈ���R����m*�l<q-0Ķ���(����-��iJ��6����p���Ç�NZ�,J+QcZ��TJ�p�-Z�Lƃe�6�*3)�B�am�(�yr�zzxp��
0C۱Ļ�Gr��o����QU���(qșKXڱ]�a�[j�[�Sf��8x<J�b����2Z+h��K�f؃0���6��m9�b"�+J�U��b�_iW���OON�zz{i��S��VR�{��fA�I���3y�H�^:���\~77.\p ��&V�I�)��[�\�(�WN:p���C�mq��>=y;̗�*�	�/����� �4DF��f�c������߄�8�mHX�Zە�%��-)Z-���O��Ӈ����WV�!2�F��t�͎�8�IVĲ��Ƥ-�M�0�n@[�q�e��IupY�Ѵ���Ǝ��P+�������ޑ�[�}w��=�ʭ��)��W��R�J���Ͳ�l)��͵�f	r�93�ĵ�r�h��n�m���"�0�AF�P�!����12�Y��]Murݼr�o!T6"�+�0��-L�mne�Pr�ʑ�R���-�0�����7�;�;��'JN�!�c��L�ek3�Wg^���iB�Y�Y������FҨ;���m�.L�6�W
�����,��2�7{�6IZy?�GS��}�	;.8�O�����ͽ�FfL��C3)u�v��j''幃V}[7Q�,�ܕ,��JW�B���8��dR�9=�䮝�c�A.ù����`���WJ�3=�g*U�\�j��ќ�J���W�,ǓKͯ}c\���������yY��_]�̝�[|��@��=�P����bF�`���������B,�۪������7ѯ	��y�~�
y�L�`�-��X������2�J�篪�����̒xt�=�w�<�'��8_�E]���L^�N��Kޒvhk�rz�Qh�����}��^��5��>����޿{�R"G�
h-X.��{}���1=&�睉�������{���o���Y�[c�eS�!/�p�[נt�{&�N���R/j�gc��5#A50(�MXբ��M3wj�GeN����{�W��n�b�6�#3f��u�_\���m��5�b2����[�0U�L��'e	�vo����k���\�V��ӥ�TG4�3�ӂ哄�}�E�n�;k�����YC>����LJ,zY��E�+�w��yU��j���r�/l/���]^X��N�_�exr�|��u:�x�e�8������>-I=Xl/���UI�1ʂ�q�@q>4w@���e��U̕�٭��ͯt���f��oyZ\��q����Aw���fόaJ�l���I^긑������V*�U��Z���7�Y}Iw���އ}����|}׋<����˦3��JĎ7x/ZZ{�Ă��Yt�����<��o�/��F�'�N�}�AV�3>ޣ��{`�����yO��u��^ܲ����5,��\����OQʫ�>bW�!�����s��������oH'�ŧ�G�T�~�dq#~��<c�}=���������;A�����fp�>�߂��5�ة{�%�y��z{�����x$�Ԇ�zŗ�e�XA<��2�ìsi�od��sQZ2�����cj�b�mV�Z�n뎐�pW��<� 0�xì�˒�5��J�i\���;�]�n�'6-����[�+��kй��Y�o3�?���b���ګ<'u��]&Ȝ�����
~�*��J��f���Z��z��fS����a�K?�]lN=꿵{�S�$<{�^x6����|�p	�ɻMJ��-ж������}�.���'uz(��N��p/����~�J���Z��kx�ǭ��Z�o�����K�3�Y�au��o��\��V;u��¹��ݞ�ƨ�'-��kC��q؏����A�9��mݟ�f$u{o���iGOl�X<����Ϝ��9n`cb�Nx�A����d���o�&��g��{�sl8׋��r���63�jv7x�0֜б�k��\<4Y��<snw}A}ݬ�q������a��aW��^Bj���M��.l�*������h�N���C/���O���w+�ԝ��U���ݵ-�¢����݄＾��%���MkKN���!����Pr��c��[�o�&
�{��ۣ��0����� �5�e9��;�%��3�L�B|�/��&:g�ɥ�rs6���z.��3�ku�̳|/y�.�����W6�LB������UN��N�<�o�eT��Xsf�ޘ5�ZП���<D�y�i���_7G�;W�-Y���z�M�I�߾�b:��R+�pW}ԕ�u+
�R��۳��z���Ú:�=�o�����r�hx{#D�vЍI_K�R�r���ۖV^��3zj5��OŴ���k�v�-��Z�as-߽=Om<��$X�gh]u]�b��ﺽ�&.c����.�|<6>�%V�3��r��z�)�J�1�Z�d��3���w�Ͻ�ǃ�t�P� �x.���{2l~�ˮC��K����G�~�v�^�I��#cƈ}]b�+��Lzmy?Uت��"϶�����>���u�@�n�=�o��ߔ�����*v('�(�n��C�q	��{�^Hp��/U�=��C9���zw�Mڿ22-<���(k`Ė��zi����Cp�ܻ������<���G��p}瘦2��F�>t{(ЇηY����^�lw��7��B9��nL@�`� �7Ν1[P�&-��R��&���y{��վ��8L�}6�#1�u�S���o6�J�wk��H��YWtZ�����۵K��zu<��nF��S�*4�.�w�ۼ0��~���LJ��xR׶$�bHUX��;�&M�`j�y�$=~�x���j�5�U!yJ�����ᝀХ��]a F��O��*f�A�o���@mh�_�ܟX�O�b]0c��]��X���q��yN�v�I�Ë�-E��!�Z�/)V͕_mD1S�
F/|�Ow�b�ո�I:�eܾ�ݗ����?O]OW��`ͺ���F��&շ�3}�՞�TF!}`��e�*�x8=�$c�����ȷ�e�m����K<�\>�X{r�`�½�+��ޙNM���zz׍K���G�>%���F2fxr�g2�^��y-_���F�p�����WQ<�n�]��KFD�.�ާ�{>^���6ev�kCdX�X>o>���~�c���5�2�>��J�ϥ����X��LKd�Ou<��-ɓ!TDQ�0����[�U�3{6!#p��>_Kh�L���#/�]\]F�횲׾[��ѳ�S��M�Y�`���tOIU��j�J�!��q���exگ	Ҡ���Q�O�\�r�8��+�8�v:C��VF7�.�;�n���f��1Q������7��t����jW���oӼ�fy�=&y��kb�b��x��2�#U=���7xzȓ.�Ϟz`E�z\��{��ޏ'L�n��yrGydTI�E�j��Pޑ��|�g �o�K�$~z��{�y�;w�.�)^Z��e�'q�{v����0��N�^C,������x�Y�2�f�:x����l������碣)�\�ڋ�]�G	���FV��޾���x�8߳ި�˸�Lz*3X<'����s`�;�G׈ӗ;z��zl�$�3g����V8�o�A�)P_����a/1�Y�/6u��Y�U�\��uؐ�߀���rK�9���]U��i�}�҇cf�cY�k�j],��1���������-�]�0��������݌��,�h�����['zz����ni��Ю�P�v�_���jۂw��:��05�̌t�xe+��^)���L���N
7�F��s,��	��=���ϔ�o
ꓒKn��[�-x�F�x�j��n�$�ݶ$[�:��順����V�=3�v���U<�vc�������k�hC[�.t�+8%Vڨ:J���Y�����>Ϸ�G��!}fA//����IL��o��K:�zu�������+�n^�g�{F��;�Q$QW���
����LxO������q��.��"�r���hR��_&��V{�����叟�w�w����;��7�y=�=<�<��'L�b���~���J���{�%�h�
5F��)��}p+�{D^6'y�?o�%w���ƐzOv���??]a^�^�.�V����+)�j�݋�����M��Uޜ��*`���}�W�Მ�#l���F�C�Ѽ��?l^�[���׋�m�w���۞I�~be�{@;�ѫ��F{�1�:?VP"S^�y���,����+�)yz+L\y�[���
�'� u��S�s3ģB\=�yG���Xj��H��=N��E�[��̚(�i��K��|,��X�u�=�n�v���u���RuV��u*ξ�${u=��ü� ᱻ�9�I.=w��ַ]^��ܝa��>�Kb�ަ1�q[��u�v��TC�[nv��:�H�u�Vsfa����Qg^�	:��7���̯��|�+Z7|m���1*���I�c�.HlD6wm/X�}��I�Ӄ=��R�n{� �a";���3��	�y��7���s��GL%�^�@9%X3��X=Q�a�.�X��z�X�{���s�o���Ԧ�8o!�`�	"�Y��R�yZ�L������cݞu��y==�+5�/N�Aw�ΐ�RW�w��m����c>Af�.ze�'�a�'���r9�����
2*�8y��	�)s�=�<����oTV����ukӧ��X�/���-uAa����I_��0b�H(�;�O����mj���C0x��uO
�ݔ��i��Ig�W+�F�[U��%�e(��%ħ��ݯ|}�v�\Du�`��p;����/n{�i�����*ٸ�{�]n���=~p���>�����07�]�`�c����}�+U�=R�\��;�HK�]��Xvu�'�5�b4;s��5��D�V�o��a��8���j��N=B�6t��&�4�,���Lʃ�[���jl�F�ד�.X�X{�"C`��r�8m������EMB�]2�g����lЫH-����SL���!@�v��}��Ӭ�
��B�X����s�A��E����g�@Y?��̱2��`tʩ��5ygujYk;޸�d��Xo�y��ڶu����|�oO�7������߬nw�)�[��"�z!~{=&�4"��觡�
��E�?����S�>����ԩ�>�r�!7���]^��x�Z�Z��mǯ#j�9_g�ԾM�+L��J�tX�<h��`��� ��
bj=��w����"�Y��jZ��D(t_�}W���zy>�i�v�7�+�ˣ�N�/�hyI�ţ�����]�l���j�|�a��~]V����{�3=�ޡ#��G���U�elŌ3�;>庻_����$T陿t{G��L�Wd�[�[y�*Yh@�a.њ�V�u*O�Pu����������g��?zA*Fv$|wѰ4p^��*b�j����=�jͫahS�=D^�����b&=��ǔ��2���^"-�Jv{��]�J��Z�Nx�;�6��1{1���׻E�8na1���R��O�GH)@�E�k�M�
\w���q2o3��>�u�ΔމΚ����5���B��nt��4�hEl�m��$������"��8��^�#����;���Ǆ������|=�����C��� �ɰ?#���{ú�X�뙟o�D׼;-�[��;��4��K��~򷝍w�����mP�ʾ��"����8d�B[����*r����^���r�yHm�Ok�z{����&^I�>�)��ᣁ�U�����{���വ5[���3���7���� �p].Un1YH��g�w<�~D���5X
�5�o��H�d�w�-n��Kv�Y���n�����Vޥ�P*��
e�a���<3(�����^>��t�����p�G+Ooz���MOD�Xj��m+�;�}�`�� �)z�/mX��b�
Y�+Qn��.��j�h9���bt�R�J�=,]6ǖ����or���[{�!FF?�<ݳ=��.�
����!����>���ۙ=+�}U�U��/����=��>�p����{xbn����|���[��d^��׸��Lu��`������Kq��]��9)��w9cE���\�yI�7W�}F���Y 8�
HN�W9�A��>��"B�&�<ŵи�;+2�5D���_.�˂����`�b��n�8��v�N_!fet�Cy��}%ڀe�Cۙ��ڧۍ�ͷ΋�<��/+�j���k�y�
�4�Y3�+zlyW-83c�j���/� �5Z��a��Ĵ�v�z��6b��6X��7�͜{9��yw4��<Z�F�Q2�:$�n�q��ahv	ٜ�Q��e�17���yFg�N��w+�^EOkqJ�\2�Bb�VT97B2 ��W=���HW�u+/�f��P!q��:�tl`�;t񳵮f� �#Ap5��x�Ɠ1�y��2��M���mW]���$��4Z'��/	��c�����h�)�oH3 �,�r�n˘�{~�i�l9�J�kJ�5�V빌i�V�6�ʚ�;�ޭ'�e-�ndѳ�KD��c�#�����^j��o��n���Ry]�]�lt�ȓ,ś�pm�9}s�Y�f��2�dӃ�tg5d]Gb랿b��h�c��ʇD��ٌ��}����\�j=y��L5�V{���-�fQS
묛���F�gfZM�rU��Ez���2�a��uC��^F�O��'|��d�����~7�-K|�p:hU� =q!}-�Z6<�zq�����j 6���7(������P`��8����p�sw�W���r�);�OY� A9��q��í��\O���]H)��sC�ľs��{�Y,W-sXuM�Sz�f7�&õ/ea�R�Q%��ǉ3`B�w&���L6�Χۼ�)����ĕi��� Y�}sz�ͤ��gcEcfK���j�Ρ!
���3_etYQ�Ol�����_��f��k�O/Li��;����t�QCV���*��w�L�ҝ�5�J���ۈ�T��.׭	�b�\N�o^P1VN�Vcߓ��1��ů���c�x�"�,s��gT�t]eo7S���L�$Z4�9}�驔ے�Ej*�2<��-�o)�c�u��R�%�Lh�����=W���½N���JWA+w�p��3\�8��ޱ'{�vY�2Ĺ0�cvu�7��R�>7�,>����c �E^U��96	�ݦ�o����� �ucݳY]Z�p���l̰݀��٭
;�����:t�%Q���ޭ��������+�5�T�Z2q�a:�&� ˱��sT�Y<
`�C���ku�(�
Ť�ǃ�[�hv�P�3��d�=!���X�]�-�VҺ~���n�f=�du\6u�\6N�uz
6��`ݒ�Mg+�ms��i�1u�lnE19�2[�k"���9�_��v�現�<9ecJ֪�^8pyp�Z�3v�!n��wn�d�MJ�)뼦��\�Q�QG��x@1cF
<#�"�	(�p��ȵm�3w��5��q�&[1
��7(UX��o��B�C�*��)Æ8p�G�U�V�6�Sm�s3��76�V%AV�UN4Q��7lKw
��0v�C8xp���r�dDS#m
��1[�G��
������0�[mA�k+-���[�����xx5��a��Ɵ\]����J�EȢ#Uxܢ"��K�(�N9�5�300L*�[�k�xt�����q��y��Kj���c�ki��ŧ-��/mwsGQeD�+-�[lV�mRܳr�L<<<<<UA�`�0Ƴ)��֪9n��VfS��f�12Ѷj�Abknڗ����=�ɏ�r��V%���2m��K����UJ��ȵLƩ��!�Yk����mjQ����N��LN�ǹq����Q�s�q�Dʢ2�k�m���B�[)�ֹ�n�C.i��Q��.b����j�7pݮۭ�l̸�fҦ%jD���6�iL��d�nf8�,̱f[[rҷ6��N7��3�5���Ԝ�F���b<�q^;vygX�u�;^-��ʇ�;�'Jq����a�
$��t�χ�C��A�9�����~F�a^o>�T���?wJDD_ÔHB�J�h����r�J޶�>z�b�[���u����?�~9�GF.�~f�K��e�'��/����Xa�RG�s՜����<���T�y����_&~�
��af��?�����ȥ���#��rN�>�ʘ�c��YD(�JG����0�;�����*�/M?��W?u�'�B�~�~���^�_���ٿ���C��s�ϫɚ���[����`����ٽ+�c��
�x��xc�U������
��`S�մ��## \Uo��{������`���H�����&�뇔ո��L��~�,՜&�#��?D��X��tߎ�E��n�r�l�D����=4�e,��}B��M[��{+�>�Q%����Z��7\wNg{]x?�0�0s�#��
��`]�RE�V��
f܉O�GPP<m���J|����C�`Kk�&Y.z�b���x��؉�	C�� ��k�|
�8��[��3��X#���^g���4>ل_�3���z럻���25㫀 ��ND3��|'�Eɘ|o�U�Ŵtf-_}�T��&��`yT͑��j�����T!�fˮ3�휡��Mq����ȕ����MH��u�<쎭	}tBu�k�ߖ�ʞ���/�+є���F��9�W��)��ot�\m�x`�| �Nt�n:����[|�v���䖚u_���*:�ޭ����a'����33�G#$��i�ȟb��r���M_P��	��ϫҵWD�1�|w'����|w�������7��}`B7U�t(����-�:�Ov����z�C|��f߹�$��g_y��ҁ֌�d���[#���X��ul�����w�#ܓɼ�5�H�
���Kf��T9;wc��}��k�c��5����g��׍|�������/_����}^��6�D��a���mH�|���?v�X�������R��ث�*�tea��ƸB �a�3�E��@@�|b�oߏ����|���=���F3��'�F�����Qq�~��3?Xo�r�-?W킒x<� O��$����2��v�,j>�jk��:�q����=���)�,7��&�������y�=�n���xSf>�DW��Wy�:�����H\��u}5՛jPgcȰ���EC���S�}���+��Ñ���G�\�(�����v�X��)�S^?E���F	�h��*��Ҵ�L��X������Ѹ��9%��V��~u��~۫��wq����Ҹ�/���Jc��Ձ!j�-���,��ʿ]��w�����f��'�%4yϯ��U�M��Wu�h+��{���4!ֺ�pl��EU�gE���g7Jd�B8�_���K��7��C�ʆ���)����8KM6Sb��~#���y��Oic����>�_At#���G��(�.<�i���-�v�ڈ>���a8z��q�aL޻�8Yj�#���ya��?�B>�q ��s�b��ۇ����'�=Cz*:�?;�O|-.��,f�a��Q�l�a���EIA����@��0��W1��_�f(�/wMU�y.����6~��mz9����46�W��#�'���?0C�a�>��3�tR�b��)v����`yZ�oӡ���e8+>N����L�7	�A�j��¦�*���Q��3��&����c#��O����,�M- f|������9gb� ����Z�F$����?�s��rǣ�R6=[�`c�4���z�	�G"Y���_�Z�M1���[�v��u᯴%Q8/��8!Ǌ>^�#'월�N�A �:9I@�{tJl��9��1�۞�d]�0DLhu?��{��4����B��
@:�,��υLC����Dm{�j�j�ΧxA��r�ff^��%}�~f�C�|��(|�NB�|FAJQ&>bA��1���(����r���/Vn���ϰw3�mt���+? F��'¸!X���v}��&�
7�a�9�\Tn0�VD\�+��y�%.�Y��f�����4����Uk�YZՋ#V�
��j���
�O0+�[�XŰ���,��K���Ms���F2#`#HOϏ˥�y��. �eϼit���܆!��Q�/`VkI��i��>��|�sx;5�d�o�Ͼȥ�Y����7� Vō���ם(XS�7�[�Ed���/�rK�Pz���lMҽ�������j����#�n�?;�\�XOnUCf�ރ�8<�+�!��X��|5���������˗�}�����^���0G��yϣ��jc�<�8��8w��ųk�%�w��b�vy�vDG�X�y�>��L�������a����Tc��������
T�s���W��W�%�,o�x���J��Zvd���zw�Y�����@ȶ[��HB��D����.��KQ#{�_y�3"��k�f���������x#5���vj�`��g2��O�<���#�O.>�p�4,�oՏvL�7��C��lP�ղtw��p0s�h��7�޹����*,�#L�q��O�ȽP� �|"}[o�������}`\����b�-���v���)�z?(H���l�&�s�&� �IX��q�i��LV>�pd��5���N��-��Zv���=��T�UGq&��F�<�+W�4��K�,�����Ɲ�)�l9[7���o��,o�Y�x�����i�v����-�ۥ��eBo�S�ƀ��vh���m�r�{yN��k�)�Kn���{�\�����N;��gl-�.�Z�E�jY��3w
�Ⱥ�2�^���
���C�A�H"H�0Hz�-Ę�,\h�d�+�D�;�b*AZzѨ�uڌ��WDB΁�Z����M�ݾ,m�Vߴkop���t�����L ��t8s1���~h�q_I��5���!���}6��2\\��u^���wvA�x09_������_.�'�<�zs���@�� ��~�%�7��*������^o�{ȍ��P�������~�yA��o�Z&���`�	0��&C�
^p{״��5mrյ�xC�溼�}G<S�#�v� �wJ@�	}�b�G�����2*�\"�ſw�SP`<�Ep�q�	9	����/�ct�DN�R��-���R���LfVm]P\�/��������W�����<�+E���e�;����'0`�NB�n�����<<)���h}0_G�϶������X�����^�8g��\'F��2��Cy�l��wǛ������zb�/F�*BXƫ�g>v��-t����o�#��Xf�b��d6mg�h4��T�͇>���I�,p�����!9MCgj��r�8���E���M��i1��p`��c?!�4!t>Sy!H��U'}����"f+�4�!ұeouͮ0�;���f���'�J���ź�bAS|�l%N�Qɉ4�L\n�gpq2]ğr9�J�Q�J�wG��ǃ$t�d�]�a��j�e1��x�#+M�U����6��萈�DHD@���#�>"> l$��-{���"�}R�����
�w�q��0˰��M2�T.:�jރ����~>���pߣώS���c�$\W���\.�hǡ߶���"����3l�:E.o�tg���P��ӭ��\y�'?'<��/��s����Ʌ���F��<#ho���ς�SR���69N3���Ѐf纣�tf� �D\��4��p�_}}>gc� t
�0�������>����^GE�A^9�~�kڷ�e�P�96��;���G#$Ŏ�G�$���6T�5'�g���Z^�s&���(��:�W�w�7��G�s�ȷ�pʌ�U��X-�Ү�z��b6�`A ?��y���؇��A'�as7w;)D���1:-�n�4e@���k���n�}A�`�c�g�����;M���X����p_�'a��$���aV��{i�eU��A���׆��E�qt��e:��*K�ۨ_ρ!��`��. ��������ly���@��)M#�h��"�ɼ��W��Q೯X�-̐)~-��0�$�@�h	���|~������s/��S�s���v�G�_lW�����i���<�B�y7�Ny[��?-����r��g��$f��Ү��Y�*MӺv�xc��L��g����R��< �i�s{��(#��gT%3t��b-gC�x�v���pGK����9���՚� @|�۵�7�N�?�� " ���H�"$���a'��y�o����}4�L~�y#9*���`��F���_��E��>a[��6*�}}T�*���[�2�{�Q����N� ^t�
-��"�U�o�62��'���`a���3����e���]5������=�:ە鼋�,3���Xf�VW���k����V���\��+Q1?z�[��[7k���<ȲA��S&�L`�轅;-���B�F�i�-������+��,�X�����w�R!��xS��������7"<'d��G�S4����1��%�G�ѻY3��g�C�~�@�*/��hy遊�`�X�ܓ#rG@��8wc��0�R�k��w=�k�nn|���B�;B���r���U�ّ>�P��>�3�8Qq�����!'Nw6��w��yva�9���u�o9VCE��R:)�k�+G2Q\� ���U��r�~�2����!��3�{滽�rd���?��=��h�{.�~���W.���B���"|�)��,Q�V��,�b�k&7��!dc�
�k���c4��ĝ��8]��w�+�r����ϖ�Z���1�����\�f�%g
|X�|�6+R�t�g��_R�L��l� �~{P�����bq ��t�i^P�2wV��뱩1���tí�#�b�WW)��2(N�٫5a��q��v5�uf�E^͸f^�N���˿>f}���� }J2�$D	�>?~�_ϟ����٠�*�ҡد��o�z��;=O�>M�x}�����&_{�!Y�����x=�0�'h6�,H��O�1ң�wJ��b%���b�����@R�њx:f,w8���HwD[1I�]GE��~������$�y��G��omt���/�ͨ�sS����=��j]���p/L��s�B��fc�h��T�P�<`�O���*���$_�H��-����q���������YB��>Z��'=8�X��6܆!�<(��>�jk��dD��T k5�
>�N.���ݘ�r�����7��zRb�W�m��JU�Y�6��~��jȼܫK3+v���ݕ�x֊2d\1,h��#��s&��9����3���h��Ч���n֐nE��T�x�ݨ�O�𺛓�spx�	?�~�'��xLC}�m�tX<�8�|����K�4}��Ǽ��y{�B���6�����o�o�9��"�dR>��Cb��_�E󮎨��]v��%��˯r�]&�?E�3\^�R���Y���q�`���g�dK-��!a����f��}p��r��95r�
�f1_r�����������һ{X� �0��gn�-Wr��v����|0��ц�Q�r7י\xA�����-�ڳ2�lp6��=�u�ݗ�eե-��c��l踻�v}���A�;w1����� �� �# #'�  G� w`�+SLML1����!mݼ/��Ce��75N��,ʖo`L<�Ş���|˨O��;{��@�E��(�w�ɦ����Υ�ƚ���1��*ʋ��|�y��������������诧��wRuw��X�ܑkκ�b�X�G�N}
�R�Ю���*�Ki�iԹj��t���~���'c��e�](��������Z�Q��:�.���.�.w37�^�{�<R��1�_�`��L&=�C���?��A}Ú�9���,?`�դw_���|����9�z�_X픎Q�s��eDm��!d:?x>�_I�O뤫��-e�����r�<ǫm�����j���骿w�����y�(�dW0gD�hg����5��fX�G_���W���IFkޡ��}Mϑ�����7�-p���T:h�.&Wc+�>���>��c�P��H��:�#�t�*7^�cúR�D�Ю�Q���kſ�p���}����5�p���8xlFIȀ�أxm`��ء���P;F7�;�ZK1���fd܋���l\x���sŭ� ��KJ��)M��J�ow���뒛Lx����(��ή����%�'ހ��U*�U�ky��1��f(s�u��\���dY&g�%�%��q�e���k)�]R��o����>w�\73T���>���
AH��F#		����{a�[|�1�H?��Y��l�lL`B�*+��b�}e`������{���G�r��8{����Y�[��&ވ�7Ր_%��k�U�~Bɟ2'��u3�u�w�^�4��xn����?-F�� ��X���!��N��7ʭ��ڭ�k�<qxj����Xd{��w$H��q]K��rVw=�ct�����}��a��!MCgj�
~�=%q�H�j�V�Oz��s1����ؑ(k�F!�¥@T;��m$l4�g�)�e���V�# �����^��v�e;<�J\�9���:C"�`v63�+j#.�LC�F�J�<7�[g�L�)��B�����;�L]9�ڼ���Ll��D��X���r���`h>�N�"��wQk����/{1D�׮���(�ڷkD!n��>5�	��Ɏ{7�t�����遯B��U����jf�!->��~�^�֣_ޝ�>�����&��=��>$u ���?{�cH�s��g�>}�d_E��h�ڻ�˭�OS�۩(�uױ��M�<�,5N~��7Oy����j<�K�B@u�轮6#?*	"%{7�{����ʾ��)���u*wc7VdU%-n��%�(�+�<ev䗶��7��)��r%mS����B�UK��G.s�֖V�m����6��o+�a��� ke�(�jA�nd��n����6����\^E{S^C�h�y�y|#�Z�[Û��W�{��f�,��p`
�jފ��QH�Bȉ�6Z� n��>�>��jv��+Wg�͊��I�X�+	�F61e�E�z���#����ZZ:�Q�:q�ʣ�����G��	J�.�%`�4�XkO��Ԯ��9ϷOەG�H�uQ�j��|(�j�LV��1�[����c�_<�pJ��������[�!��{��KKH��<����d����J�(U�G\����w�����U�.`�i�ۈ	`a�8�\p,Β�hkod�J��\y�ԡ�w�Sl��V��N�M3�KM۽���wwGm���K#�#������Ջ�U8
����:�*9nj��w�\f�4n��j�u��oe�oM5�osk	�4�a�s&SVW3�!�q��Ƨ+kD4���~��/:��>	�˽���'��=;N�Sɻp��v:Cw$�z�4�b���̜�\���.�w�hvQ@���b����ͦS���U�YsA�#8���U�d�V9b��5X\0<���n���%��^�R_n��3K�VR��3���e�nc�p��U֖�&�B?5\:z����,K��R=�w���Zm�א��=��Ϯ����w.�(Tw:�KT������N����
�veZN$6�M�V꽙���4���w*�}����饗2KV4`�z.�Ur���5�e^�dE�he6�V=.0�=1p��wa��:WR�g��;h:�o"���mEC�����`sJ׆�jk/<�J��'�*�:� �ɧ��P���ƥ)����Y��=YR
,�v/Q�Z�������S%�3�����6e7��-�6B�m�x����1Cׯ����zwJzbU���~v�����5��;X�VQ�n�������4[�K��r�����j ��4n�����E5���9o*�R�oS���������[Ҫ��t��ṇOr�a��Vk��c�i�Y�S�������9���2tx��E���e]�Swl���b�dP�v��O���}ڑ��+��q�6�1����U�Y�{R|��%p=d�����V����7gӏ�۶ۛ'G�ֹp9����:�����ȱGkK檺[����,�!��K3�orXFԦ�J��}�Ds|�%��e9|Κ�'ը�-��N2gR7ۚ�dy���CWf)�=���u���W�\�ڧ�v�}Y�q���lK�����.n���1jp�#��7%��pw�_a�d�5��!~A!��c�4㟠(��A�D@��J ���jB�= ��!���IR�0��d`.B�r���1�%0Dm57-���ܦ�b6��*���L�V��}f���8b�y��j�VR���*>�}=8p�m�On{�8Q���̭�eh��˙R�S�a�p�1֌�-1�,�5���Z6Q���Fb���O�p�cj�Kx�">8m�֕�AV#����*�Q7r�T���[-p��ͦ9lPZ==4��Ԩ�r&2��T~�cR�5)l��.9J�aR�[K(��r�cPU���m=4������Em���m*V�E�>��ˈ��mm���/)����KFֱU+mmm[�֖�#(+in\]j�5PL�a�����Z�%)J��ar�VƳ��UTQ��VZ���-��aT\�)Q��YiU[j��Щ��==8x>Z#Fs.R�-��2Ưˇv�mQW�c��kQ7)�m��1�K.e�X+
X��4�Ӈ�}���J�{�1e����Uq��+m�������ˎJ��T�mUZ�"�-���&�WO�����"�YYl��G,�V#iK[Q5q�ZT�kZ��{MuRl�-�c3
�m+X��6�hQl�L���AE(�
�*Vډ��|9����Q�R�ʘ��LLX���)m�+R�g�.\�Z�N���]��k��n�v��u^�H�X�*��7�-�uX-��f�^�\��%c��>���Tɛi�r�f� ~	�d� � ��Q��O?<�y��|������q+��h��S'�fo�f�'<GPFv�k���}�=`��	���D�`C���������2��Qb�Fᘄ}��p��Xʫ�m|���9�ض$n�9�Y4e�jb-�F���H���$��.H�r��~+�#���؍4;|���ny\���b��|n��x�/���[���OD�7ưʿ��?0Dč��4[3-A�Q|�{2g�g���忦h���İ7�|�g�Ր�[J�(a�c7��*��I00y��� X������>��'���^>�/?u�(yJ`�E�Q���	��67�#�E�g�q�g���N� �Q�C����}���
��/���������7�atK�g��ͿH�v���aOa�_�rJ�����������$oe�~5����Ts�`�M?x��K�����y��b�;��О��n>�H��u/�~ W}�/��khxS>?�J��Rي�Q@�kiN�g��O�L�c<c��a����lfn�g8�,n:���.��"�c�����
� x!����w�w9���,Զ�����Y*���&^�Gum�S�]|1�kbfu�a�|���]��ZgV
|�!������P�lv�S%	6+���J�,@�cXJVR�rۇrн�Ӌ�v!��w+�Ǌ����f���'���}�b��4�yHJ�G��W��2AA$D��aG�����\�~���l{`���GS0�	�	U��'�f}���џ	(3�?��a�ˏ���w�}�O��5,z9�.���z�3y�*�h���~�6#�՘b:D��N��yP���?y>�^�X�6�c�b��m��^�Ƣ�Ŕ٬O��'[S[RE|�N���s��f��W�
`P��k#c��N��ଈĪii�'j���j&��w�(#�v"т�����ܪ�K���H.��A�
��  ��^#cwʅ�SKH�/O')����~�瓸7o�)_�Ϣ�<�j��0�]}� �O�1��C�̫1��P67��
F[��9y-N�ek�[�Yc�|���b�E��.:,.���`��P�g�:A��\�x���:�V���Bȋ�E��A:k}�⌸�w�ۚFҘ���H���g���Ae�ii_����ޫZ�rn�>�����x��۴Hc2��ku��C�&.���>����0�l�D)m�;��}��<�=���P�	��E}(m��΁Gp�X�M��K`�XΔ���_�+�+��.7�5�����}��`��栣8=J�ޱ{�u��[��Y*�nZ/��y�C)�N��'c���%��a�7{���,��Ӫ1�`�8f��^J�T+9�ZC��a�,�N���M�(����p'7{xE��ڬ^
�`�Y���
�/)�܁ȏ�~��_����o��C�I �# �	�"0$D��ߟ3���ϯ_�m�fi�(C����=מ(n�`�wS9���bǗ��q�"^�킼��9Yr�,c�@�5's훃<%G���J��'�9�7��H�T)Ǉ�1F��%�
U߶߫��
6�#c��b�U���⢋��.���=��p�yܼ{��X���:��>`�37e`�N�����>�x��w�[��6 dh�l1ِ�.ꑖ=���>�������e2���%TL�&���#���$Y�N/]����俪��~'~o��_������=]��c�/��uv�zt�;z�c�9VT^������Ez�go}�_߂VXᬜ0=�Tcǫ��F[9"םuF��a9P�VL���
�Z���_�*����˩>�0�%��n�y�/088M<�k����=BԆ��N���#Dtu]vY�[y���{�*��"ߤtR6A�C`p��~:�j<�E�P�p.��A�{��U����:�^��Ӕ�9G-�Bʘ������@�85Bk�%3Rc�ŏY�E(��2���� �{A�%���q0�7,޽�;Z�W%Y����[Z"٫{?Z4��#�3ل��Y��t�����-�X�t��ʹ���:X�zF�}��Ι�ى�����Ff�y� ɽغz*�[➽�ݧ7Ox]����OY	� H��"���$��#Dd��]2���~�zk~S�ǿ:V�c3�wG�������"�MEB�aWH���=9;:&��>�W��w���.M2���	``�{����Q|�ϼ<��(��$��'����^��ӯ��F4K�v��J���o��GP��(wJ@�(��$�bv���͏+����XI�wۼU|Ǘ喙���*	��� ��V~�P��Z�^m;�З���t슱�����
�����,=�9 �y/�~��p�ʡa�K���X�/sw���p_��w�&~S�k�~U����
8&�����Y��Ve�P�dx�5�Z6�~��c�:}����1�U���9J`v?�l��B�{T�8��V�;U�,.���(��b+h�D^k~�M�3ꌸ�Oo�v�����^�}�8X�}Y�`2/��6p|�*�hz���}�ӱ�,��i��Q�=�m׸K�ti�:b1�����!w�q�zi�ς��^|��ð��[�s^�T�]틩���Qy�2�$����#�dT�Q�m�S�zL�*H�7�[g�L�)̘~��c����*��&���<v�A�vF�9�n'���t�al�P&YT��ϟM�I��%��]tkv/�j.L�5Ġ��n
h��κ��K����ƣfv_)7�-�Y&�v�F�J�Pz�i�eW>l)בi��7���.!�����q9�p �ʹaM<r��q��5\d	�0 � " "H�I" A>�|��ŉ��$1>�������6}?��'���ℸۤ+�#���Q~+\�Oλ=V��ٟRy��O�h����߃4�o������d
^�{�v*JE}��.NK���^���Mw(��5	�XY���ѫ�l96��a��z�����F:~!w+T~70���Ǽ��v[�=��wb���\+]~�ϻ����J�V���*���ӄ�ml������J�����J�kܼHs�����b�i�k�oB�Q9A�~;�]__`����(�b�����6�og������^�b���%B�v<�ц}�U�'�V�d,eU���\�\
�s|c��n���<ޖ<z-���� ������ض�c�PݠuOݸ�NWg��Ⱥ�z^����a�Ê�"��8��5�U�
&~`�@��=**j]��;9K�����Qm^��E�&�5���ĥ-nn�ҩ�}��2�hY>�`��y��Nz.	�0󚜉[��wd;�e��|/����x\)l��
;��	��`���C���dk��������r�������s��yh9O���N�ѻ��G�ra��ë	�p��ɑ:����!�W���9��Due'\3&9��ඁk�w��2����<�j,M����.��1t'3��[B�Z�jkP�4�ðoׇ'
zSʾ烾g�y���?�$?�$�$$FI" !��0�D	O��<��~�iC>�Ꟛ�TEIr��ek�5�~-�����W�l)�>��U�I���G����[�RԞ�"
FP�4���Ȯ����\�Z7s��=)����w�5�b���1��c�0qT�1�a�*kԬ��p=��]G�����٢����W�39۱�=��˞��x��V1�;L�;9�w�"_O���l��$��5�b�n./)+37���Y�{�^s���k�p��Χ쏣�`����A-�ȃq���xc^ ��`��9�w�m���&�3��h`�}���u�w��7�n-�R:+�hm����xЮ��cWs�E�~�U�����U��(�<!�Ti�Z�kہv��YM���B����3 ��$<�wJ+/E�K����h���pFЙ���~�V1b���Iҁogc��n���rY�*G�\P���.�Q��������u@;?)p�T��V�_��������|Zq�6vbZ���W�op�?�Ӱ+�C�_F ��*�X(!	� �.z*A�*�����֠ll�1�s������?^�mH�+�x�α!;jm���ف�A�ћ�$!�����8����u|7Z�v�}^*�>�0e���[#��m�K/�wv�������O%<y��9�^ꪧ��Pyr,6컥�s巿;���~�'�I D"B�A�D��!����wy���}S��@�=;W��1[خ���H�TX+��"Lp�����"Q.�R[x9�w}ϴy�Md־�Ֆ�-y����Ji�)��i�ʪb���W�H�(��DϘT/��r�c(7䷷�<�18z����ڐH�zo��Hh�BJ3=�����ϔ��,�z�~�=���ρ4)�g+��w����gc���XΔ��Pb�W�\ml�'�q�k^��v���꜓�����Έ�^�b8.�l��Tdkr��X���^G��f��-ʧ���S2�1P�WR����O��8f�ƃ�?g��=��K䇷2�_x���U�1z�s��ИՋg���u{M��1B�A�aNEE#�!��y���*=+��"n_�!��
B�%X/���iаrs��e��vMX#��S�d�뻻vWf��*E�5�~�+����M����6_��ᦩ��{""���}�^M����`���Y��Ä�0�[��
��B8}�~��w�I�ޛE��R�n��a���E�DzA�/����FT-8cv�6�2κ�Z� 4��BwE�W]���bope�����*��Z�nS��/]-���P����xPC*0��k�!.�h���[9���j8*�l��F/OVZ�lY�r�'�H'�UU4H
�ҹdJ3f��� �+�H�F@���"BDB|���+�9��s�M�@�?�78l�z+���c��8T�ص��䋰���6��
G���^�˙�?lE��� ��y�rT8N-�v�	��q�BxN�X�*�}R�(еm���q�Wg�Z~���D=|���TUe�����F�3�zA���q�==&c8�cP�V��>w���[���=[{��䩣�k���u����;ʈ]̂A�ØLxO#7I��'�j���Y���q��Ɉ��`Y[���������O#ѫ����t��ڰ�ʻɷ���w�E0X�:�	v�$���3��P�O�m�����^�lr�����q�9+�8�=ʯ;�w����<�h���p$̃.qQ���Gv���7�u�H�B�����U;cЅU߼�����Q��)���c�Qa����=��4���y��/��*Y8W_ԯw8'�#>ܺ��LV�ˇx:�r�1���>bGS��}>����}�/&9�k� L�I��k�~�����R�6;Ց�bo�՜}f_���#����Z:���~�n��st���:5j�j�N��1e[CH<�vl�.�קE4�~�n����9o�R�\w3��_��+5۹�3t�)
tUДT6+aYw"�N��ɴ8�j�C4A|7 ��J��9XV��(�ٸgr�/o+��M܂�C8aɨcqm�k`�f��{�r$�e�D�wK�B��H� �H���� �B"@��	��?3�����>{�Z����������V��_w~�=�S�ߕ[8���Ӟ7���8A����p�ڋ�������D�/�j$n������,��ȾSP�8��\<���N���a��c��΅��.���xp�G�M#�p�PB��R�`��-�)�e��zd�q�����UK�Q6r�߲~2����#n�G��`=�RF�TٍUv�����k�	�W��˨[U��k���5�������~Q�;*ԡ�����=��칤�rw����bՊ�m���q��HH��:��(�����C�{ #��5��x^�%����3c]��7K{W��_F-��!��Ò��<�#��b�}��8���'�h �!m,�޹0�1�)�<WT�������3��*3�R�Yn����Dn	�&#N�F:q~B^� %�}�ޙ�v@���hI�)����}��cϔҁ��3����u}}���y]��Qk,����W1��bLz��tP�
lyW	,������l��T@�{"�S�z����I��w���ϛ��?^p�0=����Z���:�mH���&:�Y{�F;��-�n�S��Dtek,þ����Ϝ��,����%�Ͷlߊ�����<��v��c�s�su���,�=ݚ��;%őU0�*9��$h����7"9��j���LFY�D�Ϟ� d �#	B ����_�ϙ�������o���o���%�|��"x����9Q_MK�YR4io>�"G�5I�a���9�w��vgi�y�l�raF�*H��N#�6exm
&CLN���%��و��}����{s�WG���V8�O�770��z��Xo�\���b��0y�C;�U�l_:���J3{��]x�;N]�}o7o�^R�"�K���!>�A_{k!�ޑ�x9��1�nY
�u���+���h=��TC~e��)՚ߟ�;<��e=�q[�j��.��w�4�io��(�1�\�a�1�
G�xM2=&Q�հ���;��b���w>~k"��ʪ)k��F��/��ہqkr��9%�O��*>eH�-�ᾣ(w��Cl���9aM_
Ӯ�W_t�}�󪾾/�7cv��cl���쿫�L?�xc_|���?l�;�Ns�;��;���o�.�����m�W���(��[6�a6��O��
�H��DJ�T�{O:�㔳�ے�8��q�� �>{�1]��򛆾-�R:�U��!AG�� %�����]â�0G�͝U����A�G�p�)��Y��eM3�����v�ۘ2YN�]��]I�ѵ����,辺w&��56K%)Ϲd	�CV�sWVql���[���#m�X�j�vY�:��
ՙG$�d�Ù���;R{��ii�f,�A���8�%��},T׫q�J�q$����oH���͜Y�*�(V��\���|{<FȨ�'�c����}*��65�}�se���ު:x��B��q��{�[n<��&���V��} ��6��S��u"�+n+rU���4��{���.%�����DY2u���h=@���8+#�C`iE*��+���Z� ��_.hn��pL�BT�>�w�Ž�.��F�JO��P�[�(1����ETXřb.x����R=\r8�٪��E���;ڼ�}wY����؏t�˙u�����Ĵ���a�E��ܙ�$�x6e��F�Ny����w�P["�!+MYs��4)�H��O�B�槖����^*��ʒ��J=��o�hk3�z\J��ݷ��۱����`+��k��%9gPT���Յ���6��0fk�Hn�a����c���Q�)6m�^\ǘ�.��R���F�J.�wM�k��r�4��V-��$7�uܿ���A�{����۔!���m�X��+Ν�S����1�Q6/&*�8��^���h���25�Ai�OlJ���G�3�?*�c�;�J�����4��EVs18���i\�uw9<�"�E�1�t�5r�\�G��[�L�L�'�Uk���Jb=r����.��׭���/I�&Fk�Y�`y�{7*�#q��#U�;2.���<̖ ��ʕ�ӣk1����}�u�p�I����Վ�(��޽��B��v:����i��_S7�������p���U�u�8��}w��&މ}GBB����Y3]'+�S�!��1(�E�Zm�h�s��dO]�#>ՕB��*��;)�M���o4�U�)7��u�\����
A�|�#�=���<�`e��"kw����ِ^���&:�ɝ�!��bH2�U7� r�Ϸ8Y��{��Wd`�hvq��q�麜�{*c��F�]iH��3�M��.���6��{x��e���\�]g5������X+ok�^G}zŖ�
u�q(#�i����;#2�sn+z�S��	9Y��g��9;]n����u��p����b�4��W��,7�ج<�]fì�8.�4;���]�2�@��W;�K�_e�v����e`�9��V�W�L���w<܃��2W'��b�u�@��j﫶kx��诋�&LfU1��[���ksjgmɳgLI��w.ft��;z�=&��݈F������*�O�}ɘ]�0L���2;Q-�q�Js��X�h���[EUQR�i����2���ku��Fۮ"��yvee̕��T���b1�Ң�VͩD�t�!Za*4b}I"0X���ɎZx�9���F�s0u..��wU�֗2�3m��,kC�2����]�'��=<1QJ��U=�Ow'�޷�����JڕG;u<�&S�͢��Fy��H3���ڙKmҾ%q(��{�8i��QJ>&`S����e�_�T��\X��r�k�C⢂曍���Q�LpTm���O4���kUS[��U
�<�j��v��M��;��w48aH���;�����8a���s�x�[̵�K�U�eqQij*�~Ҹ��n�v�f2��f`^�0F�ie�T�r�*��n��DN7O|<+����y��-a�y�`��0)�r�k�h�ZiqP�q\ܢ9���kJ����Nzy3&��6Ꮃv]�r���st�w=��=<㏗�8�e�����mJi�e�e��[W��b�ۃ+��]�0�r���&��4J��Y���tv����̩KJZ6�33w-��{ �s��Ɨ��1-�f�<i�"Vs_�a��h�'үn+ܱ�:F�;����M�\n<>T�r�"�f�A�B˱s��S�ш�Y
%��C[�u �=�UW�� �! A$���$�#��|  {a-m[~����{�	<!3ti��T*ж���O�H7���X�
�ۘeo��k��RV:��c�Hu�Y��.�q!�<�5���j�r2�E�	k� �T�kB%N��/����W�eY��di ��D�u�c��Hr��H���з�iiP<)3]}	zl���}���=�N�E���+6'ψ��Bi�A.�9�8/��j�pD���
�b�=�#������o��k�d`��'y���U�q94m���tZ��o�pAT
&x)F�p=�0'�"}=�Txױ�s�����Ҟ�Dm}��P2��1M�U�D�+��²�������0I]{�ζD���_�M#�79n�@�7�{���C]3�9ӵW�U%�t��ټ%��Y"X�8�ޖ��+�6r2�>��-�5������m�/A�L�>e�̿x4"� �2��/�S����L`~!��ܯ)��*��z��dM����d���z�*ވ���Ra+ZA���
�*nJ�Pq�q�
�$��>X~�-����/�u��.3l;]\��ӛ�)*�o�[u��MVi�2�%�TLUr�@��h�2K�Ȣ�/����ۧ~y�=���Db#֊���]DU��W=�WN��R�f�`�+|��,ox��]J���?�'B}������UL����6���|����H�$ �B�H"BA��@D�BH�>s/��|���-EG���l{>�A�ƨS<�\���o���}@^��LS
}�"����
i���f�%���gY��=�b�qT)�ϑ�e�t�8-:2}^��bV�üQ;�~�n����%���)M$��G���8i܂c����l�#5���vV�X��!�^������a�s����"@��#�2�>6(�]�N�y|�z(��l�>����E�=�%B���c���yO37�u��9�*,�X�r%�1��;u!���j�k�NH�����bi�Mu��-�j��n��>�P�sP.I�Ȣd{X[��!|t�σ��������~p�3uO�r�ؽ��7���������X-َ�o�:) ���$W�N�ꎆI����\Q�m�O%A�}Kٻ���=^](��*�R�|q9H��8,9�]��΂�����a}�>���|~{�]����ސz�|:�`h�����h=N>X����}Zy������t����8-v�޻���b�N�BMq�a��P��o����3�#r�lr��0�t;a��Fx=�UF��G��Ƈ�?����8���i�ſ(�`p�(���m��Z�}��;��:��A��Ε/*#s��Wֽ�~�Cw�r�ɝь�MB��-����mtBW?H7��l���^���\��GKS��,S����n���=�|Ɔ���Pr�����a "B D	d�`@�$�H�	9��۞}�Ͽ��y��ۑ��$�PSD���?h>DPN�sż���u}�~�b��&"nr��\`�����(1��aƋ?f�ܞ�8���|1�Ƭ��Z�X͡�V�������z�rs��o	�q�`;o,0ԩ ݺ�w)i�5B�.,����<��&��	[��v�/S���3g"�4�#������Og (�{w�g �2�E����ine�޸�{�˷0;�Ĺ�����@炶o��S�`J����eҟ@��Nx��o��f��l*��,����zO���P2�F�u�p��迏K�Jj8����Sv�+�f~���>pũG�<}�a��G��1�.��PB��R�~��[>S4������ʨ�u���tIcя|��F	쮋8���@�y�06>���������REe_�z�0 ��J���O��"5ϋ��o�~��j��@货�Ǐ�|"r����.7�T�����\��V� .�)׻���5	5��~<VXO��<�46�on#����B'>������m�����~��̠E�t#G�κN�p�I)���V)Gn㔳��3x�b�W
U��c����4�r���Ϟ>�� A!���^�8��(���!��-��y�Yk�<�KY�n���i��ɕ�; �&�}���y�p�}�w�}�O�2H#$ FDB � >�3��-\�e?#��f����gk�����5c�&�s�o�ωAM��0)<ВUAs3��H,[�@9ƅ�fM��훃jl�Õ%&~�W)�^#�v���]P�Rcow�9��O=�ou�~&"����@B9�\�6���j�oB�P u�|0f��'��~ f<�?�E�>�����$��_aV���&<`�?��_PY_�k�A��"|=�U���{i^�;W&u��lH}i��8�eF�p$q�3�zO��5/�eO�!�^nHPDVgF�5���B4�������F���(���"��9ʀ�-?V�c��/E�?>�5�O\:��ם���{���7
����)M��-��b/�Ldz-�|8�W�.�EV����;��o���u#�s'�H99П�W����"��b��ߩ���V����t�L�(p�x�Y�+��-����/�6N�(F�)�$������ǵJ�g�R�/�L0bkՒ9Հ30f{9�'%(/엇��7'|>����\�_��������H�¥��1{3Hϻ�3w�3��#8��_4֥�J�FG>�:�9m�S~a�9ӗ����c��T�
��۶8�i��r��D,�+�nzf_Uh��hf�}Z���Տs������*T;U�L�	^ɳ*ܱ�]��خQ��Ii���>����T���!�� ��}���jҦ�/ϰ�۽k�||}�n�Y��?W5��,}���yW��l��ъ$�����״�38��<ޅ�>��rz7�&Y|���>wi��𝬁c������A��mz,nk۵�;ϟv=�/hƈ���1]����F@p�}Bٴ�XEM���a�7�,f���}��UwYy�L��_F4x�]�
���+�t���Y@/ФtS�4:��=裋6C^ٌ���b#����dD�#�Ԟ�n�#�J�-[nص�|j0ye>?V|�(UoN5n���;#��w�����C�q �����Zz����(�g�<,��ex�ԝ�}R��8�eL��w��}f��q���9Z	� �v:���B.�H���P��l���	�م_���?T�D'����)�����>�Кx�K��!p�C�_�1��s�G�Qq!Kɚ���۫-�^���c�я��'5㣔�����:h�����*L�
A���z������j��f|�`����f#�;}nFQߒ����*�`��8<^#�Y��{�V(B�)�{�1{*��/Ur[~��V<�]�MR�A3��!�%�n>B��r�*����m��b䖢����)��;��N�L�K+���s1��@�%R�p�$гUzA��N���tgWnjKll?���e�^�_���+����?� ��$D��$#0�������$L?>��߻������T�dĩ�@�U9`ݸ�>����B@�r�*���G�mG+ܣ���s�~�M��cɬ3nDA
EW�N"(]{����q}��W����qAc}�����.��{��Ě�����~Ǵ����W:)�~!�_|�vE�*�쑚��}�y���#}q}���m_
�3���<!�<�o�����7%^���%��*T�xeZ-���rˆ�̽���y��/xO�X*�V-�v�c1u{M��xf(Y�1,)ȱ7v�}[��;�W�{�b��۠�[������g��3L��@p����ϧ��|oN��<bu�k��؛>��;�	zK��<{����W��^w�.�L�#5�����M[���ԗw��x{�}�Ϣ(�D?�ʞ6ء�#�2�>3Gxw��;�w�N��6���n�.���:�ЬN�vG�{�Z����k��9VT_Ď�#(���Br:�C�����rEuW�Ll�}������{Z����1��r�>�&��At�Ї��������O���m��_��s�fc=ށ5����7@�[�~Җ�61P\�E���z�p���sb�;���ݸ�b��dԿ]ed$&�O�yc�҇dɃ�K�.��iu��w\�񜅸V�i��t��:��5WIa�e"mKU��r+}N�@�=f�hx{)I�ӟ<�S\��4�\�[K����$�# �0���� $ �� | t#�|���`F[P:=���Z���3��]S��^�����$1;�@��H�_N������{�{,<㮦�m���d��Z�������2�ȯ�>0z����]?t�u����2���]��^��f����_I�]鱾u��Nfz��	Wէ9OG|��G��x�/*��Y�9V.^��A�b�D;>aP�~򟚜���?-��d���ߑ��G�ؐ�_(#G?D�',�gl#_�\Q��x$¡�*�
h:�H��^G���Eݻ{ �[������6�������C�L(�����=zj�**+�=**NCf��Tj|����|�#=��誔:�v�&�Χ�����$�=X͎5�b��Pd`���p�a�9�A�a�SY�ݐ�]�¼_���n�1�S�?Vh!�&�����qx\+��]2y�'C�M����s~��$A�d;#_NOԧk�������`J������j���s����~��[�ާH��!#�/�
�$4}�hp����xܰ��3�	��ut��2�h9������p�63Mp�!cU�
���4z�UI�N�kt��k�M�NU}�O%i	<��Nfoc+&ǵeŬJLT����K��&���ԑ���[��)ѡ��3�a qwa�X��bΔ�3��l�ea�Ó64?�|�_�D� �� � "��  @�� �f-n�l��wJÑ�3�Y���3AH�2�H>�ˀ�(!]�\c��ٝ[��x�$71���\�g���3X�������d�Ac����~��a��������0$Ǹ�7a6f��x�VE=�ݗ��|�m��#�Z���BGߏ���w���e	q���b��^K�r���~�]��F���8�S��Q��~�y�C����!���;�' %��[NGV���f5�]��"�GO
"��o�5�����״ѫ�Caɴ��>$@��TLg�w+R�Ҏ��f���(�5���9�Z��jv:�\u�u�3u6Ty�Vi[��׏`���F|�i�b���w�C��A���S��b|��D�
F���ј�>�Ρd}��Gw����i֔>���:3$�_�K=������P_�Ph��AZ��J�QӞ[�d���w��v��	�4|��=�t��#�=5��lGn}�o"��E���?q�3��JV�.+�H�ú��*}��K�䉷���k��s�L��z5`�YV�_*0���$PZ'�2��!�&�l{�y�ٗ�|�nD���\T�RW�<-�ɱ7wa�zp5,e�ɚ�g�w��a	߄�+�]p���r)nK��q.���6�ؘ�59�^��@N��
t�\���Ӄx�d�OrU���:E�+���pR:�쩲mq�$�;T\6	���H#$a�" �}�@������˗=}�<1�~��#�S��=�?o��blwSF,7YE��c#�l�q�2���{nlmSu���{�vİI�H?���0�;��u�������#B8~�i��9G��L_v��x���йj1���|i&pt�{�%3�N�2��`��ȱ�PgcȰ�^����S��4#^��O1z)����Z�C)�_P�	_��,9�2�s�ߞ��l�_{N
��a���t�e���Lo�{O���ݫ�;����z/�rK��D��5bT|ˑ�*u�Y��-\���6oo���c����R����_&�c��瘙驪^@Tn%�uz>�}s�u������.�rP���l{J�+�ݸ~FC�	���ͦ�����O���Ngr-U��;�>��'���9A��Ii{�*���1ީL�)�|S��X����e�IsE\i����,���Y��9���P��ti��T)o�m��^�)�r٢5��vռ6��;��F���D�4��k@�7�Q���q�����c �����N?e��wׇp}��wCz��/�n�7 I���{��a:w0�yad�ɚ�u��ʢ;��n�0g�P����M���g�A���K�ۚ�'�����w�zG^��nA�+v �c���-��_vnL���]��iY<��HJ�;#��d����@��	d �$�0>#��^�J�y?]ξ��o��S���WKMt�Pj��0���C���%/�>��i�?���s�����\�zkt��K���G�}nT
�6�lX〞�,P"����]�"��`���4���*��?q�1�[�8;S��3�"�s����WRB�1�Uu
&��P+
�R��e��h?��`xC	���=Bݘ���Z�%4���!iC>F�ah�9�還7R;���Uiv�P�:�ԢOG�H<|�S元R
�~�nQ����7�A m�D0Ǳ~�T��w���D�z���{" �9LN"�-���Q�}?X�T�¬�m�Y%*5�~�z����;}f��,�/gq||�5�Ίc�]�򺧆��ܫ��{��U�gُx�KQ��z�q�,C�t*�m�����
ʛ��l�p�c?Wα���N*�"�F��[�����߃f�T{]m�tG1.3RC��V��e`zbe��n�OQ�:xx��������H�?Da�I��_�Ev:�{�{�f�� �(.Zv3'�� ��ɿH�ux08�T���U>���D�ޚeCl;|]^�S�EGx��ڵ�Ԯ^�չM`Z�E:R�n���rvy5�쳓?j�M����e����K���rZ}��Ҡr[�Kx�zգtw_�]�,�S3V�+Ef�lh��5�,�#�Y��@�Sa\�w��J+%�� E;������bp��5�F!o{���uo0�aRy�q�;��5��D�gJ��+/f�wf��)�gJYZ����s��g<��nc6��pЛx�S9igf�;�,
F��LV�gA;����+�f) GSʣ��0E8��m�ȓ��A�vt��7(c��*�������b�Wh(J�����߶Z��ϟ^�bs��]�6z&�5/���.�J�����e�����:=���n�J"@�y�b�9{��f��5#�����x�M�u0��ʇw��b0rK�&T�j��b��o�N�[� ����k\ٖ�h��K͖�&.�����dx"��B���!{Q�Y$����{�z�;��$%���O.��Wͼ���&��fsiu��m�8Q�8��Ȭ̈́+�!���-�\u��;�;���c4�:P�;�v�s�e����3��)Ai���Z�}�M�4ն3qE�ßVl���TW�%T�[��W3��ܚ`�ʡ`�f�R�!��㉱צ�5������`��"@��H'���J�	GV@����I��!$�k�Tq��5R�R��x�H�)���g3Ք͗�n��[���%;�������EZM��c����ڢ��*�IɅC�og���[~����ڈ�p^`}uiR˱�gvࢷ��s�_,"k�x��A�[��n��v�o5崘�9ǜD��w�m���ĬU��A�coh]�	�|+���\����(���09�v��t�m��-+fs'���o�.n��.���O/	n����X{@�Dû��Y�d�u�.e��SB�Յ��S})��a�u,f̥�S�����Ɋ���%�9JAK���N	�֘���އX��\�{�p��[\1L��v���[$���[sr��H�QS�.l��k�G�S'��.r�5��V�ۜo��]�����Tכ�Z�q\������φ��K����m뛙���R}�J�-�{��»em�^Y�>�@V�y�f�J﷉�N��$|Ts���G�S���м�9u!܍���R�>X锆�b�}���v�%�}W\���,�Q5��Ïq�!�b��۰�����,'���	���ݾ���U.b��ḰS��r��6��Z@,b�5��[8	�w�y�dOB�\Z/ue7�t�ݹFi��]�%뺰N��&jG`q�|��+�N���w���zm����,޶"q���ȤѬt|��qA�f�h(IP�P�D	��UZL��$���3�#me�WjĀ�D�L(rY57M�`H<,����0�ID틍���Q1#x�ź'�F��c�s+l����<�]��F^^:kJZ��pMَ,������/�i�(ع�8a�O�¾5�q8:�hV�S2������h&�(0"��c�&��?�8�$BB�����nfDc1��zxa����:Rѥ��m����8�r���^sx�je��p�Yn�ܺ��h�$6[E"�CI�B�
P�nT�s(��f3�Q�Vأ��3P�)�31D�-b�\�G\3qj89���}��4��o�8-���ar��r*��Y̹mb�'_*���˙��a��m�S1���p��m�|V��J�.s*&��&��V"��4���� ��ʤ?ӵ%"0AB:R�Z_-L��g0�����&T�FEG����A7#�E�e�q��۶���ӆ�p�i�|MX۹�=�sN�l*c����Ɖ��w)��̵�]��Q5�d[�[T3fSZ��m���T��->t����r�L��i���c15��]��6�ڠ����i�Q�5�kQM�g����>�¦�ZVx�O��4��#Jx���ַ4����Z@̹���PD�r\��ۺWq�1��9u�P��A+[0�M�Op\�[�n��=��*���$�4��wmbצ�kSf�J`��-to���]��]W1^;�[W5,��?Ħ�f6�m� ��O��H0 �F@$a ��=���ߟ7���'/�.\���4��"��`���3@w�B�y_��/�Z�0�N:ouY���a�{ϐ:�X��?��O�K\_��B��@e�_ ��!����ފ�Ԥ�E�6��􋠆"�wU<��n�a�7���r*���� ����`�~�.:�C���V-x�4�[��J���w���}$y���7�q��NT+�I�E!��z���� �2����BRi�;�VXk���ݝB���c�j�|��`iڣ��������� �� �N��͉�ꎼ�F�>��o��y��o_�wѐ���K��L�n�3��.�����DW���o�����w�{�Ԅb��2��5&8�6����򬇁R�>fz��J��<�OF���{#�B�~ta�5��Y�����r"��'S�*s��a�z����r=���*�;�S�k�������d�&-��B3�
�_�HM�,c�d����N��EM:�pQ��wX�Q��إm�=��&�|�W�}"a��u��!�%s
4Y�6f���βj̯��0/�^8՟�M{��l�|�����֫6�F�^���v���CCz�\';��.����&��+3����Z�����Lc�P�L<��L1wI�
��$~�tVu58\�s��*�&��A�v�ǃ"j�eƙb���b��΍֠�y���n��jZ*��7�s=���?d�I � F# �d� }��~o�|������J��u����\D����u��Xb��O4�y/�C����
b��i��t/Foez�&�o������Yܻ���򜏴��#���1	�n�	��������xgd�R5rB�c{�s���ǁ'���� E;�z4�����KE8���qa��B�g��W�Z�#�"C%��q��FRv��'��d�tc�Z��>w�`��Ȱ��6L��{5Uqv��{�7�^��Z�F13�>�G �q��d�i�Ip��A
��K����Γ�������w/mN:�t�қ�5N.8OetX>�����"1�S���p?*�g���>���I���|��7[D��,o���J��>
f�O��-X{}�#�����тb����\OUZq|v�I��yy��+���xF��]� ������Q�m�k�v,$s��A_�����&{�=֓���4pl͛{݉x��p=='�"��-7��U�v�ؾ[M�t6�N{���G[	Dz��8�~ѿʿ�w�-��'�O�0$~�?���0�)�bq{�	J����ԙQ��R�\�]D^�i�b��m�ՙw�?�N��ψ��3j`���!������#~�HzE`��Z�n*㦳����Q���<=f:�)c}h!79`���M�݃�Q+Vq`>|֎f�B���졎B��R���L�VVo��<T��u�A�Rn)F_|��@�� �����$}� >ｨ�Z���4��)��8LC���1�	1��b�i�o��z�G�~��uy�:�N]����s��Gܧ��)_Ez���Xc��@�x�(!Ntz9�3�*gz{���������ٕ�|!(��r���w�懋�g"Q���	PbG��Y�9CtBp��)ҹ.����|�B�w�b4׻��XJ��9Q���:"��>G�zm/�&uu?
wO�-�XX��J����`��C�=N�R��]�n��=���)nn�U1_>�A̮q�B���TM;�WUo���<g��d��'�����˼���n�͋�/�_A����V�eIU�6�§v4O^�b,��jn5����ɑ�H��-�s!�c���Y��?��VO�q�n����~~,o�T>K��v�Gz�$��A���#0DzL��[}�[�/�#�n���̮�ϧ�o�#L���ݽdc�V��>��/��d
��T��߻:��&qf�oc�1^�'cp����g�`�~	�n�2/�{,�;��t���i�@���4Pu��SO{��Bv�����3{S�w1'����+��3YWׯ�R�h�Heet�D�Ʉ��ky�F������}3�=��h.����[�69L^��z{دn=��P!�H(/�*�|��]˶��η*u�=~s8�y���3����� ���DB��B�����!>w������`Jq�N""I�[�a  �}��W�)WS���!ByBٿ��zU{�d�B�;r:1e���k���3<|!���W�l3�*Bk�"��y\�w��7��!��
GAmE�����ӕ���s�t.X�n��%A�2-����w�g�֬Y��p.�^�ƾ�|���9�Q�U����1t�>�P�5�0)�$H�I��ϠBd8�l
5��Z��\���wF�S^��M�Dk}j�}]��װe�� ����6:<$)p�VOyQ��W����Y�ײ�G��V3Y�+�w|�Sӟ')��S��KlV���Oq8�&E�}Y�Y�&%ޘ�W�[�A��� �H���b;ջ}b��N�B�z�r����:,!�F"���SauT�L�B��w�WuH�/�,@�z�z�!��n�F���_@���FE�����UL)�p�*��6bg�@��5�FA�A�&x[�v4M�BM3��C[���tPݟY��ʫ];��tL��d�ˑ~�_љ�g�rt����,x����#���y�
l�)�9�ۺ�?�������*��o`ӄ4��s���ӑ�$XhrB�xT������3��<�%9\�R�m� �ي��前��Pj�t���=b�;WY�[õ��pa��8N�"�����Ͳ`��u�M;%uK4\{��sp��w��8�smY���		!�" ��� ��o�\��֣^P�_x��S��O(14�衜+p�ϕO��O���	p'L��s*џ1�M��qswk���?��cۺ��`4�>8����y�v��ctu�@�I�^�2�������9�}�#^�՝ۖ)�1$O���}�V�G}1N=�%A�ƨS<�z�`]^�9�<f�WQN��/dϻ}�[� ���J>��#�����_w��`��`Fi���@qbZv1�(��]Eh���\�/��v�,�3���X���p�ο�nػH��jo=�����B��~��F{(��#.ei��1K���!�%�WI���imG������`�y��>뮅�F�B��jU�4�&�,���.:Hq¼��͎���so��+�a,��"�*�8�y��ʄ�}JpOF|?)�f}���,� ���î%�}���\�V���}� ��u�M#��@Q�lbN�gt�v�w� qߑ�p���,w�8|<~1�\�2�W�3{dW����G��
��=�qp��`W�0���9�G(��碖_1ڣ��f~j����~�IV�1���,.��W�V����yJ�٠��k]Na�bQ%�� ���`�%hT#��/'a�g:��U����ۥ�RXJ7�������-�dy������a���u�'��|����w�q`�@FD��$D"$��������������o`�.�aP)I�.+�1����쇝N�,fy��J��zV�T����15�g�A4���	�pA��H�?!����$m����^%��5s�5�4>��w��4bn��޴In��o�SR�7
:�0�����c��)�v��3��O=���0�L�[��F��`_�`����PI\�|��?V�ܞ��,��&iI�@4r^�}�㬿��Y����qc:،p<��r���V3c�a�������(��N]���^���詑���U?K>�NEm�G�ʘ�a���Mm�~��m+���;6�ko^X�C�:)>���d`�y}>��]+���[7��}iH�ĩ�x*�c�s7զf{ �=�bhr��s����cGF_�&�eN
��{A���}X=,x9���{�z��i������MB��Ss�>��Y�8ME�e��R�:�h68]�+ۆ�[���%�z{��9�^|��i�q���Bv;�F�~���1e}�'�o�A��E��u�r�w齃�$y�4�o�
�at�,î��XP�ǽY�?s�p��Z�
�s��*n�}6e�QG��J�s.i\:�p�t9;L�;�t�/��;�����]��Bݎ�weŽˌ�Y���Y�3B�kӍ���Q����@�D"1#����3�jO�ވ��h����#����˄����3��tXJ|��PC��;��u�L=w����E� ��N=�:#����y�����߹N3�9�����u\�����(�׎��/&�ݝ��������=3�\9	�9>)S?rίJ>�;z�/K�]���&�s�Nͳ5�h/3��u����|�D�/���!��h!sW%G+����q�������� ���U)�Vu���+^�2"�&6�@� k֫�����e~��L����t� }�=4Q�-�G� }�V1�^<b6#p�������(	��6���K� �c��瀚v7@�����GO�,Ӄ}��ព�w۾�yn0�v m�;L��U��ȱ��uǅ��	�O�����V�}��X1���=�#����b4���Ji�&:4r�$W�D�68�|w�Z���3�^���E�AIb��K�S����V���O��bo��1m��Xb1���]@��Lh1���DۘX^i�}(`�d֬�傪���f��@��(�#˜�Ѥ�o_����ں���)8��S��gS��ov�1)�Ό��j�a<�X�L�9�o*��2��y�`�e-��{ց�Ta����z���($��E�y!���=՘�}��.�:$7/��Fl;R��mܶ�>V�,�A������DQ�#"0�����?;����o���@`��>�1�b��A�qP�������(]�YTt�$_��cN=�^Bз�;j��􊆚��ϭ.:kځ7���,9�'�#Xev.vm�>w7��3�NQQ��ޑ�T���e�TDSwJC{���9*R����GI�Gz�q���k���+�Zb�~��R����E,���n�23��|�k�-�nڨ'�/o���{>����<!������N�?#!�c�S�<iؚVװ葦>�;>[o�"�TX%����":�}br*JAI���5ޑP�w��}C�t���n.���rW++;jO�*�{�j�p���x>�x�"8�2"n+�~4������J��1�#؍6�5���z3*�ѪV�w�n_q�o���ʄ��s�2H���� Hq�{�F�j+#��L#n���r��9��]�f&�@��>�8��n���F�q�@ ��#}ʼMEz�dk{�vw�Z��#����ƌ�PF����9H�X�>"m	��%���#(�׾2�}K�Ѹ{�ڽc0S�*��ٶ2Ʒ[%��d՜�䔳Tj�2�I&m῵?�5,9]N��͢�*`���].Ě�y�"�׎jO��uݣ)�v'�vV��Va�����a�z�tɘ�a�b��l��`����"K�D�n�h���b �0D"�4}����!�F��c������[�g����B�1]GE����'�/��~�[��mv�uȃl]`�Е	�*LCG0�f��v�ZSH�b�^<vT��1���e��7����D�a#DyO�>e�?}c��f;*��G^�o���;��2��/��#��f<�'#`ј��A��E9-�7F��m��6Cd�&g��誗�X}yKF��-���.=�.�F�3x��
dW���vw����_+��՗w�y�G��t7e�x���/o�^�YSrV��Vu�Q����d��4z}$���G,���܄��J���P�]vP�7�z#�Z�Q���:�u�Ѩ`a���PdU��R��#ü]t!R�q��-9�
,����ˉ���y��bG�UD9�[�x�9��NI�dHE�}$6{ �8w��]�M������;��5��y�l�[�����n�����\�+��ZE���)Br�n��U��"C��i��P��u�ޱᾸ����+�x+V�{�#��
$�wE�˲$Q�ʻ���4I5���=Wk/f'�>Z5ū	�͢��{V�:��,�*�r#l.^�<��؊�˒��n۸�t��\��W>ј�.1Ľ�wk�Fԇ%L��{m�k�*z�Dv9kL�i�d��/;/%չ��}�� �B��@��:�s�qO�Z�Ӱ�h��t�;{�:ԯ�"4�7�b�C;#�ft@-Fkfh^�.�cck�B�{�Đםu9h�fc��S��ƑQ!l����Ӓ!�U��k�FC�����R�twkہ�;To�s��:ǃ��
,�.�t�к���a�yr���=}�����۱p�z�s���)�L�4�q]��\��;�d-��p���$N������t�>�CR3��Y��Ž�, =���=��YW�?t>���6 �W�" � ��KD�Ǒ��s�"#8u�Rhr�:*+�k��Z����b�'�;Ŏ��u�����394��^!�_|�s��R������o�+M���������g�lF���	{�@��:�	+�^�k���#vC7X�O����ޞ�`��������f���n��`qh)��P�9�Ci�+���Xo,1mR�3��	�� ��lå����}��U~��Vĳ��TXu���F�q�7~����U�~�F�
۬���[`���>� B�Nc�s-�=?�l�5�sB�&�d�P^^��a�W[r����idΪ�1d����ޠ���Gr��ڹg+y�w/(��S� �;P�x����ncb�Mף�M�Qɲ^n�e��vR�Vsr􇛇{�U�U�)��|Ŷ11��X�LleS��zq}ܺ[5So�.)n�]D�:X��Hh�f��͏b]�ojs�%�o38���Fj��11b�E�E(/���i��V��w�����{zV��*Ԗ考SV�V���o`j�U}@V9t)$�+�.�@t9�%���g8k�RgL���}�Z�u]1�wI�:r@4W] n�]�i�aɑ�\�E���w:��)�ci�+��;�5PSW
Auh}X�@��ޛ�/o�F�eNiu���q5�i�|�_{ �C�5�k�=�Jalj���)�z�������1km^	B���������,�e�H��)+V����K1K̨��V��`�u�pn�yޘl��H��~�Ҧ�
��os��p��,��3��NW10�g:ەӔ�V�=m�Ǒ]ؕ�N�Q��6F�RP��zP0�W0f�dVF�Ҭi�uT:�����������j=Z���d,�W|%B�;����$q�}�XQ�ah5�Wg���u.�[�ĺywh���KMΥ�֔h%�&[�h=����XB��]泺�AH�\'�n���W�gpЌ���RU�f-یnO��\�s����(���뉃A�]�P;.c�<��i8�x6�W�帷�����[��靑�FӉ��̜L�w��ra�T�B�'.:���Y�\��:-}}}'5��
����:�ܷR��ĵt���moTA�a��3���K����tw�I"��(�w;�Nˣ�)�����4"�⚮w�k�S(�ΟhX�)gM�jȅ޴�)Sp�+N�T�i��$��m )�PhGh�F懦P��ޚ��=�nYˊތD�n��x�H��^�бo��i�}U�����Zy�/Z$q�#��D��N]�l�Bea̱iB�fǩRRAHNT=,��W���,���>)�5}hMo���i�\���ۓ{W돦�tesk��{.n�q����N�Bh�պ���N��7�(9����J5��n���bѬ8/R�q��u����r�vA�k�Z�Xw-��V�g^�z�	���Y�:�U�Kw4Eڔ�ȝ.�WC��t�O�u���]�SjL�� ��wA�,�(=j���TUk�Uq(z��eZ̦+.�wBq˔�<��-��|ڨ�.=�1VisUU��^��wG4v)��	e:��*eh�NZ��x�k6��z�t�A�K�ݕ~AZXo&x���:�}rZ����D�YqXY'9��VN���q�#%չ[��Ϙ�3��u��c��;�BHS��_v̸�2\�sv���f�%���Ǘw�r�7�uD6��a�h��(=���5@Z�"C,Sh5�~yf6ڕ(���X�̴�,`��:zxxxxW�l��WM3�͸�1N8��L�ͣ*�T�e��;hn�m\1ˍAar�r��u���5���ӧ��D��R�Wn1L���kU11C-6�wk[�Jܣ�%���[h��}����WU�-¢��e��QĮ5y���S���Ç��É�^7��ZS��k���Tq��5�hմ�-����gZ!�Q�f8]��Z�ܲ����GZ��N�<8xFҨ�2�TkD˚�w.%��W.++Q�G*˔m��Y���~�-]9��U�K��������:p����kg�dq���Y�Tˉ��H��r��V�\k&$ܯ)DX*jq¥c�yI�v�me1�s)k�
ƥ<<<<<<�|�73 ��ʕ�u��Lݙ��h���2�E����h[M�¨�k<<<<8y�'�9Q�����6�.n�1Q���gq�Ab��Q�Ʋ���(T����h�L���N��zxy
ĥ�*(�ʈ�T*2��5�(��RڌcP���˖�p*��}�5H�/-�LW2��32���`4i�U����%n���M��l��e���]�0��4����+=�4�_E9���95�rvv����j��}rm3[�Ɏ�s8�m<9\�����k�g�
ל6��u�O�|��������"0EE��N&�1r����T,��FD�*\����]d�ƾք���B{"�1�PX#��B.&��Fo^���u�/�Ӟ7���60�Ñ�>��4�S!�h.�|����HC�lߺ��o����0?�������n�p��G���Y�f��!�F#.��re��R�������}ך�70Ƈ}Z�"����S����}=�b/��7t�D�#"3+'��42�u���^�����%ǒ`w����Czݶ|�\'�:�F,���	P�GMH�P�i��W~�UQ_���j����(F���3}�S�T6yd�<�!���a��Eܮ�Kٺ<S�LH�{��%�r!��%"��0��ϻ\�.�ki�b��ɶ����|yH=���!��aD� 3$���Ȝ1����l�}���8uAG�uu�2��C�]F�=����/��fΣN�f}�4���yk��O��g����C<$�ј�ߥY���kvt��Ց艮��c޹p#5�魀����ԥV�;`��$vƲ����3G�����y�7�e}���7�|�E؊f���v͈V�3���XY�\+���7:�ww�
z�p�/�P��.�ۖ�KvT�shJ���� t���,G{����G��uWd�E��Up=��R��A���zy�/s_z�������$E"0cIO��|�Ͼ�{���_ݯ��~V7�-��>y>�B���-¢�9 B@W����e���wM,J�!�~��ʐ��Y[b4׻�ń��6,w�0W����cv�����j�6foۛ�i���+>��D����⤦p	7����G��blwRF-�F�<�F��wl�'�oøx�0���R���	��|���(�3��U\�T�Y�R!�kS�t��4s|��cv�mn�6�FC�"�%B(�\;��do�ag���>�U���׏��0G���esj�ٞ������:8�,2���j�����������@Ľ�m��i�~�!��>ng�ח�g��4������=�E�S��R�z	��W��@{na��mAJ�EՓ��_�8
�vg��X���=�}�"; ���8迏K��&Y|V�����}Y �#K�и�s��|�J��c�c�|	g��ψډ����N���^�"����	������L�A����9�`P���}%���H@q���~��g@��>k��g�+�n�X���le��)Mٌ���o9܅�g�V�SCs�=�&�*��ǵ�U������0�Fh�� h�L�>�\�}�f��ޕ�MA�S���>������[��@�hu���|�Upzee7vB(�pƤ�����Y�?<r���mm\۹�����D�@�Y��mW� �S��o������#ߗU���C?��\t��}�Jȣ�d�̾��[ɷ�<��[Ƣ�H�l��ʅ>W0(3$��I� ���/�����'�E�E���������R�:�_X�ii�;P/U_T��H�Vt�ʒ��R�xu���$[��n����l�W_H�U��+��4��F%T��NR99��`��Jz7;�}u�x_��^��B���`!�D ��LB������J�`�{���"\6{9z��&�KxE��u���A��]�E	����S���G��v�$e���oKkF�VM��#%�T�B���P��&��ƒc��г�5>VE:v~��� �:�s�>Lz�L;���o2�}C��G���z3/��J�]q�W����·����s�{����NDgd1���^�=���q|x7����6�/�~��5B������}T��%��͉'&������f��v�~�{��jt�!��f�7KH7�@���k�S"P���k���I|U�ǚP���(G�T�un�/h�2�#�,��ʩQfSO��m,�/ �d�Y��9�kU�9(N�xs���5pd����郝1R�p���Z�(�*�C����Z�������-��L�J�7>`���~O��1DEP|>w��&ٽ�P	'çb��f����}[u�r��Hh�Jų�׬o�7z\�}��qN��<-}�_Z�L�P;,���EqBd4+]���]y�qʄ�/�\�BV�1~X8o�.�\J�����r������CgrAh՟u:be�;?:���gk흜��|��G3���;	�p/��|E�ʖvHS�8)�ro�<!�dy���Ѝ��8^A�U�LT�ba��X��C����x-�h�G!Y+du�ϔ�*"q��a���H��זD����5yϷ+}"�(�~�����_�]*6�8�F'*�Ԥ�["�V�=oz▷4m��{�5x��� �lWӢz*L����x/�t`�]c0jv��9�sa;���9�S���-shW]��~ ��X�Ѐ��:"_���;h`�x+��]O�|��r��D�a��1�i��(��TG3p�Ё���|y��#O��4Nb�},�b�P�!���|v �b�����S����s�AuBX��(��:93�}�ʚ㸪#�M~�z�u�u/��k�)�:���۝����)X:�8�ݽ۳�C�2h���#��J(ɪ9��l�Ӄ�Źm|��e%��%p��új �\UZ���h�#V�U�v���XPRq��۾:z�G|� �gp���o�o�?O�Yc�׷����Ͽ��������������r�����0r�)��:�h��@��A�}�T��:�TZ���}���[^.��v7l��@1]Ґ<���+�ϼX��',�W�U
_�n]��o���z�
�6}�n��f�ߍ��3��U:�����ņ�I3ӌ�a;�-M/t_�AYU�׹�S�3�A��'�P�m��67ӑC[wc�Ku�|f�J?o��/�Ѽb�I����;�V:����� �)&,!e�^���R� ��7�hS�M��l>������8f��c��^�����a)��xe��.���z��$4��;�Oc�k�'!ᥦK��\r�ֻ��Ѥ>SHN�\<���}y���t\j,�PRb0x:���l�I�(�>K��]�P�A�����Ᲊ�_|��m�q���-�\�hg�S�9��[3�v�woB'��L�L��}6�#�rsBoW���2�1�)o��@迒�"n�}��++��ܣ�����d���`@�xJ��S�6��)�:��*��)c�T�r:#﶑��'�� C'�I���#}9�e]�^�ImcQ�̠w�Mq�H��d�ܯ��x�z|8k�&WL�ب��h`�{O���y,J�m���]�tn�xU�k��u�IG%��&����wd
]��m�`3t��}eK��9�<�̿>|�|������((����|�k�s2P��c��I�=P' H`�$�#������V4�ң��q�����c�p�2.K��)�\x���	;��9�Ǥm�0�ȝ/�]
<��M���<UY33���rE�]����Q��W3Y���O��G�g��H�
�O�F��E���.s�����^�^�q�_+�������'������W�����&;L�/(̈́Z��wѹx?*��,����g�M@S=���3�p,r���tj=�E�p@?}61��)�S��]��wt���>��"A�|_���V)�`�/!�s:�c#���* �ٍ��Z�d5e�9�D�#�xa�2S&*-��ݯ�{��'�R0��>����v�����n�1,P���~�k� �-?W퀜P���솭�������麘��7�����<�K_��~�T��C�D8n�К��z���?ӓI�� ��j�Q
n��3�>�;*�9{y�]�X�u�y-�L�`�,E<���y{�S�E�7%^Ƀ�#/<���~��1!2,7|w*�n���tP�6e�5FtΨ��7�mZ�,���cuJ�賱�Qf��5a�,*=��,u�gpq-K�z���ҹ���MGCx��̔l5�fu�e�����c A�ubs:r�X�����U{���G*7z� �
����(
QE#"�s�{��|������&t�=�~��%��zX��K�a�\_}'���N��mr�b|P�U�{k��l����=i���Y��P�c�J:8��L�/V��#/��ʩ=�[6���
^�|/�����8�����Bo��ާn�7�L6(m�o`�Lǰ��nŚ�V1i���=�}�懇,�b��~��m���>�7�î���;��~������7�"4��~`��_I���qށo�'��,NU^�9��]U�$��
�TY���^,��f�)�T��ɤ;�h!��~��{�!�eR/{_e!��_�i��%��E�N�@��WC��{��خ6A�_�D�^���x�7*���|�ć1l@9A�����u�v1�SKH����_�g`5�+c�7�����=���x��I�.D��(��f����euw���6k��>�dE͗����y�8�9��XϘ�U�<mzP�����I�u����G�7��6^�g;�����tFc۰Cܺ}ǉ��B��r�B����:�)�WVsH�Q�F
�1��ݻ�B��F��S#*��V��w�5Cw_Ǟ�B����,mQ��n�_p�﨏Ňݦ�"���D��d�켫N�����c����y�|?�@ �H�{��bbK�?��1O)��~�V:FAG�I��<�I�r� ��5�^�}eW�Y���2���,.���B�K�r(n��5�l�q���`����K���i>�����6��3�������+������"�
���Y��W8��a���f~���$?@z�9�|r�E+�2+R���! 1�m���9&���7s�YMu�U.��&��(PȜ
\T�<k�}`���C��|���cV-�|�ғ@�8Y�OعA7;���>����1q�c<
�Z;bdy
���s�ĸ��R�ݘ��Fg���ofFi$��o���Xӱ�>�x�\}g	�d8hI��!	؈��dz��1��5OdO���>��#5����j� ��g>ʖo� HDe�2�=2Vc�FRuc�$�e��ow[�Dmz$y��]����.'t�~:n���u�^*"0A��A{�-��sN�w�/r��:%FX������b�-�$P^u�o��=��P����3���<)t�2��[�ٵi�y!����ۻ��7��5ZwY�rp"֒ElT�Pc��z1m�$�����T8b4Ȭ����#�*�Fv���w�GSh��&�Ȫ�^�M��5�2=���]�C�C�uJZ�i��&w6�U%02saL����ȂA �H��#�ܦI���}~��v**tN����GBπ�����k���E}�v�N�q����U��ٛ�Fh�2 � މ��u���Aa�3~۱p�uu���O�~=L���u^7���7�k�q}X�R��셳zA���]� h���M�.寧��G���wu~aw�u�9��ܯ��r�� ��T
=5�P��'���GNyL�(圿}���T�O^���ǡ,#��=B#�w���F~��7�X���o���"�	1:d�@�M�)�c�:��l��s��?- ��U?o�观=Td��7������R=1���_VQ\�:b��f1:�ls�wD
j�hҡ�=	�o��B{��&��_��-�RBq��=��9�\�Yk:_���S5@�`�a��� �Gs�����r+[w��#�s��M8Y�n�U�q;;�)L�����6�����]BɜdNѡ94 As��5�lk�S�c��4��j�8=�z�Q?M3i��+���I�b�K����9�P�1!�
'����=�
�y�m\I���|m�K� ����_o�muT��b��}��v���j��tyl���J��A��Q��R��O��Z+�o���U{�ǡ;\zp.N�U�Z	������f�R>���3�R�\k9mb�1	��d���"^�:g���/ofXF# �`�"A>�����M99%�;�Q��A�a)�l�j�Sv.��>��Y��P�� ��=P&gB��M����w�S��m��;Ҹ��=N8�3��pȶ�8�d�:z�r���i��6!�5/~I��vjOW�*���+��:Խ^�C�V�"�qr5��n�> 2�<������j3o��\b����qZ��.f�9xE8O��B\r$Gxo�,U��S1�}��8�7��x�*��.��yp%��~f����z���C���L�ׇ! i�_%@m.�����[݈s�6���޽��ٹ]ƞ��Óa9�6�"B2L�9�=#j|jK�S"t�:M(��a��ލ�C#n}Y�<��ub߅�"�e��M�K�+�� �U����W��h�^k�z�a�.����c|���|+a�C�3�>�R��z,�f�v��,����xҹ!�c�}*J�F��>���Q�4 �6F������7�#�T.�3�����������o�!�3F�paD��	��7lF��y\�����)1о,� D���3���Z��y������bY�3�D��:k{V�^�l�I�;s4�ȦL��A;T���+�XDLꡎI]�fs�r� _k�/zk
QلjNPfR_Q�ۻ���F�<z���W�9b����5���]ی$V��N��u�G��_�I�/�ɲ�J-d]V��$�t+�@Z��2�oN&ʤ&j3����K��v��h䝒�s�t��(��'!�������1��[��vt|6��g�6(.�������`���M1f�bH+�4K���I��N�!WE^Ř�kg��YS5��3P(8�l���]0���o5.v#�ȔgM��6l��oqfٛ����ʸ�mDS�g�$�!|K���M"�Vy!m��>�³���P��C�WT���p��(ς��=M�9辄�[�n��k��Z�l6��bK2h�9��L(�j����ՙ�oy�U,��NP��\�L:=
�O9�kNl��˼���2�=O��Q6����]�q�\B�Z \#hR��łD�nn\g�9�Ԩ�<��H�է���70Z�z\ݛ��E��7��,]�� lU��� 3�+�<�z�u�w����M��z6>�BDCT�i�Κ���u9a*;(fY�c��W�o�촂��1�B�k-�{��D�Z���[�̽s��b�w�X��D��Z:��y���b7v�^��3�'T"���i"JT�T��LP�T~�8YI5��]���W�U)�nJ�p�=6ᮐj�pfq��׼j|� �߫z��,b�R�����	�bxPc^I&%Jh7����3%���G(*�}G3%�{c�)Y��#�U���	E�GB���;�-�����}��i�����󨠕@�>��(����Dh'l)�놷Ǣ;&C�f��جc���f�\ēu2�=W]��;�G?�F�yJ2�5v�-�I�Tf3Z��G+����ə1s�}a���T�Oi��
�.�',2^7�t��T���e�^b�qLV�ntff�m+,枅�e�����w�R8|���X�;�UIz�/1_Vz�����k\����`�U��M�D�f�יt���i(�ݫ1i��2��m9CfE�1o�*Ԩ��%����#P�/*Q3����LbF�A������.����!��".�5�!���RY%2B�������Z+x�Zq��; �s l31�����k2�d���&���}.v�n��6y�˅�@�M��ۥ�Q���ܶ"s[���Ĳ�S[��&]-X��9�V"�eԿ��i���9�z�&�\�[qu9�f��2�����f����0~��]y[L5&(sj�̴{U�b[b��;���cרG
yu�N�+����]y;o�tV�����u��P-Ii�) S���UHv0,��]jg3U&�M�h�I	bFH3�H-TD����)�f�BWJ��W��Ei��cI��g:9�bc\��)��T�����\�cF���r��nUƳ㋻���i��[A�?N�p���fa��!�/��lʱ��U��jZ�y�֞�)����j�nn��ӧOm�)��SiSZ��ambT��B�U�����T�&M���������X&%�`�5�X��U2xxxxxxeTQ�6f_�L,����[kR��5
�B��Զ��k4U�Z�[�]�=��AF2�HӇO"�і�Q�\���Ę�R�V6�P���\|a�Լ������OS\DAM=:xxxx1�(S�U�,Y�/��Z��ڊ�5�J%(�(�{B���6�4�������)Z"/�Ɗ9_.Vʩ(���xفP����a���)��A�Ti�*�0�N�<<<��r�AD����\LQ
0�1���\M�5
Ŗ�Z��-K��9�mMj:p��Ç�aT�4([ieEg��VPb!m�Le��F�E���b�a���cceTV6�2��h3g���b��KA��0ʈ�"r��~���e�>���f�"�Z{��s�7��w.�}�q9j�c�R�9;�Z��FA��T�-b�X6wN��%���v,��TPN�w��A""D`�bx�k�pLE��?��B��>��:�,1��?MJf��c+v~�{:ȉ��鋋�$v]�t��
OhǲB�*�Q�_,�-?V�J�����?���U_����V����7�\&�C͞�E�R�(��Sa5B+=W��,�q�d`S$`-�p�h�{���r���X�6T*����,oKgc>���"��M^�G��$�7%i#�͙�p/7r�}�	�CC����x�s�ƃ��2J��J~p�?+�b��ܟE�<E�
���J�UJR_�r�����P˩l�o�p��8�>��B�)�-�&�?{x�wJݧs�\`���M�oӑ*���}"�"�z,"�"���&8G���DwS���y�dW^����ƻbj�Ȼ�H��r�g���9�`W��>�ږ�ʑ��x�������C/&��)?>�?}�@�D$���~��|�q��'8��hm��|l`Di��������!��Y �����,5���[��]E������|j/Sgr�_ϰ,�̒$v��D��^D(Yon}�~�}�ϵ�JnT5�O!�,�x�o�q��^*�k�yN�a���u�r��S��z�vQ��
#I�{c{r���^��@t �����n�� �cl]H���<�� �����N{2���{�
�|��~y�s2���y�3��	�DH�""�AA��׿�����9��?�267F�����W��ZFbN���g��`W��ltQ�X�~S �x���ϵ�~���E9"�?p�;7=C4���.��NR9Nlq�"�G�J[����>�x=��	��ȁ��!��#�����]�{���g���O1�t�Q����D[�xX�.����X+��	\>a=�	�����s>����*�V��>���\v�]�y�L���E����P��M��H�(��h�4)B<=G���g�B2�g�f/UN;�N�2����z�ف{vBGێʃ�0?�	��x{͜���N�=C%|<��Q�W�j+�K*�c��v�g�~0|QOib�Ḽ���t��}�_)�rߚW����.0uNI�U�C�W��yx��=.`�7#��A̚�TD������`�����LE���ð���V>"��e^Á��\�7��8&���7~�#"F�_�`9��a�
ۨ܅8�|��AnR�ɳt2�WO����5��翖��L�P�(�t���x{�a��sc�t�~��uн'���$��BC�F��=��u�ݏ$�^�]py[��,X]�c!�[ٛ��:�-��/-�g<�϶L�.����jC�Ӓ����z�����9c-��w\��yg>޷��o�o)���ḝ0D7b'D����2��J��Ԫ�t�:��=��?����TA��#��v�����1V��������x�w��m�1AZ�_FE�&h�,��T�Ͻ��]��J����50Ɗ�W�5T�~Fj/�CO�@�?V��2���#R0�BЅ-�6f+��;{rV@�E�~����.JF�Z50.�/��6\���"��߁"4�w�ORf6�nS��AJ0a��T;�
���u�k���8u�yg�NT+�#�w��^|���ma�n�z��А��a��?s�n=�;$�*��t����;To�v�s��R%�mo�Ǻ"P�,b�C����@�������y�/�ݘ2j���.Z�a��ʝI����^�N�E��H��"B��f�!n����0�y(���Qx7�|$y_L�~���42�^G�ޭ��gڕ}Zo��R�b�(��DA���X)��΁�R&�����m�vF�x?,KY��}�����*�Z��a��]`4^����+'焖�D9��G���C�@�A�}��*��oE8�P1��)�Z��(�<<~�y��@��Ơ*R��,��|h䣾�;^Wkkv1|��;g�滻�;�u^Zw
~�N�BC�_/Y��f�(oz��*��_M��=��J���pw���r�!��[d�bWj���ݼS$=m�;��#^���Ü�X���r����"	��F��my{X��O��&�Ή�����o�ݿ��α6;�@V�Xc*���m���}�.���-̐��x�������)�~0���+�.�~b�~���qͺ��ybgoNe�]z����LB|�E���P�kll�:<r�M�#$�`-�鿥�GF���]ދ�?F�K��tў?��+cܥ�p��,&�b�ܝ�b�Z~VI������]K~5�*j{���1���uth=,2,%5�	��v���8No7��Ȫ�ov�ĉC �	�
�>�xw��K��)�e�"��n���FO΅v��
�(ˋ��[�ԕ��E�N�(I��L��)"�u�l�L�O#�j6q�1����ћ�8��ce��1�+I�}?9PB~�(K���8��'�ϣ3���������Ra���?p�-��#�8���6�U���!t!�������G�[9��_n�ʽ�rdߌ���~T�o^��5WR��Mp��'>�3�D�d�Ә���H��BK�Q��,ݛpn7*�q�t���]:u�:��eL���#$����f9�k �{��P�xK *�3]���@����{҇=��U�6�ժ�t�4�sM)N��UO���R�c��8�Y{sv�,vy��Ԓ"�v*��̀ޡ7��*	�Lշ_���Ҡ��Y��?DB""DH�Q��/WO%����1� c�s�"�:��f}�M���W3T��uC��b=@��Z,�q��p�X0�e���ݓ�l��X�LiH�t{s�Z�=R3���JO�A�i��P_��h���ؙCƇ�>[=�v�D�ПIPd�w����hz�~�G��4	���	6�g3��\��_���[�r1>E�j&�	��@�^�*C���c͊�+�}�<�b�2[{U����y���/�a����_h*�r��?t��^|T��	7������\�-�T֍'�=��bw�3�Y�n�ҙ����fR��T��d�ƽ���ʏ{�~K�}\����s	�	���dG�@O�E�mwa}1`T.]�*p�[��s��[����uY:ȟM��/�tK�}�o���\�u�گOh�����{�"�?�u��I.qcW>}Q�<��T�bۥt3�Ul�s�u 
6WW��.{VU�5qc�_�-	�7��jm����>�~�U�a�u�̍e���r��:=&��3�E�މuz7�Ky�X.G��H�Ph��o�~ì�s��;VzX͊��:�����X7(G�;��n>[2��NI���ӣ=n����HͶ�A�a���y�e�ܜpԹ����dF"����E�}���߾�c���P���?��P�`��{(9��A`>��׉��-�����G�gc\��ow��	��Zk�w�T=�!�|P�f�c1�=sX�Rj_��qY)ꗼ�[��v�WP��R�~�Rrt���7�w_e`��K�6{�:Ay�꿱cw���[ćA�ތ���J�ݲ��v��"�/a�o���C�V��v;�;������Af�;4)?n1W����x{�%����X�R�z���[��z�]�lr��2�'Ca��������DA���t5 �=�hp��<�y}Ά���Y�fVf�O��/w��;����[��ұ�#�
<�g��!�7�ǌ:uZ���i��[�db�5<��B��Fw��
���$0��3�
�foi^pˣ~�,[����k^���D���	qK��i�������=�k�m�f`l��Բ]%r�r7�AJ-�v�z������5�a�G�x�B��쉓�Gl0e��/&!2�9t��h�X���� �7d�}j��ٽX,��,m���zTBq��ү+�=ңoY�{1p�$"�,�É�k���Y��2���9��
�U����@��n��y���x{"�߀�����{ˁ�|���C-��۸�g?U `|3�R�<�����%��^�9��2��U=__�]y��}�y0����>-��[��IR�h�OB��ʳ�1|,�Js��}=]�[�'�>aވ��ˉ���_�k�,�^?��MJ�-���*���Y!���)	��<����*q�4w�7���D����{��ΜKN��2���wxH�:��߂�/x�u��NkV��E$��9Y��[|����|�
	��Wі_{�/&	��}�4�~�P'8 >��`��a�7��o����J�o��KN;�~��1�ڽn)�xh?�ީյ��q�/3+Mj��>N�Q��fd�7Fnoq�vʩck&��Q�Z����	߫���C�ς���3�nb��#�" 'N�z�Z���J��W ���zAx�<T�Vɹ�	��pW���l�S���&��</|�vv�euC���:u��/Y6QyꬋjS��kfH7��[��d��9{Ϩ%���\��]m��#w��wv�n�{�[6�ƅ����j���+̞�'�l�~�kZ`��;�u��>� �:�O9K�V���ϓK&^*��i�m(r�BF�S۸�U�u�w�v�i���/��x�+�D��螟_�;�J,J#�ːO�C
��G���:�>*;����Sƽ�z���vM��{��P6-���dfvb����U�6�e����^n������C�!\�.��ƣV���0�������6G6͞f/�?p�����V{E��$fN��)�k;�t\�@ݎ�h���=�ȹ�G�r�4K�����3m_�]]{�Qs"���Vd��ǳ�'lV����5���v��Y?`jNezSG]LuY�\H퍜W���Q�_O���ny�"��w�����*ʰë:k�:��ɪϫϯֵo�S�N��7��F�ߒ��&���V����%?�xA�ďw��׽������u�o�)mu�Վ2�N�|�^�Ϥx�g�N���ܜ�N���y��$�\�.e!U�z�W:���ge���k�֠&:�y
��b
��E�����C������&}�gr0�{�J�c�!ʙJ��)�'�(����G+j`�n��cA��n�_�f9�r3���Ĺ6��~�}����;H1����@��#�V������_�p��r9�j3��M�>P�{w�gOzz/<��p'.���aR���1���û��?u���˅|"t����92���O}z�CC��utﻣ���(oP�/K�[�ʸ��]�F]wr�T�B�ʰ���iP��1�1����-��I�y�wvW�'mNՎ����n�������רQ�O�o���WL�c���>�Y&���]�A�x1@��Ǳڰ:yu������ĭ��=�&��y5�{{b�!l_��8wH<7\܇���g7֎ӾQ�����b�f,��Z�PV1 tƎ���.���m����S����
�B�v�w����$�z��E�G~\/huL��΂��5o�W�}*��~1���|i5[~�1?�]���A�%w��v8�9*�@��C��~�Ue}<�����v��c
<������Y�8̱��z�ow=(��!.�ZqfS��&gt�]�pi�A)������Q�P�Д�黓v��+2}6�6�'B�G�
p�I�p�{s�T��nD�Y���n���&�.����j��M��eB~�_{���"k���v�~c��\ݰ�^Ws�����"���)y�f���ͷʢG�f n��Vr>5�R~����,~�{��?{�8!^՟x��x#x��k����eg��	~�H~z}����!b��Ԡq�	���#;1o9/m^7Vj���9Y_Kbw8n=����Sj׼�f��H�~�=��+C}ʁ\��c�Y~�z~����(9�	#�LU��Lg�s��EG�������t�*���g�C�H���%��צꯗ�E҆�)�$�t��.�-1v��Oܼl�oT�J5��w�]]��*}�a�Mj���y������^��z@�u��뗟MV�}�/ilD����R���)8����(@��u���R�^�_s���������y�w�ҋ����0���dx{X��yq�=�n�,G!ϼ0 �����a��{_�sW���j=���]�	Pp�c7�A����[9^Zü�ur٭Ӑ�uٚ�ݷ�%I.����Q�:�f�aH�X*��qIH�8�ɜP�;�_���n6�qqފ��Q�'F1�%�s}���![��S�ՉV)���y�w�� ��n�h��w<r�]wY����)m�Q*s��!}]�s�Q�����k����B���'Iɔ1�p���cxu�a�t7���yҘ����åR����Ft���QΕ7����4M'O;bָ2q�KM�f�]�Z�Ë]���'oKp�96=!e�D��*���V�Lt��Y0�Л��^��v5�Dns2�Đ3��Xpq"����"��N4��{��[�JދS�{Vή%�����}G-c�q�]\`c�5,܉}K̑��r��\���C�Y�q��Y�]������V&�Eݘ��k��oh�6^[ro�.����t^{���9v�-�6�]�;nc�۪�r��T�3�.>�A#8�����ve������Wv̙�t��&�T��T
�n�S�9/�J+.J�V0j���&u����孌!\�KR�3��Q�����~���ekwÒEc�: 2'-!��o-U����(�Y4aN��n���	S�Yh��f����ڡ����j�!j;ce}�bʼ�2�j�C%۠���H���뺗q��˄:����Й%�;3�E*A�!lL��}WZ+r4������f�#-
�.�nd�b��g'�"����.IG�����gu��P�2�������K}�9�]|�:�O+E�1=����;V��]��Xo� o��{����dunkb<�M�5_��KI�J�ﻄǜMR��5M�WMI�1pN�pr��嫷[�CV9�{����]�k�2���q���G��uB��k!
�6=gI�K(/�ng�w�fU���y�N�c	1Tإ��X�2'�K�[ ꝺLo�n����_�T�--���ۂ������+;M���Z�9�Q׋2��=����m�_fP{�.n�Y�m���O�2w������7�F����zo:o__+�o��h��<ۭVN�x��p��6��Q����:��]��-�/Y�y�@9�����kt�B���WW��y��/�,L��V�Ƶ=בb��*k�CoEkHMY3����˲�ls1�˞�Ẏ%v����#!��R+w*;�9��(�۱Z��f"�}����Y����%�O3ڕ���(�3بj#�|�g*�\{1#�Y�O����דF�y�'�6��]���7��Q��;���i�%n���8e���ؠ�ݬʐ1���v%ӫl;,SS^Uku��it�<Z��SB����s�%��tů��-<�OgL��dL�m�-�f�׊mfn��P��kX���mTNڕ�R�&aUU"*1�U�z�5P����b#��t�<<8x*Ŵ��cr�����%j�*�=f�2���̱��9�b����&5��c�*1xt����J�S�҉Z��Eq��Ţ��fep�*�\Ţ�\��eYpr�"4�������R�KXƖ64��K�E1�q���j��Q���jyn5*�<<8xx6�Uq���W-S�3-�f�b�#���B�jR֛��"�J8���ˎ.xxi��DEOB	}l]h�Y`�-J�~[T�������E�3*R�?d��+N><��髒�֢���R�6ҥEjQ�Sn"�3*;$h�3qk�j�F�:t���X�#���Qqr�
ƣ�&�"j��T-�s0k�EDci3*�

"(�\����Ç�m�߉�T�QERZX"�m10c�inR�n��F�Ҫ���\�	iE����8�TUE)j�F�ʣmQZ����*�*e(��1�D�P�	�M�<�@ac�y�����365�UJ�nvf���T�]QL^�scF,$:LY.q����+)�ᭆ��"rӱ��o�;�Y<=�Z�}�
��#��u��#~ࣆ�����|�H=�H~5�Zo�kټ�~+1���d�oo��լ�x5&}���Uu���N�U/j�찯�Y`vo;J�r���}Ɂ��ކ�~#_��{����S�xz��|�HrsV=�ku�kPԼ��
��\���4�[�V?�v�xR���a�~�͏��!W�*ry�^�|/���Z��q���wW�|&cNk��S�/2���=�2z��>��m�6��
d�X����$�@����}�g�m!x��'{��o�2���a)<�-{o��NM]q""�L�^�j��/Fy杌j��K+巓��
� ��~~��l$:-ŧ~���\���{T�������gF�j���ܴ�̏f^�9�M'P������p���7{�\��w�~��.]/���wotZ�\��6`����7�2��Z�ZU{�0���;�IN܍Q��};Mʻ��_Ƞ�}�������K��.�VE�
�_I�n����
4	2d�q={+0(�5p7C�g'��T�o4�Q�6M��K�N{4N4ҫN>C3H��ӈ�X�7�q�h�����f�b���}����]�
��ǃ���,��c3�\�:i����~��6=�91t��GN�f�g�}���F��'�WyS^e[���a��Tp����+7=G�	�D��c<������0/���g�S��wܿ,˟��|Z-�^O�Ͷ���� �mc�
��z�� ��O��eQ�w�!z��^o!����;��}i�sb�ꜯ[;Ch@(qU���Տ.=P(ž�^^�z��o֬������v�C�����T'�B6G�:*=9�£�6�o�U0�>�~=}a�����7=��I�{3�-�2{�������O�<ԓo�X����)�A9�x�N7_{����ﻨ$9B'�.���h�w��Y+�H[�6]�	�����6�o)|7���&j�����-���-����g��}�w�}yn�͕C��4+��1�ﱩ][4�eQ-���̂0e�ݲ�j���MQfSI�B��#]r�:Y�h͚xP�A`ՠ�}��"����W��������q������Ӿ��2b%R�״����g�e^*!�P��s��oN�u�ʹ��K^�lE�|�k�c;�Aq:H��(|?
�m���yJ֍�g�1}�ԕ�|��{m�x6�����a��ǃL���DML��7vC�����ӓ��1#���LS��>ǿ��*�DbQ�P�{���j�%�-�ѫ���ڍs	�-���2��{0�����ݭ�g�auv�h��~��ٖ��p�����kj�J�N�^w�;�9�������9���+�$,�ؓ�9�ƽ�}�M�gm���=�K�M]�/�ԫ��|�,�>���� ��ڞ#rSk=���G����&�=��}�~*k������{/�}]�������Cy]�P����Y�^}�lf�����U ��д�������7#}�>Ò`灭�h��3ݾ�g�"��wF���;9��6;��ouL��.�[p6�e���۫����%��@CT�G&w=j���6�.��T4�(Z��Ũ�Qᝄ���^�=<z�Eq=+��%�}���l�Q���'=0b��Ͷ����G�z�_Q�oi
�_��-�{��5v!�&��,����u1��3r�.n��jsh=��%��
��e�!�'w�����0�s=��ݱ��Ů7�܄xd�WB��=�|�R[����>���XGi�����N��o�45��d��[k�D���Aw�<��\�qfh�?*����:gk�줣^�H�E��>�a��e���>���a�K9g\�v_��c���m�i	{
p��="��|�Wb�تr/aV�v��Se��Y8=�����&�Ǥ���e:ׅ·뽘��DI����Z��0�����z.��Vw_���߬g �c��m;�@u6" Ń�K��<.�@��.h��O��+��<�.���I��ED����^1�@�Z�'�0>��^ȴ=τ}�����q�8N�m�g�����+]'z��i�@׋�5�Y�.�{�CleJ|��Y�ڂ��~��1�w]��@K��:�|���ڋ���a,�v��H��tw�:7n4+�N�t�L����sE�:�ݺΧ�g~:��)�����z*�tTЏ�����{��X��[x�H�4d�"ە�n����+8�^�gNvY=�*7�Z�£B����e1����*v��J��m�fޱ_��]B�S����!c��g�S�J�I���MC�zF�ݵ;;��I��e�}���'�<��ɉ}#�W_������j۴���Phz}��l��]��b�Ӱ�aX��~*D\og�L�p:�W����|���Y���g��JQ����OΠn@�=� o����}ڭ��]�d̺���v����z����n�Jܾж��Go��GACzH��?TRʅ�+�0i/jB����ׁ�g�~��O�o�<�R�)��pPG�[�c��.E�<�o�s��Hퟳ$FW�s���(Y�OxOf�^�
w\�_Tȷ�<�Uoyzҭ�+d|v�}7��tl�=�`���
��H�P+{����4_�<�������F̎�[��3{wy+	z v:��ݰx=�+28��Υ�X������\;w�h�كat���2��OP�P_y��D}�n���}��5���XU�];*19ᮼ�z���j޳����4�S&!ns'�2]9��p����dW+�k��[f�`�p~�ζ����MC��ec����F����V�D�:�EJ�\q�K�(3�U� �ǓN���k*�掉�i�� �G��$�J�C}�o�;�"�{U�+��"�ROP�ߣſC^0��N]��6g�f�e�Pm��H[����z�z���9B�R1�����yvmX�|�_����l�m�m�q��!�hWü��w�5S�ɫӻ�0�>�"� �I�뷷K;۽�D��փ�)H�č�DP�M�e�iW.N�_2]��T6�d�{ynw���eOy�Ԏ�V��ϼ*}�����{�����Bc覭�Iua�?_y�!Ƕ<P�c�����R��g�g�T_�������1��c�7��R�["��~��b�Ww8���yM^���ٝ���/�oK1�5�}�1�u�Bؿ��?@ޒ�mwP��f��r�q�{<�������}����7�2:����f��!Дn]_�yO������l
�ޤ��q���:�^��,���|�=�4�3�9ZtV��l��=���f�k(��Xmo�.��mυf�n-%�T�ς)�$
���P]�1�Sr�\c���Es�����۠�%۹�5Wxg
�I�Z *�+;���Pi��t:�9��n�����Gq�S��|��O5>_��#i�� ��m��F�A����/4y��_G�t��*O���5܏U}��ӽ����UI<;=�$��J�Q��s�֊_����� ���>r��ٰ�7��l�� ��������!��zf+��@�/�m��R���5�2���^�s�f�wD�/|�����5t�fʯT���E�SP�|giǫ�{�^>��c7%��_1��䵱_{m�C�����I�|�K���>��wn`��R��k���S�I�@<�C�y���0g�!�h]x�[���D�������Pծ�=�z�6���ҥ���{7�̚�[����v|��#�ʖ�_o��y��*!�}�o�2�E�Ѓ�x�'9C�W�bn��cR�g�{%e�CQ�B���$�~��C�<�A�d%���bƿ?#խ�R����Ȧ�r�!�w�6#+�� ��XcG [�ϩR7��vk�""p
�%C���72�U}¤��^�H�}�׫v=x��OR��b���ǫ�m�z�v�XM���|�W&$�1�U�;�g��3W�����I�����Д���AvzJ���[�n�F:Tİ�r�l�t?}�諏dn{b����iҗ�,_/i�=���aa��&� ��{��OP+I��[�V<��=����9���h���}Ͻ�u=���cH���W�y��
x��t{�{��ӯ�����n���6)9
�����5�_�G~W����@@L@�9��Nnz�>����;/HK��nt,��1�1�5v+��r;�@@�������?n/P�o�ۚw��+b�Z�b��w_Ͻ>r{�mWX�=0v�tH�f�<�t+؅h>�-���2X ��+}�������\���Zꅃ��3��-^N�ɋr�z�׻�w;1��3اH�K�t_,�j��Hx����o/ ��>}�v%u#܆�q���χ��bHu�� [6��Oה�d��ɜ���{�7:g;yz�S���Y0#j�9���X��X��߯��*X�߲Ty����Z2.6ܽ�v��=$�4�	B_s�.�`�X�������	������V!ݻ}�|���z@�r1Bx�?��%�}{D����6̆%0�k��0`��{��x��];6-�ݵg����'�J=��S3o�U���X�ɚ����سz8z+�h��0pYF��zF<j��5b��Ւ�l�F���jؿU�fҿ��Qv�=]Vd
�!���eKbw8#�b++:wLlYer�в'e}}��e�M`ev�B��y�aX�<[�u�Aџ��D�[����wAx�a���R"B�-��6�\�6���������&h�}��Qy����������.�'�YΚ�+��ƪ|����=��F�]w�Bs�2&g��48��Y�bT^��ώ��b��7\��mSz�r^���B���P��U�޼�'[_D~��%�� @�H:��e:�J���C����k_��7ury��$�վ��������rہ�'�'��|����os3��9��/T�!kۤ_.�x ����q/���r���~�Y�������X�+���֕��W��G���=�iX����;9�㺚��|2�5P��DT}i�#��]���O��^�n�S�(H����Wfs�fOf�B.���:�Ÿ1����E`�	&�a��(T�=n�S����X��4k{�	��M�Ԯ�*�.Q(�9��8���f�������7Dt�����]�<�G{��ߦؒ��O�k�
�P�J��)h�_}�o8�7 �g�N�7��"Ʃ3փ϶����w��w{���IpL�s�j�h_�����T�&�.��T��<9��&ۡ5uמ���.�p���=�7���'�P���+'P���Y_�v0�n2�eT�_�Lz'o��9����Эy�>\wA�}��ǓEn
,^�k¥R��|�U�U�Ѷ�_DʬKz�Q�_	���w�;�v1�v,[W�VUy�EE݈�9.}��,^�Z�羧p%�^���w�P�a֩j�sv%�q�p�L�I�yV6P�'�qm{���H�p�烲��T;�����o�r�'7��]��4k�g7m>����D��dm��on�9��(�O3���=�Vсr'ۢ�X'-_��Avu6DY��p���WyWX^fw� }��Y����M}r*�bD:W>:8����֏��� ��֠�pno���B�%y]�Ge��؄�o/���U����4�Ùfa�c��6,LP�9�[܆֨�$�r�sW�qN��[�%���� Z�W�h�Z���]���P�E��Ǉ>���[f�-�=�(sR�m�ʎD̈U�ܻ���1[���M]���Il���:�����"��l�+��V�{ϳCt�p˗�;Wt]�Ԥ+*y�0�BTinZ�����d�ܡ�a����3ѹ������C���G�4���Mq��9�,��ye�u�W���I��M�y�Ef�(kC���38�	����n���N����-x����\�4��gӣLb�����a��6�=���38>������Oѭ��f&�9j��S��:��iF��6��;T���_m�h=��*�Y�Q$���L��;j��ԟ<Od�yc}U�X'��]n�[%^+�0_K0�ڙO����xmMО	�g
X{��p�ͦjK�y��t8GB�L�c��>���=���ɰl7yM��׹��;[F�.�j�6�4�����cBt�.��\#)�q��*B��Bܹ�ޫ�݋�f1�in��Uj�\0�K��m=�3.6nf��w�Z7�nP�k�x8�1D�hr\��Z�l[;��, ��=@5{xb7�l�n7n�& �����3
}Z���{����zĔa�I�p; ���T'"�����`�p^\�EPWJ�B-u���Vc�ՙ}��M����Q�B�9nB�p���ȵȺ��uс�̵]:��r����e^J{fr�xFҨ�:��wi��ܔ�J�Oub&5��UNr�n���v��m��pS3�J�㺐Q������H^M��ELr��<�d^h�u<�ւ�s��Hr��7�#�˵��5�{n����I�j�;�*�\m�\���R��\]�z�vkµ�v:m��ˮ� ͗�Y ��ƾ����h#�eXܼ`�&�Kݺ�Nf��M�#�D�㆑�9ܗ�R�u�;���qI��F��i�i����FƸ�cgM�%*\�Zպ��C���0-âZ�29Sn�m^����V��n��y��� �ѷ7z��t�\3��A����n�����s�t�|�j
6[�Ҕ�.s���9򜒘[�CE�66�h�W�,�a:���-�,q⧿&+�(u&�oUؘ�&2������=)b�!����dCuS3�9B`���[��9bH9r7��b���=qp���U�Qro	�T�2�N��9k���N��o��P~�8�^�?y<��S��y"1�8��Z5�o���H��'�euh*�ij�Sq�y��e��6�a�W�4���Ӗ�Ⳙ}q؂Kk��뽡�X|�E=k>�X��m��*����e��)wnv�ܴ�N:�.�������h�"g�SH�(EhIj�K�"�6FP_��)��� �$�r$@�iQ&R�"eK���
S��Y�9̷9r-4���c�Ո���F������0�mQ�j���k/���N�6�X,�j
�,ʵ�pӇ�xxy"3��+>�Fm�R�����܊�"����B��-�JP�n==8p�m*�[�X�D
�b�bx�-ZՉ��Q�*�Z5+�"ܣZi������fE��,D����Q��?b�N��U�J�Z0]�9ׅ:t��ï�Qc6��D��Q���m�#�Rz�F�ܤQyh�=��N�<=��QEc+����\.S1T�.2ʥ����cZ���V�p������ų�-��ح�J�_̢9w3�b��_r����+QU*����o�p������!��'F�W�r��K�QW�^e�����a�����#�US����Ǌ��m��Th�-Z��V�"���ɷ6�X��k�Բ�X���k�o��J��\��Y�"������W�1X��W����u����6��0u��TRVU��!f���^����Ѻp��y��}vR����N94��d6����?z�\��}�ܶ�""���z�<m*|�5%�����'��)��Bg�����_.Q�l��VjdW���r����:�>��z|����=t=�^yT��Dt��s�k� L��*����ﹾ��ᕂ�U>��v��������3�{��ă}bԟ	eؑ�7�n�^�:��u��|�F-�ݒ���]�)��[���)S��%gqW�{{�|�_���ـuGl����\*�Zc��4�c��olG���=�7��ć�6�]��k��$?�k3�¿/���u9��#ވC�J�``�� �n�򐘞p >٪���Gۻ�(ʛ�4;SV�1_4���u�eP�A:e�x��U;�{Eϯ��ul�NvL��_�쟵6/��J۴�Ƕ���ٍy�s�^��^���ܭwT���ތCՂ���NO� �Ra�+��Av{�ܓ2?J��]&ės¾[���g,ۭha5� X�
�_�u��ٓl�����քZ�J�j��X&kn]�����Ka\TM�	Ά��%��SDe�5��r�Q5C\(@S�9�����W!D`t��F���[\�b6W�3,�׽���r�$)矲�����yR�N�|,O�Ts�T�j\Vď?m���f�9>_Z�_;+��ȑZ!���i���>�m{�نj�/�^�ճ>�˰��v�wgrGe�CT��>-���ƹ��s�;�)����ȯ����!hm$�u��Q��1�
l�je�K��e������wu`c=X� ��#q�\��P�@~�������D���zt����ٱW���xEZ>����sݎxv=��m�}���~F7�@��59#��GW��)��?g�k���Cf˞ќ[�{�lRe'�F��gʳ_�١�@!}F�r��mT����ح�ήQ�����X}7Y�0}��x$,�ۜ���lm�N��@ߡ��k�H~���Y1��矟�+Gvf�ޅ�x���%�;C��|��}�	G�(tσ�������z�Uav:�=���6��b p#b��:}[v,gv>��l�쩃��!�p�3"T`������0�+�@�z�rx�x^G%�)�ҮS3��*�nm�)A�YK^S��2|WS�rv�..����L1Բ�N���y!TU�,��wi�� ���7�k/��x�h���h�-���L��
��0�X�E�e{f�C��-����P5~����3��C��M�+����}Ӆ?<�Q���]�wp[��
���y������z����16:�s
��	��O���w�0z�J�A�����g��8�N.�.�u��7_y��3�Y5W��T�ba���/�,(��S�n��}���R��a���	ROcƎ=ELY�??{�u&���֩��ǵ�&�K�\����up~at�+*Ho�g�2<�EG�g��j�r�Eo�G4҂�&����:�a}�X�=<m�������|�Ի�����5�`�O��k8��c��|�F���s
�!ν����O�?W{��>���r<7m��F��Iȱ��,�n��:��q��V����.Q}*#C�Q��T��;u����y�իn���j�d�a�ر�)�o�\д�Lf�^��;*�w1>Z��G,�S]::�NC�6���t��I� ��F�8$v�ֈ����X3�j��6us�����u9�};��r���j�F[���bE���ͅY��]�a�=n�xBN(L���	CR��5!`���������0l�[ �sE߿g�=��jS��~ü�R�ȤWs�����6=�X�PW ����P4����}�]D�[5���~�_����]]��x+�����7��<�9�����@BF��ǣE�CCqo�//X���J�����X�^��������ҳ/��TJU�u~�7��	������C�J����#����I%+G(^��L��ݛ�mۺ<)���w�n�ON1sx#�R�F���tD{����ҟ�A�DO�����z��J�.Q��l1
/��l�9�PX1}�K4zd�ʣ��;��[o��C��x`OՀr�����ۺ4;�����k��w�˔7ӳ�Oo��R��{��AP�n�o�����U�i`14Uۛt}���랜K|��{�;׼t�����;�w�S�Jr�˚+�vyl�dy���Wn��ۓn@�;W4.���k���VRBzfd@9Yo.��HV��!�A�v¥k�C���id�?,7�}c�T~�1엯�0H$W�,r[{�t�{˳��J�+*wr,P!f�(l�0��zz�Qk2�T��Z#ʾ�Pes���C�Q�� 	�`P�Dc�y.����+,2�1Rgxyx���}Q�:�)X��y�7w`��� ��r��gwM;�tPc�I!�2�T!;�9X��}�[���F��S��٫��Iˢ��~?�P��7̎��+�쇝�϶���ӝV�z<��=�
7Wv���ޑ��w{�t���0x"_�S=���]̃��sSs�������-|�O�槴i�.D�J�j��]��XgGb�޻�]y��pbMJ��\���{a��B�b�{�Rw�}��HZv�$�͡cB��]^�U��z$�yy'��U<)�>��z5�P�ڇ(�_�z~��o�#yБ�~�Z#��}���cS[c�5¤x���o���G^����	������vg�xXf�x�C���{��82cp]{��0d3�:���-��u�؉wO�C3��3�n����+��ɉe������SNn9#5�컨�ߥ]�����sD̴_����]m`\ᣚ��M�J3��|	�b�T�����_|��n_ՙi����)� =waA�h�&�l�#���5�����H�z.|b�k�N让���s�|��}|�;3��}�(7
~+���,8�����/��p.~~Q{�}݈�-I������47SV�1M#"���>���B�3�OPD|q�����o����]S���M��u%v���aa�2�C��x��wefyu�Ʉ09÷���zF%�}7Z�~���^��g�y���6.�J^zxY�TM�cî����#^��Ѭ'W�����1y^̢3#����e����yC^W�D�C*�KO�,�E�_��k�ᵛ0ɞ󓥝Y�@�d��'pih����>��!d6,�r�0�[[�����U�r���ß��I���F�isV<��=�#p��n�l��}Z�V��ۊxl������ƝX�"�?x������wGPs\B��J��^�	�����ツ:�[[]]}�Tc٫��r�w�0�j��.�E�+Wʱ?6o�+��V�,�U�G���e��,k�];�.sN���TT)�s2�@I"E$���^�o��3tW9���㗩���;G;���I
�w#4�uq6��U��\?U������L��B<e
�ɶ�|߆���?]oG���~��}%�@ϝm+�=��8�ݒ+�.���2�p�_��b[�]N�p�B����!�S�?b�}<���B��ѫ9~��5�����������C¦��Ǿ!��h��lW������N��ow38�<����r���=KmWX�?t�GG��O�n�����s�U�w�������~l6:w�C��\���F�Y����C���W��C^���k5������)��?���������K����'N!b<=:-��1�����d�H@��A7LK����Ǉ�h�d/�W����@���Ctn��
�]c�7_koarډ�ٴ����z�tW�f[��%���Zr�ƿ���x�<k�w�<߀XM�}�ٝ��f�e��,�V������Vf����2��6T<�f��@�3�v�=E��>�3Ax������.���J`��$z_�b�,;�X�y�xz�S��]��������Q=J;<Rg��,D��ww���
�7Ml	��7�Hajc��j�"Y3��j��/�~��6"�(�=��~���͆�\��i����W�_8م��{��8.g�i{����Y���fpu<���ٻ)���q��'ʄmld��N��wTY\���b9+s�,p�T����ϻQ��Nƪu�k~}b(*�WC%s�����S2v�u}�"���Y_8>���!��=���ϦdxL[�w��sq1y����p��C}�o�b����.g����������������c_�+�����\��s�y�v&P!�<���'�Aо��;�|�}\��-����Z̯P]�lr��-��\t�(Al߷�;P����8,e�+��G�~�����53��G=���V�,����nN�L ��G�n�X�0/�
�,�����<2~�i�+�v!�u�G�U�d�1�W���ԭ��s8=�l��5�h�g���['�/�Z��Ɉ(9��cf��H�_4*����#�����2�v�U���Pg	�@m�˘^5�:�`z/����B��W�$Fp�]��@�s���N�5�Yy$�ZAaͥ4�� n�Y��bk��x�1��Y��T��Hu#.L�Fm���M�Ȉ?L?�f3z��&�}��߅�#lM�]�����wBj�g��X�%*�k�K������ks���]�+���4vb}�)!�s):S~��q�}1��y��1����|�[����[��\^[ܫ*����u��}B����+�G��oo��[�+Qs�|��t�.�yc�V�R���.��j kj��s���o\��?�oN���3_���}_���7a5�����e�hsꨯNk���Y{Ѕ�ڨ�>�Ck���wKo�����B�7*�bt��ol����+����c�z��϶�쇝��|�v=�<i�^ꚯywlu�o��o#�Z�[��vu
6D\������׻�O�*�}OwdǾ���צ}:;σ��l����3>����t6 >�P��|�_��?N�����ϯ����tZ�5�㏷�(Gzn����mcx\дi\*��j<ei�M����4�o��ӏBɺ'^�(��~�n�b�j�C
����l�D��#B�U�0r�s���~s�;�<�ӗ��|u/�ɇ5�t{ɤ�_N-���vRؚ��;Пu��R������v]Tvܓd��|�>��� ���n~#۴&|�j�}����^��R�x��9uB�b���'�Pԯ;�a�fؿ�0�% �	������q����s�����9�7$��o��jժYN������Hy?nlz����"��碱g{r����r,?_)��]�{8�%#Cr�G1�����Ȏ��p�%�hy}Y�i&�(K�l��ኇ��P���DC���oL�fkw{cζ&��H���ԗ�i�yn�͕[Q؊��}t��C�}~���MQ�2fE�.b��U:w���ء|�W�[v����{Ӡ��y���ʹ�{޽W����y�<2�JĎp�������o
�U=�6j��d�p=ݙ�ry��<�e]	�#�ᕂ��J��z�{"����c�#��u]�S���-�R�Qq
�Vek����"B!��e�!�}������V�=�;�G���s�K0�L���,���6�f�j�4A����ݬiӍ舸���b��:�o��(AD�n���gd�N�}P��R!���Ⱥ�]�o�����⭙���9��6J�2iɉ+v�J%Ìz{^�dxkǝu+v�i�*(���5���&�B`��E��$\���d<��S*K��z=/��JcؾW�;���;�N"��xB��q;5�k��pc�	�Gv* £���������uff;�S��[�$/�7d�h�L9����[�Z֝i�3�Dh2�C�ª���F���̙��n��Lt%�c�Hy&2b����
���>eN�Ò^�c�E�X�Y�AL�y1"�R7�|�鼼�ؼ�8��}����K*�Bȸp^#?8*�8n�$/s\(`�j�t��alM	���չ-�{�����	F��MmD�,�_F)���
��g�w\jR�X��F�N��x:h��ލ���h�������J.P���e]�x#:2n�m�Y��m��]L����F83�J^�0:'��{K�^~���hS�j^�WN��T��ŏ\ģ��n�f;�����*6�Y}p�e+�]\�
1�-�-�{N���}����e�\C�w���D�i-VV�������2��4�f�e�wd����N�Nfνʎ*���ƫ��m!N�M�R��쩳.��F}�INk~mK��}�2�r��A��c/�'��;#�n��$��7fU0��nh�=�clO_.&��#�W�<��˛�@�%��0��؊�;ǳ�)M�{8���6�^-��1CZb8r:�g��{J��P*]�<5����<��p�&(�MV��C[�7gc�K��S��6��.^�K�v�p����Z3h���4�ۏD�=��Mu����ܲ}��](_EVB���Ɏ<��RWk"Ʈp�u�*'�BK\ᮙ����ݭ{Y0.�knp�Z�oMt ���y|�Y�^s�R���L�y6�ot !�u�v�u�Yy�� �/Qon�
��q�� �=+t,�E�)��+>��K7zn�f	m9����F���:�\
�Տ��M���%�K�j�JO��̫ԛ{#�2Y:��6�iP���� ����ĕ�ݮ��"�vU�d���gds���m�y�Wnօlw^�ˠ�s�D7Ѻe�	�r+�>�����Δ�:�8j0[>�2=��]��K��۵���o��x��|�>[�]���|��z�����^�)7,�����.'�g1W2�������ʫe�ЬmZ�k�1XL��N:2a;�&ާ`d���0�a�]1Y��[�n����T!�����j�g&��o�ޑ�Y$�oCVF�rV�5#%!.�rs�M��٧�^�涶�h`Q}�:�9�M�x̓-yp޼���W�)><m����͜ku�/�/H�Ki���K�u��fS�]�������u�ܛ;p5Z��m	�,�&ty�0�Ұ��7c�흼}@�uP3���[��9�/8=�HR<t��>�
���M�4>B,�+z��Q�ur��"3�%�m���ZRqz�rr��˻u��x|�"���4X�.EP�ږ��\-�Yk��[J-�E���E�sťUJ���ړ8~�8x>�jyK�Q��UE*�J�#h�iZZ�Z���%�)��Jᧇ�2ָ*��'�X,�X�eiEփr�iW0���r4�77n�Y[K-�<<<<<���rҷ-���n=s�[Z��p��V`�-Mr��-���˶����X�.������Ç���pˎ3+b�0�8���E� l������,���ݸ+�Z8�SM<<4��b1�G&X������!ֱr.1�si��fn�0Q�n&:ʙv���ĹQ��N�<<<
��k�QJ��U���w&�jL���T*\��WE+]�0*R��+��m4�ӧKx�9h���^Қ�o9�kF;m�b��q�2�0���2�h��+m�ܹ�G����<Z�մ�na�pm����k}��Fc,o����v�\[X�[-�m�&S	"Q\SE�F�*6�)$�eEh�.ccW˟a0ثN5��%���\��e����=�	�V�"�����Թ�ӏؤ�CӾvw�"���c��B�M�w/���D�p�[���^a���V9��~�>��в'g�n�s����a�����.�!d���E���=������<1}^����u6��b6�%��%�@G����	��E�^g���s�eO�ϲz����IՎV����~~���.c#h7#G3s�v�D�4o���M-#k��w�P�{4/�r�t�a��3�J;��f����LFC�(����.��Tν���)[w�Z�M��
�螾�k3��$�ջ~߮n'�4/�W�������=��t/�f�ٯa{���x�/U��'�ź��z7���,`?����=��7*�:�˙��n�e���V�Pņ!�יU����pu��C�B��#GF��bql�H��y{ܷ��b���/�X����ƻ�{~CU|9#+E�V;!Ciy	�0WL�]������KQ����8<������t��t�]�
m	�{��bz,�
�7�U؉��Ůf������n��6wR,"���l��l��ə�x�/<.��]C`�����KXqp���MŽ-s�M�3}˲N�1Ig����@���i�s�a�8<R|W.NJ���t�|V&v��:,�Ӡ�u_Un��!�}�"mJ�ea�G���A�7}f�x{2q�c98M�&-���է��3�38/��uxUuA��ݡk>~αꛨJ^�:���楙ʯ�E�Vo�%���[��^P~a��{��JX�dd�{{�c$�bw]BA��ҵW;Jv{Ua��p$�0�(����B��������{ꫡHWxH^��\s��n�N�+��9���೮�����ڟ_W^������_�P��z7#�gf춺m�h��f����t�w�Aw"�%Vba��~G����;wyKX���`E��u���ڰ����!p�{��P%ۿ2�����A�n	B���*�w���U���� �>�Rk���m��Ξ�g�?��nc�� i�{Ħ��lz�qN�r���W�뿹.w���u�l�@܁_xf��C�Nxi�N��yC������Tƹ[�vH�����]_���@���Q �O�ґ̕�T���nnQ<Ž0ޛ��ĺ-�hf�Ǹ�J�/��-wh��;b�Fe���s�����Y�:�-�����bR�U2�n�Ɍ�LT���F�`����?|>j�8�֨J$��T����������\��u5N�R�]qӿD��^{��]Vn����H4!�����BRB�x<�m_���$������_yھ�sdG�޵W��´EHC��9�ϳ�o�0d��iZT�p�� 蓛,��1]~��,�b�<�邂#F)2�_�y����t��_�U�W�`��p{):�K�&}acb�#+��$�� �0�|�)*c55u�|u^T.'��=�*�f�	C5u�B�s��[�`ua�;�a������5����'���z�eϹ7���V���Ȭ��FU�� �=�y�V��A��6?u^��?�b�{~�q�;��m���;t���O��9��f0ߣл.1V���n���{���X-	����>�z��\�U^�]�Q����F.f|�Y��髉/���	�!���!C3�7�ۀ���_ī:kc�Ӌ~�:�Ɵ>�N;I�G6������t.WV�b6����5�J6r�X�ځ�ѳ˷�3Fj�:�T+z��Z��G��K�l�m���T��Ć�.�p]J�&n:�<3���D�E�u�I�:�p��OOI�UfC�[n
�|�7��[3�ܿ�6�r����V*�.�A���n�9���U��޽�u@�1|�;�\W��4׼�*�~֞v����ȳ���8�AV�`�4fǗ�w[�w�]oȬ{>޵�5�{�[T�q�@��퍐�wp�U���d]����>��'�X�m&����dW-���֭d	�)���w��Q��r����v�|�j�l�u���X	�sb���|�Q�<{}s+�s�W�����X�!�����7�?��~Y�Yy�{<vU��΂J�jA�V��'���ѡ�s�_Hy�Q�ǆa����jv��.���oN�h�����ڄ�;/��?<QU1�xA�ٳw��y�k��ge�?��
�J�5��6l����g���y>�z�Wyywf�z������}���isx�(4��z]l��g��8xu��7U�Y��N���rFD<�B�v��prs��7*[i6/p��Sz��`��H���Q��#��k�7.����\9G7pj�� �'�P��5o&��mʥ�U��J�׽6���Y/�)�����CM���1(����.���Q�:��}���|�hJ۴��KF��<"��u� `���r���]+9=PE��ÙU/�9>�s��a&fFA�A+z�z�Lg!H{������.��D��%e	hO���X������tݫ׵�&�p�cΖXMS��U��v_��G��v>�����l7wmk�lq#E��Z�������w��^����N�=��ڰ9g��?7x���S���z&gKi�|�6�Z��^U=�>�B�d^Y9��[�,�tpN�1݇�l��ľu|����i�7�U������zbϛ��"An;�3��k���v��ǳ���Ƙ��5m1B�4�������[hc��7"�h@] �T'կ�矯�~A�I~
���Y���)�m���fy��׶�_�C�u��AO��c�1��6W	�놖�}�͝�NP5�^�˪�GG�!^�S����,�:�2Ϗ��' b�gNt�Y���?]p^�ﲛ�|��2���.��%�Kp%�t��%u�\w���7/6����y���t޼�P��"OSS�vl͔?����~�KoR�^�V�������`X��M���A�����i�ۂ0�w}��w���"7�;^�Mu�v��Q����mWh�T���z�*��Ϟ	���^��4��xRC"����ܨf�3����P	�����O����d?�����F�Nu�ˢ�w��S�jڿ{�=�4;�������)�QC�oxw�e+�l��09�-Hf5bo*��8���=j��(d�m����1{-
��y+5�t:�����}U���6�1�zJ�b|jOb�ݱ����Ӵ��|���W���y/�HwW�~{�S��w�g���/;�wa�O�9�y�z���@:RbQ��0�׾���%��"[���������������}�\�2�NչP�튚g���Z���e�(am��(9܎����������o{f�c�nFW���8w��I�ih,%��٣nm�r�V-�kDHv.h�=�s��s�\#��PRo{�d&�i���ɢ�K�52�)�[�wFK�@���\vvk6��1V����ˏ���N���E u��WFj�#ղ���,�B�r��:Vt ����`���J3A��9?�q6�Y[�J`^�&lܸU�e��4p���:��)k۔��Q���ѱW��~�7wv�[��v�����O|����{!3���!E(��l�_�;�jއ��@>G�9�;��Cf􃯼��>{H9�~��<�V���U���
��٣�'�;{�X��_,;P7 PC۫9��7y���f��\��6��{�;vթ^�k���oc��B��������9s3k��]%�"�T<��=�W�ܷ��a��X�>����|/_�꫾6cf�$�Yk�0F�_t�q#�!�}�!��2G��JP���"��aщolq���3�Z鲽�L�F)2�X�o%��4��x<���u)�\v�DU+6�\�ԑ��.F�=�b���f��{+��;Wi,Fw9�����s��z�!�ǜ��_�9��B�����gY(_}Y���l���=�MbI��ikC"�nG�����)͖�n_T����R�Z{33��V���s�t
�}r��f�4������5{gux�����g��mHm�Vt(��t}v�fvt�,޼y}o�$0�u���{	"�b�E����.�OM���<[�~Ց���1�¯�Zo�=��_�)W;�g��T�"7ٙ���f

F^D�-g�p�Ok���ƥ�t���:��J"�Z�}{�,��t�I��H�VCC5�
�>��bDP��� �*U^�f��o�4��T��e}�"�$v[hx����P���-��3^�%.Y���/�Z������E��ƇGX��]l|B���{u��߂�^����牫��Jb�<�|w��29�Ou*�v�vuQ�C=�?F׬߽{1;<�ܷ3��7�Kj���Z�+φ��i�����~[c���֙��j�d�^�}�C��::@'������ϒ�n�]�Ac��f������=ޘ̀���Br}�&|��zv�ù��ҹ�S=w���>��^�uV'�y|��|�1E�C��#~���8�c�?UPv�m�_�*2�*�]�g�ˮd�v�ѱѴ�X�3t��+�f�-Wz�O|t cH���8�@Vd׻��Q�� �&���Q�T�s�����cK;D&�9���4�4����ޑ)M��������H4�;V�������%�{�Or�n~���>��,P��]GAA�;���tq��dQ��~ԅ��/�C���������ـO�A 4-��o}��j;�ߤ�qhwfF�w�N��?bA5ߊ�ZI{��G�;���+ڢ����l��\���ζ�/���@-s5��7�f_�Ix`��m����x�v���J��f���gB֋,��[}��<2���>���o�H��{X�/�\����]u�&(�X;�.A�Z]~�k��v�1�!�C޻��NO����c�Y֩5�~�3,���avz��ذw°T�}0�k��_G�'���f��j6gd_�69Sw�j��Kꯗ�(k�����O�V,��^�ޓT��Ѻ���y�����k}�{����m;�w'�DFK��;��a����+�ɸhZ��,�����`CbLM���\m*K_%��	���z����^.�W<+����e8��� p"Iꫴ�8���8�wJۢ�4�����K��V�e�4F�@���zhQ'?P�T.�5Kdr����!�O�v���P�B�c�"�h�e������rK�y*.�D���]�zdMz����2;x�r���X��"$�Zp�ᾜ��ϻ��>��!��[������f�:�c?���]�s ��S/~����;Ψv=�튭��1[u�iD(�$� 㼖���UA���=�=�_"|�m"/�z���g{٘O�_c�S{�_bޠ-n��NB����}l�� �ѡ��ě�3Ig��z���5o޹�z��<�x_�V�W=��4X��xOK�x/�*<�u-��c-��[C�����Gi�{�)T=���W��z"�j��hh��W�f����]��-= �>�T����c�)]Ǌ���rb�6GU1g[�<2|0�ɤ���n�o��I|�xX�{g��ެ�,����~��exm2I�G����'���������A��ff��_p��gh^T��Z*�XY��걃����C<��Y������C�H �		%�T@�'�'�O�?�H	����@��O��(�#�B  @ � ԒBPB$����H�% a � 9�9��   �r� P@ @@ H @ @ $ I , � �   �2  �   �! � I$�H f`�     a � )� �$� �I"H�@ @ ���0 Q@Pd�H�$� � 	�H    ��� �� "��@ B ��"�� ��� (D� I@�	"��A"" �R(�R( !Q!0d�RD eT��� D�� I?��������B~�B�@ c?��:q�חZ�����(��H���p&>~^k��7��x�g9����H$$�m7�5���q�$$�<� �0�����?�����a�����A��'�dO����Q��?�r�O�����g��?��W����?�&���!!"I#  $ �H� X � ��I"$ @` ��" "@@d$�" Dd�H���@ ,��h BJ� B 0 0� �� �  � 	 @ #   � 
 @d �$@ c @A�� B2H�B�D#$� �@ H �`H � �2 I � 	#$���0$d� 2H�� I@0$�� A �H0���q�����A�(�E $ �R��<>��g��7�|���6������S���B���u�_���7�'����'�=��0�'� HI?���?�������!BI��		'����D?�G����B$$���|@��t�,��������2w#?��8��1�6a4��!$���O�G�@�IA	�YRRp6�I�5źIZ���-	�5�<
�!$����� HI?�����dP�D�����#g����/�|��������C���B����'���L'г����81�>���$$��M�������}@��U?����?�g����?�1AY&SY�L@^)ـpP��3'� bG{�;���r�7n+�I��nrҴUkj�n��l��a�[66��mL�k%�Y����l���L23jk[dM������E�kk5�UQM��m�0���2R���[%� 5Em�SM4ڴ�Z0���)��mkQ�30�K[[k` ڌ�-Vf*Ѭ�S[5��M��^�sm��3Za��Tͨ{gee��Sbj��j���b��U+Ij��6L��X���6�M2�����kf��e�2��[fe�U&�l�[[i�4�kFV�f�[[h�+i��ꧧEN�,�|   Y��]���v���{n�;/n������={�mܺ��t2�]�N�״חM�w:�E��k�5�j�u����[j����9A���zךr�ضM�J�Uz��WM{��MH�l�Ska�e���|   =�{���lr$�aB��|8}B�
44(_{�:�hhhݍ�P�;�K\>�
'^�[{�y�O�sU)�����ި�ݜ��W�����ںW;�t=�-�o
^v]:U'��Usm���zjڷ��U6kj�l*����mfE���  ^�������n���N���Fh��]��K������zvi��m���S���;��i�v�{uS�d�juw[m�a*]�[Vԭ��#t�+��nW�Z�F�YhD�U�cJ��  �����}��=�޽9M���Z�g�MS����=9m���=�G{���A��q��f֩�V����6�Wu�����ʆ��,�k��Ժ�E�[M�i+Z��   w/7����U�aJ���閍v�T�d:
�X�5Z�m��l�.���֙�ݦ�]�0
��6�Mh˹۔WJ��aZUjͭl��[mx   x�)�Fu˵�G]�t�k������*�.�4w`�vuHi)�v֤�ֻq\ *��k@�Gw6k���uUp�3ն�jj�	ie��   ��Uۧ L�a�ruѣu�u6�u۔�F��w�� w[� W��5��������z ��� (�ֵ�51�6��mZ��  9�A
 �q� �V @g�8 (�u��B���  = :w 
��  SɨT��j��jU�E���|   >��t �9���  9���:���  �W�� \=�  j   ;qp( =<�` 4���� �M<5�emT�ͪ�iX�]�Q=�  �_� f�g� �y�� 4��  ����z]�  ���  �t�� ��m�  �S�)JT ���i�R��  ���JU � )�A�IU ��F�2 �Q�h���J�b�@ ٪o�?��_��_���)��ew�_U��C��Km�ܦ�VE�{��(W�0 0`��Y>~_�1����m����1���� �6��`cl�ll�`�h���~��������#z�̡�r�+�����7a��J8X�5v���3]��a��u�Af� uh��'��~V�'+�m�t5u���n�q,�/��m�k(k4]+��K�Q����v�:�"j�.�(C��C*NU��6�\%؇�z�DC��+V>���±���wm��EVE^+����������m�Z���L�mf��J�����]`�u�
J�[�ğ5ׅv��Wa�+Q:���)"4إY�)���c9�vAv���=�<2�n,;��5&i
mރc�yX�c�Yo��Z���;���}O(|y�X����(�����0�u^Vfq�/�k8�K���x�W+	�ڼ{ð���Rd�ࡊP�9�Fa$�`�	����٭�B�>4%��ؖ;��֟ˣ��o��+�y�wY��0�v��`:UY$�Y ֳc��HgP]�.	�vM��5؝�@ޤB����V�'ٸ:1�'���i�_o[D���.��v�iB�I���+hj�T�3��N���<����]u{��Hsl[�nql�+��f��f=�6�h*�Tham��9N�N���x��yK���a�i����������h,�|���7|�+�Q�I�8�WR8���}��V�7�.����A�b��=X�ֲ��K��v���^V<�wCZ;�\���W�m�}c���}�����Pv1�ue=ѷ��25V���i�w��cSZ�touq��-���:��	=گ���	��:��hZ�;vP9xWV��L�K
�����
Ӯia�- �ޜ`-�<�ᇏQ��)�+r�XﺫY7�����X�Ӆ'Z����U�t�
�]i}�!����"�J�aB �c�����=:{f� �[��Z�/e<��n���'���3�A���X���n���n�}Ŗ�ح�u���	1J�%�үN�̷W�[����Zm_P�-.� c5��u����m��C4����:��iޚ<oy�k�hu�����2�ߖSē:YLاClSX��˱�V��f��4Q5�^��	v>ԓ�����J�����qD����⬃�����SN�-�w`����\�ba�c��t$��lpj�q6� �:��:�+��H*��ě�o��=�c���w��x���|O_<��}Ee�� e,�z��-5Zlj�a�;Z�״��k�>[X;ε��[�x���>I��jʺ=J�Xu��r�i"�	^m�a�W<V�e�}o9���6��YLa%��㛖5��6�4妵rX�;�W��j��&��Ceٳz����`����eW�*�J�6ٲ�F0r��3��,�f��g�*ާ�X�և]�� .7���zu>��u������(�	�}�ư�-Ď���j�a�ΐ����ʷ�*ݢJ�o���:��.�F����5�{Gl�)<ǃk4��q֡�^QvYc��֟v�P���u�����w��0�T[�|��#|=V,f�l�b\���˵�2�K��i�;z��d?��e��2�u
��n�k�(��A�[hr��5i��a��fk��8���<{�� �Հ@�;]��u<����m�(�N��![a���A�� (��ɮ���5�a�=�m{����*K6����o�Ai��m��I�^�)�@x���X�Ņ��K����Vh"�X�F�ԚB��U�=��,�M*��h%�1�ju�ke���_r����Y�v7Q]�D���4Uն>�r.�3cr�[t�8�CH�b��
Lr�r����[�@]=�y�e���n��r�r�-�A;Ĵ��8C�+t�
L��_PYO�{�;єG> �c�wm�[�؋+EB۽��$�'�ǰ��ͤw4�S�j�]ٔ�_Z�V���]s�c@�˯o��}xE�xUջo�3K�Gl�"��ݢP<��n=�h�7t�݇��Y�I��m�:!�U�:մ���^.��K�7�.ܳX���6��)�&�ߒ�����tyt�.ۥV���:+)�,Z��h����y�[�ƟWRM�f³ר���Ĳռ�}J�"2�����=�i�5kN�O�Ƴ�=VN�!Zg�*��w���ؽIX��wHq��o� ����S0Su���(�%]�C4��cRI�ŀ�^&��RWȳ��K;_!��mupu[eѻM���uܛ8��3[!����Z��"���_1��7c����o�M�(�gU�T�a<EX_�]h%� ��v�O��e7���SU[ݫo�Ǐ8�w���bi �>��=[�h[Ձ08:Z�a;���(o��h&�+5u`�G��%������4i��/E�*ʽ�-��#��V���9@'u����m��k�����o�����!F�v�}�?]i�|��ʅ��iՏ��6p�}ƒ:$�M��o9g�jm 0m;m-\4�Zg��B��N���[Z��i��I
5z5���l�̺��:i��lNGʆ�6N�M�y����K^3ȿ��ȫ�������z^Շ\�e�u����f���K���	M��gu�ۿ��vm�m�{V��;[VQ)�i�8�H��F�����{a���.�^�T�pʴ��N�EV��X�sH�l,�+���;|��f��0Z��+N�9����%t9�V���]��9��U������J�M���u�xcOU�!A=w�S��G0>�@'-�cz��]���n����QR�"�Ţ��&�wc�˶���
A� �[{�ƕiKoҲ.�>�y��e�-^�&�
Ua�L6��t���Msi�Z ����I��V���7�_&GrєI�dw��K��Vkn��F�0-5yz����v�xk�e�&���e�:ӹ��s��35+��uY�!��4� �t������<Z8��՝��4-#���FQV��/�n�u՞4���d ��f��ۢ�qu(^ޝ�� `Ab��i�cw�r����!�V�߷��S#�qή}w�Kz�;h�#�˷�=��&1�L�Gt�&��^bT���.bˡE�h���p���*���v5��気pҷie��A꽲��ۭ��:ݫ;N��'�_:{�՞�ĝwp/qWqA�i�VV`}[Kz�X�{�3e�Ԑ�Í�i��ͳ����i�p�irS�Rx��]�yW�j[�������֛�k(�����*(�g�o1��tۼ5z����h={`��X-�ok �R1i�F�OY@�Rgwo-��z��|�v���-o><i��x9Y��0�ӣj��.�˶�����V���)�y�YV�a�8z-]0ݖ�;�-`��3z�����L�W�u�v�>[WW����N�lS/i��k��!0f���Q'����n���E^s\u���e�k�Df��}��t�vZ,��>Yv��qi�Em28Y���]��M6���B��.� z���kP�p�V4Rt5�-�-�ӕ�v��m3֓b��7�¬��8�g�B�O��UG����'���4�*�E��ӭ[c)qb�~��B�Z��Wq���(V�>U��r[�^=K��0���cj�]�	�^^�7�Y[�r.�u%��.L3�!ݍ;�vƄm�$-7��6�FSu��v�]Y[��.C�>ddjdnm��z9�|7�ז�9�C]Z�zC��ܡ��L[b��W�C���0*�t6�w�mN�sZ��Ҷ�{�]ĢAj�1u,L�����[���u㦝j�t��iն�f�f�7	����5�5u����
/�#_^��Zy���#3��ca�X�Q��۱|ȷZ $�e M�2�t��Y�N��4��I���������>�2���V��|fV�ػg8���Ɨo'���v2�Vpop����@*Yz���F�ۮ=��K,�L��]�*���]5��[�����U��n��;��_�Q�1��L*��^o��X��c6��vb��+���lR8P�O��ǝY�n;�-=��=��u� ݢ(�_gn�Cq7G.���ڻ6{�{����@�(����_g#����wj�0�w��5x9�� ��AjoOf��W2]���>�����n&���
l������l]>%�L�i�F��Zs����e�w��h����j�]�㔆py��Y��qqu|1�U`Z�_+ۣ�S�g����On���h1@:�N��:w,�Z3)M��s���Ձ���\7���6�^�ci���syŌ�-��;yhU�2͗�f���)Rg���,��)m$ie��fV�٨n��=<V[�k�iu�`t;)4{�v�=Ɨ7��q^�u�66����d���Y���|�)wnR
� X�ո�����ź��C�����׶>�Æ���E+8��V.�ki7��C���B�0��R�GZ�j�R�A�9%ʭ���
�י��%o6��Y�+.�U�*�۬��wo�[�n���]�s�s*�� ѵ��ú=���u�*�N>�YF�v�=���w��վ�3Qcx�۬M�9�k�*ay��,���&�8p�������H��=�Yʝu�e!x��cl�,�5k��,��ɰ,S4�H�t��u��ʹ5$�����we%͇���Da�Ի��Mun����#��m��-n�#�v�}��ڧcp�X5Wk��z��*���A��C���!�zlU�>;�6��"�2�=�Ca���R�\ܽ�l�����9͢�`���`�/�˾�9b,s�ig'�|���`�VVmk;���k���6��Vֆm4P�l�V�4z�4q���;f�[���7��N���I������A���m�ZI�r�lqj�� ��t6�Ļ�cEe�+�{��a4�ݺF���7��RkoV�����n�f'�cZoXZ���i���W:�.���h<(Zd�\����un�<.���k��v9=!.喻X���XG��ǚ��i5��Cz�N���]!w���$��7�Wַ3m�A�[H��eh:	I6��m1H;&�j{��V�� bݰ��NY�J��EV�r��'|4%�f��'���q�!w*��,lc�c>j��y�ȷ��h�>̴���5]2Q@$�����T5V�c�Ɔ7o3z�ܐ��2�w[�Z�q�%˅�Vm�X	a�tQ�����`#.�]2��;wA
�T��u�/Vj�G��F�Cw���Qt~u�>�@�,V;�tI-]�d���Ԯ���ׯw���mf���|$���җW+t��F�6�+��y<�����]X�o�FVST�F�,�i�]�Xj͏��J�YF���,[YW���������I��I0Y.wFݮ�z����m�ܢ��"��m�*�T�<��5` ��yF�V���TFj)uj������b�����4�n��"����t�cG�BK�;|��@ֆ)�!c�x���C�9��WK�w$Pu�0���l|H��[Kz՟���VN��maܠ0ث�3]���K[xZv��,[y���-�c�{�X�M�*����K��*)��Yd
�� Ӧ��F���\�wY��n�{Ɵ�k-m�K��A��+E,aՂ��㝣�"�u�w	(��ݘ��Ɇ�yi�.��Y+P5|�ʷ΅m ����Xs���h�|�1�^��ͷKcuƅ�̶	Tp��i���S#r۫���%�LΜã^E�Ln y���,q�}l�Z��O]@����`a/�����D�,u ��)ҿ�}J����TO|4h�z�)Wm����+�5�X��i�ޫ���ڽd1�kM�	��#�5|k�W
Ygu��A'����y��n����F�6qf�iT_f����E�Ci��amف�]����c�ku����ZRv�͡|폷)X`R�-���wM��/pP�Ae
F�q�嘬m;����,2q�z�K�.�[-�L���ɗ3��ՏX���҉<�o(o�;-c+���N��.�q4�kv�˫�%�}�yh0le����hG��XxnP ����x�acD�XAu��R�qw4��c�=cm۴��Sʶ�9\n﷟&���op����iq;����;:��w�E+ޢ+��m7�� ;XX��Y�WOS[�V�ݏdZ�mZ�y���3��ݏ��y]��Y���Ǆ>�K0m���GYV��wB�Wk,y����kmp8�V���C��ͤ,w�YA,��Y��4�[��z�u֚���,%hnwP+���.��iY�� V�v6յ�IVVM�Z/���'�TC^&�&h-{�F�vr���L6z���4��ݬ՗��v���Qnҫ8�`Q�<KY�V����R�C~|�v��ΞW�6�u��xl 	��z��CV����:V��{B� u���7l��}\K*�Ջ�=����6�y�E�k��m��6��
�WX2����ڸ��g�k��W�6	l�Y�����yXZ�n�[��Y/z��g�6��'|,Sq1��4kV3���<�_V�U`
�t���
 f-��2�μN�������_4��3��Df�}�oO/�Vm:L��%�l���<-����/Q��<X�}���k��t�d ��v����;�yY�v3�S��M���Vv��g���y]�kǆ˥Qi�_Q�V� w���n����v �a�L ����F�r�w�����bJ�x�՝}�p�f;�@=˷�h뼳�жĎ,�����4��X�N^6qm��L��P��{�XEh�W��wM��ʶ��ǙwE�gU�`�:U�b��v�����#H<Ŗ,�,�/m]�,}���i�7lU�V^��i�'�x�kY̴Cwb��h�خ�|)P�Ɨm.�Fm!}�u*=��v�����V.� S[��uN�+���+��ƻm��F���AK�Р5�T�!g^�	敭����1�X����F��0;�p#��ݷ�����c�x�v��W��i X���A]�����
�͐�1�d�PI:M���q�2D�c��*k������]��s>���[�d,�RqtJ7��X�W%��r`	J�s�q�8�rw�`�F�������kU�
���֥�#"�T�S�DI��nu9[����xه��4��؍�$玥�f1E`�
�+���(�|���G��*й�H��[�h�t���(sDY�x��AO�&"!�Aй�P�յe�pR�9��,]����b�H�N�Y���k��N��YUc�%�VIo=]���x&�87�;t��D�:D:,�/�0�^�G��4Fd�y��"���+;(�W,ýSqW7��F�\q�N��n�Ti�)|/Ss^̙�Z]�Z���}��Έ����5�%�u�d��u�Д��8)q}fN:���q-��cy�̸���������q݆5��r���X⫀�׻�K	�N�+�ԕ�#B��Й)�|ܽ�d����t����/�7���U�S5���ތ̗�c�δ�v$V�;���s[�.)b�8\}Xv���!3�;��L��^moGjļgF�QQ�A.1�F;�,���\d{��@�%�`�z�	՘r
��}��O���o��-Q�eXr�8,:��L�hο\��y�-��|t�\�*��w*�6�17��}`t�秭�)\������#i�pR�&c�R�Qg��ֈ�>�+4s�)�ܮ�T!����U�wT.�^V�A�U�z�\H�K�\:��Y�V{��2O��@WF��&�g���ɵ�A_��U�WO�`#�i��O9;��5�\aH"Э��K�-ݫ�p�Mnj+��J���v�t�S���M����Ҥ7�k�N�-rs��S��tx��MX�GA�ZM&�Zޡ�#��f����X�K*
/5�Jэ�s�X�*v����o���u��F���z�&Q]9�L�98��j��.r��V�8�/ǜ����E����z�+��p��j�R�6M�c:���Q��Y�+j��9��2�Ƕ�L��,�ĪND��)�T຺�l�F݇�f�Z��uu����ޡW�3�!�؋�p�N㩌*�p�m��r̮\��8T��O�O"��&m�}�h��'enV=�ً`�2�ƃ�k�ݡ�B����:�j��\�׍�U4^���Ur���%	����O��0gR��teP6����7��N�Z���<E�VC_X�stnq�;��T�ؘ�v/z������éimJ�ǩl$v�v�b�c��Z�q��.���sQ;��7��jOHޓ2qDQ��N���&�kk�mƗ\溥bFS"�������ZX
["��[6��HU�އ֝�wv1{/U�pe�$��}�v�&�e6�'�*�#�̠�%V�mZ;�b3�ep��7/���ݹ��P[�S*;�L���#�*P� �7,+d��\F��G�tN���o/����H���d�&Q�H���\i`ˢힺ��8������Ipi�aVV5f�5[
1��Q��Ю.��Сs�e�gq�JQ�9����g��&5d0
��uc�f�Ӛ�im�4.��X�r����޽Appk�L�q諽� o2����V�g�5ʐ	X��鷋Oc��u�k�]O���ӶAq�Z���-�����0%�3���(Aa��습.ek����!tJ�7�Y=��#�w�'q��.�|�hÎ�,X$���L�E֣O9*;kl��T�k����v]�{�;
`�YV��&X����]��}zy�t*��,U�~u�Hǃ��գ�i+u�'��X.r�Cr�V�YL�K��́�R%�^�]�\�^պ�,�&��]�Qp��ol0p�F��1-j\=P&c�k�t�Z���+M@A�.m*��t-�lR���5�1���.�et�u���R&��cd�>�Y�m�F��"n�I����%>f���4j��|��c;+��8�p�d�x�ֽ���lc��©���;~��n���۝)m�#4^kå"�t+C2��u�Hi�C�b���l�����R���^�:+j9é���3�gF 8��TkE���n\���0ż�>I�$���]�˅�ϖ�����&�*T�F_f�����и�����t\˰5�Qu��|���C���ӳ��"i֬`��$䊢f��<�}�5�Y�VL,��s��]d�QogI�34K@m�Tvnb��ÚβA\��*�ᣋ��2�]q��q��n��i��W+���mD����,��
�0��懸[o�IX)����ƳY=�^�W0S(Ze+hEg	�o�e�����j���}���)���4N�]_X{�|>�3
�ؽ�r.��.`ω�F^S��T��������Ы���-ON��X��b�k�q�����v�f�B4�e|5!.��fIw��t�X�/����2彔�)M��G<%�:K�X��5 x�֍j���b��]8�\�h�<�5Ȑ��2�n�tk4ӝ�]�G�u#7���t���^�O���o��uN}��α\[˙��{�M��{��{+�fX�;26�i�t�;h�gk0���.؋�l��+2#Cv^������.�ȵq��u�y�s&+���Y¤�-4ved���HJqR�U�M='	{��U<��:_lnG3"=%�4�x�f��\�mhgi܆���� �o�QtF��3��-��khʛ���MT�#u������{����Da�3��Vƾ�ݝ��<��`�[R,���ܬ�I]�5.��&�gt��T��wu�õ��k�T�̠�;����侎l�� ^�4���(�7�T�J��HيMcSyb�tD:Mp�*�om��-bs������ݫ���V_V��ڏ�
�4���$�wlaѼ[��p�01+�ov����P��������r�l��ʎ:�KS�(B~��6�Vo*�묁�̛��I^��h.&��t\�E�챺"�h�C��.�_r�J���Һ��Ѽ�,��T���^����*\KV
m��[���MzM�:�Av�|�W5��.#f���Z�U�F���Dx�0��B���	�e\ŋm�50�^h�S��t��wȒ�5�+(��J�m4����ea
]����u!�N� ��tH+V��u����h�%���G�&�V���͓��5���]}{���0nS�d��r�I�Cۮ�`����*K��U�u-��4+_J�2�qa��+Vsq[ڊء\D����"����S5 WѼl�R�L�[�V1CQ���W:��n�lcF���Ⱥ��}��٪�F��b��z���'T��w�nv(�3��ݬ�
.�z�=�,Ğ�i��9����e���F��3�\����&�:����Shu;o�iz��.o��a5���ɑ,��vj���w&�=.��Q���n��VK�©b��}��*n�2�T�Z�|�p6�4W!�/8����e�M�n�_]F����ALxh��;+%m��&���k�Bбm��n��ݫ	���+%M�0���a[�ƅ%[F�ƫ�`��{t{M5oH1e�Y�j��8�譐����!{w҆�Ci;~�>.�*��p
ΘlSKl���F��:��S�U(���p6�	f�Y�irOv�{�"�5 r�3(f�.�7y.�hv�핦�U:���TY\�F�B��rL �qWQ���b�N�|�q�m?�E���٫���s�(&��
��w�$�3R*+ڕ�Ί����<#�V,'����n.�K�m�Ou�B0�!d��D�]v�=���n���Y�>Ŋ,�gw�3-nVƨ�w/\�a�`�
SNT����e'zl�2�`3yn����ɹd�M�J�7u�W�x��=!n�T�V��V��;nP����m�׫���/ֈF�s��豚+��g�a�[��ii<1�O�\V���pVsF�V��F��1�K�ZQ��^���v���W�+pu���3��C+�\ͻK3Hm�R
�U��j8�,W�8!t�&��6nś��B��)W>ޤr(%N��SC��^	YqW1*PB����n�n�m2ةb�'sk�q���b�Lc���p#�KǼ��l�q��m��n�bm[W�-�;�X��z���e�˥�R�*��TK��k:���w��W���_K�����3u�l��n̷hS��uψ`+b+�V�n�#f�n���mã�	�WB�=�Un�v���`��WBms͎�4�A�qX�%Z(n?�]
��|��LM{_���V�R��=���(NR�xsqz�]x9��[�׾��T��o6�0����8.�w9X��K�2)u)�z(���-P�r[��sPg[ܬ��S�܂iW��E�x����`�R�o���b�m�M ��*m[�'�g>�����G�Z�[�\�̏]��	���On���m�.<��Y�Bf�����*��Xp�!կ\�2���ؒf��׸�B����\�By^[෻��Ƴ�6�wz��d]�X�U����ҳQ�"����j`#1
��g��v�֡�z���F�֚�|�����vU�q�e7`�y΅�՛��:���̕�.�o�6��mm9WR3/�\p�jR�V&��,�*Fks2�zsxT�X�RL3�u�V�u�d�Z����:�:K�P�C|�=l�OP�o�r��7/1�׻���/-nk��ZE$�^$���
ޝOy%�L�W@V-��ֆ��D�[Ü��v���YJ�B�T}3Hn�lySb��c�1-��D���K��F7��F���5RL��剕��;l��4�~fW�*����*�Qަu�����MѺb��I#n4�� 5󽙖�����G"�t�����e^���8��zM(�y��mf�j5�cI��f��W�v^e�ݹ�t�:���$�ˉ`CZ5#�:$k(���C��듇�v�p.��h�s��뽃�q�4�Q���ָ�8�w��]k X����	��*����L��?��K��+�6(�tr��e'�9B�|K� =Zj�:n��u�Q��+t |K�zY�����̊DnYѯm��ӧ��@y���e][���l٘�m��#�gs�\+D�"��P�yc+�E���7�m�(�	�;��:l�ݤ�m�1d9��� `wGi�->����ݖEXŚU;����[e��H��ʛV-�b�9õcn����9a@��B���egj�Z6M��QI�^�Rvn�iE�RKv���B�2Γ+=MM&�-��t}s�M���8�	�n<� gv^��A1�ٕ������5�@a�6�}���W7WC�b���aTjaҳr;��hT�2�-n堩.ܷ[�+���V^wD���#:���tp��.���"�c�z�+I�� ��+� Q�w���H�G^QY���&��e�QSVu4���33x3�R�ᇭm�3�Y��a��4�L+�7�5����OAZ�5��PVj�:��,XSNn��o_Ek�����k��y]]K��f9S|C�[غS�nhk���ϓ�ev��nPݭPg�7:�*9G�i<�Z�u�сsUd�������:�f��WеOF�ʸV��:芄<`��F���:
X����}�h4�Ch�ݭ�q!���R��=���T�^Y�8�(G�Z�7Vwt5�)s��Y2&��.�ūzi_r'��C�x��mcK� ��5�js(������>�1oc��)ĭ�<�%����J�l��`��ps�V�����Q�&�I![��э����n��o%��t�ÜR`������y�n�_<,	�9>��K{S�&��R��	����eo�XF�o9�l�W:uJghӡ��U���c�z(vF�ib���P*�N�}n;�rY�W��ګ���r�)�OB��d�N�w��B��4j.qP�e]�ҫ-�5���=\Pq�>ý˩�,�G��\�fܖ(;��Zt;n=������(Y�AO)��Y�S�R�[���۾�O�s��y�����g���n@L�S}��,�{�֕J��n�L�K��Ys�#�Ċ�t�vI�h10�/-�!n�������E�R����Oh�{F���9�*�hP#p���SD�=f�ktЭU�n��o�2 ����#����fGۍ\t�J�mk;)�̝��?K#{=�t<rƵy��p��|]sr�k9ч�l>�Fc�'Eg�6ϔ���;YL<N)�խ��M�x��d:�w���%7�:����a�e�Q�Q�{�	 ���,�:7hevVk2�f�Mv'����wxWS�K�Y��-F	�[��g�%��n���[(9{Je-����V����}כh`�T7�IWp��w�4zſ�V�J�T$��j�7`�t�,���p�Y0�\�^�o4��H�6�٢½��[-6p�I)U����;Q|�Q�DiJv��t��{n.�R7�-i٠��e�;�����P�]ζ�Ό�Jj���;��+�f͢�u+�OZ�K���8�Wv0��iw��a�9]�3��j��V1��O��3C�x�k�q�ܮ�9�*���u�W�m\�G0,N���8'CQ�����ݕ\7��Slも�$�)k�sI6�w��$�>eeܽ��	��g�ڏ��&�ť=��%�ڭݮ��|w͑�ָ�2�^�m��Je��C�ۗ�^j8�p0s��J�k��]	���\�Эd ��*j��FIv,���%������9��_o5 )u\O����j8�c)Γ��u�b�]�����%2�k�]
2��=�46F�>u�/�벍�O��;P�f�q;%�"Es̟)����n�E��l�,��r���o�C,�ڛ�3'
�ɖZ$Ԝ���R�N�U�D:���Y�SX�F��ﾪ����0� 35A�|�38w�)���Վe�!������oc�86�����c5�`�y屏�fZ�P����{��U�xN�X��R����r����x�2�DaY����:P�M�u�S�V/�s��}�`���Ӗ�3�Wa|���@�s`��{�XI;
7&Շx�pYs�9��k{���_e�1�$�-��šOO��W8�l��s%���w>V�q<l-C��-�C�җ�7��4op�i�Xs-����j�� DWm��N��T���t�@������5}҄Fa�s4�8t�<�q����D�Ը�Hl]N����/�\�<�9�*������Ԣ���M��9��ү��e��a6U�{�T�B)�
0s&�M^X����t��m���z��4So&����݆V�(VA�*�UH�'d_f'eY���SLc-y1�	rɓ�j�^��M���ȝ.���n�>B�F�ŧ9@m�4 Hda���b�b�Mv���vA#Z��q#Y�iɳ;jr�R^�����\Ś8�� �<-i�GwR�b�s���[mN9����3x�GMd%��*�ZN:ܼ;MB��=��p{�,j�5F��mru
�:Z
��`�S�m�T�ᴓHU��2�}ܡ�;�˭*��﹬����[��W�:�Y��Qr+�pAl]�|z��yi���%�O
�dc<:�5�u�gv�(��[����qʔ���l��27��bs��M��;#�W�Vҵ��Æ�SZ��y`l3�#����� �S�s�Ә@�J-^mb��'+,1˺.���%��G/W+G�cl����Q��{K,�~�z <^U}������b)���9�]������ڳ\��C�w�L� �)��#H $7z�>ucxhXI�]���(c���+jj�ޡ|-A�����j36gr�O�N�P����<���jS��*��ޥ����H��Xv���8�#v�`\-m0�����z���9�B���#�N��akb�H��Y��Y��e,7�l'S{�����lS��u�y�B&m[g�_�r�n�r>�.+�J�<E�8��^���F�u�q�rTl�9��)N�1 ���=���FP^�b�ޝH蔬ѷ�#�(��{�c�Qz��|�zBۤ[�9�py��,�ć
(d�n�'�*b�r��n�"m�m'+�7M�b�;t�r^�5}�G6��[��!n�b�eeN[; ��(��t��_fNz5��u%�bz���z�|��α��n�6��A36���4��|5b%Q��X��:�B׳q>E��x�es���i�s�{]�e�뾾L�5��Y�e�u3^X=[�R�^cr.�/)��5�h5�����9��wYw�a�Nv�4A%J΋n���e�>�·��R��YhS��*]�������\��(9M�Ƥ�v�vmv���%ԙ8���Cٝ"r ��t:w1k��.�n�f����GH�٨�&�F`�����ç�͈�bʎ�3�ի�b�wGI��ww<p��/�I`�;)b�����<>Yd+�"��C�6��c��x1FԿ��ZK���Gt���폘�2R�%��3��s.�b��g�V5�)V��.�O�����[L鮣f���_0r<z�Y�	a��Q�ֶ�ͬIbJ�w`���v�<M,ɉӌ��,Rf�پ��u�#��4-r���)V;O����q�G���v�Гx��w{����kV�u:�K[B_w�y3�;�2��e]���i�mEo"�6Ww�>� i���y�ǩnF{���A
Մ**�ɝ�79b�	��k�30���#�=��w���e�DV�v�����V��Y�v%��)�RS�s%�>�A�����v�\}���
Y��6-�|ܣX涏N�֐�,�}\x��Zn�Μ�IA��r���p̑}%s{�jfP�o]�u��[�Mg@�*�lF쥠,{�	2�JC��sX���EcC��m���Ѽ�OS��;z�졎Y�e$�a�N-���;�Ɲ��o��Ռ��T�e�LYƖgv��\��2"�Sp���x�sp�Ơ�1�}]����+cHǷDUg7������V��9( Ȭ�^0-�M)q�H|3�;���7)�u��U}ʸ�GH�7�:�gNl�3W��ΚO짢5��M�F'a�u���Rb�h�%I�������{�'�2�hln[ݩ�ۢ&r��Z�6�p�1���ڌ��i�=�G�#
i|�mf.wu��043KÐ<��ڜ��'�H��M���If����s�;qA)��ݢ��gk�s��qIq���L 7/n"u��|M	x>Vh�)��W���`˃!T����l�G�M��o�Wgζ-�{E3�Mo(jP�h�w~)]�ǽ�30s[����i���NQ{N\���h��t8�a��!��Wl�"�t�!&�}�jQt�b�13Xܧ�|�/���[Y�g7ɦ;-9R�+�R�d�����J���9��$h[�����]_R��s�zf1�x�GL��v�4��\]�������>B�ɺV�M3�����,#��kQui�f᤻KC��R���2�p��A� �t.��[�a�y�2�t\y�)}2ojF��a�%9��K[NJ���\v��J�yks3rj��N6w��Mu]M���_r���r&��٥�-�܎kH�F�8sm�����tAi;+�8�@�#x^Y�;�(��]�ݢ�c��{�W]�Ă��u=6�pG�*ԗ�1=�
����(���Z�ՙ�tADfgt�����g8ıJ�h��Kԙ����,4&ĩ�pr��s4y��f�^���/nW]ъ�'�e��%�ؒ).ڝ�M0H�~��^ms�,ʜ�ݶ�Tت%���-�i]�{�^���e���e�ynM{���{C!	�ٔ�5C�X�e޼͍
�>�PCu��IdY�*��X:���ط��ϳ8S�x�yod��e���4�Q�����77�L���-�:Jd�Ϯ���u��!-J�b�hɱ��x� ê<5u�ᮕ}ݔ[X��yH[����F�@��rZ���/p��	���6�f�X�նWwo!XS2����HH/���9N�18�&��ܔ[���a��T�Ǐ)�6p�_7���*���MKr[�0E$�Mk�ʳR�z�v�W�enj@\�ĊWV���m��Y6�ub��%�(EF���a�X��6��W�[-�PQ�1�T�ru�mPd��)��Ł�̼��ز����J�Ӑʳ-��ދ^�Pk&��mgKmu�wE	��lZOG�@8�a��wm�Րݽqm-��F�2��Mp�WS�l֤�t�ow;i*f�g��EqE���!������j��&�u$z��ݩ��FG,)���A7;)cU�n����Ǥ�-m�bB��n̃JW�;32v�e^f�H��ty5�%�ẚ��K,q}��jt���?n`�\��{�z�8��Vw!�2��� ��+�S-a7���U�� <����3����I��̢&�V�Xh^����S�B7i��c��\^��osW!�Y��;E ��ﺆ�ʜ+k�j���W%��N^��/4���˷K����#W�E�'G,���a��M֮�AB��{�v�JK�k���
 �EVtc*.���f�_	I���sgs+Ȟ��m����^���Ү��	�����2ua#�:�Nm�*���mE[��F�̶4���ȉ�,*��)kRte��	'oNьa�pu��ҭ��O�B��r�����4!DL��
��T�WS�N��@�7��lW�a꺜P�I@.��ѺSݜ�^r���*:]��ҭ�y�iV&F⡮Gu8�u>�[:�T��P2S����f�S:�i�u]'���K4��k�iY,n�X��@�픷Zͽ�Mĥ�M����>|z��8d�	9�w{�4��ݬ�f�PX����)�����b�b[X�e�.�	�
��}p���@aťg'�-����娅wS�hK"/$��ޱ�3K
��$ȱ�U ��X
C���];��Ŧ���5h�����&lr,�[��YEMA����
�N�//�W`KO3�ǭ�����\��3)3)��T4q]mC�h�h[h�E��ۥaWu<Me�ች<�!�L��}�bg��W:oP���ç��6��U�[6�:��f��fG���ĴQ��i Og��{����`�Ac�-�]�O�gJ�{,�)�8�ay�t1#Ь�Q��b�7M�o9se��FkuS�f�I*�˹���;.Ƌ��,M�k�)�6���vV�&��X����x�Kcw�dΤ/whG���	����S��:�Y�@���yS%q<�e�H%�@O^���ֳ�Y#�r�܈����|��R���6�d,I��WP#�8�M�W�%�##����.=��Q��x����!v�ƻ���W �Oz��8��W�.ޕ��ͽ�V�oh��؂�"s��Y옲ݬMA1��%���+B)hUn�zIBCN6X]�$�۳����D��j�Z_S�`���
AU���$�`��!J��4��N�ս�U�_er�E��Kvx�n����J��=c^�����_�V˼�4i�}��X��K��_1L6	LM֕�YIn6�X9��*T��N�tKN��ꗸ�E�p*֮����ڳmWfkU�tGl��v�P1���-l����U�u�~�xe�wA�R�У�I���y�f����ܷ��:g�5I�Ȗ�dy^��l�I�//�3��X�|��.��'��[���R�2�۲�!�lW�_v��x\T��Ij�k=khf7�rv�Se B#4�wvYq ��U�˛+GU�Bn.<-	Pv�O>K�[�+-4�9m�+�|2S�:�=�Z]����r�ڍ��|{����=ԝGd�죪[kl4R1$�w��B�BU�⠕X���x���d��m>:�4�Lm�VS/j��wj]ϰ�X�P���)Roi�f����Hdo

·|��R�1C�G�=
�9��Ҧ:2��#b��N�i�֊��R5�=aڮ�8C�[�K�k1\bE���x^�К���J���oY{(u��ڏ�5m����\���<�쾗-&��Sߛ=�22�g[��S�qlt�@��9�ne��M�*�[���[!��c��w��C�:�b4*uᡒʗBk2WR���Va\J���!� Y���O"��My0���4�Ʋ����W.h�Is"��Cf��W3��G��5�i]p��vjn��p^��,#�Bǿ<��Ŭn���l����_
���c�b �i�������ة
O�.պ[q���Aj��75��9eJ_MX�Cr�E䀰�,��'�.��J�yݑV )��<�}'2���d�It�҆��ZZ��#�RU��ű�8Y���ɽӐ� m���j�
FU��-6���q.��5�L�'�v��%�p%���t*���R�]�`���j�*�zo��E<���=��C@;e�
��A!�{��WtT�I�Q��#ݮfe�\�	ܥ�xc]ϑ�m�����䝄�"�-�u7��uWsb�֑P��6(�ĭ�]��g1��ങ�}r���R��
C��l夷��ol;i$ިs:K[�5Ż]%��^�[�� E��ٗ����c1ZS�S��u��0�Gx�;�Zu�>�v<����x0���U
Ҝ���$����j�%)��uq�"�6%9Vi� ;������;�#�������R̒���	f�)E]�5��n|�B�f
Q����>U2����'-�aB��b�����U��1�K�c{7��p�zoV�гx�%e�K��T�k8����T�h�;�u�)f�L5�kTe�s\J�`q�BH1�U�QJqpO�&��vo
vqum�ԏq���ԯ)*�Z�.�۩V�J�T�1
&�����o���
���s���KЩ�O�Krr�:�|n�>OY����Kp�5x�cq�ۺ$�r�kʥ������k0j���XVF:��O~5w���n�خ��8T��{F�)�\���59��1���t9.07 ҝ������͈c�zw:����y��}��nh��ZX�NSiba��j�+$�3���l�Xf�I�w��3��QZ�63�Qd���[xv�<��R����Z�+��dY��9����>�su��Yv��ފ�Z
�@+����S:�∀��Ly���\;���`z7��u��'�%�>��)B���f�]f.�L�S9��E����sEd�R����\�^W/������h#4��㼭���vY���aRB�`�c��k�;J��Y�#I0��%h2����,�}/)�~��[��ah�+�������u�J�Ь�\^ֳ��:��bd�w�#��(T�Wr��"ޱ�C��Ց�L�"���VX;N��4.l͝��*�>����_�{�r��IL�n��.l�[f����ؽcYݘv�a�w/S��N[��uނ�z�������Y8X�.�Ucg*H�b������iku��`�ʷ�`(�ʛ!���'V8���+8եv��¥�e�os�wf�Z��J.[t�YK��$dvSzzY�C�pSΦ�mlcWIg'{|�X\)�8'';����K2�o��Z�թ�v���x!eB�"�e�y+���u�%XN�KFrh�}�B .U���h`�7�$e�8�XB�ͼ����nvv#g�B��;R��V�\"n��3�3Q���U������EN��ؼU�M�4��4�p�:ݪcK��Ι�mZF��5;:R�nR"���&rTE�7�iiptĬ�1�T�Q*�!X���6��T��Y%Y*Q�p���Z���p2z��®�Y�I�x}UU�}_}���A^s)x{,8��&�]>]ۜ7�L���3Z��U{���lk��4�k4��H�O�*s�[Ƹ�Պ|s�[�̨8�\#�)�[@)Wx�4��9�5��U�N�Wu��ռ�+��/(5ʙl�G���>ܹyƋ��]s�˴��t��a�ʬ40;��� Mh�)do��]�ӴS�3J�ٻ�P���*?�����#g����G����iv̲L��v��oZ��*4��V-楷����7'8Eۂ���ȣ�u!(
�,��/8��ʕ�]���u�E%Q�諺"&T��p2��dn��O���D�_v�ܮF���j��ۚX�P�':ǚp�IF�ZG��a+��2�U��-^��wR!z`�����sY�J��E�p�}2\z�ƚZ��-4����{�!�{Cq
�]rœ�q��� r��j{L�+bTsO^�&۶»V���)��Lַ2�4�")���:r���{� u�-�vBh�t��@�]x���}�m<�W��n��i���ƮW;�ٜ)U�f���n��Bjb5�����6Q����1v�Z�ξ�93�T���.�a��[7�D��-�T�Bwo��̵��Jp�7�(�v� A��L�e�͘��ռ�:�+&�]k�n�l0s�ھ��u\y��u:����d .�[+�c�HN��څ*�q�t��i����^�8	Dt� Bb�@�� QD�""�l�ӹ!^�QPI뮹d���XA#$ź;��$�I
��\r�r�*��C	LE
�S�+���S-SC14��Δ+)b�Q�P��%Mby��9D�*��E��J��dE��f�z�UbU�y9��=,�e��;���I$GI,B8y�"9�Ҽ��9eWN�(�i�Kwr=LTģZf΂�V�d�Q�AEȨДft�A�XE�Z��(�W���"���S(NXbae�L���D��q�HH�Q:�ʚuUi4��T{��[Q9Ih^�y�%1�wj#C3��gH�Ŭ�QZ^a����L�V�B��*�*����ȍ
.
t*$�9I\�3�)d��r2Qh��]*��I���v$�Y5VD����33�HEQf@�Rk#���/�����㮢�.E�9���/Bu6�x�J�ѵ��H���3ml�6Ҭ��=X�0Eqe:����a�UW�~��@���T&�����p��Yq|���(��<[S����e�#f��3=C�tz�Ï���abc��6�N>�a�-X�eV���Meˮ+����e}��M���jyT7���F�+��W�ʨ;�~	����^X�LŨL�υ��=��|~?	����y����z��*Zԅ@CO858�Zx_Gfkܫg��S��g��,��c�'W�{=�O�`Nf�O�
��kyz`�X��5#W�=n(�r���+�(�`�~�U����׳'�u�n�S�8{8�a��Z��#v��g^�4�J�S��d�����@��'v�T�ܑKg��ߞS��y`��mq�����S�X�:IӶz������R��N��;��1�&�����R� �n��b�Ҧ;"W,U���)+�}%��@�hw���*Įnc#[YݻWZ幣F	p��q�jK/���η�2i����B�	�`:�Х~�	��M?)�Kw؄O��ށF4!,�e޷:)6����q�Od�R %p�����%8a�Z)3˨�^�u4N^��u^B��ȞPB>b3����5�_f��c���8'�]/�]��V�����5&�,w�7�޴��V��Y֥f�6�u��O�.9�_MC�8`k.+��*�X�*%�AR�FU�@��fE�Ֆ^/u3�Ӟu�h�
N Kf�J�k�1�W����븛�����L�9oa͈��f�'Փϩ�G�"��Aq4���������uBZ���$ա�]"b�`d�#� I���X+|�����ȑ��c��Z�d[��F��޽���#U�׉e
�|�'.]�(��p��y��x03����}��#��f����Z��bS�gԶկ2^�u��p���	��IԶ�A9�z Զ8��*��P}�Ǳ������ԫZj��S=�9	[�W6�S,n��w�>�N��~`Ovz��(�L{�p?1Wo*�Tb�YrֵĈ+oViX�b
�-��&/vXcd�a){p�s��.��U��fT�u��`�驪N���i)3?m�٨�.�H�T b�ex*�/���T��4dn���}���/��v�S:۶�ިN�^����j�`i)�{�$���F_:rJv�B��ԳN ��e�6���pݞ״��Q4�p��w�g��J��CK�/��׻m�FQk�7v��c>^beghѕ`k]'8cҊ��ȥ��R#w]��A�8+���*Z����yFԔ9%�sG`�H̔��dv��{�9���B�Z�D�lˎ��nz�������K�p�,4�ʠ��d�tF��p;Q��'���t�C/6yV�$���_oT����.�:F��yuf-$�8x%GW�2�~x�v��U�N��<�WR$�n~U��LS�����v��1|iQ����@BC`f�I��WN�*�#��b�wt�NBɊ��t>��s��M\>�5��H�1�%����OQ��Q�0-�+Y��g$`���������k8P�R�ki��Fp6fv%T	�g[�q��sSP�f�c�u�K�]Q=�>�}ʱ|��pf���LZ�IˌV�I��c��$AB��{ʀ��3��H��T*��I��\C������~[먓$r�5]'q��Nv�E�#��������7z�/;]TH�4g+�� ��1��6�(kޣW|���݌�3_�k^�p�P�[�m�p�.�d�
�f&,黮����Ŋ�ioP}\b��<�h�A?�T�}ё��)���2���]:�^��WOcߥI����� ri�����P��\SYkt`/5�j���ـ`���txl��W��s�1�h�&V�`@,�,�\�Y�y�A���8�d፧sg�}9:OJ��p�-������o��$�<��#�p��mO�6Q�<�(���Q����1�үtP�"���j�pǽw��T�L��i�M51�3��U1y��wF�哸׹�?e\�ʬ낽η����#����bt���t����<��Qmr�*�&��*aԻhS�����tw]K��Ѹ���/�S7�j�c��Ӯ��\!��z��ʌDX�%�'\!#�5u�ۜ.Lu��p�fO���*��L��E�FN�uN(}%�{/r�� �BV���{'�0?U=ܾ���P��1�޲�_]���w��y�K_���sogx�E.(?�:� ����㨠z�A:��I�����m׮��&�Ui���Y�oj�	�,𸩔"���+ l�k"��
Z1	�Ψw\d|ft���:�ג^On�v�O(�}2+\X�+�T~�����m.�a��R8ة�[���-c���T#�b�Py��N���>󷣩��<I����j d�&����Y�<A�w���k3�;�p��&1)aq���n��p�* �# �j�»���;�+`J�Qw��ʂ�t읍��=¯�zq��M,��J۬�_ ,�Hb�V���2�G����js+E���;�`�+Iw,����-w��][�B1�;*rGH@ͭ���s��%��f0�TH0�`j�r-���ҳ��u�vJբ�|�T�J`��>�U��s��d�B3b:'S�EL0#k ;���1W�߱�ԭ&���<��{�mF��ø���
��c͖�As"�7Pr���s�-W�茵3��t����3n��Vr\C�=}4.+�8e��\~ڄ��A����&1���ѐ�;�̻V�e�}�j����=�q�U%��M��I��R�&z��)d���)�s��&�7K��rQ��*��:��e��ٺ_�k��Rj����5��zb�J�=QN��/7�� hq	΁k����t�.1�,��mB���#��Ml�-�1�嬵�&�y�]�q`"tE���}��Ld�#5=����b8iW����閳����|����8�����P�G�c�=���0�pW��T�W��D��U�z`�
�L&����"����O��[��gA=����/���o�W�W��=�5Ff����B��T���<9:����R�ˉ����r@��N,���ʹ�7� Ō	��|���y��uI�������⣘��eX ĝOu�ϖKo�ov�k.����T�o�*]����1�Mu��2Qw�u@YX�K�Iq���fp�6�9=�:������wf� �u.U��<)��z�[���K���V�r�$�=���3b]�&����R���JpIZ�t�5/s���� ����'EF|[q�&WÛt3�DTB��綜
YR�&��vS���ۢ,�n���ɇ72����r�O��1�T�mTP��@_���VT��J ��p�e�b8,��	��J��Y|0*Rl��-&��@�全�f����!�-�Ɔ�t4K7��=�{��b�i���@Ӄ��QRV�8]���.��������5�yy�K������T�t���r�c��}�F�y,}�.�W�(��&z��5-0� ���#@\��$ �M�å���h�M_�^�19�%�wI]s=�nw[�Y����w y>"����͌�Q�.T%z��Q	5hd9t�����Z��#�z�M���}^�z�\�R\��m���[oШ[��Fd�t�������q?���C)��Z���8\,	�T���mL� �ʣ��Fk��㬁z7�>����j.'/��o�mT_Z�ɓi��9����&��z𻂰x!냇$'�G[|�%y�`�S܇�m
�X���*]�hQ�u�k9
��3DV+�Nj
	A��t[=6v�8<�Wgt�Q�������; ��]up��҉r�ꃻn�����y���D`gɫTk��p2DwX����9��C1c+�S�JR��`�ئ��C�������N���?2j!��	����0��v��7�>Dvߧ$�����+��Lp�0�ஷZL^���%/n;�·�{?��^��3y�r��
�*f����O�.�ޗ\�ܲv�j��0�����h_E�bs`�*|�
��x��Fn�nm*����Rn���_��A��mS>��VL�=�B O݉Y��Ĭ��S��+]:t�����}6ڮ���:rLUO����Z�����U^��k�ذ�e��ҽQ �@LJg�z�_�&xFf�H�X��̉�IKC{;xP�1C����yJ���׫ھ�3�U��nS+��mL_�xAFt�w"l���@�z�v���@<��Ҏ����8�b���l|�9B�`3�	���Q<���*�;����{S��=Y���a��RU '�\�0���.����U,`k%���#M
�p蓶�w&|~��cG��>4�����N�J�*�n �ef_p������Ӹ�@�5�p���@�w���
��@/v��!/�`���2����{�f&#(v��>ΰ`%�;M>Wq������x��u恓�L�ޙ��d���Սjh�s4&�9�(���=�J�kFC!�y�F���[�&�z{�j�]��e���';�}R������sƀ���`N�F. k(U
�A����"�+xAv��ws/��INLQ�ok��3�!��;����V(����3�О<)]䝗س�}]V�4i��6e�p7���K�ɸnc�0�K�
�e8A1�V�qg1����EWF�(��8M�!"�pXb�e��D;/�I��N̛��#]�EƗFI]�T�v��c�t�=�������O������x�u�w�<�'��9���ʂ>��Y^��ޔ��y$�Bu��S�-���yf��
��ϭY�z�3=t$��4���jT ��{�*cV�CHo��m
u��	���P���h�T�`��l�a�%a��^u���`�+�K��1j�'_��t<�"��1����p+����A h���5��$�<��I��� �y^6��d�lV)"e
03�R�w���sO\V�/\i9g�����K�mmVSx��:����%�oC]��wR� �)I�Kޛ6�� �J"b�>oβ��/x���|СG:e�4`wl*{���\C��gZ�c)6��s e���D�u��#�w=o��)�ụ��u&FhS�Z�������$f����Y؝+�zos'J�-�9w\�U�%N�Q�ڊ4 �X
`ΞOͥAd4���
���i�g�O�j1��1�f�_:����+�Qv����YC�Pǲ��3�nQb�T!F7X>c��sUn�=\h�s䲥�t)�'--5�u|-]CĘ�Ǹ�@�{k��sW�*�ϯ�`�E���;��<�/�rQ�� <6�H�������7�� T"�B���q}����/g��7�qָ��p�ި��{���c��' W:�z�����¯�"�u��@x�� TH}P����Fm-O�ǀ*�Ym=ǖ�p�N�1���G��	��{N���T���3�����k�bH��\�?I]�B��1��XWq�j�aZ�˂B�-����Y؍����}`��}�����U%��h�G>fq�붐w�\�.�?TBJ�.��pbc�*y�7��T��)D�@?��#�'pv��q����.����	`�O٭olky��H�B2Z: 	��&*WJb��d1M��*y:��J��qv���j�+3Lj�^��m^:tl����-���كw
���,��GGOr�O�a{�m���&����p�5��9���6�@��L����\<s^���S�x��p0�>ڸph�Z���$Ԭ�=��/�ꆒ�r�i�O�k�Vk��vVճ�(��	y�E���9�
�w|sS����X�O*��y9�W��������ܐ�]N!lc� �kat�;���[/:��pT��=Y�W�5��B]m�� ��~KW3�[�M��d���XLT�늜��	Bƚ�w������l5G�`Nf�N��G�C�V��5�ƶm<��t&��f �eV�T+�|���CUvK�E�4���S<.���)L�^�E�-�䱦쾟^T>)��n�v��Y��{q�&lx}�� f�^��^Zn�尲� 7��\<�!_��1��*���tÛ�i+H�-O�Ȏ�V����X���2�afV�"D�t'�-1�v���f.*c�e�P(��tt��}Q��L��5�֢"�n��[��v�0&�������~cj"�\!p�m���o�(]��a�~��.L��G��*l�q�����l�|���P�/��G~�#J��c�uB���YA�)���[��7M�2rp֑�K�N`�B�ს�W���X��t�����o��L̨������X���U��7u�w7�P�4hd��v^*d�Kv����с��4m���R��!!�:7�U\b���pͺͽԭ�}u�5N���	9�'�c�:��Ŕ��c�Nƴ*7�H0���;*ڭ]:c�\R;j)�ټh��uֻ"n�c']�k�V�$�����B���8+��\+H�{9*Z�j����u�ΐ��"vۅ˕��5�o���ڀ7�!#3�k�����N�i��d`�]�MA��Q�H��D�Ȉ��	L��J�ʚWۍ���#��?GB �IC����6��m��`��1���������
��yW�}}���G-�.��5�E��Bgj�;7��b��E�򘻭v�׭�T����&!Aγ�ץ��b3���kR��&9������vZ�Q�9��q`�m�+B�.�>L1���Z��ei=�}׵4f>�a�ƴ�_[�x�b��XWA��8�g`�PA�]}lU���v��CY-xz�ug7���D^j趣��I��ܼ!!O�����Ϡ�mf�|�43��#1�b�v�a��1
u�<,-����vӰv�boW;��]��g�8��Ѧ��b�QG�Wt'X�4�=Z��=$F�텺�Y�{ԓ�ǰ�Wt1)���e(�ʜS�ݯ����x��c�mlun�-Wh�]t0Y��Y^ M����J�c)V���N�:�v���8SS[�8�pa5�e���-˖��O�ɷڅ����[��u�`u���u9f��V�"L�]����[#*�(@�n|��bV��H��-d7�u$H�5ӕ:a��:8@v�Dkj
�*��l̤�)�e�ǝ������V;{k���h������nrI�wh5�3X1�d�n�T�����oVh7E�S|lg.���lī@˷b�*͢I�SK���8�}�1 �����m�*��ﳇi9۶�!qc�t�e�-��1)ۼ#˖_�%p+�kJ��2���ǫ�o��K�k_���F	4j|��8NiL�$��;����/n;)I��%s�I�5ڷ��d�TЏ��ӝ�����	�b�|^|�u%X�ՏSY��;�j�(��:.<Jz����W�at��s�u1]��J����y,�-v�w�B��YY��.���ؗc��e���bv��D��Y|uu�y*�k�YL����t ���ds��a:)�|[�坢��%Is���b�y:ƈ�u�ȻEM���K{�i��ٔ�����f!����Q�'`�{�2V�p�hP�Z�=E#�O�p��f�k���o_0z���1DW�%�O���9d	^��%p�j�Fbu��k*�b�b��o�a<�sըɇRnP��l�p)*��;y��C;,[�=��*ʆҼy[��|͋�
Vd��9�O��e֞��Nek�̼P&�6�H0�! 
A�Vu�*�a�45���L�(���_;�$$y�VD�*X�fuYH�SH�"���L4�&J�e�r�L�d�ԔN��X�����9�+2\�Q��$'9
a˪jd�%H��24:�KJ�V�r�P�hD!�������DrBs(��euRs�/4�CQ,��H3m!QgeMB�Q"M�*U��T0�t�T�Kj��T
V�V�Jl��0�P�a+O��\u
�uwJ�G\s�8U�hbB�0�����̕
ʽ��I�;�N�*U�EE�H�fR��U��.PVK�NbG��Z�Ur���Y�UY�U��[��R����J!��#$*�4�9y�$Y�dEg]��.ŨY��ʨ̹G"��a!��5�,�K�D�\�h����P{��e�u9UA�L%��?�<������U�:'�7�s*�(�
���HV��͍���\�i�ze)���^K\nC]"R�Ƥ���Iq�W�4�uE��`K9a�<�������E	>!ɼ|��eӿ?�Q��v�����?[y�����nT�v�F�����0���޿��𻝤l����1��D{{��w^��}o������˷'*o������ۓ�~��Ǉ{v�m����{L.𞃬=��P<|�W���9�t;x�����?�yOɼ�&�����'�<����CIo��\<�;��)xJ��j���ԨEO��"(G�0�{޺��B$m��~����������o�N���~_x	7�$��������C��xOI����;I����y:>8���PS�|+�X��_5U�Q�C�|�eeM�W�
��P���"G�����������I�\z>���<��'�����7�99��ϯ��o����O���~�yM�	n��[��������0<��iD�ue��@�����b=�O����NV�,�afD6Jh���ܮ�����)�!y����N����Ooi�0��>��zq���&���Ǎ�P���;��n�l�w��o��p�QX
��i������hX𷒈؏=t�9��$�Y� <��	��{q�Q�]��@�O<G�oo;۴�v���_�nNT=�ݏ	��j|�h0E�Y�tC7�D0%��x����Sz?pxW�������_��X�͏>�y(�}c�1��f4F��{NC�|�������GpxL*��<j�ۏhra��Ǆ��?����s��]oH{�ݽ&���̤
�L� �� ")tC7�Zg#*��`��og�WM�B�>�$E��
@|���o��N���8��}��zO(xMz����w!����]�N��G�}C�aWy<G�<&���Ϗ>���'?=(Rq8����u:BArsۗvڞs����!H�(~�?x7��m�97?��a�~v�O7��7�o(������]��q�{�!�ݷ�r�y������ޏ����������0��y���Ǘ����ک��qd�ͧ�)ա���_���<'��ｃ��eӾ������ۓ���߽�;��n�㿿{�I�S��=~���	0�G�?pzW}v����˷�������xyۓ�'i7��������\���Mi�?))*���2�ˤzN�;�[A��U�ԩց�sU0V��y�x�;r�1���u�jT������I��-���$L����Θ�_K���ƴ�smKa��eVnm.���� �����[���;vƷ�cΊt����3oz<�k�|�����Q�ޜxN�o��xL/�߽q�����]��ۓ
o�Ͽ�˾�]`�|r�>�����s����xw����{?z���
����쾜|C�O�|@"�#�3�Y�T�����Y8q�W���Nӽ�Ӭݔ�[��������ߟ>0}M�������������}@>�X��o�����P���<'0��|�G�<���goQ���k�}��&P������������N���8�x.���ۓry:?&��v������zC�a������|v�<�����N��;�ｿ�����>�eyQ�kMz����j4�����w��yO����1;�{y����~OI�ߟe����ro%����|w��&�ˤ�u��������z:7;��n������aw�k�}����D`��Y��^����U���)[�\_?����8��v��S������������O��B}���v<�}�N��w[s�< |IӵF��p)�����<����޵;�:$G�}���6~��K!��V�׷�k�Ux�{ON9?��C�aC������q�v���pI��~v������ݮ�����S{Bt��}F$ܞO��<;s�c��yv�����[��#�>������;=QS�S�H��Kb}G8��p~�ro�����׻�`�}C�����IɅ��y����ߝ�p~�ro�I�!'����q�!���~����'}����v�܅�}���6�,��R��T��r�A����ս��{v�<���x�:w�i\}B�m���g����o��y7ϟ�<tbw������90��߼}q�=8��������E������}["+]H��X�30*����M7~������9?o��}m��<״<&!�ߣzC�����o*�nӽx��<'�oo;�z��v�P��o?�=x=&�P�[���6���F'z���6����<&}�R�Y�k=�j�J�8�!�Ę������;�aL/��>y�˼;]��7�~Nq����{O	���Z����raO>#�o����?;>�&_��ǿ�z@�����o��]�7�'}�����V�spx:#=�j�3�s����1�S��;�0j��[B���nTM�����G�� �î:����T]�Xvkv�N;�[�܉�L9s5U�,�[S�W�pE}��[�M��Ӝ��K�\쫗4�6�7G�&m��AԒ�z�u��J����!ަ�Ka�"/��U�>�>����yI��� =o�8]��Oɼ?χ���.��!�<����É\z�&�����q]�1;���'���0���ޝ�ߝ�v���o
��ohG���q���VͽNnĨ���|�U����׏�ސ>����xğ�nܛ��|�ǔ?&�������7�<��z߬{ON�v�y����Ν�ǐ��	�!u��r���ɾ���y����q��\��]wV��{���8��H�8|�H�?|w�8����r{7p�E6��C��q�%���s���> ��������P�U?��~����7�9������nן����G�<�(�ozj��o����|�}" �>��p)�;����v��1>����ߟ��}�������x�@���xM��w�k�������O��w������?~�����90��y�����.�ꢻ��-D2.XQ�x2[?�I��|O'X���'zp���v��P�{�xv������=���'o�}������.�~M�����.N����ؓ�yq�Į����o��9���r=�y!^�Y�GwxS��Ah������Ʌ<��!��]�ߐ��X�q!&�|e0�����x~;y@���y�<'��8|^�?&�훧�I$C��,�3x�-����7G:�δ���~�見T>�����?~��B�m���~�J�S~w�ϣ�Ǥ<��N���z|8�}Nv����99�?]���aWe���L&(9h-ǈg:Y�n�Q	h�fu��]�Z�7��5�]�jh�G�"(GЪ~?x��o?ѽ�ɿ~��?;r�ۏ��q�I?;<�=��㷔܄�;����Ҹ߽>]�;���çj��~'��	�]�Z���)�Sv-[p��Ƿ\��+B�6=��ш��o��}y1;�|q��~��������)���c�������~8��|���x��/����m��w�y���վ�ro	�����p/��$����;�U]��+�w�S+<�K"̈�?Q��|�\.�y�ɿ��s��$�Z�CqC�%�6N����������}�v���;���w�¸������~C�a������_��*��z[�~8W�=�!��sR���qc9-i��t+y�ؙN�B`�n�53q��n��ΗVwmd�e�fr�t��;�̺7�����_��楘Mz_*Y#yF��Z"�O{�-�]�f�Kią�g���"��99��9%�M���3q�I�Q��J�=������{ݺ�^�=�祐��!n���~��<!ɥ����xM�H<G~�;|O��>��ߝ;����~B�m���\
o�y>����o�_c{?x�ɾ��s�'8��8���C޶r&�9�˨��{.B}�� �|�S�I�Ž�s�;��7?��xO	�߾�S�F�&���v�F��;õ�>;r�ý��P>�����~����o�O�����S�������:�3Օ*��?t��#��h��c�;����þ;U������aw�j���.S
���M���!�x�N���w���oi�0�����hs��͎W~M>�xO>���0��L��Y2kh���T�EO���p��F����y�oܛ׾��'N��@���xM�	'o�^�}���Oi���y��t��ro���>!�W��ζp;��n����2gcvC�4�U\'�W��Ü}�+�˨�K�|sS���,Sک�H*��v�xW�������xS�3+4�h�Z�_S��2��w�7��x�?2���^W�5�������-��{��Y�ҽG��gS�k��s�n�(�QYd��m +�ֲȗJ�.f9��>�-��Oz>G�v�B�څua��R��0e�&>(V+�Qɀx*@.����ޞ_C���7�&�}���q�����w}�v�4�5��ω������ฺ����>�b8_X�� f�fΞ��:��Hi�Nyܱ�W5M����m�s��4���a�����(P�%3��]"Uj�1�r;l����s+�,�M�V�N���ޠ�#��Kn���v�+B�d`W���2�pj'��l ������g��<�L�}J�5W	\��s2�qMa�e_-iT� gmZ�z̮Vz�>��U�}1�[Ia���W�}+*�m�6�E@2|����ʞ���yp��3�1��>�l����Iډ��	�{�R��n��:Y����6������]�r�\-7�o��s6���E�\'�XKz2+�c�pq�Ń%?uuReӟ��4Xmk����F�q,}��[;���b.�Z���&�Bq�(� 5l��-$Ϧ��Z놇-W��,j��kԺާÏ>Ӿɭ?f[���3AZ?:��+��9����.g)����M����K`Jo�=��B���S&,1��I��.]���0Y�.#I��3l�:�Dߩ�g���nJ�S�X&1�U���p/>��!@gɸ�q/�'���7�}^��?>� �t=��
u8�Ѹ��'��}$?�JdɸM����_��I��zA�Z�R�5���K6���]4|��ja����\MF������3�%��v�N��`�x(Ƒ��扶��Η� ��`BO[!Ԩ�d�ZBE���W
��ԛ���)�>_2��i�0MϺh�j�������m���t�|� 
ir���{�w�N�+k��q��8sЁ>w����uq>�mq*ҮptpC�b�c[m^Ҽ�b�������CA���7�1:X�Y<�SV���<�J	5W1E��W���vyz�wWf�e���hɑuP��֥w)�]�l�Yu�8,�T b�exy]6��>�QV/ֻ��p�i��n�^��1�}ؾ��w����U0���j�I)�{.pov��m��y׼ק"`���"媆��s�>���U�.��yӒb���w�2p߆-�"7��p-�M�I��!oQC���nʀ�5	O2�^_޸k��4�j^��g�N�v����۾śyi�HLL��S-�_�j���[?uDT����Ea��2�ۿ����1r��y���{��f%T�."�H0���T���ל]1S
o���T�:C2��"^fS��R�Ί��(�D�s�r��i,��Iv+1#s��5��g;�3s��[X�[�]�s��w 3+�6�a낇���w>%���oO�a@	N���+2��	8�{�_m������qc�ښs�<��o<�g���H��`�zG�̼����J]�����ʣ���i�
��I�G>s:!��^�i��.%Ո5�%
��+�����w�{�3���-5����=�PĐD�p������ �]_+H�oǈ��<�'��\-�-Q�m5��GNM�;�J�0����*T)�,�;��S��!W)HW���a��ݶB]�*�k[�ʒ5���(��.&�]gw���}U�n8����xh'�!Y�Q�kOڥ�bB�ry��*��<o���G�8�$fn!2B��V+��#�9F�K�G��Uxv�+�:!�Ƥ�|�vd�71�l�y�(9S-N�d��k�S!�'����ʠb4g] a�8�@��_@�����ةz���/c\z��(5�v ԽS�@E�誕V���1Wu���s����^|����E*��CV���,gMS:!�7A��s����P���+)�K����NǞ�{63�_=�r�t>}C)q����6<�]3½��e^�5�>�腛~��&"�R=�~��=��:�{o�\�xߍ�ԤJ#LF����(�2�p(c=i����1�UB�4�3C��nz�l7��J�G�Q���%�����~cܰ�K�-��o�}P�p�)!�o���}�mP�{����F#`�Q��(]��m/
k�C2��=0o�����Z�Ԋ������\���*;���n��U_�iC�h_���+��㡳�Q}HT#�(ﰮ֎Ӽ��}܂	M`U�g&V�r�����ص ���nەlrv��f$��E_<�4n����k�!�v8�e��e�ͥ�Ițq��ksK��S�5Ð3x���Ejk©:�nC��e�JnN��4����
�^��ﾈ]���TSU��&&ˌpO\��n�#bc�]j�X��;y��Z2@�|�.���|g��[A��=B�g�.���,��c����F������T@�рq���N	�]w����S[�̨�3��j��B��({�C��;NBru�D\��eB�FC᧺�/]_A���� c�%_
��.ơoW�N�1���D357�[�<��w7-�Z\lBL=d��|5GNLg����%�g�ԝl!�Z��h�*&���3j
�u�-�U"��<5�K��J�^G��	T�Av#C��W��;ijW!�]����M.ݭ�mQ�FQ�ƵL���9�¾�&y�/��'X(L6}����J�j��U�ōm��K����TU!R5�=�LVWԸ��yq4�����1v��
m�rl!���\��O$-q�aLٔu���1��r�:�I�����&�Qb6��C����Z3��,��Y�]ĵyK��(�����T����Ry<3�x�Nz�xE��5��A;���ޢގ7Kw,n:*��Rl���Z�e����]�T� !nȬr�qYۈ���F�������A�c0qc�p�7�+W.�g�~c�
�q�SڿK���k{)�ѱt�͆�i=����vi���=g@z�55�"�F,Ki��w3tۻ����`�U�_U}_}�N�S�RL���Z"�b����f���7����\0�Ҹ��L�:�^=�SE)ޙ^nվ�HH%�yo�*����h��>�:�^2.X�]s��f�,��6���M��S�A}{�C��VC��P?Ov�L�0���*_�1�Ͱ�8�7��y1��w-�҉�X��{�ED=�n{bS��pcT�}���m$�߾G�]۞�F��˾��jSe��8M}U�,��:zph�=�L�t���Y|@6LO��$�s��S����ݼs�`�x�o族ΫZ�NDrV��RY|t|�t[�-��/�aW�����Vg8����4
�A�))�⺩3��}5�8`k.+��+*��̱��c�d�ak����h�OS��h�꺈Ί ji!�O{�`�9�|4ey�_�5)���O�_^�ת��ј�w@T�B�M�Մ���-�ϙ�kG���L�l��W��W����� X7�hc�H��`d�&�@�����\��T��v}��T4��ket�m�û��-?���mu�x���En�ބ�t�Ｓ�Ez<j����jv��r��wȘ���DUw��wq��+�"�mҎ�����{'ef�V��]��g���L�X7�<��	�xT�y[�eq��]����5TɜK��G�_e�m[��]a�����)�qʡ�M��^@t�,!`LB�@��q/�"x�{*������~������'e��p-��O#񪞚/mJdɸM����e�Œg�$in��g�c���]�Zb��
t8X���%�1CÝWP�rwhƳ�%}%���}ԶԤL����?%*jr�s����8�4XWS��beQ�2�W)�M-ۃʂ���2o�R�C���+Z���I��%���쯪$�ɗyWk�)���CpW�V ��˻@щ�<�_�|]ggd��`�EG��|��Ϛ��!����vл�^'vꊩ��G�k�ѹXܷ�
�Ӻ��N�1�	�X��sΡ�q���SS�\�7&$2t[���N�ܣM>�ˑ��}�����|�9T����(2u)�_l<��WxF�:�e��6���Z��y�闲v���k�L�Z9ܫk�0�9��c#���`"��r�X���Ҍ �+q�m�n{kճ�t�ႎ�S�A�E@(A��v�)œ&�Z폭�t�8�p2��H)��σ�1�v����1`��i��Zǒ��=�8Ӂ�wF�ε��f	�&+m�\5`�'��b�x�,���n�]*y�>?8X*ټ��x�KKk�&�mw16l�vm�Lj�݋�Ǆ011��7[4ŭ�o-2�+���k핖����[kp��k.�#���Zr7@Q�$�}[��}Q���.�^���n�q9��3m�� ��z����6���VM,�w-SqwT�c�M�y��}ݬZ胧��D��N�r0
e�u���qV++��w������*�W}F�%���y�D���L�Tp���o#'x|�F�h�����`�kt2@�=ޮ�Ty<8E��l�O\��@��}�s��W��%A�I�EgAm�\��и���K
<�Y�*"9F�-v�TN�?�^I��eq���$g0@�4��8�-ƅ&^uЮ:aG~�6���+C��In�XV,���&W�j�vN����*�>����~�jB��-�}�]��T�"�V�j���8kA]C��-��Pj��	�B5�O8�ڼ�+�n��@૴�7�,��	��:�2����4-��w��Np�������u�)�V�|��X���+J��'n��[y���4iXX���:l���}Q�L�^ty6�)z��Tsv�#O0w	@��W������T�;�D={1Nܙ��KV2�w��oJ�8��]�W�Ր�i��Eܚv���e7�-@Ԉ��(��S�ryfb�O���l�����n��n�sk'gSwѦ�̻���9�L<�S�nn�C��w*UyO�Bs�K�L1m>�}Ӆ]��ŵ��q�4�Jf��
p���#m��v�AYŗ3t�D�Bt5満氳4,������xan�w����[x��t헉݂z� ;��Fo;o9�[,ih%6nfB�C�7��`��a틟ʬV��F��}(z��I6Y͚�N0�w��Yg����)�k#2wcGS�IM!niRfn�\�yܱ޺�n�QN2M�g ����r^غ�hR����ww����R��:��r�'p���(�j�EZ2�oΨ�Сu�`|�t�P�����:�P_&��m:�֯��NPOGiyb� W�}��eތ�8�.t�9-�-�G529o8z��]���M�p���2[4�i2U73�q"[+if#zsX�6�ŰN����^T�u�_� y_+L�(P���sp.��aת^ �%ٛ[��;*i�X�.e���JW]΍����릖��aq��Hm3]�Du�O���ԭĳ&�a�z�섲]<
�4��M�:�6�*��hW:m�!
U��ؼ/��oqk�Vm<���͎��"�Mh���Y���>�c��{vي�19%[�]�m쏱�����C*ӻH�i���D-I���Q��}�}f�>��{G5Ɖ�-&.��
%b���0�Ш�F���0P|���#�����J�[2��$HYAr�΢A��I5fp��
�ɚ"��"�TDPfE��s�""*�E'Zg(�i���5�16��8]�*3�j�aDuHԨ��-�����Ћ�r9TEATA�u$)$�B�"9f�wr2TD�%p�u9Gue���eUFK(�G$�LS��hJp���SY�N��Z�+�Ҩ��YTuNgRIP֑Q��R�hf�N{���U����ȳ�UˑAJ�E�URA�TQh�;���#�
Tβu$41,��8�h�(�D��i��a!UfE�S����+*�l��DlYTQ�\�J�k*��PRt����"4�dI� �++ �Bdnl��(�����ZΪ���dw��ZEE�DrN�l����lW�j[�j
e���ώ)Z⾴�2��Ȟ�^l)���q�~�6�Kd"�a��#��̦ee���}�ծ��lӎ� Y�YQ���4���ZK!>��f$O!��!��m��S���MO��ۖ�6�CU�ʾ�JwOH�]r�X^8	Ƌ�&��wl9t�NU���� b���QR/��j)�w-�S㺝!��9�1��0'Q#���!����n��fu���+i�*f
���Wz���ث�[¾�I�G!������n��ub�$�U����*j�u'.�
EEꢁ)�b�!�Z�Ui���ą��s��8C�2^XD�d��*�g]���(͓8��AJ)�c�F }q��1��b�ei��D0�̘ߒN̘Ptw�}�E�i�./L�uY+���O��y�_k��iҜ�����*�w���kt�����l�p��r#*�?�D9�nXi���uRd�v0�v��?p�b]y{�m6�e��9��Xyj��:5T�br��(9ٿ���]wR"��K���ӻ���it}	��ԺE�T�1.�G6�0�	��LCG����/�Cɂ.����N�T�S�A+ͯ���n�m���X�A�Բڻ�����%���o�%�;@v8�vá$r���6�Qr�bG7uܵ�o(���\*��{����ֻ�vd+��G�"{�͖�,N�1��6�ʼ���jP �a/e�u�˞6�ǁI�şϪ����+����`�7ՕZd��Da��Ʈ}*k�d行��&��j��U�0�yX�م��%�]��Ac��p��^�%���FpYqߞZ�J�[T�PK��ND�bX~�qs%9a�[�
b��>�I:
t
��KµD!�51�}����$���VGT���)� ]`��S��}�|=���[;���Z���Q\඗q���I<7ۖ�,u=�=�0�V�J��bh5R�����iSp��ð�%TA����ټ�*�vJ7�����O��<���p)l�P�SÐԖco�7�{��7��Lq 7��.޾z���ݼ���f"D6v�U��![WfY�6�a�Ӊ��ݑ�摑wSB�RT*���1��h
 �n"d��u�3�,p\j�p�N�?�h�(��-�ys�Y�ߙ�^�����X�|��"Ev|5�G�Ʌx^��xA8}�-����U���bId�2��cz	��]�_D�N�n�'��3	X���:<���Ɠ��p{+��K�,U��@ތ�} ���6��X�Z �.9�-'Y���Ҷ{<�|�5h�ՕK3�4U���'���;8��hAK�_,�S�0U��E�s�g/U��J���;S���)U�Ρ�"��n$���v�����r���tn%��h�����D}�@��ӷN�	��?~��L����σ��U<�Bw(&�>�MNx��^��R����֡��X�m�!�屐���q���健�SC,�?,��~ZTD#X&l�
v��_V�-��Xq���7T��ޑ�K~nw�t`Do�AX�6�i:�hy���;�|E�2��q[m��3������n�gT�'NiL���W��Srq8�(j�>^VX�JW����u�q��*ZMc5���ł]5���.>'/��^�ex(ꖵ��>���*�]�r�!:�ZW���^�a�Z�h����,W����9�q��c�O�e?!]Ӡ�:Z���q/[σ�L�u���^�C�+��)��J��q|S;vՆ�D��t(�{���.��}B6 �<�kg���yLB�u\�7_j�\�'I�tv��ASz��T��qc��`4v��Q�^4C.�&b�*c��U��g��1�y8�grQky�>�G:�'
J��葼�hw���,Xp�|΋�]zY�Щ��y򚫇��fL=���,P[���>I��X��T��*
H�����4���ε��y���ax�1�md&V5������lu��v����Ggl�^s��`��R���-�̢�c��M�i9&cܹ[�#�9���'r��W��N�����|s?��"">�IqJ�l�]�⤬X	8h%��� ۮ���9�y�0[Z�#3U��ʾ��<�t4������c�FM�2ry�iG��0r���>/{f����.)w��s\E���3����wq���"Y�
��E	�ചU��>e
���-�>�SOJ۶曊�c-u@]\�I!'�K{����=A�\��M�����ۦ�՝n��y8{h�l���]ο�\��o*�MCn��� p���?*p\�%��7>E/��ע1�}⃄3�������7ܧ��]OGD;��2o���>�`��09B;r�l]��:\BK��J��O�A�'`C�&��e1Wp-5�yp�:�1���i��Nq9���9os����^o��(�P�m�ƀ렮�*LA^eU�f�KuA�:�V�u9$�va�=]��u�5�m�w*4�
���Ui�wQ���٩f���(Y��P�ah�I>���p �Lh.p�T��d54;�|�k�m �x��*�G���ۏ�>w��c!Z�r�����0�	�W�x�7�8����tس�ƐY{.���8|�p��씯�_�N�?Jg��(VĜ�k�n�:k'3!��v�ѕ�.TSm�VVH�A�TH[689F������8ƞ6�Nu)�P���[7Ye�v���������A<��U!��K�=�Y��l��?c����%�j0�cӡ��C;LVZ�a|u"֒��A�ڇ^��ʯAhz�p,2R<������9���W�G�ңJl^����ɮ��&���B�D��^�\�������0ІY�yO�c]j���������9��\xAE��A�`�>�.|.����,�~Z폻^�Un���W�8@	Hc��g[UyMc?\
��:I�P�-�{C�Q�Z�����z�\^�T�Q9Kg����Aéс���(�#8;۸y�_�zL�&D�U��UwCP�+$�aW�)�늿�t�8[���v�8�f ��*�S� �j9ȣ�̯Pш�:�^��uX5a@��H�ƾ[¾��t��s:!���`)���Y�I��Vq��\��|�b��gZ��������g�M9���&Ṏŗ8�vcv-�y�o5ܞ}����!�:]�޺�?�U��㒆R�W|�� �:��(:&[�ͦ�Úa[t]o>��4�V�́�di-��E����Ь�;.K��y%�I�g|OkȒ�]1���O��od�[5�帡S�N�Z�#���f��b�Ԥ��!b�nT�ŹW0���������{�l����}�D%V�)�̎f��Cs�è���v](lZ�A�k�
�An8�O�Ԣ��C�7z�v�^@v���<�/~C�{ܕ���|��$�b25�H5��������D��4�^ss3��Ļ7B/������mU1�f��;7������%?�Bx�b��4��M2hs5�-�Sf����.;e�y����;ʘ��5u�������"�wBѺ�r�+P&�p���TE�６���1����S\�'Eg�5tb����8�ʶ�o�2�8p��W����0�''_�A��_sK�8�{�P	uJ����2~�<��S;���9��9�x(�.�oP��%Z�G�V���֋���:�q�fLzT�|�e��Z���v���? �HE���{���q���B�[���+�M.���|�V{�L��ְn��(��J{z���-���z�|��"�F��J�9�m�^����_a�Sg
��&wk8�Kg�*�jK1����Qq���,���j�<�kה���&>�u���|���#oY�E~r��7��{t��a��K|/VS��������!/(
�ꐟ�q\�Gړ*;�Ҧ�R�s��%m��k,�q�����S�^)��]@����BR�%NQL����e5nrnX��}��W�b}�]O���r�T���U!]�\�bqʗ�t���,�c��ruE�dd55���s�%�Y��f����Ý�!�#kR'���b����q�[�ñS��g���G0���2�z�=7}�&��
�W��n�9o�p�u0��\Ƣ���0��߸�	eq�H�ꎍ빼�l��#&��쳄�2U�_Cr�'�'��KD��:��Ll���eZT�u[��E���o�Bt��%L��5�_X�DON�!a��A��[֞��v�dn�hǌ�@�*�UewF���eS> 1P��4����Yv~,�5����X�c>-�'/P�D�=}��Z�&j�cc�'2���7LԞ%�S�w����	����f,�fᶉ������^�Wd;tG�a�_���c�<��ڿ����/���Py|vW;�ʷu;�\<ց�i��G�l�dňA�@ł]5�����s�@:�}2�:B�l�r9�b���(�F+�nf�Ԧ��BW��ݥ�a�3P!^�v�.0<'�˂1�U�����U�q!�n�GX���mJ�5���
!��ԍ�-	͡�k�ͅ�eꕼ�~YiZ�D�a�>��k�Q^���o7u>\;wQ�*@��[�JR�%E[��a�ԏgt��w6�r���Z� d�2�^�����*rq�$v�ٓ�U}�UP����>���@�KI��Rec��t�/v�L�0�#�Hhg������M���V��:7u���U"�7$R����1
��pcqV_Ժ�F�\�'N�%��&��Y���Ԣ��|D.:#�T-Wp�:zr�a��=�L���o��:�jk~+��>���ױY�&�{��&4�{�K��?:֨�uǃ	��[��,�/O�lS�NV+��<p#�s���sj(73l��e@�����ҟ�"��3����NXჸf�tR�{q�1v۵�R��}��r4��c�t��
��h�� ��( ji!���C��4�x�o��ۯ��{%�Ƣ�8hq�_�^�3��븛��:n"����Uq'0��K����ƹq�w3�kmô�LH��*��� XԚ�3�.�1p�ɨ��h��M�,��q�qo�c;�I\,���R!��ӣ#Y���\�F�ܪ4ۮÖ �P
R��Z��SSWn���r�ٖ�b8�Bˊ0�T,���n��ok�z-JdɸM�����jʘ�;�k�c�o=}�ʍ+l+ɐ��y���W�Q��Q����:�aվƆb�WK�VS��'}oR�c�mt�oP�"1�2���s�5��/&���܆�|�:��k��Ll��*���8e��X�U���N�r��Y�e��翕UU�����'���PwE�SI����c�0y��?eǞ��4�o&�?�y(k�
�d�7b�����t���K��h^��Z���m�\h����*LL�׸u�����Y/��+$�gph�\�ֵ=�����N��59a|�~:��Pϻ3s��	�L��*���Xӭ�%Î���8�9b̓�9� */UCK���s
��>}��e�H��d���V.�X�p��9��9|4S�Vf6OA� �]D/��Cd㟱���DsY\>�f�l�{Z���UШ��CkW��A?�^3�*e�똆���p�,2k䧙}�/�Þ�۰#��#5�>��&af�q{$����΅$�U�u��SW�Yj*�/���x��1�<��h�7@�׿w��Qc`wB�t��P4���ל]1S
{Ք�S�W�ٕ8��Z�qC i��Sß�gŀ��&�d)�g�!	�GI=Pf]�Xlڡ�Ã:{)����7K��Ÿ���o�{�(9,Xֶ�1��a��ga�w>%�F���P3�B�\�o�е�Y���Y�.�`�fX8��w7ִT�XE��E��qᡘ�v�|0�Q�*�U�ώV�pc�^:�T�ν�[�>��;&)8�8�Jy]��0����#���L-���;j���r7*���ǵd}r�)]��П�����,�Ѿ��h|�?�:��B��p��p���S�	�M������#��FmW��~�� �b#O`�/2H�ƾ[¾��$q���|^�i���6{j3ZY�ܷ�k�+�AD��꒺n	�l�����Ti�cj�r[1�ͪY6�4&9m�o�\�Z�H��Tl���!�KTt���]��:QW����k����E�W8n
�^Ikt�����_oJu=��$E�Jt����]��}+�0\�xi-�j�{W<���<Qp`�i����ӻ�a2�Br��P��L_D9QO�X�3,��hba�t�v�턵ƽ����NP�ٽhh��VX�j�����<U�ySZ��yS��O'6�_X� �P�s[^j/^�p���TUX�Я�m�OT^��N}�<!��]D����;�s'2�X��i<�}�.�VT��\�\�zDTE��|�1o��S\�&$[;Q��u V;Z;el�	��$��$i��(������/3�ˌ{�P	uF�����j���.��h�[;�w���X>|��tL �]K昭n�_l�Û�q� �k��D�����EB��)����w#a�ŧ��W0����ƪ�J�
�N=M���J��^:;ƈݒ53ᵌT�iH\G@��[���#����rV֞�@��Aϝ�d�MG�/��/��!�� �;:�\�������í�hf⬳�ԌM�ܥZ�����f���#b��m`A�����.���W�`���Y��Y��h��m���v�K���4k(�Y�7kJ��i��&���ݜ++hD(	W�Д��][�_p���fh⒦�GF��J)˨��,WC�Ę*��.�Zq�-K8�ܘ��a܏�.�>)sS��O^&l5}@=��m�WI�9{�bwQh¡�8W4���L�xo#Ov��h���`��+�gR��E�7
�9�L&C��<`ӽ���ҥN�欆�N��8�`��i=l�m�����ii����Z���3NA�.�,T��w��-5�X�s�}�:��7[����l\*�N3n�":�b�]����h������yn��LT��I�ԕ֡[\�p����v�\Mw(�c�3���x[k5n��s۫�Ep��h𥛷vC'��ZqV�ph֚Bnӫd�ڇ�+^C�ԽK~�k'^�!ɡ�b���PV�Ǒ#V��)3f����if���}��Rq�*��p�����Bu�`�htwOVȨf;L��-f����,�ngJr���������3z����Y�{
|^�L.�z�	v��1(c�-�YtH7�kz��=�ZN���9�Ǽ�e��i�7����_	��̅��#���[M����cM։�ւC4�s7a;�k6�y@�9�K�����U�z�Ư�e�Q*����t��7��A�Y�ݲ�%�k��FU�R�I��)t��k����LI
�Ç�7�e��X�н����ZʎfD)������M��ёf
}�
������)�oR�B�]�c�C�sg�9�|&I�t���o�m�}(�X�!|�Z�f�zV����f���5�-��g�'��M4/��jW<�����k���Iϋ�vX�d�ٷv-��c\af�7M�8�d#& ��خ�z{{�eg�ԁ�2���tkw����DYww�4`�E/��ę 㹵i���d��3ؙ�R�v��f�,�Z{��њ��r��.+�F���G���u&8e9R�V��g����1�O�[4V�/���}�V���ŧCI8s�I��C5��#V���n�-�m*k. �J!W�����,�o�Ď�J>�����Oe-r_j���� �hh h9������,��X�	M�C%\ɇ�_iڰI���*=)�-4��WX\k��/4����X���R��1gs%�5�T��[�x-ٽ�-�ճ�Z��Σzoi���1��#iC�4��bɸ�e�*=��.���Y��'�P	����R�L�Iq�O���4�K�U]!Ve��$�H�PY�VEwtw2�!T"I(��0�r�Jh��I-hV)�HU@F�uPڪ3E�4�DI�T�at5H�J��d��)2�wP�.^�y%B�P؈烗��Qp�M
	%ZK��G(�';�*�P��ĮDF�ȃ<�iEeU( �rE�q�QN���G/$#-3"���%�j�$�͗(:�E�Z���Q١G(�Yi�E�NTs��e�ȫ��̢+fx��ݔr�VU+\��V�t�")�t
йD�
tJ�%�V�t�C�yT�ӦHer��΅�"�̊ԣ��J(*�""s-n�૫
�wEҸ�Ww �Y�TEUEQP�r���qȫ�����N���y܈/Zr����Q]P�#� <-��z��szZ��̀�@L�}�K�{�wo%Hu�Y��㴩�I9��<;;36�8��4��wmN����DDG��9�T��@WY�|ο	�X���TP6ں��{C%�����Qc+ަ�������׾�)�\���&��C������[��j��Z��<U�~4��/Yמ�R���e�*���]�X5�џ>f9�'=7
��,�\�P�JU��^⼧�=�d��E� ^��5�س혩�ϡ�,��c����F�7w�Ss��o����}�OB n�fc�U
�;_>��B��*��=���1�s���6"�Gn�ce.M��v'�Q�צ��+�=���3ǅ]��\7�T��b9F�j�^�{U.3�p\∆��
�:g��mwZ�l:#�m�&-�^|W�^J�(�U���ڪ�~��{|ȇ-Yd�J����ʭC~���wRQ�i��� ��/V;NUmږ�UY��n�W�\��?l$������%:���܀d,2���;yן�.�W��ɥ���&�³�屐���q��L�0�
he�v~.�&��7W��m��i��gj`�Y�}��;p����
Ň�V�ܺ�����\ ֽΧg��nQ�boF͠�I�T���Y/y������d�WMg�j;��1g�9x�P�x�䔤�VKq�[�9�n����q��tV����30�̫�y]�aRZD�ð�;5 kG���yJ�v�d�,rN�rn>E��ϸ*{V���3�D�V����N��P9�u�����3���bx�~�^�C\��]��-�[^+��i�/��U���=0V�D&��=(;b,���||K]� ����bK2�=i����:�]����֨߫=�5P����E���[�Ҿ��o�T+�`�W����c���V���R,<8p�_.y���uI��~�;�y\7�.,x�����%����nv/>�f�<��X�
.� �}��crG|�y��r�ru\�U���X�t�K@�������m�	�����j���0��Ξ�!��j0�Ҧ9�K���U���:M��2�^�^��`�7�uM(~kTx���aw����G��o���=u��e3�۫��zy�~�a��P62�2��*�@�E����9�}<U�R���M����x�[��A�����!�^/��:���h��"o!9<�P�H���+(��r����(�.�����v�4��4u����>��C�4�&��g���PY�캽=I9��ε���ɵ��Y쬱ۢ��O�0+p�N�vٍ��:Bc����hK;��}4U�}�L�2��8�t��fin�
��"�>��;�V�z#��#�&�-�έ�Ȝ涸h�t��l�7!:�&�1�����?T#�"�:LK���ŗ�nWn7#)(�%]QqFܸ��.�Ƥա�9t����MBn��o"nb��
�C�n�Y>�>�/@�cz��ai�������Pɦ�p/� �a _G^Y�Q2�_p�M���u<sy3�||Y����*��:��r�o�=���GD:�R�2^�!}n��ٵu����H���62�Y'�C�(₝mv��b��Zkz��f�}�Ab����_4�r#v���?2i�������� u�u9�&Q�2�r���n�R�t�osiޜ�{��#\Gj�df�C�/���ܨ�.o-����F���-���`D�u�}ʺ�K.�m���T����m����P�"���/T�����_d�{����I�.�u�HH���Z�x�\>7��V�Iz�AT /�$�.'�Cd㟱��&��_�ep�k���^Y��~�]�^gI�����+]z�n��b6v\�JGYZ��C�"+PU0۩�+���q���5�:��F����%: b�Ɉg���J=��(�`�WItKhc%�\)�q=5���ví6�gzG6ޑQ��/#ti��4~��lm[�҃��]^
�W�;r44inR�3m���SIFFglWZ�}?UW�U�o�=�:�ԸV�����y���w��H��KDYw��,�g�/�J�����ٜ��j�l�wVGP?W����L����-� �* � t�>�ݿ8��tb�%Er����c����|!�X�&�dB��~��B���OT@H=ā�ϛ�Oz���e���ί��N�]K��ţLG��8��@k��eȢ�ꂲ,}Oo��鷻�lm
͘����jrz�
�	l��
��K_\U�:w.�>;�	�M�* �(H�Y�h��[;1��{ϩ2׾� CK�T+����J]��D$�"����{X8�����Q/	?��`��3��8��!E���!ױ�$	�GmI�+yJA�KjF}��"���#��3%�si��r8��.sIy�Q
��U�h{�����Y�٭E�:���c!�a�B�;T�EH��ѯ�L�c�']D�?[A�]��uպ�W�����U�ܥ��ծNOE��&��CS:艌cW��hO.�^OդyP��D�-�6ϫq�;�oUX Ҭ��t��>Z<m@�J�+ptZ�M�2��{W�p�֥f&0�[�I��nm�����0֌�VGe��w1ne�6���$� %���+��.�y�t]�����seY�7&r�^Tl���8bVN�*�����ʕ�[q�q��Ҳ�;}�of��Խ��ᗒ�7�����|����U��lVہ\���}�k{Y:�i��+_��&y�]=���0�@��ǰ�MB�y�+ͦ���?Nmi�s�}s⨉��;ôb��i�y��,��+!��{y����ki����vU�c0*����* J����]��{o�^X�p�ܤz�:���yj��P�*γ�LwTAW?��ˢ�W6���F�j�]도,?_�����9�c�7��}p�YW�������'��s��F�S���U�>�Y��Out�����^8{P�{q
o��
�dgw4-ϝ*J�ٌp��	��)u��t�l���4��m��`u߷���S̃�h�;�5<տ'�P�䬫mo��~����gü�R[=z����C�*��m�-=R�w��½R+7<ɪ���B�9hw��m�����:���%pFVCYկJ��X�������W�V�����+�����f��JN�՝)k]�c�\y��4!n=/����١����hc[�==������*oZ�97&1!�35^=��^�հ������菟f��J��q+��X�M�.Y�D)�����y�ԭxf�tۦa�)�+Ni1QSM�;QsV�����q0�3P�=P
�v0'�"stj�̑Y�-��\�ɯ�R�\����BI�a���ʞ�Ϝ�jnC�bW���u��p�j�s�K2�%,��Ž��&�է�&�]�7��G�]E
�N��h7<���σS*�yW�SٹZ�I={�z�3����&z�	��!9I�e���ꐃ�/[ʫ>{}�j����V�%<V?s�����Ӳ���x�D]S��5'�s����l���ʵo�����nNl}�����8�a��x��.yũ���J2�W9�'�C��2���ӴQͭ�O��^����]�Q=��A�͏d�{ZF���2z��f��/�k�	��X�v�Ӑ�.:y�t5Z�lvjXݦ��\���f�3�$�f��p]	,_G��:di�w�T+��c��v�<��0.ŗSu��E�8��0f��a��y~"�߹�$M�����p)���K�mA�[� ��ۤ�|[�]�Q��&�P��sh���mL�ѽP�|0�Ǯ�� ��>6���8��U����V�'��e��m07��TF����Q����kyp�7�S�'�F;|��c���e8^m!ީ�h�Ǻ?����s�5�=���j\m���-�{�i� ObP��{9��PR��
+��`4��3�9��<�,��Jjb�Ks���]��3��e���;��0��1DN�L�W���j�a�>�<��.���ܴ��yПh�le}.��B����l��nr�v���?7�)�`����s_�o�zET����	����o����^��햧�V��l��,���[���oQ˙m�h7�A�k��[��ZJ&���K;�aͪ�pEٹ=���߻Ƨ��[���e��x��|h �oc]�su쉎��)�<��_7�q��9�}祶��K�;��k�/+m��׍�/�O*�ٽc���@�U�'Tڃ��k��y\����h�q�LǼAyC1Q������
tyk��^rn�!i�묫��S�.�#ֶr�����y�����ߟ��wbR\z�m-c��GJt�+K�;I�O�Ҥ
��a݇k�Ǡ<�^
���pfq�W������L�Kϡ��[Xv�X���U}_U+h��SV7��*���p����8�p���F�+�+>|��)��_y�<囮����Z�T�m��=�.;TLV4���<�;�[?y��$0P񴲖	)��z��mgn~�����)���c�K��޿a�u=��l���WFٚ��i�Gv�So���*���\�d�}p1GTLT%͹��a�ΫL�%��s�RA]Js1�x�3��}�y�������
�l�\��\<�7�IW!�c�Zi�ç�gr#��TV��\>W'��Gd��}B�ONO��{��o�O\ڬ�����7���Bi�UGv����)��}ҘV��I���ޯ5�ou�*
�R٥)���8}V�e}�w�s��&ye�1�mb�wf1�s�A	!	v��寧���q��y�ظ�T�uqZ�[�1/����d)ߴ��7�~�<M1�DԞ�W�/B\D v\T]w�J��dPː����9a�b���/J�R�f)�Aۣ��K=��Y��*z�PJ��Σ&-�Q�z������+9F걖��.[��OS�l�� پeovS9���܅��D���{�fkdd��l�S�J��菾���]ru�)kS ��=ܢ�D)��h%��yq�:��E��b-g�u��؆<��pw��_E8u�=�CmQ���[eg�of;��)�W�w���\�	�T�Q�I1Q��Q��#�T&��L��^��G��BoF��Sg:��י1�n�:5i�)�����$sn�vy13xmݶ�`-]�s؜�������ټ����sy؜2�\�y;��*� ���o�Ʈ�����P;��a�P���.~+bg�Ӟ^�m�+�"]���"̿���G�~7]s�N`{D��D��Q������r��;jy�u8�E����>o3b^�їg*5ʈ4b�,�	P��'���x�R�2�o"~oZ��)���M��\�;9�1�BfS��[�΅��p�ƻ�l�c[�m5:��_.��N������Q^�r��5���n�kϭ�z���S�q�7����¨�qj��3M�����mugn�:�2ڂ�+S��T+|#�9����*S��|��X����_^�r�_2�t�x�m9v�+�0��Siϸ�L�x�Ka�=���_W��g>��G���*���荮*�Z�_�[���o.1��M=�S|���"�Q��Qy\�7`�Az��+��R2�<��[�d��sזMtΫêƽ�0ˇ���1��*�#w�>�O����K]�ʜ�X��T�@d��n3�-���R�����Z��7�	�ߘ��f�}�j��7��M=�P�Q.��D)���A<�Wd:b��9��\�X�=^;t���6�Z+A�w�8�=P
�T��� �܎��e1T��M}���7��I&7�+�Sn�p��~�+��Ƭ���0o�u����NGb��x�Rz�f�7�\����6���Z���(��	"/kM�)�~l��Qu>��{9��yf�_Bi\��Ѯ�\'�i���^ ������%�V{ݯb�R��}�ݳ�p�C_��7T��5�5�<����#B����Gp��@�}u��	���8����7�"�W�ZKEʙ�U�z4�����$*-��T/�ܤ(j������ט`Ot�E�z� �e
HoK���:�MK��sh;�x���ڭ�+�{We��,��ïi�E�1D*���+�l�Ş�ڢ��M�ˉ��'m=�κ���jv4�_^���<�lX�u��Ř7��(��l���yg+�O^�4�f֜�a��=����F�^�'��vi5k�W]@n���Gu�@L�[�ie�m��ѹ�ql�U˜wt'�	ʽ�(SȪ��A�4ԛ����{#��s�y��`
K��ۧz���`HU#֬�<��J͙t�Ĝ����oy5��K6�:� о,��Zz���R���榢-�;����0T���2��iٝs��gRM�w(�,8���x��W�]W�W'HŁv�_@� ��P�Ov����pB���]�����1D<�<��&f�t��J6�Dv[R��0�q�"�A���o4�̓qb�+Z�=�I�+j��P��}�#��\:�
�@��V�*�<uS��y�A�h�a�=�z�]c��.+�/��mc,��.�.�����7'm�A��P`�Vμ˫����"��m'yӯYf��	yy��B
HwS�W�BI��ݶbyƀ������k@�	ya{�]�m������xd��j�	�D
��dF��e�ֲ��ĥ���
e��(�"ǦS�*m�.�i\��tj�[M�+����+�]�-s[��\.���C���n�-�oo��t�*<7i��·s��\6�Qy�>YL՛�)]e�j	1�u��6UʽԆ0RӍ�6m�w(��_�`�9+�g'f,�ģB�w[��Ʈ}��� Գ�O�<���ƾ���!�p^���7)P�͍�"��rW^A^���tЙ�7kCU���f�W�������P2��V�:��V��#P	����	p z��]�f۲1,Q.��>.9�feT��co���C)n�jVG˺��j����9��wژ�S�6� Մ������"�خ�ۭt�c��r��f4ɹ9*9M����ʆ���*�:HQPc�Θ��8h:���a&_F�q�"}�w:��M�[�K}���g�����֪�YN�V�(Γ����������&Kk�Y�o��̓���}	Z^��+��ʽ���w��Yk%C� ���[���n�|i��*٨U,���%�WZ��ܗ�q�������T�1s�h=�|�ǽǑ��9l�Lt���d4��=�\�y���}��,��b��5���� v ��:�z���vv�7E۝�f�F���y���5Gi��-��[q�������
��=ړj))S�*;�Vk6�6�Ƣ�k�%�w^j˧���P�|Y��܁��^�M�I�Pr�U���hW4�����<9|Ĺr�X�QR(DrxI����Tr"��AT�1B=��1D�RS�g8�r"�$��W\�P�#��������+�'

%)6��u
 ��!�(�C��f˄�W9(3"�&��K����Sһ�wt�Tr�*C�+�C�QD.;�
(�)β(�wp2M�¸�QQ.��(�J�9�W
�$�h�Hw7a"�WNb��GvP�Z�[p�ԕ9DDU!���]��S�'w;���:Ĝΐ��n!\�=,5�e��9A�]Z�:z��k�#���FJ����U��EAQʎQ�f��¢Qu+�z��G�̓�<ˇ�j.��3*���GdW�pŇ9Q4���'wOTӭE�;�":��x��N8���eET�I|�8\��Y��g��>�1���P�����T���髌%�0�'X1�I�����p�fr���h�vVLI�݄���W�U}]�pt����E/輪g7�>���%U�.�9��i�y�t�L��jS�wc���&+;��q]ޖ����M#u]YF!�״�s�J/}�s�w�r�aɵx�5}+>��ݷͅ�ԟn�y��u��ͺ��Ⱦ}��`(V�
�f\N���J��TlT%��C�պ�[�n!w�GT�����L�l����<����=��p�����_G\$۞U��"��zd�h�ظ�[���q�����>�KG�$wV��{�kCb�쉤�kۯy��^0���N�-�ʄ�m����{>*�!��|��s�$3����z�G-���7��\5�vk�ꈷ-�Q!w���qb�Nބ��Nf+��r��1��q>������ŷ�	����T��w^h7"��������	��3�{}�C�eM�	4��n���GQj�c��X�p�LW�ˌ�U�.r���חF����!�Z�0rhA@��}�tu��Jxh-�砖��Wj�R쁄�vL���ġ�fy��4m�'�{.{�Ŕ�Ä���s�\J�L�)���U��mף#���}��UT�y) 5�\P���C�����Q��oߒ�i���l
.l�Vb`�Z�H�O�P��v�r6����sس���]�<��e��(֨�#(�i�Q��j�^�n_V�w������0}�x�mfJ.m]�s�ۄ�մ�ӄz!7i<��]��5�����P����]��6��������"�����ԙ�zz�C�9Q�*����g�MH��K����om�LWmM���V��T�cNʗ���ϧC�Т��N�{j��5-P���̯���nMM�I�6��1�cU��͌u���op�~<�#\�3|7�k��ڦ�*�<�es �T����(���u
��#2vm�JTz�u��jG��̅�I[񰠿>[*-�9訬�t�Y��{.$N&p�x�������\���<ށ���C�[U����4[9��i*��yE��nx�0J����H��6�HPu6�\�3oګ�8��o�գ�������&1������{����n[VL=�H-$5K5Y�����v.&s�sK�0�;����zM�{��� +	Cqn���ﾏ�>��=Yo�caM{���U_-o.���=���Sj�����6�f���yce��v�����Pv3���IQ�N���5�>���)�n4n��Ssx��Įh/��ߚB9�}|�k��-�9�ol�Z�����wbw�fb���!uy��~��b8�I��9/ ��\��a������N���Qt�":�i���=�'��V�����>~�愛q�So��VĩSԎ���rV����Lع��ۣ���U��U�t�Q���n5�@W�1�l�Ӯua,������E��׺ϱNͣݕ��\G'F�8F�M��S?k�2�x:%.m�׼�xw�O|yA�����8��;Q��������b���^c�*��L�E��4l�-�����*���O���D;[շ�q5�s�K��6Z�3��f±ؗU�0�kU�*��y	������>!e"v��z&������@�v�~��m'@�R�\׹L�7�Hu�]�.N��pu�v�2�&Q�kE�5���I��\�Z�2���	�Q���mJOln�Q����>�餟'6�ko���?ٴ������?]�[�}�.�5�hn$g�y�Yrr�W�)ف]L�m��X��ݨ}{YvsP��@{����w��C��&��h��뎲t�mIg�35�}��+Go��KC(�W|�Y�U��N�����|9��BQ��[A�o.M\C�}e_W˰��N/��X����-T���eW�U+��[��\c{P�{{��-�"�
ۅ�
����;���ﭟ:�:{.���sL-�����t�p��Cv�HK���7r��;�O��	1�S�ts<��V�����7�	�u[c*]*�AO��ou-�4�ep��L�O]Z����;C�������le}.��D)���4'�!;���{ބK^���p�9�~�<���ri��B�'q0�3H����S�إB>��}5��u^F{bu��r U���=RɏQjv��~�i��;'?Q�fd��9�^){�8�?yoL���R����S�}��e�Ioi.��6zt��!L�t��7��]X���d�O,�\U+o��J.�ODz=�}_}_-}��_��S�;�:^�O��u����&��]�p�ϱ}�b�a-{ �wP�t.A[Aܗ�G��Gb��;�;�5F��f�J��K��Z�W=T:�w";P�x<�_�Ϯ?g���i �:.;9v%z�|\r#*���i�j{�ix��/[���K߳����V��E��]�{���" T��L*J1:���yQ���͡�: �*2�����b�T���_D���~5Bg�i��5#Q���FS�Mrp{�f���y�)k�F��M�W�y��Q1ظQ�͌t�y�*��m�}��PF�w��c}�ޛ>�0O��(��C�5��ƥ��C���r�{r����+�]�mSn^���{Q��@���@�O��>�Ϋ��g�C��7�
���yS;)���=��k�<��0���_T�4O�Ў�Ď��t�Ho�?^�ϛ��h��E	��G[|6
<u�c�}K.�,ޡ��t5;f0�kQ8��-����]�9�aR#����T"C8�v۸�$6�t]�\%J[2>�V�L�#��d�
�YqK]�H�#�S�e��y���II�1=�_Z�D}���ܷ4b�O�k{n!�j��<����}�oM	B��ƻ�Y_��A0G`;���^��O���VΩO-�k�5�u[��n��;��{����%����V���]��Ե�C/��o�-���P̫�y���YӮq:�.�dp%���ݎ]P��RM+�u��<c(,\e
�S��{݂��9��V���l`��sQ+r�'��ڑ�`��S\7��?e����@{���~R��R;@�C��DJy5�jܩ����/ۧb*i,����Mƻ
�5��l�[P��{,{+�-]U=֢]�ܸov�ի��է�&��CYU�Ș�:E�w4�M�y�m7s]٥c�U�%Nm㕫w^+��iKۈ��yG9\�ݛ���^m�pح�΄�b��S}����/���/i;�����鞌�	����L���E��+üB���`^\����^�,%�Kޜa��R�E(�+�g7�^kg��6�X`|����ɜٜs�����ϮbU.Y�(f���t�@I�&��GQ�F.�[i����Xn�\�k6h��X��U)N�򾯾�z�?Ju�����"�����̵o,�� �]v4�⧛���n�)�.�RA���w*�}��/+���~����A��:���墣U�`�{)֘!�m1n��=���,�;��ur��K�5��dë��x���qu�r���ˆ�˽��f:z�����L2���ʺV���ryӪR��V5��z��{�OO#�L.ې����cX��4���C���Ϲ��$��R^�[(�z�kn���w��:[h���{4i��MG���|_�1	w_R�O����gkzp���)��
W% E�X-ĺf�B�|�O(U�E{W<ɪb8�W)�ǙK��!.�wکl�r�m���Z�ϡr��A����M�;��4��y�f��Mu��**i�zv�歗����
B(�v�t6��;�G��сa1�V�.����.�K}�S�.382�Z��1
������4R��$�Y�k�v3�c�le����::�&3����Z�L]�jT���.��^�oP���ɀ�kT����Źp�8��*bɓ��F��v~�����ވ<��1/Զb}�?� �!>��a��q�¸���9�2�sL鵸䷬�~en�I�$8�E�����p�&�]�#k+8}��<ܣ��o��c"���U�*'��巩��I緓�㺢� ��gf��舾�m�T%f�X�o�f*�yQԴnjj/k��g%��̜eg.�Yq���m�jO��C��P��c2���l�}{�N#��L"J�ͬ�}d���x�2�
c���ۇ���]���C2������g�@�Iq���`�/��X����5%��35�}�{�2ﭿ0MI�a7ݯ�KI��OX�N���)Gx�[�⦚s�{⯪s��;f)M뵏�Q��dE^���tL�ϻ7%�-T���Cv��Ǻ��k�כ0�~�+޺E4Tg��uH���f?����w�UgN����+jGs�@�"F&3�-ᑨk Ҩ�Pξ�^��6��x�e�F�����m�ߛ���v�sf�x�/.`�B��,vtٯ�!s�J��;9)��k�:�\�km���H(4�f𚈇2Wj�=I����!�BN�^N�m���D���� ġg���o�6�������QC�H��}I�۽��wCj��֧�T�WK��n[z�g��:���.���=���d%���+(')�U{�la��]O_k-%��O�U�2�]3P�]��u<`�ә��;�A��kf��]��*��i&���;�����t�\��X(�P����������Ug	�%K!��#�I?G/���o�_�^`�
�S��ݍ�O��nЧ�1�9�ے�&�y������5Fk9�-�.����@��{�9��vD��"�Sٕ+�^-��B���r��YK:qh"v�l���j8;I���+|:�o�_�Ï9�i�XǪ�C΅wV9��*�����Kծ1�}G^�u)����:Ϊ�5������P�O�����Q5���/��\.��S�cH��G
�=����D{��,9o:}΁�[뭰j����k�E�6q���;~��_D�Y��Z*�gClI���
t�|��⮰�Kj%6�J�dQ��N+�j6��;�e�2���%0�睛HY�;:g����_}�u��2>������t �E������{B�l������Ϧ�(Jc�b��\(���:����Q�z�p�����[�N�R��"ml��!ʫ	�{�P�k��	s{C36uѸU�m;�!tԧ37��3��}Z�r����c�o� ��%�ZS���~^��p�卧�'�
o�u�U�l�>F��g�7��z�r�&yư�cf�U>O_�}���r�n$,�h0T	�ң'�ԝbSb0�ޤ�j�x:X·��PU
��)OƵ}�3�-����n$=���C�H�v@���k�; $�%��B��_9}�[����ʒ ��Π�ףK�&��d-�� 0JZ!k�媢w�������� Q���g=薬�{}G�۹L����r��h&{�Ss4s����#��ɧ��vN���6�r��^�Çl>��'�(t��9���j������O(;R��g�͆�ި�F�ٰP�Н}&��ѫ�2�,��^s)>��R���0)����]\�(-�Y{�rB��:�I��M��/gm��N^�gp�0�=5Y�}/[9�Xٔ���楩�C=�gd?3Ҳ��ڽ�iŻ���q��u�Y0����Ʀ��Ci���b
w�Iso`�;�u,�ti�ϰPt��zݪ�畸��H��Vv֦���r�Λ���cZ�V69ꝃqs�`�{ةj�*Wd�Ռ1Z�SniM����z�_�u�-��OL�7/��L�� �-�7Fﱖ� �ѺY�{�Ih��I���U|��{�����ip��F�Vǂ��Jj�j�)��!��%��#�)�M��Vf�-%<���5�_g%�&���|Wn!����W�Z�a�eR�Q����{���e@�`܄|��Y�Ѳ���ϖFP(!(�"����(m�z�C�s3���3�� F�!��j�l��A���e6����%C���q��@:%WGF�'WX«҈�n�#w�6u㣇BW���8��@��;�Rwu�G����=10��9I�3^,���_Z$<�*Hsw���R�F���s��h���>�rS	Lc����C��7����"�Ю[��}۹E.[�Ew�lő��k^AF�Y@�+n��ӻU�u�[`��i��V�S��}��Ch���A����>���v���Y����l�2��l2��)r�'Y���Į<췴��eHNw��Yd�ˬ���o)0��{��+����>kz�X�n^�u�4�۔�R,�zK�t��nk޸��If;ͩ��Gk�݈
�j���/I#[�Ck�d�����ַ2�Wy���G��r�ãU]Յ�=qp�ij*e	|�i��u�iw\9t)�*MJ�kb��bJ��̆�j��s�+1���`J0NQz8�+�Z3Fijn�l)�eY�qL����zʧ%(� �P�mJ{�*��E��Щ�;c͏vι�sD۫��-pl���ϕ��g�܊ʾ�Y���څ�R���+��ׇ�K�n��Ҭ���?Z82q����Po5�sm,�p���Y�#��I5����Wl<0�iT�x�n����/��Qt+jY�_ �\��c|8`u���k��5/V�=��+ߗ7ʖ��0Z:z�)�� �o T�.!�Dt�W}�b|�R�n�/(d3s��w��vN�ww�	<TΦ�n�b��輇�[��"6��F@�Y���sbn`,{ƶra�^s��m����z��Khn\2���FZ������`ǁJ��V
ݓ��urJ��(��P{�)�+j��K�5M(%�w/�Bwx��Ib
C����㷚��i���1 MIip��lf�ݡ]#�"[t���[��f-%<sR,����!�w5I���"qW���:b>�V%&sw����c��֪B��Ȩ�N�M�p�rBt��+-�8��� �S(�YC�Bruܵ+EDԸ��N-R�JS+P�Idr=s��ۑQʭw١;�U�����$U�.�)�$�hfL���^�Q�!]ɩ���VHG��p(��G"�NU�s<�"����E9�X��0��TD��Y.��q�w5����+H�\�#̠��f��B�(�Eun�Ы�:�+I9`����ͅ��½B*(��y!�B9\��z�q܍A�Swr���"��u.�AH^N.�.�TB�5sK���%��,�;��s�Y��H���:#�!EK-ݹ�H��D�VK*Caj�Z��"sB�9����'���T���d]L�Ԫr�m,���J�:!ܗRv�mwO
�\��U­g].r�{P�3�ȋ5ֵO$�E�W=�@#3�/Y9�rΙSKH�u��5S���/D*'9r��*J�"Ȣ�Ģ$�z�UGNɫ;���U�q4c�Z��_:&�z��3G��{�^>9�<�Ndn�&�jX��� �V�)kr��,��\�����~{~|�긚��'�T7�k�������DO!�-m@w;�y�;��[�]4���q�bTۉՓ_^v�M=�N���&��CYU���9�L�9�r�u�r[���V��En���_O-}��j/j��Խ��(�錭��n�G���b*��8�����^��Q6��J�����'pT��'�-��S�Bq�-�f��+�>�7Q�7�����V��xrU���=�
���a}ryOc�J���:�ͭ�k:�.�W1�E\��Q.r��|���b�6�E>��޵�A�L<�_7͋�I�����vu��;����j�SV�%�::�K��jFB�n�k�=�hW`K-��޿+�����3�%/��H�6w�G))*[�)V�t�V�X��ކ����M=�7�n�Lek@�neϣ2yMT3�C�Q%.����R�v��MO����B2{Sћ�����[�:��Y���Bycq�ǀ/;V��^�)멣q|$���>���t�U�+��P�X��Wo���=s��(X�9q�B����H�n��B�B�[nQ}z�b{h�&��g�Q�D�к0f7Rel�TS�Kܭ�I]��|�Z����0���}q��|�P�I�/c3|�}�nK>��*K��|��'���ز��w�½&��=�|g/:��)4e��vS̽��&(�?��&/ZP�M���L�D".Bs�{����4ƭ�v��ԤD�C������sW�/����a�OХ��;�X�k�N�l9��V�ښ�ud�ku��D'�jL8n1�q)��ԩ����Ji�uǞƄ���c�/"[ɫŵ���j�Zp�n1�w�ԊN-��ص1;�'7���l�-mD����߳����ߊ���{Rв>t��W�o�p�1�������}�t��ј�m�u-��:����;�'a.��f3�˞���Z��v���v��1�P_�n?�[��~��o��g�a��g�z�]�N!������M���>��u�����e�\A%A$l땠l�g3]�(� ���lZ�٠�N2�ڳ���y+G��Z�
x]]OFȍ: l���;��y�N^�Q�9,>�pVѰҔ�e��Wd��tw]'��XHF��y�^	4�޽�r>{R�� �}w32r�aɸ6~���K_��5�~��5�s�{�@AƗ���F�c,Lډ�ꏶ�%p6Z����[��SM9�f�jT�2�����hw92�-��+@و<�r�/��TB�J5��z�=6�f<���sYEGt��r�s|�B�Z��_II�u�T�T���=��� ee��V���Ʉ������-�6��}���(��c�x1�����{s�\\��S�.�Ʊ�_F�ΫleK���E]��^q��V8���^ߏ���ۄ�c�nZV�k��>�_[c*%�(8��i���V�i�c�5/^_�R�\u&�e�w1I���hfMu�`Ӊ��_��=��U��Z���~�[�Q��rQ˙���;��02:7/��;���-J�tJp6�zP����{m��?t�[M���4�#����zc���d�lV���ȱS\��F�9 S�,��S�Ow�-��7ӺR9Z�%". ӫ�l�	�7a�#	q���ee��
�MTVuCFcj��Y0M�$��t˼�z�U� �2�����<�N�U���H��ʉe�I%�&�uJrm�/�{���4ۍw�Su�C� Z��;uمc���)"m=����	��Z���u�'�<pv�<��f�5��]�1VN:s��G�x�3�A���;�{\�~I�+y��K�Z�Z}'\�Q��fl�gr1O/Z���~�v6�z�Z����ד��R�{��L�Y�ΌǩF^�{p�,�kz;��*u��6� >u79QS�{
���Û{���@������x2v���:γ�LvW�\�;���ꍥ_�\(�ÞlA|jm[���f�}�}�'���[U��`~�P���~[(KʬB����[��	8�[��n�!9�j����0������g�%�������eGxu��tQ?kgG�>���>e�8z�x�59�������.�ݼ�R��������T�QN��k��q�o��tڍ��x�x�YAf K��:�.�"�q]}Q����S���9݊���:�@�ʖ��KK]��)�ݝ_ %v%vx;SJ�u�j�ppv��=�k�HH���/il׿6C��71R��8�HH���TI3"x�b&;{���x��gm{1;���)�����~���AP�y
��tB��P��\|�>�O�L�\�z��{T�'xu#Z1�OR5B�����`��PZ��rꅼ2�&����Q�^�ʵ���ԄN���EL�B!OJ�CA�3ܝ)��;�V��~z[���m�t"�[��4���<a¨�R��#�:s�Z��WP3�4N]OGRp��R�o�t�Q��L���+��]1�m�AM�9�&/q��]�эr�?�Q�qN�=�������T���-���슑٢�o9�Z)�4�v`q[|��^TͩY�����{Q{V�{��*Q���-C \�o{�����Q��'�m��So�J��ڝE�&v0lz�O=���r�@��i�׷���1v:�y+X�����"�P�����b�zS����m��X�5���e���3*V��f�!��1�=�(g�^�.�܉��2��,}�[�0�9�7d�r�U�;X^�s*���_�\Z{/ 1/l��$7���a��V�dR�,����+��;�����\�O�}g��{��nY��b8h����2K��t
c�HcT�F�����}�n�û� �5�(�Wb��Ъ&+乱p�>���5�tڮd-��[{��z� ��T]9w����e�Wdjn��=�]�,�m>�u�l���RVZș��s��y�p����OuF�9W
�+�[��^8z�y=�6
��qU�S�W��KQ����މ�@r\�IK����T�j�Oq��D��dY�T��-o<����.!=I�q!g��ࢂLT���3S|�UJ��y=�YK��`W{��t���[%���Xڶ��j�\m]8���w]�����n.+-�5�����g5���l^�K�i�����j�f;F=nEgG=��Nv[�}���%�\2�8v���aJ<�FX5pI�S���<�\���<.��O����g��<꧹��$Æ�qW��Me���� �w4Cv2~m@w?���&����&����j���n�~�i���}S��3ڷ����N+�c+�7c���C�*���W�q�}�ң�mkʳIx�x���/���an�9*�Z���9J5wBl9+�.n	�t��oE��K�Qf#��c4&�1F�����5�x���)U^��AyF���yA�,S��dhu)���s!Wxj�X�*��ɾ}�qo�ix%�\����L���8.�ѯ����n!=��vn�����bR�c�4l�x9ܰ����y�vK�MU���Z��v��]#Y�eA~��n~(K�.@�el���o�N����:Ȭ|�M��X�ӭ�}�Yvr���igTR��֗͢�͕��v�`u�])����5�jkH׽�K���V;����fۧ�X�+6�Fur��l�\�l�c��܊i�1ή�*]�^C��	t��'�����g�̰��`��(ͩ���z�/2.��FR��K��2� u�o�9O:�+��f
�<�<��^tG-��ά�f��g�4b�K�����kn1�ڋ|���w����S��{%ӷ�͓:���k6�s�����\CZ�f�ί����Q!w}�{v �. �j�g4������'�ż�HN�'
x�K2-Ե֕��xȧeY�(�֯c-��5�[���8�m�ͮ�e9\���;�kr�tw
p]��a��� �oW3�-EƶW=���cyvQY��j��`���,�ǉ�\��t�\��7�
������]�9�|��ۖ��;��EE�2�]2GYݻ)*�����īb�����E���Z�]���$Ҹe�v12�9��r�J�)o,�	̇�MF�z�}�=+rkw��3c�3�5��%k�S�G�c]�w�	��v�N�X[��)��v�������M�)�M]�v"�m��m�Bn5�7Z�C�Z�t�{0o:�7y;�uuUp���y9����w�K��^'�����Ѭ�:`Z�Y�62T���=�8�c�A*qo*v��������Kۅ�5��s�{����(mA�<�Y.������U�;[r�e�j���"�o,\�wIX�8�/rYKU�mK�>��}�T<r��ʁ)���{
<����gwW:���rA���w5}ѝgj)�ʂ�`�=������X��͜ɵ&(lw1���Q�-)z�Vk*��*�w%p�N�B-�wx|/-1}�f��ղ ���H�5�v.ҦF z�0�-�n������h��U*eN��Cw��8] �,��p�j�9�ӊ��3Wp�>2c�*�s���w�s�Mj�r���.�J���i�;M\:��犣:��h���,)��������!٢�z����Q���x˄��I����T��ʿ,� Z�n�q�Y�����{*�R�+U4���������4���q!������FM�t(�y�p����@Iu�]Aҥ��w�k]��3��U����K5��v��1��R�@��7�S��%����r寧���q�힖�վ��Y.�r�&�kF,�ȅ1�.�(���/����w���r�q��B �e�o�mH�N8�o =�P�Ȣ���]�4=����g��Z�3@�����7�4�OF�|�2���xÅQ�P��Gj�WױT��{�Ȭn�S.md�n���A��vL��k�Q�艎Cak[^�n���J�/���y�"�Q�Rzas�6��A�=�};MG;ʆ��w�ú��Ձ_mY�����t�G�y^V{���P��zMK���>x�����l�|~{k�=~�;���`�g%Qj9 yF,���l\��������|u��$鰦n�q+x��n4#�ݷQu۠SRob\��j��ԒvBp�Ͼ���7'v�8��?-;V����3sb0(�z�^��ir$_'&.l�����C25~����l�����Uu�V7�vS�R�T'��5�s��"Eg���Q���V��xs��������k��P�o_��61�>SӹUz>�i�	:1_��z:4P�	�3�5r�:��\�	q����ca.l'I����[���v��r��8Cso�����%8�	dmt5Zፊ�����z{�}��..��sϖ�o�Dzh	@�I�ڧ*�V�X��ކ���ڤ��==��y��-c���Q�qoz�1�9Q�{��2w4}�ǽf�]�b�U�t���B ��=��\1�o�0�ޟ��b�]WԸ�7������t�b���l���N3��{-���D]��:hʪ�!j��o�BK�a���S�KXޢ�V���Q�4��k�X'_3�J�M��%V�<�fD�$�4֫����ٽL\/+$i�_b����/��<Y�Lv��Y
�f�t���}���h�ql���ۀ���uT.���آ�+'x�z�g1}���� c�cJ��ˆ����ӝ��M�Mɟf�nub���k�EJ��k0�	d�b{:9f�=W��R�t�ެ;�!�dL�:V[���/z��絳V�e^=����֌U�1E!"����:qv��J[���E_qMq�u��Z�e4��%��<I�R��S��u;�h��̀.������A��f�1�\�>�hqV>���)��^J��M>�Su��H߬�@6hN��u+MmYa�cV�[����NmZ�^��I��!�Z%u�M�o�hKC�����!�x�k��屛��]���V ����*b�'��Փ�ۓ��1��:͆�5�*"括�E�E���b�x2MyN`z+�=.Aox�_0���	Ǝ<F�X�릵�et�ޮ�!+P�Xr�(��{���Zw0��Ɩ/y�}���Mn�l�Y�C�͖�qsf*��z�p:��1��ș��O(.�������y����H��9�>͎�Θn�t����G4�yKL�o���zE ^g).���ұ�5[�mh�8Ql�;�eu*z�V��q�r�� �v����e�ge��Rg���4���ۡ}[n���fQ�A��Feq�[�v-q�)չ.!��(_��]iZ�vN�oF
�à^<�s)�5WN�5�'Y�e���q����f�Q��"�w��n��P.�������\�I/��
���� ����vK*�˫�ׄ�X�C3 ���-�~�"�|�s�4c@���k�WN�+z�ƱhSv�-:�j����c@����;�-m�}:���z�i�U����a�q���2�e���X4��y*N}��kL�зm�f��ipN�5}y����VBJ��;�e��tv-�X���7Ӟf6+��8/-���{��0�o�-Z8������wXF��6�ڒ��p�8�=t�H�pʺX��r�bR���K6�9�iE���DC^|�]'���:�8n�}�\ �B�����Vm�bwG�%����|2�3��T��G*ŎL�
=��9R��q���V"��j��[��7�s�:��.U�p9-��i�N���t���x/��5-��h]v��Ҧn�r+H� Ĩ�wu��7��ek�T���JMet7�;�CW#\Wt[�Vp%��`�.\:�QM}�m@顣6;�g����h��Ҋ�µ���d�y1�=����8Z�N�����-�q�NqYY�s����`�in�i�E���iiʙw��4�N��ڔa9��7��su(=��U.u��t�v̋n���ð��Ab�(�v�dc`����_0j�NKL�S�6�Yn�R��lJ��#����:��*���Rxa�2�D�wE��2�]�ʽ�(�DJ{�Q�;��&)e{��V�$=tr�D�\w��[R��֐�-5"ꤕ�6j������y�A�*��h�"Tێ룊!Y��']w'"��Ey�����i.⚓�l��E�	�AKL*"3
�R�HWP�M��5�U':g�Lq��yz�Nsqg���%�t��5�,�CKB���G�����I���9�uwi�T��ڒ�s��mu���X�\4�T��bFbh�D�R�QJQbru/-M�F�l-J��PB���hn�8�P�E��ܯ*u��m�ʽ�IV,�=�4�RNTi��ԋ�p�C��1�s�J���uq��疙�̙�͚���EQg�Eiܹ{�T	��@�S����y�ib�q��h�l�P��Qݻ��ӑt�V�B]��wrT��F�V�rP��&��V��#f�գo�ػ��]����|:+����x0'Ǽ��֙y�h���Ã:MGB�eG���9%���xr���&�TK�P:B�TmH���*�,6�(3��S���V��K���|��+�AFw��;u�2V��[�8�R�C�OGһ'�>��:�>�I&7�UNF�᷵�V8�԰;J�t�����\�V�w;�w���I��١�I�n�Z��t��i'���Ds����-TK̨�Z�yd�Ѹ����Qİ^n)ł����1�f�yO�[����yV|���>+�mICuVJ���s�s�<�yV9�s�_^�;����q�>��ٮ���3* �팋�4wڝ�ι��e.sr���Q6�����ｽ�g�#^|�tv�{���fRIu!{o!!��>ꉹʏ��}��pPy���'��w@�=�=ؘ��f����n^Ϳ�l����*�U�iBQ���ډ�ʭx��y��u|��o�����3�����Q��X�g ���Gh�H����bX��yKkK��{X�u�DT�׃aDe��\/�����?q�{u�Ӏ>���Mk��z��+p��ּ,�;�y���R�|��E#�*V�W�.-�*3u4�혦���;�]N!֮�m��@ك�~�I}[J
�Z�qp���9�ޮj;���*��9e�O��{jo�����l�P`>URo`�.P�g���kǢ��󬩨|�����8{o�s�n�+��K�2�JY	���SK���'7ԩ���騇/��ֻ#\gTE�2��W�̜�m�۴�3\嘇�Y�0B�	u�×-}����9�r���U�-����L��᧹��/�d>�v@�O-��Z��%Q��T$Ҷ_6��[G��z�k&y�U �=܀��Y���4��}+rj7y��5�׉����_6�f��cZ5�FQz��q�B(w�H�=]��w�\��o�g ���S5����W���\���mI�I���}�Sz茎C������N��S.��HjR���G��$����f�z�6�ޠ�{�ix��K�ɍ�ҕ��en��0�]��ՙ�n^�Q�m-D�n>�|���,�缇W��tP<��,9������1�@S\c�X�d2���%\}9Lɚ�i�ƴ��|�Lx+;����&<��&�ԐPi|B���(.�әao3.|���p��kZQI3;5�"Yfc3�f=�ݴ��Ѥ���{�R��k�k>}Gi�Vq��gF�{\�=��9���c;�fGJ����2��QX���K�|��#oE�����Oz��)�Y�@�|b��Qtg��r���^}�y=������L� 
-u��]�ggQ݊c��*�o\K���G)��Gj'�3/e�)��a�O��Ux�C�i~��[��g��,(Z�:�3��ڷ��!]8T���*1����z{�����Y����y�YV�I7o)�_M[�����JeD-on���{_&��)��𼸙i�.��{�Nhr�,l0�O�%��*[5
S���k�]sG��C�Sb��o4Y��8Y�7�f�%��|W�h�}]�T-}4��NS��*�_Lͬ�UR�����m���H�wˤ0~������r�X`�B��A�|v_'Mt&f�-4`V��V�]Gm;ݎo���|��v�0X���Fo���U�G�88�a�� � d�����ȓ���oU�V��s�V,ӝe^9|�j;� P#ou'/]��u婰�7�����jV��$�wWBl��Ԯ�S��ѓ^ɄV�2r~g5�p&�6�j
c�.��O�]ʼ����Q��=�z�ޙ-�y;[�H�j!��öq0�	�Gj s��)n����ͱ|���MO,�כ�èO���=��q:胖OM��u�s�ɯ`~T�z�[l�o�{�4�'�=��8F�pv�{^Զ*�t:�Q'�^}I�ʳ��=���ێ/>�?-��>5�IV�O���&�9R�)T��G�s9"���
{s*�{��a��t҆m��v����s�9�|�N8{�Q++��oW��V��T��1t�Q3[��N�]p;�^$�<�N��kw�����OP�3-���|�����f,�r��wh�Q	sb��}j�w޹�gY�N�NI���R��0s���Oum(J�l�q���\Bi���n�|ab���.�q<��0u+�f���wk�@�f��v�5:�6��Ό5(o-���n��a�)�8m]
S)�0N0J��1��Z��8��Q��:%,���|+-rN�<��&樸!p�S���*C's͔��q�j���d��\ۧQ��'����=Q�����uZߔ�q��e��7��^g��u���F�wA�������̊���yÂF~gG�lY��PA�%�y��ڔU?�	��8{Qo�St݊	}��A���.��}<�A��t��Qr;-��zY}���N/{�lc�^p�DU�o
�f����{rF!*D^�pZ�owZ����kY�{��c+�t�"ͫ{{�+�y[vِS�	]�Q/^_�qĵ�_Q������ J�0���Ñ�~�-��m���X7'=&a+��b��z���j�S��vG���q��>V 8zRΥg/�����jdyOî0
���S�z�A�TTD��ӑEx�\Fm��|����G�}R�Dắ0��r#=r}���z�g����e�5
|J�p>7g��n������H�.����u����As��?^\<���9�@zMǶ�»>~찇��o�j���vX���b���s�y�55�i�^0[���"]�l��4���e�4����|k�E�yL���R�G2*7�X��4K�kU>T�Q����q9Dpt
��6�7�r�w��md�ջ_5[zT`��d�{]�ahQ[�2��Lۧ07D�����X��:�Sv"�qT���~;<�-���W�s^�	�'|S�+������7������mtz�E#���V*[h��.PWS�t	r���L
����._���]o�ȇ�ݟy^��#��	���=��.�B}6X�s��	�>Y5��]�6���_Ҽ��c�O���~S~����ON=���!�}{^����Y�)\A�xA�>�Gi�8T<D���k�D��ˎ�zW��ޝ�����]��^ZmH��.x�Ƥ��2�џ#}r�K"�+�W:��Zc{+�Б3����iϽ�|}�����NG�ׇd:�A���.��OTL�$yT8bw%_�^���+ގ��\��]O��l4��s�O���=y�p�"=5�>ρ�Y�p@�� �Q�3>�~ݼ�S���@�(e��x�z�HU��hhϼ�����Hү=냳�a���ϗ��gW�b}b�h��@ݨ2H>�I�)�
XV�և�y��޿~��a,y�߷O&wB�x)��ǫk?U1�	b�&:%z���|}��Z�H�m������bI�Xǫ�r����<�ɽ������F���o���Qf�X=�~�W��W�C��=B�f>��U�<�Y�� GwI3"r�"ʛָa�M����U�qW;�S� a��-c���N�Ơ��H��iѰ�WAX��^�a�x�B'\�1��(���ww)Wj�]JB=D�|=:7����.'�쉷3�!�pzH�}^�t_��^3y�}{D�{�w�3��Њ���{�jM�ޤ�z� �dXC�`�)�3���񿠩�R��Ve��Y�9�;�R�m�z�Շ(�=�|o�T;M]��}�d��P��e��&M)�T��;���_{Y0:��_z-�0���8΋����_ٴ��r��i���c�K��l�O[���6d�J�u���hQ[~g�K�ٌ�Z:���B�\Ogu1���u��}��O���)����=��y��P��d=)�+�	ǽ ��1Q�R��ʽ��g��
�X	���u�|T�͜r;��z�烘��5LØ��UHN6�/s�o�uM/��( 6�a�鸞����<�fw���k������o��?:Ag���b=Z�L%� ��7
��O�Q&d�g��Z���`W(;���6ܯv�.��Z��^�aB7ǅ�I'�e{�P,/�UX�*��ުOz*ezb�j���ޫ;��W��������z�ǻ�#l�2��^�=����l˘eQ��gs k��xȽ��B��Ebp:���HW�����3GV�X��nG69��`�k�$s�-|��L�9��6hS���Y�r��ʮ.��¶s�ٔ�F.�*;"����8*��nD���ipR72��:��bJ�6:�Nr:�W��_��!�cr=�|y��{Vo�M����2��-�Ϯ�?@�<k�}QX$Y���-]A�÷�(_Ο�Fy�y�/���f/)���^���a�|�\�~�\{��DU�p'��q /|CE����g�C���֎홼�'�Z���&��!���sޒ2}Tķ2\� ��>�&[����+ћ�<z7����m�M'CѸ}�£o�{���9��. ��A���z�׌�%�U%��=$zf�\�`{�}me�"��=�^�Ru��}���m_��{��O�A���XC�d��r禥R�����=����l*�3>�qs`����E9Zj�S�iz���+�16�fM��O�w���[�[��FL�����D�K��IX�;,���⍴s�M_ٴ�r���'��!̃�b���Ȫ�����H�i���s �:|Jھ��7�
�����l�1�/���ݚ�r�5�-p���k'�z9n��yPfo�}���3�P業�+�*�yKw��ڰ4;��j.s�=uL���	Ŋ���mqѥ�R��IE��������o������P0kX8]݆5a|۾�-dv&�&��D'�L�vpĨ�Z�����~\�;8&f�<�#�N�!�	)*o�e&���ɠ]��[\��s���Ѿ�n��-��y][��ˈ����ha�W�k�a�g�G�~�2}U�%9��)qwQ=q���o'$���;q2��Ʌ���}��9���^�/s2N�Y�A�p+�wϥ�/�9����%�y������4>����"Cz��V��i�ڵ�|C�	�q*���J���,���6�/��~+�����Y�p��7ҬU�{<�,��:W��CI���ʀg�O�޷A��:hy��_����r������v�ïu��A}�W��yz+P��)��,(w�Z�]-Ź7^����w�z6�<fO}�Uf_�(@H�r�}�[����\�i�$�a���P���Yw�2Z�^,g�;��5�ΞsSw�^�V�i�����do�q���6�޻��@6K�r �5�������!�<}��Ì�⪷�d{^���\Uǫ֑�9ⴧ�U�����^�fm̂�D(#�����fح��.���S��e�e�p�R!׭�9��\Oi7޸;q^���vz���m�
*�qOo�b|h��T����* �yM�s�;���;�j�u������Y�9�\a��fv��ɼ��[2�v{�W;��"�^�fV�1m��P���i<����NC2�%tsz�j�JVs7n�A���D,M�䶬	;����#1q�J���\�W�7:r.��������2QϘ
�g9���%� 5b�K]\7*JUa�ձ�ic�6<R_pI�ǔV�X-r� yV�N��=�&c޸�b�_W���it��;#��UH��e�@�#��/�3܈�7�K������+���K'���\����9Ex�^m��:0�����Sc;��~�Bw�=�y�Pn!��g����\���Z����w^�Ӧ���d�V�<Q>��ÜS+O�o.7�r5�����mׅvD?vX���L��O�F���'F���4n�|{�1V�/1~���ۏ].'�����uG����i���)�]��ǿ��n<q����7������6����qr���P6tu�S�t\u�w5S�|�<2%��x�_����6����5_��䫋j�y������,ʖm��fc�W�|�Y5���X6�]�E���x��@��R���*B�>hߢ=uø�G����ʞ7|JWa�=P��U#�������͵���y�Ԯ��^�\`L���Nv��ף�hx,�����#��$�!x�2��g�-2aʺ��Ū E0��.�p&����W��>>��\?)�����7H5�6Kg�'����ު>6���ۿPV�������v��m���+��\�����0P7h��}��x�T)7LE��G|;*^�VԾ����|$���4���t
D���Yd�v��u�Ym-�q��O�����&W3hc�k)u՜2���sÏ2��p�m��e4wY�5�4���cf#��h3H���6�����:�
�v���}2w{_x����`M�i�i��	��vrM,��*���yDPVq���ʊ3�8��Yn��i�ҫ)n)�����6h}{����M�	��wO�"1��ˡg\�ky��ʡ'`�9Z(^���R[N�n���;R(�7�)�(q�	��aYv�J�Ԑ�1��L���F�Ճ7G;�-d�u 2t�[k���Z�ݘ[�D�0�;�qeh|�cF�u����ǳ
����z5�2�Ry@�J����/�g0rj�F,g�ۮaΗ��չw�j�6���.%; h���ȉ(��	���6��6\�w% %y�X9B�x�خיLq�]��$���Ջ�+�d���6����5}�x")ZS�-)J�X�۲�:9������▊�x�ǝWX���J�L��L��f��J� 仫�DJX"s_l�2W ��E<אtښ�<)�2�;räSSr'�0���
.�p*cR�E˹�M�Sif�521*��(T�6-6�v�jB�6�f��S+�r�D�D�t9�^��d7���; � \�M�h'c��$��`�c42��$mL��
gk�xęʻ�:��v�o	өěX���ame�,˾������E��r�A������W}���8�H0�OM�&�%F5@�sF�ڳаn�ǽ�5��,v�)@��'� $�C+����Z�����8س0Y����ҭA��
Wz&Jc������G*�+D�jG��
�XS7z��D30�(ա֟>�:��kZXE
km��:�����vs�����Vᥳp�|�+���Z�t�[q`{�匨w�s�v�3^՗��a:��4�	����*(;b��	ɨ<�u�j Y������T�&�س��p�+�$"��<�u�nԖ5�����x$Ԉ�n�6��$VVg �u� "`��W��sVov��2��"Omb�Auu�e��hƤ�ظbz/�m�5x)��]eF��G7�ְ�܎ΛCy���bc�e�,8�^��vl�*�G��՜Y׼0=��A�F*�E+/mC��:k�c@9��Vs�n�H;�������h��N�v��E-�߯,)!�k;d��t��qÖ�&zJoK�Z���'�a��@5��(��Q��-^�L�tn�c�8ԭ�gc����È=��}.PҘ]�Rj�XM�Q
�|���S*G{��"m�fS/2�K��JJ�.�x���tڃ �{G�J	�;[	9�I�ED�}�<bfW]3���DbǦ�7�)�˝"�`���56��j|q��+�s`���t>"�1B䘲t�򺻡��{��J�ä��n8�d�����(��'5,�T�X�"�Q�髚�IG��ٝR0�"�0�$�H�'��&�HX�L�%��wne���h^��(�D��x9u��:���0�(�*�T$�Jպ^�r��*�LfEU�i�RV([�U��%i��D*�I9.u[�QE��bgNp���ự7$�D(�hu��H`��t��+1ݸ]�l�U��Ad��֩���H�U���	Lͮ��
)�Y'-+GG-ɚ"�Ī��{�e���4Еe9����ꉊ����8�Q(���*�bV*QZ�)i�4��fV�̒6����X�*mݹn�TN�!jr.G�x�m�pIK�*.�)�R���UCS���T��gRB@���I�={��0zƵ<0f�d�2�qy2��s�%I���hjv�e��5�<ʴ�Z,�퓚Y;���f�����e�����\��V�SK��*��׏���^���V�o�x����Mg���Y"�˩;vo�lV��#�%���S�jm��_��_�
��W��޶���iW�����{ϼ��D���z���%�~�rY�� s�2��H��^S���z��G������_�^ӑ�����w=U�+����q>�u��>�Q:̖j!��<LL�WQ���>܀��k$hۜ��|7��]C�]WܥMj�u�=�׉�N�oޭ�}~ț���eX27�	{��n��w��ꑰ�;)~�ů�踟EaOD���_��G��@�=> o�u�9�|��� K�ؙ�{tl��z��-��+�+�<�Ѹ]/�����ΪM��L�?z��`uC.:}�%eN��&���\���+���w-�{C��u/N�����Y���+ˇ���ь�~����Ϡc>�Q���b~�����oF���8'K���&<�֏\T�N��V���=q�w��!��dgϽC�/D���	߫�����پ@�`��yދٕ8n4�wo�0�|'tÜ�q�:�uu0����_3K�������9h!ng1ָ�޼8��ɮUzt�V��]y�E������s��!z£ՎP,�6�F����MU�dSu3
].��+�HO=�[�Dn�h�k�|�6��#�5ǵ��h���H:n,z�u*K�2kT��;ҕ(�FW�����XH�ym!q��#.���a�SVUi���~%Z����p�����ŏ��� {��Y�Kޓ����~t�ϼ�и�S�z��C7闆��T+�\_��_N�s������>��8z\c}^%��}�=���W�7�O˽eL�������]�1i�u�����H~�3��3�1}j��nz�<��7���9�����w�5���z�V+e	����K�f'^xe^I�`O��b�U!}w^�.�Ю}����=Ln{����ͨ%��9#��wV.������@�>,q%i��}-��S���
_��叼�nf�i�Wn�UJ�z��{�4��RMǽ~����PȁʌÁ0[�$⯠*���]���e;�V��Ԥo��7�1Sފ��{���yߟ�'=�#;���p�K��@H�"��T��c��.u��)S^�������f�#q�B����m��}�Ϻ���נ\���Y$����7/u�������Le�cex�M�!W:΍��>f���Tu�ڿI�z|�������:�*�$glGrb�T�B�/<G�;1f*�b�ιJ`W*��BZ��(/9ά��9��A�7�AO��6�o7��7��9K�m��S���g�b��e�ǤӔ�vH��ѭ���u�!��w���OE�*��ިE�L;k�+���J�·R�벭S T��xen�Or��`�eϠ��w�
��<��J�W��|n���w&-��2}���ni��=^�<K�6��b���.<ß�:Qk�dq�%��]�m��֢ki��Wxϓ�܅0+}�]z��S�o3].8��>�~�{��P��T�]>%Pɇ�wL.�V鸥/�����8Nv����.eTR�ՊV�;�	���nC2�h:��?uXWs"�e���ڇq��h��9�;/&Z���2ǯ	Gн-�η~.��Js�R���'�ݹ���䜸��:v��xkSÌc�{��:�;m��+*�d��G��|�<�$�x�r!���c�K>�GE�΄��u�����@��� |Y~��ʁ3î�Q�f�C�p���~�^>>���X�\wuz�\��"��/Gr��>ʟ�>%+�,e<X�|��n�.8���x�W��[�&-�Y�;����h߾����h�C[R���OQ�~ �c"�R7�u�O!���?{f����Y���RS��<�z7��߭�q�u���rY�x��Á'ʡ��e��)mݼ��23�v���ϛ��H3��\��ܪ9�&g��ղ��]{n9,���$�@������J�3P׷�vZ�ut�+�E�ηP؞/ۂ�1����<�xǸu�\�#�	>���9u�īm#���w)YZږ�:T2��j�Á*��Xľ��O
�u�q�� �e�ə)��Ԭ��{�~�_����:������Dmǽw��l�P��k��J��4U'�~�5���@:�s�E׺����>�L���FY�Yu�f�̂�h��2O��^DfX�J�[وC��d�僐�C-�R>u�l�Gޝ��;��M����v�s�H�nm��
��#���_*���D�IMM�����#>����ڿ2=>V|gJ�ry�L�����y�U#҉~Q�+�n�m���	�j������7E����ǚtG����%.��nߒ��\��#+�=�u�}>|�� ~������ �zl�*��;Ex�j���/��}��ۮX���/��m��y�ɸ��Ϳ_����_{.A�>%@�����ǼDp�2���IY��O�����^-�/���\,o�h�k��7ۯ
�~�#������
}GN<��>��v������3a]{����o:�ǲ\״�~�����z�߯x��~�z��X�ӹ�3w&g�,ў?���gng�����rN��J�N�j�^�dx/�D:�g���Oަ��{&fՎ��Vd�(�
M��
���YN�dWG�3/9�C��Z6T')�� 83oL�J������B�n=咈��3�2�d�KX
�a{����]s��Xam����Ώ�n��':Z��Ze��A��̚���jt3:F��l����_��ʝ6�'v����O�b�+&��r��B�l缎�q�w�ٵ�t�������Hw~�CU����R�0���z��z��t}W��f:��t�ݴ�D�E���VE��{��~�<��]��%�5�#��<j"J�2�=���v�|x�޿�az��ϠO�;�qޟa^�>>��\?)������e��%Ӟ��Q1�5��g�}��yIK`{��u3�L\u�K*�Ф�{O�����o�x���W��Mg����u�
>�F�ks�1��X(� fx�C�@-�C-]?�����W�}�h����%���a#�R���6gb�/���T�8�P@�F@s ��E���2��>���#��lUVl�fY^��On'���@\��7=��3޸:n+�뉶d�P���@�&&%z����ہT7�=�8?z�9�m5thO�`�������|ǧG����Zϯ���������FD��QY&�<�CMfVU쾉�x���?\6n<�����Mǽ�@�>� ;�`e������2�i�i����w�y�ވ����`N�Q�﹇�O��7k��Y���L�E_k2���]W�5fc|Of���AWN�GH��d��-1�b��Ǳ%7 �p���:�҈n���n��m��h��n�ˍ���g%H�����ǍT�D�'��'2����gh�˧�m/mǱ��ɸ�/�ɸ��P��e�O�d���eeghs����[�.|rpm�s��T�:'�>ٴ��+ˇ����~����l���3ziT<�}�B;�'ӧ�"���(�C&�Z�O��n���<�:�G�s�9�|�baV:��j~?T���^O����f����P�$FT�A!^U���?��N� X�|�~��*S�ۋ����r��/W����:���-�6�d^D)�;�ò<����=;�~�����8t����v=�N�*@
zݐW�{�_��|�!��<�нS�z�|Js/�=uޓ1��33�=�33o+�W��VUx߮T��@w}^&�nW��~�\?ߌ4�}?.��hD�����k����!̓���6�L�W2���[�._��`��,�9���z�ǻn�ߦ3�7�#�W!N�Cl�E��z��$�R���9v�=�xh���1��������P+��)�~6ymE��oxǰ\�j�J�,	�R$TKjr-]A��y�4�嶶�%���Vx�ӕ�a�(���c[������k��îߣ~[f��aD{��u(�5��4�5��۽��ڤZ#x#�fvГsScmH9�}ӱgV�[Rce��v�%L9���;sy�~n�T��ٽa��K��������@�T��=�֚W�� ��R#Ůo�Mw{��ǲ��w�iW�@����B���"*��8[�&�	^+&	>��R�Yt�e-��QR=g�|�+��h(��y��C���z�ۯ]�7�9��SD�q��I��Z�d�tb��Y��j<���*:���s�;��:}ՠ���@���_�ۙ%��>)��dDf��Ț۾�s�D�T�]O����/��|�G6��T{��O����`o��w���73�7��e7~�Htnr|fa(Sc%�xк��5k��K�G�����&W�n�rU��N�	n�R�O�Q���$�"��0���W��މg�j�X��+�Iܴo���
O�JS�jG"2�#��C�7�O�����(w�d��=av���
};�Qz}�w�o������G��[9��}#G���C<��>��3~ڱ��ȇ�2�e�v���F����!{�50j�V�q=�{�	�>���:rKf�:��3�%9�֧��u����rNq�8:��:��{T#Y/�>[~���V��p��[%���w�3�,��s�����;�f"zwS�@�6��ȯ��P;m���ɲ�֧�pf�qY�km�.��t�����o�Z�݀?�2�K�ۨ8q�э�{�Y��hs�O�w�fm���0i�V��b���v\����I]aAnHT�"��<�[4>�tn��mEl+��7�u��jfǾ�Iӷ3�&xz�]\�)�;,c]����`�C�L��|V�<3݃v��BP{����f/VT񿬲R�2�T<X��g���n�/ t�����+��5���IV�;+Ѐ�g�Η�����e�Z��ۇ�"V���yC'��-�����}Ӷ�k�*�\-�����I��h�z�=������c�\ܠ���I[�p&�C�]���}�j��66��WU�޷�n��Ny�����7�Dm�{�~�D�@�?_� }t����v��w��ۘ�}��M"������+�;���*�޲6�V̝�^�1���������Gނ4�L��=��l�d#-�ʐX��ُ��.��؈P�96+`,�{�����.3���������#�V�2���|o�>'9�+a��� 'u�U���jT��O�>���'�=Q�+޿\M�>���5b{TK��d���cΣ̪�u�P��3��ԨEK"ǽ~����σ��*!��)d�!����}[�z�s����~|��>	=+�8���Ԙ7.�*����q�̣�Rݡ��s{���d����7X�x8���׽٧#�B�fAQҎYX�_�J<�{>�n��l���6�������ȓ�-%�	[�1.mJi�����Z^5��Y#sYS�Tw���i�U߿m�c󫓏����8��q�ːiO�P0>7^1��r�R��!~�N ����e=3�q\TG)|s��7�9���߶�»!����>ɜ�0��j"S���}��0���:䡛
��<r7���gZ��f}�9?Ew��+���#�OY����Fzְ7�߫O�G�6�;;s?�ꁳ���:��N(�L
�����t���OޫU�ǔ�<�RA���ＯQ���Ӱ��ݳ0��ck&��T���$
��Ϡ���efϔ���������K�N=t�q~�A}�*x��)w�W���ח䡽�]��j�L�ֶ��<�.|?U�Y�W�=��c��Hxr�^Z�Ԏ���O�J���8�f%�w������Q��G�\	f�|����W��O��#}p��=n�;"e��K�''O �3��'z�O�������u2��T̢�M
K���ȟ���G�^y\>յS˽���yдj�]�Ӱ ��2��
P5 ��C-]?W�
Q����#Ͻm���bd,��P����=��>~[C�`�أa���y�SN冶�6f���9�Q$�'������+�ɛ8�LH�x�#,��A��h{V�g����ia��f�Pw8��B.��ի\�.�f#'M�5k{�<����+��u�Ojz"�w� \�iA�A�=?�IJ����o�hp����k!O���b�.�s\EϘ���v��.'=ꃇ��~���d�P���@�&&%z���|}���l��\���b�z7=�vH�~�����R'�=:<M����.'�쉸s>�@���C�^�x�@�b̋U�����+�FF��������M_�߽�@����9�7�T��6�xU]02�վ��C�z�>�}'DKu��"���mt�6����ΪJ��/�ɷ�P��:��~��~ӕy�B����F�\���s'�zcN��:���i�q��*�6�����O�\ak�W���e�:�F���b:{5���k�w�PVf���Ī�0������tZ�\OdwS����xu�Ϭʒ���]oEG".����T9�{����=�-fT�Љ��0��b���K���'�һΜ�v^ =���ϧ���q:�z_���>�s*F#�s6��Gʡ����=�;>��=]�׾/{C݅�g�3�'�i�+�vEįR����3�+��H,��B�T䞻���}YZ�^����)����s�._	���rs�o�U�ю�5P0o�������G0<͚]�=4!�I���� �#�� w'�74h��:�QO��M:`XA`|�"�Q�w9�始��&+z�Z�i��˺��ǩ���;��΂���sq`R�Y*JmwR�9E;A���s82��a��nf7�{Xt<ȵ������D&������[�.���o�X^��
�d%]Vr�N
uzs|�F�V]m�
V��&�����{"�#����z�\�ӭM*�p��V�Z�܂θ�]��(;Xqo>�g��,�;�k�Zr�t2���q_S*����lh�f����m��0#���\��wa�j�5(4n�qv��0͘�0��v�sc1Q\�����5\��3��hV�Qo7�35����\������Y��񈞞��SY{�p���S:���;1��D��d,	��Rw�aʾ�
���	����G�V��
u�Y\�T�tZ�����V��Os��mċ���� ��{�5��b�Ar��\z��!8�6S�ݤ��@���Kk��W�q�Us���P�ֺ��@�����JG	��BR��w�G=օ�Ac������WT<
ٓ&H3��*x7a/��c������/絽��+t��	=sB+��T厝\�9j�U(�3y�Ԧ20)�8�ۑu3�z�J�[�u�NN���3����)I-�w!5�4��|��,��ˁ��N�zV�ak�܌v�3��1�UbX9[ǕX��y��^�B��㦙(Q��jہMݶ)���5� �[hl�<�f`��w����X{^�{�[iΩ@vQ����]d�ۙ��J�W��n=�8��3��:�<Cqkvu�m%�t��}���~�;��T�Nw+�^7�:t�zf��_E)j�\��$4�R���}�����Z�s�>�!��;����/�UH
zw�N#ή�[�n;[�%^��o�.3S�fn3
Y�UY+�Er-��ev�*��Ǩ7���-n�#53��Un�ג�pf�ٲ�V1���*����B�[�Y"�#d�����uc;���gRL�V�i�wu%k���O[b�YѴ3��/5�\����Ɩ�ʈj|��|�M�bݖݟ��Uc%f��iS�M�N+}s�e�Q�R��l�+�w �։��o,sZ��3�kM�I���M��TqnC����Ӫ�<69Q)n|�p��ks����/�a���:S�L���D����e����i��*��7��u���b�K<�Z�|t�-Uw�X*�%�Q�S,�B��]R��b�&e���ӊ���M"-IB_w3ˆu3R�Ϯ�*4��Ê�{��"Θy.�a1X�쳯����9�Kv�z�ȞM�,���G�P����S�V��d۵Wč�v��j<��o�b݅�R���JNX��fh�G6H0�h�E(�UE��?�Q�(A����	fXbW3D)�s�E����wB�9y�W Õ�!����e"� ��*�2P�V��:���y�jtW3٦H�E���PZU��9i"(WCL�i
`��IhZ3�����儑RQ��Q�)GCje�fQ]:���1,�#�jH�;���JfL��%ML��t�,.{��(bt���̋�s�C5#L�QK"/'g���'�mJ��]�'������&eZ�-��N�������-�*�,��H�"���9HY��8:礙+*˚�G���留m��Rډ��ʐ���O'<I!M��

snG��bHQF#%Hs�RY�Ċ9�t�Uk�wA�a�Z�U$e��E2E4�b&A5*Y"�X��J�"�E<��C	N����A%�7w�,�u�M���9O��nPp��}�rù)�y�7ٓ��&NU�#89v�Xd����{�l�]S�L��l|�ZK��?�Ϫ�Ԫ��*�Pz}��|OCr�}޺�⟭\wb����<mߦ�{~̬�쓃גIU>��$�Lo[�._�k��,�>�L�N#բoޛ�6«�W\�x����kڶ���Ed2v��X��HuT����V*���Æy�w�ll�y�~xi� O��|�GǮ=�q��5�1�YcI(��ŵ4�`�J�**<'yT�gS�Jjb��Cޭ���l��}�U��ޯTy@�>4ȁʌÁ0[�'aC�V��f�:j�ѮC�)��h���+��W�!����=�ԇq���^�bn�r��+an�y���]8�π{S���z��CF�!Q���.=3�}�}ՠ�C��@��_������Q���5N�k̖?U~h����UJy����e��>B���~�~���<s��Nx���,����҉��֒*6������*�R�h\W�i����З��\?+�1�b����[���%�#����zzz�@� c�S��,�`^�0?m͜��~��_�k�r��Ձ�Y����ݤr����D�O3sA�<��W�/�z�Ԗ;֩t���
���P��@������wηq���W%vϬ�v"�u�,�ǔ��I�3)�kl�ƅ��v�V��v���vvi�:Jp��������U|Լ�+�6��8�>ၾ���ޠ�n��O\y�Pw�hU��<�*��j]?�t�[k��y�������#�s�O�Â�ח��U�9�k��mX�t��U�Y�#/e��0?5n��V��O�Fuk	z/Օ���������u��{I��ü�~���ݹ�ٹ7�S�j�a�K �&�c�[g�/�3�h�tu�Ui�%��l�����.ix�������Qݾѳ>��(�v6�zk���9�(&Nٖ2	�"��tY�C�F�C]��J��	Y���ɇ�꼵���A�F����;�޽f5\���R�����bI�=NC*4��5�w���Nrx����R�q�^�Bc���?��C��0�&Yqg�=Fa�ѕLI)�K�G�^����;�~�U�w����!���ў�>�܍��~�=�!�R�f��$��3�r�8�*j��d�W8�,�d��{��˸�m��r��{�O��F�����6�޻��d��wLW<�V�>�ƶ�@���< J}'@��
�R=p�Xh����*��z�>'<V��#J��z���`ǩ���fA�_�P�Uz�*d)N�����7*�<'���̫YNZ�m+�x��(R KOnָ��|;�Vw�F]������!�7p�͏�90xRddhy7�\�z�O�x1���r���':R���r*t��P��q*_J�>zb��Ęm����F+�`,����2�7\��C2���(r�^��g�z�̙y�"C�X(��ҙ��)���{����^�fE��ʒCQ�GI^SB����3��Z��̕M<3~�¶��yMj����K���>��/ z� {���f}%X���Oa��}G~���RY],~�(~�n�3ֿ'}�R��=�B���w"�^'���;��,��
Y= �� �*˙��D��o�n�o�%z���3�q��'������r�?_����_{.A�S�S}�1Y�>ǨN�ڥ-g�']:�7����/��u���o�|s�~�=&��^���a/gb��#';�z���\��>�|rPWgC����WO����o:�ǲ%�{L'��[����Z}����Y�/�5�~��7���:���?��V�]SX΀��'7U0*/|�<&���Gr�v���R�
ո��Y���X��j�۹�:�'tw�|��t�T��l�u����V�������߁���g�����y�;�?m!z�����)Y�xh�T>�+#C�љ�]�����f�|�X�4E����ѥ99��c7],f�ʾGa�k�U�+j8g}I65�)�*����痺��Z�f�]f'�	;1�������+f:/�(%�0�fnr����ݪz˳!_�=A��vd2�C�ګ'rSD�z�������6��ܑ���,�}��0;�rA��Q�ҽ����Ly�z��K�A�̶�0#_�p��\�q_�G���K>��Tm�l�G\���>wp�z���O��=P�O�n�;!�Z�xA��ߣ8D�?m��ؼ��z��zp]L�#�a�T�s�]T�+Ub��{J�)>/���ˏx2�,d��u����9�6�xa�U��Y�Ɯ9T`L(�|ܡ�j���G�ԅz}H`���q�r�z����'ˏ��U�pv}T�>���e@����-��d�)̀��y�.��V;T�T�O���W+c>��_�l?R�n3޸:n�~���d����&:"W����O����wj=\�}4u�:��7�$h���2#��D�<px��N ];�D��B25���.�չ���Ex�D�ӣqGYڸ��7�q	����=�R�=^ w��� s,�X���t���������[;2Ǡ��7N
�WV���}�W����y��I_c��d�?z��_�G��"�+3T{i(/E��d���SG'î���8%��Rͧ��^\<��v�O_�O�4�dzc�&o�h������T��d�o9A�h�bi��`��ߙ�,פ�P�<�c���ن��OX��>��6[�^�J��x�����=�
t�۷j��|eN=�я��
\�:�t5��S�i�+xtG���s-ΰU^oi�����ג�دt������������>%T�j�����������u1���Mz�P�繣�n3��ۅ�F����;ooE�ڨzVu*�	���ht�G��,���^T�������9~�W�� *"���ȗ^�!:�z^�Մ��Js*F\)�;��י�H�y��=�Z��yi~����\�Gz�����H��i�)kvE��/zO�c=ҡ���)�rO\���w^�@�y�:=}�zIa�g�j�G]*�o�}����p7��[+����p�^z��r��z�����^��l%�>c�>���q}$���C�g��|�7�З6�h+���/d��ٛ�z>œ��(�;���Dz���Mb6��,�_I��'�|�R���9v�M�ǽ�e�����"��X���u��q��5�1��\�k�g�*��`�ŵ7�WҒ���~�����Gz�׹�ެ{>G��U�z�:o޿\z(��DTf\.�O�.�U�5%z����C��*y\U�z���Nב�����n3ޢ6�v��9������~뾨8�=�xq��.�%v`�t�^���'����+�ЎT��jK��Y.�ޤ�.�t=�%�yݯN�V�I�K\V���$#��2Z.��%�=�`%}ǂBGV�yO��-9&��A��&>�\�IVť9�-�}�{�I�̃� � �ʐ7 ����h�C�*9�Se�gx��~>��o�~��T�3��Yx
�j��J�V!^�e�K$��D��(VEK�s�2�m�m����ޟ"|B�t��`Xރ~Z�H��_�u`��"�ϧ���/B�.{Ƅ��5���K�G�x`�NЇ��[ѩQ�F;�ӣ'���{����2NB,���L>��1�-m�ȧ>�\�s�T�T����ս�.�g�~���y��F?Hs/Ł;��(TGz�A���&\	�0�7i�M��V9^��)��}���_���o+c��u��u^㑯�<g�4=[=��U���R3K'1xȝ3�ۚS����-g�q�+��h�>�p��~7�n�2%�{Iϡ:��9؏;���e��1ϟ|j�{JT=R{������P}:=u�Z@^%9.D-��}.ix������](Cǭ<�S}��F���]�޽f�ә3����:v�e��<�S�:,ӡ�#K!��{���w�Y��=�+�KtXx}���Tn��z�j��=gĥc(���ϑ�rpG����ޓq$�_zz�\����'��������KS^Bm)��7&�H�ǴŴ�퇺_W�nz�7dK��c�@A/,2��4+��)�'T ��2��Ի�y��Ykײ��#����Dl�ܗ�ݡҦ�ଈ�ۢ)�H�HN�K�ʉ���h{���_����x=�X�5�,��x��f�A�LU���^�ϫr{������Y�+��ȏc��������	������?[㎲�y�,�ĕ�+�F��#+r��5�����p\�z���d,��f��늷N��<���o�iQ�TF߽w����G�<U�&�3�Ϭ���;d��z�W��z���G�\U��i�L���4����_�9���˳'R7�#}J�������qD��7\�/����o�!�}M��՟��� p����uJ�O��Oi>��uz��E���|�Hj�Q%yM�=��x����z-�uӪ�����F7��_Qd3��b�{޿\M�3�*	�����}^��x�}�>����u�Ԡ����L;�vG��ڟ�=>��q�S��Y=��zTw��!(��Q�赞=�s)�Ȋ<��mG��r�߆C�q������}�42�;�r`?TsU�x���6u{c�K�����qN�M�l����R��g^\,��w�5�������^�+zU������F_A�8�����0��ռt4������J�u��H^��p,��+���ZҽN����jO. �#Vi�����'�d��VLܐ]��!F1�;�%B�'��9s4�����1_)-��ݠv�D�s���>_��a�a|WժԢ���y3�ҁF�O�����exm�����ޗ�q֮<Y�a�������~����r��1��~���~���l͗�>;;q3���:�NQ�f�~'r5S���P^{h����9�h��)V�
�=>�{ gΫ�N��ޅAEwn j �^������2*(.�N��>
S��y]��/aO��"�����;���������%����v|JWa��#��H�P�^\�ו�d��w�j�o֨�U�7޲.J���/�Ǟz����k&GU�~�k֕�#mbt�$�5�T;�2��>�,�uP�|;��9����T?t����U�Q=]+wm
���b�r65w�W�^�l��O���C�[�޺�Fժ�W��qϼ���:�\KL4j�m����<0ס��g���� �,ӂ XJ��r�E�����!E�d�בY�ַ���X��	��Yzۨ9���0�ˮP�9���8+�K}�Qh�#Do��\�r�Qr=����[=>tÏN��v�R�n>�z�鸯_�&�fK5�"T/��_S~X��`��k����҄F��n�䣔U��6�V�!
���]��Z��\���z�����'��,i����bs�>�����We������.P<-���a+�	Sd���|�iiLw:�#�].5�������{��T�x2�z�^��%z������Q�d�ߝ��z}H�`���6���.}~țs>�[�Fx
��J� �]���L��1�*2<.w*�4&5�&��n=�R���{�:����t�V�UX�b�I�y�\��"��>��W/�h�.�����{!���/�ɬ���ȷ�iul������)xz�b*�J0�H�Ƹ�����{^q�O��w5ǩH�W����vc���7�@�����7�a�<<J�X���*}�B�<N����v]����$��z�G�ν��C�9�:��PWs6{J�f��9�̾��6��Hn�=��gƶ��ϭ +�֯�>�^�#����~sC��-�5+���Km�����7��v����/�o�ⲫM�ϙ+>LK[�/��^��T�{�?:Ay�!��)]�R.��5���f�s�؎z��^
��7�u��.4�
��%)�ȇu	�W��ve�C��^��9��'����b�T�U|�<�(<�\=t��]u���{�q]0bgdϽ�}S8ggΧ���;9�Kۭ�H+�(v�l	`�Y��λ�����|���)�qyL����Ja]�)�ȐM�e6�q>��<ot���JҤ�\�E�E�RPa��K��T{�+m��t
|�S7	Q�`�(_,Ճ$�Vm*�1j�89�)B����r�W��{S��o�Vf�����|�*���9����=���{��W��4bO�W����yS��������ߌy|.K4�U|e� �H܍�z��S��u*7����[��;����B�t�z3�>�2��CJ�� t߽~��|.O�C")�c����[Or��r�C���\M�>�Y�Ty}�q^�+Azv��k�!��{�F�W�ؓq�����3���9ޮ�Y��x�M�{���/��>F��q����M��[>�>��U�֯+�2TW��������Zќ��yG|U�D�?�mD/�{��S^�x�|�G_ͫ���ۍ��W>�;��)��s�G�Y�����z�
��$*.zA0���.{ƅ��Zj�]O��.31;�,�ͻ�z�T�/��]ɋ��~��G��=@�Bҝ(m\�
C�/I����r����ɺ쩸�_�U��5�������1?]ȼ~��n��O_��A�~��z��ኧ6���ʯ�w�_�s�s�k��l�������-o+��q�y~�U�9�C�}�Cճ�?uX��R3~���=���_�����%�̅�g��L��a��������8��x�ʬ�)nG�J�Ai�9�AnZ�[�I����;ك��/Aݴ�?�E#?���J��Lw�֮Hܬ��9���U�35��M-���`[��ʍ��V��r�X�)���E�\ӫ�R�,S-Z����Q �X�v�8�؎�'��zk�(�u�7]5n���=�*Txl�{]�+�v5��|���y�KN����u�6��٭��Z:�i��/ ,uG0r�3S����2]&i��w٪��RR�kwk�J � T��(i�x�c)�UjK�7���!�빤���"�����2����E�Ay0�&�4�_'�-�vn��ot������؝6�;��X
����;�8M�{D�Ѫ�hOFG�>�n�w8����xcln#�p
/���3jUq�z��+T��v�BƪY�4��_c,��x6puxE���q�y���k��V��>5��,rԆa<���,�,�+>�S�� ���7���,C����U�x2�����7.���BSi�gfJbQ��VNM��m����(b�%ܺޭ�V_��Z���-+�F�v9}ö��j*�=�X9j����2�k��TKg(FE�[���w���z(�kA���W��vF���.t;��խ�J˕��ucH�.��&	gj_*z�]b���U��Be��wJ> l$��|���R���ɐֱ1ڧV��]��Qh	���Ѱk�b���Ѹ�ܰL���0R��h�PC6���7;D�[1��'kXD�AS�����XE�lI%�++{��H��㏅V��xSYWշ�:_"��lT�[DGo�986ԗV0�J�i�z�n!I�y�H��m�H=G7��;���+�:����x6���ȁ�j�b��b�Lb��Yښn��'{3�ًnV����V���q�57�
x H�nX�D7�mNK���s�ޱ�̵+�,�*&GV����h�z&͏(tdD�p�c<�\s�wN`�x�s��Ζ^��V��7���tW4����;Qg1NrіS�s�-�9����I��8#��2Ի��z����W"(Xɰ7/�4���	 ��ɺ9$�9·�_�-����1�,jG���Tk �.^�{�ާ������k�g R���6���������-���kM"ԬCL�6E�J
�v2�^Ȯ�ݘ�;J�!t[\�任���lg-wa�Qe��:�C~��;f�n���H���@|w��V�r�Z�a���Ve�F��E:�mf�LKOJu��C)�����gk�Rd���#�EKC	�U��w�*C����9�Dʬ�\;)j�y[�g��������o됳�\4̹���w��*26B��}yW��Qć��.K�*(eja���������r�t�r�AM�|o��$�gI�����R��F�n���0%2�(�
BS�%�C��K�DEQ�Y�tJ�R��J�\u���R��\'$��Nr�ԫ�#K�NE�BTV��I�(�B@��T���D�=T�;��C6�*[Y���RjR�������E�ZL�����I9j��aE�{�I(�Y^�z�Hg��^Ց�H�KH�ie��爰��#Sݎ��#���0s"�,�SH-�sQG#�M�K��e{��T���it��I��DQ&��jBj#����H�d�Ii��VR�%�N���GSB�jGM5���^ᥪ�u��:z!Լ�(˩!D��i̽ݹ���wc�ਙ
;������B��2�C�E]L�Q�yf�D������,-L+QOPt5U֞��X#��yA)VdKJ�P�,X�̋:��N��~�����(�vH�����Od53�]��P�f�U|�n�f�,�ȩ�����S]�==:�ˆnѭ�:�U˹Q����I��H����ݘ]YI�������o:��dK����ׇy�ǝ�O]+n�L{���§�=�d���Ú}�3��EeW%x�F�ʣޗ4�|M���Gz��_N)���i�GsU�}�2gE��#�m/t�/�3����ώ�'e?C�"]q�+��
���l���?W��9��ϝ���z���YS������� �$�#P����>�^3ׇ�%qs�E���� k�-��xn?S�Y�C��1�5�,��Oi�~'�M�s0c;�^���]W�*X�z*ex߮�y�ǖ!�ý�ў�>���}@{���iP�)K>�>�m{/z]fF��D�������C��-����'�����t��r<���g���n3ʈګs<I�O�g.��W!5���=Q� �5|���yM�ÿ+���z�9��ǽ;�5�Gvq��y�aOr*o���F�W��e�:��*�@�7<�����!پ����ggV�_����~�c�w��>��_�Ps��~2.�f�U$5p:����L�5[��u��%4�4��~�t�0�����ٌL�U�5�Wx�U0�s���n��O��)$���&6:ј����h�\]ڭM�J���"����ڌG��^�����y',4���]���
��ݩp�ŒL{4;3�:�JN��f���g$���u�5<���/��B��B����#��_����ώN���=Q�*=����3�*��5b{kw��bV_zEf��
�Q��y����a�����~Wr-�^'���;��w|�w��Y��4�Xܕ^�9��5�̪�C�V��-���6������W&���so��8�"������ћ��+����?��b���oG���\[�/j�]k�:��7�+����V���ʥ�Ƕ���T<ԪE�
��� �f���Q���l�wY^+���Ϸ���u��N5�2$5���||Tr"�vc���^�]���Vq�q��p����χꁳ���:4ү��������z'^JΥ�|�	>�=����C>��?d3l�'V;��F�T�Y;�fW�|�^�m�����g�w���^L�z��`�`T-��Eį/g��K�N=t�q�~�B�VT��R��2VoF7zb�0T�R�ݫ�)�K>�>�wJ���T����C�����ף�hx,�^Z�'�`�o}�O/�/�~����J5'�ѕP�#��.�o��<�ޯi��I���G���H�:����J=��=Gx�Αۮ�+z	u�j�اI���:�<�P�h㥮yG����8��.:4� O�1���^������FQ��E2j�J��
�+O7m!�(����^��c��;E����b>P��N�ʤډ󗱩ݱY�2>�t�uXni��g��S�i���9�.&�������]u���&���K���[]W�m�h�>�ޑ���C������ �,���`XR����r�Z�~+��}��^�E��[)�LT�
�z��hȏ{�m�yg�pv��]�>%��TdL|}${Ș>��'���g�t>�l�~XW����>�W������폟�q7�{�M�W���,� >��b��kf���{�u���dǧ����egP���d�ߝ���D�����6���.}~Ȓ�ku������O�/�lz�g�2!�
�tU�j����LTu���}�J�z� �Z�;w�h�Ƿu`�%�:�*�y��}�Z�`?dY�h~�[��t%���|��G+��ƭ�R}�Ɓ�d���U��}�%eN��:����86�ׅ^m>+�쎼qUO��=��x��g���1�o��7��	�����Y�<<O(��F·'�p�.�U��f��v(WO	^��]��ϛ�vF>���{����͜�J't��Pq~X)�]������n��캝Sp]o[���>)=�40�˦8.y�;�\pU5����vkn�P�9�2�/]�n������d���yTs�b�pLˣWzZ��m͚Vsܘ���t��6��:��&�C�l�^RP��{6%z��y��Z��1~�����U���`�W��נ�>�JyՄ�G����#=��T�ˌ�5��e�}$��1�G���ʭ2K�*2XB���W�{�v#�Q�R��Jq��1�Ej΍���O�{�rK��C	v{�=P��T�Qp<�=>��o�ĶW��)�=��μr�U�Uפ.��hߢ=}q��e��NI�w�Iꉔ=P&x;����r%�>�	�#-��){q.�ݮ�:��E�"����=n�ݎk��Xe���Q�"�}R�
�ZȘ/<.w���)��yY>�uX��;��yS�G���[��c���|.K5�%T`Y�+��øvnd�R�i�$;�>�wP]�y�~����V��iY�@������'Ǫ��W �5t�s_$r�������l	-�&����
��o��*�=^X�zv��k�!����Qk&1{�|_���CJ�&�B}�渀�$�끰_fB5��Ts~�ω�-�^mŏ�r=����ԛ�<�~�͕vj��l͹�X�RZ�=$L�Ru/���_���������YÍ_�[�>��$2����o����%�O�\Ubh����Ȭ����1�0�#(zR9"BI���V�)�D�3�L��"�\�4c�Mk���E�f�AӭEtʝS:�]�G���m���LFj@\�BVɯ��I��e�O���O�A���9�5�2B��~30�p`�s�4.�+MO3�TL�e];�s��C�Q��Wrb�m�̛�z}�b�z}fI�E�цl	��5��]��ey^�{ѯbT��+��ͤ:�]��ϓ�܌~��T?O���<�޺�kg��B��e�0~��We����_�N#
��鸥/����y~�y�{�k��mX�t�?uX�}T�zj+���WR\����\G5HWp:b�ڝ.��X�~��w�.��NBu��s��)�K� _�'}�c�Z_�k�{��rN_KN�g �t;���u2�J9e�[�Q��F����|�y�S�D_�'޹��:��w�ޜĴ_��:v����-������8�r���䳌���{nG�]��u)�P�\wg�z�j��4<Or2�P3ŉ�[���5��M\����d/u�G��8�M�}^(|=^�?S�Y�Cݐ]b0�L��g�=�Fcv �I��.���r�D��3���e�}wHSv�5��ё������c�\ܠ�	�T+�u8k�~�8�R�����p ��wZH��{K��6�eѴ�t����.9d��p���u9k�y6Y�b��Q����KU�b}Nݭ~�X�,rd�٬�Ȫ�S;�_�!�Dc㎕eb�{/�"�Y�7��@]�����Q�[�������/t{\��8��$�A�P&�C�2�X��'���r��}�'�{#}@{�4-J���ob���Ƕw!��_�]�,�'���jK~��@��H��U��C�+��W�#v,b�������W��T =�W{�4�������U�7�Ae@V́��p�C3ॢ�F�O��ٰ��d��+Uޜ���7ޮ��dzw���Oi6�냷^��9��|�Hj�uB���lĳn��ʶ��:���(w���u�ڿ<|������z� W�~����0�d��7<�ѓ��|�Ǣs)ё�&�uxz�������6�ĿO��`w�T�.;ޤ��S�rv��qKc�K�E���+�t�x�^m��r�߆|������C��><4˨��5
��ȿoy	�Q>�~o.A��P,==g��ڐ?j�1��y�zv����K��=����S�l�K��'��\+�<�,!뙽����0�(Á�exm�����ޗ��#�_�nb�vf�[��,�a�/z+�^Ǖ�O_�^�fp�>;:O��:��to����X��{�Qe�_+�z��i�ꓪS*��0o8������>���KGێ��A�~���;tt}D�2x���S�]!�����Ҏ61
����1���bڭ�;e�Z�����u�7[���VR�̜�i
ws�XEB��a�j��H_�d��_�'��^���K�쁟C��{!:�ݟ5{-o/L%�k�Wٝ���+�۳v�3���OVM3�,�m0)k��^^���~/=t�q�~�B�eO]�c�S�X�9�P�؇���³�=Q�����@72<�o�d[�^��zX�~�C���1�}��U�T��s>aṁ��O�U����K=��wz���O���[L���{�ܲ����C�G�S#Ֆ�ρ�]9�I�`H�wT�sS2�µV)sӾ�
��W�\y^g�����]�C��}�#}#ǯ<�dzk<}���C�*�,	
P4��6����i����\\����G��
��z�ў}�h���V{�;���0�\�iA� xثwV�Ȝ����+G��u$��p��z��z����_�o�Ը��z�����n��S��w �J��ؚ���b~���-R�qG�}��U޵�47�L8���>����m�ՠ!o5�1�Lm{�w@��n��>�����!#����}^�qE�ڿ�����p��I���Hw:����0"��I�]�����b<�k�^5�{��m�on�M�}�#|�ZW�{]{�c�*�ջ��K�MA�G�Wq֟,��9���J�Ow	�#�ܙ*��3��	P/+t�V��6��Il��B�uh���F�&<-�f��,��5A���E`���@
q�`yU0iM�g���~7N�tVԿ�k��K�Q��5�2�ge,�^�Ȍ���S&Kn@�}>ɒ�2�NKqӃ�R��{^.��x��p��x���W� }8}ח#��h�}��^�~��	�~����f���*�L5p6�?SѱuR�{7�=��cPyqձ�'��N�ﻩy�z<3��ݑ�>��n�u�^ա�eV�N�_��^�gl��-�}�&ю�����ӭs����Uྗ^��w��XH��s/�u�y�:���P�H�G��u��>U��*��EL����[�
����}��)ձ��F�=��Cz�~�ѝ���'}b�{�l_ڧ$��lL�4g��z���p<�A��c}^&�.�㨘ʩtVK�E%A姻�˅���Z���^�b�,G��I���\=4�EW����I��="�]���z<���>/NG�/�z�G�C��XVe���T`L�X<�����W��X�WO��
{���＇���I���P����=K;�<ISއw~P�v�"�Mĥdu�T`����+~zd���v�8C��0��mc<,^p �hU��N�Wc��a��
ܤ����=��@�n�J�J����N��b��I{K�j�DXf���g3K�WR%�$�9���`vf�����]�壜I:�� �in�RR��_�yM*�/����V���+�#_������Ǖ���^nmV�8��\�4}� n���=��r	^+0*����+���Z�Nב�~�8���8}�38}�>�W���F��o��v��L�5�<�� ���`>>�&�
����m��{1dP�n���}/��@z��>>��o�{נ_�O��f�̒�*����"b_�
��_����g�呞�]sۏcܩԷB*��=�u�>��'�����|`�d��r������X*\��_{H}w�2���^R���:���{���zH�~Wra��2W�>�އ1q���2MB,���L>Ο"���0���8����s���zj�i���w���U!F?Ps7��'��"�w���;TD	���b�H���zK�ٌ��N鎺u�eq�(�~.3�/�>���~��>١����ud;�P��7m���/�]̋�O� ����wj������\_��:��3�'���-ݛ�Y�mJ=о��?]D��/��U��R�eԝ���LTF'K|�����U��XW�]��_�6���,�H,�Ɛ��
gw�ITv5�z=�ʉ������j�ɜ�PRu2�����VqAQ<}z6�K>�J�ۚs�����<VPf���rV�=O��{�����e8��'����C��͋uǜ_Du���N�2E�i.'V;�6��宱�wQ�]�su��;0+�Y�.�3ވ~w	dyޣ��gF�IӤ�y�஧�tZ�3'�%]���(��>��b����`�L��j�#޽f.5eO��R�2�l������ny>�����|���y�z�\q����������VG���dX�[[RϷw:�W��3����%���I�A�|j ϩ���H��w^�<�{ף#�'�;���o�Ǹ�5�̟(�m�`��8��*���'���O��z �yFX뎷q>6���[�~Ӟr|睿Ls�.���
|:��>��6��dd��r �$0,7P ${|��G�\VQ{��,�K��)����e�l�>~��^{�FϦ���s ��+f@��n��Ȟ��;8��{���I����ke�ޯ[f2=;��t�{I~�A��+�~2.�f�T��t��T�O�����dV(��������P,5����x0���Y������ꌁ_{�뉶g�TD:�Y���={r���Pj�~�w>f����:��-�l�����}?{��y>x<�����`cm������� ck`cm�L�m������[ co�`cm�� co���m��`cm�� co� ck`cm�01��M�1����������L�m������� �6���m��1AY&SY���R ��߀rY��=�ݐ����a���<� �L�;f� ���!l 5Km-`��F� 4Z�( ���CBF�Ҿ��y�^�*�6�6�4̶�$������ml�V6�(�f�X)em��u*�)�h�dSM:cšy*�f�QZ�3m�Y��jk6͆Z��6[
0-��m���l̈SmZ���"ʭ-�2��g=�-d�� ����-LB�u��;wvr-0wp�f6ZRq�m���s�)C�{
�k�:�5l>  x -� -V ��    ��  : �8  �M�   p� �5;u�4ގVSc)�n��{�  �|�h��!t��{�]���z�Ý�fÐ���y%g8k�m{�@s�{��;�.�m����1kZ�  '��O\�E�k�{��)�y�J����z�ҩ+=瞯l֍z�����Y��z�[�֞�F���;�7�îR�֭Vm���dѵ�� �{��k�ws��UfJ��v������{ޗ�mC3U�e���/Slͱy����3�תZ���u�zW��W{�u��ۨ�s��4ƚ��Z��� ��ϊ��;{Ǻ���Ox=�l��{���P����k�[��ڽ[��'����S<{�z�ʩ<�ݻ{f�Թ�k��.�ƨ�km���l�7  �ʔK��5s]j���sZի��W#I���
���}�=���֝��үlU���{�:�]��u���p�53;�K%me�l�cT7� 'yݮ�V��r�u�[q�e�'i��Ҫ��l���ws���Mۦ��,���gk�u�]��@����Sa��kSm�wi,��  �F���Z�1�p�R��Z6�9-+P���h���݀ۗnԻu���v;vխ����p��m�� ����WvsZ��c�[I"�qçB���L���M�5�A �w6Q��        |E=�b��Ta10 �& i���0�)MP�b2  4@S�25)T��<`h�4` ���%)Qс24�414�4�O$��I  �     I )D	�$�d�d�0�Q��y4�I������G�����B��o��w ]{׬�\�X��O5�}���&���a(?�D�����K������P��C�H��2/��G����p�����xo�3��>�!��D�8�hAHHA�
� D��.@<����QE>D$#/��DmP@NE>����募i�_�B�����o߿���ִcZԒJ�I$�$�L�I#�)$��2I�I$rE$�L�I$��$rE$�|PM��M� ��@�$p 7Cq7p7Cp�E�dwSp wSp7 CqD7CpD7 Iwq7 qT7pA7p w	M��Ew pU�� �M�@�Q�WqU��7 Cq7Cq1p7��*&�n&�n
�(j
;� ���"	���.����*������� ��+�� ���(�*��.�)�(�����T� ����P���n��n(�n(�j &�n"�D����@�@�Q]�������	�*�����;�#���n*� n"�"n&��"�����&� ��m����Z�ĒZ�ĒĒԒĤr	$�%I$�J�I$�$�$����$�RI$�	$�$�I%��.I$� �I$�$�I$IrH$��$�H��K��$� �I$�$�I$�I�I$�$�I$RH�I$k[��~(ۥ���.����
`\�	���Q��V��R�b��g���Zn�[��������U}ق�����O����[Wb��$u3�ٲRbɸ�*�׸F�g�t%n�ܼԆPi���X��#^L6�\��ȑ��YoeЬ�����h�Ǝ�I{�����e�M���v�5S �ǅ�,��vo�����s�۔;2��M��u��YiZ��P2(r�n&������e�8�)�mn����A{V���Y2�M�yZq�?�᷸E�4��Ŷr��m y��[pVm�@����ߴ���t27J��Me��!+iږ	w����e.�q�sk	�:ŭh����Qw�f
w���e�y2�S*�Ͱ��ʡfn�i�e	�-��͗
4>�ׁ�n�[4�aL0��^S��^#t����F:vX���cݍ1D�]dj$�Pf�j��w.&�7z-��[��r�Cv@���*hq�gN�v`��26���+���*d����y�nH͸�v�N�5M:��7R{ B����Mӈ��N�2���b��OP-��K�Me�v6����KB��$����ޓ0��c�[7h
Z(�44J�(�+F��j)���32���!oN �q5��p��[A'@}���wy��\�k�5��;|]t��Z�YB�����1�����
v)�!�r����$�Ш�71���ܦ�4����@�
4U���H��I��|����V�Q�Tӵ���a��t[74}j���Ӭ��o�]f
��uj��yn���ZQi��̤�2�)"�T���g>OSϖRKp4�m�F�')Q2��i�;�d (���^��,�����5�A�û�{qLY���y$�U���O�J�@+œ֯s���Ҿ�y���c`�g/��;1��kU��!>��n���'[8NG�=!H����T#A;g^�yR��;�ih\0���B���C%��:��k���(i���G�^���טiv�h��=�;$u��z:��4p�JѴ(�P3D��?h:�j
���Qzv��E���kn�"��&�
�d4�e�(�qQr�:������ڼ����S���c �	����Q`���nᠾ�L�Ea<;4Y����&S5���˼$v�����v˱��v�x��ʧ��]�$�k�>w�����g*�("h�8Vd�7X4�c��f�jV7���[X�j��Y�଍��.�Hr�R�#� 5�BYڼݼ%;0��T�b�w�hO��.¸�|�f4m�<m\>��:�Z��ML��^�s�ak	��lQ)���
�V��̉�M SF�'mU�^n�Ԍ(,�P͎�Ӓ�:�hkS���4+0�6���XPB�)*�C#e�hU�J1�����`^�&�D�>�Ǥ�t][��
��<J�2j��J'umh�����crB��!�`��;�F���Ix����.�Y�9{[�L�zk"��)K�Al{cA�*�L�q3�j���miu�1Z%���j�#�-�ժ�N��ZF��lƋ.�U0;�����5�ϳ9�la%m����z���,ǔ�ev�[BN�R�l�}�V䊭�ll�#�ӿ,�*<zRe��&Lƨ�p�5> V��SA�ȳ
��Ͷ��R˫I=VΕ������ī�W�5[D������40���c�j:Ued��*ꢊ6�76�f�+�t'�Z��Xo)2�뺁����swu�6��E�Ii�L{�5�h��j��:�Wh��Ɗ�v�17�������wb��ph����hM�x��q��fg-���+lg Q��]|��j��{u�#`�{)-��iͦ�d׺���UÕw�d�Öx>QT͏�T��e"�d�2��&&�ݴ�n�kn+j�Rr��۔��Ե�)���uڂ�!0�%m��v�볖`��0�r������-�o)u��;���sCq[ݻJ���h+v�`��X�E�˺�0�;����d9M����%��!�K*�D=8�J��\[��G���n�k&��$*h,:���(�"ō���/"z:����Z�T36�:`,1��֍�N݇b�^2��P�% �[��ּ��bޠ2���qZ�Orn��&��H�����X��wz��@`щ����Q��!�
����4~v·��0n�Yl�.�U�6�φ=�{z����b����Ƴ�^&�:�N��WS� ��Ĥϝ�CL�*ď�؉�eR�>�����X˕ �y���F]cs0Sm#Wx2�ϣ{�ĭ�u˻ub�ѹ5Pn����^��y��R�_Z7Tu�ScSj�׮ic!�S2ݸC-�WZ�j-'׉'x�s{�<E�㪒]j�E^�(�6�J�Y�y��JS(VE�WQ��ƕ+4-�(+υ��\��	��d�R����������oDq�=�8����[�8�k�!�,�]�+:t�8�Fzk.�ɛbė�����;�;�3�2�#b��m�t5&�4�����QOw�ܭcu������A�č��$oi��D�>Wt�R�n&&VF��.�t�Q4$�otĒxͫ.��U��x&�()X�v��!��a���۳�W=�@�J���K@sa����!1�dyg�[��3owmX�4��4]�ǎѳ��Pے�'�r��6����0�-J���bV�xL�j�`��\w)eB�1��&�5LL���)�,ǃ5]�O�I�X�6w5:��� ׂ���-7j��{+@C�[��2]�K��j5dfM����X�a���n*���U�`e�V��pCt�5�����7[zG��@�c-L�+u�0 #L��X���V�4����=�;)�72���<*��&�R��.�]4V��)�
Y��m��d>4�U֢CG�o�*�o1*{����z����1�dq�#�B�BT��!Pٳpv�8Q��4	\�h�{�RՌ��^ĭ�7&cj��NM�����u�P�&dm"IY��>��	ŏ�kp`,^��VX�m�f^�Ϥb��-;��	70��z��)�0�@�Խ;�X״;뻾\�bj����m�y����`
cq��%��U�b�j׻@���hjðĤn���]��5Q�@�̩�V��2fx���b�?8�▎䛃 ufCt,& /%f����О���.LbFӂ91��[Y�ܭ�ԈnE���3[�/^���u���g:*�%#:Jtq �ʳ�e\̧�,`FcAތZIZ��4��ݘ�݋�Y���t�X8�OH��-�
=��`�eȘט�BS(���j�0�yT��]�E�,*,������I�j��(b �zTV�T#lIz�,Y��ZݪG*	�I�q��L!��,���P�V7/*�ŝ�h}op�q_w]+�'lД��c�t0���h�聫31 Y�h��Y�J ҵM�[���-i'��FecE�2�YUj��kfJ��?^d�)CV��̋j'��61��@�3��[6�g��)F�.�^�5�*VԂ�RhTҡMҖ����[dP�IZ�\���ڭ-�ۧN���G�
뻭W�,h�I�n��SN�����t���|�qm��I�;M+߸bI���߀(ڬ�M�X�TʫW�HTު�3k�V=y�5�{�C�I[��WnP���c�+h��� i�X�&�l1z3X���u�ÙG-�*��$Ԭ�)V��b�8r���f�2��v�硽��iNR��k�����������A��W�v��j��TѠr��e��2��ӭ7]PEjY��"��(�v���Ѻ�˨mPj4m���;/A�f��Fై�Y�%:ͺ�-�>ͬ/sF�ʻJ���h̋J�"m��⹛.��E��i�c���b�UcT	Ysu���jƆ<z�DZ71@vMŲ	z�H˻�-<�Xt6ֺ��<����o6�P[8������Da�V�q8�6w�`\�ݺ QJ���{�Xi%��7o33��\����T��{�7䕆R<A�D����'!=ib��F�q�+��E��B�ࣚ-��ɼ� ��{���M���x���'�6;�e]eށ�`x�9�n�v����E�h�X�Q�ʴ7*�)�ʧ�E�� ��D3@�{�^P-@��7-�n�K s^Br�N�fH7pBD�{�a�;��8]pUv��u�w�5Z�c��m )2��N��!�_%V�5�S?E6�c�;���� ��%6TR��$XJ��
�z��u����Rڰ��f�d�%�of+��{��O�m5]��ڙ!n��ݮ���}ݗ�m��4�]���7���ZY �l��i�Ѷ�U�7�2WZ���U�a�fb+i��k%�w'[jɳ�:�۱�5+	ï`��a�Y�i�Qn��H]j���ZA��vV�ޑʳ�,�ZE��i��e_�%@]�O)�{�NX�WS�G+&��I�|u!�f3�QL�*�I�`A���9klJW�J;�J85S-��&��������׵t���A3����YYz+�ś'��9QTt`&�X)��WY��d@ V+Z�Lݠ�ǓU�"���yP	"������N Qo���#mj9��,t@R ��S%�v2�{���{��ual����4�~("�#Yd.U��e�uaY���>o����~���{)C���T��J����>J�!OW���҂<ߞ��>>�뾜��RV����M�ݰev�Mf���n��5����ۀg�5�۳ֈ鍚�(��j��	�W!���ƨжI�X"V;�G%t A�4�e4�u�wy�r�g���f�K��E���-=B_��T�����~2������8�#g������\���!IhQ��O����>�1�z�Я�
����tlj����wU��Z���JL+mlbYׁ)�i#�V���.U�K�U��2멸(ѽ*,.����^^+�ˋ��3jtcY+jh��o8�M��!��S��lJ�CE�W.H��'(��Yf[������﹦^l��	�u�ň��';9�b�V=��f��E�8�S���9�)�2�5��F��7�\[V�MgwJ�㕻;��J.�L��f�ˎ�G�@��\*.�jF� �Iy[��,��'i�s1�1��Qii��r��.�]�ѿ6Lt��Y�d�Ԭ��)�n����k��M�mޚ',���wt6 �z���Y%��o��4�U�r����Ž�f`.ST�ϕu�j��N,}�t�*�oT�;��]�vAv5-6�k�-^#��ը�s0%���wV�E�H��8�EW]P�e��o�=��9D�C���5	��>����n2�0_P�6�wMc��f������co���D��`�rU��^��ui�r1{;u>�N�f�+쮉���GB.a�L^|u� yޡ��PQO�M��5���@7Z���y��Hs�6̡��2񪔚�d�G��vN|U�dZ��U��w,�<ɩ�Z͚l�����v"��O/o�P!Ѿ�S��(L.Z�+L�8���b�|]ݫO\7]��\�H��,6�۔�5���#����bYD�Qd�ݬ��\�(H������aZ�]Ն��p��\��	�R��%L\Pˮ�s��"�V�t�SG/c��j�-��^�H�unՇ��V���}�e�v,��鮞9Ls��I}���7/gf��8�U��TR7w��� .���ح:�̱)��"���
�SI���tΟ�S�uy�J�׍�}�7w� Iʵ���u� 0���-�m�[�S���C X���'�5��{�w,m�1��ТԼD���ս#\^(a{�d�>T|{p^c�TS�j��T����'3 ����j��d+Μu�컹�.ī��vp�������w�kDNIn�빖�(w�u������蘼�r��u��xRwi�[�-Ϯ�%+.���J�O�Af2JÐ�7�3�Q�9�����Oo�x��<��׈��X��J9�]qb��K�3Dݬz�WԌR�b�˜w���X�Ӗ���bb��4o�QdYY�-v`���$�I�0o��l���5��]nJo��\:��#T\6����R�n|g�V�R좘{���r��릃�f�X�.
��`禘��Hx�#;w�J����Y]]����{��e�Y`���M��,{˹ā�T�n�;�4M��&�fZ�/��{}�G��gtIRKM��X�canuE�T쬾�a�F]f�����$S����x��Ҩӕ�y�6��.��x���'�N�������}�m�Ǌ���jڰ{x�n�&6��`�Җpr��1���h:�'��Õ�����H�7�#"v���{NK�74��������Ӣ�:��A3RT��]� �H�s}�R�������2����uC��:3�5��:�c�8���b�z���Q�����G�� �R3C�)���m�V!�H\��݅@k\S�]�\�-�ŵ�7�����̫4&F�g%�٤�.�I5kh��xa�m�Ӈ1M�ea�浹pL�T��Ef*ƺ5��2M�����]@.Ø�t(���4:����޻0��JaֳpK��#*^>�W:�::f�IN���QE[\,��<�'Rt�:L�7kmS)x����ݍ;�.���{	$jA�u̢�%�*[|Ŏ�����@7ij���]�:$��-�m#f�`����J�	�)ݑj�R6���T�k�Ġd�ub�a3� �WRN�۾�i�X\q�*��-IRn;�'�(��t$�X���9��m�w+���Ǜ��ﭐ���lj�Uta�
L�Xt�8����r�z��Fe��QqqF�WC���n�b��-�ih;�)G\;��o\�e�+��`�s\�|+�R�v�4B�*�p��4���ʣ���)�q
X�R�q%���#�v�T|�]�E�3OY�RW��Yn�ΌgP��^�͑V���O8ݺ�T�)%O'Hӧ�d�d���veڼ��,)co9kj����:����\̧Cu�Y�X��5��U�;1e�-��D���U�4��A_JT �z��ZZ�Uͩ����[�.���� �6&gU�o���=�{W�&�yl��)��Vйd�<�7��,�0�PR�Ʒ3�ÐPZ��Z�P7�z�@rLa�����:Z�*��à(��V���8
�ئ5�Y�W��b�q�/�e���殏`�Y��b�:+(od�I �A%
�!�$T�d�Oh�:��֧.�8�O�115f���.R_'P�p˷*8�8R-�_�,:�o�G$�b9(�e`'�[��˵�b�[�
9�r��ة[о����]-r�-�9VVlG���&D�ɴ�����\��ڹ��:���ۥL��é���*Joj r7�W'�4��x�xk�����+�
1׫*Ew)�ڐ�v:j����%Z=��7�?i�I<��]�ȩ��Y�p�B�I�l60���|�k//*��Υv� �;.Ek//u�Q%�8q�[�F�X��Ye�*ҽ=I*�(����v�#E�V�rO�通Ҕ�
�Ӂ}4h���i�vʦ�/���9��Wa��<]l�q�F���im�*�����lVr�)�,P�w%�V�ĄV��s w�V�g;�et6x�u�(wpP���[e%ӭ�V�b�+K��211�K2�Жʭ��]JG��v���M5݊z�Ч��q��SK���В��9i�౴j�`�t8Z!	�Ϋ�R���:9���D^u���v��"U�9��Ƴ�M��K3�fR�ŝ�+��g-F��<n�\�	]Y6󊔷Xʙ���o֫�T0u�E]idFU�GVX�����t��[�v
��줊55+�00�cN�>�M��d̩�R%�1'Ck{(�����s�km���k�˜+9�U�����L���xN��r�pK�M�j6�@�ۜ2q��j�8"ܰ]�}��Cc����ȟ0�����>�6��MAP���-X��4�zE�F�5�ᦲ\�Z������:VI&C\�9P���dX�&q�Z�\ޡw�LY���F3� �i�=Pb�9P�Xh����WM$�ñ���4�b��Pۊh9[n%�m�mٚ����74>�!Vk(+b�k'�^�s�u�ڞL�S�Na�i���=�[�\jݧ+�� (^:���U���;*��;��7���	���YvUX#-m'X
JP�YK��HX;Y�Y�tuۼ�������
j��¯~Y��$W��{��q�g<��X�6�lX6��kE��1؍tW4�V��lm���R��e�A��GyS�:y�Ȝ÷M���vv�E��.�]�:��#����{)��sq[W][λEM�RU��[�v�S�e���������O�g�j�;�t����"b[�up�B�t٭��hC����*9ۑ�m\��N���J̬��SgI�)��^ѣI"J��m��%��*��[fHu�;|M�y��W|(Jf7�rS������ۭm���:T勔�qHf9����W]�]%rNm�-f�"�M�Jꑈ�v>�mba��{o]X|)=Χ��v&�k�+vX�^k8�)���Jm��,w=U�p��`IR��]������I��5^t$�Z��ι�ͥ�͗����qJ�-��u��Y�q2ک��۳��d����&fmQ�@oZ<of������e\W΍>��9I��<Ƭ�y+(΂D{��Բ=�-��n	�k�.c�C�/]*����}��Z�S��c�]����VU�t2�ȘG��H]`{�i^<�&�<Q�}����EE�Y2����J��4)⻏�2��'C���i�]X�[�a�oJ��)�9P��1�5�q�6b�'b�NL�;u��Mڊ*�=��n���7<�hټm�h���\���R���Sw�ˋ�9�ferѳ�����{�aa��9�Uԧ2�u�"�L���1��y;�`�=���7���+6Q���d4 ��6��rQZ�s���ͩ+b/���mjX]�)�X�,�t�S����{tCX�Y�����V���[M��f3�V��lu���r���gA�Q(�u+��vXQ� �Tx]^-K�e8�H"�������b�������qі�%�����wR��������f�=�W.���5#y�M<�ܾVq��>�U�Z�^N�y�V+�i���,ڦ����us��p�+CU�B{�)��<�d�V�P�z�t�$�EaE�,n���%œ M��Z ���$���%I�3C!U��K���Iot>�lNffwf�7��v�Nf��˶��kz�q��sA:�!Ƥ����r�W�68�$�I$�I"�1G�\-nNr�Pc�������#X��m�r��b�MS5hU����(;�2_.�'�n5�^j����?y�������Nϡ����g��6�����%�V��s�mE�~�Ӄ9_ԇ~|���ĺ�	�?���G������~�'�����8�o�qKSn�Ց�sZF	�WwX���w'̋n`Z��=8�KcioO��3���8��$��7��]�ag)�K����4]J�Ԅ��M(���W�<�*WT�v:���HNf��u�5��aQ����\�5���!��Wǳ;5՝G�+V쮩bEG��GJ�R�T�VbCUw�+&�ť֎�; 5�f�]9�@9��/��wwx���ʮAn���%���L��,�⡣���d�jp�1��u�Y�u���^����Q�@��B����3�%�=���-7�O;�Aorګm\��(��j��M�����ԛvpK �,̼��r�<6��u�d�֨��4N��)�Y�Wf�i:w�R_
�L;�f�u@+Ӳ���}�S��N(�.��\��h�E�_MYoNՁ��Vl1Q�Z]�5lɊ����N�oZ�%�$r��ؗo����w��N�R)�I$�$�!&H$�I:T�I$�$�IyE� �6	j���
��9m�d+�դ��W
�U��*���S2��_JdiYhOu��;E
W)�$�;�g�Kx�9Mp���fn��v���Yk8Ù�;ǷWH_r�թ�(%O����7a�d��74jU5e�9F��Ғ���u�
,6Y�}J���]�l02�9�٫"{�;��|ື��^MT^��Va��"4��C\Uԕ�n,��j�W:u�
�i�Y$;2uq��>�c�B�M��⦩���ր*�[�;�R5��^�Z1U�d;��Ḛ�U��w�v�+ڼ�t��ah=�z�H��`iz�hdb�添�e�.a౪�͖*��$�Պ�Ҡ�v�Kʍ�om�4�q�����q�6�@���/��c��6�b�zz���Jw7#V(՚6��:ɶ1Ls�[�L="�bm�|,V�K:��M�w�W1�QѹbW,�WGd�5�7�7z9�t6�m�r�N�M� $�I$�J�I$�T�I �X�G(E����[i�z�R�t���ׂ�vLM�%%S3p���L(�Z1]�C��i[��ѼW7(^*o��N�S�!����e�u����ᷯWXa-)�`�*��P5���5̉pՊ��)�Z$�ۺ�:m�
1nV-��
���9��.��V�MmT�F\n���+3iЙ��Mu	B�A%��W��6�pV��g5�h�|͒Wj�k/iY���Iu���W`R�]ټ�e�F��)T�]�u�)ƈx괱z���4k"jݥۊ�-�Vw�hж15��x%�Mvl��Y��|�7)Іc,fg�ȃ2BT80h������i��N������bX��^�>��,(@/�wٯ���eҬZ_U���F���<%��n�0Nu�Ц�#�g��1wf�TZU��!`S:�ШP\Fj�wT@P�b�qw{��l�ٸ����.�̹#rG*I$�l�HI�$�$��$�I:A$�Ek�����xO/���z���gf�Y��383���0�U�*u��e�T�`d�9c��)����/���8�oP���VZP�1t.4�'pU� ��W:j',"ޮF�c��^����ڝcn�!���Eˎ��ͩ�U��S7OEt�~˧�Eö�X�u7�˶�6 ����+�2}Еn���V�Y��L\)��Mǚg)�(�H�LWK��+����2��5(68ps6�&���l�{j�P��Fd�݋z��P":��l
Ucr�O�t���Nb�꥽h�Gk�m���quL���[����.��}Ʈ1�<hc�𵛅eJ
���%�u&x�0;K�@[(�k���KY�v��iWM]��o�Py��W'2�}b�ZahA
¯7���xkC,�����3���+[[P�q��ܬ��ĭ+�����f������Y��Ș2�.9Q;�!C��E*I$�9rI��$�d�t�I$�I�I�LZ`����&�rƄ6���y$�J9�1�I����ۼ���
�Z�N�I6��ʥs��a{H>���p��6⦬�˶ꙺ�eW�5���G������/1��bj�����'9��."ْ�N�UP�Kލ�1��#�	�W���p;��mMy{9Co�	$nw^�j��Zʶ(G�GwSN�����5��A�a�V�K�݆:Ʈ-�ֳ�\n�k�YKb�KA���Q�X�0�^Q�\�$�Y�vH���2�Q�n&�g	6����+'yp�0�b�{���V��x�!�pi	ؘ�NZ6���8�()Ko������H�RT�ʋVoZ����ͽ����LYY/��u�r��A�٘k�t@�-o+nJ�k��0%ջ=�f���=������{�P�N��Kw&��
��v��#�poؕ��隆�ƅiݮ�O���,���h\��m�`av+��.�nȕ1u6��wYm&�{�.UwANM{E^Q'Y$�.I$��I�2I"�L�I�I�\�
�+��ڻ8�NP޺n�/!�R7��&�@���\�[�"v[cr�d�#�\\�#{kfɳ*�;_n���e���u�t���sr��N*�,r�:�)Ι���5W"�(+� �6$!�]��Mq��9+�����z�S[c�
�� v�}#W�`���l�8�-շ���P��n���1���:W]a��[g���*�CkN�5j=� )�d��&��3v�U�]EG#��%MPe�3���iuoP<#5���!�A^hԫM��]�/$�.�!�a����2�0�J9c3q>��W���f� �r�PSI���]x�gMSM��?fV'.r�A�fe��ZHD�R�0:J���("--%@�V)m]������Y:��[e\D�Wz��b����)v�ícw�����/����[��W[T@��!�Q2/�>CeX�Š4��ǒA{wu�!YX:��l��/c�䓤�I$�*HL�$�G$�$�I&I$�I�f�{g��@�2$T�h�٤Qo_Z�9�����Kg���i�/�ܗz�SL_>s16�L���V�s�A�.t�}.CDU�,�d�g	�޻i&+:.�sH�rf��b�����u8��!���(��]��U���I�M��6k���5K��E�uXu-�V�[12+y�w�\r�`��}D�u����#�s����]�H`��Y��AZ�v�ۗyq�諢�4�v��ohֆI�е�|u�b*=�l ����Z{�t_�Cf�F�"����Y���d���: Z[�3r�7f�C*�Y�x+3O4D�Ma�\��	˸R��w҇u,j-n���g��eN)�����PO^�vT=	��R���ͩ��)�Ċ�@5�jn�^��^̎�k��FF�)�n�)�H�}�- ��Y�da"�Q�巠�4��n2��8=����z;
��O���S$�9Z �^n��
-N�M�L�I�&*I$�H$�Hd�$�H�s���倯s��rޣʓB��O(����+9�B���8�J��YԵ|�:n��|&����3�Y�vuL���;�U�i��W�����Jc#K���o��;NKV��r;�,"��ݸ�(�q|�M[���>*���uG�Ц��vM��Gn��zpRWv�Cܩ
�wPj����䆔��8Y�ـK��54�L��\�p��>�fԗ�)�uI@I{�?�Ֆ�]u��>;��fP�|�Q�#�q�ƛ{|�Dܐ<��mU�k��i�|�ծE���U�_)i�G��[�I��a�{*sf�wf6X�2�5�\ٓl��y�ݜ��q����)]�	*q��\���Z�c}՚��p��/&�q��w%[/c�7��bûG�H�w0u7�ٔf`Yj;��eŜT�肬��wŬ�EM�����x��+_,�2. ��ɻIԼ{��f�:%�ܖ�I�$�$�$���f	RI$�A$�H�I$�h�ğ]��s�w^�ݪ3k`�|L8�NS����f��W-�	w�וe�z����Fm��a�z{]�p*�p�M\�Q��`Ji!�STZ1f���Ns�571��i��k��L�F'�Km<�E�՛�66�v�L�<܏0�"�e氭%���&�*�H�u"��U��I+��5�{��o�D�}8\<�*��ͺv������о;H�3���r��&n��0�$M��YVn�;���:�Ε�!OX����w��8w+ 8���k궪�����ľ�N-v���/0#����_|S��z S�.�v�$�ej�a�U/;L.̰`R�#�{Kٕ��D�!�����GtQ5���.�κ4�=��2/�����(�-�zlo
,��O��\��q�Gk)K�%(�JTGיݮ��wM
U�<��u�W-��!����E��[�l���ΩJ�d�ۡ�j�戻2i.�G���W R�v5n#I3\/9ZW7�.,*g(���yX���F��S,�8�#����Y��T+����\#좳57���X9Z܆��ˤ�u��ܖ��;3���GnK	�G��3);]Ɏ�t6�v.'���k�eՔ�#q��tIi�"� 跕�+�M�Z�_	�1o)��4w��h���l�Z.6��3�Z�^W]��F][��n�����C�,�XM^B��Bf��ay�׌a�sbi�ڰ2��ݵԸ:P�f��)ٻ��v�l+�]�ʏ;{b��j@]<!�=/	��i�f�h�[�<�L�t��>Z.��q����kR̓��$���B�"֝��A9���Q*�+��U'�k,�t���v&�{5��-��[e���	f�f:�_ѯ;�}����a)�-����]������K����B��E��1���OlҌ�������}J"$X�#$�b:�!|�lL����q[}�v�W��n�6%#j��cn�6?��}��>�:�,��>�}��]G҅��Ҽ���u���L�&���S���������;�8�"�Ε��Z`�h=A�5�vB#Bւ�S�`�]j�22�����\6ܗd���R�U}���s۞���,Ȣ��Yz{D��oZ��Q`vּ��c
T�e�Y+F>b�`�
 flh��=��PV�7��P{\s�ǃ��t���/Q�Iv�p����vҎ�\�(���Ý��mj�[#/M@A��G�"c�)Nt��:n��&�a5]NM�ʼD3��qn�*��(���S�8A���JW��ٚ\'r.@,�.u8GV�(֓���fLA�(__X�oa���C�Mǭ�}VƠ�/�7G,v�D�q��Mq��Y��1�\���|%GZd�6�ȧ)G�M+T�.��V���L]τ<7"r����%j�oM)v\�}�!�C�Y�<��5d^mfęڕ���!qR���M̏;���	��r�c�K�A_'�>�Rd X������X"*�jB60����2�Z�K�5~�=��K	[*U���2 �+Z�֑�H���B#{P�2"�������`�$$W�!$R ��C>X� %��绾�a�ld	 Ąa 8��l2�R�Y~|��ȇ�%Aa�H#*,!	�Ilq!FS)h��)K����	J�ϐ�ж���$�,�±�
K()R��(���Ϟ�A.b%�����i@mm�+Z�.N�7\0Te������NK-F6X�����T	)JE���`b��
�"����r�2$R"�tX��!���b,ImL�(B#�Y2�YD!֩�fI@u+HA%C�G��,���bx�4�6�w�`���@�}����j�u��%Ջ`�v��jXxҘ#��[��C�������N�W�5_�}��Q���*��B_�/��ܕ�,���Ϟx�%��w<��HoB��'8����Orxech� �q��yf�l�9XztN)��뼶^90��&_C���on	��&ۮ�q��ɼW���%sG-Q�//<��W�ݞ��8Q��l^vÅ�����J�w�U�ϵt�ݎ
��(F-F�:�=���/���6���{�����*�*�Yљ&��>��]����S׸��]L��r�gk��:ʋ��D�`b6�e���a*ǥ�*�[}N��k���j~��f�ոo�E5)û1��Y3��+���:�0-����&^ڭ��=�J��ڵ^H��im��No7��pm�˒v��zj�Շ�rl�l����鉣ч"���)	9�k���U:Rgl�boM.��y��
hM�5��T����'��V�9�ȭkd��KSQs��I���籆��_�L�JxJY�=o����B��&H�x�U.y�3>�t�R.���Il�r�g�KvڛEL�V	3�ٞOY�8����~��ۦ���l�Q+�2��q��Ȗ���ehF������)U�������!�m-��S�ӵ<�T7/:��oQ�"��H�C�X���T�}���r�b�	���}��-�j�qy2$��/`�J�;&˕�
a��C��>�:fj�ȭ�/|��ɝp+>>m���|_�#���/�M�4,����$=(�=�[{\r�3�Ȏ�$�T_B�ƍ�u��ܶ�`�rU��[�y����پ�nf��߻��c��
���F��:�A8W����ru��q���؍�&�Ӊ�mYYd8�[�԰;�Kʣو��e"��|&�6��v����,چ�&�խ�_D��i~������y���jK}�Nl�;p��neXq�V����RS�,Ғ�Qs�i����k�΅�Z��I�_' )p�+ݎ=Qf�\G��]VS7
s3�N2�&M�چ��^����=�1��,��ӎf���g_�n�<z��ѳ���;�j�
i)�@u�A��7���Cr����_tQ�kū7�'��<��[���+4��TM@����*:�+�o�d�&��ʺ��z��"Σ�viGTQU���Ij��Q�܊���A��^��i�M��x��Sp
ƽ�z�`��r>�ʩ��e�u9��a�*�+�3�a�C/�Z쎗�xց�;��~�Zj���R�UM5RB��z��6a�O	N:�� R�B���LZ4b�GAhk�G5�%���]G�!S���F&T�nn��Ⱦ�g��՚�3uR1�Iػ������_UV�e����k�er�!�Ky�R��=�d�~��S���S9�9�?!�!��U���\�[J��_f��Ty�evdʃ�n6&��ūÓ�(.o�����q��u���H܃���2�Na��V�I<�N�n<'o�+c���r�𫕃7B�I2p�����������6N
6�a�B��(Q�2g�,��tz�+��i�`�;\ν�FQ�$��S�&����b��8�V�)W�������˴�Nn�x�b\pu.o9l�<$��o0�[tM�l������mu������8��1H�n��J��T-��C�.��|]��}�.nk������M������zN{u��?/�#g����J?\�v��ذ�M����	�Ʌ�'���<ks��)(3��<�����Vr�.�U�}`:8n��.+ML�%k�."E��R2��O]An�Z# ��t�F��`v�@4S����x���0�e=���Mu���A�T�C�w�7/��n�v�Xx�T���4S���CۈLp�.�1����G1�&��9�Z�Hs̔��C��7d���/Q]��ɒ���^!��oa�ysq��S�{��8�pGi�]ߟXY��>�����O����V�>��Eڨw���an��̕z=��!�YqN%[ܡ���5U����7j��u;�FL���p�c3l��[ڕP�.ڪ�If[��NVX���eF޶+ ���{��\�U��f#�2��ލ��C*��ԛk)�2�K[NU�q�v���os��;��1E���ay�Բ�nUk�c�e_F���
8�pӏ�P�����Qnc��npc�j�������k�;9��1�a�A��{*������>}H���$^�
,�� �w��t�r��]���T4����S�&f���@�\+�܊5�*8���R���.Sn��}N�9���ޱ��	��&!���o���}�zh<�=V�ETM��������M�o,ޭ��@7��A�"��G^ �Ӟ�c�wy��}3G=��42��1��y*]�p�ˉ�x�4
zh��D���.��;z���.�]�G��n{��V�\�����4���tJ�U��lp��I7:��Jt��z:��+���5T�U�Nj[�y�;�^��o�/�(;F��J]=Q��ʑy۔�b�/3&����5~�}0Gq��U�u$���@��O�c���Lf�\��rz��A�d��F7|d	�_�f���^45���|���������;��:�1H�v�����L�ݔ����o`�%=iл%�~D7�X�;��j�&�b�O9]�qC�_C/7\Yr�n�r�M�Sq��GS��]-&�s�����D�9��k!zzy��9�3� �An.�kNm|V8Ϊ�j���&��>�z����%C�ll��r6�T��d��=	{����WFC�����*�&gw���:3$g�d��gf�ȼ<���9w�#<�Y��i�W݉Q��l5�J��У�$�+�\e��d�o������Z��R\_��Dt>��|����cu2:	�C���w\]���u�®�SaҎ�2#��Ew59�,Ʒ�noc"O��8J����h��m�&E5z�W-�p�¬��|���!ڐ��C:�p�ӝ�0��%��i���M]���FgPUkx�)\k��ЮLT�c�_K9W9�+yHCrn���1����x���eu��׹�7-PK�;�}̿M�c���MmYز�2UsoaՃ3bm�V��4���y��C�� ���Y����[*2�԰k{"�M��Msyp��^l�ɜ��}�Ƹ;9L�TУ�WK�o7�t�4�]/f������
�oX�R������.�n2ހ�O{����s���э��'AuQ/��]\ZO�:Xu���f:eG)�ЎnĨPYx�r��ۉ�[�u2��_uH��;��`��:^�M��P��׫Ul�v���`O):��>�f�ѫN�>C�ڝ��;,�8WSy�zR�c�|��k"�v��z�Beˡ�lx1`����K{�`:l7�nH��v\C2���%.�[��rQ�#~��x�.�ȪZ��HiS�77Y���I���u2#cG��U�z�BM&,���:Yܜ��9T���d��Yr����ޤ�>�3Tnn򫌹J�L��]�J���81�H.�[y�6=�����g�
䷋SY �莣�{y�2�Y�\fV�-S�cs����^���"�7���Df�ȳ�;P����Ou.�]�DQŬ�F�\��Q=�fفz�7�9�f��|����RN�衱�n�C4��5��Ke�����YY_oz&LLct�kwg&�'��h��'茏�f6�lxW�^g�?��$���nu�w$|���U
N�K�˒�7�v=me.�fu�n��ضS��;j�ˣ�֒��^wVq��B�s~i�s�ʭ5b�:k7�����@�$j�Zm�7}��'�h:�k��B�Sy�Zu/se-3 u�Vr͂"��+N��q:�D�o;����؄w\ۆ���ۍ�A�w_iO�K��ǵz��C��wF���'s��$�|F|��G�Ȇ�ƅ.���PeZ-t��yb
���r�ܖNsjʉ�p��K�������n"�	Un
Tu}�g%(�ay{���&@ܼ�&�8�Wq���ooM]^�Sz��n�׃�n��G�]{�[7)�%�$�3Br�e�|��]g	�h�U�'[��b�p��<ajer4�N$���9��q���TڃQ�@���Z�kS����jfn��p�}R��I�E����wydub�B�z:W+�2pBݷv_ Dv�=��J�ǖ��*1�gn���S�ͣX���Fi�/j�ڲ(]���M��ػ�ۥ�������<=��Uv�o��_��K��k4*�O[$-��Փ�;`���A/N��j\����e`�Rc ��S�}�Q�[W�m	� SWR�L����CR2�Q�[r](;�)�]�����U[ji��\w!� �<�.x*�lz��&g\�P�u��А�v'�kB��]��:Bӛ���3t��Ġ��`�4��E:����%��[�Qpd�0���DE ��f�7��������bU�(΁f؀��,�SĶ�wv=�K��e����5S-��%���zJ(Ƭ5wwj)בӮQ�;�[	�ٻY��r�Uښ�N��e+9;���2v��f� hf
� ���m�4�j�1�����R�\^m�(v�� �}P��[�>���ciл���*3t�(JkM�gӞ�\7E�7%��3�e����^��ٙq��+/���s�B(�b`�|�H�_�`��ђ�[HAB�2@�+���%�C\]���}-��,�m,����e�62�KbW%3*�G����q�=󻈓���
YR�$%��aa(C022��ʰ��2`1Z��&7���9��&Dka�+�Z$I
��L2�I$�:��FE1`1#w�}�+8d��61!+B�!c�1F��K�	AYa1r����AR$R8�$�^iR&0�2*�$�\�������X���#B/�	 ő�V����m���Nc  ˖
Ʃ(@�1H0m��R����1^,�`@� $P�D�##��m H��ؐ%"q��� LU�V���Q�
e �6[��֮#}3�>�>�t�,w���0hP���Ry+�0r�[�;�C�ň�{!�
�	99:w��p�sZ:���U�,��o�Ī5qÝ�O��)��Oj(�ݬG�O��+�<Q���C8�3����#ٵ�V]#~�/@������d�8���Q	y9�4V�mq������䐝#�ލ~ӱP�W��w��$�b*�+
�� Pg	'���0=oذ�hh�7�6sӵӘ�ܻ��[���9�s��K�O�j`��:;d�U�^q�����y����O�>��mx�
2MOnܼ�{ӵt&+��G|T�{�*#�Jxa�f�tT����N��Mv��T��E/}N$[��G�5�竔�=�a9#�Q�~���H�0877��mO/x��$+�d5��>����~&��@&�b\�e�إ8"���r���xq{A�����^ΘsNfs���}u�^�m>]D70�/���Ȕ�9#��Rg�ط��:��S���ݺ�II�A���ە�����w�r�<��������5{F~���O���H>q��"��8i,̐�z�<�j"	���}����Ҡ�ܘ�^��q^u�=���W�Q+Yyq����l�jM����7��^F�ϲ�ӮKbs���<�����=⢡�r����/i\�;lǲ��[�a	���n7��y��}��#ǽ_��o#��
����PX�����A��~�B�luP�
L��oq�>U;����U$M���;�_p(��^��+���{7�" �+,e��b8�M@,�\�=�;9�����T���L���ߧ�4�ϜYOi;g>}���&;4����/l�t�EG:�jA���pk!����y�Wy���I7�Fe��3�(�+7ׄ��kb�0���g1���p�l6��o2�mΠV�$���Z���[���i��Z5��\a���{�%�"���v�W�FL��{'Q�����3��j�l��t�9t�{���(E���C���t2�ѯ_��o)��w��R-{���W�ԋڕy���^��\q�u��;�ۤ��r�տ%�5�W%�ͯ	�F|6���^����ϖF�3Q����CԞ]˭~�W���6��7Ϗ�)q��Y����{����BŇk��޳��|�:���\��TE�5�m{m����K�mÍÜ���@{}W�>�I��{j�=���ō<��ݫ��yP��ϒθ��񝝍.�z�O��:^į����86ŕ�u�{;�e���`6�0���b��vds�q��=���6~��].:׬�% N�+h�|��n��s`�tUr�gf��Q*nG��sN.^��G�p�g"��t&��
����gz�8�h�^ewg�wU��l�Z��|�O����|RsǸ�me�=���'J��PU��fj�_='�!����f]s1��d
��!L�R���p9��s�L�ח����7�����&y{*vjA�j-D{����n�`�M�z^	&"��;��' ��HTD�!�ۦ�5���߹:�"���@���ԁ�<�-B���"�!���]@;/0^�/�":�����8�����ks��mk;�7��|�-�5 <�@�q>��9� �^v�@�ټ�j r��Ƚ�!P]E�*����^zn����cu{=�/�uCL�E	�C�(�S��9�7�yf�aMZ�����"�!������1����ܝ�KDoz�1�|f�����_DC�Ѵ��j�H�g=����s5 +ؙ9���=�{\�O#��'���]G���'`5F�CQL�y8b��KG��@�tb�E�*w����-�� }�}2V�f~��kWޠ�����5�@��z�F��I�fl�x�Xú�Ks.4�T޼�9��y{�Z�zb�����:g��t��ntF�Y��9�ޱnk8��5������ H\�y���1�DLO��ܨ�!s�/`���=��P1�M�3�]@���@�ﻼ�b���ؼ�޽��9�sZ�*�ϵ�N����� ��۲��\�eC�@sD4O"���ҥ�Aا"��Ȅ��R:�ؚ���ن;��Y���O��9F��b��nȾ������^ʖ�,��&�����I���Emz���ov��m�k���Q�oq�{t!Ȗ�٨/`�=��."������+ʵ��M�1T�@j��B�Q����Z�9���3��گ
fx3A���D=�^�ӊ�yp��P�C1�v@�[��.�������*�E3�汢��}���ֽ��j �*��C0��OB��9p惑{ �h3��K^�Ayp��t��;�yd�C��19$��=�n��5�o�����E;�B�!j)\��=pC7��_LE0U'"�/�cT'b67Y�����b=�^׶3�x��{ܯ�b/��(n�{R�7�,�����qb����jJ�b���uI�>��}�&�a�)؍g5s^7�V��{[�WL�q �F����Pv+��,)�rE�*-A{p��# f��Q��$�SWַ|�u�{z�-<f j�ҧ-(�G����SѾ�ND�[��J��P�.f�T[j��P�Ⱦ�b#예3��x���"�G���۳��]qù�bI����&�r��P�nAx(R�z���E:�f��m��c�_�",x����"��i�]$W�D��2��]7���0iy�HT�?���~���$B@�$B@�k:����޴�o�RN@m� ��K��Wz��D/@��#�� ��6��&��ز�@�hd^��*�srj����w^���[��<Z��R��P�P<���z+P����_4�j	R���	 ��M�%���}%Q�䵱�k��tNA{=�Y1@����P=�X�`����h�P�bY� B٣��-�{
��s%��Ns�y�r�� �����-K�s��C�Pv r;J�j1Ay�-��X\@�K��}���kG/�k��s�����+�"����\��E�j��,��.n��שU(j��Br#x5/�\@�S��Vd�k:߱��׿�5ۤ��.X�E�G)�=1�3�y��2�ྈb�� �*�	ȋ���!��p~ë�k�b)��F�G�0>��<��n6�5Gb�f#�ո&�z.C����P��`���6���!��=調��v�=��ܞ�|��V�72b�Q7���(z�Ȯ�f�鈏{@��s���r b�eL��Ƶ��y�ukw���x/
��>�+h���0^@�m0��E�*!�;�載�� �Ӕ�T	�r.��+y�8���ޱ~c��xR�ը�$Y <f��ND.U��B���R�= �R��;�0f��^D�=�_i�Ϥ����h��-ms:&�n���l�n9��Q���o��#у�<M��D$�t��d
�U��=���ع4�:BŭU�4�:DM*�ϸ��$'�MN�_�C�o'��ʣ�� �H��Ȍ������׽S�vf�3� j-��� ��R^cT�@��R<�H���ᗴ���ؾ��H�n�bӹ��oZ��{��e����mP�����>��#��-��
n��ݶuw�* j����n�
v6�&wJ�6Ż�^ӷ�_s=����~�k�ȷ��H!i���!�-�Ѹ	nR���b�h�=�`���Ҧ]���P�Kހ�N��;�zݦy�o��趋�y�&j���}���)�T�+�� rC��7�B�Dw�rB۽�����ә�*��{����'���\�B��{P�i9�E$�8�@���rB���H�r:� r.�cu�ߦ=�cy�}�@�Z�0�m�Y2�Z���q�m2ڂ�^@�S�b���)�d��S�MU����w���H�^�& }���7�-E}|��"�f!��	y�_��"��'����`8�v H���K�Ͻ��<���=�7-�CQ{
�w�$���,���-b��p�E�B�T���z�*R5��
��W��=�n|��x�`s�I�n�F�LAm�|n��Ʃ�L����S�=�r.R��l�ي�.fكh/aȎ&�"z1�׽~Wqmf���;�'D���Ѹ^(_�`j	���r%�J�c�;�@rݐ�^�A�h�9��1���w����Un�Xy~�l��p��&���}�x+KM�,����t��]��y^������.*�=Ч)v^F����i$*�X��B��"0b��*����+�|�� H� Ȳ"�q�s���o�/�j��KPj)���lbv)�T�bn%�Gax!sT�/!"��ñ;�s�6z�3=��%\���w��5�o�:�"�,���S�G�C>�5��`�P��Sq{
�":�ؚ����z�R5R�1�z��V�Ӽ�g�3�}��}��k�Q5
����-D5T��!�`��Ȅ�Z&b�.�l�v%��[���;�g}��M�yݣ�{���WQp{�T��Xr��5
��	��^�����(Srפ�Ƣ��gm�[�g�������- ��u��/DOn���Gsq^EўXd�Gq��YRܡ�MB�PN@�BEsq�c6����j�λ�N�ax�#�Rf/�����/f`e�
Z���.^b�v~��ط}��ݬ�GQ�G`T �;U�۫�M�7���zӢ�/!DWq5b��й�NE�iI�]D�iA5�Fg`%�K�v�`� Z�J��ޱ�j��7���T���Ȅ�^�9q}Z�;^�����"j/��������-B���{ ��u�-���s\�{�g��x@���P��eMNA�;�EͩD��T�zG�B�h=/�L�q^Ŀ��u/�����{~�����f)��}�<�ظ� v%���D}�*�P��ɤ�����tp~�J�{��SuRN��X�������t={�՗-X���X��g��{d����*oBE��\�
��p�vp�J^á��[��O�_U~����	�I�Y � ��s��F~	&������Mˠz���b^���v�"�Ol՘�F'<���G�4s�.�<9��)L�`={ut��C�Fp��{&�� VSW9 ')����.۸ʎ.]��=�1������
��Y�x<�;(#o^�b��1;���4�(�6�;"���c���vܻ�T���՚���pHhŭ,�^ܫu���n�3�뚕W�&�vYl-?*��mg�u�0�)rf�*z��yO��级�K�毦lj�YJն��\���#���.Mb����c��C�W^Eθ��z`Bښ�c�7&3��GDl�o��}S#�Nj�I:E�MuH�*zԌq��o�Ņ����7�8p�9�ө�wxU.��̅��!�+l:�ҟ�;r*��_���}W�$P�@��s�wިfsf�I=:*m[ys��5vjy��}�w�g����V�)U�֚�p͹�#�坴��~�,�<Tߧo|��e�f�)����׾�A�J��qK��(z��J�18W��4]�q�㘽�^�z�N��q{��H~L �_P؊M�YN=6}��x��꼼��WL�tM��!�d\3��ݙB��Z�,��n8H�C�wV�i������T��#-nn:�$�b����L��:ȠV&�K=���:����Cg��j�~_M(���vf>��Z���Q���j��++�ɧs�& Ƕ>�" ��c�Wj�{���]\w�hb{�+0�m+�.��gGx����"X�TTF���LqSi��em@By��D=�I�2�Kw��[2ط��j���p7C]e�8�����0�ay�����S[홲��K� uw2���v�U���*��zhV�ݪ��Xq4���S^�n��䱞AB��S��.{���3��R]f�+hTv�@�Lt92i5�\���me)�������Z�Q�!�|�յ�h��B�4���MU*-f����}��,@S1KKa�t�:n�%/��H!9N���\�hT���V�
�B]f[���u���Բf���R<�M@�9/�w�ec[�ՍN�L�,��啌m��7��q8�q�����u֘���f�G�6s����������#U��*
e�'�c��s9xͬx���Ǖ�����V(�FV� �{T�#�!C�ݮ��R��፺yW� �G92��H���,9�!͙����9�[׀��Q�eH�E�ɼ9FC�Cu���� �M�;��aIwU���;�T��i*�G�J�i1I�Ъ��Ez�'�����e]?�N�Uf��s�(�Kk�n�68�
�JSv�g{z�a��ꥳC�x�"XV�vp�&�{zE�=��"d镌�}ԝe�N��<�9z8*�3���vUŕ!`��!΅�o \Y�5�䅵{�f#bN���
\%ҝ
̬�YD��5�^��]�ŋ=�S�P[�[����t��:��`69,c6�V�Eː��;8��
$�ӝ2�ཧ�6aԲs�n���\�Л.�JB�� Q��*1@��έ�cU��9�{d�FW��i�=���"�mg'��wk{��1���r�e�r�����DX�蕒,ʱ�	.�YK���T����Y܍D���S��s����w59kc"֒��3�o�ƫ�r�d�%��n�>
�b�>���l�I��R��n�j�u_>R�� Wow��7�J��.�����}�M��VXZ�
/�q
���ڮ#wEw���؏�~��jD����H �HVKᔍUi �1e"?O���w2���.D(���B���ZK�*`$qb��+P���{��:�Uǖ�b�0����+�勂�HD�0�H�\e`]���@�$V@����"[KD"AaAB@L2�wwA$���V�!IkZȁs)]�cSh�@��V�4��{�u�U���VQ��
�R�A�6Q jƸ,!�!.���6�1m"]��NJ%%���m!��ʐ�-d��BX�9J��Z��;���' �Rd�*�D�2����e��L�KR]��N� P2R4���'-VlJ������r5.9�`ֶ\H��$�R��a��R&2�-�A�X�D��Q'��#����^�Od��'�9��bo�<'��#Ź܌U͐���]2��|ۗ�1�+�_[�5�s|���
�H"��� ȩ"���9�s���[��՜���G{q��t!��ƸW�P���h���-������Sx�'K�W�����4Sټ[q��o�U���/�8U������`��u4�Eq�t}1:�3�l��"�#R}s[z�WE巤�Om����:�p�=n�h�w���.L8�6{�t*���+�t�|_]�'L�ټ��
�˝g�]���+b�+q����5ђ7bN�j��Kq6\����W끐���\cF�r�Ӊ�l�h�Ѭ�u)��;X��S����BD�0���c�P�[��[(>r�]ZZ�xT٬Nu�j��-��]s�ˋ������(��bcw�z&3w΂a�꽏,V��ڋ�����saK�Og*=5ݪ��O�kMakb�/L�ø�]��ZX�S/k	=��S2���U}_����FEBDd@�VDS�ƵſH�o𠹉wյ=��먁WO�xC��I�t=��ZVN�cnO?�sF��r���U�kMg��:�NM�(|�ơUR�AӦ�le=�K���I556�>�$X��;�ˏS��g�Caa���IX�����=p"^NU�=pq�i�25��H;��9w��v�CȞ���u|��U2qQ�G���!7��"M�Ֆ3	����X���u�=��^lm��O��I�Jc��D�]�Z[X|��vW��/�R�=���K�����T�[��%�6�_Mіh�翍�Վ^߶��w扥�h��S`3�Ð}�0j*�89Y��E��N�>ڍ��2��f�Y�܎��^�M�+b�i!30v��+C3�s�q�P[�[��,e���ȡd�ϫ��u��W|$��"ȁ 2*�������	��(Cu�ӽ�g�P�t5��[�;jR�+Faѕ��lN��K���!ɬhZ�k�C�;r$�,�� �He�ٞC"��_��͛�Tfv�����}",)�A$L���|;m�ȡ��K�0:.�U?�(-��G37�j9���#��s7��}��<�{F�ڻh�#��9T�������&�܍Uut�yW����b��sn�{Ot�H�	���WJ������7}kR�y��}�߹߽���ƃ�G^�W��c�L��n�D�+�$!�Y#�S���[�ߕZ�S}��5��6������w�7 zYf���X�,⚣��g_�f�Ś�;R��z�C�Q2u��=�TWڭ!���Qr1G3w���πȋ"��2(2�
�����s����������_��=�o�*��G]F#@F�f��6V&ԛ�t��Ao�k�v��������wV�Ǝ���TT#���4٫&��vm񳇱�f�|�q���jVҮ���
{�Ei�^�=3��*���r�ǘ�2���o�������C�;�[��8	�K��cR;C�	�1��p ��&�[V�f�M6��ޡ�N��>TR<��Y90��tO`wֳ�r����s���W:����hn���e��=��/�oYP�1	�k��j�JA�<QQ��a�OÉ�^:��+���+����6���RpAºc���eer������۠���QU�P_��mhυ��L��;ch���<�O��
�{���r�:4��Q��V���9�[�s����?�Ed�DI	$D�����{ֱy>Ŭv������$>�b���>�.��v�f�%�\6���{����P�/��n=��1�"Ec�E�#�ᮚ6͜U�d����.�;T�ҷ�1�M����gy)3�u�ݛ�U��e//HJ]^AB��oS�����WV�:�����Y�6��Pr��է/y��Ӷ�{;�t�����BN�P��}9�ƈ*i�p�/y��qZ�P�����Q�S�Bkhu@}���Q{+�\ in�\\�3ơ�W;1����+i�襴:�4�e�w�����L��m�j�V���#�~��Sm3g�twV�hVm�����&{w?MQ���k�z���U��s�bc�\g:�y�!J���=����ӮF�WNH���4&��S��p��ϫￗ�2" �+"�"�{W�~�WG��˝���Է���x��=�%���y�Y�ӻ�ի��Q`~�*<˸��O�Լ�SU��K`��j��kvFBf�+�������Dד39��V� �"�%ާ��n�����u��}�R���l^�������\ϱ����eH�B4���!�"�2pZ<�����W��s{V��������F,F�T�q�g�n)���]R���<u��y,Vi�g)�[��A�?P�aX�����~_Z��%:F�;�OJ��G�����k���;n���f�/yI�y�p�`mP6z�{lU�����#r�gY58>R�������k<A���mX�{�����t�5W
�lL×��g<5�9Y�I�ب:��\#%Ea���Ʒ��7�� I 	 I	^�8ι�z���ü�zsj���0Q6�V_-���q�S��]�Б����8���������\���gox��%��)o�`&����9\��,
�����/��i~���v@m/w/q#ymV0��;�FnyY�J~�~[/^�}F�ȜÞ[�G5�&E8]k��!l��S�Vk�YNME��[���i���<��o�Nm���K
�|�g��W�cN*ppIbd�����' �ȍ�Ow�YݑU'$]=ċ�� ��ao �퓗�QO��O3�8������(�����#鑤X�k�����c�1V�����V�.�[]O�p������x��8��6�1ҺꇔIǹ2��/���P�6ά4[�ݘ��Â���ؘq��%��5�n�ϊȋ"���" H(H �����wc�*�9k\�*��|�Uâ��
���Arl�1��+�y<.�kJN�]�5QF�!�R�i)��k��^�I��D�x�N-j���o>Wz�)�D�$�$����}�j��FZLi�q*?��*�kVW��f��6;le�geܳ��s����Kn^�^�m9�V�V��t�F��QR��}�� �	®�W)�L�;�z�3k������80-��k,H}N����s�*�ϩ����H�#s�����V5���e�oҾ����)E�40e��9kx��ˎ�f�p�D�D��L�%�o���j��6���b�{Y�n��8����ӧ�*v�Хf�s���F�po-�g,��ۚ��ə�YzX�D�����EM��@�p�[�\�PQms��y��O�U�T�A�E���D�/���{o���2�_L[6��s\0�J�5�zr�Im�|�/�*B��Qb-�x"%�c�vS�0D�ܺ�e�X���O���hm[ۅpڹނk�(��"�<�V�W/��9�U��Qu ��U������x=�U��X�>͇p���W޺�����==�O�I��l���T�c
55{���\�h_}���͗Es.�ˬq��j�g}�j2��v;�y�.yc�ý�L���r�U���n�a���̔:��qFt��Qbi�Қ���J��ުԳ������4@�[���b�A�Ȋ�s���5���BH�S�C����f�c\mR�r�cA��9�b�6�j���]�=Tf�f\���Ť��C4<Au��'
���M��.�+�嗙/��d�-����O��@��E��Q��
����2O���%���R�,jd�	8���}������<���n�����Io]]s��4!�#��/����J\��ǽu$�hjO�Uz�����y����{�7�۷��M�zg���s������o���3�XYq �^�D�{�9}�֓�<\s�r>���-Ȋܬ6�`�k�8��Y�H����7�P4�TK@�z�-5`��۵�\��N����}��Ozv ���t�7��u�h7d�X�L|��Ʀ�͊b���<�\��Tv�&v#�&�
j������}�F��'{S��S��K���U�]�(w1ܾ����۫�=:M��� �\֫�6��[f��g\���l�ƱP�N�V��Μ+�����78c��tٔ����$¯�V;h
v�t��FU���N=U���Y��5v��+�I�E���w;��u[�g�<.'`���z?�wh���p�W�F�1�uwK�+���nv��;ql۸i21�����{n;ƝҬw#�m�YW���P�=��2�n������k6��pL��93�^�0b��"�����$���SE�[ҹ����wn���aoB�^��p=��b�jB�|M����r@r[� o4~wwa-o-:v�]�v;
|�h���j�zp[ ���w+�Eh���d���T,��c�ct�,G��)%�|
|;��z�冯!�,vr�zXSG+�7Jhˋ�%�n�.��/Mt490(F����H>aR���Jq����¹�Am���SC�ݍ������w����m<@���Ыn9�S�N'��'��Վ{��j!`�t��㛝(��*�����Y���ӧ�:��S<�&�qX%5�X!S�rG����Ǽ�es���[R��ӵs�F뢀qa� �E-*�}�z^J�6P�h�)tM�n[|��3�K�T��Yynwb(v՘Vj��
�"�
�N�3�"�O��C[����S�M�5r
�e
�+�p��
�[�ab3���i;<w�WZ�t���1[x֋���S���`.��7�cv���x����X�]z�1�LdE����3���x`w\[!M��rY��떵�J�\!�O��HO�]�I��K�9�Ӥ���) ��a�r��i�e�0=��AX� �.n'�6��\�,���q���܉�q�����`��;쁌�GD��rT����$�YGF�+�Nxm�j���!���Hd�tPhP��7�M{D��>bq��QDqn�i'��\����F$�VŖ(}�fԣ-aQ"Jܶ��_�pr��tYa-q�Rѭ*"$iV!.0 2��n�vX6Ŧ��Fs8J�G"�lZ90�,+��ʍ\U$W,P ^�w NA9���PI1"�9p�V�F�`Yw�܄<�X`B�0U2�2#z恨�U�1! ,q��w0��� 0r�1V��iF�� �q�#:�)dW[(b������t#ᆛ�P���ki `d3KP�e�D�&������a9X�+H�[b
���[hV��@LH V5��Km����G�`�.�CIl�ݚ6&b�c��Kn��#������tر%��#��w5H$V$1�}���?�b�so����8o�m̴h�w��[q(�C�)쮼�5gQ�rJn4b�����E$A$$$$D$V"f">�����~���d�=|(?��>���,^�+R�D��j2FR�c]�+{]�a���Q�c�]�y�Sh+p�]�V�C7��y��J<���Ғ���y5�ݝ�����^�.h~�_m|Y�lx���-���;F
�m��.GAmT�O(wZ��֎�̛Ė-b�pڞ�����R]q��w�9
S�s���6�+��Q�7�-u垪�av���bӖ�z��,K�bkt�>�|wn8�W���X���}#��Ƣ�˞�9��/��E����w)����枰iI�׫���/�q�f�[:�[������pʲ��i�q�cO��v؞n2N ۬���ؔ��u�Ի�ۺ��)���C�j�ꏪVM�ݙ���c<�-{Kߓ\��ɼ����|~DVE��Q���P�+�,�{ӝ��~�=��g���tS5�О��y^���O����n@MV�D����+�l�:��H�FP��i�M䝃qƍ�d�m��ef�/�a���;va�c���umμ4��qN1©�p�D�]��n��3��׵�hj��zl��Q=� ~���*�ٝ䝁V�/��=�=Q��T7��tv��C=u�,=���Z��v{�o���}�Iu�ʷ5��`<�RR�ͷѷ��{��y~������bl���9~)���\^=�1�+��!�<_ea=w�s��Lh�Eɪ�8^�%��.��*�T��6�)^lҗEY+����>"�i�I�����\��+3"������ٸ.���c�v-�i4X���m)͉?���W����Dd$$@dU�A�U8g����1�������ޚ�5Ms�͗y46/E����ӂ�C��.'�ON��k��_xX+4(����Ř~�h���]˼���S����)^c��P�|0�'b�u=Q�¬D��:��9w����ߕԛ|���&X�S�7#awkE��;���X��ow�keq]w��2�L'����.K��5���P���hڂtk��`o-'��MP�r�Ez9�
�}�s7&�M`��#-����\5��yb
]eu���O#t���2�����}�s_+y%laQ&�m^N�d��(�1RӺW�9�Ro�Ln���d���cTl[Հ
���L"���Y�LjԷ�.D��ј��'5����β����R��)�_^����ܼƪ��5�s���"� 	 � # +") !",�-o[�9������j���sF�6�V�\�����R��R���jko��p��w��k�-I�Ew�@���(�q����a}�j8Ӹ���JyV5L$4�iMuQ�*/+�Df��3��.����^�����Z7I5�9�}����{�W��N�$��wuD/#����D��U(�����S������<Rݮ�*�Ol+'���8]���V�!�S�q�s%8��TOu���NLmڃ�kU������"��G[�qmo7��. ���>�1|!h�Y^/F�3�F}��)ȱRo�l����\i��� i7W/É�ڮ�5e�+���<�j�*�|������9����ھ�m�h*W�6b�[mT�{ܕ	����2*���� �,�R��N.�{4��q�Zq��c�ݮ�́�0�)Nsnj�3Z�-7��9�s��(ȈH� ) �������kZ��/�k��T|k#@R��M������X>e�u=)�FOD���d�5��h���}e������ވ�=�{y�ޘO��tM�3�A���� "�\��뢄^���"�s�gpCb��P
yQ�*�Z9�`pʚ�R����͹��ë����߼)�p�Zn<@��������æ��w���?.����ո��~x��jN��+lBN��i{N,㬗7���h7Q�����E3����\a�P{ۗn���>$��o.Y�z���"2�\d��HI=<�_:����^9W�SiBl��,��V<8N���Hnj@
��e���V����@#<wo(�*�޺���Һ�7hI��ü���}�^�t����ߣy��[�y\����P��"��s��m�:�N&���WW�$Eov�Y�N���B�y�9C8��9ބ��m�D��F;�|���ۙ���r��y�s��
ȣ"����2 � 'q����o3!����7�/�E�:�6��J�1@��2�o���K��pD˩
L�=�$ �)i�Z�j��5��f{W�<f����`nr���'����KG�ִu��V+	�Y�>J�
�f;	ɽ��!���nTYv8}�G�DگJ���#�/-F�U�w�Pʌ�*�tpc	5ҏE0���.���*�N��{����^�4����>�%\ ��	Ƹ*�EX���tFi��Y<�dާ��j�u֮�xh#��x)��G��N����w�=4�i>�BS�
c�.�о����OH0�U�x��`;�g��o�Fγ^�4Y��<4����?���حu壧ޕ�Z��HW��`��`�~��Y��"�D�V�X�=vl��iVV������#`r�����U�c��t�_ϊ�qm��-W�
@i��*H��ɛ�u�����kSp���CH'x�r�vT�;�ܩT��q�7�[��nO�}������@�@�� �A�P�3��W$߮�I".��͉��:��5+!>Ϯ7f�_�k�3�f뵲ݗ�)]������<geP�����sU@���j�x�F���2�F5��{� ԍ\5�Ot~~6���0�����xSUW�KD�t{�q�Ǔ�ެ3�J�#ιpc�كt��{DT�M~?^���W}�ℙ��sP�0�X�%�%��D��]��`�a�{�{#��x��פ��nѱ� x�k|!�8���(�D�Jn���6�]1Y�� �_**¢`*���1�ja����x�>~5�ƣhzZ4ō�l�դ)��3xr
�ԢT�N�)T���E[�k5���9f���K�)]!Я�'���8����Vs���CD�������Υ׿�)���`Ļ^�b�_$4Jo���{�c64uo�\��d&�o�A�^I�)|�w\��iZy��c��\���	ĥX]I�U��bvh�[Z���y����@�� ���EYJ�smk��������sj��X^_�"j
h�U��X��<%M�������H`S��]~J�e�"���3V�*�����	�2�ٳ���$�;�V���-���-5���&�w����1�WےO{�(q��]uk�Z`oΦc��^NTl�	�7�z�,�T�ǚ[�
_��o�4T�hi`����<C¤�xFR�K1�ޔ� V��`����サڭ�SttBUB�h�;FT������7Q�Z��q�g��.2��^��ͨ�N���ƃ+�	�A�x�q�Vv=î���;E�p�c�UB����8v�])�n�)q�'��
��^�'����GvT4#8A�(U}�S��h���
z|O��5�O=��֓�/2Ϩ䷲����1��fr%AUP�zDo��_K�s�q꭯dgf���N�r8�f��H_)��}��Ss�B����y�1�W@��▷<�i{ݚ��t�f�i[�"Jy�=]�P���B��4.�5Eԡ�&�')څ�dA� �@�VDI	"#�{d�'�#�V[�2�iJ�aɜ�Ҩw��zM�*���X�8�*/x���P_���G��tN�^�kF�5Z�V2��J�fr��W;���#��7���AE\+<�&�>GB��N��x[8b�͝�v3�V{��_it�k������c(A�ڳO��_�ѷw}�7�7*�Z���#���\h
U�(Hiw;��5⃅���+�v����]�z�A���xyţ�r��
�������������gS`����4&EDvxU���'� 'Q�� ��lr�>�b��ִ�FOZ���zvm;�7®�`V�sq0��]�Oc�H�.�*�+��Z�����s O|�"������U����j�~"g!�@�`F�I$ɽm�)�Z�{؈�G�eQ�:š�B���lw�0������(2���0�l6�ݣ�Hro2���T4ͷ�$�n5���B� &<膍rt'����K]0��)]Z�ޓ0��k/;\Q�Ƨ%bQ�9�[V�+U}c|9�o���+"��2"�)"�$��]Ƴ�w��Wģ�z�F1�_ɛ�� 9��T�dm���Rf��N{���v������ZWs�� ��\�+��)�Ӫ¼pˡf��v�W��;���y1�j����c��m��A[��W+�l�}�=����.Tt���fe��5�����ܖ=']Fucz�,WY�Wف�E�J*���p:��w�d9Z/B
�\�;DmU;�Sx>isb`�L��8�D�@;}��U�p��/���C���i�u��H5T4ߗ3�G��\T��li0y�Z<�����S��5�u��w{���~�)z��C�_j�@T�&�0i4v��9��9�fg��X���b�?�@B����s��t�x����AM�����>\n��182�U}PØۈB�NC.�)dA�78,�W�������w>f�ԩVk���u�.}ue�۽ȁh�����5|kN�k�Es.��ڪ#$�����[k�D��X�
Q>h���R�r����ص��@E�.��^V���fA����ז�P��sXsf���C�w0dZ~��&}�eKR7q�Y�ns�Η�Mtx�w�6��%�oh�W]�3�w�5�`�cFRj�w{a>9��Џ:�oc����(�Wq�������\���T�A[zr�x��D��Ov�7�z蓝�4r�i$��NB�|p^l�q��ΑJms�^Ns�,i%}�Fv��)��	��X��N_^�!;@����������)�2���%����rr[��f��.���L QE�5�U���ȟoo}׶
�9۫k�j�L�u�ެ6��u�eN��M�W��7�ޗiV#[���#n�b�6Vق̮�|r�WkH�Ws�]s���S���O`�m=#��$�m�N9������SJ�k�6j2%�CU[���4�O�QQ�b�i��)P�/:��+qtl�l��6o_i�gl�����hU�3Uz��U����8߮�Y��u�}��Xy=n��%AI�V�7����4��=�ZW�K��B=\ķ�Z�r�T��k��Y354���t�@oVXV�D�x7��5M4����ZD'�P.�;���Z�ń�*�-`Z�˩ǝN�	�|,��(��J�e P��P��ϵ+�s���Y�ˡ�yS3J�2�k���;k}��7�$�-�8�����2��U�F���١�MNU�hр�h5q��Yi'{	�wl0�p\�]�q�Өv�՗O�u�B�M�g�6�\:�1��s2��5+��R!�Lz��:�V�K��4����yJ4��j�_2-Sɤ,�k�[Y܄��V ���]�P0.�ov��)]%0哂e�u�oj�{v�(��00��Z�R���j1�+��Y�#���?�3ޮr|ء��MbI�klX.�5�(���3��QEطTċ.�O���i8���&1qLlR�+%�KbKZ2�"c@��w�~rq8��qSm�Ym ���)1K���),��b��HV��Ф��H�,���{�����c ,ZQe��p �m�A��}�C�筠�4�c���I��ll�Q-eѓM&��H���6������JK��-Y	hV����ٻw`	le������c�Z0�Ku��Y��g:K�f�����m���x�찛���{}�x|�`!{+�H,�:��6$���w��= �^���	�rxK�P��Bk��u�_k��@B8�}�B��B��_:B3Eج�#��H�� L�>���v�Gݐ��&�Gi���~���A#˼�9,�ͩ�yJ���ղ�hu�r�s�"�YL�����$$�AA@��g �K���#�Cۗb�e���H�,6#@�9	a���V�����^˓{����؈�)���tKK�n�:5�+�j��$�4Z�_�'�;z����`i}��gЁ�8�{J�!^#(eY��`�z��$� �p�T��NnW�TxY���2��.�2��M�����rm`�����Q�Q����{P���W��ϯvj�>1�]�7����r�ŀ��f����s��%�R�&�C�^Q������~��l�Ɠ�5J*�;��J?N3R���z2�/_1�wmD�8�x�n39q&�0��;x�o_�ã�J�|["�y�*׺aכ��+���I�?^��3�­�U N���]SU�>B�
T>0���32�4ӹ��4C�I��U�&ffrr�֘?PDPr���_u�;
t�  X�7��^K⻩��f�g�DfjcZ�x�T�1ڰs���蹨�}q�9��\�괓�c�����O���k�ݹ}�7�s<�/�s<�9>���"H� ,�H,�w�g\�}lZ��5���l�᷊�VqUz��Q�����#:cs�S8QE�+6�ѕ���+��ȱ���Mh3M<��n;ǝo.����F��Vx]ym��aߍ���s�
̸�L�s���k�ƒ�j:��a>��^xk��� �fҬӨT���m���3�y�nu?�TS��K"�[����։ya�Dx�/�l/� f�L���z��V
�UKd�YGl�����Re��b�=�ڊw'Lo�v�BA.2����:Dʢ��z��"��L��x�aFx�l�0�#��R�[�� *f���5X�A��d�\��Ⱦ�?�jњP�4�i�w�i��9\�e���s��R��;��}�E,/����u��U�܊�"�'�y���/@g7��=Gt�t��wb�i���2�YOw�a8�.Td�+��$G���(��W����\}1WM�l���حY�F����z9�P�rN>it��'L�r*���uBH",��"H) ���3��'��b������xd��QZ�6\�)��s6��/F[��|S�G�����ƭWGa��	��1X!����p��H�\��`B=y��ҫΘpMB�a,U~76�&����G�o����~�8�� `V�K�W[�9���3��.�(�@8\`�[}�	[���/F�Ѕ ����^�)Rc9�7�BF��鿍Ә9��-�wش� 	؜���\�# *����ȃ{֧,�K�O	+�,���x�5�d{I
�R�Ȩb1s�K�"�\PSZ]��o�R勵n�i�%��4 ���aL�W@K��e1�W���ޓ����"���h����4*�%�����Ohr�O��a-�V4a���̢�m�Qh�ʸr ԡ�vgkO&���v
�9����V��lk��8�R���b�}n��[bQ�|���s�5;{\��3�h�B��T�H�J���i��ꊙœ�g��>|�2H) ���(H�?DC��|��}b�y.~� E���T��z�H8b<1�+�Dm+[u�e��ڣ&�8����5m�b&YU]9ؘR�+�r��R�E�WX���K����u�P�Y�|�wV3N�,���*��4���~���qd~�d��Ep{��2�؈�����l&X��B^9g��K��DwH�����:7�@sd|G
���1 ��fOy�(z��n9��+}�<��K�������hTqKً՚y%1�#���Ӳe����Aߍ`�<7�d4��5�~x�؇ia)��1���*L̊ÆmÚo����S#�Ӑ��9��{�I�YJ4t��%ʓ2���d|��8	����Y�_gI�Y�����
��@ D�
tL�ߛiV�W�b��mwO;X�׎�9K��s�ѷ���� w��u�1����?=�da)��DR|�ݛՏ=�2�d]-���ɗu�W�p�G�dJ���#Ԛ�V��v�f5������|�H$�Ȍ�H �
wX�y�{׵g1𽵪/��j�*+����P7QF^+���O�d�ʽ��_�U�Y=ç�9�ᮡkXχ�B�p� ��4�U�,�+�_�kN�4@r�h�#�-����OMH�:�|8](�QӺ����ޭ�F�]�"��EX���#�j���B��
���E�>Z��IH2 �T��X�Wq�%��!��	a��+0YM����k�,�y��
��gF�gb�n/�1���@1 8�x�&�\d�0�q�J��-;u��ݪ�����Za���	�f=���绚$6�)���csZ���-��=����}^����'�1��ӽƧ�F*ju��*��C�U���Ƽ�t`�[+S�"��|&g���V���I����<�j��PY����Iz��
��<�x��Z���	���U�qW�u*~U�9T:2�U�/#Y/ �����~���Sb��EuװҼ%�Ҡ@��NN��}���[�\A�@�(�2u����s�W�D$D�E�I#��q������hL\@tB+���_�8�Mn�Os�2~\<5���yպ�nM��U��< �}�X䫑p���&B��胂�Wisͼ��g>l握��ÅH:�Q:3�x`Ϗ{ v ��Z N�j�ܵRV��D�$���:;��k��c�� !d�"�}�	����3s���{�3����I�'%W�#��9W�
�Q���X �ζ�n\�w�J`�'׶ F��|�N��!b�xTd�	t7�:|�=7�t��b�`�g��yS���Mc
T�h\c;Hב9��@�.�-�����֩W�%���hb�D�)hauXto��P�?a��ӛgM{��;��!hm�\�$�$p�U��ph�9�j۱�
��Q����"��n���U�Q*��M]eU��JK�e���%Z}�<�����Kh�9��k�k�>=lPƴkB�Y����s��D�(���G��Y�Z3&'f�<�*q�yr��0lba?^1���fr�����d�9�>A�	�dI@$P�/��}���ϝ�
�B���4��o7Q��T���E�B5���``O{��3#MFͱ�!LO?�U���L�M��%�J4�*�4�r����c�����a�-U;��¶L��:[
�K�y��U����5�,���B��+�
�Uj�x�N��O��U5�i�w��Mf#���EQ>�W^z�7�js�I�te�ɗ �%��;�6�n���&
FD1K�'�2��5J�՚3���9��NV��6��P�T+'�S�b��=��#`۫�`<�*���oui.x�]��F^�,�
�g��Wyp�.�*�\�pfR?�՘���>'�_VL9s5UPn��*^vڕ>�W���X��s&V�薷��\R�⻛�0�P�q!ɿ�GJ���X����|���~ݱ�t�c�Ş�B��J��h�O��7h�bW�քX�"-�f���\Ӿ�-|n߶��0z�g�x�R�Շz���N��e�.�:�5�c���;��Ɋ[����H�"Ȓ$� �3�g\�N���R�ƃ�D/��o���KƠ��s�wI�8����������]n�׮�� ��>Oz�ʩ�6^��3��qmT��'���΍�#��U9R�J�	#G�]C6�j�N���[��2����0�;��;B����r��
��,��L{o���K�SV�_���h��>�hU�x.%�)�S���Rt:�M�3�v��lPeq��&@�u�����g�0��6��no+�saL��?�&2u�Ĉ��<�n�c5�J�j�7�\�W����z���B�+� ���G3�*���Ю&88t �fS��MgoJ�I��#".v4d[�OvVS,����AH��7�6JWv����n_:Sq���QS� �>�4*��X{�S��2Qݿoc;\�2��+�U����w��3d��j�oV;�ݫ+���t�u����4^؟CtH2��lY0�JMJ�v&��R�u�qɅ��ť�*�\��,�o~�ޛ�w��]����	FA�$RA���R�3�U1S��9�e�2�Q����A�xu�|0��[s��w��ǜ	�+��T�)��s2(oP��S�S��Q��펡���t�"Z}0�^��B�:8F�o����@k,n���.���7\�lL�� 늎��� � �z�I��pC��X�@�d��N�[ꦺq�.��\I[G�������-��q��nV��*�����0X1�x~K<�Q�}7O*v+�A.�͘�qp�zF�)�{���-Ɯ�pP�x1h뮵*r"nc�`��|�kn���9ڿ��i���D2���h�<<�։�mh���N��O�a�AP"D3�]S4ͪ��2�+�T�. �V�H�6{��,�����.��qLV�3�+1eex�ƗO���>�������:5��è<�0�m�]��ٲԻ�[�h��}�����r��=|uΧCp&�b���Z !�Ix!�V��9�+uWnu�q؊J_���LD�}3�L�$� ȁ]�������}���̓��U5�rѳ�Q�Q�N�p(�V���^��wf{���1a����/W�=T���^��Y�3�e���?p�v��қ���7T��Spi�bn+� ��~��`�2mZ�u9o�n��k������_�:�[	<��?�N��K�8��FY�L�U��pO��񢢭����J��:���B�����+�#����v_��c �0eQ,~Ͽ\Y��!�@P�%eW�i\���W�SoB���]ѶD�PGV��j���č@k����ȃLy�;>�U4i٫;�a���Ї ����j�c<�ή��Jn�%э�0��!���&,�W=��N]`=��I�٪u���R֋�r���v�D�V'GK�
a��SR��C���0�}�DS��ۛ*��
99a
]Fh��3K)�t�.� 工^�:z1y�\r��f��\��k��������
�AV��:
�1*# ֘��D���Ayt�;O�:�+�ck�c����!���׌uy����@Mu�H��a�1X�E�T���b
�>������wN.���\�=�hQ{uصd��c2b�>��1=(T��1�nn��ݒ̲�B5#n�PTf��]}���\�,����B��Im���}ۤ��9c�Kt�L����NM�X�Z�h*�-���8mz���3�j��Se�?Xa�뭴qu��e�h֋�x��8�`^f*ǀ\e�4�4ำ��:l���ik�v�T7�x|/Bb=���_T�_gV���*"�٫]ŵ�uy�M���)����h�֚w�P]���[�-��.�mM*��a�-mM�Xԫ,� 1�����&����vxA{[� qT��^J��xy�t#TX��V7r��Y��ZU�e��]����"�i9R�u��Z�Z��Fq�Q~�@d'�q��� ;䡋�v1��*VJ$͍�x�rov�ս�ӛ�r�[Ǽ��Eǰ@p�t��m�:�R�����>�ݱ�v�=�� �N�7z-H�ٳ��hKx)(�ҽب&1Q]m5v�N���p̖�H%��<F�.��V��1��\�X�e�ʏ�k�綕t�a�}�Ġ�w�2�K��n\�u���j᳟��}�9OV�P��q���ƌ�2�s�3:k�}��)�+35Ag�q��Pd��['N�&Z�k���G�+8����+3�h^0�N�\����������KjvF�7j�[e��_a��`{��q�Rc�r��L�_nl0��ІԲ����[�m2������*`�W�%�s�f�d��������y{n�tz���<ob�4���$���E�$+��7�!u*C�jk��I�!��똧��)r�=<��B�n>}�}�WL\���Z�s�m~o���7YKZ�驰y�Ys�Ɛ�B���bJ� �����VlR$�BU�W4n[U�]����J{���y���w��HJl)�BF�Wv²�e�	�hM��g������y���O�B)��wfʫ�����A=f����]&����5@X�pb:�.vN'�������i�2 �{��K[�/���7P)ዻ6i���V>�����i�k�}��DH��N`hXk�Y�R!	��ݹ����h��cg��{{��4�y��b6�ܖ��rHT�Ym}��6���C��{���%�@��0�F�Jf��Q��MX5� O1��8b� a<!�&k,�&�ڰ�_n�B#���L��6�H+���1���snÊ�u�o)��5�2�zͽ]��^
[�$JoY��>���I H"���'����Ԡ��`����/U�g�[�8��Fb�A�=@�+&�T�ZSHtd���V!�@��3���bpT`3�Y&�f	е=&��|�x��r '���K��xFk&��w�ίu�������*�x(tBj\� 9��X, B9usJ�{KO�@��ǨW���P6�4=��E��T�]�8ST/ݓ��K�O2�r���kB��
�Š�S9��]��r�
N���K|OrQ�����N�_m?d��1]/z�
� oe���+����Ј��jș�I�&�9��[U�Fa�,��:F7s�vg��8��l��pW�ML5�8�y�f;��:\�F�9_ۻ�{EB �q1�=*��sq����F�����y�;1������AS���ha�l��l,�Ћ�ud�\lc��Mk5�f�`����uqS:e�)��[d�����YGa�%�!S	�2rrt����|��� HH�_~�9�gV�Z�ou_ј���'��"�T�wWWl����g��r؃�U��p�܌�N�f*�L����R��l�H��)T�w
}��\��{�{�~�1��0R���$P�1a/���y�~Ӓ]y�iF:���0u�;w�@��Kڈ����*C�Yx���
 �C8봨O����� �>�Ul��k*$D�FP�x�*<)Y�V#�U��aE@�gO[�\�Բͽ/�W!�`�U��^_E�_Q �/Ô�#��_E��Z^�y���!\�#�L�~�(�:GE)��F��Y�����N����Ůw��"1�M�]nQ�@��M<$�P]L����[Nw��~���m*�|=C짩������� �xE���OOo��0h���6Ӥi�x`kʮ�oև����病���W�y#�O�.���F*����ق�6�ő�aj��9 JL�qm�9�/�r�`)�x��]��)%J�kr��t�}0��4������58��wz1D����gr��Mb�%���H���9��$	D	d$A��@�9g}�O�3��L��7Jnnb��uL�I���Ek�;�����ò�0��):���/�?a��zDc�s�hK��Q��3z*^J��O=;�ՎSs��^u%"-:z�	�������j���T&�=�?F8\V�7���d5��{W{
sc����KiQ����Q���5׽p6`e�O�t�,E��xڕ�Js�8m����}ޫϽ�*��ePR���C��u��w�x��1�*�i-} �)������4����(����.��]L982I
��b�h�}�ʹ�3�
��>�W�` P�85����K��\�V�L��o"����Eۯ[]�N��/:�-H���:�~��h�9����à~v�!���S�
L�\��k�MY@
���p���AQ�&SjP��*�(wKV.{��C�b�)!%�J�AXŷm�*EM��(]'�>!��=��F�Nλ9���n�Y���R�y~^r�g�ŷ�Msz�3�}�@dFFD�$D�ν�w�3X��5k۵]��x?��࿴�xV�)U�/r'(�מ�/$��PVY<�ڃ�*���*fpTb��7��:�MǄT��z��Jw�s,F͑UHce��/+lE��9�b���7Q�U�4ݧ�H��dO�U]K�3��3l
�\47W|.�MR�x��pE$pq�m"��߶����� ��D4��u�ѳ�U�W:7j�%Jo��y�>~��z=��b(v����wMH�Aή�k(`���]7H��)L��X3���<ڍ�_Σ&��bnT)�2MƮϕ�����%�������>�\2�g�=���r��up������>���;c)�u�x�x2x0��8oߏ�_�W��st�a^o���>���;Ǉ{�<)��@���,L��WU�~p��h���{.S����z�!g��W��M�Th�8}7�JER޾д�L�����o�����5�� 
6Z���������"�q��T��[�2�Û1gU!���ԡ|9�s���ψ��H�� �"H	!��3DC������f7D/�Z�#83D� ,�/a����-�ڲ�b+3x�OFu�.9���������f��4�Vˮp  t1�f���w�v�$T�=��),yPD�3��e
p���w��/��n4ʁ1�� sP Cw�i�]f�<�z
�����P8�LNyb�ִ�1��]	���50����p*�q��'�tW
��e�G�V{p��$$fw_T�6�ʱP ]R�3z>R*-��X���0i�Н�M�A�|��DG�S�{����.�Y2��1WT��6N:�r/[��Q���F`J�Z �"U�I�YG�_�T�����5Mb���M��ق�@��^��p��h��^�tꥣf����ZL�_M&*�;�s
q��
bt#T�2��t'��
��N������[k>p���f�F�1�k�u����l�"��Yγs�n���K�	��"�WJ����S�jعL�8�a
�n�;��ä��߇��Q"� H� 2H�3|�[��c����7��8�����nT�v"��~l
ZK����9��[Jӣ�>�f�����C�S�J�pV��A�Z�����ЮiT���g�Re��;_�ϥ�p�,�b���4�߇i��w\ ɩ�Ά�z�N�9���f��R�j����g0�� �\�չ#Q�xgS��(��u�*��+רS�rn|�v���ɖ�����WpV2�|1���[� ��!Wr.���1IG)_��r��0�]�k���s��R�����e<�����4��.z�*�"#���\4
��\.��ꐬ�݉=Ǎ�{��[g�Uʱ��J�$M$?ң����B�G{(����3���(��n�MU��� ��u��d-  j��[��~5=4�&{*��#w���U.Q'nv[K���ne�u_݉#�Mޮ��.)&7/���y@����n�z{[����M��,��$�r�p�7$w�D�0 �s�� ��$ƹ��@>A$dY@$Y �B�������Q3���L��0f�	�ϥ�:�lP� Ў�3�5�NY�^�Jq"U;�� ߂fԺ��^��_Q�i�6T)�b��Jq�=��@x.(~�^ͻ�Z����q�h|)4*�<Y*����w���@�|XC���jh�VnQ�וx?~T�ا�S�v_Ox0xT �r����SCBfWY�`�؎<K�a�P��_"�LvmT�/ǉt>������dx}h����4CY��.>�_��Y��؋Ϻ���a��5L�\h��Q�֚XZ�Lq�8#��š�_���CZ+����R�z�&Oe�# 0�"W4�\���p~�+�4��àY�}ѡ�*���@v{R��wtU�7��^ӈ�PT�K��` ��KyP]{ېK���'���Uf	��]���<+6��j�ʁ>d��`P�۲���{��⹳��DS,glR�a��ɲt+8.˛�6����
��p1�����}����$REI$E�Y 
�5�s��K�'�5�ژ0+����&���M�N}B��3_��V�([�R�=�zp��]?���_^Ҭq��:��ɂ:��
'ǯq�>�o�3�b�I^�>-Ժkx��8��T�R#���`d�o���t�Fߗ"���X2M�1r�*3���������Yo����
�nj�q�"K��O�3ӈd��������:���\>' "���]�<�o�֌?�Q��G�������aR��e}������������S�8��X��#(h�:'5lѦ�ԄxϬ��F��B5Vw6�e��d����(����7����:�~P~{%�3�|��'�Q� c���*fv8I��.;(`9�@zo���]�u��"�SZ, ǽt����^
�5���=�����V_�w�N�f���$mQ/s����(��e'[ү8e��}��#��<�=�f#=M��S7VTY���M�sk-�{��.C�h)"Av�'�:��ʁ
���ag�������$�H�w����|Vo_+v�;7>�X�H���~�X�~DgZ���D=�4��(��ؤ�c�|}��]h��x�w]����~܋@�/5�M{gA�b����`����Y��L�:R�O����R����+�ԋu7J#|�S�{/��߱b 疆%��������m���;�A�M�<7l��pV�ZΊDԅ����
�!�ӵ�\٨�$\�{2��>�:�9.Wڪ�4���z���8��6�^�,�J{��h���D
��g��Rf��J�A��+(S��X
⾚�����q�󉹇4��8�؉c�J^�1ٷf\g��䚋}�6��t�c��C�D*������kr��_��&� f*�
q5�"�7,NEˈ�*$�^֩o#��K�h��쪿��!�+�⊃i�y˷5�]ԧ�ZWhg.�
�JbJ�l\�j�7�vk��잳NE}&\�+3���$9��m��-X�&b������Jh�[=n�r+�@P  (
���������F�\�f�1i�~���3P]	Spz~���U:d{?�����Di���:&�Z2�tܶI��Q�7^~^~�eKk��GG�KÈ���p9� ��:򘫸���o�ŭ�r�\tS�t='y[���0�.�Ǆ�H��"s�1���x�oJե̱�0�]s*���8.:J�ϭ��|lT�WK����������s��,/z����MY�2ɧ㣅��~,W�ⷪ�N�n�H�.��K5Qw ΁�T��2!!5�VO�]~����Od���?N����;���	�t����\e
�>eCJ��B����z�.�j�E���ɱ�x%�+&��Fb�6�����f�چ0h��I��h"���r{}�/��x����8Vq�]��[p{?]1Pt<6�����ξ�����gB֬���k����h]Z���"b�/
6y);�s�)"�bO��n��^���ޱ.9Y8*�Ϡgd/GXu�坙r�`��[��JU�[1�GKtn^�9�¥#1�}'EW[�N���W۬��f��6-X�n�Ge.�$�ϓ�h�Y�{|�v��uI�0uv"�SՉ�@��2\��Y(-���&H���t�t��Ʀ��V��=ǂި5X@�5m&�j���[|���DV!�����=�Aֺ���<��'3A��0����t=����T�N�vC1���sEQ��gm��2���N&������E�-MB%uu-g�T{:�Ӭ��X����Z}Aޔ���Ym�C�w�֪!q�ĺ�Vֱ����[�ߡ�j�˄��o�]��Q�4�i=��f�i��\tQ]�H2�k.g����J�Fvb��k
�]�����.���,�x&KqNA�R��d����7DXu�¬zmp��h�e$�Z�o%�N�K�/��[���I��*�g�tfR������b�
�i��f��׫��sq���ʊ�<�dNsS��⩔��n �Pݵ��
	�����Qsnuj�w���zNf:-^uݻ���5�ў6��	�C�!����5��@�e�P���`}�LiϷb�b�Sq}d&0+��tWxE}�۰�ި����e��;� =�u���_r�B�e��X�6��Hӛ0��pq�Ed�i���;���	�.b�#+���P$�V���ėw�����c����_wc��pm���3Բ�7����H����x ��*��|>a��:���X���rW@Ϙ���m���jd��ǳ-���[�X�������|ͽz��u��Itf�0�u>h�'jZ�}��'�7�/8䕽�t����&S�S��FN�+T�9k�1%���z�.F��"[�R5�0'rM��u9}��'J�v�򕶟)��(R�ץ(�^���pX~"�U
@� Q|�$��}�`a�"Om*?���8�f�4H4p#�.D4I�4�l��@ ])� ���{׷��;̡b3��D����e`RHxC޾���m�L!�"H�� �#![,�7����4�!���2�ZЁþ���c �	8�<��7s�:�	Y[��4�V]�� c��@��{�*�98���!�	�!�Ĺn7Ĥ4wQ����]�\x<�爇����Q�D<���.����z1��ֺ��n�wtF1�l��t3�>U��!���o���i�}�{w}�ڹ���8�Y%��67I�ha�]�f�k�pb`�m�Č����&�4�VY5��0�I�\+�͞�����|}'w?K]m5��)�.o7��N;�n��Rp7�`��okw$��̆�6mo'�&��
O���bf%]��~��>뻗2�F�3�:@�]z�
^�)R~�\ü��4����g��_a�r��<��Q��"%`�!5��o�������{%E�,+�	���{�ISs�S�X��*����H�Q
���&�p��>�q��3kD������}��]aN}b��P�ВD��䆺.3��I���Ȕ�P�ׄ~	]�ʹ���g�*�'��u3Bz��Ĝd�3X�;�J{�'��!�sQ"�ʋ_|iK��GL����\\l����%pwwq*�o��D�>�N� �VS�@V�r]��
�(�c�{H��DR����9�-�����bpV�,Z�ѳ?p��+i��xb0S�߿,���z���X�b=�&(���ML�D9�T���}xD5�,�'!��H��&wek�n],�GiV]]��fֺYf�
FɈ*0t\�Жk(_�i3��n��3)��:"Ks�g�p��W(�ޫ�9S,���.Ԋ��f&fffb^�'��H��i��;='Jb-�RR!0�9�ꇣ@s��"����-�ޫ���+e-���2�t������:�����1�<{�5�.S��mp��갭8}t,�m� L�����ho*�g�4&%<�Z��=��$����	���A�٫uD���* S�8n�/��{�{������$���\����H�<43��>���;eXF��BL����`�WE! ߺ'Z2��oiV8���0kή��ظP���)B�\UC���Em`�F��R��4��.��~�!V�{,s^��[��bNۧ/������}���󮶱�>�b*xt�	��;�R��J ��|h�e5����O*������5��!�{;�v����b��iD~�pq/��&E������$��,��s�\KY������Ob��V��?�h֮��X�u-�b�!W���=��
��W��F�*nS=�>bK�9٥Pʺ���Z��'K7�^���;�S/q��c�oS2���@� ��S$���ol@E�AʵV��" �PY:'4�[V�B<}ջ'�L';8�b�t8U�fPhC��s�Լ535��m�)Ն���L��(I����t9��K��'d
~�d���&����փUg�¼s�-E������)���Z\���P������+�L7����2tf#�c��XSy���p�2��_L���!�q�Y{�P�,p���S����Px	�[����I��X�pU��[>�8.@�S9��xa/��'���b�i)�ˇUkN����������j/,�o؇ '}�� 4y��Dgx���n�l��H�z�##B�:>;m�3N��2jɃ&�:����zȹ��B]���9.[��ȿ�3M'�k����i��wAu��K؊C��/0⠬����Q��>�;�qs:2�f񻒖�����;��<��p��Ȳ��dG;�	�����;�ō!�e��gq�Dӓ��������S��~�H?�/�3P�4mԽ%�Rf	��A�n�S���E#�+^߷�G �_z��Z�W�q����1ߐ�������-�;+n�5��z��p�ֈ�H��_���>�h@G������+}�T���"2i���h��χ3[��I�Pw¸D�,���)���4.zWB6�ӛ�*]��x�s,�dp�U������t��OA�j��g�Ȇ�t:&�\4p��(�Ԉ�'�����4@��}Fj,^90�E�(�N&LJ��� ��;�����tw��.����>�t	�̇h|�h��[,p��A�T$L=�����R�`L��Q�2��tލ��_�)?R�E���V�
�ō�Y���x��Z��zphyh�z�Ed��z`O�"��&uh�^��ƞϭ鱸%O�8���������%�YX�k2ML��),��?z�[�}	�?zi^��:�W��^��VԀ,�iܰ��j�ɇ���ڔ/c�z&�5.����wt � >7 '�}����\(�+@�ۺ̣�I�>�G���1����Y���Ԏ�Sq�5���2cA�pU]9��lxo��>��Z���Bu�[E(;�����Jo�������T+�Oj��&Rjy�Z(WsEƯ�-�}8L�����!�f�r�iK�Tl�(�vb�f�D���Dt*����P���Q�-p����
3,h�z�J����e�=u3�hA�)]I��c�*è�>R�2�&�z����Ɛ���޽�����H8����J@NF���Pĉ��`h�.k^r.U7�k=&��<.���:�	~L:W�^��� }�]�C9�^�������j��0`���t�]q���_�
u����}q�Ǽ�rfwMC������e;���)u�^��O��Q�M;�F
:�w�r�-�f�i��	pfX�欨�6��K�0^g?:Wb�"��S{nl�G*9K-���%6�y�Q�7���=jsJ��Ó��y��������d�$f�ι�z�C�}ʸ*�R�e�==ۿ�Z�c�����)����G(�ҷ��9,��3*\�3�3�T��t"�\h��=9��k�����ޟ��P�]ѹ��� zxpb��Q��
C�,-yڛ��gJ��X�;6)NT�5q$.:O�Z�5:}G�G}y*�2�V��
��_f�h���륦@i�_�_x�r{������w���C��x}eU�?,h\=9;'�T��1^4���Q�O0Z�ހK���k�a^"�o�g��G���o����c�)�ޭ�µ�~M��@�t� T;�/� �j�}�4\Mf׳=��l��	r�sz���_
���f"2��릫S邀��?�l|l��l{�kX(sF��VD��$@��W�x?M�Hﮰ��m����Kfn��kj2E��/b`.�Nrb�Fb���a�#�X�MH'�VVD�_v	�rI�$I\��\�5����Y����g��>!"H��!$D�}3��{Ȕ�7��n��Ȋ�3�y]��"�8��2�rK�������}wCZ�u����@l�i�Ĺ�4e�S�ɿ�-�������g:ۦ��1�W:��š?i3
&e��1��N�u9�"�B��˚��V�-[�T�燢����?	A�59�|"J��FE��_,�Ɨ��o�ZGK����U��
���Zk�CE(]�y�f�4�|Fgf,�y,�AT۫�wᐏ�Q�݉P���ꙋ�SӦ>-"��Og�h��M�����I�LT ��TJ�#��ە��y��px򧆠�`��/M�M\
�PR�^�xW�Vx�80ReqYkӞ}c�zoD��x9� 3�*c�Վ�F���̌I�{��������2v��}q�Pl�bf9�Z���l,x�W+�By�.`�$[�6j��D)��%�g	p��eꡎ[t�Ė{�Sv�K��h�=�(�b#Y��j`2���h��_0��ҵ�o���9�O�IFBBI$���&�J#�?G�9��u���f�n7f��V�Y<!/���KUp_�-��Ӧ��u�w7O5{�Wy�.S�b 7��'(�<�L添�A��a���i�����9
���@Q��W/��i�n�����d������P�P��9{?.��(��)������`��?J6� p�=��I�n��³�Z�+����Rv\"�&d��­�o 5�z��a��,�Ѝ�����t������oX����a���,Ht[<*�h�ċ�\�\~����n��)�����VO��sH"�����;s�**
�@��S~S��.pE�U*nw6T�1n$J�O!�#n])�b��uBb�N��]L�*e��ݩ-v�r���Fk2,���>/�<#	T V�6{��%��ؼ���s�/s6I\V'�]CLy|.u*�->�T�t�'u���� ���(y�XH�h5��Y�n	V�Fw_F�i&�[;�{�+n�:�
,ܢy�Eɉ>�!$������x�{{9������[V��WW�F+ТH9]tR�8u()��9��.�u�+(֪ڿ2EZU2
���sxPU�P������]���R�O�YYT�d��}�[�S�T��ͼ���ē��D9ًj�S.��b��Ց3�3�O�G	psӤ4ϧ�Pѹt��eK�Vhv��*\!�v�__��?g�K)]b_���7��IJ�B��QL)z�M�2����t�d��b���n�/�ޞe/���K��� �oR�:k|m��*�u'�o��S܋��7|���ɘ�U�2<Ǧ��.��R=��99F]��eM�/]E�Y�9�&�%�Y=-�*���QҦ3�S
j��GV��K�Qi�K�*��ME�,z�-�!w*�y�N�"��*è���vg~����B�N՚�2�/��j�|^�\e��7k�wZƬ!�T�Z�5]��]v�WW�7�^�gL�����ce���m���6�lH`�Od1�AvmI���ު�x�Ӟ!=��� �Y����b���) ��0�Y��a󝾳`�{��.ad�ܨW��r��@�iWy50'�w]	��7ͭY�(������Q3�e���ހ�n˨w}�#"��$��0*�c:6y���WS1O��
��:̃Y��i���װ׃�lSnas��D��s����1
u\�GD������t�ūz/��Om�C������{�L��?#���}���5�����_�~�rN�t#ܨ �c��¹�dT��Ts����@p�g�V.���i��@��VS�Vi��{Ɠ���!�P�Q�s��<�?�������7�Q�t�
���'KN�+�)�x�Rv��v��m�]C�����Q�[�2��b���ݜ�����˫直z�*�:���!�#Y��(���VED�ݓ�Q�}{R?����s�H�\���)���3���5��ޜ.+��T+�tNY|��lqaI���*7(2j��)n�v�1C�z{nJ�!�F��y[<���~��[{�U����_1{L=��tכ�h!� �ta̲�ͅ=¤ڹS3	�t��A��͒+l��&�tM���+@Z�h��u��}�W��UoJBa�p5��E���3���څ]�}]k#b���J���Ȧ�·t�IGkvn�Q������@,�a�=��.*}*w�,w8�:��=i4+���53�ݧ�t�_cj�,�"f�]�eY���}�A�;�v�Rʻ5�{��d�z&�R�ゴ�}���3��q�y;��ݬj���8����e-�vwD��YB�#�e�e�,�1SM���S���#w�]Շ�J^�ͺ�Ӱ�۠6v��\�`�
�m���n^�l���k�JF,�g+#����J�ȺV��Ԃ��"D�춫:�:��H�G8'P.�^�祝�wAO���R�Td��9Ӈqs�ƥ���nm����)���<�l�S�R�]�0i�K5E��7 �ؙ:H��ᰜ��Wu]�5�Z��E�¶]�/-$ų�����{)���@�{�W��z�oV�,J��賯�i9,
��}H���bxV�)8�C)y�̈́e����ݵ��O4�sD��`���3��g�r.� ��2hx�^JX�75����=h79��@�[���e���VoktC�e1�6���e�\�^����ô7���"�k骉�|�m��t�5☏��*�蔋���Q�_�`l��|@��v���e�f�������Q��@����2!�8���F.�%vPe7QemM��,�F�r��-�Ɯ�$�F6�7RUƙ�T�2L�+�n�\�i�$�Z��V�z�G�Y�>齒v��)�!0~c�H��F�J����6�d<�=��D�w��s��@�5��
��C�*�����Ci[}���}R��h�25ȵ���7f�i%��$����p6�ww�1�R��Ė�������=c<8a�_;��v��r��+n'Q�0�Su��G)h�m�!H����`y�����V00�R( +AJ���Ypb"����ٷ&�w��$�ĩ�+g��6"��)rk-��
7F�,5�wtu�ܰ!�aG���&�5p�\H�@Q��]�[MҞ�wp�۔3R鴚��n��FZ�S&���M�-��a6Ԁ�m.�s[�U����n�����,,�5	.�q�T)Q`����kݺ�d�)�'#,k��ny	b�'&�\�Qy^d�
L�'��UN))���Xyg�g�+��
�7��*�SY���-A�ާ`�~ ��z���	�1�`�֋�o� U�vj9D�r_� �:y�ûv�OIf���%�d��ƺ����S*�΁7�˙C%���F���&1�c���l���[�����e
��-�{� g�Ij�_�2Z��;� Y=D�y���1�����`^\v]"��/TT6����r~��S��'��4`�^��'~�z����hL�uo�\ܹ;g��������T D�֎#����]x7�bo�Fv
S�8$+s�EY���Ǉ0sQ�xRsU	"J��LP�}ט��Cm���B��}k��{(֎�Z/��A���0O5���x���w=m]�a��,U�Α>��?q�ܗ[h�qLS�D�Y8{S���j�YwHtu�ˑ?{+�P7���廥k �Y��~��YsʼC�vd��V��V���Y�n��7���8n�^�fwd��=�����x�1;5+�[5w�Ӝ4��t �"pB�&fv8Ij��aW|���Z0��||�ݪ�χ[i�Vly�R*:��;���^���fD���>IlE.��ׅ����>���`�J�f��#U�.�����s{��Dz+�1��q��돷f�٢Ł��� ��1����Kq��{�o�{�H0���j�R؃'[�V3��O����a�6~���uXA���Jwu�r�ϸ�����H���B��1C<u'����v�	��X�*ْ���a���dSO<B�
�5�u�X.��V��s��k-p�m������SL5P��)E��^z��&<2�.�������<�H �7G�i$Ak��~��ab	�6��_y�{��uz�fW�8�V��d�F�]NQ|��Teͱ�&��d4x j��QX�e���=���##�N���e�}wYV+Ұ1�!���B��P综Yq�7�R�`qNWb�ĻU�R�B�f���U�Nͬ�Ԧ�*	nIW5�pnدV��gG�y@��V�B��T*�F�pT�U�R���_�;�f�aҙ������ʿ!��zϮ��?o�Ø�P  P�#GL�M��^��ٓqV'K��B6�қ�*]���b5]L�Iu��O���&�p)�U鍗�v�Dx�@�|@���3���v��&��=�{��I���ssX��OW"
�T�/5m\y돖e����Rb �����g�J>�E'��3^��b�T��]Zi�愛�.	�t9���E.5`ˤ1D�^^ϭ���%��r%+����Y*`AU3P����[.x1�e�i�㯟U�~�d��x-�^��K5����	_Cð����6O1j����=7�S��yb�|`�CD��u7�B���S����/i)J���ef�~�#Y��,��븁�#�C�Sߢ9���#W7&�WoR�On�;���ON�[Y���mˁ��%�T���;.'�W��X�r�;1a^K�����9�$���RWVؼ�pU���>��1y�P�ј���G���S��q��i_�A���>����*5`���]7:7k�9�M뛾a�+�\���>���e@4U�
�@���p���
oK�I�"���p�>�~�~�Χ������#]�2� �S�X�Yx���Q6.ǀ�GL�3��V�F���D�SQw��5��b��oz�I�{��^f��Q��GB��U��C�S�#��/T{�4n�Uva'����B �b�~���tX�g���8��E���1���s$���ð�X�鹡i-M��XD7ƽ��2��q|�sy�f:���)J�j%��;�_]5oG�Ȼ�^LW�;��/��Wg
�1{F�@��b T�=���iP	F��wj_篅��pJ�*�7�8mE<�f��ԣ�b�S�uu�*wgs$8�;�����;���4ӎ���+3a�u��8��(�4�:�s�np�z�j�#����w��a�/��@*�TVy�1\�8:�uuߙ����
�3�����8|��2�u�5��u%����r'��t����+yqq�&��A�^�pS���Z`��~4�.�i����B�a��S{�b>��V2Ƀ�ʄ���Eᰐ�ͫ��_;�a�|����p
��t��oƼ�e!5��x�h#PQ���ԦP5"�!L�h-��\��4g�d{ʰS���o��e����n}�2蚂�vW&�s��{9�������G]��]�^�N{�EqKC�ם��M�v����k�����l���-�LbU�*���|Vb�m8S�|�`�����b\?�s��CUi������#�,��d�|���hGQlLTz�"x�p2t#F~Z:υ08����B��l������[��[��;Ҷdzi�{	��Qɍޠ�ɾ"���P�����(�>et��ċOdE�����E���Ky�q�dGbJ(q�Z%���qt"���EL��A�*5(�fP�66Z�x^�	5U���b۞��C�`���a�H�|������N������o�4����_�^���ОǽѺ�0�����O�*V���Z��T4T��&\�����o�Q^e?S��
�z�v`u���A	�p�9m��cK��szU�[��~��]�:�A�5w��K�P�X:��K��˨.U��?z��k%��\��Ǖ<�U�-0�͎qh*.��;� ��=���:���k�2�2��>D�L��pA��%}�v����.��{q�2V���r�����[.�s%���I�eH����9J��`�}|3����N �����V�8B~���ƚ��gN�+�Ux?�`��S��~1�u����^b �?z)�!��Y�ƐI��?�2�q�ki��[g�>ui�"+��ܕ����h0�+���֢~�h�ꔆ[���Zט��2g`��p��Lm�\W����afN�jpK�r��A������'\����� �5���C8f���O:*ae�-��K��r' :�YMS������HJ�ß��t�nEY.�z�?��s�iM�<�>�z�8"@B�(J@��R�����
W��S�������aV�tg�@c��������F�?��hq�3z�Qř�3����"���PR�����R���+Z"q#"c��P��\�������*5���"��~�pP�Yub�� _E�O	�~��bo��T���]Xe[�u�����"Y�(E_[�n�T�w��4	����Ms��Pt���VG���Y� �+�Aخ�=��$-!�Ao,�; c���ؼ
r&�A4'��:V�Y'w��hA��R���9hٮ�K�G����R�jx�`���BI�G(o{-_,\��w�q��D��e�lS.8n::'�v�E֗jn�֔X��ٻ|�q.�Ö�?8��Kq�ǆ�����M�jѻm!��(r�Ul��B�o�z�1��-ޓ-��#����a�.��:�˫���}��c�sؽ���w��a����
;�Y��u��!N�d�h���*n���ښ��pw���+�U�W��ΈJ��a�zT����rs9Tvд�7�[�2��ͨ��⮗7�ʲ*+]>��f��7]��Yy.&#dP��%�#�O�8�UzeJ�֩,΍w{�lJ����*�.s�w�A٧70$e���>@*qh�M��Ӕ�^��x$����ܴ<�p��ʵ�7\�R��!¸$����ޮ��
�onn��}�&b���ȳ۪��0 z�:|D�D�/�H�]��H������L���l�X��A��	����u.��e6�p�h�m�9�"@�����ЦyӤ`���[�I,����[�����X��2��\��7zJ4������	��H?��QW�{��-0���L���{"{5�g2WB�:��$�ݭ�dN��a�֤�Dќ�ȷq�����u��� 5Ը?]@s01PZ7f�hK�rQ`vF���zυ~񫟐4'��6�G������|k���z���i<Z���r*a��*�]��]x_�
��3k�t�����Y�Ќ����Oޫ�D�x>y�C� 7N48@��y�+���V��=�6w?>x��~7��*V�TV~~W u��Ɛo
��ף�jo;w�@~���X�:���i՛��*�@/�I��×��]*gRQ�n_ж���}x*�zxZ62���<km�>�]Wf�>-rS{���CG�ƣ�h�?d����� �g�����q�R��~������1��q��.����VQ3b����)ץ�(�[�ɺ���ߔ����[�/��kV2蚂�E�l��� �.��	N�t5�z0Un)75&��E�BiN�]ja�qe�����U��XJ''gZ�1��wD��gaT$�%����'eT��&�"28���S��{wc!�����������}�X"�3:�=�5�|�Po@�ӓ�u�1#�&����-�e�*��e�q����i���Ǘ'���	�Q!J��6zۻ��@�p}��U�\0X���I7�%��t������&OF���~Z=v�
��-�.�J��ͅ��І�ޫ��\�|>zh
������J�5�}sN��
H[�{��ۼ��Tw���Y� _�Tw�*P��xy�S��J��j$'+8�H��3��.J̓�X�q�P;u���Kc�0�YBZ����sy�ܜ"yT��r����z�;�%��R��m�g/6#+V�o�:1vЊf:�ݭ2�����w��=0��^>4t)՛X�B��妟[��=�� ��B�m��.�ǉ`փ��5+����GE�Q�����[�L�����r�q�g�P��^����CX��T�J��j�ѕ��/`��NR0~�1�Buk�׎�Fk��A���\)�0�T4�+ ��8i#��H�q��B!ݝW�(Z��}�z�gt�N����/��Ŝ���Lh��ګ���Wd��R��(��l�V]��9R���Cj�����(6�eL���'rXNZ����Ob vXf�,�ݖH�{j6�8�!fÒMf�;�q�u�Q���A%0�s4�*c�`�Ui�se��'hʅ��7���s;�VP�1r�i���^��]S�s��Y��ub��SM��Ó��7��m�8;mft��*[�L9nl�pq�+A�:��c�U]����9R�u�Yսê�O.�[֩u�&�y]wѝ�J�	��+�6���d:ᴊ��eoB��T�I��c��lҳS:��ڀ�/��m�AP_ 鎹"�C 6HV]�`r��\���Nb��(w.��ë�'="6��Wr�:�yǅL=�O{\�x��a�[��#���8�n58���`uZ*2����z���6�O;�<�=�λ(e�SF��c�
H�N]Ʊ�]!ȶ��U-@mٛ���PX��yPt��"�����p�怢��'spW9r���s&��3���u`���+M8�v��=03QZ;��Y��C��� �<li�I�>5��I4��h�y�r�����Z��9�3��F��P�r�9�t�J�̘:��� ��<,���r�b�b�si��ڜ��o|Fz�uǩ��o;��o1��F��!�x�<Ub<��a]lՋ�܂��N��b�d�K��؂�0��pr���b��6r����-洚�2���abj���f'!)c��Z����y�\�E7�
���4�� -�o1)Mv'��8/yM2+��v�M�>l�_�
 P͋fiV�n�.ԉ�Pa�4�M�e�� �_	n����!	!� `@8a�����@�d���%%֐ �����lA2��;�kn@(�b�{]	�f��=�{t�4��{���0T�@ǜ�v�8�!*�ȣAP'�����I����<)�(2��c	
�0��5��3�vP�Ad!�b����{����@�İY-e$ض�rII ©	�ip&�ww�2� �� �@�"�%],�;hJ�e#���v��.J��" ���0��+U+���h����&��p�`l�lQ&�M��"L I"��cH�em�k*����թ+H(�H�Ǭz�L[��y�É!]����]�T�WX/m>\[V�͗�\�M�GQ�������x�"�����ȿƷ&�ǫNNufItЊ�7;��K�'U��JwH�a����\,[۱�{��ÿ�����v�̟-n�#�c��P��n�E;���"�U�r�f6������U�K.j�X�����t˳���qΡ>o�������;�2P��~᭔�bW�=>����W�+��-;J���ͱ���!8��ׯ�;�P��VD�3����3d�
�f�n.q�/7V���dъ��qz&~�t'c�;�bns���㜇���UA��x���!c]���u%�#�5�%�z���#W<JT�ܙy`�Ҥ�Di�	u��,��z͹M�攝�d
���P��n`�+�䬐&/D�S��!,Q��\]�J���n�� _	�(��=���ۑ�i&I��㡬�c�s����x2�n�װ_����TK�ܰ[��:3U�T�$��'Y֏鋿l���L�W�&{�I��π]F�>U���wS(���G�]SGa�|*���B����<0yw=���T�ic����Ǘ��ޫ�p�d�+�����ڷuEٯ��i��Nۍ:�X�`�7�Vw�7<�gfC�r���r�)M���N�n��T������eV/''w�a�q�5��j�M���޴uzo�*�ܥ[�+�*^��
�:YV2z�ISd�[ܸkon��8	(��جQ�����7[�M�	?|�֛z_A��'����(�捽̝u�H��m�%S&mZ����r�	s�5}��K<a�L��aș;Z+3�d6"�4�l�3���Q�J�dv�N`�|c���4�(������%kǼL��^-l�
����i��͢Ub���3��(�5ջ�ʍ�=��J��@�>���④�^0(�I��։E�`}�>y�`�(�<���n�S��q�᳹��W|�Eq�۱>��>���9K�W�o���ַ&ܞ�l�r�p�ޞ��/ v�h�B��sR�`��Xu=Ԝ�m��4w(k~�Yu��䭼^��<���}�H� Q�U�ُfǈ��jF!���u��q�q*�A�uvVCz���U�s*2t�(B��F.�ʺ-a���M��zw9�A����\�����RP����k����//�#�4Ə�^3z���i
���C_n9�'���T?[7ni�i���'8&I�9����j�w+~7��{c�h��g-�z�j�5����0���u����ɪ&�S�{������NcXrz"Q��K��e�F�O3䲾]�vE[�0�[3,F�?g��8r�~*��{E,����}:P+�{�F���7e..u8��[�;��<Z��{$by}cr��U�mEN�q:U�
=5	��$s�svʌ<�+����}N����1���gwѮU�,���ej\�} �}7m�����r�9~޻O.Q�יż�{$��v��峺���{b��@�P�=h�į��B���^��6=���TJ͎3�_�iV���o��o�)c������*��p=��T
����Jj�(��f�5M�xhW^op23�oz����V�Y�TS��H����Y+(5qvƩ�Y1��Ed�scRp�<M��ֱ��7*�<���KcM�d�M("�E~�r��_C�W�Ў�t�{����9��}�����Q��;+�W�t�zZ%�o���7Xz��&��C�uݯݨ���.��������~��Jm1u���%�5X{��o��<Ձ��/k��};
��������S{3n=��O����9.ϫ��f'̧�Ϧ�~�&w�n�"����y�7����~r8�Q���z�+�x�\;yshp�`�����q/�NeX��>�G��RS�|t��`�f�y���y��=�u�"����{}ϻY��-���YM@��{j���N�H;K@�����ѴnnJ�*8 �w�j.�X#���sAt�%r��v��ޡز$�`N�L��a���L�n7�u&ޯ7���]Ph���8c���c��N����W�I�z���|�ʮtqbvzO��Ҡ�.�Ԫsn�"_}xB*�W̪�s�bh�s����l��fۗ\�ϯl!�W����$���)٣�6��rT��.��#f�;�d"�d��w�3�����!鞨��].�;>�Mb��q��/��7����!+Y2#�.N�=Ue�x>u�;Y�Y*�����\cw��{s}F��h�u��5��E��B���|�)0��nn�ؼ�G>v)^oy��W���,*���b8�5H�U�>_[ԭ��p�t���Ptv����L���FdXh.�f����&�[�[@��B��lpvM����]�������؜;Bzm��+zB�e�{)��$�kxɹv��R�=P�Q�+(,g���In���&�//���]��҇'&�>Ǫ��q���szN�$�-0/-�N�շѾ�6�b�h}Z�y��ϢjNpٯ�j����X��G$(��5 �Ȥ5�3D�V+�M�r+z�s&��YGjZM%<��s��ڹ��&��{�8�Nvo�,Q���P~�oumgb|�	�8�%�&�&-ڶ��V8����+O#��*At�	}7�;�U��;���n(ؤ��'��{x�9�%$���ü��N��.�w]��x��ᩍ㬦�9�� ���*� ���_�\�@02���4�o��F$S�6Ok�v��J�ž�N&����Eiu%��	��ޮ��7x���2�RNjd���j[ޛsw[�@�,*�y��G�5ul�Nj28��H�8P�V��Dr�:�8�v.���������lUʻ��R=�x�l̵�L'�|��ӹ���I�����C �C�j�����@�z��-5��W0����?^~ȧ�y��>�.��GM�Y�����xD�,�z�;�O9��s����/n�8G��3X��]�+��Y5�>�ˬ������4�TBu�����oY�q��p+)x��4��w�Jr^,w�t�;ݱ�c�J��.7g��ڪƮ���e�����&o㯪T��:x����"fjq�\�h���Ÿ�s�!�s%�W��;���j/�٫��U�5b��,�}Kf�Aޜښ�-�q�r
�W~��=V��V}N��y�+66���Ť�G@[�4�Q��������39Gy7y��'0&\�:AS�i����O��b����N�}}��d?+��<�����}B�w�ZQq��ݕ�K����b��E~y��y�7�j���V�>���_�MJ������8��7��B�ဩ��OC���w��ާ	����iS{��ڐ}~�_ҙ��5��W=-FL��q;ή����2�A�օJ}�S���q��"��5�� �)�/[�����'�q����v��f���^c�%ISYn��
*���y�Њ:���-�S�{{�z��{�yi��̴8�tp؍�5�+�]X���N����7��b�;��{K�D~��-�Ӎ�l7�?
2c��3�)�]}6�;QƖ���g9ݖe�'b�CNVt[�&�ɭF�ܭ��b��SNIMƌR=�c�窊�{���,!y�#�2wT*=K�u���1�~����<�3Q�����V�u����OGK���!����^[g�R��<t�=����2��;�|y4��[+9��l��ݍb�^�s�m�5�Ӌg��w�Q���{i(�>��ng�ٙ��e��\�Z:��}���Y�^��ډ#Ѫ�%�7���T"�Xq=��U$5ey̧��/����6\�y��5z%㎊@��i�j�)@�����kM7�46<�zOY��Y��=�*�y�r�vΤ˛��k��g�Jut�4�ř��Q��~����:�w�U�嵊e�^�N��J�)�S�g0V��H�r��J��p��m[��ʧ���lܝz����L�$��˾�a��k|%��v˸;I��!w��	ˉP[nq��S<����.:�Ѕ";��ԕ�$��K���$rQ��V��cY���ѝ�p�7�ܽ�q�AY�a�,����&�Q�K��BK�V�J;�gt�B�%$A��(ZI�R�U�j#���l��7�h��ٚQ�AG#ܦ�(wc�L6�5 ��Iw���mLMe���d�:K�Ķ��n�̙.����kZ�D���6�n$u uJ�kh^+�.l��Չ�U�t���l���|�l���&��ή�c��#`���Հ�R4�L9�P���o��gS<�f�WgkVh�Bs��֛ǟs=B� �i�f��{��َ���Tަ���2��ήL<����n.5d)A����_\Ud9���,L�@��ɋpT,*��y3���-���z�%@y\�{N�p0����ډ�h��8rų�_'>���wk��THf@R�+3���S9��x�����*�tL5�ݼ��̋9���l�λW((݄x�(S76U�&2���o4,��.V^��L3��o�N�
�f�T&e���"5Pܮ�Q&�}�;����7�9r����=r�ne$U�rw�s�p�
�e+s4c�"�v_k�\���>��Kq�Qs؍AZ�Dk�b��	�'�o`2R�'`�éb#q@��p�h
�s�3),�:�[9(��V�؅1L����O���28��Hs���bbM���e/����b ��*t��+�8�����f3tw�X�˻���H8�{�Y���ɩZ�,X2�%�B�a�2��d��F.�2��8��\&��e��mM�ږ�W���n����zc&s*�T��\u%���L�C�voV^eL� �e+X)�9Y˜Fx��s�?����� fd�+�:��R"��P�M�՘�0!!K�N��q���2F$ ���0��-e0Up[^��pd �p�<Z��aB����ƕ�����`1%%$X�cm)2��H� Žݾ�G͕@q�QȘ�\& �IHJ9r � -�ݽČ�Ui֒�$b�L*� ��X �" 	���傄��9ԁ �)� ,�[LJD ���(8�����{��b�"
Fse0U'V�bR%]v�� QA6�1��f�wq BY��n6�j�*�UH� ,-��FF ���@��5G%�a�5���v0D�.Ua+�❮?#�Ÿ�����F�h���F�l�+9�M+�[���)BUi)A��I)ߤq��/��:�FC��HET�n)b'�jI����11z�>�|j���c�΁y�N�uEi^��x��U���A�r��G�sf5і���|���ron�]&�����i*E�r�p��t��$��P�i�Ǣ+j�%g�zkQ���`���dחi*n��6��̕n���ҖC�Y���'*��O{}��Na~ٛ�3��ƪVj�v�p��jE���&��Yj���Z�m/=���z���n쓟pyzm��=qv�'!��y�/}Ɍ�x� ׼�l:�7�����Z�8˅lC�i�{�i�Gz��\�p՝Ɨ�ub�QV�[��Jrb����t'��VA�R��eu�k�n%yg�Ū�5�r�%��q	g�y;p�b6`��qc�\�u��Y6����(˹��\��~���>�<�S!��Ul�s#d^u�(]�J�=w:o�Co�6$F����ՕQ|�.z�N����*�E���#/ǧ:D����>Y:2W����=>��3$l�����`�*��	�vحN��0D�+���F.i9]ob��e�I��iU�S;HTh[\��cM8��J�^�s���0�zQA8���V��$�*���+u��dpԱ���B��]&ZHF?�Y�s}ѻ+יE���U����Y%���\85�6Ќz�\�7��F����'S̕]*�����=M����׋��ԇ�ʈe-A%4fi�Џ*y��Y��wsŔkn�9m�<6�R��|r[k&#�����	ud�$
Xfo�&�`�5���'�KV�0Ng�)��۠F��ܾ�d�]�4b(�J�}ġ?�Tf�Y��^/٩b�P�E[���)ǽ��S:Z��&�"�1Gg><a�*]��v�e�T�\rc,<\T��K�Eot�o;y٬��gv�fΕ�ܐ�r=��>�'�WQ��{N龷�b�-f��R��[X�xw�3ǧ9�v���]��}��3JSxಞ^��#��!��m���?T��ɼ�{����R�{qZU骵	��)_S��j$���.UZ��]�>֫��_�$iE,�Y������g<=^�QK�!�|�ڐ}+��#+��I�8U2�v�����ʼ��JB׼m�V��/Rt ��*4��3�A'Y�k
�z�]]�*����X���3/:�����C�ڂ�>ݙ�O.]0��3�e@�Y��s��MX��uEy���1�W=��kSjt����AY�h���C.6��p�Z���4�3��N���H.���^�3(���4�U��y������n����/J��We���̚�<�ka����2���[?���MS��Q��#����&w�zQ�{�,����,��2l�m��y⩶yzJ數��\lׇydG��5�U�` #�)�j^Q=�Ӻ�u��uQ8���W��HڼAl��ң����}�6l����m�{9���7���N�`�y�HS)s�,x��r�>��u��9f�r1��X�+��r�f���>�`�7҄����^Z1��{&~"��ч�m` ��2��λ�
}�y�:h��`ǽ�� ]����N�Z��[��w��9ެEȰt`b����ve̠rrZ��y�����]��9����)qbC�9�	զ�~���'�J�K�y�,��7�6&�x^����y��,[�y�����t-�r"�s�uh~�#2�Gp���x�|6�I�g�Kuq��M\`�V� ;^�9�[�s������ۨd@;�h��ݺ���M��=��[�U|������7۳��(��������WZ�4)�F�mgA���t��<o��皶ORέǝ�a�֯�*�~y�G��w��x����;ܕF�1f���8X�v���Ef�\��pk�;[����$���k�/�v�B��Q�Fs����:�be��@1Qi�n���eXwʅ&�Z_����r��Ê�1����hy�N[uɱ�(6B�+{�RT;�6��)�9(��ۛ�"=�&�~�z�[F�%*���Vr9;�wCG�֫��6�Ow�R\�(Ѵ��^^����yܖOtDQ��یCy�z��zٝ�-���:�T��U���������'��׏`����k	��'[HLN24�ӝIT>�<�#d^w�[��j�3����x��P��UF�'5>��1ǊD��n�bӇ������(.9�;�akC�[1v����I��V�!�YDW��뉡��Q,�#��!]���_XR��Ҩ%Q$L�zY����"�,�.H���WAгm�md���eֿ��O��e�_��=�B��݊�,��d�n�
�+Xp����k��wG���ʊ�-8���L��Ц�|AI�W�StCCׂ\�L�w��:⹍j����{!�P�*e����m�C����Fs�#ұ�&\r�O�u����C�>v��PLZPN�n�Z�-���XlDmM=�R��n���t�祆�noi*��p5�c��v�Du]D����"��Θى�UB�Yj�Ǘ��qr�j�V�d��&�eH��f�wZs58\=��b�2ݯ0�s>�2�xO~��WSu��Q�;��M�kB��6\c1bҝ�!��q����W;p�ʻ<K�\S������\��4O[��9}���:��wz�QP�������VVTP�V���M�Yψ�u���1��QFs� ��aۇ�Ւ&�|� A�2��3h^z�S7�VJ���ܯ ����]�������C�d���3�P�#��(��Q}0�nD��H�y�x�N.�ܾ:����	=oq���'fak�[xv�U�2�`!�P3]�F�m�e�>����h�T[�Qw��R����gjaj�䞴��nfsFX�y5������x�6#ͼNe���'#'�,��|�{���G����z7���F]��7�n�z�**e����*�VU�5`�_՜9ͅ�n�/������Q���o=���s���Gx�ez.E��
��|�^�)�k���[��{0�T�eF��N"F;��V����9+�M���j�Q�H+UEFd��
��P���{�Q���Ǣ���ضua���ݚ�ܶ�u��� M]%yF�z������o�/;&������N�WI1"Zݱ��2�u�s�f-���nn��LO�� �ȱc�]%G<������z�x��Y�jب��*^1�^���-�W���I�Y�I�0vo�p��*pg�I��oGT�d�6^�r�����h���Q�'oYo{��jBp����'���l�h�Vк��CY
n�H'u��S�%�����]]轭��h�`��FfG]�Ŀ���{5Uѫ<�&�N+���h��.LNe۰�z�}Ѳ q�|�ӵ�X��m�q*�^��m�9�v���qtn8�Ȕ�R���f�1�L1w̧��r&��=�&oXy7��ܚ1�P�V��܋=}�=q��W���]c�|��k����8E?J�*א�u8�Tʙ�#d�jC9�b�]�u�n��'�h�K�,����=(�v�䰀�rW)�k
T�q����Co*+�<r(u��gOD���n{��b	�{7c��}��>⤢ʲ�\d�T���N����q���y�h��߹�����9.��S����~[��u�MFRf�V��DM7��Fٛ���25����Һe�^�X=gy��>��Q���A���e����;U����q���R����w�y,��v�ٶQ6�T!�u�)���[�ۊrq������ѭ�E+�zlԾU�|J�y�xW��{>�;>~��	�b8^fa�'g Y�w�������&f.�Al�m�2;����)��yg�<���ݭ�O�)CZ�el�?�������?�o�?�T!��*I!!$�d!B*"$�~�� @@O��HP��^����C�cE��M�,�5G��R\����v��jd���:B�A�P,X
D*��! R��U@�� Bŀ�UP(�)P*  �)*���]�k`�8�@Q � � ��@� @# �0@"I � ��@�B �F`��@�D�@�@�@�F @�@�@�@�@�FF�� H U��m�A(�m~,3����(<žZ$�����R��%'�����
�"H���R	!�N����g������B��}�p��:���B��������A��l?#�v��n�ŰX�ETO�$�I
Ѩ��JX,'S�[LpDD���Y�M��~�;S��h]�~H '�](�� H�!"����?�/��P����!�!?� Y>��.?���������l? ��²����TDM�ܿ�S�V��6����>�I�q�A��M��� �l���uA�o%�~v?��?��UE�p���VK@����?w����BH<����d��He�����Z�% �������Lt�E�B����A@PK�@'I{(7�@�"Q�EA�_6��k%6(0
5�X0~��7�7�2����%υ�p	���@$J 
TJ�@
@�0 >���~�>�p?���G�����?�C~v�!z�۔����D�}Tǐ�T� ¿e��,��CF�� S���~��h�A��G��4*�"`�k@G���ƿ�?C'��!�~�>����p��{G�u��`<��)`�D�g�Q�g�!�����d�G�����?0����C�T��������{>�� ���m���A�>�����C�f ���l,B�����(#T$�n *(��DD�����?ܡ�2\S�B�(O��������`^`3GׁZH"X��CG��� &G(}��D��Y�m����	�Q�#�����eO���V���.G�4X�T0O�?hCb�3��D.�����"���1r�`I��%������X>��<����DD��E�$����0)�~��`0~�����n�/���>��>��~�~j�>��B�'�}�_�zy�B��ϼ�
�,Н?TOڇ����	d��?��'���s����Q?�?~���>�8"QJB���/���u#��TDJG����c���� 8x�����x����������P�@�b@�,��?��\�YqlO��?���j��D?a��H�)�����?��$���a���������>��>�Q,~�~�?2�U���>�
����C�ݠ�����}�>)�	�衱�&�I����.�����iRK����� '����,~�,������?M�HC�������|�_��@A?������t8�i-��v�r̅ ۍ!���XO�Z�4�ڒ0�h(��	��?�������rE8P�y槗