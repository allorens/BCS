BZh91AY&SY�l&]�v_�`q����� ����bG~}@         _}}�lUTDh�6)��VƂ��(QRRU��k 
��e�a@��V�ґ��*V�-�l�U�eT�$�REQPR��%l����%j���Z5L�*6�-1F��e�-FmIlm��m��k-d��ض�H�A��ʭ��K
Q�E�F��XP@E
8��-��m�	�2d�)���u�ՙ��p7l+(,��$��̀�2�&�*��M��U�ERm�[mi�4��#fյ�2�S$���8k2i��  �R�����ը;�����ݪ�*�]���c&���cwv;����ۻSU����]�M�.��V��+)w:�S�Ulʹ�j"�[h�lo��� �( :�ީ@�(///x dZ,.���W�����R�^7���+���ހ�(w�x����m�=�Uj��X4�Zw�Rz�Uf�i--��"�[mkl�p  �:SCCۚ�� ��Q���ک{a�Ѽ>��f7۠4�͞<ES֩^˼���/K����YR�7��r�E�И�ǽ (
�{��A�7���ff�֣f���V׀ ��:���{/����؟oyݞ� �wOxT���{ҁ�ҩ������@g'� ���=��T����B���ot{�*(�z�h�llʡ�ډX�[m��J+�  �׀���[���
7���J����V�^�O{TU �{K�i_F�A���5lhB�((t���[�h�Jk�����vҳ"٥��6Em�Sd�  �� 
S�L�T����)�@Su;�����{�{�]5*�R�(F/pB��������.�UIJ��u�:��q4�4Ѷ��kT�U�j��  YP y�����8 *��1@ �.v�G` ݮ�ܸwgk ��p �
�� ж��6V�2El��   �o��Uaւ�N��Gc� h.�p���X �u�7 a��u�s� w\pP�.ڐѵ��j�����  �^ ��  ��� �N�:�؜
 -Kt�]�:.�p n�p@��� ����Lj,�Q�RZx   �� =u���@�Y�@ ��� v�� 
��� 	��P w�ht;n:(��   �  50T�RF�LLF`��1JT�� 	�  44�S�b�E       S��)IT�@d4�LCL� �&��jm�6SCOSL�MM�!) �(�(fB1� 0 z���<yۜ^��n|�|F1MZ`���-�gM'M0a��s\AU�4Ɣ�w( 
��׸D@U�"��_�(��1�$���=����SUO� ���EU����������!zHrTQ~�������d�?��x��2q��<a���2q���a�x��31�2q���c0q�0�<d�8x��^0q���d�x�<rq���e�x��0�c��a�'x��2q���d���a�8��2q��<`���a�'x��N2񓌼d㜼a�<a�x��2q�g��a�x��^2q���a�9�0�N2�<d�x��98Øx��2�<d�3q�2q���a�'8�����d�L�a�'8��N2q��<d�L�d�x��0�<d�L�d�8��2q��<d�'��2q��<d�8��2��a�8��N0񇌜d�`�8��N0�<d�'x�d�8��2q��<d�'x�����a�'x��2q��<b`�x��2q���`8���0��<`W�(�0��x�/�"<d���ʜ`0��x�/�
<eW� ` �9�0��Q�(�d���^2�x��Axȏ��`�
�^0�Tx�/3(<`W0�xʏ�*�a�(e`N0��xȏ� �`G���2#�P2��P�
�(�2��x�A�"<eG��^22'� �eG���2��x�/Q�<g2��DȼeG���2��x�Q� fD8��eG���2�U8�� <`�'��
<d�(�^0��xʏ 8�``�"�^2�xʏQ�(�aG��^2�x�/Q�(<aG���0��Tx�`N2��(�aG���0�xA� `�2�Dx��U� �e@�"<g2#�Ts
�`G�����`�*�i���d �*'Dx©�Ux�̊q�2��x�/�
<eG��0�
�e���0#�x¯�"<dG�0���`���^2 q�^2q��0�C�<a�'x��0f�d�'x��N2q��<d�`�8��2q��<`�8�f0d8�q��/�3'x��^2q��<d�'x��8��0�<`�8��N0q�N0񇌜a�'8��88Øx��0񓌜a�3q�2q���a�x��^0g�����a�x��0f�&d�'8��N2q���a��8��2q��<d�x��N6d�d�/8��2񃌓d�8��N0�<d�'�q�0�<a�8��0�2L<a�'x��0�9�2q��/x��3q�2`�|Ra�߽-iw�>���qi���-��H�.�ծ�CLt���ŷ�*���N��nV9��VRwD�"� F��ZfD�MѵEշ��4�{sYD7�L�2y�묧�H��5�_j7�h��>i)�����6�!�u�3)k7�����r^�*�1#m�+���tkv�+��T�[I���kn=���Co�0�=����s�� �*��%�א�`uy6�:�+oM3rk��t��R���汮P2�tQ�E��I��,il=&���3oSWk�켢~؍bHP�!	%�6����=�U�YiQpo��J�crȭQD˵�%�ͬm�ס��3��l�Z���ՊDq�n�iu<��I�l��6�DO�Ram-�&8AՕ�;oom�R�M������X�N^U��VK��SP�[����eݨ�Q�+?�d6u��!�ܽq
�B1PY����˥��Z)@Qh�m�zB�k뷀�M��:["ܺ�D-�����UAcr�:�(	P\[RK���ܴ�w�A�`:'0�)U�t��B�%�׍V�Ƣ�d��#�Âiߡ�V6̄c���J�ؙ�]AEM��ܬ�2��h�`�Ac��u�ۍ������^��w�G��E�y
�1���ES6
�s�j�}�x�g��Q�X��l�u�sn�gr�p�wQ�Yl=8�,h!@���G�˩�A���0C��e�2w2܁�Qw�!\ޔe��h�
�m�p�N��:�����ؗ��u�{�v݀���ѻ�K�Fa3�r�4ޛ��DU�!azm�u7Z�o
�w��t���ek9��I���ݱ����S;,�[-�6�DQ���9��B�9�1�	�(*ۭy>J�0��u3pU�JT�r@┍��cVj�Y�آ�;�
�&�����
ȬBen<�r8��yA!�wH&�Fw(fK��}vu	��V������^e�i�[)֬�&&oM���݆�r��1�F��w�L��eW���hܡ7kgAG>�nt�F�Y�)�т$�Yz[�Y{P!�b�齈RH]���kB.������h�-��BMm�L��	��*�3J� ��5�W{���˻ϋ�n�mXMia��v� ¶Zh�dוx`0����#Y�; ��:����:�L`����T��̭l�v�޼��vKTwc�8ne^�MM�!ZA��q�բ���d��R�m��Um�N`:i�W��X�I�WW�1PьV/�O-�,�[���z�dD�7X�*���!I����k5FdVN�ڲ4�7|���TJ���X���nnY�[��e���z�<D0I�ódl�7Vd۬����xf;z�Ŋ�S�[�h�Ք�r�֦�\V�mB� H��ח��N텧��v�7M��K�v�͔�X���Y����h1�v��c��*Ip�H֘̣Y{-��Ы��e�O^T ��ݻ�h/�ǘ�S�"ڽ$%��(�e�SXFPٺ���^��������+;�5Ь���cS�ตf̥���m<���`էt��ˎ��z���Zj��S!/kK�˹�I���!Y����;��2�SD�/B^��욳hUZT�4�yyM���49Xɽݷz"ʍ�*�x�V��M��%֜�c2��@�eIB�MR����-V�ݫZ�}���Z���,\V�Ga���cbQiD^�zq�ɀ�l��.�j=����bt�&6#IhUI�A@6U�x�3���fBI�T��&j� �43��)n��{LHj]��F�X�3*�I[G(��l@�7�1۹�<;Q�[[[�E���l���ƶMUD0�A�-�W��c3t�e\ݙI�ss$�!Q���N&f��7�؋!1ECZcM,V�ӣ6R��6NT����rV$M\,�	��i�ї��贛/5�5�,�r�=p�svfdm������(Č�o*�M�X��1{���:�D� �o5	D�<&��JG��92���h�B��1#BlQ�E�E<ӭP{dl�)^9R�85�h�i,T�-NV���9ּIד.�Y-�+�y��|Z̧ae��Mh7*��l�B��#)��0용5��m,4�C/��:�P�մb�3m��#�1�R�c�rj#!7+r�u�lӖT��-�ú]n����
�1���F5W{D�4rI����;�-'c��{-�x��r���$�����(��+t5��)�Xj��P�wiˍ-ٳ^�i�۔������-�Ȗ���B{f扚@3F�%&2��4� ���a��[����č�U,a��91�y���ȍͫ��@�k��p�Xky��7au��m&�>Į��,��xv;: ��⛎�$��iI����yb����y�Y��B]��ˎS��R���I�UG4;@T�7`5��N����3NKDa��U�l���x��-��`�Ul]�q\iŪ^eG.Z9��ky�/�Gr���v�Yܘ���W(�j���1	(^�F;���Z9ĺ���z�kI*���U��N�Y�G��B@wRՕ1�����[0E�i�Yj\U��^Ș���VAh��Y�SL�X��2���h}gX��2Β`���2c�J������Mb��\q^�r�r��W����,m��P��k���R{i�0�p�Ɩ`u���z�
@K��[�4���ۀ�%%bF:(C�3a�SI�^+J H&r���7H�*�l��V;�kVLak�)��&u�]-ou�r��,��I����Ւ�Y3E�XiP���ku�QZ�m��5�qm�Hݛ
̡���yp��m��D��]JP�ͭ���m͎���,��F����*6rM�%�]
{M����U�j��İ��C
��3e�DU,��C����X[հRd�Ec�(��ff8l�th��y��ދ�jz�����Q��U�r�St�1I���j#2�|ˬ�G)���YWȬ�\���a��������*�I�+ {������4�p)w�b'��n�V���Ba���u-eU�OK�&�{��͐�4�z�u4U%����	^⢕�k��õ��$p2n�&�co+7E=��+)�`�퍫$̭�
(1z%�zm��J�-GX,�Nm�"�+6���oqc{��B���0�§�7b�!)�胶��y1�ǻ��I��/V�0�n���5���6��W�T3�rX��ie�	��U���X{]�����:BXqJ�Nl�x+v]IF�M1���WsF���z.�p�\�U���P��A�JީS"˽�{Gdc��4�:il�Ӛ�>�̡w��E���z~!X�:��y�S�+t<	��EM�ٔ�Z�����=�S�#E�2����4�c��*8��	�����h��)L����y��\5wu �rTf�3,��T�	��[�^[N��;Q�n�`)�2�Ռ�6�ËsZzԗ״ �ˋr����	wwR:��!<���s�--�[tT|��`��2�{�.�����;p%�ǣi'X�ʝc)�t�	��E'���`Rxfrts�%Z�n fkȱ0�"��E��L{j��i�ʨ�e��ȳX�L�j���viJ��P; �3&M�K~��a�D`yR�n٘��y���Nǲ�Zocz7ka{M[�����b�ަ�k����miv��y����%����b�ےTH��YW�fe�[or��`S�s���*ݎ9D�a(֬-��q��-�f�Rm��m�[1�
��#�b�.��j�1�� ]�&�p��3f6kp#�����7݋��J�8͌�lZͶ+&�%-�2Gw4,���
�F�b�M�*�)��lܴ��?7�Zn[jhU�&+hJyZw��`Qt�]�.*"V��f�.|8���Y�t������˫w��c�,����բ�K�M@̕��C���3 7	ƞ�;U�����Y��=�WyN�pU�
�����Ά��tSr��ؚE�kٖY�N�ta����[ٰ�u���3�����iPf�xn��d��y�63�;� ݉-I,Gxس�iG�ظ��uzD��biU�HGyws3vJ��٨����/�n�	�*=u��,�kwr�=թ�ކ�V�DU�n��/�j3�̭�˧nC���S���]epn[��Ioix�m���_2{q����8X9cE�niES���u-�v�+I9
/�Ց�{T�-C�ZrV��ؕP4�ٶݭݺĭ�ߛn?�̼t�D�:��Kϑ6�a�F\�����,�F�&����N�G�oh^R�u��X��aUn��bն����V��{����)Q�B�n��ܸݰ0lĭ�Ů\o�d���=
Cv�<�d�5���P+F@��M��J�I�!P��> ���Y{3�m��41l������rň�ҠuW�mIy@�B^ٹ���2��1��t��V�֢\��靧!�+]��[��Y�N�{v��3&&����Ťʶ��D*�o*jK��Y����Be��rƴ�00��b��ѓo]�3wf̆P�L��wJ��#����P`O+�-����?�K[&��B�%�&
&�B��Ko�r&�U1Z,���eE�%��XF��C0�n0b���Y���d���0=�A�q;š9V���պM�@f����'7&���:���lݲfjp�oq�-���VŌ3Um#v�cB+��5Kd<N�m3�Z|�*�l��=k;�S��:�Ya�[�Kl���ZQ�wUee͊���m���b++,�m��)?���S�pѻ��lNT�f��Zj ��yKf��tΚp`;&<2�H��k،cD��Q�,�n���ݻۥ�-���CM�M��pt0�`{�3�.I�3r�	�
{��6��1�cb��cd.�Vd�p��G��"\m ��F�8P��Y�F:�x��a�!�fՐf&%�Ϯ�)H�E[���s)��(�2e�b�p�&,X+/�׬�-��{tw����2��{�/�h�������jR�#(��䛦�-��7]iOA�*��
!B�����K�ݼ�2#њ\�k�Z�z�|�����~Vo
K�tZ�Ym�Aٕ�0�Z4�;{��^^;O�F7���u4i��-.��6���,ۓ"8�3���<�J�yz�nٹbb��#�� �j�5`ܺ,�Xţ���Y��c6���ɪ΁L�D?��7D�%���E�a.��18j�fI��'��y3AeSˊ�2J��Q�)�8hU���%,k4c4���ELͩ��bEk��p�`��,c)��f<B���y��Y�a�a�LۘҌ���J�1�lDp�ׁ����U[��E-8*��l)<Cn�]�����m�����i)���I���*P���X�L�{�q	�ʺ��"m+y�x$5�V�QNU�Ҥ2\�j�����`5�!�!UsiI��32��핐�"���y�w3e��G�e�m�i����]��+^'�d�-���WE9QL�Q�Ӯ�.|v6�oFa)b���D2J\�*�=!��ꎪ��N�!��Z��pRw>�r��9.���M�)իX5|�0%m�]E����SC1ͣ2�B���ЁYX�)���M�x1}�2^�td�
;g;�SR���3B�P��-���U�̩2VFs)A�d�o-<ѵ
N�%��f�r��wɘ�f]nbݹ�n���xZ7+n�O�ճ��%�P!���y%��£���[�&Kɕi��\��ouaq0S�	9�T�XQ�%��ڿ�X�;@\�3Iߞ��],���(�гk#7`Μ=B+��##�^X�2Va�M9�A�A&ݲՍo.�Z�O�Q�6�i�W�,�T\�,�=(h��d�l���L�6x:� ��� ��Ś24r���ԣy�11YV(�3ٛg8�y�&�ph�u���\{Fj�U�6�V{�3��K�2㶜�����e=�D�Y��V�{3�zj�ۨ���j���lfT�2��Ҿ�i�-�!����`@^����0���Q��V�Tjigrh��:64���M�֑W34�>�ێ���f<�H�gi�y�2�Ő�&j��ɱ�۳�}��ֵ;��ᵓb�0�la�F�<I�;E|b܏tauJ֩Da��C��K�f�X�E�׌6�є�3'$�Y�&�LV�ͭH;S��ۮ@�P��J�T�M+T�ԓ+��i�֝�J�|��iv��yyn Vд�Ӈ'�zn��"�2�h�F�mV_W���5��|�$+Mꕇ`����H��6�E�[�D �H�Y���`�,��nk֨@p��Y�X��3��LUF@�R�7@���b�%Ba�Te�P?f�D2lI-�.27�+�����R���� �����ӏ&���P��i2����˵���&ZsUE6���+��a�� �M2f���7���F��^�{_���l}�Pa��&v�KЋ2c<���v�sO��>}����q�M6X��>��Z�Di����e��E{k�!�w��q�y׫���)�ڤ����5T�s��HZ�M:R#��)ke��n!Tô�{M����֥��E�
�VQ��9�B��]�U�=�ܚξ�m���b�7���?R;����;Li�f�2�,0�gk�[�ry�㤫Vr�E�N�C4��*::')!�(c���j�t�c��Me͗]�򝖆t�#c]K�������2 ��F�ye��� �q<�F��V��ѵJ�v^]2���⭔�bYJ�+`�
������IeX\�C��a����͊�[8�_��ف�<I�P*�Lȭ#b���8J$C���X�M��R�`�e�8�w���5hN�z���1ku.�=f�,��l�M�����&71���,S�]��ӎ0)�%	@���dz�"f)�>U�#�P@�'�peL��ښ��`�2!�����Mm7��5�M�3�s��_n�k�罧*j�?^
�d��_ʀ=��?���T��vK��M���/h�L���Qc�����c� �u�R|��.�z
TF���[V��L朷�S
��ݠ���p�z٥@h���ʀ-��n���"���o�$�|�ԛc9]���u�����4�}r�m�Ԋ������q�%��׻�;ģl�x3O*�L�=�tM,�Dwm7���\�h7��Gr:�c�G]FN����2>�۠pK�rN�ݞ�n�\�f��|��=�ϻe�W��������}�J��.d�2L�Cm�O�
�z(l��&�/-/�l��֢�$+5Npj�W{��Z�w�V�P�-謭*��n�f����p���k�-�nV��lś%ۗ0���i?�b���wt�1�[�ĭ�
�}3:��\T;���Pt�F�H��/�B��6�*����D	h����[&�R� |��˳���tֶ��]7U��g�Ej�y�:x1X=b3p�@t��������t.I;\2q�В�D�6�j���םl!�RB�	����q����8	T�TӡmN��V)	U�����*/2�u(�n��zOko��S52�#=��ٙB=)И!�ٜ�鲪`δ����Dy�W:%�1�K<�i[
B{���Y��'ełm9�M��v.ዚ-�7o{���9�.�Q��,'^���]yN:Mi�6[@�Ml��(l�]Xl��F��*�LwZ�Kn2��>/G*�S�9�4��D�j��u�Ay��}��A�7 ���C�e�a�O�h�ݜ��OGI(݉@��o3m9f�I�<��w,ފ�ޞЛ�ŵ!{b�A77���I�o���g"߂(&�L�&���Uwl,�M��Z�0)�:H>N0qݵ��Rd����F��i���݇IˮV/%nl�Ը��3q�4��c��3�QɗF��T̜rb��\��<n9XWL�l���'���6B�4Kǐ���ng*ᘆ��[t��`�e�#ThB����U��ڢ�]w����Rpq�떹d�0滅X�.�jut9㖷��U�,�q,�u.g��k���u5۠Q⍪��̚l8�B�f�ݒ(����@6�d�&�Fú�ɵ+<��ܯ����c&;���?�m�kK�Ζ+lE1��.�)��u���	�X���Q��d��O� �����E����swJ,gb5r��l����w��a����"s7VZ�tՑ֌�+Tx�34}i�w\M��N)e�7/S�qշ��U�GMֱEcUm2�G��I!8��|X�Bb8hD�EK�����sr�8%�7�4��cVQe%Z�ͨ~��\�榓Zr�L0��f�p=Y�.yr�IK1���Ao��xS�U:"�2\���'U�-!���a0��v/2'-��tk7{��Z�w*)Xl�R��UvC���㭽$[�����WZq��8;/t3��M�j]5�/��w*��"wrY��]�AY��۝S%V,;4�{/iADo���(a۬�l�������/McS�[νz��]��Mt�b�ۍo=�)���+L�x�U�2U�'p�f1�.rp�;��Q�02v��髒���;�ˌK'`�q�-Z7�lh����gc)+���r�)鼖§��eiz��I*�� 4JSɖ�q�EIr��^�v3#D�34*q�����Y��on��qQϷ������=F�%Ԥ��˞���}�f�he2�uJo�� �;��.�3�3�ۈݶ��mq�OH�gt�p��ah�,^��
����Ó�coU�T���K�22�W��&��N�%,VE7��N�,�����7\���Elj�ՠ՜�7Lw�����t�@h�z�C�F��{���M��p7�m�t�����ZÌ��$֩��ڷjt���ٗWu���5]ͫ�I
3&ڄl��w]:��7+�/���͕�.�}+(tcn(��=�9���R�났�6�����y�܏�n�l��;�B���������l�T��9"�\���F�؎�F;;������ЦV�E����#Ϗ`y����T�� �E��1_�ҽ�N#������N���z(<�u�&�Ԣ�_<�W�A����U}X��1������OLY�4U":)�M-c)�V�0j�� ��p�q��.��-�&;˓�������܇R�R	%���pw�:OeGQ/�D9�z�8��\h�q��l�0�3��z�;�e �-�n�<Ρ�=�E�6r�E�sg+�&&�X˱ո#G���:�jC'`n��rhM��Ei�ˑJ�W��Ѫ��6���[�̖�`:�"��dH&X�j췉D�^�5v|��!��w���E4e�2�YCUu�$n[��Nq\����d�m�V1�DI�s6���\V
O�ssF;���.m��\��;�;j�z^�;y�wU?���c�]f�K��he��f�a�r�p+1E�s��z�j�T�0�TvJ�["5�V�uE��ã�c���-$c�];J�ɴ�V��He���Gk���j�Ew�X���Q���YST�֕��u�qۧ*W�#fڑb�b�7NjG��n)Z�:��跐�S����q���ӧ�j�[o~��ك����JZ���ݡ�kۯeWxՈ7�p���Z�O��E�ӛ[O��7�p�c�uy"	g�&pZ��1�x�rܬZm-�ݢ�_`�[��Y���M�l3I;N�׮l���໓�~��`S�J�y��фw)CL_e��4�܎fpA��8X���]�<w�%��>�N���V����:Z����M���x��h4qh�:z�3���v)u���͋R�ۂf,ôca�؆ŋ���v2�vY��0e5��SGFU��׳�c#��3�6�%��b<�CZt}�S�+X�$U�a��r3n���B�F���2��u2�^
���R�l���Wmc�����z�-�����J�d��˚J��m����̼bۑݰjïzM
G}z�y-t�o�e�t�;Nc�|by�Ō�ʓN�nh��f�+��3P׳����q��q�<�ac�2��W� ��3X6�]�e�y���*=�_X�;glon!�fc�d���I� $��ur��j�n�ٽ2�W��!;_���ZA���y2�꼘��1����F�{M��w�$r��wm�])��ww��Wut��]�Ty��޲��KX\:>�IjYw\�쀛|h�pEu�iҽ�B�(�r��%'qz@����t/R�k���W�ٚ� +h+��#(a8m�n�'t�n;Z#����6R�ܨq\��mʸ�� Ɨ�l���[��u����t�#!�DoE�lo�W����*�R����h3��)�ʠ�"��a�����e�Ȫ��{ֶ�pF��x+w��c����>�Ԅ�Y����ش��:�s�K�����ݢ�b�YX�q�_l����
gҥ��SЪ9Vw5�8m>�jXi�u�,�]�W��:���o}qK�E�%�|@nl�\ZZ�5�0�L�����(���g"��K�Iѻ�t��m�p��3�8�G�JK��5������J7:ȤZ�/wQm���W�M���OzM��j�N5,Z�ٛ�CJ9R�*io��>���V���nG&�.��͔q�[���v�1+�;��t�G�	t����D,���N64z�B�`��OF�g)c�]�=��dY$��d�M��%��9:B���D��|��-�6]-���Թ\]��*�͍��,�]$Q�����p§wEp?�k8X�yՂ�G;U�FU!��.^�z��쇖�OOkV�u�u���	Cw��ي�U�}����Gd��w�Gr�sݎ,Yf��EXE�
��f��H��Pm5�1�Ԛ����1T�aҊK�pٽ��4�K��o]��8�k�;H���-�X��J[N�i.���D� ���S�:��n�W��θ¶��6֗M�4����2������a��̉tj�|�n�H��
z�
n�ZH=�j3N�\�81K��т�w[K-�`l#�j�΍��R3z��/N�G�8�E�ݥ�W��̏gqS�nZށsˤX��������❶j)��t�]��C�������5���rl��_SmqF�u�JA8'i�����5�%Y��-�j��{1YO��R�-!��JΖ�Y�<Be��aJcٴq��%�wx��[��h��	�;V�y���I��$�<�씢JK����*[N2l�O}��5$��c���.9n�u��0m���ʎ��77_]c02��˺)M�iAeJ˓����ю��d�$�\��^�t�m7Y��;oH���A�6��0\;�K���kkDKU��\3We����!����)Sw�%3���/�Z�n�ھ�2��s�:fs&�]�.l]6��d�$�5G��P㇮b+,�7�7;��z�M�+�jtK��
�_4����^`ֻs0�^���eK �e@�k8�7M�ZGJA��PN�T����=�>�J�RV'Y�v6�����r�A��Nٚ�fZ��]@�}�g��vp�Q�����n��S/�04/�4y�����ϧ3�]6������g���"y� ��(���[�ZcB�U�6c��E]��OSǵ6���/���t9�@�
�,�3u������:�V<��ݹM�a�ef�
]N��]u�}��iʎ�d���p��s;n2��3kr�nm��"�BT�������y���{	D$z`���Xؑ�Eڧ�醺���T��D�	��wI���=kk�ԼY��Z���*�ci|��^�	������7J��e��u���q�.�_d9Y��ׯ���:��(�s+D��,3�я��U�	�C�Es�8��g�R7V�8$[[8h�,��W%��u����U�5�8�BV�6��@Y�;.'�7�F��Z�F�JZm(��lnV��E��:т��!���0�����5�7`����k�t[�ٸL�|m�n����� ����(C/V3��s�n
����-f^٠$�f��J�ݳx��}i����u�U�CF�²��xFn'�Q��&D�3}��ycP��"!��T�����}z��Z<��'n��P����3���2q\�2���C�*K�9��ޚ��v��ev�p=}鷡$�v�E:��m����	Bj[�syt�m9:�M��L�Pӗ �3�ᨏc�L�L�����&+�Cy��l���S�zG̀i&dܮ�O�N�7;n�zTj�O^m�ܝ��wW�yBn��+y�Y��'bWN�S�KNgϞK3��.��⠏+�����9ij��va������1�2om�aM�ܤ��K%v)�Dt��M�y3g36������DN&�_n���8�4n��Mssa�N�[1.�ul��2�k.#ǖYN`���$����Ĵ��0��4 ��e#�Z�;���E��0+'`XDv�_��c���>�Y�5�ˣ�oWuŦ2�\�H�t��.���Z�e������<u6�'k��a�2=��s�"8$�1�nY�$��qWi���ae�z���B����Bl`��3X��*>oBOEP���,4�J�IZɅV�狸!Q�|Vlu}5�g':N�`���/7q���qm�v��T�S�:mLwN�\#��v"Mgu�^�P�������\�tM}p^�¸�o9q�Yъ����wg[wvt�w�S�%�}�u8!�S�/���������]�	�"�cx���QlH�t2���y �i���[���ne)ə�[DCb�d��D4m"8Tu'i��ђ�?��øQ�^;��"8xu��]�6�^P��3��a�����CL2�����:h?b¨X^�m9ttp�[��7�r*�����l�|:�lc��YO�"�(�GT�Y���TPȭ�=㍰��A�3jܚ+Z3zm,�D�%/sy`�bGo��9���[6�B����	��a��l��W��t�۩�1'Y\0�,�᱅s�Y:��jWYe"��(��{��R���(�݆��:�������I�$�&��:���P̼Nԧ�iڶ���:�N:�fn�B�ك�tM��:SZ�c�vf�`��f�n�+u)b�J=䶫f�R'�����T�C
H��1�!h&c�9`���(𪗥��l�]���-	"1��8�%Ed#Ӂ�ź%-i5I�,�B�2d/"�#�ɲ��i�*P�t���n��)CJ
e��M���US*M%X�
�h�2�ME,�N��ni��(�c���)
���Ay�wn�$v�m����mEH�2"�P�Jmϧ��Z�Bȍ}�E0i�R@X%��)_W�]6���V�iۼ��T-�Gu�������IB&��T�4i��ZN�Zeʎ�:� i���#�t��m���V��[tF҆HZ&�َ,<j �� `�����@@j�$,4�X�܈���ʺ��Ê
e��LBz�V�f����QX�2�ǕO�hI��I�O��f"?&�$3$')񫺌$��q�*(��n������7fn(	e�!+6^!Y2}�Z	�*�&p�0���ir�e)tR&FM(Bp�6\���'U\d&�!WT!R��B)�ֱY�d��I��Z�ޠ"
<7��5PQ��wS[
~<MUA�çC�=��0o����zVy�1{q�津k3��W4��Z�}yʆ+U��^L�N	�r�")�Y�CvWCNt�ѻ�챓"ȍ��ݫ����-Aȑ0piV��zi��} �"f톪+�oi����ۗ�=�#�V��0p�k�v3u"�役S!޽v[�IJ��y� b�*�8D�ܨ�a0��H��U�,�cj�6e��3���9V�- 4�L�͜F�]�B�u*Y��+`rqv��,<lu��O%���}3��uθY4J�h܌��-w�L���\�+��W$�V��K��u��r*��^|��}U���P�ꮥ{����rki�&�_G�����U;���S+������]�ѓ�Zw)���6��``��u��;`m��[ߡC�3[t�V��/$t��Ύ�t6��
��\�Ӡ�*RI�r�;��'^�7�B�S�ɝ+�����""�bGQ��aQ�2��[+�8��1�a���&��]�����\��q�4�eZU�2v��hnF��`T�S��e�N`Gt7t΍�؁���x5�Ra����ae\�Cz�n��t뗴إ6!.�/��K�':�T�!7��IU��\C�8��0f��2�Nf���:z�[�Ϸ�����ׯ^�z�z��ׯ^�z�z�^�z��ׯǯ\��ׯ^����ׯ�~=z����ׯ�z����ׯ^�=z���ǯ���������ׯ�z����ׯ^�=z��ׯ��^�|z��ׯ�^�z����ׯ_�z����׮z��ׯ^��fz��ׯ^�~�g�^�z����׮z��ׯ^�޿\�~�_��������=z��ׯ_o^�x����ݬ���*$g|Y=�L'Y���=LE2��8�������\%�n�ؠ7ϘF`�.
��3u��nL�]2�:8z�_�S��5��G�Cg'sQ�
�E� y����9R�4��yR-w��U 	���7[��+���P��^;��!�̻�՝�T�͟�!��<FgU��ĵ��:�e�SƱu��`G ��Ps��"m)�}�%P��z��L��-�bf ��Q�ʼ"Wa� a`�1�{�������0���RGXn���2�a��	cJ�3e\v���c������:��7�&�^L;���{/>#�,�v��u��I-m� E�wrb�����uk+{9��w颮(D9;�F��#mN�t4ͨ7��Kq̥��6��09B��Գu����1aɥv���#���n��������5�&� R�рN���qȥ$EM�2C-�7S;z,�F��k6f*�J��Oc��0��hٮ�����H�:��t<r�9���C|�wx�8���D�e�`壊T�^���%��D���>morp���l��T��fF�Ӻ>�X�ޗ`c�m�6��㪽�wAq�*�\*�!Y�Ԇ`+Y+��s9+ƩvhUhS��`k�t-�?� ���|�w|��|}�oǏ��ׯ^�޽z�^�z�����z��ׯ^�~��z��ׯ^�z=z��ׯ^�z�z��ׯ^�z�z�^�z��||||z��ׯ^�^�z��ׯ_�Y�ׯ^�z����=z��ׯ^�~�g�^�z����׮z��ׯ_O^�z�����^�z������ׯ^�z��ףׯ^�z����?_������z����ׯ^�z��ףׯ_~}��ϗ�F��w���T��`�w�}���Xy�4�c#���VR!�k�շ���4j��}O�QI[��to�;	�Y��ڽ��n�E+O[szVP��t8�ܯS'T����KL,*WԒ�7{eD�5�bQ�dfmE�)g'�� �!�'S箕�����V�5�t��5�jH?��ֳh�שv
z�H}s����[+�ku��e�uytIkY�m�H�c��Q�w�'���C/����q��f������E,�I��[�4ӣ��qÜ(��[��\%n�t�X�:R/��Ze�T-�b���H�;�Bk=Z����W�(���X��edM7ΰ ��u(z.��6�z���,��و������{8�B��4S��Dv�,ޡ��8]A1�C̶Q�nL�UZ6�M�T/o:�f�;��u�V��J��U,n���c�5��	�c;��g��C	�;7[ڳ�����w���c�K�LY�-(NW1E������wM�r�L��
]y�
�l,(� z�����g�u\\���;H�3�F�P�T�"�$��٤�}��b,��"�����շ���:3d�^A���ѕ��!	�2�fm��i�ٹw��`:%�D��}z��]�E�����z�~�zϷ�^�z��ׯ_O^�z���ׯ_�z����ׯ^=z��ׯ��^�x��ׯ^�޽z�^�z����׮z���������ׯ^�޽z�^�z����׮z��ׯ^��g�^�z����׬��ׯ^�z�z=z��ׯ^�~�g�G�^�}=z���ׯ^�|z��ׯ��^�x��ׯ_O�����|~�_�^���z��ׯ^�z�z���>���Y�j�u�8�NI�J ޚ�!}2��4�I��㣧��e�
�#4�;c���N幼��{ί��&��	����0���J��W��=�Z��e�˝�G5Zk��J�1�qm�|� �g2�KX���@9�1��"ڼ �N�=��SV��!���W�k~��g��-�]��z�H^<�r��`�>�NL��}rn&���U�p�\2q�P�" �[k^^b�v�N����QQ��{*���[{y�õ��2�;�X�[c�W*�u�7��)&Ж�޻G����S�w��k��73"Sa�j���B������E��3��e��omc�9��9U��-��Gv�a���h
u�x�Ƅ�:���4���#��trc黭���E���\�k�>�W�������e��`4�G�=��u��v70Y�Dn��FgT�E��&K>G�b]�SG�x/Lʜ/J���{�l��u�f(3�����;��FMS�v��z�4��s���O�{�wJ��;钰nd�CnO�t::M����u�+�����J�ąnU�B�.)-��St,�:;x�����B���-�otKtH-b�Y��Օ������5C��DN0���S���>�a���Sr�g=��j��w�e��l�6�b�;Z�Ի:����e,�ʱ�3uV&���kX�\#+����P*�9G�������{�4���F��N���.�Jur0vt �����9>1 G�x/ �U�h��	��.dU�Қ!��1�!��d�Z-\��f���L�߷��2�h�2wK�[RwP@�hFF��W�rp�0LS��i/3#�b7[B�Q�oe�"鲱��M����w�J��wBo7/��Z���x`���;*u��_|�N+��g�d�������S�̺;dCجLw;A��m0�z#����V'_R���l��,��J-���4��X�-��yt p1ڿ��;v�M}���<�FS��ֺI��Z(t	h6x9��M�b�T>����f���"��(�	�((Գ��$e�]N�XW�K��"f����աzz�Ip�(E�
�:%����F�Xz�����G]�y�3��dyb�r?�� 7�`��z��jY�ּm�pMh����%���Gt��es��,���Z�PX(S��U�Wt������Z�V��
����� V�-Ji�Y\F�*���}#QK��ZBr&Ȭ��� ����J���@�!դ�TU5���B8<�1��e�3��GL��/�� �|A=ZWuA���+�kF:�BS�˪e���|l�+_	G�=�����L�G���&7���D�N޷���a�f��YYk��I��gu�0��[@���7:�z��O�]&2�s����8x��c�˅�_T����U;��,�m�����⁸V# ��1��f^�2R���W�Sͳ¢�MTF�����9J�O��]�K��H�U�C���,���)�[�9��c�n��.�k
uf��ms�(�-R#Ku�����[w�ZϷ_n�R�s���M�x�Q���by�"�E��:8�`��Ԉ�c)��%��D)�[%���l���!�[oS�>�WZ�'{wE.C����P��'z�\]�N�1)�]":�e6>����'AC�����Rn�R�� ��r.u��3)b�� !�2Z��6Z�EFwo��o�Z��S���� PQ�̬)f�ʘ zvMDn�q8k��.�kv��uT�S�{��KM-8���8e�h����5�dwȜѮ������]s�.V�V;��<�m]��2mUj��\��G����qJtE��Inutx���f�͆�����!�T���Ҝyr���ZD�ƇC΁�1sm*ޢ�V�r��]փ��/�7��yjfopr>ѫ\ł��
�!�ˍ��Q�-�~��W[�@��$���]�Q��zK+��w,�rS'��z�=Mܓ^୭��|i�s�t$�X`0��-еq�f=ܣVi��]��z}��לW8)N���$9��F�����=\1�#v4`וtU'۟Sw�k�YZ���D+8���j3�yA���y��|[�����k�W�}X+�ܾ�Elݮ��f�x�Jv�x*E:-\���C��U0���H�^I-��W%j���� �T��d�u3.M�W1ؠJ��]u!�p2��.��q&��r���;�vV�d��o3r�㒘�M���>NY�$���C�U;�B�#h6N8�=/k��G]ŕ���yx����z�cW�;0�d,���,m�l�n�q\=��M�ԶN��q��zFoa�f}�8;鮺j�ؖ�ƾӫ�s�5Sko����T$��%�F�qx.8��Ձx钤8+Kn�a��d�쀟���ohh@WC�GE��Nto�|0��V�.Џka�a��̊1Z"��G�:��w��o,Ō�}���':��!j<E��W7%g%9��S^j*V�B��*y�fbͫ�!Jz벙2��{:���>�=��04��I��֩�Zh��+�FőY�Ã;T:�	�R�T��6a}��s��� (���q����;]��Y���,�Gu��Zޭ�%�]����oX����Z$|sCލfXr�~�<yq��+b�'xsI��h��<��Y�Y$�}[� {qP���s�LҶE���|(��b�L�&���*c��� +Y݂gi.����,_9�n�Z�aJ����:ոUۦ�mmC\�0Ss8���zE�q;VT�[
v�o
��d�Rs��0u+��P*�Wlv*��P;IRBB�Ū�ޓ�X:7�K:#}Z�*.ޑ]�3-�����S�)��G_d�r�<beB�Z�u쬸i�]�w�񺱛|��L�D�l�u��ev7/+2v��[
����h kڊM�/�8��\ݫ��L��޳������u�q��ب+b� ��_G3f��0�S����4�oK��<[�t���+����Fi���p;߭^A����,L<�ط>����U��X1]G�W�6�U�s�': �D��2���:�����+id��v�2�/������5�r��֭�	�ikw0�dH��ޝ�n�&9����"�ֺ�j���Z�i���>V5�m
��\�̇�i�nTH��)�g/�܃��VH7��1L+f��mQ�
�4�q�9����A�����-��;��M�s"�ҝ��U�7�����T�tvk��1�׳���!���򔝄3��x��t'��G��\��>�`��7�o=�S�^�69Ǝ�+R��$Ṓ�B��R���7/*�D\�m�(F�Z暽n�p�l*z���|�ީ̪��ǧB�Շi&�����Eն�zr{��} r�-A&��)[m�\��Hu���:ܰ{�0zVlQ\h�)�o��Ō���q&�f�9a�� �*7�G�^T�[+�6빌#�鱐��YK�Ʊ�Uӝ���ڤ�.:BgN��I��ۚ���	-��7��\��Y�S��rKLY��$�jVkSTs�nֳ�#}��4u�ޮ�b#k��pB(�����{�S˧԰-�;������L�|�o�d��Π�Ӫ��"km�q�j�JtW��ԫq����)W��t�Z<+ga��]���E�g 9���c(J��b麃���;�:Lh��3�-\O�u��<��M{K�.�G�悡�(T���P
}r+*�,�����vc\N�{��qpn���[��huf�9�n���wc�)��Ae1���k�9vz��=���a�������w�L�G��kh�i�T�,9�4�W;fL$��胫��T�i�u,+��d�%�Ԥ8嶅���t{8U<;��#7��@�`K�؃P�aM��(�ʆ���g&]��ٷL�>Lr'g�]�9�ے�O����;s>
�т}�%�sf��R�Y�}c$�kr�*6�,[��[�B���Y�5�U�T�z``�FnI�v��Ǽ��f�(���Ŏ����3����j�RPmKO��$� ж��{��Mk���w	ww�4cET��*�t�����Hђ��HX���(���ug���L�J}��x�u_9/�F�w*M�Y�������i�؀���em�0'����U��<U]��k0U�u]�ڱ��w���<Y窄&�s�@椚��[Rd&�&;)�G�d�lJt�u�Q�:��8� �5���c,]�I=���Ҳm�����;���󴻺̓)S�ú>�&.'�ĩK2�RɗVj�r;F�����M�4s}�;�n���ӛ�u���n��]�IN)ض�������ĥY��HRA�8(��f����N( �7}lõ.v�	�����k�-\�?rg���+(��^�=b=�qj��� �$�$�ZΎ]w��v�x(�+r71%�Pѱ������A�dkj
ww�k���땮�A=�;�ʏl����[Lf���`ͭ�Һ����꘥84����쭰�*�U�@�b,��%X\�x���8����<�!qQ�b`�����渥������{��V7��S41ev>ܚCdp�}ɗ�(~D�J��JZ
X��t��Yğǟ�䀀*��*}����O5�~�NԈ�:M$�i32�ZІ��6��b&f���$�.�J��4��1@���$cHv
c!$��_�'��Ki�ؼ���6]���;9!Ze'ݶ@�b����Њ]��Q����'tNRkz)zr]]b�'i!C1�塲.n����;W�8Ԙ9FK�v�a���5`��u�J}��B,�@�E��ث��s|f�.�Ob��TB=n�6j��x$8��v���.�GC i��Y��z����KM�K���Eyx���oN���V�S}B���񋋜��`\�;l��l)��-�6��0��m���n��T���5f��P}�A���8	�	7/�m��^����$��Zee��Ic�d�sks���:���ys3T�Gz�)'��M8E�7�մ/*]�{����9I����eVMsbѲ�wf��w"݊�H��nQ��M���]7wf=���f�d��1e�Hd���r7U��3,�t����N}�R�Y�f	"ʹ�"��%i#9i5
ڙ��_86PvXT�P;�++
\j(���FʷR�$t�L�Ğ��t�U�6$㋫�o�ز����R�JK��r�3�9�ueX�Hܜ�����eݸAL9���t��Ǚl�د�<�f�8�c싲YR�Ԗ��:��1�����|-<��w��j�b&HH6@�A
��;�f��)6�4�i&�1��nH��P��Iպ���K�Ƞ��c��J�E*"Lq5���][
�)SJVDA����byr��8q�gY�ۙ�k���ˑ\�l5D�آ
�����Q�9�������}>�����3�����<��kTv<�<��E��d��Uv(*��V�*���*������!��j���9�����}>�O������9�~��W�i�i*�wyS�墣F�7��b���~�h*�fڊ�b���b�9�
�9������?O��������9������cw9��5����3y�νc2|<܂}s{�߭UD�y��7�1QS����؊�s((�w�y�͓��G�8s�0��C�j�1Gk�|�����[g�n'	cY�bZ�M:4R�l�A"j��V��N��*�p����դ�"�����9i
S���7��h�hMiV�s��N�&�m��B��vֱ��*�Fm*p�Eʹm���F�	1�;��<��я.G.X��7�y<�z��FٵM�[M���6�?i f�(�H)� �H�	�Bi��a,��oPp�W��9�嫦�s�91Pz�DX�n��G�����W�i�Q\�6�s����62S�s�og�xa��\��<�㈢+Z�g��y�jX��X�8��yǋs��nA�y<��4`���xADV؈(׾b�*#��W�Z9����*����l$$�A-"$pDI�s�/��^cl����j��9j���Y����?]��o�����"d���{zk+}}+�"��:dn\a�2\Y��XWasw���־�a���5�ouy���$^*`��T"��  �\� i�O�3���
��/D�+D������	�^o�ϷK��m����|3��6?^x������m0s�̑Ի���f�Gp{mH/֓7<���}�s+{Q����8�d�粺��:Gd��`e�3��U��sV�4�'KC��7aj����>����3{P5�3`��8�8�C�ڔ��|;�?_��ӿ.��#�;z����T���=R��y�����L��~�ef^�;�"1�y�׫�1|淋��D�'/���*�O��[
�U���y��/[7���׳��>v�)�zs�g�2�,��ث�i&yL�{�����K��[��S��=;�������;m+�W�mf������P�%��tӈel�k���x���w�y^%�͇����=;7}�n]�\|}]�%����__����7��+�o=�����^9P,��mP�Z�,����=�Y����j���7R,���)=�Yr��1T�G�n,ys��z�^F��40�z��s�G�<�6ƃ"D^�(i����	����npC��q�e�OHK�o���տ4�艳�_W�W8���K˪�_?��u6���5��v{�彉�|��ze�U�7���e��{�j���?�����_!�"�
��7vD��+���j���귨��gѡ��}:	�5�B��M��)�r���ӽ��W����&}���E�C8J���'�*�`ã�3�q�㙇o��k�1���b,��]E�sD�:F���>�C������R��at���R��ϼ|���OG�:j������+i���i;�{E��W���"��d]�m�=�Lo@7]Lf�Duq#��h�7�^�Nd�:v�{��*Mꢾ^+1�/����}�[����i?>����;"�=F$ؙ'z�>qg{�L�y,z������U����q�U�-n�&���ˤ�0�]\���S�z��j��c���3[�O�VAv	���y���n���PM�z�����b�s��Rȹ)�M֜�KZ��&�xh��57Jnz˺^=�z�ޔ�6�E��%ga�͐kڱ��ㆁm�X\y�{��YyrPB�YHRN'����¹d�c�-��y}�F�U��o�����=���Ne��M�����a��	R�r�y8{p?gyߔڒ���X��{�G��zwZ �=^��<i�NP�fn=$W68�˾^ܞ~�����҅�S�|ۡ�1W�u���0���o#�F��W��K��xN��;�޳��qW�8�9�l�=��{='��L�dц�U<O6��FEX� »�g޼U>��;��L�(�2�_`�.�;2��C$�Z��-�=A����|�mH�c�YY����Do����Ar��ez��˲��g����VR������^yk�k
uK����7�gY�~�^�����RxA�6yeP�YS��h��5;{.fԞٿ��^��w��;�����{Ζ�|��P����f}��i���4���w���S�}�6G��ꭖk����=4�L������?a���ɟo�>��k��-w����^�ц"�>"�A���.�o������X#xe�6�6ۭ9�r�2�mb��.J�/G��T1��gf�p>�"fx门{t�rWIK7��Ca�h�2n���3�uu��].����wjvDr qV��yR~���e��@o�Byh{����Q��|V�3bb�� �_�M�+����y��c�v#�{@�o���e�?�^I�~ȓ���:}�වj��{��5��z�o���'�پ���)o̦3������l�)�/��~�_��-�4=ƺV�w|�zÈ'	��d
�;l/N�<�u�:����w���QeG�_����{�>^�/���� *���f��ͻ�����],G���^�]z63�>�b��q�o���?�_mo� ��wO=���`��(_�=���T�OM���m^�qx��9�:�����C�v����)�[��گzON�c�+(�V��_y�N`z��������쩍x��į8��!NQ�ܰ	0;�F�6<�9����5��42��y�8O�$�v�ɀ�ٜk;����L]u�/�t&��m*&��J�6�͌���un�.�b��Fp��)R���~��w���uj��Όu7�K�[��3�D۬/?N���;�L��%,��;���T�;��D��wb)w�g2����,<{�'rǫ�N:�P�����0��ںLf��POkue�%�/F����e����L>-i-��x���F|MZe�`�R���-N��o��8�#Yċ��������Ʋ,���Ve8������%%�pZ��_��z{�޿m_�)u�����b��|�=~���A����xemr����Xc7��� |���za7���]���R Z�->ъ�����zK����W�2�Ca�՟�Q���wbz/�+ӛ-X#I���1��.��զ�I�l"�|��W��U�K��=�w�Uy=n�C��6�I#~��9����j�y�u������L�d�:�z�ɶ�LB\�^��}rm�:��_�ߎ�J�ڮ��|�'�՞J2��n06G���S�ހ�d��pEOy�^����sO�.tl���z��PU�wv��SJ�Nd�r�?8�݂�/�Lʎ��}���l�V��؝�:t�p�!�y� ��P����&��[�vz�'�L3�,���s��9S��^�T�j\Z]���b����{�z�6{��<RY.fʾe��a��cu	�hf0�j훲���E�]��|�e�k�{YM��N���j�m<�n��-�3�å�Ĕ1l��ⓂW��Cs�j���'�p!����
�3-Z%������x��l�Iq�tl���t8wd�u�%��@���]��q!��2)�깥oޤk��s��U&z����{��^{>��w�f�&M�7�[�g��Uz�������*�8~����ߗW�g��h����>�«�3��3���H���Q�N����{���p���x��I�15�^y<{�����X�@�0����o��<�Yyo�W��w&2owiKz�U��/��h�߱��g~邕{�.�����O\j�]�����U��j�M���}����_"���D-v����=N�o����GXN��X��j�k_�Fw8z�o�?c
����m��SR�=�x�{��o�Ho뛪��u/]$�w�*W�K�p�lG��U�˚0�� e�c��i��^C7���~[�+�'��m�������~�d�(��`�G�(z�G�^�R�P$PC��,����f�8�mq��l���\y���av��]�]������o)�mJ-�ܛ7An�6�%컃��Y�R����M�Gy2.T�U}�[��tq��}�<D�P|��u��5F&w�5�G��l[7L�<�U�����b2�Qц�;��ʯfሱ	������,�'z?;��g{�]z�mq�����'7�j�
s"��0�N�MʰMl��l�1�ꞩ{�F�e��LOr����=
�[5I���G�~�0�n>#�+v���B H[n�xvA\��0ߎ�GoW���]�q�&���	�ͱb��7+�G�X��U�|���	���y�swZ�O>�x�4NU�3F�:Z�q��N��TZ�YN�?\P�l�y��\|N�Σ���c�Ryl����q�{�=�����/8���oX-繽���Kf�[��G.ON����ho�����i���
����X=�_�{�3O�������#��[�ض{�{�lv�+)ͣ�w����},	���g,����z=��o�ئY�v�o�o��dX��
u��k/�C!���Ve�tp׽HTCvX����y9�^[��[~\�}إ஥I/zjS$�CUg<�3^�97em'I���a�f�j�>г�hv��8�d$��zQ�s�
߾��{5[������~���1�R���>��}�y�����}f��hg���R�^�Fz�|2�~5��9�󩏱�|7����6�a��9�.�{;��(��\
|ѱ6~ϕx�4���A�k��w�@���0ite{�ԙ�h�t����-E~�t����3�!���;z7�y<w��;4d����E�����o��Y�����1*k�ك4�F�`r�o������''h�7��e��`��w��~�ߺ��//���a�v��~���s����:�y` `�=����Ѓ�k��}޷�_�^������ü �N>�x'	9�,�Y[�X�Q�"}O�a�g/EuS�r��S�eY� =�5ut�n�νD�v�cY{3 ��K�Y�;2�������f8n����ps�v���tb)(�o��Pկ��u{ۭ���E�^}�����7˛e�0C�iUꇠ ^en������4`_sY'ى�t�ۥ�nU�@��w�<�����{��k\�Yb[���˛ĺGkV�C��1��>���?Z ��E���BɄ�.}_|>+��s@:��䃙�G�~�g�{���Y�#��|�56��^6X�:h��Ό'�����k��{��>�h��a��j�i��sw,�:���""Oi��T&��Q1��o����eU���o����=e�N�u��O$����)�.���mUR���������UP]��Jץ�z|��7=y��g��_�P�ʂ��7�e_�o��N>7�'�pzFi�|='}�hz3���0_O��ͭ{�M��^�=�!�yΞ��9=�ޜN!��9��}�;�f���9q���u���@�ۧ3���sX�ho���g<VQ�� ���s�`���u���$:C����������~��Þ|-��g�:C:�w�̼8�Ǘo�KK�r�������)���0v�W��O9�������u:-�K޳vxz�A[�%��e1L1�8�-\���[��:_^}teɽy�5:
��/�n7�����R1u_$��/�?�
���B�.���c<w�78Ϲ��]>�ag*��s0�7�̝BhN��i�[�c��z%�ވ�ֱ����G���-;4n�w[i��;�Mwy��竳~u;�����
��[Oo�(��Ӝl�����L-�O/�9^Πo�op��;����n;O�7�Di�9��&���OWw��
Sz��y�*V�Kp=����֥�{�ǽD���}9�������'�'G#��ns���肛��ݏ��ڨ_g1��~y��]�O}���Eq�����t�7d�<�_���}ph���Q�麟�����9����b�;�{�%mد:�{����8���//Xg3 x4�=9T�}o�u�>�y.�r�3��:�l�G��[W~_/���]ة��X�/��ǕAq=��pb��ة9��㛜�窜Oח'��@�,տ���i��x�|3�Qp%W={�z���=�c�k Δ��s\�ғx��H5���!�,��o���
�2�v���?�u�Ǚ�S|:�m��N���#��h�X,���;kij���+��3Qn�PV]�(�T4iK>kX�k7ZН�[�@�)���i��8�	װ�o
�����c�aT�W\��jceΈ>����<���& %�)��U���bF��u&�.���� So\y|h��%Ø���$���v��@n�p�u���]z�G�6-m{n}¸��Or�GL��
P�u�H��Y&1���Ius�8q�|�l�hތ}���$�pQ����F����S;�_�:]>�����Wr�a�iѺn���n���T���S!kl�l�3��\`9CF���*����Eg!�o�ᚯ�g5�J�c3�)<����i�ȏ۫!�˽R�ձ�w�rkV����-���b]=V��6�UM�s�{]N�+��R�h",�:�3����;�Naf\��j�jI����4���2�7̜�;���t��,e�rb�Տ�N��)�;g�â��)!��ohv����Մ��܌���,R�e7Y>�lC0^�v��љ��+7�u�L��mg�C�%����8�=�N��\�F�]	��%TKe,wO�у�m}�Y�N.��%�ʅ]��̳�4��[�؇Uh���jB�Vi�g�,S��5��g�2,?���뜑����)�Cee��Z��i��rp͊:�5ӆƆ��Wd=Ɓ�q:yn�(�n�:ő��`Y���[���3Z�Z���d�����c�ڶ�[Y�����,�e��1�Q42fGέ����<�8�e���{mm���I����2螙��XS�4K�P��4��s��=�FY��	����T��Aeɠ�y����XF���9q�X���N#�Ȏ>��]jx��δ�[y�A�"/Bᐻ�]�y5�`�*�	z�Ϝԕ(7�o_|xJ�/0�W_jE=��̚����8	u�m�T�2o���z��{O��/�AA���s�^-�"O��G�FTNYjq����[�.����� ��O�K�w)�8R�2U�Ob`�:�E���'f�#����L�`���ˤ�Y̧���`����~ږ�st[0�.��lGu�r��]�� C�읆5�.�7��a��pK���U���8��H��Ln�n�����RB�`%���/�xQ4oYu���b�03��o+!�݄Z"�`��5i��-���{�U8@�T�C��D�D}�U����4��η��u
�3�y�qk�kKṚI�	����ے*A͛.��F�4�$�������g5�G|��^:����7�.�GMQǖ��%����E�>�k.V\T����Xr��7B�H���I�<yW�u���7��*��,F��r���=��
�i���"���8z�1����<�z�U�|~9�����~>�o�����������j��yȈ��\?n6�Y���8����cS^�TDG0h*��ƞa�V���p��v�۷u]Xue���*�(����N4c�|��b(֨Ӫ��Zy��p��5�\�i�((�Ϸ�o�����}��o���?���~��wNF�wnr�L�G��=G�h��:���[+cTUlj��|ܵ��Ch���(&��mJ%	��?<�`�M��yq)b-n�EIs��?.�,z�U�δQW���UT��Z�٣EEATQ�h��z��U[�lTD1D UDDZѹ�͵�SF΢
���F���UE0�ͩ(��	���KDO��b��Dl�Վp��p�Q��&*b�""�Z��cm��E�b����Z(�3RU�{�nj�����nr�4b"�*�)��(����q1TDQL5y�Ey:�8"䜎h����ȿ~����V�\��8�Õ+��زY<�E��R��N�+5��6�g}s'ЪOFn𥚳�����;�aN�g��Z�@x�-�c?8k[=������'����YẈ�(��~�i�d&�ىSgI�|p9����=���q~�f�ܚ�C�rF���@���%M�^3u	��Y�yk�/�W9������j0�1����.�z���������zv��)�ʹ	�a�ƛ7H�G-�ܹ��M�{�"���}l��9��M<xN��ĵ�#��SQ���cxt�>�P��ޚ�����Z��13����='W����deo�[y����|��G�\d��������5�o(B3(���["����@2j��d݁\����+k�T�z@��Ό3c��ˑ�"�P-�y���ћ��R���mD��׎�����QM���ȦԢ����!�6�8�AeP�e�n:�sТo`dn+���w�,��]��A�>���Py�t7��pzOچ��|��������d��n�˞Y�yS�ar����{94&+�z_���U�0���"�*���<c�Y���NO2�x��c�w�������5vg���r)J����}M�S8����x`Wq��YP�EOHx���`�Q;W�˒ϔG�Z�ӷ�%^��T�u��q�"ڝ�i�1�ީ+����i7�pS�tѺśaհ\6Ld�C[J�lR�z���0�N5\�E��2�,�G!����e"�m�pO�V���^�����ߧ��G�<�{9����e!�eї{��՟{�ޓPnc��-���51����8��g�̮������R���nu9�g&.VC�=�ßA7�\�����{p&>C�\6~�D�a`gw�l`����ź��p��S{G�A����7S�7>@��]��	��{6�_{���=���_p%.ϛ����������\��r�su>0
\�C��33?�������o���[J��B�T0��=y=��m���J���������)��{.�;3��9����CY�ǭ��<z�1���ۓ6\JD#E��V��f���}��Xh�Gť��y��Q�[U�p��5�����P��������< ��ym͇��ފ×
�XǗ���Hbv�J�圢[���MQg�r~�~8���<㆘�xu�3Aq��1����.Ks�{�<��z#��`f�F��)��3ϹM��\�'���ST
�Џ�>����BZ�f��v��tW���Q����Y���_޴�6H6]�5����u�qIV;�w�Y=c�	�[�ޝ�BHu�k{5�!Q��c�M�q�q�t�Vb��+o�ְ�m~��y݋oC&��{�ȿ�΀��l�u*�)�Y�Î�;ק�����6����qk�w$�0��v�.Q��'^7�����D��/0��O1����6q;��i�椕w�k��s3��3UMmX�;�wgK��Ӡ�wu�Z���Ȩft��!I%4�(R| 1���h��M������������}���@��u�=>xR+�ܘ[��$��ɀX�-E'�;�/_�Tf��wWR"��L����1�6��{�b"��v]A���n ��S������/Z6 g�nljz�����R����������}������}��O�w9��Vڦ g��\CH�����a��h��lN�z�My0���j��=a��W���@ǟ�_�r*|7d���~lo[PwƉt˞�����	܎�~�L�WA�M�8���:�F�x:��,4���sR�vtH��
��+УZ	����b�C�/O������ǢG��zrm�����-��_��EP�N��~S��	ts���I�zv��s�y�C�v��'�9�̴*�A�t ���P�u���%�7��c�� 8�8�T'�� �q���|����ӂ�}GZ�1޷&��&����f��� �����p���P0	��X�J���~�~�CP�5�?4�Hi~�����B������L�(�����/���`����  4}B���'���f���3�SN�����:����,�|t:�K{�hC����vmz�Ck�cc�2p1�:��Ȍ�h~Jں��Hld���ޤί؇U�i�c�%����Z�^�yrV�m�f�iNط4aTAY]�j�J0�� ��Nr�6]��Xk�W��>���}�.~�-���{;yP����v�J��|]\��ٜ��no]�]�"��iq�Xr�Vn�<��{�`�	����P��?����]�����8^[�Q�M���|���d��7,�gg�8"��4ʍ��}م�M���7)���tv/��L4�6~`,�sc����%�w�������
�n�?�uoȈ���h��8����T~�VG��D�n?5ߒ�,�\�Uˇ��(l�Z�y?3 ����~��.�� ��斡 $�.9�j)���U�qnD �$q��P*�S{�5ix\�,m�07#3F�#�|5bc�M��T~F�6l���QD34Ǉ9���Mڶ];�?u�pO̲�3sx)�����5��V�����
�P����|fmO��]���[ �KՅ0�[ �i��G	�-;Z���E�ęl�ւ���ז�IL��Fe��[ Sm%u��EFdǅ㺨����jEЈ�M��TdV��:�ާ�>�Ϟ�$j|'z;���K��ZU)����y�x�ⰹ�S8�1���$C"�v�4^\��6�2�s; �P��-zC��4��+�@��/�bӁm`���[׹�� �=a��t3[�����z�ͯ]��M�ޙ.Z��s� ��S����/�i�	Tq�:�9�Y���YF��g�����X�ۉ˺��GE��{	�0Kڛ�+������+N�[c[��A��^��]��97���c��4vp�+Ճf��s&���vG�8����96ک�cA�j�v3/�n����T���S;y�FE]*RcuϷR�~�3��3���y�����������=���#�Q��ϼ�P��¡��6���k�Z�	i�y�v@M�N�]֤�6b�ۙS=��#M!���nR�>u�|6��	��@�|t�5���TS��Q-�"3���H�'����v�����K"KI�
aC��Tk@)�z�`0hsϠ�� ?�U��`q�$$>T�*^�暴��W��]A�i�h��0>�=�s~���zB�����������i���X@hw��7e����HnB���HP���Ɍn�3�hoH�[a������).0��D_���_]L�1W�gv$�[ e���SR����Ҫ��#X��=~�[k	j+�M��	�Զ���[����b�� 8��@���s��g�/��n�!���ݻÔ �Kw�&��f����Cj����^�o,ϝ�r��Χ��6~��!��2{����N��`�>ſ��2ږ�|�C��=���<�J#Y��4���;+[�yE�F��b���mö1��_���lQ��v��A~'ݾ�V0z�|�Z�oB�40��K&�eM�
�X�!ရΐ�"��G���U�W5O2JB�[Q�o���mCP��]��˧�KRۮ$�$������x.���і�4ǈ�.�s���'��g�/�ɚ�|��0;�N��p|�S��4@N{u��%@��+��x���d���Q)Z�f��NS��[w����T|*�C� �GĐ������	��1�.���>ce�k"���3��$�;"����jgԦ��Ɔ�w�KN�T��̵��v��ט/-a�M����E��c	��⟥R���&&�P��6�Y����.���B�ޗ���I�a�������T6�	��= �'۟G3\l�hħY��?��/I�5�c
h��$�u�g-�BYj۠lN�d~�� �!�1��^�0Z��f�B/��/�\�Ŀ�����s��p)�۹
�Ȭ�^���1�e����й�̛��D���?3�EE���1HSv?Bt���w{vQ��H�d����)��i 	6���{�;�2�5y+�۪�e�]S��*�B�j�a��:О����p��1�_ס�]񙼉��W
��r��r9�3Ơ��
{d%�*1�>xF�7`�`���cP{.:�m��kqzh�ț�LZER幩��^wf����!�H�L�h6���{بn�E������0XlF`=�*�{���{��]�X���b#��D�`�k��Ϥwʄ
�:��͍���zF�N6��&�����)a�\Ρ<8PWϴ'�&�����t�
G#�]l�p��mq��Fk{mxO��{��!�H����4\GFG��B�0G�~��|s����cl�30S�5��]<�����k�|��}q��&\37��ǛՋ��Ε�D|+����r��/w^�?�����"�.���B!~���w���{�oݾ��;�F,��9�`��SW�E��}%:��8'�G�����8v��s��b�m>pѼ��3.J{\X�>.k�g,�䮃q�^�|���j��!�ȟFD�����9eOt몗�p2se�m���r�s�ƅ6�Fr�)�q>��U�}!�Zu��;=vb��}p+:��K��Q� �o[^:a��O�3�J�VZ��ت"��k��V����~�]�{�S�[@����5_~{�_�c����{����yO�.F<��S.�5O}׸ݒ��,���`���e�-�����\&,S��/^��7�RmsV8��D|���\�]Z	X�zٔ+�NK�c����L0<��Q���L� �f5P���O�Q��p�[΃��]'�Z��J_�:}Hݍ�3�1C�]<��G��-z��@�Ⱦ?�͎d�"�ng�����[�����.e�HyŴ�P��^�sR�ߵG7W����,LCy���+������l��d��:��)k^��|h.��5�B�~.'�mV��6\�3,�y��yl��<5f�P��G��S��![��Wz{}��V��̥��.Џ.��m�x�ǝ��\�+y���Z������lek��Ju'W[���~~«֦�ޡ#���}}1���ʼ�gv�5# �:�7L�&�LO4�J�{I]���)IIv��k���e�'��:�S�>�]M&4�P0�(PR4�KH%!@��������dd�C��[*�n	�O�S1����Q�;فM��
9�	�?p��D)5��p�a�uB�g%{��̋�n�t]��xP*K�~}�T��W�C�:���}��B	q[91=1~"<5������!�x��wE4'�;L�g=�9ƺaP��8­�W�c*��[��D���4'����8T�^Ͽxa����Q����	�(:�_�z�ʢ?�+8���G�C�ٙz�4��y�>���gV
�BO~��ʙkoX����c��}�4o4,�}��j�[��rz� �v�yϭc�e6�h�5���7Y�hO�C��\�c����4�����B����u�_Gަ*S������:7���(A��->>���=�(�톛����WuD9��a�z���<����<0�L%��)�|!4ǷÌ��m�w��5P-2W�w�<7/�������!�s�`D� �[� ���뼪������h�"��`��J�3�S7���D�j	V��UЬ g������>j�@)�l�l�t�e�V�Q�i��e5^��xW1���u�4^��9[�-ڡ�)1lu�d��ΛXwJ��B�e<49��5;:��z��]"���w2Ei{r
N'��Ć�,�4�CVZ�v�J�c#n�����o�{��_9m���g@�Ma�*HЅT�����37����"���zɛ�7�'��B��q*���Ͳ�ǹ�T_L
���N��ԋy�2�0Cu�k\)!lK����;>7�sח������t��SM��Sm�������N9S��1a��|r'mt#�2��vC�ܸ�_7�Dj��9�o;gE'�A?7W�����}��gUi\�;.���)w/��)۞��Ȗ����{EךR���΢}��Mw����?�5�ݜv'O܃W&f�eٓ��-~����y`Z��W�TO����B=T�g��g��g�=w|�$� #enoWaʔ:*Fr���ƙ[�5�hj
�9��_}/-�ɨ#sm��8j+m��2�0i��9��;��W��y�������C��|��O\��-P�4��A=~q���_s��
�e}:�czB����9=U�H+���-�P��}�X)p;�HQ����qH������S�WHڹ.*��1M���kվt�D'n�vkM���j��5�͇r}y�hm�x���VS����'�bo������#W;1Wdǽ�;ʹ6�t&������l�����Ky��)����E�/�,
�	��Y�GM}�/y�����R��;R����z�+7<�y��14;j�m̵s�]KnvنRvI�ϝ燐G�%Q!�t�e2���	2�*�% ��<0���_r�Yj���E�cּKL>p�?kH��B�/��~����YNo~������9���o����}戳���P(=��;D�D�� V�3ۢ���Ϫ)�v�X9&�1k��
L�����2�|�K���3k�*%��e;	�93����t�W�����[�	jG_rX]iguI��3��ٱ����A���&Z9eSl���;�r�2��d;�'�u���v7�����U韫�s.��{4z󺂰�q��Й'�b���� ��{0�/�W�exnejD2�Y�;�9'��_yA��Yn���
O��_�R/�Bblb�{��۹>F���v��V���%�,�������<��>\s4���v��u�a�R1���KnE�R�꫎�mUv���hsH6m�ž�H=�u����~LO��qߑ�([;&��vzhpӮ�Tt��p����������cÕ[�lݣ&�4ř#����q�4�K6�>�y5|��YM�'��Jw����`�맹�x�z\�/Oϻ���|�o�D��TA8oR���f���y]����T�Ɓ�\�U���2�;S4����n��Hr�3��X�VP��Fq�e+,��2؜����;�Iի;���;yq��k�q�}�����pC4W\k��;ۏ6���|�j�a����
��}�^7�,jj��Z{"
!�G�v:s[�T99t{ט8>J�շ�fi�)@��i�i7�f�Qbu�/I��9[�)����u���1����*�7נ�I���=��p�p�JD�2���t����)���t��K�g?k�5�7�y�mԫ _����T뭍���z��,�j8�D^
r�H!�/�zQsk4���J��T�d�.�$��\qi�Ӗ����yvM1���{t��s{&gsε��;&i5�]�ܗ�5��\� �_4���z�� yX���^q:9��E�q5]F�9��O��R�� :V
��ŮT{jاV4��=Aw$-i���&49¯o.���6L��k�����^�W�qnڻ�!�7��t=	�/���r�����e�[��ĕ�i=[����� ����2|f���*^oSI���/����:�k�m�[S�nU�[�K���5;Yʳ,9�7��L���jq��'� �1[���Wp
�L���) ���7������e��V��b�TǐS�%.�ޠ%��5oK����j�c ��=,Q��RQaݖ�`FH�N跺��G	��]��@���e]�T9r�"B��S[����'^Xt.�A�C(�5b�*�����)����lzQ������ �GmeFc2���V�`%=��SF=R֔�mZS�S�x��;R,R�3��U���1WDXk��m�P꾼Ǯ�'n��y��5X9��(>.!fU&
{�V���T�P�X��|N�B��S��ru<r��J�̮d]�NѡLmh<������VV��yќ��e��vC�o�N-5����2vqX�L���	�f��Թ��̂�G	�x�9\X��ӽc�J�}ffv����L�]t�*��8g;��o'd�LS��:��\n䃺o�8ݰ�Rgv�U���X��h7qWM"sM9}y7����Ov��ڍ�QTs�,�[}����nf�̆Dv�H'Y�qs\�>�E�iukU����sw,=�/XKb�l�gQ�ה�b����ԩ�b�{I���y�os�ΰf.;A���}��`igM�J����5(֛ϵ7��'�0�x��p��z���o(�o��4���S̵�g]��j8w"k�W+�%6&��x�3ؕ���q�\�6�g��Y��tݻ8v��� �]��\�0�oo3 q���g[�tݶ��]y[ur�頖b��vڵ�ƕ\�HZL�mmj�ŪnN��wgr@p��m3i�o��s]�ek߳+B�ϙ|6ܤq�6n���6]!}�8���@���^a�C2�NB容���@s�:��T&�ʩnC�6E#��B�(6cA�����8c2�4�
�i"	��m�,ȕ�����P��9�0;���Y/Z�]��
˶S@�e�$�a�?}y��HA)�������LŧUFڠ���7
��"�}������}?o�����z�g����l�b
��mb�Z�-*�(`��t�**�.~}<x��?�O�����}������?C�c�)����h�VuG6b"����mwz�z�""�Z�6w��<|}��ϧ����}�������ߓRU%�5�(�N��'�mh��5'��1y�{ǿ~���!QUk5DQl��)���Ӣ��.mTQ�w9�cCPT�b�j�����'�(���j� ��(�b٪���nN��b��т�/V|�UT�4EUUL��\Mm�"�j ���(��^��������cs�<��*�&"Z��\�S&�6�S��DE5�����7�l��1Z,i���QE�"j�m�I<έb�*&娃F�k��A6���� _���*���&Q�s�O�-��3!�;�̫�,���ޛx���r&!9/�����QKo
ź�Iw]XV��h��#.O��cmF��Q_�C����dB��e])Ja�*�4�P� ЍP��@��qＯ�M01����_�^y��r׽�9�/�����|��t��G���-W���m*��f���lvy�C�\��S�SE{^��L<åӌ�z�5Ѧ(?o������*h�5�W[um�	�J��tv����&;�`P#��}�א<�qT��L0�-b�t%���n�g&-��u���J�(!�_�?*�N�&'�\~a����!�)��_���Z�p���v���Urr<�{MK�P,6 UIj"��(���_��p�a۲~G����ћ����G��/ 	�h��+L&mz%��(��nQP꽣���&y����f\ܝߕ��g���Y+oH���h�@���I��8}H2�Ll��p�>�7$��5l��A�P��35]����t�`�3��w��.e枘���2���)��H����f�{���02�S��DY�î�w��ޝ�,�D(^��u�p�����>�����=���	��ջ�=�7�Gd\3�F򺇚��Y2�!�o]����k�*��l=���2[�8�����J�b��4՝�uU��Z7s����㷥��1��L ~WG��u���;� ��c�
uǍ�t��"�Q�u��5��>�'z����T�r�%�l�+s'=\V(nKN/��ee��e�uc!���GG	4!P�ܐ���uLsf�!�ӳb����� �F�.A��H% R#B�-��������3����a=ש){�������W��n�ͯV�(W,���|w�n+��q�C��B��4����z3E��Z�gy�a�d/���^�c��&*�~J=}�G,m�I�n��|�CƑO���j:�[]�n��P�o:9��Ih�� ީ-���&�Ҩ��+q>������EE��@���%��˨��{V�ġ(CŲ��C�硏;���M���ڮ`��˹�[���cMVsl��{�sLwz����8�hj�ʄ�e7X��ţB�T��oD|�|��l��!�D�,������V�T��=繆\�ڤ<7	�%�5 �)=L�?�*Y>G7��cNM@�\�a��
��:)����|A��r����ey��(���N����3����F��(���.�_��ݾ��/F[-!γ.fלp�Bk�g����H�M��P<C�tg��~LS��˧���Nn(���6��M����A����,���ʷ��{��8<���V9w�.ik-榹
5פB���<��ol���]�&ޚ�.}k�M����j���%� ���nvTM�epɗ�ztf��t�:c��f׶��6��[:.�x�kg��[f�&�����*��T'AXC1�2'<����V��Փ<�.��I�lgJ���Թٖ�������Y���I��/3��@��.��+��F��AB�:�y�^�31���w�O�O��O���Z�� 0�� �)�B�A)�v6�Dh�O�w���dkm��^�q�b+rx�����ʹ�U��K�M!3it�V��M�6OR*��:�˦F��v|�8�*�ylC�A_��_S,(�M`	��v�Th�V�����~�]
�3Cs}M)~$���ٲ��K5�B��:c�'k�'?�����n��l{��m��nuO���&���2T���P���`��}��g~�����
��޺���R���a�[`5����8�}%�w�ff0�|����G����m��c
�S��^^|�����S�nB'E�e�Hs���t��gdN�-�j~�.�\$����
W�ld[l�(9w�����L���ߺ.F?�G~�SG�l�	�[W�c�C4_tǚ5B��;��1���EAj�j���<SF�b�՘v��	0�ך�C*���쟚Cx�k�;*�<ޑz�%O.�<r*�!����t�=��� �Aפbۚ�/����
��z�|C��z ��+��xl5�����%�Tb+	t/2)�P;}=6T;��L�ƙ[�6|�44:;�}hD�]2\�v�ϗ���;.��<xd�S��Թ)+:/,���V���.��uwb>aȠ�0��a4N���!zn�T�ݸ�*��nˡ���ܧ�U�d�c(��\�l�hy�)Xf����6�-��r�c7#LA|�M�m�! �&deHЫE4	@% S@�T��-*>������Yp˚[�A3Lx������'+����x�Fr ������
f�졾��xK�Y�z8��X��ݮ��<b ������}����ߔ̼��B�b����?~�.��y��w�'j�n]}�k�:�D��>��yh���_l��(�կ����A�/��d4%MJ;-���++��
CC�4��n9�K�TV�6��ףt��s�-��V/UYJɫ��s�"e����C�W�gcj
��T�a/��0w������G�2�b��m����q; Thl�roK��J�
��t�*���15@�;}�8��u�N3,�b�����[ᓙ��'m�0��H݆/�S1zĶP�����-��=;�z�/F4����UV��FF��Jb�׮�Gq�j�� Ũ1,�l��c�y\��Sp�p����z�g���,�R��__;x��a�B�i��qT`&�=�ݡ��^��2�b�OֵS>~�s�a��B�$~y�t�t=b�r�e������T;`����X��)�U-|*Ǆ�`+�)S8����"/�ɸ�,���=!�C���́Z�۳��N�/�p�z���Cԧ]nY�t�V�����BHF��I ���"�'�0�
D��=�mTM%�_\���7�GuK�+ޱ.�G08c��M�	L�x���t��)�B�(�+�6�6>�q�n��O�r:��<�{�{���� �F](��\J�  �Ā��R�R-	JP4��	~sb+A�f���!1�F��j'&/�Ǧ��^ޯ9vOې���d3Eb5-ݥ�q���{�;�N�f ^��z�s��搬��&�Cw8��a�V��j+��,CC`��[�3�s��%V:�Z3��ƌt츷�D��s�`7�.�����CG��kH���y�ܧ���M������.�CvbT(����v�^��㞋�ܔŬ�K$^=�X�-�61��<[)D��uR��ڳ|�	�yTS�<���7���vM/�l�����1��痷�A-��=~��&��CǕ��,���ǋ#}�яI�BtȜܔ��O@���:�sK�Zv3Yɺ3�q֨�P���z�Z �Y�� Ѹ�h���ȇߤk�P�V����-��s�n�eҢ�cXi34��g�k�Yȕ����O���_3&S�kO�s3[r�Zpe�E^�|}�1��E1��$�@���kƿ�;�Y�H���S'zh��|<��sH}�
1�]�H�[�B;$�۠�[:��rC��*�L~����:��/	��t��Vt��D�^���N�r�X�L�D�_��;���1�f+�Z�]���[�U3�wu����ط��E�e�r�RRa9y�6U���a����r{�N��:��nj�@788oo=Qq�����ޮ��mΓ[�8�q]����!�E48eT�Q !H�*H#�~��^;������<�W���[]8�/��\sz�6�0��ߺ[J�-�OX���]�������{�o�o�a$h:��l2~�$�C��P��=۵�!�>�n�n�o�;���*�W�4�-g��Tã�v"!��q���y/�|l%O�ߔ��CMm�Й�E�]��zb�m���V��e�n+,�a>���׵��K�NY�����m����0�D�n6AM
�IMz�}ԧȫ;m���
���{�NK׭��SK�HE�2�|�.��R���X�`d�h�ލקْ�Ɋe��S�:�j������������q�$�KA��7��9��,��kF<7�t1����L��i��tԖ��ljSm�n��c�	��Ny����hk�Zw:�4�R�u�!������}�^E�+�Q����U�kH�dK�0jO��<&�Y{߶�g�h��W$�B�g��Z���o���=�hЪ�����7Pz�����vJ;�v:���e�/%%���\�W;�v|�1~sɵ��E�����y����k�i�l\��/�V�oq����dT�(�釧��&��ץP�Ś^�%
��s�b�83^k
�.��l��*2^��3�v���ߠ��x2K^�ajZfNY�9C���7�S|����Y1����z2�F�j��h]��>S�A�4�a�EGH Ѓ@޾w�����s�Ϝ��+�z���׶pW�i_w�/�<�;�&���d<��a"�_..\%��U[ԩ��Ƕ�s[!9��Ħ�Zw��Ƌ���	o�D��Dz��	�.h�a~�3�3����Jʕ��O^��u.ӐXT���u��~ZǮ�������z� ]��������k�=9��9�j��U`M�f�l�}ߪ��V���ߍ^���!Ca ��.��w-r- ����t����=�$t(H{{�3Q(�>u ;��7���7��RL�8�B?�s%;�;�:���^>k:����:��.�f*��y�r�� �� ��gaL�?�:�$NR����\%T�\5W�*q�ԧ|ڵ���f�JF0D�
�]oq\�?4��_���ߥ���O�w������O�n��Ul}l_�Y�\W�
muF%�^����S�jyY��U��d*�b�_�ʒ��ew�\��h����g-��)��2˜��l���0�e8�ځc5��ψh�֑sMO��
���!{���lw	�?r����_��]0�XJ�ò��x�;y>O��U�=�608-x/ƥFXw��ȕ�ݔ��~���0����?y4t���'�kIG��#�\*���9��@A�;�f������,�Z��Wnh&��tu+W����g5��+��;�,xp�:,e8e�mu�x2���:��Ͽzo�?�z�ZT���:p�.�(
!�@
�|	 |3{��w�\L�f�?>!��Y���?-����M _t����C��^�����i�H'��>��v�;��r������s���[��~K�/=g����R��܌���3L�rqJ�%��OoH���f������'|�;^B1m��\C��P�W�_TO����ﮤ;3��0k�1C��S�k�)��M*�QH�7-x?F��C���9��4�?ϼ�\��t��`i���Ys;Lv�X��&�EV��]�0������:Ĵð}�g���O�X�R�y����Oz�!���L��lLa�c�+��>"�>�R����B�=����_�s�iFW�t����aC�z��E���l1�a�q}�s�{D��^Ml�\���tt"}~���$)���X����7�?yE�j̟g��f6`.�!�ܡ�r�;[�]!M~�-#��.�B|�<��Hw����2���L[r��mz���c� �m�P��ə Ve;R���6Q2�1�ܖ*
�Q~S�4��>�I^(��!�����^�UlɎe�j?j�B�R�E��SR��-�=_���>d���@�e�b#G��ܗ�eiU��Š;�]�a'L[���]� %���;&s�t�)KΦ�ؽ�n�-#h�*ٖx�L<�dEˡ��5[9�-�)���;{�^r��r9�z�y�^G�5���Q�ʮ�0 iD� ��)P()
hU~�}���}>=i쭚��:�|Uy��ǰ�,�J�͋G����q���;m�_����^�ޚ�{��ѻI����S]�7��B��gA�v�q4ɻ)eSiW"tb���%�k�j�1�����]�/67S�NNl7�ws�Ǯ�L��b�O�Z]B۴pg��5���^'3�-B��L1V@�
)���v�o��>0���9�U-x��?k5a�e�ƲE^�lԀ�[4j����8������G�<ό5lx�C'ڋa<�"�C4�`�'��*���A��Y:���t`M��7+�L�t2�O��}�W`/���X"�<[|�rٺ�9�[��I��e��ôWl��{6��o�'���N��W�*?D��f[ �LX�w��ڍ]�Fjj�vk�.[���zN!��5��&��H�y[<5��;�t�S�r�y�W'v�6��mݝ�pd��c`��������"�Ȫ�j�a�25�9͏Vqq<����ٗݏ���5�m_���0Y^��CF5w8�Q�#u�q{�k�X�O���K�*�~�+w���kl��8��B��HZ4��WgW\��V8���;}^�~̚�w�>e���0��ut���EUEz�W�E皸Q��＊D�r�!gj�cn��6Hn���7֥��Fp"1ǆ�8�Ѷ$'x�/�yۺ̹��ݻ6��M�����?�#�VD`M
- ��A����x���8���A���n� ?.$?��8���0,�/ֺ�<��T5�&�:|k6/[W)��	>��S�D�ð)�N(>X�T���S�mx�;>��ؐ镵fr�j|�1��S�&kjD��v��x��^&F*ao���Bz�1N�L�͆vL?pUw�<ӘSd��6,`����U;��9s�ń��r̀%t@�5��ͪc�5=h�ʵ9Rۺ��|��^���@��-a�+ �j�,a�P�m#"[)t�;���꥞�;7ޘ��0��B#���T"-\
��y�����JV=��C(y�	������ك)�Zp�*�=��+������k��V���=q�:�;Vl7'��?D�R>�O7�#��魴#��wb(`W1�w'oZ�g^\�˜ۑ��..�\0��l��rsM%��X���__�����8���v�Xy�z�lgk~7w|���TE�ɵ�u�����(��kl^�O�w�qT!3��|r��>���>q��a�|Y[s��:[0�!��*�b���= �Pu���H���[�� 3���F`��w��!3��������z�Ⱦ75�T!b��5������v��pZz��r�=��r���\���PQs"�(����k,���+�n�� �����L�Sβ� 6U�1��r�$^t1T�E��̎�w.��$Ji�[}��,�6��C��$�,�U
0	˯71Z�`$�.Q��	�n���G�zj�)��s��:�%	��н�[��ֆ�]t��Paɧe	
<^C�i,���8�y����"/m
U��ѫ5������ ݹ��bp���y�C{���N�"�.�",����=�z�r6r�-<��wM�Uh���.6pN�̥g#�VU�\���W#�;��k�f+�P����g4���]��s�eּ���1��/TM�d+���Ki��c(u[�Z�.vN�y��u1k�S9�7U�U�x9��%`h�o'q9�2�C�b5hLn�u�u 3xn���	Cx��ߵ�j�&F��w.�"��q�V,Q���nƕ=6x�A�8ec<k���Nظ�ʸ��3��5+FVRç\���i�"r���u�l�۵���3,�$�v����+�{���r��".�R��s(�D��KN;ibn���MG^�򈼔�vr����o�6Y�uo˼B�O�	k3{[ޮ�R�pN�ԙ)EAv��}���T�{V$Q$���۸rA:�m�u?�MQr1IV����Q�|l��cf3]��¥l�rK��z����9jo�ٕӠ�ٽ� &h�ݸ�}�6]Z����t���E[�h�֛�S�����p\��1�Q�(Q�o�cfWQ�b�fr��[��g�f���F�ֿ���`�����搫�$���`�Μ��Y�����F��B�1I�b����D_iU�TVcGK�\��Sf��6/쇷��:4�Nɦ�`���gA���3���Od[Z�ɸ��j��#/��u�����ìN3�5�������qc�Y��6���{t���k�������B�����QA�3������JLf(���aV�ۭ�E���2��k��ޡVw ����9��{\�l�r�ך��{�ٱI�g�u�O8��z�\<+�:�c#��gh���'�Y@R�eY��2��y�8��{���Å	>�&���\ݸ2�[�:��-��I�9�w�-�&�r�)��lD�'f?�L�Ӎ���rco�$��Ρ�$-Y]�v�=�j�Z���}��N�@� ����:ܮ��ޘ/l�y��@��bSkЧs[������Yz�U.r�IF��Ḿ$Նe�Г����jI���G�$�~ ��-EZ�b�2�{�y¢�?F����O�����~>�o���?�����U�QSU\�o'y�d���!�'�D�D�ڭ�?>�����~>�O�������3�{�h��Z� Ѡ�����kURr�k���Q^l���珏�����}?o���?���׷袈���5��LAU:�E5zv��-SUUDET�+MLEy�AO2d�ӒJf��q\Ψ���h�׹t�j��Z��Dr6,p��8k;����r�#E͠���5yc��Tr�U͉�����ֶ��,QU̚jMjJ(֪��DT��r��#�`��i+�9���Q1�-y�T��j���lSQ�SQQTN�m��-��U@E^񨤡.1i�g14U���l���j�sU�;�����:�~~��Y���껃��1oRt9#���/*���\��3sX�՚�t���y��~]�>�����eP�A� a� rȫ�����ߞ�Ͽ/�7��z����|d�d�y�i�
0[��sR�li�n���*��Y�j���;���ye�������И���dH�3�ŃR��XIxֱ]��,4W��̰Q~�T�y(���w�-�3_0hv���D$�/�g�{T�q;qӬ���ʅ{�:b�<��\n(��ɏs���'_� ��:�#�����l�1	�������Sx�t�IuF=c
�z��;΋�"��/���=����)��3���#�6l*n���'�ky����ϊ��>c���k�tj/>��>�a|�7.�d��}৯C�l�+�#k�XF�K���,��A��Nc	��O���S-y��m~�,�O� �?>�D{�bx�K��1� qv��y�[��^����V(�;L����t��߶Qx��Z�����S
���P��9�:<.�;n9`>q�>��iǃ�ҹs���w�b�=�mߪ2/cG=IÀ�0ӿ���Hu�~TR������}�Y�F�"�����3��Z)9}�����t	5�j�%�Gfe=@�|{�8m.�'6#^y������21�����������k��u�ǻMMw�=p]	�^ֽ�5��)K_Ji�断4���0 0��T0�+�ZQB�D��ߝ��B�^�*�����C�ԉǧ\�"��خ��d��RѢ|g��� ��?8;�"��\���X�m�#��66i�s��՘�[eV7��W�/�C�3-vj�5�S^6l�K��msC(t�=t6Bh��HU���L�[�*��t3b�ωL�§vc<�k7OL�/�C�M��O��XZ��A��@��ݯ���d9�*{�>0��Ss������z�~���v1vѮZҹN6K�
iMs�W�T�B�&���W8�:�z���N��#zol�˵���
���&��T,v��������:��>�W���]��+���]Ѹg²��{�]�G2� �7Uߝ�5��7�l~�=_1q &޻{dHOL�WvC��SZ�2%��9�v@0��Q�آ�@խ26�>������]"��ݰ��}�jh�Z�K�r�/,Zc:h���&�ܖO��~�{�1c��+��N_��t�~7y���y��Hy�l,z]6�zO�01��9;;36X��i�!��RB�5����e�D��	���v6q޹���6�LV��l�;ۗEEGW��+[<�d����jY��J��� ���Hw�ek@�;�䮗)�B��ⴀ�s���tt��ڷ���˨�p�H^*�k���4���R��]�jX����
#�=�j4:��%U��3��2��O��MI�E�����D�
0��2 x3S��B(E{�n&]ޓ[�~ �owf���o5��0*B�׬v�3�=Ci�+�[xA߫���o������z�����R���ャGN�������@G���vÐ=O�o�<H���5�I��gM���8�@���R0\a��O]~���	��|�_�5��)��z��I�d���]L��Bzh���������L�����@F��׹ٵO���{�Ln�[��s�3���ش3#΄�z��[�г>�잷ܥ3k�f'u�Xh���  j����l��;aD�������v�7y�7�]NM0��ܸ��[� ň�ɲ��m���+mW,7L����/��:�xd�1؟;�mr܉w�qTs�*�oH��-�̙c׸2�O�\bf�Ry�ܤw2�b����7c�l��zki��H���*1��Q����}<չ8�&*탑�,3ýΫ�IAbl걝`d�i�r�:����0ϕz��'���tȷp�c|�����'s���]0
Qa�V�n�|�����$A�FwH��_��:�� �G:��6n4��KY\?\o�nC��&�S�f����wc�ϓ.iT�*Ǖ�"mo�����DN�Om�t��b���/��0~���7��-�Z�3q;9C���q�4aaT��)���uc{-fۈ;Yi8���=����O|����S�0!�S"��{�v����� ;X�F2����<1j8�0�T��8�<�˞�Lkm�X�5�>0�˔�Ev�㪋�����Y�Q:�Ľ����#	i�lo=v\�Mi,��,g�dIK���lhlw܌�'�v�[����C�hB	9疂�<b�>�^���TXmq�ZS߫6}`�z�K���V-�/
��_�_,pStL��yqd{�mx������l[-��.�E���m�Q����{����i��w�F�"��D�+|�����M�n��$����^�����V5��ͳr�X�_�l��/�kpK�^D�&������&��+U��D]��At�8�i�!��33��o2ֵp�X���4۽_����n1О��.���w���S��;�-]���V/�&�T�y`?`�JOo�bߟ��@��f�U�i�5��a/\��Pap��1߻:�|���y�S���*U�f��dE�v�,a�ܡ$���9����E�l�3���e0�:&���f`��h�6"=���j�d�S��TS�S�d��O���7ќw��<�������K-���c�0�uuCPΧ�"����eb�o# ��w�wk�i_ja�@�9�$��H'���rR�/,�%tɊ�uzû�9d�)��%�+$�\*��ٸ�U��񩻰|�"{mcf�}�1�Kc��7������=�s���@���2&@����������zݻ�Ye]�Ư�ܱ{�3�_�6�%��Vo>
�>���'R*��8i)�m�x��z�ܑ�v�ضZ��Ǟ���~[�6���O�]��j�f�u X~?m;(����9^�W�Y�JI��:�m�a8�ˠ
�>ޙ)��-�'�`��]b����P�S1�V��%�=�ty��*�MWq�[]�����47x�Ky�2�3V(2��rz�2��J}�H卿I�ɂ25؍z�Y�2�n:�������ًCU�wR�2�pY0���oL�<'�Q�_�J�\:.3��7�eT�aٞkö�1� B�ǧp�^l8M��'@^�,���s��1�;�z��~��U�s�(�a'b�Ϧ�-I�0������F�m����?����li�R�,�#�<�����_)e��b�p�3�i8�w`%%���s�C��������%��=�#��k+W~sߝe�a��m�S��E]y��MGx�
D��cOyB���D��4����\��v�;�5;J�lX��#1c�����ݹ�;`�)���]{��>�I� ��]T|~��^��3�@��WwO��:�:�ݼlU��:�:�_@٪4ev��w!nS5b\����_+�p ;��-�g�#{��2�J7�m�S`xg��MZ�5�ۙFl�[��]�ު�*�&oZ�%��Y[�}��<���&�� �1�PJ J������y��4z���?�*,"g���)�Q���+�s�f�ƨ�d�Ó;WW�o���[���C�'����d ��"d�9=���,�7<ə�Y���0A	�w��L����?�~���3�Q~YѦ�P�]�!b/���Jy����p��g\z9`|�;��\:J46�-!�����Պ����6�/������F�3S�GP�wa۳y���_P��o��`�A��}޺��v(&~�ڂ��|�6q��,h��Ͳu��b�uf="Y��c:��k+����=��:����bS킧ڕ]
�bʈy�f����QS�Ww�GN����=	t|�dֶ�x ���qT�v��L���~��
�Q�?l�;S�������T�^�t35J�Ǹl��8L����&�Wy�Q%ؼL7�T��8�y�c�l��en�݈4�v)�g}��\cL��h���C����(��WHy�k����	���J�_J���X]1\��	�nJ�7	P��
�h�#���i�`��Ҽ|���*A�A����2�+���s��)zyẅ́��'hU4��n�d�5c�Zg�1N�%U:��k�#�G�d�6�����,����w 	nMZ�l�u+0=&�L�bc:y�q��dv�g�G������l~��|ʦ����C�gn	:WA�"R��¤[_R�O<8zڹ˞�X���G� C(� ����o��w���9��Q�Ջ�Ϭ~��^EW'�Q̺ʚ�i��_���}�3�z�)g,��(�0:]��oeu��,rb��τ��m�(I��d��5H��6^���ʟ5�rw�[v�j�6�Qq��/%�T����D���C�u�Q�v��:��Uc��.͛&�9S�����1�d7�C�%Ṱ��zN�������SMv��6p����3W����ǦZC�f���8�:��[�b���ʆ ����L :ŕ�)�qSn95K�=2���������lOҼ�y���#�ϓ'��,W=�{��vm���Q��D]��w(e��Q���sY- ��SeϚ�.a���G��6���~�t�\���s��!����j��0�fC�ga�^�6��*xz�ӮvmS�:�S���cJ�Um{=ί{2�_V�6!L����z�TS/3?���b�#��b�5�eC	�� �ƶ�7ڃ�#�����^�ր�ߚ� KT8����L)c�̈́�ؖM�VU6�w��ǜB�ù�]Պ��ST�#Vq�F�XF;e� eV��'<�i�=Y�Wo\��lX��>�z���{w4�}Q_���`��ŵ8fs�^<�Z����Nx/�p��sf�PѻB�u6�}�R"6��~�Ͻ��߿}��U�*�	���<� z���/�e!�g6XD��K�5��G��W��]y��@M���gV�;�2���JyE�w�Λ���ogu_y�r��D�%����2�\��������cHk�`�XU\��h`��Tk�g:u��� �U-| �LM����z�c
�����z���aQ�.��򯱃��B�'��q�۱�!�6��05�F)��m>�C�U���$�C	�/���rk�wT�������m��Cbyt%�2k�����*xӵ_�H��Z�CWO���C�l��,9p��V�b\�R5�ڎǹC.U���`R����z_�}���'��C)H��[�<�ܠɬ"d�E��N�}��ŏ�a�0����ٳE�l���bA�����i��w���ڡク}B�2�at:1�/B6ǒ�Gn�q�M����{���(��ؽE��
d�A�3��o�1�zO Gl�<�1����W'�%N��	8�׋�?P5Z�LY~^$9�D��_J�$p.�,����;�P�йS/V/@��[t��~�_w���M}���5�/�+�f��P�e�p�tqDd�����7�rȖ�>���vz0����˩�:Ϯs	+�y�
�n��	f��mW:k�	v�!BV��:�@&�ˉ��v��^ab�c@��2��{�)������rz��\)֌as���ݹY�VuZRr���^}ﯟ{���߻���R-�x 2nNs�#��xM��ke"��oN6�='���#1̜��SBz�}Q�RcT5Eo�<)e缟��i�\�["����M�3�E���k�-�#J��sq��#V-��;���ͼ����3@����WhY��6~��Y|�^�*m][���O���٥�u����r泫!�C�{X���P%ޕ@^���
za	B�8�W3�3r��9��4V��"-�.T��An�R&�uis� �Y���lݟ��} �O�ߑ∮�BA,�nd���i��ϭ,��k{��=�tН�r���Nᮡ��C��p}����c���Z���߼'wS��c�_��ON6����zy0�ݳʼ�͡ZU?Ә�>���k��Ib�>{���
ݭ��+,�lAn��b�vhL��B��3`�������e��(�@�n�
����O�W�[���>y�!t��@GLu�	~@��M�L��4�a#���ۋ㚕�>�T-����v:��s�I�p��[_C����?h~;�Gء��сE��� ,����U�M5at�OEu3��"c�+�=-��<��y���x}8�J�K�-��E���z;u�__!�S��ma� �~'�$QD����ʱ��.]�^v�3����WU�S�t�7�k}�)�_�ce�=Ӵ<��k-C���A��;:un�˿�@���V�
������~�uenM֭i�|����0�)����8�h�(��w�^������5���/k�H���$T�Hq�)��Ƨ����ZS^(W�9,�"w�Lheq�����g��7ޡ���w�����r^;Q��a����l�B^Xȋ��Ĕ��=f@z�45�y�~^$��\�s����ס���$�D^���*��U�2i��#��9��1����	�.�M��MY1[u]�ɸU�v�t!ٽ��!��x'�4XVz��|O�����r���>��iȡ����&2�c#-:�Ϗ�"=���J�.#��v�w�y_���3�*0��JZP��~9�8��a�_�C���@�9��O����%;��Rb��
oh�o���9{�M����d�cl=n��Z��p�9]C	�dg��2�����ߎ{:���፫��bZ1Mr#�z�C��#8���Z���_�US�EUvWL Aw���.�|�Ofm��Z{�V�KT���"�x���m��,^�D��S�픬ػ�Y?���X鿎�(����ϯ�O:�Ӹo%r��gL
��z��N�x/dBq�-��	tE��}jR�zu�y�����c����D�s����Gr���cB�4��;x �b�.e4-��*,�.�ͱ�;_(F�H�h�#� ��:������U��ra�P��	%^����r�_%fZ��Y��y�GM`&�[2�\�k�;��/vZ�Yg�����b����}�vE[j���c(�z�8�9Dn'S�}�����۔t�mv`so��8p;4\+���fS�(��#�Ö�Muܕh�+9Z�W}�,ި3�'�mUZ��\#�����ˏjX�����fEtf�ġ�s/�T����U^�wx����8eGн�C����*dQR�TSr��^��{U/Ki��<�vk���͙�tV�,Z�YCy_4g^7e#{
�f[�t�Q�+��Astga����[���j��g;�W
[+D�L'�^�r��-�֛� <[��G.�t�8��/�\^T�c��J�x�љ�:�n���{����Z�^RTW��R��#S�'F&Wk����O'Dv�W��Io��w�ĥ�W�k8�!Ù��f�t�A\���:�.i��s2�oi��)�v��37�;ۃ�@�H>냁�ɠ�udh�\�@�Y�t1w�s��6n��gF I���$9qS�{T�\�oZ#[Ju-29ힳV,�c�E� �������:W1�>��o{�q=�y��lx��e.�:�ÎkMmD�u���e�1�h%x���d���1�۸�R^!�
��F���w�z��aݽq� ��IqgE��{Wt�۱��+�n�������ՠ`d_7����y=�<G�!J�~WQhQ�=����k2,�^oU�ֈ�ب��N�t���M�s	Cg7A$=��U��۠�E�&ŞnD�?��GU���wZ�]Xǚ�T�Ӷ��u�n|�Q�[co$j]��@M�X���,�v������GG`�Ǧ�w]���*�0��F���=Eq8h��gC�g�4�u_r�Pr;�M]�܆�2�Ĵ�׼�{͘��vn��:ȣ3�A*�c4�*�%w#�U�lP]�!�����Z�R�f$�Ǖ�a�8F���[Xd[C����v��u3��L�#����tt�2�`W��:�΅Ö�����aM�X��"M�`��]p�͕�Y묽�$xp��L�}f�J�,<���ʍ���Fm��eT������߈8ZB�ljհ��ݭ�}�*�Hr	�d��˫5�`(�u�F��UeM���������N�#9��uFVSkftn�p&�����|�\R�V6�y����da��ڜ�Ј�pO�������m����D�5�u4����E���|-�!���N
�����;:
Ü½���EǶu�
���9jk��$ntGg]u�qSS1�f�̗�<'6oL<��zh�x�9�W<[]��5y�1J�����˴�$}�Rq{VR�C��q㩽�l�_h35�-v�wWT��1�|$�c�p3WN��)�̚s{�8%*�V0�@[NK��i�F�@��iSiGr$Hm����5! ��`�EU��P���. �I�$\���P%_aj08iUFɵ��c�ۻ�y�W�%-P\6���E^s\4^��9�����}>�O�������g����ٴj��5U]܍�QS^cD�AT5LU��珧����}>������?�����~��j(�9h�"���v0E��y���J*a���s������}>�O����?�����_�$��W톊�*���Es.$�i9r�$�#DU1^oW�(�*�b��V˽Z.Z�i�$A�>��<��,ch�_�Џ,�U4{�*��&��LDC�KM%kT2[gl�P�i��#<���U%�D�^lQG6)�0�<ڊ).`�Eh41E��b֢Y�-�U��h������І��MAW��QZ����r��Z��E�j��*�t�*��b69b 4��8utj�+:;/{6��&���1��P���|�	��%,��t֎77iD԰/�q��;�+�p�Һ�F������uSxh�dS$����C�0������9���o~� �A#��Dޯ�$h�f}j��1�����1Xi3)��*��{�ئ���c�{&�	����E�L�+o绘
��Pw��]�32ס���U���dA�;�t��/n���>鼰�gPk�X٨.�n�۾<k[i�C����5g��!���bSv{k&��ь�ae�N�+�l�i烹����z�8�O�S�[����>�R��Ze4x��'֩�mr&_�O����e�����z�"��Ө�|`G7�n>���-C��lN����-i��eV�Q���CT�y��zR�r��6�KHvy����sr�P�|4φUxxl�l���m�\�2���幦�~	�µ�_��~_�E�t�b��]��
�W���k;�\Fwt�
j2���m�t.���}!�=�@xB幰����`�5�_�� L��r�;W�(u����ik,FO�7�����K�͎�ٲ m���94�^���q@�+���`��Z�+��`�b�D-z�]#u�W��m�,�5����̈���e�,����K0���1�zL�,��E�%R��ob�#j�n����u�V�CX��P�+wΙq��݈`\�7·Uw�j���In����OrlS�aQR�,>�S+��Ǹ0Gt��y|oNuZd��+aЧt���c�}{|�}��߾�[��?��2��<���Hӫ�d�u�>�ǯ�m�x��r�x�pO~��
��*��i�(r����LN>"KӞݡZ��R�b����3'������f)�w��KG "���Nŗf�e=�嵯��Fnd��C����N�q�����ǥ��G�o���FS6�Qaغ�V�6z!��v��Ѻj �D�{�B��^��Mu05<���[�� ŧ�,��T���.� ?��78��o���?v�������罴[Q�^1�qIƶR���gV��f\�3�y%t�`�P�NKξ��)��)Vk�b�v�W˃�jb���F����3W>.�-#%�Uh]��1��8x��V�t��qFzV�S�Lx�U��kP+'%ο�50�*|���w�d��!Vni�[�5��k�x�fB��;L;�{���)>n<�S!��p*=��	n��tn�|�y6�qJ���/�?�}�ߠ�z��8�<�E�ƶ�n�z�F�����T�P�u�����T3�}]1��~�S��P%�WF��T,�����kh��W�Ʌ��7!�ѷc�L�W��/k�w^c��=�E��n�����5|�4u5��Z�ѿ_��G�|v���[�/W��)�n��vЗ��3�ƭ��Ղ�mQ|V}s)9����{+zPe�_-ۇ��O�}�v;��m� aBK�:�]����Γ�k�f����_����'V�a�{�~�N����x��c9Qa�t�+9�ov�_:���#>�*y�;���;c�3��S��e�kJt7k����d�!Ux��,�B�2�uiq�㦆5Y��;����7�x]�D_�A�/�4g}J!;�=\���ɚ��i�&��`g�Q�##i��
�I����4x��pƄ=���3i�<�~(�z��xS{��1���O'�f�N�8�X���QX��gL��]��(�m�5�p�aa�%Rw�`�hO@�[�nc#�gu.�W�5���ߖ
6pw�@����Ȼ�O��,���Z5L�k��ՓkEasZ��}p�At�zk�m1 ���A{�!�֙�;�k�l���P�y���L��+qi���]�殕��T�l�3p��*X������1Z�ט��*0����zk>���������v '!�=�M�T�M����6*���M˷Pg���9O�bZ�Y�L6dt<"�����u��Ϡl�D�c_����1I���	���qo��h݌o�Y_�2�T+W������w����g��f��=s.G����D�����)� �&�sn�K�y�x��z����;t8�;22e���k�vf��vlX5�jG�:s+71Ůtkxq�.�kYǎ�YW�gr��6O_9ߜ�ϗ�цa�?�+��>��78�|!�yf�$�1j�a=B��@)���(��X�~��9Tt���e�8ĭG�/�V;��:�ig���Lqz��h��1A�d�tɧ�b�s�Q�u���wH8�nw��!�hb��ݾ���p?1�O����ܨX_�a�r��yқ�{�K"�CXVìT%�M�_�˵mh�M�<��qBsC>ϣ��㯵���i4��2c��� ��I����\�%sPKK�cv�\"����K%���	[����8�h�cuy���y�&ᓡ���)�h<��-i[p^����
��I8[����A/�h��NK4;�h�1������ר��Yܗ~����x�%�z^X�d�{	R/�Oe� �S�C��W�z_�t-�B�p�!̃џ�� ��r��L{�#��w>�jT�^+���_/]+�wOk W2Q������v�m.����������aY�/��Xikv�@�s�iS��2;�])��g�~BY��:����i��������@��=��+�S�68������y~�P�^
|��ek������wnz���K����zr�8�_Ȃ�7Ϧ�PlNѧ�pW�b�wK�Y��g�V�1��h�	忂f���J@�h�5w��V���9��<Ĺ�qғ�	���1��(��\��N)M��n�`��Wr
N�z���A��I��M�L�w�O���ȼ�=�翿�~������Ѫ��}�[h�6�S���T�d�ر��)�L�6����~b��~ƛ�p��jt��ʹ��Vz�����a� Ƽ|`��� 5���E���Hv�O��[k#(�Ľ��cl�S>�]�,%�"f8�f=��Jj�2m{����y"q\�<�ӽ�a4V�Sܧv��"��cŔ�CU���>����Q�=��2�4����J׷/xuCx��2���r��6��6�"p��;�H�`'��e?���.:�s	�⨱�&��%�bgD�^�՛��.� ��3y����e�:��s掊�u耙kױ����["oT�{�mi�c*ѹi>��95�����z��jg�`ޫn��q�Qmr��j�g�U^��	���M�������Ļ`�a�
G��FZ3!�$��1��9x���Tsu%+�Ĩ��
��-��Z#��J��ni�wR�����zj���N"kC�;)����4"�U���G2��_�*:x�K���6���?�Ǭ߷v���2��6�tl�_��
���C�'�.�kiܖc�ƙ<6����8F�y�����S��	r����rhѰ\ʭD�z�}�\�{�I���s������b��D�RFゃc�N�#ýx�o�d8T�Sy������ϜvNA�Y���f^�5�-��JV�΄��#jF��0��֞�p�����Cڟ��1�K�_�5��l��7�Z�)��NO��1��K����������0�l������(@'�~l/@c�y;#=.ޡ�잵U2o�jr̲1�6����C��F��k��Ġ��g��s�_E��@?-׬|d��ۮ�3���p�M�2���G�/��Z��'��g����]�����@v~���X|x<
9����Xՙ�r����B.�[�k2�#VHڞ�!6o4E'�����M��U<����w�V_�������s��������.��xrt�.��(��5���sȲ��D^���-�T���q��<�x�,b�v���"S��:#}�� 3q��9Bf���1U�ν���0�3�]S��9O�~Ԅ��+m��cs��"iB����M�C��.��^?-O��O?\��ܥ��<�lkEeSm��*��NC�O��j��������Hw�qU�4Z�TK	��&&ĕZ�5ku���k���Q}K�Se7���	W44�ò45��&�`_V}�ʵ"h���w�j_��-r�h|�f����7���w�3���%����
Oْe����a�KSY�{;/O2�ɔ/f�7�!{%���[���勲�IX��6I+�K2�l�l=u�evtO��D��BV��uq{#T��|���oo����]c,����oGs��ik�黈�B�݊��7�쪇�ǥ�.�ìo]ꎩ�h\�Ϗh�Kj�~�/���f���{-��[�R}Ҥku#t6����g�c�<lU��~WT�_0A�0�Z!c��=��"]4}r�7�F��� ����7���6�)��J��n��\��)�z7�fY���s�_�z�	���2��'�v9����y�!�u�X��Z�_���vl��c�����ǩ����a����}���t��Pj��g��T���p#�-BO��))-�l��q�`'�!��:��|F3Hm����TŬS�F'�/,��3ϗL��JX��vD��gOH�v���c��Zgy�~���(����
�H��LѺ�A� �lhX�q����ok8f�y�jz����(�o�����P�����7-v��Á���E5R�dG� ���(wP�А��3Ys@dy�6ct��y&>I�K?y��/E���m{]�ICE9hw�g�{@kZ�`����p8��C�[���7:�A�!������$*{�9!$��O�F�I^�Q:�,���Lf���?�w{^�XJ>�0ھ��T���~�q���z"�cXQ|~	-i��D��?a�,�)g�sד�ZYǲ�ܜi����̴+A�[�!��|3�3�8��`ӹ2k�1T:�o-.�S��x���gEP'�V���8��>$|~<�����q<���e 3��k�7.dty�D�����d>�'�z��N�}8��yۮ!s� o�[� �,α�#�˦��}�nf��|sQ����B��*</��OW�\��{��Wd�:��`���^택�|����zS:U����ZE��Pu&β��w��ᵍ���k�lڼZ�2��cQ1���lxMT����߰�'�Z�(>�%7�.�ŕ/CrT�x	nͩ���'\�s2��9�ȸ�p7��mN����#ze'ԣ�x��ݯ^�fP�ٰ�q�!��������
1[��
?��>>r�)*�����s�T�0��\��2`�w����eۯ�#�/S����>G0�{w�^oM<2�����<){��xfA��)�d7-�n+���j��5�m.�jy�x�g���'��������(��@�����_��ŻɃ�b6��\��_�i��(g�g)ĎV�X`��by�%k�6�6��8߱禪7�k?�Y��Al��z������9�TG)��Q�vUc[��.�"���C?y��#���i���]>���4�T���\��7k^���4��jsFu:�N/d9��z���lv��A��M���<9�}zڵ/hV����nR�"6b���1�B���L�2� )@���Ǜ�ܢk�Qbxc×C8�:NCEj�;��[{D��R�֬=��3$7kn���r�=��$7�%$��!b6di��rD1>���#�Ǯ���������M/�W�K�����=/��4#g�ӫU&:.8�|O�y
H�󸧛ϭ�T��0�V����Z`ܹ�4=�A�����d�
1��Iaݞ�Z�q�m�̼��ۦL%��n:}8Bf�"��C����;a�Y�G�v�}��3{llN���3�UA�ٸýɺ�	���ߘȖ�����;������!�cN�S��+�����vצg�;�z����D�3f�v,�ܣu�C�;��2Y�5���gO=0���@3߃�yaO>��l��i��DH��\��hSY��r���s(z�����6Q���S��*XX��l4��_"�
Vۋ��Yz.;^��橨����f�Y�k�d&�n�cߵc"q\�=M7��c7Z�?n�~�� ��� 8���r�CLk�X��Z���L�E�/B�K-�Ugyz<z�Z։o5�6�٩�5h}gM!g�{#j�>��%v��Q���K�6��!5
[ �;�w�
�l؅2�Qۜ��:��'����s�
{��V�)�w07#0����lӕ�I�w���&��g1[����n��)�<Ľ��k������K���Dz$bXU7{oU�6�d��D���e��ðk�����\�@�ǈ`��ۓ��^痻���S �QV�·�_<Si��=��LJ΋�9B��ř}�v�}��ᴚ���m����y�y�0�|�/���Wky��K�V1:�t�Sr��wNE��P5@�kߗ��_��fߌ�0�(Ey>u���s��k?�)�ѲXOs��Se�ˈ��ҝ�^�<�)\��=���h�Ҹ>���f�Ƭ�[$K����&�S<7@�<ޟ_ o�l�Tq��s.�bF�ÈI��?3��uP�=�H�E<څ��ԇU�6}/���}� ���KM����pJ9����)�k��[�tŋw#�:���<��VĴ���K�\gI���l��:е比��r��7{�\�u�a\`��`���1�>�0��s^Ƥ��)^��;�k��x�Rt��ʊ򯛰��W�������3�ީh~j����`Ѳ:�.���(3HP����ޔ��9���de��v����kq����qַߕw�������u
�j���L�������}\#,�N��t�fb��K��<��fT0ofi�1�k��y��N
�����4K�Z�E8R����u��N��ᢽg�A�Tc#c'�^ٚ�zMS0��ַ�˰�k�X��N�)�ٕ����˯�(ui{�"����4Ů�����`������l�+�,틏B��{6�iǷ��)+e���,L5��/��6�]ظ���p/WP㍴���j6M�8������r��Jo���a���mu%�un�\�뢵�{-P�r��kr&ر�;l>�}gu�;����ڔZ6�Z�׵"�4~������yQ�{�C�l&��c�E�3T��U���j�[�%�)26��zݴ���4�A���i:T5k��垃w~ئ�٢B����X#�k�p�����ە�u%4�{	x&ŭ�bfۃl���ӭmW]�ڄk-���!ʯa�n��O9+Twm�Īn;��@gus���_La�`����A�:�+��*�ZJ¸h�8���Sn�}�IU���ϩb�����r���ٙٵ�!'���2�1P3�m@�p�������&�"��(��o,JH$��>r�i���c���]��m���q�[�;�4��c-��g"����Ǵ�[ѝ�L�	��m�����\E�{�z�j��t�k:j�o\5�l-�)4
g�]���v:��:�-�B٫�K��z�F�GR+�g@��є_M��&�"C+�'���lE�`����㽌e_O�f��OmL����Ҽ���>�-��.ko]�q�R<ʰ���Z+:}���N�9K����8勘�9Yۙ�?lЕתg�W�E?R}ز�ݐ���'����3{��HaV�Y�JJ>(�(��s��M;r:I�W��c�A�V��kJ�j�0'�+ϲ��ugN����2Y9ҸU�} ��v�.Ja.��n��/)���d$�O�a�6�X�d�cNGvN��[�ͪ"1Z���o[������ݰ��tA�ѫ#���^k�;&B��Ppcm�蕺5�CL��w�;���/c&�����1��[��/z����jqE�a����;���+^G)���C��]Y�k��8;��ׅ�cy���*��Y�����b�%�g9�Y,��R�L��+3�����&� ���8��i*�Y��,k�w_5���'V���>=�`��[yKJB�&ۺ/6m��0�Q,��x�,����������P�;[�.i"�P���bD3i<�+E���OFJ-V��Ѯ,�spv���a�U�6X��������z��<�#��q��pjVnu�kݹzz�k~R� FTF�	Ք�OE��]��Wj����ıo)����v}$g�r���c��c�tu�\��
ʛ�r��#�����听���5O\��y�n.�::-��f[W�]��T�GV��P����	,�Q�LCTSE5Dr1�(�Pѥ���H����o_������}�ޏ��3���$��3Gy�M15MUQ_�4�Qj��b�)�h�i1D�?�c�>>�o�����~>�o���f?���*R�1h�p�Ť5E1Fb��Z�A�yV�Pߟ�O�����}>�����3?z�vI��h4`�G�ѮE�6tl' .g��Zim�LG6К�(i��h�����h�3UP�I1MG6��&������i�N�9�KDl96uT�&�CQ>mQc6����-A娊��`����T-�MEDL�#U5D�QA�MQ)�RP^ly��-s:��EPZ4�\�i)#�5r��V�G���� ��TR1��t-3RО�!|�Eؔ�psi�\�7.������w�/5�	������:Z�ٻOzk������> 
������_/oJ�!������	O�T��Жl�h109Jf5cy���v�N���ۧ�����X��L�s����`omT�{�-W04��W2��P��#��؝$w"��k��u����3�r�m�r��YR�0���|�y��UD��\�.+S<�:*����&ֶ�7T?_!��� z ������<-��[c��5�:5���p캃G��b�ۤ��gmvg3n�f%�!G�}����<��6��nW��O0�j��3��^�xd�db�{B�c]�kjဍ�8����v�=�>Fe��� =��7#��b�W��h�P�Z�7��-I�ߊz�:��z�Ϩ���G
��g��Ȇ�t��р0�����ƆM�ɗi�*��z1�-1�n��2�fst�ok�֤.�Sd����|�H�?�?~�>�c�kѽQ��c}AۋIK���ʘ\��ȩ,���Ɖl��q�C�hu�?�yP ���+�ī�}��\j����ݰ��5�;;�q��4c�͟_�6�/�C;���˳F�\u��\��Ľ�0�z���:H����x	�;�V%��DU��"�J8��V[W���o �̐.�K��[�y�A�Z.�T��A�ȭ���.��yDe���L����w;N�ܕ۠
�^��.��dh��q��|<���֮�W)�HO��z.�JC��N2��j��@�U�>�;/���(|>+K $N{�������uU)�y	�?;�|�۬FqV�I�o��w?Z�;ψ����Ez�\���O.��0�;}�܃<>������,-l�a�_�矕A~k�[&Ϡ��}6���������,q�險
e٤�Ed�d�)�}�b]���kC�'�O�?;=���DT�c-�!���UR-vu�&�ճ[�+�f��gw�����w�N�5=�o�����S]8<��s�<�ɶ���#T�#	fI�'��v��Ky�H0!�VM��0�7$��5�*E;٨�{8��(���,����k������3cm��R�]6$��e��i�S8�s�+�O�����b�i�S�`����odJ�Q�v����g[�|t�z#�'�r��J��4E�[�����*Y�8��;�����������U� `&����C�:�;������GX�z����x��s��^elvJ�.�o�⚞�_���P�0�d���yz�<�]�����h~K����Sjeݬ����qyE�[ݝ��An��t�!�N��ױ,�I�}aM��^k���:��3Ӯ�^-��]�  @hG,oq��VN��bG�׮����6�p�D	�il/*��ٸ��^j[��v��Ό�ͮ�3�B]a��$x(	4 ,UH������������p��v��eYX���lo-l�Z9�(��O�>Ê��i#!�欿����N.�,?���� �X�FC�]���	�r:��	�-��:z��>�<�@�X�
9��6+�W7���L��rP�5�d�9ׇ�Y�ǙN��f8��8ڮ`��� c�x�ϐ���:k���" I���'|Ԫ��hl��CF��"
|�M0��
�^����ljz�Q������9�-l��������-A%�R�D��?g3�h,���x{��������9��b*�����c�p�d*��P���2{�����^/~Ϛ`��'>:O��+:���W�.i�L(�l~N3�_��vw5�V�����zt�Nl�L2�����a>��iP^��G�c
�h���l�P�emtk�s�<bṂ�̋okZq�3@�TZ�b��;>9ȏdFDH��u�9&[�k��Kb�\78vd�阽��O���*�KMZc=���0k�����Tm@g!��E�8���? *�^��幂G@Bj0�d��M#]1���6l��eys�K�<WP�oj]������K� ����E�G{��!jӲ���x��
k�^��k��v�f��w+)DM�m��s�U�.zjlz��h�	U:�3�sj�c���[�m�'M:y�{���s�ΓnC�G2��&঻'\9X}b7����> ���uV��.R�{	۾��ϙ�.L�����C�{�8�M��Ь{Ս#FJ�+Q���s�5K�Q�Ӿ3������5q-R`r��4(SM���υ�Y�9˸� �g5��^�ƫ)[z�]yb�f��E��w��.&�.�h��_��~�G��,
ǧ��I�uU��lڵͶ���%���M��U8�|T_L
��:�f��_z &���6N"_)��l��k�ѹ��a���fЋ�<Z�*��ؓyU�w��yY��?1��ݖ?~/�(���|jޅ��Y�[���`���2��{���1I�~h��'s����:�s3ϟ���u�������t��Hw�/B؍t�&�ȷ�������J�N����7^�Qm̯G?K��=gD�=�W��W;���Ӆ���h�L�����l�ԉi����
$��~��NZڢ�:�h���M�I4�<��ؙƆ�;"aG�X��t��ymi�gM6'M|������c��2g���?O��p�����D;Zށk�¿~Cǀ�ٯ,ۣX�}��%5��z���nP�[�f�����ڲ\���v�,Iu&�\�^�4�L�k�WD)�W����^z�|��Q�|�Qz6*� �b��2E�=Y)h��V�`p`�9��N���=r���j��	)�l}�d�W^�� ���5ɪ��	�r�W�y�0R5s�I���>�s��0`W��k'U|�uC#��q0�9�~^�!��6�d<���JQ#�x�ߌ#����^�T���ƭ���ǤmA�-F"�CwvÞx�;�3mo��p�t�����K���}���Nz�df� ��g�cSe�0�El�9w��{��������6%	��^�w��ֻ��5e�00���e�cc�(��ԛ�+�e;���Κ�̇x�n6
�t���K�A꠭�0;}�P�����>�3��_K��Y�@���vp#O�K�N׾�����vۃ�%~U�V_2=�� m<�FP�w�.���U��6�f��d���Z�t�!�vMzVU1*�4��z�5��p%f�;p�	X?=�}�Od�q��٧mЦ��5V���{�Id_4�'7�"�h��{��aċ�v]@4{�18�TS��c��WdYΨ����->��N'��D��x���t�Z�����B��z��4+��WdJQ��Q�;vv�3,[/q�?x��c��0��W���bS�@>��b�zO�eP�`6�8ݪ����S�1b�󡲡�Ieod�p֊r�S���;F�{���t�{�a8#��w��f��u�z�����u���}�(w�
���Y3v^[�s{{	���e�S��+��YV&sS��b]�ٚ�z�_��Gď��B��z�o"���P�������0�G�;��	]pޗ!�
~d�D˴�_)�R���1��d�k��W��2ר�%0�x���kߢD�0�.��GT�.s�t�vȒ���� q[뮉�`�j����1>�m�`WC�J�[�# W���_~���X�Ƨ���?�9o�!���c�O{�aC���'y��0�"dUxY5�6���ʾ�l��8�=����B4�6���t�����'�g[N��7�OS�/K�z+�ȹ�B��qdǵ����U�w���Y�Ar��?��_���+�r����l���P��������1��Q���􍮒���<�;x�g\YNH8�>?32��^|\CDd[{��9e"�ۧ3+�A�m�9�˕Ŵ4���D���7���W8��-�{9�U={@��y��;"ć�g�+�}U�x�񅴮�EN�^�m�z����ͮm�ٗ��<f��ty�@�y�k0.2
xi��8���T�������:�K�WF���0�I0e.���or�q ����?~0_OWb����2��v�M~�T�v$�͖�����<rT��A�t�sg��u�dGL7%y�d���hp�a˧>���+�)�rԊ�6n��w<��oJ�T�����6���%>|	������8��z�j��V�Ԝ �b��(�y��F�!�>}���_���Ϟ�U;zޗ�y��<v6�1�c/�a6�R&�ukxSW�\�<��\⪇�����+S�#}e��ε�>x2*��S�㵝4�wk�L��%>�[�6�*�qsl�e����̻��W�/˨6��vwx�H{h���|��y��1m�3,�zdǔ���*����g�t�TS�ĳ�rw=��Äo(P$�ڝ{��%�=�xҫ��-��b�����j�_���!U��I��ʵ��(�<����M#�6ęf'�y��?7��'5`<�R��w�q�ԙ�dXSy��N�O�#v7��GT�%��Jn<�� +p�������q�%�7wl
�5�wm�vvR���k��K͞�6c������F��2��!dJ!a��1���a/=K2���ni�.=��N�n��_��{bɡU�S��ل��w8�	I`��5����Գs[j��OV���� ��ܛ[�K��������*d�E���dsas#�[.����x��4�2E3���ɟÚÕ!Cψ~���7�_� ����G~C/�v�e�њ��f�����*2z������v	��OoVM;��,�*�oX�Ӳ"5�T��8���r�"U���칡<��2'8ܷ9�����I�;�J�L����\\_<���
$��l<ӇXSj�ĭ�=�S59�Љ-�����F�X�̛��~0�0�	��;r���m(��N+S�,{�Dz��s�4uߘ��<��L�XD������Pl�Iq��H~�˙
F7X���4�ױ��9������L�����L"|�z��~��9�u�i͋���\��v�sR��'i�70��}k��@�0JSlx�4+\�*+���X_��r�%)��{��v���v�k����N>���P��Z��
�����u6ʆ�s3r$t�K?gsy&�G����~L�2���T�=�%4�	����V;՝1��gM%�؉���L��71#�����|�fڡ�%�A��1��s@P����z�~D�����m�g᛽�\��Ĝ٫ W���Y:���X��XT�зf��v˽1�<4k��@M`-�yhn�[�"��OM��s9׊Xq���C�S"�^Z�+�`S��
�uQ����]D�]&���ފ|~	?q���ea�����c��
�M݅U�U���&r�\XK�d���e�M���M�����20�̆a4�8��:^��M��Mͼ��}hJ4x�V��)��d���T���<�=�ǏB�}�����n76��`p�+ou�U����.�gM֗b4��9Ӆ�:������IK�S5�p	����jA���\����4ܸ�,X�;]�+�tIMv��]N��<�a���^�%�ܠ����_Z�a�흉�x,��ޠpȉ�*�=�̸���.A�v`��V�L��Z�s�B��ε~aq�z�S-�.U
j��5s��)9��o�U���oy���Ӵ��ږ���ALm2�$;>�σpv���⚿�E���2�o��@r�w�j"�7B������H(,�*���>�i$�������
?ߓ<sʼs���V-�)���Q��Y�48fw��A��y�>�>{J���\j�2�����#{�y����1��d�mڭm���^��R0�Ѯ-��lG'�q�^�4^�E��<��Q�(��;Au{����?߁�a��+��~C����G$6��Ŝk^�KH� �X�_[�'[O6��5^w5�{t˿4�z����f�<|U*=���z����{Ƈ'A����U�Jaoijy;	e��
{�ˍq'hLMQ[U���_L��l�g�绡��;���y�;[��S���^�\��\DH�{.��?���e�Vdے�{����C! �M�pg=H�C_<DF��w�h?��$��O8(n<�޵Y,�`�lnT�q[zΜu��a=�b��
��#б�\U8И����429.Ns�����j�6ȁ�{b62�����S㝙��&�*���֠�n�7�1���|<�0� y���?j	'�>�`����`ɨZ�o�l$Ɇݷ`W"g��[L���q+6~��(�����++�V�|uX◌h��\�q��Йs߳�گÁMRR�������E�?�7�^_��;����?z�k4�˳O��] \��B�CR|a`a���*��$e2[��U�5���|S��׌�=˯r���*'�C'ڸ�hӲ�Y��#^��n��V �Kw��F3����,�.ة���Os�a���.���Zg񂻢3���:��#D�L3v�ӛ�of�v9L`x��������5� ��̲d�.z�P�c'����2�;O���Ջ����i�)�\�nK����<׸V�Km�w��:1��]S��#b��Z�r���~�B��eO�V���П�sg��8�ҋ�Ў-���}����P����9�"�9h�|j�ҟV[<~82�18���1���kZx�4j+^B�2�sI>o &kq�w#/3�;�5�|�v�Α"�~�GqP�w�;���y�|����N����I�N�^G�x�謱��'h�7S���h��n;��6\B��Rh��"ku��V1ugvX�푨�,��G0�
R�ݧ/7��\�PB��);a�W�q��̭�Pr{��i�hg^���=7�E��E��!X��꾝8��c2��"��h˝oK��h���/Nt�P��࢒�6^�KF3�f��2�1�n��&�Y|����70���7���PX\-�,�ܼ]ʕů�X��I܀��Բ�Bҽ�c(�q�Ұ{�������Q�˫;-j�nm�c��1;�h ���P�J
p�U�b�b�z��WI� �ޭʈ�GO�c �t�KkENw"a�lөE�x$��k:�s��QV��̋à��z�"�|H f�g���5:�l���1*�W�)���ௗ�����o�g�wZ�#y��wA�95��`��s�.�г�}`�U�o����#`�LC/�F���L�ĎW�� ��8��NKS����T�%�*}���Ԙ��)9:'W���d⧋���{r�r�9.Y[n�U�ON��鼸�sN�~��:s(Վ�ֱ��k��y\e_:_#���ڼ}v�pK�b7���&���.5�]ogVX��:�Z��e$�[��fʷ�]q�N��ļ���f>u��}t}����u�'����Dm��۝ϩD0hN�;��+�D�A6E]���"˻���t�+>*X�$/*ƙ*�HHR lK�E��T-���G�i��zNU�E}���3�L�2:���+x�����VՒ`H�~���)�j�#�rw�������|�p;h�J�X���w}�o`�q^F�l@X���2q�w�k�y8'� �,[�ޕ���L�W�����ˣanr�(�YC��$��v�>zբ���zΓ�1�0����{�s��7}�-n��nF~Ṇ��Z^^�=u��8 ���t�$����f�=\�p�'w&B,��:;p̓�e^�֣�պf�c�S����c�u]�x��c-��c&���樓3�	^}� 2C����$�;�۔�b���ݴ���s�Ͷ����T��ѕ�lp^�#�)�:���us8��v�ӷ�"�;;��B]Պ	�R�!�ҡ���W�ۘ��]��x1�M�j�+k��3
�w�钳�K�CQ.�!�NNΦ
f�JJ�>���gU⽼�S���E���5`͇�kyɯ)�q����x2�"��ƫf97��;��'��b��fr�1��tY(mA�_n"f�Ż�Q��;a��ڙ��(���ڮ܍��:;@�Ù�U�sM�|��W����,}��xe݄��gJ:�,�q��|V��ˮ�ge�<�i}/)ڧ�.�F��n_eQ��TJE/�2�e0�TZ��E[��KVQ)�b2,��!�
M��`�G�UR*�Q
!�q�J�2��*�D��ے6(��$5��'���h���71�"��4A>Y�
&(Br9QQRm��Mh(��x��z�}>�O�����z�fz����4U~��SG���i-�U%�mPDUQ�������}>>>>>�����fx����\���i�s��6��<����ZCN���"�����^9�>>�ϧ�������?���~�O�B��y�5�S�TTM%4Z���gE!H��PT��=^A�ּ�RW+a���BUQAJ\���Ss.�A�K�6�>K��[�E��=G
���A� �'���%��EA��â-�UHD����.y�!���T��ZtRyG&�����A�8@r����4�4y��LVǗ#��RPi֒�Cט"i<���+���B�P���i���gli֊5M����LԞA���9>@m��_I��I|	���i���V^��`p�#���������q^ne=r�V�hʖ!W.��{��F��\�n."����/�tKJϔE$A)H������ |@��!l��x5y��I��a�ؐ?�5儜���:���,<��ɖ\3[u���{i�/d޶&��)���2���Ͱb]Pi��I�=��hO����Z�@��7�B����,��a�6�l��4�̙�H���[ͯ@��f���O�o:����:��"c �����!vaʦ����S�ہ�Ӎdnȋ�ap��YC��A� L�l��p�<������#ح��g| �F�?J�sS�Z��/��(ŷ��V�2���)��H�]6�[3�T���u��(�Ⱦ�Lv3��&}m������Ԝ����t����o>���nP��1��:��'Z����[�@��a7�캚-�j-����S�hJ��X���)��/9zq2g�:���jʳ~f�^*�{:,eG�WA��{��'���r�k��R�`�{�f��i�ɪ8q���׫��������H卹3�1�*]��m��=z_/�럷>��es�*auVnN�Ox���զ���M��9�Z��/���Z��DC��w`{Wk��b�S'f+���S"{B�v��ݴ�R��НZ�#)K��QgAA���$�#~��elq{3�y;2iޣm�vd�4�z�B��xF$�M����"���2�E�r�Ԃ:��K���k5�5*�|����e#YI�pC���|�]X�߃�y�y�����U&y'CT5~	�[��G>*D�1��R0䌖G]s
	鵧�]�`N�â�}-��37�Z�ߜ;�s����B�j�.(��'��w8Ġ�q)��tS]�w'��^¿Y�c���\D�D�`�[�_~�YH��oN"�e�=M�a�Az�Z���މ����}�[�R�Q���I�ϛT��_d����"�n�륩�6�Z�r�cjߪb�&�+�'�W����y�6�4pR:<�ά�K�YQ�[F���	#��6+��)>��3x�- 6/�DYW��|��6�U����;v����e��b����o.���@uXFS[q�\���MճM�yгe�D���^�
7:}j��N^�(r(U�[Nղ�"����I��x</������a�I?/�4�]�F�Z���et�v� ��Ƌ������T����w�������7}r�5?q��	�kJ�W��סs7�YyY�ֹWh=9ԑ�
a����'��Hl�j����CDᴲPî��̼��w؎U�n���x�9�:�=�v��5Λ����vc9G�m�-���Cc�պ��b�J}�a?mb�W%�R�s�ߟ�a�f��ҐC;4_�&7;���+)�
EW�MX��(��lj~݇�I���C�Yc�&�AY^ĩ+���,+'�4�*�v�5z�v����heT�>m���Y�ޏq!k�Ol���z�N�R���J�����k��;r�m:�~k��*�����]�!�"���e�e��ӽMұ`��I_!K;����]M��Fw�ަ��\(ۭMr��r��P%oM�/$�A6��:�nE��<[cD]��5M��۽�j�^#������}�z }�QT�a�6�[f-�"*z���܄e�"�e�+h�M��5����p�۽�Q\Q^��vO]�Qʣ�NB9߆��,�Ū{6�y�K��u��ݽ[8݊9gA���fU_���%sڌ��ڨ�f�C��.���1�.���!�~��ǅk����|#D�kԄe�:�S�Ŗ�j����5����ӌ�Y���E-�lh���T]3*3u�,D=�T�fWD�e̽��
��{A��Y��;���7����wf�Et_��=�P�K�Ձ����7�3�̗h�A��Gv�	��<�r�vI�\�g]�_l`�.S�M���/{w
g)�s�8��[K�ޥ��Ev�j�\���l r�,C:}��1ݙwM���ř��)�r�`��	3�+�=5ݎ{���O՞���쉗�~`{'tt�������ky�$rY>3�u"�2��Yr"ј�����'�=.��u{�Ѳ������b���G+w���py��إ���a��?��3�)t����"/2�I�>���'R����a�Ҍz���8E��/��(�EYn��]GN{�\��[f��}aVIT�s!C��������[Cy������Ew3��&}�̕�-޵YLvk��co\��sU����R��1�MR�p�\ ��~���-�6��+�a�Te+��x�ue��Y��{�*:�N�{�C�K{�$���7��VE\���9o9��;�\]��'�ؤ�{�HVo���܆C:X.�.������fW�|��=������f-�s"o>��K켡Zn��P�J�xԲ���5���=���=���3��Q5��.UŠc ˺z�9�wHsl�^����7�)]^��Ŝȡc�'Rʰ��8k��g�+���k2a������7jr��Ln8 %8�b	���2?����*�������I������ޑ]E%݄�rF��6yd��x)��{�߬6����y�{O��j��:+ݚ���u����a���cɕ<'{���ьx����kȓp��t;��wޖ�<��˫�_t��'yu��� ��b����SPj�	³������r;M0��x35�y=tV����F&�A��ᅆH�����@J2m�3�V"d��s�#*�Nҽ��m�'�j�䏰'��ft6�}p�^+3|�DU&�Ыwc��ג5��s;x�A'�L*�]n�?.���6a�>�?^KDfe�݇5�z�Fn�/Ml�����^u/>%L�}h�ߩ1�ߵv ��¨2,罚�Vƾ����\Yu6��Q1��U�a
t��MOW��˻s!38a�?:��y���d��{0r�|���=W�=��p�ެ���V^žj���9�Nxe��NBЋg�r�[���[��V�/{\#%'pT��p��+;V�w�n-Ƿ�e���=�$�h�4�"\l�c�k'S���)Wov�b��i-��a�1���rf��*�TV��v��*�1�|�y�Y��3?}�]Ve��P�c���fO^C��(���2�ue���/3;���d�\��<8�s��^�*�*C[���KdY%�(f�F2�ɖ��|��3K|�>���OB��J��#��/�\��0%N�S|�T؍����Y��]��a7���@�(	�x�
}��vyN��nH��CX���sv�êz2!q�����b�2�rD�~;��kK������7����\��RW��Fü�BQ�eLޭ���>KvE�>5��1i����vI����� i�����p�t����S����9������j���*�F�ד�Zc���9�����%���ń��^W�\��a��"�_u�gX���N�Y��ā��c�ks���@��d8Д�٬��4�ߛj��2��9 A�e�v�}�G{lg%�<��r��r��[o�x�����v;R��Y<��K+��Y�wn�1Q�EEX~�M���S������Dj�\�uo�Ί����w6o��7�m��T��u:N�z��n
���;��϶\�u
�=ON��vطq�+�n�z��{��?\��r4ʫ#�Ͻ���ݵ��s��w0����.�or�-�|���6�.�����KU�6n�|�L�/I�<��Z��ֽF���f7{���o.�r^�m3��_�Ⱥ����Ut$�\K�|�k����L�����N4b�}��5�|�w���G�k|�}A�o<���O�9pg���]���o��*0r���y�Ǉ0f�vc�
Ձ��:��ߵ_\���-V��M6m(]v���q�X�V�R�gNo�ժ+&� E�g�;;0X(i�7Cwy�x\v�Yg�#I0��;�1�g Ϊ��n��r�}9����~^��0���M�خP�ޯL�$e���=�OnhD�jONVvvUR3�&9<U���_����,`Xע�+����.V���35�$l��]d?x�+:�fݐ#���LB�sP���L��y�:�,�wBP�Ƶo�>�|χc��f��|m�3����Z�]�
���Rx�;6gfo�Z��ֻ���P[���[�^\��<�r��;J7��չn)�Q-T��w�:8��*Sڶ��:��kC�<���¸ڍ�_��Pԉ[�Ω��U��mk.'��	��a��+�v]ja�@��� m㞵1�v�����7wS/f&9U�9B�q�͌��y��7�a"��6IN����ͪ�x���*S�ȶT��e9A�{ٞ����iѬ���xO��@k������iNScdC�`oq����2�zZsw�]����&�ڈ��#7�k�?|����O�R
w-����+�3���8y|_��;�.��8�Y��%��?}�ol�xT(�3B�,��}���Z)�tF(���L�6}�`�ex��@�N�bg�&t�O7w��L�J��٤O[=����c8��L\��S�����o�5t����w3�C�^س��25uE�z�w�/fC ����Pps6��56�zM�)�����f˷Y�C9��Zޟs��vǒے�v*Ҫ�U<TU�:��C2�ۆ��#&IJ��sx}�:I�[��,��ރH�d���:�[���'�FM�2��pݗ5�K�I�l����W{��(�����������݁*\���v-7fP=k)f=8��פx�<�ޔ�r<�;/z�o����@0��"]�-���xCk�-�o��f<7��߅�����V�mpQ7�x�'�,����{:D�|���ٌ��PG,׉��;�-xU��2�#}Ub��D�f.�����N�GM�R�+̍�_к��wb��WC\%��#zE���D8���y��w){���#:{6�R]^�ӳ%�p\lK��k�pK�R��L�ݘwr�\���������$N���X����hh�ʹ���-T�Ң.�x6�@Eo����u��1֬��Pf]i�q;F��xwlf�T�5�^�>{��v����ʏ?nb[�ލ7V{_K����tj�1f�rGKύx��6�s?��p��
�g�i�p�Ÿ����Os���m'��C��z��έ��Cu�a�{ 2O�� %+�F6�=Ҿ�{z�l[�K��뗮��	z�G*���<C;�ʱ����'��v�U��"Ww�s��qM���6��n��l����:W�B���#��][��Om�}y�crD���,��vß* "�,��w�[�c��A���b��LszAuvB�\ra�x��\����uOs��O���%�m�����<��f�{�	J�z��?��-��� �a*�]O�3{T�<�B��u�ö�-i]��K�l��gֲ�b�-�����Or�]Nܥ�mI��|Orڳl�'"2g�y�&��jlD���l�r38(\+�NV��=3NP�ݰc��R��w�.�Q滆���5!]X�de�zE?aj�_^�pQ.wrɼ���䲚k\�m�v�܄E,!�8�O�Q��6�sG]�{��l���gc�Uo*��U��u���ڨ4����QsҸr����|:�WA���|���h{�����ݲWM#��bN>I���,T�7�U}6d<�s���j\ފS��g= Y-i)��ɇ�mno#j�s����E#8g^��vF��>�OԮovUd��#���g��jK�<S�����>N��w��|7J(�Y��������љ��7�����5_��R���]:��v$�83��{�i(95��F[��{���Wo��D^Kֈ��nSi�yV�zZ�%r"�M:� vᬳ�h.��V)��x2��!	\�R��L���we���S|�
�[���i����q�8�(N=]QAu�e��`il���R69�d���ۥ�p�5�m�VaW����$�^�t���v$+m�хو��k����瑻��%c=�G�}.gfr��ւP�r���.�+�8(�P�L��j�d�ةu�ƳIb�ި�.��k6]�Bm@�9��)�c�\Ĺ��X2vwHs#�і�e½Q��WN�����X�<pP�x��D(2ľN>o_5��1w+H�c�U���ۋ�I��N��B�-Lj�g'V�P̺��
{�q̑���{�ֹe�HI�ҹ��j�N$��|K�N���Y���Ϩ'v�(�	��b�\�cx��;'4�YҲ�u5O�=ߖ,�J�qz����nA� ����ZFAm���Vu�x�j�C�+��.�򺷕��Y�IK,fIq�X҆d�ͅ���y�Q-��l)k�|�͓qẘ�Jk��ԁՉg��j4�(�ɁoU�Z�cTJ�\[�s[P���Sv�bzl����R�_�(�Z�pZ���,.ۻ��,��Hd���/O:[r�f����-2݅�	æ��V�u5��tj�'�u�$��6~�B��gO_HWV���1|	q+?{��� ��T'����b�
��q��v;>o-<i\��6�an�ߗY�EhU�渺�]QIp^ܵ�=��7�C9x#t�0��kw�c�Н�B��@qv��hN���K?ȭ/1X_s�^Y���ui�RW^�Y�66�Y���к\}d�N+N��!�уw&ؔo�]�֔]w>!k�f���K���|�LW���M��S]��j�,���ͻ����+X��pW�8O0uÑ�e�Z���)X�;%hh�u6biJ�d��5(�ν�9�%�����!��ES�%m�Bt��G�wu/+ox;�efP��2���[NWl�\�0laكj����YGp� ��r�7��@yn�=:��Y����Ese�ľ���K���%�{�����h�]\Ch��u}Ǌ�^Д��XR'nLO�z�֬45�n3Ou2;��X�]u%R��C"t׽��vx�%[pGYD�5BJ��2�s}@�&��&;V}ǴdN'`�
9��GfuM�L�&���Q��f�5�L�+L�]b�r����y}c��t�fK�x�m�����ۉ��+����Xb��9fR���3�'d���uB�@��bˮ��������Ԯ�I�B�]�[�i[qf�s�Ŷ!ܱ��hLP�9j�g��U�B�jV�q��N30۹U���3'1�bh��!��T�a�'�'n'&�b�����rns��~����
�����:�!AE5C�h"tQ^9�>?_��������������L�u0_�l�`�xjNCF�5�������70P訂#A�9�o��������~?�������E�h�G9�;y�O �ꚭug:Jm����]�ǩ�#IG5�Cs:փ��<s����}>>>?�����f{�����N%
�+k�T-:JU<�7��ڂ&!���.F��E<���R5��6ֱI����\�P�F��mc�(Mlj���rdh��*���^�s�8�K[a�Ѩ�Fզڝ:_������6$Z]<�<�P�Zy�j�5����cj}�p�S���;����m���l��r�	th�L:Ѡ���LVˉ�h�V3V�X�حfM���1V�9ǋ�\��-��Y|�QyQ�s���[�nj�'��F咃�����sk�����Պu�A�l�9<�m�Ey�G����<�lh�4���`�'*�("�R�U�AEU���sBm� �F�\ư� Eb$}�c��m,qU����Ɩ�9,a��P>up��x-�0��M��X�\#
��QA^�g{���$0��/�{��߾���n���_�֭ᛛ7���Zr"�L����d׃J��MQB�sr��;DY׹6ӽ�7�A�P#��_�ņ��|u���k�3�f���(&�� �>~��Vw�=�0_L�[�ƿ:s8"rm�3aG]���ݘ�E�P���-�_���k�����}ʌ�^�ƻY�c�/&Y�H����_^�wU)�}ʈd��c�� k�}����X��/8�1��{<�j�{|uZ��|�N;Z<��|a�5�V)�Jbl�M��t��_}:�Ă�3�\S����#���4� nVzz%�3�y���'e4��{;=���9�=��Wj7:���\<�F^��K�S�-��	�U^����3t�+���qN3of��PZ'����Cl��LC,�H����ƛ�O�^ksjߔ���z�P��]�V��̞��CԶ�'����������o��oƞv����~�<=6�]�����c�2]�vc΍���ń[x�X�����ܒ��Q��p�6	����&�$c��2RN�	V�Ic[Ѓ\���c�k:D'B��t�1'T}�/:�<�gmŲ�2�m�`�����5�7�w2�#����e�Ϫ�g�%KU�[4�7f$^6�㲋��~5���PG+�kG#�Ȍ�K�����]��w��U���*�����u����ӷЬ�J2�6���������x�рdG�Neww�c��.f։�[�^��t��?�s����K�<wk�WI��@���-�m�u�ސ#C3'����h���z2ݜdh�ff�x)v->���2w6F�C\!� 70�]�t���֪=��Ly�*�+$u���@�ŗ�O�X�k0�Ϛ�}�5���nϚ�}{���>��+��?v�E:^����sV�U��/84C��sǝ��`Ż�Q�v�>��+7g-d6We6����نdT�]�\��ȴsE�tM�@t��d#>��,t�i��U/gw�PrC(p�V�\ͨ�|�OsL���AVѐ^���=��_<J+����n�U��������Fee�cj]�.��k�d�	�w-,k*g�>�#3y�8��ԗ[�r�����*�x�#�P~U�`��;�Xmcޭ��e2b�'c�%��D��zu��t4=2m١�Vd�i7s"���T��V�ǷU��Wj��j�����#����	C�0�$F�}��\7H�m$Uk��q!9ݓ��+�d�n�8Ӯ�6�k5 Eϊ�͍�}�SN���4C�md�X�Gٽ�d(>%%�*�s��@ջ�5���b��]�
ٛiRo.nM�9E�Uׄ�q�]8K*}V�em�r�+*��׫E*��߫�����oJ׋�����nOý��#:V��(�x��q�����H}�mB`���C��m�m�͘�W 9P+��W�7X&�ΫЗ��ڮ�;W�Lwg��M�t�K�u�]�+�xU�4_���ũ���� �7x���U�R�yf�U���:�H6?�-r4���OSk�L_7��+�"��Ҹߛ��|��
6Ŷ�&�ǺLZ���'��������;(^`O�՜��(۾ޫ��-�6:,i��i��ݑ4�ݝ��cփ�S*#�z��-7ݚ���z��y�Rb��õ3�g��t>��۬�tj�7��.>�x�c¦+nT̗��F%��vv�],Q��=��1)��u�j\�R�RA��jrRW39�̼��QNh]�N�g`����L���6݄��Ȍ޼bp��Qݹ��p�����AtO
>IP��hdϓ�®���DF6�sRz��/{ZO���.dw�@w�`��b�
��ŧ�٤�� ���G]��z>'M�:�ęcA�=��<�O>��pU`[�oi��k����ֺ<��v��iQǄd��G����z9�i��Z�|�ѷ���x���Q7��"j�j�DY�sO�$lgK(�_8OO>��-�6����\5�>��u�T�����z�uȍ���yu��~1x�2�W��ˆ`���k�u����S�13�����Wp*�o��ʛ	<ץ9xV���~ݤ���M3�]�jQU���H��e�����֎��G���k��J{�-͠���7l�׌�C]�[q��o����#�z�f�b�)��A~�1�e�K�iq���J�y]Ľ[�f?�l�LM!�y���*��ب�5ܞ��[��J���=��NIm^:�5�o���:��r�|�쵛N�#U����Z96p�����c�U꠷��咇Ƶ���R��Ә{���]��Kf�̸�5ViP�|jIFq��%�]�YѠM~��˹~�3\�b��}���2� ¶|��ǥn�+��͡�'�h>�z��v��5iӷ9��YB]j���%��x�[�syMa���k�Vx��Cc����C�$�[��Wi��Z�'S�`m�sf�����w3t�������g_�����c�q�݌�.��xO7Cٲf�8��)�dWoj����[=�m����m;i����3��������Gs����!��׼f;����G��Ҿj�xvن�B��=�n�yg�ssĵ���;�0���/���@�k������K^ C���bуfd6�洁�7��#��z�G>�N���7m�!�8Y��*V#bv���4^c����\O��J?�%��
�t�-Sk��r��v��%v�Oj���3�i3��Z T]�S
�N[U�;�f6c�n�k���[B��K���r�י�.��v$�Bb�� ��K`��V�x>�:td�݊r]Xr�\�E3������?Pj_'�:`߱q[�k�♺�۪J�l��`��Vj���=�pv�3��UN/v�'��=����ԿO��	��:���g�P	_3%YOu��V��3W��I�45[G�S����vܪ@{���F���K����w�g�1���fz<�-��pϙW����[@�ʬX�C|��hN�8�%��&/�e"g��\��E-R3���^�%��T��1�TT�_���K��m��ֵ�ǣ�3�pL��_M2�3�����6�%~J���ʭv�=L�8x�{�ѻ�����odW�� .�6<i���Ej��h�Hm;�'j��2]�.h��3~�uIx��
V�dۧ$�9/y�dG�sV�+퓛'mݢͻ:��{I��c�k�{v�I^u�g�e�D>������Fv���_xYd��V�׭T ��X�v�����w�6��� �������Ia���n-t��R��d\OTUm[��T�y=g*�}k��Lx�G�ᒛ��
��@��E����.d��ue�@�;�]��7b)��WIS�{����O,SK�]M����۳���Q����
���1��td�honݮ��\�3cΘ^kka��Up2rO5+�,np��X�/Z3&N1�-QWS��O��_F����KM�M������|��5��o�Y����ff���hn�ޑ���i�2kn���{�:s|xvkI�{�h�cuʈ�"2`>o��[��#�a�9v���K -�<6xɔ���\P��Dt�?K��Ś@��k��,�	��t�9����Q�"�v�!����Nq�u�T�gG��Z]X�lR����<o����Cd���2U����y��NQB��^%n�ʝO��(�;v��gh�>8��ɻ;������Q+wLJ�F쁖��T������1n�dwh;W֮��t�l!�&|�*�Lz|M�fpٞ��$^��f��*�Zw�F=�s�{�v��ww%1���Ksŀy+��9�Oj[Vd�]{K��vǹ�%�)�I�m��EC��	��4�Ǫ���w��[R�
�qw�<�6�`aU��rw�;�D��5�in�̉;�!���]r[�{˼*LV����n=]�6]Utv5��w���DӁ������^�����.k�u`�T�й}����O7����f�<�
����.z���DoC"�R�ͮ\�^�x;X�R&ذ���'Y��QP$1��]�����_[F�4��:�|��xY�Xt�4�nv�b�A�J���dQ�~��;}-�	i�÷7���#7��D�2�1%~���gf�j�1}+M��Ivy�`�/��"�n���/[���zn�7RD=���7���ޚ��%cU��Gd��25�K����3soo�����k�q�R]��z��Ω�lL~5�o��Pȑ���~j���U��O�ء�;o�.j=��RLү��@YoY��_�v��+[f��/�����8m-�C�]\�y�(�w��9P&�������;�a���z���=؎��cA�xw���eN�|���X���[)lm0�j����k�x��D37����>��N� ��h�|��=�4����Z�83e�cl�4���l
����B���#���~������_~6�����MY�}���$�+����B�L����R�������2m�S^�2��� ��6��0m,�n��
��&E{���]v���q���*R/��J�r��i��p�G#��O/3�]��:�Q��N�6�����p��V�t����ͷ{2�/�}T������,�������3�f���v t���Q�2��pǄ����ɢl�MOoZ�4��-����O�;�t�ҧ9ҍ����Ǿ�rt�U^I���+�5^��[+�]�wj����!Gs`x�J7���.݁y#_��Ir��J�y[܊����s�k>^���Y�#Lt�;����ؽ\C�����C�h݉tJ7��K��m)�Zs�ɶ4q�-}���Q-<��GM��[X�w�q�.�@��lɼ�O��b�Bd�սY�:xp���)k(&x)����.j�z�
���������g��� w(Мشe#2�'y���ws��2{{#sv���'1e�&����o6�n-�'}4&�2Z��u�;_՗y�/�f$>����^�U�x�ɸ�����u{���5��f	!�!�U�Ɖ���i��ue�j����lmNg_]�k�P�;]G��A[�Ѕ}�k�m� �ğ��;��q[�E�����67qJS�S--kuA*ˠ��F�$xMN��i�V�
b�%�RZ����c�e�uęq�T훞�nYF��l��_�$A�������؝���,��B)���9Ɖ֭��80b;�wVV�t��:
V�.�e����['��-�}���ûW���� �G/J���X�4/��l����AW?��ǻ͏.ݼ����9�:`3�����Y�up��;�5�m��mq�1�����ǖ\��%�������>l6��G�
�O���M�t���Gnfh��\��q8���;�mqX����������߮��_��B?�XF͙xY(������@ȣ��ͭ�V�i�@��t�]Ԃ(�]]fe��u��'Ε�ץ�n8;�-��ro^F@&�R�֟B�غ���s�n�h����ƥ���j��%��m�cv�lrZ�n�Aǆ�"SY����x�T�����u������(pW��_s_�.@v.k=Օ�[/&t΂f��k���!;��ۘ�h[8{��W}���8�����\��f�G��s�[� e�EiS�VfM�Y�;c�ޜ2��9��eN�f2w�t`�������kok˕����#LrV��6����8�`���Beͮ��1:VՑu����'��L�Z˛K��;�_my9W.�p4�1G�SB�b�F�|�j��B{Nus[6ٜ9Ka�\~L�;8 �T&��`%Ux��Ҝ-�ݝq���ռ����\�dp�v+m���A���8��u�x�H塛�8sL'�p��MDS1��SgP��w�hL���I�owQVѶ���=�����?���4ċj���IZ^����9�*��2^��F�$�)���G6�+
#�����Ѥ�mn#�8�,М6�ʉ;��Ռ��zy̖�=�sHZ�o,�{�4%h!�a�WU·<�T��\�V���8^V�Wg0���(���1���3���
h#ܘ7���k-J&M�y���2VS�L��:N��[Il�2����9[�����+5��-���:J%�#>:];æ5�.��zl���vE�K��!(����d���6��}K(��m���15��T���-.�hD��ST�d�menI�.Is�u҇Rm�o�R�T�.���/��eZ{c����ͽ/l5����i[����_Ӹ\}q�5�`0�3�	���L�Q��M�����a�J���t�~NX�`�KI����},`�U�p[KF�G�F,)��۶s�qN)׷80f�z5�M���a���ѝd�(5��w����v��	"e�O��.���>�َ6����ڗ2}"rqz$�p�ɌW٨�7Y�8�Fq�m�TC�XK�vC��kia�9��d���)�e�ո^�Ӭ��`���'�^֒��:YN:��zP�$���y
����v\]QV`�N�}�;�-:���Ax"�aY�8�X�1֢]�y�m���y���
<E�"�lރ����4h۾��Q�(�Y�0��.�xTxlTkz+7M*'바����i�t��dx��4;q(.�'�7��偑nI¶���4�}P8H�9�[�\b �sUAy���;#�3�e���Z�T�8\����;\��k� ��[�{�9�>�o���Q�/��:wrɷY8��_w�i�R���L�r��P�	%�×e�7k)�@4X��-Ǘ�u{�R*!���+'����/��E��(g_Jn����B��K���?!a����5Pu���YuqL`�Gj��N�źص*�-�ެCش�7�;p3W�-.�1b�ȴԴ1��J
��E��s���94r�u���R�����(��"�eJ��@�Wܕ��t�:�|q�BȄ$h��e9I�n$r	2Q�F�j7 I|ۀ��:��N��ܪ0��Ei	�f�C'��	��H!��ÉZ���&�E��1�m��X�{S�z�Ԟ�mZj#X����Ǐ�}>�O������~����ӵK���b�0ih(��Pj�hh.��O#�0��������}>����?���O�~�jڶ(�S��<�C�߳�+��*-y.5����/!9�#1mp�T\珷������||?_��3?z���6�[~5�MT�T��QF��b����ך5AMhļأ�d���h4�̚�Ab�Z��Is��'I�4Ѩ�Z��<㤤��M�SUQF�ƶ��(�����B���V�E�US�aŶ(�8nF4V(���p�1��m�b�Ōi�1TE4d4co�\Νj(�(m�61Fڝ���[<�lW#��N�[��
I�X�C���E�t�^��͓Z�QG.r�;Fm��K�����H���p3���1cfբ[r=s&��.Th4c,N�%�1�Ť<��~|��0��) ��o��![�3ͮ�iٱ����޾o�L;u|Q�۽E�"�)xDW&��������L�����ˊ�@ZTtTu\e?;�.��a��(�b#��S�4Μ��o��-ƫ��d�G���W�o@��§��)�Ȏ�i�b��vc�F֮cc8�w�K���Eɽ.�q�tf���>�2�0��[۽�m�vC�^�T�7Oa�讈��^�vB�^K�`�����ٺ�ḥ<�l;r�#;7F�W���;����L�W;x�z����ZY�p�t���x�	�&�={{�D-Z�$�:�ܨ|9-���n��'j�.�>�u�\�/��`v���%~^]Aԟc��τ���ݜ���sjݚ�R��b���i�m���F�a��h���[�$��4Ge�6}r6����ϙu���%�o�UZ�zx���!�#�|�W�];Pa���r廫3�Ok3�DE˳��xz�[[n�(�H�e���<�RSs��9�GVܱ�ܽ����Խ�(���S�S�8��(r�50��;O^T�3�'yg���!4CG�&�N�t�?fNn�J*{PN�n��mS7��FW��qL4�M��pe�v.U�cy��v���e&�ː�w�kF0@�®��
�t��sZ�~&��M�V)��"�&�3��F��`��z�f�1ͼ����2ң���F*�4�K��0��j��f�j���ћ͕����&o.���5��;��b�y����ܑh�i�;Z/�7�H�otGO�3�NU���tcզ�|�EO�E)��s��u4��/�ٛş��tгY4mmY� �Ԇ��*X��ό��=v��� �l��Nq�����Q��r�Xl�٥5����U�n�]�^�lwc�Δ��6�9M�W�W��F�ur��g�x����p��cګ����
�P�Y�ǎ���������%˸��Z�i9��Y��N��ɥ�nl�N5��j��(Ϻ�u��a��8i�J��f�{��;`�z�ԠQ�zG��l����8n܋���*O�3i��7��`L���k9=ح��l��\�>�1�h-�W�WF.[���_y��O\�����b���κ��uȅ�`��2��8�8����{Kh'ڹ,���e�Y�*�T����fi����z�nh�"؅Y޻������v�*vt���պ�q�=vє�N4vifg��Qڱ՟>�Ӂ�ؾ#7'��;2or�h�e�Z ��C��=�#zt�6A����d0f	<t��xEo
�ܙ��+�b�n�z
0(��7�h��J���P�C7�4���N�m�y�$��I�-V�z�D�5����C\���Dʱ	P��{�7��W»63��K�	������)5�B�}�Zp��Hf��i}����fn�;جu���A4�����E)��i�*g`$�
OqA;V�g�M��>'szb�ڞ�xZ�=-��Z��p"��=�ޝXF��D�ڡ�NՙJ�^JUb���@�e��{V��2�`w�f
�\9ڭ x8���63a,�o�q]x��׽������xӕɧ^�~�����~Z��K]۾�H>f�_&�����9���2LĻ:���S��b����?��l~��B�]@A�Yz%�g$y��z=�rʿ_B�Q�/J��L�,bv������5c�I����w/,f��O�;��]ܢ8ـ�ɷ����LDq$S�f픹��ugk���!����<�K3m]�[��f=��{�m�8�p\�du�+�� �c��x�k'n�}mM�������=�7�b��t�m{}���#n�j��$��V��|������~�_Yڲ}��˵c�6�>�Kw]vгYl^��#�{��]从YF����線Yi���q3���V��#c��6�S�%ex�m��q^��9=���{Jh�}�f��@�b�i�Z�](�G��wg�y��{����w	��q7j,^˛N�-}+
}����������k���o��l�����2rؑ+L�b�r�Ӗ�2}v�g-D�.��\p�{�d�k�K��q�{LϞ'���f
O��O�m����m�8�mbU��~�%��q�/��#��H�l3��KG�KW"��Q�����t��=ծ�W�\Nlz���+x�*��o[^*��*i̊�fnn��bӽc�_k]�k�˷'_:���d˚�%m[g�w"q=�dfVJ̑;��.csOEJƻa��cr��8�D�Cx
ZU�ٳ�DD����$;����&�ʙ�u��&vàr�(��E���Y�䮋wTK.��Y������er��}��;N���j���]�ZN�-�*
�A6�@����O�v^zN^�T��I+�N��,��3FWq��n0Z�p����M�Va�9N��s��#�Ur�� ���u�ϻ��JWR��6E�������v[y��.9��#5����#�Y[+X6x�]�4k�MSQ�m�I�y7kKc9WuW�8}]Y=�q>�7>x*��|+1}Ćo�ɳ+���~N�n{�/��ks��� I�ew$��>�����`�xn�e3���j+i�>ff�c^x�<_IU�V)�C�2IW��,��vS��|��Zu��J �lQ�@��6�����e�^/LcVO��7�om�_��&'2���U�����\����3n2-1�80����W��z.UZ��|������%��G���@d�<�'�5_ ޚ��/�{uM��z'r�5>��k�L\'�e@�M�z�7���ڒ���Fb�eMF?[�<y�1���e�~:���+0�鑆z�Sb�1zL�ZD���״;*_��0�|' �(���6�����R��U��-s5p��,r`�Y�^�+���=���r�T�) ��e�}�8���f�� �;�3h<t��3k�}Ye��~9�{%B�Z��\c����+�Qև��œ�[32��g���ρ�h>�	a�R�����a�O�2_3�����r�+=Ĭh��aZ3��,�ݵ����jY�,v��[��GT63��۱1B�J2ټ��O�����}��5Kd|��e!X�q<��S�GaNC3v9�ܺ^���^5���G�=Ʃ�ITաƎ4zV�:���Š�mwl���D�����5UD�婢ȷx����z�E�cC�,�?)��Z_�n�J��e��/W�v�����Z�\�V�*�l��;�ֵ����7���"Ll�1�\p=�1�HJ�G9W��u��j.-m�n�x�м*����[�b��i�r ^��pq}^9M��1��`��ӏԣ����5�-qp:��Vi��s\��|CJX�Zޮ�z�Bg�9Sߵ���߽�lǁX;��[��Ց_�wG��̿.�5��8ǐ'C��q�O'JC�tPq/��ka�pG((�efK�c�ʖGACN��JS��E�M_-V����x��ଈ�lyg� JhT�Q�oq�!��iZKn��Ǜ�X!�*���bN��xjX!�L.3q��Jn�{�R��� ���{m����}���|�I��g�"�oLG�Љ�3~Z����s�j�fUf^�⫝y��H�8ї����m��v#^�[�o4�90y�+}�Ķ�ߋ^��b�9�`�������-�KcR�j|~�Z�4�I�9����g��$�@�o�}�{{N��:�c8Cd�R$�5��K�e[�h�V����[�7���z͎:!%L���0lC�=�<��q�,��8}|�������*�/����a�-c��tk��ZE��A��{�{Ȇev=�8��]�̊˼���N�y	�,Qi_�[���xNt�	�\*���U;�X
��SA�L̰�U�qF�9L)�=��o$��+�H&��a�U���-�i��oEKh�l/�f�������f8C��v&{�Yt�ͷ4�|�Fq�3MN\��k����r{ʀ��Wj��K8�A�r7HsLܒ��� �p���I�Ii�2�Z����p#UJ�n���/V�ҧP���92�'::`����W�O���=d�d���~|���v1� 3�\���SSg-�z�kf\�Mz��ZNn�`�����K؃�ŭ�_�l%���qkdR��r���4a��3������n�f�dW���u�o���(-X�F�,=+v�∮����U�Qer�WpD蝩����j8.�b�h�#��Ǌl�����U虣w�A;����r�����mzyq�����4dE6�������_�����J8���Yy#y���Y�ǘ_�}2�i��4�ڻއFۂ�A6��I2*��;������o�3���X"�F����Zlz�
y�vݘ��50a�.W��ܛi���o�>����Lᚵ�Gz�/D�	Ԅ}^�7YU��ҍ�U��/P��g^��n<2>ɴ�y�ت��E�Vl_R�Oݛ�'�E~����M���IF��Q���o�q��f믲��£�[濫�
{�Íg����]�v�f�e�a�48����y�H���̱�(/4��L{����:��̠�)��!�.�.;]�!D��.��f�4F����6��i&�Z��<v�d�Z3�ܾ�^�A�H�+�W�*��N���F(��.������@x�k-�e�%�B�1eM��"��a{.a8�]ps�9�� �ٞ��S_u��~g�}dЄ�DM�}CS�kȆ����y�
w(<��h����4��[N�4ө�h�9��bi���-�a"7tº�7���U�}�V�f��KQ/זG'z��W'%�����˷ic��Us��%����v!�FU��mGӁ�m���3����Y�����m�y,��>�a���V����:Y���2F��q[��z�b1���D+���x������2�Q٫a���DC]swF���3�W��*��
�T�w=�R*`��d�*l��kif��i�Cmk�@eב�۽�A�mW֐I�r_<z�Z�K�8<�,�4m�ǼY�F|�0��ڗ�*�%�ad,��d�W�W��fϝ�j�F�jjm�{c�]i@�X�(Q�Ǜ����Ŷ2�����ݎ���\��S5{m SV������@��G���ȹٚ��J��HO�9ѽG�\��蛽�κ�Y�\��#�,�e0fޗ����(�-�j���P�rb��u�0�JDA;�_ iY���Y�h¶{˶�{F{�������H>.R虈�ga��«n|��5c�1��|��V��<��p�I�={�0/����O�n�C���g6�1֢_7%WO��"ԢS��F���������I}K 2.�ɜ�1�����F��6+��>;H���2�j��hXA���C��
��_L�n���=��q���ܮ��]�5�a��ATdA�uCa�Hxĥ��F�;�Ϊ���w��1�x�x��;��{1�]����2�+y���n��q����Z�Tv�C���PPU7�=u Ul��0l������$����z��.�iu��jy�!g���Z�1���u:`z��I\��\.ݑ�Z���9�ֲFI�0�^%��ٞ�m�M�^�T~�\�ַ��g�ik�6]=[�4)����k0gf�GAo
�l7F�+kj�.�Ք0�� �ؠy�]N�{�R�_E�BP*oZF��L�X&
,�X�F~[�4/t�3C�:.E���wݬX�n9�� ��#@r��Y-��_ֶ�}�A=�w�Y!�*t=v�OvԜ1�Z�6\d-��$ԫA��,J��+��ۡ;K
Mά껺
��?Mvp��0<���;���5���̡I���2��U������ie<e��3��n�aB��ft��s������KY�`1�Jr�p�)D�ج��Q
�ե����[j#���u�>1^�ߴ��]���d�;�b��k���V�F-Pe�ѧ�&[*<���foT�̸[����p��&�+Es�Y�_S���[AL�н�M(�1;��q6:�E��E��s呮��*� �K��4e�9��Mͼ�]�8	��h�Χ>�5;�)�sh��epd��f.�H8Q���쵏�����Jͭ�N���ZF	ͽ�3�dq'��5��軙�ު-�Be���5.�t���@4���nN�P]�e>�r7t�Gq��h[�Ju{� ��[Ğ�oT�˥ѳ��Fm�i9�2��][N<cc��T���q�v���V�8������e)r��M�(+�n^s�Qź�Y����k����!�����I�,g�k��y�<^������]��~i�0���(]�ufE�n����r�j�<�x^������[m}����TYd`�
�w���d���bPzFS����W�yR� ��H������c\զ�}.���j�l<��M)aL$��m>���Za�nV�����ZF��m�Lyli��u���7u�VR)��F����
Rx�d�fw��5�ۨ��[�)X;p���MZ���"��$�f�&�m�vI��쇟	�9]�����S]�yVO�%�q�	�d����s���7`賲ԧ��G[�t��W+�t�iQ�r����,�9�i��o�:Sl�&=T�_BЪ0����,�Rn
�l!a���V�]mHv$B���	ֺ�e:DI��1��N7Z�\�����v�sA�:Kg��O�}O�V��_�{b;���#� q�v8�,��7F��g1���>�^�-˛�Jۿ�}x�v�O�m۩.L�Hp�b�S��Os!�hꬽe�,U�-�x��SxDqd���D��.zj]�MIƓ[%���݉}��9��=fᨣ3mcږR1й��s%�[	�նu���N�����]����x%�ZL
m�S�o*ʠ:k����I���)�r���w�9�yS�<����XJ�,2���|��:���J؄��8�d�j�^�;���.��Եc��vh:p	gn?�S7���.ҫ4�8���}�G{��!ؾ�	X�K��T�[y�3{�����޺�-�7hcf�5.o
WN�A�v��<���r�ñH��F�4���O���ow��Ͽ9��.D5E��z�xEZ�\���le��4\�浂�y���|}<}?O������?\�=N�~��h�Q�i9�LETE;j�QDj��TQ��3��njSY�OO�������3?_�����Fh�)���"����k~��W�Å��S�b<��9XѶ.}x������}>�O�����������b��E�Eh�UTLs:���uA5�(�4v�TEVՊ5���U���r�cj#X�lSEڂ�*m���)��V���Q�kw��TEQ��{�9��1W��A�Q��2MLS�Uz�#��ccl��4�s[D�`�'F�U%PmmkIX�4�Dl�r�QQSO,�E�#i���Thv�L[cZ�b���X�e��-:��j������Q^nr�v�m��.ᙨ�5Y��gMΦ�tE��l��N��Go~�<����pS�b�#�9O$�V����*��X���rM A ��@���w׻W���P.ܓ8�Dc����F�;ϴ�Ŷ�3�Zzp�r����Sj�,�-�c�u��ج�ƍ�~�@���ݻoW_Wm^��S���n�X�V˧���C31���h�v����6:6����Ǳ��G���9W���VcՕ��,|�wfC^�~�\I���������o�896Cy至�Y^w��q��ҳeueGZ�h��n�4����Wz4��b3wO�WsG��k���q]����9ڷ\�{����4�f<�X��2���y���%3���ԝ0�lh�ʖ��ʨ�R�x횼��^�
N4��g��41��z|"y�����U��4�/������H����i��f�|���E��ֻDS��Uu��m��#w��Y=Vs�7�v~3��m��\u�~˒����־�ի�->��3�~$�w��p�,,�Q�}�ݚ���HEͱ�{�p��5��� ��B�� >i�擄�F'����R�$6L�E���m���n��Y� �V6Ѝ��N���_#��sKz��UW�;��jks�j�� 
�R's��c���\	k��*k�떦X���`�V���Ҷѩ���Z���.���Y��U�,�i���M����>i��"���`���SUʰc�����5H�)ަ�@��2�i�cu<��Ѐ7'��:��Px�l�?�֟G�Q��HJ�'�p)�cS(��f�}fv���������u�F�x0�e�@UK٩�Q>�r�vWg�޴ݚ��W���A�\U=XmUz�?�㥶<�C�U�s�s.�tƺn�֒��^����ޚ��D���z� 1��U]P1��v�@:�}lnm�fmY����s;�0	�������ݬ�Y%.6�٣W�fޅ�o��8�gy��`���K\z��t�dQ-S�����
@=+=���؉�]�<�a�4��Ͽ}s�!�<�]�O�W�䟩�h/
�zj�K*�����=�OoH	i@1O�R�2�j��0z���5K��$���n�ٛϽx��:_u��;Z�!����0��j�S;,��������%OG;���������^��{5�Y"y������v��+sS�::����A^x�tz9�j��B�A�f���7-)[�e�Wo���
�HC��T9G�}0ޱ=�*��+���Mf� �������P)p�H��h�[I��E�H8Jr��>]՟lj����4h��DK����oɣֶW�ÉG����.��*��[<��ͣv�+3�P��%�'Sx&�����	�e��Ee{��*�{��<rM����u]+ɥL��{�bo�v��8r��>�c*����Z=�gB� ���y��f[�U�v������	��n-�l@Vf��y����n�L�s<������j8oc5B�#��`�(�S�z .�8�
�V^���T�^�y���;������ �7�������d횱;I����a��x��s�EO&���^f:E�g���T�X�Mv�wf<�]���v�T�F�ag}������~����'�铏j���م�R�2QtB��֓q��@c@��q�����~|��ß�~�L�ת��ܸ\�Z���@��#\o<�n��.��f'�}-�ZOc��d)�}7"B��ߌ�J��?p�kz��BT����n��y[lR�IU���+�jc��X��K_n������4�T�n�>���ݞ�֤���4`��`'�
��k��C�u�0�zp����
�#�{^�s�vGgn��f�y֛���|��͗��yt��m�R
��ƅ�v�5!����)of�ۻ�N��ȿ`�po7��i:N)w;�R��z�'ܮ�� +}a�-x�`�׷Tn�U���{���e��j���X���I_T"��,:�`���Q<��wN����.4j�>�l���^��,��>^x�|y����PKþ�ή=u��kKV��ǀ�?oo�XNL(�Y���N�.� ��2��v͝�7�d��=L�ݟ>���"#Q���:gؕ���A4=W�=�s�~/&�f���$/����'�cýy����I?Y�\������7k&�%ϙ1�I�tu�M��	�mw���1;1����&�5��]�5�]&�w-�bn\I�2G@9�l6����0�}�x߾5�	&�r�}�k_i�7=�^��M��ץ�qJ�@5~u�����8Կ-�>�n�����������:G�dN�e�/gV�h��< �{pt�2�iة��Œ�b�1����omjWR�`ui�aH����f���uA+��[B̉�f��Y���._<�5z�X�+K��n��2W���L1�����"�(����]��HU�:�֥n����V`ȨB'ru��{DnC�CR����%WL.��{e���p9����122��(�<=�͸��U2tۭ��x�,끶뗲Db��أ�r�-)܄˯��P�g�;��[�H#=�J��
צE�;�f�8�p�7D��2�Ȉ���7�Mr�hw� os���8��4⭠��W����d2�����e��(�-�{ytW���W�=*s�H�VZK�����+��\�"|u��5��"�c��Aes�Wi9f�z������f��%uf����"oM�;eF��7��e����<��i����&�oM�,����*e���E'�ˈ��w�^ӷ.�mA�:a�H���lP	N�:�e�g���֖�L���;��{��:б�$n ��W���>����e	��.	�����v�Iecb��Mł�XJ�fI�V�};�,�5r�Xu�y�Ė7�P��ԯG��V1�>�8�̋���8O�*��EP"{�����ܻ��,u�+��n&�%��ͻsY�uwLW�D@
�
}S2!3NO⾪B�*m0���g��^�G6�qq�u�g���|�1E��*c�F"z�Q�����#���|s�f��GW{8�Z�3H�dU*�v���*��4C�kˏ8�2)&�`Z4��g��v��f�ט�cQ��U��}]�f��C�v��mX��P���q���>��q����S�;��nfwzb�l��5�y�|֞!Yx�X3��<�op�����V��U�Q2$�k�[��s:�T�<h�OiLMuP�<�{qWC�u���7��M��h��RWS�T���d9�T����;NK�`�ln���������f��a
&���Snv�h�n�:]�ڪ��:U�#��L�Om�ă��'+��)���ل{�/%*�������B�5g���<��<���_��-�q�|��u�=�	e����9��ۇl��j�<��b2��YQ�<嶥���Z��]gb��T��v���c1N������#6B�T������Ԍ&�b7��w|�]5���1��\s{֞5����8����V8�lh8r���ֻ+EE��/Ve#m��pv���!H!a0Z���$%~��� ��4g�����$'���������l�qlGp6�(zm�w)��6�����q�e]�Y%t�'6���u�o����z�sߨ-#/�/K[CU�F��=��A��L�+��ߖޮ�ZmP���vCt3�e	ռ�QrW*��,�B�|����z�.�n��D��O��C-2C!<�H\@�����݂�=��*��h��:��+��.i��m�!�g_2c�z���|�iMn�B!'{h��EZ�����Nz�۹�;h�s��r��;�F�n��|�SCfmWp6�G�U:^�Ĕ�s��uU@ӗ7=ׯ�ڥ�Z_�ِj��I��T�{��/��y�8�c�3�j&�5V	���0��9��"t� ^��;Y� `��֞�f/;I��Y�D��=�y5��) K?�4�ur;��r��7�����|�g{�I�����g�n�z�#�3j�^�7+rj��,�m��؛b���+7i���t��i��J0#&� ;poj5����1�����o��{a�/\��ŁK�:���P�ffno�,B���i���r�@�2U��'Z�** ��H��4�N��Ql`��U��sg��Ou}w�U�x��Fk�<��8���;���e�ڪ*��Z���cY�{�����j�tbe���qŚ9\�Xٖ0��y��j�N����yY&X��|\��5�sP(��N���\U�0�g�j7�P�!^��b%����l'>�^����ryXds��i�_q[�{j�{a�������G'$��C����wU������s��g���&^�u�6p}�s1�-�i�m�*ҥ�`�}s��]�/g�Ȭ�̎]�x�c_����"�w�[�뻏3�v�����K�Ԃ��K@\�7H�z�v�ԧݼ�Ψ�u�C��b�4V�L]^e�j�x���~܀pZ�6R~���kO[�K�V�:s�m���7���5�j&aʑ���S�٭�꼕���z�Vu\U�]�w6�"Z#�'�l�q��L�Ι�`�I�#oM�D�cU�XLp"(H';v�1�?L�e
z�q5hp�\��I�hΖ%CQ{D�%����e=C��͢���p�Z�W'j{��7�f���RK��9�����E۫|hs���8���RblV�.',bm޽���t��"`�w_M��ה	OS�c�L{���$G`�jb��{�\ �n�:���^�eqʹ���/.����p³�6�3��e��S�4�����G�[�GK|�$1g!���}���l�3��!������}c����e5��L�Soo�8~�O*F��m�~'����Q��A�xpC�^Wu��$R/���{�)#1�ZA�6�狆�w�Oƀ��.��I�`�d<�vf.ԵF��Ȥn���%聣���#�J�E�Ѧ�Wfd{3S)ٵ=��mz��s�dI�#6�#L� ������:S��|������,�&�U��m��Vaf��r�ifz�K�&[��-�U^��4��<�̧�����4�9N�P'=ӱzU���6+�J�xl1�O��P�ZV���:�9����T�����	�o��egr��R c����˯f�I��
�w�^�Njp+�I�ә�k�Q��8�%�W0�Sv�+��$qWh[ߙ?+LD��|k[�
�8c��(�	%2iGZ��6y+M'p�nd6�Ǥ�2pq��鹵���1&�*�3ע��(ғ��j�n��Nu7���T���50n�s*�g�Li��dy��n��k�9���Q�/C�V�v�ܺ"��]���-�i�W���7#m�V���9�JG�T�3�]�x�~�2<�y�C�x�e<���7��(��b��Z�2@e9}��N��јx��_B��9#q��0g���u��e J������U�̉�{~^�d�~]U���˯i�b�ͱ�ك�5�F�R����N��il�u��l��1�y�첮����|�c���lС5��&��oMt6P�Pŭx�}5e#�;As6�=q��j����P,���g�n����t>�?�� ��+�ԫ�7��cѾ��=���'����j`7#T�G�E��T��7���3�M��%o�vр����������y�A5�m�67X�jM,i[i�)kf�<>χOo%�G�� �>�PAG��}D|�Pl""��n��N��y�����C@¤!"��0)B�!�� ��Ȥ!2 �"��CL��4ȁ4�Ȭ�(�{��(��(e^s�A�C��Enqa*@ ���{@!�|�Q��BT �$PBQ �$BQ �!BE ��"J���J���J��*@���@ !(�B(! �B(!*�B�!"�B!(�B�@��J 42 !�B�!
�B!
�B�@���0�(B�@$! ��B	J! �!"40	H�4�B)J���M�HB$!
 ���B0��!�HBQ!	�$B�!	�	� �HB!D�$�BA!	@�%C�?y�v ǻ��+J �� �������f={Á�����������ߟ�,x�?�I��;Re�y����#�A U���"*�/�X@@`�?O!��.zS�/�?��R�W��r<�uG�0��x��ӈvTI=l�
��!,A �@$0	J$$HH���HJ�2�#(���J0)Ȅ�"H0�*���@$@$�B��@�@��C�H2�	 ���! �@��)0		 �0	),P)2(D ���P���B� 
��R���T��
��)@%��R�@	J	H� ��� 	D�D(D�DD��"* P���1a�/�_�p�����"
4(!@� R""G��:�H<��uo����*@����t��� �PL�M�L��D�]=ļ��݂���8��������ӭ1���Ww�l��7���TQ}�?�<�� ��1����J���(���J�F�ëB�T
  
��9?B8!����A U��dg����G �2��	���02��*��4 ��@@w[NWB��V��N D��C����Z�S9Lo� �d�8prI@�
�Ո
��r����}M��"���#�တ�U^��m��t	C���e5����aK� ?�s2}p$%�=�Q�b�%)H��D�RB �������JHBUT�*�J�*��R�HJ�%PU"(�
��R��QRI�A�5�J�J�5RRR6aP�-Y��K��
��mS��̬�dM��%J�m��F؛m��U�kf��k*.�]([&YBҳ��ZB*m�����0QmVl�`��l�Vi(�ڰZF��L�Y��V�j�TVY��ҫZ��U�*�����(mUU)&�(�-��   �OQB��Lsp�m�*K;0ᡳU��W]ѭRn�S�m��m�L���PQ%[�;��hڗU��m����j���M�V�V�Y��h��-�Q�4��+S   ���B�
(P�{�^��(P P�{�pСC��B�
�ռ�EzUd�iZ�MX��J�۪����M*����$B���*kJHm++JF�ٳ�5l��5�u�v�+6l��G�  '{ݴ44��J�F٠bZv���§W3����[�qZ5��Wsv���T�Ԭ-R�m��wV٪�+���U,�շWu ;jS ݩcB�
���ԁ6ֻo  ����W1�ZݷF )�\�WMkU��nu"D�52����UE���:h�0l2�����W\�A�.��6+SB�&�5��x ۞"���ݵ\*����`Q��툑�κ�$I�v�EB��J��҃eu�J.�m�
	��U QΨN���Qh�U*��i��  <��USb���0�w\d�k�ƈ*.�ۺ ��m�ASt8QAIv�ա��4A@u��D�p���A6���i�i�m���]� uǻ V�8  'c�;c@�,� �.p �;�ۅ����4��9�� ��  '.��˴�6cLT��lim�.��  �� ���C@�GAJQ���5����
 ��� ��K�M��l�n� ��\ ��(��Ul�e1���m"ڙ�  y�����hW@��  �1!F�'w4��s� ::w.p QӮݵ����]��gE� t�t�&�4j��5�dm�m�x   ;I�J(�p  .p  Ӹ��C��R� uw  �v�  ��:�U:tܦ J1�]�  < �~@e)R�	� "�ф��Pd21�鉦�f�  �~%)S@  "��2����� 4 I��1��b  �Iʻ%3x�1,\�� F&�7��~���]n�5�3�^\n��G� B�s3����B�pI$��� �!$��BO� �!$d	$�����/���?��Iy�i�ml���"0��L�L�s^�ˍ$��yR�BHf4:�v4��Ӳ�$ �;Z#/x�T��U���=԰Rj8�d�{�*^kd�&��RZi27+Uix��*�@՜���	R��e��,�\�pu�����cUs�d�xU��X6�/kv� ��k�d*=�(�uP��IG��VP�<z e�5f�8�{���wz�޴�SC&��ZBAz��Urm��:VoH��pK46�ո.9���c>� �t�kͫ�4�/J�_'d��-j;/3m �yaV�7��Zu�(b,굡�=Ef`�����x�M�i:Ę�==k�`��ZVe��#�`ȕ��PW�a�t^`�{Ev�5tαm�2� ���m��թ�̴+Ԁ����KZ�C#R\�5���s�fQ��jePceLAnX�m�v��lQ`���hꥑ*Y�%5�H�ɢ�il��ƫ̦�����<v�*QA0�Ǡ����4�**^��Ejn��J����Fk7jx�XP�X�z�gI Th'x3^fɺ���Us^��dJ.��yX��ʼգR�{�E�e��v�6�Wz,�h���Soee	nY�u��X����ySC���SE���T'
�W�������րRSZU� ��Ge�R�ӱY���o�ބ*<5�3p����{@|s\�AKZ~/SwJbW��B9Sv��.H�����wr��X�����A�2��m�� 7 6Tԙ��(�no3	e�cJ�Y˻��}6�v2�%k�wx�G0�7��9W�g�
{)��Zw)�I����(0v�*{�3.�Ͱ0^ER���D?��neb�S��6*4mQ�6��o(崩ߑ;7bъ�
�6q��'.�@�wSYoS���r�:�<�fn�U_U�me�w3>�)ڹ2
�j�֗c52�l�(L�B�3D6P��@�!$%�SQ��.�3S.�Xi��ӏ`̸��O[)�v���m�V��1�A���4+cH\��1ϥ���9xL(]$�f'��-hyL-O�.�B�NvLݖ��gM\�PT�*��fQ	X��:�N��F5I�mZ(r����Ⱥ�]D�p����XYҊ��coj�G&!���J��2*j����Ke�1��r�HM�&M
b쬃N%@�swi�B�̈́��/�.��ٗ�л���O{QcAՉ�'���YWne���޶�ej���31���^\�Fk")���Ǫe@����3C���PӍLz"ݩt���ՅxƝ�R����M�1�yy�:X��j�I�n�U�{Z��{�^4����1pSj�A�� Y�C'B�E,F�+HI���V�ѧ�J��i�y��3&�6�0<Qe�J�P4F��Ȏ�h�p��n�f m� �L�b�JBf�z���ԩH,��(�k") e���/;�Ȳ+&C0��*ᷙW� z%��	��5v�T$��:�є�UWwx��N��z�`�K��t|�4��j�y.��X-N�an��BKui��`�Y�q2��=�ϲ�w6V�Ez ,����3���H^lfM�F�F��&��r�Ci�Y��{a�G~�ݗv�\o!Z+hRѐ��JX-]-ۥ
�hJN�{tɭ����83(�S�F�^�@9U(<GS�
٦��-�k m�u��Z����B��WGF�ł�L��a�a1Ś"�H^��,�@^�u2WkN45�[�����BT&�)-K���b�fV���!U����
�ڙGc̫�i^Tȃ���O�wm�II��u��軓޴��i�m�m��K�ٴ-ᔃn��Fn��kH��su}zR�i���`�b�Q
�E���=���q�y�,2%*�5�bQ4h�ۑbRMY�Bh\���,e:75ޡzq��j.�Ic
jr��U�(j8�S��|��ȝӧ��[͓so�f�:Rԅ�u��u����%�X��1�R+!��EԣZv��h�"ZX��iI�3 6��t�x�)7���F2Y�wrA�{����A#�����.�'�®ηM�k�ԛ՘���uth٬L�����ˉm�w�A�	l*�z��,�G��/	:��o-����ח�d��œ$J*�m�3D�QF[!au�%m���7#�Gdp㣚�($�����_m�y����#v��8���^�E��/v�&�� m��q��Z���[׃iKt4�3 (i4@4(�xPz7p�Jl���w��*��8] ���æ��5��0���B��W���Q��zi���w�+w`8ra�Q��֛H�2�(�VF"C�ue$���z�
���n�j5f����Y����t|��D�	S
���2��0Z�r9�٫�fR��v���B�D%����2�*�r7`"sr�^J9d����sNbX�{�P,��P��Ԯf���D�I�K^�V#Tv��"�
�Ui;��h��b�4E`�{Va�UmkUI㠯vf �6�,��>n�t�b�rӴ��`d�k9���Y���5��R��@%m3�X��{PnHJ��2�7�����Ӵ@�a�S9u�顼�V�}�źU��`:�$B��5�&T�u��5����jⱚXq��EJwo;b\z'ζ�v��Iv�@�b�pC� ��,{JN$&#�։�p�7e�5��R$�E�ɹI��cLشܿ�1#gt��+��,���n'�,\+"��v��<�x���*���\��Y���TEXb����5Sx%�Z۫��r��X����;�"�;F��	�oDr�lb
�w����n�m"��,�]��x�x*V}*k�CJţYPޛ�H��t�)�hQ!�b@r��Va�%��*���%�v���G�LM�I��8����uq�+%]R�&�M:��q�p��{n�"�۹��F����ep��0���Ґ�V���R�$�>GT',��ݹ1�����Ȧ����L�oU�j3L ��VAC)i�Mf���-��f�ѕl:���Gl��0TR-�.�N�dǘCxRWkp�ܨ�ׯ7T6��&�軻+4<�rݷ��[��9T�3��A�̣
/d�F�Պ�Bc����&
�-�,m�3Z>X2̓idH�ފ�2jIML'&�Z�R���V��ՂQ�x�A���2���1
�P�Xk�"M۬�#Q4�n��d��� �Ȕ�<��oTPЫ�,�б��SSHyJ=����܄DEME0�f�T��iY�f�n[+Z�++]t��j (��*ݢ.���[��4�=��u��^��뎅m���0���ӻ$�@���+u���V�Q����7r����b�9��2"�p���4�Y�IaIhA|X�����Go1�!һ��7Vl�vƐ�o����d-&�$�hɊ���*]�I�J�W����jE`]��Z2kŚ�;�&���"��t����-3L��S�d��t<�'u�c���LІ�3d$��K�N��`�x�z�R�N���,��IJ�XR���e*O$r��h$�Ѯ*hɟXr�3oE���k�#���-X���f�N�hQ:����6�WcF1k%��հ^e��RF�B�P�` �@c��-�ۺ�5T���;�P%�����؟*.��#*���.��:��MѱG�B�X���`Y�!a@��6�V���[wZ&�!�.*,���������r�7+5,��b�ld���%YsFؼ�G��ڨ]����gv��a�Ҍ	�4#�C,��nƊ�l5I���P��ۓ�&+�zsp`y����[m�����5����U ���ly��[z���d�e�@�Q��+Kz�Ӎ�od�!�N��t�e�SN�ˢ�Kð<�v��y��mr���Ϝܦ���f��c��Co�MVهF���u�zeְΝ
:My�a�ZS>�)�-P܁d�CW��]ڨk@kM+�wwr<�NS�b�r��c\0K��`dY��G�B�d��WN�MbR��y��ԧYYgi��T�04�6�.���g5��eh��㧯iL��ʂ��#�V0�s���ܷS�҃#�J�Z�@d�B�X&\E��kp��Y ��ݵCY�ٖK��2�&\�F覕k{X�oW��2VfAʆ\��!`�c٨��,�̦s\�vj	�g��[��L�u
t�0pQ&�К���L�%Dk2����*�!��ը�%1�K��sbvᵲ����W-�u�*���ղ�j��w�Mpd�G镶���y�VhT3��D����Y(R���1�C�ѧv�li�2k cW�(��mCIA�Oh���Lݩy�6i��H�
]��y�/���Ȯè%=�^=)�B�5��«F
��F=�ѭ�6�v��^b��F�$Uֳ0c��.[P�h5j�ze��Ãn���6����vJ�tBZB�+������&��0�H5����͚�lk(�Y��F�Nf��*�bf�ۿ��9�z�Y&�.��M������6�rekǫN7s�kE���?'6m�	�2����7&V��8�R�hd|�HB�#DsoV��72�%�M�
�C-�.Ew�s#9/���o�l��0��&�	ܦ.�e����_67�v�����	�Ń���\�݅�V��7U@�CC�f���I:�cM�x%i����X�m7Kv,��S4JY���/,�0,Z�c,ڠH�,v	8m�6���-�q�Q]�MV��6��[���Z�֪{�ASB���r�cp��:m��9pil1Z����̼0upUދ� �A�-�oZ�SZP[��7�iU�`�IA����ݷY�L꺭����{u��J4�2fL��V%jɤ�q��!Z5e� &j�L��
�0��{��#,ٺ��3"B��Wn�5ú���"Ӛ�+���J��0,�-�>S3P����bYQ�yJ�cB���Ws)6[؝�/�
�,5.�VٖA:���F��/\u��ڋ\���n0V})�������1;yEIY��m �`���u����Y'"�KƮ�	�3�����+s��n��o&�u��V*�T�6�����D�V��ŎAj=l-i�e��ܩ�;Xe\�{ldY����S-m`����D�gl��-4�y�� ��h`F��À<;�s�)I����ҤZ_$ K�*Ir-�gMkour�J�һ�s]�r��M��V�'e譺ȥ��)Ml˒�퇛U��F�WQ�w�/&�d�84�V�N�m��њIt�$5B7��SAm��^-�oZ[f�c
��чl6.�a�X]��ZfJԝ�6JB��۱Hբ�e�E��rhCF)����l���ˇ]���� �0�M2�M�^,1VL�*���JV��"ё,yj�t��`��՜x�O2�vbV����cE��hB�cU����ȓ m@����U@��;%���F�� ƍK�7m�M�͊׬�,�$f;�WSv*mk����1&�#�Zu�Gi��ۣ�wfнv�$D��J�L���'Y�j�
VlC��JrZ1�����j����/6����BR�i$�b+`6�
d"d��K)Q�J-�Y4������Ϣ@A�ouA�M�9�-�i*i�P�{0	i���Y Oi�3�Z��e^��z�^ ���2��B�b%�n<�ڬ؞&��z+b�f��X����M4#�LY4�v��2K��-I��*,V��¶U�idR�q&l�O5�[+���S)�U�3hi]�6��|�����N���dH�Wqϛkk�:#"V�m�L��֤f���`�	�͙j��jZhCGe�dJaٰ��^ZuT�D:�]�����j�bЁ����jyQk3"h��_��ʷFFQ*��10���N2����i�H�Q��,"@�j�Oj!X��:Rةܒ3q��'��� ��3��p̒��p�q;������a���"%J�P�N��q��(�.`C KªHj�)MS���\塕���V�e­�� ��1�6�ɔ�W3.�h���tc���ӆ^4Py��4M�!_�5ث_
�-��Q�*���3*�Zo1֊����[��A�N��;r�	k-]8�<��TMЧY>nh���X�ԍen��v� -b�̸	������������ڛ)�r�GN,���
ӣ]�j�dQ
�ݗw�I��:X �ܒJ7�#������v��q4%ifҘ�1��(؇	&6J�-��d�G[4\�r�%���ܴ����n Q�zeM����r;�WL4�l����b�_&��%R�V�HA�r��h�J�4u8n��z�5��'7 ��Z�1��@�F�n-6��HV-51E�hr���A5-���:_���C	\i�(�jT���L?��MRšq��D�Lp��d5N�VbuoӬĎ
�ˢ2�Im��.��b7Z��`��d�/B�7q�۱{���$V�0�˩3iSA�P{,32�B�[��M�p�v�T��қ�[Rb�:K��^+dx.���{@h�d���wR��:��8en7-�
�H!Sl�8D�V�n���-݄�ATedjs�5�`�ڊ�
�4��+ifd�YR�6�uxV�p�`C� �t@�soS�Q���[��-�X3y�fV#�ȉ
�I���;ZZ&�H�k2�]B�9�+����ՙ-��-Q�F��-M�T���Fdph\��Ɗ5�FX�ݣ���&�K����XR���vтU¬a&�+,�jm���&�VL�&��|�iY��hX%J] �M[��:��ShV����1Ժ��VH�1q&VE0��	{L�SsV��o�[�D���x�)��zj�D�M{���O�7�V�ոf�3m�4�\胋�+�2�m�/��fҦ4�u����`UL��@�t��{��J)u����J���6���8��/y
�D�Y�۫W	��k\��\�+8W�@�����)��/�{%M�w�Ѥs��M0��T˹s+V)��`����Q�|��^ip�8�x���]ww�`�{@ø�b��;!r��.[�x��i��\��$tҰ�cJ�nn�VxTY��c��),h, ����R��ͣ�O�7����mmwGwO ���Mc��JV�ځt˔3j�<D���z��N{���9�`*��3��݆Acc�L�Y���i6��,N�6��}ُ�g�T���mJ��m'd�E�ʺN6�IY��ŁCq�Ŗu1��c��f�6�=�m�A�zb��#x�+}��@�ݠ��InO��w;q�&������Y;e+��؛'i����r�7�]F�;�_�K��\�
�c��v�v��m������(��-���`ObܾۛOkD��S{��f.�g�౽���3�
הL罁��FJ
�hRp!P*$�c�hl�ɘD����<�`���9|r���՘�7n�����{�]֣7*�ΑǶ�rǠ�rzFFV�ϐ�B:���0-J_e���ר�А]a��C��2��U��ґ���|8��!��=�w0_�M@��L(uf�e��hQX�d�*YTl�R��)�\
�-�W@Њ<���X}�9�Q��H.��Y|�N*�h1�����ouk�pj쾚�ٝ�op��06����fM�kRuzޞ4d�9p;űn��T�i�#��Y.�z��Jn��1��F���Zec���ޞ�9Y�G��+N��p��+.��z�Em,o8uc ;�7�l#ŀ�EGr��j�SD$EvcU���}���y�Ȩ^�8���pO�U�uzimն��9�'t�]ͻyyV%]�u�YA�J�����T���f6�+���*Ńwl�)�JNdW@�;����lm�"Y�:�5�j�2i�;��Pη9�z�u���&>�k��ץ��Z��1�܍�0���z��Z��k�.��S�c0��y�	ԣ7�S����}�[�K���k��Ƒj��3~�m�.�\�D1n_A��E@r#�q(ֵ[(m��@ej���Yŀ�]A����v*���q(e2�,d�mޞĶ�G		fם�HC�eF�r��Τ�So���3��'P{��U�NG�沔��;�f�����֒�{��.K�]Vɽm���
�fu�{����_S竄j=q谂a1H����/�ӱ����8g�+.���=ɢފBwǊ)�3��wdjRw�L�G�}�譙u/��v����d�њ���
v�ڭ-��^n��˘P5ӏ�ܲ
FJ|���pd�՗�rJ�Ψ��s��^���}�z�ͷ7��;A
�t&�� �&թ��p��W+ 
�NY�}��犸-���^8��1��Z7^���[�,�C;A}��ـE�$���]^)����֡�aN�v�����o-�u_p�S*�]Άb飩�X�a����uu`�X%]
���e�V�ug!��%L�>�F��&�u�l�.���z�G������Q���X�s�����]9uB���܊|�8��>���"qP4ۮ�R�&���*� �]*��A��6��N���NH�6�U�gt�Q�y�^mNM1���h��8��,��4����7B��ˀ4fvS|�L�k2�B�Ts�![t8�(u����_�)a�o�D���c<Ù�x�J�z1�|�ӱ�ڣHu�be��9��ԗ���oLyf7���k�H��y�x�YC���ي���t��=+3�s��"im���ۏovS?`�}���,��%g�e�*o>��Ԫ;��P�]Ħ��Vݍ����N��Vwl|�E���5��چ�������x@;%]���t���!Z�^��^��4+�1@�״b�E�&�R}��+�/Bg�;�����TA��h2��˂�T+����N���@�s\=}�׀��4�*���Er ��,�5V�	Ύ��+�$sQ#Xv�.�8�S�q�B%�)�&^ͻ�ۧK:k'
g��n�a�.np�חw���t�G���r��fA��`�Y��v��h�
��(l�XQ���秴>=/7�=�tt!u�M�lLUt�G�X�;�� ��t�cs3����	y�&��t�f���f��U�6��'r;��Q[؁� �(�Q���5�Z�p+|"јm��u�%�SmrÁ�,��R�;�)�M_�xr�&gO>9`ܘͫ�������v����C 1M���VQ��e&�E�Y�䕂��g/�;���-��Ғ�e��$[59s�@�>�b���MY[9�=���M�� ��41=��������̋]I�Z��T����U݉6�j"�COtu��B�
��
� ����so��.�_c�a�C+W�/#�!�Ew��N҅7�,�u�n<���f���,��R��f-T᱈�����u9�7��Y�]��t@�l�%�\�k��2*��Vrɭ�n��:4D5:mt�w��:*�>�{�NN�ƽ��H`i�Ð�שi�ϖ�n"��ʠ���q�զĢxed	�n+�[�K�d:�+@����W��7m!r���Ԑ8�3��̵�^�6�u	��7M����m��\�)S$D�Wj�/dbOu�ع|qe�=�XPn�٪���,�f f�ve]�2Q�yhI�wd1��Ǉ1�9���>�{·�����ޮsVJ&+|e�o�d�QZC/O�vp/��G+� ��7w8�71����ߤ�:���69�;r�P���N뾧\�]pֻ81|E���w��S�z�Dz2�S��kF�Zǩv*�loӃ{��Uvn�Q��.��wf[����i@����#��жv�7�P@�PϤZ��t�(vs����͕�i:�
ح^K��Ƈg^��+��dD�/*0��,�#vWv�P�1d��FM�C�b��b�]�`I'g�v\�4u'�������x�]S@G.�o]f��@�f����*�z�[����os�ѤN�vd
���f�m�b]�5K,`㫱`AP7���(�"��⥽A�Ă�B�'�&�WY�b�b��E锂9��-�ޙ���Sy��U�(��YQa�V�����īmn!�V,����+������sCv'��:���9�񋷘G�A{F���Dӻ��/A���u�Ɉ�u��ɽ�h�Tuh�]���$T��gQ�"�k��LQ��K���n�fL�����4�v�Q:�E�+sx䥽Ξ�	UΘڐ,���7%E�Cd�8;���zyFp��-cܠ��j���,���r��QoJȨKN�w�Z�Iѱ"Κ6+�8Nl.cy�ֆ\�^ p��3�C�7]��62���{}��B�.���j�4��"WZh̎ob's�r��B	��0��(O]+��@��K��*�YB���adGU&�[גwRvl].עS�KP�5v�+=����D�M��I�ܗ\ʚer�N�X����X�V�C�W'���}�0��J�Rۼ'��]5�u8�ԗ:�ı�C[��sAP<3�I�͔���w���[b�r�=�u��]T��pD�p�<�X1��}:u.@�����!��)�N�����'��n��Oj���^Vꕖ{�J��˕��I�BN��+�Wnd����鰁w�Q#�#��`��!3����S^�:�ޒ	*�@<��X�ٹ-Z��6J{�J6�{L ��k�=LeI45ۻ�u����X�GJxx�s;}7�� ۩6�:ě�
��-��۵���R�.+���!��c�<73�痁Vsf�r��Ycl����ko�Vաt���U��g�Z�K�����ᔰ>��3N�4����ǭ��e3.H7(��tb���X|�^I'HJ̩��N�|��kp�i����״��j�9����f҆��S��	�)��S�)H�Fs}/u�s5�hN�+�KDuYj,�`
T��r Y��[�EE��N�4��n<��r�i#]|0d�ۈ�J��+�p1u
�R?B�Z�ꧣ��Y$ə��"�_elxo�>�]��s�oI\�)��,*��u.��ҙ�'ڰ�e�C���ݳ�+�U#���ŎW٪�w�aFs�W.��Z�c�o��j��}��LQ@>n�.�"p��R������L��Xy�O�N�:)v���nܧ�N+�)4�õ�r�>�-s�&�wr-�7Ϩξ���Xw.�^Ga˨�Y�k�8�&�4�'|�7^���1�@;9���� �P�1�"Ԧ��hnX��3-���ǟ:�&��xc� ��-�d����6��P���WJ+v�Lu�W��w��M�hsr(��Ӆ���]���Yy����B���O�*D�^�k�7�
Hۇ�Y󧗛mEÒ�u�r���	
+���Oz���Sv�)wQ��Z�C�����C��$��3yp�3$�U�X�el;�kң��U�����i�4�\W�$�A��6��|�o)�x�N\��eI�<;{S���ё�l��2*��*�3ϱԢ��h�3)���(�-h�}�uϫt^E`u�}����v.QcK�%f�*>C�PԙZn��m��ʼO,_}���sX����Lt������w	yaG���Լ��[����i�V����ۗ(���}!��E��4�ᛆ9Duk5������1�7r=��ˆ2eE�� Wm'+\{Xi��r�K��XL��i����8�*����y�v���.<	2\��R�.X�y���ܜ�V�!X�� �4F�h�&���v�F�T�t�|��9�Vq�cC��s���M�5�s�:�6�#�N���c�]�c� =C/��%eV:�6���ާ{����e�xWt��:Uε�{�ј��j�}t��+�0&UfG�Sh*�E	��ۜk!����}���i��L�t��/{��u� �:�s�Y|)շs.ڳj��U*�,+���?K���@���z��ӹ� ����\�-�ǳ�{y2�5t�#Y�$�S��:r�4��8���@�*%�M�9<o-�})G*v$���|겸p�4�o���ǌs���C�c�+��:��yo^�-���܎��cX$g�ał]MUor�w|�u@&Ѧv*N�9�����=,��޳n�0�緡\��#Yݦ�S�IQ,6sڸZ�{Zno���<��E�-��޼!�Ք8���ڄ$��ʸ\f�ؑ�V��(:�U"��(��Z	�<��*�]�"�m�w-�� ��)v�����v�iC�@�f�;��,���.��˛fg����	:S���o2&�^	��m�:�Jf)��U�x	3 n���}I�]�ۨ^��-ݸ�v�j���vIz�(J]u�9\tݣ�ܽ5k��|��EL�ۼ&f?�	�P����'�¬��;��er�u`M��.�Ji]��q=�)�Q��ʁk۩,ܔ�p2�2.�'�WL���Z��t���@�ZUكXkAdoc�n��D��P�;�6�6�)ʉ�Ř�����l���]��z��Հ+!���tW�9�2z>FKĖ7��.�]��u} �<S�7L��u�w,�	���[[;��kN�M���ޖ+�[K9������|�¾]s�x;�+[�\ʅ[�mN@�)rs�S��pQDH5EL�M
����6�\��4iv!Q.�v�T�z�YE�`l,�%�,sk9��?�\b
�ͱ���ۍEr�7�ZS�����5/"O.��S۾�3:�-׵��)z;��.���Au�APV�����[�U�����'ECR���c���Oa̻����{LLU�e��Du��sk��]��AP�����lW�5u�άw��;_H����Is�� ��[�H��z����1�%
.�fs�b;J_��
v�+���^̭|a ��eqqsԱ.�����f['�{�nH3���])��¹r���/k)�0�\��rٝ&��uqgW3�m"d�jY/�(�Y��+yԈqʷd�Iv�r[Q�'&�Z�u�3g���TuS!�������r�Œ��:����JZ7k�yt8��ҹ�YGLS����L�C���?��V��] �2�K;�������X����vpU�A�v�F�n�bUa\�4�)�5�d�bd6Ɖ�n7��ɏx��#vv��'u�����B��w���3�eB�u`ǥ� ��:�A�wL��6�7ق������1�S���1�:�
K�ɛ9��ʔ ۰�\Vq�e��s^嬙$��vR��=�d�8p��3������8�U����yն�3�&˱O�<�W]�i��Z�^�-!��C��}۬������ݼ��!�����6�
[U�]��npM�ۚ��Z�t{m����NP��;a�W4�փaoj8�>�;��N��j�K�{�4��&���<T<1���9�3^qmCۺqޕ�K�}>8��k Z#\;P�f���ĉf��q)�5".em��6I���Q�*S��Y<:�}7{�&;�����8��V��}�k+] �R�����)(
�׶�ueېP��JΗ����W�#u^;���)�^���ag���Y{����u_T.�<����#����w]�P���OWs[-̹H�(��a��|��R�����Tod��'	����y�h]rP;6(���c��ur����B59�[���#̻��h��ys7;���]��[��{��}�s�~<������HI$$?���������\}T�)�7�����o�=�LfVRw��m[3c�U��,2������1�t�^�L�tU��X�%�����1��z`{�GU>�\9��C-ʰD�o�K���ȗ��g>���a���5�ϲ���l8q�]�S��^������tzīU�%� ���pZ�}���G�x;68R�{�g#Ha�����k��7uݕoƮ+��@�U@9n��k*7c��ءu����M�v�sw�1v1kk3�Zp�z9\�pX�<ŗ+�0�Y8�Y�tϘg~|S[X�K�x�W55�=zf�d�4xia��	�j��zӶ�Z�t6~e�t�U�h��3_��5���2���Q���2��۷t�H��ދ1r��3$�/l�8�	b�gwA�sv�m���O]E�59<m�P��"�� �6�����V��O}§e�|��\�����@{�왝��wAϫR���J�r��v.��3�k��7'Z����f�D
��O0��bA޵�u<��f�^�]�wB�s;
�Vj%R.�����co�|�c+���w�����O`xx]wK��rJ���}�6کH[4H���1s\��I�t�&3NJ����q��Q���7��oK��:��(�k�鲱(on �c�Uw]�S�����u�]7e'r��T�j��S+5�߳h����	���#E��'�tU������@%q��o
옗m�I��e:j�_)�Z���S�	%`�0;rL�خ�JJ�
F���V�F4�ˬ͈YB�h�옜�4|J�8)I1���n�Tm^sYV��Q��W>�-Ib��Y�]���ŋ��U����T�|�Y`���9�e`�y�4�W�M�b��X�Ew���<o��\Œ�s  FR7�����,�T�F�Oq�'J�
u�:׼�C��NqY��\��X<7��֥�
�u��rIһ���g�t�K�sq_:a��:��T�u7� �Fa�
嶯C����T�r�n[2WQx:��7J.�[+��12�7,]�/5���p�ܒ�Zr�n��_'ٔW�n��3)۰�,�8��[- y��Gq��ve��Rc�Kr�c���rQ4rȂ�,��e
Љ�ǹݴ��GL�Зj���Z����4����E����E�%�^ᨆ�-�W��z��F%n�v�8-��o���k1=�u
��>�4�/����CW)r�%M�r�2��,�y8��7*���v�u>}������n����w����W�s�\�Sqb���sV�nN�uLE����ǔ��7o�m�F3vY���l�n��n�fہ�U�7�]qJo|R�զ�5�+r�]�F�J]H�I_�/xB�A]fP�ӹv8	�b�"&
T)oj!�lˣ��2�L�\+zg/�ZѶ�dv"n�O1�ty�M&�ͣme�+j�BŰ�h�ׇ��h�E������1�Y�>4���c���(b��7{�N��`��6(1͆r[����Xo{d�+Ә��uq�2��l]�_H���ʚu�4_k4��7����lb܋,[@����@C�A� �ƎR������+�0�
:YC�q�X�c�奥+�b�{��P��Z����P� �˛Y\�W�����5edb��|R[�Lp��^�A��MY���a�t2���ȲN\���X�+͚vrl�{���m��J�����}zhB�����y즖�R�΃�M��;��/�����YW;�7pg)�V75+������M] ��J�����������������tC-����.��X��Vڒ�۪�P��Rsf)��ĳv�#��wWז�����1X���� ��E܉���3/���](�Ag.,�
��՜�>R!+�	���V��	-�v,�	��C��3��Na]�`�F�t��#N`[]Ċ̅jXG=�ceh����e[ξ�wDGL3nlԵT��P��F�,Q��L���@����\�.5ȵv��Q�Wy���pѴ�}������H��|���|��T�̩r�v$�S�]�^�;9��pt;J���U��v��X���HĽ�)^�rY�IϜ���/�$�����C7"PU�Gՙ{�P��4֝�j���6�-	w��W)7^��5�;���[Ƃ�U��0���ږ��c�+��\^U7�Y�M�YS��̴VGw�a9�������bmT9��{suV�[ȶʋ1��溷��ʺΘ*�9k�rj������2���7��,ɕb@q�ɉM��7:��.��9�vXtN��U��HhgHr���l��k�mB��+��ϔZ6�q��WhK�m�J���ce��^��m5{RP���8�um@�n��a� �$��A�8�!]LZ�{����z��!ɶ����=�=Y�,"��t5�2��3N�ᙺ:u+×��(I�����lݤ��g�Z�(�kyX�"�fr�-��]Jr`S�.���+@�\s��[w�~im�sd����2�fTٵ-���Z	mn9�F吵�[���s��4�	aӰ�n�@�����Y7.Ȑ,�o��i�Τ
��K\�4�I,5���]B���)8�̧q �`R<�L��싻w]�Y��f���Yo�5�iq����e9�qUr���47�P��m��#�����5�T�R7����pp��!��vq��Cv��O;� w\��=��n�Ξ[����U���B���0�½ْXw� Q�iҙ�A�C���v=J]ޗ%�/M)w���i��PC�Ŋ[�ë1l9�J�A��n��pY��(��6�7@=t�®��Z1hv,@+6�C�����2.]a�����2dF��_(�GOn�g�d����C�B�Y+'^Ԯqv�s�W�٩����p�N����j�]�6��lLR����hW2�a�����^�8\�qY�ɿ+c붾df�{�ʳ퀳|9���ܥ.�]n�q�2��aҚN����N��;/^*ϋ�ch�w4R%M;]�@:�i�+�(WB"
;�7�+���aL�8�pٷ����9G���'�A�y�
T4��C���1�B݂���7�p��Nb��	��
��oq�͞쬢��2�-V޾�7,�L�S�U�o��Jn*m�Z\������jb�c4)[�R�.K,�R�`b�%nL2 �fL�kB�!4�yS�z�j�K��7��X��Ve�Y��
n�:_m�N&���M�Vfm�(�Ҹݭ����,4�ƸZ�W�t��u�O��S�,@�tV�䡰ɬ�u��kX�c�C{зf�VM��T��M�M��0��7�5���ӭ]�����Ί�r��j�ը��i����걏C=H�=�Rq��Μ����⡖�|��e^.�4s��t�QH\�S4�c��Z�܅�gt�=ʏn]��b��L�u�M���
��ǇG��bү[����U���e��&SWb�!	��"����7D�y��n�P�%9�lrg/��-��ղ��Qy}(�Q�F�=��YJ��J��]�5�7�W��t`0��M���%�~s�<�� �I��Q��Ѧ\T��%����A�A��W���Mnd����ok�5�	��K��v�X]�/��u���n���;]��d���m��dWT"��#d��O;a��*��;�hY�
#�7�Oe|�*ۥ}}4����L�̥{�Y�,�!��N�5�Rf�ح��).O���&��W[É�)n侭�N�A�e�2���d<��Ǥn�QV�kx��]ټ%;�� "�V�̨��.WYZ���_!פ8^��Bw��OQC,��_[O�wl�J���-�,�ս�Qb�CsYg+U�䅷m�6jU�*PofYMj�S�r6�^�G(��D��B��]��d0\j�hs�Wi>HGeP?u�Ԙv��Gl��Zu��ŻX�0;�赈�Vu�j�
R�ð�����ң�0���V����p�2qƯ���z�r��Rtڰ��5������1�L�_<�;C�\���C$ߞT�-٣��8���5hT(�:3Ip3���FV��n 2��p���k�eU�АR��`�|ĩc:f����!��:�g#>3�B;i���ʺz��%J�1�l��������{D|
�`��#x�` ]��L��J�iΤ����'��	��Gv{%��=5#�q�s�T��77���&���H6�=�gp�ε��Kt�u��@Y�7�;v!]y����R�H2%�g�IGj�܏X�I�gY�+_��c�VV4a�;N�n3�Z���ńj��{��uvKb��4wj�W��ṑ��7�SX�{ƒ��Rݾ9�ًk�G��F��
΍l�9b�|$��j��0�V�1������8���+�u�呒���`��v�n�x������e@�KB�YA[�tSF��뺾)p��X���
A�׊
��o)�KK2�ᗪ���W��[x��N�a�0
S�	;Sz:���5 ��U�V
+I�ʥ�9���(���N�Gt��c��-\�fM`}{n�r���ωu��۷�/�n��S�_,[I[�v(�x^AYt��v�Q�'*w��sF�9h*I\]YG��y��������U�9J%hj{�W�<sk�ϴ��Gt��̡��;Red]�S:�U록����TՐ��'�M���|��e�ń�M�Q�1ض�qA��32���$FnY��y.E�q�%��*-ǒ��Vy�c���M%/Q��\Y�����mі-VQ@ҫM���	^�,6�9��eI�u��#ɻ���9�Q�H�AH���Q�uv��l�"� ���XK�d�S��3�kIwIu��h��[A>`/.�*n��mJ�.[[�:(�u�/
������_`W�K�^=qr� r��+�+JD`;v�.b�0�������n+������l��ô��S�q�.&�љj+k-��U��U�=ض�{�d뗕@�Afuĥ����O��ا�0�_5o��8 ���E��u �&fGi�s1��b���b��׺�]@!k�43���[6^E%*u����I%f7iVE����5���Y�^)9��8�q��`�yu��i��*y_h�K�㹷���Y��7���yL=#5�kr�b�\��Yc�ΨƩJJ�9���Z�FX�i��ZS37F�����A�2!����N�-����	t�ҫJȊ�.��U��Z��n�'%lu,�q��v�؛�R����P����:�k-t�ue�i=!�@V1-�2mڵ��'B�PPh��N��&�'&�.��3��8��y����(3moTHٗ#S�o^<SB����LC����f��DJ�}�	�Ҧ3Z@�"cS/sHL�r�F�����Y��Y�=�Y�q���補t����m�uz�	�PgS�7���z�ڶ�Jr����4Gс��+8]N��slC����T�YU�r��j�Gk���iս:�X�bXV1n�w�y te�[?dO7u�n5ɷ�6V��w�!��-96��VZP�<����U�2����Loca��N_N����t���x��9=���Y's�,*�#��ZNZ90�*�0^4V,�j�Z���wz�gM�P̅�e��`Ϯ�]����8���ZH��
�Prqu:X3��,f�=%fjQ�����l�&��0�5��Sd�+�V&�EJX�T�ȁ��gCy�M�z6���㾑a�寰�8���Vm�@���9�k��r�%o9�6u=�z��zY5a�j���[����=L�}YD����N�Vf�g59�[	֙�Ɏ�ݎb�,�YO��n��G��fSSd��_��%�:�m����#f��g3t�]X��y��I�����k�叻�p}h}w�Y�9�+f0 �`ڀ�_�(¨��WI�m�]b�ӝS\��*�(೰v
uCM���L�_'�)�r����p�ʓ��]0��䗋�r���닊�b�~Ď�����{ѐ6i�VM���A �0�%�7-ҾŒ��o3u��=��֥{�{��/7R[�r־MO�ޗxѤ����M+�S,u��Nh��5�fV��	ޮ�&WE5���ڮ@Nn��[.�Gj�Ld��L���,�׈;LL<mT{��VV�l�+y�76�5.V��V�\��t�'^���rt:��:Ф�C�ƴ!O����U��E�F�ő�x�����I �	j�x]�0q�/��;��s�ubc�(]�<g[�WK��B�(fbK��h�]�V���s����rvv���Nt9mK��k|�e��rr�>��e�u����iH�U�P�P��ax���s;�d�W
af_L�;�d�	N��)R	Pԋ��.�!��mvM��%M�7nM�꺱J�v7eM|�VM ^���Y���vLe����,)V�MvӴ�����C��$\�oEAʝ�X�w����qM�E�H�\�{OB�*`U3��3�\9G��0;�Z���Ca@�2
��t�f�?�+]�LR�U��:|��6����yl�Y��wP��=N�u�1C-l0ܿ�Y�մ�ÕzkeL�H�g8ª]�M䮑FY
'�[zУm�fPc_[�lk��\9]C�lS	wxN�M�
�w��*#f��Ü0K}Ьw�b,N��/	�)[0�L��Y2Vۘ����K�R��w3��n�
G.�6�뽣h`��σ��Vk���Y��-��WFn��ָ�l�G�+��/6
�"���BSY[�4%6��]���R�cɸ���Q�̽U��u�}luĥ+���
�q�;}W9�n��Z�͜��b�yz�����S	���Ȋ4T�J��T����U�}_W�|��%��3�S�(`��yL�ge�p�Ҙ��懠�M�Ϫ_l��P3
zNB4&�-䙄���<D���5�@�U,�Ytv��3�oX�7���	+)�����H�vJ�+)�&V��n��-o)��u���a�m`�"K����k+$d�}.jUq�ެt��WF��dњ�ꡎ)5,����c�D��u��-Vep)��6R��41�R����b�U���p1yZ�,��yy�e�*D�E%S�)�7*U՚���r��eϜlL��$_F��a�e�"�=Au���A��k��FR$��g` h9/X�����ҥ�04ф��P�R]h��3wz�8��
�u�ǍkF�nC�Ի��\�H����j67��;}Q}zUd���E(;�t�d�rq�C&+���>��5�q��@p.iݩE���Z���^�xpi쮵r�,$WF{:��K�1L�*��H��:�33X�|eĭ۝x6֞�/J}-�Xh��E�˙�z�S����i9N8�!3';�l�n��=d ���`e����M-���N����v�v�l�ҩZ��X
ƶ��Mn�g-�gfE/Ĭ�k�>v�ح=���tdRS2�$4�Ҭ*�t�"���8Hi_j�6V�Q�@�s#���A��~<���������Pm��&�qθ� ZW$��d��El�:L-�GK��.�X�b�����
�`ѭ,�,kEFڋm*�Z�-������UYUm��
�"�Q`�V��b�QLJ����T1%c�R���EH�b1E"�Qj�(TD�DF1-*LjL[b��(2ZETA,1���be�-h1X������@D���QG,�b�j3� �.Z��R��Ƶ�X�D\��m�cQ�*�@�
�l�kZ(�",̦D�X*�T+UU�ef!������Z�QYU��ĨUAH��ʣ-
fd��J��`�%�Affa-�l�B����&5Q�QT�R*!iE[e�PD�j-��h��KH�,Kj�X)�����ƑE��ņS2@�J���bWf1j���Q��,U��UQV* ����C�D�ZX�PFLJ��U���SD�+��.4Q#Z�AU%dP*�aE���q+�UI�n\�d��Lpa�m��hfJ���#Z,�LI�b�DADAL��m"���刨�*c�k����_=�������4��ι"T���];���4�����âf�ީѻ���4��E��>����E��L-��?}oy���ت_ޱ�� ���?-�lϬ�ʵZ)ҝ{\�[�]���4M���)�U`���q0���f��*��%�-���x��=���5ai�do|ѡh�Oe^�]������� ��uX"²׺?#����V	A�u-�΢���3(ºU�3�1*�0u����$m��}�s��f��m�ǔl�� �ܖ�T�8FY[�b��
��n��0�b�����6uׅ�^粪g�R�X���Θh�xH�1�2�.2��܎׭)�S���,\����6P����q��7Huƪ�c{7����䮨���1��Ղˠ�򑳝m����s�y���DxU�e����>]w���X��\�9���N��
�f�_>�i�W���U�3����#ز�p��N��������n���t���ǽ���4�!�͟�7��o U3ҺUZ\~u{|�_f�G��U�f(��/9ʼ���K=�۔�Gc֫����<w؀\w�0+"P�Y�_�����k��t��$Y�e}�^^V]Y�G�%$^5��}����qX~�GCZr�.ʉ��JSi6�75�J|r֛7[���a�x���6f\`��ĥY��	�re��A8�mօ̡r������;�^l�9;T���#����
y�9�z͇�(;�y�ƶW3�n����?\��#rJ�Q�����qs,�qY�׮�Bq3 ��ε5�l�Np1|ڿ�5�����0ݼ�2c��������$=��O��?�\j�r��s��"	���]Qu��s�����rCj�tw����|P�������uO�dg��|��6�>�[���^�h�Q�ݿ�~��g��W�u�*�tE#!ITB��c+�2�gcA*������7z��|��X�@�_?���.2]b.N��Q��z: 3�Ӆ�O"<�m��Q��e�Mg1(
k)^Q���4L:��Nna3��ҧ ;�+��rU��c�ϓu���!���Uxī͜A�t��}&00�JHs�j���z��wT��^��D��9�W��uӽؗv�Zg�s�Evke��/���V*���_L�"��'i�� 4��(k����X�+��!'M۪<v�j�W׆ �=�V> *���׀w�����;�-��<���h]��R_�N��4��#�Q�=]��T �#�&�]�۰��4�uٳ 
��P����.Rz��o�R�Fɏ����ݶ�$]�D���u���R����$�g)��WP崸<ge5���(��כƤ�R���T�:W�٠�]�/�P�x%vڔ�vP'�/c���PN�@���.ͩ�q���:��k5,�?3��ip2i��-J��s>�en��6u���_!0��⃳9ܑ�TC��\IC*氬'\�@.�=�4�{����B�OF��f��Sk7��=�b�n��_O�g��3�5b���n��n�a��Am9�j��-���Xq�8���/�Ι
�f�?g1/Nd�1y��?_�ba�Q�̸�j��݌���U�G������C�F��L���Ľ1m�5�v_\��;��O�Ƹ��q��~��6)��U�>_:w0M[�����ު�C��?Ʊ>~��ʹ�ͪ�	:�Tr���]G����@JC,�G�q�a�>��wSu��: kPU;�,�Kb���$�"�5�t�9��	]���e�e;�#H*���(�u�
���pw��f�����e�il�\��%��8�C
�t@��ܐ-A��"��J0�'�.�պs�F���4 �Xb�1s���Ϣ]+sD��H��n{�Qu֟�-��t�S[�s���X��^�h��yT>��U�;n̶%���3���7���S��[[N�+�ָ���tj�	�^y�+ԓ�uy��t����^t�(o
�S������BV��;�țw}�[y�i�Tl��ܼnJ��5َ�&�2��0;����}�me��z�Uyַ�!Is�g\����9�'G��'�m*�{N[��9���~ö���u�~�s�k
涘��FP�2!��� �����U33oEA�jU_c����!z@��N�p�X���y��i�4����_��^�ƭ���rNXt���P��V
��l�7�P���d��w�A��Sڕ'7�}��7��QM\��8�J�cs\��7G���_?zٳ+܉5a���ڷ��Zb��;��a�uȭ9=7�OCU�(�������*�1�.ܠv���:X�/>/��2��DV蹾&y�����z.�@o��NҮ��~��f�����)V��^�2⪞g8V�93*���, NR�J봚�
dKZJ�T��6d!��j�oN�1�/�t��f��^}�/s�OD�g�揳B���>R��y�JY�]+�F�u�7�o��/j��Vw%`j�K��4�:T�	^w����hVJ���ܟڮ��ϝRg�˯�Hv��+~&�=�eL���Op��������GV��{n�\M���o	'��f��V��WE\�:�֮�<�i'�x�K{h�����mLv��h�)Gc�o����ӨWq��ѐ�d3w����D�SsoEj̇�e�Zz	�L�Vw��ӌwvU��p���F�!��P�s��s(�
��}�˦Ѝs�
�s��"�ghr}"��҃�:0*�N�1��s9~�1NP�pӢ��)`����j-�jzsN�n��<C�'��qxr�B�2X���l5��{\T�čww0�T��M�-�{4����.�ҭ�Qˋ��ٞ&$hV@Zb�pu�Rk��PVX<�`	GTZ�U��W*���1��� ���]8H�lLLR��7�ݱ0�O����U�t�u枝�53��HAX`�@p�X�܀L1��Ϻ�X/�Q����hwF����(D��{sִJCVO��vl�>�7��T�����G�y����ǅ�o��8�3�K��Z�`�J���3/Mfg��`3���M�uZD3�6lp�:�:��\�4I<%6x�vW	�q�T*;�D�y�������c��ϟ=�S�\�J���J�d8jW��cq�"���<z;�f�U"��88s��aYw�
�\�U> <�d�U�z7��9LҒ��ٕaU�"�AsRm���zF�׍f	�W�8oZ	���j�X+���Fۉ�utd.Vm�:�10'c��7��j�W14�l�#��-�:�����#�5��ݡ��MeV��W{G7z`��&��\ݻ�G	m}}|.�	��S%�!�N�"㻆�Me,��Ћ��m�{��as����}����|8|��O/�Q�[��/U��+��x;�q+��~/4/�>��g��gV���}'����j,����@ۄpwl����h�S���/�Sv�:�t�(`ߵ�N�]��(8��3ҺUZC������F�f��:�r^s�������*4\3\c�s�� zOW3`v#m������*N��m��C��e�&�W݀�6!C9����W_T�#.�VY�]P'6:g2_Sv�n��^%O�5\ _?-�����N�;���6�dYߛ�y]驗�w $��k���imf:��hB;'�=���h<���eBꋨЅDJu�[(hb��#I�ܵ�s�t,=_x�yϔ����Z��0�;��7D��V/�nc�UxgG�{3�J��aGOe�V�Q�*!��0��rG�`�T��93vn�)��ƽx�����v<%��_{�.�b˛��传9��;n�0x ��ҏ�9�E�^ �� �?/kyܑ
u��1_Zޔ��?:�b����ov�53��K�7v\���wL�����e��),{��Y��*g��),v�I`��*\����ڂii������x$ѝx�Ab�opʏ&�ٱI}������Ź%>O�\��+�kӅ'}�a�]{g��nܭ�Տ�1��Igur�1�~{Ӭ�2��T*�N�6~vuo;���ϻ��>iV����R��e��d
�m�`�(l�a��
�jJHsڠ!��tA�N�rܿW��w��M�M΂,ϖn+ƖW�֩�f��w]0�}
d��O^
�|ծ�=}#pu	R/�hU,�bk�5�k�{�<f����Ku�~_8i�;��V= H�sN��,TJ����E�c�qw1�?�����2 X��'LW�d��JδV�P���B���N���Ɇ�bz��@�J�cqγ�~��mEo���Q�!���rPʋ�ª�S���j���,�p�@�:��x��[I��f7M7��F;���,Gq�u���p���v�k-�nwk��\bƇs8�����:dN)l�p���v"۱��_�O�G�zȱAt���.s�e{ز��z��$��f*��2�<�x��0^9za��E���h���T\�R��8fj���H�5���]U[r�΁�������y��~[\jږ3��d����
��M�{J�C����3́���p,�*���2�1�R�gݺ���^�":���P�x���
���+�&��s�W[�*��v&GW2[]��"�ƞ1�Z1%�z�E�ޤK�W:�cɼ��9ו�暼�˴�I������]&ŝ{Y�)2����k,�o_P %!� �'�=�A�̼�H�}�0�|+$�[W��s�z���4q�!#Qn'��o*$,�<��"���=�ö�r��@Yz�����:��g{e3}�����|�ƈ�p܌*�吲eQ���a
0x,UOC6����	t�4��1��%وag׼��s
��Ü�M���A�2�0bE���;7�+�z������侵Ma4�~�H;��+ �? ��g��A�ȓT�PɅ�����B.\�2���%׮��wdR����}�O�у�yg��Xn��t�W�k�2��H��G��:��	�XԅɌ 8JG�2�nD�������cE+���ð8�9y��
-*�C�p�6�i�n����� ,�f�~e����g�F�e]Z�I{3U��l���Dޘ�s���@z������Ԓ
W뻖A��9ף��9��N�V(�c�(V�r5O��������F�Wq8�j@�$}ʝ�b�@���\��n�Ɯ=�6�:*��-���sr�o����Ǆ_vNa��*��7^��tK��ZYq}�]J޶zQ�z��*�{N`e��(����2��<���Z�y6�w�y)ѝ�z9��]Ö6ξ7��,��D��}na�� b��n;f��]/L1c���^�<8�cY`�~=(OB�FY�VԴBi�ƕv1�%~3�>��f�O�1� `8���/mt��5���B~V�FKs��
7�`��gG 7����#�'ħ��oW^]�f����<c\k�8\D�TSonD<�s�O@�WL�檊>�[u��ncR�ē�e<�/K���t����6ܡO��x;Z�W�
���X�M�	��Lo�Ԝ�s�*�@a�FY�P�����g��W�1O�,C�.J�Y��f�)O<�}��]��YpT�d��Օ�T��qS�`ch���,�����y�N^�F��ra��i��a���)��g��Oi�����&�(���߯����= %��Z�����g�>�v=`;��|�����G�nR@v�<'��J�5�w(*�J�5�`��u�,���C��c�yƑ5���/
�G� o�:z "_e����![���iZXW�e����btވw|եs!k���]H.q���%LN<pT�8��� *���'קfv#��n������M*Q�oE�R�k���d���D���Kb�YN�GV!��x���i��7�}xr+q�qBtH�F�CEN�WnaW2�:�u46�����0 3t�
a����ruf�(��H�kZÇ>j@h�X��* �����W�X��E����#1m�l�KA�X�"��ޫ2�Rƙ��<%w�j��D7�S�۪��ʑ_Q�R��(}=�SO��b��#���,S���Xf��"�Δ�e '��y53��R����Bi�gLQiݽ�n����F�ݿ��EA(�C����G�X�[(1(�q����Uݲ�r�~5l��d��]y��_�CU�|��7�4l䤾aS0V��� �?�1����Iaﲶgs�Z��^�n�z��W�]���^W��*Q܇U�OL�3~��_3S���3N=�ǃ=��Z��Ǖ�[\N�q;c0��݅D7(h�׆�N��A���v�g�r��U�˞�s<w��O���)�b�.@8y�S(c��ƴ�_:��=�%�(F�:�G0r��U�ʹ) �OiW,�k+���<�\�e�W_T@�1�32�FFè���+Z����\5��V����m�_SU��z�Ǟ.���?��_ؠ�9ŀ0}�^�x+/��t�L�U�2�a@����������N��X5�+j�F���
�˒6� ����df�܋ܦ��ٮ�\"����20�L霟P7.;]��bc�&�3�S�i�7F�T��k̽�^ΰ�>��&��bLdǟu�ڠ�msi�_sc>�gj�:V��6�j(W�ܦp݊�3��t/Id�Uj������٩�B�+k#��J�U��v��|����ͤ~z�����N
��K�F�>�Z��a���q3;���@1��;� ��z+2���:��[	N���`ӫ�w-v>sP�>,B��R����l[i��m�M�ͩ�5�+��5y���2�����<�Je��\q՗K5b����fY1��_QNi���mc�2��+O��Ѹ��m�7�
���;\'N9��[��9{+�
b�Bu����U���Uq�6��fݱ3&��\��&R�61g ��ǝ�|v�����*�nP�,��Zo�6���w(�<�dyM�n���P)ܛ��hn��PfM���ZC6M�c:�U�D!��I�ռ�N�fؖ��
�7��V����V��&p�m;7��Q
ell��uD4vuL�(�21�K���ݶ{�[�-�Rh�z1�o�l& ��l������[oΎ]gnd���> �/e��U�E*�O�[�����u�����鎪�J2���
wEPBQ���r���J�:�YV����vKyc��P�n�X�Ed�͕�0+��iZ 1rW+�\8b�K���	>ʻH�Yº�NZ{(�.��e���Omv�]�q�<���.��	c�ID�Wv5^6^nG�Q˱�ښ��9v��ld�u:��4�.ѓu/u����}^ew.��!�X�io�0;ً,IfM�Ք���%�t���Z�}3��*���.����t[�qe۝|%.��2��	��U��Ԕ�4o���(j�^m{�Vؙw�E:[�'�ryEu�W�"\6��Q��s�NT�����ȥ�i���=hZ{��;C@O���1m$���g#r���b׺���oʽUu��ދ�)�ǻPT^'��Tɗ���ˮ��;y����[�� ��#�s�(�of�ґ�h�����B�ک�(�e�޺�ռ "��C��C�=����р��<�Y���-��81u��ЫyQlTU�Ʉ֔U���YD��\@lj-�y��m*,�*b�b�ݝhJ`+G{���GoN�H�N�3z�������>�}}�� "܃�@�\v��S��mL�7s[�Y8p;t72�o<E��oΉ���Q�9���\�^��-�Bg�eŠa�S9�����X_ z�v��j��=��L�Ǡ����+��QS�)��`r��n|�h�2�^����N��v5v�f�74�Tɚ���I�6�9ja�����f>n���c�rX8+��k�m���m���j'�o\�i�h���'�A-ٻ������%v�ᆔ��λ��F��_s���ut1AW��V
Ŋ��Q��U`�VTd�����TU��i��(�I\d��*J�(��2 Vh���
m*��QAb�b�r�Vc%TP��X�,ƥk��X*1H�PE���-�EH�-�
�TE��W3 �
ʃkj� �2T��(�U�J 6�,D��dZ�VeT�QTc���Z�A\l�2�AeB���#[����aDŊ(T�J�YP*�,�UEU2�K���EQҪ�"���
���m
Q(ř��V*�m��B�d�X[H�H��
�����EV,%�
�6��kX�Qb��-R0U�RE�R#QF"�bE�����,�DSPeJ��+�*���"�����U$D��Q�	E�2�(�rڅb��X��R
�kP�Q�TUDR,Y1
g���������;��c�짏8`:�����.�d5����A��7б��A���Z4��u$qZθ-J����%�����0�g��RVi �js2DI��bM��O�P�<O�t���8�z���O�*Ԙ�z§P��H?Xz�+<IP>J���tG��>�DB�X��7VL4�!��Γ�>C����b��Vq�����L����ޡ�O>O��2J�UEX�Si���0Ӷe}C��gy�1�!�1x�@ G��럹����[�ѕͅ��7ٴ�����h,��Ld�wY��O���?�q ��J�;�I1
��٭B�j��+7;�M�P�c��J�weOU`,?���?}��}�)���~�'1��<kт!���$�<L{3܁�|����ru�a��x�I�+s�w[�@�bt����<M�VV|��D�Ad�|ɥf$�+5�eB����&{NCW��B� ��9P��
�\����Ϣ��+'m�z���u�'�4���c�~�Ɉ|�����Y7�ĂϘl��7�'��{�@D�|f3���M<@Z�S����T����:�!��D��6��9Ib�����֖㈉ Dx¦Ӻ���A!�8~�j��*�����%|M2b(
I{jaR|�z�����yt��>Iy�ڛa^�H,��LJ�U'{�+x�H�U����N?D�z��p+�'�C�|\`W�Ͻ��*m���1ڤ�|���<NMP�AT���wHq8�$������b��1'�*c�=ՊAa�'��OP*N�S��rm����"DA��(������u�/n(� ��Lx����l� �߹�1�V���J����1�N�hc\I�r��|��?Xu$f�C���B����P�?:C�˴R��>"=��J�;� p�}����G�5&�
�o�O��g�*J���M���xɇ�6�8�;��RcY�����J���d�Sb��Ǻ��4��+�9��~S�����vɶc"3�ך;t:8g�Z�3xmX�H� �����~@Z������
��w�|�?3�bx���ͤC�;��<Ci���B�<IY6w���CW��;�!�q%�jy5dğ!G� �G��)��jي'k+8FF��,��e�w��h2V�m�oX�x�^Rʃ����*s�2�s��l������,��v��a�*�g׺T��eٴu���Zo"҂Tx�멶v�^��f(]��ն)Vj1��˕�åԮ�W,֘��#%��\{'�ߞ�a���C�:�Z�|�� ��S��J�U��*Az������W>���!���'���ϵ��=f!���i�`~�&���`o��K�
�ϟ�b O���𤋮�yu��m��W�;_5������ä������4�ē�>݆$�&�q!�3�9<�c$������d=C�O����x}X>��U�ﾱ_yW�������Oo{�u�J�^���"�I�*/p��'���4�f�6������ǩ1 ��a�i�V��I��:���s�$�%�c'Z�̕��d�|����뻜Vm#Zww\�|�%�0O�����~���B����}��&�M$z�1�Rxg�H"OS��Av��3T�=Ch*a��:�}d���$���a�?!���X�o]ϣ\��������H�8��Gg�Ȧ��J��0�y�H(x����$��g�ԛ��C�?����ΐ73�i�2T��Z���T�=La�
�P�=a��g�_~�69�d_G�R��B>�>����Nb"�
;���3�|�!��ex ���L�p1'�ӝ�d�Af��w!��
�����L+
����b���&?��vM3L�&��O��m�3������<�y�ϵ�����c�j���'Y�9?d!�q򞧩��ϐ̧�I�+��sH%I�9;�Md�����j@Ĭ�>��M��i1 ��"�C䕛�s����i�����o~�;8��+�?'wa�(bL@���iN���+�,O8�7-�I��=�So�
Τ��so̜�4�_�3��3�&3�i1E'���k��""IS�+~�Hؽ��~aMҧ�������R�f��L�����?j�I��ѻ5�&!�w�<a�f�V~�a�i����~-��
CFy��!R|�~��d��X�s��X����������'��Q's��}�d�Y;<�zR
A~�YSl=a\g��h|���=OڼM�|�����x����:�!�4�0��?0�/Y�7�6��T�����q�i����@��"8�&��M<��`z���[���έC�0mi���]C�S�gqל�;̤e�&	�y�+�H�%��淺ve�.1f�jUq���e�Q艺[(Z��Z��]��48d-��b�ڹ�N��)(�>ji���_�'g��l+
��'��ECi*��cw`c+%C�~�j�=f+�XI�/�O�]<`T:���'��Ag�~t��VO�����#������P��yz{����en� ���N�w��@�+�3ǩ1оaY:ʬ�%�p�CI8�z�_�j6�T���Y=k8ú��
z��Ƴ )>B���P�X��AE�Ņ�VNd�g�X�K\F���L��g̗�&3a���a�m��H/R{�1�'P�
��{�v�g�b>s Ă�~�y�m1!�;��C�.���"!���{Z=��=v<��r���`�(x�;C^Z�Ru���:�w01���dՠx��=��|�R�����8�P6{�i�����>v��=C�������Ă͡�s%CQ_P��R|;RWf~�[����8��W�|P�>C�Y3)*8�zj�@�T�M��o�LH.�C�4�P+7�ϐ�
¿���6��T:��|�?0++%w�쁮�?3�;�&�x����me;�9}n�m�x�V�_�`�"��<��q&���?[Ę�O��<��CJ�ĩ<xj�$��7;a��f�M0�?=I�9��:ʬ����M!R|�p���:���!��>�eq��Ǩ���8��*[��"<E����;��m ���;�mX
N!]��ړo�
����tM��SL��̋8�~�blˤ��L����6�_P�V��z� y9�4��_���"R;�S�ߐ�;�S\��UK�u���<H*��0�
���1'�O�|�����p�R��J�����'
���M�I�'{��+%���C䕕�ώ������DTE���� |���]M����=X��4���]0*!����:���'���i�T��hU'YP�<C?O��q�Af��ܜ@�T���&>�b��4��U���O��c�#�!���R���گ9��z�V����$�|�5OSo�
ʓ�$�z��I��L����C�n{�x���1 ���QI󴞡S�� U��Xk�ϐ�A~d��4mD��b	Ǐ^V#�˂�B��;�w�+�9�7�V�k���؊�۩��E*����	e��۸������IT	�Ї�8�d���c���˹ܻ.q��������vfԴ`��g�l�oV��(�C��]J��)��6�=������I�N+&�+x��q^�g����X~Ld���'CT4�HT�&�i�:ɞ����d�4���}�#O�L+�Z���(/9�ཡl�<��z�û�p/��}V�X����-��F(���+�e�(:�:wJt�s��fy�n��}l9zըx�X�řE�1�uL����^V�ƃ�i����>��&����^榑j����'k�< �^X���%\7g�}���#�k�[�#4�ĳ���M�%Y�,��/�ä��7�j�h�K�(* L5t��e�1,PC3*n�M�`{�{C�{�<'ѓ�L�i�u�Vo�S��oT]q�N��\5D��р: ��V��F>���7�΢)xs��U�"�΃9(޷��Rf#��N�y4*�.�_%��Z�^&��(Î@Oa�#���B^�,XV]���j|@y���4j'4�-�ͫ��'����-����/�oF|�-�+�=>X���U��Y� �?���͌��nf���bB����qC�u�)���ī��޶�����a�l���k?��Q���8���z��;
�0q�D�V��+N�e7��
�[��n��@��C�\Y�7��DVWx��x9�Ī_,v�i�G��8�S��MFbv-97T�!ֻ
��E$���N�.������o�3c*�e{u'\/U�:��B�X����n]�q�cr�}�k������#��b���Q�ؙ����D/<8�lэL�����ީ���^��2���&4W��˄�=oh
GP50z�U�ҟ_o��e8�Q�$�Mn����&x;�U|�L�pC��t�^�)W�p.mfT�`n��xu��+aݗ|�ۤ	��k��U�HE3�����(/.�K6ie��zz$W�tظл��}�� �.��?$C*͊�*%*D�a�/*T]F�mn.p`Ύ�V�kS�A�E��%�]�����:sp�
i���KJ��'����ˤ�CC��jq�zt}��L�;�0����`=��"���HϚ���x|UbOѽ��0�z��9��X���\����������%܁��ydW�*�@���S��b�:�w�7���D���h�^���¾T����R�(zP�`[���v1P���&�S��=��w�om'ͪ���u�*�ՏYcd�CX����Hsڠ������cK��a-�y;i�V�>�X8o�y��K�*��t]���s|��=�w[�r�o�;S��=��Oq"����� ��ǄkI N�v\�*��,t�e�YxO�Cn�BJubk:mƥ7.nJ51��f����v�3��_Vx+���Oa�U-�Q�p�5�V��^r�S�U��Wv�	��0� j�l�óۣqg9�bx��'eW$<8���x��6t䥎�̿c��-Xv{��g׈��'�y���@�>�����(_��C��8z�2+��}H�^H��>V�]�u�~���%+�k9��ʩq�#8֞��ڬ
�u�;���w�4F�MQӣ	���8�s�?a$ū������.0t-C^��lV�����.�y�xHQ��yC��ʞ!E�F��\ޭ���p�NĈVb�~o�Z�8Bo�U��=}͍�����:[9�e��3j␡�V=�tz�j�re�~�پ?J��¸n�X�5�(\d�!_\��6�8�,<���^��ɉ�=���wf��h�M��<��=."T�-����R�-�E(گ�n�ޖ}8���o����!4��1���t���u�p�A�<X��R~ي=�A����=VQ��.�U�l��
��5�6�3Q}��rt���\����V�Z�ą�d��#�i4��m��U],�J���\���\�t3��3��C���(;��a0-Y9O�s*�"��}�j$�Hƹ���Ξ�|mtU�M{����>\^(nx9���W�ޥF�Q��;�ѝ\sw�t�G��w�����ظ�kQ��/7J�4/3�G�FcP{9��7:�\@�7d�7�0�gC�pۨA���xV;�&!��tP5����ɬ�S��w�`��
�<K���/⧰ňL�ܺ�<�J��c�M�s�	Cp��W���jL�fҒOD�t����-��Q��܁��ن!��������$�w��A�\�*��<0�k���Z6��mG]���?*~V��<+��!��w2E�=ۊ%Gc�r��P���AUC�&�:(Ē�`4�ok�'��|]�q�,p�ϝ�ϻ�]aȘ�^LZ4�n��K5��p��<(ٸlL!�,,7&���c�<����7�WPᶣ�C�Ŀ��LF�������3�����O��z`��6����F_�T�篻t)ʤ3�tlM�Dc��+.�+힧�x�+��)*��p�*wER�5��Nj��#z@�7�"3�1Tf��H�@��!�� Yr��W�{�%���k��C�۷�g�Rl����9�9^j�lJ����J�g�~@Wa#���ʠ��P;�Z|d{�9�v��,㶳��ٻY7��{�6CA�Ż6�5�la!�dQ���?���x��g����b�m�k�J��̊N�������6��j;�w9��v�#���92���]9��rZvu�0�y§u�fݰj��5�sghҮh����������햬V�����j�������Y_h�z^���(�A�bQ��u��F�ʿgU�'�Sg$t.{��V�	�}��e3��ʔ08U�z+�#����l����J8�{g����M�=���H���HL�ڶ�_KNi���m�_%V���|w9Hz�}i�|�W�5�oޞ���7���Ў�y�Qh�5,��GY�ԺH/M��ja�OFHY ��ObU��]v��TPjbZ6T�Q3#��g���T�y(u���
������.*�99�NS��dI�٭1�T�X �zo�Tb����+�e�
�vJ	'g��M�Fe�4�RZ�U����NP��A�"����L��X��z��m{���g�Y[�u�Rn���w�C��kE�}V�w,A⅀:�o,�ԁ�0�e����rC��Yٚ&n��p�\��/�A1b{�­��p�R���� _��9����Ӱ����egb��d]7�̾��}�+L�ZL�4����5Lb�����>�7��^6�0���ڍE� �N]�;� b��<�O��|0C�����{ŋ��j��|���U󾙴��9�e��mmW
Lw��k����,<�u'��μb��]6��h���yf �8���5&��:�'-Yw��GR�V��Lø��cW�7�}�U}�V�fG�O��]�?=�b�y���W8��:�����NTE=T����lQ�	Nj�v�����C=���̠�h��+u����,+7�V.}��=�u�nn�"6��Շ�k�.k p��r��P��q���M�捜��?���<���q&�7��8U�I:� C�R��ֳծ�D�����?oЛw<{fpa鸢���~~+�V�=�ζ��^�u4zY�1��jvɸ{0��C��Ke������x��X;C��QNm:��;��Si��@8��	��5��#�,�)����8Gq��N��1���8�q��NL���@�N�G�0�g���P���#U|�4�g���1����i}ُ�]ZEu�33��#������;m����
����c�K��c��]���]�b�{��{o�:ŧ\)�F�<���
����6l���H�R�"n0����ħ��)/t�:��ɨ�!�Kt��7��r%	˚�Q�B1Q#�L���pn�A��9��{d��jL�8dY#|�F��ySj+�o����fk�[cU[��/�����޺R���B���.�i��L9���:�ԡژ��7'm�;�ܳ�pn��Z�$=-��-�Of}4,��Xή���Ru�W��}_}�"�5-���4�u|��w\,�&a�Nz�����T[�"����C(t(+��Х�����C�3��q��/�?��������,��.ND��:ἲ+�� 5��ok���f_՛|�p���d��1�~��KӰ��4L*��[�1���Q*zt���6n�l�98�f>'I���r�u�n�s�����wU�B`_t�����,��<OL#L?W0��"�{���b��q]��V��_��F�xX�KTъ̊���{��3RZG��G#����u�K��B:d�gNE�������RՊiѝ�6Ԟ~�Q�H<��]�Yٝf9UC�R���"��0Ts�:b�ɸ���gZRU�?�b���竗��]M��V���P2�U�P-�gKu�������yQ���7�w�m�y��ыgxNdN<���'g���*����k�R|z�Y�a|Es�(~!�N_ty��9�י�+�����ժ�_n��FLPB�g��e�Y�#kU6~z��Ώ�nx�d�3qt�)-���̇UM,f�Ʈv�UǎsS)���6�@m��Z*<���W*mD�!ٶF��zݡ0��A���`U�B[��!a�����K��ӱ�GY.n��#&Db �v�(��}Հ�4��J��sT <�������a˓~2�u�ضh�]�@1ī����6�J�(�4T�x���e�=�ڋe(&�l��K},]�(�0Q܊�_)@fF��mM/d��C��F.�W��V�-��b]{}�֑*� ��=��㘱�e�����v\��׻�"4:���a�M4���umJCXg�������q���K +�㣽.���`j[���4C¤�]�W�.X���԰ER3���ۨ��hd�s/ ���:�x�"�2���;e�d��0���p��E�� ��[y�.r�`V�d(��Ja�ūhtpu)���=��QL��OK�4a��s)d]�w��m�� =a�߶0��i�ܨ�'�.��v;΃/��-`���f�z
�=��gd�90��v����㬼�$S�\N*���P�q�l]��l�!��Ϻ���:-���zN�:��gr�waY/��	�(I�twZ9s���,��C���Λ5ܙZQ�WbF�s��[�2Z���[�xuA��5®p[�{J��4
􃫴s����G$م�����x��ʨ�/�f�t(qc����4���Z���*��xY�ʝˍF-�坝��1�(�+x���U�|�^�6R�S	�j�樂-����ķ�Z�q
������);���:�N5�6�'�j��O�	f���ʹ�wAX�G;��;UC�d������K�)"��]D��y�*[P�?��Z�:ؚ�K�.�5R��\�����Ⱦ�(0��%�D���6�Z��;;nt��ʒYnAX�8�4�ZӅ���<�*�7K:�q����#�^,����}�uϰ&a�@�g󋊕�-�m��2�C�B96g0��:b-mb��si���i����X�p�f�gaU{W��� &�H��ER�uc@�gH���YД5:DvjRm�}c�in7��,���o^@u�-̜McZ��<��{�G��U[��2^`yB��ˍ���:ټ�v_
�O����r7K�%]Xg<R���ZW5��I���6�c��g0q&�_o�#��D�^�[V���H�e�F����w+x�y��_H��o����mY�B��WIz���$�v-�E���X�@��CE�f6{as�nՆ�,PG�a+�ro�T��F�d� ͧm��B���*8��{�mp��K&��B�ޡ�AH�U�I�����Dr��z��.R�g4��f�j�g����h��)u*����[IM-[k�y�Y̵���&�8�I #�omM�q�j� ��x�83��Ƈ��r1t����FG0Ctb�� ɱ���������{D���Zʛ˫T��_���{�7袔j6���X�Q�Tƀ��\lYP�IY&%Qm�
,��X�*UdYP�(
ES-XcQ3(cP����Q)J��"+�`bIPV ���cTb�Q-�P+(�Ŭ��RV�+R,PQjTm+��T�D�dTb��1U`��%F$�R�(�)Y*�`��V,mY
�e@�Ym���*�.!P
��.P�X�A����� �F
(!X�[�ApeEԬ��b֠*��b��AH���R,SR%�ĩ"2*��I�TTE*�aBb��E ����)"�b5&2�`��PTUQ%J1b��Z�"�X�AdY��f!U�!���V�1�k+%V�dQAUS�EeLI0b�H�\d�e����j
*ȵ���,YlUݼѵ)q��@�H��ô�(��y<�Uҫ]���{T�"q�3q�%��q�a�hd��\-��]:����DDD}�v�j��H�����eƼ�OӲ�p��,��k<xJ�����\򧼇^=��˯�u�k�Pw�C�&�`�ҴâåWz�l���t)M�)UvJ_:�s�-��̞7�C�#��{R�1.v�T�Ö�'��p����k�89��$��ySE� �\I����͸�ս̸RQ�_N��>��H�E���S�����o'+��8����0��|��^.j��Oa���[�}���	<�_��o�[�	D·�ۘ�\c��^<�L�ާIh}��j��:tf��11.�Ș���,��?hA�ڐ��z��&�*d+ץEE��n��7ko��V�Ku'�W"���ǯ�K�Mx��[Q#xs~���bjv��r;5��Fg�0�-�js�1`uCw�LR�f�m�iۥvJ��������*ܥ	'�H���e����˞M��"�P��H��Q�`	1E�X�8o����z���2��;�7�C~�W%�# �G;�-��UE��p0O��S ,�f��0�\G�����9��Y�9{\F6���2���������TJ�o��� y��&��~��I�Zu��	�w\]�]�U�^�#�v2w WT|��o��d��[�ˤ;7F��7�i���Ae�1��t*9�	}��� /�a��s��u@��cTL�z���_}��W�Q��7���L�F�鰽���q��2tD^�;�+���,5���Q�o������齾��4��Z&�h	�V�\�?���!�SJV]�V��s��T�R+�.�)Ҹi<5[�g���aT����?\�.1�P����d���hxxj�/���ӱ�)�{z�bB��[./��z�r<k��%�6�AZ�J�K��D���@���4�THsy���{��n5�Zr:���m���E��\;P�$E#�������Z���n�s�|�����:g���qT~�R����f;")�.!+՜7���B͐%R��9NWY}œ7y;}y�W���#�^�}�$/�V�+�i�����b�Li�G�[Κ�'���S�]9`F�o(�$VDOS�x4c�0:�6c~X���ѧ�+P�q�}� �=�x%��x��tO�/q�Pn�C]%�;f��	*�p�S�����s3.���^���,o�EEK�9#j.i��˓
��A��lʓ�:��WˀPs+k�<}+i!:a�,VT�X�����k�����+�=ۨ�7��g=r�;��~�J��{P�k����uij����BM��Ks�W=��>�&Ym���m'��:���K�� gI{y�$�7�Ӌ��Z��+�w�k�E�W39��v�L��h��?���>�脒��m��=Zh{�n��d�+h
�����ʘ���5<H�|&)t�ndq��lk�:©�Q�m��B&F�������� �(��K-� L!ٿ�Q�)���z��y�-dfG�����T��1[Q��%������+�҉Ր3K�0�ڡ<��z�F<�nl��,[���]E�S�׆��xʮ�_δ��w�+9^��x�KCM����e(�[���������5>8�d�Wg�Ec³�[����y5&b7jV����n7��k�o����͚��PP1��Y�\.a�>�|�(�\�}(�5-]�MaR�´�����ӁSܿ�'fldscdہk�oh�u�h�5پ��9F���9;�1��V> R�^��1��n�ECW\(\c�_Trʝ;��F���������''nCR�^|юf���s7�!��N�(h�3-;�ń,o��M�ݢq2�	8Wi��Ʊ������w:�U���P׷��Lt�Yxm9L��w1���i����'R�+��ٱS��:���� �c�|�rbQ�}����e��`Z3���B�X��"N��Y�aWU��f�In^2���김`乷S3��y��'C���.fV�˛�E,���5����Y�n�2f4P�������Dۮ�b����U��}�U�Ij9x��e�*�X�R��g�0Y�8����KG�d��J�`��<�H�o-���P���v�]��yut4�y���ߛ�ve���n ��� '�}��.��X���B�|g���q�{}#_*Jv/�q/N� ^�v��=�_�~H�*���7����+�~'��J���سBE�{�y�.�c��)G�� �_B�� ����B1?�]5]4[[������y{w]g��\|N���_15�P�%T6m�փ��#��H�RCR�l���yu�1�����|�7�8����=<�d@/��Y�M_��P�s8�I�{P��q>��x&�x��꼗��ȝ���æ��R$Bg�E�� ���Ms�~�Ut|��N[��%{���{|�t2��=�l|����&�U���卓Af+���TwU�CP�薈�N�A���uol�hdÍz�3��im�Cl�XHh��T\�Xa���:��q��4㍖¬��a�6�n�Y�'5��ŕb�|	�[�;0����1M�K=I�=\y���b�rS1y$x�������,���J��E��y$w��R��Q����,�Z��c0ҙ���SKGi"z������v�9k���fG�0D�6):qSwh��r�y��9\p�}w�:5����w�|��H՝u�~�������V�Ԑ�Oz�G����A�@
�(�\���p���7�5;������j��Ifv�^�5�<>������^�k��ׇ�1�iP2��X-�gKu�����pՊ�-l�:������a��OY��B��sX^�c�H�~y[���gp�1�g 7N��z�7�c�_bj�y�R�f0CeNM��Lud�+�9��Y���L�{O���j�Y�t�f��Jм]��|lM��'�<~�[:'I0'�g�	V�pD�o�i\��{�W�����˲�8���3X��2�Ү�g��Sp�
Sq*b���)PP.���#�o[,�˞�ӮW�Tkڅq��Q�����k�8\:��.]J+>�@Jh�@#o������~�Ob���֐�<s�9�{]�L{���Id�V'��)R�D�JI���W֓.Z�=�]�=B���̼�3�b�!���d�5�ơ�Cs!�!���~�X��\��L����x���880t,���f��=f4B{���1�5���O�Z�NU+ =�w�=:��j���_A��s� �:�M�"{(�9@�9���Ɨg�G�ߋ��n�C�oI�6S:�q����rs���s.V>�Y��-ߡ0�X֝I���t&2N�ft��Y�=�t�wS�w���b���d��e��	����}�}G�<���9�U�>��U'�@���qۥK�UMx�_S�t������|%�x�t�ڞ�x�W`ZQ8"�i�ѷ����Sw�LR�o�ʪzv�G]�����Z(�����$�$������6�L���+��ň�M��DT1�&�Ӣ�]L�۟���xna��bn�q�=�M��1�l�wn��q���4T9���l��&�O]����^�U����k�������*�<S�>)<5F�[�x�k�#�����O�|�	����+�y��f�MX~ h�k����J�	�h�s� �e�Ef�>r���K�ky?y��*�o�q�|�3_f����g�"�MpwQ;<%�S�}1���-2�����W�n��9�UOd�~�3./s#�A���+�k2�CY��W��/_,;$��u��/y�j|�#^�PCs[��Q�-F<�;!zO�[�z:��'H֍;)?��b�ꎪ�\��٤M1dclc$$j.e�g9U}_iA��3�S�4)��	mH����B�Һ�$Zt� @yc{PNq�v�FD�X�;y��Oy�%�
�MB��u�z\��/8-�.H�u�茭V0�;���
? �
�v���_)�q�MZ�����zKw1Nr��<r��z�N���c;���j�o:��qf�ݱ=�V3����}�}hT>qZ�r$��̀����Ϸ�]C�^v:�'��ڦ�8�?)�x�3_j����;ckG���غ����1���M��*@T\�h��C�7I\�Wq(���mK˙�۳�ӂ1�WJ����yV�CZ[�o�ʼ$��s݋(�^�՗��ڔ� (n��*\�
1��Ɏ�� hKb�Q�4:8J��pk��ES:��w�@�Y�GL1r���΃�ހ��y�@�h�4CS���փ�7FU�-q6[�K'8�ZR�D�v��1�!,TB{V�AyLA���������+�C�' eSCeͬ8��9n����jvNƗ���b��I��N���j�h��򀊁́l��=ra�=�;�\Q~��
�*�-�y�^Z�'Xxy�����W�Y^���VnOP�u0�fS[��	Jƶr��h�
�Lq�c�e���xS�,:�|k��O+Х�d�:�O;9܋���kj�_�m�1|�-��ͪ�u���^E!����y�(� ��H�x�n�p��Q^��9|us��R�d]�̾3J��C��a��nq���n�#���ͥ��}~_b�pf�t+�ߖ����6egL��һ,�����셨�Vu��2���+�-w>���B��cz㕺(fvW��6�o]Jt���Q�3H8|?}_W�}�NR<r��ձ]��)*'���rLCο�Rxk�= � Bu�~7�+���׈��0����7V����1��
�(c;X�4S���%_�����^��x0�MW6��:�-���{Ovh��v��^�:#ʍN�7f�j��<�*1�O'j9���<9�Дk�#�<��#��ұ`�P��]*���k��}��VK/���Wf06����Y/32��_����GNϻ��Q�I��ir��q�<ƪ�h)�rأ�Q�~j�}"�5A���xj���C��L��S�2�s�ۀ*j� ����x�W�����u%��uq�NV���A���9e��a�Wa�*���?$j �P̑C)w>$T�2sث޼�(���U���y��hb�S���4/���dg�ӛ�������G�ЭU�X�M�KU�VJ���gsg�:2��+�Pٿ���VD:��tEB2:H,���-�[��<Gn$�8z���T��0p��\�9��;�	Xk�W���\7��ϥ����=���t=^�4���q���{ǣ�á�d�02���gR�$ęԓ�|�X�q���߷�����5zF{�9��S}Sq���S�͒�#�&��}n��@
0��DGJr���u�U�Q~�������\Z�z߀Z@�W��
� ;M��9�B�p�?;��9`�Z�5�7��*�Ϭ�c�`��g��)��)h�Ч}�|���u^�����LɎfa_}�\��h!��_ή���BT���]��a5��xG��A���,;�+��h	�6�Z=����Wf�Z�aH祵�p;[���'���hB���B�m�qΡ��������-2y��%R�]f�2l�H!!���9�1ia�*���a�vn6�`]9c��0�	��ِ�n@�\�N���|_���{�(�R���kƖ{^�*����U����7f�x?=�u�z(��� �`�����b��DT�̈́n��b��R>��;=-,�F����ʍň�m&{��p`<�w�#0h��W�5�O"�$ze`=�Le�C��J��K�z�R~����������Cl��>��6=~�I�U>�����(�C�q�>n ���J�#��ֈS@�G�C���㷳�w���2X�q����ܱ�j�*=$#P�
Rx�u���"��jm�O,C4�P�T�)J�v���k��n}�)��A.�N��
�z�E׆b�GM#wv�vU��W������㨬d�9�w�k`ᣇ3�o&���<�Jy�^���=5S��u˿u�/[�A��Fr��V��װ�=ԑ ک(���+�ﾪ�腘�l�@��R��h�گ�V��WUGP^ﵫ��ʆ.�EY,��E豔w�)�-n�9?XH�s����j5�����$r5���8�nա��0���|�-�������`�;qS"`��1s5�d�4/�a\N��71�;]t����P��J���d#�4�ȯ�۷E�0a	�BWU��0Ō*{_�}���1�7)֩���7���ʬ[� P�ۘ�Q�ྴ�����;*_Z��M*}��uW��o'���*N�CZWi��qoZ|#?h��ҼgJ�ԑ7Q O1:̦��sX��xf���>�������fM�h��5\0TwY�.8�+�� �)�l�@i�F.�X��q9�_N��B7�zL�������O}�X�t2�ew�wfZ�K1�@�	̰�.�g&'!�Y{��R�W:�y�L~7�T�iȓc��z}k)��OQ���^���������n�:3Q�y����/��l���MA� h���V�+����E�`�:��ڪ9����s�#{Z��L�J�����r�Z�йF�|�wA+�A���vm��ǞgGf�AW��·6]�7V�>b�+�ƀk)d�����t����|)|1�:R�jn�B]mI� ẴP�AK'�X]',�1��ݱ&�r8XE�s�[���SY%k��3��[z��u���$|�Q�ۨof�W���A��.71T�|Cn���WD'3�
�F����w��:�M����f3���۪��N��*\ ��N2��y����4��Z
����7!u�9v��B*���.u���lJK�S/�����Ƀ��5xnGJ]�Z@J������L�m�������>	��U���
��H�"�����7�^�4�h�a*���es�GB�_5���sݬv��({���:�T�l^r���N��/M-�J+P��ۓ�^�����̼�������'XRwٳ6�t�-��6O��o2
4p��0���gn��N�����0������S�v�tu�ޮ��f����7K�h&0�-�PdoNM�M"��J�a��gt	(M$�8*"9Y��e�[����#�Q�����H��n��+��R���ɒ��Ƞ��34���j�KCy\���j�ug,M,�+H��Y4�\�R����+�RԖ���=�q�9k�#Tn)��b���E`�Gۆ�_Ü���l�z4vN���n�gTфb
cAWg��ǘ}q��kF�i����!Ρ��n������L����*u�WYx�l����̇�⸘�{7+[U��B�׸R)f�ƞ8H2t�g�ڴN�F�o����wo��X�)��a�����yɩ��Eɛ����_I9�Y�3"�h�"�V=ܼ�?9�f��W�&vG��+�>?IF����jv���bއ�����${/7�Պ����|�+YcP|v�,Kr?��K �3IYc2V�lHݾ)աh����
���,��C5	*f�O@zx��YJ;��l���Z�G�������5�ib�r�֚V/f�\w��6Ds�͵���p�*���+�۽	����T���5���̫��.�ڳ|C�ܹ�A�m�+��9�RrɫXk}�݀�[4���2`���i�c5¹��w�LxB�9I՞/B��Ĭ��_G��� -t�P�K��#)E��om���n!FQ��ӘK*ʱ�1[ŭ:�����&�Yz�j�oC9*X+�U޽��ۭ���p	oR��`$K����xP�C5Y��6cl�#N�K{*�7%�)}�^��t�N�fZ�IoGY�Xv�lˡeRv`6��QF�m��º�,]��l���t�=lb�	���
˷�c=њ!`���V��,�셩��WN"N�}��:d��^w]M�	�I�>�����U*��-���AAa�*c
��"A��`�
�$E�Ȣ�IP��`������j[eEX��!m�H��V7.(��(,QQQ�3X�)��7.E����*ȫ-+T
�T�
�����b�E �X�E+*-J$PQT���1"報�DXԵ�Pc�b��L�Y"�2(�`
(.0� �	iY�UaU�f2��)A�PA`�ŋ"²�iPFEQH(��H�(�JְF,"V�+�I\H�EV�����h�1���"�
AF0QT��ڨ�DH��*���,PQ-+�*���p��EEcln WW2�11EE"	��z��ն�f�ľ65*����դ4rì�""y���;��D�e�IfWn�"�FUֺJ![�f�5��jC�F\]���}DGJW���󸻪��s��j��w��N���+�W�W�vx_�!�|n�� i�3~���8O�Ǧ���?��hŷ(sY\7����^%i�St����U�̨qncj��;�qn��q�/�@�Q�!������Σ���i��?;4��ˋ�n�5yf�H(׻�RT>�X�*t���SG+�T����ʫ��4�/ND>��vEKT*��	n���N��+�4EQu�1K��Y�����箩|Ϸ�]C�]gc��i��n���g��(�$�0���	n���r��x3<�S��,�ƪ��[q&��]�N.觎��m,�ɷ��)=�N�OX�.z��лR�9n�nz��*0�C��G�5Q����?w|��̓����u�y�[ѓ���ʸ�}�W�3/���������9�s�̪Z�"�BȆ�Y����&!�iY�����GG|ku���`*0����k���,;��]'����U�BWNb⭍���BI�z�{B_cܾ��Xn�I���wC��m����g�.�%���A:�U�7C��
:'�/�[�eu�+�Z�yMԥ���駊��g(9' ����I9�}�Z�di
􉸧%:_=/z�]Z_m�m�&��˘�_*�;v�Bњ"�k.�_mvI�9[}ߪ�������S�WM�CfU��Ëls��)&g�Cl��
��.t��DÚuV���L�jDe���4��1[�j���纊�R��x�#h�
��R:�捑+�믜��:�J]�y�󱔻懫s��Do�*{�޶���(��ڈjr���z��Ñ�Pq]A��+G�ㅹ�����'�}VJ}B�vVӜ�F�8=�K6��-��5쳔q\	�<�_\�y׊�i*�q��\d�(���g>o;��5�5��mqrE��t5a�1�i��(k�of.q՜u�9TiyZ��=�Y�ݭ۞(�O3���G^-�w6i���)�q7"�����qܪk�o*!4֬8�P�+�u�Af�N%Y΢snU��|��($���c��o�m���ǅ����A����m�P�n!7�
o���+o���@J���lWsR�b��`��\�sv�![LM�F�2����Feq(~�؝_v4�jV字�\B��c���Ĺ�yz�E���j�S�p�m���`99�\ݵ�9M��{y�C�h�;��ÌSNw��"쑵)�&�S�y���9pĐ�9*jhG+ATk�-Ư2�YJ��U_UW��Sw��v�wzKKm�tc����,7@�{U���c�<]��$����9���Wt�n�)�[qگc�R�s�%1aE=�m:p�'���G�)�����W�]���n�+[�VpY�UE�!71��nG����V��gV��V���A�]��}w
�����/��w��u@�//3�IV�Auم�qϕ��nzb�C��-����Wy�|r�M�txDx=��q���5��7n
Y�Tk�s/���ʼ�s�U��\ش	�K7���o��]1��򓍛u8}6��&����y�)t�7^��u	�,>Щv�>�s�BWn�t���nq�V)�[���^�ޑ%���#=Eb�^�7��:���S�5b��Kv.!�s��c^F@�A�wU�bS�P���v��~�+�S��֣���Q1������"��jj;C����+!��Ӊp��e���`y*�B�F�\"7F�Qx�;��m^$��놅1��Pg�6�X�N=(��g�kI*N����S������>2�9����gl�Ͱ���q��U2�[���ȸ{�W�_}X�*S:������Q����O�eAڨ��!yulyjo�[�b�wn�2��is�R���0-��u}�� ��J���+���*���m�� ���sr��S�:)�#kWm�z�nS{Jo���ܶ
�#sQ:Ј���Dxx�֌�~��궻iC7�'#JN�V�	���շ�B\�OM��[���"�7S�}���V}�~�:J~}��H�����Ӛn�YIn��[�쉉��l�%Mm(�q�ܚ��>i��]]ں��I�\�{��7����MՂ��"�fH��wˢ��2��&����^��1�ҞԞ��5�4B�������S�M����
�O_�5�+��bV���2�v��du���}M�;Z4Nc��[�q�p�*f��PxVP�t�W-��氼�祖�s�	
��d�
��t�S��>�*㩻��O�DKہt���U�C�e�hނ�;�2�)!��t4s��hw=C��+(�JS����V� J���^'K�r0�ˑ:7�vt|�8��Ģ�Y���q�Z0Vd��O��ci�$,�Huܐdᵷi��3s9ī��sV���8�:�!gi/�>ɘ��uz����֐�L���着���덒�7"P]��#7:j5d�u����CY�8ilݒ��B**cm�������.��x�4�2���]쐞/���z���2���u<�kr�pT�w92��;���;�ڏ�1�^NTb�3��c���>� *�����^���{�>��:k�6k�m��\[�\t����WR������*�Ol�]Wz��39R��>jM�35y��m�^���=�\��,���ө���I���t����l5���TE���>9c�%r�2���Gj
^����qʾ�+57}���q��G;[z��Zؔ�e��\��l�d;�\��p_M���;��稬	��s���OvfL^tҨM����N<Rd�8މt�Bۛ���E>K�Sի��ˌP�r���N�q��%7ʢo\t�m�e���T�mĚ	E�sSq���6"u,U���/2�"�i��ڒ���]�W�sSvD����ס{�YrK��L r<��ދD��jlɡT���q��6Z��r�d��B���Om��&,\�YƬ��g��$�ų�f"9�S^p�۲"��p3,˹
7R����Mq�9���;o6�{1�}�}U�v�˽�݊ uz9�ݸ�q�[��U�a��B�8s����k��A��XN�9��z�.�o4+z2i�1_&ʯ�5P#VU-W�|9���M�ZW�-_����e����TV�z:��Un�¹SC]5A�r*.��tmOr}8�GK��Sˆ��+��e�ɪ��L�q��c�f��{^��a��xx�ܯP��46"������*ܙ���>�����\�ԣs7`�剘�ن�����+��r(�>c+K��It^��dZݹ�}��Va}�*r�\spz��!�
�ˌ�~{�K��=��b�+���_�G�s�+b��Ժ㜇�����KV/5ճ�ˋB�|��i�m�g@�robs�&羜���*�ߛ�����l��g���zϲ�Y�EgT����o���.�<�N���X����Q=k�C}�����YΦiX��׬�m���5XM	j�m��[v����wyA�P���ɚ�.;q� �$��݂��n�8���'�v�:�f��+J���"�E�^���)G�zK֜)�W��;�Ք���c���kђX�h���ygwFn�)�ҹ0s�v�O��UUQ��Z0N�c�[?D����_Y�X��F�����i�N����"cK�Ү��N������	R���nV�QgY|����k��Խ3V�y���nۅkj!�v\'����ßqϓ�K6�?o:���|F9A�U�U�p�[܈ׯ�!���Mެ�c�����͉�1)E�Ń2�6����\�#��,�N�}��j������z2[�㨥b �=�Y�w�%�[ֵV�����B�5���+uQO��m��E޹D'.P
�u��3�S�m�^Rۊϫq���O�������Ekwގn1^ޞ�6�⩍��*E��ȇ��'�Е@�YQ<%k�}w�VTs�_��j�#UX٪��&�5�Y���*�f8�.�K*-��&�݅A=�����p�d�|���&ut�^�ƽ^�?{�����%Q}n]��~~)�N�h�r�fk	r�1aeC\_e)u����lJ�4ڳZZ��ÚŠhN����.d��+�}�]��r�7�h��s��yŠ�P+e�g+�NL��W�[G+�mi�Ws���]?W�_W�b�?7��;*}���\�D9�����݅`Kl���	|pj�ri�hKVÇ�8\�V�m��ݮ�➣��㰬U>�K�����Ju֬�k$*py]E�+�yޚ�5A��T����˗e9�K��$��Ѿ�Ho�v�[��a{t��������,��>���ѽ�OdJJ�st��T�������ͯ5o��O�e�gm�:]K����C��Q\����D������T������iz	��w9�r�b��E�Is�k���d�v�����"����[��r��k�s��Nt9�3��6��my�^�����0tUu:<K��g��R�Ҟ\c�ݐ��BUjn:�m�q*�B݃��]E��OyZ�����N�����|Hz���~�N�W)�s�<�Ӊ`ѯ�T�}��q&��¢�Yx�kqW&����)�'4��Dr���Ձ���+q�Q���vW��TU�l������!��Ԣ������4M���<�b�����-M����	���j��U��	���L��X7�4�����N3�T����Js��:AR�Y��t�Ҙ�љ�ö��}�}TB�/zx�m
���j��qB���E�Bz}<J�E�y��t�U5v�"��歐�^�é��+p�:���5P#�TO	Z� .�}/l�ǵĭ�r-�6�m(T�7q��v"U��u�Y1LWns׹Ue���xM�&�[-��}Ƚ��WW�CV]§�b%S<.&Z�X�GD�=��C%=�Sz:b��ǎu^}�Ejbv!����:�si��ۇ�q7#zM{ŹW�&z�<��o��K��ᔹX���[��\�wcdA� 쾐]u��x�o,�u��W�?y@�2���w�GoSus@���.R��ܹ+����Hm=ʚ��O�ܧ#����ު���Q������L��o:s��YWVڍo__T]��E4�g'{�ETP���(��@a�z���@.Ns�����׫!�犽�6��3^����9��%rQˢG��e`�-�>篵1].�%̜Ch�cXUq���a���5��F��VnژR��g�
ʹ6tw	yՔ��|.DR����+]���� � #x��N�1�'��\�X�fi�;s���è�r�>#:�XLW�š�����R��r�-_�>�"Of�<�'y�^�*곎��:Ҳ�7�p{�#_u4��^�O�+�4��<k��ܮ�뗷�~�C�֪�*����+��)�i�v��q+�up��佲�k������Կ��wR؞��\��(��w��|�~c�T�/lPb����+�ظ�Ƶ��ݍm�u�-���R����1w
�}�Sɭ;�zZ��{.9���ftc��n���*�._�����ϯ$������ĻN�2��{�z��}�����ߩ�5:r�CS#R��M�2A�������Wc^e����UV�aގ�o!T[������pf�T���sݨׄfV����̸��w�t�V�=�]�y$1S��oR�W�YO��3�x�I�]�]�E��+��,{a\��EW&kn�H�MYO7Z�*6��P��vz��٥���ޙ�X�bo�D9��+n��"��=L�sM�zWgf�}*9���Ѥ�bB���B�W6���=��ګUǿ7��V�vT5�
[����ҕ�2��KH߻k�2θfb�5΁��l��mٴl�"��e(a��Iq�c�]7��!P�}ش��2~بY�����T��p���Z �YY�|[j#gU���'.�\e#'�_S�4kj̆�����K('Q:9vS�1����<��#���m�Θ��գ�86/�\��ǵ��r���޹'p*�p��n�v��;�i��x��@�f�q��<17���zkxJ�!w��
u欨�����
�a��-����a��v2z���K�%t���vr�L�ǥ7(�s��E�y�b�V�p�;E�|#/;f��Ʈw:�k��T6)f�ﻍvoG�-|������V�f$���������Q��q�DO'�웖��"[�ڲs8oo��d7@���u�;N}g�eXn�K��a��W�H��2C����8��V�cj����51���N�e�T嗀�6lWS�:�-�L1Տs8����(��,ˆ�P�ݲoD��1�˝ԑ`������|�0t�3�c`o杻�o#T�[��
�6r�A�noX�_g�=˚V�pc������AT�:�:�0����5��L�-!�ge�{s!�*�e	��L��|��shk�ݓk)����oN�d&��j�9¦s��"�Őd��n��j2:�|��$Qj��dZ��V^%ˤ��p#���X�;q�i�)c�pmJab�þm�^M�a�gu��a�dMͭ�rk�rj\�3,�PWE��|/�B��;���q�W]�//+�fM}d7�]�\���i'�\�׳��"�gq|�.���o��}t�T�v�2�7���S�a)��Y��� ��Qf�ۓ�cY�^4���nՂ�Jν�[���S$c�bE9�
7��tW�(�&��IDMwr�.8����� ަ��z^R�܍��g�k��^���K�&Bi�ΐk����żڻ��\0���*l�yi��"ȧ�Dn��K+r`e�V�y����%s��.���7˝ԃk�� �٢�E��J�������'ί��E��6��`���3�n�MU��/wj6W�;�c�,ϛIV�ܚm󡦋�_J�	�A�78�T��0ݛΫ�9W��.K0hM��/2<��
]�&=���0f"�ۇMM�S����ZPh����@Y���U<f*t�k.]�$E11S���E`��Ȏfv�$v�^J-���)��i�\#��R�k��y-���{%9��;9�ᘜ&[�Jd_Qn�Wt�ڤ�4$�D�c��ohP�v�AZ� m��Cw(j�}rtY�}��I�墯eȲ�S������$3��g��[����U�hp{�R����c�n]�N$P��vú$�Q��`Z�
'Ts�'u��Bsf�gF�ک:ܶ��s��g߽��������kE��
"�#iF�jV�EZ��eq�" �##F��E��)H,����"T������2�T�E"��X�Q��I[�J��(�Z�X�(.5��TUQ`�b$X�X,X�AB*�E��,X*��B�XR���U X�V*��ABڌ�(���1`�d�9i1�EQX����!X,+&Z#������\`�[j*��b�� ��G-����""���eee`(�X�a��PD��"�1�E��cX
E�Ua�F�"(}�!��]lӀN��_pB�(�����KJb9�)���s,+f`�sT �qv�9��P�-�a�A
G��X��]���������ѻ���Yh��7�Cz�z�u����/�ν��1U�����H�mB�U��[�*�F(?5\�5HqP���ySM`��n���.+t��A��ًPO�d^]�7�E�ط�<ƾ�s�Ӟ~�^��=���[S�6��T ��{#Y�]n�=A;���V��c��_n��O�a���WٝB�;hI�җaj�����M[f:sys��=�QʣK��د�'�ni��/E�h���ѯm`Z���?W%}ҫ���JS�s�ogR����T�
��M-�� �tr�&�ܦ��5�i�}obUAV����;�4�m�Z���{F�|���D�GK�3��_ѥ<���ݸM�)�Sq��nTд�íU0�=���%%ӳ�.��]pt�/�rK�vw���
:b�^�Ru�<;�4�;_`��V��S�I���/�]1[��}���^9�[���v����}K7rRH�+^�Z�Hi�z���>k������};�B-���[� 3�vi�ʔݪMakO�;�ƽ�<):W<��Y��*�Aʹ��d|.e���jq��x����t���w���:��] YSh<cn��l��}��Y4�5�g{Vvt���]O!��Bo�'���zUB�闚��%�|n��[�8���>�WQQ�J��T�1+^X}�p����*�܇�q7X��V+1��l����+.c �.���K*ؕ�9��C�@�y��3K�rqoWT�9��T�5��<�N�&���Q��y�l5^��-��r��ٚ#=��ŕ&�m>��P�ʛv�-�N_lRֶ�/t�K��y�ģ/�y�vR�gq>=ˋm��e:�e���f�k���R�/���h��O--�(t��+����K���S�.#���ZJ������@���tDW^n�V��U�����h����F:�=��f2v��˅�]r�jJ��F�7���f�o+��\��*��|q*���b
�R��*-hʳ��9�oRA�y��7�������y1|��S�k�rĺ�*�b�z��Q��o6���W��M�L�Y.V�~�w��ʷ���+����c'�d~ۆ��\EϮ0���[j��{�Z�xT�١"���&�43��d�z�a)�ޮ�;*v4�L����o��ֳ[�L��.(5��l#��@�,�ɧx~�����'�jd�9���~�='���{�o��U�y�.Q�T�I#K�ƣe䞥����ח���p�*�:�,�z�v���>�v��:�����H����.��Z��=��1<�%�d��ת�zRY�v��B\șcb\T���P�E���pt.��(7q�mIق�
��b��+qW&��.`�빃y�rឭ銎I��d�SV�W�J�rʓ����as��=�2ev��f�ʷ��+ܩ��\6��x�-ؘ�(��}��"xJ�up���U	X�Â ���g���{Ư����Unī�1G�vم���ǵd]�{͔R�[�H?�Қ�{��w1�ˤ���j�K![�?D�g�o��[�j���v��jZṶ�1r�o��90s�yUCni�1Yp�;�Nv��L���������]�W�.V2�w��'�ϲڣ�`%�c7�����J�:f8�Ϭ;����q8�{1�n�w�8�(��a���e+���O�Uw)IWfxi�4;�'�
>��.l#��=1�l�c�i�G��71U�x(njn������.,n��h�u#z�l�S6��}C��)=ـ�׷��b�~	e�|����ڋ�uy9X���1'���jeI�F���Y7��Ny��8�|��׼�z]���qmP\t�����M���dI�҂�%M����mL�g�_�wS�騌xr���nE�\J�{nl:��7����m�G�.I�^����-��յ?<_w�'B�ս��sh��+Dm;�8����=��TB��}S��쯵7�S��{����!�I�Z�����6utj�lKf���nkUg�Y|�5J�)�֟uO�`�������]�Z�
��3����Y6gW3XhV9Y��Ɩw��>,}��u�>��c.Wf$�n�Y[q�T@j�7�J&���7ymŻ�1���WLtuRu�5�ڒe��jŎ3\�53�����O8��2S�-ŧ$�a_�z.���3zO���V�O���\�EBr�^j����7g�<L����S��}d�%�
ݶ�{�<Ht�u��giû]Jā�;���;��L7��K�e����Ѿ��]W^9x8�n�|hAա�Z�|���.���֦�\��%6�4�]�;�Rt]K�\�;�j38d�;왅����S�gY����<�*�i��)�,���.��	�n��
�o�
�T�	*N�xX�ˮ�[�7�A^��G.��ĭ̸	�B���e�}Nô��]e�m��+Kc�ܮ6�C՜{}~�؆}K��v���ǵ�53G�Gv���8׮�s�el��鸂�j(oM)v�1�K��������`/\XY��慵;/�P=�+��;C��SUŻ�X��K�Su�p�X�S�Z�ꉎ���RS�v�����v���C����t�K�'=��;|�i�CϨ}�m9��5���y���y3F�
ɑ�:Oy�n ��,���v�(}1��z����Q_r���+�0ۼ���oN�[l�q����v����nqU�x��h����d����(�s$������-��~"J䯸�%p�~�TB�=:3�&�^����~T]0�(��j;[(] ��oJ����ι�:���{1p�>{�ם��J�ߞ�f\���e��2MY@��=�&����$l2U�;���M�[� �Ļ�TVһ�Vb�G���i9s��j�(3�Q"��������A)����}_-���X{�nJж��jn7�
{��O뇱*������+U]�W��L���H�Lo84���U�	����o���=����%Q�ԁ5��z��7}^ƫ7��I�]/���ͯu�����͑Y+��u����k{�mTf�nP�,��.����M���jf.p*t�i�63q'&Tl?}HW�j����	����{>��AZ�L��J��Դ6�K$O���{�r�+�����.��U;���Ӛ��*�+�Z��g+n�C�f����+.cB�K*"�?D��2�ף��|q�Z\y�ǜz����֎W��\�;C�*��Q-S<.&_m����<����xq�p0�\}�p��5�ɸ=_"�`4U)7g��ͬ�|M2|৞0���o-�)2�t��g˜��۸]%�|���M*��I�0�/����S�b�J6Ν3.z`���l����ZП	[W�\��*W��»����ul���[�u���a^��;�("��s7����9v��pQLض�I�.��'*��j@,��|Oy�N��ē&�;���k��w���}�Ң�9�X��f��א�to����U-[��Y�c����U�/�kUE ]�����Ջ�W��ߪK9]�ix_����ԝj�ZEH����{�T�gu�ۯ�}}/�c{�fO���<ٜ���Xt�7���&����w=�6�f��ee��*�yt���~����+\K�!5(�Ե�*�H�㊍��Fs���^������z�l����-<=�bS]�ëEƮ��� Q�k{�1�F���{j��o��W(��Os�I�K|��P���Q0��îͼA^��̌���;��mD�J&)�⳦���������s �sʃ���͛j/in���U��Mv¢�a��P��Ԕ�Zj��]1[�Q#��\Ɩ�z��u?�����)Q.ܯ�t@�J���Ր;|�H\:ܚ�Xz&w�n�rj����pV�b��b'�HuC0�@�V�h�VR`��j:[q��LC��Qi-"�ݸ!tv���L�&2*6��N3��m(���a�6����fЂ���.�(n�I�ժ�Fuq���p�G9,.��P|�֣�-3Knv°IQ+���w�_�L�yT����d�[�ǰί�}��z$$�Լ��ߠb̰�n����a[��j0ՠ�a�RD�+�<)���施�+����E�K�{
�;�u	�;��=�*���)��<|�KY�� <z�hw����P؊�:xg�X�VLwe�LmCe�u�ɥ׶P�O`9��BUc
�D�ߋ�>�)q^�+��R�J���YƖx�X���C_5k��b���%����;�����	t��y��9��J2_Y�5RW�k�hd�<U5�ʇ�n2:�+��+@��Ի��&��K����ޭs��׺M�C1x��ܭ�첤�˽Sr�X�˟F�8�=���c�]K����!���yHj���9sW��h'2��tSX��׃v9�%s�N`��^_Kȳ��r��F���{����̕£�/R��g6C�1nz��O:��T�����=���\�z��<0�E�b��k�G��w[�WX�%')�j;��/���2ߪ��6F�i�q�7fSٳ5�c���`��*F!��HP11�9�	�v�����IM,uY}IJ�u�t���H@C���$E����X$�T�e-�Ϫ��[��V�]���V����׋��J��J����9Y���gz���!��FOf=[��������.��oM'Ee�R�P���J7�ASQw�]�A���hoe���:��J�\v�����u�Wa(�We�������!���w�M]��+W4��Э�?K�j�/8�3�����!�{ho2����<���]	��M�_AZ��w���\7 W:��kX *L%3"��b~]	m�y5����	�B��y�ɪ�j���o���3d7���/��9t)�1ǡ-�K*�s]�qcۀ�h��d����IP�/R5_&��W��ݾչ���yiK�����nǖ��Dw@�G�V��������Glޝ��+T�f�mL�΃�F��y�|�F��/aÊV�纴Q�������o*i�Q��k0P�y�2�M]�8��D;h%���EVD'��qF-�>�����>�v�ʄ��xHU�f�Z�7�����E�*>�M���z+:-�^i��}$��r'i>9ա�*\��1ɤ�Xs�\������3��v=^X@XGUn��)�}�9��Sͦ�B��ߋ|P){�m>�^�/���>=�4����y�}�EJ���8�#�I�9yPW��SO����OԳ�����癶י��bS�y	V��4�mN;;�`ݸs�8�r�8�H^ڥ�;j���`�l	��ɝT�h�+T��q������Y_v�=��+\�֬b.m���+t��=�u�G�ѥ�M=����k�o���V�U�7Q.]�M�Mnݺ/Pؕ�Ԭ>}�V����ݴ�mB��cB�oC�(z!�����wv:���V�n%t\S��t�<U�wb����%�mJ��RS��	%��ɣZ��u���&�
\*-s�������n5!�*�"Y6;�w@�D�oh^�{hV��=TuR����jU���O������LbSH������U�Nchu��b��bUʘ����^}<�+^C�.���%�K���]ej��+*a"B�.�k4u��R�����ե�	 ������kKy:�2d�/����[�d�ov�;�P�`��;lr�[�8PY��VA�8*T�T�f</�X�NWwD�0��Ֆ[CC��ز�#k�o(a���)��o[�-9C]��'[�ME�<��p-2��v^�t6��I�i�M��s(M�	��ΩI<���3ݙr[�a������)Oeվ<�XdU{���G�]�ʎG,T�񨞧�����c6��;�-e>��A��o���J�d�8��m�x2s�N��1�V��"%��b�l�wb�
��˭����CkNùlR��'SO���;�˜����qMw͢��VV���E�!S�=K[�X)D#�f=�r
&vS�傕Ǯ�^J�81X���{W(:8;�&H<J�ʮf�93��h	>?@�z�>%�Ĵ8t������v��l�U%�W�;x���9�\*�hw��u�vy*1��dT�a�5,=����]
Ҥ�j�ܾ�b���8�zhn�M�Ԍ�j��v,_ms��UF:�(M]%K�/b-wPB!t#�טt�7�	���֫N
<�����:N��9E@�s7GF�v�Ub!r�{�e�ʗ�K��1CSkd]Vd��a�+ƷmF��/$��	�����u��J�¤�>o,uՎ���'_-7K;]Ċr8EZn��O��)�wM5����ђ��'�+�����Q�v�]	g�
�[�L�ʬ�G;�+��`�%3��{� âbm��0����̜����mu�N
��2��T��w�{���.�6i��6�0� ��2���o�]��֙�II|y�ٟ�};��o7��,�Rқ7x �=�c<�XS%+�k�{r�Vs���Z.P\�9L�yO��$�\�&�^�p��P�Mڣ@LS�K�2��'.����tON*��7CY;�M���p��X�n.���5��7z��kqv�/�/_V��]8��u�n܌Ԣ�K/������s]?*E]�G�-��V�Τ�U�B��y3�u%r�{D���F�i���Os��`��F�]��w7C��q�D�mM`l	��e�!�gH�v��י��6R�X�g+�/:�bvdX� \��F(N�ߥt��Y�?�*��t ɜի2
�Vfv*O3��p�xa�{��T�وn��ap�F���@�`�t����Χ+�ִ0��p�`s��8�s;����1lފ�2PX�Ţ��JU�"�����t݌�L̆*�=�٩	��XkN�S�X����x�bܴ�T+d�LU_D+H;9��}�<�yD�*��-���8�Y��(vĶ��V���9��a��C���M,��ێT��Y[�i�X�3�"�n}f�����P�9�G ��7Q݌���=�Vw7d;���6h,���%�|�<{�8��#�! �C��9´���i����� ��lU-��EQ�(����Ȋ �R�X�*bB�Zʨ��Tej
�el���PY*��H�h����EVe.2�&8�YTX�T1�ȰX����Eb�(�4UH,,E��fZKh�]0���*.eF+���T�TհPQc�QAVЪ�b�,�[�b�JՑU,X�,`i
8�R(,X��!F�c�k,Z¦�EHVQ
�ֈ��Y
T����Jʀ�k5l"*EQEQV
��b���f+F,`�U�*#���M&����(��M`���R�`��ZQ@Qe\���eҲ�ݕ��9K�>�LQ+/�>8�;E=�gv�������`�鏶�j�xi]��Q#����X�,�Ru�W�}w7#zi���_���)+y���;[���� �ʋc��T��L��]�]�k�Ke��o��=�W'.C��	�Q-S<	}��3}ѧ��B�3�v�RǫZ�1������Co:2w쫝v��H�,)^NQ7.j����G������q>=0z��Y�DX��y��ۻ�_�@ߴ��!�/����j�_{��?l~�3R�R���Y�\�.�!�GZ��ߝ�SB��W���}�uy�/�����oeFs�r�F	V�w6-�q4�m���fך���m��YPv�8�m3+J�9���S9�� :���1��Vn4:'���o�1:~Bo%}�ؕ��vr��B���Kռ�N!*곎����Y���ϟ&�=�ٮ�!%��u=dU~�jw!Frڨ�W����n��+�F�U�<�|���v�Ot�P�#sa��V���*R�.�[c��ݎ-���z��Z�G�'����-Zݎ.ؙ�N�챷LU��,'��X���
��Jg�.u��B5�;j9]�[$V����)�����
�Og/�^ix;��gY ��t������r�]J�~��}\Dys�����Gm%����b�R���\d��ת�;+�;EL�]���M9�Saf?��������(jl���
���^.��%ǵ����|�Z�,q��(t��:�r	�q[�:���Z2��꒔e���S��Ҫ�lބ�bqj�☆��	gie�Z�y�4J�C8 �j��w���tVҿ��:ἅQn���粘��~�����1���F�T),�`�/rkݰ����MT�>��w�v��y�z�<1��g)1�L�"�=�T_�������fu��y�w���T��X��<�֧?+��g�a������ð��#|�����^��K�)=K��e4��^L5�+5�WE\CjW̧P��w�sˏO���m^c���ɥ�s�=��w�YnX/�PZ�K�8ﵡ��*j������b���b�w�*�H|Eu���q.Ԉ���r�{�=v0�o���ף�]{/��#�X����7�Ԭ9JQ�0�����՚�E�;# ^�M��Y:0(�YY1�GX� �<��B���i���nA1���V'-�m���.Y�k�k
�W�է���hw���:D�O���t,y.
��S��1V���������OFh��6�q�����̜Ö�n�{֥<��Ҭs�79�oj�F*��eC��{�mW�Gp��@���.]/;�3V�	��6�f�%p�r�3{H^ߏ��Gt�����7��]7u�֒端UA9Gk1��R͂��:����V�c��}�ô����z�{����%�}�Yq������f�k��u���\��hUc����.�t.��7̵T�V�6��Z����q�wͽ�SM��x-�n���'k�����F;S�O�ܩ=�֜�b�x�9��\v�8����r�0�K�fv}����iХYX���q&�N�.wx�kuQO���7���b�u�sy��x����#�#�W��!k��K�����s���~.�E~zC�� S��J���z�O�r�+䡪�C��,}��5W�H�<=<O��bHt�z�%��S�L�b���~�s��≓��gԿ�j�xpT5�y�X��b�Wq�nE�mJɒ�̜��^uO����=g5?0n]#��Ȯ��
�;���Vv�	:u�E�N�7WJ�xũ��c�T��Fͫ5ϡ�UTs~�س��+3��fॐ�F*�1Pzm�YQl:�9�,{�	�J���r�PURU{y�uI��UBnp�L�m8�|��yiK�n/�Ꜽ��D�m�|�y�?bS�E�!��q��+_�P������e���[��igT^=�ՠ�(?o]���8�����vymU���1������X�k�,��(O>�b�]�R��s���ͱ�j�q��7'�y{/���s��� ٯe��qߎ)���]K�O԰���PY�'F�7�k���-o=��:#���V��%p�,���!{j�G �&��ꪬ�ާC-�HT<Ow>�o��O��&�%}Ǳ+��ֿv��*j������sn�ާ��i�)5�>��;)�+|SȞI�OC��d6n��^V���ȟ�k�/�ƫU�<��z����罆q�G7[x�6	�~��<�)�y30P=J�� �z��w>Ӕ))ё��a��`�i��+~o6e�����\hU�:����v�]�ˤ��Gvk�>=��[��T��=mL_E\�z�:�μG��N )k�>W�i#�w��X�N��0�I	~�"Ev��OC{9�𼇷P~�q��{���el�:I�跗���V�\���Yh-�{e�3�m�j`=��$��K�DZ��~��U�O��U0so9'Ћ��Qp�8n2z��Br�^J�G,��	���.������}����ݙ�pq�����TG�L7P���x�V��� A�����r�NGS��;/��|��]�7AQsan(�Kv��o�m��J�z�ٔu�׻p�I\��1�}��	��Rw�/r�Yg��P�K����Y�m�֝�X�5��QU�C��>�*m��<x;ז|�(ZR��W��G{:27�G���F�wS�T��[�B�xtm�Z��Kv�#OuV�*�c�uӑ�Pq]�Uf�1=5�;3�u�:_>��+a�Tg5�)�����MCx2�r�r;*�u�Vk�3޿-�n8�"T�G��ӹ�`�
����p*��,��N����$Q��S�?9G��i�Ut�}ʭIѲ�Ɂ�Sz�Mbص.�:��KJ��]��l�:&�_<4�,9����}E@7�4�{k�嬩e�?�%{����O�(k�����B�]�Я*���FLC�诹c�m���V���rY�gy�.{QK��q�_ �8o<q�����Q1��E=��c^Ya-yjӸ[.q�b�TOh��rb�:����W�n��!�G��{�.E�[u�Ǚ�T҉t]�n&���UyU���ZН�я�v:��(�=Y�7��=��Fkٽ��;/m�������J'�|������1�=R��L�ujE��f9�seN�;��А�3�D/4I[:q�A���י�R�5f��|�椹��c�����)�-�Xa*�*$�V:u�!^�f���Ò�X�wq���U���	Cъ��R�[0�yx�3���[����6�yave����A]F����*�ݍu���ޜ����R݉P3���CW�:m�Qf���k6�w��
��{	�;C�4�vܾĮ.D���Ђ֠�MSA��;lDL<��,�P�j��	ڷ���e����N���<u���9�����K�EK+���̲��\-f�Sn2EBJ;���]�w��I��N�7�:�Y���Dɔ�^l�
����ou-;�c�?;Eek[�l\o�`���ԃ���_T��.�	�N��oJO��_[�X��f~Ŏj5gwT�mLո %�e���N���K/ZNT2�*�j�SqR�l����E�8��2.;L���Κ��<�|��d>��A����aX���%��=���.��3��mfT��_f�ﷰ����N�%\��o&[�o����`س�jº��6Wj��=N��s[ߵA��\>��{nj1���B��T6�k����7�_�z*����7W�|�Ľr�:���76��ۓ�cXS�{q�������z�l����Vq�[�U�eF��]����qN:�h��-*B�v�+�n�c���bU|���Qu�U�V9���o\TJ��uk[9<�*�h���|�숦�L��f׳)���Ŕif�i��K�=�BFT�OF9ݗ=�������=��r�n�u���O|����$�g��qA��Eб
ʺ c���gM����^��htXܔ�Y���[�����M����}�wP��%IOrfY��I�7jl:!�F_�����/me<k=t#�\�-�)l����'_0y$1e3y�f=��Y\��Pnm���÷)UW���z����n��c�a]'�x�K[u>ݧ-���R��aU������Q^��I�	�M_O�V�	�
��p)ͱ�B������)�	d�_F��*L���&�}�q�����[.�t�G�i�9CXmb�3�5�a^�E����C���2�2�'�a]k��9����v��z�;�7�W�F+�1Pzm����خö�U�דo�~���⥮�*>�k��x$�CvVC��&w'�>�+[���s��r�
�".�>��
���38��9�;���5Htڃ��S����빩�4���<qȕq��O=��ߨ�{��cަ�T�����n��|2��s]�:�ϔ��#�c�x�/'6�y���*��<�JcP��)҉U���D}�)��|�ߧ ��Y[T8��M�Խ�Ԯ����s9�<b��K�m�f�'9�pOZ��|b��.�U1��u��L��ը���n�&�̧��e�%ˉ����|�-�GmQtN�%j+�V7�OT�h}jo�=%X�:��t�����ƣ��
���K<I�Ck�0��������y��<_x���w跧R���sys����#O���)�Җé��؊�n!����fu{Ǚ~Bo%}��Į�[^j���:VK��|/\Y|�4����n;{P�Z�w���JG�QLt�����J2���jOtS�Y\�ya���}�	�����R�юל.�$@1�ی��T�Ύ��	Bۚ�)D�sS��)����$7n�0!��+j]�-r�~��v��Yk%��{q&��
��.1t��rN/�0�b��r���!yڟЍ��qn�JeK��rʒbz�uу�PY�&��9����TV��sq|�݈�V�KP�Օá��I���������K2���ys�-�6�&n�T�R�* �%���Ä��㉻��w�����'VMc{�\�wQU�'N�P�ેA�g542���E�g���`j��,��r���u7�(y��oe��V�k~u�x�Q��G+�;Om��zk�X�ƴ���o����9Ԙ�f�����V�Fs|]�FQ���T4�ǘ2�M�me�j�2�1����ɬZ�\Vx�[F�F�������1���V>ۺ�:���"�XC�Vg6hlE:>fqc��q�wQ\)�n']Q����Ӗ�������~�4��U����-)v���V�8�UL�Eғk��|67o�^�|X�;�h�58��U�믜����"�*����ON�D�k���4�#�e�8ն�3�j�I��۱s�l�6�B��|G��ϗR�}�46/<^碥�NRϢ���߽&�ކf��{�Vٯe��<���؃�t]�9ݷ=Noj"�:�Q�����LF��=ކ�*;^�*C)�Hh�<36We�o@X�8ճ�Xf����N,s�}�#^}����b���q~N��J��Vh��e)�k�h��*��h��	��2ru�l��A����v�K��%��ti��Bڈ��J.�%q��jjiU@L�ҁ[Oo��qKf�?��ㇻF5�i��u���0��mɩ��g�� �*�u�(bĽn=�A���M��� ^Ύo��R�(��g�Y��f�H�6tƷ�;�l�Ҳ>oV�*Ư�0v� �It��z���O�T&���$�X�ma��Z%̒]���ӻw(�w��UgTI��-f�CJ�![G����'nK[Nn��(�b�PT�0Vر����	jA���1Ջ����[n��}��E��e���@#Gg���/O1�Ňo�h���q��J�4tE�"�D���zWgU�f�sX�A���aBW+�eC�&�2`ajn����%p���U�5q�u	5��pS��44Q2,TOn�ƩG��,Q2nf
To��<��{�h�WT,}�uX���Gk���ߢ��{�����4��m�&M�]��6���fR�z��vNbӭ�5��a7�G1�B-��ΦNGyxZ�j�;ُ��t��9^�RM�n��D�z��'}��g������[���6�;ω�1�1M�h��cGvwp�x�ƞ���PP�k*k�w<Cg��:�ݬ�0�׀r�L��5� �����Fe�&ځE�H�4�à�Z�t4�mu�y��Ŝ`!���+$n�Z����`s]_m�R�W-��&6ta�];z2�#ϡ�
�G�����tn�@9C�K��׿>�{ǲ����`��n�I��Ê���"vJT�ŲL�oy��g�v-�٫�T�U�#m՘~�� �1\�7��xegk~PfNOd��<�^=[5۫� ��1�y+xJ���"��3:��唝��F�ňo4���]���1�����k�PL�<��	�s-T\�h�����6�V_j���:�̶��un�ˋ�1�5L{uч�����\G����́/�q���P�nb|�!�e�a�u��r>�+�t6# ���Vq"�8�>�Z;6`�ۏ�CW���Qff��S8�2�ܮ����I�"3��yp��2�L���`�Z0HH)��H�m���*PN�@��V�U������Zb��Y�w�#2>��H���U$�*���93a�A�2:[s�vd�Q��ٕz�n
��6�*
���s+"��#�xP�y�����w5��+��,q(vH����1݅�ؙ�,��� s�X�d9�x���{MlaBy���>ep���J�\�K�w%	nY��ձ�q�O�̓l�@R��NYv*]"�]��.9)
r�l�]�]����>�xt�J�/�-����Y�|6��A��1�PKɑH)�cj�8�����l��C��g6;��?���t�CE
�SR(�DعojfM��y���G0ZZ��\�/���uh9��7U�.[��og='�
�6���mӛ�5���J��#1]�=����3^��9�{�[��(��j��<o���m�et��az��c�U�n�u�:W�%�R��>iq�q���F�FR5�!�r�f^�o�,ι�N�Ӡ�a��vS� k�vN<k+L�'goB��N��÷���h��">� �����#QJ�e���U`,�T�13Z�"bڥ����R�D�X�@��PDr֥V��!V:�(儨��TQDH*��CN2��]8�bi%
"�1iPD���%QDQ:�Ԉ���**�IX(��LL�t����2� ���AVmR,�˧i�\t����V�¡��X��QE�QPTRcQJ�WB�ֈ�Z���+Y+LCI+�	�V
�����.f,�D�,���+X
���V�Jj������LFд��X���"��(#j*�ZbJi+Z�$���q"�m��$��m5R_}ܤ���e�[���m�-�u���u:pL8�	�K���<���;d(�xH�&^,�[�Ӧ��F�$.��z59��V�X�RQ�2b�$�+�B_jW1T�>jj�:�qňbgu]�M]���Ek��OF*��	��Bb�z��\"�.��}��+b���꺑mV;�ʺ�����C�*)��mB�5ѯpLR�sS�Z���H�����.���Ɋ`�ܚ�Ov�
�;�i��VօG����]\�*2�ۍJ�)S1Py��YQx�O�,s��S�`��Rߦ��!.���{xK��P�A6�lg�S*n���yQy����Wi1�.�;��s�; X7\ۻZ�}z�m¡=������}���K|c�	��͘J*�s�ӕ��oKy������{�:|R���h���b���jSP�v�f'y9X�l����T=�}��h4$��QW�1���VU��z�Vٯe�x�Q��G�WQ�Lym5Ր��ã���qo۳z-�O�61�$���	+���Wҵ*	u���e*ֆ���4L���L�{x
�EP���p	X�6�	csK�������` 6�.는�~`�X.E�x�����6�!`�\��K�w�[0�P��5ªM�K����C.�ws��L��� =c��+��Y���O��~�%p�r�3{H^ߏ�v��4���SG��un�����kr�Ls�Z���-�T��뉸5�X�W<蹖0�{9&�֜��-妟vC����&�p]P�%R���79�Ϟ�9�;8���	�?u=�(;��^�zi��a���9�|Js�*Y��❕�X�4������w��y2E���L�ͦ_�G���0��+�f���z�Q�����!��wv��O�z���A*����T�RÄ�}��Wۗ�X~)�m�-�MeFI|����e��+2���v�F)f��r ��R��{|KGv?�]��?{��	e^�Mk�V�t���
�z� �3�dT<�tE���b���ʆ��g���UI98c��j����|h����p��y���l�J����y���$��Rgnn���Q�5�I/=���P5�ϖ�j{ǰ2��p�:������yNK���;�ITr�|�A�ܒ�ŭ�xG������N�UJ	*�"X�ǖ/u��i����kUW�f]$��r�AnulSr��n�Xd�c�&�L�5�;׽ٱ_e&dǭ��tF.ა�ŋ�I.��73�WuvGf��j�>����-*�%��_k�j6��SRX��}p���BT�2ϼ=�A�[A�\�nq�^鷗j��i�uK��y_4y
�]�c_��s��?��o����G������Q��|��U٘������މ<r�TQ��v���t�Q�U��K���`���^�1~W�x}}�/y\]:�=�?]�\q���_�BpS~w(�p^��쭸W>W7����P^�pu_�]N{5K�-VW���`{=7����F���\o���H�=���T��f���k��<�u�^���8�F-�}T���S���xy��"��g�ʟOu�9p�˗8
��=F��u�}9�ȶ��(\d���L�dGL�Q�|σ�q�\�>�ի�~ʟ�N�G��i�RRԶN��1��y+�c�ر1ؾ�7s=�_�3����� ��O�ð�N�~����Q�p�c(�����ǧ�:�������g�8J��MG@�n���R�]f�4o�0�I�i^��UN}���aB��N� `����2
ʖ^}�CsK�9dYn�6Z>�P�Gn_���3F<1�k�Y.1Ev��f�R��s�?[���.,n���MR$�̺vߊ��]���Fj1>�i[;k~R�V(� r��҉ޛX�7�_B-�.�w����ِəDLp�SW5�=/�tuv=��Љ�c���-f���o#;}]�T��5�����m�?Pex��uAze�^� 6l�L��S"K�q��W�z�,���{qp&E'�w�6��B�񯯺��K���A����F��dSʧD�<�|͘(=�v��Y�w�Z���)J��2|�y���w ��z��O�_�2���rW�@y���Mz���a��o��i��=���2�^;�܋�"��h���ú6XΈ]W%������=Ӓ� !��4����]E��:��OlMV���@'۬W3)ٺ�m�n�y��=^�U���*2��:��ڄ>A�e�t-����T3�z��1%��W���͏i��v��ٵ�<=�mC��7f�U���cޑ�;�.���z=��/��cQ����{>(ٿ!%��QM�챙���2v�}c�en���kK��3f}�ǲ�C����'S��ݻqW���p���>�P͝�3o�qٱ�u��,U�zw��Ӿ#�q`j�y����@�?W��j��#ݶx�Ǟ��'^͌�/xbh�<Gsfp_�ɭ>�;�q�@�}R=��lK{O��\:�=�;�kv���v�2fe�ԟH݁!)�璸��Qa@��X�x:����R���᭓T�WF.�귪(��U$z��;1�ԱV�Q�a����]m_��W;�xk� ��tH�;eP�������9�W�}�*��?euW��e�[u���y7�_m�v��Dw�ۛ1���.Na+��=���t��dγq�>	�T�:����<��2�6�NoF:ˎ����S�}��C�BBPV�*��S��3}]�FL�L��r9�C�Q��@�Ƿ~��=�~�^�>NS)m��89�LqYR�g��L9`=��`M7p,�9z�cK��~�.:��[�5�TO�{֑�dx�6���ϣ�~�*i��	����"����Ĥ��E+�\���Xt|���t&^F�
��C��m��B�e�i������^��}����>>�h p�ʫ�>��я!y�S)a�.W�g�>
���;��x����Eπe�>˂7��ݑ]��U��n��O�Į6`��LLS�������=�
{��ľ�g��([}oe=�u������]���Sp
��:H
�𘟩�m�?x6�U���<3��{��;0�ѽ��׷O�;�X[Հq�@LG��7 Z���c�6�u���MF���{m�)ߧ�.�go�J�f�y��'f�\?;6o�y�D����5u�^e�x.97>��z�=~��o��;ŝ�7ں-��[�X��Fq�|��rv�8�l"�bgj�R ��M	�|UL%x��c2>\�ٺ�*�i�R�����ϩ��I�����{�x��β\S�U�U���2�_|�(�1h�$��p�w�8�����A�ԧ^[��V�S�q��̥�8��ޅ~�_��LZ=:I_���Ϧ/���{�]����v���^��S�ǿe�b�����ޥ�u��9z}�D�؍R����*�ǆ��w�Gz�鿽�V*���:b��4��sݻ(-�[�[�D�r|�׮U��|%�xeg��V� ����@^���Z������_��7|Mݩ]hl�3��Bo��vN�ՑUDemC�OQ�� k��q����[_4�N��;�mw*B˭ٯ}�H/<�4o������Uhҧ(�����9����	�[���=��ٙ[	�Q���sv�皣�c�ơy���4�ϟPٛ����Eߧ����g�y˓l�^]Y�N|�&<�Wzr9�|]{N?K�H�}��*�ߚۖV}�)�t��4�;�VI���^�^��~?���=����ɔ?^��񖎌�\z����TC�Tz��Y�om) J0���|Ԩ�#�9��"�E�L�+�R�]dm0�s����r��D�ϵ��N�H�
���[�&��%<��'��Wdy��=��T�
��;�-fF�5_]w/��H����=Y^+ֻ�3;��9�͓(�3h3����'D;2�ʾ�]0S���ôm�34��աJ��ǳ�v�"� �?F7����j�1���P�N\pȐ�-Kx���̭�.kB��ړU�z�n��c�t$��'c�;�݂]�P�U����m5�xc�	�Z�KnNH��X�{@��v�E�W���#�TA '�qJhQ}�B��uf��A蠖m]f�KK(��'�zv�8�NO���W�^��Ȩ��N��:,Y���TDӞӮ���g{ۻ���V}�>L�y��/����Iw /z�n��Eʠ=�M����P��Bo{,�I��	^!���u�X��j��y��&3��P��e�C���%��Qv6P������(����쀍�H�BYCd�}:��J�K·�=�"vz<����}�_KQ�J��gy�NK��&|A���Ɓ��p��mzZد����f��`	�~�Iݟ~���M���f���#�M�L	�l����B  �Ee,7���ٵZn4��P���ԜMǣ3:c�F[�΍��Q����R����U����p��<{=TFi:X��ۅ#����[����͛�t��\<.���z#ܬf�Ut/{#��W�����y`������q�w֎�'�@�-�͆����Nb�7��㌏o?_�Q���w�=�޷Q��۔m��-����~x�\�N�]�1�}u��f�sC�*�A��[�Y|֪XwT�k)��3�N�E1"����u�:�_St���&Z�p����-Y{o��U�4�2�^vVw3\��]sn�`��N�y֣<Gi�3r��y�sWG��c�S�shý]��ֺ��b��}k6A(�3���b�~����D���}!Ti��>N|����5��!˩Y��r �~U�Y]�:��;�t�{���������3�D
�Jf�&X^��xX��~��>Ӽ��6U���w�'�ޙ���V_}����W�����D�\	�n��R�]dmCF��mC���w�d	f�.�y�O��B���Ǖ��q��x\L��el�����Ⱥ�[��KG��ܱ�]9�H}�=���=���П����G#ސ�3����Q�t��KZdȁ���ȾG[}�f�����1Wy�^�x=9��+��w���Nq(�y��f���\�*<�|��!��_���m]��ǐ���ZLӕ� �V��Xʎ^�<}*�0����r'Ӑǽ������'�}�9!ض��,~?Q�4w*v���SU�o�s�݂X����2��G��z^�y�л��×���w��{��psY&�$�w��_ѕ�a秤�x}N:�4RVi�Oo���eqʷ귶Q5�[�2-�Ay@y�Q���^�����3v��f׸���j�}�<w�IZiv��$o�^�W�a9M*�]~d׳�t�`��j`f�v� ���T;~��P_�]e���EJ��E��2�o2qtvV��}����F��f�T�B��f�q�+m��E�8������2q�g�%/��;\�֠�k",�7���܌�AVg�a�y��G��u�3���Q�U1�X�!%��QM�챗���xz;��g���Vi|<�Z�c�f�o���K�7Ł+-�y3;��L�{�n*�����J��8����/�N�����%��q�o����ܩ�*����X���h���C����**O��z���v�2}{��^�'�o\����f��lK{O�/�È��tz�{]86*���3���,Ǿ���z�t��Q�5���u�ɟ�Hc{�~�i]J_ML�eg�V6�oZ㞷Lu��{�p�f�	�r�\�nrj,	��\;�2��ɖ���y��1��A�	L�މ��Zӌ������p��d�,�{�;�.��"��4��Y~�vԓTk���>]��SA��}����G;�Ѿ����~����e�Ѧ@l��5���>�_��}��ב��;Z\��}�,*�����{�����x�3^�p��.���=�`Ie?{$v�峑���Bۊ�_L����>
�x>�u�(g����q#���*���N�7u��Q�oO�*?���]Ex+[u���p��.��$ۤ"��<��)�A�6.��.�Z���ָN���:�$��#���p����]� v�r��͕*S5�	��K�c������� �h�R]���P�� *��:9��b������e��;�3>�ѫ�G1��`�{U"bb)�{NA-�ǫ�=���SW�pōp��T�Y�C�Ǟ+5^@�Zj��S����g� =5~������&N���SZ�w"o\��鞾��Y�Gy���:݅� ��`T[�\�q*�g�l1��D:��l��%N'�pv�uo������wK�3�ն{��\W��{"<r����.�χ#�7>^��s�>�V�͚l�����r��|	����UH����0x�ל�,m{�Z<������%��kG�n�~���fgt��妒�s��J�;�}����o���Dm0:��#���\GJ�7����W/�W'���uެ3=��1�&w�����C̟qaf�i�� o���0���/���V���0ԫ'$~���Byn`��y�\(~����m�㟪NS0��FV�<��� k�#����7Tߵ��s�����eW?[
Ӥ4\.�Cl�s�T��9�6��Wp�&w�1�d%����b�Q���\}�co�{��9�~+��q�W�֊��QV�����@����lsɛ�wn�F���tm�A��5�h)�"t!u��8����d %��z�;4�I�r�Z�h�=O�nK��y���o�è���k!�!�D�L�Xn\�>;b�CXt\�K˷��&�H��8���jeh�y�6���2�/K�Z{��u��s:"�C\��>F��4�bm��@�O��[f��i����WثT#E	���֧��Yw�G� ��Ue��Ĝ���v]19�h쵲�����@ֹa�t�ȩ��kl$� =ญ��h(-t�i���4!d0]IoCyGw(�gYP�ۻ�f���&s�V:X�*�X��@`�K�FD(WS�=(���������i���U���ԕb��)ӱ��r�өu�6�h[1�@�8�ƚ���u������p*��j����q	�ڋi��_52���sqZ��`���]�3���`J/n�s�$�t�9WQұ��4�IDE>�o���ms�.w���Ze��|�tt��|�da��@f�gr�,��Ԗ��YQv��ミ ���a��A�1[�=��lL����YQM�������c9���X�!�n�M�;��#i��2J5Y�%�8��z\�|��f���΍m̥]��j�z�`H�CD���k�R�@�puj����qʽF�%�	|��[j���R74 Ai����'߅��z�����	4��]i����ԭ�.��,�/e��ko��9��%	��+r�-��� ���tJ�I�Z�m2u�*.��uඤ�X�#s��1�]	�U�݃��eZ��u8�f��L���XY@|C�_n}swi�RY��q-��{H��1*�:(5W5=���v���Y�����8�]9d�]g����F	+�� u8^�$Ѳ�1cs�F�e�P[��R�o�kAJ��{�s`1�W�p��+�����k�%Z��E�貺'C�Q��°���)��M�.X��.��UX@��LCHesw���5��GfRx�����ۤ�[���"]�1�eY�[֖��X.>�.���ek��v������r�ǎ�G+ZkL��$�jcO���H�f��)�tP�~t�w+�1R�Kkc���9��W*Hj�;V�>r�B��4�v�y�\Z)c<���*������vfPe\,@�HP*���e�3�(�#�� >@�[od��+�C�u��o�}lҹ��4��ޠ�
��ڈX��hG�	��@��0H��;���sw���8h���LXγ�r��ՙv{(����!�e5�Ky]�w�l�v�������bx�Y��{�0���+xJ�vg-K�Z�]���5�	�\�]�!I�.r�u"�ۺ�v�׀��� ���L�VV��n��L�3ӻ����B�ng^��{]�T�6 !>�J�������v�e�O��՚B�H�o��5��sW_���U�PX~���X٤����+E5�(�H��kB������b70�

.�c��,UlP�jV(
9s.Z�k+S,̳ZW(W"�[VZ]!EJ�r�QK�
�-��Lj�Ȯ���eQĊ�P��mF(�(�,Ә���Q%�f\�U��L�*�ۙ&."ʉD+%`Z�h�J�k0tYeB�Ņ��Z�bəb �
c�%L�j�[V6�P�mPQJ�Z�1�9�b2��BҚ�`�Aa��˔�SL���J%B�T*TbV�X6ŕ�Kj�DU�­�72�31��"�F��V"�m��kmQ�XV�*��
�cr��10QG-����Z��,TaXQjX�,����(dyڧ
mr�16���s{�=�-�{��'+BW�>�9My�`V��H[�`� 2�(�V��[{Қ�ۼ�8p�l\��K�ɟ�O�����|�~���g�q����;�ʿwX���=��W���Ff��*ݎ��������"*�ȱy2��5W���-�=]��>Ҟo���РfXݏ�c�i�~=�0o��r�VCrْ+�[ TZ���6�U�|<1���<���lz�O��I��9J3�^�mƏL�s��Al���!��X@h���5W]ł�,vxW��\�u�]��z�� �Y��^������n�\?W���sd��̣ >�YPKGw(f(@��t�2�A��Ӿ��н�\D������U�{����d
�S�+·��T|�r볩�]��#����>+�Gt�>�_rf���������@]�e�V�$\���3Z�W>�/Ҳͼ�{�W�=�GT\�25��o|���'^������󝓰=PPsw��5qø����=��I�>��ǳ麅����|6N3��J�%W%���\\G��OM���� O�o'�E�V�Z�^�����W�وo�����4y
����7ޞki�9W��U�`{��E�ӽ�� �gL�E��L�4��jh�]$��<��`�([�2�W�k����ʞ�z�4��5��N ��	s ���n���5�ʗ"v]@�G���eܽztS�`N�5��+o��2�ų�7�H�HDѹ�^Zj7>(�'NO_�݊��;�O��QGn'j�L5�ZoK��OA�;��d]���+ǳ� �N��Bs�"��^��,��ם{S݅��E�G�ֵgmN�Yu�wo��������}�<�o���ް*:���޸H�y⸫����z ��k�c���_���f�~M���������;��!9��#�|���sʟ��u��\<�m�5�0��hc��y;�%����w�X����L�73�_i�3����u�{+�T���ϽC�26��{չ�4AS�D���.fh��D�L�L���O=O٠�����&�v�_R�b̏.=�z�8�CÊ���#�*���j.�7@W֥x�ͨh����H��-S��+M���O�v�������3ⲥ����|},t�Rݠr���b���y}�~�4��Ƣ��C�~��ǧ�8�;�:*�~��r}q�@l�-��D�NE�\�ŕ=�z<jq`,{Ndl���q/��9ӜJ9�H��#=�E<�z.�g����#
���!
��BH�m�[���y�'u���Y}J�����7QN���Ti��K����{��mI�`/�%j١b5!�k�O�q�;�E\��[Mq�wL�;ʏx���w�V�]�Cfe��i�[6&�����x�a¼���P��2�7��mT7����R&k�����Zwxj;���K�����Np��f���k��]쫞��A�D=� V�h��7Q���1��m�>�%�������~��5t��9�;dz�o���W�d�6�wp7~6���#��\�w��>�p�mS�__})�}�_������^�a�}���~�)�ǽ>����Q��W��6=��v��ϴ�q����>���M��ef��g�Q���e���T���S���z�G�<�f���r��QM�챑ZC�^��fS�n���л����UZv���2u���[�^U>8�.�ɞaW���#ʎ~�{�o��m��G�5�ޥ5�/�.�e�֟a�8��J���Z�"�w����d��fV,���ΘI��Ϗ��fx�����]��M�]�Uxed֖/&w����̏f�S J�^g��܁1 3ᱽ^�}��k���K}Sݯ�K������*f=�q]1y3��>	���nZ& ^�������׻>��}~��Yhh~�(r}B�ܹ���ME�5޸wgxO{�߬.>�'FET�/��5z�y��Hw�>�)�]t}�U����w�H�2�;e�I�;r��%��.��kA��ګ^��tv�Y��9�
3m�v�-n�]o��ۋ&���d��n@�-��l���7c�1�W�5vk�C9isg�=�X��V�
ȥ���R�^�H���_)�����ݟ_����u�ج�TY�����@>��<��೩�,L'�2ډ��*g�ܩ��2;�O���k���s���7�_��,��2f�3��Q�l�ǻ�B�^�����_D�`U�dl��/�C��?[f9�w�����������:Ð���w��ו<�%�q
۪��ex�!��k�Q}\ĺ�=�\���*<H(��ͥ!«��[�	����0���3f
o�LLS����%���ǜ-�_W��Ϧs~w�7}2ې <�x,�
���pڨ��+�p."U��&@zo��E>�������¥؋�]p��~D�z'��q�����
� +��E�Y�W�܃6�͢!myE�9�8&��9�d�2����Zi+5��͛���r]VC�c����.��q�<�j���{��ݳ>Ѿ��Bþ3�/I�ZX�,[�9���:��{�Z=��T�V�P�^ț�u:Ǟe��+��S�{"z�;6p{�tV��s��`gܯ�N��.�3��4�݃ �>ظ�M�]�/oa�do�Mt�2���R�Q�������jؑE^�`Z�(o�R�VB�p�'"�'�7��ӵ�:ˎ���p�ݵ��1K�l���xo��6꽫Xwh���o�AS���t����wsJ�ն�Z�O�*R����Vj"�$�^E�Y�}y�s�p���v_�����C���/6kM�k�7�L	�n�2�s�m�Ǎ{$�^�����U{�Nxo�U1���kE����&�.����+j�z���5�/e@��j�����JY���x��n���z�ǫޮ��m�{M!q�jY��V�*d1���D���kZ/w�x]�|�T��k'��T���N}����{.�u��%�@���`�2��Ɛ���Q^W���2��0<��,'�1ѓ�^9�h;�.��!�_�Gb=��.iTf��,�2�9^ɛy^�ts���쭠eV5=�*�ȱ����W�7��4t8�XTg�M�^���@>�`�eOz*��l�P}'���o*�]D�d
��+��Dm0��Z<�錰-��ۺ��O�=1Q�|��w�+=7A�����HB�z��%��ͨkq�����r��!>̯^�뤏�;H����{=�<Y��2<���ٸ�4+�����,'U���͸����le�p�xL&j#����x��g�z w�{,���N����x�>�%��՚�sz	��u%Y��)q��#�(q��I�R�N�R/��2��V�F3�M�4����Ga�0�vک�sȠ:�݃>��電P��[ֈ���Oq���5]��6�Icf
�t�"{�eg-s�f�F�w�z��Ŵ������׫�}�L{8��~���������j<���Tuk>�����@O��u$?�r|`e�FY=������,ƍM�����i�Z�|{xk��;N�71p��yNK���^��Ys+2<}�ss��a��`�ո~��5��;��T���Q�t���=jh�*9�������6��\��Q��j}��V9����!XG{�k�y^h����6���s�및��*�-���g�im
���7TYfν��7��d�~�[��5��^y_.%��%���R�6-�J�]��*`gZ�;����o�v�п�����\��gFi���0�O��)�:���qx���o�=�ٽ>}7��6���Kg�V��	��q[������;ۂy�]}���{ܲ���tg�&���&w��Bs|g�o�������_��wt�� r�k����Uw����{�mh+*�	��/��n2gȾ$,��y�ב��k(�S���e����>�>꾸܎������ES7�s�UXy2/ҙ��a{#��b�{�d撥����N̽�z�7"��oȔw���MX����=1�&����q��D�ը�.�.9�"4":�GW)V)�����n�U��ּ��ېIz%Z�=���R�JC:��,m��B�S ��Ef�nR�qW*3��݂��Ǔ(�%
.��B^��7��W��j#�����,�.��z��l�`>Ț��4�QjW��[�/�T�s��E�
�2Uz7O�{����Q�'û7����xQRYO��!�(l��6<+b�c6����B�E�F�4j��~����#�����[���W����X=ު�>t���+�B�a6j��xEc�⾴��ϥ����\J7��#K���dk��*��C�~�_V*�t�ϕ=�R"͊VE3�8�È2�z��D���c �)zg�le�[!��J�Y�X�]�7hv��]��>��;��m,�i��:ϴ��TB]yE�\0w�-=�>۷���>*��|��'�����<���9�Uyɺ����a�z�MF��ՋC�j��)����ꮗ�Y�4z>N�h���q�:�>��x���%�Ux.�3c�o7j��~�r(��yq)�^�>���5�	�O2�17w>#!�a#�ٝy����=,��>ͭT�>�f�˵�#���n�z���ٽ)��|X�������S�7�ۊ���}�O{�����o;]����E�w���CX{Y��j�V�)
�TD֞Z�}��0��UƮU�qR�=�[I��k�]sj�f}َ���
2�[��oud睙R���Zд,-�U���,ݾ92� �m�Q�1�F������z3��INwղ��i4�r���:yh�K2oq���4N�� ?���8�	�V����Ug���-^ms�s���r�~d��|�i��.�3��1���3����g�D���T�)eS�t��3�:��H�/�m���G��C�oc�/gͅ��;{�e�Oݦ
�{��9�_T{Mb�b�gY��&|����VN�{.���r�#F{�.ޝ�u�z���ν���P�B�\I�ܙ�>�����?P�`f���ͭ�����e�������w�x�;��psj�
�Y��P�`>��� ��~~5��}d�g�6V;�y`,ʁ�ޗ��������:H�������+��L��e�|*���9y��}�|qr�DUH���dE�G�XJ��;O�ٌ��
�����Ͼ�q37���	N����Gd�Sτψ��h��:�$[TK�ؿ��f�[:S���[s糒O��o�cQgȩ����F����3���Y��ٔLdS�������@�<}$���A��կ<ӣէG�ί� �)�����fA'�P6U��&@zj"�&&��g���-��i��g�1�j��5�ǭ��2�7�via�`I����IsV�K���	Uڹ�=�B�o^B�+���fH��d���t�Z��Ϊi|�M
�cꛪ�ӄuL�Y�d�����vn|�GIde2��u����˾�T����xk|ٿ���@{�� ǽ�D{=�r���u�A�s�t'�Ō6��/�צ����_�I�=�Q����Vj^����<�D���(
�;�Iu�H��{̥7��6�*.%埝���s������m<�lfh~)]�=WU>���I�Q�U1� ���V�<ׄϥ�G~��ӑ���=�=_�a�>��Y��G+�G�5]�{��E�[vZ�(_v焁�r|��b�<�Κ��nK�rR�^�o��	W���{^}w�%�VZ�L����1bm��w�M�mW�z������C���xrvaߧh�y�� ��lب��]R�����mǵX=[�վ���<����4��=�g�>�V�*r(���4��ϳF�~@/Fy�o�&n#�X�����r=��WlG����׏8o���VC��ќ�O���;�s|�p{L��j��2�1y3���N�M�o;��~/�G�_�Z������b�˸n�K�Q�N��*�o���XDdEϑc	Cݪ��q����q��2�>��0]�S<f���<,�cѵeK�8�8��)T!�la[v�'[/*7湼�3WF�9��E\�j� R���됋�Fz�,��u_\��i,�闖�f�p9/�M�G�Ur�T����O��v�u�/�ۇn�uClE	�ع2�*�c�a놏�Ǧl�j���Wdk�vn� �"�E��dEy�(�aW۞�k{��zp�~������9���H�^��ߏc��f��
͊�WҽK��tQ�ҙ�e��v�u��'~\O�$r=��P+��@^f�{L�9�@�R�j�;�.�>�OF(����}�;�c�4��m_�����.=8 }TC��Dg�T<|=4.�_�ꬿz�w1�+��&�^�ρ����%�^5�~W~8}8Ϥ�r�������=���2Q��Q:�^�i�3.��6�1���V��|{���C�s��~��R_������zrfi8n���\�7@V�*�I|WM�=�����~���,b��ܚ>�4�m�*���z�ۅC=�:�y��@yd��f!���/+�B��}�?`���F^M�a��{}�N�!�aVg��]�^�>!�*��v(\;�5��I�s��W�j���󧦵�������|%'������"���}Ԁ�݁}���##ʘ�>�ʡ�`��ӯ�Df��>���~3ST�Y�Rڅ����P*,{:�J����:�V�x�΅`Țƽo%N�Z�}7b=�ٕj��m�&K �9n�(���BŢ#���e�!��$�b�Ҹ��uw]W`Ȑ��+��mzFm� �VdƯ=޽�Ӟ�&�h�7����T�F�Z�u�j�Nt���v�!g8�z�	��b�,'y+X�8��uZ9>@�iuV�5� U=�U4pQ�@	ڬ�\�b�h�/2BI\��#��g�<��qA\����ʚ�epgu}mŌjz(^wS�����'�AN��95IMӠ����]w�Yl����'n*��/��1�Y�vr;N�a�����Ks�Ĉ�`���y�J��{k��e�l�.�O�^�U�*r�L�C���`B�T�nNX$�z+	�3U䇅j�uzx=�������Sj)◫mV���r�6^���RM�
l�'��͝g]c%�Q���J^B�� 1�5�[��������� �ܥ��ʺ�|�m͇��1����&<8HɁ�v�V���[Я�͕c���i�d'�y.��@t��n����r�ő�)��\qsPd���4��I,T�5����uӘ_6��T(��Uvj z�g�gw-6�/1�f�1S%51�3#��_k������X�<����9b�W�n����e�Zඌ	^M��qeB]�� {�]qK�*��(� .]I.I��/_=���r�X�gz����.�"�ζl�M	�ԇ��!U�x�����T	Y�Ս��T�F��YG��T����8�l��E#X�>���/��X���<�i�����7@��YuzO�7���[Tpq�&
����&UpqYSf�����쬙n�gZ�WԴ	p�ɨ.����+'f+OY���n�@ ��4���c�jZ�Фm�����3��c���e�c��9��� ��u�4B6P땧�p�6��X�W2������ĝ�ѩ��Ȣo��l�#�*`�2����Sa8-v�b�Z���Y�mٺ�
�	5՝y�����%NΑ��yZ�:m��T�k��GYH�]��*h�O�3
������j=Z����uA������l����}Ն�����D�.Ve/���ɔ�r5|΅�C�2�3���ou?���aJ�t�m�v����d��w=��D�����U�Wb�.�fF�v��3�ø�GyL:� $i96���IYoVT��V)�zT:�sX":h����&��R�[Ineg^Z�y�t�8je�b��&�����{�\�:&�V�w�r�<:�tc'\��EiJ������~��Jɷ7����b�I9τ�d�xM�����[ʸ,r���;s��yY](<�����N[v� �  ���R#
�(��U�Kj�m�jVڃ�T8��3*ш���EUEeaJV���\nR֣b�1��I�ҙ`��,m��#��q�\k#mUb(�na�A��Z����(+Q-����Ub��%�QLh�j�\�b
���J��e�EƋ�d,ADr�2TL��*e(��Z�.\�ԭ�m��EKaL�X�h�ы-�q,ƒ�T�Kq+�cED���\�b ��VZ�2�jDA-*�mƱ�T(ʍ�F� �c[m�ml*��+ƬrʌAj�[eDeU�R�F��&9kTQQqmUcFX�����U�Ҷ�Vը��j�n`UET1��J��"TX6�0Qs)0Eee-�-�m����m��Ĵ��[+QX*�am�
�fY0E�"�UQFo7Kv�l����ùmn-�;�P!�Sa��B_sw��������.��E����8sun��O��ZR�H����{�v��I^~��v���j�����@��v.�}⫣޸h�&�6����G=������7�4�j�4?^Ϳ�(�������ɝ��된�#ٱ���n=��{����o�z�S�U�5�٘u����/�*Y�{gIl�ζ�3`d\���L�73�^}�!h>g�}7x�Zg;݋�F[�/��v8߽��ʏ�/wER*$�.n*�	��D
��Jg	a{El�x@[��vh��)�=|�FF�%�����n] ���vG�C�!�ޚ��M��N8O$L���
G�E����{��k߁O�'����>s��_��"ee�/~����~�>���<�b��{�O����!��@�2_��چ�}}����>��9�8=�wA�g�^S��V�{x;E���/�z"�D�s�>���}/ƾ��r��x�9ģ~�_x\Nu>>�x���@�Gut�)(�������')�x��>��r 2�z�����ǯ��c�
O��L{0)����Ӏu��A��Mz��Z=�M�=��1��5[F�χt-�*��ڽ]P@
���+g��W}�ǌk˱ZvcMb�M%�W�;�y� ��W�b��b��a}�Pky ����D��uՌ^)���Z���R�����d��Y�"����6g*��7�U���#�Gi��˞�\��Pݝ��CU �@���5�Ó�.�hŊ�"��j�.Ż����({d��bu~9��;S�lW��p}�~6���#�7P��+tü�t����)�s����1"�|��zh��FX�uG���t�s"�x��*<Ĕr�U����8j����^~}��M�7����cX|L��{�;��ߚ��q�'�ǻ�|=��,�y	(�y΁T��}{]o�e,�B�x�~έ�'kgG��g���b�ǳ�g|@��ޣ��ݻqUg�����Xs�1�O�p��e�|8����9�j>��z�o�����Z�|����w�_^TJ�ZO�ߵ�V~�?8�֟ё���G�NYT�a�,nL���@�uH����۵�$W����:�j�^����Q������;�r�_�tSg#�;�����i�WL^L�-W�tGb��_%�'\c�^�K�:����W���:�=����Yhm~��}B�ܹ����Q`Tc�{��5�t��߈��F~F_��/�.��|O�w=(p��^\�/ސ%	��������[�Z�dP�j�Uϓ��l�h�w���I�r<{�}����W��p�F)�z���8L'd�i�bn�OJ�W( h_�/)F[t{9����ސvp�%�6�Ի��3[j�a��u�O;#�z���EM���Ԩes�:�U�t�ؼ�����y;.�|�s��iN[Dn)Ǫn�2\(�S=[y�R���9R.�M���`�M��#e��}U"�]0*�#��aU�_��ف���E�7���O��o�d�a�'j�gå�b�b["6*�"W��^6�g�_O1eg�
B��\�{��J�=:X�ʟ{��w�̂K���x����T���}^�G0\8Tz��4�������O>;�/q�=�\�}>\x�������p*��n&@|j�&)�G}.��}�m�ش����vD	�aI����W�|�v|]`_����H*�2ih��g=�zn]a��^%��/��}n�MF�i����Vj�����@J7�X��x�lYZ0r�z����Yo$�{�cx�M��8=�;�5��fk�,z�,̇�ꏦ.=�*x�ǫ�9��Zw�(c6��N1=������Ie�ȏ�?�x���;��:+N���`.W�ت{<}6�盼��z#޻sӐ��b|�ٍ��w�����<���ŋ�6kM�7�i\�Um����>U���s�d��_�ϼ��_�/���Z/�Ew�T�:�"���}l��n���^\%".�{c�ǻ1�k]�����`���Ҷ0���݇���t�p�+zN�ʳݷ��D�,\��c8��9��s�v��P�J6$�2r�JlzM�Ɂ�*5�ZM�aV���Y���Ϥ���7>��*�g�����~����{z���,m��*^e����0q�.��Z��mL�=�P~�w�6�=��s�2~��{}�y��#��w<��oȘyr�̂����^�T��,���`�{*��T=�&S�������s��������>�d����<]b�f���R3;���(��L� =��T�"�|�2��Ux;�-
hy�m��Z\µ��_^S��HW�}���YR�vDk�vn� �d�ɖ���^.�6�N4�~�w{�Y}��q�b�t����M�0��~��
�5i����=�6�K�>��K��q�O����nT�
�oЪ�븱r�I���/#}`h������>�����@Of�U�h���W�|�^C��< w�g|&=�P��}^�P}������� �nV
��N���io�qf��WO��Z͵�^��2��f����c�ઃ?pڮ���o�g�����.�w���:S�.��nM�YZ�3��7i�*z�h�D�xm稏T\�2*5����WЕ����j`�W���ʁ)���v�R`fc�=Z�6�{���=lj�n���3#����j��������R���;���#��z�`�t��W
��R���l1q�&��`��#�]�E�E�˥�k"��nr
�V��$�}zM��dbv��{ө��un�S��]���x�����̌.��r���?��`;��}%Q��<ja��n��ä�8��=�9�V�熌[�)��d������F��9�>��"�����S�{"z��q��a�m{���"��x����Y�*m`��� Lyڶ3�uG�_��Rz��!z̡�G���.=TQӳ�22�Է��כ�̡�݅�[��7U����� ߖn<"W��FD{��<o�YZ/��׵S݅��4��؊ݞ�j�3�h���H�W�>�z��^.��_c��/���u�mH7�)������z����{���#��*��V}U�gKܙ�Lk!9_q�����7��[�H�ԑ����Y|������w��T<�Ke�N�l���b�ɝf�&|�Ι	o^7�{5"2'.���X�r}|ps�\w��q��Z����n|ag�*��s��Ȫ�'�D
��Je�Y��og�9�S��ڽB��x$z'��Fz�����^��*�ǝ����������]n�U�K����&�����}Y��mC��t��q>���G�^�+*Yznw&(X�5&4�3x���=�P�}ZثPf9�COtN�걗�u��"������u����E��	{4*%Q�W�q�:L ���֠��ަm��y���YF�\�}��Y�݂��q4��Xd���y��zqfJœ+�q��p�3Aa\�L%4���+�@^L�+�-߁��Z>��j7�0�Z�6v �qg�,w޿g��xp�Q0�8Q��O>뮕W�������z*dL>��XZsK�_E�T;�__�r �s�G_���M|6uI��u�,�x�'Ê�s�"�*�-��3(=��LӞ��<V�����Cϖ��h�j�zz�>\�}��<|�ߦv'Ӡ;�3�e]Q��_�u�|Lm5[F�\�w:��cO�������T����z����=�W�·�r"\�������H��#�uo+t�6^Tm1�z�7=\���o��}�+���
��s�>;���s��Ӕ;����W��t�a��]���:S�z50�Y��T��:����ه��x.���xN�{�Z=�Q��+��b��ϯTt��8�6oɲ3	âe_�O�c�0�~ԥ j�b�ǵ��.7΋<��R�5�ٚ����j��]�t�䒴��Cnv�ˌ�Ү2|+M�k����,�� V�Qt��k_�E��{k}��Xǫ�M����E���꓇VESY5���&w�Y�|�Ϯ�r�\��it%¨l����ۮ��.��6ڊ�(��5(l��fN�9��҃f�;�J#�d�����S��op�*P9�~ŧu�t7���E]G\0nw-=V�뵕�K��,�E�M��gR��.=��P��,G��˞K���=<:��v�w��_=�M���;����=��]0��}�3�:������:��x�5쐆�t������߫í�Z2��	�L�Y������Y��g�	j|�������F�ɟ��*�^Ӿ+ǹ���x�����g�;#����P]��W�����r�t�~��_\�9y47��p�F�;�����1J�Ioqk�Q�	��
���YWd3p|��U"�]0+�<��e�Wա����1���'Ǵ��Y��R�������}j��χ��E�ىlق�ۊ�
�ex�9����g�,rL*��/e���9y�w7����Q�{��U�>>���{.�e9�^|���A��R&&)�{I����\�혝���vx����Y�J�Oq��l�y^g�z��dO+�P����������u�Y�+Φd���w��=::;�vz�ļo�#�����΀=j�?]��� `���Qc�I�����m��a�l����>ׂ������zj�P��M���K����.�`�:\�YK��[J��^�鬈[}1�ɒh}��]�Z�N�W����=)Rfdu�q��G��[�j��m�A����C��:S]x�N��S]�F�`�T��W>�w�a+� �_*Q���tᇰ��K�t ��z��۸��j/�����S����=_BY�!'v}02M�O�џ^O{V���>n��\5F�|�Ie��'�����q��ްi�?�c�]�����i�kgӽU�����<�s��g���mX���Θ��{I���;P�'�XQ�5�LvpQQ�4�~`�[�^w�4��͢�{^�Sv����޾�>�l�*�xIzǦ�=6�r-��+q���vo} o�H�͎�`,s�٧����-��H^=�g�Y��� mǺg����|����O�����]ǯ&w�x}3t�s�_��1��{���@C�j|�͒��o�0�V{���U��U�L_z��d�sO��G9�i~/���>�9Cy=�o,�N`�ǚ}�����w���g���\��U`SȊ��,a({��^x��E�!�_�c�R�׽�ߖ��A�Gb;��7��Tz����z�]��@'2EdL�@�W���>�p���f�v*����w)C����팎�J���;޿dz�D��������hp�����/W�2uL%���k4S�4H:�-E�!/y=T]��/r����l'/��{%���*F���C��.�a*�rq�]l���.PT.����[3�-�Թ_^�c�N6�v[�[ԏk��5_)��l���T�;�ok��4�͵E?���)Z����m	΋W+���A<��چ�.���R+����/#}�#��ף=>5r�*�]�^�T;�ɪ��{�����d���t�3,L?��T;�}~����p+ޭ 5�� �ԾS�S�t���hF�zV��*#�5A/���j��{No��ӐK�_w/MǼ�|W�-�I��f�ϦAq[��Q�J�,Yu$\)����q��=Qr�ȯ����/R�p�	�r�ɘ�%�o��k�W��^�w����Ӱ=p�w^�����ɺ��[����=�A�R^��&�Y�z<�t��!��urX����dg�rMy��,�+�	Xo�T�m��vN�6���Y�c��zwmzh�!�`�m ����g:��/�JO_��U	��B���9qꢎ���&O����s��&=��W��fp���zzXae��z��g���#ە"��+C��ʾ������>��ɞ�}:Q1V\NKrc�ٞ�(t8�@��U��Cu�罪VA13�Z� ��]�=�୶ע��n||�H�=���T���Z^���r����m�?g��VnD.�iQ��\��	�/��
�`�`sw.5�dN�o&3'�v�d��:Q
c�V��MsQ�Ế�CD�yVj�G]r��]�^k�U0f�{���S�[W֕ۇ�o�Ǭ�{�ט�����Y����%�U��*Y݂����\\Xy����?ނ!���^<���V�p�t�˜�tEV7=���3���3�_s}bf
U�y7m<���_=s�w>�W��*�q������tU3K�e�UXSȁ>�`W wz���[[,���쎧���~��>ӫޯ�Wh1�Vq����6\�dlϵ��$�q�y�ʳך�=��Qn{���4T^��[.6v�;��	~�_�|{*Q�f�C�ӵ5���~�����'@]9dYN�6Z>ǵ��q�i�ސ�3����1�c�>7XF{|T��Pj��i�<���3�H����ә����w)������ʎ���!���&�R%�As�VG�'�uN��D�����T��s�:2�i��1Rp4�>^�'�o-���Fz'����'�G�U����ϑ�`��(�Gr���m����Ou���tzj�{Eg�W�u\���k����+�!ztX�\P�Ƙ7U^Ed�C���73Eu�y}�������7^�ZV�W^*!+4��:��q�:���^P�$����ߖz~^����`�`�I��v�c�򓂒��*t�E��5K^S�`���yOo&d���PNM�[��4����+�vظ��=o[�Qjք�ׂ�� +�cс���՜8����U֘�tj��t�ň�}�A\�Eޫ��n������f����	I�}o�"5����>�&m��6wAwv�����4l��W�V��c'`��n��]���éo|�r�T�trH��ᝨSU�i[τ�M�m�w&4�Vt�(��z���E�ޣ�������+T�j�R����o71�� ���9��$N��uvQY� )?��B�����B-��ltY�֊�ߜn�:���W:�f�'D�'LuY,�L�)21�5�e�I' ���g��Е�T9uv�K�:�|
���ĵ�	��G_��TC���7$�Y�ձvo+��V�)�ѡ���ʼ���*��*V0�q;�JE����,���s���2�� ��$�+��9}9%[�HqLY�	lV��y����<[] c��gv�g�
�����Q%=���Ė��f�w
I-ʱ���/�.�=�\)U��H�1[�׷�_`ɎEPɫ������]٧��R�X���h`Y�8.�ׇ0D�U+���vЃ��=B���;���c�w�t��q���We؅�l��k;�T�w&)j7�Y!���Z��sw�V2�$�bU32u��"jsM���W5�8',#�Rء[�l�N=�Q�4i�VS�s:4�X���l���Tfs��z�3u�a��T�W��ww1F���Մ<4i9QUJ���B�+.T�Ț����H�%�t��m�]�ZX�T�%[��[iކݢ��/�����c�`�� ���hUnG��P���[��`�ttkWQM�}n���3_��<��08��*!5R������)��$�s0�s��ʮ��55d:�Z��VN�W��f��K��Mg[nu���A1H�!���	��.-uƒ�9�K�E>?wQ�Ō�'� �V�M���32e�:���Z���[����{q�W*KuB�?����Ǐ#15X,bOpa��U8��w)�a�P=�B8���
l[f�aI���t�ˡ�������1n�bijU۽ź�ԛI������S��0�rN)]hs�O5>��j��&#�)G��7�Z�H��"O;V�#\�r����\�۝���;���kl���ca;�좮՝rd߳T���o�j�4���7��n���u2[ޥbV�� �m��XwHV
�Á?�mGZD���h6�B	��:��lu�t���'&��5F�,�|��˧��� �7��r�:�$�\j"�eK�v��1�2�����ֵd��R��n�Z�V�;[���\qp����v̹�w6���^t��+��hU��Z�RyI8+���T���yئ�u��r�������_ł2�x����3@٭n) 
v�%ef�+<�0��e)̵h�� B�����T�A+Y%D���Y[m�b�pb������e,b�6�b�J��X�YAEV�EA*�EUm��V#)DZ�J��AAb[DJR�b��bV��(m����ʖ"%m���E[J�"�TED���j�eeUD���ܷ[b"Jڶ�TUUDm\j"��[s0�b���lPb�"�Te�L�eV(���`���QQ�Kj�U��#U[e���32[*�ł�ĖՊ��*�b�J�(1�5�X�[����Km,�����J�(֢1ġ����E���J�U�"���1X��hTe�V)E����m�-T+
Z�k
 �b��V1�*E���b�
%e�A�J���ְ�B�EeETQkX�UKJ�\��,�Ȃ������*�[
(��bʑQ�lm*#��QQVȋs��e*����(�U��R�˂�`���J�Tm��E"��P�[b� ˘b�Y��t�V�xtd�cv~�jt�o;����jT ���U���9t&ؐ��u�_{k��QmZ��ٻ�5N�x2�*�>����ˇ��a�0S{\i=�<=��mC��w<6!:��/eF�^����_�k�&�����L�|�c��E�9iX�1b�_��8������>R��G�9������ˏ.�_�BU!x�����U��7rON��	Cnv���&���'´���o��[Z�ߺ6x�1C۷��F��=�v��ޕ���Tm�˰�D���I��5���&w�W������k���j�F���$,�{m )b�i�߫�\{�hvG{nQ��zi����&*���,�1[O+0x���o�;�WU�`��g����O��7_��}�u�{oް:߶���
�}�-J���Q�j���z����:{N��a�ʗy&W�� g�T��9�C�.��7ҼR�W����� �~��Տo�2���'�/�5@W����dP����寶h4o�^WqΤ���G����;Eu��b����Ǫm����z�� '�ET���L
��#��a_N��jgmI��ty��Y)Nt�Ϲ���z����H�__��<�{+�X϶b[6`���B����+�.��s<��'j�;�cl+U9]9�XZ�@,הF��4�ީ3���	�iJ�����v<�sr�dz��]��C�����m%[&��wY�����Cl���՜7�\��e�Q���/���"b��]�A�n��5��a��U����x�m͆򍲅I��3��Ie�W��rզX�l����$7y��0*3P���3p`�{uH�׹�q�*\iؿTt,��g����O���>���/+�����@y�#^W��!���r59���?'>��{���Z�h����	����~U~9��;�L�{ʀ�cc$��Y=��_���ldפJ�;�͆6�6���vN�z}F�����Y�|�F���q�Y>WZǤ{�M�� ��%z����<���Y5��Mφ���fׄ�cL�<�K3!�ƃ��Z�A1�y]}�8��;1��*x�����Q�;�%��#�O�Ȟ�ï���:'3��L��y�8�^
�7����9�Ѿ���ݵb��l鋏 '���B;q;P��+�X�_"�_rG���YY�eSZM��]-�5�RVU���_���{��(o��<�W�NU�0�Y]aoV����1z��A��&��]gYuH����]�����(�p~W\���C���jQ�[ލ�vr6���e{j�i��>X���3�����X�^����~+�=��<�8���X�~��CH�
p]WE^��*�`���ӹ����n��V�!�`@�[�Bc2nZ�3��]Д9 ��\Ĵ,�����cXܧ�7:Dʵ���Mc���%wm*�)�%9VI��R�Y���M�-lfA CY��dD/���٣SN�����R��wr�f�bs�=���g���9��X�z��d�s3����4�K�q��u�}B`yM����8����蔪2�knYy����n:�́�SȊ��"����jv:�i�wso�sYW�����}�O���Tz̳�\S�p|��$V}2� e+gaVAWW��^�n�C/��n���V����>��;����dxa�j=q�%�d�C�/�T����s����!�{� ���6�����}/ԑ��P-���4W��w"߫�p�������ܕ��7��}��f릅Du<8KGw��I+�Z�IQ�<
��^��~���)�=;�\E�ǔ�=�4�IC,q���'�s�v�� ;+�^5���ߍ��=X�ެ�����4j�l���'�@�}�e�Qn��ARGMK~�=땦F������+�7�#}��'1v��՟Ez!s�Y1�ޡ=6ˁ����`[���F���50�Fm�w�O�I���;k�3P�@��kv�4�/ ���	��(z9���Ǽ�OM����A��7��<zc۵�#x��ٿ�s<��Csp,ZEk�g�V;y��w���^�^��wΑ���`b&x}lCP�I�/�KT��y����[������ʖ� X���4�ƻ<n�	����`���,[��iu�[���H]�7�������s�SUz�YevꒇVWt�!�4��
+�5���:�6�R�_�Ds�>"��+tV}�U	��^�4x�y���zl��ѻ�)m߯;�T�,�3+�m&򼸔;��g뻛�eܧ=]�3ʘ�7�ۡQ>ѺuH���E�i*��ٿ;�?�U{0Z�8z��gmD<�{K}7S��@�n��S�����{g��9=������/**��3�����*�T�fp����Lk!9\d{R��4�y7U���ˌ�,u�3~�|�s=�b=��o�{�g{nQ�{:Ke�N�� ��{ŋɝd��C�[`h�������=��G��B�=M��#����uj�i���r�%l�D�E��U�V?NuPbj�n����U�dB�l��3��찣���gѾ�����\�pA�X]�d{�=s��Ίfs��Ԕ����\	���L�[PѨ�mC�]$r5�^	t���g�����^�mW�K�=�kv�:�6��,t�"��n�7-n�4W��P�_�#��y���!MH訪x����A�c���B��T輍2d@L��Ș.}�� ���l��s^���k9]QO�T���p)�tUj����Y�ACNJ��X8�IN��ZZc/�^c����1B�\,l����[���]xv��ܽ$gX�6�hw�އV$�Rn�{���5í����8��W@g��k�>:;]_��Xbx�ay��6�4���;67������
�B��q�m֊��N���O���T�5Y�~hx�G�ܽ�-4W����8_�w}8}�~�
�s����+ޙ>6�{2S���*TKGr&��ex�̧���'�q��^ui��O<���mY����#�ߓ�_���.pX���^4���<�B�oNm�.g�q�����߽KL+��]&���>���d�	̟q��]P�+(�W>�ت-�y�Zż�bǃ�y�[j�����kڏ�F>`5��'�~�T��t�:M�{�:ʳ���U٘������ J7ު!i��c.#Ӂ�ו\n4����[��Tc$W�מ�>��9�k���|@���xެ����Λ�Oi��	CN���ZV	ú�o�X���z�0�璴JU��Ԯ�����;�$o�,W~��/�=�}$���Led֖@�kQѳ|x�:��F�ٜY�X|�@�t�� �ίi���!���ϹQF-�-���T��u)U�.8w��Ezsk��K>���/&w��g�{:�1��?_�������W�9�C����o��E�@�7�N���=���eJ1�yp�
�U�{*aYϟ�Uw�ove�s;���1RXݜ�gP8��v��{�\��S�ZW��o��Cn=ث8U� d�د�A�� ���D���+-d<����T��oV����l�>����	�.M�����G�Ͼ����r&�����q�3ѓ,/�On&��Nx��~�8>�oFB�sK{3�36�,��P�CUl�r�s\s�p
n�e��/#f�G��qt��y�Y+&�Y��^�Hdl�]��o���ȭ.i�������@l��΀}�R.����#썖�#�;H>;^�|{V��oyy{=�Z�e��5�_�Yr|,�H��̐�^*�`HˌW�ǲ=]� ��Y�Q~�c�}\ĺ�=�\��t���ِC�sP� �`���������WV���3��1��= /d�5=����g����^�ր�<���{.f�f/@������{6Uo��x5;��Bbk�[F�O�{����t?*���@{��� 
i�{��rkf����)�s&|�4�_ORr ͏�͢}~��_F���o�_�P�u��l�~�쀣�<if�(��>��w����O���躯G"&��sg������ɭ,x�>�C�P��<r�%"��{�ꋘ���*x�G�U���Tٸ��,�9���=���u�<�Z��[țU��O��fE�_]07!��8��� ��2H.u�X���f��P�9�Y8�o巎��oZ-��J�K|�^�fuҵI�xw$�5j)]}����}���f۔�*�7u�Sz�;��k��M��q����Ok���t�ԝp�nKu;E�Y�F���Ys����J.W�j�\{�gL?0%iQ'��v���xU�R�z%݄�L�C3�OCsZn#} k������.9{��g��\:��~.7�kE����>��>�ד���~��f��Q�k+j=q����5�GT���`T%���W���'�ݡSUz��ȯ�__��ɻ��~��=�
�F�9�6�]ü��N@L��6�����_�o��/�ľ�N��%�ݻ���D��bξ�ڔS�Z�U���*�	��\;ɔ�/'Լs�sA�zB�Rm:�[����[�t_Z�^�>^��G}���v�6�r��H˕ -���<����,l��7/:�2�<�Z���=�W�/|�փ�|����{��6��q�ϊ��uƸ�f��P��E��;�惆}�9���.�O�=�>g՟m0��Z<-{����J�پ�6�=��G�AY�y�Cr�o��yQۯ�������碪F��Β��dF�5Qj�,�l����������Z��9��'E��Hb���䏪�ӣ=>�����Ā��t��}>���w`��[�����zr�M���0�]uTxل\��l��ёږ� �͝�˺M�tm۽�Ӎ���X9�T����湪�D�aP�;��^��'H�],��i
w-�Bo "6$�F������f�l�ݝ���I�e8�ހx�)p�SV���o��ZF^�]x�� ��ȮʧD\Ct<X������=�p�r	xs��G�.��W�E��{;��o���3�5&��@U���}n��Eĺ��t�礏t\�����P�G=�r[ޘg�v/|��w�����[��9.v�;�y׉Xr�?p��;^ekcĕ�~�?��jp�(xp{~B���A��k��J�O��Nǲ3�s������鶬�&<�����O��+�XŇY���/_u-��F����
�k�n9�5�����9̟����ǽT$W��i	��W���mwyY^<x�j����
���Ou�ǿ	���]��3���;�/�_�"���c��Dm����QxW'��븀av`��y�Ek5Ɨ�Vt03��}k���-gxA�mzr��ww�de~�z�C��F���qW�nx�7�F鿿<x]7����V�~U>�!�Z�4s^�W��U��9v�����Y�j=�k����(�=�D�NL�wŎ{���}��Kұv�zh�B[L��_i�φ|����������+�~ʟ���*���s��q۵P�������^�w���ۻ�D��:����e"�]��bR���#�݀�j�G9��ʔ��V��Y��F��>�_.�N!�]/�ޱP�R]��ч!eK"��k�3)ޘ���.rz�7�ӈ���2��G�Z5��mլ�*�"��vsQ����|���^�*����ς�K������doz+ȭ��xuʤ�x}q�ƓO���AK�N/3b���ޟ��1P2)z���J�u�mCF��P��]$s\O�v�����&4I�^������9�=���,��2<����"�[���F�4o�a�K��C��{i�l���*�m��'E�u��zg�]�7gd�p\���ai̍��^־^�03:}�y�u4w�&w�^�S��}9ģ��.��d<�t@���"7�VE3�8
�/a��=�fr������*9��{��<�&Uzb��R���{ِk�ں����n��T+�����݆c9�g�1玝����Xʄ��m���y��J�\������m�5�ߥ>�#�r?���g孊��:4�>����E|��b㚻��<����s���:>ʓ5���s=T����!�}���P�~`�&��~OA/�����'�~Lψ�7�y����炭���v`y���g�rh�愔s�$,'ޜ�ON�~=&����ؚ���&��z�Q�|]"�,�$��*ʓ��{�*��﮵��1��0PmT8vl��]�f:v���\�[wZf�Π��β���wB�\1�od������֣��Gb!\W#ks�Fq�OC�_7���zm�.٧K"�s#s��|��S�A�WyÎ�o����Q5�+:o�I=��BP۝�2�ʭ����\�V��B��?���N�Q>�?Zx�]�{�����z���A���y�S���]�>�Ië"�����LX�Y��q���}K��ã��S7��7��T�m��l �O���:7���o��Z�^=4�O+v�d� �to��*�u$�v�S1�}����ɝ񸌙�O�,�����S���Sp��,�{"�����x�u��ҳG�/��+�|l7=5�]뇀��[��;�k��i����43]j�>��;Z��9ԏh����eO�g��N��0NQ�)���s���������O�$Œ�geo�_���3�q�ӑ^�4��~=�(�#L�ٸ��@>ʩQ.�,y=�W���hs�y
�:����q�z�1�ޅ\�o�i�S�t=>��ىlك����o��{F��[�rs�j�L����Fς����;^,k��>��.���5���ﾾ��,)�S�(���^�v갘�]ON�݃c�t�Q�K���|������Z+���$�� �!$��BI��BK �!$� �$��BI�0BO�BI��BO��B����� B�} �!$�BNBO� HO�d�@� �$�����@!I?�!	'�B�y �!$���e5���P �=�!�?���}������}�H��UHUJ����%J�**�wT
��J�Q"� I$����*J"��)T�(T�)
*T�F�{���h5�i6�d�6mhk6VPM�)� ΋��%�8  �  	��%V#*RS[ �ue
����F�-�1`P���(.:�q���Q9gwQ�'6����uS��]ۊ(�K��p��jsd��D��8S��);����uk�ͤ�r�v�2+bQ%(`t��٘iF�J�	k6iV���IB��t���EP٢��kd�؍(�AW ��K"ƫB��e[b6j�"�5�)�`�l�Qi���X��f�m HP��v�j�U�i(6�V*�h���m���@ �JD@F&F `��E<`���@4d�i�bdLs �	������`���`E?�J`L  4`�L�4hLFD��Rx�OQ�a46�R	4�T�4`2yL�4�6͹�۸����V�:�[j�
J���@6����Q�AAB�|�@P��:�g��c�?9?k� �C��j� ��`�UP4�4H�b�P-ǥ�ΚԹ���e�
��jJ�:��������`�e��/���>_���1�f��[�r��uy�*E;YA,L�k.Z[��r@#[
��Z����� ��0Xx^׮S� v�U�c @1�[�`Q[�� ��%ʋ,T�ܴ�I���D"j��ǈB�eЀ�j���0Ӓ�@ԥs%�-���RLCp����"�̳xt!���[�`J ��T�Y��1d30b�[�F�N�:�mɛ���fh�H�hm���[�]��67p(⬼���5�l�a�t�v+nI�M�wG5�Ռᖦ"kRf�=�t�3x��÷�o ݒ]���k]�5���U6M��fJ�EQu�cmXl�#EU�
�*����
ү ��e��B��m�H�t��%�ٺۻ�3j^'yQ�Z��xA*شԧ[O4�4�����2�AP�5�Q�ՉڧH�ܚk��u.��h��I���Ɣ�6ң��u�n#�7��ѧ��j(Z�vB��ֺ�oJ�4����pn�4v �*ݽmU�������zU�Ǣ����e�J��8�bkV����{J�8Ct�"qj'6�A�D���gؕb�E։��j�y��U�Dϲ"  n���a�m[ta{�ު1-�S�)K6���i0l�"�W���9��]�l@�m�:�A�Q�nP�Z"��i5���mn	n�حsHy��nZQ ����)�K �2�m�)�j�q�b��7�1�=e�ݷ*�)���ږ˫�skrU��.��'p֬�km���ҵ4ᳯi��b�pY
��YJ�;��X����E+�ZKL��j�{��S����IQ2ܹ1:���d=���5j/3CY����Rf�\���M�R����EQ�̺��$�Le�rWy�8�:��X�U�5��ʳd��H�=n�47$F�Mn�KMe[w��n���[����f��q+FD+Bv�#�/.`��Z�/V���ЮHHa�%Re�����A$� jjj��Bai�(:n[�r6��̔��i$�ܫ��l!cyؕ��CT��f�m]%�0�u����77�KMw���2��b�mn6/e�Ŷ-l"��z�V�����4�s"(�i@�Vn�cu�";zR5yE[Mr���M�/d����-�R_�V��ݭ(�e��e��)��1��.� 13u�Zș�&Ѳ�#����M�k/0Z�N�0�tA�[RT�8v��;);+,ۻ �m�pe`X7*8l; Z�,���{�]��x̚E@��T���Y�́����0�F�uj�jŒ�4�E�F<g1){��-ÖB�xh��A׹�E=��+M݂-XM����DƁ�9u��F5���Y��v�#M�e�v��`�)\+s%JJ����E�郧4"t�i���˳��^�ڤeo�V·b��-%��j�>�ih�&#�T$zFV[e����T�C�)P�:	b�K�U�ae�%i�]n��PT~P�)T�n�ؒ��k�F@���h��E�𼘐���0��vY��*A(m�Bh+�ƚ�i@!kw2�2LQ�NSa;EP�/n���N�f�2��6�/S�9x@"��kZݳ�-�f'A��
77t����k���Т���$ �S0�z�16��4B�]*��ͱ[Z�ˀ�-��
���ԇ�WB�70��Xr�Q��G��ʻc�f!fTy��� �I�dq,���kDG�b�I�Z�P�A�ILD:�V�쬎dkj�]���@�@tn��yO4��7%eȀuZ%6������8ĩ�����l�!�Al���:nŜ���2��3�m1�j4m��P�L�����h�9HƆXz#�+"X�,V\׆�oUӤ]m�� ��l����6��ֱ-�񶮌[�m^)X�'��W1KJ#�̱6j,�CpVR+�B����ř�fJ�%bc2��`�����D��f�jL�'�M3I�ۺf�ee��c�a6.�H�T/_| M��cnjt
�[`
��'[�w+v+bN�dUCz	��"�'[ pf��[�J�
͜,,L���˨�KP��t��+um(5�9� mʚ��#��2)XDH^���t33%(�����^��ѤGE��K��"ޠ��2a�c�H=/��X�ۄ$2��Yv]�7	���h�	�k[B�27��r�jCf`���1�#��o�� `�dF7�@��&�E���5$����͟�:��QK龋Y�c�k�W�*:7��� �(�֊cU;��x�C]����ֽj[��zM��"��t��YyQ�ƓD�[�K�(���=x�@VsT�����` B(N�-�S���Qa��*�E�M�}X7�d,�[(��I� �;x�*��{�f��ǝ�F�i���KfP����'��Y��M�����fX����a��\B��氫W�<�t	�-�p�MF��4P�w��6���]�N�\ov�K�ΩK��A�)+�f��&`#x��,����_V�6��谷(�6�1�u��|gDU[��XK9����\�uu^�5n��WS��i�G��h*�z4�9�'���}���J��r�[�̆�+�`ue�C�ẜ�y�i&��u�\���:�nإP��=.�#&bJ�7+��<MU����]y[��;����n%��@!�ڭm��n�>w�ݠ�[�-���x��G_s�8�����8��Eqꉴ�'yC�̥}Vt��r���R�1�}g)�4��3�;S��]�p��n�Z܋U(�2<7�,�V��՚;�@��(%�2A܇@������V-^��H8оJ�N�^uv����U�UeN�fFE�f��5���O|�ؔ&\�wj;��γ�{���3�X8��_>Z;��v�շ��]����8CH=�`���c2�L�яw����U;��D��7)�§	��}L| :��t����U�VX���(���7f��|-��]u���~�L=��{M����&�G;ht��/Gu���݊�g���7[��2�m$:���ws�K��e@���b�����O�n�PؓZs�o=���p�J󃨊�� ״c�r-�6�r�c��X
� �B��������Ap������\�l��Ϲ��y�J$��$\������j�f��J�	��':'b�#�m6.�����dum���v��
�gFzP�Bh})宜��n�qiL�	@�����M1t�'�\TWY�,�����얽��t��o��}A[X2�c�Io��LBsyZ�d��G��uu��豗�E���	�Wn��*�K�U�I��Nֹ���&��9͏~��%E��Wn��mZ�rbfٮ��:�Ƅ��!_S܍y/�xF���ʠ�`u7� {x0��\D�"�h]P��Ӥ*�kB��4��VU�*m*sP=[\d��r�v���[z��cU���[��[}g�ң����'A����f�}�.�d��M��;���XVaJ��ݮ}���i@���c)k�Vnb����b��M��i͊me<b��*!s�[��:�F�q����]�v��4�.!F�:�?nI�NŐMCf:�|��Pi�r�v��sΣ؍R�]K ��Wds>Ɍ�uk��R2%��lM�Nv�9γ��ƴ�Z����F��h�A���*](��w'ĝj��(Y�#���x�K�lM5ۼ"Q]
Z38��6v�ܼ��d&�wu��e�&�ttl_o��G..7�	�Lܟ�!To��m�ܽ��ٲy�w�cy�5�V%Έh�\���Xy�\Q��y���DWk۝F�EK�+/k8+)��K�R�R�s/3j��Fr:��<1����:ˑJbvQ:Ӝ��E��͢T��x�9Ѭ�csX^f����	v�
�Q��M�B�����uڰ�Hӎ��ga|��V��zN��(��s;�z�ݠ��҄�k�B��	c�g+7Q��$ܡ�Sxl8E��yڙW`�QR�d�Pֻ{S���]Y�XOJ9�[N8�Iwm
���`Zk8Qv�RB]N��4b�}��uڇ�ֆ�R԰�Ȭ�B�j�I �[x:��"�=���d2�M��B�3V���Us;o��P<��ZF�G�ٸ�	X���r�X��.�9�*ޠ�1Mra�|�����a!�sK��9W':�ص�Sܝl󳳾�
X=:�pI/1�n'���j昦�"7����I%6�So��wuI$��Jm�rN�Q����ے��z�rus0k�^*�Ǧ��D2m,��fj��޵�,l��#��k8@��Y}YV�Y=&�W�v΃W��tاg"��+�)��:JcV=�=JVY}�g%$}��֞�q�l�$��S��A%bQt����-�}�)V
2'M�s�����o�S��+2�&�0AC-	5��EP�jQ7��B�  (o;Hp7��-��V�����5�UIĄ̊��oQ�43������~���V�+W�f�-)�ϻ)�����[xb��ٴ U�;l�%��p96��y�i�鵆5����kc�p�]`u�&�;��0�į����7��F������wD�&��u�
8+>J�]'Bh��V*��
��u6�Jq�"�K\,b]�Jw��p\x���s+�M7)U��#.�C�Z�|.�y��+�;e!��L(ճ��F�K�z�q�����[���S�	q҉V�=��G���[ӡ��3�7��:�G�s;���o2U�i�_`�2�j����:����'ݒ��A������p��Ŝ�:6�0�Ѵ��Q4�[w��,���.��T\R���w����-t���`�G�W���Lfq���N3�B��ZSu��<�W�u�m��L9c� 3Y��8:?u�>.	B�Û���nSE%oE������Fi�V��*��듫!x�[�]쮠ûY�>I����S9�:�K2�������9�z��P�2�@�;[U��R�=�x��-�|��;�����4h��4A�S�����,���zZ���4;��i}}��{�e���S��]��E!��⧋���z-e�2�l׮����n�5��hɌ�i��L�����[�Q�},�@0U���\"��ŷV|n7�;�]�N�s�]v�Q�d��ɹ.ʺ���*�y�9�uǊ|�wt�����k�V��kYN��A����x�����1�BD��\�j�;����.��\�v�=��bÈ�ShZ4����x�HU��{�+Qķiּ�
��;e�·A��Abξ��i0��Z�[0.⑩c�L�y̚�phĦ�܃���t�Rmp=ie��P��2�u�{H#Y��S�5�X���A8���3��J�7�6&l|����_vN�G�L��ƽ9�n@��v��BG�r c����t*��:q��g�VR�֚���1e6pX�F��"/����L��|l�����u�* %2�	5��ۓr%`|��Kojsݸ��5
:v�ۡgt��SY-G��),�r�
b�F��%ki�tq �n.��Fȶ����q��;��QE"�>��`m}�7F��;"���U��J�;���p�1+��ͺD h�Z,d��Ln8�j]b�k9��˷�f��Vm)tg� �YVgָV�t�̫��P��N�$��6MCQ�R�[� ��	��Eh��
:�5/�[����ضE��LD�WK�f���7,-��P�C��������ȭ̒���;�J���[�[z���*�=)��pwF���[F,���na֍��#��G�+��X;�-�のJ�)�����.�]F�dJ˝��Ҧ�_A��8����nɨ�s<�`u
nj�R��,Zs��l7$w�>;u�39v��`t�p�t+6��ZV8��G�I[�%:y{�l�����;�2X���ek�]��\R��_ef�.���IU���9.6�[!I-%�T�PQhL\��9�7�3�m����vu$PFSVJ�9��v�Z&�-����@�:��:{4��R�݀����Q%��(M��u3�r��6h��ur^��Q�pl}i��:��]%
�Vk����k/�� �(5�a��;�Q�)������M��7{��(s��Ъ촺��7��,��c�yN���MY��[KMv"����Z��}uh�++y_�T,�ZRC6
1���-j�Q��`P�CQ���ͬ]���f�6.�!}0�A��HP�z-�����FO�s�R�w��VmxO=2�=�&��� Fdu)���+�VY	T�W-�^GYVk��	����^r�)Q���u�x0B�](`H�ƃ�;䲦�E2�`<C)��&"~�T&nZb��R	tÅ��}bg0���hR�q˄
ڍ�\��X�j�{M��&Q1-���W}�Q�w��=��\ӳ.�M�mb�B�������RJo�k+)ϛ�ks���j�j�1�Z�7�I��x86��wݕ��ʱE���3�ve��3 �|��^P��6�c볷�֨�zD���u]h�)�=�M� g.l%�.q zS̨�o�!u���,Y��v���F�r���َ�ٙ�j�t\vA[����U ��,��9H<��9�F�
����Js,�cN��^��f���X��mJ�9`u��G�6��q�v��ez[�����y�Ӥ�$�b�mÙ8��Jbԥ����HwI+���0$�v���������W_Y��$."�B�p޹Ӱ�4v����0�wJ-6��-��k�����{P��q�����V�jν�sj�de�V��e.g�E�JKf7�,ͬڳ�)Qq�KP�xq��r�-n�ܤ.�*}k�XPv�KB��"-�jQ�ť�l]Ȃ��gV��.G9�n�JdS��Ϯ��WX���"E
�`��{p�\�m0��˧���R��⸹eE��b(���p��U&�`���M&qp�X�YiL[��*�-\�b"�*��*��bʩbVإ�l�+1J��*0Q�T�QX�mc��am3J-AjV(,͘��p�����~<{�^�w�����:���x�}J_�����1�?eGٶ��Wt�٧�_�ν��qw��]��7 Q5�+Qb�7-��	Fc� <���|���Ѿ��A��G+,"=�1%y�I�ۤ��l j^����91�w[ύ1����.�G7���&��/�Kά�̯�pE�H_�l�����7�nPg���#����'+k���Sy�"�L���â�����L�w�x5AT\-����餠�#Pri��Ko����5w��m�G�B_)�~��5�KD`�0���)��;	�kϼg)�{u�������$��A�(R[���	��w`�g&n�Ҟ���y�\�'�ur�а�f��"� ˞�TN:12h�뚈cTs�8�K.��ά����`M+��usց5���Ǥ�N疁�"\T��u�#4��rG8	��q�����l^�jUm�u廷,����%��O��d��po)��,޻�Ӵ�\��^삦��j��3}X簈ҽK3�4U5�ղ�~�#E�2*>b/<�N���V>���_{tS�9,�\�χ���٨X��{wV	����	�"�<ϼ�S|��6�=w+=x�)D+J�^�R`��ӈFE����(��cO��� ��y��̷KRܑ������D]�oz���>V{;]A|�4z�u��)c�OS���sԭ��ޑ��b�v�foW,�ހ*f���\�[�v�0��"��u��0�QJ�p�䰾}�j��S���a*W���(���bNo^�yiB�qHe��3/q��ذ�p��Q�٫�@���Ař�����0��^=��򌝳��&����BB���(�K�\L$0�`�^8�tj��;�5���7�Ņ��/syk�=x��O�3�o����M�V�.q;��<�/��\\�¯8�}4�QApNu��iY�1'5"Ć^�7��|�&���Kr��B���ʸ1�䒴VEW� �Ыu�]57b�m��c�T�Y�"��%�Q݂ϔ3�Z�ˆ�j.N�����33ث�7YA)���N#�e�ϥ��x <�*^��ɰ��	��Ra��7.j��7����"�gZ.�cGiw����q�Z�M���QDJܱ��N�"&�.΀f�p0v������:��jX���P�(ˌ1V��n�j/Y�˿,Pzg>�*x�I��cIL�[į?9����Mwoa�g�C]ʒ	��f8��W�����i^y��9P���H���!Fh��ِP�c�.գ��.��Ұ@��3�nkU�_��\�X �[�]��J�h��a ����x�T��Ȼ)��3���Њ�^���B`y�(�^u襀.yO��o��b����H�$�h�Q�jc��52F �aI���NM*t�]�)������5�����#��)�g��R��=�~�ʟ�g�N_����>�c�zWVV��$���\�}(��[~½����<c�ݒ���m2v�S��Ofv�/.�_�0R��b�������4�9�Z�.�Y�dWg��-8"{�^r����4`T;�0�|�+Qv <"�JW���
��%�q���ڳ�	�	�	��W6lWA�qF5K�u�j��=W�^hIhn�Y��<0�L���﷎��r,�;(��/j;����kN=�)���7�p�p��#|�j��ΘT�xa#�K�t{���xd[|��B��P��閠r���	G�%���uԫ�M�݆[�a��]j鼑n�+;��N+:�L�/�*�%aW�J�.���p��=9�ʋ��W�Ͽ��%���d�~�X���{��x�0,-���QNc����,��S�
��a������w.�6�$r�: ���4R�Q7�l(C<1�e,ϳ�z��T5mJ��a��Lܾ�&���T㝹�6��\��0�5d�����v��s�(�+	s��u��#;'R;{DD)QN�Nw��vc'�?fX|���r�zfIg���M7g�c�|�+�p�Z7�yg�����t�y&�S7 vm�Fڽ	�{n�Γ�~O�/�r���0��f���7A��h5iD.^b�nܱ��ʒ�]a �)j��RX���H�Yh�j��#K!
���at�232���>�8MmۍV@9%L��.�� 5e3#�l�QW�Z�(eCEcYw��T� ��F��*\8�!&�]�������/I�ۥy{��Ѧ�U��ދ,X6!*��q0�V��U�8n`��.^5��l�b,�Lj#b�W�xT�l(q����5J*�J���e,͠����G4���q�����1�%p��j�,�i�ኸ�)cV����+mKl�IX��h�)hV
UfR�81*(UT�
��2QX��
�&,�
�lp��
!��S�YW�C	1l�U�m�kqp�eAFШ��!�Q��m��P���R�R����S�
���͢9V�R�����0)h��
TZ�UAL-�ÌSQQQ���TŕAUqj�N��>q���?t�s�Ǐ�ttA/Q�7d9ҧ���+v5iU}"�s��Si�A��]�#J�Y5��3�<5]���mU�,�~�ZmOȇgo�Z���C;k4�p�0�5ߘ�/H�k$�G�Bu#v�t�z�N��G��Z��8ꩥ{�f�Q}�1��2#VC9R!c8�+�%y;Ep�+�B�ʗC՜��ͩz�j�t<m&d�ԥ齕ޫ�����d���}Z�j*��DT:��[��]��k.�
����Q:~Y�:1�8E����ݑa����T�h��$���}�%'c4T��6��А^ȁ�}ˆ���ۏ_�D�;@\|o�W�	�Ց3F�xL��ӛ�Di<3/.NR�,ދ���=�hʝ�-�&J��+!s�w`�p%����&��;�Q8TR����hY� �evaÙV�Л���(��]/�]���2�WAF�Y�JGqf���K/Ǉ*��9Z�N`�̀�t�b�5�W��n�u���+/m����t�+�p�i���<�犼���/�����8U�:'6��^��K�V��G`i�SXGP:z�V�*-�o�����c.�0�����k&��I�C� �JɶH;�)&����Ǹ~כ�C̒e'���X�cT2M���`d�YĚ@�e�g��d��XI��$�d�i!��~I�̈́� ~M�2�����sP4�| |��"�v�<�4�O��006�\Y!OY6�m$8w����]�]��O!��C�)!���@��hC�$1�I�p����^w�ChO$����dRM�e���4�2�4��Ha	c$=̼���I�$�y'����~`a��B`i'0��0�V@�a�����I+"��,����d>���'�T�C�8�:��I<�f����߷��VB�'&����$�dP��q��Y��O����{�4� ~`L��I�H)&R|��0�"�q����ma�7sw|T	�Q����F����B��Q����W���	Qq�x�l5۹�}}�g��}�s{߿e$?o��8�T�F i��R~@Ӥ!��Y��é�~��?c��d?$�I���$<��4�i	?$���@���	�M��w�k�$��@��e��'��c��`|��HI.�>@1��~����2)�!��HC��'����'Y2�=!�I*d���������H�N�~`em�g��8�8�$�7I�	��>�Cw�����2�0��C����N��Hm1�$�I4��4�m�����;�I&a$�:Ƞ!�@�`i$�M8d�d�$-�}_�߼I�L��솒O�i$�dRC}����0�!�C�!�����g����f�ēH���m$�dR|��0��N�L��9��g��I0�i!Y&P?2C�!�M��8��qL$�M$�HM�w���ݺ��j������4Y���n��h3��}G>7qЍz0v�>��O��R� P���I<�~��C�3��HI0�:ȲCl#��{��Y0�B��d!�OZH^RM01���J�8��T!��8��������;�:Ϳ�\<���Fd7մX�Uw�a݊�a1η[��NR��ֶ��]I���<����*BC���-{��;��װ���ג�;�O���>�iTx�9z��.B�^��J\*6X��-�0��o��VsnZN�۶���q�:`��WdE4	��ud���UU���LFV��ӂ�Ae��vS��h��5���/)�9�"Ԍ�4#%��/ݹ�j�}!؀�c��iV������%��$�w2�������=V�Ӟ�������{���{�u���F�]/-��8wL>�9�7�:>�Vn]���������0\�[�`���q���8��-'7�EN����z#����乏��np�����p���cŀ�T9����U�s�J9���Fɋ	�xWi�|)�S�L�<�ٍݜ�	*�Һn*o�'�o�Q������gOj��%:�u���9B�e�R��$��#��U�d��R����,����޷7�Z�z�u�j��Rҽ�}w��MEt�R�+�H��Q��K�=�DDb����Gƽ�}[�򳆥�z�Y�r��}�<�M)�c�5�/��?G۱S�ғ{�����W�j��p��-x��$w��� �n����޺`չW7<��m%�;�����,����)z����'sM�څ�9�fz �os	f�8������-�vI{�"��*%Y��{9��%����s�sG=R��%�R�����U�8s8�`�˒aˠ��)H[=,��<�.+^�/�Kn����M���k)D�D���W�?w���--��OJ�a�C��5���⮊���;�q��dO�*B��䳌l�޴l��ā95m��}܆>A`�*��v�;(��ix7>���g�&�(�z ��.B᝖`��) ��oX�	�|u�,����?ps�>(X�.����tq��ˮ�4ѝ�N�M*��S�TsU^2�����6��E����Ы�x)MF��vq�U��V����q��s��[�8�� OvuKJ����|խ2{T��,�=WV�F����9�#c^s���4����|9�8_ V�.lh.�=��(��nؑ�m��Vy�����;\�������﴾�~�����J��u�Ѣ�un�8�	JX1�#�%�]�6��+���je�Yk0��2[ww��ˈe,�Vg�*V/��vV�:5u�2p�i��5���I���5@G�:a��7�t��,���m�N�C��2�:��e���X�Y�Z�Us.�/e��!����yv*��]*���T	�*�Tݚ�X����v^7�fa����<U��_�ߩN� �| _ؔj���Ae�?XV�.-*\�p�b!Z+m�2��D��(�eQ����(��Za�3�F�R�#X��EETAAU�0QJ�ř�\�KA(Y�aD����L�L���G鷿~����t�W��s+Y��/����a��?L���~T��Gߟ��2�V�P�v�㪹�V#"�(�ָ<�[�s��X�j�dgT��j�k���r������������C�u�l.a�v�&��^��˭�[B��8b�l\}���yiˇ\���v�T����7��Ss�°�S=��̚:9�c�Z�9u���;&�y��w=j���GM�[Gb��_��D{�eeNi�{�>��e���kt����m��p�����Q�1%e-�Z��[�OB�z�E�qGU4OiZ�#x��J�4d#4��3�0؋-9�jkF����\N9�  �_m�b��Fc-�:��b`M�	�7ݫ"�*�̓X���8P4E� �C�1L�;��],�\F,����j�Z����G��n�_�|���FV�	V�/���\?"oe0�������d<�
�e�:���[���{�tu��vz%M秠��+ P�<�g���؎�l>�W^���QJ���N���]�U���ڊ�&��9��P�Q�Uׄ��N�+�.��S�T{tU6�@n������r$\��|�.�4��<;�}UU_3�G��Q�~���{��j�oTI�l�^�3�_���o�!��gT�xbD��׏�P
W8nH[Jr�<q=�x@���ԯp"��.>� ��T��P�LuX#��L"!<���;�ms�*qD������`��4q"��DC���͍�<xj5�9B��u�VQ�����s0�3��&���#0jn��²[�j����9Ҩ�{��#����Gƹ.�X�w����w�٦���SZ3q�M(=���[m:�I`�f����pӚ{E����V�x��=���S�ٵw{��qZze�j+�Y�uB���XT;��ٳ+�s#���'�Ũ���MZ�
ƩY�u}����ٜ��t]Ӑ1��i-�{i���A����C�N�i��P�\0�|X��|������5�כ�����������G�	��ɖ�d/�a��%"M�i٢qdcX���]��+�i��F;jXl�.�}S�,�`jy���,��Z0��Jm�X{j�����P�����)�k�sw��]��[K��W���DZZ�sM}�p�h����4��j�W]GJ���������r%l]cǏ��r�M��6��|�Uoǈ�����0��\I ��&ZA�J��)5��yp��I���3hA۩X%��K{N����6�mͣ�m��� <���u�s��}�b 4x4@UvMյ��[���M��5�Q�rƻ�E��Z;P��;_a���S�s�#��{n�>��c�m<�Ʒ_����xWV�<���cjj5�It�X�y��ݩ"�Gfز�;�zB�f99�u-fd���.�=ƻexn���R��I�q���ݥ4��Qگ#b�K�\�;��-sv�_�˕ճ�7%s�aw���qH�f߳�;�7H�U�lli� u)����G���͛3��}�-
;9�h�/[�ռ��TL�;x�o�E~i�%�X
B����$��y+ִ���
���]z����=�b{dR�rQ��qy���r1�ͬ䆭�b׷���pv6��[���W���[:p�K����'8En�����ʤ��3�a᝶֪�RVu_w��ꯊH�n���[��ⷷ�=��/�+��Q���ހ�H6��X�;��N��\�0���/O�H�ֽ��Ɏ]�y���(r���!��4�c>oy���!�k�e��n�Ւ5gl�u�ڡ$�'�Գ@�~�g!���}�����G���
/�Lu�D6�ݡ���jY�:�I�q�h�Bp�]Q4it�}H�9=oEL�-�r�Pb�T���|w�S��>ܓ���%\�� �3'9��$�k��J����1��hY�2,��m2k�c��7WٚKG�k�u�s��3\^8��D��x #x]��� �d�/n�mɶ��LQ��sL��|kA(wʖ:����x��+(� �����BhoR���2r֤�S��<�D)��. >��e�=�0��W4d/MmV!�E�,���1fJ��F��+.�(	BU��k�Q���b
��J'Dϲ�YN�,Wt0ڒR���q�^��mˁ�N�ń����J��T]KN�̒\�p�^4\�J��,��Z�	��  �U�!�,���6m��Z;��3�~1�J��E�Z$U[kKK��Ķ��k*Ԗ��TQdL[mDh�V�Er�b��DhѣKB�X��kX(6�\Z0űUe[b�+Eb�B�p­�cPUE��J˛U�z�f���,�JR����iBû9��R�;J�"=�z9��r���F6;o��k�wa����yuz�;;����IoGk��	wN�
�Y�F�uau��E[��tf��3U`���V(v�C��������󡣅V'n�8L����E�u�?nu��u=ݙ�*d�w����vkD �h��>d��Λ2�ʇ��4kƠ�_/{	VL�^�#8E�]��'��'�)1=̕} �+��q�}+��rK[�Sӛ���B�v
�3_ꪪ��������<�7 ��f�t5>�{��}��8z�f�M�R��|�WC۾X�Iuz~�L�u�v���t:F�O?Ng��)� ��L*�Z8`���*��z_3[��]��L��g�sю�^�"���e7.�.���B�9��yJ��*Ok���1DWA�ݷ��کa���k���j���5�E'�5���8��Jw��\\s�N!��	���Uٺ�ZsU�n���׌�^ݩ�s�{��;�gg�By��E��?��P}Yn�*���O�l�O�T�t,xU`�<+�,LZs`�޾�a�Y�C�3��H/�"i�(馷y�{݁��ƴ��i.�&kb��=�:��>~L��[7�~�}�ht��>����}O[���/j$��ς,B�3�r'�0f�5>2{4�ؖ��,��۷3`m�Y�W*���|�w[��9���綞p|��
��T�W.ɿ�!g�/(�j�|��m��Em�MR~�F�X�������C$��D0�Η�.�l։�j�Z_z=��'UϺaȘ�\�dWN7��]^`�_ۻzk�����I�nٛ����'n�N��On��+0��g�\Mn��g��v^�����5��Q��둘N�ǭ�s�o>��i��U�D��1�4�������4�.)���"��B���~�p�)
��*q��U°L���j�~ǙјO�=O�v�4s��G��(ە���>B�UmY��4��	�=ۜ�<i��1[�ˍX��>��Z�N�r�L���-L�^����U�P͝�­����E�h	GQG��Q$���k	�~�w��§ɗRi������>��lM?]
���g��ǛB��(�p�T�*��~!��B<��{*��~�Y��`�hV�Wq��K�)pp�+�Rƫ� �:7���S�ܦ8ڤ*�*�3_!*>7B���8��Zs�޸s.n'�&"�O�u��I���S��^wQ}�BEJ���z2jpx}�b�F�饇�
"�����-��WA��Ơ4������ګи�X�~�f�Y��2�Wۭ\�@w}�nI5��ţ;C�g��܅�޻�'ܙm#���U-UsT�6��'-)�z=�b�"������zc�4d?8h�ee�5���	�5����+S?}��y^�f�N��Μ9���_&�9L�M��3V���u4�r�ҧɧ?S��.��Lc?��Ps5(Jy|~i�-]�mA�~��>�cŚ��^�I�]8~�\#�f��<|1�V��ׂ�}��h���*��i
c�p�.�}�{fhܶͧ�$˱�J��ε�O=�����7z80O>9��&��)�����(�D,�5�h���s|�-��ُ��?}�}C_��M���.��1gɾwg�b(e��V��|ţP�@�X<4�Eo5T/w$�n�h�U��*�S�N\~V :�Y���+©�S�����V���w�)�����A�b�G�蔏(.�b���&�3�~�>�;y�>,�)�Xk6g�a�2������������ӷ����Ä����}�np��\*�?��,o�}�/����~CE��G�xz����L8��>�ѺpxY]��Ⱥ�8��K���K�6�;DR����V�Uzgr����Ø��ڇ&}�?xצb)T|j-�0����k�ys&S3w�4љi�}��9�5�Ʀ���׌�����D����6����ߝ������3Lt�>���q�(�u�<��pp�N�����L�^������?wr3��:��ӟ��o��>�3�ep��O����P�+@�(�U}��&Q��<�L�)�^j�x�*V�b�*W���oèW����jaC�h���]C� �3}W~.���V�YՂ�3�}���r�V��u$��q�������7�﯌*q6���^Y���q�)�o��7�>.����Q����O�v�5�;�s��7�q�12�C۳.��1%�E�=R�
��x]
j��1e�7������ߓN��V\k��U�Ǝ�z�>�*{'��';Vt�Ҳ�O�f9�����}x����Ʀ��<>t�����4P&�ɚ=��+F�)��o�e�||Gվj�f*U��y��1��om���t���q�m�ҁ廪p++cH�|��k87�~�'c�	�O7��s�t��:��� ���s�����o_'�Y�e>f���6��P�*�xtVi�����|=�.'�`�*�mZ��*�pxQ�U����ϸ1D1Z ��X�5u������}߽�y��\�O���{Njϭ�[������*¢5@u��5L���kN���k4x��T���������,5����`� �=�^����zb�z��X�}�43������fF
�?f�\0d5AEF�ޤk�7]���XL�͠u#-�Vk�B|�\q��qe�;Lb)����K�j�Ii�ې��ONX�w./�=K�XA���
�Cy����������*8��R�ö��v-}�u��u�(�
��kX]��K\�G�}}ӗ@wN��=u�v���٬ɘ����!���0���*��+��U
Vzt�ҕ��:��\oIh����p�c�&jmƕ2�.ؒ2:�HǑ��P}.��lZAjV;�-_^OE��ܽb�#%�U_�ݸ���!��^�}��4s��I�Q%�c�����۷[׉�s���|+xY[���eenQ�v�����ESb[{�ў�S��R3����M��C�ʷ6�䥻.��;�}�����/#"��-�ﻹrT\���7���[�W`��e��X����k�t.�YZ,뎧�h�v���wQ�w��b�^r��9��؋�b�U�`�F��("�Q�Uw��¨���"���bŕ�"���TA���ʈ�GUEXb�T�D+Pb���b+"�҈���dR��iH��R���ޕ�t��	.���ި"s�e��{�Ǎ���s�꿞�N�e+��_�K&Sn��J�)�eޜ�y���L߾�]�{�`�)�I�6�e��ϊosWfP�k8���i�4U!L)~��3������m��ze�we�ޫ�F˘*ķ�`�/R�z�b�g�y�۰�>��1@SqR�hu���Z`N4~(�����C{��ϱ�y6�;�C��^5c?V+EnrOy���Tf���5�Pp���%@�����.&�a�Mofu�1Ƒ��ٗ�����'11�+���Y��_������]c��o3)�t����¸L&��)�ѻ��b�+첄c��ۼ�톈�?X�R�5c�� ��/l���!����E�_����9�w�u�ot���8�&}�+�5ޞ�u���~�SI����?Ή�����3�����5k
�ؾBnϞ3����}�M��/�ǯ���5�2��c�9�h�y7�u6?=M�x!o9^6��W+�)�?o�,��+3F�9���]�l�D��q�,,�v�[��9��kD]�)rNP���(��� k{��??�������p����}�~1�譱³O�8<~�)
�}�<f�y��N������yCJ��S�3�4��sT��)��=G�8�gy}�u��2��e��R��y�S�����֮7����T�Dx}�P��>�M6'K�]Uك�4@G�z��|�T�v�˝g`5}^��Ӕ�wI������6�o0T���&�sN�L��ɷ�w��9��ۛ�4Y���b9Qf�|���W�\~�s�=��1{����Y�b�━�9��ǚ�ګ���U턴p��{�Wn��O�?'��5�m��Ӟ�����P���>����׭��}�&L�stŢ��Y��o�O3�=�*i�yuI�Њb�
�.�k���*�	��w:B�hT*�����KH���^?{T��:*���+E?jŃݶ�2���\6������F�||h�n�(e�>�>���4�NC��&F'�S���y�M�ï��p���u�؞W���5`��"
�PU!�~g��#�����:M"[��EB,�]��r�9��]W;"�å�L���X+b�1/��I�}ԦT	�1�g	����O���9�t��}����5l�2�x���L9M*|~ˬ��o;N1|�|��*Cㆬ:��+ޘ���*�r�G
��N~��;�Nf��9����ٌX�gԦ�}z���o���_�l�|�Ѐ�4*��o=��h�ð�\�{�h���L�ݼ����f���|���s��_3/Si�=џ��0�/wgݦ�>�*�W�g�b��(���E@x1^������ 0V{��o)�G6���4�Τ8<;o��eJ������x���:�Z�
'c�n�H�{�ś��}c���>�?0h�pӍ`����S*�!!��
�?�C�V��
�]�4����)�m0��&�bs�s3H-Mt�U�+ ���+�á���՚�7L�q+-pd�s�}��T���0�G�HX����4/Yfq��h?`�=g���i1�o�7��ǹ���0�r̰(��x�L�WY�+G�`��"����ڽ�u!��
��Z��!X8W�]n_�]�/T�׌nu����X��t�|6���������<5Z��2g0P�ʪ�}mȋ�/�_`���w�{3¾�H|��Kゖ}��{�%��继�iCL����x��}����@,���RRG��uS�w�ɑ۴�;�j���}��A�qtd���'^u�3)�|����w�y2����q�传�CϽt.���霥q�'�o�_;�����k�4�T�\�3�kT�6�����5��m�HWY�a��r"]t̝���֐�T8"�^�{}$>�����<`q<��m����(�߾��QL|7��t�?������;��>�y�q��ي]5�0S,���\�$v?<X�(����4�VoUO�n����ϼ�y��^Y�y�s�����s߱���,۷�b
��T�*��1j��<�mQ������?h��a��[�}�(*C\,|E	Y�َ��w�<c_wNߕ�o\'ͻ��й�Cn[����<��7���h��`{���ֳ�}�4<j��*c_���|��b2�"�VT�P�A�ˠW;�ڣ�/�z�����<�&���Mҏ�K�1���1�A�mˮ��>�!�g�(u��ֵN�	X=S���P`Z��*��|�+;}�ʇ�>�v�	��1u.�Ձ�0E����w��TG�V*٬����Ej��n;n
!�f���,*�*�>!��i*�4W��f�|	�6��7[�1>ͯNm��ʊ�^�o'�vt<��G�ez�L�k9�`�>��z{�w]��Z��|����?Q*����w�ے�%����S2�͆߯;�3ю8��N�۩�{��:u�	V���_$Rn�<�׾�]t��ݭ�ڃ����c�'{E���yS�n��r���<�8齦��ۜ�Qx�vo���}M�ϷO��Y��v�x}��а�U���� ��ς��t�T�TH}�LP��u����P��*C"8�&U�l���s9�S��]�s���p�����l�������0|�6%niwp���/}�cӆ����_L�����ZsX���eSɷoP˧��n}C#��7X3��o}��w�&&�@�D������ĕ��n!J�z�vQ�c�{92-LHYu���5A���E�j�iW�"�X��F�pT�:]q��D�X�hS]��qT�+�fm��B��wl��z�>�-IJ�ء?-s���^�{:m�8�	��-%�ݽbM;B��ήlm��Ԭ�ҷ%�v6�`�f6I����c�sF�,�Zn�++Ҕn�`3%^�V��*8e�Y��CM8�X�����ƀc7J���\
:\�ǖy/z�=��4C�fv8�O6N"��/���X���9���m��hM�
*�:X}.�(�Ufa�"r�X6�k�nVN�ہ���� i�И�fث�ڊ�C���	�/�G��ׄ�:�����\7������A�s]���s�Jp��]�v�o�b��k��W���b�e��H�V6�ظY�Ňo��!G�7Z�����k*ۡ�By�.����<�3�	|�R}�h����y�����QfRZ�+#QR*Ȱ��ȰUX-I-����Lb��6��!��1���"a!��+	�e
������f��0&�%`a$P��V̡Y�a����x%	Fu�:��շz�(T�$����ϧ�͌�i����ƩSy=�۾����x0;O0�,�uo�x��ͽ~�.����S��c�t�7�w�mm�g�{'3�^_����m���8μg/�ޯ���;x�n�y�6׏P����q>w��Y×<{�7_r�e�T0Ï٦�&Ǯ��~6�����S	Y�o`��c�ޱ�2�9�����q�lR�B�]-eT4Vi�� mq�Ш*���?>G�/BYj2(�<+�������W�2	�׫�s�t"��ϳ��$����9>����?=�7˴�+3��ưd�r���������SG.&���������) +E1����ڭ�}|���������}��V��^��{}ն~�ׅ{��Lb��YB��*z�YHnӿ�tZ�tn���u�J�k�)�i�ٍS��z�c�羹����Nv�f��=t�+�3�s��<��}�1���h�
�LA������ҘʳT�b�"��C�f�����G���R��q��z-z�����{�+c8�@�ݶ��Ǆ}	
D��O-<���0a����+)�W}%�ꢵ��V�;(R��he��~�t�dYΖj������-���)�?V�Pc>�+5Mn9��ʾMJۦ�X�l��W���	��=u=�#h����NF���g<����u�D���9�/z�YzsM@0*�پ���6�X�:���^� QO�;R���U�e,+�3�S�~�!;�٧���{0�jAS>�&ѿh��S!����CL��K�2Mk�2����`[w��3�^�+�1S90e�Zh�uޏ:Q��y�TSV]��ǝ"�qs�r�6�����3IC)f�������v�OQיз�1�%��^"��c���dȣ�P$�g]۴4Y��o�_p!�WυYFwd�'�~{�w*��[�2:LZ�|_hᰇ,9T'*� ������X#*�p��f٫���YB�61�� �Y��+,,d���1����^_"��Q1����5m��5<�t���{��\a.��ucr� �7.�/�=���W�i���7��3^�ћEL��G���ŧ�k�[ň��n�%T���胧1��>�8ڻxu�ݻ�&���n��v�k�g!���r��L+�e�}���|�L^.f��B���!F��F�I�y����ޅ�m�Skz�q{k��_7kt�6+���"�:g�D0Ѿ��^Ϳ�q,\7G������S��<�Cu�]N�[%�=.;]F@Gr2U���^&�Ipa���l�J@�M�����PY����}�hP�dӖ����H�R�⣩�oƱ��V���Plڙ�c�Ү�|^v�8��T_�V�P�[�{�g�-�"��d�W�9����$���α\��ޥ�̍���^T�ԗf�'�O�k�ߎxVM�}���ʙ���~q�b��S�(���>Z.����uK*�t�KN!5�|�e��R�1v��(l5оw�|��z:�q��z�Y��0=N�u���<�,�z2��[�=W���:�Q�IM5�gA���PفW���gO U�ݳ/��4�)�)�.`��s���4+<e����]�u*@i�S$�P䮋����7�jp3z�:�Z�"1nh��}m��GT3 Uwn�\���v�WMq��1�!���
NC��ws�sbVTE�'9�jgo���h�)`�^�CZ�tO�͙Unhzl��DzW<�S��C�3%&j�|� 9G�xD���6���gSf�Z��AO6�̙�IU�~�뻣wY`)mjg�}�bK��VCu��C��r�ڒn��t��O��U.I]u|�0-�?g�E��Rvl���b�<z�lS�NΈ�!�s�ͻn���
��;���<ݪ+X����5��R�f�kel܋��%QJj��z�,�ׯe�7Ek�S�d��(#��4�w���ʲל���=�tSYI��
����O|�$'�O���M�f;hһ�;�E�x��Q�5�\�5���|�/5[>�6W>U��	�.���%
�:�(DkT�2�Z���Mzl�Z���z& �kaj�B�ά��:�8�U�(s�%-g/{)�F���J+�>��l4[\�U7r�wC�qܬ�w���"�6��N���=�w8M��PR죚�B��8'ϴe�jr�
�r=8a�+�vS��$N�y����Y��V��f6���qb�h�j��G�]�:��Ś�����Q��f��q��!e��� 5�~"d�����	g$l��3jc!}(�/,]�D��VW����vI����7�<�uh��ZX!%�x!n��F̥vj�'���X��#�`x�Rc˘�bP4�*�*q���H��,U��˺H�m�y��rr���)ݪ��UCe����r��	.,��E�P�
�� �Y3�*`I��e&Z�a��aͳ���e�p�VB�Ynn0��W5�QIP�m2��f���E2�Q����
��[Jճ8���ʻ��gי��U��~@ĸ�%�m�]$�W��Sz�o���Uн[�l+�TP�������{�p��؄В@W�_ÁW�Ȁ����h2�f�ҕy}���C�'$>�7L4՞�:�=N���H���^���+u<�ϥ.�j@�ն��;�7���G�ծ\-�CF5aE�c�ָo����o��j�Ե���B՞^������M,�ZjU��WP�<R��.���������t��ٯ~�yf�ێq���SG���w{w��yj9�Y����.i[9eA�B��4�X3�+5�k�;�F������'ؼ�Du���J䷚�Ko�(�^����~����lup4>7�ǨU�[$W
k�{�B��vE�OR��M,E�9ǜ�wn�|���\�W+�x��9Yu����I$��/�q(E��:C8~X���P�53-��r&�[������3�Ɨ��6�-i��&���>��K����}Wu[sq���dŽ�QR�v����u�e�^�����]���F�D�2
�w��Ij�!y+4�9��=��)^���K�*V\)B͵oX�ۮ� �����c�{�G�e�+�:���}�5}&�6"������Կ�^�6��YP4��f��]x�T��НreyE��T����g���c0:pp��SP�M|�R:�+֞�ъc���=�̭�ci��P�k�����C)B�b]��L})e�<���Z��1&�6[E\�d8�-�p�0&�޻G�M�w�&xN�H�0?�yc��G�L���	�6�QnC*�W��+J�&б}}�.��29e���*C{��r:��2+d5�,D��zu���˰kod���H�6��@���,��j�e��7�O9�r���Ώd�P�Xqo�.�R��y�����ߜַ3D�ʡy7��ccxW����Cm�게��Na�1w����U�f����>M�5�.�7����]��e��})G-jF���M�����,�5��������\�j�ח��o�����J�(q�g��>qx���6��w�m�J�!�:\{z7�N���Wbp}�5�H�e��ue�9\D}�G9x\�}��Z}s�%����}|T+����/D�������~#cL��Ñ;o~� �K����[�Yʠ.����	Ĳ�ƽ�j�����1t�4��I�Oّo7S}�`c��)gJ͝x\�Ȳ^�.?ry·��_�qOG�+�z�ݎ�Z�q�L���~�&��������e�]O�9������p�%(��;��$���P{�7�U��ʹ��]���/.s�sO6�Nb�}Rh#����O�d�V-R�b�Q B��A[���ˑb)��54����O�A�5B<߭��_��8������;���n��6f�O��J�걧�W��o@x_Xd���\i�u9fwHx��ܨ�W;��Y�;�e)՜��{,%Bpd'uІ�tf�d��۪��ݔ{`D��C�I��\j��S~4���v���Z�'T�ن����:�������^���0�K�i2��>0���2x+���	M	�"��t��V]�xB]eҞϤ���W��@z�/!/�u�z)�u`�#�y�gO�GM҅�� ;/�cx����Z���G ��XQ��٤�7z�����=aG��=H�=2��2�{��[���<����B��w��cZ}@�{$���X{��������Ķ /��pt����Rѝ�T~��ɓ�ެ��BGF������	��m-ǧ�Ծ�u�Mb'�o�;��Y�3�'JW̤Y�}ۡn

�H���UwL@u�\���/��xX,�W�i�1�j�s�=8m9�%�Їv�5Y��f6bE�$�1L锵���םq�J�@�j؁�j![]Iu�#�Eq�ɼr��Śx[��uy�Gr)HQ$l�+�)W]�\l��k��K�j�d_��`�{W.�[î��O���iJ�VK��i�R�o!P�rmLe*k1�wGmU�s�k.�V�I�:8����X���X���J8L��O�l�0��������Q�+
�U��/�VX��8qx��S2�C�*9��� ��1)M��hS"�9����4 ��*0�Nͦ>Je�Ķ����� g�h�$�Ե���ɬM�ɫp����U܏[���n"�
o4�j�n�.�h9C����R��Z�[oiU1R��.c*�8��+�ZJŬ�q0��)��1��UeKl*�Q�Tb��Zƍ1q���PDQ�����AT.aA*�ԫ0�F��%3��1\5R������X��"*����ď����{��Y����d*ղV�_p ��Ԟ9�j��Ky25c��q�me�q�8]^(��7V�F=�T���Xܥ�tI�hg�Cd�<*�&�-(�c��䂓�~-���"!�o%�3w��� I�6�Q;=�wO!p�T+,�t-�m�FP�x�-�Ib��kϤ��ᮛ��$�G���{�{7]�eK�Uڜ���)��J
TiZz�^A1A�\.�����$���Lj#=+ 	�s��LO9����=Y �V7O]�+��{��u�of�M��RI4��Ćk���ʇ#�V��F�k>�˩�S]���N�M�������a�@������ɾ/�)������RNE�}m��w���+|�Bq;��5���p ���Z�E܉'7��k@��,�R����;���=�K{�٫�����J�F͹�VXX�]��q�����Znj�|s������v�C[+;���E��Wv���V�FT�w�S EZ�'#�-���p�s��Xc��C.�:��i��K9�d0�jl�����v����C����+ڽ�`�l���Y�ծ9�z����ӱ�V��7ztf�+���x�*n��)��7gb�e��@:��">�Qd���ټ���g<<R��'�fmlv�2��*�H���,�1�ci@��bu��3�:���ø>V�~a
Z�n��]>�vK`O¤B�l�0�uwZïT��2#:Fooc�� &��8z߫�'�=0�K��w�roî��}����Z��A���H�Q��ip���ԍ�[Awn�@˶G[+z+np����z�ѵȃτO��y��rۛ�q��YJ�2%!����<�}Ӡ�;2_�l��x�S�Q��Zj��h�;1��&m7]Ԅ5|vV샤�ܕ��Gөa4A#��(��N�$ `�]�[ޑe�x

�P�p�c�jT[�.�[]��n7p*\�ǫ������ƪ.<����<�*x�Be5���c'�R���Y�X��&*즲L�[y���A���5��u�C�n�z1�ģ�]na�r-��B�ʊ7�j�7o,��*��Y�x��f,j�s��ol|'"r�f��@nV*�i��퉺����-�{3r1ԭ{7<�tsK��:��)��Wj	��r�]��EU�{z8��F.���4D�S�y�}�����t!δ5R��m�%\D.Ĝ!�/,�΁՗wY����hX^�u�f�ս������o8�M�n��p�B�4�֢���[�9%%�5� gz8JͩH�M8"�;ǻ+��:P�IO�o#��{�2�r��@B�Y1�~�|If;�;wّ�i����F�K�g�����)vWM4=���5��vd���l���/i����Y{���5����b�Mw�D�>I�{^YCo*��]��,N�ި�x�`�h��{l�H�tTl]z;ӝt�z���t�����7$к��|*k~d���xӇ����S�����:�t�Oa���W(�U���{ژ�ֵܬ�}��4����2��f�[o;Y[�x�k�.�W�|k���,U�^�Zӊ)x�T��#�t8��orH��a��v���,A8��=��:yɓ=9t�<�P�4�e��.\�l�י��Zm��}#5"�������pT$sd�	0��+0�Ȑ�����דj�_F4�t�.[T|�hn������sp�^���U��Ǜ6��;*�Vf��O���Sr�Y�Z�v���qd�6�o$:/ϑ�kC�p!91ug�ku{��x��9������qtKh��� ⅛������8�	f/��y�xJ�YKo��=kp������t�����B%p3�.S(cf���3w�]8�Y���K��z��z٪���`�gDzáX�}Վ�����9hp
�� MCXx���̨�owb��QBÐE�}�RT�u'B���n��� ���.����w���R��-�4n��V��$P�����K	N޽l%r��x�7�@�YRʊ�䵂�4��2�XyV�%�0L5��\��C��-\?�g�,C.��G��h:@T' &�f9D�s.�8�`@�M����r��z4֣H���	U����Xʣ�*�Cp�]d-��7��k�kwnn8:�3��Ar�KV�UX��5X6��X�IV* � �(��*c�QUJ,X�V�Gv�Q	T�Z��!R�+3��E)*��UEf(��E�� �(���U�*���0V" ���6�ۗ
�͢"��"�`洶�!�W�+��P�iB�1QF+F)C�Z��A��T.��n�����ԁ$�����m�����_�K9N8�!Zv�Z�=���y���Ԧ�fG�S�up^T�������&��q
V����.8Es�K�K���S��n�ץ��6��j����L�;E�V��j�.X��QuR�Zp�,�F��ӼZ�b��8]I{����[ /E<��|��rm�ɴ�(��v�Pd�J�9=��G�ؽ����y�8o�^qɼ�5{x�
�6E�k��K���}|�����6�<��v�_�C�Z��JrQ�\/�
|���..��Ӝ����*;��-瓖w�E���-��,���C1Pí��'3�]׆��W(��.t��)�����[�F#��~`ײ�Y�)�j�Q+��Df����K���Z�/�}�nX�Mw�M�<�
ƪ5#�Q$ĩ�>u����]����h[޵|�X3���3-t���%E��j�좤bA��~�<�}���Ygi�"�zq�^�W��3n����k��	HV���8�ΜQ���$����Y��� (2�5��]�)n��;5R�]��3���U�nIޣE��� ��vU�ޮ�W�*�'&F6�O�n'Ƹ��ڼ*��9����7��/�Q��	p�j���W��LO����ǫ�>��EYn9�j����|��g�.���Cg.X���|d��/��Eu�V�u܄�m;	{GrJh����2�^Y���υg����.��U�h��@V����p] �sҳafCY4;�@ ⹀������*�DV��'���Eq�fk|���~��9��̥)f��yQpj�g+3qR�S4��ǉ߷b'ًս7��Y�"B�e�Y�(-	�]�L��v	1�8�%k��W��<��su�u����4#8�e8� 0��]|�P������S���"U�T��~�k��Q�S��m�!憶.F-�J.0r�mg'�"d��|�T��Gʷ~�`���^��q3��;����ޭ�{bU���y�n�ji(�$>�}������s3=��RZ��N�»F��
���CԚ^�MV)�0�f�Zo��>���K��>3m�4�a���;iP�'��U�uo �ǃ:�OJ�ȴ ���0!�b�V9��	^��+�"]4���5"RG4�C�wN�4u�8��.�5��ٕ�*^qW�v�u&y��!"���-n��t�.�.9*�U$ (
a����9ͽ�W��[S���ҋqkTW3�{5�3��Ih�隗�qc��l#�Aev�w�i��S4���O�nڱ�
С��P�y��`ɚ"�&++���n��hy��S�oB�8ysT�G��@.�u�ܚf-�����q~z�fQ�R>��?�K�C��.�5���װ�z���=ǖ�u4���/�"�I�YWp.���_�;���P�����>#����-�-�"�H�@<����ëb�r��QQ]<>Ӊ�n_���c�6��C��w}�0l69Ku��!�ewa�|�U{<�����d�/�HW��6f[;���9�,u��w;��^�I=7s��3��FY�c��f��o��\Jt��s��H�Wk(GΓH�NI�������>;^<��_^�	�yU�t�g_+�9���"��\3��HQ"P�V��[�Qtz����Z}aG�7s%����;ӵ���H};����<�]�;n����!'[8N�xox�'�:�)���l��:��Ej{yWA�.���,���� 噱�Xyb �ṻ:� U��z�m�-I�Vx�ཀྵ�n���,УE-vۏ#�J+���t{8v���ʷ%��QM+�t7z����液u�oFL��U��z�����@=��b�k�w�(�N���5AR8Ӯ�񌢭��7� ����{)ùCA�f��]s�\���x�\����d8A��A��|�rLhU�:�m=`��w����9W-=P��6�l��j,�nʄm�Pm.N���m����V�r��tr�r/�,=�s�U�Q�,���;��[�ey�6[=K��|����-�ێV�j���v�P��������iq���sl���h�1� U��EL�������Y�iQ\j�T�v���c�s5,���q�����Y;9*Τ��A{Bkr���p�ZY��G��j��Ob���8�:y򷋾���}��;�uT�ekQR�
B��cQ�(�:�EUTb��p6��aj�TAX�*�[b��DbֱEڢ��EU��&sk"fXV"6�pb�Y��J��Q���b�J�����т*�sn��`�,Ub֊�.��ͪ)F(a1�
8��J3K�qi�ܕ�_[����oqn���%~F�K�u�g�����Uջ�>��5���&�nz^1gr��zۊ{�̗m��\��֖�j��k72�ޝ�D)��Y��U(�qhut��������x�zSI�CC�>��YT���{�qx��Q��+k�"�T'G�ڬ�}�4���))E���[�e
�6�����1�yfm�m�℡RpI`;9cT��gH##'��'�ܕK@�Ƹmin�Ȱv��yF�{Q�l4�uگ.�)��d������h�)s�wj�@]E�=�C�Ǡ��虧�Zu�S�Pce�(91s���M�6���m� ]OS����N<�py͡hk��A��O&L����|����1k�^�n9�w�[1�u�ػ��0^v�5iHp��-���U+ȅ�T�ؾ��q©�no��4]ǸWL�����^ ��{j,�Lc,vؼ2���A.����q���iy���C�p�=���r{ ���r�Yٹ&��@sxݕ�sn����,�3p����V�Ft��qLqɪ6�]^KЧ�r��t�}���F;����Z�7�����)rnw��zP�SW����1q�=f�O�&�fR{Ց����Ԕ�cztVb/^�{�I�W����B�v�\�1�	�5:�`���c���**dV�i�ƶ�le���5R�r��>�©��ٓ~&��@ڦ:�}3Dݜ��*�t�o����܀b���v*���rn�҅��x���/�2������F9ĕm{整pA�✇e�gOaH�m4{G|�G�*�%��Z�r�,�t���]�qh񣪃��VE��$�=���U��T,�p�F|�N����sѻ{�/2�i��yqx�Qo+a�̚㷚�z��)��<�	ɣY.�S�a}�k��vfE)`(I�)�}�3�w8�e��;�$BVH*�ؖX�U<���x�ס�T���m��z�`�l<4Y��-�Y�+�O*��k�j�q ws�x:uv��j�|���݊o��=�����h���e�d���6�t�i��t�+EˆOQ���$�^�5�i�ڇ��*C�(�4�d�"���qɐ�N��.1ɼ�=
���H^f�vg0P���&��O�w����� Gl�Uz��Yk+^V�͇����L>��9��F��>�~spB�X~�}�V'��[��25�)龰M�h�W:�Qnc�%��z<��k�Ã����K}���ukϸ��S�}��I�^D��U��b^~��fM>;[�vB-��/���N����	#�KY똞���	�~�I����|�Ӄ3"����D��3��H����r{kdӰ�t�ҲB��N1}���OWL�5�u�;��k�_��Sw��^T٣��MKCU:�"�h�]�'7�/s�
k1����ˆ@��*뀙G �{J��X�jZh[c6�a�<��3s�a0��ή�ɻ��:��t��f;���yہd�U��:�bm�y�<����_�D{z�opQ�ܼ�^;��ñ���A����`!WR�0{�lG��\�&i@T�b�Q0����YO�BZ���j��(�z���������WX��/s����>r����YgH�$A�]�l��((�LYs����[ǒC�����y�Oe�H'�x���k�=��KW�r�r%b�W5�_FP�n��\t�0��/��t�:>��>j�ҏW�k�@�	t�`]CY/3h;��`h�2Pb��":�?5�Ծ�2A�okk��:�N���ϵ��^c�n_����?�h?����T�UV";�dTB�'?�(��zK�(��f��E��b�˒���t�v�?�?�&�g�:�d� ��$B��ۂ�ጱ�C<���?��������&�RVp�����.�P�#(L4Nq�
뮟�h�/tb�M,�눡�a���r_���$9�����z��Y���&y�H ��MӞ:��ŏ��� ���* (~�������"Cp��,rzT�媘4S�W�O4���(�p<��G(b t�i�0W�B�c%��� *��y�Z@��]pL���C]�N��"#+�������b��
�cD}���͍�� H?��u�d���V&5(Mr��f����xm*�i�Ɠ�CS`m�-�3k��]��=�ܒ��pK�/�H�be���Aw�����_�u"�ߴ��2* �^�]�0�&V������,]'�v�h�Y[���=8s-���DU3Z��y:������|�cy�� ���@Cn�����j�a�W
�I4Y;�xH䪀�V(�"�(y��`�.��bW:�����^T$IQ��?�P,5�" ��4hF���Qx ���$j^@�M�`���Ħ�	���)|p���1{���al=�Z3��@1h{�ûv��P���Ձ#[٬О��&��@|M���4�'>[CU�����fq^�<��1	�"�bS�Qx]��D��(o:9�a�f���$����;Q@%}*�c���=s�G��BkMN`��;�Z�K�l-O�\A��y�_�ݧ������#ǿ�aB��\�ܪ� �ˁ��c�/ݹ"�O�&ׄ�k��04;��C�K�Zv�T.C֕�Hl� AC�`_!�b��{|�m��d ���v�Sb@X.�`�ꑳZ�fW���G�)Rɑ@=Ađ{4�GNm��rE8P�k�|�