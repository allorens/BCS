BZh91AY&SY�[���t߀@q����� ����bG��           �� ((�����F�T�  � 	 ��T�Q@ ��hj�hhP 5� � hh �� ��j(�u�mUAZ41�A@El��TZ-�
�m����i�e44V����&��
�T�M6b�h�ـ� <�� kNڝT�[j(8�4�dN�"�� ��M4P% P *�٭@ �B@V62�4�#@��S�Pu@��E�  �{�l�VQD���f��.��-2��,¤���[cTj6�b�� 
���j
�=��+C"ٴ�֦���JP�o}J�h(����[�t]����E�V��^�h��(����w] ۋ�Y^Tm��yw�Z^��������M�3}��G�1�a۽gݾ_i v�P�T��+� �T� b�޽�w`1�Y���@]�ʶ���}Y�`]����ϥ Χ� ��^�N�<��Zh2��׾}�D�5A�W�{ﾸuvִ[�}}�J������@>N���4E��i��Ǿ�J��|>����mj����T�b�..�}�����A��ҹ��V�U�y�zk����}���ڕ�.����mmm�j��x W�{�敦@-�v�x�ʆ���֥44��b*���T�0�����%����Kb��n�S[df��m��vU����y`��{ӽ�ӻtRθ(R�m]�{��
��r��t֙��{������袄�v����/}T� s���}jB3��%/j4kb�-��aˆ���b�����O`ӳ��u�V\�A�T]��eF���w��V��iUNJ�u�PU�@ � >}T y>��� g�4k�_pzuCݻN���E^�j�-�q@V{�<��U�͕�s�{��A�t�n�4	�lִ�
ЭU��JR� n�|��l���{J^���zz�����饧�ں�k��㣠ݳ{�Pz&����-�zX��n�:����4�تϢ�P a�B�������v��,�Zd.�
�n���Z=L4�ؘ�Т�9�*�%����=W�ꩥ`� ��Z�ҕ  {���6��� ��}�TzkZ-�849hsW�����N��A���t[�� �4�CN�;�
o   �R�@� @ L�)R�� 	��` 501)T��     S�2	U��     S�%%Abha �2 ��) ʥ 1    $��ҒAM�
y  Q��b~?G���~_��S��b�ڳ��y�<��ỀU�֤�+�
�k�[��  ����@`� ��aTW����H ��/����?���� @X�RI$ށ@\`l"�� 
/������������ؖ����m�lb[��-�lM1-�lK`�ؖĶ:alJ`��6Ķ�-�lKal��	l�6��%�m�l�`��6Ŷ�-�lKclŶ-�m�l[`��l�:b�ض��l�[`Ŷl�6��Ķ&����%�-�lb[L�%1-�l`�ؖĶ%��1�l`���b[LK`����-�lK`�ؖĶe�-�lK`�ؖ��%�m�l4��%1m�lKb[ؖ��%���lb[ؖĶ�-�l#`�ؖĶ�-�l`��[`�-�lKb[ؖ�0-�lb[ؖĶ�m�l�%�-��%�m�l`[�L`�LKb[ؖ��M�i��[ ��-�lKb[�����K`�ض���m�la�����-�lb[6���6Ķ�-�l`�M%�-��%�-�lK`�ؔ�`[LKb��6Ķ%�-�l-�`[ؖĶ%�-�lKb[�Lb[Lb[�Ķ�m�l�1�lK`��6Ķ%�m�laLb[L`�ؖ���m���m�����%�m�l[`��lc���%�-�l`[��Clbi�l`[ؖĶ%�-�c�Ķ�-�l`�ض��[1T� ��ث�[`�lm�-��
6���M0m�1-��lb�l@m���E�*b�Q�"6�F��`�l m�-�Q� ��1؂� blm�lTm���Q�6�)���A�(:b�lm���A�*6�Fب�؂�Lm����*6�F�(�[b�lQm���T-�lAm���1@� ��V�"�b�lm�-��	��[`lTm��F1U�(�Q�"6�cb#lTm���A�*6�� �K`�lDm���`	��Kb�lm����6�� �cm���� ��؈� �"�[`��lPm������Fب�[`�l#-���"6�ؠ�` [[b�lm��� F"���(�[b�lAm�l@�Kb�Lm���E�6�Fآ�`&��li�lm�-�� ��� S-�-�Q�[b#lQm�-� -�-�Q�i��A� ���(�U� ���*�[b�lt���Fت�VآFl[bƘ��&�6��6�0m�l[b[ؖ��:al`�ؖ��%�cLK`� ���-�lK�Ķ%�-�lK`[ؖ��%�-��1-�lKb[����m�lJe�-���-�lb[�6��m0m�lKb[ؖ��%�-�li��-���-�lK`[ؖ��6��K`�ؖĶ%�-�ld`[ؖĶ�m��ض0m�lb�#�6Ŷ%�ؑ�lb[�6���-�cؖĶ%�-�l`�ؖ�IlKbi�l`[ؖŶ	L-�lM0m�lb[�1��ؖŶ-�-�lKb�0��m�lؖ�-�l�b[ض���m�lt�ش��-�-�O��)Qߞ��0��w�9��,��Z�>����-'�N�K�VwwvnF���ޔr���^�Է�ȏp��ۗ19	�*l��R��]P(�]ېi%�	T�H�b��)3S���j��*k2`/�y�[�<�X�2��^Չ)�6S&m�J]햟�g6UO:��ݽ��koc�:n�:�]5!��d�O�,:a�Co��Ν���,rö���T��*42�uoS+'�nd����x.�r�F����%݅�ۛ���J��ku��+36�RpiV�5#���)olid�����C���#Y�Yy�9z��C��qCpub,J9|��˸-��=��S֦��H͸EJĶ�sU��wCV5���U�E5�Z��H��CX����X.�ѫ�heS��)B�kY�M2��� ���0���ظmX�f����id��k��nbӐ�YN\�FW����R�ސQ�GKj���xQ�h�������3�L�ٶq\�;W��ݽ���+n�ś�������Z�s�i"E�U�jj̙HlP�˹3���J�Q�
�(K���+3I^ ��y6��!��6w2�lV�;�6�S�H�
���BU7u̶uefWR��\����Ov.�˛�e��+�������R�&5S���a��:4VI��Z�o��H覲ʗ��'�]�Y����6�1e=��:��vi�u�d���P6fѲU3kq4�Ê�3巖:�Q�N�n����÷A��M��`�������*;��9�iTQ`-<��X�t���KǦ�D^諪k.]Y�kB�)�����|�#C�U�+�EӵUd�.�/��,k-e\��	4cfjڂr��Y�1M=m
%��P]��m�˻M+�yE���uP�$����QTбp�1X��\��K(�wM��h�=n�{l�{м��k1�a�J�Gt�3p�H�M�U[��\WKM�H9"VJ�f���6��nb�G�"+)�*R�k0۔0p���57?P4h�۪6�vN��V��<�Y�Z�΂����)b4��C�6�����FX&,�	VF��2�� ��]���QF]�T�F�b���R6�%i�/\�(γr��d���i�)�	$�KkZ�6�-����B�j;"2����!�롕^��G���/�DF�!$�Zi�6.���Z1�X*�% ��$�ʹ�K��ɀ�VM��n�+p�o�B:�f��q���Q�̶јt��Ʊ�n���9�K$���X��$�EY��6cL�Y�qjhaM{$��n2%j�K�h,>��t�EPgjʤ�F�7�)\�ed���Z���J�Μ�:Vk6@�,�UV1%nj�kv�*è��A��tA�R5��v���̵U��ي���)SFإzP����A��k(������jdK-�-W�RrhXE�{�,�,�9�����\b:A[E����-J�F��Jw��+y�c��{-Bk����\����VjL�Y�d�K+j��l;�wn�*�e�P�ai��Gw�(nV^b&n��9��"�ə4[�AM��[&Q.�Ř����X��ONU䅘�8�2XYb�Ћ�.Е6FRSo.�x2��-��U�cc��:M C�-͠vf���˺�ƛ�E#�b���WI)��YKK����B�M�rR�<�V̲m�˜�T��9��J�N�Y
U�#9Q-"0�¦/)$����q�{�m���.^l��Z2��5�1n��:�*f�J�;��+i��j�)�#��$ت�utn�8Y��,ĠYt�<j����f-�++v�6�X�51q��ɔwa�'
�����XL��j�[U23�^^ek�P���Y�F�H����c��զP%�B^-���D��,��CSt��4��iAN�	bܑ�5V��N^eލD���y�]0���d;�4���ӓsl�~R+ ���BG�%T�M
.��PXS����i�4�*�Kh�Ĕ����R�e���y��VmKD�%�h'��e���>k�EU&��0\'�
R�7p\7#�<��ђ�+T	ӵ����vr r�IrVX��q��4�Mk5v��5P�'�1T��j��C��ɚ������d����:V`ذM�BY�K���qc�5�7I�������#��in�G4�L����V$��̮c�ו�aI����6��LpIV)n�aw4hYyR�ZH���f�`�v��7��b�ˇ� �x�y�	M�"��rB���T,eUlX�6J��v
�խ��	�+l;�/*���Xܼ�)�;�䧍*�.���W��l��V���q��o"�ƅG��QjS�e][ͪV�;�Y ��p���2/0�V�{��[z*+��T�&ifQ�~5�Դ�*��7Xi��hd4eꔬ�m�ml��]^�gpC�Z�V�F'PEg6$E��8��"�8�cd�*��X�8V�ɗ�2�H:��[����U��DBu[t*��gI�`�WVúY.�^[�*T���(\U�L�y�b!d�sE0ἆ�.�clޫ��-f!#	
�ÇDW,8Ŗ��V���5*tf`ʬȆ�������-�˦�Y��r�%4���T�2�&q1eИ��Uz�	ͺ���&�Xuk5lg�n�2���wj�J��c+[z��Gp�;Kme��q�2��<�Z��Y�B�f0����y[�� *[���r��Ͳ%�),�A�z�VAʩT�Hmз�Z;�-�0��=Tݝ��f��.��LB���@����[�$[e�0�S�-ۋ4��jJBm��mл+7�hH�WSk`���X�T�Z�D���4Ē�f�mu{W+^�u�딲me`�i*��n�%w��a�6��u�f��	"�{��ї�7^��mk�V�n�Q�^��{Y�X�%n��N���qe���B]�n�R�A�V�O"fCM��Gm�4�)!T��Va�uGD$36�%g.�ܓme'Yi�J�D��Õ�!��E쩫VJ5J�כ�h6�$r�KѶֳF�X��>�0�Q�����1��-�ve)�̦K��3JX�/f��sq�a��Һ��T�4w�Z���!sڶdp��N�2��isWL�J���5��%��vڥ�flf�8��dl�eeܺ�p#F��A���ה��i^	Y~ѕ������&��Jp�m�bV.��F��Y�u8��0�����hܒ٢�Q��G$,4��Wk*�e�L�oUyzQv����1�Bƻ�j�2��M���5:*���f��nV2l����΢�-�
N��5�L#Z4d���*WOU$�a��*���ׄ�my��H�9������;
�ˣ���b��p�N�%%f�Nk�V�Cq���Iؼ��j�����U3M�Ҫ9�x�n��1�H��C����03S�-5�D��(A�r^e<��]���%�E�9r���{Z!@㡴AҒ����хn�U�*Q����Ed��2 ݺ"a��r1���.0�<M�ʢ��9Lû�j$D���+&��)Qāʭ�t��%l��2����Iu0����^�{xri�n���6��
Z�טnn�x͈�XP���-��-k��ۨ�fnQ{�˱U�iR�j�f%W�v��Zyl��sv��M��}b�����b�;x�[YSpf#-z�C,�b��`�U������{g����D�b�F]�z�<�-�0
-]SwxT�,�+h��mЊ(��8e,�*�iCN��gH�]df]KQj՗D���.[MNY���c�fDM]`�$�P��x�,x�,A�8#,�Sպ�]�0�j%{b@���őb�i0�ZɭRȭ''�*;�^��n1�$�˄�ݙ�7�uv�j�6���V�M��4mV��hF�%*�R'r���̛#�ǭl��(��b	��������mn��6�9wZ�9�HIR�B1��*�\�̖^�R���z�I2:���4��-��H�E�,[sb�.9g"�!̹ܺnB�35���oA�{�ޜ�4��2c{E��JL-��*�ʥLTSYâMF�W^v]Esj�X�n^$�]ZU���e�t��t�BUINO�#a��A*C�j�,����r���J�"X4^l0M����y�2�H��i��bM˰e��d�Eab4���+F�1�A�6�0�Ve�j�]�f�,��+�[��N�#on� ��h��Z�V����ɧC��0�[Z0ꪷN,�i�uSm(��%F]�q�]	��n��+ܪ!�e�CxKq�[FR�ҷI�ՑH�(�p�M�+LT�v��P���m�.m�^�e�T�\^;�q,GW&ܽ�2�:��R��N�Ɇ-��G(]�sN����_��:�6�yv7G1���8��u�f�ZY��֯7�F�f&�j;�`�$X���	��[,�u~;����If��F���mV���qYZ����0���{B��+EƵ֪w��J�#�.�=6��)SdV�!��H�#�afb���*�M�h�lƪ�
��{��!oi��h#�]���n茽 ��TV��aJÚ-)b�V١�Ѹ3ۘ�Sw*�r�u�e�/Ύ�j,��q	L��-B
C4�]EX��ᅃ.�j��"U$R
µ��$Ne�	�)d�%-���܉�ളZ�ge�%������v%�8ܺ0%�=��Vo�R��׎�MŠ��d����GA��Jm�X$��t��u���S������Uzi�PZ�K�m}��e,��n̇�r�̃աjA�S&�f^�Ӵn�j7s��uq1���O�&,�-ܳiԼK���\��jB^��XH7B���Ce�׵��j�T�J$��]xũ��׶eگT�q�j�mU�ûv�p�#��Dp�kT�Ԗ㡒�䩇y18TbPr��wyA!J�㬸�-��4��;�
���[�ַ
*EE��\���g�1�2�DV�J�Wڼ1#�1�Y	9a����C#%%IV�,��u;An�0�J�;[I���xh�ei�Iut1�+C�-�J��ךM�7 W��b"��Lf���\��3��T�e���O�7�)��<�%�j���dS�N��M�fA���R^�N�f��.��,7[�h�UmGS֙M�ͪ׮��^]M.�� ݫ���[y�km�FU��lE��W-E�����S��%ZN]���Ù�<�ZJ�U�8��*�Pr�]��������3�M�9��݊��AJ�)�9[Z.����M]�!�HFwi�z�M��lWN�<D��K���6�^�F؅x�ֹ��1W�^����n�̪DR�n
N:H�`UlR�9��T���VjnK��;J�g9cv彂�R.�L���%�ޕ��m��Wţu�f����!�{���2��j�M�xr��1p�*�-7��W*�7�ε��b��ݙ~�7�w@��O)��@�),�Jl���ю��q�\2�nջJ�Pz�d�j�ԅVwb�Խ�l��T��dLP�6�sPCre$.�0j����ADdᚵ[A����S:��	M�C&��$�l#�@f����Y-ڡ)�[�l�f`7�Z�B�b����اo�[Y=�t6�,KmS�����.f�����H��+U�M,y0U��Tv���`k�PQ�Y6��8m�F2\in*�אbٚ�pK�r�1����m��uy��y��1��-60�F�!����t��a�uI�T,�QڣSE�*e�7V$����Y.m�.�	��96�8��o�M!����j�+�k��JH�۔0�I���&�Z�[N��5ʣG"�7�ln[yui-��3g۷	IJ�������D�g��b��]b��o2���mK��ѕm��I2��4���ʺ���-�[Z�m8�!V�C$9R�%��v�r�,�m�m*�k�\x�[̑:��9�\�sUy�ӈ�m*T�����EP�D(й��ͽMaull �'sc�<�V;��Lm]̉�.���7eL��#��QAЗ�hcuL�!Z�z�q9���]�y�U�[��ܠYr�d©Jh:��iö��Q|���-HX��z*��by�����ۺ�i!G�-t]���{��mltu�5��-WZ�K��B��U���Ez��rT�$�Z��"i0r�7��	����!�5D-���U��}t��-�Q!���c[Y� �����AT��=�Ql���)7�L�3���6)N\�"�[R�2��-u�J?[1&�f���M,�ԩ��m�v���#���Z��)�|���6�_5֒��t�t�B�ު�#6P�7#�U�ށ�uԓ�JZS��6qA-!GR�X(.���թw��Gj�M`%.�T7E��Z�$	�I\�L�����e��:��s��>H�K0Roq��y�)�b�9�:�AU����j�;�=�ST#�{ϩ�oh��X��n���%�-�	GGS�F\]�`�����"�v���/u��|�WZT�A�$!���&Z�����Y�N�y<I�Y�B����HY��n����@��*J$�
�|�r�ȁ"�i[@�в|o�u�(=���N�%�,v�Z��EI����� ��+`"�c���BԚ�H���fRQ*J�(^���[�}b�0�hQGE� 먐2�k!�bݭJ�I��QF��+��K���5k3�P�!�f��*������t�A��I⺮42�HH�YF,h���Ԡ��b	��TQ�œB�6�Υ�
��#�[JX�4�ZƦ���+o�Ε�V��*��U	ҠDQ|���$�JV\��t�X��Q+Q*{N��ȅ��F�x^�yZ4Z� �kn�[��-A�uL��vΓ�$Zi*�\�(�N�].͉P�N��Y�Y��.�k��](����ֵ��Q��E��:��
�a֠���w��k(M�)��A���[�EX�K��7$!�Օr֮hCԓ[KR=L�i�&�8�d	E�J�ī��UUU؄#�G&3�:��q��%McE�4_N@�m�ۤ��\���vo+39�z䮂Ir۾ A��Qr��S7pu�x�I���Ϟ�s`ۤ�����D��cR�YŸ�p?�,�2�#������?^�{?@�*��K��GIφ�G��,rbe�3����-���؝T^�j_^��\whq2�����SfK�w$�Ol���3jV��e ���iYqޒ��G�����3����r��Y���Ch�N��VUl7zS�����Yp��V��zf��B�u�
�MT',��U��9	�B��	��_#{�����ÛV֥�y*���]!�S�u{�fQ�;����mM���w�d<j/-��ٌA��h\�+��ɤ����c2['i��d3
zq�w��G6�r����b\$䅶�1�j>���^�ʬ�3!��K՛;/4n[��(f�gb��k.��V�X����Q���Ĕ�b�$_^�x�-u׬M9�v]�Ol<��h��yR������u�	�Ά־̌�+�����%.�UB{Rْ�7.�o^���^�n����n����q���m�19���AFa�(J�N�;���VMT:��(��Л{Ӟ�*!��Zʙb��=C�vY����u2Pw.[c�������N�����!C�V��m˔�Q*�X�����v�JY��_�Z�tq�r뱊pn��?AJ�=T�Pq��2�Dq�w�y�h��<\����W�����M*5.5�qTV�p�s�Mc;	���w��fuA�2cj7f��ay�B����õ�`��%�f���ӈ�|i<7uw�����8�X7����z#PwW�u�R5V"2�n�q�f:C:>���'�d������%P�z�[͉�p����os��{\Ѣ���]n��f�ou�{�	��;�0xr��a��W���i#T׋��쁍\�j�/k���Pg6���t��g
9
�H�^*|����Y�X�_x�\����3��T�r��1:5��{M�v����Lv�Շ�
�J�Rh��][l��f�ۏ|r���Ʒ���Y�0u�ǌY����Jgk�n��}�k)cկ�(�$�t�@�'��S�7Xnv�b�4�b�����i��wj]d30e�M+���UC�����:a`�Z=n�Y�U:��P;}wln�$�.�Qsd�om��]E�2�FE$	s�	��{r�*m���[NZ}�8ȶ���doB ��cSD��{M�-�qtuR(�R��W��[��o*�yk�J��yM�}�R�����$=O αX�}�YȟtVr�x���Q�xq=���6sI��x��\�i�+ݰ�b����[0jE��D;��V����d�}3/T)\nT�_ ˏ˱ݵ�XB3!ӛg��N·J�b�g�!\34o3�+����1��t�Y*�z��
�trxZ��6RWGV���{s�6��Q%DwFTl%H�އ�{�V�&�����t�de�����"��a>�ЅťǢ�ښ��1%������Apvel��W���wv�F������wmms����\uXeQ<�e\�N��jfև�N��ՙ�I.�Kr�V�Om�^�����{�,��-/��W�S���9h�[z�f]QZ��"7��ƍ.���U�[%	DC˰�9]��ZΉ�ǖ�I��(��kM�Ǜ�ܸ�w-�R��XSwZG�'or� ��1����Tf��pN�Ń��@�;��<�6��N���4�ؾۯpy�Y�<i�OS�*u�ۘ;"F����9�t$�yz9�4��jՇw���S�������Uc2�Pi+]p�Sէo-:���J��u)�R%`(R�9��c{��6�`[YT%�N���i�tK�ɚ����༛3pB���wK7z��0�����fuɉ�Y".�	V��K��L�,�l��1�E�$��vsr7�cS�Y��ܫݏ�R��וU֮�qt|��+�Hà�Ln8�ʻ�"�'V���j.ܷ�\c.���]̬�8�f��,���mbƝBj_��S���m7�궝����q�z��������-�N՝��A��"TnF�&S�rb��6�ܽ� ��hwV,���z��P��0�w�/J���6�[re%��"�wwfu�ݤYP�DQ7���B�&�Krȅ
�6t��BNʊ����i/X�L��Z&dU����B: 4�+:�f���;U9�%��)ȸ�[X�ֵ�4�4U��0�֤ܣ�v:�9���-�ےe�P���5�YU�3'U��g.U�r-�kp�qwZ�@��˗:�wY���Q�n&M%D���{�ۗFT��w�4udw��ue��p��X�I8]꼲K9!�T����8�Q��Rؐ�HD��P��a8�D�鸻�鹆��몸���T�&��5�:��$%m��Xц�&6��J�f��eљ6X[b��c�\�r퇑�E���Ӫvo6:�b�)#Q��gH���)��-��S5��&�����ퟖy9�	��#u��[���FPf�:ÈTP�ƋHT}+1ɹcd[(r�,�ܛK+�%յ[mUM�t��Ր�p^딍1˻���
�l�8*��
�5BR�p���G(��Z��e.�C�c��м}C�Ml�q��^u<)�@�KV�f
Oi��w�2�|~f��z���J惘����\'�혱Vv���V�Z��3��BK�[�:⻫/mh5K[5���r�[�åIq�W�����W-�cOK̉a+�SPoyX��R-������3��	�s��cI�x����ʉi(��㻅6NԼıF��aV�4��k���_[�9�&�٫�(�d�j�b�g���e��n(��ec�Y��wk��t¶*�4y�.�ᴡ�)�e���IALc.���l]��SP�RB]6v��TՐ�d]Vt�\�嫮lN�n�j�t��j_Myi�/r�)_�բf��Yu������S�ȇ�LRL6�)��>�4�u�ݻ��BL�O]���	*��z�u�9H�uL�r��B3(�����ڴ�A��:6���o-��tm�h��s��fU\$n��A����9��(-��[�1e)N���������,�l+��+\U���wB�gM{�o��f��9i�� ք����T�l��S��*C���o7sR�SO�wd�"�q^:��D�Ֆ���ŰZ�ruom��}�l7�FVk�^M���ԕ����b�=fd�ӎ���J��M,9�e��oa�-�ީyy{p�L�q�*Z16�9h񻹢�ջ�%�AWک�Zs>��ܝ�ŝ�ے=��jcRK���zx�	c���ͽU��0���y[شA�EP�4oY����k���h(��N����LZۻæħw'm�s��%���i\�JXb
g0�9��U,d75>J.�+2�������I(�]�x��vS9JMZ�7�������2]0�%A�;�w1�M]�Op�}f
9c��%�!�`5\�˫po]�t�hUc�8�ꓵ�k�������+`.���s��U>����W
�Wy�����j$h�mM:�@�ѤԆ�rr�LPY�Ƽ�r�$&�J�4�FV���g	��(iЬ*��xQ;�5nڮ�X��Zֶn�1�nuui��ZeP�7EF:�7"�*�B�E(hj�)�rls�QL�E�v�ne��s޳m�U����n٭YT0�*8�\�R��X��ּ3W'5���5���@[�"qL*��К˼���Q����F�N���7��t�s���`�s��8��{���Y�t�4d��-�M��[}w���i����&����
'Eai5K71��қ&� ����ŜE���<tG>���"�7\-��B�%,��_U�Zi�z����iG���C��I���K+��/�i���[�V\�}�j�Q�+��M�f�9`W��J�cq�-WUisc�q�@��MY���DΝWq�j��`�Q	ͣ#�Vx[}/����ֲ̳fB��*���
G�^��W�3�ᙹ1N��Z���U٬PE�U
HU��/���)q9[��ͽ�s	D�zɬ��f�Ae�6JX�F���/)]�� k��eJ�u�r�b3P�w���'q��ZX{����A����Lw.�늷[�e;ʡI�wn�7���FlUG9�<ZVwscWX1b%�wc��͖�;U�x꣭Χ���oq�Ʀ6��8 �E����d���Z��tdq�Q�S��S.���͗۲�WU�a�;��[�y���*��(�ٽ�u�+$�DS[z�ɉL<W�S[#^�ը�Ω"oSDVޕs�1��|�ݢr7 :�Ivx0�Ǳi�M�4l�y;W�'t��iړajf2J�"��;^͸�`F��M؄���
�������yR;�B9��mQ�v�j�L�]�����I�++��K��fq��jLdK�Ưvj�QQ��Zb�m�@���!��������=Y�ݣ���*Cx��ݸ���I� �B�R�[�_�6�����i�\�i��ڕٽ�Z�%.:�s�*�wv��Zn�d͗ѽ��p�skV��t�.�.�-,�044��P�S��o)f���G'M��v)z��2�i��G�C�X���!���zm��d��Y(���Xi�179r��9�"���)�5o��c9D^QƎvwc�k}']��j�Qh��	ܟ^)z��r42�����V܂�WQ�V�d�vDS�C;F`�t��R4u���]S5�1�r݃�֤ژ���5���|&�����e�p��t�Xu[i��V�w���gb��<4�d&���_�Kp����=r�^u\�����>�qngs����&J��e���t�ƹ�&kewQL�*�FJ�kY6�1GX�Х�2�C��L�xa�4��%*
Fm�Wn��NI˶V�y}ef	\����K�݆=ɘ�F�P.�y���q�r��d�+V�@ZplH�ͭ�JU�S�,���,P�X�e6N�y�-튭��
(�Z'&���ͮZ*ͷbI�\&�ݯ��U^wm*���E�ni{�u0��zP��lOF������mF�Ά�\�������i+
��������3����fRkuLaB�2 �=�d"^ֿ^m,cG!B��H�����(�gq(�b�C���*Y9��Y��iIXz����<��B���wo���wi�]T���V���%�*N��y:#Y4�f�L�/�S��L���yP�ZXh�͜�]U���)sx��(uo:h�{��a~CS��!��}�J�n��l�n��k[�V��n�b�Qҷpݢ5�H�@���	B�9x�St�S���mSv"���n�h�\�\.�XO7]���.ډ�w+&��jW:\�=Y�qa��ڋ��	�S��J�deK��>�-U����D���K\ۉ1�t���pU=�ͽ�3�]k�V�dl*�q���wl�8]��,�a����8*D�����.T��[���Σe	��q�m�l1��a�+��b�3�	I8���R�"cf�5Q��ج%0���'*̕�Z�}��yWSjh��[�5l.��*�ɣ6��f�sFtl�6�pem�Xh�ZFf�J��f!"L��H*�T�lV�)�#e���`��(K&6�E�0ەH+��"q5�v�*���s�������]��1WO�զ��9�n,\�0���K�57u��6�Y&&�����M`��Y2�����4_��v���+j���ؽ5��j�l�q�-Sڙ�z�+|�{xoV�М=��\��Δ���{pe�ԱS�м���u㧵�³��V'��*joN2�$�.�-�I��zx�׏���]��GM�H���&�+�DԢ�M�e2��;�!�ˑ�w��p�Ao��\�X&:��--:�|��y�E��Wn��Q(�^)�յo��Պh��"�ST�<���ŋA���Dm���x�6+%�U�cuh���1�^ԕWi����2���"���\��$�7wFF����W�����iI���-�9X��^b�ҡ�ͧ�`�RV����Kz,V����!vB���K��`��9u�5��j:�6�fJ�J2k �H���c5Q.ZyP�i��;Z��v��9�Yp���T���%�)��m��Y��Kʈ����e�,��Π��.�U�k�)�ݓ�s؟�ҁ�-N
���].�K���^�Q(��#P�D�%�R�:�=�vm#Ԫ<ܨ I"��$B��	>�/+qZ�yg: ��;���p&�-bb	<O�|����d4+�ju,1�a=a�ĉB9(QGV�7-Z�T�J'�ِ �4�
����WmT���ye��P���LM �n�	C����f]�4��fB#���+D&���)��0LH4H�%)��$a�LO#�#`���9QbQv$ؠ�s{i�D�.H`��C��1/	f`�M	�fN����9tM������� �À@�ꪑ"��P�0�.����d_��� �lw*����1��2շ숕�*w��Ͳ+Rq��6 O�<�N]_J�h�����OTH���H�&&�)�MP�jͤ�Ɍ\�k,]n��&��f@X�@r�-U���Vɻ�u7��=a�ĉB
�#R=h�hQ��0�n�c�V�%-LA'�[NPm�{,q72wk'fa�{Д�H�D(Q!1���d�Ʃ�fM���~l����C�)�D�yr�����A: :*YB�ook�I�A���q7ⶲ�VLn��Ob�f?2�T6#T���2�)]�U5z�K֦���v�?������DQC�t'��������PG����x�?K�~?� _��o��Ӡ�s�P3:b̭�}ƍr��A���[+��uQF�f����5ؕѫUB�����=1%F�ځ����zء���X͚y�� Du��>b��U�R��h"��(�ÞJ��[kE�Uӷ�ꛔ��}�ɜ���ךn�b"��lɪ�ٌ�l�$�F�E+��ݙD�"��Z�S�y<ڭ��%j�����N��c¢D汩��[ץ�,�f�.����M��}7$�Du���Wx���b���9�4�$�c��[O;�5�EP�{V��Jʄ�[�Q	���]�H��fV�u`���1��^����i`��љZ!&��f�d�Y��G��WG�9p�ubƍ�ij�v�N9RU��V�,�
��^�5n"����=�bT8!�R��ɡ�R�m��v-��um��p˘�
@��,ծ�6v�����k���b	��,����4��7���+¹�2h�ɵb\J��%��
�_q�J-����/{*�v�lU�E�-p�(K�]���[�2T�cVt	w�&�X��Z&��,�"�K��26��z�y��2����_U�i�7e�mcӫ;����}�<s5Y2�\*�-�=f�1��{�']�պ�5Ě�eU���v!���֊8��V)c���y��j��n6�۷qƜq�q�n8��8��8�q�q�n8ӎ8�>8�6�8�n8�>8�8ێ8㏎8㎜q����>>>8�8���q�q�q�q�v�8�8��8�n8�N8�8�q�q�pq�q�q�q�q�n8ӎ>��$�v*a���M���\ť[wx�B6�o{z�H��ԩ��(lnLU%E�Q�%Z؅omc�@ڦn-���
.�F��|����r.�������=J�nU��ֺ��j$���;�<���fp�HD(0�R���%���ь���a5��.C.ܻ�¶Т�Iͧ�6uw�*�g5aS-
8Ʈ��桏���m�ʓDe�5r��JGo1�u9l��n��:p��a����#u�R��k��\���f��;H�&�+gH͸Y�A7���ꪋr�T�*����뽓�b͖���qb��"�+b���V��&&qǥ�^�g�U�騞(q�]Ln��5䫹��1Q��Ӳ��9C4�(Xf�9���\��T����V[V�̆ƽr9���UT7��_W*Sc�:n�"ܑQ�1���S�b��Pm��"��z5��Z&f���X�RŒξ�	�C�^m2���	4V�).bl�.�"�YzdWK%`R��e7R^3�A��w��z�N<��j�Mȵ�/qw�����Ǽ�-m��7�����5�UR��ls0Y����ٴ����z�D�՘�n^��Y�\,��v�fv�ƶ��j��n��4A�8*D�D����UTyi�ox��]:\�����Z�a���_^8��q��q�|q�8�8�<pq�q�q�q�q�x�q�q��qӎ8�8��:q�q�_____]>��8��4�8�;pq�q�q�q�q�n8ӎ<q�6�8��8�q�}q�t�8㏮8�q�_��������B�)�xv6J0��ꡳ-+� 輽�d�f�"3V!���st�YjFt��EYj�]Or��g3��9����/���3
2��Sw������ci����8:�kz<��q��/]��m�����r��ej;��si�]m_PVf�b�!��e�7k.�J�j�4]�kV;Td��y-m��[��d-�^$�Q��h-�܇���L=�
I����A�sy����_-1]Z���T'L�FJ�^0�e��	a�WCv��e��(��3r��c���i�Yn�'uF.�6��)=~�|��F3N����3wN;��KKK������:&S�G�NmBr�֖��[V8ܜu�a�+hï���}2�Y�T��h�xدJSt�[\BO\��մ��GhY��9��ܶ�0�f��'�痌�����-���J�t��g��i檲��|��m�����X�֛S-#�[I�S&�=G6�n1�bo/6I�f�S��e�lB�/���5�/x�5i�\��a��*���m�9��u����uݻ�瀓
��&�Ҭ��	�i���\T���f�ڲ
k1����qf�გ�nhU�����[�U�ʎ4�o<x�q�q��qӎ8㍸�8��8��q�\q�8�8�q�q�q��q�m�8�q�}}}}}}}q��qӎ8㍸�8��8��q�\q�8�8�q�q��qӎ8�>8�6�8�n8��>��:q�q�����ߨ:[��;�Fm�����Ά�i��Y�+��\�n.��>QEX��+ާ��tէ�&X9�i�K��X��"�g+ö`�%��d�S��ͫ8�1���D)����h��j�-Zi�ݫ;	]QTjf�N���ʹ�d�=SuDo��.ªZ�f ����,Y%7rL݅�W[���c5|�aDa�^�Òأ���B�ˊx��L��Nd�&�S�BCH���R�������*�v8E���G�յ�l��L����7ةS瘂Dt	'X3m�pҷUhJ�C�<���<�w12�'�6Vq���Bt�)zM���Tۚn��B�%h;"炊�I$�l1m�wkہN�j`�����j�A���A�BI���b���Rs]��t⻫��Q��5��:uhvc��'�J2w�����Cz�����P��p�nԢ�{��헗�Y�̠X4��"�v5�F3��+o�U/".�P�5G.h(_;b��gT�&�O����Ȇ���Z�w��sqA�\UfX����2(m2�ХU:�W�r$�nD�-ӂ)N�ZpKU�s���&��pxJ�"*��M
�S��V��J�F��d�(�P����x��|v��8�8��q�q�\q�N8�8��8ێ8�q�}q�q�q���q�q�8�q�q��������8��8�8��8�n8�8��8ێ8�q�}q�8�8�8�q�q�x�q�q��qӎ8�>8�6�/�g��n��ֳ*s�7*����uS��Xΰ�R�]L���t��͏�� n�d]�|s,���M8�����vٛB�EV�.�6��4��FK��ek��B8��\з6���*��U(�I�8u���/m}	:��n�^��5z��Ǻ�
�Z$��j)��̓�b��p��;^�O5�mu�)'H�jf#K��fe��F�A�3H*HU*(p�{q� /js�͓��iF�)U���;�t�f��|��_;Y��Eb62�]��lR�8�4]���D�4��A��<C���Aə+�ۃ��¦&B�|�H]S
��"Y���pnԠ��޾S��ia��cYWp(Ҥ�$9�w%'�t6"^
Q�����"ԅ��/���hnt Y��u�ke��
��6w�(U��S*�s{lK�����w�D^Gz��h�	�9y;�%[�uk��@�ή�>�׈�5�&�5�׻�^���uZP�̜��t�[6��Bh����?YL��G�������{t��I0N'���̸{�'��Ӱ�xhdCd�Y�+͢p�j��Cu�V�=�E�k-�\WVY������d.�	�Sqn�I����V�i,��:oB,�Y�!�V%Nma���&�c�pp�����zq��:�H�����`Ғ�u]Z����M9H����1�)0��@��W&QL�Sں��I6�,�U-*+O���쫻�@�a����NT)�ˣ8�=-2�:��G��P�N�Yw� Cr���F�oX����Jk���)�u�{֪�eؽ�{���q
�esg����M��	�)2t�U!)�]@
$�"袴�&�NX�P	N������+2.uw�QMI�j��Gn묧�X�n,��4P2�|�����c�A����-��B�U�������6�k�԰�;�o��擗bL�U�ϫ�`"������++�i���rt����pY���a1b�b�vh�q�=���!`�z����t�HP'(=���5�������)|NSʪ�a�n���f�{����"�m��r[ۀ�3b,�6�({zђS 5ی�+����	�t)yP�/4�]ޙ�tی�h�{�l^2���B��ܠ�-�)����M��6mu)�r����~��@���x�u��G�c�s���c��>U���7E��omV�'U���n�;���3ҙ�";��.�/0`Y�2��n� 3S��u�c�ɂ��F7���ET��n�̜"�˕��O���oF<���ZM���]Y���Q�Q�-^��e��)�Yn�7.X�xڍtUc��!KB�͡9������f�kj�F�u��RZf���h٬�6��K/\\��Zk��^��t����@yw�T�æ�jR.h�0�,�x�%U����*"��L\��skd�ݥ�GI�e	Z�kr�7�}���(���*����`�DS�^C�fa�9��P8e�V��I�PhN�b)����ĵY�l;��r�%w�iN:F��.�U/z���Τv�h�PK�ge�S�ٗxt=�
k�꽧g����ʆbɦhVę�N�vk3�ޭ��o=�35$r�˃��⬒Vg���lǷ��pZO�Y/6E���%��r�G.�vT4s���[��(�����Jj�F���������vš�rJkk�s��wv\�Z��j)��N���8'�ؠ��02J�f,z)�Q�s�F����V[�%**�T:T1Je�*�Xt�K4^[e
��Ƭ}��t�Tzgb�^3��R6��B��m=�Z���� XVI��+4�1ș�1I:�֨l�ٯ8����EeN=V�ɼ(�N_t�qh˪���[��%���8x\�s�~"��S��eKER$%�{�F7��)P%vG�w7�b���,(͡�U�t{�՗�D_Lz<vߝ�ӑc���ה,��[�	�X�-r��p�6{��꡽㑺��8�h4/{FnW����pI��82�4m���[���{���٭��[�vn�C�[y�_�#�����l���tS{�Z�5�'��<s�q���h��1�[)4��=�&\��a��5P�؝��t�rs��!!}��v �:��X����O0l�;spT-na��e�y��3fe6��qR\�"�����coN���M5�&@�\+:�^��&$���-P77&�I�l��IfE�YvD�Ӭ4R�R��r�wfL�X8��]��.����$�R9n���^eWt}�Dj�E�+F�<�X���4D�H�ʵ��Ɗ����2�)n�)#��Y�Y�SJ��꠆���]a���L�YY97/mo6�ۆ����gL���S�]��%3v�
{C���ӽW#����2	�.����GD1{h�f��"m8u%"e��ɜ������ت�����6v�5JE�6ZR��\;���1𶵙^i����nͷm�;d�V�M���MY�������v�R��&s&�nqw���dgWo#u��L��ޫ�����nmY��J�p��[]{�'�]�쵻�fb�4P���UR�d����WY��r�k�8��v���hu�,n�Բ�ɠ�
�'�v�dۋ�!)�Y�H�h�ӑ�q�hM�ˉ�Yzk��ȝK��{�`Y���=��5��Nf����:[�A��rrc�l7�	V#[��S�\���G��s
gm�a(8���m��u��dn�1�V��D̄*Ro<ґ���Of1��*-�|^�v�^�Ơ��j�p+�y�y�Nك����d<�A�#�WkT��=}[J�Y䯤��X�����f�Lˑ��f�ƴ�B��Y��[{HZ*uPW���ve���oc%�5.�
��VΙ!�EuU"�+U�s,�y�!kc6ѩ�嬼kpͣ9��i�WK�8$����2�<,JBMq܂�M��3��Z�)˪�,#��l����BY<�n��W]ݎթ=�����&�9��.Ǜyj�i��:��<x��H����V�wT���b��kB�z�+D�6�Kx���$��1%��Swb����׺����ek�޺��a��2#�h�`9W��4���3������,���3sp�Z��m�a��"��'�N^N�l��f,�YA�㳵h=��.�����"�.��������YM�X�A˪6��Cx:inu �^[f��kC2X-����޷�Q�h��
4��z^��t�FY��ot��=˓�],��5��=Ѧ�_nlc���?f<���ȸ�4
���r��7�CQ�:�eelƓ�'�N�<6C�e�r]�ӖQ�Sr̨n(K�Ŕ���ډ^���)u��x��c�c��.��Q��m�q��0���{��ح(W7�2t��]�xe�2i����v�y:�gaκy{nCk�|[��fh��+a�ؔ�.P��Ħ��w�؃M�̫��ua7Ҵa��j���Fݕh�4������4y-��1�{Vg,w�z�ۻ����L:J��(�H�7����dP�{�2�\��y�{6Ե��O5w��5U��g�򶓮�w�:+�g��f�81�21��;���:���}�1�a�:�"�:��[)����i}e�E[�C]9!y�V����p��wь�s]Is�Nojv��R��A�eW��� b�n
:�uW�5��%w;�oQ=�bet��GSr���k^څ�}�V;͂�G�e�p�EN7me��ʨ2r�oz�:�xVʚ��s*����2ve��C�g4�Y��y�B-�ٶ�P�쌧��I
��Fj��x�GX�m�
���B�K!f�y'T�x��k<���X���UCX������K%y�J��;2�����H��5 ��c畁ua=m�	�"(fU����F�q��N0��^>OY��
�2�4f�9#����5j3�\4��)ڇE<睢�eJ�5������n;���M�GA5��M�kJ��5� �YiVfc�[�!y�^��N���YR:�;x�WT���=Q���u%{ޱ�<HBg���7u���� @_�����������������~O�G�(��I��Y�Q"'�H)�&�*Eh1�L�TZ�n�8h���A�Q��TK��?=D*��7g:�JɆ>]ָI�]YX��n��'u�躳�+k)L\]�Z��޼�:k'rĭ���4�\Ndr�5L�&��iS�Ɍ�"��c�ڈV[;1��8��u�R�����K�X�wWv�ѵk$��Y4���W2,�����vG�^u�]� M��K�{�>{�Л�֨fui&�u�&%��^&�U�nW�g���[�5g.Q����j�'_wQ�jX�4��0���[쓚�*o5ҥ�(\u�=ra�˰�8��u�Ѱ���b\84�d��gA�t���ޝ�v#Mz�����i�U�Ē�=ȸ�b�z�R1��G��vkE�A�����j�ŻS��@�oV]���R��1�/�ٸ��Hmv�;�mn��&�&v�����e˅۹�o/c�3N��(�K�Ky�yKk1賍�u��d�����W13�Rk��_9�f��q���q�YQ6�-۵�J;�T������ܜ+R�{ݤŔ��0�/wqi.��5w��)�C�vN���z�{w��7�U�b"X�)8����K=f���n��8��/79�|2�G��I���f�r����j���j����;,>��mnJL�Ɇ�)1��4] ]�E���`��:I���$ѢS`��P�B���0ƈi0��D8C�Qt`�����ӯ+��Ң*����0�M��[�n�O�$�H�)Q)$"��(�E1��	 �QI	��ݻ}q۷nݻ}߻�ow��fEc�ۅ�vIW-�j1�(��AQ�s g��ZI"�BI@��:q�}q۷nݻ~�����{	2)		^�4Ii$�0�w%�bbT�PFo{����{�q۷nݻ}x�d�	$$$"�RF�=���0��sgw.����zx�a��Nt�:z����nݻv�۷��gj�(��w]�ۻ�q��Վ�vt�����u�����2�&��)�"s���֮��ﮠ�&+Ƌ���di�\��(��G�x�Qr���Ewt��3�y��+�����\Ĥwuk�k����u٧]\�x�;��9��Ӎ��ܮm��K�wN���vj��]E۱՝ӗD�uwv�v�w,wn�1�k�ݺ�A��9�ٸs���RM�r���7r:��r���g�͠�g;���'��t�<cI�+����Τ��S?[��t�AT�M�`���Hl���3&h�ȯ.
J��c��1&a���+�t��q))��Q! B$(������N�|N��ېys!��FT�:��]���4;�]1J8l��bu[�m�3��D��j���D����z��s�u��f�m�fز���c��;�u �e��-���k,��o]��/��D�nB�����w-�W�gZ�I�I}��>��U�w.��'��kv��s�ͭ�єk�F�*ʞ0;��&�߆�:	&C�"���x�K	vn_elL9k�H�c�&�и�_;�^�Lr5W6�_(�s�b�6�]�q��׹o>��;� �P;�����(uQ�2o���wwkC��z�2�4�V�;�?Bۜ41� �q\�1l͗Щ֞b{M_�IM�7��g.�l�B��(����@�ʙ��Vݼ�q���ɫ��+w�7���*�:���:Y��_�R���,�]NeM=�]�jf/���+�j�ha)5 ��E";v7j꺤�a.~���v7��j�n*��X�׼=�N�_3����3Z�!t�VЋ�r���.��k���É�١����)����J�m��(;�Q�벁��?��3�eC�n[���I�N�[��P�jef;l���ab]�Q{Sh҉˷J鋘�d2N��S�L��H�X��wX��Jf���UG߱=҈���7�5����"�o���E��^v)k����� NUˍ���Ҟ�8�]�bo��[��A�8n�o�7Ls�%�t�&���u>��|��<��Y/��tQv��(��+�:��5�Aa�|B�INwpw}���V�b��Y+}ؽ����Mh �yK�[N%I��mhbK��c���2
OW�;�(�v �wo=_.����	�۵5;"U�/�Oer�\.�sZ.}�����3=��~���u�r{xጚ�qֲ�1���w�MB#O�>�'�x7�yy*�<��-_�ݽ^�T����]������i�7��
��[���MqWK����8���'z�5��;jY;ǫU������}�'U����#�#�r�:y7��t�����������8�w��>
���Xo�ؓ�Y-�l�\қ����(�·=]��Kۓ�S�o]ܻ�M�iM'i�#V���5�:bQՐ�Ҵ�{�-�λ�)��
S���Uԙ�T:s;�����n��f���p�y��DnM�V:�WB��w��VB�ʜиfYC�VC�;W\h{����ǭ
8߽:��g�}zR�Vm�.��k[D���J)D�+����3Q\Ǵ5�J
7�Ӕ����j�)l��w�0�q���-�Ef�uLO�ĝT %����S��n퀛��/�k�PG0ѻ���ȝ�@�`9 ��v��Ph�xmɌ�<���Dm��Ϗn]{�d珮�@M�>�9VV�<�LŴs;f+N(��c�1�^�|�i��o�[�<L��(��������޽��9�t�Ѹ��TӄS�E�p�J7Jjz��\%q� �`�1Q]������	^����c
�L���z����M���"�L`�絕u`v7gPpn�i�qP~0�J�n�0��p����\v��Mc���B?<��SgW>I��V���u���y7�2�n4���˻CM�́tҼ��6{��Hi��p0A�5#�S�zi
yW�:�.F��f�l��F�*2Qu��j��em�3hfH��a��9Խ����㊼{-���"vlY���dRq�����gS�Y>�y�5�ք Ge�eB��($�w�cW:����q��R�v�پ�B��{�S������J�ò�.�.��xb= �緯��z�^�4J'�owP��(nm��4���t2w:�U�=]Cr�-w�V���CF)�E�7�8B�o�y�3j�ku���Z�W\U(s��'�z�%i$�(�tz]����47��1wz��s�1&6��c愩 le�C���r����׺4@�нN�7�{)pm��W�l��s�G8�P�*���\�wUǪ�w��"�0�Q�Y��,��9���Ga�q#}�F������2F{�OE�`�}�]��}`JLmq�Ls{�e�*� �d�2d�J-�Vtc�O�H��0���ڹ$�^瓣m��]ꥺ�n��!ָhI���h��V�/,;Usv�]T#HV�W.�5�&ed���v�$�3���'(�MO.�b�C�#��ꂔ�g\$�!c�V(��K;m�r$Y�m�3
ʘ��S��(�I'!ݙ�įp��M�ʵ���W�*o�0@�"�n8�0R�F0h(��K��*C����]�W|�i���8|P�;��X(>�"�;�n꼜g�����`�N�K۬3��v|'�u��W�rױT
�D��&I��/.zS3�2��!;rUWn�&�^��Y��G���ҪZoܗa�Uݣ�ذ2���vp���k�vy��Q�Ǭ��;f�wR�F]����*Mz�B/d`�Z��e�e5;rl�c�������	�(Oz�������^��g;���R��*� K��ԝ�Jm���(�؝(uezy�1"�vZUݝܹ�j�{���ϟ]������}ĩ�&�����4H[���Y[\�ʸG��� ���@;W}������',����:�����ga�@m�����u�N�!9ﻦ:�_,҂�;���*8w�����z��I�g�`/L��3�1	��2��8n��1*���r�i���c��F�u��i7�"@���3��I�V.���^<bϢ*.)9�R��e����+2�d����J����&lu�+�*$��k�s�]/JkzR��"+sv��'�e�d��� ��soh�����r�o9gsg�R�^�]�6tU*0�%�b{�Ի҇t��R}Q���l>u٪��+�>Vȸ��Q�4Y�]�b:�o������={�ꮄ��R;��>���8C�F�j�WW��6��LF�Oxk���py��P.�e4$�G��PU��k"����vb{LA/k9�j�K�*dD�2'�9ԝv(v��B��UJ�t��ꈖ�^>SU���I�^V#"��)r�5�փQ�)��o�uﻁ�&�I�w�2>\�B��qcy�7�Qp��ND�����%������gݟ	*�-yzS�����9��17l�U�Ꜻ�X{����r,\�"3����#�u���;��k'>{2�AY�|Y��������;��yLK�uF���p�����n�̎��xua����
-]��4�a��1��l�a�e���a���hs�9n
x���7��=����Q7H�XhTS�Y�8�5x��r�=�.l��=��������J�gX����2��ƙ�$�l"�đ�ᣗ�X�ӎ��ș>���)��u�����{�\?�������w���?��ñ#��D�^62��ا�����t��n��ҋ`�>>C����n��s��bY{����ث�_<SO�ϭ��}����'�Hy�	�7�С,Iq�v�fp�B�.x�E�{��X��
���p{^�Gj�7wY/��kW
�����k�)Y=Vz0����h�_i�f���62n�)�Β�_V����3R¡3��J��>G�W�f󓐒�hmO[}O��t���DV�->i�z���T��Q�$�]+S:�R�uN�v��O�LZK��E�.����O����
�!�(����u�X���R�-޾�b{��rC���R�/@c�%e���c.�nsFT�{��xXf�v��,r�ӄm�@5�،b���1׵��|楌m�MB����JWZ�㝫��ڐ����fCf�����.}xUh�P�<�Q��Z�u��n*;���@�w����ILNLZݹ�Vs�̪�����+O3S|N�\�v^fvu
Yb	hR��޽v\T��l��{���q{ӬD���vz�v��X�i���E���%^�|�����k�I��E�':���6�����Ҋ���U�qC��:d�K7����7TZ�6>l||B]�J�����5��Hֹ�y�X5�ȫK}��~	�����l���)L^����p�Se���{���1�N;�,@ʹhf���	��s�b�+,�U�yG��nl�ٚ��3��yS9�j2�*D��ZY�z���]�����L}�>�$�[��g'x�72^��Mω���h�������m=&s��4�qN�U�+�5�D@�}2����u��E��M���-,��zUm�d��
-�����TOU�v�u{�s����e�I����~�<"�Z��.����r��X߭�t�TӸ���c!mҵzMA����N�Je��"��,-�r]#��T�Y��LM��9��>�Ը�6�����f�/�<�Q}B��;���u����Y��5��f���ظ�JVʾR�j6J���:nt"�����5�\���l���)-��!��� *�������L���=!�f�ׁ�vy�������v�bZoF�nҍ�����L���|���`��T_���!�V�U/,��坖�@�"{��㮄��hq|��ᰲ5T���ʒU-��wؽ�=�!���ۖ��cir�9W���Ǫ�=��Κm�&w�&ƫ8]���8!ߢv=�,>��&�;	S�]���q�,�����¹�F3Բ��Q���lɘ��Y5� T�9��3�M�
�2��Stf��s[��R���W@>"n���cr%�W��;���r����P�K��o�{���4/+�����FVZ�<�Ԑ8���WW�~E, �/��?I!��u����Vf,���r�;��?:WT����G�f�5wSp3���dQ�4 ����o�ihƎ�f]�w��5���2�r�R����i;YVk���hQ�wW���j�S1��lr��+��]nN�����Z$bC��Z�k�g]徥��,�\�&dcƦ�;
np)�z���w,��F���e�9���:�}���v��� ����L��J)@X���p9��fHEOpsqo���ۼ��:�̛ۮ[h[9?R1!@��hOt���V�oX�x�#���.�x9��8۰>�V�3'����W�!5>-BTL�LN�6�p1>d���ϩ�����a{(p�`���(>��:\��{b����x�(F9��oNw=���1�n���&X5Rѽ��g�!t0rd������w�܎���]_���t��:��Ƕl��3췋�>TX,���\7�׸^���9;�;b���]�ϛ�16�Tgi�it]�}n�Π}#L�U�^^&�ihx��f�6]�m8Թ�LP%��.�\�k)X�@B����u���/�[���r��c���{��� r�JQ�,%{�U����=�lA�
����^s>|�T��9vF��Z�f��e$�ɕ��&ԙ�C�i�Z��ش�n'
���H8O�ʩ�sGfun�	�)�6�Sϳ��f��y���a�%*��^���v��Pu3��3��ʄ@����0<RpV�`��X�{9���:��l#.���8�5�J�fԼ"�%el�!�Y>�+l�sm�����M�u%E�\�a6���Ȫ�gj���x��{���ug�@�\�J���1���)c�o&��5����؂58(������dE��oL�s�Lo��Ô�ݗ�̓dm��g���M��Ђ�MbS�ඖ��pѨ��I*U[�nˬ9#2��ܺj�(
�;����^k�:�|���LB��b���t�x�q�q�p�j�a���zVcd�UjqLv{�|�q�Y�EK��ۮ�V�e:�:��&%U�ݫ��3��tW^
��{���l�:�-іrf[�Bg6hQ�m 몋=���T������-�D�L�il�r�q�9_HA%�a�e��%����6�����I�78�-4c#�L��/��sc�k�&��[6:�װ(�]��ve�ҬgqJZ�m�+[w�;^dY�w�i�<��n�]MfcoV^�Q$N)��e��b�#$�:�Af�ұ��T��&g�Q���~Kz��m�{r���Q���pa����\ ���b	`�X|2�t�p�WA���2���66f
\�S>�N��)̓�=˲����ݹ���(��0�E�u�'KZj���4c����4�];��+,0M�*��`�Lnu�{m�J����Ԭh(���mq�����	]�i5�L��$БK�'"�bM��c[��f��)�ƭ���"'�`��R[r�D�2�Z�#�E�	Cː�g-b-Q�5#��eZ9�C�xH�m�f(��r���9��aع�/(����2�I�R���h�+J����!cy��X�{u�[�
V��ɚ��R!�mt��3e��ob����ꡜ�6�V83�Z���|���&��	�R�A��<�(��Ȼ6�[����6�F-�V��WU�z�%��E��ts(7��Ɨ��@98mn�śGUG��5n&�%�:,\zjէ�TM�{m�c��,5y�E��Ӗ���\�i՞��g"��f:��{.|`�.C��ʋ�^e�sY&�X271њ2lY]�a�(b��-�����)ٕ��k줢�i�Bfr҉���k�2-2���%ObX���]Օ.����c6V�����ҭ㙤��cmem꺭�wQ���1U��7S
d9�7wO"�N��UFf�y�dG�u��
[$��Ӫ�T�V�MR��)��J	wh\���ѷF��r�~� (�M��
6d�6&g�na�!���<�AM�z�ݸ�۷n<x����ò20��"Q��;�E�Ha�EDQ�|��q��v��׏8�p�	# �
1�
MDQ�*,F$��5�z��8�۷nݻv���ΐ���h��ni-�i��'��|[�XF幮nX�hBm��6����v�۷n�z9�$4Q�����A�9\��sY4�+���!��E����sd4��>��d��6ѱ�"e�F)1�&���-�r1�*��EoK���Dm0��Z��X�m��XɃ@�^��To���h��BBFI0I/�ɬ̅��U�<טnȺX�;Rv����Zw]ކN=��hj�����`��א�	sy1Y��y����5*���0#03�}�r�G�1��}�j�z-�����|���)W��h�R��44�}��q��m�'�2�{�W~h/�[߇/���<=��@V61��ip!��	7�S�'2�O�c��[�E�9�)�N��Ua>�=������
.h|a�9�05��>_}�"��UD�2/�o�ݐC*�S���b|o��������*�ڼ�������6���~8f�(������c˴Bj�ʖ�޳EKr	���ù����R�`����e�ҁ��o�Z�y�|����ɐ	�߇�.���m�}	��1e��e�b���n%�c4�P ��.���wD�Oa% S*��Ф�n�x��	��x	���L?����uN�����������Y��1�C�r�a�"�s�\`Ksy$e5���'� �u@tX��g#�:�Y^��
d!y4�&�ٛ�c<c���K��*Rr�n(7H��U�`(��e�%�<�&��i�TN;Q�����8���_D��gA��ȓ�=Pi������H��y��l�w.nz���ۚ��4� �M ��0�P��&��{b��os	��X�$��^Y��]�;�ܴ��A�}G>���r�M��p^��6�0��Y�P��m�9N�^�C���vZ���0�eʸ3[�m����b��1��Yʼ/�r�{���=PL���=u�gMݹvq�Uմ�G.�X�����'{ErTn>�X�Y�ł����2o�Sp^ s������
z/���PHp��a������H����$��LxKo��O;�9w��3-��xޜ ��ӛd��.t>��%_P�d��}oy�C�}`٩3S ��i�(�U��=J!� SH�g�L{TM��2Ǿ=>��W���?�D^� � �����K ������T6���s�k��G'#g�Ѳ�y)8��~�a^E8�C֕��ۀ��O�8=��%�<�Ec�YZG<��xs;:��;`.+���޿K��VHl{� O���r8÷C�oH�
0��Tr�w�����[�~����ϑ�2�[��鼚�����G���ovIw)���bՏ7�6$q��n 5�s.�O>5��sͼ�>|�%�縶M��t�y��B�ڂDC��縚̗4�A�� �pu���f,�d�C$b|Ϸ�V>c
�>@RLX��a~>�bG��1S��w�B��[RP�/��AV4oA���l!J/�8�
g�%Ռ����.W����t`XP,��ؾ����k����'��/֬�Z�'��&/d<���^W�����43e����4D1���q��p�-چ�3P�	1��[oi��Gj�&o4��\{���G_31����/2i��Ϧ���G��(�b֏Z�^��*K�$�[pc�L���Nh�wh�L��S\�Y��]J���Uz�i�K\��N�@3C�]�1Gj�VsV�@��n5!��I��"5_� >#��{�� �Uy��jձjf�n8��@ �g�D)�H��B`� �g�%����Ͻ)�z�Rz����-:۲ �r\TL��Q�%�G޽"p��|�Y��N�cb�3�P�5�xȑ�U Yk=��$�����ɵ�:f���s�?������{�O�#¼A�k�:O�*~6|ż_i��!<����ꮯOe�K���;��)�:��	�s@N��x6;4� �П�.z} &;�x��~��zT�����<3\I[���U}'��ܢ�T X�2�7���q쾽y�á����MlbN���=o��9{��O�۽f�柽����2y�.���9ao~�˷��ʹC���c��qw��i̔ڍA^���0��8��`c�`k�Հ�=~04�,p
~�2���ηA�ٗ��ߢr��l1��6���С�p^�߼�@��	�^���	��)W�X/�X�|g©R�©����R_n��O��E-"�%��z�����P9���Ԏ�ghɃ�����k$��� K��\Dwx�����VL2��;L�^��p"_mݻ;��|�xM5c�`�k˼�c����i��\����a�`h��0��Uq���/���\����aR�Z}w��3p0J��s����|i����,�,=ϱ3m�K�({-���Sq�C�����D-N}�t�8�5HI�o���U��d;�;�}���q1�2�)SnA�2oVw{���#���||������k]�d�<�l�^���u�Q�ް��&]���x����f��y	��
I�Ovoct�+��-�]K�x�5z��\$�KW�`��I�ty�3��t�f,�4��,�乱����y�w:�5�I������քv�f�L��*xQc���W��2�Q2u��l�y��q&�& Jk��}ѱIxi}oCqL�0G��X�M>���=�T2G�w���݌�6&�ݑJ5]+��l��Sw}�S_{�yJ����B�Z��_ĉ"��H-i M�A�>69͊Nh�LC^�����c <<{ �DZ��&�B��6s����i��=!ű���� A�GK��}�<y�&�HE�)-q���^\�3/�� ��MN����x���HϾ�TR`�����Q	�p�<#����=��`)�\^�O[��|�y+���Cn\W���iފN�_�T����)�Y�Z�������_� �ң�>u�n�����}��C�p�����ŢcmdxAWԝ���|k�� g��'��X��7'�50���*�곶����  �A@�_���P��v��ӿ��|G˨]�gɌ�,����q���ljm�����y�]M�Gh�PWh ��Չ�J4���0z���qvm���S?[�g�O3s
�]��n1@������me��EF����[���-ɬ�U�EG��yu7�V��3jT�֦�{ �\������R�=<�����4�cMPX#	3\���>|������h�y��}�ӆ��e�4��N��lU3�,�9�77�nV�	<>MJB����t9</��.����H���l����5<#����M_��g�f�|��N��y��VUpA�� ����$��-`
ޡ�\.�M}���-���L?��`&���9��3����������r���1���&ج�o�9?C<;����{;C�Ǩ$lb�7?�~���-�q@�]���/���%�����?Y������VJ�v��PT��)�z`u��҄{c֢*���q<r��M� 1��u�$Q��>50ؓN+�]���_0��of�y�­��\Nt�Ě^׀���jZf@D�/�?��n�/��GFہm�W�vA�q�|�fqz�j+Z&�O�q�/l%���p�3g�L�/�[��h{q��pM����e�E����{���@z�����CB�It�-��z3i�[ �fA8���0¯��<��&��Sl��rWW]�E Á�nAd�H~�5�+LK$�oK�*|XR~���h��OV��xy?H��K�$�J�6u3C0�W>۝7E�Wک�w��l����)�Y����1��a�����D�Ų�nZ�8�3"Pn�K��,Uf)[��Y#Z4�N�!y;�Ղ%z�n�3�]u���h�ɽy2x����i)��iJi�j
H�O6�$�%��j��o} �{�Bb_��EL�S�$�[����d\:�/}�rUU;w�/�{����BF��kP���"�SQ�9�7���zL��b LU�H�EPÛ��msTN��h<���głG�=�8���R�s���1��M�0ٸ�4��:��	�̡�zo&��[=� ���eV��cW���K*���Ǧ�z�2��;���X��I�P>C�L֪����q���g�s�d�r�wM��y85��6ɶ�r��ˏ�~M'�V@D1�1��ܣt��5�:��I�C��V�s��'u������
^�oIo&�8��V⽌��,�6��i��� i෕ώ�q�_�1�g�u[f4�^���k{.���&�Q�^�Z~�T��+O�1��C��UY�j��9�A � �ɏu&q{S�P��~oz��jz��&���I���F�#x��or�]~g�B}?u_�V�͍�/k`w�;: ��F�g~o[u���*}^�=���ؾ0��v-�lJ��x)���r~��8�;>�W ,��z�A_��d��<5|S�7�����?��+P��c���Y�ַ�!9.�㚲I��P\��͉��++*ޛ(����k0�u˱�tvgr��*U��������b^��t�-����:��t�~���"�����f6�dRY	�+m�ɍجeeQ�JpfUi��T^���kE����G� �C��>��H�%膏�x�4M4�4�4СPP�@$��S]��_p�0����� X��-���ﾈ���\]&~�N}c�Q����t �9$�IQT'�8��kp����h`Ƚq[�C&��{����Pz������8����K��0 Xpw�/:�uD``����~�%�j��
2<3n)����q�/E�!�%Ռ�c�������3l�Qrҫ{͸J'��%h���d��w�1d	5�qfE��<~e���ǘ�y ϫ[�[|{'-�YL��M˾ȅE{y��p�����??�������T65;��}�~oo�
�(T�B���Ĳب��XL�J��R�����_��|oHk`(I�Ð�)��}���<"�U&*�_9cgD�g��w�<�	�`I~���my�N�޶��,�0�ѫ�h��p�B�I�
�j��괧q���b����3����7��Ĳ.�6�����F`�~�H d1�ȟ���|�}��gP_R�uQ	�ؤ����G�jD��I1'O��g�V��/ 6/d��PnSx�NX��v�^O�; ǐ"@�i�0�������9����LD+��4D��5�]A��?q7���%���>��7�]sxO��kOO�����%m��=u3�N)�ehnf�"r-�JN�b����od����j�{c��U�n�M*�$4��VM��S�
l;*��ۼ�4Z޻�4����!K���gb����K5=F�gw�� 6r��{�Z>��hV�� �hB��ݻ[uiX֢��m��I �5��_��k����P����ߕ!Dq�ӿ�HÇ�}!x�q��{*	p�=��a����M�"{�s5b�= w����xx�~q>*��O�;B����)�@�ҦG�<���X/�X�;y�yt͕��Ő:�9�|�^_������]��x|��a�!�8�ֈ�>�M�vG�R�Tk��&4n6b��S1D��T;v�{�M�fz:"���1�9hw�;�<K�<���;��ҝ̖�;t��}�(�{�~�f���2/~� ��ǥ�|0��mg^� 3 ]���.�i�Zc�.|(hk�
.:	�,��s�S��yH��w/�|��x�ۡ�K�Q�k�y��h��"c�y8	@�/���/����%Zd.ʑLu@��~x�B��4���q�K�8'��&LG��{a��Lz���M�H"4�#�q����y������L���'��n�j���r��S�<r�����X�_z-������Q���!��5'ƥ����q+&�=�jR�
�nЀ�,���\�10��	�H6'*�0� }��P!�=�*G��v_�;���䩷��3V>��3%��	]EW]S��.�Kum�&��]�'v-Y���)�Ƙ��Mt�����\��T�gGws�|Mì�sgrt�iɶ�����i��'�9UɖY�}�C� > ��4�P �4ҠSM*=�Z�m�kj�ڋV=�{��v����А�pA���zd�9��=�tS�M�a�Yp�Q�����ji1��v}�yF����񊀡xC�Oy���N�]0�ʥC�X�uxqܳ0mw��Ԙ��9G�J���ϖoN���;����>Mƣ#�;2��;�V�l9����PZ�uIw��;w1��p^����R��Z9��r`屧�DkH����kff�c3�Uzdk��:`5�t�Iq���s�1�)�A%$��y����1�J��^%���>�c<c�]^��R@�k�ޡ���Z������*�9� =�b��~�t�*�Cb�l����� �^}��L3n=���;$]G��G���O��V�:]'Gu���K�9��j x�L�aP���雨�"}�m,S��=������ex�#r�~�m�O�����ܠ;��v�G�u�"3��\c�Hfh��(�lt��3�Xmă4�i�_,��۾�x�}�	=M�3d������J��1o1\���0� <i��ĳ�p�<.H�,�Խ[Ѽ�?ɭB�'��T��������&�8�ڣaJui���cV�5�]����ѝtr�����9 ���«#�[/)�W�(��^�H�E�*y�;����<�������Q	��ʽ���3gm�ёM㫫=*�Ժi�]��;"Vc��vy�|�n�^棲���`;��?������G։�u�m�m��V�m��VR�"��"�H��~g;�|�v��=��Br�����31B����|l��\lj~�1�א)�j48r5Eڜ�������^CR98��]Ao;���t���,/�)�o�͑�A����pEF�/i�����=���t�����A�U����JgP=p�p�OBpM����M[}�>�m���Ս�����|��2=�"��a�J��z�qx��$f�X���w���\�Ξ@��|k���_'rz��M$�c�g.5Lc
�]B�.�}�.��̤SH�kgۀ�f��k�����.����J�_a��@Q�m1�[�>��ʟX,��w7�RN]��t�9Y�O�S@�9ڛ�J��lW=`�#� �	� ǡȄ�Bc�l�/5�]���9�<�.`C�����-VɆ$ =���/e!4�jN[�gt4[�kS�P���I�m�sK��QRs�b��L]���C��P��އ�y~hcb{�&�����<�a��y�MƏ^�FYN�����GI�&�a�5!��w�)8�����k�3��>y���{Th�M2�NB,�T ������ȣ�N���r��۴vm裨f%0�]�*Fh;Ѻ����W�2��ɭҙAbg\��s���㗖�D�7iq�u��
��kZ��mD�ʸĩ�2f�^�8I�c1�n�.q,�bdf��Y�Ȏ�wIW���U�8��D�8�m�+�	s�h���D8Xؒ�ҫ��!�x����k�u"lW-D�� xql�H)����-�i_co;��RN�TDカPA[��C,]�ۗ��*��âлI��:S�w�����fY�SyZ��6�r�u�ԯ<��Odc#{����=yO)����3b���qQ��dϥ#��ӈ�^EL��0��Ѧ��M�����u�P�����n4��R�/}�nL���KNh�/nRΩ]T���b�}�̛1qê���E{t$��[3e@�͗b�vF!��vÎ�W�։���/���9q�Ɩ��i�
6֗&�̾�,��Z�J���[x�[4ᰐ�pK
�U
4���oC�ȵK�N����̳�H�)�aB�����'VD��yf0Q�հ��<��Z���E�<7#Hk�OIQ�n��ٚ��tc�}x�r]�*I�y�/'>Y�T��^*Ŷ��H�8Д�USvƊȏhm�l�ɚ�j
�UR�X������;u(�p5�����4vT�N�Y�
L��(ܖ�^V�������L�C;���vT�p�-PYA�o8��h�T.��L����U��EJ�O�]^���D�w��flB��a�T�2�t�8���N�|8];h�4Y%C	�T/��z���muc���.l��B�u�RG��yS��c�.��r��qIX��	�b��l.��9�+�ي���P�&f�or2�Ƚ{T�]fN�Nm,�ٙ�f�oh�xq���!���C��WYu���s:v`�R��3)fz�/)�ӍRtԈ����wnD-&�r֊J�l.�D�[�jM;���+�*�^k�D�E
�S�tC�5rɸn	�1�rk1$�J�oq4�^����.ؽDAwi�nU���7�3uu��v
�J�n�Rk���N����.���7U%+'�o��eÓ!�P��������Xv�4n�Pł�ԩnU� ��FNo5*�6�@�[t�yp��A"�YXa�KO:�of�;|�h5*�c.��V�6�l6�1�^R�o+G3�Y�K��:��t[Og<�Ih���Mڪ���Z�{O��cٛo^��A��k	Q�#�gj�WTu��Yz/ec8���.VwN�:�����q��K�Y���'��"�gz�,��$luw\pBY�%��k��;i`��L�;]��X�h���\���u�нQ�SssnQ܁���,���}�ʎ�!y����Ǫ�Q��7x�cyU�Ek�����u_;�n�5��Ha��L���QvS
�D��א��-� �/R��N���vh���E�[e� ���&x��x�y-դ��"�jB�̦#Rc���?�z��{y�}�(�W�cX�ƶ-Y:z��v��ǎݻv����8��b��M���J��C%I 5��N=z��׏<w�7���7�{�m������1��1�6񷈓78�=x��Ǐ<v���a@���ASv�v�M��$dZ�$��[�M1�q�=x��Ǐ<z�̉ ��! 2,m��)�^8�7mSTbɂ�V�v�U�k�%o;�N�$�(�1��ll�6�TcB`�5�],�ۉF361���F+�nF)��ٔhCDFœ��Q�om\�Q�QX�^}}8�]^�	<W����Όw�D�/xL��p<x���:z��ʮ'�ZO�˙��L!FҲF<�5l]���;�ä�B?���ǜ�<����r�&��*AR
4�R@FD3v�r�[E��v�V�Uk��{��AB:��R�1�eT���ߢN�P^B6��@�������.��E���Їmy��S��u��=Z�2������~W���t�h�~=l=�U���H��א3˜X��n;l5�{&��>g^jOb�|e�{�1�8Agh�`3���p�.�Hl{�23z$�J�if��ژ�oD����>
���%zC+��"@?�煮6~]��~W~���{Gg�eѓ�c"4t�͔�i:Ѻ��@A�q2�[��<�����1С�3�c��S$�v���Wa�4�rX�/j	�ӗ[�+2d��^A�	��y6˜S:|����Vճ�qEʧ-����{��_�c��1���# �m��%3����'6�K�]X�_��\�Lsqfu�Ε��^�P��N@��诶�f˹��;���?yO�y�-(�:�DT�R�����&/�|Ϛ_K��QLh{�^�>���g��b,@-�u�����x-�M�ӏ��7���U����:�����J�r6Ml��x�Ǫ���Iñ�Ts�� D����nQc�{)�&�qQ��S�����u[hz%�����F��WNlcE��/�67\�iyN�(������Q74F$��P��[�1�V�p܉eR����6��ڇ�0Vҍ�y�Q0�뇉��gk4J��Q����J'Ѐ����hQi��j*�)h��"�H�# (���Ϝ��o��f���̐�_@+�
��W=;ݼ0��Ʊ����K�F-nʍך��!��BX��;H�)�S"�s�ִ����j$_���l�v����K!f㾩Y�ڬ5ӡ.�g�dJ��,*����P�r���.�`��B����g�]�5��J�5��q�6��L�� ���K�:�&GO`���w�QaV�y�ںXHOm���1͖�4�F�&�l��8`�Ώ��Ņ�ͳ�&2��+�����r���][pl��tmOG>�ȟS㦒��>�C�~&|9�c$I
��y�!��6L^��2o}.��q�ۖ���ye�F'��@#C��Ť3���	CG�&4?�Tre.�y-������9�+v��'�X'i����ג���]�=x����s�j�]S˾	<4؏'�\���FV_��?K�G�u~wD '(˹���8�ڃ_v	g��v8f�%c9�5KN�E�Ѩ��v|�����p����"�'��W�4��#m��}�t5�g�e�t3g&��U��3TyWP��r�m��I�������z�Cp(�4w`�7i�2U�U�۪�N�'����_#YZAs2M�Y������eR,@˫ف$#:�	:��c�9�.1)����.���y.��s�W҈dQ�X�h�H���R�h�ƚ����Z�Z5�*�������Y�u0�}���X�X�aA������Wއ��Mj�mCr81��C��0ĶS�K����4������P�Q�c������ۓ�n�,�A�P��&���fp�^�+`��C�R߬��`���^�(~!�����Q��;9��y9��<!�Y4!�ɞs`�L:*Ell�<�؆u^�w��D�-�"�
5,�,������'����0>�旬F�x�����5p�C��ew�> ꚇ�/�̩��z~X2Z�׭��}�H�XcNKa~}�.��ƻ��Quq|�Qu��)�]G�lDrεۆ!-!�5f�XCC�~k��[tL�7�$о����XO;����t�X�1{}�h��DC��r+q- �":����M�^���B��,9��*J�/ق�3����0ȶr��Α�����-�[=^Qn��{�������Tѿ*�G�i]z�z 28���:�k;���\����4��R�/*������8�c�����=��*;�|��;b-mg�)[s�b�b.�ƥUe��i�v�i����կةㆾ};�4�_TՐ������Vyr	-��F�|�Ѿ�**����/F.���;�m5"u�4F�Fl��
,픅��"'��s�a�9[��מVo<�'О@BEb�X�4�P#M @4֭sU��v���mEjƐ �E�dE�y��_9���όѯ����#w�ѩ�ɟN=c�O\�i�װ�����\sۗ�+v�X9N��g���ɇ ��׺1���S�F�y�hVC�z*DJ����:���u���fe���XFZ������J�Ce��l�%��d��g��"76n��Xx��_���J5� �Lps���_���$���^��l���(Mn�a���/���R8�6���qx�ll<�󆆪)�g�5n�/�?>P
T^�me{��4Nv�W<�̿l����ʂ�q�j�F|��#z2�}��ǅB�S�Xqmo��{}�M��t�l���L�aҔ��6���~�(2kO��q��|�o��3��iB�R�v���.d���w�0���2ǯK�u���>����Y�#Fm���Q�Q����Ξv���T���i^�ծw����q�1�����p��Dk���[�SSF����bn�;
�5����Ǟ�l�\<{������{<�$oR^�tG�yj}�i�u4����h�(PYmf#���BF1�Μȶ�j&�Q�p�J܁S��u�J�dŒ��xe�ꬪ��j��*TDBH,�E��!���n���l�ܹ�tN��5�n��j�vgN7�J�����o�Z飥f����Xw;��uKvW�a�a E�]h��SR�Z�*���Q#�ҊSM)P $A�4+P#M
!QED��Mnn_�����V���:�W޼���M`�������C�	�����^�z�����cUc,��-0�:/]�O0|E�N��L'����ݚu� �Lk��3m:ݨ����5*�Y�R�ݡ���4HM~U���>;���#��@t�'|�@0u��,����Rr���jڊ"S��!��ݢם	8"�O�\�G�J���쉑_8'�f�p��*\va�U5��0<��T�s�=K�dّI����j��n��7G���O�̴����f�1x���2���n��=рTEZ��
����k��Do��<�����i���TK|mj耽��|t���V>a��Z��c�������4�c'u5�Mٴ���"�U:�b��4C��U���D��e���8�OP�֜�z��rr��E�^Z��4�ߙ�w��2f�O\�Ty~��+N~_�߳��(P�Ā|������v*y̶ٔnU�Ӡ&��5�� �#���Hj�H�i��eW�$cBz�?[�{�=�әX���nC��V|M9Ȳ5��P��]\���Wq�X�0�k���,�5q����S�/����6 �W����ʖ�.3Ac��7�U���9ta�x�i����1�SNi��O��(g[��婲����eVtu��~s9����@��ҫPA�B�M4���J�Q$DY@BD$U�7;�gu8bo7�C��z�.^�=�+EͷzA3)���n�A9YX�K�Y��c���iԖ]C�.9i�J�ـ�\��Јn��:E_�+���gM��7 N��������U�cV(�F���{�5Zy���ue������(:oe?�\:O��{gEA���(|�.&�:8��7���)Ĵ�U
Jqom��$nE�*8ސ�ԝ($�s�'ZP/o^_!�5�C-�w��qO�.��_7h�-���(Y�FOQS�`��1=x;ݼ0�qha����JS�|k6tÿ�o
~�Pq��>ܩI�S"�<���g�zz&�C�mxw�|�Sq��D�}��q�����,��l =m)o[0 ��W�y�7(���,s�5s��]�P����j�荅��]{f�0r�>���R�JuRhmJ{Kށ�ya�:z�y��`D֌�b|����Qy����U� ��W���5�8PZ�Le>�"����=)N(�.gbO���N<�����p/������s�<�F�5���3+��<Uy���j�N�Vt&���A���7�J��/����z�P�^�y*��J\ssRk:J��H�hS�bש��%��������s��T{�8�2�鸝����[S/v5�d��'[�]�N@���G:�}ni�/��-�s�Y� tF) �� �4�%E�nΪ��ծm��m�mFک6�m�b��m%���x�!�[LͽHW�ݚ��0'(�k�G�@�d�V��A�b2�4��5��,���ɚ-зf���L;���ێx��,k�[ ��k˼ `X6�n���4�]qS���¸u <Ӧ�R���[��?��7a|�#��ك}�Z�ȧw��x��2);�M�'�9�w�X�+��Wn���l<�/^J� ޤL��IMD�-0����j��vv�R��d��μ��t�Iϧ�°�3�"�匊�}cab8���m��(��y�z3Ur�?'f+�`���/}�L�8����È�Ml�����þp����i����[rǤ7(Ф�+���v��'	Ĕc�|:�@��L���{���Nv�P����֑�p�~}��eq*}�A�g*��f=����Lk�]j�1F�SҘ�X�{��S�6e9�x�)�ˢ��4�c��tW8!��9��m��R�6DJ�A@���9��2 �o����Qt��T��!�i�������9����j�.�;\OI�jݗɞ��)2�7g;z-����6�[�T*&.
�j�^��ى�yLn�
uF1��M�&oR]2�ejMhɐ��ӄ3�N�����B����N��Nh18��i*��O��y����Z	f����T�>�S����$i�J��7n���v�V�5���l@x�6K����k�|�^�GG��h�9u#ů��+�"dS[���a��Z���jsKY?U�?���靏�E�����B�p��=1���Q�o}?U+	�����|i�& 7]ʓ1�e������4��\Dcy�Љa�ã��ֿTĶ-���*��%ߐ��&�
�2���A/r���U#*u�������A����'i��l�&�6/���u�8��s�b[������LsI�<�ۧ`3c���sOR�,k�1��.�d��`��
�����d׹?nr���(nu�w�O��ƥ���|�:�O5
��$m��|�&�U��'�Mm]�@���7!�dI����B���OǍ�[;����@�n�P��F/A��]@� \��3�� k���%�ލ�0��"j�P�DnP��m����G��C�ޭ��~�/A ʸ�C5�SD�DsKH!G� ��X�sx ��/��1�c-׼
{ʼ2G��3{Cq�e�)�����[Ӛ��l�GH�x@fE�}ѣ|X��3�-҇��+��j��E��ٙUm6z»�Ac�3ٙ�1��8�9��
��%�K�����]�1C�6�.1m0`(�>�5U�Eb�e��e��n>��Nw]�N��iˆ�`�s����#�⺋��74��z������R� �Mmʪ�-H-�Ѻl��S�2��< ��~4��J)QcM�AdcZnݵ\�[E�jض���ȂH�"�9Ϛ��ߗ2 z�����8�"S]�2�&��c=�#��,8N'�8&Ǹ9�1
�$tb;��4�Z���>ّ�^�9�5���|�.�$��^�gG�l��œ��q	G3뻪��LWm��(��Ԍ�<s��,/Ր4MAǟ(�Ǽc�ES���P�-趋{٥m�$�ݾ�a��/Q�燐�͈V(��s ��+ҞDÐ�|*5�^�;���V��fC�m�(�=�6���׾��j|�����5�9�����}{a^AG��D&ݖ��F@��{[uM�XD�H���`vjvcX�׸ŧ�e#�F"�4�K��-� �ZD9��e���k8_&���V��6��A ���(M�D�Ǐ8���r>����~�e��ٱb���T���I��B���J�|'_��R'��m��s]�:Rq@Z����hz�[�	;�rX��6���x��vo0f`�2��{����i�_[,���~�a��cέ�q��a��=X�p4�˽\��5O?�P�e���`�D�|d^��>Y�����Ѵ��=㽛�tYF*x�1���
���fѵS��4��Yt��W���Cɳ!vت���'&�b#}��s�Gf�ꧧ��Hh_ #CĊ����M@�_Q��r�;\Aᙇoe��YKo��v�����ay�,Y�?�}��Y&I�1uƖN��W������i�4*Ё�HTTcM6�n�[k��֬bԕ�ff����.���
��w�msa~�Gc���hP��t���	�ֺ��<���}�g�����g!u��� �)=���|���V�+���~3��0S�0�������k.Tӯ��z�4&�e'�%�A���<�>/�i�������3M�zbrnhv5��[�˞)���NN�ؐũ,����h;�|��f=�-̌� �{�8��޹�X�ء0�"QB5�>��ϫ�'��:�҂{��^K��<E�f��i�����{1�LT?V�f��,
���lx�? =�jg��x���l�r�d5AVd��~�`�����BM&�f�rq��ɋlg���"��|�'�*Sb�ow!>���4���rЭ�9ȴ۬T�@D���^�%8��d��m9�ߵ��Zt�L>��i��S�e�~D�9�3���A�Y쑽g���������B��������2�C�A9�<,�0ՓUͱ�0�?!0,7����=}t�1���S"�|�7�s���Zь����{�x
��Z�ʩ�P���K��˃	�ۡ��ܐ����9j��+/Gqv�6z�a�fc)��:�;4՝�1޻TN��Q��a�d�vr��Xkq�ݕg�����	c)f-ݥChU:!۰�P{g!��B�J]6få&�),�F6UQ�pF��(��]�t���w'X,e+W���F�&�����>(�`���fj����{�,mm1���u�S;�/��I�Bx������w��N.�2�ݗ��UU�y���5vn�W�8�}�*��Ha�MFC��	�0U�oq<��c3U�]!ݴjr�3��VJ1�p��W�Vd�Y�:�m���\4��j�XYP��o��r�eq}�y�è�Q�j�[aD��s.U���U/0�%�����蚴��B���M�1��ڊ�u�g�J�e������Y�#
)���;ws[���8�� ��p@�aX�M\��u�*���1i5�C�[��q�b�N�-�Qm�&V6i�ɛ��`Qm����p!̌qcf�j�0�W��f���c�YMT�qUe�C%��u���m����e�][��mḳ��,���4u��Tȡ��Z튯f�N���'��x��;��ZOz�&��s1o�ɚ�TNf��@i,ㆪ����)"0�4�q\�ӏ2^Ԩ�D��]qU�5�P0	9�,�m��6��3&�+Cv$�8Ž��Ӹ�u0V�{URv�3)�}wK2�Pm�JŃ�ف��}8q�1���|�4�sd�{��k��!���)��C��l�3�2"�8;��ˊn.U�t!���8�eǷ8�6�䷉D�L�
�b�F�7v�Y��%ٷ�PZ�K���n������������J��R�l�Hf�yJ	�k=�+�����e��b��|�+�L4d�٩��ۏxM89��v�J���G+s�,�Eμ�VL�*�j5r�h���2yd���̨j���0�!�B�&6B��C�t���{���)ˬ:�̇���\��ӻڻz^K��f�2��U�0v�ʗEf7�BM��W!����+���Ո2�GmR#B�v�h����uR�ښm��!gf��dDV*N�B��o��˪[X�]S*�N����Mw��X��tA�Y��.k4�P'�oQzk�Z;$�B��䮕�p��RkDKXO����
�(P\9y3w2(�p�[�w5W9��;����圹���aQ�}3tʙ2��$-�C��G�N0r����&���zp���
"���k5R�̵
W2���=eF�.q���a�AG\�[6ދĺ�b����.fU��\��e��8c��U���f�wF�ؚ&��Ż'p;i��[',�2n�&��� ��l�yL?�u3S�n�r�9�+0�Dn�I�̔uZ�l[��9Pr��7���2	��"E��v�mE��F�����$�F@���o�8�Ǐ?��~���|�+���J� �61EF�� ݣN8�8��Ǐ<x��ם$� Qc0�fZ*1Q��*Sq�q�o^<x��Ǐ_��{�����&����sW�V�(�`�����x�ǯ<x��ǯ^��E�d�E�9Ez뱤�i*6+zk����HUm��Eh�)1bb,���F"�65�A��ܱB�F6CE!�EQ�Tlm�WQTV$��Fѓ,wu�ĕz�k� �'��	���i�s��/lE�+���UM}U�{�rF5;�▂5a����B�9q0�e,�ѱf3W�Am�h����j"B	eћ�\���ضƣm��E�;���K�=���������.[�����L*����PnQ{��Ic|��T���J�5�k]�;B��v`|����ixhN�������RXk����-j��UݑF����,�x��ʖy�.�qE���-"(LhLe6�R���ᒴ#�b�C�Ȭ��q�3x�tB/maTW��x�Z�9��]\�C��+��~J�,�'�9L�n�d�3C���};^f���#��9��WoH�w!��4v@f�`��:a�8G*&𶼞�7o�a��͟C�H�T���1�O^!��q���s���&mM���pAՊ���.�t�m�K�
��bo%�@NQ��n��H�homA��%��a���q)ZIo?}������5��'F��C��~��B�������(�-�s�P�.�U>t������w%y��_l�jP�*��D�/ߐWnb�}��[Rꑍ����4�*�{\�v��Rkt�9��YוdPu(	�_d��a��מG=��KKS�g-܉g�kN�R^wPsճ��ޞ�vl�\��7R��xo�5Q�v���Y��;$ްk��ع:���ɬݬ�P�"DA0jSb�ڋ��fw>w��a�5��0��h�]�w�Ε��"���Į͇���]y��5R�ލe�ff�����J5
��mr�Tݺ�5���r�y�{���7�^�"ƚկQ�����ʟ��~G�훸f�I�Q����G>�_��������v+yx,�R����Є���g����L�ʡo�v��ǡ��Zˉ�Ⱦvs��a�xCCi~��Z��f}6e=�g�b���)�FS	#gq��A�y���;���:�qtF�Ƙ}�t�7�o���酂�Iu��Lk���=��c�r�!�}�(.��;�6��l�S��lT� fH�^���'��O��J���庾��w��;�z��,�mӧ�\s�����.�R��_���3�Q����F��/.��M��*��Z�|�����3IP�zY�KӼ�F��;	v�]�=s����i��Lr�l�g�M3�@��͝`�����%�_U�U0u��K�"+�]�{bd���<x��1��ǌm�[(��dL����eã����3����=�npD�7��<�!B���{HfB�@x����g=K�|�p��7��d��b,�zGa�����o��?L䝎����#���1TÊMC�e ������Nκί��z��J*�q�E�c'*�k"�طy���g^c�Y��L~'*�r�tޒ�9�y����2ʔ�a��D�M�0&՝��#C�{T�=���z�KXJ,b��nY²c��Z�ޫ�3"
M��8Y^���5��y�J����J��B4�Unlݻk�6�����98x���.lo�؇lgw�XF%�Mg�W�u}j���2$��6���'���W��DM��D�L76
-��~ǆ��D��:`���`T'��|c�'qxT3�nQ���Иvl����u�)�3zrB�*���ʰ������l�N^��8��\՗P_����zk�20vB�)��#��l�zǶp��S���n[+Iɾ�z�cϢ}.}�g���5/n��ɪ�IzK�Q�1�בx�_M��ndq���^?>L�<;�w�Gd7�Z�l}����:F%���/���s��DF�~�Gv9��N=�֬�Tm-�PL>O�.�T��h�0q�D&%���F��ԓ�gM����ބ;����Rkk�gm
;�K	�pʟz� {��BǕ�fuJ�؇��:�1�c��v��l`����렡Je��h��o75b��|�>��8`�{0��Sc��[*�|=R���ʜ<��$���v�0Z���y��i�g�m�fi����D[AF������D?%X��Nf/�4��-����̿./�f��d�~��YW�V��V/�ː�ѫkk1=U[j�2Lʻ�֏�	m�U4Q�G�a�yZazq��ѫs�w��͵V1�6���[���mv���i��Lȕ�o�r��J.�N?=���#�Е�#M �MT�4)QY���w�u]�y����އ6�����P���rFy9�I�s�|w��}�l�3z���*���#1J1L�)�(N�[� G:"`Kl��s]�zRqV�y<ڹ>a*�F��;Y�2�����Ξ[��6(w��CC�����=	}l�Y�J��<�hؓSA��>�F}^��t��%�q�o��ݍ����?
_Z�A��w�h~y��~�З���`�9�:��Ԓ�S��Я%|U��qɷ9Su�<���W4��־5�cS)�|Qc{�z�O�,���.�kh�M�u(m꾽��=�1t���k��?uTË}S�"�ʌ�d�#T߾�m�J8�h�&_�ٹ�B����
��26�	!z�zbϹ��G��7�ef�/@%�].�_��M�V��<L�ȃ�r��J���g?'K�J���Vz�kd0Q��,���hH�i�lj�K��:B��N����vzgX�1�F�=�A�(s�0{p{EͲ�I�v�
=@>�{���s�Z}�p1,}���i\�Q�#��Qw�`��X�aϐ���~Vk3��yƏ%�3ᗭ}:k�p��V��^V�Mh��K0una�s�X�.^��%\�s�y~X�+?�|^�/9�7>��W�����j�+GUl���j�#EĜY�p�x�K�/�
�n��2آ[`�ն�-ǓV4-S�3y�2w}�c湳U��J~������i��i�H�Ȁ��<��;��LϞ��o�\��WmՔ5K�E�����q�}^���0�ȷS�I=�`<Vne�=9����E�9/�"i�JA�'�-N�"�e����{�����]�\��H�u����z�<3aJc���3	�K��*��N�o$f@��ݜ����m��%s(r��L���_�z��nT�{��Rg/��j-�b��xq���*#��h���f|>���nd48ƀ�c�^� �O�Ȟ��K�.�E�֮t�U�,{�lN'z�i��s�#���X�$9���g�����	,5����ܕYh��62��v�U�q��[K���e��pa7C�e�E���1G!n5 5����h~�p��]Γ�ʏ�O�����.���x��i�����V��f�^T��n���@e0���c��+��"�w!��d�5Ё_A�����}:~[���9egպ�X6������_iٮ+U����0����,htg.�۴j
 M��!ˇ�Ge�C�)�B�4�)nT�8���U��ktd�mݾ��`�z��#�����.�p�u�����
�/������aɗS�s�j���]�̼¢�g�Zz��6���D�,[UU����w7h�r�'�������ܳv��U�E��\�� ��H,�H���9����|�����v>�|�A~�S��^L�޺���H���W�}S��4L�\4���X�~�(K7�KK�����yxlC`3?��>&쎐������P�_8e8��6�{���ZǋC3/*#+0�j��g�w~�q$P�����(�\K��&�L�_�"���DJ��:��?a��J�vp����v���^��u�?���^��LV�z͜a.:k��E1߄g�~��>/&S,�\j��E�P�&=y�9�xi��U�O�����?Fcս[�M=��Ꮷ]�J��>}��u�g���c~�Ҟ�.�9���
�0L����8�b~�pg�I���Y��}��9��C�h�<�9>_@"lϣ6e9��=��	�7�&5��9(.�����ޗ�~�N{r�f�|	�qt"i���t��+�.����)�to�%�1�a�R�-;cV�+�AW�r��L6C�=�~~k��q���_A>�}Iߚ��䙮�P<�I��VKwr�tv/�Л%A�9��K��'Ѽåy���y���8F������t�8���1�˧g���o*1K��<�D��4a���ɝ�s�k�WK��٬RxCT��'b��I�Tq��1���`��E��X�Ҧ�7i�FB�{�����ꂝ��{�&�w61S���r&Z5��8�D��[�,����j���u#7�X9��M�M�)ĄA� ��M�ڻv�v�b�۫����9;{/��yjq�"&t�i��ʅ؝N�{[�i�^P�����S����Bu�K��k�F�VT��u���۔Ĳʙ�s"7h���+^�W�j+��	g�[��df�A�׎^%�o�3˓�.��=`�n�EP�T6��S�dzq���"�s���v&��=}�1�~�`�)���:�P�?�F��g��~�I\�	�+'��&�[yy�vr���L��NwU��������.�{����\RX�`г�#�����}�{��- ]hS뮢T�+?ǃ���J|���kFy��5PŶ��ꏙ��_���[��~_�+^*���=TI���^]��'6Ԃ(F��sA⯖R�0b�X\Y�~A�����4�~y�ƫ}��t^������sս��|q��!�U�����6q=�c״�.c��&���"��
m�7�^�v�hx�1�6머���[��2|�a���eMB�It�-���Ǚ�L���a��w�M]~ؒ�g2���&\�α��"�*֧� ��\M2/�H�2�y����>�)��+.j\(�Z+Z�UPxV���u#��=��q��T��cN)Sm�ܴ����/�d%�J[��{s��C9U"uc��$�p�qj�����w�j�Q�FSY!�B�/�ؾ�ט�N7k�`V��ϲacO|���ɼޏ�1�h*Ih()�?���a������a���%13�w�{#Z�|gO���6g��edY�:��Y1��7=�T���f����[�H-�L�Iw���v�c�E��?��l�@�C�e!x\���b��+���A��n�w����9���"��ʺa�@����l[LG��Bm��Pi���.�)�MA�=:�.�{	�?����ÚqsH���^b\9�#[�=��o;SpΙ6:�ֈ\���"}/��1�/��ٮ�6lB/M#�ˤ�����;�����5.�~b����0��K��wmm�2']P�������I�X�^4a��Ϛә$��K6z�D�h)�}�Y^-!����MQIi_�~�i5V��?]������b�������8�4�G>��[m�vQ�O�vb�����){`H�"�H�3�|Y5��ʀ�d�6d`�O�u�ƻl[5z~
Ʋ�����_w��i�8�CFD��^��vО<�"a[��V�:���f�Ŝ!x�Cc��T7��v���;W=k�l�;;�yA�2At]����m���ג٤&M�lH3,�{˝~��H]��������}zb\A���ZɎ0`M�`TVN��n䕜��r��M�_B�?*�wb_V��֬�V�]�Y]�J��k-.Vs�ܫ�:\T�y��{�Q�Ꜿ��z��ě�xa��////"��^^AI�5/�/��ؿ,'*o�1�ݥ��܏=]Y���J<�]�cR|�x&q@F���޸�Bl��́�O�[��bh�����G����S���q�r85����C-0`������;��%
�:��p-��sӼ`P$1؂۔D��:fG�}��'�ѐ���6���F�s�,m�)��R5� �ݬdU�>����%Ø��@`��i��{d��ϛ:n>�����7�{8T"�ó;�fv�gtCN�FuF�+�ZB+����.b�P�xG��r�}�;B�HBv{�3�u|tt#g�gOllD�E�7�QN2�m���%�k�B1`7�E��1f7{`,k�ފ6��(t�Tkv���@\\KJe��%~n�E��!��_�����p��b�̓��<��R2}:�%ι�k�`�K�nT�x��E�jm��&�E�t��{ٕqo���ԣ�;M��u�p���MC�nn@��t�"̉��L$W8oA׆4nQv��R�U�SW�u�ڞ��-=�3���D�-ZS�`!|v�㤂3}�<-W��zd^c>�<�_� ��rTh���#p;����Ӎ�w�e�ͅB���*G'q1N��SZ-f�&!eF"��L#'3!�t����Gz�T����A�?@ 	#b*�H\����TΤ$C�Lv��&�9J�[��Dg
Qީ���X3r5J2����c�N�2+9̽I�}~�SMPS�Bw��o�k��C��0����M�+�a!=��pffo=C�����1�qn"t8�WtݥE�B�o�������;�������`v�NV�No��φ�*e�}�}k/�*ǘs�;��x$$���/�d��*~#<��O�fm��Ƨ�C����1� �{�g=�9����1�%�b9ǘ� ��S�\����?N��뤝�C�:"X�_x��5.j5o:<5g��1�H�o���t2��s�D�NT����7s�pC"]�Y�PT�N��Ƌ�N�Q���"m��G�����p��䣫=�������%�3Y7�T�M־B
�ӡ�r�k�o��nsӦA��D�_�{2��}�|�˩���z�у+X� �(�܆[���hj��� B��"�J��1�zx�]��wͫ%q�=2z�U����2|�4�Mw�\PL��J�'�]�Fc�Ǽxi��ޟ6�<S�  I�F7j�E�d5Ā�>��6m)�I��Ȏlׄ�,!��n��o�����K4��#2*��~�t��g1z�����/o����������G��]wU8\��5�=��ܺuzl.���i�Ǥ�#���%N[�"lD�OFQs�p�эz�^!e\팳vwmC-�bp�8;�ފ�gn�YC*s:� }N��^ݝ�:�4L�1�#:�c�7n_���h홙.jE��g:�M���t����n�X������[���@]�y�3PB��J�\Fht(6-J����`�X\<�)����]��T�%��	<��r^�74���%V�QQM�9viJ���m�����w���+O�Mpّ֋�si}Ã�	���]?f��`���9H�Ӛ�a'���tu�,�}Z��[\+hK��LԽ]�к��v�;���j�RO��u����w�������ՖR�[�=�uf֞Ye�\I�B��N6��&(�1Γ��ۃs,ޙ��a���7x`���Y5^��\�k�f�5��x���'Y����o�����)���U����Kd����;�7Cv�컢�Z%ܪt�}#�sss�+Eݭ:H�i��>{s����d[s1�	����r��AN|���Bɺ��&�	V+5Z�<�\��DP�SU�0o\�ufL&J�Ň��ڮd������,c�-�K���Im
���`�ْ�y�"���*0�^��喴��9>�@�[Z���#������-�9L؉��"Z�rH���dL�x����I�>��.���a\v�mF	"o�f�d�Ck�J��лC�r�U<�m)tvI�*�m����(y��u��l������N�LS��6T�Ҷ���MiosN�޺ҁ/j"�2�9ۚ:�6�d�;m ��[���F<��rns�ۋ�[��4�+e]i[uH�S�̭�^�G��.��屮�ͽ��]�;;hj�U_:V�Bx�2	���
��NxT��Qe,�ԍ���n�jw#V��L�Oa�
��4�+��H�)�'S��[lt��ۧw�+���Q)��v�LE��2�d9�s��AP�i�)dm�\�a�-d\(�m��W{�Jc#���1kq)@7mA7�v����ȏh'�p���+�.��T��Ux��^L@����>�u������f<�e=�L%-�fe�W��쬪��I�Fag�&�y0X<&��t����"�
���5
W[I-UX�����ß�ia��Vٙ�ɗ�2c00�M;�f�;�W�Qyuu�L{���K�;h�M�̡V˵���U���T�w����2m�#q`v�>������ݴ�U,�vTJ��**n)B�JYj��k���,Ԇ,ygn�/VU����#3J�MJRЕK�F��H�U�Ku���;,]o�΀�����ݢ�_�!
(:����p���.D�O�~�S��nl���00"�L�I&����m������H�i�G!h�Xl��HE2�L92[�D����Mv��W)X5P�D��R�ae����B
��7\��ܘ&y}�s���옱�la#T`!D�Y�$2�)�N�v��o�Ǐ<x���ő	$BFBA���F���M۷���q㷯<x��ׯ{	j��bE�o����(��E	M1�q�x��Ǐ<x�ͯl��sB�h�sn5	$+�Q�Tj�i�}qǎ޼x��Ǐ\2$����P
��ܒ��e)"ӻ�r�����ML�7�QrF��
�\'��Z.]FŢŬk��k��c%�fDDj.j�cs~]�5�b�QU�]���hM)o;�i��<VZʮk�[���EA�5�j�t�,�$x@Dv��� ��s��xm^�V5��;����io3ו}\�(��ʫ�Zf�hgj�e�)m�\g��e���ޠSd�
�o��D)��{~�^�Y��4�1#*D���}�_��䩼�`M����)I�Ԙ�/�-�cX~��\޶3���E�sıN�������VKwPl���|�.�%�d����3*\!ZD���2B��E�DF�ʇ������t��"*��W54SWA���eN��r��^�4 ���kz��m��k���s�����w	����/��E�-��~W����(�_t��s!~:`����>:��Sj=�i�L�6�g�vJ�/K#X�R;�����N���dD���Xrk;��0��[0N^`�\��ljdK)7k�V��Х�z�>W�S#(_��q���$k�|��ܬ���� ������~��G�����9j
�G�{���=�M�L�' ���i�CF5��;y��
͍AS��<2�63�
����}l0��>�� ��}ј6'�>�G;��Įo�Lg���|�m}8�
g�P�7�1��8l��)��)F�/��d�3�n��۔�	��i�7v49Gb��j�`S@$���_E��b*����]�=Xa�2�c�_���'P���Т�\������PS~�xR�U5B.j���UN�nB{5a,b*)�b��H&�Y��n�Ȳ�r�՘���9|�!v�#f�fW��|���'w�1�սw]L�W�S-ot֑zۅ2.Mj0��#�y�.�����Z�cϨ�ߕ�\B�7O��O��yqBkvS	�n���jP��*��@�)��4�;���7�Yf���_��7������c��P��A��7�ZK����������f�=<{����e퓏����0��y�\zy�5���Jk��R��:��v�w�/~J�(�x�xH\_V^-�����_�����v"X�.z�J'�$?r��E��n�.".+�K.u��b&�e�+ᵰvW�J��W�lt���1�M� �:G�t�|D�r0R��zl�]R�Ѕ^�]hWSȴۥ:��Ja��FSSdnH�z�X:�<�c#�#ޭ(T`+�b��CȢ�\G��1E�"*��g�{�]�j
�ʨ}_�𮜐��Ѥ����u~n�F�U�9�z/����ۇ(���<��&2�$��됥�zk�>@�^�C�^�1��qxOȁ�����7���(�;�~���O,~HM�]�'c�s��)�C�fY�;����3q%���N�J��9>�;K����O�����,���9ko¬�7��>����+~=�W��b������/�>��3�ӑ��晴�s;(;܊[�nQk�n��὇���y��]V��3D6-�i���7��OPOf��1)�7�#v���ՒВ��J�I^�
*���Q�KZ����«hQ[��Z�u�7|��\�)L�c����W�x�||���G=���Ki�S��n"��c�gд��~�S��!�O�Qiα�B��_�:���(�=�T�1&�u<�s���Ar�U3����t�0�nɆ�;�M�4l��d^e�?Kr8���x/s��wJvN~/�L(qh��=��tu�<P��F�1�D�lzC�>�0��R�kS�m�����&��3`Z��G�|�!�0t�ޘ+��!lXp�N��*!��5yg�iۘ�귞g'� $1�'�2Y�5=��}=7"		�B�c�Y�(7.�l�9a<$���iZ~1ӣ}7��X��{8�� Dd�{��L�h�ռ$�=��	���'8RAl�Z��^�x��S8�C1�>&-�q��>�{�� ��6��O����Pq��{��l{����
t@�����]���鯫X[���?1��~|	�<C�޻�hVy6�_h�l]�7����c�'� ���HE۫+���'����T���������8g5�{|*�m*U��Ŋ~llwL���$��#� P��~���$nE�*��o0��Is���S���+7ATۦ�u�u#}s��}��V����t��S�^��YoVm�������z��_[��V-˘�wk����j����#F���;�W9���΁+6�-���}Hi��;�LV��n�(m��.AԲ����"�i��c�1G����ٝ��|��ɷQ��=`�f�1���ܦE�&�t��Q��νb���k�Թ�8�1�8\������˪1��-V�F���S��S"��Zx��M�e�Fә���}�G�ސԎ����x� ��@P���?th>�U;A�
���Og��YK^`J��,j;���vҪs�!��7�ԍ��-!ږ"E��e�:��z�������W{�G�Fț���,U{�����>�>$�[F*�XJ{mniwƶ��BZ��5�˗��f�Y��]86V-���dVW�9���	2��%픿0O�u�c��!��G�|��b��7���5�U�6f͋T��x$�aV���Ctڥs#zEZ�4;�'�v�� G�"x�^�?I������;~�QB�0���7�����K���s�X���'䡛��x�u4j9����d}о �1.^M��B��311�B�C�J,���,���dr�����(Ӧ�ma#GG"�@d3�'D\GS�]�>1'�����1���+�Ep�s\!��ޏ��s�h�L���i��4sK3mJ�b%"�!R-�f%O_iG�}�Y:�c˻w��1А�T�R�����A�D���~�[m��539}=vl�W޺�t�Efi�h+�2��yq.�YZ`��e��1y"��rS�:�����������f>O,!h�ma�4��P��a�����1�ey�w9��+]2�8n�Q,���OC�*�}�t0*U^`�26�Z���g>�6��C�=�6��O����攽����Z��c����`��U�=�CB��_G�;8����^��P.�Ժ���1>,����gZ6����p���%�6���κ�]��-v4�L���/C���l7�17Q��t��\C���<��x�X=<dEdA4p��Ŕ>!��I��O5oD�IBa��!x|�������<�M�dL�́-YE�w����v*��A��XxK���O�w��0�W\c�����|?C��׆ߗ����7S�B�G@m
�F�>�2HR/�����J��o<�u�y�����r5�_�Y�
����-N��ޛ)8���"�	�HM�P����677�5(��k��|g�������ƽܜS;�PN%��솏_�XBmh�uRܢ��`�K+�#�z[�3>Ze��"\	��|`[/x��fz
�/Adk��祐9�K�{r��V<�=�c0��'�ȏБo�-$>�ڨ���?�vqyJ׿r�^��֮�D&t4�`����Q(�׌��ϫag�6eGB2%lĵS@�,\�4w��E�ŋ)-d꣼��j��2���Ut5�_ZUזϬ*8gRMҷ9�d���b�I�[�s	R%����,�ʹ��3M^��mk~nj��sfìcČ>�ߝ�9�|�SkX}�P3�
 C�z�	��L�T'�Q�3�C�zwW�p�<>�eW-��}�Q�
w�D��8+�����G�}�;�K�|���qY(���G�eN\���.�B=돀f(q��F��
�Ǩ%��磐��
�x�����M6^�,��,��*�˱��w�D��w�a�`��8�>$�4�1�]P���^�0���=�W�>�!U�<	��ЦI�mR����Vמ���#�ByP೫jd;�ѦTI��(�
-�G!�,�����˞е=3��縼�/1�O4��u*�2�%8��-��yv��r����q�[��]ZFS�@ȉ�W߆AI0,!eد>�A���x}�� \Bj����A�E�����K-ԭ�����+��">{.�'
\�E8'�yk{,.}<��HU�S͞��ޔ��m���Z�w�B��<ڮ`Fi��Q�Tu�5{gOT�C����\\:!�nO�n���P��{_�9�}����~w��T��.4���{�B�c�˩��Ϟ��2����b�B�l�̦(����BP�Wx�
�Ar亅]onPyoVb���c���d�jJ�#�(����OtĢ����2�_�]�4ma�n��O^A+.2�N@C,�3q{�9��"�.�V8e��wMh��������o7���}��^���mC1�c��;��ԩ'�Қ���7U�`�b�sxO9/e�cC�[��;�4������_h���M��p��V�{v��P�8ŧ�k�=4�uПYL:�������t�_���0������3�,��OD����~�o����+�$&2�?oG=d�;&������Ve�<�S˼r��;`���K�&(��=����~Ξ�k��I�L[9��F�R�[X#��V"�7��O�랿A�t*���{���D3���������}l�{4-7u�*��
L�U���j,
`mǿ�,+����e�Oi���D�\�������2�z���hkպ���L��-�ބvF�!�#qw- ���WC�����b�3,�U�Ю��~�����N�爴��3�ͪ�F�kS�m8��1]�郦��f�+c
1�N��=εf_V ��hc����t����zh�Rhdy�뫼�k��X���4��ϑb�;�<rZ$�����^_�Cj�[�nml���	bN�L"�����h�S�.4�F�6����2��E�+}W4�6�%Wl;k0�d^���sKQ8R�TϠ^Y�Z1���!�^HB!SɢG*�$���s^k5�l�ӗ���	���;��Ƅ��NPJ.1x�8N"Q�S��IUE����Үy2��^yy^�[ߙ~���c��{�����$�>u��6l]��21��}�N�>B�/ܣWj��l}���E��n�Ka�����;��5Z��z�X��.m�7/%եWϱ	�^��������-�s�#)��̋���oc6-f�af����>p������|W���]�T.5C�wq�Le�Y]������\��7�N�=n���6۰؄�m�w����`���[�[#���B'mV�B�:]n�4f��_���s�0�, ������6kʤƹ�Ht	/��45�A�,*T�]>J�t�h�S��ռ�����y��.>��r��g���vܘ���)�W�r�]�3���	؞�#��S=Zi�'�]þ�;��ڀO��=z]7Y����
YX�&��Gz���i�;s���,cڍ;My�����:�j�Cg�A�kSc��w��@JS��晕�k.J��Y��q�f1<0krTXW��N?�~�(�?$p�*I�L!�g(!���uY���}V����Ay��l�Z�J���}��&=��Hl����v]"�F��"�����b-�Ka�7P�:ݺd��-6�{�z�m �Ra0���nU�Us���j0g�.QI���L�bl遵bٍ�����>m�����x�`�>s뵵{3
5�L�T����k�_Lw[���X�y�K��Q2�	�����"e��헢��0�Z2HR���Y���[����1�c��9޸�܆�"�g�d�q���1B �jx�7��y���F]oFs܆���1�tS��v،�Q�j~���П��(p��.{���-�%9�댟�=�5ΩM���%�0����hO���ǐ4L=r
HoE7W���5��x�#�O��|����"��D ��7�����v ~;�����5S���C��*;�N��]���~1'���.���~��znL�ϗ���,��-G)nǽs�{���\�)�pk�o�>�ۼ��p��2a]�kj�h{�d�2�*���U�uKТH���7:����[�9,~��뾵B��0,m�*{<���Hw�Ю]�Y�Mam�cB�h�Ƙq�^�9g�}B�x�M��P�V�T�*�M#�=��eڌ���f�z�+/���.�S�;F�i	���� "����S{�� �����J��1{��(=�U��/3���u��T������o��㋈��@��틴������.�
�~�����L�>\1OT@+(1hv�m�X�)�i0�����1���ݙ�	���Z}������%�Qay�s5�U��ݓ�K3;4�=(�r��el0�Vк��H9؈7Թ���N�u��t�#�5QY ��b-��A�� �ϼ���G��m!/hiY�˻*�����4k��:%T%m�;��Ѵs��b���K�|.o��=&L�S��1�����p�s�����w*��8aƧ|�-c*�C�6����Y�?H��|s��Ǜ�fJJ�'
�/��YB��L�ʾ>�w/�OK�qq6���w�=��.���h;��.������>��ʰ��gB��^���`!�hLsk�ey��� ˬx���*���6��;�t�lir̗Ewv�ޜbC���\>뚺a4خe�Y?t��R��%�*3� Q�b�c�\=�,�A�'C5oំ;>��K��2D��L�K��B`�qAa�Q�'<���8<��T|ԭs%}��Ϫ���ط�*�B"Pp�]�[��$��y��Gey�F6���C?��`�F���Y�ih�_nGJ��SsQ p:E��p�˰_(��X��$�XO�߄�m܀�[4��'�qh@$�5��ٵ[wM5��Q�΅0]�����;�����0h�G�����5��'�C�����H��&�I"�I+5jS~>��"ϤW�������D�%c|���6>uA�EO����.=8� �T���;!���af����0Oc4KU��Q<Ct��M����ʭ�-�=���r�s�g�ֶ�9�9����Q�86�[�Ƀ,�g�[�:�|�c(�}�6�Ky�b��!]���G�%=����vÚ�F���3m�+z1�����n�j�.Q�ک,b�aV�,�S���r3H�si�����TW}�iV8;��&{}9�W���v��h����[�wCkۭ��rl�b��5*�73�˫J9�j��-[AFf<h��c�-�̢���K\ڵ�����~�S����=��u*ْк3���5�1������^ߙ�����_:O�;a9���|ܐ-{r�G%[��Y�Ѥ�,����u�}5!�uM�Z��e骻Z��j	�7�������$��Dd��N��vnĝ�bj�ڷ)j�|j�l�&���54�â�[���V������Gv�9=���R���YN�J�Ϋ����J�x�������hu_V.Qv�ܤ��zy��{��ON�Ke.ԝ���ݜa*u�n���Z�3I�z�|K"����A���M���~�d���*��H�aR޸�^n9�J���M̳	%9Ř��9M��;Um�����#N��-��˶S��ө�J5�݄�0���K�8�q��ċu޺��t^�S��d�`P�n�ڗ�K�0u]���9Sy.��Փ��T��|�L}Hg#���l�D�`*��7���o�å�� �<��sV(�[��DF��	���X�4��1-�,�3w�>�Ufb��(N�Ρ���{��m�yn�"OQ��+��<!�Q��\�-���/0��A��c�{��n�.��T�Q��cQVu��霤C,$5��E�s��Ώ�9�r{]#5����K�ŇuG��
uڙVGV#�W[d%�*�!�eNif��S"�}�yЛ~�͸�M)rN���J31lW[��tJ݊����z7	��{k�5u{��.:ю�,�u���3�7n�Ju^�W��Y�-���)�!�N��uKi56ԊS�;z/vƩ��5�'5)����n=�A5��%u�Tb��vE�ݜ�c�6N~�DX���x���=YRŦP�7kG>���.�%m.�R�[v�AR��ծJv0�*�P�ܮ�W��+_gV¸�MtI��ܸ��{7LÃj�ۭ���mѡ�s�
dY�ɦI���g&����Z����>�؉�yA�}Yy+N���-�+����{uf،k
���{�ܢF�m�̱֘��6�Ml4
�o6vr�I7q�
��C�Vٔ����T���T����&�V-���yR���Z�����\�P84�2������,���E�|�x�S�]����/vV*�o���]���F�n�X�bk"R��7�E�3�n����^2 I! $��P
��*��&��s��n�ݼ�����;q�Ǐ<z�E�J�I����F˜E��j*,cM8�8�ǎ޼x��ǯ��-�n�5sn9�ss����M���p��nݾo�qǏ�x��Ǐ\\'a%BBB9���u��m$�7ǉ�swukTjIH��Li�N>8�Ǐ�x��Ǐ\{�IQM@$��*P�wtl]5�yU�W��sQUӔ��βn�WwF����<��?ͼ&�����ۺ�p�k�t���T;���71�������\�wr�����}�c�乢�ww�W�sb��,n^���;b�p�wqwcN���\#[��wmr1��4��.��=����ܣ�^��_6����Ce�k�q��k�z��{��p$��a�ÚP҄ �\���ʔ�H��x������s2��̻_w�]�+�����-�7'�`��T�����b�I���Aݧ�z�M�1:��yc���U|kXX�y�
�V��V��`~��_	Dw���£��$b�j�ؒ�#Rz�uS؅O��<D�����+
�
��}kr��)�V��D�OD��Z��؇#2��2<��9KiF�	E�4t9d^�$�'B�R3�퀁���p� H��64��7ʩa�y�������]{��©K/H�m�s�{����$�Bb��E*��5�1�#$4>K`�I�����`�cǙȋ<��rC�'�A#�$
���:/֢�)��\�6�u�6;^)<]����B�B>�j�D��祆��i��\�ڽT*��ҹ���	��u �^���s��s܋_�-�}��(�~��x��c��B������#9t�w�u	��-df����Q�j4����a\�fUHǡ�n��a�8e��%�����}l�]�6'��j��gsORZ�b��X��=>�g[�)�z�"� �(p�R��k~EJ6�����3�2��a��5y0.�n�mS�Z�p~�r�Ϳ�����:��=�d��J�I�˝r�Ս�6~o������15�WYV�Mf�Dڂ��ד[p�V0�zlۗ�h�D�`N��-�ĵ[�s��r�˼�=�����1��3̭|ϐ���Y�������[��,Զ��Om�h*� !�dk]��&�6\�C�>dND�y�N߯o��Mcױ���=	&e�����\÷7#�$>��������qwa'WTW�g5c�Ǽ`o�V<Γ��kA�?}�'�+!1V#�&�M10y��Ӝ}���&����Pj�����4���ʙ�ᨌ�Ԁv_8e�!�N'�P>��2*�%�0��}���T]?[��o��WLګF�����J}�CSe�pe�1���{ m�d\?Zz��5�G�?`_�F��A�m���Lx�Q���h��\��`ڥ���|k�ז@�4��r�n2�*��ft�X�.%Z�O��(�Ju׵�[៮g����{<w��E
�ז�����ꋇ�{g0�)H��c�yʷ�U�;ym�U��ۘ��t�ב	����:��
qOql!㹌gP�%v�x'1kE�sO�6kߗ|���@��?������0Ҩ��x���"���BK'�9�x*�^����Fʸ*�"�����\Q�������0�ވ��;�ʔWu~��`E�*�l���$����d�bST�]�3�k}ϙ7����Z��P{l'� T�*���670�r��6h\�s2MQˆt����/۲�U(��\鎸j�}�w	�r�vD�*L5b��/���m6�sB�[��"�k��8�)^u'H�I��G����9<�@��F��:>��Ņέ�"�F���}�$Tx��+R�k}N/[З�\��;��XXA�xj���\�7�.��P�]�^C۳��]�m�̈�&bgM�]���d��4�d����%Ů��T�u������@c�\"�{q4F
��V�����X�ݚN"=%��(���A��W\ܴ���K�g� i8c_,/b�7���'s�����<��O���>�$F�T�6�*�,Y�R��!ˎ�ǰ���f��ń�����%V6����V��B
z���cY��A@���TTӍ�'���g�a��ArN))�H/�3a�w�'h�Y[�+���D����+���D��hY�F}�*Y�1tH}���>�>O�o����sB]#��0n=��n�S�u{3�"�0%�s� D�*|B���;��KY�^\A��;ju�f}/2���_p-��5?z����%r�My��]6y�mM����"�E�Rg�:Ϸ�N�#�z���ۑG*�澰`�b9�5������4X��&�*��s�ҥ5�(��fݥ�vT�X؟�1�l�}�>ۣ�@fc��8�R�"�d}�Ҿ�ccG�y�dQ�]�#�կܩ��WU�<�Cq��f�S;��%�=�7t��**����(��j��ʦ�u��C�Y,�����ޔ��>>?���;�ۄ����,�X���#��2W���+F�w�#�,R%<-���'��|U#�oj��mз�xn���#�<3����O��=���V#��Jt�-5bjp��_���XK-�`�����;��@JX�Y��~�2DO�'�����z5_�+۷��m�eu�ֹ�s�|�xm.��Lk�L(>��(+��#����5�I�i�ep;{tҫ��
Q���݂��2u���^S�ʥT��)�{�E.[�ř�c�� ��,+Tq�����?lɿHR�v�H-�i�*��Z�$_)�z�����5�K�5'����4v:�;Օ�Ovm���z� g�O�-5��́�i��^��z�%Kx�+p1�W�����4�:8���;�"*ֻ�	0���R��y�:��xmXXHfO�<�r��eA/uf��MF��6�,�����|�\_;#�֊{�0��Q���G<���<���T6{Bz�����[��D�m�F}8�3����@��A��F��G?y��Iݹ�<3k������lۛ�z��Ƿ�0�y��l����!����(����,�㵢Ԙ޽�m>'2�$̥�]���ɦXD�
��C#�V�EQW�5��@��sU��N��-تٔ��9]I���ZWd��TW��Z�B̫�9��|4B��1�g5�}�;�}����f_,�U����7�͹]������u�v�xw��@��
�l&qss�+jW��}����5E�[xCn�/��Z$�z�^a@t�Ú�ϥ�������Ѻ�	>��0x�E���s�"��ޡK��P�:ul@�r�XXu5�}��v��:~9>{��<�������F���l�OS�o)��P*m�d6��V�@�7(+��`%�x0�o8_]�ꭁ���֖*�8>��C�L0��Mz��h�:�%5�s�x��m����iR7y�ϯ�|�_v��t���8N'�8%���@ n,�
��@�����CDW�W�3IZ�Kׇ:����T`IM5ߕ���񹩝>SۼH0ТS���;�YFE��F�T�{.���~wL��DIu~*[�Lh$i5��ܑ=�p�G�����'2�+E��Z%d �~|���m����.�'.���7泔S�5�
�?�/o���>%]ys��΅A�8П�� �И>!��S�j�i��E�q�O��G������<�'X긁UuOɡi������'Yھ���KZ.@f1��F#������(CvVUêT�U��1��d��>� 2�u��Xkh�Oi�1K������e�����MV��|c�Т��M(꒵'����'s�Y��}�������U��g2XϘ�3L'T�h�yf��KD9!��Ρ�_���z�Z��W<��k�����a��%�]i���;����яp���7�o�k�t�bk�q��ډ�̦��;{+w ���MH$���z�O'�\�=!]��u����C/8���q�7�'ѽ�� �����+L��2+�����e�ǣ�b1�<�q�P�8�I��܉Ə-���[B����)|d^��}ѕ;l��C}��2�K�6���˱����zw�H�>��B�c���ƍ��>�;@��!��[b0�@|Ź�I����O�:pl|��//��g��pm��_{c�\2�0�p!���*Q���^�V�s
�{�=�b����Kr@ߖqc���Gㆹ`�-?�`%`��I�;"���#0�MǦ}QLjK�1��n{a:�������41b�46����oE[�����x�`Xd��=��6�i�Y��;��`�!Ҽ��lq|k�l ��&:�V�ю�0�\3b	�\4��5W	�8e��ܵt7H�_ri[݂�s�;ܠ��
7���+�_z���L>֍axյ�s}'Ɲ#J���ʰt��dP�`,Ŧ-�S��85`���)T�5�oH�SR�oulJ�,e�}�]2�#3'+�7�."m���z���:����~�������ѫ2Z"Jb����gg�x�Yó�Ǿȶ-���b`=��ґ*�	O>N7S�<ʝ|�{�=�Qv��d\Ά-�����|�#��!7s�F�i:�IP@T))��K4S�4��]����Ɣ[Gtc{$=�.R�ò�`�~�E��l�1�� �Y���)����۩�)P5�q���#i�!�I3 @ �4�'� �y�H��)���ޛ����/��;�u��M��7@M8��m��f�n�N샌�?&C$�/LWq��<�h������$ԷgXM��<��f��|*1�U�p�	��_�b)U2�/Z_,�(����ۿ�i/�OH3�<_���IaKcX�WZG�8ll(�4 9�P���:=jz���!�2�6Q���a�?>������'�k�PK�)~j�iܜ��FM5�<ONa����g$�D�f��U�#�@��C� �K���^aٕϪy�h�p����k߀�NQ�c�T�]H�ǻV�Ě�L���ksHgV6C3�A��01�o�z>�ӂ[�W���h�5��04�����Hf��{˃����S��E�kr}x�3��qͧ��>�����WЃ�pB��Nr��I%�q�4�'��In�J[,F�s�	l�I
MV���&���k�@�Rj�uVVh����F�(���ln��w~���+Ђ�>���z=�G��w5�������6V�Ů�L�!���1äFb� ϡ�r�}�lQ���Nus�����]�$.����H�x`;�	�TJ��n�!��U�&wx����I�<�|j}}��U��/Ug5�Q�P�e���-���/A+��y^k|�T<=���e�Y�Yƥt��v��ل�'B�`~�-|����b�������<W���o7X��^hތaH��U�4gaͭ��z[�a�<��-��/K3�~t��om{zK0�׃��dޯ,R):\Y�z9�����t��s^!���M|��:=�I� ��^s��-F����gp2��W��2�7/,p�D�d̍���}ZG5B*�����S:~�=�ćɑ|ɀ�υ�w���8��o�Ӝ��9���<޿g<K�:��KL�QI�͢e�eO����.�"��)�������{\�mHm^ܑ�s�0��)>0�0���n�c��p`ۖ��^"�xI�[��t���F.|�
��Dq�|h�r���B�z�);��g��q�O�iAc^�%�J��(��P{>r�b;�:Q�q�E�o[���eu�i�M\��s��X����Y�%.��}(�γ��Ot��8�F���ec�Uku{��j�hP��C�Flxx���oZ���|��'�K���ɺ���4�c�3�	���][q�2���G1�0���* Lsi��4�k%*T�u�@jvU~�W<�`o�{�r���i�^j�p���;2}���#���X���<6��cv��w)Z�K�������[�P�[OR�n���m��a���@hƠ�M�Ö}*�"�f���������u���]�=��Lc5��r_[��s�g=�OH=���|�Xs��R��	��=�O�pܢkH�8� ����c4ǉu�}���P&���353��z��j�����fI</�+���^k��qk^l
�J��w���u�t���w1���8���	��UEoc��X_�?]���gO~Z"�U����u�&lt���#Lk��xT���*Ewu��j-ǳ#�)Ě��b���kEA�^
=�뫘�sȧ�:���C(k}�n��N��`�	e�zv��i�kyچ=�z��
!�@0c����2;����{�[%�1�+m���xmAt�څ��.��ߺar�#�W����o��2`p�� {�n*Mj��w˝���C�]�MUˈSV��� ������M�(����j�M�/ȧYK/L�$�sj������W}�WUn3�j���B�k� �uf��]�'��N���h�����xN�j�D�+�ъ+�h�wxpͥ�	��J��8�j��h�:o;�DT��WU����r9s�����}�)���I«e�U���\Y[Ǣ�8���&��fT�MZl�j��)��+`p�50���Ľ�����R)�$i5���싇OF��ж(M�T�u��%�f��x����<��������k�@)��_$�sz}I>��Xn��X����ޛ���U�WR&v�Z���%�uxظp�y���ׄ|�,�!?*o茴�*�����rO��4�$ơ-4Z�/�� �at�vC���r��S���;%P��RЃ�粮��3��r2���?��
��	ܿHm���dF~#XVO�sס�y����{���h����uaWX������i�mHW[#��<��i|���G�����ј��g_\����|p>���Y�,�/1�(ݕ5�0:-f�m�W����G��9�m֤�� c�E5c31d��l@j
E��.����}���P�}�ߡ�]�+��l�m$x0���.6r����f6�M��6׋�ܝ�:�1<�/�P;�ǥ@lo7u8� �!���mF/őF\�+J�@�'b�W�RɘF�j�f%iØ�B�u�+z^�݀��|��'���a�4�wP��Z��/E��E3�V��ÍZ�s;��ZU�9��i�����^�Q�6ow��f;��Ѓ�:�v�uL���̬��OTm�떴a�W��w����R��d^I����J2��I�&�������UZe���Ӝe����VW<��̷/�!���OnU�:��� kt�)�K��2f�Ւ	�R��0c�S�orw�R!�D�J%cԬ;�OB�P��#-���f[H3�:+��f�[}w���Q�E��ܼ��%A�\�fJ�ي�-}V+2,��>��ݥY�{����L(YT���[:+�|��
��T�vȻ��l'$b���F*�A�ě�L�RR�eE��^i[�>M�t��x��a�n���N�Ԫ�*r��[�]��nuI��ҦƲ�����)��YR�`�G+��5�d��l�Vc�k�����Wv�R[/�����zf���[��^%�[�%�{��m6m�Ԕ7�$��٦6>��ZCf'سfn��uG4���T���s1U�rɬ
b��w=:�p�����S4�llЦ�y)U�J�U��)oK�[����U�9���][C8�=lghV[�F�N�,]*Z��1h��۷M��y��kT����pn�)h����sJ4K{��{Z�ا8��:��i�l�n�"�i;u+�f�έ�"
.����e-���Ob�-n��z��Өu&���u�7u����s������಴��َ__]���z^����Nin�R����5��,f YOOU������Xu:�mݝ��D�fcK�39-UPd,m�p�Xw��rΗԳ�v71J��O�)��I���٥NU0�I�!u�4p={�$YD���"��{+�ˊH6�y��[�۔[	'R���5���*���^|��ԒVR)t���z
WU�Z}��ʨ�/h��P��{}�h����[�C��O�{;T�� �����uƹ;;�R�{D�ɓ��4-�	yzp0E�:�b۩�w�޺��'Z٥�i��w-(��\�4�ٱWfI�{��Q/8J8d�+V�q����V�=���k_6�����lyդZ�T3����C ��w:�q���L�d`�3���V^uY�	��M�3���y��ך]VS�TXy֥�ј�+9�6��E���'����b`GB�1Ր_R�0�(�
̽�!	b$^��i</ie�n�I�Y���&ܭ�8��V��bʼ��V���ڜoXۤ7��B�;1���a�[NS�%J�0���Aۃ�:P,���.�'M��饝E������[v�z���e�W*�8�4#v��J,B#B��6��$Q@��>�(S��s�U2Ij�@���웪0,�Fêm"��(�Hc,��Y��mp��Q�l�C��5��wA,L�a�G`˕n�L�C�Z�;����ё
�Nnl�%��?��nX�.W(�ƚq��n8���Ǐ<z�����}��kӕwn])�2U3T4Ɵ8�x��׏<x�{��39h�ᱫ�x��P�j��1�=t�8�Ǐ�x��Ǯt�T	�(�)R���FF��RTjT	R��i맮8�<v��Ǐ�bH��@��$�RS�����&H��r�� �s]�N�#��������ƊM���痗9Fx睹�D/��9-����t�3BQI�nvs$.�]��e�۔Q�[��9&(���b���]�뮼;�����>ן�цY�i/�4H\ɍ�t��K�[��QDE��;�B��Z�@C.��h��{�:V�	�mA�/E!�X�P�8�e�4��k7*��m3p��m0n�Ğ
0�DeJ�]��M�T8a�z��^�	)��"bGLJ�@�����������\��%�H�����U�_S���/ʪC���!�_��G��~��]Ơ�Me�!;�T����ME�߰:��^9��D�x>��>�]�v������_[�H�h.:������J\*張S���d#dF�n�u�c/4�L�asK�Ϛ~����w���o��\��`e\���l����ٯ`r�W�$�
��_uغ�}�8��D�T^�yW��cl�L�����k�����ٸ�O���sv#<����{���	�ʜ5M��oU�=3Y7���);o�;}^ݫ�)[��[�����6R4����5�Y�ՓI����lm��s9�oC-n��ڊ��o:�b�]�f�e]�͎#�ќ��{�ڕk�l���A��5���PP��,�hYxך�n0�E�o&�Q���j��.�:&!���D��	fx:_eR��f��	`��&C�u'��ru�rk��C���h�x��7�ch�d�s�-9��(��}m��Z���Yn��:.d3��{�K����K�c]�iβ��KeÕ����E��LݣKɲ�$WQ_�����}2y��y��o7����ZQUέh�����;Ƿ�OG_�\�Z�QJ�d���^e�	�OM�SKDj�L���`{�hwl����Oj���IO[��h�[Gq�k͍���g�	�0����Ѐ���5}���y�@�C׳�E�(�S��8���cCh-�uy��uH*~a5��ǓU��=&<;�x��{~Eg���������h�g�gTUD�-C���/]��.^��C|-�]<^?��c0jb��i�f����~@ϥA�ʝBx^Ţ�b�9����7����犅Uuk�kT��Gn��I�Ȯ�x����4�b{^�}�_�u�5 �z!��]jT��y
��O�y9�r�Gl9�ɚ�5���=���}�Ng���U��'�p�*�NqI��
JA0�/Uۃ��2�t��m5i�� �j��ܙ
ȁK[r6%<U�>��ɭ^Ii��f�Iƺ��e�N�nufE�%�����k�V���������mD��-�PuPN5��55��V@����`��Ͷo;8�{��a�qs=+g76��튷��Z/FY�Z1�ɬ*������m�c�1�k��xy�1��o}�6��-UA�fP�k�����u�����9�s�<P�ͼ�֞�|��P7��|�[ʂ���A���@>Y�*,e���	�5Ƶ�MU�y=n�B����h�l��k�H��t�4-mwO`b�Ov�֝W�8��h�Z����۔�}5�&�k�؎����CQn��y-�2���|��Z�*����WG���w�-�_u����iuۊ��g]�"rJs��c�W���FM3��pv}���૯�#�}BA-���a����}ٻ(�Sb�?�W/��V����R^��0@�C�ޘo6Xgvl,�<L�D��\�����%�/ܽ��gp������6�s8���!*���E	����7Ud��"�dz��[���;'v��]�(�4t}g����J���O |����_�A��X�ot��s1����.��͸�Tݫ�"2�n'P�D�r�B%�A��ٕxiΕ�̊Q%��������o�<iT�
6�\�.��,��� ���ֳZQg��0��n_i�؜Xndo��ʻm�Y����7�=5�o*�Q��=�BO_�1�c����53]2��_|��6�4@(���R�E�5;xz|��>_c��,��᪩��p7���3.�%���Q�GT����C�e&�]����q�î���?�9�b���u�fڹe{,��=�*}ّ�ZOe��<�)0�n���\�$���������;n���$r�R���sx�P�ev[�F�ٓx��-��&�R�T��|���n����3X���ə�UVٳ]��9���{"=b�E�ps�T8���EU��#kcn�DkJ���z�{~ȺN6�~���l:�g�3�^���Nz�[��uc��]�ͨc-,���z�u�{��)�H�;=��,S���Yܢ�;.�S��=.ʎ��>���갆��['�}Ka���04����7�[>�I����'��*ާU<K�o����w�f�<]��mk7X-��M\��;�J�YR���j�L��ݦ5EɜVhM��f!*H]���(֊;Tejyq��{�F�y�9k����"��\�dl�K�V�F艗��y��0d��Z� TO)p���J'5�t4�������g�9"��.��Hq$@�ꪪhU��$��{��������������M:�)�~��I
[�(PVH�l�zH�n���*V�c!�!�YR{D��H�룸�J_'�^����Y̑���ه&s)꧍4)�$5��
�`n>I�C�C;=񁀺��U��5}�<r��jW#P����ѡnJ���dK�����5�zp�^��+�ϻ`����LȼQ��}���A$n3�c?`�#�'��Lw������Y��Y�3�H�T��2��q.�p\�����{��c�B�<�o�a�zn:&o2�ֲ�r�e�\�H�)�d]�G�)O,�F[q�!)�۹�=���W4׮R�g)��A*�q��<Oe����~,R��TF̫��W�����q7�G��2�`�|�^�q���q2�8��JK'�5;ۂ����i�r&��Q�&��W�o�+���֚_��d�S���"�Bsc[;oq:Qb�j��p�I����Z��OX�b��@�f�'t���N�|W�`�����S6���ڦ����QxnRuw��{���s��.��{��(^)j1�	�$�Cz���9�u�����o7�ߏ���D吡?<G�|;!z�21�V�����t7"U�.�"��@	f��nH����:�A�
�6�07k�?j~U2�ل�hʩ��?[|�A]��6玘MĆԭsn����']�4y�9��o�V�@j��_aO\�#[�}{5�X .�y���Wt��Iڼ;3��b�S�����d�[a��B#��-�]���B�q�U��oH7�_X���$�Wb=��[cdɘpFpp������FL��d���Ǻ�U�{�3=�W��.��q$9������3��1g�'̮E�Թ��c��ֈ��&�6�_gO-��>U�~^�Dc=�!B���=�p��-�^^j�DI����@�o�f9���L��{N>���]
�f�z��-:A�\Ѱf;��S�YB�&DTQ��[�w|��e)���Xt�hK�=�{��Jj$j�g��ܤ�k�U*��Vf���v#%ll5��,܇-��غ� ���P7��qՅ�(�"��@G.����D�g+$��ݡ��w��2����KN>�b<���t�n^s��;m\�ʮ�컯5~�9u<ԕ�?�1�s/;��N���|�YW�M*�M>٥�_{kF��w&QE2��I���1��.fQ:+b�{�4!�&_��onp2n=|*��FaGo+xrk���R�!�j@��2:@gS���r����8S�иZ֧9��6�4�ʥzɒ���.�oSNdU��>�+%ɀ��-��S�SJ������a�Az#v}<oĔ�8��۽�Q,�F3Jb��d�q�7���wJ�"��'�l��qV����Шv��qh!�%E��}�_�|�[�>A���iw`��l;�II}F�1|@�14ήv�q4/7=����cV�Wf��
h�Z��'Wy"N��b�["`�-�p+We�/�v :�1	��`r<�6�O��_�m�꣢]�[s��G�mq(uG8Έ����k��d/]oC���[��� ��������+%k3׹I�Y���U��w2�j��I��u���{}�3������N��0�%r/!Ƈ@�UeMwN�x��Poc�+098�Xcbt �n]X��u���v����}f���_S�y����Mi�3�u }����y��o?����nzs��TrU�K�����^Z�����[���f�gWO�S��ލ>Sr%�\vXmә�_vm�A���z``���%���!Gm=���P`k�>ڑ�i�"%_�X��'�j�݋����sp�ϑ�SXp'���X�����&,�bR��~u�����YL|��x1��u��ѭ��|�q�}/d+��{od���X�U1|Ԓȫ�B�j{�7���hfݧ�Q�evX7��8��)��K"$�֥Ǩ`c�6dxzKܧgh%�u�w�UDu��:��3`�����A)�֬�@o�e�O�F>C\�Y�n�7/_��s+�]����0T�{,���~�v�̛�s"����.&���8)S�Y��^v6��bh�4
R�L���V�
ҦFӳD%{�������5��V��L;,'G�sƪUH���Jg-��ꗒ�X�;\�P��#K;/��.2r�,XoC����/WN�G�[�$�Ç�y^.�@��[jJT�S�Sges��B0��STK�V�ryM�̷�#�I�/��ץ9���a'y{��I�Mi҂�u4kv����r���h%�Y5��#D/$Xd|��K��J��Mi��1�c�������ES�h��+>���\�q�-���������)X�\cª*e�o$n�Y/'��rH�)Q=�4u��ۀ����$tz�@�Ƹ�]����=׍�h�fmj7�[�����qOc@5z��cL�b�����u�!g2������M����#�<��
���v<���V��s�OnA�<Hխ��e=�s/:��R��Y����e���]�۸��ֲ�ga�xkv�{�l�6@�^ptȍ��*|�rp���_u��{ݛօ��ԋ��d�u����B��>��t��4 ,�wZ����ϡ�����Y�'5�Wb1�8ِP���Ϋ�8�^���S�7�����h��wf`��T}X�ɥ&�����gB���H���� *(����p��F8w�ú4����e"#N��-W�F��bg'0Oe��P�3�Y�8u3���4��m�t�{��8�8����YrR\�Gt�([���I9ԡ6)j��qIl���8Y,��|PDIC֘o��.a1�>+�N�u�͕�P>�JӋ]މxJ�Y��&1@�B0�=٥U�w��Sw�Y�Z�D��7�����8�3��P�@M7��,��e+>^aN�U��N���l=L�S��F�A�rEP���?;���vA��R{�������" G/6�z�1{���puϻ�%�;�*Y7�1���pMFK���х�7j��ΕT������t2�H�c��9���W�`[r���(����s:Q�^N��K\�]:�̉�+r�$+�+d��<5���c�a�a�L�Ƽ�;�k�3�����Ԗ�혍/���8��J0��2�I���_c0���J�5.��>���5�LH���]a.X=6�s[gB��u�(�ȭF����F�^&������XOb�Oa�f���	�3AA�vC�ޡ���X��T;*����u;#�蝭[��kfP�g��w�p�Ç�G�;���yɮ����N�8���NM�+U����%S�y6K�X-	ch�ײ+U���H�ۗ���H
�˃->�	���4Um�eu:�f����To�UǨD��O�C��vҒ��v�]����U,J�����\��S�E���eV)z���nA[���w�b��c)��N6��]��u�^��*��"�U��4��vmXRyi5u�;<����&D5.��:ݹ�m&]���G~�	���Zئ,�U�;Du�JBë�GL�i;֞��<�5�ۗ�~����%�{x*�.�*������T��{I��d�p�s�3m����T��Y[&�7-<��Ou�9gCx�B�i���lQWYp��i��[N�,��G]�<kVN�z�a��M[��Y���z6��*���[��ٜ�f�8�R��Y��Q��-^���̭�6;,�W������[gu�m�l��FGc{\�J]��a��1]qr�wJ��آ/�rnu�/XY�.nGuw#�v�`���z�|{*�qD��G|�/�쮲un�볛�;:�I6\�	e�FY|&gVB\�X9�\��-�Gs�&j����[i�܋k����%��t��Día�w������u8{A���E�+#�9mҕq9ޕ[����W�d�s�9zU��\ժJ��ΊX^!�J^Vm�U��O��,r��d�#��)��8?)z��W�7�qZ��q�h5�6W�)Q8��+�k��t������k\���uCM՛��d'w�1�Sڂ�Ǒ7i��-L*��l��[��qw[�����e�w6�p��
��YvPXM�	4[�1��]���5��r�y2����ױ��C`�ħj!E"o]��n��)�.����������"�[bT"�v�]��P4�,hb��Ķb��A��4�}����#z�"�L9��d=n8��뗼'f᪽�f���ا-���"��rY��2N��5a37��v;[���k�NA���K���T{	Qs�Kf�ad�T���I�w�]0��sF�"�r�i�����a�z��*�P�������m��Uj;��V9*p��)�U�����EeEsu��쪱6�oЩ׫-�TZw�)x�f�EI��i9�]2��N�����ĺ�귮ɮJn�W)U�1��V�4��c�v���C[��0Y!�V��zT�;U��ct�6%mͽ�w֎
��ڗ0��tN��C�7}b���5:���U8����p��e�b���U����N\ミz�X%��;w"ڛ�ka[�Vzn��]Wv�=5;S�$ݞz:���X�ܜ�i�c%��޶�֢��{V+B��w(��U�:�l��VkL^G#S6v�:°��3������|��h��s����"��c@��j)�H�E(#z�ۏ��x�ۏ<߻���|E&���-%��"�t�ܻ�x�y�&Ŋ(BI
�D�i맮8�<v����~����|[�e4F#&��s*�s���E�z��qǏ<z��Ǐ^���PH$ɚ��6��H;0D�l&қ���qǏ<v��Ǐ^��� ��#0IL]wM�p/:�m"��ώ��٠�;�7��u�_{.�c�����F�Kdnn�}�׉)7��Tcy�s2'9�	)$��]��{<<r%�Zu$�%)�&��_J��Ɇ�\��3�R3f"�rd����td1j (�0 F�ۜ�BD�1& �$��12�K�vL/]���%	\��4����ur��5����)$ �&�U;�:�Ϧc�sޫ=sm��֍׎�936�JB�8	K�B8wW&�܆����WX����|||�o7�<Qg!&�ɕ���;kzz�<��37�����2��@\�91u��X��T��N�Ϡ�����l~����H@C���M5����S���.C-<�b�sU�t��p�hI~�h��8�>�hք&��Э�9���lS�<<�#�x��U���t�$Oc�hdTn4�گ�y9ڻF�38"��#ޑ�����իb�z�ہV�&���;tϧ����}D���N.wd������PFr�*��ɯB��z�@�pw�0-����ٮ�g�0�+�����~ڹ�T��}�֯_��r��m�:�w�+�]sW����ҽpɜ2�~��'n�ET9�V���n|�ױ_56*��\�I���baM�q��΄�Ĕ�UaٝL��A�5�	*P�퓔�.�A�s2@����%7��"y������LZ�3���S�[�.�"C��ԌU�]c3N�P���D��m�2�z��CA�W���/W
}�N�Pl�[�P���W=��wB�Q�"�!W�U��.K�B�sr�0DbN�%K�W�wEŝ�o3�D�ξ��n�m�ӷ�w���K3�,a�i�7���]xBO�1�c�g��Ծ�޿��ut��pS�,;֨eSf�%�����g��ͭ^��;�mlԽY'���$2m����o���˦�%e��F�\�7��탋�0�	@nDM:���=5֙f=��W��Ά���-�t |a�墤�'�_%J��+C&(M\m�lB��ꓳ�$�mq�~�ׂ�,
aZg�3��6����a�Ek�������W��j�L��r���1��8��S��d�{0Y;M�ӽ�ǭ!!TDS�2eA��f*��_wl�)�&���ׅӟ'�q{�z�ɍ}S|�g�_~�6�N5������O&��Ǫ*�u��F�a��r����[b޶�7k��tqk��0�K�:˸�?	�=:+��ɏ�+��O5m��MGDgKԵ��{���n����[]y~�d��y'�À�~�Q6I�f�$�˹}��
b��B�f�ӳ����_�^l��e͵�J�/ ة�k�p��طlܨd���hga.�(����d��J�P��� �dx`��Q�+t��V��#"�8"]#�nB�^�Lf�"����L�0���Y���n$Ii��j����1�c���p�Yϟ:p޾f��Fv���ܲ;A7񤎴��St��8�s�>��y��9�n|�]t�wL�R�Nfm^h��W�w�*�R��=>�ʷ����͋!��e�oE-�������j��nG�D�]��1wR���w���u������!S>�A�S�`5�񫌟J��&�9�T
�<�Mk�����xļ��cmG���H@7��]y
'5X��w��i���ڝ�h��u�����=ڸ�:ُ�B��HrL`������74��9H��\�*/�9���i��-�؜s���$��5���F���:� ��U!�^U�ᎋ�[�Zu�u�e.�w(ǀ]�e�߽M����q��KV��Q(��=�F���ep��2^�֬*N���M-�i�KUVt�#��%�qW`�U��#�e@%Lo��gR���$�a����Ռی4(��8sF�rѫS@�y@��y�Sr.������̡4Ǵ�X�+T�];�=�[N�V��);j�V��C���޻*��]%q�n���ۇ�w`W7;���:�{Y�YDU�4:g<�k�j�ӷ��*n��Ǝ���3$�n��r�"|c�1盾�9��y��d1^l��y�<݈����߅jZ�]+z0_Y��ǧ�*i��OڗŅx���=�g�WTe�����bU�Zq1K�v]q�r;��ك5����>=��m`bw�?l]i@��'���K;��2��Ɠ&��t�a������ZHG�-	e�=f`�$�tTB�1A��"jK��kdg�N�Vm��,k��eH�y+�:yɉ13!�E�_]�����] ���8���{���Ⱥp�Ձ'dpx�[�MGY�j�l�v[���+���&��~����a�is�_u�L�(G�0��Mq&�F�U�E�zѷ+:aV_R�9�n�o#�4��U5WJ<�­�敠����-G���I�QI1ޒ-nU�����J�B��U6q��_��4u��R��|��w8��G9Z�AҸ�l�����c�63��<}7�h���.Pj�ڍ�7�Q����t��V�LAݥT�r�2(a��rL'�:ݸE;���b٥�L�Y+M���U����R)�|�FA�FX�{-�}�&�~���9�:�;�Qs�D��;�� [��o޻��b���o7�ߏ�R��`�|�Ȩ�֦>:iq��ع�D]�f�juڮ��^�g�uR杣|`)��9h�b�6kQ��<�F��U{��ecN������U�o��ϰ@~vq�u����A5�gq�/B�q�3�����9U�F��������p6��}7��k��F`�*��_Uy�-���g�3�q2��������mZ��[�c��o�G3���6+�EB���,.GOJ+�S���^@���A���Ԃ|ڋ���Wک2��kM�g8�_H�A*��n�f�ҽ�����3�֪=��ԩ��4���#�?�4l$"���3®��"D���R�QODߦ��ui�0G=����ϣb ?4Ҙ����7�
��"���O	ώc�Y�����m�>��~U�ATH�`ˤ����C�	�X��B��K$7Y�(~ʠ�Y0E�a�{/��Q��[ǫ�*F���m������[�XMOQ�.vnb
c��$"�v뮾f���rǆ3\ی������0��b��6�7�s2�]��s�ڝ�Nc����W��U�n���|%w�x�������ҥ�a��@��]��q�ٷ���s^间!��Kk�ʒ�E�����Xt�SY�n�C.�8�P����>;w"���L�sC�M��Dx�O�ǔ{w����h6�C��%�L�m��z�H�gV2� ؓwǭ��:rȾ��G�z�&��[=Ǌ���[k�m�i�T�|�3��!�J�]W�W��1�Q�)��r�U��=%���K���*f��w5j������6ǃS�]�,����
�|�,λ�pʰ�7ۏ�ȎʙHj3�^�[�a�y�����Ӱs�P���WҤ�ebw�:��ݶ|8�E���mv�i�7<���?G�-�L�f���k�ɞm#ePɨ�^����w%�1ʟ�n@�[ o��M�`K^shֵ��X������1�VЌ��9~hf�,c���>�������z\�w��7xf��5��N=��hǢB<v�v�&t�T���c�Gp%J��n���s�3/��~z&�2�a�{n��4�@�_�E��fc�;���ŭ�H���f�SyqH'D�[��ǀ��]QD��X�!Wla��a�X������۰N	���i��D4�)7U(���K���1�c��9��|�~�_ז%�����<=B[�A�!��Dp(�ǫ'������WU����J��U2�CǠr���xVYG�þ2�C���r������wOGZD��E���I&�g>�i�ؕb��qz��+�?�l
����$�f�Y�ƍ�F�p=��>5�yY�<�WDN�?N?���Dx�*��"U���W��7�c\��AS��26�R	�k�#��)�˦[l4�r<�IO��U�.^�@؍����ߩ8���^ӾAU�2��=>̠"i��M4V�gY>u�(v�uo�w�\{1��w$� �*�.����r�G[�4��&9��.�)���n�o{}!�۫���	���|{Y�k�^�� �z�Ӱ��Q�UQ�3���}���\��@7�?��^�kBQ"8�ے�m�7D��l�^@?Q��x�:ُ��p�>Aly�.u�8�W�ڵ� �Js2Y��!'W9����i�ctSֲsE����KR�.nT�Щ��G�_Tq�]Ni��5���vd����Y���nWV+u��Ӏ��8����s1��fj��8L��U�^���39�>��c�1�7�S��V��v��[�/)�U���Y���W����j�|tx�Sn�V|;��#G{]�d܈@�s����P�}Z��۾ێ&�M�A{�߳��b�����7l؈�"����y+]��
����?]+�ѐ�}~�ɏqZ/U�E�;���� j/Wb��}�>�煔8�S��ê�\�b���5/�D�Y!��o�u�3� ��Q0@���Ժt��ia�Q|��8�Z�gR^�e�t`:z�4�Y�[�Ψ���ea���E��#FL��7o���312;4���ѩ�C&�K����^@�{��y1�F��b��9�x�]4����;����8΀�R��F��=f�w��k/$�T�6!�w ���;�U��~{�ֱ��W���	�9�o��f^f4Þ�-��Y�5Tu���.�)��#�>�%_W�׮˨��V�ظ�/�b�ʍ,q/Rک�0a�c1S0!�	V��$����.Z����T{��&l�mU�V�1�B����D�ӆ�����bZ3u!�T	���Z37/w�z�U���+��bi��?��珛���y��-����D��}Q/�13���\ؓ ;�*Z���pUQ*�k����f��L��wa���{2}�5-^@�J��账��3l���P���}v������/s�U䒐�Ŝ0{�۳�R7m���7�YJ�&�ZxT�e������d�"5�g��>\i^<�RM�d��-��Tsk'2���2�ay���1�'�fY�^�ˏ>)��4�r:eq��g6�1�n�/a�lƙ,mv�.\l`��h�x���Q��CXo��o�EJ��w<SƜn٩���;�D<�C%P�e�t��V�z �z�Kzs�rV��9k-wQ���N�G� 4j�}����n0��L7�s���2�Z��}�*=�ǙK�\���w7�o���,�x��Ѓ��+S"~�������ki�C�1�m�+z�c�u��p���[� �O��<u_���NM��T��q�^����5����o �lp����݇�꾧?���!�UÛa2�֭�Q�f ��@Ha��R�@�.{�&��b���'%;��cB����X�z�6!ם���N�W]%�1r9Ss&��'Ml!�;��}egumP /7����y��z�m��b�y�E���)��v��}H�2-��2�ʚvf��ލuV��t8׃��y�w�����|�p"H�q澛`^Utfe�\����c���q3�: �0������=���K� ������m��H>��ӛF|S봁C��&�>d���3*��ϥe��M�ݙ�R�	]q;mW]Δue_=�:3�NU=�ZU6�!tZ�1�|s4szk9&�JS��;wQ/�V�>�����=s���i�[����cK/�,�t:s�*�%*��Pó(s-\��Zv��ٯy���py�u��}<��'���&�ॱ�8�S��]cV�֦����4���>�ߠ����A\��h͞K����&v˃��2�4���-�5��d[n��<�v!l�����ɐ��zլ�`Hx
22p[���!�s_��H���T!������{M6��5�5s��q�$���D}8�D��S���I:�t7&�Wv.ƪȕ[[��z${�l5R���m��uc�tנ]��E^�ږR���(�9�Y@��mZV�5��U���n�)̲Z��3�hqP�Y��a�=���F��^RWi�t�͠L�v����}�����]֫�K�Ŗ����zMb+T��aus�y�����n\N�mmi�:3krQշU����d@�i�����HP1w5m�Ɯ|J�������ݕ�Bc�W��OV]n*���{iT�k�0�]M�W��-9-��=��2M�ZĄ<7i�	(�G�7�w����8���"�&A���م�V�p+9֗b{aHr�-��pk����m2n�q��[A�[�u�T�dV�����Ml=�1�sT�SzIWQ�)�XtY�ݾz�;K�l�^��0��������6۳���'��������hX9Ĺ̥MЂ��j��fS&�)�ٙ�:^e
��y����Һv����U�d�Y[u�(JAN��Z��l��afޫ:Va�6��9�eu7wsb��H�X�C��h9U�@�eң���ȂJ���7[��=$;���k."�!���U:`� �*��:� ��j��z�ͯ$���逵 ��p��(�S2���M�(��ܮ�f2S+UX�AH>J��J6�V�v�O��'e4��n�~~% �;5X�%K�"�!cr"Nۂ+I�:*�k�ۏH57n^�[i���w7�2QR��:�vbL���n1Gd�w��|GD��m���L���MjoG�::�L஁�)�J�`Uƶ^MX��)�;'r�5.J�_<Z�$�x����l.�%�4��o(r
���@Ц�VU�ѻU�aJ�u������6�͛�CH��(�s;�c��4�Z�)z��U�����غ54�/∲�^	�Q�5e^S)#����N���jD9	.!(h-/&*1��R�N�G���vv�X������s�,Vt���8�J�"��D�K\�R*[�Z�ɵ*�d�o�͐8fL{�ǅeլf���G�`�c����������&�G�ѡ���Yw���j�vuW0u�m�A���Ҫ���^����j��'r0�/\6"U�{��qئz�^�U��Rr4�q̤����A��+˧��C3^^A���W9U{���*�u��>�V�8��6����9uύqm�2��0䗑�|�ٮ��v5�6�Q�[�)Uƌu�:��񜎁"�bo����7�h(�^�זs3u�Q��q٬/�Y�5w�:;^�+�z���o���k�b#^8	�p��sՍ��I��˧��ι�����]FlES���0�$t+�I#�޻�:��$3��"IN�档M ����_7#vz�m� h;b�h(%8��r�rD�!����B �D8�.�?����P�� �
I�,�6�NW����)����nʆl��B�,#ӷ��}q۷n�_��oǬ{�!���䑈�
"�dLĜ����MdA��^����v���n={�I� ����̆)����cc�(��Ԙ��"hHȲHB��ƞ�z��ݻv����7��{��:�JQ؋�왒&��!2�"�!���z��ݻv��o^���	# �uM&�d��."1�	L���n\3S$`a� �H�f�M���K�Hk��	�7�$ID�ztJ	D����Rd���4��a1�\%�\ �H���H��!FHX��ӦF����Lę�&J�
}N�$�쯓)�+F�J�9J��3b��QXh���F�:�qķ��]pw�i�o�GA���Y0�K�ӘJ��%�ݼ	�(4��<*�i8�QPd�O���~?���鷺m��u����ZU�L�E��f�j�P~ܥ�����D�A�C����ۺ��d�����ݓk��>�?��y��L�4A�Q��l�}\�lV���M�GC�r�䶊&�Kt=fR����1�7��39��g>��aȁ<ñ\?�.Et�}X7`��ݲ;/s��>�9�Kv7�:]�DJm����o��z�ei;���oO��r�U�7�x󒯮㍑\i���]�����úY՛�ZV.�����إ�t��'���-ps1��}�D���1�W�����I��dpϯh}�95g1�Q����ʋ�/9H�\�<�]�ȨX�,?�P���X|v
񫽉�{��fx��;���!FϪ��cl� �@�6�ڛ�Q�ٖ��-xs��t(X6�=������E'�AN�jjϗ2c���xը"V�#j�
�a���e�)�9X��E{g�|��Y_fGĜ��E��!m��b�;�~��ܛK1A�{�4�ٞ�ڇg����s�.�����cm����ĵp���5
w�*���;˫N�\��}U�tͺE:�4u�!�w+�=���������v��[#��@kE@\�G�)�q�G�+���EV�c�A��c4�ꉚ��O�m��2�;�q:sSǫ4E�5���7D����m���GGfd���I"������u#���2�͞p��=y���Tb�;g�z۲���=zހ�d+w�}!||��i���R���;��G�������k�;��F7�:�I)<ir��mkgd ;���٦"^:z��ۺ/���i�LFl�>���v�u��3���X�o��.	��=u��b����0u�mvTq���"5L)�<V�3����]Q��KS|Ik������T�~�`̸o0H�0eWB^|ü۬�<���FƩ���r���l1-يW�zed����-`]�� ,�Fҗ�2b��G���!,r.� d����e���\l{ylu���-��T�l�<Uz� ��`�Jg�jr���T袞k�svcvc4�=�9���Kpa`�5�uᱢB�X��x}P�NӌYD��5�,�p�I��Gn�Ε���1����:�\��-<�����0��n2k�u�����v4
����������/H�)�}Z~}mWZp��葶+k�&;�$kUv�u����y��L;z��ں1�N�D+����77G��X97��<�w�,\���M���͞��n���AJ�+E[��W���\l���m�/��me������Bo��Q��V�j�I+�U|�')=��w�'0ƙe�!���+�?Cz�I��M���P�g�
�:^����y��r��f]�ڏg�s͝�p���6f�UPG�&%�[����V?|����ʕf{�:3�1�/#��J���<j����B��t�J�
��R���ne(B�V�B�G9ҵ`7I�)�w��z��*C\���F]t�f|Ы|A|,^�p���}�9"���i��^(LZ�=UO,#{���5s����������;.��:�zx_�D��~�j��h��So.���Ha՗.ɾ:�2V�Ҍ�n�z�Ō�(V:Ǖ+���m�L�U�S��ӝBe��j8ɧ5A�['�S;ֻ�t��;x���o,�t�a�ț��]�)jFNG�V��w�ڂ��m\mI'-��̔�c"}�����{���zVt��;��5��c f
�308��3���{�{5*߫5�1ɋ��ǂE�^�ŝ�(�Y��8#���]�ح��Mˇ"r�J�G�?30w��3�Ov��$�S�v�GWn���X���qwS�<<1�f�ky��@�8�����{P=��ΗW�`���t�u�@��X;~.�KՒ."Ujn�j�v>�J����"�<�'�#Cy�8�6;���nٶ'F����v�n7$jǥP�0e�s޳��Ĩ`ʺz�&@$�����kT3�����o�7���=Z3��:=�{�2�Z��\�~���<��\� �Z��T���ѷ��>ʞښ�V��;H��O�&���K7CXǽ�S}�F��#�������a=�7�d\ә�i� �������Nq����ֽتlS(ҝCs:m�HUC8�V���k�I�Qə�"�}5/eڻ�ièo�����ጔ����k
b�����U�l�'VU3���侙�j��w����fa����&��|�6���H���ID��o�A8&�V��7j��Ҏ���O�_GKj�j����GTfgLj���b�*eձԮ����8_7�PhVA`�DC�[,�bS�,$eI��>>>>>>�P��A5]^�ȇ�,�{T����dE,�#�gBD��q��۶��]�X�;��)��g�춒&����<���P_Ӽ#���N�}�f3�s�]�vf�Q��۽�5[�-�x��o�͐2�Ύ�p�F`U����n�+�j���Ln�^�3�ݮ���M��Ёp���nT'�鍁�WZ��	�s#�X��yޣ��D�{����Q��~�{_Vv��M�����D��V�����=�6������ȓ)8S�EUu��)8��-�9���qiO�0k�B��&���%qB��f�e-����d�*�p�5�2�&��"]t}Y-����œ�cb�	��k�N���?0�b$K�r: �x��X���b5�Q����݋cj��;�3V"�����DvW�6�#����3��p�tv��`�^V���E�6u7����>������fs�斝Xq��Vċ�\Ʈ:_������J���~��F�G>��_K��;��D~=�����!U�	=���3��/nP���������,C��5�n7�e��f�/Ox�ދu10��Bi�{��Y�oUW�*{{��=%��0#�|�;,��1g
)��@#���
5�z�j��E���wlii�=& ���<	͑���w˯�\�s�ܽ�}��)�,ٱ����n{��D4���'[�=��;d):��'Z1��˦H�mE�ӹS8�����y�Μpz���L��H|t_l�֔�Q�	�@s���Os�k{qI�wF�dPa�s�6%c����͝���ET����20�a[v�B7�GmϯU��g�~�FsF�8�6;P8���5x#�(�D�ْU�3�v+�A*UO����u�p�t��,�{��Q�/*w9�֢�coAKy���uwl���쀂��=�V��(�70�"�S�^�-qi��E&��OF��nu3a�n;l�R=�Z{^L��:7|��rC����
���(�ݪ��$72ujo'i��g��ی*;��9+
���!��b�&���3j�䕡qR!�\D�m�j�����ɰ�4�e�T�Eh��s=I�ɣ�h�.�Ѝ8��VC�4T6��9\ռaW*�r�D�8��nH9��t�;tu�eM�e��X-�� ||�o7�����"��7�y2���]~1��@����T+y��\��z�f�������1�ǛR�FM6z�:3`��^����M��}ӤU��V;)�Pz��\�M�����f}j�¬B��C}|ߧ�>��c%
b��V�~zx��}��G�'��t�1�/9�»)�Q�k=����Zn+�Ã��*�l�����v���O����N'�o�憻y
�B�V�K\ʼ����X��`�0n3���D����D��	T"4�_,�Zg�5�0�7욇Ie?=���#e���Z+���sO�u�����e+�֔��x����gr�k��
�P�g���Ǟ�	�=>���r�_��F��\�r��"v�zu=�'�*%��gAO�}bLa�_zޘ���֬����͒V�\33�q�^���̑�Oi��Nofe��7-��%J�JUDu�-EWl�]�,�:��n�MVB,�6o.��P��B\�8�.�]��ʝ�O#֒ۚ��*��]��j����u�?��ek��i[%Н;Ƅ��\̚Q�-uq\3��y7ub�}�}[���Io�x�������D�:GQ�Ŕv��%�/�V$�����Ud5�m�e®��$����x7��j���VuyF�>Q{�+��Iy�L����cć��:܄0�<�{����O���:�,�b��K�K��V�El�2��m@mN���u�.��#o��z��n>���0�.8+����`�+!^/�}�/����H�V���_b�5��WUY�Fe>P�;#ͮ�dռ�[���t��NA[�;����x��k�������$�k�V���xk^�O��l�d�XW������{���o����.���:,�`b&ښ����ΛV��qjeOa�Գ��iz�wl��a�iJ'1��[��N�BZ�*x���2�58����[�|I���l������d-��I���������J~�b�&����촠A�a�w,�E^E��'��̳]3ĕ*��ٺ��&�uE#,�7lX��ۼ��G(��q��2(ح�(z)h��"��X�t�Ò]mr��	veE=�Z�j;h�&MN�;(\ɋ���40��D�m��4�q��o+E��[}�������*(b�I#N��*���=���-{D��>��V���cl���_x_L/`4�S�������+���5H4UV=�������}yfz)�a�w_�%{�7���HA�"����_c�n�3W�����7U��g ��ժ��o'�w��ͅ4a��h|�2+�tT��Smz��)u&��ֶ��ryr�{P��b�M�ٿ~r��1p7X*�r�Z[��r:s�*���(�*KFW0b�W��T�����=����H��Ӓ'��w�l�o�
���٦��Tʧ���yH;�.o�s^_vr�rz��4C�Ϩ>GBF��qlmm�f�Y٣��-���F͡�v���9�[Ϙ���^�0�n&5n�,�wv�G:�Wdn`m"$FĈ0�;�mM��������Mg���z���Bpk?x_c�uK��D��n�GƱ)��q>�onɵ�9�>`�ϣ&�I�^8�//"Ҥ�R�h���͊��:a�v֗��*I3[s��H�,=܅w��.�"��x��}�7&$������-�|a�?#e��nnY��A�U�l�/��b����wjoe�Zw�y�����A9�36#$��j�G�F1�c�3�3���~f��kfbfwo%����O�3w�u�sLt��7���W����8�遑�.+��������8�`4��y�Q
K�5��u3�r�l�W��ff0���:���ZU�vY��ڕ�ݓ���^�S������f���˝u0r%���f��N�=T�}�T�ch��n�H�{��`w��gR�sx�;٤d�6��t�3�4�}�t�{{e"Fv�Mu�r]��az=��T���n����QU|��u3�Z����^�R�m͵eKk
���"����v=��m���%z�	�4��̛&t[��+�()���`M�{���S�i���k"g����Ȧ�A���0v(z�����Z��xo��N�N��A�p��%�/N�ٝ��[<��A�S{���߇��@ď���j3�0��k���l;�i[�z����:Xk��>�lVVm�����δzԌ[ݽۀ�b�*�hd��l'S@�v�S��gz4dmWY�qN:�ҧ7z��V��8Z���]H>K���L�A���u�i�7B\��1p������2�8�*ثـ�gp6�\W۟"lj\Z^��<���	�9
*��$�P���?�x��QX�SW��u�Çleek
�:��p!խ��eQs�/�B��[�=Y[ƜK���C��5z��)�ly*��둹Ucn���St���$��	ond7J���S�r�S�4���7�����T�g�Q��<h:)����j�%�Լ�ZΥSQ{���n��v{q��t��A�v'l�ӝE7�ۜ��0m�6�s:���Vqr�ٻ�&�t9]��*'|8b�Sb�Ty^�}��劖�s��ܫ��X�X���Ms��|�;w�,��j�М:�$��ka��{Y�EZB.䓓��1D��ɑ�N/Y}@�
�0���h�e�I��EQ�r乓b�w|ru�/��|�E*X�9{|N�C1|sG֯����jn���I2�]�(>+w�,���#YwEL����u��(��Mªƛ�s��g�r��{T���t�e��"NZ�a4�9��|h\���p>(k�[#�����|;1&�����{z��#ٺl�qNݸ��7x��Td��Gt@�';��Rv"od�o5�*�j�X���q�Iiޖԭ+ҽ�C�ג�� ���2z��Nb����um�T)����r�L�[F�ڧ
��g����J��+>�C
�+�����!��4'�tЄ��<6��tX�+^��a�����;��j���ZhS>�L�Y�f*]J�QQ%8�Q�um�)<**�R�n��/:���¤��e��V�Y0��ᚰ#�D��!6u��w+ƧT�г6µc)�N�����X�f����89`v�Ɖ�>���Z�׷��K�)�;eVf�"�v��1���'��T����w�e��˪���KR�$�+���ܭV�U
�S]�Bl����q�u��yj����"���s��w��;jc����~�+���d1���;��N��7F�t�.�p�±�Z4�Գ9��_T:b6:U��
R��HP��>�Z3^���CD%{��Uì�A.-�ܘ,�U{����!�05�j4�Fܴ���Tb�>�,mM�NR[n�V
�sݫqݻ��+�8�_B_[h���YJ̣)�T�^��k�9�q	�Y9�"![�ǆ�|VUN���[�l�Uu0]�ia,�=6��l�ÝcFY��3�#pU(w*�p�aǹ�!��v;�˖"ِ^�
�^?%����sFZ}�vp}|�8��HV>�+R̞+l�G�ܒ��3�N�mމ�p�Q��E�
iuܺ�풦�w�*��r�ٲU-O�����ie�Z��W�S+,=}q�n$���f��g��Ұi�^5�l�V17�[L��CI�T:�떛Cc�':��[��}��
�Z�JA�wB�����:'��;{�ŗ�r(���{T45cQ<x��YRR:н�3l(�L�A&�P$��#37� �3(	����I$d�)�8���ێݻv����o����vQ�6e"ϊ��!��I	$;AP�t���Ǯݻv����7���o��"�Ȥ�6(�:�I�*M�K�dHB1��^�=q۷nݾ�v����$"�@&Ybf�i(�5!	#	��ׯ_\v�۷n޻z�����BHeBi@a�H�ι2"��R)�G9�WXœQȆ%1$0��b22	Rdj�3 �$"F�I���S� ���]%0�df����$�,��K��c(0�%��i&JIH����"J1 c@0�d�wtј(*1c2�F�#oϾ�&/*���ؤ��}�bK ��(e�.�խ�p�w�?Z���^j����
�-$�(��XN�
�aWo+U�G]5+�0�t������y�"���.//���g���	T�p:���i}�rC��S��n+�z끇-d��j���� ����8��s���t���y��$r�H����#�8�<�m8%�������{e����*�*���%��2<�����莍���@_N����3^ww���l{~йDz�����0" �\
�O��r;6��3�SvtF�V�[W:�J�D$�L>��n���ַJ�ȑ

w�"$��/�W�ͽ&�&��H1?i��4�ù�εA�*�-м��~�I��L3T��Z���:�u�g��.U��C��.�;��!����U�����+m���8D�9����A׼|���s��ZE��Gt�z[UzƫJ�`黶4G� 8��y�o�U�D�!"(.Qq=�e+[[Ӄm��j���Mrj	��V"�w�hA��H�ͽ#M77��Λ�+M��^k-�a�z���r�U�Z&[ps�ҳL\�)�3[�4"ejUZ��t�+�d��٦�SP���2�Ry�=������4������f7g��0�x^����>}A�mW��dWz�}�������(�����q�jBY?	���iǺJ����n�
w��w��=��W�%^}�� �����;�CZ��	�i=pD��,�qa�������Э��&?r�uϥξ]��ƣY@<p7����0uUx��2�m����U�gCY|�Wћk"�F��P��>����&���t�%x9�*�-HܷX�����uo\ޥb�i똯pS{0�f̀�u׮@)[l����{۾�n�&bΝޗ���=�r}��[�Ñ�	�5�ї�+�L.&d�qWs8ӴIi1&5L�b���5y���Zg�tz�l��*�\cTWo[����@��s����e��h
��`���ˎ�R|�.$����o�!�s�����Agq�;��i�\�F�@w�{)��v
�j���5�� ��1��Ia��:���[��V惄)cMhw�e�+��Ǧ1�JS����)�ʉH���*�4f�&��'�f[e雐���V��a]���̛�bw���H�szַ��ڬ�T�q��:�]�Vӊ'R�Q��*�����R?Č�ּ�]��v�F�q��k	������.3}&@~�'�|��l��a��hx��
	���rP�����V�"�a��Or�Ժ�.�w�9�ņ���ܗl뛳�i�L���j���P,k�Tx<e�z�)����������x{���F�;h��t�N�ݳx:����;����gE�uE摰��j�i1`����1�����=o�$q�pV��b/����>��Sˆk��g�*;U����å���#��%�W�3�	�{��;�nT�N����K훽�ZXk�j���d���v�&_s�{,�m���S]�Ҏ��hq��U�,�����leC��ʑw��/&t��Y�W+p��Mzz{;��qmW}h�w���� �����o�=9�:+0_��,�#��$��h�n���H���DkmVKii�@VQ̩aQs{��t�`���]�w�7�{,I�P�0f�;�v0$�]�w���=�-U�7Clڠ��!�8g��x�1�m*l�[�+)�����Bμ�$�ʍn�Ǹ轑�/n�R�*�8�L��(����-�-�]���ٽV'5T?�^��g���W^���f���>>>>o7�74l�"��̞��$��g��e��H�����NLh+�ܷ���2Q��,w5��M��(���1?�{��m��!�d�m�i���9v���ڝ^�~�|Z�s�&�`�+3�1�fG0������VF�A���Dg=hR�J~�U�ck�(f�U��K9��6�@4�ƚZ���Ij"8�v57L
�FE�	��v���ZV���7$0�q�7��p��Y��ERR7�Gtw����r�Ft��_�y��-�#mi�2��Lw��� y�
��;@�ޘ�V� �1C�Ly�˅wI�FDCb����|a��c��"%�E��?]��F�mSB��������J�Yr��{���c���,�wV��@~��{yqby�����S�Ƈ���f��Ș^؋�������.����S7sxd�:�*���?����v=�O�m�Ť��ٮ�\�M]��vlڭb��.�s�\��"\$n���GS&qU��U���L��Z�}Nz��f���Yʯ�\��QM������^[ڊ�õ���|��C"	�e\��~�O3E5�59��y�e@���1�cy̮���k��z�͎;�!GH�Z���B&�Ԏ��;X�)v��27�t�z
�o����>�Ĥ
��7���+��쪇�b��f1|�}�~Y�t(�U P����%X�&y;�ų<'�A;�#������'n�S��p{�E:�w��֊�9�Skp/'QD��&0�f�x��pk�IVWE"��n]:�p���7N������s%Ϫsh32l�.��)+�\h6���WQ6g͘�s��W�^]focD��0-C��c�Ǫ�
jSCe��U�V �l`��kb��=3:�i�|������n��{�1V<9��p���Q�kV���f��
�=���1���,��:��Wo��x��"1H�a>-���[�D'�1�{1�N�2]Y���a�P2O�p�C�t w���q3��Bvb���4Jf�B3f��*���Z�u0�����5�a\�8�fR�Wxޮ�֢��0��̥Ț}4^�ܓ��Z�.���r�I�B��
��s�:�wg���Ei㳠�X�C�{���{�@k���7�1��o5����}�>o/�B#�j��
�^�!��:�/D�V�"D�[J>�=�f�`
W���_�uUqn�'g��m��Q�wwKe(��%w�Q���*9"%�`����y�[Y��N(���tQ׈�)���o>�6�����?*z�24�÷�y]ޚ�쀑] ئ��
�e�S��u�ګ���
�_@|�j*�R9<��`�|YGy�$���=��j�7�V���z��J�K�}��j�P�w�0el�9]w&�ɵ<O`����0lm3���|<A�\Cc�����]�ݓ�S��w������q3�FMz��ـOM<��竇2��e���4tZ[�Fl
!�<�E�.���y;��|����d����Y�x~��g�Y��kH���n_��x@��Ft$ls�y׏<Ɔ��	`��K%�,�L�͍#e���u>���u*��X����U[�B16VW<ò��k!jn�8�,\D�N�V�[�����F!R�)���\'U��t��d\�Y�㩷���_:�m��5ƥ2v�v�on9�Y��|wJ���))�i�!)��g}�������F��t��W¡�<�cZ�I��%9��|���"�V�G�l�kLϣ;!wf5>����� �t��c���R��;&�,���1ݣanS��D\ڲ4ù�伎k��H�+�p�)��l�6�\���]�s3�Zb��ѱ5�ދ��3� brrW�	-�{����-���ԧ�gcWW[R�Ð�Y���w��,�=ԬQ�,1����C�*��5�s�dG�
�4�v�S�p^���϶����\��w�k�|29Ji�p��		���8A0���3�l
7�s�ݿja����}T�Ā�������������]^�FŽ�vK�c���e�� ���s9��:�y�	�5��}|΃�\�b?���mN��.��uKH7T���>��\�-p���q��/"����*S��=3�Qn�\Y�Z�}HtZlÃ��T�w�5�b�Ș����Ɨϡ�O�YrN���[��kt�#Mųf�5���jp�=�%7EDC�W��szd��z�Q�Z�{�U۫�y�����1��Rɼɽ�20���roVM���������9��s�N�v�9��»��^�k��O��5��[�4��mk�ToY���W��=���2-আqJӔ�������z��C�e/!uo4�j6c�m�_���,��G/ViqT�3��*��V���n���}r�z�n_�7M3�H�0��yl�[�a�ثq5΅��[��x�Lq;��q�N������Z̒�����xΪ�:�kx��Ƒ�6W$R�d�=���,�NX����yD�Lq/�2foc]�e����m[���+�<��qk�
]�Z��x
�����S�le���a�0n�������)��"��P�F&�s�����_k|��㱵
�be�x2}>�n��E�[X*�P��֒��1-Oru��
�S:w&#��&zGR���4��p�O�.t���N��UX&L57�J�[K�6ԉ�جM�tf�O����)	��5���H�*Ԭ�k�ƨ�᫫��{��M�K��9(j�s���u��%kzN�Az�sΥA�q<���D,�89��G^<r0Lך�����Վ%��o���۷w^�7��6y�8�ΞGT��UbiQA\��BW�X����;䨶�sѹ�����y|�`�����nOv��_����c���|��0x�WLe:�M�[����a��뼈 �h�;#x��$�Sl�>d*}M��i
��n���0lA����y�`Z����Fa�D�<�S�*vL[��l�Mj$&��私�TETK70�t���#�}/���oѴ�Uۉ�r��Q�Gsk
I��[���o A٭�g�$e4�vZ���	.��o�	����Q���]�Ծ��>�эؾ�:M��g�/�;��Cj �ǹ0�E�=��y�/�["�1U)�"\;���]M]2��V7� �gC��E����𝜺84�u��P��d�@ׂ���"��Ot�}�R��;���9r�W��|�h�za�dN%>��Fl�ls�4l���{S��Ł�^�ɧPc�Z�Զv>lpi��v�٥��/��r�5�8s4�D�4/FTe0���ɨA�!��`0B]��Ri"�$�H!�+]�W	�J�e!hy$�H�R%y"qJ�e�(��	MN���d�ŧw�um���;²��X:�,=r��z���f���j�{ƎS�����L���7�4�&�%�>�[�׽��9��,rq4V7r��W+:y��UM�N�]��\��F���XAo�zw=��W�]G�~fg7غ��u��52��_��t���m"�������En"���۶׉�L���eS��'3]�]�Õ��^��'zE�(
�a�X�0r2b�a~+�Hw�[OuO�l����l��ߎ>`<εA�6�+�xJ ���%����V.HujY�6\q�V���G��OA�!��:�����1�4�/'�^s��g���O��|����l;ƞ��D��-1y�x)n���5M�����/�D�*)>OP���M����wu�f��b�O>Ӄw�3�Y���6�ݚ0@�ha`-+���T���! zx{��r��������9	��=��������������$G� k��AA�����)���h�@j���{P�P���E 0T�Ee�,Y[KVٌ�Z�������*ٶLc5����,�fږK6��f��,�J�Zc�Z�56�d��m����S3)�Zb�Ͷ�,e[Lc&V�ɌզMMV�1��d�3m���j�-SkY�32e��Ɍ��Q�Zd��m1��Lc36ښ�+i��6�X��,YV��K&Uf�ͭ1���Vj�Y����ZcSkJ�VVU�5-iVj�Q�VVVҳZ����f֕�m+6��եf֚њ����f�+-���V����f�+-���R�m�Y�J͵+5}e�Ֆ���Vj���Y]5�����YVmef�VV��YY�����k+-ef�VU�f�����YY[+5ef�Vmeel�#�� ��
�Ue�T���JͭT�ժ 1D@ 0D���J�Z�YkU++j�f֪VZ�J�mT�����((�kZШ(�++j�e�T��j�f֪Vkj�f�T���Jͤ��@ 1 @ -mT�ժ��Z�YV�C@ 0Dִ�15++iY�Jʴ�֥f���H 1T�A�Bt�
�@`,���em+5iYkJ�Z�<�y��e�+*�R�V���j2ژԭ�f�+6�ƥZ�r͵5���kJ�m+*ҳV������eZji���w����G���x"���$b*�F'�p+���������������������~���o�xO�~�����~7�������
��������Oܠ�"�� �
��?�?�?H}����Q��}������
������#�>i �=���~������?��}�?*��-�-�ZJ�T֤�Ҵ�K*�l֦�ԭ6��֖U�ij�զ�kSJԳj��[J͵-6��eZTզ�kMVmi�Z�Mm6��J���-���֖��5-iV�Դ��e�U�֚���m�em+MjjmieZSkM���kM*�M�*Z��ڊ��V�[j6�͵�j�kZ(E$�
 @	I5�ֱV�V���ZM�ԛZ6�i�Ԗ�ҭ,��-��J��*jK���%���_��
Ƞ"� �H (�_�?��~?�o�@�&�g� U���?/����~��0O��x�����c�K?���@_��b~}u�q U� @_܇�A����DDUu���Ј���@)�?�P����F�E@��_��G�a�,A g܇�}���A �H���3��~���C��}��@�O��!��cB ��p���� U���z������/N~i��Pb]�~�������<A |Od�`og䔁���7A��^�:�`EQ�`Pa��₨�S���?���	���e5�SQ��U�ݘ ?�s2}p$������Z��ղ���UH�"6m�T��*�@%!*UEil)�$SF���b���IJJ�ow��T�QRB(J�PF�5,�Z%�(&�km����ٶɤ��Z�[F�#%���]��ɲ�lŠ,R�j�#jX�V[	��-���mki3��4�Fh5U��w-T�gZ;*��ŖZ���%���V�+T�Ͷ�6�[j�[hj�Sc`��[cVU���M�fٚ��55M��KEj٬eJ4���h`��Qݡ�M��   ����em7�;E�mv�wwV�Ug:Um���u���m���V���Oz�k�Wn�]�������2�ع�ڦ�m{u��n��븷m���Me���g�=��I��u�ͳ6����wn"[m��f�|   �CM_b��h���t=��w��ٛ�"G6^��}����Ѷ$-�6=���{uv�[���m��يֺ"��N��j��j�m�O\:�]��x�9�k۳����h�����ڛk.���k3&E��6_   �|�i�a��s��W[]��mm��n�lh���O8����e5�^�w���ٕ5+[65˕]aW�˵{��GL�MM��.f���[n�5�Mj�������jJ�ک�"��  8>�6�}��A��ʮ/]U��:yd���:�v�m���5U������J�-�'+��G�׶uj=�L�^�]U�u�^vf�i0�cj�XL�fSV�� ;�d��jͳtݖj�$2Y�̠׋���SO44�Uzw]�^��@�w��KV��oZ�Tk6�P��*�[n���,�ҭ�1�Z��m��k| ǟ`��GhjUu�a�Wz꽶���k1R�U�UU r����]�WN��2�n׶w�]]���
u�Z�{U�%�{3�n���cdښ42�F� ��)T���qXt����^��=*�� �w�� ���VpQ�=y�D��1��J.�b���=*�
U�{< ����)*@��Hkl-���6lS-m��fپ  ǚ� �Sp7ѥ.��ozT"*��{�ol����P�(%c��)"�oQ�$$�,����.�]��z]�(
ow��GE^�W{֭�յ�F���Rm�i[i�g�  ��H�4g T 燹�zT���=��kT�z��Q% w��QRUt^���$����@T��뼑J����ק��Q�ɹ���ɳmmm����d����   =�*@�:��D@�9�i��+�A{�W�UT�{j��޼�V�����%x�:��9�I){5u,u�D:�w<��(U��S�	�T��hF�4Њ{FRU#L�Ѡ`�=<FU*�4  ���R�� � �=��LT���Iꔈ�*�  f���?������?���������n��	�m!�����M�2'��>�|>}�˪�� �Z����UV���[Z����[Z����mk[f֪�m{�>}_����?���^�z	6R0)G
y���b�Ypuvj���AGwuxq�k	�*j/[ה�xE`�2�;Ěp�I&�F��卛jJ�2[�W�� �3�H!�n�n�B�ec����8i���IYj|���t����)�<9)Ñ轍ɭ�-M)K�,��v��'4��73q���ǷPEÜ��4M��8�d,�L�w-e=��)Yt�BitRɃ^P� ���32�R�Xp��>�1.J���)7�A;R��q��n�ժշ�ؖ��J5��[���1�i"�rQ�Z.�*62�G�h�͢�ob�����tv�p'P�
��=��e�E�D�v�Fba�Jn�ɱ�&�f<IXU���ж��VnE3r�@�Ź��R�j�Ƀw2�EB�gw3X��.��h�cr%N:Tor1[��Y�H�m�L���Vk�
��,�I;��
n���[�9G��{��}�JlE�g�Kt�ڹ�,bR�E��/jl��ų)C
TJ^61���kChY��/��X{�V�VK�A�6I�Z��p���U�$�u���Ƣ�}a�Œ��Nj�ԗX���n#H
���v5�	<݆�).�s���C��HnZ��������1�4.:&���k�;7T���1�@Dm�lٶ�n�	Lz�a�y���u���i.Q��1k#8	������V�&[�2*�tf;�qѳ��{Ki8�T�fVAx�������4���dO,Ɖ��5�;�Z
5��;ܢ@Up��u`�5�I��&a"v�;�<��C�(����ݭ�2�	���,�:��E��n��YT\8����I�tUãj�p�铞���򓰹<3{Vx��`�X��ub�����U�b��f�<�/��|�jO>�,�uRYi����i��QX�jn�W*}�f����X�۰	���Gl�y4Yif[rĖ��W���<�Th��Wl(�ua��1Z��m�����.�$E�@F�(�-RחYr���,̫�Z7���)��c����d�
˺[ס+��n����-�e��w����7�`f;��dc%��
�� J�:^Mɲ��И��ylP�G� �kq�P�r-́�dy-DD,D��r��:��\����sR��e u{�6Z���8am#YQ�ii[�0������yY�9&�Zc��ح挴&E�^L˷�պ
��${����t�X+#X�ӹ�ì�
Cv����Y�3n�j�ث��R�n=s㻙r;��#c,�2h��.���S��VM���1YNJʋj�m��8��
���-�4��אk��N毕X/I�T����bn�+k)[Cse��b)!e�����E-�6���,����+hհ23������������X�����Hu��IRa|��cV�F6�b�	<�V�6�U�2;�lb
6��oDE�hP�1T�R���H7����Z���j�D3NU�٫IN+�VF�Zc�re*Z��.�- ���`e����5xʕ5-�
�n:͖�٨�;-[���7FZWӽõE۰S���ɏ3	��f�Sͺ�����]Ե���Q@����j���z�Vh[�h�m�+��d�7A�B��;��F��ʼ��v�2���;f�.��#aHI{��e�hš�i�cD�� �:��[�e�&v�M��c�H�)�Le����x�Jpd�ITT��SV�^�="n��p�ՊM@�䞨;h>3pw��vtj��5M=���q)⎒�K���vDHZOp��G7-똑f�F�f[�U���dE(ټe<�����C��h%	��4�2�nv�5��zJǈ)c�{Qwx�ƷCtlw4��q�@d��BO3鮑wg!���cZw�l�T���v-\��Qwo+*���B��cmEb�3��mqȀ�&C@h�ZeZ���b��u����lн;B9M�s3j	�`���b�Cr�`��9@�lKf����Su�B`⡹�B2����Ϙ��7[�J��U���a��(ha}��5ǎQ�%P�j��-}m�K�L#j��S!x�q�iP���7K̻SY�T]Hn�)y`ZA�w&7tV�`j^�ý����!�LUr)��%M#O]i�ܵ{iR��6���H���R��T76,[6�h���v3���y��L*d	�a��d���Y���P#(+ U��dH]�i�b�Q�#/�k 7t��R4��^Z��-�mm%�B����oJ�Tȃ�X9���n�$n��L�lު9���ӑ9�ظ���Y��o�v���CbL���
�B�f1
ҦK���Y�4i䄳5Ӫt��E�r��7"W5�) ���9���EAX�j�[�o]���i*������I<�{�+�2�f��ڬ[���3��;��˩m
���($�V�ϭ�橢�(&V�]G�� Ц�,��f������YP�ZC�b��UyVr�#+��6�?��M:��Č�v��b�'wtpa��JŚh�g�իM��!8��[��eFޕ󎅭�
;�r
Xv	��-� ��m�]�&���iէ���?�`��yJ��F�ޗ�&�yx-,%��B�
�s.���)�CJM��	l/]��]��·N�Y��ׯC͙�bt$80�V.�P�J�%,���e�]Y�ɸf7"V���PC�q�/i-�-���%��`kC4�iT#��EQ��*�df�A�WQ�&�)͋)(���x��9�V�E��6e��V۠��Ӄ��*̣�+�]�x5fB�h�eM��DY�5[1$M	id,�TvUƞ�L�x�Ta��!I!�C���cwoV��c2Tx������S%�RJ��sbn�6��)Ѽ7��P0R����Ų��u�
�ZY��3F�Gv5\"� -g��Ћoe�iQ-�s�h�F�a�;V��d,��Y�\l�U�u�(��E-�j%��f72���El�M�0�'N�`LD'-�^��İ�j���*�[R�J4�ϡ�1D�
���UzM�܇"�A/1[�p� �� Ӹ��ڍ4u\��3^���7x�Ah�Y�I�n������ɕ���*�r���S�a nb��ٷ�m�u��n�@����ux�b�;�^�le��F4m,ͧ��#0Tu��џCޘ�!����S��{#8��fA�[�,��R�r�0 Rm�$R�1|�1	Q:�$��?�݇m�e`���p�|��i�|u��A�*f�cFIv�{��H2�����Z�Bf�73QX���G���v�i�S*S�t�٭������ �U�D����Vn����t��?M� k[�V�&��F�M ��BT ���`��OX�S�ư��3^�N�܉�R�gJ���2}�/�yO
ıӖ5湙2U막�H*�G9Y(^�@�4;w����v����C1@�d6\VP�u��R�s����05\�*7)�ݷ������[z�c�Ze!��6Į�؋6XTi�D:Ï3.k&�j����Ң�,������D�Xq^F0�{��r	�f�ƷS*��z�-�<��"2�[%b���u1	
�5Y���n%�ə*�&�~J,��� &2n��T��{\
T�X]��.MK2Z���(��mlC���A�������Ω�e��Щ $�L�WW����#���9q�Ɏ�z��q]�4HJ��5(c�L��C�7C'�>�׺G0��:�7�Й��@n�s%��ĕm���J�$��H71}vӛ��M�R�[�f���n<ɮ[x��U�5eE�Z4�z�ê��(�ϵ*���We�r�%���B������$"y�ZM�j-x��m�h$�.Pp�$��~J��fC ��1*VU,вX�kl��!�f����ˋV֖>H�b�<(��f̈c�NF�:kZt�0^ڬD�i2(���ܙ�E�^����7�]K�"m^,M�'t:E�+^�V`[�tCOwm��d�c�B�V�mX��S[eܔ����m����ɇ�;Q�P½���`C}4�X&R��v�kU��(fZ�ŤC�l(�I��E��x|�V�b
��GA�,I��[�Uzv&I����+&"���t�Ǻjء�*ΑZ�"�
Ǎ����ԃS`������ƬK�{cr��nI�Ц.+Q��x�	u$�vwr��orJ��In��ǩ�8�Ci3+~F���i�\�]��k2T6DP|cXy[��3P�j��Xac�y�TL�<6�È"�ا����P�3�jǸѰ^	��`��M�U�U�ԩ����Vn7�s'�i.5��9YÙ���g[�Զ�Gb�U��f��E���a2��5��泘,@�$&�Haq^�m�����8$n�R5Z˴F�o�-x��l�1��v4*˂	>�������6Ցx#�,V˺�M�!Βy�mk�5���swf��'Fisj2c���չyxE9c;��r���_Q$�/Y��*,�t �c�{w�p����$�t��F���9'ʢ̺M*�4�¬:���X��N�\��'�cj�ݹ�X-�:(J��M�����ݧ)��whXj0�--�7a�ˍ��p��b��ۛ&�f�7XF`���[����T�+�6�m�إ��7{2�Y
i��=I圃"��PCm��Ҳ�Q(�vD�"�����-*��Efwe�x>s`6�&��*v�"q}��S:�#$݌In]����ÊLˋKz����Z�]K"�,��6e���bH�^�z�'{��@�YY!AQ"�V	I4APF
�ے����
G�MMqV�Bb�����cX)��� ����M�"��ꬴ���2�;w��|00���)R�ov����K����LL��m5@�q,��Er�l��6���`G�4ԧa�Ux�[5�k3*�ތY�V������&��D74�:,��u� �Y�m�r�C]�P��An�-@�f�Vm^��I ��z�W>��C3kV��#(Q^��8AjJ(�Li�=�3B�G�I:���	2E8p�Y�I�LH�)Vn^�&�-��t]�n�f��X2�K�2V+��H�����$8Ȇ���"#����P�Y����l�8U+����xۙx�i��a�U��k]�/�j_����,xKa�*��n��eՌ���S1b��nDf8��wI���)�%�d؃S{�k\;��i�!�[�IZ��f�3X�-����&�h�]cj�R�Zaf%��Gl�z��M����Ù�&�fVPVY�/u(�I�������$I�@ ��v�Օ��Mkx����0YI�,q,��(\Sв�m&��+d�Q;�,7�M^J���V���@aBL�b��M),J����۵.S�CM�#0<�4��q�v�Jo�,��do)#J���]��*P�ݜZ���a���r�ӈ^�J�9��0�wS�׌�Y� ���h'���e�lm^�V��h��$- FE.xPz�ca�YV�dD�Q`�he4��`���ګ�
�ifZ�R���K�mm��	F� Ȯ���J̩�����5�`=�6��W�#�؟C��"u<��)ޘ^J��>hX���N<�2��2�3s0�di������.bU���V�z���ch��r<�W�4� ��KqB �-���%%4i/X�P*n�՚c.�w1Q߆����QrRӣq�Zw ��	�7mU����bЍ�F*�4��IXA�";`�`��E�&�
NaX�ʵY3z2�F�KTf$�k6,vt�e]��)Z��(&nݲf6ۂ,��"�iˠV�t�qX>hD��ئ#͆`��$n��a�b�H�/"MܘFȢ�y���p��EU銢I�V �I�6��ɐ��5��`	2յ�Y0\1��t���rD[U��A�I���T�fʳb=�t��a�VSC.ةOVf]Ҋ�`Bج����Į[���R�����1�v�.%$�v�\
��7h�˰��׏M�4Qu�IIc&��ю�J9+/`��Q�[S�R������s�˻�`�e�0����s*ۀe�ĳ�Yg�Cz*r�� �N��i�,22��u�m�[���$�҅X�^��ո^�ޚA췶��G1�t�`v����[��"��!��[ٙ�D����G>=߲!��e�s4��,$JH,�v��:�B��z�ǩ6h�1ɧML�����%8��Ol:T�	�7�����T���hˢ�	t� "y�e�����0va�� u�k�-]����_h�u��,=��}#�٘6n�j�ɚ c��kF�Y��da�)�n�cw�GlD�j�Z���r��A�MK7C(��+^f��@�8�]��U�[�-�,[[I>����c-���b![fK�A<SN�XX����Q9��Q�
�#z��ZUU��ފ�WMhۨ%H��c�T"�6�P�1(�ءI���L�<�5%�bA��q�%�Fm�9�~{[f�a�j�f.Mv��<`D��~p��Ɠ��:���Y[��2��L�Ŵ>�Mi"+w��«$g]M++^��p-�Ƀ74#��P�7.M'��{W����XF��Ęp��h�*v��><}��	��t����Hr�Pöͪ�k(�.�	��R4�wJ'6�/*f�ܭi2��D9D�Y���X��b4�F�22��F)��N+gS6�	��&�yw��E5*�@4����76�.���/*����V\x��ݐ�-P�Y�e`��I-�q˺ɫrx2���3�k����x��(��-�;U��=��o��hc .��½:7�{ZO*s�No�L��$k�iLT;"�g|i��9�L��y���v�C�����CbҖ6����}.�Ov����t�k�e��4�z��y�y^G^�6��B%4������?Q˪J&��A�r�h��w����{F���a�)<��uq<�_Z��J����mB�P���!)s
��7��gA�^*��#��6�/ ��}C�ݹԪ
�Ad��#S�>�����R�뙄����7��h��g�$�@�RJ-U���B��|�4���7>���wè�t��;�.�X�]3m`\�Z7,!Z��r������_ ��v�~��Ѷ09}x91�y�>@kVw��6t��Q<�U�O��]M��������<c��a�6�;{��%��ҵ�Ū�/��l�ى[�����dM��؝/`�Ut6��[��n�2����0��]�QǸ5���4]�e�yfuO���%�[�G)5#���|�'c��X���x@�KZ��v4F&�ӏ#�@����O{��#Lq�QzT�-D/!R�f���5���-��!!Q�Y]��ܦ6��w`��\M��޷4�px�}�b�N��x�I�˲�!䯕;9���:���SsV�9�9Q<�9���;_-,���)#�7봹ջ| �q��&���P�z }�XoUΉVN̝�o�X���}N�w' ���]t��
����q�1o.���E\ʵP}״g�h�ަ �QK<�+FK�g:"��{3����㗍��ՕQ�r�_�E�:��-��q�(ԑP��K��&�0y���b�9慻���t:�7��o>���㾠��{�|�㚌�+��L�w^X�
�P��f��sv�*��W���K؋ZI�Vp�j�
/O&�Z�6E�;Z�C����Ĺ'jdv��
�BQ���Wr�TፗR�͵Z�7؞�v/��ֻ�ʎa�e;<C��)k;25êr��&�⢐g<�kZW{������s1�T�ozR5�t`�+�:c���ʘY�}|r����A���(&�a��0u�o�E��ݖ�x�Fj�:��fZ�39�M-�'Ê�@'wm�;���2�HXeb�;��<6���[�p_xۏ����	sk_D�
[���G�<u���Ī��r�3(�8���kE�h)՜�E��j��Λ���H&gz�����=��������g��K2~�$�n`�+ה�L�v�	vM���P��؆cɢ��Q	0b9i�:Ɉ1�k�[��r5T^�g���^���X�0�hn��w�d[3�Jۮ4�[0ᰦ�ư�*l�|GN�ݛ��M�R&	����dmE��v,.�aɣ����]}��Ƙ�c� ����_6N��9k왊W�>�I������ܠ���x	@����.��d���;�"��v����]��6�rWP�l�25�v�)�V�G��RL*=�"#��j�F���/w�g�c�<���JA�S���:�33�Fv�S�ItW%��O�Q���^M��vS����,�k(Z$�Xǵ#Ώz��&�M\��]5}y�4��Y}{whM%���,ɹK=%������t�{����Yۮ�G$u� ��XS��ƋuLd��Bb�{&r<��j����6	��̤2о�������	9��Of�}�E	�Ǹw,R�,����s#�Νf��z��u�.�����[F^=]�^-�����k-��
���;Vb�f,S�����t%�"�B�"�Z�SWb��r&����ryg,&Ua�}��Uպw:��<�T$1s������;�r^S��5s���°_^;\Lc:5�j�)u�9�n��{r����#��6rc���a��x����Nm��Z�KA���{�PI�k4ly��d�u�q.��+�ľ�����k7�`��A#�j��O�P��f�XMEoo�r�*�{��n�Ǒ�jI������م��a�j%
��7$�'�eJ�wa�v�ڌ��%���47-t��gƝ�Z��$��UJ�ާ�-����j��S4CN|fcq�8�ckT�=Z2����'�03��xN�ք;�K�aYcs �a�p�ؼ�_zOz٭t(�=���8��}7ii���z�K��c���+֯4Y�s���t�W_���y��첗N4�"yx�3�z�
W��lŪ+Ζ��K<���8�m�X
$��br�"n.6����;4�7��)�KT$|nk�i�BI��T�u�-�+�A튺��<I�w�e&���.�Q��{9���o%ς.V�:��`����o�h��t�tl'����[�r͞�9����m�Ol�2�,��ˀ�}�b���2��^�Q2��Ԩ�A S�˻���n!N9���Ol�;���%@C��ʃ��]��j9�@��������;Dp{|z���q𹳻�9�������n�b\�Ќ�Y, %����rf��<o/Jv�6�^d�w��۾��H�A�kM�;i��`��Ws��㥍R���8S8't��3r��
ڶINˈP9p(9�P�$�O��>�%dSu�g�$��3e6��3�=�	k:��yx,���8T�����t9⧱��`\�ӝ�ڃ�"��Q���Pv
�p�������F�u�vd��f�OZ��\���-��s�u��+�2�����wd��m,���)��f���Fj#TS3�cԣ��;���ĥ�J��ft2젖.����7�/Q�ڷ9��>ώڱB�:��o/�\�Z�s�A�Oڽ罬��р�C��@��"2+�G�u:���T�����mSȗ�
*l���Y�ns�!� Z�4K{ٟAZ.�N�;˭zIv�DZjZ˹͊�򁮟p����t���l�\s�M骂�������iU�����m�[Ǚ��#g�A���P�.��,��3i ��
���Pl:K���f�%kCq��BdB;������� ��z�����ʼ��Ul��\;{)��مS!�55�'s�:�oI-�\�#-u�oV	��n�`I���8g���Z�{�׸-��F&��yR��W&�C��<r���{�d���R[gr�lz�Fj�r5�k�E]�GuN�T�@\��9���c���-_0;}V��n���噂�|��W��T���{[�lN�ݗ�����wH��7�t�c!���SU�HhO�#��vG�k9��G8��
v֮�-��9Wk�"��Get+>��;;���`\W�=��ݙ;C�cI��U��wW��ۥ�L������2���8Ƚ��;�_3Ai��r�R7������6d�}���:�U���%E��rri��N�1���-q�[+(e���R3�E˥:.��G+8b�Utd�iis��Ju�#�Z��N��5�M�Ǧ 3V�f�2i���<���p-_lG�ۗr�%y��{�!�L�1_#��+ۤ�ķ��I7�=}(�n�8�1��ts�!�]ڣ����ɛմ��K�ӳe˂�{w3�M�6.˓�Rޓ|/y��ٷeC�+��̵��`�r���Ү�܈�e��}�m x�3F�Ë A�{��<�����VWnc%6��2ǽ�]@rܢ#��xt�D���ep�8ܶ,���->�,����W�SY�Y����7�>�9D�F���՗���:��S�Ҝs-h���u!���9N�SҶLk}p�+�;Z�ڻc$�<6.瓧^%^�b��݆㕺��U�m���������Y��B����z����e�NB[�Rw��7mGw��n"���
��l�ޙ;��y�A0�h�2�����fs)�ќ�)8�'Z���Z��pt�,v5Q^Y������YA$̚(����0m@�j���:�+�e�B�k��͖�H�ͩ����w��A��V���س�S郭绣�!>��n�C�m��iK��ԱWۄd
_A�����]�OgjY�8�W�����Į��l�W�M;����f��۳��hVE��h�.��0�Z�>���0AQ,��5��]Is;����F�j���������0a��P��+�D�ʱ��;���"�4��
�#-�fJ=�zw=!�kN��D���0��� [V�C���'T�Ld�rw�g��&���5�b��7��gyE��؂R�i��gN�Vm`�^s+���1���E|d[�`�z��'#�9Fvv�F2�t�e*i��ȳ���p�3��.9��Q��j��]]�|1�ma�tr�,|�6���Z���*�H�V���X\���Wӄ[��e1�KD�v�7��يŉӇں��7��s\J}(���R�DUvc���Dgn�`�3ơ J�
`�����.��j�*a1X��{��Ƅ�h�Zͧ�+y>a-�]���n]p]��C1��&���Y����7��ov��W�Mno�u蝋�t�rϴJ�]����pZ
�� D�Փ�px,
��軛�4���Fjh�D��s;�ܸ�5AS"秪3v+��3w�5�4�^.]E��"1�>���z� �`�sz������w;���7ydh}�kW(V�<���f��\o���y�㤰Y6�%ؓ������V�7F.�w��r�7Ȼ��[ʎǧ=�8��Km��:���M�'Q�sv��	�����=`���@��ݟ��z����c�p����{�%��#r\wnWsO8�L#7gD�����Z��Y���P[����i�D=���)�� �M�7��>�B98/p�y�R�|4rS�)zr���vZ� Y�A��&����Q�d���6����%��sGb�{ے�T�\��P���*��R�e�zC�N�ՅC9��3.�Q_R�D�L^�9|Z�]e�g F��R]�)�6ۻ-پ�e����V�i�g^�O3.jG�([��32�z�s�=�P/;��ur��}fȍ���7x�̀��!�#�N�S��,�щK�(j	���w6�]�]9��}.f�&�^a�(S��I�^Lm��+ef6���ly�1!2��Qœ�TED[��z�ǎhZ�S�oq���(6����)���(��(t۴�6rN9�.e���艣�����9�ڒ��
ԏІZi�[�
��r�g�n�	�ka�[��d�����߹m��غ��xr{ވ��C�]��;���*�1)@��R1�Q�B�Ǽ�e�9���֌�����̆��H�	�l��I�S��om����]�l���H���u�=w�-Ý��6�ۊ�\��{��N&b0�G�<ׂ����rk�{,�u֧n�{C���zٰd��r�>r<F�ٲ����o���3A�Z��9�|6�u-�~��o`�/��o��(}����4޶��7]����l�':E&��R���ܸyS#�qO��A�hu�I���Ӳoe_ 4��ݠӑ�oI�B��x�C}�P#4̒[��ה!�0D�On �o�v}�v�ASg����VztC:E��J98��sX�w�QT�8��ls��\�1M�Z��Ӥ�Z3-ҰÖ�-�4Q�@SY�`<��zJk�+빏:ӗ����
���]�r��bO]���d]��2����|������l٬����&8��7F�6"��Yis�r�Vf2���#��),pi|�j�:�������7ک6l�Yi�M ��4ba6O�o��A�ȩ�,����h���H��Ȃ�v���3�C��+q�o¬j�2ܻϕ�[R>@�ڸ&��1�ac:����;s��y{���<�c��ûs�;8� S����nU�K�B�j�0<	ꆩ���*�3`���2�ڛ���Xnsj���K�I�T�Nv���꿳�_S��ȵ�
!�<��.�v��;:��\#�mvܔ�yu,���v����stBjL��Q��]]�v�m�y�
��*v
iw���wJ�"5�� �k��w% F�����F�HM�N��1���]*��Y1��:��}y�C6Z���r��ոA)��@��Cն�ҧl��i�_���@�wj���C��у�	��~�}}P^�ש;���f�*�Z#[Dn*G��֐r�d;��6�0��Ń<{�|��R���V�l��oS٫!YKE\�dPUz�ŵ���RE�G'q]���0�KA�y���;V_����G���|k�- r'�s�5��A�;{`]�K�����jSx�]ؐ�����R�&��s;�c��`SF���3�6Ոrs�Y�
�ۢ��v��kۓcJ[
�-ܲ�(�q���ɇ[cs!7�<7w	��f�����͐g2]Hiほ2�mNY݉is����>�(�7({}�f�Š(�|�U���w��;Y���jp�4o�PN��[�%��,q[�'���m��	(�b�DF��EIN�u�d��x�n1ω��x~ޯy.��s�ʕ���]i�אO����TTC]��+�����QV�w�WX7�XMY����DF������,�ЅJ1J>�)=3���,^a���������ї�f3�w�nF��4�N$1侍+9lff{;��žox���Nc��*�X�CR��>g"��Yׂ�v�9}�σ�5x�ܻ�STᖭ�����wpqe]����e˷����|��n�eK���T�J��?�^�����S�&�y�n���z���ڛl~��dO̓U7ѱ�4gHo^
1���u�i;t��R��A�YcBN�w}v��?e'�s��a{�М,d��^��Ѿg�E��<_&4c�Q��q�;����m.n�p�p���H�7k/�;r�e���t��gD�DVh/�f�ڳ�O^��\��~�|  ��?�����}�ˣ�Y��k��a\I��^і�?��JF�]O�G�X���A�f���G�t��5�0�f����}���Dp�ɽK �Nz��Hc�1�I�c���b���)l�L0��$kU&r�]�n����w`�Vb@|�RB�L�5`��ս3Kw�8,� ^N��6�t�%������u�s]ڄܾB��Cb��N�
��V����k��-B���YїR���4.���/uV�j� �ݗ�v���)T�aWr��^(�pjiX��쉅u�K�|��.r��bf933���/%w�#ǗJ��Zg���� q�����XG(��=���@o�6�p1���:e��%�8=�vһ�E�{<�����}8�-�-1��u;��_!�'����b��7D�M�q�{x�`����#W�T�=��B��VA�}xc}G��*�z�ł��5x�]�qz_+K"�9�=����S�tZ�z�?l�L��#�9�fp̶�.����삯_\���s�g�U�/+֤���bi|3vX���IP��r��db=c�i��Wo.����6��C,Xa��ga4@M�8WN���u��(����b�ض�K�L��e�iM�z�v��L��w��0`��ͱv�� �[K��h�5��˶Ě���x����'��t��3vi�3i-�X�ہ ӻ]J��{ֆk+�;h_(x��,V&����t�&�6ط8��ő����H�"!���
Q�լ�̩�ceګڧv���(�,Q�vo-U�e��N]گ]w=������Yh�[YF�$����Dj�+�9���h"G�.���=�k]J>�]	:�Fb$HW=�S3>�خ$�ӻh�k�[����e��[,�8Xl��y�L�F��Xh6uqJ曭�g)�^�s�Zo0gƣdޤ�κ��:�
��tD����cu ڻŖ�W^��vi�kVM���^��G��T�\����QS�\΃5^�(�|ҷ0�����������W���\ÙذƸ���X�{���<�4�癸Mc0ꅸ�n��s��f\��t �vgK�4<�bv]���9�wx��K��y>����c����ZGӟua*P��F;�N�T�%�nLn����o��
EU��p�G������U/�
���g�Ĳ=�.���:K��?k���W�(��7->n�B�㺺t���|����y�uh�0u�k���1��d\8�Fo{oT�{y������-��Ieiҟ�K�3&ajv"�[Ù���[��L��0>�8:,��]�]�7P;Gu����<�C�Q9�3�]4���.��#&q�+k�ܴ��U9{+��ܼ��*�Xg�v	F�\;���b��-�,�����a=��rk�YYy$�6��K.S�!t'$�³L��ko�t�ElX��[_[��M�6J��3w`��(�ZWo(q�2 Ep����i�3�v�u��X#o�$�o�� �7>�#�S�9�Y�;]G��@Ѩ��ߥH�m�a�B�k��X�vvl�3�Çf��@�`v��:GG���V+�/ypx�|�l����$������ۺ����N��W9��Um��6�^nH^�SBO]�DE�N�8ƵG����T=..�����F������}��q�4�]�]�]�!�:uKj�n�X����}1��Cz�wNGq�ˠ7+�i�k
��q�c�Z}ǉy� $z�v��^1]�c{�پ���[�8v4tjF��9�l��d�g_#A���(Ѳ0^�4�t�5"�$���+����V���̵u��^<��������R2�tZҮ�C��@�Lw+klU���V�p
���.u���c�������y�A�Ǡ��/g��f�]8�h)=��ؙ�O9�ߦr�.Ḽh��G�y��v��v�ظo$T9�yU��e<Ov
,%�HyZ���˥|�f��r[��FY6a��:K�%�MÝo�{���!� �f>|&(�:a�v�C'Am0쫜zjS�2�'�ك�2�.���*u�Z�Ұ�j��V ��מ=�ݧ�/kS�������.��Ku�g��h��(�:�ܮ��ל��w�9c5̅ha�Y����~m&�\����|�_l��3\#	a��.�ϛ�����&�V�Jj$ua;�����ʊ�
�ڴ�f����KTa�	��j�=�Mp<S�NR?���=�ڧfo����YI�*<˻�k�����{9�LX
�����ś�y��I�O�,�[t���P�{�憔V:�!о��u���*�B�x�U{������dr���R�+�
�<q�X�Z��E�qR�j�}�s����Z�LZ���]넝TT�Q�-^қ��(�O.�FGe�%)HXu�;��/l�e�|=��8�`k	�bus�I�� uŦ�R[`
jQ�b���֭6���]u�S\CXp]��_n޹�qaY�F�#�=η���d��!��Z�m���0b:����y�A2�g<ۜ�N�
ac��Ĵ�]%�80�j��c!��*qbI`�+��N�X�"��������هWތ��F{rk\y��_���TB��JbW������s��	�Z(��{�\��h��Kve.��ΎS��f�ۭ�+}�ARc.C�.�Η�X;�{���(uK�w�:q�ww��k���y��7�ea{��흗L
Mc�Fb���*�4��
t�g�Wr���VR#���v�O���-�n�e��4 ���ӌYw�b�{;�ӈ;e���ݎʁe[�}h�Pթy[�{k��LF+����(DtE��]�v�5t;�7���]��8��0���e*x�r�6)��w�1!Q�u�eEk&�����f�W5\��kyK
A)���G�je�sMs�ŝ������B�F`$�3d��Gv�}�5U�����
��mqY�\���8)��g9�M���{t��@���X��{A��J		�8n�e�ʏ�;��[3�f��%�j�ڒ��Y,�cJ*���R��"Kw	�����_C�H���ǵL��� �[���:`{��5٩5��H���޲$�,�ؤ�8�����tS%��^���V�ˢ��A���\�$V)gS�us�0mk��"R̭��=��ĥXڳ�#dݾ���CճTK#9Q�xK9���'
wѪ�J�N����n��tƀ�6�X�U=�ֶ�糵����k���\�'�:��C\�CM^fiW���=�s�[�����7%M�};�w"x
����D�g�C�s��߲K����+i۶�bx�Pb���wv��#-�w>�L�9��ʲ텚�qD��=�r��f�]i�@���u(��C�;�����JB�v�d�����6ҟٍ�`6��U]�C�h�̩��\��C��=�H��.C��<,�ݯ��w��U4T5��d�V�LfI;%�X1y kd���TM�s� ���Bl�5Yvw�x��g;-���>�&�4M�~��!�E�w��W�mʪ�Ѩ�'��ʑ�%��;LNGz�p"�{f�G�j�=!v�$,��d���j�Vi[�`�@z�
�r��[k��ދ��f"���MR��E�<��׺��bՐ���t�A ���U���A��(�S���[�����L5���.�zs2�q^�/�k���j
�}����W�/��o�6lX���+y�m��H���L�;���:���y{��.g{��������r^l��98�M��-�.�� ����-��1k��)=γX��yt؊㲸�w�g�z�Q�
��4e7�.���&�*��2'	�@{Da�|>Z;�/f@�_�Aݚ��6K�5+F#��E*�.�o�u��)B���-!�a����������Ҋ����C(���gwRٽ�اd��A���D�˦�QD��{�'���8Y��Nu�=�j:Cr�'Q�yN�.���$½��{&C�g���GmtF0C�H>����9L�9���������+?9����Uǅ4M˵և۴�3W`}6dtЭ�nnb�y�fL�gx���Bp��թ�c����aYr0�G#j�\�r}���l��	v⍾��VT����Y���3������2�C"�j�����he�ץ�(�ͣ4����,��"8>��	�D��j\����,���m��v�����((�F�L�˫��}�=W�=�vUI�����
����Do{i��t�٦��+����;t���^��!a|��b��7Er���!K��6��K{F������MU"˫(G-�$��뽊����u$�.n�{�k�)cY�WL��X+���s��X�u����s�+ӀK/j���ܱ쮫�{�[���'lN��ON��.@�{���vv�u{2{3��]������(:���ف�a��+m�s�Ve.��zɖ�x��ڶ�(��\ѵ EY�f�p������Xq�gnP�vop���C��q���<�`g�ݚ�g��E.Iف�$��}_H��i(�;r����ۧ��2����r]�n�<��E�YT�A6�#b�#6��͝Y����f˱��}.�"���ef�B�ͼ]�r�=���f���m^#�bpd#�v���:�e,ʛ8�:����X+X5tmnav*�=���B�쨍O��&	0Pn����Z�¸��]g_5�\6]�y�ێ��w�U�[K����=�5�>�W�U�em7\L�, ���q��t�B��&�6�1!��e�?Y�{��h偎|�p�w}A��Y� {�P�z[2�;=�2��Э��qn���AZ~T`(y�,��Tɵ����i<�̭j��f��Gym7" >g��N�.ѺPr�_}��L�f�L�v@N���h�X�QԾ��-|J�-��-q+Ȩ�+��f���w ��X���;;�^�oU��Y��#2�U�8�p�6«����!�6i`pֲ����B�r����j Q�W�RKo�x%�6���u)��ݜҽ*�b]�7Y%-tÚ�e��#ڬɉ���<Fp�ݵ���ǃ9��5�h{|��ps{S[���F��YB�V�ÑI�-oՑє즑�f+5��}�q�ۃ���Co9`�B`��� Cк�u�
���F�ݻʝt"�YZ�n+znV��61O)R��"���ݫ��]��	Kxh�@kr�pG�M��yJ�N�� H�+.�n�f�hv@��9�_aɼ̷�w�9���J:M�R}�QxՁ��At���1��5�Z�'@�_���c'15wy[��%{�Sķ�-�s8eM8�����V�i�'�0�kN2U��gt�n�3y�ՓM�~C�_��p���'$�`/����F��r7Gz/�]ν7�͇Tɦqh?i�6�J�R�~f�Xz��G Z�u� c�+��W�m^-w6x�X�X�b���7�����^�}��泗4؆3�v5ɡ<�P�x).
�@j=��eI�wkJ��>g��Y:F�ǻ_�{8v�(o 5�Q ��E,ev��'�{D=���Z�.!��#�Y#(�M�=��d_5q�����dɀ`y�Qچq�@�����k���YB����;���ZG����������@�55,환,�C,8��x�sb����s{�?��I�.;��B�ͳ�̹O��m�nǹ�w�T`���kI-s�Ō�_��������>�oZ��M���>�w*䊿A܁�r�v��mI��]�I��ߛz5�����}Ia���Vv����f���{���>p���2veG%
�U-Q�zs8�i2��	�ո�V��N��)u��5w+i�ګ�p<x�3���m[L��O�L�:-�v�LW0Y�ѣ�B9��4�]�!kx=����z�Ql3��8/"wd��y�jd��"|�uщ�Kxv�Ɏ��>��쭲kxq5{f�qz�>o0�%z��w��x�,��azԠ��c	���8v��9q��[�wt&U�8'/�y4S�0!.��]=�9�b��V����'�c^�Lǽ�(`�����۝��WJ��H�۸�ѩH\fB���*�
:��P�k�x����/�HoX���V�wnQZ�z*%-�/V�c�}��I��'����Q ��߲��+��{fg.�&��J�h��[M�����ɴX\J��ރ��:0��炸�K�iӝ����n���N�.C]�nJ��to�-w
&�%���߬s8b"�Z�i�Q$��ieN�Ϭ����me��@C�oŘǉx��'}5P��WP!��bņ8rd�B�;�]!г��Κæ��+g�3\�v_3 S^%���
���E���W�ZO�=�EX�:U�Gn��j�:I�X�Vx�2d���z�HE!�*�puO����%�T������y������u��b�r�LȟX|�sW�U�H�̎���v����z9�R�{��
WU�U�4�_7�9!��c~��h��t��z���_����[��S�\�,�=��P˹Z�m��i�a�����^A� ����֓�S,�
�#r�Su� �B���r�w����� �=YNv͆�0n'm�9v��Ḗ�3J\��[�����)�*{ǎ��P-yV��Lk���RZb�<�����y��^�|��՜}�e� V��ܒ�e�kp��6���\+Ua��V͕	Ŋ�A`,??��g����ȥg�3)D�2���iN�K��Z/�e��J�i��B���/A��mQQSojD>�.�Z��ڳx� `�zlVmf�D�="�O�	R�!_+nneڬ�q�E��'>kx*��%�t�����J��|�;5^��:l&��=8���4^��fǬ�5
߬�t�犫{�~����������kffe�|?z�7';��@��}�ztI�0�
n�655�s
ǘ/S ;��<<�K=��N�	]��;�;x�&sw|l_;s4tm�`T��{}�v[���޶ ��E3�e�+CWp�-�}9�pe�|�}�Q���ʒ�1h�9;S�0'Y��t�f�Y�v��N���Zǻ@A}�m�5ݛ6F�Uq�IQ�2�ěyL���cS�`�g+���A�M��J�tɞ��4��;xE�fݟT��G7L�a�P�	� ��ډ�=x���4r�Q`�4��S�f�Yo���Fsth��,���I�#G�U��t$d�V�nL<j�&�T�4B����A{e�1^�`�J�mL\����K60@4�ͩ�r�Z"���rS���wyh�ϙm��u@=���)���㕙�&��Ku�)5mA���x�j
��Rc!r�=�i��Ԩ.���6�a\_�Ũǧ�?1p�]/��u$ҷ��C�*\�c=g�Y��~�L�މ���1@�T�v���4+ǅ��ٝ���q�Q���Y�d^�̼�Ѧ����W�f��$�n�'�zh�,�u���B�b�1�^����V�����lr:�2�ܕw�P�Vlr玃���a@�]ħl\�T���gTj��Ӓ��%�0��k�-\�w�\~�F��3.�-掲�J�VC4�{�f��qg[�΅��°��w��n����
(|*�CLĠ0�R�Jlb���a�$�ߎ�� ����%3$�!(I�2�� 	w]&�]ɍ)���9���%L�F �3�$��d� ���(
�܂Q(�1a���`BI13&$�Rcr�#F!��f!`FA1�wI\��	*,�1���l�h4LӺ�AL��6$Ȯ�r	w]"w"�%":�H��!4��\�����.ss�P8�2fE!��٘����t̒#\�eD �"d"(�w]
0�A%���r��(��Q)!��Q�L�,�']s)i(H��$l2I1DX�wn��� 1���Bi�D\�A�Bh$��2"bY0�`L��L(��m�Qhc�wHID���1&A���'�f�����l�zhY�w(�<yZ��M}����d��/��;��+��8��x�:�{&�z���tZz�b[]�_��>�p�v�}�x�fG*;��B�Ev�E,ι[��� �~��dY��Ac�:�B��z��3E�B�������(=)��(v3�)\cn�w+:��ם[�[�!*&\CԵ���@�CuC/�}3va��,���}�ج��`1*	B�n������׋g���S�z�~5��(�s�l����[uX�]�P.2�<�5l׆�j�^dR�2��j�/Q7�g�.t�����aWn뿏�;�<�xI�<y�4�C5�ϊ�=f��\��E��KUc�
zx(U����C��M頍^�J^n��U�ߤ�%�xG2����9�av�S>8]�>���}'k��Z]>@=�� ��I��D<�#U�ϡkw7����/<�ۖ�[��s;qQ� �bJF��|D=9!@�1����itnl�wS{!�j�o�e����7��[�Le�]oC��|�JgA']%�*��u��zv=����7h�u���{E
�/��v�sT�_�G��y5P��)�eǌ�i �����.�ƫpp��輴��Ě%=u�:�����k9z�wL���tpf��r�=�&����L���~�4�2�Z�1:1�e�p�9�^�8U�f���o4��Ml�Җ�p�7��Ѡ�3���`��{���J����}��K���m7X���vj�LƳ{n��)0k�KJ�#�eZ�����xW�P�׌������k؊/C�5��~��Ƽ�L���� ;�k����	-���:=�'[��7p|m����nc[��P�8��5R��(^:�����0 ��
�7�{��8/+Y���&�=c�d�A
�{l�VO�Y 2\������0��z�N�>���;��;k�*�Q�j6��׹Y��1/�ɰ��wl�U~j�"�K���G��9M{N30���QZ#DjX��������~�)�N�h�r;���tTV����^�`�}*w�u� N�;���ӟ%B���OgY��!���#@�?l�����b�$ػ����Z��n�KJY�4$��_��zLՍ��a��_�|-�f��{����*-� }m�W���z�g�S��(e����^s+����Y)��5�+)=�0��L��uK���N�c�f=�Rx���Iw�)#��va9���.�c����G|N�U�	���\ۯ��s��'�/t�vu5u.��ӸWcXu<~X��.�ޮ�}�[Ư/�ɝhhX�hgu��u�opC2�ֲ���v��ئ��+�/,��X�vK)�Xr����m+��&]A���2:;�c��l���vi+�>��M�2q�i(��y�K���e��-�~��Eh"�ʓ}��]W�t��������KW�̃�����^��#!�|��K�[wcS�tU��J�X:SKڨ�b��z�\��;o���ܐ01��.�TD���'-��W٥ҙB%������Ϗ��%�̓{�k���
cԖ=����1]+�\c�Lf|X��5p�>�5��p=fC�^'
�;���x�o�r�P,P=�D�tkKxP�R����c���n�s�����-���{<�N��-�2�վEVPT{��w�K��{�$�Q�J�z}�f�$`N��^�{Y~wH�ո�gY�O��k�q }���ڽ���5^WA��C�Q�\E�9�<w�/}zT{ַK���	�/+M����ʑ<kG�B@�7�E:�{����H���)1߯c���}T/��:׶�ϋ��Ysl���M�3"�UD�_jDv��4��ބ��wүw�7���	�+f�}�CGDɏjN�6v@���7Q����=��TNΗX`*$�]�e���)��w�����0o�	��F�3��sY��֜Y�	�v��̦�:�^���w+�)Z��<���Ʃ��t��v�R�#�uc�1��m($��E)&�h�Ś�vz�J���x����>�g���s�g&����ݜ�)��z_*-[��y��k~^�d4�����X��=>b�Wt.!��nX�#?`͊�Z�W���=�L�f�=W��8�ʐ�Y��We��|,?�p�pT���]��e��m�S3�|��J��@ =�j`'��A�� ��W�ֳH��W�O���[����]{}
�l�|#5�>��7� dV���uq﷚C9D!}�&��(i3_}Ĳ$LY��XA�H�n�b�rUy�W_�{��L��~�b�3U��VM�ؙC+�~V��t]B{"����%fǩ��+~�Z>��u��)�g_�j�g��i�� �F�B;�tL��������]ԙa��i�>z���;`���=(E2�'r�܈wZ����H芬���@�2=l�av���h
�?{H:�%T��t�K�!�����8�c1���s'����=�o�?a�gz�}aX�߸�'YU���O���g�/�b#���Q�>z�9����7y|+��=��ыi�Y8�)��� x|�$i���N� ISSO��W�M%���e㚑A��%��'hǡ!�L�`��{jҼ^�B�Õ2�C��S�<<qѧ=DO���:n�۳�JǺ*w-�L:���q����d>�X�P��|�v��ч����#�˛��<�v�#Ŗz-Oi���"9�����E���ja��>�#�m�qN�����)���@ew*lգ�=Mm�̼Z�N-�p�ѱy�>~��	�u��.�n�^���cS����m�e��c�X��K�b��80j�и�0�@C}���N�Cj�8LZ&�w�.�g�c;ݵ�qO��[*����괈͢M8<����Iծ{���~���i/!�`y������zVF�zkR�����w����L;4� ��t�k�c5�j�p���\�ws��IKTH�{dE��Z�k��y�ְ���r_�ϼ��
�|�������qA��#��4ݕf D��zQצ�q�z�By����P=_7T2�{G�����l�k�u��~�V���]6{b�eoq��V��4z����e��dPǡ{M�Kb}m	�vEA���1b��dA2�3vg�7**��T�65���8M�d�&2��!������S�g {+Ng�z��j�ٷ��4�MX~T�U^�[���Y�~^;<�z�z�����}�]	��Y,�c/o�ӛ�X5�j��]�z���%��.v�76i��J�wȔ_��� �s>�*�S�x^[@dA����e`�C��1��M'(�>�L�ch�d/��h'��!�I���K׽�n.����4py�W�Zl@�{!�ތ6v:�dR죛L��W�ɣ����bׅ}�pV��ി� =���g�7�{ɻ�P�</��4y�y�fu�l˥��v�{���/s;sD A0w�3��}&��
�_|�T�@��H�qΨ�x�k��a��w�6b�*c-u����Hh$�6P���H�\��1�S<q���K����C�g�=o�5�e��|�l&��S6�ȁ��(�w`�wn��-��F�<��k} �@������Fժ�BE����z�xB�_�k���ש�g���-�V��8�n&|��P�2��00��ճY �7��ݳ�:yhˮ��&_�(�x��Uh�3F��ٝ�!�B��.��|$	��@T��0�Q��MR�/+Y��{o��h�yg����PD��`z�m���E�t��U��e3�s/��[xvv����G�T��K�%ōP���.7v�/�p�&!�<�ny���ӟ_#��>�lͿ��{*P�5�gi��G�߷�6���4u�@kȆk "���ua���"� �8��} ��r��"z��7:.��T�pA�������G�2>y���t� 'p�r�����`W⢌���_LZ���0w�#�����))}�f�{��cC�+7c<��J=��0�#;��>�t���eXD���@�FS�-�����t�^�ue�d���ˌwn��>�t�zVF$ӵ�����~rj!�p�Ԍ��Q�G�l$J%@�R��ک�։��p&0!��8�O���`�3_����T�'��bX��z5�A:��r��A�2�n����vk���_Å�n���yq�	c���o���oE�>��-g7���묇ݘ��Hؗ��'2]e��?���:G|N�U�U7�<3�&�=B�)m�X�]Mc�k�ɄɆ<�q�V��k+E�<x�p��-.��u��aϙ������}�m�#��5�"�:�F*���+2{Ҹ_�[:6Z:i��0�j�5yN;�#g�}���.�����m^��K.��-���_޲��L���l�v�ן�b�Z����}���\ԗ=%�Y4!\x�c��:c0��D&�o��a�9qyDFε��ۖRZ�!FÄ�2�@���U���Ѿ���O��֬��=/e�i�k�����vo^y�e����g��\k��j�gǹ�P\�d��7Q*R��һ�{9���1���5V�V_����?Vp�>�~����:Ol~�|_wb۵�[.�BCS!�����z�#cE�����r�x�����v8�:��q^���s��|����	�M�s�ߴ�0r
��b�y�_]C�M�nrXէ��r)���%8;��۷^ʻZ=���BuR�  B#�U�zS;X&��4zaz����E��cZ���xlCE}�`6��=q���LI(l��t*�xK��J�f����ݰ|��0�-��f4C��JblC�%y�H?�";E�W����Sf�c{q=���Lh��V��d���Ʌ�;,�9��w�Uɢ9��X2�L��PƍV�G~�����!|'Z'e᫃f���zWt.`9�� ;�z;{�Ws%�R�o�>w�J���tD��E^�Y�����+ט�X��+7�
=�ijM��G�{;e�ŋj��P�{��)��@�`��2�c�V�c.�ѷT���K�v�^�b��Cl�ϯC�%Ḇ�[�S�۞��1u�����b��Z��S�u�罪p`�"��Q��dL���Gy��鹺�Y�v��׊�͆/x_�$���%p��G�Z�=��K36�Fs~�<�}����!��x�&1V����`�#��I������;�=�:�ebVv׽�@ɉ�X̾#����Ԫ{'i��^��[���-�;�"(�*Y0Q抬�#Ŭ�+�(tn��\	N����Y3��o�	��ߛ���n�q�ǂI3�����s��ux;��ᛡ!ݳ0S��q�o�ji��}]�P��ͥ�R��`��V	�>LS�rv��{�x��+�X��ܶwև�a
��P��|��Z2�%��U�^��r>,P�G�Ҋ��SK�e>@Wv$8v��i���i��/����o�w����g��O��]����	9��_Q�
AH�L����	\Y���\	�eL�����/�R�\c���=�5���ъ#Ӑy:G@���Cø庙����]�_�<י�9�������s�
���B.S�z�`B����� 1���G��o}+3�\,�+�N�U��=�k2=z�m�;��E�L�7�!���U3AB��DϤ�����B�p�0%�hX d��4%�B� �����N�Cj�9Ţk���
��w����C����X�^T��D����#G��tW�MFJ}�B��7:KW���e��^�O9�M�s��a�&z�?�������iD�L��t�v�fS5�iպ�K��\�z ������Nը�O����.�`���`x�Fhe�`N��%\��G�a�����=�{s��P�YH��tU�����K�B��W��+z��F.���+H�W�ե��]�w^8i�WL�a�q$�M�O�˥[�&����ڛ�x�
�����1�`�|�FX�{K�0J����
I����}���,���k;Û��8���L·�]⧺�-g��pNz�hm��O�Oeߴy�+{͋�^�q)>> V�F.��|����D����y��>�<�������A�iT����5�C��/fv%�D���,o�A1�s'T�G�h�5�b-�S<��'P?PjF���U�s�^|����]�����~��o�s�<�M����3�m���h�c=fQ� ]���-(dE\��,XP��{M<���<��
�C�Yr����R������o�,w�Kn��8J��g�O�h�t� 6�=wu�u���i��P�7N"�j�ogE-��K��n�v׹�������9 :j"JF�3�����Q��-�
 F�~�n�7�&�py����'q	�6bW�?�]sD��z�O���t�^�]���6������1usdh�,gQ�����C/���=P��b�Ͳ���iIo��W��뚼�-4Y�k��q[@1����m�\T�j6�W�E"�x�i_k�㷓��n��f�D��������w��(W��S�xR��x$_Җ�B�:3S��G�f�N��n�,�Y���*�����`���g��wF�P�f�WI�M�b��Ɂ�F�M�������o�xxN�G9���s;��%��jޮ��e��Ɋ��jŇ�qg��E���v+b;@��}��+�U� "�f�����ur;�&G���rĈY��K�{Z�Tt�z�q��O�1lŗ�H��/iI�d�]pw$�~7F�W#7мM䏟�{�X���Cx�y}N�3\�[8��]L�l�_o�'Q�m"����5t�}uӋ��x�=�_>8��^�4?�mt;4��ǧS��/o�v�^�/F-ט�G0h�6�K�z+�	ZwX7p��=�(V��o�4����lf@T��M;[��i��k��>%��МO3�m�ϖFs�sւ�X�H3�a�u�˽��ф�%�ȈW��H�Ij��{ggvO>-<�5�9��D��7DJ���A1�9d�ڼ6�ij��z�ʘ�'���������t�fy��;s}�Qd�0��}b�7�R#qt��{�����y�1��D�z�z	0�D<�j#C�G�[;=��v���W�Ə3֎s��-,�Xz��-W�W2P=ˍmh#T;.1]ڕ���دYo�t���ԣ����.�a�z^�X~Kyvj��Y���*�`M��\b���w�2�i�e��6; �u���ӎڌ��
�tt,�j�0��Oz��-�������H�5;:�����ޅmy��
�>�׶wR+�B�IH2u��z��yF��tܕS�y5GL���#S�<�rp����[i�I;�c�0^���L��i.�<���{�,>�32����\�_2~3�8b����u�8��UcM�6��]~4��S����<շ1�Ļ�Ȏ*)/�L�F��S��|,�W������̺aӫm��v�M疑��]-k��\3�s�ۀ����A�,�me*��ش�b)u6�y��k5�-'_�k3Ƭ�5�ŭK�=�;�$и�	lf�������ٻ6���܊��ڱ���u��o�W���C��d�
�^s o=R�JǇ�<�Z�	�^��8l�:�����ۗ��#o-�k��4��������@�^𧦂��Uτ�����?�a��T��`u\F�(I4.�D�ܨB�ۙ'���N�l�`	�vq[z�[K˼ե8�:|��ʳ3ٱo#�8�L�Y���U2^L��=vc��A�'�>��*���ڀ��V�u��=�eg6%gNܻ_����\��Mz�Sʹ�-À]Ϸ�:�R�퉋�	[lf�����woR���E_3%����U�{�-&m��}�껸��O/JIw�:�DT����coT�]B�c`��<Sy��Ń{+(������Ӵ`]$�F�d����s/9ϼ�������-�(od�bS3�[�y�(��p����\oe階�J�ז{�<�Clջmܤ��v�	�I$��R���H����fBD� �RT�I&1��Z	 J)��	r�dHfgu�(�LE�K�Ή��dI�4$�F���Lw\�p1b�̂�DH��2��Y���4�!��Ɉ�r�I�fh��&RlAQb��Q#��wt�1HNW)�&��"�9�Q�&%HXfLD�e��bȄ+��DSII,Qd�	�$R1�D5��e�a�DD��1�IQ�#E.�Z$��m Gvᘁ�S�		ˤ�Bhؒ�]ۅ�p�h��s]���9��ۉ�B˺��Nv!3 �1����P��-�d��K��|@� w����o`)gT�����z�5a��v����VB�[7�n^4�-�&S1s]u͗daw�vh��&�w��xQ��w�?�[u�x׵������߫Š��y�H��x��������E�\�����;oj�r����_���[��:�6���ṷ*��������6�"|�$g�*���8�n*국�o�p.=|^}���rߪ��o�����k��wv��W���Z7������mϋ�{��s����㚻�W��~kϞ_Z�����[�{��/�_��Š�����1�~0��u�p��ԏ"Ͼ�u_��_o��~�}^�x��߾}^���y��߷}�گ����y����rߊ�̻���>>����p>�P>`A�[p���^7��_�F�W����:ƈlNa�����so�4���8���H��b$w��#�"4}#�u���k�����oJ毛�瞾u�����o���6����r�}~��[گ����y����r���{ҽ��{�o�B���"#�E����mWn��//^z�znoM���]��~�����������o�w�ߟ�������^���=o���o�~�>���okţ���׭���Ҽk�������|G�4FB�� ������B���(m9�h@�*W�_�l=�?�~}�.m�u}�����_��z��*�.��o׍�ۗﾷ������W���������?}����\�w���߽����ѿo��}m�nz\��ϾW�N�7ڽ>�X�a��2��M�yыO���x����~��z[�x��Ϟ[�r��^����h7�G?Z�W�O�z^,}_��(����y��_?{����7�˱�@�F)���'M}B�˥F<��:����JxZ��E��_�>=*�����{m�o_����_�z�������W⽭߽o�xߪ�W��yzZ7�~��~u���������W-�����x�-�늾.h#�"G�����T����gޞ�����r�����og���s��1_V��|m��~�Ͼ����_˥�}��[�6��u���*i��>@��B���W�*��ڽ7ſ^7�:����h���}^���]e�T"�u��W��_�y����e�����ѱ�~+����y�����y��V�W.m��������{os��{���_w����ו�\��u�o�z���6��~��{_���7�n��<��zx��x��0>� �@�>��/�7��պ��ڶ���PH���>wFf�b�J�e�A%�=y�P��{��n���	Ɉ��E~]�.m�yP�벩ay�#"�#��l}�j���PL�{1�ۉN����|�Y �c�B�7Ξ
�T.x�u�E��ͼ]wy"[����	~�J�~o���||���Q	v�ϋ�������������?|��W�-��~��U�iݫ����^7��^/�{^?/�|�龯�x�/߿�W���W���n{k�^5���=|��K�oV������zkA�w��H���>B��ѯվ]��W�kμm��k{�z�W����d�E��x9��""7� C������>�js}��Dh��w֮&1�<����\�>q��8 \1o��{�:�u�W���sx����k��<���x�����Kz|j�x�DB�G��k���G� �9����x}�s?A<~���G�=t1o:��EN�״{���N��|c퉁��p� �L�����+�ţ}?����7�����EDW����i���ߝ��oj�r����zo�;o~^����o����G�",G�(Ð�^J~<Ҏ��Y�Em��h�|G�ҧ�b8}�>��lwLZ�\�6�^~_�}Z��+�����/>u�oM��W�]����W��^76���p�j�9^���ίkN�{����.D�B>�蜿u}�����_]$7�#�7��׋���|�o��h��>}�oo�|W���o?:�c���ϗ�}U����n���=}p �>����Y�_!@��ǟ:�=��{m�x����~W����񈏅z�G{ӳR����m�ڗ��׶���w�~���}[�x���_�⿮��z�^-��|����_�NzT� 0>� ���� ��� ����T ���\t}��@>��P>�Q�>�q;;y��úޒuw� �W�w�{W������nU�������szm�wv�v߭�~��7׋�����{�s|[�z���{oKţ���/�}_�x�W���}yoJ�����w�7����4p��q��y�[�!|�U˗����[����5�v��-�^�����Z{����m�o��ߞ�_�������<�|\�m���}�~-���m��`��Ac���$��
B>��{��>|s(f���o�4|��~���+��M��5PW�	����`����5�����|_�~w�/�߫Ţ��u�oOֿU�_��^|�叫�����U�D}�q�c�
#�Z�
�d��^���c+v�
ˢռQ'9"��e��u``��eE+�핥�"������YLڵĝ��(`a��0({x�oin�;;�����Ut6�/�$�r8Į�X��z��ܼo��z�Lڽ�ý.��.��^�!�b��ˇ����D�� ��-ꈱ}�f+����/�z~�?�~���{m�{�����mzk�����^����_��ֹ����_�ο��/kF��߭龴�L}���1�p��	��:mH�5.�*���f�c���h���ܭ}�"8\���^�k�����_��>������j��>�����q�z��>���x�^�ޛ����^�r�;o���y�& �$82>>���^X�2�Y�����Z��������#��,�����H׍�^/�_����W�_�O�����|��"?}��k?}"3�c�^ւ�/ߝ�_�o��W��|���� �G�b#H�}�G�.נ����'������_��ƾ����5��<~6����\������v��ҿ�s}m��}����" C*��q`| ������}_Z�|n����hߋ����~-�">��4�o��YJp��Q�H��禿��=�r�����;^�}\ߍ{��=v�6�W����_[z���ou��z\�������齶��o�����}�z��o1����������p�|�­_����n� ����:�7�~�������}�|�������^5����k��=^v->u���<�?�{U�s~{��^���o�����G�~���X��D�|Y��W�p�x}�zZ�wO$=���M�K/��/�o����m����]��_}������x����~+��Z�����5��o����v��x׍��yޖ�b/.���W�O��w��oM��o~W�^^��p���?}3���x��Խ���&� \	����y�靖��	���������5����ڮ\�6�<~_�|��{U�s��o�����5��?�W��oKϝ�����ݷ�����]W��ۻ��v���@ G���.�7GwJ���}W�W�^��5~<o��׋����տ��h������r�[�x���^�n|k��4rH��__r���1󏮺D^����H�����\��*�v�b~;�lyh:�WP F�B=�������ݶc>&�_�Cs���;�f��[��J3���}�F3piי��9��_��;!-�Ҳ�iU�R�?{�މ��6q	����<�lc}�*M,�oI63�3�|1�9P{ܢk2[w;@��f�ub&���s����T�2)�^WS�8�w]�3l���46�����+�VF�}__�*���W�X]+ b{�*�7+V�jv��e����J%���e�C�f�B�W3�nW����G~�Ɍ�b�Gi��Iծ{��o���k�nn���vޠ�ˑ�@/S�o՟�]���Q����2��Mv�f3^���%��cK3F���x,Λ���x��TX�X!2���2-|�a�1���W ��/�-Ye������6�Vyz�~�h��"�Ct�������Q�}g" 5��ع���J +F�n>>8s���6�}П1>�,|.S]��}��L�>���k#�zq�[�hLn���a��C�oӺ�\��z�p��c#W�����r�Pon�U^js�W��)\5�5����/��{���^�
��@]����ݧ�Ӊٔ�x��
���,Ow�_J~��y~�(Ǹė'&�Ωý�M�@g��~�È@s��٠���Z_ϐ�U��L�����7��X��Y�57� W�ql�yLF�:�k+����ۨ����=ŕ��+�b���>�rX��#�c^�}�[�,34���G��&Xe�ݶeb�C�]���;W%޿I�}:������0���+u׋�{<,���c~���Fƴ�V�S�W�n���X�N������`�9sJAY8@P@���[ZE�`�W ������$|�����q�؏�R�\C�3�ݥ������l���S*�F�v��jS:	:�, ��S3'�So#�׋�3�rH��%F��f����2�s��<��cTͲ���)�&6�/�c�v�K`)�H!�4�:@;�b�cY�V��	,k�[�ƹ;q���PPʁ�X��wk�0�&������5�h�Ҵ@� Qž��p�����}(t�ыƶ�$�
�3��T���/}����?&`��D@j����
�cV&�7�  P�ܤ�"��[���޿n�VSf20��u�/�w�>(!�E�@r�y�2��Ә�W�Un��L�{��:����b�\CUJnt��0E�,	n킦i�ǁ����^����׾�|Ͷ�5T�,S��G�o�����%�"��)�F�t��� ��(sA��vVja+"�O�y��x�|���.��^����v\����T�����%����҇�Y��d�n���
�ZF�|z�Z��AU�3
�8�_�G(�C�/�]!u!���{�
���7�5���_D��/�s�����9���ܝ�b�Q�φe�Kk�ʯR��]d�
����jz����u1{Is)-��{:���E>d&�F��·6�9^���lf�Ƶ�x�s�jظ^̛{In���B��}��Q����<�ܮ�ߔ5���8�����ֳ�V��{��5���p��p�z�rڻu{�]p���ҁXK9��{�n��5�>�Gm/�a9���#ؾ,�F���^L��q�w�ٛ�9ʀ}�y�^}\��;R���u�9.R�ע���C��jg��x1�|6�v4�WgQYBΈ��� LG�ֲ��f#޶��j�GF^I���ʃp���{N+*�n	P�\c�����=�Ɇ6�
�uˢ�l�v��YB��)����/�#6Bm\���
L�� �t
���D�׷�������Lf>#�+ލ�b�S��#k��C��u��3W
����� g�\��$���Ş.T��\�ҍsnp�" ��5jq�*��p�!\45۸yr�F���z�J�������	�z�(wva-mZX��W�+b\JwYWOO���8�a�BWЛk�}� 8U`g������o���̡2)�upA����~�!����\���AyX
n����X��P�%zr�ܸ!̛{,�51P�1j�ʯw�vi��˥9��ty����:�&�"i��BV�CP\��n[(=4v�Z�%Od\Xٺ�����.�v��ĝK���gR� V��c���1���	.7�rp�ZBǪ�)�*�ER��w�.��">r<ڰފ�>2tAJ��43�¨�[m.cC�����w��~,.�l !�~wwA�C�;�="�|1�|k��p�4�����GJ塣O���>7����d�)�O�m:Ό,�%�k�h"�k���~���m�E:����\�e�5������FT��n�^��9/L\ ��+��h�A���Q�f�p,��^Wf3½��|,�(���\�m0}�ɽ���)�7O�C4��m���ʑr	ڀl8��y�v{9�yok��[�/-�L����`�/� C��+�ׂ�f�^�l�	��5$�Fз�g=�C��f�G�K4 ��C,yJ�������K�W��
�pG�"�3Y��;��|�e��%�n�������R���'h��]k02"S���1�"��;��f{4�z�S�R}`w�o�{�Łx�n�+�?�����1G������\��X��]�^і�E�޽M�.8��{�|���0V�{��w/����K��H��B
�33\#+hl�**lXG�%�w�ۡ-�t�12��U��i+(�:��-.�)�]�vҡ� �$�4��m��e��Nq$_Hr� ��
!ў��$����rŇj�z�H�6g����5��.���`|����VELH2u!�DG�}n�n^�c6�h�_c������r��(
>GI;Fc��H��|
c��0w���۟Sq�0{ŋ���Jg|�3�t�{HnC����=9 7��JԪV��Y�מ�q�*h������E���*��Cp�ڦZs�@�T[vF_���Y�s�G�q�s�2%�*KZV�*��2�@�j����wx<�%�l�~/�����Yb�@5�|�-��^�e�}���u+P b{�xJ3����8dF�#�l۲�7P��v����n[����Ҕ柙�jDwQ�i��P�4��p���Gmo�PO�vڞ���_�g�{҉N��@��右�7N����0�t�v�f|�xZ�V_{�ǜN��7��2B��<��^�?#����`�!�r��y�dY�����V�MA��2V�%�[�~�}�>�l�����5aV�u�w�a��0<��� +��b���O>> V��9�xz�g�)7X��e��_s���ƻ	�+��q�f�~1k�+Yȏ:�'r=Q#v�n���.M���a��Hp},����s5av�X+�-u�J���k]���Ah`����<!�*��Zy�/r�nV�%Y��m[v�x���y��s��J�,3PF`�z�lx�K{]4�'�Q�7��]��d���Q0�9tD}�}�U�+po�F��b�!�'��g�y�����b���5:�g���h;���n�ݿS��QI��n�e�fW�\½����)��"� ��	�:�:���3�H�D���fQ�������[-����\3�xT�X�}��~�^��7����E˟`a`	�t����b6�V�c^��{�ۚ 	��X���y�X�5g�{3b��?d"�z���]Q��N��vP÷^j��4t�����h���	"j���P���cQHģ5����r~9?!����m��&�����~�&��}��x�!�W�IL\T�k6�W�E"���ik��u����v}s������yK]�|��b�����@�eh���}��²����9��Y�h�Q7���K��-��^m�V�l��0#p��QE����<��b��X���妷W� �~J�p^V����7�E��҅8h�;H�Q�=d+�� �n���Iԯ{����Ӗao��ad�ӶL�޴�ݞ�f.���o�V�^��+�t癷��n�R
PT���e��Z)V��A��uf��97x��V���_l͙+�#;�o�4z�� �ީ���`�Z���8wr�F�#{|rMw~�����{">�L��7�~bw<*�rk��h/ :���@�'��ss�T�]����JT3f�`�������=o�G8�9����w���̏F�L�6۠5Û�DPS�&��{�xN��z���A����?\�X+
���˄���
��&�� =��=�%�qa����{�l���1w���5U�U�f�f�����ef�No��ՊEI�>�T���ϡ]w��WXS��{�8����EVƫr�u�|���ʻ�kS�B�퇵�}-���������l���m}��H�S��erC�~+�B�9B��#�3����'�0����S3\�[���{��+�^�5� ��"\5&s�;�z1�y��%
}3���=5�@������~C7�,G��B��:�	;�V�6�v���,׉�KƗ�T��C6��e�t�x�3+����^<~j��W��ֶ)�M�.�>������z�:�P��药nM��*P����l�V�������}V�l��l'ۊ`ʻVv�5(en]��8�[�շ�5I-��sk	٘A�� i�E����>��b�=cOK<i��W-�#c�Qk�p!�8n���誺4k9ov��6ݣ��{����޻L�R��Wh/����M˽ޱ(�ko�3�6�s2�m%�+:��G?/���뗮Ї���+��#T����j�6�^�WJ� �����đ]���A1h^��k혌���#�t���G#;2;7n��Hm^ �TX���[��AM�W7
7���9���lX��6�>���Uw&]+\��=��J#w��q��2�N&�����Eh\k�{�F�¶�j�=☏Vxq̅�1��gÔ(��iW!�P�0�Yh���(���k��x���c�6/�ƛwf#gM���4�򢯵9N����.z������
�zۨ�ab}�T��������25�mh����%���;���9Xb��C�t�dn4�7a�
�E�R\��*L�q�e��K
�NД-��t ]�)���䩧C����h�_A�Ρ��"9Sn�.%z-���W��Φ.�<�n��&h�W�B�s�Y�f�D�R^�۩}Ye+@���c	i��:$}v.�/Z�&������痖%8C����2���:ٗ�;���@�Q�<(�r.Uݓ&�e9��&֌R�3�O��˸���{w��Vݷ��͸���;��iu���[�B�$��Y���|��HH��4�))��މ�*ႁ�YN�*>����`����_�WBR���ʯt���ٚfG����J���W9U'�8ŝn?$|�*�ٞ&v��ڈ��z���lb�n��a���2*ۊ�Ђ���M��,Z'S�ّT�k@� �m\̂��:۲�E��t��ң64���!�u���b~�oN�,;�TyE��@�T���Y�6�&�3;FG��7�ùc�r]�1�M�V)���êڒ��}	�e����E(���n׉���
e/gzi쏠�@U��%��i,��FE��Y����W]�P�D�v�Y��&����V2{}�	p��J�6k�%�-OI�93̩=�u��q�(�u��1�N{ޖ�����I�Ύ0І��n��A��J�����%EHͥ����Q�ͭ�8�N
��ut�+{f�"����ŏ�\��ާ��O�s�$��w����w�@����j���D�{e���.��ٻx��8�o}p�̱Z�ٴ拮q
\1_N6�E�zEwXcVr^̧;�VՓK_H�^�z��ܐ�\,aJ��sZ�-}�6,�C����D�:�u'�n�D���jBzN��`v�E2�����֨�p�q.�������CP;J���WF%J�:��s�)��R}�@��Mv�E�-�W;�XlԼVGSKO��=��{������?�~�Գ0f0d$���"(� Pf��؈Ȉ))�(��jbL�T$��؂�
I)$�,ɘ�I LKD�&�]$�����Wuڈ帐Q1M1k��bKs�$� RH�Q!�M���t�F�"�(�4�a�,^5ه.�MfH��$ �Hd�c&RY���
+��l�ƹh�)F���2B���x�("��P؆<r�$1�4j&b  �7Qd�R`K�"o��K�ll��)d�d0X����fef$�b�hŹ��c�:d�
��la�	�A� ��Pl':Q�>��������.
�M>�2��tiX���H.^oz����
�ձ����������rl�=�l�E��d�@��}UU��\u��߱��@���JݾN��(d5���I<�P>��SJ�4������b��
��|Ր��a��xh�#�r��45۸x7*Q��ѪLǠ� �E_�y��)�Z՝^��cԯ�)�����3��7�`��5�T��� "<#�L�yll�H�#�Y���gjW�X�:�0�������.pCG ����ݑ���E�O^{ ��s�|��d�D�2v����_�� �43��մ�Q�h�,��Jbl
+wӿlZ��>s%���͑�GP��-ݬ��f�L�CG�N��x��5�Ӗ��?�w��!��8�L. �y���?Zut�5�@ދ��%���j.�VB�!{�w�4�|&�[�.sq*�ܠ���e��3�
��*k�2v(��@�a���a���?m�q�ZhJ~H����Xp6�t\B�V!y�f�6r[sB*R!�XՃ~�����q�^�'ɡО!�<��Ϫ��a՜�r�Oz����ɖ+�^�z�F.����u�bC_����������#m�N��۔^��33Lձ *�8Q�s�r�A���:)ζ��FƵ������#L��վ��:��f�n]"���z�b���Ϝ����sx�g��Ϧ&�J�i�(2��9�nr�D$ka/�}�G�}��3�ܚYg�78�ZL��	f���3�e���᡻��4�_��<�K'!.�ڴ����ոkD��=�\-�_s��6%>Cڰp|�|�y�]��$?JD�xy.>�P�O��
h�\+ϱ�A��H�u��	OɊt�;,�=�9�`��z��k��.i�;O/'J��Q�wZ��ji���M�4h�����4��S�p�X���N�9.>p�-:m[�A�k�8�c/��L=�w��WZ@8
4��&���_����>v�oR=��k�B���%Q�ˏq�"��"���l=��^��f_��ۯ;�z��{>� �I��R=/��)J^Œ⦀���	�ϖ/\Q=p�;+��/�������k}���[7&�̿X��/K��@Y�U$*��@�5�p!x�9�{��m��^�+�]��?�1WS�7�,�=��P��&�%smxϺ��1���|����6c��w���)��>2y�C����ͧ�1z�"��ӿ���q6�iѽ�Gu*i��_��N�p���{�]ݗ�ڼ��M\�ҩ���Y�������ۭf��!a����°�.�����B2!��K��!䃊j��(Ԛ����u�L���î+���M�(�����t ����cF��Uc@�$�`���P&�5����n�g;�+����d��� >}����]o�=�E�ħ�ͺ�\2�ƾ��?'L}Jn�2��}�kUk���xc(>^{�/�o2M�\\�@on�/3#Qxv/����FheÑ��k�rU��K����$�=�x{^��Mk�u��5��H*���ΐM�`s0h�}��v#ix�������t��y������qt�Y,�g�i�_?�Fz�������G|KiU�<������_{n�z�U�+�jٮ�Z�Қ���dܫ\���so����F�f<x�sB�����/M��z����օs��#������Ņ���g�{�#��Y�����Y�`#�,���_�ip�������f���!���d���-*�c|} 󙝽Wd=e�+ L{U&�)��uZ<<�W��5뫊�� A�;�#�Z!m�{7��^U��ƣB�/U0�K�+�'p�Ǽj}���-u���#Q�0r�@GS��=��,�	=�K C�u�M!��<7��1(�bv�u�ͅ���j�r���|���h�T3>j�g#�95�}��Pe��8�#zz5�8�(z�A �p6������UŤ��Nq��Y�s��3��z�<w.@�ֲ�vu��5Ƹ:�CZ'�����pu�wv��R��vk���څ��*�M.0}}�{�� \�8o
ĵߝ���O���FQ8��A���YM*�]9����g����fOa=�s�_�zck��8�C�Ja�z=u,ڂ�3�L �-��`�7�,X��>����u7ܠ�[�{�-{�� +�45�x}�s�,�ȈT@�<$�@W���e]F��wP�z��|�d�u�Z}Q���������@c_6��\KǑ �� /$x�+&i�0ٳ�����R����}���
�UC�_&�Ap��o�/zO+��j�a�ڣݪoֻo9�D|b�^.�i�ea�.�|��1#Q�M۠5�u�8b�|=7:�}hSZb�/U�}��K���.��ֻݗ+���#5+ؾ�([W��Z�H��D��OR���]�A���j�'�U�tk�l7��jVꍳ���&�ؤ��7�7%sjM�]����+�?{k{�8����Ea!\~���}j�B�o�,b���My������!3,�7�뜆��O�����{���c�C+���ǖ�۵��+����*f�S�z�(���.����:�f��ܺx=��{��B��E�{Ӯe�`�0�y��e���ٌ⡑��L&�;��g⫍�O\�x�L�&��#|�kX�u֝�nB�?.���uV9[���o��֬� �ƺN�U�U}_,1�E7��qR�s�� u��c"UC��[-��F���ey��G�hN·��������QZ�%�
�õV}CY<@Y�{�%�C�������JwC��{�#}*Zռ��ў���K��/l��J@�Pra��ªD���r�U߲��m��38�����>6�`�wg]/�u�W��
��-z'ͯo+�LWO���|��ʽ�~2��I|���+�08��/?��G��0�#�����i���I-�����������/U��r}�b�҅� V�q�B>�ƃ���p�nT��T���	��p�xxV��kܔ:�Yk���j��X�Ɣ��+D=��w��_�c��W]�ה� ��[�%�x*������<St*���@�Zk�����t���4p��7Dd��n4��������'��e�|HF��O�{���.��5εm�s��4C͢T�-����l�P?e�~�e{ْ�n�+[t��H��1�xׂ��j�x��:W-�;]�|�G������▛5�+��\i�ђ����c�}σ4g+Gv�.(�]`�-&��)��gu��(l���iW{�4�YySv�P*�0f�{�זpu�O�C1�3�,E�f�GfS�e	y�+}5έ!�F�\W�n�U*(���hbP+W��:���#菸�lrAO?3�G����{�4]��fr_k�!�K�ՉK���F�Y��'ʘ�SyV5M*e�{'�5�п���������蹁��,�أ|'�~����`Z�;!���3�z�K����[�^�����1���c�)^�b�{��)�Y�	�@��!�ߥ��=�2jV75�|ĺՋl���a�Y�.d�`�a��[�S�����p��2�i�z�8E���?rs�F�OatmX�iaϙ�%��~���_��a���/n��R����p��W�BަoOE�YD�-/c��t�f��=�j��
�����xU�1鹆ϰ�f�dQB���|w���H�ϼ\����ԛ�γ�X�8J~LS�rv}e1��0iվC�{\�\���i�\�vl�W~���:�x�'� �uSMw��Ӱ����(�|#K�A�>{ڳ[JL3}�y/z��t�����x�x3�8�c/0��|��J�г�pv�@џP�X1�]J���rz1�!~�W�Ϛ^��G�7_�o<��d�0;����ߝϽ(b���W�\�fi��L���ݲ���T���+�K�չJ��o{ �t;��W�d��G�;+-j�Ż�,��Ê���2����=�D<nh����V��<vz�ف����ŭ��Ѷ*Io����d
,*�p�������P�=�z�~���QQI~�"">��qY�H5�	�"��t}1F�_Q�)�X�qW�L��uax�~��"�F��or,�K��~}����7f�C�)��� 2��	�5�:"�/�u��%�l����N��5�t�^��t�j��VP^��}����� ��P�bc)������q���t��W:�8�߾x����{��?JS�~f}��( (֜EdN���Q��Vg�m��V�~��c�!�\�P��%�r��υ}`',}�n���b�D����{Z�]c-?��m�qF�Ɇ##�Yld$���"���>���.y4��^G��y�%�U�p����T{B�٠����"�kqA]+w�a��0<̫< �u�6,'Q�z<ل��oZ&�� ��Q�F���mg�Z���,�󂼅J����[ק��09)�μ��o����Y�	�f�6���j�~t�Y7*�s�+��Ղ��g2��y"��o��l|��u��=�e-u�0�o�B ��3!^��������ǭ���3m%�Jc�}���ty!�\�j�ߍ@��9w�ܚ�;�1��6s0��gw$&q�{L�em�Pb�d�z��;/\奩�W0���ŋW��ػ�k�h�f$&&�L����<;R�������%��.F0sT�9wv�������OZ���W6}~w�AM;��Tb:���כ,����B�����JJy�z������w-������z��J�� ��0��Jni<�#n!�h��Y_n5��+6��x��L.e����V�$�>��Ln��
�K�L,�.����	�'pه*X®�������c*gq�GX�6k��$����õ�F��NK���J3Q����r~9���ݫ~�^��J��#q���q�K���/�A X�ՠ�}ܪ|ҭ����;��
�%i;k�HT��;p�v[��&��S,� =��! *�^�`*�h.t.�z��afM�E�x���}�޿��Ώbu�M����(�?&`����|$	)P���wZ�cs���60fA�'���ՠγ��&�m׀���"n Ȑ�F�iVë�ͣ�H~Y��V(���*29��?!1��P�5T94���u��.�����0\�3�Y}�+���mW���Ѯr���|�2����C3�H�R�4n!�@k�$B��9�t��\�N�\a����2����<���Z;�&e�Hl^t�`7�;skgk3gl�H�{�Y���%�H;��Qza�ߵ~��fZk$�� z�aɛ�Z���!f�T<o7�����I�J����_��x�qX��k��n�4�2Q0_/������n��v^��``��c^�1xS K���.��Z�/v\�����/US��aֈ9x�X����E�����d�3�����B�vJ
�uא7��Jc� �37˹e�U�o�/QCD��+�^�0sʸ�{ҞMg�p�k�O�d�� �W0����	Ƭ�Uq���y������2:�4g��jv�{=�.�	��߶����Jc���,$�(s��Ĭ���̙J�~��`t��;p ��l𿹷^}ʼzln���ע�Zh��n����6�7^��,w��a���� ⭺|�*���Q}����~C7�,G�S��[-��}q#�gm�Q��ɣ�r��N���ti{U. hύ�����ڽ������1�u(;+�8�	�>V}(�����_�/M'(D�q[$��
��עSk���1]WƲ��th�}Z=2�А��h���:c3��GԚ�{�Ub1��@S�|�\��/*X+�M����K,>����T>Y�{��~���oFStݏYT��=�lK�0V�[�e ^Z�YN�e��Ь��1M�>���{�o�79s��`�>��x�2T|1nһ7Mp�4���2�t�dF�ȵ�3��j�u�r��E���H�B��3�[�y0���^���v��gp���<�V�t�jv��Q��K��������W�K������VTz�����*{��g��Q.�L�I3hB���{�JR���\�����l/n{�JiC�5�4���'v앯{
X�����ږ��Y�mL��3�Θ9����ȝ�Ξ�~��ktO�1�P�����^0�7ُ���1��%��H�a�~����H��^e�q�$�GQ��3ٲ�u�Ë{�Y���v�C�|=a{
��,�n]	�ۛ����g�8�Q�Jgb8sM��g*��t�ꁇ��-7:��<.�b~<��a��VG��h����������g���1?U��$z�Ga�C�Ͻ�xw`)U�7�<�%`��5�O��jq�o��o��ذ��k���`�*�O��֚�*��P�V�T��N�������Ynmj�v�'��9'�\��/��q���8�0o��8?
z��^&A�؈
a3�Y��7F��0&�硯R���X8�r)mMV�o��4������(3O��[�'Ӟc�
�'�;���#뜆N#��=��Wwң�Hf��w=�x�ٻ}غEԤ]+F粊T�'�m뙶��g�<�jP�19����Щ?^@�o�T�;�T�kV�O(3;�����̑Fba!�E9����@ �E'i�拧�)�ʠ(�V��6��Q�d�g���y����"8S;`෋�X���0{t� f�6��Ų�M �v�l]12����U�,Uu�4����tk����E����m��RK��]G';��f��Y()w�6Q�$T���M���mX����J��=i�C���l�@����
W�,5;8��(��w wv������_w Y�SV�d�K��NR��ɱv�p�d�Ѝ���U����|����É!�ZP��}*;��W9=i�iTii��P�a�/k���YՈ�F�ٜ�ܬ1�:P�[�MQ]B��l�#�!g��!-��ξe�/K云s-®����kM�¯r�T�1p�@6�Lq�ct�.|{�]��i&�m�)�,S(gB����o��J�ɭUډ�<Sc�%JAw�4�AܺɅ�w�񗚑�KЍ�3)]�8�8��5)��93��HV��پ���5�5�{��\{��Y;�Z']��/����	O�/j�%��(>/�o�.������7����#4�p�� ��˰�q��^ޣ݁{�+�o9��XQU2l�Y	�tX)^��X[�����;����Me�����t��w��v�Z^f��#ݽ�3�����84U̰�>��*ݪ�]�z�gd�/w�dA��k[K�7tիx��Y�]v`xp[�ԅ�+rP�� �W�ؿ����4���u4��Y'hҮ�ǂp�|�ٰ�9,`�P���YX_(�r<���������"Kz%sw���a�n�X$E�{=1��YĨ�\�%��s,e�o�1��x*پZ�7�mk0���s�Q,��T� �R��i%\�u�q�U���cqy������ĥ�V6�щR��
�Z[|��H��c�k�=��3E�J��,�ҸB�
*WXï�����B��ə�°��n�X�6�^�J��wN=��,��z�y��v�b�� �;�,�D��� 7�jFYw_��ë{����	C���g��l骩l�����w#ᦽSP�5:�>�o��8c�A�o��ռ8y��\�TQ=-��W2]ɝ&"y=��)G�i����K���B_"�U<���9m��Pn��|��r�E��kYSf%Cq��� fj��2�a�y��9[��;��ˀ�Cd��a��hw ���u!G$�3*�vb&-���z-�I��A��l����в��b����o#˅�$w���~}�����<�McL��"��cKII~:2�d��т64�5�CD�QT��,X��(4�h�&"��b�S
#DjMEJY�nTQ�1�U�r�Ia�EwtX�I�Ō��X$�`���C�s�I�D��FŐ
���Ik��d����b�1����QL�*
)�r�b������QDf��&��(�h�.nZ+2��ܱ6�g�PN^5=w]2�����/��1c�\��fݷg�ޖ�5����'����7�íU�Yڭ˨�ky���������:f�����J��?���ϼ���<��7&��a��{&��]a7�8ѻ�i8��YsW���~�i�ϝ���~����Mzv�@����Vz����y^�X��B���5���j�Ż����6��'�*�X�_-X�&q^��u�X�4ȩ�-��)T��Q9{���F�э[�t6kt�VA���7��]�&��eqc��0�	*����W>)Dg/tT�I�bt.̓�$<�~;��ꆮ��vP�/��=1�<���ƨ{��Ꮽ|�ٍ,~��ȗ;���=�O۾ͮ�>��O<9���}1�/�-B���:�5W��P����hT&�(�f�L����/9�����Յ������QK�wޮ��M�k��c��%:b�۝韎N���;��V�ٝ�:nn�r��c嚹c~�i*����Mǝ�6�\n�]�3��+򫆅v��������w�5�.�塍l*��5c�Śy<��OE��іJ��w�t�� K�=�1��'c��8pʾ�"-��Q\�Pv!�|Qi�r�==�:%u��䜝��u�3�É�y-�tq��T���?}��U���7�P���i�u��b*���W,�����>���i�U�4�Xˡ��rC�<�*2l���Үe�M��k<��e)�Y���5;oxYHy��:]�3��^����8�U���*���絜�j�w�YEj�^��k��㞯L�������qﲣd�vx=U��Cm���׫7��>GϏ���(Q}/~���yt]�!��6���:n-F�2�F��e�,5F{~�8���!g���cړs���o�5���N�$��LS�gS��8����/jTj^-o���	;�6��'�wS�B���/^F1���������r�m_N"�����]��^��;��3�4ko��c/��Ǹ�֦۸����}�&J�N�q�7R�}����8�^������TE�P�7p=e���(P=�e�e��|s������чr�e�(���d�<g��陮�\н��x�Ňt�Nh̬�3�Q3N��aw����1��7F5����#�g"ge!��G�����1�6�6�1����hǍ|���0�<)��̻ޚ��3�a�������868��������m	�ۈ
��!?xW����%�)���G���s���o;J����K��>���_<�g���Aߛ�v<�Ȩ.�D��"��'|2�v�*fv�����ٹ�#W�ʨ�U��oC�H&��y+�l�̵7������a�k�i��cT}�G�陞�Kju&$d)�"�9��'�;�yǭg�gS~�k���}����9C�F���W�NN���u+qS������3��ײ�u��&�z��9OFDǜ��_]�g����	2�o"B�w�=ޙ�۹Y���C����ln�[�f�=s��3i-yO�R���e�;*l�?��=��_�L�Vgzxצ{�ͭ�%����t���3Z���M/L��&��
�l�U�\^�Fzx�ٓ�k�Ϣ��R�s��oc�|gް�b-�޶�O%imH�t@uG����O��t����;eߚr���TĮ����7�^��w�"
�R�"�+�Q���gg�Ř��焩�.����\%p�2�sb����n�i�p��������ެ�Ѽw���v$�E�٠���i(��"��>�;m�X<TN8�A�U��wcA0�d��0ѻ�Z_�e����>I�@���Ŀ/˵w<��#r���Y��j�zC��vfm����0ro�CT��ڶ�k��{I�K��4=��u�G�'�lѹ^�[�r^���<�����+���6O�U�Y^��)��0����5l$��������e�=���6uB��}j����U�Q� �ܲ���L����7~�o�"y�c����5ތ�E�2�]#�Qo�*�y�;]�(�}�F8	���{6�}��
{���(0�!���F�(����U�=���x]jGε��V���]��=���sխj
-z�Y�-��X1��A�#t�����^OH�c=�Mvھ�P�;�x��l/L(-j�z쪟x'��k�CN�є,n�ճ~;��wx�l�c�̺j���Þs�lK<�oǝwv��vq恷��u�;B��M� ǰbPSzj���.�Y�ੴ�A�}ᶥ���ٛ�~�I�!=E˲'0�%a�ڍ�>p[mL�)��fUϽ)P�s������|���D��GjI�]Lc��|����{�\F���� T�h{�T�q�5���?^��A�E)����ﾈ��V��4gM���F�Z:x��s�{8�x?x/u�����Yx7�y�c�\6;UX�Yo~���j���ҞʭZ����=ީ���{#�=g�zw�4���/��&a��KhzR\�Ë~��֮�G|��̝Jp�`׋�c����ϦGń�]�^+�V��s�z�nr�T=�W;뛨��n�x�js��eb��^SW�ͨƽ;ucv�����Ђg�^�%d�c��5X|���.&�&��~s�
��Mzv��ۄ�����h�0�u���N�bO���ңUB��q���c��~P�?\z��P_!x�:����f�kN9�ү���D���ɘ���<�c���z@Ìg��&��6n�H�UZ#�����tO��Ru;V�j
[��Գ(���d�\��s������蝭ɾ�U~#��Nυ1��V[��o�E��s>Ki��fL���t)�P��bgR��Ԡ��GrřB�{�,�:2&
:��W������b��Cv�0�X��2zKu�jo6�jw.�.Q�\(�*���.��E%��(��]ha�z���9��g��G�%��$���̏����T#���S}��y���Ke�8��zDc��	Ƕϳ��a���eߕ��h�ӏb�I�;�ШM�Qt�|�\�i~B�c�Z���y�w]J���&��h^���oCP�p��B�s:�KTjWU��UH�p.�nMD��_F,�y�IT�,LM&�=8���h�;�ў�=ag�l��C�Uk/!��M����Kk9{7��<�_T��{���8�.(34q:�+�q@ܳn=��_u�b7j���_�����S��V����Ҹo���Sɨ�ߪq^�@^�죗��h��x�����e�F�(�s�5��PО�Pٝq@{=<~��H����V��9~�j�a�+Ny�y>a9�|1����5�]����(��$�q7�g����#OX�r(�k�S�o���
=�Z��;����Ϲs���m�l�YT�A�=�����Z���9���<w�Y�8���z�{��{I|��BU�w
����Y+3wb8;��v�ǡn�EX�u u`w�h_Y�Q�*WpZ��L�Qc�t�Xi����]�����Te���s��9�n��������B�>5;ՠ9/d:������j�\Z��izR�1>�y�"�)��s�>^�����]��Ҟ����t��K���,����v�{1��j��[=�r}�	k^������ۿ����!��$5�U�Oq���8G�E��]���}��5�nDy�zދ���q�-}�>�(ݘ��X-�o\���<w.���	{������V�ʉt�d�B���R|3��Z�w;q��z�QM蘗���?@^���U�V���<�I��.�y�D���&�j�lWG�E�0٩^̰��x*KYM�j��ڧش��a�*2[��)�=Z������5G���/m��Vg�wL���?
�~�3���	o>~{����S�5��{Y<}���=#�G��,�X�1�kqQ{H{$�Y~�N3Υ�;ہ��9OFD����_�R�1��$�.���W�ژ�*ە|g����N�5{x2SG+>�e�����"�@�O	��Yh���	�c�wK�7�<��_d�GU���d�Q3�"�}����N���>�'� �5v�@�W�鞹��^{қ|g�D{�,e��;�>5����N��K��W+��y��{;������{���V�Ϧ4���Ht6�>�k�����֯{+V�539Y���^��f����X��+�j�,l���l��.�r7�����/O�d����^򓶦DM����u����z�K=�d�k�n{��^��:�:��==F���D���Ӎya�d���*ƽ;U���������T)Hzz<�TS�z�w!�E���fͯQ��m�s��/�^�V��^�����cgٻm��L�'�No�\���Z�Ez��{���8�[C���[��c�^�M�-3NKڒ�Z��E'��c���-��n�����c}�F�N�g��ޟFĺ��������JʏSsE-�T�;�-��y�Ccq]c�����wg՘��7�b=P����l/N缬���~j%���-$73�<ZcT���F����М��q���e�G���&�����x���{�U�#�s����{z;��-U�(���-�3���IW�ګ�V���ɶ����<Y������gt����"J����ū�������+/2�s�<�h�����K���_���x-���|��Z�k�Xho�:]��Cڶ�w��̋�>;��)�l���y���������D)�5�-c����m����2X��hM�{.oKs��ZmmMF��aŽ�,���D���l�l������h�f?1ݻ7w��f;���p���X��n1���TCё:��c��l�/
�/�\�}d��%���_,�<\�����>��
й�[5��Έ�善�U}�zR^u��k9ZS��<�;Y�=����r�w[Y3����S�����no�.��;b�z&�����+�Dש��.m�l��o3%C�%�&q?�?j�X��*��N!����j�]Ģ;M���^*��{n��h��g�轥�^�T��!�rmP�X}���yї�<�"�G�}��Վ���C=

'�ě��m��Z�e^�kӷ�h!���w[�y�+2N5�Yga"���.k[VR��/Y�.�*r7S����{���bOa��q��ǎ�R���W�Niz���Wc��Fh~#.��v�:��-*��/�I�{��f��w@炻����4�K*l�E.�P'�+�ok����<�Ӟ�ފ�����ƭú�[����6��x1?9Z�p�w�C�Yu9�+^�-H�4S�� ���Z�JU%�rou��8k��\�ݽ�7K^�k��7��5?U�˥��衺'�ҩ:��s�[�~�ՙ��s����(2�OM�vw{�{ו�+�����%��n /zi��޲|��9 ֯	�xߋ�]����g�o��G�oݪ�a�[
����Gu��ba���[��cs��i(�p�D6�*�iL�����~m��2⵼�;5/mMD��_F5�м����z���q-�	D�ܺ�ՍPed�#v�yH:�P�syW�{y_fb����t=W9Nd�ۅ"	3�(/�-^mՋ��ԫ��O5�o�������7|�+�._�[�4���]��Z�{�mzY��s"���b�y�`��o���Vs������ܼ�w�HԬ�,cv�^&�&0ըv���Z��֭<r���ȝ�WB��<s���t�h؛P����j8�::.�v��Ù�Z�Q�hNB�=��|�L��Y���!v4(�������7We��9�K�����+0E<Ǫ�?�/ݶxxg��z�t���A�kX�H<n��52��Uj��.m�[8�F�C�ɷ��9�zV�A�:�@�N�;'Z���ҏh��F����7̧���ϰ`���&�c�@���ae�:p���/�;� V�R���8mҐ�����z8�ꂋ�-�Gf��q�t�"�8g記����=�4��ؼRCUɖ�,%��`��+�#9��Q���gL�8�z�۝�`��o�Tu�Cҡ-�v���X#C�����x5������G=��ҷ�{{�^�E���\(��v}���V�MFPp�/�-���Ut�k۬!�
b�̨��2��9[�c"Ǳ��B�R7����܌�줩/����3Ӌ	A�W��Gu���8Z�ͭI�c�8���x�(�n�g���`�.��uuꂘy�)W}c�o���4��p�158Jm�� ��'^�H��cA����T���R�k�di�l�յu ��$%j�B�h�VxHe\�g��R8d�mKWj�n�R<���SY*��bL�3>�o�\�Q�E��^�]yW=�0����dݣ�:5�c}�o1��L�۾�mԙ�c��R�Zm�M�"m嗿c�0.����x#����lI�n���Z�v��XA빤%��<Hv�vc��J�R��u��}��5��[}��H�G��^�$$#�>�sӻ�M�9!��Md���kUl�ႏH��W �/�ȳ�����<Ɔ���X�㱜z�e������),W�.�A����fU�42M��oga�j+с�A�jG
��<�;C�'�m�eŚ������4 �F�N�� #��Y�]\ʊ��z�唛��i]����sg��Yڍ묍w�v�y�Q�<3�϶�&���/��7�9��SPz�F�<�5���Z�A\�w5J퇟�*i�j��N�����}�ڬpi��6�4>�1��Xժ��`�Д�0�>�WI8>�˕cnKx_�[>��|m�R��
ӨG̯a �״)[�QWE�7�'��o{Z[u>}]r�o�%o��,��u{T��*���o �ރ�uN��K��Hhd��Y��W%y
U�TO1����o��ni�*�X�QͷNE�-��l6��{{0r����X9�^:�rv�r7E������<եV��
ƺ	��3 F�3n��7�`>ڛd�[�Y�۳�v[�v�$�s�&�l�F�A���)���3m���(:7:֑����]�	�6�����J����bu����/H�>��k<��V��N��;�q����e�lVfV�y��������������ZM�L�I���\�AX��16��%�k����ґ#IQ��s1�F��#l�"�4X���1�L�2�
LF�L�Q�12�+�cj5�b4�d��L�cbň�	r�n��F#p��w\�4d���;��E'8����фܸ�*K��5�G5�Nv�Lm'+��Hg(�t�Fܫ�S������������&��w�Wu�������6��Ŝ�#�Ȝ���½���e`j,�8�֙�T�
��j����-�ͻo����^h�T�sfw�إ�ߜk�Y��3�i��+�Uiv��G���X/�q?q��y|w��y[�ޞ>��z4�N^,�Q�&��<��S�[��D�6�^�u닅/�'���6�ƽ:#�
����l�2o���+�@�?�N�D�{X\m}�G�&�;o\�d�*G��"^�������c�KY�J<�[.��<�K��%F�^����ŨI�����7,����z?0;|��#���q�W�(�o4w_ԗ��t\���}8*����3Y�����l%o/&�lB�n=Ev�r����l���¸���k;�śFz�F����5�[���cr��=c�U�N���������ч�/٧+�Z}�7Fy���!����y�>�����y�W�2� ac��xm� ����Y�bC�w�^���U�P�͠�n��t���l�t����Α�&���9��8����r4z�#u.ۻj���T�4��[rL�N���"%��yk��ن�vJ��q��Oi��)qN����q�^��:�1��C;���'>�L�o�>��gby����"7�����a����{R�?FL�����x�of�W�!?nx*KY�M��i�Rْ��O��ڟ]��9���d��8>O�@�X{<�/m�U}j�<8$�D��S�����l��u�m�=��'���x�!���gD�Vw�i��p�u{^�����Ono/W�}�U��{-�E��P���B�_S&�zIr���:a��VG��z����9���G�����{�.�=B��S6���^z��|�h��ʛ���eR�gڵ���y��3��y�u�ۼ�T|���H�a����`̨*�bț���6����z�
�p���vX�[ϻ�o���O�oˉ��ZW�l9��[�gW���Huy�� +}I/f��y~�J����~���!�7h��ʤ�*��[3bo���z���Õ~���^�ܦߓ�~��SY/~�w/Үu^\�H�����]qjqn��[Ee3;�P0�������	Aϳ��w��mNgb�h���p��u��O#�-.��m�����w'��i�V����V>}гF��vX0�p�8>"�Y�m������y� fE�-Q���p���{�b�
|+勀bےN�_a�Ċ��`	��s�i�x����F��Wc�w�|zoA�y�hn�"dP�j�����i�K�p�d�I��A�^8^���*�����1���-N`M�4�բ�
��٢�nbr�n�3ު�>�Wz���:]c���~�h����&o};:}醯�M������1��w5���/�����{�v�ߓ�?���
�7ڏg�W��W�]y����fݭtoV_�c���7���VħNQ.s�!lzn
�F��Yp��뗎����(�(�z��r���76wz�|=K��W�yFx�6���Q���{ؚ����+7/��ɯ�d�;��M,p桷�`����m�Lݝ��=R�V��^Ƕ�܉mg/3O�|��s��?W�h�x9���	ɻ�����T~��ޕs*�M��Y������Z��+��-��b�%�� ��r�o�9٫)a)�2uV%��6�á��V��XZ07�=n�N� N�\�I]��2o����èҺ�]k�h옡���>��e���ǹ/[��12��8wG;�VK��	u�������!��vV:���Y��D��ˌ�������v����g�@��.�	��'���m{̛W=����%����7�z�c�g�{\���yZW�j�;p��i9��^T+̷>N/"��f��-V�؅-�sY���k�kӷV7B�N[�z�{;j|U:Q��-s�U.�+l(�ě�v�s�4���5��+Q�l[��6gm��p��A�@J�������J�[��p�\colj�q;Z�dfo�JK��b��5��]�*���h'�B�RR!�TN��g���>�6�zx��=�?&��&���zb�#M������>�tCK"N�j�J^�(�bō�R��]]B'$=���I�leD�Jò�}�Lx�����j�U��"ol�f^)�����oU�Ҹ������b֥����}���<�"��FA�	��Ҫ�n_Ӊ�-�ѹ�54��@v�n���5
e���eL��8~��S|%���ʽy�&���kɃ������v\Jv��d�=V�xEr� >�tx�j���L���C�K㸩��ޅ)K�hZMG}��G��V�¶����E�֫y�g`*މ�̽�����еS}2��{V�v��v�u&�4d�;E��Ք�6�9��I�o�*���)���q_T{�G��f?$3��~9�%܎���~��,�����ۛU˽y�q���/Ƣ�f�:�67�Z��{�<�o�"C����g���J�r��F���K'�Q�4%rf}���u}�o�!n�=CP��w�K�o�X���{R:}�xg�ܶ��}�QK5�E������!��ioÁ0p�q�G�;=wk0���sX�^���my�̬;�ƽ3�*�ix�*�ZZ��S����:�b�TM�T�X����Pu닅/]�!�Rz�y���I��=��Z81S�Cm�U��(�P��aq��D�Rns�zW��;O*xvl�OP�/9�kԢU��n+@و+`y��*5T|�U�Mr�����w
x��#�v�k�?{{��8���y��s(?�8\��=9d����K�]���nMWX��l�Ţ�V2��^i ����鵚�Y̥�;�͓<5�ʶs(t�%�ǈ�!~X;�k�O[\t�]��GZ[ټ{pp��7���gi��l�묷>�|vy�Y�{���q��@+2ۋ�l�'�(.h���ҁ�����N3���r9x���ߒ��e�8^�����۸��*���ϷG��O7��<������'�s]��ɢ��vױ��z2�����_J8"z�m�;j�g鶙��(�S@F:���9��ž�}��![�hN�5D�9H�w�x7�v�߅}nD~�_,k��7<ji\@w��݇�L��J�P��n߫�<���=�����;[#��G�=��w�	�nx*���9����y�U���JX�p2�w�7ݱP��=#��c���b�&�N|[�oϊ��UO�5�k���LKn1�q?=���g��f�"p�;��_�e62<]�?v^ɓ��&����n��s�FD�qs-s�w: ��d�K�����Ч����ې�VP~�u�=(
Յ���� r�`�Q:��ؔ�^����V(��I����٫_����;���=�6H�}���E�0Tړ^J���6�H�G�WN9��"�m�B�U����@��]�� -x:��J����^�g�%z*R�}뜻�1K\�(�upw���Uv��;L�e"Aкu�-�ط����2�jr�M��+�燺MlJ�!���j"��"�e��B��.�Nr��qϯ�n[�O\]K����z�Pۆ��Y�����柡��;�-�y�����k빺��у����h������v��v�#rm��^ע��c�1ku�x�{��=P9Α��g��'7y�+]�o�{"m���\aq7�76�{p�}��Mu��^���&��ԟv���O*_��73NO���Z��#Ż�ݺ����3C����;���z��NPSd�At�Y���j�M|Ry4���s��k���<��sN�n�H�U�*�����J&J�J��75-ۀ��	t�X�aw���7S������	�����N�N��j�za�yQ7�x������2'5b*3��1���0Rlc�s�Q�v����S�vzР�+l�Y.�-;�];gVz��ֵ�h;A\q0�9�|���;Xǹ�����#�H�b~c�'������e�$WGw7:�u°:��^|+�z�U]t��F�~�Z'N�e�)`�J��_7���q������(��h�]*䰹h��u8��	�)��F�ӣX�{���}��LqK\�N���D;��]���o�tj�SR�MF7����[S�0�2��Cbb�ۗ�d�\N��WM�쒪v\�9����b��<w	*�������WJ���s�c�v��y��ދ4+�>_Bm�����N^��ժ�s��?W��yV;W�|4C4L���8�y���0�}�d[ځ��鷕�ef��Z��><��a��9�Lٚ��ͨ����r^����ٺ�v�zD]⚛B}�]mF�N����j��מ+�3�x���6W?/i��Z[C�U�u?yx�s�,�V:�/�3G1ϡ����Fl�q,�������:nN~~��fy+9�c|�5�4��� �:|T/n{�G��I��m�:�~*����)��崩ԕ>5:������K��Tj��J�Ż����н���q>?DCZS{���[Mc�5�֕��P��UIH��Q;�����Y[�!襗mn^�����#�5&��W��GT�\�p�=�\�����DT9�5��	�G��F��0v�=���0��Mk��T�	�}��~C�v�<�۪�cۃ��³m�}Ad���\^�PK#�aeҪ�zl��`꽗7�'�mJ�٢o�e�smǨ�/�LA�`4�N�.Ç;�u���8�^~+�7���Gܽ�U?Rz[R�+˥���ǌ�=��u$T����ġ3W,yN��-���S��E�2�S�IY�-���e{��U-�RZ&&�z��f7<DjiCzШm�Qv�ǹR�\a�z�uD��+PP]]l�#=B�~rW�r19�hU�%�jz߽K�u�S�u6g�և���}�U��6f�A~����k;�ߗ����h��uU�IA-oϞ��]OǄ�Cё���@���y;�Q+�,q��U�7:��T��kgg�S�u���9����x�dn��W2�JK�Vy(qV��T��	��G�gL�nK�R�՛��y�׌���9nh��8�^���^C#FyVz<sl{l�V>�U��.�X|���T�OL�ڥ�	���vpe_���ǁ��jЮ�[��7b���5��}��T��W���cX:ڋ'l��p9�a�|��Qˬ�D��R	���<<r-u�0��W�T�7n��ܧ"���x:��ݭ�[��:��%����rgx�d{z�Z�ݞ�q�^��|�
�G�P���ϼ7*��M�w==R�<�w�t��4I����}m��/�)��'�b�����_��k�;R��U!�����ǯ��Ԧ�C����km��/S�6~�yv���!��s>2�>߰z�ι绶��@W���̡ReH�b���ɶ��:O�U�/o�]h?P�����}��`�<��`{�P��*k5��}��O֦ۿ�����r��0�O]^��ʽ
�t�@������W
�M�\kƷ<�=V�e7M�|=ełr�_�b���ڋm"�	u�.����[6�_��[���j~��V�  4������̵{��0�q�%"<`%cV�7<ji_�ߛ�k��k��_e��˦u�|��v��w�?�sH�}쨝�~������&h�>�������A0톅F7lWЦ�֐�����y:^�^�/o��c7@�
��D7��5�/����d�{�d�KG�+����*vmc]h�1m��B��zm�kB�L���ה+�S�7tl�qe`�����m��q�VC07�V>�Φ��F���Њ�D�0�Y��FIJ�&.���ږxyӿe
!k�)ѫk���n0%ë�岑���6nb�|���w�p��Z��oi�}�|yF�_X����#�X���=�x-՟<�?IV����n�:���!�U������Z:�{�{,�q�Q����Զ"Iנ��b/Ү�������'�1�iF�:�����vv�2����)��H�*;�P���:���q�;6y��z����ȡ�W3TUh��}�@7M�ԁJ�3q��F��A%���.��;q}h�yr���{����7[�9bG,'����w)Ƨ�X\�������O�������\�Lf垹�t�G�o�w6�O	^�#�]p��.��u�ٲ�n�^��v�5 E�j�F�Ԯ\GRkH��Qj� �����u���jWw�6�Ee㱝b���о@jB���5#�I�X�x�e�p�$�R�p�Qr߰5�*"s<z��J0������D}��Z�+b�l���c+)L�`<^�;�D4%��ʰi���-�ל�C&f%�� Ѱ��cty!�h>�7����u��A�p���R�U�Go��]Y+([��㰹˪�uD��H��a��蝜�#zN־�qt�#��4�m��G'U�{���֗m`� &���T�̋A�o�Z2Ǻ���p��M\U뮞����~(��ˇ5h�*�⛒�9�u�.Zye�R��`w�m�2R�ti^Z���"������`<��Sa�X�Zx�S�z�ɰ��gUN���v��7G�ǚ�<D����0�o5��Ďmp�]��k�;0���͝��U�]ҙqs�(�}(��N���	G�;q{k�&��鸜�(8�7��
oB����˻b�'��<O�;�-oV28~'���ʽ���y�,�yj.T\_Ay�yt,�v�B�_P)}ƥ���Τ��Zrp��.뙳����5c�T�Vi~i������ݧ4�'��m{FH��P��1��$�G��
��m���o�����1A!>��gr��͡r릝1φp��s�!�Z��Os�뵓�9Y��^�l��/u>�9��X�	�"%�5C&.,C��f*��Ջ�CK ᕘx�ta�hs�vb[�&����Z�0�r�u�{L����k쳽�j��[$p	+��qbT�a��T��a;}u��i;y����+>��,�t�㞾�|�a�Y�q�x����pAMt��_&-�׻N�-d�!����y��������|���8|�Q{Q�x�|� ��ӯyOJ��m|�1l��y�,V��]���KI�ɶ�j�Z��s
r]?&�vw� -͙��G�M>F�\q�:i�ZY��>yӹ��`��cF�Gw��w];��:��vlV*- �F�ƍaѹI���ӻ�.%Μ�諛�DlR]ݮ����.�ww.&,`��F9r�m2]���R%r�m���u&��)�s;�;���5�n�ܹA-�W#N:�\�Z#��b�ċ�j(5'-�wnkswq�gu�\�F����Esk�6f�����s�wm͜�QIW5%�b�N��.s���)���ur�5� �������;��MM���Ŏ����Y�ݕ�k��49^��!�h��qŘ
쭏�)�m�$�sOd��z�~�M�ɉmF'�WED�;b����?^�ǉS^)UmU?�nMFno��n��X���!���k}$=�5�)�^ȷOJ�Ӏ�����Ks�̾YZ�����<�^����{��9��7n�O!�����6'�N�e��V�����e|��Z�񙜬����������}�ζc�s�z���^��-�s����-�'�m.��ג�'��ɅP� 鼚+#]�J�*��w���sW��j�Z[C�U�7=�uzJ�OV�n�1��O�w���i��=YK�\\)K�^g�ōd��Xݯ��R�$�N��{�Zۭ'�K�;�V���ɷ�u��W��k��"����Eϡʙ{pm��t�k���:.�ޒ�7��f����Փ>�����F�T��q~�A��W�R�;�լ�����{,���h1��g`���)K;6�<b �&f��K��3tZ�lA�B�7���>�}p7q[��� �H^�EBA9N[`� �̺pL8���(%ն�6k��q�nNl�ad	۔pcu՗s���ק2;k�q�6�ʽO��H؏\��舘p�!W��R}�	D��D�������[�R�-R8<���o"\�t���޵�V{xw���ڧ�!(�Of���Z����˝��ܟc��g[p��1v&ǩ�9�S'��_M�鋞�_������4a��������u��j��v������(b��C�6�4��_���7w×e}�N7��B[SZ��e�;��'��
u�a�ZH�T1�U�����~:�.%���Y;��%SK9��q�r%b���P��CS#���G�V}�ؕ�tw��|��ej�Ʃ�k�������Ϣ��c�*�=����{�5��:��3}6����ӡ4���ی�콛��hs;u����v_��7�f��"�|?JK���ͪ����ز�^s���R�w�32z������H��|�V3�����z�hڵؑ�������)b{x�Kh�>R���F�nV�gm����q�S{BޟzK`���8&��{z�03���)�[#k�V�+�T�>^�l^.���S�m��{6��8k�L
*��M4��n�J�w5,в)��➴E/�A�e�Ǐ#�~��^���Ŕ�܇W���k��i�=�^�I���73iyD~���r�IBڌ2��£q&��Z�ֿQ�^���T�>ǵ�q����y(�˹��\�X^�ңU/JW-�8n��͘�ʸ�Yx:��7��;����Ì�V���w$�z�H��B�?[��]X)��.�<��hx7]э[�u��n��?��d�C����k>�^�������O��:�.5c[��m��t�:/��B=~�Jwn!֨��ǃeT�W��G�^�:Ұ����
l[��9D��=_H��7Ui����*���d=sr���-��Z���v�Q��XRJ؊�^�yǪwU��g�D�:�;~uY��t�-:����Ϻ{6�ޗ�t������3��p�:��ٝS=B�,�����=#����{�_˖7���+�g��3�2��^�ܿ;�
ݦ�z�N\����,k�1y����D�ںv�KoJ��`�]@���u��Ջ�(��Pǯ%�h���w�F{&�]��>���b�pۘH�Ȑ��}���绷B�M��O��1�i�΅;{��c��
::�N�L�{���͸�@��q�k�*%��ȕ�^h0S���NR�H���߲k������͵<��=j�������Cʛ�f��-xӴ�Zf�eĿ��󘬫w��^q�g-�Օ~p3<jt`~�����{���|����R���m�u~�U�Ϗ�39\�?w����}�����u�+S#`��O���{�v9���Ee1���Z(��
^-��.� ���S��k�����K'v�nTr��������^���}�<�튧�͒�e�"�v-q���>��ܲO�]��l>���:�+þͩ۳��K���9a��Lz��I�&��:O�U�/o�N����!�b��}ũ��k,J���=4{�y7Z�p�I��Sm���K@^�Mo�|+1Х��"�bY����Z�	;��}�&},���o5f��]��*�˵,(zI�<G"�+[�p�Kb6gx�I[���Bp>�{���f�Hܹ}�C�4M9���l^r����c�rWd�|[G�D5q+��K�K<h������FԽz&��J$�U̝���B̓I��z��<���N	�~5�w�T���/������*���W��C�N��R���d�G"JVU��p��ܿz�9��[�]/�����,j����N�v��ة�~WhR�d{�I����/F]�<���S%V�[Q=	�����u���>�ΚQ�,��G�[z��h�Kv�B�s�-��A^sK��
]��=��>\�{�g��YM��G�mM}�15ۏ8UD��;b��h�Z��)>�;�?nng�5|q�,���W��V8s�6�{Y�z2&ho��������=��V=Vc��Ȑ���է��g��~�a�pNf^���3�6;�3�G��J��zm���:�V����Z���W����/��@�r���E��Qw�<�?4_y,P�(q���ÈO\k��oD��{^g������<�/yHjy�^+%9a����b�Ūmr�V�])O3��1ٝ��t-�]�)�X����d�V�L��v'V���9r>y�kk4���OJPa��e��2�w�lW\X]YmU��Բ,��&t��8PF��la���q��\����0_ff�鸳�6������.��]x1[eө*�]/!��:z�gs5�����{�C���r�ݫ�*Uǝ��YOC8U�:�\=���𨘽A�����ֿ\z��wp��5����5�3���J�Kډ��QKcŻ�z7n���nk��y��%��i��zi�+�V1�]D-�E���$�J�ǻ��~����A8�jY��I��9\�[�eBT�z���P�T�`4�J�Kr~ƂcofW���~�Jn��Z�t�E+MV�T��>فφHt��;U9��*�.߳�aM8�ĕ�҇^i��������ܑ�����`��eW#��g]VMK������s�V�j�7��v��Q��9�2�۶$#y�-z7-�W����ޥ|l҆��	�*�W�Zö\c���� �݋Ʀ�ֵeԬ������rR�������T~^�������Ŵ�x
�=����d���������R��.�V��{q��>�)tt�[d2���v@K�0��a9OGf�[+����%�.��q�]��Ь�h��o D��~�s����Z�z�M�gP���Ua���z;�2R�x��O�/��Z��=�ͳ����|�-�JU;lE{�m��%�g/3��7��Oh�չ%|�W&e��|�M�G=�s�ha�������ŵ��r��]�W���]-2y��ڢ�U���S�+E]�ϱ�.�v;���Rwu�)8��\�?i�>�Z����>�g�2u�<�������8������Z��N�Գ�%[���:Q[�����joh��z�&ߓ��7z�_����.K9;��SB�>5:��u�s �T�ڈ�k�2��
���I�t���*�x�J�fsY����f{k��L�q�:U�8=7:�sҘ�����z�c���q����-q�ն�?\z� {
���h�T��ʰzt����6�?3;��!^ ��3wh�qн�o���nЇGϽ�X?\�h���Ǐo��Y�į������Kr�c[�q��leD�J�;-}�N��O3��S�%�:'$̤�me-�zk8��4Dᾮǅ�[X]j .&��B��叩�g.ﺖu��r�3=�u�\r��Q��
�ԐV�Չ偼Z;��n�l��5��z�)�X�xz:Sv�������s��]��ztLpaEq(�|���]f����~�{g����6�:Ś��n-j[>�R6��Е��ITF��1R/~�������MD�<��s�{SJ��p���5�i�5��[��C�rry��KS2d�����|���Ļ��r��{-;����xc2�%,Y�8��1�q-׃���u�{]h�Z=����Ǆ���7\��g�ܪ�zu�f������Mǝ������V�yt����O:��c�؃��9�:h�9y8��|��6�k�{ǣg���T=j��l���HSK��P7rfl6�]�4o\�eJ��׫*���x�=����^̍�G�ӄz�¹�y����?|9�ZLo<�.��\��}�N����=!�5�V�]�ì��ȋe�=�z�K����8�_N�8�;�R�3�螞�갯�͆�����y'w�)'�>�V���O�߫=�j���z����R{HА�9�m��ݼ�w�^u�C�#@Z���;��̂�"]��K���1t�.`���1ð�5)J.�،c��b|���9\�����R�0���sO�t.���W�f��)ڴ���Lβ������5Y1%�;��q4�>��^W�Oy��v�ۭ����_c^���f
ـ|��JCj�⏰?o�{�*���Bǫ(�wx���������Mgc�|=���,�7��J�"��'�J��W*q7{p�c��	��6ݏY^mD��Ж��1&�<�������!h��ꯢN�T�BN�kƷ�/6ތ����'#�.�A�R�}��"�V�{��{�}Ֆ�W6c�)n����1�J���*H�vۇ�w�uHz�[��S%����G�J'౫�1�޷R�gq�؇��2�k�w�8�����&�(�f��U!m�ޙ��+]�;�W�ׯ�o�HrP�:���^������a�錅4槲�Ɗ��՟���$�R��˥}�'�yP��֤��Cn<�+��訟�߲1�����;�bS�{5ͭ�P��sԖOѾ�W���c�4ہ�s���Xً��!s>�wW}��WEH�s���Z�bK��b����s�z��I^���-����Ay}�=���kz��5����s�!���*�ʶ�.Tz���hR'��`6y�'��Va�U/�A}�Q�xAm);8_ �6�۱���%��s�su	u�]�ܨy��u�*�U��/<����_,�Zxә�~���g��Jf��hp��1c����1��/�k>��Is������j�˫(���}gȽ���ڊ�ߧL�3^mmWz�\�l�C�����N� ��^�q��&�q���?vytU�)�md�n��_��@�gg
G��k���2sB��8�£���������n���PU����z�Q{�)����qV�b����Dޠܦߓ�~�*��F��18�|�-�TT��U��,�'��F��b�e#2x'���0�Ou�Ͼ|'������{�5\��NQv�]/g`�=;������l�K������ʡ��e�qS(.8����n�Ĵ��\j���Zͯ+�YŹ|��zn1�#��wðl�p� ���Xn�GϢ����hP��׏u����x���j�<vo�x��0Ϩ���i�阞>a� l��G�W%��gv���Ε�W�8�X�N�予�y:�cŕx�u�o#o�V[f�:Y��MᏵ;���J��V%���'��s=�,�[Z��fY�`��ky3��1����<1�K���q a�p�[����=V��C�)Ad���Ͷ5ѾdW�#�Ipv�{{�1މ<�c������
ܩ\g�v>˿.�&i�U�Zp�8f3� ��0s��K�����s:�%���X�Sn��ܢ��N��n��N�<�X�1�s�n��r�1F@��6��A�72�\��s9�'����dGP��qkOgsi�mo��=eiݩ/p�� �+GT����0����cv�)��s���yI���B�:{8�:Mf�u�ͷb��Z��.�o���Ej�~��n�Pj�^�.�^��$n�h�ԘF�G�u�#/��l��I��x�W\����m�&��rθ�)��h���9!ǃ5���"�=,���{hc�%D�p]ʗn�m�O�z��:Q���&/l+��I��+� ㇍�}׫�h[giI�+�;k�<�Gy�chTH�u7]�ð�u�N���.�w	;hH�p#�S5�}�m�ˁ���[��Ͳ�rli:�)�;W�[X'l ��w˻"S�A��c3P}K���y�z����%�tN\?dz�g:|8:��x�u��N��F�/�*����F����ܛ��Ɣ�^�/��+�h/.�7\R��/���
ⳅ���9���&/��BȠ�^S�Rh�C�H����Ɣ���q]�ۭU�K�eA�LL�ds���6��P��c�����6:��f[G�QzZبhs9'2�։��r��n��|��Z�0T��Q�(�Cy�c��έw���5KA���l��b7}��M����V����n(ʣ�6��Y�)�ak;�;��mV�e�Ď\������6���{���Z}v۰���=@�̵�M�s��qTtyo�㠕����gQ�V��N�&oW��o^�[�G7/�b
��>cC��e���z����{6
�P�FBދ��v0+��^�p=<��7�5��nꯧ��"q���=PU�{ނDV��9T�ɵE�.�I���G��}.���U*ﳯ�[��hc�����ؕ �t����cG=�����a�n&��uڏ=�h~CMyw������n�����d�ն^=;����O\|�j��w�fn�T�=H^gYYhq��a��s�W�z�>ԩ�b�=��/��W].u�wL@r��!=g�Bz���S�tq�Y+�gX�v�R�+*
�?�����?j yѶ?j֔P7��'?'˳R��h�5���bu�K�Z�v&�Da½¥�o�5���ڣ��4�=��/��
��ڳ��~�3������vy�Z��8��NB�Ngavp�t���b(��E�2���2��p�)�SR7da��w7����M٘��6�ƻ]��&.�|��B���"��4>ܺ\���5��w\��k�I��ܹQr�n�4k�]9F��(ѹ��ܹ���7:N�;���r�M˚*+�+�wn].j��Pm��27��gw��%�����Fwsu&��cr.�\�W#t�K��ۜ����i2wQ�[�͊Nsr�h���E���w9�����2�k����r�ۆ���#9�71")��rs�"���lb�b��'6��떹]4V64p��4m�����Nn�4k��\�X���N�nEc�M�s`����Ꙝ �ޕ�l�Q���mfo9�X�S�u1�.$�1�`�Ha�O�̋ut�{��jܟ����y596��I\�yc���߆�/��~��#�˴�L�M���uUqQCRS��U$4��Ea+�c�_=�W|[�]/����^�!���=���ӌ�1p<���w}T�|��W�������G�d��D��S�\�|��_9���!�m]и��q=��ܟ�+ީ��{V�-ftX��ۥGЌ�ȏ)��f��-9gZ�ѻ��w�C��f�5=y�|2����W�:��`i�fT:��B���T����g��h�=�C��k^չp{ӣsM�ř����Nv��n3����롷�s��ސ
1G��\m+][�"^NU)������zU�Y�*+��Gg�׷	I���E./�z%�~�3]�_�����Bg�aE�Xb��G�:e��`ީ�:%N{�K~��Xر�f؍�ON}�+�c�XȠ��/������T�|�v�7��\�N;�).�k�������N�"�r�N��}J����� �ވYĜ�w��{�\l
6Nd�l�K��Al�j�j��.�^r���{*ww�v�/΍����
Jnvy�\x����z.8��:�}T@�sћ����}`ۑ��$zhN{ǲ�ɗt9����N�:�Χ����i��E0�b���_K��S3� 	xɾ+��V�س�s=G1:�Q�Q�,��m�fn�R�6J�ذ� QSSo�������o���.!�۠��Q���j�� �2ˈ{T���u���vpz���xf�-=�q�g��NG[��/-�g�]�9@���,r�w2��ϭp�.�7{�.��]���3�e�ҩ�W3~�;�a�v������6pK6������&��LJ�[䴞��D��.*e�M���©ݬ�3_V�c�0ϫ��]�ZF�֧��Ļ���T�I7��83}���G g��02 E55�%�2'���o��V�7��ǋ�'����mzg�Ng1S�й�R�D܂��N������a�^�!���r�zpWo��yJg_��^U|�4���x��K���_#$�n	g����������s�6bi��>���%*�^���r��*�{W =���U���櫹#��:�/k��5���vbH��K���{�[٬�v3�����ڤk\�E�H�&E��G�R�����qf��dF�Yh��UL�>۽��\�Q�<�9e�������#7�#B�tA�Gu����6w�%}��w#>�-`emj$-K2rڽ��^���c^}��@Ү�[�u��y�mݳ����C�KkE�]J�_���51j�C���喬�z@��"�wfpy���4��b|���t2&9q�QoM�J��+��9m�-,�����6���W�/�Ӎ���5��l�w��Uq��j�܇�#z\{����{�+M�b/���M�Q��Q��-����[�dn(����Z��l�.�[��[�Ķ��5r�b��f˳׹+�kֳ���%^촢��d�@f;$k
�fcx��؈_bjȼ�TEP�%<���h�F���r���{���k#,g:ȧڼ�]M���&^vadEuR2F�%Q��@��U�{���]u�Y��{�q����r���w>��b���h��jI(�|&t3#{F�L�Q��3W���X�פp��of��������=GOqY��;s����ei�+$��Y�3�j��Cނ�������K�.�y9ϞMW}�<3z:��{�3���n|泌vĴ��v������MS���=�z�΁ �H��$��^<�r�_�.�s+zF{���G�5��b�`�*���g�׷>�<o�d@N�3~-�eqU�	����]�r��1�Po�e�z�ק�1O���-�/��CI������퉷�S�l�9�M�[�e���0��ѳe�����!-��P���#�䆝��۾��^�[���''ou<�Z|�ER��o^u���]<��lC�J��<*���>�iw]"�)B�_I������<�3����l�a��~렅Ǐ���v�Ʋv�LZ⸫���{-��9���O.]G��Wq��~=��{��o�}��.z���Ϊ�����~$���B�="�n\v:����e��/��/h��m_I|yŞ��{!�������5R�k�1�Q�&f�N�l������<�.Q�N�Ң|v�aβ�����۹T����E���,!؍�^��Sf`�X��8MӘ���4k�T��>���N,.�e3�o=Uq���(�|����/ޙ]�il��7�t8�^ʾ��7Cr�����vF�M����޿-��-��K�]y�j��ٺ7}�������5�fՎ��}46�{$fr�Zn;�J�a�u��w��U�C^����K�Þ�r�#��\ɱں3��ؗB�y�ǆ�Mc%�e��َ.5�I���}�s�B���/�	�d���DO���t�q����ӏ��C9v�5{?=�~@ �g�ihM���.���|7n��T9��;GD��|X
�]���Dl��>��t=�S��,4k��3j*��"�kbzs��}�@Δ.�y�rV=49g���1�³���V}�Hv��G��b(�@�>����#燛4�]C�ǪvL�[���W�����RUw��7ȗf��Ҥ���93�Ef#�<ೞQ��	s��W�m�Iz9g��%ڦ��7�r�!h��7�!"���k��H/	�!X}T�-�+]��6R�=1��!�e�P�N��4G7�����'��P3�bI�,%=�6�F�ߏu\[�=���c9�aQU�^_�� ��/[ND��@�T�l�K��1�)� �w�Aqȇ��מS���ȹ�H(���R%��G��zn3�����6rK�r Nj$�����|����}u7h����Na����\J�H�s�V��a��=q]V��Ϫ��pB,�5VdPӵY+��Dz�;v߁�G�t�z��1�z4�-�4�Wi}2�47���uUqQ�3:O��e�Kz:��z�G�U�$����B�x� 
���v��gǹY�zq��uF@\ù���y�B��a+.s�z2���$��Nي�{k���5~�9j����M�֋Q,w��@-���΍���s7�z��TF�w���6��ȍ����&����j�����:�Q��7�����j�z�Q亀uo���������z�,�fg+�5�E����٘�y�aliOd�m�Ӈ.����e{�|���5�^)�PG:�����t6�����oP9<�=>�s.�u;�� ,Ι�L�����5��e0�+����;�:�QLI�Ź׻��qkk�Z��:�vw�ू�pJ���XMYޒ��Ku�[{K�յz��G�un�b��h�� s�'��/C�3J���%�l֕�k7Np#�-��I؞�d8Ga��
{ĳL����;$�Y�್��.����^f���)��`�~P^~��y��~���v�8�����D��<���8ɜ������\s��������)���]ߺ%d[�Xx2�n����v&̳,�ڽLN�!Oo\����X�eB���Sq�}WP���[�g�5�Ow԰�'2�������a���A���/�uD9ϧ��ވ6���jry]�͕�e���8nD��-�۠��Q���L<�3��3��9(����`>=�i��ڥ�=�<�͇�y���<�zD��i�-��'�(�֘���a]٭F�U�_���o&?T�/�>y5Ư���ޑ���t�v��Ws���d�͸ '���zݘ.=l^�f�yu��k%Eu��'��[sS=�8�ׅ\�hxd'���1e���@�]U�h,v��qd<�>�;[Bz��� <��1 � W�vW)����^���'��{6�o��n��r^�o��{���Z�����u�X�O[�4O�um���ރ,����>v���;�"��4zؙs�����'+�Ϋ�=�@�ճvvdժ>��"j=X���q=�P��v�x�)�͡/���y-���j��Ί��0V�|}YNq�˳�}C0D��K�E�/b�d��.0󴁣��
=]�jW�5}�d��g#�Q���u=��[��/��Ɠ]��EOWX�R\���$���\�|���@47�s�y��)^檞��ۗq��<��k��Y�9tD{�:�;��3]S
��7f�}/k=3�y�9\�߫�5��1}��{�̧ֆ��ʤk����#ݱ3�b,�|��u9�s�U��5�]s6�޽�S*yFr���|��B�<��c3��E�.F���Wú�:��4{�9�ol�&��Q��b��d"<��Ó�7�],�q�C��w���]�zF����\gr�B�f����L.���~��"��^��7�#|�w��������_z�/�Ki�����;���1�/����;��1Z�;�� #+��L�j�c/�d��i��y����q�J}����{�X�俆�Y�k#j�9b���t&v�3�2zgSu2�����Q�W/}���Vx3�������&:�w�Ԯ7r9��s�P�RIU2��_�m�'�~�g��5�l���
g6D����W���c�<z�|�{���w�ͣ�=����A��t�Vs�d���f�vHl)�}�}R�Cb=��1���6�z$��*Ns��ҁ��\��n�m�y\��!�{Zu���7�	�%��� A�h1N=��b:l�pƞ���s������]�y�7����W謑��t><A}g�H)�/Ꞥ."�Zs�&���ϳ��F�u1�|�O�{hw�O��fȜ��)�5�v�K�������$���D����d�l<y�B徿]��TMX�n�ʭ�4�����Kw�=_k`�Cv��T���:�1�$�@Q�\Ud	���vؑ�W�Q�>!���՗�B�>�w�6�N����o;��_��lM���� ���!G�|yy׵_�Z�~����H�3�[u�oEY�BcRt��Ni�>=��7��s�|e�̖=�KSd��VԌ�8����v��UJz�I�pg|q�^�P�W�nO"x�7��`s�d�uu�jF���dSɦo�ԓ�<FW��Y���^5~���C����M��7�={��u�L]�_t��Z�ɺY,��r��Fg�}d/��:q`-�eS����UXc���:�z���#��.����ym�]�"�oP�@�yfJ�0�a���f��{ޝ��S���3|���t):�г��Bޠ�\gU�;9�46�{$f{���n;��
�a���Y���zȡ���ᶉ@Z�Ÿe[�s�۾uӨCt_�/���}x�s	`�hkgl��Yu�C�
�ݬ�������D�:Xr��{A,^	Jl^)76��&Wl�|�ĩg���{�ה�U���4�NKk�/�����ϙNd�_R̹MΛY&N�wy|�NM=�����N�,rK�9���;ؗB���n7�md�,�;e�[��Ng^�&�^,�*y��#�O���7(vɜ��j��8�s���~>��y��^�,�l>��nv���M9�&Pw.���S���x����ָ�ϝu���ˍ��3=�0��\5Nn�x�KbJ>5ԏY�_Y�P��qS<�Ӑʿ���/P�:��}]�kм'�2�t�F'ov}���Qx�����iq�8I�dv�L_�2�����<�<�Ou��?{���%n�>�[�}z���e�6V�@^��;N}�y}R��(���l�a�l�T��팸������y^97�裮��t�s����zo9Q����v@��.܀���Hn�*rX�	��-��)�P�:� ��<��qWݤp��+O�H�ی�=u�l��>�����b]!!{o;�8R�\m��W@���<+zi{kCȗ�ٌ=�|��N�>냷�wƇ���&X6蚾^ƨ
����#�b@�54.)���D�R���M_0�+<p��%�w�'A��"���c��A{q��v�,F&����;k�6<3'QRUa&==T�-sz^�s�#\C����8��B�dB�m��8��FX������NR��5�9Y;�Z���rSq�����(�����b��Y9����n�+�n��[ן�P�w6R��>fUrD{�[��}E�M_ޖ:��!��U��+����7to�z�9���؇�P��tU_g]r40�=���;�٘�6���f�Tc
q��Z���U{'��sT{��Wup<�fhz����]XfU�a����K�w��[�̺���N������3MR��U�{�Q�_R؟w)��&�S�� �Q'��
�o��ޤ�C�3��Ó��7�:��R��f�Y��|�D��~NϾ��|S'����'n�C)�v�M˫�fw�e����rrO���Y>���'/�!�UI�=^ewMqJ�v��/��n�?��;�k6���Uե�bɼ�ȱqY5�qN@�z���^.α��C�Y�7�w^���j��)\?�d>֖�d�AF�3�6�\�7N@k�dpT�=��Q�z�b��X�_�%5��7���r�]�hpܗ����Ag�(��DIhѕP��4�˙D�ut����7�x��j�Y�����#�c��qܧ#��ȗ�����.��(U}3�(�"O��6S�سb|�N��c<���k]�.��L�ٮ�l[��e�x�K(�aE��ww���r���+��f�vWd�k}~�F'fy�zv\� :��7e�c�"�an�;gqa�ĺ�5pݨ�f���7p���ok4��}�E��n<� g8K�0�zk���0�m7����"��ϤԈ�}gP\W�h���q-ђ�sf�2��1T�k{	&d0^uL�Gtuϳ�u��|Gd���/*��  ��&��wG��졃r�
�瘱�]%ؓ<��y�V�c�:�K�b_B�l�/�%ȝ��*���lÈ�pa�ͼl���t�T·����u�g���yHkj���â�7.�a�hVp�z]w��\�>4˜����6������n$��?�N�1����1�{�ս2`�I���E�mR̃��d��&L�0Q���y���@L=��`����Xd�=$*�I������	"�ǂU�*S;}��T���$|ޗ���^�y���ӹv��y���#{h����ͬ�5�`"�!r�ԓ3 ֣��!4�G;Q�3��Z�#���)��xT^��� ��U����~Y:�y���;���{��[�h�4�<])1������GTڜ�؈{PL�_:�d_3+A�'Q_�F���%]��m�Wr-�L�f��F��鈅�Ӱ�c�nS8YK{���t�ǁ�p��o]�CWyw���93����u�ˎܱ���Af��sW�cD=q+�ܕa��ʁ��`����gګ���Z��S�ǖUꕪs��R���݋�,��}(GN��>+�W�T%�v?`W��z����pO{<�A�,Kͩ	s
13}\/Kr��R���`V�4���2}Kji�--�j��l�O�:��
o�Ӄ�ʱW�9�0��c�ڥ�S��9�
���{���r�`]��ޮ����%v��cc�ᛧ�v�Թ1��g^na��u��N��2�@b��-���f�㎯F�aI��ݝ�a��S�wP����L_Vc����y����69.����/�V>�k�N<y\Nk�Ε�S�V�J�뛖��VW<�lv�+�Xڛ�le�Y]�i�f�(Jy26���k��N��&��d�|��%��|5�VѶ9�]��ɬ��c��ʏ��,fWY|LYwy����&�b�})ܭ6f��жf�l�.2���P[}�5�4zRAWR����q4�7�d�;��oc�J�.��޲�ۓ6[ނ]�\��AIr�k�a�hlܻ�����:aƂ\�>�
�Xi��
����^����ܱ%�=w�z��u;<{6���{$��!�x@�]�dH�;�y�бl3<|��h�5�B7\y݁��r�;�s��V8�\��X:�[|)FxF�X�0�5tΚ��4:]�o�����\�^��=}ƞ�֭?b�	�8D$�U�Y��X��Ү��������upb�x�J }T �QGBr�k�䓳�Q�ᓤ���q\�s\��\�]݊�s���\�wn���Uˎ\Pr��t�P����*7wt�W"��[�ɺQʹ\ܮ�w]�m;���;����L%�t�-ӻ�u���nqwnP�r�5Ζ+�$�t(���5���N�r+�ݹ��� ��N�]�N�rn���u�L��j
�Mݸ�Q���u%Ic���6
��;�f���w:�Ĺ����w\v�s���]cwrU���]ݺ�0C��p�f������uC�Ib��E��wu��q�9�����(�I�]ѥ˭�n��.�peˑ��Q�MT2�#Y��wu _�� k����v�w��V1]��]C����:�|�޺r�]�{�㎯�պ#�!@\�'
�ΐ'I|.�/l�ud���џ��T�)�=)��M3^n�
��^��t�v���3|y|6pK2��3`]cҖG�I������%��yp4;����]��[ݡ�B~�h�����>�Ėf���y�>�w͐é�{��F@���vW)�n��ף�Os�2f���}��[۪��l{n��/����p|n����SR��"P@�N��/O{�Uۄ1��sP`lޜ&d��k�T{/�@ݖK�t�d��D��D۪��@���F�/k��zr�E$cv���^ͺvϺ�G��*5]E>�@�|:��σ����m�_T�$�;6���\�d��������R��]�T�}E�Yc��C�ݪF���(�ܢ=�4��&�03��-�=�_)~êm/^*��;)�Et\�l�f�����Nu�3ח!.�������K�w��a�
�.���8���lY�y,��=��0���'��`-�K�9��\l_��ޱoz���uu<�xa���fzT��rf_<��k:�M���0Ktdv!�_k�il�.�[��[w؂%�O�Hp��]���Y��)PÌ����� �>�����yv:���j�;���{�Z.�V%w��n�V��7z�-�b��6Y���)��펝}:�r�S�vLs��0b�T�̐���t�K�fN�O�X�]C�zS�6��Ih�Rۧ]�z�/[c��rBB�/��?;���fϸ�w�8;18��7J�&�dr�~���/�T=ɷQ=6�N�b�����U� ;����{�qg�-�}�Ad.��~�[Ed\�(z�^3�/X����h/_li��ǀGw�3�13�!c�ǫݗ�gZ�����:�(e�$��9눉/��o%�^eo�?�O�ѲJS�!9zg������=GOqY��;p��zbz&s��򏖫�4z}�f���]|g@����R�	��μ����8����,��~y�!2�]�v�n���VtF�f�Y7*x�(��΁ �H��Kf�P]����[���`a��e��쫿'���vi��qC>��R����;>�<m�:�3 7 Y�\U`�z\?���<���N�NWD�J����|��!����Dz�؛�}U=7�9�|H�%����^}'�]_x���b�&O,>�1��������9�4�y�{��x	�\f�%'b�Iܙ��^�2��_��\b��Mp���\T�`<�/h�w��6�y�q�'�2�!�|LOEv�p.8U�r�Nn��y�d�I�� ��R1J��>{��2pTF��we�m$�ԭ���b�%��c�$5�,H����OL����M�A�[��3�������;T��g;6����h�̈aT��ߓ[Ҿ���߹q�,+���9�*��&/�D��7hr��3��#6p5�o��Ҽj���kw��ڪ�	��G��5Y�ï��5�V'|��m�
�Z4b3�*��s��-e`ا=�W���T-���%�t=����U�x�N�[{�,~~��{���A��	�솄 =�FNF��zs
�/Ƿ#i�v�-b�y�Y�Uu[S��.���U�Q���*=C���]�����@��ҵ�rb.\fQ�cK�:��ءr�Q��q_
u�ȼIs&�j��6;�^�:���M��ٿD�¼�w�[�'+����3�閠:�z��M�L�o���ʣ�>��N��﻽p�|��q���:��x4wfu�oE)S��L�-��e<�����v#ghB�ug5uw}WC޼�Z��'���󃳶��y�ZlQ�s(صt�qS<��9������X���,�A������V߫�GgKjv5���a��W��I@�"
�6�R7S�<yts+N����9B�Vz9�����{��#�@=}Lw�w:���f�D�_��9L<�-�����1y�����PO�������d�@�PE����s�^�����S��B��q�=ǼWv�� �:Ky���h���b���yP�O6�Fs��2VngY�UG����H[�.vc*��V5a�fŧ��p�и�o\%��Kl���n�9k�=q�{/�S�\��Lvϭ���)#;��>���]�� ��D�t���T��}WgBr ��s�]! �<�B���_�-�G�ⴾ#�wY��f�U	�4�z[Le�<�l�UGg�d�S�wJ��_B�և���1�{6��GL����;�t��S<�][�9KQ�W��4;�U>7�!� n|
jhK;�4
���w	���}�Y�c�e�,����v�N������CB�!���R�i�fW$G�U���{_�c>�Nb�媈`������剾���oP�q=c��C�\CԹ�I�5�>��f�;Ů9>��X+"����yy���|1�=��ݺ���#�����T_�Z󕙜���o�7�������.�ϫC���#����,��]C��^*��o:���qΏ�oz@(���z�s�J�tu%^:R�x�3�d��V�)�K.3��רm�̋�೏�g��G�׾?��?~�+)z��79�v��̭<��_L�b����M��p�7���}�b�O c��fu-pcr���V+{�Tw�i��L�d��Q��#,�]��
 Ԡ,���[#w�-1F�	�s�4Ӛ�fh��e��n�bK��\Sϯu��Z!e�}��p��ےxd��58�I���l�}�x��� �:Y��"�v�b�m<o+}g�����g	�2y�'��=��?dS�t�o�,��j'��R�L�و�q����_�w�7TdѯM�f;n�}�:Z���:����(>�R�tp���3ڇ=2��٫�8&柲v�tnn<��7���B�S��ep��Hp�wZϞ�EQؒ�L<�dK�]��$��缽����z(�Ɔ�.���ˬ�}1ǝ���vM��]����NIl�$��+k�<�nʎn��0�Dp��6�S;�)O,�`m�ҩ��3�1�Y��}__e���|y�8�[(�|oGz71�5T�:������������}.�୉n���O�moHg��E�:r����;��+�df�<n�2�-�(�SX�գ��{����jm��N�o�����]��}V�7����uD�MK6���	D�մd==�a��:y�t��{s.g��[�+����.��;��NM��N"��u��Ir�d��@��wˑ��BN9��Q��7�ͮ�{��:�m_Q}ҁ��`}�u�TGu�n���Pɓ�;�qZ��|[���Ӯb
���C����0j�M>�r]
���wz�`bta�$�}RS#����0H;e�gA%���èTRr���n�N���\����w9�嗆.�r���D�/�aE��W�9D�{��a�0Y-��KpwU��ݷ��7�?R�?B�>��q�_�Ά���#Z�x�hor��bd_)8Gf]T��������P��Ǫ�QѼ6p)+�����qo.B]w�1�EuΗ 蛶}"���s�>K}�7�;:��e_d{�h�4k�ɂq��σ��p/�ω��P�]�c5WnG��J�l�S�޷��y�3�}Ax�u��>����dv��V�Ɩ˂魈��(=x��]y8��{>������r;WgM��GfK��>�J-��Kt���5�I��w��=�k0^���V��|� Lf�dZ�K��u\5��ϽH,�w��:�+.p�<K�w�r�q��RcF(�.gǑ���:#��C٫8�c��q������{�W�������5h균���N��g�Љ�FW�g�D���{5���z�Tc�<z�>���C��}�^J49�G�a�>�O�7g̦z-IQ�E��T��O'9&��>�����a��>^އ'%ݦ�ǥ��t3��y�-�5�c�nT��$�3�O�
D�ų�Av<y�CnX��w-��k�8���^z�����C�W�=��Żdܮ3ǻ����0���=m����^rE~!z������%ڢᐵ2E��w�B���/F��N���&ŗ9TG��m�:Ŕ 5�x���݇62Ü�
�a��������B��c%�x`�[��k������H��Cr���"`���-�eqU}r��/s��-O�=�=~�q7�b�+��>�4���#��u�>��� �����ܻYZ+|��Շ�w����q#|V?B��t�Ǧ�{�<Ӄ[�N"��q����S��y��y�iI*�;S����LU�T�>�񯗴T;��}&���'�A��'��1M�+`�Kp����E�O��$-�b�zw����^/�z�m��1���(ñ��{�Ń^p��u��Oi��~�hXC؍��k�ˊ��B'�B�wxg��j��ǖ�Xc"·��+��l\��qY�ޡ�%�M������C������R7��Arl�:�{��~y�����>�\vz��,v%�67܇����g;������#27��pr7ި{w3���#{���e�.l����g��4חG�%����8�b]����[��4]����U��ͮ���T��}�V�57J�f����b�dI�����2�޸K^�Q���ύ�$�,}���Ձ����T�����!��9Sz��#�U緼�_W��Sɮ=���H�7�_K��<�w���y�I�*H��������#2�kߨ���6{Ŝ��\�,����j71v��S���(k3p��;�]-}B�!|�&<������f#�"\-��Қ�8#��O��Vp+�]k�=]�^ߕ�C�w���t7�������E���B��3�(����#t�2� zhr�pח�d_�s�MMf!sԲ�o1]i2��C��F.=��e ��"
�2�R7U<x�
��j����M����x2<�{���@=}Lw��yH<���f�D�Fc`LU��c�IC6�;�5Nߊ�cU
eǸ��/]_	ݮf�;g�(���9Q�������9���;�$]u?)�Y�*)���T)��b�*n�(��+O����=u�l���2�:��=�r��U�X��<_D�0T
�}(T�a{kCȗ�ٌ����K2�'��s]��l�j}���F\�K����G������(>f��(��+a�"�[p�~���;��y|Y������,B��&��\��!��;f*%�udף��.b�>t��U6p�fV�˩���:<���u��3��F�qА��:둯��=����=5���~�b��(~b<ɍ�zZ4��[���@�P�����V=|#y��ѫ���3�3+)�+�89|U����@�W=#��H*�B�xz]gc�̧E��u;��������u�m�3he:��x�ׯ��!��C�|��f�+�.�m������)5��]�<����ō�T�k�ʀޮ����������]XfU�6���	�5��*��Mm���Y�G�gֳH����̯����Ϊ���G#WԶ'��G��L߾�6Њ����
��g�;Vu�����p��p��z٭����*�2���+��'�u�]�]|��Ό�.T����xMf~|����ޔ���.��F(r�iM��p�&�s�uޱ�bY�#���%��R��u������{O|�W�=Ռ����^;M���{� �S4�@�q�`H�M�f]Mt=Sh�p���Oh#�]��3����^����=�(/sۤTQ9�F�_�K��m��꽚�/b<�ѿ^Kz�3���24{����^t����ep�v�ȗ���>{t\�J5%��d�ǮT^>�m�*Z��=�gQ��&u�S>���s�#�{#�qܧ#��ȉyh<�>��eHwf� <"��v��:A%��>~���鋊���Cɦj���x�oH���C;y���+���і�Ա�;,Y��8"#��΁1J���.*e>����*�C�>O�m�S߹F:�˦9�DВ2�	�x؋�{�+M�7�,�V�8i���ڽH3���P��b���AlU0Iu�{f5aҰ��z�7r��6��ݳ{�F?g��o�x�<���la��G����ےOb��G�M\%Q���jl��l�����Rs;�h="�al�y\�gܽ��J�8�����A�6`�J�5�����z8	�z]�yS��R������8��c{��%Fw\���:��P��H$���t\��~K݅��r����Oե�"������=�:p2nux���țuU�7�-�F�h�ޘ�5�t=�N�T�wFF#�ި�4�
�pھ�o��=��DC�Q�ꮃCR�R���=�K9z��yI*��S�&�O�xT�g(�xww�p�uTT?K�h�>�{!���k��{wp�,,�{X6��(-�l��8��Z�B���(g��ng$�Ϸ�#��p��S���Ys�.�.��9�+�����"�ѡ�'\��Ӎ��.)l�rb��̒ǆ|׹��{�#�� v�p�w���{ܣ6m��3�}Ax����l���0Ktdv(��ٹ�|�\~��C�3մs������ :��lgUu�9	�.��J�̖;18���P�l�[�6��؆���2�ն�\�|6�ål�;��ǩ�'VE��\F:��������Eڼ�_�6NC@��4JB|���{K ��}[���]�1s('%�� �V�{Cx/�\uɱ�{�og{!Ӛ�fj�CMv��BB���}���w�YA+�c���C�����h��狙kD[}��&�u��i�6���6x7��`����P��������������Ag1��<�v� ��kz'�.�T�yAS )w%���4.�Q�@۠��d�fÂ�{U��<�$�.;mbt�Pז�B��X��Аn+�W��Wt�itc��<4����<C	̃q$7��1WS�%�$��{Y�	�;�Θ�E�z+��yy9>��4���f�W�vQ���A�E��<Ɋk�ZXgf[�5tB�3�#bPvx�ZD4e'��V�M�]L=�f��)���vT0:=S����\=�u�߶��wgE��k�P�)m���'�a��8��p�<�ٽL׾د��Q�5�oOx��ٝ#M\�|�
8�\��|{��un[G��[�Jz���`oe�]I��K9q�ť��n(�=��|4�c}��;x{�杼B{/�d�D#P���Pi$e�}�s��7��o�f�U�9��É���&�sC�/�h���z��ʳUވd:��v�Oj��M���9���%��1(�Y`�����;�S�k�uj���K�B�%����%bX��P�z��b�S6���"+�յ/v��)�hM���nl���yкy���	h��1x�d{�����tԶ<�)n��dӱ��;����1�K�1s�Iv���Ѓ3��w[�Xt���{-��%��/7�vT0h�&���u���z{�*Lg���i�`������!�(P'K�Z򌥢��}�=�帪�fa��RQ}ڻ�+�9�27�3�%cJv�ŧ��WD��t�s!/#*M�a��YC����C��Y�˻�w0�֎A�FW|j��:���9SY&f+C6��{3�<Dw}������IȺ0P|1Q��&P'jBU��\�j��u������'"�{܃�>D0���8�I�?k��Kς���mYa�YMuuƐ�\��ŗ3g<�l��sS@%���Յ���#DGNuX�+T�t�:��ۚ��@��z"_o�Ɲ�.�F�~(��Yʹ�b�xYu�J�w����cWN�\Ҁ�� J�+1�{ظ�;u�u�����ԧQ�{�}z'�{��0ъ���]t�`	��t�oT��RS6��7r��T��uά,2�n#`a�;�Pe��^���}6�	QW]oƉvԆqz�Ǥ�_ϗ��T,�ݨ����)�"�{,���Ǽ�u�LҼ|��@�7��%=�Y*E.Υ���&ݴ�P뛤;�r-$i`4
�4X vQ�J�F��:Tq�fA�b��O�'����/�Y�
�L���5�˩T��Y���:5�}��2^�S$@�zї����Xv���x4���\��{4�C0�v����n�߭Uۘb�Zj� ��DAĮF&�\�%JW;u�"Kwv.nV]�e�$HiΓfs�b��@�AwuwuB�;D̌И�EDDXأ7wL"��"	+��5ˉ!�Y�F3a�1DXw\+��']fDFJ	!��B���ۻ�f��ц���&���c%�RXd�1�m% ��hbGw(�8�(��B\�Da.t�v�\�F��K��Ic$d�wnd�%�f!"�lA��!Ҕ#��wW@��bb!0uқ�����ܹȐ!$HƓLs����*P����͌��A�s��PI4��ܮra�Ji�������"�3]�]ݎgU��t3��qʩ��ع�,[N��j����S*�1��hC��
��x)2��L��Ʈ�<מ��y$�i���0:l����W�F�g�x���kǠ*��t�+�W]Cgz:���s�19�B��_�6t;U+�|z�������QgG]L򘸧!9�{5��iꀀ��<yޞ㚣)��-��t��{i�J���OEg�f��5�>�$�`�,IR�����<���>��r�l�x��VҞ�鳴��s�[A���qێk8�g�r����Itg@��"�Kf�P]W�p<��s�y��^��'��8NwS��v��q��Pϯ� ����:�{*x�̈	�����.�wtƱ���7�^�>��9\&5���q7��1�W#��G���#:�퉷�S�p����Y7I��(t�3�\�x�B����#|P�no-�i����Nou8�Ҹ�x�]ҫg���e�Z�O��W�'GeI��� lwJ%��� �5����j�M��D��=9�������f�=X��l?c�ٟ����95��$G�p5���q�Nu��r1���#�����mW�����e�E��z5v#F!�\�X���B'�B�w8���2��ü�gc�ol)�L�W�L������!�˝�w=�̌��??f����s���'���Pz�}q�$���scɐ+�_�g����XnK���w2�v>��WAo���\�]�l�B��rͺ��S#(cjڏx3���Wg1(���JV�z����kl�ܕ9k_�dp~�ϔr�>��	��Ѕ�2r�����"[#irl�Moɦ�Tow���ݥҶTWj9~�0VU֎�U�q�P�W�V��t��w�"��@�@����\��ŏގ�^�'�W༷u��3�W��ձx��M殌�}�t/w�\{y��~]�{(�51S�9�F
�\��|&v�%����dv���tD�v���g��{N?����wmm���|	�Bܧ�O[�jz:ɳo靋�2��.'H�8�]���]k���8��q�uI��y;{O,�-9�*�{��OH}�$TY�R�2�P3����FY�Gl8X���U{s�3~Ƚ��	Ml��HSr���;p��b�=��AV�c��*���H���h9��nc��h[�!����O�׃#��}���;NK�A��T�l�K�1�27�.��v���k�Sf\_E�d�:���[��\G9���@=7ʈ��u����Z�4�]�u!�fv�Q�]p ���Gu@��q���/N|��qE�H���������#��'��H0�&Õ��[ ��R�b�g3�6��t�Oo����,��W9�uw��qv�c�N�K�]�t��"Wf�!oz���{�+�/6�����^��W����^��Uyk.)�v���n_U�<��eצs���%l�KBp��Z�nN1~lg�M�� �o� l70.�҅`/N-�K�l�A��l��P`�����u~u�Ovl���I�ǒKǑ#����ܘ���g��U�d88�}a�.'�������2�2�F���ǧ/ uF@��뉿�MuIl	�1R�����5v�O.���m�3����]��!���YsUT7��q=�g��`w�U@�]��m'��)t�bM��>qؗ�U��j�n��c�m�ѿ������i�����뀺l̪�~�8�R�򭮛��OB�(�g|�6h#�����*�]����}�Q�κbw>�M曳������(�e�3�mD(��eC�J�C���/�s���6�J�E��YŻ��H�eʕ5�}Jg6(��{y�]�����♱���Bg�`eư��q8vv#�}�_{�S����w9(�y�;�:#���67�q��/Y�}n���d�_h�E��ɯ� rb
�7��]�m��/2�W\GW���]�b,N��c�\?����9��%+3;0�Uһ�hyt^��=Bm�⑺
���io6�=w��3�ڻ�(�����B�s����>x&�|M��缪�.W�#��LT�5�f��1�r-Iv� ���;͗h��#�FӼ�ΙlX余��bU�����\��q�A�p�����N���V�Q��w�����w�R���Ψ��V�J}k����#��t�����Yr�(���C������wEW]���F�-2��S4�v��#�{=��r:�pܗ��xU��il�;���^�}�����,5P��nb⧩3�&���7}�oH���{�3��#����>ۭ�!*[4��⯶k4���	�p���:�(�Ē�Kx�®%�C��q�O������V�ΟnR˭��}H���\]u�0�eO��:��0d
��SX�ٻ�;�;������]�� �m�����;���uD�MK6���@�4O�umbaJ�l�b·9����&T/n�>ձ��a=`GMƓ[ܜE	��_jK��`���s�����/_��vL��E����-SC����Chn�r;�9�K c�����g�.VYݱ�#��5"�>����!=��PS�Z5�:�n��6���|�/��o����c��5��f}Bq�����man+�[6OFP�M�PS���sЬ����2$�B��~����Ǌ��W,A�^�퉁J�/n�`Xu.��ݰ�*f)�6�/u�w,��Y���,(ﵴt��K�N�{7�4vA}s��ap���T�xJhӱ�ݶ3i���3=w%7���͛)Z5��k��V��͕+c{��rv�@=<�j�z�}�.��u��)8f��ꁓX�xl�fᅲ�t����R����οn��+�ꌎ=]���N���|�	g�w[��~�[�#�D�Fҵ�9���h�F�,�t*�A���p-�!�$���WgM��GfK���|�(w��lv{�.�x�n��`H{v��P]���M�E�*�L1��"�UԸ���p֧ϽH,�޴.=ζ�:�m��Q>��hƂٮD�d�0\�r԰�GDv��A�Q�f������9�o������ｓ*b����gX���m2-I%TD�
�·qS<�/�r�{5��遱����}~���1Q�ޯ^�m�yggKT=ϋ�F���L�Z�
�3�@�XʕH]T�r��u�.Ps
�Ϊ��æs6�hh��\=����ϝ�nC��1�7*Y�e]�$���*x[���'�;�{S�C���,��Wu`]���}�C�o:�>7�u��`ܩ�l�	��c`q܍�w���ў��Ц�x���z��i�ި����/+��>�M���G�+�؛��S��ԍZD�`�[�`X��Z4��+�����v���5�o6��'���6Wm�ي�K+Y��.�k�����2�8�`�gH
7G���}�!�)yק���2d����ē].sWL;Ȃ:I}��s�zY�M5�w���4���̽J��?ܴ+b�3Օ�����G���P!���`L=5�����Sdq��y8
n��p]]�btڢ�1ߌ���O��Z��@��wRqR��{ �{D��m_I����O����&�K��mG*�7դ��5�V��H�uu�o�2CWj�gx���.�eS�e{��=o|�Uf�Rͭ�b���Qn���xwO�X�B���1:�#����Y
w8��y���}^�s�y^�=����k����C�����՝a3_vCB���ʊ���ai^WY�H3uм��c�-M�U���졃oח�#UWiϞ�5FuXs�}ңݵu1L{����#,O���=Gܶf�ó��C(+[��:�f�gx�^[
f^�xk/fX�wn�c=,g��g��ة����E�h� ��eЙ�(�QYU�aq(�p21s��&W:��}u�+"Q�ۻQ��k-Ώ>y^�OfڟE�Ñ/�t��3�?!����;���q۝�bR٩F�xǲ��a�5՚q��t=���}����'2��Z�>;�a�1���1�۳r�~���=?.����Sx��n��Y�H�<��͉�`�%5�F��g_>뭒��յ4a8E��,i�+���Z��;6�c�ǒ��jvjqϟ^���2���e��wz�m�:�-���,eXh�z��r���jn��2��'u��VՅ�����.z�oF����í�ϟWqY�Hv�u��������*��r4eS��Ǹ��-W.��Ř�*h�UN��.����(�tOq�{�����9����K7�(��d{^��cW�er��и!o��FwM)���{v������9�纀zn3����<;��|}N�F$��W^uɻ rG����T���E�ŝ늹n�!��WϤx�\y��S�y�vv����ʿJdO�"��fu�}(V@;⾼��m�ޭ�$���������v�_]����L�Mޠ}_uUqQCRS��U$5b@�r��x��=�i��C�V��oV_���G�_{��9���"�w.Btj���2cr�J����4��,��OW��ئ���O�-TCڻ�i��{��3��`;���]EOiΏ]�+�]���}��mMT��:�31�6�CYC=κ/��T�k�����{!����T�m���|k"�Wj�Ff���+�{[~c���~5�ˇ���W�z��7�t������)����vd�o�Ͷq��Q���X�|��=G��2*�*��veN뱏YN���0zOv]�R?��<��I�=F���%^�����ޡXI
����t��b7��q t�쮚���${]���O��6)���=L���,�@Q�g��?����	�m��z��o��V�:�f��(S�P��d)&�1�N=Uj��/ۏsc��yUp�����P��\W��˩�с�E�,�ĺ��^r�C�B3��7O��[��!̽�˫�o�W��d>�K��id�heyP����Vk��>^��ƻrS1_�\���tz���.!S]�2]wt�SQl�w5�A������FF�cg��C7����GC��)��=] r���ϼ]Q����ݕÖG]��r"^Z����bW�C�=�ou �:I,����2���n"���{2�_i�c���u�r���\5\�ͷ����]�G1����~α�=>��P$����$5P�*e����L�2�o�n��#zG��;�u[����?Kw�=_{C={*��Ǧ�tӂut	�)@�<�Ē�N�u�R�b�<�79�LXsݮ4_z2;����X�L3��@�������O�A��@fl�_��i�dX�c�l�齄���u��|팈=�|7���I����u��n���������q�*�4 �~�Ca�śk�6�)Kkc8E�6��VV�7�_	@ka�wuyS�ĩ�SUD/�Y�p�d}o��!��纏u��#��ฦk�"�]��g��v͙J�ǀ�]�k��Ѓ�:�L��״~�I�8%v��|yI�{2�j�����)ϛ�$�?�~�N"��U���\'����H����hwrq=}bkR\��S��Q�S�V�'Y�'�-Ř~�F�;+*hL=���}ԁ���v3X��m4���kۘee��=�W�1p�NdǊ�ޛ��;ţA�e{��Ĵ��;ģC�ރ�sz�yV42�:�i��虊��E�Y��̓Sуƣ�S��]?W
��/Ɩ�\67%���-�������
�vY38-F�������:�E���q��Ӎ��.+��t�Z�Axev�˅U�ղ���{�m�29Wz����k��Ze�{���~�hA�T&����x��v�����3K��ҍ����@��Q�-�p�T�AN{z\oMGx���x��C���mٹ&d�剻��;1��W�Ƥj�J�|���S]#+�zW�xyl�>� �z�舵�>�᫸�� ���[	q�O��#"�ς����l:G�x:��e�@^o�x�����L������x8�~�y�g�L�1)�d"�&XU���S�e@�+�XgP��U�����V���x.�HL/��锼��X:�W��tS���Iy�zNT�Xh�j�ӑ.�+RH7\���/�>�:�{C7��wq$�^�&�~���:I}O�W��%�D&n�&r�[��f�����Wo���!yn��}^;��yVs
IbL����M�*a��E���;×����zmt�4�"A[���b�RS��MG�=M�S�����y5�=�yu���<3:B>���!�`�]J7�%TA�A�`�F��hFS^�FU�����S.3���
*wz�X���|��q�H�����"�5Z2%+���Y�t�E��5t E#"���-�A����G��gu��'���4t�[�|���A��tNU�K�b#�A0̃��/��i�b$o������9���<���66��jo�w����?�~j�f�%'�$��1qq8��v �~��ܮ�C��B��~��E:��u���%��XN��q�_@l�����#�(k��-�XCaW���ri�}�}]���`�E�1��Iݻ�b���>��P��r4bu�F����O���8�.ߜ{�uV�N?d���W��+y'wB�~�S}��m����=P)vY��\���Bi�}f��ݒ/�Z�����K[f�-���t8���gF��qT/�FϦ�t��}���x|��1Ew7�����ߒ��D���t�)و�%�N���ٷƦ��nֺ0*e���'׹|�\lĪ;�)n�1F',���ڧ���b�L�;�H+�0�����<֗bwe�r��Z��Z�u��z���;����R�4F_��Te�4<'��X��y&�ڠ����
�fV)O;"^�aӀ�F�9-9i-GH�Y�f�4�h��.C֎�(�g�֔��.V�T2G�ip9���E�� ���m�v�ۘ�K�}����ȷKpU���98a(c㹠u"M֌��k�\���y��|p���@]�Zp9��Uhȍ�+˟E�{�'Jy���wb.F����u��	}Yw�{T"B4N��T�X�+�*Q�V,�q���ukM6��s�H��r{�U(%�4��;-w}��X9��	���1n��[�Դ��X��ZgeN�S`\�&�i:���4jVi�t
<�.j[�J,�T~+��^�!�;�� �Ga���4^�st/n��;+l�I�������k��t��9���Z��f��7�[
�m��J`�ዣ���J�Wy��.�!�D	k�n�
�˗_��م�E�<�Q�4��8px3�ȗe��u�{�@��[��J��a�)���p��]�vTZعt�k�@$�����M�t�y�A YJ���W+61�4��+��������jD8����]ͭ�+���ǘ�y�hUN�gu�%؀m;Y�,Oۈw��$'���^�_и�j����S�W�5���R�|l�����AN6c�f��:�4@���뱜4�iw���j�{�D6$�DSii�5�Js�H��R��uH�;�=����$oee덖�}�c�_t�Y����}ϝ۠;s������^1]�g����1��a,�p�sUc�]D�h�j=��B�O)��;��͙�7����D��viܟl�4�I�ʊL�����4߽�f�j��Mg��}�s��wȓ��X���#0A3x������b����!R0����a��Ve�B}ܕ�f��/7��^�Ne��ois}�<�97�2�S�Vд.�O�5����k����8]�<v�rQ�t��n����L0p�N	݀��u0:&�j(���Si��x�0:}��i�����:b�&�5y�d�h��;R���X�tB��|�^CC�ɛP}k('��ғv25pu2��f�����D��� �ja���c��4���r��y*``�>U|y���I��ˮ����F��O��Q�3��Yok.rY8��Mp|婨Y{É�����ѲPsn�Ŷq�Ieen�9V��&tڂ�ٜNrl(PݖE�2uZ��.򵜑c2p�(���\^�������y�{��$&�e%]3���W�)(_n����§#���l��R��j+'�}s��n@N�x"�{�i�B���
��;t.�4I�b2bT�nr����urF]�Q��X-r��(E&m '8��%#4h�(�L%0�"�CC2(�@ILa0\�R�]�Es��R�;��)�I1#
�F�H�v�(X�b�	(Ц���,&Y�)���d���i!�E�(&0f6D"2d�fd@J�H,���bΆC	wu�AC!B12X�Q�&�R�#�"L�wwrY��D�$F`���D$E0ibaA&e($�H�Q	H�IiM�($Q1IB�I)I"�BH�$ C�I������!0зw2F!���H�F��,)n�z��_
���GoBDs��q�tR�}V@��q}Řճ���
u${S9#�ɼ2����b��e֫�w8��k�����?:��]���{ƀ-��V���p�a\k��������v�p�g��n���z�Y�w�-��w�#� ��wYU�B�G��7��I���w���k#<��_��og{Y�)��{O�>�j}dٷ2*c�є�.+������׶������==�W����uw�H7ܮw�&{�6O�"�����6�ח!�j�����w�G0����؜}]�uJ��u�����п��'h�=#]��.e`����yb�73�:�u�,'on�#�=׃=�=���{p���9���@�T�*���&0�����T8������B�2���e��Lį��.��w#�@=7���H��e��Ŗ�n�i~V�}oHt��B02JF��:W�gz�[�/��8�4�:w�i��MF�V�$6k<�x3��=R��o��pB.��g��@���:&��FoV����W�55���&��=���Vu����&�u�ު�4=�f�����
�Nw��@��8�߅�i��V���d�4��e�����SVL��� �2r�l��,�v�v�zŜ+��e'�U���V�.��"*��l[]���5�4�)b�]�t��i"h�NA=�^�zgu��l���/�NJ��/Ň�����ߍ������6�:����ϋ��辍�d+k��{��8zq�o�2������+���1�B'���/:��bb:����$�uU)wFF,��O��Ȅ���}����g�B��P�3����z���֯��$��N#�� ��N*Oi�V����ζ,n�k\�r�����hb~}@V����*BW+fia�;��d�Ct�.s�E��^�z���j�8�������Z7!��l��׏�y�מ}�s���:�"�j�� �@܏!7Ar�t�Y,�9�
t��?����r��_TU��7}���O���'����g�����r�L��@C��&�O�X;u��h�G�9��]q^�cb�.��oW����1���҇�ɻ��҂��D ڷ+=lozz=�����裣���p� G�U˲D��u��[=�>�}����l����>�z��\S���UC�3�Y��
��tjt����ÖG]��yh*ҳ�fF��P��J�E����x�Ȃc�&{M�P5[U�枨��!���;��
W��G���E��;ql�қ2��-�nk�m�t_�f�8'J���DwN�E�Z�C��݊��}T`��S�^G�4����ζ"�]�%��m���6�Sb�-��^�w�+�g�vָz8ۓ���/5)��>ɇ֑���Ϋ<`wz/{w��%���_e:�;����}'�!��N�p9T9%'�Q�3��yu��T�3n-�}�mU����,t/HG��������d�Ͳtg@��P71u2��هf�u�Zs�ޭY�����b��cs�[G�����h�#lGZ�5��f�#����z�J� ��#����|��բ6j���y>��o;���L��R���H�C���.͍���D�(q���{K�i{p�.�la��=l2w���\�vD�s@W���!Y��uWT��$�4	�d�.F�;��!񯗴T;�����H��=�.�^s�/�J��鿝����՟{3���I�H�%�ʅ8�B�;ţ_3���#|7r�����d]^�ݬ~x��%��{>f�+��G�]X:���
�l�>�q@,�Щγ�:%ù��O���Ϧ��ӹ���s��tA��P���Y{�	�F�9q�S̸Ço۲�a��=�6�Ӂv�]�@S��ȿb�X���h_J�.���}�n����}9m�j����η���#�%���1N��f�EG������fv�9���Իl�q- ,����M]Wg���,�9���[Jl� :�s��O�h^������������bjwi�X��P����R��!�伭8�Y��6�&Z*m=z������p��p]���w�b��נ��\�s��4;OnM�������ɉU�z{C�ĵ��c�aS4{�{I��"/;p��q�kR�'F��o'r����<�<�,�w�f��}�d�2v��>C+����.�x��u.6l����+�^�f&�������uz���S�^G"��*��aP���*g���9���\R��e-��K̹N�̫c��^Z#��������WT�`S^)t�4�DZ�
�1�"��*�ݚ����[�g-��پ���A�ή��|9t7�^om����ЇJp�:IUt�r���cg3�Ϸ��|h�D��72�y�Ǟ}X6#��;����@����#u�!�`U��xp�]�2,D�����4��W���wr�#j{���A�о�a���;�.ۈ�������w�1%��q q�G�J`\Jg� L=+�0��O��8ߏi-g�M��X��nMgkp�U�����SLϝUIb�Ijl�6GN����[��C��i�V*�~�UW�X5�[]�3�}䉗�t�y���WK$�������pvk�+�n�\�r�p:99��%]L���a\�Z�M$������Z�X���y���ɋ�w��N{j��7`��is4�g���� �[붝A��c�Y���̝�^�R3/�rR��9�8��k ���Ƨ�����C\yo��gl�w�1O:�������-=�D;�j�Zo��q��dP풌G��Q�0��|�ʶ=�VI	Wy��w�]Q8}ew�E��ǒ���:���mu�x�0]>^`�Y�3~';��`~�S��&�j�Wf�<�z�� )�Ч�]�c}�8�gU�;9�46�W~;�6uŚ���1�mA:���@��V���l�g��AD*���9���� $�<w=s7�^7��Y��[��i��7��(���ii�g�Y�Sl�^�vd�r���^�컾Zb.v^����O�ڟE�ˡ2*c�є�.(��y��Z��6®u�U�a�U���G�Vqs�]����N��xأd�l�@Θ���^��nz��zG^���U��Y.�
��؜�}]�g]!��1���	IԶ�������Z-�b�����B�Z7G�wn�>=�q`>�[���F�r�я2m˫�Hq-a�oFJ����#`�N�(X�$�`�/vz��\a�k}�N������ԡ�=��oאi���JM�a�h��%:l&�,{)2�h��8�4�@鴸��n�2�Q��wې2x^s�X�չ���*g�%f��$/W=aqڎ�h���~#$����E_���F$�1�l�ȣ)��x.8�`�bW�rH�;���9�MϹ�������t�{��M��و��R}!L⑐t�)gz�[�=o�b�}Y��]���o]m��<7&�ޣ��Z_�~pB.�@ـ�@�x蛈x�]d`hu�={�s���α㮛1�{6�ϻ��&�u�ު�4<�Y�@j���
�k�{�Nʷ�3c^���9��N笎�N�1��Y�zq�o�2}�}q7󩮣jd��gt�]`�(���nwN���8�{��z5��03=�G������g(��W�����~���1���c&��T1�U�h��'0��Ԃ{��	=��Z��:ؿ�uR45�G-����>j+���U'����ʾ�wqhG�rr���f�X�f�:�E|��Kח>��zU���g{�鬒���o8G�͖�.��T}3w�Da��8.]�S��\g�����Q�g�2ϼ3+'�7����E��Y��|�D����B�������?��O����t9��Ѩ<��J�sQ�|6�u�2��`����<D��I�1@{�5��>�M��g�\f�n�g?�>G��yU�˵�=q�/]�]�#�W:��X�̙s�����Z7�����\)ޡn���O]�w�Pi#��pzMe |v��Ϩ��q�2ߩ�A�j��ʉ\�\��������z��3z���t�9��uc"�}n�7���z��T��s���f��*��uŝ�>=Nxq�`N'hp���Eή��=���l�+���Xz�����p�h������3���C�uH�9���\ ^@�jt����\9du��1ꃢ=�go����gNj�|��ͭ�.Q%�-3���#Qp7j�= [!��g1�c�S\��O���z%��z�1����.��/.P$���`r�wT�S]I����4f_)(�]�x�b����#��q��t�v���㵙�<��	f� �������}�)S�����r�V�ϧ��������T�WC��9�n�g�/��t;���dʞ7�ut��z����]��s�o��e: �u��@<5{�E�mZ�yֆ�V�7���z�D�3<mP?>��dY574�[@OW
xHyP���0���a>t�=��{ç��C����|;>�/%�ʎWj�O4�����b#��r�hwŻ#x����������H�)M^e+�.l�G�9a�4��8J�h�5yR�����𵦞�M�,��~���k��[����
�p���]k�-����]M�t|�	+���dl��*u&��p4��K�=��V
^G�uٞ,������j��>b�Kfӫ�B�0�*�^�X`�|=XF����꘵2w&���	�.�@)�-�e}�t!�z����:r}��(�}��d��wLr���+�"�u`�S��
�l௥�2���p�Ѽ<7���&��r���Z}�xg��e�ΪDP��r5�< ��u(}�p��A:�za�W��]� r������}Thwԧx�l������p��SW�Zg�u�_v۩�`{�	ncv=��iU&mhsYW���4�;�l�����ӟ��1��[Lj�w��=�/�R����{����ʽ
"���<�ǥd[�Q�l��Fٍr5�I�G8��؁8�_3+�s<<�{�y���QB�{U���������tg���ע*�0�<B3�2�_�f�������w�3�q!W�r�.�.�{�2c6��a�!�>�������1{�m2�J(�.	���yLRٍɧ�}��6�޵^��g���EF.�Ǩ�ϧ����W��u��>���� �3�P2�
�����7�S;G�j�~R
huT���Y49枾=�����;o��n9�FʖnD�g�����D�J�uwQO!�H'�$f�	s�b�cWe�B���תv;~K�+iRÈW���Jed!��-�c�E��Vc��d64�3k_K�U���7{Λu
��=|�F���S�^`�2���[}�u�v��ɢIJv�u)M�%V1*�EEu��X��l��3�<��<(\K}~�O3�����H�=��>�s4���+�.�t��0!�2<"7�"�N�25���r��3���Ϩi�a8�8�fq��^��s�F�-ԗ��y:�F�E��P6_Ya��ۇ�/��|�ѓ3[}�ne�i����ř٥�㾯s�#��\g��K
Ijt�6`.�*�^��p{�Vd=�9�M^�n�{t�p���e�,�ǧ8��q�������U]F�L�Ս�.w�i��+�Ĝ��8��No{Ƽ|�|�Q�m]ыM��9����5��h�,�\�;=o�;z��/מ�}��W$GO�S�zu�Nv�u8迷v�Ek����l!6_d4 g9�ҴLZ�;�/0��V��]g+���hT�ƃ�G���[���>�ߥ3��Q�U������0����vW��17������E� ���h�za�VWx���%��N�[�$��U
ƙ��Ʈ�_l��qno�{�\+r;w</��Mc9D]� .6ngţ�K4�_F��W��?SLj��oLT4<�����wc�r�����W���� �%�����CA��J\Z�<��s�ͭ=�w����`&����PFg�����33�>\׾���L�02�=h.�.��if5
�2n��3&o�{�=-��<�z:/�/i�䇽a�{�>�j}dٷ3�j:r6��E� I�˂9y�Յ�Q�²{���ోk8��'z��1�t�wS�kKQ�R�,fO�ts5���-"���ml6/���L�WH�����X���^����ϣ�������|��h���u�3��Nt�X1�<e�S<��9:�Q����W	�.�����ls.�!�����è��G˩�T_mOӄ�Qc`���g����TN%]�oH�;R/��J�͞wW���a�����qN�t:���g$�� ���X�QӺh#8w���t�79�����ELt,�H8��G�j}ţ�r<v����U��N	�nE�L�����WJ���S; �V>�>�m��j	ݜ�:K�l�A���>��wI��;}w|h9��|��n(��^r�q(��:l,�뷾��\�&�W���¥��}l1��Y�zoI��,G����4�]|���p�B�~�������{���R��2����ث����H���i/!�`yLX�#�Z���kZ��j�ֶ��յ�m�Vֵ���[Z���������:�����j�ֶ��j�ֶ��j�ֶ��[j���Zն�֭�km�Vֵ��[Z���յ�m��Vֵ��������*�ֶ��յ�m�⭭km�=[Z���Vֵ����d�Mf���V~�Ad����v@�����[y�#��U"�}i
��I�Y����i�dm[F�E6kZ(E6ƅP*I%*��D�CϽ �x��&ҭ����lֆ���m����� km�������f�Zm0fX��V$R��[DW��acT��QJ������kCj���jflm)k�m�4$i����5���em���M�lT���IZ����V�$*�n�n:��ۍ���uw ���v9�p֭���V�u��=�i����f�O x(^��(��5��:  ��� �7�  o^�z   �p  ��AS�^���d����FS��WEdz4��4��0)Nf��:�F���U�v�-�7Nv�m�����*�[c^�f��w��՞cm��;�Mfn�f�����V�S�����;']��@�9��U*3`h���f�*��8��F�&���m��(�1�(<ⱘ,��(�n�uQmmh�ei����k���s��U��ۗu�RtێݧAݹ�mUʮ�9�9uQ���kk�q����< 䫶�[�˸Cf��s���U�C��]*���i�Z�ݷYUU;�ƕ����n��K��sn���#����h�i��mM-clk�  �w�uZ\�n�ۮ�Z��]�˪�*���"��Xl��lٻ��;k��7]�5G%۩�MkJ����[;�f��ULL�O  y�jCZ3V���F�̠u[�.�m�#��u��1��i�G�ЪӪ*�ۺ���p��ܮ��X�eVm�g� '�Q�z�t������Q���+wp�csp �ں ��t��[�7��wN�[l� ٞ =�
tk��
�5��Aβ�)�`4#H�u�i��j�����R��@TJ00�H�� h     ��0�I$@ h��  �Odɤ�QF0&L ��&`M��@�(� �2 �M4@4�RB�4���PО��Ci���f��y�) h����6F!=MOS� ���duvWq�ū�׾2��m�cL��z��MzU��*�Y�L�-X�"DF��\E��BDGc�RX��" �ATD�'��,�"2H�td�|���~v������*($S�@QL 6	�>�4�R
*#:Gg�>�te��O�}����z�	��i�����Υ�s�e���4��S�[=Q�Z)*��WV�y튫�N3Vyn����W��=�[[EZ�ӌʁ��u�wZ�ljɳ�,z�-�*�koI�[��[�x*Ah��I��͠.;ѱ��n,�jP[1��/En`��e����Y�hh-j���Z�P�8ň���;�f9Lܪ8)@�nb��YBa���է6�����Ð��֘�޷��P��r��Ir^��͸`�s3Qr���U��p5�>����`[y�`��2/ �aqɶ��Xi�m;:�QB�ݣZ@SK���in�r�7R)��̈́�o�&�0����f������Hk��{���v��tn`�Lf��n�OEa�hPXM�섖U�"���ܹGT��,ˍ[ƤU(�d���a�vy�
׻J���n��;T.�sd���	��s`��ŭ�9+/�X+Id�*m��ȑJ�J�a��⧲Un�T��I2��v�F
�yZ� 3-��te�5-TW-���VjiLl��hے[.�Q����+5S�c*���u���F�),�n��;1�Q;e_ڡ�	X��C)Ix�;"��R��>����S[�l�/f6��yFT$S#D��P;�U�]n�@V�z���uJ�<��Ҋ����wI�;u��.2��j�4$ӗ*�zn����G�6�o[�%�,���t{7	XQ��  �{z�C
脌z�KvwU[;35n�ckl�q3��Y:��j�zd�u�fU�DQ�ue�T�6c��g]��N��#Kt��Y�����"�S���V�P%���j�槍����N`9�6��F�1�e�PS��Um����N���M* �����2�m	�TP8YR�dʫ����i̘F�d&��;q�ʊ��AE:z�2O���z	*��藘p+f�W�+ S �cP�y{�d�K%X/3(A&R�U�Xh[�y�=r�ƚ�y��هD��L�X�N���d3dC"7��é*�)��k�%��R��X�X��T�O�8�9tod֫q<qm=�Q�"86*k"-X���`�f�̹�nc	<��K�V��`�R�"��V�ɮ1��Ìf�a�ѠI�tԲ�5-�ݶ6�aKF��*c���e�ÙӔ*�wz�V"6���xK��(6�ZLh�J�YN#U1�Le��dt)KE���X��TÇsc��~Ǹ��zeaaa�{��ui��2���R�Z��fZ�0fi�Z$y'�X�5��WD��*�[�<�T��mfdj̿���R2���go-=5��YV���FG�B��G-�x�j�7k{:��^KZ�G%єn�xv�2-҆d��8N��w�ݘ�M��eixCq+��2�J�<�Xi�'YѴɛh4�q��qn���NL�Y2>N��}�f����_�p���
��Y�8�fY��+��*�aux�F��F�K�"�+Z��!�Cړ��e\0�t;y���e=�v��-G�|��z�Q�7Es*�4�}��
���}Vj+�קb$9��r{�4hi�-�3�A�y�J���7���ն��u�/����� �B�*�"��'~E6teՓ��m��y�߳�)+W!;�2�A	�[���13�u����)O�Q��ʟ)��%����KD�(�G�*�6^a�pK9k���J�HmR	;�V�f��R�oIT,;r��H"q�r�j�8v�J쓲�[1��($�qF�Gn�ɭP<�������p��}� 8��a�Y���TZ���r?�G���F��Hm�0P(5�$�6-�Cqͥz��DT$N"�]�D���j���P�x��W#��Tu1fE�,CIUy��)�'n�HS3{Kh��F��*�&�F��u-*?PGآ�a����%�U�^�4��Ԁ�f�]��6�����Ϳ�1Ŵu9�M^��{��6����d���M�����aԙ�Mf��L��4]�ԍ�¶��{��X�W��0�ʐLOj�5I3r��w�n��H�Fh'5�D���&�h�I;���F��n�c�۸���Fi�g2�hiK(�RPi�%�͢ńoeC�gm���d�o�f����b�t�I_@ղi�[v�iJ���YSImVZ�"�O��y��՚�Ǻ������� ��>��p��h��nU�*M�Kє~��*._��Stޣ��)Z)����)�d��Uj6~�l%Z��%cߋ���Y�(�U�9{[�,�^�6��{x�Kn�*b4�.�xZ�����ZY��b��<�=�p�$�W!ES-[�kor�l�RX��@&�uWv�UcX�d�R˼:ԃa��5\��Xg�������e\l]�h9��
e�,n��չ�N�a�lc��k�y�m&����4+b�x�"  e���TJ����Uf՟�]b���d��%ራ ����YӳE��X*mx�?]��ѵ�ى�Hk��5��W��J4�i:E�Ť�����f����13�Z�kv�ʦt�*��E�Ч��e���ff�x)��m��h7��V�-קXq��rdGU���',F�R���Õ��������.�m�ȍ����J�R`���0S��E�1�Z�baL��Ht�ە<.A���%5V#j�
�,��+D��ܧ3miC.���IV��LV�q�Ǝ�p�rX��G B��ŷ�˲v�����.��W�ދ+�Si�!��w=6VT�q r�t\��#�9v���[1Ӻ�XV�K�Ð�Y9|75.B�C���M���/����)��:Ѫ(�YS���Xב��0�(fFZ J���xjG��A2��65���M���U�U���J4񳮋���ET�u�h_���qU-�Z�]����ܝ���Ǔ)I�f�ɇa`Q���rXeBj�v�Un�ɅeDJ�%%'	���XE��¬�r�&k�7�ㆉ�Y�ǰ��{wj�K��f9�-��V-�h�R�uD�8Û��n�aѸ\�	Xm-d#�г�0�0sI=��K�+)̷Ec//Vō��"��n��u,)y${�k��a�[x�ʔl`.C�RI[!��舵U��K�Ȋ?Zѣ���̪�$s^I!��-n��k[wEVCvH�]S�T̙vi��uY�c7O��'���x�9y�c��0��F��I�d7��@D��;P�̱r��tl�ѕ�U�v*�@�J����o��TeW���lʎ�� �+~jc�B�Qk�/U$�WI�Gl�4���F�ՅU�T �G&���Z���bZZM�e�ܓvu���Hᰁ7�:ʵm������W���H��f�:�*n��ʍaNA��5�(4��������PU�d4�̹�D�8�Ѳ�#�C*�������giSN�&�:v� l�Y+kj+Qڢ��F]K��'����)@�r�Ѻ���el�4N�l�)ֆ�
��͝�F����#��*ݢ�,fC*�ie�A�!B�F�I���,�&L̑Cs\ܗ��V�E^�VI/C�Bz�͵�Ee��Z.Ҵ!��d�1	+u�G&�PP�mD��e�5m��iTuD�Yܭ��M$�#���=T�ڼ7��0&���I��S*���Y[zN�*�LX�B�7�F�,ݵ��5���p�fc���֫�R�op:�����f��#ot�)�zm�1k1���ۅU�X��c4J	
�,en��j �-U��y{��S)E�[K2�Y��1�
଱����)h��e*��Ū���� ًi�kyrP�^�o]�o�b�#G6D�Q6��hdY|��t��*V��`��PU�m�v+�q�2�xovG��5����T�U��je,��p��<n�
��`�G7E��)�TNn�fVe٢�7Xޡ/(�H�R��R3%��,��e�fn����؛:�}�K4��aV��e�"b�kE��l�a�a34K�Z��� ��`�Y��l��<��q=Б%<Ҁ����;鴖_A-�72��Gf+�i�Pk��K)ה���b/�e�W�K�i�Q3�(�*�V=6w�k�pՇH��f㙊J@[�m-�#uDl2����)��ב���7\,fe�f�^ҧ�	B���T�̈́2�W����G$n)�b��K7�y�i<wt�K�֋�^���mLQe=��4%�#Xa[�Z�6[���z��s�������U`���3.�L͂3H��A�U���iV��Y)����}\� ώԕ�3s��6Q`ڛs#2`0,��Z�-�������'� �5m�d{7NӒ,�9*"sAMV�1��U&�sV�f�S4��k�ݳt��Mj��Fg�\�4M7U��ip��ji�GU��r�F��ïtX`�r�b�Gtki������YX��)�T��j���.��u4Ȟh�����{�B�tM#��ҍn"�.ۙ)���-B��cU����j[�KJ��F�56�����=���dP-��c�X"�q�Zi���$���̒7�aқ�ˉ�k�]�Ɍ])��%z�4@/uŊ-�ǩ��x��fp��������b3�6�)����T�n��x��a$m�J�1c��f���T9�J��衏2��Y��Ϣ?2��r����c4���f\�x�M*�����HNmv\��<u�^u�'gI� �П���'�G�����N�3��A�����_�h�������#����8���eD݅�v��RI%$�I$�I$�I$��ܛ$)"L�$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�II$����S�I�uw��Mm��J`�YJ�r�.��L��E��)��]Ka���7;��5����˩X��������*��
���ˈ����U6��R�fK*�\��Zj���`�t2��s4q�2�B_E��8b���Tǆn��7^�Y��ץK���\���Dm��}n.��ov��Fig3+����f�@&5���-�)�A��5��EfC���NU@�={6�+�;5�R:�0@�[wu3L]m����?8����Yrw�ʷ���/�S8�]�����{|m��sf�%��YOV��x��Kp;$���K	�N�c�9g+]����lm<g[��
��Q|�{�]��u9bZ���*mV��ڮ��@����D$W3��m�Q��yk4	�v �*�F҆�t�=o��:[��B4�$���w}:�i���y�o��Puҭ�T-<SU��~wR` �F�V3,X��#��$v��d(�%�s�����vK��h��0*���
VC���͛W�0Օ����`�)ٸ��o�!���	,ӇX�ZQ���[��%c��¥�&�,���Fu�B�Z��Ef�&�ߓ\)���̉��ޒc9��]�*����Kg����J�^��D�K�@{1+����z�.�R�»���G�G���Xew�,���B��FV�R��j�gv��:��vt��So���(\�A����X�҄��T��-�jPQ��꫙�+��ul!(�D�����3-�k2S�;��̠v�T̂J��d�I�е+SQvbؖ��e�A�QN>�E��J�vv�;���&gq�E����}m\=C��֮N2��.K{r�BZ<�<.^V��.�F	Z�N�v�Y�Mp����j�Wn����Q�X�K�����kr*�Q�d<
�o���yթ�!S�f!kX�ǩ��1ɱ�l�e����Nۡ͝��++�B4��lᵶ�]�gxp=Ac�����V�۫�b�JY�S���}4�f�WZ�,�p�.�����P�\��3QܺN���P�E[�ټ�OpZ���9�Ѻ8�֎��|����je�ۏ���H-��{,ʳSviE6��4GX8��v�G���֎���Wa���y�仸rGʲ�=Z�eݮ]�޽F^��Sh��7Ov�i�SEȻ#�sY��)ض�`;HT��u�^0���i�m�2H��ν�Hء7K�b�����
5w_1�s%e=���e�F}r���rK�V��k�6*�I�9���4N��l��+�2B�ghMW��^jF�*X;m�d5oRv�F�����9\)]ɫ��3��$k��c9�gh;��C�ײ�E��]Io&p����O{Y=�ظ�Wi�o�&,;�/�;NnvlB7�}eE+Mȴ�I�E�jE+� nm`�q=j^�$�u�!�����M�P�yz,�������z˰p ~<��Üf�.9�`�FT8���Ѩ�`]�N���o�.�-��8��8���CVT�g���.�dmKܯ�\\G�ՒlԊ���^�UG�E�T��WA���ZN�ѓ }WG��i�U=��7�%Dqw���
qՇ���V��;j�F�,²�x�	
ΩYf��YZ��g�k�j�R�}[��:�&�#>��'�z����{7V0F��r6Ô7r�8P�s�i���d̾{;�w��k�F�os�8�k�
�Z[6���Q�LjD���l1���wX��k�{6V�8����Q3g�t�,-+����ǙiIyO*t���v�>%.Bghj7Z��������[w*v���v��xӌ������Z�qvt�yL���%��*q��{*v�S��i�y@����\�Swe�)u\p�9���"�V�wJ�]\ۂ�L��f��7�V3�I��=�Ӝ�֞�x4]�p&����v�KX��N��3��<�i��z���U4� �Y�0���FAY�)٥	E�Nd���orŵ�� �}�F��e��.�I9u�I�EO��Q�H4Lŕ�v�Ӷi)İ���+��Ѵ��g��g$�a0��YJ,W,\h�2��v��#,^�N��P�З�nQ��=�T������`�!X�MIw�L�.�il���g���M
y,�pZ����w��!���7�z�E�Z�d:/\�ye�R�`�d&�a���m����f�vs2��Hd�K g\�K7:�N'��M69��ق��P4F�D��
��O�"��vc��g����5�ٺ3�.H�%��t.M�W(Ù�ȋ�s)�=��]�$�vQ�?,GuhWˣ��G³:V����1XU�Co,:77��Y̳��ؠm�zQ}HG0
���䍗r�c�gh���0.²<��2k=݅�u�L�6{�L����efy8���L�7bM�k��	kӻ�^F�F�R�җ>����G1$��oTb�v �#p��Řn�L扎�3.p�	w��*eۢQ���U3����|c�8=��V�Ìn}ȣ� mM��EٜFܘ�	��[\'hQQk�c��Y�f�;���Qe��a��VZ�o89OWI4K�k�4�Sp
�r�eR��}c�^��k{�=a"K��M�5q��ZVN)�'�z%��GEN��*��qݜ.��Rq�v*D0V�ɛGm����Ғ9��zQX�sT�+���k(Y;�uwG���;_K	1�,J�Z�F�GO�L��}p���l���@�J_	�eK�7��Y[���10�v�_7��K�R�\���A�E��qpR�Nn}����Q�@��Ckn�&���d���p$-.�C�GtfA��Z�!Q6�˓��c�^��۪*Ȟ0��$n��I��ݸ��Z�Z�����E��7�^�Bc���7��ۥH�����.Wi�b�WCt�mr�\�yo��ꆎ7��A��$���\��T��LL̬�l����������7���3�o�UCF�X���[!�,[������ڇ�%���RA52��wY Ȇw��m2�nG��:�.��w0�V�bR���pZl�����Fo�`���Z*�O�ڙq�.�+�����խ�9��C��u3]E��O���Q_���6<���띮�F�<H��(�UE\��,�2u�^�[X9
u��@�N�瞎���^�3U�wBwUz��nU����b�(�ٓ4�7�uz����c��裚5GM'}���/2M'���[;@{N��Rr��VA®S���m��w���ZB�T;qV���B��sI]Y�j�Ҫ��7N�����
IN[�vbVT�+��Y�R�FVE�`��W��;eS�����D|M�������[}�٥:�o�b�rz&˸o�'^/���{��X�s`�rvV�5�s�%�+Y���]�G,�/{���6���-�x�vu�;jΨio��y&���%���۽�G	C���y	�{k�Nu��K׈Mc�κL/�u��kt�h�pԼV�;����B9�;,/��sk�j��vUs9�㮾Z4���%�o�H�MT�7�O~���Y�kZ�4�2�oR]�S��($��!���K9U�q��p"�z�(�H���]u|�&����8��&��bo7�x♡�!mlN� �21����7K3�&b��mH���bU�h*.8
�^�tk�6:�]�z���"`׃�kd�
c�T�����uf��᧛k.pmv�ɔ�*���5=���y�uAO!,ڼЩ/:�t0�oHB�y�V���şc�¿j7re�餶�ˢ��M�4�W��a4�G^��&�r]�ĺ�ؕԥ�KcF�!�ޣӕY�V�4Qjf"��s!:f�M�39IE�e�RNY5m;0�5})`l���p�u0Db��T�hun�&���(���g�i3�������J�h|�{Uܓ-R2�Μ������u�k�+:��Z�j{&JS�z�v%{+�������__S�H�n�B��R�� ๼:7Ԟ�drJ��!ͬ���n���טB�%�P�R�X.��EZnH���b^V����XkY��Q;zݝ�R 
ʬj�M3V����ob�t�wLIN��|,l/2:2h�v9E�|�v[㫶h���{K{+sz�G�")w*Tf�#N����T������s#��5��zy$��*e�#�9a�8-C������*���T�@�G��ݹ�
fq�od���U�l�:5ip��X�Y&�ױ-r�sV���䷢���3ː�W%��d�7F�Yv��w�<c^�hvf�����b�;���r�v�:�%�J��c��K%�g��֠�G�h�kv`=�J�|�Q�|Ep�i}g��7,��Ħ��Kd��+f����U��֎}��C�9�u����\1qIms�79M=�-���R;7� �br����1�kp�J��ؠ�2�\'���Obͧ&���72U�G��z3]V��{e8	Ju
��9�:v��S67$d�$I$�I$�I$�I$�I$�I$�JI$�I$�I$�I$��rT*K��JC*n�*+�w��
�.��9��J7i�!���$�I$�I$�I$�I$�$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$BR�wB��l�%\Y�uw>�����Z�Qھ!�_�i$���?��������W��;���?����&�	s��TQ?>�Ш��>��FO��Q�c����矫�\��>�����o0�2e�U��k�2�Ɋ^%�{2�E�B���2�(e<����c*�IQ���u�L\��JY�ӈk518́%B�Dz�kάN@Bʨ��A��VkM��z.�m*��uڨ7�ѐ�Wvo�hP0.2$U\uo!�uMB���b�<7Z	����u
�NP쀽�4ُr��/kֲ��58��l�n�4�<$�®�+�5�M]$���M,�/7N[)h1_5�5<I�9ٱ�E�C6*�a�ș}iξ��Z�Ɇ��ZƲ�\"�R�&2�Ó��n��^��k�vT�z�^VI���\]j�zbz+�Q�$�2�{�R^6D6Z��:���ݛ��������'J��rw�Bt)֬��q�߱%��f^���>�MY|-iY3���Fdμy�v����M�6O�-�xl�rH㰲�T����V��b�M_a�H�
�Fnշ/��4�-n���;*#�Wv�㳶�����
N�E:�o,�E�f��%��wx"hiײ��r���UP������<k�R���rܮ[u�K.���Y1!�{]%S������2��1�5��1r�:�Kdhde�c[C��仫��A�B��.�><"�f�[D��Y�!@�ίy`c�3wM�(�V���(�f��g@�ϞD��˸4U]\w	��F�u��r{e)��P|��#=���Qut2C��4)Iwh0���	����o�]�(~]['5�w�F��Q��)��գ��
��@�
&VՔ�&���]Y�-P�G��"�D��Y�{{'aڽ����9�v2���s{ gSF�͢짖F���v*NL�2��[�9�Jj��9X�2��{SJ���
��Q�\d�@J�{�2M�4��ʄ�4��Q�R7�Jx�[ʏY����?m�L_-��H��Cq�*���\�>7]�s�;�{1b�G�`	f�6tT�x���TO]ֳf��T��CV��蛲Z��n�|�N�K���5ЭZ�����XP���@�-�j��_];��	I��ˬ����M�7ʢTu��+73u	n���j����x�Oܗf�ȗ�E��8�C�Β���Bd��`$��A�*�i�>���:�t+g۹ٔ |Vj%[xk0�գ��9�bh�!����iv���W7o����e�w/��Zb-�u���u�ծ3��0�	P]��<��n����̟e;�^J[����񣇲Q�k�^�&���I�F	����-�1+���ϳ(Rh�P�p�=�S]�!�@n
���������,r#����v:�WQ�|m6�>1`�N�gZ�D������8;�_Uj�˨n��K��.d�1DUPWV��X
��I.��/(��;Z���]�yJ!k��4�?��D�$)n���ԥZ��Af)i;P��J��\i��u��)!������L�n��0�p!�3�w���j�i���e�rd�sK��+
Z˒J�ާ�0�kkw2�s����Lڷ�$�dw��ԌgջW|�l8�˪�ݘ�q�j�ec!$��I�^ƩT-��u;�ɝ<Q���}Hh�a�>�
.�!�����rWF�M�\V�X�b�!���p�E+'�l��V�-+���Z��b�+���
�z�.���e\���uZ�H<�4P��Ǒ��uw"���c�2cJp:i��P����=��G2M&���f���h�0�����8RzZ���Y�{;br�7��	��TS@�c�ۋU*32�E;d<c5P�\Äf�U*���l�hu����wEWٵ�:�4�2�s%(4B��f;=\f�&3;��(��I�]��&�4S�o6
�, (l�)ѵv;�7]eZ��ݲgh�jE\^���t=���@<P2'�&��)m����Z�}���udi+9�l�ӻ�#���c��0��l���b�d��l�6�*�Z@�{u4�]�h-V}đ��6�լf�����f��4F��!�e٥�n��P��R8�%Y�q�e��r�� ��]�Sͣ���!��^�V�aΒ!drOv��ї�m+Jb�ֱ�-_��Ui5�e���P�n���f�J�D�������im��� T�����$�X�
�+�M��w-̽��q��|	�;e�OT}��u�Z4U�&��W<G	�0]+ v�"\�����T�mދՊ��C6��9��6j3|`��`�[I̺1�ց���K�v*̬�~W�\c�rqs=>�lh5��&�;����,�ۊ��h7��`gGe���C;T8ѫC���iq5L3�����ꗃM�J�.�]l����dZr����i��YZ)q��_Nc3�+��<ꀭ�e]G�{���@�3�ob�����5�!��P	��V�MbK;��֗n��ˊ�]R�o����a�R�����h=9�ض���(�,\sU���}��j�4t��`�S[�E5S��4O���W�U.�"3�����e:���;w�X۸�B��&�'�E�@]=
3�M_PXP�j[�dk<�˙_V�v�2kJ�v,X���q��k���e��Al;;/h�U'�=5��N���(�M�:SŸ����Uؙ������Q�YV¯��}��'��$�n����GT�|��+n�l���~�-WR �5o�ܸ��K>�.����]��f�wR�v�jf����(�����C&e��p���ͥJ"(v��7�L�A��n�����x9�w4-'��yZˠ�48���P�Tx���Mws��<��s1�풣ţM%t�&t6c%���lu��O��(�s�g���]z�ݰ��J�
쨥W8%e\Cx�^��|�}л�]���=Λ�3J��a����Z�s�����g�`b�Xi��rwS��@�;U|^�UU�˙a.���Qѝ��S�F:�8��!�.�NC+����$�_Vj=��wS��{�
g���h�Q�6b�cRz�Lc�֕7lP�y-�G�Ns�~�	�[��7�1�S�R��Y�z�k�
Lr�?�Cm֫�J�֘��Y�2�M.�I'�j���
��ݒ�2��]�C	U���YJ֠���q�h8��G�ݱ��gGk4�n��YV`�u�>X�Tfb�,M]�3/���/�Sj͓�L�V]�8�k��8��>�Rɭnnrۗz��D�����`�ld�@�`��J�%!�	Jmw[�5���7��G�-Lh�,�鄒�ԩ����k0�gw}�ޗ��2�e]e�d^/3���(v�T�{�n��]�<�*�%p�RW����E�9Rڋ!���r�Q�Rdz/�Z�{V;9%�%K����k*�_��8��MG]u�졶՝�$|:@��m�da=�H[�!�ݢVrCC�L%/��vۼ������e"ws����\��Cf���O%L�m�K3�'�������X����S��jO��ҭY\�n��_̊�:*��SR�WCPW:�2l�UٙM�����۾�Iג�V\���i�#�#���E;xN�hDfКm�s�]≯U�V��+8�\kz�-���{$#eY.*U#�|����p*��F��JT|�ɣ���Ē����Q��6��/��V	���CX���^�qc��
z��r��^a �H�v�誺�+!��v�cކ,�X\j�5`���=�]F�UK.��F]1S�3䃀	m@�]�5r4렳H�ѱ��F�`��U�$��U��p�E.PĞS9.K3>Qm7}�`�S�K���d<��2a�� ����i<?#���]�I@�����k�Y�nWP����fY���"�\��e�b�R�>��)�ewcWzgL�wjq#{��nR��Zv慑��ʰ�`�1�w/T4H�ιDÜ�[ut�2�r�V��*�7b�V�v�Z���a��4�=�På��5bڐ���9����P�ɭ������1	����+6�'�M�`i�����R��Z�9cpwG�5͖X�mwG�b�k;�wMd�̘���v��;;�R#iCs/,J4�������e���_+�ZŴ��"u��{�Y���	V��7n�0�M�� Xg7ܩ�2�����э�����gY�R�GD7�t��٢٭U[x���7jʹ�m;{����-��1�K/]3�[ӵ�51m8��&��Wm6��ۑ����9�Y���ej&�"�\��`��D��g"_L[K�F�M��&�%Y����碍�WO�l+��8,Iw����А1�UϺ91B�-��̸&%G/i�U�v���Aul��d����όS���x�j:�������*vZ_.��ʧ��q�F�Y��k�۱v�0���Nu��uS�6,�:')���5o-��;�(�>kr�6b#h0� �ap�N�Vm��i=�=�WV+�: ĸ�E�Z�Н�hs�vu`�:���S.���[W��'�k�zbe��"�U�����
g3��mV� �˱A�T���CZ��i��X٣S���*Q,Ӹ�!K�C�jeZ�곴ݫ���maԢ�����b�3Ag����cSZi5��.����4oۥ>޸�v��pKvZ��eN4z�� s�yr��6%l�_�$����K�9[u'XO�mkӰ�Dҭ����P�@�'�\}�s��hI�ʱ���uL�o�`������DH"���C`�B$�����>�C����x�����=���{��$�I$�I$�I$��7ٻ�3��ne���ݾ,֑ХO(QA��͒��TZ���0����OzIVBVN���0���a���P7(7�oR$^���B�*Kp 9d���u�f�c�_4}�<r��*�,Q��:�"m)m�&T�즷�3�r���\��:X9SRJ��=��ܠ�C���mf����{,uM���4��5�e.��G�/����һ��]uZ;	�
��Z�y����}���v��L2&'^Py�`��j�v�ޒ���J�(Pb�q>�W��ѽ���z� �y�R���}ϵ5�[E��+��f��@�{�_w-dJ�M�٢��zn��#�j��&���V�$��-��/�V��R��R�:Î4�e��Ya����cLnoaqDovnU>�Z�Ͳ����m�vBQ��E-#r����\�����R71v�q�>���"o-�����i)s��䓷��o{�������{��ʜ��(*��9��	H�e����
JJ��)�b�p��(hK��9Pp�%
H�B-	ԙR���AԀ�Z���PsjZV������
ZZ��rd*�ŉh��}��Q@P0d�PI�%PD�%�C%h��5d�M-%�y�����#5w|&���s���I
��hu�$<+��	��p�[R
[˙�i	�������ғ���_W���|����N�{e���Z�;�\R~=�׹�G��.⊺J�D���7�����1�ߎ�4���?X�Î�45����k�s-a��zw޾�e��r�-��Ԟ�=ZL���}�Sw�]�G,v���3r�ᙯ����,֝�S��)�RgFo�:up����V_v��O-h4�K�%�P�+�RrpE�Z��S�}�%����D���?uu�|���}�":ֽ��&�o4�;r3�uw�Z��貒��=8n�����˱ŗܩ��ew��ƣ8�p��Kr/���7N3r�5�����>�!q8+�0�1��J�r۬]ƞ�N �ؔ�(N}�H������;(�fÑU��}��gJ�Jq6)��9����V�Kcm�q-�/��He`�[��N�9��3����#���)��.���ڌ}j:7�@�JnX�TQ��kN 4���N7]��4�zߺB3;�*;4/I-�Q~-����z���R:{�*�X�����wq fI#��<[v�쪌
p�ʣ�����~�:a�w�����Xs�t�]�5���Q$��h�����;�N�Z�WT�7VS񉡅2��ºU�
D.vb-�8�a���_Z�����M��7k9��_�.5��󒻥Q*�����]�e̸��>h5���`��(���J���tn����%utt�JM�w<�	���t�s�w����Vkw�io1��ewn<3�ԕ��}I��}|3
���ү��7vd̤��.H�itr'{��w2����Z�ًk	�rr��]��#)ĮձsZ
7��~n��G�v2�����	����^�N��{YQ�i�uw�"s5��t3���7�C�&���z:N��֡���=��d|Sj2'�S�^�/t]G~8M\�^����k�s!��H/�A��˃U�f\<�D����S����m>Y��0
o"D�ml-6w[��9�uJGJo0�\�'�L���t�e�Pl�eɂ6x�Pŉ!��:����(�Km2۸�"���f�"�ܑ�%��41��
³=��®ح��j�;]b@�y�eflT�fcns=)�q�q#�y��L{�pp���tYa��*/,�/\"V�ѮE��wT�+;��^�	9�^�jIt�˞��ܼX<2��+�s��7\4-9��\Jwݘ��RN���v`��7� q��5O��ޥ|�$�@���GF્����x0�ց���^��X�R�m0�A�T㸺T�Ť����ˊ��g��c�� Τ�Z���i�h(��K峫`��g7b流�����;a��IlP՜w�+��a��g:lUv9�����(�1���mͦ��-���d��U�]���@���P�߸�y��D��މ�щ�N���y�-E7݂��|H�+9_a-�Ğ�Y
N�(��m�o��v|D���3�yd��^ZW)��6�^����Dm2��}0��5}�.���n�	0��+=�W\�[k�ܸ�t�/�ěͼu�Qg!S���D��H�U�V�/��]�o�xz��̧f��d��H���$�D���q��jc!
�V���Qَ8���	a�Aޝ�\R�/����S	���0�ګ���q� X��#�M����F|\e�7;11��P��Er��{��[ͬ�|�\`�����A�7�wu`$ܽ��~r�]W��M����|�$�@�"��Fϵ�8��<GOmz���x����r����Ƨ�N�a��5F�,G\��	Ff�c��3������z0 K�=����A^�=:��G6�2�'��[(�����T��k�ٍqUـ��w�_1������fs��ޞ��K0��>��LJ��0���Io�=Q�z�nS�Ǭ��I��Qmf�e�jU�7k��ͽ���5�c.S&L�7�$.G2���QV=��2P�ԅ���]�-�GG����#�/r:���p��`�N�gRy���gH�֥��yPWs�V���w� �-Z�d�g"փu���Ef�D��S\�CQ�w��r[��Z���E�e�\���WB'U����#Q�q}#�M�����dG=�w�ӗU�_U�S�֬���\�,�X�+��4�zM�LuK�F�)3ӼH�)0������5uƜ
C��r��$��L3p�HY-MA੾}wjs7ӛ����S�I,ЗM¡${9�K�ȣ\�V�ķ64dA�WJ{ۍp���1u*>��e�=9�2����=�n5S�^W����3�3CLDPh�ZNrTz�-5,$�Wn��uref�w��$���ķ���ή�f$��b��23�7��Tre?}*~�([�qնV�]�c�د�$Ә��"�S%F�"�Pw����={�v�6�>�S-O����7`ҡq ��u�yQ������XCa:�{�C���*�@���Q��Ο�O���9����������z`�C�F��cƎ�3=+�x5���8�`�Umj"M���tG@�F	@��竢�|z�S�T�=.���-�����>~��	a=Ŭ���Lh����Z��cq�˾��KؖSi�B����W�rb��7X�d��m��}�gOx�֌����>����,:B���b��x�R犼���?/��?kի݅ə<}�э��,�,��[���$�V=[8q��9Ǫe<���愫��Q��g�z�Ng:w��w:�+�Q�J��+d��$mg������*�����P^��kSt*�Cљ�1'������r�e�)�F�q�Y|1&�UME�Bl�Z�Dۂ�\�v��3=$=�u{�)yn�Y���D�=o2b2�U�?��~�s=C���C�H�Ix-[ '�	Y*l�Ec�1��v��5����� ��0����^Us��U�C*��b�o"�wQ�:����`:�)9km;��CB�>-�O�X�:ߟ���WM&r���Q��f�`����N�����2z�l����F�5�k�>�J�c�o	d���0*Q�ۥ���ɫ�,豌��yJ,��'��뮰����e�R��M!K3z"���E���{���*�~�,L��29����J�i�n!Y\R�5�|���vXO�M�&����y�K�L�-�+��
�;*��mħqƽ{j�SoF�I����6�&7�縙)g-9O�zx�ku:��p�9�R��C�t�Yq� V��<�PE� [��x7�p�Moc9��-�aI��n��o�%ɫ��˃�~�	�{Uy�9 �׽W;�u6�34+�R���.�%劲&�;���Ȫ�ݭ�3�y�^�JϷ�OF� z��R�\%�DiiM;��>U��yxe��*���e��K��n�ڶܖFsvxHk����dxy�Q�ټռ��u�ȸ�7�oF��B��K�A��/&I�d�U���t�`�ߺ�9�ս6ђ��}ܶ��{��E	�ܰޞ��u�$)��{:��u
pAt���D4X�\�Y�Vv9�C�s����!̂ĝ#MJ��N��'��{d?c?.�}h���ؖ�	�)�:��T��c�
�����\s��!�u���w�����ʘ�p�N���`��Gu~�ܷ�/����'0�Y��Bp ���B��xL�uޫ y�>�$���2_?L�p�HW����[5=Ǭ�@�N�">(�c�3�`{CL������-�z5��i����~�rV5���j[����(����X�b��0q3��/��Qќo��l'������:��c�]��tDl����L�&	#;S�<[�p���_g=�v'�/��@U�G�'�}�����\��5�<s�w=��q�٧H��k������qgE��jj�M��ֺ��hj�]eݮ����
u��VE��s5p�i���kc3�ɼ��;M_i��`y���g`�<���N7[I���T�Fٮ�]W�bW��4U\����(Qy��2'�v�}�E��Y��\J��ٌX%����8�Lp�@%��X�æM.K
��:Vf��n�t!]�:��t���#0��4���59֢F]n�'^&�-����r>(%��E`��ӹ�ӗ�%�a�|k���������ϘL �� s���Y�y�<�5��{a����CpM���u5.�VĈ���-����4��zW'�*�`�y�j���M㺗j�ʺ�'`��CR���-�p[g��7������ꕒ_n��q�#���={6
 ]�b��bͲֵY��al�tg7+���^��f�:u��[{�>�0k7�ٻ�A�^�JN&-���kt�i�X8 ���GK���<wk:�Ul��EI�y�S�������˓ͤ\»�ض�2αwѽ�[��1m�3AQ�o���i	B���I$�I$�I$�I$�I#vN�e����Q�cd�2��2�#Ӷ[B��y{ri6ˬ΋q�4ރ�fv��fMgf��~��y�q��e����B1Whܖseb�Dv��d;X�ML`��`�4Ԯ�#��Q嶡��*�r���wY�,��ͧ�8���C^�ӛ�1�J$D7�]�;�3���b����۸^
�'fk=�]ɝKz�Y��=Q��sgj<F�8YU��R��.��C�ŹԵYu�l�}��k�F�D�9V���uj܋u�{�]儣Af(q��H4�'�)wM彭�-�{�g��Օ׺��;��''f�-Gq���2�{���Vˊ�'z�K7��Yf�q���s���VͪGZ���v����Y��eC��9դ�;���P��Q��}9=�:���'R7q��Tj#�f̃���PM�f���]j]�2r�r����`�X���i2J�!Rw�v�M�{���7�~o{ߧ���QO2H�Q@�B�P��%'2?C̯�MR4!E	@uS�BJ)E �%��!�дQJPdjA�GP�#��@�% d�N�"�B��F g*bI��NHqș!�f!u�jJ]HP�34Js!�G�$���̤h
V�3 �0�̂�]��g�c�5����ٛL����U�}������	�i�$�"(VW@���K�u���M�}p�/��SyR�g!�������Q��i<ԯ�/�y|~��.5e}K$����g�D�+�'���#���������
���:����l�ˢ�~?H@�}]$�}�藍%�j�n�zy̧��
�G2��q3A�9���ҵ�\����i_&����f�%Ԩ�H�A�ZŒ�oI�G�a'QR��݉��n�B�A�����XDc�&�i��φ|�#MF9�[�]@����ݨ��+tu[�������L�����NX\>�kj!�m�b��0s}x'�ogqFuı��+~"M�0b���+sW����p_��gEFz�+X�H8��ӛ݆\7V�Z{�I:"��ą�:&U���f��ʭ
�^&��*-R�.+�6Lm��7�/���l�7��SX�y�݅��e�����X�91Y���m���{oQ�~X�[�XJ>�ñ�c/�n��Uk�+��4h����oI%�^��]�:�z}	�Gze�dI�.��9rlg��a;">��q�7�V��_dYv��㋢�2�]��Q_vF��՘ȾcG�=(���g`��E����&I{-�WH�ߓ�$F5e��$����t}���ˑr����ܱ�$=�hL������k%��'t�}k����s�w���n!�x>��[z��Fnn4[s��K�(<���.�%pJ���z���!k[����˞���muK]� �4���6�`8ͦ� kq�����X�(�o^J;k׮�<$�=�s��o ��L[���N֢4 y߀F��bJ�9��mAk�s�m�S��k������Jr�iI"=��y֛�ڬ��Ұ�v�|��%p
�6�'75�h�3-Ge��yg+N��3�Tm	���{��|�[�d����ذ�1e�� �ت]�g�"�2�QFJQ��`��G6�����V��pc)/Zpu��h�AZP��;*��m�S�<��KܨYWF�a��j��i##t��dAKqi���xǦ��b>׾���QB���|V(Km3�o[��(�\�]ʛ�r⪤��y��
EI�^Q��:�������Ѵ���6�G_9���>�����{r^�/��{��]}��{��2�#����{/��� џ}�>�s���@���837+�>�x�O-<bn'$>��]��xq�~����+�z��=:��wyj��1Rr����$1�ٱ�b��E��)��(�4s/�Og��|�;�����Ϭ͝4�4�p�˵���'a��gL���x�M1�I!�|����^w�}����9�o`O��C��=f�}����^�}�w)ɘ4�rh�pw!���Ry>Ò�Z��5�g\��~}���ܧǘK�]A�!�5�H�]G��}������C����2����J�9�3�^]{�]o���G��'�����8��}b�˹|�üC���wyv���>��5#���^�B��ҳފ��:�r+���?z���p�/Q�	��`yd����'r�)��>�}W�u�C�>c��y��q��p{��_s����y�8��;����WP|��xT��{C��rG�|�tb;��8��! ����w+�����pf�����Z�g�]�����}��)������k7&������n��3r�/�'��i���$���r�S����{�]��={�|����FJs!�Jy?�e�2Wrs�{���q�vkr�/qΰ�{�suc���~W^��s�;��>C��S��\����9��M�q�	�
!(w/>}�0'>�.�}�ޖ�r�O`77S޻�}��u�k�>��;���N%:�p<���!�q������er5�Ț�!�B��0�t���.�97և.�x�����Ƶ���}��Cũ
M��~|�<���O;���MJyps���q�s:{��
��;�p�C�|��}�|壌���5�>˫�u���
�9�f)���V��fR� �oB;eй�ҡ:l�����v��~�rз��	Aw�"Q\�$�:޸�H°˓M�gI��D�ꪫ�����}�7߽��k���7�v�}��ش=[��0C��x��d�����>�����bjW��=��]y��壛G�{��{��>;��|����_����!��Z�J��w!O���GҦ�ރ�M���q�;����<��{��{�[��N�C��_n�wK��K컀�o������nZ�:8�9�$83:���� ܯ`}^�ֳ�|�޾�q���|w�I��<��ܜ�c�~���C�y���|���H�	��@��:�ӕ}��sr����&��[�ܒ��d�=��>;��>K�:�ܻ��p��P��ww�=o�����6�߸G�JZS�:��;�8������:��
:�7kR��k�{������u�ܧ��&Ü<��^��=�H��}/�b{+���}�m��u�����w����2Srq�/r�>G'؞G`}/�2���~��O`>���w������?]k��z�w�}���K�C�8��	�?y���^`���>�}���]�2w�R��)�<��ΰM��gîK�y�w���Ƥw����@/>�{+�ߺ��ɒ�w�{��2G�|�$��Ru\�u��u���u�s����{!�|��!N�,=����J}>Jne�=�<���
�3�2_$83�|��0�2�s������b�����dM��f����n�Y�ڂ�<�ѩ��k�%ۭfE�i�8��S`_�~��!��7N��ɷ�IC�;��X����V��9�v��K����g�N���H��#ވ�Dy���߾�߽�P����'����XF��]��N@�IA�M��0p��B�����x4���q�w��_\gzg�s���{���_%�2���y���^�e9����9�"Vs����ܔ��	C�|<�O�]q-vZ�:�����~�OL{�~�z�wP�<]F�~�������N/d
N��w+�����I�
Nw}ϝ���㮾���(}����
��Η.ez<š��C���C�z����MGQ���S%7�:�=���~�<�������������zu!JnI�}�r��w��r���\��;�-7RfuGp�H��O�b������{��wߟG����5�?a��FJq�C�~��r˹{7���|��j����B���J����������|�n!=����>���~��15h����G���p�wG��=\{��C�i'R�N�;��}=޼׾y�>����ԁOϘ�u�n!p{�r��>���W�7��۩�=���}����ןiS��������{�{�_��>O�`���a�.��u�^��܅!�=��I̧����X���7/����n��z���5���|�w�������S���䮼�=��
=�=����^�by/q�?b����Jn]��}�9����JU���̣m�M�}}�~j�ݵv�n���Y9y��rH�ȑ�K͕z3�#ັ���ޯ#����n=�L����F�y�[�U
븫ivE��&5 �\�bi��/ڪ��몯���]�߿}���na{� 7/2y+�~^��
�o��O!�1`�B���_b� �`}/w�����`�{��1M`�߸����C�G�Bzc�3�1$}�=�{�%��&�|֔�{�pd���<��_!�u�&�}�s���޺㟽���z=K��'ـ�n��X����3��%�>���� 5/�{���
d�)y<�7'r��F����zo�y��מ}���GRo1]���n^�8��>���:�*w��}���`>A�r�y�!H��{�?{��־����\��7��Ò�/��G�|�q��/qԞB��������`���^�,5"nJa=���w��ᾮoc���y�~}��w�o��x<ť���`��>\G'	�s��w]b�@�n' �� �W]a�M�Z��ﷇ>u߽�������t|�#�&��5+�?g�p�+�/�Z_.`2�x��Jy!��/�����<s��k�9���Mq�7�~}.�r>�e<��x������_=�@/��:�}�7�K�'����ԩְ�>��u�=����q�w�������|����:��|�;�d)O>ǈ}�q�nW�{��J�]󋐾�{����B��������5ߙ���w������y#��wB�up�����o�P�u�;��4y�{.�a���ٿ��p�'}h{��Mk��?w����S-m�D�(QT�R�,q]g+�a84��Fd�i�`mT܎�	��=Ɯ������=��;���c���P2�AW*���lg��uwi
5�}�;��/Ջ
�l1�{���� "Р��|����~�
a}���:����ԧ���Jw�#ܞI�+��u���G���]���>���Ύ=����~�w�s�_u�>�|�r?u���̧Q�'y���{��>����܅9�{��8;���<�e��G�z�L�y��[����t|s/�/r�!�y�~<�S��n2�8�)��!@��t�1au�'�����%�29z�d���>��s�}�^k�=��]J�'�xw/�=[��o%�_ ����>�s���@;�=��37+�>�N0Sˉ7!Hs�Y���3/z˿��w���y.�g�x��A�����G��y#�Y�_e���^�}�w)�`ҝɬ�7rf+ԞO?j�]�������=�G�^o�b}/Ҝy����ۨ;�7�uw#�uC��/��>G��u�쁮w�
d��)ܞf��Yw��׼﮾�7�����~����`��n_z�(=�r�'�x��A��;��8�/�����#�������q�q��w�oϷ�|�@�-_o���z��'}�_h�A��Q}]5�n���0O
�=q�k��t����e'�i����YN��_���V��R��Ŗ�)�3��S�Z�v'��Ei1){{5�.W��譬��/��"tsy�${�{_*t�G�q��e��b4�.a[{Z$���i�q�}�.m���{�y�}��:��2�h#ލ����/�@t(\8l��tnB��an\[�����q�v�y[�ɳI��1��0 ���B�ddwN�ڑyEuk��c.�1\q�N�w���UC�9<$4��׀7�4�gG�(��k^WIW�9�kf�zI[=$zx��Y���`y^�M,!� ��B<ߤ��u�}=SН �]~ ��X�B"�a��d�rYOȽ@�^;#��^VN�r�Y��T��5Po�C���_g��F�g�V�E�@`	=�-X�a�n!>��������Ufb�2Y$4c����3��S�S�IFe���d��ػ�~������n��b��r��+�ш f-�'��������{���9���;��TytCy����2�"��s!lpb�'7�;�cn���BK�c{"k�� ������4
���R�H% �J�@R�P�5H]w�~tSsH�
{�{�0����$�Ƀ�tfA���)]D�=an!��"�0��I�g>�|8b:�����8_��˪�����+��Y��I��r�^p��EOn���-��_��B�;����he��bu�aV���H"!ЀfoE<}���relX~��)���jex�#�0����%m�N�߁�C`�ۡ�F���Wc�3��:�yI���Ojw��_*��#UN3�Nbf���92ژ��-������X�yS�Q����Xp�+1��\_�	��"CXp��vu1��쪯ʊ�ߛ�p
Z`�Ҵ36�	��n��pj�ܶ�::�ջ�G-#xF�iR4��4L\YY��cMS��� N�Bo��U+�f������I2�fnb��\�srVK�b6�9"�-���t��E݂l�#�ɑ��٦�Yd�� nK��%�ef�\��uwq���v���`�F���ي"U��o�T$׃f�/�f��#�,�-`]�H���\��.�l�d�sm�9e���
�x�q�R�oovf��6��eE�o��g���+$g���u*nH ,��Wn�6�cN����,7F< �I�uo�9�a��p��k;X����W�5eU��!�{�į(Q�ݞt��,x03����(�殃]�>|7E��WA��4ڝv�v�mP7������[Pǳ�@7G���)7���8�w���ܬ�V�^՗ s{�j^�r�#w�����nlM�dkCW�o����o%X��<I^�һâ��S��u���Q�L�Z/Y��ՕS8�� �l�M�8��	���m��I$�II$�I$�I$�2�>���=3B�p+ʰD�בt��_+G1�U�s��ƆV��ߒ��U����	��a�O8J��ϳ:�(��75��IEY�s�������)���դ۾�=��=adEXj�TY{|�����D�udH�X~S�ŽA��v��P9�`��3�����+h��ݒu	��u�;�VEC�Q���e�%��y��h�fR��h#qj��]�����nS�
Zl�<Ҏ�NޗYL����-�E��^�޸�ժ�[�c���_z{�M��T>5d<��ϖsө�Ff�}�o_`��_ �\*F����L)oX�oum@0X[jm�y��q��q�vm'�;]ܬ辫�O��L�sGB߮�!ܙG!����fF��D�պD�S���"�ܱ���Z�q�j�������v��ʩ�{kAYt�mv &1s��\Ӫ�͓����٥u;��źF�&ܣ*N%)$���$�I#3��{������)C@QC��ʔ�	�u%T��$ru�CP���As�<ږ����R�FB~!2R�a�.p˩�h.�G�O0�����̜C��9�cS���:��8����#��D�G%)a;�DCHq�:� (��u�?��M^�kyٝkTү��-�X�m�;R�Fe���=�Ҵ#�jM��J�Vι"G�}�}UU�x�M?���G����a=������>cT\<�~����%�\(|������@�ƴ"�կs8෪�o�W��8g"P4��j�7ȡI){=����\Ӣ��;�%���-<>�rG]>v�!�1c0�V-me�r!��n���UA+n�|�������]�iul^�s`��WI�����_��:M�Z�qtwA���J�SgӅ�����]����Z>Md���?yj}~�M��qݓ�
ޚ��lpe*0��D�:�=z�9�L����A���e�����~��O(��ˡ���e��k�34��N�|;
/��,f�"���p՚�ts-l�۸3W��]t���7�D�������T�>B`Ǆ��-p.�w�:ف��X1l���h�i��4�����DDFbn�)@�uY��z��܋-�f1�H��-��ҘP�Jgb�Sh�������G������Ǽ�B�i�ʷ�l=z%�g��Y������,F�W��)a0[8�B���:��]���fξ��k]��z@`�۳1$KF�5ǹ�\�ڇ_!��*�Rma���CL)w´�q:|�����ZOrȲg��+j�Ez�	@�Z��W�2��5������S�Ȕ�ٰa��qt�F����~�D��G��>4��\�����ڢ�ڬ�k��2�E��&�4�^�7""v�h��3�N��N��s�&.����n��M�V����x�<�+P6�o嘧��9zF����V�~<;u{k������&ޑj�b,�:��?#��z#�u�lL���Lr��{�(���	VS&lWE��X ��^͏Lp�
�ɼ�~O;"�G4�37-�Y����y3yI�2�}��V�QU�a�jzj'� ԁq����n����N���[A������u�-�VUG��R�[m�8_��ck�vx�V���K0 �VF�9��0���P������p2���]���
��VQ5Wʚ��Q�q)5�����2ּ�.��tV&��+��� F��wƢ.��k8��[Uc��+�+�ouX��*z�㖺��c�=]�y�j��G햤6�{���si�ِ.�y�o��#��a����y�bN�^�9��u�uwrT���[�ͱζf苝�v�u�8�Y/9�]M��*.bI?������^�Z-�t`����0ZO��c/+"uUE�;��,|��t8�L2�y�)����nLk��5��ۨ�3Ѥ�7�������؜�:�.����R6��Z!���8��&�^U��w�'����1�ػ�O2H|�\aw���r��z��KR�*������<c)9�
u��9t��U�1E(aeM�\PL��T��r����һ����g��[�&䄾jMH���{![sB	�\�ة���ʭ�h����K��w��S4c�0��Z7�^^�_U�&35�s�[2_�3��-�}���`�*��#1掮�-�qb��KF�_)1�Iݹ(���U���M���K`�e,*�fb6��姎�MC�G�"#Gcm��?AWz�{�J��7z*��N_cm����>��1�Q~0��rs`Ft����z��˾�X��[��ַ�8����*�c6�_)�롧�N�ޒ3MC���&�Zp��v�=������Y[.�)%�����@tSj�����FA��,�:�Y��ܨ�*/���=�VsZ4R�Ξ�St��<ʝ��h�7��Py�Ub�Ю�&^�w^�Ɠuz&��H����C���۾�n�T��9��9��#�;���\"�(G.a���sKETR��ho�&�]D��˽7�����#���L��Os��	s�n^,��w���`��1aC��:Dy�*<�r˱*��T\��Pd�gI�~I��x;eb���ύ�F%��o��Ԋ6�z΄������.��Zo#l�`g�3���5S�"T�׳�t�u-�a3�GI}�^��t5�R�[3�z�m,���PT��4,��7�z���s蝘n�\�pE_�-2#�>�ˡ��]a�xfL�:����ss���3>�W6���e�3ϑ��^9�j��\&�+j,�	M�;:�(���5�0,�)��tc�P�1Nќ�UP�;*W�{�/@Ɗ{N�D���k{�{K�Qͩ����5stws	U�p�S�f�+gN��z�7��֜A��٧�f�I2��S\�ޥ^���g�V>,o��Z��"����Gh�+-�����f�J�x�f+��h�F��klXW�����:J�ot�<�jS$	��┏�]--�mnT*Q�`ݪ�u׀앆�&��P����}Q�CY曘����!��Q�&�ێ[�E���\76u�Nb��z�〽O f[=<�d�s�V]�������w��&����J�+>��[f'"R�c�"�q�F^��Ưx�[�;�B�`i��Z�,�7=S=��J#h�c+��U�^�B6O9�o�.�zxpȨu��>�OF�]
��[��dZ��#p���e �w�g����~�`4�Ġ5�ҷN�W*$�3�C���¡�כ��*��^�ŒL"�
�F��M��l�𦞁�"��3n3�8M�0 ��.��+�@��|��3ݖ�v��\�����������gn�|�yO7���bث+s�}Na�ʘ�����*^
���%��ܻ�'`g�%RWV�J �����>`�m����RNm:d�e孎3^�P�G��Z����i(L�+!l�͆������B���Xf�cSp��|�YZk�5�wT��8.?/wgZj͠�殝��Is_?T�;G��&�_��Dh-�L���|.�=�`�I�z��W�����K�K��Ѽ
/��g�}� F�B&�H������!��l_X�:M�}p/^��ꩊ����.z�Sn���e�� n�9��&�3�b�;IkD�[�9���O^�Gzz�4Zq)�D��{mkQ"�
�M��*/���pV�j_&������
�ܮ�^��G̫�37�%��_�^���!�W)6�xfk8.�ʊM=I�ԧ*��^>�&+f�u+����9�;j�(e&qN�mڊ��=���y�Jm;����\��r.��pJ��(�]��فܳQOg)��;z�=�����TY�z���Jq�y���b����6*ojd]g� }V�ڣ���y�]^�ĭvڢ���.���|�>p�#���Y���nE�g^^(�Lu*�z�$����m�����99�z$�[u���B�f�K��<w�R�<�_B���^�֥�
P���VL'A����Y�M^�!,��}��L{S�XS��x���Z�����fQ���eׁ��|��+��o]z�|�v�>H�����~�Ŧ]��O���3��"1��f�^f�[k�Ъ3.����G2�J��k����̗�Q^�7��`�Έ+�:QV���ƍj�C��{T�&(��7W\�E����Wh���`[�������K)�u�Lt��»،�B'��7�\�L��p[��D^�n��pm�1��'v�襢��4��MC�`�Xm��%�ٰ�a�]����&��9��*��CnD�5�	�I�r�	Q˷Y���X�W���}�)ua���}�b⛬0+$F}�ѐҰqgԗD}=�^_�	u�Fe;�7��Re�y!қ��]ù/�-�ཽ�m}ȒV���}��=#������uE��B���N1�U��o ��hz��"�z���>m�˷��HW���9�8����:�ssR���O�͍'x1Xҍn/JR���"� �([��Ȫp1�\MH�����qgLX���h���ô�X�+Ǜ�]�N
zn&[��v��)�S*BW�{�c�~ew�?#��߄q}����U�}gE�,9�oeX�V�@F��b�u���I�t�[�+#,Y{�F�B2> %���L���ݿwT'~t��W���
��1ߨ����mn���v��`6�V��̬�{�p�:�%f���K���=}R�`t�{wF�cL+ˁ���j�+�BU�]'���j��G���ʌ8_`��iW��*W�J�����^Pw�$���g$ &�%0F�#�sZ���r���@)TY�SQ=%�h��+Ov�f�5|_,�8�3���M�ֹ�*�L�[�E`wZ�MT��X#GY���=�����g1>�#������cF�Tm��4Vf]�2`����4Y���d՜y�3����ʙ�(`�"PK9��k�O>:띤����N�\��;����E�t��Rk��:���#md	#9;D�M,�l����}�]��L�#u�M�
d5�Ҙ��l��w�vD�vY7�PXM�3�gml�k	�{�ҦR�NQ�Q�o~�0Ev
Ⱥ�#��~]և��͘@���I$�I$�I$�I$�1�����+�e���	9)�xs�÷6����U�f�f:Gn%YRMy���!��]X���i���n���$��j��YQ*Sw��[Z�@#�\�v�+�I��R�6�GL�1��ӏi8�U�o"��֣��I@�}>h�Ԉu�l��K3;sm>���b�� Y�+��j��Wn��:���e���S|��Ò��/�ei�oY�wr�r_j�MN�j�
R�.�)������ϩ�;+��m�\`�=
�8u�w:���zB�*S�WQ��H��v]4�8�d��+��Yԫ~<�[��>��L��y�;G�V�v���̖�i�CC�cviI�+m>x��t��.ȠK�) d���#X��U8%s��Sq�DH\(^!�7VwSp���)��gwP"� IPp0�r*��)�'L6�Rf��h�pE˄qb<�*N%)$Y�RI$�H��I��/�3+n�"&b!�}#���)�2����u	HY����I���=hǨ9�EAL
fcA��Y��ʸ���Jb2]A�Z�$����Ƈ� ��us)Ԝ��-E�5��q��1�,�F��ֱ��	�&�g	ns�:��EEfV�([1��VAN�!(cXkXd�γ�s����i�0j�C.����Cď��:���X��f�V��fY��9,fE}'q�Z�5h)̲�� ��C�mI����Ib��:�¹��Z(���9��qݭ��}3�ؖU���兄�6I��M�P�Ј���
��.�� 0�����#)x�y�R�D`���I�4x�۳�Bb�F�o�r�y�"���o�Zw���>��)S��8s�=fն�Nnx��o����GD���w�zW�x���PT&U�t0�e��;���̇R�'�ۤ��[*_���b���K��#��%7���`L��P{(f&����}\+�b; M�1N�ny׳0zi���H��f������꥕�I�
��On:�������-���LQU�%�fpA� &�Ja�TοMi�N�_6u!�Ws�[���WCj?g��]d��]V�i���.�D���T&bU�sG���P��u��(}:;��{!���!���y�<�`$`$�k-e0Ƹ��X�s�������i��Lxb��D!��i*[0�/�+>ں��U\:�GJ¬���q����Q̓^�,/m'9�,)�r�dE�AJ��V`�sݗ�f����X�)$��G�=�m���ƌ4F�^>��<f�!�4�w�+2����5�Y�����xP�0�Z���G�<��sY6t�$��G�gq:4ܞ2�۞U�L���_�~4��\����<X(�9�v�Gw�=}�l���:�IPC<�
֒z�B�ۣ36*M���i�E��X��Ex��u|��^:r&hR�ش�z�X��wjrx�F�o��w�D!NPL_�}{t����E_o���Hh{�R^Qr��s"����H����F!\򼪎x1L^]��*��u7�9vka��վ����`�zf��C��3��V,�\
�)�z�9k>s�H*Y�w����$_�Z�k��~?Rܔt��"3�z����N��UY�M���j��V�z�ׅ=O|�!�,H)�7ω�:<PC;�D���qf�n�ۦ�EZ��`�����/t�Yx4ↁ�ǌ���FN�N�D>��dC�N���П^يb����H3n����U�T����DC�JL7Z!O�N�'<j�U	=��,�ͳpg6���D��7�Ŝ;�[�A�~�<{���&�	z��ԑ�MX���fҔb���wZ��)���VC��N�������d�++��.~ڢ���V�\�V�5����ܹaؙ������di�B^s'�N�����;���FtM9�0��Gc..oϟ���扡P�S�eg{�"!��`qZ�-x�<��Ɔ&}>�;�y�޾��r�Wt0��]�����Xo�D,��[O�5������������wHO��!0,�ׇ���R��_$V`��rw9W]��6�>�}�LvS^C���Zj��.!�ŵT��ם�����A��
=�+���5���#�F��F�Ĵ��?���]-���T2c�:Y�	,����F�qq��h�IGp�܈Zqu+	�Gw݌03p��
l�@�t���pOEB�[���fQf�[�M3shW˔Ȓ;�G�"
e��uv��*�mF�s%�|v��g��xQ�M��[ܓ���O�f{�vXp�lxj�=)�<�qiW�JWQ�2"[��e��i[t54����y�'�ʴ/�x|e�=51~[��1�/ꭙ/��V�y�݅o�NW�@� Ԋ|�ӆ��a9O�;�}Ly\��97Q��p�i���)�a}�f��<�z��&�k�]���-�o��bD��S�ڳ9���:�j�Ü�7Y�����G�ty֩����=5/jӝ֥I�nT�
	\<�r%�����ӓ��bm���|�4���ə���S#�m0=g�Z��p�B���E�%��o���{�uR��ZF�#=�%(֟O�Oc.��755n����:��nxŵ�g"I[����L�<6GLh�C��h��Z���oȪ�;g5�v�ڜ!��|�]��6�݋>�Hԗ�&R9����ǎ��+z�gk\C��$��O)fB��U����`'1� 	Դ�m�,�H����d��ƫ����{�	�jX����~<e m:�=�=�d�F�f���	^2��=q
v(9[J�h8�����;$Up{5��ۭ6�;�r����.&�K����"t����2F�9��ն�Y�\���-�.t�^�`��a;��������;�7ʈ���MU�x"|V��{��d�x���Ulo���AJ��!z��X��yK�zv�wʃ��_!rv�S��B�+ʙ��L;�+��j��]{�`���:��H�����s��L�g�o��hj�"�=58}k��;c����v�~��ʃ0����B�Mt	zj�'z�R���1\�M���Mj�q;��70���w�ݸ+l�d��s���X�50�$a��J�{ꝛ���IF�Z��������_K���]�Ɩ4J�e��u�YW<�� m1~>�K���X�L7Þ�ٱ�J�fɎ���,.&�+�䔤n�j��.-��"u���
�[�h:B��/l݄�!��)~�G��&�������wP�2�M�z��|��){r�x�	�4����f���� �}�ffC�2&g���5Q���5[⚨��|j�ݗ�޺vX��=ƐŸ��d��԰�g���ԼD'��=j_��6�Hv�)LvW�U�q��ZFح���� ����cb�\n�����Y�%s�M)���ĉR�D�ݭ=��\C�h��9 �N1�=Uٝ���5�/��x���z`��O��ͱ���	�"Ν�G�smGs3��v����w�j�����#���x�����*�m_nf��b=ﵒ!g���z��t��J֒jS|t�y���Fd̳m2��ɧ��]U�����|�t�x�NJ�A�J�^yǙ�q;0���NS�<��+�0�oT\�~\Y֙i��ViuU,.��X��ر�7��A�V	b��Smk��G:I���c��'�1�@fV��e@��X��J�1H���y����%Gmt�R��z��՜gv9#g���mo4[s��W6�̫�3�kdrG}�i��k_��d�&�� �lq���� ��U��獘g��L�|EP�g���#E\��R���ԓ˹�0��x�'�Հ^H%��^���\~�.Q�<�N�)�+6�����ن��s��9�*'#i�P{��%Κ�yB�7�j�Y�K��4<>he������ѓ���׳8ʬ���V���fe��~�;�����D�iz��6�g
��[��2�k�*`�[[&_�cf��.7�PFJ�A
�:d_)����rj��u:v��S���ܹi؜�����*��L��&s���VFE˃��Jٸ�%Ʋ�|C��"ւ>��d��E��*Lʵ��WT��3r&���mS��i�������Ϧ��W���<��<��Χ�o������Ѥ�WA��PL�}�o2݅��By	mp{`BN�M�8���D��em��o"11�m�,ęZ�@K+����=���y�#
mШ���9��1y�7� Bθ���-+<n�lIjo���s=�����\^�6ؒD�Y��������潈�/,�����`>��0.:I��8;i�!�ZGL����i�yu���e{7�;��DXQ���5��$_�vwh���f��d�,��75��>�/M� Ϡ�+�>!f�^��hk����[U�&��U߂C5A�L��}���)�>H8��Lg��}��q��n�*~t��Ipi�������s��ؗ9�+\_;.���T��h~ˠ����t���
jE>Z���Bc�Vw���U�
�Z�9�]'[�_3J�z��#O�M��;K�����I�?��U��U���������sx�-5�Տ�f�#��/��6��EƢd����v���;1�r�.��A*M�Uw���p�F��ۜ�sxh�
[�Gu)o�u6��
����M��������ݡ��܋���R<m$F�G��	0����*�4ewZ�8��U+!+��nD���Ԙא30~���}b�oh�8� �!��Ҷ_}���Y��)��i�$����h������C��2FKv֟H!�e�t�u]�ۤ���,˄n+*G"I[��|}H�#��4Ee8-:��$�������b�����H���H�����ǅ mv���iw���LOB~�2.j�-�9x,ʘ3%E��6��y���vz�CYљ͆�Y�z�SXI�q���w�&�#-��5>ݛy���]n2�FF�����X+���L��q:��3�"��,߽e��ͽm�ٌ�jd9�'z��QQ|�k��Es���R{l��#-=�<������Q�̋�TPT<k�̼`ڦ�������^Bk^���� �M=��0|��mة�e�ԝ�`����� �j���z50��P��Nރ���'Cj�r��|s�GvyvFkp�(�Gt�զcu�2[釣k��r!�ElLK�Ϊ�S5���;�^�1�q�g&�N��5i�^��IW�%7w;���!E�P�5��!񬍞*�H��x���1����C^��/���ǧL�1Gظ�|}u;o��X�9�J�Vm�8�^6�ڃ0{�f�Eu>�si�S�[�u��ħfM��U��d��#GN��Oz1�p4G�r���c7� |*��kW���=d�{�䥠.�Վ8I���ԅ��羷`�������Z�8���r��h̬�-_�V�y�O==K�Byi���u]b4s���^w|���_y�����6�`$`$��X�S��ϻ7�����P*�i��۸E�Qþ���#y t����o�f�o�¥�X������Z[�>�g���&��>�W�'�@��{Bz�vj˝jK��|7���<r!��=Oh�+�6n[�իm�]x;��
�#S&u�\eA��a���.ko��f���� �@�A=d�m����]��<Et���6j|y����C��U�d˪�u֍��g�zd%�zE\���*hU�*e�N�_p=��1�*�k!S���cc.���t��t�-m�u1�ڳ)�ɬfDK,S��ԧ���7���GkT[g tM@�)��vh��B�0�s;AC�p����@�&Q'�gu5[\���j�b��R�e�3��}��ut�N�{vD&@���n�`e��<k.�۔����^R�l�\��WHe.S���!A�]uԱ�S�y\�޾r'��7bYr��4j�ј=�Kݺ��^�]yi�\��.��r5�u�dYuu��r�U�*i�7��mT���>�4v!%^��{@�N��Y��k2��W��{�AP����Z�����U>��Yk�ˣ�,�fQ=�i�L;�or^�K��}:�S�aبEg㊼}6�I$�K��I)=$�I$����pv��s�
������!����Y�J����Ffdv/��a���yaV�i<3�]H2-=)�y*�RKybj�y��Z��k\�<-��|�f�Y���^�<;aGˍ�T��{h��]�s��&su|�m*ǀ��n5���Q�ۗ�5��tԸ��R��o	�(�W&�:��-�O�h8c��k5ԣ���5p�����������1xj�9oX�8����I��a7�+O+��"f^Y��d�[ݱ�b�_*P^NZ�)�ۭ�ƏWR�vc�Wfe�"q)ɓڄ�����I9�w����*6�䖨�iQ��v���/fVu�+n��_AD�b1�}f7&��:��&�NB��S��Y܁H� �t߉1����
�M�ڶ�w��� �H�r�
�MW[��L�PCԎ����3m�o���x��f5ɵ:ih9��Mhq�����&���O(˓�JI&�rI$�H�����L{F8�!�G�B�����Y��]s�sΠ��:�FA�U�hMO���\q`�Z�FA��&q�q���g8dZ�5����z�Xs�SAͅ��YO���*ծ3,��LT�H2���?"�),���i�ˈ
3�Eqh�l�0
i��˝5�ea��:�9'6TZ�F��38�ʆ��ʪ�ֵ��� ����5�F��"�"���#�u�(�P�fEQQU�q�k�+�LJx��q�;랎	՚�+..'TTd�fTd�&��F�Q���Ph�}��s�u�78���aE%g9����x���<׾K쩘t��ʊm�=�wݣ��n��d��X��,��4��ݠ�HZ��{��l)����컘�߷;`oZ�}1.�9�_��jqT�y��
�&۬�ƐI�g�m�o!�>8m-=%A�Z�OP*��]��W��fo���>���گ����5�����1ş5�S��=�7e�6CSf���7N'`ҝI�_ST��Uj��<��Ii�+���2�J~��[#o����o;Lu��#?.C*:�ff�o,ҷ�C]��Ik�t�W﮸�ED��
��d�r�����+#�v�n���N]P�رp�ʙ�i��29R�fԽ�>ѣf���a��]��̖x�=I��9�n��}K�g���إ��=�����#=km�i&�f�2�<>���k��4�Zt3{�+.�����[�%k�yޡ�w��$٠��1R�gL�N��?���/���92�L�̊��W��]i9�ĕ0uj����/lv�R�ҋ[1l�\�8��$�����9�j�Y��X�w#c�	(�B�������NBH�7���zO9�Fc~�nNЗ%��S�ʞ���0&�n��A��י/\ՠn��C�ok}N̡N|w�J�r�	��eNu;��^�\�R]Wo�g�Q�,d�qR\k)>#�ւ:=ό	�xP������-CbD�c�<g��8���k����g�P!ӝr�fz������C5/!��;��Ӌ�Hq�9��G�lKGɋ\n�+�=QH������+D�,^/͌��Đ�R�^���M�)�,�/0�ە�4*%�rgW��O07�;n/!����kM]I�v�˷ޯnf�C�׎W��5�P���D���#�F��F��g�k6�׻̣�i��^�jgԄ�"��q�Tt�s�s��>��F�b2�"�x\e�+����cK�b8����Z!�W�\��� E&�Y�+u[vR�Pf���z��-%[ef�W��Df���Y�݈�!�N�I�:{إQ���R�u݅�M��a���OwC��`r�c�P����_%��=��.�tE%���ʴ.;��������M�Di|����:�����;FT��KD��SR#�zf/u�I���wg�sM�!0��6_\9Zo�^�{��f�p�O!��8�ut=]������ ��fY�ԥqҧ �3ʞ�s ӘR�M��S��A�}x����L	��wps���NL��R�)p�8RUi�I��!�.�͞>�y�{JFx�8��!/;�_$��^��֏�}2��� ���W��Kd��,ʒꧼ)I��3�n�y}B����kϯv�č§.�nAI�g�D��c��Dx�N�<;M���<��'�%K�t���:x�m?l[���F��3�fk$f��hk�|r����k������VG��;B�g]	CǦ==N�b�+����o��O�QFh8���o�1e����8{���H�Ob��؋���V��ꨰ��#f�d"�}��F`1]"�ԥ�7�%5��quM޷�E'��\�/��-^l�y��|��Z�	�$�q���\^"u�6t�D���c��Ҝ���l�h��������JU�^@��+��8�5����vj7��{wsܞj>�DQ�D�<rSd*��k��E{�w����Ê����2�@ˣT�a�icnt�ԩ���UGY������RO_JP_3�fK�Xq@G�ϼ���O�{P�N��_ x����7�r%.�ڬ�D����_�9���+��,p亜硥}�����ʉMЮ��x��S��zDȈ��2<]��1jJ�/m�3Q�#�z�@����������s�%5x�U���c�NO;��xf(v�e��L'Uy��GN�>Ϗ�F6.�#�9Q�Y�d@Ѻ�B��Kxdf�0nU��p6I����;C�=�����}zM��
��*�۷
�>d��j]�֫ڞ�b>��3�׉A��� ⛕s�����E�3t�8o:�.%�ֵ��]W·h8D�Ѯ�[6|-j�un�ˮ\b��O}���E��́�_q�o��0�G��M�,=<��/��F �ճ������9�-Q�;��c�t�h��K��.�ƣF���b�{p��j�ˎv��hثsb���55&P�R�)�*�^��ۤ�M�t���P^�&�j���<E����܆�a���)�q2���M2�g�&yULm�dw�f�WC��wW<���Ր�T�w�`��0���D�o�������Z�4�U�����ލm�J�"��D���c;����ud�<�uLqA�[�]�h8��}�vQ1�{�ˈu�%Ӈ��˞Ԟ��B쮨�1[ՑJ�n��*��yO�Uggy�Lj���Qc5���4�Tr��_n^(:�����'yo=�w�Ğ�1��^�Ʊ��e��&��WҧX'�����S\ޱ<e���+f;�{D-/&���Af�XT3d���l��y%,��rn���7�6O*�	Y�RgPٸx;�ɽ2VCN�Y�SV�f�izU%}b�ޔx��C{\Jm�T#�@�˞J��xƙ�ğ�U�ϭP��>�Y�{�Y��?w�uY�Dӎ�1+>�Z�4綌����7��� �>��t{|�N՞5��w0ֱ��I���ܸ��32�A�s�����Nc��ހu[_?CZ�/�6Z^�y��D�{8���0AUFYv�7c��AO�lFy:\n�O��aa+7��ŭ�{�:y��YB�����'�/O<0���4I6y�r����-�߈C��=+'��0�"��f�Ό3}.���R��o��3�}�1��/_��9s�"�nZ{<����$�Х��w���5F�s,��3�M�7���#� �|�^�U��L�v���Fx�F<|��9�$'�R�^W���\a���I����\^	7o&���㷷Q,��TsH�3h�t��7-�I�r���y9�,FZ'P�֕V�Y��d��g=[H�$�]S�a,��tr�q]��q-�>0lg��I�J�#���;��Kh�����n]M_��j#^�0x/$�}�pO�n/!����:e�;�XԽ��E�!��הF�u|rX5�y�'Q#f��Ѩ+6���ލ��A���ʞ�������[Q����MҒkeJ
i�Y���	Uꚓ�R�L�Z�1ir�yYHi�6!Ӊ;����&/lت�������g�����0�VU[	��X|v֞���C�*��� /۰�m�LO�U9�ih��!@5"�k�ML~#7���ݽ�qa>��<�7������i�ɾ���.���L���7*�ީ��G��OM�S.1X��eqҤ�2#��6�	V��M�B�p��-��u�u�I5�Gq�R���R�5ۜ�Q�b#�ȗczF�@ǋ���;�YJLL	]S	y�"w�Y��y8�_v��G%t�ɘ����Jt�#���LZ����-����˭�+�L�y��V6[rT��Q8J�����ZWY�z>��R������FN- J�g�`P�L��� ���W.�t�d�EEK��C]����Z�DK�b��
�'�����/���c���R<I'yYԸ��+(OL�G"�����u1�j"5�5�1���3KԣXy�'��^�T�p���n��,���7�q���	sV;�S�r��_h������k��3�} �N����I��~'N����H闕KK�g��p���r�"廋�jzg����y���x�8���ǁ�>����D����D=��¼v��y��w���r�朝=~܏o��ƒ����}�k���@_h��Í{����ή�%d<Ę�ڇWZh�19)���{ϼ�k�r��q[^:@�"�,.�f�	��n\�Q�,ڸ��tr��A��PT3Ө��ck����Э�4tIOZnǠX�Ս��Ff=]���[���k�{�˺��l�
Wqd�.�d"�J��_��ِ�I���$�QJ�� ��㹇)��o^�aui(�s<4bY5��H��Ot-I���CHOra���g�aû�Q����s��}�t��<�������K��K�Q�\����+{!M�1N�ns��FT>�u����A�x|���.8b���t�DL9
�I��C���5����F�R�@LB��U��'ӄ�;�HY՗�7��!ۆh�By��v2�7<��~a�H���İ��zz�cZa^��]��
��{�^ڝ�t+�k���b�v(�B�M�Vϋ��Ϧ������q�Zo��z����8YGn.Zb]\whu^xz�1�9_�;m��V/K��A|���]���&z�tP��pY��A�o�-��wF�^�+4^V������xR���_��v}��t�������b>�HfΜ,	|�j��J ��2���;~�H�W��٭JS'����H��m��m��
�v�\��*�^��U��M�7p&�:�Vr}s+���v�p���Q�S0NҸ�}Գy~jm�ߑ�z������̸پ�3"d�k2���[�7r���%F���}�e�I>���7��b�x��\F�?5x���]qZhUj���^�=�w�����iC�3�J���/5���Ƙ5Q��m}�x���~����zV����L1�$;��Hq�EytƼl�|����*��g�驛ٻ��H4�s��������S�\�4>,e�F	��ƥz����ek�0�,�G	3�:0�g�ό��t��0R���R���;�a"�7j��B���E����$�L�D��k	7Y;�iekԂ%�1f�S�
x\a��٨7��$�$���7N�K�S�vf{��Eu)~.���)Y]*C����S��w�*`H��r�o�Vnf&gTe{R��0-Ϭ��7.X�br|�{� �R>���}�^�\m�[�P���ܷ!�q�)�e�а+�Dy����X�"(���f��7{�g=��iqʂ]��n�ͣ��VZ�>(�e�G���ב=<�
�<�j� e�&W]��嚚��a�9�����鑶�*4����.�V�K�T�Sop�ES�qc-�A��Č�!ԶA�`�!������g5ٝ�a�ޚѯq�M�&>B鑵+��H�}L�(�����Q���
�V��٬GBx�`�Z�ې�Y��	���ݽ��C�Z�3���s�Zξ�}6����6�0��	j��=�hk�6��k�2�mu^��!>�t�%�=CE�b�s�6'�;6��y@N��,�yJ�<d|�M]�ض�4�gF(�̜�X+�ax�M�r�rpu�ݱ|�Գ�dD����yt��
&+aΣҧ-���d�=2T�(��
��<�j�g,�i�����i�	�h��~�q����5�ʇ<�\�%�h�L��đ]�91i�Ԋ]�'fh�` �0�I$�I)$�I$�I$�I>�Y+��_(iSnE�.J��{cU^��f�,+�X��I�
��D�Ś����2Vy�{��/LLR�'3b�y��N�5z����Y�9`�ZM.l�z2��'�;S'-��!�����ۣ�wp;�5��Q�1��Z�iv�Yy ���}�o���!15ɾ�uxglqj�X�{fz3���N����ݰ�)!�7�8T.�_Wa5�:r�Wv�i�t�>u�Y��!L�.��b��Z&l�vjx�	�XDv�
��܊@V'Kr��9�;bRg`�e��k�Y���j9*�y��v���76�S�����,Ss%�qE�㚇�-���N���ʚÁ��uLD_�-�(�G�tZ�k�Y�L�yG��4�)���8��JpE�l�q�E��we�	->�l6"p���vP��4J�j#�H�'�D�G7"	>2�ɿ.ZVs�Z��������<�.oB��,��I7���������*��s"H�����y�d<q�9�dNNf9j28�Y��h������Y3�q�#IZ��0�s�Z���5k�x&8�Y�U765qa59ej��������5��&��d�Ffe��VX�f��S�4QITU1E͑317�QTsN��]a�Sqa����(���

j5�ucu�s�ڪI�5�0*�l�f�`j�x���7T��Le�TPq��c����<��{�}w޾�v�3x�U�-��>D�jk�F�=��١%�F���'n��Ԑ#��/�I�Y��?����G��17#F1[Nto��G�-k۪�֜���`�>�L9�1�h���#L#�0'�ڷv��z�.�<�!J͜��|�jb�I����u��>�Bf����i�|p�;q�[>{fbP݆��A��*���7qp�f�3 ��= V����~]^���W��U��^$W��
|t�<lj'����P�E�����<ؾX�cH/8J��q/T� �zQb�����5�&��n�i��������Q�<9�Zv����Ӎjg���y@|Fj&l|t�e��{��ܓ�U�����o ���RB�A�K� �7>�4� ���p��H$�6j���/�au�Ȗ�:���F�+��(���د�!����T)���Y)��ŷmV�O�|��cKD�.v�0ejό�{NX�Z�	tJ�$��EZO�,r�ZC�%� �� ��\�+�ދYr�W�C%�dݩ~�$2��<a=A�\˸,d�e|WZy�j=��ɹ���N�)wnAP+�o+�����%&�Aܘ�39�&.�8,��r�ى�/���3Y&&*h�o)׭�������sjgpZ��f^;��%Q��V�ۘ*�ܹ�̧���IM�����G�ظ�ZS᫏��3��H�[�v���嬽���Y�������0�H���;�Դb񗏎���u��y�b����y��N��P�G��e
�#�V�a4���ͽX�s~�)�cc.��75%�2�ڜ�S3%P��j^m���i�gz�5q�"_�I��g���!��f�D�/R�4%ۍ�6ƛ[u:�ʜ�ޭu����t����)]�Y[�[����������zA��K�hZ�Ma'��2���u���v��u���6͟|��/��4.�Ћ���,�	�AU�x��D]�>�I��5�y�&��פd�Tl�̾���K|�Ү��xAY܍����>�&�k�d��n�m��-��!��7\�2J��� �3.�w�+oU�Teoq�
���!y7aC�=  8���3��sq��I���\ng\v��,;�Z�!F���͛��{��#�d�~^J��oe3[m�48ט�P6��������������o,�t�'����+h��c��6���F޲�UbZ��8:��u	,�9J� �b��ڞ���x���;��ת�oo�N�<��C�|n֒�<>�̙®6s�Z��Kٽ
ΚǺk��7���x{Ŋ��"F^���05x�P��Cc�V�.ީ�kns�M�e�s�0����<l����ظ#�9Q�W]j&Hf吹��3:wYu��"�\_t�q"q�V�$���Ԇ~&��o�Pjb�.���܂��w
K�un�Wؼ�p�p���qx����ʮ��k3�k�b�ӕo��^/��A��w�5��Hx<�{�nlD�&۫���R�:�V���ak!�^]luz�<�vʾ����ͭDO'v�Qi�^m�zi����rIv�Aٯ��r�c;�/5��=�4����\��[YP�~��Zec�3��¸���ㅖ֞�6�I�)�U�� KTfۨ�����E�Z�_?���\-��G����}=�����5���Q�ZsѲ.�]�|����!�ʹ������>�:��񲎓�����t��Ҫ�N�G�s����߮� z������&�#�;�vҥډӟ.JC�x�P'�gq!*�,������nj�[�����Y]�T}灊�c)r^�:e�9���s�r�Ȧ��G�C��Qy��hi����eoHv�w7�[���+�7����~"�|~�.�cq"��L�|E:�-���b��e��sU�(mo��,��'�i��l/�S�^Hz��+^g����k�q�������ܫ5��qф�=cόc׶�U��L��kxx,a��S��H�Xn��N�IN���)"�a�P#)�K`55��.��� o*/t'��G`��"a�gF��v�Y)��7���w���zA�e��$5�$?�_}�ra�����A&�WK�a+���3=I���Ň�F2�)n;^�}����7j6^ђ���ƚ|�L�9Ȫ��}X6tV=)�P1��ʚ%�s�d��*p�v :�S����c��=e=��v�!�J�!}2dB/>�K��h�>���e9n��%Lݔ[L��ˀj#>�4~ӔB=���kB^5�qD��G�ī�A�:lI̢�,,�/����D�|F�q�!�n�i����M+@��\]d�W �7B-�%�M��GI�����Bέ�y�_e��k�mY񰐿"F��K��O�lHVV��0÷�0�y@2�i\�w�W^�<����Ef�U>:f���'���3�¼}f>X����iq�V׫ճ�D8�)<ABޔ]skI�d�>�E�]��V���^H������Ԭ6��۬��J����{s�s�[W�����{FK�4f�cP���тD������5\�:��)�"�#��q)�����{cMN�ȪS���;��Z��LW�>!f�W{m{����?w�npW��v-`4^#�9Г7���0�jX�:���!���<^>�������-K�SZ�6��K{�ȉ7�S^�Җ�ܳ�a�/��Q�ָ��{�����P-`���:���!��r�+s���m��j+�6.7�/G��\#7�c�� �g2k_�f��F9-"��e�7KO����6'"-���c��p������~Y�q8��դ0x�-�2<���U>*Tk�9
��Y;��������1G8����}�h�x�(a���RZ)�t
s[;��jgZJb�3s���e=B���ԍ�Ӧ ��;X���}�].,�y˴��:4+wBA E�t�DL����R<I&��ô����6�]��#����,��M=WP�/�aE!E:�R����Ox������}��VG>�S�.���m�GOF+H�&��D����I���.ls���SGN�!��Hoވ�A6��u;��O�*N�DX�;F<�F���A����V�@��u6�W���~Q�oO�N�Ǣ6�)��и�ǧ�cO� ���ʧ��_)�9�W��\Cڷj_a�d���	y���:w3M�}jz�o=�N�F.d���SD\��mWP���
��(0�}Р�QF粶e���]��r�wDx�!��N2��[���1�5�_H^d���^Y0��[w3~U��V�+�j6�"�V hq�1.��v�$���9;&L��ұ�m���t�U/*pVSE��PUn���d�:Oy��=�K0�f����;�j��=kz�C�5�ӕ��\�2����r�����w!� �Ӎ�&+=���o1F}�|u8���I��
��8nn7!_eL��֘Ėo*c�{'{̖� ����n����*UƦq'����{�V
WIS�
�����;��zU�0�\�jح�3r��/og!K����AKU�5wYއ��tQ1�ssq��G�8�4�1d��^�3ݩ�Sx��.|}B1�>�G�r��]x�=��5��1aV�J�S�Wz�;�32NYZp������z^�U�����a!��U��E��Ɨ�'���E��=T'*���S�'��ū�ٶm��m�(�Zr���|��sVՌCkX$e{n�]�����d��B��\;��T�E9�^�>�Sb���55&Ub0�	=8�jP,�r��h��9 �S��a��_/���^c�鹝|���)���
72�c��d��H��Ӟ��v*]�o���K��sz�Y%zTeVˈU*��s&E�+E��L�fVz7{`y�z��R%=��� b|)��;��-�^�_m%f�t�_:��N�$�fw���R�q3T������^O�����Y�Ow�ݥ�Jb^l�Ѭ�X{�.����2�r���c:ivy��M7�32;�Dw��8�u���v[��Nr�=Dz�O2��U�8�Ckxr�:�I_�}�D7���K�[_Y�����G"���:3Y,mTt���0�7$����p�N�qUŢ\p^]-�xن�i�e�Mu��M-�m�J�~�&�\�V�v�~b�˕2+�h�w/"�Wg_����r���}���[r�f�F�Vz>3W�h�j��-��m��Q������]�b�4ĭ(l�qa���J����y1n���7sh�Ld�<.3�m�f`�N��T�L�T#;5�8uQCRGO�׆��*��ǥ<<f�7b�����a��[��-X
`K�阘��]@�v��)Y��-ϮS��r�d	�)pjK���9S��O��L3}����{>30'�mjt�7�u��!:q��a������Z��0�8���jߧ#G�M��e��?�5�A]��uDn������Wٕ�u!Nݤ�@�+�k���$������x/Z4�)\{��I}�p���K ��K�Ȥ�囯k*��i
����}ڸ&[����P.U��r�Bt-�Z^���GL�y�.9�sr��MgW���^���%��Λ	Q#Kť�c'�6$��z&�Y�ʯt�����~n�qJ\h�3�*k�:�Q=�L]Y~P�|h]P��]U&s���ʃ6�"� ���F�
�zN�KbU~�{�=��#/��&c'�+��;���GF\��}*��l��ܙ~Yj^���<�q#׬ղE�^-.\�yY��]�"��E�)j�3)˪2��m-#�Th�K�Lak]��#g�͆�= ��W)��s�F^��v]lL^�\�o���,ƞ�U.G����*����O�="}X��Ov������~���kP)�����b�EA[&�5S����=������ ͛垜#X.&�^:B����K,뺱8�3��S̸o��:t�̀�K4V<5��B$�]J���D!PIG6X�n�i�\�c��]l@����M�6L�Ζ���q0*�v�:2c�ҎM"=
t��]!���~��=.Ww3���D]E�} udޫ]w�{Q�+ ���Y�( ��ӥ������ʅvk�_�^���nܭuf	��{� ���ݺD���+U�E�g��}Um�{DI�]�y������&�T�1 ��L�S{�KiJ�,��g�6��ė}ͭ<��Y�d91,�E8E�:@���/(}��MI���F�j�`�S5hΩ�`̮7g�{�R�e���������w�om5���x6b9�WAS��<�.�V��������f����{7��9����g�(iQ�䫉;/:���]�.�I�f�J�e][�.m�M��KY�ttY'sd�å�t�F��+�6���s��	/�f�K�z����*�en����C}��s+�l[��̹�}�2NYxR��t��������6�vuwl��1�$�I$�I$�I$�I$�CBw�(�+.�3���ܨq�n�l�ٙ3�4���T���ZW@�����A���wҦf�/{�."jwQ�^��������K�n�*Q�Wٯ*�*J��з��\u"�r{c	ք��GD�]�vN�Cb�6��)�o�ݡeNE��cL�3#� grOmf� ���yV�p�w���L���c�QQ��Eo]=�)BM�.�Iܧ>�$���C�ͻ+�����F46��PgV�P˻��1�J`�GB ���n�Qܼ�Q5:t�CO�~������<;��������\2��f�(I�m��9��)�GL�֖�}���J��`5{yÕ��w�8G�SW,	�LW.9x��}�u�R�K�L"Jz��\�O���5+=�S�w��G�ʁZ���9Ӳ�̑�T����]����fL��6�aYD.�J6 Ţ�Q�<��H�&��L��2��)�"�.I$�o{����7��r�x�A�64�UQjrՔVYfu��1�0�ֳQT��SV�(��Y�9�SM���QfeLEV�#ELf�TYch�j�2��H��1�Y�I�Zɪ$�����32�
����uU]Xư�F4F����s�*J*
(x��4PU:����
!�f!F�S��ՕUTLED9�Tń�,��5�2*h�)��eՑ��3QUDY9$QME�eFK��NM�d�8EQqaUZ�(�������2�5�EUUZ�}����;����ƺ�����BvR����c�f9ܦ�I�.�wң�J5���o��$�'�j�����b�.]K Q�Zj�җ��T�s���;�O#�Q�"�C|-��;�	�h�>;`���D+�N��#���qL����!�NϢ�_���P��7�8p�p�b�'�%�eg]��\��wBI"��r�*亇ГڜU32U	/!(��	,56�'�����4,yō�!���36������Wu{w��R^Nԓ�Kzx���1��Q�z{�$�v�'����G[Z����[��b��6~��$���GI�af�����;��z�Ggѳ��${��un�Yqg����]�nYƊ�X���������:�� ����=���Js�P{�Ό����[�^a]=�����j_q�[�L�${Rk��-�Fa���.�����J�%:Ѩ�uh�JzdX��G��b4㨌��rl�uZ�����|��q1�7*�؆����v"/t��m�۽�!5v���	���I >�B�YL'H��^H��,�_K�wp-Dŗiֺ�Y
��譯�^�Q��[�Ё�r�E�t�x�HV��e���yc�AP��j�쏝�}&Of�J�^,mo��W�*]�N6t����=:`�b�j�G1_y[��?>��;'�6%v�|{ؔ�j����0>W����hf��!�YMG_s�u�Hˀ-�r�hvf'�v(]H�"eR����(��̌L���NP���P�)f��W1s��M$N2��&Ώn(c��BX��	�3��p�,;+� ���QVo�*�<1���E��x;�o_ YL�7{7�����|z���NZ��@��V/mL�)�:e>���#�hD�[k����\k�}�VPMM�r�ԅ��:��t�VE	5]"X�!�M�w �P_��Z����������O�WS�#�}�����t�
�Y��2,:t�;Z���F�5K'z��u;f�ѵ\8���$� ��OLh%�R�u�#��n�}ãչ��{0,�\�e^j)- ��y��M�V	�g�C��laaf�`:E�ӝ"����֩�5#����ԋs��Cb|O��Nz���H��8m-=R%^���۝�n3P�i/e1���U�	zw|���yOW��;�A��?jϺ�Y��"f{=+�j�ߵ'�bɒ�oi5�Օ�i�5�*~�i�i�����plcMyL!s0k%��E#�c�d-��yU�)����+˭���r�m���9}�z��}Q�]%�߯���L�Lm-���@�9��R��w��V���r��2���/]��命&fs�����])Җ�c�O
smZ�W����G���:L��$�LզSI'�{2��WZkюG���cL���d��%k�yޡ�.���zL�7�V�� {D:�{��ƌ]r�5���:�U*9,��C*�KX�VV�L�ta9�MG��T����^[蕬���jp���f0(h�E���7.����ݚ�;�+kI��5�8�_�|��-&�L�́_P�UU"v݉�J���Ԭ���r�u1���+ZZjs%'��aiYa+5�@��Z���c��������ϗ��;���+/�/����|g�LT)Bjh�*e�"�w���ݽ��!��[4�.:w�{���3�
E�9�s�6�p�l&�E�q�$�h����13����K�wy��|���3�����Zy�A�ʝ~�r�,�\`�y;\n�cQ#N>H`�i!����5m�X����ӽ�&��\�R��50Xb�k�[�W,�w&�"�u�众�7��z��c��P5����!hyH�ǈ*ޔk��{q��9�˻��2}̐�l�Ѩ/�p%�o�ϝ��NVmƺ1��z� ����Eӗ��T�sM�e�	򘴹rG�¥o'�^`P���+;bR��6�'U]%I5P�\�밉��3��f-�a�ܦ\̐��ul�i Nԏe��3�w���]��rn�1��*,�����B���߽��M:�S�6.�'N%x�z�}����+2д�Ha���>2S�.�o<���(;����:`���S��;.�`}J\�ih�E��+X�^�m�#)�;��pY��Fg+���9�euÕ����،�R�u^�����8l�0�O!�_I�&�^.;�zzy�<dfr�ܕ�$^b`���]mT5NảC1x�x�-�.�����ǈ��ۻy�d���2���N�����r'܄�:�h(a�	y�*i��_j����֓S�.����p�7>]�q�Y�h�F��h�Ӧ�-"�����y����������N$2��Ƕ�9���&^��A��Fr$����=U�އ,�|ݝ��;6|}X�4,y��<�@֐u�+��;�)Q0�M�����s�R�r�<m���x�d�OWd���-VQu��K�Z��(��n&�- bΥ]J�JS�u'�B�pNy�pu�m_�o�f{$�ٲQ��R5:ᎅ�;�Uc�����v >�K�;('PN�JWb�q�s9i㤓����4���&�2g�X�j$r���ʗ8կ����ӈf={4�{�]_g��B�����1͝1c$L�7���SL�ۛT��+���_��˼�w&���eE8O�Ù52�=(�D=z��x�b!y�����7svx��"+�+�xRpݞ� ��)�nN�J���.�']A�x^��v#\'��-��<}j��y�x��ϼ��+�/�RT�jSZL��ق_��\��<X��3���Xvkf�#ַ���լ��������4���Y��N��T���Hw|�����DɉOOxVeu�ߪd����X�3��נ��,�,Ed6v����o}C�Nx|�9���aᘿRx�ET�
R')Z��pJe���G\K���i��20�Lq�U�Q2w;��U�W�T[���{zک�Y���
{V�d�JR�nC��3��OS��]�1��{���v�C�������wT|E�j-��K����GHqZ���נּ�b����$i~U.u��l^N|n��@�j�ۈ
/r]��5w�����#�7y<���ZJ��XXAa�Zz/��NP���+���8]�ʡ����ycd���
�f���B��]:�+E���iOK�+=�;��u��	\)����b\�0UTN���SB�������dLXYt1��'�DD0�6Q�!��1f�a�,��=�s�p�2��N$a���6��z��U��y/Ncł����=X���YuT���\�5{�dY+�uo"��� �0��	.�Ŝ��;b��+�N�m�ﱒ����1����}�J"���<�e�B�;5-�50y
e /�����)z��~K�ۤD�b��*Ө��s5SO�A8���*�ʜ��3���;G3\�C=�����.�����_v��,Rk>�j]�x<�%�e�ݛl����u����s0�$���s2��p�y�1�k�C���̋5�6m��qO�j�eY� }ԍם��E
=�y�O�g'��S�M�����OMWԊ[��� �렅;R���`��軿P��?9�X�������~��Y�L�����'z��Y�Kr������~2�R�`������I����@ m�Rf��]�SҲJ�z1�#�K���RӾ�A�m�Ǐ�]*t��3nO&��wwf�T".ccl�\�߹���o�Jxx��m
��Yě��r����kڴ�ʯ��H��VZVOL�^�������k�!Cy���)���)�T&����,�����`ȹ��(MA��M��"��6�7d)VG��<^,�k�e���o!��;��#L �9��XEzt��^�4p{�����E���s��Y�N��"�e�u&n&�����Of��>�]���g�5����H��i~lc�pWD�ܽ��J�ڵ�*��f�����+,+=���w4�^W#��Υ$��D�P̭�|6c�2E�@�*��uwdv�B���`��T�/�kqqn��m�&�r��҈#��KM�n��D�W֬K۷!�)q�����LkS����f�>P�?{�]�9�Za�CU+!�j��s�EP��.b����۾bX���g2D�a�n�F�����מ�_<Rf�U�P�N�Y�H���F����/��3�n$zƳV�|5u�U��[^I�f�WG�vV�$ӉX�ǭW�oL>��iz��t�l�<�em�p�*-ٓ�Ĺ�2�ÿ=��5z���=�XCG�	�iVJ�o�
>�(���LzEb�pS����euÕ��r��.V��
������.����g�N!�d������B����\���u�,|�A�na�P��C���� �qik�_�S�ﮰ�Y���)���u�S)���܉k.��A^;
x�=�n�C}e�n�񇫰���P�q�m�V��(��sO�x��<Ȯr���<)5�䩤Kw����qSM�5����k8"v'w�����I��Gv�*���3�U�y��Oeл�.�K�+e��L���G�eNx�d�n���:�;�w�!;�0N\��FY"��r�l����ޤM���ޥ[���i$�	��z})�|�xl��Վ�<�bƆ5�g���N�һ{�1��z�8z��-��6���z!�`� 6�~�ɮ�w�!ؕU
w�Td`��"�nd9���;^�7P��f�*bƝ,�]L2�0-/<���q6񜦈�n�õ=��u���:�f̾������,g0��O�P�O�h�C۬�ϬK|sOk�;w��")?D���èJTC�1z��|�+#�odf��<O��~����rN��=BeD�ӛzA�'c��d;��`�N��T�-�B��v�fo��C�����"���p׭��ú��la����y���U�tS�m���%��Z���%$]o[�p��t�JEVӒ���j@�V�"�h5���'�.%��dLN2�i�R��Ǥ�E���K�^<�:j'�ڭ�����׭�'&cv���a��BܽR�AX-���ID���NpX�P����{�܂X�)pg���T�uG�YҖ��=Γ8��]���TK�&�3��
�n��M�Ke@s���b�k�~#z��u632Q��L�F�^���d��]�Y�u�$Az�vj�A;ᆂ���ӥ5i��q���f������`G�����r�;4E�N��M|��J*t�<z�iQJ�B��)́��搱d�·[�pS��y��[��<�"E�w��W1�2ot�[��K�C�V��T٢wF�n��:������e���'B�ѧ��(��)(�a���ci �Ŷ뫨�I�}�SX���t;4���ʤl]N���hRt�M�0�hfo=��1�;B�j���b�uaP�����$�I$�I$�I$�I$�XZ�kC�����@�ټݵ�p$�ʷ�L�� ���kgO�_J�P��g>kYdU.��<y���9�eef3���%�ܚuL.%��]�OJ�JҌ�g�iDK��+F�té�p�t/5s!�k/Ma��]u���W�Ti�;4V�}���#� ���wS���I\���s��T�WnJ����]q���p��o#2������:u!�s:=���Qq�������u��u&����'{��!9p�l�!ݸi�1��t�z����,�v&����Z+e�h!�H�,[�s��/uUʸJ%�A��������QT�xYMq[dNU˶B��2*�2�.��v,�u�^��K E�)��+:3��h#u����J�:���]$�w�4O�q��{:��4����8��f�+J���R��#���}M8)�X�{�4�aU�Ǥe��S�E�d�I&����������	�����ɧQ@f�Q��U�eYaE�dSQa�k'Q�0�(�3
*"�5�\grrK2w��Dqah������QX�Y�3e�DEEd1�q�TW֜�����)� Ȃ�ԙeT�4�4�o2(��N��*.,��2�F��fAT�a�E%Mfa���e����dwdUE\�REG%��PQWQ�L�MT�RUq�UE�rZ�0�����5��Ys�Q$��\fKQskX%�AE5AM�F5-�a��cE�N��q�Y��QIE3�T�ȭA�0�(��)3�5R�\a�M��"hhh����0nl
iN3�*�Y���1ip(���f�r#VUTQPE4QW�ָ����h��3���{�k7���
�Z'¯��m�H�]�S��n���RI��F����kc�諃\+)\M�)����=&dm�[zp� ���/͚W�O�/�5Y����ipd0+n�{�g�5yx�=Kr�{�\ū�7�q���~_L�M!�ޜN$lb�.|}��fo[\ʺ�f�O�B��h�]�W��\��A"s��˩S�����0��+ܼ��1p՗�E�l�[�UY�(e{ƤF����V2��uFbXH8w�Om?D�Ӕ���������u޺���m_����Ð�+ $`$�Yk)�=%���y}0�<͵��#�N����#�0�����>���EY�zI���Y��!��n�<�{��{����V�p��y3���'5�gLt̙.�5�qr��Q<�j���m�r�>N�������{���Q��tG�c$C�����,���~�ջp��v�sUOgO���ת��w����-�}d�f�5�F!X%
�}ܲd�޵X�B�s`���mYڲ�yx��r�Y� j�ˠ#�z�ʡ�R@���M�[{k�K��5X���B 0U�F��˙�&�Y�N���unkxkz�)���k�R6׎��ᔨ�-*���?F�z�虇wZ�$ڌR�'b�쮨Q9�B��O�Zn�9>�G��������LLm��-eÜU��=᢮�s��m-�ZVx<<l/k��Q��j -�{�Ǐ�w�������������JC�QL�םh2�A�R�)��r����׵q����$�GF���d�Z��I,��-M�a�;"LH�S`lp�ծ��J��߲C7���4��P����OX�&��؆�����/S�����o$�I�2�U3Ժ��X�g
���=��`����V��������,{�8�ݐg>J�HVA�"������3�x�͔+Ƀ9S��4����;�"����OU���tjﴺ�����F�ïf�sst.����=�T\�C���}��cQ��)��4$ٔ�&�M;�]�F��e���i�3�BV+���*x�O�����7\t��L��DS�\k)=#���mF�.6w��I��5�9mQ/��oug���GǫϚ����U�������vi�%vu#G�%�$��!�b�lQ�ƂCF�F��M�d)�uY~�*�BhWIya�o�ӋM<f�T��!K��=n�R�V�ٽ������O<�ݸ��h{J�շ�_�|�����/���Yμ��{/����Q^%�d��a�5�-����߰��W[����~���/Q3���C�r��D�p�h�^��b����Ɨ�-Z���n��X�#N$�q�]KH���D��
Ԉ)�KKO2.];SY��Ju��eܐ/���z9[�*��q������K��8�9�5��]ؓ6�ur+jPB�ָ�}H�x���-a8�r��վ.s�&�ڰ�eprKIr���t��<���:�Ƞ��7n0�#�y���6�9	�}7�=Q;�M�c��ZK��~�3u1=�E�?+���=�4���q��RYW�t,P�Ǯ��K����3��
��w{�Ep�]�0���~A}��q��Z���∻%�p䢻�fg�Dõ�:k��B�A��O�����M�+�B����g�g��1�1.����.�*LgS�^��Q��CKI�z9ԗ�{�Q�|(u��F�z��Vt��@��x��2���X�NA�(ZC-Q/Ъfd��h����4����!8ݘ���i��	�qB��,�6j��K���#:���TN���
y45ͤ�M����ӧ}Ϗ�h-�d���R���݇|x��w�`��x�
8_��x��GI�H��SD]�p�,>���'E�������e�줻lmK�aV����阄2ѽ����X�{�Ͼ����YO�Z�"E�]:���/gsٸ7i^s�y7���� 5�:+I#����e��u�q�@�5�n$� Ut��V2t��A��_��ª-̂Xŷ���y�w�� ���,TyXfW� `}-s���]��wZ��z+=;��-��i��|X�ᖇ���w(���V�fK�UB��\�'�xr�B�mi����1SK3�zߌ����Ⱦ���:uh	ddT�i�����G�׊)^)��	 �=7���Xޘ��b��(&���-����e�V����Q1d��eTt�5����.���^ �G�~��j��^��������K,bDPbgdt�K��Vw��y���Ř�{ �,բ���![�4�d�z�c<�w����8p�!筜����w�߯�Y���|i}�x@�v8�'{�P�l{W%�%����s��^"�ׇ�-��W����,[�&����j֘�W=2�.�.�)�+rF�=sg<u��h������Cۇ��/E5jT�j㥳�����|fƂ�[R�U����ph���EY��������D�-��h�(j�С�ƪ4j��:���_K:u�U�ߔ�����>�F�K,�?><gڸ���:l�CmO��,H�w|�j����u���~�nr\�CO%���L:E�t磝�y�K�o^�K�o���u���h�j]��P�Y�p�ֈ�rق���������d�>0����Ut ��֒z�B����P�l,�}Өf�)�)�U{�	��h/��iMx���;����1ͿV4�9<h�W���;(gsA�U(-8�j
��7�e��D��ќ=�����M�4�U�������Nf��/דH��]7[.u�{|~�Z=�^$Y�Zt���k�����������S��^u���oxc�^�%P���7>�\.�-�ͩn�/���:jg`j��{z^�B2|�y�8�-E"�s�J����tq1��%y���9뫥�}�U;	Y��W\urVx�]J���/J]���6-�{�8�$6w^�p<i�ݺ�*]ګJz��C�D����zv~��pmM����Xt)x��e��^>5�~�`�z��r��^��V}�/%�.xv�5���c�������;#����u��[��<�yxĉ
׭E�jH᦬K�1yFJc�7{�.:iU"{�nc2p�]����v���#J�HVN����h�=k�r��*��Qob���*s�" �،�Fd!��n��>ً����o��/���P>���|"�4K����O��7ݳ}u���Q�4��R׏������/�B
��Q��>�w�ې9w�pZ��	���C�������<l$/Q#Nx�{{�`�����R\��3 j�G�+�_W�8���bkE?0��.	Y����E�N�{�|�������5u&���}�y�;�+����Mn�(�ͣJ��:��9w�j�o��=�8܍]��լ�^:����P]�#j`�$������e���)f��)k����A��'��\�Sb~7�S;�.Mk$^��۶n�b8�ӳ����:�9���2;�{u�u��T>���#N�1{�qU1�u��%f2/+ iz����D��a%���d�k짹o@O�Rl��ͦ<��4���mB�9������$N�11yr��x"��0)��	��e�a��Va1�������=��B��7v����Z�N;E���>)���\�y����[�%�"P��el
q��t2gS�*ٵ�B�������y���
�lצ�*~9��� �64��Ȟ+���ܚcBlL޹�V��2������r7{Jٷd��1d��S�P7�N�@m	y�3I�IH�ކ[�\�3]w�D���>ѤLv�����R���0WY�lF��L���&�Vd�6��n2�q\����Z�����ng��G�h�}nNs���O5��H�$��ֻ�i�+����dM�:�ۮ����z��oT�� �5w��@4�!W��r´T`ma���q��b�{h8`��<d�����b��{����U���ga�1�� �j��� �0on�z�ݾ�`C��|�
��nN~��.2W�q�kIKy���Q�1V�R�f���5�W*8G1쫛�%�/�J����ԄA1�4�з��Pbwpk�!�m��`7��g5oU�o@���Y�&��4���Fqj8�|Z/(p��:�d꺺����������DC��\I�]Jb���f���]�{4�*h�kW�k��!�:R�
�q'����%��!Q���<s�m6�����bw4�4�d�I�gv��~��)� �ם�B��&��TT�	JՌ���Qb)1�t7�Ү7v�VL^�i�6/��:®�̧�+B�|�NLs����RA�M�O4s�#���TLkb��<���lF7�SI�v8����5�Ȍ���=Pk�nM�8�ȗ1�:�K01RF�r�2��K_�y��' �Q��:L=Q�8h$�K���,Z���d��Ś�ՂWF­U� ��<�f�ʬ���L�r��5~��tfD"ژ�T�6�d����s#�N�H��Y�5��b�q��*ã'!��5+�Y-�5%7����O��5'+��;�2�n֒��h^��V�^�T��79]�ov�I�����p��bWd�]��_p���k2^@�&f��J���c8��k9Y�iM�WQ�̓�� _6I�xZ�W-h}�e��m��w��7]����)uy9f\�.:{{����������ʺ�Z,:;]Y�npt�T���Z!�he>�P��}��Ýe��5:� ��[� ���(�Z�8�V۠UܩY���̓gGYGbHO����z��We�m�mJOBd���4�6F=�V��o5����rny_%Y�g+��F�+j��{)V���}��ʐ�N�_;������y��hwg7I����Y[N�������4{au�3�J�L��c�H�����|�X����Y�Y�+v�uc��uJ��B�A��a��9s%2h�5-�]��j[���j��:+;kIZ���kmn-{�63"T�C��r����"a��V��֊��sc�ԒI$�I$�I$�I$�H�o7l<9����2��j
i�d�o5��������^vv^n�7n
Q�����RlT��5g{��z�5�� ���� ��7X�Ԏ���:�gi�牰`�*��F�����ͪ��͝ �*X�<n�ynm,cp�cg�2A�����P�3Q��N��,���<I3D��/O:Ne�P��2�� ��J�Cމ�@���v��K�9���w9��|�Qq�'����H���}�Fr�x��x�31��_(K�S�Y���^'W��{�ƻ�b�AK\|e�kor+��^�{ٶM�����L+[��쵺�ڀ��B �xq��T�Y��S�F���K\�2�ng��&6�p�7����:j:��wiv�P`���Mw|lΙ��L�dS�\ ;R��Đޭ\�ke���aU �w���'��<5�G�0�a��ۚ��S�i�l��W6ޤ"u8�NK��2�q1�'o)$�{�������|hufEBQĆFFF솊Z��)*���N%����D�KE!DE.�8�*�'$������X��.4LIKINI�b���L���H�NHP�e�Df`�UY��ԅ#�2

��),�Ժ!i"j!8�$��$(h5du��-KIAM�!�(��2��*"*J)��eMR�%T1Q�r`�x� ��%�*��ʓ�Ȣ�%�r
�*����@���0�(54�4k�5-SADP�SKIk
��h��\�q��cAIG�uΊ%��J�y��Z��x�GbTn�O��J�긕2/q����Mj�gtn�Z���C���~C�lbSd���(���zF��KA����6�18Mś@a�Hgl�1��u�p;�d�ZU����!WE�M����O�W�J�'4u�t�Գ��K:/!<�G$�vFR�ӡ�����J"��p��5ർg s�==	n_z���+ܢ)/�*�C�B�o��d5���s��Q��b<Nc��qUһZy{� ����u�֛�0���b�l)�=S�
wj�-f�$�7�z��i��9�g��I��$}�so�C�=5-���c����Pc�i�t��bhd�鸲�*�ns�I���+���"��h�hT��͎�(��b�vsf�;ծOk*�J=�*K(�hVgI�R����.5[���;�EgD��u�k��~}�̳�gߖeq�o�t�{]Q-t���0��jo�_g&�R�*Dq��=��9��Q�b_7s�^����ڨ��ˑ�=�͕�4���������.�s�!��T��p@ˊ�ܱoW�{��o���KǨb�
�OKv�ު�lc����rWoqh7O��s�蕢!�/�w'<���}�9Ճ�l*��i���i~	n-(������ap�
��.+5J�����zt
S[}K�����2�m�GyE^d��f�؎������d�˘��V������ȳ��9d~�r2���&��ה#E�7}w�D3"j�u���u�d��Q�w�Km�r�_1��L�ԛZR��]HQ݈�Ҽ���|;���Ж��wg���"z��B:)$I���@��ł7��]�zL����]�0ώJ���3�3 x��%�\��1�|����c�;܄\�~D-�w�z-D��O2J[Ǌ+��-�x���.�s��о�{2o�P|�n���Ǹp�tz�?.�;�L�k}޺ݤО4 l<�l��s��ɗ��\ĦH�MSlޡ �F@�t���ҤS(�v¨�-f�0�s�x��2��8:"i֫�{��\.zMrl�X&��`��K��C��㠵�8��RNmJ��2z>�����B�yx���J}C���ק��ju�9Sn]�laxf�l>媮!�=F-�j��t�_Vr����JƷ���6��V�zę2�F��T�S���gO4���=:«˖��^��i�,�}�BN�=|�Y��Lg�z�S�N�z�&$z�斜�j���'��g6�f�H��t7� �<[�6�Q^�W¹<���Oh��N�7=�	ɼ�|D����.��bQV����1��T�q��E��X|3J̖�S�� rc�Һ�
�r�绾,ar�Hcｧ�)=Ɓ�8k#���TƛBӽ���mTP����k���"0�8mA�%����m��@M�Ppt�O��i\�
���#���{�:^'1(��;�=�O�N�8�n�V |�����;w�% ��<�s��u,9�t�8Y|�qt���Mݤ�b7|:Q[��ٷH�ҥT
��c�f͜� ܮ��R |��&�sL�bv���ڔm�u b���S�{��I�8�pȾ��V��[7	�T�.���/� U�9=6#�_��ILO/������HcO;=�@��}y��5�Ѩr=O���՘u�x�z�J`��4��gI����눒� �c0����8�I�Ө��6�c�P�2��d�юi��x8�Md�{�7��:%&G���O��E�P�^sC�n{=[��;.�-�`��3���l�J�r�w��J��i�|�qx������������ܢZ^��!������,���}�rʎ�"����F>$9�t��<����vi�}��T�QŨ��T'���8�5���/������J`�`��mN]����x�$x�1��u^�|�M�LO=�F�Wm�w9ɧO2\�X���|���
E�T�V�+��צA(��[̖!�M�k����m�X��ш�)���SV8��	� �HJ�g���|K)Q>asȤ���_n��tD�}X(�z{�9�$�q_Thqc��U�mέu�c_��)�n�N���g�nF�F���"��g�s
e�c:B��$@��͠|�"��) �ԗ��*:����}}��ՙ��Z���##��P�6A�T+����^�xk6�f��o�^�
�	�k/[U^�J���{��%�{J�cu�邳�-v|k2>���NR>����8�-f�<8G��\�^X�����.|UN�71�8���%�)��rue���25S�"t%�O7a,]�����W�͡�DJٽ��B޻�*�ִՆuO�Z�Om3�&�6$�9|�@�	>���%�������ۃQɩ�G+�j�z�]��QQ���Szpq��}5;˲-Պ9x�er�K/;I�a��F�J�n��[ΧS�1���B������u{�"-�γ�;8n2U@T��������$uƖ9��W�O&�
�Έ3p=<8Iط'9�'��+Ӫ��H&���ɻ�J�F�7 ț��T{�谭;��[Kˉ�ZI��v��Sl���NF�@
0*�c�sҢ�X{k1��֮�4^jAdc6��΄��(���.����mj�N �}7��u���F�G�Ө���տM&�t ΍�}��n��ZS�Sٚ#�5�PV��م@ӡs�Lnp�bG�����;��M��E�n�hC̶�����j�
��`	G6���w�m��P3W��[��:�˸�2Ө���yr]�7��Č�s����H�V\8捍����@��y�����w����-�"��Q�w��X�cެށ���*{�p���6���sY�|^$��1]�=�` %��u�Vr�	����/]������h���N���'rP5�b)�q|�^�ڍ�S"B=F6MT\ٳ�:��T�,uLyR��Z�=�FAȮZUzU޶N��{�z'{-N]JJ����
�6[
r��{Lf�':+�WkKz�̇�i�񍹵��@%��TJ��)s)���h.3���P�����,���b5W���)�ꉍ6��u��mk5���jq�Cz雃�~��>��`�����[�,�����\��rZ@�~*bz3#7��üS����xf��ƶ�êZ�@���q�1���9:�y�B��㞽��bw�	��X�s��k�-VG)���P�Y���K�:�J&�(8�?w�`�z�J�A,�zu8=C6��6��z����:8o��R�E�td�E�ą���,U���7�{Ц3����D�i�oa.b�G�:��$#��}8<�q�ФM�'�SE���u��L����<��V��y=��0���}�h�ڶ� _tF�3��Oo]��p�I}m��2�n�L �=��ls.H�s^6܇1��&�Oe(8���c��9�iH�ͤ�&�*���͚�1s����#��}��XWE��s�-�<�K��T^]ˊF���p���d�l���n��au�~?Tw�L
���:b���C�qiL�X�4oSѬ�D������a���M�⋨�.	��F���w�}p�Yr!	�����Q�nH||��,Ha�lj�9�C���ߣ���}��H�Ȣ�;��.�]hm�����
��Y����nU����lWTKL���L�p�֋�PA�dOEs����c����GE]82uK��2+�i��2"W3B{�,���t#����N
{:����c�d�&�Ӽ��Cpn1����G-(Jyu�$y]|e*Z�]T[&#��o2��%	�)[Mt=��6�	k{����QsNy �Sn��Y�b�x�v�!VX��V�wgJ�����a<����k@ŔH�{n
�QG]��Z��5����!��"�ʡ�
ד�	�L�v霺��-N��xPrps5bv5�����VvTM���s�k�:c͉<� ���$��k{���/�Zݷl�n�uwͽ7�j��s���[30T��yn��V�I�&�=J�@�+�wlGO�J{�)��<E� ҫ^��mj�iF�dvU�Nz����dclM/�@�q���;�M���^�� r�%�xLT8΂�TW2++7{.�@\��]�������vxڬE��Ik+s�sn�ި�F�A�ǻ_t�v���3p�ky��Hw�耞�h�.|乽� ;y�ġ�On�}����G$�I$�I$�I$���&�e*�]�7�LrT��R���*Ӷ�z-�qM����v���*��38� `r͡#Us��ܺM�M"rc܆52Q�ݝ����4mϜ���橍���ܦ���%��*|=��\��Z�n/3��-�����q0B�\�MO��g9>Y'hh��ӂ[Gh޹z[��Gk�C$�@f*�77k�Z����p`-�X�5��L��.�9fh��v�}X��+;l*{�ێ +.os��҂��k���]��]s�±i%A���R�e!�\&=�S&���BKMJ7u����0�U�M$����mP�j����*5-�6���Hڌ�h��X��Uo�=���].��F��D��'{-��bm���������xza��T�q���{���L\���	��t�d��:�l�iJy,wS�"eu�nd��WFF�#u	��S��';��I;yI$�I$�9$�Q���h�aԧP9-E�-P4�@�9S]��P�IF�Nm5)BҔ:��g2��ՑG0�E)̮HRR�!q��#E*ѩC�CQI\�s.�,.`ʖ���(iSR�$K� y�JV�Z�\�!����'�j�hhN��eD��Ԇ�hJ )(�JbV��#*Jh�y����`)h��G�c�3�'ȝ�P���+�gl����*s���j�M�4����-u>�:kj��J�"p�����4���Lw~�r2�eۤU~#�q�Q�E緤��:�6�� ����=�.+�N�׽jX�CV��w��cb�KZ��
�Sh��!k}�Օ�
(D��..������mq��h�D3F2�����S��v�������n��.K�3�g��s<�e��ް���f	�[7��c�q�y˳�:�GWH�e{m���3���j�
��ӛ0��s�{���W��#�z�%'�A3c*5*4��V��{L��<'4�'�z� �Jk"zMa�&浤�"�q�Or�DH���i8�=�Jq\��Y��Ѩ��
@��Z�1�*64+��J���wf�ܗ*#�����
� d��2�H&��$�K[�%�#�S�/e��8�X7����)TP�!�.o�IY�F��(8\����$7������H�4^��E���d���V�3�α�0Yw��뛎��������i���1��y{vM`3c�ÆT�&󛘜�+zG�*{���APr��n9n�(p���"TԾr�R�]T�H�cL�QJ%>^$�6�Y��Z%l*�[D�E9jV�z{��� ����e����*?P�J�f�qZk{Ŏ�����ࣜ�q0jY�صl����w����pm��L�%\k�v\���A���X�U{g:��3xhNK���Qs����OnmcLk��7S�T#q������1���'��~��S�U6�����ęT��K�[o�J������ҏdT]fi:�Y�r�1�v�8�o�m�v��L�`ݠ]_.�$��"|や�όV:$d�P̞�O�ǆt�y2�/M
�}%i{.�-�Ğ����rZ��U��%��&sS<Az��)7F�������6��@u�#��s�K}��1�)9&�`�Q��8�zAm�Lt=�z���[)�΅�Z{|iLrq�B��C�)k*Ⱥ�B)r���$~��Џ8��Ym��+���1dٜ_��2߫R50���`�)��q�vT�ZBeL<$e!�k�;�W=�p�L�"qM�
�B�6��t�~�k�����n��u2���ѿ"��9A��م��O#�y-�U���9�z:�}�I�ZbXX���T9���Y����3�8�dt�{�>P�j��x]��x�#"veg#fj�Gk�Lآ����,�_�gc��G>��3V{^)�::���N|������G�Q��(n,0Q�WF!����+���O|�19����k�L���/zH�^ոZ?F�D/�tg�_\f+N��h�W�
��QmL#Cju�h��t�+�/k"���������4�Vchӻ�<U����]�e�^~4���+�!�X��dgNa�'q���ۂ�(���I�k�g��;Y��j6��	���z1��_B3�j{j�f7<:k�ޢJ	�X,�erƧ�b�)���Ĥ4GM�9R3�M��d�. ;��n1����_[�9\IӾ�=�\>��l$-�j+O��sq�c�m%�+��G��uya�1��v�rϠ��Gc��/���*�h�v�s�Fd���&]�ʬ�F�ZkM]�R�&�O�w���UA=$-��W�i%�	yE�:��%��
�=�����z��p-���Y�x�р�z�e���
l�`E��:�ѱ�ܧ�S2֖�*b�ꐤ�X2&�U��g��"q�&�nbS�E�T8o7�b9����f8�l����ٮ��fk�V�0���'�:��N��yė�k���[��F�3�o���0�S*ꯞ� �v��l�0��[�&SbM~�/G�i}�������sYi�e�Yd�͹o����Wf��m��ږS�Z�g���}+f�7���?k�1�ս@K�ԯ�
�*5�0i�֕3������uv�VF��]8�&k��E��Wc�R�U�]X"����`o):X�Kulf�e�=�Z�������m�%�	�Ţ�7�LT5%.�UgE�Q{�"�A�ਨ�W�XOrG!'�d_���;x�UkOMY�@���v#/��|�ާ�a���D��؋��&^�r
�D�gs�M�����٭� M�l9���ѣ`Д/�����Ӽ*a�lP�kֶ���p�l9�Y(�նbe����O�\z�y�p`2=�ÆEA��%k�$�����-\P|��A0*J��(�3u�x�oqHс��u򚈱;z�.�" T����=�t�הS>��-ξ�U�!%w9��Ys7�-'q�6wH��[7f��v-��v=��
>�U/�Hb�޾�wC�SJ�D�n��|S@ԛ�%ҥ��F���t���w�Nvl�í�i5�uǓ2j�2�e8������)���3r��ȋ�Ssk��@曨����zu�0��Ū�o�/-HUC �p�a�������
99�x=%�YF5�C,$"�fim��{�"ZY�m":�[�F=�1������G�0��]|�����~<Ft�j'p^��nn���Vq�[�n0^$�F�3uͦ97|9Ì�˸���U�&sS<xј�o6�i�7p"�#�Q��{i{k�T"�����0M��1��K���(������\�D�����I�XZ�Y��z�^u)k,���q��������-S�t�<�f�fS��z��y촯�"���;�W�o2����{V1R����V�vS��`ͣ�{p��O3co�v�k��n��m��}M��H�3Ÿ
��J�q|���������%n'_�7s�1�'�F������KH����6�5!�	J�[1A([�};~ҹ�CF:��b�o6{J/ +�#�y���s��Q�Vo^۵��jb��:�r��v]RWfj�i65����5$S�S"9
��	f#ӫ`���w�yG=%]�m6�t�0�]�D5	�X�jո܉���wD�ԴS����1Pm���
�2��]���)��q:yo�l�#K��-I�����N'/O�xr:�GE�>u���]��%��1�k�oQ}e�{F@���f���Ӈ7�E�*ږ�)|���H%�t9�o��C�e\���Uu�J�����г�̆N����L�[�k�y�s4��c��H+z�5��h򋫭�1L���3��n�rA�joI/�(��.��0��YU�D�u���o�u<�)���ɾܸ�Sh��To��,��N4_�-mb���U>���i�3�@����;W7�S�)������x�wa�R"��p��SQ�\L��`_uc��-g<a�QO
`� +��*L�p�x;���l�8�O�sl������v|��{��Qi��=^$������3~�ܑ��;�(��ȫ���F�)��I������;��fr�X�L�8�@�Ζ:D;�
Y�����nc��vm���P� ׯ�<��N�뮸7��S�&��*vw��M7��n��Xw�.���`�_=�i����U��1�(��3Z�Q�:�nU���mNo���ӕ���}1#5���-o�-i}�6���.����/�f3nS��{[��^K%܂o�ve��!i���ަOJ�ӷB�|5�Naτސ�,Ijgz���1�h�t�w�k�{H��Dsѽ�k�I�YL�G��P8q��{��u��b��	��P�X��l3Zj,�e � ���'�@Yp��&ސ�J��I9u1�Rl�q��VNv����J�����G�PؙS�Y�ir�Ƭ�|/����<�?�3���	���T~�2Ȫ����KDMXg��DO���0v�
"|bɒ'������֎���Bъ��㥇�,�ئ�k�.�JE TP.1E TP(Ac�5�	��=�y嫓�:��?�g�����x����S���q?�?U��DO�C_����M�������!�A�|���"4����Qy��_�F�իM,��e���x`����׿֘�A���w�o߰���损��j�yI��y%$�8"?�%�D��؉I���I�?JǡV;�O�d�#�%��m�_��q~Ӝ��n;�*�7� ���H����Dܩ��?��Щ��G�Nے����l#$V�{�d�$[��"��_5`��~��A���@]ߏ����GNj/�C��&"�����c�;�h�5"��'򿫁�WasT!��26�ҡk�2��գ����a��?%���\?C��~�y�����#��9L�M�?���?0�d���)����� ��C'�s ����W�=f7rJ��$Deޖ�����x����$r���ٰY�S��}�M����䷣�6|;�4��7ɑ?#�Ө{���9��^Ǹ���$Dt�*������J(���܇���<������Nb�~B��$��耢'���#�`���?��X�	�������<9L?#��'G�DQ��ը��}N��`���&�A1%���{��/ q�6{��u����؏�	�z������o`s��㠯����t�
"z�?y�O�#�Oا�D.������B�o��!�)<�����[7����\C�7��~s�M�Y+��V����)��G�=������u�Q��޴A"#��ߗS�߬��0��/��/�D1}���]�<��5�΃�9�v'J6������?˿D�< �t���ه�%��c��C/Xs�km�3G9x?.[|?{U�D��oe����	����1�4�승��l�TjSӡe:Mf�������a�ÿ��~����"���~�DD��_����h��	�¼g�žk�rވH��'ro�L���W�`����!�z�:C�u�N������RG�
g��G�����.�p�!4�J�