BZh91AY&SY�Վqߔpy����߰����  aR���
@ @h P   (� �U*�( ��   � �   �@ �   � zГTVRKB�$i���#�8 ��@ �	P   
�, |	y/��A��A�qC�k�]5C#@��A�&��HDa{j��R���R�[p}�]k�B�z�s��TS� <9�=Oc���:��9]QC��J��  N�t !ǥUk^f�.@�F��=�SL���
N�J8�]���@����\q{>�y���G� �)�Ƚ�#YRM�d�s|����:��` �@� �, �<z7g���h�� �����r��0h�3!�I�40 ���D�<�Gt��c�@����9��n�A�!���   � s�ZF��S���Cpe�4d;����H`+�2`���np�=��}��o��۹�֊d���!�F�4t �+� �	< B�ݹF�vz�t��;�Κ��F��y�g��` ���.΁���mף��f4���5�齌��L��                        @   �U?B4�UER��`� �L M`&a����Tщ�aC& &�bM��E!�i��F&	�����)U<��� 0  MRB4BhOI�he6���j=#&exl�*���T�J6��4��&0h47���?<�n�t�j�k�>����t�_s�Ӣz�>,6l.=\��sys�s����xla���a�K��m���~�}��oo�?/����[�x��c˥���aRa܍�lͅ�Q�����8�p�{o��m���=������۶UUTg�&���o~o��W������'��3���ן�[k^1�B"!��D�"��f�"a�(�,DDI�""	^��"mDDL(G����q""YBd����Y�/��3�BxG���DDG�0KDL��'K�:"mD�DK �K��"<��Dq>���+��E'1֝DTS(�"{�e�G����K�r""'Y�DD�""h�b%"DN"#�a�.DN��<P��b'�0�G�e�%1��)DLi���X"'��0~�̰�0�Ek�]GS�S���GO�8�")ϸ�#H�НM�sK(��iD��b�"9�Gj"0���YyF����!O���Dq�G[�Dm�Q�eaO��DF��iM*u�6�";F�~���F���}E!�����<�DS���B6��yM(𕥈����"%�D)�GQ��De�������1�Dd�8�y�G�:D� ��aC�� ��b%	�w�<'X�e�DD��<"X�����"L,DKd,��h���f��?v"&�Zb`��؉gDOv'��Ȗ"o"%�+�DDD|A���""u,D���t`���t��""'��" ���H�D�K:"��#i�DDG"#(�7���DD�	D�	x`����&�;�Dϑ:%� ��(�~DK�DDD݉
�_"%�M��""xM4��"h�C�DJ��""'*}�"`���'���"#g>��"bh��1�DDᨔ"%"""y<P��DD����0KK舖#�"'rpJ(N�""n��X�""=�DLDM=��\�""j%	�!H���~DK����?""�Ȉ��L��DL���8""a<""&�%�D���MK9W��WLOH�߱b�`���X��x�<�?v%��&�8w�bA�Oz!���8&�""u�,dDDN�A����0DNܡ�����""'숉`��P���D�JQ�ġ٢	�X�DDOvxD��y�.H%|�"7�v�A �8���)��4���y>�m�DD�+�DAUD�<$��E�<YT'
�"'L<2"&��N�DD���"9M���#��O9"^Ĳz=�aߎH�d�D��{Ӧ��pߴdO��Q�� �?"P�=��N�M-��D��"%��NI���"%�p�����+�T���9��䈝٩Û,M;&�/"">����Dv"x�A/DnX����#Ȉ�P�8_��}]9+"u(J!��_y�g�H�=G�N��!�P��""?pNx��3�"A+��E�,��%	F���<7Ǆ�N��;���.D,�*"&d:t��D�p�G숈��8?x��"vƢ'������-�*HxI�D��"Y� �j�"q�(Dj � �|�'��M<&}�ܱ:<���8M+�N�#�GӇ�'���L0�ƞ����B#S�'"""N���,Dڈ�,D~O&%�؉Bi�.DDD�iB"&dDDNg�DN""`��""��DL0�DDN3J0D�,N���4�L�)�DV���Rֵ�kZ6�cq�Mb"#h�SM���'DFMA�DL�C�DD�:�"";K���f	b#Ȉ�N�""#��8R&�&�좄Dn""#&���b"`������#�:�"pD}���H����K,B�Ǒ�?x�(y8t��VA)ex�����F�"X�=ň���BZ`�$N��؈�`�DL�P���:y��B"V�K6�'����g�=؞(L�DN�휅nM4�ȉ�2�Dv ���,�2"s�(O�L�Yb7ı؝��N�D��M�G�ߡ�8&d�0��b�j:X�<�N���	�	�(B��e"xÌ�0L��Y��iJy;�S(�)��#�DD��D�/�DDN�Ȉ"s�}Q���&O��t���r���p�'3a<i�2��p���x�Q�Θr�9��x�}��+�xԆ����}�>��"](��Gx&��0Գ��¶A��'�y:P���"<����"#s�"y!�B"#Ȝ�I�+��$7��t�Ҩ�������y�:ی"8�a_qF)�J8D�,M�ǂ�H%И'��A��x则�a��P��h�;(�:a��B#��>d ��rQcȈ�;8p�gY�G"">�^<P�b`�DDϙ��Q0D��tK4Nԡ:94J8&��x�N���bx�N	O>��(~gJ�ı�DO��Y�"&e�̐DjAD��,�������f�'�nY҇��0�䮞9"&�=�0DD�D舜:ϡ�x"X�Ĉ��%�DL0�����N��`�9D�H�9�"U��b"z�x���P���DL$DJ8,�
�1,DE�i���������$�DM:'�D�m�3DS�6�";E	��,艂&H"CDK҄DGH�"m�%�"X�Ȋ�2�4�Ȏ7��#�DD�<&rQb",�Bh��X���xJ8NĂ&?""'D~DL���%vt�D�7�u��#����Ȉ�h�n"#l#qO#�O��D�DD�Z%�B&O'��q��(���H��m�B'KD�NL,��D�c�3Dv)�S-Dq�4�DJGۭ�T�e�<ی<�!ޖ7;�K'N�"p�o��ˍ��}�i�Ѽ";S
��iza��D��%0������hj"DE3���Ty�z�B����1,��i���	�,L=�<L�͸���S�J-+>��ı.�!g�(��ģ�j��!}�J�������.DNP��K�<?\D�y0�4�����g�HA���n7!�C�N�f�=��xDJ�"i�P��:�����m{�>�
����d�8'D�:P��"qO؜,��I>~�{(�,E�ha��#�(D�2�w!e��P�b�8Y�a��y4}J,~D��������tN�q(蜩@��%����O	���"X�9S���M(~g�,J/"�;ř�DD��D��d,F�&��B�F�'L�N�J �"'Kϑ4�2H'$�����"��:�!:Q4�޹�YT����e����7��G�}�p��D����_�����׶-z�j�����x�s����o=�os��i�-{2���W�s��	{�b���%���	oK
������^�2���V>���~~=9��t��2=�f�q��Np�6}�6; CHg$�ؽ�E�����Sf�}��M򧏛��byK�Ȝ�X>o��fC���ڏZ~�uz�a�}
�����}쳏��rs�heO�=H���w,��	�=^��l8��wg��(3�{�gL�{˚�%��Å_v!��9h�q[¬���$���<o���r��3���[l����3i�|;�+���pZ�%�{���ި���ug���\,������i�ù'sT�mԱbײ̻�����N-}��$���"s9���=�'�'���]��]��N��}�wr�W��ᾷp���o>o��B[J�Rxxμ[ݒ�fF.fಮ�ٙ�}38�rN�?L��.5�{ɐ�[�*�g��fZ�x���}�y,os���������~OJp;1�)�8�
};������)�S�6O׼�VM�n"�=�sq�_�Sq�����3��{~�������wW���y��#�9+��FD+��˵��^\��:��=~��;ʹ瓜�ǐ��������{D���^]���9�+�gs3{��Q�ݟg7Z����2�ۆ�d��w�+�w��D,Y�ww#�����H��N��"��j�]�b�NT�|f��8%���1��<��իd�������t�:o�7�5�ٸ�.5��Wk���0���z0��u��qm�陳��Vy�y�,��g��8��R�ݞ�����R3��{=/d��΃{}�*w�ጼms�0g4�H�qkyENO�!�~.z��N�û�`��E�ONN�zT���k�!9͜��Ӳxçr_gs�&1��N��>]���Ja���i�8x<p���e���a�<a糳�X�~4�i�f������ڿx�h����ړ0�� �z<=K��' �L8g-�qjLѓy8aÆ��U���iz�Ӄ)J2��DS��iH��l��Jt���:R��ɸ��<2hκ���!N��4�y'sUJc����t���w�ᆝ?�(v�Ֆ�+�(��(N�?���Ǐ<a�����%H~�4�.�d�Xt�+>g�x��oq�S�(��� ���*��:%�8t`h8��,0�� s���gL8a��b��ԩM!N��-S3�Zp������o��m���m��v��V��l�0���E��5�	h�4f�F\:&t�e4�I:�/�x�~��7�殚~=�g�L:~:W��K�)� d��n��8S@��?�SK����{�8h�4f�?Xw�u,<tӀ3r��K�SaM!�$�9c�@�zn���a�(�����^:te h��ۛ"])@�!O[�y���4}3y(h�=�(aN�Q��Ů5ƕ8aӣ<ar�"�	�hΘx�s���z�8�t�):m��Լi��:0 -a�`,Tt�<S�p$^>��[}��3N��Dy��idXs1s����~�v����dOO��t3����ծs>˞��ukP>���&�ߗ��ϱ��c����x��I����;�#hoK�>��l����{�s:t�y(�}ם{��w<צ���˦�$:�&�+�G�tt,�[���������ϧq�7t�um��ݛɓ��Xg5���~�{=:_��;��Nky3�S>���+�i����f�	3�ˇ�U��3��}��Y�ss�N�G'�y��������o3.�=�sVe76s����s���\���ݙ��[����o�^Yg.fn�� ��3uG������3�I����&}�v_�9ܔx�d���nx3k�7g=2vc���97�o4�V-Upb�硫�|o�G38v��ELV�I���|�>�'n�<��cٞ���F��潇{f����bm�we�=0\�)�9g�:�MTKk�ƹ}{��{�����*�:f��]y������,�͸� k�;{�#�Ja�7�a������Ô����)��猏LΛ|Tc��ʷ�=˵����u7�y���̞�}�2���B�̧N���V�3׳��P8i��{�\��4o�Sw���Ѽ�/'B��/2��re��W���u�,&]�<�?��~�۹�N���vK3�6���E��M��y�RӮ
dQ�ٯ�o�r_g;�_j�z���������:.����l�0/�<y<��\��S��o�5�y�n=Z�#�x�[f�a�s.��K�gd��3M!fN�+�2Q��r��3��������H`n{��ҝ�k��9�3s$�ّ��/���>������_���7�r3��g������w�mof,6S�o�W�Z������v&��mk�O�{U�×:Rn;١ߗ����ӓ��d��d��Zx��w7'Z��3��x�3�Ǘ�o����9y����7��χ�|-�����}���o�9����Xd
{��9ow�����M7������{'����;����y�:^���./�,ܼ��à^����)Ι�ʟ_7�t<]ɓy�Z}�z{M��������ӌ�_e�=�b̊s�y^n��7�y��.��Nq�ze\�[r��������~�3ZA⛿�������ߺb`�ft�NΟe�B1���>\b�D߸���s���$��܃3�g2g:b�ɹ���K����U$�m��q\힓݆k�����f�4�S�GW��3������G��3Bg_s�.Q�2/7�:$���rN��p�~+7�s&��0˗�Ls1t�����?<z��uU���h��N>o����U2��v=ƛ݁r/��ON���f.�l�%Z��Á�\[;F>ù������3`�{�g�������?s$|v��~�e�-�^�y9(<�
aҜ4����'��3}<;=rxK������9��i���b�.��=�f���fNx=��p�9��pT�ΐ�fw�|5ӓ�����{gs��dB;���36/����w������k���WgT���VH�9)���[�;Sj��9sw�s6��n���v�S���N�i�E�3{q�s�;�������Շ2�?.|�/�8zI�{��0��j���:L5/\��9�gx��3<b�z�Ft���x��N��g~.b���r�5q?v�
�w���}���W��`��>��X͗�(}�M�M8A.�;����d�¬���S��K�ݝ���}>�\q���z|�$��T�'2<ăǹ9�V/r�r����3���l��;~�K��;~�z[�I'wq�!�]��k����1=f�g{Js9����������;�{�Fw��/��	%Ϭ"�^�O8{{��d
nss8e9�+]�gƛzi����'Ƴ�9���}������}�n^Y�[�r��i��������=�{=�s�8��Og9�}��҇�M�_L�-�=�YF���3�Nm��?����|S�q~n��L��{�.y�Ay�ɽ�f�{#�u6�݇x�����7��&(�2�mF{�w/85��&�-�N�ƺuy�w%���Ż�_��c�d�}.��o]�|_E�\^���f�xzo���o���2t�Á������<�آ�rɞ���s��x3��|���m�vs�_O.�\��� �tKl���;����vOr,��kr��$ѾZrÞ]�I�����Gd���>�i�؟��LӜ:���͢S8�o7���_E��v�뽽�nA�z��;Ϟi,��^{��vU������C��{�N�����xw&xV�eu�e�E���{�Oan:w��C:s���{6Cw��&�Ύ{zz���� ���|?��3������k�k�Os7�f�8e���7��b��-ܜY����9U�����9Ǉ���
vSm��w����������������q����ϗ�'��>l�ꯏ��:��ߣm���Oў��П�����e�mP��rZ4z楯1�f��S��V%r��b�ɃT2Ϫ- ����J"�u�� ������eR���4�[�l[���fZ�hC=Kl����˴�g��:N���f�Bp�6������^�n2ʩ6�-(�.mu��v]�1*[��)�@e��pV�Z��R[l�\խ�J�p�Ne�m�Qd ���Q�A4�L�!��ű�6�&��K�1�i	u��]x�� �,�k��&�lē��Y�0�[]6t׋�uV�a���-%%��^K��T#z�e�N�HY�*�������%-0j
l����J�[D���5 �+��WU�\s6���5�MKv�K�R��M��BB����5��D�5�$ʭZJ�4,l�]B��F�U�0X����S�n���D�v�Q����D�
���v[��E3�ˋ�gZ:SF[,�h�Ή52�c:6���Z��Fm�CE�k+	HV�H�C�[%�$����g��$��,�Y"}ADY� ;���ՙ��׫��)l��������0Cm�-��v��{d+1]ʪ����a}�ƝoĞbXj�w:!u���7c��F7t[���U���V\b ��6/s4�js+LW���#�l��c�!������CM]Mf�f��GdM����Q�1�qFf�X��2ջ`F,d��-�&]n���b�W�U"�؝J7I�zRb�>�Ͽ4!xȍ�h���Q�?��D���,�˹Ė���Z�:���_~>_R��/҈�AX�)"����G�� JX��~c�n�F�#vu�e��yZك�n�{黼*F�T��:�.ڡ-�[v��Ea[�R�I8�舢+TC���*&�� �>v��+Z>�ʗ��shv!nn�],��u����8�։I6���[p�0n��Y�]�ź�١���{�͒�,y��,�v�l��ȷ�}z�fF^��hi�5��&�,���دq������cV��.���1���#G�2��t�>�Y��r�M�]�i[�J�˝s0�4��Ж��^�Zi�gjR�kj1BS���k��Y�N,boi:Q�V�s�/bYCC�Qj�XP>�p�ᥭf`�Q��Y��f��\KK�<"��1a�#_A�m���(t���`�`e�V,ڼ��t�~_m*ŗŅK����q�h�C���L�m	�b��_N_i�5F����%-�*Q��JW"x�Zڭ�	W=ED�T��¥�����6��j�!0H��F�&�!�Qȃ/�>�E��r�X���UQ}�錵�C�S��[�m��ײMs-�l{�U����]1���X4����J�)d���&�YQ�h��<�+|�޿� �������4Wp�f^޻ޯw]�������t�[�����������Y�S�M�>7SKj���ԐVl���4������	>���W���'�����U^*��UU��+�*�qb���UWV�U궪�U�UW�UU|�Uz�k^��Ȫ����UU򭪮ff;X��/�W�UW�ڪ��*��h�͙�g-��&6��(�celVm�����fr��e��N�7Vٚ����>?�ή�www=I$��2-��V*��UuiU�W��J��򪪊������UW�U�Ҵ��}K6��W����U�Uz�9��X���UUU���EiU]b����m�7&İݦ��Ǜ��d�����}��z��⭽Vޢ��WW���j��UUեU�*ڪ�ZU^�V�W���\UqU�*���EEUW�UUTUU\y�s\Ux���W^*���U�W���Vأ�9��9j5)��r�(�yL����ܱZ�R��n!i��-U�$۵�*V�M����H��rV�%����9j)��κ��M1�a�7�DS���F��ef�{��_w��`ٛ����?��?o��O��g��>o��>����r}�/.興�""6��"��ZB��ѤDuDQ�8���"<y�u�"""""#Ȍ����#(����h��#����)�DG^F�FQi�m�y�R:�uaaB#���"#H���""6���M4��#H�"#hDDm���E#����#L�L""4���0�m4�DiH�DB"8�HB8��"")S�<��<�h��"4DDDu�"6��6�<��4��:�l��0�
iDi�y��2�0�E_Ƽ�����#Y�sW������UAf��My!-��+3��х���K\��L2�F�-�XɫiI�av����J:ʩ� �;&�V1m*�١�T����-:���%n񷯲�ń��u@�lXZ��V�f�ꒈf< +kP�hpj�X���5GkV:b%�$څ���Y���e����4�޶X(�h�쁡�қLL�;ru�/4��vJ�Kk�7:6�\1��mh�h\�W��	��R.Ԅ����嬭�ϟj���@���ͦ�ڮ&m6��ix\�m�1Z��mlƵ�2�-��`vt��1�ŭ�Q�B�l�͹(�%v�%7m�[��eS%Ŧ��h"�\Q�����e&f��1qK��5 BW5�l�-3��Ь��Yq5 �ǚ[����]�����+w�A�.��1����k��eh�r��1�f(�ǘ&��u��E��1�
L�1?�Q��M[��4%�m��2��J[��
gg�n,޵4P!3v���J�sP��Q�%,�e�["���0ѕ®� �9v��gі�oD�	��p��J�mb�V-M�>|�u|�ANnA˪�qf�4_�D+�r�[��Fb�G"�`��5�.e��L]�
�\�z���i,u۝Z�ʋ����lM�snl˄�mn���ݱ˺�iv��j�V!5cN��α`����FhLC[t���k����˰��6`�i���fs����u�\1]��@6&��m]e��+a���`��]�ٌٌ���RFu������-�`�Df�^!lM���b�6�7W^ظ���x#]3D�t���c�&�Cf��.	�hҒ7c�n�⸙is� ���T..��XMh���*���m�ifΒ�L���m�M6`[3���Q�|�䍪�3R���Ԗ-�nv6��H�Q�3X�`@��K��ִf��ű1B;kfô�HHC�f.� ��TJ\�,f��o
9�r1�ۦ\��--���ŭ�����і��;v���p�Gmb�Z���mɯP����2�7�X��jkMA�YJ����2ƠY�e-�2�,�ޚz��Vi�%j\����V��kv����!KՕٓK��b�c�)vY��nή�������V���L�Q�nm��z��v�]�)��1�=�TX��S"�Zf[�ϧ%�y}m�*V#�v�ԗ5�����9s��.��#�J���k�b[)�ѱ�U�#�t:���8�����i�J�9�TYs������.���WXZ[�X��`V�4���c����v�%��U���L�W=����|w?�?4���U���9�s��ϟ>wuw���I*�s��9�.��w���I*�s��9c�����-K[�G�ujFJGQ�"h�(!�,��j��Id�����fֺHL۠c2Pu����[���c+�jD�:���{@R�X�44qi��5e���
�P̠X:�Bb�A�W�^"&�WG�k���e�tڲ��]ׂ�P/���4�`�t�źe�#2]B�P�ktY`dس�u�{Ĳ�&K�X]K�m�R[M��GMv�K�F���&�d*�G%���H��U��Yh*j�,�4h, 9�YuE*�V\����.��6�F�؆JjOz�^�	24`���"�W�7��W�#XcF<sɄ�ah���dXˑ�O����K����vܭ��7m�,�cPT����Bl6�Mn���]ݼ"V�3�>�g��0k�n��<ڔ�P�kV�0h:�����l��V������IYHk�!B�ҹ#��l���F�^B�,��ʨWJ��R���V��t���i�m��% _�n8�\� ne�1L*	U�2Μ�e�-1�Cr*,�&~��6ۿm��R��G�ujFJGQ���:ɇi�����d���ӥ��Xa��h��0��9CJ7�n6�j"��$�V`1iu���x�ҊՉd�KI���P�ʦ�v;�W�K�;��YFt�NS:1腭�T4�p�p|0�_�s�_��09��e�(�Տ�n���hͺ;>�$.V4�wd�����jϫC,���t�,��)r��j� ��mQE�0�Ƣa����5�kM4���ƛy�L��Z֏<�"JGQ���:�fQe��$6�B4ة�RJm�ӅuJ��g��pf��h�G�� 鷬<h^MP�EMb��׹U+Z��c,�-hf1�������`����eշR���ei�u�1�Z��0Qb���[�
)h�\0�����Gy��R٢ΐ0k9M���"�����;\��$8>��8����
#��Zn��s���XCJ��|��S��<�E)DR:t鳦���,�Q�'ʪ����!��l0��t���n�R��y@c0Ң�=�b�]�v��qێ�Z�B	7]p�jmen8\X#�����-��f�^���`RelѬ�n�����k P�Qi����cㄖ=�0�@��3va�<gOn��i�c�0��^6Y��m��ay{�U)��V=z�q_:O�m�1�LF1�_ɴmkZ���έ�R:��DG��Ig���L�/����a/���&��0��|6�R�5F��z�>v��+w]�lݱW��YmV*,�$	���c�X�����#bX�k�ȭ���\e������#5���J��4 �z����j�c���P�&IuV�FnU^cK�ի(d�j|ϝM�;%�A��I�����;g};�2���K���m-�G�g�ICCbU�:Q�^�>]U;��#�0j*��Y�L,��82EB"zm�I�:0ڢ*1EYd���r�#�M���6�(��[]��6�!g���`����|cP15f���a�s�,GX���p�AӞ�f�S�f�ꆙFU^�$(�0����-��K�Lij펙���a�ά60��4��j�u�����SM��R)y�D"���)�u�6�m����ު�㢁+hA+zm�km��7hڰ��'�� �G�eS|!A�!Z��ƭ���Wm��1Nc?i�����iJh��s(�m��1����C�QÃ6C��d��>��q������ڷ7�<�:��٧�١�k��w�E�#�tݔ0e��T�lkF�F��K)��(����]���0�K�8a�MN�H�΢"0�#��E"6t��YE�X�r�+Jی�m*�#m���E2m���H�Pg=B^h���R��6Pp���ܱ��,T�z�.��'��{8�i͓�nihd	��8��R���o��5tcn�Ր
*+h��Ae�:(�j�42cta��҅�0�JR������h�����qB	v��0�fs�HkYYr]����;�
5Ս�5c�{9E��2ˎ3�����}����s{Z�yh��yբ#
R:��R#gM��Yg:����:�m�C��3��!ʡ�3�]u$����� @��{�e(S���C�^+!y���ŵ՘Ϧ4,�c�ǔ��<�(��R�`YDM3�FI#��t�������8�YK`hB�`R��C�܅����388�{�]:{�0,��hoZnY���T@h�B�l��`Y�S{B��i��NT�C}o����g��j7���?g��l�V���y�V��)H�"�JuN2a��mW��{"��+g��i���X�����í���*�n�ql�Ă5'#��֊������x�G~"Mn1b�7� k�˃i�;M5�in	]/&�u�L6����HcMH�(,e�k���Ҩ���L��
�h>��,� �w>���ݮɹz��ڰ�Ɏ�9����	���x]�g�ǎ.͕N�)�i�g�U�}SU�#k�j��fi.9�P��M�v��;;MPB����Y��E�Ś�z/F&4��:Q~v���{�ӻ�Hl���dq��'D+=��3ƊI%E��Mh0��y_q���q�w�siJEL��:�ꅣ�m�<�L�׾���M�g<Ԟ[0���y���z@���f�(��cm1�ߘP�I�T��Q�����*k�y�����Y����F��dHA�%���3KF1ai�KǍ,]0��.q�S!\�R���DG�uh�����8h�YeY�M��N6��p���a��&��xh@���6X���]2�t�21�%�J���%�Vmi�iXQZ
�q��T�m�4P�F'[{���Tb�$��U��q��v��Km�v�&R_����-̿�P��~G��f��a�F
�S��oS����"���$@�+
!q��:׵못F��-l	�:�������6�ͱ�:�f�fל[6�ml�Kj��-�ym[l���-�mn5l[�k+f�Mql፱kf�[]Z���3�<Ǘ�qkjص�kf�ͭ�FV�;Z�Zٵ���ml�ٵ�ţV�X��ճkf�y�-���E�ճ1�g���#4��yųk[Q�ml��m�1c��Y�p��!���3c���%�<CÇ���L<N������cxųkfض-�ymZ��ٶ#L�l�[6�k+eխ�b�f�ͬ�0�a<h´Y<?����c��Hx���G�^'�ñ����j�<B`��ه�c��8?óǊ���6|O����F�c��r���y�u�imZٶ"ߚ�+[q�3�����6�myŸ��kg�-l�Vűųlu�c��83��l��=��Xl�2���G��A�OJ<O��>���������~4O�<V�#�;�:ҏ��~���1f9_��OZ��P��}׺_�_��WTc��o("�[y �}���a��HBM��m ��)Sm>�wIV����1�(�f��cv�5MFV$�,�g�Ϧ���5��f���T�%�Y���͇��4�:���t�YHoL;!�u�D���,hN���t�������T����Q;�m�oO ��9��s&��;y���q��W��_{��������rI*���w�e�o7wۻ���*���{�|qռ��ky�V��eH�"��:�M���af]HI	!�b{u��nUo�fF5�M��-��i1Y��nzF�U^�R�l��T�dK b�i#��ѭ�q���[�tB�2����S6�qC�k��pTдwc�C/���w��1SH���7x�Y��7����g������u�rU�m1D���C�����c�J�����S�I?j_��Ky$�wUY�������f��/ 0�e�@;�7,�LGF/�ݔ�%��b(b�`�Z`�h!jXz9v����9U؉���g�b�:N�;�����q�7�gu�ӄ=m�������66C�pix`�am$��f� ���i-8le��J���"�@(�5�#�"2����1���;�c��sb��KZnc��R�9�%��a��0�eO<�����uJS̼�)�:�)n��2�N6���1��$�m���+b��͕ ����ѷ��&�hKt��r��UHߌx�0`S(bZM���n�o/gM��]�΅�\��0�LX4*�00���J4�[��d�܎ݐ�bZ+1{I��55f�$�0غ�,h6�����Ņ��=�7����vM�3m����8"��vA�nFJ �i0)�o>ˇr�zk�OA��dOW���9���=�:�8+o鎊�%G`X�h�#�_Ε��7���#�����.�"���R�x�e�KI��Y���9:�%x��a��-,F�����HT#�t����sM���(���*�y@pb��@�nG�:�S��6+����^My1&���E�,�� ���&��<��g}8�xw{�����<��L�DR<�T�Xh�C,�9L9����aJ�*yQ>���8�O�L�QMx;3#T�p�#B�3��M��.�kJ�rL>H��ǖJ�|�lYZ_�`�Zڇ�SD�Z�#Ƌ��a%Y��dRU*ܙ�o�*��4]�te�k5F�t1Im� �����)��		)���x��i����5#�?v\՗}��<{��ק�*��n�f�&�m<����1��s�A�G�ﶫP���Q���8Ŧl`�3��H��0�Mm+n兦w�i��͞Zo]+GgC�l�g���vvf�[b"J���A)I�gYeңM���+�����_41j�gt�j���B���3�4~�sŋA�4�Z,�LX��!��, ������L)���LO�RG�I108��\X@Q�ф ����<`}���<3��6�n��18�ɗT�nɎ����c��<Zs��8����7D���{��B4-LeڀA�	ǮqQq���Q�̮��w;[�	Uc�Yv7�0�K� ���CB����9����k3�Ht��t/�1��1k���1��b����������<�DS*GQ�)�8�L0ˎ4ێ9�p�R�&��=1���A�
(��3�ֱ����ci���\9�vh���KI���B��nq��Ќa{��c�l����p!	c �K
N҆�(h��P�	�\T͌a)������CΛ8G���8����l�36-�D�a�� 0K\!f�H�-QI�������ww��<�;�\!ݙo<Gd�;t�DGKc��]�oy�����ݵ2��#X��*�Om��"���RQ�"�QY{��L��T �uܫˈ�N�`hi3�цƕ鸵�wfv��7~;��O�8x�e��m�x,޻�s:Dٲ�w�É����C���҈:��"����x�-���jݓz�,t��tyM�m�ӭ>i�:��ߟ�y��DS*GQ�)�8�L0ˎ4�=���g	������4.Q�9)#c&h�g�E�4��8yS�����T�jϓKDZ(�a �(�C4��܇����v��C���=��$&���Ce!RLV�I�041���f�l�m�ٛ�	Un��]�n�o�>Hq/A��P�M�m�;6kl臿���ն֜��f
��2�6+���~&YsUR��T\e�cH����D�v�蛝9��;���߅��t0>pj�#>e���.���D��w���f�����αR�4/�@�ŊƌL9��P`���`��е��㶝�:@�g�b���3ca��%��h�7�߳�u���z#�`٦����`��m�Ė|0:�7V�Ia1�(�.0���7�1�����??-�<���h�eH�"��:�i�qƜ;���u9w���<JTXIɾKMz㝠o��X�� B�Ęha`�Ģцc���-1�^i��*(X��YM.�N�aGU�1 �DMJ{�B�GtScf!&th�<�����Ώ�@A��3[�f���f�'�
Z���m�!4���g�C(g(P0-�K�#-�#k�n��̓VD�-���YI=���wE]�A��
N� X�U�jՊ �=��F�]n�GXk,pZph]jP��C��7*��9�h�AH2�!���4a�at�I��Bؘ֐�o�ꪪ�f�p���G�hpx�`X����hh��hg@�D_.(���sN���/���mn�h���Z����E#�uN-�\q�Uo��l���W#���M��r�[Y\���r�PNeY����X!2 �c�q��c��Jk����r1�j����j�չٶ< ɶ��MMT�Shj��ta���S�6Q ��ؿ�×�\��s�|�{�Wj�eɺ�Q��lW��|Ϛ�R/w��cg�z�<;t��U�9W*QOO_�-߻�,�ۢ�v�@��%�	F/�~����S�_}�~h���1�Dqk#`_G�0�J�뤛�7����4l�6ae���;��H�g	f���G%�il��C9��ܪ��<KFгJ��coe����� �CAыc
��I�i2G��p��Hc��2�IM�)�Rd�&�@L s��Q���1k]e �M�v��]��c�=����Q�UU$�=|a�#�umӇN�GQ�z�z����X�z�7tt��=�{Ɩ�
�K�Ԉ�WRk=�j�8��t��S�ZIq4�Ҧ�T�CJG88/n$hb�e�v� c�M�g�`�_s�sE����1��`��ik~[���ֈ�4��)S�qme�Y��F��;i��}�������ha�IH��F�h�}��m���' �LwN�{y6�}(6�����/��5�(�F�����A�L83�������3�y��S���,6�A3C:�y24�&U�R��44Y4���щB�l{�I9��;��
�Z�{M���6��0>)'E((dML���7�th�I����1Y���\�&�+V(��8�B��>Y>ď��ē <t�Le��dC�r�t��i�3��h�@��I&��E��M�1x�7C���8ZG��
�7��q�vY�����!�ݷG���P�&�0�A��D�7���B!`racG
ZߞG�)��)Hۨ�G���0��<-6�ёF�1&��kLlm�4o�h��6�3g�/����wA��hf��Jr��H���@pjƎp���G��u1y5� ��E�[��q�����@�t�w�B=^�{�<�)\;���&�N��wt����N��4X0.3a�)ʨ(���pdq��A>��
ϡe��k�ߴz�}7�q��1�a�q.�|4_�!�;�=�:Ҷ������'�n�:}��Z3�nj���GS>"5�(ĶQaB�W�	:m�J_��c�L�ѫDe�4a�8��B�f%��_/�ݫq��|b�p���A�>oq3E� ��be���G"��[�'�>~������S�ԥ-kE)GQHҝS�h�.��5Ө��l�660i&½C�-.�#��qQ>��� �@��ь���@���� 1���UUiC63�GR�� 07���cFhk@��YrGJ�0}%��Ӻ����F�dJ�H�j,#�s,�t��ӎ�i㇄�}c���h����@� �2���<��5�d�[x�ֶ��q��w5K��$v#�c_y��L[�(�0h4xc���WF�/a�#p�h���r�A�n��kyY�Ӿ��:st����ҲቝL�G�3`�|n�D�}[e�w}z��_�i+�g��P4�;k�4iD�A��P��������T���V;0�6C�I�l[��ٵ�kfص�V�+[>[6�ی�fikkLZ���m�-my���+jض-յlZ���St�>w8�ml�ٶ-l�ٶ<�ml�l�kjص��-�[6�m�Rڷ�j�f�f�[��_�S�e�?6��3N���m�ml�l�ٶ)�cZ����oS~�����xe����?��x����OÇ���~4E1kf�ͱ�7�Zڶ-l����՝�!���d��g������2x�<y�[9[+Fm�x�<[�el���2X�~K<O����D��<O���h�4>�"���C
��3�e�մͰ�ٶ6��L2ż���b&��g���6|V��鿏џ�Di��iO5O��m�X�?�ͭ���V�ml�l�[����g�l�<3�<=��׎�Xl�8a<8Bpg��aD��x~'��)��ٶ"��[,-�-�-������TN�g�ժM�9��MyNfO�y�Ƈ��C�[�h+�fj���q�Q���/�mpX}������w��������u�=���������C*׊n�v�3'��̌G�9��͚z=y�T�@O*����g�nm�>è\��3�.js�w�_E��>H�o��K�}6K��wΉ�{����c�Z�gE�C����\l�kVL�ł�5582;�s%t�y��|�q7�{�,w�|qʮ���-U��=�5�ŉ�\���L�J��g�`VŨ���{�kGP�9�>(PTLX6��%$�ܙ�v��<b��M�	��%���ӛ��;7*o���XCp<o��B�#�D:�F�Uq;�H�ۙmw%�,��}�t{;���,�h��s~�\��j�C�Ⱶ�9�ۜ4��Y��'� �iE�q��=�?�{�b�;�s&�֘[k�+�>�u�Zӵ�*b6mku�g,�^G����˖S��n��.s���6�[l���V:b[*�%�;�M�/1iSh�4Pk4�;j45�:=�	[�9ݝ�ز�Lq��JHm��+Y\@6��v������O���
Z�`�l֓k����R�Rjmm%1.������$t��ę�m�F��F�]�4�Ri��0�!�����4|*�X����4a�i�Lm��l�D�1+�-l���%D��KF=�1͹;�WWN�p?�>�s�߻������o~���o�;���������W�.��󽻻��ޮ��䞫�����ukyŭJRִR��G����8��2�.6�K�Ų[r�2��S�
]
��ȩ<�p#N�J��@�d-F��c��и6�J@?�v�OYj�e�ΓǼz�Ў�s�f��KhlX�.�e�.�٦(kcil�֦tLhL��6-���U�2�"i�$���\m�ij�L��2�ӭ��b��h�q[tܻr�Rݦ��-��(�PٻYa�:�*��+�vt%��0��zzw�c��j�6��V��m�f�v�3����f��M0i�K��C+�{-��l�Cp�
�P��ڬ�		�ۗ����'�_�=��6�ַ&����/�G.�ڶ���:By�T+{�=;5_9�Y�ڌ��կ͍�'"ŉu1Q|DpaVDE��"��}�L�bZLLi��]&3/đ�O�P�n(d&Ę�l�[sODq=��7w��;�<0���7$�jV�[phv>RJ
`ű	��YIz�6i���gK[<����z,�G<{�9�rD�2vT�(� ���
`�=��ic�˅��ow��m����t��p�8�r8��kƅ�x�sxG�o�;�j��N閌��0ic�d��I�|��H.�+/�r�MFX9S,_�����+�TN'�Ih+dy��a�m�S͋N�Yb8MՎ�6ڲ���;��PƇ�`2|:�<�^[򔥭kR��E"�[Fq�qre�%5�+XzJQ<�U͏(��t96��n��'y͋�:[yx�:r%��P��M'��<Y.��Qu3C�(����g6�r(r��`Ž�5�naц&�(Abh)P��Q�r�P�֔�|$T���F�� li/�`�-�%%�ϓ<x�6�h�������wV�]�U�
ِ5�Vƻ@^�����饃=�|(14�L��҆0�`q0����
w��g��f�U8�[�ߧ��Eg��R=v��{��m�9��Ov]l��Ch �{���; �Ѡ�T+�3��-���S�u��Z���kR��"�
uN-��ˍ��m��ȉp���mT�5�cb`��iz��+:y|b0�׸62������8�:0�0�d���*^���I�H X0�������3��S���8�r�n��1���Ӫ��62���0`�џE=8�u���Q�`�X�̭��VQ~�Dz�%�UU8K�w����h��c��>q�T��(���Yͫ)ta@������em�A�é��n�a��}��T��yo��XP0aѐ�v�t㐋z�"�|4�4�8*�|A|p���ӧJ>Cx�5��b�0>��A������:��3��<����JZִR�DR!N�Ŵa�YfB֐�����,">��&,9��$�6!�M�0g:j7b�{}(��&y4$����2|E`�8���l�;qA�84ih���x��+^:��!p����̎hr��C��0hb��G1yq�,I�yOJ�1�!�j9ALl,xہ�ѱ�a�=����� �r.4���&���#G�&�5c:3���$�alJ S���DVɍӪ#��Ig�wd h�� 0�S+��A����.�FT��ߑ�-kZ"�DR!�G<P2ae�a����զ2��0�1K�5Z�$�f'��j.
3�E&�TE��Je�E��K,�
�	��e�D�'(خD�J�4���`3�2h���QW�ªܨ\��f]@�|$%��˳S�"�ն'χ6�
5S�H~��,�r,��Pm[�=3�T�;^>a���<�db��,z�
����l�
���X���1$S@�81@h+�x�j�DE���iɣ������x꘭ߣ/)��Nc�1ǭ�~4�A�H1�t����G�Ͷ�+��I��a�߉�`�|s�[�;ז��.��@��-��tn�+4�+K�Jq��b<2����������=� �m>%������+nTl�%U^=6qC�8mh鳾<�롳�~��T��1s�}�g��yh��?#ȥ-kZ"�Z)�T��0ˎ6�����0���	l������Z>k�:=-�l 0�a�p�FΗ�����!�v�܊��0ag���_l��K��UN�UT!Ü9i��ei�e��4p4.�;7�ߗP��]��8�6_���
�����f�^49��'j�ImV
��hV�b��
/�T�_�eR��m��ԙ�G�6JMpg������>������J%�u_����:`��y�"�꩔Z�`����/��c�$q�����2��V��Sȧ�h�ukR ᣆ(0�
�hllLh�E�#�_;�ʩn.lttGN�͘�ln���B@���$r� ���UJ�p0a���E�����N����\��HTm�R�w*�UUTITRuR��nT��M��˦4-$C��srTM����"�1t��9�3�����uy�tɂ�
���5�Ӈ�6l�`0�ln�Q�k��IP�>4p0�ha�����|���CG�{�o0��y���)O�Z��֤B�S�h�.8���e�K8��NC�,:���2V�����h�W�US�>ֆ>��e�@����o�ΛJ��{��P�L�:ӕ0G�>K�#�4��!In#�f�IupÆ"�ӣ���}�me6Vt(`���%z��{�s�D�����OX㮶1:��S��ㅅ"yJN՚1k��+������0a������i�z�X@`ÆY���$-�5���
_���L�8�����og������ﺧ�i�Z���S�ZִE��hS�qm2�.8Ӌ�7�e�h]�t0�5��l���_��I�@���ҷ�wj�\*]Ye.�T��L�ܕ�3��be�,�f\�kf`����[��%�� �66&9{�������/��q�&����������0�����[����Ơ����������g�&O"89ϛ\�&6lq��uyz�kS�y�����aA@�6R��GM/7���V����V���j�|���{��h�3��+3%���aF�~����u��� �ϭ��;�� ��,�Ѐ����(�m�m��C�q$�i!*,~��?Ce�.��`�6|�H��ѳ�p,����C���$z�:�#FX���[@>�7�_�faְ�j���=�x�������X1���k���FG��$�8p��(�F�E<�Zֈ��jZ�[L�0��H�Li���aψ��Q�X1���EIW����o��f�|�Y�`Ϲ��p��)p��W�GGO�o�c�:�[�9+�9��7ã[-lLf?x�q��=0�P2,��\��r-����P3����	�n�Qt���
�io(���:�i���~�8�q�`ù7���r��8��~q���;�]��p�x^>3���$���$ቶό:���b�[�7����q�8�^g�3L[�
j�Θ�-yųhͭ�[6b��V�Ql�Ɩf�melۋjض)�[>m�Y�Kj�ͼ���b��1�<מf�ͩ�8��l���̭l���Vխ�q�bћ[6űkf�3kb?W�ǈ����r7Ӥ���1kf��V����~�?3����������z'�����x�����O���;��~0�(��x~4n��lZ3l<ŷ�[6�ml���l�kf���gm��-l�ٵ�kf�f�ʹ���z�.8ͺ�Vͭ�1�4���Dg�����(�x�!�x��=���<<(����4x��:<O7d��pq��<O���j8M�#��������g��l�:�1�#1L���?6������o5l��cL[Ŵ�ͱn�lyi��583��ׇ����T�d!�~�C��g��xOǣ�ºt�TB`�x�7��~:O��7G�FF�%����Y��\�	�˸-��~��#Xt:l~�L|�/of���I���ڇK��7��Kܗ���l{8��
�^��b8&���%&�h�ͮ��U��z_lۣly���'%�p����駳�z;�����ܑt����vYz�e��O����Y<������� �J����=�.N!q{v�׻ͷ�V)~Y�^ݼ%J����4}��Y��&ww��=���j�rJ��{��n�RI�$�$�����ݿ]ޮ����w}�xm���Z�O-kZ��-�8��,2�
0֕hllL��ߋ?�M�����޿g���.�v�h60�z�a�q�P���P���m}jh#�H�n��`Ƀ}�G�ۄѓ��|\�-��3�iMZ؄!Tr��wU.\�9
9Ë��т��/�a��c_W��ջi�ͮt��I�=н}���<ލ��ۓo6�4�><x՜EQ1��ix��OQP���%��&	C�!aI(�6�Z�O��%���0c������<�̻�^[��K~E)�kZ֋Z��B�S�i�q3y�,���1�e�6}�W
uR���]��,��1��.,,�C)���o���r;���S�m�A�5�G]-0��K�3���^U���9��-��j���2�9�Z�,2�#d98�f�c"�����l4t��k�41�c�m����������1.�1���t�e��g�/��8z�U��Fc��Gy�I<{��☚�J���|:��3�4Qd�F��6Q��<�i�F>�}F^�����𷔌4��<�~E)kE�h��k)�8��e�e�c��&��N9q�ܗt{��F����ro�s&ń��T��KaWZ�r}�\g�q������bX.c��i�ܮ��ID��eծs˗�+�԰R��+�Ncg$ǝ�@�!B�W�"�9���ə-P{���{�ǿsI:��;�߹�t䌚�7!���[��$y;������4�iU�f]��<��1�c<�u~_K��*�r�M���81�˦�GR���(�f�

�e��ʡ�,�����C�3�na�gŘ����_[�;��lcK���|���6>�,><LFc�3Ǖ�lf��4lh�C��E��4m�ڱ�����i �qZ������XUUR��UԻ�RrJm@�S�9�f�+���,�C�nѥ��o��L4���h�-kE���-e6��,�㌸���k`�Cc`���*9��W��)+40a[5�@���${<h�J=*Pc9���.�/6���ߴݯ���l��7�֌���|������Y0t����y��6G>g7m�R�>m��Fͤ.iQ��
>2=3�v�e�%��u1e�V��)ee���>S�h��|����×�]�USf��[4B�x������V3y���!�ɽ��Ѳ%����7�i�V�����"���֋Z���S�i�Yq�\vLk���s���`��7&�5�lvajm���G8���]]�UU{_�1�>[!�鶔0���va*�c>7c��[���㮵��\�[[l��=�_��J�y��ԝ
Bj����Tp�d�0��#X��hß7�e����㌝0��,��"��������t �	|�E)t�cZ6D�TB�e1m:��͐z9���{ͲM���G4^��o��)�2���d۫ejDE�")kZ�h�����6�2�.C�W#�J�$��c�6����c"�9���:G����
 �E"X�񢙵f�(��	�n=���fZ�7�C	����:92Eո�83�ѽ ������F4i�_ee�1�/cc~��i����~�s�8�߿W��n���8�OV��A�8���~<a�z2�f�}����yN/m�g��c��Ly3|�'���vm{�Ea������m��*�]�:h��(�a�.�~S������L0�2��:���h�Z֋Z�ڛF�e�C�B5�Ҍq���[��0n���ܔK�X�$D`���E* Pb%,��(&��eiŕ#rK{�,�'��lkXۖ���2��,��an�'V
�m��J�kR(m�ֵ���]���rKb�e�ll�L$27T9�Ƴ+ׯaW�o�d��ߣn-�F�c;�m�<r&r���
�#�$�y�gd��ŉ��	%H���?&�T|tz_8l`Û�g�G����P�n���e�����Ls����U���9��43�W骪���3G�,c
>Nh��3�Ϳ�H�NQ�C
A����ӡ>���	d!���N}-r0�cz�R��XÀ�s��GFo�*��R�(+$�-iejZ�m[n��gww�|7wdn��o�:Q�hHF*�rȚeV�n���6���B1�Q�G�TmP����QFf�N��~��l�JG���Zֵ�kZ�kYFѦYe�q�R��
Je6�HJL������1�<_U�<3G��
a3��Ҝ�pz�H:C�(����"l�P�q�6}��H�0`��������v9GJ�ob���ڡa��8�a<|Q��0cZ&���3��{����J�G"�Hb:Z�M�˿�S�,��'KҊ t�ş�ݲ��Y��,a���g�e���I(��6Cttx�n���T���4Y�Za�����")kZ-�����6��e�e�>���;���c3�I��g�m����kW,eG%l���;��M-�0܃d�:���F0�Mvg���9M�F�8}Hl�6vǱX�o������N-t3��i�Xk�>�V���6=Uֵ��]F6Q�1��-6P�!�j����d0��a�Ä;�AL�T^�衈e*>�>��L�V�ճi���(3��
�i�{�G�>(�F�2��TS%=�>l��Xƕܴõ���?6��)��KZ�kZ-h���ѷ�ea�0�덷�A���A���tllõ�ӕ�G0v�"n�rN5��(��#�����JÖp�'��>���đ��#�TKu>�GDW"��+ �?gY'�/�D5�B 衆;�ن�m���م�����v��ccܣf-�6�����c���%:�o��M&`1�t��h����)ix獔V�/��|1���!�[>n�Vi2��t=��ʔ�T�,���Ҽ81�<����u�����"�[�Ȍ�DDG���"#l!��#Ȏ��a�F��E)�m�T��6���"4���<�#H�""""<�#M�")R�E)O6�����"8�Dy�Gyqa��!aDG[DE#��""""#��4�(���������q��m��,��0��km�����a�F�C�GYDmS�G�M��"4�"""<�ԥ4��[K[%�h�����#(�#��<�<���#n��Ha�#(�6�N�B� �DJ=�T��n˛�}N4���d�k4��x��n�h�6�3a��䀧"���3�*%��%�U�����M̴��$ZR7뙉�?E81]���Ѐ�}U�w��zЍoD�77��i�=s�Z�M̺e331a�S�W���d�C��� ��j52+�L�v2р���(�lcM�k�&�aa-B�dگ����3�u���0�UA6�̼���]9Ř�_�8�A�wYbɒk�2��iv��nf+���!��5�q�w�>�7�.�PQ�hD�`D��P�Жx��X��x�/	[>eS�խ9�ڂ��Q��L�-V�V6}2HQ#��A)�޹q쀫ߢ2�/F�����K\Y6P�}�Yl����8���]@��,)QS&�{d�����Zeq�d/�+�A���oǬ87V�Ũ:�i�a�[uλl;c!mS�ih�%�,�R�bm��-]�2\��j�Ѻ���t��ڛz',v���d,m1Iftq
M4���R�ba�c�ء���=P�tQo[��;$���2���9�(�M���-7h��3�0�k��\�µ
%iu�lC�+�����bi���I%�~�4E&�'�\B��6�*�/�	"�_Z�'�� b�w=�}�z�IW$��{��n�RI'$�rM\�{�߮�WwrrIW$�����n����)h���h���Z�[h��2�.15��}t�Yc�V@rE[lV�ZB �14%�͐4h��-�ԩ��f\-�c�@�vq���⤲�<�i٭�L:�V�i1,��lE�h�%&�l6q�^m�Pű����&��^����`�4\�P,l��f�bR�0���cne.��]E�uM���Q�Y�j:�t-��frJ�M�-�n�c7���j8}~�@X� T
�D�[V��7��V���\T6Y�gTf��`�����060�QJ��9e�QM�	K���l�w#�Z�'��U�d˜�q���'U����q��L��5��3�����˙U��Uڞ��b֠�l�M�.>��h�dq��Qh��䨅&A��%F-�[�[(��ӮCF�٥�0��E8n�6l��Z-aTP�ͭwY.�x����Q����}D��j�t�)wM��$�J0c+�a�Fc&8�F��ې���v���.B%�
<�kE�a��=�7��6��E�`A�i���[�l*By�ֺ�Mk~��E%2��UT�xC�0�CdP���/_E�:s�ʫ>��<�ˮ-O�R�KZ�kZ�KZַ�Ze�\q�O��/3��R���qU�0ຈafqi8��gFP��7{�9#�T;$�����8��cM0[�g=m�9�pd$�NF����4�7��ކY�Ѡ����E��۸�Q.퍌���o.�huDlK���JiY������Ke0�kޫ*�#����t�K�����Ő�nٯ	Z�5�0����:�p�7���1��8��$�e�/�%��"΅0jsE�ʾ5<ޝ0��q���m���u���~e�)�E-��-kZ)kZ��,�D!0��+��4SJ266`�5��r���F!��f��O�ű�T�j��e���{����f�� �s|�r�|a�63��2�c=[��V86R�Ж[�kn�`�Y���Ţ+���(z�a�(��k��Qdrh�cC^�1�,4p��1p4A����9)yf��akMK��χ��w=ݰ��X���mF��1�=�	�0`��GY�u�c��l��u�[y�R-�-KZ"ֵ�KZַ�Ze�\ah�y2�J4-���{m��q��n�PrB�l�s��D,��Q@����챍U:.���C�w�;ʬp�p��:xjU/x�0����h���m��Z{�{8p�Eb`�{TP��Qҕ�z䌡��}�d_����
�yLm�x���j�7���lݖb�Æ� ���6pѣ�vq�)l��͡��:i�GW�p±C�d8�y��:��)��-kZԈ���qƙe�eƳ~�U��w̕�*^\���[J������d�0�p��R+[>ex�&���b�Q'Vz7'sK�o|Y�d��62Cư�P���7E{��(+,�в\ǘ�>����m&ЬX*��U�+��J���H�m�e� _���Z�W�m�@�!	E2���nG�L�+zw7�7{>��S���=Y�>jy��b�m&]k3A�{�j�ufd&����g5v�1e�9IeE�>����Y_����cJ(��r��q�ǜ��`�ƌ1�~c
u���F��7h��jF��ሳv/-i� f�k���F�MŢ���mhg~85�����2�P���e>]2׌!ç�#���ᲆ1���.Qe�9a�j9&�J��(�[��YJ�=�*�ӷT�.�ǥ����=68P�M����j��3�����Sud��Ciӑ��e-�>����s�	^L����"<���[�~Z"ֵ�H�Z�Gi�Yq�\q���66`�Ժ�k�ݖ0�ps�$aZ!����c*i�|ǘh��"��E�.-ֵ*U�B.QL��B�=��f�O���7/��{}0�)�l���w��M��w�S,��mϛPN
�~����2�4��zIA�i��0�x�Gǎ-*�s����������1�-�a��=/q���A�-WR��c���^��9����mմ�E�JDZ���jDZ��8�L�ˎ��d����RB1�{0�;�2�(��^�q�cd4h��K�y�:���!c|fv9cj�ϱ��~����)�ߏ��q��=���1|!	s�Ϣ���j��\�t�V��Ԥ�m[
Y���!s�Q~VP¥6��~C[{4h((c�m�o]m�����ҽ|eU�g�9��i���D$�!e��o�S���m�C�(��LG�.,��3��oE�l�Cj�Y��8|p��Oȵ�-kZԈ���qƙe0����f0Uz0l���|��n�U#��w�G i�Y�>T�A�,��cj1��̬!�Ag���
71fJg�:�34ݲT�_�W劆��[�(�k�[��#�{�>M��P�Z6<!�Z�졜����%_-�X=�64�#v;(aB)Yy�k�F���>zdp��8��L����-��"82�������/b8���~ӭ������q�m����y�Z��Z�k[��M4�,Mb��D�$��Y��.9q�,���C ����`�7Ř�����7f9�\x���3�-2�>�"�mj*ܒ�����2��9��)�f��V0K � ��6��5�9�����y��愖<y�R�?~��7n��wy�M{�>��2Vf���=��޷��&<����U�a�)�ݹ��m>�Uf��M{���+�Yɧ�kRQU(���k�Kl,!��0�<Qgg�6ʪέ�Y0l���0k�ƕpM�a]]j�[{���xl����~�D 1�	�ѽ�6x���u�h�"ú>2���?5�A����޾�^���l���1�q��=f�+8\>Vaå0����(�'�YKecT%$�F�Em�ͫ+�����3�.�Q,\^Z�fYG~$�41yh�E����L�7*��F:�G��!�
4Q񇏍�H��kE����8�$!��$	�|�B��(�B�^c`%N�kcc`�(��E�c�_��y����a�����k�d>0ٴ^�0�ˌn2՘0c8KV�vQg��``��&��ŗg��q��\!D �/��x�,R$Зxb| ���m�ݠX�Cut;�MT��f�Ŋ��a�	?�ލ��� 3�P���Vk�y�`�\)}�Y�i��6g�`ÿ(Nm6�/r6ya�K����ȷ�㨈�HDDG�GQa�!�DE#��DDGQE)JyמDm�DF��Q��DDR""���DR#�Jy�DDG�є"#�"8��Ȉ��B0�#��a�DFфeHDFQ��DDDDDDDi�6��YB�e�Yq�R6�]ye��VQka�Fѥ8�E")�#�"4��""8�ԥ)�)O-l��Ե�kZԵ�DFQ�G�E8�:�8���0�FuDGH�)�!�^��O~��X~己��`��ko?fo�|�ݏ��Zo���{����<��o���q�d��%\��Ƹ��1@eN����$E���[�u�\11q�w��ἂ`ޞ���Z>	���m�6Z�#{�J5c��.�&��b.Zq��謐�4�BTMf���w��o����i��3���{|���V��������UW��~-~{��?7��U��ߋ����mխ��JyjE�h�Z-h����qƙe�e���1�G�ǩ��Ώ���W���WD(���Θi|B�[mB�Y��'t7�e���h����kM�<��#�s�ڤ3�(�������B�%US�������]�H�B<�a�Ų����<�.�w�s�m��O�7�GU����b�B�1����E3�:����#�j"�X�]{<i��F���|�_G�T�W��3���6�l���a��O����H���-h��"ַ�e�\q�+�i��6urͷo
Q#��4cg�5�':1��!F�
1��]�/�>Th��e�p�v]˖�ܪ%9uq�)USN<l�:�f�!� �0��,}o۪�)��h�\�vP���>��Oİc)��5�tIT7$���aдld�f����D(�E�<E���{��1��&ѼQ��!�P��>L�I#$��;Cq֍�/�n�0hf��7�)E��yKZֈ��kZ"ַ�e�\q���pi�t"�j5:K�x�U[lj
1�"������cV<�Y��P�(SBz��E^�mw>�e!v-�Meh��HM��[I���)��f=A4� ;Ͷ��i�&�Zb�`,I��il�J���E������s5�>D�&3H�)�c�{�X��r4�ev[�2�)�o�g^JE��ceu��p��1���E:3,4XA���K��W|�3a��0{�����g�2�7C<l��X��Y*����)Qdca�hm�g`�����ttQ�|�sՒUp-fÃD�>���B�Z �\֩�\sG�F��+!D�/P4td0�~�_T�H�6�U*�N���PFGNG�?��ೈ�K�0�.S��,�dV��*��6|C�4|Q�gy�ִE�KZ����8��C��m6�ii�]�͍���3C�����D(M����.�7DbX��1���p{4a`��c���$�ٳ����[�6��S��)��XA�X P��j�Ӧ�U��,� W��O߿>�	?��;��'#����W�y{	V�Ir�/~��.}�|�x1�����\����I�ûo��C	,0p��J"c2ȡ�'�R����w�>��hl۬��JE?<�֋Z"֥�kE�h�2�,��*{8c?g�Κp�v�Y���5��P��if��n����'|oz)h�E`Ŋ��6����t"��a�;�����8�Lc����`���7Rmu���cm��U[S�٨�ʩo�c4[�7�uZ�g1Yc �"��@�d0΍�P�QG�]��ϽE��/�|��n=P�!��Q��(aj�Ge5���͖h�y���!��,(�:�k��\��-����y������kZ�kZ:㌲�.8�O��%|0������B��ݣ+
Ǚ�U���oT��j�籃;�裩�a&�9	S�(����`ʎ:&H�8M���V�%���xᑺ-a����>DPc>q�8�NNY�`�."�t�Ta�VP�xh��!�q�0{2��o�D=M�C6c+^n`X�d�|t|�#��7��1)�
!�<|��9C��0}cp���o���-E�<���E�KZֵ�h�2�,��+r�Ʋ�_"�\D�V���Iac��6}�eR�B1\@����Y�u\����,cZ�eok�z��c��r��.v�	���-&�	��k��r|"&�0`��B���7�����-۟��j4����unw�Q���������������G (Ol��.��W��:,�������f�c]ɞ�����U�U��Wﲦ���c(`�^��$r<�����Dë�--a�og�/��3���1��X�<�R�qO)��8i:(ٸih�y���ǟ=eU�U�h��g�`�������J��U!N�cz7�9:o�42��%��T|�d���z��Q�5`8F ��!��o�x���z�՗��Ϋ4>Va�t���>c!�������N�Y�e��-甈��-jZֵ�kGL0�!0%�b&����+K�<B�ha�^f��#nW����m�l�������yY41���3����>0 ��}�֋4P�n��)���N��j\۪��m���A���<�Q��&��[�ӊ�����u����P�FgQ �Z����p�w*o�������eyɡA��>���[��Qka�3ؖP曶$��l~6���1�xB=�ih鵚m�a��<������E-kRֵ�k<tц�!�Q�,�ʪ93Ccbc<p�cuQa�E���9��uU^�pT2����Ǝ�)���e��{�tt�t�8�,�Y7W�����)ݷm�J���VT2�*�FO��?��y�uu+���b�
+m]�a����4h������6���!�h�֛���D�i����n��^�T��h�8��9���G}�Z�O)�m��yh�Z"֥�kZִu�B�(ΰ^chpn"42�P�T6�� ������u�JTQ]�4l��F�ac0�������pTs 8����s/��FK���	�Lk$x
:�/���e�Y�^�~$$K���8O�XYϡ�ݮ�߷pd8hs���Ň=>=G�(V[tuw��T�g�a�3�
���e.9W��Z]8m2"�8���n>[��"��:(L�Z�ޜ�e�]+�{ 3A���D�+#��\�tB͇�Z8���G�Du�ya�iDueH��H�����)M���DuDDDDm�"8���DDB"<�)H�)�H����"4�#(��#��<�"<�8��FDG�GDFQDDm�"#,�L"""""""4��.8�hDFYeDa�]im�YuZ�e
-l:���6�#�G�B��"8����R��8�-k[�Zֈ�"#l�������V�8���8���0�FG��F�H�6����Y�s��l�tڣ&*Ƚ>�ss���:�D�f��4�I�r�l��A �6M�ڌY"��a�&���=���9$�f���q4C#LRJ�7�T'��3י��4�7�������ǯ��ɘ��"&-�V����okF�3��,��6�g3�S�Z"2f^M�6!�O�M�"Y6;�G�o?�o^�fw�����Ce��ܧɓ,nEm��5�4�X5��u���,
���%�in}6t�3�5~�W��9L�/,�-6��������]3���7���k�����W~9b�f��%�Nf�MNJr�ꢗ���8_]����э�L~�~k��$�
�ǟ�-v�py�̽(O�3�{�f�s��������39�U���Í��;�긎�W����� T&\�no1��q�&�œ��Y�>�V�h�F���X��^W�^b�&�s%yd����tx�Ѧ�f88�1g���s��Al��PVl��R�rf��2V����_W��[�,��앮\k��5r�|�]����:�B��(��,*
�Z�FM�ͷ9�s��f�RSMj6u���@�JM(ˮ!H�L��bm�(U�GMc�&�8r�^�`]qfm1JT.�p�ЗNJD7k=�d���]��KMF���m��W�uI�,��+�3k*��([�i\ �]U�m�j��}VR��|�GGZܦ���U�"e�u��%@�R�rn�㔒�VA�ɜ~礓�UW������^$�I�*���s�������'d��_��skZ�ڔ��Z�KDZԵ�kE�q�Ye����韾�\2�."��9�&̪�j^��:5*����mH�SM5t��e�v��4�iE��E�m-�YkLZ�/`���b��k��X7[T츢�qv]*�ڍض�m�0]�f��-���2X�]mƛU��1Ke�4����PʶѲ�n!ve ��]����16�n�Ѝk����5�X�lX	p���"���2�K�]5ׯl��.�l�Km���ؠ��Y��ip�Z�˲��6�*&8���gn��l�9���8��N��T�w'ύ�Y�;;��T�f�2�����dͷ#�h���`�j=��x�-o1���^���ꓡn���x�xf��
����h�"�H��b<@��M������^4a�#o����u~~�;��}�����OEF����}�+kF���b�e��P�J*�gƶ�7�#�F��U4�����$����F;0uf+Ș�?�lF|+TM߭�����ptN�( ��m8~{:�Q���:�)Ǒ�h���-kZ���MYBa���I������n���}c-�4��!>L��z���Cͤ Q�y=$�g.\�L��1�����O���7�OR��l��\MQ�^�E�v�g����Z���|�������~���}c�V��:���6����M3�Ǔ�.#�2I�'f�[��[![߰����P�P鏲FYg(GL,4oE�P�t��c|l�CL��G�8���?"<�E�KZִZ��!C0�h�cj��cchg�qt�oGֺPO���*�n���:e��SU�����>��>�ի����c�G6�0ĶC�;�����-�_�������rbqG]�' 卺�;6o�
<h��N.}Ӆ*�Lu*R8g�-�B��Kb�����8�zv�G�j��W�	U����[�mҢ0�l��J�(cogEE�u��k���uǔ��ȏ-kRֵ��t��B�)C'\D�6����AW�cchc5�������N\���)`�q&m^�G�_*G)��t�0ҏ�&D�$ܰ�ˠ��VT��X�{~'̤��{�h�i�dPmiY�̓T֘i�3]ߪI:2��YR��ѥ��oǸ>�f�X��,,�2�8�:��-�s�ƌ>�I�������ܳ���p�sa��2�tx�e�I������,�o^�t�fDL(�!�r�>�rQ�{����u��q�8��<���Z-jZ֋Z֎��,�ˎ8ҽ3��ư.�1�6J@L�t*���; �]J4j\�B�c�}����'m���WZ�ػ��6��g]��	�h*s,q��Q�p@��/�.MpS�o	&>d9����qW��]��멣�Cq?����$(�cN=�..e�R���͹y���c���Y6���ZEf~[�9�Z�6�,��cy�-#[;^4l{�&��1�͌fwMC�c���3�VPxk�:i8p�y������US<6��Cn��^4������(!��of��;O�*�I�脚Z�e<Dq!�wc��>�W�ct��7-�4�t�����#�Q�.&��s�5��Ka���C��j>h�V��3"8��#��-E)jZև�<tх��!�Q���6&A�8K�(�7M����66�}�Ҏ4|YM��VB��QN��˕R�����!�>�UU���3�J�YkF����ƒ0�B��g�M�@���Q��O��L��6��ZL���mY�����tP2��j��I+�p,VA������e�	�L�l���l��>��񡿏�,�4loR7��s��ѝw�l����gR�`�;���/�1������<�<�<�:�<�q�E�kZ-o-q�Ye�aG�3��i��y�`�'��l�=#���v}��~��8ap"8;f��������KE�+��n�`�kk��0á� ��M�Q��ͥ"ir�n@ŢxޟSʁ���s�%�l�Շ�Uc��V/�A�Q���dV��CVp(Ό!�4�M�3Ag "�ϛlld�״=�l`�����gL
>Y����q�Ѱme>�-'�~_�>ۿs�~i���~[��uռ���R���h���h��B�(��Lo}%6����2V��lQ�(s�Q��*W�8�!�C�pP����~^|��:���n#�����F-�GZ��'p�1�U��<B/(Q���B�$�k��:ƕ���M�#	���D�?��Ã�]n
���UU��e�7��X���޸?h�6:P���׹�����P��>��#Ƒ�D{�\0ß皒Yf�����QY�U7f��y��Z�E)�kE�՘t��!a�y�I�%���b��/���G�[����p��b���e�ش�ESxOz�h�$�b��n�]A�erGj�;#m�̵�(T�v��.�tUk���V��W���H[�����>�S,��]ܩ�b�7���d�:����F�iϟ9?6ǆ�/b}źw9�w�7���7�}=�η�\��U��3M�L7�ݙŁ��d��ѐ��r�27>V||q��#�_��1������ |YD>Zn�ɓ�����O�%派a�֟�G��ٱ���)W���>43<s�n��iil 3ɭ�p���#1o��U)���
!j��|i��
(e���mi�(���T@F��U�rQGl�.�Y�iyCj��P6�Z���v8��m�:�<�q�G����V�8�L�ˎ2�/c���1�jkm�0�IRg����Q}��̪���j�n���p�|""{(�a	�>DV��L�U�I�;�R�^՚���۳�^ǲY�m9O�Ų��Rb�[�GZ���xx�����h�gK,z<ۤo��ւם�n�DTq���~�4�/���Y��ey�3��*��i����I�|.�f�&�wu%Pp����X�k��� ��m(�5w���p���>�:�庥���""2�"2�����6��F�GQH�"2��"4󮺏<�""0��DR"""�FQDDDDDDa
R")�(��":��"#-"8��#�)��F�B��"":�����"4�:��QDi�P����������8�hDFYq�D�BYe�ܐL�tAKi
-l-KmjqŢ2�G�B�"#���ԥ)JuJZֲ�Zֈ��G�Dmkeo-�8�������#,"0��<�"6�Dy�Ђ'��vl���*��sܾ�|T�C�V�6rf��B���sd�ݾu�y��,{�����m�6����[;�|[:h��C�9�)o2�7;��L���yؽ��y6��gyZ�y��Ʊ�}��Ў6T�1�Hy��C��}�,]6q�k��kM.���H���i��H5�3^�W����[�ٻ�Ƅ~��ks&;����u���~w�������*���z��s�wwI$��Uk�9�-k[�:��-E)�kE�ո�6��C,��`���,a�ݾ6��NB�;�UUFϾ�D[8Z<��C��^>���2�1�Z^L<iX���RnN�S�T7Ye��[[��X �4�m.��/�3CV˺����DZ�QE�}
65�!g�h��8k��|��!�g�G�>(!��{m�87	)�˩$Li.V�4x a��x�niXsln-,!(}t(d6C�~3�}����y�帊R#��Z�kun#���,��.�ؼ�cZ���sM���{���smϋ(΍P�5�n��Xh��u&W���r�֊���Ӯ�Y_��w�*.��^k{o���(^E���5�6�x���}�,mЈ�Ƅc(62�t���cm�J���ߩ��B�w�?N�(�*��لR��A�Kd4�Ǖ����0~S�o��)��O�3��庥��y��q�G��kE�Ÿ�UD�Mb��'���_�U�S��*��G\4��?�&BW?5��V�����<R�ֲ�JF�3KS\9!�\f����u��@͌.]��ԙ�1����z��e'�.b�^� ��77�ڵa�Bծ`�#>m�fs$��$����G�����󕶦Q����r�bv@p"�a�bcŎ���I��OF��j���D�[3V�����yu[�wm�[mBJԲtA����]���,�6���,�2�3
]^
�͒�RW�x��
�>���N8���F�s�`���n<m���=���,^�~,�J,iC\��OR�F�ԅu��v�[�e%(*����N����Qѡ��63���>9'c)f���6�?#�<��6�R#ȵ���8�L�ˎ2���!s��%M�nQBE�����6�u5ůYhٔނ�g�R�M�}fi�1�ᦷ��7'ˊu���������|V!��L!F)�����7����ϔMtݞu��7�3�i��b��y
{�-2lb|v���l��Ԏ�����v����QDq�V�i(p：~��7a.ˣ����~��d; x�]��cO;Ԧ2��W�f���#έ�yH�)H�"ִZ�[���!a�.:�"x���`�P���Iwm������e6S���a��A��a��H��-.��׆w���$%U:���|���0�ыĹ�����1G�R�HF�]1��e��n�,�4mDl��~B�uD]{1l6��)X������kK0e/�M�D�S}��T\��t��eAn�N�������2�agA�5ű�4W��GH���y�R�E�h��<a�(�!�`ٮ�9��l���nB��.���4��5�����6ܪg�	>��}+��[(��[��v���r��qb�|0�k����m���6C����i��&u	�Phm;~��Zi$���oΤ*CH���Ϣ�t��������m�#�q���ے��}G����׍�MꇤY���ncc�tц�=�Z�՜�m�\m�)o<����)H�"-h�����e�\q�1�^�GS�l�Go������J,��QL�#����R����6�$�JEQ*F�	qD]c л��մ��X���Km�����\��ل^�V-q3�[֦m�k ����NW���n{/�G��8<xw8c��,���yyv7�8�x�K��L����S"���s��rq�3uʳ���E�Q$ҥ��oagV�*=�̟��\8 �4l��H�2�`z�6`�Y���f��{ I\!zZ'���.������t�6��
Ms*8YK���ѭ�P��ʭ���%t�*��W��"�X����D�k��6눖*���
�a�o�˘7��8���F��x��`�0�L�q�3�S�#�8��y�Z6�R#Ȉ�Z�[��m2ˍ8��o��1�`2�hgl,񭛐����Z6�{��+5��N��G�Ŝ�"�,(���I�{>�QM��X��AD�V�cN}��+��x���ޡ���I����%YU������[r'�L�U�5jj}�~�.��Ͼ�0�����}!;M�-1�l(��,�ѭ>�zA���I��ȳ�Ə#�<�ȶ�JDy�����YD!�3�7���[ci��i��3^"a\n��!~o\�,��)ʥ��=7
\Y�D�ؐc@|�w���9~�b��߀�%�3kS���x�Y�4����p�l��Y�#�zQ�P�ђUd�i��mr�ˤ�&��G�\:h0KTQ�6㏭�Ë��2���CIiY�`�Mh״UT~�nJe"�8_��@�q�uR�[{2������Th�})&���Zo͍��Et�<��-m"���")��YD!�3�;m�QM���/U�����������?��Þ[6��6���F[�>jIn�ݺ�J\��k+����^u�.[��|�=�x��x|��`����>9߽�IWDEG���b�J�)bݷ��a�|NDt��͘61��'�$D��G����������|]4|��m4l>e�3HZ=���͢����>��pѥ���ݔCc0��[H��DF����mF��:�"#�""��DeDe�]u�y�DDDi�˨���#��4����DDDF�SJDuuN0���"<��"2����")�"<��BDDGQDDi�q�2�m4��)�DDqmqƑDi�P�De�i�QFQ�B#O4��Է�8���Dy�!B"#����R��)�-h�����"<��"4�#�#ȶ��[�mŶ˦�Y�FDa�<P��� �&7�Sٜ�+j��(`��&;w7F��nZ���Y�s�Z���R�O�g�����pj�L��g�'+�d�����k\�U��2f�*�o�Ŝ�����e+�p�7t����1�J����(���_?=���>s:��XCr��rd��5�c�^��P��Y����}��NfG���;�߯D�J�F� ��ęҕ�
l��՞��8��̐�����Y ��ޫ�����vm{���^�q�2TC�x�~/�r���}&�܉�Yd� �Z�mڛ������z�]�;��Q�X@M�L�Z���lF}�&
�c��c?��>}�BN2��Q=n�rFW%O�i�ϳ'�'Uq�>Ǧ7.��8sY�"irY�&w��'c����7ǭ��R��s�b�B�n߱��9u��;����2-o�w7}���:o�\.�sr-�w�@ղ�j��M��(�.17���{��1�٪b�AE�Qp"ZmKv��]G;I��fT�a.��fb�Z�n����|�B����9f��Kf�]�3Ͷ[l%8u����ac-�[��v�U6���xt��;R��k���X�]�5��W�"b�CL�TPa�9%��ն#=��$��m[iP�3i͆���]���	y��q�ʛM��a������5�g������ު��Ҫ�������ĒI'�U]��7wwv���OJ���y�m�ֵ�JyמZ�E)�DR-l-�q��eƜa�N��u�c�ε����2����v%��6-�]��1l�%��Ks��)1P;6�!#�9`�SSF��㉙W96�p��[��5����J�E���XT|6���([D�|�Y<�+��r�[�5�jGG8�[���)69�=K�WMpmb����ڤ�Kè�b�	lcɋK�u��QM]���ڡ��Ze-�l�.�l
P�Ce� ��0��UWi�f�Xͦ(LU#�"����3kY��o���Y�3��:�M�=3El�*`�3e9��<B��Fk�.��1�� ����:��e��m����w���vY���g��yo��f�h�t�M�o�[�q����e����nfG���<��p����$� s�i?!��UW{\[7C�;�Y�o�F���S���t�T���~�2�[���у��m��x}��{�Y�Q%�s�ƶ݌���tlk�XN�5m�uUu\`�i�&Q;��.�2�!K�8m>������*�U��mt���j�Æ�(9�uU߼%W��F��
딒+����5՛M5��
י�8EG�����σx�W��m�=��1Ƒ��q��]y�F�JDy�[qm�Yq�wLc����*֛m�:�P�aF�k��Ԫ��������p(�����r:�g��<rG;���gN6�4۱��-�C�I9��1hуv+5e��Kq�$= �窆6۲]6P��%��=���b�~k��{���{-t�g�>���QB�o���K���XI��>Qx�m��:���>�UUS��'��f�?:���u���)H�""��c<aY(��T��6ci6��[m�f�$��c]27���S7�����h�c9��|J18l�3HL`�)X�,�ŁE��=� Wf�\�5uc2!^Z&���s+P�u_�����1�:�4-�Ê6hpf�߅�~4l�e�P�����nrS����$�)?O�-'�g�I'�����撰�;���~,ٰ�5�X8a���hg�����<�i�G�H���2�YE��
m��Q�����m����k')��9*J�t��WA��|R��>E}�v^3<	����0�
��Ek��b�6����.ߛ�C,�E��Ŗ��F쳻m�x��ͭ� C�^Gf�f�gw���$����ٳcbc[�_H�"�7��MV�&uR�ow��9������:��W�a��:�>����yמ~F�JDy�[q�5TUyF���n|�?�L�%�Et�S�e��J��Y�$�cA��~/F�B{�m�@�lȪ��)��--(�|�x�����A�6+�f�mT1�(�LU�qr�6�Jl���Z�~�Yr.�B^�d����뼓sg3��pm`���3s����3���Ry��p*6��>��Yȋc߆a�U������7�{��.f+����t����DJͮ/�
���}��6p���W�p,�������ç��)>��o~|��|����g9z|�ٸǍ��2�qI�m��\Y��X��[Vo�"�cXF���V|Y�!nqztV|(��cT��	�$���wU#y��s�������
546�鯜�&R�ޖ��l��u�E)�DR-ke���Qc;^�Ʈ�m�:w�Fͫ4l�{�M�+F��p(��D)2����u%>7�~����E*ag��4�ݷ��އ�	�Ɩ����W�W7d}�FX���}U�[��*�>
4a�������>}ٖre߱�ԍw�g���e��S��`3�N8���k�8ql���>4[�κ�E)DDR-ke�d,��Z�i����"<46�L�ƛH� �T�lsҏ=���eWe���ӷ"Ѱ�xч�4�D�kX�m�X��X6R�ey����}m��܃q����Y�}���~���jb�Q<��DJZ�Uݔxن��eV��ь�͒��2����ߓ�Xt����(p�ņ�h�x>�pf�m����5m�6�"ƺC� Y䖎p�dw_y�8�+�h������هM�Rߞuן��)H�""�k[&e����ȃ�$��f��3~���9UWW^<>�������)a��0>�lz �>���)?��62�h�u�f0o�3��OU�����ZK��:����\a��?�l��֜�����0�Spkd48g�Y^�R�������I��Ap�m��)A�ō���U�ѽL�8p�+��������-�h,��˪u*�CcM;�]k���
�|��h��u�-�R��DE"ֶ\a��UEP��՝�G�7&d��7Z��>`cx�I��ٟ�Ң�fV�GI�6I������q�����يX�F41��'�֛�뛛cH�"5�*d��f4LX�YqmbShlhcmØfs�B�>���]���Ym��LϙjL�*�Srn�5�~d�Rd�W�?���YEƳ�{3hE(�0�0x�����U��f�b�����X��7�\7�r�C�,�����Ѯ����@�3���6��D_lR,�c8�\O��� G�{_GD�����ܓ��'>���d����#wn���%��i���@��:_HJ�⿵s���KT��P�1�ʩk���[��\�G_�L�*���v[xh��T��40g���7�Ϙ܌�sE����G�)��uז�QJGQ�<C2�YE���a
�6��爡�9���3���'#�Cu�6�l�Ɗn�(��t.F�f)R��,�'j�����4-s��e�7��_�7ӥ�b��PT|�����"�w�_.��bn76�n2RFW~���Z���-��B�F/����Eҍ��3Hmae��Y+�� ��YP��6�l�(bҖ8mbc��k�0|�%U>K$�}����cgﰵ#.)�l-�DDm��""<�#͡qFGQGXq�GQ��y�Q��B#h�""6����H���<���8�"6���
GYDF��FQ�mDyO)�FB��""'����""6���""4Ӎ���#����ӊDDm�q�DaaDa�i�QqFXy�O4�E�Z:�ֵ�h�HB:�DDE#y�)JS�ZԵ�����":�aDq�uGT�m�u�ʍ,��[(�"6��M(NA��I�\��,7�9\����5��8T�e5� �0�3����l�4Ό4h.������2�l|���Y1q��;�ֿs���?_ֺ��g�����N=�mY92�q���m���9��cCo켶?�I�(��SlkBl�jV�NG��X��E5��\a�%����VF�4!�Ĝ��V��
Ѧ�Tf~Wy�6^��BU`�]�v_��x~{ʫUU���s�]�ݮ��UU]�<�.���$�IUUw����Z���<��[(�#���DZ�q�m��a�c�yU,�죆�{m�4��h��e6�l�gv��;�㚺d$�62(gq�[[!gG�3��Rj���&�u���!3>vK�豗*����ͦ�.C��ݼt����q�?�κ��m�H�ϕ�:5�p�V��3A[�{,yE���#%�)+ �6���#k�}:�u�(������μ���)D舉���!��,��FF�m�[����M�B�8�{�Qh�}n��5�.|mӎJ�v���lQ�l` �v,��TT�gHp������d�rt��f����8 Aj�"��S��+8Vު�T�T��M���>~�p�у_&c⥨3E�ˑ���5遡�KD<|@Ѓm%���E���Q�=$���N�Q��m��>��ɴF���}��0��}��-o?"<�?-�R��DDDZ�b�UU	v�ϲ�6��|`�I�l�#f���\�P���^e���m�ɕ�^�+��	1�c��ԅ���@�"��ї\��`ڦf�Bc�̅m╮��um��Sd��s� $w��Ӻw�x��Y�Tʙ^�Ӗ���m5s���{���\�f�Hn�i��(*�I��z��v�~)o��v�SRcD��}��Ɉa���V5�o(�[��ЩQ�}:��4sÈ�r�hk�p4�e}$�����Xx�¶�S�t��G�|=C4�ϽR�g�Ѱ��"��ӧ�ôy|pe.��=�8��bᅞV^��X����Y�{�yC��*�k�CZ�p��9���KC�W�?(�#>�0�a�2�}>+O��*����[�V�M����:���(�#�����ǆ`�aeX�m���7=ٛ�$��8`����\	��l�k�82�|P����A���M&Q������G��oU*B�WF7E�K���J('�ݳ�l��4�yr�Qj�U���`���V��ê��Yi]���S,#ib\R�f����^��.��m�͗���S��6�����(XCg16�)U$��y�],Q �&_^j�s�x�#�)��8�V�y�^Z2�R:����[0Í��n��3X�CkM���C��,�7��D�M�8/�,��7㨬V�q���6����8����ﵗr�-�qy��ߺ�5��~wY]j���C,���n؊�:ܶd�&V\]@���1�h���!��9�A�|0v�_Pѫ�s,4o�{��(��nC]����Y�}�ٴ�zb�<Yҍ,�j�����i�\����>8����yh�)H�"""-c0c0��,tu�6��i�t�l+��Ze+c{KQ��A�f��aP/Ÿ�������&9.e[&E �}FݥN��ܩ�����V��mm:���&�r9(�bم��P[!��cǨ��Â���a�m��#��[rh,�(4pn�N7�5��5ej�ꜩ4�4t�QC"{4p�\�%� Ca��a�����Y���M��i�D��[bM��(ҡ�YAG�R��<��FQJGQ��/���QEW=ӝ�G� ���BT�Z��A\+��6IQ|V44dƛLMV[�T�̴q_����3�3�i�4�t+�lq
}-�m����1�A�����U�
�-�(��L�w�W�gDl��\d���fb��ڬY�~�z�|X.b����C�L�u��1�3���N�W�̊�&E�[�8�1�(5R��e�:`m�7�vb4���%S{�t�!d�Y���m����6N�u|V�)b�gil������D<3K�HQZ�Qa�ϼ������.��rxf�/-th�J�bD6�on1���K�3��?��㧊4�Z��n���H��)���ccYe��e���O�.� ۩�8��8�!��m�__�l�e�7Ɇq��G<S�4���V�y�QH�)H�"�<3C��Qc4!��� )�� �:���l:��C,ٖt�~�D��<~�ԏ���iA��~�#00�KD���{�����f��x�Þ�j�x3i�f�B�ھ��5�}��_i��w�7�dSi��c-N��E���*��)Zu��d���L0gG*F]kY��StG
(�����haθ22,6��|oD9��a��yhٳŇ.��Fꪔ�na*����Ͼw�k?g}N�J[ȴy�V�a�uH��[�Í��n|m������om�����x�sc�Mϻ�W	W��0�e|�)B1%c55$86��ֈp�AfȎ���cta�a�o(c���L���#���g�44}���@�Z���n6�W��|�q����󰪄p�6�t�â��~>��fc)�s����?7ͮ#�[oŃE��XY�Մ6�c͜��vꬽ���6a�k�
k�F���6�-�T��ujFJGQ����ɆQE�7����M2������l7��uR��8}\n_B�)peB��iw����[�P�Yh媪ȫ�QIj�c��4E%��ϟ����B.=c��G��6���x��m�ǋ82�Tq8X��Y���)�EQl��$'�齟3y���">8Yϧ߄,�t۲B��5�˹�6�T�qQ�=tP��tva���9)�xp�8B�E�A��1�v{�O]������w�iK+ꪕUF�l͇�����m�{������=��n�/<q��cn����ݻ����Ӷu���}��M#b�g���h�DX���h����E�����"�M��-�h�DX���"""�DD,���E�4["""Ȉ����h������"kmm�dDMD�dE���"�4Y�km4Y�""h��"�M�dH���h�",�h��"""�H�$Z�H���h�"!m�DDY,��"-��4X����$Mm��DE-��m�,���h��"-�E�ME�H��$[[i!D��h�"%��""",�������"h�mDDE��M"D�dM-���"�"""(��"��B""E��dDM�""[k""""E�4DD[[i"$Z$M$KmdY	D���[h��4DYD[k"Ȉ��dH�"-�""h�$DH�&����-�h�����[i&�DDD�-��"$YE��h�&��h���""�[DH�-�H��&�[I"[H�-�H��m"D��"Y"D��%�$K$H�H�X��$��$Kik5���i�4�qlsi%�i�4�E�%�$Ki$�,�H�,�,K$H��i�Ki4�d��5�$K$I����,�f�d�4��&�H�Y���D��H�I�Y��H��"Y"D�ki%�$�H�"�d�%�$K$H�C��	�m"D�I��M"Y"D��"K5�4�m$�m,I-��"Y"M,�$�"�4�D�d�$��E�id�m,�D��E�%��%�$H��II--�֒-YZ�&�-$�,�dD�$�Kmb$ZIm,��-"Z$Yf�[K$Ki%���m"D��&�H�,�M"Y"D��BY,�D�M$�d�im"�	m"M,��H�Kk5�4�D��I���kibD�m"BY"u͎�[I!,�H�Kk5��m"M,�,Kii��%�$Ki,�HH�D�E���D�E���DȒ�$�ZIdIi$Ki4�E��K$�K,�Y!-,�H��Y���i%���%��Y�KH�I,��i--$�kD�֒D�D�I��%�%�H��k4��KI$��%��Ii$�D�XZIh���K$�KY��I!-$�ZBK5�h�M-��I(qlq�K"%�%�ɶ[?ә��&5�c[&�l����l���gnv磤�,����ۘtf�Y��Y��[f�[6�Lke����l��c,r�����!a�m�Lh[2f�f��!fθ:�t�B�� ��	�����B�X�͡3BL���������4&��m�!6��ַ����Y&��PD-	B!i�d$-BBɲBА��$-BBɲM�Md�7�3�#-1�M[X�r-"2&�i4Mi��&��5��4�Mi�h��D�5��kMI�4�Mgmn4��5��LZi5��e��֍&�Zi���M	�4�Y4�i��Mb2�M4��M5��i���FI�4M4�Mi�i5�I��D�ki�h�D�FD�5�D�5��5�I��K��,�&��i��&��&��#"ki�k&��4Md�MhȚ��5�M5��4Mm4F[M	��&��i��i���2Mf�&���k&��ki�2�D��D�5�D�MYI���Zi5�D�5��Mm4Mm4�YD�FX�&�4�[M4�Md�Ml��kD�Mm4�[M4�Mbm#"ki���4M4��M5��2i��&��i����4Mdd�Dk&��ki���i�&��h�d�4Mm4&���"kM4�[M[M4�MmBki��ɦ�[M4�m5���&�ki��i��hȚɦ�[M[M4�MmX���Ț$[B"h�E��-�4M�4:�éLL�h�&�""h�"!1dB",��h�&�&&���"E�DY1dH�-�DE�"ɉ�d-�E�,�-"$Ym�,�DE�����""ȑ���&��ֈ�D�"�",B[kD�DB�"Ж9l�ȑhH�$-m�&���B�m�-�Bȑm	lZ$Y�![iБh�4k[BE�Y,���E�d$V�"B�4Z�ċF�E�"�-��"D�t�$!F��$Y$Y-m�BК,���h�mh�m��"DD�[iE�dH��H��ȑh�dH���,�BE��m�HZ!-�"��"h�,���"km#�ۅ�Y&��-���!"ЄYeۛ"Ț-�DE�4[D�Ћ"DD"h�"-�kmdD[DE�DYD��Ț,��dM�-�E�b,���",�����4[D�dDX���"�"$YD��[h�DE�d-�H���h�,��h�-��""�"-�4DC{i�h��\z�߿>۾󹳌��<��~V}�6�-f�$f٩&w��3����s�>�?��������t���������a'�'�����_��_�������ӫ9������ݸ��ϧ������O����ܾ-�÷���������?����?���u�g�m�����6f��_߷��<�:�����7�t�� ���~9���#r-������o�vF���}�}9x7���6|:����v�y����������|������lͅ�3�/����4���:���}�9�����o���5��gݞ������~����nn�o�����>�~Y�>�㯗g�����:Օ�g�^�����ׇ46f۟�c�1�l>p�6�۶70ٚ�e�l���[6bY��[m�[:�vs��p�s^�z��\�~���zχ�v�_��n��[�Zc65	1�zLBCl�&��	l�6������O�}�V�ٞ�Ǐ��o�o�zz>�|�o��������.����o�����񾟯"���s>������-����znޯ��>��������<|6���;c߻�Y��~�~w���V�vo��?��'�Ѿc����߃����������8ٛ�}�F���>��~�~_k�������s��^�C��;�a�w}�fl?�׿�mm�����?E�]�����u�n���������&�<c�7˛f�w۟MI��i���-�Ώi�l�s����}-�gs~��C�v�g�l��>����;wޝ���'Q���?m�|�g���?�z�ٛm�����_E�?��f���x����}?�ݟ�F��>{�c�|�t���������Ϟ�u��6{�+���߆��ϥ����}��c}�6}�?=��~-���|�흶l͇˙�g�����~?�������7��}�>���c�~�~��>/��>��������{m������l�������wq�v��n�|[���c�n�o�����_�5[���q�O�w��������j_�x3ag�_6�7�ñ�Ns>��7��&��7A�ݖ�t�6�7�����=�z���s�ñ�l������VϏ�>s� ��~]~q�緢l�O�w��F�|���s;g=�o�������/G3�}����?���ޟ�9�:��g��=?��?�rE8P��Վ