BZh91AY&SY�����߀`q���"� ����bH�|      ��$������ ٚ�+c*�ҚhV[[e� 6֪�j���5f͐ d����h�UJ�����S�د@h�J5�-�fض�Q�I6�F�!"Ձ�-��keQHP���Z+m����m������dUih4��ɥ�P��4�嬷�ުP��F�+�Up����׽ޡ^��[If�lڭ�dI���͖�ZȪ�U5�j�RURM��2��6�D[h�J%[k3UKV���7G�W�֢��`    \��T$.�6�%BN�R��.�u����mn�j�m�\��v���hӪ��j(�S���t:��V��ު`�E��ڭ�bت_   =�MSl�]�[��˰����I�M
)���{��Ka������Yi��[��OF�{�z*T��ݞyJ�;�/���������R���խ�j2i���� �[Y��  v�>�;�+GG���r�N��/1�Pw=>�Wo�����] ֔��7z
 �p}���P}�}�����c��P .+�4�v::�
6� )Jhֆ���֭�  _|�_Ow��<+N�m)^w�����v���ꗰ�[�� U:t���=.�M��;�y�K��GCu>�����{��O\z�Pz��P��)�$��(�(_  ���V�6���{�aҀ�S�zh�h;��
zӠ���:���+��Ӷo/{����փ]�^��vM�緛j5K;Ӽ4���w���J�`�MH�mM|�h>�|��Z>����tP{���h5B��.=S�s���֞����z���۴�t�� �A�z���@7�n�W`н�7�W����4���BR�V��� lɾ   ����
j��s��J��iǏ������Wu}�����h�]���<�4x{�Cw^w��[{m�J�e=� u뀣�8:)v��c2
��|  ǃ� ����uά ��I� �����u���w��j� G�  o]{� t�3K� q�J��h1�YJ��&�o��  ӽ��=�N4 �W�� �����ǝW�z��  ���= 8�����S��+�e�t�C��q���Y5@���R�   �� [*�] >�y& У�\���;�k�(�7��3׀ �\���7: r��h���    P  !��2�*�0  M0 �{!�R���  � L "y1
J���&�4 �  j��@��(      � ����������� ��2Q*{)�M2OS2 ��=L�����~��?g�J�����q��͊Ś��kqm�]ќ���:1���3ff͟�` *�T?x� ��?�?�Ȋ���@�����}O��j�截���-UW�|���0|	S����+��?���/_Ʉ�0���&a3	�ɜ�s)�L��0��̦e̓)�\�fS0���e&3�L�f2���&e3	�̳)�L�f0��̦a3	�0��̦a3)�L�f2��0���&a3	�L�f2�`�as	��f0���e3	�L�f0��̦a3��\�f0���&`s)�s�fS0��̦d3)�L�fg0��̦e3fRes+�\�)�s��f\�fC2�c0��̆`3!��f2�̆`�̆d3	�L�fC0�̹��d�̹�̆`3��f˘s�L���Ps"`A̢�.a̨9�2*�A\��Ts�aA��A&ȣ�s�aA�
9�2 �UL�	0&aÂ9�@̊9�2� �@s`Q�s �aT� ��0 �EL��
̊��0��D��@s
�eA̢��0�U�U3"�aT� 9�0�ȋ�3((�As�`Q���G2
�P0+�E� �+�@ʀfUʣ�Ds
�Ȇd̠��2*�D\���Qs �dI�S0��Q\ʋ�s �eÄ�� �$��s�s �e̢9�2��U�@ȀfBd̂f0��̄�	�L�f0���&d3	��f̳!��fC2��̆d3!�fs!��fS0���&a3	��0f09��`s�L�f	�2��&e3!�L�fS0��0̆ds�L�fS09�̙�a3�L��S2���&a̓)�L�fS0���&a3.be3	�L�8��-_�h E����sFk\۩P���8F��hU���J�{�B�T�
�7v�*ڄ��oDAe�w�DŰ($l�N30���M`nf��T�z���^l���&����aܩGx��H�-H������jS��< �QoH��mjoA+f�'B��x�,;��O.řhֻH*�rG�m��t�k5(�۹����A�n�n�T�qQ�(B7u�J	��6�Lݥ�a�Z�ZS*,�7,Vw�%B�¼���bìeJ��Cښ.�"�/Fa�YDP��&�y�!.'4[$����j���Z�a'5�!�)�m1�kO�Sj�8Q�̛���r�>꼕2R"��bǴ��3�������nl�sUhb�I�)yF��՗d�S+�I����2�Fȃ�2��;���Q[m��b�;�xعC �o��;�j����\:<:c`��wSF���#���O�ɾǩ>�=�R�j�h��IwOe�Btmnਗ਼ ����+Y��QN�ˣ���� ��f�ُp���2����ɛf�6�d���M�f�B�$u�ttY�m�С-,�7Yطk=�]-zto�*H�I��ʎm�������a��^P% F�PI˚�@+\m�+D��PZ�r��7Vꛔ���j�ML��� �b&��t �GekX�;��т�nՋW�0�4��Ʊ��R���LilD|+0�1��f�h����Q��J�s2�l��5;Վe���;��4�v� �U�/pf�nF�=�̍���YCZ��mx�D3�9��f�P�[��LIX��"nP5�f9o{��t�)��I&�v��4�c�[���ԙi��Z��
m��C��[�gV�'�Ŋ�fm4i���T�h�ņ�W��mْ�ǚ/a$��&�V�j-�;h���'k^�n�M�İTT)��nm�s/{O*D3w1���Xp�E�t�2&^ē�r�WSH�j���8u��hsi�V0�C6�����Ҝ~u�l�e��QC�-�u��3*L������:��:P���̼NC�1N�m�2rf��r�Z���=�#���wv�R�F; m��]Cl���0�h&6�M��0D�+u�Ƀ.�ȝܖ��1M�L���;[l�`�܊`�}��L�W<r�E���{n�Q�`*L9";���gqP��m0�U�}��ͭ�p1��]k4�x2L-p�2�,�!)FQ�X��łV��1�]���(�
���
����!��P���<���E�(f�V������\e�pl��qd����|�vx�6���bV�E�a�F�XsLf�g7wl�!�ӵ��F�K�^��z�S%�۠l�L�s��q=Q�p��<b�$�Lފ6��r#(j��y�YX�	t[�j���s�Z�m��Y�\n�Z�\�`�ۊ�35]e}n&d�a]od�����4QX0`����K-�6F������gqaђ�N����Fû�a�CfS�Vi'ma��$.��*T��`jb���ą1w%%��6����I8],�sq1b���ъ�mlT8�,iĤ�b�4��
��~�����̳�A���t޼��r��um �5,�8�!�75z&�C�,^IH��#���w��N�9X`OX��ŷ76�G��V���B�2��[1e�^
ӥ��<�Tu���S w�6wP{��v�2�\u�^ѶCY��%�3Sn���B�:T��U:��P�/r�I�jQ�
��vO)A�o�)Ҡi����j۳-���M�U��CX12-V ƬZ�S�6Y�;�qә�eȤ�V�Æ�jX�x ��V���ı@�f�E� ��l���M�{Cv��t��(K��z�D�:�G\�L�AS����[�N�"e���]��G7#YS,�N�}%���\�9�O���x�2�ȝ%X���\���ﲁuxS}���ZB�ѳ��n����i�Gv[%�B ���;,�S���[���N�Vz�+w0�YD[jHk�CJZhj&���/�-����x�����d�V�N���ʊ���"��Y�m&8�3��;���ʚb�2�V�/A���F�CeA���2��e�cADm�=�p���(O	�EE���E�9(ʻ���SZx�*߻]���7ɋы��,BHܻ:!"�65�n�6-b~�whdČ��ƮǕv��qBq��5�(��ܫIU���Fޭ\A�.e��J6=���zc�QJ"�Z³m��Z͍���<�}��$�׺3��%�)`��6ml[Lȶ&�S�
����q	�갔�E��LSI!d�Х�34P8�Z����k��W������Mೢ��i�P���j��cE��&n�����݆�".4�"P������yR��t��lS�Yjf�F�m n��ө����x�ţG%�m��eL��M<;Rn�5I��/1Ni�JtoP�b����,���͊�C����ښ:���%P��D��-^;�1�)���Z�QD`�(Wϫq��x�rZ�૖c؃���G�3AZ�`jPvۨ�i���Ԇ+��v�h�/E#A�AY�M��Z�u�l�h����ٛ��Vւ�����	��J8��4�5�#�*Ki��vkS�i!H�5]�� �5��7!)�@���y�����S���$\����SX�H�*�I�%2�ѧXȳ(f���oZ�SHU�eVS�鷵����!83.�,v�pf��w���1BK ��0��K-V��Xr�`����*���Tu	��	$2Hׄ�c*t�{��e�"["ͬ+s� <%$B�[����9����UՊ�!b'��KL65K2�<�n�mi�u��G�d��l���M���y�,B�/��Tt齭ڭ� i�-vD�`���؋+R��{w�n�(
,*������2�P��)�+v�F���gv��C[y���t���3
��jǙH�5���W.�94�/��[�
̴�Un$��<�(ڂ���d�]�U�({(Ӟl;t�T�ŧm��ƃ�(�̻�"��7i��u��ś(�J�*X8��flxժv�v];2���M]R���զf0qY@P�w_=as�l�ū �jO�'i�C2�^+1���đ��P���n,��j ��E��t��-t�*�2�F��I�㵑�,����p�o/r�;��÷@"4�u<VȮ��T[�ᛴ)�X����kE�ʒ�Z3,���4���1 �ݺqJ��	J�=f^�m������5c���ֵ�M���O/�Vn��p�bn�L��A�o��e��ʒ�S���% �CNXC���[&uy��M�j�nԼ�ܼuGbR����U��Qn���!r��m<o[�aڀfa��oFLJ����;���/+Sz#D�f�Ӕ,�3482�,���y%�׻*D7���h�h�뛪eK�ص f\�Y4��q�(S/2�.���,�Sq�-�w���-�S�ͧTn�ūr�MY ���M1S+%Vh6t7����uص�����E��@��猵*	aGiP���a�s�86���g|�֝�tbxU����.��TT;
�5�Ñ՚���t���(��ㄐ*��vJ��l<��Ùe�G5����Ẋ4Y��
f�J#G���!6��H�t�Gd��W��D�‬y�����z/
���։.�V��u�Z/Y��j�Y�ǵ�u��𬫚)�.i�4�S�[gr��Ro���DU�_
�'�9
s0뙩Jme�!��y%
�EXt�kB���f���m6i65㽏.�`fI����I��{6�r�Q�Uͥ��V:˺T��Itr���
7n�ͫ6$ʶ�N�efH��0+c��<"�^�x��\Վ"�:���Z:�+0�9�tӍB�Qn!�Y��1�[56-*�y�$yiQ�&/t�[���<5�M��.�u�oIX0�����UKRccn�V:D&-E�&+mn�y�tu���݊^U��W��ps7҅O���K벩f�d����t�f��ᙬg���F��L�m�*Mc�Ue�CfQ�)42d�GiՓ �l�ϵfj�g@1)����:���#oKA*Z�uT�l���7Y#5��hMp��!�4ࡋ�M8c4�0���Oui�ET�+��o��Ky�k7H�G�0^�Y�����o�v���c���j�����36��f����ۼ��]��X�nWm<@���~4���=��u�3��+.���Vi0�r��o�3Hu��Z�,�D$�ں�gc�9zo&��^�Q!b̈́:�D/l�6a�T��R=l��k)�����Z���N-Hv�E.m�x�_b9���OwS5�lm���nV��^�6���ĩL�`d��=@�4���B�j噗 'l��f��_�Z� CMh͊����6��.�0H0�ZET�n-���Lav��։��
���S7��Y.�ǹ����e����l��A�.�V	��y��{coa�6&0�yڼX-�ܕ��2�i�7
�d�CT���hǖajjijE!�CV������Dai��2�6������ek[��f��0loR5nO6^�Z�뵩�ZTh�L�2��CÐf�7��Ff�v h+�32���6���CC�����Kp��(C���B�NB���Yl��TF�nV�f���V��,�n��k��a���Vt�@�.���+^޲��)榱ɲ�5h�?M2�|�� �8��o�Z��(n4��C����p�\3�)���-��i�r���^��~S�)�V.Xj�D-��c���,e��T�ɑ[�����oikT#oC��2�6D�Q��a1<e=�x�d��i��)���Y�H�� s��E�pn�Qj��k�"����-8�n�x/un�{{P���R�	dݴ 8V��J8(��v��iW..^;*m�n�,;���	�ȭ��*�k�rx��ֻU-]��C	��H4�pi6F���$P�T��mq(����i��"\�vE�u�Ԑd��ĭ��8�kxTr���m��Y��dyN�RcA3upQ�;���U[�Wr+"f���V�)n��/�vijWYy�]�/;7@r��a������Y�̥�z����X*����{v�۱�92X����+Y����Z��Z�[�W|W^�٩�Y�VLa��Is�0��P�Nޛ��Ǚ�p�7s$����ơ�YY�v��
if!Oj3Z֩�L�M�%X9�M:S5�9�ؚ!�����~��tS5�XZɮ��,䌛�b�bY��\�Lc�RQ8oE�v�p��M:���S���̽�J��pG,;�+ksS��e㵝}���S(��S\Վ�<�����6�6��0]�p�z��8���W�[��̋P��jb���`��)�\�-�v��41OPw
�i��nj�7Q�Y�,#M�Q��qm��ĎlF�eku�-c܍$���:��� �i�ţv˽v7�|�4���=Z���h*��*��6G��Mv&ʓt'��nm]�	jI�%�w&�:J]����Q7x-	[����ƮS܈�.���a�&X�ɫl�[��+�;L��)�M���HF�T���%�J��u�GB��JJҙ[��N�\D-
c"AhL=��&��r��n8d{L�˱��lzj�3�z��WP�6�\{R*�iV����t\m�U�S &�L��T �嬵�������	N��^х�yX5�YD!��R�X�V��K"�p�Z�x�#N=`�~:pe]^��st̅�R�ݡ�T�5ב�U����+��%	s/W�llfOc�Z�����I�Z@�)U�7S5bN�Ď[E5Z6f�l#n��sS+n��ǵ"X�P��YS�j�
T���
1��e;HUͫ]�{1�XV*�Ӆ8)�Z.����m���y��Y�>����^7'�Z*�0�u��s���!բ[�ҏys�t�uESwl�k����������]�J=x�գ*��qX�P�E`��J܅���فQ���pGS8θt�z�4u�QZ]�%3�%fV[�d��̶�-��8ح�m��r�J1e�lK�'3���,�B��v�FM��W��䭷A��S�w0�!���m�i5yp���tZ(��"���z�M�D$�{�x^
I����,F��)�-��s )<��1m�M2r�݃yPZ�.UY0�X�׍����b����1�F��LE��	J�<���?M;��&	Yf�T*)*m�H�Y�V��Âr�����$ժ~�Ȱ��i�U6���4�Y���.̢�C�Kt�݋*�0����(/|�OZ���`Z��oZ�j9��)�#&ȥD�ѡ�R�,Di�"1] =(�ߴ/pr0�*ɛ�4��2���j��<;C�Hrr�A���.�Ng�]�j�҆�"�>eT?���Z�ة-�v��D��|�ȼ���"1���/��i����K�ic���1n�cj�,wB�.�A����t����H.�����@z��9�R�l�vLq#Z�ni�S
���� ����;C
�8�6ռ���T�<!�=d^�9��c6]z=�;g����w�+�����@lsQ��D	�h�n���t,�m]���Q��
��+Lk�<j�d�8����S��uw���G%�-�B�v^��.�E�G�iV�����XՂ���Ղ�c�©Zb�qs����J ��g���mb�� �u-X-�B��g,IQsUi�I^�i�x\-C�vn�˼4�n�\���@��wt������x{G�w�h�i�۹,��Ko��4��K`��<SQ�W���9w�=[�+��i������`Z��(�*�4q�@Ϥ*�]	�gp�L��4�
J�r^���-����������|���L/�!������Ko���Ԏ��*������܇&Ʒzݹ���f������0��ȥ�TJ�T�u/�nX`�.ӽ������ս44��!TN�Y���:�plY|zo]���� �K-9Wk8��m'\��D^���(g_d����6�����n�H������4�r[�r7uK�L��hn.!W�u=�,]J���V�\��a������դ��&��N"I��KCP�	�'sy�0J��e`;�m'C��z�é#tTP�& �g�5}1��5�O@�Ǝ
N;bf�/�
�L�Eѷ1�T�WΥ���Mӛa��lB��L�Kks,�3t��t�v��&w>G ���f�����A@�u�r/�@{�[����C�.��L���Jl�ŷ:����2KaL�(y��0���p��5
۔ĳٰM���g,ŉ٨�3��w����/k'+� �<��O(�ڑ�ݹ����vR�:��I\���:Q���U/S=a7Xt��B��,y%�b[�@=�c���&�f���"������\x�����X���)��o��ΰ��6z����˫�7�3��6P��@��[X'L�(Ǩkκq�_t��+h�l:�Zޤ�n��E�Ue���f���K�Wtz ��sy��af\�sNu�䔬s����;�Fºt��,ۼ \o�J�ر9��)�����iR�}c���%��i����׌�{��K0�m:�ǡ�U��ybx&qX6.��g%�&�%���YzOL���=��Z��BV���m*�����-��:D8p��|$C���.�~���H��z3��)=�\v �Pe��i����ɂD�jՄ9\��Lٴmg-�\�,�NL�k[W��z8.b���='A�5MJ�Y�ze��G.
p,��o���"x_+=�[��7�ð��0�O{����4�؁ه'Ѯ��]�6k��s*LÊ;G�7�B��*T�뷠lP�_L-�b����X��'�8���D�w>���X#�W(�u;e�ѡAN�b�����oFm<Y���� u�(�!�D�J�mm3�Cr�1�1hA�Μ�Ed����Ӈ��e-�2��uz��5f�3�h�ƾ�z�.��8(	�xČ��6��s���2�NS�,���������U�9m��[�u���i��Nڷ�XA�Sq��Hof�Jopqw�P����[�k.�n0f��u}��ij`hU��k)�|����0݂MrW�7;)%������Y��x�=����q�reV����[l��;U9��>=h��-�N���u��'�C�T�|@u��.�}5�jI
��e
HҶ���tѝ;v��v��q�z��8��l�hp�L�5M�v#��M�1��$ݮ��Qi�k�tĢ/�h��m�o�,.k���C�����V�f��lȀ��L~�7���lBIx�Nd��}5B��U��k8��;;������������7f��J�i��e�0���O{j���6��x�����S�F����O�[�k�g$��=K.�鷚��8�S�%�Ǽ�W���)��@M�Q��D�[ю:V�4a_>B�2���պ���^=p8�S���XtqqJ٬�t�Y
�pqޣ���z��([Ty��oQWP��Ý�w*��$��dii����XY��ol7�,4�&������Ń+�*2����k|�R� �n��E�twjAr�c�i.�΅�u����f�3o��g�t�.�D�ֆ��w�&�;j��mԵ��n*��U����;�\w4&o���u��xۙf�5�V��rop��S�2�ay��n��15�M��$�J4�>#�(dj
\��E%�����9�قjR[K�)��q��oB�w�*�y;fup櫺�G���UL0���^op�8Ü���G���(�'&�H��WK��p=LmwL�^����ʛ{!B�����],Ugu�1nB���v�%�Ä�Cz��sQ"s��iZ64�N-'�m*&�se���W*y]�'�0��:V�G#����n)��5�Y��Pc
@��e�aV���a�t7LU�;ӂ��t���q�>��{�3[����~�WR��$۳�X�!�y��ڴN������u��Q�٦�Tz���v���8�y��7+�:�,�$:�V����w��E����K�O ]���t�8w�q�5�����Y�lJ�>$���=�]lY8�|B9�UBvnqf=����Z�5�
�f��o�G��5�.�ߊo�δ�aITW�k���f�k>7[֦PnI*V����|j@�3-��.#�,�%���d�n1v�c!,�VR���84T�X5��l�|�H��]��Sk����Ǵ"�7��`�ݹB}k[J�n;�ڃumog7�k:#��2]��)/X+.�� ���7��g6��{k�ɜ�@ь�049�\��Zsm��Ĥ��M:�f���G+iQM魬nU���]e�y��Y������GV�
��-��I(=Ҩi����vq�;�T����9Gv�9It��#_GC*Q5x�-Z�=�;o��_I!;U���1���۰Uoa0b���ںN-x��\@>���H7�fu�#yT��.ݝ����wuXv>��U��n�z�6�i��@��6 �FF�I��C���R�F�om��n�;�!#�ٷ��I��`vd���z�ʎmJC$���)��N������exV�U$������T�k���K�6,�kJ�$f㸔�L3��yR������]�W`�&��"si�� ggh�&М�RWIk	�-�������4�o#"F`ַ7"�./w/�+W଼�N����ԭ�%�5�:��Y ����N��u�HK��ю���]{�w�^s�+L&�R��&�U�K�3�a=�wr��vod�s�lm�[Y�!Dw�0�I�A]��%���m�]-��2��{^�ܫ2�+�����<'�=�Ofx+���5=��j��������fgJ���1�[�R=���[�"�����ZV�b�}f�r��W�H�a0/kWs�}omrI��k�]&(ӟm[�m�ռ�ig#�D�v��.���;B�	��Sa�3����l��qŧ#]��i�Ǉ���F&;�uu��>���d��V�*;5�i��J�`y���^m@�,[�m��4[͆[0�ݭ1��$]�o)�Ρ8վH���=u�ݔ��B{l��V]�{�_��`����hp��X��Wm%h��/n�r٦�ę� �M����Ҍi��hv1/�t�eCo�E5ӊ�qecąj��sJ�ˮ��U�5��Ʉ'U׻���sU�N9/jN���X�,�{�ˬ��Q:~���^[@M\�u�e>��2�#pY78S� EPK�L�\�i��eٿ��BkJ��r�̲����/��4s�5·s��&�)`ښ���R�k�L:���&�@�Һ�R�^�%���a�Gp�n�WN�)�"�n���j�80B9q���	��4WR�̧L�,�m��f�����7�)�I�˻��� R��wQ��S��Vv�tf��Gygr��وd�vb3�-��W���h0�1}WyQ��H;Ih��x
ާ��ۋq������l�7*��Y�$�?�b`��[���r�j�,c�[o�.���1 �����=�iA��p̵f@��
�:�f�ldA�k`+A�[9�ƺ��x�%O);�`ٹ�.��ȶaZ�/qc�JaxP�y+��Z�!��$�4��5�l��Ji���
��r�{R����j������]ѮW"����[o��o�S#A�nR�S&��boSZ�.��'x���5ຝv������ � Np*�øy�ή�(R$��{��P�L�
�^�ьҳa(c'p�e�T�1���L�vE���M;�ܠ#6#�$��fı�� <V��N_Q��Ԯ�U�ϖ��˥c�o���		�[�q'�Ve�1;B�3���{·jv9Af�Y�J:Zh�-P��q�љ���j���p1�dӒ��ʹ�
����ծA�I�Q+x�z���Uv#	ۮj�j,,ov��3[���.�KƍLݬ5;���ܖv���1�v���#�Y���.��An��������O��P��m*�O�^�=�ɤ���{��
qh�}�>娽;1�5m��^v��y��$kD3-N�[{$�g��yw�q'X���WCu���h1���]�i�v_F��gf�`��v�Ӕ0�Q���N�a�h��ީ���7�D8O.���&ԑi�D����J:r��Ww��U3*��5m��Q����;�d��	�Zo4hK����в� �Z�e�;����+0k�plފ�i=��UߺYs�Nt�-[�^+�#%�P3@�l�9ܫH�2�F��ބ)i��f�b*�����n{�j	l�|~=�{gǶy�(�,�4��u�/pf �G�t��!m۬ƾ�[3;�KNR8�����2;u��(d�6�:k�� ^�ⰝI����R�e-j�h�p���v[����u�d��p��S.�'r��r�l����hq�mcΗ/&��|�;8�tT�²���%Դ��L���w��+�\�,��������Ci��YXN�WZ87	�센o��0D]~U�\��;S��K%�Ү��y�u;	Ni���4޲�;�r�݋a������#Ʋȅ��T�����Ll��gsJ,a�;B���(Լ}��]F�Ԓ 9�6�"�wsG��u�QѬG�'ӻ,-��u���r)�]�]�Y��y�c�ٕ��	9m+��*8��Sz^R�[��:�N���8���]�j�\�v�R��ʅ��������E;tu�r�Lԩ�\m���쳩�S�*:�:��ےs�	��y@��(o>�>y)��k��I�[MqJ��o J����rP�s��82^+��"����]8_e;���ݩр�Y� ����k����iW�Q�gkNز��a�rhB�l��F�ܡx�_Ly����_u)�S]J㰎�h��X�{�c��p��X���/�=Y�5 ;�4s��P����`�q�[�Q�j�#f i�[S�`��;�X(u9B�P���]�o^�8��1�Ɵ!]ɭ��QCX{�&�X	}���ْ�=�6�����c����6M���p {B��� ����7(b�"��[�ϙ� �t|��������MY���u3�os�W6��o%�]�c�J����Zcۚ��/w:���89iF�@�Cs*R0�ע�H�+��v�U3�^i��na��+�qF[)��|T�O�+�� ����U���{c�̥GN�;�+��N�F�-���<bVd��i���z��k���F��G/W�X	����S�=ˑ�$��VY��8����oϢǗ�5\�ӓ2a0d�}��e�����`X׺R���[���ڊK�Kղ�o
��o��}D�����C0v�}4��X0����r�=�e����LQ��n�L��I9]�GYH�b�N�-�M�X��3�}V#\�*��If����he�ͦ�����
iFE;����U���(m<�7w��r<�,�Z��Yw��R��n�$`�خ��	˺�zK�6�k)mr��7/f,s h�Ļ��r�`tyx�쭒�R��.y�P�co�U�3V�Tb�J���n������S���L\}�qذi�\D��e�D�:�וc)f-S�O 9�e���ʫ�o(J�=�Q	�5��X܂�.�d9�+a�\튕����n�{Ph�t'+!�*)Ж�J��ֹ�#Ӻ�ݻ9�q��K�d�m>pM5��bu1�k��ԹV��S�6��$���t�F����yn��Zz>���z�n���Z���&0����@_;���:�o6b��$<=�j�r�=��U�\�
}��·W�E�\ͱ�wa�ѡa�t��Li�1�g�������@�K�8U��^ݫ��k���QX��L@�؞��%<+�[|tE��Q��N=��w�w�A��Țt��0-��N���3���઎�h� �=<�,��>�\6��Ưv�Wi]˯CښE��n,r�j���1�/I��`��(2�ʝ�-fd�fp`XP�Ш�紳%3���ɏ����ne,jS���)$�e	�|VU�}�9�BQ�{�3:�ec��F�^.r���}��z[T�.Θq谛�<z�rE�n�J��oB���}6�[xtb(A��K�D��Ʋn#x���)��]�`1���׃�0f:��9l$^�KL5t��I�&�bם܆LgL�x9�l9k)`�.�������J+8���/�}�h'	�sG_i�\ٷG��ro��
g��쓗e���K�:�룃S�p�JG7�	m!]ٚXl��q���:��{��l�<�j��E9�/u�{�:���_��L{���6=�Q�fJ��ŭ�k"+ca����(KޕF�2SI�6���!U�j��U���#9����j�Cն�i�d4�%�= ��(�R�uy2& �^�waiI�T�@:5V9��Eߑ^B����<M1J��-����4��t&�M�S=��.�\˄`��(�i��B" ;�,)C�Y A���b��Ex,Q���3Q_�6��DjdP��D#g�U�WYn�b�6U<C�(N]��Kh X͍p�U��]�-2C9��0�FZX�)�橂�EVܿj18���l5�0Ǫ�]S��@Ֆ�ș�fj�T�*�Ɯ4� Q_�����Q���o���_�O�@�0`���?���G��/�����gߙ��/w��e^��PQ��;6�T��LU��w�Y�z��#�15�k��շ�����]��kr���j�@n���EwqOb��}up�\�⳦9��L��Hdu�����e���eZfu���Yм� ��.�5�Y6WFu�Ņ0p�=����z�w0oMمJͷ��;6��ڔ�^J����-��lU��(�<�b�s�1�泌	]sf;�b&d}Ύ9]u�7����D��&�^b�^�v�Ⱥ0U����<w5'��.Jh��SޮJ�S7�Sj��ݩ�P�i�L!����#��dU��`*��1�ē���ɹ��aV����bv~bv\�q]K�.�\v|�]�A�L�h�Υ�w�^7B�rtn��|��0�ż��>�دl��Tq�l�U�4���d�Í��p��g�|�\`��u4�m�Vզ:�� ��sK�E $�z�>�����p؟��]mN"-�[Od�Oq��.�8.-�]�-O���\/���]�P��\h�q�M�{U���Scj�R�Ce�QXc͹BEC��FH��>A^�q��ϥ�܂Ծ���.�,պ��BU����TV����m���f1�݊F�e��p�1����kF���ptc-�ċ�n]`p���0�����
Ya�),R�"��=TN��64��������ֶ��M������-����������-�������������M����[Ckkkkk[�~?������~?��~?�����~��馦������֖����v�����֦���������~?���~?������}���~6���������������6����������������}?��?������~߃��ϧ��_u�]�<$[�o���q�D )�SC��r﷘ƱLI�C�$7�{uf�!����K2��^���x��Cgb�,Z��ѪR��ZU�n%��mej}����Rt ��n��Kdb�ы��WN�8���5m[Z��WH��)Zv��>�J���j�e�zsx4��ُE����^��WR��F9�i����&�֠�i�rѷ��0!�8:B�Q�l��W0E�k���k��ĺ,}8�ZdV��;��K	�E��WR�r`�(wE|:4�핑Ά�p9������ ;)�3��� ����sw;�����;q��C�l���Qcf�o�]k�ܶ�f�[���c�h`�f���^.B����i�kx��qtj�٫��pR�(TC�e���P�cŲ�����0u�t^0��k
/m���B��m>PbRJ�x�(��A�hP¢�@�Υ]�o�Gt����I�э��w�8v��/,� M�5h��9[��Mz=áHR��TA��n���4��-NbŽɺz�E9��va`|F˱�]:���cJ V�7{9�g����e.*����k �A�0�ii���O&Xۤ�Z�2�s(���ʏ�
�q�*�ĉh:Λ���=7&���&�Ѫ�`$2f�[	:���o3'QŦ�m2^q��;��ֶv�����֦��~?������}�����~?�����?�������m���[[[[[Z[[[[Z[[[[[Z[[[[Z[[[[[[[Z���[[[[[kkkkkhmmmmmmmmkmmd�������~����������|~?������g����~?����~?������~?����~?������g����~?�����y��~?������[;.y���E�m캺��m����X������D��ax�͸�x�u�o��V��[�G�d.�W�[FS5�4����E7��'Y[������b#o ��\��Ӡ��l(��#neTm(8�b�I.`�ûkt�����U��:IS�
y�{��h�Μt�u�[PZ#��b{��v�Buz����#[6��"����$6�"�<U[�t�����+��W ��V��Ŏ�>�"b���c����%_�2l+�$3�j�=�o���b��I��K���G�6oYA%��]�<��sH
��n?n�i
��W]��g�h:�0Gс�qo���3]a�w�O��?*���H�ںl+�3��D�<䵽t��3��s��T���M]�m<��c�'\���nr0v�yҳ,�vf���f����Q��b&k��l���]�f֞����S���	F�,����4����6ٮ��w�!O�Ŕ��]X����^ʽ3�U�+0�y�&�t��81��6�2Z�`Zz�7z&s�.��WVU����'D�[��H��Q��W]�7�XX;��[��V�i]�U��l�b��3wk5܄*��G�ů��c{�5R��w,!�|�c��N��Ѯ�(�RTRW�f�J�ڙ�$v��ݑ�`uؽ@��K=|ﲔ 8�XI�� ��]i����^
���.!{æN��ɳvJ�B�|���y���dr�������U�tuKTu�Ż�e�3n�J!{c�:�F
�Y���C���f�"��Od)�k�+V�3�sA��<'z��`��,\=�C7��0h6�Ѵ��Ѥ�M�mAN�ĭ���ҽ�b��6��L��l7�Fhv]λ:ȫ%��R<Ѻ�ј�lZaS��r{FM����wZ;}坔�u8�"<+X���4d\��I��;�PX1s�(��2;fWkg(u�Y�k.E���Kz���zb����4�oqol�`,9�u�,�0�VfYi�p�+/z����;0LbԘFX�[��̈́�XF�c�:-����w"E���#T^e��FNZ�7�5����������ʷ���%��t�^�Kg�8f���7k�clZ;���3j٘0�����֟Gp���lnt��)��ЭZ��|��z+����զE��"�����sT�Ӌ�x(H�]�9���BP�
`�}��!>Ӧ��V�CK��U���[�yk�����ZYHWb\�������V5.i���t��K:F�����V��%mv�(�v�ob����I��8t���2J�# ��(3�����8���M)��;���29�J�^l8���KXm��Uۉ�s�.Y�a��:0���⮆�*za�E�$���Co*l���;����c��]U��$���8�H�Q���x��nƅ�f�t����U��ykxcI�F�z��]�
ٻ}�3�xb� ���Q���nRᓪ[���]m�4��*ו=��1dZU��p�y�.���o��!e�/J͝����u�7��2��ѥ0��M�۰�3�i�)���ru�Ao(9y��P �[}9������u��@O�Wu���Q*̎�]�rr���4�BL(�Z�q��vK��S�BM0��ک&\&ʭ6r�"��-��N��n�R�#���ҁ\�ekѶ��Cv@�Б�
Es�N�.���]6�.JX�呷�h�vֱ�e��[`�o0=��N5Թ�E�[����ʆ"���p_)1���Z*b�P�QXԷ4N沅y��|*"܇�Uk5��v�q{����5��V,,�C�& tS���,Ұ�b��\����MwI�]�,`J�S����L5|�!m�]�\S���Cl���S��5�Ac��H�:*�*��K��7e�r=�F��'��;�Au"�W��6C&�02�S��Y�/Z��Z�7�&k�Kr�-�Q�X���Ͳ����]�\4�����F�w6;{��x4����6����ޏ�B��1ޓ�{(��m�0�.��5�)�7ywxV��:����b�f+�]%X�6j�'�Ht�@�+v�XpU��}�Mn�y;��JyLԮ�Ŏ8y���	�fAo��Ζ$��9�`*��n.!�SW<9g��V��5b땥qqr���	r7��}�t���wPt�eDgb�mr��Yp��v�$D���:kr*&Iż̜/t��+T[�q�l]�1D�ͧ�Z�J�fq��&���'n��ʅ+9�i��x2Ŧ�ȔJ���뫙[�y�XJ���,�����Ŝi�R<��Gt��K��� <�ւ�yת� ��� W���u�i�{Acer�]������FV�5��Kqv���/R�����xB�Vs����m�5�㼤X�" �x^M�M�<�D��K�2��;-��2��N�[ǎM] �.��5�3�/g,"'q��E�:�M�}�7���>4\�H��;0DNu�f��dʓQ��I�^�pU�}A�dwݍΖ���G���p��ņK��@�lǱ2�ݍ�v��<���Z̒�d[fbw���H͡��Y [�	�ASo����7�aӠ�
�7^�C[v�<�Ղ�c�[����;��MTx�s�YyN�vL�}� b��q�3v�Q�ݧo���ir'��Ą)�H{שDs)_M4���.4s*�]�X�",D:��k�ع�mJ��]l��!�����[���]�]Uk%˓>W�w���cAD:�8q�omb�C.�25���@�ݒ���a����kR�;�kY�b�i��W|�;�g�6�+��i-Zp���&��.�g&���r%�u{\�'4�YIRM��76�:�^Wm�^J��p���	��w�::{���(į6�n�K\�!Ey��2��'P��/��t_�������]���س��Y:�ݷ��.���.����`��}&��nh�;��t���v	91ۉ���Dy����Κ�i�EJ�c�Y���n�GUm�d�Ƭ�W�p�	]���T�g_+ש�f�8�r��^�t����*�r��b��e�f���e�m�=���7��h1*K�ZB����@���lʒ!|�G����Z�܁f�Ƶ�=��F͍�ݚ�h\�f,Ko	���@*��}r�F����PhO�-؍]c�N�IZ�(�x�Cy�����C�rek9�H�e�]�q�w�Js��B��zµ,�n�M��ʺ�Uf��A<S��ۙ%И&�ĖU��o�+=̛̈́g��B�7ČY �I���,i��f��2�4�q:#"�pfҭ�Czs�Y��Z�m��v�c���ֱ��̖�ve�D���ۜ�F�R�����j=��8ɽwϾ���[b^�5z�$�ޝ]ǆ�5�+0j9�Z����P�[.��	�mY��GM\*�`�҂��)�I���X���l:=��A��v�KJ]ޙo��_X�k1�5�@7��CC�4[w��M@���V1C~�ГV�b������=�-jX�Q:��\>��p�-aV���Swc8�z�'FAJ�nhwwO9�E�:�Q򝺷V�[B+��0w`��n���M��lճ4kn`�jn�.V�ss�,<�/o��A�-6�[.��=i`�skr�Z��ݗHn�9|vmGb��'�Di�`���A;��Wmd�c�̬"�F�K���ѐ��w���X��l6L���R�Ho�Ɯ�����Q�C�e�˸jd�����p��ّ{�Ͷ�=�n��S'Il6����yҳ^S�&�$�����T�<ؚ��1oy�w57�YM��IZ���!��q�73��N֚�s4�Px�}��?�Ǹ��ޡ0���&��+U��3.]e�t�jӁḬ0�Yh'���ǻp'����ƙ���R�{�	�������Z�m¸��Ӎ0�h�ddOK��RY��;�4��/k%�pO��݆0�.��y�l�>(��ż��X�5���=ݼ��R�7��vv=u��%[��$Vމ�(Q�[�����h|�M����<�q�F��b/��-���U����^Tƞ΄��N��H���q��Sj�Ђ����"�L�M��������VS�(Ĳ�L��ܥ���<�痴-��%��dX@�nE�>�2� (lõ��8���ǔ�V��6�UɴO���
�e���,:��޸X4;���p�ܷ7p�Ix�K�a�mA}`�>�Ba��U�uy�U�޼:dLi�DH��ad"�$�MVpl�zwh�r��r�t���']qH��_m�t�}�t��da�Ӑ���;/Q�����)
V,Xo�{�U���.�7�2�6�Mۏ I:�蜺��C.�����0�ssGL!Oh� ���؛����n��TlpU�_YP,W�sU�+��dZ�I�.� xzg�k��*�̽�}�ˬ�c�ygwG
1B�s���Ņk��W:�t��H0@ԃE�]uӭ5R껭c��������*^��t��Q*Za�WRH� u �y���f�Ga��׮+`�C�c���IGX�z;�:��P���>�J�=�fvro��o�0ڧ�M�h��
����k��fjf���.�n-����e�}�_b���J�up�#��&�/��n�̰Oٓ�fh�|�Rd�#�u�vT炕[��H�݅;-�L�]�&��h���c�;���3��	�CۊR�[�NE�ȭ�m�8�7�r�GR���U�{����u�P��4�o�ƃ[:^���yut0��<B䬳�)��tY�)E3W6gi��g��M�ڗtu��5t�K�����O%VE,a��4���:��9|����ŵ��H�T�$#��g��ͫ"�Z����:V>*.���Z�w@�d����ukC��J�k�]MW7;-��U=�':mM�a��E]֞�Ag��R̩�5�*�8h��fĀ���n���_U�v���B�;k2��1f��>�:����vKנ�g4��b������N;����`�S�n9�6ދ��	�pI_jɊ������M_��I�.
�xr������΍+��j'`m����k.�]�TKG������b�w+�r�Ή���:oVn\*�}�V�'e��`CR�FG%��T
�r�;�D��&����w6�3�NJ��V�.�h���B#SY�`�Uz{�f�ڵ�;����3����us^/Q<�'��+�Mz��ܽo%*_�!��t��Y���]_J�m0z�W݌�̗M�mD������|��+Q��i D{ҝ�n�ٴ�u�����t�[�%'���!eepYlj���Q�M�<M�	_^��n��t�cs��C	��a�z	Ӈ��U4�GD�h�05@*�z�{�4c�%�V:��R�[�Pұ�:i���hA:MQb ���8s/��J� �spR����Yt#��u��[�+Rju&�H��� I>�8�Q�eǴ�z����k!�64���)<#�?���󀊨��������������������8-��?�}z�DY��H�l�ğ�?�pQ��	E��D@�bܑR��
I$#�J��*�8؈��b�`��l��A�.\�9)ÁD'&��`�����S��};����Z˝k�
y�q9E��`�׌��ztT{R�m��q�Zl���7\��\�;Nc�O,����.��#�dT�}���wps��; �7��f�Gv��6�Y{y���gTW4�"�t����{k�����W}�=Α�8X�Ҭ�1�ص��#$�ڌ-�J9k"�<����uqE"�DR����1�$���^,`���=���XΕ:�js:]<\2��5Ԫ[vy���O8��g%�|��P��F�f�!��X��������{7f�K�;�e\��lx������{҂Ube�)r�Ǚ<	6���]Ϯ�4����OqM>�9�g�&n�ˁ7���dSR5c"QkZ���5gH7h��:�r�	�h�A�J��Z�Ս�k�Gy.��̫�zd��՗3o���S|=lZA˩��QF�r/K�N�n���*�� Ȩ�'D�%��5u�
��X�WX��Q=a��,��ph9
�Y6���U��ENTz�V�cX�E;�(�m�[�'*L�ݴh���o�B\���C���;�
me��wp�ր5�KtLV�Ć�$�K���hi;f�������+�l' s<9�moweI36NO��G���	[9��칙�͝���7c�C�,#nL}0�r�oB�n�V��E:��T��_����)GE�Sj8��"p��I6ˑ�JI��l%A�����B*�u�H�D@�ˌ�.4,"ʈ3��\q̈́K��!L�Pa��@!�0�
�%A�G M���%?Ŧ	��,Ȅ�(a8���5J6�3
- L22��<�~E�UT�+��bmm���;m�b+m���h)��z�N}�O���~߷��~߷��~?��h�e�|��4}���ГEkTP�Y����Ga�Tl�s�����~߷��~߷��}�����i���G�ߙ��:j1����1�9䢞�U����F����th�[V�(�#\|��TSV �5UDTE�7�ܔ�[.�W�����-[m��QS�J}cv��ۉ��cD[���EE�AGlUئ�cT�5&�E��V��Vى��Ol��F�u5�&d������!��N��[T�֊i?KEUt5ѻ�b���j#M&���4Q���آ�wu��>�����ti��Gn�w'\Z�`��۵�qqت�Ĝ[=q�-�.�����\�Q����wc�q���k�j*7c����k��^�7����qlt��y�j<��u���%Zh�u��-�k�Cf�t;Z��i��:6�fhfv��v�j�#�&�h,�A��.ؐ��C���b��ALo�F��O�1Gc���t:ڍ�� �h�͋�PqVچ5Gq�Y�#cN��X�K���Pѣ���`�nE� �dϿ
��hbo��u�W�"A�R�M�E�]����q�ױ�b�@܎�i{3M;���'q�V�(/Z�z���=j�G�H)7��!��� ���P��9%�`�T;�9L��{Ք�L9�� j��;�-�\�E�ϻ�'�ݣ�<e�T�3D_��݌��'�]���^D7~�gI2lɡr�v�M�>T̵uV��ϻ����==��6u��&��Q�b(���������*��L��	l����m�Y��cգ�V�k�y��U�	���p���mG�շU==���׺=�
5*��}�%>�G�Z寷�'�i�y5F�] Ԓj��~�Ou1�Ȼq*�
��W��כ�>h��xS���\�E����<\g���4h�7������׌#��ˉsIc���5yTR�F���+���s�f��}��T��K�Y���9�a���W9vUz�����yF�����D�ryOI4�5��C�Ň�lm�L���<&���V=RXc�n|Վ'�Ż����i���ht�O��I׆Uh�F�A`�kv24�N>6/�{���\�i4J��EdFk���n���q�"b��.s���Se�s��'��vL)��� >��;K��՗���_,uh�{;����Zܧ)Q���/p�ɔ*�W�4���M��t?z��6~(VsOoh1�f�����[���5-���I����dyW6>�AJ�����s{�"�[d0;1ѭ3]�86{-���`H<'z�_�1�V�q����z�>�\h����H��+�f�W(�W.�}Q6D��htdlS㷙�a�ng+4�\`�6/a��?]e��$e�:M�I=�<���B�/l�NL?|��nV���is�6Md�f�9����57L��_�E��UK�{Ѽ��������c��5�v�>����z�����ܷOa�4��8r�M��>���ߏٶ���^2�{]?�rkw^)go����V�zK��k��	�T�}��~���f�1#��#c(�_Q���8�]�y���A���2w�Sq�ʾ�ow;��XOu~�}᪆�)?��k�:ޮya��d6��x�T�����V��P���ׂAP`v��G`������δ�V���q̚mmo�]R��7�U�^ە�����ؚf�ǡH(˹���r�ĕgf*�]�Ͼ�\�IKW$
#�hv�ڌc����y*�j�}^�uxI���:�v�������&�7ǁ��W��4%3@y"�U\��o�ߡ��lP���'׈62�p{QJ�~ݺ�E�x��Xt�b�ꭚ� ^����u?y���c���;�ç���C���s�Q��L�xj�H�z1��o����\ZN�^�qt��s�}����8�����8��a�]�m}�*v%zO�q�]�s�k�i{{�'f�OW>���3�!yUtɵa�J���x��<�����ڨe�pj���n˩T��R0~��f3�d��k�p���e9��G�҂�zĞgx��ok)�O��W�����N�Ţz޹�{��Î���t@6��T{��4��N��D���4[߷n�r���U�i�cY^q��v�1��l�Wp��ˎ�z#�r��Tåxb��JX/�!}�ЬȊG �-�OƳ9Ӧ��[��A�/��s�R��չ�sm����$�XC��:�^Z�c<۶�����Gi�GZ���ۻ|�ﳆ~��������1�t�}BU�ׄǈl�Ӎa���}y_U���U��7)r������5y��L��|���Wu[I�˦tu�͟޽�ΰ����9�	�M��ؗ2Ī��֒��5ud�7�����0t@���n��mohs��&OA�4�r6���b�3�:���q�XM��}�G�y������z�P��h�oO|�|�L�y�K�롎�քK���@{�/�����6l��+g�W�履k������7�V��ѓgK�;}W[+�hJo(�<�.dޞ͇v}���:�{މ�YuS">�zJ��C�ͳlx��� �^#y����t3|/�F7��C�&���'n�ޛ��>ꩇ���|��I��=����#�$�͝�5��sf�$�q�OI������Sڶ~�I�*�LZ�ظr�9>�ur"��Q�ƵE���~y��g�B��~��h�>%^�m3uu���L�:u�v ��m+|���˽��v�LWrZ宜lo6Ub�q��/��7~�%�e��֕�m�e�Q8x�v�:�PF���i�������g��k��0<�>+
��hNY�:阞�Mw2o�Uc!y��Y-Yd�)Es��*1�#�U�{s7��c7	$�m��8����W���9OV��:�6d���%-~��u�^�7���3~n�g�ۇ�2��<�z�+�B��t��~������������5:��진L�B�r^��u�>�է�Hv�=yػNt�6ww(��pD��g`�6��$H�~�������P��wl~���Y���W��3��мq������s�/W���l�v�v�>Y~ܷW�r%���)'I9*+���� 	�&��mM�u��:M�:�[p�k\{ؽ����<��O�|}�jwѵ:�	[��7ǹ����ĕ��kk_��哙y�����[�(�~$\��b�p�V�f�&���.ZN>8����c�.�b��3����Zן^��$jW_��L��E�P�:G�7��է7��6o'��h��&E����z�4���#ݳ�1N���.�X�ټk��{����Ú�Y�ٽ�������l!«�b"��'ό�>���i��(+{UZ��Tzfz�Z��6x�u1W��V�����#�sJ���>���Nu�}�<�e��,�"Z�m��)`FhF[�Zu2�4����4
�]A��Y{�=�۹�W5dߞ�_z2@�;����0�cd0�z띮;������I�g��W�B��u&WI۴�Ϸ�õ�o=���=.��Љwj���^���N~%{>)�I��9C��'\�?��|؞�O@��1>᭄o@q�כ.EVѧ�x�%�{b۬y��r�k��{x��+�Sj���өb�z�]6�yo_E�>Yw*�g��>n)�����}�!5lǵp�3cÀ @0�x��ɹ9������U���j�u����{��I����ʓi�i�~�z�����)�a��~�s!}�j������M�](�>�=��g�~����6Z�̩tM�y�{۹��֏��z;wْ���1�+n�#+������;���D��e�t��2Ǚ4�~�X��;��h͓C&#7��$Y���5f��x:ʝ:�H��Q�P��n��{Y7�3��r=��u��K]C�DZ�Ci�7D>ü������y�O.����~���^�ش���l��q�/Bқ/�9��od�e�L���}�74#7���%8�{]^U�̤���7$�G<|�}�ݕ�������ye*<ht�����|�����z�JF�������0v����G��x�mU��0�<��.�X���c떛���ݷ������I�w��c�ƨ>^Ϛ�{)��Pp�X�t��8��o����FT:�~�I�����1�+��T{2��Y���ĵٽ=�U�ԕ+���y	O�9��^w��?g����W���3�����dݳ����v���Z���<n���3�H��?=ޞ�7�g�Tv�bū�ׯ����}Ȉ6�¿f�FƇ��+��1A���/v����xC=�,S��Ή��<j ߌ����7p8o@�2�.�51�k*y���f��*����W��?<O��7�մ�[���unʔ�FXۧ�*��wO�t�Kdo�O�ױ�j�/}�8��o v��wIh���n}�ڴ{=�_]G�6���X�w;_\��9å�|v�R�������c�y��2)�����EK�w��Ū�o+��u�ė��n���:�T�v�ɔ�Σ@Y�$�2h�0�9,��������B�x��D�me��m[@	��X��&N;}}��,��$��uw�O?�Z<�s%c�$bud��=Gr�{b�9{����ؔ%k�g�3�_rok9I�Y��ާ����gtޓw�v�hr;k��)����,tA�w�ܛ�)�0�wOy\��ˁ�M�i���Y���0����6�ί{Y�������^��_��f$�O+����o���4�۹���8՝��3�򲻄rC�ޯ���(�w:2{�\v���r��4p�1ч*��4�EY�|�~K�y��L���ssۀ��Y���������$׹��'��g�!�"i�D�h׺�$�d�?��9�~*��S߆R{�{�'��J���%A&��Í�ľѼ�ok�qt�2�E��ewϘ�μFxﯝ����id{�=���ȯb���D�ȱϴK�vW���o��<.o�%���������i40�H9���I��o&��dso�U��:lѵPR��-��T��bS���*k�])c�t��.��bhN6R��j�˧�6�氱�hUڵ5Ш�ܺb�U���!���5=av�Z�����]���ی�3r���L$�mK76��3��tc}��y�z!>��QZ5t����I��2o���T���7�w��{��Dq�A�x����&N��ݦe֯�'��.�9��[��q/E8��7�Q��|_�7���\~[SӾ��jH͐��Qq$��6^b�����k`��x3�wz���@&�v]oF5�<ƿX�NxR�!���$����Tz���\�<9�`!��� �"���p��h����ܝ�<	��$k��=-|���6�?�����_0���{�^S�M[&�լ����l�E'Uw��+�{]� s��ا���:���'oE	x`�{��k����T�ޒ��Ҟ{����)�^ᰫ����D��Li�Ѡc�i��"nM\���;�A��hگz;�O�5b�컼�O����瑋U3Ҋ4�]�j��ߥxm?{�z�<��-�ד��X�5�9@����v�����aQ5�^�;��*&���X�� �&�D�>u���X=�}j�t�����r�ý�H����8�ܛ��#���:�<��Y��g. �]"��lS�ׇeڨ֊eld�a�q2�n3®枕U��Z����}��L�6��9S@�� Mi��^�>�FoU�O�W��>m����\��W��~�k�NI G�#·�[�[����H�b/ժ��>�G�O}���w�l���s�b�v��ގ�fI���w5�t䝽�_�Y�x��05Ӡ�i�t�F _����&{����vT�sy�s�l�_�����M����<��}�{=&W�+��Ei�YQ7���5��z:~��BRxL�&t��Nz�7�[�8�+���� �E�\��(F
���=����|��?��7~ϊ��vU8����*�Y�{���7g�H��M����;�q���>�g<��y����J>�gp���L�|����������KU�>�k5��5�Mf��]��g9e�C:�׃���m@�}�Y ���ح��a�`�|�<��]�&�}�75�n��zs�y��F�����V�dUyx�Y��uD���J����w�5�vBd �f��"i�絔�+QV7fЧ�k7EyirP��°�shG�9���n��yV�N���Ҫdu�1�h.�q�m;�,:N������Ng`�YJE�sfv�m��ƚ�9^��fl�� 5����tk��JR5�[ݯ*[�*x�.��S�����-�c��M�wST��y23�L�
��Sn/��Z�Y���Ce*mF�>���Ip�P��,;�ڴ��wԻu$��^!�Pԧ��4�i̙g+���X�SU�9�q�>Ani�X����r�OCg���,��@��;��������m��0����ҭf0�VT����wԢ��B]}x'$[����uB�L��j@nĳՑ���)š]37�s�<�?[W]�Y|\�S}��ԙ�ɦe�Δ�r��ls�݆S�ZG���J=@�̬]`oa�����zS��T��o�o!(�fWX�g"n��ʢ���Y���ռ���}���St�-�
�t<\;]�:���psx�CfS��.�$��% �DR!W�;b��j4�j.7����C܂g3aM�z!m���]f�}E�Η2v�N�%�Jh�e��{+��4�8�5�����2�*�ƃ�1�3Q
��m���Ox�x�:�4�-u�;5t�cmf�t�a��w:���U���o�ႅw�Փqӏ��{�z�l�,srL��deݾ�c�`��*�i`��S*m	ם��<և��V���?}Z4-�dt��(�[R��6o"�ͩQ���"4��o��^�U�|��t�1g)��)���#vjs��+4����:ó#�(՚3x���tU�ZNq_\�A�j'�����Ai�cu�Eʤ��F5Б�K���ڛ�[u��9���������r1خ������[���om��	xӎ^�<��}�� ->��������Ğ��\̱Ҵ�{�m�<zU�M��l��k����-�ة�ɟ�>��O��Uj֛�Z~;��U��[�˙�Z5�oe>mK�qN	1��W]��m�cO�Qдcl�5�*8�`e3,��$/����N�t�d�:,C�q�+*�M�N5g/$�57b�ü�ps[��6��H�0f�	X�=2ٮ"�L�K�1��JmL�Z6®�Y�����㷸2N�Dk��2����u-��u�Ž���p�=�!z2�Ac��k0};x��3�-�2Kk)$�J�*�:��`	��"�@�>��T����b&ZgU`�x��v!��K��c϶ʣkz��AKv�y��U�rٖy�լ�C��hY
\��%c�{�o��M�����Q/��GKS[���X�
���I���\s��`��Ւ�p�yd]t�]s������"��Z������c���h����?����]`۷t�[]۱���I��፲t��������A��kF'F�x��V�Wv���s�X�Q5v;����ŉ�>>ߧ����o����o��������w���>v8�O�=����ƨ�[�yQ�M�ˡ�շ��U^o,cvN��Wv��'<�������o����o����2��IDlcG�&a-75��V1�����t5_V�Y�?9<���Ǫ�i����o+�_�j�:.,Dl�w�ϕEZ4ӧA�y�y%TK�`��GC�������ӭ:�qUD��QA��J��ht]�btFѭFѶ�j�&�b ���vn�׫q�bh�wWU:��V1����:�=�Ӣ�F�k Z6�9�w;m����:`6ζ��i-�ll�Z�h�(�F5���(��k&�DGܚ:-���-m���^MW�M4�ѫcA���:��WٍWZ<��"��>]'F����LSZ����j�k�������v9�L�F�����Q��mlQ���Ejт�iւ6[��ڵ��l�z>����}*@L]y�*�R;]a>�,҆�DΗd�r����Dt�/�8b����H�̇�JV+U:ݡX��b���gkz(�� �a5 E?�^�걽A�skCHނ_��8�'���i�}����񹴎/�����������W/'éd>0���^=���i��L�@vH�%rЌ�p�y7~P���?E�p�'2��7rx5#�ต;x>0�<�d��>���&=��1�b���v�9��G}�"�`��A�2�L�^NN����hσ��'�M�� S�`qm���������J����Jm�������v3�H;H�_N�_�M�����ތ�B��~SJ�v����Xx"��!�v�#���q�IJ�⺚;U�F�Cن5��pok�(ıR�&�}�����/�B�$���|��\��X��,�y��k�0��BG	�'��"K��b%9�j�
c^Ԟ��ٯѹ<��\:���'�e���mW���7����q��a����څ��}��0oQ��$ˉd�g��Q�b�oj�˩\1�Oi���s��Nw����M�B=�m	�86���R{T�M�M����U��+��#����t�M4kڬN�̄=yOP�J"���G�>zQ��-��
����)���U�v"�G��c����h��̩ݏ.��𘡍��^u�A�V���vC.uq�%J�H�����loN��Ϫ[��Fn;�"m'��.�WY
�Ɉs�;�9�[�r��=��s��2ݶfAX�eNos���-%v��b�u��#��</b=y�Iܹ1ɪA�1bſ�5��+7�c���HA�g�����yċ��Y��X�-�G��Z F.���H-In�L�8'��޼k����8V|�����%�`{ϩJ�Oަ�XTF1��Ny�v�,�?#�
�Zȣw�h�gC͌��+P��2Xu1�e�|�}[@�ym��H���}��v�Ԩ�?c�f�����<���ru]��K��I�,��
Z3��d� Z�1�g�娽�p��)�눬̳���H��3��-�v���i���n`c%Y���󝆄���C���	�����<�Vo4N�jsQ��\<���:|XH�Q� ;���	9���so~o��&�$�c�(k���cAy��{�s��-A�]0��p1�ʹKO�6
I�w��� Ȱ�����\���kY鋹M���v-ӝ�{K�3.Ckq��ptQ�g͊`�gO#��`X�}�5���Ó:y�S�}�)M�:kP���:�TV5%'����M=h@��n�N��iQ���שi���i1�t�=�P���p&��F�a�7ڤw�{��˻:�3�%�U�w=C�/}x���k�P��~�FgY�2�n۲�"�yJ�y'WW�3��B����:϶`,G;Y�Gru��ޠc|�龏�7SX�{�X���2�Ӌo%��
�>�Tkp��\K1ΧJtٴ�ܕsk���RI� �-m��l������6���n�Π
�!�2	� D��;��н���e�׺��	J��f%ӑ5��|Wư�-��P���9:.�<t�k��M�p%9)H� )�⟇]���ⷻa��?n]<c=�m���Jq�y���i�9AĎ���2�},�4�v��T��55���^����I���r�pi�EP7���"r��v� �<05��������,��N�|X�uA<��]��8>w.δ=�P[�Ҁ�6ɼYq��o<����!���*/�����h�y���.��8�R��k;mgL(4�UZ��j���x�,Qن��p�|p'�|ɻ�L��{"㮪5og�a-�ԟE'7�7^o�̜qv8�,(Z��3* �8�+;��O�@�bU��J�ӓN��U^]���#�5�����Q�hL`2E�i�q���r��� �Q�'�m	��@�����L����޵R.��G�J��q�Oelx�Â�T��~N�r�q�Ol.͚ܹ�ްG��4�/��˦��pȗx���4?�i�6�4O�/�f�vە�7&�ص�E���j]�P�2`��Ş�*e>��sW���?���ycS�P��-��8�\�Cf��>��y�V���K�BX��d9S�;32��kAPP��]��36�����AmJd�Oa��G�C���0�ܗa^��;8�@P��y�k�/,$L?f��br�S�8 7�DHz��fK������_02v#G`�3X��&5�������2d�3���\�;�86�DN+��;���Q醟l��m��Ɔ�f�G���<�}k���o��{�6\�'�N��=�Q��j-=��0��	m�dΕ�CB&��n2�5��u�,���݈yt��;���C�����\H����&���T�0;���gaU�B�����=���N��7F�e�a�����.���ג���*��OBԹ�w����!�m�P
N�3R栦�������"���|i�sR����� H�"��C��5��Z�O0Є�Xy��N�d�x���񻜐e+Я�li<��a8�jF,���R��hG�0� �Sy��;(t�dr�u�'�7m���{\ǐޙ�s��zR���5�O����JǭBB��&Äy��7��oh���]��Ϳ���������w���%�.���
cX��\7�r���^�Ǳ(;`�@�a��כ�ݤ{�;1d#�pX����~sv�������֢��X*��@i�"�B��|6uNU�^��g�<��?0��"5��zKx�a9^~��е�f���|��j����Y�-���5C�[o'�cw�X�\Pͤ�Ȉ�2�n.dŝC��r��9�pUn�bC�jo���2��ʓ���y��%�Ӯ��=ʟ@���!v)�!V$2���i�.���B�Y0%��{�?��?�����m�C�L&�����yÌ�����ָSتv�[+�kW��q�/*m&W�&�r�s/��WAi7R͵�E��m�AZ4��*�/q	�N�Ƚ3m��_B̉{�|Q���l�;�{xŶ/2������zc�NԳ,3���xy�����U�K�KqA�=�L��j�NR����mVd��c�^���^}�D[�Xgc��jA�D�/R�uUO^_�O����4��!�q��Nd���6B��8
�:�M׼Ұ=��� ޒza��-���Ǧ�a�������/����hg@�ZF�	���|��ǳ��:��n���ӣ�K�����L��x�\By;��f���e*��R�3�aqf����X�/d�?O=�ƕ�S6�;*��_2�I��%�+uge�{�_��'w.�z-������!+I�{�CӴji/dwP�yjͬ�뼯%�9��C��F6/r��,SI�	�M#ܮ�-U��B�%�����-/CΞ���ꌅ�8�����=�����.��/r�d^�Ji�#)����|j�Er��E�Π4�qa:�^e?���Ӏy�z��-��L�n�5c��.1n�;}g�d؆�;C`�Hl�{Y�öq�w�Q�l71�K���l�\w�(}���Դ���|�^��ђM�VB�W�sc��Qg(]	���Vw��F+�7���U��8����� &L����}�F�C�ӎ͟L&��8M��~w��? b ���H�4������3Ӓ�b����k̢��W!�op��/Gf���S��f
o��$oQ����y1K�|*�qW2kk�)�a���lc�c�w$�1X�&^M�Q4pvu����0��Zu��a��	��\�����u�ӵCd���]�l��N����m�TBm�zB�VE7, `��j��b�;ŉڽ��TE�����Q�
o�No�{�������9HM��f ����'Hν�1�!n�tyio:��)��S����c"�Yf���Cۮ)�z��Ґ
~lF<ʏ%S &�����pr��z9=k��n��S�ڇ����Ի'dz�гa̖LoӬ�g}�?W>�|r��u����e����O)�9��=ݨ{�K:"�D9l/B\���"7s�'",7�@��U^�߼?q�e�U�G_~nr^��А���<D&�C��L["ak�*����{M��rh�q�`\@:ҨVuUFJ�ܹ;�G��Í����ͷ�ƧH����2ƌ|@M}����/X͟�<�mg�ϔ������%P��ڮB��1���t���.u��*F�$r�o>T���ރvK�޳�K�c�/v���GZ
W�5zןZN�����ICTX��r�� �E3ie]��rpɮ�>�2,6�9�z����n��jL�ֹ�l�4��bQ��i�����s&`&@ ��2���_����ɐ�GR�]��3���jH�4��Zz�m࿫\RL`�|ջ }�r�~�>��Q��G����uZ�Cݯl�c�?�����!�gX�fͲ��l��sӸ,��|�=��M����2ȶ��s���7P���7VTV5�B~>p1�OAd	b�N �>��|jʋ�5q�ͽ�.�,Qz��]���!����Fs�,��d�2a/.�c��9E'V�W�+
�����8�#�����T��vm��/��e@ZZG?�S��lVA:"�8鑮��9w��"�8�g?R�N҄�ޖ8g.7�n(�'�bȀ:ދ��YhVk!���A�i��`�to6zx���ĻM�	�~=0��C�.!�W�����X�j��}Ɯ�')9���fp�<5Et	d�'�8����E�^q�0��Nk�QL��^4��:�f�����?<�V_��@ׁ�Q\9���(�}����D�Y۰�{���mP�c&����\���K�N�m),i�a!<;��d><�|mzͶ4�lfK�Z޼��#�X��b^9�	�B͇2q��E��]<�eN�MX��@?Ϳv�����!^�P���vX}�w�2�X��.��@�U�7!Np����h������~�+�W0FnC�v�(-e����㼣�{K�״O�:c�;��t��'��ǝ�Vrv�M�{�T�&v����2csrZY���k�Fa���l@? `>62̙2�3�y{[}�� �BG>��H�>R�\����%�2��922u����Q���h�\�fv�����*	tlr���Ŧ\,�����d�t��yHpK.������a*Zۑ�<�m�Ї���C^$�[�@���03�8�%�7�8O@�]`����r��Ga�7_Wh���㳸��<�{�O9Q�V��v��-�{�[9y�חt����C�|a��>��ө;y氏m ��K�i�G�"��z!�p_����<��_m��P&��D���ۡq��Vwha��Pk�W�����C�i�:���i�	-ق瀖HA#͠\e:j�<G��� |}�ÜQt��.�W�7@�"#X@!�L]���Ʈ���Ơ�H\�veAfP�n�x�F�I�fS=xث������<i��1P��Y�Z�pL�p��k�%�j�����M��R$A�k����2�v_m�C��	�BW?����VF�U�h�O��p���,�#!7��E�j̣��� �W�۽{�{���(�J~)�	�c�%/X�zs^��O�Z��Fg�pW"xr5���#��X]����z"fW1��i�6Z�=�h��[oAX�G/��ʖ��Dԧo�K����'��!b����< �ua�}���C7,�N2���fE�Cj�M�rY}ɭ�3�u)�x�e, WI�e��w&&|��~��s�\�"�y�����޿O��������y(��w�Ĳ.�s�1����:���w$��ZX�̜�N���f.x�(���^�,�=m,3�	r��ҝ��(�a�aHs�1���ۨNY�6���{���x��M�����;Ʒ���d��ne���w9��q�S��*v��N'������L?7xo�5s]�����iZ,)�N�u�^d���By���%=����oq}���0��Q��G�����~
~jz�=��
�G��A����q�<���5�� �vp��]B8s�Ə���Մu�X���|�{)�q�o�kq�yv��0i��=��(搮�;˿Z�?�Ga?�H�_h�����町����,({vc=nTM{o�� =�O���4��f%�<3�@fp8#���P��T�����t�cDWK��l��@N^��]����]���LP^j�� cb{�8!�[þA�N'+�
^�3�7����JL]y�Ъו�P~����7���Y�	�-��ې��C�6u��of��y��ĳ��-$d�C�$�%�߽gz���4�5�%�%r�Q�Ы�޺zjf�ث��-/��ſ~c�����v��n�;]�ۋ2�᭽ɻޝa`�J-]:�6!i�Y:��Wo2e�uu���9ї�t�:�3K���\��ŅViEM��~X+{���D��y[��ؚ��2wF<\��א��x3 ��ɀ�&L�{Ñ۞7�v�<�����e�y����
qa�`�m�*�¼0Ѫk^�7o�53?�=v6[D;B���j�+��y�6a4{�AVlϖI��$�!e���n'���l�5���;�]��vn�=�����lO7X�(2jX�������<�_�U��A�Ġ�|��j���>+����K6�x�c��R2���j|��Ƚ���B2�����Tc����^�5��;0���k��J�5��Ț��l
��k�V6��$�����H�44��k����cY1	�+s��i����=x���Ôy�����FY���S��f
}}%�N�I��Rr�y�6�E�d
�\�Ef��Q_�pV�z#���q��@��j/�C�Y��.�M³��/Qku緫c�G��e�y�.sX�Fm������� G����G�V6�Q���l=�7�棱eD�a^�1lQ�猡j��j���*��ćA�<��+�t.�h����(��}�Y�__^��(I�LhA5mv7���FM�ʏb����"r�9���0�� f�(�~KJ��U����u�"���Z'��C�WQ�s�͡�	��*e�;%'2���ytv��l�
������p��{afXk��iYrL�e�]`uTm3N�cF��Cr�I��7���q\�\�q�i�ދ�]��{���U����܈�t�ggn�ԋ4�}L��x�.���S���)4F��c��ژJ�.*fR��-\1vB��
��v#[w|b�dwCw�-���F�Mڥ�����PQ��X�>�@k&���}��[���c���S�m�"̦ݯ�d�ב��5��|�W���R�tp�tF�|3��ȬW�NlU��9�d�X}�:e��B���v�IS.��6l9ԍ�&qWpL�Մ�O�	\6m�٢�o��`��̕�Ef��*�^�
�y]�Dn8�z����dUT����vV�:\���x���q��Y��|XqZͣ�������N��9��B�\�J+��9�i�A���ĸ��a=��ϸuj�|RW-��FVEftK��)Sc&^q��ʓ^]������z��w8�bs���V��B�����7��D����Jm��������E���"C,<��m�:��1Z0��{���O_J��+�wіt�w�rK�R���[��1�u�[����jB�]v�8��:��ḷ%�U����'r��V�0�<ud��w,`��wZ�+�.g��Ic����e�2Ç6�����t�X����Ȧ�L�]���5���*�3x�Z�W+��䊛z?S0f��z����).����S�Y���v"#��ܭ"���RY�L�F�$�����{�롼5[�&GnYg�����ܱE���k���O���i�aV��b��K8yJwζ������ِ)H��Y�i�o^���*��^��)Z��6������4��F=�d��L����醸�ЇVU,f�X��5��J����C3�-��wŒ�n�!Y��J0SW�F��y���$o'vya�m��ry�0h�[[HdR�'rs{h��v��nM�*]C��nD�	�sD*�*�m)��_MB�g8ni<�mh3u�[�o@�fW6���Z�[�u����8��PG�TN��O2XG`��sN���q]N�a;�[|5�ʶ��v��ҕh`�;NpU�R)VN��]%��[���7S����\�77}u1�z*:Sxd���!J��;xJl\���5/Z�ri�֘��+�㭸utUy([!�\��'�T�C.۹�{n�wn6��/D{�&��w_�O��g6VJ���%[�&�t^^��b��C2⛭f����
��J�wgE�d=����<�L8m
m��W���4,�������Z֛��o9�J=��iT�]N���F�/
݅�sN��2��a�g���ܤ[M��ձwvsR����5e5MӍ�e����?~�ЫQ�d0K8+~ps��]�[�!�~��.51.��5�����}>�o�����}�߷���ϕ�b ���CAƫ:	��\N������c]uA�~?�����>�o���������o��h�#^N�j���3٭4�~�7bڨ4�Kq�nԄWY)i�4�5UDE0h�4��Q%�:�I0�V�tDm�b`�A�"��'BQGI� ��5��zӶ:s!z��u�A^Z*�����0MI5)I���(*�j�h�Ӷ�K��g��LJU->'����(��gm�=�F��"|��Z���4�QQE4���i�@j��4�W��:�'F�3���b��/�h8�Ο#�QMWd�4ꝰSZhO}��4V��h���7[E."���Έ��MW�XtDu����l톚q��Bcy�����G^_�~��}��w��hX-��q]i?Pwba�ݹgS��uYݕTr�E�[�М��Q���LpY7��0���@ �o,�.=��5Ǡ���Qd3,DR�5;�uԝv�3���/<�UO��0`�2f�?]\yǫ�J��fU�΅����J(��&�;��teW)hG�υ�j��K�1�e�c�O�nMsO���l��r�vR^��^�ɭ�ݵ����g^7�D#��=!�E�� l23L+�h�3a/<�=��&c�K�m�G#g�Jsܨ$8������c�h%:�s�`c%C6���v��8ԗif�mJ��,c�ᕼ��1�=)�Y���<�>wʱ?p4��po��?~����O>����g{�߹X��.�"WT������W�3m�I�sͼ"���	A񅇸�E܋�Y�Y���v���ޫ����ݙ�|szq��H88�77�Hj��6m�dgO<���4�˴0)�h<���g����l�#��¢nF�m��X���_��	�,�-�}եW�b�G��vנ���i��0�|Wyz�{�f�\J"'\eL�Y;I��MY0��tB��r�N��Q��Y5E�4��4Z��n9ƮZ�.��e�k���Y�zf�C�#�	���N��Ǔ��D����:�ԃ4z(���[���5j����GN0�Iɓ�fu�E�4äL9�V�7�ޗfU�kr61�.;߯b����v�G,�ЎPٶ劼�۶8�����a\�W��!���꧘�Q˄,}� N���#p�C�tCX4	���6N*�~��e�.
�e&�t��͍������ClE�X6�c'Ή�� f���3 ɓ&ff �ffu�ޮ��ƍ�0��p[���k/i�o�Ӆ��-��r ��"��[R�#T�ܾ]�~*r{oP�+�U;M���yE2�HK��-�'��BZV�nv-�I���n����ݑ���Υ乃�$ٔ�M�\��j��Ib��0�	L"a��C�����U��)�X�������}n/�8Ȣ|�N8�Uk���ҭa)�ZM��m�Sju�R���t�á.3��^b��� Lj`kd��Bչ��8���A/l�sʞ'�/rޖ�[[Y���G7�Dq��A-�{b�����E4���Pl
�e���L5��J�A9m�VR����T��Q���������4fP�C�ܬߖ�,z~�"O�0���#ɾ�8&���ڛ��s��[��vZv(���z$�z�˱�&!��ǜS9|����\F���F�u1�`3����҉{`��6�ͧa�i淤"�J>F}�,���GD����-���̽��3Y����i��v�Fd��4�ض�7k�mB2��' �z	d�)^i��S����@�k�%)ۙ�:8h���D�%/��BUfKL%;�!�}v����<����g�݃��~���nvp���.�R�s+�>女���w�p�ʘ��S0���8w3msݕ�,�R��r�ΚgKV)�k7�h,,c����ofr4nPJ�vBx]`? f�� ��&@���}�vww������/|��W�����Xʩlj\�.s��"�(Q�l�T��a��_F���"�#8�E�T?k�=�	���i��+c+کnj��M���%���_�f�J��\Unv��C�̂j�;q��!ʅ�/ȰE���{��\r�})��P*Ԛ�o�|�y����;����j���}�S��B�ѓx����yN6;�aM�:A�Zy㔩�����̾U�5����]��Y5����N��K#g��&<Q��G�c֡*���Xane]"Ϛ\��t�j�=z-3k�0<�K��7�D�}Eހ��.�X�ީE�3��iۨ�S�I2��0֋���Z�6:w�#��Y�r��`&�ƅ2����]i�?7x�,��c�����T�7;6M���מ�a�!	?[b�]�y��}�]��='=��[ ��gT�}8F�=���ֲ�%8�YOR������Ӈ�p��:[��:��xlY��ʫx���Y��{vZ�m��V�j��{J	{��J9�]K6�3��23�� ��v������9�:3�"�����r�l��R�*ڰB�wszo��cSƣ�t������.f�yX%\MK�~�7jr������CC\��_�U�j�tj��l,���-gHh eY�q����ڏc�KfV�E����W[{�m�#i$|>{���|��_G����s������m�ĳ-3i���u�&�eO�9O����'jY�^��ȷ�;Y
��Qڍ۫�WĹ5Vˡ2�����K�>���}{(�[���ų�;l���ų�C�.�l\��m�;]��T��k`��)����{�����ٳ�!�z	C�@"A=P�|ڱ�k���=�S�^z7�H�򸊇�^�h���C\�����d!�+��P�nu+�x��&�*��A�y�3���jn;u�{�����sAK�~T)i�5B������<�g������ߍX�p_��Pbǒ�䓡�p�obfժPcK'H䅀^@�E����le��B��]�Nѫ�#"zVS`Ն�Н5�5����/>^I	M�8����M'�ь����[�z�^����F�/�l�G]�:��to�)aj ݰ8nJ�nwA8�Q,��Ji��F�[���W0{hNj	̋��<�]�Wڥ�
�pƄW�Ivm�7��
�Z\51G.񮋣)��T�cIMmusIM�����Edu�w<,d����s�0�	$C�=�ZQ��J���ʷ@�Rr�h*^���s6�)��ǲ�i�{Y펬֒#2��MRgC`�٣)���:g��X�fz�`���ImO������:a�y�!�n�W]Hs����y)�P�!���G_qV(��ɒ������۶H�sL��o�F8��W�P�]s�,��)�6�[�}�mǯ^�TQ�Ws���'4i�:�M����U<�ݵa�**��C�)�ݤ�5�/A�<���q�y#��M�0Cl��5'��K�<wX��N=B�i9�R�l:���M � ./#�vđ�Am�����u�@(��O}��_V�.�û���*���J/�|׾]ˀ�bC��H��
!�5��.��4�� ��e录��Z�
�Ȕ�BzE7P�궻ޒ���#&�lR��T���ͳ��p�*S1s���7'637;��2���;'��%�_$^��9�è1�e�|�}[rk�c��=!��CjW�7a�Z��Z�r�'k�`�1g�幐��^��>H��n�����X�i�qh��e�K��YY�Y�{as.r1�R{�Ƨ+Ҍ���x~����q'��Ń;	�Ř��Z�=E���q����#��\��=�ߕ~�-?V����\�dL$���z�-˛8w3(M�����'t�չ2%d�Ql�j&a�������C`���$z
��zD����q0i2�/J[�v�U��x��N,�֐�
:��d����=fͲ��l��sӟ���l��)��H�0.�v��;�aQ��O'n���+��S�,����r�t�}���^�o�u��46��&�F�A��i6}�\��7���}gc�����Y��H��$�:��td��u���R�u*���8ۭ��ph����ͩ&2������&f &L��30�7��ݶ�d�ZmݳX\M�J򢱫����렝[�n'g�1��λ3r8VD��,ݬ[z�]Lw��`3?�3#h`��S]�#:ū&=�o"�!s�E'V��<��`��k�S\M������*o
dNNǞ�E��aOe@\Z@��
�~�a� ���NlBd��M���q�u�u��;94�/�{�Y�TS�����MN7�A�i0�qB�U��Cfʩ3O3Z���+�m��[yѦ���Օ�p'����(�y�q���:^��[�	�G�D�#D9	�K5�6�Z��h�ݛ��7��D`.�@��&]��
yC��"���[���v�����C���t�8!q�د=�{����(�7ѡ�=N����4hQ�)�х���r��PX�Ɇ���5����gQxss�^�:�^b�17�/:꧍7�\Sc��*�
�O1��k�0;��Cʕ�_"g77n��S�#~e�y
����|�>�Ɯ���j��N8�zV�q[+;�/u�����2��5yWދӟ�����w0B���%�a¾^�rz�#ņ���Y�2]���ve���Z����c%�^������B�!�ec������Vf�j��w���O;V�oآ�{�c��v���+�����^�yNR���z�"���
ZP������\g.�|Ƌ�׋CT����5���c�&�m�����_T{?P�W
&s�PN�篯��K�����C>e�X�P�秧�T��#�@���"Lp��Ƈ�&��W}�3�dw44.�;{F�V&m/K�:Ra\bKׇu�Z��v\�a�l��������ý����)�P�����~ͧa��p�u@$:Nd�L4�l��m�ilԝ�S��#����2�&}�
q1�%=���{l�ƫtC�-��5�Ȭ�W�g֪"F�]���w
��9I�Ә��\���yE3�r��$���̛/sQ�F�2�[��!s��A��Y�cӯ>.���Of�gjK��s���8�u{n��Pג��Ä9�!����=��ɘ:�`�ϕA��3�O3����!1��P���+���=;�^�o S�; ^�Ӊ/�&<��4dmi9<�������Z�PD�V^%9��0MAIR*�\U�9���r�X��B���w����Pz���|@L9�}���g>�~r�<SH�0���qOsu)��g�sC�W7.�n�޾�|�%��DA`����7M��xi;͘���=~�t����L1���۔KV�1��[}�0ϐ��2+����k�<�����
U�� ����3�L.�:�.�!�[X�Ơ_����)#.[��9]k�#�ss�^6[=�[�cT��n�%�{����/�&zT9�Y��C�2�F���{��aS�&�7K ���~��� g�r�g9UG���w��������r�}f`�٥��
��A��`&�ƅ�N�Y�+�|OI�ģ*��N}{4��,ف���i���EĻ�p�a��̅������>~#��납��~a��=�I�����=�9IK�}R3T���R�|�?�6�v��"�9o����N[�G��ʵ߯}��P��A��	t,~*	{��R�es۞��:C~���/����!�SWe��8wS�(ve�[�@7o��&ҙ��m��S�נQ��T�,Qa���f�%������5V���(:Fk�<���%ؾ�@v̽�Lu��I~,�oA1^:
b��C�S5
U���of]��;j���D�� �\LJ��{�J�z��f�0�����Š�5'Dɦ�n7Z��s�aC/s����z"e��dK< ���2HY��̵=�f��nu�'1^N���&U�X{0�ˑ�x�0���m=y����,�b9��N�de9�MO����6�T�5_����s�{c�����VE�,�d�#6q=z��]"��`qmâ�_k������l���݁냜�]�֠'�֎�U��U��Ѯ:N��Z�lwF>͖pCE�8�2c�	���i�3��G�.K}2��e�6}���r&7&����'2f�"� ���8b$Jޓ^�W����,���vQC0٢�hV���	�|�%��3L�0 kImߏ�י�Rd�Y
#9��j�7���"Sox�ɫ�M'�]:E{�b�)?,�#r*���1���O"r˓�x"��!%�H���l7%W5tB	�+�K"�R�ebQ��b#q�a٬rP`�Zv�T3�{w�#�d�D�eza0R/��&�O={�%:N]�9#T�b������s5�9^���\�Ϸ�22&���b�}	ָ�_BG��y�N�I��6��]`�;�Y�����0]/���"�a�Ú���#ϲ-�?��M�1��@��j/��詸C��ҵ��W��w��ތm���]yG-	�z���]4�@=�C�8�`|�[!����K
��Sf����ś����3Lla5~����E�7�7��=x��zO��ûP��v��롕�,u�o�R�9�w�).�;k��\��n��mw�)?5�2m�T{L���we���,�+��+����h`�2�L �E���z��k���еnd��c���ܺ}[rk�ʰ��l���)k��Q���vR0c�Ag�"����axfO�/M�Πpl�(�L�$�(��6Ks�vf,�4}�W3G��u;�����L-g����6�̈�;��F�
�[�j�ނk.��r_'2��qYjR�x��1�Ք42`WJ�}���n�e�:�ڝ}#����|�yV�Ó�������2f�&L��ڊ���>S���+��׉��k���A�L�����``PY��9Ɂ�������,iG3㯻;��C�ֻQR�ZA1��|tE��y����pC3�ylmzOܬN�ᳳiX�˻�l8��[]Vb��zCL���D���v��D�6��Zz�<����W�1�N�w	�N{�#J��_�~B�5s�V3kZ{a �JZĬ��F0�kȣ�n佔v�Ӛ|bk{3.�ܺ�ih�+���Y���z��u��0�~k � ����)�����)�h���=��/���,�~k��~W|�q�-���;-�d��0����-{��%[�ô�u�w�F��wR
��Y�.���Ʈ��sWޝh�[�)S����Y�M����̥א�F^?*�l�ݲ[�30���Z�%8���a vE�*��<��N��x�4,�A�eyK����_Bz]}k�d�=.��I����h_|�@�E��|����B1�}��o;��nڑ��`^��7e��;��_L��c��"賎n[�#k�f������x"�/�[�k�~cC}K)$�vgs�`̔�y��u"a�SNN3kh]�-������*�-������4��[�pm�sy\}��/^E`fe���Ab�o��4���e3at��ٶ���'����0"Ň�I��7X]+*pW[����ݸ���[2���	�u0'j��=7�K�qVA�v��R�F7������20��r�@\�6=5y6�}��(�r<���[�dn�U��ҍ�ͼ`9���#+������#��iQT�cԚ�*k<껐��ɡ��{+Q���S�e.�O55����bQ`7$W�vn��C9�\�Ox�+tlmQ{�{c��%aõ7rm2���ǆ��.�����^�����y��*�b��K)�ڣ��yx��\sz�R�q��*Ǌj�K����kaY�s7{N8�Zʵ��T��V11�l�&kt�3�v��q	Y�jj�(��ܻ����n1�k��]Nvv,�"�F��z�NS:�0�P�d��:�v�{�Ԥ"º�
p:�s#Ь6���w6�&��{jI����#��鹺4�S�H(Uv9���r��p�K^K3
CX�2���K�.����"�;	;�=\�!yF��j�V��@n[&L̓>
���vZ���,�5��N��&�ږ�Pj���H���L�ZՇ�GVr��㈶��k���H��P@_.�R��6���.��[�Ҧn�s�kX�*��wH8�I��F���z
�Żvz
,���m��	t�	[��b��*���h��$�t֣i��R����X+�i��{|^���#�:���ٰ�95�d�nT�Q>��nu��%��b܃Eء�҂��\�2�um���8���3����s�0H��lM�J�x��[��rNJ*��\�S8j��u'��8���"Ƌ�/�������I[-֞���9�
�{3O�c�t��[�Au~�������X�F�
�ҟK�W؍v��2byF旳N���z�;L�oS��R�mb$�;Fnpl�RwI�f�ܤ^.8����W.u�Mz0�H����C��fe���7fT�<�J��v��Ȼ���A2�aЕɢr�4ٗS�́v;�͍޿@�V�g2;��zx%B��;2��[�r��yf�.zcfp�T��]�p�1�e�#}�X�ἇ@v��u���ym>Jx��ޱ�F΀��v�h��Srl4UұBt���8��X{�0^֤7�c\���N(���E�9_K�\m��֎.��cGXr��1SO��@�y��(���
�I�=Hl�)��)�J��-��+uf���r��:��į@�"���WԮ��@,Z"���V�Q.]��>��UͣpXS���-+��e�\h+c)M��(ԗ���������_r��liְ��=��e�jL\:mZ������췼��l�;Z�v�[���o%I�ɺ0������%��%F���<A��C��&�ڴ�:
�)�w�y������}��o�����?���-��MQ|�QKHm��-y�<��t�V�tS��m�o1���kT矏�����o�����}����|��ZZ~{���:B�H���A�쏑�͟�f��|�Uq���R1Qyg��#m�7n+��:����� )�펶���u�|�J��䷘zM�"o��ռêu�:JX���c���������_;o���bO��#����T�OW�����|�¥��ē]=X���hti}K�=	��
�K�;gZ*�qT�}���	T�R�I�4�4U��1����kF�Q�u��i�l�Q%h֟I:^�4�;b�G�_W��Ey[�C�4I��)��Z��S�����RW�v�PyC�i�l��TѣAlR"H� 	�t6�rSh�՘��.\��1Kuue�ٜC�0��]��W�)<�N��@h�R���x�ݽ5��v�-��<���`�7�@3ɓ0�)�/d��z��.b�|�ᠿGNL*��熫W(�ߊ�Ƒچ����^����]�]|��/Nç^p��l7L@M��]`�4,ߜ���6gI�+ם<�g�dhg�B3"'w,�r��w�*�/s�:j��|�.@������s����ke�I�q�֡C ��>��vY�Ȏ����i�()�Ts	m	֡�aߤ���@�3��� >'50̳s%.�Ƨ9��i�S�����0
XXw�+�k��y�:MKsW�@��^�9�"]�w���|���mux��W�ݴN�zBa�k��s�����O\����&e��j��y��@~+J$���}���L��QK8�w�a+zs�=k�
�T[y��f�Ȳ�[�	A(4��}A�E����=k�}��⿷w�n�"g~�	A���U~B<���ħx����Bq���
@j�G=x%�&�t)��YF�&oow�E�&��}�g��<���}G�Fä�b�h��5��3m����s6��骥�7|m��I޵!���(Q�'�+ע8T<��ly)��f�?�:��a��ݹ�\Cæ��aiOv�^w>�6"LVЩ�vFT� -�Nc �U��2��p�*+z��[�sz>�N�ϯ1EC�8����o�xӿ����g�.���`��ԖOێ	R�x�Y��U�CM]�O餌5-��*��k�NʗS��{�2H�� �7� ��&L ��^���|��?CDa��	�yY�%ץvлXun��zǆ�Ol����J|ܝ�.|�]���y<sF!�(�y�B�O5{ �L��JrT&	���B�ѓx�5�з�tOf'ب�VZ99�Gٛ�c��g�	�h�+C�/��=�2��/Ⱥ��Ƽ��¼�g��>����o�4��xK9^7jb�Cv_	������t|ઉ�+��L^Y��X����D�[͖r�;j:�Ƃ@������~�B��c��P�x�;�������㡧�K�[���
�j����Xy�sk*�#x���;[:i�zz��y}S����w���ߥɉ��\��9��aց@iC�~�t�����#�Ƙ���?�6�bk�4e�FY��fn�2���i��q����W.��S��.s�Qk[R�k�-��pA�Ѯ�	�m��'{.s�hzs��M C�m��t�+��
����P=��9�ʗe�03�(��\�$���M��S�ٻk������ԋ�^��,�2�C��B/�Ǥ�-��LW�:鮴5�!0�L��-�l�V��vj߄y�❧_XC���B��$W �s;��*'4�33&���!k�r�'}e��r7�e�5|�/�S+�D',�^]A�8`ǈ<��[P�K������н�B�yzu� z��w�d�w��}s�ϝ�ݹ�D}���s�
�{�j�v{�Wn�E	u��C�s�ã�\I��^��M<�}3��W�����f�4y������s�/�׳1�E�-��� �}�L����J5׎ǃ�h�ǌ��ܜ�(���yN=�Ó5l8�}w������gv&iBԦ^+(!C�@<�W��Y�ZgK*�>0χ����r��xC�t[ͬ7�
��^6�LcHI*f�;(1���P	���i���"�]w��	˰2`�n�9��(dmT��W=�F�E���/-�#�Pގ�=,SI�J��Fc׭��� v��Ι�B7�zf{���`\��� r .�VJ�j�D �P�Ƚ��4���i5��3��{Zօ�.O(�,��?<�ۧ��.�x�M�jM<GP��[�4���9w��i�[q�i��W�[��qԼQ������O�p�}>�H01�(f�2��f
o�����2ng38�+�r���_uS�oHh�1��hx����F������[y��6����� t���~E��#��sç��޵	���-?,�y�./#����[
�����>�[���D���|j},��u�s?{���ԟe�}��+*t��2��MQV���7(42������L�[����+ ��c�F�<^<�چP�`�[�qw��8��m��M�Q�Z�/��x���${J���rTė'3D�\:������`5�2y��� {%wr����q�����:�i��r�k�2��zԍc^*;�6;�1�Fzj�Ѭ��0�1�Ev�sL�����1s��}11t��v_vh�t$���o6)O�T��-p����Xr��+/;-��Q۪7�܂���09.���<3k�ު�9�Á�F���r��߀"b�Yhx�9��w[ǚ��;�G�4[:�7�q^��Z���:��K��/Q����c���۴.��ur��c��θ���Ƽ�$&V�k�����J:�۔@vfU��d��e��װ�P�	Mn0�[|Lt8��,��Z~��$�2�h��N����Ͼ70n֯lq��aw������y񥿲������dQ3 [�Zz�<���17Q�v��r���b����H`�a��<MG��[h9	吃sRY$5gY�F��-2^�ƛ�v���[��C��zt��_X����,�uI���^l�]'�vOAd�t5�V��1��{Y۲K:A�Ƭ��~������ǐ���la�"��T���=�	��y	�D�w!�"ڰ̌�z}f~���0ʎ����X�l@�:�4l7�8VXWoI��uϙ�n�_{}���/�..��\������q��%��Ӫc�Wis�'h��UҼ+ku*d�[($3l�(�;U�� Tٶ���"ĝ��x�AR[����&&A� �^�Zb,����2����aIa-�rq��.[�<-�Pd]L$�"�Y�=�q���{�2i��Y���l�[�΃�kw:w��T-X�E8���a=�m
�Ӎ�cL:A����N7M��ٖ�e�l�6�@Y2� oQ�ɽ���_���(�%Ɓ�p�;�0���8�6j����_=ע��^���Иs�8�U�]���%<��6Ⱥ,㛖����ٮ}
��m)KY����'��k�K><;{`� C���B^S�q�&̦}fW<5xZ�%��ǜ�[?.{m��GNt�E��9�'H?]4=�(>c�i�q�)hQ����;�2q�߸�,%�vD�� ��U�ꛞ�sºx��F2��1��t����c��ٸ�m�nZ�:q␋~|��dn��Z붻5q�2��{��+7>|G�Ӝ�%Ә#��K��؜���M7Ŏ�N��mv�oe�fҽ���5a*��˦��;�_�� �/@�Տx����+ƇN��~/r�sQ6����
X #K��I�;�t�t��I���v8�	�v�tE��tg/k:�M+Q��Y�, �;����φ�U�__4�`����b>T{�Pêrĝ��u{:��n�R�=�`EV��d#��R7�s�4��3.P�c�eE����꘮p��D^A��V%,�ќuX���U���3�Q�o��Ԡs4,:�)�v"���fa��ə�dɃ30��{��8�eC��t9o&�y/�+e��28�;�e��$=%�za����]{ǎ�?K��Ŵ󭏨�Ӥ���%ϐ�.&3%'�&���fƵ�[Gdη]�x��-v�����B���o)x�T��Ίc��!a�����}�<�j�U�����}%_�R'=O]P��"N�G�={zq���*��&�'�P���!�d8�� ����l�X�׋q���j�:��Rū���c��|ÏP="ySGnH�kݬ���Ux��B05^w��篩	��&�>��pi�y��	L��No�J`��"�]�c���`h��7�;���S�2��|_fN��][�zRM��5wS8yEhpD���ze'E�Z�-�#Iy��~:���i��/U�y�W�y�ۄ�c���ZBvl���sԹ���"Uz����EL/ܪQt�pe9�f1a3v²���(�F>��8�%$��M�a�C�uL�"�У�S���]�TU�e�k[#��vL��u�-H�s_�PX��)ߚ���?ka�~?4��G<�7]�^��B1����>+�����昳���o���z�yP��ʴ6մ��������@=��c=�8�N�l`;u�O]���e�:S7'�I��ʎ���f#;ш�Ek}9G'k�-ӱ��O���B���%\��|[��p*^�$��I�<̿�`���2��^V�O{���;���eRHT]�,`[���e*0��}�����z i�)A>[�p|#[SG�3�"һc����
��zbkζzL�1�kXV��`�%�^S�j��m���2<ϊ%����������,W0�������nf���z@�ǟe]�h�M�}�����=qK�Ɨk�{ݽ5�,�ds�`�������55g�'�y9/g�]g����:���isGgK�Y^���7Ol//o��v��GD��ņ����E"^�Ұ7�?Hͬa�Ŏ�_�^��|e�Y�^��~�Z>@a#��ZZP�,�l��[ѣ����V^[8�՗��<�v��C;�����I��r�>#ߨ��ìٖ�����N���	��]�--	��T륹�Y���MO�^��܋�f�e�[Z����z�e���P��9����{HI�����@8A᧰,ԩ3�`�&������ۜd�v�ŵi�a@oFc���n�3�p��Sg:�^
SO�}w�O�D���l���su� �W�(�E���*w��ZD�s�x�����ҩ�����2��!J�pt��'����Fd뎓���B����]t��8=8;���h"�r�f+�u��*(�|����,�6��C��Ӻ�?�B{�e�^.c���M���B��o������ϣ��}|���\���8�F��݅�_Dv>5'�t�8�M�!�D�f�t�`��}'����'���u~Z�74�Tf斔e�:�"��a�N4g�}|�&<Ř�	ڏ�)��`��h�/�鳯65pl�a���]i|��g<�4���5х�ϸ-� �z�M�y�2yȜ-]|��o����(Z��^�ĥ�l�n��r�O�y�yqyK��p������3�� �9yۚ��B,�8��:���4���s]��Qx�Z���3T��2K�\�c�d�x�o0≡
��",j�GV�@���\kJVvh�f�r�c�o2������{��hy��]wJ�P�@�wluJ1X �>C���.��7����,7���-~����G(읅=��|���=E��A���pt0g��)���5�<�#���@�MI*;��d%����񐷳���l�L(���@{θח^>4��+B�`����X�q�2֠�&�i�U��R1n�4�}yqSy���jeش�c��@:"��E<"]� ��cA>�?�����ms��b������S1�����T��M+�3/�)BTݲ�����wEn<��+kV��8�k(��D�ǁ��m����M)�F.n�m8S��uƥ8;������q�]j�ht ǲ�L�h�و��ٺ����3ɐa�xM�Y�o^�R�DƗ�zl�;�>��4'z;p	N2H���|kO\�o&�- �N�n�� ��Æ@��a�>F7����έi[7�����ȣ:�(=�X��Z曌�y�П0ܪbG6@��I����\U�c�Hu������r�l��O��;']Lwh��� K(�=�Y���CJv���Mv�ן�Z���q��B��šs�k��N��zY��T�xi�5l�U�c�D6룱I��"T)��.-�T\:�\c<�-�)T2S�2}��.��"�U�c�wm�f!3�Z�Ad���s�*�J��]��Ə4���U�oD���a�%�Neэ��3�ö��[,�E�iޥI�����E�.4������x`s3�V���ݚ[���1x�A"}�R��L5�@��ӵ��O<��@�<�5�����m�UH��H����m�׵tJ�d��P�*3�-|�z򟣌�;��
�fW<5xZ�E��[�#Q�U�XY}gaSR=�dO&�}�b ����h{��򨦺�2(��n+���Ƅ��ۮ�]W���'�x�__��ۻ��,�v���N��n��8`�s���/���:����{�����k�W@�g��֘��;��Ű[8��5;�8�����s벯�K6�+z.���me�L���;k̹֜�H"�A�y�����x�9�CZ�^yc���c4'��ʥa��g�
1
��5@0�TL�l�-�>+���mF(�ss
-Ѷ�˥k�*	{k��O�Нnj���0q�<��#c�̪�g����m����o��2پ�a�Y�%A�m�U���Ӕ=ƥ���/E�3��.����s��j��P�v�����<���
�\��]P͗m��Ë�}�.&x�bɗi�[+]3e�vF��}���۲!�]xS˼�J��S�
�T[#b�@�a>ʋ��	I@A��Ea���o=,˸�Y��]��ƔM�2��7����1�Fd��騼{k͍i�p�/$�/n�-�9W>O��}Ht\7rF
��M�S����u^�xZ%0�V��°奼��*�U�L�z�L�����Z-�����Z�2!fP�`%G�=��sO����z>}l�QM"���3f��9۵ֆs�J9������%6�E�!2X�Jx[�(��׬z���S�;)h��Q��n:���k�O�����/��s�	�x�Js~*S�!B�2s���jlM�Y7#)���K;�e�W1�
	��feԿ�Y�]�֨�>	���]�,�{�ˑ�G�]���C�~ѫ1&��4��7-IoO��[��p.��\wd`��f#/T'�ݶp�����-���[����)�Z�*��Fd�AbE5%<�*TtK����Ql����X���Zʳ��֢㥢����.�'a׵�yGyx%&m=�y��;G�j'l��/Ce��uq݉��-rwW�����]E[��gZ����p۹�n;�m�1n���n�(@Hs�:�q�2�PVՉ���q�Ԉ[Ju�Q�S����`C�h;�D��ײ_�w*��c;�+���A�HsD̼�V�еe�I�!K���s�ZTҍ�v�]�%Ee����훠jNG�ok6%c	՗%�nw؎�Cc��V/�kCnPy�Ģ��T;9�Չ׵���^�W*l�9��uwm�1����t��\��u�G%�;/d	�6]��p޺�z1@�iE֩��1C\�eR�Atc����'��!:�+e�۲sc�I�V��@�C8���;��f����
G`V���g,���'{!��07�i��6�������p�d$���ރ���i,���N�!�9��]����n��L�u�s���g�{,�z{\W��\��z���`V�[6��X��@�!���ȱ&���x�6�R��eŦn�P���M$��ϹTu�z����ήVjv{-Zw�h�f���rяR,:�w4m�9LD[��7�KS4��7r�yJK����	�1Iu�u�j^��9#�(Ը+_\��S��ץ�Pw�fL샥Z��[�bh��.�&X/5;�����t{�.�S���c���׷n�'��+�h�X���kA� Rw��Po�j8�n��ze�oAݳQ��j�,��bᜨ>��v��w)f�Ci]`GF �=|�2�r�@�Rl���Lt��������T�;�*}�麱�c1��"U�-�K�u��7}S-�v�CJ�-�s73����
<ξOd�!��8���b᯶N@=ŲG-V!��J��1�8J�i��Օ�_K�}Fn�oQ|7�3ɩ4!���,��G٘�>y�2n*M^���u���`Ų�C��e!�f6�U�Y�D�¢��9VJ�&����6N�wtm�a�׶�% [�J_���~3�hf�!ܯ�E�9s'WWegܹ>�+Okh��.�-J�p�Uc�k�fļʄ$)�N�j���8^�tE�M���7��!V�'&�*HO��=�5�&��U+�9&�)��u�z�j]��I�hZ&���<I.��o����N�7����MgN��o��~y�N!�먴��QN��������r��&-�eB�Gu�����B�k�{Si0��+B+���0�|J���]��ynL�q�Y爨�ZX�M�1$�|�I@��@�AXP�2�+L՛Up�ES
*~z�����h[a��GO�m���#���)b��5I�PX�A���~�����������}��o���'�К�����N�E��&v
�c�SFښ"J������~?o����}��o���~~��]QKE!V즍����"���[c��K�4Нh��"��u��F�'�������]b����4tz�Q�3Q�
7�4�[�vt�i�lTm�Q�i�/[v<ً�u��i��!���v֎;i��{d�B%�;�lGA�SK�T�ֲj��]�b��ODv�]����:�0vɭ=����5��vC�mly�E��'^�
k�յDh-�������.�h��X:�}^�<�fehQ�5�d�la���Z���CE��EQm�E<Q]((8���"�:�UEۻ�A�~���حP�颣E~M��ԭ3�t�m��Fou�n��4�Q�힫=P*�]���cR�ùV/;��5��i���\�W��!�Q�:��U� Ĥ%���IE"�6�.(d��"
"~��3ɐ`�
��Y������pg=࣡G���!�Rb,�_x,�L���D��C�7�Ru��YX9��m7+�i77T�-��ײs!v���ߐ�eǊ��0"q/����O�����]��(�`���ull'�w�\w�V/w��������2@⤨�rp���	�}|hQ9���n��*���U}y٨����k���Z~kAc��7�%�Am�!��B���zy��ټ����u7ǲ���:��ULV��/��}j;�́J�s�O�a�%�â�`@��9-"YDo��a��|�>s���퍒��}�0�б��%���b�sO���H��<!x��:=�|�y�.^�����(C����;3m��Λcqʓ�(�|��}8�8�6��[D]'�F[f.{�O	�Qa��ṕp�4B/"u�3'���E��lc�]�=[5���a�0�������X�'%�)���m������G�s�?��B����K��{����m��Μ��xWݜ�e�P�=x��OT4���l�T�T?c�=����7��|d���Ūh��r,7p�
����}�F.�!��ߦ���8�)�X 1:b���Y�`膩�����x2F������M=4�G,i�=h�'m��b�eh�ݎ���� E�Q*��g�t�\�7^c��
�q'wZ�
���t���IB��O�`1�2f`�2`�eE���p���]45�s��tvJaԖPB��^h����s޲����(�f��+�ϝf�eY���o���e�*®����W
��%L�`�ƖN0-E��3f��=[�Y	2e�g_j�zzЇt88���^�\zUx�c�mEzF��yB��SI�J��u*�_c����zp�VLf[���W�N@|1U��B�$���d"�c�<��@�E�\��q��>��@ě�nnY����-HJ�MvF��W�헕J�c ��"r���c���)�y�7m�"=Mc�͕%���T	b$i5����O�p���l���a�2�����J�k�9�:��\'`P��.�BTi'.�9������z0�>G�d4[W}�
J��[(����v�,mB`�2/���{�.�]1oCo�-? ��	|�R�z+��X̍Mo�˾>��fu���
��D�.(C�z����:�f</Z��a��Gsד��Nsc�N�ۭ9���t�߭��O�(�?��r����T�j���z;����ғ�X��y�N���d�2�^L��o`����P/�f��"�:�EX�
�2F��s��+%�:/Y�t����%Lw=�1T�zr��نݭ�fVMC<�&�|��-�"���M����ڗ�V���;�
J�=��C#Z,@��wU;�݀�}L�k|d�ɓ <���*�6˅�mHT	��;1�`΃�����k���k�ޚ�̞�vd�ډ�my��\A���ԋu>w?�>��Nx�u���H���AZ�!1i�����v�(٢.Hj3w�r�YU-�B
h�
��Y�Y7�nh�鐐���C����s�=>�[;�&���v�zB`&�C6���b�;�h�Peر/�������x4:D��:��I�W�u������ᜈd0da���]P�nWS^C8u�"scڏs��wș��Ƥ��p�w���\��ȩ7/݇{v�<�^6�K� ��2�a�-�p/�W>���S2�H8G!栖I��H�X��c�]���m�؏"Ђ��X�˖�}��y��z`�p	�eE���O�C*�k���mklU��SǶԎ{��{�J��ذ�S��hc�$}��4\mLIv��u�UEV��4��*ETf4^m�Fܣ��؎���N��U
W*�
j�ܜj=����H��N`\鵩�Y�w�[׊����K7	������{1���R2��q��$vE�*��N��~�*fH��M�YW.���(r|?M�ad�����ޡ�Xmʶ�G��X$nj��&*�Z�4� ��y��������T�pٗ��W���̭`5DE�R��s�3�. :7Nt�$JlA@W���z.��&��4�cr�G�ať�&�2` $0���2�#��آ��Ϥ8����́�^��O��Re��&*��QzK�b:p��m��]�/U��c�I]�yҌ�0�p�"1���x�3.�����%<��6Ⱥ���j��l:��XNʫ3U֠&�s���O��A�|�P���=K�~�<hQ��4�UY��Rr�����;Ž�+j;k��)�Ƒچ	��W�ƱD�/�F�Ǽ�E5}S�B�1卩��lh����3ً5pw�y��z�zn�h�nU+�ASb��a�bi��S(�8E�8���r7��V�e�q���{*	{k��HhN�{��	��ԡ��;˾o���]�li2]X�,������~]{v�sW��T]o�݀�#�KsP=��/��3�����P��n��"�ў�: ���o��d�Vl�l�e^�v�rb�������-m��p1�Ϯ�˼ `N��,O� B���ћH��|����\ٝO�6��qoU5�sm��#��0ҴE��bm�lg��`L�\LfJO~�s6�:�b=�go�<���Y��~����p�]�n�����+���ً�=9k���G���t��I�p#���b��y�t�֥as\��I�k7�葼Su(�x�ǦZX�C�+h�}f��(�:��9Ӻ�I�љ����N�ȝ�����YoY8?��Ͽ�� �2N�t������[��e>i(D�^ŸRC�^?�Y!
��H��t�P�E3�r¬8	8�sE�a�Q�3mf���#4�h�C��vf�$�.{��A��B��G�=>5�(dŵ�ؖt6���]�,��vF�����8�y�8ڶf�����>t�b�I�vM=�ܷN͌�=9�����1C+�76�gL2e�A�iėʘ	��E�j�BS+/��R�&����]Z���h���Ⱦw_�G�� o4p��_�{���^}n8EoW��y�S�9��-�w5����k������ô�RM���c�}Ɍ~ml3gW�K^��fȑ=}%�����<F��y�U���wvB���j�Llx��;.˅ּh;��J�JK��G���>˞RVb�&�cN*��C�M'qUiWCը���T5�K�5'��v��A���ev��ڙ���%�,�ٴ6B�(LJ~�OI`Z����5�*�=Z��3t�w*��<��cQ���ܡ�������0�ã��ֿP���%���0���u}�;�W�ό�� N�#8]p���Z����!X)�;eѬ�8ۉ��n�R�ŹMC�ӛ�v�_jQZ���ۻ���.�Q��v#���꟏�����y��tp,�T4��i�/��)E )�y�ك%.�x�²�BgMޓ^�X��)i0Dy(�r�@n	�m��a���2dɘ H�3�{���zU�`xb
������:')@��V#�&!?KގS�ǩ����S(	�eN�̺�ռ� M,�X�;u
����`Eh�^c=ϲ����6C�����$���.��̹�E��t>�py�W�yc�c|������	`��г�H�Se�^��2vd)w΂�$�vZPkXCHJC�@"I�-����0��"Y�!���d�Չ�<I/t�ꅚGN�)m�^�����፹�i�hvo�41y�#���y�P�q\��E'1�
�̘�U/ʫv�wuփ�,�dsLde:�MO��^�1䥛4�Ƽ�s|��H����.m�K�������y����U�c��oz��
.���E��N��np��8��p���u�R�&X�=*"��X�b��J�#k�� �f=���>x[� �d��as	+�A
y�tB	�R��ȦP�M;+�z����Zu�����񤲕mTW(�I8��&<yʘL��H Z�P�����lS���Ո����1��$�i�-i#I��F��6=C��G��m"�mP�vaQF_:��8"�4!�:�N����m�Xk�0�������q�ţ�z��eB����wHʛ1����$�ghL�˱.I���6�-i�w2"������u�y�#5(��lba9��b�1
��8%ޞ��q��-܍}��722d���fÛ��nҽ�������N.�cy�$����g<�5�Xs��=���}�-�
jQO��GGs������ڍIhgIjOx��O��n�����O ��ށ��8EM�py[ݹ��J�8;��1����ׇ �	��^�J=�~�k�EⅩ���|�gl���ǘ��W\�i	��?y�D?c���k�މR���|���ra�����:>�6v�1�����Gg�M:�y���S#+b����ഇ�����)���D��ZڼZb5�5wnk]-��j,0��t��m�MsI}���Լ�T�p���L����㜞����t>~�e�*��e��M�PÔ#���df���8��&+���Z�񐐭NS�ҍq��E��Փ�P���d&Z5:�01�f�}}�hMq�.��]�O����^��6�zn;��,ٛ��<��P��B8��8T&����l�9���47����L��j�:���naf��γ-E�)i�~��<��[� ��O֜��{}�ZҶ
(��N[BǤN�j-η��ī�2�S�+���7[��A�ۏnGXh0[tMm�M�;A�����*G�fot�A�.:Xo�eq��Nf���u��Vr�(.��L�(TV�������!���4��sr�ë�5�V�t��|@�z����� 		�rv�V��:2�A���¦�(��ΞQa8���=�����r�l���6<��Ok%[�� �G{5���(@��%�����[�\�C���$.��<�>G~�<�Z���_�T������56��:Q2׿P�PX�R�%>��{�0R�̫1����z�W�R|6nxʞ����ݝ��v7�_��'_�7tBd������R��RS�|�a��m�kS��ʭ�/4�l+�@Ky��ć�rMl�pi���*�"��y�ޑ��c�L{
���{ئ�O:�t�v��}i��B5�C���@��c��4� _T���)�t��X��؎��ff���=ܘ��5|�:�*,x!�(�\�ɻ<V���ŭSl%6V���W��*��vL���+��a(,h.5$'�A�nZԄ�!q�,�jƅ]��n���=�x�_��ь9�̄
�t�qv��­t�y�R�a���8x\0g!����F�|���`֛����]�U�)��d_�6f��q�Z�
�^�������4��it���>�D�nԎ%�%5}���D��:Ů�Ƒ�%���侃`\��-Q��y�[x����g��m��-ԩ:]��݈�S)��8��+���߮��2�Ǚ�v�
kvx�S�6�m
ح#LU�egj�q�L�5!�Xn�:n�n���Y��[��k]c��w����&dɐ`՗�\�=���۝��R�i�~'�����{��r+��v�g%@�.�ǰJ�[eT�j`Z}�պ66�L6��[A���]�u�
�pOp�x?R�[B�%�^4r^�^"��yP�bX~��6��(ke�^����=��pzlA@�r��)|<�<���Ƞ����m"/���q�FQoq�fڔv�u�{�'��zm�OՐ������'��d,z�x�֡6lKk�R�*6�������#�yҸ#�槹t˦.Z�?0�|��4_ȻzS�ݹ�9�{^%�b����q����R̠i):��6a\t׫]�ݜ�2x˙�����CFF��|z���J��Xo	�yHL�)����z3�i��.ޗC����F�����5��!�;�����4�|���L��%9��0Ms�}�t�wn^k+*9щ,kxb��\ب�Q/o�����y�V*`$���|kӽ2���O!�6�)}7V�Q���$�㡦)��G�9���+v���N<��3�ؤ��x1�>xN鎼���U��7��[_fu��B����J���{��t@��W[��+��ݏ��e[2ݺ�kj�.v��c��,2}V:�~X��]-5{[~	H� �V��n�P��-�Ac,���J�2n�2m�v�L��\�E���eJ{�2��f�6 KP���&L��0���{��ά�]���V>���My\�,O�AG[��p���L�vaA�Bm�И.�=��[f��t�b��泪i�p����r�O�eCx��R]���ı����)�~�ӻZ������i�$�w^�vB0Bi�_�jy�5g-�v8�0�}cH�t@�^�Z2��t�8��5�;+�uD� �����Z�Ķ*�)�Gu[
��e@��ߞ���'_n�zl&Ũ5f��5 b�:P5t-����7J��أ�Ͻ#d>r�!^s��2��ת�yt��,��z��X7�h����:s�"?,��K:��k�s[;�v�:�θ$�{q�h1�\m�s�Ӵ;<k�4X��~�c��|�	��/��6[s5��_�%�^$ƾ�Ǎ5�!����8�	ꆐ_E��lEC�<3�B5�k��^ј'dDO#}g-�M�~�ΰ��g�ג�u�L�;X͟�\�4q�$ȴ��6��-�Yy�}�y[XaWi���i�׸F4��b x�s~��O=��`\�3P97PH	������>ߚy.2�v�^�.��Ƨ]�
�N*�,��R�4k5ء|ܲ�Y�w�����o|_W=�/s�DEZ��&���w�-�6���JX�P�Nn��յg�s�7&m��������)�aΆ��f���K��U�4v�7"�eḑ<3�,��ް2�ԤpvP���j�	q_CXm�{��h����T�J	�����.�@�/u֤�`��6�`-C �����šYO��q�������3!���s�b���]�����v��FL���ɯ�4�)���%<9�2�J�+m&��ӎ�s6h��\ڼ�q�'�Ww��ov��'u����J���*�v<(Z��qP���x�39�kq`�Jb���PO�M��ܽ$��5γ��r���p:���P�O\��&���2�IȆ�N�YY�35XY��A���;�:��B�	.5�(�)�;���vf�����ie�*kd�og4��y�߃V�]���`"\:�et��>��G������u�կ�G�2��ډ]����f�67�7����>�x��d���[�vk/[�A��+.����D*M�Ʌ�c ����n`]O\���YK��JV�Y�8,��Xsʳ���c�CF$e��f����tR�i�;��iU��i�Iȧf�3�Jj�q�*�3]�- `�[�c�$�*���޲K�ɰ1;Ir�O-�cE}�6p\�=��5|>s�ad<]+:H$���e����eyܟ;����ng�#��N��
�(m�[P�q�:�c����0��soI���b���Rh�Q{��^ҭ�EX]�G7&0���8��@�Y��v*�
�9]ûw4!�5ȝ@
ۓ4�\����0B5sjũ�8�EĢ�7�4-��<�j�Wō<��6;p��ʏ����9��\�Ym-D1��8�q�Jݛ.�neM�ƣΖ5�[|E�+si�˔�I9tCyľ�&�޺�MRHr���Z�5�%�V�f���{��t���F�ٖu(�}S#�5t�@�L����*��X��m�vi�Fg.�3[ 튇��^��^ _N\p��sZ��%��v`9��s�H��,�^�.*+�Y�f\cs���쀮;�tET =���caj�8��P�qq��f�X�)v��r���W7qdb���	J����K|�Fh���ڥ��E]-��j� �b
u�Zp�# K��ˠ�i#�gg-в���ū����PVmw���sh�T��9-\�-���p�sA:�swc�L��Wi�"Z-st%4]k�(�]M�Y��Ɯ\��^.0\4k�6eI,�r�&��`��j��ci�Z:Nq����\]p�oh�յ����yet-2ch�%�6���*wq�/Q�)�0^��0�9dj9V��7���n����Kp�&h�o/����2���r��Roo�-Q���b��KB����Ij�5�UT�W��#�ƭ����'<�}>�o�����o�����?����ص��:t�����Ս�N�9:�c��'Tt5AON�3�?O�����}����������?5�::^���ulyEFڊ>PW�ѓE[�7wv�d��"��iuC�@o\�m��+Zb.�<�#���(z���y�*��A%���֝�E��z�!�EkC�*�V-hi~�零-c^�1���BuZ<��y%ڊ�ݎ����>TDR�I:��4��DZ��\f����=xj �� ��$�HR���@��=/A�Plh��롵�*��:1j���u�M�}w�	�&��Z(�QA�Q�cj�v-Z�"�*�%th��b#cz�;e�n���D^�O� ���(�	l��{�!\>��y����ղ�bkV�j�n1%�yN-�r�M���`�������O�}��t8�<-t#��.Q���?���"A�{��y�1g���{g2�S���,9/1q鐦m�7쨯H\D���(2k�����/[ei�����Q.�l�
�1�ޭ�=[�:
ȱ��D��v�{|������O4�3כ���^�
SL�Q��R�CEd�e|��V���?��&�G�O�ִkAi��>ܪU��G�oB,3��(��=�)ͱR)���&�}������Y�זq�KF_yl۬��t�n��~h�3FY��^���[��T��D&*�<�T�sj=]���%��t:=�o>d�a�|�1���@r!7C�m�^Ȕ���[�IߔR~D'�Z@[�#z�1]�{~��ܫ<�!{���[AF�<5Q�W�sX^��qm/-^����R�L��8���_+o�S��q�/]�C���ܣ_�a���(�z;���ꘁ·m����]��8^}�=��#�;�D��)��s^�-.!��z��猞��M��Ff��c�E��
�O�Yc����:���A�#O�L7P�`�4x�LX�h)l�hf֯�w\Z�q,X��q���&

��`�hSL\xϻ�,\�Rܓ�]ݪoq�^����/���X4�i�����V�6Sj;�Þw.��hm<{+�SON2`�{��l6ΙvY��\�&����0�m��o`�$U��v,�b�@���ӳ�쾓P��*������'�t�
��;	y���r��_�BA�eP��} I�޽���{��vC<2<B�W��Uf�}y�hP���.^�꧲Y^�y�D:��,���ٶ��3V�W�w�P��4y������֜߳gח��;�uإ!�bpAS]���EtL����{aC �Yt�O�f`0&|�[{�d^�}U���X������q��½��`)̆�O�I��/&�s��<'�%�Տ!V�(�ڢ)˃�Knt;�yy�n��f����孚����@(��YX�]ZW�Rq�^�5�~!t,9�r�f_09n���;�gv�q��v���d�箈!��'L�X���R�aMG�q���\<��?0'S&��*�[����-��� F������Bo��[��1	�{���J��Rs�g�gX1��j�'���]w<���8ޏH{h	�'��2�+e������oF&�K�LU�Ȣ�)=�3r�X�{�-�^=�U��S�P��ł�i�:O�'� ���0%�*���}�}����\.���%�.��R�[#��b��i���7#�5�XYx���� >� k���~�T��p��]��l��Vk�^���__sq[�$���r0�j��=1���i�I�Tp�3�̶:�������z�B�F�����l�o�;�O�����<V=�Y]e	��~ޢ�=M1*�s��{�_�-1�T>�P2G�%6�����(<�H�=�DS?7Vq�Y;sqJ��Ѹ��Y�������Q����0�3�������僦��	���Ô�/�R%M]���[�u�q�P�+]�*�]�M*��i��*Ai���(bۆuל��soXR�Ʀ6Ƚ4-Xs'q�X�T��%G0�a�X�b��{��;U�.�3���-�`��3�1�"��̮}Y\���e�X�	N+�J�bІ�z�vu�G|��k��"q�Pg % ����H	��mr{�5[��e�Ba�D�s�����Rms�=ԝ��S"p=�qEy@�	?8v����r4���"��wa(���vjU�z4{9�؜P\��!�za�胏\�ok�����<ˌ����Ml��T��X�����f�gh�9�/r�׎Hym��^�	�Jb+G3�`l�:�PS���n��g�7��v��p��6��j�ن��ܤ.s��%w#�JN�z͜a71P�J_u��>����O4�s���q��N�YgKe��u�u����dX0�,m�٭;��@��чs'�e���x�Gc���]�6��x��*Q3�؁�V\q�����F���{�c�Ŋ�@5��s����N�`�y��o���=�l�(g��
h��iBs���mT����E�;�G2���'�]�.e�^�?]�(�W�{=
K�1M'0%QEǆ�� �L=�L;e�V��W����Q)�@���k�Y+3�wr�'̺zET�6���`J��]����'ʾp��9����W�]؛]��^�m���G\��,���ƒ4��z6/�9M��Pc���v���P���U礰����+�����0��U�ac�J.�s�1�b�F:ܵp����%��T�b�;��ջp7!0u�&̧pE�=��?7>����%�����h:�z�6��s�\�K���f�7�4�*��]<rya�F�޸=�!��ǸS�����2g�����:��ޝR�Н���c>`���ֿTĶ*�)�Gu[
yJײ���v�E�� ��Ezo�f��7}���,ʼb�>�d
�p[��.6�!ݒ�{y�ئV �5�h;]�w��ywt��kL�qW����{j*�X%h�����GNy2~V����-ا۪��w�kvN�w��Sں�d��VB�m�R}d�ovN��S���&��_�-FZ����}�sӯ��׷�Lp�xW*?�	�Ȣ:B<M؜q�~[be�=�Af'�^S��ڧ�os"��'{Y&:�����5��s�
ɺ&k�`��+��&�y��{b�.�1�|��vY�z��7ۥ�T6�z:vBF�:N���]��شd�h7%k�g��1G�q�]:�M��h>�άa���qhIꆒ�-�>؊���v~����(і���������C\YG�ܲҝ�������&$_Ia��W��$^E�1����L�cQ�=�Jeᐧ��|D�KH�`C�Zs�s|�1�#J��:���a�n��{����WZ7��#��r�t�|n��Z�MԣP\���a���是����B�%6�d�����ϵ�os�ݻFCi�O���c�kݩ�5�xJZ�)�s��������5C7��[�^v᝻㍎�1�/y�)M2�g�S�ϟY���Iz0�Oțy������љ�^oVY�ȁ�r�عwMI˼'�⧼���Mmb7$Od\:�:=�=6�flF��vUv.�����k(�,��������q;ԩ'����~k)M0��z0����鈲��gG/:�<���t!6������i�,�ׇ(���'����z�\ �3�:,�J|O�F#)L���X�ŗո^:���k[��v��h�sM�X���AnoW[jɎ�a�Z��� �Yz��(��W�jZwZ�	�FQU2��cIR��'Iv�̄�wQ��.Q5�oA����t@����y������WF�4���l1D;p��x�-=�#^�)l��k�,� 彙�ݩ]F���<���,H1��/]�C�c?��ǌ@�u��^fn{}7-��M+h��9���V��x��]<^n���
���vh�`΃�A��}��te���E-�زs-k�Z��K��y�+�c���Լ�s�C��!#��\����0f��0q#��=aKC;cw:�l�F��ғ�a�M0�M��1\�~�,Z�����36���x����b4E3�0t����ƽ}��( ��8r�0[�9i�]j(|O8���u��c����el�����)��LLG)Ԛ����Y�}6���-�o��,�G#��͍��"C$va�'Ʋ��6���6w��>��f@p�C���ܫ@ڼ��͋5���4���œ�W������t8X��VIE��4��c�c:y��#E@qAv�gUJH|����Ք��OϷU��[#7y� o=7�k�'-al��p�]Z�F:�M�T9��̂qs��|7�!`2�
���'�mv��B��u�o�.�<|73B0y�w�?x�Q���V��UQy���1zǪ�"�x����a^x��/?G�x�~Ą���W�Ǌ�3��N�l^�֍��m��M:Q�\�G0�`�o��q.�Pp&����~����v��r��� �wԲ`X�n��y'h�Ƭ�j�#��;>;wE���1���,}�ҙ\�J�*����ܜjQu郥��a ���W׶ǧ�K>�x���GH���N�{#���M�C��S:{"S�)PN��PzƩp��<��x�i���}ܺ�0�QmAN7�5��@q C��}[,�ozD��T�p��mX7Y�!��`\�9�{���A�@U
}z�,�Rr"��f��r�q�k\K*�4훓]�q`�i����Χ�̟]QL��g�k��vk���kÇ�A�Ƿ�\�%�s�4���y��Q�Ӈn���թ�����I��������#9:A�mе1؅�U�.m��D�41��7[=���Ж��^S�N�qH���-t��R�a)�sӇ�;�6�5<b�u�L�_]��
��I��p���Le7����8���r��������Ǯ���E�.����;�Sx_�,�[ ,?ġ���|�'�VW0M���C.��oX�"q�Yw�$TP���w�8�o)nn�μ��9�!���SC��!�
�5y?|��h������~�Q_i��#}(��Ewx���d�m����gtݪʤ���78f�k1�.��i���xt��u���/%�r�qI�xS"t��@�8.`[Z��՛���jǘZ�1lr�ڭ=N1����,���Ñ���5��x7�{�i���x���g�9ݶ�z ~lh{�[9y�<��\W�>/R����+��z��\:�3�A�sXm�az�м	���(4�'����x;3��3��6>b@>��^^�sn�LUW�N�B�t$ŧ����y��v9���HB���4�e:j鋇��,��DûJ-T�+&�n.�������c2k�I�ږ�{���ǡEVW�J8}�l��o[�]^�rk7�OK����M��0M=, K���d���W���I���P��tωt�X�����j�27��U��ji9�TQ~�c��P�B!��|���Є��s
����K�z�����O����2X&�#��T�h��z+�J��]�.�V�w,�=Q�v�q���k��u׼���������)�FS�|�=�R������`��w9�ۧ}˘�G�Z�����$tٓ@DPދ.�^�*Qu��)�b�@�[���k�w�8��䨒��.�(Eeӧ{�E�`��#�hI�X�^j~��\�&ʞ���/|���*T�~jN=��7Õ��mƻqVͭ �Y�v>�W�D^�F_�W��+ʇ/�a� ���!��%�.�Ju3�Y|2u"���*G�>.����+�>�ڽf۝˛W���JJn�
њw\�ZX�ESP�ìsT/�y��B������w�wa\/MH7�����|�oxl���q�4�C�y���昱�	�ۮa-Y�h]�Ta��k�C��0�Rm6U���N��2�K ��<��Ds���ֿTĶ*��
e_�uY���Wè����>QVu�����>�Y��T��!n-"��q|�@�!Զ��5j&�(�UW�!�Qױzo��N�Ά �3�-)���X1�=�	��P(��:9?x?�����dtq�������d�ݚ'*�k��B=/��._��7�t;�~��3d.5�G>#)���B]���{�œ�~Q)O�k�p��Sܾ7*�g�Ռ!�z	\Z�%�\��1�>芇�	�S�1�ѫ���{W�{{eC:@���ϥ5z\�O^��U��uO�M��3MoIa�\�����:8�`���#��[�1\*+����P�,>0����j�^�P~��^�䩚�97,������_�j�Xsw�V0�=��l�z�κ�Շ�zE�3l	���56�y���Ņ޽��[�(1jY^��N��Fb�-U��Us�F~�|�Kq��	*�X};�Eg��<�62(��|6�ۉ�&�e用�vb�a�R֤y�0Ȫ+W��:�{��xfM~��0Hv�xkO"�Q�<2�r� o��zu�[�H�Û�`u��G��@Ӻ�c�hֳu�Q��z�32�@�:����ò��<-�|L�g�������~��Qj
!�(�`�QN[nJ4*�v>1jg/�����!��^�sL�������N;6E�YG�@��(�@��$���P%��� ��kk�xN�
틇Q{M��,(	��7���p� ���Y���&�`	�Ј��ԆoT�2O��'���S�5���J��S����Q�[�s���*vO�D;xpvvDBm�1Ř?WkzD��(v�,���-?Sp�4%�N��qR��X����=��k��Q������>zc^�C-z����"I��:�ΌKhf�n�m�w�?o@㮻����iN�q�E���wg�?���a'2�=�۸�lf8Bب&����O>j�O���|��s�I��7q�����Y*m^������k�B]6�u̖@���}����ye���٥�~�H��-�v���{��E���7�b�Z@�^��I��,��;(�5��Y�.�=�q�oD��w�2ԇp�%�<EzSCH!@��
�,L�W�mא3��l_������ɲ�1�����>�f�����u��(�[%�H��E-�o�\��J������)�.�ZU2V��e�W۱]�[Xױ-qe���-�7�`��sX�<+�ܳ7(W��˅��&� �uVIh���5�(>�X����z<��,�8E��y0��PBH��X�!�λs������p��8�oF�10\�-�/v�v��z�!�87P�M>]w./^:v%���U��U��*���T��wX��*�{5X�cZ(X0qg]�]��o�',�`�(�9�Vb�K�T�*�<��n��W(\NF��I�,��Wô�ͽ�)t���
 ��/&�� �O�@��]��D�O�`��۶A�2�f���f4&.C)�B�t�{�0um�襾�Nm �G��_
�6Ȭ�i��ؘ���s�9�Z�[RfV��:�ʾ,�!j�uf�5sy�`n�ز)2�Z���l�Q����khe[�4wk{��]J�r��T��oml����9{�;M���7�7��&��zv[��h��f��Ws��cnY։�|��t��͆8@^.ޝ�n��%ݦ[(>����<I	,K4]5�!d��v�+�Af�^$vH,
�j�z�O/4x��2�]���������.\�k]-��a 42�BN�}������s\��va��\��S�2nZ-N���H4y��Bx&X�K�-�⢣7:����QA���\k��t��m�D��F�_3��(�.Y@!9=�i>�D��LY�G`�����ͪ��0F WV�׆P+C�������lu*ͺ�X�&,W3���������&�(�W+�g$���5���Ɉzk�H�^P��r�.�]{3I)��3���]�m��V7���FL�'P�M� ���Mgs�3���S���������h1|6�Q]Nv�&ك_i���������7Y����&�ɁRD��M���\�i�W]��lE��࠻*��BB1̛s]ru1_���!B\�c4�kVHC�FJt�sT8�#woH�&;�.�{�T���;B��D3$��|�E�n�͢�U�i�2��RJA0ۗ%���
G��x]�X�j�w��&ҙ�J}6���@���|�>��]Nh�C�C�5�ܭ(�� D�0Nev,��iŊ��Y�%���Xwkx��!}F�å��)Z�9���d����wKE��=i(���D⾥��+��`�;�.h�S��;*�%���̻��3o��7�]t���'�� �W%��Y$qU��[9ajP�dg7��+��م��3���(c��ٸ�����r� �e`9�:��������@�.<�<�ko��
׮�>���HM�fu\a��X(���prb�}�g�/g��u��6�O/+�ϳڗ�������5�ڃD���3��r��d4u�MV�5��#g�7T��@X5�^�` � {��������L��X?�3�0���u@Q���^��8��c^q�����j]8��A9�����}��o���o����ϑ���d��<���{��AN��ͱl�Tţ�ADMu�1>Hs����?�����~����������}��3ݴA�5�����uI5SG�ۭRAF���"��4�lN5a̽۫m[oQݧ'���j���T�z݆�2�CQ�]h�z�;Vε�J����A۹���׈��m��̚(*ŊtvwT����U�B�]��%�<ؠퟩz^�g����M;`֐�E[=��m��m���c��ɧ�f��M�Q�0k8��:J{c������`��Sk:��)"��i���4k�;��ޞ��h�V6"kF�6q�-��w:�ڂ���5^w7gA�I��ֶƃz��U�{����a����E��V�Zgǜqq��f��C��������y�!��w9�ڪfZ���BzMg�A���^�2�����U��H�)S��Ë�������t��;�;gz�<0Xq�ch�!���$�NI#�4 �!���� "?~u�?}:�oٝt
u�����U��TW��$�pA˵�j�2�/ܥԚ�����f�DVb~�����|�[;��G; ;�pi�=,�ᯖr����py�TA��ݟ��U�Wv�Q��XTp�s������l���?����a-��R}y4ʇ@�t�9��=`��������gc�M�ks�l�>�B'dw[V\z�.�����	�,�,k�ukE���0����6#vl�7(t|n��>�s�H3�r���ٌ�!�>�As�BeK
V%W0�:Ŵb��	?UeU��ZsneL:��cƅ���q6!���YD
��R�ܼ���
TĦX�Q%df��W��N�q+��)/�ز��A{0Ô�Bx���n>��o4�J��.�=F��њ��̩�f?����3{��r��z�-wʀJ�2&c|<*?�\���C��'�-�y�x[���zwy;!�S��䢙X5q��`d��'T���A����aֆ\��/y�y��q�r���(YT)X�I�Y���Z�E�rĂ��r�;�ıXA��,���#2��y�T��(ch�����səۺ�YAJ�ܺ��y2�-k�����S���i�\-N����}��˽��[��-+��kJ���#��`���f�'p^\�Aa��@�4Zo��=��w2��n��	Z3b�eͺ;!ۛ�ŘFj��j�e��@�I�^K�
��a^�Z��2X-t��U����u��Û]4&z��:ku�*;��]�M����	�Le7����ua̛qC�H^ʂ^����fϝ�;��-�7���X�K��a�@8?į���ߔ���y�m9*�t�=�#5�:�\m*��ͭ�5hM%�,Z��������Ĕ8y�Ƈ�&��X���P^4s���Z)����c�,����4�k�݋�lw����,�)�%ߠ�&г���Ϭ�c�%ϛ����M�/ՙ+[�:]�[�E�&\9@!�� �0؞S��pO -�_%{������{�ސ~��������Q�ٯM����Gdt�5�\e:j1p�bj�N��Q���;�j���\�b�h��@��{R��)��B'�2�x�J��~��c�4Kg����������1P�^Qޤ���:��Qx�ֻ�f`���c	���ɧi�M�m��y�؄ӡ+��.�ǯ[ռ4�{gh�-�k��H]>���נ�z~]������nZ]|�DOe�X�WlxU�b"���u�[Isx�5��ҮU/Zt���g�X��՝�}�N�&�J��;{{���P�Lu���r��M��!�mM��(%���&_T�Ya����j��-d�z��|���������љ�PUS5�_Y��1_^�m����9D��JoΊ��V4\])lTW(D=��$!e�vs�Rz�v�;9NͷT��z��}���Ju����^4��(�䌦�_8��s	�\@.�qSDٸ�4e�d�n�u,�R�9Թf�H�ҝ�z(�a~�R�����/�jxM�[�U�߫;	�4�zs�T�oK��BuLm�{�)X�I�O�
�~9��ʟKx�����g��~t���77v�ؽvw�`�5�
�7�����ç��ɍ,4�^�P�Uz�k��2�lj�=Et޹�Wge
�@���Ӈ�p��a���yí~�1-��P�Z ��+��:�x�>���*�M:�()�^S�U2͕4�d=����X��?�S�GW�-��͝D�v4<MF��9ِ���v��<���z-Ko�L{&	��AG`c�ts���kC��I
^S7@�on٦�\!YX����[@��iC&���F��nf�"��߇Vh�<a�=��S(.��d����>����`f�!��8��>'����oR`hԄ$ƌ�7���y�J��ͭn��-�0�B�R �K��x�1�]����M�FQ�W]D-a�3����P�3��c/�t��Sۯ���vaۊ�~���󽂯=�k<c�Z9fJ{���[&:�;��K��:h���������a���	K���٫=�μ�C���S���/�O�:��4��ג�ח��47���	e0ӱ{.vN�d�Z����0��/I��q���CP!@�������y�^�4�J���Ѻ�dhf���Olu8T�b����Iuފ��VW�t��0b�ho˝?����f�᢭l�,٨�Ç7+���"u���5�%�%Ӭ(�f=[ռ�[� �]z���5ԭ��������VR�ro�w�R�
FA�3͠tA	�r��:����L��F��P�t�On�/{�U��y6;z0O*5�Ȭ8@��jԸ�- �Js`�ƒ4��==#�B�y�ix�׉���e�U.K�z�tƘf�~��Y��{&�+z�$���%���yU��
�d��Y�#��u����b��4�=���=:1�XB=D&������ ���Ϻ_����T�c��{�8��9�H;�#k�f�w8~�E�A>�C ��C�.z�3Lz��V�(�QGz�Na��
�;�jBc^*:=�A>;��FՔt��k�:��G��E�OI$���]5V��N��ɔg�	I2B�Hд�U+�V�!�q��5u��=��+yR�=���؟3Wh�PQ�y-��`n�AA��j{�:�'6���U-n�(�+;�k ����g^S�kת���B:��������ɨ�&����Te$�p�Gy�b�3
�Z��׮�'�V<7�6��X�����_�1��?8$l��BEv��Ds����r���./�.~a���=0�u�o�+�s�)�^�lr^�/͓��BՇ2Xux1�e�c�a��_��,]�v�b豇$���>j3�k;�f0t����9^r�.�'�.�� ^�Yғ�a�M0�ɠvQ1\΋�Cm���y�NN�~����H|12�h`�7���#�́j��A��#"[��ؽviǅ�g��J�a���OCU�l�	8r�)��H/ܥԛ�3g�l�ж�ʃLe�gۮ���%xb���T��l �5��x9����	�"���["����N,�Y����͵��dW� �栖I@�!�^M2�WˌJ��Kp�_I���}O�{罻Cӝz/MQ7��ɋ�w%�;&� �֐z���mRE��u�bmd��ی��#�$E/! >�-[O��B���2h:���lQ�{4�"�tE�F2��M<zi�j�eeD�� 
պ�%��#�ǧ��u����m:*i��:×}��M^Zj���G2f�u��]����nR<35�9D�6ӝO�fc1T�*f*{wa��v���X*dOi��&)��9[]��N񦅐mv�9ze��s5�T�����rlp�m����3�b^�Fp� y�c� ��������9ަ�Y�ngݙ/`$�L!qZ#�+x��m��N�����/������dx����	q��[>j�3���.�#Dd+fh���7%�����k��aM�)V�\o]\۠�����§��6�"n�3s�ݙ�w`vq���z�U^���J:Wt��I����4q|�[�Y�ݣa�tw��~$�����i�ҥn���e,����f�R�k�ki���E0#�uGb�^�U�&��ueq���25��fJF;g/��o33v8�d�wӡ3�`����P*�N%՜S��������b����d[�eH^}�4l12�p-g��~d�s�Q/���W_v[u��A)3�-�>&#�WO�۞v@�/W]i�._�Y}���I���[`^[��<$�D�y��=~<�5�4���	G_:��*X]Օ$��E`�8��ɿv5эw�@����5aCn\�;d��붞�#4L߉߾@+��cJ}�{�!cV�h��Y��(eZ�]�	�K=[�19[|$�2�%��v�`3)`�x��l��B|�Y�q����<�bb<=��v�K���p���nVf�xH���6D��ג��*uYn���rfv+�w��D:��� ���b&:k"֢��o!~T��T���؄�-�j{h�֎cV{U��Os�������J�Lb
���54lD,��gN�)図�k��v�EM9��p���������!��1Us�@uk�
������n�
x�8��:x�w��)���v�@�g:�#5��I��[��j��˾^�4Ew 7����Q���/���Ǭ��]:���r� tLw�k�����
|��T���6>���Gx�^z}y���jU���Wy1�7L�Bl^l#�A��j��*�mV��ME�d����x�j�ܸ���7@aF�HRGO��H�$���{�����8�*Aޮ�){ϲ=���0q|��;����#���+ޱ��6}Ϝ�E�W�H��/{�ǥ?l���5w|*�e�X��շ��#�v���]d��׳�klMʰ��ۡ��UdCL\hv�kxU����D���c�k��?//����')�m9R𞕚z	dG�cػV�O/���P0�<������9�O]�sz��:7��D�T�,*�Z|���3���`���(��.��ǳ��s�{�.�=];^ؑ���Ң��@d@���CG5c"��]&W�-�'�9��_�����o�3�-�T��Tu�eY���A��
�;��<v#�)G����U������o$w��ь�J~�$
p{��re��o��tl�2�u�?$��(�W�"��D��{1��&����@��M�^��5��)�
rYŎ�A?���OOU�6�����tk�8x7ewgp�4�GJ:���9�Z�/V`��Q�S��Y���]�7�Q�����M�Y���� �2
]}��eĹ�h*��3H�:CEn��
Ѓ�v����@��(�)J�B�9Uz�Ծ�%%�.V��8r����h�����M���t�[�: �xqTh$U(�Oa�u�e���ч� �Uy���a�&"V2
����VѧY)�u�އYo:�z�<
�-������+�����y���񏶯�
,��}�x�Ҟ@Y�������b��#��Q\+�gL�*eΉ�"2�%<�y72��U�a��j(�A�<s;�mXm�ގ�������2������r�?�T��@ޔ��t|Zbf�8V7\5�2^6���w;g��ʺ��2u�uϠ �C��c����"�3���C�;��vg�tfwgeJ;r����,����Gst���c�F��-L6�Hf��~��ù.�7��3>�u�`���vmhf��2�'�	������M�dF����⦖�E	)Te�7t8h�#���%k<	l7To����
K�2�ټ�/M*�xW����p��\{1�����V,�[�9P��0>m��#�V��|�W��M֝��7v����Y]�9�{cH~�������=�U�#�U����.�������?E�I��v�;�:���ܧ�.s�OK� �}	Hy��7t���Sw[Fִ�u��;ٻi�ȐI��N�I�tI���Npha`�y	�z����06�y��u��e���|)��9S� ���}d�-:�,��*c^j�q_WNK.]���2��с�j^�y�~s�T���+J�y~�hS�o��Y��9R>�E8Լ�/���U�ĭ�8������M���-��vhW'T��y�=���o{��^���M*�셜�W�䨌+�\+U��t��� �ֈ]��ǲ0iL��\�T"qɋ��mvdRhx���׏]�P�_r�q��Úr^�2��߂�GrWO9+�2lɺ�*��ldo[v��L���ڳ�(	@�d����Au(7 BB���ղ�ҧ�������K�b�44��M�������Ш�ċtH���գ��O�Dn�͗Y��y��{��3g+��EsCx�	q;mT�2E��2/ *�?����>	���s������I,н^�z���t��5ё��d��S��������s�ե�ݺ��@1\g��*�esȥH׊�B��x��+�n輍�0��gL�6�K�tw�!)�͞����Z�0@���շN��Kj̦�퍛Gv����L�k���;镮MΝYL�<�c5�;��tӒ�v=0�w�dl	{-K� ��U�t��G�ǈ��PY}���2�1ۥt/q[�quG��I�O%	���N�+����w�qW`c�*����G5�r[�`ZW�G\���<x�1êC%ıZخ^���OX+!y+���os��6<���r�ux�S���N�]���hoD��{V�ش����v7���&�++�-���	�D��۫μ��ܵ�Ƭ�ud�*�em-�]消=#͜k8A�e���%�*j��6T�i� �Ӷ�V�X.ͅ�ֹٸ)^���Dݎ{"YJc�¸,�I�/S�3�T�K�c���e���-�՛c| �BWd�ֶ�@���1_uɛ6�%�<�Қ��L��|�S���x/�*��1'T�ٓ����es���;�!T�vf�K���bٚ,:��r$�tM�r�b6�T�u:к��Z�&��֫3�<�nu��]]d��A aV�����.f���vմ6$�KNHq��V��k�uL��y��q�Vu��%t!јRg�H��6uv���2f�Wd���pH^�}� oJa��"n[\�nj�Np��x��oP�X/$�����o�G�hRvej�vRyB�N��� wV����{xl�����Zc�9�+jX�� Ւ���,�!(h�한 Rq9X�%h&r�gl%+"�¥EjM��:�سK�ԃ��w��(��i4z�"-Uo]�(fdgz�����:3�ٰ� �u�v��� �J���0+�R�������w8��+;3��N�})�h��ȰTb��Q-:��Z�6�X��כ�>�틆��^�x��k2��u٬U���;i=�����OV���e�n��o4n�0.�sQ�@�uER��7�Ȋ�����u�@�S� 5BU�5Ӹ	�vM��� dдJ��2�������bQ��E@��}�Z`�t�M�i8��m�奙� 4)Y�EJ��8��[e��॑E���H��I��%^`�{�+(�eՠ����P�zJ���(YPo}�.�y�!^w't�|���]�-���1H���m� �A:8怹lޠx�ܝY��8�@��rJw��Z����Qm]X/xk�m�t�����\{M�7&��0����@h�*u��w6(C���u 7�,�=��m�<bv��[�5�(��t��6޹2Ǭ"H���պ"�ރ&U�r��(�;�+�j�t�]���eZ�2l8'G�����	�=)��W#٨�'K	��1��cX�ْ��#�����\��m��dt�39ش���]�R^�U��:i:=mnS�py��O<�Z�:۾�trl��^cNNخ;�7��x�h �lR��%`��u��a�2�l�M��=���]�Wmq�mk��Z�.#����v���,kmmfy�|}?������}�o������{8ߐ[V��u=�ZkU��u�kX�|��I���j�lcA�g��|}?O�����}�o���������	����̚��[h�wwl�j�Dlgk�F6qS��Z����΃Z���h�����GywcX5�������hӝ�Ey���ۺ�c���֌��g5�jm`�Ptj����Q�j�k�}��޻kmiţF/S�h�(���N-y�w��m�ѧvwVv�3�;U���b�67���;v#S�Gh�X�ci۹�wwX�M�F����Ǚ�w��=t���_u��"����G�k�1mA�ֵw�8�>F;[�͈�F.�؍�Z�v'lm��c��7X��g%���AZƌD�۱����(�\`�Z�ѧ]tE��D֠@�����u�����h�X�>\�v�,�vF@Et�ټ�.�y-�X"Y����U�]��D]w��w�#��o7�����v;�q�.��i�7ͣ���ut�S�
�t�[[j�=0j�d�j���|L\����VMI&�f�2�Ҋ�I��!�U��WvV�����*��L�.�1�'�i�<�����$_����m����������������<f�	�Y�y�<��"���`��r��yd�nc5��H؎���k�GU�^n��":Σ\�raE�+TR��;�9�:�y�x��i���=ܚ���VE�Ek@����0����st�d��ƛ�W�a�
����[�PɌ��k�&e�qq�n�7�>����vF����.�nڢ\߮����Y6ć#f:���{�2�����̀!EH�r�0�������˽�Q-b\Op�S�w�ՐUuE�1��D{��\b���k�<W �|.]N�qt���.2�&Fkkj�ޚ"/�::u�˫g'�->�[��`!�,'q��P���-�^����щ0s��*�u�5�n�A��oE��
2�v��6�|M&����X�;!ј9���Z{|�ds�iGҷ^��<������b�5yy���"�v�q��тP}GhO�(�-��r�V�u5uM�Ê��/���d�<ad��� �bLjom�A���Z�dꇳ[�̀sF
������͗Hl�l�[`0��#��aܬ��M���/f��`�-܉�y�.E[��h4ñ����a� q{��T��<<;
�^���n���M�I�(8q��%%��R}�P#��6g5헋���;��&���=[���~],u]Fr����6ǳ��۸ �P��Mov�	�͢��6d@7�O�/I���V�ث��_{����}=��~������o.E�hf<
��x<5账�k�C��Y��~�� D����ۊ�% �����srK"�$�ث��O#A�hV����7V�a�u���>$�
�S�Ng%��p��z'��^�����!1�ݯ�4v��U]�(�9l��.�%��v��C��+$����]�8��Jwy3R�喽�e�� <��[�Se�ô�kX��'&�
]u�.���`RCl����b�MĲ����-s���� e�]\�
T��S���u�36j�<��#ㆬ�Ȭ�Z��7A6 ���6��ȷS�XW���=�))m�<[���5z���\S6�ApW ��G�$�s>��j�ONb�5���N��x"ϰB���T��l�t
�r�k�)�+
���������.��Ngە���8O�#Њ�p�[��.}��T�j�E�n
)n�9��y[�F��/� �9�~�n<���S�Uo7oJJ#u��Y��lY�pԳ���P��c�;��������Ð�}6)�>^��f��5a}�\:�/7/�?˽Ӊ]�i�<�0�^�;U���Ag9�da�"խٻ��Y}��Ͻ�˃Uu�F
����F�\z���Heeyh�5}�#JG'U�����=�/��v��"��D�/%����m��-�{U�i�p]a�J@����(.
6˯+ܻ��N���{R|���7ω}YcN����:S�<�%9��:Z>]vw�pg�홣
��]'>�/�O�<�ߌ�����AE}Xj�Ҿ��"��8��1)`�t��:U@j��H���'D�����gS�.B攱��?l<�,6�\t�����y��'2�gLu�z�bD���;fe��{$V��K��vV�+�:s�N8���9ӷ-�H�=�g�2������5�(hVh)�ߓ�߷��.nm�I�rd��3���^�#Lc�x���x��Fz���g@����%$��Χ�c��e��fNl��y}�AH���x�Z�`sc;�c���f��*���ۘ!4oZ�����F�#�䫂��7����#��,�f��x�[ٽ���F�|`=T�6z�b��r[^� �Pt���xg���vo2Tv�&�0ΰ�"��693���n�Z5���+����=�w�a�_���l�_m�wdI���nd������h(7 Dy!>���cq�U�Se��v�g��G
�u���Mt�n^CC�dbZ+`�Kd֘���L����9�Oe�B���/&O7Ȥ9��K����R�����x'���0;��'����,�藬1��\��%ؿv��ѧK{�Y�Ȟor�-'-��n>��=6@`�m�R��+[@�,ʃ@*܌=Ou����RV:�U��v�BfWQ]U����L�mՁ��Zԏ9޽�~�����37>gw��� ��\����VR�޺3��d���;�ղ���u<�7���V�]�i�.���vz�*�es�*��ߊ�;Ό�T,�v[Q�ݣ},Dc`p3�O�ASz@��޻�Z�0����.wbF��}*�ene���f��]Qئ�M�󜸢�:z#��v�9=��.���F�4�J�[#g����8!��oSL�
K��7Oy�5��!�҃.���.w�a�D��	�Y�0"�9*��U�z�mה/(��x�q�4�@�%��q�>��u�1�Wi�9��n�b�q��'�"���]�.����yf������$� �x��J����e���sw�o�x��t��@(���)�u�n��"$gc��M����9�5�c���m�����E<{a�w��ܗ��� -EoY~�`���O���[Ba�C4���T>z�@�� �#}����Ϯ�N�&�����xT����z�e~�fsA	|[֐Q�/:뎤��Ԥ�����Mu����ɆÚ��Ѳ�:�������[�fk�uN�i��m��3����ͼFM��j�����>u�5ɒw��֭�Ɛ/-M�g��KRV�?FJ�K,Ѻj�6�+����q�3(�X�:��54歟���U;��uRg���Y}y=}����W.�Z=̂��T�@):*u��u3ؚk�U�-��L�]��{s���Ȏ�V���IX/��= �)�����egoOvl�?sLQܞ
pQ\[69.R��y)��7j��h��%��.0�����2�~j�l��Zy��4,��Ek���~��&h�����q�q8+�-����m��,��6�쥒O�^`̈́��ދs"_��<カ*�sϸ��6�M0q�Ά���oi���k�$��E��ml�sE@��	7��Y��j(Jp���O�����;gsf��<_\��m^d+{\��mYX��� �],u]r3�ǎ���vv}&-֒(bkǾ�h����9�d'0:b����븃�qT�m�ۛ��G��\-����a��y!�}3����1�Q!�9y�aKpv�[���Ƅ�C�Y��Cz��8"���)Ne�4�.�lM�LKv�b�)��J�v3L����ň/��=7��m�1A���׸S?�-�?Y����/�z�W�����Z�-��^�û�Yq����vq�T{1�e����6@���Nx����g�K�z�-���y�Y����ج���!��a��^��5z��m�6o��o3���ݐE���X�HD�ܫ�rY��^5!/`|����mNa��|0��j7�h$��:��i�G[6Vxv��o6������΄���HZ27�_��1x�\�Ory �>�wٓ�®7[Eez����ɹ�q����Uơ ��4������+��&6�%�n�W_��eP'r���K ��8�T�*oD����t󤫞`�k�D��jg�':�wL`݈�+�P��NkK����"�j�/���^���3Lٽkkb;8�5�= �]@����6X��C��Dh���a!����휜l�l��w�-IQ3��oR��Wr�	�0���Y4-����
���c�r�Ä�yK<��5*�^��0g��0M:,�}׮�<Â�̕\����M[����36���8u��K�<Ҩ�����Q/(�tr&����������"��Y�۽[̨����4_ �l�R�w7Ct��a�uLDwe�vn��DGl����򫄽�֩�)�u��z������x��k�1�nÜ��F�����U���[�\)
��Q|⚚b4Qu�gyi��[��SN����Y��	aH�����y��SY\���T��ȴ��y����Nd�#�6Ƿ����?b4 ,�ӓ|�[�����+۝7�8]�������ͷ���G��1�g��$q����,Ό��~ �3ްq�Sc-�k�6[��.r =9�^*��ǎ�1�f7�΁��|�&��urm�������X/,�������nM����	�����;�]�~�f�B�=�qW�B� ��;�A=�W���G����C��¼�=�]����:�T�z�l�CծKk�� ڒ)wn��&a����c9�K����1|�����c'�.����;��oz9l��4��fy�>M_�&��R�-�ʍ=tiLU�X<F���py�Ѫ��w���J�,,{|�,Yi�c��Cu\��a{6�{�4r���nR;+F<E���r���ŋ7�n����a�oO2��Q/��� �,A�~���-��H�,T�T�[զ��;�7�{��H�����8�w�Y�:j}��(����	�!��U��d�^���2�F��u�l'�hO�2J��,�����[�2$ZHXlg3mI���Yzk.�#Ew_�c��ΑV9�^㭷S�s�Y�����峧�k�����8lV�U���+���+�뷑���OG0|��b������qd5��.�rO�uq��JM��4���!�;-�F��7MnI龋�H�X�;�����ި��Ps���r�x�3P��X���i}[��WI(��K�`�m�\�xQ�>����ŦrՌ��W�tv�oQÛ�Ou(]>ж�ɷƩ��Y�8E/�4.��[ɫ�����r�g���@u�%e�Wzc&�c݆�`pn��53;��C�5�%�wu�s&��J�����<��iQS3;�S׋���k/~����:��g�Sl�U������*6/�|��ެ\p�.D!�͊$�T��4�w^�`^�\/9�]Z�A}�+��d��U�7�` .��i<z�3F���7�ѵ�ݎMU�,��@�V��C��ź���t�f�}�t۞wk{�OZ;��ydR<�pU<~o�W�Jr�V�����#A<��M2��sg3�l�'5�6�Q��#SzlP�ֲ�j�59�Ӟ�9��9C��TmC�;�|��Oo�
��h�S�9M#u��#�+���3Wx�u���|z���~��)��Z�3�ve.ƛ�SsU��
�Ø&VmN����]���Ounnvd9r\sJX|�J�B�v�ji�[X� _��/-�C+謫�w�D���}��Sl����M���-�2�^��R�U3�*�m�q�����f=nZӎo��*ZHɂ��![|tGJJ�^��'����\�a���T0k���j�(�S�`�� �����*��3g��T��.W��I�0���:�v�I{K�g��l0�A��cNϯzM)�����!.��D�j��u�k��Z�sn�S�]H��3/zs20�q��j�]�Xe�B,8�s�o�����T��f��p��CU�__<v���-�"*�H�1ZNcDwo.{w$͆�R1xL�ה�����tX�4�WIZD�A�+�].T@k���p�U<�o1_#6�t�\0%a�쾐�ܱ��W��+;���؏�%e�r�S�����S6�r�ˠ��}�y�"pܺA�n�G*���`��ji�Ŝ{/HV�e^o,��"fuva��3F�$�;���w��C��)��E�6,��M7M���[�Xm�� ���V5d�8��󫯀�afd�S;��{+W�f 1��L�2��{�Z8z�R,���|�[��%r[}�w�F�ިg<��Ν� 2%�����;�ȷ3�a�`Q�pX�\��G�KT�iB�sJ�(�^'3X�}Ǭbgp�ԙ��dqc��
��۔��@�,���n��Xk��p��6��8�-��{����f�<���WQx�����7u4˹���vd�2��"��&`��s;�H]N6e�BBd6��C��|�C��'��	�vo
�M� cB�ۀ<��p� K0w[�s+m[pռY 4�6�Đ��t��Y���Y{�8���۫�cRq�y���é���_Bz��4i�r�[V=�MmͲ�Y���@A�*ɭ�W����N��k+H"@�5�a�.�F�`�nT�s��S�P�$x�'s��J�z�Z��lY�Yuk�V�vu����;kF
X�翏Q���cg�d���O�����3r������~5�ƨI����sМ�5:<)��z����7F��Mi��ܜ���]��X�]�u|�)�����"Q�Ќ�9<��� �Ζ-���m�q��N[P�]�f9X_�1Z1\P2*��I�n��{�g���X�wԟ=ԈV	�JX�6�V�ä�Q�{�H�ູ.���ε�F���>�\F����Lզ�o[�8|>#�S�f�鼺���v��U$ꄺĂ��`�5�pUɗʗ�X(Z2-�шt�/���u�Z$� ���:Q j��,��g1V�O�9�;��2�zZbs�N9OD���[������%�u`�fɎ,�N`I�X+���c��Eۺ�V����SNP�vmgC��l�)1t��+:,�W�v;4����:Ò�m�*&���y������_P\E;+
,K�T+���M���E���:1G[Zz�6��+m������i�1Z�ys��`�~ͩ�P�����R7�n���o'�tZ�=kp�X�q�2o��N\����x`��r�t�ږIy(͢4Ak{dO���O0�ῥe���	V:�sw�)Mp�)�����J3V-���u�1���z��9�	�M�Tw�+ש�6u1%NV����E����ݨ{�=\�:���Y~��~��~F
��3p$AO*���^��������QU_��wFI#m����{��>��ѣk��$�����o<y�����}�o����o�~߷�G��~5%��'�F���;��v1���5��ݨ�Fc6-m�����v;���M斖�ֶ�����[[ky���(x��ͱ�V������<��llk��)�F�(Ѧ�O>^]Q�Ɗ.�^�!����SF�ݯ�:��kE��U1Gכ�;n�7��3�5mV�6�co;�<�=l�9�hǝݻwdӍ�^F�F����y��I�v�#�ݏ8��lU���b+�]1�z�u�I�1lmY��5�l�ڒ�Ŷ��jj)&.�vq��Q�����;�Ӌ�u�F�Z��j�LMU���mM)U[�v�]6�khֽv�5V�UF�Jth��j�̺lglb�n�u�Z�z��բ�b�m�����b��h��f��}񊂚�m�6ޭ;8���^xd�lz.������5SQ���+`)�km�1��mj��0ľN
��-;Q��ΌT8���E�@��F�
U%}��ќ%{�1�dU�:B]��v&uu��b1�v���7�6lۣC/�v�������
�`&�%�Q!D���D �xJ�:�� ���`X�͵�v����C[�X	�lW>�\���C�:�r0A���w�G���]���\�Qѝ/{�0��BI���y$^ig?�KH�?c:��7m��T����;�胲#ggϻ[�c��(����/u��g}Q���4/ٷ�;�D���T�ˬ�8��v+�*r����w�za{�6||��j����=0FS �Aǟl�p+�ޣ����a�* ��L5vNg�b�����j�k4�+��³^�JE���Fnt]Q9���d�ղ�g����ԥ�ꊷ�'#����ܒ�"�OsS�ݭV���㻶En\wr��X��K����tS��k�
3�_>�@��&�UKZ��r
�ˈOZ$�4GZsiM�(�`폱���W	�z�۝�����`̀�s ͥW1�x��\�@A:��U��(�b!��	�4RޫZ�v��/=5�(���:f'ۯK�J��A�Q�y�`�2w�yˍ:n㭬�t/5��z�]����a�]�w���7S��k%+A����Vb
*�M��Z����'�G$�E7o��U�.٬����no����9��M�o���ŁՙI��pf�����{nmwӒ���F���b��*{��@�P��2����7s3s����W]�؃�W>*�M[8��'5>�T��p���i��^#�Y���&�4��݀�h�����45%M�}u��ߠ�!�@��^�t��N=^T-ަ�yѦ���ټ��sƵ����21��n��-�[�@�;X���l�Xꮌ"���M�.Y��}+������Z<�\��xn�d�v�i�^�)^���ޛ�|�_��^�F8��]�>�2�:U,M�3�;s�dD�@��Vt����B9Q��U-ގ��Ֆ�ƝZ"� �#�ti��S�h� ���0Hϣn+*�z����M��
��6r2V�E��#�{�$d��w��^=؍+N<�Q�#r#��:����#��u��u�T
n� ��s� �Q��J8�wj��xy�[o@���C�˹�ʊib��9�,�&W7����4�n���o��t�T��ݫ,!�\�ܑXc�t�)�iIz������X]9����8.��l��qt�9���̪f��]XmXA�k�]��k�t���u��˼�BRw�]��"�K%-�ځ=���a_�������2r������j@���w���tI�c�!�f������Rs��I�ס�󢕝W�=yf$o"<{^9e��'����tw�rsx�޽�)5�5uB�!b#����Iő@�������:},�\��_3�g��s!KX9�����D��1k�����j�%��v���}��w�]���ʳsu�5�p���,A�~��ѯd���Jڔ7/[�3\�%�O^���4��P8f�A�T�H駏M3�z�	8��mr���`��z=�zHk��.�	X/��<j�{��N�� H�X���[(�/l\�N���s�(����DƮ��JJ��+�
[�͕��Nmŗh	����l][}��1���8lV�WŶ�J��5�r�p~َʈ�m[���+g2�<Q
��J�!v]\[���I�ȥH�>;��S37DGQ������A��A�q&��XV��]?�&]`[nl�����0f����c�He��/n뺲:T�s����+�������(#�4�D��߈����զۀL�f�q3c��w�"E����:�9S��bo@Au�����`�w����ױ�;sWy���\0Y�oTARq2���;�����N�ݑؗ��b��$,�^�F�a�8b��zD蔪gqͧ��ܖ�f��W'�� �9ǺQ�^�hWD��Go�n�p �AA��so
f��Vv��>pn<'68�H��n����q�fI��=ºT$��X�=�םD���ǆ(��ڡ�U����0tqn��`��'e��f�8ۯtN��ڇ�*��:��y.�P/-�4�I!ф�'$1[[�kk�\lDhB4Tx��H���,õ$��(�lոHI��U���,�W��\�*I�����:Z���}�
�z�q��!���E����t՝ܺ7��o�H2��a�.ה����gUR�&�{a�����:pQ�������&�b<3�YZRK+�-��������(��7��� _�Z{�Ep���:k}����s�����J�m��vf���z�e�m.�t����r�S$�1x-C���L�`8����Ws(V�o&����[̶�5�ǼRŨQ�)��j�Y�h�mN�T�Խk���АQ�\�5W�o7�~�K`d�X��}��]��X��$�g�:�uq):9�M�op��X�	~�p�J{���w��6�}o�G�:V"�7�g�T���Q�U5�Y��π���{25/>�Pl�29�pj�v�'���W��<�)l�����F';U�E�מ���	��?�W��R���4/:x�~�ߛ�ow�(��/ԟ'�GU���E��H�V��
�,��5�ox��gf�����7��t��b>]eQyW���A��h+`��8��{O��&�Y�2Փ�soX2�a5��
��]��qD�B�1r2��TS�*/;J�N��o0#A~�8%L��gE~]�|W�\ &w������q�N�/o��U��Y�م"t�cB�XL�}�0ǫ�ް�=Lzd���&��;"�Di����lI�
Gh����:�X2L�Gbҵi���\���q���!n3r���7oq>�{�������j2�{n\.v���0��8�
��e�|��]��0nTtz�C[`�[#�=a�G{{K�QU�ݙ�����{2�ވ��@nR�e����D�mmA��1��'.��'amE�W{O��_��a9�N�������9����(��?NC?�t+��Lӭ*i[l�DY�!��r�exg=\z�k4�J��K�])�鸌��X�wS�b�[&��A˓�wX4�����*��GrC�^kCdjKx��9���.�hΦ��u]��s.��{����V���q-�d��b�o$�\t���&^�'�E���:b�MK�޸{=��4�4�t���B�x@]��nk�Ur�I�ɇyJu����/ws��'� ��s��ȫg�S����p�39�l3�(?495�x�n�{�}|@烵�QH��>�u��a���t�pQы����z�j���uPk�Rvx�R����5礝]^5��7\
��\c+p�a� ҵ�gv�^#�V��ih���T�Z}�k�d,�n�<_z�C�TZ'	��H����D�����xYM�jX�q]����i�;V��.�58б=��L ���*$�	z����R{�v���8q�����5�c���{CHݤ6�#��]+yV;��l�V�R�{ |�y@��sۢ%`�M����t�9�	�f�q���R\wk��Y��C�ھ��ޡ���w7{�v�l��_|3�}�;��ki���y)���"j�7U�����t�O]���^ԮXP�0C6 Cz���6�Ҡ�ǽ@����t���g";;{k�o�JvO�O���3���0��O&��fLz�2㟵���ˎ����\��A1�v���2a���;��6+��=Qܞ����������275����i��_6���ELc���UPl�l��.�OgpJ@ab�<�.�E^v^_D���R"k�,������Y�y���ͺ�|4��
W�����y	]��)�!��ba5��koo�Lߙ��=%[��K=�A&�UL<Q�ɋ��k��rr(E;gZ���z�i�$���c�b�]CSHWV ��a��@�ư�~0�0�鍹� c�^�$�.p�s'��=4��@
�٘���E�_���.�<�96�䊻��a�js�x�6u�DfQHۇ#4�u�w���K���AǏD2���� ���&n�ty�kg+�EW2a׌�]J�p���ͩe���ڹ/�����,�+ovid�)H�e� =΅//7��w-y�xl�糅r��Q�t�������T.ԍ�u�3,|�#U�Ŝ�����
9�)�b���!{�7�%|�9`����>l�ƙ��a1S+��h�7����"��2�oAZae�h���ڥq�tq:~�c��B����l=�d0�.K$?�!t+*���UY\�!�^��Rv���Ξۃ��Y����(g���6��x`�˽�n�..S_�Nn�ʙ9�7����@U����#�L �(��x�F&#ݹ4�E�d��ʳ{�Jr�y˛ӫ3�u+���L6��v����R���S���'Q�R�2��*�-ĉ�����6���^=W� �d~Uj����^s��?D+�V
g9C�^�K*��V"k���u���X��;&0�7i��F�y~a�l}q��y�Q��G7^5�\>o`q��M�m� =N��G�^jx�P���V橥c;:+�/��5nt��Gx���6�X$����NTW���aC��1Jf���j�t�i��Gu��ԉ�M��|ap
˽ܨXt��=��s�`�X[Fq{�������UJhǏc
�	��'��,@@<����zǰ�m;�C������pg�u��@�g~�=��S��� �˚�JR�t����Y;<l���My+=�O0�v�B���eUےw!\�ej=C��wu����޳��J[>��Yy)v4��S�s;-����z17�}�hF�Q�<s5PɈ�,���y�F���.�oH4�N�Ӣ�2�-)��eë�]��#�a����)���R�?���"^M�X�9�:�n�N�}��ȓ,�ȡ�!(�G�x�ޔ�����s�y��o��L��L�����>�W�?c�^����d�h���|M�)+ �)�p��=6w��lG`JyZ*�,�n��b�*B;pY"5n�e�ʽ�S��z��]i�r�l�c��l������y�����
���~섞՛���ߓf��@��\�Y[˟��y�۲������֧T]++ʭퟗF�Hb$�E�,sit`�Kp�nZ�����/\�����B�`��ͮnƮVm����Z�U]'k�Y�L��Ƒg��d���K�xI��3�`ŷ'3�f��&�c��k�&�{gm���Z�ƌ�����z��v���]|�Tza�Fʐ����gx��%{�1��hdS<���gx���T �Ю`��r	0�Du�{<��G��]{J��Bԫ��e��q9�ۧ��t���16�i��;�.=�fj&.�q�')�M�Z/���tsV.��|��[{ Ӕ�сuf��(ٸf�1+*#�w1�����:6�|�y^���_�I͊��jA�
�v�umᾧ�z���hE)5}~�[щ�j=^K��zka*�-�ܵ��=�����u�S�~���`�/��1���Q*z��B������6�GFn��Жl�We�w"-k��0[F�~ݨS�ʋ&��B��$�o��wf���['d�\H�v�Y�����2^G2@���z���ȃ�v�g��е��'��^����̌��4��FUΫu"��@.��Њ�z8x�D&,Dh��b~}�Aʯ4�.�9mIv���c���/����N�I�K+j�ݨ��qv���[K�k��Y�G�f��b�]��[$�Q��n��oc�k�8U�|gOmQ�pc��3gm{�zuc3���3�-aQ�pl0d-�X��\�*�;f]KZ���ok�z����9�Xku�S�V�^���)ojF�B��Z}���Y���N�O)����|*J�O�2�\��슆����qU�ٺn�Z�f��;=f��VW��V(��n�ޒ�۫8%��`T01�=כwVȱ��S�Aj_5;�fch�,'�Li�y�Fs�v���v��x#��u���б�ÒvcEФ���'�R��ш_2x�b�l���c����z^�ޔ]{j$��=��T�n���j�M���]6;U{Q�X#qFխ��y��m���ɽ����1�4)�3�`���WWRUᕥ>&H��S�բY�-gG�*�]�k�Z`��lڒ'�}���*9[�t�h;쳚�t�m�-��H��'�1^o6�E�&�a
Y0A�����V�غ8(r+>G�p�)��+�;J�&�nh���aғ��-�ff��!��d�vK�^��M�u��C�wҖ�R��|�Vm*�ǵ�D���[�o�=�Iw�.ΰE���R��Y�{�Sǋ��ȭ���
+�u�2���)��)�(�o/)�սy�Vu�dp3S'a�x5K�Gau��J0�-sNrޚ�cmP�D �X��T��կ������G��|�a$9�p[��\8��Ǚ�os��p�Y�N�R�\��eNlv����y�)�+���3zG]y{�+����c]�lN��+�Q��m��0-���od�$���+��9�&���W1<d�<4kt.�.��zݡ�}��P�M��I4�1.x��I���{g0r=�r=\8�li.�̻ݠ���\�aeЬN�[p�6�5��Uܶw�o#�om����(t��N�[���%עd�����9���e�$*i�.���T�V�=���{M]�W)��op��,�x��ཋ�#�xW��]��AW�Lk���"]$q8�9���$j�
������CΚ�^lɸ����w.3�o9	��Tyf��Tj��H�L"�x���'���Ps�{Y�1�r�{�u�tK�;ZZ7���Wde������70�����\)fnU��S�̡Y�y4b޾�Z��n<hD�V̒�g���we�J>�;��
�(�b��RLb�)�6�2A�ĩx��wY�9TQmu'[������g
��,ܣ�[Ȗ�vh$J&��(e��=�Et�[�(�m�ݻv�N�|ܻ�v.���¦w�RIz�<{��;عo;�N�>�s5	O"��U�R��ׁۓ���3b��0�*��@�EgeYӹz�����_G�����V"-[TMETQ�����}���'Ƀ��`խ��E�N�v53�|~������o����o�������3�U�w��&cZ~l<ƪ��"$���֨4�,kA���&���wg�����~����~߷�����~~Urk�,bv�0��ض���l�à�-A����$�IE�t|�'mZ��kN7��b����[4X��ɢ5�QZص���b`�m����EM�K�7��%�q���Q��h�gQ��}w\cQkb�֊��]�1���kmz؎ Ŷ��#l��4y��J��h#6�h�
#gN�ڴSPDSkLkQ��݀ڬ�6+i����J�V��[o ��Պm��_Y�g:<��n��k��u\F*��(�pDU�ζ+n�\liz8��m�+X��u����EQk6�mkA���;Uw�����+�3�z�{f���z^�5�E�ч��TYη�`�/�yX-�F�z��Gl:���*�f�"�J���"�[Y6��\wmi�&�T[b�`�v��*�Z��+��hbu���_>}/�F*ݵ5���{��������A���,:g���fV^�d]*c�x�^��;�S���
�u���s�}�|Ω1'��UrEOێ�u>� �$/D�td͖ˋYz�{��m��,��N;�%.e���H'W�.�v�f"v8=�$�z��kwo����="8mk�Z�<��Tr�\���<�^3�Q�n���B{����=:���Zuz=p�_z:�A�^E�W��;�D�Z:���؆~�9�U�*S����l�3c�;�;.0"1>���r��WH�a3U�j����-�[��;IQ��]m	��4g��X!��F@���a����;}�X��v�7�&Ggݯ�O�P �����|�|Â��FFo_K�,E'�ʽ��c8�^Ⱦ��A�Ҡ97d�c��l�6:����ŧv5�r�#�N�t�a�1goa.���em�:@�m3Ǟ���Ƴb.��E�j�.~�Ȥy�%/��׿g�<�7���Ѽ{�.���;�יyp]21lj�>@��Pz���*��.-��O�,����Wp��v��Ul@hk��NdOylJ�������M;�O7:�]GqU�s�@��$�Ғs�t���ɈQ�ݡ��;c�z�JB���{odV/������U6}5v��x\Yz++�q��C-`�dH���F�j�2:��hIkR����_���nn��$.8M��o��,���3��O'~���w�|��<���נ����}�3�fI#�:WkH=P*%��S뛬�&��0=Xf9�e*)����x�tW�(-�fK�[M㹝�pޫi��X���Nz���]Fs�N�x3
Ӳ5�J��4
JC�5A�ԍ�u�ː�,:"n����7��/6�$]A
h������s�U��L��V�\��}����y'�(�S��2�� ��Z@�WŨs6�O�R�-}�zczz�8\������ʭ�d5�;=,͎�� ���p]Pʞ��U�U����Bg�b���wg�ZQM���;&{�4v�;��٫�(�tr!��v�b9Y[٩{��{��O�˶���%�NH�W>������b�nʽ������Ȁ�����*o��N���{={o{�P���sT���ത��1n�6Ɏt���&�*|�mZ�/m�bm^�f����\*!ٯC���a�
�x�v��S���w�v���$��6�<y�g]Ϲ7}�T-��4a����tk���]����SKV���[FP~����o:3m<�w>��)J$Zz�\�,6L��s�:��Ǻ��%t��/��ƳyK�^m���M��������ꩾ�C9+�]����w����݃�쩜�,���鬨P�q��x�����˼�[.�BO�N�c{넮*��["	��+7Olw�E�
�׺ǃ�ㅘ�£^��h����|���:�͌�UYe�F�s�����'�����|��!e�+�m]s^�G�F�,����k}ͪ*)=�(F�g������T�6*�o���SmZ��|�,)nL���=Y��bgӏ�gy-:�>Wd%����SsNd�w������{;ݓ��y�d�n%Kjd(d{+�R���ޤ�����?,��`�H�y�s�����n���v�]�_.�s���T.�R����+�17=��{v6K���c4�=��#&��V���IO8s�Y>�LF�lG�ټG$�-o9ϲ:�V����fx���uq�U�Xt��FE�.��F����`�8��ơM�.ٕ���[
N3zf�>�wA-��;�[�W ��R]�1g<��*e���fBj��f����&����+=����EɈ%��-����f�(ׯ��6 �iT�}!�}P�n��[y�-�$�.$�#5�Ν��i��ܤ�U�y5�m�h�5Áhe�vG�@1Z�Ĉ�Dr&���⅕&�&�+^t��`L�-��Xk﮺��kB!���l��s{��zX�����;+�y��2��K9��wdڎcL#FFN�\ӛ�W5{��C��>�z�i��ceO�_k�y-�Q5%/n�J�i���.�^F��=H��B�9y0)���p+:��*�/��C��n?nf%y�-�2򙅰W)q��:m�}���l��a|Vc��Ŀ-��x�[�3�,�RS=_H\u�\�� z�?*�����q�/$��G>�<�+Mk�����|Fqc��Qח�͐΃�xJm�Ż���y9}ooDA������ϵ��H�'�,�,藁x��Hٗ4:t�'����_'������(����9dE�\�_/��z��be��Н�(���12��Ǭ!S�ObZ�Y|J�;r뺐�U�l��qم��V�͹g!�B��ң2:�3�fs���x�z�^���	c^<�7y)��WrU�A�jm�=����y��N��7�E�h�j�������(�=hl�%�{Sܣ�ZT@�P�S��b���<E�t,₸��]&��@\B��W�1|���/p����7Ouz&�1�W4� ��=�v�B5Zkg���3g���iR���!�y]��H�R)��	�L"�-�u=|��}�Ts֞��p9��~&���8�5䊚}�t�K�X�?@уμ�;kj��M=^�*��Spޔ��u����]G�ϛ1�n�O^����mq/�||A
�g�g�+aMjh�i*+�.V�x,ׁ��u�^�_�1�=e�l�xH�P[�/�d:N�lF��_)��4R1!�m��..������/�l�L�\�;8�k#6�.�댈�S�6���P5��ȗ��t5͉��<zfJ�S�6�>y��A���g�5�\��uH�ࡍ�ia7x}�]��g;��+�z�9�-�t�s�0�P��oN�KS�uw�7!C.|�D�}�:I�]cAr?���ʇ�K��`��J�'V`����>��Z�uh��U����t�Xi��90+�0l�1w���>���&�>�d�i	�u*e�9wOl�'hl�����@�ն������}���w\�6�{'��u:�MC�v��l�Pc�n�W)�6�WFU��v�ف��R���P�m��>�:ݥ�<�tQS슁0%��r�^�n�m۶0��"���y�h=��hJ�����V�r8.���f{;ݗ�}�yu���4X/
-v�D��ꅭ?��QyP�����;�8w�q���C�����L�]>��pXJ�N�Y����,�ۇ����o�r����8A6��+��Ǫ ��3�� �",1ے�MO������Wz} ��T2OH�!g���5UP;�=.C�*��;�D���{j�v�`��>���>� V��).�xF�I���C�xUcC�g���Z�=w;�u��������EنO���9�s�6
=΀I_��eН��Fef�V�L�ӧ��U�����ָ�t�-s��t'|l
bl���s����xv�|E��V���`�{�ʩv��̔�c#�n�y2�I��حf���q���xMi�(
Գ��
��d��s��o�Ծ�mR���5�	�$8 �dRN�9��,X�V"u�O�v�_F�oEզ��j�1��:���h��:�b�M��j�+h�WL����"w�޸Ƚ:���Ӑ��0�jp$��\��]ޫ9�o#y�r����3�y�y�#@����t����>{|������6ؽPQ�n5׷[��zuȎ&ɬ�yX��b�nʷXt���[#5&�۪��M�\+�9���4��H�lޚT��:���W+��C��ؽcV�Z}힩3ٻ��� `M��8%����q�K|Hdk+ݑr7���+]�����ך�]N����?�Q����(�k�X�x��Dn�tMU����/v7#��$�1pQ�V睩��f£QV���ND�Tk<Py��xu�M.�:�:�GD�os�C^_}�2��,Ǟ�y���QQ�-L���[�{�M�o�y��0=ɤ
8�q��`0�=CKV�mSl�*D�TkUTN-�4�g8�|�����x��Z��k����N���]���D��
��}Q��A��֌"9��	4�b��\�BV����f�̉�������һ/�iR�\0�hd�� �*�"!.ӻ�%V�V^���UW�N����tL�Mz2�t��$���2v4�Z��6C���O���6�t��`���:�9��'1�B�<�IR�*�v3�x�T��\�nC�W0�ӂmԊ�t�Y7!�� ��]!p�T.��e����f��wu�B.�ߣs'�Lbi��H��%����6��p��˪�[��of;;Y�o�I<zVV����YK�7r���J6�dL-���0c��ގ��n��
~T�惢�����mH!ڢ6kevC4Z��ۗ�wFH�>�}7�$��Ek铋�3�@./�L�>�qf�Z���=N�vngvS���[��mW@y���8��\.�-�-��;c�.�|S��k�l��Sͼ��FM��&�9��M\U�Fm]��܊49�Eo�!�z|�Q�=�j�
�7�П�!X�g~��t��ai�yY��v����»��e���)��V�B(��ĸ���o����Q�fsNW��a���LSI�Tr�����X��3�rǎY���ʑ�\4���fnA{Y���e��6�{��	U�)m"�O�&j��k���c�Ϋھۘ��P������ه����:�g���;Ir�:Clg3y�s�m���!���W��/��Ӝ����#x����v���
��w1/�M �دA��֝�x�0p�6VҎޯ"+��ׁ�(϶)�}�Ϯ����[��0.j&��'��9�U����W�W]��VBD�7��\S&g�瞏<G�7��n��H����8e1�P�o#�d��F�v��o�ݎ�=�#�D<7B6��q^+����@���tl��A\z�0�d)�h��\B���)���/���I[�M�v��;wQ.O�0*��0��uګLs)���h:{m�Y�ъ���E)J9zt-��YV���S6�#%h�y�=s��/	�=�v��z�ծQ�����T*�j�����n�ie'6�hY�6�>�������ё8����)+��\hk�H'WQ�(y�,8tm�e<�6�~S�'hYIॸ&�=sZ��͕��ci�� 9QKif�ι1��
8-�֩�dC1V��m��7��x�^RX��X�q�k��|���c��u�.����2XRtj<��ܺ�BW+;��_�仏��{d�.�k�.��6 ��[i�V����I�6=l���M/[���嚸|=��.n�Zh9�"�㫬O)�]����kă
eֺ�۵=��?��
�Ǳ����������C�1P�5��(OA�tmN�����y뎝飻�RR��g��x��#z�������q��ݼ�Ùyյ:_�p:��������)e=�f���{���N��#����!˭F����&�.��eP�����l�������.��g��R��7mݎ
g5ٟi{��*�m����kg���F`Ff�|S3�w[��7��޺�#�<3���:M��� ����;�#F(ڕ8x���I����g�<;� ��C�����(�ݣB&���8y�����tBX&�sl",��8�	C��3�����#Ty��g�������ߑ&��`�������" ����q�	B�/���1��
z�G���2�7� �*�(Ȅ2�2�0� C °2 C�0��C �0�2!*�(ʰȄ0�0!��C � C �2�0� C �0 @�2�2�0�� C
� ʰ� C
�0��C"�2�2!�@�2(C"zdp�0�0�0���0��S�(� �� �� � ����0�0�0ʰ�0�0�0Ȱ�0�022,2222�2�2��}��9@_L a� !��� ���#� !� !� !� !� !� !� !� !� !� ;�D � �T �P �A �P �A � � �P �M0��( C" C C*�C  LL �102�2�wC  LL����4Ȩ310 M2+10�4�� �.eR�P!�e �@&&D!�e���&P!�`BP� !�	��eXefe]��0!� C�2�2�2!��������o��
�0 �(���X �߯���~�/���#�������������p?3�n����������h"�+��������g�PE_^�U���x�X~��2���%��?�>��������������?^$�C��S�G����{��@�a�,W�ʨ�,  " P* �Ȩ� t �B � 
 I  L  $(# BȀ�  �  H $�(@ ��*B��$ J2!(J���JJ��K���D�P�A J�(*� D L�� P�2�*�4(>q��,?�����S�j�-("�B�߸~���~߿������~��g���EX32�@}�~��?@�E��L��������~'��TETW�?d?�?����O�U� ��������?p(�+�P��UQ_� 3�z`����������='�=O���x���߽����Ȋ�����>�������?����<��?�x�I�O�����ETW��������ETW���������/�Կ���P��?�W�߀���{�}��H����������I�?�<�����A�����??E��"���0|}x�(̏�}����T���?0�~?��d�Md�a��
r�f�A@��̟\��m�zJA"�T���"�P$�J�U)E��QT"�$J� �*�B�D�(
���@	D%JIJ���H����!#�IQUAQEU(l
Jh���
�P��T�"��TJJ��Q�B�Ru�*��Q�B;2 �����A)U*�T$JB��%"T��	$�D�*��T�*�UUEQBQD*�L��T�!X  �ٶ�>wR��L�C�MIr��:7cu��wCu�j���]�wn�]����ݻ���[Ī�K�tmݮ�M�36�:I���Wv�4���r��(��UR���Q$�  0�!B�
(P��xp�hhP�B���ý� А	4=�\:$H�yf�5:��Z��������8�ݢ�����q˧Z�WS6��vî�]��N�ɵ�m@%@H�E
�J)'�  ���[cG]�nI˺�d��k���Tک\�4���n���v�:��u*���Vj�2���GK��ة�kv��i�.�N��ݶ�3������V E*EQ%�W� ��خK[v�R�Q�
�[����[Z廻Vi�]�JSX��ݝuG0�aҒ���M١.av8KTt�wc��:�� �h�  DJ@HDW� c����7F�B�d���up�s�B��*�;�ֱ�kH�9Z�5N��;4jX�r5R����
�
��J�"�lR�� 6s��B�`uMՆ��S8�uN۷F�D��u�cb�FZ�I����R�5V���]�ح3A�Q�V�����	U%D�� v�x���d4���m֙�b�h4��k�U�TcQ��j  @��� @k�j  �0P��D!�RQP��0��  �  L�5� �  �p P�e���u( F0 �t9�0 �0 �(:Ê�*A)T�!%J�� :�  �0�(7U`�FV ( �,����A��` :�j�  &VCJh� P@�D*R��5B���  c�( ��  %`�ۍ\:��0( :� h L�h 
mK�PX� x)�	��U#@24Ѧ�S�0��� ���چ��  O�����di�M��1T�@  �eU�Fh�)<�@6����Ps�H�UL&���HwO=��R�UW�U�}_}�,��� "+�

����_��"�������~�����������������C^^�O�h��d��K(Mo���NË�s]��KL�����^��ڷ	��-Uú�X{�DR0�ơ$l�jh��DI{xuݴ��ؚ�m��) -X���/Fbh�R��S�]�Y����VSĝ�lVò'kV�J��V �ΐ$�W��60�5�V`C/o~5��hz� �6ʺ�ì�`��x�L#��x
[�R���٬�q1��;�I��V�wBQiZ���Tz�8`x7c��qT�� "���S&K�`\ Z��E�.� �"�և�塎��7Lj�`��R�ڕ���c(��@6%�R��H͸(�4]˘�c���ӷV$If�n��A)�Z�,�S!c9�X�As7s@���m��أ�A�+R�v�b�\�m���>���jK�鵲�el���Al8[F�8A��0H�%A쩮��-W�a�Pk�j�A��J�KÙ�ѩ�t�[$U�[HJ�F:)M�;F�N
�廝�5ģ�&�m*��UM*[�	+*"�5�,����{(\�sV*� ʆ�͌ݡ&#��ɱ(R�[�6���c�u�fd+g�{�j�Csj]c��X���W*e�rj��"�6n��)I�&JFL+~yY���J�H�hY�ޙ.�k�U��0]dM�^�E]�r�^|��9��N|-,8Q�����2�,��U*X�r&`��X�t ӗ����W�Z&�+��Yb�kB(6C�"�jz���]jn7E8#�m�6�ȍJm��f&ˡu�X���w#2j�FKW���j�äkhcyl^�PvtaC�s7c�N�G'��C7�5W�t'
�G��3F��c
OZj���Q�P�#�%c�X,��ܥ@�Dou�v�-otPJ�EtR	�r�S��cr�(��@��Ɲ�/CsR��J��3%��yd�潲�&Z[)P��$�Յ��m�0c꽳N3��aL��n�C6ݧ�m�n$�`4h��0�?�;�|ZL)��N�K�ds� z�RZJ̭��������r��qe\�^�QFnL5���Oj�,����i���2����؃[�쭹I)m,;�)bX��X*�b
�+�t���f$�V�(cq�B=�O"q�YD���n>ݩ��D�����M8�F"U���͙#[
�$졠A"ʕ2)�0���v�!x]h[)h�� �a@i���-]��(�Q�4>+	@�e�o.� �6��/u��v��X)�^n-�n5�[����8�`��8�H�5��Z��&î�Br�%�	-Cf�$Ѩ3�ShYq7��+���	��LJ��2)���;Q\�.�}��F��ZpQeAB�jRq��^��0]����Q��n�2b����OV�
�*HE�=<�*P�Ry��Q���W�P(�I��[P$9� ��
��3d�4\q�`X��qPWJ�P�, Ն�Xb��2��ʶ��l�`�0�kU��k$���ۘ�I�g�*�`R�Z^��ٕw�m�u��CE���j̠�PZ¦����9�e{�րҚ�,b�&Ǣ�������{�=��r����W{t"	���Xk�Q7p�2���fK�:f��gZ�q��'J��*��`��̵N�-0k���]��=@����:&�x�eV!�`"�6[���pj��������������1�LU�FY�i�Rӵy�]䤝,�VJ�t��ʀI ��f�{ObF�Sۼ�ͩA;{������(��Ƭ��x+C�V�M��ac2P��qz�:Vt�% �C�B�Z�����Y�R�P�Cwp��FQ^�y��:�^��f�i��$`�:y)��������J5&�a`]mM�ф �҇DBbe�ۀ�iT���� ���Ie@nMQ��Wd��mL���*�@gWM;�Tܷy6�XY�n��Ӭ#o
PM�p'��e��(��r
��6���h�\*����#f���6f\��m Cb��Ն��72�Qb�������A=1��r���Hn���YB0��J� ���cE�d�H�ief�ңB��ȶ-aKӴ��V62:)�s	/[0^�7S�^���:�b�1,mZ����S�ˌ�^|��ŉ��y%EZ�E�X�6^-�y�X���;�ڿ��f��8sd�+2��\Z�E4W�L�L�I�3Z�ڕ6���T��=��Z@E\�6�ʓP�d�����XQ\ca�ޗ*��N)�޸�����A��:RukY��X�,4�����o	˛��@�ںQ� 7H}�Y�̇+dh٣��\ڔK�F� 4�k4�%٫B�M�/㵬���4h�(1�����Ԣ(���7uj�f劑�Y&�f)s]$�� Vp[He*ݍ� ��ո*�A=����IZ,X�����YH::[{�t�J�e�ʋ �(�rU��쓮t݊��bw�ݱS[h@^*F�� +'��6�pD�^����12�U�.P�AdlC*+@��0B���rY1�l]Qۀ-zd�N֋Y ��gcu���X0)Bsh�b� ������&]���n�:!�sm}����	AK�H�YE�y�=e����jˌR���V��7���7�x�BEX�5`�yY�0����r�M�ډ[T�'v1f]K�/O`Y1,֝w���cӵnV�̙u52�h���FL��ܕ������:��C��R��-_P��s���b�W��5�n�,����I���=L\j'��E�l����mÆ{�-��.��ID�nS�Z�y��B�M���V���l+6h�6�P�6e*�l+��{�����OH��������`�+U�l%t�� 
)DE
r" z��Tz���5)y5F�6��Xenȭ���Y��
ӹ�H�d֝�ת�jp��U�EQ���J�2���)2�&�ǚ�Hԫ�;;z��՘h�6��y�t��
;�C�.��n�Y��T��4 ���+)�K�V4�)MTnYUy` K��Q��KZ[�Q�x���v�l#ySQ���T�]8q�mh6�	��Z�E^���6�U��M��Y����Ğ\9��?<�L6+7C�8�8�Y����Fԩ3kz���m'4f���5h �7��u��� @r�û�؛�!N�d�6[rT��)ӭ��f �0J�XU�F�f�hr���	fem)mn��4�ؼ�c�+m8Cbf�׊�ԫ��ӻʹ�%Ö��R e�(�k<ӹ�d;���0��Z��0:5���"'4^�m�e,�E@��Y���J�IBdӘH�Ö��Z�!vKC�0If��خ��/iAti� �(���Y@��շ��v[e)�j�#FV�R���S��.�ȕԻ�I��>��Q�q��F���#PU�2��Lb���p��haI^������줴�I�x�si:(��aӀn��-D�#qK!\�k&:�1�'!��3'�E�ܱy��cD�,4� hՂ�/+2l�i������sr��y�u�e!��]k�-�Sw��h�hP��V
[����z�&i5v�R]�u��eĩ�¶V7N���,���)Z�~ٷ`e\���OO\��5���B�,X���P���sKPY��*	6oۻ�X�X�L-��!���ۙ��2�r��=Ԡ�n8a߷0�GE�D�	�]Jgoh��E�זk�,*�bV�hyZh�ג]*�
6�\eV�D�!ϰЀ�Rf���޹w3uLZLQ!�ۛZ����Բ��`�
��PG��Wp��(i���U��l^X-8a�yKN"P��v2�y�ݍ�K�RPJW,kwc�CR�mkJ���I(}z�%�TJo"���|Xo��/��ZL1�Y�rց��`�3r��ח���Y�i��)v9���[����:)�B6�c�xqL%\@ESؖf�ѐ�%n�wM�6lH۳V%��@S�+ZZ�Ж�lZ���R�L��EV؂��4̻,껙��ubL����|M�G�Jm�,� M ơ����b�6�۩��t#w,F�Ǣ�1݇��t�S��
��=֐$�&���-&�fW��;o~FB�mҤ�ɿ�F�b�`z-��%��&Á�	��;�n2�3PpnJ��2e�Z��=��F4�:�N�-h��0�����[S%�WW���Pn?��./�m�����X�˭8%b8�a)eF#j�(��V�t��gn�V�Å�E�٢�^��0mV'Ifّ�S*�rX���V7�9[T��fV�S
��Q��Mi�J��~7n;F���!M��a��JE��k�Q�&92XǮ��UKEF$�YnԧF�[5]E"��-�h	��e13���JX��@���!�r��ɴh��_�S[$�r\���HU�H��M�oAf����]m��ea*֬Y���rJC-2�J�qެ��M�ְ��V�ֽ���,iks3(ݬ��7�s-�J��ح�r���u�ۖ;N��h��E	��YZ`��L�_2T`]d�W�n=�H]f�n�jn��z�}t��x���87ʱ{H`r�,9��ݧ����kJ�2�)M�ᆦ�e,��Y/"�J�fϣt���g4m�f��-0:�n�E����K�ױ��(^���Y��^T;�N���hɈ�́-��h�l%AB��H�U6m���*wv�ŭmH�&Z��aM`cF�;:Pb��΁a�ؕ-*�5$���fc:���&m<���yt�9u(݈N��Օ��V%4�$��:���Ck洬��-�s�1+]c��,��3u�6	w3qLϬ� 㘠!���2�=����1�Fު��Ð
�r�#ûy{X*�i�0MҢ)9BB``�҈�뤩9��&�[��t����rœ�F�w(ЧS1*�5U�G�]n��U�C9�ջ��l]�l���L��7W��jU�V�b6�����/m%��2^i0R�lFdJ��M��U=��0��t�B����r�="��Yd����6��Ί041A�� �&�)�H2����.���ņ�G�K��j�),�*Y�P^�G����F�@�]���EK� T�t��5�En�M�N�j��U�EMnڕ�F�8Jf�$�� �jP����Ʒ6�d��J�[fŠ�l�{�-��7���M2�f$�V��F��hK�e�7�0[�^�S�[�+4���[{�⹸ړC�NZ��AiA�BmpJ����jeU��K�+͔A"��,웯s)�N;P]+�� �A�r��w2�թ��YzI�"J�L�Y+`�T�T����JcЀ�Lm�4�v����%�H�Q��Ge)r�e���X�d��peF�m#IxvJx���
��c
�tiQ:+���9jnR�GSQ�w�Jq,�u��>���lT
���r���Y�������g+c"T�B�u�{S��W!�k)��b�,��f�׀b�F���{ 0>W��ve<�Ք�=r�,������[ĳj!MݗJ�����\&��dz�ұ_�l��,C{���)Tgr��;V4d�N��ݢSBl��4���� ���]���Y��4vձ��ň�b�����L�sD/h�j�yZ����;��� 7G#c��6,�`���y����=M���F��i��k �C��~qX4k&�P�v�-	Nbl���ɘ%H1�IA"��7E�����5o,��V˶����l�xiۧ��L,��	�u�r�
Ǚ��hhA�8+L�,�V�����Ӎ@�t�j�}��TĶk�]єq��\��%hƝT�����@J�$�U�:�M��fP����:�F
�eY��WEµT�řC �h��ݘ$ݢ0#%�&Pu�Q5.�C�4���f����Dx"ǈ��Chѕ05���@���4R��j;�JVq��j15��&kDVl J���e8�=jL��[��ԗ(:D���+L� ;Y��ő��a̕�e�������]\U��˛�E��ɰn�e � �+�ڔ�k9p1���R����	�!qR�X{���`�[v��&�NV7�ӥMmd�*R)��wd`��I��9f".�ЧN�Cv���R�[y{nh�ڽ.@ض�`�U��yRl���c;z�����f�C:	��mjX�w(��0���Iܹv�(��& u���S�!Z�[��	%���(�J�@�-�t�l����v�Iw�5閥���`�dr�!��x�*����_B��+X@!X ;��{V��y(kZ5\Q�EIM�,.��ݩb��G2�L�9�Al��[�ǁV$XX��b(m"RQ*��@�]ޝ���0�%�/N�ֱD�g4
ŹG�^���u���f\F�!h���8䰩+�2��kM�������6��U�췗t��̑4e�/��hR0J��2�s"���Y�K��i�ĭ� �������w���dn,O���m@�ABLM�OgΌX�
�cUm��d��N��)Z[S\��tʛ�����'#[�l�t�Cp=�I�T�k"�]�˥%�q6t�yh@�8r���-���`���o/C͢��&��T�:�3/3BB�p��GS��Z:�JV}���X@�bݝ���c&[�j�@�,n���е�Ӗ�r�]9�ur��x�Q5��Q��L��$���+,���ڬ��rn��T�M�߬����6ü4M�[����@D��Z����r�+m��,f*��5aI���$����G]A�R�wn��4>�7�YGc�[r8��GPt��a��+i܇���_��V�8�_Z�ekC���bX�qa�
�ט�Z�=i��0T�{n��Q��'ܬ>p� ��;k'}.�+ʃ5�`ܹ]�1V��V�c�_T�����cWh�z&��T�Ju�u+&��ఐ�+F�<��2T`�z�eb�!v��Cs� ~Q>��*�s ���.�.Vn�/`5�7����m<�o��\��erj�����j��m������i�Sٕ؊�ۣq����{���1�J�z��4��y ��u���m[1�N#Aɥc����g�ij�`{+��i0y�Y|7C��y���;g��.��R	$��:a���̠�	�_Q�^��eq�m�"Vв�ee��U����f�02a���K܅�u�X45��[+QhZ����	�;2P���b�Vਹ����,���뫮���ۧ�C(\�sr@��Y��Ћf�}����m��3��=ʗ�:��k1�;ܧ��$�k�Ye�V�Rnڶ+1\�Sx
osx��o�ԒTgsM+�}ٚP���g]���Hu�ක��Ƴ�N��NO5�+0�'ɗ��l���6#zUʷ&�Zs7$��[R�V%���u��Ը\��m�.j��TW@�����"�\&��@1ue�bƮ���ʺ���WyW)����8p��FZ��:��V�zD���g-@�v>�7�%�DN�9}BД�]�cc��C��ݥ���-� 2����/j�b8�u��e�l@ḥȹ�م�nՅ����+8Wg]L3U[҄�	��o�9�kV�+On&�f�v�_]�N1;�v��V�U7�U������V�i�Nt+��4�7�r&�?t��ǅ,�{A�<nTPd���}��l�^[T��Ӂ�twu=��U�D��u�G[��J�m�7�v���ܡ{*�c��%^K�. R�Ǻ�Hs�B�[��U_Y�_7�c��:پgk��T��9Ȑ��'�ÛKۛ�Գn
s��X�k�tv�F:���*�� ϱ����Ƣ�p>%�˜uuI���.�ٵy&Z��X[�ﹺ�鋓�nZ@շ��h1�|V�vM1gz���z�T�9��[�i
	Nշ�(��8rv�늒t�2�P��&r+WZ�yYNU�m��գ���	}��(�.�)lY��p>�C]f�0	٨(ʝ����v��Jֽ�Uʮ��|��*��4�Y�1+���`��9u�}�)�
KW-�o�ٴF;��d���P.W}���lڳ׼3�
���!����v,��o�ZP�+�jMMN��ܮ����!��ՙN1����ur��c;�:��7Y?r��83E��w͞�T�հO5r���ǭ���m���7S��->�XL�1�liV�|=ھ�n`�j���g�}�x�{p�Z ��^�7H�;����H��<\E:+���/T�krwgL+��X"@��vaK{M�����A��X�X�`a�p�
�a��f�/��Ѽ�Z������=յ���P�[��ͳ\Wou�v�i/xj[8Y(X�ř�u�h�}�v𤳹u�v�u��[���6X�|X���t�We�����s��(e�5����J�����[�51̔X�r]�bB���u���;;�tfjN%[�ڸ^U����@�
�&hvS+�b7�VK�t`�z.k&'�)��=xPT��l�� �\M�Y%����$�/���;�x�YY���̮��WV����Za���#gj������F����;ɜ�s���)�Ԫq��n�:uvI��gj�|��NZ7S������r�3E��Xmch�i�yγ3�9X5 s�*x߄X��ʋRgg���̒���M�<��<��1EӸtL���H�u�ϒ��ek��ٕ�,-v��1KTQ�����Q��W�_;�����mj�,#����9���8�E8��Ք.�(� MupD��^�8�ׅʺ17Z�[�nu�Yu�w����Z-�����s�{�"���u�O��a*�x�T��ͷN6�-͎���� {F�\�Js�f�j���27BN�C�
�NR�̀�gUk��K�|�������Ҧ�R��d�+�e�p�6C���Q���˂�V��H��ˤٰ=N���ՠ���m&x,�5�|�p����n\e��*s���<T���x3t+���F��o2��>	��ё���k.�عk��fX��Po��;:�n���2�(T�0m�i+�(Dj�Wo�S��Zʹdr=��`r��.��v�X�EJ�8FK�Y �Ѹ�;K�h��.�.3m�;kw9�]���R�vt`���S+4m&���jD��������.JL�}��n���.� <(�]��Yp�����K�P�T�7%ÛH�%�&:�bC���r�!bH�3\��u�MmN}���������q�[����UvI4fg1Z��Qhϭ�oE���J��:�Tu�*�*ᒲٓ��g ��Wp�����e]I]#$>��W;Z5%L����lq�V[}NR��'�է5��#��Nt��<]j�(���=K.�:��q�(�i�P��^�.S�u#�V
��fu@Wfs���R�8�E�[4:d�7���]�.Ōu�:��5�@���hcS+�����72�o����cj^�/��*�h�ق
��O�Fgm�R�{P�6�"�����8���ҨVc^&�Φ)��wwV�RiJ�ܽoP�8��w�}���Q`"���u�K%!��X�OE���
;Cl=��9uݎ�x�X��5xƤ+x�W��P�N-9��,'�u�7���o���N�ۧ���~z�2fg/�S]�C:��;�2������yW[.� ��HX�j�6!z�K�S�+JK����/B),�(�īZ��]f��X�,f��]T.f�0�l`ݺ6i9]�m���QN�3�
�b�ֲEX����o��d��ƺ���E8l��B�&���固M#o7t�n��\k�h�\�H�d��Qj����نS�_,�{Օ�[�U�ϴ;;O@ZdEV�*ܕy+�Xg�t۳/-���b�ʌ��[˭ls�C��b�;/�C��%���4e�f�ɭ���i��W�i���ό��/V �v]J]�+�����Iã���۩�s�x뤭�:�wAr�.�*���#�-�q��U��Y+f�7��� v:E����0�,Ԓ H1ū��V�U�y�{�aOU�6��w�w#���c��22j���,�4�#n����"�Z����g(��]�̕�t.8J�=Iv�=�<��Y ���uB��E-Z�7�ڷ����uc�`5���bYE�`�l� K�N��+��;Oxᤤ7y�	#��OvWVs�g�yZ� 6�$*�����R�*�D�?v`+g&>���7`c���=X�Y�����|_W<V�y�����н���);V�L��>�LN��]u�G�b�)�*l�{��΅�+nʅADP�N�.�k�L��s���tu��t�N5�N�pc:�,��_U�<5�O�S���Ƿ�&�n�f��I?E�����R�q

u��£��&�e�zy��S�K��5��O(�:�\0���m�r��nՔ����s��F�z���gFzh�֌W���*]NVuD�[�BQ�,�Op����}�c�{��F3��ŉ.:�)��:-���%0�wr�f�J�������F�&iܧ��w�̷��7�]*C�N7�{CW�6uv"`�i�_	%�J�Y���U���i����C�C*��x��8-@�V�M�8`�XE]�D���9����J�;��R[fh��ӗ����x�Ǐ �a�Dn��6�X�X��j[9�����UaL9���;U�ʛSt�QK����O��"*Ѩ6�̪oY�ԝuȯ4GXVm��������W�[#��]O��֗�s.ڗo�����DK�y��&�J����պ��Ùy]`y��V��X�*��POa.��ǭ�����O�J�������ݿ�4"�k�+���)Ce����F���V��b�P�+�=�9y��ؖ�c�ꅬ���ZpR��i�BV��aX���}���1sW�|;NXO$b��(�m!�m�̹%w-lPR86�%8-�ۘ�ޤ���HhP������!D�����о�CZ�ݣj��X�=ܮ.�n>��ϭ�����Ƹ1��9������E"w�t��39��2��EZel���E����K�b6]���hA��Ѯ�z]�����gZ)w��7�k;��mNF�����7�V3d��l�X�ʳX�/P����u�"_lɛ!yw��� -����`����"+�܊����\M���:��Ø��_Vs�����J�YA��[�N��=6��d�ҵ��X�څ����V�����[��X�Xs雳�f��2��i���<`���γo1���N)�
�}`ԭ�:L�IqW��z�hLHY���H���*����A����"�R[Qc61��U� ǌ�G���*[ݻAZ��ڱ��Sm�ʁ��l�����;b�9���4��(���ʑ�3�9���I1dd9n�T{_5���3�l�da��s��:̽�����/�'�Iaأ��d�8Q�U���*�[��؂�
��k�Ӿ줮�=YOS��u*�ܔ>�J���.ʶ�)�(�oK�o^t<�,S��<<� �9JN|k9g%Aގ�ø	��V��tv;�P	n���`�y�Cfu�Vc�fɇ$���w[��d�w#S�����s.��@��^�M�[C�5wơ�ξ9�[���U���ɞC/�H��w����i�H�����g+�@�Y������}�几��}���PO��ّ+7v���w=�9p�1,��(<��Y��j����\O`����};*��͞�&�f��]q�)�=i��XTxÝ0*|��ZR�]�IVf�c�jO�o,E�Z��P�����/�Tgѡ*���f���w�ڭ���uټR�|ѫ�]PU�w� �Hv¹D�Xٽ��JZp�b�6��V+��w��uk��I��D[-�|��U������X���Wn9g(b��_GL�d.�k=���F��.�x&T��'*W6/p[t��q��[��U����:E�����F��i�b��+Z�Ϧ�խGl��A�}�e�94��h��
Cە.�0b�ee����'mo*�2e��*!YjƖ�c�lL���q������l��J���c�¸:���CԱ������v�pt�v=�ɯ)�XX6A�n<���iH?�����u�t�5#s,Yua!�(�f'<������ it)pp���*��Q�x{����c��p>�ɓ��Y�!ceٱ>H�1�̢�M���ҜӒq�HnR�/ SFۑ�5u�Ɵ.qu<�+8�豆v!wF<YW�Wb�{/�wl�6Z��j��6�t@�z��;$2[rv�$hز�����*S�/�n��dV�p�!�.Y5v-���Y@ȡӕt��\7�p�4$�V5h�b��	���]f�ءR	�U��C>�ϗhQ�f.ǒ�}�6f�%ul�sp�)���u��*�41����9�7V��>���v4�@]���rOL4;�\ݾ��-'�pj��kkG�+ǽ.�yY
��-�7}\�M�z-S�r�&*�к.����{l7HV�)�[�ȷ�R�v��C�#qd�n��|��<]Kٺ�#�9"[}��{^���iCn���BKwa�O]\�GN]&]9\D��k(Q���;iV��T���2D�r�#�.�V5S��n��ǧFg$=�*'#�c�U�;�n���l\a;(�U˥v��諦�[@8�s�\9�6`����^��[�mgݲ�n��ٝ�i}��5
��0��js��A��p�-�{�3!l<��V���t��%��:�єK��H��=�����	y����� H'F�n��a!͆T)%ԯ{�W�Bӑ�u���ޫ����6#��Y�,5��1ڶ.��o\4��y9��`�Ga��0�.�>խ��,��Ӂ�;ҍ,/��|;.rz�!���ه����3��o�9_4�ѶgT���mh����5+�/������������sz�1�S2���e_m�Њ9���О�;iR�u��i�����8܏�~��������quP2-�T�aZ	�O0��T��#o��q˳z�v*~�_�K'�U���� p���*��ɤ�VL;#u�z��i٥9��}���G�2�X*E�mo/����He���Sv��ۍ�r1<�݅U����Δ,|��Εy��X��Z��$�X�<3,�����l��GĂ�(�����[��]P`�z�Ikh�r;�C�W`�"� �Ut�����z�*���N)DB��Z�]br�4�YZK;����ڲ��6s�\�5�͘��awDT���U)Q�;d��fc�-��F���N��[�0Dj�ݔC�L�63F:�%*�\�|���j�bd\�6�dL�c!�������NQ���=�h��Ӭ��E]�h�%��$�n���U�&��O.y�����@AZ0��u��fe���2q�@�e���Ҕ���]��%3�L6�<�r�8��ɹ[|T+��؏QA�[ʧj��ϖdQ:��zӭ���;����`
��0�w�}�Z��+\p
����Xܮ�0!x2bi�u���e�kD�6��|�0.�4FR��C��3��:/S;��q�5:8P�j�U��,����u�V�K̜�)i@0ꝉfH6[�Y�]^_P^#��#F����ܶv�I�]Ξ��t�I��.�;/��Z$jq���	��41;#���N+�:��d�fv��l�ث%Y3d��#�K}���)9��i��֙m69jn�*�wϓ/t9�t1f��S3��wuY�ӌ�����w��� ��� "+�{����w׹0Ѵ�~;���]t�;��U��jQ?[K+{� �gZ�gMZ�H�A�����vGTw9��ú�����4��gF�ŭ�5Vݗ��U �)��B�g߇a�t�v�³���0r�ZlS��UO��:8�;}O���;�+[yΊ�{�\J�}+���Z�b�6�e�fK��om�@%+��H���V̧`��&���U��k�>��K�qT(�9�{[��U�c��Ê��a���T=d58����Gwl�aw2�&�t,f�Vw&��	<�����jS�:�ٲ��c]ի��]��Pv�p�*�Eҳ�ژ�f����dM7Ҭ&��[ڹ2f�ؤܚ���`=��L�Қٕ�R��˱՛�y�ES��
D������y�ok����Em�Z�m�M�V�U�_�D�Yi�hG����&�ȚN��~��"���$k��6��Є�hX傻���*a*�Yz�rň��&Rcc���-�G6g6��Xb�Т1��sJ�N�v�I.Ĭ_8.���[n�p�NN���� m xH�nr�}6k�S��m����L��
��6n�gJ�}���4���ZU���U�Z�sT�����h+̾K�:L�pB����}Pm�ɬc��}�QW��t��70�ף:M�V�	��0�sq��R=���v+�4�����qS|C�rѨ�G_%�]�*'����Ф�]p�땀��\��.���룕.��6 �
��7�"��e���Lw�ʂ�{w���/���+B;&
J���-�F�΅�|�I}OK׽k�y.�X�U�dӭ���m�e*T3>V;3���Ū�u�,h�|�ӷSF(�U�����c8���ya1fmH*�f2N>��u�Fƽ}�������ݪ�,��Ժ���Ơ�yÞ$yī)rT�S��7c�f�x��Y-@i��o/�Af�26��fN�cN^�땢�'SuO&���Y���ۖ�#����16��1�I�w@�5j���]��}��J�v�#GXL�!r]��C�+T�cL=���J�N��Ħ���ОR���e�xl�qӏE+ь�L�u�����>-)r9@�;a��<^V1�k^-��͔ݞޢM�We%3qs��i���S��C/L������ޢH�[��}»d-�.�壬���D�"���/�Y\���9��� 
���S�8n��-��6��~��_\�+��N�ԥQ���/u#hk�sA�Ws�%�wi�������*m ��|�'���y�����yV�f�ې; �ٷ��ʚ���C=\��2���m��pP��3��S�L���YewY�,�8+e=6���wӘ�<��0Bo	�k1�KVqh��)�w�+p�w��;�p�:�`c���I�#D0�b�S�Y�m��͸���LAy��ժU���z����� (U��o����|����a�'@�$��or���V�wl���R�=ݺ���ӥb�����ψ�lTy�ܶ��2S[V�Jt�?Mz�������r�<��4�s�T])�b9j��f��`�E��]Z�N��R��GKf�AG�Eͫ�;f���R��	瘭h��E�z�����yf�8�>vT��հ�n����������rV��.빩��l���T��lq�O�,+�wR�0Ao5ot�+-i[[T�ZR�z��+�r����d����&����}�[��^��Y�'V���ū*�IS����zq)H���ްڽ���[`�>�f9��Q.����F����˴VX�W�콽�PK�N���%y�!j5��Q��,�I s���+tZ����Ճ�n��:��P.@��':�X���bim��M��`��{7#�T�-+�-%��7������`��^X��'|���E����7J����$�&�*��+��;���5k����+��&T��W� ��a�'f!x�Z��5U�<����N�!*���ugH4Z��f&���V��Wz,���%�56��Y���)��ի�N��J�A�J�[O4
�+_[N�ث��� %%������b�&�囲vY��ʆ����f#7z��=DZW�x ��Tv�@����r̔r�={�s+㪍�|�K��2��l=���ǚx���|���e�cn]�歙�{�ܻxZ��}r������}$��8��e��V)gtj��oF����|���h�2ѥ,h�65WXu��Y]}���6��_|
|E�F�����.w�hHJ��� V1�ٯ����ǉ\����v�+wR7���b���[�����VXr����7�;JK�6tl���33��}�.�j���hBl�4��]W�n�l8���֦,�r��C{�:Ԩ[K#�lG�U�wïm�aP-�4;t���s�s�Y���1�����<���,��rB�1z������'��f#��2�
R]�1B;5��m�G�Mk���oc2�D�B�:.��9+�-��ѥ�F�w 8���y���o�Y���t㢙]KF��U��r��L3O:&3���0*Fu��EHR�H����9JU����!�]��|H���B��)na[S�iLخ��U�V��j�J|�n�Jե:�ct��Er˾I4w%�q��^K+jwLֶ�=���嗟aH�՗A��lohMqr]^V�#�q����U�v��U�Xik���'m[�������4,����\�n�BJ	�����oWٯT�Tcὄ[�SZI�{uϷ9�&Py�E|��2��jp�6n�ݷ2�����}2&D!JVzr�pT[�]�P8�U�^Cy|�,�|T��#3$����n�Go�2A�n@���w*��Z��;��4�m@��LC-�`�kiIK���r��6��X�ru��Oe�۵}��ہ��ڝ���A�4��na��j�-�hZ��x�H}�V�qh�D�nG�������PW��v���F�Zc�2(Bd����2��ly����fJJ�R\�4l�a��ef�XxuŎ�졥0�L��ݸ��r��1����BMР��5ҵ�-4R[3��9
QB�d�(��Aikw7M�fU��/�k�2r��j��;�Ȣ���DB]��;�V�	���:�9tk�[�:�jq��;����β��	y����z�
�S���f�AU�h�vl�X��H�����*7�6��ӻ�v�W�"��p�I��Μ����bp�-ՓDJ�N2V��ɻ �u�"�;C{�u^SȨb��H�̽�P(_&b�kY�]wt�n�I��]N�ٴ��yY�|�y]PDkZO�n��W����t,e3�������t*-Z��)^|�n�J�Yڅ�U�T�$�j�٤�9��Q��@J�f��g�����_c\��PkE���+ċzk#5�Q�Y������h�vd�x�:�v�g�X Vb�X�8�ܹnՎ��7�;;I�p��]*S�U�UIO"R���tb5�`���f��B����E#��rf.Cqm���mfTՃkT��gH��վ8��}f1YF�o�XB�fU���˚D��ԣm>�Ro`�����ђ�b6�d$�����+iR�2�c�)7v�h堤X�L�t�)��{1���	�X:��wX&��wKFu(Gj����zx4E�C���$��c`Ɲx���wy�)��x�+8E����;G$t�������-��Y�
�u-0�gU�`J޳��5n�6�>�����R���&+ek�Q��A�8�*�	YM<��J��:�=���N�:�xM�g�K��e���լt�*�2ʻW�C��T��Ic��P�k\�ɒ���]�Φ��{hP`A��_r�a����	���9[�uҬ���헅p�o�Xtqq|�;ʰS��V����x.�Xo��s9���JZ�ӂe_@��@nbҟ�G�]�
��������H� ��\2��3pc�G,@��Sb���XG��ծ�n���l���z:�άrݶ�{R��wm��q �u����W|1,t�ܱ�.Sr��h��;�M�����ˈ^2-�;���j	|����W��K8�a]\�$���Ag+����I�w��;q�v��ֆhy0E$�[!�����0�b7	�Z3�Na�}ĭ�f�Զ֣ǩl��Y�]1{@1�5ʻ/�ϷCW�4)�㛝z"�r���V-7��n}�Y�����
����0��ډ�|Lv��}�����|Ja�jΝ��"o�a"Su!tx +9�8˴�[K3M�'���}&t���+�@��k5�`	�lQG*dtu�F\;ۼ��B��Ӡa�ܫV�{�����ܫ{Z�91u�0,@�C0�O��؟M�B�x�&��P�(�e�V�ٌ.�}�5야sv񆩮�����̿�C����W�Z;bt��ڷ�;Ld�F�*�iDŁ�e����DF/���-ű/e�l���ad�Y$����ڰD<a;�zd���D�m�\�c�ف�d/z�r�s���cg� G|�<�e��܅ͬ�G��]w��f �7/�Щp૵�� ���g+��ɣ%�l:4�:����6&��b��tȦC��ëcr�\�e�ذ�X�2�H��Yy]d(3�UҳSi�F�.�t��:6�YI�.�I��K�V��J����qHֵY��#!T6�J���9){Q���]�CZ7$��rh�ohs�6����co��[\i��*ú�dۥ]X�<�uƘײ�sf.���Z��[�va�BP?Kӊ�}�|յ:�V�=%b� f>!�z��_]�v@z���k,PV��
�݆�Ŗ�C����Y�Y�ykk�-������*��;���j��8�uƟn}��a�w�V�.2�R�)T��tV�3k.�|9p�)�م�Я�u�=�պ�FA�W8�[�0l��i�D�(RЂ}�>�,X��u�@�2���-�8
�]� W���=t���٢�/df<�
�:3Ɗ�)�_i��Ӂ�S��E�6x��G�L��/-ƴM������h����4�m����M#5���;z�g
�K�Vw�bך�K�
�᯸&�k�(B�p��]檋C�y�F���*]��B���؞G6����8S�Hۙ�Y�F�Y������>U�q,��ʖ��/r�y�5�hʹT`n�d�@Na�{KK�4C�����K3�_W;)�A�#��h���i�6/?�͢&5�ST��b�L�fK��v�*E�wx�����x�������׍�A�l
�_0%e�"Cgur�o�;�#�!|ӻ\1�g	l�P�N�i�(f�����G���;2�eg�VS{�y�L#����dO;�@]��2[D�p�ׯ9 bDO���-�+7'�E�P1*��ڛ��̾3]����GTk����(]��օ�)w�6�e`��B]5���L҇L��Ƶ��Լ�˥7�_^ŤX�Ԗ`�:�ݭ� �t_`ٴؕ����Z��ދV�E�ε�U�����R�Ԡ8zn���ޱ�iF����I�a�VXmgcCT��c�؝w�c��|ڱ�^!�̇���޹�H�Z�vg��l�F>�}Ү� �P��r�<�;���V�z�f�j��N���u!Ʋ����f/��m.�p>���wV�<z�E!u��ap�z��r(1���� ����O^��W6vECq��Mv:�Prj���҄��-���V=��C� WǙ�xZ٥��/��{�.� ŀ�ꋹ�̼B�P�J�Y��;ѻ��k��iLv�R�ڼ*f���|��ü:��y�/�)j� 9��)>��4Uե[D�wQX�Y������}��3c&0�8J] �u���s��4�����Ee������B��L��c�`]�"u�����WmN��K2-w�#�� ��k�AC]H�I��[U��q��yr�������سCAY�3�j'h9cquݶ����K���a�{"���-$�#~�����Ӵ����i7e-�T��3;:�xm��wx��⠑����kF�]w��_f#Qb)eCAaw3:�I�P�N1���G����ϸ�9`ES��ve��#�y*����B�K�ľ:�hW�ܫk"��ڂ��8ԻPܹap%���2L.��i��;�12�9:�}l�[������t��/�<�dVK��e�7RN���z�Ó�e@yC��PEK���	7�k+
b�uf�h7B�X0#b�4����n��D]��U�޴JV���t]E�$u*����逜��ƃU���U:˥�A�+o6�̽�ȷm��qc:��4L��|);����t3}}f�JWS jwu��*�xUf�J	%cMeHؖG�l;y�j�W�7z&���M+7�/ˡ�)Vg����*�s��sT|Ү���=v�8g]u�
N�v>��v���t��Vd��K9�+u��Ս��1nC�^tӝ��bQd�,S+Oe�*׆���WPY{�"r�#e���T���n\��t��®����JY=�E���c��46 �+{�²��j���scg��ם5�o�]�0`�������|��m���Ԉ:DS���H̩�Gnr�8��VL�Ǒ]ڊ���4ol��,�C'j����]�XK�w�q�8�k�}�+���%�����T�=�t����ٽ�8NB�C*�wS��� �e��mħ���nT醞V�'��!�6P��Ι���#'���aY��5��'k�h��Y"a[�iS���C�N��ɮ��Y���&^D�r۪��V�&���\�՟f�kM�m�B@���45\�p
�PT�%����YC�`� �ަ��n�����X�kjA��W-)l�&��?����X����"�뿿����]k�jfl.��sݹ��8���������BwƯf��q��x��ŉke��D�L�˓�3�L㪺,܇���ܑ��m� +�� Y����6��+k	�����S㍌�tgs���t�Ո�{c!!4��Ej���Ü͹Q�b��S��L.�o-�����k8�c3�U�[�������^�>�K�����v�Ś�Jp;h�ʔ�*_\�U�B��n�ʔfhfL�����<�-%���'1�"G>�1�M�]��`��%�3���AĀ���?-�46�R�"GRC#JJ�v�9���������J�NQ����l�A��z�$U�|ō#)���Y��^��iL���3T�om>�:J�]qf%@� `r�@n:ņ{&wr;�l�9p�G�/>�oT�)���X��|���H�9h6c��}N�V<�r�MN�GI�h�1u�noa�i�]�L��z��I����Z��״0�9t�N��_]�ٷ��ƀ3�A��G��z(�tgXTq�m۫F����tNm �����:�����k�h"q�aô��
�����5����*^��'�.�Fҳ�M��Z��f1)��7V�ө��﯇)��Iѩ���+9�@導rz��GO(_i�C�%�����L]ck�Ư]m�������S;n���}y�YK��צ�cK�x'Y�Q���{Jp�$f�4@5��mlh((�D�T��lb� ��j"����lM415T��EQ3F�2A[d��c4@U��hrDE��"��'l�5mX���Z-���cTTAUTP֜SQULT��cF�����Ѧ�mKCLC0[h��5LT����Zq4UPU&�j��T[��)��F�J���CMTӱ��t��H��k�Tr1DT�S��Ta��"jAE;d���Vê�vӱ���))��(�mj5AT�4ִ���&����5��k[A�Q��(&b���� (j*MVmb
"�h-�QCZ̕�[bb��J�*�)��Ѫ���Fڢ(�
KmRD�QZ]TICMEm�(
l�����־|�ހ�<͹O�恻ivYСm�r�;��Y���J�Jʆ����{jT%����2��I(����oXf��f�����-���eP�+�R:�[�od�����@�dk���g�k'����Uq��o�+Oԋ"/�}�hXo�o��Y΃�p�yHẞ�^����Xp����D�$t�mߙ�-�
�z�Z}�\�ׅhF/�_<앫-�x�Ա�p_�b��/���B:k߮
�)άV�O�hG�Xu0��<M[5��Z��߽&�pS�߻wݹ'���+�i�_�'|;�Ug���J߳�ƨ�ه���m��u2�<*�*��?fĭnux*w�pW�9�^d�� xp���F���U��]}�m/V���ʬ�H0�;�3b��.g
���
�D�uG�iy9��t5��S�~�5��Ik�ܔڥ�F�ۦoZ(>�u�o/G9ޭ�hd�	8Z;��W?�""9�1F��$�ҙ8��M��-��������)�;���*~x�l�$�K�C���.?:ƨ�,��aU�~u[RR����/D[&���]�j�u�e�3E��R������(_w;��<Eާ�'�V��(����M�V �o�;I��J��iV�Ln|�w�SC㷶�ءǀ��S��h�A�!��m�Zs��C;q�хǟ0��̘^�nd}�*s�n�F�\�{�ǝ����j�v� ���6��$���]���.H��w"�:�+�5�t����앙�}ꮍ�~_-���b|�O6T5��ە�����Yg5\��tĥ�=�WؤV����S�!2k	��u�3��*ّ�	�Z�s'ӧ��r�_I�gx�3���e�(�ª�n�Ă�����>G~�u7:1�<*W�����L!VX��eҼ��M�~��`���ƢI=��G@�ԇ�[�I�;k�n9�\�r.����[��Ӡ‫�/�1`/��֩�|�����Q�v����r�����7�lgnDѮ�z��s�k̸M��ʥ7ꙕ�V<I��u3k�1��[g�W��=J��(/e�B�ͩq�����U8��{|�=�F�K8&�}�=�>�7��T�W�4%�|����=n��8 i��!�t7��|�3��R�ϪW�-��DxN���*͘V��%��3�w�)���4����n�z5[��O��s���3��*|ꥪcQ��|���{"�g��G��^��8В����Uzˣ��0ՀOx��\ ���M~u���8"F��<F|�X��WF�Q�o��]tsx�&�f�o�/�js��P��=�t���]m��X�]���G�i!�6�U�q���Й�N���0�9,c#s��<��O��*��a���"(�K�i,�|����W�����ZK���=Aނ�ӧ���<��.���j��3%V�]�9����L�V#(��N�����Rߔ���{kI�5����y�|}���5תb���x �%T�*��1X�{��b���w��]v��\~�[2Q�L�>��/D�����iu�E-� �+���{�+�xf}enߴd���SK��l�_���L����Wx���.�[�=X��,G G�IՓ�[>��s0U��O��t	�D�yWi�#����B��,Ov?q��!eBL�]�L�OoL������4!�Q���D1Xy�����ʰ.�5��o�K5ط�9�b�v07���v����kN�&�*��J�Iv���P#y�E>3����o���/�=ޘ��ie�Ι��|��y�):���֏j����N��6,^dڨ�+�Kf�y)��v\�iAp1���S�	UBb��TͲi�Ov
�]7
I��z�������ZF�ʺ�����$�ԅU���8}%���Υ<^��O��wF,��~7c:�I����2�)�ӫZ�6ۏQEAf�e�6�W���S��Pή��g�uo���)���*Iq�qzft��9�d_J�
�EE2{�=@���Į!�:Ni�;_Cabu�n�9`���Yj�����l��'���Ν���3�ׅ�zsHu���t���A�U.�9r��)`������	C �y�M�P���b��c��{��z���[Li�2��d��]C��<��v=�����{�Ӿ��V2���>&����2��:�N߸��X����6�o�[���xVj~4�{��ʗ��]HGq�먜���h�s^�������u�7'�8e;�Ɵ���l\�f�^�ǀ�.����'�et+��������ٲxJ'�s�I܉�GZ��*�8�^��T�]�X�|ˣ��+FZ���=̏}�h��BPH�q���^y/I�k��L�RYu]�ز�{]yQ����Uk�
g���Qh7F��3�B���k=�z��i�=�t��g���鸁TP���ށ�k�����i{n���*]ы��ij;)=��e�>ZN���V�gD���TD<m����}X��e����$|}�(U9踜���S#u�R��]����	� Ո�Ʃ��9�Lv��I�0�
���i������?��{��#����@���W�-�{*��
y���?Yr�K/{tb�s�����3)����aB�\�a��N���=��`]Y����t���H�t,;�ԱP=G����&TY��p�Rۉ��H�J��Պ��R�U�E�Awrw��\ ����)q�.�v}6z�}#�\�HJ��ä��T;���O]>]�!�z�wm���Z��*ZOHF��c:�6����	�z�Ig�Y��>$��x�e��\w��k�${�rrbt��(u�N��ݴ���YD�Oo���>t�(n|N~b�`���t�8��eB�W��=N�-x�u=���W�E���BfԹU�0��`֭7���a��#߲�O`œ�F�i����7BW����4�zV���Y��2�\#VbnT�h�*�Ku\^�y[S��S<���_��ﵰi��=�p�u]��k:�y#�ff�C]�&��t?y�@TTQB2�˱qVL�B��Zϸ���<��Y+k��.�$� �܇V<�|]��y83�jf����p2=Gǩ�=�:��,{�j��S+XaD����kO����{��+D�~k���i�'j�\��ae;����i�j_����Υ�.���U�t(U�DT<8	�}נ�����*�G}
��ƫ���{+0y�~�a�_����{t��R�`����Ӣߑ�{In��/�Ax�5����\�ç)�3����VfV�W	������N����7����賴�+�����h�s�e�bV��^L�R�Q�v2� m*�`��Y���.o�yowL�о]�(�E�'��Y8#�
��/�S{�,ʔ=[%��Z��-�Vqr�����
�}�7�F_ˮ}��p�o>4":8�(��[���3�p��v�q8�ū~6�v�}�9 �z���<#���\^�+ą[D�b��X��?�l���<�[ro���މb�e�U��=ߣ�Gx�+������l/����l�K<ԮG�ݏl����֜�+5_�{2C�zg��^�	���+|��Z��ߛ��Dx��3}�{0�G��ｩ����uN��5Tڿ*.��*U�#�ީ�r�~s&t�zq����Y[70��we����w���L��Mm_.�Ň�GT�V׀��Qb���?��Б�0%�Ɉ:;7 ��>��I�h����qD%��̪c�zjC���^R�/==Æi/{e�ް�v{s2<J��
�T�.8Ł1�\��}t�u|��;�rvq;�ͫK|�ftO���"���ǀ�;p�7�P�P��Œt��g��PCg4a�5����j���>y�]򡵂�%s|�sM>�Eӣ�]w��q+q0�W6Z&�tR]V��뜙��y�]��m\{>ۗ�ڄ�;����e�9���!*l�F���_'�f^I���%�k�Rxo��m�V�y^�n�ݙ�x<6�<�[�G7���<�4����=�9�"4EK96��'��TCAWsS3V�ۅ�	^�xwV�U�]�-;X�q#���x��^��E���5=��nt����������k�ӷ��M�m�!�{��,Q�"x�0�'��w��3μ%^V�?o���
M{��UΜ�l����g�K>�q�&�'2]d{��J*����x�����>����^k9����{�9jA�<J?k�m_P�)���U���a*�����3��g^XЧW��z�J�yz3��JQU	ϓ�\�})¨$����1`vh� VP�@;�_�.?%�n)i�jCӗh���G�db��Tup708���<�z��,�5tA�8H8i`����[K�|���8W�9\/.�k���b�>աWz
�#��~/:�-�u,ǘ<-I:z�4.�:Ixʫ��5�a��,\�oUX��<-vR����U|ob�d�S���挣�'zx-���
�r��np�5��5���rۉ�J�F�"P��T��.rw�X�jK�U��r�gi���n�V5���J�S����mzhYtn:M>x�5�Զ@�|׫�������h�r�TY��}P�<�b�J<�.nvX5{]1S�c�D�s_`{i�Tf��,�u/�b�d
]K���Lx/���İ<��������
�U����x�ӱ��>�]Հ��*��F`��+�rL��d{�o
�1uf�G{�q�	 �͢�ͪ�yBۻ%ҲZ����T:�������(�kr�j��m��)�7�TGck�σ�	UBb����#����[��躡�_QGۜ�+&2�(�
����i��}�SHU]��G<p�@��u�&�]#�wf�R�W�n�c��-,�x�Ǧ8f�W�;�UP
f�J�:�*X�OX�Yj���.��z6�u� t�zPH|�ؐ5uע���CQ��̔7)���w�<c���{Ë��c�)ܩ��4)՞&�0w��A߮"��Ck˭Ú�힗+���彗>�`Q&B�7�u!�ꘟ7���TDu��6i�B?n��3Ig'~�ꎺ�z^��v�;��X��7���"��C�����F����f<5f�����GoDW���ܨ���o
����=n��� �y�E��<���2����<��rk���6w B�t'�S]��r�s��	|Ŏ�:��Ȋ��Y�j�O�Y|�N�k�=����������{�M{5J�Zq��#��c���8��wm��]�I�޲��k��Y*liQKD1��H��:���A���4�7��PJu�E�v�`�yL���7]=�V�.PA�p�ت!���J�zRo����`�nS�^�m��C@V����|#Kt���>�u����hU�ߙ�
ML��B��s�,�s.�����V�g(���Q�er�x\>�o>!p<�v;�_pr�ܰ����l{zB1��� ��ͩ|��V�� ��.��;��\��eZ�ɸ��cN���5�v����eR(��]P��D/�>/>���#�� =PL�<�,�s��I�<�]��J<�P�Q�*Z�zB4��ߌ��0&���8'ܑ��Ėdƶ�޿	�n^��Eg�j!#۩�����^+����]�<8_�G�P�K�	2��٠���Z�+7�������Wa�U� �T��ah��Wq�r�����J375U9�)@ԏ$�/C��|����]��X��'(u�G����y�ٯN��p���!}����w������]ݻ�%D0Ir���o+|f��J�G�ƴ�=ɝ��>Ҍ�*�x��/�zT��j��L?o�[ԭ���ys�Y%�˺Ia����|1��+ln�����֘�:�.8m"a�׽�u���!����52� ��_G��fꃋ1S�,|��O���v�˾C������l�%C`]�Koy��xiߪv����ޟ}ڨF�z���Yv/Jɟ\(*�}r���2��xf�ӵY�1n��(ռV}^:��gx�<~5C���G�)�=�WX�C(�_qd��7�s�&-HC�'�wW�(����-��Z>��uܢ�ʽkۼj�ݘ�5;MȧƔM7�p�������Oz��g�'���[���Y�����m��D�~s~�1´�7۳�&ȸ~3������/�g��߄��kL���E}�pW� ;{᭏
���B��z-e��_��VM+;pM�A�f*������[�]�=|I�iCE��>�"9�1E�hj�霒�{6��%�u���u�0q�Sݘ!�y+��T�$X�{>�uV*,���އ֯�g�EZ%[��{)����x��VU��q��_��lW����"�X<r:,�P�����wu�q�2�UAJ��
.+��/fHtd��R27�_q�R0��P��f8G��Y�u�A����L���U���(������m�ϟLT�fG�Sz�v��_����&v�Yv�47ң�w�:��8�U�d�뾷\;&�<WO'k�^�n�X�"/zlf�6`��u����n�u���Mz�;E�(��!��37�´�u9G��Nb��/N!,��N�V�P��O��;Nj�u����m\���c�ӥ�ɂ���u"�]��+r��E4k�:oG'٘n�\�мr)������K$R�T������՘�j�E[z��&Y�C�wݔ&��'�y���-�����LnӚR�K��j�=�i�4��ܔt��w�h�u�BCYι�1�6dM��P���t�k0�¶���r����Qu]+���b�n���]]�n����y]��<���a�2GPJ�.BI�vS�2,�ל"WWA�C(�V͈��y�����ʖ��N��thE]����ػ��(c�����/.�N;�k�1��t��W�cp��N-�u�qE(٦��&-;w��c��}LT:���޶�5}�N���;�SɁݓ;1��FsT�Su����u�{F��ݺ���P���\p�ǧr���Tղ�MU�ǧh��y�k	�T��L�hFm�1b��c��Mu����|v��سt���L",F[��۳u6��I�l+�@�;.Xs$���<����X�\^n"��:ٛ�E�*o,�Քk��I$1�Pr����T�f��y�)�}�m��&��`,nfPO�Wl�<ުy^�K�M�|�]P�9Ӻ�����(�)ư�\T��ს5t���R!�a|���a�D������yJ�|����Zf⢓�DL�F�}��y��(k#&�-�'EC$�/u\���QԚ�[\�Un������WfP���厗a&VkX�;r��Ria����SG����gA��<���zD�!ҽ��f�:ɜ�l%u�d�z�|���.��A�Y�7�\�qC�Ż�5\�)N�8�D�� _A�-e�ڡF�+�X�ffڰ k�`�������F���颍m:�����v!i�ƫV�lѬ'5[T
��8�nX���r� ^]�W��E)ƺ;C��zm1[�޻���r�G�me�:j��`��;(�`�S�	w�j��ݟ�o��,j��f��V�r�˫��p/>���Н�3}h�LS��EwVk8��r�'w�~���^��W���/ml�+k6�������W:i��OwA���(�O��>Q�m��s��4��^�S1@�6���Ӆc읇U-��87/`G�M��-�$�sX���ۧ\���$�R�R�g;��]��9u��e ���\�ni�\P��E I&�usW�J��[��\R9H�S	�
wW@G>ܹXri�[E�r�=���Q!on<�ngn���f��P˭�n	���a�fv��֗dz�b6ìroj�1vÂ�7q�}�8!�<���pP�702�D3�sϷ16tl��N��{UJ���J��u�9%n�mj��Y�f�7Z�V�IMPS�����m��(��(���Zb֊����&��hm���ACMQF؈�4�i4���( �j���4�B
i���������������@h�*���)*�"�h����i(TP�
�9I�`��%���5�Al֫Ze�.���Ӣ'BR��C�t&�h�4n`4rj��)*��֒���F��Ji1h�%��Ƞ��N+b��J��Ѫ�!�4ljR�(9��KcK��F�h4����`��i�ִ�P[GT�u�AȠ
i��I���;5������QI�4EC�EUt4�@iқcli6���4��t���kSEQ:�)�"Tl誡���+F���QZ4�U2�%��S�g1��|�x�0����t7@*�)���.Y���1ܤ�5�c�j��X�>Us����^;�{���
����R�}PA�%Q�&���?O�9�ӧ���uK��%t�����������]���B^c�y�x>����E������"#��)�y��oݝ|1�\R�=ݺ�E�}"$8>����^K��o�=�N��]���oc�%=Gg2\��ɠ?F�
<��G���O�ל?��=���?;���?I������w	T������o<�ܫ��#r��������@����ױ�y/o����K��a���p��.����8�4i�<��ߘM<���z���uu%%�g��|�c���~����ב�A���{�|�t�w�V1[�/|��",}"#DE���}�O�~�O�<���!*���t��4�g�9ט}��˩y|<���w&�G�����ph>���z��y����%�俣����^�<�I��W�wz<���}���]C��8��x}������<���}��_!��~������y��?#�J|��=�ܝ��r�_u��A�u'�~�z�-:z�������#�ۓ��^u�����8U�K�%�̊��tt����ǌC6>A�%���luS�]�b?K����G����wK��A��'!�{/�?����&�e�<����}���{�\���p:�
}�^={˝����V��foy��q��|p��Cf<#$�:��r��O��9�|p:��|��n_d�!/1��C^�������y~˹��|����|�N�|����(}�G��]/�_p�y~}���l'��V[���G�`����������G�s��Γ��ԅ?g��:��wx~?�u>����|yèJ|������P�O#�9�4?^u���>���������h���у��x9xp��7�Egv�������{���/��y}��4%����u�|����~?{��=��t���e�yR���<��7��S�?nOo1��Gp������N� 䀿lp�W�9�8�n_\� }�G��~�~�N���sއ^��佾yǩ��^{������J��w��{��������ʟ%���G#�\��w���\��ʎ�e�?�װo��p�D����9�T��1����#l�Ow���wk�:�G�pq�J������@�R̗�9�������2��J�>:�`S�M3�%ح�s��JL��WO�j8c���'��L1m�[�;L�]��枰�Ȍ:,��sr�puc3����k�V������~��w�����u	_>p�^��M=��������S仙�sN�$�y����x�S�{'#���{p�g�<㯒~���n~�����H��GǗ�Bv���"n��:Q��4�F��-�ϐ�:y�K�H��ﾐ����{��:����t�@�q4y�~O��%���<����uN�v���e��N9�P����}��? �%��4>A�����9������i4��?_��<�G|ǰ�y/��?|��;����מp�?��F�y�:_gO�t��~�׹��G�Ĩ��eXQ�_xk�q#�?�C����&�C��ߞp>O���o���N^��{�(
(?���su	y���^C��/#�|a���/<���y�=�S�]��z�w	Q����>��T�^c������w����S�]'��q�ǲ�r�������/#���'P�5�;��'q��i�{�]e��u���.�|�5Ӳ%�y����s̓���D1`���q>+�w�����G���_<��w	A��x=^I��Þ������e��{�c��.�>{�e��t|��'0����uK˞a5��w/Q�|�]O�c�S���z����C�槻}��Mx"G�ܚCӭ���r����8�S�'�|w��G!)����?t��g�9!��y�?�����=�|���^��y���i4vy����y ����G�$}�����וy~�,P��������!.���>Gs�]�^p����]v�A�e�<����'���~���M>��޿u��z�BW�����9w ���(���o��=�_���=1DL�^��7��}�}7R�9@i��^d��r��zl���r�z?K�O�t�:��u�����q(|�_�����G�J ��<���;�i�y�z]��uC��}�7�EKuynYW�����U��>��_0��������쟻���.�߸z�#�r?����u	O��'�u���9	Ga�=���`�?|�u�{����p��i��}���^C�yy	���#)W~�ۜ�Q�&c<q�LԐ3�{p��	v�g<��
fs�Ǩ�mp]v��5�m4�����S���n9�1؟yh���{dsVF�>���Iލ�7�^ԣ$�N�ď!ݛ���vR�t�G4�=!ͺ+{N�,�%+75���7��1��rWt_�^��B����Ɨ˝�>����=_�W����.��u�Ru&�?}��|�G �'{s�O�{<��1��w	O����{�g�9/�w?P��D}� ĭ�u}T:'�G��Յzj��|3�|����q��m ?P5���I��켇��?yø=�W�|�}=��p�[�=��w?����|��y:~I�c�}�s/��w�!�|����?P�|}+�<��X��_��7�������~�#��;�S�O#�r�#����KEG��~��%�_��}t�?�a�켎|O��y�<���!*�������A��x�/*~˻?pc��nO߼���<�7�;��|��������5�Ov:��B���u������&�����_��7�O����w�BU����C��O��c�8s�<���z�F���`����#DB#�T��kpU߮��_��~?}��O�u�?����`���yN@F���c�g�^C��w���ݤ)���>A�i|�����u=ˣ�|���z�%%:]v}�G�ܞ�A |���G�C"#G�[�痟�"UA����ʕ�ʪ���>�>B#D9�#�<�BQ������>��;�T����hK�>�͎_������I�~�K�>n����uy��<��=��/5��/����O�����������}���������������O�xà��������HP�?�/�^q>���&�/����NO��{�<��r9'/'\��Z(�c��!/2vw�OS����p����G�} }L�����:Q��'�<<�nޚ�DP�� !�WW�[1�������e�O�����F�e��{����Pk���㺐�����伎y���u:]��_������\L@����� #��T.������k7_����x������_O<��bi�I��x>Gp����9�A����I�z��Bu�hk�=����O��}����|���<�SԻ�HW_�¨�k�[ f͛����}ս�����y�z?ӥ���חrRS��6�?��9'�5_7���?G �<�����	��u���c����~��<�g�9y� �����y��\5�
��j�U���(�tV�����.�_�7����6oM�A,�,�#�x�	/6C�����#�ښo�N�[�C;& Cǲ ��(���ǽƌ��`�D�����l�����<5��[�Łt�:�����`<�]�sCǸ杁u�x��CSnM���Y�_X�کhvmN��>����C��^?AT�r_�;��C�4#{���u=˯�y|��}�?o����`�e��_�uHP��<�����G�=��|���rM�Sܞ�$���˞~�����ϲrk�+�ju�b>� �� 8sb0DX�=��9=O�P�����u	O�d�������͏�w�z��������OS��������~��u�z�Q�x���� � ��^���uSx���Q����k�8}�?|�G�>�l�oק|愧�c�=���>�r9���f�:�i�>�Ϗ8{���μ��N���9'Ӽ��b>#�B/2c�>��A���ޖr��^����=}ݖq�����G��ʾ��~������A���v��<��C�4��=�|��{�G����nIIN����c��?A�ܩ
#�9�1�G��A��tѝ�J��v��5��
_�W�Ǽ[S*3�Q������Q���<�K.ƅ��0�h�7(h�g��oڣ��?R���*՗<WÕ�ucϐؚG�pgB�)��`�8��Ý0�O��vUZD��u����� a>[n�6/	PL��<޳ۼ�ݧ���X�rWNG�=��\�X}�x�l��B����Y����(X��b��w��;��M�E�U��ͩ�{�w����Y�ǹ�<q���+�^A�����ǅ{&V�GI�[�(�������;��G��Z�&��3J��ܺ�<I�iCE_�Ȉ��=�Uc���^i=����`^d�'�S�.9P��){d���,�l�B�'`��9nR��k
��QKEݍGՈ���u�<���wQB����w�]��S)d�	�%�ڏ_M��-�|�;�N��Х3o:�#�I)��0�}����1rN�ᯄx����y۪������S'~���g��x\y+�[��!5�pq���ެ�}��e�~֝,��|Ǡv���,�*��~��va��}+P��{�/a�(�O.��C��>��S�#/���A:��������.R�� �O6T5��e|q`��C9��7�`��.M��8x�t1\��5l�F��ثF�B���%#]��WW��Ժhq��pmnj&�����`dS*�SZ*��b�Ň�ꚪ�z���4�7%9�x`��h��U�ٙXOR&. !��IO�V�$@Fi���$\�R�Q�9^�J�՞iq�Z��VN���������D�G%Z
�(�b����kf�g���hL���UpcQ+��|��� ��/�R9F�:{M�-��9uQ}<��q�eR�]׻�cěVV�A�UJ�Δ-�͑��;8v�^�xAm����<�pw�5��z��#~���f�*�����h^�ʅ��o�x�0EW]z�^�ON�/<�F�u=��+��Z�j�m{wXV	�<=o;E\��K�9�)��ދ`RB��nޮzjEY�F:��z�Z��
��״**�t�	%D��@a��N�����4�kz*�V��s{frV�����S>mI#������Y�3:�ʈ�wX e�,st{�����7N̛^�ɟ�̫6������+	
��nW��:�7/g �:�h���+�ݍ���� N�w�e��"v7]�g_޼��`+��O���/��5��K�N���f���<�/b]g^�~��U]�^Y0HN�g�N�=7��KՈӦ|N��u�V:��X��C�gz7˩E)�����S��pS�P�n�1Ogғ���gڱ`vh� U����ֲ}
�l-�V�xo�io�k��������e��B�LOO}����5�N�9�c�8kcU�j.ʠp��f��*�(���b�t����v+C�Zp��(r1	�c�:FW���~�37,-��t eJ�x��g��wI�;U1+���$_T�����n6n�ys��=ȓ�S�d?vT����[f����a��y���{��ʞɞѡ�w��nMS7uw�:��ȏps"|'X5��:��;����E�7}FNZ﷗�קI���۾Mr�G�Y�|���e�	�f�ѝ�LW����H���ڂZg_��[��E�r������R���e��q�`��^Jp�s��+��h$���v����U��Y�]�$�$JP��7�6H�l����lgR�r��'0�8`��6�*�ݯ�7�D'�՝$��S
a�kw��wf�/N��Ty��%I7Bzs&��8���y{kWZ�S�`7���eq���r
�Dvץ�9aT�)�}včVEӄR��}�=��Af���me�����7�V��,�r�e��G<p�K����l�m��poZ��Ɍ�V
����/�?�k��/Yvk��ٲ}ûͱ����3}4h�[�n�Ϫ�����8��tm�x��5��f��3b�^���b�O˖m��OF�������k2P�}�<\�<�OyS�ƅ;<M�`�E��:��+��]����ݜ'�JND���>J�>�����u4��P���~�k���b�6hf���nge{i�G�)^����K:X�ؼ&��P�xVWB�y�%3Q�3�m[i~��^��]h~�l��%���֖�b|_�������CR�՜xkx�8).�vF��������Ġ�(�+�؇�+En�+�P+	M/
u����CTz+�����L�w �q�G��׻�/�mV�ŗ\;}b��m���0�upƖ�A��]>}�
�ӈ�w����j����� V_͒��>j�X��8i��f�����g.65�aPR�	��W~������3\i��G97Ky��r/���u�mt����ػJ���]J�f�. 39f�XV�KX]�&�gX|����� ���ռ���|5c�yK<�>]�STC�y�S�����=�Y��$�7�"�!��m��vj��qI��^�y�����]Er���T�c.<���Y�#.9]��'��3g$��Q���9d�%>�Ȅ3��y����g���ؔ���]]?/nYu㧆�.����Tz��P�j�q�.ꕊk>�Q�C����Z�_<���'x�w�,mc��p�[�xbs���E��=��c��<����B���{�Z�ӵ_nץ:�����^3S°�6j�z�7�ɽ�����]�<*֐k�Y�-y��u=ϮBdUe�t�-� E���#��V�r��y	�*\��hz���"��n�����[Y�w�"Vگiii���v�g�毯XzwC�$}�Zy�#a����R�£���*��~�D�|݆��lp�ǈ'`-�!���T	$=^9�ps�ugo�? �����ʩ�ոe�s+��w���AT(�>����k���{�~��|��fny��c�ٿ\�S�X�\���7��n^蔔#i�Z�1��K�WX��/r�&½�X�����9��e�csVV�&�]B1�{Wg״"��L>���C������z�M�?��RX�U�2r�ww���ᰱ=��'��%Cj��b�E|i���'�=h�<�-�sݦ��x�U����z�z��{�χ� 5�$LC�M��(�:H�Tk���Վ�ճ��->&��L�]xK��2|��4�]e�k���U%��Vl�<jd��ϸ�`�	�i��N�/�_�À��^�Z� ڔz�b���r�H8�뙏�����>��eǹ�!-��+���*���ʦژ��ǝ^Me���n//6ye*�s�P>�%�_�t�7��/��>�Ȱ������s,e�@{���f�=º�1�)�C�S'~���<#���]�[�*{GI=D��J��ٗ���-��,�T�����vX,ऎU�M�#�ن#�q�Wz,���d껊�v��<���h�� `�P6t���Ed���r�my��l�R�]<��o-s�r��W�\C��p����n*!�5���ut1��J����)�g����+Onv��'rFc���\�ia��/�Ui;XXM*��z�����`��[.�|B�Eczm/q�v�n����)U���C�I*��y�V�,���uG	{�U��UX���p�Xv?(���4č�xp;�%��O8^�r���T�����Ɂ���s��S�y|W��vie��{`w)�阥/W�wQ]Q.{��ΫY��Cy��{]�����$h�+��p��6���u�5�v��]Gή�Sba]f���������	�$F��Og�=�:��	����=����Դ�9/�����qw�맄L뙏w֊�z���5�r��l�7�o���E_O"d�ܕ��<ع��$LM��[�?kݼ��<�b�N�9��^�������ϻ�L��Ͻ�k�:��=��IYa�ʃ���ڼ�7ff����ޟER�+�"�ciК}K�#�]Ha�J�y�en�j��f=+w�U��ח)dW���ඌ*��9�;�%c�u��q���/�xX7*�g 9=nq���U�Gy6�V�ׯP�R�{E��,5/)#�tY�nF�����B���>��QX�v�!=7=�qѾK��7�gK ?U^T����Ћ�ɂBw�/��w�����8a�����v���
��bM�ż��¾�F|�`F}�나�P��;P�=�J�%��ϸ�^��,���[�=�]{�<�yn�h�	h�M-�Sg0�:쿖
׎�:�_�[�螞������MSi���w�C��x�x�8�¸4��VH��]NT�vzx}+�<�_���m�E��]p$� 8jN�&���c��Ix�������s�z��W�=oV�m�ܤ5b���!C��<"��Ք�t*Ћ�������D �qw�.EUѺ���b���`���h]�Nv�3v��K�G�W��z���'�������1�p��Np�G�.�3�g.��W	K��)n��i���"0ʷ��vl���=4	{Ƥ�H��zD%j[�\�E吳|�S��؀Q�,��yo����҉#�v◵��x��8>�,s���U�"��V>R�3&� c�Q��WV���&���5���r�w���Ř�3Y��C�-�M�ua�d�n8��ŀ�Gy�� �]���mΕ�_V��n�QL�9h��O>;a�-4�ov�Y[2�S<���xY�q�,��>��0�iQ8l�h�ȍ�;o���*#TL�o k�f����j��;v;�ەX����z��!w\1`8�%C^��j�Km��A����L�r��S`h�Ä�AT���g���x��&o��m�zYT�1�m9�v�I�4�)wVl�V/�"]2�,"Gܴv�����ĠL���X������5sD�V�=#B�yaa�����ҍ(ڸ��$pP��"�����Xw%�D��#���k��,�bs ��m�a0l�e�pL
��KB�Y²��݄"��[������杻'�ǣ�F�l+�6Md�l�uͥ��$�w\yˣ����(~`�s�Y���z�iK��p#R����N�Y*���{�4�0�ܻ���n�]�e�x34Z`tH�+b�?{�Y�t#���ARܷr��� �N�N���o��rٺy�:v���8Yy�>T�\��m9��Nr�z�s$�-����-x/fW���g��;�ڬ��tԄg�T�hرp��V�V$kh��N�L����4�;Bmjj��M���˅c��\J-͆��(������ʹeW�*�;,6B7��kA9����Q_c�i�Ǜ�,#��mmn���{7iH.�$���x�W�[��8Н�8�u�f� 7h����C�f&ށ���'f*˦�4��>R��ߴ9���fW@��}wp�d͏:'�i�E��Pa��-|��	7p`��ge`�\��7h�/f颥�4�4r���ݮ6��4�	{�' ��t�+v�A��B]t��{�)��������rJTCۙB��˜�YE��
ըͫ4�Aq$2*�ܽ�����\�J%:�1��	&��l����EB�Ǖ�ka��kvU�c����]o/�]:-��묎��I:P����#��tZ/��ùY/Bto�f&�.�����2.�����tΘ���y���qN��F�D!�r�xwx��s�nb�}J �%g+�[݂��>�0\wW�����hl��jF	q]a�]���N�\����,�k8�짦�U�M�.V/Db�n5^���O��_n�� �9����V��F��P��,������Z���F�� t.��bh�[cZ
1UQ&�B��D��H�t��ѥ��B��4:�md�T%��@�i�4PPPPR�4U%5LQ� P�LAIl��l	cضl�t�b�4���)�F��RQE,AT�%�f�A�ѥ�WE5��R�Mlm�4h)HkF�أF� (H��[Yi]�4hJi(����AI@DR���CHP[�Ӊ(t:h�u�P�it��K�H���m��JM:t4R�����4�M�U#P��
y�)��+���N��)(y*�b��AQA��*���%)�h���Z-)APSH�7�럾}�]$>"vDeZ؝Bf�g+��K8��skPyoL����H�ͦ;0�9A#p�W[���(h��%['{ꯪ���)�a1h�3w�r�Q�|;_�Ƭ�p\p����P;��GʻL�/G�j��P��=;3�����ۛ�<���O�쐍�u�xK
��s��oնa�+���3~=Մ�:�z�u�����s1m^|��X.<�
��ȏw�c�O��`ֿ��ณ��8ҡU�^��'C�|�l�nb���3�<�ݳB#������BD+�BJ�U^52O���u��P^�4Nxr����x�M hn���ktq���TG6�YNXT%x~����mS�v��\i\|�'��&������)�K6��%]g¥-#��7���������;��\]�/@Cxr����C��:֛'0����e�V=[n���u�/{�Z~�[���wnm�M�kT��U.�Ir��b�S��XC�7V��7���=�P�]zc#�!�a�Bʞ~�җ�׻]Q��V�~;<ǋ�Tǖ/x�Z�B�q1}`�x�v�4�{�{S�9��k�3>9aP��˭ý�%:54�o%ϗ]D��~y��`���`��^�"Q�mţ8QPd�<�+����Ӑ�s��������q�Q(wd[��Y|:ˮj�t�n�v�wj!8���k;]����V�yRG�-!��)B���e`�.�NqR�\����>�,,�_qR�wb�{� �ui��dL���}��_U}�}J<���w�7�?�.�/f�q�-�����al^G�/0�u��?|��Fi�M���,���V�o;�'ޔY�=����`�A/�Ҟ��f������:�TFi�<����Iu��ҵm���f�;���V(�A^�<�7h��p�P���{���[���`w�s�s@�����~2
NX�Z�hت*#����*�Y��`��VJG�fA����iy�s����xW�j��K���V�Xu�ٕS�$�ӏ���Lx�]q%�o�j"��W]_��=����Q��9�U������g>�R������mHˎW+��� r����Q��^�U�n#6u�z�����Bq�3����3��)bR�}�c�_�+��-��S��U�s��UV�@�R��,� j��Q �:>T�O�*[����w�gL�����yaR�����=�(ߪ�$����#��4�hҊ�;�ԮS���}����;�Swv�yd��Z�F<�n���ʖ֕���%[�T٧�8<�g���c�����<���"����,�	�Q�P}�;���9��봡+f�Q����M:=}�J�
ީ�۲4�[���Q�;;�ͩ�Ʀ�ik|�.��ڰ(���s�ݻw���0�}��T43�Yd�c�&�mmr���\����Wj����uz<�y��^�G���  ��[�5�JܺT]���K�T�U�p���uZ8���(��5�� 'ޓ�[��S7�1�5i]s��SrS��J�D*9J
���*��ce�>�:���y���7�����4%\U�w5R�����`s3��
�M�V}���v�4m�z63��T��O��p�Zϻp�aހ@����S{~���gz��s�Y���hZ���o���S���c��F��+�Ԃ�[�O�*ф�c��tz%h1�
�k{�^�R�g����~���~��rN�¹��'�h	\>��N'f|_0<*��d�>�a���֧%\��wBS�/�zM��f8V�����M�\���	n��^!�v�^A�֠��=����h�`˶�K2�
�,�>�%�����j�j���[��0�xL�r�Gؾ��k
~QWk�{�} �$9C�(pk~�{�)�����Ov`p�.<��o���'�]�w�ǭpNL+�b;�h$�6�o�l�����6�g��������kh�5�O
���%i�`�T��M��p��Qn�P:�Jּ�%[�V�e���g0gG�ֺ����M��mLV�[���l(�}Y��a敂��'�h�����r���T�\�-�Mˮ�3�> c���-��#)ad��O�{���;�������r@�3~f:������ h���&΃P
#n�����)CG��b��R4½^9�N���ȼ�ݳ��ذ}n���"<^�5�*X�X	Q^�ۡ��*U�:#�b�b��y��׊j����\�ߜĉ�</����`dS6�M`��E�-LXn�T�ku;�gG.^�}����yu��)U�ń<5	*�.yz*��������u'��Wf�s��R��G��r�ΚucܞN}$�����%q��o�z�%Uy�mvyn$�b/\7W���n��F[g��Fl����m�q˪���L��^�*��ߒ�f�uj�vod�?yJ W����6�S�h��5�~[���������"4EK#]�����7��9+;�ŵ�x��Y��1PU�ʫ9](R�b������F�ο[���go��	���������^��ۂ�y��p1�%a�s'�}��]>j���<,�9� p��J��Y�� 
�B9yX3|��U�(f�c�ۍ	5x��k�CݵF�_��z�����eiʷ�r�ģ�Ը6�׻7����{���i��#R�)�6�(�Z�d��}��򖩆�0�Lk#h�P�^u!��;&_pR���H�].jn���+�yZ�;��v�kh�H`M�Q��&.V���;{����I6����}�}�R��ӮFz833zN>�-�/iT$O���_��7{U���a*�zJ�Ψ�D�N�����|n`�ḋ��f�J���("kzu�������tFe��Kk!���$�F�*��eTVIOW�K�4����9�i�b�]P�|<񿒞G���ڻV��#Bͤ��^�����G���żD���p%�D��+�r�����g)J���y��ș]��kF��.�[�Ո��c�v��� #�>ۺ�H+k��;d��"�p�)y��u�u���d0:]i^XTt�s��WÕ�l1Tݰ�=���z����sy�]�!?|�|���/�'��{�����B�&���Q��q�5+�底�'�p}=�@A7���W��A��>U�W�ʻ��*pBG�W���$� ��W�M[����v�~���W�T���=�4wT$U)��e��ktW[�¹Q��K.�J`��&R��3)���)����W��V�G)Wt����r��[�)�Ğ�~�d��D]ɴ/�%�o</q� �S���]̰ov��װ<���59��G�C��>hѱGz�"rv��8���;>�C���F�'{����iO_E*,휆25��zctD�̹��L�z8���A�L�_P�����I�V��p�(命N�-����}�}U�u�I��QD0��K��g����T�\+o��3��z���9��n�LP���i���>������t.8�:f�9JM.���U ��p��[a {��r�I�F'
\�n���w��uB6�-�0\U��T�\v&<_�!�k+�TƦ��L��q��V:�:��<��2}�#> 卡�������� ���!q�.����ףU�spxur����>'�;G��<��0��8�����j˄�Z@�N� yx���#���ʞŕ#r��ie�Rޏr�u��3Z;	�~�.�����/3b|_1�Vqp(c�Y�8�&(�Av��bG�i���#��'�d{���
�@�p�����:��q롉�tx9�z�=�z���˼�k���T�&J9���*��u�mq�����k���*xW'7{G_�ؤ��E���]OoBl-�{�b���2�t��ҭ�*cĳ��Ix�.o�T'��u�s�j�����2��.���ؾ|�����~`{�f�2w����a=��m�;V��Ugv��f{��e�-E�`��b����Zݞ
�E������ +�vfJ�����z�H�;4@��o�&��T�\x�-"��7����M�]2�̝�wZ�����JPUә]���[��j�	��]`�5xq�[�4���}_}��D���C/�b���\k�ә��4t?G��H�D��9uAM�u��|�k��x:Xޮ���C`,@��3>��v)�����P�*h�V��y=!	�1��u�����j]X�F��ݺ�^�c�r�Iŉ�$x�h����B�wژ�>U�s�år���7Ҳ]���Av��7�:��nxà��K�9���۳���V��z��Z"�`���eN�r���N�ۮMeӠ����}H��
P���*������i�����P�xVߞj�a�N�i�u��w�P���J���YڕU)�괸MYV~Q;��{�6T�*b��T=���{[��{����\����|��5h�U�{� ���~n�`�*^	[�&o���Q���6|-}���%�����S"x�N�^C�0����%��Ľ��ָ9}��{�>D@auX|M[�\<�Z�ѫg�Ai�7+{V{��*�<mw���B���NT_j�W�y�ݛm���L��:��2�}�<-���/��g��7�w��"�C�i�����:{Ke�e'�f�	���h}]75��+=���s�u�ֽ:��ZS"����k�Lm�w	���Qb�m+���ޭ�X�x��5k���RW�p�R���SVgv���8�E�"�9$n�Xcq��"D2A������}�[ݚM/b둀nex����K�L��L�M�^�-�	o���`����e>6S�縶H�V���1�eW-�*W�%�@k�%������U)�;��-��0 :�Ҽi���&6u#>6��9����}����)����Q�aD��3��z:��aB�8Le����<R&�@I�x
�U�iq��cTQϩ#�x��F2a�`~����<�=yֺ>�q��,�9���u4"x	:|
�y����)CG��Ҙ�J����h�S�U�U��w՘Tj���҇���uº��@�tP@�a!���J���i��<���#9�E�~��x	�Z�s'�N��³%���f�4)�x��jb�0��kxK4/7f>��.��:�Hpr���|�δK���[P�L�	�4g�0�G�z�vWZ*�O��=�����y8_���A��tK��+��G�z���pT�/�X�Up<.��r�U�^j�];����^Ӏ��7'½R��7��o�����+���L�J@Ŗ�=��B0�/���==�����Y G�^z�:��Q{��FٹVآ*�?e�ۢ��pAQU�.��8���+)��Wn�T��~*rzb"Į�ф����٢���[דU�]f�[���٩����g���L����$�폝֪fZ��W;��W�W�}�[Ժ���"Gk�ϥ�Y�ߎܡ�_�߰D>_-�}z�;�6��F�wx�+EbT<���z�W��_|�Ζ�_{�Őj!����Y��o)_]yj�H�.�tu�+�'�{�����i�ڃ����Om��{M�V���6~�e��q���s{��Ub�u뗏���ފ�Fm���UX�S�oU-S�t��7�����hI���B���1�{Ս�̘�!-#ܾ�݅TLD��N��k^5��쿺+�q���}���|���Ւ��ݭ|�b��J�.ޜ���3����0S_
2�8�O�#��d�n^��|-A<�ҿzb���$�:���M/j���F�v/�����]��)�e�ڰ�{�"ݯ>���Z��p�9tA�_VI*� �	բ�$~|�@�j�_v=��g9ӻ&g������T�[�Ud��-�C���x�'j��"��;NҼZv-�\�.��/fv�Υ�zhCQ�m���.��K
��s��mm�Gܨ�*�(W�X��j�MN��,�/U��w�^��Ё�Y�u�� �Շ��6y�|+���kw�<ȥ{0R������LR���W
�M-筨.7�ۜy$QwqTv6�;N��9��9*^�=�o5�e�;!�Nu��L�l�\�n�"�0�k�V��| ��^�|���v�4O�p��|���/�L�
��r#����,�#Ԧ�	��=' ċ���M��۪_UU� �('��|(�3w�48*ϰ71��_P�雛G�I��w �dQ�g>������pK�]c�-_�"�HU/�֎.\��md����J�'�wr/���}��wj'�5�+�D��&5h�鄛�P�+iL�$��J��Q#�>�{�q�]^�"nx�����pxg\�d�,�_c����v��/Y}��8�vA�X<�ǡfLX�޻���ܮ�p@t��Uf2��2��ۄ�����kzpkWs.��x�o���'�Pk�J�u���+��
���<\�ʘ��=�L=q�V8���b���	ʽS���<=�ucf����Z\/��/J�54���8�d5���q����p���~����yDg��/f�>��V:S������7G�b��yx���ՕЪg�<r5�y/=��R^�����~�#k@NΝ�Ip��Z^f���cڮ���:UuGﱺ���KK���,��^��]{T(4\8�-[Y��^�39��:Q��w��Q3z�O��;vAH-�CY�t�I�b[
�����g��}9�H)c��w�2.�ٶ��؄�B=fXiVm��7,n�\nĳSi+A�,��_�q�e�Ž"�W䋙ǣ�׹6o>Xbb�[Kz��B]4*���J�>��[�r'Ea�1��/Na�\����	Z</��r{Ot}��m]i����wO��zě�:�E��Sh�f��-��[���ز�.��ݭ�Z��9@�lI���Mvt�[�N;����m��H����=�ه9�I�]��W��nj�>���#T"71���:u�#��.��we���)��B��X�s�+9�9���+	d�+��Y��64ˊ�Q�ۺ��մ.*�\�{���[��:^��au;r�p�q;=��ژ15M�����MẨL�Ha��9�P�b���n�$��:d�Cd�|�^<��լ�4lb ��+�]>�|�8�z0�WN���Q�O\ߘ���k��\Y<	����+pCf�̖KX�S�e��#tT��֗
��[�q�IP�@�os5J,���+�d���w]�)� ���d/�9�L�M��ŉSY�B����j�e�6����E��d�6�*r�(�Br9�����k(�C��e�VUt�2"!�z�iS��(�bM�ǲGW9��.���u�8���5���CMZ����:���:�=.9��Sr�t����\1�x���.�#�9De����<��b�[xjL���l-�r!�	�G�`^7%��K���[ �l�IY�z���mk����yӚ��^Y�u���>=�{oQ�ϗGe�u{ՠ����.s �$�"�u٦���pW�2SK�\z�T=\N���imbO����t5��⛽��&�,u�]�U��6���:]�*:�1�=[k[p)��C�'eM�F��]�Zi�\x(�É�a��6�c�P��z�������	P���v3ESۅe���ָ.��ob�B���Yf�Ї:&��x��E�h�:���6��ƍH����Rѥ�gyQV`��5����|���JeO�K�WN�%��oJM��v�kȋ�����o��z��j|\�� ��䑏�7���f�Gi�Bd�be�7/[�X��|fƠ��)3��#�_����`AQb��]ԎS똭�݌��- j�%�[�
�h���6u�FҠ2�6��wE�j��]��E�<t�[�v�b�;]���Ȝ<�k�c�A��K�b��k���t��6���\rGj��\��K�K��&�s 3�r�چvu_�pu�LR��Z��2�o{w����!�C�g1�*��ZUgs�*+��L����s��dw�3*��*��6�$�W��@p�ܾh�q�.�R�����C��t�#��;��uu�5��;���DwW���Ety;t�36�v^�ևo:���R�g���럷��@�҅Q@�t��F�1@��%	EP4�RҔ�)JR� �"T��t:;�TД��@U�CE4�Q)MP�%Ƣ�H�h�C���� 4�M�&��I�(�j��
�M.�K!KE �IEt�JІ�E�*Z�ih(�)hR�Zt���"Q� �!%�����LHQJRUD�BPҔ�d�����B"���(+l!@�IT���U@D1%�@�L�TKC@�UL�CICT��Ҵ�
�����"����ǎ��ݺ���8���;j�a}���1�'�re*{X8T�E��\e9�R��j��F�!�J���Ƿ�	ǿ��ꪪ��7g��{Z�u��㳄C`��ڸT��a����W���'¯�|�r�(��%�{��"؏<��7練k%-·��U�D`n[>�C�����9h��{��wQ-�W�0{��N"+0h�U��G{�^���*e�,7ۊ���,�(����W$�l_���r�y�;߄����V��������o&�
]B;�2�q����k[[kC�Խw���iF��5%�T ��_?G�7
E�%-+�����z��\��������h_��r� E-�0뤀�C��=㢥��>X�;�!d�w��X�-^�/��ÑӍw��0ch`	����9^we��Z����7ژ�|���P�����g3�ZJAY�׃��ep�;��Ţ{�}W�>t�G0%[��[f�8<��o�5��},�N�t���#�KÛ����_ou"W�
P��=ʢ4q9/���y������'=�h�dF!V��	C�S�+\y�>L��X��0��rbǙ�/G�OM9�gL;�bܧL��]m�����)�m� T�a-	��S�Yv��|��,ʺ�T��BڂE��Y���0y�<�,OSV�N�5����������Pzʝ�V��s9H���Z���B���35�7� u�3L͌��r�c��B�������\����x�	���������l=��8)_5�����*��]�E���Z����6w�k$�}��b��R�G[���=eC� �5n���{��M"��KTn���m�V���r���x��~{I��F�Lpp�Pi�{���?eZ0��˱�A���OQ�7�!�J/^�@����{@O=IhO�������U���ub�Eӧ�w�w�zX<w���"V��F�Q���f8^�����M�^�-��;�}����{���l�;�O��
����eTa]Ԡ�l�k>�jK]7%阪Wo���`kr�Yi�]�=��ɝ�d�Ĕ`Z8�����Qg�������G�=����WQn���@�UbD��:��;�U�g��媫��?�g��
9�$r����N���Dm�J��"o�5��eBYp���zm�|� h��:�����c�FI�X����t��չ�#�������9�a�Jz�UQ�:�%��X�K��|MU(�ʡ��|:b�V+����is����쬾 �A!(�+]�M����2����ab{ؽcN���ê�:G#�7g�{�x#��C;�;��V�m[c~�:���#����%B�^�9�7��B��L���{4	m���k����Bü�u�{
�mV���Y��_UW�^|�u��o�3�!�up�Һ�དྷ�z9V�7��q8ePo��ƇZE�Aa4�ѕ�ؤ���ݻ枌�l��ᗡW�k:Qw.�R���x"RS�3�^^�����\�7՝���53﯌٫��ņ�9W�m��v���T"RS���*@�@�z���y�w=��)�|�������WS����{VW˗T|zd%���}�B��SI��*�`�b�ڪWժ�u<*�y��~[}�Y��>-g�5}�
�ٷB�
a�<��Mg${����.S�I�^��9|�,�VoǀDU!��*���&���/<�~��Va��0ߕ�����n{�4����T�{o�<�-��Y�
�@���T3�b����i:��]���oki��-���(��#�hW���ҧ��کj���&7M�{έƄ�j�9����#%�I���=�4=C��n�z3= ��:�Z�����ε�|�� FOO@}�آ}�hי�p\K,�����g�z�����1R�=�v�����6��Z=3j*J<&1Hc�t՜��o1!s���JQvF6�y�Þ������t�?f@��9M�s�L�[SOW��v�g�������cP-	�䬑�<pz=���^Җ"�˰�۷��h<�^�]�a�n>�6Z9Y���/�)A+�n�U�=����O4ݻ��E)���+���h��LD�D��A,>i{Uk���_kρ�Y^�&7~�k'bčR)��^����ב�tQ��"2��pik�2G��4~�+��#3s��h��8e^��U-ש���Qؾ=X��,G	ㄝ���H��芛1 ���]y'�%+=]#��:h@�C����*�aoN��Bѫ��6���?b��t!P�ʬ�Tu*_k����
���:���d�-�1�S������io�B��j3U\E�@R�:������f�GK>ϛ�٨v�����I�9;$��U��Q�w�;����݊N�"t?���T&� S�U���h��b�Q���f�z�/��l�2%1w�y�;���C���JUpW)ć] ��V�3�\��<6��V��gz�|�m��c��T�M=��εYdg͹�B�V01�4�b<N����WP{o���T$�ܫ���M������̷�;N@{w�DK��&�?n?r��˝1�� Q�k0X�.�;{G�.���U�=�����}t�J/u����c�r�O<���{F���Q_-��vШ�r����Z�sA�
LC�v�X1v�XuݖU!�݊��s2>���q��[�m���6�4+`���χ������.�K����n,]򝝹��A-ž�k�{�4��jհ�[�K��K��V}[��"�^_.s�jS3�s���u�p�v&��ν�=Q^�� �l�t��~/�Mg�tU�Ԇ��lS�ݩ(xNϪ>hV���:6�l�K�=[xwB���E@��l.�lխJ��R���xp�]Е^��޳]����6{˔!����+����.����y�EM�y��{d.�����+5�7�8���;��cZ^V�yd҃4��^�	P/n!����J,ɋ1\���?]&Ψ���;$s���Be�8�	q�vC��M�`���|�-�/a�>�ۛ���	�&�j3U���-�罘�z�j߳���E7�]�tƼȮ��]�{�W*��=�c^ԋ�t�� �%�f���P�)�����O�ۼ�v<���/�W޹}�EVF��z��x\]�f�'/%l畸)�h_����D�����e߰|��0m3
��[����4%�G���J��ΰ3�]���J�>��֕������CFN,,u�}�ʘGɜ��҈������/�����������SWw~�G�7k>C�3%������7ڧ˳��mJ�f��d��{��/����]�-
�+C���W��+�*`��Bl-�peWv����R˂�m�OZ1���9�H6{�|-�뻼4�{[��K��+�S�W}?X-��|7_g�N�q���.A�3�m������Vb�er>�y�[��"����-����-���>ϻs��'1x�Kݞ������wD�h����ws��.�OO���g�}6��|T�v��j��`��S������둇��fMpsqY�Ok<}�s��.׿_�pU�[�2�]��}���q��{�?̞��b�gkf�|�����:��ƽ:e�Â�bt&��-��O��Thoz�[`*)+f8�1s?{�(C{����꼯J8�o-R��R�>�sb����¶J�jN����<�3-�]�~�V.�"**(��ս"O��Q2sH�p�	jE�5��@.�U�\Ў��1�d�u��I?���vFJ�@��l�ιljz�����m����_���n�����T�Q9���lpJص�:�b2�̲V�>�*�=�3���UU��[�������gU;��S,Ń���kx�I�6��c���^ɃJ;�v�vy�(��r�`��`�=���R=��h�[��Qέ��lے�JSX�UX���[�=��>�3�z�N�����������{����WO;����O�A��҃
݋�^RB�ʫ�Ŏ��6b(��������ּ�/m締e<��K��~7�k�Փa�2^3N��SʻV(u���9��ϊ��|��n#Pw.�:��?}U���I� ��~���=��;�����L��Ы��w�}���4���j"�#�+z�[�X������c=��ae>������g�N�q���;�]����Y_�jX})OU��:���:��}�-[��i>u��^��KP��k�cɮ����{��K�5��z��y�;o�|�^����h������`����p^�=���co'w��b�*:TQ�(�vP���Ա3�h��,�ٯ�p���j�(f	Q_P9=�+'
]зy�c�Y�Uº�W�e�{�g�a��fcה1>�+���r�פT�O5�ygU���[{������#�=�{���U��
qں�i9��~��>x�[�4��Z[Bv`���9XA]�ӯzz����>�N����C�����~�����j�-�,߉bS�j�j�+c�Ct�޺�g��ܫr�������%l΋�8�:����V���yy_9��k��T��z�,-`�b1�5[%bjN�:�>�3=���l��{͙˔!��ݼ�=�o�=5�P��Z�xZ;m@��I��F�˫��	^�c�O|֗��]`��~R�O��uUi��Z;Y��k�8⻨�,o-h]���^����U*a	@ԓ�l���̵�;J�=aŗ�G����Q��ֻ-t�MGq̓�W��K2��!�����=<���@�M*�m{ȵ��9.$��k��&ï�-�j���}���v���Ӱ�j�Pm��>a���o¦���k/��o˽��8O-�����$���j	��C!r8�.J�%���n!#K�	,�������2�I*��ee3��")Ⱥ�*q��aW'oC�ɋ+w��1TE�h���M���Kt�6�X+~I�ծK�M��	.�GG��}��U��i*[H8ו=�8��4�|��ϫ��nsH��o���I���R�cx�m9���ǒt�OJ��[�W��{��^�o1/'Y�wʔ+�Ϸ��N>}eR[S_j�%%Z:��q�2E�T@W�(+ESz�����Ý|x�nz�u�����,��ne���r��wc���W4눵(�˜�f�]��ߖ>�yN����n��}�r_zNȻ��c��5�ZИ\�>6}����V���y���ngݸ������F�5�jc6z+���r��~�:��n�z��~�D����m�Zŀ�)��!�f^W�c�$�ݴ��_O�i)����R�p���ݪ����K�:/]�Jr�"}�Jn�R_�������w�Qd,���9a���z�щ{זgG��Kxwz<c���?
�+>�&��^�b�����b��f�#њwo��������֦�8T�t�Ī��Ⲱ���Z3���#x+B�@��`D1��P�;��������f���o'U�Ni�0�f�;t��n��Њ�9E��@�c�����r_����O��7�ouia�ic�ʨ�������ﾼz�B�����X<�����
�7�N���'g�9�����Ҏ%<.q���ɫ�j�+�ಔ������}�Mgp�79�㼬E{V��O3s�	���T��ܬ������f)��+ϥ�w���5�N�Z:߮�~��tPj{�f<��ܨN����k�ou�`y���o"��~��)��t�����D��ʟq;� Փn�����]l�if��P
�oz��H�*EPL��xXx���=�Tȷ�9_>}���#�X��O�k��ף�L��7�}/r����|,<�px:�7���-�zUS��� ����p���'��Jt�<9���Aә��2�R�Ulة��>��V��>7v�E��>מ~Nb��Z�sm����&�z�Gc{�M>�K��d��=�3��I���x}�A�mP�K�}��'x�^��a�{=��2R��9-��Aw]V/Ndx/�\j+��V΢nS���`��)� �Z� �tpm����5� �S��U�;�s!������G�4�t�x�<�p����0�7��o�Vz��Ͱ�`06�r��<�I�TJi*�f����k%�(�b3���[n�wY)Ԥ@�h���k$�bv�u��6g
b+���Q�trU�H�ӥ]fZ���B�ָ7� �8sAK��_��z�Y����><��y��,�Ժ���mx�&Ed�=K��oQU79����*�ټ�����e���8K�5�8�V��U�\��:�V�W���W�5�Z����"�zw�ɊZ]{�9\{sH3�������(�a|�[��>�r�]aH�u7�E��q|����Ф&��0�Ȃ-�	Zdt�P��_.���saM/�i����sl� i$ؓ;�:��ź���p0�7��o����%@ۥe�v��ݦ�sK��w�o:9f�Zk�Z�P��ʤ��شz�!WYN�(Ą����D�2�+n��z��'�N��t�ǹ�t��j�����yy1�3��74�l3hq��O;��J��tɢ�>��c|��)F�$��8I�u�r��F#�k�g;�^g���1҆P����29%�X�}������m�A���e�l6��{O�:�3�[����89��)t�v��^}�_e��O�b�mS��K����kf�yY`Jon��[�
�D�t{0��()E3t	��9��(=|5:}���ʵxn�gvHF���ۖ��$SazVȋ�I	@2��]]�cF]gN��N��ﭥ�`[Fw;X���u#-�f���-�cg��^�����4��7N��.�G����^(��ᐺr�v�Ù��-�XA�9p�&�Z����I9�P�"�5rF3�zn�Y/s�䛄��:��d�@�s���-Z��s(^sΨ��w'V+��y��!��_�R����}H�m 2M�5���iv����cU�Q���]��Z�®��(��;�X/7����ϵ��\g��mɘ�`�,{��X����}��ݧ�"��E�@S}��3,��A�d���(�ȧ�l�^0�5`�뢬"w��.�]�x��.�%v�[N�Q|�ʔMͺ�Q\hVo+�ɬͽ.�,qyc�.�qv��0����Yv5��)`��D"��A��ǜ:s�tM��It��U2m�����ր�[��7�8�=�:�i�|2P*TV��79˵3,�uv�r�e�ʻ��`Xܮ|ۮ3hd�CZq�}����]��4�M���f=TTE�J&v�l�$��qޘh��	V��0Q�;^��q=:�
;H��r�O����BP��E&��V�N\���u�2�Yq�ƭh=𝆹�ۜ-g������ۊm<�k���-���[�q��}SR��a�{,w-=q7�L�^asJ+�s+#y%�����EE�M�)E��Z)hT����"D��������
@�)
��!�h��(JP���*��J
���l4�T�TM$Z4�%Q&��CEQKT���T�HRV-1%4�5TQ��EJUQM,H�kTEAAIJSE-%)J!M�PSAB�m���mH�RQAU&�KE%DET�$TUA@PA�U-R5TUT+T�Q����h""JJ���J�&���J�������PTE�%D�--*RU��IF�P�
��,F�(M�F�J
i*��*�������eX�4��7�-�2��K��8��y��ùg��2��̚*��v_4�:%.R��tG
�z��T]D-��$�]��U�՝�GC�x�������:=a��f�f�k��P{�s��A�Z\�Å��ޞJn�egw	��w~��˙�v�_)�R�2�Y;C��eK�\�ĥ���ݾG�An�=���ʊJّ8�zMX5i�L�=�j3��Y��	����T��_NNVV�u���[%&������^gv���ٻuӕ{=���͂-2�����U;ۈ��u�ĭB��g�/;j���+.�^`�wek�}x�X�M�Wi`�Q<U��=����O���{}/�{-�]MϽ����>�7�]N`�%���Ou=J��7��i_� ��+�|�F�t�h��Ŏ��6~(�p�V0\��9g�w��vԤ����>�>�%�Od�wV	��	�UR����V�N�������ݟ�������o�C�xT�Y$߮}/��<��]�U��N򵶱l>ݐ�wY��\�0SWy�4-ڧ��*��|T�TV�����*�>���QvW"i%�ڄ<��:�vGf%1���v�wh%��5�n���c"��]'W�69TF�f����j�������ۋ��Rgu����^1�ϭ����>U��6��*�|��̕�N��.��ܷ`�Z�J��`��V��soS�	H�l�=�W�����F�x��$��y����u�^|&x����Jr��q�+,.��+2o˺��;�WyD�q����}�ǥ-�}�V꛽۬^khk�?���)�2W���'߷������5��$�sc����ګ�皾N➪�}{:� ��3{��k�_E�[ګ�V���S3Ԥ֚��͝�}b֎���|z}%nឿ�;/��Z��҅���Jٝ}�aҮ������wog϶g����{A~�<����m����k�]�P��s�]��"�f��c�LQz�ww���x��
���Y�;{k1��:����ōkE_A]Ҽ�~BG��7YػJ�ꮰa���5���x��|&g��5��qӻW��`u�f�ykA>4l~�FPf�l��>�;U���#��Q�W�!�V'zӼx�� R��w�!�=BP�Z�w÷a,�wxt�o9��[��^�����3$A`uՂq»�u'���u6Wfmw��}�Sz_��}��;��{!����M�Q�	�#������\��cQ�[�E	��3s�$�'Զ�q%�_[|p;s|#��6�	��&ea�묣��W�{�Aѩ����3�{�Qbֳ��7���|���'h����ޘo4�e�Y����J��G�(D��R��E�|���1�iY�Y�wxVnB�K˺
�����~��3N�WMeug�o��fU=:�쬛8�o�])�D�hu�q=]��<�s�Mu�v�֊��]�E�Ԯ��0��C�/r�I��hsX	�_��YuO+2�*���X$�jn:�S��im�w�>̷�;A�;#�0�Gp�(s�;1O��S�>�v^�|;'E��v�%'G�K���,P���R�ƤGtu�xr�~��;�*���^����o��0v�.�o������,��q`i�ʹ�IJ�S�M�vN,��g�q��JŤɺ=[N6�|����e_�{��>6�U㞹$��ڝ�u�7�D&��Ρ}1�G�]�]s~�I�=�i�Ž2��G5����q�YF`�#^�����������y���wˣj���s�}UU��f�_�]���Tv���R�7_l]�w�~����Pد��M�O)�݋��,�5Ӛ����IR�rs��w��ηp�9e��$�4	�q���r��̨���Y���s�s?v����Y=m���L���֊E�:��'�x?t�#b���7�8��;�偭:�.>[޾^l+�Uy�JՊ1K{!y�����o��}�vH�k|D]}gkܘW�Ybs:���W~�B���r{���l�9�PG݊�o�l^�F+�~�u��d���2���+/�.��e��ȯ5sc��>7���6�x��kd�jɰ�o)��*>����c
�x{8orKO������1?ww3�g�����C���C�3%�f�����,��H�{ɴ��k�n���+z��'�Tu'�����Zx����jsz�z���a[Euιm�X�U����� 6��g���8���F;A<j���PX'��y�/��6�����{�ś�{U��S|�k^c�^ѽ���
[��y�\mJ�Abd�T�$��z��8�)��l)hT��4��W���(�x,u?_tͪ�=��g6m����� ��*���Y���Sza��׼�g��ikj���S��x|�4=݋�Vpl����c%�S�)�k�~õNq�C]�<O|���o=�y����x�G��ز��|�d�8��{$���:R��X�yg�&�����t[��L>U��z�݌�����Υ�WM~\��4n����=/��{(%�GZ��Q�V�z��G��Z�=;3ճ�3S��O�Y�βM�U���`�|�w��=�k�Z����'��D���R���c���MY����٥8����2M��+�We�Ֆ�v!�tx+d�Ԛ�IA��J�5%P���Լ���x�����]e1O &vn V)olj����+3�Y�g��KˈI@���<:��O`;归v}2s8f����өv��{]ۦ3촊��X�N�l��2�s��p�Q���'o#���'�ś�E!l�م0�Ĵ5�õu�Z/���[�ܸX�����[�bw���y�.��y�]�Ν����p���Lŉ��Ԩ�wz��ե�6\��|>��!�*Jfu��{���=�'�zOW����V_�Tv�>Tienb��f���Γذ8�v����F�E�ڋ�U�p,v����6��@\
�T�^g�-gL*V�YS��D�t�%�{'hs����3��Y��g-���F�?��R�}O�r-kG[�AI�SeyX����1�^�?�^BS����Fc�j�����֧=��Z��ᆟM(�ӂV�>\V�{F �:�u���(#��+e幷��Cp���y��y-WZ��9�u�{�5�F+��8���xd�젮~9w�U�W#z��ڛ^��U�nke%;�?�g�`��8�������})}��wNVU��-���J@������f���g�=<�Ϡ�m�`�s�E�s�|r�s|���F���BNt�c��TY�O|]ͥ&��οr5�Y�� {n�ya�Y����Xg��a-�&��d�h���ڃZ7�u�ź���gVdy�v�Y&fq\�^��΋��x-�7q��T�1�û�o!g3a�Q�'G3�{��a<Yq���uۨ�f5Y�!�=��*�H��8`��嘆k:�����^�����b����R��iB�ذ#�����LJ�W�;!���O��.��r�H�ϫ|6�����Uk��*��h4��c���B�H�۵9����y�wx9�5i�;�OQ��H�B�mw�S�rr�*��o5�aw�W�� ߤO�ɴ��.ҰgUu�J��k&�u#��	�<���>;�dŘ�{�oI��Q�	�'y��onb�dܝܺ���N��i��Vϊ������ao� ����g���򀲛�aq2#����Moz��W�,�i)X)E�kY�#�\K��.7y��W!�<��&אqos�>�s�Go��ݱ�R���Qٹ����&���^��n���op^m�TM�~��iڻ�n��md^LQw��ޫ�žNx3��b��z��rZhu�q1�ӵ�+�g��F�\��GR:0l����U�j���%|�]�H)b7��]o}������E�I�͸�9Y�(��Q�t@�_�*�f��9C0<�p��[�qe�������=��duM&��4�|Nq2Ҵ!gun�_L}�W{N$�]V~j��V�[����������[&��R�����|��E��G+$�g��,9��'\�~��o�s��0�T�Q��{���n�����̼`w�A���{��|��ǜ��Ol����V�nrK9��9��i����^�7��LŚi�&V{�����v��Ov�r_�eY�ڴ�j��l�v�}�kg����J�J>Ʒș��eM�W?S���h��y���j�AN`{�Q7>��x+G�x�~��Ék�枞D�2T��΋�������u��������¯�=U�S_{_d���%&hV�kb�W�Ӵ��n�5gڴ�d��wq����k^/{�u�)��n�Z�]q��J�jN�<���:�'��_L�|�^a;Xz�]<2�X;/[����}:���,�|��^�m�]3�מS/ضԆS�����j&i��{��4�{��K=�;�ǵ�Wm!�$"�P3���s���l�����J��^:ٮ�R�6-ڨ�_�59��y���aV�T��Ue�2�U�p��7-�܏���^̙�[�_T�A�����#]�- {J��ntY��S�~�ox���7v\7q]4�'a�����+�osD��C[�t�����'���ܷ���������:_��>����9햎}���ܦ���/��7ѭ�5d�w&cc)�_r�!���!��W���"�5�bݼ��Z���\o�7�k�Ղl;�fKuM|����S����6�&�۸/�Â9}59��������a-
�
ШIz)Z1}�d)����h���qW�T�݂�_;/�z;��͞�ڗ�EPH==M�=�G�������� ��c�u�1�޲�o-M�O{�O8�Ȋ�{ރn��y)n ��|����N��'\�ϰ
�����q����nh�Bo
��R�\�x��/��W�>�^M`�	7:x�J�+�g·^}sv�-2���d�{<�5��p���t{͛����� T'�t���~��}���\$Oie�ֲ�mo���*�zx�g��ϡ����%- ��t�>��������+8�-��/1�Q�w�72S�7��7[�"U�<�1&��Eᬮx/-.��C�]u����P�{j�.7(l��77��u�m:�o#�g3SzN�z�9.u4�X;v�n�sC��a�JzV�������2�FhO��Ń4g?�!�V����s�v��׸[��ZŅ�U(��~}iRO�:_J�*�#�Y��܇�\+��*Ùr��#��l���;�g�3oEU�GǦv�Y�糟���f�.P��ݼ*_�y��Gc湎Va�.��-�^o�uMb=�/\s��z�洼�:����zq�!�~4����7�Ⱦ��z[xs���`���w�/�x
�;��19�'b�II���*W���������}F�t��V� ʗա���=�����^��@��e6���O��gt��s������v�����r2��W��l��`�خ�O-h�7��ITs�����+ra{QT}�PE�1_����[C�������=�Y��g�4���X_��3l�΍�+��W�W�'���(Q�;����x�P	a���j�碹leu}�,����,Z�Jy���me\s(�P��{JqIeۭ�g�%�K3���!�� ��x�/�\\ ���gv��&�gJ����Sc�@/{.��}��1��qR0�x>ÒN�>���v_u�|�P�+6�9���n�^��-�5��tX�*Ʈ	C5h0�Y�d�J�`k�����Gt�|�=��^��z��J�X�&Vk-��ۈ]��wOVw�0KsU��ۼ��io>���t����Ev���ٗG5;�]��9Uϴ�-}-tU2��'d�7vP�A�!�*��pL�9���٢�̠z�ػUp�mg$wdzf��;:/Q�aД���������i]B7E�d�(��V%ur;�7}\��H[ٍ�d�Y.��.�9���@��e��c�K��W%���*�)m1hn�:�yw�'f�NLf��N���׃�ŹL#r^6��T�貜Z�Q�݂��]���P���^�>Y��9u�1Waݢ4�����\SK����=�5�����̡y��Mr+���u�u���d�Qz�M�1��F�����{	���el�A��c# ����SD�se;�!��R�IT�����*�&�[�Z����bw �&5<�cVw�nGty�Z;�8�#Y]f�P݊����Σ`ӷw�����"iK�����҃�V�vw:���iw%;s���������hዣc }0Ʀ+�r�b�gZmEP�� � ��S૦6�堑��K�fq�"uՋD%}��1-��(ki��Y��q�T��\�ݺS��1Z3U΍pw�&�rY�fp�w��VR%���q}e��[,sPYo+o�'-�8�hS���i�>�0]���_��]q��R���J���G�-����Oh��j��S*V������IyR�Ö7�v��Y�;�+x���>n�q�]��	�ar�]��0��Ӣ�[df�<ʕWn�z��AkR�e�T��]���;s��'y���/���\bM�U�*���jNǕ�91�e�lf���W�������g�1|Ee�ʰ��V�����r�
�xA��1˓:;��c&4�?^W.�̊��Z,Si�;)�'��;�r��\;�������ƨ0�B�����x�xoA4��ua�bv��eb�uf����7����ehLz�_qg�y���Wv븾�-�)͎��c��k��)N�>z�K�Ek{�u�Q�%�k%c�t����
�.�A�5�L?�Z&���j�r� N͗O1��l��x'&�bV�Cp�=�t�S o�`��Y!�_��(es�[�������M���e-��� �\�ެ|���(��
8����ԕmA�X�bu`�3Y��<�σ�O�m�FU��b�<	U�:�Z\2�ٻ���{�
��λ��uDKT�QV�֒�%��j��Z ��)JJi(���Z�h��T�-KMV��F�P��҅P�E%���)]:��
V��*�*b��Jt����6Ԕ�!K�Q%:�14%TD;`�h"i��h�(GH�ti�i���CATR�M��BR[�tR�P4	BQ@Ҕ%�BD�Ў��EE!Gr�]�
B���E4�--<��HDҕTŧ%R�_iB��|Hu�'%o�X}�`3`o�l¹�Wh���2�l�u�����'���7X���BM�V��F��;��ůd��bi�������G$�������'Z1���o%�ދ��E�ݞՇ�4�U�T�M�Wm__r���`��xG��t�)o*?j�K�f�]���쵻�c�r��ݞ��;��A/�;�=�W�h�,�g�OT�gܞ��mh��n��_��V���js /g��+����Ѹ��y�d��I��V�c�n�=_:Q[���e��[~��t�h*&-ļ%���rԃ�����iyMY���R�p��,���U��M����iݮ���))Xڒ�&9ŭ�s�Z{2RT�>՗n�/��`+�z�8�2}���y7�=צWr5^�/LS��洼Ϊ�)RLv�י&N��
B��j���n���M�Q��=m=��O��d�ډ�^�h�����M\{T��S�[^�{�o� ���uz��ϑ�os¼W�޺ՙ|��&��Q��w�տ�y�'�*�iۥ���cT�YYW�$�v$��R��0<>x���X�{��5o�b�]im�Ź���d�U+3y7V]a���xY�7N���KQǈ�2-;wc[�c�
�R�B�e��z�mv�G��i��[�$��>�'d^�Tr�����ϖ�^��G%į'����DwmM����o�l
�{�����i�_r�����q{��ʖ��%��n���}�Β�b{�`TݬC�3%���+��WQ*+I�"�3��ԱtW�~�H�*�6��I�XV�!Q�:8�K��a0�Q5V��ъ�B��Z[z�C�3�/�T�����\O* �v�쎬U�iX�����b�g�ްWn�\�y�}���#�O`v�<q-~�|�����q݊��yf���Y��Fny%�����֞5��y�{�4!�(����B�v�Rۊi���W���y��j�ռ7�QPuy��O��k>����n�b¿�����}�)Z�ߕ��Xq�a[����}�D�NH���!y�O;�%h��y�������v9�]�����Wb�\���$v�n_7�hz��ee���g8�9��KOt��9����S"E���U��ұ��ͣ+9v�:i�F��&��|�A���x�T-��\��;�u�ԑc�5�5���LE��=}r>"Ӈ�(�m5��)��3%vm Ѯ���q�)��Wܿ[��|"�լXZ�#�ӾZ�����V��~5��%��0o��
���/�(���g݌68ƅl��jN���5p�7��\긼��S��`�L�ꮲؤ����v0^�m]&�u��� �'c"I<�<��fs�d�3C��b�v��>���Or��=��7'N�X��{�<��sv�5MO��<z����e��`��-�����tڏw�,���w����5d�w>����M}�EzOi]��`�Na�Q������2~�}�.7�Szv�;�l>�&d��ˠ!J�Ю��̭�}~�?CA=�8.t�}I��n6�H�z��d�C[jw�7S���J�JFϫ�qF��N}�ܢ��gͩx��{V����R�ݽ��=��l�íҕ�E̮��k6�yb���~�/���^��u����1XI��n�����ss�xG:N�=��VY]�'	C�=�z�NU4?4L^	$ O�f`�����X�9z�����(�t��r>�u�v��w�*�
���v������i���U���C��E�����mM�?��}O�I닻v���BJ1X��dLo���B��%�-���ݭ�Z�`~n��s��y���`O<����}����s>��)w�zmZ]qcܦfW��lNG�7l�3]w���^N����A��X{��xp�����!nb�0ӹ�������u�aoo9Z1�ej����+3�C�Ml�����������Y��'���~�ʷ){��,-j�E%13b��V
�?C��_�cK�5�Q��qm�6�T�et.��(��y e�fcr�ژ�������b��j���Ϊ�w�揵��=$�}p+�'�������X���g�b=�8�q����֗��]Lg�WC�{�w��,���nd0�}}0�RN�U�PqΧ���|�W��x�u�r�<��,!�wjK�m�������kGA�=n9��|O#"�57ڨ{ϋ�p�3�����ie��F�3��*jв��k},MjcXw�eg�<0'��C�n�y��C�oD3*��Z]�lV[0+]�P���S�N���W����DsV��=��E�[�r����:Lvu�"��cB�����M�NhG��U�����Zhf��i��}�*�*>��Omv-���v��]Z=��K�?���mȴ����,Ё��`�دGnǻNPn6G^kF�Jm�~םU�!����;ksFK�n��
�����}���>�}<S�g���/s�KQ<����BKB��c�'����uPۘ=�g�,k�y��)iTY/���z��x��bR�}"��ܣ�H:x
~:a�	�]y�K��^���f�ˊ��:�C9��]{�SY���^=�^|��G����7oG��s�l��]�窬���mdKf΋yN�^D�լ;~��0��"g{�����w-Wɗ｢�	��]�=�zĻ��|8���한ח��z�\擕�n�׸�)���{����J���&��{�jR��K	9��ۜ���q���J�����^��{�!��5ig�!�P9����ҋ�H.�>�=����4�k���rx>���3�%s�Ͳ��+��}0G��I@��fMv�;w�.�8(��y�nVS�L">4��P䞞sC(��+�L'e�8릞A�yWrtxf$��}W�,s��`��#Ӑ��j۾3z�y)�Dx�Ғ+d�ԕ-=��s�֭=�%%�&�'N��zi���}��iH_OM���և����s�b�O���K���׷Ɨ�W7j�B����e.����n��b^��޿(YP�,:�UwuU�^���3\�N��`��~[^�fo�;s|#����ǖ�W`���=�^����y'��S��ܯ����Ӌz�� ���;�{����Ŷ�I�#�s]Eq�{2e9O��U���t;�����}U��u�[Ӯ��Ͷ��¼]�{¹!��U)�;H��7�V8<G3&y�z���O�&��y.�
�T��=)�C�a�6g��^L�p�F־�7z���|[W������٘�-G*:�l�?G;k�N�0V��_�rz����(�ϩz�3�|-M���9M��F�����ǧ�����A�}��M9%��F=1��{��pu�+��gYչ���C�u����v�\ŪK ������|Bɗ/���}���`���<�=��g��W'T��u*6+z��A���k.�>+�z;�|����]�C=B�e�X��6�G�&^k0oK�I~�f|�ʝo>��Z3k<����s������O�B�������9�9��ܗ�vb�}�t�u��9<��v��^õ�8nx���|��b��3��]�r��T*�u�{�S��w��K�L~�����^Ws:�;�͊/��%�j�=�l����δ��&���z`yէ�2�|=����{�U�kլZ֫�t�=@<]�j~ۣ�d�ܥ�s���u����X;oº��ղVjNߧ�Wʚ^��g�-#��S3S�{�>KOg��]��E<b�������>��5���;�����.�ۉ\��{zŎ��E}oTI�W�C�|�7�Q_fi0��w1'f��}$�lG��v	����=^�o�T�J��~��;Sy+;'xz�|�'�^|%ŭ�}�{���]��W���}��x^���S��q��U�E
��)���uR�b�v�r�(�ۃjƃ�@y���6�3r23S=�r���W_r�#W|,��R���f��^m������p�:|��XԾtd������W)�Z`��^_pcv�[v�ˤ�l�)Y�hn\�;X�'���2j�*z�N�����|�.���b{�����̗B�{l{h�QX��"�}�(�ɯ��o�&�*�q)R*���W[����[�ͼ�0壂Oi�0���y]G��^[�����s�I�v�&N���.߶�o$���U��']�\�]�/���ħ9��)�>",�'���C� ��盔s� ��<jӥ
���"F��"�Õ���~�>��������<���s��={�/Ub�Cb�=�K5OQ��>v��}S��WϦ��?'�m�ǻ<�?S�*��׎.�:r�X�f��,��oŔ�I��b�f��yY_Gի�ӳ<�r�>��S���b���~�t��)3��'V�|g��M<�^�r���b�Z�R�Jyu{�>�U)��sؗF�9MQ��P�XpB�؉�@�y�T�n��X�t7���ϡ��hZM+��c7U��f�c��2�h!*�GC]�n����׃��j{�uyN�����CS��F��X���HW6j	�JȝO�7u��͸��k��	V�X�9o(h�a
�v�>��\7:[�̻���ַ<�t���J�jJfn�+���5�ކ��>�ڢu�u�s�������Q^.���eOM��+W_A]%`��q��u?.kK�ꮲ�Y�n7�]�s7�C��Uٳ�� �&,�0ZXs���EQ��5 �hq��U��A=�^4�nm�s<�ي�
!#{��n����5��ֻo�Y�n��̃���*=����I}�|X?S}AE�kEpĕ=��jznXi�r���mޏU���oˀ�t���s�|�L5tVU��뤛{/1J}��M��ͩSv�94g��[�h�H�� �۸�֊vm��r/&���8�����jr*�=*�]������W	��8O6y�B=�{�CsR�	:�"�ϣr�	 ��~�Zu�/I�p #��m�竈�p�����nG׼�5�~ne��%��� �|��G�y��ߞ/A6{`��V�2
���s�%�7��K	�ާ�b�^���c�Ѥ��[r]o�+i(r�f�zb����'�grX�J.c�o&�8�Ӷq�A=���#�0�<���nP*1Ck&�s�J��\�9[\����g�[�Jnr[7��s�~/O���<�^�R3��c('���y4����e�U��iv���V���S�=ئ�e��$�g^V����j̩�s{͛�x�:V�머����!��'���wX�dΓmv�g�#K���rV�3��q�ভ�;�J���+��n(�*쨴��zƭC�O����ll��&��	�qkw�� �}rK�˾^�\sVU��^l-�z�x,��؃~և����qxLS�~[��du�=KW�/@��9>ͪvK��)gfK~���]&Ψ��	�$��OQS6�d���l\��9W``�ED�6�/a�>���v�Ӥ��5�\�Z�v���@����'���?�S)�X)��-ƾ�צ�<���y wV���d����.p{P���w�3N�_f��C�w`�����E�/S�Ya�sJ���('�¡j��D��/c��Xݧ��X�:TxX��ĸ!�R�۲�]�a@FE�W�[����w[.ƂC�����"�͖X�,c�MV5����+���n�&.bv�M�B��,��u4�L=�2�)hc[������<�.�Η�ٍ�N���-fT�������Wb�[d$_2>���kW+ܨ�.%�>�f`��}˸gG�2[��J-��l}��,�w���W`��e����i�-sW1��̃��&m&�h�v;s^�u���T�^�}�f��X99>t�Qխl���x�\h���3~Q�h&.S��E5�J�/�I��r�D�*+��N8qY6�c��j��r��thZ���;E�\�v�.;�e�Zia+y�-�ye�s�6�K��5,$��F,�}R�i#�4��l��*�\�afw:��˵��DGuG�[���I��"�qK��!��M��8�#��+�T�Sfm��s���W����|vT��A�&�j�\����[�vP�h^ٚ2�Ca�s&q��0�p�mc�0Rޱ���5�[Y[]��kN$�䓱=P�r�����9�1�ŏ�	��Q�N:�\�cU�aZ��C���W��S��l#)V��Q�f�m�3��6ڗMt�`���\u:YO1�d�o>����58���聕���]���~3�Ռ9�]-��8%p�B�Op_	-A.er�6E�1t��gN�f[R��`��p�Ȕr(RO�������h�k��{�)e"��H���&WZ}�;S3����wm��6�x�Cʂhe�E�l���QQR�����Uؕ�9�eV���R��P��:�Mtv�ϡ�4��y;H�d���x������1�K�vJ��JpD��vt�L��R��3 �V�T΀��Lč\ت\-���Y}%�Wg5|�Y�8�qF7{x}��;+miU�'J�F��]6��*깗�t�a޻�n�gWvRG&M�:F�Vޙ jܪ{]�{��v-)L���#�z�9��%f*�ؗl,��r�㻚�9K/";3qgM�3WOl��".]�����'+��i��`�:	�F$c�&t����)ǣn邸7�\2�\���:�,�m^Ed.3hTė,#^�Ю�N�ͦxֶ����Z�0Tf�Qה�z�����j�4�8w�z&�s�45V
�Xju>wY�`5ϏR������d�Q����75����W.D���&�`	��]v%�\\�O�|wU\9�Pkem�LJ��kE�H��B���I�Mb�&����8
�����Qn�b&I����,�K�C9U�gdfT�(�r�D�Z�i�(�.��j�����޼���YF�H�`���>�a���`��)�:rj��.7֤ a\]q2����+5��[WGV\���T�T<ʝ�k]!Ί
�
��R�)� �
)�d(O֩���
ZSZ
G��)f]�(
�i9QN���iJ4j�:JB$�&�F���U4�#Ei��ti�DD�2�t�[jZkBh�шJR�� ��u�J�(��bf
�F�*��(iNA����[�1�6ãN�t������Jv���jуl��T�X��
4Б��Ѵ��*t�ZH��M@h�)Ӫ�l[bB�l���*���
��*��@B���@Z��W��e޺׶b#�D�[0A-qҮ�l7��p�Ij���in�w��8$-���2�z����n�����6o��^i��B����<���/q�Sz=7k��&b����s�ɒ�R�_WuU�Z����A����\]٢�WXKB���F㧉�V ���M��>�}���ܨs��-����}͙"����R�
�w ���Y�a��$��\*oO��}�������l��<��hRb[B�y��׭z�ހS��t�JWmyv}[�7s���s����W���K��!n�yun�/|�	sn^�vb�}��+��R]�|���<o�-�^.JOf����o՞�C��Do(�ޅ�r�o�P���~)ς�O������=&8(��� ���U�h�ի����������m�ȴ�5o��E9Yi�ʑ{)����Ⱦ��Q[���լ-j��|�x<O�.���֝������y��Sۊ���,/�G��h���(b�J������qQ�u�6�ߪ!��𵣚V����r�[|�`!��+1��f�;�@y���/y\ħ}o<[����L�_{�����͠^�@ȲO;��g��n�{�77�l�x.��P���S.T���5�l�e#���%@��V�.�	�8S�Y���g?|�� �,��=�:�����,���|5�}�L����g����Ә�v9�'����^�`>���*&i��{E��*����3�K�no4��<yy�N���@�}�~^�}��9�:����w�񸚘Rw����AZ� K$��;�>�oA������;�o����޾�����_ݰ�i�X)��I���cn���q��/R[7����o���*��Ƴ=�q�`?��� �ׂ�M	�5���o¤��s(1iʝ����ʛDe�F�����P0�7=����_gqː�-9�����E5�޹�nTD�-��vZ�[�Z��[k�o�D��.�n.��&�>�G��<9��A��M�=�d_e|�c��U����o��>��G}�&H��zv�<�����K�5��$���O�t����K�s�n�e�kx�6e�ݔ�!��R̢�!R7+�Υ3��]�`�T/Et��XN�6:2��9q�����4iv1�_q������ײ䉇�ڸq�4�pڤ4��ep�Xx��E��i^�u�RWOX�;]��Τ6��u��b7m�#H��f�Z�n�T���������>�s�=3P}G�,=�lܝ�>�m�-D��S�{�.�f}~����b�b�wsk�>hV�̭C�#���7�}^�I����gY+�ƽ9VT;�(�I�U��ߓY�,��~y���ҿ>�H�S�Z{J[��y`�k;����z���ya���u��dj�W5'l��L]ޏ^Z{uW_�K��0�U�|!o��\�T��oP{��5}%g��|qx\s�՟5��Ϊ��9��SU{˻&��w�
z�s��,�gS������'c�w�~��R0�M�/�M�WL���:�%WQ�̶��7��j*�y�����R�bj����}t-,���O��l�z����4���W��^~�؞&�B�/5s8�\�w˶ �u`�3���v�X�Dw;���j�*��+��ج��x��p!��Fh��fbgưm��6�lW�q��]\��춘�R�j���Ze
�Gp�԰px�ݵ�M=�]3��;r�,�iP]�s�iF�'�GOg,�����Q���BR�ܺG6d�Ȟ��h�f�Ն��r\U��姮�I���ɹSzM7k�3�y/>f�-+v>�ޙ�9B��m"e,�{�c⧭-���=ݨ�%�XV���x_�\r�I[�n
tĕ"�_�y�\edk����T�JT�\nQRA���,t�MUx='Oy=; ��U�{l܈���JO����72��K� <V�n�=}�`:ͥ����^�B�.+>t�g�ߦ��jnm��^������zs�]�~���ѫ9��o1�z-P��.������[��sNߣ�y=���׫�*�׀ntz>S+�l�w�<J���u5����}���]����~�~X��sE�TZأ%�NgE��K�{���s�+wd������އ��+:A�9�OVL���kk��&��Ls�-��9�>է���R_ޣC�n܃;7��yIB�tW`��v0߾�����<�{�^�vUb��zx|Y8wB���tuF����K�A��	��f��L��kp�p&�dH�\T]�n��v��	�f��Ğ�O�ZO��ڟ���D���`u�˓+��}�3�_�2Q�Mu���NV�$��:�ë�XƁ��Me?���5������tx��K�ꮰ[�����-�cx�]&Ψ���}'�{�˝���[K܆R��R��TO>���^�0o��KR���W�f�׾�o;{`j��jQ�s$O_ܯ����`�շ�ݣ�t��5��Tk{���(-�Y�*{8=�M�s���[�j4鵘�=���B\s7��oGv�չ F'�r��o¦�z*n�9+s��>#�c�[n��mzɷ��K����T@-+3���Q�U�mG�R*�d��>i����|�9�?i2:)M޿��ymm���l��(�H4�zѣY���S�*U��{S�ת�k���5�K'`��s���g�~�X{y�5^�r�̇#�G��|O�����t\G'@:�큥�অk��k��� �v�9>qN�������xS�E?i�����4�%�K�~�\�V�Z�F�]1[�o}c����`�X�'Z�+���Bs�f����3n7�m_����Y]�<�e�:M������zT&��bT��Eu(�*��]o��N������s�QS�Jw�ޡ�������:�+�[y�J5�N����5Ky�טN��6S}�a�n���]]�Æs5�gf�{$��y���qƭ���~:�>�6S7�}p�2�����k)�TNw�א�� x~I3?��Z����U^���lqю*}G �<O�%׏�<킝�3�N�n�]����gCe�N.y�����>/�'0W��P�Æ� ���Dv+�GN�@���Zӊ�����︪����x+��L^vT鿬�{��3ƌ�B�u\v���d�c��쌊�N4Mw�R�-�W�Z�)�Wއw���ҽ|-vT���$�<��E|onT	D���{�3UWZ��l���8�;���)��;��}MS�Y|��*��$�D�`>�U��v����Z���z:��ٗ:?C�ԣ��hR�O��Iei���3�:�o���_��B��V��,�giH��E@~��;��=/�p:pN��wM�C�\*�;�ܵ���a����uT�%����^�?%��3Uy�6_����
Akd��y���:P�Z-R��cs��t���@0�A�F����ꭗ����V�x�u	�`�鶴/#��ۑ�������c�or�������'c��Uۣ�E����
�k�7� }<K�g,�759sur<����(,f�HVu��8W1K��v�:�u7g>Ƴmwe&��w��º�o ���Uuлc��`��� ��9�vɗR�̴rv�oS��^�c��_����+�7��o��iL���BG����FB���ێf��ݤ<}��tn������7ۮ�:`~�k�T+�Dt�tS>��ρ[8(�\e2}ܧr��]��Sgh�=��ʇ|��M��ɓi�_������Q����҆�qޕ���r���9���e��X��81���%�F����N�{�)Ѹ�����w�o���ύ��x]��k**j��D�{t�'��{c��Χ�ฎ�ZN��G������}]r���bu,Ӿ!j�4��fm$:���n�S�l�9��P}�k��٥X{�������S���߽+�nz�Q_��m=�M󟷃�L�l2[��h?����k���u��Å��\ ��]��Ezih�'϶���q;խ�u1粟N�|��\gNIۋ�O��^4gj:��U��b������R�ܵr�ig��X�L��S̽wP���7}�Y�/����$�L�i��ED�Pߖ=C=�����%t����������L�Y^<��{����|Ug;�Q�}Ի�V�O}z��~�U)�����B�@Ր^sXk&'�-#���y]�f��E��I%|����oa�v���-[W�6������8���u�}y�g#����#���(��Hb�4론Y�J���. VH�1J�.4���귂o:܄	�;լ��΁ �x\T�p�ۺ�7]�bo�n�������A�MT<�E�z�N:U�+������'�Q�㤗FP�=Ċ.R�멉r����μd�;��J�|
���g��{HN��>��,� og�f	)V����L.=_\Võӕ�z��#7�x�-V�nc�ଦ���֍&��tF[��)T��� �h�"~��A�i~���C _�K���*os��Ǵ��#Q��'i9�������8uV�"IC:�q����Р��}^~J�V)�N������*2�.�&ӗĳ�.|�~�*���"��j˺�o��Y����l��
��a\he)�5yԴ�w:!�7�tb��f��r�k�U���d��C��N֕a���a�\3��Lv؞��x=j���m!���=	;�S��gR����dd��u�q��`�{�Rl�z�zal���0�\�/���
=��b�E>�*���= o_H��ۙ����#M�� ����?B�-1�'��}�C{^5��%a>&nR=��_�}1�E�]X��MX�]
���wOd���u�놥\8��gP��]MCepAWz�k��Ӳ{gk�����-�DM���q[�1h\�.����N�t����{Sk�U F��	J���1W�}J�����|b)oV�J$Y�^���z=��������׶ǥU<'��jr9�A��楚�X� �fy�����'t��\��|WbΩ���N�}�.v>�~�SI�N|�u��ɫ��u{O������e�]����-������\|&Xˈ�tp\���%�1[�W2��L�u��;�b�ii�v ��n�q��y׶�K���pg���gKS/����R��Hg���p' �^\��D{;L�[�|�;^F/�*Y�:I�a3��!qS=��ۺb��/X�聭�;�{*+8LK���΃;�8q׮�{p����VW��(�#���0�I}P��lw��Y�쳗��ȼ9�|x����K����Д��q�<ꑉ�0��*�Hzk�(	�%LͲ+�{"߹	�5z��+���	U�G�R}q6��q�S���NF���e��F�L��@x��h�^]o�}�r�x0Τ�=����\V���.��2�m���a7	������٠֑�=�̣�#�E�Y��I��G�K]4.)N��,+��de�����Yg�>d��*@Lz7����W�B4�k���޵����.�If���_^\��(aI�9}�嶅Ɂ�(��Fu�R������<���QN�������y�r�z�7�ۑ����}4��j5Ȯ�y�˄@�a��:ƛ*��Ɗ�4CV&�T���.v-񻼲�<��{��ߦ:OJ�'o�3	\	�+e����울Τ�R����L�۟����v{|��p�1z��	�H<Q9��Zn�E}+k0����fT,9��K<�;�	��`����Urmc�\'l.���\�����eQ�c�?�0��(�M��Y�v�}�V{��>���/�����宀to�LV������ɟ_�,5�� '�p�tV�7���)������:}�l�or��e��ⵕ���v���4���3���o?w��d�����>Q'�O��J�9��@^>�c�W?0q�c=����?O�s�;\]u.����|c�T��s.�������J�}ᔀ��|��V��	[�j�Ku#�ѱ�ُ�ܩ�\r��geN�����3�
��q��mP	F̆(��;��_�C�o[זs�/wo�Z�%8���}�w|�J��]鑻s��$s>3�
�(��7Q���뿑˭�����ǲ���ڨ�5����!���p�L�,a^��Ĥtw&PF�,1.g�R�Ѧ��N�;�� e�VJ̑=�D�U��N�m����n�0b�oq�GS^����{�K��϶�d�b�Z1#�m<��h��k����F@<jXo�^荖`Y��|�����Z�̶لX��.D�[��Tv�+xNCwf�I_f]���!R�L��.SG-fb���iR�nQ>맲�^0wo
�7&V0�G�v��W3��<�H�o��癹�oU�2�
*��u������<��o#W]:�d�M��g.��5��c�S�nĽj�J����c�oxl��k�jR��]�y�c����c�*"Z�k8��(�J�^,�/�Y�`P�aՍ�o=jT�#�0+��2ΫT1Uɳ/-m$1>�]�SebN� SUf1X�51Y+�%�a,'V�4>�GȼE\��}��<AmI�v�n9Z`��	�6��S�n�������ΤIUu��c����\ΛY��x�
���J��B�5&$��5�y��ۛ��(QacV�j���
B�W%յ{v��o��cLؕ�}0��MK%\�B]�G��ᛆ��F���*��]�>��6;�G�fmx%iN�U����Ȗu���a�w6�[0��|�� 'Y��L�ht��c.������ظ�%�h�D�� /{:��Lob�ǆs�����Q���9���XhWV��(���R�E��9o
�q�]�uQٝۄծ�u`�GZ�O��6#�SXhq���&Q`M7t�БM����j5V[���W|H�C��~�+֗i�}K�u�I@�إ��릫'f��P�|�=.Р�f��6�h�zQ�#�Qj���O�o�;ͧ���h��;q�r�:�y�w٘��1l|���s��֧Wgq�5�4n�>�4�v�g�nX튘i� ���p=�����glz��RP��/{0�@:Uh��N���R�'��鮩:�晦���M`b�*�V���Y��`���/+�ξ����l2�����r]]����Ά-%�� �M}ݢ7�]��~֎=].��3��й�Pm+J*�fޱE@�ϴ늝>ݜA�<�WU����/{tQ�z�I;�I�II�h��$v�n�\n�ecVI[�p�~$V ���we������ʂ���Z���R�*X���˽�R��H�Ы�ɰ����._cҫX�3bY��	���{�pa�汤+=$�.C��E�oU��S�uo9J.��n��'��u^�n�opv/��������Ojՠ���ެ�@ݱ8�8H
���yZ�E[��nWVv�Z˟p���m�f�߻��m�::L�CV=}��ɛ[�"�&�����T��<�ƬW-���F1�9��^V�܁��V�΃eƍ ����P�*�89Ck��f�Ô�{;1�7��57ם�����Z�y��/目�"w>�άRQ��]4����!ٶ!�ډ����\���W߹����:����|��h)ŶH�TP���G-4�[j��4V�4��@i"�1��	4��i�����i��Z-�Cit�����F��P���mk`�Ө�i�E%�뛜S��+V�Q�w1��ƗZv�ք�4�f��9h9:F&�����C�H4:��t4j�l�]�:1�Cc(���'N��6����щ֌T;��M��PmF-h��4hD5����ք�ys�bj��	��&���Z�Z�5��cZ�#�䦨�Z�4�Q��CF �3�Jm���ith��H	$�h�Vu'�^��,;:r%�T�S�˨��*`)Z��dѬ���:[�;�6>���T��r�V��Z=|���s9;G�������u(�SB�+z|�K+N2�y�|]c.��H�#'��nU�/w���|��g�����q�z��>�n�U�w����\s\�;y���t'��#8S�{���<c�IF�A]A��)l�d����Jk]���MZ�/6��CG+���٢�T[�[�8��n'�ڸ�	G8��N�ζ����P��.�;���Yw[��o_�1�pR�J�>���`��&�˙�d$l�1+iѿ��9RϢ�4sӎez�m��Oe˅��h�o.�'�7\�t���x
WH��N�3)����}���c� L�s֮�+*sI�R{�����7ܶᦪ���R�2m7@k�2/6_�Mt�=&:���c���!�T5�>%a�Ȍ���z3ii�W��N�z��F����w�z_�
�p(�m�׋�g�g	ځ��X�KÂ�V���v�w��ǡ*{���]r�m~�W^bc�z�W��Y=�gｳ�P�D��c�	�0��OM�iV���x���t�L�J�a�6I7��+;���N#%�s�pF�8P�@$��rqs�)���3���͠K6'D�?ǘ��+��I�e�[J`�D�0�n�Dvs�v>�؋��#��k�&"�b�׺�	�Õ��v�A��;V�Ġi����3��?}��r<���+rѮ� �^B�vW�ڷYS'�b@{ܼC�ջ�i�\� 8]�d\D�nN;�����p�~��t�g�</*����Z��1�Z>6����8��c��W=x��;.���7�)�?G�����ǍH�����}��F`ڥ�N���u��{�}\����
���s��P�7�'V��`�<�����3��CΏ������)�:�ʋ��������^$ ���q=\/n�x�EwU���>��}��;�����\h���K�]^�q�2mزQh�'�@@�$R�]먗q��H�T��9=��'c��/4�Ԯ�]��[Tp����8m;w�If�D@���i7�<�{�j�G�w�=f^oz��)��������F�q�茷whU��J�� ]5���Z�n|^���g�s��Zs���.#�I�EAs�[8^Vi��.U�V�IB��q�aNT���uخR�Y��*�*{N��6[7��F\%���r��|\���W����$o�t�B�q���u���0q�T�>�?^!��`?	;Ӈ�	F���!k4+��p��C��h�W��s&�>��{\6���,����as"�(u��g���J��8Ȗ�픒U;2���'��Z�^ԝH�]��!��on�C��٪Hp��L���&!�e�|X�������uxTJ�F��N{^u-7��p�]ы杚7ˁ�|�6<���2�V�!�⋆��d��(��釷W��^j��͔1mU�	'w@� >�p����,�����:��';��ו ��'� zam���qN��r���޶4�a$�gӓӯ�L�Dd{o��S���T��k��[ʰ�e�����(�g��&o�P�+����!нޕׯ�'W��z���e���}���DJ�xO9cJ�wPw�F��}'�,8J�<W�*�*b�^G�5�ӊ�:�6j_�	P7����&y�O�\�{К���s��xo�8����W>b��#�?�eT	�qS�pY�A��J�0w�s,C�L�u�����\w�wu��/�y_�ᅾ������Y�=P�B�_�T^4�v��1��'	U[)ܿv,[O�חHv�����R�$�A�L��B�{���1K֗�B�(yu�H>�R�+&�{�ۘ�v����@=����++��%GI=Pf	/��W�{g��~)J�_�(�֘vkz�e���	�J��V�(%��	��삮����
Ұ����{�Ew����]���g}A�����P��́���N���ݤtS�����U�j,�w��[f��*��0A��^�W1�ƽx����j�#%:�r��޲�'��vu��uˮ&�����jw����uH��}�>%" ޜ�(^��U[3JoKίǀ�u�YVR}q6��q����'#��r1��5��AD��ZCA��f�[��\�ϯ˦ӎ&@逺�����+��-���T�#/6�9�s�Jn��� ��p�`�뻟G]�yF�S%�RB��m1ytкS��t��oYp�[z}e�0����7bY��^\�P������f��+�TMq�'`��w�
�tr(�ɫ�:�w�\�9��x�<�mv�{���8䩒������܃_t�v����~�+e��w���9_�S�xm<�ѤS��\��-/�����\�X�V��4���ח �K'��a�����o�;S۝���?x�)��z^�������;�>Z�E�K���Q��ϴ�x�{�ս�3x�W�v5�r��z�e��OI���L�n_\2��1���<�]�����:����:.�;���'���9�(x�|�Pt2p+��k�����@W�x��ǢUs�!�c=l&��o��辗r,��n��^���Sҷ�#[�$>!=c��Ι�~����{>b����m�����X<*�g.�}���^�!�����o5��͜�]�뼧ӟn�cf���N��͏������x�RwV��9�꽂at
��5\�ƭqO,�c0w+��~�B�
5L�� ١�巟�z�aХ@>���+�E?b>��<��	ֱ~�����h��C��}�p��ʝ7Y=��^5v�\S��m�-��nn�����Z�U�k�:9��vE��y�܇�A����c}�|zdn�Βt�_��G�u2�@�*�^7���j���.ʁ<s�T.���c���u	쨦�������T�A's��WVǗ�����{�`,�WS/��]L���U����ޟ>�����go�p��Au��[�~��̝������{��h����GO_�����eӞ�Kw���;\r5�ð��`)����o���˕�ݳ�� �ȃ )-�,�}>�å�Z:j�W��w^w�OEN`���գs��mc��6���\|��phTxZ$X��a����I��69!�����c�V.��#C�����-@s�ɶ�`��&�˙��	��1�� �I��N!����D���3�x�8j��֌�r�r_ɺ�_�� Ƅ���5�M��fS&<�YT���q��tzw��R�Y�`�	���=5,�B!m�P�t�%εe3h0�R��'�Sۭ�5�qL��0��@3%卬t^bʱ��c4;{�_Gz!wGo�4��4�z�#5J]]L��]r��-wґ�2��j�8;���Ooq������B��Q�Η����4�T�G�2\&�~�������Ai��na���z�������>
Oa��<�+�ͥ��_�'U�8�E��p's)w�Nx5x{��:uV�9�|n!�'��\�
�^j��ݔ���cЕ=�zo�0��~�;�⯴y�_��?�ߴ�CO�ٳU�w�t2���0�������� J�{T8�����O��q���%O\�sCt����L��\? �^CG���,����U��|=�ٻ}�+l�p:�Q��ȿ��srq�F>�|���y|.3�$���'�\���z�J��wgx��w��f��WU#p�zG���p�t�H�/?\&W��������9'EKP�q�,YN�����'zq�y̡�g��T�t����J�Nh.���7�<����z��{�WS^S��<j����.�2��^�j �0
���p���)��V&�k�4z!�t�Vp�4#�9�=��J����a���Uy�~���H�'��A�$R�멉j)/h��ջ뛲�|�:�v�p�3�9�Um�(ڗ�T�AO:��0r��҃3bk��XiJv?�}�}<��g�YW��h�br�sC=
���SȘ&���M��ժwl뗐��/��r֎zM��'݌���Bx�CW�ɖF��q[���+�*�{������g���ՙ����l��>;�+��N�C��,� od�`�ZM�����I2�ۘ�]��o1lˋ���QO�O���e>;�֍&���n�ЫS%MG�.H��t�������ݽ��`�;�}ơ�q���'iϴ�W��`7	��-�[5)�P�ٮ�+�%��`��>4�l���&{��\T�83�e3-�Q�u9<��%�As�K��W���)0_fW�����מI!Q���31�:lz\�4.)�a�Υ��;�����\sN�>
[qC�]�Q�3����n8��P�'�JD\*�i.>�V��������������|m�dٔ��vvӠ㓠�m�`N�s��*A��OW��n��u�z���s�;�~suٝ�x�mg��hq	_��%T���ռ�
�~y�8��Lx�+��~�{�x�tp�-�M.Y���Ǩ�S�'�e3�
�~%�5��wPv�{E��I��p��XQH)���r�<�Iگj/0����z����>%@����}&y�O�\�{��Wu��_�J�R�����,OVÖ,�1�?-��x-�r8����Y}���ʺ�ڶ+J�$���Y���_ZXj��鞕�F0Z9Փ�t�ץ�񢻀͹m������ܜk�M��*.�K��r���#�M�<7���w:v�8e���N��di���˺��u�+��s/�Oz~Q+����Ih�::�Q�%H};%�1[��\���3�����5���CT���c�����vT鿬�{���t�qS/�Ґ��2(�c�1�f��{���q�g[�5���u�����M��vT�vt>�3ԅ�S=��n�Y��o�����p����b67Ux8Z%���t���A�+��E��$�3
�}P�Wr�u�� ()���Zʏ<����'��=��T���9N��t�p�FZwl8Jϔ�7������B����ˎ�̙r�3ip���V{0�Ӿ��*q�Ӊ�ö�܌��գR5�B�OM�n�UO�p<�e�#
��Hj�3���qY���i�Mπ���i	��{��������>J����H�F̐��Q��fEON#qP���#/���̧��֭�}Z�vﵝ/��ș�C�Ed��y�7,�U��^#n,���
욼�A�8��M7�O������pq���ZJ�/��1�+� �T���D�|����ED����x�܊:-3qS�o-��ap��(_:o�	�e^�[����]U���<�&��Ь�&V�����^���
s��W�p>'I�GW��x��:�s�(�Zx�h���[!��ڙ�+%��5��at������lIP��ųc�8��^�t��1C���N�y�[�ө����~0��o=�<���k �:`a|����kːk��� �-=<�������y���5ة�狌��/�oJ�{����-t���o}b�ɟ�ġb���j�~�{��h<\O�\@���+��:�i8w6S7��Ҧ���'���wpt&����0�Ń^�f�s�����������,�����,�ճ�����ր��z����
Y�&��{iYtf���ˌ���k�����1�s8s���̳0�P%�B�5��ҠzR�͸v��я��>]�~|��V�U<��w\7O����;e��pf�A��WN����y�I;4��Ǧ��{�%���uP���cvE��nw!��i�pc:W����w:I�Ry��jQ����i�C2�g���Q��Q�����/t��!���>�E5Lo�e�^�|J~}���:���mi��y�3�H�Q��L�,u��;�U��\����,�8�g:u��Z�"�%+>s�|k�Z����&e1���h���Gz�3�n�Uķ|0z#�;\tɹ󺞔�^Um�8N*�c�uk���)$Vs�]A.S91KT�Gyq�7�+��-`mX�C��Q�X��Al'��[�Z:�/8g(��g�o
�.Mڋ�a��u�f����DΧ
�[����2	�71�L%��t7*_qM��.�M�;���d���3�{m�:�������^��t7��AKd��y����P녮�p����R�$�ϱ��<�=ս��zX��N�I�x�'ûw#%�"�:LO�<�h���������z\�qa����`�MZ��\3a�X�Q8�\�@!#�d���9�[�������@�T]�q�q��Fc9m9.u��L���`:�G�_)�n��6o���x��(�J�,�𨔫]JG(��{��?|���yJdɸM��P�\��1��rk����%Ø�<xn@��WS�pe-�+�+
�W��N�z��G�>�����g�q9^��y�@�=��i�7��#	xm��+��Y��k�~��Z������Η��L�}�wٵN'CT�}V'qׅ�_�|o
'2��:�a\W��4���p9+�U��6��_gYx o�m�D�w��9S�+"9Վ��׵���R=},�˃0�h��U�=X�FfrΜ�=�爉7�ご���ȸ�u��ϝ�c��j�w��_���;w,�QƮ�Dr��Qq���Q�Xq�2��Trr������aP�Ϋ�?{��_ ɞǗ�:��ҝ��WgJN�e�o�����:��ZsD�76s܎�Ȍ0��5���l=M���4�ǘ283+;Zٹ�h=RѡqH�2�j�ym��]�@8�F��`�o�Q
�3.��vʴ��-��Q��%�]/�_R9N�pnY2X��l��}�V�]ѫX�s�r��^�d1	ҧ�j�C.����m��2����ã��}�t4Xj��ti������u�vfY-��c��,��>�Z�Jl�ݔp�	��6�d�f�k��'�Xƀ&�'{e�e��c�9�8,5���-�����f��:��V�y��õ��u �)�7�!|�n�r�#e �3jV�ʓ�l`�uy��N��ݷݛ9�*e��zV⧩��U5��&9i��1�mU���a=��Q�O�[
��]���S3�
���h��=Qs͢������s9��Q�
�a�6�Z�X,��їR��-��KN�p����Zp�����S2��*��4�fn�wD�o:����]�a����듮��,:e�Z1*M^��O�7��n��|",�t�Y��ʦz{�]*��&C%��R�j	1�%Z}�oW_�n*�ۤr_,6�����wvU�M�eӳ{��4�?,՜H�3��9�]_>.-��E8��cO&�l��Ve�E^�n����x�z��9[҄�i��b��lI�x��T���681���q���~�U��V��t,�mG���\0�$���O��8A![r�w�.��E�J���K����z�q����U�-����F��٥��x�o�b����r�o��k�cDm����4z!�ڵ�<aG��&�k�<��6A�;��.�ܙ�p��j���Z�kh9�8�h���]�+*�.�t��|�q;f�wE,�n���*Ӡ�Åէ4]>�	��Ř�GHXƱ����M��P���b�2�Xh�)I��>m�qΥ� �T�"Yީ�&�S���/��繐���W�μ� �������)�<h��q&��d�g�zOd�o���� �ؕ<�S!W7�ۖ{�=8�0U�e��T�QT!VX��tA���qT�ݙ�|��-\�Dh���PӃ�=�|�<��_dF�cY�.�r��Գ9�úl[�������XS��'uҰ�鮘m�l�:kkQ�:�)uA1N��J�$z��42���^���e]�G6�v��NDHy��
:����y����2�I����u6k�1�KnN�*бs��+��gc�#/��1�)��]�iW1��+W�Y�
�)�
�9��\l�WY�{r�U�� w�@.��=o���7�|�^r]+�(�N���'Q�ľ͋�v7�m��m���])˚j����ʏS�t3��{��hev�-�J�u(�n�*NFW ���-\AM�q�ղ�e��
��ڛ��JR�t|r���f��fI}�5�bň�֜N��m��t��P���4�-h
gb�����E��N��ƴ1�����l�V�V�lESAc��qΗl�-p��63��S�O#�1����&5��5���(5l�3F��)�SS@hJ[d�����M(��1Plm:+U�j�h�A���f���6�rĜ6X��K���QQ��SMm��e��C�4�b�:qD��l����9��j���b��M(�&�%�s����TQ��h4j��i���u�d�E��QX�b���"���@
���Qy���\7���m)g��N�F�>�ãe�tei]EWm؎ʑ�#���o�|z �΀�wCD��vsgPX������X�R�������$|v\c2n�e�C��e{�|jE_�ׯ$�ߙ��JXVY��o����C��J'C�	��_L_Ѷ�J��N�/@�L�Y^)�GH�c�8���։��>�N���U	����g��0X�C �(I��R�J������lh�캚��_y�.�zs��EOv�|5���;6����Ë%GI<
��$Qr�O��Q/WW������fݼ�ތ��s5M[�#g:�%���}G_�+��N�C��,� o
 Jp�j3!���/.�;쭼�~9�&7��Z����p����Bu�I�����Ы�2T�q .����]�7��Y/ݑ����2әH�wO{�ơq��c5'iAs�[8^Vi���3QP�����K��f���΋छ!T�ٳ�D�)W
��Zpg�l�n#��K�ɴ��,���%֦�y_O�ע�u��݀��a"�nT���J�uxu�N{\gR�q���UQ��s7��yp�z'7�g���G�g?���TF˳$�qD�x�܁/�+��x=�Z����Hn�6�_Rq��\E}�M�<��_�x�[jϖ��QHiN��;i���N[�xf^�d�������-�2ٛ��.�۾�u��Snحnh����|����Y��$��r�;��q�F>R(����jX=y�Y|�1����&�%k��&�d�:�vHȮ��H�A�]ȸX�:�NX���,^��K'��酷��t�0����ׄ��~���n��5�Ƌ�=��cЕS��k��[ʰ�g��X깑xQ>�|'=��Zf\�<��u�Fu������IxO�al�V�"US�}ʘ֧9�A�~�
�ɽ�k:�\��e������<Q7e�s�n+�X@L�"ʁ�}Pک�e���Y��F�>s��*��Ugq�~��(U̠����	�u.�*C�Ӓ�����y�V>�ZZ�c���S��[uJ>���S�-s��}S�����(z��(\T�㴤"���~n�s�w(��u�,<P��7I�u<t^��*Q�������f��ROq��Ĩ�յ��u���}��uw]_�o�׃��KG=���O�VW���8!D���b{�~�U*��6�j�[�tgY�Gz�%����n+x}�CS�� ��<ꑗ��� ���^jǖ�{�2N{��z\D�B��o�R=vU��S��t︄|�aL�^U#�{�U;v���M�1彚ǻ�gD��:l�����������59?��{�V7X�� ���ܩ=�# ��}���,?S�!��w[�w*e�
�C�<��r�':��Q�aV��g'�=0�֧Nħ���|r�]�	����=���1�QL�s(ws��53ن�C;�y�<k��@Q w�	V�`�x{åq��\7�*v��D�m\\�i��&'��u���[��O�T?��Ѡ�(���$.��D�y�кS��K
����0�����=����͜y��h��C6�\�G�T+U_q�'n L�;�1_J�tn�욆���B�˕o�ۺ��B�mi��ŷ�t/��K�,p�,N�A���N�!i��5J�����yA����G��l�@jr�c�&��r��N�_����s��ѹ�:᪺�=w��@�$Z�#c�+k0�\���>ޕ�r��jN�ѿ�]1[���*70�%��^��xןd�?��:h�X�Á��^�2�륤��l�n#r���%M=1��ⵕ�]���:Q'�3)]�5�����p?���=�,~�8�S�8��'��m /\1�uh��1����{�;�m�>�����|(�+q���6heyoן�z�j��f� ��}��,���x��{;�^۵���S���L�ј\7��;�:h2wz��f]��d{����=�V�`
�K�K�']\�fѺZy
��]����4l��ļk�ӱ�b�R�cj����w��7�-��~��i�4����Ձ8m|I�'lC.��׃��{�}�]�IT{���mc�!m;�<Wsa{]j\��z sfE0�F�WP-J�]X�]�'gr�v�\��y�����owi���~�Я��ِ7D?��7;�?Rz�4���*F��N�D�ј)�r�����3�
�Σq�=Q�J���x}�C+=���5Lo�e�Z1�gG��>5=�b�"������I�,	�
�e)c��ER����>��YZ}�9�0=2wm��}1�__�Yu�U�p�d�`�j7��bOQ �����I�C�\*���u��\5zc�P�y>����u��'pr���0�=%� o���O>�{�+Ú�O<���P�㙷
�޹��hq��/6�܄�t����pۻwp��k�����13ζ��JL�3^��N����-9Ц3^.��V�nx��9�d�6� ��q(�3�H�X��n����ݼ.:vu��{)Q��}Y�pٽH�m�r�rm7\�L�ЍxR��~�����e�ݬ���q32�3>�4����
��[9F�:V��{p�UR{�)L�7	�\�`�~G���F�;�^8s��5
a���co�����=��Z�b��KMƫ���rw|b�ap�s����÷�v��X�ԚB���n��7���;6��qV�!�jF����uvܣӮ�kv%F;(:��ƭ�����B��`�]Re�ޗY38�3ֳ]�H�仯�n���wwZ]�a�;�G*ѵ�Ѵ�ٽF�N�˻��:�]dI;�.\�ݣ�����~�� ���@���]8Լ8:��9�(7V7�&1��l���m���cl��p���+8����ڳ����QUߝPY����탘�����z���`ێ��}x��*]x�T��Ȏuc��5�pʹ�~�d�Y�^4�	|��dϋ��a��Ә�Ԫ��A�|O{ᔀ������srq�F>������_Μ��:xKUqwV��`��z˲x'3� ��z"����ܸ��]2o䧙{��	��3(��4u��Y��7~��=K�ӒX��$�L��L�W2�b�mP�7�X^�p�+	<Μ���SוU��}��}��·&߀35��p�yY���V|P����R�NťV&:��8������庻�wV����Lf9�Bj��Sl����#���2���H�.R�]e�a�t��u瘷f�O8�^�"㩻�涚<�O��<��ӷp�=%�D@ޣ0�,�.K�Hީ�����y����1i,�G|����-}qV����|q9���RG���*�L�8�y�>Y�x�y�w��^U�u�Ӣ4����p�Á7�D�� 9����`�Ӥ;�ٓ��\#�!��Q�`C{:a]���p�=B���ȡ��	�j*�n��k����ag+Ur���A�4���\�'.���YxsH*��:]�sOQ���Þ�t��=$L���z_�ơq��q��I�G��il���;	��3=���NW{:��m�ǔi��P�RWH�G���W�JӃ=��L��1턺ܔ��Y��*wM�/,ݕ4שPYj{1���׀�(��s�	�q�c~�:��=��3�i��D>���=M���O��՝u�=9�^�����F������Tl�2MqD�x��.�l���(�Q%��Ӻw�@�ɜ�y��W�_�4���}��ȵ��������������d�@����c��oǐ�������j>��E���7���[J���-t���a��ߦ�<V�<�+W	�yK}�����(�Qh{K��Q�^��f��8}���m���UO	��ʘ֧>�uq��WKU,�~�F�}��p��x�I�P>>L��=8�g���ҠWݍ\?B��e���Y������L�Me����qX�m��0�K�#�	�A-��	T_����9(��b��R�{�f�U+=�VakJ����E.���'z�\FvT����(z�҄���ڠ��F�9 K�����5fV�(�`�ۜ��96o]�C�v��t�e�g#�{�����`�ɪ���*X�l���(��x�dk�9�e�rt�ݔn6�Y0�Ԟ��z��F��]CF�o� �[�ZSl#�&�U�/-x��qYr�W�g}����v�T7�v�!�(t�z��:�:
�q�ޙGbΒv�3	�3Ԅ�����M�ո��~ڏ?Yp��
�E���Q�ׇ=��F:��v���Y\���B:I��Ϻ��l�����[��\l���e��w��Q���T�~.9�jw����uH��;�װ�\	�$�� b�������#��VR}q6��q�8�iȄ�a�CwA��~���w'�L�U��y��f��Q΂4�}2��h7
g����\moW�*v��d�U����ݽ{��\�i;���;�f����I!v|6���<�h])�så�ٰl�7A{��)w������o����2W���
�V�&�ʓ�f�U� ����4E�s5~"�1��<�X��i�Lu�W!������S%��偏�\x
�;��Q;@�Z}k���~����ayi�����K�XdwV�e��{�m�Bj�M��@*N�_#4=�� ���DK�΋�ݺ5�|%������஺���/K�Ҵ����zw|}] 輩b�+�;��υ֚�zp��R���o�7��un�vp
��
T�=�$|)>�x/���Li��v�%w���̬�X�_.��x�E�!c�[ہ�:Ռَ�fЃ���I|a:�4�r�����o�{/�zZ�k%m5�BPJ�����,��B�W���e�g��՜:vh��dϮ�<j��8�z�ΩZNaL�V�7*i���l]�����{4c�z�������M�hϏ}>șc�a��ܟ5����Gm &�v*y�����]�#���\hsկ��u������w�c*�p�Ne��^����^��'�͕�T��2�gWḛ;\��;�"��?0r!�&{����7���;*t�Yd�\��~��q�ѹ�������⺩W�^��A���-�nuܠ�C����%z�Z�W~Y�j�T�d�K�O;K�.����ۗQĪ�tt���rY��=�MS��7��`�Iγw���]=	��U)�I�x]0�*e)c��Fժ�W��>�Iei4�Τ��c�5]c�_C����p��V2� �k��(	����Ҟ���g��p����M`Y�QGuＲ�:�/���㬏��w/�wv�/@��k��A���� s��E�Rd#�޼�[�[2�owW+���/6�܄�t�x�'ûwq�F�8���1�3��.1�Ұc��h!c�؎�za�.��DJ��oq��Ō��`5��/k���������z�R�w:�Vn�������az����?+wԑx��E�L?	5��{��mO�3��]�ݺ�;j�Z�Y+s�����,'��B����kg��(�;���P��.�	5hx�\K�s�ɿ�u�_���j˙�U�ە�N�����2�V�T�1)WQ��,zs*9��I��]nJnx�� ��=�QC ��)����l�.�������f�O�K��W�Jg(��{��?.�gȦL�����u��,��|8%t;FU�K����>�֑|���ͤ6�9�r{�FZ�b������N����ޡ^��ݻ��������n�Eixg�C'��FN%��m)�s��VK��f���o��ûX|�k}w��G*qR����?b��3o�x�6k��@��ݘ��aK[�/"�{g����-�z�5��sٶ�x���}*��>�t���46��oY�enZ?v~�x�.WN�:r=���.
u>��$�'cҀ�u�sι�8�Jjtn�V���9Wr�~p<��֎z 0[����*���3.z�@�T����sЮ����fUA5�7�~�]W`o��پ�����琿�:rN����$�<�΅$��϶�	���A�~�~�{�mQi���]6b�B/���[�Vt֭�?��v%��j�.繇GgK�'k�Ŭ;]d<8�O��W����d�ݨ��`���%rO^���9�ݺJ�K�ŝc� ����p�u�gV�RVś�����a*I���F��-��U���ʹj��NEW�Ow�NP=��w^�g�qq��;W|U{���e�� �|e0℞��t�N��n�Y9v�Ӻ�З��Ə.��c�Φ�6�&=%�t���,�C�G	�X��w�1�{���/e���O]s���;��KGT>���O	�N�Bc�Y�D�s���YpZ�I�>z�+c���Qq��D����L>=����:}����ϓ�M��#U!Y�;����π�T܋��<���7f� �5Z�+K���B㋌�o�;H���4�C���]�A1S�'�>���"��?}_��\ԉ��?ܡ�A�����Ӄ<6S8��y-�&���n�j_���V��t��ȕ�
�)�H��; ���
�S�Ж{Ƴ��Zvt���M�y��;V�ds�]ы���E��c�1q�ђtq8��ؗ�����9.Q��y���*}h�Om�|i�>�6����ܝ܅�C���;G?Ew�a<�ڵ�ѯm��� �W�O!�N��>�����}s�_do[.=��c�U=>�Z�3W�ʰ�g��X���H�}�ݙ���|�"~�$�vee�U�/��E�3f���#����:s�$�n�`�����u<>E�w�]�9{݀�}���-ME�����Y�m��L���
=斦�fm�^V[.��󷩽G#]R�����T�.	�L�m�����6�J���FE�DVÈ�Hu�Hj��u5j�SYjb,�2��o�;��S{ufU<�0���'hV�ӓ�9o��׀twy�r�Z���n`��*�2�0�ɶ��F����%��iP��Θ:��L��YWq+�Q����mܾ�Ew�*"V󹈉iv�tl��eJ�����M�֪� ��J�Q�݉�U:��`�����`��*NrY3s��k)�:�:��^l����J�u�z�\1��o����:-U�\5ڴ]�D�"�����ܰk[�s}***ݰomǔ��X�yXI87!\L�[�]����ц��n˘ˤs�5u�/\��}{��sS���$���[Hʚ�n26Zāǻpk�����S:��iZ#���v����\�`�9,ft�0���.�B(Q�e�z��\��W.��#nA���\?E �o�K����:o�μ]�J��o-�U&j�u܆�zTu˳��&&�qK����w[<�"�@Z������Ѩ�nSt������4+\	���Zr������U�\�c6���H�o�ֲ�૞���o�UQŕ�9�����\-Ңm�����·]i���qW袽����+��;ܮ���0��U�º�]z��*H��;�o�ӯuxɅ��wh�x��wY|pWr.�ѥ\���i�
go�<��=�g��J<���)LIʆnzb��.��fC'wS�59{ց��IXI�� j2ٱ�X��|�et�5)a��
��5��WK�W���ˠTu�O*��[yOɅV��ʜ��>�37�~���}:6δ/Kw��D�~|��f=��U1�)C�+�7f�h�;�3��2g�<o:�(�@��n.��ü)_
���o��-�\�h���Kؔ�w(�-�mvS�Enk�7a�ʣ��0C�+�6�nW4� ;Yt�1Z�t�����:E�>me�Z�m���.�mu��/S<�Yrf��#�	5��p��wS�ܗ.��y�'�Y�e�p�厳WqL�|���GV��8dHw
�@�ӒU�p�D3����K��	��f�*�Xݸ_*6��vѫ-f�x��%M�CUr�r�yh��-f�&[0o����w��6�ͽr�)9ı*]'��FV�7r�ڜ��*�+�vT�9/5CR��c*Z�{.֪+`ׅC�.k�\�:���VAС�E�H�;CCxw��O��GQ�Z�&+gs,�{C,�[�x�;����ώK {�@*q�I�S&o �����!����5��u�vf����Ƕ�3�3�Y�R���k�7铡�j�� �P�V�T��檡��mlA�l�V�cMMZlh�gM1M;glDMkEQ�&)�"�`���J�؍����m�L��j"��J�����h���QN�i�N�i��E�c0QD�kh�M��b��h�����E��S\�s:Z���m5h�j
�&*�1ED�[8����j�;bض1h-`�*�((�*"j��l�٨��AQkE��Q���Dkh����.�D�UD�[X�գQA5UT��1��m��UU%IQUUEE1[J����QTZ�U4ZtZ���EA���
��m�AU��#jq�U,�m���(���cL�Z�CQE�%LQ[dѪb(#f �L�MS��c��Ll�*���%@P�MF���_+�\t�/T�1�{)C��1�t����G���R��r�٩�cT���-��xv3
ݍ���K�x���Xr��u�vp���6s*׫������v�f���ǢUS�}�*cZ��us�odQO�}�^�����}qt9q�~3Nu�7��O�@��}p�
���O�����s�f�󰍌���=j㻕{�F���rp����::K��*��%�дP����
w�ӤU��~pb�e��y���;�b�MŖOp����z�ng�g�%E�,��Z�;��gfL��X���;`��P��t��S��AU�0��(�$�A�L���&s0�s�����vT�f���O�iz�/n�=���:�t���J��=%��΀�f�ȱ�{��ޢ�����g]G_�e#�uQ,�R[q7
��>�!��}��zm�T�>�P����>��<'<)�fy�L� sQ%	L�w�uaq�R}q6��q��ó▯z[/�,d{<m��_�v�e�][5p�AF���=S 9	V�`�x{�@�\n1up�2,�;$J����*����ec��9��n�廻f����GT������}4%g�xV���ꢮ�hd��S�]���Pc�5n�$�fsą�ʺ\;-�����-��[\̚��p�}fM��yU���y�R�Wz�tio��"����~{�8�\�^ݞ8�l��-���N�:�JU��q�v��T䫇���d�>`��������˩�o����̕�f��*���2�����pv���2:�܉ ?y��Q5���c��wFFo��GmpW��b����Z�9`c�W�N�Dt�v6���!�o6���
��TWҕfQH�_ٗM�����&���� �:`a}�h1��~ۋ�<I����C��@_�+��ﵰY�A�����=;^����腮�tC�����Y3uc/.+}j��4+_Ϸ�.8����>�:�Nu�c:�i8w6S7��;�;���i�w*�o5ݘq�V��]��߯4�3<U�U��Œ��?�cV�_?�q_M����Μ���¯��^��r�*���ه�����T�|(�+q�� �^[r��<'��l��{]y�eyOw^t�y�k���`w�h!GS��;��{�u�t���\geN����kr�J�h��n^
�|�z�=Z���̺���T���P	F̆n�Zy��s�s�w|�D�_5G�g��b��g^���)�t��D�f��C�_�ەQ�Į�xk����2��c�O�=�Bb��r�v�tQ���V,G�cC�ˆ�>Y½�o���ԫm]L�ө�J2�}!���<��LzFʮe��u̅C}B�6������t�\[ QB�&��Ow��<	<T�ȃ;��l	\Ǽ�FM��D%jYրsi��ٵ�E��2�'���顎w/�x��I��e0T+��R������q��b�����ل�d��]�̔3W�`����Q�.5�GVuBΈ.�����J��q�`4��}޺L�ʶb��,�wb�>��uo?�m���G,v��v��w.ݣ�IF��d0
[$*��¢`vWn�=���߲u�΅k]���tա�/6��N�I�x�'����Z2Q� .��gkS�}��-_�DÜ�*7Gt����zF����~�9�d�6� ��q4��k�{����]���h9������&%m*7V���v�Ԍ�o.�&�u��@t����E��FҎ��`8wXFͩ�e�8��Ҷ�UԦr��J�}�n�M]�rZ�h,"l_U��af��&K��P�E���ɮ�G����l<�����[LWf��L�z���sW�f�/t��	�Wzak�tS�p'[�Q�/�ޖOTL.��b�����0<׳2z=���뺾vM�J��x�%O}�k����x��vl�[�c�l�2����sCo��D6^�Dh��~ҍ�9^b�g�s����U�9o�C�q��YR���;^��t�z�]�3<b����ݎ���=1|�NƄ`��+�;�����;pi4:	�Z����'�u�����ۥ�j�t�83�\�(r�����}R���h�s��3Flv���1S��\u��:�����T��;�땜��q������p|��qlo�a�ez�N�KE�<��x�}Q��6jS'�) ;Q��nK��=�MWr��z��"|:7��O�'5^[��Jqs��ˉ���w��q�ە�胲�(�,����c?'�0�`�K�J�"�vS�G_�j�w�G,�ӒtV�N��p��	h����U+g�^S<��� �M/?a�ڻ�ٸ��(��g��\=�^�B=�Q�����P℞�{�ң��>���}5����u�]�B_���|!��3�ڸ{���[f�^r�N�d�J��l\�����Hgӯg�먕qI{D�)׃Y/��}G[��8n!;w��YI��#z��M䘔���O��l@�83`��$�_	��b}q7�{���|w>N�i7�茉�x��VU��Ev��y�WzZ �_A $�A����5��b�Q�	;H�����O�G�{>;�{�����ss��$O��揹J:�Kߟ)�G��3�}��7�ִW�̭��w`�#����壋io*?)�-X[�i�%��\ F�3��Ų_L��v�}<wV;l����Y%dٱP���^i5�����}�k(�7��|믓&E.�NZ���3S�*�S�����u`n�z�7��f:��|_R��h˵�DD�������t�fc�.9Jd�2_��Ji*:�N͙��6=���h]9�4����������z�:kKmQ��1�:4z�_�
��[.̓��J�+lE��C���e;�Z��a��(��~��5q�6����rwr-c��m9`N󸑮�A��d���fr��z�o�y#�+\@��m�Va��Z_f�����߭��^Z�3W*í�7�a6.;z���^�},�wxۑ�!���>	�9���S�$�'�#�S7�=���TƵ5`V��q�zd���7��ލ~��X��t<�P���un�hl�'������҄|\��\I�����>��Wx�v�#��q��w�o�7��N%�tv�K���4�>��XQ��V/}N}��fO{{���u����P>�u�쮨��N�����M�d�Y�=P�C�s��;���o�ՙ���nndc�
�=聳A�|1�\F(t�y:L���)�0�eJ7gI;juI�A�^}��7�Twg)���F�n�/Z^��[��z%���@=�n�z}�Ҳ�*�\��5}��I
�]e,� �a���g/,ǉ�)�����e��R�sL}:�|h*_����k��܂�~�p���� �.c�9ӲV5Y�!�%@{�}����ӛ,��E)C��|6��K
�V�gDcTȔJЧwY�Wfv�Ud��HG��%��te#ވ�]ĳ)mD�T�_��5;��@=99�>�ݚ��X�Tygz��z���y��c��t��5P*�@��uaq�'�p��q!G��
cSF�\�wW���:��Ʊ܌u4�d)�Q��4� ;	V�`�zҫ���m��gLg��^X�v��5��hǋʹ�9��n�廻f���J5�T��6H�I��C)���O���������_���P�����K��=��Ϡ��%z��Jb}�T��3�G�:zk��jGN��0粕�=�5q�L=J�1���䩒��1¨�2!;�����>O����p�D����6w��Y��E���P��<�j�M�t��;`io*���8�b�w�B����\�_)�z���9>
��a���i|szV��r�p�uZL�^Q"��d�������{���/�wHV���8?L�l�x�Kp-�Sq�KI���L����2�l׽ǻ|�}�5�����N3�5��ۏ߯4�6���rp�?G��ڟQ���S�{�/MŻ��u�掾�m�t�Nλ�6��	��{k��*� _��"��FR!6N�ǒ���׺�-�R�H�+����X8����w����V�����圦71�l�-�{n�__��+:��V���N"�>[}'k7]��Ro\o$�Ӊ��wWx�ᎉU��<�����X��^�~����d��׀S��Kk�Y�P�^l���xΗ��}�H
�W�����.��������p���5ul��E�B�0�z�E����.����3�u�\omP	z��7dZ���q��k���1�"������5���h�ܧ��ʐ�.t���JF�3�
⌾7�*�q�]���O��e`�N�}=��l����k-�-��<1Ĭ������I�Ix?s�F���lmq�ӜϙP�o���徛����=��t�^�d3�:�o�.���|
4���_@L���<-Bh��{ޣ�6��v�m���Z�*�;���]�:����w-��0�=%� o]����GN���w��sϺ���C'�Ͻ�c������@?m1��n���O�����Z2Q��9H�߅�����Yb�<LLD���qE�y��P���H�$ա�-���s�ɶ�`��G��y�Y��M�c����q.!��f���n��>���n�s=��ێ]nM�n�1̘�������Ek��.}�_v�7�Ol>1����A�ѧK/w��q+kkZ�>뛠�R�����t=�˂.���w�]S�~��s�Ù�ﭑ����9-�J�L�{J�]b���Hޙ����v�&�;@A4ड़��G����������x
�GM��fS#��DJ��RS>��+w=�kg�j3�Fzp�7�����2d�n��
d^�s'�a�>�6�|��Ki�=z���G�>���5�ڑ<�o?&?W�Q�.��`���:6�\	ۈn�·�6r4�z<av|2�'��6��_�M�������)��ݤ�n�1�J��<���/L��Ǖ�q��O�K�c��T�+��j.=�{Ly�^��piV��:������N�s��W9��z5�p��ϕ:.�>�D��h�k�܍E�?����+�XD��큔�����u��u1�n*�Q�{B�{����F��=��3�Cܶ.3�$�OdL�vc�N���ܨA�p�1�&M�\�ϽbliF��o��o���ƴ���Q���w�g��Μ����w"g��t)%�����J��\�E �2	T��u�k�[��%��̔�O�m�g�*��U{���e������|P��� ���G�5P�*m#���﷧�|����lh�k�Hg��g[U�3	�IF��O`�7Xf�C�q5�3�Xn6�(Kz��E������;;*��q;,�kˡ˭؜�}��1.Ϭ
	�9�gѬ�����<\�osy��5��4[;�:ܥîT���M�xg]��;��S8i�Xռ��ɘ[+RO���"�e�����l�F��)Z��e�������<7���$T/�z�bV�^�"�Rw����G���p����8S�P�&GyϏ^�n^4�>�� ,��" a����ZH�^�\o뉷O���)�|w!:��%���y?w��Υ�yVܲ<�ݱZIS�@��$��;F#�]X��ќ
O�!�E�?4����ށ^�Wv������Ru�6!�[5p�IB���+���1)�
��V��2�WZ�+f��{̂�V�x��zܛn_�f�.��4��\�ٿ���;���Q*u�3ޚȵ!�Uޫ<�m�;�O]-=�H}�����vh�r�/�S�W����a(ii�եk��ɷ>����Y\�×��{���5~�C{��!�;��SМ�'n9�(k��ryl�RS듚غ��R��zc���
�0�G\�/����yly*���-t���Xu����7�'�y3�sj�z�N�����z��9@�$l�T)��;�a8}�l�}���J�xKNJQw��[̝ފ�ѯ��Z�|�v�g�\B���^�C�#���m酮�O8�C~��շB�����񣟁6��s���9`��)�h�E<�A���E lr���gM7�՘5W9Z9]6���;�h#�oFͮ�Z�v����b�v��ˏi��������y�&]>��";Cf�|6�cp==Rf��uޭ��:\�`;{;�T�s%vɬ�P[��➩��se���Oü����s��xo�8/��9s(z�::���YO΢���>��������/�;<\w�z���#����N������?�hg�i����
��r���l�a��Z=]!�d>_v��1��N�<�x<�*��ze\��`�������u�3�8�R�O30��A�Z.�{���1K�iz�/n�=�厀{m�O��y^\mT�z����KYT�(�x�t���(_T)��W̥��S��B��]�+Vm���zB����ip�T�J����U) oMD����v�Յ�S��K,s�Zq�nx9̿nz绯�<Y��+NBR0�w#-�Z5jdk��=Q2��A�)��m@��<X*�>����s=�Ŧ^iq�R�N�0��!�x���9p��
d�_uI�d��0nM፿����ꚰ�rh8���<:PV����K��=�o���.|�^�j=�Z������zņ���R�ܳ���}>o��a�>��k!Tgu�BҪ�Q�ԉ^�
P}Q`~��E����PE��N"���� DW�`����"��PE���� "+���������E~* ���"����� "+������"����E�b��L��N��3� � ���{ϻ ����`<�zPQJ���� �*�)ET�@P� ��<�DEQ�)*���m$T��IJUI��+��B)!J��T���T���%R�J�(�H��{�*R8 e!�f�" ��&��Z&�,��i�4]�AJ�h���ꝄP� �p  �   6�  m��m;�]k7�UT�-PI� ��6�J-Y�m�c(�2��f�֬�&V6��Dm�(p�ښ�R6Q��DɖU[44:�E�iJ	�(P�IJ��nhYh
��$�5�T�EP;�֨ * t T�
��R�p�D�P�UE:ֶ�[ 2�(���H�	)Eim�jKC �P�+Z�P� a�kN�4�(�T[b ���  ��P(QZh$U P$Ũ�Rk* ��V�3j��Yblb����kZ��k"5��b�%� 0��h��hf5��L�m[k�0M�,m��l�&�%$6e*�p 3 �a�� m+j��5�,0V��cUe�!6���H�@ M�
�H�``1M)�)JJ�A�14i�F�&MLL`���~��%*EC �0# 	��h�L�h�FSȧ��H�2z���H��TP�'�h&�	�� ѯ�O:�T�V8c�8ׅo{�e2�oi�K�h���©C����A�A�����t�����>��**"�aI��_�>,�����hC��� �d�XUV%�M U�*��� aUo���j���!��ǰ��d�����tbT(���W�J04~���?�N�������7��K���?���1�~�H$x��y�XuY��~�����j��Y�>+��N�H�zzЦ*b5��A.�u��� j�T3+t�sf���y�q�c@�I@@����i�y�[E��;�wZ�o�=��QDN�jl�W��4�yJ�:"�۔��Q�"x�t/�H�Ňw���7^�C�Z�ʇu�y;� �Z�f�>��f�F��h��Z�c�i��4�A�RW`��7{O,ubʪ\p�W+�Yt[@��9��6.��Ysp]�ƫ)��Ya��ũ��ea9��N�c*��II,�h�rL�?R��%"���Kt�F�����(c�Ŏ�KH:��o����8�nkPݗ^bzr���:ƜZ�7{ekj�n0r����� �2�͡�z�}�k�W���N��đ��WfTQ[��lՋc��7��Ni,�U@ۥOr����+���ݓ��	C	Y�Inf��j��+*�j��(�NV�80� �K<��4�3u�YF��Z�$40��d�iK۠-�΅��J�5 .QIm��0R�x4��*����1M�WQ�ԩ�F���5]�(]	YMe���W
ӊ���B�nз{�`gb�Ж+��]-� �--��b���l,X,]��sT���B��H��Vt,�)�Ŧ�Ӣ^�&%�z�٣ ����l2YC��vb;Hj��#C�71�7 �Wf����i��4���c�ٯ&f�Z.�a<�7E�4���~Yω'ocB��o�6���-:7�h����`��_a��u�̉7R�Q��'��Z�z"$.P�l�ѥe�9����޷�})L�ޓ��+�$t�7P�P+pm⎭U��9x�f��;�x�r�Yv���!7b3]nR�I�[d��RCA��ݍۙB�f�b�XT����vS`BҐ�X/Y�I���ߒ�X��+�ch����Hp���v�"��4<��O��݆�x3tq6�8���v#���j�ɩ00Q�^Sn��.�G�m�omdx>u9�aB�
�V�,B���B���b�����P�.��B5�Ѩ��m]cAF�!iL��#J�f]���d�b{x����V���xrxj�u:�B��ޥ�r��9�S��9u�f<�]����3&�PB����)c_�F�]0b�J���=۶0��M���2�Έ��D�di�X	�k��y0��];��e����k&3%���0e��{4���WB�;�HxW�>ݻ��E�LuZ��RL5s.��
`d-��������f����4-��PW�$;3u�J�(�tJ{����a8$"�M�.��@Ͱ�J5�"6��[ٮ*2��P�W�R��t]�'2���� .��˦��.�$mӤ�w2�ɀG��˚o�V����Fe'�jR�Jss�Z���ؖ`gj�:C�\�  4nP� +g�$��ͤ���f�wv������KPFZ�>CN��$�`!���.cVag��%Jf�[���!۫U���5h�guj���MvJTδl-u�RA�q��ӑ�X�ߡ�&u$ʳ3sr�-�^n�IYC �A�J#��V�^B�eV���: ;9E˫Uh�K��o��yJ!�X�[x J7t��s4iI$n�{L�	�6�Y�N<�:�"6Y!ۑjX�j��h�e,|ia����ƜJ�;�/�h|Q�MT-MTw��%Zڗ7��w�A�qu�K��:�Z-u��Xz���k�R�3���)�n��[s��De-MLFj�tL�LY���h��]�Gh��%bY��uMz�WL��M-�N��P�uԨ#�&U�w����Qi�X������f�"h'��&�����]�pۮ��q��\�b�s�������p갎����ᨭ�H�4���F�,�7�t�������
�Psh���[2��d�7*]��09WV�b��*˽5��j[�6�.G�i�D��t��>;�n0��t�=�-L]h���ԇv��)m����r<ɷiG�i7����ʔ�j�4'1V}�����d��r`��cy2�uwZ]�cN�1x��.�T$�U�\���;�;��e��U��^�"s5E&����(�)�����T�X*\���y�< �kq�zVh^-�v��:M�GQ�}d!t	�ov�7��Q�ÂRf���Wa��5�x�8� �6�Ѐ���cf�U�ħ��qQsTn;��	�.£��y)=X3N#G7�ةbh
�xMkݣZ�uwV�*�X2UՊv�����Mv`4S�Y����b����4����F6}oK���f�M°�yR��+1WV��5�K4ɣ�R�)�k0��Kh��wgz��Y=�sG9,������P��M�kk��K&,R��d
��D��;���6�J_V�'�U�,z�]�[�hf�J�^���:�)�6�6X����*6j�s/^��,��n�HU�m`��If�c�cJṇ�X�O3�m[��VcW� A�l
�w��I��҆��s ��;��t�L��
����	�Җ,a����H�AWw�,�FJ��I�v�a!e�x��&!.S��A��Ā�@aF�Q�H�]L+#m4i��j�N�6��۫2ml%��8 :s�k�5�P�כO>�#�eY5�faխ�������'���W,��M���J�%պ�6v��peٗ
;�Y>��S����rԬ�2���y��ܰחt��hm�p��L�ц+V�h2���]��q�;���"�3K+Jڰf�����tu�$�k���eK�D�/oo�*�ůF��`���W���oj�Qɀl�������S_�Q�HV���\ի(C��\��c�����=՘�k8q#v���	u������T:��ĳMlKm&��e��H��4<RP�S��,��׷B�C��Yf���J�PB���1�XM���ܬ�x�Yɴ�v� [Ea//�',ot*� ����W�z��J�m��(Ֆn��b��^����`J��D�<&
�DS���"�unܚ)3x�S6\{�N�a@��B���C�ͺ��z��m(+p^�5v�X[��op���'x�Z�K�:��}�v��iK�!�-�a�2� 㶓��w[�7�YWYc/4�֔�f�� fL%5ԗdYo�!{�$��f]��,�״-�T_O�驁����,$nX��^��QHM]�rȳ�SL�]&��HM%b����s>�l���j�ڐ�Yi��\y+5�@�[��eŔs h)ij$ӱ� "����51f����b��V7�M�"�ʼ��`!�2����^ųE^�T�U�k�5�:r)yW`�)i{D�Y��ha�s��G�=w��t�s��h��le���݃�;w��,)�k�N�� �aL5���Z�O;�=�����ng�^����;�d)�ea�p�Uhb�cW��͕�zd ƔM�ٴ�r�c*P�P�yL-{��tr���NP7����y9@�o'+כ��^��%ӫ�����6�m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m���m��q��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m��m�����r��j�����iм�HT��;�\0��7Gf]�lU���K���+"sLv��8؍��ˤ��J��Y҆���[��YV^g7���)�h����w���+"��FS�P0����ԉg�n��uB�v��Vi��])e.D�Ǜ�$^ɓ.f�+�PI����(h�;�yN8)�Ugt%�u�p/��B��hX�N8�w��s�ܦkCbue�g,�ݣJ�e8Uo2wlՔ
�Ҵ�Y1��5��i��#+������g�`a.
P�C̊n��-_n���TA�h��}�y@P׎��\��"�@T��O M��������CG�4���ճ[y��%�g����U��*�7�y��]g�ǚ*^���'KE�ɼ��V*ۗS;6Q��!��F�Q:�X�W�8:�>n򰱐���1`��i��o-�᫪x������<U����R����y쇺���m�8�n�f�Z�,�Ex���m!��
Mخ�٠eKyڅ�K��`�m�c���Fؾ.���u��V(�(�Ի�;z�w��(��� ���_��r�u��w=Y��ol���Ze2�fp�nK�t�py^إ�,��-e�Uc�˲��H�[�0n=k6ʊ��Y6*.l��m�t����{��t����xq�!\q��I����`�DՒ�2K�J��̷jջ��)[9�!��;�Bj芵x7Mr�Q�Q�!嗂��CM:�3���e��碘�G҃�S�㻗�#���=N%*����b�ǻ2�iqd�]g�W�֚��B���故g��WN���g6�Q�٪���Wy�՝�#4����db���|�^wH,�$0��fMV^v� ��:3���ۡ�-�Pl�8Y���n�=��$L�x���r��(���/y�bu�"G��x�.i�� ��b���J}���ZNX&&�	u�¢�ʽ�5�e���6���-��)O)j��J:��>1���Q'��Q�uWd�{OW�d��+Qw%�13i^��/�'J��@\㰳ګjgi}��`Ś��#�5�P4�U�{]{�S:8�WӸu��m�Lv��v��'�[�,�.VU=鿨�IM��J�.���vܻ5n�37+�I�����s1Vq/h䩂�KL�R��ٲoM1񦉂�j���lM��E')�u�gVoJ+o\�G+L�D���sg�������
]���-�~MNY�ɑ��{����g��k��3����M�	�bY�v� D��׽:��K���/vi�]u�䳺t�a嗎��*��8v0v��9'
r��$e��<��gh�CK��z��Rs��kY"�(eL��l8�{���>%ņj� ����(�od���Q��\NU���z�k��+Y�ɛ�t��β�HlNJ��tuC��(g5��L��3����*��;*��yG�0�n����,л��E[B�}�C�\hn���Yv��键�wQ�����OL�-�u��ۭf��g��
�}K5�R-h�9 �\U�3��8�aƀ�YV3�����N�Y�;(II�ΏngV����m㽹ٛM�4�����Y)U��DJ�܃32�kכ	���tyӧW9L�8��4�s�A��
`6�V���&��f�Cu�3�E�Kh�an�%��
���y���a��{�ϐ�n�s�/z-�4��X�lm!A�vm:��+3z����rXx��f�0p{˺�j���Ì��I����K���K���v�N��J��{��t>Z�[I�	��1��G�TR����[���ӣ�V�:IZ�ݙ�DǍn*�*TC��:���w//-gdyQb�꼔pX!8����^���ns�=����*��Sbu��J��^�up��J�s�.Ь�b=��4�EIʷ/���u-��u1m�veixۧJ���������T[ct���=LI';x�x{��>Y��a`�
Y���8�\�<�l��sm:˶/i�ff<6>s�=s�\�ڑ���W[7a��J�;�S�V��+�t}b��)T)������Q&��}sBȈ`B�D�+�+���)D�����ݛ#�	�Ck9�*���3f�Mcμ��x�hv�Q9�I��5�_��Aԍ��n��!$����R �K�I7"�H�';0��֥�u�,�p�j�!N���:*�7O�����G㣺�Cu��LLgnK��T����+�-�]�;���9o"��"�m��$.n�LT��f2�-�T	��]�Tˮ���l�y�'c������HBǯ�3���\�ir
�ڮc8����Q�d��Ƶ?�X���^��� �Db���b��u��s��kU\C��Q0�r�J����vQ�R��F��B\�5���t�h�"�6��X�,�(#�&8��}�:�6�!��C9�4-��f���veN*����Cf�VfS�XHa*��-Ѳ��C�N�D1晒V�3:ׇ���;/v:f���䜺:���o>��Wa�QJ�!���网Z��(j���Z���^��OZ����^�fgk�$���H��6�30sÓjZ[zh���nB�w���+�"��7��2�MOt��sN����GN x�e��R`=X��<'E�hi�ݮ�Y�%a�36��O2$�J�7Me�c��o>�K��1P�M�i��]���K�%݃�P�V��	��_H�ٻ�v�&��V(��@�Y|Ἇ��'	y;�*�aʹO��ө�g��S7��k��w�����Yd��x_m�
�T� P[[����-f�Y�37{�=ˑ�-.��
��4My*a8]� e�]�Oy�3��=�o���9h0�6AZ=��5A���iq�c5���v٣Y�/�î�
7�(���]��F��͢�.�P?[����y)��M|�e��d5MW�%³���P)˫�4Ї,F�\c7��-�¦�(�f>�A��N\7e�ڎ�5��it=�(pt̾]�r:<z�LS4N���6%go�[�����B�OFdmts�"���:XL�M�1��a�fv��T�4.�]��\s(���>ŧ�wVڨn��H����r(�1Ǯ޲�i	¥�����t�|8d�蚫
�t�{I�J�n��Oz�:�ZӃd㽸T�}}Y�ִe���·��S���_t�*��в�K�ᦋ�mm���J\\�y�0�l�1���Ypb�꺼*ۻ�,�\zK�Le�❜d�[��Ӏc�㹖�HJ�ض7͸�u��_s�=�F�y�����ȑҦ/�mJ���E�J8����N���*T6�:��E��lܤ�4-�V�gwe�a9ȃA���+k�����]��m�F��e6[m��M��m��m��m��m��m��m��m��m��m��m��m��-��eդ&�mҳ�r�޾jɜ�tn,��l��m�������k�����g��(�����UT���Ia]@ 5�EEG��tfB��A^�����,�Ѷ��P�/�0����윚b���z.���ܠ�Ծ;6��x�(��L��vG���r��R���9���.+����,�u�L��>�YQݭ�e�;r�#�y���VWJLĝa"�SOJ��B�����d�y�k��.9،�z4-ΣS
mjD"��_e���]�Ci�+�!�f:B�CNL��{���@S��u�$Ww�'=3)�V�sMi���f1x���4�|�f��*nڠ��9dG[E=jɂ����$CF�pc���8q����v�pR�AΦ�-���Fnv�e��i�k+0�~�9��t�P���X[°���L���#�K�*�B�J�3_K�읜6��62ik�;z.n��j�ڱۧ�[8QH�%c3(a��jr5f�yuWT�uTXE1;{�b�P�,�t�G?K��d[H�\�딲���(�:Ph�7�f Fɦ���J�%��� ���Q<nɘay�
��i�&�l���,�*ȫ��vφ�y��C��zPS���b'��oi�͇!�z�	g�׸�]�0^���D��I؁U�[�Y}h�toe���x�W�Ux�=��ٷw���t���h���C�*W#C��#�5;����B�fs�
�S�]�t�:�1��`���>�#�`��.[���B�(QU�K'6�.j�]
y\�̀�[8�{��7	�񳧡}37ǭ^!ki����.��m�����n;�����Y���t��c�<�ג],=x	� f3��d##ܸwaw3ke�X<J�0�]u�ni.������с�{���>ـ����8|ګ��&h�t�Nѷ�l4Gc���|7.�$U`,i�0,n�]��sO<tM�L��@g*ZVю��8WY���Y����B�v�x�uc�v�cn�:j�r�N�=Í��Y�&�+]:�VT�t�+Z�D���{�>��u�e���*R�y%��Mj-�Na��w0�fq��Ϟ#2�[�쭘
㎗E�.[���ө%zv�K5vK��ӣ_V>�cl��ur!]w�;[��D�Ϸq[��]�%�M3	|��]ݓ>3�$z��V ��-A���g47Qź���[��v
ug8��)�Uҟ��왂u+�h���#�ti����
}Mq�k��3�"@��A=����5���']�G
�X�hz8�SY���N>Ǚ��n�a�vjƲ�|���;�Sus�6}�f]L4[��sJ��4���:Y�M�ow+�����4r�%�"9��5�ol�cR`�N�t�!�`�s&2�b��6�1�{{*�?�"���*���ɥ1��l���y�%�E6ȳ���wA���a�!��o�^�2UfcF��\�e,�Yں���zX���S�+F�p�ڍ�vl�3���7БV���uج�v�z��B�gs��f��J2�]T1f^�͙4N�f�Q�O:�cL�bcq>��Nn�8պ��u��W2S�t �}�u�,��[%u�t�����P�{�ZF��Tv�r�H�:��V:��U�����Eun� �G*��Z:����%;��v@5,�3�8v<D��6S��OH`�|�<Rj�fu�/͍��w�F���]H��H�I��
�k�U�Q�쿐�X�t���]�B-������s)�md�Twf����B�G+h���WgK�B`Xm�>��7�b�H�,�εx+d��\0񮎕�Ne`dE> .\u�[3s�N��QP�ԭ��rs>'Jls�{5@���\Q�ul�����0�w�N)V�&��"&�QBa�[��7��m�%���ƛ��ioEU-$�!{��Cq��|��O3�?��4�w��f������[�O'�8��y���ם�$jWDP�Ҳ���jg���u�w;���]�qL�N�z�S���>�VV5�䊕���a	v˳��w����8�lx+2 M5}�R��:���u����q'���\����l�Ik�Xd6o�rޑV�\Y�d���`�;N� :�!,���e�F`�v^��2���}�ye��7�(^�d^��N.����D�P+��V�IZ;ll��]똃���K7N���\�.vLf�dw;V���@��+�F�[HCΥ'�kEƔ&��.$���6^4:�v�.�;*��:��S޳fU�k�;�Q�ū��C��f�D�����3ڭ-p.*LN���ɬ�Y���[�t���^��8�4�72�N=GQM���;�Ʋ2v^�b�� �}���>˽b��Ta�tp�V�{ۜ��#F�3W|n�\:XX�FѮ9ͮ����L���QKg
��lo}���T���f�#]Z���In�ð.7���0VJ��2�O���ȑ���p [R�t��jH�8��Q1�Q���(�t��켛\���v��U�N��q<v�u�L�ڹ��zT�k4��w1�,�3w��[��oR?w�.��V�lF�-����m�'�]:����a�Ҕ8[�1��2����McU]���'�GQgc
�o(��0ene�,��`�mC�p=�
9Y�e!�k��WYpɩ�؂�8��]��#�b��t���_V������<�O^ИpW;���,��2�Wp(��7s�$4[;�W���ßq�53c+����[�J�'P9��\4�u�jN��hP�0Z������+����/C�'Y�lԳ��s,���F^��U�%V����\)��-��p��%:��v���v��w��$��\G2i�x��IV;��Y���Gz1X�Ȇ\��Km'�I�0ܔV��,6�qY2�gl�;A�8�����&R�Q�}K�qQ]��bޕ�n�p�o����B�ξ�e�No��>�e��jWv+�[{�|�Ê��V�߯b�2��^dX5d�r�Wȥ�2����Ӧ��j���+�ˎ������]SU������'+�{>�DG�sN��zU��ׁd�n��ǥ���iS&���:E��D+�����/�@���}��5��tҮYzM��}�y]�=3[=�]���u�;u<��Ʃ�y�I�l���{�x.^���6ͧA�l�఑���(�C�k7i�i���J��CՐ�U���^�d��g��W���G0�bR��=9�ڳ�e�ׁ�/�r�k�Ǽ��|y�e�җ�n�];��NU�kq�Ő���P�
��4췕�g;98t�1[�`JYX�-�$�Q�ݦ�Tuem�5֟j܁�uB��L��+��T��m)
r���
-C4����dX�az	�%oJ�_#�UH�������4w 6���ˑ�o
xuVỨ��{�k쭊�g-�5f���	��f�F���DOw09�R@�k��*ϭ�fm���B��Y�5fU��wȂ^�J�rt��;���,ѶR��`���HAv�0K(g�NXT�
��:��7Tu���pֺ���q���μ�����Da� {!�`�'���!�za�׾��YNw�k׏����m��m��m�$�/W��1LTx<8���r]��r��m7g��j��jݖ�����W�Tˡ��͋�tw)$Y��ɽ����f�<�\��*�������E�D���s�Ү�t��:�
�B����_L�ǔfl��ne�F��jTL�z,P4'oo­X��Ru�����m<�/�7z�k��Y��\�䁣G�7�=Z��R�#>쳠�xG������Uܐ�JC��d��x��8ی�E��f�}u0�6h��P��]9N���2�3r��7�#��;��a�j�K�_�[�f[�vn}{[M*7y\�=����C�v�L�B��M�,}�$ 8���1�^I2[wݴ{w�9�s�y�9�}��0=C�̅f+Y1�a�N٦j1Cib�UՃK-,���b�j��A���DL�¤���ge̥m��NaLWyfb�E;M&2i�"�°���"�J���*U�a�ʈ��fZ-��%T���̲��PSẒ�B����Y*���CL�Q£J�cRQ�X��dD+��+P�ʛj�)��f��kJ��i��-���R�)Qg�*:���`)�����L
��H��V��Q�YU+-��T
�eKl�����g>��=� �mJg������t5/7�������*��5�Q����qI������&�fK���֍T���k�f.��g���8�T벊��(�fM��ƻ��E�Y�=y�Ѳ��M�iN�����j�4)�^>���O��n������eܞ.�m��U�9�5���\]"�������������)��jZ�����{A�lr�T�)'���L���kW�_?40˒p~3��˺{3B���ma*������ߥ�m?c=����_���F���)���{�w��N�2c��sur�w"t��{Ե�Բ-D���p��33\ΑWE��q�i{�J��d ��o_�	�]y�l���J{������������|J����Yٲ4�aف�=YҸ��R�M���8�P�]zc��=�j�Sމ���W�v�f��k&��N�H=k�'r<hT�m�x��_�|�i��q;�K�^
��w�U:��m�)v&{1򎷻����.�e��D�J�À9$��TFH2���Dڻ�-��.�ZP��=뚎�iQ���>>�9�M��-�@^�+Ao�n��2��ͬk��Auj��o�:m�7�LK)d�wvfo�"��x4�d�>w��BA���%$����]�~�QZ�TE�s��U�	�Sױ輹��VT���V�T7/9�|o.��9z�yV4�[�l���[���q��2.5۝���������켙�t��Rd��|r�r���><Mo��==��i>����g�:�{�+��\.&,d���O)�/���doeEu���^��&{jV��"wM�j����8�7ը��3ǣ���Uߪ��wݧ&D}�VV���b�lV��S~<� ݾ��,��ef�\b�����h[S���tjw6^vtI�sZ��'3��ok3]�U�'���^k��5�&�6�u�{sygM����o+}||��1�L�U�
���w��Q6���S0dn�j���gP�2����6��o&}��W�CL���v%��d��~6z��yr(��Р�M��ד͝���p�ﯮ>�g\F�6��V=���o�)�39�\��z�sG=�y'P�Il���Y˧5C+�B��+���-�PCV��ؠ=��Mn��
i+b倘7�#�$�*H�.w֤J������e���r}��{��&]!�d�1��/oN�*�^v��/f������(ޒ>�uA�&�ORڅ�ތ���8�0��V�ӛU�]V��q�A`� ����D�芻���t���"3����Eg��R�Z�%���J����{���sH��%�
� Y��sԦi�K�#� t2�n�q�E��f�2e9x���k��)��قJ��$�tQ��^�=~ɎîS�EL���KūZW�>�Y��R.�
��fv���x�>�����A����ӽB'�f���|�Iԛo2w6;�5c�[y��6�N��ث�V�Ϟ[(��V�Ө;T��s��>�����T��_=��ZJ4�����]gn��4���U��5:�v���jNΝ��o����ޙ����.�#2��S��������iz��^�4���O~��n(��~ΒOfK��i�KV�r>������uN<�x�Xޭ��=�:sٺ�c����=�臣��x�d3���!���l��R�G9��Q�g� Pf�ٝ���d�W+`��ۧu*(U����;���1>]�&eŴ�N��r���䃔�5]��sA֠�{�P��kI����u�T������E{ڬ�Ζ����f����Ө�]xv�l����u��^�L�8�yw��b
Ʋ�˸��F��#V���W�TFOLʔ���Z=˘r2��]b����j*��pw�K^ap�.�D��tY�y���<�����Y�gxs�n�{Sw3��d*IXy��6o��í�K��ݾ��#����c�m�[���:6�z�{=Z�ռ�{�
���_[���}Ս�ye*�Y���ypY/ML��gl&��VV�ח��Q�6[�"���7�h��6�dWo[I����-��uj��0|/����٦=Ҳ[�I�٧�^���!2�~�iV��F9�����R�Q0Ə��e��9$]
���q���k���4�h����r �6��O�@X^���rwG�w��-�n�cw�}t���QЋ29��{��;R絥O��p�{������ڸ��麎)pj�Y�����Ō��RM����������yvĥt�;� Ǣ�b�ֽ�,�N���@(�4��S�t�7}��#y|����!sNZ#�X��֮T0�O��qn�M��L[$��޸��6����iも%������]�;��^���]�-��u�N����|��lʴnS�_0c�~�n��B���j���r�Ǡaܺ7~�(���0�v�l��gN���3M���(�5G֜�����̬�
�K�#Y������Y��Ǿ|�����!��W�ѧ��z�o�[K�k���#�-�SvJY��z/�jqߊ+|�\�Vi'�(��@�#�g|��1C(w��5T�"�G@��/�B�W&�sit+4��[m17��4M�;�X�U����Ve.Lem����lz�w!��gյ�ZU�����.��{tL:B�ъ�h���~�x��ke�;I�*
�&.4�����y����G؊�M�r�e��Y�v3�%�F���7S��ы�C�n	��j�i��v���y��Z��c���������u��*��1�4)#s4f�� �w5�h���F����g,�S�޾R�l���}o�]]�^��Y��g��V������,�@ ē[����:��o���;��-����7t��S�k���c��쬟��gO(_@kc7)c�\6)�8>���+<�3b���'ZI#�<��T��2�]VuY]xl�����9�ˑ�1�u˖1���N��/q�9È��%�x�Nv�q7��<��Vo;*k3Z<q|�L���T�w�CAୣ΁KoA[׭Tp��7�eX]E���:��D�N*����%���
��&n�k.��]X�/�j�Ǯ͆��^T����\w�ﱐ��Ҭs�/@ÙQm�.����b��v�L��1��A��J����ZԠ�m�|��#x�Ӻ���;���ʓv^�J��{��kל���m��m��m��nHT�Xu���G�R_A����kv�V�W�.c���"�`0@r�+}\�v7��le(7w��B��n���͸����[˹De��w���G�S�d�l�ҳ;�]#�+��O�
�XD�����s��뻅	0�Rɺ��4�����:kNoZH��2^#2�e*`&�&��B;���÷wk`�T�O&f;�����m�Fkb�;�6 z��;�]k��M���Ͳjv���/��ń��k�l��InRg�n=�v�@�}�o�����tzT�Gz�$�A&�SHEm��v�81�QW�����v�h����L���s\FrW8%�G�zI�s�yߜ�=>�^�a�:VEG�W&�0��j���Ņ@����B:�1�I��%I�M�i������Z\@P�H����Ud�f0ݲN��m�
��fP���&k.�Q�hbJ� i1��I���B�b�E��Ӧ���=3N%Eb�E]��!F*�UQEX�@Y6���]&xL������b�c(�/^7=�.������7��5��[�hJyZ���ʿ�n�/��+{�w,,���Q�_���ެ�7?N9��~���{;������v����I���^F7_��Y}�̆wo��~����|+���?o\�����=hw����d;VO��q�^�V�z{T�Ws��R���a�ߗo��M��K����XP;��f^[����c��VÍ�[�|G_l�ƙ�8��'��W�y?[��{Z�������\����#�3���𬫩k}�2r��,Dh���!�m�7츻\��"m��&�d��1q�6�����^���'G���:�Oy(�t���e���$�Yx�/��/�����~�Vf~Y.�3��k|�y��Id�@������jsߺ_��_W^~�~��%j�S1>镲���MN�o���M7�DJ~������g�L��u���F���	_���?��\�{X�M��VG��K�ꩳ����N�����D�絀ӟ~�?U{]�5��S>F�e�7�߻��_E����ё���m�tL��ߒ�ꯪ�W�?K����x������a�ǳF�b��=�R�$"���^\�m�
��.�w��{̭e�����Ne^j]u�6T�,��(�/)�JD⛲��}U_}W�nX��u�P�4�P�b�I���z�m/�����KK^K���f�;�t���t�ej�3D3V�IH��t�=��\8,䝵��y�u����_5`�ͩ�ݷ��I<���kU� {�n�ݾ��.W������f���IK�3�s.;&�Olb�R���ʅ����*�n#���eE�k������l%�q��n�U���?�rY��'����x�����֥�L�W{gҦ�,�Y�9���FN����Qi<�4��Z�����佼�λzq�w�Eu�%�yw75=�Z���[.��3u�ಫ��_�i���v�h0�`�4��н��|��*��jg�i��-�W���v�iL�JP�.�U���=�>@<I���9o��{���i�8�_Rx�Y3�	��v��o��j�]�g���}I���g~���z�޽���m�Bx��$�I>��@6��O�1�Y!�����!�!�O�sݾ���}w�ށ�I��C�
���P�$醻�B�m���'L�'YBx�f�i� {���9��y�=����� (}�����C���N�)'1$(d�k��d���tϷ�w���w�=��C�Շ�OR|��b{�!�OXI�v}f�q����N�'�$� ��g>��{��Bi��a�$�����g�]YY��C�:>�C��5��;�4��K����Ƽ��� !��c���R����I�n�m՝_�yOߪ�A��WC�=9�X��9pՆ�QK3`�֊�A���T�_�R�u�|��a%a1?:�������:Hv��V�=d��:�����d���C//~�ι����'I=�|ɝ�M2M=�M�q�������B��=d<d�	�!�'I=a������ι���&�<a>�:d�'����v�N����VCi���=N x�75C�6������f��='I>`)�@���l0���x�h��4�ɯ,��O	�v�uՄ����2O�s�,����C�����C5d:d�������C�;�2w�t�ya;Hc%@<מ����5߿s���CL�=O��c$��z�=�2q��bz�x�����&���M��@��ӿ}psY�<��礇��d;a�I=`e��$�x�� q��hx��'�o�$/�oL!XBx��}��n��;�y�N�l�2CiО���@�'l���!�6jä�!5��i�Hx�y�:y��o;�~��>:a����a5��LC�I�I2t�Y>I=`,'l�O,�(M2����ߺ����O��yID�	���1$û!�d��$�H���2T̡��ߟr�?9�[ËsK��1��?�6����:���?'V<�#�Oڗ[�ϕ�})-�����G�����>�ې�-�z���TE	&���}�z��'�t�/l�蛤~2q�tʄ<`��C���0`��XI�/�s�5�����M2m��Y!Y\H�:d>��T�=In�$<Hk�ԓĂ��\�g4����y�zHTI��+���	�!�=H`c=d4�>a�t�d�:OP���8�Xs�����7��ߟz�O�'L�t�&RM�2�� �>d��OXOl��c!������CZ4��޽����=����}�0�$���&yIՓ����݄��B�IN�a�=�m�/|�}�j���󿽐4�ӻ i<��C��I��<d�Hq&:@6�|�Y�$�T�r��r�������;H|��!��Н$��T����a����d�$1�I��t�c!�z�Ѯ���}���}q� z�}��H7d<`,�@�>��t��x�|�m'�� Y!ߜ:�]{�^�<O�O���>��z���Ԑ�0�;a�I�>g�Ci�'Mwd�|I����qw��~{߾���<H$�T�hx��i� |�2��a�@��C�!�C�Ow7OP��ݾ��Uޯ�;?~��^�F�
�F[u��D����6C�qJ��;��&"����&��eN���Y��L8�|�ޠh��vO��!@"��zߝ�=�ޒO���ɛ���t��d�!��	�E�M��4}d�-O�x��OX{ÿ��=��w�COo�&�zj��$��	�=d����C�I�<@:a<`#q<>��Y�מ���7�9���$@���I�x�8��z�x�Y>>�!�Hi���w@�민�7�=����}x�0R�C��d5��d�}B�C��	��
�s��8ɡ2B��LϽҷ���y�O���@���N��$H.���=C�2M�0��$8μ�d�u����{缀i'���d�~�����yI2�:I;CY��d�=CY!M��C���������y�9�6�{� ����C��M�v����g�C�C5a�@�l'�MM�0�_;�����w�~{)��}��a�Aa�I;d� �t�'��l��g�HS(|��'�ѻߧƺ���p'����M!�Rx�uݜB�|�l��=@��q��O���ݰ�ɭgϷ�u�y��>a>�M$��$<t�=a� c4|��@}�4zS��y�~�so%2�;u&V��|��4"�\a7�ݕ(��rG�L��l�vW�w�B%ߎΉ�o^gF��v������|�����$"�>������Ӈ���G�o��8����7�>�V>7�
�jڊ�뺃c�WvQ#�W����&߹ggx�49���_K�rȇ�����2��ڵ�V�Q�<�vC$rn�&�ob+��xm��A�Ai��.��F�c��Q��ALl�Ǔ�fS��\��|��|�"}-:�t�����ϼ��r�ݨ�v����D�����ò<��&�^��x!-�v�f�%����HJ�W���W*C���R�/�ʂ�(Yyw}��%��c�C��ݪg��FS�ᬏ�:���V���$nQ�p�0s͑���U������,�EAd'��:�9+?��?Q��U�.ǻo��)�F�z��CJ�M^ר�yZF���O�C*nj��T
�;o���s��3�x���?TS�����}��-�dd�!��?;���c`��6�]xRʵ�]Ȉ����Z����},��Z�\��Y�hΝ��D�e<� 掕���[G/$m�2J�+���T�u9����<�`�YQ����Y��n�{�Ng�y�W}LK�*���5�lS�ʻ�{grG9�FWư����r�}��8^���I9�>��BE	"�	 Y(� �"�, Y�
Eb�,��"��*�DX�"��(��R�}�5'��h�񮏮*!�ݮ8�^�E��q��F��7�7������Ӌ���(���_뤮�����er���2S��S����F����aP����8�vnR*m>咘v,s��b~�E�z@<�G*3K<����2ԯf|�⺙6<���)��}�t��;Z���b�W�="خ�1�R��"�@�S��t7�[������s�,+�+e��Wx�����/�vdvz{w(�a5|!�H�9��)�܍���.��,�:Q���T6aVx�)�;9����bP7�G
�J�k�K^��H���SK�+�9�X7��`D��y��NL@q��P��w0(���@��0�� �X����G�y���{��û��xԔ���B���<E{�ʠ���j]���R��nԴwm!w����\rG�X����]�7�b�ޠ�ş	BcjOH�O��T����#W�n�Z� m1;Z����i��Tt��0�0���ⴣ�k'�G)k��F��q��$�]�2�[��r�۶�twL�h5����1�&l�ܝ}BC1-E�OT<�v�rqz�
T;3 ��,%ۖ�霺�l�SM��;����(C���s��Ë4v_��E�(r�h4wm��u�į^i�~��m��m��m��k�a�G�=�^{��i��;F��<m�;qp���j�I��w�h��;r��,sV�N.ƨ_'ݘ*�(D�zy6��	N�&6؋��M5��$�ùd����Rǌ=�����pt얃���lB:�kҰ��J��t�Ʃ����E,�10b�k{��fٷN[�:{!�ؖ�t{
V���Tn��YxO\3K�s:����@�wi]$ŝCG.}2�2q�f�0P���m�=�%�M2�060^a�5@�Wq{&]Ѩ�짹N��k켗�[F;L��ٸ�5��_\���.��{�;��{洺�eH�IC`�>L;v6s�j�N�J{\��<�-)j��ޒIi�?������ >��mV�T���������j�6�Z����i!�"�*E%���V
�6�fF��̵"�	m��L�$ě�ul�"�*%b��C1h
(V���&8�P.����)3򁌚`VT
�yf2"(*�*�6ʐ��3Y1�¦���.�*A@��@$>7�����|N{���ã�bM�ۥF��YI�Y%�����.H<]���ﾪ�a��~�]���{��ϥ�/�f�n���{��sS��3�]���3urd�ׯ�L�]"hy�U{����<�lЌN=��U��g���z�m{��ޞ+���X-V��~���ާ�s�b�=Ky�b<���Q�7U�A�#��9r�*��t�_�V��=�k��꒝^�1��YR��3�	�!�Լ���y��>o�N���6�<��5�vr{)W�����S�bEB�e_ �ʉYyk�P�E���b5�����3�t�|��e���nC��{���@��8���_W��UW�L��#Fٿ��j6��2�;]:� �T>Tj����ʆ�\ȇ��}d���.�L���-��^�`�3=��D�6�f�S��Ai���5~1C='���|�Ϊ�����(�/4#<����xwҮ_Fj������D�&��w'��t&�5x�������i�4����������Y��֋BF7����oZk�74���;Nvj>���a��S��o��SQ�)ݗ�YI݌W{Oh���x���?�j�L�h�Pr���N��O��u�}�����ݷ��Db�CF���dsr>�꯾��w�}?��Ч?an�1{ ���:����g:�t��祪9���==�e�c�ѻ�{g۵i��o+w�ܺ�8�ZG2�*�n�l�$췜q�R.�|�X7�2t�6Vx>��ݹ*<tk�al�?P��x����W�eO}l�����u1QG�t��h�r��7�WB).5�Aa�Ê�<~�~g���\�(�ׁG����n"�$��s�){a�ފn��U���?��e�[4{7�6Gw���]�3V��i.Lq�u�7��H��xfoK�6aX��%#2�/:X/��>�ﾯ�]͖�¿�ﹹŚYu�3�*okG�P���K�+6\�;�ܽY����1�'��^��9�_�3���9d{��Xj/,��HhRGy���@D������7(օ�g�}�c<�}�7�j+��`O>��/�=�˴��Ff��j͖+hW�گS}���|�$���osx���\s}�>eem��{�$WPA@��*�Ä]��>*o�c�x��δ����kc�"g��j�ya2��G�^�Ke��*��A0��{�&��y�+��v��m�'=��}��UTsQ��.]c4�Ӎ�nˠ�n{}a!���8e�m�Lw��
[ތ��Ga�U-��6gޗ\�������E���g�Y�z;x����\l�MghY�x����A�
.�8.��o��9�׽���	n��
�4ՠ����������)e�'�>x�x��֮~��:��G^9�6��o5b�����SJ���k6�4>����G��fvf�����q�M���ڲ��OϽ;F�e�a��c
=�;6��8(��ԣ�xI{%�I\��ՅT�ҫ�&��}qIg:�g94�Z1N��K���W���v��r�w�����S�5~�-�g�W6Ae�RW��E�_���W)^CMon�;��>`�۩.�.�� ֆ�<�)�y�}=󭃠��2��	w��9x�%+D�n*��y�� u%k�hQ��j_�I��̹�O���Kl���Jc7�I�S��޶seԳ���42��|%�k��w��h-M�����J���*򗳽��	�v���u|*�3h��9K�J�)�أ!/5a��W�*~>9�W{�Zt��ۛ���x^f�S]k�ᓃ�{8ڶQ"oQI��c�>��  W�
W���_{��S���G!�@��ڶ-��� �[M�t�
��'����#�Qz��t�N^ �P��Vw,���kh��~�r��e��Aο�M~p��]�����g��[5\�?����fۋ{��E�X�RTob��j�����,3��u�vIy[��7�e�ʊeQO)V�"=��܋������T�V�gI[=�GS,ݫ�#V�ƲEOm��G2�A�۷��,[o�</��v�v���cu�uFRD;�s-԰Vqj���n!Iu�ci �D�ŤL!Da駏r��꯾��M�a���(��<����W\�b�8�J�)��y<S�}	��*yap�h}�~�ò��d����5���u
%]��%
�TB���y罱d�$缡�[D9�c�4�	xn��eiCx,��G��t ��P�����_��T=�����N+���x?�F�v3Ϯpm/@"Y�1���0��U�[����1��SumN�	�W��6�-��㾑���uz)a����Z�H[~�y&,sD�-��2�LQ[�X3�+^��#�3;y�Zų�fHd<�G<֡o�}_W�Zy��3��Ἥ��j�Y]^�|^�o�\Y�̨V>���J�n��a����W�$ڝ�=�4�=\}���6� �Wy%�zG]�u>��m�Ө������d�K2��B�)��-��#��M{���a􌘜���[�p#%H%˫��%H.�l���@�Zqz�5VMY�q�%[��ʩp�7�P��8 ��C^E'i���|�QslO����Q�������<O�m������O��aAb���J�[2�gL��3��%:���ku�7C��)aŕ���@�;��������v^/�MW
��/�O��ss��t��Zw+�8����i�c��O�^	Cy�:/��gc~]`� g�S��㼷�b��j(����x�RغĲ���-a��.�`
<Tթ6�e
��%B�Tyᱯ	�t�r^���e�p��k޺4��z2�\;�K���N�"0��A�n��L��c�`&""���>�:+��aj�*蟢^QG�fuP�eu#\�T�S��\�`���{��8���@�������y@��"��;zS��b\���h���;DC���V-���h��.��PN�YNI����<-���qf�뽡ve	6�)م���y^�1O���i]��3������n�f��4v>�\�౉1�#[�8���1m�N�ٸ�INi\�� �%�W�����/i�V6�t����S��ȱr[�ѽҍ�y��:'P�i�zT�p{�h'���A�b�ᕜ�����F�� �.�ީq�զ��Pz�»vV�ѫ5e>37��(=��v�F�]���Y�s�k�O�gs�6v��ʕ�#�-��%���^�G���*T�]a#���h��i�Z�1݂VSvw-��i�2'��hvk����I��4���� K�;�a~7ܥz�c.qm��I$�m��m�wk!�5��m
�@����ׅm�������r(�m�N�f���X�I���b������!���D���݉�s���af�Qd���Ǵ�y}r.�Y����˶:�k�@���r���p�n���ѵ�w@�s&ț���Ȩ'������\1�m*ǃn?��5�7��Zq�vvS�:�r�%�d�����آPD�����'���н��,�]��%������n3�hYl.��x_s̖ә�2|�ܢ�h�)Y�+pa�)����e+��Pq�܃�vL��EM���H�R�&�p��5ܔ����n5�w:ærn��qM�ؖ���RI�w�<�9�O�kL�)E|���X�
:IUgz�V��0n\���%E�B�2T��d~��Ы혁��r�
«�3	�ȸ����)�m��2CT"�[�YLB�
�Tr�PX)R,R������Hv�Y��U���bt����ϙ�6�ۓ�vhٯ	���Kgf<�ui�>�bl��s�u�W�Y��I����t]�,h=��h�*X���]����&����AE�]˹A!�d����[;���f�ЯP���e��I���A�������B����Y+�&w)^^�����<~��E�7�/�zno���]�^���I�L��H�/k�W ��
�몚N[��2N4�P���H�c�������⤬�k����==S��:�v�I]v��3���Ts�Tοm=�Vw�^ w�@ U��<V0��_���x*� �k5�~�ˎ&�Õ�뤺����ӹ�N��y��sS���_V䛛�e��t}�ä\D�8�����MB����}�wJӑ<y>oi8+�����=�:��"x�L���;�TkQ�Qii�!k�/��=x��ɹ�#��G�HȑDWH�gf�}R�t'��y�Zx<M){Q��o�/����X��iM�Pzס��<�"����/k&��t!�v���qj���PG�}��ڼw�+g1|L�	�^�/�)�9:�,\:u�l�f`�֛�Q;S�������s��#�:��{3N%�yw����)�F���٩������u�3Y����?}_}��g�Yc�˲�Gz�C���
qkrI� 7����xm��V�q_�;���)K̩�F����-�~�͋��"g��'����អ��s��H��;*��r��$v�m1�i
k�G^�1>��K�e_�Y7��̊C��=������R���{�q)��o� �u����!����|ԥ�.9��6��}�f�倓e;��I\TV������(!��Q�n�.�(�/{k��B�7��!��'�	u:�k�ߜ�xdk3��8��5�X�Z9{�����W�ۍd��ij䝡����w6Ӟ]޻��_�T��kܽ��%�9��+y|�]Ii�O0Vf$��������@���u��+�pN���� b�ŗ�+ަ9خ�>�ݳ� sR�{�|.���5�@�.�j�[�J��\�^	EuX�^��$������Ю�ߢ��5[�3@n�v� �V�{���=Tf���l��͍.��r����I�3�����'��!��� �X���l���g���r\��V*}}Sa���S���r���{L�;ź(���l�^��4u��v׀�a|���O1v��"X�{������ͅ���｜�%&��W[��|�0���D��_�b��Һ�g?{��`�b�C�k��ѣ��Ю>ۿ��b�^?\oT���hz��T��� �Z��
��c]Z�o����C�.��F��e]
@��\�v���ތCA���t}u���))t5}.�.�	��`tU8Mqӡ;!���&k�tW�e
�ˮ����)н�=]�۞ڡu�����~>b��N���䟧�#T^�gQ���]q�g<G�d����}��ѯ�?{�pg��ll?!M+�!Kna��}�M_xU����>��a��b��뗁�����m���v��LZ�f�R�z�L�ߒ��'���͙+�VL��Zu�7'9|���2���f�|�l�Ŵ�]���}_^NI'���k+��T�t>�=�$�Cx����Æ��{��Fx< ��MQ��5B�wm�W���w����ˮ���"5�C�^�5f ��,\�r�o�f�Iγ��X�R�֊���y,
� +�#�Z��L��zVp5�XB�E.(QF�u8�\{�\�Ͻ�7u�i�?A�z���	Ƙ�~�UpE���+ڛx6����C�ZhC~��Y�")�8fL�V_,^񩏬�ݽ9��ǉ����7xv��=�z�d���C�������_¨�8es(1^�/��n��+ڎЃG�ڮ�*��*��hЬ��x)~H�K�[B�ӆ��KXm��S�k�x#N��GR��oW5J�����-�ҫ$:(w.䦾���*�9X��'n��q������I��8�����6S�������hT���ϰ�.meAQ�H��ׄBC���u���眽�=�`r�z�4>γ�V�������3@ \ּ��l�o� �
�i��v���W�cG{}ޞ�|>3WZX��5�X�Ή�t��+My��[fC]rаEh^:M/0�W��ۭ;:yj^��^4=�^၌'�`�X�kVy|��vs^���م��w���U�	��B�)+��9TU���H�*c�Ҽ��_uQ�*�ơ�r�0�Q��*U��򉁆�¸K�]8<�
�%���A۩�C��� RMq�	9�\#�>�J����^�\V���BVLɺ�R�p���alcv*�Y ���S��׀�W-}RM�����vn�<� �u��I���^�< �k���ЁV%i�����P�(x� ٪�v��nE6s�Y��x�@�g��
7-
X~�R
��<��}l��������i��yޱ��w��<`����^�>nˬ#^c6��R���+�=/�D�+q��5�o�]e��M�:]�1�uH�zt���k�̽�"�^4)H�t4u�f��F�6&����� Y�iB��+C�/���r;�:{��K�0V��UwY!�� �����.�S����^�4�,���`B��V��=�}=똁���Jeu,�;���lJ�������nx�7�� ���u��qi2n��R�
�6V�m��y�Ӿ府UW�glrOuw������� Oƴ<�
����=�͝�����U�) +�up�0o��ŏ��e��2�'{��׬1�3^F�ƺ�M]t�)0?CG׽|5��h��j-�K��48 w� )�<)��"�7�۾���|��[>�X��Ƹ0M�{��EXw�w��|���]`��(׊|iB����\|MP�0�����%3�
=�N�H� }\/���c;w������uu��4#@�̪@eu������Pk���m	�A�G�6�p֌�w]o�B!���^���`��V6��.�b�5Z�4�E��ַ�k�~X���i����= t�h�ꝍ�ʘa7���f�j�9Rd�@r�ᝲ�=���]�T%�ޜ�9��}�|7c�'��_�����K�4���>^gA4ga�S���y3=�G�HZj��i��h��;�Uк5RD�=�w?3 ҄G�iBz\�!Sm~r��	?{{�h��ׄFm�L�R[���k;!V���K���,S�f��n�Я
��}�t��s]�墬.���j��z�b )x����1�>.�!���'}�i��Q��4u#�	@P���ub(y���C���z<?jx��f��H֎G~4i۰��_�f��y����g�C���)lѤU�A!�zw�u���f�w{�&r͞���y��<��]�'��<��3��4�]�^v�Q�Om�`���'��TZ�&n'���o)W`�v�9@����^p8[�����0]M��wh2'ԩtX'E2�%����u��)V��;cE��N�������Ҳ�J�oV}:/�憲,G��x�r�E%�z��AS-p�)<�7\=���s� m��r]L����T[�S4R�.A:v��DD�K1��u�Zf�T/�� �tj��?]�D�=��b��nQ�z1<o��Š\V1�ݜ/:�s���y�.�L]5���1��6Kۜ,�s�N+��@��w}P��љW�L�f9=�����J��֥s������k���Dua�د�8G�ܷ��xzgtvW.=��wu:�͵�C0�ʤ�/��N���9Ŷ�m��m��m�ת���{�q7�S�l��n��ѩs�-�pä�fHl�
:21�Ǯ>�KnV#�.�k��C��gƤ1n�E&�8]$��������U�'���ͻ��g!���W�7Q���_-ɻ	�L���^�M��`2n�nE�i�r㌌��)O��Z�$Z�i�/Z���g�`g�p��th)v�$9і�]���zWk��c
پ�,$� yܡ����tД3�ǒ,��љ�;��N��消u7�%]�8Ӹ�܃-l	��Z�]:�2r��޽<kWs��W/"�Y�5�J��HyjB����p��yv�:�9�L�͹ѿ�b�(�/�e>F8�
��-��i����}G�`VB�Ƴ����$�j�]eTQ���"�2�f�q+��.�����2ٖ�AJ��1
�7V����0�������Ӊ���VVVq�i�D�M�������br�ݨ����X�Z[�ɦ4�0(˫ ��ed��^�T6¤���,1]2�7��l�GT��
Ő�
������i�	�Ƕi1�]�2��7i���1�*T����k����֮�2�L�Se1�v��[���~�����\��ξ��RΟ`A��Ś5�n���7Zhx߽u��2!���\����3���8R"�b�T���J]ݺ�B٭
��}�oOL���
�M^@�M�+�W��]H�y����}��K.���]
���4�q�1Y��h,k޿F�yމ�������g�4��+}1,�n8�}�uY��[t�"�x�R0Fp1��ۧ׋���z{�J'���� ��t��P��b?c�z�z5��|0L:,M+�4��h���������Dv���S���ץ���E�tl�G���my�fr�GUp��q�z�e��X���[��I*>4�8+�{w%(aT~x~3(l�o��u2�ʷ^���#1b�Ν��t	Yq��ƨV<�k�'��h|��N�j󠵄���W�|#����:&[�T��,n��� @<9�fL>������^���lX�ʖ�
�e�o��#�>k��yؙ��b���_eՋ�X1`�D	��ފ��AL;�WV0d,/�]b\p�$��}6y��|+�@A
C�����N�ƚ��0r��S�:9�^D
��B�+Bg�wtl�4W����ė��������T�:�ig�ѺO�s4
ƅ���Ӎ���k5)Ц5�r���s��~���:=,���Z+�`�j�s�a���È�H1�ɥ^+u��}t�� ��	e��wFװ�[�O.� ��1�w_WZ�V�쭺���|6�����/[M����l���q� � ۧP�͹���<Mԍ�5���u���U}UB�WG�8<>6^�C���9]uc�﯇���X����{���Q��[��
�M�����ح������E	�4�p׆��6��h`� ��rͬ!�Ӝ�����]^�L�*�z��PR	�Lh�;t����zq�G�芙�Oƴ<��5��JIw������|10�F����СJ���!X˒�/cY�G�^�phc�0(p�1^�wt�W�ӍI���
{З|�/Kb�9_�6XgY�a�~m�}�O.�_�Ո+�K�>5�@��hw���f�g����{MOc���V���5¯���M�@k�����8�T櫠yV��:[��˱�f����1;���W$����yy����W$��'5��d;G�K�7�{?}_}E�����_���B�\�(б�F)��Z�m�YK�ܖ{
��
.T�o֟ Ժ�pT*�}ii��(����ǃdP�*7.�9f�`��;�����Qs��z�>����EU�w��x�iaCxEhu��ɮ*D�T��
l׼qr��,u#��{N���W���n�/|�]�������[�W� �4���額?	^�f���T��p��m������X�?z�����}���i�SG�+�y��^����g;B��&�U�\�"�+�#�],.��Q��ޙYL�9�=�8^�{��ʯq��� D��!U�����m1��H�y��݄�l�xNæ8j�3f��Pb�]]`�Tm
�9�%�0����ua�Qz��]��͢f����T����|35s�ǫ?R�3Y�ΗVMJ���8p�>Q��������<$�?��2��{Ɲ�b���Ȋ�����:A���?],V|_h ��n��P�:S�<pz����0����c������_���˾~�@U���
�ˮΰ���4t��jN^�-4���b�M��Kyu��V2Ib��E�g����8�B)���M!���
8i<So��k�0��n]^�T�*��3���CHg��W�f���i.m�A�/-��� ;?p����v���n�#��yb��Z3%R�`�k��3��0&��<����U㞮���MS'׊�0f|s�	��I\��K�n�Q����������������W&�Nwj�����$n�����=?��ߓy��<z`W�2����Ë�%��W�k�g�&o�h�����m�c��0}��ښc}��^k(VC�|>8��q�A٢�~�^%�I�f˪�GJe
�;b�F��>��������r|���m�M>'�+(T�w��z ��w?x�~�A��}oc ������&q�Uǯ�[X
bxӼ쐁W��Z>U�л4D�B��弍\��Rǵ�����+���~�&S�ypWi�0��zzm�q��mBE
�~Iъ��D;�<�6>����j +���کX��&����-��f�~�ݢ(���k5��̙ˉ���[���S����I��}kFk��Nj�]���t��e���r���y9Ko�UWض5'��a ��]҂�� G@�,��9f�z����>���^G�(q���vS	�`_�����@.z����d͌~5w+�`�\=���g��Sɞ���yj�`��i���Z����EU�߶�Vy����ð�p�U��5���Ʒ�>Ǉ�⃞���j?H�i��yS5�ׂ�Q�������eu���jw���z�k����x�����A
 �KҮ�F.��d [0{M{���τ�z��FB��{+��l����#�**{&p�=,0�e�Ǽ�W\ej9=.G%����(L�<$Q.��|}R4K�{ƼP��ͭ'������X�H\ft��[*�e_Gvo24v"Mw'��l���J�њ�hl���Lk�,��=�8����'?�_}C3WG�]��uՒ����b�4P�)���Va@ݜPݵ�ٴCG����-�@�pa5.�����ދ��d��Ċ��,��5�X��i�����,P�7�y�'����i�c���5"4ġG.����OH
�\������&��Vb�тѧd�3+�����!���5�L^���.��O� eз˂ ��i�=����(R�/���\	�����zZ�NدK�<���g;�ޛ^����`��FU��W��WY.�#�p��jM���2�Tf��>r��ia�}��Ag��m�D�l({�;�v3MW��P���[WWXwĻ�D/;���I�v˜(l�Z9,�o�m�Q�b�ͨ�_�^kiNU�V�e{�\	����d70�6�,��sr~����<�q�U�Ő~���t0{Kr�����v��˭��a4�{��
��#MA�Pi�*�X��;~�^$T�a�8Se��X]=�=�__�w.��R.>��Ui��|(ρ��/̪�۾�I۩�K�j��a�O	|��DDte��<�*V�m��8�'�ر�~>4��=�N�1E5��0��o��)�G��lxU�,*��PB�٧e���zX��S��M0Y4���Ձ����}�%��D��yʗ7;Y���P�a���VH���,�c��Ї�5��=�4^lo�i�5 A^�8{���ۨ<)V;$�y_>��zw�ñiV���L����h淺&++gYZ\���7���ޞ���s��RS0�u R�+�}݋w�������ټ��P�e���x�I<8��ˤ,x �|ÿG�8�y��z��\����⡥H�.�̩�U�'�eW~,@G�8'�܈���|p6~�I~ĺM�6G30�jz_�v]�g��W뱃�� +�4TŻ����~��wpU� ��Q�kC�n�|�������i�P#XA]���֞h�5�G'��G�����������^���Yz]�����`炬�k�y����]p�|S<�&X�Ehp�tȃD=����{�|&�ۂ�|��T�~�kC�[%_W�sJ<�i��Em_�Qv�����a�$(X�����~\���R� �ӓV�}@���Y��!��J�Y���r��;�Vr����j�.)�2f�y�飛hhSD6P�Ꝗo��3�'i��r,�`�]�R��h�oW��C��
CZ��+�W���j�^�o��i0p퇤'�����l��\{��V0�u���٢�7�dGssM���a��u��P��W�nVM�P��{(3Thc`���z��[�Ur�Z�x��ߧq��c#;D"Р2D�0u
�C��XZ5�����CM���P�ѐ'��V��%IƔ�ݻ��c%-��^Ce�y�[]N���q�6Z��B�\aޣq)f���̵w��޼1Y:�#�橃��C�.������k��Y��7���@�r?k�Im��m��m�����\�¸���h�\)��Kx���C	>�jE1�W�_[�W�GO�fk`�����+�9�tv���B[}���p�I��n�����{ ՝��r���(�n^u��xNu>J��O�Y�&���ոp�}�a�٤.��N9�a=����8����ؖ?B�@����z(gT|j�5ʠ�M���m-t�y��jv�t��\���U�ח\߶v`�.mE�[�W�R7�]�|�|I�j�Ͱ�f֮؎ؔ�u����nk�拭?�Ŷ����y���y��hsX�}�hә::���xM�K�r��X�ZgU�	ù-����Y�;�T�N�I$��`P�+�
CeE<f i�jb(����^[&�)+EUY�Lq1T�a���,Б���� ���dQ��W�`��clU�&�TG,��쮙&�XbbAB�8cE+1���J�DT
əAH(��&ݡ��5Q��w�!��*��՚j6�Z1Y��
��b`�#X\��&���YSI�׭�����zo������C:���DN���3sV[����S����}N�/}
������*끮����Ab�}ᬯ<���h�W48�>���WF��ax�]wm�~�7�x�9O{3���lי�0������^�WYKS����!�'�4}`W��Ŋ�
Іy�&��������S�o�Z ciт�%
c嵷�p�G�w��r�1X>�g8�a��W� ~�
�PR��绞x�S��B�^_]��B}u²�H���84cݞ����P�,Lw�p������W�
Xj�Y;���r�g/9�"�
|l�5�(��x�z�xb��G��=`�u�O/�क़P"�������!�x��P4}%�	�꽲�����k҇Ss��W������*U�0Ꙉ��i�h�ܩq9���cW̧�[�������_
��y|*���ٮ�������P߅=s�Y�Ϝ���<*�X�Zjx�0���s�*C��u��ucA�H]j���Jf]hN��\U��[Y�3�@�.�X4Y~5�2�ׂ�x��YY��b������<��L
W�>5!��������щ���l_�HX� �WR{�������pוx꺱AYR�̰\�3w���>�q��kè^DX��A}WV���7����I|��b��ź0!M)OW��RI�*�-3�L�Ќ4�o֟ ԺO���m񇼺��!k���j�C����n0�/���<Maɵd�%lR�%.��9'j�\�hվ��Y\��슼�;�~����=L́�	�	A�¼j�i��Y�Eiݜ���^�ux� }ᰱ|P�8B5�X�6��VM|$q̩�(gyk��8�ԥ�R�')˫��X�k��o���}��ԝ��{�����BL�]v��ջ�&����8�����وl,��=��5�߶^�O�)WJ�~��j�<�yG;o	�
^5�
�Ȍ5z[	�i�����Qv(+F��AˮჍ��2��O՞��)�lh��I�*��]V��[,3B�@��O����yw�c���5^9t�o��x�z�~���%C��aEt�S�
��G�_��Sa�kƝѦ(�Wr{�:$�Y�umk�b�s�N�o2���Y;Z��X�V�����6�����+Eo���!�H�Sv*���۝���~�7:��k;�|`�.��1ȉ�֟�W��P�|.���*x]]au��>ʅ��bg+���觼�V���hA�"���$G�i��~��GT}���t�=���J}��CD%��Y�s&�#V��#�$�4K�/Ŋ�D3tME�� �f�k�z���4v�4����*��(1�WZ���6�fx��<�9>������D�*_�; �G�G���~O{�x�����F�)z�f�����5��r]=mdپ�M��:3Mn,�'<h�]!�P��8M+��%�?M�w��O'�⬊cM�F��x�<�(^Q���Bz&>5��T P����	�s��wK7k5ĝ���\�5���<O��=�w<wX����b>�D\|��UƷ��ssS��c\����>m[��⛺���^���EG�E��� ίyQ�LQ��L�4��h~6���6q;�x�Rw��#D�w^L,<>G�+A��ۿ�2e��~�X<L S��A����^x�#�mqИ^���n�,}ҫ��ac��5�~4�Тk;(���s9�#��R>�����p(|� �ʳ���ㆹ��/w�'VW+Ƨ������n���^��.�w���xב�:�� )��x�X8y����u��~:4T	*]���|���~����vOOu�"���!X>�0�[_�.�ŀ�~�}G��Y0�}k�r�EsB�ͽ%gX��vk"6�y�{-u+��5�ڝ;*@v�Uʑ���;�W*;���$��꠱=�5���-�w����$�
�^8 �D�枞��xN5�h�h��s�^ŋͺ��K�� en)~4�x �{
S�^Ƽ:
��������O�G�����[�B�gW^�㇮�jϔ�N�=�n�
�� i±������_������n�N��(�Q�l�zXZj]K�9�,T��]�쏣�DM5����1vib�_��O�hyo|�o�g^鳺��J� G�e<��A��_B�x�O��{��Ǖ���4n�p�`PB�)��ѧ�^Q{w�:CF��tG2ǰ�� # -�����v�9�9����)^��V+eYAkV5�XM�oM�ϸ�c\K�oL�����5d�Ǥ�794y`��67����k�� /����1|H�f�=f�B��L�~�3���w��7&�e
��7�����Wx�1[S�1B+O$��1�}��WX'�Q?b-h}]+��^\>R���2P��� � C��5���_/2ed;�.�b�����c��{˴xR��eu����m^�:�V��{�
��f�x� }��*���zsz��{��\޺ۥn�8i�E���C���!S�d֧������`Yu6�uO���R����$�y�^Cޫ	Ƈ�Q�[P�.�И����Ͻ�ǩz�cޞd_�AO��i
�;��GV�A�Xu1V�녯��xh�ˈ�7h>�v������J�WX�iDx��Éӵ�w-3��\�rEc�Ƥӏ�V�VA}�쟨}�ޏ��~Ϫbp�|lp� �����}l���+a7�$�WOexr+]�t�C��h^�i�#Oh�h�{���^��׎��Qˮ��ká�.��"#�	A
���'ZC���Gև���yƢ�q_�APWy_�D�E��u4�9F�;����\|
��,]�cr߫VG�ʬh�B�xA�����4�?x}�
D7�����i�Y�}��;��v)y��ZG�Ӻ��]f�/nVH=�Px���8x�.�(����KX�k�����wy.�}�|ǅ TM �ߺ���m>��w7^G%h����c�j#��^�( ġS���ۑb4f/{�]��糱&��qV3L���J�$�WS�cR�b;��VK�_)��L��e�1w�����p�����3L)9����մ+!���oG�~�N�v~���y?�_��Eg�[�$���/V]�d��B]���W�L�h7hp�m�S4U�O�4�Uj9㽆�_jK��J�<>�|9��e
���a +�p��Z������F
�޶CY������6.��$��t�k<�Ѻ����'��*�Q�Lҷl_���@���m���Z�6B5�H��L@���޺�оձބ}�� )o�F�2�����A�+V;<�׳��U�e�/�17��a5z
���W��;������.�@ƳDpև�)��oG�q�mz��Y����5�wwS��ۼ��S�ęcy�d1X�V_n�s���nQW>z��N��:��ɭt�)�r�\���/�q�gî�K�v�~6-p�PȡV��:����Ӗ�t��8��X�&���X���Jg������wF��>B� �tt�á J��l��I�Z�̿(��_Y��
]?�p	}��)��^ވ
���@q��:=,�����iƼ��YC��xj,Fs�ัy���<)^$󽞋�X"5�P ���=���zk�|]�9�N_�ӱ4o�<�����A��	��_K��XB���TE�����$���"���<X��px)׮�������"�Cٷ�I�/5��Bj/\��G�E��a3૥�7_{S���έ4��n�{{���.�O�@p��&���T��uجޙ��Ir��-��՗P�r�
㵝��HWv�a�aF���t��}��n+��sp>{>���0����p���\3���I�̣Ť�*��wo8 ��N�NtƜ:�b���4b���V���{�����n杧b\�2azFj��@z�֦�h��M�;�T|�5��������sy�;Z��D��Q��k�� �b�K��N��\{ �0��`ٽ'b�� ^p��=m���l ���侳�U�It�t��Q}��C��a���6��K|��<�n��w������s>db����+l���9�����ե�R���s(�t-o2�&�m��m��m��^9���d�³cj�)���K��%��x�Ep�� �J�mП:Z����Գ�ٲ�3x��L�Wt@�4��4�b��]`���9��u�^J���:�Nb=V7�W^��.����ɛN�Yr�h�v�	�[����È�-��y.Z{uVGz��S�	b霮�R���.�qm���v�yڝ�@������n��f��ֹ:#����cBZ��wn��:V�V��R8eI�/:eV*�t�*Ue��3�st�T]\�)�b=�z�O�y� +V���6U�1�q47nvܼ�����Q��T��<�8�]���jƌ�l��q��.K��՚m���]�o� ����c��ъ�mA`��p�TW�*��b��i4�e�)wf
�@��,TQ)Z��{h�DĪœHS�T�Z6��]fd���y�04�e����B��[m�a�34�,lQEƢ�lU�-F1oM`�FV
9B�v�[*��kE�pJֲ�	P+X��uB�K5Zʂ�QD�,����arᔨ�ݨ���^���cN�A7�%�;OoÛ�=���Gq��cܥ��I9�(gj������5����+^,�`y����C	:���?;�=����C,���C�p@
�0ׄ˃�	<=�{�{��Ka`��R�6�!�4Ś(U׍9=�W��JZ|MAxtzK������� �98��]$���\`�8��k|i�z�!��h���SS��:���
��4�;����lU��bC�'ww/[��4�&�����˼�߶i{�N����c�}���F�5�Q#��}�G�B�pCR��u�Z|h�;�*�N{7�P8p{�H^�<,PE��Pb�j�i�d� ��^�͸k�Ί�5����r>�]�e>�}�yg*duj�#$n���>[�Y ��^s��h�&�Z��*u��o�A�͵�y-���*P2��]���e��d�~���m˞����zpN��ڷB�4Ţ�"𠋃�arNI�<~�>��������M/MW��P�&�X��V'�n���wB�Q�ll,(NW��pe=�ֿ�<�~�X_��������`V�����F�	g8e�8���݅ǆ���{��6.���vĳJˠ�d�/��PQ������R���a�x �.E͢{{'��]�z�O���U�X���J�P�K�>���{�M�'�bǨ�C�R��P�`�x�a���x��w�D�5�Sw�P��^�<*�c�R Gi�}'V�4RC��]O��[da�;��~�>��>@�"�֪�n�_	z�imW���.�C{�^a���@�2��g���L�IjΈEK����֢mN�Y��8z�t��蹪s_�Ặ)=��p�� ?W���0��c�WWot�~�P��i�R�C>�u��_�AZ0{I�B�f��=�zHk��B��Y'�C�*��V����ɔ嶜�L�������S��o�
��A��W�����zxSÜp��¨��ōV���װ�j#��/(��d��^�?Z���Wu��
�D��q;�u뱀ǵ���w'��Ñ��
���� ���]��ÃJ{}��yDLQ{�N]�	^Vǡ��o�8+�у(���c�u��̙�E<��
�*��؆CY���8������wt�䧧��O#D@���x"�ThSg�K�+��}����t�xs�A#�<p�"���AWI�����ˈ1t�9f3����kM����3���2�5�\�#�a����X-��˧%ߨ��
�mK��(�4/��p��`��4֊���w��g�'�q�KMod�<X�_�������͡��7�=���������1~4�;���~�*���D~5P�n]X�X�~�.�h}b�n�zׁ��O-M�=�C�"���<�iÐ� ]"�]#�-�{7��w�C^�i���D�21t�v+����Vf���~X=���4A�����A�!.�*�(��w�w+4���8<(�`��_��a��|~.���'��
�"5� ./g����X����4,�{�8U�YBW�xA�,Fs�Q5�uŋ�̭WC�Me(�O*:���U�Jk`�q�۾�`/?=���(���&�h|3�j��;��LJ�Rmy���4��E��{���<K��������[t��5������+~\Xk�K�~�&��O��-��(�{�(y�]�U�X�V��]
��)�ΰ�������C����V��pW
Ǉ����4+��w��+��=��4x|��<y�X����S��G�%��ɷ��f��4���pB�"�1`<,1=u����KU������`@�A�P�+� Pf�9�����(�Z>�5����\i�A
��~ �^R��k��5�O�+*ʆo�K�ń ��z�w�jnh� /e�c�q"�kְ�Yb��wq5=;�w�}������`��4�;�
���lU��)'�3�Y�z��#o�Q�V(�o��%p�C����}ս�K�����+��c��Z�ϕ�Ա�E�{��}�ۂN��Q���P�G�p|o~���m>�4=~�*{Ȏ�o{ӆ���� Hb>�G�t�� �5��z�@y�0��"�ΰ%��i�jZ������CO�Z�NدK��C^����\P�8^W��v�/8�z��u�h,���L�ʼi��:��¼+G��a��W��󿮇�^���L<e�?i!*f��}/u�C;�;�^����F��#Ɔ����<m�ݔ����������4������i
�ֈ(՞D=Y�]�|��&z�����S�*�C�+Ë�%�Y�ϴzE���}|g�kC�[uHR�8(C����e�}�d1�i��`�p�r����x�P��Ǎ�KcW��[��t�6�=[ەhn��}%�/rʴdx�{./չ"�{i����~�p��ז��
�utM*��q��7/�tO��Pbo��A e?�౼~0��}�-�+��׽]�X(�4t�E
�Ӱ������6����|�#Ⴧ����
|]
�6��?oLV�ogc�{�J��G��<>``��4|i&�����f�ȇ�hx���j��%����)u��M�>�:����d��B��e������Q�+^k����U�p���W��XxQ�=AK�L�#3�W�zب/H���"�8���?4�
aB���&�jH��=�W��׈����j��Jۥ�猖��S��RC�H��v�#���HKս��wS9�w�xj������EI(���Ǜ�9�|�Z�W�wi�@�l/��i�M0�G��u�ux|.�CI��B�V�	���'����wW[.�+��q�P���Т=��Ӕ��2����«��^5�q+��g&������s�tOeѳ �z]V
:S.��׾�(�����(
С�wP�ۗW��4���A,��dx�^RU�Zpi?p� 0f��`2�;����œ�������=�+��A�ЬE]@k��X�m�eB�3d��Y��
�~><�ڬ��l����W�r�.�iw��R���Y��.5p�5 !Wε��^��I�p�"ѧp��4e�Ph��*�yg�H�G�v�nڱ����6o�wc�<w30z�ז���^Yk��i)���U�/�Z���u��KZ��yI"6&����V[����y�Mց_��(M+7���^�ư@á���wZ���%��U��U�*a��
�����vO'�kԊ+x^�Ѡ�3�W��!z��{3�ӓii�+�X^˃� �Qbe;�9Dׅ�ck��7]�{��mhb�B
�Q`1�m�f��/�x{o����}��WF��0MS8�<�3�E��~�yz����Cō�W�YZXxV�5�c5��B�~nPz�L��(�M/g�
�@�Wi����R�t�N^��G׾>�\���C�)�+�X)�]���y��1�t��w�y�{��@�0ಉ�{5z8�����ޣ�ך�
��ku~�V�q:���/6^�����2�ϳm4ud׮�Qe���_9i/5�Z�x��{�~E3�mq�ʹ;�Ƶ�3\J�)��y�y��zS"��4�@�XP���B�XlxT���]5���� r��&��r�A��ka���W�Nǽ���}^6@������EXvT5�\2��Im��8�K���EͶ=���
�4k��yw���}b���r�)���^!n��G�,ˮ�P;q�M�%WR����UE�oCŷ@B�����l�-��mh6�*���`5���'�ٜ��ｆ�QL��]љ��4cնU��t��*���l�J�Y�?n�G1�j<����Q�uF�S���V�/9ŲsO=����P�'�:��.̹!�u�K����c����Z�2kF��P��1�6�{-˝���-6���z�M�4 3T&�P�gQ�1@�o*��e�N�e:y[ֳ)}��}�*I�X�j�:���,�Z��[�[�����C:���Z)�؏vɇsz8Q�������8�4宫�����#�a���n��^J%�"��mr����6��;�^�8���2��;���u�?D��FPw��yW�%�]y��{:��]6��G*i�%�ҩ#k�wc��`�2��P� ��v����"�3�������[w��Ai��fgj���|:�WP7�I9�$�6�m��m���u����ֱV z��ꅓ�jSqi(e�3n���wO�=���;3���Ғ�iU�GSx���5��
1�6�*f�y�BP�l��.u�W�|73KKK�[Υ-JJl��*�U�x� _�Sz�VgMc5 muZ���Si�N�Jb�����3'<#���'�.I�sv�drVgNT�ݭ�7+cv��V�WN������2SY�
���Unw+`ܤk:؜f��&�+w%��Q�)Y��5d�l#J��U��{ejeC���lP�+ĝs��z`X7�L8s/|��՜�k�u�M�"���k&q�{w�\����$Ζ�\:�w���t�I'�JQ �> x8�5��-VQb"��KJ*�D��ZUt�C��UUU݅�i3,X(�1�*�R�娬\��**�TEf��mj(����-�[t�(TZ�LrҢ&XU̦6ѵeE��PuM0ƥ�s,��n�a���AEUJ�eEEDD�L�EaYwF�1�A�,U��VdM�����mm�DQQD=���oMq�\q�F�Q�e*�%"�(��ejWHc�[�E2�`�+i�QAT�+�68!��L���QG̺�S*Q�b�Qj��Xt�ch�Ȱ|w�Љ��u^>{�;���5VP�@pj��u��s��=u'?�ܜ����p�'�^=��i��0�٤��`:D�s������{z>�*Mf7θ��(vq��I�BOt�3x���=5��+�Ư��^���G?l���5�8I�=N�&��c�1`�y{=�G]}�-��v���1�v5=��D�f�S�+yX�]#{�ґ�͹���O�܏�I�wW��������۽�p5��N]:��dGu��~�-��轥Si��b�� �W��x�z�������G)iH�Ҹ�`,C%Ԙ��4�;��3y�ϩM�+C3]<ǭ���j�b-����5�߫ٳ�g2�[cYRL��b�nK̜&����f�{��w1T�����f��1K��?����/Q���\b9���ËA��s�s�"=��<�$�>�io�MZׇ��~#�[vl�YG�����+���u���|����B�:t��l�
ºp2��q��{Pp2�z�3=f��lv�Փ�Mo�t�M*����q�:�q�1����^��$�ή�V�jTa��W��@2�.T�6uɰ���az^e�e_S�.�ă&>�m58]ci:޹������`��{Î�O��9pM�؞����4i���S��eÝ�ޑl�[�D��Z[K�^�����G`���\	{i��
ī~��R�9	|�vzH6��G��4��f�y�C�Ml��a�/�^��֍Y�p	U�N�Δ�r��c�X��.`B�3
�q��z���$n(��*����\w�9Z�k`��oX���_*rӊ����-�л��'��}���8-������_���c�x��"�sJ�U��y�9���Qޭ\��>�B=�1M����CR���s�rf�F
�[j�}RG?+=&+�VV�v�i�s�:[����e~�\H���x�on�^N��k���՝��^t��u��x�K���4�Զ�9���������3����埨�qO�r�ԃ8;��w�����y�-?�о�;t�O(l�h^����[Pe)���Yˢ��p��*K�+���(`/y�9�K��t�V���s�Ŕfܽ�IW��^��j�����d�ǅ��b�]
�q�ٺ������F߬��^��y��)r�Mi�eo<��u�9B��j�<���w��-�z����s����U����:*�gj{.%��n')Z;T775a�u�[K��í�(��:]��g_C��:�j��'άj��\%^.]�y�<^�����ni�{��y����z�Qc�q���.��0f���W��նk}��}�3&�G�e���|Y{��-��S�=�`<
VU�`vi�s�ȃ��� 8&���Y^��(����+ w�5nMH�{F���=�����H�]ս	�6?J!�݃�չ���%#��Ȓ]���B^����;a���V��&�����[��MYdVs|��U���|�L�j-����Q��/�շ~�ǣbqL�HR������/� @���Ϯ��Ke1J�pVԳ�W�95�,�)��I��v�-�VC�$����*�6�{��/iM�m@0��7�Ks����߮/Y��sU�La.�;��T���
�v��O��*�=vD{Ȓ��h�^�>�Z��}�l�=�p�����9��ϳ�N�
>CR�Ïre�No9����˜#ͽ�8/Sol�l���ի쨕��a���V�U¯W�a�w��a��r&c���U��1�����.֩�������6$���?�7�9U�k�W��mu VC;��:���j�G�/�����#����o}$���V/hj��,���/���\
�'�C��;����v�[�@ɾ�lp��Չ!pR6����G��ǣ���,��[���j��,�:4.d���c��P����S���>\Z�L_&�|kz�5�r�w�#��53��5��m��u���.��0��mL��#=F�%�#��c8������:��MLDo��ె��^�o�nK��P�L����7b�2[���䔾/z�V��RA���dz��խ)��߿+����^*���DsI�Dߗ1w�`Ȭ���(�0��X�7f�眜�4�gG��EA+���rA�9M;=�|�r����<z��=��ܙ/^���`���9A���[�lG�)���\�6��V��j����s��i�Kl{;�A;=uIJ��l���_��M)x���s׈���\�N0�J���q[��ߝ(fm��Ӵ���q�u�bn�W�����g�u%>�^���]���W~�p�7v�����5��l@hm��+RyA���ٽX�R���������dB:��gR�)�ί�r/��\�CJ���#��\�i���8��|\�0(O�enᕎ����rD�g��*�p��K�sG&8�M�����J�Rf�%���Xn��$��Ǌk�5�kUti]QF�*+�^�U�,���ǔ77#\�*�\ �a�<��jNJ�:�3�1��^���˝�:}y9�1\s�W<�W�2��7�!q�#��Ez��� "�̞�{�8�>�缤G盆�=&4���U�F��Ip��H�u,�8�g�\��	�JWB�w+�x���L>�Y_^�f��]4:':WM��oi�}�SP����I<����Y�诔���\Wh+�bޞ^w���v:r��P���{�K��uؤE�W���/Ν�Ŭ{]r~�@��&��!�^q��J�c�~���8��<6S��o>C��t)�H��W�Њs��a��K��f�4�uz`[Jo���5L�5	�ԓ�5Ca��.,���%��m��$(��������m_ٚ�b��֣M~[~��A�$�cי2��x��J�i�n`��t߄ݠ�i�A���5F˺�7t-H����+9�]Բ�Rk��Y�B�T�6��Cs�t�B�Y�Q�xE6��->��f�囻p�ǃ�k���s��(���ϥh��+(մ�]���%��'�Z�&�D���]�w3r�[��ät��u�R:	���fdn�_[�VJy��z`hu� P�B�s^�L^r�؛S̓���7�
ݾ�ob�j��ة�n�P�͋���uE����-n*�F��8���'s�x���1[�Н2��8��{��԰Y��s��f��b�(;�f���rS�W��Θ��Ym�>lËsJ�Qώ<%,'����+3����qbl�:�r��:�	x���4��p.�ݸ[VU��h�T˝t�����{zz�xYM��m��m��m��h����R6���b��Vw* �Z�ǲ4�q�#�_fuL���Q��oJ�-5�򢚠]G���އ�K��r�j]4��,�љ�m��`� @����x-&��[�pPɢ�m����h&�?mAml�j�;�f�Xn���w6�l��I�|�C���wwt�ݳ��r���ygf����7���=�����EC�'ǤꝜ�J���'7d��֧�iDJYj�T����=�#S��v���w�0V߫�G���Ty��&|(�\5)P4������iG��U�F��;�Hݔ	���5�v�Y��<��8�J�:rA�H-N�d�P��u^�|�l������q;�3[��y�s�s�{�8#mc+��.+k���JZڬ�W*����UChQ���*�m�R֖�*�q��&	�F*�b�l�[f1q�-��ċTe)X�Sv��Y�,Qc"�E��IU�RŶb�U��X�Ȫb7Y*5��A�#mAA[ERҶ�&5S�\��"V�Ci��*e���,)�i�V�����UV1Uq���r�b�`-�E�-��AT;�U�v�Qv�jҼ�7�VPR$`6���1�%b�ETQ`(�/���7�禽����A-L�A"�ŝr��R�n�����5Ns�	��I�ǩ�Ɇ�����q@NU+���Y�T+m/Z:�c}|�Yy{�5���|n�a�խxo��P�\ ig��_G�p��k*���;�0�u�(mEx&�CS���~��� ��h��
C��f�ʦ}���'��ywּ糯}��#@b�����fd�9��s��Wu�Ի�2\�rvvdC���ޛ�r$/��Gk�-��ǋ���=ҽB�x���]^����`�y1��v��*v���)U�3����v��<���P��3�+�R���{���Ǭ��e��ڣ���lI:�����~jq�#�L�D��E�SyQz�v6��{^c�'b�E'*�\�u�_���z���Z^�'{�����h�X�Q�|�qȲ$2�/s���k�}��إ�,�9\cڗy�N����S����*D�o_3�.g*�,1��QA׈J�*b�o>Opm9E⠸ǝ�	��6řY]��ʵ0=}�����[?�~�N4Х�Ku��<"&_fS�}�|�� �A�fGg<=��lM:��<�(�S�i&d�t�h*��35���	�&*n��Ǵ���,ԛNt�d�n)0���F��X��_�^�UN�n�a��V7*ĝ]0g���e�J4u^h�ϔCf�F&_r/��o�4�����G�Z7���S�1���o:x���x_���P�}S�+=T@P^�h�L��kc��K�]�
`����^_����$Qju�T���x��.γ̘�<�0��5���ڙ�X���_*��^w�q}��x���N��d��L�c���[�Ñ)���t�a�\)���=��"�'����sE�8�0�rL���Z�k�5��P�����Wq�\r���^��Ws�+W�Rx9&�J%X>����YgN~ë(�M���v��7a>����V�_tz������ٵ��
rs��y��1P��@�BLXv��/oQDf��yۣ�,�N�"�Xi��2+�of���k��R5"�m��g�.&��<�KZB�Q�ws���vX�ex�.����@.����ۉ$x��������2���IT\j��J�����W�҇r�Թ"lF6:��ь�-��Yk(s�FeD�S�W�:N�K0����l!� ���&��+����-��aP޿wA\�=bEҭ�٦��{�B��cһO����6�)��������c@�9��jt���P|�����}�_��
S=R��Rz]��-{�^��{j��&DLQ�:�92��Xr���$��RI�x�Lw�J�l(�j��E�S�%�p�'yd��L��h��� �9;���Lܢ����������4�����7~�{:gv�j�8��#ފ�A<��>F�1�Wu/��X�R5�� z���p\��=/���dҞ��~Ff�r���u=�l�}�KI��3��gp��0�W�w6�_��gw�V)M��H�V�/{s%��-�M���4%��LC޽^�}��O����}wQ���K=�|�7��ώ*4��[YwQ�Eң
<���Cfy,U�ƌ��5��7�60=���:Dv��]G�{�!wc��N:R7Cƽ��n��\���q�{�2v�+��*#<�F�V�bP`ϴU��m5WF�+��T�=ƁE�N+�O�b�����)Cw����ةZѵbV��9�,W���4��P���W�����{=[��4݁q��pr�ܖ��k�W��h���ǹO�P%=�}�s���Q���޲�gC��#��^�y����;y pꒆ0Y�����ɛ9�~��R���*u�*
�4�������~\�h��Hŗ4��WI՗�;�o/^���۽B�����<^���i;l	rmmm���Z�R��� ���E���'�n�1D\��8�&�VG[�bg];��_I�tճb�\%%D}��=|�=�.�Y�
����ymMπT|��+���"ͮ�K:�,�th��XF]�vsas�h�v�t�؂ؙ���Ԥ&\���d���j��2~��-i�*v�����`��m�5���	Snkci9�k)S���	I�b�׷@
d��ۘ�P�&f�zt��ߺ\�J����pnn>�+�G�����j"*	e�/;��W���o�g��˛1gTjX�W�z_�eq��V�I9�;���A{m���e�Z�Rf>j��:#8���8��RǺۋ���]���dd�8�/��.&��۾t"������x��̗d�c�z��.�.E�Ee�s�q��
�h+�f���}��h��{��j=qB���#(��I+VA��,�9�y�z����'?�|/ut~�n�����y�u,ykM��C�+ߺt?��bɑ�sb�OMx\�����#�w����<�)-1����p�KK�7��߻�;*��%�
J��`�sg�c��όO����y�!��h<��q��/��u�I�Sy4�؅y7�J`�i���n^��}9�c<Dtj賝/ט��K.��t��{��h�⫒Ķ��;���� ���KOf��x�ì�v&�����}�M�C�8b�tz���em��]<�4�=�b�T�����B���.o���y1�w֛-�ܿ��1�m��w��ġ��_+��a8�A����w�)��ö?r�Oq�W�K�\F�73�h5���1V}y��!����/l���OS���*l�ӯPG}�3<�U��řpr�:f�WC�=��5����.�gH';�7�>�m%�b5��2H{�ש�|��,[P42�/(�$0I�^���gʽV��^�U��Y�ַ�������� ׽�S��������e�p��x��u��MQP�s�Y¬
�4�+{�mEq���F�6��d=I~	*���鵔3w��K=�է�h���9��)L�sv�}Ҭ��w��YX��]�@��6|��HU۠��xo���]���Qћi���-�;����Қ�p�������̭:!����?	JW�ԧ,����M)%vi�R&�""͠���R�<��vC�]
̱��Yƒ��b���N������୾�e�*Uգ|�-���E|e�d�WQ�:ޠ�θjj��af��9X�<��uv��q��ӈ$$��v�Ӥ��F�ڻ�n�y-�G���0<e��ԺiM����)i/�=Ga��	�k%<am���v���9�(+��0���xQm��m��m��m��i���9�C�����W=�������w���_|��`��=���8�1k͔�t̷���6����_W+v��&���I��9��`m��],����A�pu�;�ճEѼ�n�-�iv��KƥZ�f�<cg/c{�K���&�bWv�dU�g[J� ��9�M��VL=���vt�}9���%=�1v齄Ԏ�&ڥz9�q��*_9@�`ܫB�v�k����-\c�����}	�Rn��u�ȷ\�*u�>wNY��/��-5l�:.��յ/)�t6����$��{��3��t��<�M�6=ɑ��O{]�{8��s��a�������	��i��~<M�v��GMr�C�eeĲ+i�$�\B��܊��`�PU�Q�{�1#���Ś2�{�f�X(����U�
�.Z�q�J���AUb��AE]�,X,�5�-������"��b�l���H�X�̊��YZ"�H�&�H,E�X(�T*[J��;�LLCP�@X[H��J�UBQPX(�V�(Ъ�T�C
�-̑qX%�ő`�
�U��6�Xnn�5�߇3}g����U��BP�zL��v1S��^j�D���;5I=��].���b����k�A�M�ѧ��x�(�����f�\7�Ѵ���<�A�����J׾*��Rx�4�ߎM�џɍ�R�k>�f.&㩼����m͇Z�u\�eɅ K��w�꡾�l����^��J8yrF�ۗג�q7���BsM����AB���vF}:
.�U㙲2\�m/!�O�{� 7�%\�u<�+��7���4[�.&�����G1{}���(� �(�%xz�پN2;P���2�ޚ��L�o�|�]i���J��;m\eT������~�kb�Z�Ѽ��Q�^����mg���E�X+��f����?p�����Q������Cy�f�+�uZ�qZM4�Mίa7�əY^7㍨V��y�Z[��P�'::�4{9���=/�g��Rhn�|���V_�5��>��	|O�/)OhR�ҍٞm�i���Vw��ΧF�j{�g�nȜ3!�Y�<x'���2������̮��{6�oI �u��Q���A�\Mk�{t�����d��϶���̐m:IִVФ�m�LQa�d�%"��#����g.X]�p+KO$��_{@m��"�V/5Ni%�cse���gle*t=Vˊ��k3B'��u���0�y�%�C]�s�^vvι7;�OB}9_��;�5t����m��1��ӹ���~���m���^�����ӪA3�Z���A��ҊwsLupZ$��؉->�{�:Y-Rb�%�L��s9�%�r�w��H�J|���U���.���Ӷ�2�z�I�GN�jʛ�=4Q9�o���'<oX�}6��ږ�\���{�N�oq0oux�{�y�x8��,�Ȯ<#j�,S��r�bgQ�W��s���ٓg���=|��s�2Wy�w�8g���׼׫���w�W���ڂC/�u��b��rϻ6��^rèv/,�8~�I{�ͫ�)-�����~�2�N}�t�."^g0�5�4n,2b>B t[����d5��#����g���ٶ�9nnQ�p,��C�mOC�_tA.�J�
F��s�����<|Z�X�5�����o���͇Ƨ��W��R޹=�j%���*�^���'�n^����Zr���[��Q���y׭Dv�c���E6>J��ON��#O�bct��o˹H�Ov>�絛'$��{�����q$/��@{�D�7�D�Sj�^�X����j�������������X��ۑl�3����{��y��ׅJ�9 ��MT�nF/	3�?\������"y.���L[�m������?*d������@L�
�+��]�\�4���O7Vu���O�ٵ��Q{Ry�ǻA�{<����u˯Q/��1@�;ý(��К|ȼ�F�d׃��;��*
��&�e���`�=2J���ͼٮm[oe� /���s��� $�Q=B�JTUG�	ܝۼ������'����o4l�7�ԓM{o��^Q{�ܪ�{u�[Yoy ͽ����rN{�X��8�$;;z���K�P;��E�N��
��N]����~9@��wS* �׃�ɾ�0�$�Q:����[�t8mz������t'W$�lV���IQ�vL���HF�o)�6���\�Ve��:����՞O<<j6S����X�*�����5�Sg[�ڙ��i�xV?'�f�i��&<��Vމw���*��Q�hs{�R	ã�.t�;2����a��d�fwp�T2�\��I6?�Wk^��W����*�����a�։�޴s�S��R�Y��י�����j�R�g�#cL`V*1����	�ױɡ�DpQH;~�:3F%c�V�^�-M�=�8d�I�W;͜�'�^>������oҟ��ֈ7��Z�9���^���Q�Ã�Kgz��~�{u��=�H��J�ke$��Q�^���[é7�$��r������[����bMo�����(�֪ ���q]=#��x�d\��x�7��EAq�⿢V�+f���:��WǺg6��ؾ��t�o�4j��4NM�LM�log�R��Ӽ})v~�������v�8p���<"����*��S��M��5�@�͑:[A�J�lE���Sʈ�j|:>i�{]ܽ�leE[#�h���H!����`_s�{���t|݁��W�T�2��z�U�*�	�����h����L��{�x�e�����]����cz�LA-�W��LI�hN��{��J�5�&��7���6q��>^���3�$;~��l��[�;��ne4J��Β�2�e��:��Lt~���M�	z�'��FJ<�Fgo>�qL��#o��B���K%�� �/�^M�-�u��.�bh�o�p�e�u�+��.�Ք6�r\���"<&iԺ��}���7H�����w�g����l�f��J\��O�yt�^r�V�D[�6v����GQ�^1�=��"����ĘI�K�j��ս;����&�1����R��e%`��gx<Rn�D�S��.Ͻv��(a��:^��͜���������bT�>#�C��&���&�<+��
�����| �׻�G��z����fp���s��sJ<^S��Ǳ��:,�k�ck�������c7���lb�TǕ���j�hQ�K�*Qk�*�,ԿL�O���q �TӤS��(3s��̧V�^gȃ���Y�L����ax�~�x�L������R����E�}޹]FɯvSovI]��lY
J���C�c<){u8�pg��7���E�a�[Gb��t��|hr�������~�׌���}�����^�˥���*���/���� )
w��C;��nk���?p�G�~�슟��������%PUk(r�UAU����UWPaD��!��P�*
Խ\���a�����M��7ѯD�Nn̛��P���KQE
P	?�3�̛�M��X�'I�A1���v�],�J-3�{�mh*���A�\��l����}��MHo
���z�Q'Rl�~�d�A�<4C����}҇}L�0�)I���{��� �*���b��PU�D��9fW��tS���EW�qU��D�(�8�G��s2�������b��:�_�U8�Ͱpa�P��UAU�>�yS�P�$B��T1Q��c���п�m �h�P�X)O���+u`[n���$�4�ǕC����9+UAU�F�t�m���hVzp�p��
���`5U��H�,��l������qt5�����*���[�rH�7�Hn�͆���=��JV�˲���l\M�-�v�K ~�����p/����/񡯈Ƃ*��4X�*���SYs��!8�Cgڥ������(QJ ��%=9����K�>��2�¹�Ϳ�q�����rAU�,	�G��`@�I��# �d!pOpp�J��X *�T;UPU}��p$4���d��ʁ���h�.^a�%Me�<Ĺ���*�����"@��
�&��d:�?�B ��H�(����H]l�'�~�ì�I@@�P=���!�N���LIiN���L���: U��9G3��)ЧP�
��'���+s�`S�{��34�3�:@ޟ�6�*
s�뙅|�@�7`�j.�q<��F�	�L>�L���PUW����t� ��%(P@���$��TZ/��~��5?p���@nA�~�#�L��55��ߎ�1�1@�R�t0#�����@-��ϿA��'54�<ǦL�=�ULGA�7ׇ`k��
�xp�K�S���t뽈���(C`h{�٪D�Bex^��,&P�S�Rm��A_���W�
��M�o����q�"��zN�ܐn8at���-f\(.LB�׺�z+[SZH�����GV����"�(HUZ 