BZh91AY&SY��X�֑߀`q����� ����bA�� ���II�l�6�J٢P���ٛ4��*�J�ٵ��$����h�6+-�k�� փ3U4�X%�T�4�i��S �Y�uq�Y[m��ڕ��MI�d��mcUF�m�6�df��[-�[6��)�Y�04�2��l�h�Q���m�5�Q�[��f�V�h ��uJ{f�ڥ�h%Bت�kkY3Fڈ�kd��6�,�jՅRն��*#-U����-6�eM�Y��km*���1R�iM��Zԍ���5�48V�m��n   �w��v6�]�A�uEk�]��-���:n�mY�M:��u�ݺm�{�������'m�W]wt��v���V��]:�Y�RcmQL��ڤMl�|   ����iU�=/oz�jlk�K:�4�7�=�K���+��^�U�k����6�-�G����J�B���OzT�RJ�zx�R��Ǻ�\鄨V{i�h�m6e�i�U�   ���EN�%����m�JT��w��
S��s@ju�n==�UN�U�{��IT��{�ܢ���.{��m:��R�p�r����޵�u��%R��VeJ4���ͱl�f�O|   wx֨/��o{d�P��㧫����zw��4
]筻ʶԯY#��rJUw�wT�U�c����U����)�����5+ٽ�{L�-f�1%�ն[m�7�  ���������Ri��8Z޺dvr]ҩT�*���=I�nƧz������UJ�L�c�t5v���=��*�W���a��P���6m+4���ֵe�F���  ��ۯ�T�t{�R绩%M�I�R����͞�Q(a���+�UR\9��צ�v�޵�ꪝeJW�W�x�4՞���&����UR�K�추��9�F��L�2�4���  ����ڈ;�מ��l��������]���s�罹R���=Gv�R����8%"�V�)��oC�*�ݝ*s��R�R������h�Sٵl`*���kcj�5Z͟   ws�������@h�U��Ѫ�������W�U���Ҁ׽�����4l�ǳ���T�t��� �q�#m�J��l�*d�4   ��5������ot=V��ܷ�I�{9�+l��S�;�[��������u�U�=Q�y���Q��g������U���k4լؔ�2��m��  ���Q����4��n=h�;���� �^�^ G�ʺ��N�{�p)�9G{�n�k_  4  ��2��H4  � � )�4b����@�  2B)���Pi�      �~%*�� �    ��&������SM �	�&j2&RR��CSP�#(��&jd�?��/�_���B��9?��(�N=;�a�ݟ^��f3u��~��=�Xɨ��   ������6��m��o�lm�y�0��������������������cl��!U?��m���ߞC���)�1����w�����c@��v�gm���`����3�o�6�Y67�� ?^@�&6��m���9��v�}d��Y��v6�ɍ��m��8�}g�Y���CY6��o����lYc� �� `�v�Cl`�q�7�v�6s����L c�8��}g >�m��q������>�1���`���6?60}gl!�����l�pcm�������Y��Clc� ���}gm��LY1�!���1���Y�7�pc�8��}g�Y��� ��7���-ژ�y�����x�U�����ėPf��t�z�	@��=cm�ұ�O�m�����[�Р2���N���6]�LLe���RIHC���A�[1d�e���U�w u��/by�Z,��L �vO���uiݹN|UK�H�d��EOMؖkR�G]Go�ׯX�w��^%�z��ϥ��wNnh�f�aݵ���!���n��J�%��|�5��_���[�!D�]�� ��i�-�M*��W�cf����P�X�ٓo�z-C(=�su���+Cx�I�6�f��wq�)[�蕆�Aֵ3�����&��V��VC�T� U��X�Y��*е-.,fcv�Pr��Z��e��� ;u�P���͠
��ɴ�Z�u;�1�z��0�k������c5&�����q�1
ؓa��� bb��on��?(h
y�9%d4�{uli�rk{�v���"2�&�<��ʅE1,�01y���n��#�!jb,3V�m���V��!��{��d���Z���(�8�t��ku-�D!^%xh,1&�`Ů��Jգ.�̷$R�&ы`���sf���Vk�R�6��Z�ɀ�@�n��R�y�Fh�2%�gs`i1R�x5�S������/cN�q��Hkv�Z֡���y�+���Ԡ�4��x�h���1f�li�1��ks/G.Re�N�V�AZ{H�v�bNCDޜ4[;"!&%ⶱ���֨��iik5V��][����,`��x`���5���6�ۊ*PI:�ɫh��[�4cbE��li��0��#I�
/�7L�XwF]m���4��¡[�����ՅP'0�,���A��KzH��`����V��A�x(�D�ں[�b������pnn̙��Y�$��2��F�s^n�%�Jce�wA9WvA��8�yc�.�I���.c�F����X�Mպ��6��pQ�n�Yu(#Wj�����q���Q�[�eEJ<�7v��Am�)�Y*�U�kn��:T���]�T�"�ش�v��Գ��7���1-��� ���f�"?\�|$�2�S�x_��`����qh�n+��M	U�n�2a%QU��y�-[34��©a���r�Ң�S�u�T)��M�/D�1)��!� �-�2��Ә�u�Â�RDɸĥ�5Su&jY��Y��[���
�l�զ�N�df2RƠ�KdQ&H�JcT.�ާ��+���x"U�q�.vЩ�Y�ڱs	�(U�tQ��jd$�d:��J�',d:���
#��sQ�z)
vV�;R=�T.*9�KF�:6�l�3+(Ğ�Zk �Ҿv�0(�1`١�j�R����+MB7a�y�[3�
b&�B���p�o&4v���'Mo�nCYA�i�6���W�3(J��Gv@@�͓2���C@����q<���U����kL���1��3/��ɮIn άGh�5��=���6
H���LH�ͩe�Z!���E��.غyyj"��,5�����p����1Ru01[�_�r���B�6��v��7�f)Y��j֤�S��E.�/�3*3�
�oN��3h�W���imMV@8�w3%�`�u �ٶ!MTz�-�Ph��X�2�4a�1ݙ�j­���5����;�k��r��XE�K�L�Uy�����y�"��u����6-�m��E���>���S�6c"�Ĭ��Vi�4,h��p`��MFi��k���u4&0^k�^����[��U���Lh�P�0m��bl�����ٱUx[k���駶U��I��gU2���ލ����/B�K�R��PK����<�ɸu��KO0s	ע
'�b:66ԸP�����`� � 34�k`��V��Y�&efAR�7P�X�ֻ�X�^펺`�6�����m`�B��]Rݒ���`����#r����Xc
4�l�WcE�V�6ګssn�8���K^;P8��V�upE0̡�n�S&M&�;�`� 7v�������Z�^cn��t$7u+��N���6E+y�9��D���,�B|���af��gv����M��M��i ��� ��6��Q�/黴R�b�w2M'-+���Fd8�Z:��0�N�RIA���Z)1��lï�+v�Yh90S}�ԛ������R��K]��Q[OA��4̄X*KmVb��1��m
t�m�:i:�m����l�D�$�Qk�b�i��!� ��8.��iQ(J�Y��:R˸J]P"���9Qen�ZmϚ�K]A�@ �������4�.'N'�ͣ�6)�JڡH^)nG���S)C�]⡻�[���1`�`ͳ2c�44�A��"X8���n����Ҟ�oX���7��ǚ�o��֝-�ΝA�����I]�UiZ@� �����(�{��ff�;�X���p9��u�|�e`/QޮT�>�����yJ�Mt�`Xj��lY6�'r����«����|��V]k9$4l�x�r5��P49r�a�f�R}\��[w��bT�y"�U��I�O d����a
�5�2�W��=���cv� F�讦ݭ7{���T�}u̓�,f
�͚h�޾*�u�E��W�x�v�vy㦠.��%�Հ�����A+�ךKǠ�q�8���{�4�@c�n�vdR]n�ț!�k�2n[G�m��Sp`�b$E^��1`	ڃi;�*��(���H`K�-'���Z��]k�#iR:�эY�-%�U�b`ï!�.���nL:��6�4@����v��/�nD�5i�&��v=�����f�)�i�2�4��2A5��,���ܷ�r�j�q*�J������6 GjC4�wZc�Y�w��kf=Tܼb��1���]�0*݀��0M`��I��恷{6Hn�%wF��Q�]u�_hޮ�u�5X�;PR`�[��oI�ԁ*����6�z���Pݥ*I�kPD6%n�nm	;�iG��"*o�M���f���	��\����f驩��4޹4�43uT"S�*f�5�P��T���{F"�x�F��l��Û.᥄��h��t�+2����"��JR��lk �7XBƚإXSR`��R�7�oE`�s[�%4�n���`����4c��6�FV*�E���B(!���ª4��Z��6$�*������̖�b�x�VaP���ۦ�ڛ(F XTfZ��B����6F�L
�AD�ퟎ��M�8�/4�����z_P �{���I��y�u�vN>��Z�0��Ҷ����C�XرcQ�n���:�ڃ�oa���w�f��ը�K��L��pk�"�����mJELm��v�7T�����0`����
�(Uٔ3r�7���N��]����,�:�%�E7͌o8�I��c�V���,f&�0.5�]v�3���C���nT�x�h�fYun�Z�k�x-��e+�8�K��bv�a�7p��5���G�t,x%k'	ͬ�����b�� ��[����ZB����-٧3�u�<��T�W�Iw�/ u�Gc�t&e<v�ͼR��O2D��4����)m���o�$V**�;��Qg0�X7���7o!�/gܷ�>5�p�&�)�h��W�^Ao.��T���nV�+�w��6�r��Ta���]�Z�V�緖U�^cT�7E�޳W�sX�;F�y��b9+4��Y�ڊ�_8]��˭ǀ:����i�1\3mR�b�ln�s!qqkїH���.�I$��+�i�Ć�+x�(U���c}��|�h�hR�zĔmr�zM���So1l��JT�C)b@<mbe<��j*6H�W� ;`B�`u��˽{N]1��\t�)���i-��(�5��k
�UuV��]j��8�)
|))�qՄ&ˊb7�D�>W��W2���+( &�0�H�NUn&�(��tv�=-^)Z� �7����qƐ�[�v��ert&�h<����ޜ"�J5�o)j�&f�"�n� �kl�Wc��w�����9�B��M[D��ncQ�0�%A`�.R��SʼI�u]J:/��8U�K)2n<ϭ�w��7Phl+����lf�u�BWNVe�nTiesi�Rr�+U�����L��`+/%b��@e�2�-��[��"��~�Cx���*�Z�v&�N�$�n�7��{�UXF`s$���m�+rjuu��UI(��w,�ɚ�^Ic^|��Uk�t$����XA��h=J���D�ܔ���1�/2fn��j����j㨃Z�1�F�FEccwf�t�GoUi�B��f#�����3C1��3�d&G�M�Q�V�LY�wOd8�f��Q���ѵl;c��
�.��@ӫ���0�[�eI���Ɂܭ��[�������:X�1w���[�C0�&У�3�62k7>D��E��n��7��:t+��N�[yut�:�G5ݣ����r�ICJ����x���n�ӥ��k1& otmJ$A
7
�9���%Zʆ��
�bT�L��� �^Px��Q1NF�L�E�ۭ߭`�/9�%���d�V��d
����R��,�,��*��l����8(���,{���]��Rl�`�{G4[p�<�ǨK����4�Gx�<��v�:Bqk2j�V�s7�A0��uX$������W��ub�%e^�73#wr�)l?Z����w`����ݙ��H�6�����m�m���_ib��k�V��gSY�]��-P��9Yn�ջ�
�R���HpG������n�ܦ.����&��1^���C(9�H1�*�n�R�d�j)�M�4�b�{w�3${a���ō�n��$�3M��~&��B�2CV[��B��
�b<p�{&:F^�V0n������ф]f^�Q�ID)��,+.�j;L�Xl�'�e`/hvnnn�OkdXX4&���.�e5�[m��RH/@S�z���7t5�×yR\R7vvcJ�N���7c�Y��2��pMF�E��s���;4C��kj9z�#4=���ȋK����ұޅ��pu��F�f͍T�P�eʙQe+GFl�
w� �����ߥ[Պ#*YQ��nn�7$����ڐ���N�3kje�f�
���!��֙b��CSf۩��ڏLf�okksraR�`k����C�6��6$q��wY(�����x�,E�c4@wm<t�ٍ7���їG��S�$����{խ�n��w��86����M��ulj4�zVe$Z�Ëe�&� �X���7�kqT��(���'���k吗�[�.�nd����+��*;Y�\�����ne�ש$k^�����rV�,(�ݭ�p�)l꒦	@i������cb5����V!y&���T��4��y�7mX",A���&ح������l'��l� �aX	P2]�(FU��`i�钣�E��Z����v���8�������<�cCͽ�������Lpc�5����u��P)6�Ncp����x�AJ����2��h,2�c�NK�)�^4�����,i_���Ɋ��V6�����M[�+3w�.�H*xk�_Y��?h�;� z֪b��A�C���1@Xi��]��j�C�m��������*JAQ4����2����;x2�)&kp[�7w[� ���F�j�sB���4�*�Ud��CJ8�/�Zٹ�e�P%>&0,����`�)�l���7{�������kiP!܏#������\߄Vp7{Lڋ%K-�1�i ��0T��$�M�]��Me<[�뺙��V�`��܆0��Ŕ�W��u�	kp����VVbx�ld$T�1ū$kq�D���4��^ʷ�$�0NV�V,��K�Nc�$#XlRܫ����kN�vfVF�?0w�z�)��� l�{��u%S
`x(��%3���1@kh7��F#�ҝnC
p'u̤�����1�[/-9p��Yyxuʣ�*Q#�Y%�x��y����_M���@�6�Ș�sl��h[ԝ��覀f)��c��0κ�"�ذ�$頛J��ش��f	��j�Ӣ6:�y�S��l�Xh
y-T�Nb6����ieᨵ,��ZCM�^ҧ����GHp$�ʀ����d�X�c�xXY�e�"���+�����݂h��+ա�
������$��fai��d��)�`���҉�&����0nG������ۀ`8��R��fe�c0h�z���l����i,z5<WgEɗ�cP�#A�F�� ��Y �-V��|Te��ln��CcN��V��^d����F�7U�8[�1�����n�B��knE�wH�UG��[.�e� x���L%YZ]k�쳫1��!7��_�R����5�����3J�ޭOya��O+�W��:&+umX	%��+.��K
z~�vx���Ѡ��ǜ8��/m�4��(TA�ȮEk	jm��;D|��Hn�M��t�[K>���h�p:5�X	,�/HɻY6��1HX�5R�J��,K����5ͅ���I'b�ZV��Ĭ�5�)��7�C>{�԰Sӷ�P����a�te���[�M��o٧>M)���PZ"��%9b�eU��lfD!Xw��a��w�4�@�`M����yq��OJ�VPj��PG*=0�V�&�T����R�W轏��U�4�
4����`Р�z�i�zmb�ʼAZ:[h�� `�
Lb�b�V
}R�������ɇ����vβ����aZ&����	��(@1B`�3��w�  �����dZ�Ŝ������
9DN���]f>��<���v�||������H^�
�����~��� wB�f��w�ҷZ�`+�E�<��`��9+ǣPV��.�J
�X­t�N�j�7 �m*q��mk�[�%/��E��U�7�jQ�����A�|����[�zEi롙��J�۟��lNPTse�	v�[�[�~M��aN�Qs�"��H
W���x����Mdd��
����=i�Σl�.m��3����c��,f$����E���n�^D�a
h�Z�킱Z\�,*��Y�)m]z��)��X�&�5�n����ϧX8*A��:`b�Bq(�y)��u��f:-���CB|�t-Z����f��,��U����z �j�-�a��N jڢ^��1K*�3u�ogW3����wA�xM���9�8�Xs���:�鏐��&��~޷6Ҝ�`q�Z�׭�w�$P۲:�����@f�0@���团˕�1 ��F�9�;�&�m.(�Ʊ�ϣ`����F���bU�M��.�W�}�n�e<�S�T��Q�=����S���=��4}|�;����q���9�G-QĪ$+.q��[���Ʒ��ׯBHLr]2<�fk�o�9Nϯ/4գ7v���X6n�L���9�5D^�����gh�p�J�T��0仝�f�Lwi
}w��fl���<"(���͌�:���TUp�f��2;�7b��c��MUdmJ鹡Ni�E�}0v�q�B9���ED����
IPx���~CM�#iT]2v�]+r�� ���$:{�&��%ݧ�L��go�dQ�5�v��ucm��Z[����Q�,�	-���Ծ���[�i��T]�x�T��룥�+�K7(��5�6D�gIo�X�J\�fma�2ئ�N��x&Z�˿��.DIt��N���ͬ�y��}{6�uj��O��M2��bVժ0�bZ2��c<�ŭT��ɚ���2!���"-H�GY�t�6�5W�9�7��K.�n����i7��$�^J �N���0U��ڽ�'������tc;�n�V[�B��p��\��|KXm<�j��J���u�˧i�ymF��"ŸcUú}�����o�/�K�Bgn���XuؐX #E`q��+�PɰMѷ�z+3�qai�����!��8���b�I���f[��:l2����ʭ(��T�I��;pY����XX� �04FQ�(�˺�)X��(!x�zwV��>ݴ>C��w�n���-�]������\���˙*i�R9{9�Q�5��H�J������Β��#l�ʆ�_ʙ��/p�]L����rZp�S�8 s��շ��_QQe���>�h���L������q�:����2��-t�dK+�c7t2G,
zj1}�ni�t��aB�+Omp|)[qpY]�Mvk�	c��1�+Z���h�*����3��n��88	��w=eU����0��#z�y\��2	݉��"�3+�m2q��(6��n.�3�9�7bJrwut�/f݅8М�����,n�$t"�]��*��hH��H�d�o�����|ռ��medA♏�%�Q5psz2���޳s��A �e.�NK��:ry��h9��c�v�r�Mh]k�{�MXQ�<�7��*��m�,�v4G��N�	��n�ꖺ���SiF���U�E��҇IXfs�1d$��o1B��ȴ�̣N!�Z�M>�o�o*VM^|t�Zz�����c�6�H�V��jAb�;/�w�t�79���w�(yp �T���=�։O�:�됓�aޫ��:J��&zVк:!�4�s�S��m�(�#�`i���D�m�l�j=[�mt?w���=�v\ey�\��]�oL�mJ��]�r7>�|r�KaB��mKӍS�[�3�掬O&�m���(�Y��c��M}�lڈ��A#:ڄ�:
r��!�sk�T��`�0��2�-�[[���u`����E���;�
��qcm����`��9Y����2�e!�G�o  �6��\i�z���B��"���v�J����n��B�,��aic���,�ˮ�h��..M���0����m q�Q�7!���rP�<����5�CZ#�++��.����z��������5}uq����G+{�r�`����N��pT�7sjƶ)�r�C����TuHu�Pлn�@����T;�n�x;]�ؕ�q΍໔UXv����/�e�@��'2�����`O�`���+G�Y��cL泥R��E�}.������t�IK�/>@�jU��ʄ��qe=��q�mZ�b�x�%0��3�v�]�3�X嗨��&t��;��֤o����<��g�!�ᆶ���r��viщ_P�b�Ձ�@�:�-7;i1�l���բ>�)jk,���r�_Ϙ�S�ʂ�]ԭ�v�ˬ�J���Rq� �J�m�V��m�����v�bJ�c �ƞ�;x��:F�ۄvT�����e �Y���f9	�@��W!�s��m���� �}&��ڤ�åݑ��\>�^�{�}�H�.�cM�W+�����h�B����t����iA[��f�}[��
�B	-�ml5L(zJ��3:�S������v��� `��yu��hJ�]��a���9��łb;9�X��Ѻ��ܾ���8Qغ��S�݃�@:Od�X*dl���,�t�Y+�S33�{:
2Hv.v����я�u���+<���p~��	N��e�$ 꽊X=~�����$�-�J�W. <�9�S�U�9|�[������=�Ws6bɚ��J�o+.fMY�W�G�]�_WS���;\�X狭T��od]v�ͮ�Fŋ�t��w�qEZ�)�܏�?aě}s����okM��$�7��3��6�-�e�єEC�Tr-Яa�By���1�G�5vn,�.5te�W$�+c����
�G��Lmg62ں��D��B�S�W+�'���T�]��Bp`ԁ=w\6�9�W\+�ԛ���4A��o��\Ӑ~ed7� \ŷ<�v�͆!�)hA&|�0t���qP�8����OS�A*Rv�9{��N5Y�� �R8�9�W4p�[bQ��9��/��������ц�"���̘�OF�rj�e�{��v�L1"Vv�K���B<�W��c�6{S9�	vNW^��I���[�v�JSa�\�֦���M�ߕ�l�	q��9P���6�D�(��B��ƭ��Ɗ����A6V=����V4��Q�>�d�[Fq����6�N!�{�F8][E)75j���#��<x٭�Y
��2��(�ڎ��ܶU;亐5t$Ug���s�]|�:���s�^7ѥ�.�n��S���ѡ.wj�����{��R�Z�V��OT0��B6}u\�\�`�/y�xQ��Y�d�m�N�Rޠ�Ie_u�K��)���`ܭ����J���}�x���F�����.�C:��t��2�����T�J"��˳7L쏍�Sth΍�O`�[\�l��r2�Qa��]!���+���T�:�������`U띪���M�VH�P5n�fARc\V`xF^������,
{A�ǪT��5��E��J���SF�*qǝ��^�̸,�_U.8/B�]�E�(㏉�Ee#[q�>�I�c�A�<�Nɖ��2�,1�4���+X�Q���W�a
�%m]�ˮ!r�tN�щin�eދ��H���	#4.�Z�*oy�:��Nϗs��)e
#*�-�Tc��.��;34��.�E�\�J�ƭ�`ʔ
�ߕ�Z�%Z']4g�ݽ�/�R��3a�J�	��h;�]�mE���[%�p���Q�9��v��\w�'�2:ت�˔/r����-��B�Y��<zvM�MK&�Θ�R��"v�7!x,+�;�]ҸK�d�� A� �c�έt����	���
W�e�ՖsP�pv��
3A�į�X�ޫN�tӒ�`D�0�q�]83V�M0��G��:���|x��z�l*_Nє��*���E��6���Q�e5�BJ�Z�65H.�çA� ����{���8�64J7���Y$es�{c4�(�.�ؕ�c��ԁTne��6CWQ��%v�(kz9��v�����x��"�u.f��;����YٗٻYg{Y9<�$Դ��(�o���fhF�ic�n��wK/vvlH��kB[����c�K˴E[��8/8�y�򹙛�KA��5�T!�c�[���4f�
�v�Ɏ�g5;+�Yu�
})�n�\�Nu�\�Zq��1��S4s(�Mv���T6�U�5i1C1���=#O�P3T>�w���l�H�K�EgTxl��u�FD(�ZMl��\�s���1��K��Gy㩶)r�qG՛܂�-̱%����̕d�>5�����:��('�U�T�����,������/����5L�foj��\t��|PU�_2�q�d�]S���;�n»YX��J�.R��oS�mRW�he5>)��!{d+������;�J����*řo+
���pP�#Mp�⤷�$6����/B��.V��E��Fk'��{�l�T��#�,QS���N�qj� v��/�a���U���'.�;��V�'C���.��=�`���m�x�e�v�c�E��R��X�/.'�K��*�}R:�q�w�Q4&�Rn�"N�l��h��[�p�r�!]� 2���rvn����0���..�{�{����S0���:2o̶ۨ$�.N*ū��+=�34ڴ�r@�y�[��o�|�����s�)����i�׺�#(��j�2��9�49&u�� ��(aRiQݔjx�.�p3�3j�u`�fKu�){�ܛ��
<���*�"j�0��}X����EN�xٮ�W;��T闭�Ӛ:��
il��*CJ�l츫,6�jȫNe�{���n0yQR��ph�"A�ܽ�N|x]_��)D1Y�_w�"��֎�����o�7��8^���[���o+�r���҂vY"��&�'nfj�L�
��6����Xݒ�T����!J�;�����m�]���F�#YQ;�|����p�"��=p*p0���V=�c�`:��� 9=B���`gm��њu�_l)^��Bt��"�����G����<=�b�i��7�[�{[e�#lAIm��60ج'g�fr=F�ub��<x�z&l�Y���Jؙ��)��@�[��yR�u�x������I�7�Vd�܋싺;IP����i�͛�S�pX�Z@r��/�٢d����u�J@k��ߦ���N���.�=�I(�	[��4����0���%�C�l]�PͼT�_	`m�N�;��ā�L�������/�n������Xf\4f
U�/*���u�f��Y`������|�Nm���5PL
�lf`:�A��,�,:��rY���̭2�q�lrӏQ��9Nv��s4��'45VP���sj����Klψ�]��ⲷ��#��������h�,�Z/^�Y���<zK�Rf��nW&�r�:a�ݟ'}m��K���i<�˄�t�L]�yR��5$��d%Z����|�ݮ�.B
�en�}P� �c%͙��w���q�jn�X�t�)r��ɼ ����{�3��%ӡO����XC�.�Yx�e��}��!�:�w*o�љv?��;t6�P��.NN3w�S��|��*���JJT�5n���V���^\��  +��'�g�6C+�e��rfM��	0�0���e�s�]��lo-��@Kիb����g.0�M�{��ffC�V�N�AFġ�Ϋ���)��z�V���a�6ؔ�7N�s�<ڴ���J����n c⡮�Vwch��h#{�^�2���-˺l���f�j�E���U�{R�س��;�$_DK��H��N��Ѵo+[-vt�T�����yB�u��<�v#�u'�(���_D����pO�/��kn���A�v3rIZ�S�T�n�,�!}���
u$�q_Ί;C�����ܰv䠆��cy:S3�>g��9ܵ�+G���1w+U�9!��ND�ջN�j���T1��� ���̉�+S�����3��]�4�ҧu�O�Ag˦o�!j�4�1�l=��+hc9��3QT˖�]�+V�Dı.�nM�xv\��u����J��S�W�K�<�Rc!����	��ۧ]��31i�n6�szP|ɯ���GD�1E�ᑛꂴK>����B[�,�k��|�54���Z�k�f�����s�k(�NA����AN׍ɗM|�i$3Ҳ쩦Zzk-ɭV�d�I�]Nf��Gwh�6@(�Vp�훢1�n�#���Z��C%taݬ�>����&,�Ŕ�V�F��*jc_m��&.`�#0���2J��	��x CiG���N��klL6�V�����B�.��8��C6�q���:�t5 ���N�n[E>`nX�֤�pe��nr|E��97X�l{�����y�[9a�އpH�w�]�ζ��v෠�5˹YW9����^�Bb,�/�v�8��]c�?
���Z�%*�v-NVB�4[��o�=����tn7)G�����4�r��Ev�d�4γ��o��T�|o�>&N�)B5Q2aWB.�bZj�R��X��;v����{Pv���vmf��E�H�Q�7�P����Hi��EbS�\���5>�n�&M�Eӑ��H�R$�+���o b &U�M�Tq�.�y$�z:�f�Qq����4+�4�C1���w�y{�Ѽ��L=��d�$���$�S��E.B����+��r�3t��9@v�mC��;n�����}R���:p�؞��+���ꬫ��]c�l.1�y����y'�p��������� �m�G��'���~sc���~�c��}�?�����������~_�?7�P��y�Dm���2l���v����e]7�T��Gm	l�+�U�s�h�Y���멅X�/p�EѮ纪*<
;�C���GUj
��)�J��s0�(��J������i{.�%k*��Ab�j���ӂ�:��{��F���j���٦�"yV�S�����*��ud2O�:V�/��5�xΎX1��U3����K-'�p���텱Y������ʕh]h��_J��h�/�"��pXszB�wn0Gt�O���UՀ=�R���骷�Uf�,Z��P��4�Ӑ4Q�\���v�����]�3GY�2�����ij�t0��y5n�ePn������r�d�-���o��]γ2u*�u������&s+$�H��q�,ʸ�|�=ӹ��غ�������돡)j��`Lw.+��]�MV��'2m:��|�c���n��#+#mh����X�vM�&7rW0���{x٥7�����0���V�p��Q�̻%��:��+V-(b׭NMi�[m-=���{Z���jY����f�
���#�q��yݫ]5�4��oq�ײ�N;�w�����{�Wt�KU��\\�u�"���X���m���s@�w��j�]�͓�0�V���G;v�F}�,f܂��)j�\��*n���iL�-��k��x́G���߳p[cZڵ�M��67o;�9��ȹ�̂�hVB����w]7r_fQ�md����_o��E}݁�"�JƦfn�Q.�+�����3���#T/3����E��]� ����w�@�z��C�q���v�WN�������Ful�y%Z5�Q�;�ނi���+���p������sh+Ur�)y�=���8�X��GA�u�w�ME��Ьql��ڧ��wV�rbE��j�4g(�|���_Q�E,��G�>X#*�5���w�����Y�ǉ/�eb3z�b��b��e��["��ط.�eXG��[J�5�}��gSW��Y��:�\o�cA-��O5Cb*P� ��t;�ʈI�!ǣA�^�v�f��x��$XX��Vn��r�՞��z/^a�[)}��`��jʊ�}�qϐ� ���smM�l�S
O�q�X4K���_=�W��-_8��X��~Ñ���4�i����	�5w.3����)�(2���20�Ŧ692�^��1K���1s�⠫o7�1�������f����X��j+�b��
���1V�5��8d��Q��䜠T{m�&�\��R �j�
�~;������|[�N�Rn��Кˬ��w6���bÆf,�y�1�����w[��El\Iyv����,;@�Env���\�yV�j����;[k��:�����V%f��(��)��*���� _V�k�(P���+������f��X�����+�,����e�mGR��ƺ�Cw��&�t d����if�9:�w��W�����"2�뷕h����E���{!��es��q�og*�CYH�T�V��ײw��Y��M�ΰ�)���6�ېŦa��+2�dv�8�y������,����_nGx^J�(�v�mȕ�z����L����
jޫ856��\�,��:��tJ謯�m�ܲ���v�V7B�nV4m�,־��`�2͐E>�5�qjMG�[�Ʉv�e!��v�<��KP��D�Po�&��t�%fͼw�P���wi�F�R�>{Ot�o��͠�&��0�R��m+ ��'T�@���vh�x�1��y��d��Iێ��t�bx�Ð덇�K³/J�8Z�F���hgꝀ��nò�G��	���N�7نCڮ#0�p�H�d���>����Ss��&4a5**.�v���8=�w���(Z��f&��V���.��������jǷX3EkU���S6��L!mv&���<�f5I�S)�+����yÑ�W�Q�![��`gF��qV���M+$�"�[tp�"j�%�F���U$M�h|� K�2d��Z�vc[S��Lڽ��"j���ݚ���	��v���͋�k%7R�)�b����5�6� �u<�ַb�ڒ�xЭH�Y�g�J|���5vm�-�r��ƾ�r���;�� [E�zM.��5�Gʷn&�빀��t��,}CVv����!sjS��*7y���{��2]qĦ�G��YGD�FY�{ftZ�|�+Nª�� i��[8����pҗ�/H[7ws�ٗ/	V;&���\%F,җ��I�u�m�s����l�83A��; {�aWA�ߞu��\��f%���s�x�S�8��-i��+(9�2���TB�+�5i�t�s9t\V^Y���m^M
�L*�1._b��Zr�k28��v���۴d���V�e���d3f�Ѿ�*5ó2�K�Oɴx`�G�,�3,\�ʶ� �쵚2���oU�w�[ G*(����󭁈K��Ԧa�+�ټ�dt	�����C�8�Ko��ji'T���V��\�]>u�- z��J)�j�$�4+��pQ�(dc���%�%���;S��wM����W[{e��u@2>�Lk2l�]^ݞ�|�*���g.�k�$S�YMn�EK���rm�x��u�υL��k%�cK4�N�x�wm����T6H'/d����4:8��gu�B8KǕi4d��xrkIK<Q"���L<of�>��Pf��7��%&.�M���[ӵt2�żyGv�&t0�;��@�Ves�ƅ'*8!����I�%3[Rw�X�r,eD�M[	^���psK��a�)к��ƈu��+A��;�/p	��v�VGy�������T�CwF5W�m���mti ծ��BP�/J:u�u��s�v��k08�F�x�dt*^a�
R�_\�n��]���Y}&P ��Qا#���!��#���M�Le���z��F�М�WD�yG�.�ˠ��f��X��℥����%���"�vMBu3ը�����ѕ�1S]M�h�(��$@�1`y���e �b\���v�u�9P���k^�����MФ��ݺ�t����9xs�X��y��*�ŗ�a�#u��b�.�u��.ri1,��K���Yv�ތJbH7L��Q\��Ģ�\�K�	&m��ڋw��FC37p��3�',:.���fS�ڼ�Э��7����؝��B��<�JuK�E�w��μ6�LQX8i@�7[ĳ�e���xDP�%�J�	��g`W r�A�&i�۸h
�n�C�k$]^�Q�u� b��@��M�fJ��J�ū�ws�[��7���6�*�}%p�{`�1up�<�,ӂR���e�����ɞӹ�l�m�B`�4Ƃ�:m�3��;�7�7H�m�������ʵr��Q��R���w%G�+��@��ú�A&":�0���'V��wS��h�-*z���}��Z:MJ���I��/�{�uyC����H�f��XA��2���/��a��$*iJ��wpH�{��)N�����p[4f��-�Cu�y�p��ٷ`�
˶�T�n	���t-��-V�n���
���S:J|d����쩨bf���bt���j��v��5��L�=��0?�$��_su��w̫;%2�c"r��.boT�3x͔6DE��۴�2��R��a��Ǣ�v9�{�����TՃ𩩵�N�[�-3�t�V�t!�iEǀ;`o�Q�+vC�-靋4�� GSp��:��Y�n�usJw1���Y4S�/��d#z�x�!!�-�-�k��[���1�B�41�k)�����9�H��	0��!4ݖ�QO���)kZ�,i�l�x�[�L5]ݷCn	w�]�Y�KU��l�ngRN,N^�B���iYr�>��0���[��f�.���"��nst)L\�V�AD3l�ro=�#Tv#�,����� R��B��w uWsS�Ck-�}�fQ���VÚ�����(=��L�ѴE���quv��e�V	E΅=v��� T'WlMT�ۼMH+e��NW�N�J�3]�x��yj�񫺄I�v�ȶ�5�+/�c�*��c+������u�[y�I�εC&�B�Y�u�&�m�v7R �L<�.�j�t��Ü�y�m��,�<��M���	w�'.��dp<�d�t>ۧʤ}��0�).V��wb��ƹ�s.0	��M����{v�ñ�ր�"q�r�������W�e*���Kd��΋�Wc��N���8���X3,��>��m�W��aR�*�Q��fu���V�q���ݗ��A�4�Z�@Z��
�J`D 6´��c�ݜcI�٭����gE�Cf�>�\r�|iYD�W��=����*��}��y+@�A%���gJ$�����G!��l�~eR\)���a�R��K,Y�b�_0�V�>or��fv�fX�[x�˺B���ۥe(�3������4��{�uj�iv̀<�k�K�o�%���4��lzQ��d�ow��DH���ԏǆIv��U&e��\R�����'|m񄊨 [/�k_"0�L�(Q4w�g:˛PAS':7c'Z�73$�\�)�hl+������XBbW"�CkV��c5��n�&e-2.q\bf���W�*H���&�,g���K�t�"Ԋ�s��=db�7�	Prp��z��0�ƀ�yDVG�yˀl�۷n��7k΋G5�/kQ�+���b�->�$&��ޫ�IgB��`���#F�&r�N�)\n�|z�����60U�����H��H��l[{�BI]���3C��ۂ�Ks�,f-�v�{��I�+���۪�)Ӻ)�HG�gs�(j�$^��ܭ�N�s�d���&�|(���oB�xJ�O�`�7�ͽRR%�@uXt��B��F�!;mX/5. ��&���\����#X'u��%R0tB���2�>�s�� ��1떓z.Į�����<��t0�f�C�pb�t]o-84��5��p���V�VԸ�f�
�.8�5��B�uX��� kA8Oq(h�NC� �x��X�@���K���W<�.��b�_��/�jvfƇU��&�ٻ[��-V����ٷ�7��
�V���η.)���eB��n,7wxp\}�L�s+��[N�:A����
�8�r�c��7��V��V��m}(ih-�'���yB��n��p�����'T�����I�F�ҼT�L�0�qFt���%n��N�d^f�c'"6s�G�!|�� ueVM����A��U�&��C- m�R�M����a|h�l��u*�^ixsS��oJ{�DG�p�8k�;V)l���b�Kr�!C���vKz���5���ڎ�t�b���qo��3�/�=�����ߟ���ݤ�fk�r�	>T��a&���%C�mC��fmi����|��r��,��NV8wV��No;�;:Ʀnn�9l�bʦ�\��$�_=�<0�)��Rv��m�)Y��mJH7e��&]�ܻS��a��>eiOH�6����	3]�W!v���gb��h�L�ED%qyE0/`�ڨH2$�0j��\�Mmi&�fA>`�#�ؚxF���" O#�����lje�8�5W*h�f�뮫#�!BanD�:��b-�n�L_АC0	����Rr	=�w6r��F�[�H ��n���fZ�Lf�/�:�D%7�năm��)��Yw@b��mq�n��Mb�bVĂĮJ)�hS�]O,�Ѓthf^+v���U�9mv��ۂ�=�dK�q�Ӳv�H�M��yrK_���WWӞ��2�����3/��$��r�}�  ����%��(��"Inh��q�:�'����^����R�kM������(�T)v���3+*g�x�3t��&ۧm�mh��v�7�f7,VT�#�z�ǀ�)��p�[n+��N����'{������<G��'p ���o)V���3��]KheB4_6�l�Bfͷ`��g86�7ˠ����U��{D�Ik�l��*QnS6B�j�G|벹f�8^Ρ�X2�;�-�;��L�09$�X��L�P�}jF��3���OJ�¹��zl���u��+�9BX��m�u#�J(D1����3�fиjPf�,��O!W����۲�v\ї�[���kS�LP�W&H|��c^��6B��Wd,�����^�ᑗ�K���,XJ4+�bd\�gv� �:��o�F�M��l��Օ]���=��ںIX�PC��ÐʗN@v�uevM�=��k9�b���eP��uu�Qۤ��z��ev��w�B�j箵�(	�kD�Z��X����*j�I k�+��3�x�̭��%G�2�̈́��sM��7
�'n��2� @YT�i��<��iV�]ћ�d��L�XZ�S�e���i��c�oMB�[���0.%_Ko�V����37�p�Q�у��fE���z"��H���4���j�a�h�CLT1r��:��c���s2+܁v�`aX��Z����$H_-4�Sɵ�
���R�],�(�����jƠn��v
N��Wlv��Ρk�����T
�>-`Q$RU�K=�Gs;79�\H���acp��u�A�]�ћ��#�IE'vAOALwΣ[G�w��M�W}�^d��*`A���V�l<r�g��R�����Mғ't�N��AJt��`Ú~�˗��v�Z���r��+*�M�˂ޗ���gq�֑b��ֻQ���.l�,:}otI���aQ���`��V�w'���ʽݱ�f�o�f��S
p�]��pɹ�F���� �_v>o�� 6c��.���3��[m�7@�n+ܵ6Z��7!�� p����*m֧��@x�B���kTJӋ�նja�Zh8V�P�#8G�y��c���y�r�u���'HwD:�V���7J�J�I�Ԧ`��n������������oޡ���g��o�������6�[�7�߿~��7����߷_���}�>#�$/w����-{��wp�M0d����,H��<V2e�@�F<��2�Q��*&�Lp0�;�Rec��W��� Pju��:��v�5���㏈B;U�`,�Ui_���q�qNH{v��Y�b�wpv*s`�Z��!��q�w`*�v慾�y.�s8�{`�S ��QN��Bw���0��r��fS���E�9B���Q����ڢjfj�7��|o3��șy����	��-2��5�����<��uU�Ʈ{9<�!��yͰ���Z.Y|�C�>Bs�Rc&�Xjrk9]n�ܜY"� �@\��K4��M���ܽQ$��f�;��l4 x��di#�0 �]V��X�֔�jۓO.#��C�A�uf���v���춸M��o�sd3��3yԙ������3��C;!C��f�EI����[��u�a�����pI�y��g�:T�i.w���ϟg7b���G4�$"NU����:L�}Ю;A.v�WV!W���`�L�kv�m�su�.���52���0���.�(:��9YG�#%��6�+��37v��W�n˰3�#B�;�2��������Լ�/h:V��ӞJ���ɋ�w�$��6�y�J���u�vo,>2*}eIӲ�wrN��
������vm�b�f˒B��8�oN[�A"h ɤ��a��)I.i/]�z8W�=�{������zE�UI�}~>�ڊ���c�s�{���W��"��!7!�Ü��	qs߆�>���~�q���>�^MBS�Ut�n�gQ=<]�w<��tw׉�%�t�o[�v��:�Pp��z�Tg�����DB=뼈qY�w|g͜��W�ޏz�(��>�|C�!�by<�9Zf��]B�]��4S"�\�s��׎��sGq�
��^Noo�+��<v]����a�������ܝA/$M�E4�I��G�$�˹�IY�9��r)�IZ�u�_�w�|VQ���Y�b�)��;ޏW�{���9E�k,E�Īx��'9&�mYeע�:��S�#��y��{���P���D����$Y��v!�����sXR=ܽ?:�B�|�NQ�2���
�����K"*J>��*���J�H��V�ZJ�@�(�2��5��{�p�wi�#���:��Ak��^�p�M��ԯ:D��r�N���&�~D��(�Z�Ǟ�-�?>'W��`� ��!������12UO^d�+0��B�B�v�g;��P��mI���Ym�������m���n	^iʾ�����ҩ�4i������zE��sG��Ϥ�Ɣ��Ju�I�}tU��ϛצh�H:���}�77�^��d�I��g(^�^}XN�38nϖ��o������[��{#��j'=Pm"}C;/G��<a�<�k�F~��{��Y=�V�Ca^n�Ŋ�n������uU���Z��s�������Ǐyx�d�su$�~�ឯzEU�.*r����&���g�
�q���}�K�����>^��W��1��{Y��O~���,nP��y�{�x�߇�57p?l\��o=<h���wr}���3��g'�~��7��M(�V��z��v�;����A�>��O?mxI��=�m{��Twb�md��FY3��M�ҮN��������8����^�>�<j�����W����ޙ��ɞ�g�WA3�{��]3�W~�����	��������v��b�U@�5R����~���L�P�V���9���K6���z��ٯ&���۾� ��@�ST⢵�4l��B���*��&�ϫ	�x���\Y|J����.q�}� �S��,�ΙZ'L'A6�Tz	}x$ۚ��}`���� ��u��d���8��-�ϧ��Ʃ���A
�/*נ��%����7�`�߇����z��R�~�����m\?)u��2��+��R����WC��rD4�Om�ӕ̚��A;�K5S�S���9�U�^�5g��^����þӺ��5��٬�q�^g������	w���mt��ț~5O-e��w1x�~����gI2wn=񺢧**z:��Vf�k�OOSڇ���צ߱��O,^��8�Hrn-���/}~D>�V���N��
���5T��X�]�����R[�Ǒ���uz���<{���y�z����n��M%,o����W���vcnX�~����{����&fj/�n��cm�����V>���{�B̝�}9>&ǟ^1��0Ζ��qdjk/M�<+�/yO6J��ֺI�X��^�����Lu=x�{A�����A�)����H�(�+7|�Ǹ�h��HS��E�XJ�n]9p�y��"͜��t�[u��̞��ʢ6�
�ޜRWce�fvZW��.cYh�F:���fQ�r�V:�6���k���_����z������so��M���j�9�AZھW�N���pl�*E$�w�_���v�7I�Ǐ1��`�MY͐ ���粇n<d������_�x�����C�_|���==�_���Jf�b���Fn�'u'�=�=�1z�]�g�̺o*�����u�&t�go��=����;m�J�R�4�{���K�ժ5W�~s��~�D�x��޼V��_!y�y���$[�/k܆��,�J�'è}V��J�}ǎ�Po�0Х`v6z�{�i��,��s�$1�M3��,f�e�3T��h�^x��{�I�<�S�%3��A9z*�ȯӕ�jٙj�p_3)� �S<cG�� F�7�݃+�sN��&){7�=��+���	G�žJG�-z���®�Y|3_�*m,�si"��]���s1Y<[:�D�	�h��~U[Y��fw��'��ջ�!�r���f$n��z�+�oq��vU۹�C��΢�T�Nr�*��]��AY�4�X��J޳E���9���c��*V6��w�qwXt˛��Nk�]��ʢ&7��b�,�����P�s<V�7������ԙ�Hs"���[���H]��d�9t�O9S�7�Iǧup�U�)H7�{���leSb��Gy���O���-�"�wxݯ�N�����������^]c)���㽞��Q���	�Ƚ�lYG��O3��{�痵�{&�f%�O@i��@C	b挷/S�x�9��0tQ+,�V�p�'���7��ﻖ)��b���`�����[A֘v�Z�8�_���7A&؟7���$<N����^�q��]5��	��c�{����)�׏���=����C;�ݖ�x�t��Ey��r�x�{��.����&�=����:b�W��"��/I-Ͻ[��Iމ��q�&�:6*��^/�.�Ͻ���lHFU�Z+���&gv�8���8��=��rov��#=]l����*=w�ˮ�����':�^w���&g�2E���dΝU�{�����>�p��]��3�dڜ�>���0�2&yr�[�8,=R�c���a���]8��7Q�o����|x���oFA���Emܦ�^>�N�y7A=>Z�t�'��[Fk� �"-�ط��5>��֕�V/�^#!!N�[����K�Y5$띲�s�� �P��4��
ΕF�k˒l>��<�}^}"h�~8�^�r�<���Q���|�K�nA����+�r+��s�{���A��\6M�jx��䖟m��>�������W즈W@��l8z{[��YY�wk����.��E�g��R������_��ȣ��v�dy��������;jW�>��d^��5;z������=_��4x�4m˿H�jH]� Ǎ��c���럼�^��U�����g������I�ͺ�-��۩~��]��J���D��b��:ƙ=��L{T��M�#�}��5�z�f,S�-��v}�c�3�O}��faՒ��S���e�9�I��mgz���c�&A���V��o���*��
�����τ���=(k����MPI�=�L������&��ݲkdQ���y�T�8�����چ�6/��l�B�{�ڮf�#2���h�4ÿ'�Ώ����k�s��*���;�c��*�d��-��n�|U�,*	�A3�:R�(ݎ,���(Ԕ���"7@��\2�P�{8����E�-��K����"}�J�҇�qcsyXlܬ���������-4�����ё�g$X����t7����˧��	�Τ�cϟA���jO?o���������?Gw4��i�ܻ�pzTI����+��5Dp����@���`տN��s��e�/je����0��ƶ��]z�`_y٫��~5ģA2ߧ��8:<t����Cփ����<�+�UO��|�*���g��u�����n#�	yE��rv<"�^[��oY��z>�9�k!�\)u���+���أƻ"p���;�8�ZA� uvh�=����ɶ��eŋ�	��k�]i�|�0c��(�0!�:�����I����H��KX~�2�f��,n�v�� f�M��>�����T�y�B��O��6��X�S>^۶�A���n��
�&��vתJ�ھ85����i{���T��R�>�3�v�6k���zkr0(�g{�c��	���ގ\�9M�c�fΡq��QS3/�5�'X�ں��,� �ٙ]���.�S%pm�j���{Y�ie��Z�(���p���y���������ooq�Җ��=��r'،��D���0O��yQm�f��v\���ud��0�>Ou�}u�����=|{��Վ���V��+��d�{p+ڄ�t�oz����V�y�z�ɚ���1��g����OP���&dH�cR����;Gy����OS҉�7�߾�C�<.z*����y{w�<�S����B��nӳ��FĖ�����7}O�K��@��ruX��m�=�n<h1��Ooz�́��;Xe�����j�O\�?X�-��O4{*��yᗚe��ǈ;gN\�3�6��q�]����������#���g�ӏw�\�_z�{@��z��N�ש�s��I'��ϝ�����0K�9�w�q�m�g7��o��y{{d\�����=9��B�J��'�:�Ϝ�Uy�1��m��8|%����s�q��/y��F{�����t^#x2GB\3b��ʧ��ǀ<;e���0Ȃ���|J	������\���U�:��c�t,T�◥e�'��Һ��S.�ǅ��ә�w\���{��73��/U}���y�m�V*4��&��۰$��n`�p���;�n��[k��G��W�����;x��*o7y�3.��o$Α�zK���}��Od��-�/���~�&ӥ}�5��W闳�
������r��j�5Q��:S�:\��3�B�+�:d(�a�����5�E	-�����䩺Ii�/��A��B�BwJlsu�^�����ʓoƝ/eYo��=�EE��ޥ]`���>[a��{��e�*A�]���K�w�lk7��X�볛7ɷ��#�n�=�����������>�=�	�������{,v|��JR���L�-(S��^NF��W2ɭ� ��5�7�N����n��ʬ8�껽�NQ"���g��_�x��������M�N�%�{��[@y`o>��Y�%=��S8�فT�F�B5�p; fp���t��۳QϜz��M�ګ�߹�y��d{�7D�����k][�׶��6��tC�OV��K��څ:����6���3�M�F��:�Y�\�pq��	��x$j͗���ā�i;ٗ����$@=�-�$6T�ϊč7�xkz�j	��du�m�J��e*��3�F��cf�-�ԫb�`ܭ��e���q��U�T�w�6ΆvI<}��5�}�ӍL��Z<j�c���s�/���}�XML��=�'�ױ�-�>��;�����9�,��Se�}��h��^O9;��,��jz@�3��,>sd&/�k��n���)�;��[g�����$&�Ox%�Z\s���N�yO�O(5�g�����]�� ���TyN�i�V����6�V�ˣ�:OH.ml�l=�=|?K�|�.klo��~�j�Je
B��f.�My�y\כoݽ.�RW_����X~o�w�����̝Y�{���·�jΈ�/�^�t������FOOeCv��	��;�E��E���){���3̬B���'�Ms��<���G��V]�E��P���jz�V��:�X�'څ��;9��54�
1D�qn�2\�H��ʚ��3�/�/D�W���K2��1���H��X͡���/�V^v�^�)�nC�S�s����jʻ��痪�P�A!r�gQ2��%�%��cȴ>�ьV�S��9m�`ʳ�f+��6��i��|���M��rj�^8s��������)�w������bk��+{rP�B�d�b���;���2�w9c��[f����zjO^U�[�j������G[��(qR��ל;����X._j��ծ���\���&�u���;��ͥ�1��h���G�(��y��}����$7�M��	��3�y�J���ٻ{rNޒ_�'_��jC��f��=��C�cr�OZQ�8nxӝY��|��Wo��r_ �OM������9y�E�}\�u3�^��^J���7���@4�ʚ���>�ڞ~>�������}���-w��(���t���{Y~�[�'�G.���d4q�s,��و׽Yw�b�6/ �7�>���S�����ӱ��ϳ�bϖ'��y_�0��x�_w��ϓ��T���������Z6���������>���(*:�j�w�c۾s}�����u9�����c}��H�/��7�߽�W���Q��m~�3r��	JX��CJ��ofl6���:���w4TQ.�4ηI����(ֳA��H�6�`Η�-v)�,@���5����;\���n�w����fj4Ś�3M�1��)���ެ�R>ˇo8����I���n���II��0�
��X$���[�7��%+1VI]��\�5�7+��W��X1��Q���U��WG��m]�����9g���b�\�K,�/��خ���	����kg��4Wjy,�(���,�8,��կ��f>�_f,'�ˣ׀R��є�W���åm�s�eH-횚K�M������2��*��T�4,^�jbp���yyx{�=��1�+7���6GqՒ͈��R �-��;c�d�=��R�,��Su*�r��ῶ�ih@��c��!�}�;��6ޮ�4�	�� �M��G�Ĳ�e��7�A[�t"�0Z�m����wu�`��j�f����gfd�~�EXEdCk�Xf ]=z՗���[3�4�Dw��-Yu�yZ�1�-�����m*��U��9u��8�6za�V_T˅�̕���L�J�6⩗&��f��S	��V��HPɛ@|]�\�;�����;��k:Y�;� #gynG�(Ñ@V���c���E���ٮ��2��h�O������]HsO��W}9�DeE�>ڳz0W�Kֺ����Z�rN�'�L=�=�f5b�9[Z!A��=d�7�;���5u1m7�^�=��� VV��l��bſr��J�o@��к�o.�X����S쉓�\���A��C��^�f�jb3�x,��i1�Jf�w�;����8uh�W��dj�.�%�*)wKV�1<��״"��"i�Wt�ǽ+vq�2�g�\�8:����aǂ�2�j�;�&���T�P�[6��P�I-�{�����XuU�)����'���4�75n�&���r���i:4��
�S��e>����UfG\c�n�8[[�P7�jp	ooN=��G�m�=��.��]�&(>ݗ����kkaFo&���d�_��7���o�=�Fe5���ud��he;Vi>޸vet�M����:Y������j�t����ƶ��Z� U��7��R��uf��E��MApǷ1� ŕʍ��2����9,:0a����	�n!�����=�t�����sՅ�7q�]��#�Xz�[���s41������r��j] ��٥��9W8�*u=��z��{8i�-Ьlvf�o�/��q�*WL�r�1��KE��(A'd=�f^^V%�j�Wq�Ї.�j���8x��oz�j�fe=�*�p�V؋Y��x���]X&<	�p �ڃL��E�VYhp�<���#FN�ovVu��9w�e�lZ���d���v�S]���2�^���-m�KCtJ�&�x��\�g3�W`�o-��p8vf���^�so�н)�ڈ�_N�*n̻1L�C��gD�5�����%t���D���sQO����F���n������:����'D�����u����^<��E��C���Q����_)���N*y�".����!u�;I']�~qȋ�R���E%J��H�|��.Uzn�w����EH,��Nr$<�<���sþS�����|��q-r]i��'|����<�C�"�	]�[�c�f�Z����m\����ܬ{�ڡW���}���s|���,,w��=��O)��"�=<ֳM�.'��z�s"�G^y{>�da� l��PS��NT����5$$��u�W��(�M�����q������%Q>�^OQ��'&=�壛�wn�"�$����)TV�!y-2���e���2�T��]MT��̽۔:�/B��f�t�(�N�S���绎d{�ʼ$��=�=!B�������U ��$��\����DT�JYbHa]�ֳ̉-��rQ{����ҕ�ܴ�K./6���'U�s��V��刉�e"'��O����t�4����%j��T�O���HӤ�3=i5)Su����]g�9JݛΙ!�ǹ��*��Qrm��x���[����W�����6�]���G|�Ⱥw���Q~��@���H��P�ׁ��ܧ���7v���.he4�K@��Wl3i���`�ͽ�{�G�����'����T��q�����יv��ܼ���iiA���X�Φ�Z�޿�+�9�3�s���X9_k�E� ��m�Tx��m�t�,.�B�u�8?P�N�{�V8�앆m�bQ>��,�9���luNROU5��gB�\�q?��qP� "$��T������H���`��AO"������м�/R���q�n��L>�5�E���d�s���|�q(> ��K����O�|s���TQ~V����NHO�-(�j��oD�'<��)9�R)����=���ò�����[ �΁��)�}{��.�����G*�A�����|�9�G_�NN{U�Sl5�q��}�v�޵d�[-�'�R�R�<[	ɧ���w:L�{>(��7�>�8��̰�^Kp�9]#�n1��ˬ����9}.�A����hu|%C�BW�~�F�<�nr�h�2���ר9k�=7|'|�h��i�಺���:js(�j�̽���ݵ�t�U�q#,3\�@HRr ���	yabd�����_Vї|5��u�LIw����:]M�d�T���o� ��8嵄$�Ɨu���\9��K�l�;��vu��v�ЧP���Vp�%'����z�u�˪:=m�wPz�@Ԕdi��G:@���;Ѫ\n�u/�U׸|N�v�"�K��Z̛ኹ��1�(zy��u�ɹ�
�Tr��墝/-�U)���8�/m�r_*�#'��dV����r;���_���+�Ў-Jɣ��d<�7|�������0��q����]�@���q�2-�gH��]V�ǂL��A�!��,Θ�7\b�n=^d� �Ԍ��e���=i�G���[���=���J��<FT9�C���%q�<�Ls=ñ����߂5�5z� �­S�3ν��`�ݯ��ش�J%ߛ8i�t�^���ɥ�O7i�C.78N)+U��R�A@�R>W� �2�P�y>{v�}ջl�%v:"������-�2��o��3�,��n1�J�vtb��tz��D-
���/~�
�����a���>#��g����p�ٛT����y�H�"OP�6������+\~��p'��܊K�x��quƷ�w�*c�/\yyu�/t���A�?z�Q}J�Nk�"Mۄ���Bg�\�æ}����'�.�?9��P�ق�
����{:��W$$~�y� V��Kڳ�cH�X���n���m��	V!�cٵ�4Ayv�W
�aU�=8U�[i�0Kpqcw(
�u�5��03U
��i����º��W0�-}0é[�3$��"�vL�^�'��o��z	��j�p��Mq�|�`r�R�ྺ��u�.nl�ԩ���QnYQ�=X��=�u�z�1����6hJl��Ļ�n����4Y��>�
�.R_j�����s"{B��B��ra������K-2,\�Z��p/n���ۮ_+��p�)(iLFu6no�q_>�2�c���x�록1Y�V�/ʾQg�L�T%p;���-W��1c&�hh<&���o�upO7)�A��k�G�*Y{�4���]��iD�v̥G:�Ct�C����~�/��MaT�5k�5��T����҅u�֑�ϧ�w���&���"�%WrS�]Wf�B�&��m�S��1��3	9��g�8ػ%R�~[�	�?s����!_c+U���Z���6i���ݮ�F���>.	�:׾����.}Ӵ[�I]cp���[�vQ�z��)D�:�J���yx�Lr �(�[��Ȩ� ���P�u��GM���5	�=v�T�K����m���Y��OT�Au	Gk�NrD⠟H��|�����,E����u��s1S�*
�1t��^;˝�إ�}��w_���	����V����,�W��Z�k��gv�V/T�\����龩�*�K�m�f���k����p���i�� ��%��m����+c�V��.�����c�cN�؈|ݛo�mǙ�Lŵ)VQ\���f�8�����^�p`A�%��Q�F f������W�[�d��I��J��@��a�*p�nA�7�EY�X���sɊ͓�c�!���u����+X�c�Qϧ�5��&�eu���1m124^4f����s)s!�L
�Y���߉5MB�&P�P�m{��9Z��
C�R ߉�dM��#����F��*��KuG�uX�u�Q'|�;��6�r�%[H,�+�X���R<nm���/��]S�'��c����B�T���/i�6�!�S=�md׋PޕX�<J�Nb���Wz�O\�m�r�i������H��)V�5P����j��Ѻ��4zs�3����'	�p�w�uuW�� zd��fYs�(��k+RQ��_z�?E,�3�w��0z�dn5p���nb�َ�V9��M�ħ,,����Um�h��_�Ż�Ѿh�j�l:��t��������{�f<\،.�$sb�c�M�q~4����)?2���J���@.�QmK�酹ל��-il�"�*>����qm\Is�ۨ?H��@���Q�9�;\ʢ}����U�j,2t��=��Qʽ|���<˓.Jw^�\��U��%'Uݬ�&7�]ED*R�[ä�/yb���S8�*�aŦ�rV���䧕wǘ�w\H閂��ν|�gI�&�%�)-L$Vv�e�\��3��,�u���7}�>��~xU���|v	=C��Q�H��s}ު;Y��͛�x�C!Ü�g(��y&/����{���1%��(�}�	ޕĝ�5���S����}L��v��1u_W��1��+����y�ӊ<���p$d�qv�w�	ހ���A:��w:��@"z�f���S1��}��ƭ�4y�A�u3��9���`��A6���7�C�s�o�[P��9�e�jzn_\ߏ*
[�e��D_%M�:]\��@�2�!��{e�`nob���I��Pi�hi�,Д/z(nA9���2��u��7C�b[�4>J�1tuJ�{��]]���X�jO�ٟ�PnJ�PdN�j��Z�yr{��I��o�?okߏ�诞�w�.f$�/m��}U7�����H���T=��+���4�����;����:욲7����3�jT�Ɗ*����D��M��mz�+*�s�q���x��=8���4=��nO��_��]�)�Y�ob'<N�_�ꬼ���ױ/���~%����M�YT�emk]�t�4��D����\e�?ީ��j�2�)�[�ۭ���կ0��E�nB��-uq�6�	{��ʌnH�<1��WY�vOgx��4[�}u�y����i��F���� �­gpL�P(�1n�<Ė�&��7�IϠ��HAm,����ٹ}g	ͅ7�o�ef��󄑆@f>�f��l����-=V���-ȣ��sv��s�%U�*N�=�,�0<���3��v����R^58����aA�J.-̪ ��Qi��UWҪ�L��bՏ�#����_�gOV��S���|P�"Fi1�}ȵ�Q����w[�'�{�ӊk2kǷ}Jznl彼�O^���'rABNT04���Xkѕ��g�8;(~�,������F��F�	��W���\��m��l�;��OxTI�a/`p���oP�΍ӢN3�����C�%�e�,�fZ�}<^X��y����E��H��a8�[�7�5��g�B��t��%��/@AR*�Ta��4'��>����s���κ���,ߖo����,B�����z���a�#ڠ��0Z��t��\Χ��֚�%Us���U�Y"!,嗼��I$���#?.��C(A�7�i=��.Dn�ci�[� ��29� �-�5�7��Z'1	Е��JY�?dx.��FE�YǷ$�����~��Ĵ���K�FCEy��B�xЩ[3r͖�nB����482���ɸέ*e��ؒ��s�ƆI���d��w9TA+ȶ�f��i�ڤ��j��<�9�e��Ar���bM�0e�b֏S�P�R]`��ydּ��f'�?=%�w�9�f���o{���6v��}��㻨��f�սr��E5_R�2�b���DC�#�DǏ'�[�}}{u�r[6^̆�tKY2c�E�/vsJ�6�X�&~��EK��tޮ6��Cμ��ȸ�)� ���i��Rw��C�k����T=0�z�P�mr$�8�I�RPwj����;��w�e���Zz�Y�wT�/D^��k������9v�j`�SN+Wx7t+=��XE�b����;^wT��ך%r=l�7%g��~[�P��꺜;혖l�wC,��O׋(^���*D���0��1�����Zިa"����z���}Z��3��>3E�+�-�`�2�֛j���l�j�m�͘}'J��о̡��v��>%DJ��1�U���r8���Ey(:�Q��{gk_�?�L��jKŚ��ȧ��1�Dn���(�3	����iaOѸ.E�qV������Z���!�ni����b����Y�x��J�
�M��*�(�;�]Tk�X��{a�l�^Ǟy�e�v8ɇ�N���h�x>Q�y�%Y�ނ��j2��V5B� ��ĸ�����
���s�:@z����2����|XIwU��_p;�x�
B�9�_*u�m,+�F����Hnl�IP�-]��4o�z�#�u�فn���6u��ec{�q�l���"����ﺶm�N�ӘX��0�|�zv�e	����s��9<?�n��y�� õTN8<G�T�<�/~?��,ڄ���q|�.3k�b�[���r{+�nP�V��}�( |S �s�@LƧ7QL����z�:�e�=!��n����2��U6���<�Pj���v�t��)F��D�������TZ���s��/�\�njh�;���>���C���*���Au	G��Nr�G'�"g&�WҋXFf?Z��#��u��g��HUsQ�C���0���L��f�]RRu�4bP���"c�dʛn#�Q��g��J9鶽�P��0�	���ڈA��	
�`֌�:}��>��sG��=��-���k���a"j�^��7��<�pjY�l�e
��(k&��ui�{y<�*n�(^Y۵w����2;�(�Lw��%fq?(`Z^�][⪛�%��HM���52��:�|长��c5�_����*��<)�+2�>3��>5�!�W�c����9���YL��Ѽ�1��Ԯ��ܩ���Ǵ�c��5��Ve���<=�;�v>�~C�^~�����/[��˩]��_��߄5�d� �zmA�s�1�X�{��*#�@o4��{I�{��Y^�)�2n@T�s��"���cR412���{;&��:m=�J�p�\kd�6�G9ly������KwY�)���x�]�@r��:�ϋ�9�YmS���{��FƠ���G�{�_B�L(���s�U2.sڕc̜a)E�@�^C����"���meX1����@܉��zw��=��w�l�"7���ؖ酌*�1;��M�J{o�S�����m��+Pnt�j�r"��:�kZ}��˖#���f6�Bw��]N��|֛i��=k�sQi�ܣ����1Ȧ�p+��Db�Bv-��=?�w��v�Q*�=�K�͵[:^b�H�ȬjDSܽ���Ɏq�i:�����:Ĩ�L��¦NH�u���v7Rw�_>���,�������*.P�����Ɔ1r����J���ݐ���PcS6.���{�Ξ�=p�ozٍ�ێ�ZORNtt8�|�$���������� [����b9�;ʂvbi����YJ�Y�O흑�=�6��G������׽'�uU�� 7�����MJ>����{��m����emQV/���1m̃ܬ\k"�D�I*�zb�DO1Z��ek�q7��w���(�2�L�<jP�q_nA9ݻL����_.��@g+X�`����j+V"�D5��Q�[�����p^ݑe�}/�J��hn�o���W�����hŵ���N����K��ynq�PӫU�T�19���,*OVeIww�M�zzP��)� B����}�c��>Gv�ѽX�_@�
�U�d�}��U�h���>�S� ����V�R�(7 �5D�sU5z�S��d嚊?p�HW�d�<^��y5n��I�۾2���MP�Ic�u�KT\"�&��U�ɬ`J�u�ӇQ8�϶�l��/�^GL�<W��,��U�^�/����+�x>Gt?��*��ۅ�
��tv��0�:r���,�r6�����]-I�-K*�l��k��u(3�؟�����gb�Ş����ri�o�7B�a����
;ʇtS\����O�x�j��]a�V�=�R}{aI����3�<=a}Z�*1{ߖ�{MsN��0�K��_�j�}"$v��8�`1]�͍��Z�Y�r��{.��,���~����lg�}%�n����\c�Q�t�Q��j�PN+ul��U��܍Ѵ���l�h��C�R�>(��ڥ�-�i�5}������ܸ��옳}��'��jJXFOduJ��BT���]eT��5t��h=���M[��i�ơ4'��{ax���+�\���H?}��}g��}�wʈw���'��!G�-G�mq9��;��f����s���$%�x\�6���¸��#�:n�h6ګ�b1'[���b�;�,k�x�7��"	�  n��6�J�[��������dmg-��8f��]=rܘ�d[,�Y���n��U�!�n^�I�ڢ�dx�*ȩ��cݻ��[�- ra�"���&W05�M]JJ�Sx%�%msf�h�P���ĉ�K!���iD�͇&��L��gd-*�>�/��u�;��s7�j�.�͑*!-ܲ�k�J���zee9R��&��8��ν,k�8@�%R��Dҫ�%����]�Hu4,8:Z6edĊt["�#����q/e-��0��%d!���>�3��Q%�{X�kv�'L� 5]�e�#�D�u7^�Ν�b�7{Ss��3�L�W7�� ���ۻ��$ؒ��q+���WP�̵�\�r�)q�cK��y�fƨY��3KyOՅ^U�2u���,&�����S)��[��R��NS�����U��� OO��G9��"�ǀS��pp�mMޕ%���7.o-#�A�'m�@;�ڵ�����O#mTC���Z���k+^�GTyW���a��h;�{�Z-U�>���G�쫁Kx�oM��]��p�/8N�M�����2�D^C���Jr�.(<֗L��r�B��Lġ��֊qm��h��C(Ay��d�/2T79��p>ŀ�鴾���]��u2f
���/ƥo�։���E>�ｗ���Z�0�u��GǱ�f)���wn^wu �֞�O����^�@ť��#��eu���*+�DX�ѻ�NK Gֵ�P�RI`G&[V�>Xa�k��.%X�UF���T%'P�H�N+k2�1����˖ò��.TF5��d��$ǵu�Z��탬h�h�aAzsW���mleK��.�%e�!m_Z�\@�g���vf����Ub�)��Y��[�%��ѧ��J�V�K(���n�s�u2U�a��/J�f������%�NQk�y�L;��;�+����;Vg������+*Н��.�k|�(����Y��)׆e'��F\w/P������FZx�	��0qy��ǽ�;��`�ךÜr����d�ړ'J�L��Km��.��p�Y�D�7|��Yj���R�P$��k��,#Z�I��Ŷ�=-���P6&U�Rhq�˷7�EK����;��B����@0qTw;1�=��ڍvs��['7��C$Z��clMt�Y|�� uf�y(��)�nW�4IW�yN
��u�w�ޡq��kG0k!X�ݥ�]�uK̬ͧ�DYlLj2~FT�o.s�ra�wtTL)��3J�N�r	�Aik�����8@+u%` y	oXB��@!�O��e��z��R���p�-pG���S_L�@��׀�Fc���tU�`W_8h��J���5��7gH+++���O�l�,�D�����YqC�wXl�%x朵ZkW%�ܾ�S�b�N��h�S����$M�F���:�X����TqD���Z�I&WeQ"R$�W���]�Н���i����1���3.��R����V�$�/'#�5�����ۜ���,���i�H�[ܺ]̴�su�-dg#�r�{O$�rT�~%�%�#>�V����
�T��9����Q�̈��š��J�i�ҩ'P���������T!<�9t��=�W8���sBK)5iI$fg/t-��Z���8[YgPʲ��c���t��f;�a\�Zw��{��P�jP��z`�=�a�L�аȸ�U&�SR4L6w��E���J/��-MM�;�~[���4�y��Bj��A(���L�JL�tr��|�{��Vc���E9����D�"B�FX�b���Q���QG*(�G)P�IM�9�Y}H�*J#�J{���E}�9�"B��9̥)ݤ�fr�:,��vB�(��Ci�Q�A�M*�Y�%T!�(9��:�h�}��B{��P)p���A��r�x�5��Q���Z���X��`�EC�����7'�Xqn�E�N.�a�ؒ�����݂
�(|�� ?�_W�_R_N��`��������`Sּ����J�F<�0� �'��tN��l��B8�;� ̘�3�6��})�\̚`�ϙ�~j��8b��<����\Χ�H��7妄u	U\���q�-㧍�����V
�����q��8<���tq��u���W!�:��i����yd.6l��\���S�eGr�xG.��ȅ�%z�����R<�nQ8z�n����T����>���P�Y�2�.l��~@?X��O�7�d򒚽R�uqJ��"\aܝ�Kf�S@�2,��Y�!{PG&�����6�b,���EK��N�:<ڢa�^^̋X�U�;�%���gA�|�����������Ѓ)~\�6@�x�^{>JJV��شy�x�^�1�#c:�p����Q�i�]K]M���+^��eB�M����ʱ�6P��USw�S�����M�#���7 �_HN%*�Қ��wJf��C=��[�kpe{9��+o�,�����bm�u�ޝ�a7��=��ǩ��g}2�&��>3��
gǬ\IDʿo�|W�@��,F�=FgXފ�[ղ]~)2�o@q�/)a[��Ykݺ����I]�u)��(�;Q��	��&��[0QǯE�&y�ܒX��^q.%����7�^���+SizG)���}wutξĝ]���S�������޼�[�3��_~�S�M�x������ZąWr&9ʵR�5��#�"<�Gi�Fl�B��t�y[l��;.��)ղ�e���t�9cl�ȍ�+M�R���/T�ۜ&b*�od�Ɓ�O�)�?e�m�27��,�����ô-)#juO6(��複pj���ܟ��;?��kNT�ᴄ�ϳ�=��O8�r�s,���p|V�*��N�CO2�k��HI1�QlhLF�h�	���tvq�v	T��nϸ�|�>�%�A�!�g�^���5|v�s+U}���?( � ��j�Nlmת�?Aoh;���^�l=[�#NmoN�u��mΘ���:i��MW܈;ҠGz�5�������L�Cw�gM���1s|��F�GѮ�Ŭ���vD#��'9H�(O�D�97ɨ��nܾh)�z��[)٢5�i�e��g��x��01�@o��邓��%b��0zO�I�$UN7*��k��:�zk%�~q۰q�;�����H�TS�#6Ο}��-���)����t�^V�P#ty:d��MZ
��8s�;/l�E�31�}�!E;̛�u�2�r�Ǝt���t���%�Mۚ$e���,�������M�B��W�X-���hb\�w�(�~l��*��n�y�|i�Qx-�U�/��}U��US����s1�>�}�l	����P(ME���s��b���zgˁ��9LO�N��n�S6����͇�� ��H����P|�Eyu.�4Ԍw�Y��2l���3���Z:U��[�2.Ж�3��cއ��l#��'��;R�2������{�t$ji����O���K T2sC�'�����_7w��<�P�+I�&�XJ��R��b�<#G;�[�^>S�y>��B�t8�Gm�1�U1�9�m���Րӏ/@�q�1X�Ћ;�z[�S��B�;�`Q|��6=ݴ�O��1)��]����x�c ���n�EZ�}y�r�Q�~��8�4����s�pԱv�����!N�S�K�k�N)�>cN�	�D�Ĺ~����ڴ��@h����B>�(��F��g�D��S�dĈ �\���`��j�U�U�0�yԬ�OñPΏ�������u��"�3� D��\|L��R�Y��Қj鶘3�Ƴ�iH�Pb��srظy<k�Gk�N���l� 1�Ljd�ܡh�맻������J䆥���6GY��9�AVVkH���G(�����$Zj��:Vغ�'*��@͡�K��Y�6��աWW�q��lN��ν��[�;8p�ֱn��{��Q%��L|�Zl;5�GpЧ���}�W�}Ү�ڹ����ln�3M��J�v�Z.���B��3��p�G����� a;�,ͯ��D\L�b/>��LJ-cU��山N��W�U�a�+���a�������<�qADSg��IM��ۄ/>�y��dO�༁Bv/��8�������/��u����Z����������t�7��
!��E�D����G���7d���f��)�(㧗�Wk7
�]��f(6�ڂ��MP�)a��܂���.9���=~��#3*�賝�ʍ�;�(��\j+��;BFHm&�.�۾����Z����A@�R��=�{*�݄�a���7k2�6���v��;mS@����2x�%)�=%sM��i�O�0ր��=�Ty��x�R硏&Va�UN�Ow:Ӌ� �Ȭ��{�N70�f��,�y��N��M�~��15dU�������z���@�s��M�؛��w���U��ՍK[�܊9A��^�O'ΐ�^1�>۽�S��e7���,ؤ�k�nQ���As����|��].��q滗�k­)F;Q��;S+�`����Y�;��+-ۑ.���K�s+0�i�^�wέ�)�\�m�Wk��|��(�y��De5*6�=6T{AV�cP�Pm�oEƤAw`��گ_H<�8�Ō�PS�$���cGcٗT�L+Lvq�͎9��F��P8���P����W��W�Ip{�l���9�«�X�j�|z;�������1�Y"�t�آ���7�*[��[K�f�\-�	�):�&�/id��wBP`{h�ZBT=U+��#�*Y�^b���������lf�t�{=s,��%�y<{�E���Ա�9��k4{#����!{�S�ּ9�;9���n�*D���M�z9r�S�K���Q�1��E��LF�}p��o��ckLt�`��'�y.Sا�y<h]�Urq�IhǠ�g�tL�5a��_cv_���%=����|�8�Ԕ|?.��ɡ�a���@��C�LE�o��M�u%�KZ��oETv�'+qu&9ǁMWڈKJ�"nY�}nBv���3�vk����S<�um$���Yz��^z�;rj׳Q�t5N���Y(WP��qL(�b��#FG�W�<�e�i�d�d�����]�ɺ����3#R��Ԩc�l���E�j���e^5������{�e%�^���UM��'`�+����fW���[�	��T3�Y3�~�S褝���8�1R@H~���=�ߙ��I��M�F�^�i�$3�=���M���ց ����]�0Z�=��������=srvxK���g��S��9�yk��\�9���]�'���Ev�He��#�r�ȪX�l7�O��|���b4���kd�Ϫ����r��TQ�?
�MM�Խc�j��>�S0����`޸}n<�o��AI��y콍��j*�E�f�0�_P�nR*�"-\&���ǚʛaY�V��0�(z�_=�wB�#K؞�d�3q1�r3�^�D�DBۨ�����QP��>�)S\����u�Ħ�%�.uIlnu˺�+/od4]��٨f,�),�{h�닽[P�E�;k+��}��6`����y�9v��'�iUT����h�wu"������~�{;���+!P��
2��-�V��!�n�P�J�����"ߛk��j;)z�3!�d�c���,u���>�r�xuM���Zn�J��u�`�3=M/D����Ὓu�:3��`�UjZ���B���ȡ�R�5a�K/�F��r�
cJK0žu[#���Q6 /D�c�՞q�,���7W�&����}��U4e�x��� �6�c��ZI龢��mN�x������ex�M$,����ML�Nv�ݠg@�J\iޘO���e�#T��[U]�p�1T���T�q^�2_���;�
�	-f�3�xTQs���|獲L!��P��f]u�|m�����U�O
�j[ƃ!7�B���VfL��W��ىg\Ε����L�����Ǣ��q��+jl0�gS�ы�
0�k�����͍`�C��lr�.���y��W���nCZ9RGK`ҹg^[��eҌ�4�]��Z�Mf*㧆�+��/���'��wA��ٿ�� ���+#�{D����{���j�"d�-�bdT��v�O�e9�|Л��O��xq�:���s��(`�=k�e�I�-^sBQ� �� B8����Dq؊���먃����q��F�=b,�nui�� v��_]�,����T���+\�-!�l&�-y�*eə\Ǻyx���=8С5s��[�uY��Ҏ��ir����
�`�,��6������ҍuff�Ӳ�70�eDI�i��W�	��\=��'Ě����?6�p�iW���1m�9����Sn� �jQ0��Pl��DdzP9��s4�Q�]����aQ/��Ӕ�FU�1!SBdTMЬ{�Ȫyt�H�IY'���\��І�^hs���iˤ:��	�W��2*wj��X�.���T�sx��u�om��av)n��е�<T�ڐ�j��y�*�-͚r��(��З��&����#�e2�J��s�T�uz�V0I��^4Rs�|��Y�ܸҷ5��~+��&=������/��i�K;���9:���d,GJq<��U��&�m��ٰ�~�%`	&�m��*�X|H���+��G$n��3�K|F��]qk$�T�D�5|*J�4�n:`�t�B7(����>�R]�a�����1�119ّW�+�:΅[�9륮�l��&�R��?�U}���-C�~�;M�}�0�'��;kh��� &�/���mC�4����)?4�+�e��SZ�C�)VǷ�rs{ǻ�-q}P!j���_y�K��)�zV&<�g�C���-^��*`́�ə�����n��u�g�l��Z-Ǌ�C��I( S�:�+�?�%�o4��ַP�"��?a;����3���Î�]�w^1r��@'zTݐ�˕&sGPs�x����v�O%^x����;g�Z��?֕[ޯ���8o��r�Wl�Q���x%y�V��9p[I��=B�X;�/�?<�C`�2��3�;�^��+S+>;����gr�c1��<y�1z�?^����	�0��
_-�qv��M9��(�N�44C5\x�m�\<��_.�u4�DO��`�P2Th�d˸�"P�8���P��3�oi��+�rM�?K��y��ǽB���H�>�N�֘J����W�A���f��Y�z�]���h�2_9�y�ݛH�wO��Ig9٠��)��+u�"�O��Z������n��d9Ҵuŗi�%��֬�C;b��ꋑ¹!ZF���J�s�s���s��3ɑy���Sp���y��a��*r���+��2��r.C�d<܂�뇜��.fG��[��Gð�G�j\����8�b�J__ʇ>��^Ӭî��e�s{� ��M����܉��|��Ṿ��|�0Z�O�YR�⊔ͯI\�e�Z����Up`OF`��t�"�����MwREȦ9`T�{�^����xX�1C��,盺����V=�J	��z�D�t	�~���L�ix�Ma�8z�>�	���'æ$��1I�|����m��H(�t��x�ʋ�r��G}_�褼jy�9Y�����N�j!��=���Z�+�fmOaj\�2�a�����8��Tj�cV�NC�;��x�4�}����r�`��d�����o6��n�A��^OݡH<�H��I�ʁ����ZR��\�n��|�]v�Y�����iv��z�s���������R{ F
�0����:�2.g5[�z��]���Au�y�ݺ�<�;�46�zUu�Y�����T}\%��E���#�vz/�-{�����"Dln��Wr�U�o@�|���q�w���s6��ZКg��j�We� �>]""ɀ\qS�\��6�(T���Ōbq����[�R�E���$%=uU��ƹ��u�(Ǌ�/�Ә���o,_F|��N������Y�z�m��)�t[G3�ܧ(��@��r��R��#����zB�Q��Ҳe��ۭ�:��u��iV�e/�^kkS����5"ĩ����:*�6�}U�}�N֮ޢ_d�n�#>�4Z��Μ��ff���������w�G��;u���Zn�U�b��<�7뮳�5Ҧ����S�Cΐ�}>,������hY�險Bg��W��L���`�gI>]�ـ�Jf��r|��L�`�aw&�6%r���@œ��U=,�/s�~S}�ޢ6Mx�ܸpB���N؏��D����(kL�R5��yԢ�O�u����os=j ���/�z���εR�У��!"MK�لC�PCo(מ�8����s�٤�m����Y�;�[�2���G�q�U�f�6���y�l'Ϛ�c�A�9�ΰ�³��'�fɰ�kFk�B�XE�1
F�"���7%w��T%4sU�û
��,�62eEj�K�d_W{��e�n�������F��a�L� 1��gx͚�W2��q+������ć�ﲟ��[��ko�>���]bS�M�j��"���Y
�bB����+F&W��0	��Ck��\��,Q��[!� ngPf��(��BN��Sr�{:��f��9, ��T�߷��}�uE=����K�*�dw�|�n��YY̔{Xb�[' �]�NF��Q��4f���T��o,Պ!�e7�����=�Z˾nt����B�p&eZO�Ν���7RR�ulC/rt��;c��J��gSm�\��=�Aa��o��,�iM��a��Q�D�	�s��$�ͮͷ��4��C@��L��Mn Ĳ��1K:��BB�g�9J�ކ��"�=�(Ff��bly&�I�`+�7�c�Y�Cdsɏ쉭ҷ �B�}Í����%����\���߯1�u7�jk�b�ժ4��5��)����� *
�ޫJ��L៵��w��P�L�5����$%\��`4;��Y[!ȋ{s��ru(�y��^�Zh?�ڃ��WӕK���S����]X�[ׂ�r�o����gY��B���t�ʖ�t�fǔ,=���,�+�2o��GEom6�[���,�M��]�����2�L�]��j,���5�Z
2܉ŉ`�l��˄�,�e�صT�\�`�][0��^�JYaДf)@	�]�8�uk3�B�e%�+��v�fY��9wQ������-��i���(�k>Up�EX^v�����lHk@�/��co3�윮WwӉ��Wc(�\7(8�L,fˬ4�C�>nX�I�Kz��[{�n��	�2�P���{��R�r���tN\v�Eeub��J*�R�E=�YZ�u�͗��j����P�	F�q��z�N�#����WF�\�s��9f���T[�d ;�]mΆ����0�Z�r|�"cΩX��	x
r�!pȖtJ$�R8"*Y�x�3(܎�	I�n� (��M��el��nWg*�eS֑6��xS�N��n�E�T��)ښ���e�ըт�h�;�(�W	��4�7n�o�)�9u�MOf��Q1�f���kEk���|�x 1��\����!��O�u�P)��c����(�%�wf��>j1Ӹ�,�vw��>�i� �͵����W�p�T�6�����d��J$�3��Y�(�.z$UI�����}��G�9�t�lfkx��jQ��P4�Jgdyj<��YI�R!ˣWt�V�6�ҫ��	Zo�}�	��P��`qJC���I���}8�]o'o�G���E�(4�74���F��5a�;�q���[7u ��\�*\Ρ�#5.:]r��+$]�n⋁N�=�#��K���HɭȐR&a�~2qg��"Q��������L|�����ee�:��-@A�f���-���p�烛���Аt�Й/`&Y}��,�&,<`�2
��ĺ�fKܩq�w�sW)5�[/m@q72����<=��Yd��*Чq���C�w\xs�D�O�;��"s�*�E�l���1�(k�MwH	���w2R�`��S�J�s�I5�W��"Ŝ?o�L��@�D���N'4��=��V�7l���az�����Qh�<�4�R��K�D�I$*�!*bG���!������Q$��Z���!�H�\������VU
��b�!GJR�hА��e���2̍�c�w	
���qZWy�A|������|�8�
O;��)+v�2T�W�AC�s@�4J����		Oz<���!E�V�QE���U:���E�P�$�dEh�H}nEUz'�sı� �"ʕz�U�ĮUY���W�/,$�Ng1,�w2�D3𧈥��F��C��نIºA�Q
? �)�
�J�h��O��w*+�	Djb�~G=��NXY����S
J��݂z�y��'#���+ZʣG�=1��]D�uL�l�GT/�xN�j:.m瞪���k�Ds��D��P�P�#��O�e������?<dv���տ��6�Ou��`J�[a��sT{�$�a�-���u�9�@ӝE���X���4Xb�9������;� ��O�����=K�S�<��v��ن�3	�{*Y{lN������-b��������qI0�*� �u���0�UjuH�jEP�}]H{�Α�cNv6�u�{��G��z�U�T��I��
� P��$��e,ZdL�5Ҿ�������9Tu�ts����v'v�9�QN�0S����!Xř�\�;��
�	��f���NlTS)�:U�v��\��lō{{�y���TZ�<S�ne�-�)���z~ȐR�@����C LaB�z1����>�������!ܬ���ZcOoޮ>SBQ���$N#��
	������^���	�z�J<�����}��O$;
�����<M��L�꒓p}Hx�W�ؗ����9��=t�Z��}p]�v��Fr&�q���JHH��p�L$�^�B���Fs�2�au�����9�V�l�ŵ'$�B7��u�ȼq��n�Q�^�e���z��:Fd��z��罵A�*�9]Վ�䛧a>��B���`8ׂ�w�rX�����qj���PyL�t9i�:�m���͑:�7M�>��9�78��Ô�S�CW��]��&��_Wa"Ṵa��7æ�&|.������v�;b�%���;M�%�sK�[ʌvu��{��k�{F�����m���U�{�32'V����x�㹬h�w�lo�<D��JBm��Dڡ�~�B(�J�T��K��B��Dk�7m�xz�.��{z�w{ܽ3Ӑ�d	7���)��,_�b�e׊����w~�y��O���PJ�mH���SFz`�����v�&�\�Į���rGh�%�1	�pJ��s��۪�V0I��M�ݴ�x��Dھ$e�7=�3��7L=��dp3}�ۆE9Y�ZdU�����m�fߵUK�a;�Wf����Z�M��_b5 ��Ҏ������!N�S�~>u:�|��r�O�����ΙT[{,����M|�"�!���}�a�G�Ğ�/q���W�Lë��v�6����!M$��	tqč�X��j�Z���|^�����'�g4���D���]��/^�����u�>>�Ԛw!�kN��|�O�.Q�@��@�an�B�E���l:=�s�ŧ*Z�WQGM}�F�������A�|�OuV�
�OAO0	�ʚWL��y�W.Ⲃ���{�喫�T�������i����?�"6H�Ѝ=o�t���c�,����+�qL
��g/��&�2��f�<�	����R�ѐ�3��im����D�s#8 ʱ�5��HZ��|�9u�/+:G��d��3�;6��tes�J�}K�����޵պ6y��o1�	HY�����e�ʡA^��C������U�A�6f��Ԇ'����ߐv��f�e���`W�(����mrITN1�:�)��oDq����ru�v��7��X>�G�P"�jDgB��<�t�c��aQ�P���zξl�&�V���*X�I�#��MwV'j�xځ�$���P��&�T��R�`�Tk�٨��g����E]�l��smz؁�f�����1�დ�Iqр�T���T�:P'�,�����# �����0�m/~#��͚��}Ư׊>W,����c߆��a+�q�+��o��ن�CYۉf�0��
.��*f�nL/�VU�7�ݚz�Ld
q%��Ϯ�����ёw
v!N�iN(�}���v��(,4Ȕ���6�
��+ &SY�t���������5��ظd��C��������}7k��^Ea�Y\��?q��h	�(�\pk���\NN�����yD��rOTq�+1����/jV0��������{=EE�1��ˑk/Ѥ�n�ĿƱoV��ge�w���PQ~u�w�Kд��\��u���pdy��{�od�����ڧ��L��/.>5:[4�j���>m/�>��޸���z����}Nm���6����8t�c�I�$�j�	�rm:��\^�o+���;�g<6���ST�fQ���R�"Y|��N���O��_}_}[�^�]�f:�|�����5���˴�r�j�r��W��;�n���OJ����0���s���7��0r�ymy�r�گ�N��
�<����&^�\���FK-��"R��ZL���{�}��s�z�6��LF,.����V)9�=��I������g�~��dK��FܗÙ�k-����~��"|L��*J�Z`�j_p��p��!^�~� �vP;\hy��W̾s��ٛL��.4�L$M�+5#*Þ4%;][��7�ޒ2���B�ڬ6u�uo!��e��v��N��PHɇ4�="��r���@8�'��j�8j�X�B�����cz�+�ם�x�/v>���W�ږ�@�~�h.�)��,�P'���n�7�z��os+���Lx�Y�}������ȍk���kd�Ex>�$���ъ�ȘI�ߴ.^l�P�o.�E�����1�a��]T,�.��p.��ng+�bf<q]��N��z�c��(3u
�%��_H�nnz���eM��f�Z��0�(p�\+����n4�({V�[�t���V@u�R��PK�Ne��Ā�.���Αu<r����`�V����������;EMѷ�Ó��閭��2J�`�.���Ȍ���odцWK�VF.�[�so�B���v�ӝ�4����W+3���F:u�V�67�r��T=�����5ג�Fg�O��P���u������mB�ҳvWy|V�3N9���K��s%/U�1���^�E��{W�����P���u�ޭ�a"��SE��M�١+�B��q�:���vfVV�u=Ӎͱ<���xǏr�b���e�v��l
�T4)��Y�Ƿj�L㎓�2�r�������CA����t�xl�N�<S.~�%>��X�59�g�D�ه*7�[�o��&�<f<���jS��/!�݆�f�)��l;}��T�r�:j�/E�<�1�����E+;r����/շ��_Gb:�W0��nz(����p���b�L'D��
����GF��	~>ؾ��4(�r�dbl�6��zÈ�Ւ�׎�CT�7P�79�c��9��(�Z�Q����e�����s5'��[r���opv�=po�d�L)���%Μ���6�x?/ɍ\���J����>�+3+���Ӿ�8y����4��;��+����*���zD#��W �wn�T��z��';��������IV��R��˔�7s�7V�p Vb�iL�����~R�t���V��٤�ZD�DP^V.�N���C��h-��4�E��@[��ģ���Β�5�������6fP[��e��f�������'y���<䈑9?�K�>��n���޷i�pq����z����i�I����ڼޞ˂����Y��D{`6)0��Md����$m�҇����A�0o�ֺ�s�3=�=r/�Y�	\a���QMXܩ�N�E�"=����E�����fZ f�svam��n�,���{���m� �m�H�9�|�Vz�	��D�¥��.;ʄ�����/Yw��>��8'wm��vL�/�P��V�&�+�X��Z�*��<<���ix��x�C9�{|B�nn���3�U�}���՞���sMo�����Y�.��<<�[㾧�d��]�b�^�ފ+}��:)4��U)�7W!�>y 莉,(fS-��S"�=�m��Ͱݼ��ˍ�����2/k7����'��V�0������v�\#]>^�Z�<:�wcq����-:�0���f���8�t�]ﺦҳ\��Ɉ��5:!��p���B��z� �1i�1������943w�w�1Og&�է�i����Z|�"��9��Bkj8��7Z��
�[7=���f��Ѐ���^�,������<ח�۬ )y��
���v�˲=�4��"諹l����ro ���DR*�5򚎉��0����OU�N>i�R^�5������-\��+oK��'ó�-Wl[�:�Yx2n�j�a��Z�͵M)�����������}ǗmW�) ���Ho���+�P��J�=�D觩��=��䗍�� ��uJ� ����`�((��s�;�wh�iCn����jj8�KQ�
(7u�\<�5�1r��@'zTѨ���K]���7�	W�ʞ\`������g��.�єW��I�֠H�v9lD�Y�3�<��M1(����P���B�5?nV���#�;���T<s�l�޿cT�/4��N�/!ʥ��P��"	�ˈ��e�
_*�qu��4�H�E���h���]o=�n��޿ZL�C��#�AD{�F���n(-#ҲKT� ����1�z�Jr��uZ��A"���oE��X���O�F��>h*��&�j���PnJ��3���W�c�LF� ��7������}�s2�n�b��+\�,�y��5Z�,t�N.�oƧp4��(�ud����j����Q�<��{\�[�KT~�9cVӰ��o�\V>Δk���4�w�u�~ǐ��]FH�9~�<�ʺ�tD�x�2j�ɵ+�loW_��Y��u��{9b�t���F�U�A��Vj�I%J�-��`����t�-Eo���������偌�r	�c��%�p�\f�#����o]��v�Vd�潝���������������+��9��)��M܂�Y=i?�_}_|c���-�;~����w��-�wD��X~�s�y#up����GZ�R�ģ�b�Eel{-c��[ȣ��n׏�<��W��:#���KrNUƃ��x���u���f��
U:4-���7Ns��&��y(���[��cjrr�v=�@3�0r�=~��WQ�ǚ�r�9�cMn�fC9T3��wx�5���:�O��J�/id��YP��t��Dc��wm���ޟ���ή�<x����:�xlil�;P�3#���8(���F}k�We�u�r��9\��5u���x�޽/GC�c�0,^nFԼ"�/<��5"9��T-����w)�=�L�[�'���ɕ3����߭�h� zR���#�`4�i#�yA�O�
U�nw�{',���Y��*݇<6P�_�m]���2s!z=�s��W�l���AKd\qiC�&��;LW�='1�G�*XQ��W�������=�B6���Tq�S\H:l$M���Ԍ�nx��������X�R����<���ۈ%�9=�-��Lp%䩹dbqM]BW*܊��!/��!:�<�ɼ���o�q3�yh9�6�,�l�Y7kSY��fTC6���4��M�\�Vń(��u�q���Z���N�z�ҫ��a��ч��}+z�Z��*cd�ĝ��j$ub7Zh�+��v��\�Q��<i�����M��v�S-�������V��u8O?Ϗ�ݠv����uzI3��e�9*��I�g��,��tQMi�����Է��wc��@�%Α11㼳�wFdR3��
��q8�b,�o�C�u���|�!I�1<Z��7��ݓ�^���e�[+�@��UP��fcEB�o���6�.�Ū��GsP������6�=P��=p�^��p�r���u�����E{�l��ɓX5�S�v�[�<l6K�b�����ʵ�5w1
v���74��}#T�MsJq�:x�`b�(fռ����t<�\a2/x��������;�*�,�a>��y��Ѧ�q�;j!9Eav}g����W���z�u��!O3t)M�L���Эy�}CQ��{lw�!!v駋���f�^��r��1뀃m�ǹJ/nfRu��m�s�Q�J뱚�/�5V����kM=�����b9���*Qf;���uP�)���^���)�3	���\�}�j�nm�Ω��ڷ�i���ܱ�JwWL7�0�pvS+ãU�w������ԝ�����ԝ��ڨ۱��{9ѫ���̠&�Uyv}����N�+tm`���I�m��2_l��-7��A�cB�,R��)���(���sy4�Ո�X,�Yg�x#.�>�3r��أ�Ւcޫǝ�°-��v|>�A��m���E�ޑ���U}UUUهݹ�N�W���K$�9�P�ϭF� �i�����-<%Skߏ�����u�1=�m�v�廷lc����Hnlc\�7UA��B�1r�W܈;�
�	-f�qQ�h��\Uz^l�OF*b��H��-��'U�Ĥ�A��Z2����I�X9w���aM�������u��MP�MȂٶ2i��j�[��qD�k>���?G��2<��5;�B���31M�;[����/`Dt^��ya�#�ݪ��� a�^r\[4�����v�e'���6m�_��M������D(���d���]���݅p�'r�;6�Te]�fNdc�Yj�[�㔆��Hb{g��⚯�abiA�k���SQf��T�ac�2�&&KE��<�]��1�u�E��z}��#X�7X��
C�R"F�#}AD��W5�@E�yb�w[��%\u�0��E���Mz�+�j��s�)��۩���ĊO.�-�\�	r���N5���+�+s�Cg��*g�p{k2�ɯ�
q�ĩd���ղ86q��
�b�зm�׼��������r�y$�J�t簮��
�G�EE�1t�;b�ZAP�Sa���|���6�q4��Xp��0���`�����5��|v`Z���LIշX����=`B(^�Tgu�Υ��uʱ�T�8s�x�Nu8u3����D��P>��+j�N�q"��+7^�n��P�I�r�J�,��͕����Y8a)
JfF�2h}�Y�7�Сcn���-�dW����ֵW��C���C����|�7zGsX�el5t��w9BZ\nm	��գ3.b�V.��4�=��WD�i�Kf�]�lmN�`յ3rbt2��1�S��z���=n�Q WZ ���gDG8�[5�3�	ۡz��m1�B��)��+�T#'9I��{�fv:�[t�ߥ�8>'^=���(�pl��թaR�Q��oZ��vV�Y3��t�J�@>:�2���݀�.)��:ш��8�v�͛0� {{�zGF����۵,�О�5��$�|����"��`=��aO��e��b�D���9(iz�ղ�B\��K���x��{�����t_l�z�כf�ͩX��q����t�8�4[\�����k!R�tF9��t[]����T�ݬ`0k`�:�[Go����mJ�"����+,+�Q�L|z�@�ۋ<��x���;X'�=쉃��&o��S"��L{�vk�-ξUn�y�ꛗ5!-6�8�����OB�C7{Ѝ��`��k���e�{�v}oxp����P��F�=]u ѶX2�{'�)�h�
\tb]��۾j�C�V�h�����S/.���e@�Z�!?��0���xq������r���<�*9a�l�/B���o�R���X*������tdw��(��	��N�,�e����\�۩�!���7�l��鮤��hq�,iE	s7��&�%2��*�!�/vq� S�fS�{�݊f͂ʳ�nA�>Zx�.}�g	�)R�w�T08�r��7�uf҉V²���Ål���0����W	u#�x8����(J�J�'��u�ܓ�u��|�m���1fb#��w�� �;����ֲmw7ԫ]g�n��H��Sh�O9��՝�$��{j�L8��CX���Hb�m���/�Ͳ��\�b)'8�u�[������׹��]�A�$7jn������:�ϥ���#Dr���]; �`ζ`�E�2`xn��>��Jˌ��ae��Yt�]d�_e�0��ޣ�.����������n�U�G��i6i5�Z,T�]FT���E��e��)4��fB�R	V����i�YlǱ:e�n�p��Cou�Q�؟ٷ�I�Pt� ����Dhq���Հ�*��x����9�ؽ3���GY�>��������sVz��s�O��x�#�s|�,����w-e�BflT�_]!�R*#΋[S>ˠܣ8��@r%�r.I��މ�*��[(�|\��9m�t�ut�{)

C�>B� �@O��̢ٗ��K��td�t��$��#��UG'���*��Qa�2���Β�<�,%֜�8��Za)u���\���gU���V�����н(#����.P�,6�J��8��rr�P�YQBA�a\�U�r�r�I�)Կ:G�jI��G�ܝ��9*p����N�v���������-���(����n�4��"�zIRe��<�">L��~ZW����f Aʤ�UU~R��i��r/?.zVVl�Ȥ��D���UʹA�E��*�K
��(�uT�M�[HQ3.QG(�T�w�y��J�Zt�Vu��<�%��q�����T�KQ9��BC �$es2)3:J�'J���t�`F�Zs�R���U6��'ez�'/�Yq��kN���hr�r���ZAG{~�w�x�����8���Uh@�����V}5!eJ����bۨ��۲%��) �]�-.�Wͮ���ĝh�
����.u57����U}UUT�GWY��A7`��1D��%�R���	]�]}p8w��8!ఐ	�L�%Tȹ�j�n�ibL$^�#Zg6r��.��?���ǰ���Ӷ�����<�.w�P��O�������9'�-�u��=W���6��({��o���B� i@J�G9F�ptݹ7ax�t�1�!Xn�gޣ��w�?�����k��ӴܼZ}������T}�&�ƣ�tu�{��݉����
�#��� NT7�na3b<9δ��V����@c���΂���$!���X=�=��9N���o��BJMS2n~�������M;��⛍:�����;C���l�^(n��0��yy�c &��Q0�q�Fl��ܧ��.��y�[^v�	Uk*�#��9Y].�A��_)�^���CF�A�d@F�`O��^��5;;#}��m]�O�l�6Z���8�9���3�V���5�3.:	��NAq�H��	/�nA?a�����5�ٻ�w��
���R��,��ƕ7�3�s�tP(�I�PM�ň�]��=� l{Q%�o�!�U"���aоwF��:���:���n��|��]��vy�������j����Ψ�SDv$Kt�7�-�T�͛�>w%�}��v֨��"�	�ؓ췇D��o%Q�9��˅v�lబ�zFh��|.!L���y@�������݋9���G��mς[i��%���5���H�<��_Gz�U�R�?%��PR�>��e���VV�k�{�˯����6|�#3.�ۼi�(�0w�E����/�I��Ic9�;3:nOM�\m����;�=@��!A/Bj<kr'�>�q_O��j9d��Q&��wH��#����S�,y���ݞ�a�J�P�v�?B2E2˩3���<Ωȳ1j�ɵiu�b�W�6���X�e[Z	mk\�r��*�q��A�^ʤ}�:�&�M��o�1'5�l:!�������Gj�}�%�/b�M��n�6���y����8F�2t����S4ƈ�s����0���;]N,�Z��NN{U�X�Z���=���1��
i��j�5<�Sn���F�gI�d���q���ꂎ�9㫠>pZ���߃j���~���r\&jc���'k��V?bĨv�V��~��}�����8hoz_&��^FB�����=�;�I��Fܮj��5z�kԐ8D��X��r�ϪD���E5{�ɗ��)�=�d���3/�.�XSx�c�QV�ɏ�;��^�R�x��8�u�7�b�u'�m\����i���U��弮����$"�5:���F����������]uI+��|�	e���d,5��Y][�2%L)�gB{��F��f�ģ�V�J�,��r���ˡ�݋$�W�U}�9���Ҧ�����"]��ٻ}���� ��y������B8Ȫ�­0䵞�����6f��v�8ݎNG��Fk����e}:ųd��ҁ��҆�E�kgM�
D奈��^?DT���co���7H��{"1�uZ���)��:I&�Ԍ�nxƑ�>�L��b7g0j����'��,���Lq<,w�����)�*�k��z�Z���?[;�
+˫^�h;(��z2�ڧmcǧ�	3if�Է���l�E4Xݣ�+��k���������^[t�2��r�}�j(��ݞ��4��#��M�0}��G���=݆�>?{��[���>��ʫCƆ]<���sX}��Ł��zF�vW*���[�m��n�� {� mN���J�~U��ܨ}xԺ�pl ��I�y�O�~���忦'ˁx������Y᮰ɢ��B�H���
�/�-�J����Z��͉�Z�R݌:��ɮ6o�=��KW��C���5�ߣV�0�{e;�� �|�jv��\T[dP�(�,`XM����i�������Y� �Oeb�A�Xgtn�GDc����0N��:��t���S�e�?:���*CsZ��[�ık돒��&nq \���M�g�!]dE����m�q��E,�(&���Wӗ;����PX���ꪭZX�^^��\�J�$+&7�XY��3���Ck9)�&�%���{̹H�w9�E:,��ȉ�����Z�H��*�J��h\o��7\�^t�i���Y���=	���G2��h����Ȍ�/쪀��%����S�-u��,�ل�]�w���j�QYku�n)c��0ܻA�Ғ��~U�DY��o�vg��cV�"�`c%:�m�����6�:�vU�����Qa~,��1C[>�X���� �v�8���{I����K����=A}^�	�b�w*R�l�P�q�����ь\�T9w�@� � �6]��ǜAc�r�S�Nf/��=)�|I�cRx3q�(,�>�T�Ԝx�L�w�Nj9i˟�������0y�	��H��ξu��v�<docZߌ�>�]C�\j�d��苨�U_���v���\�>����t��97ʀ�Z�&���s�GD��ڠ_t �
y1.��)Ԯݨ�{�S7�fɂ���%b��#�}"!��>�kw`�7vT< ܄��=
.2��9����"�
%m�k:nP�WJ��6*vB̸ef�Wj���7N�n�ūXPM�Y�o�±�J��{2'��K=��6��"/R���w#9��5}B���ɋ�q4�O0
;8��[�ɼ�������E���e���<�]��Q7V�#QL�3l��]TD��d��@ɨÑ{:��V��P��/Ps���W��ݴ5�P��W!"o� ���#f�ȓs�\׏�|���a���a �ٽ����4��ꭕ�J�8}���P��6�B�m��˥
uRVL��<��mJ�U*������7�l�#��@�Y�^-�
q�P���K-X��U�
 	���{d&�[�s��}�U����G^��@���U���}�u�ँ��4��<w7�Nٱ�T[R�pw�Ԫ|�����v޸8ۺ�+z-\I�`Yg��J7S���#���
�����&����׉ɉ�9p��WO�7�5��_�a����b2�j�a+ߑ3�ԙڸǏ��grvW����2���`^��n��[�y:u�ZqMi�{v�9x���EBp�X����T�ȼnn�@��������`����e�����NЊ�u�{�ܟ_�$n*�+UrԔ r���!S0�Hl�!�ո�/�}	��!�=�h���J���ƺ�J5��d������vA�}�e�&���+2L���.��Q�:�5.���t��,SJ�;�Tz�o�UŔN=&�%���xnVVK�[��ѹO�t~k�u�ߒ�+������o3I/���2J����-��x
�l/eX�E����gT�
�{�pq�B�#�wGy��}�{í��͞��3���G����7���^u3BT�2 �ͯ^�~g�c�z���1\��S�PT|Χ��r��SqŁ�A��D'z�,�u_*�MHۮ�������K����Y]wml�����蟽�RR�[�
]*��r�}/�b�V�M�kW��^�]��`�TO6�oZ��ш��E(B�Oo�@�1$ouA7 ����{;�o���P��N[�p�L;�'^�!m@f�Ϛ
�w�5[�P�ق�&���j�9^���]�c�Z\�_*j,���}�j�٘5���r���\�,�s�AWzSQ��"B�9�;���/�t4��m�P)�ܗ�5롹5�:ƕ5��%���N&�$�:�y�I�)u��Xg�bL�N�x����طx/B�����$����M]z�xgC�7ɂ����D����G�u��M��e�#��k�Aϼ���������<���g��|:��(���ڭ쫈pϛ���_w+�O��|��)���q���X�8rU^B/�#�䒣s�p��F�.���]>��D�y��2N��+}.17�����ܾ��V�;�.Th���)��,�D���T�L~M��1R���0��ЅWTX��ᓃ��`��;����b(����R���c�BQq���Ǎ�A���'��9t�ln���S�]Գ�K��+"�u6���eT4Ev����xxwO�*���gX6�%ƹ�]�������j���9/�@�{*�<cI��zb}�5	��RǺ�v��|��F�/�}
��j�6�EA��� �Z[C�d�b�6Q�tn�/�S�>�7,E0b<�W5`�:h��g�J3;z�'�{���W��;�<�z�;-��
	�M�]nou�l^�I�q�����uP�-o{=B�U��f�]B!�=��b%��6ɩe��Q���������h�K�.5$q,�N9�/^�΋ا�y��B֬#4�^���&;�V0��e4Y���q�G�}cB8�b��L��I�g�(m���ɍ��	��������㣵��Yp��{C��|�lØ�mǁMW"�	p
�H��>���V6�ۄ�!^'@����]<;�3��m�M��|Р���U�RΞ�{��Kc���G���[Q�\��g5���'mu�|��ͫKA�%��<ߥ�W>Q�09��DA���=�K�ד˾���y
܈���$Dǎ��ۣ3&���5��nMۥh�ˎ�V;��W���}�A5�p��}�h35¶<�t��H�jf;��Y����u�m�쩽��%ʚ35��V����x��|(��-ժW�B���#jHe1����0:':,6=�t�����1'4;<.�:�c��������5&�e5��r�T6m�ډ6ц�E�?�_W�<��I-��G���J���ݳn�ͪ6u�=�S�S�k�lŒF껇���)���xR�T�v����n,���$�s��� o�=��_�*l��^���_�f4�{�%*��rNA�vn�!�{��z�.y�5��
�sdIǗ*��E�|b��������������v�\8J�bګʔw�f��e�����ֲ��Un�����a"��U&�c�e�i�K��[1���F4��1�Ɂ�u�Z�L�-a��Oؔ�����܌S�I�{j�
��g�C��xx
�!#G�-P����r8��N�\�[	���/_�
Ȩz��/V2����ܕ�� �����iR��"/Tue�jDm�zY	ˁz����oc�S>��e��~9�ӟW��7?s��+�J))�V��X:S+���~�*��;;ܚ&� 䖞�fAV&O�z�ӑ���Z��,ݮ�"E�>+X�������i\X;�oL��EI��gv�k��tu�X2�9r��<�Ԏ�f!o�����Y�C9�����9aSz$�S����ƌ�W�Uõ��=���J�f�;����m�h��|_X[��O��K)\��q�7�tY�ZWI!*���9[yO�J0���o��z�Y)Q�-���X@nXۋ�*,��=���V�F�MA*C�^����᲻rV�����=�{����?=�t0f�<��3��QM�)���V7 JLd�Z/�U75��5�(�'d�WG�YS�g�5߳f�|�J Od!ˈ��ۗ4x���E���a�Ƶ93͒���M�T��z�4�G-���O�%�="��d�W)��@���A-x���v��u�� v�WN�"!�Y*�=v�f�)��L��3AuIIꂱv���ٚ�9
�� ����m�7�T�Y����@�(1ټ�'��j�Dp9Zċ�|A��E5#f�[3F&�q���ÜǄz��^��Z�4��?J������	5M^�S(^w���x��ޤD���W�%�M=���<Z��
�7��^q�Wo��z3ʄ����4v�Q���%��9�|ߨU�xdU<�P�}�nov��os��Kť�ŭQG풪�:��������s�O�b�e׊���[����ê&/6[��B��ſ��(S�in�	]�J�Z�%sJ���i���P�,���b�mLc58EA�/�H�Սx���n�7E�kވ⥬20�w�����B���G��fb���~������i��i3�#D��e�>��%ۧ�vo�3��]�6��;����J��3b��E٬�z�7��n��V9e�\�vK�5-�CÐ��G}8�r�7.=�znD�n�&u�&qi5���o	W�Y�n�Dk���ί�� C�VgOm�V_�1-2/�K;��7 S���Sf�qf���^���R�:��	��ջ�6�a�u���8v(=2K�iWb�[��9�����~U�y��
�g�{-�c<�LV�[R�i�{ÖS���^^~�t����������D��Q#��ڣ�j�Z�t�>*`:��j�ǃV��J�!%�6��G*�xѯ�1�Q���J9�ld-�ʮ�8�9}�3s7��|�h[FۀM���B�Ѽ�Ʀn�6��.o_UI���/���Il��Z�muUSTN�t�/;ZU&�xd�*��`Q�aoHS�9�	GU�j��7+hsd�[ȍ�J��T�wss�mY��k�>T���ʡײ#+�鯻�
\o���*N8�r��q|������;"�{�)�)vk<�z�c���!�F4�����Ϛ�E��2!�
	��42�a���0�������[}./>�=ܷg��������9�@�|��_Gz�T5JXww�6z�<�w�11=a�	�'U�D�1*˫���VdB67s��4R�1�U���G�������$��lC���\u%�4r�t���y���h�sR��I_eՕ�1����WEݼE�v�"�GY�z���_iݡx�N��P�r\��H,�.���ö���K�Ff�d�c e�)q��&JKxJ�&��
s8: � oe�	�r���fT噊��/)�N�����Ym�8ܼ7��b���"jq��WfP���=��2�A�Mu�3�������N���V�4�g�҈:�8HKx^�ī5��|W;Nvݸ ��w�><9g��QF�6�>U(�Wo�PهI���8���"��AT�8iY�r���wT�M&���HYT�r��.���dW˄�)\�����-t�U��t˘�p�Sq�Z��i'�u��Mpk��#��X��6n���l�Ҩvk�vP�"=[��%[H< #��0�ν��j7,Z�x�gf������0)�wqVs���6֎։ƒt"�Zs�2�x�Y����U��ep*�b���ڱ��f���bk]�����'�;E]M�YYx�;�E�oT�r�˓��J�o�����Q�=Ol����"��t�VJ��!�i�����{R�y��6����F������+�j\O�#ܳ}��'5,ꇹf�#lU���$1_>Ts���1|]�J�V�e�[|����q!�zr� �X"�F�û3�y(�y;�C7�����%}�b��=Aޢ�h���]�8�N^�ؠ�TH�A�ŵ�NT��Oc�L�<�]�\W~���󭂦�NX؎�6�PJ��ÀTSҩZ��˽�q��|�^q9en2éti
[*�
�,+�)tEj��HGz��}��/�[,Ftnu�HŲ-u97k��*��|�Bl�yN���~���
+w-����^���@7	��sv��V����R���m���`��鑗�)Y&�M�Ҵa�7J��f}��S��׶E�Zo1w}�F��퐕��n�!<#���.�W�)�FZGc}��kĊj��o��"�����N��r�-i'�`�*e��؉�ñ������e��<�3�L�ˬR�<�Hl �%��c�=��d-�ך���A�w6�7�%��B\�P�7[/d�lj:�ܲO%�A����%LO!wR��rPu�geJ�&����%:��1K��5c�W�.�#�M�٤f�;O��y�X+y�+��r�T0��>W5�U�i>e6�ioS�|p��jN���Sp���
Xy�1ֱ�k&|4�H٨��U���c��kot4K;R���"=]-20�Vh#$�q��7[�*5���۵��ܖ������
�x� L�T�����v����"�\bu�fYk��r��.ڻ��ggoj�}4m^L�q��@�~Z�lQ�B6Hlr��t�nR���-ې���89����}�G�~�.�DQ��Y,�-CA)5�&�ʥ�AV~3��;�Q�9��|C��q�Ε9b���˥q)2Ԩ�IRM��A�ReYHj�U���S��}�|>{�󻖉QQXdA9K��*T�uq�8N�%KE�"|�~>E8T�F���s��{ǽǘAމ���REʢ�!,���U�����s)����2�Y7��{�č��T\��t�Ir�l�PJ�4HT��igg�;�
�2���8QM�sUL������K���'ȺV�RK��?�-3(��)6_�n���ΎEs닷8�%Uj� Tu��_x��4���܍D�=n�#�˜�TY��{�g#��\��"+|�����DU<K��G>xy�[QnNy=�p���9%UUg|�B� ��[��ǅ_!�(_�O�wT�W,�hDQr��8�Ȃ!
��"� ���^�K)�����Ra���ilOU�w��L6��u�t
lяx�y'(�>��c�T�߾����ǻ��T�?��Ӿ�y�N�����u5�U���}���'��9d���ו�N�Ј{{��j�vz�:4��DOݑ�:�+/B1�9R.�$S,��SϪ����xX2e��-C�g���Xz{�ܔ纭_��Ə����~�5���(4�$%����^���+��}Rz~P�M�7�s�ӛ{��B��C�S\�5-or(��f�Ͽ-����P_��`L�?\-zkK�����ذ����q��z���}�>xS���(���j�}B�cj�;[	b�U�W�����r�GVvp���ǐ�����=��0�݅Yf`���W���]��ĵD���Ma���YNUn��� ��z��ZBTn��3����F�z���J|�5gCUo_�t8��a�sw�����o/�{jH���}�b"�T�R����[�N����?qam1�s!g�4Ӯ�RYn�@�"R��91�H�q��Ju>^�Q�V!�{�j�K��&0��ճ��,r	ual�Bu���L�50����ql��'ҹ���.x�k��W�FAC6���Lu�`��c6��|ޙ�/R"G�d���<��*�yW��`]*�]�u�Z����Vn;���<4M�J*��i:���t@a�u���v򶄲7qu���ؖY��ã��a�wxC��I��v����.���4�d����7�v��u8�	�=�uڗ5��@��r 鄉�ŕu��Fn�x�N�A��W�wu�$XY<����ϴ�<���f�c�<v:������zD.S�ڇ>]��vzMf��۲Km� ڀ��� ׵L�ǝn�6���^������ra��El� @�*._���Oa�ߥ���6���G
�'�w[�:����$�BV��D��J�M9�������@1t��}H�褝�|q�R�G�M�O^��qM��BB<n&�$L��5�
Uv�I����*����A���)����>9��@���p�f�ee*��]�t�wW�~ޛ`���г1��QMg�n�~>ۗXE.T-��м}\0F�����������w�~u���	M,��eN��tĖ�%�.{O%�b��*�q|;e�moZ���,�x��n�f�������?@��6`�(X��&|����Q��$�~J|��V/^g2/�kNf=;U9>�q��,f���v�!FU܉�U���r8} �����-�~��#d�C����]���]G�H��>
�����ZOs!u�.�O!�,֦$�x4���k8�aゞ��>��';E4�DROރ�<n�_<;30
MˏbS��K�8�%��.@U��Wʳ6�d��S6cn��$T:��L�)}0�Ohr��O��U�{�$�(��&����f�����J��/��똽�����%e^��������T�'^��b*L�4�͎���Ͷ��Ԗ%��&[�l��p�sRREZ�ghJ�vgy�su˂g�L訦6�^�(��������YFKs���Z�]�<9���G!t��κ�|Z�^Wv��P��L�'�r=��D�­S����������!Xř�ă�[{�y���:����c>0A,/C�Bf3S�%���-��'U�H�[���R����h�,.6���~�<Nm��`üE��T4�r�<��a"�_U�2cC�Ֆ�9��L�[� j�n!5By��1��W4[����P�z� ��"�	􈌋�r�XF\����t���x�pu�ުY�]����H�+��-̳˪JN�IX��G� �H�����k7��Ӣ|����ћpj�;U���-_���b�|A}SV6abu''�q�T�쥙����j�Ss	�����m��G��ci����V��Ы�:Ă}R���L���#��I��{I��:�kSS�E��
�ͬ�٣wd6üZ��_�[$�X��)��r :�a-r `1Eٛ�;��K�mݻ��7*PQN����g��rv�}si����[� � ��B5Mr�q�ݱʮ�,F����Ee���蝹!S3l�qo��6K��ЪKT�-3�Ul�F��1ߜ7��B�c�z�wQZ�]����U��Ϛ�ڤ��^>2����7
��i��Ҽl*��ji��dN9��5ն��nT���V�j��wB���<�PŖ����Ҁh��<ҿ@�r|�����`�)����eoE����W��d\�Sm�2q�O]2�\P}�i��l�0.z�9b���Vn�Ռ��]�K��sXK�sQ���9Գ�a����:�]ơ.B� ��l�8V_���V;�ű�s��U@ƌ�y><i�sW�qMi�{v��ŧ�:�ȩ�l�=;ת-�M�>�=|׎�L}o�b"1Q�GS��ĝ�s�����Z�Gr}n$n*x�Y�Uۛ2�W��7���)��B~.���H'�o�L����q��cu&���qA�Ӷ�_�J5�kʦU;��nu��G��O�vB��yT���J��FNmx��:��%���eQ[�׽:�v��<�O��Ua����A��"�	��:��!����~��@�Z��S\��4�����?�l�=?I���]�7��gG�{�=|����t��8�P���]���Y�Z���f�bX�ٕ��N�fC����uP��dt��v&ώ��}�6B�㩍{�D&>ܱӽ�u��pb$�-�'{����m��<V��&zk�邖���' �,�	��]P:���=�e�w�7ӯ��,_���1�.���H��^�t������ޔM�1�>���\�n3���nK��5Ӧ�Ѷ���vM��{�5��bE�Ϛ
�uRiM���P�.�T�:�;�i%e<PdN�g�B���l��wv�4�f� �!�{��97�[��{&n�_G�:�"��a9��v@q��,+l�vO��oSGQ�nk��9-E�"&Iu2��F�e��zܓ���խۄF�Q5R^�P�� 9R.�&�,��Sȭ���R�֢{*�T8{�k�qϓ���x�E�����k��u�E�e��mvܦۘ6��Y�ڦ�R`ʼln�U��X�,i�@tě{�'%�QI��M��-{��s����"�|ؑ�u�j�Ws4�Z%�Nѷl���zVK��n���9���T�Ŏ�+^ҋNN��k}z�޹�Z�zґJ��X�9[5��2��`��'���j<��Le�AF~�n��9���	�>�@�o ޲����4������T$��r+�)��l�CqM�ژ,`y���׸s��[tU����D���gPҳ�[�X�<v�ýJueϞ�173�唶�ߚ�Ut7��D����pJC�YX��E�i�֭E{�a�E�d���[��˰$ �^nu�o~������7W؆�?em�7�/��86%C�BW R���/U#z��}��|�v�������O�H�k�����-��w_������0��쎩Q��J���+ _E���w��o�΍����*Hr]nSI{H�d��3>�-�|����q,��\8�PcS�Nɐ���m'o.	b��8�]�����c�S�Y��r��8J�?��~��F�ihj�f]�.+j�]�w)��R�5Ec�~��BI�N0��m�:Dl�u�ú�=���+���Y�>>��cx�Č��<hH[�k�}��ް�$ܖ�/n��y�Ѓ6�"�Lͬ	��{��y�mx5I�ԥ{_(rV/j�Y�$������tb[^/]��
t�=Xr�7s\�s�i���c@�9�t�RW+�P��$RW�E	sf�럆�Y��$;�(�z:���Zw���q=��$`�k�"1�AWN�>Fm�P���ɢ��{��fa��/��(�uln^�CBxU6���8��ë0�(z��`θoy%o��Aۨ�]~��l�K�EK�|	}�
����#��^ܭQ�����P����^��ļ�����t�Z��o�ZvAXe��Q��76h�y� u�^�b��� �1u�GN,ٕ����:�R��_WCm�8�$���G�ƞ3BY{U���(�1��'V^�C^s�?�}T�������ƻ?ї��8��ʛaAj��xa�W�qMg�wB����O.T)څ��U4�]8մnjZd�D�����g6�epL���Usw6bY�ﻡ���"��w"�J���ӑ�.
�3{�'�C�y@�����f�e�����ƣ��f1�=׆�7��ǩ
�xq�b1w{�~6���X��$$ʻ�?G9V��e��C@�2��(��x0ƕ�&g�\�j��Oǟ�%>��X��b]`��3����ƽC������B�M��g��]��:Gk�P*�1I��^�s�9u��Ɣ����@(�;BT3���b\Y��t�1�ۯi�Y�#���V�9"��їZ�arQ��o�9�84U�W"�!d�.��c�z6��jA�^�}��*b5�W�`�V*=�;8زT�q��z�:��q|�.(j/�b�s�^��4v߼.=z��m����#�ho����1I̼�잢ŃWP�Jz.��[$�i��a��W�kVWb�E��<SU����@8��!H9�����sL���U�F濃`d��M��soҲh=���]��{&x���Ͼ�;.w�O9Q�;�~�3�%�˵-���h&�]�KU�d�R�^�nb$c�.j��+��}��rn���9�)j�(0I�o�e&Ւ#���vG3��7�s K�O�o�KZ���;j̗�k>a�u�L�N5�.��t[�?�{�{���Wv�ߩ���Z5���)��hJ=@ls�''�"2/��(��M�	�����i��@���Z�uCZ/vdf��
ʑ�!�S4꒓��+TG��DL��B%�����������I��'�"s2zwG4�y�0r��"Ďs�����X�DI�]�Wx��7�ۈ�^��̤�/C՘�s�cy��N�`�e���0]}�H���� ������Q���k�O�s5Y���us��\w�Jk=3Go9�7�C1N����{����<:�K����!piY�������_BEy��}s_qѰ��x�,��O{���v������7V��Jp����
��)B��icU
�JT]���9^ ����̮7����vw��]7��� ��e�L���������g��M9�~��;j����k�����L����b-��r`�++ÎЪ�l��yNXP*�7vy*�ڵ'_�Ż�aqm2b<f��/
A�~�6.�wl�G����d�x�C��(���q|�A�/��Ӝ㼰�~��3%�Rb���D+��b�ڴ��v���s1��ͪ�R}4���7?lʆ wȺ�eZeg��C�g�V��__�=Ay=�
:��j��ZU��m��[��^�����c+]�c�u���]wO-��T�Q���:{%�Ͼ��Aa�rx����������zz]c�,��pޮ%�D�U����D�׺�\��Mܜ����;­6�% �S�:�F�""��2rFM�q�}ԚhZq]��p�����~���xD��gU�����_�<�hg�v��� kvo/}*q3_J��FNmx�B���ʩML�u[{�s����qT߫�k�g��r�P� ��zB�r*���]�T��uUc���K�f�=��3r1�`���Ϻ��W��k��|���>� O��
�K§S,�qL]���X��� /H���]��j�Ōcμ�5;�U�cEOA�P(��b�r�u9k�ˉ�Q������Q�3�,��P��7 ��{��2�o%e7�@�a�V�]z�ɻ�U^��ۯvv�5k�%E����-I�������y��i�ڨn�2��ۖ�v�$[��S�:�לH��~2��Rj�RX��u�ϐ)�E�'�&��u� V0��׏U�q�A2�k,2g1����޴�𼌖8���F�1�"'��#U%�U
�Jl���E���s՚^�}2��1m��]�`\w�`T�$
N��i,8�nEv���}��7o��4��zg��e�W�y,��֧�Ot��[A;�p�cE+��>J�Z����#)7g$V�XΖ7&Df�-Q�
�k���´&A�k�uӍ\8��)��h���Y��-=o-h�p`��j�{��{���1�1��I���W���� ɫ�$����wg�ɴ�����$ٻ5�g3]٩׈�W�EM�5yێ�#�Hx������^�SO���>i�@��۫j�r�\*N��:Y�]샶��=�p�b���dn���H����<�]v,n<�s"�@�^"�z����Z�5�U�,���0�.�e�|aq��� �k(z4��:G����,�����wgE��hX�
��=���s��h+r��P;��:Ĩ{P@���<��9�R�;��Z�t6*#f{K��3]Z�'���l,>�}~����jJ
�0�Odu	Q��J���3�+T#^���X��<�^����4��-��#%��'�hD���I����P��V�����5=EҦ�Ր�]
z瞒�]��I���憩�O����W�l��B8�~��o�g-����ɋ��u7���Jia�%n+�T^@�61�N2�]Cʄu	5\��x�Ux�Zy�U�I��˕���><&`�Č��K4$.��7'���V	u����6��)L7}����=޿/;u����Ow�	�󋦱�;C�
cy̽�7�w�6�،lx��mk�ׇ5�D���e.%]W�e��q��2�I�u���I��@��?)[�ڵ��u��@v�m����T����b��2ܦ9>N���Ȋ�֚1̠��d��Rʇk._׷Ke=���ս���9R��Ȕs�����\����x���G+�c{$U27���دõf,� {S�2��C�!�9��"{ǫr�P�2�boYV��]��<�eek�د�k�Yu��g�S�X�X}צ���&z�qR޶x�z���Q��(�!����@
��no* ��HȋߧPK�u���� R'L}u��\��Tf�Fvd/A���q,�k����h�ڽ=��o)�a�H��Ցɉm�|��GzgN7r`Y՝�I#i�0a��q4ED��<�D�m�r"� �S]@G�Ño���uԺL�Mo	s����1�q�=s��t�Δ�[�Z��؃���z�zv�}'p��Gh���(�uj�K��C��� �Ӗ���3�Wr����|FN݉AF#6�S�7�z{uȦ�[��#*��[.oIX��
�n�9ݥ�@'dL�4Ԡa`*Z8��*>蛛M�����o�74jU�t4���J6�X{vq�_U��F����X�4�NU��8�]>��:6M�WR�2�U�Uw�V�#�m[��e타I�[W��\�0�6`C]���P�&�˪�F�6f��`Q����_U�F�kYպ�)�V*2�-��t���u5WAS�����v���\d�h*:�;=�*km��[�C�f��ձҿ����qW>�VOIf��|vU����X�!��9�X��JQ2���yJ��Mq�����X7��	}��P0mwHȆ&:.;
�����E=�r�b������o\�mo�Z��yq���b:]�&��;�f;��4[:c".QIl�J_P��N �rZ��e����/6���Wc{:hW�6M#��eֺȨ�U���i�8�X;ls��x�%�'I��;���*)�ԅ���0"w>�.gv��N۾1�u̟E������5�����f���\v�0�m7�n,5[/%+� ��x�vއYʑC�ԈD`z�t&E�:��]�fZա�u�Ce=��V]�n���KO��+�\��G�7 #3���L��{H�E	v:���)�g�;˄
��0�7hL��^Q�"j�gq��}2:T��q7�2�6-��ܴ��`˭����GQ���So����j�n��꽴�|0�I�Ke*���q1�+�1V��n:,��|wjb�w6s��+"W������[��]!�l�3�aӼ�l�YL��fc����̊d-eL���j��}ia��c��sv*nb&Q�ʁ-��C\�<5b�U��T��6�u�g[?HN7r��O�/�m�+�B�j�����4�z���w��9Y���Md�������;%����K�HG3��d�A��ۉ��.��,��:ĝ���y!��[z��A\�}��xP�W��w�5�*�k�W8�JjЉR�o{�>�%@�6ԋL��RR�'eQ��Tɚ}�<U�G"�UO$����
9yiJMK$*��.����s�/�gymO��XG�u��Zs5D���*�	o�/y�%GC眷�]���V��8Z�E�5�*����e�!�����k�{����U������h��hz��g����"�'3��r/9aȐ��u���$�W�qpB"�\�9f�ʜ��׺L�s�@�#Qh��]8��\��u9\Ԋ?)Rg�DZ���s#D�2؁Y�r
2BTM�r֔V�.g�p�,�-iDETEt��MY��z���Β �I$T��\ⴥ�PDUz���THC!{�U.��D��1��*��'p��������u:��ٖ�޻ɔ��ll��޽�ۜ*	2�f�]�x��1����?��SB��TUQ�}��BY�Ԍ�����?�
�P�)gPP#�#"2=��b�{����G���;�����Όl�ЧDX�CKΧ�|N�+�s��C!��itQMV�K8����F�:׾��m	�MNu��p5c+�u��E���
������~�T��|���>8�~�8�/t�P��i��F��CE�;h���սP�{�C��UB�L�#�p/\O�O��q$�)(>�k�D}�/��7v\|�{S��̓�?6^��4
���5BǠ,���LQ}�r'hr�*	^��
;3�����\�f�y���G��c���o��ĥU��Mz�Xu�6�	�{[��b���c6D�M*A�zc=�u޽�|����?G��3f��-�5��W�[<#d�k
S(Ov���ۢ�Ӝ����7W��y+�Wٔ6����}ǆ��T>=�\�]Y ���d�*�1�F�(��=�9��|�]˟������E>��T��o��~E+(��A�s1pzse�+t�����,m�N��R��{��L3�x/���+������L�dz�Y����|�AH�~���w���X����I12o� a�H(�V�L�+2����"<����u(lS02ʕ���Mb��48x�<[x�\�A�ze+㽃�M��[mp*�)o2j�+�Z�@�x䠞/|7k;բ�.����h5kt�f�����,�����	ֶ�R^ʆ�1v�$���a�5��F9�x������U�,�%��9�����Z|_]���ˤ����l��3�ycK��i���^��.e����6.�*����ިO@,��`%:\U��L�UȒT+��ݔ<զ �ND�!� ��f����*)��t��uX�	I�����6���'�s��Ǿ�\�?pX����0��
�zB�r����#����=[N���� ���^�|���c|s1ՠ�kE�y�Xu�?|������.�Q@ȉ#�OX�^	K`T�k�������~����<M��f�]RRu�%b�`����xڳ+�n��cZ��vp���%��̕^�ir��:X;�ÜQC��Ml%��kW����q��(����+�Ql'��T��Q��S͇ &����e�%(7X-R���x෵�_��D�K�S'�&�t����h��S��>X�f|�p����u�2���(O4U�	��:~��Xv��<�4�©�Ɓ?�mĽ
zwƗ{kiZ�Ƅ!�W���?q��> o�2�78K��FU�/Ֆ�ΗKz.ksx��[�\�%wegL50���k�Nҧ�k������vD��p���k�\[���n�&�/=
�q�*l�͢��GGF��.p(Y��V%tc��P�q����5U�9�t�s>u��I���S�t=�#��l{���1�3m��V��n���c�Ձ+�)Qv�J�U�C�^�[� Ʃ�ex��\Ovj�OMb,��S���굕�+�Fd@�^C��}�g7ً5-]�q ��.�Y������ǳv��Ƒ{bS�UJn�	+���Γ�}1㰤r��*s�Ϯjb:�<.��B:zX�;B�q�Ήz��u:�G���C�Ӽ���W�ѕ5^Pf{y����AFЯpG�DDb��-Ϯ%���T7�����W'��	}P�!��h���ۀɵ0z����_5W���Q]�uJ�"b!���Qʷ<h����G�2`�c]���"��N�����BJ�����Gk��*n�Rq��J�Lԩ8k٨�o��v=��D�/��t�핬�����t������S�j��FJ=]=?D0�1>[S����X��5G�OXG�5�Q�ڗb�;�_z��g�-��}�4	�ʮ�4��@ln'�6׵9ѓJ��t�R�C��
�_r�b��t���/U�l�%��0L9��)���Y�"���7p��Ճ/�.�h#GN���qа�q�WՒc֎���t��^@�����=ܐ]WFl�1�W��]�)�\ٱ����7��!�+5��7���˶^�d����d��b���žT��(���t����u����շ�&ɭq�'��Gy�����|=��~v�gf���sCL���%���G;ݴ��]�(3���#G��Vlo�'��L����;�v>�K�V�V�N��(���������͓��s[�>�������q�^��~�䗘��m��E��f���Қ���(hG;c�l��^���[�6��qS��*QSۼg��uJ��s�%�^�W4٫%�;T�4j��ʾ�v�.r=B.Ex�(����)����{zg����g����:���q'����n��`���A��y�Q�U����v2!ћ�;T�vmĸ2��[�u{ kG��k���8伧\�ڢ��[�;�j�s�;)��fi"$��=N�h�h��/��)/�(���Xp~R��s*��%��R+H��{1H�� `������a����Ё�>ɠ�0�Y1�}ȵ�Q����Ҏ�s�~]��f��9�G]��X�7�N�֠�ʇ���.�A�o�(�C��P�A�teYC�{|Y�j*��$F�̌�~F�7wZ�E\��ǹtX�l��\����JXFLl��B�A5���i�,�G?ۘq���C���� �\3�j7{�e�t»zr=S8�s����Ti'���eX����(��(��UF`��XPT���f�k!:�H^`�IJ�53ts����u8ym້�#.���;�Y��	��c>�ޥ�Oس��am9����S���Ypo�-��_GK� ��iNQ�n�(�>b%+��m�`4�i��c��Y��̧���<Rk�A��AA�գc�Od�L6��4'Y��֓5�^��}#�8�����-�5j`l��p�]�����Ҥ�X~�q�yS[�5}�X���H�װGL�k��2yU�;S�9s8�����v
��"�H��F�Xd�zC�s[�^�c��%���}�~G�܂ϛWnro���]�5�%r�R�u|�Q�pX���<�������ɯMD������Y�5F�CI'MT��ı���.�'��~�H��)��)gP
�7�#���SS�7=�X[R�ίD�fNm��{��s�P^-a	�kX^&��H��I;��㉅8����䶫Ӷ�ZW������F�&N���G�5
��u���L�ۆV�n�9����� 7���oka�4A)��}=U�������P�	�ǗR���<U�~/)���o�k
h��$�Pf��u���r��P��1f���WD�T:9�?U����|{�=��y֟��o�W1���hCt��0�)S���nFv�j�v�ej�������J�V��kb�0�Ҧ��J��x�N5e���S):�mZ���ďY�G����8����}L�ۊs�W�wW�݃��J�(r���ś����vՙ��Jz�V�9;q�����w>�2�]W(M|պ��i�H��c��m��m8���q�24ڝbՓ�n�΃�2��E��5�2���ϊ8��X�-fP�rr�Ķ�̑0T�U��m����f�x)��E�=Ҟͭ���	>��^Ne��^���ퟩ��g�T��o��~TE��z�}qnfz�}���y�����y��*�Y�uK;���e����+��A�Ғ��/���F�0��<��m�2Ĩӕ09�z�y�v2oH��4e����X(�f�|�t���a�E71�J6ν���E0��CXz��GC;�lm�x{��:C͝j��uY[�غ;G�:����v���5���d�\H=ؠ`����F�Й�NlTS)��[�N�&GC[�Ib�M�q�.����F���Ĕ�E���GM��5C�+�@�P� �& >��\�$��n#����}��2�����N�'dŗz1��O4c��,\З=���B8�'�*H�YW�\��U����2V�w�y��)!�x#��_Q;�v�9@�܇��ߩ��uII�ۓF$Ll��ƯK	���������B+�V|A��p�^b�9	w��:+��B��wk�4��¯(�x޻R���v�x����X�e�7w_>�b�r\n��Z��$�*WP�p�{v�Q�>TS�Cr�Vu_M��,����|���/_a;9��ԞqSY(�n��'�̞�]��.M&��$X�s���Ү������F9ݼ=�,B"[~ab�SQg#uF�$����0˅_7�bD�N��S�'��*���w��Ԃs�"'뺘1�sEjiY�Ԡ�3�=U���_1,¤��n�{�s3s6��Z#�ĺ�Q{��(����RVg�|d-s�B�^����}����v{&]�eUtu�\^���wt�e�T�s`b�e�1V7����-�xy���\E¢K�`�J���]}����w�7]\�	~�˦$�&!1ҦX�����YXQ��*�TW�cY��k��OuB|�K|�w^~pVڃ����3D?A�BD��]�ܶՙ���E���M?�9~�>�P��ٺ/�2�1d9�(�������!OoS�<S�jӊkO�Ɲt��7����U�A���o{/���2��b:`+�I5�5Y�fM�nl�#p��8�����1(ih�����3�s��[�@�Wʊ�cW$�!���:D��$DC9�2rr�q�X1����;ܽ��t��4t֌�\d�b�5��U����;LI�e8����Z���<.�z��-P�{˃���X�{)��/o[���c��TK/�D��v���|�ҦX����al@\�����	1�k��]tt�X<��w_�:[��3�����PcR�<��.8ͱ�G(l{�(�!H.7�J�L��.�]S7c�cwє!Eu�ϫ[�W�����g�.���C�&gZ�#%��0����h���f6;c}uWJӊ���7fsoH��NQ��U�jG��j���O�O�����3^�MIK�hG]u��yǹ<Q�=z;�+����
�c��Ks���0�b_|��|WPA�R{yiIꦣ99[Wq�z/��
#�Ȅ}��n>.8��=s��q�����f����x5����n��5-���J�J���C�v���� 6�h��2��{�����S?K�m�첤����jG��ڊɮF��t�,�{����kL��	�!\
2#����x�TYdɄ�gf��=���=ح�$vk��9-Cpɵ��h߆<�C�J#�j��ʡ]���U���T��Җe��;yІ�@T��>�n�X89��PPdőf�7uG��٧�iA�����i���e3��9CZ�crYX�͕쀚���LIǿ���)9�R)��S������#;��7�jd�Z���x�B��Aɉ�/Nl���Z���MoR˼�HY��ҝ���;���N�M5��d,���¹]{�����d�	��m+j�Jf���[zS�qyku����p��rM�,����.�dȯ��P�Ƈ�ȭ77�_�3n��"��t���\�p}��޺�?fW��/���lR^4%�Gk#�)�<����paF���;�Pi;p�­���R�vr�*��8�={�>���Ș�g�G(Md�4�������m�cdvEYYU�v�p��+L!������<��H��-�5�}-�3�W��L����?lT�����M�����-醐��R.�<x�E�����c.5%�a���n��D�T��.�5��1�D�^.��W�
�<�7(ж�0eh�a��^Η�:'�0�+�ܔ��D޾�ǭA;���;!����J�[�ԫ�GO*d¤�p(�t���E��j����+"�6��*�`Ԭ�m�l3��E �҇.,ܡ��J⚭�������֚"�:�M�q1�b�FV<wYoi;�6
k� Q�PTlH�����xvϴ��`� �f�b��Jp�u�����ަ����տ���Y��r!r���K:������^<�ݴͶ�,�����CM7vc�,�^G�u,⽩f�&��ۺF��I�9ءg�D;�3bGP*�����	G�@�T)�t3Z��l���eH�I֮]�e`춈}���ݼ{t:-�Y�7�<�P�`*��N�/`m-��;Ux�^Vl�^������Fd創��QP�2�VE����NKi��W/\�*�jz������J����6/X��s�`=��c8��3��E�O����Ǒ?����ً`SQQ]{p��P��s�FN�9CV3B4�|��Oֶ⚙��EF����ݗ�^ȵG+�n��Wj[XPO"���I��=��X]}���Tȍ�[�u�E1�q�>�u�`��_9��I�g7�E�n�OF��<h���Dv�֐rs��Z7E[b��q��&6C�/���ch����wN�����}��+�;Uv#v�/Զd9M�-Y�{y�By�}'&��݉�i=>c��|����G6�f������)�,R�&z������ev~g�F�R.��o��ii�.����#n�s�� �ՉŪ�c�⊫Y��+�W�a�O�5���Uvzx\�T
�)�vlj38����ѷBڻ���-��w(�z ��TJQ�k�<�G����}�Y���Dz�R��Xƻtv�xe��8���̆�|L�@�`zH����;�VK��D�Fp ݍy�mi�y��!7�\��(�.�n��p��[SF����}�u��kk�`b�ug J51%�z����_�i������$L�� #k��&��b]3�th%�ʻ3��au��Cs�쉿gaDb���k���@�A<j���4�e�s���&ih�y�r�d��As��t0e�)�Q�Ou�Z"괥��-�e�Z^]����ĝ��m5P���H�ܮP(�`v�|�c#t�72]�z�]WS79����j<�(���YY���s��]:��a���b����^mn�B*���䰝a��mGY��.�|Yvʕ��1�Ͱ��ۥc���$"�|�Jqv,�;t����C"��#e^���0i �j-J��r���7�rɗR��{���B�d-�ƻ���[G�&�w�K8�hr�z^�d�*B��	���38�"S��e��X�ڠ��fS�1����In����4���vo��*���u����4�.���͝�f�µpoL��)Ϻ�"��m"ˇ^n��Hji   [X�]�.[��%+�2:ε]?3����T�NYc�J�n[7K5�J3P�u0m�f�n�oY��)�AC�K��WR�*ud����B���Q���u�A%���!"&j[*���u�Vޒ��%��^����pq��#q��9�6RI���)���\Y&�6rH�T��Æ�c�O;����j�Mm��)��8�[7&`��t�"���%Ӕ2�1�n�`�`�5�5.����J���X���r$]XEe�����MR�����īʘF���B��AÉҩh�.���J�_0��K�[*]^�Qܜ��W*f��&�w?���Se.b�L�Kz��
=�v0
���w,�Pg�On�ұ�l����Њwk<�0d��n����+�� ��Ǆ$���O�����>G�|�}׸s�צS����[ƛ~oޯ{�ŷ%�e�p{���<r�,�n��܊��,p��SM!����Sם����W�j���"�ݍ�yu�0+����z�^���*��g�8*@������C;#zI|�Y�U�ǭ�]&�N ��fh�ŴK'�Yz�s5�A���L�-^�y�����+N>�f�d��;I�)a��}԰���)M2�姟o�Rp6侤���XCX�
V�]N��f+i�ѓKU�'�^��NԹ?���R�>у.�(ie�Ebp=��S�U<(+h�V�q�\�m˸��}->�%1��-��m�+s;$hYy��1�H�Y�@� ��%�B�j�v�k�7�pS55U��o�<e�R��i[��A�ec:1K�L8����T�;�``� sR�a��vu��f]y,e*�6��Ϋ]Az.��X�`pĳ�t��Һ���g)c�A7v���^�Djf�[�X�Jeά��t6e�LQ>�������ۋ?���Q!����ާJ����G**|HQTr�T�dJ�"�I��Jar�"�2�7R���Բ$Ⱥ�%%�*9���a�Y�g��T!4J�A!��D�"%�QÑG�I�9APA*d�"ugs*�2,5"9j�Ȫ"�%�TUETPE�DGWt')B�FF���Ԩ�H9]2��QS�=�=���p�dG΅gD6TEVa/�<ʓ�d�FIDDW(��7�%\�DM̪,�C�hE^+,�C$�\":dp����(�\��=ۜ��L�5}����r�><���/S�s�sG<"#_;H�PUr���T"z%�ri]�(��=Р����E��F=ز"��P�m*s/��p#�We2�|�����K)���*g?)*~�"�$�ٹw��:�����p⵰������:��N�0��K������%�N� ���v�p�,����5�]'�s�2?u�p�����t�n>�k�X-�}G�2�ۓ���`_Ԥ���y��瓭,��?yA���s����z��1��{aq�|L0\�5���nY鼑�و���	����s��5�~�a�ز�w�*�Wp��f#��⑇F�{OA�=���X�#V����lsMؖǺ��L�m=�Ȧ�xyH���ۣk�Si%1����,@�I���1�î�k:ɼ��|=sMdt1��!���*}f�����O\Q�)r�s��6��F�wKoe�	�M�@�R:[�<d*��f���S��'���l!t��DO�M��o��]��&��j2F�iGm�M�wnU/}Mt��S\`�c��=;3ػ]���/'X��%*�'jͭ�VeW��=[-ƻK�����4z�XW����ܤjhp5��ܮ0���j�9��ڥ1�ϔ�|�ʯ�2�-��� �x�3@2��� f�%hҺ	m�<�P�?,�a���X Cc;�6�A;k:8�+���/z�(����o���p{��@�nR�b�_Sk��Q���Z�]`X��V�W;q���IW�*h�'<�ڝm�{nK�6�!�g�3�U�ށ���;���-p�a.X�Wi��Xv���y����)>[E!;�n/0�V��L���c�پQ����e�q�1�����{/b�5(�љ{ݳ�||N��Ms��8� 2��z}p`u�3�L<��ptjg��/��蹪��˃�f�q��l��*ߧǙ�6p�Z]��Bޡ1�j�v���F��-�q��N�Βw���\�r�������g��3�������=�OK�ɒ[����d���V��I�;$�b}��!��x�j�9	�s*�{:e��l�7�.{_V�u� ��j��}�A�&C�#���)rXS�<f�����	>b5I� ٞ�����$s��4�p\�[:�2�[��:�����2c�q�����T�*�Ѧ 붤ׇG���{&2�]_n+�~����vs,�l6)x�|�$�&�P�5�~��n<�̫�q�]�McW;�Y��*C�O^��#�T.��&����q1mº{�3�k+��35;�J��Yu��%4�����d�A<�Kr�G*���æ�uṷ�I5[�-z.BH&�J�L��9�G����'P��F����]�i�ow��oE��,�wjĝ~�����=�#�5l��+-�|���_.��Ֆ��w�b�R���s�i~�v�{��3Ey�$2BU=�Z������d��C1�,���U��ڃ��izTrIٹ�C:U�Z����P)nݞ���ͭ���ξx���f��d7\6Rʎ��|sִ�Ι9`l%�c���cF�c��Ԙ:4x@�D�ONe�N��/j@e���$���6=}k���G�����)�G�w��8����k��e;�y�k�Ad_���]�ܳ��_�	1�o���PN�Һ2�r'��en�	wR7�iG���g�0�fӕaj�.�e���
�o3Zf؃��Gu�e�F�����X��(�v�n�8�Z]j{��G��Ѧ&X����ԃT���dƑeL��&h���]�,t(bM퓌M��3UA�G�*�t�wotu��T�DϢ
1ccMWr+V��{�?yvu��'%/�Z���i��ax�/�3��GMu��NrQ�Hٽ���p�d�[�%l��3t�\��!;�;W��!}���7����%�sl��BZV�_$�s���Û6^�����)��,ȷ#�d>h8;�nֹ�����ۜ޹�x��,�G���p�#N��H����":��\-쎜�{Pdχm=�Y���p����y%��TL֛�wO-r)������i�~�j��*@�����2O��2��`��Y�=34��ݽ��A����-#���l,����R̓2�vlJT����~�X{�춮�������!��"�J���Q��Ӝ��k�fØ�k��D�t�M��é��-r	ᓥNPՌ���\�)v��۵���n-�-�/�8�=�Yb��M�n�Y�u�Rp�}��ԽE�V���i�R��ɂd������,��;�>�˘�H�s�^؅n������f�������ڞ����j����dώ[)�dd5�6�0Se�Hc,U}v'2�B��wn'����0x&�G�{m*���c��9���3dMɻqӏM&^2)8�ݳ����[ԧ���䀲=ˬ��QhU���ƳC��m]i��l�R�o6l���SH$kw3�DC+&��[\�dvl�Q����9��p�9Fe#&Z�c��5c^����/�p�OD�L�|U�#mL�:��q�F�,�}.��^u�c�G���X+;���^c�d��*����ǸM�yb?���+�X�)՗U��wh�0:˴�J�M"�B[ϻs����A>j}fy/.Uy��wI�rj@g�ݰ�֞,=:�j��*��x����B��f�fݥ�[v�ق nޘ}�(Ԟ�;8�R��g��R|��=Sm�|/���X��q�[t��l+� �� ,}��C��q�^���피��m�/�.j�3�J��^�b;�>�e�;誉�y�l�=��s��4�ݭ4v����tė��2d7Hh_��Цƪ��/���_�ry�p���3�����Ŭ��{T��d2x�f�ukqY.^��Ƽ�Uw�\1׏X���V4oF��z䁐���(`ܳ�2x�E��!�q1�6ٮ������S�&�������\R�Fe�\	k�� ;��翋Ȥp���"�s�A��[6��r�<]){>c�ە�gS��ݩij�gt�1~+��L�v�j���:��ħ%ك_@�f
�;��Z�!O�Zg�薥BSwHMh١Yg:k̡³��R4�(�g�w���˟n�4wS)�l204�t]�V�F�T{؊������U��ō�~��x�+-�6Z�����ʥ﩯�D�pv��eM}�՝C�0g�^�]'`�(�Rv���(s��,��W�<�]�M���4e�)<wf+�^���z Wa���	m �zJ�["��J����
�k[шh�Xp�m��>j��kt�n�ǚC�]M�yX*�u�Xwl��Ʋ���{{׽�|:n�J�l�k�XE��.�GB�r30g=�bץ�ps�%/$y%}������]��p޷7��V��j�P�ەn�ݡ�����1�;f7d*ߨfpۢ-2!�Ϣ򝚒�{�+:+:�I�T7t��[���u�j�@�(��;Ұ#�x?�e�w����"�ɖ��I ٜ�i1�?l��w��܌�b{U��lg��b��0tս�=�J>?3��D�*����k����{�<���W�^�*��*v��A7@��n��Iv��]`�l�P��ݷ�bv�_Lu
�Ә�)��*m�ܦ1l�jO��*�}�yy#�ro!{�
�-��,͋��Gc�s��.������	�^n��j�fnQyOn5���7�ӍQY�'���_d�_oVU��޼��c�cp��G`�=��IZ��>&8r�R��7g!����ݠ@s[>l����2��B�0p��d��t��=�����w�f��W��K}ּ9>���7L�]%��6ʺڣ�|�{��79���.�t��#X>�_��חd���9!�2F��u[4#L�vS��d��7t*��&�h-��Eݖws˘�n�N*Ҥ�A?$�%1W�J�g�t���^g<��D(���C&[ae�+�NM΅�/�*�jN�J�(�L����6e�;;rﯺm��v/S�Ė�R�u�Vq߫���{������O��%cx2(�s�}m�ݹ�S�Veq���Q���k�)��
ե�"�"�fETA���y��xot�/G�������1���|N����+COމ̈́�;Faύ,5�ᐮ��eĬ�q���H���P�x��NV��x��^\�;u;�4*��qn�Y)��k��6���'�i8�.����0��Q{�Q��)y I�N�4k�f\p��V,��c&�C��bYo!�4��.�E�+n��ݢ�ƾ�k�V��ٽLR*��V퀏t����a?��̆|3�emw�����Dv�Y�������}m m�ޥ����텞��}���Ϋ5�,��AҲ߆^����|�}�ɍ����c�7J	+���(��M��4YݲrXJ��6��^��r�$y�8n�0�O�9�轝7~�VP5̃{�(�n洫�ٯ;-w�ţչ<e�Ձ�?�o0Hߠ����	~ŝ>�l0��:,du�
�]�%��y)p����-�����>�.66���`�+�SluW7�����6S@u*�+R�c=�C�	<�6�-�8����P2��9���WW��v�n귰t�+hW���ז#������}.WnWA��ӻZ��<�&�h<���wu=)�|Q
G!b<U3G�S*v��1��^� ��N�~�ߨge�ߟ�<=�ػMw)y�@��I:T��)�M�9E��&L�Zl=�(���� �g>��l*�����\�ӝ��'v�� �v֋��}	bVi�1����@l���(�,`���[��{�>��9��D���e!�Թ�ts����`�xOm�z�N�y����R��#�x�l�O$d��pl�o�=����\o�΀�Ԁ�ieѸ�ʾ�K&ܠ���U�Ryh� ����Q��}*<^�N>ߤ_���>��/wc] <p������rq���;Pid��R��٭�ݭ佯;���U���o��M�dس.���)�p���z:��t���3C��P�7�U�)]�6ׂ��l�8a����g�2e�������@�ע'y?(���|��'��Ӗ�=�:��{�SE�4�Q��3�K��ݾ�<�a�o%$��`���w!Ջ07X��#Kg�;6��W������0��^����ײ:=�**�9�ұ$2{��2)��}�Z�\FS�v�����z	_^�5� �Rzgj|z\Z"m�����ua��4|Kq��{�t��-�}���|KG�楏���}vI.����oݱ�t;���,�cgīu^<���p6?t�N�5���J��l����YY�;��=��3
�i���(P�&�5d�feV	o�6c�:�8�c>��M:7����*�&�bbz�z�L�̩bΥo#�Я��%%�J�: 2�Y��9ͣ�qs�,FG�G�T�޾J�نc�x�»�r*) �ߠU��퐤��������y�}L�Hn??[�h*���V��ٕ��é���ޘ�|7G�<���_9�q��Ig��")�����h��O��t�U��P����'������7�ۺ�I)�y9�EL�ʩ�ji�8Fu��M�L�t6�|��L�0�6n���C���ȭh�m�f���j+yfB$��D\�h=L�tǟx<d2MSf�7����j�ۈxQ��wwej��z���Rĕ�!�s!e�ǶZ����)V�i���B��mކc���a�5��q�Gt,�Agz�Q�kd���n6@�lN�*��Lw��{�7���k�e\�B�h<R�Cb8�&R�H�"dl�	5��\�w+�lx�{�9ٜ+&�m�u ��YG�!����t�S���u!ʗp�ŇlOTUDj�m\���4��j�W!�����l�|���GqF|7����yx��d�kSE[�x;*�j"a�;r�ڹQ��*��|U�Sk�T�����N��K&�'ɭ;�7�,���m�V�C%KǪu3|��V��ҩU�k�h�*c�T5ۃ��S���Qk;=C�q;�׫�b[:�౭=\�oz���}��+�Ii��@&<����f�K��+k:�]re,��C����B��xGg�֪�S���o ��墮�+�t&q��+.���P��O�0{|s_#.͓0<�P�a��Ȫ�c�x6�<�\��.��+ ����n�70p.����[yp�ٛg	p(�ۜ�Ab�_Jä�kV�Z��m�<&��X�s'����Yge0�L��8��Ĺ]��q�0����d��A�viB���#i�"�R<,8rΌ54Tpضܔ��#�j!Z/-��܂=�ܴ�N�.�d{ˎک����ݤ�;��Qئ��9��	;5� 5�9z@3�67�T��8��.7*��u�w!K9�"̕w�������V�֪JW
�zM�"�%�d2 f��e4ȝ��Ӌ��W�;�e9=w��{��Y<݋�,���b�aҥ1�����Fq�T�w��-u��P��r�ڕ!]ƃ͗����n�wU�[�1P+#`�g8��lp �(�k�]M��2Y�
�oWL{�T��αq�0�w��#��
}�pc���%��P%O��u��c嚸�t��A�m�o��Y�� i�d�se�ӑ��
�����ȃ�ev�Ly�Yń�׊P\���Y�۴�>1��t�0k8~��i���\��$��c��Ϭf]��l�d]� j���	2��B}�d&���ӕ`�D.=��֎
�̵�p���f��b3����vnd�*Z7��=��p1��sP]-�7���(2�e���A��H�S���6�F�h5�'e��� P��]͜M��ՇDC�ɐ� �辏�n��\�^�9�볻ٽN��2<w��}�ةI:�R�
�1�3�顶�J�ʑن>�u`�G��;#����f�d'q��Y�4�1uNg�T�zݙ�(���T&��B��ت�w(�>9��r��as���\��s9�%Ҷ
��Ygi��V֍,��k����<��w;�+\�S��r+a1zx��S��ђ�oA��N�+����<̜tTq�k��SYҜ����W�7ٸ�V/?$٥S�R�W�N�u�3������29b򦾃��J�bl��`+�x��h��k�ŋq*��{@S%i�Y��`���P����vCjw��WZ�@5!J�p⢹�����]��ǩ�j�9\먆{��Lu�@) (c���Nq}�T @���j�9�U�ے�%��Ŷ.�����/�f�8�ޛ�������U�Bו��+W]��K���i��Q�M��Ȃ�!��:��T|�u�U�ś�	{Wؔ��Xвt�$(C����~?+X��Dܓ�r�!r�TK��t�"
<�Tp�A	�UEQ����}Jg9^dEs̾a}�%�Z�U(�I�V���QD*9T˕�s$#$��ι%.x�UT���UG
��r��9_D;4A̬�'=�ͅU�D��]�&&G�>q�%K�:��"�*"��G̍y��@�|�W=A�DV�aU!�U9�(����p��Q�F�NR��u(��O�q����jF��>;����w<���z}�s(�qwB���Y�]*9r�̩��9��U˖�n���q��wx"e�%��#8RԢ*�(�Qy�'���R�=�<�=����$�$-QbN�'�ۓ�9�(��[����j�p�������S��"OA9��ޔ��9���Jy�>/r3�F��ą�	a���N���u��9�G�QT�q'	��
���0,����.��������#v�wP'e�l�����p#�L�J�gQ̊Hl�-t�6�sT�m���^T)B���opr{��tp!DР)"�cԗ1r� U]�Ow�U;�`�t��uB&Cuhk7�@��d�=3o��WS�B[s��H"x��\�̷I�nϰ�~�y��n�e�a�Ѹ�yW�+k׋�W�oV?Ж�)�8���Wa1&�¯%ܲ�Q�8�6���d>����	g�7c���Mx<y�]ߥ9��ެ�k�Ry$Β)�KJƎ����+;o���DVj�q�s�+_N��~k�ޓ��,��~n��3��MkN��/i��1&}�}a��kںAZM7GT73�D�_c�'9]���,}�D���n��|69�Pd^+3
������ۋg�y+��L�̿}R'yZ�`�<,����6ʺڢ?V<T�ľ��6�3ᙓ٧�ED�}��@=�OC�3�+���f�#L���>�&�1�)9�S���_�S?|T�gr�"h���Jb����=��~�H:�*Z�%7���"E�7[�+z��^����aژ;7�Q �u����<E�S���,���&X�VWv�<z*=sxu�D��rP]��A�|��$�c��҉�8���R����%$�_U�0m): F���M�{co�u�un$����:��݌.���"����|�~�x(����`s��~C��d%rb��=�����q��;��OW{S��P��ʖP�Ms|�UZ�����;'��� �ќ۬����7jh��[H�U+2)� t�]Hmϸ_�U~w�5�	��n�F�z������GM᭐(��7k��XU��}"8<�ָ���1�[5{����l����TJo
G6��m9��m@B�6n�e��VK�+�7/;���RWl�^���\o��.�лQ���� �E�MŤx�{��n)�ڽY����7���UC���\k����a0nT"�z��+`��iT\a}�Ҫ�MQ|=�Cɶn�d0��������T;�U��O�*�C��qu�����/�T���fy�����ᷘ$o�{d�~;I�Ƹ�5x��tM��u�����D)�1�b�8���6!Yؐ���s=K�L�K0E��ⶄ��Be�)*y��*/�ܔ�R>H��0�5�rr�AlG>8"0َ��f^�3� h���� �©K��W�	;�wQ���-���� "P���WLy���.�2�Y�<� ���].��oH�S8uy�D&���Bv"��-�x���:3cGv��'5Y��>��6�d1���Z��{��r�_C���0�t>.�����f)�:�@��c,#FCr�T:IƜ���6�����vp��-4���R"o�ѵۮ���-�$7��(��w ?��
��SӏV��Y�����S��&���������$c��a�-f���^c�c.�⭚<z��t��sp���ie�F�nk�۩l�Z��FE�ZV���*�\;�n�}7@i�T���,�@k�k�?KT�*Ny���u횣ns�.��[3�~�W,���VW;��;,���� }��7|�Bz�D�M&!q�^+F��;۔�u���fm|��n�r�)x��z��Q�y�i:⧬����v��QG
4C�1�#�ȿ]�&�y�.7��+v�]H޸��V�!��y֜��9}��jHg�K� ��Q�]��|�H�	�jS��2q����ce�YQ&��K7��-R�	�ˬ�n��Fo��sx�+��봁��~<� į�rw�cV�*�p�p�ޱ3��\�1Wֱ���3,Mrj�o�<[��C{ݱ���V����U���
䂧e=�L{��'��jV}l��>s��9q�n�H�sه�놴<5�'��SƧ����Hi\S.���ώ�F�@/6D,��#�GlR���t�¼���	�K�����p�t�w�(�H7���Zdj�>>�l�Zoj9m))�q�[������|�3��;��'VP	sڠs��>��[��XlT�lnT�ЅLNl��9�,"��of������N�<�:z~; �ù@�M�{���e�.�w�p˞����\m���9���eE�� ����{����Q��j�#z]᷑ KΟ�n�d���ǝ������6u5D�Wפ��H����MF�@�u>��f-+�zjn,�{�oJȓ녁�y$��O�-�{����g� -����t�|Ny�Լ��T9����(eax��~U-�\�i���vO�����P��|�q�l��"E[e��K,R#6���u�&u�2�>��\r���"7�y�y�.vQ���o��E�g_o�+��;=#Y%�N�]
�ew�q��|�^M���f�"�1�pS����9���'�;���xRy��+Z����u7�d,	�`	w3׋�#6��kdj�n�}]h�ۡv6�|����s� 	����`	��]в�AmjNвqu�ɕ�γ�.]3�77b;����i��C�2���I�ȿE,:��A2�%w����鬝�y"粛�vREf;^6�`�,�^�}d=Y�.�T��k����թ��G/��XI��]����y�)��Ô�"8-��p�"�B��ɧMN���כ���OXd�.�RΠ!-ղ<�,�`�Fhrd��X"���ȭ�:7t�}��p�yW*e݆�_w
��p6�2�7K�ͧ�]謙��s���!y�1�|g=،I����.������DՙW�3�n�t�6�0pfH[�D���M�-[`�t]x�La;6e�s�*�������)��o�aք�j;��cٔ�N�?r�{m��n�����Zj/#��3�� �Hm�aak̉��2 ,=�y���s�u����>^oO6�[�z�0p��$�u�:�Q{N�$�z�X��b-��J;��N2�,A8}3(t�50O	SYJ�gn��� ���g
O/T�e��m����y�Ry�R��{����䩈���k[��M�vn}yΘ{�Y��A#�C�2�.FA����䟺c�����<��g�|���] ;;9�݄t���܅���fWIs�m��.�(�*6��	��e�����7�ؗ����Y��dgx��^��o*D��D-6���>���Ҫ}��&�P���q9�XP/E��z��\N0����_M��/��,�k�{���C�Z��ZhtdgB��C�jN�Ž;Tܵ�6o�1<�K[�[�ͩ$�Uv�<z�.��q�4�̵[\�{���B|�x��|�;Ȧ�B]M�݋�,��	fU�/T�p4�\�)��.�e�N�o�^��(���6G
7�2�u);��5�F��| ���>C��؆��q�/�&�u�I�aZE`��ix���c+v��o\Ҏ"�JuY��.�z{i��Y\��I՞��1�T���h��Ҹ�ZutnO�F�~����u�h���:�=�W��(ONㅱ�𴮅t8��b�풥=�Ssd�:�5�+b��k���u6n���3��ׇ��ՅJ�Ⱥ/��I;�&����O!�.�4v9`*Z�^R]�>6�j��-p�j2���o#�Rfe�=�p�P&a��X���P��h=�=��yɿ���l���{���<k�iU{�I�+����a��x�`�h�y��i�f���8�m��G��oL3���mΛ会��+j�6���s����6���E�C�����f� ���}W,\L�(�u��q�4;}�w�I�ai~uiPc�Վ1�9�[�l[�ZdΕ�t�p�b{���o'��\���kЭHc!�d;�v�Rm���<hl�j�m�8�.B'�`gpb��2	:�E촒,G�6�ʝc疳3����蛹����������{ߴn�27v^Gr#��!���X�r���wY�ۂ��	���y�w��3�'�ڀ�z�{���Zk�K�r�gkƍX�{+��,����Y�w瓻 U�@Us��*�=�Y~�񹬛��|���q�k����۽�g���
2r�M�Pӊ�-��_�UL@~^��ovz
h1����緡�V���Y0D/�+n�طg
�{�Z���y�Ü��:�\�	7̄�b*`�s�<���Id��y���Y�-��%�ru3";42bn�t��/���{f雝(�p�s�s3cN%p>���e��G������+�ֲ�����)��.��kmނe3�%����=X��9���z�8��4����R�8�gԮ��0P��g�{��u�,1���Ց��8�Q+x����EXc'v�$�e6������˳�2��D��n�3�"����*}f�o��	�R
�2Ry���h���g���m�I�T�hm�fα�c�������c�w\�s%�E��>i<��Qm�hQ��%v �"l�Ϝ�nȽ뒕�Z�A}T����r]�5�ݵ`%�u���:>
�9Ǳ�I�Gx����`��sfww;�"�Й�Ux��l$^���{���V:�q�I���X��y�������a��@�R3)%`N��#�	�n��1���{n��ph�t�,��s�o�m��Mx��vE�6��@Xgۃ:Gj�.N�X��Af�,�n�g��ľi�1Ն�[��2ib���OzK��kGN�=:�T���<��A�S<���<�� ǜ��eG1���Ŕ�:��g/{�7��Ny�]�m�1�'��33s��:=b��n)-�A�]��m��k��Z�#%v�'�[$�{�� �	dA9����.�l���|�Xj&��4oG�wS�G��c�0��Z�v�Tɚk>��p�i4������ <d5���+=5f�EH�~�;C�Q�a��ݕ��<��$��Hl�B.F/�%�l�⮁�Qɂ�']N�PY�ݱPa�ǖ���n@�K�GH�m3����_�8�mK�4p��%z{o4t���]N�x��в�	Amzԝ�f�׊̭�m�[�\DN�|Oٔ��u[98�Eݲ��I�=d(�û�A�z�Q��I�������=~|�$Pt���l�^2�l��k�亽�8����wa����X���63xv��@aVI���Ҷ�uf=S�Sd��E��
Y��n_����M#�Z�;�\�L���q��צ	0��e�����}�����F^^:��a�E�C���&|��fϙ���,̓5�x���qw��J]aE����:�α��註��4�Ꮿئ�a���vq�1���mt7����T�X!�)�ZWe���K�9�`ǖ�/�
�g��(Et�����j�����8�I�k�b@���y5ĕ|r��f�`r��^*w�����M�o��'w�#��{�W>#%k�Kt�ӈSmi:�{0f�fnޙ��h=�,`y\F�Bgu�����'�cƕG>�ͳ7f:&�{5]_l�
n��q��8q����n�cN���Xt(S�Zc�'$Euf�������6�F��i�5�`,=�/'E�k�ݼc1�v��Vns����}->(���蝐\�{"����66E�ϥd��<���'��NaH�n��m�J���Z�2�7�-|���鶪۾�wk]�Hx����wa��LQ�+�L���\&�u��\��qe蛑^��pU6z=u9}�ZY0�VPN���Ŋx��]�{�
�65�zH{�d|���5�g����t�O-�e�Uj�"K��S����N9'鸍I嫸o�[����R�EMr�6�=�x�|����g��EÛ?����V%�c`��HC��2��g�I
'�����[���}#�n��ӕ� u��n_:ǲ��p�\M`��
ߘ�](�]31,�ݛWyp-v�XR��gc�l�T�*S���c�-���b�t& ����iwS�;�5����K�}J�q��������s]�X��]v�[@�U,F�Ǝcavl���<�6U�'":��,�Z��G$h�ӈ�dipB�0��YbF�f�ې�N�R]�1*���3���d�/�w]� r�MR-C�9^k��m��e4n��2%��4�I[8gB�qjLkEbJi]�鴭��ct�lݎ��9D3X~Kg�9� N�yi�,h���j����sqg,��㓚���S��^Ņ��7�Y�U)b󤨫�k�����s���ˢ�/:��&�wY���"�L�h�`��;#�k����t�'\>�|F���`<�f����\�R��aq)�+b�h`��Φ�)�T��&��اY3(��e����ڦT6���s���CO^�v#�AwE��N;�:��Z�r�N�|Rx��ٚ�J�c*��V��<�p���U�m*�a7����s�'Vu�DL�nok��5�_>��_Y�D1X��%v��F�eݠ�YeT|潫���F���$���R�=}O�����a$ޭ�ӵ!u����.X�3�6`�[.[BU�\7X��n��+��:,�G6l-�������U���X��(�`̬����IA�v�n�F6����+���C�d�3��#������×�i���1�����
{��,�v09N�5M��VƘ.�B�d[7��n`OBȾ(���.�%��h���k����<�*��K�,��39���n�@�k�5�̭�k�;���k%��l٢�j�#'vXWМL6\���ëF3(�U���wD(���Wy]A/��eI��=}-^�o(�+w��L�s�s�-^E׫p��+P�94��q�B�
��+o��*+�)K�/ '�m�}��w���� �
�K����õX��+6��Ŕz�V峝�8�V!�d�b���b\����A+t�'v�+($=�-�Ge�|�Z4=h(n|���P[�Y��h��$2��.�*e�o����e���\L<4�l�FWFrY�m�_R�'�7�j錺��ܵZ��R�����mjrX��ɸ���E��>}}ԅetEM��9��g8=��P+��6���V[�y��ܕ9A�� wJ;�&B�u.�JŃ���.sB�Q�9s_=j�}��r)�%5v���Ę�xUe�/5��}G�]��ݦ^r�M��(٣a"��ĲA�Lq���-�@_*��2u�,?X�Ԋ�S�㏳(
�HS]%C-%�6��rQ�U�#�WpX��C�{o&M<-�ZⰹQ����.%��y��|ˮ�%��w���H8[��ԁ�bSm�"r�;��a]y��~k� *�-�ʎ|��\��pQ�Ā�O��>��,'��x�:�BNy]Z��rwstL����`�S�K��*��^�%�xG�B�^�<�蔖�W��T|ʊ���CܶTy� ��6B�wR�OtB�Z=H��M޹�ȷ7�ޥ��V�^WN9'�Ч6\%4<��EY)�Zy<��tG�[��o�o|�:d��Ї$�dr�p��FDAS�C����I.Kdu���tU�O�f�BT�^/{�}㎐^�|}�>qu� �Ֆxu�i�E[+7�dr���X��P��'1*W���s�f�<�9:������0��^%.�r��k�>�=kq$]eW������[���ώ�A�ww��^	8c��P�.N�EA�wُ'���W�z	9.��֐_t*���ß��{���8�����QE�6��k��tTCu�f�Z=_g������YX[���UV��O"�����.��!��"�F��0E�/i�\Nn����"��P��ʀaU	`�
�lba�-��6lԥg<��
�u͏�葲L̉ՠo1n�&��&M�]�}�$�Y�=c>��U�W�ǁV�d.���=������;a7'�t5����$Ϙ���uY��Q����ve�4�[�C.{S����hd���8�"7R�nI+e+v����G5i�*�S���G��,0�{t�T�<��p�b�T��h��T:�$GF�Ȣn�K�A�d����l'�#ݒT�46΅���<�z�`���a1 �$͐��cVa���qL՚r�F�0��<�Gc3��,����1���}�?v`w��<�-\��A+��u��(�~�{�D�a�����m�s��g�y�����2�"�6~��y��yYZv8B��%L{��8�m�Ot�̝�uB������|��ĉ�c�l%��h'R�V���3���uڱg7�M)���[��Ƅӌ�03����7:	8�E�4}�FEi��n�M�@��~���r���?qۜ��14�V麒�{N2y�Dld��8Y�+����,��3Do��Yd�t�#S��E{S)�H.�=W��No��<-�fG��5շ���K5��<g�殮j�XČ_^��`��w�a���r{k{{���߼���}�`ّ|�tln�� B�����2ﭓ����g^�A47&����!�`��U��]{2���Qj��0׶d�ē��V���n�#�d�V�]M �Y�9���*�Ε/o# ����\uAѢOWe��չA=x�@}S�}n�<��d�	T����ܜ$��ǳ:γ\��j5�j����J��[f� J��̷];�v�����V>���$�$N���d8�:[��O��sz������]P�PG���qD��6`�y��6����~g�Z篜IgE��T+vF�7m������ވ�\��a�k�zg)�%�#����;����s��R:�sg#Zv��Ǜ��9���nwy�& 7;%i.�<ݸ�VS�hW�H���b�ս�A��~'WJ7��F+m�f��ކ9	����}J�����6,���u�Z�jS��S�Cxȫ��:���%�i4�F�K�t��{��2��7M�kha�&ޜD��ޣ���j��ۛ��n��U��}�eo`�Źi�:�r����h�h� �2���h�c���a��=��7Cs�HL����x�F<quQ)D��2	�Yii�j�>#y�0����̆��d�gz�S/4��" ��v�um��{���Β��ޞ�f.M��el^�����)kO�r�}73� l���g|N�H�<�ߪ��a7j�vE��vz�Ҟ��f��}5�H}�a�e���[<�����,�+#�<�{�|����|�ڰF�c!����C�G���,��]7�4L�0bF�2��c��mrv�:lq���S��g��Wt�KI͵��N�܆�l=9��/��zF�<{�-��Ϲ�b�c���[>>ٙNٞd�m�OfN4U��n+�J��r䔶������)�F���Пj��De�9�g��=��)k�@�n0�t,�AD��D��E�n����666�%v��������j�����ȴ�)a��k��\�5�nE{H�i�����(�T!kO�t=9b�e>vc&t��G�Ygޜ�7�]H���)Ŷ&X�AT��:[Is�}���RI�z����r㻄�Z��� t��dM�Q��.��<aP��Ig\m�E}�<����s*�朦�숯}��߿l�eʱ�j�ѭ�^�/��g�6���
��g�����;���.��R���v�8���hv�&�M'D�[��=��!��Z'�n�i�q��ėox��P����f�y9��H�Vh6�aWG�ȰOz0d��֧ۛ�^�\��y��������udX�BhPS�KeЌ��DAޡ1��gmth�*%ܲ275t��sW��PƲSamˡ��Ԫgocy����_W��s(΋	wv(�|���>X1�k^*Q�M}������~���k����n�M4�q��=m��tA�W��Ͱ�d7g���e�1���9{����Y����w���8�ө,��$���9; ��7��2 ,�R{�!	{P�~��&}���i�s~�#��ΎW� �m>2�쳧q��u9�ַ�n�#2V��,�en�����}v'���IҺhY7��k��yiku�ɭ+��Z�U�Nvl���s����"C����b�����C�[�k�{�wh��ړ=^	��3*^�f'I.�=�N]�j*g5��.��XH�A8{��j�<���ׄ?m<V�ϫ�n켎����Dd�C2R�eƱ���)��۷r�/l�sf���Ћ�17F��t��F�����5Dvb��<�.��4q�ݙ>&�H��u3�P�R�徛��J�{.�.p*��é�I��'n��L�%\��+�x���k��cJ\�T�"_oqͫ,��Q�����7\I�d�*��Y�@�x��Q8\If�<�e=�M@h�f��K1Bj���l�4���G������n��f����,!�n/S��9�:h�>S'C���o�Һ��J�Jݰ�Į����i��l���7��}{�-�޹��1P�u�u�ޅǀ.��
ؤ���)[T՜/^�+0�A
F�#(7oL9��Ǳ���������A����>�i?��{��l?1����E�L1�!s��x�w�Z�U���)�]�յ�E�G��$.��OW�[�B(�M����?8	��^�o��%�%�p�3�^W`��!̲�ocô=�P�k��,��{�KD���K��Ƨɯ=g%iW����x��qU��u�B����Wr�b�������������!^���i�C�����m%����9�=Q��=9��W������r��<��/�!OJT�G{S�(&ͦ��;rfڭwwL��.:�r�'�L�׼{)�����0m�9Ɨ��T� ���ۛE�?��s{u#�ؾ��G���%�lc���;�B�a�j��m���^��m2�-<�Vf&�V��������-Ƣ�f�����X�ն�5�
=���#ǩ���ς� ���tߧ1j/�luY�;��ݏ����b73u�i�A�X̌���!�@UO�٪3�&�Yr�(k8���m�H����)�jn��[����5N�qYB",*�����i��MH>ݟ�
͓��.��J�Y�
��9�����6��9�V�f�fq��9\�^Sd�!������F���������e�yBG�U�P�3HC���p�zƕVn�ֺ���Fʑ�Ze�<��.��z�}"�U�ISp�e)h�U�)�X��V���VԬ�X:��'b)�0�xfŃ\�^����&'�A��n3;4��Z������v��Ȥ�˜M�0��Ik�T)��n�H���o�1�6X�Ϭ�{ūܑ?_������B�6�\�L�(�U(�6�Wr��@��Ϻ)��?%�p]"���n��9��U7g��ۻ�$��V�ݹ_[�:L��
�'km��f��p��S��C4�"��֓�k�#wI���>+�+e�#�ψ�� 2ޱ�*Vt�����ff��|�Wu�+`��e'�pW�du���-�F݌�\�lzڔᵵ�No�O������Nj�|~�9�~�).{6к-����M�x{n�z@�>�"��Ĥ@��P6�<�vѡ�.�2��y~�cïl��R٘��;��q;�a�ȶ١Y�݋a�+�C��z�Om*�I����!+R�CF�_H~��ǡa{*ZZWmE�m1<�x�8;C�� �'�R���"�4�Q�]��w���k��o���Z����~IZ���WKr~�Ҳ��{�!gKU����4��=�����J��]����#�/ �K	�E{jVM����t=.Q2�./zY%U��w��	^ު�ȝJ�_Z����1�������ܶUN�:�Ҏ�v��'���Wy.�p�xc��Ꮶ�@���#�d����I�G��1{��R�zYd5�$E�S;�<�����~��9�Fg�sh�����%�U�j���Lϊn$���s��^��g���Z��x%��]�S@xgǡ]0%)Ϳ0~�;X�&����j�iμ�Dr̮�g�a��Q̎M���K̞��Y��)�8{���͢ԟ����H&�PK1�^2��3�v��E����z�m�qwk�v.�0yYT���+���mb���RW�̨�`��ct�5w�+>l�h+M���h�n\q��\�`o\��C�kRXs�o_�g���!� F��w��_�s�<�+�'�ؕ���b���5=�EQl����kq��ɀ�y�U���Bc`nb���>�*]Լ���Ί����S/3/���k��"-6v�>�n�xʙ�U3������nz�٭F�fzX���W�'���BJ�o�;N*ͼ7�%��]�|S��R�r�������w-9������:W$�>��NZ)+���O�А��R�>:���lD�����޴��I��nd�fu�B�:Vi#9Q�[U�3�l�64Џ�7)>�{���z�շý�݃y��3�)ц��.����_4t�b���1�զ�˘��4��k����ш��D�C�v3S<�۫��h�����.~�Sbn	�:�>n��F�gHq�i��ؘ��1_f���b<�"�oA�${��6�.��F	R��YM2G�<%��g�A��_a�Í���^(��ʆa�݇�<(��!d���� ڸ�GL6��4�#l<`�5�bn�FYδ�Ȭ(���Л��A��9}͎,��t�v�I6�9�̽;2����_�Օa�Q0رN_n�]��8@<AV��UJɟ,�x�˧�w 1��Й��g�x���ֽ�M�����&��~�4g�YU��*�ǁV�e�gcÎ:a������44mX*'7�D�\�-D���ȓK9�^�1w·��3/c��V0"7ٿ�\:����K�\:cD�M 0cGT��[�r��ɻ5�Y�q�qV1����i�h(n����#tM;�n�AeT�\�i�R>�q>��uA
��5���н���4�����u�u�@C�gEeLj�L�&�v3$�ܣ����A��5R��pq�|$r]>nI+d�ߒ�fl�Y�H�j����������m1��ϐ��i�\&��k��#�o���Xc�Ψ�B�Kk�@�RiyA��r�fh����'��R��7C��dN@����,��ݵV�/�z;O��c�G�	l��abfȅ�1��p�6FV�?V'�{8��5Cv	[�s(
�,���۝����nл/�_L[��Y���a^��(�{�^��Xmi~uiS�{Wn�_&�F�;33��u������>�6������V0�U�=�ӸrF�\>K���b������<
��@n	����_v"Oci��X[^��J�y��vH6ޥ�+��i�S�{��K뵗�
���*tlfar=��G�j��$ɺ��3,>� �khX�c[�=�5[�������O����k���6��v6��o��I�;m� ��c`6��|����`v� �6 r`�9� C`?`�����p`����q����m��Cm��7���v6�ɶ�9�m��m�rm�� �m��;l� ���9  rm��m����9��g&�l�6�:�lvv�l�6�9��n�q��Z` �v�m�1��u��m��m��Cm��6Ð ;l�� �cm��m����9��v�l�6�9�m���m�� !��ɶ�9��@ ��g&�l���r97�X3�`=��1gm��0��[���Џ��ߵ1������r�!�ߐ_[����������>��u�(���O�������8~����%��������G��m�����@���g����?����6ȁ�����C�g���.����?V�x?�6����C�����@����~? ����&?/����߯X����� &Ã  ���m��lle��a�` ��C���`@pm�3��v0gc G �7�������=����)�2�`�~f�����g�~`�����<��?�O�~?��?� cm������?s�������������������c����lm�}�����?F����8��cm� ��o���~��������-����ߘ~�w��66��~@ [�n �?m����A������M�w��p�cm���H��?������@��o����(�����A���_������~���?P8������m���I��� 1������>�<�߷���?h|l�~��������~�������o���9ߖ�����������_��[�~g����G���66߸�7؃��66ߛ������������PVI��Zs�� �j6` ��������� ������(���JDP�T!T�	TT*�D!	((R�JEB�UJ� 
����$�T�B*��� �J��EU*��AB��W�jHUH��d�$�J�	"��"�B�Z�V��&�B��DD� J�Im��H�AH��$�	�$�2��%
%Q"���B�HT�T*%)"R���) �J���E@)
��p  �v�fU-�b�h[m��Z)5SB���`6����P�@XV͍4cb2���45e� پ���T����ѷnt�U **��B(�QB�   gXh]�
-��a�s�(vǡ�CMP�y�z(v�
$[Ҝ:$vč�!��l�ԣl)BʬmYZV�SQ��V��h��(֩�fFK5m
JԲ�-�ږ���U
J(���kT�p   6khf�������&�m����H�4�a+5��@6�j��wq�ƫA�-2�YZk@i��&�ZM��M�cE�B�)APR�UH��x   s�V���Ԍ�m5�m�3@�jQ���%��[Yf���j����RV5��h5���S*� �i
���EUl���%%T�*�Up   wp�E5�icT��Ѣ��
Փ��QJ	BB��f�U*�)��F�1� ��D)#4�J�KMH�P�URT�  �
��X(
U��I%	�@���APY�բ����(hY���ԃ*�	��
ڀAPQ%)IB�(\   m\�%VZE �C� 5j`*B[( �4�*�����F�`(5T�J�r�E
�v�8��QHT
D�TP��   ���BJK�r%J;N8䦴�.8�UAR�gl;t�R*]�UKM9L�̔J��ʡD��v�u�v��r��R��w$UH�Q)T�$%D��  6�zB�T����J]b��%RE7Eg)�E����m��7D�Q�:� ��n�)*����V�ն�%R��;�ZД��JT�QDR�   w�-��hn�X:��T���D�QUY���jUNu;� D��R�܋u�넊��u�)wlv��6�\�Z�U���R�(0� )�IIJ�  *fI�(bh  "��	JR   �o!���A�F�e*	��@ H���"2q�Ӛ���Khr=ȡ�Oh��arՊ�XA+]ؾ��_U}�W������f�o&��6?���cm������l6ɱ�m��������{�şʓ��L��V����na�`l�v,�(�k[�J��(9V�6�%���0�wn�j����4���ʋpR2�{���2����
�Y�|B�)|������@�Ujv`�GrM���È�U0��zl��q��M�c+j�Q��:�^�^�������PՂ��1���R5�Y���e�K������eks/r:�w��b�(Vf��+
zw)�L�Z��`f�ܖ���[p��dY�nna&��l*�+F�QQ��&��v#�˫
���� *�ZcD����J�,S�Vo�V�j��6f4�u��#&Zva�zV�)��~]�I��*ְ�mԭ5Y����˗Cr��׫���Ϧk��Օ�YgR
���D������N�G��!�%RP�M�k�7j�̢��K2|�f#3R�P����ڗ��p���P
�(f�w��r6hը��0�cB��T�kP{������uɺ�����(f�G����BR��l%�AL�Y+
d]��Sr�l������Pԯ*�1�3N=wGC!����-�EO�L�t��uQ��a�2�cR���
���(ݍ����uc����6�����ח,�{�)P0���(�+ue	��LA��f��6�D�l-�F���V"�IxL8ޙ�U�^C1i��jEj��I5d���+4��N�-8 ��njW�M��W��fd�r���=�-*��w�UBf1*^b-�E��N.��7Wf1�U��R��amӷ���S�M�נ ��ͩ�-L�Q��iz�ʍ^�]����x�Ex��7n��a��X�)j\��I2�=�.%���F����T��j6�����U��w%g�Ncw0F��ǉ�JX�S!�����9f��a�9�v��`A��麗""�lø�R�3��CY�^��p��a�#n9����?M���=3%X�i8Bn���i+t#n��uA���fT�H[,֭�O �v��T�D���veM�N'�r������^T�i�����y𥒖^ޭظD6P�ji/��a�*;���ʶi��l�B���e�k)`]��&���N1m�-n9�@��5%�j8r�x,�դk]��F�w�%�)�g��X�[Y����r�ጞ'Zխ$颠�C�5�c�l��Jܙ�ݥj�m�m�8�
1V݌B�%,�0��1l�/��cr�a�o���v�YtѪ�+E<�D�G�r�`��F�1�w��c�mZu�
�G��[)Nf�C	h��t(���m�G��,���KA��V��^�%mYi�g/ul��V��rRP�jw ˻���r�0
e�;V�4CڳӧG@6�2f+e��a�D�f���P������2	zU�Gyx]�]�;�v��S(�p�������+�V��J��N���66���&�VK���g,�C@WcV���L��%����8���6��D�E��l*��H��'F�X)�5b�n��;�y�	/V�a�}�l�|�-��U�dU�:�`��S��0eU����%A��
޺�Yuj?���WR��0"T��U�i7W��d�5a���C��w��J����vp���� 37@�m�:W��%f�j�R���j�f�P�j��d�N�8fS(�P"�"~�5��76��ЫT �j��2�5t��Lc���o� ��g(�I��5m��7���eZ�d8�ڴ��U�����yQZ�`\�,�A�;y�p�˗���/��n�9x�њ�d�-;��j��jȫ���N�1a�S�q�(&�z.�f��4��ސ�U��� Z�5��	��3nԡ�i��S���`֔������`jU���D�>�izN�]e1[IMI�̭�x&��_�TzY-h�S����KOEL,�\(�J���ޜwln�j�B�U6%�ڄY��-�P[rY��j�����W2fo�p�v�rc���8�VC&�tt��Z�:�)@��yN]Bn��"P��LJ��N�ek�t�2�e�e4�H�N�ki�e@��X���q��m�X�f�p���L�Ĭ�<rc�B�̼+�]m�跩Ղ��q�T�w��:%dH)�jP�Yb�2C�^�����(�4ܤ��V�a74m��nR�qi���7tZ]ٷI!�[�x�K�W6�*�./��a�x�I�JTڰ�AR����h�Ú�]ۡ�c��U�1�Z��#"���n��:�M�.jY�.%.��)���Kenm��5y3^����1�3n�-�MM���ݡt��3(�j �t:7̚���w�l��hF�X��#wA�m]u�w4�%z���3wGs0����Z���e����5l��V�	Y@��銡��@��nˠ~�3P���%m]ʁd5�L����
�m;�Cʗ4h:�[!���bX%�='(�6��1�0
k,�H%2*{W�������	�v��`�C�u�"�^n�L%Z���Wu���FX��U�m�����n�Z��PI�)���Ej*u��t��6�th�"�5L��f��)�t2[������F��h�,�Q�<O~up_�R��eh	K*�<���썆pA⛵�-�ͽ"�R���yd��[��'K�K#+5�T�A�7)c+���������)zkK8�����1%w���2�]��#�Ln��i�N�.�۬��/xm�S^���B�˻�Gf���K/asn��8��oB3Sl@c�x0����\n&�����܀��[nemm[I=N�W���	���r��-��HPv��b�e#��w&�r��wp0���ԍ��\�,軎�Z��HI�ě�ݬY��oLIJu�#a����K%=��5&�a��v�8v���4�b�Y6��SLS�����n<�]��yz(TH/v�;=��Y��Jr�j�%]p ^!�̭V��tMÅ'�&n͓2�]�#\.��҂Z�YN�Ix�r��Pd[-����d��M9n�P(��	9rclA{M�h(�KE����B����eڙ����o5eb�
��[����d�u�e�؛(b�:�)�;�4R�����%P�3c�%�um�����VhMx�$Zm�%]Y��t�Ӻ�n:b�m�5���Ե/������u�Ժ;&�4*�{�P#%fT����4@)G��bղ��iL^�UD9���HKe@��r��ܰ�U��%A|/@Rii"���jil)��Xv�kC>N�Է7��z^<s7�Xv�ܶ����++vš��J7�3v��n�������5n�k���Z*^���!Q]M��$�����e�Ր̩.ɟ0O�m��a}�F��H�tv��.��Hfb���cRtm��f��/K�a6�e��F�f�-���r�'p]@$�Wg,]N�f�!�k\{W Z�{�e;Դ3�=�KV��tk����x*]���zi���VP�mR���If	 s!��9v��*�V?*Z�#�;��0F�1Zl���İ3Nn�kV�e�2����6��N�y����K�(X��yd����ZAdˡyZ�z�)��"�{Plml{X4*5��`��܎uVmTt�KbZlZ��9�ޅ.��Z�[2�x,8T��)�!_3�yR���pL�I�����v#H�J��sL���)�Di�Wa��N�ol:B�H
�cx�=��������B�yIЗSF����i[�.2G&�h����B���Sq�m�n�l���n��4C��&���-�sU��\���1�Ú�Q�v�+DGV�1���-��6�e�[��^��谥�ӽ�^��c������ܫ�)*Pcs�e�f��J�V6@��!�)6YPM��&Զ��6q����n�9*d�Z9L��GE�AZ�YX�'!{�[�["�cmnH
6pR�#�vV�`G��m7�n�d8���LT�ә���c���ɋ$jS��c���ywya���Ʊ��v�]�A��Q��(�q��&�Su�9NJ���D*O)V^����fB�*��͌lO6�Z�ڬP�;N�օ��e'u��vH�LQ
Qc�Y@0&'��eB]��퍣�"xڸ�kd�����1V樒�YdeY��En��-aW�c�J���	�n^Lb��i0�ӌK��ӣPR�A�ZW���V��M]]MK▭=�KKo]�G/T��N�Q�%����`	����vr�E�ՃBؖj-}c���]*Oi���yce�DEș�x��;0��$R�L�j��������6�JآPw��M�PF�K1���<N[����ڋ^�̨��:e�3*��3]0�mII����
�Z�y-���m
�KKx�q6Xd20a��8�ͻP�.�	�d�&�����B��P�3M�+B�X�*R��
xe��,�ژ��jY����L��&��v�(PIF�hS0��-���i�d+Idi��ȃ*���*F����M�72R�BīQ�� �PZV���g�o5����a�KQ5�չ�=L��7���tL�6�o.����WI+���<J&�e-�J�(�]e�0'���ܴd�l k))BLϲ�7��n�D�!F��~J�-D��iS��ǁS���M�f�K0Q�j
9�����є���̢��kp�{�e�մX�yLF���Q�q�Z��k��zc���Ʊ�n��A)�Rԕ��tg^�Wsy\��P��ႜ�JUhcH|�VR*�@%��,�D��9p����<K�['E�h�Y[An��Z�Q�*�Dڴ&�u�ֱq:���X��9[*A��6�� ,Y�5�AYK3l*%wunU�%V���7�N+4��*$�
�pˢ�V(O	��M��T�1f��r���˼����NҼM�aH���+f����olR۫��볪�`�1�.Tq�0jj���1,D0 ���j�[y�y,���fl)!��
n�t�����[�ۂ�)�5�$&�[!5Q8�|6i;ݕ��ђ[��๒|�K#!bm�4M��i�Z��g�b6�k��rn�ܛ�&�"T�շ�O�J��L2k�ȍ��)�: ����%�˺4�٤��0��X��e(Yfa����G),��i�7!$�(�F4q�]ٷ��1q���(�$�R�M��*P�b2f�bz	�w����-�]�G,nby�oq�G��Y�,ӸM?�m�nӽ�zE,�g!bm�w�wgGEҟk$�W*�V���","�P��׊�hrR�1��,`d�q�J�=���Qbj��.b�w��H*H��M]�hjƇ����UkV��]&m��ի��qkva���^ �Dn9%��(��e��R�]hDL�������x�K�{()ulF��\�����j��e� cAܫFV� �dN��t[J:���CKw �W�N��c��r��.�@��o/Aˬt��z�#^��!�<!N���`���T7�-�k��I��Э��r����Y�c�Z0+�xK�dj���}�!n���4�szIE�Z#�#jM��R�Sъc��:���F��ſ^JXX�p�&ӷ�&T�ݏ�2�����4��h�X���O~(�L�5Լz6;ԑ��U��"B��R��me�B�v5�qRAݜV2�x��w��B�.b(� ���k$�#��J�m �.�!�����9yҔ��$�J����օme����Y4J����|�0��(�ta���}�N���oN�3Jye��hݧ��a�� +�R2r�ٸ7X1��9���l��͈�!R�t1��!�E���-/��5�1��%�

u����7*n<��@"�bcK�۸��Ef���q�H�ͳwY�B�e��`bR�{��,E��*!X�-(7y��K����Ac6Q����c4hNg��ʋ�[m�Q�Y7PMP���m�ŵ5�{v�e�'M���K�r֗f�k�"�[�
�K�J)#ln��ݔ�Ly$�-*��
T/m�eo�6����Z��x�r�M��u�Qj2j,�EL�E�����`��lR�VEJ�����5��P ��������9Ku��ۚ�㙢��д�4*��9t4��YH�,�aV�bm'`S'](�(|+n�ܴ�8�����,	&����[�mS�-TZ�8B%��R,ϠZ� �@�����@g1
�Tٳgp�Ly��V���K[a�m��b���$&�1��܇m+�-��p����X�7Wrm���)ҧ�h
[y�ԕ`!m�N� �wd,�Ê1�e��S�۰pY�=*��l�7����S�����[t����Y��*�M�*PA*970��&�ӆ�WYYc#	$��)�I<f^�o ����C-l���E������b��� ��b%P��ܨ#ajB؎�z�"�-�+~��=yxMZ�*�V�L+pn˷�e��w�Z��j$!�)ֳ��͋n�K��j
�A2Ԅۃh-?<�������L�t��#�ݡwj�&e��qQU"� �eB�k]޼��7�X �hG�n�֒��ܡ@�Wr��)uN�b��Q1����4H1�b��م���C��R�r�Ig�VjjIm=r��MkDN�A滽���4n��QEVq=�%8�%�l+��n�-�c�A/ELotIW,@�+(�]������Q��2�7x�"͖�c�p]��F䒐 TյOq�U���"���*��p[W.�W�
w&7��̓+Qс
������L'E�L�T�q/�^!�۸�ʛ P�ri܆-���D*<�b�0P�T�Vݿ�����%��T�@�귻L�]��C�0�N��8޵+���i��֦�na�8��_fEh�;��:TK6��*�K|[�[���i����*���V�|�&n�!A֛8��Î��rg�j�7M�/'w����NZ�=i�������T�\uyP!bkfo���a]�]�t���e]��@��Ȱ)[u�z.��E��-S�|GS�J�P��n�Ǻ�ؘ��v�hw(LBt'����vZ(�.>��]��T��W�t������z�Ԭ�
SH��>��ngw�e;5Ȅ`�eИz͌y�6�Md�ܺ�򱮢���η/=�lm1Õ��[���6�ۻ�GU�zv��]�4>�����ȥv"tz�>�w�{����vk�5 ���7G�&*�sh�!��jI���;JpzPR9�U�FU����e�ں�����7�7J�O��,�� �^�b��{V���bWC��W)����0��"�'Z��wl�HG�-YF��zƽ4�@(�4
�S1�<p����*�j���i֋�y�Ms�Y��ؘ9�����3�M1�ⲮT
�쮫���;ˇ��du^��X�z�m��ӭ��޳�����m�J�;�ˢ��e����5�������Q�hZ|�!��
e�,}|�l��NY����Qyv��9°��`R�)e�0��U����x� �t܋.�q�*QT�^MԎ����^�������Q�\WU��RX)h�,F�>Nl�k$�T7��L;�殧�qYb��^�^� �U�[tE�^F�/�Q[ף�a���n�J�j!̌� �� �+�h���9k��yo�����m�LY�#FN&%Ъ�����,�:�C �1��Kz��lp�d�{#t6��c�l�r:���.M�+��&�C��D��#);��\��Ns!�k��T��.;/S��p�y{k4�����Y�4�� X|U�3�)��:r�6��[h.��ӳ6��7	º�K�����[��\���ڹ�ڹt�Kuö�:�zu� ���L�|EJ
���:�}+��F�q�]�K��"�6wMe>��9(�6�UtB9��Ρ(EW����r�����f�A�rgR��]��!j�\g�B7�X ��W�;H�e�,�(s�l��l�Hyg٧P����]�b�k�N�w@yX��ݽ�z%y��h|Z9��?j�G0䬬�Y�>��B�s�N\��nr�΀@�D,v&/yi������E,�γ5�ĸd�7z��Y��ۣ: n�,�d[��I����i:�,XL��-d�%����05�Xʸ�5G\��6T�0��dYd����!c�m����ξOX�z�8Vx�]�k#B���s��mtǩ�Y|�ޭ�(����N�J���BX��t�m�������R�ȸ�P�<�&�.a�Ըw<�X>ݢ��M�Y�w;zA�-�� L�}2r�]��&1���:h\'^e�|X�s�V���{��4��v�]8�f�ߘC,�|��qn�8%i����뵭S%|�c8�}}��VlX��a�y�ڝG���h��f�,�o��ff�!���l�/�t*3��h�RSOvE���V�9\�m��*!��u�M$���l��Q] ,p����b�A�6�Ka�	k�x�	�BN�tլ���4e���DLY��\^�׆�[@�B+X�`
R�$�″��C<�,Tid{���m-�m_R�ͼ����^���.��p�x]`c�8n��
5h����/��Ѝ�+���
����s��8"� ��o��;6��ݤ����,�%a�SB����,�W˚����b�	,�k���p��q����V|l�}trC�(u�k�N,L�5�{\��̓Fc�$[�ƒ��ɖwW3�h'��R�F��N���%N���r��+J٣����0�7D�>gVe��@N$v�m!=�.N���c���{c���fД̚��N�X��Y���8��P/�èO��Zh�ɘ{VJ�j��<yks��j6�ָU,6mn.DU���]eż��6��A<�m�K�N����9U�b=�s)�����u���t�m�y]DG���(�K�g����]���#x˗�����x��둵�ޛC3���z���:��g&o��l�v�FT���q��j2+�{G�5;��wυ�r�^vsy	��$qލڪԊ��0c6��:S�竹1��Q4h�o����K.��td��>W8{s(j'��gj;�Ċ�]��=�P䩛ˮ�+�����;X�a�k�\	�����^��k|�	��V�t��"`<HwJa+$����
�킷�D6�vd�W��\	�B�ڀ�� H��-kege�*b޷K�⸪�ՊB��>ך`�v�})TO�is�S��c�'e˓0i��h�5��J�� c���4N��r��kПV��W�S;[��3w�[����GlN�h&x���u3�2����54�"�d;�}�z���3��J�w��t �D�<�R�����Us[�RPy��� _eb��r�
;wz1tI��w��P��}[I�R��b�8�NpI:��iͷܥF`N���*��:[T��jO�2���p̀A��`����p���MwPQ�����v�8��wyΐV�gT9��4y�������a�z�vM�J��y6��H\Ց٭̱2��:���>�=���	m��RXK�<���v��뭭ޔ[�ý�f��!���f�(�蕨�c�����l��2_6|�mx�n����"��3���]}v��������zD�����-�]P+kl�r,�P�x�C4	ם��Z:�;�Sh��w��e�*�94jEٚ�XS7��ʈ�����ج�_-�]j=����Ցm
=�se���i�o�[�P�G��3vk���P
͑�:V]2;ˤ�]ގ|Nn�Z���)��|�_
T��n�qZ�3��{j��C)=��5���Yt�"�ò�Dt��FU;��\��v�N�X*����i��,şl��J�
�X���ܧz�q�)�`JrB���6�۹�7-YQF�u��i��]�}p(;J�L9���bn�]P���ۼЩ
�����nU�Ź�iz�9�1�E�Ō���&R������ޖ1�tnc��*5ۘ�RҸU��v�������(�6@ڨ*�e񠷐�y����PՃ;e^�qf���G<�t�irRSC�a��e��V��G(�ݔNLo*!��\�Y�9�%B�x�=�����|�C��-�wm��.�y�%�,WE�6����T���[�g�{8�L��w��+z��8,�hѕn<��RJL;���Gp_F�Q�(�Yrv���¾z�52YЃ��q�b�X�⠱I�P��ch'R�خ�1ǇS]ڮ�)0��r:�v\��љ|H�q�7u�:$��6n�Z�V����I3m*C�"����e`&��i�:֠_K]Qb�x��o\�Ӗ��_e�z%�������fv`�87�ےAL��4�g�ۊ���#r��źLدrE��̵U� �Ww��t�4��h8g<�f�u�!�)�	�W�����8��֋G��;[�ݘU�{�W+�Q�u�ݪ� n�5�n��jJ6�v��G0,{H������^������~�eV���'C���@]�T��p��e���x�9giC���
}��)[:�T+�5���%]r�i��5v��В���S�a�"�4��j�!�
CFϡ��\ά`�GA�x"���
�d��Y]\'U,��&ه"���o����l���S]
}���}�����"���"zm�\�΄2<��W,�*����D��e�1�xY�m�Z�X�T�	�]�+�]�p��WV.�=�­s����4k�%-�Y��;n�>A�b�޹���Z 5qz�Ӽڙn����k���]oP�|�(�QdǤ�HRQ˻���޶/��WKO�;�3�PrK���v:7�Mc�G�ڣ��ޮ%�W,�� ���L���u���U���*�MۚZ�H��p�Ui�5ڷE��*I�0c��uwV�aj���]�F�ݤ2p�NX��II)��J��<ՐVWX��x��m��㵶H�r��Hw1t��7-��λCy��}z3�5H;��K�Q��"�RC%,���PYWq۠�e�����)6��ݙ��F��Y��]�y' �#6>�כ�]�8�ݵ���G5H&Wl���ŵA;�}�ʼ
����c��u}5m͹ܷm���,Փ%%gzɈX�C)X1c�}����f���V^�.C�	���j��lF�͖{@f�sz�ZΤ�}/�ZR�-��3�}�a�BvIe�s�^�N�[�b�RD�eAюw׊�K�
�;�c��n�'OJ��mlz���t�6^�
mj��x������6��|�K��
��t���6��:#:fwsE�Y�۱��/1c���2T�W��V��=�mp��	vdࣴ���: ������<�J�df�l8�l+$��_�%�U�(<��P5���L��@oS�`ޞ�Ǭ>z��׎8�p|ސfC&�ˡY�ƹ�k:�X�!�e����{�6�<��A�ň s���S��zk;���������q;U;��[�Sbw�UAv%s��dE����X��]Ktҝ�Ⴏq)�0gG��/-�n��Xzc�/�ͮ�c9�o/�"�0D�H��M��.�%c�Z7�JG��\�uF�,';���Z���t��v���.�Y�j�MT�'�8�ʹ���B���`��u�W[����[w�F���:�gIښ��!t͕���NͶE�;���vMi�B�"���uӤ�v���{�����vP�NH!Fl��Zf�1�`H^�����g.�d����r�u��I!\cz����J����mg-�y�iGÞ#k���=�ӝC1e%kR�t&�sQ��v���k�ei��=��/f�9��w��S٢r��X��;�����t&]������[�@�L�W��I<�i�����v�9�l�:SVSh�������<ι3{��T�o�X\i\b^�� ���Zf5��P�m֋�3�N��*��1�H�:�e3`F>Pi/qT=֨a�3h���9���o6R��yC��׃Y9�)����T����>�_.9��g��A5k���������3V���eҭa���EN3�.�Ȕ��q�����ReN᷒nqʜ譭a;f������]ةm���a<�7�t��*�+P�B!P�-�^(��i	�|3"�Yd��:d���Y�9�٨J3��#F�J�պ�*�	v�F`���m�gp��,�O8�FpQ��=P������}�h��F�ݭ�Z�4R�47�uR� i�,ڎ�R���>���5�w��I�s�E����՘���FtL������.u�Ѫ��ʳ���Sm��5�����=�%�\�ؖ��^H\r��۝�	�-��TA"��V�Am,�24�0�{��--Q��FbUxi����d�gk��/m�N��=1�9�Ab�2�Dqa��̶��GJ;Z�j��c�>�����=7����gVw��H�żDI�:Ɔ����l�`�JY�o-\�ʹs3M�=oK�>�hD
�0DX�e��w�,,���J��=|m��u�t�Ӱ�Pݽ� �!՜j[�9�ZF�Z�JI��|�M�f��Q�}Z���v��5�Z@����,퉵�E���z՞nvF6Еp(Y�4��);wqλҴ�:��i���/-�WY�qֱu
U��so���\�[z�We�u�ޫaAB���]NW7�b��.n�����[�	w'�u��������y�ZoG0r�v�s-9G+1f'���ov0���Cl3m9��e)�n�|�Q�]�+�=���࢚@G�Z���Z�q���lgc�:��X��K�l�y[��讘U�]��%����d�'n��
����3;�8����hOnm�h���֥�ovT/�E�Y�q��%rK*M��r���JQ�����7Z6Ve�r=���Q���'u��:�b9(�PhL���m�v��w\������s��C�i?kU���z��ۺFC��;�=��f�y�¡lo(��U4��m��n�ή�o��0^������Dg�o�8�[[-�J�;�L,Y�t�q"���clH��et���9��c�r�>�";�;,P4���Gp��a�'2��K��<o�;��������]wj�7��1P�ؖX�JQ:ܷ�vS��`���s�, �m���<����h��Ƿ���M� �����,r\f���O���e�w�X3:�K����cn�4�꼥V$WO/������4q��z�捗��o���F�󤊣���^�تV_����Y��խ�0�,p�.와)�����/�s��Ѯp�:u�hcd��L�u\��\].ָf#�dZ�*^�BiK�)(��)vv�C����w3�{QKEӬ�I�
̴%&K��+����ۦ��������,NF
�0ձ�h�r�C{op���9�)�`=X�� ��B��;��ԩ�c:��j�7��SqW^�j��Lúd����ٳ*��d�{z�ud�;��lLw��!�V���\{.��gv�*��t��0�K��J��e�I��M�lt~Ӊ�k�n�����ǽ&tb�&�w3g�]��e��ș��.Kay>��h����� s}�\Y�Kaa����w���&Ƌ\iP�}urr� p��[LDڽ���k���պ�7�)"��{)�K���pk�����U�۾�3�it\HLNu��k=K;�;�yn�L呝����\�U�{/���3��gBz�����+x�C�"g�+U�T,Ыc.%���P���� ��:N�lN��s:���;�M0��_>{���M��m���`�1������������𻙷e��EY�)f�̵�sD\�˥��<�} on�W;
<�i��T���s{��iQkr������t�J���
�ně35*�����.9��T�s��g�����W@`%p�[�����H�86�I�k)�2^���
u��2�w��5U��x4��bK]�7/z��čM��kT+>lXduf��8�ݗI6��c�Eӛ���'�	g��[�v��H\٪�)m<s�}�q�'�M�al�SiM�4d��cNV�1��*�Ԟp�s�btO��w��gb��N�k9��;�;Z�#8e�m�%��,h ӷ�;bue�B���⵪zЙ՗O`�к�K2!����5]rN�ǀ�Y�))Z���![)h��X��{)Cɞ�Y�q��C�D�u@ww�M(���|u\\��5�g�5�i��l���c��=�.��W0)N�V��v��xw�S�po��l�V���V�s��<�p͸*P�wQ���zU:f�v��#��N/�ۃ$7�Fr�/�)���0U������������u]bԗJ�ZǛ���.ޝ�v��{�b��D�`{�9���
=I�q�
����xn��:����w�g��M�VhZ��(+��JbZ�I���7�oJ�*V0+vv^�sQ>Ƃ��r�p[�3>���Z胏�V��w�^�KY�x���ŉ�+��=H�˸��� ي�^&�u�n����Ż�!������8��.��� ޔT�CJ�+V7\�.{q��ږ-7W�q���L]�2�(^�3��ae�qwb㤛���n �me8W4YXzR���u�p֐7sc���/�-�^
VaF�W�z/yX؀�S�8I�S9��-kL�eh�t5wl��T�.:�[1�9p�@���H�gk�����b�� �c2�����V��o
$�XU��N3r�]YT��Bf,ү��mu�2���H��/*����ѭ�.�¢\�h;n�0T����wVA�%�2c宎9�c2���c�B��k���M�t�ٯQ�&L�>�G��R��Q|����Su|Iݲ�u�(ѾV��>F������1�-<��w���lũ�[MD��X�X��o#P)PՉ�A�3���#��ЭU��P��7��ʒ��U��fki�YV4S��yW�g�z5+���*��%�fq vHX�|.��H��yW���X�gV=�N>
��N�h:�wM7oN�㸸8"�U��)�u.�9���C�ϰp���1Yޢ�p��M^��u,��i�Y�_�7㕖�0�u
��и�����V�Q�H�,ih(_|�C'\�ݾ�([*�UÖ&d�tS�B� ť�lANmY��^q�j���f�&�ͧ�-t��پ�k`�S��-��q-,�S�+�W��W#r�K�1#@�Ǯp�m%W�����Ź�ՠ�LP)Siu�Y�&A���DM�5@�e,N��K���{�h���֛�/9����M�u�.d�w. ��5י���-)��ȭ�&hTŗ]�غ:Y�S���u����N�ܝz�[*��m��7]�r�*U�vb���:wWYmNŦ��r^�	&_]�l��3s����/V։�
�JN��V�j���Wh��d��/zūC�o:��Zv�	�pԕF��#Si�� ������"o�\�0�v/�ɷ���Y�Gf㨳�W]|;)p�T�،�D���r�޽.��)a��N�tƼ�k~Q�*�jZ�5V�w�p6�toS�r�(�L)"1�z��/]ξ)��-t҃�Ŵ(K�7Z}�md����V}{���mĤst[�#�.7�@Gs9�R�>�*%�A��Ƿ-�z����qc�ff= ���%j�X��ѣ�N��m��rA��f�v�r����3*�8�����4D��L*�Nΰ���:�o���֫�h�-��ҥ�
�SM���e#]�X?�R��	��b��q���z)��C{�j�����8Q��5v���xS�Y��_h������������wV�խ�@4I���@+U���`���q-���C�ϟ9Ƭ��G<s��˞�\r6����Y����Bj�w��G��Z���l���u]EWy[@�,h\�l��Q�7Ճ.�[��i)293-���:�ؾ��8��kr�U�ޡ//��k�Pڣ���u0AoW2E���|�4��0����z�9hL�X�U�]s�6�ٵ�0�v݇��5�;zWV��m[�]�*-�˻8 t��h�Jo�΀��z�^%�6�K+f�{MQttn�V�V��oV�*�j����>�J�ui���n��U4�<E�wc�.��	�Ӡn��TW��r��V��\�Hq���S8����b&��]6\lp]u��:��2�F\��ۥ�����n�nA��Y!�vm�2[tXUO��k:~M����#o�Q�x/q�/IXD����w��
�:W^0���l��w˗]�,2�:t�j��I�{+V���!�`u�, i���;����{�9R3�uV��X�5�O%h�91���l	Ɔ���VI�h����trY�t���`�]�:�;�}�͆��}֝8'vZ�:U��B��K��Qo����J2fu�:��6WP&�h�RUr:�j�j�"�?eҽR���e�ݒ6>e���H�c�G(h���;N��Zۺ���S�(������u�K,Qߡq�j��Z5��lgmڸA|�k7.�G6�zR��9}��܇������t���Q��f�G�VEGd������n�/k;���h;u��TO[g.�V̦�]hBe���*L��Nbi����R��bë��Ć�ȱ����F�����;ux*�<��S�M�Q*��T�z+1boI@Kz�Wu�l���C2�L�ike�{�ًTq4�M�Mj���}�ye]>�WV��}��*8mrD�|��I�nD�^@��԰}zh15:��wR��rV�Zjc�in��t�Ŭ�#P�'v-��m��b��+uh��D�;Q������#yY��ę�e��ǒV4�!����/�]�`J�."�D��9=m�V�$�ku�}t�A�&�����Z�fķ��_v3�֜rc��Y�����@���YIkuۗ&��v4V�Z8���mTui>�9z��8z��%<��!IaVF��\�]��+ɫQ�zyZ�еr�Gf^7�P�@�Wn���Y��N�]e]�G�R�@�®�
0[�v���6s�C�J���ai���-T���ti���ّ���5�m��:��1iV�`0�owT�+qލ��*�5���x����>�\�
��7/{�hnTq��I���ESm	ۃ�l�@T6�+��H|;(�V�S��X.��YDàv��=�;��ÈY���S���j�`��w17c%39����Zn���V�W�j�Ц[��vڜ'j���9�`V�f�P6��63�ٟ+���z���]B��Ȋ��E���`��/2L$������6�ZoZ�F(���&欺�$pS�W�j�b>�T`̙c+X��kV�1&�>�B��u�m��*HOƏݺj]2�G��-�,�vv��,��5Q�h�=Y���DvQ}	���Ry�Y�.+���^S��������'9�j��w�A*��.�S+V�M�w������Wb�J��]����k���]GI��LT��c/��\}�P�cbӃr�k�RmWf7΍�֞�9�"�5d���kc�ymk	_0Fo+m<��b������p�U�����ҙ��z����ع���#6B�
7c�c�w��� _j�y�PJ�1n
<v�]}�\KCfv���o�%ꙇuk����4�Y��>�&�:��1�_p�z����I|�٨�EN�7��ዢ+X��]S>��\��Y�bG�/.����G���W%YU���Zoa�4Gr&��u�E���x��/yӰ��J��o8�6�D���3�T���o�6�1.r�Xхմ-}�7`<���ڨ��{)g���y	���΂s4��Ǻ�CX����u��z����G�
���4�G�t��k�ˋ��(G�7G_*�&cBb�����r���r����/5�W+෹PvA����V(�+Պ.��SD��`Tb:<�Aoo#F31��F�R	.�8��̤��I�9�ʼd����v3Ъ<� �#ΠXΡ�E=a�,c���Yq�xIH
뽭!nf�T����κ�;b����f�y$��b��t��X��ۥ�]Z'{�ag�;�������҆I��V,Wn�[�R���u�LgF��:XZ�j�<;\���zF@U��������a��V����
���잎�h�/�*T��`�D�W1_V'Ώ%о7��N� ����ǜ����
�e=�b�-(B�;f�*gq'�]�g�S�x�N��}u�G`w�Wܦ��u�-���Ƽ<���/0JU�`�0��i}���4�Q.�_Z�:�\'-�ި\���_M��W N2���dU���4&�1As�����Ƕ`nSY���et �F�p�̋`8Z�J�`�C���in��tfW@Dv�\,	�Uwn�Q�7%�=��{7�T�ƤV.�]#�ko�sR�(�λ�ܕ�^TRC�l���v�������X�k��d�pd�g+z�Ѽ������ Fs�oe�9�On�k\ϻ�Ԟ�.�����N�ZU��W�}W�r�/{\��gWn�w�A35R�{z�ʓ��&�WM�h	uw���ÿui:�#��8��}G��溿�ں�
w���e�ݒ�e��vT��ۛ�҄e:f�1K��;;�f;{�d�cm�	$$ǻi>�P���T�M�H�`T]'��9����Tj�u�΄�TX���l_r]Қ,`�
�:]�q��M�a4er��yL�Rj��D�Myu�v��]�������ˣC����[|�;C.l�����ejÉ˒�������*����V�;&�r��{]���cU�м6Ue̼ɒ��%.��˛��vt��r��v����8`�a4�Q��_.l$H'lG��$*�2]�OR�t�+��7�N�lu�й�ہ��(P�0���Vǋe�Ŕ(BsU�.�N��̬yC�I ����y-�����ɨ�5� ��/�p]�S�u���:�e����n���)���3��h�Kz�XӏOp��R�]��)*٦wm�3����q��+5u��e�lŲ�e�;n�m.�z#��V�qt+5&ە�.q��pi�y���|�VnJ������Eǯ$!��Ǒ��k����p�G����i|��<2ݍ��u��]^At֍�;�n�Ccj�,C'�U��|�(���7+��Yc5'�0�hi�)̨���Ȯ�_@���t)�q���	ɷI�x�����k�f]��59Z!/fq]*.��Nܩ�T�%�;�����8{v�RÊՃP]�	�Ӷ���f�[��Z�Vv���w{o�.!CZ_6D��b\�7�V�����Т]X�+�[[Cq����F.�X���S+F�	����Yj�Xls�E7�S;��,�Fʆ�Y�W�y�.�ҪO�g
�k�w��#`R�TBc�V	:��m����=��a
��qQ�jz��Z1A�/�xAJ������Z�=�����}�jMЮycNn�']0%Z�Uݺ>��3X��4B�`8��hM��3���+[�̫��4�
4�aG� �A��i�t�v!�3�t��[�9�;k�[�&��Q�s~�W�ٛ�����K�k.�M���,�#x5nY�ѰpL�û�tW�28r�y�y�ӖtB���Շ���b��u�*�K�a�`|.�'$I���/]�F�?�́��:�h�a��QCDZ#n����+�.����G����nWT޻+���Es;�6*��0���n�|�b��aU�U��R�w|�
�-��Y:+�HkR���;�ͤh��};'$���wwU���Hbx����b�e��ٙ���9�P�=�t��k�y!X/CYٓ��}of7�i������A�k�"L�Á�����q�>,��#@_r�{ݶ�vʷ z���D�U�g)�HiT�e�}yn��׍Q�՗��a�k�ܩM�ʮR���O�&��8u^wR���zgS����"\;�Ӂ�ٹjNv���(��72�s��n��:4�7'S�i�glw�ϴ�P�q�R<���R0&%*WVF.����u9��[�q�=B�e�b�lw-P�Sī��G$��t��[L�]���u�b�j�Ń�R�"�q��{w%�ھt����ֿ��b��%D��/r����z�0��Z�u�z�
k}cj�d���v�L_h[�b�ɢ^U�]�I�[�F
S+��u���N�[-�e*x�g�sH�]b��#u�&N��).�X����f��k\t1�N��vp�m�ܡ��xW"y��2���=�`Μ%��8oJ�T�.���wK{���\�귮!Ժ���,۩Y\�����1	Bj��u��γJ;	4�9��0޺��m������Li�C6��m�������{�IN���@�;>�xg�
��:j���.=�.��t�_V�qH�п�w<ճ��$G�Z��+�������;7f�kc	4��;��ޮ̙xr�l�2�c��I,�y
7|�)�,�Qˊk���Ǒ,��2����JU��/z�����Ѽ9�y����j�'��%o&����8
�v�`��/��c�sE�R��g`XskTIY�+78�-�!��<R-R3�����,�GjvH�<�Yw�gq7jr�Y"Ř����tS���N��e�W+��E*4B��!c�:C4��j�\�NwF�nI
���S}���pG��]��|ͧV����w���W�U}_}���ސ�1��H��3H�޴Vr��[fH]w09�l�i�N�,חP��SvRk��5�1P�H��H��%IY�w���f�	k�젠S5�9�'7�U�bEN�6�t3w)��R�)�Z�Y��y�\�ڼ����ѩ9�_fjI�N�k+����W.{��ݫ���iv���R�`*`<��㜗�L_l�ra|�q��z��C]��ڼ�8�EB��s��u]8Yr���u�o95�ݷǥb�Z���l�u�9��ƫcM�!Q�Δ �睤iy��-vv��ev;���Ƶ�X�ҡ�B�׻�1�2v���8���V��ί������T�&
�od�Fʻ��o�Wr������د�z�rqK���qB��;�qgl뻺��L��i|z4o�[r������B�i��F��
/�J^r��;������n�uA�U�Lu�0 *�{C��8$�X�-�<o���S �wƻ�7�͖7\�A���\����yMT�&bhs�i��|�a�h!j�t"��s�ڕ�ۻ �8�9ˤuY�" pb�m�cK�Q�6�j��pZ=�uA|0�q��`(�S����4�&l�o�XS�r�7L��û��^#t��e�[��*9	K�=�Is��,�2�X�ty�;:b��j��e��yӵ���W˲�],��/�y8ui7ֆ�.���(�dtC[r�+��@�a��݊�.���W�j��j�+@�@i	UT��v�w�^c.�Ir��T͖����)��DRy'��su�y����3tuY{���AD��*E��Q����ܼ=O!#@���*�:��E)#H�� �w\��Me�/�1��Y�dn��En�O]�-n�n�T��'q �r�s�,Aչ!���ibl�;��Q�I�1�6�i9���L��au�P�"䧝�wUh9�y���u�������V�W=�r=iVu''f�"��r#�Y�G�l�AE;��Ur�C$��N�DTE�2Z��xeI�:9ⴏR�d�#�.s�V9��U,�����*�ԉ�uHse�U��j���\<tJs(�\�J"���Yr���f�g"�ᜮ^�WuDC�Nqa���:e�Q#�(P�� UO�ED�i�NT���K@���Ax��[B;��woy]��u\Q�\�]��@ �bøC�;�z	zjv;�)�_|rLs�r�Ѻ������C9��i���)�+��^��)B��@����';k*�<�fw@�˸Fi"�Ѯ���c������^L�<B��S����'TVs9�A#���g�OR:\ktG"m��a$�D���W�!�\_vE~*�p���QM��rH�=�������U�u���j����B]�7AV�_���fZ��ҟ��XSwgW5�X���^� %+x��j8G20�cʱ7��b��ב��
���]���J��ר�z$�`h�,\�Zu�!��Dܑo��]Z���m����U���)�;���g�s��!�_�w<���X�"�m�(�ku<���'L�Z;������;����u�Cһ�^q�~����p@�%�g�gG���:�j�}>���ki'o�[�V#�3���-z��1B�Σ��9cF�<s�	��ٔ^�@^J�Db�L�Ԓ�JR����y�q����le���R;nc�*��U�Zik�Ip���T���u+��7��r�z)u/>�׽l>���
�)��gP�V��̈́�%���j�+�A��T�����7lE��3�N�w]K���fhK��Wj�ʇ�}7;��ٜ�e�ɼxr8�r֞���$�ڀÜ�����ʔvGV��R��UQZw�i|l6G�p��7%c���a�Q*���KaFR�ٮ��5���ǀ�l!�c_>ۺʭ�n�ڿ��ӹ`��;ydf����uɛ��Ϳ_؋�Huʦ��twϬ��خZ��F*u�S�@����X���Ȫ�����`���2�B� �
�1	��hTA[O�����)4�&�uQ��a�����	_ke��L��{��@��B�.Z���h�F�ΨK�gcA;���)��n��ϓ�5���m�џ�^�C��$�����/ƀҾ*��Q�<��F���w~���F���Ⲝ�\�1=V:��trR�Ll'?>6�(@YD��(��>F�y�I��%�
�	�J���ֺ����$sr��C�cx��:�X���v;�f��~g�+X�^�^D�*�tv�}�}nM��NI�Ŏ�M���,�a7<��� \Xc���7��(%6�n�kIǒoy���2�ĀƁ�/c�Xq����+�S=9����d�s]pl�2e<8=YX�%:�����':-sRh�Sęl���v�ӻ�G|�aڷ��$���ɼe�}�c�o7�֑k�{x�c5��Di7Z�Dڸ�Z˄��h�+��-�VD�NJ泘�o7xJ��Y��zB�|;��n����
��Pu%����~��+8��/.|�cQR�I�ؖv������a�F����+\.U����{��j��gy��N꘼t�s���fZ�go4��{qW�O��n&���舻2�+4tzg�7���Y7�M\�q��n$��:���W�ۦ��s,��}>���t�PV�t�@rS�r��d�m�]wv���ل(8[TS����:�(+����̂��d�*�̏�R�R��i��zn�N�sF����734���ɸ�*�w	�-�0^8��	����)�X�ge�=���p��Ʉ��RF�D� ����<���C�*7\<��8<�,fL����L���l�2���;��B�����!�s��H�5����#U�F��|`byy:IY���b�noo<ly�"���`V��䨍t�F�ʹ�T�1b�6�y�|gV=i����%΢n_Z�qƈ�P���Y�0����a��&9��?y���_5*r�$����������{����[��p�rb;Sː)K'������k9��|+qQ�l|+jVl_E1�xC]D��Z�X�Rڒ*�XN˹�n��8m�ԩ�ΗY���E@r�`Põ�����:��IT�d�}X,���+u�
��[��弥�wg��c��x�=6�l�w�:[��]�
����~�[p��H�w���]	� l#�{�uF��q�ʩ፬��D�.&[.�������?[;'~̔!��+cE�ݚb��R�Z��5
rM(Y�E!U�tj�C{P��� N�<b�cp���B�ͧ��z���f5�[�,��s���H��}�¾O.�ɳ��L!�Ixu��xG�A�Q[�*�p��gE�h8�x����IVw�5^����Ok���F����Ɍ�ȉ�C/&�hQ��A��r��Y�����4<9�F�j���?S����9����ȑb���3D�!�nsJ7f~8����S��5�Ma�d�!XPƧ�;#U1 [r��E)����Ϛ�(��@R�ų#�y����ԍA\үi�G���q�m����(F�-�k��0�]:c�{f�xRt�ҳ�L?=N��0N�c���.u���"��&qSW��ea,c��4���Jj�U>�����φ鯆��Ed�@-e`�*����b*,�(! ���R��p��8����{<:�V�Wbŧɹ����[]�V8(n�3l
�]RVΕ��kP�Ȳ��	d�u����J���9IO�p�o;�$_uћ�D֯�G�g�T-rIb$JMMD�Y��혳��y�j�}��ۑ���S���Wq�]��%�t�b�ns|�8��\��^���;B:N�ώIG�#�D�u#J� f��!�e�����=��z�+���~I�F2
�9��)�!l@�Rx����3��v��B���fg17ڑp�,��.�S��9�������G;˸��Q<��o�+/gS�R��]��bauE�&&���qH�w�*��!�8[�͆'X�"�P�z�ZVZ�Jo�$1�8@��d���&&�VѸ�c� *��3c~o�٠�l]t��'V�mp��WVsٌ *��Y�:�"(#^����9l�s�y������qT��ג`�&�>HwV[��͛��f��]�u�K���<+��c��������X:9ԍ�V�^��4̸��:���\G9���uGJyU�=����f�J�rPo��w�$��Tw^ʮjaY�38Ζ�T u��:)mGl�;�42��:c�=�,z��J8w����y]v�.j�a��j���xFg#9P���`T-�"ὤ _:���#gLJ��wMoG6�w���`+B��i�!�|�7|
��V��9��J{�$_
�`�We�Ɇ1��}�f��\OUv	�d�:;;�����ޚ`�R���LT��_|�K=v�V����*)Kc�{p$��s|�W*�Z�q�t��%����!ݙ�ڪ'*�u�nҐ5du:?U�H��3� �.�z��k�Y7sؚ�Z�t���~��B�r��S:<��O�����lN
�;r�25��û����;��/)�ȽS-ȉb3KE�h���d	J��H�P�%`��S{O:�q��������z���XT2�\s��Q���V&��ҭ ��� +�.���=V�i�Tֻ�W%�n��q����-;�2���c��8��#nJ��w�=�1V�2����7�j]��ף@�5��enF�&"��.7�y�q��w�)Өc�;�
5T���94��BґϜ|>�.�����WQ��Ζ�c����p:�-\p"�:�9	� D<��,�Z��K&�0���+fEt���!��!#\d�����v����O��se,BN���7}}��)G����w�v:�"%��p�L����K�Y�3�db<�e�Y�Ԕ���7[����;�}_s�.�"����dS03O\M�QnH\���8��}LM��e�R����1<� �z����H�o�Me�gP�v����T�H{RMj#������V���3��F����g9u���ge�A��J}a�͂��x�
�ub��΀�`��r�f���eX�sz���3u^$[o9㫣Ҋ����7S�=Jp1 �Û� ���b�=�.���~̹\u�SmáQiK50���k�l�@��x"z��"��Y���ŋi�y8���{Nzm ���:1oBud�a��ԑ�~q�$-�t#�cj0���*�qBj���ۈ�����
�<=���� �Ks�+��`��2�l�ݽ�����]b���{��?``���ǵ��(ڏ;�d���@�x$��-�탟��1��%��I��Y��ă� ,=�٠8?�Z�r�䭟Z�E>ƪ���ed�
�%��z{�d�<��ْl��	���Y��JyX��؈�1r�C�tz�k
�}�*�T`x�ZO��K�o����[*��N�+6{�ٌ�_Bx��q��<�6i��J^��۫���y�8S���jr6�<ꨠ�d�?Zn�;���n񌯛�,����㛞�Z��o�w�����N��'M��ǉ�0���� ��N�b�����ľ1p���꼬�
�4����qZvgY@��_GHu4LF� R�'��̭و��I��Ȁ�Bl�[�9�n��u�o�5^\R�L�������xW�aoj�vx�l��X�7��\f�KT�V�__��x	��m�5.x�0Onkי�e�ð�T遻�0�ӛݭ�t2ƕBvpo^Z�P�v��ׂ�`j�p���\s���1��=�0ҳ����(8�2�\;��������s��_>5|�^暈�}Mi/o/��3��Z�g>dh��8*-�\�L��n&

�����|�\>k)���q#���I�������t�,��99:U�ː�RQ;cGT��=�0�觻٤��bxQ-^�!� ��1aڝ��,*s�)T���GL'w R�J&��"��[�s�����Ҵ�u�W�<LS�ʘ��
��.��sL�9T�015��LΥ���5Ag�����n��N��m����B�T�
��Lr2!��𮗬���]6��^��<0P�GM?��(�7Ħ�������.����0K�uϰ{ס7)u?&�o���%�����eR��z����m7��0�\�Ęb��a���kŌ7fU;W��n���p�w+��z��ʶ7����J���-mT�!�7�S�O:��W�:/X}����a��N�)�],+��P�U��:'�<���@1[�@�ͮ��/�wZG��nP�%�����j.�:���v�f6�~7�f�it�G��nI��,	J��q�6 �$���K���u�[lNj���`A@�E��8t#��U���h�����s�ݞ��ն����k�Nτ��C��W���;#T���MϨ��������m(��7��4��W4z��R���F�]મh�Ә�y|�?s�)?�k��[�ᙔ��h�BVgԯ�M��Y���r����)-.��ܢQ��|�U�zcu�3�~���@���%7ۼ�f����J1ٮ��{��9DB��Z��3�S<ϕxTǽ\�E�.@��nf'Wdaʬ��ejN��鳃D!�o粄Tnؼ���|�"�S����ҕ����UW�4�K��Ĩ�q��I�F4&p>1���
�ʓ����^1<����B{��.	|^*a���T¼j�,�����qS���w�M����ze���3�xҎq�Mp���4;8zR1��w�'m�6TЊe�M_[�ss�M��K�I˧t�@y�s,-6����V��0��|F��I��c-	���vj����1�t�kW<=��p��� :�<6Bd���?!��Gm�x5��<E���7Λe�]�k(��gQ�����u��Sp��`�F�#�92�Eԉ5�r�v:0V^M`��D0����k�)\VS�Ħ��7+��]48�r�����
���$;,XW(�^����Zڻ��I�kf��An�44���W;��*u�MEG+:�U���k1mu)۶V�/y�=�r��k���N�!X$gOe�B�W�4����Ӓ��:��2-�-��Wh�t��β���ϯ�s���On���p��`�QW���N��'�-�MoWon���0!^���\�p
����sڎ��avdOC]gLp���;���9�ĘC+�ʄ+�/J0N<�zX�O����� \s�������'�����+�p�h<���T6+�T��eP\@���=��<ޝ�}g/캩叵������o8Se�����o�o�@���δ�����c/������8{��m�0��oz��bW�}1����4�.X����4[��o�@ ���\���6i��=ev��;�a��ƣn�Xy ��o�岑�s+௦2�U@G�$	�t�RKx��`ܭd9��哠7+T��2x1�H{m��>
[82Ξ㌽5*��i�#^�NԴ"oz鬽!֫��#�*�&�j,�+sU��h�ͪ�>j��v������M��QE<�U���̇Zol䭳t3��pR�D[�Y�]�'�9���[�X�����4�̩�[ܥ�����j�`��%�d��t�8��������Ѥ%A��e��.��T���t+4�bTj>:`ק��u6�;�%LO�d�TB3bw.�޴1��Z*r�`���%�7],Me[�����6>�d�NEP�f�&�nt�_u6��*.��fl�b .;��Q{*q�������_*��X%��lrh}gW`�j�9���Be�K�-Q㈛<��ˮ��o�'� ��0�e5��h��yl�g��Z���-3pĶ�4�V3~���:�y��M��dZ������\����s/d�2��b53���ՔѺ�n������#>`���v+��뵈�`�����a'����ѵ��N�_Hn��Uԭ��;��]3�AY����sfbe��e:�p��Z���|�g#uj��
���q�"tm̭I�Y���ݜ)t΋A�[�fY`R�h���޳M>�M�:�؝]Л���Z�0]v`�k�YJ�VζL%TB�����!�Y{��,�k�l���Wkѵ� ���E��6p�}N��GY�m7GZ�����0
9.j��ʚEy_SC|��=��"S�t���d����8��j��4����UE��]]d��,�]��]�yI�j���Ιٔ%��,��V�*3ͻ���f���'X��'��A��;�j�W�$�Ɋ�B��n��R��[0kݙ�w��Ϗ���J�{^���=�y�~��Ev!�(��!���v0�`Z0]um�����ᣳ�>ű�wA�6��H�[����l��E��BRV,w�wucmn�5U�KiK�-�*� �*��v�ʕ%]үiӬ�J��]	Ǐ������ϱ���ft��=#�$��M�a�#(��d��×H;J�y���Gi�( 0S����jH&�̥���](�\N��Y[��j�G^�Pոrh[�m�3ff*,�w�S%7dM��4Z��x�u�cnJ�M�{]}d�t%���m]�@ȟvg7Nr�}D��@�6e_.ε{��#� ���&�euN�N
[o
�r�0�Xyֺcm�}�����,� 5tM�����{��t�%<���&��S������J<�Lc���^���z��$q�W]|n[�=utj�le�OPz�:�Q��ԄQ7VE%ن`�u���y��'_����v.0gϋC$5�`�z'�u6+������]զ+h�]2'��s%ƨ�gJ��K�g��J[�y�E�������W�;]rF>{r.olvhq�A>\�(�]�&�#����v\[o�/�=��8Һ���i|�T��yt����\���y��X��9׭k��V���8RA�ǀ����Utt)8�pt�Q#:}ת���Ɍ�
�v�e����P�H}i�ڤ/�hVn}Z�η���Y���N�|���s������>x��IT�F�'u���NZ�.�
��z���l�M��]	"�9�#��*'SV���ԶE9%R�*&QUh�sGVEܗR1
�(ʺN�y�N%EED�\��3�r�����.*�d�Ue�u,J�2�dr�u�+�r�J�W]�%��B�����J�\ʫ�]U:�"*�C��9�N`r���D�HFe˕D\��*(���E�Q�r�dr:�ʊ�)�p�p�92�Us�#$(�2t�9��IS��f�]R(4H*քtd�*"�dR��2U	���8��L((��ug��������"̈���J��Z	��(��.Q�\VQ���b:��z��I2(�b�wCvP���%A��\��p�uێ�]W]e��BH���%�j�Ґ�K����,Ӭ��fM���PM�r�Kuȍ����@WZ�ڂ���v�JwD�^p�F�vR�R���Xq���<��Ww7������>&8���<q���&O�&��w;������!�>����<'&���ߐ�P��!F�C�?!�����0���>���w��!n�G�}��c�DM�[�*�o����������'*o�����_�;�ü;N����}y�]�=j�&��S~O'B�7������.	�C��'���97������?���f�} x|C9�s�U�ZY��Y���{�*�V���5_�b�*��G�_!�޷��<��BN~&���zM�	Ӵ��~�	�!8��9����<!��x���?�|�eۓ}B�i>8���Ϩ�\~�G�4}�1�8~�c�<�����?�|y7����;�x�;�o��~���A�0�����������Ϗ>�?'!���a��m�<�N����7�ӎC�����t����	������=x8>��D1@\���R�9/�:�����_�����&���)����p>?���_�P������O���o4raw�O�x��7>��0����0"o��s����xg������]�99��!1��F����%>ُxM�j��m�"�>�!��b>�8D{On���@���׎ɧ�<;ry��~C��Mu!���&���v�~��������ˉ��L.���m�7���7 }}b5����\ۍ>"��٥���r_���}�}TG�?X�"����Ӑ��7;���'A�0�o��������&��{���[r}�p~O)�!'>�v�}Bq8��߾<?�DxD���c�,��B"Cxs_��˵�v��
��DAG��v�@X�I����N�����t�s��!�}q��oi���ǔ�墳���c��<�w����yM������q�"DB"2;�DxA|G�A7gXJf}�~�]~��>���"#�n:����F>���ݽ&O���~p&�i'���Ǎ�w�iǓ��	���Wo'G&���v�����xC�i���x��)���Xj��_xX�������
��{/��y�^@����z9:�"�D������N�㓝��]������}�ޓ
��Ğ~~��>!�0��~���%w�i��������=�w������O'�nM�	ߒ���[ǿ���`��|\�f@Zk��fC��b�-��9�U�b���j�.�.��&�IZʛ`�_�h���/g���=�p��G;瓥�m���Z3���ɭWqظ��k2���jr���t��������F)!�h� r�WrQĕ��,��"DE��q��<(G�G,�coI�:Wz���<&��w߾������^�������9�z�����|w!���?!�0�|?�v��'�9��R�����@����G�I�w�����ǯ���ɧ�~�`��P�͏���<lro_-�����;�7��Í�Q���6�>}�}C��{w�������������`���M�t�y�w�{��M���~�w;��_�ݲ���	e���9��y�o(Rv������7?�r���rS_ly���!�0�S�{��>_����=%�������w����
�+��pB��6.��1"3\�߶��9�#�1�ލ��F>�"0G�i���q�0���}�O	��]ɤ$�&�'�Ļ��	8�S�]��'!�4���}����粘\|qx<��~C=~���~����b���^�U6�r�iǽ�����q�|�'�>&������򛐐������y1�7�'z�]����9��������G;봛�|�?!�0����������<���G�����E=������ǉ��]�����yL(y�|o�����;o��������� I�7�$����]�&���=lxIM�<Q�'������e7 }I��OG� }C��sěd]Fo-���A�巷s��Joh_m���^���<������?'��]����|�8?u��&���>��<<��������~1��N�w��;�����nB�8��Fz>>�3�J�wq9�ߪr�9�����a}'���ǟ�97 x?8����w�i���c�S����}��Пo�i�xF>�#�#��͆>�<b�} i~<��>���w�=�#r�o�������� ��)ۭW}7Z��unޥK����NC���''�x��;��]��zC�aq��w�x������~C�*�	�y��x������>�±�7�$=��qy�I�!?���oo�	zJ���<������ey�L⽽�����G�_A��M�_!TE}@:Ï�Ï���x���'8�����yL.���z=���O�90��Տ����xC�{�c��$�����H�M������������>s������쨧�0;_��ϓuKw��hD�l���j��q�a��n麗B:��q��9+psGbj�����{��Sl����`�ڕ#M4����q=Ǥ��$r���ރ��O3p�L��k'`X%�+�5�3$=��o�w.���ވԪ"��G�CG���Ĉ���i��o�v��G�<u��r��&���m�=x}8$>8��z��'��ﯷτ߿��o��;xWo�&�![�=�w®e�9^��#f��]�8�����>���ǔ�8��G�xw��n8���y�L*��׃��^M�I�����1'�=��z�r.�ޜy�7�$������݁M�	��>���>�"!��������w:��?]�}����������_�~@r�������N��2o�v��}C���'}��9ӿ���y���&C���򜇴9����!ʇ�ז��"!��S9���޸5�~+��}�7�$>'�;�8�]���ߝ�7�>�8�����|!���7�~v�}}w��M�	P>��7���������<!���<�~��|OI������nBDp��@��Ĳ��n*uR���<�i����ǋn�Aw����XP?$��x���ۓ~B}c�xW��'���	��}�������{C�i��}�/�iN������<����W�G�_m���}|Z�q�?��gyӯܕ���0}DBF���b$G�`�y7ϐs��ŎWoI&�yܘ~�~N�.9�N��<8��~�����®�������P����>W}�?1��>m��՗w�yo}~��bOH����]����o�I��׏��\
oHO�޻i<?�	��7�v��<;y<[������=o�®N� �;˾�L���(|O�s����戴��xDI�ۂI3�z�e����~|�����&O��9>!�M�������9]�~q��H&��돎�S}BC�����I�\
o�s�k���xC�4������s��B"��1� #�� ��#�Fُ,*�<�5�G�#�H�4}�q�DB#�������|OI�ߓ�����@�{���M�����}��9�H.�~����P?$��'?�7��G:v�DA'�b"��G�G#�.i8S�|���*�fj{�#�C���$h�⋤߽^}B�c�W׿����<�����Cü�~�����}NL>�}��_)����޿�	]���ǟ��"�} 1��nb�C>��P�����_�	B�=W���nw94wah������z��Y����C�h�(E�����mfa���+�U�VۨL&	���+�73�_j1����oVZ��:����!�$�󖫕6c�/7�a�Z=3���g5�Vhk������ٜx�	R���Gl�������Z��-����
��x<���o(r�����۾A�7>���xE��;������7�$������7�p)��{�O�o������~M����cÏG��1�����/(��]��Ui�~�.���]�We���;þ;L�um�|O�s�'�Ŕ�]�ߓ��S��&��?!�u�۟�}q��i�/�=��������>�ro�O���~b>�$}By�۫���:&�3�ڡ+������]}M���ސ�M:q����&xv����w�iP��97��Nq�=x��pH}C�;����xL.�����ސ��P�J��=����s#�����'�5�S�-��[y�w��D}�",Az;�|�F����#�3��'���O���P�@��w������M!����󴋤<n�����ĞW���{=G��z1%p�U�1_h�)�3���u�{-+���Y;C�+�P�D}�D}�b'��} ��G��vP�_N?�����O.9����˴�ߟ�������zC�aWz/���7!ɼ ��s�|�ۉ��"��"8�|D|�A�>^6GNu�ܛ��U�f����� G�~��b�DxA�E�y<���ۼǄ������c����ޓ
�{?���M?��������NHr|C������������<'!�@�4�D}DW
�H{�D�ʗ�[���^��ʖ{�",} ��OL}B"�����{v�����i�4�SϿ|�����y���猡�5[x���?�i�ߝ�g����*���?@ri�#�����c�}C��$OvȢ��׆���V�����#�">���"�DG'�9߼[r���i�x���0��I�'~�rԟ���	<>ݹ'��}Cˉį�=|���$ߐ�Hy�x}~�����z?~�'�봋�������i9�}�D�Ӟ���V��Sd_?�݉�a#�����T�\�y�2��+��n�El�\�=��p��U,��w�X��`mT�[���n�zKߴ�#Ip��3���O����f-��o��4�<`�fę�p�n�S�~������oX�W�|2�R<���:�H�+[I
����ң�Q�%���j����׺R��nB�%�e����p@�Cpp�;�|@�}x�L�VtQ+w~�����sY�;q�6S���R����'gX1���f�4R/Ve6�wq�;����5[q	˷ňc�D��5(h�}�x�l��4���5k�K�>�b��l%|��[�R�1��eK�	���N[)�1���S�@�3�uкXp��c7y� ��P�kG
��؎n�v:Z83��W�^������Gr�y%� s�YWټ�-�т9�D�; oK�L!����+�:�D�u�E�h�~���1�^x ���yӔT��}T�۬q_e�O�HwJ������1���j��N�<�("Z/1�l��u=����ԁ�}R8_�Q��3���BFb�hW�m<8JGv�6�Y�w�R�;��'�B�/�1��9��y7�
�]���E��E3G����r��tf�+5]s|�WJ9w��m�)�2��:Ln��}M�1ngrqV�'�$�JJ��ohݖ!S��M�V��p��HTaa�{^�������J��ų�f�U��vQ$n1Q:q�'T����� �����:����ʌ�卓��6#zPv�\�. 91P�2>��ײ��{�A�x�4�Չq黻Y9�Ht�ɴ�:���oI�Zu8��3[��z2������Bd))<ˁE��)�fm�����z�T�9nA|�^Z��
}= �r�5���Q˼<Ӿ�ˍ��&���3�)�+ �UڲwS=%eG�f�n��CR��� �`���/��D�|��0¸ʨzo\�3Q6~]�������t�޽�{ʦN��qΈ�`����#�D�NU��_�����=��:�ѣ����;�ִ͖x4�-}�Q��TN>�U�L��҆��ă��@Xu[0![TY�5X��,{P��-q�^zN|�K%�WQ�}�@���q�g�~yp��θ�:#D���ĩ�Av�*W戚���0��y�kݚ�4���Sޤ#K��'H鲸Ћé⿟d�&�Nz�6U�=Wy}�^�*3�P��0�s8���w\|��X��T���nZ9�r����q�
���I�9�ھ�~�q��tt!^é��*k4���*�w	��i��⅄�]�����0�$[=�gV���)�-:�_�+�iHU5�k�� 1)Wa�V�F�G�/$��o�y���;iz����x��7��?'uY�<]�#�h����<y�ͫ�q���ynb����ޔ�=��R븦H�EC�8*ݫ�jf��R�Ξ���)���f<�I�������h0���U���ˢk��Si��A}�d������-�ty:����c�����t�N|��p�Gv�3Jru��s�=ز,��WI�*�+X���S�^#x \1;JԬ.�M@f9�hhO�J�$��ZST�r���1qNdl�j-�q6gKf�j�8!�9�c�"TʓĲ��΁36Ӂ<ި��v;�L�9�0r��|�5�!�eS�_��ͺ��wx��[���}�� <�'I!�{�M��e��bGg*c�BV�a�a�4�B��{Ssں]�s�U��p6��J��V�X�����e[�?:�X���u�5S���7�<}:�6�i<�9��+�j�}�
v�1���'��+~��0��)��O<���^���V�����]�S��U��}��Ù,�x�*�I+�C��3��\6̤k�4z�7��~�&��[e:�Ҏ5U��6x52��R�H�j(��9j4ޟ�沎�,���I��NS����l��`�=Z2�&�m�&�}ʇ9��¿��1[~w�A��/=�)5諢k^g�-s��V�H�j .8Vg�p��vxK2!��R+���f�b ���|c�:��[t�'�~y��S.y�z�t#�H.��1�U�.����J�����>�\�a�jvh��rb�ΕԚ�_nP�n���Jw���\m��c�9؜'����#Q<�r�n�_.Ԩe"������<�z>�B�²�/o����4m�z�L�C�H�����XCtsm�\����S	U��\RIFg)�gEE��}�	
�?��gLYٓ;��\
L�k�����>6��{.*yy3d�����b'] /��u�s�[��y��t^kyX�	:��k+�c�f;)��`���p��y� ����<+�K�9'��u��tU���Ij���4R.�@������6ph�;M��P�.�ذQވ൳@Q��)�mr��3|�0ϗ
���5*���w
B�i�-�#>�{s�� 鉸�*�����' ��S����WU
��g��a���L,j�,�iоOk����0{��r���<8��W��%����bc�D]"b��xt��e�S��vzr:?;s��0� Sm��{�w{�V!�����RTC�ȑA�b Z{>H�炥O��3��^�3�{_1��c]k�󭩱��r�D8]ư\r�qˠ#�� :�<6Bd�a�����m|V����#v?2�7�w���f0L'y;6z5���~��K��ɵ�?=���|�.��Mm}�8���0��5�(;Os>��0�4��=�Mz���$��G��uF��Ʒj�sT/�,�.6c�!��(�R��Q�˩����(�Ǻ�5�+gT�8"��j&]�|��k[�:��an�uw#�vib�V�'��/���Xö���[;�����4㝹B�Y�����}GLݺ���#pY!#9(+80*��B*�Sn#z�_.ǐ�-�B5�8wF Vmo���9ڽ"GZ��5�
�O^F`�h,����:�Z�CiN�!���ԑTˀ�`Ȝ5��E�޼�Cێ�J��O�u��l,�=g�t��*�����!�����;s���t�?3:�{fF>pK�{��\$u�wK��\�ᛁ|����\,����uD���]X�#��᳟Ta�����W��6�v�湆�K�i�CE��<{"�i�A��b����+�и5/;ݨ�\;ͮ��L�*ua���|�K)�sP�1u��"�e��m�:o'q�\
��s�e}3�Q֤���WL��78�ѱ̎=��9|M�v��h�Z;w���?Uj�
��R�.��3Rrs�a&��2�5,"*���ͪ��,W��ȽJ�;��9�{�8]PF�:w\�u���I�M�4��Y������C^��΋}�([o�}.y�u�V�[ר�}H���C�2*�Q� �D$m�a��~�1ݥt���.�VsC6f���W����Зq�k�&�JZ7�<v����;��V^֕�X��&�mh�]�)n�+#\[�`k��Cٙ�O����t+�O�`} �&h�B�.�y�V�.@:���\�7v�w��"�\�5U۝�P�k;��X�����l=�yv��V������6�D�U�><���M S�]�r\��P`��$�f��n����39��!󅳈�i�g����3����Ù�\�6�ݮ�DK�4�qt�3}Q1���[������W�B����U��"����ĭ���~zk�J�a�1�tj�
�9���H�\qD��1��&�\}�E�1�n�(=���p�Uy��3�{^��#p9gY�c�&�^����W��b/�S��8��B����d�@\�<BФ�a��՗��]i���U�9��_9�L5���x t	��k�4�7���W��{J�w��C���s7�g_^�~ *����T��y�:�ȨJ@�Q�'Wġl��gZv�My�]*�O˳��E���{]sj��ژ�GS�7�;d��;����`�X|����ഄt�ǁ��:q��y��_��.i�CƖc�F������;��:`���Ӗc��'���������~�m{^�p��A]ŭP��	��a
����6�.���K��n_�U�;'v{n����S2�^r��SW���r��{֡EXOiַ���<01�¶s� ��B�)7�dk8�U�T23*�nyK���:�j���Rq�v�A��q�+��m�,�S�`�|%�y�A7�'K�x�i��=�}�V�Ô��X�j���Y� �p&�k֭��h�B�+�r�U�v���D-������:"y+�"�_n�xr��k!!)�����Pvn�)BO�(m]<�����n�:B���.�o�8�cq�����=!t���++7`�ʅ��^9�]s�;
��|@\fZx.���!�Vسwq�hazu��2�Y]�K�7�����B6�I������z�O^�B�he1r��Q=w�3V�E�z��	���ɴ�#X/A-��|��u�[�վ���=� x\�#F\�L�p��	�+
$�dm���R��XF_d;s�ka㽔�3Um(��P�O�t�G�h���5� �Fj�����k� �Bps�}=8���w�1��,�|{,aJ�AjtQ�'hPc�Ij��C���X�2�֋)怸�J`���G����ŭ7Y�m>�j=���Y[��f+�fm��(�&:�n q|��f�
n>�l_8�!Վk�n8Չ��*nI��P�V
��Z�u�����[oK��>t�D_i����enS�Ys�S9ʘ�%]o7�q�E[��j��7��[�@�<���J�S��E`o^�a�Y�|&B*�<'9��.믺ɶ�'�W,��ӕ��9�m�.���ਭ�b�phǳ��w�}�֒s4<b���Vf�l��TN�Sk��M�{I�[�KV7�K�xܼ���m�c��3��)u�!���7iʶ�M��Hs��u�.P!K�`��^|acZ�C�e������|1���s�Y��>N�)c�	��Yy/\�9M6���DS�'v�l���`:�q�5H�V�"qV]]n��[� Et�u�B%���M��W.f�Mf³`D�R90� �z��p*%{e�\�2N9�	�����Xi>�ym�`!b�s룴�訕r�\�9�4�'^^*�C>�$J)�g!���r,`�S�/>�w3{�������o��6�ޫ��`�Ƌ$��8q���P{��?�,W:�-���6�tr�ײ��L4�$f���G\Ps"��^v�95Q���Gci*ͲF�K,�ҕ��z�EMLF����2l�i�k1Ae�h�W]M�m�4�u9����g�ZVZ;�҄qL��EҬ��o�8����3z�2E��ܦ��V��2ӷ"�F�N��v����jg��Tt	]10�wϤ��	=��r��F+�u �K*�T4�[r`�kp����$Ӯ̭.J�����' 5ve�/N�X�����g�:Z��v2��4�%]E���+���3��c�6$d���v���b��D�ʟ'�)�dZ4�Cl�,��_wf..���~<�����.y�%@��:a�d��Q�b�wnQ��(��Ei�$եE��Bs'v.�9p3��D9��B�.�T���r�D�$�Xi�U˙9$���ԏ2(�=�)��wBL�͡AJ!$��wJ"�$r�9U�F��)�*((s&T(�b�;�QED�/vТ�hi��J�$S��@�Z������ �؉�%�HQjWu�;rI���Ad�����P��rI�L��Da�-
���\¢��ER��@�)�z�EJ��3"(���A,�O]�M[-"s.x���.-r.��rY��8:$Ug#��,�F��B(�4��Cf�fR�r"�DY�tp�L3+E�E'[�ܬ(FQUQ\�:PwES��J��$�9�FQ��(��wn�^�x���G#S1U�nm5nNUr�L9����I��!��ʳ!-n������@Ѫ"��H� �9�7Z{����2�aR�uK�KpZ��+�t��HWG���{��U��5��,���cu{K�vKT�0�GP��;YQS���������x���#^��T*^Uנ��H	��x�o�0��S	�h��c\��!�n1�fQ��~F�w-�΂���o��`�BUy�sO�j���U���pHO{�rK6���;+�m�k$Y��w 7P���(v�>�4W��G��:�n�D��N���_E�+��"=O�Ѧ�}��_oTj6;�ȧ]��rD&l�V=26�� �s����0U\%'z��[����1����vΔʌm�M���ۙ��2p���r(�T�O굚�uQ��):K�L �ba���'�S`��Ζ��	������{sYv�w����n��c~e��[�8�����=��(��Qx�}����O�l,m�(E��=�⤐[Up�Tz�Yt��>0:�f�y	�IZ[õ�������t�u׷�e��o��':� �6�|̈A����s���>�:i�<2����u�Cu���\��Y���Ca�Km��kr���]1НQe��7w�8n?za%�e$��"%���X���ص^�+�Β�s����5Y�-����;)���HFORl^͏>CZ[���&#b�+z�Fe�s�ֳ��#��<|��㕽�y�^�{ s!mu�]=n��vT��A���n[��V�6��g�q�C����K��l1Wf�ҳ�ꯪ�K��5C'�5ѡwM��ʭ���JeI�1��-�#ı���k(�ۭἝ�<#�|��4L �`C*')��ʯ��X�9�F�K��q����s|tN���	Èg)���u��
Q,��?��v_��l�\"���*ү����ce_?
&
�܎��VD����p�ɋ1A^�5�Uއ�)�8V���X���a3Q��_\�"���W��6�=�XK�8R���
>�8�	��]mo���]s����m�S��U'�Y�뺃]v��d���!5����&�������c��vS�4_RՖ1l�Y9 ��Xy5^��t,���/ua��_��A�賾.���y�N�84B��{(@t�d��ng*
��V�)�4�y�@�=�@mǱ��<<�(�RW�q�:���?�*Lƈ�0ޮ�W|�b|���#)�D�F��EOQ�y�ÅL1w��W�5cx�u�~>mk��̞�#�V13�O�\��"t����H��:���c.�+uUޕ��c-N�C��=Q0.P�c.]YQeأƗ�_�J���f=��l^'�h�s��������g�wޅ�f6�s�^��L͹vf[��[���p�go7�y��j���b,�Җ{u��ۄ�&�or��D
���T���d�[Yej3r�u{�Kƭ�}U_}��ض�Sͷ��M�m*��t V:��t�
�H�ñ ;�5t�Zp���.aQ.�N��l��r��3�	�-3L[}V�|�����Rxl�NH�0a�6�g�nUQ7��sZ����_v�F��#�ʐ� S��loj���}���5s�1�)����o2�pb���v�Pf��[�MM�^�G��
0w�L�*7�TwH���])K�a��HÂ��|�i�F�J5vzUԾ~M�@%Nፎ{Q�w4�MZ봚�{/ڶ��M��d1S��*Z߱mu��:ͫ�컯5���3��ԍ�^�w.���*b#�֊�_����]af�Y�[@��y�"](K<�3,��$V�U�
��X��d�b�mW�˭����;ϧ����C�U���I����=�\��|�fq�#��L^.�!��j�e�ܣ���C��P���sӁ�:[=9�`�`�Ҩ{��1_b�L�*ua��a��/x迟�`cf*����J�,�낞�n5�����ղ��L��,���mn�i��٧�Hd��w���61�%ʃ��9�G(�í>�a�q�u�h#��jT��N��6�8`��+>5�(h����M���1:5l*�:eD���v�{P}UU_}�w��{�vZ�,��P�X��t��T�o��s��J�Cϕ���/��e=�����
��T(]=���e�D`�mĪ!7�\�!%E�jw#U�'Z$K�b&kr�	�ޥk8s�lt�_8Z'��B�'���1���}�UD̄�*��r�����;�m$n7�+��b����H���W��#:���D$r�h�[��c;�|�j�3��K�n3Nc���+�M+��U�1`;�ޚ �^�h>K��>K��D�%^l5sm=�bsy(�	�p|c뮥�vl�!Y�L�����6�I�J@��8��c_8�uu^U�X�u�*Ԑ� �a�{Uk=�,m�@��%L���s��+D���"�䙜�Λ��g�[$���;fR5����vϭՎ����3T�1|Pt�\�+P"v��{��ڒy�~RǶ�E8E���[�oM/�"�t�߽�q!\�y��X�K�[o�K����+W/�p0�5h��H�#�| ��t���a����.ӑc��~��[5�zw-^Sk���&��Y�^U�>{]��;��^=h��F&"�K뇮���-ͼ���=���:�&+�v��Y�Xoz�n1�C]��﷓�V]��1L����h�g�?�:�4Z+�ۣ ��5en��ꝥ���7nU�Q����"";.Ե�eo4���G�#�� /�l�i���s�j�ք�bí�٦O	��]o��se��k�Gt�Bd�smLF3z�ڝ0ְ�w���yCX}����#XN�橥�rL{+�`����<Vc���*B.6]}���`�9l�9���.2�<Z��Y�ݱ�K��bz�z8�u4��ĸ��88����G^�Lt���}�ahVyn��g�]�O y��)#ro�e���g��1�D>=5T���Y������{�G1&P��jo�n/j��GC����TRF2!���<���B��b5�� ���e����w�<��[�����)=�x�BމC����;�b�ܔz��Gt�(!L"�ķj�;+]Q��ޥ�x��e�Dj��E���.{�|����7ƴ^R��#�D��`
7��AV�.�7vL����0T�1p!�w�֙ȍL:�po��%V+D�#��R޹́2�Dm�ץ_t�7.Ѐ0=����ʜr ���g�-1�������V�9e�T�W\����g��f	��b�&GcxrQV��>�,�=��l1_��Ky��%G^�+Ɨaw��:G����H������i']C�ݑϷ�Ge�7l%���%��Wh6'��0�ͫ��\��똺�g�Ĺo�4�R�}��}�|����}���?|�*�k}q �x�%��z(��|M]S�t��ަ;�*cs�lNB�-�t�]�f�"�Pz�\�]!��,:��#��'A'��u�-����_���im\'�����N���#)�;CE�f����R�S�a�'̞1�J�f�3�P\D�v�h�'��UG8T�qϸ�3�Pٸiv�g���#D�uP�\�?�k���J]56?A�ǹNs��h^�#^l����ٿ�e��qt�LZ�l��QD�F��zb$��=�fbN̆�ĸ�I��a�J��,�[�He�g=z�����PcTc�B*�V3����;S�^�=z6�tnzM��h��R��4{�`y���T��Q;<%ZU��� /��ŕd^�`1{�0�*��Ȯ���/�؆���z�(��	Hܘ�Q3	���P���E��ۇ�!G�-�T�L����O]!b;5�|r#T�/i��[l����� ��xo)I�B�㲽Y��e�nq�~®�fQ��2����zˌr��ȊtƋ�Vu��I��	�`@��(KýK۾W�������+v_@��@0���Y��WL}�������gd�S�ϭ[��*���Y��޿��P [	���.G���Yq=;���J
�ͻq��owQq��'i��sMvZ���4�H�˥�F���ﾪ��F�N��M+z}�����2��ƣ�뇐
e��F���>e�.���䚛��uG4��Q�0�6�+B:�͔�0�<�Puq�W�t{����v�����3X��u��k]V+G����#�;��R��5���wǰ��P�dF�
���dY���_-=-�'�9۝I	g��;=Bc���m�
���=���4;8zR1��0��J}&�;+vN���V�*hGC88��@Or�F�#�Oĭ=s -5lO�����&s���gr\�����σ�p���ճ�]�� <�!����Ձ�fl�h��S����h]rG?�Vɨޗ����4T' E�th����m��a$�R�UN3+c.�_Q�2[��5s�xW�c��o�8���Ʉ4�����1>������TQD�|���px֕�����m7ƀ�Z>�L���WdV�|�
��\}�|��k@1�<�q�Cϊ��x����]��
{�57�n�h������²����zĽ��d���X���uN�7y�%%��+M����;Ǝ��nE���W�}Ho�%�6-�۩j�c���2�r�b]+���<�^9 ���n���nܞ��b�f��[ԴݪTq�[H��h>2I|�Q/��]�YϏ-�l<��fb�Ԥ"�X�o^��j��J����f]���T���}_}Uq�7��%�2���,ǂ��<�
����l�����Y�R=g�t��M��ھ�sV�]Ӊ��K�q�� =T�����a�Gw���}¾��h�xC���%sĘOwS'�ݒ�4�����˪�3�$���s&��)�xu��9�}[���Y앐�]�r{�,8�hX*g@��p�Z���9��1�u9L�v-�p�;1}������}�����4�����
�IGyɳ���!�n�v:Z8"�Z��>l�"Q]��+a��S��痷�R�
��v@ޙrp�C��̬�V%s�S�w,�j�ʔ��fy	SW�Ã��0,��ڸc>8�}C��&d%u]F(�ƴ5IQ#�2ո�:�2sZ�+�����\p"�:�9	� C�F��ȨR�GX(C	��X���V�{�C��]��d)��Z7|�;�yG�����
U^���-\���u~Wۇzq5��uJ�����F���;�3L�{��v93_T7�[��\�]�n抶/������$�h"��za�5FɨTI3p�[�ђE�]�NV�/�!z�]�U9o�z�y�]���W���7FU��*�S���ku󼜕�W��_v�	@99�b�^�o2�h�s�s��ꪏ����;���xZ:G�� i�1�z���"��
�v�;u_2�1h�:�V�&k7�xW�W�=9��G6�2�|}��	���*�ǉ�3�k�ɺ���C��GA�(7#\�Tꩨ�����D�:{y�Pcdt�G5DG;��+���X:}�Tq!\�y�wN��t�H����A��x �KZ��Rs��#�Tm�>K~ߩ��t��k�Y����r�ѩֽڧ�����2��s��&��ȦQ.!�������u�#>J@�Q�'v�&���=��=)b}���}�:ь���-T�F��c:���S�L1H�5����׷H+̷�f'�ޯre
a�#l����Q�*��1�J��.~��v���M�ƫ�3D���`N��M�K��g�.�}>��:`�+t���� �*������+ƴt��y㮰�$��|�l�m��̎����~��M�}�K?d��ӳ�T���w�&� ���
7/&��W|�^�yJcql1�zP�q�'�ŧ,m�����c
e|LF�U��ƝZ�����ǧ��(hk�(��R�,��ռ�ng��u0cYv���r3,9Oz,ˤ��0���3o��zî�m��Dq8�+@��fhEP�7&8�eA���;η˚��n����Z�__\)j�O6Sf>��%��ˮUw�.��F#����_N��c�DD}��f��ˤ��Wd��+?F�!Qoj��8\<�r����W������#u"�^�����K�Ξ{�0C���ะj�q{��5{���]�>NH�F�z'[�r3d�Qg��>�p��1��o邂���|c"!�n�3p1�Q7�x�e;�g{by��=�7�3T��6[b�6�^��`�
w
�_�f��0Y�KLg�_rv�Nf����[{�[T���q�ɇ�8uLک����R��H\V��}�rɉ�]Q"��1��KIy=Z��T�n�]�MZ�>7�{����=�PC��x�#��.��J8]��bӋ��cYog.���Z�迸�5���a#��j�}�
v�0�9���(nSƦ7n���친ޢ�fI��s{P�{�2��o�m&m��c�,���#Cs0��8r3�i���1;��q��UF�'��0����;���͙C�3�!R�lj��NBr ��}>�כ���~k�p�c��p�m[�r���(n�y��W�L�
�U+������N^Z�ʽBD=��VT5���k f-�vQ��[Q.��s�4�`��ZNO�ު6�ru�l��͎�*F"�im�ï%�/�Ƴm��N���	�Cn�uwY���	d<�U���]wS Wn�Ҋ����#��=��oW7�ɭ����]�'�{�8�:�P�ots&X�<p���ʥCM]�o)ܺ����o�*Ӥy�U�;oV��w)����iԠ���K9��F��%=�!�q9�����J�+�P�������H��]��B!�s^:r���Wv�'V����{��
�uv�e�Л ��B�Lܫ�E��Pv�v�Q���ےC1^hfn���p�u(�_Pe@n�h'�hbov2�Q�]}̵�SΕ)L���*����c1'���tj�����]�hn�r��
��B��q|�{��������L?J�ۼ\��+@�2�i��sYƣ.����s�Q�r��1��;®�]�v�TU���(ڭ7��PS�����m�l>ͽ:��C��h�g)��4�yP��l�������ޝ��Z䇻�f޺m�\��V'����;8\�Ӎ��yQ@c�ӣ�DD�[�gs y)�e��}�DL� \�h�N�\p��wftٮ�3��ꐪx+��������wUu�x����n����ܟE�*��(U���ʹ2w���5y��G�<�2�S`����쥥a�`��B�����b:�5.���սSm�ČF]�9�L���:;�sMv�Y�>X�"d�Jfs��P��Q-�]q`sh-{�!e�.�a��Z�
�h��GKWq��sCmw%	�#op��{�T�쭷�zqY��H��`��B�]�9�p0`H��אb�:]�ޘ1Ԯ7�sK0�m��/K���o����nw	�{W�}�
إT��걵�X�#�w�1�ꭉ\�R���3\ښ�񰶡�M���=t:����L�V���|��}w�;Xk�9�y�j�:�������P�]�Ⱦ�y ���QWOnWtֱ8Y5�]��w1,�3�8�:(A#'̖�"6�H��Ї;^��ג�9`}x��ۥ�t�WWM0m����i$���Gm�6�J-����rRsI�q���f�j��C3���n`���F�� l����̓���#)`�i��`@�{�3�4�Q#:�K�8�(�³[Osi��1.���o
�qMΎ�r �E�B���z�V��:��W�0�5]�]�"�6�1�;o��v]��+Kf['j6��kT���ۤ$��ZD���zZ�X�Mq䴽p��#��i�4��IJF�ޘ��ز/�8���L��9�"Uo54���1h�z�@�dTf]��3D�"TR̐�s
�dDV��'�U����)�U�0Њ��l���:!)��TTC��r��J�a���"�CB���L��^%�$���X�%��i98:(aQ��p�­g,�$���#�f�9�g�tжB)Q��QB*Ȕ9�2V��Tt(�B�J�V������%Ȳ��X�"m-J��r
9s��Ψ��E"u�'C�1@�!˩.����Z�]��Ȑӫ*��QL��5������fsȊ�*�:ny嬢"�r�#�L2��h���g�c��eZ��,���T'���Vn{�*J��"�MMM������CՕJC�%z�EȨ5R�"�����J�%$�'qQ2�4;�s����OQ�s%����E��i`N��jTX�T�$�v��A�:$jTA���"h������V�RF����95���,2�P�Ԓ%v�[�au�ږ�0�c�gs�@[����r��KA��1ͱ;;]����\�عnp1]�ĺҶd:��}��W�U��1�^������o�*��V��������y]gj\d�1_a@GD�z��	�T�r��x��]p�Θ�*-�f%�'�ñ��Ƨ�awH�����t5�E^�ƻ��|��5�q�R���]���مF5k��F�P��E:c����Cz+�f�����67>�s���t�W���Y�UG3Һ�cS��5�f;>����^�Z��E��oݺᬱ��y4��=b�r\Q�1Na���ȫ(P<y>�h'M�!�=�"�H�ŰM��<��F�Z-����.
�7�Ԁ�:/)�h��q�5	[ČLUWd'f��jo�f��ͬb��wS׹�����J�ܩ�e��;f�*���q�T7�4S��M�wE����م��x�P�Oy6"D� �=q11���\a����v:K�2��uVO���<�ԉ�q��SS�����]E��H�ó�H¸I�u���L	'~�wڅÊ}�w`U"�f�\7�l�@G# �O�_'$@#C�&�
�(�����y�{ ȱ�m�4aeo�B�����(�u�5C�CG;]%�m�V��^��gWA�(�_J�Cv���ʶ�P�q)���v���3�T2��Z�P.bӛtXycm�bk+n��3��jQ��z:���9,��/o��7Q�����q�r��[薜J��������w:йQS�U-K+>��:��ɯ��qvr��Qi����/���\��or��F�wk��]�#�V'.´:p�-�΢���]lfm9�~=�Ƨ����4B��V�`Y}�.}^ը1�d�W,K���|�i�mp𫇲�v �U|�
un��'y�
�+�mV[�r�M�hV��p�U�`ciL�G��b���`�
�����xP�p��E�g#tf��HڽN�����jH����|��k���[�ؕ�a�H��u�����oԑ�8��-v�T#\>�f�m9Vu:?Zy�K�>x�yq�G��=�v��ϳfI=�XY"lQGܧ�o��a��xs�K���b.��#�ULm����a��,Fi���4@f��ͦgU�P���Ϥ	OfX��(�B��L&n9[��<��R1�z�.��V�z����n�1%��W�g�Zik�x	T�o��Z�Nl�O�ޟ{>8)�9�]ͥ��LK�`����^?_�pB��U�툪t@�8��<�������T|_ļ�����t�)�PV��8�n�F������S��'�vt�Sz�p��_3pP���֍E4D<)%��s��I����xk�{u�'[��-�x�"y�e�д�@	/ ➎Z�\�/.�b�U��<�%vt�<�M镺�vȺ|��ﾏ��-er�۷/�d��wR.5����Ӭ����vrX��}�UL�Jꦊ����gQ;��P�%�y�f��خTZ��EB�]�=�L'�F���E��j���U/��fs/:y�Ei�2�g_0�U��9�s����@�L�9��4h�<��^�)��;%̰�W�Px|~�;�4L����}M�C��\��BZl���^��$�#W}��%��
�W��s�)�����gc��.����IT�﹨������3�����	|NÔ�`�J�n�X��#W��`V=���Q��x��Np�\� WLdB������l�x-��9)c��+�]�wydw2C�zڽ9�u�J)��e��@�s�=�T وN���u���#�D�Nd�F�`��%	�䖾|�5�W�y1���S=9�lQ�8�'�a���j ;ّQ�RأF`Ѐ�3yJ�u<(w0��zN/c��?,�?=ʥ���v�� P�}���W�d\��&]���V�a��<r26�vaJ�ܕ�`��j9b�X"��r���fb��55�~�L�w�2�W��'GY�X�_;ƶ�wM��p��ǫ�[5v��`�Xf�V�5|,�����S�(�����G�G���7��8⹬鬉�NB��f|���u�ү>U*��
VK���s�Ƿ35n����'�y�J�nUws��-�2�A[����� ��%}�VH�u����쭛�=ԞV=轎}U5��q��7M߭�D�����g댃'��MDU �>$}T���І��X���u�e�B�ރ�Й֬ҙ�Wp���۹A[����b%����d+w���ۢ����.} �{h�J#j#��'�>	� �7�BwP����:�A�]z%&���i�x�q����3��\^b�R�H��H�@��9�X,�)U�[�kaӶ�1ƍv�6`�jL\ĉ�*_�:�nu&o�m�a��O��R�d��i,������7R֓g�}�. �.\���t�V�G��}��v����(���VԮ)g/U������9bG*��>iJ���6���H�+����k�LM.����[p�Z���M�������Ĉ����g>r�58$`t��Lr�����n�qh��+��)�a�\�#��Un	� ��LYg3N�W`�=��j�@z�j-)�0"f��?�@���W�w�W���k,�������kc�oV��1%�u����2��}չ'/������k&����5���䭵���.�������zm*�s�����������[��V�y�Oކ�ɨ���
�S*!�4���E����;v(X� �:iR��G��m�w� �����f�C��\{�p��	��e��d��uDh�N��g23�J��Gt��"�z����Ŀ�)����cҭc�>�\<�qWTEB�Ln��&����c��17������_ٓ�~�y9��&,o��mp���+\^̽�7��W�*ٴ@����yC�{�w�vv�N�Ԧ�=�<���@1[P]��ף��9E;<%�^�ùd^���ߺ��{��������n_��8:�����]c�����n��|�����NH��g7��F��3�����F�*1����kul�czV_�.�\;6D�͖�]��ŏ+��sW��$^O�+u�	F��V+�L⦯끬�7���,h��wN@w�K9���7��]����ը�΁�7E�F����VA�ƣ��	�e��v�`���'�ʅ�GiU�wW<��!��z�ǻ�@��7����.Ph��:�
�C�1��@�2'N�����;��SY���#��7b����n�hB2�P�`L�۳�
����\o���3p���P/S*v�A{%H��l��0��cMMͨ���g�\ ٣#�u��#������c����K�=t�o�/6��6A��/�����L�#���i�f�1�ARg >1����(Ҥ�;KQ1?)�� s=g~����9�u�r�L{�u3�fO{l�������]�򿽨����R�@�vR�[踚�	�rP�6�.�2��q$��\Ys���s��'I�U�������w�+���"�1"~%i�\����y��m�mj�X:J����0�v@U"�ԙ�ګ�pԁ�LX����P�����X絬"�7Pg�_^Q
����WG!9�	�z�:��7�gx��E�r�$��m�]8��I:8���(C(!�y_*��Q�����M4��#�)���v���*��|�1��v�Q�p�T;�<��D ����c0���B*�Sh|Z7�]]69C[v��J�<����������׹��s����&Ȳ��L
ФdoD�2ubW%<�:sePϥ%
jHֶ��՝�ѩ�~��߹�6�9tG���B�E�����ؾw�״�dP���V��q��&���U�5������+�9���ofy�w��}L �oh{n������'+!��4I���E���j;�k��u˙*
JU�rV�oޫp��N��
��~�tVDm7y-�G�z��s���n���.�B��&�Vεk9�y�ظ���&ή��)Q[�C�T�-�_���������Kд�w���dز��Xx���1��˪�}�*�r�OK�0�Ì���^]���R��v�����ǯ���|���]d�V)��§V|�9�H1�F��M�yη��=FeKڿ���� �8@�JDT�97�O"�U��w�^(�i��̩ůjW���$tl�V��aq����h�~�̿� 3e?FA0�m�V���\&�ȕ9�%�^jv��s����D���W�����f ����1�q�����W�2����"��VoR�Z��K���
����~I�)��p"�S���`�4`�Q�H�R�G=���Z���W5�{��´Ud>�Ɇ^��G3�*���Ҹ�uQ��|�+A��f����mpPE�}7� 8�Gd��P`����ye3�@Cp�ɉ���b\��|��-Ԫ�������X����0����l���Q�>g�_g��;�}���Ms�¢'s��%����~zT܀��I���s�k�Rn�mT�xb6K+���r^�^�&��2V��(��G�n�'v�akeh[)fFu������8�W��̊^�}���8��2�)o��;��<�r��$�_�t����qf�X�,�7���Q
v��]�}Ԗ�s�9�h%F��xzq���*d���_}���k��]�/Sʣ��F���ٹ,\9QI�"*9�|�,�����7%q��v�yz5lM���66�	|�����=5�����0����Ψ��7��(Չ�Y8iuS�������or�
���'�א?)7�+)^Ǟ�>�����t���l��,�H�i�e��I�t��n��8 ���`z˥��5Jo���R���۶i� j��z�{i��޻��v(����I����X�l�>0t��B��ZY�S�|�T���o*r�kR�۹l��{��T�-t��l��r�*�>���f��
��K�����+�ק1w�.���@}���=-��畋H��$(¸��Bj�;��C�Q�{�x��hB��S���)���K!� �� ���6Q�\#:�w	��i��|zP�c��0�c::��"ʘͅ!T��R��j'M���nDf�� ��d�a�V��G����%;�/��{dh�wP�0%=��1G{^�P�q�pۀF)��A��s��r�q{��6;�ڥ�q���k�&*�HQ1/2���J�+U�
�8TH�'�Qd���_nԃhM�轢�H���L%p�
��V�a_Q�:�	F�z���7-����ɾ�{�s�H�(%u��B��������sCmQ0�5t��R�������h$�>��W�D}�X�{i�dh�̾��0GP I�9]�Ne��5}?R����"1���fS�sg��J�<k>���uwJ�#*8�@-��Z��5�HGl֥HYW�Bj�8��{jz����7���+z�-�b�ul��܋�VM$�6e��ܒ߃��n�$�����៞�:ݑ��a}��X5Jջ��Pz[�}U}�c1뫎Oj��9���5��{��v�mB�S�]w�f��oQ���ѳ�E.Ҽ���y�w��0u��ި/��T9�I�K�͎��3��w_�{F϶Q����~+�AT��ެY%�f�o���7�Jy����ܭl����m�N)�}�iN��Ww��Py�A�a�m���}PI,��=,׏d~Pf�WKKGC�p��}����m��#�l���\�x�Zq�W^&�[o�U槝��u}v;���u��Z	I�O�5����@˗2�uy�^�KNF��CV�f 5�W4�b�6������.�����i�<flJVu��Z�!���v�vgu]�T�4�9�O&�Q��K�Hx�k�`t3�s�YT4���b�N�nvu��lsʛ�����~����":f58.�9���T�k���Q��-k{kYkr#[U����o����rW��9��<ks�,n:��gt]I����e�IvSz糦,��������d��@샑��Q����贬�O�@�ݴ���Sۓ���}���Zڜ��g!���`]�v@Q�R�B\-5g��xT=Fm�)7�+���Kg=�_$��p�d�;����;�DJkfT�ݿ)���u�̛fOozx��|���6͝��p�j�v'�Q蠷��>���n4WWKT��v��5���y���M-�=N���	�*y�1�����3�sҽ����:O
k6^y�M�݁nRL涩���B��Z�X웾�d|�	k��������2�:g�oڵ�j{�Egѩ��Cs^錛u/f�`y+������w:檡��7��K������N�>()h�������w�	F���n��B1��
��)=ܭ�!7��/�*�	b�� �.�t�o_L�4�[q2x!|�v���Qڨ)�cTxwm��F�b��+$Vetqi�G��^�WB��ݹ�W)YRe��J=��r6j��tںR��ꋲ0��hwփ.v�lp���Y��,q�O{��3�7ҹ:�v��5��T��i*3N�ZmP�XԷ,ry��e쮹��x�'�6h�f�j�uI��S���0���le��J{,�!��=qv�Z
�ux�����`m.L �o��wooq��`ݜ�i71[�G�P:�X�c�.���VNE��L�lT;��
@_k�s_P�����l�DofǗGxu��Cu��X7�
*�{.����uZ�M C�wb�e��7۳�Ua��wg�j�.����8:�PMJk{�:o[z�ёA[#e�B�GR�/[|���֊�Rܻ�����e�[|���b�m�]y�le*�q��ۛ���L�]_rQ��-ޚ��)*��+�ý�ƒC�Vϕ��<�;�����c��*|�t1-�����<���NԾ��i�Z�%(C��w:��]@qcd�Y�r��,��smQ�]� �RS�4}"�,�U�֭�y[���3��/n��x��y�D���+8�t��osXjb��q*h�@�;����c"V��D�o	�����,k�Ϫ<�}��lP��;�e����&�n�h	L��#y6���2�7i>;��_<��Sod���V����Ь���W.�m�q�y�2����7V��n���'ssDn��`X���ģ����J�E��sJ���O��'I�,��3�3�r�2Rꝷ���[|�!��g)�.(��bެ�}�H��z\Χ�d��y�+Tpf\��Qۤ���u
���1��+�̵����� ��+N�Jv�5��}�f�yvt����)*��٘�^[ig-b�&%�nM&i9�GV3�U��F$�
z�#r�T�£[�Ӿ]G�*Ev���e��#�oQ�®�]���gՉ��� gl��c��qm�:�H�^�u��/�ss`���j:Z$:�
��Nh6Q���v$d}+�N��r��/�v�ˤ��ڋ0���� �nr�g3�U>e�zj�"9�Am%C�J#�s���3p]��M���x0���ƴn�cO����λu�(tc؏	|��,���t���̓u�QJ�k/;���-�m�D�����ܹ׻��!�k^L�`���/�P��.�'���Ne=����V;YA��7��B!�/&�h�D�$15�M����������;/�oq�/��8��o��سjf�s�+0��f��s-�3T�Ѕ�Fr*KB�7L]6��v���%7Y�];O"��-証Ԕ�9�����#hn⣍vԝ*U�Ѹ�t��J�%ԫ�.��˳X�#���VM%�u�xAp�.��i`�����e���quy�ϝT��wPPZr4��,�wr�/2�aaJ*�^E* j�6��U��qҨ�)n�ExaR���eU�U:����/ ��p�ʠ�z�\�]�^�]=q���\��=:{<(���B*	��4�&Ne�z�z��{��+�ZI��)NX���N�u��6뺲��r)�Hr�=]M2��Y�si!�**I�;���f�9�"�I;��;�0N�hr<�Ч4�u�qLMhS*B�BQ+M��3��!�$��C�]$�:��!��I��$j@��jR�!$��]H��CM����(��H��]���:��#���\�I,��N���t���˞BE��ʊ,�(�e��,���-	!*SD���ȃβT����n���^r�M�Eh��^�+
��p�$M�����1ȗtv�䫅�3D4$un�#$�5Ξ+S=I�t��:J2�	֒? ~0A?| `D+s�M�ľHF���v���b����1��Q��y%���KDؚۧ(9��ɱu�ϸṸH�b��,���着�]͢y.�j�R�r���5^9�_�k�{h��Eb����~w����%�M����Mެ|.9��-X�c,-�����0��^<!�W��j.=���T������q�-SC~o��ml��u�-�m!�m{��a%���N����l�QiF�wع�u�����;HȾ��M(��6��k�s�dU��pv��O9���Vq��2���9�ɽ��i��쮪2�uxli{���A��M�GrT$��jT�Z�O�')t��"�%9��ln���{�o'�o�0�5jл(n���if�:���r����IM�\&����m�5|�wm��*n���G-S��3���]���칗�i�5�Rb��\饐�.�ǻQS��3�#y��"��yaԕ��&%���e���s�Q���j���P�l�S�R:-Ĺ����I�-� �5Gi��Gt��L9��e��[w�WM��i�t�5t�iµm=�b�G>�[u��9�ނ��d��Ny�w�r���C'AA���t �[�N����{"}�`1y[�Nv��0�ʲ;���W�>�>��ε��5��ƽ��r�酮��ˁܝ�����7�5�"̷��YV��������҆|^�A����k9�４��w��/j��ݗ�?G�Of�q��Q���c@��=��S�D3���y���QR��o!��J��^�p�5P��� �m��
�%v^b"S�E�6ys�=N�[]%�hMkn��.����͎yN��5����(��qA�ԫ)�����|��v*����{-D��n�y�\2����09��Y�^�Rz��|-
�����c�@j7�����|�\�á�hp<��Jk�n��mS6�Ї��.;G�麞�?*��G���sB����
��z��35]��iKrZ(q����qv���:t���Q���!4�7k^5�]o�!Qm�5����3^���Mɣ����V�txG����ʵZ�H��5��){M�y(���\�I}{��̫Y3R��l�:WG�r�\2��ޅ�2�JѶ/a���bѠΡ��zU���k�>���ܗK�wՒ
T�$0�w����ecy��y�()WY]x$]�l<�+zg#��U}�}_Q�%x-�K��G�V���ux�)6��{ǖ-Ǻ���=0_q��hm��۞�D;�mn�K�֪-Rv���_ю;�7�V�8���b��+.��%��c#��zJ|*����I��y��n!��Dh���w���MB�Ѵ���1���U�������T�t����.I�{����ڛ��1]H�B(�|#���������?_DM)��~U���s��1jͷ�Xl�'	N�X�UC�2�<(��1�b�����Fnz+/�ou'y���-Y�e�4�[��q�3nr:�OLBcB��k��'E��⺼�U%/���
U��8[�j7y�g�<���t��l�|���bc��v)f;��[:�]K�{Y���^gU�3����˟5%�#}P���b�A��m�eh3\���]Ł��}�*s���Qx�up���yn㜅�+�فa:�w~�3S��k���Wd��Z�/l\�_#��df�l���t�:S��8��0<��gT�  *��H� u�Ok���}�]�䶰Y,�o@�]��wu��߰�{�F;���8Sx��>��yܑ�kp.f���� :[��KOd�ٴz�kJ�G��"#��nW!��;��D^];���y+�Pq�E�^N^/i�������vo�sN��}���u��]�b���������z-������1�	�o])�f��K�j�*�m$��\'�Q�8�j��i_o���<�j��)u�n�.���8퐫�Q�S����Ž����eC�Wc��.\�Պo�B��8�T��'yU��Um������܊o�⯲:38�����3k{��yz���<�<�Ը3�E_%_bV�Ά���k��u2�e�nƫ[�%�q�{�4,����F��bRb���#�9>m�L��B�k[�Vn'�v�X5;~ݎ����i�.��8m�b���+�dK�]�ۖ���Z�p�D9�!��BKf@��[9tݻ�'^���,����Z�w��i�;�'���j�v&G�������t��`;�m�i �/>|���l�v��j
)hw���mz��Ga��E��u�9h���Ɩ\��p�X�0�;m����.�1��@c�\t��n�
+RƩ,�s��Fc弧֫.(_u5	���^��\gU��b����:�Pl�����򾪨��Ge��O"�l޸��Ó�M-jU63�%���S��r6�Cs[��BX��n����^�/��m�;��L�<�6;�4Zދ�?�"��𒷪)l�`�xs�W:Ȅ�~N�ܸW:vx�ߎ��H}�m������Ź���T�hs��7���h����J��o��{B�w�޸z';cs��r���[�����h]�L���!�Z�7�vw�%I�6�;ڣ�����������-~����U��;�g8��o��N�W����]�k��մ�w'�ߟ��5igo��>F=�C��r�\����U���*-n�]b�ų�s�:w���;=Lz{��~Q�i7��'���B��Է'��g��(uڏ	��ѝ������ X����ys�C���=0W�PkZ���&6c�����S��0���H��^%���0�(dh��(,��z�W*L'�e�%l�HQ��B��c2NwLja��IC#�[2W�is�>ܻsW�n��vE5y�Ȕ�[grH�;gq=��i�ϛ�teC:`�����w}���t�}�}_U���%�/y����E;���{�(t��s�T&|?mVus���53q����A^f�W���mSO�sW�Gv�oj
��XY����t�]S@�{���iX���/U[]{E�#�꙽�5�6���۶��-��z�dOv�{&xwx��Fտ�̯�fb>��.w����'��'���nUV��`ErƔ�s�=ALʌ%?WL�Z��.̱ɦ�a?�K��4Ni��%�����S���_�Ä���B��l�Y�#T�y���PP����,�V`Ŧ�w���4�*5�I��SqԞ?&8L�F��[
k��y��]�Q��kwyi��Vnke'B�bvP��NC�
��6��tiu��Uo��4�����ݰ/L��J;Jw�%r�)�6�$^�`O�·i9����k��z�������.ߊ紟���Q?%m�9���N��8ﮩ�~��9B���m|���s�ę34ّ�LI�瘍�V���B�-�V"�zw��?l :�B��J��(���Ǫb�Ҵ;�jv��]��^VgF��H-��+�9�詑���ݎ7�xEu�q�{{54��q�c�r����#�q]=t�-��>�6�ʃ���z��s�����R��C��T�̋����������c�3�Y��-}�8���Ud��jq�#W�[��(�O6�_�J����N}<��6���W�mUd���*�8�6m�`p!�k�(���v���k��b��yt��8���ݎ�nJ���j�J�	��ʮ��Ur��T�c�M���W�_e���@�6:^\_l����4��nx�#�k$����ڣ��Ծp��Z�.�o&�^���#WpȮ��E�#\�{g��`��S��)�Y��
��wE'��i\|�.Т���Z�	'�W<�9���;�Gt��d�t�+��jf􃳯��ՙ׋rF糩Of'�I��e�E�Π��ٙ}�M_DNk}~�b��ͭl�N8e��iN�g4u�cU|��LBC��[��o��N�"ze8��������)��e���r��~]��q;v�%LJ��/k��ݮ֫���E�]��,h�mG��F��dL̜��%Zz���L���6�pc�Iή�zVZI0�q&⧹�u���4	��4��%r	�7^u�BV�y�����S���k�U}UV�s�9v�KU/�w[���s������l+y�?&8��qlI�ʯ�qr���k���N�Oc{���tn�t�P��㯙���Z�X5��V���؝ܼ�V��b�W�'���p���>�Ț�:a3��I��\��{�oԭ��&5��/pO<��E����r�?#�ŧ	�Rc������)�9�Ƕݸލ�wN�������;��c�7���	����o'�����;^�t'�;��Gх�V�����[T�8����~_R����u�/yw,O�Ѯ��6:���]�ߌ�����>�m�6�:���y&�i�7Y���ܧ��.C��������������(����LQ�X4j�b�u�=�^� �K�UM}�����T�-kq�آ��{b�EPP�Kr��.���y���L�jT�j*/��O�+���g�����	��{q�Y�5ɤ���if�[Mk�xx.>����=�wV�;�w�����X��R0��D��v��*dwZshݝ}
������|�:�k���b��A4 ��]��,�C�����V����m]NB�����k�4v����f&����f7?osٞ]�,��r�c�G�I���H�w���U���ޝ��=ζ�S<�ۅ�O;h�N�X]Q;�u9�g������Q�Ȟ�ٮv�����I�K���_C�ܞ�ߝ�V-��Π�Q׻ܔָy�m���{�������U�\�+�+�	M;x�u_��Y]R�u'ʹ�c�~��yave�N�KY�|�p��Á7;Py��r%��u;�Xd�����k�g�`�Jܝ�O�@ۘI�M�f~�T�8�*�n�[h�UJ+\)�]�ccD����ڼ4���s�r{x�|�S����m����M��|�>F��D�rXV��҅�e�G����NV��-���ͭ�q�W���}��]�Dc
� ��8�7�շ�uH<��Yl��^?����9�[�%+o���6cѦ�eF��>8x�Kj��y�����kܝ�Ӫ��
�Dod��.x�k�h�ⶤ�5�b��1��))GoMۂ��̳V��2K鷕���fُ3V3$PcQk�\�95j��#� [	Έ���`eDK���۵ڈ�M��]�W0Hd:��m���j]���L�J�꯫���ק�� ����敊>����z����4/�Ok�'�[��،�o/�/�\6�}�.��}oj�Tb���6�[�Yx�ޘ�2{vj��o<��BZ�z;��7�C�؞ٝ*�����N��Q·llφ�˗�����'=I����^�[^j�*�����P��|�ݣ���$:���Mf���)T�ዲ�6�e7��W�W�ud�9ʄ�w���+)<uy�2��VU�uՖ�5_e���ncm[q�Z�
g��M��e�%M�����?b̾��3ܗGJx_��O�ftCѓ�t�3�i���3k��P��6�b`%��09��\��GO����z_�������!�m�r���}D��M���]��~'�葡��ɤ{�"JY�6��玵�w5C�1�sCo!s�(#�"
ޯ�'?Ep1�2�������1%1�5$��������c��n��<a��s�;-�M�8��-ka^m��O1�X����	Y��V{[s��ڗƺ�:�9�k���r���Tv�����e�]O$2Qх����^h�J��{s�w%�k��2����1L��:�З�Rq�Hg8:��-��V��ZU^���jr�Ny��Ż�Ko�#{���2�s�ʜ��u�,rI�
�����޺]���^�֋�\�)��M m����zƭOW*Gf�jGt�y�;Z�<�F�J����]A���$�z���\i`'�/����l����T���c��D�r�C�s&���0�K��:�*hӢeK5�0:�ި�َK#WbiǷ���2�.�Pﺺ�]Ef9�VUu'��u*iG�Ѻ��T��t�ۮ�p�eF���W�uQ���6��v�Y�P�Ȏ��tu���Օ�Ռ�C�Y��e<����Qr�|$�o��B��c�m�S7^�>�+��2T�e�����n+4�&�_."���[����k]���,:��^�ׯ�L/4e�d!�J�zs-�,C�m�-hw\��I(�뾊�KW@
o+�����Vr�X��_�$��|!�W,��ˠ|�
&��;����;88r]X�=�4Wv�$����c�[V�w;��ED�TT����׷1LG�ܷI|�F�n���⵮�̩�M�a�jҲ����G6q�R̹@�,/��[�&�ZE��$`#�+oFE�r5�pT�Z��.�Z"��jR�� ��� �.�wFre�r]�O�Y��al�l)M�)��[�1�E5�EwnP�t�D�33q,�3!�%�*�z0��-�7qG��0��f=v��!�]j_Yy
�^�u_p%��Ꙧ�0	y�la�t/��6e"�Y57%��3C�י�*=9KnJI��k�o�u�F�M-�d�v1.�54H��������>�b�� K3c)�(-��/ ���������崨�^f�]�q�
�cVgmh�}�� ;���
v'3�]�zI*��_4��̡]�n��U�9R\&+Gc�ʇ�ͽ�]��븓e�����Y����������͚�z���T��T�3��;�r���o�UR��m��Z��F8դ�!Su*�:��eֹψ|.GC]XzN`�df����)�X+��V�{V�b��O�fcYE��@���f.��;��ƧA��')�C{��t]G��������[)ʹ�fEM��39����+�f�hH̜wtT�vu���Հ�TyZW�R�{� M'7��3��j�0`�rE��X6��n����"�A��_6;Kci$�m�R�eK%��H��J��OIk����]��r��f��'])qK�	�1�p�֒qe��X)����ԭ
���RL\�P�p.��W�{�኶��h���ٸ�\p}5�n�;�v��ջ{C�.�;��z��uؚl>�k-ݺձ�J޻�C�ᗖFU���+Ag7:�rt�¹umގ�nwu	I �p�@�,+������@F�8��H���!;S��E9�d�������$D\�b
*��,E�S(�tsu9�!9�Q�D�Ցajk$�D���3���ݓ��Q�e	�W�H���#�������0����E�4eX�RF�I���Ub&Y#&Gs�GNa�)j�U�n$[�M�Gr��PTF�D�%�dk+K�F�ӧ5�Fgj�0
�PG]��<��S��"���+�U$�
,��AuwʏP-=�E�V�t�+2���$�9E\.G)Z�Yt�(��Ủ�TTE^l��b����j�����7�a�W3'�1�����)�E٠��x�ޅv��G��;��p�ܞo;��K�3���(Ry2)�Y�iu?����)��n�~����T��o5o�iJ��OLp·���a%8^]-P�#+6�NeV��Iky��P�I���>�9|��Z���Y
���k ��[�ᩬ�kN�b�5��t�Q�GU��:.�/,R֠.{Y�:գrP]�E/i^{H?K�����!��yQ�p$�/D]r1��|����ַâ�����+}�$~���޶�`���v�M�=�vd���S���5��6��>и��4�n�Υ�!�*hn!�-��SS��z��f����%�k��x���[چҾ�j�{(�.o��wgJy8*yα<�Z�J�No�6*-��*�a<[o�u���*Ǝ���fO���s[�����%eW;�eR�������SsV��އ�z��J�o�8֟>`V��Ɔ^j���?u�;�J|��e��ގ���YQؠ;cX�i��ܖf�S(˼�����ލ6%��R�͢Ҽ�$��i�ž��mGGC4tt�A�)3+�*u�.gsx����<c��9!U �\��7:��7Ԓ�,��6k|0s�;o]&�f^<�f;嗲�O�[�Q�N7��C�@7�]#����Gӂ\:T�d�s��9���L���Q*�¢����O_�H���S{i�j��,��ƥ8��oBH��.���(�u��x`�r�Oosړ��N��Q����	Mt����f*��Ǟ�1=��8�����C+���	��}usǊoW�9�>���+#e�'���fs�� ����w̯�5����=󜎯�<10��{;�s<��c�K#��O���ʋ�e�Mv�ݟ�9p���%YN���ֽ��P@<C ��^m�u�;���'�	�|��iN�i���������F s���w���kF�m�N/=\e�ˮ�J��a�'9����3�V��{#t8N6Z�QX���Ye��o�1~}��t{&�r���ð�%{���Q��\/�q�����`��7(������3��]��"�B�wָ��re>���ܷ(�:P�f�n��WԽ�Ņ�؛Q���|H��]��
=�{`ԫg	�/����\0�<	����;+;:u�ÈQHwb�I�ZFb�����K���� �U���ۋ~�GW>[Ke�ؖ�����M�NWF����9YK��W���=�,Ev�UއӘ�]ϭ4)SWݾL�>
[��o���;=C�pr��s����=vq�Yί�Tb��{�M���y�w�S�Jg|�r��GT��6!��������a��D.�̝$�1?rߏ�{�M�6&�4K�_sճR�+\\�n��ތ��_q��A�j*"�*�T�/�D�3d�h����͟NF'=�s�-���3�
������Vwz����<�8bn35wd�>Li�Բз	&�M����Dm��L%P!)�doTK��r2��՛���则'�r�EuLތosJ��oFO��+�h��b��{�'����Q.n�!Sj)>ɟ��w�\��Um#Nw��'�<�sU[��a�2�v{��gx�0�jxlJב��8&��=�|k�K���x������[�ަ�r媡�4W<�X�9�ߛ�H��ڮ����t�PT׀<7�_'���w�t�{5��Nmˮl,��q�<M�"�ؚ���L�.�n0t����a������mk���J��k,�Y rn��pJ�.��2�r=S���"eW���:�UW�E5����DٷQ�NGz`��	���+r�t��1ڵ͝�T�r��[r�^�f�µ�ii{���YU��֧)��`�!�Ek�4��1FSBتo ]vUe�����z�	���|�[��!u둩ܽ�Ѭu��Wg4#�4v����<^ow�s���zĦ��+o�<|.#�Lc�5�弤�^��?�KD��u��x�+]���m�j5��ūl7kG}�7c�Z�(���=�غ	k�(��~V3*
��*��}x�V(�_ju����C��\db�UҍMR�z�W.ڇ�6��`T7>�s}J��w�T� �)��c��U����_m��m��>ܧ�լ�}��� ���j%EkP��_^�niR�y��kS�#�j���m��i�mlS��W��,��������H��+�Z�1v��\�T���W�u�~�A�G7��5��wm����n��l���Q9@1[�"�]�r\x*�����P���m�n�&�v�-�h�M�-,�}�7�JX�� &%�̋g�>X]����nRX��ۜ�p2b�I�k)>t�X����|��'���^C}6y�hI^����# �`E]����G���o[!V�����:|�|��(�O�-%5c�s ��ӵz�.��Fp!�G�����tb����og�yGЭ�Bď��ս�;�}o>��iz��J~����ّ݅ɵ��{�bY(���]<���bg�57�{��%�wF��B���Ep1+s([�b��.[ڹ�9�ܦ�\�M3��S�q2��jxBc�Y�iih#���n@���	��f7w�(uНI�ش�5�9�3���jhVE��v.�a�����{�T�kJP��Iy�m9�ߩ�.��#�47�˹��^G:{iv��]ٗ~f������ߊ\W�^v'�>��y�=�:��kf:bSX2E����U7I��$������h\w�>}��j>����e{{��4�K���vYn�S��x��ܭl6��8�B�B�����%���Q�iD�@�}�&��3Kdf≃�IcѝX�r���	�Ιu�/;�u�it�Hk����#4���mf�k:�9�#�/"��.λ��F�8�ɧӾ+(��������$H���_,8��ۗ�s�P�}��6e�i���C;�ҭl\�8����g��*��7R�W��tU��J;ls�ܸOW;�챏`�g����y� ]���s��-�˙���c�yTd�W.��&�E��������Gs~&����p2���{���7�I՜O&yaS�c���[��I]�Sٷ8���\�P�t'��pw����#%:R�\@����qݥ��S�_��9i�2t� wضYԽ^
����@��T_җ
���1GM'��t,V<v�F�?g��x��)�\��(weU��n���ve��h�ʥ䖦C����2�,e.���t����7�7U�ѓ����H��Q�-��0m�A+g�����֢&�{�G��kӼ���	�U�[�(��-�:3U�&���}�3��#���3y7��F��i��TBx`u�V�����݌#dȐ�:�ݫb_d�j}��n��N��̨}�b`�.��.��۪�����/�g;�3LH�Y�#��	�v��&:����v�W!�>�2>�}�/�j��B��Izj��Q
�әz�6mچn��p޴b��3���+f5��A�i�;;Ú��:��wyк����L*��5��ּÉ��)&%��S³Y[/��UWO�{�����l��&�F��^gT\���Z�S�]E���M�b�L��&{*���R���X�u��'�E�*�ǵ���5�^n�n�牙]��&3��g��,�rq��wN�����k+����xu>���G�1\NQZ��w$�4�9�*j,|ʳj!<�K����e���F@*vn�/���[�����F&�[�Н��k�5���mĉ��R��wʚ�r�\K�8��:�Q��S��͊��]6�6�p�qWs<iNV󀹩�]޹k>��*���7ޕm�L][p��HM��yN��:�0����m�>�d������4�L ڬ�ڋ�O6�*��s!�8��]ܳ&�ڥ��ݏ�m��njU�ȁc��Pv`�k*�����1���u����oPm>q���лm��.۾8��lo��E�Kބ�m�^m��~7�VM{�JFp��+jdBe*���-�
ձ����fjn^�B`�E6�Od
ZP������Fh� ,Q��;U�i��դ��fB���_��qË��\=�W/o����dMvt�����>e�
����e������[�$�M�Ɲ�r�|)���F��9|ht�V)�Zױ׏��]39����15_[H�9���=��Kcj'4�{�4��+�����r���+]�]�qrw�{��{��$�2�Ҡq��ٺ�[��]���|����+;�/>���g5�����j�cx���/2�9%�O&��l���֧#��2!1�=�+4����]�O{`���Do���{y;ݎӱ�	��O���NS�`g!�Ek�©{#q���{jTO��,U�i��Ţky��<�|�.��#i<�p�c�jt���ĸ8�����M]��7�(������V����pȇ~��s#"�N�.�a)��y���>��v�>}����S�����g�]/���B#���#��'�%ך���W����8U���u_J���7"��Ѧ��yYu;u3sVs�+B�(��ٓ[������b��:�Q*z�:�s�,2��иL��uo5&mB� qܭ/���l#Ƣ��<�����'������wq�#)n�)�SG18�	��/1��Xx�����bgy#��˿���8|�گ9sI���{��Fo^�ݙ��;�M�x��A����/{��^縩��CX��}��� �\7>�P��j��y<�J�Xv�ܓ�t��t�>�O��ޛS9sQ>��	�z,E�N����X�[ꅆ��;�T_%Q���y�DOr5�o{��{ݻ�4Et�%�F8�
6�Fs�鑱�_K�	p���t�zk�J��4�Z����h���W�OOk�P��Q�)TOLs����(�\M���}�)[�3j�d[B��8����-�]#QǊ��L%\o�݅ٓ 7�
�'���)W�w3Jw��9��=���g��[�a9�.��Q���y%:r�KT����+c�*�m�7�S7��Wπ)�R�U�i�%
�\_=܋��;ˆ��)�X{^��yP���&*�P������p09Cw&����e�y��њ�wl��k�]���(=�C���#�N%(��j��؇��J2�c�=�b����Ī_&^m��Y}�=��u4N�ݺ�[)v�v���vi��T^gr��6#{������;�Y�7b+ymO�Y���R�9:�w,�#J�Z�A���y�c��E�'�/1ս3�D�ojmIhV��<��]� �	�,qz��M������a{�s�孋ǹ���Q�Mp��2a�6j�f�c�s=�m;��x��+��f�>}��j>��������ės;^�)/�}-�_��Vr����h\w��k��������r����x��T]�\>1�U�sg��ʹUcYc]�p��]���q�qy!���.��sac/s�oz�YP��j�GvB���:�x��l]3vD�����'q�\�6U+�-6��7�'�O9T�j���ǧ6�#u��z`��T\N�|��A�|���w�ޛ���-�ɍ�q���[�WBʅ
g�]J��
�=Ȯ����q:�7�B*��%�ϣ���\��]�FO��v,.��!%R�~�=_Q�A���H�)�����G؈Tm2�^����,ͷx�U]\�����.�po�X=��<�M�`�Й@;o��nw�\ΜޞYЃ�yVk9acj�Ȧ9�a�E;�\N���'t��Fw�cYf۠�f��s�]��"WƷ�����	Xu\ͭ�/�>�b�D��}\�m*G�ox��|��)��L,�^$+����D]���fo5�Z ފ� 
����E'һ�.V.�bR�:m���_<�n�Skc8�a���P����21;;�kPvʷD�le>	�{f E����õ�(�Re,��J����g:��E�Oь�ᭁ������K�sykdU�f� 9Qfo�F
y����Wr�Y-�
����\B�)�˙�Ӥ�H��=VC=Pv�rq���4��#`)��\�HC��n%pL���n�,�ڝwoM>�N'κ��!g��J�o9����5�� R�5���˷X�uq�r��:mD�Ln�w���)ufngf̓vG�5��ʘ;*�J�S��dUr�63�C:�XsGh��u��w��$;O��Yc�h�i��ŏB!�j��̻�(gC�3�$,�B�\�����x�;�m�Kڈe�x<'{�����{����M�[��Z	���+q��U��7)u�:$�	ؗn��W�e��d�љ̄�,[HpcS�ٹ�2
�WLb����v�G��g6Oc��5��>���U�w�a�*X)(�]i�Ĝk^rZW�I:ocuo#7��u7'k�ҴW`	>1�6��E�;v��ً+�s�${�I��-�F�F�H����txZ�1ԧk5��<�+2�=����ӛu��c�̔"��mRzG%[�خ��`vz�K�Ţ٧b w���c1�/}�{�l�pmh�;�Q���N�7QouNg)�[�@�9@��X����,u�gwh,uL
L��C����R-r���*f+U��B8��gRtR�ՙQ*f�˱G�A�֗{������˧F>�aW�}��"� B�b����\���%K{k^a�5��kw1w�]������P��/�6"樢�@W|�g�O5|�l��&��[r�d5v�AT�0��S�V(��A=��H�b��=���l�;�ϨM�N����*E��͆b����+�����_u9�51u��4�J��X��_-_�������f$]c��{�E����b̔�������]��2�31j*���R��
]�q̝u׬f��F�*�\-N҉o:����H�e-ۋmJY�20v_v����Q]�C\X��w���|�j���w&��}��q 5�8I�Gvv/�'30\�o�T��������W�f���V�����4�V.���o��$K�ᖔ�҅��˽+h]"����sy���3n�_��h3�\�XB""y�fP�,�j�����3}CwX6������s�%ҵ��9,���|�1���Avdq(c+^���l,��,���#����1R�𦧌�T^�ʹ�wO����&�4 ��i
@L���#���V&�d*�*�$8*	դ#!"T-(�A�iP"u���J�E��dkY,��S'u�Q�I��&�\��r�*���IiJU(Ҩ�eWL�;*��Ur)F�h�#Yr�R� �J��+�""��L	2����(�{���ɥ�Q2�"+�D��LNY�����,�Rs5
:�Z���*��Z\/0*����fDȉJ,�f�*�
��Pr%�Q�ʱ]G9�29U��J�I	�fE*�u�!\�E�
��(�*�պҪ���H�QȌ��զ�9�����͐G#�e:�&t"��	Ա�r�TQȢ��, �$N�TEt�U��ι,���"���.p��' �$���r
��<���)D��Ց&A2�M��r�
��R����ð�*R�\��Сù���h��L697�l����Qw�ؓOd ���}��8�kzڇj\Wt��+�}L���:��bј���އ+}��ZH�}��cZ���&�#H��w=0�K��d֕2s\��f+��]�rv�<�y�C9���ƪ�݉E�S�� �������I.]�-��Kחŭ܀�+�[|�[υ�4�Gj���F��6�rjo�=��boWƞձ��gu=�	�%F��6��
7�dgfd�HN�q��b�=0�����g��_c�w�{|�?i��zT����䉉v�m06�t.f��\�am���^b�ǤPT'Z���n9ܮ�Yt�K�X�.'�}Qڥ;�z�>����^@X.�y,�-e|q�e�u�+Ĥc9�����LVf�;�[�S���>�>��f���'���-�zڡ�֍K������2Bl�-����}k�{�5��8��i�z=�����ǁ��|���<d5�H\��u*1^�]�����h��e���,���۪��j0�n,]�^�%�Z����P�ugd��]���v�4�u]�K$��{t���V�h��a<����f*��sՏj��;�[g��>���!��ہ��*pVR=�|��T�΅�˛ʳ1��������F�Bj)~���nM�q��g{��!w�ݜʜ��^ˠ:���ۉ�ԍvb��{�SaN�7���I]ƥA��j*�+���J�in��8R���^4�dS{K�3+��	�?npj�+��}���v���o���p4�8kn!�ڃ��G�r#z;`�җ-B�)Vur܌�921Q�ˌQ�K��M+�ù[ѓ�Iپ幙Z��@�n]�-P�i�m��b�韇>�����M�!|���E��
Ǐ��j��.[��nA��W?F�.(=����!u�rnKZ��ʓX��f�w%C�1��4;�Oa<��ۃ��\�}b������ּ���*k�e���;�㭩/a��u���;�>�e�KD�؜u�gU'�x�oou����vs�����u��)5z!NS��7�����x<Nnk@�z��[Ox1}l��Q �p��S��wW��8��CX,VS��.ٍ�TX郱���a�3��J�N�U���qɦN���p��F�(��.��A�t�G��.i�{yd���;���:]��k�;΢��+flΝ/z"�qvo˝����9e��t&F�R�+�5�S�QJ��Rk2�o+�Wט�������P�J��kGs��ꙩ`���qƹ��y�G��8{�����Ǣ�ڏ�iX�l���%KA�ƌ\39��cU;Y/Պ&~�.
^��-}g*>{�:��x����9�K�ka�K���׹ͩ��Gs~&�����O�����'������.ztj`}�8�]�-���k|��{9s�Q�B`�n�m�z��<*�e�6�a�Z�Z�Rv�ӌ}i���)��*�5`[[�+��!7��(�vf�<��n7+蝃��B���!���;�	7��ݷ	��Ľ5V�L��o���Gg��d��D(sŝ	p���GLRzZiii�gf2�V��5t�g�q�d�M����ܨ��zg����x��T�\���B`�������t�}I%�vY�)l�/�h�61J3 �Œ���X�d���\���k�L��u\��]�{���"[��Qe,�ҁ���I�m�̧q�f�sS3c�|q=�Vn����4�S�vI�3���ڳ��mǸ��p�tC�B�o8�!�G�9>A�n���:E{`.ta)��Z�v�+���i���r�Z�z�����|�[�g4u��¯�a�Q���N,ut�z��T�'�n0�fpsۙ��d,������l�e)�\�c��Ᏺ���!f�:��WM�W�nWփ����v�}�=����O*�7��uw���ا���c��.Ե���M��i�Y�D����t_2;��f=��dC���mIw���Ԣ�Pݯ�\:9��
{h��y?����ug��F�.���T���}!!���*�����^WQoUE����AmF�3��k[+l��M�l_����3c�KWX̢���m^B۫���ѱi�t��HV8���,�l-�jW{�gG�j��P�L��q�L��ޢfL眵�&�{#ʣ��D)�,�ƞ{v�lT[o�U構Kt5���t&6E��YI�	��P�09����VWvwv'v�s1��qь5tqG�N�D�R��AU���+���57�t���b&�[L8�ZS+��{.|
��Oi�vCr}����-������K瀦e_nfati��qΔ�ell��mu���ݛ���Ч�Cr\�j�'�]aj*-��7�*�A{K�Wi�s1��w��,냳�k�}*�1Q|��O�K�0&��w�Sn5~l��19���
�W�n)�����A�K�}|�@�}P��ݍU�-۝�ﻕ\Ҹp�+��Ct�j
﷮J�\�q�/�+c��X�.�x���GOԻ�)}֘�V�d�N��Q��눷=S\���wk��Z���u�e�&��j9�'��9�\C��Ќ��34�۽����8�yN�71\%k��-n�@[�ɭ���;g9�z�]���[O�]��5��O��11�8I{�im[%vOn�ܢ����7mH;0R���e��u���������^�3��T�w�~��Sh�����C�=r8QH޻�.��m��C���MC�S���'��lO>����=���(���rKzV�b�}Y&W��d|�z�����QR��"�n�eã�����ݩ����f�eρ;W!�yH��)���7������u���3�W>#�|���5}�1��QkZ�R� ��GsN7��Q���MO^o�4�l�anwvOO{ך�<�_s��^��Z��@̺���ծ\�eB᣾7ߧ�]�/iX�.�>�=mE�x�s���zi�F)y�i��"h�泦E�u�9�ns9F=ǫ
l\:�	���h�-lv�R}��h����ʂ��ʹ��c�J�W�u�&��:�az5����%�{&,P�)�k��GU��
���/�TY��g�y����jmnӺ���	y���;��~�邻���z
�%E��P���s#�������F�;��qӪ��w����)�F�omA郱�Of�7��*X�:�^Ew�Yލ�h����"��^�c�W�лZ��:�L�G[����V��=����c�����r?.��e4��޵���#����^��1�D�x)��Jk�G>�\���]żr]}^̰�Jн^>�0M:Wdע�a�H�%b_b�f�0�@��j�F1<u-�vJ�o�����.n�=~�~۹��pjԵM끞���
�I�6��2դu�!��{t���6���Z��P�o貹fk^� N��,���w�� ����9�����/��)�ױ8�w���~��:z2��"+��V���z91�
U�F��B�*�����5	p�O!S�3�c���!nS�$F���D�X�'�Z�V�r��r�l����NGTBxBc�|^𕲦69#=U=T�V!Κf�{T֧��Yˍ�m�P��T�`�&�5w����CN�r�/8����p'��o'I��!u둵	�<��]4[������ݓ��wLˌ�ی���iK���j��7o-hO�K��(�͌�
޴��E���wR��t�	��G�iX�����]Yy��'�`G�N��v�]�E%������\խ�m-}tQ_9�w�]kѾ��9(*Jw{(�����{<��6�|��mZ��w{�c�����e�xlط)��e��ve��k�eW�rw��[roq����m5�nm�U	�a�Z9�����_h�,����3N���4����k)��ۮ�p�+�R�r�;��K�뙫���-y���|���!�R���t�?���ٚ���Se𺷸�>Y{r�-N�y��'}W��7n��1�7���˝z&��u	|�p��v<NrV8�8���}�;�.���kr6�)���{�n�_bˎ��̾yz�
�P�{��ި���b��*�A�7��5��;�LG��{����e:ч���Xx���R�`%��Ź��'�j_������]vm���� �dk�r�
g�o*%*��}P���qoUr�;T�'�����ݝ!�9|j�������O�s��	LEt��^�
0���=yS6�v�/��\�J��s���֓�yw���-�n���Q��-�.���]�É����g�\�ʆ�����S����扷K.��N��od�a�u*5�V�3ڵ�|ʍN�Zc2�ҽ�tn��eM|"�{�u����)1�G�TA��y����Z'cy:n�rŎc�j~\[�C�{o��{9o�_+����e=�R�����w���nvIX��������3}j���)<�����N�-Ɔ��x�b�:���tX��9��3�]�-h���-.�k΍z�3�vR_𒷒�$��S�b��{>�VS�OnCu�N�t��}C�.m�H��ǽ�Q]C A���qԢ�2b�Wr;^p�by�\3�STk�ektW`�YoR��������+�j3 �Ƶb6��(ؾ����.�q֜��eu���
���|�t�Fu{<g9���&5�����5w�z|cj����UyK{l4�s[ê3�S�~�sk:e]����/����z���qZT��y'�*�d|u*t��f���Mɣ���V�r�x��ƞv�^��|+[kެ�F\8�B��5]���S9s_y?CT�L�mgP�<*�*�I�μ��Yh��v�u��vZ�g�5�"�rt!�?@�����t�:���Xw9�Y�3g)�W�{��C�O]�Ҹzm�ђ�7�����5;K�7$kޥ9I괥��1uL�����P�qt8����9��Tn[���g�sh�Wt�W�5�[3*���C�O�z��}]�P�sY�eN7̏gH�����j�ZУ�Huk��ek��gk��I�>�L����W�n������V��͗ZՈ�7!&e��g�{���J8d��k�Cٱ�F�5����r���$��@�j�v/8U���+��l�\�7�U�᦯\+8O�ꑱG�!#e�o o�2u_t:�P�}c��D��0��"bb�W��)�[	w�xe'^E��y�I���3j�����>�MWo�'}�e��Е���'�%��麇�<lSU�mt�����D���O���2��6VMC�g*�r�,sZ<-�=;�`O{^�eE�Q��:�{ί3͍���)���MSG>�;5�9�F���	G���&�^�Y�;M���"z8�[�U�:�,O�ϥ����&��_�D6��޹��@���Ɵ��=$���VQ4���M_W승��ЎK�%iXtN��y�]L
�O}� k���9
u����dM���.��ْ�n�>2��1v�!���v�2�,��fP�[��c�ܧ�\[�n�x��avN;2�<L�r�_��ӟ�?ۻhM������k�ܪ�k�j׾�I�z�3�Ќ���9��g�������^߸��3õ:���ΐ�~���̒�ϑ�3������ig��C�ݦ��`���^-s:�!�fa8����l�ؿ_���W��ޠ��[�9��X��
 *Ysz=����ۑ��bP^�Y� B�I�ƽ#F��J�ߝK�3�T"{�~�*ۛ3]�4ȫ�ʍ�vS�[��>����d\�Ahn�^-���36�/��#Zm�V́0�+�k�	�6�����1j�B�H6U�}�Yj�ok���ծ��TG=��篝���@�̷B�-��^�6���w������,ʺ�>�Im�Gu����uzV�y^�Go�N��u<ˏ.�7S`�pm�B��a�*7���O�S��z�jp�Φ��M@�Q�u0_u�ok�}0p�=��.9[Տ����fĺ��?�%�{vU̪n��tu�u�QJ���8�R���+ju�x�)�n��J�7t��g�!��4v�vp�z����O��c8�_�\�Rkq��5;p�+�KlmgI��&S�������ἥlZx�l̥����-��W���i��m*ɖ�O����(���V��N�8tԻ���_t̩Kyp�+�B�|��Z ι�L��-pݖ[�u:�9rR"�Nې���3�l����+�*��!`2t��·C���c�Y�JM�n�]X������V�V�e3R�\�P�	���N�,���:|U��B�jE*o6��kX������jS!�@�ɉ8l���`���>�S�ow�=���X�7�֝�6֡/�pL�;�Зn���R�����֞%�oh�����@��
��%dv�d��; �4���7�2rE3�>8z��l�ꇝMS5 ��n�7�7��W�ɠY�)�Z6s}/��[N+� �����v�51�u�<��zk�#�0&�GN�oW:5��f��Z�±�,#u�N_r]*ؽ�|o8I-oo	���޻��v8�䫫���-���pYU)ż���������W�"����|��[�C����0��]wu�#\�SM��Ԁ٭��O�im�l�j����E�@�*�L�3����Q���éy��: ,�8�Y��������aG��<����j�@����eax�%L�  DPz��R�9�x�a�����goo���1��Z�F\q��͘�����Z3�ullm�ZO(�<T���:�ٙ���ࠫ!��!*۝4��P��Msv2�P��A�!�p��Ҳ�{[��<.�HoʗX����Bw[��#-��PR����R[I��!��JЇ7�g9�;9Uy�Fn�j�^{��4�t�#v>��.4�n�5k��u&�"��N��U�k��v�K�1�qU�����.�%�(�E,竔S�+2m������"a��������vmۂ�gL��Ou=ڳl�-�k��0@t���&�M:��[���-��:��r$3��mM���.E2���f7Y��#Y���i�:�+{{���nlL������OW���A�:�h�t�!J����0TPu�\GN-:�{v���SC�`��4\=\�cYNCx�<�;"� �g�����Wdf"i5��vL��^��������q
͢�s���Ȋf���%E��Na�"�+��eRq"�
(#:D&p͜��':���J�SZr���Z��A��UP\��L�3(�U��!K��r��r�ʈ�b�Tb�Ή'���W9r+�İ�@�W �'2�P�B*��z��!#��IQDTvUU:,���瓑�S��vA��ATEՉh';�ʧ6.㜢�"��B��,�T���UTQ\�&GuL�
&'K��U�(b�XUE���%J���WP�e��EA�����
�!'$�I���&ȹ&f��'
 ��r�r�S��3aAfTRKx!H��%Ih�uwxC�ù��$��G��(�I�@�i\(���*�I�Y�UQQ��d&Bw�p�9r�2�׎����fdQp�_x��GţDus̢�W�r���.Ds�g.�+����갓���K����FLr��3x��ֱK�&�u�X�|�I�g&�ұo�m�掝..��[��Zy���t^�3�lO�s�9]ڰ�����|7��1��f}�s�\&u�Ы���k�pzK:��5b�C%�P��9���3�lz��d��o�wD+��h{"�71���;����Әi[��뮘�9[f�r�>|�Jܭ����x�ǤW�D�Q8σ�t5������'��jn3��Kف���.�/����3��+R.�&���Q��
�,8KGّ���z����A��#fPg^Kŝ'm��^G���s�$k�i`�*�@^5��14���"	h���r`�9�V�Y[�w�y�>����t��Y�@������ݹ�%_L�ȘuzH����G��~��8j��QMfmn>�-��/�<�Gs
�ڦ.����6}��樁<�&	��a~�Ǘ�Oݧ��G(��{���!�Zd-�ר�����q���/���PnfG�d :*�@�WړF�/�)��n�	蛤�mhw�N�I��v���Lz��/·���Q�!׳���(Zr2J���\^�ow���R,Ec��CЪ
��_\�;ց���K�5���z�7̋��5�"2�c<3�[�kb�e�������,.�����M�����.�j	3��!0�ov<zou��4u`�]��u�h3U����E�i��D>���Z�1��y;2�7���#��ً�e7��7ðl�ݐlwΘ}��`�+@0]�����nã{�����y0??m��9�yj�޻5?`�h�Ђ1�[Ɏ�M�\}��ʣ��=R7\{��5�C}�� {���NC:�=�cGw�\��'�p�,_�\Qc++n:2���7:|��޷�e��.9�3��0*پ�����Z��=Dh��O��G�FUh�4A����^O�k�VJg�j�u�9�^��x�x1�cP��f������(��{�)�I5����c��|Q4l�~���/�����3�E�^�n_i_S/A.=�}��D�--[���ʵ>�pQ������'40*��p�o�Yz�}k�O��
w��纟N��-�C}�ǅ���C��k�xW5�1P[�M����hx����,����@k>x�/������dh����d�HVJz����Q:g�s��_��s.Zuv٭�W4�i����T^o�G9�ū�Y�xJ�Ӭ�T�`��o�Ù���Mg�_��WʐG���}���xw�F�i�+�}���V�l��h��y>�SJ��#@�o#Nj���8(�)��*,^��g?o����Xl��/>�	yF,��"Ԗ�Q v�3 �ޠ)��Z�X*Z�`::R�t�˫�k���c�9���Qˌ�.��K�vиk�N]�RXÛv��3l�H]�q�M-���+|�7�К+L�f�J�\.��:�O��߲�\ߎp�F���{�!Y��F[s�LS�̚�9ԯ{��,Č��oq:�q�	[�38g��~#4m�yW,��iDN�Ny��u��d࿛�eM�EI�n�>}5�8�Ut�)�V�����"�1=�����mE�B:���H�\s����?>VwV!%s}�T�����w�T46���uC���DV�K9s,v�Aڅ�q���ԼT��+[�ꥌ۬ �ή��1��?^���E��	�wT|�Ȱ����=|�Ǟ�o7gޛz	�ʚ"M���q�!���=礭�1]N���D�>ҽ}Q-�8W7m���h:�(d\�^�k���箬�Qe�T)��f��ڹ��߭������k[Pl�ӰC���ۍS���pǻ�'��b��9�2�z���B���^m;�j��`z~��ŚfgqE�=}�g�䥊;a�r1y�R7%�=U0�ަ/��ʙ1���z�{������Ǩ�8����-憻g�b�r��z�|����t��桁\���aL��O�s�}/mƛ��l�g(�J�b�iIX�r���8�'_�7����e� ����x�H �ϫz��(,hAu�5s3srsZ8p�smq�(��;�����xR�+t^,R�h*��]���m��z�,̹�;q�Z"w��9αC0j�/]Y�In��A�O:��Z
�{G;��r�[��3��3U �鸧 >E]�����ؽ�슥���Ձ;�)�Zu�\�a�{����p�������%����}�la��4=9wU��4]�J����
�������k�n&�z�1�ߋ��{M��H�P�%z����f{�="|�����s�mO����lX];�/���=���3��b�7��_w�]�n���&=����Li�: �����k��t3�-�.{G��ޗ�<��ͷ�%*g�/oܜ��E��8���g>n�~���<
���\�C�[�=��V��7^��8�<D��(��φ�yح�׍ǧ��>SZ���)9<MD��3a��ʄ��׫raf��˜�䜐��:��ho:��V����=�|�n���j!zJ9s,v�75�۸8ڸ�e���:�>�^ڲ�Fa�E}���CO��̆x����uP��8kQ�OQ��3C=uu-�F/߮�i���;Le�~�����u��g>]Lw�`���h��o��鬐�;=�ن��Y+2ѹ����NlJ<�v�k+����k������_qܮG����<�.�>�~�uΕ"�̿h�iW�pOn+��!�j&�f����D�B�HUӹ[�*�5�	y�΅�_L����Wnm)�+�$��vʫ�\����-�/*s�7�{�t{��Y��2����`_�'�=��K5����0*�˹��_��n�`xL�b�[B�����f	w�<�xu�4\{�uŬ�n$�>YP��V?	V�~3���M�_]M��L�3�̼���ʑ>����v۽����v��$�7��0��Qcت�����\�/��G�i�qRy^j}�q���.3�c*!�����*~>]���B��VǑ(��z��W��Lȕ��)��y�=������,^��㎼�=��ONF�[-	a�:�w��Hᙾ�RĈ�o-+�D�V��&��:%ɳ�#j���'��U���a���;�x�wb�g�j�u�˹�7�bb>�i,��;��F9�{��mW	ߝ��Q����]1o2��c�Q�8=ܧ�#<��Cq���\LL7Qt��A^��"	h�5׃���؋�pK�W�&��U�M����'����z��7�3�R�0,�\�	���1=��궉^�MU�!/n�3k�'�b�o����a�;��:��n܇�Q;����:gU1�����޵yOb��#ɺ��Z.�0��#�11�y]Щ �2q<K�u[X�l��#�7F��	fFR�8��7q^�iV+F�S�`;Z�	K����3rW.�͕���t��N��6��G�e����,<^�TD����w��^
+] �Ĥ���X�G�}<�o�ޥ�����L:���bӞ�y�fϽ�H�800M(�]~��T�lV�mMR׎����S�UjG�h���Μrox�ν1yŉ1�s���}*�7���G�,��#��B�)�h�6��mA�~ڋ)��'G��ۮ����ǳ�V</��طۜ��]Jʮ{�5�e_��"�EF?�q%��f�+t�y�Zs\�_Gm�d<�=�sf���һ�҅vz��`\�u}�˱"���Z;��I�)ڇ��=����~9Cc*��Y˩�=n�q�~�g�� g{=~'����;ס��*���Eh��IӤ�~S�E���Ӟ�;@[�����e�8͗A���Ϊ6�\�lW�~���]���M%�����{y��Fllݳ�g}�}5�QJ������e�:x/q�cp&��
+�z����^��]
���{�%�(��_�~��w���1q�{κ]W�Ǒ��9�}�������+9�X�f|4ۭ�ʅor��PN�8}�u3��a77��Z�y	pSOΌ�d�˹��Y����=͛m� Lx�u�o�*���gG(���5��V�o)띓�X�V���kkEEd�OcWI�yז+b��f9��儑��8�࡜��z�l�wLr�p,��c��}�̓��޶��\��D:�_�~zOm�	�n�^�î��.Sw;�Q��·�m:#}=q�jx;�ȇ!���r��Q���H���/R�����gs.{�+�@���:�[g�<��%��C��ӧ���ܽ>Ix�ɏX����ۋoɯ�5���������'�׭#��ԁg=�xTE��ȿ�˒�ax����i���.!��s�:�=S>�u����jF�i�7�u���"�c��O��ң���H*��M�������'I��|ϯ�A�Z�)�Ӏs�i�΍��n6���b�<�ٵaA0�+g��v������&��Q${�ٺ�ו�X���u�s�=�>z��d伮p��r�յ�������6�OM� zITox튂;��Lv�\�#�"��	t��嫛��d�S@�U^m'~�8�;�s%��Du�/m�����(�����S�ZS}˝ۇ>�\�gUJ���\ޟW�L�u0�~��N�����r6��W݄X��BD���]�c\�qҜ󋩞���ƽ���ueJ5�ncH����v�l_t<��A���6>�~��x�UI�꠫��+/� ����|�N��\�s�@���ޔ��ٶb��:��T�: �v��3"��}b{�:Z���Kz�ӆ�T���sI-�3�����xH:��l�խ{��[��dԭ������җ��Ǝ`.Q��\���C���I��yh�α$T��+u��EV�l+,(w��};8:�k�.2kJ��htm:	���^��k��Qf�j�_쌤��8��Y7��3v�ˎiJ�~) ��(yFMib�g|n6� �}T7����}|ǔ{·>���oZ��pYkE��C���vyu�c,�[L1}�b��W�f7��t͖�����j���w��=e�R;�ܻ��yߙ�C���M���D��ʑ���]i��M��ut�z�൓0�8r�����<�p7ض9߇���ϡN�g��D�w�z^�ɜ��%
�.�g,�y��;�h��&����C�{�s�v��s��/ސ8n���ՑP�^WdR�����A�GF�uP�e��] �-��7�i��3�$g����r��G�Ҫ�B{��F�{�o��x�Th��Ws�Yg�/⧰�gu �JN�y�{�������8������쪌��H���������.�14������:3��C��UVY�Kk.r�;.��?����N�Ϧp��� �P;/�����	��c�?&��8�
��֏�Y�W�������$�AV��V����2W$9QBhh�&�V����S�l뎊�$���|3.�z�����ϙ�s���bs��m��Yi�5���UqZcu�쾩�ѐ�X��w���yQqaRv/�?Dy�yz��K��s2�3��7|ey���,�]�t�����A�U������B�M5��C��<C�#�:���x+�u��^�(��<�Gζ�=��j�����ʄ��&^n	ֳ�3����co��^겷f�j1b�m]C��T8�	� c�UCY�3�˯H�m��^�;�Ο~>Eiϧ�Ɲ���'��dΊñ��8~�}w������~^�`с��<X_j��2n&���8�{P^܋���QB��c0Δ:#=5��S�;���{@�I���2B����g����Bw;�\m;���$=C�:	�7^,��xk+i�������Ջ!`��^����u������W���n1��]������hp�.��d���,���X���'!bv2 =붨�ku��~��dm��g:��e�:�	��b�O��=}K������p8C�ڄ��׶zs|��3��@���o�)�.5�?�N��/����l�9L�v���Ø���|�c���f�A� �t��謁'�r�M�ٸ�wD+�Oև�)�s��q	B4<��}�x�:'���pv-Z��6�{�������wt1vZ���a}�U�N�\Ù89Jn��B��Ժ��yσ��7�c��V'ս@)�����S6�;�����]�QWQ���=V���^d�9wlE9<x~F}ʶ`c
�Ek�A��vF���ou���}9��<v��g�H��Q�%���|�(�t�Ư|}�,��D9,�Tv֜�=�T��YZ���>�ya�j�!)��L7WJ�W�z�>�W��+
����}��+�H�>W�"�u$s�����ds7�6)�[ /�&4�{�#@\�+���n�s�m:��BO�lLsݶ3��y'#ϩ���@�ʈ����$��1�S㾚N��]+��]��h�:uI�����
C����S�HG!��
��nI���ǳ75:��<@��~~bN{֤{��@�cs���Η�uꋨ�-Q��|��O���z/Y�դ�f��=��� ��:������Ray��B]9�5�]�����5J����v��Ŕ�Z�ҧ��l��Q�M�d�p����$4sgj�2�K�l֜�>CR�ڜ��Jt�䜼oo� �FrՈl?my�)��_�0HǢpw��(�਩��os�S�اf�rU#jO�{ʀ�d.� �~���N��D/^���r.!���p�N�%����2'�B�����hˮIBGm������z��q�]����>�Nm]�Rv0=vEqY[�x_;�8Rt�	�ʉ��\o��+rtck��wRJ(��.��
ɶn�|����uw��ʽ�gw�a1��x���K�Lk8���e�e��jֹB�k��:;�ޅp�6���~�f�Y�^D�v�Fuhf��}*�eC��A]����I��W���,t�ĂwǪ�ܾ5�H��H����[�q���7A�u,W���1���c�ʵ�oq�s��9�5r,&�<o��9̃ۼ�^P=�+F؏��2x=���>����u�pAf��2�wm��u:Y1T��V�����G�&'�����I�'�
4���2�$���:<7�F��V�����5�,AWZ�xэՄ���U/{:���bđ�Xq]t� ��鮮��J�˶�6���]��1I���ӳ@Gѵ��HWn���-Ŏ�,�i4��kF�Ј�����
��e�4����Iq�rvۇ42��}���tw�5u̔7c�z����2��S.��2��}��e������N 2u0uաy�L&��ҕ�ʹ;D�P�WV���NYzt���C���[�j�܎c�N�$삫ufH�S@�*�â7��E)��d���r��"6��`c'l�V�ArZ�ϒ��=<.��_t�j��`tǰ��2cB�(�{��3K��Mv���O��)[=���/4U��2�
T�Cf�śLf軑�ò��_5$�2*|̹�s�Olo%��f+Ǎ�h�j�{��� ��.ռ7Ζ��BG\���᮫s$�s^�}�Y�� I]]����M�P�c� =��g<��s�|�Pz	$�K� Ɏ���/Z�J��+d���ڙ��U��,�_e�**TDt=F�2�jl7Q��0#�p72�9�S��b�s�7��S(SL3z��M���ꔅ��HB�ߓM�lr}�.4J3^���Ls�8n��]����V��]f+��;!���¼aCu��E����7MM�h=�z�tE�V�7:w���*��F�Jּ�K�v:���(LۙQ�k��&�8��̡���1�dH%n"�F���'�*sG46��SV�|��q(���軤a�@�KW���djg�k��`�5�{�f���{��,s}C xL+Vp(��cf	� ��w
1��͙��wT9�����E7X��������V-L��� )f�\n�3o����g�k���yT̂3�Zp���Ŗ�,��>��Szv�fZ]^��De�2����;J�l��r�������L|��3)^0�a+�/��J��oZ�F���k`YZ����9kl�j�򀚌���9�5;Ͽ~|�q�aȢ��(�Ȓ������Ч'tU$����*D�EDG ��*��H��.Q9F��G*N��e��ZX�&m�"��t��eM;%.�UQ|R�]�л�E�B���U�E�\����ɭ:p�'2��ͪȈ�3�vU\("#�ΞdG�Y�Ç �͑\� �s�>̅U"�=�(�j�p��e:�d&:,�5��׈	S��MD��I�|Vz�P�\�r�2(.��i�aQA�d,�����bĪ�Va������(����e�G0*/��T��'��E	�E��x�TG<�g��Z䔭�Ĉ(.r����g�(�"�RlՅ&���R�!L��s�$�T"�����W
�<�TDUu (� 

���p����ظ1�ݛ4]�zd�yt�=���h�-�I�[R��M��Jt�A�8��R,�b���@z֪I�wV_t7��}���v���'!�.���`tG')��n����U���m.������Be�����gZ�~Q2�צ|Ւ�~RN�ܞ��^��L�7��X,F�������Np"�N)����)�B����+H�J���s�,^)~7���G��G���:7ü�U�Yxq���޵ͅ~|��[tQ��j��j�1ב3ƥH눪`Q�|�ï�a�}wx�>(^[�w&�r�S:<SW�5Ĥy�}���CM���
B��'�����n�>�� i�9y�է����7�<���|����3ܛ�#E}���H�Gt���	�q�J�_T?V#t����9����V{��a���[J�o�^��?J	��	�Q���ϫ��4���S��\rn�L��2���g�7����/��*����~ _���|��K�޸�;�c���Fq��8~!��0c�`:S���\h�_}��ge��vǽ��{���^ʚ���K�����t|�804	����Lv(�d�q�=�|=Ч���4�w���mA�&ѓ�sF�:�gZ�5�](P��:̽�y+8��wX�{|��b�N�-�Z[���
L�����<zJ�6-]6�uh��PMHJ�b����"�'Z�N:���J{Z8\|:�Z��y��h���6;�GA�Ù<œ.�����9F}���	[�-�E#]�)�)4=�Ub�kv<�bv@�@��{�=0`bLv+��mE��.�`�5I;]�dy��!���RW�����2|z>~u��Cà�E|�%��X�3Ư�f����^�+74�N#�{,;��P�=����̎�1���]��b��Q����o�g�<*�Mg�j'K�f6h������LF�t�p���Tc>Ba;ʃ��>�S��\{n��fx��X��C���g=�K��Y�6����oz|���9Ͻ���O�٭���Y����e��T���:m���x�`����^yQ3�s��C�QJb�OLr�3�*�麆��
����ٞ����^�!�������w��l���nJ�z��b����γ�� �4|����ekv�\b|z��\�ul��)������~�J�ՠ�4|3T���r��$ǚ�}7j���jv5ׯF��1�T:�\<�<��W��7���J�.�^D9yU��2�*�C�j�Ãe׫+R�h�8@�7^�%x��u�O�q�s��p�����v���J�)��>,�[��5���P��0�<������������N)R�7���,���?��>�8s2��Τ4C�rn�j��zT���!,[�ɱ���QL)u��yl�]Wi؈t��lbM���ۤ6���WڮM�R��Zcj`��-ޅ����} ���0���P��q7�J�܍n�w��_�#
���*�0��Ϧ6N{leRj�o.=�C��0��8t)\��uJ�|O�Y���s#U1�}]���\�צ<;���m��Γ�!�N6�ηU��<'}@v#\�3�얅Ɠ�I��[��M��l���Ȼ]��O�\���P5�~���b��$�V��>7�b�qK>�Y�+�.̫�{��C����<�/��s~�fYQ�@yc���h�NO_L�ދ�}1�[-��U��O��g���c��ά�_ ����9��;��Yȇ�P����XyD����Q�j���=w�I`C�e��_�
4{�_Z��VS�G��M-=�_6���$q�lc>�6yF��sJ-Bs���ҳqU���g��+嵐�%�ld����'Ei�ݧ�Ζ��� Ǝݡ���3*�gr<S�}�Z���~ڃQ�ى��@{�Z*b�(�7�l�z}�}�wA�G+���α��e���H�/e.'�Gw���ϴTW����/�fk�O��C�g[���/�2�n��k{yӠ��E�lP�y��u^��V�pJ�gr�vg3�1���&4��U�nb�P.�w_\jk/1��~��]��_(UǛ2�z�/�r���a������u�~H��(�1�����f�c7|��D6f�]EBf��滧t��k�v�?����E�P{�X7��q��B���Q�]0�>�fn]b����W�9�az9�GTY)���Lk��P���`L65u:������o$h�r��du��u��id.pU�	�����_ծ�<����b��:�-u�(c�v�)���:�Os���}�V�y��U�pOO�tIR;��&(�Qs�#q�����C���+�1�(c�1tw��Ӿ��SB�o��|��7��Ǳ��[�٨= r���"@�X~ۨ��{8�hn��k	��{;;�#ўn�����N��wa�j�J}s0�EңW�a�D.��e��ǖ��X�E��~���}ş"����=�G
�]�3�@Z|�dƼ���S���G����^��:F%=b� �	F��7���QP�N�pʝ����b {#v�T28�D��)&,edmN�,y������)���,��y���t��bc)���%�ཕ>��gb�-,��3ա�/h0a{'�2��܏l����{�Bs��?X�ˆ���:�(�%~�=�>�W�;&�F�hQ�5�me��[O-�.�q0N�aj��j�@Xk��o�P����4_#w)]�R=�wx������݆�Yw�P��{�Ё���b��JR��`�)4�ZeE�෹K�����fJ��-�p�ɻ���e���Q�V�y?���x���u�K����1i�)GZ�=_Y~dL%ӞQ�]�M�r��m�Q�s�.�b�+=��Rh��n��zI��Ш#�**c]�b�e�MU��XF&�c�ϳc�eާ7^�g������ᐽ-}�i�.ď<�c�'��ˈ��xK��wy��a`���r�КUZ���K��Z�����.>�1���+�ץz�l�X�U/ W'>��BuNu�塐�SSu
���|�９�����.t����ј��f��Zڊ��s�B�|�s�Yˣ\����!鸞���V�LQ6�z�YuGE�c3쯷�?W֜���� h\n@�U�e�,�p?�YP�#�j����{j�s�,^㊥Щ݇3�O"����������ۃ|�l��e�;yP���C�m�'D�O��0'�G��aL����B�����\��j�Kָ���߫�q�/\8�W/�î���RE־uӐ��o�I�{t�μ���LS��x2�v��2���'Q�W<�|�p�y��2��/O:u�$��Gt��%{bD͏�arD�vf�ࡈ�Wr�O����6��3}Y�\]p�7x�s�er�(h����~w+��Cxy�Vw����T��7n�޹[�gl�s'�"�t����-���:0&wM&Rs�����.a�w�6b$q��um�����+W��u��L9c�=E�0�Gb��f����譚��-f�����W|����,ﳃ�?g�����F�V~�<N������>!G�4?���ma>���w��{P����}��s��[%`�f�����3�n�7�K3�6�T�B���I�蘘���4������ȮF'���kg�,:#4b���㽯f<�u�3����>�����O�wc�\� ��&;UxyW�W�ˑj�5s��姪��)ǃMI���V.�)�[@z�{(�+�������C���0��������3�F�I�n�nU%��䇜w�q�??s��s#EG71��Uy�bR=����-ٲ�-(3�~>� ��O����˲�_ٴ��oKD���q�Sy��^�,�_w�n���C+��xa3So���-�J��t�{���\�d�v�S9Xz���1|4
�g�=;!�u�~��lgMָ>kl���(�{;Le�֕q>*#7�ɛ�s�m.t�8���,��!X��u�*�`L�ho�f��1��/.FͿ�^yQ;�6e�E��G�rwl3�_�Ƙ<��;=�V+j��N��pR�lV�f+�j(As�V�����{+�{>7ʱJ���1�ޮX�XyX����-=�:�
��,U�E#�L��ݭT��cU���7����u�+�;��i܃H��Ǎ�]]Xz&u��*�|3�ަ��Ƽ�3�y��o��[v�������T��Þ~����3�nA���1�L�:�=B+�NZܾ����Ǯ��ͯU !���/��Y!�t#�ږ��<����w���:���=;�j���p�x���OQg��k��M������%���pɸ��'�~��x���f�y\{�#q���s�t��W��A���T�xk�)�L�.�<�fO��|T�&�P���k�E�p[�$a=��+�p����הqM��#Ȝ5Ԫ=��B���n�I���!��L{@L�aYu��]�<��ە�̵�˞�����mE��"�,��/����ꋤLO������֡G�w&���{�N<����_��9ٯ�C�h
��r@��ve�W0��"4�S�o���-�w�py)�������0Wؗ�������uJ���"����ǳ}�g:J:���ur�S�-`׳�эȊr�������[�����(�?:��:۸�\+ۥP���=C�r�HrɌڴ�Kݺ�>5���X)t���T(��w�i�Uq��r�p��wbi�QýA���	�^���$��ݲk��l�tބ5K��=�Kfr��"�{���A^n���q3}��3L8�N��>�`k��+�v$lx�qn���n&�\Fmhw;���7+��{3!�rwg��]ٝ C5���VOK��A��#�v��\wQ��~e�嵐�%��?���'Ei��_���`,��W^W��;8����e,�J�7� {�յ���&��/�������GhULT�ho�ٔh��Y��N_���G�j��q��n0�w����g4
���oeZ1��T+�Hv}�0��!L�8���^�]�~�!�][Nü)K�yu�gS�5��Nx�9�u���myp�2�E���=1a���թ��r�`ҧ�PU�Ւ���S¢2z�ps�t=-��a���ر��Hr�z���ۭ|���C����%����>k}h��|.#]O1Řql��g�v����zIJ6�f����9���Jw��{Q_v�2��ҍOH�3�+��^W�F����~�<�r|F�oÍ5�X��;�3�8��^���Z9E��3G�WU�4Ke��Z]��O�O˪�%�sܳ<y�lH��{���!+���o����¯�	O�f��Tc~�v�(�Y&s1F׎�2�V�3.�5Y7y]<ռ��#���A;N��A�ھ��lKdUG�[�t6�;ltmF& �ċ�\!��>]������.�k���6��Q3n��;[7W_]���ǰ��9ʉ��o��o��/g��6�/��J߬��ډ�s���	�^dky��H�s�H����/#�Y!���P��,��W��@.��<5�Sw9�]�-�-��J����~=����N�l����Y�{�T|�e��S�ջH�N{tW��LWH���a�3q
��*2�̱P�����x-|��K��Mt���~�8\��1�@�0/d�fw�����@�w:q������x��俰���+O*��R���ï�+�j��9���Q&�Oa�/��&�:����̌��s�q������ʟY"�ڪR�v��c��^������Oά{ <dS��t1�Uߢ�5*/��#������Y䗱��}���Y���^���H�?eؑ~z+E�ޓ����Z��9yf=-l������?�rc��S(W���yuxn�L�G�:�9K�.#��!��w�L����Ur(S�^�Y[��f&��R>	��eQ�4��=��|�_��&ѶsS��,��zRE��'O!泦���ͼ�����=qT��&����K�U��GW��b~�sc@��"�t�*7��l����0��S���fR�{𸸥�e�9�;\R�3�+y9�������[���QN*Τ�ٜ�O6�6�;��Sm��(FD;�z�}�[+#�O슞��f�[o�$e�Ku��rsC�L]t�vֳ؆���=��fe�/-�;�"(� ��p��3է���S�n{^Go�� ${�(��`M�x�x_�b�A慒eB�W9�޻5w�J��ƹ|3��|*%��A�ʅq�(p��PN���c'��3C{���7*o�Ӊ]V`ڻI�9�o6�9�z��;Ѿ������yp��Nq��U�x��J�7Ef<�>�9x�kB=���+��%�Ѱ���\kr�B��,�:@��W��NI��o�cc.�Y;�-B�v��m�ğ$*'�G9�U����T{D�m+��^��|�(&s�'�>}��X��^���8� z:Y.��'7��a�Z��h�G���<��ݨ5���\�=ҕH~���Vnv����O��Yo�����L��"�$�U�L/�t���s�:2
s�1{���|.�v$����ݪve�SS;L��S��rT{j9�>��`hv�S�r���*BVǶ=����&2��Z�7}�X��=��^9��9�a�r-����P����K�J�{B���n�s�ް�PR��}"7��!#�]�w��ޣ>�E���yg�v�xg���F�"=�hR���~t�y_	��5���at2�d��̺��s��r��k2F��/Ek������>S��#s�%��jr�T`��\]�wlGbQ�Yc���T�z-�wlJ\kx�3]k��B���oh�)��0��`�r�)rC�Q:�c��N�p�t�s��F:��7��qU��	ȗ�1)�Nw6�ۨ�õQ-�4�[Q*�1E��(��'*s��)v��f@ۂ�e�%s�E��G%�ް�t�m��dcJ�����$�0�\@�HΪ�"�gr7�2��b�';c"�;O�0��i�*�7jpݹ�]y�wΧ!W����H�������J�Y������C���/rnP��vs��Ά�tYh�HQ�h�p��pL]յu��}ݖn�t실�P����Ώ����+�4N��:�Z�Q�|�.����rs��<T�;q�[�7���d�;T4��5+X��q�dIfgG0���NaQ�p<��R�`-b%���EJ2T,Ӡ���r��5CyA�`��Eh�3��(�+17�����(^02��mvu�4��fN��q(�ۋ�+bk�gG.�I�ܬ�*��dVfJIR��ciYOxvl}�[��3Mr.�����Z�#8���r��M��=A�yG�)j>��dͭZ:$:�:Ŏ�����U(;��,��Ÿ��钱�T�Lq4�ڮ�O7� '��ٙי���8h���`��O~�Ms��VS�딃j2�|(݌7͔�f���ft���Y���d�M��w�"�g%Lx��tn�>r�z�!t��:6q��wD�̚�A$(�C]Œ��쑃�wov�씮�}ɼZ��,��}32X�f��K�1݃���hvstNT�.g�"��rV��U��v4�C{��\��(\k��1�_:;{Hp�s���«[wR�}���-F����`Wr@���QL�)q���p���B�8 W�p�]�w��հ��ݪ1�=�t�6(d.�sYkE�1��5��͙�Ҡ��Krj7��T����H�*��ų�LԺ�2��q:�u����]�����5݀�]��8�۹&����4�p���SG��$sr9*����o���G+y'��r��k��֬|3;������z���1���3��<#���5�͉���V:[ٍ�q���/���o�NB]�lN���a�u��vK�])┴��|	x�����|O�r:�P�א�ݞ�8��\�jJK<WbxƀN��.X��م��ۥ�*��V�-Sx�J��@P�H�.H]^^ꥢR�=nr���ec��3�X��YN��2��N�7�|p�C�x[�3��5�zhq�:�yœK�3rrY�쐥u/H*����uC���a��V�|Mw]]jG��� �LJgkB��{�5�۠7V�6�[��=Or�[y�;a3�&��������'^�S��2:�c[L�WcN.<6E1�GWQ5o��t���z�cÜ��F:��������L*�&^=d���3r���_ t`Qǘ�΍P��j�-@G�L !��  V�!1!.!�UD�R���B*/2#�#�Ur����iʓs
��dUZ�J�(���Q!�
��eQTZ��I$Er3D�!g.QȈ)�"����2�]PHK�Q�u�(�� �s��¨��Ԣ�����&:�"�Q�u)�TQt�EV�G�-�EU�:+�r��4I(�#��r��D�5e¢)]��=#Պ�J*%�j,�����Q8u$C�`:��˜H�SZV�q\��r�T��
.N���S�3s/J��A��P�2�!�@�5u�ΑD���NqZ'C����W+n��%!ʧZU�*u9E�!,�QdE�s��ey�\���Na�B%@�XR�sed糗�rIv���-=�zj ��*��Ȫ�$%�w, �KJu�Yr(C0�*�=<�����N�^o"�^�\&XD�t@Vǭ��|R���#�e���|��&*����6�[����뻳�9���R��dW�zr�6��ߐ�M�x��������Q�SO�/�̆8\d��1���S�^&�b�I�U��h��]���a��N�~���+��͖<�W�y���r�hP���+��2�)���[	
��O�)R�/�PB�CW�;�PT���Ci�C~�>�k�{/���|���K�z�����<������Tu��<bҼl��?r����f��4��{"Sv�U���U{�9�V��޺��r������s�z�����(��	H��ߪ�����=�B���)\�ˬ��Z��XD�/�*۸d���<��/Bu·��U��]~�θV^L��W�f�3���W���ko/[�p��1`z"��q��w����*�?�w����Ke����p�x����xr����Z��}	�d�����g��3��>�2�c��O�"�z�7�,��>�x�L%��n<4Ί9yU�`�V	��W^���߲X�;���Um_	������x��Xe��c�i����pT��t�7�u�\�(\)\LL7r��+�a��ɀǶ�j��9���y�$n�2�M)[�&e��&X/�5���e*�_w`����$�����x'�x���!C�g�!�Z�'����-L�є�v{w:���>6�4E���ށv��+-r���uMȶ.ħb��G�fն&>}���;:6x����)VzC���&ӻL���E�ǶH��d����F/T�c*��\�Z�]ެ��q��z�_���ឥW㞝�
�����ܐ?	@��/�64��eŧ��]*^[�5�a��R3c3}��}�įTC{4����y3:!S�6Gu��]z�=Vg�%jX<�_��g���v}NQr{C��=5�*�?Y�o΀�3f����� ��4�5޽�
��n��c�a^mhy��=�Lq���,z߷2=}wêG+v`��kV��e:s�	=Ǘp��EX���B���QR�����uW���<'ԹH�z\ U]�d]�r�w�z�� g�U0{�0�o��M�����=����ۉڇ�>���|�e����"���N,��|s�����w����=q�h�^�G{m	�N`��K��3�0.�ה<�R��8���:����Q��|��c�F����q�{W����_3˅ $@�������R:���:0��1{U��S.�U3��q��Q��s�����c�\Š�5���}U�X�,��3k�Ж���R�v����J>Y%��U#��w�lG��څ8������V�j����t���z���V��Զ6L0K����֛�!���	��kُk���8ru.�yi�����		����T����{{�<1��V�4�����#��#��_�=U0&�����L�gT��^���</�:��8]�̫Y<�xp��7Ǒ�J�.#��Yz@(���z⩉�<�&�Pl�#���g؃���ʜz���o�����!�T��i_K�\{�,�d8="~���ͯ���@�s%�p��bW�����]X/3r���u��[}=�Ad?Q��G��f=��-�3!��� �¢�NIe��$���O�C��XûN�+t���:�$_�P-�{���u#a�4���#��������߼���i��K�`v��=��o6��^�_y���^����;��kqr���|��3ۡ|`?9����Z��3q
��&{2Ǣq`��A�\�z�I���dV�FϽٷ$�� �&X��Q�Wϫó���g֊���_x V=�*}�5jxQ�۟5�}�>�M"�XnK�뉺��#6�;�����;�9�JG(�~�Y�2��^uo����>�A_�~�<o��Ȁ��"��%`��;ƽ�A	�����}��^�:F\��b��]o�D8��f�f��{דi�ɬh�LvPtg�l��m�;%4~*iI���]�z��Wf���L�!�q`lD�+�y���O7Fw&��6#�Ny�� ׹x�Y���_i�kky��gvR�&us������z���ާhΦ �����yI��u�es��vxW�2�$1��xS_��36��9wOc+�~]6���������r������0�9�!n��.��\{�O�~�oaf�S>}欍
����E벦6��:������y׽��X�`���p}5��>�;�Xzi��F�TԬ�B���~_L�(�����uI���X��,;�1������E�iW}�1Nh��e`�溣.�pY)�8]Sn{ŋ��H�Y�ޓ^�ɡ��.��$��h~�N�<���M��\S����Up�y�څ�x�S��}�
�]=W~ঞz��>�-nf9�q����c�^������TD���:�c��_���	�f�lR�s�o��p�����W���p��~�`~��D?!^oW���<��c����3V�d8�1�.=�ï�O��K3���Hͦ��z�Q�i\M��֑~%d�sۍ�rvҧח�|�����H�����Qj�T>G0��/���n�R^�z��v�R���#��oNe6�ַK)h��X@��In5._���Rg#����)�,�..��$�z����Sޥl]��S�_]���q��;�襴U=��R۫�U��K�(��_��{�aS�WV���{�^v'�h��!{�TG>��4���zI�:�A�V ���'C�R�<O�W�v����D�S��ѐW������bO��k�.��8P='qK������\5��b����d_���Y��8�4	#�h��X��eLc����[�g��,ǹ�d>{=��e����/���0�<;*}�_1r|=;�9�0O`mc�dE\�G:)L���g8�HGU��	���S�z�۱O��dp�za��u^~��#�^���]�ܛ��*���~�_-�/�T^��è�/,=��Q�7u/ٮdp�c��_]uʾv�33ة�	�w�k���(.8'��W���7�s8��؏{�{���Q�;ѐ.�N�J�9YX�/4��a ��̘U�o�c";�_=먳(mY~�*��ٱ�z�O�~�Գh]�5�^���Ź��|�`�kjv*"��RGX{�LeFMi`PC��#��m�EO���>�q��u�H��[�2��hV�����b�Д�ė��Ő밦+6�m�N'��T}d���Tƻ��ˎ�]��7/�/������/6�w�y>���ak�Ύ�-�����RCv��w�k�nؾ�C�)�^źOBO���b�0-�V�Z��;�x�|Y���*c�Dz,s1>��g���uoV�ޏ�Q=�j97N�-���e�(�I��[Y4����F��������̽��i�i\�������Հژk6�����/�˿����ϓ�<���[ӑ��}�{�a �@o��x���홛�
�8{�@�FtsqN@�n��]�:�Q�O�����:�p��Mgf����+k�����V�O���rK*��Ar+����M�<�=t#��6���K׺������n��!F���	�X2�QRX�#눘�n�H�W��JE��k̩|�]wo�ϕ��'L{<�^��P�~�E�{��w�g� �Y������^���J���M�3���c��i��=���t��ԑc=J��!z��/G�@~t@��5�6�i��dV��;ȯ7ϰh����xT�C�̍0�n�o��yU��G��L� ޅ������]ۮ���z9��je�W�y�B���"V���oix;�>1s΅f���4�r����u��3����2a�u7PO{����mZ��`�S��͖=����/��h^�y�/k/c2W�Nz;�oU(dw��~۸��p�����"$������y���:+H��~�>�X,?\Ǯ�uf[�Ζ:�7�_^�3@��a׏C�ߜ� 7�f�S���wY$����k*CZ*!�Ҁ�f�kt�#G��3�"���U��.�_Lzn��S�}{8,
�RH��n�G��uSx�V��*�Ș���k�W���1��{������(�}t6+�Gr}���l
y�����t��Hg��V&��=��V?B��Ђ1Ԗnq��j����y��p�_�y��W��<����|���៙��?z;�g��bG�X����J���l��&2��S|rF)s�.Η"3as�G')��7屏�}���r�dLÉ�9��l��Kal��^p��
%�ΩT���J����~�Hw���+;\�;��c�'�s�#�Dx��쵩ْ�=�36�{�.��͑%TL� z⩁7޶�|5Կ��c�-��z�К)v]yn޵���G�W[�n!��欲��%���qT���^���Zɮ}s�$My�eo3|���uzϓ��~wE���9�̼z�C��3���]; r������L!�j�Hw��9����Y�}�-�nF��U�|$/y�>���G���~�dxd�W�!)m{&`>sL��x��zu��xM�v˱`v����*X�#%��9�J߶��__�\�ו@�cc���uv��tj��y���;�d3h��/��r	h���T?~n�m�V�l���zY�n�m�� �z���\�u?xp��p��kVV㬬�p�>J�.�p���M81
dV��V�ٜ_6���澝M��:���Š��r�1|�c璵�=�XF��|�S:y$��ܙ�fҨ����"���`��:���iCO��]��N�[���}���yr2��7�T|?:��W<�F/�9�����V�3Q�����L>Y�iJ����p4���>��;�y��@�|Q�c��CQr�Ȩ�λ��}ѵ�C��{`���ҝ�q�^���<(�>>y*m��<�J���_�j�0�����pD���{�/!R}�7��7������Y>�_�G>~ڱV�D������s���Sys(�<�����ͯq���e}�lM����Rs����v$_���U���u�r'�f�^���%pULm��y1�je�����������E�~�s���[�j���%˯&��fN�p�P�N�/~�ۅq��f�����~�;���4�o�F�W��e��N����9�T�B@z�i�~N���(uE���\eL�����Zٷ۪e���z��2��.�#I�^G��F��%#r��c�(���i&Mn�\�����}U9燦}�E�^�����N^�={P����>ؙF��.bK��Ǒ:�I�]��N�+�oU����L-�R���{Kp��F�H-�b�Փ�^�cV�J�yUX�����.� $,��"���2uՠ�=w��r��.�[�	���֬����|�υi�\v��g��b ԠnLt�Ӝ�ktdy��4�^���y�<�Qh��j���5�>y��.�KG�z�:��H1hߺ��y�&��>�b���ƫ�t��\��vzi &��D���5�j"��C��9��ǽ�q(yzF=i]Q���Q�7���p6��/�#��<��L�l�����KGۑ��n1*��^���n��Et��������#��k��:�p�\�`�����,:�T*������wg��2w6k"��mVߥ�)���pl��%`/�:�����zJ$��t���}�������Ȟ�d�Q�:=mUO�MF�-p��W�Dc�oھ'e��g�Y7J������#�h��3���;�fq&6U��ʑK6{F���_�|������O���T���Wɉ�U\�k�w�g.�}t�i��Lb��HGT[�"a#�_�����n��f���~|}�Ǫ��Q�U�y��W�nv����댌7߁��ü��q��2�r����{�ᐽTYE�?ɏ�z��-SV��F�5�~��\n��n3fV�G�ϒ��1b��X�ީUx������b N�X83'DI�;7I����M�OMj���5��0��.�_M�:�r�{�ڵ�g]c�{Ma���7���\��F�#�՚���,�t��N�k+��.��u��❙x��p�͝y�Ż[�;53{WK�Uӷ9��訮h�|0EP��n=�lO/y�,��b�\�:Ƀ0�h!Z�Ag|�
���+۟Y~�:�{��z���ղ6��/�3g�m�@�g����o�*���g�Z�;��g˪�ʞ����s#_�z���o�u>Ay�;�}���w^ۅ�������W���o�<�F/0JG��V5�>�S]Y��%z��/�,���*���ݚ����O���w/���+-j/��[,�kW������ը/'T��>N� ����%ZATbw�!וǰw��Ϸ��jP�Ǘr�SU�Ki�vX��n��JW�̩3�*���@��������4
=�ۇ�JO����wS���>�|zwN|�����w�$���Ar+��Ш.Z&�X�;v��MXz��G���3�W��lK����*L�N��[�t%�#똘n�I�w��/N�{~�9��d�����P�d����'��x��ҋ�A����PF�Y��;��!���e�����v^8��l5�KNA)�S9�8��Y��{�N�~����� � ���`�1���0l����cm6m����cm������L6��`�1�����cm��������o��6m��6m�����`�1��M�`�����o��6m��`�1��m�`����6��6��1AY&SY&�����_�RY��=�ݐ?���aT���(
P
H� PP" $ � *�(���E����RBU *�*�
�)	))D()�U--�@  
�9ET���J�T(�������*��)UT��@�@����|  �� �R��V������f�,k�RF��4����( � ��$��f�*��r���)JP��@ )^���Ҁ�5�R��@	* �f�M� wpEQ�Q(�VZ�4���Hl���
��m!V�l�&B�"
 p�Ԩ��V��mը��[4��1$Qb�Hf�%���8 9E$iQfa
�Vj4Yb3m�6�٨h�$,iifb�UK*d�Y�U)
J��� 3\����[)�ER�,���f�Z֡*�Л(�i�L��ecl���B� P�� �+�Jn�*��Z����K�3�kL��T�&ʹ�d�P*��R�Ѷ��-IT! QD� 3�f�R��U[ڊQU�V�dl�U�յ���QB���ZTV��Q '  �(WmS+e6հ0�
��i��m�`�2RF���J �8  G̑���,�Sf�P�%Ykm	ZP�E	@l0Ǡ    50�IH�d4F@�dɐOhaJR����@�M4`�L� EOb4�      S�A*IHd� hi���%"2��&D���=G���y56ԂM"ST�      ���I�,�&յ����`lk��oS�@��(�9(��pPT*��T�@@���}��g����~���A����
@��AD�5H	�L ((�x\���'�ӿ��~J*"4��Jڍ6F8=���v���Z4(BN\����?�x^Q���J�JJ��v�e�������t�7A����Eڥ����OH̫��=j��,��-��)�xWR�z*�+�DD �y�$������٫H�:Vxm����"u�'��Z�Z�9�R�[ͥ.!��z�nP��+]��X~�6)i"�ѐ	P�-Kٖr$K��1��4���ɖ�h8V\̤�ͪke��5dx�lY�ELn+���dLKv��H!�M[0�,Õ����x�i���ZsAze񽧘IF�iY+-V��[7�5
���!�v*C0ǭ,U�e���a�4��`�6�4��O���#m�V�E�-V7��w�	A]�ٵ��ʙh�+F�ǹucL�k�K��ne�U�R��Bo4$ԛ%�4M�v�Zm!Wm��������U�%m@4૔ b�]��ٔ
�DX��N�Y2�����vV�+v���b��7u����"�n
bYˎ]�l�Ĭ]�F��ԛݩ3m���͏f���epZj֞j��tBYu�oV���$P��f*�>˗��"9GX��h�EP:+N}��/N`�\WJ�An�B�������E���ګ˳�^�*�A4��Lc8ie��YC5�dܰ��n�:/J�������eZj�`�<��_`A^S���`�Z��	�/(C�0
ʺWgv^	��\�t!�,�蜘Z{�X��
m��n����K��ⷮ�!*����+nON�ɠ-h����v��ݴ���̻���;��| �0 n�ɏM�{D���B�I�k�>�åL��|,U¥]3�NF��/!�)V�DHU)�uڌ�m���	�2e���WI.\_qu����{�k�Uk�8��+"����e�2�{o\�eᲩ,�mF�t!'0��b��ݳ�1��qܮ���kn�r�'�^��@.�7��,7�)�����_&����Ūl�U�x4��gv������;�٣�S�p�	�ݐ�J�0�EȂ�K.��6���F8��ǲ<��Q|:�s�yd"�������J����=�@mժ!�
�~�aԍ�E�dҍm
V�HR]�*�#e����	���'�B�j�K#t�[V��v����_�i鴐T$1Ft@��ؕ��uJ9�h.}C2ͪ�5ԁ�k�Ш�L��E�ѶF!�1V��Cw(�*�+�ld�mk�*
&���o�R����U��o-Z�qZ�5=�44f�W�����=+sr�V#n��1/u1${Z$�q
�����n��\T<+���k��ޞg�C>V��05��T��g�ԩM���׊�.�QJ���wN��ُl��[�ȴ]���-\p�so6J��#�|h�L��w95u�U����Fmn�V�����+Uc*̭�Ss2�Em�A�BER�N��@*feCgÕtZ�Ú��kŤ�#*�Ջ�z鉻���qc��q�Xl[�5���'��[@�);ŷ�y���1�����'���\ʡǬ��o)'�՚vE�v%nn����`��a�k'�`0����e�2�݊d������E;Qh!l��Bڢ�՝:�C1�q=��eZ��RGZ�!̭��JÕ���TF�{r*	譏0�I�r�'�亴�;�t3FT����$�Ӵѽ�h}o�����zN���8=�f���ejuڑk.�SҩqL
OW��-�jDaT���A�{���nnϐj���X��M��i�ޙR��-�E�w�����0È$��7CDmeJ��="���{"ؼr��S�*�Cj��LDiF��W,V�d��QGuy[��U�[3[N�]a�<��j���:sB�׳@��nh���U���U�s�v}zNP��B��ҷ���e�-�{VR(14R���A�c�uN�b��������U2&f��$�uiPm��øԬ(��FR#)�+3�W�Ń4
s5��kK"u�")<�cv�a�fnU�ws*V1�L����nj�6��y�hAD�6�m�m��M���Om��)]m�j\ذ"Ұ��/6ԅk�&����|K���d�M!A�f��Y&�ق�')];�N�YeP8n	k36��++&0QIϬ�`F��va��՝���F��w;���+��:�i�*�Yl��o̰�1�Vl:�!���p�� f��CTא�D��.��t�i
8J�B<1�Ȑ�6 ^e�U�,d7��bXpiٺdG>���Se����,<{I�a�7I�甹n���ZzV��\��v͕��s^<�c�]�j�3�V��O1��Y9�J��eJ�4eG4�LR{r=X#,��֡s��MbL)i֚%��VQ܌|�� ��V��t++�S�X�>�yXLʔ��)ܗ*�iҳ9h6,m��{Kh���j�"��Ʒ0XT�!�l,-J�݊���8 [CM9gv�yZr,{Cl��LZȵ��� ��d����~�ō_MV�B3���H�4l��J���=ʇr�0VKB�wW.Z�Z�k���f��=���B�Ӂ��r��i]�N�[���N�4���4t%��2��h�������3J�>{�������N��y��1�G/�jţ}����"�n��v$1_�U�tl��eї}����]㫦�A���hE�^�b<�K�^\�q�ث6�X�cEd��4�Wowv�bV���*���^8-�� �#�m���f��Ʃ�J�;"S�!\�ޱM�/
Oc�&���!Q�wqD�0�S/6Y7����򝼖.R�ڲIf�	�N[�8���qXj�h�� �HM��[[t�v�w�$,ih*��-[gXVöow(��e�d���/%��l�:²�B�Vֆr��6x�l%J����.��x����B��Mzi���ֺږ�e�ѥF����2�*���y����\��gy�끸���[Z�0��n�Ғ\�q`(�k0@���Q+Q�����+ͷ�wq֢jK��*ܼ����k]\
驋�����j���NE�Y4�tr�V�-p07�z@��D�Vi�r�������4�H��Y���̂�١�Y"�D��-�;�
fY�QX+t^<[z��&So��xti�hX��-���*޺���n�1OdZ�j��������MQ�T�9���{)�T�df�fTՙ�[y�֍��F)Z��^���wSӆ��G�iY�R��fL	+�NYs0���sK�q�̬�H�@[A�R��>�ZE��Ѳ��]��'{�H�E��9��@��2i��ydh\�-����qn4g#3��捖L��ǘ�n��֦��qJg	��[�R�f�1���[��Z1S@q&�YA]mj�9h�m`�HJ�x����g���Cj�M�2�iY���x1�ſC���c�t�Xkt���1M�ڼ����0��/me[;[E�b/v��m�0U��6�*Uux�^��S]�j�)��^�� �JO�W�F�)�n`��,_Ζ�y�n��mؙ�n�it�)����V�dE��7��o��k7,�UX�HucM���a��^�H�5��s@n���G6�"gln<�ہ�*âuԩ��H��f��z�T�omZ��f\c>ą���l�b�������L0Rt+����,v�n�V[4D�0�H뽫;�qZ̦ku�p�te=����3��%��0�����B)����t6�+���haܽ��uK�v[��^4E��F[��r1���n�AS��˻������$[�.�EP���	��v�4�f^[�x�]+-����%�]kۂ��ڬr�%c��GN��hi/w�>,�yЌ
���>6ƫ�9�mc׹͑uoc�
�//CJ���uB֬�j�J8��soXO",�BQ�r����X�f�-����*Bբ�Z���J�+��f}����\*�I�^��O�U�mwge���������?�C�h��P�%�4�CB�)�wK�-ĥq�X���ҟUݍu	<���^�eKr��� �6��z:lEm����8՛�v�E���q)PHˬyx)a㳱9[-=�Ֆj)�*۽t�e˦)�fPy����R�f�؂ɱ�wW$L�9��L�=������.,cԔk7���ԗ��yIO�r�ܙ-�i�6��I�Y]g�k|j/s�M�UEZ�v_����"D�	���rF��-BW8;7�
�d�����kU���y:9
��d����϶}�^�)��er�&��urG�����[���+�s��W\�:M;�' �-^,�Ӥ�5�qaPW]��P�W�L/��Y�-=|+�S/�hRf�ɳa��mBn�����L���Ћ@��qE��E�"��k��*��#�w�-��w�ݨP���(u�r�t��ɮ�n3��9�y�/q�&���m��0�����[c�ϕ�cά��y�].�g'��\��I.�y�u�RZ	o9dƏf֩w�!������"��v!S�'�+�0��]=�p��m4�j7��^�w{:�nù��i�U���j�K-O�o$5�S���z#�`���6��l�m�9�q���'\\�U�w��ّݡ�=s�ǔ�]�j��t�%a�u���׆�=��-BN���f���3��PnL�d8sNħIսf,�8)pi�׹�o"�>&���r)֣���u��p˧�Ңz��4ѽĎnWrY��c6��1m���fn��N�:�p����..�@� 6:lo5��]2�^ȍt�1uv��onu�o�m��[������������P��q�ۤ�"$^.w�8�w�X����Ƶ�r���qlJ㹥@��i�F��H;�ġ��g]�HH�.`�ͷ#{D�����-!�K!JH6�^v
���bx�j���|�P0Y���iK*�v�R��J=&GƟ�
�z�[�*�z���5="�#4�i�w�-�mrz;l�����֫P9O a���вш��W�N�<�����G��{��^�8�����ˣj��l�[ �7���7�1�>�*WE��N�ܼ��@(B���곱خF�w&�t:�7�3����YJ��-%J�N�7+�$��W.!����X����i(�d�k�>	\�^Ԃ�[��sK8�#2�R�RQ��z����zۼ���nZ�Ά�¥;�t�g�J�⸻|gf�38J1ڶ�92\鷯k.Z�@t�������#n�[���Rт�Z �5"�ihs����3ʹ�3,<v�c�1rN���P�;N>��Л\�woj�!3\���ٽOxlAh	q���D�9��
��>͢k1��vٮ�wfMK>�u땖�2���٢I�+a˫J:(�����E���{C���Z'� �A+:
�l���Π2d�캁F�ˡ�b��Lo+hAW�d��LJ�+4ea���y5�q�s�u)v�"�Ba��ܩ��4���1I�-�[o1���9Պ4��;M�N�� ���ت����QGT�ٛ9��'mkҮ�:JF��Lc�q�O��Z��ֲ��h�]�a׀�Sz���\'h�ͼ�s# 36Ø5�%K]թ6�2~���^Qô�/-^�!�3�D���譬�v���1��S2��t�o߶+��z�rm)���;���W����N�1�S{ٝ���^��dw5�u���w�`��bI��!a}�$�6gf�/�T8��}Ytܡ�i\׳�jA���
���?�7�V���v%����}w�3�Tˋh��؆�h {�ң_v��]�k�e�l9��m�V���T:噽�P��&�������#{�Y��Xo���cӨa�Y6�S��(#(�Ll�\��o�k+���p	3����P|^t!��i�#Rb��BwQ,;$H��׆�X��?'�1T�4
bZk�L��7�]6������/��B���jF��S巐gk��nҵ{����*e�S�nv";{�R �
n�Ў^�M�D(�.���$D�5{��E����Q��ϟ>�t�}��h�IN���7%0E�qg�n��{�3���x�	ɲ�mus��M��Ikn����N,	�k�EQM��xtm�E��\G=Y+aVpM���L�gn�l�cA� �6�_N�u����q���I8U��X�k�fi�������öɰ��G.ےK�\?���'aD�:=���һȿ`|#Jx���WJ4[��am��Y �aysN�\�e�k0|�اX�˺JK'b�4)//��fK�Mݲ��]���6q��3��d� �.�6��ѻ�.�J�ut�CUaq��xD�]v��tz�5��'p�m�u��+�9#�{1����J�r!��j��"�[��������g-/��k�c;�{3.���Ү�Wh�+�*����J��nc7��GY|�tV'�:o�Y��*N���"���ȓ��F�ܗ����>�=���ς���q��-�j�+�Wc@����7�C�ɬ�n�\��'S�20%n�'��a]�*г���#��E�lBA�ʔp3��O]1�#����6&\��!Y����;{1��G��e��s�K�rkqgoU���c�n���>�h;����*t���X��Wu[T�s4%Xs���v�1�\�؂ʰ�����	ݝ֫9]ln�A>ˬ��4�(��ŝڐ�u%P�^a��(:��]�nI�h����f���V��ٮ�A��-P�Og\�� �*���ƀ�[�f�bøB�N�]7������ ��Z����=�oң칤�:9A�n��(��X�����yP3l�[�f�v@���ڍa���'g>rc=�N��i`Id�v�ô>�T��:op��75��B��,����%-�^�RlW6JTxq���i���Ա�n��J�Tp�Rq�,�P@6]��m�y�W��T�o�>v�fB�����ruf�T��`�(lZ[��T��+`�/f'���[+X��YN�ꛮ'f\./:�L>c��4�Ѥe���fq���!Y��{P�a9��\R��*���1�œ�J�̧�隭e?=�sQ�������R���N%����,㢑Cs:�q�gr���Xy�s8To��L����vC�6U�u^Q9Q���i �mgW�ʸ�G�X��۵.+3�u��N���=��	�̫��K�+����yp@�
�^9�l��q�R���ްU����c�u�D�y����H��G����ur$Z���D�SӚwF�얊�vs��p�Jv�]�\L7�����ԞN}5�c"2�r��	+w�x��f�H��$톲�ЕjM���7h�u`�[h���M��q,fG�W+;��m��m���E�Zղ���wv�'�:���qob�w(T��c���nt�խ� Ȧ-�;J��e�_N�f]�k�����ynt�����,�}�:77he�csr�o<K��ۛ&��yLL�vS�n=�$�̺�SnD$�Ӵ���cj�g��7N��7yI$�I$�I$�I$)G*b2T���Im��űl�Q���Y�q���|K|b��m��F�y���r�7��I��9�أv���9����Q�v\����.��5��]��)�*J"��yْA/L$�$�IRI$&I%��1��۷۫�i�Š�]�|ox�̛{/,��xf���2��R��%Yt�veN������8���+����� 1,R�(N�r��n����ej���D�wɹ��3UC.KM+�=��׉U�7�˛�'�-W�B����ݠ�2�&C��|`0`�6����`�>��8T�[���l-�D�e!GS5���17凕���m�W�q+6�P�R�Сe,��1��9�X���R]�ɖ4�m˹\�s�۸�c,�ٶ�0Я� &���+��(
��T@�L�fUQ:Q�:�$ ��Ȑ��R�F��=�'8@�jk������FR6��+�/2��jXp]�L�:�-��F٠������װ�{g��YfI��0ٺ�+Z[�%�D*�('��h����B��֝�1��X��4f��<h<{r���e�F�8Y���gl�J�·p��&�K���{���z�>{X����s��J�b���U�G.SwC.p�E�;kl+�s]TF�]G��ث�rxWh��,Lk{xL�[t����xK�2>["�sW��B���l���e໹���r	kI���t�7�p����4�+h���Ō�.�<Y�(C������{��h����8���T��uw�nM�]X-���"�	쿌���|����*�Z�v���R�B�S��e��C����V��>*���m���r
Z�"K�(��t�Fܷ�>Ɉ�S�I�-�fN;@���Ĕ�C+x8�r[j��c�R�9h1�v�|��#�Z���N��#e�V3-��P981]�<W��&�6�7�����s�[I��^�u�����z���򲬠2�Т�a���)��s�+�p��wZ�v���F���|��d+N'Ԅ��	�5_1�u��R�rLdWP�t����.�� [}]�������ڻx謡g䍊�+7&���*�����������k
��),��%�������y>��9�xZ7�j�zo�3:��u�K�%�����Q.��r�֦:��v}���:��R�Wug]�ί��ͩ�`��#�%��s{��4�t�U�x��GEu�v�Ŗ'V�}\'���ӆ�؅��ՠ
v���ʎmX�z�z�kHB�ye�q��,����6����f�,ђ�&R��4�����U�=ˡ�`���qU29ԷB�	��0 54�h���vq��+*ާ���v�ca�<@<�
:�0���%�rZ?,�I�p��!�����J�AeN���,��u�U�B��F�ˡ�9�;vʃk]�`Wfh�K��V6�m%����g<�9�|�p�]�̫"�<3
YV"B�m�@��	ʋk0N�3���\YF�]� ,3��!(杲��;f��%�!�a
e��M�)��ãj>���˾����Q��>��VX�/-�bk��l�/�ͻ�#�5Q1*�Ɗ�Oc�A�Fę��;z���۸��Rv0Y�:��woW�qJ�t���YV��;O2��lU�K�r��i�Ql��3,�D�p������e �z��"��b�/\}��E��;�����I�I�(�&�#s,���7��u��m�\��Xw��x�2L�
,6:��$��K�����.�����=I=Ѵ6�	Z�^!"�xm��b�.��7c��kR��^�0��)1]z�%	E���l�iI֋W�J�Ϟ����p��\�{�GWC��⭬�ah�x
�h5ո��n�SD��ݶ�'s����iX�2wD^Cw��y1���9KBwS$���i�8[���J�9i�ܨ!������38�gb� �� ����-d�e�]h����\ԃ�y@O�����S�ΫS+j�IB5]#� ֖vJ SY-U�����PȰ��(ixL8;;� �`��,?�Ha�K wu"�)u�4Gt}:��� �/���y��sP�q��L�i'iV����)r��6b�x̱�Kv�&%�e�a���M�O���80w�k$�ۇ��4��Z)f�'(P
��lE��3F[��lS��ۦ��K*��O{ϰт����m�X;�2�2�@R����RT�;+�]9��TEU�6+9�6*���TO���g�i;���`��Ά3���r�lV)��&��5I�6Geh����£�䭷�{s��	 ��z4�sMYa΃��q^o��Q,����uK��.��)np}��vpY���wg8!}v�?k�6���{M��5Id�c���w��]��"��f���g+
�ֵ3ǹ��L�ճ����ܮڙ�79�V��W�����0V��O� &e0��XK�}���m�������}�G���l�*��t��"�VmcE�l��r�.���y�ȮQ��)Y8����/4����꧝�kPhA"�����mu�H3�k2�X�WS�K޾�NL����v��˙���T�r;`���4��D�E���3��n�=H�����q� ��ir�T�3�)�	��+���m����h.l���v�w� ��j[�>�)U�ӆ�[�I���1�kY[�]�]
-7�y���L�4es�豉�p3::��-Q�t�^�$p���e�ׇ��C���d��4��cU�q>���ro$mܥrN�fa$A�c ��J�Y=�4��0eXm:6z�rvI}�p�\��hE�eup��Uɘ��E}�L�N�˲��9CWH�Ϊ��l��ٶ�գ��#�g˷oؠ�{���Qq���疩�|�5R:��q\�2Ao�p��������f�i�U�z��D�,�)��Z��+κ9u�(�N0�7`Vq1un-�37m�O:��Z�B.��%-�*�.�d�C��L�C�ިiN�lR�ξ�S�oc��;C�nR9g�kxsܪ@��gu��Bt�/vɉ:�W\�3����>@�9�<��[�=yd[�.<mp���;��a+j���P��1�{�et�I�N�H�밣+��Jy�ۙ��<�ݮ���z��
\`���[�>x7�.��lAǜ�LY����m������ [}���Zil�ϴ�Nu�F4��Ʃ�ΐ^�� T��S�-}����Z��S�^�[�t�`.�ň���z	A���莇Pƃ���pM�����ydl�c.�G��j��nͽg�%�-s-˘p.�ıI�M.�sop�3�٭s+\*�X�u��j���k&t[I>|T�YWK�\ ,�(��°ԧSu�3bB+�҅��K)�4�
fIْ���v/��'a�@-�tN}�jHfa���_e�^>�u�a�'7,t9\IO�A����Q�xRY��We�wV�[u��c�80���=�nw=�[�m���&��(�5�e�-�n��E���ki��&�#\+ݫm�W�Cn�6���V��I���	��U�E�=}e�F�ޖR���O:���;�.񾱦�@�'\��v��ٳC�2RA�W�얥��4㕪�t�N4���c�[��+�J],u��Qδ��׼�s��Z��h�����]�e�㊯5(�Oy9��X��Ui�{���B �*�ٽ�0=Q�ӷ-�\���K:�p����J�3�5�/R�T+y�B�K��'%�C��v����1�O~�ǩ���W;���9�?-g
��(Z�w0�t����E�d���qP�4ҋ(��L8�Y��ҭ̻��viA�]L�.ս��F�����]
5Pؼm���v������Ѯ�)^Jt�����Ƙu�&�豽�,��F ��]�\�zZ�l��
7r)�+�V�q���Ҕa�)�����5�r�]Ғ��woh�h*'no'{�r����c�Д����@bW��f��#���i�}�`I��Y,�w(D��z��j����ui+H����i$�R�c*eҽܗ5�:��dH��T��*_GZM�VwPs�ua
��uӕ�CxQ�'t%�6�`�C�`��9�p�'1�3��iq˩���̖k����R!,�.�Wb�[��hb����L"A����w;k)����JݔUFh���]��͊�8�Ka ���C�z�\��7}��!�V(C�M�p�~��|��i�,N��%d���S`�w]�ٵ�/4d���5Q���(Jl�V���L��Gn�5���a^N�;�ݢ��^��ʏ��@%5o�Ca����+W�1��kP���"�T�V;e�15h;DTD�$�!��ij���U�����w��'���M$�n�G��li��]I��E�I]�9�vJ �;�D��&�Բ�"�E�|l��<��y�'@�2J�H׉���[�,C����`��?�̮sMLT��]�Ǯ7Jnu�,��Q�ymX�2Q���ĂW�CWb�\�F�e�b��#+[��(���CR��}ӈ@��r��H�w4}3�[e�m-�mln��ƻ�Fr�J�
Tl=1'��ۖ��h������#���{�F�7Se�U�D����-�Tu^�]X��f�[�ܣ.��h��o,�>|�U%ѻ�s�`|�l�Y��F�Ҭ��:��xĬ�U��UJ�3&�d�޷ٜɜ���.��m��/��J^���X�za@1�w���Gx�Js�q��N�[���r_w�7V뎺�2Fl���Y|�lڕ((D͕%���arD�G;�[�zT�:�K�ہ��	�rS"��ﮠ�]�ں���V;n�Z��Q�;L\��T�Uv�T�h�eżpC7
����mT�Une�1F�S��n�b�q�mUE֕�mu�u��r�.DX���[Ʋĕ8�jJ���X

�
+�a����2㌨c�m��Q��bu��k��Ԩ*Z��T����f\eSŒ�7I���~ʬ?<y��4���7
�ULLfT��q�#��ķ)����ԱF)lZ��h�p5�USsqMv�R����̉����M�nk��j�e��bfPr�E�k6��8�R���7�WM��\廦�ㅵ*�2��ˆf�4�b۴�M)kQT�U۹WZe���;������i�Wd��=�u�jj��4ʳ0ũ�i]���2G��svD������ϊ*�����gn�9]�L���F���u��o��ͽW�+��
��^Ἃ��[9�V���~AI���[T>�ꄻ#m*��l��&|a������昌�{���7�8)���Q��	3�~�N�w����Zw�5bI�4���U�ӓ�\w�	J�*�ݢ)�Ftm�}���
t@DO�'k;:Ĳ2p�8�i�,�x�:��oTQ�����F��:�QO���0i�C����XX��.�vt^\�{�NE�ܡ�M�ׂ�IW��F�dK0s�Goml�ɤ��U�.�4�d���M�&^�."n��j�l3s��9�s6w^dn����q\V����5��=�cX'��*�H����]�X�H6����g=(���:�TR.-��kN��*�{V�|����x�7���+�o����Ϛ���{Ap���/8��t��Fg���aC�.�N,݆��/A�YTHb1%s�8�h*�y-�	=�H��ڎln�P��QٓƵ�1*{�ZY��ȱ����֘x,��5���\��s��&)c���V Þ�f�Ǹ��śvk�x�&�#�Ct8�d�3�r��jj���| m'zi�ϛ���Z�	�s+C��Ϯ�x���OE���k����[RM&��yѳ!w��;PXu��U�n��hR�ڀ�:��qø��fN����R5�5B�wNmE��)ئ��=S����u���T�sd3u�d��S[!SYx)��#����Z��qqSŶ���SZj�#�b��Zj%��[�1W���❝Ł*�rMؗ���F��\�t����(�+6*NE���*��yZ����>u�|MǊ}�{]�+���=�KF�<ߏexg�G��ȶY_�E)Zͷ�ܧ��h��� �����p�q����tl�?-����7�N����Z�-DQ>�`���{�t\5�]N*g�����2�Y���+�oHŚ��m ��� �ې���.���9M/�m���%�$}��N{$���N�@�}M���o���Tr啶�h�$�b�W��Z�2�������^����m�@��L�o+o�>I*����W1fKةbE'�r �b�r]y�R�j�Nö��!_���"���Rj%7*��Yw���3Ϯ�1��	�w�S$	�E���f������k��$Ŧ �*�:4ن�u�c ͛<��<��y���Ϲ�#�f�����,΍��ev�mI�*Z�.*�-�<�d��O�����*y$�a�)�<�s�{�ڸ���0`�[�փCֻ;(���^2Y7��-]���hҚ&B�T�p��f��s�rSnqr� ���t4�m-V�<�+y[ʢM�.V�ȷC�s��}�X�>��c)B��Mv��˲��И���Z腨WR�3z���n/Gub��]�8^�^�y�;��f�I\�:<����.3��s�@�^n&r��g,���,�W��ok��Gf�>���޵��t����jؽ8�L�4R<y�r��
��!`FÔ�#m�2�y)��Ȍ��T!4/�*�:z����0�ƐD�h��|c�d�VO+�O�R,I��p��^��s�/n��blp����i�붮q �)�kFhb�c��s��ۛ��mG&d3Z�!Š�N'�S*�����/�	����Ț��3t\o�x��̊{��Eq�@���ӕb�(��9Gw�w�~�����]��3=1�z��>��Nf�L�������0>\ >[�9R6ow/=ju7ѧ��qvwJspg!��S����g�ĚCe��3���,�H�(�����~(��,6�<��{��'>s'�(�aqu�=}��}^J2֩/����d�̜�M��ٖ�:li����]���Sb�/wp�?z�[n{&4���v����b��켌���{��[���\�9�l]�tͣ��B��D_j��3�r2������]�%�f���*��S�ǂ�������Vk����JF�ʎ��+�z���g���,{쒎j�(�{�M��f�Y���ʳ^�w,=�k5/"�3#���v�:�2#-����m�]���vD��kQ'����Vp5Kxvx$�G�)�Ӽ��m���Q��Ư�&�d&Fp;�;r�>��;^Y�L�z7�D�fzc�1Bzj�/��˽�+��зu��n-��v��8�\�ڦ�ks�S�c&��=��ʊ��W��פ+ �3��W���uՅ�n��+�S����I�w�э�m h�D�0SR��1I��2ܑ[[�L�~z-��uv.zu*9;]8�]<��B�ݳHm�ю���f�m#�<����::�Q�ͬ�W�ζk���(���טJm�V�E�)�ʬ��`�o��
�gk��Nf�梚a��{��F��Z�e�F?As6�{��f��l
}�D�,�l���_d�[PI���ۄ��Ҏ�Gau��qLS�Y!��xة��y('���'{��H�"� �Ꜵ'aT�41=�K��'�,p����>�!S7���؁ T���5�!j�nZ��"�R�^c"��n��Q���z7=��S_9���������̓3[�Ş����/��yi�鶺�]���fH�=�_~��%�k	��MZ�g�e��|�O=�,n�uD������6hv)�X�!�׮�+]T�x��\� ��8;%xuyl�;�vvҤ�:J`t�"���I\պ�s2;(�EZ��GZ��xj�ޗ��8�%���;�eg�d<���ޕ�|��bvl�23��ОV�U���:\l��##i)��ۚ�fu���B5Ƙ�yg��E<��y|��]����n��y`�cE�b�[I�9Ķ��;,�1/3��ٰ�}hˡ��ڷn:����5���zuu���q-���)��@/�a�oy坒���z`�R���Oˠ#c&�䋍e�ۑۛ#��m^�7=��]�S}�noM��4��o�df�ʪg��r�P� �ָ��3�v/��r��Ònc^u��DEٞjp1�4�4"M��r������9�'��13���>�L3\w:&�����ɲx�'�6���x0=จ�R��TCJ��_��&x!GdyD,��y���4�ѕ�\m���ۚ�sfV��!f�	���s��Qsܱ�FE�tT��=�s���������f�\�}�1:�SJ�H]�w~׿#��4@T���������c���"�E��W`v$;�(Z�r����d�����_j��ѳ.�w'�LtE���h<̎��y�˗���J�ڤ�:%a��_p�&�yP�����CG+�7+��.�xz��/��ު�[���urI�4�l��"�]��J��#�����`�6�P�Z��%Eڵ�V�0U��j�'v��Ƣ��Q��,���yW�D����M��r�9�0d,X�	�l�Y��\[35�r]k��ЧvS�j�ңh�w��N�ذ:��<�t�!
� @FsW#�y^��\�Yo-2@uCx��ֲlM7�v0M��_�z�+j�Uw�zJ�U��ӢM+X�Rt\�h�}[WG�Yb�-=����˟F�w^�N���h��[kL���v<Ҍf�sD4��i�v{�2��y���K��ǔ����+��;.C���b+�����B뗁�3���ʺA���8����m�#u���-'��ɍVH�ƥ�W�ʁ�9���C�At)�6�]��r:�6�2�T8�,��Q&@��3h�$�)S�U j�]�Wn�c��[�n8*�t�)W�CvM'LS&�)D�R���5R�ʶ�b�1x��S&��ѴLl|@̎L�W�Vi��TwW����ĪM�wm�[FQ�n�-���d�ҮD��g]�X� G&�P�r�lb���J@�P塻to.2�֞��6��2�w6W�͇/k��ev �ތYU#��t����U!���-�8�S�J�AZqt+'v��AV��$(Yv���N��#�r��H.�t�J�7eC��y
�$MJsynHI�`o(��*�	�@D_�����W�� 31�K���lع��8�[j��J�-�R�V��U-�ܹ��iPֻ�cwl�-h"*�G71�6��7]��6��bn3V)�����&"��୥�\Y��ڮe���:Z"cX�*�)Z�Mʦښ���q��։�RٍLF�J�.n��cV�6�i�]fc\���i��4��UEE�������ʆQ˻[��9j�J����1�V6��5n�is��c]mcj;��*��w0�L(�����S,1Ec��f7]��e�E�u7h�[�fW2�K�eim�v춙�3[R�-m1��+1��h�h�~������J�I��Do���m���vD]C�6����7�)¤
�f�Q����r����H���(���1a+ğ:����mEa��z�l�q�������{��=�����+hɕ?(��f��_tO���`�c�g���_bW����6�y�ؚ�;S),�c����Q6d�܌�H�([�7=�*�4.�Odq��d)�,�˘�J��[��y^Y�d}��	9�wg�,'q�Ľ�Y;���|7�֚�{�(*m3��Γz!+��fT1{c��*�"���N&������nѕI^I൑��ͅ�V%�b��y&�2�'0,>C͚�\�,gEs J�9 5�6�ˍ��6ʾJ���D�AW���lXsNw:��u���K6�[:j��u���M�usV`��]�\��ci-��)=�����a�z7��A0�۷�܃�X�z�M�a�{U�{8�O��Y��(�̌�+	�l,d�s��1��}����3Z��kn�k�'jB��!���Y��;��o�˿`�M�Gk\^�V\ƪ�BH;����h��x#�|���/���|@�������i��>{��"j��׫v̛|�5+���g��к��� r�7�z(-p�^�Ey/"�/|��4_�óbj4�#��-�f��^&9�9:�D�'4�lgt�rz�hm��W��r7��a��D�p��g�Ը_e��#T9-�����mrs����A���`x�]7j],*0�����{�t���&B��v�V�.�܄@u��Ox3r:����u���|�W&uE�QVl!Ӧ�˺�]Uy�nC��G�ܝ5e �x�A\�T�KBٝu
��(W?"���Y�|6�=�J�<����3,Q�*Ҳ U�սk�e����JC}��{�d:���l8(}�'˩r:�H�㼍[ض�euX�-��6���FqP������}g�}���0��!3.�E��EgHo's�pJ�ۻq���qI��K�!}���`Z�'�*�Z.+�nN���S��	�Ǧ�ϳ:�X�q�Y4t�����zM67o�J<�l���S���t�⥆"��`I�r�b=��|S�L�u��&�팃U�F�u��ӏ�E�E7O�]4��ڝ��3mH_*/��꿶������Tr�T�j��$^ezb��4u�(І؞��7\C'��8��7�}|�����O��Ić̓P��E'��'���`z��O-�� ( d�{A�����g�O4���O`}>�� a�a��3P�ROP<z�)=N��ϘxȲ��G��S�"�oMQmLIګ����Tܣ[�+!w�{�خ���H5�����d����(�V���:�C7MLH!��8��Ծ��^��]�DnF�Ҵ���OjN�#����}�|�(l��a�߰��N�VC�O�߰�>a'��
�+;a�O�N�Ӿ���|����ö�;{C�H)�'���x�m�?!�'Hx�l���0��<d�������OYL�v������>��b~d>���zɬ���~Bm�ćhnY!��[ lj� `{�� }����:�����d����C�|3��I������,��~a�&�Nua5!��qI � ǽ�����?f�q����G��ċROY:O��!0��?$����2y{`0��������� ǆ�������Jw����G�q�����d� z�����Ě��2C:��	�'�3�C=����=� /	�W�?S]���\��{`xǀ�����&nd��K哤��=@������N�_�!�!�C���s�O���ם}��O�~a���t���h[��@���'<�t�|��ԓ�ݤ�0;`3�a�!�	���[�߿{�|}��<�̓�8�O?!�$�NЇi�l�E ���'�'(��� *}�c���t���WŢ��ǀ��~��=�!�C�d1��=d=d񐟘
I��R~d�,��<I��?W�����ߕ���W�7���j�w���b��x��͕ۘ������%j'K[-��0Δ�P�f���b�a��b��8�]��sѸ�.R�"e��Yo��1$�Y���(v�z�|{a��$��:6�<dY'L4N�8�,T�#�;�~����sw����O��=d;Ag'P�2y~d���ܰ�n[X04��x�ϩ� ��S x@u�ȷu�_Wˤ����|f x�� �����ԇ�?$+��z��XOY&&����P<dP��fy���Xx'l'̞�c�$XLf�t������X|��'J��$Rz��!����=���|2,��(�|����'ïhC��'iXL|`u=�!�~���T�dԞ0<�?|{�n<����=~�8��a�%C;��O!=a����'�Y=g�m ����2N!̲C�s�L޻k��gZ�z�����s���}C�C��0��/��Sz��iN�z���OS��u�$>q8������C�T'�1���{���!��ROǷ�OP?Rtô���x�Շl'i�!��M��z������{w_��3�&�=�|Ǉ�!�� ��wN�'I9�$5��E�Ѿ�? |��~d;`z�yC��~� x���Q� Kg︾��'��~�R~�1�R$������,��7�W8�D/�����q���n���,�X#jy���1�ct+[��b,9���7����uj�(:��c���s����Qe;��).�d*4	�f����]solP��]y�=㿼;�`q�2��|æI�?&0��x��i+	���$�{�uh{I�N?0?0� �9|��^��o��C��x��&�Bz���$�a�`O�B,�'�'-�I>�������<<c�銬,Fֵ�)`Mq��@��S��MOP�L��v��� Vv�<fFv�/��E�� t n8[�^��R� �hzc`�	��yg���|����Yd>Bx�l��v��,&ޟy���������'��d���M�����OP�!��!�:`nP������c u�$��si�_>�o\�9ߞ���{��ݰ���+��v������h/N�����o���*fY!O�=@�!�t��w��}��~��Rx�z2�|�%a��'��̒/��uB3�'I=@:���	�_YN������>��N�'���䁓�!�"�>�<@�N�O;E&=$��I�G��%g��������Q�=����U�x��ǀc��L	�5'H������x����@�u;a<d�݁���(MC�4��}�:����y�_s=!�'ɨb��|�����������d<d=I��:��PІuI�8��>'�������&���Q�>۪�Z8 ��=�-U��3������������'�;H�֪b�<�w �eu���^Ot��0�}K.���,?�%�)��w^��&0=CY&��9�4�x��'�hI�Ol'<M뼆�a�'��)��x}�"���F�l�w��~@����$Y0����2[�ē��=d���E3�	�&��t��Ǉ������\}�7�����~bɌ���?!����v�@1�=��f��<I7=�<dY'��;�c���噐��r��/d�lx%�^�Q!�l��'IHa݇ԓm!�O=O���!Ӽ�v�ݰ4�����w�^��BT���}Bz�a凉�������;Cĝ2O��Y!z�2 <&�������� -8뫩'�^�"�>d�N��Y&��'�T������VC�'����� �XBal�'�'�<������ϻ�����d��/);I<N�=I������l'I�>H2t���o�P��<A����p����7D�q��|��DT�c��~��}>��������[�&kԟ4��e�}�[i�*<�/�8��0�-���$[^����x[��1}7�؏�E7j����DY�g�e�3n�J�(�J��qc�J�+���v�s4u�W]N�6*50�����2s앑�.\��	;�˗��rtѲ�X�{T�,�ˋ�{�|�������'_t��LUR�us�&}�N	s���q��gTQ�i�LD�4����n��Fq��ĬB�x�x���r��%��v��0f�«#q���0b���x�\��0:F�cf��D�>DӰ�:W5�S�YG���쵼��ECJGc��Yճ�uQӳm�tS�vrq���|�e�`g��'�\R��[�W&�g�J�������ڣ��KJ�}�:�Y���!@����\H�o;q�xՂ�ٙ�$�ۚ��k�u�����#W;a��0�����v7	M/��jn��D[���;BN�t� Yիu�y�+�.`�2dǷf͵��/�次�E�RK,�����L�<{�f�W�Ȫ�:N�B+��reҗ��w���e����B�i5�楔�+��@(���(��kv]	]�/^{�c�ɶ�*�{^o�=�sy�Jb�\�}���2��4!OQ�\��!NY��v���T�A��!`�-�ΊYn�>��i�c��@��c�7�uBw�Zja3�QC9r����G��f��~7��#4����J��-�6�.�.CJھ��n�j�؃�E��Æ;�r�۵p�R`jv�]t�Й��4�f�]�� ����_A��2M��)�xe���뚶f]hƫ��#��7�XC'���ۮM��w<��91v ��v��I���="�\�d�I��G!�����솭�:]��f^QVL���;S�BZ�X��&�8bTV,R;{��7�d�O,�ٙ���V��Futm��R��=p�I �"���~�o*[��u�S���qp!��ύ�}�k�\s����Q��Q'x����E��	Cq����+z廛�h�1ު�f�%���[�V��啭!�i�k�����KFe�;��
Z�[/�듁R��þ="�8.��3�d�z��<Ж�O��U���'�)��BiЇ(��Q�Aٽ��l�l޿��,E���~�І�u�d1^;fbw&1�\�c+�k)0�b�8�,E#��D�]Y}ի)8�Zpv���)X��6����75�rI�C�JɎ����A��'17I�S1����v��l:D'��x�,��ǀ���̅�Y������Z\���uf��e�0�)�p�4l����0�Q��]ѥtr�l(/�ے~��b�eK.��=�f��Ӓ:~��=�.��b�HN��JC*���Z'
wJ ֩�gQ�`�+N��M�b4�tT�MLY�Gw2R��,�r��GNp�ZlY�H^P �ѷKLN�hm�ft��i���$t6�����w���B��R�((�M�����*i�H�ʲ3adn\vV)q�;;*�oFA\�"2W~����5C�*6��k���ݹ5�-�ͱx����!���hL��˹�mh��]��ܢ���p����mܸ�jf4�]±��\kK��̣mL�0UV�Qjˑ�%\F�2�Ȉ�5�Ƽ��Y��!�r%˘YP�*��X�%��P�*��jR�F�k�R��*)A�j�q2a�������QU��E˙Qm��Ԫ*-.%��ǙU�D�`�J���-j"R��6��`���Z�TQ�Y[Km�V��2�P�Z+-e�
UU�	�~�f���*���m�Q'�Q���[+Y[�賲�tT�Ȼ���=� iM<�ώ]Kޛ�~��C���S�o,ک�q�]��'��د8w�J��~;�i]M5�ÑVз|.���^F���ڻ�tTrp���.�+|���*k"�ތm��R�*`gr��V�ߦ{/�;؃�*�����9\�zYc=�T���P%ߖ��;���-mx'�+�_/^=�Y�E��}����Z����x��>��6{�v�y�i�1Qcݘv������˗�3bۙ�2���}o[q
��+�����X�vUý[��8���m��j��%0z�r,�z���S�O�F>c�bՋY���Iʕr��m��\�[�3y�:�x�d����/�{�x��4�C��꒨F�#Eퟦ�'9a�SL=#������;�O�[�,���V�9�s�D���Ǵ�ԡ��,0i��x���Mq(�D�Q��՘��d�0��LK�A�[������-7��@��5�}�����d!��H�==�.�[��>�}���C�)�&r�!\�>DM��W��'�b�XJO-=�UQ�[R\�Ī�5�d�{�F��9��y9��5���%�V����(��ŉ��	�6f_n�*L�f����'Đ��ˌ}��̸��܎�[&ٜI�Xky)FT���U 䴿�yU����i撗�=�'��k��a����;�Q���'a<�5�{Īq�a��u)gi������J���9��&��e�WK�'�D�V"��"`�\U%)�1lt�µ����<En�P�9f5Ѹ/pI�7K��U��������}�َ�o�ｇ�%�Q���v*��}[@*|�Tտ0:i���ւ�n��,��9��o+���gsN���5P���a�(l��O�Ʌ:�!�T��	�:!=zD��������e���V@�=h���<�6č�'pCnd�h�ֿ��=b�z��4��w��7�L�r�7]�ݾ}�.L�kk%�H�5$W����
�-�p>S��
Zծ�}xu�[�����g0_x�?'�/\�ر�+:�j�tF��z�׻�S�Iˬ2�7�=׏Q�A�C��T��ʕ��u'�OA��W=�w��d�F���T�ù��·b�>b��A�d/+�2]�P�j�y�g�˴���z�s$&������d^�n����l��-?G���I�F��F�m�D��
�BqЖ���M�Ll-;:;3f��Ḹʮ�H��Ȏ�.;W63i����#��ykߑ�+Y#��L�i����6QӻR��B�j����Mn�; ī9\Ĭ�d\z���Y�=�f�\ٴV�$W�xx �&\�~��|�8��T5\�Z�G�y���ǻ�^)�l��l�9�5��M���WO\�{W��@��u:Et�tKU,��:.Ld�~}�0�;Bߗ�j�N�Y��J����N�w�B�^ޮT���l��(�sa>��}Bf0=���*�s��J��2�n��z���v�fF��,Ϊ�g�7�L���#!�/1�o�
�2Ԉ�6��mR۪�y��1l�ޢR��[8qTl� ���wr9���=I�'"t/jY�:>�Y�)����r�J����֎/4����PͧG��,[��
�Y�.2uJLn��:͘��+�Dq���W�xx�9��Fj<|Ej���LR��^"a���YD�Z�_v�5a����
��:#��e�1&�9ia��F��mS�*�Y�����O_���5���w"j��JƊ�F`��Hz(M�k_I���L�|�A��Ӂ����[B.F�,z%�=Yx��y4���/�4�q�;0΍;\��f�����^H�̇u�N^6���w��1����x���K����7V,]y�Xf��+�b�oz\"���2Mj,̍t�y��z]������y���ʾ(N{����j�̛��Y�1D�7���Y��J[��ԗ���4��=�U.6��_�'�1W��=D�"��f�G�.{�Ǎ�{��_REc��g�!�y��ě}��{�o�؅/ϒh�:��Ԧg5�;��ը�VM���LWr�|ėw��=��]v�p2��wa��J̌<��e�[ۧ�3ٸLQ�p8ĳj����͇�ƇA���s�᫮�,S
���i�ޯ_���]��nEB�u~�/Rx'����+P4:nܓg;�5{���9�V�'8|D�Mx��b��k�.rz5�{L㞼�v�.��
����\��ǳd#�$1��9�.m�é�r��y�}%Ks9'Y���];���LϬ�Z���N�vtAѕt�6�+7&��,}��s}X���)| �
U�m�-}&}�Af��ۃ�p"�bxm^4�Qi�芮T�uV��}�O�.-��tXK]!wtU>�hvU��n����L^9��L�sbS��ŋ�ä$%�燳��:N�9K���}Su�����kq������sW��*p�.�
�1�{�y34�on��������<b;�B��W�`S ����Ŀ3��Oo���ɘ�o��X>$�/+�e�,��I��~����a�ܳ��獞��p��
f	f�J����cGq8�yTF �p،ӣ�)�Z�(!� ӕ���/u��<o�E�+�[�$P�dr~�ꯪ�y�͗1��u�'�ِOVox�
��3�}/�oK�9ft䅯}���H�%��'~Y-f��c�>�m�)�,#���|c���������<;�����&u�
ӗ¦��8!�;�/���b�z�k	�P���V�����Mlm���e����SJ��F �н�:B�`���i0�yE9/a��	3,9���=gVY�+4]J.�%ߓ����`��l�:gI�[�-X���<�8.� $�Jݬ���J��[{��c3#'Oa��9��=��aV��
3x�9d^��׼FF�O�T��8U�����-Y�}�x{���y���ț������V�gj)��g�q�d��0Αs�ZyRc��{kss&$_�����/_l�L���m�Hl�^u�G\<��7�������"4�S��vo���]�g�X�ѝ"�i�m���]���.��$�*�o�p�jp1�`��RK��y��p�ݞ�A��ԩk�'�Q;̫f�{������˙X�^��{!��qÓ��K�F���ˍsSQ3���S�,�O��Mq�:)�~��Ѐ��E~K��g�56I�F\GwFWdZ�Ǹު����:����e<[fc�J��v$���J?J8�/�Z���4w�4����C縏W1X5���&�t�V�f��N^J�Eof]���܈����b���{�0SݒQX�a�Ҏa��,��ڼ�k�1juh��5�s��t�>F��;!@^n��y.�5[	m)�`XQ2�=�
y�T�)��v���\V`��l�PVt7\&�ͨ�7�_K�ݐ�Ԩ�ѝ�M�
t3�e@��ۚn�=�5%��X�.�����gY�r'gC�+	60����Yۗnڢ0�OvĦ�#��������a��[y���9>�=��,e�Im4f��~�����T��%/qD{Sc��4�3 �K��NF�Y��a9f�3����ǆ�I�c/�j�,(\���t>���S�-��0b�gh`.�n
��n��]b�;9/�R�D��/C3�B�0\Na�Lxs2R�32F컿�r��ȍZȷX�a�Ȯ�&]�t��l|d�HJ�*�qѝ��a�b� ��i|6�ew�J�5wd@Hv-,�v㦕�Fe/��'�����&qn^r�c7�p�4���JY#2�R�.�!R��"������v���Î�һ�L��m��pX�0N�0�rc��ެ槩L�)J����*�4����f�Qq��΄Żҟ�5�:�t���v6ŝ���I�#J/��2fW#��eJ��1�et��e��=RI����ݜ�LB$�dΨ_b%.J����G��b7n.Z�ZTU^8�T�h����Kj+-(�[F�c��"�e��h�*R�ѥ����*��V��-������j����F+�ڪ5�y��
�a��JU��S�ܩm��Ug2�Z-�YX�닜L.�3m[5����e�ZZ�iU�h�ˑ�n��Z�\�̸��6�V�XУ[mk�o,��ݹ��4\j�[b��ږ�p�ʘVҴe)���iJ�ʳ)mF��P���e�(�@� 5�~~{1�f���L��sy5�c1Z��=���s5����;��2�Ғc���
V��#��������Y���"�
��FH���p��ulJ=Sb���<!�#�87f�OKXn8�n���T�}�1أ#�K�&+�%��E�#�b�a��X�g��s5.N;yM[{�����2Q92u%eN��;��O�U���ĭ9ӷ6#M�Poг4Y�O�TE���Y^;�{c�$R:�]��$���V�o}B�6�'��ٻM$�C�ogi�㎝f^�J�{;����v4g�c&B��4P����#.���Ci_{:�ǣ�s	z'N��Rfj�Gn}MGLu��/>Q6`�����ͲN�{�F��ɭ��]�ǈ��={�͒4,z�8X��W�/�ˬ&�
�z��\�t$bn3�_W��'S���}2���(�2Lwox��=����$�|׈��2�WChT�~=����Z^з�pI�+���+s#��ՔC��N\SS{�_�hg@�k���JC����Z^�5��MX��R<�<�2]yb,Z�y���9�{DK+'����;���yN#���S�<��XB�r�@k=2�X�Ks^9�|���P�X��;/��^rIM�э���Q_0�.u�ܩZ�β*�O3�u�s�ښ�]Y�J�����hE#�boo+<�@2�B�@�lTwܜi>��wn*��ZR��<R���)7���Ei}��9P���}��4�IFS'(���U�"��6w���a��7x��b a��Q��j�YL*���nf�d��}�;��ף5Ívf��}���c��E�Ƴ<��|U"�$0�t��nvL���-�,���m-n��W�bx�9��^׆{wh髏#O�Y�%�n���Ӡ'7����mLY�%��e\T���}V�u&��z�~��?[uꈔv^n43�_�:�ޞ%��)0��'��+�J��e�gU�&��K��F�Gy�=c�t�&;��X]����K�TYp]�Ub)=��7�:�(��[%��$W��
�����p~9
�����{F�D����Ԗå}<Y�OD�X��(6h�6�rZ#�2h��{^'*�mW�T�X��@B�r�Ի�z�&��Q��O�Ө��0�]�3����E���Cuu�s|$U�r�x����4����ݮ}�u�p >��A��R���
��L,d��#g×+x/ivy.���̮3�&������D���fz�{wp��^���hv�'\����4�n9�yV�^��<+�F�ᱲ��.Sx<�m�\1�M�N,��fE��V�b���#l�j��8^�Q�瞬9�fey�䌣x��8
gf驌_Z��������&q��Nj�3�����H��K�0�}/�� ��D��U�Nx_^Eng��<]C�G7�!$�@�{BCѝ껮�P�;����%�
eg�Q��$V�ڎ��r�i�s-���H�`�p���';*e�6_r���T՘GG]W�b+}��,���[�pw�Q���j�qw]�E��,�ͮ�.�x�������ٞ�j!�Su����[.���Xg�	�\��ثZ�u�o�-=Sm*�q�Z������(��Q� qd�lV`��+] ������Zv��:隷�MU��
$� �2jOpj�i<��b�3�.�x�r쫙eJ�*Bq�Zn�˩ؽ�]�W�yV�R�xxx5xҬ��s8}D�mH�k0�u����ڵ�o�(x朕薬��0���h#�s6}w���h�$B������N�of�/x�=ڍ�u��F����k�kW3=�Ê�q{3{�硓n������=���%���k̪��k��eI�ky9���K �UfN(6��%7yMK�����q���$vē�<��T=�����C���Yy��><2�br̘̬|��ܷ�M#��;��8��;�������œ��I+��vv�@(zV]�V.�uiܛ��'�)�{9��\��R)|=�xi=��;:�k�P=>"wz�*��@Ң�8��� E��k����+f���k[�P�ۼ"A�[�ʓx�S�R*����:\=r��r���X4�a�+58� �3�Mٞ~>=Z�r��ex����|�l�\�[�.˧�46z8���P�V����Vmn�fj[t�]1�B���ȹ���[{���fw�JD�.*R�5�/׷ޝ�a�=<�˚ը��W����@}^�(��Z��0�Ձ�z52���
;�]���H�E]h7���MdY��:�β�� ܏	����u[��EL��mw��Pjt͛Ы�]1�΀v'
nO�U���*L�l|7;.x�YV{!o�H��u�v�fU�i)9�m����كz�e��ꌚ��A�\���=��9��s����'pE�[�<��N5*k�P��CZŧ!���y�����~T�GJ�`#����� �]�7&�Obh�w��i*��65����KW�7�qV��w�������Xc3ǘ��ϙ��6w���E�t*�'zGr(�>�ω��b�UϽ��rk8�Oa�7��J��W@�����mZ���΅ԭ�����^�yK��}-��<�s�t��s�_e��i;L�-C|��34�e�ۈ�I��4\���O�}�{�%v[N�k��
��ڎ��T��=���a\���Z�L�u��y]*B�����eg[�>��+Ul�*_V2\�\:0x��Ռ⇇�&F�,d�n���8�v�M��nF��F� š�k�>�b�4�ӣ����ж8
���4s��0X�}���j^�hV9p����z��������W�V�5�5g�(΄��N�4+�m�EÏ#&'�Ɏ�
(T����1m =�!y]�s72��(�-�S�Ј�tr�L��bq�����,�jn��pwǝ0�4����CCY7g����<=���:1�$0h��\�PU�w$��	z�S$��n�r#0\���#+r�dz2�OjPUԂ��s�5y}��znM�e�*c��]>�9N!�ܜխ��&M�أ2O}U�{���ۈ�F_1��y*&=���iQ���#��[��re��4y�Q#G�97�n�ڥD��H�DhCe�g��\0V�5��a�����ᢔ0a4h��|���}j�~0W��g�m뽎�����7�SP�Ţ3���FF�t�26�<�Ӭ���:gOP��H�f4��ᎨH���EÁ=@#��
��6�e���x���� ƀ�����||.@�����ZҎ�Oi���0vD�;#n���,B�����6z����\����4{�0�`�GE4hX� S~�S�����+ݝN�^9Y\��!�{���~\8V� ?��{���hˋ�7�"�<V���˨�u�}�f횗w���3��uש�8\�:�Q])X�H�;Q訃Ooa靓,]޻Ҩ��bhj��ۧ�������(*�N��Q�J��Q�V�`��ݾ\{�f���=��,�b��w-����"�b�fj���3"��[��沕	ז&�@$F�^��2+ʻ&X�۽�֔����9Vf3Д5�%F��!d��w왓��γG,;fc���ޣSx��� ����̎��KB���N��S$��"�vgJ�g��T�JWN+���ĕ��oG�m�ޅ�5U�X���U�����z��^Z������T�y���H��u&�i�m�Q
��]����1�i��^��(�q�9"�޸�c�3�����Li��|��h��$]�kmt�˧xk��V*p�D*IT��i�b`q�|^�I3rB/z]Ŵ��˕�R��x�y��xa�3�\�PK7oQ�Tُ{��te._ItnT���:�� 6lйa�r��v��Y/p��M�r���q��N��8eG4u���ڎ����񈹵g�vgC����A�ˍ`Y�:�|�@����BM1���ԑ*�]j�0\y+Y��Oq*]G���:������y�m�j��u��(i�K� ����B�V*;]�\��GM��T{KAy+*S��g�,�د����[Aj�qD�q��
݇1J}fg8F�+d�+�٦9TR���WB��ϳb�1B�6;;7��`9�����V3���	p2�J�&d�B�����)��;��/3������f<9�;�λ��-���ZZ�F��+��51�1n���h�K����ʍ[J���Z4G0�;h�%-l�ac�Ah�(���J(��/2\+W\r�UmZ%��kRۗ1�6"��[�0�R�m�-3�\**Z�-+l���lq�6�JR�j�.cK[cCr�\�-�\s-�ܙ6�,QZ'3�E���������p���+�mN;�6ڋs3w1��TW-+F��������Uv��m��i��+RҵF�+�x�)��b����3���=�<��I�PWf��t�I,"�E�QU�Zh��R�� T�Kr�_HQQBNرS��(�9�[��.(l�Z	�-�&1��=;ݣG��`�>TF�cW�H@�ʂ�U���x`;�"m��.�X��R܎;/*��*�ު�׆�����Na�y���j�Dm	^5��]z�R%2�ʓ5�x�~�3W���y�}ٲ�� v4����������
x��{Ķ�0�E���� Fi��8|���䨢�y���պ�+�*�k����T�����M)Y!9��ۛ�SD\(�Y6(ɅN�}��cnC���S�3s�}f��H�
@�٧D�Z���X΀6���r�=��wnx<����0h�RV&
#�����D��ɺ �ye���1��ɂq˒��Ǜ�mu�*rR�י��Q�� 	�ʼG�"k�$��J�xe2��B#Ɉ�G��^�T�YZ�+�� {�'�=V���� �����c���c�p욫C��Pܨ�n�*o���i��{F}AC�;[rtl_�T%���M��O;GO��2�W��ʳ[o�UhU�[c�Ë����*`&h�_�@�T���h��z�p@��]嗪���{��3� <6,r��@~4��`�"'B�Y�S������tW��t*&��ʞ�ٱaʊ
c$VK���qR�Խ��bA�`ÍRa!d��N("+(�QiɅ�^��BṊ���$qE���x�Ō
�� Bx�o�s7�,�v��>Z #����(� �Qњ@�l��[y��O\�^���׊�O˃҂e����>��pZB87�N6=�����S�YS�dK+d�V�5�zw�P��e޴OR�O�B��>���L����!6��z��Ȋ�j!�d[��l_*�J�*�+w�_ <<�j\݉}7ܘ���n8eЅ������#hYv������췪���tz���
��h�X:�
�ŠO,��6�;�}��iᏔ
��~R=+\z��°�g����������,G��u��thZTTɁV��^�7���� �n6S�����A���';���^uS�Y���T�1�������7�k�ǻF�ۗ��}�Ҡ����DB�f�������?h��X&�V���2�/�j�ʇ�P�3#}�b"��C2����S��Gr	�ˮ�X�F���X>Utx�W��A,�������q�{ ���V��]5X�Փ�*<�:7�g�Pý^�3�Bg#ˍ��R1��v��:�Ԍځf�l,ݥ���`/'"��u��IxJ����t�f��vvV��Ƚ���G�����������>b�c�vר�٩�JT��1P`�$Q����1<�}���o2�<�� �el'#}�[��� �a� ���9qU�{ޢ����"�*^|�l��KM����s�_x��,o��?"a���U՘���u�}W=���I��v�HN���I�*7=P���/�ŞGP���y��}��6W�r�ZڤL�5�q��:�y{�g�j����Ls�X,:�κ�(�e��;� ��h<x�21b�zB��p:���z��
+�^�9pL����h�UI����oj��ˎ�.�t8sۿ�=���>�7v$)l�X�^P��y�ZMXc����>����4����q.�/��A�����4{
<9yi��q��Q�h��֪� �,.��"_Vw.��]K�����Ԕdlձ ���̐�1�\�����_W�/ߗ�֬߿t�,*�����Pg��d�������G��6�|�����iG�>��'��h����P����[���3�}|��V�cÄ�L1Z5p�վ�J�gt��{~���
 ����=T&�
� Ŏ�o�TP>�+�h��b�\8U�h������pkr���)� �_��EH1�<%FEÆ�Fm��\��0�D!�ea��l�5���j��F:(.K�8g.��c"1:qJT
B\8���sa�.A����[-�5�
��"��<�l|��,Vu�@z�sM��~���U�\*����U��H�p^E������n�=Bߡ���	��q���(�k6���f�=wtB�ySQ�����1����vJŝ8�2"��:�}�\�SF[�6j ��V��xp��)~x ������L�&%���X�)׭M�����	�X�]|�����SƼ�ҁ�-����q��p������wOL1}�9�0�Gx����"٠0v�Ӡ>�[�?/\��pႬh�N�0�����JX��^A��_y=C�x1�4k��pu�:5��*i�X����v}:* �]�`���x�/����a�����N$�ݗ�'_� �m�GG��۬z)CZ�e�֎]�>���f����n!����FP���õ�9��C-Ǜ�9�3W��X ?L\0B��c��5�4D�{Ǝ��;���P_q�\5����C���5)�p|E��s���)��F���"�<@U/1�TY��^�w+ ��H��oM^c
It���uj[/�-J��B���Fp�����Dۘ�In~�}�}_9�?����g��#�C�uPgÂ�:x�����
�[z�b	�VӬ��\Dˀ�Hq�
E�b��ѣn�C�ceʳv���r����*t���+4!�t� #�4����cŤ��<�s{�%���E�n�+W/�YT}�A�| 4��y;7&��Bd8�72�=����;�s�c\�,8=���c��W�\��!Q(����{d��������i��P����X�?)��PC_˅y���G�w���p{�����6���k2���&߱%@lĎ�j�v=�Ү�&->� �*��]O}h�c��G��h
8(߶VV\����֨���}L|��hwǏD�Z�q�}$�4��g5����>�BG'p�[��R2�X��/M_��Y��ط��(VCM��x��j��*Q�h�@dыc�Ƨ諭��7'�&��ࡆ�&�\�#ʰh#�}��J�����>S�8�&-ME��*� #����yAN��=6v�){o�s�`���ަ�*a�V@�R����lC���`�.��v&:��7 ���`���xt�t����H����=�>F2=��ٹ�KT��
U �Hc��>�n���� 1P�@(p.42!˷B#�� �Q��*����i��
���|ͭ*z�s^f�� Q��m�W�K/�vY��C��x=<.���iC�yh`��39jklތ^T����]H=��v*
L�ƨ\L�6�`�PU�����Q�0n�%i�F����a��m�TL��P��cˇ䟐�!�F�ɛ��_l�MX��[���2����/����OY퓭��CjcA�\���{iE�f"r8��җ�c��x	E�?���nũ�����[=ʽ�5�C��Y�-�[RM��������lT8�Z�>YR�M7���W�^�|l\C"!C���U�yD@�:�.�v���2�b���v�dlt��f!ǲ�\'=-�A�{���@���7`f��W��x������ww3F�@nB�y}	�
8�
��$1@] &y~>͓7���*�<.�A�
b긱 ���H�h����� ���n�N5p햵}cE_��^t�G��w�qzLDtz�tL9T*xe��A��N-r���Q`b�z�w�:|�xb�'�����x@<k�h5�$2&,�'6G���9�XTٍ��M;"��lL���U��A��9�$󻴔}p}�}����p���CoP��K�����W�x q�����$lW���Ab�*��e̡�v���n�헢'�N��qp��p�!9����3W6T'$[��ˋ�i��0���7�!�@���j �b�LV0����{������
�x~}��D�3�gC}>}�Va��e�����L�wJ��T)���B�؎��iOUNr�>���]W蠯;T�KO<�W�����������`W.����X��d�]���ִ �PA�c��3������>i�����u=;���9m�{�� >�{�v��tm�F����0�vm�H��p�P��p7�Z�RJ����7��{߫�Ђ\fv�G��\t�L�#�������C�#�X�S��qNv��/��t��dj���V�W�$�.B�=�J:nX��M,���;�fΖh��xVrTGd����G��3��sTv�'q�g��%yَ��6�}�Jg\_%h�S�.��$�E��ʌ_X�f�!���^���U��.j���PB���L�T"��H��V놓�;�f������m"�SC@�Mc��5Y�\o���ХY���hs9�bmp�ՆslG-�t���Ү�_b��W42�c]��\vb(�UD�ޠ�H�&( ӝs��]\�b��K�O^EV��v�@�L���W�ɝ���g�ojhf1e����uH�Zփ���8sx�v�*"b�Vp#6����[W��Ь1��$�]�7q]kǟ4��x�ֹ�v���IS�s�����}>u-W]CO4�`u�5��'Vm�U�qȦ8yZ�.|Ĺ�)k�k-��D��=��iꗻ��z�Θ��R2,�;WGt��mcY�|�d�1+�+�ӖS-GVfZ��hP�Wu���С�Y1�����3�Gk�Oq&b�QFh��N,ݭx��*�9�]�hv��+�2&��5�2lZ8�6��11W�fh.st��88oE.;�,f���W~����ũ�1���
�S
�v$=���R�����Z�#���on����2��G�ާܺ����_+Y9�`�l����ȫWԺ"�S�%�+.��oE]m�X��zÌGӎ��m��	���2�^1|�l�$�y�]-�x ��u@��'|�鼪�����H%�u�Ԑ�U�'�U��,�/�5eu+t�<��lnp�@��"����5y���%ީ3&�d�����I�`�X���m<w�̨�u���eI,Cy�����Ҳ��e?im���P�ۘU���Pw7w,���Y���o�u�Kmڪ���ј�,�Z���2��+��r�ѭ��C��MTY�&[���-5)��s1�����˛��DS�`��p�eq)r����ZU��lv�K�ff�wnfr�v�.L�L���6��U�ih�r崨���,�J�3�o2���[f�\h�V���y�ݚ���+��,��9�F����.7�`lE���8�,mQ��r��:�F���w
fUJ�Q&���UT�
�R�����J��y��*��@�/��������>�mr��f*�wv;���\ns��n�E\h�.ܟ�� 
[�Ӫq�Ɉ���=�R�j\^Hd+�Z)�SDG�>�����۞�
?^��S�ZC��%�F
�0*}	{�4m��P��o�C�Z�BRf�xuvf��/W�
��Z��Wv��u.��~<��CW��2�.z�S׼p* )*�0h��x5sh�S�¹Db����ܳ�=��P��4tW�pц��G@^_c �']��	���'�f����n�Jݸ�#�������2���8��v8��qJL5V@Q㣦��QB�Pfs�e-\�ц��H�Qbɩ���E�Ч���	k���*�k�q�U�}���P�Ů
���
��Mj���,��u��n)�Lu�N����uS�9�W��:V]-��R�AfJ�T�v|�ƹ�-��T�;�.ǖ�$R"�v̩�.�@q_I�*����ON���ע�g@�u������aў,h���b(n��@�5;W�� ��� ч~U���R`w	1q����g��g v�@ͳ}��ӣˣ
M9�}�;I&�F��z�c�G]5X)��o��txX��o�C����x�܍4}B��Y�����*TM]���~����w��>R�ߠ��aߨ��꣧@	^���()qu���{=�R�ǝ��R*a�.�^����2z{Ӱ������
���4`���:8@�B�������W�E���i��?zr�O��ᣇ0k��.���R�.TQXu�!�
[��BFw
c#�!�ܲ����4��]�F�,�E�u�Sc��<J]9е[�*u���U���s�5��T�Q�9�JӁk�]4��S�N��S��M����\���{J��5����%�j`�} ��AʎQN����B{�Hxk$U֐>��� Ԋ��h8B%L91nLU�Pc�uP��!Ɏ���v1w�t����R�;�U�b�r�@��R)m�p������|�������Z��?h@���\6a��9LZq���\����p/�8������r����ǻ=9ж�kr���*�P46.F�.)��:՘p�b�%�Sxy4�X�G쉆N�V��[AUC��0V�R&ESm��/'�@g�m��N�G?����K�8}���B[���?v�K��
�V o |*�_�W�^��-�;�w��)՚�����X)
P����fgc�ͣ��s)x�W�3�3��;�r��H-�����23D十�+Lf�-�ęSk�J_x �^�n�~u��R�ƹz�vS�j���
�Z�טJ� f���O�����μ�P퓧�+֕�15�~�p:@���Zi�3�xe
�'�r�fa[=/��ő�`yD@KQ���</�@�Jz����*5��!�PL�"rI�
�5�"��ї�y����#b�&��f˃
�%p45�"&�[W9q��&�@�.v�X��Y�=��?b�+ݍ[��s���o��-�4��°�?���#t�U��A~��{�~������:��c �9е#�-"X38������qb�֩�4���a��~>X��,�^���f}���˰.:��ժ�����໩gA;��&�ŗ��@��m�K\s�J��N�6�_��%�����5�7�}��Vn�H[4��`sUf8���y`P��j�C�����`Ѣ�,P�y�19�_�{�J��n��c�ǅX��ӣÆq�(3SA/_;���k&�w�,V�6Շ���'v�=l�߷ٿ`�@'�:$} J/ۧ  �O)��������,W0T��{�j��xJ�r�
�՜�M�-$��)@��2����+ ��j� ? ƌ�
Y�/[4LLd&*�W�P�pL3���I���8��Yy�ލX��,��\$R�Ϳ�؂@@�wW{>ι�ʲ/��@�<�ֈ.��
�UT������랾ˢ�~Ƿ��pz�Q60P[���`��n��{p�h1XJ�řݐ��m�s��O� 1n*}R�b�z����;��'ﾯ���gg���X����矟����CS�}�� o�I���n�3D��3�4���P?)+|~�{7hh�z[G��>�c�W���+Ё^�q��҃�b������ܛ��D�]���Wk\��}	��"s�{���b�x���Y�ߓaя� gD�ǓSLèB2�e��3W&0)�6;�R�A��ۣVWs٢�%�=����dt0�H��H@�U��eE���K4ǐ8�c޸xxV`vn`��m�^�dP�2t8�@ސ���x�nh�����~P�������T���ܷ�L�!rx}��g�9ee0��� �Mr�F΀���xX+����J��`m�Y!�7HF���r��V�kj����b3�;Yy�߂�9�|��������}��Q욦.��s�{� �ob6C�(e��.�A�,�.5�/�j��u����z$S�}_���HV���p"���GB����ԉ�tV��;�cD�1�7���X�\�
:tj5��Ҝ������4d@qs�Q�ź�&7'�����PC� �����l� ��~���4Yo
�G��� �ʷ�2���v	u� *�.���m`!��xl�Ht��	��(���t)u�ũQViE��W�y7�%ъqBoF-�Wȵ��8�P�Pu�!�6����"GJ�Q1�g��;��yHtL��Ō�Qjr���>1@���E������_�9g�wƭ��LO_8� F�X0:�()��Jsi{�<�����+&����;A
�q�9@3�!C@��Y�U�ݽ�A�4j���jK�a�^����}b+2���*T봦�F�+��S/�SF>�@���f��*��z9T5��"2N���Ar�MÌ��8Y'���VҫdK�P�T�\B�]���^����zfߘ�~"��Pߚʻ7�l4��AZ��_K�z{�Ej�z��1PT�X��®���i+I�)X��ϻܔ�"#zwdQ�Ra���>�b�]W0F�h�q�n��1��(L��
�����1� ��hzwO'�La��8<+C� ?X�?��*�0d>���]Pڅ0��Sن���n
v������G�S&Q�>C�ګq�pM�:׍\0VО9�飔U���N���!�6��a�(X���5�����"���h+5���ɪL����Y*�y�����]NKrÃ��{7��Q�#%��&�x��X�t��1ap����!�IcJ���X���E�	nO�}&N/��y��*_��iP�����Z@��i_{�Y �~zkLW�僢Z8Ro�%��c�8�!f�ⱑJN�����yXǯ�dӣ��D�`ʳ��g(PGŞ��C*�F�4dg�r��"���)0C��>�ogQg5Y!@O�t��i���UDѠ0J�X2M�\��!��>0�Z���N�������0e�
�l|�q�,�p�].͸�/%��xP@ڽ�2\�qT�������en@Oht�7h��Ji�)6��(��nc0�-��lj�6��ڻ�iX��|��x=d�gik�����Q���O\�7�Exȝ�1 ]$e<�~Кk�̿t̃^e6͡�ac�X��˴��ݨ��7I���u��k�+���	�W`��8B��g&KoC��i՜�2E���$�.s�c��S����5;�3����~�˓~1�O{�����#�KÁ4V�*��j
_GǼ�����2��!�Ԣ�cdVI��"r�p�0s�B�D�o�ؙ��� �
N�i�iG¸V�Bʡ\MpЏ*��&����6f犪��� !,�ϩ��N2&�N:#�8�f%:�Fǟ 81����I�i����4/g#�x�D�g�W@�W󰃫�R<��^K5G�y���v��ƴ`C}�R�������4�g�
�D]�^u����ɬ��~"]gwh}�X�B��l�8|�q��m����PT,U�~L G�O-땏���U��r��ۻ]8u�<V���i��4Vz�f�U�8'l���B1���u3z�Vijڜ�PKgw}h�������G�cS�2B>��˦!J��h��g���(3�&W.��ճ/&E��	re����d�k���lng���̬��N�P�)]#�o�<�FN�E�W��[�4�mu7]��]{������ވǝڭ�����aMR'�r̴���F��C��n��T>u�,±���Vs5:9u%b5�;f���]e^ф�4���\ONJ��R�B�4�<+���|���6X��Lǝ[��[̻�
ώ�2�ͩDg}>oM�F��{�n)ELz��g�{yV�n�PvV�)�z�"�̜s>�MW���¬I���٦��\91Cr�wi)�M=��F��l.�vce3s*'ov\����aWT�;^Q�STH�ζ�V��]N{�f�N¬�1<xn��\�n�G�Eľ�j����w%ܲ�0�ed��/qL�6м�J�U�7Awb�g)����c���2p���@R�J�@&;�fX�*"���l�HB�Ze٬�|�Ŋ!@�n
3)+F�������f�/1؅���$n�H� #���Dݬ`c#���j['�o�E�i��
0$5K˻C
v�P��Ŕ��BD�Joò�]%Pvwgtsk�T�,j]��;Btn��d���T�~���Y�v�dZ~���ŋܻ�U��nB��l�`Mh�+e�F�;A�q�Va�������!5 }�yoC�4��c�i�0ܩK��ݔ�sn`�Әt�^�3$�p�������<��W�h�����Rj��KB:�ټV85DW��g� \
ep3ɅR�mZUƩ�R�*)��m-�6������V�d]e��r��32��-A��3�V�X]s�6�1�8��yh�嫕G���Z�6�qܱ�nSim�7lYKf%E�fLJ.Ws8�9�ٺ�\������f�.�&5PܸV��*���v�nnd�TAu�\3*�A2��kGE�ij!�X5�G)�\n7--��9�E��^f��1b�J���76�tV��2ჶ��7sv���h�U��*"���F���6�&�L��2��3�,�T�|a��B��9�w�)�;�xA��#�x�\��_2�̹��'�Iؙn�9�hꒃx��})[�;��j��z'�Z4n�p�E9?�}��C"��S���S
��
y��6�Y~x+��+~.�V�b7%��l_s��b��t��=T]�E
�]^I��W��D�Pvo�b���עW�حU��mh84a4I���Xw�-��+Ù�/ʱþ��wQ�$;��%����V�>���)�P*|�=(����� ��E`�.�,g��y}�o���Ç�����rʗ�e�a��K��QP���5^��}�:m6t'���>�ʬ���.�o����G�x�.�*��$�����{��	�ȣ��~a��on�W�˩�6������t��Z���j�g7dL71{hW*�XF�8_�WZps����V.�T@���Xsm���/���(�}�#�P��V<�r�/�S�k��؟<.��t�Y=�IYקJI}���.q{uP�j/�!G}�Ȋ���-: ����6������ڦ�������������8�$F5{be<I���LЈ͜�B�\)�Ɣ8����G�qb��v��:�+�����7ZA�s+2�t�W�YR�.a6��O��y��j����X�˳o@W/}2��W7#�2$��E��G����v��Si*6`Ɩ��8�]�v󴥙Q<b@�Wg�24�u��6���ݽ�c�c�]���t�X��ӗ�b���zxU����4Ej�x���7ʼ(�fi�S�����c�E�q1��A�y��ݺ����G�("k��u���6���Vɀ�l�p�piwb/#b��3`H�1nS��	�*�ZN��`�9G�Ȃr4m,�CW�/zΨ�Ð90���w;i9�oD�T���d�e��*����{���;)0�A�b'g� tLXb��ַ��f�%^�udx�2^��h�Ne���#�0k�wAv���X���Ȍ�@1��RLّ�&Γ^��!��w�<`�:(!��>�
�%�#�5a]�>��������Z^r��pБ�+�p�ҭPڀZ~ǅ�9��� ���J�X藂�M�xU�oE/�����j(��x<J�1qaϲ93�z���nH�FN�s�5��n҄+d(%V���(+��ft�:�-;��tv�sц.�#�y��d-���*H�hYw$����˃�ث]� *��U�«���၌��P���t��Dn��3�4�h�@�+����/���md�v}�"�A�l���	�&��A��ɔ�&I�i�v�f�����%/�JoQrlL^�̏��#c�e�^߈�f��/`W9������H�a��ϭ����SCd������e@/kם�bq���+b�HQ=;
.���1:�����wxx�5����b�uMx6`2'z�@�I�����S��j�sU�)���dI�j*�
�JB���K�kO�#n_�����1/�}����Pz%���z���
�`���ɿY�Y���|+�|�b�th���xv��^��eu	o�K
G��+E�^?r��B�ʠ���|k�5���X��Ѯ}+]���P��s����6w;_BG u�>�0a(zW*�S���MB���2����1{f������j��ox`���oMn6���f��m>[���:���;�x(���L����]�-̇cH�"�2G���Ø�{~W�SBp:1B�3a	
X��jd8�5�c!��=/�`�7��8!�Vw�x�����*����0+�z�Ƣ=�J��K:����s��1yh7��>��~�>�j"��®�_�:�3�&:®�gc��`Q��9�N���g��4��ʫhU�|�:�׳����\���.��

�
��
�=bB��$H�vl����,�lxWdX'�~�V��t*�������o��rgwGH?3��	<�iѕᗟ1S)��wv�׈֐��z{R���|'�X�D�N�eQB�YѨ���\I�{��qq"�S�v��d��ug��k�T,!IjѴW����\F����|H��W��μw찺�{s݋:�otG�Y=�F����%Y��7�鞹�	��W�*���n�G�{�^�˦.}$@���W�-g�A�k�����c��7c�P��!۲9�G�Y s�@(lM�����A�,U-�k#9WH�JAb
R�*A��YE�T>vp��Q�e�{i��,�T��XRDs�R��(�4��s%�-kɲ�9�r��UŌ���d>4"]1 �j�Dt�ɴn�$��FW��/�6�tg���g� ����W�-j����;����"��Ј�o�e4�S�<iC�YCe�&N��^�B�\kV�5�~v�a$p�9��j&��yv��z{���^�P��M}u�Y `�~�Oư�X�Z^Z�z\��w<)��WJY��k*���mY�X4O������ɔ&�Ug_�Ӎî�h�rxQ��g&�V+�]��nq��:Yˍk��e^G��Aq:ի;5Vَ���q��UU%��$�μ���ꈠ'��:&�(jޏ��Y�8c/7�^'Ƹ����y`���
vj��*�p�0p�4p��+�n��*xV�]���@���<�+5�fFԸP�i�F9�-�I� ty
�J������_�hSʔ;e�_^S6�e��v&%.I���l���C�K��\Qީ�!Hno��ŉ���];@+�:���`��Q�$��7�6�X`��5V3�5�����_ox$t��q��a���уΊ�h]���<+z��<g(�f�׽���/Q��>e���hC�g���m�f!Y;O\[9��[Q
9�a��n�Tb�q��{}۩�N"�4;�wo���O�b��3��B�a��.�@i=�"�J���&���j��9�i���S�5vF����Y�bt�u%�� �Xۉ��fre8���Ӏ;�h�ҥ�E7}l�w۽���[���#�[�;A[����79LO��V�]���f� �X��{;Υ���]ȩP�
-��N+����1��X��E�ֽ�8_�`д��=��T�������,yYp�\����C�\ ��c���݆Bll>���a�Ơ�(�U«%"��s�X���*���G�O�H�;ĩ�㠪��p5�� ����b>��K�6���#��t`<��GT�;���W�@��bѳn�ܓ��a�D�,Wm������
X@5��01L��;ۮ��~A��k)<N�^(,:+CF��_]�
*��Pս�ߞ���i��nլ-7Bi�lJպFhX�o-m\�+�-����+Xx��	�\KF�؁Vw-�ļ�o�ΗRm^H��:V�)|��)W���}9S�blذ��H|Ă�e�t�㙂���9q3B�h��Y>K�i���Q�1Y1R�,����ǹ���DdF��[P �����/�^�mr/�sEІ�*��<1�;0cIð�dU�1rH<&kp����@;>��vc�$Ρ#�E�Y4&C�g.]s�A�{<�;�Ԉܣ	�p��Κ�ӣ wt��Sڗ�g|���ׯY�tPwi����\�H;W/m�@����q0���S���ѯ_LGx[�PF��P|d����۵���twN|=r:D�0bb�ɀԀD�W�`l���Y�Qq�z^mנw..��جغ��ۉW*j�=�L�ެ��x�K5�RW��Y�7W��ߜz��^��o��A�f����(�����z�X�4U9%�{�t[��H�s�����̅2���\Q����c��m��E�l��&���1f��7���T�{������^s�V�w,Z��W1�7�"��
]�Z3�Ŋ�׫GC��xh�'����S��78��[�Eۥ]8pORm( �UV[�f4�T��tp���V���u�#(����.���[���&�`
� ǲ6��{hDHQX�2�W�^K�y�G�4�U�yR�: �%VA�;X=��]�-K�=XM�chT�1P�$GD1�ʊ���Ӄ���V�b���́�=]��c��DH�,@�e�X�tg1��[���p�T1S��U�j��r�G���h�ҕ��.�z�U�0ߊ�fV;�L���VA�Fѷm��쓃wlU�lS#gv�U�ǞxpUհY��K��h��]'�-%1�p��=��6�GS�gt�6g]-Rc���4���9ݣw��Y��z�8�w
�TŘ�wSuY+�m%�NS��8����gr�[W�g>l��xƺ[�A�v$�i�#w�6��j��I�����\Kqhk��W>�b��F���e�o�ݷOj������DnT�b��B�fQ,�̸Ξ�}�M�ӊi4�9�y�dɉ���|Rz%�M�KvU���ʍۭ������������ݽE�s�1Ty5}&�f�t��i�\�.��|POo���,�wP��D7�A��"��A�-@��7)Q���B��l�H��ZgyN��i�tx1rn��V��ݩ��a�K���Sv�+�o8ݻ�C�bdU�y�a������+e���	�+�B2�^� ��#�3Pf_�&)�l*�+Z"d("��g�I���jȩ2��G�l_�����3C0;r��x�	PP���ږn�\�0r�����>�Ùk��ТCp[�"d�<�.�*Xk.�Bae�*a�h��Qj��v�u�1�n�خ�
�YV��*�X$�+	>����w)Lˎ���P�WXrI�~j��8J�0l��Ӯ�������.;�Ԩp���	Ceѝ��[PS����mm���f4l^튌�+p^Y �xh�kS�@�y���9��d�S� ,8 �lzh�G��R��ʆ�"D�*�!2l9�2�8���Lmr��2e���tc�`��͍�2�y�(�|
E�"�U�̘
Ĵ��N&0ǉ��U��yKR�*�XۙU��eT.ٍNs3T/2]�l�2�6�-C(���3�.8*�ܸQ��LlZ�mh�;s
c��e�j\E��eh�ͭ�*0F.Һ�q��b;�1]U�cXU+(&���dv��2��n��52,D���r���������7C1na�q����V\Leh���b���S9a�۹DF#�*�-Ll�*�E7)���L��L��[-aZ5L���6k���3l�-BUF�#�5E �vi6�]�v����N�]KC~����j�#����V�W�����W4�kc6���v�L�7Ƭ4tS��C�*��,m�u��V Ѕuq���g�j�FW�X��>�ըn���ĳ`������p�t��_�LWe\\�B�j����=��]z"��\��CzWN�dY��X`�X�7׋��Ӗ,ux�x@��F\~ϥ�H;�D(Ls}�eb%ž�s�::�:'\�l�/*ɫ��F�@l(1��yk��kh\�P��͕�)M)1P�t`6$IB�׉��(w°r:+!c([��u���voy�|�s3����fDÂ�ARI��>ڑ�Q^�B;x�6��:9�p\j����^'�i���k@�0���k�{�	>;wL�s�Gڞ��x$*��2��H-���μSη&%;m�I۝&��^��-tVM��O$��d�l��3�*%�NO��UT��ﰑ�����pI�]#�B6A͚<Dc�f�E�23���S�PqEЛ�A��5Ch�9P(�B����m�\�H��.��5<d1r8����F�%8�{��m�6�j�̠��s���0�U:p6g��r5,�u�\[8ڏ_��b��.N?����a�c�v�P�g]a�Um6opT8W��@��k�W?���Y��J�)<���܏sԺ���qq�b;�!�v3d80��^!�����P�k`�|���𣖴�<�/e�8`�)��6gzI��4���D	��z�����ǅX��y�^˞Վgx�����f��������b������i@{.�P�N�3A�7��e�e�%X9W��Y�|X늓ۦ(궮���|��v��qՌ �bee���-%�͓y�ԑ�d��U�������5�����:�<4@Eh�Á�	������Xu��R.�C��ҁ�#��y�^5�aѢ���(UG���y�軅ǾF�ipႧ����q� $��ƾ�oq���σ��H��k.��0�c��1� �F�/�(�h��#��\ix��!��¸@bTp��;S�����B�֓��a��ފ���sNB���t�V��RL0�K��΅�
ځ�QV���^\�����fJsz�,���V�#���<ke�1�Ly�/�r`ͭ��܆U,LQs��dE�J\(�6��*���k�f���;Hw��#SOE\x��J��z.ly/q�X6�@�:�f��{Ձ6W�R�;Ž��2n^���@S�j�d�X۝8��j`�1Z"���$ו�Z�G9Ԩێ�Y�\-�?W�I<����_&!��D�\)�Z ��6-�1��0+�LU�]�(�3�����bŚ��Z�U��T�ќk�U���מv>�����>v-X��u�;�]���ɯ$�)�ɐ���V�����5��S��ңr6=;�s!qM����fh\��"}�^	Z~���C ���T�����z5�EX�~%XMX�F�l��~k���:x��u>��'f��� �c�iqB��{��P� ��C����C$�W^�V���x%#��xVm�e����l��y|�Í���p�#�x@�JpT��>�2�dz�ñf�.���Z�zLdpEc$}HF�\�4���%!ף�#�B�M�}+ۡ�g��W���������=k��$ެ�κ3F}$9�Dᆠ�9V	E@�ٕ�{t\��.K�缩l��#���E�9"�Gt�1���^�V�;���Q0�H�>	+~��Ä�ӡ��zxP�.����=�p�KS<�c(Hk��T͈�Q �2My�Xy�%}܌���h�~�H=5(x`p��Z���vnɾ�����h�j4ޚD�-5�;��������tjt�4��h���)2Ҥ��0P��b{����8jZ����Ar�@{���1Cr�,L����>>� T�KC��r����3y���h��0_&z&��1N5�֌ ^��T�th
b�X)W��1�o{�矝^���%bX�S�^Ь�/��`5&���r&V=YNZ!�]�t�q�]�Rv�wZ�;9յ5�CUgCs(��0��E|���֩�m]�TE��ZQ_xx�_6��{�B��b����Gb��g�YF�d�3/��
�㢗U��O@��@
��u��*�F߸˼K�E�<��Z��ζ�飣|xv|~@5�U��"��k�\mAc��>:�R�7Lo���)Z���Y�}�O+��XU�x*��*�T,��kB�5��t��������S��&�T���"+(�Uǎɇ
�q��yP��6vQ���M�[=	L�M!��^5\7R<�Vn}���y iO�T�xVWL�z���g��P�^ ��,�<>�����!�sQ����E,��t\¡l�������x�A��ԣ��G��Į�b��K:]RJry��߳(d�P��:�.�S��Cra���j�]���>i���^Q��P��ꗃ�yTV��2V�)}�RٲE�s�����4u��^1� ��9ƣ<�ka~��������`|h7y`u9R�@
��ҭ�r�8���,�<��u�C�JL�� �]�D�[~n��o��A��k�� E�U������j��]�[�Ʊ�5X�3$c�5�`ǆC���: ��#��E�^�F��yp�5��E1��4�Ы������V��M��Ϋ��A	0`��X+Q���Ft@��v��Ɣ�Cj���C�8m��ઑ�__�M`�Z0�����x�b��AB�Ҹ��_ki���IP�=g<GgL��=�x����6D5��0Pj<��i��7�ʟ�0�&���`�⩰���_fu�Y�x^5R%}�����R�T��Ǖ  ү�v�ֺa��n^#lG�.�J���ʭHD�|[Ru�{��ȮjoZȱ������Z�s�4^�֡Er_{�;���A��(���6:,sPSN~UW��$^r���{o��*����٣A��gG���_�ƞ�[�0����T1�QqP	���4h��z�<|g�J>�77];����wF��"�Y7�s�>�U�=��	�#6�(�t�ZG��I��Ӡ
c�Ts��Ǯ�����e��'�I�5`�e�F2�r�,��;v/% ����=}�i�k���3�΃��~�!�
��-�;Bw>vV�8�g޶s��p�*4Z>�� �N��l�s���6��_N\35�a���h����.OO`�^[�vL�s�{�~�'M<R�Z�6~��/��u�J\��	]+�<v�K��J��,�>�b��/�}�M6ij�qf�_���ҬUyq���CC�n��f X��O��Si�v��^9C�<*�K�hw�+3M��Pz��]K���sS<�J�_s������(tI�S~��f�E�]��W�ޣfر
1�\����.�JYs���R~�$r�'�eMB����0
zӶ�vW{6{�3Ơ ���T�'.�O'ϗ��kA5�R���c�(lY)������x�R�����4N��3Y�%�pৼu7#�ί+�4��.�!��p34��k�p����t\���D�l�v�ћ")>��n_U�'�:�i5I��eBo������.�0bƍ'�B^���%����g6w����=,�w2�DV6�Fז�T�c�{<'�x݅�2��p��*�
�Qv<�o�x\���2$����TCEf�h����U��Nd��ުz`� �%������A�<I�W��H��N<��H:6e�nek�v�YP�\eTzWp9��I��70��<f)Nm�\(	���c20�8\�|�qt6�*�MY�n������{��Ec�6vӕX���F����|j�#ZWQ�'%��β��E��7 �a�vRt�fI+�HNX��%]��"�g׺FV$a�����n�Gi��V�O��򫙃:�O��P�����ڻ����.�6Jw,mѾD������5��ܾWR��[��m%���N:�xtwK:Ͷ{/���{Cn�A� ��.}�L�v�o7�˳i��2����Փw*�3�R&�k���R���ʒ�=�qA/U�W�1'X�M�9�m����Jn�����˷�1����<��]OM.�O{R�ZN�X�nv^d!^O���	6�|n�Hv�Ǌ]�q�ÙG���%���ӣ�b?\̭�Gtǚf����[ֈ����T��$Y��ZYYm��Jn
�xm��"Lh�zO��¦��8CM�������&��{Y����վU0�%�6僗R��x�N����*����^Q$`APs0A�n�
����wB�D�7д��vr�QKt�+0@#YCDP���JA>��+F�?o�jG�Z�Yn
P����lfŒ�J�*��fX�0�	�%R�ʀ2�!�	�n�r�3R.�P����Kh懒�d��N�M�4�������l���p�.^EB�W��Xssp�x�=��eѼ;����[5��_�]�`�BKt�7�cibo���������:2�H��]��;GQ���N�p,�^�\����� �U}�����1��%fZPGd7Y�V]e�Հ*��|'2�֛�q�8\����m�nQ��k`�cm���h��m�l�3TiGr�������:Yy�R�eichV�F��Q���-�,W-Mh�3��J�Lm��(��Jյ3.5�Z2mƩq̣f92��6��fZ��*�q�UDxٛ����pEm�����ŕF9Lq2ٍ��ƪp�d��YZfU8���+�.\�#���n�32�m�Lq�(cDb���1kS�8��m-�U-�-YmQQpJ64��YDPm�l�m��R\�Q�8��ZV�q��!D�cVѻ�ʣ�?u�Cwq
Ӛ&�t5BW�{jࢶo��K��<G&ͼ�2L�)bQ�y���6 򵎭�r9d8��E�Q���h������54˻�O�r"��;�
}�Y�f�)5��=��G,���Z������3M+2i���*��no(S��8Yp���m��8���Y�E���]T�r����3:��E�:�6�T�dU�W�E�!E��uWI�zc��*�fR��q{z�Hen`��Έ9�=����[����%1~v�u]�Q��ζE �7����ϯ�yuk�[P&�w/��[H;o/W����M��3��eH�ܭYj��kr;����.�tn�\и�8#n��l�%�6���%Oܻe�����>��'R"�A:+�B�\d��עY�4gv�����)����M�����Y�J#ב������Du�-e>�m���a�Z^O7�K,�J�7-�m�7]Lp��d;�}5A5���ֵ��A�!Ή�,�"ARt��Bb}��!�"7��oAW$����{پ�s+�Ⱦp���Cx�����w4���˳�����QVP��j�mԮ��ڵכ.{������Gh������T㐇�T0��gt2�wI���G��k��}9}�+.�dMDF�a#z�<5"�[y�/�{yO��{��6��u�ԝ`5�"�8j�T�$��D�#�fΥ��&ugѷUh]�D-'Yi�sb@�fҞr5e�{tLm���[��o��XiE�OC
X�.�ݝx�U"���3�`�u+w�Z���n˪�KO-Mm�˘�1�{G)�[ҵ�^��s4G�ķ5h�/0P�;K񧓽��������Q���q�Я9"�,��,魛�"��P�-F4b4�
��[	eUg�m0�#z�N��c�R즠��q`VIf�L�8n��+t<���]�-_%�nŴ���F�u�5��n#��y�>C�詊���6"/Q����X&^�r"�꘷#��w��Xٻ{�8J�;|�Su��j�N��ٛ�Pu8t����wc�@W�`���c�=0���,�``��E���'����.�}Ո����ܧ��7��SX���'�wac��^��cU���Sز�rVP���.�@�򌛖:���V��;���ŝ��e��x�2��"��_S���D���gQy��En���ٛ*��͉�:�r�\Ɖ�g1\�0z�lweA���e�E���6{��o3l��g���-��a����l���L�0����z9��=��+��{�x���A�y������+.G[��]�d�=��}Y�^�f���S�qR���q�mo$�����e����ID�	ͻ$��pdcV��T�aΒtWY�r��W۩���.��FZ�j#�+gU�	W;3�{x�,W7&މc��&pE���E�m��S��3���N��	���SBaz�V�r1��Џp=DOenziR����U�/ӈOo�����E]�#�f���%��	^���]�s����Jt�M�2�"�<�}��y�ab�o)���
�7,��6�n���tM�5P�f'Y��7B�/�D<Z;�����zw٣j r��ً��	�@�vV�*���l�@p2��f�	EY����0'0K)Vω�R�=՗3�Δ�B��x�]��Uۄ8��Ue��k융dæ��
��>s���W��a��������ĺ���/��$�A���|q�{�_.V����v��R�G
6o����7c�Ky��Ҏ�y5��G\sgU��Ͻ��=��ʯ �jJ�]��z��N�p��J��Fb�>�}2�Q��k��*<��E9ءι�����W{Ռu��\s�V��uYhk��h�z����{R艽k�TS=��)c��s���<luuE��̙{�y��R���Y	���g
�����Y�� -w�+ůҺ�7K~��u!fN�5����� W�0zx�>r�D�ND�Ɍ�<1��;&���}0ъ*�r�k
�_��S��]�G���������l�.�Jέǿt�����RRz�);�<&���ftB�'�����x��f�6Ӵ�����BZ�w(��z&��MW�_�������`�wr��g���啾�qbΌ+S���˞�F,��_�U�Ded���>qe�^E�������- �}�{� 1��{G5��.B�&������܈��%�����=��g�5�*k	��Rf�v��힙�ټT�K�Q�.��wX�씐�Wzа\k6c�d�c8��s�#���)�z�o�/bߣJ�U�ChQ�uxŦy��;� �B�դ=|�a�jD�7��Y�M�ɪ�g,�-)~bl�a�	<j�YKWs�n��k�ES3L���x(R�1����i	E��3��⩦�;��A޴O��`���F�z����4�A�k��]�V��5h=�x{�ʕ�T���Aηʯ�(�.�'w���v,�ܕ�ח3Swj\����ZyC/�խ�yfRg����XU؅����{V��j�}��TN\0��H�J�{���n���R��^�hq��ju,5zm�Ўfs�%mʔt��4b�ቨ�E���da��r�P}��3������7�]���q�} ���`8�L��^���v��=���
�*��9�{3�jr�����Wm�}�֘��;x(��im�;��@Ods��z��h�齬�vs����S;���Ku��47�,.0�'��7b;�[C��==�-[k#'�"9L����qƊ�:';%O����c�j�<%ף�j�N��*���s��r�.a{�K�����W��PQ��R���X=��x������ҭe�M���a���=�E�8sm�M��x-�5����C,k�8CR�0ژ��ݒ�zWB#0�E�uɉRJL�8���ֆ�20E��IC�e�阦Ij%�|���n9�<��OC�:�zU㧘�'#���W����Ǐ�o��K�����Du�����2i����{��"���N@�rي�%e�M\�����29b9�S���vS���f�yNߋ��
�q�������=V�1P�y3��@�ϋ���3��N��㟜{�n�����Y��ѭp�52���k�D��d3NNf�Ոo��V�ŚC��c%`�k�n`�n��T�Gr���:o%HgŜ���ug�ʔ:%\�{��3�fui�[&����q�ė@m�9����M#.^iT՝$U�
�U3{O>����tOT|�ҸGo0�m�Qf�C��`�f1�t�V],��0!�
b۹Vfb��+��,��i�ó[}�-fM�n��1oV���Nr�l��BRuJ�T\�Ճ��ϮS����+�����,-	����ޭEd��T%��;�k1[�5!�/!�^�J*�i�m�ܙ)�L�,y�S���z%���Y��u�D+^yM�}`R�r�0%f�Ű+{t3�Rɂ����LLͽ!��C�J�b�V�MQ#y�7���[x��捯���nN��{�\�x� ���wa����Q�'[v���ш��Z�L��H��dY�΅tF��Jn�u��=
����$�3b�gY};W
�'D�WX�r�򛈑�y���U���sB�
#���=W2�R_s��_V"����G\�~����,�;Xt���=>�pُ�K�I�;�-�����["��}]E���=�׃�^��BU/&|J�	�����a+P�vl��]V+�%�XݬQt�\YX�w6h��Ս�'iNR{l��jpEh�ډ��Ym%ܯ�
���R8��ռ�۬�8uu�3g"q�]�/�Ib���]%Gb=K4�9���v��e%ɝ�5�Z�b�Bm)�=w����ٯ�0k,jme�493�Ř�@R�EhB���-{�/Vt�R�<~9���DdF�P@fn���#�@�&N��q�B�B䅨.� p��m��f�r�ov˖x�^s�g��:d�yZ-0Ec+B��(�Ҏ�b�Ղ;QQ����Ċ�[S�Lt�7.U2�Wsn���[�f�-RT�2ʪ�j5���s7(k(�h����m7�L�p˘,�1�[1�KX�[�qod7)Xp�ļۋ��	0l�X3lu�G]L��m��nn`��
��s.m8m6�Ԫ*�;����.��F�5��Զ��ڪ[EQ1+m[�vSRƫ,m��X���4�^P�0n�LS-�6�\b�m�bKe�V��PjU��h̥/.(�"񨢮^&�h��b5�"�QEUQ6�U��ED2�D�1��LNb�0v��EJ�(�TG��Z���[�jT`��т��.f�|w���:<Vc�8���l���p���p��!�wW���ql���ze��#tMۿn,�������ŭ/I4C~�ֳRMD�!Ό��n0��ػ�5nky>��ɌD. ��^�Ӻ��Q�f��xVGT(��z�R����l��j�J�L��k*�wm�Tִ�;���ܰ��ل�U�٢럷8�cXL(����?��^J~sM#�;"�[�m۞Z�x���N5��>}�鸉s�eug���ozE�����+��t>s;}�0�د�C佦vS)�yr!C��z����ŭ��X��,p�%8�.�{��/Pa�v�x�� �]���=��o�ܯ\j��f<{x���s ��y�{�$TM���ۑ����S�^ �6=^���|f�wM?�B��b���lK�R��^��+��B��ʳB�T\ǘ�]\�ܻ��#�ku<�-���f�E���j�
 E��G�Z]=[~��W]���ǐ)�9?F��M��#�zc9L��UW̘�H�f���a�C:��FV��Mp�.b�"snW�����Rls
�e���������c2��>��q�0Q����0-1 �\Dm��y���)�δ�\ﰁ�{[�{Dr��-���VQʨ�"�,jՂ+kڨ��t�ˇ�^-��i_[���U��DQ�ٕ���+�"��O:Υ�-�n�����S�:p[��#�.y�=����7����_1�6g�O_o.=�B�2�H�������Hg^�������*���u�M��y��3���%����so'�vz���mogQ��D�n8��8�8ٹ�;BN���Km픓��*�׼{Feu�0���-5���o��gep�&���m���)5Ȋ��ڏ�z��>�����ea��	Db�8�)���;
U��Tg�mw'��MY��/wb��J��0̄��kFp�s+X���$�o7nާH.��-ʳ[���])`:��b�٫�c�[.8�Hdbމ�ݰ`�tֳ9��5�n-ĉ�8K��CR&4M��s�7ɚ㎳�+�:B�>�ѵ�tZ�Ѵ:Du�--��J�*c�YB,�V�69� 5�Q?�}��Ec�5,�{�'�J��.�n��͹�����6�;�u/Xz�JޛϦ�����a�2�8�K�fT>�Ӹ�)��V�{�e�+޾�L2SV�w�@���6�QI� ���j-�g����5��X[�n�+�1Q��{�1��9r��5kY�h��ϐgf���I'f�p��!-�<���N��@4�ac��y�]��f6�c���6�t�Ł�|%aKtNJO'jSl=��Us�3V�.�ʥ�S]
�iS�7z.��S�;Y�{N�o���Vr�ҷ��$F��M�g�\�ʁ��W�%QB�%��yQ��o����W76���f�v℘s��\�I�����9r��M
�̜1\�q"0^�q��w9Q
�<ކ4Ϋ�X�r��Mq��J�5�u�-��NA�o&xf:T�d�YȤ�����k�����p�%HKv�较��:������買g��+��>U�g���MlT��;���*��ZV�h��uB-�-��<��#��A��uf���-��WN�jY�۱֍� ��m�6c�)zIk����C�Y|/}�a�T��̇�q�4�i_k �fᓀ�T:+3�d㦇hƗB����Pg(�[�(�k���T��ʫ*Są޾襯o<Y؎tM���Δ�;��#{	�T$YZ�{�+@[���
a��dA�~B�E��uI.��fr����n��=Vq}n��ش�t�B�.�dz�y�Ю)^ռ"�x�fD����@nH������û��f^�qr����[�}��JL�/����b��|B�Ն��a.]E�1�k��V��WYT��i�x��;7��8�S���9ذ[Z�͸��
ب��:��$�ƢU!ˣ��l8}\���t�*J]-:�������8Ċ��f�p8��è�Ž�A�������̽��0�)n���kJǨ-W�so��f�5%��,��}���)5�ql��_&��x��Lv{��k4/��U��eR���Jx�g^�y�ލ���7��.����oy��?DSHYܴ�љKp��n�B�.^w������hU�/gn���kvC�Ε��O�������B�'E���3|h��t4�i`dgNe�#�E��Ť�Q�O�����f���F�;��7ˮa��J8�H�����nH��6��n�DH��8��'���[��"c�3��9=��\�������t+��b�\��2EFO�;���u�Oή�V�V����l�W��*La38��T��9��7V���b�����P����2��y���Vsnq�g����2EgC�&�Sټ��̲֖�� ���_�:� QC����Ƭ�߫˂[p���I[{[`��c��<,x�q.�&�HX�YI�cӲٝsq�Oy+
]�T)�WKZ�J��7��o,�F���U�}�5�ݗ�����}+Vs�_���N��5��Ѷ��KQ��z���.Y6,�{�Dx�V;a���'�L{}�NrD�%�^��[gD�dбP��~W�帄�ݣ��-<ЮGD��A좳bGT��^�OT�H��	
Mz�s��s���^��s	ڗ���ul�R���n�E���5���wO`�z0��՛|z��rjGt��O���-�[�霭��s�y��ȸ.� �cK����%n;�rOsn,�I}�#4�ę�m�us=0ﴮF���A�j���3��$ª�Ȃ����c�<v*a%�A&#�nF�Gj��n��.�'������w:�i�,D?��J�a�S�6w:������v�k�����Rd���8�IcJ�Z�`���E�	nF��R
�X\�}�Ĕ	�%��7���*�~Z�uՋ�*W!���D��ff&�Yd��:f�MM[�f:���[�yL��㰧���w9.Z����BPl�w#}.�gŚ��Xo�D[�5�_S�[:�MeZgk1�w�.�;�U�(#���֢H}5��	�]|��e���H�ǃ_N��հ��r)�_tb��>fi�ӆfL'���5_����h8��Z���^Q@���<�gsέEtʖ����]^'��=AǴ�(RRI$�O�TD
���*"��QԢ� LمOHIwȡF4�F��HV��nx�a�l�������MIDIw��"x��8[eQ�Y��*�tJ��A�Lh���8j����LÃ\\�>�����*qX�
9`����E�<��՜�;,T3�Y�ظc�ED@���y�V�t��� �����0�p@Q�(ȔZ���a�8�8��_�p{��������u}Ne���$	C��ED@���>�z;#$�5�2�[���sB���n�Y&���`����)N���w���2�0�W��/J� �?+�QQ&�Ms�6ׅ7�R�&*"_	P��CS-$�eq�R��Lbҵ�zX�8M3�gz����p��K�M�4|���`>����f���7��?��Y��҆�A(���h�*��ڛ/֟����j�0���m�Ү��q��N}\��v�d�M�`>/c� ��]�_˳�����B*"ר������,�d�ʤ��J��z�;AD2�r���� a�����%}G�����bX(	�a�.Z����k$�`�F�I��>�C�b�� B-��H/�\,8{u׭%�IHQ!�1��*��C�#X��jĵ�2�P> �"�����;��8���3���^�q��|4�3^�@>F��m��*	˳�i��:a��u�N}�vr'�=��rW��C���Q:n�n7��2x�(Q^^�xd��"� Q},�fMO��=[�?���ZmM�����i{&$n-R���BV����A�����PZ���G���'���eSV��[gk��*"gQİj�x�I]����dC��������Cq(c�zpȰ`-�,/na�	 D���7 �o����ǫ` (��<�ܐ.ip��ݵ�v���5�W�kb鰄��>E��Ds����w$S�	m��