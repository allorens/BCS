BZh91AY&SY�\l ��ߔpy����߰����  `^?}�     �      �X �ǧZP�����/����U}��ԛ��9���ã�݀0p@��Jb�)Um�!��:S6B�b�\`�\ �J]�t�6�Un����ܕfY�������NX��WF6�TΚ�bCYP�:� ����%-<���gk%Z`�� � �kl�QUPHQl���ɞ���&��L �  �OЉ
J� d4 ��4h��IE2G�dڛP ��2�2i�4�M$�%UM04 &� 4��M0")M ��d�j6�SD�!�M2��MR�6��?)�~���Pa1 d '����S+2/�,筳ng�?tT0�
�D>��W�/���~��%T�RX�*����������鼍rx.��G폱l�)Ln�o9� ��2��JRJ��*(0;I�$!�$2
����?}R�(+ȇ���`|����_���_3��g<���ϭ�ϮG9�s�
*B�b��/ўg����v;��Ly�ʊ,�LyH�Kb�SZÐQ
-N��TR�i
��V6�#�5��6����K���$��p�5�^y��u��9��6�����b��pZаx����u�pr�q�W��؊b<�Ss�����s��9��s��9�?��5^_�w�\q�X�!=!=!= ��x)���A.��&>��:�k�2�u�C�;��������rf+��>��SO�5�}�G������M�Se&��J��Hv�8SN��5�s�o5��hW���|8������kb~B�B�L��~Y��bՈ���	�88>��C�Һ$�<������f�E셲����c}�[K���t;�ǣ]x<�z��!��X�"�:ν�q���U��t�X;t�.D��h�6Gu�q��zy�N1�]z�/�գ��Q����h�N�K5��R�1b�b5���R�-UDs�@�h�+l�db)�m��#Y��1K�@��,�ȴ��6���_P�G������b�����@宍�8���hE1t�[��ֱV�-++WD���G��7�pi�������b�7hD~B�chZ6�G��C���|�5�5���E�Q&#ʺ�jբ�G�+0��Ӛ�5�����b�mb�6ţoʆ�SG#��N�p2S���F�G�4Y��-�ɔ�)�.E9\�g�����.J�^}��Ko�lZ�=�'2���J�W��x$�1���n8��|�4�p��\5���!�!�&�I��c�C$������S��7��0wd�[�[���666;��ǒJ���Ho����0z�h��?so<��g=��^vrp�L��ŋ���qtKɊ!1t^�;z�U���+^8pGX��Sթ�)y:B{M�RJO�R*�6(��Bm���ꔢ"�	;;B�b�1yP�cb�q���#�G���Ӛ���i���{�d��V��??�)�س�6����?��W��bw��Y+a���5�s�e!�*{s1I���kw�W\�$�[LۚLZ|"*y��r��٩�~Nl�<��;s�{ݺ�v裃�B��z���v�U#�3]^�7:��'�I�KiU�$�'�b�mwu\&�!�nih����y
��s�S(��I���㟝�~-d^��������"�@$Wza~�~�c+C�Lߧ�w+���v{�'�e���{���'C�l;�;�}��u�N�q��bٻ.�GpBc�j�d3h5�t���ȡ��]�&��K$�哻sk�[�Щ��o����ɛL͛�ɕccq���h�n�I��n��:�{���K]�,��{ޞ���+~�"nN�,O�j�M��ϲ]¹�+GɬO��۫�~O>�.���*t�o�WI��mL�<���̸[�oL����˘��Nd2��j����~m�`p]~.�!o��p��8���{��ty��`�v�X��M�^^�z�]7���t�x���r�f�ݽI �IwSGO�ɺy�,ɋ��0�\5\sM.�����h�2�	�My`�`5m�m�J�^�pfn{$���{�׽��u��ٴo������܅S��7L��ҩ����{<��wz��]a����0�#o��qfe�m������b�cN{�O;����-��ݺ��U͒�3S�hj��MZ�\d�e/`�9e�r�;��雉�eQ���fr^���i�ޗW`��$��L͐�Y����۳N����)��ץ��&��01wj���;;v�޼�����5�g���;#}ܿ��%��t�jw��N�IN�7V�ɢ<��sn5���V�f�&�&�ޖӣ����`��,5n��n���q�PɋZ729�(�'ݗ�C����ʞt�}Z��^\Oɸ�kX�Bf�X�M��Fg`���ͥ�fG�	�,���f�֕fI;�,Ly6�UC��g+��J�
�5 �964Da��2m/004�ӢY֪�s��h�5:�L�[��Q����مɛ��*��M�=���,��}�b�x�Ͳ2h�2p6��v\8�H��2��E��U�_����~K�	F�i����pHk�@�S�;�a9�����]t�t�:Z���hȶSXL �̳b���� �ƨ񲱃hm��T2
Z�qz���<u���1��G"�^�#&)���1N'-���n�Ԫq�:8)%jr2�KG/���U�,-P/,nDw9Vf6Q�tn��Jr�㭉X)��#�hg	#pLj
7#��F;LU�AX���n�N�b0UƜ;��Iq�S �nZ
�`��*P��� �i�N"��T�(����a��#%��t��T��(C,��T>be�
���Hې��rW"%WeO���H���фY�v[-M9YK j��d�-(�B+�=}3f��י�����ƛ��b�l�Q����6D�Q�̰U�2��4�=w@��ά`�rEY�Aw�D�`��C�g�]H���TO��}�����<��N�D��(�� э-��T��r{�-��:Y��XVv����{OS��FP     �`  $��.�N_}��]�����o�� l ``@�@ 0v@۽����Z]�Q��Y,r�O�N�Ĩ;w�  � �XX� ��`y�M8���i 5T��Y *H#}�q���h ��  �. X{���{ͧrv�!C��P(0jD�q�R�\i�9T�x �
 �t  �PUU@�Kɂ2"D�Ȳ�"1Zc&��� x� `@ F ��zU@�jq[K����Q>q7M�u��Ƹ�k� ���      � ;ޔ�-$�bLV��	�&`�	Lʀ�Ҍ��4  @       ��Dk���q�s���M�. L����n�����~`�Y�؊[E�?��������>��O��������~O�����^\{x{q�Ƿ�{DЄ�BB���(�/!�P�4$+M��u
�P�H]Q
�2`ɓN:Q���"s�g��R�uj��V'#�b"��X셵�آ�v7U�H�,��B��t��%u���,���ɯ9�v1M*���8��C|�G��ɍJ�m�(�	 �k�̘���UJ
�r[�x�-���Z'�d�VؚyŊ�V���*;H(ۢ��*���vچ�Ȃ
���,((�jn�E*��;���#x�3339�ĳ3338��fo{��C{����7��{��C{�����{����4p�,�Y���~2�	���`]��P���	�����ԫ$(C�'t�԰���ʹ�H�	�>���>��`ЙK:2jr8��Ч�*j�vS�p�6Y�{Jrۃ�~8h���eZ8pD˷�3UUP�o,����iOS$,�M`�o6c���-��et���[sX$g����N�6<l5�lJ-�0Y,��Y��L���a�s��TF;vڭ�����DN8	g�4u0�;�\<5���醄y�W*�����ƍɠ*��V�n���^H<nDn�"��ZGln
�T�CQ-�K�\5�oSȚ3O��!�t�2��˧�%�jI�Jj�U��F	�ц���������e�A�Yf
p�0�͔GRy$h�OM��q8t�8Y�A��f�8h�m�rd��u��L�(Ǳ�Xd��d�F��������E�9�IX�OMC^&�i�L��Øs�Ķ�&�����9Wn��l٫pu퍦��L�ʐ��ηg����9g��q�����w>�=7�]rEi�D������d���i��㱕J�U��r���S�"�nq�E�5;��4vn4燼�{OGĳ)��;q*���ʅ��Rl�xa�M���]�֔��z	��76x��=��i-x�2�gP}�>ǧ}�-[ӷ��w<'���Ǥ��ϋ�����~0�����p�0�x�NIҝ9):.�N���Ν9�ӧn�O�:yxv���Ӊ�ӷ��;>=�h즏�����B|:���뱽���{8rc�x>�$��6��>���[ ��jVL�g?���7����(kZ��8����i$!qn��iĖ�����kZΠ�Zֳ��!�ѣE2A
2�a��zE=Hd��&�i�c�)m��WN�R�5r�9�;{�%�5�����H��[<L�<Rw�Z���ݞ]�����NVE.V-��U-��A9`q���մ䲚�����aL��<pm�8l�t�FL�Nˣ+8�߶c5Pa\����	 �̸�4�lD���naF��j)�Ӷ�*�-�^�Zȥ�D��Q����OC��i�0Ƽ�M�0D��ɳ���H��=WP��Cz~G�R�ц�Z㶷'OO.<:y�y��o��s�2�����:h&���y�c�J�	-Em�
ND>U��r$��4���٠���ޯu��5gP�Hl�2΁��s�P����Z[�8l�FL�z�sʄ�/��L&�<cN�Pi�r�mpy;��.�b��.��xD4���/l�zX{��Ӹ�H�X�"e�zzs?g��b}:}8��
�x��k)><��U��c���4�lm��H�tR]�fξ��%/�^�N��-�J2�	$2�P�����M!EW��^~j?	�'��K�[q��,A%���0�j�:;Z�ʚ�-rZ�XR̲�O���GB�Y�S@i��Y�Q�My�Ha�[��Lׇ������
b/���}MkX*C���>Q�c;�N��.<>w�z7����yݱ��8��S/9_7�:rE�҇� ���*�y.��׶�pm�ɚ}M�'�p��J�,!�&�2d[c��X|raɆ8���N�3�¥@�xe�֓z_9o�V��(4���!d!f��d�4�Fmb���%Ua#�<`u�InR/�C��H%:H$z��: l˒�	~�m�����v;>)��c}</g����C��j�U�����S�lS�?|<8^9�Ç�pxz]/E91�Q��p�xzf��h�z.����M��|xgg��~���=)~8d4����"��(��Ij���x
!D��Yj��������,���[��%��d�֢L����N�-u�sX����@�H9���z��݀I
.:[a@,۶KQ�p��
3b��|s	ki�[ʥE+�U4
5 �
V5]��8�ʙ���b�m����|w+���V��-��&Уj��B�HՕG��k2Un���2�ƚ�qE�>>:��y�,�q�D�L_�I��y�����Ż���n���KwwwR���Ԗ���n����4-Mj�/=Q6�2���Zo���P,V����Cbv����X�˳b��cd$+6eل4G�!�����;!N&ݖ���P`�P�1xe(K,����3�U�������4'�Xhᠢ͔d�&7��e4P�����K)�S��I�,Ka���� Q:���X��'�E�G#!��`Y�Y�OQ>4���S�=!�̖�dh�P��!,��~km�R�p�M��MZ�T�G�["��%Z9k��나H��icƜ��H�U6��٠�'e0�C!�g�w¨�"����D3��<=ŉ�S�ֈ��,;�ƪ��聆�A�	g�4d�̯�����W|�Fp�<�u�2E�������&�m�ߙ.���M�@Z��+��Ǣ8�<Acq���a���E�Wt����'^���J7a�C''G&ܳ�y������>�=l��Ŧ[$�=8Qd�8)o�HJ\$l�Pd�;͡��
x�t����v^�5��l��0�\�T�Q�O#0�}��L�m�G���<^	y<�{�
0�х�D�i�K�n6�ap�=�{��Z4�l:>��8p��,�d�3�����qr�\̶×O`�NV��IqxdM9L���CGY����+�a��n�����Z�\Qk�v�ioI	A��r��<��ګ:���Y���7 �F�uc�&���Θ:YF{�L�X���X�dqR�*-%C�0��֤�+���ps:$��#lzUEG����e�[��)����}6Z��l�$C��!����m rnD�M�}h�R��SR}��CÆ�P��h��M�zj��L&bw��dK 鎝���dザm��փ}!"�֌�d�/2a���({�Έ-'H����P����6n��-��?����z0�C�+��x84x)¢z)�?��Ə��~>=3c����
�*p�^8\Q8���N�����ϖ*�Z�OQ�������>���7���P��V��A�(��CQ�Og��"� .\<;W��>A����I��kZΦ����7ww�����������Zn��!0h��0�I���I>,}8Sp4�>/)dbTB�'�4��%?e���fLUw:;,4�&��� ;<`�O_\���:P��I�h4l���#(�����K#�����o�1jvn�$�D4�FȆLM6��)��T�|H���0��0`�nNM[mz�ƂҰ�ԥ%�����t�$x�R[�
�Pi��IMK��Mk.e�inS��h����0�%bQo��}i�)bD�2�^�^0c&)2D6��4ު�r�3)��ԝFCz'0!4
|tl��� e��5�4Bt�I�S*E$��˙f�2��%k�.�������;)6f�D���O2�9��_s2�e�9R�W2�b%�R�%Kfz���Z�s9��q�Q�Í
6��ART�8�������U`�3$���}L;Cq�O���8!�2W/x�.��_&��֓�/a��4���Ѣ8d��P�a�t� ۧ/��g|�U� �͗�J�ҭTEl�_�l��L�Sq�@я$�N}���oN<x�txxOO�ֶ:Ja"m���$$9�H��sÅ׺���A�&ia�� �^�㶽�9>�|�7�2�Ogw���P�5��Q��Ơ���c
+�I*V��R�%%v��-�*���*��6�L�����iҬ��9rm5��<'\+GM���[��\�Ó�#���=�f`���7�U(�����o�a� �O�rxC���)t��4�(����u��)֊L�)v����_#P��'	�-%�7�#�K��%0Zd�0�Inؖ,�NeB�<"�5�%��)5��Q��LULe:�{	$��Xm�$������{���P9x���FBPƋ!���G	붊N�0�e���Ģ�X�Q�����;m<�0M�X̖C�th��	��?�����
x?�WE8R�xj��5��(��bz<4y�����ӳ�ӧ�on�}9��Δ��ӏ��a�~���������^�˨�b��#����jw�-o�mL�J(:5`�@pe��*V�!q�	�(�[���'T�0i��ډ!'�!�����AF)��Q��TPc]�1e�%#{$�Ox�^U/%�d�*���撉1�Xº(�$����<�6��VEvIi�Be	���i���9��k��)����2T	ԝ�vG-��#*��Vړ�hR)��ӑH��UEJ�%c�6��B��:��u���8~�>��w��׻�V���������ݻ�wwwwwn��݈KV�j�%�=H�Wx6� !�TD��)K
��>F����CU0jb�q�ک�L����I�8!p��1�z�у<��ٗ����,�=�5+�e�^1e7	2�<+E;L)0߰��a�d6`�B�q��!$%<7�̽���S��)i��["=2���I)�0�=�N�7(�����m�O �JM-�
4a4�0$!�̆�H&M���I��[�Eї���\�=�Z#Ncs130yKh2�gS���Լ�O-��(�G�6���p��8W�Ɂ<}�&�q�����+��Ys(u=5�a�jn}������η���<8���ӱ�I����,q�w�ϖ��[��Reb'��$��#Q�Wc:5E/
��:����ՂaQ1@���UC���*���D��4�1�^��(�{43�a��o��߻�Un�u���d=)�Ӈ�a��=,�m�d�O�=8�6m,��3�0e�Y��j�s2ܹ�PX^��8��^����C�ʷ��N40C������<�{�V�J�
}�)рm<�+PxŦh�s��X�.��ܻ�7������`�pɤ����8h�O6�d�[�����v�!�	�>�{�}�C��M�(��)��F�u}:���6�xb��X������'��`[1��ޫ����Y�*���"���L�«!�\X�l�۶ßq�]|�E��ғO�:t��)��G�)��1g&�M}^���L��Ӣ�]�a�4Y���0�-xΤ&&|ˣ���i��xhL�t�U�����ЯC��g����nl��m�>��ۏ>ӧ�=/����|s������z_�pt<.�W�G�����K���ӎ��]:zv���K��<�/c��x)§����cѢ���Ηu�t�.���/Nz^�y|s�g��F{�|����߸�,���{�w�s{�u�n�������������������[��w�F�h�f������̟���ɓ�i��㶍s��x�B]5|J6�-��=cҝY�o-���$��rm��<!�FHuMz������߮�?WO�1���u�2FB�S��c��0aɄ���	6��;e36��0�x��������V�E�ϭ��=0�̲"������S�a��cR�2�JG��U�R�I��1�4�m˂�8t��KᯆSFR>�}0a��ܒ�f򔞱颼���nK�CFI�X�r����\Ƿ�����v��\xo�w�t���~I��V(�d��@�|-j���8l����0�0�n��{�֋ӏ6���W|�p���ɢ��2��RF�h���6�`Ɍ�����Yk(��t-�l�<,MKOagǪ���J*�����OCzxl<,�&��}rAۗ���T�-l~E��ã�l�JY�)��&�jvh��K��d������Ģ��y��Gbt�V�@�t��B�$�u�_e�Œ"K4
�).�h�t�+B���/�a��f�[[z%�gC{��I�)�o��\꫷=�r8;�`�k�R��%�l�o�!�B��F���J���.:Q�و:Rd�rQĄ��W��U5��9O!ț��z0�� �	��!˞W�ɑ8k�f�v�'ϲ�"[7�Ԧ���3�VZkZ����nxY���k�1#�N^`��M%��̜����O��RtkO��L̸^W3(���zP;��^zn�OuF�ĺ|�$�nN��������8<ys���_�}=>v�9�|ws|vq���x:4p�0j<x�x4h�xS�pxp�<9��Gg�����S�����4r��K���3���.����ONz^^�y|s����/=��A��s@����Q��Z�M�ZF�n���O��9���KB&���v�Rq �HYl"��db��:X!����ڭ<�؛tG����r���(H��h��D؂+aEG*�#��+�	���M)#(�+{���T[����t�B�ѸF6�8����i��2:"*!�^��vÕ@�8�M��$�Q7+_!��l[�j���wv������ݻ�����wwwwwwwwwu-Z��V������Ae�m8�j1Ic��VU�&���`*c#L:D߄��ͥ&Ӛ�SDtO!N����z͸橧3٭
�8gX��<�;����N�5��oi��wN�͛Sd�G�Ů�us���N��M�'M92YN	ƀ�4�Zd�f�gʮ\��S�������NpA|o�4�p���F�8CG���K=Ϗ]���	���(tzu=�yKmr}>�#<��C�Bxl�o���_�K�Q6���ْ:`�Uq�lR��0�˗"�%R�dP$R�fxk�m��C�h�t���o�}媧+�T�<Li��眇��1.�r��xM��24h��N��P~9�d��q�6��ĉ���_'*�@�c�\��w�﬷��w;>�������F8B�7��{;��`��pg��ه��w>H)���>��5c\�lB�|ꉹd�FJ�
*()�F�mV�l�����ˊ�LfIb�����K�U����9,��ख:3��V��OC���S+՝.f�����=�4S�R��﯉�(켄���9EB(i�R���!Y�����L��\�*8�؍�\b���p1� ���=��G���:�x�ٲ�\k6�M���`w�5�U��Nd5a����5��p��4|�*��J�q��+��PB�-��(�X�1�b��F�(���$U!�)T��R��5J=I<)ʞJ��jc�9m:�i�:Wi棓����SG�s��!�7uu��r�J����s�l:l���|����tB;�Ĥ֟	h�uѾ��ۗ��Tn�ܙ7�˞Ra�ih��÷E�'����K���/��>=9�|wq��g��g1����r�<v"p��t�K�K�Nt��ۥ�ӧo)��΅8T�xp�p�9W�4p�8%��x'���ǥ�{=)���>��@y�#UC>.֣$�H'��2(��"/�E�%@d9&2�W{�Ϸwww��������wwwwwwwwu�kZֵ�h4h�F����H`|��>��x�I��dj�3���^k�����]j�҈�A=ڮCZ�h�S�3�[OS�mlɲ�����y^��U�.O!������%��2�n[��>���@�`K+�^���s�xմ�SG��͆=)���j�~���­�F��KKl�WJ�*�i�U���G
h�����N�I�:z-�R:6�Ρ�K���,=!�'OL�
<2d�k�׼y�N�у��s<뒋�e-�ÎUUb�99Z���ϳ�C&Il����Bm��~Ơ��$��OSP�h��|<!����$�#��&���̔d���gtH�<3��y��&M�J�!S��13��㶈��S�S&�%�(������M����ʹ�`�n8$���SS�O����
�Rz���'�4�}O��9�q|�/��_��^;;�9�Ə.�w;�\�V�6�R&�+K{ �<�ۈ�]c� �>=�f�)(���y2�9��m{�^�}�o���~�`�(�k�q�B�;���
,�F��7o[�OY$�)����"y��'�o�實�}�v[��Ҏ	���<M6h�xp�GL�vo�M�6y$6�s�d4���0B�R�048lG9������3���I��R<ē�r�$,6d���'3�2�#޸5�s3��.�+.���o���q���f��P��s.�L��K���x>����_�)�.���GÇ/"�18Tx<t��Ӯ]9�ӧn�N�]�<��t])������u�m�tp����ɢd�G����F�OK��Z6V=�3w�X���z�s�dɂ�ΗB��EV'�uf'�	����YQ�E�6���#�T�k1�X��ȣA$��GG����78́<�u�V��-��2;(�RD�|(�&ԭG�RX*�M�F�Z�C���^;�`�����G�4{g�>��cG�-�_$ry+����QEF�N��d�ev�(��������hc��UP�U5D�e$cm�G�fb�c�����x����]��������������������������Ե-Z�5��K���il�R�23�J^
��mت 7#pa%M�_%����+8Ԉ|G��q����=Zlÿ��M�y�7����C}򲭺0�C�����v;<(ɓ}�&}R�m2�I���M9<$s��gsӸ?N�k��9��\I�2�����3']�-Z���
xzSgCЋ�G�!�������+�oW=�}�KSSɜLB�6��2�}��=�	4TMS�$��0Q�$��Dl�s�g�R�U�tD���sS��u�!i��ʄ�=l�m�	N�N�xeg�]�Et$�①�2$�䨙w��@ ��+V�(P�;�bl쪾O����S��Fک��<lȝL6��9ʓP�S�__ON�͔��M=���0��?+����uƾ��ju���S���-��Z.lLw�Ǐ�yWTS$���<(ђ���bQ�㷏��y��.�IQ�������P�T���[,ӂȸ�Yω�5��b]�i�=)�Φ��#dzø"q6�`�F����`�i��(��T�GG'����zx���2�,Ι�h��E���+w�l��poڜ�L�Ye����a"�y�2Ŋ&�l����#*��F*��b�� qM�qu���Hi�����OG\N&����n��=oZƷ:�fZl��p���	��Jh�r���0�y�}h�Î����M��_1�^j�WU�k/�5���κu��N�^^�N�On���ޞ�]<:qӎ�{q�����������Ǵ!�B�Zk�HHBhB���;=����g���<:yt���Ͽr��2w1f����;��������������������������Bժ*�pݺr�ɇ�y�(�����vM�=�8�������}�q�l�d2l����*�*p�3�{�y96x]�g���t>�E������:wO.�ʼ��'o�ŷ�b���8�ԱE)"���J��(�NV��+SXi�&��QuiDjC'�ϡ�:�n	�vF|2���f��ۢ��!ӥ�0�e#�3�&H�|M��^Lr	��M��1+J�`*���>A�x�0�z��Zu;�s� ���֋K��3ᅞ�]V���:F�4p���K�y�owwa.�I8=�̯�,��ᤑ	�\�g�{��d�f��>յ��C�4���3.��fB�&�CM�F:INS���������Of�|�t��z���f�%N�Tr�5��Gd�K�D�w�S�c�9��{��{Բ���lޞNvj���[���|��Hd�̖`��/N�6s�Z�7i��&OK�]T�/�:�p[��O2Y�f�h�f]�Lz�S�̞��M)��!��];}m�L�Kr�er�<|6p��ɓd2h��!!���=������Z:�wxnnh�p��o��$�����Ii�	�~'I�_� ���)F�E*�ƃq���/�����>����	o�|�fvv[���m��@��ow���-)��j�3�BD$�E$�Ô���A�ZdY"dL�E��s�-�DD�EE�sD�4Y�"h�!��nh�Z&�"��!�#s"h�!E��#D��o��6�4[Dȍ"dL��b&�DD��Y�dE��YȴDZ&����4Z!���E������7D"h�M�ߜ}<;8����H�dX,�&�`�"dB&DȲ;F��"Ț-��B-���2!E�-�mD�h�ۆ��h��h�-�k96�E�h�-�E�h�n�vК-E�h�-��rm�E�h�&�E�h��ѻ�B-�E��m��n2#D"�"b-�[D#��dX��L�f�E�L�h��,�Ԓ��#s#Dȱ"�[D"�&Dȶ�h�"ȳE��"���"�&E��&E�Y�2,�4Ȅ[E�E�,�E�F�m�,E���0�F2��# �1��i	�%���BZBL�$&�$�d��&��BY9��m	d�Y��0F"�c$�*���P�Hdb1�F#QPY-&��KKE��� � %A��� �`��kCZd��L�d�$�u���	$b#H#
Ā��2	�E$kk9nJ���#[F�hF�Ѥj!�e0E� �dY"�,��9E��,�"ȍ�ی�v��D""Ȳ,��ME�YfS:���Ҹ���'ëO�Bi�;����X(*0��F(������WГ����\���������'�?�?���΃�4��?�A������3$!	���~������
2��y��8)��6����<���������2�7n|;�wK>��R�I?���jd>���;�����|�P��~_�������������h���>�LEC���$D�4�C������p}/�C�:��6}�m�	������o���������4�����
~�Њ�����g����� h�P��B�ר.����p1"������"RRZm�g����Z��4n�'ޟ%3_A���S�a��~.�O�Q#�E$EE*�M˰a��30�3�`�p�m���õ���٤6�6�ܶ3�魘������Z�@�zӸ%XSa����ɀk#���ۿ[�n��ۡ�yCf�1���D�l��7����"Y��$c]���L�~��#�����L��5��~G�RG�<����Mm��ټ����������a�����ұ[~�� �
O��3M����ٶ���9��?/�~�zG��{x:�ݛ�J����o���@|��O�L��	��,��_q>~�����9�����>~��;���~(�(|}H~�T��i?��!���W���������� ��y&��~��f�P�r|�@P�����"�pC�h��e�O����
���4�}	4��"��E.Q���2$I.����}��3��V�ᑣ�;g��?�y���G��;�f�)bZR/�E�(p��41 ��������[�	3�8�A
P�?]�RI'��?���O��W_j(
�/��W�� @�>����N,O�[����ٟ�ۡ���?�v��7cg��y��A?@�C����ǣ�~�?4�����C�����|��0 ��ɤ�} ��� ����"���~܇�sg����G��m�O�>���}��c}���W�}�R�R'p"D??��L4$A�*��4Z������L$_���Ϣ�B{�a�~^dK?'��o�#n�����������ï�? ����2rϲ}/���M�`=�c��~��6�=�Ăt	
w� ���<+�������/���>�	DZ)����@��y`���?������<~���
PD�0��.���6R?i��� ������F�((F�|~7������H�
3k��