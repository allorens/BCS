BZh91AY&SY̷���<߀`q����� ����bF��                w�T���*�)R�� ����TU$��TH�U ��JP�I(WfIT�()U$J
�"�IT�T�TLƁB��
R��R*�
�Y)m@T�% �T�J�"���$�D���JI%T����:R QR4����!*_<��()An`�P�l�	�V���j��wT	T*,jER�AX�*UB��%R�*�B��*��(�ua����� t[)CA=�w_=��Wf���5t�wT�Եus�����t��#wi��j�AV��SK��5�S�u�v�[������6�u���w��
"Rֵl�*k"����V�w��}�P��R(���;}��YH�R�+��MR�D�ij�AB�o['*B��8�ޞ�TS��{�<�IUU�^r�{����N�=�ρ���T����Ԃe�� ����*R��s;��U/Z�u���Wl�J�5�y=�l�%M�}=	U(��s���}R�T����}�(P/M+|w�jW��j�S�w��}R��_CW73�^}�R(�M���򪪥*\�*)"�t ���ԡJ��\��D�*��x�UU\�>|�zҖ�*��y�IR��V^^��F�T����UU
��{��IT�mjϏ���(*UU�}������Uot��T�+�S�H���FVf��T���RT� ;�u�*��ַ�����H����^T���<��=J�GU��s��T��ڭ�}ވ��U�w��֔�[x��AUR�����T/mRKUT�h�R4`��$�)*��)JTQ�>�DP���q�*�N��u������u;� �]�B�83 -�{�P�/(�ճY�w����[`*�r
��Pt`(��ҥJ����z4=iw �@���֋��n�( �n����@tt[I�v�@�bN�뭎 
�� P�	��H���O|��)@���^�A���r Sފ��h(�,v�7�)�X���pP*M�v�(\L�9v�Ȣ�UT�5�U J��4�|�Im�y>�PS>�p���hB(ӻ�;�WC��gRƁ�n�p�
�ݹ7P�:���t�%ER͊��^}{mS@=���5:w-j
�:�@�N���w�@�wJ����vv��t��oxV�(��WCG�       } 50��$hh �I��шE?M��SP      ��d�*�       �JUM)��d�d �)H���2`#hdш�� �Hz��*$L
zi�i��42M4��2~���?�k�?�����DG�������b푪��L����n; �1b��7� DB���PPU�TEO�(*�P� ��ǠH��������!�O�;����������U[���_�����t���C�A��������g�06<g��cq�c1�8�3��3���1��8�1��1��v�1�1��8�1��3���c8ǌ�3�c1ۏg�{`�1�c�q�c�<c�<`�q�c1�q�0c�1��3��<q�c8ό��0c8ώ<x�1��8�1��7�1�g�g1�`��g��8�0c�3��lg�q��q�c�1��q�`�q�`�q���3��>1��7�c<|x�<c�g�q��q��c8�3�8�1����3���3�c8�3�c8�g�1�g�q�g1�c�1�g�q�c�q�n��1��q�`�q��c=3���0c8�0c8���1�g�q�g�1�xg�1��1�g�1���zg�1�g�1��c�|c1�g�q�i�`�1��q�c�q���=1����c�4�3�c8�3��8��1�g�q�c�q�gc�1�c1�c�c��q���1�c1�g�q��x��l��1��1�1��8�1��8�3��><q�3����c8�0cq��xq��c�q�c��x�3��8�1��8��1��c�q�o�x�1�c��c8�0cݱ��=1����c��8�3��1��<q�c���1��0c��1��8�3�c8�3����8�3�c0c8��
L+����eaa�� 1�q�q�q�q���@���A�Q��Q���N�SG� 1�q�q�q�q�a\efWGG� 1�d\e�q�q�q��GWC&E���A� 1�q�q�q�x�������� �*�"�"�"����+�������U��@1���A�Q�@;ed\`ada\`��@��@1�aCG0&0�0.2.2�������������D.0�20.2�2�0�0.2�������0�WGGG �Q����GG���E���Q�P1�q������#�����(��*c"��������Q�E�Q��A�Q�za\dP�U��GGSfD�E����D�Q��Q� ��A�Q�A�q�q�q�q�q�q�1��GGGGGSOe^0.22�2�2�0�20Ɍ#���#� c� ���8�2�2�.0�G �E�Q��E��W�@�Q���q�q�q�q�q�q�q��q�q�q�eLed`GGS<`eN2�2.0�2�0�22.2�0.20��&0�2�L��c*�� �"� �+28�8¸�8¸�8�2�2�0�0.0��20�2.0.20.2�20'd�1�q�q��SWG�� 1�q�q�q�<e1�2��cȆ2�� c*�L
c"�0	�)��8���ˌɌ�8��1��8�1��8�1�c�L�3�c8�3�60c8�1��1��8ݱ�c2c�1��8�38��1�g�q���;c�z`�q�`�`�q��g1��q�blc�q�c�c��g�1�g�c1��1�g�q�g�1�c��q�`�1��q�n��1��g�q�c�1���8��Ɍ�10�8Ɍ�1���c8�0c�3��3�oc�c�q�g�g�1��3��8�1���8�1��3�c1�c8�64�1��8�3�c8�7Lc8�3��0c���q���q�`�1�cg�q�g�q�`�1�����1�g�1�`Ǐc�g�1�`�1��x�=3��2c8�3�1�c�3�c8�0c�m�c=1���3�c8�3��c�3��3��8�1�Lc��c8�1���3����1�g�c�q�c�q���q�`�q�lg���0c8�1�c<c�q�g�q�`�q�g`�1�c1�g�q�n��1�:g�1�g�0`�1�g�q�c�c�g��8�0c8�3��lc�q��1�`�q��x�L�Ɍ�8��3���c�m��0cv�A���o��~o�eOy��;�P���.u�N�L�ybC[L/iݛ�%�iׁʸ�Y!X,C�T�̬���:�v�͛�:�Q-��b�!F��x�ē),ۘ�nDs�o[w�I�*3Ԫc0�����V��T�aڻ��z�x���IлT��ѵWZ��C#�6*2^�qa�L��9m���%�[N݌(b����mkq�̵C�-S��P�2�l�5�gM��P�g!�shf�+B"�^T�+lش�@M�Z���0X�R��ӯe�'�ј�a�A�l��ԕ�ֵ��<�w�fXʇr���m��?�шòV77�"+�1�o!In���V��ʗ��k��]�GYR ��D?`��ط��i���eA�#���PM�G��՚�!��]U���SE9���+����52���EU�F��Bb�e�[�Fܭ���f�i\���e�zC���d�l���c���`�,�V���D�3[���C�$8�ʧ`�V��-�����YV�UU[O	OT��9�IJ^��۱ ��K6���I��*�>8p=;�Ub�һG �ob-���4�^(d�Ӥ��uv���Tf��n�-�w*#{��ʶ
.e�j�`{z,��u0^1�V\b�?�"��WYw$���-��m=���pm�t�	ki���ܽ�C5c��2�$���r���K��-��cz���A �@��fe�k%f �cj�����14K8.��I�c[pˋ3�(�ڌ�n n�tn($�yV�m]�r%Er̲��R�Ֆ�y�pJ*���Hq���:�**3Q��u��Ɏ�=b�Fb�Z��]����Fߑ��JS��Ҳ��J)��Pʆ���eF�PZ�Һ�(Q�X�V�)!�e��C�HUǚj���yn�U�jܠF[!]��[����J{V2�dKn��xD{M�Un�HK��죈ڙ���CYl����Nyw��*�R6r�mR$%��a��Y$ RkH=߬4�[�6@�+���(�U>r����	Vt`a��u�kMU��laK�UkB$�Ë숛�`�*��n�!W�(���J���S�,H���uH�vޢb.<&3�sv���9W �;5U���@�
���`�4��E��^V&��j���0�薘�u�t�&^��Q����Y��p+�W9W"�m�q�2*�/7G0\���D�
�r�j�;&�6���U�
�뗅iw��ۉ�w�[t+/1��!�x�̨
�k�(ٳ���s+2J԰c)!���ǰ�тA�w�w�Ʒ2f��EN쫼���VY�����c�q��3lø]�4 ��Q l�{�m(i�Ű�v����Ǖ3L��A�IoH���7���F�����F���7h�*C6��敮*Ä�7I�����v�d�[QR��V�m%�-��1�+pQ)���ٮ�y�r���(��-!Z�mJ2�f��LZ�A[�ا�2L@�Sf�-6��w�-�79�)�9m�w���Y��u�l$h��v$.�ïV��Z�R�٥SYz!M�y1b���Rj�T�Y��1%L+�)暇@�Fen]��Łl�%������ޛ�*���tVS�荠-�۳$:`X�n�,�f��*bШ��@;�0�Z�e27�z�o�[L8�@rfn�D�� �սlإ�lˊ�q�"�Y/,����i��;`���c�[��ݚ��KB�Uj	��+)���^:��{�fZIZ"���T�:�LX3,=�Ф�	]#W���)��7G)*�lm���Cq���)��r��N�J�`�-��i)�vP!R��aO8)&"ݖ�Ռ��;Vo
�:�y�6�60]��f��/[	�F��;�cV"x��ŚNGPx��է6ú��K���YcHU��2�q�NQӕ����*S6BvGt���V+i����uU�*˻,QM Qm�������q<n��hM�T&�e����vHu3Y��	������Yx1�M-dM�V����A5U�9�v��F�ҕ�ӑ���m#���XԙeI�,�`��0I�3Z1� ���D�67�6ޔ]Zf�n@��0!.���cxu���m�`�v�bXw.���P�&J��wP�kf'�t�x�<�(�2�WeTu�	�q8��]�p��B�eũ�z]$�ԎF*�%I�w�.�b,���f�Ɲtb:o^Un�;�2�Csiz�]��M�u�rV�Y���I��2d1�+N�sl�'r�Ǘr�Йc6,n8�R�1��C��Z�yE�WW�nZm��6*Gc+[�y&L�&�t�ګ�W%&/le�|�bѩZ,�j�&�аX��zj"اXb���P��+,i���JD��&�($�GYF�3;��Y�b�d�aݜ�ƻt����)K�t���=L�wnJ&<ݡ�[�o5aa��p�/���1=��j�rI���0*�V:��Kz�˫��p�M��ް��Ö��Nl�G��~z|�k)^�Q�%�$e[T����4F<��AiScq�f1�������&�õ�blԅҲ�P��NV��ik��!���vR�l��)M�p��ق�r�0rR��7O.$`Y����w2��+&í�����3e���J��V�3l�#9����W����'E�d�M͖��,9��*�K̍�7�+\%ݔ�����p�r{p����tl�Wf��MʹC��R��7l�R�|-!:��9D�d\�'���i���^�dC�n-��ɻY��f�|�Jߦ4pcN�1cs-�"Fu&��AgP�sNj�C^K(��4nf���Q�H�)z�X�-�q]�h��
.��˷3챴2���m�
�hV����[��'V	�c7q�&i"�1�Q�AB$Y+i������<Rk�!ĉ	��!H�ޫ7����S58�)eܳ]9&�p�
�L�!��n�I�[��i-�V���h]��Q��#4�Qi��j#W�V�+�l�Kc p�0��9F�L��h�.�<iaV����d9x�4^��%�"�mـ���2b�u��E@�׉Tx����liu�����G6������[�#$4wn���o(mU"����c[y�[b(4kA�	�3�%d˚/mٺ�V)V�tn�MǐK�3t)=Z�%�R�d�n
��kE��(���8.�E�#9�M�շ(-۵A���)n�B�����b�Ϸ���^�D�׻3G.�4ql����4��"5b�.�G"4�Y�����V�*	(,Љ���ޅ�L�:��P�
�BJó&����*�Z�s�Vn]dE�pmm|�S�L���nK[�\��-�U�+6B��W�BE��e�bL�V �f�m�1�ӕeZ8�R��+-U�%- ������L�6�{6�B�Fü�e���b���$�@�J��Fٷ&�kF��鱺�eC�',���q�AK�S&�0D7�n�G764�Z�����y�
�[i%O6 �n�(�Í��=����R�3z����ro� rgBѫD����X�Fܢ�rj^ʓ-�Ǵv��\�����%9XS-���6�ֱ�[b�8S5\�ucHN�!EGS]���d5�����n�RG��i��2|�\V�Xc]#�!���y���űt�U�&�Ѷ�������QCOk^�sh:��H� b��)�n໭̓���W�4�f]�����'2���D�/$;7J@�V�4��SxƳ��7�L����>�ȭ3�	6�c#0Z�Wb\Xl6^�{��f�$��q۴5bq2���ʬG$�
D�Q�-�,��8tSS]�dz�ZJ��䬒��U,t��䪼ShJu�9�r�"��L����w�����h��mBB�Q��3*�F���A�����6��yTD�1�E:v0�2�q��1̀�F��&��c�n�by�UZY��Ȧ��8��kr&�/JQ֨s��	Ϗ���ѧ��Z,�v�:�d���f4h�*¨Y��Ӕ��k�tT�.�Qa��E�B���71U:E$r�f<ۋ%�c"�ə���Y��b٧A[)>��,#���s(��K$��J�=ݱlKV���=RS��V.l*��z6F^l�3h�7��Wrf¬e5	x���m�i�%�(�	��{�c��ïF����d�@$�y���ث����阴�eÚ,��A�����S�v�Uj;B�n���e��:�Ы֤ax�X�f��̻ݡ��%\�k�E�3a���#����	LI�g���o!k�*B�v�3v��4�kr��=W�na��k��3J�<��b�&����sUL ��d�����[en���a؞ME �ښJ�iwj�]@a��[~���܀��2�oM�ؔ)�ȴ��(�e�m�5[g[���Ȉɬ��+{ Q�B��x���������Y� ��fT�����TX�0����i�-�z�
i%G1,r���J�c�d�Z�9�Ir�m"C*Ъ��%������HʺƚchM�Z����yKMi�J�jrE��Ol�!K+sr���`��C11�V
{ݳ%�{�oRï)n�m�n˳k"2�B��[m[J�b��5t�e4SXYQ��i��M�!a��$�Z���i�y	����M�ʕ��Vj�������� ���݌�n5,�����-E!�N`�]I7$F�3*��t,az��nּ����ܧ��.·�3NG�t��n]M����rB�#[;6��� �yi�T�R�8(ի�Ѵ�,ٖ���	���y+j�7&먞|#��
Y&K&����p��)`B���$���0jU�k%���z*����1M҅L�5r	Yy�M�5t��(�{�aI�Ŷ�F�B�ġ;��l,ش�,�/h;b0��3U�v*��N��c[�;Ǒ�W�Ր�Uɺ�Ke"R),î�(�MZVڿPYV��ݼ�wՁ�n
�e�A\�x�/4c��	�Z��,=�r��_h,��Tݠ��C�2$A�P��Ҹt�ƯhG	�]�wm��s1���u+��FUû���de�X�s"�hIl�ǚr�X/R2d�¬�e^8F
!V�P�׫7u�Gv� vj](�P{.hW�͈,�z���n�b����
6R2��iu�o6<��FсT#bn�/SD�l���N�&���(�l:�+ٱ��q]�b�tM�6)�Qd.�UZ�lм	�!z�ܽ5f�[���S�b�n^��MP��	�e����ycp��
r��
T��F�2<�mĄ���=:��N��H���|f��u�Uw��9��1u�98��H�i[�l-S/U�M-5dFZJ� jFi��Jǀ m��0Vcׇ3yf���\�Ε�"�]�?MR坧
o
܍�ڮF1OUb��Q���o4;̂���T�i�ai�%qU�U��JD�������2�.���򿠷�Lr�l��Zz���f+�`��%o��i�φv�,Z��{��}x��u��=���Lo+S��2]���&t�X��n��9��Ij���LT!���3�*�f�2���I|��Ov#t#Gfb\�;.f�L6�m��M����n��q��p��l����;kf܇i�i�qK�5��
sV���]Uo��2w`,�`�մ̐��"�r#�j�|����͊��yH�EEe����x�0�U�2'X\Ɩ�������c��F����V��;hC�Ai��Ț�t�P#�����a{tNo^�f��2�5 L�ZL�篳�&.2���}��hV�uuy��F�V�ii��DMwe�u��m���z� i*��J�]��t��Ku�vfLw;����E�0m���Dv�,�j4�ͧ|,��1TMqZ���<Gr
c�_$�;�!3Gj.P�T�3�R�on��I�}}ܖ;���e�-�`&20P/0���\[ɱN��}�÷L%O�=w�eE�<�*�1Q�6J�Ok�-��W*|��PZ�s/�>��pv�#V�����f��SF���hQ�j*)D��8�֎����Ja�X�+ʡL^^��z�(O0�ܡz�w&�X��\�FQc]8%��,Ҫ�=��"�h�.1I`�h�91)���l��P���O!�����2��̼,��t��2��$J�������D�����U;8p��#m �w5l�(y���/"�UO��~�I�g�%z]X�A,X����Pķ�b���+�0s(<|F���Zݵ�N�#e_�+^s���˲󯹥��;efu˺x��T���5ܘ�~���_.��,�H�y4�{�hku�0:�*�"\T����Y�3�K�����a�O��{�́]��Gy�4�/A���J�j��7YW⍙AK�jWݠ{���a��S/UV�|(��rP��o�ԭb�h��h�G5��aJ�[�λR��<��8Y��4�׽`��'\�1�'��
{��XW���w�}���&�U%v��0+��wz�'���Nк�X��+�����}a�	��&��#���Ѥ��ާV���[�2X���Mc�QTyh��z�;�wj��e�j����kv_t-S6��_o{�a�e���0e_m]s�������*�l�٦}��.�E���5��h��Ϊ|��g�A�~^I^~[��x4�X��ir�q�K��MiD���nZ$z��EYm�i+�i�Qb���́��YJ�>�4�%�����Gj�M ��am���b�;xd��}Z]o'˜�����PY�ñ5Uc�� L��9�Ukwvq��i5�؁�5�ݒ{{������7V�;ݼOA�Vޗjq�v��J-�}Yn�N�-!�%�8S��d@����AWH ń�{�o�v�T���J�p�5Z�¬T�TӚ�21�q�U��x�˒����g�R�d8�ҥ�F)]Co�U��L�jM��ff_t�8Υ��QK�JHăj�_)�r�c��P��jي�v�fYV&fBŒVa���i��D�KS��rsӲ_�!ݼ8��{[�g<ɬ�x�_*�"1�M�x�,hkD���:mR$ֶӴ>�83t��^G��0拓����O�~�w����2��W�y��ͣ�ɼ���4�4u�\��«���:ݹ�����xl�U/L'%9ք[�$��b��#�{�޴E����#�|�=7N�s�j��&�sv�EAoX���ʹw�^�$w9c�jd7�����H\.w�����ZC��xh"��%Q{�3��%���r�_;��1��
=}|��5p!�n�"�Y0�9vN�g������o=�n_Z@�k pg���툃�a�X��(�Cm�q�}������,Ŭ� �[�q�ȋy�݈Tx2!�T�������:v�T��SVH��R:�;���G>tWh9��g�Uj����ʜ�:�}���݂R-e_F�#D�lwv��˪%����Ժ&L�{���t�������}�;Q1ۻ�.����l�t�U��ܾz��2ͤ�A��rq=0���i_�s�Xw��w���(�}� \4j{��|�M�k�+��5��މ%�f�u˭)N_6���Ů��A��{���:�k�W��C�V��)�|�:���Ԙ�U�D������*O�w�U��j,md���j��]v���X��&<��,���doc�׉�j��&H9�X���I�wyE^��]��mel\��̧w� A�;:$��Ż4�	�{î[1J��q�%�� 9n����@ik�4��br;:���j��Zp|����!__vV��EĈh��gr�T��.�ɣ�栳�3�B���+^�/4�|��	;;�ȮJ�8��;ٺ�H!��b^�35�6���G-=�{��Ws���Czu�8���fd��@�>����*����ds���4x��[q�L�c�.�!����[���ߴ\�Kw�P���P���l�+7�̰e껛���:$ʓ8���:�|�ae9��P}�nP�A�>\�l�U�swGYx	ќ�`]G�;u�v�����.�dLC��v.�s�B�x'���l�l���14J���NR�C�]�k�\����7Q�""�g��&�ތ���P.���ug;��<�'�y�9���VF���v2Q����8	���̷w��@�S}2���s������k��#r��W׳� _�B�v���G%)u{t��mӺ�V˾I6y󑔭fS�\����
f�WܰJ]�c9��B[v:�v�r��pR\u�4���}w;0С�����s{3MP�3�J�D����Nq�^�Y|s��`J��h{�o_6�J�i%�2�޽�ִŖ�9/lm�w.�:*��w����ʎp�b��ۤ�d!G��c��{:�}ÄW������Pte�;�⶛��݅�M'rF��s���:�����/iV���p�����n�v�"`D����N�gn0o#U���;
�z�m�h)T��+P�ż�C�.��q�6��qTrh�JE}��O�
�]�B`�d������(�^�X'*�o�xom���d#��-��Ԏu��`3��f�z�b�&of@E�-s����&h�t�Q�t����{ݰ=U��f�eJ���˵@Õ,�`�ێiu�3eB�ܬ3�w{o!8�Z�|�����S���WZ9�������"�n��}^W�Y��9��b�I��w֜Oe��r�L���]kJ�c�G��8�+L�,+��cOVܽy����N�g�E�l-a�ksA{/�J�7h��Vwi�]���n��G3)�!���3r�S�\��fS�f�(�M��4��պ��sq������(:�lua�&���7mwp�w�-A{pt䷮��Rݎ�GL-��ƅ�5�uG�]�ր���/{I�C�e3Ab��3�(�k��M+Q܃^Xt��g1���W*6�Yc���.��w�k�2�K�8E��BvO�R�X�������Jxm<��<��<7Lc!K��fۙ���UcH`�z�# ��GS!�ɝ��,��ٻ}|^%��UZMY��Cۂ���:�0��#b�ofj����K"����G���S�`1iE�}�K��f����ه�m����"��3�j����N��Y#�l���w��s��ϩc�hpv���g��tg$
���1�d;]�U�x\�;r��'��rɰ��p�t��:ݣzꩍC��yX�m��P�ї���&�)�vpi%V��v��t�Q�r�L6�t�֒�������yw�4 �ҧݓ.vI�e�7�
���]�)kE&�z�u�*�ξ���fW�f�v�����w&NI��zwkA��ӵ��a%�on�-���'jVJ��L���)x�cȆ.HubX�dP;כPe��N�"8q���h�u�����,�����	��Q����]���9�\�@c�w7A�t�5mdݡ��1[��O:����O7`���ۆ�bЮH5Y�F���W�Ը�^F�|7k����ƚN*^�����˾2ߣj�t}�S#�Nk�F�]u��s;����1���LgJ���q�����fV��
]h�uֱ�M�5Jzr&���e��n�����be:D��bҖ����nn���� ��k�M��>�:�l��tس�R��ˈ�������@^[Z��u;��u3��vλ�)�ݼu�LvtWU�wx�x���[�w�d�9�slᷙ##>�� >G6�Y�m��<��
�_5��[�hT��ۻw���gF�䜣��z�*��$RQ�;��B��j ��e$�0(SS�����}�֡�3�䶭tG[m�������V;����=�Є�V��n�}�dۼw��-N�H��72㪳BUM������s�{�Θ�,*��?�<���Iլi�u͛��3{Ӌ��*��A��8kZ��s`[������gI���
�p����|��5:�t�|e\HB��mcN+��,���H����4jΠ0��W֨H�y2:��E����Q��}o=�_>"�Z��ďn�����[��r�b���bV u���2��,v>��EmEMWZsyܣvȦ�h9�b��Կ�6�I���r[R���길%D<tS'siU�4��!�'��gBUc�eݚ�]Y	4D��k���4دOH.U"��}H�>����;!�� �Q��6����VM�񩱍(�g�U(X8:r�nd���۸ц�l�����ۣ"��,Wp}|w���G5�b�wA��r֩�W¥wu�-m�B�w���]��A�@Ӗl4��Dt�CAWݚ,R P.^7�@Vɉۦz`�V(��a��$���]�s��u,�tF�vsx���Si��)f�}������*��
�co�q���ܹ}{t;S�������.�-��\)�.��mL�c�����o�z��
Po�:���ӭX#�U�[ɪ�	��$�y�T�U����k���9T�On^Ww�Su�ޞ�#x�-��8έ;%A|yIO��n���zEѲ)�4lԨoT(%�J�9��o���X��,S�j��(rp�OrU��|5-)vSC-�v�s�]sh'�/��ۺ�kf�xm���芜�8��JOhhyR1[k$�\���b��.��l��C�Չs�9%�!c^[��&�(�i���E;w�p��/�Ŏ	2����-I3�"��wo!Ůbg0�=r[��[e�}�Xe�Xo�b��L��PŲiW|3���4�i*u�܌mΩG�8s��B���H�|f���Ь}���7nu��-@����Qt�M{&�Du�+�@g�2}���͉~�Oy�,���q|�������x��O'.�Ǣ��'T�\��8�'����^�kBn�i�.S���rܸ�^��>i4��R��'D�=2�a��F�/1��i�7��m�I4n*DG̶8�
��ֆa��k��I>�PP|~��.�@iÎrm��v���ii��s5��v��J#G��ԤЧ��fZg\���m��Nf��-�7Ѷ�]��@�;:��Ԙc=Qذ�d��R�p��ݓ��w/��a�Cu6/��iT\M�w,ۻ�s��FK�V����V���9I�.ȷ
���XBய�VD���o�W\��z���{}��[��H
h�v�S�R��4��o%oXN�5p�4^�T��_KY[����9����ES�Y��4�<�Z�W�ʜ�v��X�#��]�t�C��($�p��F����B�ޫ���sk�t�t0�wd�8�)Ɗ9c��󇰐[MЭ���T��5�pm��}LYtM�]�$p��uiF�>Yn��p�X��TM�da���Y�>�Y�X��+�=HЕ��mn:���������.��;��Tp��s�Ct�dv�]k'��W�����w ��#7ų:��DAjT,��7�!˷Udbk:�h��+�ˢil�ŚzY��ip�z�'O�TNe7��p|�eiW�������UEOtJ[��xؾ�Į�mJ�8��{V�li7�mEAZ�
�zp���WT(&�M��mn� �s�w�R ���>g3���̹F���˲�4m�����4r)���:�Q��D�eoF"�tj\.���c^�O,�h��xg&ӻ&��|s��+Y�˷����;�Ө1�}1C�V��KWN��s%v����f���Qh��5fsc�Ĳ�v��ʽ
�Y|��&+�(F�z�(�#59��f��lJ�B��j��;c�N�^�I��}��=Q'���<�86^-Á�|�Q��D�q`̔��;UB�����C���	�)ٜ�Yò�7��Ξ*�;[է����� ��V��(������ᝫ��%eD�����"9�A=h&�֑ÁL��B��Y����Kn�}�$�N--�%擗���+x�J��r2�@��"\����`ŉӱܴ�%U�6��n=��_Qޗ�'�Ǟp��1E�[�)���c��+2*ݫ<�_7&Fi[�r�N�1Хx��`â��f�������in�_�;�����8ު�І�wj[RD9Lo �h;>[ف9uPk.U��z��l�c�j�`��g��/����_H��ݚ����'Q�&���0�|/�F��9;�%n>�7Fv�C��+GM��~YQRã��8,2��F�m��V��VE�+
=J��͗��Y�;T��Ӯ��YUȋ�[�B
�r�P�m	�T�6�6�g��Ew�2���J֥Ν�Mg5C2���許;��oF���B�Ы�3���+*�1�Y��� 8�����Gѧg.�A��.��UNf�S�"���x�}4[�K�<��|3�]��B�X/�/�l�"}Yuv�&H��'+2�;�FI�p��'HغD�ޢ�B�����|{�p-Vu�u�sT���y����*f�/�do%*�6�����'q�T�s�}�Ap>���{�B>�7�\�t���M�2�I3�ghl��f��ٔ���S�;4	�!�\w6����N���t�\�h�M���܄&�ɉ72XY��dCl�	�q�[x���3�Y'Ld5��/SuE��$��~�mĞꙙ��U�ۻzh�k�{�@�O�S	�,�T�L7^@�Q���O#�䋂����5

�&	
��S(|j�B�ۧ*AICNR~�0؛�Ww\��{YW��#�����b��Y,�u��/�D��p"s�Co<-'^4�[ƅm�\��>���]A{�}`��:��
h�t�/�Y4�TPH��i�Tʦۣ
����zI�z^Is9]�+�!��qK;��D���	VX�ԹT�����ʻ�p"g�T�%8-�b\-r[w�*�dQ�~J�L��N�UTB�A��ȫ�곖Q�3:�8ų8���i�2��j��]	T�UM��*]0�r��3,��T����P�UA4@AM�����ֹ{[`��@�a��,#,6[ræ����je�̠Ym9!4$\�]�`�Fțp�8IM���m7�5DUF�j��&Ӡ�%�À�4�4ʣk��[�Rb�5Q!jS�PO0� �)��W7S��OŦK?8P˕dUW7"96���{B��僢]�cG�E�y�$�6k�[��R�Ayud��R��&N�a���'u��;�*�K��*�ETD�تN�b��ӛՆ:�A F��	�h��1�e4&M"�J~I��H̷n����F�ٹ�p��B����,ՐZ�L$�tR-��^e
M_+��m�W��o5���83 �fmM��4��%IL'2ԉ-���	76��ȣ+��[BP��ť.�9u���D;�M�D�Qd�QA"�	�]S*�n��A�������Zt��
��n��^�R>���\�*�r��J��'>yt(�e��Ƒ	��r��E����ƺ�7��yf65�Z�h�PT)0HMʒ��%U
M�r��4�&��$<�=�9pc��W
�Xd�P!���b�$�0Sא$�R7YvMܧ5gJ��3���]Fόd5��/St̅%��fa��B��h3d#Y	),�A2!��$���S<ܬN��h�M����2�Y2$9l����/:.9Nx]+^?�'�;���������Q@����~��
��OUO{��߿�?@�`?�>���߱��k��K��6O�|��w�z��,ˢ����c�����%/U�hc��ӻ+5���Ak��kKgE`��!T\�I^�T�w$��od�w�n�+J�Ok�+w�m��b�]�n��eE�|Ew,����-�fi�`�s���xY��	_G)fٶi��U�s�5}��o*V�F�'��E�&�o1'�<�e\r(���؎N4�@Xu��W�qY\c����ɻ�s�(
Q�/���}���u�mpw�Zޖ���(:�.���T/yc�E|�����w�8l������W����O�*���y�������E��ů�SU\p��*Z��r���$'������6�����\�	׼�;��R"�lޝ�ڝ(69���lsݮ�}q��NF��3Dq��f^�֫׃Eۑfj[7UXU�I:�P�%d��=��vdd��rv�۠M���:$J�9�՛�w�d2[+�>�V��\�յ��Zr��=ϸLi��I�0!N�[��������=%�"R��9�aF &"����
��=xr��{��}�)":ɥ*\������]~:��]u�]u�]u���]u���]u׷]u�]|u�]{u�]u��]u��]u�^�u�]|u�]zu���Ƿ�_u�^�u�^�u�]u�]uק]u�]q�]u��]u�\u�]zu�]u�u�]u�]u���]u�]~:��]u�]|u�]{u�]u��]~�?_�������u�^�u�]z*::::&::&&��`X�v�CC��$uC�w���>B)nd�xW>���[i��q�$(;K-���,�<��͒*�z's.��#�ee�CP�͎U���)1ap����Lv�'�V��mR����F� �ue�<�;o	`���@f���iY'�puv��qؑ�n5U��ۘ���Wn�k;�L %����j��Uv�ܭ�S����Л$#�G��ѽ���R��z���!�n-�tA�3�,�`_<K�z74J[��-�x�	eC�7Rڜ������n�w��M��0d[vY�'zIf�e�aMr*8f����a�f�2�z����+��I�I��uh��C�<�N�O���w1e�{�5��Ə$�5�AGi��Rc�o�Y�ʂ�gs�K�y}�bݛ&�G�3��gp��P�'D�&9~����j��م]H��N2�D�S��+��E�FY��330�
�mdu'Js�X*�&@�*J�&�u��; 3q�gf��pP��15VU>;��!�1l��%T�2�̺�V�Z�}j�e���R�xJW�MR����X0�̦d�9[�v.&0F���F�GGG:�뮺뮺���u�]u�]~:��]u�]x뎺�Ӯ�u�\u�^�u�]u��]u��]u׷_�u�]u��]u�_u�^�u�]u��]u��]u׷]u�_u�]{u�]u��]x뮺뮿u��]u�]u��:뮺뮿u㮺뮺�׏�����~�]~:��]u�]u����q��A�э<쉵K�����Q�x]�:xĴ��hk��w\!wa�{�����Xlv�(V����;�w���73w�6,���3�4�sq%K�,��\���u��}���1x{�]r˺��+��ZQ"��+��*`ݺ�$g[{�L�DJz�TۇC�WNJķ����<:2hW�,q���w����N���Dx�dn�� �Hƨ�%X�j_2p��7*Ê^�}���^�b��}��&W&  )���#��9 nk[t���̡�L��� ZB��i9�㻳�2����b  uC�� 0@� Q��鰱2�e�t�A���qGp�A�x�Ҟe��\���4-�@��Eα��+A�I�;lq}�M$i�J4�KP�����-�F�D�����7q�a4,�ͭ��C�v�Z���������uAG����m�
�sd��1 �8�n�d��:��ҩ }���N1�ۅY��x<t(�܀���t�v��B��@̖3�"���2�z�aa��"�!��`wk&�s�1	�+�x�|H��-�XޢY���^�����D^��
L�3���a��i\|��y�raeGT������	 ݸ 	���$�
��6���6U V����םχz\�T%{
!���C��Pc&:�3P��^�'S�����3F���n/.X���h{�c�����d��.Q�"�	sw.C+X$�" ���wi�2GZ�Y`��v8��p���Jw]��D�KA��&��}꽤oP�t6u9�:����k���>B�������(X�/����u�]u�]~�:뮺뮺룮�뮺��Y�]u�]u��뮺뮺�u׎�:뮺���^:뮺������㮺�u׎�뮺��]x뮺뮺�u׎�뮺뎺�Ӯ�뮺㮺�뮺�뮺�:�κ뮺��G]u�]u�]tu�]u�]~?Y��~�_��뮿]g]u�]u�_����s�\�\7������mA�ú+��I���U)1�b}0���V�.�b�a1I�#5�p/���V^N��%v�a��wr/1^�ʹ�Z6ĥ��@L-b�n{�t�GB��ʴ��[]y\�����8�u���#,N�I��Z2Df��60!˰��ک�:/q��^��oWe�)��N�gh�F��q�-�6uwJ��}^�l�O@�� �GG�˕w��������4E�O����AT�pQ�����i��!��yY������;�sAژ�Y�˱>̖N�}�j>�>�|q��jO���#c/1�#�˂�� �5�}_}����[`�yR� �,a6���]�[�M�.v3٩���"̃�w�^>�Mƶ`��8J����LY� ���Q��RcL�B�T"
fW!=o��ƹI�V���Z�Q�LէW�P�	�d��o)n�Q��Y�Y�0�|�̽R�:����\���s��zOT��$�M6���P��z�׸>ׄD3)������)�Kn\GXyx�U�[��%�}W̓ǘ���#[���&��Aq�����K���,�����h�Ы�j�&ut�ݷK�9ulH�;�[DD["�)�n`iV作���蘸�q�Ѯ�뎺��]u�]u��뮺뮺�tu�]u�]u�G]u�]u�]tu�]u�]u��:뮺�=����뮺룮�뮺��Y�]u�]u��뮺뮺���u�]u�]~:��]u�]|u�]{u�׎�뮺����]u�]u�]u�]u�_����~�_��뮺�뮺뮺�����{��iAb����s�l��P�=cPa���LBI�- ��u��_U�BPS.�r�ӆ4�oRb�!]mP��=�6�����:ȴUY�!�����t�΋�G�Q�B�u_fG'Z�]bd�t�bȮ����f�������=�"��t��w2�f���o���q�
���U�.S<6��"�#p����.�6)b�E��4ʵ��1ۺ�7m��4]�2;ۆ¾xC���K�s&�9N����, ^�����+�Y�b���jo-#[�ۍ
����i<�����x�#�̦,����QlY������[�B��IG��0��0Uj�:�L���=Yb�����g�W/�Z;�e��Zݤ�&�]�8��*;�O�P63��.su�Z�4`�%���y-��w\���m!%���u@�<����+���M`�tK����0���(=tz�l�D5��.���Owkp�ZU�JW@�IWc�G���6=��8iAn��bfs3uP=AA�飇�d�*\�0B��됣|���J�|LԤ��Q����e�{<��־>8��Ƿ]u�_u�^�u�]u�]u㮺뮺�u�u�]u�]~��:뮺뮿]u�u�]u�_���뮽����ۮ���G]u�]u�]tu�]u�]u�G]u�]u�]tu�]u�]u��:뮺�:�N�:�n�뮾:�u�]u�㮺��]u�\~�_��������]g]u�]u��뮳۝�Ͼu�\tt���]ġ��2W��J*��f��7S�"X$�t�W��&d�/�_P̀�o;*�	SX�hm��F#���m��9Yֹ���C3 �:��T��e �:��љ�m��^"�51W:���7�h'靸�Y���y��v���.�ka�o�Ү���\Z7F��Z�,��]������K�
�d♬WU�-�����.�v6�[����������'ҫP�e�����TB�U�M���Z�.�Eʣ.r��(�:��zt�q문i���'r๐��dq�>��M�3L� 2�E�_s/֋B��.���wT�<����[���n����(0ξR��jo�X��r�]��i��u(�;+�E}}9������9Yq�ri�����<�68��{B�f�WIM:�}�t�'ئ-�1ɸk�zF��^��4��łQp�\Ww-��x��&²{��U�2sz��+'Q�TNl�V:��oe�"�uZ��Ti�6]�G��j��>�8b�Y�&�Ibi�,�����Z�Ṟ�(0�u�LC�sG���jPIK���#D(��0�$�Nq�l���9��Ͽߏ���㮳���Ӯ�뮾:뮽�뮺�뮺�㮺�Ӯ�뮸뮺�뮺�:�u�]u�㮺��]||{{z{u�]u�]u㮺뮺�u�^:뮺��]g]u�]u�뮳��뮺����]u�]u��룮��㮺�ۮ��n�뮾:뮽:뮺��~�_�׷���믎��N�뮺㮳ۿp����s�oB�gZ��W=i���K�֗�����[/�aZ�3l�$���1#O�E�[}A�VV�5.��6}�'��&�|�Úf��h���"���a�V�[kK��$5fd���`ɍP�,i;��C]�q�yZ��<40[ݚ�:�a��Nu����o���|:�f��Lޛy�}2g�<Q�;�m�~�u[������㜫i����Q]8�1<�S���(7�B��C�ԓ�T�ɔ�`h���_K�3mR��nt�3ڴh�����RX��~��bu����l������ZЮ��"\{*�r	��j@�S�j&�S혅\��՛�����1Qk혎�����)�Z���K��j;�!�� ṱ�/�Z�Wf�6u��Sg�+�E�~�Q����R�y�Ξ:|K���md����D� �S	Q�zN|9�y�Z"(�q����UeND�̊vI��5R�s	/M���ؕ9LP��pŝ{j�*��V, �~�`]	�X��" ��;9��P[�oz�\^{���L���b�/�'m.[�/���������iU�e���[4���d���0�c��,정�;��ҵ���sXc�K�C3�J�L�3��^�^Ζ�UƟwrn���8����.\kr�P�P�X4t{�;Ԙ䈸'nfNYg�u:1���n�f�;y"rvl]�t���>� Z��Vͱ�hA �gd�^>�����Xigh�(�5ٍ�\�Ѽb�nc�F�ը�Tw�f���3��jAÉ��.]q��k\�㗅��Z� �U�|)�=���59O��y"F��ו+�i�wp��+.|Y룂wii�v���y7���$���1C؍SL����T���H".<�	����j���ͽ
��ȧv;�(=^�m��T�ŕm���E�坉0��Y4d���^�{�Wm�,�:�@�r|&���9^�W�l�+}�"�Tg;Bͪ���!vME卻u^c5Q�V���Z���8Zk�B��CB�\��5}��+7�D��(fb��l¸�`��}Pl��:u3pc�_Z� @��^Q�4kwl�#�EXdͽ6�]+���e�7�bcr��2}�FJ�,��]�����#f���ͥW���\��ՕdJ�����9��m��G[�j����P9�:�:����dp駲���p���}�m�Nn,Znn8� ;J5-ug����d�lVP�kU��rA�[T�f��}��w�#/�ر��'��v��9z��@�~n���8�YI��r�ڧ7�[����t��7��5��,�kd�[�}5��t�TL��7�^P�|I;�E.#�F7�B��[�O2�˥IR�)NǶ���a�X�[����aɶ�ⷼ��-K8��F';�����4�r��6���!q4o�T<iˊ�t��<n��
����Q��!��i{��@��v)���tU���蠪��4]Y�}zt'�7����n	;Ay룄qF\�b�igj���*�w8�=���r�%�(U�4��^S���'�;�Z,��]�eN�H� �$�MjK��.��C�nb;b�Su`�.��wy�!�>CaSd$������wk����T�FXx�����b�R��[��*o���`55����e��<�R�Ɍ��3�Mb���+�S]���VS�.ˮA;�Z0�nP	��ތŴ�C>�4T�ipw�ȭ�
��I_#�P��M�ڙ���ǥ+	�wK�ݒ�iݭ��=��*�fA� �zc2We��e쩘Z8�"A]��0d����@� ��ɔ��e*
w
7}͗;3vpDp�x:�S������9�&ޑ�(ꊥ�9f�
"��?=��a�isk+�j��r�o����q���
޶���7��N�b�PuI��N.~���nM�]��` ���_�� ��!*c3��C���>C7��Y���+~�o�zY$T� �)�<EP��m�|y�����ˬ����e+�a�wkp^�'<��,���o7/����<�n����+�Xy~�Qч$�i��x����U�#����;w��`s�a��a%.8�.Q����f��TSH�'%��I'k��,���!�%�*�P+U�V�y0Nq2�]o,����{Zj���rx��f�-���؅��Qs<w���<��RSu5��\s'��QsNR7��WFH��K�����K�&�O�a[�{�q������ߒ�9XP�̓�5R����_ ����L����������O�����U��p���<;�G|[)�%���Q��u�y5-�'��;f�Y$�*T
.?�m�Hny'*i&
ch@XqU7�$�?�ѳA@�e�\h�B�S� ��w6�B˗A��hX�����+[��]�x(�&��&z�;�a�'�h1B�Y��h��t5�An��s"��6X����V� Ŗ��5j���ui.]���B׻�;�k�� ��#�NZ̃[��DV��K�d���Fb��4n�����ۆ��gu�����E֐
��,����k�p�A�N�U�%���/v��jJr���>���!vR���A*ѵc����^ww�Ldj]�j�{�v�M�-ީ������s�6;��魥�S�Ʃ6T������)1&��X��]p���;����N=d�d�=j� ;4mY8������T[)��,��bя��o��OIU�<�F'I��p��Z���$���,(�*�c���U/���2�,J ��,��o|�2�*�G`��Km�+�F��UflȎn0�j���D��t)5X�.1���ur�mj��b�T�wڂ�Z��qL�F�֕�H��3k���:!kx��z������{��o9t�����^�Ngoԗ#MSI"�ze]���Ud4�1�8W�uj0�ף�4�����o�>����D)׏�b��p���	�@˘	ːA\�@�f���RX��&AI0��yo���	%��ƱaI�!˂A0�I����Jl7m�B%�[NX�e%)��vO6M�J���)r�$L��IR	aK��Kq2%ɘje=��"��f,��$V�{�u<��:/:��B�)»�N���ߺ���~�7����Ƿ���׌������Pr�O�s�5�=�ד�ސ�^��y܊�kdO� �	I�V�2E>n�9s�2����׷���������~�:��ϥ��44#�U����
m�ƜcH.p)���t���������J���v]���i�!�I��'yl���w8�TaCN�˲�*�T�C�"��M"�IĂ��BM2ci	�s�C�y7gfy�`~Ɯ")�9t�i��(ޙ|�+i$�Wx�����~o����������lz@{�x�Ay��<���оlP��:م���8����P�]��YJ!H��y��!<�ck>y��($���*���h�9
T\z&.**)���}}u�Ǐ��QTGκ:��\�z���R�wg���ޔ}P>�p�>!*�!�OI���x���q�������}}u��צw�>{ݾ/_����*�ODH��)��5ug><u�<�c��/�OOo�������������|���B%Ԟ��f���x�I���U}ng��w9p���P�$����PQ[�N������q P n^T�*,�V� �ķ���^�.Q�#\���Q��G?����!;�P+��'�.Ry9�8��F����땓����%U^g��y�Ԥ���s�^�Њ��;��*.Ć����I��!�-�R�&[PP,����+�)�V�M�RȻ�a�2��s{�K(�I��NE���	��}�bI�CeR�u_ �QE�J@M(�7$A�TB�2)��_t���4!�!����އ�ǿ��]6A��!�����ПqYA�ol9��lYT>�n?ׁg�dn�\qS��GOj��+a�c���c��S�0�Y�-7���NŽ��<LҨYc�Iu���Rd�Vkb%2Z�����^ �Y`�������1�Ħ�\��yfZɵ+�7L���啇>S�����沢��t�q�N��\�6������l��95�� ��Z�����C]�;����5�"��w�=����B�Е�*�R��YJ�-�5Zt�J�)��F�L���_͡����P�iA��J}�}>�p�;w+I}W��RS�AN����K�I�X��-Ý�}�Z �UPF_��˷;��y̭�{��y�H�&�mkt��yh�(�C},}~f�զb5;�<[��U���#��{Țac5ݲ���e�E�S�<�Rh���!l͜ғ1��Ə�w�v�WY�roD4�gM}"�6��h�)��0�� �*��Bl��o+-����p�L�gmmLv���9�
�F��]ڦ��8� <H&^<��Qw>����:Ƀ��#�mR������t�u][�'�`I*f�G�aq>�X��Z��[U%�,�.VF< �2��6��Y'�c��uc\�f���q�ԊEg����F�4�hjTr�2�j�A0.�)����u�u����ȟ<��߹�ueo�z���]�����S��MD6_��Yz��[k�e{uU&M��.�~9��X5�;US}5�� t�8����n�^b�����XR���dK������������T�˕ZHƬ$6�(�i�"��u`/����pb���ey�T=��]�Ao��l{�x7=�R;��:���WU��/ڞ�J�����_��=�>���<o�C�׹�+�����/a�!��m<���׾�f�j�t�]9���{>�o)*���g
J�H�+y�)�|^����ܧ�u>�q�e��4����Էk{$m_r�Ubq�]���j�f�ӕ
��M[»��m1�oY�̬Ե2�W��Z�Ks�.��n��\�����x�[;��M0��
���ռ:r=�b{�Ea%$���>�'�%6�6l�P�R�K�q	��_i�?�{T�ڨR�L)�f��w��E���Esc�]�[��VeffB1�!:��f`��t#w���M���/�kRZ�'u,��-S^;ͮ���}MFYw02�
��ӽ�ȟG1{��z�Ȟ��(�Ҡu�V�ZY��cH�Y�깁��m�Y���$wODw�{teY��|ʺB�K�,U}��W����<��������2�-�
�q��F�f�i�ׯכ��$�"���?��ʧ���5�^J�I��g�ѡ�3���>�S�G-z��M��ٱ{�7}��u�	�x�M�ql��S���ׯ}�7~�%�kжk��c#L+	:��,!��|�z�F�:��ɌT�5��^�?=uƾ�lSoo��3��w瑊�ξ�ʹR��iC�Q�J���WQ�F��jm%δm��p[�6���Ww<Y]]2.X{�-��d�np�fE��o���Jەã���xSdO�Նd��ꂹ�H��m��5�$��r���b򆔭��Խ�dfB������ٝu#�o����p�,/�e+��͋���aޏ��џ?=ϫͻG�'�O(��ʓ���&H�MU;����i6͗��L�Xd�Y�ED�s��O�����\S�6���M���+�sѿH�`E�߱��a�mg�i��(�//b���xp��{�n��4�)�z@���W@Sη����W:���8�ǝ�|WNM���G}�Oo���#�V�y@m�i�Dd���|��w�2�=j)�a�n�N��tW�P�F�H�p��z�q�\���(Z�:fȅ�AD�}�p�'$��Cc �<������:�b����M9��Wq��-2-�6j�f�H�Ʀ�#w����Z8��-:�{$֤��Ɇ����{}ެ՝t9�]oMƷ�L
�FMށ��XK�=�������ĉW�]qb�sZy�P�o�B�2U!��1���wH�P�M��Є�܊K��ؒ}�	� V��\ݓ_Χ:R�Mt�#�veZ�q���m�"+�T�j�i����(��`@���Ջ�H�]P�@�� ��LL��bf#�A A"	i3<�v���,�J8����!i��$�~��ͥ�F���Ŗ�}�H̩�v3����G���Lwjb'�.}���B��Tr�Yn��QԮ�va�EV������D
�s�˰��|�e�Edq:͢k|פ�.�T���|'�Wu�]�\��v��:���ٲՁi��L)���l���
�K�ˤs��*�OǶ�h3ݾ�RozL-��l�٘T�Y^��r�08f�����%C�y�Y�1bXW��0��)�{R����5]��ޝ�驔P����w9n�V���\S��>eq�UP��)��ǭ;QIU=�
1Tz�	��(D
`�kgfͨ0RUr��pK~��>a���)���>`�ϥ���'�
 �3�2s/��U���&�'ď�����+Zb�T.�^�u:�����#��`��O�gӨ͕;�����;��{L[�T��p��糃�e�)�9��X�M�a�� ��0�:@DD3$�O���o�W�������W�)����d��
K����b>�m��7zWc�q�����ﳘ�ݖ�l�Ïk�rKx�!���3��	��&��e%u�)���Xѡ���{���QS'�+��wV> v��Qy��a��9�
��^}h��v�s����KњP�I��rg^Ĭ��"���b5Jc��.�^)+e��5�W�C;�`b5;�V�%HU�[o�ω��[�b	�TV
�T�-�����6�{݄��mfx�m4}��ַS�ܼ��e[3�|�Q��{��X�����.�wxt` ��JT��r� �e}�exwpʱ����S��E�;��uN1����!z�S�D��0��3r�sP�f=w@_VI�+0�T���K�v�m=�4e♕l�j���Z'�%Uf���8� ����1�4Owi����ȶ��L��s�{�t��<3}L�TNٙa]���w�����x=d�4!E�ہ��Y�|��u)��"����dv5��نSmq{uhł�r�Z��@�C	��{&>�����;����������kWA�Z�DgCi��!����.����<���t�4�t�4��@�s
 |�Qŝ`ݤLc�Q�*l��jO��:�k����^Y���s��^ee�]�M@�)-|����n1P���M������o��p	�b�~�$g8���w+1&҂"�p!a�fZ9��x樓��R��U��L�[�wE��sfn�BY�@��B�Ɖ�w��*���Q�Y�S�U>�L*%�bݖ>��R��s��w��Ҙ��[�
�Ak2�u��Ѥ��B�W�m5m�hD9�{�t�|5�lx9�/�y�ߴ93^k��	Z:{zv��u�o��9V�\�[���@3�������y�F�8����%9ڽS��|�<�ES�bi���Sv��&9T�xK�*�nF���{b��'���w��|��By���3�r�LF]މ��0�'�{�_|y��v� ۗ>��Jn%D���ɲ�w*������bn�s��}O�����hFw�gY;w�m���EƋ4<����Y�0`�W}lv����wε�U�I� Y�o7tr�z|lĸc��+�+�4�H{C�W�~�Zm��19�V�Tӻ��.��3b�ex�.|�}�M�Ϡ����p(!����t3f��]V:���_y�N}$^"�^�Ά��;\�[e�λ8��vi�Ϡ���Vu:0��h�jI�ck=e,���p�v�w܁<fČ�8�r/�����;��z/ u���~t�E,0�ҍlLϑ㳕 �2��`3Ct�z��{�Ƚݞ�R�I�]�(s�ވ��} {ۄ���<c	���߶��}�p�����F�A���
�W�]ް�Z�E)A�QY(�Q�g�o|��![��<���~�<�f�z#��F[�u���,�i2ǝqS��J�>*�»ty����*՝F�#�������y�:��݅^�-�-Q~C���lu�6غ,X>$���T�Z;��"������5�K�L�E���Ҩ@� |�{��<�DS�n�Z �WeF�H�T�ҏ�������M������2+Z�}]3�v������GL�s�����GS�0��x֍�:��M^d�@�%�3@��GI]�mD���y�����n�?�������[�$�H#�j�ܓ��G���s��C�q��j��Y����r�>��ﯹ�c�ϧ��U�>�=B����h���
�a����u�����h̍Gj�ӛ�t�f�G�j�X n�D��ӍziN仦�>-�{>�v.��ʺv�\��^�O	�jڜ=G<��[o�X>�5���V�����a�wu�'۲#C�ؼ� �y��!o�	��j�R�ը��Ƌ(Ŕ�!n�.$VKY��^����Vl�F���q��� u��&�a�E#Xa͍!�X6Y5��vq��a��������"P�IƼ�r��y�bq܅�Lv��"�ןe������א�޺���
�\tUTTI���Dp����'��&�Q���)�bM'_m�U�
�t���/�^�b�>6e�9k��mNp5Q�u"g�=p�s��n���9wn���p'z��b��1���-��f�*<��QuZ����v→��l�DuAʗ���N���-$��T���9_U�`J�r&�u��F�a����s�3�3y���S�f�����\��_U�!����H���ђj�]�6��j�@7��<�~�Y�5x��m^䣒Ł��	VUS^�֪Y���'�34!��i�Wg��f���rS���Rj�j�S�
��B�t����8��8�vVO��U"��Ō̫N��+^PS���t�/P4ccl���M�Ŗl֯%8M�׻��V�ii�Y~��S��@� D!�=�{��a(�re�\��l�09#�ͩ�2)@��� ���y�sGd�8:���=���v�E
�(�-z��`&�yY�n�쬤ϖ9{�~���:+��RE�g�h��'Ӆx�s�,o=g��ޱ��`|�>�֪o1]��"�3|o��|�{{O~��!�	����3魧��Pn�_�G����y��7��TT��23+[�$�(�����{O ce���<�^���A�d�	�o�D9�7o�p�
܆�Y@l�hv����v����޼q�%@��W8���rR�t�z��\�$U"�q����Wv�y���t�e�u,��L������S.f�`$�&˙\����ǡ���%M!{��eK�$@_pu(�͡��-�y������WKW��"�[[z��X��j5t���7v�<�	+���κn�7mF�NN�%��V{�<��鮕�M
��թȸۮ�Q��V_iɳ|u�2��b��T$��Ȗ,`�;2'ǲ�w}�$�[�YR!��j�k��Q�v�x��R�`�� �	�$�}�lu�`�`�X�u���n��_V={�&���K�������,�\F�:J�&��+����b��]�J
U�����k�N4K�]�(_"�ʙ�����]�6���<@t�>�;��2�Ҧ�|����B|7-��m8�yƳ�������e�҈�Etkl�a
��T�{�}��N�ot����
��1 ��*ҏ*��]9DX�;���F�13Љh��s���Y=g��^�)m�H*)��e뙩PŖ�j�a�1W,/�_� tH�5��IƲ�Ӓ �4�V���T\/w�j��ŕN�ga��5q{F]��y0�<�Ym���D�oTP�� 9��(������H�YqRYA}$]���/�5�h�w�oN�ӻ�Wt뼻�]���qPO��^w��F����%krvG�[�a�r;A�VX��9q������9ͬ�)�4�1m�8y�l۝���!-��(�ڊ�=8ڔ]m��
'lW����s2\4>��k�������}z��B�_b��)66�mK�foQ�oKWӔޡ#����Օ�-��F,�[z�B'�P�֧�^�J��VY�tr[�J;�-�]�o�Y�5�t�%��w5��#���{���{�`�A*��m
�|l����T�����(��N[[Fr��뵛�|��8��Ӳm-cOTҘ���Y���4�G�����|��o�=Ү��2��m)��'��*�֧������7��׹!��K���[}�����9� �Ȼ�s70��aK�dp��Ԏ��mЊ.鸁w�2u-��Z��]ϱk��F�=I0��=62��O~vz�LN���Gw^�
��tz	X�Z���To�q�+�}�6J]uT��U>��&�vA(l'HoW>i�u�ѣL侘N�i+�{Z%�{�tF�h"�$ �$�A��*(�ϦȎGs��{�}R�&�E��#���Z���W"�]�<�,;}��@�����������������������>>>>����<޾|f�D�G�>P$��$�<I��U~xK�������NT�9QDz�zzq�����q���}}}x���ry�wlwo���áúI�����W�r�$�M6K!�H$}
&*2.2*2.....4G��cР��g�����IH2p��ȹR��yI�s�P\�s@�f%��Q�%�:8�ظبȷq�����^3��s�ʪ�r��r����xG
����f>u�´��D��nݼ����x�q�q�}}g׌��O�r(��_;�O�+����''���NI(�TE��A����£��=B�Z�wyh|r�	.�Ȝ�"��Q(�:UQTp�z,��:�W"��xݡ��.^E���>�p�*��C��ω1&)�A4\DD�>>�Ǽ�}#������ׂ�&�p���lΏ�/�sw�M��U�I���k}�"᛼75���za�8<y���<Լް� �x�����>:�Y�I�[�� ���t̃�(�|�	ϯ�Z{,�s��/�� +P�����Kp��(Q�]��7w&���[cR,j�~��zgL	�u/��K��,^��`�������!|���mj`�|\_Q@��1�.�p�:=��_%� �bc���M�O_Zܒj\7�.�p����P�;�N�(�	$��&������+"�l����#|�F2s��w}���g묿f�Le���U�d�$�@�O;�#��ن׌�F��4���?	m�|.:�ܥ��y�f�UWs���+���MÜ V@�r��/���P*���� rd�z">�'��s�"�?�@���"�k�٦P�sr0���倶,[�<��%��,��*�
�x��?rIC����Iݼ�;�Xz�p��L��uϠMm�b�cxf��,p9�k{�"��|��Y�����g�z;��茣s9�9p���~o\@��s�d�k �P5���mo��x��ǻ؅8�M���DI3�qr�\<���WO]o{y�hO8�ż�3���J�k}��	F�M�� �F=%�'j��)t��;+���R�ｙ^y��@j+d�ZY)t��ݢf��WZ��WJ�gV��G�|�������]y~���0����g]pɽj���.���q�K�ORݷ"u���9Iq��t3(NMa��[��A�B$!Aa!
V�vp���{�&6
>驁�@Ȋ�NmS��V�q弣�BKǛ�/�S/x������6��עx�Hp������ !�\�1X���°Z@2;�Q�|z�>�>����m���ʐ���[ �Ԯ|+�c�z}�
��1=�g��p�A ��.c�/��b��ũﷰ��,i��p��(c�x,���T����2��|-���{k�vuP�O�E��{�`�C��)K��mon�<�0�=�v���n�Ǘo�f��������*� �"zD#E�������X`Q�$��$���[@V���`q���H]��<���%繭>Ӽ���nu^qCA�H��?{]�5)<@�V�u'KY�ȟN� w�����f`���$�m�4c���|\�0��>���OҀ�_�0>���0��W8&7�Z�@HW��>�NML��$���w�J�u�2�tN��;���|+�>,�O����H1����s��g������G��&%ڣGw{����	p2��=���`�0�Z�����~���65�@n�0��Lx���r/��@WJ� �J�3KhtTkV��8���W�)��D�3��b�;P�����ħE�`ņÖx��.�Ey�N�|�37C�p�n�U��N��v����v�$�v��9l�a�\u�l�*v� 3r�*U�*���'t+�W��`<@d���$(T�y�m��TCi�I��i��t��Ϟ\M�?��d���L�1Sh-�ޭ��*d�R%"���
�TB}T��x�s�s��A�l�G2�ow=[�뺺��ղd�m����[_C,���|Q����@Y��|�LO�lNy n�?rMB�8��	1�ꏚ1�yE���J�����Zb��RJ�z�%�O�	Y�ТЖ�̏������6\j��h����z3�y<����|x�5�Yp%��lXҠ슟�� ��Q���(�h�QH����.ivfʺwq���'|��~&�@&.X
/��n�-� ���{t�D[m�@W���
$z��A=��m�o�.me��'��0��@H�8�$_��pz�|�Ic��r�=��5W-0���^�cyiƫ���g�`$�ϝ��mq� o�N8Ì��6����[؇Z�>�8�TH�:�L{K�>�h�@��֭�w�hx���܉��8�À:��>��1��(	 |��,gwP��b�)�!S5��y�ܵ�v[�i"[b���$��
?� �����W�G���0� 7�j&"���t�!�?��-]p�{~���-�TgQM=��S (��b`ny�@��Li�~�����9 ɨ������!}�z�W��k��} ��$$5n�&u}�u_��m�,����7���7D�%�{P��*������Ԓ�85>�F�oX'�Q�1�/V�3���n��/���Ʋ6w�u��K�����c'�
� ����	�>+�ɝ�P���a�C�����3<�hq�}��g����s��́��P$�p>�F��ψT�@V���}	�=� Y��͢��(��p8��&m�1�L���. RXsTp��D����s@-X���{V�)ٍ$�+��#�|��� �o0d)�f7�a>���� h"���Ԃ���;�>��-�&�0���;�<7��40��>�T�j��:��NA�|\�x�����������b�2,f�� �e��@i�� �4MB��dC5��H����$�O�'>D�W����}𺫼�#����m�-uk
��*=B�-���	;�ƀ�F:H8@F���1�=y�L,��4O��`�d��&��NT� l��>�c�Qşyu{�,�b��ѵ���vX�-��(}S�7�dWT7������'�8�c�3cLiز��_K�w�5	���҉5�#�W�>�z@��x�@�r���o�l����3�d8�%r)�������x��P�
/֘Fs��at&r����p��I��K`�Wv^J��@L�!J@�J<@�̟8��7���>y�|c��ނp5�R���x��m2`!�e��X����Ž=�.[�}Z�˯��:]!pv��vq��hG;9��Ԫ�$��jf��ɳ聡�W|Y�����e�F!�KFk8��W�9�#��fNM��1D��nN���n��g�wق�n��/�����H:�s[ķ��� ��!B�b4!Cy���ZSUt�I�m|��� &Yi���q(�~;�/�X�Ϧ���S^�	���ӿowO6gmm��	m���f~E������\1��1� � HZǌx� �~=(	:d<� ��Hהmê��OVF��,��kr_����{�!���0ED����`o�� @�n�;��%�-��L�z}U/m��UֽoO�~_?321���Y��I͸�􈱽2Hx@���,|��+�>3���!��e�����:�L	rD�&Jǹ��>� c&g���,Ĉ�,� ��m �az^��ԁ>��v�L�׫mWn�ِ�w~���@�C��	8b}W"41�D\$<x�#F� i��歹֗���xk���J `U�d	�~ Hr���/� ][d�|*=��~�܉�i@�Z�mx@3n��ðǩ� �9�J�G{�Z`i���ߐP��t���0>�>y�����Ɍ��5'���P�䬒�X���oРW�x�����Ā��h�����H��F�T�ڒ-�>홡c��ؔ=�#n�yx�텖;�F*v=�P�]��5D�@��qeO�x_~ K�������Ky����qZΠ�f�$B����T�L�7��|�/�Xx��M���gp�7�	�b Y��I�Y�@�:��R�jM_Z�2�t�;+n(5�MZ}w�sbf�u����5��֏
�Z;3�bs��;2�K�S���hB��(@ ��dC@�~�Y>=�hO�@����g��2���?�qa��Ⱦ[�~Y�}�ǵэV�݁�w*a6e����栏��#f�c�CE�ī!�ׄNo�k��t&&�P���a�����k�ܙ��Pj������}T��YrjP2�j�`��_��H:����>D�8|�QZ7�u��r���������Q�����{�sv��rn��/�G h���֔��4����t��.�N�z��,K������xC�B��i��l�w,�PШ���$�m��zd�a�7���<�����1�\Sr���׈⡼�X�z|W��>�V�
	6����{M7RT�Z�>��q~���]qB�~�#jޝ�W"ցQ�n�iN�<X43�����ab�+�$�K�����)�\%э<��yH��\�,��[K��U�Uk�Ų��9��Ƿw��� A�8ʽH�_zD���k�G��:���b�/��gs�����y�h}���P�q���GX�9�fޗ����=��az�w�2Y���8�� ���1�K7#��ov*󁿏]t�.v]�s�%�PLHc��"ε���9e6r����ĸq�M�!�����+�R˺v!�mK��⢈��r�t�Aɣ,�S����1u���Z�|;nb�QKޡ��wy7�.N%U$0�\��B� z\�H�tCwrD��a�ﯟ1/9~����a���aEi47�Mz�_v�<4!�s�1F�\����st|t�Y�i徟A����7�#��?�P;�I��j��Y'8�����Л[�%�h{�{yϢZ�9�j��!�H�FD�t_Ga�Zzwg��\>0~
�fl;�Z��:ޓ��g��{��ă0��P���m�yp9�b��=��9����b��cL�O�B��Fq}PS3��*FT���k�Q�Smz�<o$S�B��}H:wc����F�gI�!�KU{򸢠v�ШZ�����]��N\o7��ݬ�<��e�I\��|�l4K{i�s�d�2���'��0��c��Q��h��E�[zUp�OB�e
+'%�CD�]��K�{�%|{��8-T;��tS�>]NHt!Y�_�o�y<�2���R�a�\��ܩ̘_���yw�^�#���@�V����j(�wD7��۲�ޓ�dH2[9�e�!��W��ʀ��<��6����2�s׷����?ٿ�%���t[S�C�wŞ�W_:������ܝ��k�^��|k�� p�@����
�����+�R�Ǟa���C�͚�[��
�`QT����mD��0���5ҕ��xc쭨Ş��q\�+	<��ޭL�{�ih�8�V((�
���P����:}��_v���s��9-���뺾BT�2K���ö������o�{N36q�͎n��}�yߞo��/�I�9��pd�paNpx��7��g�������O���>:�uĒ�OόQ��s��w�>|�+�W����@u�!I�8=a�������^��>'�"q���$	G�ǅ�����@TϢ}�q]������]"�ĖJ1���3�!��v����,��\PM ������C�qn���kJ��alj�@}�H���t��_�Kf��dt�f[���6�[Zw�gZS�q~�	0z��'ōGS�Kל�Q�aX[���k�i���9�[W�;�qJ�;���(���#�I�Y��e=�6
[�3��ѥ�<%���o��wď�|���m-w,4��A�$u��Нx�0���E��=�*�_1�5��-�Q��{B��OՄ+5�:􉆯�b���o%	��:-x��\Р���%���?=�q%}U��uze�G�~t��+�>d����\�!����|u�p�� ǧ�1���.�S<.���{G�HWG��p?��jG*J�6l��	5#���8��&^�=O�븜�g3��l������f�6z/)�"�=�Hj�LShٓ�����ʗ����	���K5��*;��`%�5��uoU8���y�iu�l;��VZ���BƵ�)�s�\��6�g�WV:w�đ��OS�4Z�b�����/���J��|^v��9����ve��-5?� | �� ��D u�����hɀ��(ϕ�غ_�d�χ<@���/�@c�Aa��(~v�Eg��kS7�DQ�<��k��.���v���Ź9q����{�&��	��bqM7O���9'��Ͼ�1�Iv��*�Omv�OA��md�����x�Ty��5trO��s�w9c^�;�k����9�U���K�n;��q��s�Oș����O��L}�3q]y<�_��2gM�_v�wik~�,��r�lXo�Ue/�}18p�yZ��`�#�ʼyg�������2�]�c�ɂ���I��v^mv.������c�= 0ǰ̌�!�u���R'k`ϕyl�1���0.l��}�<�"NSj��@��c��|.1���&��[
j��.���ls'��Y�)���goS�D#G־�aެdsW�$؜cz�&�fY���1ٮUVBC'&k�;��Gܹ�K��`��GF���Ý#{�`c@�/����ثu �q*�ٰs'E��~��.�u�vj���
�`��t�3Z˟�#(3�с�U�ÅڼɪxVj�"Mk,O���u 0Εe9hm��M�{���{"�=��"�ozt�tY8���$�	�I�S��!�g|{'9I;ϟk}OǮ�V�[C��'|C���*�>]�¸t<3��X�ћ砛����H~U?#���2�C )@��J4�@� �����_�Y_iP��ڬR�!�R3��$��I~^ &���q�붋�HW��[�o{VW���H?D
2�D�E�c��~�~��y�)�`kP����<O�F	��.��{�ǲ}]��馉W��?`�T�B�E�!B-(&P$��۾�2%BZc�����,�	1��L��U���CU����LI���r����ٝ���~Uq���kss,���ήy�w{g�a�LLc�Fc��~&��aLI��3!%��"%��w�����duzh��1��y.�@��Aua{Qӗ��W3���Ee6n�^�55�!U�鳅o7m`,U�"|�����+�LMT/���w'ܑ��Vv)P�Z}"���NJ���T��H^mqA�,W��>47�I��`�����$}�A��57�lʣ���oT1�Z�}ZǻD���:p�P�7rӐ��8���vzhp�};�g3�9���fl�c��v��e����`��9�)a�#L�c����<&��3"��9�a6��!��]:^�.�������(�OcD����e!����XA�q V��}���Z�4.�{��E��&���C���XV���y�+��I+u�e��ޣV 9b�Y�2d���|�f�6�LՍ.����!z͸Y[�	������N�K�D,�]7�����P�WSo4L�-��	��%���lޤD���t�vF�����Q��͐�e��՘x�n�U:�Ըs5hM٠yE����t�F�@:|��.�U�Ӝ��{qDmm���R%⢶�>ٷ�7�bT��9�u<�s�!��Z�_]yIM+�;���uŶ��'��J׻u��1�J��}�goK�E����ٳ�c3&[�`�Bcn��}Y�q��Gr�o����Vݤ	c3,�Y/�.�r�v�-���\r�S�EJ�7���A��Û�e�wWv�H���Cn�}+��Z+�x���3{+��0K��w��+	���vo{F�9��O��'}V���]P���t%K�Y\O@��ҩ{ p�,��!����I���_���:[^R�`&�������Q�g.����w�rYJ�ަV+��r�������全-+��EdW%ʃ(�1񇮷�F�9�ـ"-�9s��U��73�s0��y-ڀ���#�Z�Dà�4�}n��y=ʭWۗ �MֵKi
�w�-��t��e�"�;Uj�)�.���<{B�䞆	XN;6Er�GyZD,<�����〸�@�)�͇,�8�3۷x�0��
�rbk��.�;(�䴴�C6�V2�e��b�4�YMRV�pܐ�����de��W���I�롆��Ѩ��E�����/��֛7�_�^��簶�Od�^tf�5�=��(���kg[S�R,��:�y&9��{.�UW��s�{V�HSa��,d:�Ԏ��ὶy��al{X�i��Jk�ZZ�O9�H���e͘�행eI{�,YL �t���\;�F	y\���ZI�l]�ެ��jhR��]��9i�ӽHAb׋J=���W��^� ��(8�rG�Ժ��K�9kXwZ]�r Ke�3tEC
��u����F��r���f�u��jrb��M�����*ǅvdʖkB�K�I��D�w;�X�Ը�{N�3.+'�,�,�2�eg��Xy��T����|Nb��.b�cr���B|��y��k-f����b_שG�2���#�.���U��&qz�{K+	3	�qE�\��u��YPՆ�֭p����C�Ho'�n���j����B�Frc5� ��ۼ�s��N�{���L:7k\�h�`�	=g>�"�"��Q4n��uԾObՈ��[e�ޝ�H�Ee:=���ӌ;1��9)�ɐ���5:�w�����'��*fhN�t��=W��YiH�+b=ܰ�2vN��}���W-#��F�R�BW�)��$a�K�m2$��Ih9����#&�iCE�D�8ڧFS`���e$J�@�v�i7�-UPH)�	X4��Ql*ۦ(	))d32�,�	��[7vZ���
��T�2��d�ZYI-fS�<�dW^�0�������6C�@I��Ka�M�F�-�޺v�M��f;��E������iQ^�R�qȩ�z��U�"y�B:루�� 9���~>?q�tu��^3�ݣ�"9<�"�3+��W yk*wG�]�z����������q������Yߡ������S#��S�UAJ��<xL���{x��㏯��q�G��}x��RW
g��>$��K3D��E<HU��O������{�w��8㏣��3��=��8��8P�0"�"��\��:F(��8\�EM�OO�������q������|��{�8lw�:�MAH�!+��ZۙQd#�"�W�nF�*��~nݼ����޷���8�>��>���D�p�*RK(��HUT�"}���7�&�Dd,���(���ȞD%�w�����,���+�!CO�Wx�EEGe]3���D8FFӜ洢�:�UN�A�
aP�NeTF.����_���/�'�Pc^�g9-mt]c-əy���6rM
�2Y�XC}�;ӹxd�ه��Qoc���<���iŗ�I���M��u�nCe�2Kj-�y׌@�����bL��@ѓbpg8�4�(3�9% ��/�����s�~�p0��e)L9�@������뚥����N�|`_E�k�'x�oN���FސY�['Ͼe����}���>�<H"CYt��)����7��TE���gd[H��Vz»if��R�Φ�uZ�U��w���Fғ��<�#-"��3�E���}����\�մ��dmxؽ�~K� ���&(3[�gZG�0q��^Z�ٳ�10�% ��h�橁!x�1l�"zE���5�V����xGLf������;ό�n��j���6��zp��)�<�o5ki̤l�tc�� �;B{��
O��f����
=#5Ew�:�B�|�򜈈g�3��݁��w3��=��E�B׷��/�%�����e��q��y
�T�uM�'��/U��Ɏ����Z4�N�O:�������T����+Ҧ����^\�<�t���z,�G>�\}��2�v�'vq��{�Уq$2��Hj%� �!�EU/����6lń���sQ�צ�_JqB��[O���{��<#���nl�i9V��L���M�y��rFjG��]�J͌g»� ��4��H+�7���U&�����D�=�*j�������/�R;�(��
]ƹ:�Ӽ8.��N�0��EW1���k�̕��ju�2�kݵ�qY}y'@�_tI\�e����m�.�����ޖy���o�WX�ޓt�OT���X�?1,�� � C �܀)N�^�$"	 36w��}7�*������1�t3.����W#;��w���D��=8�!��F�T�bx]��./�f�1��0�㶽Lw��¡s��-e��=����H�*���{O��<$93KN��61�'�x���h[��4����;!�G0��m.��㫩2�: �q>��L�t4,�}U��w|�Ȏ�~n�$@M�#����M�)���v��-�ܟ�3�ɟ���\���۝��(�_CCIe|~�͐�d|����f�=1��V��/y�_�~b�-L�Ći�S^�r���,w��3��vy�a��7ϟ���a�|�|��|�\���Id��.��M@��הqª�aA���ݜ�] �����(��\ځ����<n7�G��}|��}�����%���d\�w7�̍��A��	�Y�/p�:��B<N)��������z�cަds��0�~S?OU.B��=o9�C��c�M�����f�8�6w��w�kٌD�6ba!�)�29��c�I3�����������d�R}� o`G	��zn�)�@8;]��y�BmQqkw��l��/;
ɟ-1-�{�B���N��V��^�m�������3G�>�����jG��`SV�|��wX�tNS���O�ڲ���6E���C�>��׾@{�Z��y�tuU�um�dSX"0�g�u/u���o/:cګp'|K�����r4�0�����b��E��f��@�� @"�1 R�d�%BPpdRC��*ЃB����g��y�����K���������Uz���ؒůX����h�Y$��߉C�w�s+���K$���N�ݏu0��.��Sg���w�Zc~A���H��/L��,)�ފG�u�DC=�Ƕ5�g�o��,^�J$��ِ͚��H
A��49J�v~�O�	�tc/wz1�������3Ck��J_��7�勼�+�f�B�"[_L�m�&��k�_|�����"�A0��J���Q�#��J*˺��`��T#[��5M3"Q>�Z�`�%Z�l����2��2����2�L;���1�����y�u⪢@�v;��g�s�m׼�ໍ�?c���o G(M��^S���қf�.���2.���{���v��j����׿+�@��_�̐W3� Eτ4VEǟ{���E�{�z���[/���gXV��μ����zn���>a���W�v�'�RQ�жA"�K_?[zSzE�M�i=:���RTBʙ�Oj`�xC-����N����شx'.�#[3�0<��g�ǽ1��c%Ca�f��\M��Ļ���٨vN3=�o�ǳ�K=�dek�1�h-{gl�P������:���zQ����^�;P[�\����ѭ�wc:�*��@���4��d�J _E,f�'vi$T?�]�1���>���}O��W�ƥ�8]�䝎{p��Q�q�D`zNL����������r�"8�� ���6����j1�4bChɄ" �����\�ﾷ� �G/֔?zj^��t�c���&�{��{MH�Y80�
sa��(j���mu�64���ऍ�P�>�Uly���mj}����dLo\
�}3)iq��>]�w?��<-�ᵹw��P��T"���@˄7�:�"` �}Ϡϖ��1a�ꍞ�`[kS�.z���S����*�\��!�����S����p��� X�=�z3H�T�̨y둔���,z���38�1�����w̌�yԼT5)a���^�_��'5��{e�4x�5�;*�T���mn�q���q4<_��b�vR���R[�.BcY�RV��i�r:�gY��쭃��9�K�C����`�1���U������3}L����jGt;k�ߞC�oR[3D�w9������y<k�-� �V�^c�ѐ-|q�Y2�{�l�GG�&�ɸxj.���oJ���S��V�Ȳ} /� �-�=?+Q&��$��ŏ��@�rdZ���x��Q�<�C�"��(^���{����1��ݺ�M�=0���z<�m�;�GϝH�*M�$_�9���S�t���˰ӕ��*�6pH��Q��k��;�vq�N�;0]���3����w/^h�
� ��I��ֽ+��W�GwiGڸ�����u%��c��8���
���Ͻ���<8Ut�@IB�-Z��ý�{mi��m����˘J਺q�V��Qꅻ��{��nM�}w���̆�xL=���p��
,.�UM���̴j��p�4]�&I��-/�9�dFW�/y��(C(�8<"���- ��S���{쓨�*M| -ȶ�i%?�؟V���7BLz\L���s�lT/"w-�ELq}��ݾf�Y��M^�� K� uk�~�	P�C��ZD�]	=�U����ƤH���x�A��k�t�VU���M�op+Ə�h�]�2NK���0`����~��ZLT�q��RY���7�Mj�\��Б�Ƴ1Whw������Jy���<�U́>}>Ȗ[1��Hŝz{�W ��܅�k@D��`?I��ϲ���_���9��~���
.��R("Iߧ�"�<=�x��A0����}��ʶ�*j�
�;{M����;;��(cϏF�G�R5_�Z�l�f�������	v~�#/�m���w��S�%}�g�F�ZQJ�R!��x��>�K�y�A��Ƿ�
\��c��f5ݨI�� 7uC�����*���%r
���ba���`���1mT7-�ws����}<�A���^���D6f~�6�Rl�-������JO:�~	{��)��>6i,��<d-����$e��U�� ��n[������(
�B��*���%|��:�!D���]�(�u�!���5So�����t�^~�y�a՚h���zF���[�"�᫭i���{��2$(g�����T��b�s؋L��/���_2�_7隯��4/�H@��.}�HWL��t%��.�NP��M�x�Wl���*L��GdO�ʡ�����`#8Ӷ2	�v��<�� ��=G�8�1��G��ԛ6���Ihhre�W��.���b��qQ��c(�.{��N����F'�KL�UG"�L���&:]�H�DH��̪��ĥ�qǕ,ʸ��ɸSC���n��\�/{�w�<�zf`Idg�(�dI)����!).��{�Q"��ҁ�D�k���0�ܷ����:�NZ��}�bWw��6��)����M;.+��c��n�4mH������*��]��/:r�N�(�Q��K,�v����4(w�9*��HQ�����؋ҁ����=�s}�4�}�����<\��cL�_�08؈K�]@{T�~Q_{,k󼜖9#r�%VD����}[��C͎+.w4�U�"�$���I^���ƾ޸���D�d��|���e��ZAj�n��,�������$�眫�e@�������`�3��$���Pla>/:�z
z�3�j�a���lg�k\90[8�khg�6���i@��<�w� u)�YQ�sl4;d,��D�b�ZQ�C�G�_�k��4����tI<�beTA��g2řx`'�@������]����Թls0t8%X�8��>Q��%�}%��V9ٜ�~#�^������d���麛�L}L�zڈ"�u*�)����`����cv����+��'#�/8%E���Mf��>�����9>�<�M�u	R'��E�f��\�W�K)4k�POF���� @{/HdB��dD�P9"P/�
%��L=�x3
�)γ��~�B��\�܀�b�CJ��v�� ��q���=��Ks���ť:qݝ[<#�6��k��y�$����"'�4���"6V�lO����d����*'�r+��';���,�.��lF� K�<3[�g��֙ϧ�P���\�-��T����,�!��ZU�`qOǝFD�Db���_����A��	�ڽ���
��p�DH�`is�i׿�x�D���Xj^*i�܃c|�x������hgR���P����u��e~Sڦ�a���L��}.u�SKȝz�g��3I��K�:��T��$�ǁ�n�6�����|�L��������NP��K;%2���Il�S���T�����M��S������o���,��
0�Ƥo=�w��[\e*��+5j�}8j!�3G��B%�zn�}�-��ü=����4f���9q�������?Y�i�캥1�uv�J�Q~��y�~�}�)/
nװ��sE�C�=j����5�^�G�|���>ϒ$��1y����x-�##�Ot������Ty��[�Z.0MZ���S�:��E��S�$���r�]aD\}�n���g���sg�%���+�/�sne�pΉ�?�F������N�ؖi�}�6 �˞��ncϳ-��H3�U�B�.�vD�ƕ3pp,���5���9�T�Ku�ޝ;�����^Vӧ)���v���\�T1������o>��9�O%�i���1� ���b FCP!�82 �� �@�=6w}����f��Q���<.���8������ +X�z_��=��T<��5�dm����Q��]�d�����z{���"ǹ�(W�l��H��:e�s9m�S�i�y@��_&i��s3n�2{YL�Ӕ�ߗ�h{�?��Lw)�vj5�.S��Vt8��0�  g�U\��k摰�@��r�+����X�P�}�Ȯk��c�����+@`�z��/BI����Y�W�~�ܼ��y9{�z���)d]�e�Ŋ�~�m|��;��S�1���Þ9�0a�22O��f��;��׆1�!O��=D<;�J�{Sec�+�n�.�[�Lz��f]�o_=�R�����(��ܫxB������y�|A0j�q��:�L�����zk�y,�U6粷����,?|܃�*|��se��|fv��;�N��1��0�K�̮����O_�|��*4!��'L����A�	���I��U� yM��Hr񳭲'�^��?T�-�v�;����� +�
&�%�'`��o�d]uJ�(�Kٔ�x���]r�5b*�NND�Ҥ��`�ïE��
�/[�Ĝ�V�~��i}$��oYk2����fvvQ5��8���U欴

	R.Ӊ�xJ7���4�cE̥�L���݂�i��Z��
��%u�3�,U��7Y�PwR�5���:�h�j�H�K�<�@���(��Tg�ݡ$�kz���:j��~�)�!��) 81��0F��@ѝ�& �D� �JR�ݟ�����w+�5d��n+��u
��'�+|C$�+������mqi_���Q�F��[��9<�b�pȐ&E5Pl�6u ��P�*F��"���BO\��S���4�U�^w<�=�|�#l����B���4GN'&ix�*�D�@Z�g0!�p��pM⵼S�[���cȪ,U�@�I��b. �T�����$���d_�2o~��������o��,�[��u�	��[����s{]���6|�ZY#3�w������H���f��A�*��\���@7r�?yo�q~}=r��ï]Q�=1d3��3��Ϻ�!�0wZB�٠�Mj�2�p��P�vEz��+_���s�������^P�p�����05["�GwR%p���x�%	ڧ�Q_zpη�-�->��~/����x�y[�nlc���J��#Up���u���0$YA$��}��JHy�`��^����Q��2R�<��z\,ҟ�9���ٔI�i.��$�������\R5����2����L��{�2�N�B��k�f����_�<���u7u��.V��`{��1��nkER���Yy��u������$��Z�|�t�B����#ŦE�D7�ݽٔ;	���zq'l�8�x�=�*��Z:�B�o���uf�7��˩����l=�80�� �B�F�Rp` ��)@�U�T�Px�� 4��!�3~o���z����<}���@�H!�Aܗ�0���� ?[�\y@����4��)�6��N�~���\�Có�a�:g<�z(W����S퉄���t��5��<�rS��󡃝������
�]��<ơ�����Q�P��Y@��a?s�a�
��2��l%�;��SՇvIV����)C�R<�ޚk��;>��l��I��쩶�`_���~z�n%V�1f��!�v&ϊ8ˁz����OfmU�;o,.3��e�w�p��-��<��u�����ٵSb�����z�i�,ك!�N�M�KNz��<'2H1�}v��_���4� J�`��*fg�k���t�BNo7�"�`j�s�L�d�`�lb�Cٹ�􏾛�o>�dP4~���T�%��^���E�J��B|��,)��o�1O��7y�"����u���[����ꛢ]|��^P���%�n�����i�V���}{�9��3K_wH��:���iMc�bSϹ��sc����m���V��V@ ��FpK���i	&Vf�YQe�t0��,����kV놺�]]
ս�.�%�ȭEm�Ẽ�j���Z�M ��i�����k���vf�G�³�*p+���7��w�p���w�C;��*w\Ի��I�8ņ�ݼ�	�t�m&E��of��붻FU�q�l��p|\	�>K�,ԪÜ
Y�(��N�lV��2�;�]/�ᱮt/Ep�1.\(7*Ɗ{��[q����ݲ�ݸr�.��x=!��-�5RU���H����d1��)��'W>VL�/�����~T'w��ӽ��E�b�VU\A��]W%܋(��p��ݴ�a�GI��vN4�O5�G	��)C�)�Kᔹ§�㽶��X���K�ba{��ep��X2���EZj�ȖW�\�(d.��]�ݾ�Ϗ�KU��k��$�:��c���T��u���20^+���p'�~ڜp$�ړ;E�G�6��s5�VOM�`�f�2)�%;�=6��S
(>���n�n���K\���SǛ�%�i��kWK�J�O71���N�I������ղj�]mSU�չH>�����h����u�+�ɻG~\�|�c�}m�E�}�`y���P���t&���ݡS�N��P(EK�L�U�:�c��/���?ש~���`�k�qr�J� ����:�V�í�&����r�r��wh+�]���;/�I�T�td���E�dY@���;�"��%��4�53�L<��n�t��=+w�lӛ���6���&���s�,���� V�#w�8S��PijՕ�]�ѷ�Liv�X��UY�ci�9��~j�=#%.[�9sBӧBp��d��t�R5�{�ּ��3��ƩO8+MJ�-���}�h�j�b���s2��콡,�o���U�V�G�B
�ؠq�%rB�[/vcg�'�5.}Y��YX �D��gs���"���ěv���!��)�7�Z��v�t�k7�#�e[����.8>�]�5U�����o��$>zW�SV��޸WZ�eVƈ�r��f<���mU�2�%n���Y��0r�&�g-a��Hِ��hl]�0���[�X�Yy$�$�c��®��x�ys������)�l�����.��#xaSD��j��0�ˣy`R�Y��+t��/�ۛ�k^�~����&��d�9���L��{��w�Ơ}��������X�dN��z�����~q�EĞb�w�gn}wu��r��S�|���zߛ����8��}}f}}j�r��8���^:h�7�ɸQ���T������������q�}}f}�Jں�QUUL��Tw6Z�Oԅp�ǏO��>�>?q�G��g���>��{Er&���	�)��a�c�z�wr��*��ǧ�������8������?4�n\����PT8gXp���O:T��#�"�r������������8�>��>��\��Q5^� �������;��&D�E\�룑W9� �oOoo�>�>>?q��}�s��ߧُ�e\����9)�i�O\���J�6|#�E�r�PY�q��u�Q˟�**^��AG>��)*��.]:p�\�CL(�;���"G)��@P�($�t!�Aw���{Y���������F.��ј������K�K��:<�΅-���8Ϊ�d�����Oj� �"#� )82"C
�$80+��{�zDz�JQA��o���}��|����gԸ�͐�+ߨ��O��Q���X��۞�yY[z!G�߇v��_����"�[Ld��|v��M��b�fO�S�� jwC��e�0��Qu�1L8wEw�[��üA���MRD ��˥FW���w��{��ȇ��Q�x�/~F;��Q~a�X�.5Y'r5�\,TT�;�Be��R����6���/���eVzL{y��~��Z�>��P�>�G �"�n�B/Ax��B9�D�&���<���"��[+�j�<r�f׎pu���ix3���hM������ᷫ埃������W���*�|���*�;��1 �F萆�3��ߤ<�����!������\�\��n.N Xt<�������C��qC���c3&�����Ӵ��<zM�����J>s��V-bq0ܜ��'�)��t�w_;�9�Ő.�'�e�����ƨ1��S)�;��}03g�}�E�	gRrp4���z:QV�y��<�ù6�n��2K�Ǭ��X�=��U��:�
�G�����ba�1%����z����̴n}ςQq�a53j4�=�F�
�J�F�)6��c���s�fh#g�u'yj��{�9�_w�������u"<E��*�`�%(�S�(RB@��f���{����{���r�F��ɬ��O�
�\��ʒ�?6-B�~��PГB�z���}!aoܯ��'�pk�>�ؖ����ܴͷ��Az��5�U ��=Lz��/O�v�T�줚r�},L���W�c,l���7 Qg�[��)���^E?�.��>m��h�{�]�?7I��O�{�{ku���H��_�(�b��QڈM!�G�s�^{����k�h������iy�x�T{Y�V5��@ik���¡�6���oLd��q@��QVfಶ�kf잫�C�Z�
���G���z�%R9Rp�\@µ_->�_O���V��Śϼ��}�\�9nN�@Q#u�-��jM� �06a��4�H�R@x�U�ř �]�\�B��~v�r��SZ0�C�S�N���!��20V�{��5y����F�s����B^G:j�.���4�@��;�r$�}lc} a����0��[&��:���W^g[u��8�!l���؉^>��zj��Y��Eكe���4��jMx��Ì��=y��Fn4w=�zf�z
&��fH0N�h�nM��p���͚]����FO��ʟ3+,=Ét�V�����4z
�M��D�W����Pat�zl��yU��;Un޺����+��A���o)��ls�"չ�m"�g�+��}�{�iz���[Ab��N����JO<>w������k�w���������L�nT�^�%C��A82'%H�80� iU������Oǿ���]3��i���<����JF�=&J�!,|�Z"<�9�E	00��*�\��Jo�#D!m�Ҥ�>���8�6c�Q ��c�U	�ܾ9�ߕ��������Om�� $DD0�`C,ϏB/�য়����ѽZDڎ�W\:fD�{�J���MYߧ�{ճr�E)�͆��y������4(A��0���a�L{�m���L&'T�n=Rl��/���Uxs��r�M8�Z�Pw��3֥4;������	P`��حf���f5�,�ڔO�];�H{�<�^�1ۓ�C��Ȧ'�;:r��ơ��7.���Ȕ[z�P��]/��?D<7s�����|��O��.m�~>���� T�Q-�pYSϳ�����#7=�p�W޻_G{�ң���t(n�=*+T(2h��D�w!孄ځ�95��Տ���:{N���,�ܻ"���N>]������f}RJ�Q ��1�G��9��%7l��K+&2�>���[pƯ?�By��*bǇ��bG����b��D��a� ��?")�q��_^�n��9{��nBiM�_+S�k�F~s'n:��0�{-��[��;�Y ;֯R�D���F�w�I�Ѿ�+f�*��0թ}st�4�%����I��&�d��;�a'��t�{7�vU�l���"�@� B�4	���pe;	T��'P�AN@�(�{�~���u]ts�|��ޘn]�@��7��oq��=;Cｖ(45&!�#\��N�\����Ǆ!�I�<0�����9�!�׼�i�~5����?B�&\c���b��,�8��ӻ���$>`-���s	�?G�X�Ƌ�4�1����N0�e�~�W�;/A�K+˻�3#��R{���*���l�5	�qf�S��{�PS�ض큦_�h<���Ӝ�>v>��ӱ�Vs˄M\4q�c+|���Vp(�
?�}n3���uJ����υ��b�A�m���;oM�:��<_u�s�}D0�?/���u��/m���{a�+�8�l�wU����ك�ܵ�'Ǧ�c7�AxwR��Q�x���nJ3�+�Lz>�u�@�V>^���߽F���;>"⥳���1��9�(�@!��-�Tc	��\���0���\�(�����fy~|��Q~*,R��Yv�H~�l��Q��p�w^n�-��&v��W)n�p�&���332��`��Sa���e7~�����H�D{�*�����ܴqW�%`t���]����7�л�p���k_B���7��ξX��O.�IՎ5V��b(��+n�:�0#�f�T07��f�a;{�rN�
=��(�Ւ7#�u��-ov�m�Od��o}W�LU���B1 
���2���N���@#!&�(apld�2�oJn�x�Sgг,Y���������Er���+>����R�|�IQ�7����ZL��aU�B��2	�c�~����>�o&�>�dN"~� �1gѐ������������=ߤ��o:�S<(���ĒL����-�0���`��G��|��(W}��Yă8pW���V��e׳:�7�ɖz2ُ�
��.�q���C�[��ҟt�]�%8��025�}/�>�ߗ����Ze)0q"|X�=���p5�v�t�y�z2������MԌ������L8�x���%���p~a�T���c"����?����Q��aZ�td��G??=y�p�a;�N��6���%<=�Z���)�``�a��k�4�{(KF�2�r�/�e��RPw|��8�AHԆ�{�f�49�XZ	Q
;�|�L��-l�磚��v6ң��yI�fy�>����{�H�F�戮F�0)��~h�}�o̐N�W���#3�#�֟�۝�J�4tb��K�xs��,wH����U+חt�-��&��د�5k(�3v�H?u,��u��6�� n��F�����U�����x���$��Hl�1�n�P�'��;�{Z�{8�:��ζr,QN�<u�N�Ť����շ�4PrV
s��U��q�0����0�G�4��P�P!�J�pd@P<@�NJ?z���>���DN��?�P�|����LN��R,�7g_Xx��%����ڈΙ��{�LM��~�Pr��1���\#5�}�_}�U4��qd��呫��O�ѝ�0�<�Y/7;���aӴ�UR)�xX�g�迖l��F)*��!r��������r1��>�ݣ�������1�{k�z�����)�ɂ�H�wy�_\�� �20�h}!o��FYc��.G����=��"{��E���l�8v�g�����A��|�Y�?�a_FzB��{R`�Icc�8'ޞ {2���H:�]�"�<�u�ͼ���՝#���������'��	�m���U���0`�)�5�_������<!��U<��#yIfi��q�Z�`�<��6T���!KAsn��y��=3��s�n�cxZ�3L�\R���u,V�1��N���s�1�!�E������{>�<㊁�=�&�^�Xz���n�պ'z��/X�Ԕg�{�i��J���XP�G�����ZY�9n�4�j=�.ۮ�d=��WZ]_c������?��ސ�^�Z������YS�4���祉J��Y���T��$�W���LF�#3�B�]��G8���]�˓���������D%�!��Ͽ�� �a��oh�J��6A�݃��1����YC��Qm7P�׎qY6&�Xl�ȟ�̻���<���W�a���Z&vĄfM�3��
 &	���C�������F�X#M�rõ�7�u�R��z/��OD�\����r��A�ml���\����U+��m�iڢ:ڈc޵ kSZ1M��}��;�ޓ?c�He`����`5�L��gӵ
󴇊���5�^S��ӆ%�:9���1���C�"����j���u�����Ԣ�P���
?T�h�����<���-��E��+1cTIsm��V��ǜ��{e�;���f���fl��;?i$���	b�����ZO�ט��4pL�����cej�z	a?S_q�9��29�0�}��6Ϙ@�qgr���>Jc7����!C��ٳ�����l���5�����5=G\�������U�����	+nS32�cg{D�	�h<2{��m�ɱq��t�8��z�P�~^�N�aPz�y8X_���[.��R_��>T��B���N��N��S?o\��N��T\g�WkcaV������ͽ�<a��k��M��ؒ�ߖ�SVj�s��_C�2�7~�c��w�[�9����(Q��Nˎ�G�^#���|#T��A�e�*�zf�]�o��iR홨�w{t�j��i7>�;�v��]�����j�^�e��b9�qd����>��ה�wO{���rww�ϟ<ߙ��~W�)�@�@��h�tg��Fq�;A<��ݳ�ew��r��a�zN�=C��AqP��W�r�)�K��8a
��=��}��:
�J�m�x�A1�W� ?}�f�//%�їp�iy;Gh`��զw!;L�9������c�	�q�-S�����l+�w�9*�k��L�@����^Mo�/.�_ZSf��~�e09�{gX
��&�ϓeP��U#t4��a@����`���~�E�S�L��ăg,}�a9�3��*�S�_���L�c����s�l����;��t�:B�k���u�݌�fiὊ`5�c6�"�{!ت�bb�����ݍc���O}E���� ˼N�'f�u�@��}D�|�*3*�k��>g�fZ��J�
��z������n�U�n8��n�-ie%���t�Yc���6/m�:ŲI����'>n���d�:�1�=�;�rWq�\WBa��mV�}>�i�y��� ����r�aK~�,.�RE�h�������ǩ���% �� �L����ҤZ��&c�L�!��K��aO�y�������0�����ަ�y�,im������a7���ˏ����[ux�]n�6�e[���̾�{2L�&14��-��Oz��/����ɍ��I�ě�ݸsub�D0JǗݏ.�����&��<1���h��Ċ����A #���5��2#�3�&q�;lI�& /�����c���� � ��ጐ,���6�����O�H�2ݘ]���������
;5nB���^{ɀ�����V~��'ē�Q��+��shj��5PZg7���-���������{ RSbؘ�����,ա�
Yꆑ���>���&�vL�ڢ�Q�?	�_�~���P�U1�#i(��ވ�0��4�=0���Z4U)5��%��zooOӞ[-������?�s��؍ ��b�!zf5\;?�����N��`ƧmdE�'�0���ə�I�Cp����u�G�hg���^��\�2�#1��C��T⹣���*���Ў�g���O�T�kk�3���s~���3�G�_Q�]�O�i�Ԥ�{�#r5�b��fe.6S7̹����8�sM�!��󭃏Y0��yn/�(��*j�XkHY��s�
+J�������f����|�T��w0�p�����H�zq�^���Y[X�k��~�Ͼ��� ��Q'*Xi�H|E�ky5q�E�0�����]u�暱�fT�S�KD��s�>���;̵�?��#b�u޿�dt�fu4[�,vmǫIVj� �0A J��:@�^�ZGT]��Q��G8@cT��T��W[7a�Q��˓7��%�n���"���nO��m���� � �a0 !��FvE��Ho�
l���OBҸ�V��m�o��5�*(�㫡��Xx$E.qPw��n-h�%\�{En���'S������.��"_�uf�c8�z��P$/\jyM�:���r��*!q6J��0�R�fR*C4�1B9k�*O�;��}���223�����9`Wz���:#����oK�D��&����nݤ��gx8�L�n�C�_[����N�\���H��ui�[��L��37>_gMZ������-O���r&(���^^�2~VF�Uk�f��q$M�E�#s��> 	0"UN}��}/.��1��� O�	�z��q��Q=4�Bu�z���.�[��)��fefo���?
aB�7�^�/ʆ��
�7d<�YF��Y�h���.��7��o�R�6���:�߆�'�VF���d��<�#z�:��)��&ÿ�|�vu��^�  (�(E�������>�DHx;���5�}�^D��!�;�3
i��RݤvLޛ5�Y�l�ĵH�Ⱦ�4���H˖�lr�uN7��]xU_v\�� � @&{7��f����}���n�e��Sk��&1A���!Wq��`]`8������-<���㊳�յ�[Z���z�-k�\��q:��s�\uƵV�0��^�. N�=_
�n���X�b�Ӊ�9�{ǱX�-�q��q��d.�V�u�����ZuX�^�]N�4��i��b�f��2�	8b	���e\�
]#��7�%	�S���r���xn�w�ɋ/�S�k9���Q�δ0�d�j���MN}S�Tvw:��;
Ok\Y�J������Y�T,2�R��6cW�!'�㝼���œ�;�.�՝�sL���ʲ�B:��i�C��؏fc3�M�[Xԗ�Vv���Gُ�vI:V۪<)3k)Ь�C�{�Pq�p���^[�A�{���~��S��Vyͬ~�E�5Ve�sq6��,:Yf�S
<������FD\��u#���%g#�$�� U&�q����uL�Y@�I��F��Wk�\��^,�����)v��o9wᖦڇ�U6���ھ	H,����LI�6;ˮ`�=M\�y\�>J�.�Ve�L�9dstWu��.M.���S�mT��kR�P�0Y�V@��=fX���pk41��J�t��Q#�R2�Ȃ��0��ƛ����)*wI4z����,Mm���]�N��XF�dԪ��$P�%���0n)����]@��h������v^���.oq;�NEX�l�l���žPm�}+��g,��d=��� �bt�ZM�F�FZi�NA�Q� �|��|�EQ��Yq������'>a>q��A�1/R�����)e�-c��[���]0�Nɕ���]�f�{�O���\���n�j��I�bXƯ�f9i�V5��e�d�|yַ��3VӢ/��E䁆B2�4C�Y��R/�Lq�ٵ��B�*��|����ΰ��}��^��\��CLT��#:��K�ݻm��S:�q�].�r�u�;WLh�����)*�M=M�=8�i���tF�p�ÛXq��1�\����I�������5y�c��[��w���0s�EWY���v^�!��b�Z�J��L����fm�i�1�>�2�j��h�K�j���\U���MF��3�f�IP�B9��3!�GI�c֣
����� �0�֎�bݒ5�&L���a3d�-I$Wao�+7/_'m�*�ݞ�޳CF�ӮTh�B��c�D�2��yG��}����P���GX��#k/��x�;�frg#��sG1rW9��n�ޭ��w#X�g���V֬ݕ�7H�f��_,YЭ�ݺj�^ɌK+���K���+�(����u3��$۲x|�_)0nv)�d�����{��V�,Y���X��>&b�x�����S=Uw.t�2@�/z`��К?i��
���4��s]Y3�ov�F`*RJL�HSi�4EԦ�h��B�d�h;,0XUF�QRlR��pZ�*�,$�ST[�q�(Ti���(�D��͕��L"C�1�w�t#P����k�(�9Ҡ���$ѹ	�4�M��!_t�.�)�\xn�W �5U YN�A�hܦe��R��A*�Ca��L�&��Y�[E��iȗ����<#ધ�e��nG������9�"���7����ǧ���������>���o�����/$���B����'54E$QRU7�������������>���ϯ���fQI��P�
AW>�A㻑L�����NL���5���q������:>��>���0r��Uª)�Nx�t��3����������㏯����q�}}f}}_b(�/c�ESR�DE+f��fJ��!A�#���>�_�8�>��;��Q~ЌE2�P��dʢ�]�Oo��C�_#,'�}|=8��������q�G��g���ih�(�=�%O9�EA��2rYG��U˽$���TU�H�"��/����(��u�O��T�imVU�;'ȑ�UJ���\��Õ��)��T^oie�RT|M�ey� �Z��%Ws��*�A'�;��2���I��A�U��#s.�\�v�Y�u�!׎�	G����]�ᓷi��CL�fѣ/�Nn�7H�!�M#ɺ��$|x��ѯ?-�u^y]υ�E^%]� ���,2�E�0�C	�T�E2�<z���y/O��%��	{�&�F�RdJ�5]~c���mP�<��c���!�>��S,��a9Y0��:�2�y*Mu����q�p�	�#�k����I:!�26�	��ouQ||�4;���f�y�n����k����V}z�Ǡ�z�NҶ�Q��\��d2�](5X�GG��;+,v]���(�ns�kK�O���E��.}�U��W�?z��	�+6�Or��vn���������|���C�F���~(�7VǾ`Y��P�M��"��ڄf�Tn�)݂(o�8Z�c7�%�ԶK[ϥ��(q�g�)�e�Z������0�f�R��	�q��/��?T?���	23:@����ʸ�J�@�1��{q�����(���|OQ��|>D�nL�f<�_��Rp��f~�y����x8��ӝ�Beg��/5(��~�PwtE��^O2�� 4x�$���p~\ �y�>y�����}xVv��eك��$�t1�s���� s��c��bF+��H�Q4Ώ�/_�6�W�ă���(o��)J��e�U�����S܀�N6��cRa��Pv�����^U�`����C��e�N�e<��JM8� 2����h�L�f:�ӋBY8��j�4O1['T�M��F�o:��:���@�A�2�2i#;N�@#���[���?_�s5�3ＫW�m�f4!��O��G %�.-Vp$|�F�D���	(�I�[���§[;	a@E���``�Z,����E]�bӳQn�f�k[�9+� ��y�J��<�M8�N%��F�C�gĀ�>t����f�M�^��ʱ��!D:hJ�|�׽"�ȣ-�LU0��:3h�� ������z��ެ���rg�&��>��]��@�{�r�Bnޢ�|П��Ԡn�*/���'�>ͿN���0W;\��c�9>�wU��gl;@�h��hrf�#�{#�����>�~^J��wfs����a)i�	3%����>ő��}ڽ���_V7�.��s��A��t�>=��>���\� �oe�KN�(��ż���*m˿4�.�|����S�XF[_{뫶���{�ُvP�g�k� ��3�f.N�Go�ခ^q�\&�U��Ǡ`َ�6c��;��mg�WC��?hգ"#���o~����Ʉ4�\�H;�������z��iVy����������+(��#����-�pBG����g��z���M!沯�/�T��&�b{�F����9wU��jq�ӆ��_7�b�z��3)
��yC�^��f�F\�wBp:��ܪ=:���o���[-��@�d%B2d�!ɐ(�	�1�_��?~����}�×��8�8	8[�[��~�����驰h���Ҙ;���]|{+1N��f��/�c�:gX㸗��'ua � m���ƣ�\�5����v!X[c;�-!��\��3p&�864ȳDw�h�� ����=ON��A���Ro侅O�Gg�Y/������~\Xt����̌i���V���g�����cT8(�PLK��ݣ�R�oĎs���<ĉ�Rْ�D(ߣ�M�I�+��4}�:��F�y�8y�!P�� 3#^Ry�#�|~FR��	�������bgӄ#g��J����f��b�-�!�[7*k�(��Q�jZ�9�����>��0��sY�!��H_.�q*�6���������*w;B��<J���ܜx��!����FC�/��/��>W��F�����"J��|��f�\��G�������>:��{�R���0U�~+�/0���v���A���'���?L��dH���,c�:�9��
-�9�-���������?���g5���?K�g�ͱ�hrъN��i}�6q�@���o3�t#����Z�NH�C�>Q�W$vfwg��7��h��vg!'nv�yy}��ij���,�Κ�L� {s��(wS�.ޗޏ�)��2��&H����}y�<������ ��b�����;�N8蘶�|a/\ύ�����
�Ѻ�<X,U
^��RϪ}K��:U=n�x�Q�bI�֜�lh.�.��G���$�-�Kv����ک�qR�s&�l��Rk��� ̹OFxo�=��I�Ԇ�����&)����^T�?}?���#ͨ+a�*4�n7Ue"�����SuxwO؅�D��ED�Yg�cL��X�����î}���93\6����x�2�M�2���j�^�e�2'XJ�Sޯ�#�9���hHQ���������Mu.%�oqd;��r�1��8ex�o=�6'�uQ��So��ѡ�Ʊ�����4��ϗ��sn�k��xK�#S�-�]���C��%V36)ĳ	N��/c��s�Ts�������Ć�	�?�p��@��粿!m³������w絔�Y/���g���Q��4�Qu��l"?ԣG��ת�K���w�,�K���6E���[�GCw��Ͷ)e���1OL`j%�0���aY�z>�k���� �/��
���y�W���v�h�Y��,PT��E����m6Q��5���x�=���5�&LPN7��׋Az��)�(ʢId���M��^���rL����-�Sp̼ٝ�1j�	�X�8��Fj:�Ѿ9�w�úoK���Sp� �Q�!6�E�S"�L�n�ʒQe���A�C�d��#!��L������.��Y��29K+��*S�dH���о��r��za�9�YDkS\�%1+���%���ߚlo���������Bk���|��v�j^�6M�N�vo)ٖ2��^�n�LT�k��S��x��Eiw)0�\��%ץ�

�8����)�U�y�������lU��G�uuf����[�>r�2+af|��1ri�n�
��Œī/��}�ޱ}� 3��?><��oij�k��N Z�wh��@@ZL������C^'i���Gn�2Ls����~�]��]?c����K�8�u�=K�_:�u��b����{���wL���W-/��Vj1�կl8-�NEY�<��}K�&�R�|�YTX�Ϫ)ȁ��	�����ݯ`n���>Q���7����K����9j����o�bTh�����_�Y�(��8O��d.��$bg��C ˨�,�e.S�,˘U��Oӯ|���O{T7�D�Ǘ'�z��L5��w�=n��s��.^���N�A|}�l�Z�-"�d�~���}�:,)��22~�2��~��Nu��uA3��X߮yp�ǹ�����L��vXL��6��\��Yq�R��.�Lc���]��r	}�{�&i�8�Q�#�w���VNY�k�V�����o���'�fa������TDAj�(��s����LB�z��~�k�Q�ޙ*3�_c��Qf�'���7՟}]�L����[|�6�nީ�nO^���s�3�>�y�#}UD�V$ܣT���Ԫ�b�Ǟ�v^}ij/�A����2�un,?}��kj�63�s����d1�ڧ��K��#��$(�H�≵�^���Eg��	�T��N��`�~N̛�n��P쁲�ٞG6������ԾT/r&ړT�B���x�u� �z�ז�;	�x{mX2@qU�Zg�1���E���|j^�)29��OKN���^�%b�;4�@��£�g�1<�,pռ�	�.�l���^:g�L�5^�y_�����ꆁ3�[�����Ԅ�${������mϕ�D���.�أ]%�0A<�������C�;��ᬶ6���G����2���
���ƙ�����a'�UG�|]�������|�����km�x��u�ϲ}�խ������ �~�SQ�+3#��ki���v��d3Ml����ԺDZ���
�K����F�۵��s���+�����5�ll�]���s�;0������6,n���-k�F��.l�YԊ�e��v:�wL����|��?|���+���5�̱���d �=ǟoҾ�������A^���1n�j��:�����SH�Kz]�ͮ7����q�;���ͽ�w-s��v��Z)0\�@p����#��+��d�i5h�Ƕ�ؼ;i�]{��a�(�;b��A��"X�`Ѣ��uK��\������o���dGJ��ٓ�<��i}I��H�|��~3���1�o���5?��-�~!>?oٔ��ʺ�j��ltN"�k�$����T	}t���Rd�`�dW��H��ly�Ԟ9%�_����Žu�9+/;Xg���;T�� T<j�N�u��(���&�Z{�K.*�����c\~���7��K#/жD�as�;��p��*֯QS�ޅ�B�1��� 	s����-�3�`�������_N�ٙ��qp��#L�.�
�W�ÌC{���J�,�k��
�B��TMq�#C��:v��=G'�����>_X�d��R�܂ ��ܔ�W�t��#y�=�^�W���iKx�d�����B�,��*���/� �n�F�Z5h�#3���i|.��$��V�fv�3�euA5s�+-؟�t��XJ>�@�轸�v�˄U�Vi�K�ø�+:l��Kஆ��;�e�A�����v��|@���&�_q^�]�,�{�c�&�8���R%�Q���h�����"HAC`�7�5�IZxt�����ٸu\��z�s���2�>@d�;�0�Eﯩۼ���K{��v�-B;ۍ�03b�_�q�1�6Н��rQ�1����󁾗4�{��
��Ղ�'�ja.��	!s �G�GѶ�E7�����VɆ�;k�'}@Kjz�96�d܂��a�8mcC�D�ȕ���e�cRQ��n�>25�S[&�r�n�lA�s\]�7*vc����&8�C��c53v��ȶv�>�e��2��ji"�|����v�z�̠Áڂwǫ��}�}Ӹ���{�e>�Wj`�AL��UV���u�^���(d�����ӭ���=�2¼3�_��zV���14�/\�������tS�c������[>E�>m?}}�����(��n��TaKC��/��{����10�F����+Ea/���#��j:��#N}�Z�(鳧�%���
�3�s��x��;�.�J�ތń� zS�TC��T+F|���Y�_����5 a��јڍ�G��Ӝ�����~4ܐֽ��-ff�5S�V4J[�ogs�����{2v��[�w�y(�/��o�|Y�S�
�F]-	fq	5�ŝ������k�ܿ������L�Ơ�r͔�%����^*{ZM����gJ�fk��RE]l���c�T�7MW� �R�,�%9(�mÖ`�$Ȕ`9���n<��>����J3
�j!M!����|x5�D���Tf�L�O^��sB6Kz_{�^������:x2�P]���I�P�j�w�3�� ��cW��8&����}���[��ϡ[ٟB1��^���[t~*W_iEy��Fy�2
 R��y��1h�9�~VD�]�W��cB��(���^��EN]��1�e�$�<�����RL�!���i
������A�~�Ѩ�Vg�����	�^���}��KЇ��mE�$�ٲ�m(�!k�
ui�M#�<��z/��4+չ�}��������b�C���XRx�$8Q&x��{�-���C���Q�??8����$���*&S?}�����x�d�}��	���b���������t���A%������@�4��G`"���)��3@�M�@���z=��Z�D��5�t�{�>ߴK;N̦&P��{�-�F 	Z�J�L%D4��b�cケ��P�aq�,i�f[*1b��V�l/��ɽ)\�����=��8%�����I|����o�üD�7��g3��l>��[��
t^b^�`놢�-Ү��r�v�"2��Ú!���Q�ݫLi̶Dd�[)��y���u��݊�a˧�Erok�+m,�b�|[�r|�6H[��{�Oᔢ�(v	�/����F� �%(��B����}��g�_��)����cTKj@���m�����z�L0zh���r d�f�{e�x����gS�n�9�-����?�*<c�g>5'W�xoMyl [�zD2N)cG�v��2�F�^v��E�����7k�#{,�E��J���~��\�>����:����l)>��G0{ڑ5ֺ���g��}����P�o�'f3�4W���_�=8�ޞ~S�z�<����������B/���`��Ǽ�~_n	=Y��{�M�.1�k�Y�ST�<�[�]L��z^��,}��7P�A!�����$���W��FG��_oK����H͖ݶ�x$,�(�}ֻ�N="-Mc��`��Ǹ"{V���G�_<"c�!���%�c=���g����de�7�\�n��*FI�d3��S�Ǧ��1���MI=,�j�N�_��F_�Mw�����V!�/�����W�C��g�bA#�rt�b=M����(S�ބh��/���L����?M�?}{1&�3�H��ᐶ�D���?y�q ��[^������s�}���ݼ�h�guL`B���c���1s��fa�K�R��`�{c�B��1v���وnIwn���P6��ض��*��5���T��і�c-�ΰؼ��J.v���N��i�A˳$j-m�t*�O������P>9��hM�,�J�EG�BM���b���ܳ��v�MP{�|��͞���ߊ2��1�J��d�Ԭ�J�E�O�S���a,�17��_6J�$0�`�p���9w/����%�|��Uu��.����S�)��6'L��K۵�C¶L[����Y5�&\'I��B'*!s$}��n�Vz]a��uN]�^��meH:_X5��K%��7�s5.yr��J�����\e�2��KK�FV�5N������4��^��J�7t��w:u�Te$���e�Al��;saj��ݾ�E*	� ��{���w�+ݸ�����x�n���Lx�����Q��� -��>y/�9�2�oVŧN�&3�A=qg%P�Z�9��6�-s�&�J�8���D���ܸ�����y��z&���n�u�`������mq�B]:4���2��z�$�$��h]�Q�\$�SN�7}�Av�A�¨|	>�����d����q�I�we
�D��z�I��E��W���{7\Q"I��d^MՙH�Ijٔ�w�tj��_Uc'�Q�Z����uD.^)��;D,�hXb�a�/�<%K���h�(��r@>����k��KkTR7)���U��*':�כٯ3��E�Bl�AL��e!"��9�3l`�ղ�H���`�'U˯R~�x�"��]x�zd�o\X}����!�Om��T,t�Z�A��8�"7y����&�"lb�9Y�׃���ꪹ9A �#����f�k��s����t��;F��9��ݙM�1m��:����	Z���㎴�OG��^�p�s�O&ܱ\N��7"0�,�*�o�T�{I�9��OP�Z~vx�8������{1�|��������N
;9%e�7�׽���[Օ�bh�o�
j��;%���#�v�k�!����$�L��-Y=z��	��_+��ǔ�٪��z��<��7Z��{�!m*ǋE��Ҵc��/Y�0u��]�h�9�7&*ۏ�٢�D����&�L��Q�,�7g[���L�Kg��3�MP�b�woL��;좯+)(.0c�Xq�9�,CI�:���ѥΒ[}����iȖ��۔�p�e����pmw'p�����Cm�q`��p�7����try��q�x,�*�1�)�����gU�bYp��?pȾ�AOQ{�.�B��#�)eL��+u�"/Ãǧ��㯏����}_W;�����.�"�D��^ܚ(�(�����4r�8QO��������||||~8�������o���U�z�h���:��J��EP�N�
*�AֽOO���������>���ϯ���n@}�>	=�G
\������e�H�F����A�(/_������������G_Y�_}��)��
�~!"+�2�X�ʦU"����&�\=>>>��>>>?q�}}f~��=�����&�O!L��H}dJ5�*�\N$�U�*�~���������㏣�}�w��Dw�fS���ߩ8T}�Ͻ�קּ�.���q�HE\��(��Q�P���"	SDE�D!T�QKA�/I.vQWoL�$�����>Au˅��~y.\�(�.�"���bq�9]��2C���T��lr�j� )���.څ0���2��E73���7I뵼D�A"? � �� �� Ԟ=�yH�|��I�(<F�~
��Dӊ�$e��0��2S4��k�����z�px�[ɔ�|6qZ�X�E�<kťz�5��}"��&��Eu��WE��m�w��r���s��z>遦�T2�;�C;�NR���:�R�b�u�]H^�`1�B�:��]��{	c�煆�<�0�@��O��彩^7�> N�P�^4~�.r�G���mvqV�#5O�{pw����$��
�'�^�
�ǄMy˅�{W��]"���{��^��c�M��G��sÉȻ��Pn,/.=�<M�0Y�Ƶ*�k�ff����4s��#C�Er����R]�^MJ�5�Թx3�N�]�D��V	RA��di�]B�����}�JP���L�n���"8�pXr�T���/-����lj���}>Ϙ��I�����]������eK�,+t�����s�ba��N}�=hl5�����ˠ�f>>/t}�3�%R�4˴n��B�lކf,Xŧث1�o04��*7Q:�f�:���ukqe4Fb�x��,U��6I��;n�m&�u��#hc@ѽhm=��dެf��FF�JJ���y�==����o.���C{{��q��8N��O�{��s�F�"I���3H�G8^�ܜ;D����AH������fo0��(���S�9�==#)B�x[�-��S��*-�Rv����ŵ��}��=��7���!�,~oe�0�y�K
��W�05a>mx���i�=_h��ULi��^���ҋ�a�|Mo�0w�\����:��Ň�*�K65M��|���l��g)�\ ̖X�S�4��wn�+;;�E����i�a;��3b��"E�$L�+�1R�b���u������k\ˍ���r��MA��}8�Վ�,�8�OH����P��qMl�D��y3*�k�f�,qj�?�J6�L�
�`��w��J����C9��d2�.�z��g�貆s$�l�I�q�=0���3��mܩim#$�qE�9�L]J���z~�?�����qQ��D�k����*;�Ep��|���f��Ͳ���wVk��|�a�����yjF���_��~��w�4X�j]H�N��UƱiXL���"�o�O�We
O\���y����M��Y����������(�Y�קl���X,R� B�5<#vݻ�We�t7L�3M�])I��n�]��\5����-�{���̹��H�?�Wf�yU��#|vu��F^��0��j�1�g,�&ny�A�zn����+W����}�"C�6V�ur˺赴�sj[���۲תVU�i�c�ۨ�f.s{��u�X�_1D�ڂT2���!�"C%��2d�t������ż��y�L��94P����0�D�QY��|~�� ��@�Y�Y��Ƕ?����y��躩!��X\J���g���^=�<n��e.�H��w�k.[K��&���,`����O^�� I�T�H��D�uC�:jƶ���ej��<�:��j
��g������^\!����@M��o�D���SWS�����:y�s�.|�4�|�GH��t�qB�=��-x��ӭ���R�g����q���U*�q����<�g���3	<47>Ao_t
ˍ���Hk��[LO8qX��v#ȍ��횃���+??�G����Ltc69�q��04����Pݭ�?�����>���G�/���CJ�2_����1����T��)���jKE����A�<c�����u'B�Eb���@e�Se�'\�)l�gyu���S�lC�1p�wZ=t猍��t���z]�{���~��Ζ��u��0F�n�bcw-l$��Λz��x���E�իe���~	��O}ƶ"�ˈׄ���q���ɾ�{-�Q��2��.RϺ����԰��$>����]����s����˷7Y7t���R�{��Ċ�v�,�7�9`yʏ*K;0/߄ �Co|���}�V�9F�_��3�E)�&���ʌI�ffѵ1G��/M�h�N��3��]�K$>�z�2����ӈ7��9w����a,g&{8q��cw"$etM[:�c����l3}�O/v�p��g���B����Z����y!u�z����qD��;;�%�9GtV���҇(n-��ܳM�]Wzj�Õ^�;���֛h���ͮ1bF��v{ ��ul�
2g��s{{�j�.I����5͵CZLK��;�$�C54;�3�8wvw����ؿ@�b����a=��c2B]w��_e�v����M����u�|�n�Ӱn��������5ۓEq�f���}驪)�Z�;�Z��M=�پ���Q]�1�^�V������<�^����^��|���;�������Cz�_�d�ڷ"��a��ͯ�7hѣ/�o����KۧCjɝ1���΁"fgm�5et0�Ѷ�2��>~W�m�˜���'mU<����]�L��J�_+NO$�|B���s�'S�25��S�e�	�v��N��u����BHB�B CA0��_{�������r
1M���7�dt�^&=����w}�4�����wJ(A�7��w���T�F��Twӻ�^�?G�g�D@��O59�҉<��΢�ߒ�X���^y^���W����j7}z���ٝ��G[�$S0j�ɫ1,��x��fk0�|G]os�=����Z���f��*d��MzS|<�t���|�ë�W�K������`�M�%�dT��f-��m^������5��ې�꧹R �Ey�3���(f{���+*���z�ԓ�-[��u6�]�c����U��������b6�J��5�9kw�>Y��,�Z���v<
����N�\�_��V꨽��r��9�r���+�Ƕh�nb�f>�~̃�hNwMr��W��,[q^c�>�Q�u�D<�ݓ�Gy�4v�� 홮�T���7K�"x�g��T���������ACcAb�]�s��1'�Ɔ�~�|�	x��'_���X���u٨�G�a��;�d��Y��Q�1p0��e�J�wk��U�t�+�x5�D����τ�@E�!� ���Y�=x����5���uD�P��*'&�c��h��ё��v�ضOf)��*�zz3�.)/^�kߤFT��χδ�GG�;=b.#�r��`cUԉ쵦m)/.Y�ܲ��!C#O��X�ߢ���U���vx�h�aQ}7�y���`8P,��ZT3�����b��=`����F;��5y���#�|�q�So:�h�@�ݜ^�J��=p�TQ���{��B[QM�'��s-�r3-�%��I�;ڡ䴇ve���V�9��+mR%Czd^-&xtE1n޽�K� q��akǝ���R@��Q��q�W����+��$�5m�9MQ��w����,-m3+Fتc�9�R��R�v�[/X�y��r�w�ؼN*��x�J��� ���m��ӳjɒ���i����d�{��o^���'u�P�Z>'��_���2�I�*5�f�GzpY�9����=C��
{���WgUtX��n�OW.�Q�IU��)��3+���m:��#��4�˗�>�\�)��y�R��R�w���!t��,Ί+# �\��E.{�{/���|��M�5p���y�x)�ށ��<�<B����d�DB"=�������ߪ�Hm��%f���)���f����1�+���c:���[��<MMEF5�5�]�&Y�&=��
�g�`V�����v��U�S>�i��OG,˾;�Zm��<=���ԋZ� S�ۧqZw�{g�Jŗ���8��<�;����Iq��x�2ں����a�Z��"v<�yLe�F�9��bv�E�-p{���Ro]��u߹��E���ulf���R#�y�{��Q0�f��J�%q%w�������b�7۹#�R�����]x=����0��+ ������-\�2M0�-!��M=��:��㥸;���̃Y;S�^�(��rk�_��u�IcF�WM�n�}�n��lT�)�����S�-�r��}��rl�u�z�z[��-dwkU�ش�+?�:uO�狍��Y��k��N���<|�?��/g����̺���r�LEY�t8�u�����t�T~�,�e���V��׽��V*k�&�0���VJ���m�w����>�xx>��HL	ջ��֋�7ZY�; B�.;��m�؍+�:�kʸ��tV�sn-�nR��(�f�j���D��{;��o�I�_���1��і|9K����S����<��-�A'�Pn��0!��7e������4���l���ڥ䗜T��Uo���JC$31��q��h'����+5�oHk)�F�k�+�^tY��π*n3�eG��{o�	����XܥPwCl:��r�T�k�܈0c�C!=YPå�uF> �J�YL����g�c�����kIYg|�%Bٟ���~m@ah
*�wLR�|ܗt+�O0��}i�;3}��"m� I�.C2D��11�-���Ρ�\����H�s�S@3�� q5u����gp�m�So�r�n�S���p�5��sd���ow+�jn�m��j䘋��1O��8g�Ӕ�6��oe{25q��]=�Փ�����FXO�������~�8�zZ�F	�a��ҋ�<df�ov�q"��}U��?Y�o�}��\s%}#��s�!��`�{�t��Y[�Q�� �uh�U`�y9輹5�n�Q��WAnI@~�t�ٲS����ܲ.U��fW�T�sJYElL�~;}�6V%Kt��l!����;�/߀�D��"�8m9(�N��<���x������j���Ǘb�Lᛑ|�l})�S�g���3%gN�s�CU�se���`Twz����{�
5��ofEG+�.fD�7���l�[|�8½^�"�'.��N�Z���8�$7�1�_��r_��~ㆿ<Zs�[�q����R}�)�bA��b�"��l���V^IH!�A��W����ܘ�&L�4ћ>qQ�x���̘תgA��M[ou� ��Պ��ё��`|^|�`���PdP���mv!�����F���*F��z�Y�w���mOs�p��$�ť5�S$�##\4z/Q\�*�(���դ��L��ɕ	i�@볾\Fv���֛<L�G����a��:��1�n��Ė�V�5�_s?�mnxOv�{��#���d=�0�S[ʷ{//��L
��~~<��́��]^�P�8+��K���ç��ʎ�|�" t�QD� �0L+ʜ�γ���çs7�҄���B쌾��k3�܁��^�@s�0�WmMK����B���#�����A"��}���{����'#�����0��vk�B��n/ԓ���TL߂u8��o�|�of�O7(0=Z������[�x��v��.�� kpN[��P7��v ��/��s�Xh����@�|f���}Q��lgL^%�ۼo==���&�⻄=e����\Hn1u�~��AS3#�z{-������V �[�T�����nT:�c��z-� �ѱ�N'u��y�X�ڈ|��I�����jq����k�|�������3��w��:���lf���opEvx�yqD�J�������R��钚+�ϱ�p�5�NRb��Y�T�A�$�Wz����.�76����=������6�~�|f�_��X٪g��:����P+J�,�<�8e����9j�u�`�����ؠ8�4@u]rܖ(���Z<��xx���~_���:pi<?��B��e�w�n�ܣ��^\�G�����]�ÝҝO�o��y���&BX�����ot|�3B�:�mgw��Z�M0���WB�W���+y7�1ٲ����S�n�c.��i�=��˗Z����J콕�W�����[��|�/�r>�"�P�̙�=��ӵ-+0��:m@��L�a�89I�'-[���8WX��K�0����t�=���47��<=�qk��a��d8���+W�8T'���oF�Z��z���X΋y��]~;��J�u�&g-�Ί�%�0�Pk�n�5ݦ���Q�X���i������B�u��4��n1VP��o��xVt�:�Dk�m���F�_$I9���O��u��/�0K`���C��~�u;�����#���v�]�����9�Sb�o�\�@��ʁ��۬
�xM��˹|]��M���᫻xZT�ı��e���u��2�1�q,��Us���՛�ՁĹfэ�hw._&N�5Q�ok�m�髛ڥt�����*|BŷU�}&����c)��t!Zq�}ӂ�`y��kqi�Q�ʩ��ު'�S��^L��vU�����m[]N�[��##�5A�[pe��_��:�D��K��z��;氬��i�XPC�E�;T�������/L�Ȫ.V�����#�
)�E`������X��.����w�6QHY�IS�`�*��Z�ں��Kx��t�]�[r��V GM�
X����ŵp�,�]l܈

]�`|�]��E&�#��u��=0�L]�t䓈5%gAd
9�������N�K�9÷m�U�	L@�%�����F��.A�M����b=�b���H�i���E��~�?W>�[��M��K���*��
�N�ҍ�X���״hp�v��&=Q������N����6z���W0��ֽQ��[ᗄ71l�O"����D��n��';��ӏ�=���n�n¾@��U:^!Vj\�-�̾$N�	�#yʖ�����Kv�;�qP�(]\���P���V�p����;�i�&n��7�o��3s����T|��ܕ�"�fm��s���r�����ۗ���S��M�=��{�a���5�Ȩz�9�.o7�̜ɂv��.���|3�O��S���NsYY�7�ާO%����W��̤,N,"f�F�d�j�X�mU㭳�"��Ǚ��`�Ө�څ���W�N�f�������loZ��i��E�㊝�Ls��;��D|����ޢ�ʩ	iH���A�%Ɖ�L6�v��f�$*��"̡TR���l�%QH�H���~��-7M�[tj�D&E6�F���CL��J8Z��ۢc�EE�QtD�%���\�l�Q6�%'B�6J��.Tˆ\��l����F0̙h�i�������
��$;����L�Ӥ�{7�(���G�r�(���
��T�N�����߯�������㏣��3����9E_�9Q9'����S(>/w
����?�5�����������q�}}ft�=�9Ǒ���r�|�ʯF,����y<�s�'#�TZ�<z{q��������q�}}fw�i��8Ts�^��r�*9p�F��;w���p|x�On>�=�����}_Y���PW�6��͕�������"��>2�(�}ݬ�|q�Ƿ�������3��{<�e;(�S~��8HWg�wPk��{{q���������������q��H:NBED~ҭ)�8�t@U14�P�ǒw{�){���!��;(�(������;��&{9ƒ�(\�ɋ����w8=�*�ϦL�.�E\,�J�!5Nr�	�<y0�z��Cܽ�������qwyOwZ��cT+su���u��͞ä?�6tN��Pج��ÂÊ燈��I[�,�T�q1}���b� �zT�
e�]M���=�]�T�S�x^2p������匳Ҥ�[o�j�K�
T�CjfCZ�`��:��!����^�]t+<o�Yl:�ǝ�iayy$�[�Ԝd�+��[��}��S���#�!��k��N�Lýǽ�U��8w]a�g̤jm�{�5t�#&��v㽹ي�;`z��Z�^ܰ|���*� 2�s��P�zӦ�_P(�ϭ���g�9C����}BMEU{���C<iɍ��Y�\=履�0��7d�c���5����x��g���_�=�-�T^F�-S����u���?VP�)i�� c��	/X�{~�+���D;��w�)��}��=J��(�̚v�>zϨGm߈�1͍���SN3ܞ:[��c3,�:Z�ۭޅ�׉UGyT��쬙U���������vo9S���Z��:���0�O�ݟ���9�>(vޟ��<)�P�p�%��F��9�dHMc����X���Z��ʎ��(m;b5��!9��qDj����XCP���:С��kQ�ԇt��GW0l���|n�kS0���p2�Hc7x������t��?� �� �`y������Ԓ�~?�Y�,
�#�Gw������AV�`�+x�vx����m�l$��ϣndgI���gZ^t��׈]���&M��Y����5���M!��O��~x�h�o\��gvz��z���u%&�[㧫��vվy;�ck�r%g��f�[w�FZ�C[��o.�6�z#�m��U��A^�q���,��B|P�cG�c��/��R�}�����KpP�&u[�_9zv�7����-F\����鉝z.�;,�<�o�4n��]��9R���~�9O��j�ͧ%����6��M\u�92�_���"3}='k��꫃C������&V�x`��f��n'3Zv;y��z����&V�!�q[V_c+d�S�ƚ?��r��7s�3�*��y��STM}�U��Ǖ�3��B4�m�i��Zhsp�o[���{�z���)�G�z�|�,T�X8�YWٗ3ps(��-�7����P��y9v������X�h���ˁ;B���Z�wg
+m���ΰ{�X��mn�?���D"� ����ih�qx>��,���뛖��n"���u����Ū{�c���#�J�c�D5 �=�����N*%.�8�'�>�n�.��U^��ç�4�rگ��+Y�k�h�M�v�Lw������r:@)_P��㞵��,�چz!N��.]���!�\	���n���ў����S�R<E��ob���?���P`�`�*�������GB`�@��6y�z���0�
��E�P�ͯC��:۳�o�vS��z8i�f0�w�qٽ�� ��Oi��lȶ����YW�_�3�Ҋ��sSlz�͍�ݳ��"v�OTQ�m�������\��{O�msc{o{�q���zc!{J;�w�u�^J_���^v�����~O���*6��1����
��@B�U�������F��ŗ�����{�]�|zX7lo��{U1�PwY�s����'�zn}z�]�.�2�kmR�5��}�R�mW,�L�b��[(n���).a����2a�����JW�n�Xi;z�z���8�\GB����5y���M�7����3q<X��ǂS��DA"	��G���sqs:����T����ޫi9w�v��45^�<��űM�=1j��(���l�w���g���5Q���\�dq����5�PA.�{9zwx�!9���������1�ݲg�H�Djɐ���22�F�L%b��8��3L@����Ho�E����%~�
�}&�m���6x�\�[E�W��Q�nN�KӠf���OyxԝCZz�1|��j*�2�Ë��<W����F�}=�u����x9��âG#JV��ޱ7>MC��%�D�����Vq��U��f���l�:�+
��9��ٌ2M�IE$�5� X��/ٍ���'۫��Tv�C�\0sgg�&Yb�b�D�k*�N����
Xv�P�"W�+u��p�=r������z�a���7������<rGZ���7��k�C
������Xw��C�1��x��q7a߷�ۿz�mr.)��#�#̺,�+�$�G�s�<��;b��u7�;mgR�H�K��$�b��0�:UՌ6Gۛ&��L����w��׺G��z=�v�v�jo-9�j:a��6�yX�
��V�Kl�N|e�o9�<�
"�<���ˑl�%�
i�=�DB"?�bq#��~:5�`����K��S��s8�t�@:3<�~k���s��r��wX���uT���Zo��Y���ke����m�ك[Q�&�a����/rT��oٜ���}۠S��漱��;ve�Mk-�n|���^�f��5��/%_[z�a��Z��<�;�u�n��Y�Y���쎝��#X|��ܡ#�:�X[!�������L�e�Ciދ� �;�=�����f��4}�g��y�o��x(N�fc�{� c��9�U�K��`�E�f˭�z�},Q%�|���"��F���*3w�ޚٺ��MB9���{���O����4�E��)�j�OZ��3	��Q�}��}�3{�Sz���3�¦k�s3�����=�ȇwY,{$�f�o	tQ��ϓլ���}˕�"=�f��v�	��^�X�|/*43�S��w��íg�5Xj�J��U��W�^>��F.��Y����wg#y/���޵Ǔ��,�Ĳ���/0\���N����,�Ä��c�[P��.���΍OOKÌ���D" �����-�)��2۳����1�\��l�}��Q��^�\bu �f)����9Jr�}]�{dP�ל̉m�!�\���V��3o���e�J����վQۚޟW^%>��f�ӻ�r�WEoZ���X����mD�t]U�@Ep�I��v.������ܡ����f�!��]@~���O��o�>�g��a�c2AU����2u搼�y�k���_}��BT������������tz��N��mv\�}yc-�&���<���87ۧ�[t^����;���p����S�:���#eY~����F�T�7�������ed�*ϊ{�b{���g��tz�ː���`��ƻ ��&ש�z�ȿM,�^l	6���4齫�*a��0.���*�6��|y�4���V���#B�	��dÔ�4n�kk&��Rn����u>��F(o�ML>�L����|��"�79��C2�'#M���Ӹ����h�sVe��l\��Z;V�R��P���n���;���~ y�7�-���wkug�>z9��
�w�vV�N0H��L��f�r�-�z�ܙ��"�:6��|���?Y5ʨ�qZ��F�]���-lϋ�������%_^��2��J�=W'i��yE��E��]�n�]M���L�O4.��A�$8W���e��_�5�?}�e�k�c00/4��C.k+~�쮆+L�D4C��|����Mw�̝u�e۽�F�f�T׍)���j]��E��z�z�z9]���m��=sѨ������)u�nнc�bY��'f�3ۺ^��� `PE%����U4_�:��q� 	�O���ӫ��J���7?�������d�P���D��{����İng�i����
��E��ޣ!�㱴s{V�28cI�ע���P����l�p��҆,Pu����O�}}�m�>����{ZGT���Ҫ��o2%TS�;q2��G5k��<G���[p���I��]���uMxNy �i�G�V�����ȗ�:����-Y��Qi�[[#} ��8Ns�U�� ��>8�	��V֔�=���ѽ�6Ro�<#�0���iu��۱?P�p����\3Ҹ�h��ۃZ��}�y@�C����ͻqކp7tGMϪ�7��^��-=�چ���_�[W�:�-�pA���5tF����Ǝ}J)�U�!<�37�Pwo��z��Dޙ3����_� )U�Vs��V��@5o>�Kh�Lf6;�fWw�p;<׆��2��w&�h�C�Fx8����k���f��s�UϘ��e�&yK�9�qJ�}��cP��TwQ�[o�\5Y�M	]>��kα� ����Ʊ�2����<�6����+F�tF&�E�@o�*�!��;�M�8���������4�٭g��(X�)*ܻZ��̺j���s���h7z�F�{3�;0q�72h�X6��56�Jh��%����m �(�����q��/�B���
�j���=o�O�8�3&�q�*����i�oK^�W��	�#o���t��6��N��&�B��Y�M��nNϗ3f�<
/�k1��A��s#�u��o�'ȼ�p���3_��1�M.|.k}��wRnE���2_��L����q�����׷����_�w��E�:[�y!�(9T��'R�4̠mkM���~"	A����_���X��B(��f�L�~%��|f��q�i�R��{�9'�zjUy�^=�����ܜɖ�=w���Y����5Y�Z�Z$��c�pܔ���ƻ�bRۚ�]���������;�C�̩��3W=�Sf������^��\�E�q�/�x]|P��5����㦕�x�^P#�DVwz�S�-�-���\N���nf��9���Ԫ�Hj�
��0n�w���oU��H;�u���i�v�����T��qB�K�öL�`;N�ty�0�����4��Nm��VoJ��xSL�g�z;�с�bp�״���Kb�p�:������0�f�"a� �5�ټ{��ZBA%6��>�@�t�<���ތ0�=��y�zD�3�SN1�{����P��s��nڠ�}�Pq��H5�^!��	�����aDs�fk�v��0�"�w�j��K̄b�\UM�ۻX�DQ��@x�u�H����h2ǅ�4tV$�l:6�����jY�B�'���^�����{���v]Lt�[�X��,�Ewgvv�O�R�2n;n��ո�n�M�A)�F���ǡ��y���N�9O^����#��SW+�ݾH�������xP��ڑ7.{�I�昐۶��^|��\�����{x�I��^��OE���am�T�j����_1C��O�T����`K�0ھ�Gw����;j
N�_-�s���cl�e��Q5��ϼ��� ��� ��{�]�h���xk�*��)�vg9�c*�~7 �Y	�R{�fk�K��>'6��J��G��OUE���	��ݞʮ6����s�6c9�J�Ğ���z�E.MGP$����٧�Ly�c3�q����叒�!�3��j���N�Z��Ž�E�w��wN�2A335wun��}Q����"�\s�Ue����Pý��������^%����[<r�;ݵ��:���$��wF�<�3� .����q�.��Frbv�ːR,�~�U4`;��Emʻ3A�,��tqM��Z:��X�h9D�e�`�U����2UǤٸ^��`6�s�ӵ�d�ڴ2�ނ��Wp�$��^���u�����;&��"�"h��{��8��cw�f���}�f�\��s�$l���V*\��8�q�d���vmG�$2�2r���*�C|�V4���;�[��m�y�g<��5� �gy��͋>R��p�L��;o�X�5�1Ns9[�n�MU1�/Xc0��MV ������`�ӦA�gxynG��æ�q�O��ʴ���45C>��q�0-�2�속Z����i�٣HL�.�,7WJc���s%�NtW��;K�r�O�ne�.�I�F�=���7��v�����Ւ+�޺���'�yv�4���N�&�f�G��l|��7*���xI�.�K4�ss��U&;���ha�.�)�4_5���7�GQa��2�t��q���CE�Ќ!7z����a�w^��tP��]�ȥ�k�;O���Z��g�gq�S"��3Y�����N�K�kA��̑ⷽ��p�T�+D����ܺ)7!�e�#W��_���P!j�U��)�L�Y�J��fVJ=%#g�����"�-��MJnM��t�'Uw�kiNi3��I�s���[�����z�a���Z"�=��#M���;��ΊpVk��*M�}�~_	�{Ȕ}�KA�8��#���Re��f��	�y��1�$�5��.�	{�q�5g�����Ǽq��Gܙ����f�W�zԁ٢���i�g�2���g��)|��j��HT�tR��>+�KGwb��@k3�rW�����:!5��-a�0�,���m4iü�:M�W*���q�]v��Jf!�[��[�lߓݕ�NipY��́j�sI�]C8i��lWL[�����p]�8a��TPcd�DW
�Y��L�J]\U��
e@��R����H�%��Qt�)�y���B�]Ӌ�c��EAb���ϴ� �f�.������蘒�X�����W݃��۽��87m;��R1�l�v�M��{�-�Ws�(%NKL�R*�μ���'�]�K��7rwqǄ���+�X�V`�Q;�;P�y���B�7ڴ���B��N46�L����֘�2���ob�����]en !�z㾴ɦ��H���'��6��",|�)�\�׏��Uc�ԁ�����N]�}��FK��d/g;�]����P�cu^+f%�z��S����cF�[ۤ�0�qis�m�kN��m;�ъXl��/�A yӋ�r̳:ސ��j�#��|ZG��(ripҨC�L���pM��{��,zx�N?|{{{{u��������"q�(��
Ar�+��q�F���#���+��O�k;���c��������>��>��{�E�u�C�x���.�:AF���n��=$��#�֪~;��Y�o���oooo���������ryr0L�Đ�u���7�����x���NDѡ�E~�<zx�����������>��?>���TM��"m��#��fUj*U�h��5��kz޷��zݽ���G��g��Qs�p�s�0�H��t��r�ۯ8�������o����o7�����}}ft��{OW"���z�G�I��}��U��mR�zyzP�rdA�$�s��
wX�B
,�J�K�BjڢK1��#x����H��D����ZiS.����O%�u<�J3���.�3ä�$� �A(�zy��Y$q?�t�y#	�3�et�T�o����<g�מ��^~���; ��f�t�c�R�Z��rI���v:}���U�1�0^�}-�f�����w�M��_�����a�"BD`��|�;�����9�,����ߥw���p��q�B�xP�vhv���,{�kl��ҝ9��ǩ�$F��-�޸C�v:��O�U�8A��Z����+�tb�e��.A`5<�|P4��vq�݀�`=�a��M>�[�͉-۴ǣj=������L_FѶ�`���Lp{��څ�d��o�	XhUK����.K����z>? h���}�`�rn�����"�����&����`cկ�AE��yCk6>S\��*^n���0i���u�=�q-:���J�r�r��ϊɃ��w�[�"����y
|�=x�5���Leu�w?&�U��4���ǫ�^��s\��x4�c���x��iP+�edS����>��Cֵ⒈n��"{wX�\��x�^h��q�>��K��B��>۶���m���V=���.��eYy3��־�f��#�C��$��e��Җwy��]��=�Ш��q\fhDq��
y[��K���L�Ҵ��5�'e�I�W(򗵘�'+��,sa=\s�H�f����*��P�N��9�/~g��_��w��h ϟ}�n���o��XM뭏4*`���&���,RUt�Vv�H�mk�{�/��z�L3����<� =�]��{�&;kǌ���u;j��NYL�˿�Ov��i�Ina��aRA��黧��w�0��}�pS�x��Ǟq�9R*%�gd�l���8oQS�&��K[<���j͏�Z�w�hfny�ɩ��F9�¤
�i��X��}'�:^�<��4�/9�i�70�[��֪&w�?��ݙ����"�yu\zZ=�#K/T�n���f�g��=k/l�^�漙��nO������&+A8���aR�lk�������nEer����_O���o��d6V� T�eH�ƻ�����Xn�Ŗq�0Y��5\�������e��_z0�baR96* f	'��e�Ubn��e�|(�8$�//>�	�<��LߗK�.���N�U������_>֩V���8�OFG7/;Z{\M̃�f3\~��Yd�r�ɛ]��d�gw����<Rp��!��j��+�����r�3�sb�vt׫�TGZ��P=I�X�ܕuؖ��$�ܨ1��*�`����.��UwzA���I6�����	P�)(	�P�R�ʟ�DY7*˱��f��VV�`'	8q
�aq�?���a�Do�V�ly�L�>]3�"����� �a�U�=�;;;�Q<����
�-p*
����Łψ���%[3nVi��'y�r��T� /"��tzgԆ��[ ��A%�Ymkբ��tN�W��Vϥ�kƌvר<�Fr�\�>MV7�6�I�^ZC쥽���`���f��F���0y��Aּ� ����:�羣��s3M��ۙ&�x�F��۹�5���Ӛ(����,wz(�f7� ���B�����\������$��[��m����mZ����y�-]瑨������w�d.Vɶ�&�q6�S������*�Wl������yyj�d�-y���&��Gztπ ����^�'z������i��ݗ�y�'�v=h^m���$���P�Ûڍ�㘽ZQm���*�0���ړа�oI �Lq�s��[�/���
O�\O&�{���V[�q��צ���c�}���K;��_u��JJO"�q|�Z�57/k`k��\[����x�{-68{X3 �_N+ЉhD_���E���|7\��q_�#�Qu/��7y<�m��Ԩs����6t8�5��ϳX�Om!���[��R�M p���C�T
�����5�U�z�u�a��orc�l��k]"�JX\��Ӥ8�5Է�)�ϟ�w��X7W���v�;��
DX�������`nZ�e�E��Z�Y-�r�Mm��A�ځ�f������*�~���
p�����~���?^n_oJ��A2�Z��9����}S� B��3�Ț������U��f��ӖF�ɉZ��f��ȗ�>����[�}T�ӒӽYU��x�I�Wo�Ғήje]�O�q��ʶ�Z;��Jް��F,��Q ���s��Cy��pQFU�OsS��p�l�W��a}��z��g_�̪�$��T�y�H)"a�z�>Uu���ڗfd���)�{9_V��R5�`������*�1"o�Ł������x��w�V��f�����R�-�h�#�q��w����Yה��׷�n_NWbM� �7�+'�����<�d�"=���ՔJ�j���̓�b��C�4��M�'������,�����]���<����y_4B��i�mhW��K�P�ם�~�Ha���^[�+�(��9��0V��.oI�1����������wl� A��͉�}Y�Oό�G����|k�0�m���ޮ��я���ln��S���L��Z�g۱��;K\w-6[ I9��^)��0a�:�}�`��.��T?
s+3tTLoc#z�O��)���H���_ �v�zL��Qٚ%曏���_Y��v�ř��M�����_����<��r��"q���lg~�4'��=^g�ǲ�Dz����U|���M��ԇ<����OW��XV?h��5o\a�*:�t£Ӗ�@ۭ�x�/�ć}�h3&�	�w�U���B�T��«1��cxav�I�%�$��ZB��W�dӔu1��D�~��ε�j�>����el�����7�])���¦vnPwo�	����zX[�a��+R)�0��;@�O��`<eyߦ�Ϲ�^�����YOu��*�g
�FC<���y�<�u��2��ުdj|�5�����j�h��r��F��`g`���筘�h�w)��F�\���ۍ�j����8�+Y���%9�̕M��V�_�F��D��q�v����S������۶(���x����]�c��?���c$��=�T�e�ݢk�kv���wG��>�8�
�qf���p'R��;#9%� �1����+��.�)+^ _T�0���E��@}�@�ӝgee�e?gqgҜ^0�e�$�&;�6��\J�p���������I��Yp��Ö��"o<�x�;�>�] JL�z���G>p�>�Y��t8k��m���W�r3��+6�h�l1L�~���Hp��K�ky�P��0�ǫ}���_�;/�+2�2J�3�k�^�܇;M3�d+����:b/�s-�]ݖ7��Vl}�L�Zj���b���~�Z�4*�8j�?'l����k��orp��i�W��=��ޙ·\�u,�%�W���Fǜx�΍�\�ľ�0�%AYp�e�R�E62[���f�LW�n�(ƜH�H^�<�� @2&$�-�U~���v�h0�M����pmvW��,;�ˏ��Vr;t�T�G�H�|�9�+K��)��P�������gC���nỷ&�o]i�vv8�[2���]�Y�� [���ۗ�;���F��{�����B��Y5z���(W�����A�ۥ�����z��������6Cd�XfS����"�׵�ATJ�S���!�z�ֈ�;E����76ޔѸ�W�ۻ�����(�g7!e+O�H(�.ց:��=v�I)�1ɐ�=��X��zz�?����������+	�<I��z�Zw�F^�5��NBH�|q��h[^ r؜��1�)sڱ�t�UW�9Ŏ����ðL!8̬G�ޓYl(lкA�~�m�����1x^���F}?huQ������	�^��=Y`����WT�W���NeH`,�8�܎ǭ �¤�`�}I����]�Є�'&b&S7���A{G��'��.i�AR�3n�#ݒz]��������$۲��&l9��46����-���\�W��U��5����.o�S:6a�`ɼoc�Eғ����F�&ԝ��qG}����J���);��"b�����y��I:�)g�^طkw�6�P���5;˨t�vB����-����ߠw^l�_�:�9���裦6o��6������D�Sļ��>�2��r;��ݪ[�S��`C;�O���\g����rl�٫= �Q�hǁ��C�g_^؉s�枑����w' ���/_��9�����@췋�m�lV�Ȫ�t�1}&||�mk�&�^<}Q�6��4fy�҆S[���@��!r7�S�5�T���eɑ�������� $��,�W���½��27��OM��F��r`�=�7f&�5�9���qnKC޺�etŕb�U1�����8��qP�V�y�hiŝ��B��������dR�MX+ֳ�����x���b���7���;\'�r��n���K%�Yg����t���黻,+/4��Q�7CT���A"��dU���9�e.�t��5�� �\n�U�F�I���c��{T7'u��R���fՠ�:unᐗ�&	A"���g���N,_e�G0�c��ykQ�Z���D��h�*T��/�Q�
m��]�TA2�'��ǶC����Ҧ��	A�F�ڙf�ⲫ�	vFi�U,�����/�8��ѷ���:	lx�����{��Y��U����"��ʩ��_��V.l�b�r;&�1i*TF4����G���2B��ݖ1�}�n�.����d�MDx`<��tm�h/�H�]����d:�5a�z»�q'�qv�)�fU�W9lQb@ W�
y�����V�΃U��R�PL�]�*�wS��8�Q~=DK
ӡ��x����w�B�Boٳ�g����cb�բe����7}u��4f��t�|�py�U	���ޝ��/W�X�e�]�37/^��mf���F�S�^�W�`"���Q��*���Q�QwDВ�67pr�C��w�l������ɋ_�u�Y�c%��^��-Uط��!�-�{�jO{˾��r���Z�1�A�����W+Uf�7X}���9�T��+$_� 0"��ݝ��>�2|�r�wЙ�Oި�"�&>��9�:G �e�(,��������Ҍ
?�F���c�fX���`
�c؎���/5���7˾y�);�.e��K	�U��<B�X���4,ǳdղ��l[3wU\w]T�>j��t�:�6/ϒϐ׶~�)������~�U�$ɼ͡�8ΡoEf-�X5�^PCGz��K����9癏2�9�ث4��9TF�a�DoR;�/Xhx5чV����a�[�1�I�оp��[�
R��<�|�=X�b�_E*6�]s��S\�]sC�J6���r�JcH7d�7��n�вn{%�\(�z�8�>�Z$<�k���h�d�C�^L-$�[��G֢�}�����I᪴H���/���yZ�[ԉ����@��\�ޘ`DجUu��Ҽ�3͜�e,���Qf,���q"�\7c��F[Me@��wh�����eqѽ��I[Sx|vubͼ�s��dR��;'�e�ރur�L��Y�ήK��ff���.�a�6&��ս.mP�ݹ��-S��-��qY�v��^�����:F����u�4��,�F��z�S���m^��c�L���mDj��^�VN:�+�2�.U�oX����<�/�Ѿ�,�X7��sVRb��Y+�S5R�_2��^�FV�≲;ks'r��XqdG$�森���ձڨp�p]˦sx��j�m�O��7z��T#:u�}�Ė ]\���ə#N�U'QG�ɷ�k�9=CHhK%��a*�a�F�:�9Q]kWu�2��˺�\��k���хgc�6�܁��J�O��iG�.�mn Ԕ,���8�xfՎܷ����<��5��%ي�S�Яk�;��֞m��{9�>4D�[K4T�׆��*Q�'-Hn,wy�������8fwi0���q�5���ܻ��i�����L��	S���a�M/s��q0^'w\!<:.�:���Z���_1�4ZRH���7&��d�k�T�x�Iw�˹v���5wed�1�8E�n*��Jx��2�-RJR���o��]ܐ�A.�sFw+(^�C\�t�Q����ꩦ&�s�բY�J�[h���܆�S����T��O���� � 6+*�Y�ޒ,�����f�T1�\����3u�6�N��y2����c:��b֘��6��
S-T���>��h��Mrh���j0�k)������\��̦�Ka�zEgMeq��3a�[�����~ R�����q�o<���5�n�q�C!�-� &�e�>�f.��y6����hھ��ԦBMu�U��RU��$e�G9��dgd�6�n=��Й�#Y�-�b����G�	d�c�r]��v�C8{U�y���dV#�f�<Y7f�[��+��2�c���-fC���g��t6t�eq��2�e�]Ժ̠���Yw��a%r搯$ۏ�Օ�V��,h��Y}�V����j3��w���3ox��pU�R�\�p�,�eLU�i)չ��f;���/�_>Md�Y��D���5�0n�L]�TR�M�h�m�������lr{ֻ��*I]k,YZ�R�����>q�M��q�����}�U������`ޥS��
�Y��ח\��U֣�B�ԓ+���FM2{ ə���J »t�vd<����b[�F����2��]�N�츸Y����ℱ����^���Y�������2�K؊��������"�)�%������$�*�v�d���+�c`Pƥ�b���;�`����\�ڋ{0�;)�ŻS{y��D��u��*zu]�Xm"�Y�ת�%Zi�_f����j�C��iQ~R�;[�m'I6�`���^Cd��;��1B�A�q�(�g�y#M�ΟO'i&�9I�R�**��Tj��L���ٖ�ė:�:�P�dӣIeifB��Ց�;�ܖ��,&EESMŒ���40�In�TӠj��:	�BF����rԄ��e�|abPo4B+���z�_��\�8!<X�Y�����n��{�����_�����bOxs��\(xu	�V�qMUɮIJk���v���pH|ַky����z�n�ߏ��}}ft�}��u���p��3��|J�2iD������1;J�B~]�����{x���������}~���3��^T�����Ъ�V�S��bF�y���r�O�xp{���G��%V={x�������������ϯ�Ή��U�9%��3"�B�\#�q9W)(0D�P\�dL8q�qQ訨����z5�_Y����(��Pu��������ƑS���$S�V99�(
? ��8��U3�:�������������g_Y�7�'��"�E�D��5*�
$�dEwP��[�7'5�L�Ц\4)VY��O�rC�.�]'۞3�c�eú�I��F���q����ʨ���h��Bw��W.���ON�#�kǲ(��$�F��s���*eDD���"&S#8n^&�˒��EI�H6���˸���]�S]����'o�w�Wf�v/kv� ]\�1�Υ���\݃�u�>�k�'2�4�i�R�e�L9�A�ClK$.X��u�E�1�5�^]�%���:��&�{�V��β:���a�0"�Q~
b� W6�/��yؤ��2�:�/b2��ѧzI�.�(��4�������L1�^���%dU���U�6҃b's{�-���7Xw�X��m `�*K0L+A��(R1������I��q���^�y�9ZY�h���xޕn$W��.��ܔ������yC���@�H�Q1�[��y�*.1�1�ae���=��]+�0S����8�4�_`�m�f��5�˴�?�q�)�.�̇@tޭ�]�,S�r�q�C*��s�eϛ��L({{O��VSY���z�U{��ڃ���;97�[�{�RRۜrQ@����L{��z/����*���|2����:�y�i=sVoD�W���8:@�op=@J��^Ls�vE��������b��{�7Φ�_-�(b�L��zcX)v�Φ3]�ݐ28�D>A�	�TC18�1'f�]�^��gmK�--;�:��uĻM��u���ٔl��+�hvf�җi��'��4 Y۝�6����Ϯ!ɀ'��7��w����Dn�7L�j��;2��k����zj���v��UC���;��gO^fK�y]�KMwmh^4�o5Zsx�SuN��Fe��l��}-����ծשԡ�'o8��`oQ�f���f�)�}��{2%nԵǠb�e��l��=om�Go:�S�����wx��8-�o��(��3��Ñՠo��}j���~�M�Clpr:+�h���~��˵q<��x�����u4[k�Q$ٽl���R)��Z��X����]�Ȑ��]ݚN?rA��ї����5�6�mxF5;7�a�=Ƽ{�-}^�<��+I�QT����_ǽ -j� ���Ȉ*����k�&f���;��,���~���]v�|�qжT�'�p�<p}K��|.L�!���s[Vw\��_a�b��A�h^uND.�����c�]@����,��*�sj�zk#�2�[��W�7��̔�o�|m�q�N9L��s�{X�Ӹ�gr�Hfd�XH=�����z��
p�l�����_Ue���R�U^�$�1]��2�I��26�g��K�p!�����O{Ta��t����B�)@���x/M���D�/s&��e�N^E:���$o)X�	��z��2�z��6���$�9^��q���D��½F3v�/ �K�%g����Mí�4n��O���l�(=['���E��I�,̰��1;ݘ37oT�S��w�e�Ct����3u5�Ry�83KzLM@վ�'�n��s 1��C3�<`��^���N�H�)���j�%Z��n�,q��W;�m}�h�
�݊��'j������cH����yeX�C{�}����c��ouf�ݝ���|�=UK�[��������\���2LĻ:�Wi0��P�[.;7in�P�>��������9�;��ff�G�$���%�/A��lЩe����ةԻږ4�
�3L�������aG��飫-;� ��MrF�i'un�p�ي��%���bt���*-����G^L鴻�.Z9a���Xr���O���L����O��g6f"!��6g�{��J1G|���y���qR��dՓWC���_;{3Ǧ��8��޻߻~��{�C��k�`kۭ�1(�������s��ၗ,ͺ)c>h��g��`��Ȝy]���W�7�"L�\��_�Ny���mYO��f������F����x��g��_�}����l��;e9�Y��;���,B��ܣ����s��[�<��m �����s��UJ�'vm ��;�uAO�m��<���Y�ߔ���ߘ�ۑ��a���x�N�@u��Fa��m���g���i&`�s�n�0�����m�s�!��U`�hV,;̤nd�<��h�t�>�� <v�Fl��Q��O��S>����ꅐ����*��*iԊ�X؀G������B���ع5��R�ۋ�]L���9�k2�b�s��2ɣ�Os��Gp�䗫��@��Q����ZF��:;� K4̫�]�X6��[	�uL��!�r��iN��2�J�e5��,�"��ĺ�8�؜Mj郶뻺7�k�gZ�H���Gj�8j�m i�m"i�yL;F�Q�)bM,��|Q �"_q�����b�3���0}�~����������N������Ȫ�N8��d�<��xS�0�}K�b�M�!�����u�Ls�3��WD�.n��ǌ��g�]4&��[
�+;�󻚦�R�j��{"�-���m4W����+2'��Lz���3��Ny��f�Y74]]i��ﳴ��H	YԻ{��8��\�>�^w�{k�@�3�4<����fz��3�'���E�{����W*	�l��P�'��6-��N�t��ȣ��(f�:\^U�Q P�7����y(^/LcVO�ڷzom�Uu�x������؄�P�����wP�������ܭH>;&O���8��哴	%�)�Y(&c���g�{���?��?�٤S��}�s����aj���vY��nҐ|�8d���{{�b�Ƚ���Q�4�z��8%���Qyd:��kcs��;Gi4��P�s/�O�����y*쫄�%��Q��Iv����a�W��-/3��Z߭7�^>Jp�I�6��]�u������c<��w��GV��l��	�AlwDѼی��x �cS���q��wY���=f\[�v�������y��0��m��v�8aO���[#���^ד>�>|y�ㆽp�" �	�x�;K�R)N���v�ݞ�j��E��c�ƙ�B#T63�ŗ�{q��5y����f&�j�$,|M�م:�<R�zkk9����ѭv�3A�?G��6;��f.�o�o~�Sz6)�N�g5�׋Af�����:UML��ȟ��{�ب3W�!y�9�ו���y��-_����U[&Al'�Y���|���}k��^7d�k31|��R�ּ��4���"TD��kQ����ugom�jN/�0�C5x��z޺�Շn�M�Q[�Uk��w��F��POO�ve�x�5�|v�P��qq�`��'Jw|�=�>"9sy䖏a����]�و.��a�/7zYz`@V�$��Fׯ�8iq�^U����ಡ��j�k\�a�j��:�'�8��5#wy�Ne�2����n�r��G��mA��m��r=W�\�M���*o0��R��x����(���}�ʋ�o����Z��	a]��_�ڽ�bwm��T}�(��6z�o;�~�b@ٮSc����-�H��mL���c���No��Q�����{�����g���]1�գ6䬽���(��QT��86	n��7��֦j{v<�G+ǝVC��*C8�i.��[y6.��H���46n����s�jm(���XW4����[�75��ݚ����p�R3�i�k�B��_ON������ʝ�]�k��⨁]�����9��^��f�溟E��^�^3bd;�ֻg�s�{���EW���/<\0zz!4>p��:N'��!��d���v-�z�s�B^��۾���]Z�1��=f3�RA_y��d_%����0��V����l�߭�
����ì�8(���ds#�d�:��6���,[9��Y#9�_>y_�yQnH9�Z|��ܕj�ޅ�:\��!@W�l�|�n�i��j�=�����j`�ږ����m��6�:���:9�}�g��/O�� �D Dk�]Sd��,�̻;k����w$)nwMM���n�h�>Op�����^���û�M��{�tV/V���cҾ���Q=#��|z���ш;���-�d�߻4m&f	���}T}��{`�6}��>�Γ�۰��mCbzar���_��b���hx���
�����ts37U0k^g����i%	�ݹ,o���>�P8���5��kb(����͋f�x}�H��z���%^�%���5�e����M36G3^�ӏı�܀��"��=�,g�4���	"7�!}[���n�D�*�P�{;�՛�M)���*^%L��L�Ŭ妍��������Z���o���I�����~�Ҫ�̷���X�2b�k�t����ތ5�4�)�e��_x��d���Cv�1�j��.!����]˘o�uvYx���N�]��,+T�܈Ur�U���1͓9�٥���>ʤpA1Ő��D&z�(�i�H���Y${f�x@�jZ}�k�T�1�`(nٝ!����L(
�ľ������,�y�{�2��a����ku@�l��4MԪ�#�t���
.Cs;;3|L��l�)�V�5��������e�t���%�b�s4->�Qϳ�Yq�7Dhm`Ѿ���z�Y��A�3��*���<9ak�c)�JT@GY�vA����0���I�R��FCX�p���sGr���@�Z��4&��AT';���yv�虞ޭ���;�=���W��5VR�W��k4�w}KՁ�k�U���b��g6��ww>be7TҘ] �7���5c����32�u��������q�۵�v5]����4�Ǳd���A�DC^k
g8y^��D�wa*�mWONi�>P&}4�����f<z�6[�����zp�+m!�{���6c��Tz�#z�_=�����X)ޜ#Ֆ#�mu�J|���ܿ���oGY��.�ݜ]`H[>g�y>w��R��jjn*�U����!l����F\�/Hm�t45��_�I,k���;�h<Y^��TkSy�n�Ϧ�\�_vtV+�o�3���H�[D=��=v)u��Lpc��:4�aNI��N��@_����5�kR�߆�C���S�{4���a[=��`���7a�EO3{���A��p%�~��z�#UG��&ffi0������Z/}0%��樽��p6��;��+8ºc%�6�W^ۙ�k=#s���ޫ�%�G��8tzv� ��2�J/����5��3��"ɬca�g�?�:я,��j\��j��+{BqŽ� �%��C<
���%7Z �R{�^�hf�Z`Q�6�]6)���DCkH�n��|�4g��r7d��&�z��
�����N�������c�F�u���-���*|�gg�ȭ�r�6>P�û�e��@�� �E�{x_��y�E��x�ݕ��jc��9�,���}Z=3^�wTY.n�gY�R�y��z^O�3�\�Y}Q�8
:�g�q転�`����}"������&r�U�Oё�t�К�Vs�F\�� dR�A#o:��̠���|W+��'{@���y�.��Ww7��K-�=�sf��^6h�lQ�=K������|�+z�=��RSR
�ι[ӯ),yq����s+��)�B{�Af�N&��T����{ҳK�y�L��	w{C���cJznQ�����+��ģ�}D�L����lZ�w"Lk��"�1$�=����j�Ô�k�[�T+��Ε��C2;6I�{ӷT��&�Į#�+d��=,< ]�]��W9�f7�(.��;�Z�#o"�!b�}�
ާ��38~�u!s�_=o�nj�y/�i�v��i����Y�H��/:Yz���rq8�U-�K
�¢�z�#�k̆�C����(Oj���8�=%�\�,�j�绩,k�����}ɬ�������f��-K*W]�5��T�iv�к;�V�q��^��׃�E0�ڃ!�
��|ճ²��6 �6oYD�p�#����(�$���ʺ�k���۠��KgQW7+0"m��{h֡*�J���kH*Xyϧ=�Q�O,C9p-l���W�%�^�wV�ȹ��0�*u�P!��j�c�T)��b^�7pbݫ�n��Z�Itt��*$CoM5���=2������z���	ug�<{)X�Enܻ�eu$�:�t����jB6�ƍw�a�
C�&�T�obm���
���q-FR܊�+��v�ƚ�U�ʻ�ec��3��$"�U�^��V;��Sj+�A�`*���]��_xoy�,�w��Q�l�q��['#��C����9+%{8��9[&��Kf���J#��u�x,M(SAצ��fl�**�K*مb�h�ܹ��@ԧ����tu�8�ń�Er{dc�Qh�f�����k0��C�.*�lr���Y9���f�]�{x[\�}�&CorP�_��B�T�F�?���z�k��.���?L�!�ګ<���3��,X�J��Hl����ٗF-�I�*K����^۱���H��°���F�z�ܹ�����[p�Yo���=W���iW57+����X�wa1L��p[[��X�;k����S��Ʋ�*ЏG�W\�Q�.gu
����`��D{4�0��fc��/2�xu�����a7�E�]u:vIԫ:�j���:��<ߵ7��c5��LЮN�����=����ћ���K��r�'a��r�����s[�y�g^%��\������������v��m�u��1�s\�	V$	u>�����݇��_[j�:a��Ûϸ��з�k���1��,��'�L�9�'�i ��$E���\(zO�I�-^�C�Ğ%[N�	�ү�s�������|޷��oo��~�}]=�ns�W(�y��ȅ�"�e�VIAQD����E�	�|�A�.2***;{}}g��G��OH��*���DB��n������@�"�	�a�K@��\8��������������w��҅�E$Y$UQQ�����:��Ԉ�J ���hUQU�aI���=>�8�������}f~�����^�#�!y��z�'(�TjPS(4Owp�E>3��?7kv��{q����������>�M+�yɮ���*���S����d�!_�
�$���r��$������$�L��5��ED����EEED��s�w�}���GSA0�Y&PU
i��		Y��"�*k����5�.il����v�z{�,�"̞ӄQQy�MF�q:-	+�=�������*�M5x��S\C��Y���Թ�$G�h>]��K������`�TV@;��!T�����ySzw�����<���,�#(�޹ˏ_b�"�À�a9u�l-�Ǡ1�Ux���T����gvw��ԡ��x���3�:����z�{�97�)��z�oz��{�}J�v<U� ����Z����/]��y��|�{��ٷ���٣��]�i=or �̪+�ϲ�B�Na~6�����%�>����`�����o8��YPo�4�k���3xz��ϩ�"�FG��պ�����]ݽ��$�㭫waN]�o�n%"MC3 B@����g�	�?;�}�͊~��Ǯb��P'gg�`���R�%�39�lEW{z:NNm���� ��mS�3���1���D�W��h�p�G2t�rtk���Y,p���v��"�����Fa��+��{5Ig��I>[CK˚$j#��ݽ��V�0�6ׅp�{�N)���Fm,q@�"�,��5�*��:��?v}�����O�Di2 Z�B�Y�li�#�C�Jú��|�w2��[F}Й�ʛo��|��2H�Ʒ�����m~k~����i����J��Y��hM�l
=�s�Z{I}������_�>�'��+���d
��ǐ��֋o���Q���]Щ^�˩Äͽt�Ġ�@� B�U�%΢��ʕ-E�n����<طM[^-|���<�Sca�T�a��`X^��ۓ���wX�us�}���u������a�֭�дy�+󱿷��,ꢢN�r�`�T�^���ؽ��Τ���N;$Ug�A���{5�g�Ye�-�v�^�K�������u�~��NyB>��5����l.��P-�{�f�p��|ԝz;�=���,*�z"^7�P�`�����ʠ�m�e������SUs[��/&�:����ђ���;�T �{�O�绦���`v묥�5����y��mM��1u�Q�H�v_�n��zZ)e�|�������o�#,���>4q[�������4CP�a]�hv�p
�ھ`��[�4(���u��2�w�j7�$�M�N��@a&���5�|]�#aK�[��=R=������z���['Z�a�ü1���L	�p�����
�56/�ݿ�>z~0/����>��Z�,����͚�8���Z�.�ۺd���������#v�MV���d�δ�q��tk�g_�'lWL�c�s�&t�9׊�97���l��7c�͢J�1�ε�pwdȭ3UE��aF�Un���R�}D�N(�
��!V��P�3�W����-�(��a I��?���n�ސ7�Vwwn�q<�i�/a ��z��y����Uzޘ�B@TF�>��w\�@�S��xT�v7���:0ᾕ~�6����=��WW�|�����K�n#N,��Y��:��d,�:��Қ+�c\Z��[^��0m�d�ɸ܂�i��ꧮ����;��>��E)=�JA6��7����y?o���Q�u2}�������X!s���N���Q����٤5���s:2��?�H�v�w�*��1���q�ij�9h�@��kݧ�z.cFq@o���>�����fg	ȝXV�і*z�1�1�[���g����-�;��hv��-R��s�s.��T�4���\t|�9CWzhϏ�\��~�B�:l�7n���'յ����#R6�B�2:q�T����l��bɲ���7*�\� ���ˣg��h�L&ݗZ7]sG�U��us-��v�
�2'(���P_LW�	�W/W��#[�����f���*�L�+�ʚ����谽[6NW Ϥ��1��UnV��xx5W�J�u��EQ�f�B�{�� {�j��@t
�A��Iޞ]i��ۍpV�����S����=`\Hbä7��]~�#Y�<5gT����ͧF��)�;���Υ�ʑ����,��O1���K�ŝ�=l��vN�Y�����G���`K�k�<�PV����Қ}M��Ȗݫ�&�jz'��zNa�P�^F^����5�e^�=#�ޯG�=��Õʧ_Նdguȫ��A�R���J���������UJ��D���svq��c����2��=y��,=�wQ���ݬ�M�s"ru�w��M����pP����^�F�ؘF�\g����W�a	��ƞ�v�'=�H��#�qN��Q���{{&�n�y�j;���?D�C��M�����C4#�(�A��-7c>�-�t�j��t�rb{!�����H��ܘZ�.<o���]mW�#+��}��҇xՇ��LT $Q�B.r}o�q �".\�PjQ\(�%��?|$FJ�~��o{�V�7����E�d2`QNZ��^��K��Ce�-܈��}=e=�`��@=�{���~�TǢ�)��F
�}\D�0m<���y��n�zg:8�0��܇����=ǻ�XUU��������t��Q
G]�u����`*���Z����C?�\4q^�W��o7�&<�ĸ��}����hr���X9��u��L��w���mU�C�ތjn�t����N~8yKF�ɖ�&S|]�}�ҽ�����wMM�u�{/7��[N$Q����h�tܮЉ��hBc�h⮸��ŗ�����-;�q>X�ʚE�E�7�{3���v�*��E�,b<_���U�^Hqz�&���������?G0�޸��5�*`q���r�׋���Sv��+�B���A����jۗ�FE�k��~�*���è顯���@��0x�h��K{Ȣ�d�� ����$/w˞̣�[KMU�C6+�xu�L���X��1Yxs��^��p\��y���b�hy�7ny�-�"��q8�� q��
0��q���]zd�>8�Z.ޑzg!�K���ٓ��zk�&]�a�X|jg*�;ky']�7���0x0�Bֵ����?i�j���A��w�'Լk�8rꌊ���}��2�T5�s���!л�Ҥ9���aݭ��V�S>4||��v����rcc�ݾ}�͘�%	"d+�Eס�H��0���^ߕLYR�����4��׫�o�Mb��\���wE�������a�>h��Տ!���9{�	��A?NKYk���֜�?`�n*�Ͼ�sOQ�a[_��<��U.�"�<�Ծ��lx3�N��e���"�7s�)��׃G{e�l.����ѽi�7�d�E&=V�'�|��F!�z�?�?h���m~���U�[�
#;�;�}���1��E�R�'iE�w���9z��Ebұx�S�WT�۬����]<��s��`Ӊ��	Ϳ\Y�Z�f1����jY^ȫ�q���n��M�FC}��%��zt6k�0����m�}���(su9e��nMY��%۩X����y4�ǩc1ͽ 0%�V��FH@�1Pp�KH� 
 ��dlL�X�	��ʜW�7����{�<�������4=7�����!�A��mA?��9,tz�G��cp�K�<Sz��Nq��R���h/CI���2cHb��sL�m+b����;�V��w�>�'�����e�M�~َ�����缲o}B ��r�F�yn�w\�ꍜ�I�T��K��W����6|�->1 	��Q9�C�ꏝvI��_��޾;��]�?���)������}@GG��!��ʍCd܍�R�%����^���Vq�E��N-%�}>w�d�!����kq۵���A��i���c�ez�?�i�u�xݶ��;�l�g��4 �⏵u����}�Z��P�=>�:��6Ĵ��ݒ	��e�#���yrݞR+q-�g�=�m�T�ދ��~�m�UQ��6�޹�h��p��2*�c��o������$M�N}���\bϩef4Ĺ9�3KvY�D�9b���_�I��W\��j2�2�����t�7f�hMM�i�� �$��e78�C�(�����>K}���t���z���������u����N�	
Y�ᗃ7D��T�6�n���}�,}�Y敕�o���Ӄ|�)ݳ�W��K���u�Wf��e[d��Dt]��kW|ݳǺ�D�ǝ� �ev-�}��à��8Cp�w1"�s��Zo�v�|�쾿O(f�:�1�LgFڪ]x�{��nE3���-[���W�yy�n�ZTI��pGL�l���Z�`��eTû�5�����j�d��|�v{�;:��ᾃQ�2=�ӽxY��uvu�V� !T�oT�]7�>�n_v���s��b�M����M�*k�� 0hf�+~U>���#`\m�%n����UPZE�^?th�ѧvq�� �}r`���`�R+Wr|�<r/WcP�vgz�F����W��@�T�A�	�t��D����?y��M̊.0Ld�2v�{�۽���5�`�K"�4S�c7�����;��D��+�l�����`b�]o gs��	�E��~�
�tγ^s(R��:������٣� ϳ9Qއ���N]d:��4�9���[�,�wd��3Xû%ވ��{mQ2��{*��!$%�vGC��f�y����hp�:�m:��U�\:����f��f���Q""#����ȃ�|��N��Ȩ{j��
��O�Q^������q��:qwm�lp�m�J���br�j���
�n����sz^f�������nmm\���"#�����9�n�F�q���՞z��lm��b��x�\p{���Z�Ԟ�ez�Wr������&r=���_��%U��0����7Z���[v�o� ��p	D��Kg�-D\lw�;L.�u������Q�,3Y쵸���X�νi��Gg��:�1�~����_`��xRx�s)M=��8wq�k�ZE�%��{�z��%�Su�Q},R*���C��ޢOm���5/g!��<d����*�0�o]]������փ��]��" %�7_�S�>����'��^�~�����=-��[������})���z�ck��g����8�v���?U���S_fR��ꅝ%S�pU�x����D�]�SuL�-�<�Ny��UJ�;}ƣ0�4C��y_��R���E�J�'�}u��V-�Tf@��x�tBNh����#V����fv��|���y<Juyf���G][�g&��]�x���)�����!�L��K��q����0]�V�]5���ѭ]3��&J���� DBB��e��Wk]|p�	`n=���~=Q�]?�kk���o�V��2eڅ�M���pF�C�����t�_�Q��;&i*���,`�cy�;>��	o��13Ǯ��5[����9�yP�^���[ĝq��1�va,B��ڿCaۼ��вrw
��AH�����<�o{j�S�Ȱ��U�H�B.OP���Hç2�J�ՁW(�TgN^.o��OW|w]3ۈw�x���z=�7Y�O�;��yW������tM�nq�ڨ��z*Y6����,Sy�u��p6�7�<�y6^�@��X��IE�Pպ����� .�+¹�_l��Y�m��N�ub �9Y�Av�|�@����CZ�2��K�sYW���.��{"ev�ۃ����_y{@��C���64�פ<O�%DW���?�����?����9�h ������~��_�J #��@���::$���t8y����������������"���������
<a	Q�%F�XBT`aP�D��D�8¤J"��P B�	TB U��{�Q BEA�	�Q�! (��  @�����J"�!"(@�*!�C�"! @����@�! �@����H�!�@!* @�"�
H(! @�"�*@(!�@� .J/ BQ@�%A`B BD`BQ`BT`BT`B`B{���A�	Q�E�	Q��E��	T�	�C��B,@,J�B,B�!HS �����#�] �@,@�@��	Q�E�	Q�	E��	Q�	Q�!�F $V������H�O���A��8e���TB�UU	�X�?��s�������o����_���A��L?O��?��P��??���8C�3���w���Oן��pu�������������  ���*�
����� }0���2��?��?��U��A���Ƿ�����?�>������9�h �w
��<PUPaAF�UJT@��F �Q��bQJH�hHA)�ZJE���h�hH �Z���ThE���e�fd`X! e$Y X�eF$X��Y�d�eBA�Ye!YP�a YR�Q�X��a Y Y��a U`YR��d%	E��d`XHVXVDH��a!HQ�BE�E��` Y  Y $	F`X	A�`Y X HIF�`Bf�I%A�U�i
AdH�F�E`�a!Q��bTJE�Q�@`�"(AR�TB�zJ��� @�ZT�������t~��QR�B��EJ���C�G��_���(?��`���?������U{����������N����'�N?��c�������U}�֟����I�PD�������?�����gB/��?x��@����ÀI��8��ލ��� � _Ϭx&��'��xJ����O���~�?��Oڪ*���?a����>���������?��$�����C��U��G��j����~g��<
Oڽ����@����~��h�����$���U|L�&~?ܜ@�a���������~S������P ����� A�w��?�����!����e5�
���:�]� ?�s2}p$���UU
�R�TJ��H!I	%J�I
�T�P�*$���*�!ITT(�DBP�T��QQH��H�T���H�E*��D�BR�
�EIIE*�A(�za"E �JQ)"JT*��)*�**��!HU$P�eP*���
���A*�T�T�����DJ���DH*�EQR�D�D�!TE$"���D��J�J�QH*0   j]"�Y��f����S��Z���I�͕��m�&U[m,��T�22�emRVj�m���Qʥd�U�M��j4��eZ���@�D%PI
(
*C�  ���
(P��۴84�"�
(P�G
NV
�T3m��3m��Mmm[+
ce�)Ul��T�PiZ�Z�*��F�ն[cR6����P��*�%D�)B�  5qhU�E�[4ՠY��E-�&�Li�X�$�*�*ƵEm�d���FZ-�U��f��06T�����(PT�RT�R�8  J��Z�SBIh�Jej�"�H
�X5`AUU��
�M%T֭�D�&5��)�kR؄m�a��)E @�)*��  #�`�ҁ�j�2S$�Ulj��&�b�Ml�Ѩ��!UV�Y62��hc*"FCU���lRR��dH"��JE
�8  Z��QR����QMd"�%Z��3� �` L5�  5�`J�  ��������(IE$P*���  6�( M� Z�(�-�P��`  fU�Ҁ)�M�[j��  	�  �XP&R

��TTP�8  ,p  &�� j��f� Pf�U4 �4�e h1@��0hR�5h����UQ!DQR�p  � �l��M�(m%�MS2� ��U�
4�6� ��, �Y���ѠZ� P6`  �$��UT�(�*���   �  a���  mF �A�4�(�� � 6�` ��� �մ  n �~A6J��  "�ф��F�� *x�����  "��	JT�  d��	�&i�I����@��H»!��	�������nT ��Td��,ֈ4w��-X�?�_U}���}��z���HBI�!$?�HBI��	!	'� II$ ������t����/4�6ͭ��PdFyI���׻��I&�^T�ВY�N���-y_��$ �;Z#/x�T��U����L�u��N+eڎ]���R&#D���dnV��6�8U`��)+0�,��\n���wZ��n���W8�I��ZjՃh���n��V�2B�ؒ�!wULT�y7�`Ѕ�SǠf\CVn3����l^�w�m�N�42k�դ$���W&�k�a�� U陧D��3H��#�¾��8[��X�m]��zU�; t!kQ�y�i��u,ʴ	��Ө�tCgU���+3���S��vn����Aӡ�i�h�+H���YΒ1�v�Q��E{���E�
w�Qwi�Q�L��Y�-`
��f�AX�Z���B�=H
i�{�����w	F���)F�٠Ы��ѕ{p��匰�gk�&�`+�v��L�Rͩ)�rG�McKf�7V5^e50K[���ܩE�{���ct�8�a�H���0	4��e�$�n�/dEaB�cU�-�$Pa���sYVl���j�Q'5��&D���ǑU�J��Z5) ��Z6Xq�'a��i�w���/n�6�VP�圧X�X�"�LO]{s@pf�ѳ^�ʠ�8VZ��H�E`��nV���ү*����Ge�R�ӱY���o�ބ*<9x���n1�woh�k��)kO��n�LJ�<��G*nޝ�E� 4p��>v.�SSK�4TШ"1�]�4m���i0K�w�Sr�34�RdńM˺qdC.�ڠ��,�y�dkRo�s3{���q=�q� �����qէp���ڸlҧ��2��#�U(8
�C�}��V)�1��˗"�F�Sj\V�[J�����v-�ЩqSg,Br�dwq��5���$�۔�ש�У3wb���ڭki�s3貝�� �v��iv3S*��r��$,�4@�a� �4RRB���u�b���O,4��aiǰf\k짭��;�[uy6Ս+]l�� �`��w2�voV[��H6�iݲ�/�IP.�OU�Z��Z�%�\J�n#`I�2�^G(j5��a�6� e��/#����1�$`T�vբ��Q[YxYP������C�k"�[u#XXt�qZ�;h�UձPMۦ���Ա�]���)A���H�ۙ4T)���8� #�ݧ��6WP��S+f^B��&�=�E�1ڼ�w�$R{J��B�y�I���&ə�֘�N���3YM���^c�ʀ;V/UK�f�GM�����L���$V�wJ��:M6�t�E����bj���$�]�aV$p:x>��a,�2���#MfX��Ev��::�)b7�X
BM���V�8��U�L�N�̥��7�4��/jTj��4��fDvD#���wK0 �oY�`��bR7�̭f�JAdNiG CYH,��x��(ZN�����hb!kt�7{,�;Yf'P��-P�t�wFSiTi]���4Xi:Su�Y��.����Hһժ���B)`P�m;�!��gm	-դl:�[z���Գh֥�9���H�k-d��@YWe�gk3,���̚���v���Q��M�Af�-�<llSv]کq��h��KF@F�c�Z�[�J�������[)�=�pfQ�f��r�Py�c�
٦��-�k m�u��Z����B��WGF�ł�L��a��1Ś"�H^��,�@^�u2WkN45�[�����BT&�)-K�н�YIR6���rCt�F7B�Gc̫�i^Tȃ���O�wm�II��u��軓޴��i�m�m��&Q��tF)�g3FH��J�RźI��su}zR�i���`�b�Q
�E���=���q�y�,2%*�5�bQ4h�ۑbRMY�Bh\�����Uey��;!Ŕ;��	c
jr��U�(j8�S��|��ȝӧ��[͓so�f�:Rԅ�u��u����%�X��1�R+!��EԣZv��h�"ZX��iI��@mv��Ro!�:�d��$I�k^�.æ۫��Ĩ��,y�6vu�nP��^`f�ެ�7V��R����8�Jm����WztL��V­W���ͤq[h`"����mQw���Oky{�K{p�Y2D��ΨF�#4AN�e�YbV�܍r9�vG:9���Ak)+�K�����Z�ݗl\��f��*8T�@��,�v�����ד��+�j�2�
�u�eE��AZm����of�PAI;&l��a�٢+[r�eլ�d�c-� r�%���(b��M�@;��� �*�<�MĴ��c#�	�;J��񽕮�zv��>ƫV
v��4���(�64ы.V��)�t����8��]�[���[���yL�Hb	:���B�Vh�B�x��yCB]�G*�Gm���*��.��VM���H#��倥��rn#��Z^
�9�fq�`���`_1���Τ�իh$�p�ڕ37&�:A�:0KR��`�.�U�%�Xwq�1�I2n�-�dI�RУڟK��z%�!�W����l���8�!W���Z�e�h^=����0,�L�G"
�y5��8�[�Xwa'�M���w�h��g�^*1�1իXԆ�`Vn�"���oFĝ
��hP����%�m��f��K	ЮJƔ�n��k{��E
�ŉ��w5ӻViS˰�OPB�f���Lް�2�Ӧ��ֺZ�F �Ք���J���%��V� �9��a!�[��$��Iz��i?l�����cR�Z�]6���*���*�˷
2鹬�$��H�X�Vmix�Jǵ*���ۉm��#R���*.����]nN7*��4�K��5{P� ��᠆Xj��n�7uc6����z����m����'�m��D�kS��E+8��c_Z�݄B��Z����Z`}���x$������_�lO,|����(���Oic�L`�����41v��̈́�YXk ��V�M�����vf�M:��7��K
���M4Cu��ǅ�'M�NI�-Q�51��i���1��^����9lF�*+Ƶ����i��:� �4<�rݷ��[��9T�3��A�̣
/d�F�Պ�Bc����&
�-�,m�3Z>X2̓idH�ފ�2jIML'&�Z�V*Z�V��ՂQ�x�A���2���1
�b�����e�ݧ ��U�El�-��(�y��5���Q�HY+r�Ŵkp�z��`�c�� Y¦��S3~*C�S4�ֳw�-��-r�f���Zn� ]ȕn��P��=r|(A��edװ��E���[h�u0`�4��I! �9q��5���V�Q����7r����b���z���)�65��IUڗv��� �� Į��;x���go[���@�!�*�#ca��ZM�I�ѓ7/fT�ʓ>���_ق
+d۹h�"�$h{l�x�<���uB�G�,=�I��(�b�4���Z�9&M�7C��w^f:[�$�j�6BH����T�
	w���.�4��J��o�]���y����m]J�$��4�n_����R�RWag���e��T �j��c
�(�X�����N%r���Q�b�d6�V��H�H\JlV�`2���w[.e:iӺuZ^�pو�M����p8T�^n8ۺ
X�6`t�ƅ$�r<�Ŷ[��
�Q���5^�ۺ�0���1!qQd�/pe�:ڎ]f�f���SlZ-����D�.h��(�v��U�L����lf�`N���fV��v4T�vVޤ��O(][��m��N�=9�n�ˊ]T�-��Zێ�L��^�*�\�X6<�K-�Z�n2X�� l��a���_i�ַ�d�F��
[2�x�skT2��!�rĥٚ�K�9R\���nSu��óKȱ��!��F$ź!х=`b�r��u�3�B��^l�m�Ϩ
y�T7 Y5���5�5��ѻ��T�)ݱm�x�6�U����vA�U��,�p�kNC�Hq];�4]�Kd��:�R�e4%3�ʑ���������~��S״�G��eAKm��`�F9�I%�+r�LwJ�	+Eh��)f�`�q7u�� :�d�ۋv�ffY.+Pʰ�r���U��b�1Y���ѫi%�g�E�l�,z쇃,�̦s\�vj	�g��[e��!]AB�(LI��&�V0�qR�5�WN�e�S����c��%�乱;p��J�	zګ��:Oh�-�d1��Lr�$�������J�z�U�	Y�P�N��Vn��d�5JFR�d�m�F��a���x Ư�xQ*چ��r�<�SkL.J7�S`��k���`�e��NG��.��nEvA)���M���-��Z08U<�1�ƍl9������,2�%�7U(�"������rڅA�Tou|�.��t/Ѵh͖���"V[����]�ŕ�%�5wvN� ��Ҫ�6j���f^-�9���5��n��D���V�d���u6Ch"�r�k��w�ɕ��8��Z1��2����ٶ $dH�˷��#`ܙZ��L�0]K����!(�ͽZn���p��6X6Hl�r+����x��M`�X~#f�����4 N�1v�.NP��}�q����Yy�:�VnR'v�I[k4�TqA�d��I:�cM�x%i����X�m7Kv,��S4JY���/,�0,Z�c,ڠH�,v	8m�6���-�q�Q]�MV��6��M�q�׮�S�
2��(�f�-�wH7�t�A�r���b��75,	�x`�૽�ڃX[b޵����m4cyV�Z6Ԕ�;���m�u�tΫ�ُh8��]��ԣM��&d���ĭB4�n5��+F��@�[w����^ae��i�FY�u��fD��.�Bj-�u1A�E�5W�����7r�L�ȟ)��]]MT1,�¼�b�� �B�`�����-�Nɗ�|�G�u+l� �vn�S#Uy��:�bu��kp
���i}��	���CF��;yEIY��m �`���u��ѹH�qZ���Wq���zZѕ�R�Y�p��0,Ŭ�RKWE#�����YBa���h�R�J�u����{�0���4�j�=���4��1�E�kX�` �2��
YYz!TJ�V�m���I��{hP�l�jL�8ù7>���k{�]]*E��@�� d�"�vtֶ�GW(ĭ� �F��tܺ9Sn�Ն%	�z+n�)w>�SC�2�{a��`y��e]�KɹY.�*��nS�[k�tf�]$@����Z�l*�n3z���6�0�m�чl6.�a�X]��ZfJԝ�6JB��۱Hբ�e�E��rhCF)��V��3hر
�Y6ΣO xԘR��F�ʏ/�&q�J[[�+{S��hȖ<�Y�SN0S[j�<�y�֍@�-�i4U�ZΙyjcj�����d���Ҹ*���gd�ع(Լ�ѩ|��	���Z�� �	���݊�Z��'��I�H�֝E���f�����ƙ��/]��/,ҫ�� ��7��`ڽ��� ��������m�am�Z��)�W��/%�ԳI#����{B�^ JǩVm]c���0�4
ª?��#�m�:\a�ҋ�qM:M��)ISZ�Z��ݕ��i�y���n�Y2j�I��jnRwy�pn�Z��ܵm��q��6�f��5K�[�4^B���T�i��`2ɦ[��ђ]��h�M�Qb�]8.��+K"���3dZx!���_`0dM��N2�Q�CH��A�F0���<(>�l�vN�k �\�w����n��2%n��aD�]-jF)m%N��@�W�^�̂��^QFD��
�E�PeK$C���;�/eBղš������fD�+!��1m	�n�"��Ub=�ba���2eͥ�XӨ���{�$XD�X�֞�B�}zt��S�$,f�U�:OU��AgHgBh�%[�&�x�iy1E����6��DJ����,s���	�/
�!� �4e��!+*��Z[�<�k!\*ې-�mn�ޗ�΂�-D�ݠ)҇D��Mf֜0�񠲃�v�J�ݹ��Z�U�lMj��T�X�љP8��y.��{R����[Mձ`�8����$m��t���7Qn���O��*`�Ö25#Y[����@j�f\�xACV�JWr��zmM��9`#��tT�M�iѮ�52(�An˻ͤ�t�,V�I%Ǒ��Ն�BV�{d����3iLQ�kn�`��%`��f#��.h9c�\M�ZP��lu� �ܽ2��V	f�૦y�Fтc��aL���ZɆ��٫[� йF����b:�7L�h�t���Cf'x�Ly��;Q���M���G��MLQ`�
Ӯ�ֲ+r��;͇
Wu�!Z�l&�S�T�h\v�m�ɎZ,��Ђ*�N��:u��wF� <�#-���1:�i�v#u��V���Lb�+0�w���A*X�EnS���6�4e��3/�)%�LH-.�U:�t��VԘ�Β��x�/�Խohl��Վ�^ [��e\��V�r�+����6��I%h���<��AϤFVF��0�3Yx��ؔr�/r�vͷWR��P�E�Ł��Z�ÂՁ� b��Eͼ����ʎ��Zݕ�m�����0���DHTZM=Q���6�DM�j��!`���{��U�̖�F��ңr��ުT�ӣ28	�.RwomZ���-5����r�	R�*�1+ ��\�����0J�U��$ք��m@���^4d��ɒ�љo��+2�`Ֆ�5�M�D�?�m���Ue�
���ܾ�kS@b��S�N��{RF��f�*�"��������糅s|�+ǼU��+8ln��0u�P�wY���)	�ԉ�ؔy�̺}���}Q��J�'�f[ڸ��Ƭ2��wN6��It�����8O9)��.�}hn8	�^��a�鶴zA�5wjx��e__
�]7 ��,s�U��d�S8͈�v!6�q����l8��feh��}��+��1��n6�*�����l\�(C6��V�#���n&`�w.er�9ق����l_5� H���A�k:�����7Oe]��x�ჺ��j��U��ִq�|ث�	�}�%��-�n�y�L�&�K�u�х�����,h-�×�|���6saQO�7����a�]����1N�"����	A�֔�W[�3�ΥZ����;�J��|�^3�����9�`*��1�Ia�X��a�2g1w�-)}.�@+*Sg7n����et8.��� [@�b��w"�ộNd��I]ϋ����,��)�-ޗ�|��J��kӬ+��f>��t֗ȭ}\���/���R꼵.��#?\�w#� !7�]ƛk=�Ձ��^�8;B��7�ɜz��9jf�����lW)¸�BU�w@��M�r�x6��Т��؝���&��ۛ�k��L�ԡ�r��<:�����	I�ܙǀ�����c���C��/s:�9aoX����2QZ�:;Bƹ�D�;*!�.\ܭX��&����HJ��{Uj3p����{l�,z�'�a�?���!Єu��`O[���bܻ<&^�V���X���Pঌ���k+4��$�s�2���n��|��`ζ���U��:��}
���=E��Q�����[�p* �Y]o e�]Y�]c�y9�[]L_0,Vһ��Mv8�=��Q�^[�!��ͻ�K �;��yn���&�m_�e��ž��F,J������ֶf:%��n�޳jn�6Tk���el����):op=��̛ԫ2��;p���߽=�s�.���V����c�Zct�̳(m�1�k1w!H�Gi}31%s�Ĭn�F��&�VEv�3/V����T=v�sOܓX<Ϯ%A�{5�b��˘(Nʊ�+�0�Թ����: �v�򑴥Yy����NV��P
X`ݼ� [
��F��u�;�o���)һ���N��ԟde��wU򹍍��K=�e0y��R��Jjv�}mV��=}��4�����`P�[�K�k �7��˼.�a���`��w�����Ej�Ǳ�*��;!"��f��͔�f�)獻��j�fl��8�y�k�Y7�Bםso^լ���72r�<���j���8���L�Z���kx�;:�x�dG�)�Lt0J.���$u���b[Y#���Hyz;\h��M�uqJ,�6s��sp���
QS;��8�5�[/r�GWRu3[rM6
R�`w\ڭ]�̲����櫼�y�%�gL޶��Å2�����)�*h���w�M�@Z5=��8&Q������v���x,�WP���.�+u��a���O�QH��<Q�p@z�Sӣ1z�)�Y}]E�y�;���,��>T,])X�vv.^��;���o[=e9We��U�QY9���fԩ-�-�Z���7��PV6shc튴\�th�r�a�6����f�E/xj
��B��К��� v�H�^�p��\�(+lm9c�v[�7�*උ=/\���=��z��꾼��Q�t��gwD�	�E�,O��ߎ��5qV9��/���*$�*��}��^uD�A�g{j�Y̮��K	a������@,]I��\D�W��u�ucT3�d����lwa��G\���4=��L$�ƒm[��p��P�^���ޕ�����U�U氄 0p����ެ���2�KGU j5Wٮ���5rlT+,A)��u�m�0b��c����=�;�z�u��p���kU.����A�$[7Kxs��]^�o���+R�%����"�T2�	:� �-o����!��1X�U��!������/�֠���u���'�וg��I���)T�[�l�:}�e٬���������E��:.\�N��������֙=�v�¹�:"�S
:o�>����cvt`{�H��[ѽ��}O�(�3�s\��
ɗ�>l>+3�Sy�?j�U�����0v4ٷ�d5�
ݡz�N��Vwk����@鐎��2c
�Kw�f3`4�a �W]�q�Q�����4u�����J�`+��a�qïlJ�y�D5:keW;헩p=�C���}�� u�Tb��m-�tkWf��r�N�z� �0�5���9G�F�](���@�����v�i�U�W�cϾ��4�Ū�N]�:����B�!��W$��۰N�.�:iorTM��פc����5�+� 0���p�M-<�sUO�;Wc�L��Xf�A�ܣ}�D�T`h�04�J=΅�*�Lf��TFr=y�+.���� \8m��F�R�6�e�:(a�]�� Q��-i����}��&.�m�<�]��a���Eo�#���+���J6�ĳ��>ܞ#nXo�ӰS��Ü�b�|����YX�����;Oӹ�"nF�)��5v�^<Q!�+޻��bu����#��P�[hK�tj$q�ܙ�2M����#V�����/���%�&fK:�̙"7u��.(k�v��8����I���C��<G���̳oGS��s2�F~yd��9��l�����/�p�^A�3���6 ��K���WV�/�-q�Lz6�b켒X\��
���T�Vféگ�r�5ݴ����$��k<�A�.�='q����� ����:��㹭jt��hK�Эf�A��nj��%ѥ��\�l}e���U�c5�����g�R&*����ں7m��VmX�O�i�6d��N��߷
�{Sx]
"	Wuo�����f\��`���[k����t
C��^���9���G35��+&����4:9�f6������`�]�t+w�:#l�y�3O#�f�{�gP|�~W�s�w���0��v��D���}b�]���=z��Μ�pU�]��\)Br���g�w�'R7ҷ�H�P�v֕)�<�����sW�v䴷�W�Z�|��eEb�>f�!ݢv�V:�; �**;u����/y��`g0ͭy���μ�^�L�U�V>[��P�f��gP����Ź{���h�ɳ޹��|~�Z�TFU̝��Í�D^�ܩ٨v�j��Iq��'�]���?9�ht�X+�~:�8V3��E���g�����1D�QjVz����hf81��\{{���ũ�cS*����V0;E79�7�l��ǙB�Gj����1�#7��I~�&�C���2�]�{�X.�/���t�h���C��ȠO�4�o	ܰ�ee���zDk��3vDR�a"�6�B�P�Vk�����u���4o:�Sm�ꗨt�əT�
�P�B�n�en��i!r���ɢQ�<Y������R�v��]'Z��t��B�m��9��%I����w1Ӧ��PEZH�\y!U��T�R �LfIJ�-4�2�3�"��/�������G0��/ZkUw}��ƈ/;�H��,�D�f�Y�AԵy�^[���F���Ҟ��sɦ����E�n4{� 2sǬ�a�-k��r�Ll����]awk�F�jT}��핸yc��#�cm7�{�.\��Է!v�Z�Y.�W�Bn^48/�5 *�4:�Ժ��]za�(>.��H�>%�J�{���|�N�	P��]��U��RwFrЍN�n՗�(�4a(����Q�Ku`e1���;�o{���j���|�zL��������:�ղ\���]���;�ru`�Z��$���c[��:�� ��8v��Cr�4VYV��r��.��͞Gj�Uזs�rͧ��)&�6�h��/%gqΫ�X�&������Zi���v�s�|�F7���d�+u3R��w6��2�ڭ��\.�3�oQ:ý1e�лu���j�u�k�ӈ�3����I���0�A�q�F�����<GC�q;)@�ʼ�,���fSE���e�G0�,#�)��(*۽�U��N��2�;n���<��n���_n���MW�:%��wvԕ�>��y�(jUy8չ������54�ԗ=oS���]S���b֮�x��s��(�;e]Zڬ�ʈ��Wh9�ds�w�X��uY�Y�9D"�Q���v�����<��3Lڑ��[@�xg��=�;ݬz��Y��f|�PNY�y��2e^>��n6��}t�]
`��sh�
k��+���B��FAoL�����R�S�X�j���H/6�-T$�t�A��]Bq���v;�w�$Yǵܲ]�孋^n��$T�Z�a�q,�@2�L,�x�N��x;�WE�Q���%YR�EgWe*��{e���=�ln��(1-
ˇ��5����Vm���S;��m铟pfC��D��l�k�E�8�64��u�f���r{�z-�e�R�IZ�ͮ�:y{V�Nbgy�!�6�5�*d�8�݃��L�7p��쳓��i�ܖq� P03�[;�0����kŷ�;y,G���ը%l}�{���c��Q��4j�� PȸQ�u���@�4������s�jMA�W�G��<�yG����gQ��&��W�n��\�y�Զd<;Q8�ܓ���hz���j��O�ulr�fn�Q�Ꮨ��2F����p�(������6��CN��O�}�ڗ���ޭ�}f��{;����C�+B�0ڋ@�p`�#�ޱc�76�5��̧�9�& kM_T�r�s��V���U���@:���a�9qY��Qw�����|j�z^�y�l�2�.��	�p�{PS���=��w0NIM�JG�N�Ϩ�Ԭ>k��x�n'�,}�[��k�^�X�����?�+��>�[��nۘ�[�f�����\���@3�t�w� ����ެ��&��e>����V�k"�\���i>�j�d�\�s��B�^	�;3�U��+i�kN:�T��A;t;�Q�Z�0nV�&��n��sArͬΛ���Oj��]b��Juڮl.��r�̎b3�ۭʕI0�t�r��s��]�F֘�	���5�]qww�_*��9VV��������%cv��z�m��MI}7.�+��ېc�2���`Y{V�sg[h�� �>68d�@\Bw:s_Մ'�c��󓈳]�,͛}��rX�=[�y�w�����Ar�D��6+q��+��P��}UJc��hѢ�
m�8P��êId\K �	)�v����bÜ�9��8]dFKC7��\�fE��8&�Pi��h�!)��rˠ6�f@���]I镺����.D�$sE_pZv�X(X�JlM$��\R:n��N�\�9���yP7��0�jB�vcѦ���3&?��9�n(�.4�b�j:%�����%}1�x�^j=�4=��Z�|�m�뾵�И�s�#�p���6��5v/IS�Iu�u��['�!iUث��<v�ƅ�gq�g%.�g�55Xb5�	����k������M�����3��V�  �}�����軻vlӜ�h�r��pj�1Q���u���1�N�Y2m�`T�t	F���ޕ}&�cK�t�g��ƶN��xo
�'̫�(���@�)r�!U�l�۟g>g ����q�hU��{�!b���l�[��pVsB�]��ek�bY�ǝf=.Z5[s��d�+d
�ʼ��f�]�`mwQND:�F�=x�9�Y-Tn�������_�������ހ\�m�\o�Ȳ�7&��{������q�]2 ���{��c���3=YOb@mi/;�^�]@f]�o�#%}��ma��+Y�&֒�d��;��Y���U�z�ҝ���7#���K�`��q�ls�ܤ�Oa�x��{od�)P�5̑К��գ�	K����ʯ�7��9��J��I'���ԙ�1�5��#��r��1|
���+�K��v�[����Z�ݥ��5��y��͚�!/�+"�MK]��\��.�V^�3�+u�82rn�������e@��o�O����;������wݯ+%��،]��޾�(�g(�0�9̣�;.��y2y��l�5�kU���@8vѬ�~}������[�9���3����v��xn�w*�Fɂ���{N��"����0
諳UX}m���wgڻEp*w]tj��9*�㎇I��h���뫆�6N���fC�n)���W�v諸L}&`i�l��C��jRS���f�O��eJY;�r����c���5o���oO)�a�<����ƌ��v��\���?rU��{�nR��y׶7F�N��OQ��cq��x��-ͭ��ܮ.�r �w/�V����ͮ޶�ȫ-E���W{�=��U[�>���
7	�aHqԚ����TMM߈���v:g��5]� B�U��;Ÿ�W1	�m�{3]��gk��`w�i`��JЙ���8q�v�;��r�5,v]g?��.��������P�uu<,�=C�2ﮤ����Y�y���3ⷺ*LĬ�bW̉]��wk�me(l�� �vn�_ ��v��+��)��/{x*���,�t
��V�Ć�$`LM�Z�؇_�z �գ'd]W�5Eq��'l	�ٵ�s���2�ovô!�w��5�܅L��}��ۛ}V��}�a�o��.􀺸n�P�y��{���s��ī�	�u4<�-&;�a=�%�v�w�Ŏ�_��z��C�w����{�A�w��]����=�����$�8s3�_v.�zr;4�C����Ϸ���[*�R^oQ-������@	!��	!	'�?}��{��ʝwO�m�L��:��u����P��v\յ��KL�P{Ǖ�x��{&ͧGR��x��_R٣�����.�O��L勊�����NEȐ��\�:�`U��7$��e.Nh���c��}�#A7�R��ÚMK�^��EK�Tz��6����&�j��Ogj�=�^	���8Q�0��i�,��#8�T�JB�#v�1U�U��h��jE:8��4]<�u{���6�/K��cwk+:�[�x(��SZ�(�7�d�fVZ˸��Gn�L�^�3�Ʋ���bk$��3���w��]���"ڙ��WQ��u*h�m�N�j��5.���o@��z��������r�۷ta�E��Y=6�̙GuǼv���5�h	��T���׮���)z�I*����.�^��g/��Z���}§]�����U++ k'�]�s��ܥ/�cH����;�+���t/b'��Z&C�R�W&��އ7x&qGB����؜�}��f����]�"��4��T�en���n۾��\�C�������dJ��C�V:��\�E֧/N���T���cb�M@[4�l������ ������yw��h��r��Q�n�e��-ۣ��Xb��u��VһP�G1�x��m�����J3���Jp\�:Q��=�)ͫ�(�1��2�8�u�i���������oe��gN�@$n�m�]�sH��ÃeJj�_)X�w@��݆�:���)�.�3�A�Uu�9�H"��U�F�5f�j��(8�
a˚��d�H�^n�񾩘��[Y�[��V,ub�}u�hXTJu��K���n �wb]�`7t�!��Y����g��Y+)�V��؄;b�\j���w b�r�W,v��S�BJ?_]K:�at�.��$�����B��JV�}��� �h�]�A��|N�e�V�8 `t�u��\&f���vc��u[�݂�i�@4%�m�,8P��i�}��nxc]�a�v��YA����'8���02�#b��K�$��g_]�Y��Nz��׼u:������l����z1um��@tO��*kE�Y��ne�c����Q0�N�I�#�����D�5!�$���|W=lFz�w����F�59v��U�p�&��v.m�ᡣm���*-,wf�<]�m r,]}�#�X���\�ޣZA����EofZ�ݵ�u�I÷�����M��.�F���]��*������>cw?�n�E�;�6��K����Q�4B����fqX�	�_J�Q|��:1F��O5�����ENj�R�u��H n�Z��M�zjW�Q� h݋�b�n�I���KZ�(5�.ĭ�Qr6�ӑƓ�9b��\H+�ʌӺ�+�KyV�P�D�7�ٗ�-QA�]|���]e�̎eɦh��K�s�3-S��J�v� �U��L����fWa|Ɇu�],����G���{WgAtqWkO@�,��/��3�����{;qKٙ���g�&n�Є�X5�F��tv%n��v��I�gt�N�z�0�wy������������^�F],VںgA`��pgcQwm+����,�Y���F:�Z�n��4
 U��2t:�P�Ü�ۥ��2`j�52���z���XsR͝��aZ��/fhu�,����ݽ�N7��:S�lR�9�pf�p	�-�@[��Udަ&��ؙ�(X.k���A@ �*Y��!�|�@S%��6�v��W2�wƮ5�ȕ�UVe�����T���r���YK4�$|n>������R��ʖVZ.�7�0e'��Bгo-����/,t��(]Պn��a�[���X�� kH��Y��n�ر��]�4�7$��땧�I\�B�����9���M��¥9���O�_^A�>�J�zX�blmq�&�r�OZ�[wxRb�/V�����{J�{m�C7��+m�NŔ�j�6#Kv�9����r�9�+�n@ֹ�]$�>�N�l���[��8+�,�&��3�e�՘Q�|�`/;��x��vM4��Uk�:pn>��^Eʕ�H�Snku�M��i��S
YU��g�j�݄Y�+�F�\�s]+�z�S���E�ba"�r����λW
B�d5�q��.����x�^A&r�u�ƶ0���.����@;1��Ը�7�А�5;8�xF 4����2���HC��S���Aͳ�������f�>R�\N�Ƨ����W���L ��f�vܗ�^�٧w�r�Y��U4��
�|F]�K�v*zu�f�3ju�w�Ƌ�^��b�v������n�C8��	{)�9ѷ�y?�j�f�;,2(p}�b�pY������+�y;a�3�f��9N"��&3�h�A�u$Y�W[m:���F���i&�0d��5�NQ��Y�o�"��7�:8�'9X���X�0�n�K���	���rF�ڜ[av�Vo�'fV�b.��1I�CDđ*���[w�k[xQ�}	�]��rm;��V��=s��cJ�*�t�㜎�z/&������Z�'��AA����pm��%ikH��;f,Cx懧sxʲ�v'�ikm�įz��ǵ�b��w{yS-`��e��D<�E�E��vJu�da��*n.��*���j���8[ʽK�)k�k��3\J���>@{Ǚ��D���O�)
�MgD�SF6��Wl�:b̤N;�@]�qx\��x��x_j�v�kT�v��x���+ݙ.�[+t�DWp.v��Ø�,@���c�R뫷�v�W;�i�i�H��a����.�Tx�2�w'P��+�`p��\7��j顈��x�FSb�b�@X�)���_v����]������F�-V���J����t�6IX�F�J��{��{X��+�X��Of��W�l�b�]�t�a��j��R�:ؘ��Y�@l�Wu9uV��+9�r�ڻh��}�m|�{E�l��Y��[|t#Ia�����E8�0�&��o�q;B�)N�ᕪ]���s�Kn#Krq��mlڔ4�Q�:��
�J�P��J:Luld��h�u�7��NWc]�r����LV�i�
4,����V%��B�\Q`�\�n_)��`������A�I�7���VQj�	ݙS�`:�}X�-�o7d32*3����6�	��	rc�P�g�w0H4��sz�ҝ��D�Z4\�ɆD���]�jB�mm7kx��z��"%5�82�]�Yw��et
n�:_V�$��od�7�ZqFr֝.�,�t�9;u�{��Xi�������ˠ�au��D��6qN/5Cw���.RwV���7����ud��A��S�k����[h�6�����B��!	�r�Fv�
�d��KwϜ�
��ҋƥ�yw5�,|��dN[�Hἢھ���h��owp��tP��;�fǴ�b�]��,�7G� 8��9�*�ui;[��I.���#����v�c&�o����$Z�q�O.�����6�[�f-�u�C�.�	t��]F����M�F����j^NJ�}o�.c���J[s����o>�Gq�t�����o�-�@Ph**[Lo+��'
r��L��E�Vf�#7�*�,U��ڎȒ3Ѐj]mc�wL����C��Ƕ9���y�OwM�5@6u!�%���^=A��6�t�t3pЧ\�w�>�Jͽw��)wP��۳t��:$ޢ��V޷N�+7�=�B��S�x ��,��o�Պ�h�w��S�w��'�Jʗ���L���բ��q�.���h-����9Y;�Jmqw��E�J�w��7�/�6�6s9����[N#*�V����f-��}�Ϩi��<e�a��]j˅�n��j�*�A���7I{Z�)(nk4�V�8/-��6]ϥBܣ�Ǵ��)��x�@��ǡm9)Q�w�tJ�bB��]Y((A؜ʱ�] Ր��vU�\��VAt�u
Α=��&�[�M�v�`;Crd�#����&���+���A�=�	�M��t4��m����v��]뾸懇��pr�O��
k[�v�n�;;Dat�.�������L'���ʽ��X�Z0���,-�u�Զ��$��x5MV�M�(�Xr@L�GH����$�ި��	t&�<��9�<۟%t�o.Չ]����ӋVϒW�R��3(Bv��JE�C��:,B8�d�w1�k�yWjwQ�]���Bv�pu��FP��-���{�愍�E�'5���[�����z�ֱ��ic�*
�c2�|�v8���*R�����)�L�L�z�.�Y������I[8&7>��%(0fV!�S�>kWws��i�[��.�jd�*�s^�5*8��72�7M{4olwB�@�=��5����\,]���-�;�tw�k����̼Y+��Tt�g<���%�zˬnV�����,t�2��F,&�0�6Q49�V�*�p݉6hZ��kЭ�2*2}AQ
���y�VWM	c��qtg���U����4�S�\�7�;k�^F�vVWv��K��h���M�sx�}(ڵx�tv�2c�P�t���#��+j���Wo�q�m⾅����`���V���nu��;+�,��C�/������%�N}�I���WY��UE��\��3i�/F���KG��C)�Vw�Z�\��6��߳{"�JqV���m�i�pX�R�Rz �8���5�f!�`5Ig/�W8��[W)��gw*�bY�M����xGn�e�j�A���������(��6j�ٷ�Ń2J���.t�d�t��e�`�J��Zl�9���x���^`��Rj��܏&����zE����U�C"��/�HC���B�v��'iYFe	��TY�"�M�
�N���n�@+�z�ӳ(�AŽ�Veq��w�]�vfSװ�7���w�����^�!!��iG�d�$�t'7������EJ����X��7�'�V:f�wG@h��y��u�V��M��r�a,�F����ms�}{�I��h%�s �1t�i��\�{%'K�F�_3� Zt�i�[|�;�-+����h��2��k:�!�ge�͛|�R��h��Y� �[��ErYZ^֗*��h��86�-�5��LἔAb�Kw����y�5t����{�@Q��"��*�-<��u�N�r���,U�˽b���P׺)��E*�<gp�o�n��Cw*��Q��x�1�Xu��Iܻ|Ѽ�e@��lX2bb�ud͟��� ���K<�.z�)@E�!�]�����`�z�&�x�s��ܣL�t��|����i�x�sB�Q�Dh�Ќ+0 ��	�:�h�3��A�����xk^��N�Q��ޖ�Au����9̥�)m�1���|��v�6N9��JCq�9-�m#0FD�qb�-{�;u���;[�fAkP�ڸd�޲��,�V*�s��+g5�V8{Dee���Z���'}t���X������R��t)��ބ��y�&^�6R�]
��cVSz���gYJIW�*V�A�]g
-�90'6�W:�D.����6]��xS�	{�eM��{m��C�(N���M2:K��Аm�)һwr8��$4��Ly����w������tcƈ�&�n�:�>NB���J��� ���i�V�!D��2K�-T�2�s��[N�ބ�o��O뼀a����N�ms#4���H;.nV�ML]�Q)f�NH���[�>�d�fV��nr�2�phѳ!��b�p����ܜİkK-�
�t��O�ћw�6�i�g%\���wme�f��-��M����(�"�W|:
2 ����Хm֐�i��C&�]�34�iWP�־+k-�e#{�����ǜ�9:����v���Q�t��i��zkX��
�G�,ءp��s�pU����
�Z��ʺ��
�Lɣ���6t0���N�6c����p���(}�v�ٳ��JX���Q����+�ʤc"؍��ܼ��B�hs@���r������Վn�1�����w7.���\U�ز.K�
囻e;�wa�yf�	�����-�L�,��@�ɠ�9�
we�v�Nq� ��/7(҇"`��E)2���]%�-W$u��;:�Wf⃥�su��ACM≯�l��g^�yj8bɁw�yoq�"Q�CU։��2	�uf��ZІ�IV�H���#O��g%��0�E;x�&[0O���6��䈻�0�6��ow)_�.T�y�����:��0�iP̼o�$�ٓ⑁j�|���%���H4�Ma�sh�k+
�G�^Zrp�/9���f�WV�,tķw��.SC^+������nbO>���v��^L�ܪ��T�T5"��)ܖ#:fm:�^R�׳]8[*R��|�9A�����M�Xk�;K��hw7,J*Z�8(���C'�f���m;gKW�̖�vT��\6���r4~z&�-�JU�2�p�gH�28#/D�X.Z$D��;�V�+����c'�#��q�<�a������\&j�W+ݻ �(�Y�:y�o̨c���9��t:�&+fmkAy|�7!�(��&��FT�wM�\[˓����JQH��X]E�
�'����h0�v�Cr]gj4G�Q�������K�K:�b�5���Ú�m�(��1F&�9��M[���v�ھ��@����R-�����,۴;�Q��P$���}W�L��`��\,���#�}��o
�9O�ֻ��a ��Mn<�	餡�;,,:��w��2ˡ�Rwbc{hi»�[�[C�fC�)��wu��y�>0��22�5�]ӵ�����|�j�[@�I>��%�H^e���pQ�Y��J��j�c��J��ﾯ��Ͼ^�'�nb�T�o+}�fe2�=v����V�.^Ա0��Ӫ�qz0l�4��	�2�y&a+�|�r�1(P�9T�`�]�}a���|3��܂��
dk�o>��$�%����q��~q7pr�=��;��Ef�Z�4��w��Z��t׺y��)U����B�Z��-RP2��u�@�Z䳩7�����(R`��N�m.��}؃��nl˴#�Cw�1���+���έWvszk�!����( �(a�R�7,V<7gk(�Qmڗ���h7�,Xs�&X�H��6�F��X/(�Դ�ĭ$#�Oc̓�;vm�@m�Vo�蒦p��駮���Ɔ1�mZ�:�Dho���t�̶1:�<%�}����Z�,�N�5M��q��+��~;�Ć�6�ˊ��e_4d����c����g	��i�S�L9׀�mi�<"���:ڥ���x��c�1/k{.�0���2���`�101S�P���RPk�}��J�Xmֽ��6�Z�͢�VVg_>�0�+<˥ð��g%�7?�sīql���|r�\�
��� �����h�KU�tfu)�ܪ�u%��:�7��ֻ�ܾd��Y��/ys����ɖ�a�u�7�17�\Ũ�� �W9�Ѽ��X+�h�ݸ�W�Z������*��TQTXV�b����Ƶ��UR�U��Em�"*-�X�U+!Z�UX��rE+D�R�*1I����)Qa�TX�)J�AH�"��,�Ud�Z�j�DH�"1�iRf�kb��(0RТ�� ��E�����f������**���2*"�fB�SZ�dڀ��**[j)EE��D�QB"�Գ5X�X��PD�b��ER�QQCk0�R�U
�V
�F1
�a�ETV,���ET��DbV
#+*���&K����E�H���iAVm���Z�aU#�@�TJ�b�&@TBҊ�-R��j(�����KejV%�m
���b��4�*��TQa��!Z�UDX���%ql�Z�(��ֱb��QQTP\�k`���E���sPP2V����ژE��J�Q��(��֬X"�b�%`)
�dUT��Q�\�Q�%��
R�g2[fb���V)�X�Z��Աc��3����������E
湈�Q�E��Y��d�ouX�d��ض��t{%4\���uzR'x;G<W)�dn�a��q��L{ÃŻWشM����6�g/���foH�V*���1��<?|�,����WZT*]*/�h۴��gMo���?gw<a������f��/�6�~�����J��,�Q�x�8LX�*̥�IA	:u��\�f��l���b�0)�d^����=c��A�r�2}�V�
uk���G�!�옕�X>z��j�#h����b��v��� ��B��*&r�ܙ�®��M��ub�N�4�ҷĉҔ
v���xO��UJr���&1��e؆���:$F��:󠑗㸳�]fᬘA�s����R��Jvi=.��J��Q���M�`~"sRY8�4yn�[���t��p�C�~7�yc�w�[f� ?K F}� j4��%OL^�>�nll��L�Oջ.c��!�>�Y�W���U�? 1�x�p�����41����^���?o�S��7�X����,!q�'MC�ք2	�`��y{"������=Sk��"�����"��*h�V��%��;G!d�N��N�������
3[����*.�����Ta��}���f͔H���b
���������\�x�}�}�����'�Հ�����h]������m,nk��X��vS-ւ,��d$,�	���s��U�t�g�8m\���^1y�c������i
5ԏe�[�N�#ɲEǵ
�3)ߏ�>�׽v!�;�a�zn�S��YP�n8�F�.V���}��d��uJ��py^�'U��k<T��q��+{_γ��� 2a�y���d���뫲���N��>zx�]���1b-�J����^�i�^������/�W��]W]yJ����u'�
�&e߫����
5uO�y�6�Y�L�X��	�:�{�FG�~�ⷖs �_B�D_T���H�_���W�U��_?zX��g�f@r1�;e.uǨ�S>�P�]{Y2��9.@ڈm�ꠁG@I.�Y�D�.b#�~���X�Qs�Ym�y��s�s�@෬:��W�*��ū�=>�s^D�u*��G\�c��W�.�y�lՍ�#�/�<>�2xTl�QP��b�����ª �k�ԂN��7�u{C��r�Υ��a�n��?i
�j��<�k��������r���1E<��}��^�lL���B������^a}���"��;�᧽wx%�+fa�7���Y�	�eE;��5�#�]��R_�N��ʛ���:B�΀o�v����w��\��%==�`�|��V5��^��~�"6L}�x��g�$]�D��zWWZ�����$�q�8ۍ��v�h'���c6��@�ee�k��/3>x��`N�P�;*f��=��WB�w�zkA[jq��+��>׹h��b�'�^�*���V�[���nq���b<���Eǥb���f<<�Q�ϛ
�	戏��.ZY�N��8B=뺽ķ}���=?,�{p'핮d\Q�������܀��p>ժ�[�v͙��}���#�.�R�2���S1x�/i�HV:�~<�'G����y���^u���k��F�|��F�=]%��]e��J�8���8;��4¨�KLb�L۫�m$�S&��>�v�_��	F*~�����ʫ�Uk�P^��è�(G�UK�Ɖ��L{�>�T�4w�,3�s;���X�o[�	����;���k+Z�3�j�/��}j��J�����xf�����j���W�K����F�N
�v�/*$+�2F��5[��uG9ب)�Т��K�a]e'�޿-�jn\G��W�m�#F�T�wD	O-�C ����o�&��a��Fǟ6�uo�3�~��|�+�_��w�T�=U(�������(��Ó>[K��U�e�g2�/5��'dU�r�vΚ��M��X��z[ŭ�}	X���*S�J�5�0@�y��} .ׅ�kԓ�uy��t����^t�(o#�:��v�8�Z�w�;�Ȑ�TZ�m�s��5t�!ǈ!�u(R�_M��w�{;5�]�Lo
|�{�r� 痆e�\-�k¼�zp��~�ن]�7�\�`��zUҸx��R��8�j����i?:�l���*�R6AC 1%9ZIm�����f˥�m�WV���	� ��p"�.C�o�%�ѽ�b��B��}	޿o�u��h��"m��Ǿ��K����-����6�qxfLp^���r�>~)R!��������7��"RUz�k�<U�}��|eF�?z����5b2�s�c=���G�nȧ�u�;��~քg݈g)��suJ��yP����U{yeVy��v��qܺ�|�b�0�/���|�M��*�z��(u��TFl����!�e <�"�)~+!���UO5�+nrޘ40��s��c�۔�d^t,��P��_�� +�$8\������߻w�y��U"�{{�����-v������eyh��`ӾO꾾�NW�\��\��u��b'��:w�5)x��)z�9�;>γo�!�T�ۇ���O��V�W�J��PQ�[~��{���+��Wc'�_VSv�	��p�Wyrے[v�!�^	ۙ���2��X�:�R��)fT��<�i'�x�K{h���ښ�����mK`v��}]ON*�P��X�ܛ������fN����7��u���,��9�wa�����4�}����2�v����}<ĸ��0)�Q{��M�\4���<�:���v�j���f����5^�մ��x��~nX�p6��C�
E*<����v۝����������/>�b�3���.����װ�W���f��!�]+��N\�R��
w��Y����ޥ�YU����KG�B��%x������!�b$1`�*`$��E%�=6���X�%t@f�ݨwe�-��k)�\� �
��o+����+rkMS�b^x��i�{�:J�B80����ODK��y}�9y�T�C�c�]��>;����o��C�x����2���.�y�O����~EO��?:�P�7~�>��W�+�|`�������ܯKT���@��B���0�N$�P�����Cl�5�Dϩ�	$�l�t��/�©F�
�r�S�|�2z����jr����m{0E�XMma�1U�)ڻ�*N��h����k5,���Z�W�;���p�O�=o�J��D{ؾ���iI^M��ʰ��W�滼��<p��I�����[O�
w�M����$m��7WFB�f��XJ�ͻ<��q�GKW����&�e`�<�C�vf:u'��ٸ�D�+p�����n��نPҪ�ښ�U��u�������: ��\N	L�']O8L����>�.�#���ĳ[��B�1�Z�^���� �<~ R�@*��~*��}qN�}��d}�yg�W���oA��[�^�V,��~@c���_?���q�@�`-�){��Z���p�Q ?��h4��[(xo�yS����B
eZ��w{Ϛ�5K1��g��8�����T����=_�ν�W��4�k�|)�z�̿
;
�!�� �F۬��^�{��۝�!��"�ǧ�(P���Ex�V��f�7��(<��]�o�Ô3 �� �O:��5�T��q��������s�C��c�b�ƦR̰	&�v����&���߰h���z��Ul�h;��ˊ�Qx-�ʏ+�s�GCU@�x��3�u���^�B���PǉY��W]aC��>޼�m��?4�P����z򵽮�H=�ܰN��u������;�`b.!ԑ0��rF��3��"+%�ѐ)����W�
�K[�sn�@^}���!
%2�ܧ@kwD[� L -5���ƀ�q��^�i�1xsX���S����i�jO��]�K�ov��ە��+�Q�'�Nѧ���V�g�>˷�RX�s����T�qtRX�:��a4��W�n�"*WZ���}+f�9������uc�=+���\[�;B��x��D��79*�|/�.��pݹ[]V�"�G֓y#����>��#X�z���^|�Q?o�Y��=���b� mge�;w�w���N<��Q������]ǆ��0���,f�%���)9��a©�5���NW�39^ę��m�!ڶ�>�F�ٯJ�^���*��ƚWѳ%�2]�W�`���^0��/{�{���U�W(����Aer1���^aV6�Ȋ6�������燭��O��ف���[O]�� �N�J2�`�}�L]o�kO��f}�=�UySǯK�6vV��ڒ?�9�����g��/�,B�(W�/xSYD{������h�u�����/=��V������8NG�x|�#��N��2.(��7�~~9�uѺ�u{V��Lo�Ǜ �O��8��+w*aD��U��>��!X�X�~մ��E-�\��4ǩ=���@��x@ʸ��r����9
,8^6��
���Mpʉp�^8;��M0�����9��՛h�E�qꋓo��LfoG��F�����)r�앯�A}��K��eZ\+D�kåg:�gt6$Ew���5��M�{J�C����3��NNr�x�nxX�0j�[^oB¡��n�ܤ�l�2��nc2��|�i��܎�q�t�,�z!8��R��
�[�ă�qk��s�1p��%�W �b�V��X'`���؃ׄ�lb�t:*�����I��qv��۹��;C3{�F{��!+b|z���f��ts�P����U��m�\�~Մ��L����1ؘ��׸mV+>�LiyQ!` $@�㩑�`����0����N �����W�X^���{���X��}ưV�S���~�C�o�C!�L!G�^UOsg+�"��M	J��`��A��5^ߦdC��U=\�S��*uPv̺ L�z�ԎÍRկz���Q�>򥂲U[`XC�4���3(�|>��+M���)�#m�RX�&�bkҬm�1 8m
�Q>��77Y��vO���e+�>��íapu��~Y�٥�H�}ͬ]��{��XԆ#�]���<G��R)��"��t�o}��+�Ew�`��I���kmH2����J5@��uL<���\C�5��#�ÿET���ϥ]Z��Iv�O-n�l����˄b=���ъX,�=����h{vrL`�d���J}Y�o�s�������+B��r�����G���`��{�����n�ϫ�:� 3	_?ICƧ���j볨�`Ӈ���GBS�����WyΤ�u�ћ�}�Z�j���X����۴|�P�Co����d�P<�������j/���&���Wnu��/�Zh���3U�� �l�#�X�q� �^�0�]Vb�_ /�4=���}ؠ�������xr>��`[��yյ�Α���fH
7Ss���\zJ�g��s�/<����}�񷔳�׾�܌��uc��3���V�گm7�R5�s�]}r�x�Y�����ޙŹ�ș�6��Rq�H1N�`��܈y�UD�:��8�~�T�{��׎��vt���3θ^z\+�j���x��pܱ���Y;G���0=������'^y��ܧ�>�>�O�%Yb@�h�Z;pb�u��L_ڶ���<��
y,C��%ɱIoB	al�b~OF���n�fY�=Fs�����^?������؏��H�?R�v�e�%x��SS�c}��-�1R����*���%�M]����Y���X�)��rʷ	���݇���������Ws��*�-�5�}��Q��厍[��C�^r����İL�u��z�YPE�;��П{ȿ��4t0�y`U�w \��m?k>L���M��~C���C��ā�`��w�ZW2�?^:�\㌅"�Y�yw鎋<�`]`��D�����v�5���ܺ�i�J;mሡ�z��h����9�������2Xe>{R��{���W���'�uн���`XkxZY&[rq���jV,g�k����*$,�&�p��tl` ���+X�nt��)�^�Y��Q�@����\�����D-S&���#��������VOLבRy;�؛��{�_ō���ɨ���P��Lb~N$�Kj�x�Pa�^�^�O�ڷ%�~ޘ��ڜ�����l�%�	��Տ
u���� ��;�#!g�Ӝ�g�i�x"�H�әm�;Tֆ�˪D�����
�p��W��@a���xQx�+����;]�=@Q�R��9;��N�>��j�����ݸ��1���u��_]�����K9��o_v��K/s���&�C=^��(�;M��ߧ��ۮ��o�f�/�T5~.�P�8߁;��Z�ov�4B�`h�
0ǑQ�.��^���G	�X�v��`����X�mҦ��B�|��򳇳1��s�;�~�(Liz�h�Ɇ*!�i�u�@�vVRwC�T�L&�-y���S7 8n���zX�c��]|��(P�m���>���ϥP�kEf[ho*i�����6��I7H��� ��_E�F *"�u����U��V��E��,���kx�ϗ�����is@�,���e�͡L��U���=f�k�V�f����G�$m�<S鳵pov��eh��W[���!��20�L霟P7.;]��bc�&�3�S�i�7F�T��o�r�ް�>��&��bLdǟu�ڠ�msi�_sc>�gj���Zn�	�%��؞sm��	�SfԔ&d9�3�U��Vmh�KB�q���Q��õJ�U��v��|����ͤ~z�����N
��K�F�>�Z�����.\��oaŹEt�n�ʈ0��̈́@�6O��^��q�ֳb�b[�Y+�i��Ȫs���4�������\eH�q9��H+�����rm���q���!��cʕѴ���LB�>�TS�c6�X�̸�$J��(tn%�[wM����w���㚭 ���(×���-$'Z*.j�ϕ�.�ݾ��y�d3�K)-�2$�[��,�y�󳯎ڜڟaVm�śثM�f�av�� �ǜ��)�V���*;�vz��p�ɻ�P�Hfɹ,gU����"�b݉0z���٬�C��XAQf������z�}ը:dI�8�N��5�F��F�ô�WY�W7J�j���;�v��!n趑I�i��c���MACV��3y<-��������e�5�� ��{.����)P�|�}2�ϯ\W�����7LuP�؊Q��U(��/�tl�Ne4���+k�y�%���	�-历�B]�ic<A��K6V���ga�h ��V�
��+ a�3D�z3�:.}�v��»���9�CY�YZ:��)���������(s�|�T$����z��X��rL�FǏ1Ź\�W´vV�=ښtpى���K�^�k���w^W>��r���d���Q��\^��%��CW�oݢe�:��Hu�ٱ�L�:8ZY�kmj�k$�9��Ζ�W9[�L��
��.�e���(^@������4%�C�|�N� դ]�9��6��d��Җ�[��3F`��Sr�(G��9Rj�2�M2�5M�U[�YW�Yʝ���Ҵ|X­�	�	��$��Y�ɴ��]��i���g*�'s����+^T��͝����Qt*6d��Un�0��[6h�+����v�nVIx�^k�� �ׇV9�+�l��Z۰F��v&i|X�rVF9����*�4Z*J�څ��_K��׀���0�]�7@��+K��xt[�)q��|J�5�m7t.�H�"��]�gK�Bm<]a�ŝw��Y��L-��E��ɀC�[Q����qzف<G�
JoٴI��
��cf>���Tk{ld����5�U.a�h C�,���O]�%�w�Blp;�K�Rl�0jV��.&\8	���O�]e��c�i�P׏l
�ͪ������mvn�%�6�
Z�a�p=�JyA>�b���i�3�ݶyd��V���m�ϟ.�j�96�Tz�\b�m�u�i�Z�
��^V�0f�uݴ�;WCq�|���~��U~��,?2�1b,UEU��E�b�MB�� �TUBV��-2efJ���̅T��`V"6�C!R�P��H+�aTE��Z����Y�-�P�*AF1��DsR���IR�PU�c.e.�H"�cX�T
�6�TY"�:`�Y�PmmJ�Dd��6�E`��0�EZ�
��V�,U
�R*���*��"֫���\�QE*�H

�((,)
AX�&L��EQ�
�""��*(��()�J� U���DEF,P��H��XUeaDm$�U*ԙ��"�[h,P��UV�+1"²U+��dU,P��d�ְU�EQ(ŢE�dR"��Q"�H�*,��Q���� �
)A`��+3Qb&J�T���*lF�m�AAEEb6�j�#�%�(VB�ň�\°]i(* ��E��H�b�3(�dQF>>��*�6�8_Kސ�R���[��Q+�Ő��{� �4n�IW2r��f�H��o:�'˨�t
�>�#����:M��>�J��$N�ͤD��3$�opq���S�|���h%`|k�?c�}C�
�ϔ�*�T���@�/����Y�%@�"|c�}CDh�����MՓ��9����9ߡ�?!��T�[��Y�%��\���8�Y�<��C׏i�'���8�'�T�*���q���q�_���P���v�'�Cwg�x�!���
����}s�����Ώ/4�:1&F]O}�"4G�0�u��&d�5�8��3�'g�n�*Vz�U�ްI��<�B�r��V~���HT=L���５��(x��5�V��������+���4;���;]���p͛����G��B$w�~���|s:>}����AV'��?!X�y����t�{����钲�ǿw���Y;��qY�T���j�I_�&N��v��O�ȳ�>ww��Nt�s�f���V_}>#��(GON��}NV�x�P���g�|-�!�J�C��gV�$xã�9퓧��A{�@D��Y��s����P�;/��:@�X���=g�*w��9��;�RX�ۙ��J.�| CAfb����>'����Y�%@�;���%~�2)<J�ė�P�¤�
���~�:����%���N�W״��Y*T�9R_<��`/�8�q�O߿=��8�ޏU�c!,SBz(G�"G}߼��T���v}����C�w:��iR~N�|����_�P�=�d�}C��>�S<C�,P<J�����H'�T�?Y�w�DH�#���^<��^㾅��{�
��@x�L����8�PP����w�����?|��u�B�a���2���>�p���;H,�'�?9�C�}N�
���>'|B���|a���}�$CG��ݞ���0N�4}�˼�����2Ĩy=�N�ҳ�J���i�O��L!ĕ��v�=��p��V����q�㕓�|�I8�|d���Ϻ����~�w��=g���=?}�c�J~���c��I�B���(���V$����`g��|�����dSƳ���^��t��UC�=�C�8��W�>�Ϝ�V}IY:=�|N��+�>�oy����>>$F��?}B>�G� �����t�ߚ�ة���諫��,Ge��R�*��bJ���;�6����-��Kה�'���^�[����s'g�̀+�P��S�~����6��g�b֛��J	Q����(�C��v�jc���5m�S����z�SV���>��vvP�;�ks���,���NM�ӏ�7���!����(><H/a���q*O�V}d���>��� ����S�J�����>��8��}�����N���N!���מ��
��_RdHO�����9~�s�yoC���(����2:>""�������P�݇L��V'�Nڐ��������'ϔ�;�O����f�I!�1��rcG�}�9`J��ת�ԧ��~���{�q�I��=�H�z�C��%{d�3<N'�Y�iY+>|���L��T�|��8��+��C�<B������T�'��?c ,������}�#�wr��n��5��S�LOD1h�!���#A"W����:��H,�����>&I��~p:H"Oω�r��jozǩ��*T>0����̟���Ğ!_���F�}b"�Dp��otUOF9��?���u��|Vx���{g��=I_���1��P���θC�=B����$�b�
���ǈM�8�*T�9_ܰ2Aze�O��Ak�"�c��""�:*�C�w�ћƔ�~q �g��'��1>'I�l�C�~C2|e|aPY��M߸2NЩ�߽��N�<JΓ�=��2I�u�c�+
�做�%C�&~'�ܟ�����" ��M��,���⒫��>�HV����7��y��@�=}a�������$x�O�z��0?� }J��:;�Ʋz�Ϟ��;@�Y:<��'L��&@�/�H�"����A����~�W]�3=���+�;OyօB��>''^�ôPv�^�C�x�'�O�g��E'�W�S�q����'�^?Y:�N$����N��g��=��
)<y׿�;H"DD,�ҕu��I�O�����=�#���R��������f�ι�Ĭ>��Yĕ
��^uw�}a��IY�v'�%~���[ x��tj>�'�W�|dܿ��5�%���B>^F������s�z �}�J�����|R
Az��ɓ���|���������t�Y�Y�޻�}C&H)�4>3�2qé��>0�/��i��R|B�~�Md�Ay��ryȍ:�/D�Q������ڼ<��Ŋ�^�U�pf�#Pq�z�j��;����e#/�10L���+������g��s�g���ry��г{�Z�O>��uve�is�V+[�uhںe�NwH�9���]P��`T��~���|�d�n~�P�%C�=Lެ��P���z�RXu�0q����X�n=0+>����7(|O��Ag��$�8����Y>%k캬��30�ī��љ_��#�}V�a�������hR�VVt�I�>��+%eVz���'�OP�����t�i+8����Eg{�8³���'�?N�� )=B�Y�>`����D1����#۬x���C��`{����a�Ή��>�8{��yWIf0�Ἣ�ܩ�.F\V?Yz��ZoX�ya��-ĺ��y8+�9�>��/�����~T/o��m�Ǌ�Ci��bRY�g[��~\���}�W�΀��na��4�_ /�cC�>��ŏ
uܽ��>�S��&�������v!�}S��
V@��ܥp�{j��J%~2���bC���K�X�]z���5Ϸ�]o�;��o�׈�}�^�)�5��>�U��)�7�}��wN]T�Ǻ�k;�SZޯL��5+=sB���1�T��6�1��n�
H�zw�C ����ڛ�wyu�ou;��!'7��*�T��)�7N|���v�A��;x���1�׮+��������sY�Ԗ��Z<*�(7_j��������m�;t�-\�A�F�V_2�s	o�����+�*��3�E���j�C�Gک��n9���{G�qe�����2���fϔF�8%���</ƞ]��v#¦}4�pn�}��WZ?>�����#�_�*hO�iNve�'�d���C��,e�m"wg5���܉.��2�~���U,}��|�9Q{�ʫ��3��tJ�é��G��*lz��o�=���2����.��(�4pwnH���A(��c2A�����ň[�*!���h^k.��m��VJ�4���� ���#�/�,�o�=�5���p�z�7��X���9���̾�a����>0�_ڼ �e�*u TL�+��Ϯ2�2�C�{'@��?/uf���	�Ľ S��^Y�Y{���]�:�殜����D��9d�s>6�ǟ�hK!ϻ�пZх'�����*�Cƕt�9f�U1WP�� �p ����÷n��:5@[�c�*���.z�)!�N"����J=N�A�Œ��fFU,I��1�ױ^'rgtB���0Dh�o%xCj��aYu|�(�\������Gw�c�t���온�=3gـ��Z��э�/���{��{^G&�@@u�`.=63�ˬ��Znئ���)�O���j{�̫���k_{u�x෿�>7K£q	��v�����4�ҕ�	m���G����]�C-�t����.��W�s��|1q�TE`�w�`�q�۷*�V�u�%+�oi�}v��e�W���'FP�W@�[�r��R�1c�!�Xw��:1�ͷ9M��P�+�x�-�@N��)�1��BY~[��I��@+6!�.�Wvq�Z�����VjTSS>?W�a���&4�S�rL1Q֘�N����@W�R:�9����gr�t��G���򗈼�҅��hw���R#t�Sc��߹��k2�3�	 `ۭ�{�v=������� �[�Z�5���7���.�ư,�ˎ��iǫ)g��۷�aw���#Eʀ��dbĥ��	Wh./�V��{���φ�[Ɯڜ���nXB�^t	T���W^8�c��^e	�=�a {����ٖj��\����x����nf�ٍf~.lZVV��$g�Pe�a�d�fLKɭ�4���vo����l0<��M�j��zxt�����ydTCʨ�*����lT���K�[[ƽ^htf�G�S�x2�	�îy�ѯ�|r�j�A����'6�9��'�S���>^��1<�J�:wU�VY��xua𷩓���!�Rr��P��^z=X&w�nz��F�,}���.�{AMيv�cs�T�`C��O�E'4O��cj�3�s���E*����){�j�fm.<�:���i/���ԏ }�� Ƿ��\��s�|+0m+�R�76Q�s�g��ȥ���>�/_��~�~���
� ~�KA�r��r}pػ5ҭW��gʸx*�Px.��)�'^+��k�ݧz�P>!�L�q
dC���fdO��c5톼�����X�P����#�k��ofs��݀=�����qx/�-^�7�%����f}��{+Ϭf0Ȇ�.|	��{���kՆ���ô-�0��%.~�}�Ga��;�����v�92���%�=���Of�l�ܝ�	�U��0������(i���h�.�^�g���܂���m��y�ó}�w�r���TP\��Wc����K�z�!X��λW�/����r�׶�/Ѿ�ŉ�Z����x|i�����zK�����Ү���8;������_I�/2�1��s���E{����M 3ʯ=�)T�UvJ���ʯ#v��%,κ�܆����m��U����+����!�_:̸c ܝ.�}�	�i�_k��u�UB�wsVv/�p�޸��0���j��)W�_V��7��P���8�nՠ�H[d_p5@]�s}��E�*��v%I�a��.^�{��Gw�*���`��Z�x�`��*�@-^f�s'hшV�������#�S��+3:z�]�m��}�R�{��:���;�:1�v��x��[n�{��Tk��gc��f�7 LhFf�rf�]@�a�q-��i��f��n�}DFy��E5rP���X"�H�5��{9�0������4!�ed;�'����@ׁ��]�ʠS�6�H�8�
��CA�śk羟A>/�٫�*�1`�K�����^��2��9��������w��Ȁ�m/q񣢯-�,?��4��r�̰�[�^�����Y�'�^n&}n��r!X�K��@�F�����НP�[�u�4��K�Qug�y<h`���$K�K���c�V=!�!����v�6s�l?5,ΐdc�߳[5ʛ�`�.�8�8�kzsj��"�{1l��֋ْ�}�!�n���eX�o|k�!���*�ݏx#��ӭ�ko�7�׫��*�Jϫ���1.a��g��o��8"���q�j���u��]c�u��i�S@h^���+�`P�_!�R�O ���_b^�T.�v�{b�>��W��501�;��ubl5��a�{ѡYƠ~���4�� /�����xV/��e{�g���;|a�{��B��櫑}<�p�dC+�U��΅�ǡA�D��}W�v8Ln��<�x����G�3�Gn����{,d�q��O�Ɩ�(h1�n͵Mv�H}�d5���k)>���p~=��[~璪�3"��pi��<�|x�Z�]]����ڋ�[X�z�9G�V�LI��R�;+�;��p5�����n	N��[w���W�_U?�޻b;��{�߻a�<��/W��~�)H�w��W]}r����r��k']5I���1\��je��9���5z����{0;�2+}��Vػ�ŁYt���2��o|�7�w1#�:�� ���G�a+�v+1�6���Uo(dnM#�RHqP-���s�=�,m17��UzF.U%�`:��p�;����ҽ�e���6�l�d��!��މV�a+uF����Ĵl�P�M�>X����������{�o�	�q�Og�?i���[�hY��5���ˑ��G�v�R��u�H���A]��>~�IA$슍>q{p�K�$�֯p̈́�`-��T���nCSg$��Ǵ)2��h
�����[,wo�V�K��m��eVL5��P�kM�,A}�V:�=3�P��}��ڦiw�տ��z��ІW��*,lW�f�2���;�~N�ɓ�Ϳ�ׇ�sl�K��'v6�&����j�=���xy���i��K��#�ڗ���m�Ni�mݨ�^ ��� ��	*�h/^����\���s�0�շ��G˨��}3iA@r�ˉ��ڮ��E6�`%�s Xy��W7��z�؀��1���wN
��/˼Bޮ�e=�W.��3�_�\&�����;4B��X9߾�����ߦ�i����f�#�gR�5��/�X��a��9�3���S�a���.����u��Q��۴��F�=���	�0E�XjE|4V�y�	F���t,+7�V.}����]���J�����s�ڸv�Ӏz�Έ�^������J�f)�s�n!�����x�[�����'#�0���R���0���R��C�X=e�?����#�V��^8/�-y��]���g5�W�?{.Q}c>��3�P!���΀��0��Sb6ܡ��<�M׳�S��`�E�:��c����3��7��|~�Ǚ^2�b�凌2.���[b��Ƈ���� �s��x8���{:�˵���G�E�����hw����R(6�|r��\ǡ2�^fcM-����Xfk>�X����vnk��K�u`Q��R��q��jtߴ�S�6������o��� #���y
~ز�6l����Y �qV��/ܰ�׏�W3�#ϳ�x�ʰǾ\����U�a��(>���XP�N�X�{�B��+��b�)�Ny�����$�ړ2�h�w<ͮ���TW�ތK�����ƪ��Z^I�ك�t�[L�gA�z�䵪�Sp�c�ƪt&�:�^l�"B�wR�M�����ۤ56�!�jo,Z����|����ڴ�7�/�}�W�}�jc7w��qz�K�/��u��J�ş+%|���T[�"����C(l�
�ǧՏDx�{��	�����<�Z_X/��`�5���JeI����o,���TH���0M���o�H|G5,բ��x�??�/a����s�W�*�O��Q;.t#.��m���K��L��t���+C)X��zJ��j�"�p���]jd��<�L�4�T�o��{W{�/�Vk��C�k[�=]Ж��!�Q&���5ҭW���X
5���RR4Rgvl�{��]U���9��.�̈c{&��Fe��m���a�0�g�Ib�k�گ:�u�=o}��P+,�L"t�U�W�{�������P:�@��H����^�ҭ�>���O�^�<ޮX��~���F�T�T�b�	K��x�6����1�A��1���r��� ��":����K<�}���L^g����̊��=Sm�}G/.��$����nﻵ%m;P��X���݃�O�u��J�ʴ���R�|>���_�\���Pfn"N��%%����`Z�ꩥ�Ը���
���je6�[�乸�}OQ�j�)��rC��a�`l�w��oT��[D%���n]\��\�;�p����B;2#s�Dؗk���V�+���>ߎ>�\��3�.ųE�{x }�������f�.F�^ŋ��%}i�|nv��J	�[=�R��K :G��z��Q���V2��$.Z�b�=�4���f���e\4w�V~X[����B��owr�5�E&N=;���S9v$3�x�j�u�Z*�r��i���p�L�:�n��DC�w��M�"�\唴�ڷ�SJ4x;Z^؀���j^<l��i�'�ڽ�rŇ�ޥ�*�����G�C'k�x����M{���@���GR=�ڌ�So_0�S*Ϯ��V\�n���ĘL�÷�V����S�	m${�����林�h�U��R�7Nh0,�m����3��� X��B�9;���e��.�y�e�ۥ�x��ѯC�]Ƿ�����&v�m�����ѭgw.ܾ�br���|���i�Cb�ީAz��嫇CǎD#b����n��ѣ;�KZ9�ǌ�����Gu��;�˒�;za:�nf؎	]גܳ������ˠ�(���3s+!��xuA��5®p[�{J��4
�3����vMv�Pfl�
\At���{<+ǝ@&Ğf�Q�S�ϓH�2��Wg�Z��ƣ������
�ݵ2�>���40g_<p�ھW�MB�I v��`j!ׇCԭS8�p��Y�u�k$��G�W�׶�e�V�D��J�Y��d�r���b��
�:8�b,���̬��O�-o�bb��$U+T���,#��Hї�e�ϟca�p���y������8m��W1�T���zhX��Ģ�ySV���Zo/�GҸ1�]�x+/��e��ήfw����
�&���S-�Ε�Q?jF���A��Pw�ash`�T�!q]���3)-㲠?<��LT7����RPl�5��1ڴ�Ú-�S�Wq3G��3I1J�e]A]>7�7R,�Z�K�[��;4_*u�S6�5p^�s0Z�oi��hT���"�A2�����a.9o.ȫjeer��+<�a�+8���p�S��?K��2t� �ܯ�� ����#Ygv�L�9L�]��3����LݺnM��U���9W[��F^Ayy)u��u��r�1ݺ�V���éa��Ҩ�֦���k�h�*e3�qnTP&([T����N�ז��u�T����9.L���WNo�L�[��ή�j��7N5k��].��Ҥ�n����X7��`�<�RCro�뽣�g�_:�j��;t�8�]>�c)Adk̻ie�=8P�a1q�C7��(�8J2�[�]�ۭ���Bi�$j������.�5Rh�)����霦,�GWLPn��7mJ;)���Z�Un��R[�]�]�9+:�/�4�R�Dm*�X�Q�E���QV
怡XV0�FAW4Ab�m-�,�*�,�U@TMj�Z*�Xf�U�m�"�`T�9��a*��Jɚ�U�#�ҁQb�[b�"�[-J�V�b�Q��KhT�m��Y�E�]T�*�T]eF$E��2�0X
6�Ub
�E ��fL�U�*PUs&L�ED����A,P��#"��0�
V[e]C(ᕊ
DkYE
*d**�(,���ҤX����B�*H�QUI���TH�� ��U�,Pb�* ��F#P̆)R,E�*Q��
 ����+X[E��]J¤ib��9#,YZʒ�R�(�UL�UVd�(��dY3 �-,UTJ5��mE�"*%+Ϝ��*.����H��'������G���utM��ҪC[ϯf�B������[����:5�So� 6O�������o�׳���^�����f���>>u�¸><��I`>��X�iWᾼpw�7K-LQ�S��*w����}�+���������a�UvJ������,�*��7P��S�k<�y�7OЏ���1���X�g����L1'd����.tb�ڟ�`�ۛp��ҽ�Ϫ���ly�֫�����X�����j�d�\[Y|i��3��6�x���Y���4@�_�6)�}��O�>:>�������eq����<z_��J�3���{3vg?z�Q���T�C6�e� �_?z}/�٪��v��|qj���}�[Gq6�:g=�o]T�ړ�+���^�<�xVKl�HN>A?�u���z��f���{�f˞�;��agd%7��`mCw�LR�n�g`�u��^p���]V�[����XB���Q�j��C�>��B��5���3� (�w�"�q:�Lg�eRy���ߥ�W�r���z����ʰ�K�F��<�m�1q�%��01?7T��*�������q~!�zs�2|�R}�g����*�̽�|��,����o4��֛�	WD�[��X R�&�×���qv�t�W]z8�����l��T|9��}�6rD/_n���[�Y����\S�e��x�Iؔ=�3���[�����o���S:�6z>ݬ��������~����t�G7ߞ=x~bp<"/���D,��ByV-�˶�
{a��/k2ϧ���k��ȍ>X�\W��Y�Cw�g���.n�VO*�ޞ��'·�q���rC=G}OU���C��W���}�s��*a�W��Dz��Â��c/}�{����.��w^�^��Z��
�S/NI����CK�Р�W�~ WQ�ExS�����[ݫ	*��*���_��?!�����Â�����ܹЂ7��݅�S^M�7t�E�q�C���2�TyM
�\�1��� ��7~Y��߫D,�(�:���#F���e�{T���2���EY�t؃�q��\�W��Ta�=�Ҕ!tǎ�J;��uS�`M�^��[�^�A�ee �����\Ɔ"�Gg¶��kb��{}�c�w�s��9���%�Owi����㌌������@V:�ll���ԫ��.�/q�W��tk�p1����O-�^u�z�T�p���"~5]��k���mR���б�/+B�AF���}^�{�yz��g���tfW�p*�[V<o2�[������B�������r_V'b�0��f�c�)D�k����uij����BM�uy�R�Օ��Ko%pem�t�6ŵNj�n���fc�V�N�^>ꓷ)�Ӭ�V�����v˾����E�to,	���}��}E�~��e����O�P�8�u�u=�D:r�u�C܉�F�ϕ�kn�rV�����c�4�����b&7e��rkM�T� ��o.S��[_Z�����~��B�Kwycj|�n\�<��:�؆�����uG:��?�xs�V\��%Bs�_��v6-��j �ۅ^����fc���U@��<����U�an�x��e=�_ ���+w'�u��I��^o���{���k���(��7�N��@�O����V	hm����*��'���:�&��L�ru^gf}�r�/��̬�U<�G�q�ck�_��Ν~�od�ˬIlڡ�"�ƨɇ�cU:���^�f� �yϰ�~�ڞ�?6�d|c�,�,,�p�ߗ��Hx��ܿ��j���9P��뉖f�9�kƱ�XA��<w9q�Yz��Lc�����y֧�g��[��{�V͊�=��xl�N�8`kc���*�^�n��MB,-���!W	,��{�N�
n��2˝uwz�S2���`9.m����}�RZbK~9&�u�0pB�p�MבȲ�.fA@t�h�Z����!���]Y+�i:�v�w�D}��}������7td�D-�t]i��Gg:#��'���5���q5����p�f�z��g�u,�O��Jw����2�umϱ�UO�t��|�v�����u�&"}~�(�C}O��!�Ow��Y^���\#��ݵ~�L4U�g���X��c/ӓF|ӹ-|ק�^i}e�TB�!�W�j���[n���l��Fj\a~�C�U긣Y�&Ѵ�Y�PqKx=IW��@�.N��(|ʻ�e�������t�U?SYw+�q�����L(��e����+��i������oz�<��*���}q���S��1��f�ES��?dڿT��+sWB��[�\��s�*�tt>K�k���^ͯ�,�e��F�ڈ�s�dK^���4c�{n
�izt����,��ŀ�X^�Q�^��n����]C#w~nq��]��j7��wiP��s>q4��EQ�h/cZH^/$��=�']�n�´��m	
+36�>�)�eݩ����'�+��h#���B.{�3)�x��4�l�$C�Q�#<)_]9ݱ����λS�N��Pǽ8��<�]V��#�5�k���`�<e�[�J@b˩�[s�">�菦go��ǎ/��!1�ǥ=`�mG����m{��d5�`�:�����W��~�mtEU{�x�X���^��*u��I��Ь�5z�>��ճFhP�1�)�"�դU�O�y^��j-(�y��I<U0�%X�Y:�7����R�#��W����Χ�9�D/i��9m?m�~��E\��&�p5ɏVyv��3޳�+�K����U�m8s_��|;JV1ӵ>�"�K�x��kS�t��w6y�kЎf����{���U�T�Pt
le���}�O&a>�'x��v�O�R�4��e�l��P��y���L(�C#ޞ�u�fh����V����ͨ�Q��*���R�m�c����F6m����gۇh>D�{�mQ�%	�.��sOW�����i9rN6P̺�.��Z���՛�#YЗW���U�Oz♝&*>�0gsUռ1�K���g�7U��W���	n���Q�B_Q�r��s\'-�.ϒ���l����Ja:=���V]�/�;�>|&�����|b�o
'�:��kN��J�3��y}�����BV���d��V�]m��V��{��U}_WޙⳲ{˳`h]�cmP�rba�-�c_�#*2~�����O2��uam9N�NӼj7�p���k���6����L�A���s��^N@H�/g���O7/=�Z�d��\��|�θ�Q[��'橒v��1�qW�̜�1�/�(�Ԯ�@�Urfc8��Av�����
�����č��:~�g�X��Y�[]���̄��=��6��n���L:nrP�t%�{vߚmɝiY>�F�8��3�,ݻx�Fʉ�<qN�N�ź����o�׆�O�߻��ڨ�=��5첸^���'��/ky2���	�v�9n5D�Ð�kƢ1�;�t����{%y]��R�Z��US3��f40N�5����S�7C���ݝ8Lj��Av�7	�k솦
�p��^T�-��u�����"ȴ���{�����	�u1�V�JM��'�m�D�"��m-:h� <���鞓�ǈ�o�Gʘ{]��g;�{=~"�7��z��/�\^p[�\����Z�a�wŃ�>&�7W6���|����[�,{��S=�-��:�"`�+�r���2��8�M�dG���j�lُ4Nag興��ηW��t��VD�MdU֪���$Ss�]�>�'�c>\t�4�N��w�.�n醷v��uv:ש�]?��=�N��ڞ��kM���t��"��5�W�M�*M��W3�á�ߎ�G�4��_�y#�{�s��+�s�z�xpUC��Ȯ��m�:�oޚ�z"��Ν!�]`��^Em�Ӄ����j�-؉V�5E��1Q�K��e[����t����8�y7���T�;����nN��\-�nV3Xk' eRB�ͬ�=�,̓:���6����߬+����9����tFU �F����-d��.��=\��1Ļ[��|3��ɗ�P_����D̄w�.��}/طj�	U��m\����&^��Y��^^b1�K`-� a�̑V�}��KX�Udjӭ������J��垹���}�"��o8��y�(� ��H�x�n�p��kՐr�[2j��D
�.���]v�hP��u�ŻW��a�K-�������ͦ�R�Ϻ��X��k4̴��K�N3ڲ�p� ��Ȇ��+��d�MFo���l4h�U8S�΀�L6��aS�u��tÈ�P
G��}��U_W9I�ۦj�v\��\kb^�'�Q���W�'|��m����A'���]�#����>�S�������Y���ڞA��*��Su��m����s�{c��j�!{~]]��������]<^Q��{jvs]>�r�ڏ<r�A�
ڜ��6�\�X]�G���^̪|��;��c��,�~�+�A�a��9o>�Y.k��i�*���GO{ݯ��4{�Zߚ~>�KFL.9�{Wa��~��3뒢/Mex�g����Q����yk�J�M�:�[{�n׹���{��k��u^�۪m93��s�+} �qI����<���g���z��UY��T,ofԩ<'(S�#�ڦ_nz���?�Bj�����U���N�¹��nSwO2�#}�;N�ޣ�O�~��e[<��d��^~߂ɴ	8�h�Ʈ�����"��i�i����N1���EL<-����,��LI�I8�w�u��/]�y�x{2�M5{c޹�����n�֖s�F�r�@��C�p��G^�He����X1��>��mrv��:�"�N��Q}�@��~Oq��":<щ��[_<�-կ��)��do��n5;���zĻGrO���K���|=��U�B�S06 ��׃�Ø��yg�s=�")S���}�^f�E%h�-��Ge����{��k���������$�gH���@��9����
s^p]ǜ㿙�ߛ@g�^�j���ه��+�w�$�(�B�º7�n3X3��[�J2���ם������m�u�4TT�g�gr!'�IbߗR���Tά���O����*xt�D�r��^t}�a��s��"�"��m�������WR�~+��>����+�줋��<=4���|���ؕÝK�n*!{O�v���˂���ښ����bž�{��ܧ���O/�.[ag�PU���:�|��ۃF�_���W���3��/kʦ5��g��fv�!�[^�\;k�5�5�C�g�6�]��b����u�o��e�\��yQۯ����I�t����Y����S(�n��Z�ҕ����GT�T��ߺ�|o��t�.P��n�����=�3�ۚ��ORz/����ϷE�\]�>9�}��S�}W4�	�RR��V\NQ����舅�~[�w�W1�֝�����-�Os~mǩe�p<���B.�����q�K}ۊ��J��T{��w��oiG���n���-�M��4�x4�\���u��J�5�ô#Y�?��io���ߧ���7x��u{�[�|g�z.ϓ�*�)X!���K>�6���3 '�{��=^�j.��f#ՙ�?{��6���kГ�Q�J�S�P�}�5��*2b�a�������W�V�ݫ5�v�3���ק�O��v�h���@��0��'�וpa�6�8V\�����:,{�y��*`Sbg�q���
b�d��=�-����O���"Ip����"�\�eR�f�ZT�E�b�]�y���^�W�c.�~�g���_�>~���q�ޯ�����HQ1i����wF�ҿ$�$S��|�����.-�?#�I� ����gT��)���gvT�R�A�57��v�k�XB��i���q�V�ٶF�y���\b�:�vl4�@![����t�+������OE�Ꚋ���Ƥ�HN\�2���
ڒA�uh�@�$�N'��$�s[K��K��sz�� b��.Q�琷YO ��J�G�f'ݺ��+���]���]ܮ�<{U��g�m�Y��a�!�
Ja+��݋�Z��}][�����V����oDd���x�۩\9�����,�Ղ�*SB��kI�Ŕ�֬�V��0R��V��}à��zF_S:�rk�5�-��NS�^>l��ֺ6�i��d�w: ��2���3$s����Vo�w��~Cx_ךL��a�j9���E����W�ov�3Fij�|�Uչ���r���4�k-_\�X(�;�P�p	��u��*ؼ�5�*	{ԝ5�^�[x�V�m��'DJJ�@q���[KQ݂u�'�p���n���ݖ��)�<��A�QBx�l��Z�И6�&�"�� �)ػj::���W\�B������jAɌ7Koӓf�H��nҼXk���JI 
��p��`�v�$ d���c2��=�6z��/��锯tsrd�vr(8�f���x5ڸ���W)��ڰ�Y�K�yF:%|FVM=:ԡ=��'
�T�u]���'��<�-v$j��e:a�nԱ�����p���s�8m���F�g�<��z��-��{����c&��_�x�6��ѱ�a�{9�Hs�y�wEra����M�W��r:����i�+�xF/^�]g�z����d<��]_L�1w-�s&u�1��.��s�h�7h�4.jh��-�C�r�L7�%������)5:�Mҋ��%���\��=H�F�1B+Ubd����iV��O�"���6���Ԛ~�}�����wc�o4lZ;�O��rbB<�w�|���@��[k`͉�ω�G[���KGfd��T�ZŔ�Aʒ[�#�я��|s����oth��D���}�;�����6����+Y"i���[kihMxnI�M,�Iך7kY�-��L�������
[�nhNu"��
���o����4l���ָG�n��3@���4�@��r�lb�,E;��BsH|�Z��V/F$:�e�ZN�AX��Y�I㕳��k�l�\�Y���%�rX��d�Jj��hBk��.gS���ձ�KD�9����yv��]ҍ�X�.��WN#y��*��)�Y}ԸPN���Z��`ٳ2�N�io]_ ���yG�s�/k.r��Kv�4���Cs�k�¨�ڨ��(f���X�I�0����B�1bI9m�@-�Y�/��L���nk��ّ+k�������N�q7�rt�sR�^`�ܳE�(��;���ue�Nu�t�`-��J�Aed��h�[
�a�Vf@b*��`"�(

*�m
Ԋ,F �b��
Զ�E�-��E��X�r��L�((�`jڢ]�@R

���f)F0S$��ebđ�X	**��(��%a����QEZ�`�Qe�J��0GZ
"�DR(�Zڋ*(-c�F,Z�Mh�H��F,�b��(�#"��H�R��c�n���)A@A�
�*�AaR�iX#X�(��R�5�����,Y0�WR�mE�E�Ֆؖ�2d���V���Q��U�Z�dQ�U@m%���0U�k*����	j��FUGZ��
0V-�[rfU�IQk�"1E" �ut�@�����3T�_v=$}C�"��h]�v��D����}���uZ��fzҫ|�:uS�f�t-��ϰ|���'����}U^�⧻'�mpU��c��X��r���>�+f0w�_#1��� ���#�{�;���yS;k�cⷽ��v��ս��7�M�Y�Y\��ua��
�7])��N��}])�i�-������^��i�	�J��v%r
�։�����vE����z���TGO;��~ܨ�z��Rs
k�p���:ؘ�㛗�i I�X��#q�&)����U����IWϷ(�4{��`X:� �wcv���jn��D����87wW���+\����}G}�U7�% y���~���R^��U�߽Q[���[xcU�����|��@Ϻ��\(����-�VL����k�[�Ɋt�Br�\a�����V�z��q�:F;<8��y�)��O/�z1���m�$��WQ�LO��5A_s"���W�o����p�0���%��y��w>~trv�&�N5�	\����4��u	&%�)�	}�r�gQa�<���*�FJ�ix��g�.�%��H�����ј=,=���W���Y2��J��څ�b���R��rދ���jf͏����{!��.����#K:��遧�K��\7���R'��t5�kn�3����i�|��f:�~�����\|[������Q���O����
�퐽�'kE8������&��W��Xέ��S�J�T/5^��Rar�:~Y2� �\�NLŝw�yt�]����k+��2��^��o�	.)y��cz��v�ɳϪ�\�R���r�4D2�@o/�D���^�>wF���'3Z����q�u�����p2���UV�|=�ef�y��a�^ˋ{5x���0�^��z�`]�,[KԻ_RʝG]8������j3�ғgv��!zeXt�n�����\�U��B���8�1Fv�Z��������I��{@l�2�����;�ڒ��~���l�������G�c��������V؛�����O���y��ļ֖����w���	�B�zf�D�:x�=����}�"�ۀ�Ӵ�sw��SN�޻�m�����P{���k�ƕ:]Z�v��;=M7�![LM�F�2����F���k|>&�P�/_x���-�u3l�.µ�~�/Ǌ/�ToiM��Z���Ƽv��[�z�����W.�v�L��fԻ�B�9C�2�ź&�ӫ��k�y��\5����*r*���J彾|����*��j�y�:��<��\�y�����
��"">-��)��d�e.�=�'���z��r4%�Xn����Q�;W��G�?Y��$��ud�NW��=�~,����?+�.�+��	LXQN�	���Rw�jޮ��7�������>��������=z�[U��!9�0�w~^��X��q���67�uJ��^��mݎ�|���Y6�����}���{<��3͇`���yL���+ҽsɭ�����=��+���p��Rf���ە�t{5�6:o�OW�Y�®W��1�^�~:���؏�K�1X��/d��v�כ���c\k���w\	����P����-:\0�{ۘ�C�M�^�<�j�F��c���v�=�L�5x˸q綻�7���p��K�u��u�������?NKwQ�Ϛ�����V�����6�w�-���?+E�U%�~]KϪ����=��o�w�i�h�x�{M5�_<�5&:���5֩\�[��_u"Dn�/Qx�;�]��Yc�|�`�W�y�Z�|�a���[���I_vC��o^9|�9B{.Jw�ٽ�EH,Ӎ�&9o�*���80l����Y߾����������cw?Tj�Cm>�*v^������y���g���R6�È�~Y/�F�{���<~�p���D�3]�\5�K*�q͢���v��~�����VCY2u{����y��8nw��O>��	<�v���g����W�l��tn�N�jRm_�o�I�9�Qt�z�n�yܜ�F'Wgw�����J���y��5��,�����O}ITym�{���B�n��^�� ~�1yY���<2Q�}qW���߃�Zvxm�s��\]u>hM˭ـ��u����W���b�fH��u]W��|���6���o��t�R\��ݣ�ֿk����
b���М�Wa��.M�yv)nf��^G�nB��j�h,G6��Z_���¦h�ѧLL9p��w��kO S̐{����~��w�~�w1��N�h�덦�&)S1Gal9א<�
��H}l���_Gz�]�$6��N������ݛQ��R
h���)L�M�*�� �u�ƼN���a��"to�����h'�6kv�W_g\͎3o3��5ShQ}��s뚳/�c��f���t�Υ"��4����׵�0Ҷ�-�ڷ�F��c��J��s���H�Dgu��"N�����e�$%�r\n��=�뀮cd/0omƻ��p%zn�5��L:��3���<�j*5 f�¯y\fx�c�q<�d)����e���ӱ.�^����j<�L�k�T�͉�?\|s1�g{����-�
��ub��Ɍ�Dh�ͯU���R��������%�Wy���_�43����s�c;�z[��o�Y��w�m�һ;寏�M�pgK=�����YtS�}�S�����^��k�[ک�y"����N�2�S��p��'�/�9/�:�k����dF�F�<W��i�	�J���ƽ��P�|\Y|I���!VD���՜ue��K���t�����D�}�v��e�~���w�=�un�#�p~��.uz��q�J��b�ik�jox�A��{�-�/�3[5~!��uP���j⼮2.���Kj�p_r�Dk=i����^jXJ�����hr�0f:3��%R,�XlŸ��;�h�ՍM�4*��Cn0���Pi3�	�̘�B����j��b��kJ�,��BN�5��2}�h����U��vٗүvX�g?�����'�M�Scٽ���k�T9n�����C�ɡ�q�t��؇������+f��,�i�KޝXտ�(�|�*��]΅��j�L+���>�9=���� ���ܜo~�yTj���J�v&ʘ�j3!�N���R��my��
验�o.�x+�?:�g�5�&��N6�n�<;2e]CW���]b���Â���s��U�V�N�es�;k<��V�S��+�8u6bԴ�&��	��������J�c佭�����t�������+|2�h�o3���D��%j4�_#p������?����q�l\P<�O^��`7��ګ�d(��]|�㰎��3�qo����	Իٶ� \�&�sb���c_P����z�S�^>�i�Z�}��C����ջ~e���ve�r��N��Ib��^}EN�=����>>�f����m�nb��U���ۊ�hXKV�m�r۴�آ�E3�4up�&/��i��:7q� �$��%cV
�ol~����Q}�p��-ˡ���������E��[�}�r���fNjAR����DB�u>�l����8�Ʃ��h]��Qβ��FAxJYE,���䶭�W�r�w�~������.N�z���e���{l�<�MDY�X�}���(��ꦝg�W�o���w��w��V���F����<Ū����8}�������(�k�sH��#��W����֏Ӑ��������ӭ?��uo�����	�]�heT��?�������)9������{��6Vx�RJ��;�������o����������mS�F~^��n��K%��션��%eM���g���3D�EZw�t�Y힓~S���9HNP
�m��O�S�m�(�MD�f?`9A�&��ߏ<�Jh\���p�{�,TB٠�r����?0f]z6�p��V��[K}㵝	���߷�<�lZ�=TǦ��U&�T�М-J
��:�W�]G�*��Oް��2pj�2<m��]O��Xlw���О��m*���N�׵�����z;8*��S��e��r�fk	yb��)ϯ��ev_E]��_5\�\F�VkB�[�sX�	����E̝AՅq����NVe�2��ԜЦB�=�TƬ�]
�z�]"r�umoҮq��os�~�������А�g�d�:��'��;-�q-�$҇��c�VMh��{M	�8p��녌��s�ڥZC���nq�WT��:�NEGh`�ϳ�:Y^�k��+�n�e��l�1A���iBa�>�\E�Y^����/7=V�nc��a�������~��-�Խ�O�L�ϟ��}y����S��{�����fŵ��³k�Y�6ӯe�v����V:]K����@��/9-�'��Xk�WM�v���ڲ��|����ܨɅ���4�����VS-�V;�7F,��VW�T��jS�z��o�1��x�Ѷ��R��B=�?B3#ڞ/�=��*�P[�{_�[U:�o��i���澅t?y�qY|�c����9;���|�G�f��Yw����)o��i�T6�[/��+:�����ng�T�"�~�V��N����m�{���ߩG�������u��"9Khm���C�����N(�qW35M��Lr��A��_��M�&��Y>�ϼ�u�n����#f�׹jm�]]�P'C��W:�Z[�%�\��\J���6�m�woEf��6��ɸ�pe���s���d�
�ΈY��_W�U1ܗ�{Ч�+G���=�P��R����7��������S|�ԋ��W�U�͌�͡��˔[(�a��1���9E���1�Ǩ��;��hm��[U�����N5�n�+F��0ǟ�2��:�ߞ�x.�����0J|O��������M)§�b%S1Ga+W�S����{){3�Oy�*r����w!y�F��G\:�*�֣bF�Y;p�a�s=$Vus�1ī����f#?b{�+ S^p^FJ��+ҶY�yt깴����{��3�_�L���'Β�ߝ��)罛�\��G=�}��u�!���MNM|�]C�'�NF�9�˃��.ջ�a�/A?N"�n�}���D�zd��e:~~�z'��r���|[U�������x�V��Cq׹ x���K��>���S����>5�/6�ս��6kؐݨ�B;���V2�S�z�S��b\���{���F��v���w3�r�f�aM)]���?�e\�:;����F��>���Z�v	�+�*`"�o��we(Ű�pl��	�#��НVe�w�����aQVnNd=�ֽ&�#;`b�?���ܒO{�r{�?|�d���Q��^W���F��m/R��ޚ*6���	~c������6�R��zf��j���}��~���%q�@�ǖ}];J�d{���>V�0�{���u���p3Ux�D��:x�=�ߟi�<{7�]ߓ���t/A��ϭj����y�Wc�{J��]:�|]T�� ǩI����瀏p��w�?z)KԲ����iJ�-_���ڛ�呙)$�F���O��EI��u���?{V=X-�N��)ӕ��g�'��<pL�go���Gŗ{q>w>��+�Uq���z�(j��w�vVm�2�p����=3�Pz���]���k(��F�7]U����W{��w�=(�<��}�ݻ��4:�.���
���P~N�m<�<�m�f���/��o�u�$ K�����y
���9��ʻ�1�a����=��Ŏk�<q�!ϣ 
v�~��af�y9�ݽ���v����O��U� -U�Z{��z�*"3�:Q\����;Uj�X���W*خ�ꆸ�Ka���zR�FST)i�mv�Y�˚�4�Vmt�|sF�� ��A�$r����=�Pr�%��t�YWf����ie,d��P��9I��X�0�(u�JV�w��{pGu/�rq�����L��Dd�K�v�mY�(@�b��Q������͘�Bj��o�����LJ�����>}�Fv�d�6'Ck�3E��tq��e_CFa
�ԅ��3%f�����n�W���㙗m�Gp>����c� �ܮf���r����r��JT�If�ry�6�
X�+l�è3�����1�#�}{y��^�I溳;c�պh��=����WJ�v�oR/��u�^r=(ovV�|^���Jg��5ٽ�U��b��wHMZ	�����N�Q�{9�Yh��r�jܓ�1}�-��Y9�7��en2�liy:��>��2�7u%����0ʅԫ�om�!��\wDZw+h1�p��v*�e��W�m���e
�@�\��ζ�v�Suc�����.�J:x4lw�t�ā���71���w0�sr�=+_=�<������n����}�J5��*��e������@�r敻X�a� �{h����PF�L�\�T�����PvQ��3u{��;.ۘ��Pԛ(MGze�3;�މ�x��k�uz�+%���oBj���*g9>�(YK�6�v�#���n-�%e^��(��@\���jJ�0%·&Jh��073H�zҚ�ޮ6�pmZ��������: ɕ�#��;.da�dMͭ����\��-��v���]�ջֳG�H��[��K�"�J분��Uֱ��	l]ip؍q��r�i'H����u���6*'C�0�RE)���򒴯��
��Wa�%���#��Y�]�OGc�Oju1`�]� *��<�l��u��t%�+��;͡L��)�ڶ�����O{:�}N�Ce)+]n�� �0C�]eN�MT:�ù�JS�\����)*|��[�T_�h_%��K쭓�y+s����JxD��U:�8��tJ�3BN4�B���x6�t�Wua�(�u���T�Ĥ����]��rD7h�K�d J'�)�$��Vp��ͧN�[s0��^n����i*�RJ�q�X�F�7"1�M�.�m���[�9�.�"��;���d���JC���!�k����M,��n���苣ɹ%%��L�4�K�z�pu���4J�O3Ze���k�r_]faF�ms�=I��+^ʍ����Sy챘��!6�l��l��׎�-��z�9����5����=�%�tŌ���{z�)7�k��إ3>��Ve���S��p��Hg@�5c�y�@eAͪ�B����wQ`t�j�e�r��-�+�3rSl�K�kh.2�5�T�E�wwTo$[ѝ�c�0�Y�
]/D����֌�j��z��t����J*�F�`ҔV(��F�j[b��/��k*�b0QDE�cmaZ�T0C9�X(�)[d*�&�TAE�U���őK�E���b$��B���E*L�m,\�XfJ�b��((*(�X��
��PQ�*���V��b�C0**�,T�"!Z�m��j��Eb#�R�ڎ�2�Qb�1R#(�
��#�
,���+E�m�DFA2TR1QeJ��Z!��:��UJ�eJ�Qb�+A`,��mGZ��dF,3XA���J�6��d5|�W=�#͍�yt����N��_u���:���[�d(p�Ɏwa���pwڬf�ݼ�K�,�)�E�q����,�f���}��Y�R63@��
��	���:�q e{�ќ��?PIqK�9P`h�P���{7F<(�۟��j4���M�;
��-��Ϟz�0�0�zf��1��u��nW"�|���}Bg���l|=�OD���=,4��;J �V����#��{؁ڋ_�j�/k�Y��C�	=W��ɝܝ�4�U�F'O�X�V�/չc2V�/|��1=�}Wΰ�k�N���
ݻm-�x}��L~\�~"J䯸�^Į���v���G�;�>�pV���2W�V{Y��N��O?�jfrs�҇�k�k*���s����L־4.�ߝ���^�f�v�b��q��L[��dRN�޹���z���PV�s7��~��̞��FN�-���B��I'{��)��GB�N���T��~��oZkE	K}Sp���U�{�~=�h��=&���+Լs�O��8�]����gU���H�+^�����Ӿ���,9���w=H���U��W ��vi�ʔݪMakO�;�ƽ�j����;YS�UD��}�oc��F0����2Fv�q��+;�Jݘ�S��^�r�+��1pݧߪ�﩯j�oyiǝ.��V�y�T"oz�<�Bm.y^W1�WY�onzN��+S��v��xW�j��5�Uo���蒫�co܎��WB�Mo��vKN ^�RN[���������1�וWЫ�����!�o��B\��3��2~��M8�?N�Y�z��^�X���.[x���'���'٪_�ܝ��5��N5��n¸���R��y�Ue�-�{�B�'����+��ɻ�*K���e:�e均��~��vA���������y�U�j��eib�]�����M��^e��Z�
L�E�x0�g{���8�#��l4}�ױ�<���أG��	����K�j�q)�P�Cr�����xT�m�����*���'�K�u��u��ڐx��<�f��J���]��){C|��}�\9ԕu�T�Oݯ	�����Y�\UG E�ډn��wn5�*��N�u��m��;��=�[ۊ�}�y��`���2?m�pk�����}*,V#��q<*\��"���IE��߄�o��o`f����������j��9z '��k�Y��n�,�".r����n�d�}DJ�ZZ�d�)>��u/<�5j5)��~Z������-��T�Z���"�oޞő�]z��y�C���w�nT�����B���M�-��x&Uډց&�c���\O��E֯}e'~���-��O}p���	��K���>}��{�W�&z��{�~&��sٹ6��[Gg��e8���5��Fr�I�fl��:�Sm(�j��nU����	�n�>D���t��`38;���s��U_�z����W��)�4ܲ�0�Co'�`8=�v���y��;�<��^8	Ͻ�G��p�-ؘW*b���
�~�.��׏p��Rٷ�s4=�s@�<��;��w'h&��
���X�K���r��9��am_z�y�e�Tɱ�����9��ʞ�랯Zoi�^�<���Mf��Rm��W��I����|��S/��/�
�k[�i�^����:�w�K���û*���ލ;}��@��L�7h�Ĝf�P�n�'�J��b�8���]�RUٞ����.�0z��oօ��!����h��-�P��{�n^�;!��1]��Kijy�u�/�3w���v�K;Yg�}_}���'�
�-�W\/�Q���~�����K�/�_���u.�=�H�ݙ��{�K�*������795e��^:�\[U�~D$����^e��ɫ-��ȝ�3Eƨ.v&<��F�P�y5�xw�m�^�+k����c�6�㢳�
�Ow$�W��c�󌟽��ٯ�4�iz�ս��6;|`i"D;����S�7�5��K���Y�_b�U/*#��F�S�m�ܭ�pCY`�9^�����tkԹ[��%p��Uˎm�dzq�;��b���g���x=/-i{��LZ�\/S��j��M�*ɳp55VW�*�gi<^�)כ.�����}��{�J�������� %�5�ydUֲ�U�Q�*�U�J�2�ӝ�8��I��ߓܥ���w�KGl��^��f�a�Z�>�{����zP�gq'+�S_��{�o���֯5�/������	T|1�MV7^b��!���o���ջ�+���g���w���n�ZG��b�o_�T;��L7��K�e����Ѿ�D��4#�6
��V��s��u�y��+�r1�q޲k����z�B U�*�VU9]h!�s��ّ���Vvf�6���l�h��}��7��[�\̅u�o�-�Y��]���~�����J��o��*N�id�Eq�7�z�Q�5��/��j��?z�����g���w��C{1������<��c*{���*�y�������f��uھ�}�R0P��g��L�ѣ٬^�ۅ.�AMܘ����L�{7�T�{:�xO\$5�}SU�gVu�]҆�
��K��i>�ޖ�F�-\��������,.@��j�}�(���~u��o��M�욭�_���9��TZ�/��%�iNc_P�/y֙�nq��KN��pc�����X��ْw�����]��ױ��Z��)uc�ϵA�]8����5��t��(�cw<��y\p"��m��Z�H^]G�[���ߞyWq�X��ov��l{�j\}�7�$�J���+��k�n*�m��g,MĽ��*;-�v���a�QP�Ր��l-���|)���z��~���z��#�S��Ҍ˖1�̿��I�(yg���<W6�wP;�e�߇	��v8^�����;�v�J�7���]��Y�+����#��['�Ź�0�|������U���f�{��2�����;*ch�9	s���y{�f����߸�\��m�绢��L�Uğ�/)ϭ�o�&�y1�W��A(X�c��׾�2'��{ �w��%��t�}Ϥ��ѯu)���1ܑpI�}��|�� I��ǲ�M�,����}ijL�������G��,�������WN�,&�a��B��V�����7��y�ՙ��g5����5�-��ظ=�����r�n8�U�d����]������PY����ʿT7����)Q�z=)8Un²����5��2�&"�a�.�}�KޖC-i���Iҳ��/�g�O_���rv��tu����M*f*�ڀg�2��<��tZ.w��}��w3��u���+���M���r�����a��pU��3K�����FK��|����Tiac��6�iVfxM&(ØŠ�;:���g�g��f�
�q�pk:��w-pO����J�+���]�oR���هB��+z����rW�)�������8ȫ(Գ���w�ͻ�hϸ�$�$bˆ�N˭������ɹ�o�]��2W�����W�z>s��ѭ=�@L��k�>~�9���̜�L�P}-�{gW���ʢ�	�f�ѳN�����{ߪM��@K���c�?��.��}\�;y���y������|�>�l���b:�X̕�%� ��KS�a��!G��ooS^;j2�^?���{��Z�aM{�w�����P�pmĨ�!i׳R�ث�Z�YQ����b[�U�~~ܩӆ�w����i�	�g{��5S��q@
:�o�����W��o�uXz�-_G�OۏR�M9��6dL*Q�<�K���������ǫ�ֽ��ʴ��Gw�����:�����SX����Q{�$���Oh�v�&��v��\��:*9<Ǻm�yܵ޵�lZ��p�����T9l�+�K�g6"G��`RҼ���^���v�{,��Sa{�����H�Cl*�0�U���V���j0CUu-��e�
��T���w0{���*����g��D�2�(g�^ƨ���y�J=ţ�M��Ķg� �,�˼��®�i:��O�%��
��j��.)��{��e-��]���s+-n�f=	��<��m)һk��7;^�
���{�?W�_<Mn��M��
Ǚ��{��q���F��T=�����FSǞ����0���8�����d*��b#rv�&�О�����-:y�ʴ�w�M��M�B�=Q���9��M&�S��j���/����P-z�:��fY�����	��6�n�}+�|>����˕���ɗҲ}>��;�z�k�zPC����v���QF��/\L��2��3�Q��K��n.A����ǚ���������a�Cr�����B��xs4�����W/���z?o�����wsNP�gV?V���^egx��h�,�*.�eMˁ��',�unz�]�f�c�~q~Q�,��o�>u�/<=^qe;��*�{�-�<֠�$�p�+g��/,x����9_�S�N�o�uk��{�WC��(�Ӟ�c�����s�J����\�h���:1ݴ��=I�*��W��=�i[��Wܶ+�Ԛ�)eh3ڢ�ZG�zd6Ǩc{/=Mu;7!u����KϚ�/lQ걄��e�[��pɜ��C�3x�%������_Q�º�wwx0����դ�Z�%+�d�X�}��}U�W�z��^�s�<�SSK=��D����0��Ǖi3�����#I���C'b�
UMf#���z����j��W��:�s6�񧓯h���=�x�!+$�:�J�V�G��\F8�n���R�0�50�^��K^�B�o�Nˈ/r+��E���+_�:V5�,ĺF�9R�NK�^�T�x�vg!�nk�{,,;-{ۊۺ�[si���}��z�(kG�k����#ŬV�[3"n��l%P0yz�3}�k�v�eS��2����Е��9��Y%T�5h�R�(�%Aֿdz�'O!������5k��(�jm�^w�{j�Ƹ~�b�b��������u�;���gS�\~�ѹ�z?{�a�ِ�}�B����l�p����?f��<�д�q!�9
lٿ'��^�[T�HQ1u�;���<��݊m�D?fW,�gQ8��D;h%���7.�R�Y�"�W\�\�;G�޾~0���m�A�() 9�;���J3�еz�\�-��\����ݰ�����b��X��\XW��9|�1R��VPy�8_R�X��������<3oR�y�k()�E+1
R+Nw�}g6mo�E���q	.)b��1�>�=�U/S��y���.���G��:k-7�]��~�w���\��c|��OQ�}K>�F5Ӂ��~�o�[�jw����o�y��7�r��{,�}�r�k�!{iu.ڦ<�0w��7v9��w��U��׫�\�y�5y_o�����N���̘X�j�"�(����B�OX��yhϴ,G�j�v�ߦkXju�·?��״��{G_���&��1�`�ss/�v��RU�So�}��:y��x/S~�����3#<Ϝ�aܣ���Ux�Ңgm�=�W����k��R���l���I(n.���x����>֣��t�>�s�]L���m.~�r��LދŻ�p�u����{o�Pb�'3�	x�`���85��M��B~��4��Ju׸g	E��)����qF���CUn²�|�55g�*2~���:��F��C{3��K;��L+F�u0��!tw5���o)��z[��҃e��HV��Tm��5�	z�t��K�҉������:�ᵹϢ���0����F<�7��¥Rݪ��Λ��ʝM�Kޭ���˗���LYO��ַ��ԋ{x���7�������œ�ئ���Wl��Yy|�}�-��ג�	pPVA���2̬�-��G��f�NM���SB��{9`�m^jꇮ�<a_*��U�C��Sf�s�Q��f�,T��]q4���.������UӣȽ;V܇6�j��}���`���;���\6Ew��M�Ѧ��:�F�#�| ��_��Q�{�9�^�
�cw�@�3����<���d��U���*�-��k�m72��|��-A
�A�Z���J!c0Y���P3��,�7�S��z����(m�������)�1�+ƪ�J�×:"R2R�KG8�MM"jB
�ŋ�con��$���J��j��o[�4+�	���e8˺]�(�5�.UJ�=�������{˾��J���DqU�Tdӷ����m���A���1��Bh4����Y�7AB�t�w�����)Pv��Ʀu����Ϲ�!ٵ��|�_GҲ���U�DuQCcV�j���꽕����	��ǰ�J��+v�j�}R�Kz�i��g,tj������V:�;�̝|��,�w)��ahLA�7���<{���u�4�ӯs_FH2�� ��W���yF��A>̘��$��� ��՚��u��w��T�=�a�16��Y�v|���Tl��b�g)Χ]G,'tgYCd���s5摥���/���9p;��A��7C���*sxF2�n�&��ޤ�+��K'R��i.��o7��,�Rқ�H�'"�1�Vɒ�գ���)���-�vj��Z.P��Yܵg��xx[��촐5] ��w�\�P��7j�E�b��Pe#rM�u�7�uq=8���v���p.��03����Qn����/���t�c̻����։Ԟ��q�m�`��;v%aγe��_T�xW�V�)e+��7g6��7�G֝�p+*�vJyQe�n:��X�N���P�# U�pRC�����ͻul.��v=U��+�����YS���6��q`
���(դ+�M�:�WG��k��v�,t�����j��"���Lf�M�7�;}��+7t���2��^����e�Di�t��cz�Vw�V�R����c�ͼ�3�Dn��ۗV� ��'8�u$f�����J2��:�9�c6jE��X�8lZ�4bܴ�o+f�)���=����Y]�eG5*��A&��o��+����r��է-XX2޳����.�{��b���@U1J�r�핻֜��9r)o�|o����$NC�B����#C��I�"�v��9��)��vr��a�P�]��&�k�uM�>�~�ޛώ�b��_~~m�UQeJ��Uu���E�d�3+U,��
�++-�̅@Z�(*,UD�u�v�*"��ȳ2�U����j[c����&�̭{H�N<�E�c�
�T��"�斶m��(q*��U��2
��j�&J�$R�a5ڢ
�F","*����<�yB���T���T�)*�S6�%j�U(���E
b�5y�0�R��'���ee`��V[hŀ�( �ZʜW���i��*,m��(��S�P�PQ`��Q���*���v�P3�/"�B*�k[%h�E��/-��YG2�����|��z�ݚXӇ)r��g9������y���[�����&t҇7-�|U0&�|��o��x�.0FL�6� �ʾ��Ӻ��+w�5�Q�U1�-�v"b8�U�_�����;NWZ�[�؊$>|d����ړ-�������q�yǛwY��r��o��� ��2w���Q�ok��3�ϕ��!N�*�k�z�c�8���W��):��E�@	Q{�'lm��Fc3�,�ڥZCX�y(����y��;��ݗ0-��ѿl$����`?'�Iq�K�.����>y�xQM�'^�i�)T#��Қ���;�{���p�����$��b]G�F����3=�$f��kH*���QY{�[�\�~�u`��ȼ�"�W�ߔ��
�N��Z��)Y�j�u���8�T�BOɪ�g�{�\gؕ�޻�nB��{��}3(8���Y�_[�~
�<�cqj7/k�W�Iv���T��ȩ��Ȏ�`̤m�������6��o�ю�}�=:5�+LJ� �hG���t+�+݊�>#2����{�y`����y��s9׋�X:<e�k[���4)�ݖ6銽%����늸8�����P\^f�Ѝ�5�1w%�}��(v=�|V��ۥ��Ud+J�j@w\�L���3���u�+y�����ws��qn~�;�y�u��S6�x�gi�?=�߱�E���0����s�OqY��p���{�����J�B�j{jly\dEֳV�����Υ���Vo��d�M�ӕ�a*�+�����
؞b�j���E�V)դ�q�����T����n�{�S���.�>!]�X��j��'���u��<9#Y��Q��j��p�݉��ʘ�@���>��	Az�e.���4��Ui����7����{���s�\2GNN3�h�э榽N�ؘ���`*���^T�:�x:*�9}�
��{��˹ǒ,S����]O-����k>�����4|����j�ar��w� g�v��y�K���!¹���G����[�e�~���Ẇ��)x�_���wc�Y��㾷,�����z"��������_���p�k�֒���!�+��t;�v�G��v��]h_orY\`��t��},�=����]i�;��ޮ��(��^DQ�v�!F�$��j��w`�n��a������gv>����x�wz����%���o�:�����	9z���t��s�}�#�����z��]��b�<ƾ�:��;q[�R۬�Cڟ�ho��l�~�f�嫛����yO�M)G8y^w��X�?R��*v�mN��U�/& k��/�2{��!�{�Q�LJ��Y�^i��Ꝭym?T����������'���﫼�-���o���
��L6���x%WtkWHl7b��4�S����ޗ��Mn\'������F�k"b����Qvۡw��*g���Ѷ�L��-��}����w=�͝��/����M\�{������GǙ�͝�����q����ƾ���骍[�������7p6�W���n�|�� � �	�R�v�x�;�mt-�nN����Y[������Q;�~�TLٟO��3!��;D>S��ʝ� ��+~�C�Q{��}\��������hP�^o��3�o(~�wߧ��S�.!�X�>�܏]��Ȁ{�A�'����,2IJ�76A�?L�b���~ʺ��U��:�&q����;W�CZ��� ��,�o,�ܚ�][����i�5�L�wQ�;~z�j~`����لS��
P��C��{5gj����Yu��9�T�(�]*���&Pc���΅W8s����*q����V$Ӥ}G߼��'rn%.�vU��o�"R����>�w+c%��,e[�Ӫ��T�}�>�Yy���ת��N����S�]'O@q� ��D��F�f����w�z�u��Q]яzםiZ�h"���<�,u_�Lz��<0���t������ɩ�G)Պϯ���c�.���wǫ�0�=��7�A��S+�w\/UQdx��ǡ�U�����J}�V�N=^;l�(�4:D��Q��xNfT<ɜ*<_�� �ʺ�"o�^�'�X��l�"�T�bĈ̙wE�z�\k���uF��훖�ߙ��&�Xw��%A귽<l<���]#��v�5ZP͝��#�S��c��S⾎~�7OH61o]����^���g�1qr<���ɪ�Z���w��G*�1�ә��9��z�s��\�?O�l�W�����#���нe��l��w�m��3jOm��2��}�#���X^j����4�m�ƨ�
ߢ���痻�@�:�d4w/�ޛ��3�wS�d���#j�f�\ب���-�}Yhp��}+v�gO{�e����P��?&f
�S2���n��(���p�F/mb��`�s�g@�t-�}&l˭��常Ыbu�5ۖ�:�I�I�YMևݣ�O�#���\� ����j�5��D��t�̮b�����F�u�xaC�;6�B.��]p`W�PT�ߢu�I���D���W���X����e��F��wZ�#��^~�cFn��=�]�ؽkNL�B�ꭲ��#��ǧ@nr���~��O��L6���ܨw�.���=*:�`�o]�R�W�Gc4�GtO�B��c ������@l�	L�}�T<u����(M�'aP�9�z��˩�t_}*����J*]��#ʒ��M��r�]���_u�`�t�Qcwޖ{�l��>���ݭs>�1p\�ٿ���vd�z�AzTA�(v�=;�Z��Τv�;�I��vV_#�v���l���xe)�x/G�:���s�;�W LwfL�
���˱�}�ћ�XNz��g�����O����_�LxR�,T.�E�v�UC���;��ss�wF�ɞ �s�.�h2�$���ʇ��WI��~&k��+�ax���{��Ʃ��{W��T�M���Cb�]��O����7KW�����ǊVq2kŁ1̽��[�s�w�Զ:����C3��}����mW�\wz�\G,���9BP��շ�����{���&���+d�qD��*�"��r=��n���c.`��2��Vs/��gc�	x5ՃG��6��AU��Y�*�'F�7�][�:ˀ�f���@!�:9�ۭ�_�޸��<���0��U��,3E�
�Z�uD�u�n��Bժ/���������rq]:�P�Vp����W��y���ޜ�]쳦-�h��gû#+i������<{'�,��G����jGz�i�&��7�i|��l{��L?`��+Zj/�����
4�[%um���<��>�y�w�!�oMB�)��s�<�����"�O�ֳ7h�2]��n�tۮ�/�5�Ʋ*��o&x.92��4=�.���;�ݡ;ݚ�ר�����;k6�3��T�Y�@SXӰ�p
��~��N'7�e�͹����vML�	g]�����H�i��,������
����E��_��A�P�w�mze�r�{:w��7�lo)�1X�OO�w��� ��,_�%�g�@=Ȏ������kם�wg	Uu��������efΆOx�o���#���H�wW��1<��g�������1�L�!��R0t�z�a�h���i�,lJ��7���Cw�;�;2޽�B]*r%Q�<�z�z��\������c�JĀOg=q11V��ND���&�x{��l���0����WbO-�Vٳ�MA����cLo-Y�t�V�qjv���[�vw��PMr�'Gp0|&��vޞ;Z�
�xr��=k���C���,�b��l�<�wV�@���O���V�v 1�1�6�i�C��3A��l ���b�T6�f���=D����-�Fm����?������m܁q�qV:l.;�۠:�2̚�/Ǵ��Q�u�Lԗ��fGt����������],�Ϥ�R��3qN�.'7g�~0����������^��~JIru����®�*b�]x��Up�(Q��,ظ��?�ܪ��7"}^���ejTc�����&<|��*�Cr�������i�p�����k�����kWb9Y3�>��ώ�D��t�g��>��Y���y��׏���؍���@����˓�����7�X/�ŷ�����ت�Eɕ$�Ύ���7�ێ���Y��=��� =Q��
f��BN���<�Ч�>#����N���`�<���ǒt���9] z�~�Ȭ�v<\���\oP�l=Jq�����(�.�3��^g�h�dΗ���D9��� x��L��a<��������.�{���F��z�}ޔ��>���ӮŐ�$���`Z&�u]�*;)��e_���]i�3읞�8<J�~4��C���|[/�:�p�,�f7�'���t��݄����s{��2�h�"�YWDt�.��j�\#�ڥq*FJ@�!��F�b��N��(�fDN�J���^��[m�R��8��>���זs�T�}�I��W�EV`,u�mX��+:��g���_> �c�A��)���j0�4��q��I��έ����
����=����2���@�>���e���l��&�3i�CS�g_*ѷ��	V]±n������b�͓>�I��]z~��b�Z�.2�7�������':9���� �]���|F�����F��8&w����W�#��I�s��f )���T>5{��y�w=Ȯ m{��i�<����<!���u��˒+����D-�����i���J�~��@y?v^��/7uK����]*��'�rn"_P��<��"�U ѿ�].;� f��I���r��ԯ�����|�#�Wb;�D��z���Nʞ��:�
�ݗR@P9f|���b��M{��
�"�<��:d+���|�äה�:���=Q
h�*!H�}!t�J���G;&�f���5F�P�����;ݮ����?�I�5A�b����@~��A��1¡]�S2��'�#��> �F=�T
B��W���
�g��Q$OD.dxA2�1Fk���X4ǿ	�����WS9�c�r�l�9�b�"}������B����}�Į����l��*���w޽�����7��{��p<c�D�Х���^W�I��i��ۖ��)ree���GL���#��v3��ѹ��q����q54��嶨�m�.��pD�E{���i�-�����Y���iĤ����*c쫅V�/y���#�~��}�y/n=Nۛ��Sh����Ǩ؝��۝7��F�Ρ8<�����^��}���5�w^��egj��V��=��d?\G+��]2�/��z�r7�r��O�l�uz�
��=�%���Ӆ�~�_�ڐ+ʷ��s>F�g�y2����1.�3�����<�#�S.P�a�u\����ӓ�u�Q�Oƅ�L�o�av�ʭu��e��t��β��xt���[f�o�h��$��Q��Mt_|�
鿢zXqU�@����y���Xh�۞\�|��ܙ�1/,���cDeK����z3������ǥ��r�����y6�f�&SF{}p�[�����m����8^դ7��D)�g��A��N����E�|%3��T=N����BLs�}�s���~�H�wuC��-<;IF�WFvY��9(_LO3g�t=���Q�^��7�k�a�+ٽ�w��]��} ������nf/�x��3�;�pe��Q�%D�Aq�>��(��z�V;̓C�w�v�E���q��l	c*!O¾^�F�H]7��Wݙ k�4=]��aY�=`#�&�yn�ֆͦ�l�R����.c�`�f�γOCF]B���s���{n���]JƖ5.��G�s�L�t�t���F�;i=ް��D1ٖp[G��b)[ږ�t,���,�2g�Z�@����7�m`X썐����O���+8�ө�2�w.�ʰy�������o��t.���?}=A�ٚ���5��(̯I���m1ඌ�����{���&����	��2�����3OGNP�dO��;L~�kْ�y��/�>�V*��ͯ�bfk^�������k��ZP\|{�΀�o�W�d�b��5�s�������.��=x~c��f5U?~~_���i>��W4�}��3�gczw��Wz+#��o���s���[?������ا�
y��z|�>�z���UJG��F����=}0<������*=W��8b��V�Ω8|���x�Ճ�4n0����+ٱ\D�u_��=��7r��Ԏ��L1O/��=���62�}����2��g&ά��|==�륤�UFx�y�иɟq��=��F�X�MSS����'X]w���t�O���t{�Bx+�Nn%�Vu\`�.+цS7�<%��}����Vsp�?����Kއ�����g[V�������E�����ЮP�.�q9���o�r�n���Ml
�?_y$
��q��^�eiϻ���:���YR��G� ���@=�wC.']��UV�]�^���LPŉ~�ˠ�w�j|i�C����,Ɣ��+�Y�VgqٽR;͝1���4����շʱ��L��;R]6���ჃF0-��ɶ0�I6�6�Xl�V�s$�z8����6�w{1�EVuAt�m�b�JdV-캔8ZLrv䵴��I�B�� 7VvA[bƮ4v�r�%�0:���iZX���[n��}��E��e���@#Gg�%�K��a1a��*�*\{�R�MzȥQ<3�^�ٽ|���`NB�r�f��yF�Nu���dR���1G+ǣ�S�����������8^VV=��T�X��x�����We�7H����ŪfuJ�u��&U��wP(X�j���ǽ�z����Gk���ߢ��{���rg\�u�&�U}�]��9�)���iU��Ȫ�ŧ[DkIr�o��bR�[%L�L�����jw�3,�C�0u�4�Wy��C��:�v��x;�t��_H���ܝ�I�i�|K����0���E����5�w{7UAB1���9���v�o$�kv�"�ɬ��39ގ0.B�0�ȳ��uɶ�Qbp�0(̛L��l��/�����Y���R�F�Ū�\_���2�m��1.�P�i�Ѱ�)�G�C�F�>�U��Y4���u��h�����[�=�u�4���v�M5&U`�òR��v-�:f�{ͥ;8_}��������U	P��&Ϯ���+W*���Y��ߔY���*��-I��f���wv:��t��MI���V�2qv�=�=}�{׶��5Q���T"�L�T���7;a鷵�4A]��	�t�8iߦƐ��}��;�U�{q�Z�/������a�r
�q��`���4�糓�5'M$���by�\FH^�LKG(�f�Ź��JK�g�n��e�6Wu��r>�WZ�lFA�:Ɗ:�l�͆Y�]t�����۰�sa!j���I��hE���e��WC�Wr�kS�#i���yK{�KVt�����tQ�<x"�Xi�kw�]�]AtH4i�q��W[�\�u��я���:�v��;
BV�g+�1�;�v�6�XA3��r��w�������T3�x��+'�	J`T�n��7L�,rT��d���*ㆣ*MT"L�-���Z����.Z�"��:��1s�������ڄ\�넵o�C��]��T��t+���ШS�ՑiT+�s��Z��˧+3q����*qR�/Mt�خ��vs$�9�E��\�`LdŬm\�$��Wq8$)���Y��ϰf+{��i�F)��n�u�����_]]�Ԋ��@h�F��{sq�es��`6�K��Ow�z�	�;St��:�\���Ǥ��Xę}
�C'{�'�V��WVM�QV� �=)↯�^nr�3��fv:ɖ�ir��[M�J�TÁj�f�n�����A�cC�񠤮ַOFu�!fG�O�_[��u�ؑ�:f9u]�p�=���*B���9��O�y�΍*t�-T/w�볧'�t��"�>����]���������(-�Z��fJ5�Ģ���X�79������g)E�9&eTX,�aU����WRfe��yH�1x��TT`�,�a�PD����aR
 ��-�#��
5�ETEH����)QVd�,U�g���TD9�9C�D���T�R��V�!E/6C�D���b4�9x��*f1��"��T�-�yx30n�'2�EEX���UC�g[vȡǌbA�EPԼT�8r��nr�fTQ`�-�N&b09L��9Z,P�-akV�Ëe��Eyj �2U��J����-��3Z�8�R,XԡL1_P }��"��br��ww.oT����*+�Ӣ�ú�l�K]�9#����jgk��Y�z�W�}t����?��z�luj��[/�G����QaA����@wm���ښ��o!�I��ORG|m�	��ʼ���g��\t�O�GTE����\n�'%��%W%�l��-�**棓=ap����~�b�^㙔���xJ���#���n�vo�{��
ݗ5;�y�8:vz��
�Ұ��ā��q�x��ω|}��L<5�x/Dm�'�e+W���H���㵠�����}rĪ���aq�F����Y�Q�����w�#�#��髭�]ʅX��2{�͠���쁟s��3qJ�.&j��z:��vz}�X���ٶ�E�e���1��E��GR�P�'�2D�-L��w /��]K2.?tO�w"�o�޳}��1u��;�|}�_R�����>���:�ަ�Tp�R@�uǦ㷪��v]��䉭�9'f�9�}�ν�,#NUF���;ޚ�t�ٸ�`L/U��OK����m`��v3
1�f�m�����w#�9�_��+�¯ہl5���5�OԬ��3�6��t�7�j����W�~ݛ�-�O�61�$���	+���UWft�SYk�Q�9ׂ�q�.��i��*B�w���%�͂��2�j��j��X�m����u�+O�﹂�z.ZG��	�*�^�y1:��\h�L9�1�-���5����:�+|6K՜���i�:���nN�VdQc��(o�������1��~c`۪��<���?dۧ-,���}C�g�3�ά��S҂�ib��Qj4���s�#9RǸ�wy[�2�������xx��~���Y8�/�l�Up������r���q�v)NU�����Q��Y�;h
f�e �߀W�@���&�'��sj	���e�zX�ɞG�#f�w���t�s�9ZJS`,�f}��S¯�u5n|�ٺ�͛��e���� v\�f�%��&�2��<�i�{�x�WTp�!���
�w�������4k�y�	L��z����b�[�K��T��{�fME��aK�l3�����$	�������z�20v�W�Y�wd76}$7��u�\N��A6���0���ݨuI�e�ͅYש��47����;����"��S�/�,_��S;����X/��9�*IY��W�^�}��||{��Q�/n�����J}`<��_T�3� 6h���^۠=�u������[���6����S�wC)P�u=Jb�=!t�J������w]$�����Ir�ר���*.�c��UR����^V�q��X�A��L����of(Rt��U�A��ulSr��n�Xd�c�&�L���W8pZ��y-�\'q�Z�Oud�fr�\fVY�s����'K����3K�O�ɯ����q����,":c~{�M�<{�e@�]ː61���������9'Bvw&��O��lG�]��΃5�c�D+���,�D?WI�����#'��<��^��k3<'��s�b�{¤Ms���:��O�*ǽU�q�����up^ˤW y��e�I�o��{������[&��6)��Ӥ�xu�Ԍ�V�r�O��q���K��'�٭~�=S�<��9��쁜��i���g#�W�_��h��Dn�±���&W��/쩗��N�׽��V�ncQ�4��^���-tȸw=�9]�do�z���%���������7���h�R�OwS�B�&}��&y϶d=��Rĺ�e«ۏ'�(ƾކk�}����wY�G�� �9��9��>��)�м�L�,.[V7�������Lr��tyïFQ�u�ծ+�`�=:F�6�ۜ��{q
�
��X�d�o&Xh�F�H����}]57UN{��T����:>Jtxtu__������!�����{9
�yp,���{ܸ���
�e3_���M�E����"�A:��E����%a�{=gk���T3 *��H3�t��w��ϲ�V�xb3Q���sJ��[�깽)<���Cm%/�f+�6�r#v��.��E��'}����f+u��mg0qt��.��Qc��#ѻ�Ak�	3�����W��V�q�-�puӤd�+�d��ꈩ��:�w��� ��!9�����5y�_����c�7����Wi���J8��ﮈo*�3���l�Jz��Y�}�-z��H��/^�'��_��ڮ����V�h뉟R���ʹ����e}&����El���e��fW������ڷTW�sA�s�w���]'�ǌ�_��nvx��57|��"�/���?g�u�^%X"��=��n��7Y�3�M~�ou��z��<��.�G�k��[>U����;�vquCx����D�S��_�f�aϗfJ��?������^�p��K����u`�u�jL���ʨ�G���7�^�U��XjD�:^����}���z}^���e>K�2,�in�ř��aV�+Fs�z���mW�\wz�_�s�wǤ3z��{mL�66z��p�4�d��}�
���v4������q���͹����8b㟅n����-��Ԏ�d���ś�"���^��Nٿ9���w�i�&��7�iyΰ{���${�߳�L̷ړ��$%>�V,�<v�]'YԻe"��t����1u�U�QD�b�#��ٌΥ��u���@6�^Z�j�����hj�Hp� 
��s��e:B�+^���J�,r4:�c�i�7�\�4���7\���J�v������71no����s��v�[��?<��L���t���Ԇ={�b���&*����Yq��݌���Nr���m�25�A\w���8]5�~~ȫ�0�f�g�㑳,>�S��8 U����K�S��c�)�+k��7���z����@SXӪ� ��~�m9���{���ͦ�e��+�*�5�V�/�����h���}t*�[/!��A�UR,��|��>�4r:)_z��h�#�u�)�xM�O2�&íU�c�e��95���eu3�LKg���f�� �⏪�Ouݪ��/����~82�Bn2y�q�Z����*q��i�vD�}֣�^�X/={ի*f�|\>f�-8`��ywCE��z�g���Ac�F��b��O3g���v������w��|x�wv�9���#	ޗ���E��N�_{>�0����x9�2�"�����vR����=��Rp����@LG_d܁jC,���ڐ:b�Y�Z_�i�r9����OV�t�=5�Ǿt&6����t����hw@�u��ҡ�����}����Ǡg֐��_��س�&�W@�����K#�6��ɫ�u��Ѱ�je�\Ւ�.�hM#�:a+Ā���r����Ί~T������L�5�efغ�M=^+�e�β���i����/u_}���EX7v+!ډ�B��(u�cGv���]X_1��b��ݔ�>Wƌ��<�����
���2zb�D�8�W\r���)�d\~��(����M�����������W��؍s��}�`l�G�Hu��\zo�kƯ��[��V�t��~^O�[5�n�Y<���\:ۇ����3ޚ��7Le�7�x[NO;v���vgT�۟W��)_��K:Xo�w���A���� k�0מJ��� {�k���@n�W��M=���S���'>3ϫt�sc�s�ς��Y_�]�ط�]�=������z��?kQ)� t:�]����c9*{Uf��3q�ݡ��PQ���tׇ�j� ��dWD���*�z]�����=9Yj���9̽��29��ؤy9Tq�.iTg�}�+>�)�u�Ý#���f}�������W�������������&yٳa��b�}�����x��j��@[R�k~�R+�whb�m�֏A�P�w�T^���.W��ʿ�����R�y�iܪ~۷:�bU��?���7;�Y���Z�h�
cz<ds��Ҡv����(F\�f�'�W�V�b����&"';����/06���&�t�t���:�.�UU<
�5f���ez��bh�Zfi�ǫB�ݯ�g�rEVAZ~�od��rՖ"cپn�<	ˁ�dHX���G]&fх.kBպ6��2m�&�^�M�e�s����(ZŁ-uu����,���6��I?p��0,>|����n�ʈ>�������f )�[)�{�c�����k�HsߵހJ�����zOq�;M��vY�ʧD_:X�>�܏]���Ύ��n/w��Op�z	�:�c�}T��K����!ź��.U ѿ���㳝��y�Bo۞��w�*�.��43Ox�Ac*��;=*b����zx8�/��I�W�x������]�&I��������k�|:�xg��,R���];��w�_����v�ܨ
g�lN��̙��rhS�}�ۤך���^M���K�=����w\/UQd��յ怋��i��Ղ������ƣ��${I�:��W����\���`���]��{�����v�k[���S}���8��'�����}��{���ۢ��d̲�3~_<z�7�}�Z�X���n�ad�Іwݪ��o������WX7z���F���W�]��'��[�M�~�y=�d���9���2;���K]2-����fT{w�r��O�l�ލ����~�RN���Ə>��{3n��՝����ֽ��:з�au+�r��R[@J9��V�Y�;�.ԚqS��,-�r��Kx��^vVr|5Wc��DR�I.��ז�n�kGDZ��`Av9��Z崹aK���G�}��Z�n�a����b��,O0uU�ޮ�B�g�p�E�ِ��k��^j؜�Lҧ����Vvg *��+_��
��f�W4��DI�\�]�+��h^L�n2e��V7��gm4ug��]�Ua�]�&GxoB��2a��o�r�{��2Ggz���L��2�G>۞f��G��K4�K�Ws��=�\�+ᠮ�+.Y^�Bsg� ��2.�'Z�6�e_cE��s�����7�*w:.}=	�B��I�����D�Tv[�,����d��:Ϸ��{̝u	�z����E%W}Cz�<'ӿ_�P�'����Ǵ�n1:{<n�[�rP�����X܈4`TK��u�c���v��_��ۥ���Tn֎'Ҧ<\�ٿ����3�໣���|�E����Z�˻�3ޢOD�6X��z�
�����9ỂX���<O
^�Dq�bm\��W��^M��ii���]����,�p����.[�Ma1֧�p<=Ki�
T%�՝��*z�r�_���|V�������]R'�S��\I��>�^������׋�3ߗx����W52�fg�'8���/�fx,~������%�Z��ݻ@<�7Uߦ8���MzyC;�-f3S�N.���{���W[�Y=ǺS<+y�.��#�{o����u+���çI�z�bK��&�\��דF��UȻg�t�n?�����uR�����;ʱ7�QQ��	zr'g��Nz�����}ޝ���!�=��A�^꺞e�35����q�d���������=;87�({>��jp�{�{ݬl���^����^7�y��M���0��=}0���z�d�w��x�������ڋ��8}�TE��W��G�;ǵ��Gb�`	N��u�Y7���}Yu��j���~�W��Y��xRӎ��%e;��P���a>��w�!�_��c�7�L�'9��1�����Ϻ�q�=��Avȗ*"\�egU�O��xe3q�<�:r��P>31��Aՠ�<����Z+��}n��p��g/T�����q����� ������M5$�Ώvn從���29��F��=t��|w��t���W��>+*Y܈��<��xut���o���ڇ��O!]��߀��oKq�̫��`h�����da��뇃r��o�5�I�yݒ7mL�Q��A^���wC/��~80ۤ&�'�Y�����:-t�R�H��Q�}��ޫ
�:�[];޴�����Vhn�a_�9}R�e&���"�B{��=t��}�.�(RS�{�S"�g�|w��:�$��#��<Pw�nuq��6�Z�ɺ9�	�̬͜`�}�1��a��a�(�HFd�5�C���]�묑	9�
N��.���q�����d�hT/-��LN�����x\D�z�d����,uDl�.%mt�1�r��8�*s�ݞ�׈�@�S�jڂJ���r��7�B���Ǫ/�p���l	��i�;�ʧ�~��7���#�)�nJl����*-�\�q*�*�6;�����"0,����?VM���MVݔ�g�Fa�GNQ��x��]@u�q�����S��E��Rg�/|jT�p�}Y��і�UG�.�~�Q�c�f�ǇTB�P�L���}x�5UØ���̩fA�����5�p���ߵ`2�&f�Um��ӘV�|��ޝj#����	IuG���k��m]v�^�Ƨ���<�ww��`\��~v�A��o5����d��� V�Wu�Fw=5�rG�W��(�/(L	�6�O�U�y^���A�&�Y�Gz���%Q�9ݳ�T>>�5J�w��<i�;s|GZ�Fs]4{�zn��A�:s{�����G��~�ȫɟt�?di�\����yGf_��)�=s�%9Lͻ�g�h���j;�D6���V�߀q��&n��L� t�q;B��"�4l�R�Y��n�vB[�G��S�L$�*ը�������m��`a����kRM«\�ϖR;��k9���%Yy���r��,�:j�֖���39���T�Ct�52��qm�Yt(ɔQ����=��r��{��X��EY#Kzc�6������Jf�H˩f��i����WثT#E	���֧��Yw�G� ��Ue��Ĝ���v]19�h쵲�������p�	#u]��Da�;l���L3�X9���u�1SÖ3z�u['X��:@if�qĲ�j�*i	Fg �Z���r]���q�������V�hm>﵈�L��λ��vQ�[��u%Z�;�B>{:�λ�+�d���2���1S�Li��k�]и*Z��7�j֪�}1W�����8�8t�)���1��Q��-U�3;Yn�����W>�M7L��u+k��L4�DS������;�b�{ݠh`u�{��M�G��r��&�:�v�gr�,��Ԗ��YQv��ミ ���a��A�1[�=��a���P�׬���t�Z�me1��cs,I�Z�E&��m���r�%��̒�I_=.a�Bu��Z�Jz.ܶ5R��׵a�t0$YTx�˩Q�5f��|%t���A��Գ��D��PtO�:���� �L5�q>�-�x{�LݴlI�}��+M��.��ڕ��R�����`������j��l�x�U�kmu�.�Q�:噙��T��`t�J�u��1��@#���Gv�XA�U�ݘ{i��!O�&�a|�ԙ�y��À��@|C�zϮn� !��RY��b#��v�i�r���2�۲Upxhk���O���޼��#L�@�yK�;����h�ܿ��K���tU�ו.�>q$6_7Vv2��jW��Q���s-�v>�*��;��67�'%["ӠN5�E�}p��n��ը��n�-�%71<'o4<��E����.�V��N�*�-��0^��Q{f`�ɵx�v�6��H�G��
PQ�/j�vJ]ak��`��Ƚ�JPe�E���3o�6T�ש^��nnB巴6aec�D��ү-�·i�g����HWr��X�sΰ�R+	�쭃����U������6kRu�`:�.��:t.��\P&�qB=�����J��'Y��!�&Dy����l3�xpU�cp�I���u*9)iBxv��Ƴ� BK��*����=̎�oz�n;}]|�b��n�]�< Π�t��9��ۏ+V�{���"Pa��r
Z%A�a��a���OM�8�gj^;�p��*�bG0�r�8�*Ҝq��43x�`����dt9��ܜ�<i� &A�ҡ��s��K�o.��n��<���k�QQ]%-f���O�q�tU�'�͹3�P̭���g̉��o���-�בګe�7x��UDQ�P4VUE�=^nm.L�խ�
ؼƣ�0�е�33xܜr7�r�V���RdU6keJ�m��X+��mR��mjlU�ݩ��(�
��ѼL<���%(]�uD��5\ʬi^7(�U�AUJ�X�ҵ�Ţ�b���Ȣd�.i�SX�5�)ys��Z���TeTV�eAF�[Q�Q������Z�+�X��+���lKb�Nk�����l2a�VҖ��AJƙ���V���g8g9x����*q6�Z��hT���
��3Čh�4ek"�*1-�k��l�Kl*[J��-��[�k���5ͤZ(�b��m���0��+ڱ�emeUX�TɳPFj�v�UTDunfVf�a-j��)Q�E8��@a
@G�"R�v�G�o����Úr^��io@��"����m�aq��@�(�+�1s��N��_V;�K�5�TG.),�䢝|-.#s�����y9Zd7�T<�'*�C�C��>�q����۶��<*7�뛋��{�)������;)��6�K�����+��l����;� �S ��ꕾ��P+әF�p����d7 ?*��/.W��ʸɱ��&�g���磝�D�o�l����6�8���+d?-�=*t�N�`^\�f�x5y[���X�1��������9�87��e�]�¯�܋��t�<�������Q��{.�&ڟVP�	L�ʖf^�m���A��]�O�q���v��8;�� W��Q���cgn#.��]��o*�l(�H�����9��׵q>�F�|\��@]�D8�U�Eʠ9��;�+�g:w����K�"g�9��T^u�M��ѹ�,b�0�#g�L\AΠ�rO@��\����x{Į��)���@�藦���м����pzJ�����,W�GTTC���ۍ���=�X��V�~��t� TG+&�Ts��w*��=9�ǽ]��΃5�c����7��B������=ݯ2�RY�C���n:q�f4��]H<��k��`�([�2�W�k����U�v�4��5��"�`����Yf�vw�7���m���E ��~eokE5*v���@��}��ɭ��*� �.����q��֗�����������uC�Q����dO��}qշ��z��{�^7����noP�G�%��NR�o��J�w��"�z�Oۜ��ެ�L�Ι#p�u�#;շ��N]z�[}��v�t�K�O�7�@�'@O˦���놳��+¯�w�t�s�:2:����>��������Ż��+��\D�5��#&}��#�o�2;����5�#"(���w�p����R%�E�<�s����^98����?S�B�ɟ3q�<��C���	�bw�t�ى�ix�A���=��3}]��]�2�˜E�UX���h^L�o&X]�V7Z�\��\`�������V��G��LqR�+�}�%ʉr�{�
�2vw��̔���W���;����+*o�s�|��t��u__���e�ܨ=,���yp.|�,&+�Y�A�lv鮩���Ʈ��o�t�j2e��>��>���˓�d���ΡD�͗f��9X���IT�+���d
g��d���z�\�����i(�c���FvY��C�����ٳ%}��!
��BH/[�u?�h�8oa;x&����V'����1M��S���x��R��5^�y�.��|����-Y]ٳ)�(�<�3�rF�P��n(Gԫ/����$�# �\��*P)VvBӝ���e͗�A0L`�G�I;�����J.fg�	��dݽ=��V������&K�s��c��.x�l̝�M=�~�W��O�A��I���>��:9z��~��x��D	c*�<*��fj��ý����vΩ�mI���o2 ��|nR9H31狪�Lv\�O����_�Lx{�l�~�����vyrP|�U���%&�kT�;��Oz����T����'o�hv�lך���9,:Y���'젚��7�^��&yTgWt�<_}�\;ʱ|�ԉ������Umpح#�v���:���Q�]�������C��x�'k�:��@�WWq��q���2w�;�?����ɼPk����c�Ӛ{	Ì���,	T�l�t����ޞ�ݜ�� �l�ID�ob��I�m��Mv�
�=$�űvFWz�Oa�;� y����`	N넬k�@�&������Oö��6���B�#��n9�=%�����ˡy3�9��$1���� �J���99�7rtOE:~=���C7�i��)�˜�������*�0�gy�|
��tdP0�M2�
{�W���L�gN�;��@Ts��n��pm�3H��[�.j�;�������Z�h2�eM�m`�/���wi�=��֖��2��%��ع�J�`�MC-Ӭs ��N���nf.|1�W)���\S���k>c�l�s�um��u9�w콃��q�V*Jeo��lp���~�ʋ*㒰-�ٸW(
C��<,Lm<mB����S�:Sg�}Fq���|V����n����,�}�@;5�_�F�K����1�5��+�wC/���i'c%�����Un���OO�a}�����s&�Mv�[3Uޣ��Ĵn!λ���]N�G �(N�<ʸͭ�g��\t����C���YN�}�#qz���#���z�GCT����g�
��N۳�~�ʵT{�:�_��d���jx��U�M[������m�x�v�<�;�Qc�)����t9͟I�}Pc=x����3p�Ut]������ ���g���W���l�p_ϲ�5��*�*�t��;��z߶.�ݲrk���<d��/ǉXiP�u�F�.���C�9�t���C�����R��ԣ�zwcH�}8/ߌ2�#�00k�ڨT:�Tzb���j��d3�������H��u�9��T?_��#��Gr*��i�V�������A�K"6�ㅩ�W����_�>�Ł��*U��l���=�_�Yfa˶�롦=���g�T�i�m$QW�����ԵZ��
&��w����cڱد_��[O��-���vs�L<��J=�؃C&Q�"�][�(>��4e�j�ƾ��ڲ��.�P�j�L�ʔ���9V�y��})e��]��f���Ѹ����n�4�=i���������z|.��<ݦ���5�&�o۲��j�����=7|�����+��� ���� k�0ו7�ϙ;A~>�jnw��.��|���3s]�'�ٶe9���X6����]�kN���a�/=�n�D�w��]�k3ωɥnv�x������@O�Γ3�m�g�pk��b�Nk�����M�˿c��^�\�'|��������7장�4�n�z�T#�ʣ�%�sJ�<��<T����&��E{a�m��y�W������O�^N"���a�������;�$y�L����tWv���s�����a�='b��WxE�?/�˕�o�ʼ��jP��6���\��|����=Q��#�V]C^2������E�N�X�\�f�x5�>��9�9W~�L�����m˭�@��WvvP���(�t[��@of�h+�w��^Nui�����~F�f�k���ݨg�����;7`pw�vY*�q·. �Jgf�/)MY��7�B|�%[���O;����csHv�@j_��e:έ�R�gL��i�Ϗ�Y�] �
A�
a�v�^��۹���϶�eMݦrf�*���9�/��EI���gf�=�Ӈ.z�'�3(嶫c[���w�b�9]KQU��%��Df��yn�D�Y+/����~xݐ:ʍ���}���9/�qʈ����s'�/22���ti��鞻�$ھ�&��9�;��5�0�g�L\��n%O@�#��wG��[/�77&�ܢ@蝉h�3����=����5���u\mp�)�X�R:��A���g��<ڎWi������Vb� ~�2�*b�;_�[��{�S�,c�_���Op���w&m�Q*U[��d�+�JO\wUq�9V/{¤O9(�O�;
�{�=��&��b���uѳ�I���~�1������:��T�&��-�'��ە�7�w���(�|�í�n����g��aW��8y>����tgGz���x9�.��%t�m�g9exW�*t�s��s{�'�����S�'��Q���ڢ/��W��2g�1q��7�x�����L�C=�7�s���,bKɵƶ˝�]sU�g�ω�9׷��Uxy�]��&|��L�/#fCݞ<��'�{c��z��ݹ4��\�<��ǳ{�(��{L�K�e�}�x�xhz2e3y2���j�f�;rd�K�b���$��H7o�]>���s0*J�`�}.jS%2j1�Zq	G=TJMZ�R^J;}8��9aSp`t�U��6�YLn��aɚ�q�^rpw�$�=Nt���WXa�]]��[6y�����M�D+�LB��� 3�M���vke��%;Y��>���߹�p����q�Hp�+K�܎�����*�����2S:s <��6�}����f�\�%R����W�Q�<7r=��E�__
*K-}2�� �:�hg�x4e_�;�^~䶮���W[�n2a�7�nT;]I��΃���ݱ��u�@l���Gw�.�3��T�H���uC�<��0e	�����
�'����_[��_��d{�m���Ht��uf�7�3tg��bR#����]���9Xq�V�h뉟R��.x���{O��������j��ۓJ�*'���	C�#�`xU���g�}����]'�����v�v�R}��=]	Szx_wf@��~2��^c�)E7[�Ͽ9���v�X}��;����1���J���\��G΄��4jH��*�w/(Ϩ��:Uę��rW�p�Lk��qY}�h��c�O}�&j=Q�һ������muW
�j�W,5"y���n��2oq>�k1s̫ۺ�b�{�������ɓ^,	�뎸Fq�/�=��j�*�׃b!N�w
?�p���k2��ofŇ�;[�Z�OՖ�-��ycw�nc9�8�&��w���k���YW�W��J��m'�ů5uͫݙ�7f:w��w�(ˮ�n���Ԛ�/���0�
(6^!��u(+��K��� �YވCtZ�������{CU�w՝[ݛm�S�zē�Y*ef��W�1j9UBk�Kg�Н���>�i�O�x�G��tޖ����:�`{V�}'�ռ��+Z~����u%���b�s�����^$Z��L�S��2?I�� �Z�i�D�Z��m�5
{�S�x��X={��L_����T�q��x�;�Nqߣ:@O*${���'u��]�퀲�u3���S'��|���5v�S�'+���+G�C���{���×[3ه�6e��l��5Յ�2�N�����=ɔw�h
v]0�m� ^�q6N�>��9�e���\��鿾�<_�na��k�{e�h�z{M���q2��}[^WlnI��}�Ⱦ�Ⲁ�R,�W�&��8[)d�z�t�����y���Ur@�t��:MMdY���_G���	��U�<��	X�pto�m	�u�%ZYhٗ����%��%^��yÁ̹��H����ǌñBy`����{�x3�r���X��ěw�f�����x.�y*|����;m� �;2����_:���H]�����^?d��xG�~�l;�sv�Q�#X��|U-̽)�Gg1w�����������Hڮ��|���@x���V'ZUe ���һ�w_\�Wr�xWb{T.X��jf�{�Z݇+6��e.����57�#�����Qt�FS ��.����Vz|O�fhJ7f����1�i!<���烛���
�,
��원.�UG�z�.+���Ō9�K_��y頯�}�fMx�ӄ�4�L=�2qt���Һ���u�g#��ü�Q�}Zf�dT\V�K[�ٛ����~aA��<<f| �Jd��>�<j!���ቌ�m�R&X�Qf����w>��r}�����M�N�>�F�\pD9��s9{�/�xz�'��k�B��rS22���tk܀٠���톿4�=j��f��xl���fW�b�R�]�����a��@��t{:lzM>U����;Rp���b�ͯ%�A���z/(~���T�Lu[!�����ʀ�]7�m:�/>�YsA���f��r��ۮ��U������i��=�o���Ίh��~=q������z���37���r#���}ޟ#}�Q׆hjߣb�3����<��:BUV���dU�L��/&y9��,�������7%q��U��(��|���*��]�H�������/�t��o�D�X�KG�͆�#i������{���0HC����꒖��]��
�V��(.텎����S�B��G���R�\�e�b�ԉ5�,n�BU�v7�C�CB�2C�coY�c�E��v9�Nvk�+h�vl���N�,헷1�Ja4"�w@�R�]�6p�`�0�I;]�˖Vy���L5ʞ1���nt܅w�U�?2��;-�q�`�w�R��)N�M
*���GOWi�t����8{�U�g���q�ٽ#%-�@%��+)g4����O�؟rw���;�ӝ��
�u .f�`!)��#^�}�4=� �[�+�3�J�7���o�>��Tw�ڇr��M��:
�68=��!�ˢ3�T8��~g�u�����}o������w��<�a�%���U"������"���&0��.yo��V*�OzH.@��t��}�@z��ߤи�=�p1z�C��S��P������]#�t��V�5��ޮ�B���I �/O�j�~�G]����������L���F�]��>���o�4gB��DJ��\\욑\�r�ʫ��Na��=�΃:+yT�7��ϻ۵J�y�M�����d�7�Ox��뱴q�ؖ�(�f���V�w�O��[�Q�1x{��[�
���̤�N,=Tz!����H*�p��S9�\-�'�m�Q�ɱ�bg�U�f#�]n_��v�7�s��ذ�����n��3+�ٳ��㱕�6E3�X3)�x�����S���̫PGN�h����*Z'7:u�n��X:h]:�n�z*Ia���u f��[�l	g���#6�^+2cW���\5Ƕ,�h�7����T�F��i�=�O�:B���R���]�D����"�s	�B�
�4,��V�A���'	mV�5� U=�U4pQ�eݒ/�Rޘ������і��� ��S9d��`�J�0�r�2
���`�΅����r�F�ŷB�p8����;�슶�1�WSq7�w:����:ɏ�Q��B�����6].
���!!��.S����dw���p2��r�j��/i��
��wF�C����0!C*s7',k��\��u3�iAװ�U�Q�mR�W"k]��u[���Z�!ӕw���U;ש�2�w�o�:�m)y
�\ �,\�g#�LP�6�b�q�@$�Fa����v�9fΥ�u�9W�v��/���/j����d��y��vs�W� ;#,���%��HΘލ����NRX�<�;����.j�Y]2&� ܩ%��R�fs�~�0�m�ԨQ�.��� u8}���%����x𑎻5���y)��Q����_fo=�n*����9�]J��tU�d}3.���`J�n�^fڭ�<1rK�"�c�bW2�E���+wF��cA�cڸ�mE[���uIA9��ȸdη(��Rj���WQ��'c�P%f�V7�
QS=&��Cu]�܂���Fp����e@mR)������f���P�K�aW��J0�/���.޼�����?T��w�Ux�	��f�M*�U��VQ���m*��U���e!+o(u��uԴ	w���j���W�Y�������G�fs�@�	n�i`�����F�R7�����X�b`�9j��n�W]��x��KV�8��3^�Uܶ,��(Wb���K"ҋ8q���eݷ���ta�t�/r�5�\plj��sF�t��Gea@a�O<ܒ!ol5yj�.I:1fe +�kw5u;�Ӝ:qԺ����Ȧ�4�·P\]���ڷ���#�rB&�X����ue���Y��3{:,j��:���WYu����x-�un̽]���ީA
�V ��e��+�'��~L���Ϛ޲�+ԥ�4p>���v��@M��>Q�SPK�V�.R
���il{V�X�Q�DM�[�������]!�e�T����ZomR���2�CM�Hۨ:P�	[���ӆ��K�jHQ�pn��ї]>cyfk�\��Z�b�r�_/���앓nk=\�^Gbs�cnt�\�JMx��5��=8G��Al��Պ��+��y���FZھ3�\�t�f�9s��@` �$	Q��Tj���l�E��ډjUZ�����\��֖��ʱ���kF�J��TEQF�X�[Z�6U�u-j �T�ҕY0�Ԋ�Q��-Q�L����N96�U�UDn�(1��yJ(*(�&�������DX��R�՚9(��UT`���拝�����2r�1���5�m+m5S6���`�m-�3j���Ym�l���PQ�F+i���1�j��X�D���T�c-xܑ�(�cj���Tq6�ʶT��h�VdmX��V1T��f��Վ�� ��T����DeV֪Q*-�L��QEE+UT2� �EF�*�"�+Vڠ��m�$�ڲ݃����إ��*":���Jʋ˱*�eJ[.�f���(��Ae��[U-("���+TT��Fڅ�,E��E�   �
����44f�=�u#�l����H��Ce*l7Rs���n��A7dw�q^ƞF�T��7;�]��Bγ���Zط
����E~�M��?ޟW��z�ޗԝ+�Y�d7\��c���nR9�p/D����7�p�d��)ќު���U�ɟtǙ������d:=�fV{�oVu
��-ũ��ټ񚾋�eK=ޟ�Ϻ�^g]���xh_�3�o&y�l�{���F�l�p=���T+�	���s��w#�a_n��9q�7v��yOƅ�d�f�e��+W�����k��ѧ�Y�M��ݤ���>7WHp°����NK,�Uq�;;(%]k��߮���k�g��a��Of�2��Xk]$u��ԇ�꾾2����\� ���=M�e`���z�FV��������Ɇ��ٹP�u$|�g:��v�잢��;�J�oz��~�+#���oN~��ld���.��<�]�o�ݨw>��#�J7�G�.'<�q��n�g�#z�N�Sb�9���`mE�_��n����,un֎��R�Ma�1�ns��PUn!F`�\�5(x� ��&���Z7��(v�����7��-��Uo��.�� ~����j��i����V��EX�D$fu���'nCk[��gk��1Nc�Kv��Ψ5��v��"]i���/�p�-CJ��+�_]�z�vN�wz)-�ޞ��@NN�,��|77��V^s�C�UI���淔v�-�0�7{ÇLI��-��6��EXN3q�}5lgW>�����_�7��sh.��$�
��Y W����T9M���.݉�&:��My���r���;i	Ӟ�vj��^ ���h�>�2;���G;�2�qD�蚘<�c���1߼�hۅ��]&�_���GqUR�|�O���Q���4+�ZjD�)���<\�С�Dz�<Fbη�.���׎�3:��z� d
�Q�}�^Vw�5��I�y�|�L�!��L��Ϻ����_�{_,y�������!���O�\�(?�~_���S�Y�8�P����+?MY�r�zF�k�w�_����<�?\o!��~?M����Ļ���J{�=� �'� ҺB|W��U��#{�(����=9S��"��x��ˡq�>��p�z!��C�Լ<�X�'��{���j���]��������Nn%�R��i]�m<����rO��i����oX��ɟ�q�ٖ�Տq/g1N�)V��_l�,NϵLT<:��j=(�D�2]��� a��~�!���na�t��x�+NGt������p�F)�~q��Y�6Mw�$M��~
Kû]Y� �ٔ��}�j�p2ۣ�9̥�����o���
�^�n�]K��5���v�WY��ȳ^���QSe��u*<�]�j���8PV�� ��]��5[*�]���J�_uj̔�0��20�	.Zpuf�ꀧ[���@K�0pJ���=�DU�ɮ�7�΀Vl�@=ϕ���~�my-�y��ݟC��?Wx�#[��E�s3;|��Փ�Bv�@�rX������:�\�?��;<�͝bϐ�
b�;ʵ-Ժ�N^(<(�������$>������|`������q=޼�G0d8Tj<���y~C����#����=���C.��w	�;��@�r;����S������p�炥���\�����J=�+���c�ֱ<)zi.x9����
����]R�US����z�1������2M;	���<�=�2j0��i�^ ���4k˨	�.�:��e�\谞����ɺx��]=8%��y�����]U��
N�Ŏ�B�ҙ=1P�$��GS���E�����ԛ��B���R̋���?�ٝ��ʬz���;����,c�]�����J�o~h�~��j�/�tGw�ON>�-U�{��hX�?���������~��z Z�Uz�ڼ�隚�B�D
�e /��z�k��ϽX/��ot�:��ۇ[)Y��]~�4�l�����J6D]���7���K`��y.�$��w4��>��$!�#��>���
/��ڼl��2���d�378�'ʜ�EHm`8��Ę�m�9w#�@����U�JXM�-�=״���z������']��S�g>]�1����4��˟T+&������rmn�P���슿�g�>el�\oP��e���w����ɔq���WT�꼣4�6ǧ�жL�d,�s^z� x��dϜ���<��i����v)NU�K�b��D�;=	��������E�oYE4�
d���j���E��,\d�G�f�{,Pޠ�/��_4�i9�#}��3���~��U�g�eK1���Cr�^���.W��l�kp��ܽ�4�y��b�WW2����aw<d77�OS���U"�}:Հ��k����۵����ߣ%i���=
t>��,(���p����<*"���}=5x�nn���k�]��Q�lW�g%�=����� ���߽Q�k�ݨg���A��;q�#�g��T<�tF�Mzn�El�����p)�������L��ߏ~.Ұv6PCi?�k�y�j ��ɹ}@'�S�i����t�-�.6ɞ tG:d��G�]���m��u�hz1�i����
���LS
���Z�Jbk�ݧ�����m����%�;*j�-w�?65_n���3#۽G<x��l��g'�	��X�v	`wj���R�-iF�h���U1P.V;^H���U,�P
S.�.�h[@gX��:���1;��wnkcX�h/�$U�a��2���,�ДkWW��GRfD�l9����=弅/�jD��a� �OIҢyft<�Y�~a\����T���bf�n;6�==#�\����ۋ�!tԩ�=�e@�ɩ�G)܊���dW�a�]�������Ң���شb�1�3ʰp���!)��TC�t����,���G/�5�>�ڎ��G�u?L�<i�{s/}�\+�}���o�q��`B���ȩ��.!*w���s�?W�=Vj����t'��V=~�yV�*Y
�umH�~������>����z��%t�p�p�s�W�G+��n^@W����M�Qv:#w�F��T'�G\"�{�奟�g��-�J�V�PU���26��[�ٳ{��U�O.�\-RQP�Q-���uQ�~����L�����Z���ӓ�e�<ܺ5��g�ޫ����:'��7ӟ:�q��r�.ؙeK�e�G]���&S/�>�]�Syӽ��u
�4���X.;e�������v�Q��}q��%�g@mME�WJ�^��χ/y-`�߮�x��|n2g�G6烿��F��#��cæ��ⲥ��Cs�b#;�0�d��}9���o:�a�Pf6�L7���N�m��l����͂��F:iy�L����d2���3u%�쳖k<�u;�}�PWQoS7�淍·��½}��Ɓ����'���%�]�a���7¥\�S��V�us�r�*����d��}3d�jsna��H�A��<�@������pQ�!8�q�ݫF�sU]�_3tC� .>��u߆dl�8{���7j�>��p�i(��<'l�)6��_U�����+��#reQC\��7�����_u�`�àX������쉴��ڤ6ssG5�o��͝;=g�w���vU�-Al�L�9L�c�onh�c��\!-�^��j�{��v�ޚ�=Ч����#�];*x}ِ	���
�R�r��5Q��u_��Xz�"rnB9�=�z�x���'��z�i
�BX\L��} .UC����*�H����wȍ���(�u���WwL��G����Y��rn�Mx�>�|UT������x����d�a�R�r���Y��;�Ϥ�="z���)j�K2`��,x��'C��޸�����\�t�F�����ٓ���9��[��+IoV�dO��{#��^7���t�i`L*w�ʝA�蘶��*��#��0��YQ���y��߷�x�k=0~��y~1޷�9�¾���!g�-���UJ؛կ��^e�3��*�KyW�A��"7ՙ8<@���K�J����(�e������Z�r����n�����kN��1�M�ށ4�[��&ou�:���Ku4���鯋���HQ۵�����F���u�Ci �F���[w��W�fwR {���s�.�`{��(�������t�画<i���O���O�D�䮭��)Y{gQ��B�495LMӮ���l!��4�퉖T�������I}�,���=�~ȫ��;��g�㑳,;��V���ث���YY�#��,����W�M�I���W����;�������NneCnU��y��S'᳾�����s6)r�gy
��,���@u�<����a�X�ɴxM�U���#��ר����{��kު�]^)�����d��X�LKfϕ �#��e��?m�q�̥�%��QV�{״%��@����_}.��28�R�>��q#�zj���+.۬�����,9��Ŵ������}�vW��sg}��:�wK��l����w��S�sp.9�s6}$.٧c&�ʪ,B����4�eeÉ�]������1�k7�p�F�:���� �2���X�J_s�=Q�s�{+\���m�����M��~C�~��7�L=�2qt����>H	�#O�(Ȩ���NU����#2�8.�0O1&�)l���{L�4��jƗ{���<k+,cl�De���Y�E����`��+ln2�g��}Qc�S���"�ir�V(�`n΢
n�.��N黏dUj��KQ:��2g�=�L�����3U��g�G�ŚS���Ϋ�u�[͞�%�{���'nk�پQ�j:l�uZ*�a���d~�?����4�so�������g���ڲb<Ѝ͞�mW��Ū����!T
��g��kƮ9��E�,&���_���_��Pz�����ޫ5�N��w��r�~����ޚDy?�Ki��ٱ�.;�X�;���:���NB*ymM�Geg���4�d�p���;7�=�< �}��L�n{žu��o��Z-?T��vmw�b	����ݍw�A�A�OEr~ɷNZY�L>��3�K����`.�>fd��{���ׄs��>R���w٭l��P��MY��_]�)��"�&|�0�NW�d7{�aNU��i�g1�G�yG�':�{Y���Y��~g?_���\ܰ�U`�����E�%����7�jw�E>���װ��B�D,ֱ�������G\q~����5-X	����h��W���Ҝ���V7���;��}��G���/\�;�3{��:�D���Ξ��>Wt0o�Lˇ�=E��K�Jy��J�#�:{k������(����l'/��{%�ĉLa;�+���|�ݞ��*����K;h��b�_��i5�̮4��U��hw�i؊�lە�T�a�g%K�֫b�Y�M�ֽ;q��&��u�^{��Aå!g�\�Ϟ�`����x�
�x����V�`��;�':9�{��y���ǌ�Xn�r�*�'���QQ��uߪx�*��-e��m��ʇƢ���}\����:�����K�2�z��ׁܼ�b����Dw�PE��J����X/�|��>�^�v�uϪ�����S�\�N��e`kWDr�wRE�����\V�H5nԚ�9�;�es�h,��ߓVX�=�\��rJ�d��������\��tG;��ʉ�nf�C����Ox��;�>UIt�y�����=~���z1��(WHU����M���\�����\+���a�9��oý�Լ�}�X:h���k��
�Z�,�~����T=�!�U���R&���سU0�_��goԎ�]���==�\v}�Ux�x�vvXЫ������1\TuϤ�r��+4��(�~���m�X���5p��<hz�:��N�� ς�z��sl���<�ϻ�=�"\\��u�b3[�s�gv�u��/\��,���[���]y�P�T~�~��~ɾ��?�
��iQ��\��	�/��
�`�`s
:�s"�VP��Ι�lĉź]�Y9�N�B���y�y�e�k/6
�9rK
��4�u�(Yw��5�]Sn!v�ܵ�q�0��{i]���Dю��_S�y��X;1�]L�\aP�N0���v�t�Hm�y�ػ;S�v���t̿���/�o�U~Z�<`{�~׮�*�ċ{�Cl�K1��O"�[�0R��7�vր�F���B�BR�Ӻ�Ӑ���wz�Y�L���s�w�S�~4(���������_�ٞ�=�,odFՆ�ƹ�������1�5Hp�+����*���,�3U�;D��0//5���Z��0:;���d�%���̮���K�����]W��"�J=Y���óu4��wG|-�AS�;g:�yp,�镓��ܨw��7�����{�|<�����=����i�3����RU�� s7�	�w�da�X-@6�d�)�ݨw;�Ȍ�yC�5��M����؜]��O��"����GFG��6|%��z�U�_��n���1η�q�Z�D�߱Ƽ'9
�Nb����m�@w�pi��Q�D�l�;s�]��W��4g���6{+���R���
�.���X�^�'�ǌ�[=Bzn#\��\P�ƠT��F��B~]+��|�kY~�ӽ!e���y]&�w�U��ǅ|�K�Ѩ} .���q�/(
�w�"}��Y8����X.�n�t��۶�n�'%}�T�֋i"j�����31e�[-�׸y�Ϋ�2־wx[�u*�U�ݿX�y�6��;e>���խ	���a�@W���]�@��6e�#����p����+pl�?��]3�l���du�ȵ�t���١��R�0%&���T���k]��4�a�Y�&
7���5��w.	�	U���X��(����D�i3'}��5��K��x�L�
�o�XaM�b�hZe�[{���j�q��y��R��-���9]� �����<�?���Z����ZYj�I����M#|��DH_9|�uXϥ�7tl�`t�+�r^^�G����>��1v�
SʙM�)$�@ӑ���Z�J�!ή�i|^O�\\=x�࣪�3ç}�.��� m�#rA(��M[f�}�i���,�N�Ah�X�+
L��ӥ"��f�X�pw��luobht�DQ�	���l���h1��	˴VL<ج-����n�t�
3�A�w7�;x��1sADT���N�Z�a��� )$w36�Mrۿ�Lcޮ��X�l��i\헤�f��sCǐ_��twf���YK�b�Ύ^ݡ[}y��a�9���X�*dE�F'pz�͵�wE�$-�ǔ���0��-]j��c�[=}E���T��ݫ�t���u�(Zbs�˫O{��J�wx9FJ�/z!]!P鸓=��Զ(V�["ӏiTwMhՔ�\�N�4V<gl�Ee��컔��G)Z�駐�Y����*|�;u��C���+�������XC�F���m*�;�ܬ�:�e��r8�3B�p �:�8������:�Y��n��f���C5o?�o�[��Ԟ/U�D�*ugR�{L�6�r��%J����n��p����*��\��.��-(8������-�G{̔d�Ko�[(PεAH�f$�u/0��+WD��T�RM.�,�#3��ξ8���@]o:�G���k��t��W0��suwC��<���N�u%q�jѣ\�_r��X��{@�n�+f�Qm�����H�~�u�|�+v�M��e*�Y���?���Q�z���}Z�MeM��|�A#�u�Ǻ�f͹f�bN�t�mKЅ]��A��� ��4�qtI�����*Ν�_nr�j�	�`	:�˚ek�װ�6	L�<iR���=�3VzŋzK������g+D�l�\ۨ��n� ۫�)��X�^r��� [�)�VƎ��՗w�i��g��ٸ��PI;P�5����?�ڌl���i��M�{����r���,�7(����CZ=��N����S2^��uΧK��b���̈fR�;^*\G6��5'�j+ˮf�}�;k��r���Q�O��gwe(�:Y��˥˂#�@�L�y����.��ڥj��v�r�MKs�6搷N|DY���\�Ù�E���i�a�C��s2������뵲k�N��Wҁػ{�v�7U�E/3^g�� ��R��"}h�dKO���
�mh"ɣ�fdS[%QB�1�+CZ[b��S�r��h��D[mJ������G!m(�[i+P�,K�-++m2��
�eb,a��T��3m�m֢���TVҋD�b�m�eeVjm�7��Z�3j�"�UDm^5G�[*�Z��
�TE���m�]��E��X�E���:ʊ�b���U[e����b01�ڲU�(�ZV ����u�Q�KZ��lU-�X�V+l(�ֵ(�2�h�,EX[jV���Q���""&��Q��XQQQ[lPm+-R�L�0PU�P��u*�T�(T�Qdk)A�B��+RZUT+DQE��j�ڭB���W2�֔X��j�eE��**�m* �km�(���-ػ8�AQX��EKJ�+p�U�E\�Tb��QH�"�XV*�eV��fV]�7�e[��D��n��$�۫�i#�gb4��������tYVvV���ǜG��������g`Sd���znjۮ����q���S�X�d���|��J��^�_�#�o6��Q��|/�<�ԥ�/ڹ�.1X<��>�d]�/��\NVy9[>q����\u�8��5�8v
�&�����|�W�_?^�YS;>�%[?���V=p~_<w�~����������H�1�=���R����T�f){��ۘ~�^Æ7��;�|�Ź���^���]}^���^�]�M����BΎ� ��M�]��s����b��=9�>�+"+��!-V���sXk��M�����L�ΐ�!���X��T��5}���_5����vũQ~�.��5�@���_�=�D�8�Wm\0;ݗ�2��L�\sfXw��R�L��LpqՊ�7`��yV;û	V�A��/�j����S�6��� a��~�!������5��q���+��I��}f0FM��ܢ����P���r�g� ��*�]N�@_�6�	�����C�=*g�P�,'C�yW�����	��1Ϻ����#ƣ�����,dG�%�gʀ{��t2�i���6�	�G��9�`�U�}���
�V�_��>�� #T�����j�q�ҝ{�x^�4�CO���v<�sr�dz��]��C�����m%[!��n��2�{f���pvs�UӖ+[b+�K_�>�-�<���̳K�j��\�S�Jo!�y����u��m�zMw:��3�tZ�Ҧ��H꾷�0.q�w�b���C�˺)���г�٦�ƞ��q0��O1����{�<:�wK��l�����y�pG�S���G9>K(k��o�k3\BW.:�c��� w�o	�K�H��ps�x ����`���=>����7b�:@.G��$��������fO��ӟ��*zL���vr��~X��%�^A���L��]_=�Rf�P��{㟞<����xaK��aא�����c�����C���|�IF����r�~U,ȸ��?�܊���s��{ǳ���M�N�#��esͷ]Ss}�v��G�U�q鿻����]��,&���HG�[q�Ϗ��Xe}��ށl��W���z��8��Q�卛�@J�d
���˓�����6�Ճ�a��ީ8vr9�sk�����{�&�u����Y�3�6���] ���C���M���w�h��v8�o8�^����>�b���e)�}=] z�׹q�>��p+fx{z@�r���u�����擛�b��^")�t�������c+UNʹ\�tTDY�\1�VP��&3&��>����	C�
���KB��zn)OL�5�ϟ�i*���v�5�_d��m�m,3௚�W"S^W��ܽ���8)�U&d���P��e[���N��oxR�[�6������W�x�w�D7�k����:��T??dU�L��^L�s�d7~���*�;�	��oٛ�})z��٪)��D�Q���<^GmL�β�r��Ge?q�����y|��$�W��}���pET�`֥��|{�{M�Z��*Y����7�ꪰ=��?��t{���m��ԯl=�SنyJg�ެ���C��i�t��;/�8aЪ:��ٸ==�r��$��f��7ټ��-�hP輪��._�������=;�3����`xW���E�������y�=�4|�tN
�*z
�<�s�hz���f&ڟVz��ݨemt���v�7`pn<��٢�w�/v�<@jH�cN	�+#�@z������s��ݵO���4����m�啥z���^��EI;����dU���
�#�w��R;�~�CO��1x�U�Ω�\���/86:'����t'���_3�`[�� �N�%�:�4v}���3�ߩ�^3�%U��f%�j�vJpf�'GB���.��4;�<���5"���S�5Q�+�G��ױO�vN��;vh�0��o��i`ĺe���������EwK3��b"�&ԾY-Rw�����Ul>�J���ڨܶ"Ǹ{ø�P��X*�s�J�v�*k:�-�Q�2�d��ͧ{�I��e_�b�'`��%f�jgWgP�eo�����l(P��p�Y/����W
�xgЦK"�~��=��Cd�CSb����M�hTh-͛<6=줽U��-@��5��B��>���g�Ǹ��� J����"���������^IR;=9]��	�+��v�:}�uQǧfE�;׹㓓��n4�N@��|Bšŭ���gO��u=���u,�ϗz�y'O��Y��p[ɯ�ɟt�����#�����M����t�Ҡ*9�;eb��/�9�w�q���n�Ķs���VG]������>d��y������j��k�:�dv����%���P����(Ư�(�g"$�.o�@_��@�N`=�n�
�} G9߭�?W%�V������G��Mw,wMV�;ⰻ���NGE��>��w�[�}W�;�YL�L���۞��F�S�l���z��N7����Z�Д]�I��;�d%7����"���Y�&�L�Ԩ�ܨv��7���71�	�ب����-�[x�u����џ�:/#�@l��������~�����=�sva�p3����z�aP3O���9�U��:2�mg�\�<�p=�<}�W�`<�ħZ�-1��^c��j����W_�lس�s�{�(��g��$[x�V�o��Ǧ�ï�k����c��nv4���a��i�rR������y���{�Z^J5�(eg���� &�n��w<{{ʭN��q�%��=���yT衝1<��(?lG���}�~0ۥ��f|�f&��ۣ����><�T�����W�����wِb�WI�D�n	�۔ɻwy�ޡ�"=��??uY���4V�=��*�xW��H�!t�J�_vdn��J��[�ܕ�9����kȬ}S���,
�K^���~ٞ�T%�]&� 8*�w����?^Wd�U�觜��6*�UgH��A���45�L�Tvd�����3���2x�� �7A�}T�7s{�ԗ��'^t�c���>�t8�3;<=�NVfUi��c��G�c}}��A'����1����:�w:�7�=}޼�*d�Du	C߲o�S�?0�t���gj~�Ϸ(�ƽ�Ҫni�;P;�ئ����ϹeG��,ُ}�·OI6qk�#+�W��(Y���x鉧u�tj�4��М���!�� ���9봼���odj��U�i�Ω��S��ނ�7L\x{���ĸ�ٞ�'��yt0�q��u�Ԇ=oU�Ա:�Ǘe1�݆ti��!��G��.�Ok���YD��@�\-�uK������%~��Nۻ3��p�v���b���9�Πq��1���o4i�6#�F��������P淸� �:�Ro�b�!���
���;U��t�I��N�>.�wV���W_4;��n:� ��b%�ҸX��?Ug�[W�1�TC��E^L�d��6e��ucc�e{��f�F���}޿{��`����WCu�� �k@nU���Y����!����v��;�� �L��32�uGg�5���f�y�zzk���YR��y���y�q]�˝w�/&��7-��ȹ���ړzw��^��f�'z�{]��Y}ٝ��˓��	h�.@{�R�xl6���X��_�@�qD���JG�#6�;��:-t�S?IW��$>����#���#��UNE��<{�V���C�{޼�윁Þ��`��;z��� �9\1�}9�w ���p3{�vtU�9��#|�`E�*�rp��}�0���н4��s���UpM(�>��^���䫣((XMp��d
�v�*��n~�;v���6�1��߻D�ޓ&���wa�R��ܔ}�Q��}��|���=&k�v	�A�L��kÔz}�k��L�8�<-��Ω�ulV(��FN�)���lI�QUp�g(
���,ȸ��?�ܪ��7'޿���~�^��M���i?�u��}t\gw��;Oj��A/�ȱ^:׻6�:���Ͳ��px�-�t��mm��R���sTį��A`���=Zo�	�k��������X(���w.���M�O:���:��d\j�8�dT�]�j
��a��S�Ť<z:�;P�B�����������J��8���!Y�z�=��D��LÍ��>:9�k��<�������SL�Q���_ж������6�Ղ�w�7�zsVx����f��e�i�;��p�{q��R�~r��6��rB��,��\��{
��j�����x<[�?�O��Uw�����[�3iɟt�8	�3�׽@&S2����� ;	��1#~f��^��������8��Yy�����O��y3�1d�&s�2�~!o���ηo''ӗ�J��u�EyJ��ߨ�v�=p�\�]����;U�8��.2q=1���ز�_��iZ��}�����+,�(M�u�wOi��WY�TY����7��+��9�i�ʬ��&g=W�Dۗ�n2y�y69�MR�y�u����Vp��Cr�{xyQ\v��{��Ww�'�_C����etZ2�2x5q��X�ޤ�|Ύw�u��__Z��veh�TIU��u#���j��z3!������9sC�{.ǉ����ƽ��}\͞��������.���񆸹:*�9��#��pu��m"��&�jW������0�s\�����sT+L�7�t�*��)Y��_����Ԍ_P�7����C��P��f��n�s�FiPn�p7�8*�q54Ȇ�#�]u76d�Q�������Oqo(~�w߾�,�ܪtE�7C�|%3������V�7�}��%��q����ϽL����U�k����g�7�_we�_[��"�] Ѹ=t��ԁ���&�3�>��=�Z�x�����? Ǻ#�iLY����=�u��� z%D�75^����v�4�{�q�����(�o��=e���iW�h��u��gH]7���Ҷ�C�&�Ts��uz�h]ya?FD��o^��]��;�W�ag�]���:ש���$�<�]'�;�����r�����y�9���uBh��ޠ}>�[p�r}�\<���o��ٸ�`	�����B[LWZ�ݯ�՗M�����܊ow�A��r�qL��y�Ԍ��^�v{�^>�؍.�:ޱ�/HbW���� �pz|GGuh�r9exUǻ�:o���ӑBpydu�O�zj�&}����9׈hM�Uv6]
�F�*�1ޤ���=�7ݻ�ޅ�(�>�2{��`��#S�<4]��N5�r_��q�4����S/Of̎ۈ��b�MSt�NC�+�}�(ƨ튦n"\�.\k{[�����Ύ������;2�J��0]���� t��Qެ4�X'̢8ܤr�`-Z��Q�zF&��(����j�j�)�)O�m��� �h�B�'�8ޱ ��
�����n���Ӥu����]X�>�.�8l��E[���������ƚJ�7� <q�׹�INN���;��иɝ�y3�vmXl�F��Q��M�k�:�R8�=qՍ&����)uӊ�F�s��R� h�T��`\fJf�ɖ9�<ƺH޹�=�Ƅ�wt�m�U���r�%zMoh��E�q�#��A�@=��W42�_�T�3���͹����!�ѐ�W��x����m��j�1���������S!z']�f@6�q�ܦL��{]�`c������q��]N����u�7{IF����;,�yT衑�̏��Ǯ���V�I�2���Vg)���x_{������"gԦ/���g�k;2wz���p��j&xR����X'E�ط�F=R��0��h�f�i��T)�xR��6zB鿥O ��2 �w��xF?���\�ot]pnx�Tg��_��y��5/Ǫ�i�
T%���h�>�\T;�c�>-;4{*L�{}���ɓ<��vEڝ=(7د�O2W��1�E���c�q�Wt�$�}���O����f��\���
�|��<�q~3>�S�������d�x�=��F�� e�D��T*9ϋ�P��1`��>���M�Y��-�uj�	� ܩ��j�ód�J�;1ӷ��Z��:ۺА�7����ī=�ig��7���z���	Y7 ���=��-y�{-�}��b�a�n	j����;$�����QN/o����2�mǹ�����O3�=�����Gp�~ap����2�Y�G�Ł�n~�4N�c:���[~�]S�x^O"���p4�����#�Tz�r͘���·NDuI��;�2��%�c�<q��y+���c��.���u�Ԏ����	���[�w�w��~F1���yATW�b�{H�9a�'e�=�B�ɟq���;ڐǯ�ׂ�bj�3˲���E��2���8g٫���3th����WM�NV}�q�W���xe
���\t��V)t�V�x#b��8�s~k��:��R;�Gmf߆}��+>�)�9���s�;\}����_�ʆ����f,���{z��z�ql�9�/�M:���J;����<����e��q�h�$�X�M�=���9���6�v��׵�s�#Ǻ���)�(8�Ķl�h�U"�t�I��Ȏ�J����,OFKe_ٵ��N�"�.�\�6;�TH�5�1<;�o5,4�z�/V��]>'mY�y�h�ЯJx�����X����^/^s���$!$��	!	'�	!	'�$�$�@������$�$�� II?�� II?��$!$�	!	'�$�$�؁$!$��$!$�����@��R���� II?�HBI��BO��$!$�r����$!$���e5�I��'
��!�?���}����!��x�*�(����(�R�$�������J.�"�!U
�`�Z(Uh�D�+F*P����Q�¢$�$%*TR��(�"J"u��"��%(^X*TXΊ���2�kR2�6�Z5Sb�M%P�hҢSX C� wsRU)� ��  n�  ,��i`����j�aR\ �X�jK����v@��A�5��� �B�TJIp`ó���Jd `@�B��i�X jQTT�i����[Z� ��
�@P�� �J ��b�h�QU6Ȓ�pC�6� 5�B�)[b��S[FT֥m-kՒ@5B���g*������Rm�2��1F�4aD�, �R
���ذ&��$�U@��ڕ�iQ3j�T�"RR��Q6��UUZe[m����-6�T��6�6QA "� ��&f�&�-P��YljZh���0�"E7y@ @ D�M2�)H�@`�h�����{FR�� �� �0��F (�M�ɓ"4M����h��f�j��	J�z�      �12dф�14�&��I����!��0	����9�מ����сKa\q�+�S�GW�R� UA�"5AU`)�!EPF�����/Տ�������P0�eA&~�#�#D�*��@��@�u�/�s������ƻpT�F��&��0��&��S��2YJ"��g��˟��)�^_3��&��h�B�N�Z����x6�\VR���Ԃ%���ӻ��u�o{/4���-��0�Z�O�a�Np�j,�a'xcB�:/P�b��]��2��83^������РY��#Z�6^���z]Q��1O�۩Z�Y�l(��k)&��)��!�vh����b�Y�n�+�:�g��̥3����B�Kw5�
VeU�*n�D0��`��r�eQB�Ŏ�Q��4�j�q��BЬʄY6h<"���Q���.COAb�Krɦ��(3DP�	��f�VֵT�h.�iU�fbR�[x0���?H4�+���5+$3Y�t�8��5�Q�w�1d���-�qeU��Eʤ���-�{
L�́M;D�u1�Z����kG��[�PNl���D/Zs^�eM�[�Y�(�v�+���H4T�v�%Ǣ|�mhY��j�6.�;�
�Ǵ�D�@�rb?M�!��x���5���m"��BO%n�$Z��3b�r��č����X�:���=����p���ۄ���zЫ��p�%f'	Qa�L�f<.��a��'c�Hhd�3e���Ĵa߱��6�hLz ��cW���>�=�W�t �ci��`����*)�$�Ra3��:�=8��J�]�i�6&Y��H�p���ڳ�-&�WX��-ô��Z8�Rw[I�`t%M��Z�ʄ'�,�V�&mQ�t��(�V`�KQv��d��P'Zo�)m^Q�u+PR@j��uBr�x�ۓ.��^��li��+��볆�TBh�G�4��)�V$�n��&���\Vf�G(��
�捉]0��CT2�v�jA2I�p���O�$ݍaܼ[ɛ�����'�ңd��1nǚ0n��b��&���n�Ef6��헲�D/t*xN�����(n�wQ�,@rc4���h���ЩXŹ+�W��P�mR��f[���ŔZ�oiͬ�x���7�f�`ݒhX֒�Ƅ`��0
]`(���:t��{� ώ�h;34:Gkm6�h9n�wz3dos��b���;�@䙍�-j.�*JXN�C�a���mlǤjMbL�'�.�Rk6<@�ͻ-���%�٬���3�/TD⩒d����.UC��VU�g�*�L*h�LpP��XU�[�A,�p毭��Gq�w�zٺ˻�3jXN�G��C%���{i�N���M��+E*��2���j��:F�	�����O�kM��E'q��/fZTq�Wс�u����P!7:�m�E�d��[W�P�A�'�ú
h����1l�t��TU�6��;�ɤ;kw]e�0΅��q��f��&�o%�# y��=if޲�VѠ��'��61�Fƚц����wT���4Q4fF�(f��Y�s��Sx�Ĳ���r�^�G��L��R��y��{�ս��]���&&��9��h�͈��OvZ,��;+j�8�b0^�2�1�s/1Y;�kM�3r��b�����.���bԽ��M���JX��g4j�i9Ev�ʺ���*3K�UAA;��
&�ց�ۧV�/6�<c,��J6��<Y���&��iܺ�04�i��[y6L��ޅIQ2ܹm��h��2s�z���
6��Fm⷗@���)�BQFr��6�Ջ��"(]�&�v��[k��BkX�ʂ��&:�*כa�[�Dha��܉a�V��E�wXYP�ݙ+ �uw�%	q+FE�����,\6�SSS���*\Fve��C�Yq���&9S.���w��(�mV�2Ӣh$���k*Gj^e	�De�����e�a�\u�r��Z�WIC��df�A��z��0u*�Y��#ݵ
h�V�iZ$�˷Q�{��:�:�]A%��R^˗f���&�����2F���
ڳ�	��fAm��2��i�Y��f�hPenbh��Z�pa۽ݑn���JЉ�D�6/O�ݹ[��ZƳ��X�(��E�uB�,[t��r�r��W.�VN+�,80�;��+2�+Z�o6�ڎ[&'��.�ޓ������!I�{n�.g��֍�b���i��CsC��T��"�0м��܀�V�Ͱ�їDj����.Ef�K�e�X��!��%���d�w��%�cF��@��5u����5�h��USM�b�
@ӂ1��Q�a��ƢK+����VdYy6�B����(\Yt���Q�dU5r(f4�2+H96��B�3�F��,�/.�Ma�pe�nAa|c�7P�s0�+s�p�:.ܴ�K��"쿍�cdW���BvZ�m�*����@����)f�Z��d��j����LU�c!�nf��KtUʥ&lw.�i��i*8�+Y�A�3�t�w�L��mӛr��֯-d҄���#7`��U*f�f�:Fn�M�eK�S��l�e�ˢ�)$u��4[�$;�b����
�"7h�4���m
�z� Ӱ�*1�����l��G��i�g~�9�2�3V�^�9y�^�s#��pF��ߔ8�gքӛ��b5��˿�4�9w��&4Б�n޹Y�����Xve���1U� 7E��)�w�F����,�d��Q�ńAAl�tCe��G	��MX��Y�n1V��`ʨ`G^*3s���9Vh�2;wA�l,�c̄'����-�������)�ۢ�J2��m)n��Y�#O�NƑt6�׍�ەge�
�	�IM��D��f��L�'�L3	�ۺf��F��ݒ�!ض�D,B�M��Lg]��b�2A�
pn���h�����LR�)	PڼeԔ3bb��
��f�/PL�V �d�"���y�ina���x���6Q6�ڍN�#M����0�����I�ٮ�d)p]���$��[�a�x���2�6��,)�Ǎn�y��SHjccS2Y��V6��3�ٺ�&����,��j�������x�����F�`��&،����̚��,P�����i}�b��l2ˠ�x��u�3f{M��y�j��h�Ɯ:ĺ+�]ǂSѥt*�]cƥ�O	�>gkxa���{Ֆ*-�Op�:{mn�NQUɺ5��U�ee��N�`=i`�EH�H�t�1IZxW_����@u���
Fo�ΡZ[(��Y���`����')jw ����N�����d�����%�틻��/��f��N�V�wX���+�"��='vYڕ���rk��Q�j4�dͭ���M�tc+'v�̡�Վ�K�#Z���ҳD��}W�(�H��&����,���m�{��6�Έ�U��'z�g?���n��p�\]�S��5��E�\�L�.N�pd�viu��&JSI�)Ш;	��jb�͐�b�Ow���LL� �sN1��Mu>��\��t�ݞ�ԛ�Z-Lzen�Ү�FJ%D72��7���Χk�����l�v��tK�4S�b��U�����r��3�Il۰s(�E�Y�hM�{��M���&��1|��i�&�I�uW`�;8�a�>�2�r��!"w^Ѱ��}t�HF�����F�U�iλZ��z���w������{,G�.�94�x��{�gIZ5��:.��;ӱ;4�a(��]r��]Ν|��7��o3t�6�A��qgp�;$�S��-O����2b³�e�]9���6Z�x������]�'�1`�2�l�jq�t"Be-�-�I��oH�����N6���F�wU�(Ζ�b�^�1>Ⱦq�|<������7g6zD5r$��P�L�N���/k�)ud�J ����fѰ�+b�1�e�3'`xPQ�*f�ll �8ú:�b,��k��J�h��+H]��r�=Xh��Ζ��#��.�<n�Z�qT̾�n뱾+�U�z��wv�����8*o-�ݹ˅�Ⱦ��޳��f)
�b���DTs[i����N�zy�]�<�br��N��:�3m1m�ip��m_9ݭ6-}�+����W���3I¶W�J��7��Y
2�d8��ӸᶬΘo�p@�o2m$w}9l�{�I�w�.�x���62v��(ֱ�	.pݗ�`����<�ځiL�`W�1�{�ɕ ��w�caiK���U'
 
���]=�����`S��W�I�Btxk�<���6R���q]E�{7�]���Y�
��a���Yu�ʓo�>
�B�q�s=������U���z�v����:u\��dyWx�K����r�&v,��I�AZ��s�=�<�-�����wO���t�����X<3]#�7n�.���j��n����Gab�ss��l������$t8X��V��++�2Ec�����'\�C�fB�Uꮷ�D�b�l�≻������;ϫ`jM�W`<ȡ���},P�]\HW�#��U�]8c��C��"e��UB�R�\q7Nݾ6͎��D�EGd��y<�g���X��Y�Q,tɬ��+���W,�w/k��N	�sm���*�'#9�nk(U��{���[��.&d嵐�j�⓹����TRfk*ͳ�-����7�?=�E�4����k��V\�1��Ϋ6��NPߋ�]�z����T�,(2���4IMe��Mj�5%4��r��E����ʰf���N�}0Ҥ�B��Ɍc�r�'�m��:(�N��f�kcL�z�*')�,��ֶ�7���)��o,�C�*��KS٩h�)��E�|��i��T�}�M�5�[�V�56�yc��4z�N�@�&�bT7Zz�ع��;�+E��PN:x�DO0RF�XolX�j�_g�`.m�RG*�I�1KW��"*�O�,�d=����> _e;=4��as��,�h���Q��xI��{sY�]�=
	�C���N^�*k}�0��T��#��(LK��2-�)�nl�3Ee ��&���Hn�p�&8ݥ��-�8���^ő{usұ?��[y��R�Ls�x9w+8ݾ�Ui�f��X%ެ���3O��`v�i[�Gx�e�!���V8�R7l�gou+0KY�/��`�mӺ���t���5�� � �4�hd�eKz�v������ZC\����Qq��-��	����}[����{��J��Ks~ӕ����
�@��VRwj��������*O���U�ZÇ�����J>�S���:&� a3h����I�v)�������8���MQq
Gb:�����;�V�Qy�ZO4�on�>�HG.o"6��/����^���uʱ4�5s)vA�s �9��`�3z�k��=f�'�� ʛ�S�G+�1�A��Ϻ�����lֵٽ3k�{/#��k�'^��RR��겑,�M�%]��J�nX���ͫ�HD%�굟.��lN��&����n��C+�1�o��{{������d�L���⽒�� J��
���m)',L+�yf�dL͓Rn�=%�]�Bj�Yۘ'j<���NIr3��t�mj���0ѭ-X5�\���A-�cjuW���2������1�*v�t�,��',�z�ⱗ��.�;(��&��4{�ǵ}�u�OP��8�<�,�|5�(��,�����4��u3.*�:�ګ�Z����-/k�¥����U��ǀ�������}8��Rk�ݫv�N$���g�.��u(�6v�Hyi쮲�������;k7sC4�)Bf+}��Vřm+��텹���e��f���ٲ�CN�(�@UY��t-���x����q%w�B��q�u�R.?��.�]�+�#�wԟn���9݊ךּ/���Xd=Fs��I e�Õrs�<��x'[<���j���P��l��w��Qa�sS:������IM����$��RI)�қ}���F�x�}4�yr_�\�\q��u���Ţe!Q-fbםhQW5�v�O��1׍u:Y�ĻD�E໋JL��5�m:��	��z-N���8�(Y}�dJKQ}թ��}8�6U�H��+��-I^�.�4��<��
T6����C�ί��9�gJ���TגA��k("��{Q9���y�A&��4�ٶ�mK쏬��[���GPޕ������T�jv1]����	nIQ|El��]�B��[��{x�r��釸�.�g'LT��=�&��"1�B�v�d;%X�	�X9�Ƀ�Y�T�5n������Ug���þ<�"q=�gb�k��EuF�sDd������NǸ{�35�w��j-5�;����GwI݅ډ`o4�Ypϙ�o���Q�/��7�I4R��wۨ7��̮���mpYۥ�7��5u��jQp���Ǻ�gn��K.�h��7�(F��m�7xYO/����AH*GD*�e��B)�s�J���������\�s���go�;E��͋��wrWA��B]i}�̷ZVGǐ1M�J:��ohr���
��]�ji�ͳ�,�:�l"�V����F��Yfd?&�yu&fi�r���Bp�&��U��]���ؕ��bv�<rs���igv����7f�F-���ﺄ�����d,��ob��]���$5M�ܾ	\Ht8���jԑF�6��|�cH>�ɊWf���Ε;4ZMHQ
�9��Kәʹ��敧��ŭ偓�a�ٯ�Lù�m�
ϸ�I�V��4:x��p���2�o[]�z&�u�?FQ�CnB��C���A�U�)+/M����ܕ��R�� �U��q뿐����l]�K��^����tvw�� +7����oNn;VVY+3�<'p��$+{�+[BAٕ��5f���Փ�>4'R��F�B�*�7��-��tl�F���Nvf�'�&Mv�H��Q�B=��g�UQ[5�s���ٸ�%.qˆf�Lc����."��:���=������&�m���X횷CW������`��Y����M�o�:̼J��*�A���I���&W`��N���	(1I�1j�/Eœ�P��*�}8����E]c�zm�k#lUl�3&��4.��[��MN��;���+O�0�K�Ak`���ޞ32'[�7X�)kW��j�g1�<BD$���Q��㯵_9\�����g�rK�k�7&��ݪ;	�e��.�lg�rY�������ٗ5�mT�m�\�+���q�WV�5܋�}�1�͑J9;e&���͗�Ŕ�[85ևqȷk2\��h�ҳ�e,��J�+�Ρ����p��l�5A�b��zT�^p�1,��},���[ǝ���-7ʝ]���c�,����V_D�{OZ�f�DD3ٕ +o2�F]��:����r�w��&��/����S{�7W)vR����g�:����S�0�OS{fT�|�W.�w�t���,o͌=9n�[�OKN�[��v�Z斕��9�����V�b�=T��,Ud�FS�We�nng�Х�Ŧn�Y|��WbFt�|@�o�+�ܴ񹴥}��E,r����ٴFʉ8�6�^3�Lv#���vwF�X@4"c�Oy�F�e�����)�\�N؛�X���uB�������IB��&Ջ�r*"��2Z<x�����]MZ�
��9GT��,����f�oX�7�hj�l_20�/�N'�����ږ�����2bO*:(�P�Wq��ё�7����5�.
N�^�:NABGP'o *���.S]�馸-�M�Ǣ`�Rx��Kwy��]�Lt�|���U,�i�F�5d�U��~��+|z�3^��E���=�喐2h��}�'+&y���������f����cF�.�˱r�FnS�Kt�8 f�dC5ܭ��\t�kW*�s)�v�Į�_e�mb��+����C��դ�|�K��+2���ٽ,�,���M��^b����ck*�2�M{�gL���J(.jQ��<�˪����w:���U�X6�>���b�|�nn����R:k�[+�ػ��um���*CMv�m�#��W�CLx6�<��\���m7� ��eq��Wq��U^6���l�lqif32V��T�����]N�N��"SS�(ҽ�!�8I�K$X�D�ꕙHI+�]D��M#����[U�º�n��A�ٺ�&Yޘ��sy��{�[X���K��xeh�C$tn�
!]��hށA+Q7�"���՚��R�[���vZm��318������0��ׯ�1*�󚰱rn�mc����3/�{_:�*�)ϫ�4&������+r%����W�;Ei����p�.����M�7�ӣ4�2)��5Un�#U�෦�c����<_[�Kuy';�U����U_Y�������L׌j�żց�G�T���P��n��}m1&l�彛��Ulo5αU/C�2�d��W�L�;��ڤ�2���K�e��T�T��컫��c�g����
z�i���dO{��r�Z�����?�[�Em��&e��u����˹�y0< ����I��-�vC�q��L�E8��Mϥ�KV�5�7>B�ǰ��s��u����?<�u���"�c�fJ���n���#Q�뉴w_کiW�o�Y�d��b�t�.���	b�R���\o8<����bW+��$X�²�Q�e� ��Kջ��!-�ʶ��	AU�c[r������5����f�yH6��Ƀ�o'pĭ���s�6��� m�:Ɩ��T���;�H�*B�&���"ee7Zok��Xn��}��0�����(�p�0臺A�m,j,f��:�X����F��uI�.��)�9N�5����0k��+��wwo[�7:��+q���"��o�ksqL/apr���a��A(+V���4��y�<՟���g��J=Qͩ2r�o%m5���Fb�3�6��2�Q��b�Z�7�N��V\�Ǻ})8/�t0o�:r�e.���'8��D���{�6��;��q���z�	�f��.��e���q�V��CYWWk��0QP�ٗ��QrH��U"KK���KL=LfP���k8�nTf�VѪ���h
���B�I��viЇ.�xaؕwJ�[��S��y���]��{����$	 B ��$:�=���?��я����7]k�G�r�:r{6�e��j���4oo!�����m7І��_���o�0x߶�����32��{�c`:��z���=jQ��.�R��l�.�C����]�-N�Z�ݯs0���D���9|aж�R�#��P]kK�-�%��-|z�쮲��wFH�CV��gX�,��t�ޮ�씖�[�slGH�˺�Fʿ� �_k���%0p;U�߸#f�j
�Gq�n�Ѫ�3zkZΚ�h轛I+���Z]ʑ*(��X�MN�R!E�:3���L�m���벵��[XW97���sy��%hns�c�k�,R[�m��=A�}� o��k�-6���V��r��ZX�E܎�����#Y���9�Wz���?gH$���5+`�F��V
*"++Eb�e�1X�,�:�[h��/V�ڪ�R��+���4�`�"��j��U�*�̷-X#d�̋+S���5�mX�"�Je�,̦%D2�ulX�������*eT��Q�)J�T̺j�R��"*�c���J+ձEPq������-�,��Vez��?���~��p�z���U��Y�=�EF��ɠx�j=��M�������c�Y��W1-7��D2���~�6(E�1�V�Fj�8��xwkFҽ�u{����dm��(0�ќ
�����v�G1j��0]���j	��д�m]��԰gIQ��V���F��>�]$V�T	b�38��=��zZҤ[���O���n�]�Uؤ�JvA�n�w�R=�ʩ�Y �G�,_���8g���
��0*Q�u52]]]~c�����;�2s���6��}��;Oy�v�%,̑c5e��tَ�Ě�B&�F[���ozox����(P"�П(��ip��Hq{����噺W�����M3N��F=�w���=R�������ٖ��x�z��@�Y��f]r8�{!�&j�<�4��$"�����n�Nm���'u��j<���Ax���)p�{�_�f�z,�ɍb�tr�d=k�+�Ϣ{�����G,��|�to8&��d��6���}F�pKy�P����r0��92;����J�����9n�3�!mǌ��W1w:ާP�r��r��ŉ�nur��d��F�\34�_��L�އrC@�znꋊ�B�#;˺u樓��:/��\ؽa��]�S���'�Ǟ[�.d9���D�t�C���|�bnJ��-,'r
T����űm�۱`�C�;5�gw�أp&t�2�+�^�g�᝕+�� w�3t˺���]��e�O0=9���Pl�v(k=�N��O(VQ���[�����٬���v,�\�H\�5ȳ��#yn�]4�j�S�p��Y���;8o%&��Uٺ�fd��y�z���ҩ�������[���V�Nk��L�mb���x]�XUq(>b*Et�mS�����%��Ы�%=ӺOOU����է�z�� �c�g�ȅG�뗵�P�v� �.�|GD��&�{�HA�爇�6G��Iv�M���!�Ү������Pfe��-ǩ���-k��4�UdR��:9�Es|��å�cs�wQ��wQ�Ӆ�k��D[�oM��s{�f�`ݡn�ƨ�ծ[�d�秦om[�^�N{m�0)��C4����7����#3���J��<f�8yZ���[��P$��c%`���+l�O&b����V��y�u�΍�t��La�a	�uk(H�m
t�Z�v���e���T�@�vT{Z�(߷Ͻ�h^O"fb������ܾ��MO�ˮ���-�})���{t���.�Ѫ�#���k�	]Jޓk*T���ڏs}ׄEQ�zR�Ov�K���D�'ax�*{�^r>�`u���6��F6";�Ո����UG�<I�2�CoޒIqAʯ϶q�@��3w��Cŭ��C��Um
�5e,�<�k֯S�^En�;(���O1�ފ�1�4��؀�r-�ȡě]��Lw]mbF����xX\��>��F�g;�+�3dE�x^`5�e�<Q��ro]�5;]Դ^��z�-�s�{���F����֞����ZVr3hf��-��^��3n��y���0'��{n+!\�f��_�
Т�`4s6��8t�=�/���f��F����f�K��3�&�qۭt;S�\�+�˂!j���髚�����Uc��oa�5%��#Wk�w�E�e�Of��"�5��n�V�Ϟ�5�-ڳc�rU E�cvlZ3H9�N�*l��:T�wON�U詬�q�͏c�Q�f�q����^�˝���VWhSd�{+V�g�ni���K֏��'�g��n�Х>�n?zΊ��k�>�7J�W +������*��]<��P�X׎M�y�:�m0��=5�|���ޤf$�wzzh�>
-e]Hk�=o<_pv:�U$Tx�����q�RY
ƹ*�jB�3�@,U���3,���wo7�]My>� v��.t8<��f�q�ɰwd{�g��nK�=�ß,0z~�a�/�.�Y�������Z�5+1�׻� �=g���ŗ�0��'tʫ��D<�1E ��	�F��zC�.y��s&i�%�ų��I��§֦,+���m��;Pm�(�:ൢ.����[�-�s��������㠞��}k৶�f`W�!Q�epL.A�!z��tXFFU��3M�b�'��*}�@�k_��<}P�W��bH�b��Ί�����u"�=G��P��Ӹ����a��,�N�@���;�T�g�p{J�].��Ł��I��v,�.��u�^kXB���q�<���&�7h����`���E�软>��y��JLHz$�m���G�=��� Ϗ;O��X9��b�ͫ��b�R(::���w�\Wu���llW=�<~�9t�9M�m�ո�<k��/�Sf�霂�J�vNZ� �J)��
��j�O�n�����6cn��ʹm�>�'\\�)]_�I��Ϸ��^��P?+ȓ�3�����m�AK�ѣ�zG]�Ka)҂^�uy���j����UXjB��>?m�m5��S�ቴ��2f�%v�Ư;{:&W|��G]|089��v��e�y��a��ڼ�^×f�izds{�k���N�޳��nj��ΥRL-����JtN췢��3/jetY�*�/�L�,��ע���2.l��y�mq��q�ሧ6ض���O��L�|7s!�L�]֒ݐR��w�u��G;+�[z�C	�t�wճ����N�+wx:�d0H�ٛH�U�ӎK\{'Q�uZ���-���GҰY���ⵢ5]2؄&�i��]�o���6k[����_��?+9���&�qw^�zi�#wa�E7�a-*���D�i��X8u�J��RAt�E�����g�c+�4	E�U���&��1�!!�Y]E����R<T��ʆ��3/*W�ID�)ZJͣ,Ɏ��w2Jܵw�fI�8�nf9t�5��f�˗tbX�a��a/�Y�r�݋��8�c��v��o�2���.S-����ЫV.e+E��C�:TH�/��ZO4��W���ǶN���ct�Y�Š�u�j��8��,nx��zjѢl&�Q*�C�,��T��˶�$X6�M�)�6p"w�q���hJ��fl��-%&�?YUF�5J*�2�mA@Q4��Ī�h��c�QK�S4�L�)�E�Ki��1�P�R��U�cƭ*%Lj�G-2Զ�ܤ�3(4mUAe��`�Z�IMk�**�V�D11Km(�V�Z�
�5̙��B�8�bҵ�f5���E�s2�r��*UI�r�5nf&2��hTk�,CF����J�B�m��JYJUX�[cYi��(��S5u����m+���s3-�D)B��[lET��Up���DU�QF1Ls3
)�UDX媊��|d9��T���nb�7����ͼQ�*��XճN�U�w��3X�cz������Tf9V�+�=R���W��Iv*l�q��a�W�~'�H�;ٛr(���d���;��>Y�1��Q�k�1�q�#��d0���e|�k}�rɫ�#���hÙ��O6K|5���Q�MEp�}���H 0��/����n���s���f���Vdؼ�Φ�s�-�ʼR��(ۜ��Ezn�"��>��VMOʱT�F�~΢�hejvFR��D��nQSd���񴙝N7��#�S�����YN�a+��%��]�α��V@���U�uj����zJ��>(�A?s����.N�O!F�s��{\�Z�>ʚ�7O ��9���lq�̃�i�9!�t ]��-R��&&��x�䝻A�X��xrr��N�=H��Pk&,[��h7�p�Qك��VՂ֯A�EL3C��X350�[ì���㱤�����Pݫ]�5�%�'`(N�;}1cHHe�Fs�yt������17I����H���^��A8^�Ouۖ���:�]���V���>��>���2x��B�L��$1ߞ�����k�}� |��ߙ!�&�0�%d���ORN>��h��c$� �$�$湾}+o����4�M�|�g�$>��m�a����8�q����`t�$=a�C��}{���]s���Cl���I�N0'[��d0��	�|��8��l��հ6�]<뻞����N�|��� ��� t�0�%gG�$��m&�k�@�9I���?_uÝ?o��<`���$��+';@���'h�u�IOP6��Ӵ����f�: |��=�@�0f��!>I[l!�Hx��"��Ω���g�ί��i�t'�i��M0<d�$8�'��H|�$�Oud�T��}�����B��u����c���1���S}4�u�vwf��o7�p��E���H��-E��+�pK�VHI�
��/w���鼱r��_;��n��Ї����@��!�C'���q8��!� �%d��$)l�I�u���<�xs���f���I���O�Xa�!�$���'l�Hq�$�L<@:d�g�s]I*�a'I=I8���!�^����o�XN �M�:By��ޯW5������o �l�$:�q22t�OP�0`v�m3VHS�t��Đٿ{���^���ē�=9�I��"��$�M�M�+�'́�!��C�)'h���w�_~:��������� N���:I=a4���$<����6���M09���o�}�>d�	 �䞠zεH0��m����VI<@�ԜHv�M{C�����=���z�c"�M20>�	�!��2q�J�7�B`v�T�1�xmy�~s<󜐬��IS�úN2N��C�xȡ��'����M���<ל���I>9a�!�&�C�IĚd��i'=�C�2,��P8�|�;aý}�߹x�޺Ӻ\4[-��0!	�3�+��O�οw��£��~��vNS�i��׌w��bq��Ջ�.�N�22bVA�=��ǽ�B_l�C� 钤<d�bOP:t�8���Xz�f�ϽÙ|���9!�N�LHq�d�ɴ:@=Ht�m$���R|���2�퓶s޾�{����<H0� {9M0=B|�6�n�,>��C9`t�d>d�Ci%���v��7߼��I:dS��� mY�N0�n�|���M2��d���z�b�$>`������;��H�M�|���3�@��I���@:I���Hg�Ho;�.w���{������!���	ěI<Hv�k���C���&��x�q���百��7$���n�tɞ�'+"�bd
!���m:q�v��H�\�^����=�'��l���!�!�;I�I�L��Ho,!�c'�6�c!�x�q7�����]}�~}��}`|ϒO�Hc iS�!����x��'� ��t���xs�k���y6���mi1�t��$;d:d��Cl�זHq�l'��v��xǣ���5��E|�5�[k�,:R'f�"d �,���I:ֳ��}C9�9��m��p����W�hG�	ػ�}T|���HI�T'��I� �$�vHwl������ q���dRM0<a/����}o��$��0=d��bI�!�I*v�ݤ��$遜��&К�@��T�z*���%� 㯜��TVP��]���R���f��'��%1�EZů J��y[�V2n�m<)�dL4���M�c�[�]�M�����<GL#�ݳ���ьbd�7׋<`��9��b�;*Z���\Ø3��'���hM��־UA���\V��~�2�eZ�H�$���9Y�e3�^
��Nf��D8�Ūm͉��gV���}n�iG�ވ��8���^���[��y4���%�5��Iy��$qr3�o3�V*����Sv������2U=�F���1E�8�s6L�u�h�,�Z�=:af�A�f�*��y5�c�g�6��g��	��VQ8�Z.%���arT��Wթ��V�}+W_Bht�ʞ�o8�O�-��tS�pM���H��S�q�qZN7����VVOsۼ����C�U$���e,V�AB��3u�Ң�-Z#.>��=us�����鈵����'�7���k��u���b�n����*��0���Y%�L�v��VtiR�V���0�,y�s��X��=���,�7��0l�wVy
�9[h�}�D�!B����܊oC�I�<�E(�*���u��m�,����8�*��xy? ���M7��6��a��Ч���!_s׍�8-�ʌ�[�h��֭���@Z�)J���|9�_�Hs����ĄT�Ӣo����着�����E~C�'Ҭ2��&��q�,�k}s1����L����আ���>��0_$�s�����t7�v��7�{f��n�h�[��v�n�B23�:���֍/8�j�0bt��^KY[�o7���͜�']Hk/���	�Ҿ�3P�޺�����Xy�EMĝH,�^��>�����[`\;�˺���j5Ԧ�Ӭ�nx Bق��u8Iy�z�lT�%D� ����@p���������~��T�R@㉙}�,�A�~��z#�4�|��}��r���%B`��o���~y��xZ�>bj2+���P}1�[�#쏁��$��,�UnZ��F���7���LM�ڛD3=�y��S�~D����g��Y{N�M��B�Z�ܞ`�\>v�Ue	YR����YY]����,ka���N���F���QX�\�u�s�b��F�5U���:=/jW�����׶x?߾�ImK�_���z��K�"T�A/\{���1c�)-C��
�u;�w^Dhu�;]��GκU	�����,K�7IT#�=�Gdwx��hN)v�n��TyEv�IWZgl\�ġ:4\�縛9s�UxY���/`�S���ًP�חƟdS,p5�*��Uja�\�5�ȧ.�{�JY�x�=p� �u[�Ў���X��Ȍ��N�4�-Ϊ刕�gQ�7.�<�L$�ݜ*۾����'GoN��.w���B�e�F��,9��Ǡǳ�˙�a֤��}�ԝ�ۥ����iw]q�Ң)Fw�{#��U{Vy�6����;\��zo/r�:sW}�{��Y��Wӆ`n�d��)U���-U$~-&���kU�8��VӤ]���O#6K���x�I�Ue\3ec	��)�sC�e��VH6�U�w���%��Utگ�wp�%��2�*���YB�V�x����be[�F!P���1Pa�us"Yp'�,�YzJ�7�z��%�dYGkG�vut��ՊQ�2�`#,9,��:��a��S	���}J3P��YaU��(�D鼷����x�
�J�7�p_�*��ĵ��c^���OU3YGX�C���r��2Vf ��&1�1~��cG����X�ZU,e��T-�mC�b�*,Q�Z�E@����)��4c�lQ��&�p�eU*�iD�V�e(���AU*UTDETV�Zc��Ƶ
�EJ�6�Z%QQEUD�(���	mV+X9f��t!el)h���m��V�ʫ`TYTC�u������_�w�����9�2���+i�{���H����������R���C��UF%�D�����#7X�v�^��yՋ�:���7��"s��<���y<���u�৖j �.�*��3�T��+oJ�q�/�X���{�9�l0�q8S����#�QN�Z�^��h_��7.N�C�M���ƪT��5��Y�]�	�o�6��*�2���=>�T����C��Oᶱ/P��:�:�\�^�w�c�%���f�s$�c�ˬ\(9���tÀ�S&�V��w��N9�����������_#���VB7��c��X�l�Z�Y���U݁��T���Ӡ*����'��3#;��z���@k�<\���Ql��ޜڳMfD�@��CP�z��'�a�<V�3=ش�"M����Z�ë s�ʻ��Bh��:w�3�k0�X�r�!Dj���y��8R^�G���E1��N���q���hq,iN�R���6�֩�E�&��b�D�'t�2�I����K��%S��]r�(+�7�>��G���~K�_��<D����Srcr����[]�lܪX�w�非�~�A�C9���L\�Cb�,y|b�HX�>~���!�X~�Vr!d)�j��U������km����\F�/'���4�.#I1�C��6�G�V;�g�:�dQ�$t�¹���1�j��[pu���YÇ�6~V��!L��8yi����U^�s}��s����6�
,|��=�47������A�qx��k�JXF�p�r=��>�&_;��R�d˘�FGMY�h�E��|6�{�cyn�v�뵧���7lk-ɘ(�y/Ok�/������D�Wt�R��X�9���j~D��9����o���g����|��-u5�rq1�Yv�CG�Mt��XF��֡yl"����lA�V[^,�ӿ�c�Hu���S����\瘿T����S�2�#��UO��h�:�3;3O���O�B>6e`�G����n�qb��kӱ�~T��qY�!Y�C��j}�&�#�j�6/�Û��"͜?O!�Os��:��X�V~Ը����N����G�Y%R��2��;kk�Hi�5	���0אŝzf�U���G��y��R�a���G�Z�"�W+�[���罆P�p��Q�܋�0b��[�}'<�d�5�k-c	:Quw���B�֝H����=�$��?ؘ�Ǉ���^-!�8����El�s�6b���A�13�Idr�'*2/�+,"��u�^��g0͑�p�C��q7��h��f��N��}>!��2�<p�5e����cݭ_�7Uy
>EQAyxд7T?bɻ�j�Q�e�3��)�,�GǊ��˫#��g�'�*��3>H�_ �XCC� Cԅ��6Pͺ��P�mn*9��^/��YR%�*�]�,��O�Ŧ�gs�j��+�ݱ�d>�.�QC��߈Vn���A�b����|���֞P���^H4}��]���*�� �}��i.O��yfu5�u_n�����s+��&�Q}$���s�!���>zzOoz����{:x�եyV��j��4��l6�?y!g2г��%e��K®f�;���b&�C㦚�?�za�V���J�,{�MX!��zg*9���5�ʱ/G۩�A�htÅ^r��A�q�p��5-x�ds@^���/�~�x�}�^/�^,�8y�%��]�Ck�W�#�@���_8�?e�@��儗�O�M�'s0��=���~��:�1�>#5u���]�}�z��"#^TY�k���l :��$MC��W^��wݑ�Ec_x�"͟	%��ẅ́�fR�9n�"��V�m�	�{�p6�3�XH&���8p�ՙ�9g>��˝������]��;�������> 
��d��U��T�F���_q����C�-�~W���Bʵ��ό���Θ9.���+G�VW�0Ǐ�B�8r�ط�����g�}��D*`LC��^�&��{P[�����t��F������R#=uV:���w�؅�,��gM���hac��}>���W����Н��z�2Q��`�Xk�ԩ���k��U{�*��xEg��g1"Z���Zg��G޼�G�k�;�]���4��SP�RGiԞ�}�(��kb�E�iE6t�g=�Q_���<�����Μ�mW;�Һa[;QƉ�q�f��[�Gg:F��
�G��F��6��c�T��U�*�ꎞ��C��i�ȥ%�:b�7�tMO@ߢ=�D{W.I���*��T>?G�B��x�?,�]ν9��=h�:��8G�0b~`��y��Zo�����Bо�8��4�U�(�E�>O��'��&�0ya|�������¬�����1_�N��8�4����U.�WL��xQ��/������4ir��EJb��/���Z�2K��7���[�g�Y�x�?2=1��x@ԩӯ<�:��x=����Z�<Y�c4,�$xѳT���o�XӚ����}�"滵DQ$/ �x㏮���{ހQG���yi�,�)Q��Ɍ0D+ϵz��`:�,Ol���w\��%��$��!��D�"�Fu)��DD{�{��Q�G�2SHeS�{�6~�t��F��3@:A�@r��5u0K�w��*\�+q��ǘ�w���,�DY慝5�K����Vr���3"�Vl�6_�z��D�^��K�ݹҮ�t� �.+��t��H���Ž�L�=���&���z��O�/��-�\;p��Ծ�0pXN��N��Mx�/������_!��2�?a�Y������\��޼�#�LC�|n!L�������ThHE�y��4�mŸ���;0�Z�7F����0����a��Z4���gV��j��$��;9]p����u�"ȝ���́ %���Y��ZQ�P{Q��DG�2���S�}�j��i�	�+�a�b	&ߪߟV����3�Qּ<�����a�y�F��N��|�eݺ!2��/�����f�<@����lm���
�(�b��Y�[hQ6�b��VdެQU��;=b�Ё���<h�"-���,ܿ�]Am�q��vn���#"�֙��1�X�p�_�j�u���x���MZ���a�Y��76zi~��!Dp���l����k�6F5���8rf�Q�k��g���l�R��t����~���<�x�'��>?aw32��51��_ʘ����}�=HĖƞ��C�[���F�#���.�r��EA�74�α�֭�It*`e�����90v�f����K��B��Rt�k3��*���u���8���s�-κPg[E�u������R���}&]�m�DޜB)�����i�ʝ7v]�Yz�4�M
=�T���|s�S�}�N���t'^ʹ��`��\�${����������[f0"c�L�������7Q�{�[N�b~�r�*rMҮ\Y5&)shs$�9[Cb��I��ͺ��yp�b�Ս�P�=aER�l�f<��˸.v kL���}j���U�9��uyq^�L��u]�	��X�5qW�/f�q�ע�h���4����Re�'w�n��`m$�f����,��;�]b�X�i��@���~J�b�.X��e��	�m��{G�8�]1e�*��vƋ,���4�.���a��ah�33cP���g
�n�\��h�Y�^U%R:N�^q(E�)��4�+��[�[������[�N�3��k5��mH�MQd���OFjz�FVc�th��!��T�7��� �I$��E��UE���ER�~�m-jl�Z���Y
�kݕ(�Lk����J0�-��":aGaR�*1��b�e��E�TX
V��Xrʢ�e�(��R-AH��aF(%b�0Ĩ
�X�E�UDDV,+R
VJ�e��*۽���O\���� ��i#7iE�t.��*
�W�_���}�כ�p����v�?��q^6|t�F���ROnm���vyل<B�����=����K��|*v��bl`Q�&5�Dxא�l�e<���A����Y�����|t��BL�u�2�"�
����l�	�kk��	�����~�cг��zt�Y� �����w�p���]墈�@����Y��cia�K:��Ω=��,�A�;�Y������+�ޗ�Y���1�م��aD��&*?m6,߭�-���Dh�x��"���g5�ì��.�0*��?x��0�1�I{����g.ͩ	�H&�x�:f��㋻G#|�T��v���wvN.]��Rvm��/��^��@��qI�U�j޸�I;���9��%���>J�r��?;1��m�7�3�C�؆����+9�%�ھ��%�{����UוW��PD�I�=3#ˁ�[�����;|��iZ�,ġ�/�Vt��K�p$�a�_�:���p�?&����Wy�^��p8l�?@�j����!�F� �{3o&N���e��CA��]{��q4��
8D�<�<sr�	C��x�t��H�eA�S��Wha�>�(C�b�XsPI��*y�Z̭閇h@C��E����acь��/#x.n��6�kôc6�@]פ��p����W� �f��:�����Y�8�?�2��c�YG5M�<�.�Nx���E��eF]F���K����\��x��������e���Ka��@��g{|������Ś�|�����S���fj�&�WOC�깇.`�\1PO��������Y�V��=�^?Y��E|E����f`���S��M��)&�w%ZI��>(�����w������o���X�������tr�'�:C.�dJ��cF��e�u�7]1n�WD�:G4$_b�����s��:;0yaӤ�W1�9�6�#��x"��7c��惺�^nVoI�B��8�)a묮O�2N�-Q��d� ��d��=|/B�M���w�> 
��8�E"͑����a.����0�d[��+��#����g�x��!�a{?q��c��9���!ڜ�?C��]i��U����=�X�����$H���R�F��?p�ޥ{�}�����~� �Ǝ�4<�	a�a�e(3��K8���>�j\h� *k�w��,��j�$HdQ�b����Bj���@YHSxO�=��x�x���fR�Pn�#�_+
�
u׻��3�G�چ6[�N�KM�����1x��VC�:3͆h��:�C]�٬㽣���"�CX���կ&h�J�����f�N��l�7J��o����:�䋟Th���z=5��G2�Ͼ��r6L�
�ɹ�vz���!�T��W&�o��G���(�!{]6�֖�B+^g;8J�v���*1��1��3-x鳞����\�/��4P�0���醁�t���=�M1���a��"l��|/��O$疔7û�z{4Y�צg04����ï�C�/%��O^�=��g1�E����d|l�L��G;}��-v/s��d`C`�?o�Vu�:_���V�Q��H���j��5�=�NU�^z�z^�ʈ�0,���-A�X�}ti����=���i���5�mi���d��l٫<��I��Ʈo!��ﳭ�&>�af��2v.��I���,�f&_$�L����V�/-c��������@Lp�z�^l�z����x�jw�?]{�2�D�-�&H�쪵E;��O6�z�<A�ƌ� ����G�D*����;����G"�c6Y��8Q&���F�9�"03��!���iE���@��#��<^G^����˫`��!��,r�]�5>��T�y���5�+-������Z�ú�+}3�g�a5�*��C��>�%�.;5�,yq������I�\E�C�y��q��iE:yN�ߺw{/����e�,�"��,j��% ��e�G�����Dv,�[Ar�C��<D�H����W������sВF�B�#B�L}���l^�z��~�� x�����ҿS�C��}�f�pk����(�3�Q�c�T���Z�	^�N$��7���l�ѫ�����!^^ ��LPEErV�Ӥ$�\�7үw�r�:a��}��N�](�2��X^R"�˩{|��0�<�c�R���.���ɕ�����af�#���{gW]dvkB�21;�����:l�@�C�WU�����a�)a��������Ԩ�B���ܼ���n}���u��j!OG�������s�_h�f��Aha�H�ՙ��<O��Qr�^�#��u����ː��\)ёu`�*\����n�n�t��6�:�B�;�;����RϢ=聥��W�V��\���u画dȇQ�n2��;�B^3
SW�s0�@��Ez�uz��4Am���B�s�Qcɍ���^"j��Ǚ��^����C&���9"(���7�Cm���y5}�ZD0E_?�D���CR�A�c��Ȩ�_pV��ǟR�[s��53S
b�(N=�`SZx=>��a��lL<Y�0���hW�wK-����
�����C��� ��dx�#�Xb�U!�a�5��[#Oa,#�X�e_7	����0�!X��;��+ٔlZ$�����'At����� ���Bc������C��nM��
Wv7�R��']]A��ޏ{�*\}�3
c�dq}^�/����w맰���p�+c�j����P�sWD�f�	�u����^�쟞R����3���:J�(d}=+{�|2�v�ٲ7T9�6Cʏړ6t�Y7_�F�Y�#�}k���_c%څ�ZXj�Ý�$�k��͐��2E���7�n�F�w������U\X70��;A8q���i����My��ٸY��8�g��Y�'����JHe�u]w�邰�?4���������a�,$�.�l����YJ��9 �s���yB�����ېb��F�P��f�em#& ��������rNcħY�{�n�԰��y�X{^�n���~���_q[�1�3u�⨢0�'��d|m��~�`�v� �H<��sWݑ�"�2/�$�yf����"�Ú-����zp�/WR�g�@�Z��$��<>:lj��8`�*�y���U����h#`�g��G��C)�ݞ�a�U���5,����/���U���d�/�3+��}g�����f5Q���D��Q�enu��ĮbDtS�jP�[�3��B#Y���g��?7�\�[/��-63)x�^��_�����b��+/�a�����+���G��ֳʬk�kz�����;1�.Y*�
�z�oZ�*Ag ��uy���O�צ����}L�P+k�Lp�
��ç2���y��bf*��\3fk����T����p��Ү5��K�y(�N����x�^�w.oȞ��/V��|�B��2�Cz��Zj�ED.5Աz�>�3b!^X���ozE���/�f����u���=�lG��ni렷�k\��KR�{t{N厩:��ᅐ��{lc���u�q�[Ʊ�y1pP�o��V/��_,�r�J��%�FC{s�Čb5w�o�γ�y�f������~��������E����k3�li��o>��֍ӷ��kg�L�}&<��JͮBҞGAV͵ٍrq܈��P�����
��V��{ϙC�*��]���*�3�I,�p�:l��p���;���o';����W׫R�M��=1Ăt���vLJ��Y�S�m=�5��\M+,ݹ�'u�y}|Fy�Bٳ�-a�o��}�V�o�>�ES���t�J9>���R��kuo�XDjS�&W��(G���JgF%����y3M̶p��Y;�!n�̝����};Nh�ѣ�uʏi���t\����;]ozy޼�|�C�J�Ab�����*�H�E��b�j���
�dU��ī"���˔�Q���E"��#"��EU"�V�Ec"�,�P������J��ɖ�VTX
J�H�U�b�"�,U�"�E���T��*�VM4dQEXi�P^��:�o\5;siQ�g�)��S�	zz4I˾�F~��ze$���^VH���ƫ�s>9beOu:�����nz�;��Y�{6A��E��H�!Fe+&�=0�ʡ�&��g�����C���_#�j��%/���e�I����-:���܅#�Ƅ
(�E�{s�>���!����q6��k|�W����o�7̏���l�9�HG��g�O_�X}�]]���G�A!V��=9_y�WE��':0��Z�DC�����ݘ_��<F�M�:��A#�(���/�B��z�Uy�~ y)hcp�\Fg��6I_o[��HMz(��P{����2I�i��	���l�F� ���u���:w~�ބ�B�/�x]��zd|w���_WC)���v���ߖ�ԅ�����}_^�5-�^�iv��E�Z�耣e�b�b�gᒝB��i��$I��/**WW���lh�U�}����b�E�N�Y�n��Z��˃u����aܒGo=��j7jVfg&2rL����d˘�%w��H��U�?]^6���m]:��˪ćZ}��� 8�V�C��Ϛ�1��>b+��!�ݾ]�-�@�3>��BzT��u����w������o��t�l�<Gb�,��S�r��=��'6W�:���~��>~a{?q��w��v�ws{hwgA��`h<�W��y8����s#�G����t��OWp62V�H~z=K�Q7?x�����2&2����0��TPSڗ�l6��Y!���>$�.�6��FZ�<|_+�Ҟ��!��U�z,:F�`Ər��8B�n����'��,�!�]u���;_^�����E�gM�0�/���!������!7\�m ��o��k��1�F��j��U�k���UM�f
7�N��w�)ٿ�[���;g�h���1w��8xr�f�n�3�����Z�����cb~�����Fk�T|t�]����F+.������5~a��]�0�|]��w�B�u��J״FB��쵷OL0�)i�9������>3����l=�9ڑ��<!whC��G�r\��D��}9&~��>5n�ӂ������xp�V&@��0��}�����g��Ӧ߲�]b*���!�>8x����EB��E�oo�E�#���(w8a��+��Vvz��FƼ�?t�:XJ��T_���Uuxd����/��� 1kڦ�oy��"���
WQ��eψ2��v�"��cX|F�({X�v��v�����gǍ�a� �馁��*:n��]ogy��!��*(�$�<lʲ3N����7Tt��,�f�L",��3f����u�+kT�ޢD��}�UlC�j�%����3y�v�����g=S�)���
V
%(���z -D�|��GƜ���ǎ�g[�I#�}��-�|'���gN���=��Ɓ�
)��V�d:�g>H_�[�}�D0���<r���Րe/�7r6���Q���f�W���OL��E��0Ѻa�){��Ȍ����g�5�%����[-9��,K��Xgix�U�D#|�� �c Z~v�@�w�ۓ�x�6|���rE9^��q�Z��=%ݸ3�B�VC��ƭ;��qx������i�	f�;#5
�|_̌�c��4�R�!�����ʈZ�:t�Z�6x�&�a���ɉع�b���6`����ja*Fe#رa�rQ������n^���W��jT]���u�W4a(;vi+��{�s�X���ίd��d���5Q\������f�{����5HNU�A��s�$J�p2{7�U�05�9MTt�Zg��A#�<�<D�����6� jP��8Fب����̭��{2����9K��c[�����q��K:N�u�$����
6n��CY];0"|"B��.�@#�)��Wnc �/�de���O��^U�E�x`"͜?O bh��Y����[ެ�L�C�C9i'ŘX8a�B��Y/�U����c	�u^ٸ�['������]����}u���{Ry0r{c��P���e�᳤��h��i�oF��Ru�c��M+��3�O��Wnb�{��_SM(@�6��B�y1�H���B��q�g�x�#���'�K��	���i]4��������$�8E�F�=�Y�)�'�aȷ�=��L�&���-6a��gk��"m���"���?z������ő[}��w�3}�f����}�P��K��B^��-x�#[�K��YyDx�G��PȰ�!�0�h��K�'tz�T/�m!��b�E+�Rbh����8Q�v�z���w�cc�#Ě<Y���_f-6C�Hy<�o�#����!X�v/���r��`Iu�v�"�fM�io�V���^,y}%�c���J��t��49
���bwzDwy�ݖ��}UD��9u��X��Y�/������P�����z����}�G�E��j�f�����6��O=��cH�n�7+�xS��,��}}Y	��pa�g{7�U��x�B"͟���X����w�s6��Ts��Nz&:l�?C��cM�6u����_d��ţ�?y/��A"r�<��-����٠�y!T�yad6��Z�.�`��B��"�����=�:t��ZYR��j� ��\_s6�C�X�@��F���]���4�Mx�F�۾�W{�]�<FrP{o��]� �	̫�3�	I����s%�G�Q<-a�mL`�eE� �ow���*�9��+���י����H�T��b���M��7�����,�$E���5�H�[$��w�|��Y��f}v��<D:a�R0ك�zt�:g'(��Amlk���k�Y�<� ����e�����W��z��.��%�r��Y���hn�;�m���x�B�I͙��u��zeV��Qq�iE�1O��"�Cx������4,���Y�_l�/W�5'j;[r���3��~��9P�!�	�b����\��ֵ댘�7��P6�Q��:���f�#M���!ba���}�ŝ$���~�la�(�V��h����y*�.�Z����e�)�/��Rc!���G�Co-;�f�9��R�/����=�&˱�.�~�����������h��5���1�#gO�j��,�-w�5�
��U��`,rө	�9	��<D��uޫ߸CŐK3i��:'�Tq�p�MGS��[�	)<��S^#`��9�ϱ1q�N:q~��^P�o��*�Bj�ex� �\�|�]��5��Y掑���Ax�$�G�yv���w4�Ԭ�4�U�2�Fjʊ8a�G�̮��>�GV��XF<Ӵ1�p����B�=�Ý~,#q4���?�=pQ�ݩ��GzƇO\��MY�;�.\r (�Lq~��џlgkI$j�vDfvȓ���Ykj0&�M�BێF��a�U5G���7�TZ]�O�T���'6DJ^�+D珯:6���������B�u\#�nMy�r�ѓ@��ټ`��ٜ�;���a��W��R�mۮ��d0��3�*tiT�6��m�bf�6��F�Kq�"ͩ�Ʉ�T�s��;�uh�U�sqbVL]�\rr͒W��-m5�{�NJr�4(�B��(����<ќ:��E���%�K�Bj���N��5�CYXK��y7]1T�����ܒ������K���n��$�؍I�+4����:V�(#�(�J`�x�P*��/` 
�������VL��C�u;���躁�g&Z뮧�d<���3a�l��1F7g�٥_��o����0�&�OHi��5��)W���5!����]�x�ʜ�b5�i���M��X����W�;h��*���i��sG|ۧQm>��.�.��J��oF�Z�P{@�T�ȗbV!�f�鹼�]&����]�VN�+tQVp�������U��N�)�\갗��q�}ۗ	1��.=ʮ���+��C	��w�:s��R�^?�+��NPܵ�#DP<�I gw%MW_T��պ#��|Yo��\�jV�:���Fe�;}�ŵ�Xw���I^�����t�	�۲��$��h�]C9�n�ыꬱCJŶ�
���H�F
#VE�m�*��(()�E��X��
�n�̣,F�V"I(����+!Y"&5 �Fc+
�+��bd�
ԅde��t�CAzb���1��T�+�@����!�����8p�{�^�5�9���ۭ�;V�;�5UH���̌7�P"�#�F��u�lc����}�qۣl��H-0��}uL����o�.�Gڼ^!���n!ܬ���TX[_jB�V�o�N@��ن��H0�'��ڱ&a��2&:OMk��P�Z��sa}���3����h+ީ���"���/;6t�- ���r�:��[��t0��H�>VE��k��>#�OY��,���I�8Ʒ�\l� ��ȇ��gG��wn:$CDsV_sr�G��@�L C�i�*R�M�µgH�@^"w��DA�����k��
:}4YC�8�/1�:.�}z��n�8�(���;1�N\��q��w-��.)v̕'?��ir��mVu��-X����`L�dx�v�9��H��ϒ�? ����^�~b��M{s�����Ig�HBȄ��Q�3��OI\,��?YO2�����g�E�k���d{"�;=��?T��_��i�YJ���Yda�L�n?G�޽ߦf��>#ǈ����,#K;��a[��^<~i6г5��+�����`��-��^<�?9i|�8E�hn+8E�`�����=��x{ct�1x��1�DYEt�C7��ɇ;z���MJS��A����,�HNV|��Y�aN���j�1o"��72F�B���qo;O�/�Cܥ��.HsVo3�G�ӹRw�������2P�E�3,�&IɆ�tf�c�[;ҦZ}��޹c�Q]�ϗ_�}c�em.� )z�*aj]�/h�0TS4�7�Yqv�7Jh��\���t�y8�%���;��:^yJ�^��J<����l�2��חR�(U@��3o'��Q�x��pK��dgV!
��6zcYpjx+Tܱ4"C~�;n�wl8�]M�-�@�{}F�@}[:�f�.�}C�>�94]Exg�u��p�n����3���OqjG3�@�}4R�g�\��^���T�=�XU���+�꧜�����<?F��5����%����"�S�y�Ne�۵�b��ArՋm������7f���:P�����
�{T�%�y<T�-���1��gvH��(��Kb��o����j�o�n�T8W�����}$1�bַ�w*T���;Y]Y�����Ly^[�\��Y��|oY.�,Wo!�^�4��f��Ix�Q5/!�Wz�2����p�p�}t{A�;�m�v;�ᜅA¶'T
쟷�sX�<~ˢ�2G�5�i��B�V�O���E�Է�i�bb��X�{k�Io�p�EV�n�j\+�.aT��M-ڸ���ֽT^Nv�D��!Z��,�C����1�ų��R1��:�`�a�W��X駓�p��{�sj
��޽�[`�pt�}�/�P�{Q��� r������ Ƌ��ܾذ�N��S�n�لm��n^���M<O'�ʛΜ�m E��3(�-�ш{F�jL����P��XiwFd���k��v	,5� �=�I}#�ꣀ��y�"�]ˆ����u����|��OZ���٨|�n.nV��Lb�ۃ����o�^{	u��or�i��4`F��}�L�+ee����;KDYṺj�F`�W2@����PzvK�s�^�Ί[ѧm���VMnWf�6Wbcї��S8�Õr�[�9;���>��|Q��Iy#zk��x�5��T#y~#y�{���:�;]H�{y�뷸k�w�\�9��a����h�죖5k��*��G��,�����4at�?Q���z�~:	}D×v:����n'�GW@z4��X7�'MU��8�=�����oy��9�k8g��;{͇�wɨ�f-��U�F�:�#�6��[�+q�y�w�b�*���r���b\��a,���bR<H�3ZKۈ�E�Ey+6��y�/��y�`�}9��<�:�[����D�3�U�[�l.S��>�rC<GNC�>�"�����vFڮ�$
>ˣʯc�.���\�,a�#>� ]�l�)r���	�Yz��^��u�EѨX�=s��K���wkX���M�E�����bK���xw�ON�Ӭ��j�U������Q����n�#�{LV�����3G_���{C���f�5��|��W��fa7�ta>sO��7�n^#���k�~��v��wn�Z�w����զ��A�o����eA&��B%t�ݠ�woj�܇tAB�0��w^�9}h��"
-rd����A?.ߝp��xH7F��K�W��j���"�c� k9h�0��C^Y>�S�ۮ��%
P��}=��N�2��=�Pc���I�}�J�yӢh��UJiC�Y�{e��è��0f;R���ۛ5�1�3��h6�'	ŋ�5Z��^������1o�/W$�v���[v���.����X�%�BзM���F�)�R^d��.S|�.˻�#�|I��mbd'��*i{%�n��:�t9�:�>��	��,ú��i���j>�߾�R7�?��ɕqƫ�ӯQS��X��Oe�x�e��+�]lɄ#�<�똿�z���F��f��+���Tr����d<��'���H��/'��W7��g����D��������=P�\�w��4�0��˩�.�,����Y����{��6\b+�PU���p�O�*�؍]i�Rx��u�ժ5����팳^��o/�0�K���qj��8Nt����-W�p���U�$�֑�R��u��Efw-U�ɂ���,Q2nf
To��<��{�h�Fn2��[	��/��%S 0;hһ�8�7j���F��ȻN-�x��`>Tӷ�P�p�ӌb�(��7x*���n�5NקcX�P[�ݔ�ˋzf���p��7zk	�Q�(�rF5��)���l|eu��aX�!��5(ޮ��)[���M�CE���f���f
��9�۾wkDB(�iP32�6����6#���&Ѻ�t˨Q�b�6t+�)�i���7qҭ��*���2�Q"q+�� mѤ!���cj��m��E�TU���qӳaeb&�<�-U�uQ�A�JAȝ�9PR�-]:m�/����P��t�e��K�G�VZl������ŋX)!�+E!v�c�1�vȂәk��BU����1P�ᒤ
ɩ�%P,���*⴦1��r:�I���9�pb���&S�̈�4c�aB�Ճ�\�mЪ*�UD���B��N*P�q���F[Q���3#r]�+ʺ�ݙDƚN�a��(V+.*QRcD$��I4R���wP����mX���U��}�{�E�Y;��J�T��Y�Ӥ��*\���*�Xc���B�Y4�*�b�I�2�X"Mj��V��%�)4��j
V� ��J�up�,�]aTu[F�Vd�Z���I�uK�Kh���a�m+Y-�&25�X��������V��RI��I���{��Ywՙ4Po��@]�)���鵽!wr�Fh(��2E�몴�=�.T9�j��-�h����:F�U�G��X�AVm��|hz��<x���kg�lA�ݺV���9��������Jӽ�r!��x��	�5;�Wc��n�v�uV��0�Ҍ�<�<^��=�YZ{4n؊��m�Q:��:j�a �(��8��YךT�I�qx�8X���+��������2�`��P�R5�S��+QN«�J	��^7&�ΐ<7���E's�9ÄN�����~� ���u��'C�/T��C�]��GOWf1�j뎃
�ݚyȾ���S�P�P$!sr�{�U�]�Vp�@�l��$v'��x������1"8٠�aW;�����s�:1U9��9��U���b(��x�!w�E<[u&.�89�>޽b�~6�:�\��L���S�$��x�4^)u{���߅�j#i��rs\"�ԧ+�H"�oH��t�we�(䣊We_P#�1E�P
��I�}�q3?U%��v?ߔz�d����m��%�j�>�)rq����=7 ���k�՟g�^A��5:��szS���Wұ�2díꭵo��>�e���L6aaJ�$���Z�Uyen��B��r�NY��p�v5gv������[ѝGp@=�b�)^����]{j&�`�H����䂓���Nɡ��8u�������9��j��.�Lq�"F�(��R�ŵl�ع��nh�8#&w8k9�:���wJP�}]Ԧd,}�-1�W\#�pM�*�)�Ì~���NW����^[
�1�L�'ңw0�f�6�����]������];��q�e�[ՠ�wl[��Bx0Vfj����o@Q�����Y�W��3�T�nF[
�R�'�5����w+nt)���(���f�
��s�),���P���MA!���2CY��۸e��b�Ěa�ރ�eΩ�-E��9>��wn_Z*��ţ��ű�x�����S���Q0~�t��[�ʉi(��sE��-�e_=޹^ǔ�f&�Z����E����Ȕ����\oH9���5Wfo^=�>��(:n>���àw�.�)-�᷷��c�ќ�L;�4��B#f*�vU��Z-3��WFN���|��� ��b��ŋ�c6���.1�=�3�b|��	�z_�7Y̻�|�zTo`�5AX՘{�ư��+*���cq�F�QB�3۴�C*�^fN7l�}aE˿����?*�D(��M��^k�wf��r�
�ަ�ԕ�c%]��@<����Z i�Y)y�v���F�ͩ�3�O*�Py
s@o��bה<sz���G���L���>K<���/h�t9Z�:������|k��+#!�P�O��[�\�bԙ�-���[Н�kC�ă��J�*�(B�=��b�TM����T�T��h��\�}��i�����2���z�vn�]׶�>L�(%(,P^x�GO�îx��i8]ӇVn�1[�w���{��Ƃ�,�&�>�|o���������P�(wwJ�B]�9���s��g�B�ꞑ�=�G!UhwIW���Ċ8�����9���
��oJ���7�Nܠ�GM�bV)[̙�A���zJ��X��A����oC�P�pr�y��y��3�����ƍ���h����du�>��[6�VU�[ܨ H8!ASH ���6&�.�ԱQ�t]��f.�ǡ���:زe�����a�;��Kx���\�h� U��q?^��)��33^͸A7�ٜ�>����������s��P�ᙐ�f��$4��[V�d��}�^�=����B<(�j m�6�uU�������um�h�+)��a=D;;���c#�V�/	��缝��n�*��c/��.�lh�=~���r�תeogM=�׺��d�n�F-���s;��{�ɜ�N�/�B��y9���ؓk�쥅a����G��Z�w��S���CpM����v1Y7h�=k��n�Я��Me�n���)mGۃ�p�\`�����J0ן���O#�$BA��=oo�^�Y�6؂i9Zx�y;d�ܨx�kDh�e���ѻ)(,�sP���X�AC��Z�X����V��w��&�9���(-L���MC�|Q\�[��&���X��U��tS��^��g0*X/�-�;�gNؾ��7%I��g�M �b�г{34�۞�_Z���ٲ�3�J��4��qM�s:��MB��=cz���2��z]Y�R����}̴r�s
�@�wF7haH|���d�}O��]cЩ�\��A\����Zo����|�3ya�L�D�$<���ݪo����}�S�˘g�b���׺}�ן��c��><K7�@H����w��=:��������U��F��{���w�kx)5$�=�бW�z�:vN@�z���5��!������Z^��Ţ�ӽ��!}�U�%���(��ĺ�nɏbx�v�c�*��N���H�9�fj����H�/sЪ��9�� q6�]�޻��h��V�HX�s��6�K5ovE���^��1"��*�Pv�o)��N�$j��ە�Cn:���w�ű\w�g` ��ֶT�F���)�d$��Dq���fV��C��T��{�Do�յ����O�����A�f���z�S���c:,�i�w2��ҫEdM���,"��rR
Ҵ.�6��;�y�I3O0U��i��l����I��b����;u%&Gk�V�B<�㧅BLM庴�
�FZ��k�n���F���t�X6m�X�[���j�b�.%e�M�!��&R.�T�Å�~Rˊ�v	mQ���S�p�#�# ̢�7�YВ�D�O+*�PЁTSnc�fe��(L�\��a��s+ǘͦr��׆��wB/����[h���ef��r
 �����xj}�䣅���˿�aѴˡ��m��Cp"��laX�*��������E65 �T�Z���ԨJԾҠ��e��ˎ8��im�P�-+m%C�m ,(�,�3Y1b����-&8"�mJ���XU`�ԩZ�
ȚK`�4Je�ӋE�Ec*��H�AT��aYKm�Ъ���Tq̮5�l��K5�QF1f%VU-��V��Lj�U����-��%*ج��sn��A��䮃[�l�(�Y��W���ڏbէ{��*����چ�638ikG��p�نn;9��6K�V�L��Y�lvܠ��}p��a�s�v���zק���;s��~������ʇ�GN���yEL�e�>�'��31�w�X�g�s+&\_K۞
�����eT����*t��uZ#6˙��V�X<�/�|�A�B�օݪ�1�r{/9N���B�vfv��.yQE��6=R�dxWg���[�@�U�j�xf;Fʗ�\�6nޜ�d��2d6��v��赘 B��j��B�]�FZ|VU��*o�s��J����/X̮��$���Stb�fX���h���k�'n6ZW;�ld�gf�]��{K {����D��Eb���GD�b��ԏ,B꣧;��GX�卜�z���>�lR����ل8�z�^M��s�j���#�̉�|��Z��>pmޡW�.|o��u^�G�Ӗ6�Td%����y�.4�
��R�uYξ��W��GA���@5M��:��M���5�W@� �ॡ���7h*7l�o\�n9�S�{��en��LI���W��1�ua�bX>T�����H;zMt�E���ׅTi2�}���ts��oS�����JGq\�����՛}u0_N�3����y
���z����� �eg]��0�sη�d#�ܮ�!ܾ2�gh�II��|�"�Jr��f]��-��ߙ�Ǳ�2�S7a�p�����T�Z~�H M�	�w4�@q*V��wAӹ���c�Nd�m#$���� �x���HF�n�.�q�=�%��U�Ȏ*܍`RvF���w+Zr�����˃��{3�ѯD�f� �%��Iua��i�)��v��	��k���Oχ��|�y|j˧%`���m�A*��3�۽]�s�b�����d��p��b~��ܺ=�mz�k��6�;kG���8¸5 ��G���{$z��M�L�N�"^}�,��v�^t�f�=S����R+�y r�H�rW��7�x�����-�Vٛc��=闦�4<����\>��{�ܴL+M.��_��}�X�hj�t���^q^	��k�����@$`�lG�׼��;@�Z�o1ל�����h��kb|,k'��Z��]�r��3q�:�P刽YmW�[U��3"9��O4w$�)P�5>���*�}kC�"�7AߚK)�Kr��Ɣ�Ai�}�7lh��݃(���wR�j���7��Ò����4z����\�u��:�>}Q&�I�T(�h�՞��PC�r����������yl���w(��Qm�7j9.dnvze"��7ɫ_�O2��mz��A��<������`��yKPS1�� �զ�ЮD)����f��8>���p޺0�8�J���Wy�l�2-9�~���k�=�\�F?'ۺ�4R�0�܂WA���Պ>Ə�1�ݕ��_e�бY	kWr�ZAU�'VL�������ύ)ۈ���5>�V+Mf�on�A~Y���F��W������.��Ei�솙�ag9;��z�e�^��L�p.9λ3��6�b|�ky��wX�ź�)�^u�d��������M/s�nyn��=���{�g�m��K��E�䒽�s纫Mb���S}ֳ���5��p�v�~սv�DW��<��N�s��a֟}�|C���}6�e��[^���/�v<�8̜�p6/8���x[����w&�Ѩ�Xy-\�iH�^�w��b�U`=@���_לY[/�۬��w�<KJ<�2<�$���x,�{l��e�V�蟝:^c�)c�d�yy��n����}�<jM�l�h�D4�G]ոG{�bN�{qؑ�����V3�'��xNv�7�	�\p=���$ʻ@&o��<Xr�����)�=�Ǥ����u2o��[�p;Um���!�;���/��s�����\p�\�;q"���sZ�q:�` ��I.
���!#9<�r�`��*�H��;4����Ts��)�j�����.����5n#��݋��Al+y�퓢�K={{!�ט�e����J }�ߓ�����<������Opl+W	h���[�/c-�P�L��+i��+a���˔}���z��V��V$(�B�mn�6c��뮸�'��OWD���>��2k��*ݮ\ҭa
)a��;�;�t!�#��*SQwf��ڍ�m���Փfc�
š�q��m��䫕�*�c�n��7.'Q�ͥ������M;!�g�[�R��bwNc#�ya�Lr��o��E\���:��1p~��<��QK)��6ǲE^��N��7�8��Ѕ��fY{�{5[��pE�aQ�4��@�N�p��i�I���ӫ'�/�k!>]o�^nB������xċҢ��|}�h/]z\�>�-Y���\:^�����f��/"��rZ�bv���)���&�)�t�mgY�2YF=��8m��鎜r�6�q�{ӱXo#n�bӵ�T�Ko�Z�֙1�%�ikbC-v�
�L�-{����]�d�9o%�d�Y|d\ī��4��A�֤�|2�VLT�;��X�-�?�ʼۼ*6Zoo�����}b��	�x�-�z���WK�h֌��m�i��nN�U�G!Fh�Yݹ6e ��#��Nd89^��:��d8_}ܲ��]�����\��h�� ���j�!�l�d�f��,��x!W!�u�a[c�z@)��pn&�إn�Y@ѻ�Z��I"�s����	N�5�jH�j	�`&����Z�1�IUor/�Ĭ�4��U"��-�%�³@�#Y��yL�"��h�n�Ԗ�ßX.��$Z�ofZ�E�� �1'PfQ���^+��2�ݳH�#��s�Ln��h��ZmRĳTv�4��(�8q�aT2��.�w+1�j�17�;�];@�|�]a)uV�ɏW(��Qyl7&��oJwyL'H���zY�i���=k�f�F�Y(�z�j��U+U-*�X���jZխE"
���1QQZ�U ��R�2ⰣX�Qb�P�EPG�b��D\�U�Q�kF"T�UP֩�&�E�TTR�,uJ"��b��X�)V ��R���[jf`� [X�R0b������8�.���(���d]-�ZYZ(�+�����Ѷ��B�������(�B���<�-��^�)oC7Was8��o����}�uq���\�~�d^Wyc.������6����S��\U �v����w긩v��	��3�%�a�:����Y1��sm��6�㽉�ȼYiB"p�8�f����xú��j�)��ݛ|j���hP���J����ɋ���Wv���[��'Wl�Ff��L�ͩ4��u���g��}6e��O�OWe��0-�����oph���Y��8KjЄ��<�옭ɐ��wb�}dunI�u�˷ء����Z� fp�B�g6&r�`�(������k&ے�Տ�YN�o�b�䗧�I�ۆ5��j�O}���A,s	-\��1O^�����������n�\�=�X#��O���)���9��C�C\�f8�U�绗�'ڹ��ʔ�ra�At��Z�gSfW�O6�orDbvlϭU�M5���^nn�
�gb��!N[Z�kI�E���w�����nP��Y܄);���x��Cp�rB৸���o{F���q�;^�h����b���Z�f,�7��9� Rp�
���� 7q�jB$�.�I��쭾�סz<x�g��9Y$�l�T� ���Ik�[���]^S��Qh���>J.��	Y0�F{>��*scU�^�f�p�B"�$��6�'����r����ς�(���v�S 6���.Y[7��t��RĨ�0�KGj�N=[e�`�ۢ���kYH]�}�M���{=�Wj�/C��C�G���#�Gi:B�E!`-��^�Ŷxċ��,w���à�r{����?{��C�y[b����e�y�u���8�Fè�M���W��\�F�ݿ'zk�;�|,��Vr1���!�����%Z��U�^�|7�y�\��{�]�ʇ��G%B��^`�[w��\ȶ�kk���'6I�y#��^y���pm
��n׃��;����آ&��L�����˻����.^�������m�K�usN�wk����v�M<b�$r��{	�zw�4_���E�iյ&�=%�c���/������r�o��X�r��j�n������7��3,e�{��4�ޖT6LS��fg�F��=�\�qx�{<��.�{A�ba��gD �V�w�8�,��>�UTM���W����_�)�/�g
�μh�<����|[���J�+]��ǝv,|���:O�^��^T��Cřn���[�m�As&�a��V��g'�QjSՇn���S[�<y��w=�e����tGk��1[Fh9ۚd/yQW���=K]�ء��rm��[s�}����.X�x�]3��!]H����m���n0�
th�`�<�ǈX���o��g����43�Ap�>�(��#��Ha��Ӑ�"f���Mz�T����������p�,�W�AK~j��ݿ�魓7�w0Ͻ���yH�]�f��ZG)G����.69�E9����K��I<J[�H���'���<�
���;|P�oC��PMop�Q\7����0q�Y�Y�7x�g&� �\4r�T��ٚ7�Q��ATqyQ�(ć��W�}9�w�V���[�ON�,�*��y䵑�^�+��L����_���Հ/��~Co�:�G�@��Ѹ�����Fa8]M�mn�}��<�^
/�e��x�ͣ.��.:�U;1z�'�0MK�}��wu�� �=�r�s�m���r\!�|�pє�E7o�oBU���m�q4�C�N�t�����9��k#9�U��E)n�u	��ϵ�f�n���t�pk�EL�[�u�C�'���Jy#qC@���_D�s����
����wn���f73��z�z���.���Î�z3�֗
��%19����=�[�$�n�|T׶O �ǹ�ZE�Tk�1�yҍ랠"��ɖ��>bD_����ށGH�y#"Ů˸��q1���3�M�ڞ�D1��>q)�U�W�O��o'ov�R���B�6d�Q<x��^\�*��t~=W�fWNR�R����Z�`ٌ�mu��5�����t���t�5/)���R"�DU�@��ni�J�fr��Y��6Pb���N�{p�4�T�l��;vGC��R�T^�y��hx
,����v��@yz�kϰ�!M�X��q���Ԩ�&�^�`҆)�e����''[c ��/"��N��ӻ6� �̩�*�<Ve�j�V� k��9Iu3�@wD��T����fM�����U&|�(�%��GD���ɕR窾�])�t�f��8�^=�j�w��؁sK�5Y�Z%���ss$���5v6:bf`�!��
��_�N�Dr¯uk�3�iuG+o�$K����W����x����D�Y�bHrC[^<�Dk/'6�$Ѻo�����;�Y���W�f��J��Л�s��A����.�lkX���Wz�)���"�mm##��5Z�T� e��[��y��0'|NfvI;��S�꾮t1�̐��*�gT��3Ok�����le��� ����8�d�6�+�u��vPlvD&�uqGH�286K�/b��n�à�j����vZ�Ԝ���YEBƹm��u���˫�;MΎP�n1*Q]e��G�ob���o*�-�Ҋi\�����{1�'[f�D�
��@���4�2���|&�(,S{s�%)�Zi�3ڑƝw&�*�Z�sӤ�����8pV摦c����X�wgp�AW�;VҩNp���S��n&f��saYs�]��)�k4��]�u�6�[����K�T;�M�\�,{��_3uҭ��G�7�k�k�\��<{��y0�v�G$p<���vG��5�k"�$�+6Z���*�IX��Y�%1c,f.�|��V�Hۯ��|�U�(J|��Oo,ȩ�$��J���bK@�K�u�8����yw����a���������I�G���,�Φ�����1�.voJ�AywYQr�,p�u��/ .��4_\٣��g�3:.��
�Cۅ�v\ݜ�2h�ۡ�tP�0��F�cj�Xv�t�u<J�d����`����nk#K��
<�[
r��7{o���'��-�
�
�*[dY�X"�TQ�T��'v���Z�Qüpm�X���F�UTT*U�m�B�m�J+c���(�Ulb�����V*(V����#�R*j-�e�F��-*�+Z�n�1�X1�UE��X�Z\�X��b4�G-A��Zڲ��ch�ՕZ�T)@Ub-�UR)�F8�#�U��.5��_B��J|�{��̧��m�x����U����"ᇡ��[ǯ�8�GJ�1Pؿ����Z�#+so�z׭��
>۲�کQ�h�a���u,>.{���v������e20Oh���m�V�����SV�\��`��{�M�\�.��ȋu�w��N]�U���&�]p�ų�m1n:�3U�;zQ��=��
dlC>�J7��5��T����5��\�����#��Z���{�62�% �*�^*��5�(gqX��ge��!�P/����i��<Z��]�܋��d�݋m�Aڷ�Ö�j��]N	��e��E�m�=�$�o�f�Ǵ��P[���.���	�"�2�w��S���5^��=b.�VE���i���be�uoH�C���^�O{\��O c�M�ۓܚ8�=\]#Y�ӵ�R��25�~�_� �����r�������K�-I�1���T���L�2$�:��=��ċw��c9jh����I{g#b�=)lȐ�Q</�	��S�)�ǁ1��Vu�B�_��'�⑞�G/��2l���S���^�<��*��E�9�=�=�y5Tk�U�ǃ{���2�1���3�z�Y<t����X]�����m
�!�����'ڐ����w\[��O�N%�8�(3�p%���QP�D�b�^4��%ݕ�0�r^��H��k�6(�1<���31�g��o��z�o��{o��b�o�Y�,=�b��P�6�(z�fՔ����e�S�;V�<O����lv�ռ�$O(_r��:�d溤I���nM<Rq�5��!V�˫�m���J^��{����y�f��펥��J�V^�	��%�ʫ+P,E�9��J���|Y��=B��Q��j�q��K5nZk�l=�^��0(+����PeGr�1�o#�n �8���5:6�OA����Ϸ���<�Wfy@35�u�<��r��u��%��Kŝ~�7� ���p��������7B�3�=�"1�Uɘ{
�y:���X�T�p�}hn�Vrꤲ�!Zᇉ%!{���h,v���{ԽiM��Ե��b3�Y��W����Ex��U��.ó˒&a����k�H��ř�p�j���Q��U��>�� �9W�t���\����i��汪��-G�����]u,[��(Vdl�I[��`�wv�	i�`��Fs(�.�B+�m-��b]�k��^�!��V�GN���~�tX���k�/�T<pߒ[{�7�3U�UP��v�{�� �q�\v.ە֢�w��"V�h�ط�6���q�E�0cT�O��s�1�BC&�5۲Kq���5ي�����i�c�%r=^�׏�Z�2���y	.w����زEsr��6���	�\h�� 0�r�nD܌�R�P��^0��6�E�e\�eV�Y���A|#F1uo à-@����H�����YH�;���w�W]��9e+��S��6�Q�(G.���U�P�$����2ӳ�K�cBp�T���t�]���ۮ:>̣�5�2FHޚ�V>T��H�����eA(��ڰ۸0�[�q��9X�#g�������Me���~��AcS��<E�K=rm�ܣ�ik7�*Tl�)��ߝB�1Nj���sDH�10���h&eq��}=X�J���囸�ƹ��XغA�2�U�O�Oq����ސ�����*�xNևWE�W�O6^���¹TtN�]�i3x=Z審��ڇ.]��{�b[����y�'�\�Kq�xR�8
��>Y;yn�R��t�7[�)�Bf��*��eS�z�|����3x�2���7���rw:�lk����a~۾n,��maEOUGKۼ��87�ޓ��
��������_�W\J'j\^�*�S���e���jEF���[�<�V+>:ݪ������v��^n�GX����ƫ�_����K^1�Sʨ��v�T�<�)k��IMSŷkÊ���r�����A�z;V	0�;WbP����t�=Z�Dy=}�Z�.�EoM3�p g7쾝�e^{j�*f��k�/9�Bd�Q�O��5��mly��&�Ŷ�5�`ff����f���іtJǱ��d��^Y
�k^��:�|p�.~M��$�n`�G"c}�5<G+@]��z�Q�/������H�=�Z�+ٯ~�hRk����(�q���:r�ź:�����1�D;h��9����I�����p��[95��>�GM���[`��#�CmWh��RK;E�S�uj�!��؏�os �uw9'4�!�7��zzC�����nB � �K�+���\����:7���yk�V��Z��;����Q����>�g�:�}L�j��X�1,�g<G�m��`�j�jG�n�'�,�n�䢏wl���#O	�1���#k��^�㲕���
�v��I%O�"�_[lP�on1ŧ;�Z�q��ٛ��UI�ۃ�.��������Oӥj���xZ�&4����>�.J
�9�����$�Ԗp�x�V�岧�K\��b���QQ�R@�B�sxy�G��S���^\!)u�[iDnegT��v�T{�� 0��ln��[��3�1s���.�
�C��JˍS��!��^-�F!�����p�p�APG�M^ӎZ������� ��誂?�pF!%hu��$�!�?����ڞv$�k�?���r,�h�@�:{�q���?Z<�P�@�a���h	n����K�� 6�Y#$��j@��V�3�K���9@w���cW�˰^iā��K�PT���+�'mOU.APT�銅D2b�
ea���I�iOG��yd�0����PT������sm���I��!��K�T4�@f%r4ܯ󨯋���O϶��{�M}�*ۭ�T�E�I��S�:{gօ���e�MK K�>����Ŀ7[�DY7-��/S���Mhr/���<��A�Acÿ�b���Ɏ-�hDzI���C�#�lD�x�*��2��!8�1+��\H΁��`X$2��\�� #p���0>��B6�G��t�@D`��#c�sâk��g���+R�?;���2}��BL�X�\h⨊�94��!w�A���́#cٰ�g�X�����������'�᮲Ǽ��n:W�>��8��O�jS߿Y�W����#�rw[i�7 �w��*����)�A_;��š��O3-ٟc�թ6&�p44��I{&7�'�*� (�����Ǐny���{����ƆZ�qm:�,��#��p,u8$SI�tă� ��:nS��ra�y߉`�����y�� U��6����lp�Ѡ
��@�:Sj@\+����#v�b�$!l)ʏR��B�y�y"�g��8?ػ�)�8�*