BZh91AY&SY!.��N_�pyc����߰����  a�:/:P� (		  @��U@ �                  w�yP� ���| @ r @ @v�T| У����Z5��[f���
a��Thd�"ᜤ�\1�G٨ё@$hX���D��J@I�]4� ��  b
o�+&�ɛi�B�2��Ph�ST�4�e
�4��JKF��d�^�w�jy�Q�1�[5�N��@�(fiPi�E[U��$O`Y�o@  w��+eZ�M��!��[&jV��VZ����+m���r�{���VSl6���X*��)��UZjM�R��� Ī�6�*P��E5���i!���1B�ރH!��"�=Q�"��a�D�`�2�mJh5�	��R*���ө� )#�ۤb����ol�ƘcK6��kY�"����j��q`�vԭ��ٱ[�h�`j�Kf�6ʭ�x                � � *�R�!�R�S@����LF��4S�%T�&� G��F  &F`*H��4F����54L��Q��S� IIT i�  b   ) ��)���R{I6�O5	�����UT�h��R�J0F F�� 0F�$�)��)JB}������o>+���* 
�J����=��� ��@W����Rʵ�}8D��_�l�����	���Pp�O@�f��]�UQa0�����*���D WrQ�2��	:��%B�t�B��s!�OW|��w[���ǧ��UҪ�et�j��-�ѷ<�g���"=�՞ú9�g6{g��5�WA�ڋ���l��������:��G��� k��$���Ǉ��<��,kT]b8L/��!=�4xߗ��ў6n:0.����+��/xg�Vf4���Ԩ|8�?G��<p��a��.�/�}^E�]E����.yw�痞I�mcjE���G��ưgx.V�w�k�%�0�����x���q��X��+�ǚR�<�JW:�]�R:��߰o�p�I��;P���4��P�7>I�N�ñ��r9}��֛|�v\;|w
r�	�vtx<���;��s�ԍ���Mܜo<'�S�1_i�m�7�N߆ߚYIz�Iw��Cx4�����z8nw�&߆�bi'�)S}�M��6�x�L�my&߼���o������i�Л����%bI��6�$۔�=��j�n=�H㞤ݏ��w�4�����M����4�G]��f$�3i�Ԧ�7/�Jڔ�7�I��ݺI���L��~�K�z�n���Z\�)&ܻ�ߚY��%��z�v�d�(��t4>ZOö.ˆ�M�O00�[T�<����J�c�L�ļ˱������]�1C�s�Y�琉���iW}^"��������-"L�&�>��l�<d�z6;g0�<�â�*��?�'�q�G��X�y/�8��I[l�,�b1��g�I#=�2Fy���+�KK=-+G���-����.��`��hx%�cĊ���f2�x,��GYiz#�v
��Jx�Y�}�|q|qaņ�-���ѭ�����}����ٛ��1}"������n�*:Ĩ�����:(s���|;�Yx�^b�J�B]9���-����J9�rG���������O�IGa��N÷�W�<icK��9i&�2+Vz������=[o�sȳ����Y��f��g�~Sq#Ĉ쩢i%C���ԟ�����Gg��4��1��yb����2e��L^i/ifX�k�$���H�RMɗ�y�g�ԑ��G8c,Θgq�̛��R]H;BJ�c�<�q���4�y��n�&�RY��r�Y�&iOW<��7kz�����1S�1��ˮy{����SK�K�O,��y�y�w�y��mw۵��u�U������_{���֔ά�C�LS^}A�{��v.)g�<��]�N�yNmM&B��p\q&�~%�%2��b����C��M��Yƕ4�Ği?�o�����!�17���I�R��y,M/`�ȸe�,�ٌ\2Kg��.D�)*����1�Ɩ_�0�Z0;ڪi�Rm�%��T�$ߚY�Ƒ�r�e$�wi7X�]L��q)n��y%���=i`�����$���5��)M$7�$ۡ�3��M�RM7��q��7��I7S"�p�JNYĞ9�M�y��B�>�6��o%�����,��K�:[��3Ne�դ��K�1��M���v�8��ߥ&�%�N�c~a\���jWc��p���1#����o<�c��-.q���=I�xq���I���a׾^���5j{"�d,�C��Rm�i'h�bg�I3��ü����8�I�챻ᖖa�������[
N1$���ԟÇ�&�d���z8�,m�U7<q&��`�ߒQO��C��tn8�M'�x�ē�NPg�%�v4X7��R]��]J\�
0��*�M��O�w��܊E<�i����/|���)��ݭ嬬_i_iWW|-�K��Z��+�=����WK8Cd[���\_'���=�xz��?���֦��w|x��F����Kyi���$����IЋถ9I�I��b�&�]'�	ip��=Gc�!�k�y��v���S�||}-���H�q��g6H��ԓv7#��X�ڔ�v7/��M!�JM��%�����<�bI�#:�ԛvc���v�o��7#�RCBF�<�%���S��|I<^I�$���p�m����;�
bM���I��i7v��[IWi�I�m�bN�)��I&�)6߅��!���K�_q�+B.�6��6��;L��C��L�aޏ�Yfe3��9K��\I�V�w�`���D��Χ�$]r��9���H�U)
��ıߒ�Ѷ9b��x���3��G�)�h�&Wj�g�Uxe�2��A�a^�-ɇ�yfȞyo���Y�Y�X�د����G��U��t`�.�zF��ݥ�p�J�`���\L��|JNJ��
����;lL�8�^)����:���\c�qpO��I������ğjlL�(�C�;=y�ql�_O��<g���1WWI>�BT�\u�"_�U痽9��9�.������3˭yo]T/�_k�o�3��Y�<���{�����n�ѕj��0}�(wԭ�
G��/�HU8:�x�����l�pސC-="�>ի�I�;i6�'�V��劐�H�~:?�>�9ixi[I[Je4�����7�K�I����J���c�J��G��$�vM��K�+�H�q.;3e�����>v2����X�*�Ga��xHwiq�bN��X�V&OL�˳����I��o�o�Z["�[E�س��ȶ����i.�iX�Oi9�TN��k(���/�_��=}H��ń�G�GI����f��ྕ|8�٩V�]�yl����{d���:�O��±#u�f\�o<���챊�O�n��0�p6�?{~�bI�ȸ���9�G����G�	�|I1%�sěn��o�}����M��J�ē�<JOS]Hp��	w�F��B�$�uԛv�m�^//��^<�n}R��6�n�ƕL�ԛ�m����i���}�I&�)6�7/��nG�z7m!��%�g��ko�R��6�~��fZ�M��6���N1'���!�\W�R�A�9���틒��$~�=�q��VIWG�rj,~K�x��vҿ^d�;C�p�R�]��<�[�K�#���Ї�1�RpiT#�~8w�m���.�F�x,��I��U6�x�܍Ǽ�:�~I��t�>$+He���i+e�l�3�/�'�����z�<Ku�y4�Z��m%~r�3:3�64p;�d�1��ؕ��Xe�΋,��>��5FQtx����p���$dtX�__������:==��bf������)��ێ���|_{<��0��+�uw��+><�
V�����w�ј:}��>4�Y��T�=^��6�=HP����d��/��:\~f���s۳ِ��	�x��GJD<�lV��������&�����&��{i�ٍ�w���RMj�\Zh{���������M����S_Nh^�B�y�W�v���&"<�����������9m9��d+�0�['^d:vn��N�t���%�r_K�Ä�/�a'D^Y�]#-��Vm�V��7��Fd��BMby����=#���۽^di���V��O������+�s����ٝ�#���n�a;��嚳���+�]Zv#g�|�W���u<��.?}���1E���Oi�I܋5��%��<z&��Z�Af��K�J^���M�Խ�M���:s��DwN�tM�����?���}R-��|��a���`>��y�:�\����*~�-;0�9��V�f��dG�����LC4~�g�P�/�G��}�X�ߧ�Yo]�͘;��Ts����.����\�_�ї޷���mO�,�a�?kތM� �Ә�ж��a �>k�<Wi�v��A	r�Z��T����k�}�ҝ��m��SC��H��;��kZ������RI��۞���{7;Ӈ�	*�5`��3�_R)h�J�������ZN_M8�w�B�Ϻ}�|gۈ���Z"��9�)p��HdJϯ�f���v
����_`�t�7��0H�1��yp������,aA��Q_}������f?�O麲��*w6���2ؓ�*�:f�@X��%q�t���氂���!�KAvF�S�א�M ����e�3:q�{�����J}h�4@�q�l�6˓�����^�Jwћ���bOa�Cs6a���c�|Q-T�+�'�LӒfbN��AS��%�3$KUX��)2�פ]s2��w�Ǚ2�ǭhl� sW��Leb襛�1CB�y�������@�O�33{�oX2��W.��i�ߓ'L�>>��uw�:Y=�����E+t�8��b4�EZ���ʳ
�RIڍ9���ŧ���`8SG�HL��,�׸~CwP�k1R�ƿ;�T�)�����5oGAIMR�Vp���a�*��o���3�{JJ�Z�=�x`��$'ǻ5e���̺u���kfc�P�I�����k���{�M/M�}�3;Lߟꉽ[�T�;uˌ�ڝ]-�q�Xɨ�i���\Ɲr�O|��a����9��5.��[��j�9;�S����BrN6��}�s˼�=�'�N�l�I)	�A\��k*ߩXs�����[�O������s���R�kZ���F~z��:�`���7ԥ�rߌ������tN���:z�m1����{�����:��;��$���~��Sޑmɾ1��[,�S`�<c�,�A�j�-���1���V}�틧��W��Jʌ=���)��=�ә��tU��I��r�p{��kxPz9s��3%��J�-���ز����|BY�[�^��,�����r>a��Pډ�Ė�a�l�N�4�x$��>���/'�o�O�}��^��,��X"����ʓq�i�����En-�d�!2+���JQ��o�<2�[6���HBnZJ�!Jp��J4�^|����z5�W�R�V�|^i=sVD�YS&�X�p�(��+�Ε�U"fzU	�����)$=3*:���hx��/y�|���I�w7�qŽE.�������{���M�c9�iő�K��׻�j���K1`�Jڒ�F:\G�ZO)�ػw�ui��3��ƻ��E��̺5#��GTTĵ��\÷Y����ޜT�L��}s�:snv
��� n��.coݭԻ:�7������ꀅt���W��
N��F\���~�̙�ʼ��J.�sc7�%���GB[݈V�Ǚ��4�4�r�Y�2"NwX�sf��]A$z�,����,���'����_��Q^�Ͻq����80��o�jw�n��?A���Q��c�O����;�+:�����:�T�6z��׎V���,���U>�+���4L��c��w${�f����4f
�\Sٍt��x��	3;<0o�{�u�w`K8�[���b"��W/K{�~y����~�s7&�D3t�`Y�k���G}��p��X��`�ش��ꊬ̇�I=г���b��M�V4�k�3��~�6���-U�<er�V;y+M��7��M�
��k�'�J�r�1nQ�D3��*�<�;�JJ�MM�k���z-����9S,a�ݾ�\���gh�<�;�V9�&Zp��X`S#��뛚��XJ)���jn@���)f`�S����F��?kW�Z�3	��YV)�LX�Y�f1�Jx1�M��$�l� 6I*��M�}�k{�!g���&^p��y����9�� \./���P����V��Ql��Ig,�����ef��5�"���ջ���מ��}VgR/7~���v=��V~�ߐ_=�h#6o�@�=�na��}�{_t1�~rַRc����MJ]"Hq3M��W�rk�l�s����}�U���"��4������;�WY�*��	�TZ�Fm/ꨀ�s,_>���k�U��1��,҂�����a~o���j7=�t�`�;��u�m�*���-�i�_�E��G�آ�<y�<z�FQO>���v�P���jQ���f���o~[�o2v�S�ڰ�l?z0V�A���,"��"�e̸��V	��Ku����Ӹ���D���o%�"đ�w�`ɯer �=!0M$0�ToH�;�i�`%�R�\��>z��0Z�.�3<�S�t��Z���lŤ�a'��c�m�}���&�㖱���)�{��H���7��������Q�7��w;Ր1�Y޹j���0�L�-�jayAfe�m��9�g��^���61�̾�fu{=�=��	N�N`�,�S�%��J6��"���\�ٕ�a�`˙�W,�>K�����0�yA7#RǍ��n�'yh9'�q������v�=�^C�\(wj�RJ�ʢ��z�9�JFb<a+�{��=噞�k����+��@�a2�>7�?5���W��J�t�:p��3�#²o�ְ�����-]u��#�L����%�V�9\xb,�!̼�����ȰM�ψ��cH�=d�ڲ��f#��0S���T\�r���O�]_yL�J�y�侪r^�'DY�4��>��;���������ȊXe;���X{�9�P��q+�̖��Y���ɨm�d܂1��<ԋv��p����Ɠ��&����ObWt�8q�Ρ��K�;<u^�-�D�X�}��)'�hd�ms#� �}���g�celUL~'�O皿ui������5z����ſ(�?��!�n�~���f^Iޡz"�;A�x:i�٣�ޢ���ɵ���K�Xg_g�Ŕ�����e�[4���L_]�����@����?�
�~���"ܺz|�T�I���DS���e�0c>��R��)IQٯ*�����]َZ�ke'W:U-:aԥ��mz+5k��qvS8�-+��U&(�)�^р�#�>YI�bQ�O�H�2!V����
�X+�}���+u��H��
^�$�X�����F7� �e��F���d�1��㌻�̗we�m���X2HCU�Y�2�`�S&0�4D%r�]"��T�����n6sc�1(��,D:�H$#o��Bhl�1�	�W�$��Y�6	�F�j����
>>PX��,��"$�p�� �|���I���b)ȕ���ji4�#�Q�3 HF�c]�ǩ�m�ŭX�l�%�t�I�F /���R;��"�+P!xCi�U#^�a&b�9
�HPB$�x�n4�RpXf$�L�Aܗ��t�PmD�Q������d)r����"��{Ɏź��H$��i�����Sħ� �n&C&�1���ƈ���K�lF�i��$�G���1"��5�>�1�R`��$"�`�[P�'��+K�QEap�"1!a��8� H3���1�L&��PM%<i)(&��n&� \���G.BD)�h�c!bN�J\��#r�%lk8�-E����v%r@�a8��#B�	&�1��L��&��|E4��0\d�Dz��p�m��""ʜ��%BML��D�AT�(*�)����^*��p1..gof��$l���(�c� %$+�Iq�� ChFۮ"`� K0��]S�C��q,mB�M��.a��������T��B]�+/��U���%��l�&e�wn6X����Sc�8��K�t�E R9\���(\fq��rD�Qpu_��q���G���B'_=��>V�XP���$Yi�E���q)��m�6J%�[D�!<�"����'�1��I!�S��a����#��kS�l����j#v�BI�Rd��^������1��Bb#�mw�1�ʺ�ݹ	��$*$ʡ�t�AD�?�31ò|&� ���a8�Q��24 BF�n�촃Z"�'��cd�\�܆D�&���E�SK�4Sq��*&S)�bg��Ctg_H����#ͼ�g}�E���S�^��s$�mG�dβ��U�������S�������Ip�T:�9�jw091w1lf�ͣF��I$�i$�I�4�I$�I$�I$�$�O�'I$�}D�I=I;I'i$�ԒM��x�N�I'�'I$�}I��I&"I�I$�I$�$�$�x�M��m$�Ēv�I=I��I&"I$�bi$�ORN�I�I$�I$�I&�I1�t�I<I&�N�m�n�I��I&$���I�I&�I<I��I��э4�%ܱi���(5�_;�$�v���$�$�$�O�$�$�z�N�I'�$�$�z�I<I&�I6�I�M$�I$�I$�$�I$�}I�I$�����m$�Ēv�I=I:I$��M$�I$�I$��N�x�M�I;I$�$�i$�$�z�I$�LD�I$��I$�$�I:I$��$�I$�$�O�:I=M��v���m$�ĒI=I;I$�ԓ��v�I7��I3,�)C$�&�8@Rͅ+�����|��O^=}x�M��I�I�I$�$�I$�$�i$�Ēm$�I14�I'�'i'I$�}D�I$��I$�H�I$��I$�ԓ��I�I6�I��OI�I$�I$�D�I$��I$��N�IĒm$���ORN�I$��$�z�v�I��ON�I$��t�I'�I$�m����$�I�'I$�I"I$�bi$�ORx�_@c#T��d� Nظ��Дj\ I�)"C�9����^�8��I$�LM$�I&&�I$�I$�I���I$�$�I�'I$�I$�&�I$��I$�LI��I&"I$�H�I$��I$�ԓ��M��x�t�I'ԓ��I>��I$�$�ORN�I'�$�I&�I<I��i$�&�I$�$�$�x�M����I�$�m��m���I$�$�I$�I$�b$�I&<<�Z��>yӣZP�--R�'2:�(���P�0�J L�hP)�Ei�����C$�Ur � 22U�Ns9�6�u
�@9 "fb�d��&B�4d� R�A������֊��%$_��=�oݟ�7��W��Kv9�sa�c6�ZM4ҭ���M���x���2}�w��Ç8p��nEt:(o����ñ��������xH�x6���:�t����}��y�v��Xڧ~C-�g{�NC|o�o�?L8m�_V/e>�����۾�S���s��ÏC�����C~]I�w~-�Χ�t7ލ�����;�p�Î���Í�����O�(����o{�(��wܣ���"��I�.a"��cD�2Hfc���<S�X3�$;��X�������sX��I�\�$�P�DE��!;b�����1u����H��
��0äO9����1$�m�p�d�����<���,2#�8�ቧ�-����"��O�ӃW!��d�
���"���0� �l.$�3�n4�Q�l6�"3j|&���B����Q(�}�M�`"R��"&)$<��`�0��r�Z$�@���'U��w���NѹE��B���Ngh�#W��١4��H!�!�QWY!#�����d5}Q$�Y�][X���p���zd5y�i#��3S0I��-8��1''W
|��Eo���!�
A��j)m�� \"1 d�J��rCd���DF%U�'" ��d����1���0�b�M#�b⸖BD¡JcQ��3�a|��eQ0�����!2F��H�T)FYi:!�\�ca:�ɮ}q��Lbq�8��I$�LD�M��m�|q$�$�}I��I&"I&�m����I:I$�Ri$�I��I��m�>I:I$�Ri$�I��I��m���һ]��?���~�?�~d�*���)O�����>y�B��a�F��
&�"%�Y�2��VM\��k�"V�5�f),�K,�9�F�F0���#r�\L��-Ȓە&I<X�����K��q��� C����M�0a!1������X@�t{���i�o��h�hh3�AHw�@d~��Ӈ���+�A<�j8v&�E쇽�*��(ӻ¢<�_l�ӻ�y�Q֡B�=���!mi2Ž�r��s+���/`��	�ʷCj�pQ�&���2�������ñ�x����;�ܣ(|3w�o��l��_�����W}.fT%�!Dwy�5�7DGF��Ѯo�8B���}2X^�{}�h��'�@k��/�z\Mv��<�'!8���|8���w��_Q�k���v�2�D&�YZm#Z�!�"��x����gn�Ii�F=�^��ÿ��IxuSB��!QR�t]���m��~-������M�?O��rq��5%Y�"""�ڶ��+z�Z$�h�,��KW��y�-;ؘ"�>zۧק�"x$�C #G3K9����	�ط2ܕc�q&6��xd��,r�L�5�PଜM4��>��`���&s|��[r�!J�J 9vI���Qc����%�	٧��:����Lƕ�/����I�2��=C�o|6�x?��E�g(m.���8!B��;&A�ކF��æ���v�#�cwY%�-ƌM�с��u��8j�����3|��ũ޴�tO��(��ų)/��2�_����çP�4@�wܺ������c��W�������^q��囮J/�]�������['1�ٲOR8]ӋU��q�),�(56��$��7iv�u
�,���X���AQ��H���čI�%L�ҁ�Ղ���*�P����R�x�!qHB-\h����1]�-G����C�T��yur�:"""0��D��y�'��!�M�"j��s����ќ���4��sl�·�w6�K������N��C�_�+<�ٱf��9_�>L��s]3D�mi7U7f&��\��BB���ΔZ��&�a�H�����5#�c0��jҷ��O,;��ir)��P�n��Ųss_v=���� �4���9�� ��м龹֚��.'���ۆ��x��J'�{�UΫ_:�ƐK�x�z[����]�"��Q���LR�������Mq�\�F#9�CL�IV�ދ,w�Q�xq׼�;���L�a��``u|����(,����)(9%F�9��������o��H�G��x`���fI�'�A��K�7��Cbg���k-]�sn]/W���ظl���QԦ�s�X��h��c��.]�B�f%ݑ�T�h�`�$x&��=�ڵ'�kx�^�'j�Q��3G�u4�I�/�F��@m%��y}�R�Y���˙���\`�eə-�ai�/1%-�L�5�8^��77������ib���D�"��7��s�������h�Q	ZC�s���K&9(�(�/��������,�[�˷
��Y���х��m<ƹ&�3����DT|95��W�J_z|�޵��Af���K,ln�H5�޵)����NV��|e�r�2����3E@�kZ��䎤P�h���u��,3��wf�8W5yD���ٽ(�Sޙ��*;F�sB�,�Iv�\;2�Ô_(tgo�o��df"���P�篕B^3��]5�I�Ӊ��07�&��r2���_!K8�[��<��(1wr��(����0�(��L;S�c�"R)���Iq��A�z!n7r+��k,�JL�2��St`���̍���zbj�V"�LU�g���R��rT�)�.��8�%�!��h�_k��ޠ��?��w��'�s�gC0�M^KS����ӹS�'eh�k���.�^!D��gk��d�y���U�U�v�n\�$��-�fR4�Y��j8������ue���|_�&̹�xR&=(�Q�{�c������q;��ԽiEW�"""3�tV�:�eS�E�*d�r�ђXf?L Q�[�1b��]�C=B�B����ZkH���G翳��j흿�u.�8,5ɬ��kTWtx��?pt�A�<���	�Sx��\�#(��p�|3�+�
�$y��!gs(ߴ[�9c݈}+[Ú�]����7b}`�Z�R%6@������+���M!����_�V!(��5D��F셛&�P���2j9&Ѩ�$�n��$�#Q�b5z�`o�J���
�Ȣ�¸!�%|��"!�W�A>B�N6�#����5G�A�d��c\��9�4�O�����юtsI��M9:sF4箓��|t���h�j5FѨ7Ě�F�P֥�QB�Tl�E!�$�j#|I�5������R�H|9��>u<I�D�j5�F����̣�|�Z/�%(B��>FѴj7Ě�F�MP4�KF�CL���F��4GQ�dS� |B��b
��I�~T�ACB
W�'������5�l�5,�Q�F�G�F����(�j��5�5D���<I�j0�@�j4����y����
���h���� @��/�p��t��nO�'��~���__No��yw����å�MX��'��An�8�Ț�8�������҉(�ɞ��z�p{���駗��QF�T�̑��ڳ=},��398��G�(��|t��a��ǆ1�i�q�c�Nݻv�>|��1���1���$�q�c�pҊ(���aFa��xc)$��1Î8�nݸ�c�lc�RN�I$��i��iEQ��⌌�gh�3�n�m��v̌�ɔW�<���: ��	!�J�i��<��y8�6��F˚�s9�j���q*6�ݵ>cU��_4�n��4��Kk(3u9����V���Z	�S��]<�wxw�E��y��?�Q����A�UaN����Cpy�Q�pAB�ѭ-�'��./�U��okO�ʍ{��N�p$6�\ ��
�N�V�
EZ�h+z��7ܕ$�2�{�"�U���3ޢ@m#��a��_�QP'1�d
��LY!�&8(��0@ˊ�D��Fv������e��fi&M��K�}�7e��� B!����U�u(���Vx�oV�9HjwL���Z�5�n�~�o ð�S.2˺���f+ͥv��49R��T�������Gd����W~���@r�A�O�ӛ�d7	F�5Ё��3�B��[����T[�IE�6_bT`�����&#�v�*rcS|%m����{�f^�5�X�S��)��f!��+�V��^��2�ł�JGn� w��M�+���Fp���ّ���<�xf����A4 ��qA�zĕ��"�
��@H�f,�7�� � �	R2x��.NF��,�D��q��
z/ǖU�r��I�(���x�0��al��EX�Yf`f9O�ÄB!�u��nf8�-���m�e�Yf䚠h�eW�y�$_B��4E��3�uF���L�R\�s/tVښˠǴѪu�r��5���5ֽ�ʮֿJ�(]I�5BG�h�R��A�j��kҏt��q�P������z�lZ�o�9k�-6c;�Q�th^4:���`?5��w92�`�9��D޺@x�j�k~��}�e]B�+����X~��쵻�IU&�&�C��.��=a0�[7�#�8���"�E�|3�������I�\'�Z��5N�V�^�Y��!�J�[UY��hkаv�b>�(4_s�1Q\�@w���?,�(,�\�&�J���U��mQ�/G��}E��:j����5�/������W���Q�ƫwi�D��(�-.U�r�e�H65�.�E���4�G-�l,Ļ��lƁE�W��9�V'Z,q0Q��`(����Ʀ��&j4���<����g~����e����*V���C#){���
 ���VU�A��`����TeZR� 4~���PFN���Q��v��W\ )Q
�~YP6��I�P}�Aq]F�������m�����/}��egE�(�C�I�J�W^�xc�d��qR��u��Po�:��FS�5�}������Ъ�<?y�RJ��z6�DԺ	�P�`(4`t%�I�ɪh�l�����Ϣ�[|��L��dQ̷t�Z����>��v��C�}w�k7�I�i�D�����x�e�TA��	(8	�Wʀ��dB�ܲ�cg�i������	_��E\SA2l<Ѓ��G.��iJ�5X�;�A�Qcʁ�u�����`��CL�pE����.Hv=�}�.������o�l��E���'Uy)����w�A# B!���XQ��|}j+�e#��0��>�)ڻ�H5��G�Q��#�F��ih[Yw�$/i/�	*�S�DW bM����(�"`Zi�W+��uF��Ј����
��_�֥V��Ѳ��#[�U�v�`-Y�B�Rhl��y�c\J��<U�~h4���k�A��Ul�ƾ�9�Q�O�-eQ���W��5c��.��V��j��H�� a�?'�[_���5i[�/�%�]��4@y(A>��}i8d�%8�+6�՞��M���#1���:�s��%f-ŻE#pul�il[f\&Yy�~�X3�X	;��F�
�xڣ�CE�-�l�D[�����)�a4��]E�� �6pQI<!+2�r�n���a�5SI9��flK��!�BTi�)���SEm�$D3�V��zM�D8X(5ux""�!��P^�¢}`qw����Ё���?4��U����@֚�B����P?�[��~x�������{v��d�0DP�i�S�'@�0��t��$�i��UV!Z�Ak[����u��]���1C���\����6����R>D!�+��as�e���������ac$d���B�8�&���89��f�{�t%!Y�bVU�ƏlSQh��;�>���᷃c�df"�Y���*ѻ��RI'�Q�:@� B!	Q���|�����w[����<������f.�B�rSi�.�1�v��݊����eu��=���aT!�jB�z��X1r#�<�:v8g ��ت��c&$g��)B�h}0t;������
64-m���%�3m�	v�Yx�a�6�yy�%���wr��	\j�i+{�?����u�ޔ�+M@���5ƨi�k�J-A�'�
�8���xPp��Y����v=�=�.�Λ�x6;fFb/L��9��!ӄB!$�X%�h�(���:�
 A��}��#A+|O��1�b��bb9��e�5溁ӡ+�%�TK���%Z�����4ct�m�!�"����/1�5J|�ac�WW��~����_l��J��p����E�D;������QF�+��5��kMf>K���P�}��D�n�h�;u��)�8qԞ���X7���)j���=�`"�Qi�w�:5�������23z/s.E����$H$	�Q��~�h�/(�kgQp>`5�� o҃����1 `.S�����0�6��1�LsZ��KL�� �A����ՇYQ�d!�-.��� ��P��b����y"����>�p�ƺ���[�����SU�7��?��*뉹�{s��s��I�w�Q��S��q�Y���/�(h��!�=�1�9�Q��Ɠ�U��G���v�>����"`�1�A�:�;���3N��Z(�����p��Z�J��+> k�i��LJ�A>�ɵ)j7d�nj5ӴJ6�$�5FѨ�x�ɮR�@�j4r\��ChiO�S�C�C�@�WR ��"!�C�8�!��%#PtA�:l����,Cd� �Q�#��Hk$5�j#k$5ن�Ɇ�:H�e��$H�n�Fɨ�jF�P֊�(Xm�)J[&��[&��x�#Q��Q��H��3��!h���Hq�RKdh�$ݐ�j��Ѩ��D�al��E&�|I��`���"�t9>2Kh���|vC��G�g������� G�AO?@D�!_4+��-?!�4!���*���@�!������I5����5F�Q�I�&��ɨᮒ�C��d�.C�I�E#D$l"6h��D�F�B����C}����N�Yet�U��ʩg��3,p�^�n�IMƑ�[(��_xuO�e�
�n��Х�xw|^���<�V\>��i
�󹻻��.F6;(a�<j&� ��NXIeNam�l���da��1DS��)�b)�=7M�k�EnG�Hm%ND�,�� ��m��Ij�\�\J�cA�lL�j��R(ę���̊��͑�[+h0޼�!h���׽C1y0�g	�a�^n1�҂�<�""M��	�\���;rwf&�n�6qf�i������wSܽX�?���ɽa��+�:�a�B�0�=�
�Cq�[���h��ڞ�81d+,	#Ɩ��B0@J����p�P�k���S�8c-�A��XA�63�(^I��L�}��m�$	�	���Jm��p�ˠ�p�\����aH���Q�%)�B2��[�#xShF�J[��d�,���0�eǛ.^�bX���J%�5fX�8��.�#r�c.�KU���\qr1� �E&Ɋ���a{s*��'��K�(XQ"��)B-����&&i,�BJ-�*�BKt��h�5�Cd�V �f�Bi�ϢD+	'R ��A��MH�
.#�bB*đ�		@\%���˼1���9Q7����K"0��Ԃ	h�"�B���r
ˌ+I�%�*EHid	f[	���nI�
i�G� ��0���>4���2RI$��I�x۷n<|�1�m�c�<I'i$�ԚI8��q��c���8�Ēv�I=I���m�>c�1�㍤���I�M$3N�8pӱ�1�2�Λ�5��#1�u�oy�������
�OIQ.����GT�#M*%
�I��(���j�NR�*��`4��L����dԕ)
��Kʌ�yM�.�Z�6A:$	�A �k5͗��8˒^f�ˬ.�0�/TH�+��Q��4}Ӧ��4ڍQ(1�����yĦ�(�Q W��t*����*c�Tj�p�����F"+[��4l���p53y�eѤ4f�L�I���]c����c�>�9
Qj�@yA�h�8oL�h�O�a�~�+mQ��.����ނx4>���c�?��~5���j��4���DG���+������׺�5�r��RF�ԕ���u�n5"BEfz�h�K���&��Y�1��������.������l�ǜ�d~g����bX�H$	�Q�@��zU��{+)����k���f����A�2��lp�R�zC�uĪ�}�%�*|֎���%��j�5�$v�1�٪2��e�m�5���c|��.�x<.w�<�H�a�D�(��_d�&PH�|lS%¸�@�d�Y�� }ڔt4J�Zta,@���]��4
�TtA?J v�%oi!���Pb!p;��Ӑf��O�sEz����/:n���lv��zF�R��bn���9DH1�� D	�A�ҁ���N��(���;	�Dx�(<5�@�Р���P;��+wC�A�`fV�n�!>�0����+M~�����9F@�?��m��L����B�HG [}�o���ùa�n�~���@�ˣ�۫�#zk��C-ƍi��ƛ%C��<A��S�����W���<r>�3��ȥ	C@p>�*����"���5G�*9���=}Erb!�u&w�����x��lv̌�\ԞS�$��^�bA �H$F��I.����Y��)��:�r%GT1 �;�����&	�P�����bs'꘩�0à�B"r()�$ l�����?�[Od,:�Ѵ�Ƶ�PF����ۣa�'�:5Z	�����@�2'��*=TAy���Q��s|��N`�9j/��<�� j>��YG;.�}a�P4:'eG��u��S�8�A�t���)(<zA��Pz���\@��J�0Q�������4`��:�Y t��(ڊ�
1A1x���t|�}�7^�ّ��~S>Ȑ�Li�K�4��M�Iu[+��"�J�m����YkqD�*D
3"�s��O-+�YS��bp���A�119����0gXJc�A&��Q0����A4�VL��KU�U�I2I��p��&�i��.&F�! �H$F��C{%�-ę3����dԲ��E�T���������eS�KEց�kyX�ڡ,�{(���i+��tk�Q����6\,���魵��Q�U�=�db�Hj�򤃡��8��@��	/*C�CbR�n��m|��7~�V���4��@>h�sb��X:��wW.<�t5ϿOH#�tA���o �eJ7�Ж%�uuZk�[����ۢ�8�$�sML�`J�L�� �Ѫ%��]cX�����f�Zk�[p}*4��	�y��1�x�x6;��;�7�z��ӗ=���r��u�+���� �H$	�Q�7��6(��G�γ+�񡮥��s��K���m�7���]�Q�mQ��U��j�Q�k�=��EBH�\Q�B�W%P��(��Yh�!ё�`��?F�����j����r��o%��K_�rM/f^.kB��"�	E&�,(��@�����I�ٴC_��j��B`пfI�Ee����`u����Pd�q�X'��{Qܐ5D�8����-30t_;�Р�z�����>������23s�z�淋5_�'�A �H$�U�������ݙC���y�AE���;\	6:|�Bf1C��	�!��${�W51߉�Tj�D��P���Q�J�Z���5��v9�.I��Uv�F�_�U���&�������F�]V��J	b$�׋��̲1�]n��-u��h�x+�M5�b�Lq��[b��Ix����.�E�yv7p�[">Hh$ۂ"���3�fssY斻��Nl��t�����W���0�TNQ���0����Z��aԞ��'3��#�d����0�����C�7�����|n���ާ���vc�咾,H$	�A�ҁ��d�7O���K�I���Q$� �; yG�ߒ�9*�o[Z�ϐ�5R��Y�BJ>���N�jg��{0�.���/,���!c������!Z�½��xg J8�ε�+���teS�����Z+���҅��r�5���=Ki)uE��g1T?4�N�v�~j�2q��I^�{韷Ym��e=����o�+�a�F��r~Pj��pk淟�t�����#�[֭�
�h�>J;B�'�G��.bC�o3�p����u������7����C��M�y,��"U��Q�Zb��)m\iq�f�EpBb�$LF�I��p��" �c�^) Q9r>C8TlI�АH�R�j���ጶ�yy��:$	�A �ksQ�w�jN�$���&\����_ J=�pj�&g�G�^.�=ـ6�<� �c�
�%X�l�k�Q(�g�!GZ�B������i��M��W䦩({���(���(8�p��R%s����0�&$'B���q��ޤ��d��kCGG����e��k�maa��TQބ�R�`ң��
%���W�ͶY��8X	q��m6HA(&�F�� D5#�=����$�ll��i�e���+8���oޏ|n��#1K&���*^���/�`�H$	�Q�ֶuU[�h�-~�\��5F��` �趾�\GE�����TyF|�^�n�|����Q>���Jq�S
Ƴ=.���~�Z�W�i�Y�>�N����0��}�}3y��&1u@yD��|��|7�|f�$��xW�^��Wp�o%�d�J%	|��Ss��R�3G.!�5є|�5+�x=D�5�����~;��ޫaq>�^k��d��i��Q�Q>!���ڟ��?r}�9u�L]Aj�~>I%3����AP��%�`���B�AC���3���k��4���ĉ�'�5R�욍F�&�P���@��zt����9��:f��k�Ni��i�@��KO�����QJ�U��B	���|�䭦o	#��j��G���j,F���vMi4������ӚM�s�h擎�Μ����:}��8BF�vJ6F��&�Q�5I-���(�E&�ޒjF�&�5��i$h�K�i�.M�=d�DJ5�1FѨ�j#p�t��Q(�F�6N&��$ݐ�ɨ�&��G%��4����i!ʝO��1��:5�"~�?)����QJ�$�	�+�І�ڒ�F��ͣ�5C���ɨhl��}�|vIG�Fɻ%!��x�5�H�1���#DyQ���b(;0v�(;'f��8�Qj>M	D�A��`��J2��a.R	��yX�|�x�Our:��(7p�҇%h�@i� W�-:�J�q)�����
��黀eʪ�eOCڋ�3I[m�Op�|�h��y��ZGr�Lh��F�'�u쳾���͐�ģ�v�rzB���&�B� cUīx�8��J�z�Ѧ����[@ĥ*vN5X��~����ܪ���r�u��(���0gF||�I'i$�ԚI6�m���1�x�8�i$�$�z�t�n<m�c�1�㍤�m$�ē��q�m���c�<cq��M��tc#Æ�8iPb���p��7|n��#1$�f��]�6��ď�	bA �H$!(�_��>��(�}���J����%s��S0>j�d����%|��f�:�����K������DCMgg�kf�Ǝ�����yA��ͽ�V�18�2�$&�#,1�@&�HB8&:(�G�HY J�ݙ>��dt� ����Q��jQ���[m��%�#� e��V���+�eJ5�Q�`��7�#־?}?]��ܲ��ZO�	��^ӭi�1��6f��i�<��U�8��s��ʡ7{ڹa���[�E!�}�p|>~�7^�ّ����z���H|h�!�J#���h$��T������?+^ȒW��s��9>~���B�\+�-A*F}Y��I&�P�&���a�.cP�j��	�E����ݵ��O�zI}x���q��A����\W�P��)�R�|��7GOK���.�b�� x7W`�Y��=2�D���Y���Ĺ$+��Уå"�@��9������5yEϋ!������8$8(݉�#��{�}�~�6;fFb-�:��K����+(�	��Ium�S�$�E��TD�QU��I�,Ʃ
Fp��rca��D��
t�HCM#�j����j�[z���/�"d�	qĄ	2\���U�M$�������B!�J"L��*՗�$��J��r�2�����{݃֋� �We�֡��/��o����9�DXB
`C-lv%S�g`�u�4�G*蕷���fVWz�B�C����(�0r%�H���nC������r��$�C�D(ӄ�\I��
Q�*�N�iE{��+܊U�V0��yGa��.`�N�TORD�(P 򿏥���B4�Q�"|�B&hҌj�E4zV���xn����j�I��Q(����#��i�"����Rr�tw~��ٻ�k�#1
6Ѯ���X�<KJF� @:�:��x��$C���z��U���w �wb��[J����=a][m���5�#�B�Q�Uo;�oV҆Ҷء��Rh�4�^bnC"�^�|l�!�J#��(����,��*/��T|��QjEi��A���"_N#g�;y�����M[*��_�g��W⨪k�gT�[�f)lV���.K��e�wm�!`Lawl��n\��ܵ��L��-�X%��`&��!���K�\�D�n�]�A�ld����4�H�lvF`!:�G��R�RRFK��$�ܻn���F��ܶ�#.�7M�T��B��7W��Ż�$�ȫcr�w%�B�]\.�I%ݤ�	d�!r�!t�2KK�	Ct��ܒ2�kikvE����/\�%I��]ƮTmbƑ,��1.�r�7r�M˂6L�e�|�MY�D���x	E��׶�}tOu�J
���5�ʮ�H�� �%�|ю5��I�e	[G:xN}�5�j��"��a]"P��Y�q��XY�:�-� �5y�/��u8]?�΃�%B��$����v]�9�J�p8с����~�����@#_�zFz�˳+��{��Aܜ����%�����Ѵ?}��wY�v̌�_g�����{��./#OHB!��7�Qa�i�D��<p�[cӤ�꣤��ڜ���y~%�E�x��\���C����6�6h4j�&:.����J�sCB���bd~��&~��ֆ���.]�fr���.�CVJ�m���t�(�.��~�\W��e�;�%_5�+�G7�;0�h�e�U`]5T��G<�����^>���%��g�5et�
~��h#����xCcP9 ����pd��4Oīy�hh���F�Z����X�q|�L|6��x�l��k�#1��4�t���B!(������
%҇)�����4э�W��z���Mv�yCDk��rkd�	(�A���A@��� �X�(�Ƥfd�Np+i��@�Zq�@�s����g��K^	k�iE�4�)�۳����w�������*��͛��V�89E�U�ܢ*W��л�ce�8T@��ҍ!�k�)[?�|ە��MƎ%��0Ϛf��lC�߫@q��d���$�HG�$���#"f

�i���ڢO_Q{~7l��n�ّ���ġ��D������*���P�a,(�M�����[( �b��L[^Z�˙1[��9��zv��m��%"v���6c�U��Cp74��F$���]��Y0U�D�Y��@� B���8�,�E
U�"!Am!6K�Y���*�_�+���n� 4C�r��>��tv�)�"-e�;+�4N(�1Tj��ށ�i�p�I[�)�Tq��ӕT:M�x{U��󼅅�7����S
�#fʂA9 P(�48�h9E���B�r��J��Cau���㡲����\�Y��z�H��C�L_�E�	Q�g���Eaj�rDd�}��ⲿ!ˁѯ���D�>j�a_�N5��s��U��ew8eo�훺���23t��R^��X��Y�#DQ!$�I!$�`~eX�i����6CMWQDb������fQ�뱁Q�A��RVPד�8ɩ,�H�#F����]���$�S${����BS'�m�ԡ�6ՕΉ+��q�{>��V��Wf;
MM@��iK歘HaSK�4�����LP�\EV���i��|���m!���@�cF5�CP��~v���{�gl9Xлh�x��CXWy��X~�Q��xeFﾣf��4VTi�i�5�p�w���7u���df"��N���R��U�9�4��!�J"�����<��\n�tS$�v�F���=Ϭ=DX�o�o�F����K� ��V��r�b��8*�>��0�'�&)xy��;)�6��m㕸HHp�
=�1G� ��&5e�&��?�B	��Ӳ���46]G�5�"Q��F��������W���0�A���Q��u�e]�]��Tkf��_2�~��X(�F���銃�1h��|3������7u�����ߎ_._�����|h�@� B��=��Y�%��p݈5i��뺣x@:��nX2�ŹY-B%�3wZ>�;C��7Yd0k�b�Ӡh�Hl��3���^N�E�[���Jz�F�W �^��J?���1W�&���TZ�f����k��o��<��:���S�}��T�App'��CV� ��$�8+�}<���J9������_�2I�G��F�_����P��R$�*Z��gH�I�C�C?Ak�B6MF��(�j5���b9����M�7��H�j7	:�C6CDj4�.C����Q��D$6��UJ���>D�
���,C�	_h���>�
��*揮t��9�q���9:1Ο9$�1��ɂ5�[&�4r^I���6�!��RZ7��j5F�P{I5��MB%��zI��d��SKd��i$h��I��G��Z:���P���J6MF�Q�m����D�cd�j(�5���Qn��9Ӎ-��Ϻt�Gy�y�ơY��	�|%��O��O������u"!�`�̑��Pj*�DQ��p�#�o�'#F �	>�LG���#�}$�}'�$�#�$��l���i��O#Dq�j;0v`��؊�Iك�"�����X��>���n����Д9"J2�1��f��3�R!�]�u�6�Nx�=C���o��.��D�EAm�8kPQE�ؤ%$<���s�QīȘ1&K�T{#��[!�^�L��+�#)�]�K�Tȩ�>c#۠S�4o�$�V�H́8#(��S�y)#��In��v��l��bvG���I<\T�$�#*t���Q�AxǠ���\72�XEb�H5��,L�F@�E��w�8~�q�E1E�$P�$(�hw��B6�7!�(�*/
��B���)��8d����v˨� <n�nC(�d�X��J��\q@db�NW��0�˄DbH�[���u�]?�^(�,b�1q��EG	P�Fa,�!�P�T'�ᡤ����	��2dH"<���@�J�Vp��Ll���B�8����%��������Qs���zVH_�~F���l.L����Ym�%H�#��(91��4����؂S" �'�t�lB"�%��h�o|G���A$�5A+6r6J��IG"I"q52A�đQ���nrK���$�0Z�D�II��e�m��*0FJ�|'����c�����i�Ie(A'�	H5Pl�ۑ�D�I�0R" ���b$�bH�m�_'f�eM�\[4�*��S\�\DҒXx��Yјi�I&�I<I:I��m���cǬq�i$�I$�$�&�q��v�1�c����m$�Ēv�mǍ��c�=c�;I$�$�i#(g4ᤆFb3�p��=�f��ۼ�#�x�JI�p[�E!Zx����96?P���#��J"ҁ�L�KB'L�j0o'�-�-�ae�/T�5-�d�,��	�.�f��	z��@� B��{�w6��\���)��)p����������P��q��Pe�{�P�<��+����PHW�ܫ\�q=D�{5�[��kt~���-t��HHB)^�R���W��0��CT}����\�n��F��"��Pi��l����R:����T"G5(�w�8�����=FL�b�uq��B1�����|B�<�\��i���A�nxC��c�\E���w���wY�n�7H���6����� A�F��P�Ꭻ�W�Q���4m\P�,��d�c�9�ή��XP��|}��q(�=��e���6��%*��"e`Yr�T����i߀�d�:E����y
��@��+O㏓���e��'��"ޤ� �t0��9�(<���B���f����e�n�H�]!¡����Zu\�⠘�
;1��(倗ܿ�G"�J��@�yP��C��_�>����n�wh�F2|*B�Ij%,R������DB!�G�<j�#ރOrz	�F��w�%�.�!�-����Y�e	���H�$D5CC^C���Q7��k�.�#����e��A�O�, �cl�W�(�?Q�˔~�������ߩ��c�M�ֽ�zQp���;jҰ5��{��}��W���2���K|]h��G��)h������ѝ���r�U���-I�_�|5�w�n�7M���z��=�ۯO��R-8a!@� B���~4�ѽ'�	��e��+	뭹�k�j�2~��2���?@O^�s̿̓����:�J ㎌���K�l�(�x�Y�����r	����W@�b����G܍�yB��5�9c�0�%sQk吜����J�}ٟE��H�Cn��P�9}�CI���qG��Xi�"����T
�У}d���Eo�gǈ�܇����HY�)�t��LYQ���Y���`Qq"���9�x}�M��wY�m�]�����O*f�yQ��7%^M3!�j��A��e���	G8c\.#e<�xLD����ؼp8�D�A�#��c�]�.JIY��&c�.2���$�Qs%^Q$�^`�p��aw�O��B!(��)�����s2�fJ��KA�P�R�*]u�n��oJ%L�*<� 0��@� _Dxw���a�:a��G. �X��<�8߾Qh�&)��5\.c)�f䯣;��j���t��7g�����\�'������9}�\���$!}Lip�ˆ�ݗw,�MԶ얺T�P:s�>	νb�j��߆��=�jjR��ގD���oΟ^ٻ��6�/�����|p��@�%��!	�v>��ꄔ����9Q]�|S�V�(�h�,�AK�IyJ��z�?��Z)QZ?P}ϖ����>᠔���WS�m�w���@&N3�>[���ÜևPo��֩u��.�*���}Q$��O��=�����&o�y��uWL�����2%.���n-9��>�-��63���A!��ts�������O�w���������n����D�a�wޒ�*V���!�BQ_�t�����G�5��|v:���Gd>�*:��8�4�z�V���〸n�����̺\;��ߊԃ��jm�X�N<S���k�rr��x��,7V��%���,�_H��.����D��Rwur-�CQ"��\LBc�ƫ/,���$	$��i �I��m$�s.\�2(�[.�q�4w�g�"fU"T�pg�F\���p���R�G�A'�0?}}�ʅ�s:p�����7u�����=��'��I�3]�DQ!$ B!	D|w�Q��ֶ��ˍ�v)<9���m8�z�{��]ó
ƤL/fTLd��,	��+0����Ȍ�|P�8��h��^�><�)��	0Ш�/��9">��C�n�����,����{���o���F�G�a�ꙁ�V}��s��#�R�|���/����v����z�[��u�5'���s��S�?%��s�u���r/��Q���Y���n��.���ˁH\��"%�~]���5��a����'q�U�JxY'��Y��'!E�Ee�������ڜ*.&V Bb�RI�a2�R���L�	q�`aD�	-(
-N	.F^C2��Ӫ���� B!��7��B;�Ļ��n���6�I"Sp�Q�^
<w������ED�Tپ����U���^Ro�u���r>����4R�k_J��졆Z��.��R�}A�P��Yߣ!��C4ѭo�{y�*�;D����9"E�T�J�:	�AˊO�����NS��{��B�BL�(2���`�a��di��m?l����Y�j�;���L)EAq�ih�tt|5�6���n���r{o�_�9;�w�o� B!��.�;zU�Ex�i|�9�#Q��2ε��.3[�}bf�w��3W�rUV��};�]�#��O(ܾ�BjgT�RH�t,�h��v��G�u�5]�8�:��߿��5BA��ɘk9a&)rp���*$��|b�:�u\�H���=���Gu����2�/PS���˯"X�J�R�S$M�2�����p^E:�$8x�+|s㕥,�ۡ��n��hm�m�p�ll�{��%�p�Çxx�O���7ѿñ������x<�~�Ս��6�r7C���cx<g��q��v��ޯ��J��oU��oŋX�L�:��9L�M2�,��%c��������tr�軽7ܭ��n���n�t�[=�w��8p����6�{��U�g�B�\4M'���B�^�����|��;[�L��~He��l{�R���WK�6c���j:�ؑL�R��:�}�l��5�nY����_�+���^�=>��L�3�0����;I$�$�i$�6�n6�1�c��8�$�x�M����m�ۇLc�1�q�I$�$�I'i��q�1�c�>�㤒I=1���cÇ6�\�tt��fݛ�����.O�J�����r��6NqY�@�%v]<^��n��\r�{��UfQ����~r���,���P��J���c)tӟpNt��/x���T���	֯,��*����;G�O�G(᳡a��p��o߇���>1@H�k՞N�b�^��-4St�ۿ!�ŇT�~e���\�I�cϊ��z���_m%|RW��hq{�����"����g�f�twv������)���@�!Sz�P��ҷ���.�_p<�\Y�e�C݈�Q�B?�LtӦ�љf��P���k��*`�#�����k^�2�����������eQ��yO9��9�������3`����
:��UFٜ��8�!��q<U�2�� f���xA�?�>�r�y2���}�}Ja� ��"�A���#�v���������x}��f�>oc��E�x�F� ���HY(�f&�K��2)m-�Wb�DD�����Ɍ������d�2n^5���Dc�y%�d/��-IL�ԉ�$a6T- �'�� 2J		arȘ*\����B!�'�`Q�Z�ێpF�,��\(Es�qv4�����o����v|s�}���L��lQ�%�9�p�D	��B���(�	듃Qp��(N^~��������*����v�3���}�c̿����&#ڢ���F(�~=[��ƯZ��KO1��f>�7!�P�C�Y5�2!#	8C��J;�x',�D�1ȇ��K���eRS=&{�(��I��m�]������.OoiN���9�K$$�BI$$�`���r>A=�tw{Xr3��$�!�?W�s��[�d&�M>'�P�/��0�x�9�6�4B���$����߿Iqߚ�e��G'-��e��J�2�Qƅ^\Dy{�X��̔�h��q
��
ƟW�U���{#�$�*�*R��z}�r��n���}�Ǿ�Cd@�eqH�$�Ri+��&������=+�~��9m)���D��M��d�A��V�w�wۮ� g�\ :��]ޓ�$U��}�����s�/h��7�}vn�7Gwh�1��qw$�YN���ЀA�BQ9�X@���n���V�2Wh��G7P���N��������~�wᏪ|��P�X;e���OQ��{�p�f��"4D��N�zͻ���@DAڍ�	UD&f@����dӉ/R�����l���gv�G"K�:P`^���=|��A*:�(�W^{�ȿ��E�䅽��$=V�]R��лaJ5Dt�.w}sd�4O���/�J�kހ�#�����\����g޳wY�;�E����=��I_<@� B!	D��^��C�Z�B��A��pv��+�+����#�ż����8]؎K̐��`�|:����\qs��r3�g�*�Qu쨻0��G�r"#�9�g�9�P\WWK�o��.E��.���v�4��N�|����1�թ>�}���G�+���HΕ<��T�1�(� p\����QPf5���rO���7l�4}��|=��j|�D��,��m�"E�ut�#uLj)�R��QJ㍴ �,��Bz��щ��DH*(�d����\�Lb�d�R�I�`�rR��GY<S2�XJ;4\]5u���dˑ��x��f�rbO�� BA ��L�C1 �r4$)$\�k33!'�D\���Zٚ�����S ŊD㟑�V�㗫����s�OC�
3w�T�3����٘H�w��҆�m��,>��7���o�����	ü�4�M|9�rFE��9�P�ϣ"��>����������#��D����J����,�)r�˶����7H��Kls���F���}p|�ݣ�=)�HD�Lw�	�9/�_���77Y�{��r�gX}"�O�� B!�`��}�:�E���Ƃb ��Đz;��'�k����&���I�4�!���4��E|w���%�~�@�N��Ng���Ei~%v�W>i����Nhl�>��R����/�G�Ǽ�cЏqns��? �G��SH��m�# �/~&~8�Vb������/�%�7�2%�诣�2c5ą�.d�I�EQh������f���3>�l��f��-'�QRJ2a)�ʵ?$�������Ǎ!�Bj�e�4�v"��U>�������ǉ_�G�����ag���RL�JXd��s"o�VOxe�.@ ��~��azd�U�F I3+s�&2�,�/5ϵ<|��xd�{C���_�(����.mG���ޅWk4_�U+�;I\�G��i�2�A|/��fd��Bx3J��z���!�?��7Zvg�AtPo��0�FH�L�O^���t�:VD�*O�C��>�Ϭ��f��-'���?��3���B!�Hcyߗ���IN�*�oƆ.��d�+��__�J �͂)�F�am��2HQ#CfԱ�fE�H�\b�6brjQ%O(��+;��7��e�����|���mLL�����a�|�8��H��h^�KeW�溡%JXJ����Cb](H8m�e���BG�$���UA�ƲO���oZ��J~����zB�RӸS��8ޓ�p�����tVO�4�,��札)d6���w.Co�o�x66_Y���O!�)8p�Çx:(����7ѿñ��E���v;����}��ǃ�-��p�>�vc��<γ��9^q8�]����w�ҭ���N�����L�L�K'��Jcq�p�7CO�~)���]�wm��ln�wxk~�{N�ڝ�668p�L���EOR�c�#�X�&��䀗\c�-Vc��͉���*=hhZ��NH�^AE�2��נ�Ҥ�B`��TDyd$�aL�a�k:B�D��Ơ�"u�D>Y
F0�x�p��dB�1��@��	q6�
����uz�3K!R79q���E��AD(x*2���t����X���"1`(< ^�Y`��,h2u�0J�Z�;�Vy�mA�،��0DI6f�^��[i��+(��4��S�ZWq�������� �JC̘*���H�6 I@�0Z  d�`'d�ʛ���#��n(J$TX��`x�pщ@��c�Ah'�#���C@$��0�`�!,����`�BYJ(�{Eı�(��
D����	�w�������F�!��lX�Z�J���E�mbF�����$�<i��`����f�8� ?Zу#�!T��i�Z���Z��dC�Bc�In$B�-��$o%�e��e��Z�pm�ٍ�#d��[v��6�1nCTz�M���Q��;2X�b$�S�q����*Xf�I	��֒
��Ӹ6Di$�yDf\�&�����K�(q�I��N[ac-Qpő�6\r��x��.l�	D��E�����A3�z��.�ϊf�h�,f�1�$�����m��m�c�1�}q�I$�z�v�I��m�i�c�1��$�I�I�I&�m��q�1�c��I$�z�v�H�Ç�.K�.��fٷ����i�W���	��S�a�F]aX�_"�J	𖺰�$B��TmB�Z:܆ȃ� %�ȉ�	DT�a&+a	�O	
P,�M`DT�_$.rF�a�L�G� �@� B��)n��wI�!�C<��r��b	u�~��4x~VNX]���J~�����oy���b�i섁,4(8Yr�3��{?}��(��wc�ǃa<�#岯d��fEr(�␑�:�܎hPz8Y��°�>�4���������ɔ�멹�DL�Y�4�mZ�4��f���M�!Iw,p9O8e���E��jAWO��-j����>�G��l�6�Y�<�E�����&F&��B!(�ӆiQ���+��Ot+�$D7�89˸Q���Q8רŇǃa�Cz�%$�s����>�Ҵ���(]s~��J��}i�� �����ĕ=�
И���'�ȇ9��}�f~Z���!d�e��0��@��B�cGO��F��r�?h��Az���(�)���%r::+\��UyG����Eć�p�_��h�Gu'G��gۅ�t|���>���p�'ǈ@� BI0J����m^��Ӵ)C�b��rg����u[��C3۵Q^�Ǵv�{�2
���Ǘn�z�/�5B`ʴ-?6���Qz՗�q,�R�|�����=���]o�-��Jz�e�߫<��zEQ4��>$��7�?�*o]��)w��4z��~>�-�H9�k��#F�w�rQ��$ @�l��P�'� T3�a�>=��>ȺEIۣ�}g�gۇ�Y�;�Eɽi5�5��>ㆾ6h�@� I$�:G
뭙D�t�κM4T��g��<d8=�c���BN�.��M�da�8�d ��o߉@9�^���P��yo�z��G�ӆ�SG���?U�q>��}$�dp>=�H�.�I��EN�O��,/��y�"�$+��9Aa�2}3����,�G��GmX.����g0�@�b��m1d(�;�mf}f�z���b.O1}X\�=�j&���$X�l\l9Q��R�)�t��J�l��6�eam��2U-T�i���a2ir�(p��n�d�UL��Z�ʖ�+v5�B�x0.��l���$�� �N(�*�� B!	Dֻ6�x�~�ޥ�6�2q���!W���1_-�D��gCL�}�v�㧿$���ov6e�Y5��<~�x3�5O�r++*�j��l7���y<����U�[fM]�;�@|o�Pe'�x:�3���bFG*�x,M��+�U/�$S��;g���e)s.��$�K�T�+]�A���%�:���6A�ϕ���!�H�=�G�?��p��n��z����Y����_��@� B!	D��W��u�{��y�	�F�������Y�����n�!	-A����Y�b �(f��K'��x�U_(^��M�M���gd0�)�W���a�lӁ��o's
�OT���$8L2Q_��� #�M'#* *.$���p����*
���(_GYEɅã�,/��P���`�'Q��ɮ�n.���l�JRD״3Q� #�8�I�Q�>�v��6�����\����7�o�ݦ�:@� B!	D�{��vy����2�~�����垮�2I'�b�w}L*�A����w�7Y�r�˶�$�TG�E�dD�Eh��Tl6�V��p|����⣣��Bq�5���z@U՝L���HRt(>>�Q�Z~����A���f&$Kmn*Ae���nϪ�֒�#�C��"�������H�]��f�Id(R�{3��T�Ĺ
a"&#e�aFl��HF��
��"�&Y���q�و.7�P�$C`��R$�s��*Vj$&a%M�N �1&bj��\PE�`����bB�@�#�D�&�*8� � �F-�̖�ِ�u�,Yq���|�<lQq��h�K�*���@d dq$A��� �Ԝ)��H8�aI"p"S��i���A(-���=~9|��u�8��cR�淡gc4�=,G;�b�*NmE�>���vٺ;Χa�������V bV%��Q�"�'2o���7�8�!X�W� P�4Y�&�[Zm��EZ!���IF5Ah[�B��(QmD-�+�@U��qܼ��Սi�3^8a�@�%�̠����Q��;�$w"=]Ϥ�x�f诏�O����Ʈ�.�J"M$��zk
alD��֋�ĲC���*�L4y�G{�����YhH�H����¾G�����������>�o��� /�L�i|�KS�Q��w�p<#�a�����ǟ�8�v+� G�Ax�g�,��aW��{B<.2�9�rN������>�7m����d��d$%ڔ�SIo��Z��x�P�%ۓr��z�4�,	���J��n#`Q;l$�UnG�AQY$)D��5��@U�a�v7&^+be")2c�0/�������1L,�eݬ�� B!��lޛ��K�-nD�2e�Y���� x־k�U��q��#q��U����?�"=(.5P q\n	K��U�Gg����|����U�/���3���/���'��uQ������/�c�EB繼�p>��D&��xf�?���0���6uQ�=	��Gg��>���~��.D�>�lh3��BK ���Ǹ��̣hof�����b2On����]��/N���B!�M����v�Tk���j�or���������s<G��֡Lė\�qY��0�I$� ]B>a��PT^���{))�-˻���h� ��|�5��#m�Y&e�mŹb�+c+�p��xƍ���k�� �}�H�!R���oƣ{��] ރ����feJR`p�d�]��G�||W�|{���y;�6�6��ܸm�����}gY�e(p��8p���#����7ѿ�X�xX��k,T����U�[w|��wNCtq���ol�:�3��O���[��_U���iV�z�I��,�<�ޕL�K'��Jcq�pӑ������7|.��[�����x66_Y��ܝ�([?���K|�5e���J�V,��w�r
fB���~�N%u:���2).1i�y������h)�HP�S�2C�x�s�=�6ם�Umi1,|��VЯ4��~By;}H�F��ե-~@-붌ԣ��ָ��P��+�V����%θ��i)�)C�D�o
w�� �KQ��DR�<� ��U*e��t�����2e�:ih��\*�%W�S�YW�WP��]M4|�C�Km~t��)��\���{��*�ZE�$���1����I$�O�:I$�m��p�1�c�i$�I�'I$�m��N�1�cc�$�I>��$�m��i��1�c�"I$c,c$c�p�Ç��]�t_�6��7m����d�u�}]�oWW���6p�@� B�Fs|��?�v�~�q���`��>��.W?�w_V�[��F���T���r�����_0<t�_�s�p�.�O�l0�rcV�]-Da���)�L@�P��2�L�?��}=���:j}9��YpI(e�d艗g�i��t�����8<-|������*��Vk�J�eM}S�V63;8]�r�]�d�.a�nR���+�ߡ���G;� ��`�i�>Q�=����pݶn�����Q3! �]U]�M�������!�J'��;ҙ�D�P��Ux����y}:����k���_��H���3�ԙ��RHG3�y�!��~��.K�{ʉ��0���W�U��'�`�*6"	�>��#A��lȃBNIpiw��A��yI*|*��R$RW�MN���8y�����q���N�/0��3��,��a�O�Rs�m�;>�7m����g�}�']y�5u*�{HR�*	�4Y�~kS��t�2Y��aԕ�D#R2�l@x��1V5ҸA�Q��(PH�P%X�!ײA3�
����	�(����"Fc�eSi�C[v#r���B!�lލ�����DF���`�$�܍��Zlm�N�]r�ra!R���BQn:r
d���wQ�1�8Xy{�`��H�O�xL/��>���>���`g��d}��0�\˪����S=�u,��XR�F��.47��8���S+�d�n�ɌH��?~~U��M������ܺQ�~��p���!IHs�M���vG�.���7pݶn�����|���b��X�	$�@�%��N��	n���Ua���>��>���al�̔e�Z����0��D��p�8��C�2������_i��*��7�w.�ad��-�/gSY�e�Y"e݈��1r
FD�ql֡$�����D�x+���9̚��&(�+���3 � �x4O���;_�$� 0ĳm:��2Ŋ6�K�����F�<�'�� ���s�T�K,�7�9\�!A�7��P���Wy�+P����\WR��qx��{FQ��Y���n��������\���HB!��[j��Շ�x8j��j�<����%@i����Nl#`���l�7��YE��IXbY�y�d��a��0�%��$%��$`O>��6҃d&������a?r>*�9���K�\;��u��|_��h������ӂ�3#�dx-��g��TL���=Fp���w�^��1>^�9�Qؽ�d�q\��&>�^kW�����@�%�=��3�r��3�Ь��V�=��EuVo#����:͡^���bb$�O0�ٍ>W"k����}]��F�Q?j�^�AA��ߢ}O匣{(<�_�(��@�>_���������{��I9�G=�|�l;��ۢL�|@������p���H���K�i��W��Pa�hHOI
�gQ�(�n���7Y{���g���~}|;R�L�T�ʚ1��rzD�ăf>B�@��H%	��Q�K2�*�S��дW1�1�d&˼�^e̋eܴ���. "��k*$�[,L-�R��H�IR��%��|@� B!	F���Iml��ԩ�)ԎI�Ļ�Lʯ�;Z>su�SMo�ty�U٥U%Q�m�pp*2U��$#���w��$�>��G��_A6J�gi���C�}Uj��E�;:I²\� ��/��B�;q����#�+�tL̒v{��.E�p;�@ˌ��j�=�6LXTd��L�J0�y�L�"���Pt,/j	<yAq��$r9ϰ�1uH\U��^�tn?��u���#=D�]�z�$�!$�I!$�`$T(�vຨ��ɻ�d�;��w��G��=�\Zq��ޕ~��3�B����iV�Gy��Pv;��þ�����cG}��#����Ƒ�s�ާ�a��+$_�Y���]��E.�.�jsqQcJ�0�p\N���4���^HI}�U��w��`;��gޑ�ʙ�:x9�I){*h�3(�����7Y���b2MɭM֟\���ǋ B!���y�+�g\�2D��~obM3���m�t�����E�A�Ye��u;\���Hq ��XŘî3�Ϧ��)*����}�0f�&�P��w��������a�n���d��6J����*�
8\X�і��eK�4����n%��(�0�k���I寔a����O��1�bZ=�Q�>߼3w�{tw���c����J)��I2ΐ!�BQϸ2��-$!F���<��p�|Tf�GǦWǣ�����`@�m�Z뀉ĩ���B��44��|^PT+`��Q�]	\��y�x��0F
3_&wd }�ֽ6���C���1G �y�a���2�%APeWp�	e��8���t�N����Ջޯ��[U}X�=�y<���C�p����C|�ѻ�̱���c����b��g�:��m^��k�W�4�յ��:��{7779L�c�T���ˆ��������ٝ���gH�K%3���Ç�7CC\�M���}.���u�����ݏ��u�gjwccc�����/�7�z}����#dzWD2����Ʉ2���lP��2���F�C0�hY�bO�=ΚlX�$f�N���S'�ޯ�i�MLw03�A�"K���j�;u�!a:b3��y��3QoqZF�l�[U2����q2
̧��nn�C`���@��9m�,�J$NM�a6��1S����c�-s��{�gH`��XE��@D$��~�sSm��y�q_4F���4$��I���6�p�����l4dI����|��Gُ�9��%ܜH��<'�9Gq��fL��y�Hj��4%��_Lb?I�(Z�%��/��X�C`�Y/�`u�*����`� m�HI�`��j���1��[$"Q6H��2偷�C���Dd�U�Ϥ��
�4���)J�&�`��(��Af51� dTD_%�U&�`i�h���)���ئ�M*&?�YL�U"qB�A�D�20ь?��^E2�\!�leݨIc�Ù��W��L�$i�!-�b�qSA�h�J[m� �`������ !y�����̛��-�"IL�r����L�X��&��Kd���dY$�m�&����H��֠��مAj&B"2H_�M�1b�\g�A�C���
Al�Z+�(�qBS!3í���co����'�q���$�I�'I$�m��N�1�cqI$�I$�m��N�1�cqI$�I$�m��N�1�cqI$�I$�m��s�E�.����|3w�{tw����*�_�D$2�q���*��c��,�b.TfU�1W-�8��.g��&s*��
��P;���+@D9'J���	"�r5e.���͐!�BQ�{sv\�Wc.KnL�2I�v��B�����7��N6���~޹N�Gt[	G~�������'��װ\��z��..*���<v7 �>#��o!�
���x���(����vO�����A���9+2{?\Lu7W�%�W�9��]�C̔����i#���E�G�k���u�z;�F]c����8f5}LO�%�h�����Y0�8{���6��TW8M��$�A�َ�x9�$�]\b�2���h�Q*���J4��wW?M���$�V���Go9��*�������*��@��aW	����A�����/��~Ӟ�=&IG���[��o5�[�4v)��������=
���h|1��������F�w�=<�	� B�̚�{�����nE�{G�3��p<|�7�lOs�����O�B{��1�1*�p#U��UU��r�F�D�0.1�r�f
,.0Y�*�x�a��z�n��Ɋ�C{NԇB�tس7þ�;Ԑ�;'�����n��gp��
JJf�*B~��aY˩��g�o%�ܻ	~�-�1��g�q�%(�B�w��֎�#"����|n���7�>w��Y��%(�:�뻨?|`� �#F��w��ڰ��kxľ�����P��t����7��3�_��S rʈ�D؄�Z���#���888a�B4����>��}�u��^�p��P������o����q�:�b�K�Ɲ�fQ�#�6��i>7�R�B�֫�6�Az��4�ۣ�~�����D�L�,�!�;�s�z�����p�f�Gy�ˣJ��ʓ��Y*�*JHԍ�
�$�l�	��H^��e�8Ԓ4�!FP(@A���~]剑RD$���Q��K�'A����+�Z �E�sVL�e�%��ޮ��Ђ �#Eˣ+w/1�QK��ċ�1�����v��5��H�]?�
�Q�#!�HC}��É�}ߠ� ��c}"3�Au�r�w��,?k䈪��L�+����X�R2B���ӛ���xj>$�ӟnr,�Z=	AQ�9��{������E�;ݧ.���'�,|�`���`�&��x2��}���+Y�xeN�r�&eC�����7�o�w���<��>�=~�o'�"R �gBW{����U������P(�X\J;��<%�oђ.��]��e�hK�����
���U�ͳ}'zf}�I��I�zw�q���T$�C���^:zB|��dɅ��"�̄n	��������;� ���s#�m'���0r��}���F;��	�@#�0�tv�����M�u���#.����'��AF���|!�?	��L�CT�m�	X���}�,�n��،2)�B��|����h�/x;�{�A���P�P�Yf�$�p@D�K:�Q?M����h�(�6]`wC�}�� �*�(Z)Gn�5���R�Y*X�r����rˑ��2�l���E3�����wW�z�]�j[���~O��)=W?3*�Y�4Lz���
�#��(&Q^�ќ>������7�;�F]�T����*��DA���5oW��m_��7��W�t<�r.�n�ӯ$�d;����qYr�$r�߿3����+��� ���b&c�
�<���u�>�v�܌fQ�ٺ��S�C�	g�Gp�h�v

��őn6~���Q�>����V�f���c�ި��iqޢ��Q�/��p�f�Gy�ˣ�,,��L�t���L�ő���>�V-D����-$�i���A�	<I��"�b����� Ԑ�[��dU���Q�I��8��
��3��T22ADM@y�>(ݜ��"j�0��,�w2e��\-�A��s���R�n��lK��!.�K�G ���<�����F~;3=��R�0���T.���~FB��f����23�P���tR�on����r�.eB��]���L:}pO
�B5�jP��I8�v�����:�E��`i�,����
d��B�<������gAd��eۅ�(����k��8�NE��S�4���*�^�&8�Fz�������L7Y���b2�N����v�B1!d�K���z(�v�R�T��K2;�,������/��pN O��gyF�]��[tkO�կ��Q�۠�v8v�GP�7�L%ߤy�_�.Q�����(t��b]��+�4T�;�(��ݼJ�o=1£���u
f$IB���z��&_ekd��?5��bjH@�(���}AY!�.<X��<.���sNsO^���ϓ�*�Ub���]*�_U��e��gj\8p�Ŷ�t:��[x����}X�bŅ�*<�_e�#|n��ܸ~Ct6�47�l���8��ʗ�[r?���.+J���c�S=���o��;�N��2S�1'�ˡ������˾�m��:ln웻�v�x6c/��;R��5t������ݛޕB�M+�(�͙|�g�p�!�&��D�����=�ws=lWv�v2w|�����#=�'�r�s=��Տ{��1xE7�¨��0���i߈�ܹ���=�g�=��ﹴs;��H�3Mbbq�I$�bi$�m��i�4�1�cq�I$�H�I��m�8�c�1�8�$�I$I$�m��q�1�c�p�I$�`�1��Ç�.�/����f���h�1tV��g9��-��F���=�2h����h��������{��4$p�an��R&T��#��%��WϠб���0SK�#!������^#0h�~���l~Ϗ��ϗ�H�U0%g��������0�N���Q���Ma�?"��CW����ҳ�jM���j�	Y�8�T���O���<��������Ǧ�kOs�N�˾���r��yC���S�C�t�(r��t�×��o��q�[�vJj�>B`l��aNG)Mr�SZ&N�(���`Q� ]Q�aGLT¸��J��e�r���C����(E�W��$����{�w��	�a��:j`?�S�+���B>p>u���tm���]�Mc�����wXaޏ�J�X���aO�����D��\b�,|hZؑ��jp2�U#)�K5E�aj��v���>�R�DrSL�aM8�j��n<el���j|+"ܧ�%��ؚ!d�ɆY MvD�#���Se�Xf��!�֢}��0��e�m�e�6�x����k�����NH"��Z���F�����B�N��BB��xbA_Y�v2;�r�w��5=A���	�5k�7��Q�+��>����b":����6�B��\n�lW�o=�R�hǺ�!�:�����f�p1j/!u�:=�7|k���8�1t+���fy�&����!Q��L�D�fs��ӆ�W�΢$�/�}��e�YWF�dd�,�W�������G��EaĢT*��� �2��8 �)�b� �&YA��� �!vH.7�hU	�5#1˂�䰲��i��9߮1���,�Y���!߳����r��qDiߢ�="<�3�uG�W̜Lq5+/Y��� &j���i4[:\�2C�;;h��5dw+ޮQ57��υ��%7��/ ����`C�R+�z�������r�~�,�s���1��"""7��H|��w=)�D"Q"*�`���A+/���ҡT�2����]Y/�y����b@Ĩ(��@�[-�G���"k>>	�=}�ɔg��6�W�Ш����!1giy�Lȃzv�G�-_l5�(��4���O��$0��8��Ѵ_���c�Y�>��F9ny�ݼ���!B���dUs&a�)�32K�;ttw}���6@�|O=�����ԑp������M�h���2ba��xR��9�/;��\Zs0n0����=���������,g�v����\���f$P}�ӨÜA�xP��'��Iϻ��{�Ǿe�=����^���Sp��A�HB��v�\����]����ӺF��ԧܫTʑ5�"K!�⁵x�
-b.(�*�W�l��Q�&�Y~��Zuszrl���""��)n�A�r� oWc-0W`a�f�0��1qU)B�* �FЈ��"ìA�<�Y+&U˓��""#x;f�m��$18�2(�IJ8���o,��M���W�Q�,��?^VM'���f�!�J��NdD����2�<l�8$%�
�xIq���<<����i��6z�s�~ӯ`�]�3�&��g�uJUQ+�U ���ќs�r�~?�gP�!B������6����cz3sNe��Co:�N�k�i��!	ʅ�c*�+�=�,<�����% �$����BK&�t��s��g�CLk\�k��^RD���Q�'Ls!`�{�hH�,s��7�Ux㭂�;7�,������H�K�� a2Jb@Y��������	�gym����&��Q.�����4aNwߛ��<���i.�®�Eut]�3|k��4�Ҳ�~�KǤ���_!�B�!3��
�ނŜJ�(�r"x��ˮ��#�)D���28*	�u�?��%{憏�I���P(e��l��Q�ǖYtw��IZ������3#d�i�m\���0���
���I@�����c:F���Ct�U(Ô�ZLR\�u�'8���,h�Qھ��FQ|1�;�M�+-���z��9{��I��DDG��~������)W;��@��	8;�|�f�T���ی�E>%�Zd[Nj5i:8Z��1�ճ��:�o*�ʊ/�qp{�0�:�l�P�&{����뚣������̒a�7:3�J&�G*�;D��ò�:�F�v��K}�����g�<҆(�������  W>���G��������Ѣ:�a������ɸ[�����÷&�l�p)��
�o�㡀�2L��L퉂L��0Ĺ30L�3332�D��0DT3�3,E,D�H�́�1D�PL�D�33AS�1PD��D�3�3�4QF�u H�$�"f �� ���@��f�� ��&��@��f�	�� ��"	� �`�&		�`�� ��(�)�$	&
� 	(�")��� ���"
�$����� &�����*h�(��"�H���)X�h�(��eb$����a�@1*���IY�*$�j ��"I�f&	�Bfb 	*�����Vj��j�*�f��J
Jj�V
��$� �*J)*�*��%]�d�T�T�S+U!UIE%T��U5T�+SUIUMT�U%U%�+U5T�RT�IUCT��ԭIT�M%�+RURUU�IT�RSCP�r����J��Z����J��Z����j�	X�������V)*�(����(���J%d���h�(������* �i)��b��$�Hr�HXFP��!aX��!dHXa�W��!dXT��!a!aHX�!\VV��	$,�,�B��;f�F�( �VB�hC���adXHY@����!d!�+�B���B��,,,,)# C��
B�������,�) B��Ȑ�
��,�,� B��,� B��
�$,+����,�B���,�(@�!B�B�0��,B�,��,�,�������,� �B��$,)
B�0��.(��0�, @�*C �����0�,!�)�0�����0�����&� YVBRBR�`�`�`���� �FRR�p%H$$!H H$%$X%aH  �`�`�`� �`�`�`�!FF	V	F ��@ �aV	 �E��T�E�@� ���dH!$ B		H!$ F��T�@�A���D�P�XF`��VB	%aB		!H$`��@�V%a�l� P�@���BJA#,JA�B�,�B�A,��,0B�,�@�A��A,0J�(A+0KΈ����`�
�	��$�h($���H((&�d���H(($� �(F$���H(($� �FX& ��(($� �V��H((&	 ��\�L��H(!�� �

�
	� �
	�($�h($�`�
f`�a�d�`�d�i�bd�bd�d�&�&&I�d��&�&&I�A�a�d��&�f�i�i�i��I��&�f�&&�	�f�d�a�i�b��&�i��I��i�&&I�I��I�Y�d��f!�i��!�I�ff�d&�fi��d�fBfH`��fb&fHi��fd��&&if&i�b&�f�&�f!�\��Jd�d��&fd����&a�a� Zfbi�i��I�a��hfU�$"����fA���ffA�a�a��f�fd�&fHfd��d�$!�CZ�H310CC3���L�0ʲL�3���2C0�ăL3C3�40���3,�@̃1LB�0��&Be�do�8�HI�!$��J�HD̄��C$��JEL��I3 II��$� IL���$M%	�%(N�n�XaՃ�^��	���pNC��z��  H$R�HAUJF5"��p�����<��=�v�}_w8�{��=�^l��_��i�����)��730�<R�Fݢ�T��\aeQ����#nƶ����)�/m��5�Y31�4W���7�m����q��ѹ� �}���޷����8'�пg���""~���?EUE� �D��9G�?����'��!�p�L������t��{�y�g�����x���(����G�|p��� ��q0<9WC��'��Ӏ���9Q�d�L�:t���bbJr|��=0��瞇T8:{����1��?Ѿ�t�7cQ3/���pw�F&�"�m�(� "�Ў
.b� *��P��(��4�m .0�;�p�F��b���3�Z��<�C6���>'�v��@�b (bAUNT1fA2T2� �!E ����pH�<������aǠ���<��|��6��;���1�����p}A�G����W��!� q=��ܮ8��>tlz�c����G�rdn��F$ߒ�Aܩ��<!�`{Q�yI/��������J��a��|y>��~�UT_<偺���`��;����Ǳ��v� =���&	��>\b���GҊ���C�?�W�ǃ�M��)���}c����Н�=&�X��@QwtsȂ�z����l,=D��$\P��@|8�t���� ��#Cq��0d���a�xP�&�sÏ�:�A��>Ǖw�	ъ�:	�E \^�}'��^~H���UQ|�_Y�?��`�d�|�^�:ߓ���6��Mc�5�JE�m<c��+wjx�I�y6�����D�����I��{S��6� 	&��菄H!_�����}誨���}���3;]Q��rj��oFs�lGV��88r�$������ �5<l7<�0,��a�T;��6���R�	�LQwGͲ6oF)y�0K�ݧi�I$����w�!|�jĜ�֞' ���`��5�u&dϧQ���1���Rw)�<	����~��NA}>��$"?2T��^x�H���>?^I�u���DD��v\����1x>~8�0/Xs�m��?y�Δ�� � `^Ǡ�z��?Qw$S�	2�p