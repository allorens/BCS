BZh91AY&SY�c�8��_�@qc����� ����bF��      }�GѥQkF��T���+T�+L��٤*����
Yh���ٕH��H���l���R"��U+fkJ��ƚ�J��䫘UZ�n�,�f��Z�ڬU�ɲ��[ҳ3�#m�cF4��@�f��l��2�S0�kKZ�f*1�ʵj*Z6���4����|������)U����[m��U��l�5fըC
�QY�5�kJ͚j�3UZ�Zڒm�&�2���e����2�U4�kU�D���ݩV��%Z֟x  ���$� �U4z  0��  ����ݔAK�qӄ9�֪t�cT�W@�ꆃ>��V��Yj�6�)�J�m���  ;�����^�r��S����@��=�(᎔:���u��ݼ�{��E;ާ��l�ׇ{���K�Y�� @�g^}*�D��j��6��jmV�<    ��>��N�G�/8z
���i����7���Ϡt ��aϾ<>����-����U����O�z� }�Ϗ7�J
6��R�����o!��==7e��YZ��m��խ���Q����  �>��ל:=R����� �;��+{t�u��;oJU0��:Sw�]����g{n�42齴w{W�(*��0A���w�f�miZ٢ҥ��mkZp  �����ݶԻ���t{����M 4w/nJU�����T�^i1�m�Q�x�=m�@{���z��s��Nz�;ޫ���>�>�4i��m4mDBT-�ָ  <(�>�x����ж�Q��v�WM���ҕER�ޠ=)飺�S�uA�z��zU.:8�A��^�*�v�8��+�T>�e��-�d�#e��ǀ ��-����T =�n@���=�OJ���C��Ü;����`QB��� (6�n@��q� �U=��i!cm��6�ZN  �(�l� 1�pQL�X ��AA;�� >�{o  \p���uA�'{8ր��Ͱ��[Sem�j�1���� ��Q��
)�u�< 
v8 �,��z
=�P f��(n�q� 7���� ;ʘ��jZ��l�V����T�� g�*���4 2�A� �&Z� *�L�c�>� R�y�� �g*���9B��         �*J� 0�  �� T�aJQT�@ `� �)��	J�~�      �%J�      ����������    ��کT��S���@b4�M=����;�~�(�������+𼫨�Ǚ�f��e����|}�?G��ϯ%DW�EDYEO�D@U�o�?y�_��a��H�a����C����?i�O�EX?�UU��� ��=	:B�>�DD����������ş� ?��� �{���L�������YG� u�:ʟ#��(��z�=e>�X�#�Q�*|��XG��u�8��� ��zd�X�:�=aN��� ��:ʝd�Y��ʝaN�&`�
u�z��eN�XW�#���z��� :�=a��XG���Q����� �����(��z�=dO�^�/XW����d^�XG��U�"��zLa��YG����z��a����
��z��d�Q�(��3�A�(��z0��z�=a����֘G�z��e��XG�����=d:�9�z�YG������zʝa���X�����z�=d��X�W������=eN�YG�#��g���:�Y�#�ʽa�/Y8�=e^��YS�#�A���~���s��zʝ`^�YG�#�A� ��e�S�#�Q�
u�z�=eC���T�"z�X2�YS�)�Q� ��z`�Y�z�9�:�=aN��YS�a��Y�!��u�zʜ`�����z�=e^���=e��Y�+�ʽd^��E�o�P:�'YW����(���Y�+�U�"���e�/YW� u��/���z�=ax���z�=e��YG�#�Q�`^�u�zʽ`^��Y���U� ��� :�W��u�������U��e���YP^2 �`z¢���"��PW�(�Y^���eW�@��.`z�
��:� `Tz�*��D:� dz�!�e\�XG�#�A���z�=e��XOXS� fQ:Ƚa�/XG��Q�
��~��
��x��`^�!����z�=�����k�)�Y����C�Ȫ��MK.҄��k7
�.�f��'mް�.����K6�չ��,{�h��{�v���tV�͚<�B�ͷoe�k���W	�V�+K/q�*��kcowS�4�OH;{�/J{B�,��nKe��	� �WS2�a��͙WY�3$�҈ �:�^�I�QQ�4�TqE-�&��ʳBHՌ9T2NXZX��o�i��6��k��Y�+1L���X��U�Nf�b�1�ܡw��%�YMV&��m�!n�J����t
{&J�:����LȃH���
9��.'��Ŧ^iBQ�զ]� w�%��:���e�+RPf"eat	��%D�7��SjV�Twi��S��S�^P]*Zk0�,T��g(`W2���s(��#[4,�I�j�PL�0����f=���7�qM�D���SKYӐ���F�B�(b����ZhRF�m���-k��d�هsi8���*��-�Yn���ޣy�Fq�t�����VӰ��-�n�-c+sY�.�0^�
�o��EeB���4�m���krjgpR��^Ӂ%�rn�.��C@��Z�ijt��gj���T�%O+�7"4t]��R�b:��i��&�d���a�6e�W�:W�k�x���f���H�7�����[ ��U�b�U��ư}J
f���4����[C*d���/�YZ����E��]������F3I���%I!N�!��v��'g�]k�nh�w&	��N���	@b�u�����3qY��9W�ҁ%#2������Y���wV�f7EɁ�K*�յ�5\�,�Q�S�x�wcu���6ܶhT
���3p�#]����oNJr]�&#�-�z6*Ժ�"��[E�X2]nC��z�h<�F�2��Uf��鷱æU֩�hec�5�;��t�N�P���j�fnSfZp#��,l�Ԗ ���{@���N`�&����1�m]ރͫ�q�,ǣ���cZ�[��(d���Ðf�1Z�5Jd�#t�CC5#��qU�ݡ�Pj�̥W	�a�A��xW��c�3Fmkk^��7�6r�,�����2�<'@[�Y{���S�]�y��qK�Kod,
y�2�QիU�����^��{��r��M���	�X�5@��+\5>D#Wx$`�p�+mG�A`�f�wN��U�X�Pń����䵔q��:7�st�+�os -���^7Z�,GW�s}sh��֥맏�ݼ�F^��GNXɉ��B׊����:�a�[M��k-�u�j�ĺf{N�*�mQ��ZU,�y�1ȋ�uN���D@I���h�,B]�,c�Vn4�mV=��<ze��h�N���n�	��T��	W�i2Y6íU��E�[dI�7������ P��Ɛ;����*e��Պ���jI2�D���kN��F6��۽��%ܭt���QU��u��k;P�b��ܫ"^�]�#xrX�R�Ԯ�[���P)HQ�쎥a[�����
�S���h�B�2��a��];����+[�ɩ-� (0�gU�rܭ�V�Q
^�V�'{��K�p��Ŧؿ���Vl>f����*�һ�<Y#놤������67r茢e�͗�5Z&hh�&�B� �p���O0����7u!��	��Z�?n��0NT�����;i�/r��.�K.뭢��Ŗܺ1�);�z�5���檶�-�k%
��̧)J��a�g_�Qm4���t�˴V-t���Ǻ�ޒ��YV�xUB���ݦ(-̋S���:�XB�I��4�qh�d��JU�U�0V�V�;ˢM��
�/Na���4�!����]8��e�ځxwu�ͳ":>;��W���j�ڂ�&r�Rl�kγI��]���w�� ��g����Ϭ-�r�,�3Pk�F��f�ڇ^@Z�v�'lRu%�@�lZ�ګqޤ���J��.�1��[t2kv��Fmh�AA�J�ڹ�eˉڠ�̽�L1F�PtAjn����k.���H�U��	�6�P ;C]k� ���ȁ�bi����ufk�"Sɂ�K��k$[�ㄢ
!�g�עZ�Pd�F�G sZ80Xř����;0�DD�2۴�sd֪�C�ѩ��ɕ����6TY�fơ0Rv��wsHY�c���yA%y�6۶ %��Y$R��������*�.���	�cj��
��2
8�*'Jk3.z��ffhYF��~f���Y!��--swD�v�KY��� ��U�[�仙a��
�_�*��Zsk4�j�(0]��k^1ׇ����������b���xH�}N�Z�]�*J����&�fa�+7m��2�U��q����c�8�ڧX�[���Mܕi���/&�-�fM��Rbtb�g�j�0�h�Z�u�	�Wu6�n�Nn��`nhU����آ�)݈&!��R���d�p�ڌ2�2���$qF�e[�U�S�9p8��Y�rT1`����L��P˵W��x���x�����UYHMā�QC4<�ø��wEhM3y�bg(F!�ƽ�d��i���J:��c��9��if�7%J��u�,�P݉��A/u!�J*E�N��f����Rׁ�	��f���n�s6�T��f��@�qTWI3�ֱ٭�IZ�J9����.�˷u�Y��,���)4��H95��Aˈf���	�a�l;u�C74���ᩍv��f-��ӌ�-8��)��R��eWa��v�U����[��0�F/N�Y&X�J�anmH4�jW{��{+&�^Q�k3n|gf�N,�&���[�����ùj!o��wZB)�����6/N���qҸ����;�a̬�݂.�֝o+T� ɘ$7�5�h,V�i�ES�d��.ޫvTsr�c��c����KVM�Y�#{R��1��:]�u Z�7X�$*ˍ�ز� �R��)�T�
M�W�L7	��f�r�f�N�p"I���ut��l�aY45x7j{����0d��!b��blJ3�^�&�����a�n駙cL�Yq�i��E��%ۑ^�՘���5�ĔL<RM�+j��5��j�}L�EV�<.]�N*�fM̭{��f�jc�O&�Z��5mfK�0m�[e:ke�D7I��@B�w�JxSWnc�$�7�b:$�L�,�m���r;�F�z.���Wu6�gj�����(!Y}��"���B�LF������[��b���r�,�LX6�(�Z�p��+��WQ��E#��Vu����5f0����ݠH�n��e�V���v�õ�Iy�#��~�՚��7n
��i�e��4F��K8(h؅^}�Y�����Q
����6�,L�E{����TE�G��J�0³F����XKn�k� ����m\ʉ=oQ
���5�9���Q�1�74�F�6l��,,(�(�ש�]Y͙h�Ӎ�LZ�N!V^7��ve���nS:ƫ:E���{�ɪ��	��jB)LŻ"!�+q�	հ[����J�9��%
�~�[#^�&,Ukuk�$Q8�a,��)Pr�mh���<(�
9�J;Re����5G#�Z�1�� �l�b��[�G�!�Wr�h��Q*-p]#9M��X�;��I4«[{���S\ŷ�u�����r�iҀa��ӓM�l�9yv�gK�W5iZ��9xE�zڀ�٢�p5��ʰ%6�a���2�N��0��M��SH�)Xn�$��x��/S9��"�I�������ʆ�T��7z5���"�A�ғ,b�ܺ2��s/5�HEn^P���1����)X�!���0�$Q[pe*�]�FL�9����[�����)Cb�%Z��"�9S��s]��ո4��J
�-�y�Ee��9�:����E%�AS����Bҫ@�W�Ġ�$鬛�P�3rJ�c5c���)B�Y�я�TB�n�@bnIw��U������3�-�$��Ҳ�]0�.�a��t�w3Q�5:�@��Ld�:V-�1Y�L�iX^�*�lG\*�� I���#�[u[�V�v��jGy���I�eM�0[(��k1$����MP�vJZ-6,̄I�Ԡ��ܱV7f8�iYL����锲��:!+l�y�ce�m^VJR��"��X�tY-�ø,n�����u��6�1�f擹�k_��-��q	0Ysɒ�+��!F7���1
Y-�q9W/ט�E#�nš�ͭ̷O���;��V0^j�6��v�奠�<٢��3C�ӻ[m�w�Xhn��^������e�Ǆ�ٲ�eA�w�n3��^O�Z�Ɯz�i+��O�����j�u3Á"�����6�nmh!��{*Ax���2Pp�#��p�a�[��^�u�Y#-�	ے!��tB�����-٢��z��d��|�谚�h2��n�j�m��kn�[�u��$i�o[+)�{���]�1��6����dS@�����;VA*�M$�A�Cl�Vk�;��@d���=���[��(�W�n���5�ŸAZ6��Y�t�8+ku�a��6�үBv���`ͳ��'H�C95mdD�PX��u��VQG-嬬�O����1�����t�3@�x�-�5h)2��3}��V^��rov����0c��r��?d���eǢ���M�Tf�v��1I���2[۩������4`�#lV�bP��Cg-�g��[��1�tkD���Hw1�H�K*��(d7*n�dE�����+ub�Q7D�a� Q�L,u�h���XϳEnF8^ɤ,;���E���h�h�������	��н֕�m�`�L.e�̩q[��D��kCK.e!(�Vl'QT?K���.�=U�[5"7W�Lz�2��#l�I����]E ������h�+^�n�TX�5�(��K�Ch�/l���ti-������a�cU��ѷ��,ZT�Mոe��F"�z:�r�~��osf�7��%�-����>Z�"{bo8�T1_:)���!�����U�7e�N�Sכv�h�pROPkZ�����X�������b��Aܱ�i��ӊ$"/*A$�����a��T�ŕ�[աT����k0��i���+�ad��d����v�ǯwW���he1����g�D-%OGZɃ73[��CN����b��5BÚF��9Z��D���WY���T��4��1���N�^��nI��P�ٺ��c���!"VY0����{,]��u<,��oS�,;�7���Y��R	M�!���%f:ֲ���d��X�Gw��D�nJrB���5q;����q��MO/q�&﯅-80�Q�xJ4���B�q\f��6�Fdb�kM�j��P[�x�7R�A4rZ��y�����MYr�kw`�G0����E�	��%T��U�XO���.V;k�Z�i\���[ٛ&���h�����63x $�̺��dJ�T"�R��h޽"���l���m��8˱�Ǚ)e�G�#�9/\U��M)jhm[:�L�Z0�y�@7m��v�Te��@�nD��~�eK70��u���diT�L� b�.�C3C�6�m,خ��4Tc�IN�;�*b�x0ɠ$�FբT�sm�&��#Nfe�J�2�&ѣ+)�R��l�wCQ�S�iʴ�yOP�c��iT���ܱ��GF�I^:{Or�k�!Y�J6]u�iui�EB[;Yp�x$YŮ�
�����0��O(�o�����f���:�6���e-��M��7�.3�)7K��U��3.m<D��3u��L��F:AD�.��������R`�Y�*:��HfbP��G[Ƀh���Υ�R�|��h���m�-U��FQiuڹ�KE�]���SIY�*�3-Ә@�Re��:�����okI�X�+#`�ģS'���#g|
�zs��r)m�����hG���ѐ!�WYY+"�wZ��L���-�R�P��U�q�N� F��b�/Q��!��F�Qؕ
Z��yI�g7J�C7%j٥���[,�h��&�	H�yxu<���m�n�=���DA�K�<-�,k$�4ԥ�תd�]�o%��f ��e��6v��ͼFK��BLi���{��XfL����Ҡ�O�SB=����)�̵���ZY��ef<��:��͵�V+�e��q�;n�!��	��S+A#7*�Ө���Y�����7����{K�4C���Y�y��+c�`��ҭ��8f���JR{����wt%��kXS+$m����V�T0*Lٷ�<kl�@�T��-�ܦ�ӱw�SD2�����q^�m�#/5*�75Fż9<����Fjc��]��'"������DIx��9Wvf�I�qC�tZ��H�r�*�EQ���h��aO����N�#��q�֍t.I�SA���5CHl�f���6+-�b�#-�����L�XѢ�tj�uH��٠T���١�Վ����7R�f��\{���̧;n��	�ֵf�a=�n5�:;��ò���vV�4հ�f^ԭp��V���f�!e�؍�*������;�|_t�4��vþ�E=�b�W"��ߛ�
@W�f��.�!C�m��+�D;jݙWY��d#���Ű4�H,4^�a��-�YfP�n�@��+�,ŏ����5��)���|�Η.�/J٬k%�3��͛@�@^�����c�q�]����Q @Gn��
-�LC/Oh��� �c1Xi�(Щ��F�z�:�i�B�ʧ��o�.�`���m���p�J-��{�������pM�&�<V$�O���|�F�Hfl��W�V�h-��S����Cƈ�1W/��f�u�f�L�q�[���h�G	�Y�Ǔ6���]t���'>+^#����!i ��9-;H7V�$U*U�)r�����ŋ�W�r3y(vri��D3Q�z����B�c0mɖ/e�p�6�V�(If������,5o�������
��0w����y�ꘆ��RNc����nq/Qn4�9�2�^S�c�sDa�F����wTm��ݶ+N%j�ΓF���/�F�-a��n*c�8$�sI���/(�f+��LO�m��r�ƃ�O{+U�k*����/�6�i���%�;6B��;�ӽ�$�I�}
cźT��2�mAt;8����;���N�"%<�Ψ*93l�1y�9>zh��4��Q�u�N3�V��g��J5X�3�ᗥ��U8٤¢�^�7�_<z��;bF�i��ooX��2�V$�tǱ=BK̝4�W���c�[��L���m���E�ͬ�i��o4�����T�a.J^���̔�nei���}�-G��O�S��wY��멊�MRh"��ݶ71xk�m�=nI���#T%�q��,p.[�B���|1���v�˭�C[qW�����Gm�RP����d@�����+�P����ŤoΘ!��I��u�Ų��5�k93uNN4x���'m�8Gf�8�A����C�@���*�P[��J�����#wo4��>^{���e����3���?.�.ᝳ���]SU2!�5ًCjo%	��]ї�̍B���Q���;�iz_l����vs)�m)S�s3If�	QҿX-J�7۔��蛫m��N�۲�u�@�!jdU]5�����5��=�㐲�ւV���ò>�u�r�#ZF�-�O��d��}�T�$͐; �5e�m�v��H��&gY�Zn��2��)�9y\�+�Ƙf�=�;A���%oP[#n����a�Y�S�ɜ�g]f^ǈ]t�JN��Qfj�t:s��yQ�b&n�+���u��̸#����β��}q����B7��@�Y�L�m�ڲhd��K����9AU�	8ҏ:��`���-<���/nZB�t�8�QT&\��qޚ� �I7U��:�s4en�P]����3���C�J�1]-/2���_[�;�Bm�X��9 w�Hh*�����iBfv��Ei��o����GJJ��ܱd�qY׍�c�W�_!�\ƫh�2X�7�^@+�$cmLz+S5��� SjN]�It��y�	�0���|%ҩKs	{�*��w��i����5���e�M�°��j� �x���Jᒦ���,�0ݘo�1��[q�̽⩭gN���qΧ��#ig+|ީ���"������3��b�S2��Co_,t�3-K�hshKr���;���t�U���o������u�'O�Q���B#W�r_T7Ư��n��Hμ���<�r�R�Ay\a�J<��j|p[W��m�,_F��Qɍ]���.i4"}	��bV�&�Wq�=��0�.��U��3N�n�wݛ��\���ۺ��m>ˆ�,Σ2sf`�5{�pWJ��2liAB����+;i)7��I�0*�(ez�x�(�w��,-�ڛ`e��K-�4-��n�r=����f�����N�p�{�t�������es��� |m-�4O��k:�G�U�*�jƅ��j'���1�&u�� � ��0���[�@��<_@�r�� 敊�Z��S�J��:t���S��1������iKu̕�v�T�Wg������0�r��$s{���_SWv��Q�Y5y͸a�f�:!��f��CZ��X �vU�SH��IöpKk.��_t�7�U�l���o9�	�U��+U!r��Wvm�������Wr�od�om,����Q��+qn�V��^�V�È��ӱS6u�t�D�Kct:�Kz|*�=S;E+[�I���qo3`.]��bƞ9wr=�����\s�n"'ʗS.��::�#P��pH��jm�C�e��
�V,�6�d�#:"u;F��\��=�x*:�^eI}p���k"���Z]jtD�WKR�-�sN$�_]�O�]�=�@���>�=���p��%l�c[[-�Z]N]*��O��T�d�1���Ռ��c
`!Px�麇��slа;�Fvͮb�|�#��Qjb��֛8x���T�ڝ��v�!
Ȭ��.8H��7�&1{��v4%֔�
�C��kl;X7F^*'Z�5OxYW#]g&K�/z黣�k�'�d
�Vf�g5��G�AE��VT�D�VR��b,����Q��;��d5:�Ӣh֪*(m�vX�]��6�T�>�ba�d4��E�4M���&����z���y���'Sk��(%]��n��p��LU�k+R��ݐ�!�h*�+SWv>mj���/J\�;4���#��E,� ��^.h����6[�L�@���Q��lј3b�t����%�V���!Zavn�r<�:VMx���,�P��S�}-����e�L�ǣ�8�g9�V$_���:��/rs��8��<,aRj��z{ٶH�g���s�)�Z�n�ڽWV���C���Vj��9(��s�|�����k�r��F\�إ��0�-g*�����x��q4���Ff�Ka�+t�c�Q�/��d#���v�[��w_Ia��b��P�f2�I-�6�;��R��2���Dl�~�e�j�Sg���^&{5�=���eV���C[Л*�!|��0�yu�%c����z;1���ˬ�I�5Z�D�$uiV�
]�(� J���u$AQ���SV�N�Z�-ۭ�WF����&a�;��� `ZH���L�Έlѡ��,k0�c��O�ۓK3�(��]������;,�zءǦ�]�ӕd���>ֶ�?��n)�5#��]H]��y�p�}�M�4�Y��j�%�5颩�7����iKy&	�Y��y��k2��p.ռU���v>i�UpYٹ�,�V)��7��1M��2�5j�8_a��2v%y��50�˥����`���e��&\Sj�]�UY~R�	ܲ!�a�?b9�mH'^��u���d�uDo>��f�n�gh*Q��(��g����R���i)��j�(a������Ԝ+L��7iT���[��̡�53�핆ބ���2�lIt�/�j��c:\zV�kH3(�겴�7|E�|]��B۔ܼ��sy��3�%�r��ע�����{a"����*�^��kH�W
�|�!+]��z�>�Mk�"Rۏo���Ԝ&\a����Üv�4p�r6�d{��x#L�����sf�m]LY�ȻL{�����e	��A�C����>@��J=�y�6T�W3кi�'�f[���>��\��	��C��������2�ln���=7���l��,TbfJ\��%����":�;h���Nr��h�:m��X�V}�z%�f<C,���$ҹ.�3�۫��~��&��Z#iVV�o�-mkep��);^ی^a���wP�f�oIu��gtS�>�>�4�pܙ �W�D��k��6=�v[@+�`ռ���Emk{� 4'<�VwcN!��ʮN�k���f\
R�B����]pLԓ���f=�{x%�7����|-2tk'k;E���!�6T.݂�[=st��0��r;��� �V��9���'k��giպ0��9!=��ˬ41Hlm���a�$��0�=�y�w�������%1�͊v�4��.9gw�sn��m����Yƣ�i望�X$N��*��c�܋Vdv�)s�7�*"�ǫ�U��^Fs��Ga�"8\���M�Z��G.9\�d�0*}M�Z�V���͖�<<*���ÌE�}Y��!���Վ�xzL1Ъ�ܐ��k w�d6����E��q�:���k�������M�=��bSw1:@,:��5����B�8>���	�o^\Ѵ����Re7h�7ZUB�᭻˻��"��p�$xR�A^�g)Z���Us��F��j�ˇn�M=��EȊ얞�[VۣJ�����C����<r�T��4.!U9����ɣgZx��AHZ#t�a
�la*�������S!��"K�L{�鴣��?H�V��M�Ѐ��;w����V0�v̠:R��J�J���n�M}:Qr��g0zN���t�0��������^����ڇ�UU�P�ڠYϠR��vΤ�/�WMĪġ�sEqڏi��W��a�zN������X�2"�.�u�ڋ�nӱ���f��t̘��h�5۶��v�<�*�ѳH�Y����,�;Y�u��-���1 ��G]�B庋"ѴL����ݼ����%��yW��pE�)էi�������P��j�3�oD�Ql>I2�?�Q�z+��⫻�a=s \c��5�v�Aql���Ho�:�;<�GGMݑa��=�;FF�o�8gw�R�֧MM�Ӭ��m�L��J��[)U��[�:ŇR��-�,��Q��7:Ճ}�hI�I��<t����T���4�F*Q��a���*K��Vse7JGK�a�:�[.�@d��۠���sq�Xop���2!�����ΦU�8��]�^*��0�1����e.�#�Ә�񜷷!������ݰ��x�u|���-9�3�a�}��v`3��o��LZ�u���c���f�U��η�r-�)�o�9��qe}��x�B�z�dm�83j��m�!f	����k3xn�v����C�ތ�/mh���C[|�-ړs�u$����?{f�����c�\&�P��}��_N�g;��+Rd��z�pv(�YY�(�������v�1�]���}S�*	9����wau�������zS�J��Nm�{WIԮ 19#��][B��l���{�c�J՘F��Fc�D{6�&ֱ�*���i�uu��M��*;�P�nnv
�Эm��1�a�����k_�:{��P1���.�*q�y���>�Z��:�\���ɴ=ȩZ�*�^�ӴT��`�"�yrQ���|�5b��=2��l��q�-^X�f��8z|�eZI6b��K;��JyՔ�4U�Zb�37u�ZM�7}W(.��0���UZ�����L�y6�Țpt��F�(k	�Յ�͙u��Rt.�a޽i<�h����!�޴���i�^=���0C��H.�m��olJ+� a���q�%�H�k=��#��,��<쉿H��Z�E���R��y
�ԙ#a������k��\H�e�7R�/6�!5`��[Ԡ�����`��_���P�I7ݔ�q6-���s��Eչ�Z�t��C6�up���R�@�K��쑿�4K��a�78DQ��g9d��&�	%��%���"�s���gW^��c~`��pIXIhf7�|q�,Y�dK�`ݭ؉yGw;���M�o�׊5ӵ%�r�s�2�,�X��/1�x_�.��P,�޽��9��B��ddP���(�HIr�U���v���Z�t�ś��dA��(no��b��cr��3�2�okHz�������]r��G�9�;,M^}��ɀ�ֲ���h{������a�\�kQ�X{��%Ymfɸ����w�����tf�v�&�q�w��W���qݣE��b{��Ԩt$뼇k+��!ۓ@��գ�F��,� �X���K�eVbSxqj���}�x	����!��u��JCp���w.;�g9���Cr�
s0J����na0WNVQ-���M�SL�5/��+3���/�P�n�yB�,Ӥ�d��1m�CC�9̬d_vXT�ohT,.��]�Yz*�i�������WKd��Ojm��:*sG__^�%��d�IK�����B,��oN�J��<���ۧW�F��6z]Z���
[�kL�rW^,L�!�w:�J�t�ͷ�J��h�T���%XhL�7CyG�V��L�&����e퉖�>w�3@���W3�� ;��P�7�J��픥���w,��d®��׍�ZR��'S�s����Δ	�o�X��kp�]=�ix��5G�QJ�5�G���1񘌩��V`���	:�T��� �ۂu�B]��xx�'hK�dݖ��ć\������)0��%�˪@�<6��@�ז�&�v\�Vue�����ʥ�_/2�U���gnM'�v5jQ޷-!�u�ȸ~۩�͘{+�Q7��
��a�M�ԑn�a�Uf6�2ҷ�7P.K�l�M�܁��<���b�2���q*������h�a�but��γ5�Vf!��2Qέ�˭h��-ŶhD����h��q�Y�R�Ό�a��b�,5k'n��st����&�:��%G�/$H�p��6�3Mt�aF�D7�U����s����H;g�zȕq��sN�N�x[�t��mN�lv��i�K|�;ɀ(�� h��G'�f�@�ѕ�3���4�Đ���,F���u�i���J����}�to��Ӧ1R�TU�:�sWD,'�t�8��*8������̱��E����RvX�Y��I�V�rAQHwSpfB�����p����H�rG#�I$�I$�I$�I$�I$�a-�u�dnT�X��������%��/����G�g��PEF�A��X5�t(L=�\�>��$o��nA�&!��<T�h]V#�kH���W��ej	 @�o� k*RT �L_�ܻ����g��.�P	<H���D�I�J~LD��o��P�B�n��ÕwR� Q��T�}ce]����*	S"�!
��>�*0��.GSʣG��Nu$��-<ȗIXh>4@�� �m@�"Qh��L5��8"
���$��zR{t£@S>&�F���V,D�5d�t�(,۔%�TE]>f˂z P�����Ǌ�@)!���I�A��D�6� (� /�YvW��E��(�Q��[ ��o���6W�f֘�����e6n��cr�R����G���*�?3����
 ~�T_����O��i�?�(/�o��������;��U��~|�o�����������������l��A�]0��d��1�19F�)mcv��$���5\�n��
�1��4:��u��m[nt�޲�nLj��]����Ý�������99]�O^Q��ӷݘ�{G.�&��f�ӌ,�؍C�V]e�����f�F�{�r��-@ܮDr�Ou����^���ϩ��}Zwj�<�^��CU�!����vF�A��2^����
Sy��y��%Q�`] �� �Նwc(��~Z�m㽹��#�4�y�U����e�t�eL�����Wci"��6Pޱ`��b�!���mgE\��㸃�M_Z��b��3��4�q�j������sm�ɜ�	J�դf�Qˊ����I�J"޷{Kՙ:
��.�i����yɀ6`ݕy��
�Rp=�3uͷ.̢g ������w㕗�Wطso��MB%�J�����H��ɬ���6�-ݤ�U�W��QDn�&���Ja�Ǎh3T�˥ ��(q]j����g(�]�\;̻/;�ل����a����kV��p
�T)څnz�%L�]x�R
+�i���*��	�X�z�nl	"+�*�u8A��i�^��}eMb�G�KK٦A�nPף��Ѭ픃�F��s7��n���9�'fq�B�R�"uVY��|.nἲM��[_�u�^�L:ιÂ�ǚ�˴�slօ�VWi؃@�φ�Cl�+5�!P�%Ui���m#�.5R��ʝ��)Dki��Lv��v���(�T}Rn��f�Ѯ)5�PU��H�p�'��4`:�w�����cU��z��n��cl�:�9��T�uw;*V��,��+�.�:AD�נּ�б�T7LRL�]fb/��᠝V�A����r��v��+�<\$�}T�����ҙõ*���l�{��lFBh� �O�L[�ԣ$sx�Ut�:�;{KP���{[�F��u�Y	-�rV�0�\�fe�u�������
�y��r��{2�Rnwv��A���ûE�85��f�nSI槐�K����\�6솜J�T��jK/0F�+-\f�4�G�}�r���s��emx���m�K�v�/�gV�:�)�c�������4�Q�앝6pd�����F왱^�&q��<�(�+9;y4ִ/948��m��R� �r�1-�
��k�Lk���j ��C�/x�dW�X��ǳͫ4)k��আ� �;BO{A��X!Q�-m���j7j�!Ok�N�]=�)��4N�j�sF�dUN�v;hJ��ūZA-k�9��XUk�^�&�R�F��[�@r���ۺ���"��XvAD��l�B��CE�c���Ə��hU���j]�y�ch��I�GsٽBt���D�3p��V���aԚ��޵n�����`���������F�i�Y�B�R�s����_�Ps��ěT��fod(V �fək-1X ��ky'̮V7�<���		��5���HsZ�wXyor3����K���Bvj��=J|L�~���[���kҊ�I�p�P�v�6��gS�BW،ۻ�����{JH�T<Uޮ
�kq���Y7'pvv��`|'Bv��Q�,���:�䶂rb"j�0�}�]���o[(�Fhqd�r�Z=�`�V��,��;b�Һ�����u�X���톪�c�Z�ktYU��Ո�ڮ�vk_��&�zMbw�����ܻ�+M1Ek3p
+h	�6��eG< Ǽ�'��Y�*�R�Ec��7��C �&��^�w�}�^����v۱$�rf��p|�#�)eatSM\8S�Nq�k��՗�5W+s�:��
�ӌ߈,�W��JA~=�"pڄO,��DK{*��30�՜̧�4Z�]�KM�Dq��^�����X� �3�1B���e=���
H�k��[x,[�����ep�[���Z���.�/S���o�[ҩ*�cT3�@Ѷ����%�[}������\�Pћ1��6+bN�]���)���͹tcV�q��D��jc!�j�v�E`ܓ��:�k�"�� �*Y������&�zk�h���okbwZx?Y�G�7qZv��t�RCV*����f7��l\]���ҏ�*���:�#-��K5t ��q��FfZǯ�<)��!��;F��l�Tq�P6l�V��_wv�mZW�Q�p^�VyJ!�m�ÆmN�����I�K��j�T�d�X�p�|�;���u�P�LC80 ����d�H��b���w��)��{\J��9P���"�#R���!7B���eE��E]�CH�/�44���'�ma���f�\y�jE��n���(a�BuK�b�]Y{�e���ީ�N%ԥ�����C�Ɍ��ă�)�Sti=��
,Vv-���Ď ŔhҮs"���)�*�X1���J<j�Հ�ͽ趦�z�;+7$2v�9�iM�T�je56a�G���_c�!�[�5��L<�V�蒧��E��_J�zf'�OAf�r��Ӱ�ë4sJ��NN�tf9����"��ag2��S�-'�j��v�4�<E�v����pEΦ��B�sV2�J�7N�����,��C����� �_}Z����N���t����i9Ǫlʝ�������1�g,;31�
���EJ[�1P��ru�ӄN t���nfWWY�"��B�U]�/)&_Au��7��|۬�l�:k d;""rJ�Ž�ZQ�{��N[��.��s��Z��/r����9r��[r�R�ܔD�L�1�����I��Y�.�l计[c:m�أ���*�3�w^�q� ���{ɪ:����vm�s��&��YY��0�T�]�<-Y�Q�b��)ᘅd��Y3�B�g��0v�q��x�5�Ηi�K�ӵI������S���R�F�B�#t2�l̟#����sI��0=�&��o�^��S ��S��)�ˢ�V��'�n;�-C�e-�Ǌ�z��R�N��n\�f	�u��`��q��.����'���l��F�e-��%��&��r�B֎����,;s�FХa�I��*q��h��Gm��+r�P".Y[n^�n��I�F=��+B
4{��8a�Z�ޝ�6i}���E91W�0 k4�4�8ܜ�d�uj�u(tfa��u�Ul�-N��pOca�Y��M��y��Wo�F�e@�[�{����3��,S�y��G���{օ�p9�����a{�Mˎ;J�|zV�ٵ�8�ǐ�$Aĩ\���I�+.�VU��� :!J�aņ�PɝC0���39<dv�굧�S�<�:F��9:\d3�u\��L, ����[_Y�
Ю-m�����H��{xEUY�s��*�=V%v�7A^��[��C����Y����")8�C�)v��ͻ��M\�;\��K�����O�ek9ld6:���'�Fh�-�F�:u���_-��X�pƎ�v0t�ETS/M^C�ꕧd�VKt�	s������_�3��0涊��i�p������^F1K��S`�f�D;����G�\�P]��Bp�,%�QҢa'JiBX���(�eL!�R[�9�S'\VD�/^�H5N���_ZR:��������+wke�5i��HdC�$�Bf[P���.�o�,a�mw*@����F���3���\!ξ�:��% ^�3S��J�r��tD��ҥUG�F�s%�r�u��tN��;.���!�2����5�v��;ǵ���F�-�F�ָH�È�[{{_#K������-��jR�-MHGR�k ���9��`v2R�D�U5��{��0�S=��<�#WWya:3�އd(朐��VZ������v+~Nʎ`G6��.�<5���.���8��n��L�q���M�]tQuV����b�G�5H˝W��y�w˛(jS��A��M���j֦���y��5Ij�4�`��L�MU:"A&ݗw��n�˝˕.Ȫ��t+#���d'�9J..��n���*�$s%e�� �^�so�]�GEܾ�c&X��^���w7����i���Fr��J^C��]�Ѣ��Y!��
�O�����͏{#n�X�\��M���]M&;+���Ø������'Z[!�+��|lK�ew5�X���J��nٜ0'h�$�FГ&6�=���t��f͊���'+��:��,V^����daR�ip�U��a��e��UKL^ڱ(i�
�޵W�c�*p�1�9K�e�/HE��ub��TV�h��g/����a��6��A3��k��2֘�o��̰+���y�3 ���;tnS�(+�ѻ״��a)aI���&N�����u��%'�p_&�+�[ut�{)�$w`�y�L���dl#p�]�v���x,7t�6�
��i��NCbF�y���f[
�%*;k��w=Tԕ�p3Ļ�3�9����E�K=�yx�Igxn�k�j#�ɛ@���pT-i����
��ʑ�w-37�e�bQ���Z��H7�6>=f��
��.f���|�[c%+Fvu��yAN�n�*� �ךb$^Ҭ�}£�y�RY1�$n��Yb�iM<�����wA-�"�������H�[��{V�,��}�`��DRF�%42�m��h)�;`�|����ώh�{�v䃡;z�S�c�s��f�	8�V��6sƖP��+�@c�z�Fl4���5��3#�z���ɷY.֣�P�w"�sb�ӧW���r�cR�kc���׏P!}��:������5��bue&�T�-]wi��M.e>*VNr�d�uFY"�X$��Ol����+a���+�$:�,5�:�b��Q�!��@��\c�u9�.��T{�1���O�渭$��{�vm\�eẙC�N�����dfVO:�!���}L�tt�d�Yk��Ǯ��T�(r��B����H�)�Ck�.�	�]��xV��_"jŠ��Z�j�nU���F�L�j&��CB�6YT�q�Z�$C*7�:�_�7ub�VVd�S9y��&7|.��CHn�eh���GH��	��X�;>�a���n�GBi��r˱�L��4����V�U�5�1[�JR�#����3�G�ZqY<��_,�Xo@p��)�����Mul��5+�jd5�9m6�b.�<��Ҋ�0���I�[��YV�N
y�[�CxVYDh0�v�-PP����֪bD=Y��]nU��s9�y�˫�=��4�:�%ٍ�����aV�-�ۨr���L�TG�E3��i�����@<Y��9VqD'���QM��'�9F�a����{n�=>����B���:�^SV���:hV6�cu�f:�p-����(�,^�k�����-U���U�ֱ����R���O(���OY�K��"�(��5��S������hjg<�t�b�tA]X:Mu*�+|sg^Te�}ȫ\کsbӳk�j�V%s��]P߳{�_h'd¯�q,���M.w���#�l�Ku�+���ɏz��,�X^�Y�E����J:.�c֑�ᣳ-	\s�vfHD�QlT��;hFX�`��8���,	��h�ȫpa�cgNn.���Q�odk_*-%�f@��L�$��Xvؚ��/;�C\���R���t溳f�POQc���a�G1^]MQ4i��[�p�kf-��M%��� U�UJ����{{3}q�eǀ8�a�m��ӳ^nh���S[Fm��4��U�vb��tcV_ڄ92�\*�Tv^k��*������N�u i��moa$V�|+l�x4�7��N�*e��)��̭	3SQk;!8[���no~�����%rӫq:Z8v��ϋ����֜zh^����7x�0��o�3-�kN��n��R�ױ+׬T��m�`wF�f)6U��	�aY�k*d}s-;�<i�B�E3uIB��T#\� �t#�Ș+��֨㽪��4iGI�4�Y����WO_�aJa��Zbݜ�+	�D�s5�Y������B�i�L����T��j���
d��v�Ut8\��ۥttk�v������e��!�:M{3�E�T�f��5>���9=<{�V�]�`�A�R��8�$G@e��<<��׮�f��z��;[h>�n�.Zʝ ��ԩD(��t<F<�լ��\�	1=wZ]��>
�-fN�����*[k49�������a� b(M�Yu�wiܙ:��&��)��Ϭ�۵}��h�4)-�
6Up�r�ƺ1����k��%��]�2$+��lN��� �R����`F�]�P��/t����L��~����`�m�|쪩C�U�9ܷhG�l7�E,��JY��i��$�}��K�]��U"���y��ͺr��@�v�Jn�L�ŠJ���1m�=��t��P�&/k����΍���K�6���P��z	O�Ag�<6.�{2���Y"T6�ֹ9���^]k;)%D��N�_U�j@�/R���ZHfn���`��q�+hz����)�����޻wS=�ɆO���)X���g5�ս5(���}�3dPӸ���V·[ΤjdEш�y���	��Db:%wF,���:L�l�>����'7x�p�4�K�f'�3{ps�i�;W+Β<�Z�UҪ��XCa�ݗZ�U�-uE��r�PO��k�ý���8�,��G�,����r.W�_�+��������������k����������{���_������������}g��������������p�mAV?(N�A/������(�[�ɦ�<�S��~���_�5Rܩ=Ě��7a�c�[vu�4g���蜫��[*�kf�������t��y��i)��l퍫c(����PT.�/1F.]��n^0Fn�	��+n�싩�o@���f���0wFF>�=pi�mty`��x�"�jjZ�����k�J��X�]��yc����9fpyw�Ɖ!���s�(A�L����LtiL���g���B�۬\+8bL�T��u��
f�yP�rZ3U��M�Vʋ��ή��嶦i�扴zj�8˼71J��U��E�fi�7����Q'�����ߘش��[�7M��G�A?�|z�tj+~^Y~B��a��w7}�s�zwض=z�I���T�3G55]�RU��c����f�(�v\��<p	3� p��X3�T�O��G8M�A����)���.�q����c���S6���L���,��tXA�\�p�8'�i�/�㚳"-���m5�tM)�B��o�^gl�em��4K	^t8�������$�
�#�鼽��IM�VjX��u�@��s'T��˾2��RbLm�9Ńnb�ݵƞ�s�jj��=x}��|�pQ�לsv�0d٤����Wyzb���H��m
��&�	��A[�oS89{�|�ޜ���+�2����٧��[�� R	��C	e��DJ�6(���t!P�߀�n�`���a�x�m�=�eAEI�$
	 `��15k4횶5i�PFƢ)���EM��+4iѰ�A��Ө�h���D�m�f*����Q�3SE�`�֢!����#�qR}n'
�"l�F��*�I��Z
c6���Xڶժͭ;i�X�[b��DUZ3�ju��΂�Ŋ�֢'llb5c;>n�J*/��f�|s��ȱcM5V�7
��1V���mEQ����t䖚J �Z�m�h�f�b�5$رAk6�ڦ
��њ��l�C:t�٨������d֋�b~v�4[j$�vն�M���4QYjZ6p_I��Ϫ<�����>zy�����aݶ)n�k(c	>�m@�4F�X�����/m���w��n��:��!���6K�����{�9ŽC�(��R&�T�%/U�l�����^X�l��+�����y�6n9�R{��6慵'�=��"�#�3���$#���h��q����{�7�bw�{�tii޷�~4�O����9DG�z�;n`�Q��v�~:O�k�n���U��Iĵ�f���^�O� �3Ps����%�z�e�Y��"'29�%���~��v�)`����r�c6/}��s�?d�i�n���\�ƫ��:�7��
{�)m�6o�>��`�g�~�~V���5����|sZd;�棵�[��oU��W�F��SR�R �sW��;�ޞ��DA3�3��ʡ�z$���d�Ϧдk�rO����q%'e�7
c���A_�;�ak&�\2G�����=�>�����rn*��3Pio7����}�Y��q������G�����G���kU(�=�Y[3[8�_���U�1Ч:c�.è��C�>�ks9������]���_�g�.x��¤T4�bƂa�����"�i�KI����4�A�	2��_Jm�e��������v�����y���9<�sw{��dm���!l�S ������y�p�倐p}��ʺSs�_��E见�$g�x5�fD:=ʿ�%��/=ӂҽ����=����Y*k��nV�o�G��09+"�-���3>�3���+l�b��×��v�1x�}���Do0^��M��?J��7�|v�晪��4w��{Eg���0����o\M��#h_f����/+��|;�jR�d<�~M;��a|H�b�M���7�O	��|w֝K뜘��v���7#��],�!=�sz�'0FWݙ ^P+>z)�z�{'�2��q�<{j�z�t�&MA&�>�챹�x�����f��
����o+�ٰ�Oq�k7�d�F�7A4ɟMS��P|7�C���y��I]��x5��Y�w���vT�進I�����yG'EF�Wo��'�%�=����]���6nP��&ɐ�f흽7|r>RVN���}@�/#�¢�UZ)����cMY.]PX��J�lUlU�,�{om9�L�f!�46�2Tj�n��]}Yu����%4��)��9�ʬI)�xh�4,�2�|�ģ��D3�*8����)sR ~��;��з�"��|�d�?^����ޛ�ϺWqkwbA��ӊ���9��\�%�/�|izd�S4{�����g�X�JF����ܡ`���}�B����1�q�^>���CS���L�]�$?E�g��{��˨,�;��̰�78��`s;6l_,Gܣ�ǚT*����}��.�z=}6�q����.�/�Pzz���0��̝�\�"�I�=��S�\ݐE�I�D`�p����n����o�W�N��x���{���TV�l���:���q��NQ[�_;�dʮ?<�����[q����y�T�ԏ���P��6����es�{k�j�3����'��w��(����<�;5y?}k��Q���gI�{��Z
/~=Sڱ�=����cQ:�U�;)�3����C�������]�����wb��+4���$ڧ��y�����A�eǋ��>�S�U&s�O@j�tT���d��!/�G�A("�s�seҮ�1VȬ�����:<Ĭ�<V�\��|D��gn[{ۈ#��<�߷�)d^T3ۻ��Oop<���������z���w�ov������?k�4�{�zE�쿨�'e����OY�.M�p��{f���x���n�`Ě����fX\�i/�=�L� m���h�I�7A4L�?��{5�g���g���TY~��'�g�x k��˂g�u1��c{�x�S��痽$�*���wZ����`;g��A�r�絙x���o��#^G4ZK��ϭy����_�Ǎ}N�
�\�ٞz�l�=���Y�M�52�_�Q��{��p���Ey����h�VP��󛘽��v�+���"W���p�౮�OM�ſop'r��,/�@�}A<���W����L�{��xn{3��"}�J����l��>_
x��}w�f����Q��ɯO��ܿ���q*kޓֵw�Z$������*�}]�����3.#��{c6��S��~�޷���}�%m��{E���{l��\ʧ�|4u[��q&��^�+25f�Ũ�偺+����QxkP}xf�i�;�P��Ǩ�wf�v��v��0Ȭ8�쾱ݢ���p�U�wF��H�U��g�i���	B~+>�[����'��$ њ$�6A�D�T���j-���ر�����q�:�}�k<&`ϯ<ugB	�o��&�X}-=�S�$A�^�w��sB�P"fxt�}�7x�ʻ�x[/H:}�N�;�܇�|ؼ�G8&�v|�?A���u��p"_y��~ʞ#sB�~/��Tɯ�gd�\T�<r��2(Ԛ���3jD�Nmm>6�Q��2zF\"��������[�i��'��y<�yBO�:��B�����q�w�_ןX����`!�=���¦{��OZ����[�7�w�\�~~\c?fC�pL��P�{X���w�yq7���w�vp�ߧ4�B���t�t6��U9̸-���m��ӗW'7���������p�}<E=��)nI��ˡK��<��Wʢ�ȝ k2zw=�9��75�[�����]��}˫����)b�	�o��l<��6�w�\�����8/c��//b��@��.�}��.?^s1mѬ�NL��w��p�73��p9�v�.��Y#/l_d	B�TY��me���a*�f8y{y6��IK&vC���c�����&�?[�eXj�����Z˘ͳ������ߣ�FY�'��߶sz<^	�2MW�u���^��P�#g�hz�G�e��o{�E�H��ޓ���93��UH��&����\��q����X7q�eE�笻����96q�d�e�\\תB�I��؛�&��A_1)J��`��H�}�G%@���\��G9����^M�E�LȆ}Ӄ"� �����Cf�t HM��V?I8��rK����Z�k�*`H�|܃~�@���w���!�a��{3w*6�/�ŏ��o�J�fol�ͬ $`�rOl~�Y˽��Y�M'�)��"(�y^�B�;+��&cgՑR3�W�h����4w_&h�A���g�gc����� �S4;��6D&�"�tq�|Xfɪ�C)�&Ӭ��׾����:�e*f�ի�	`�@�uw�/� �<�iȝA��>W�7�m�`�iݭ�v�u�N�����˘0wJ���U	�-
z1^gvG.����/��s��&7o��)�Am7;�:�|{wc�wr�
	3�-+s�d�����5���g`�^��v�=�W!ݮq5�U��q�7��v0׉�4 �Tn�m1�4��>��3�$A;9�dO�3�I4"�����j�o��x��7A4F��>�T������<�@"ޫ��6)��傭[�c��#��c��y�k�[��	���=��G'EF����f���/y�^��[��tЂ�#7����|���N��I�~�9[�O�ڒ����=~�}�����yrׯ�~y�t^�7�v�z�M����:z���<�'_�x(7�ǜ���Ǿ�w�a��[�ò9������3�Ovo����]A/�������/�C�����⑘|�=חH��ןG�>z)���P�Y��ջ:�r2��c�ך������Z_|������zf=�&����~�i}y��7d��M�HW�0�l9��vwlMq�Th`��Ҧ	ʛ}O}�=7�8��ul�tb��1�:)����䎾9Z��Z�Oq��8�#���z�
�{i蝝Z+J^'�ol�"�Y�v�o�]�vhY-=J0k���ŉ�F^�&��u�3�%g��dyj�Wl�gs��:��l��W^��D�~�?"��<屄���z�cg��G-#Y¢�^�J+]�Q�(;?{���l��dL��lWw�n��������Y$wb�Ϙ�6��I؜�z����Q���g�j�hW��;�d��"�j����f�9^&7"��u�8��'��۹����@�<�"X�rM߼gm�-�+����cxA��j�I�̝���NdU��_C	���S��v�4�������<�4�5��M���l4� �r�ws�m��^.:v|����w�E�����{u��$�ǈ�9��=Y��O�3�m��g|��]�Q����\z2��3/>g�Cյ^�-%]��{Q���8��<�Z�#״����끽�����c������W!s\�T6�Z��{GX�f/-�;�eg��YZ��y]�_߻�����.���]۲�;���5�)@�.*��1)n�u�<��Gu����#r���G��&;.2���������S���n�]�j%���e]�,T��a����r���Y)*B��y��ٮd��4��=�+y���Ow��N\��X^Cp繼�F!��J;M�kN�sy�s�����o������r����k�~��㔓!>�>�z?'
G�^}]%��w�N'>ߟ�&��|}�>�Y6�N�%魲�M������q�� @�e�n�m��-��Ϭ�^����*?4a|��/���sH�\3�mz&@�{_��������پ��L��{�S���C���bʿ	���y�8��jd��,wVΑ9�٬7���$�y�r�{p����,�x�u>^}��w�h�xOp���\�s�l�xo�z|Քc�6á��,q� �V���=�fy628�o��|/V��g9�
�Àɘ�'�Cf�{.i�h�tc�V!��&e)�ֆ�ş]��ye��3]_gt����1���ۻ=20F�Z��ʱ��Zk���	���n�ڶ/���;Dv�5�<�os��0]j��HXrb�r���{TT�}5ˬ�u���rPZ.�:
������Y4��[�K���_0���/M��R2�[uL�Z�0Ą���Hw�\�fsޡ;���.u���ݓo��'�vʫ`��X�{!�x��u_xz:��3_�鮼�Os>��6K4��Z'BF�������7�f��,?=;%�uF.�RK���-ѼoͲI'|�Z}^w��Fc���� u��;�ݒ:�}������7��<oͲd�>�t���a.�x�n�+�U{w= �'Z��rD,��y����!����{�y���U�v��ϳV��{����q��OlI�2Md�@I��߷���.�4�<��W�pc]��o�9��H:M k�oEeg��z����>Y7�	�h������\��ɼnk�sS;��q���l����up9A{��}@��s����X�-z��^Tt{��F�Y�pط��D�¦O}V �Xt��g`��0���Sj���o���D�<[ȴwp��~��	��n��p�8�}������=~w�����z�?���ׯ^�z����������Ǐ�>o0��z��/�M�[O0�$oC�] ;�x�mAfgq晴�_o&�>�h����$�ݧt.n>�`o^��|u���kP�\������{3��y-�±�_=����ղ��mY�L5c���o^�]�-�c5��B�b{z���v�v��ޮ�yQ�7�kB�3��@�U��8G�E�
�	�Y]��FJ�4�n�՘ƪ�Y���m��.�/H�H�2,/7WkZ��YkOe��&�������f�b��鹓.�*�-���N���g]�aS!�^�W�w+޸��j��d�j�;u�
�f�S�����d����
���k�P^\��k���^��������;{�$�s��Y��wE�q]�[`\�kiͫ�A�^/Y�N`N@p!B�H�
YCF���3x�;#t���8(�X�o:W�)n}�NP����]�<��Y��[4r��uv����""�3[�o��lM�e4���~��n�Fj��Ŷ+ ��»AʚWa�)S�e �i�8��ƷWi�B�a&'�ehR��ك��=���{8��+�k�V���/��Ӈ�Ᏸ�2��z�[�x`Gzj�iǉ��v����GZ�uvq��[�T#
������ݫЁt��8c�eh�8azg`f���3}\��*!�J��D�a�f��8�����+F�"�t6�u#sT��!|;����Ol5WB��u���'s�05!�4�Y��`���c��Z�ͱ����Ȳz�ud��u;�p�(��4�y��5�MV����&ʬ�3�������Bv�2�]#�/��Y{eu�A���q��Ҭ���,�3����N�>�/+����Z����)���q�^����hL��ޘdت[���Y��n֖���z6D5�~��,��x�۳U�R�e�K{:��E��u*;y��	�R����Vq��lV���[��]�O�R�We�Σu6\]�CDiV�G�t�DE��oE(ԫ��\ƥGӢ��eM��9	2�Z7��+5�Yś�>f^�7���ݎ��S��x��Z	5�շ1����/�t�Eu��T��֌�Ÿ0�����:���wrjr�=m�X��J��M�K��S}�����|KE�٥(;,VZȧ��l�����.n�OD�D�F�M覮�*����4	��=�,	��1���u�@Q��M�K���y��aK!���
�ݥ�Z�:1r4���E@	�V�Zm��g���V��������$9Y���YٕXpi�;�tLs�F��y7�B5H����6�b�q����YN�;ʳ��]�v��si�m��d=�o��sP{�ض��Hsp�Y5�-�l��¦:n�҂.��hќ�i����3����Ov�O ���/��5�-:�{,G�bH�[b&��ӊ~mE�D�ԅ�PT���J�s͊g�KC1D�DBLTQ�Dܰ<�Q@Q6��(��ƞQE5Eh����Jbj��%�-b�c�b�j6Q�AUTUlj��Zbi��֨��Z60�SE�EM�b��F��h:
()�(���-4��tQF��5:�@k�n`��d�D1��(h(m��TQ톊���4#D�RU-4i�݀�0�jh�&���;jR�$��N*J�f�J����T�ڀ��Ѧ�����a��"��C�tE\�)h�*�����h.lE����� ��gN�H�j[������"*h� ����"�͢�h�����y.G�:
�
���
�� ����[�{���t,^�`��r�k�9F����j<]��%�HL��s�ʓ�׹�
�Qk;u��ٗZ7j���[T�fl�q����ats�3�����H}$G�L��O�}oEC�xdK;{�
Q�\Lw^u^���[���UѯKBvg�N�6��Y����������=�Rpѻ�z�"�+��{��xe�yg�b5���a>��y�*���^����E��aL�ް0�����Ai�L������e����Y���S��~���~�//�xGM0J�;��qƤ�ި�F�4>EM�u^ZU9�����Jk��a��1�z���o������XfD	!�j�7�ª���Ԭ�7��7�2s�R1,��F&�JR�����K���-��$(�|@����s�����v������+z�H��H���It�ħV�E2��&�|�/�8�?�W*���E��X{^��={�-3[!�����d�7�]��Q���'+�R[%�7c��3xv�づ�VCU:����|��xC��<�?6��mѹ<�\�n9	�\����)<`	ƛu����WԜ�f�u�b�|=�$E�ψ|�Gx�va���Z���M��u���<�wck����ݦz��ВQDM�mU��c2b�a�Y�MdMd�1�5|\���S��]Q�ک�S.�Az�CJЭeil��oVǜ&5�)0۱��Q�=��q�)h-1�����ñ�ǹR9��s�����R$l������j�ՙ��{V��ʒ_�`JF�D�3㘑<�s��c I��?E�v��t����+	Rq%5����Q���Z�F��0V/b~+���z�V�*�L�tf�˳*�3/*$W�r�V.�M��^5�Z��zw�5\�_�?���#�Cq�ϥ�W��cN�Lb��gS �x�����f�e�7|�~�\ю�~킜Nf�$�g�B�	E���t�z0C�d����sq��֥wv�gX"��,�xs�vc<����w�F�4]��f->����4q�M�z��̭���p�'�p!.#�>�{&(ߑ���Ѧh��<]�غ�ltĽTc(����Y9�&��wB0<���'�p% �`L�#@{�d^�����ٶ���c���8��j�����>�,��A��b��Wx�?
C�r��JO�b�.���M�j�U�Fl��E�Vl���ݤ/`��!�'������x́,�2���`�j#�QP���T��<m_�����uP���=��Z�`�:����齈��
K	cOL����O��vf��3 ���2r��Z:�����hU󠩨�i�c6���L�
�Ee����N�����t�;w����JV,��ڰ�)���h���q֙�M�t�$̛MmXkwWUB�Fƴ�l�"ٷ%�'71�:��o6�i��CBv�.-;9:�wV�I�`5�ƭ�F�T<�TԻ�z�_-N�Vh���z=Ϡ�L;�`]B8#�p�X��ܼ�)Մ�W�T��oJM�Ӣ1dgVN�VZ�Ցm
��z$(Ɛ!�&�R6�� ^��_s�T��ۋ�I��{��V�y�w���okW�W���;�7�`�1#X	�F����8���a�`.s��V��Kc/�z�:��xů�n.��`sJ��~m��v���� ���8Z�!�n�yQ���WMj����u{Fg8uV���Biyms
������/6;��;=�,�8��X�j���������>)�:Vt���	yN�������E��<ʬr��P��}j�� �p氣ɫu�������魤@���q��7VI�~/ҹ�I�zc�Q�$�:�0Ȩs�Ƭ^t����}�\�Ђ�8l.aٕ��ܰ��Ԩ�O�Z��a�u��ɍly�u�'�X���r���P3^�^�9�l�t�a;�����<!�ܺEڄm����Sދܻ7Yep���=��j�nנL�1���1�@�	<<�/�a֨o�@P�U~��������*��IG*��!l%)�4V)��g4�W�Yu��X�9��6�Lǳ��}��k�{��6d
�E�_�=�X���mhЛ��q.�!�����3*r�aϘܬ-��'�:��n����և�`����*��=�c�)[Sv�n�`�����x���7��^�����!��yv�Q�8ʺ&��E��m�H{/ỽ�5�o^�V%=S��\*���i���v(���� �{Jq��^~�a�u��~�UP��A�ϧo�k܉���{������y�Ɠ0��4�^��eB�Х`G\=oM���m6���H�W�����K�(����ъ��A�5ΏuD3gh�7��d}h���8{��u�?`�Sْ�۽�w�|-{��b���@��v�[O��/~˩		���;�S����H+�$��wј�)g�{�k��r��	�%"�;��6���>T��`r�
���>�7��'0w>�C��9y[���f�36���7��ɷ@�ht]yei*L)�/|e�!�VX���#iq~���f�[_J�3�3qser�؇�4�TWC��N�#0����PMCux���;�ׇ�If,�i�"k^�aP=�[��- �,�P��B`���2�ěS���Z~k	AcAt�~d����+i��u��V��u���G�5�4�y��bK��T����ZJ�.���QWC������K�x:�Y��hH���f����*��N�3���
u�o/���.Gf`d�eb	�[�ֈ_d�ܜ64j�ݥW��=��P��[�9�t��}�$)g1R���&�Y��
����d'���o��R�7��{/��X�)53��d�>��٧v�a���T���x�@#X):=Ý~�1-�����0gh'���\�w5:�b���J�Q����y�)���&��Y ��apY��\`43��_E0	���-s%�=�ʳ3K����X���џN�3�G�Y�x�Q�@��
���T��j����&:(���+U�v�i~T�3����^=%� %����,{�C���.�����6_��3¢�X3O_f�hg�f	����]��tpq�懑�X��{���P$@'�@��i�}��y���M6�g�e�9�u�W
���0׎r�SJv�'�#w3Ez�K^*�!��v��g(������ν[Go)qt���N<��r�Ԃ�ώK�S��tgDX��3u�7��p��L5�_U�����4�?~�E��^>GK¼�钾�?T
Q��j���%V4���y���b����Ow\7o:;w�A���5Z3I��z3
ޭ�z��&�K�����j�Ά�f�m����J/wd����:��N�)���<��)��R��q��C���	X�q�ʴW��������FK��c�I�T���/�������SՉ��3�)̄�ܬ ���w��kGF)�sG�c�n����U��ô���8՚�Ӎ�}���2�&����0�.�o`�xK�.��oe�9��䪻��2l��35�ƾ��>�����o�^[t҄ŰR=���= @~�N�㘔�t	mI*ML��$���|o1�S�����2�.�wn��/,�����L�Gd�"�K���4��yNR�)Ph������U^���]��ܒ)�N�� ��Z���X��9���(C�rTi�^T�I�M��	�O��������a*.��{��	�_'��L�	=�XE�1p�-B��5>E�^��:}�����˜��e��͎���eἸ���r_��'�cc54���c>9��4yf�E|f�A�/:� �ڬ}�[�AkY;V�[�����z2��G���l�l7���u�5�������܌=Jw�F�i���l�np"�K�:8dR�Xqg�X�	��u���ҏ�$;9
I���2�4���u����>52�?6�.��@�T#{e'�3L(� �x��b�-�nզ�v�áK+r����\�3��P�-��	�D��7��X�İ�}�B(k��(�v�z��B�|��m�氓��KǙW9���:�H�OW�-K���\sH���.ͬq��tTzCO?��{۷6��� ŗ�����G�`ҭ��0F��h+�ֵ�Bă�w⟬/^C����^WR:V8�f+"�NY�@^��ٯ�n�=��Ū.�쌇s��x���3t�K3�E�p���O���x���C��+k�r��ݲ':�@х H?��<I삥��s�o�ͷ�L��Ϲ#y=��)P���>^=���;�K�/���Ģt��ߪK����'wycO>hp�}75x���f���=f�2���Q��������z*ٷ;���/�qim��ʋ�3�
�y��oA	�� �Ӊ�zYhHֳ׌|l��s�\`V��,|��z�Y���9�D�
��󴁪u�PɅ�OЃ-{�'V1�ҩ7�5.��M�tt��I��V�gmv5W���9Oܹ�滑���`eJnj��&I��bS��ؔP���Uy��6���r�9����l��q���Шt�z�����rNܸ|C�q�i&�ҟ�7�j�?'��A�yS����́և6�e"��h��8_�z�Xf�� �cH����� �y�	�M�mD�(|���z|�W�IA�Y�ء���/]��ǵp�0�bb�r'8V*/8 �݈n��6��\�f�n�	G{xj��l�h�""1�@~C(Э�X�i���dâZ���`%%�v����vh��T� �����h��kx�e��xu���yNh�B̓uœ��:y�*�a�/v���n��?�E�؉hV@�X�G"T�M,��x���j71fP�h��
�[|vU��!�[Ȟ=����V�M]|��xв���5��Fz�v
�)\5�[aU�Z�߫��+-3���WMrJOW�웥T�e�3��cz����믞��(sU�������o!s�ēz�Ő�����!�� ���eS[$�C=�Q����\�����o�p�ΪFeQ-W�ٳ�Sc�K��,XCH���x`0�9oC_��g�(���JA)�k\ռKi�-��7x������]fa��t/@��vhB[�����C�m�\�2�(W;,�޻�׌ʚ�v�$���R�%���M3z�3.���C�[9y�����jE�/��n'��+�?OUy��&[��3"������ �9v��-�{�m����3�������fݨ�E]�qW}���qAYp�ݑ�� �{k݌c���B�/E\�(r�xY�F#�y�k�&��9a����6�Ӵ��Wd0,-��1�{��]��-mZT��`a�P�t)X*�����6w���;���Y&T�C��+��.e5�h���i���+dc���Rn�2&��/�cN�9u�׺k:��xn:VP� ��4��X���0��BI|�&BGex��ا�,�S1�e*n�}�ތ�A� �ulp$��ϻ�{��U)���#ʒp�c�p|�'������Fϐe	��e�E�G��؎剽�xQu�E�u/���7��7t��Zk��h7LM����#�	�v�ph&!r�/�k)վf���@�^���(dB@4t{�o�zŭ�T-�7���L�3�9�"oi\h`0e;��_�k�m��v�j�3�
�y��o�������0�7���z�J�Gv��|;�Ru�bYX�ʂJ�|��%���iЮ����q�u��w�w\zU���΀��pe@i�rvGdQt�ѩE�y�)������V�"s��.gL���&7n�iЀv^*�O��P��e�س�M'qU�����o�O��Ģ�^�.���g^�~E4N&�ǷkP�u����q>R��uy�l@�	ј��Nл�*��)W�.��+���E�����w�w_C���+����a��c��M�n��l[2Z�3���s�lk4�=�KK�_om#n��/>�u@?6��f��?� �N�������h��|�7[��xƐ��n�İ|5�K���E�l�Ll'���N�3�ע`���f4Xg;�+��.�����Z����H���q����Ў��6���nr�if����D����zb��!��ø�}-�b\�B�4;?2j_���A@}�~ޚ�deFk��q��vq�����H�D����5ю=X�z29]Ufλ]]'��@2�Px`�
|Q��T2_�{j�E���L�}�Ra�����W.�e%e%�˳�/AC�`�Pb�Sݿd�p8�%�d�>]��ywo���,�fg {���98{9�H����G8]��܀����N��9�LWaԌ��ռLD.��R���$��!3��}=��gJ{�&��+�/���(�+JR�H�?~����ߏ?_���{���f�� ��� [�<z�sK�3�ܹ�UO����^��:J��������N֙nk�=Q�԰7.3l9�r����q���.F�с�y��I�*��O�{Mv���G[o�v�ݝ�tQ�֑�5����8������[�z�a!t<0���y����J��Bt:���2UsW���≉d^���e��*L����ֲ�Ϗ"����ھU3��-7#sݛ�
��a���¡0��9���_L���%?G�g��'V�E0
�T���vO0���q��GW`9X��.���/�Ø�Y����ʄGG�4����d�$�c���ct�����+�L�U����{��{����5���A�<�>h���D&ژ��#ry��� Cp!7K�u�BN��
��ʓ����QϖΗ'���f�I��E�3��F���s���M�m��no7�O�X�׸��]���h�E�W�K�e�˸���*wIו�ܴ��-��B�PG����1��_Dm���u�i��cAOU��AO̳���+�A����n��>�C�x0���[����}��}}g�������ׯ�G�S���z=>���2zȼ�l�c4���GxWg+f�p ��7iN#�4Crhkf������"kTlӣ�iW���2dչ4��-�r3�^�i�Er�p�<�cOT�s*�ëj9�4�t�όn�g�AG��y�3d�`ť�_2`Ü�c5��ڄ=�\[��ضF��U�w�U��R���vRh2����&v:j	@�:�n����;�#���Ƒwt�;�f�p�kQdY����Y���.��)�0�tQ5�K船���[�qPI�txZ�5q����QM����k�xr'^Ƿz�hµ�Ew��.C��+\2�UQ7Nw[ʷ���� ܔG���|к����^�]�JB���6ľ��Ӽ|��v
P��e=X�(J`d�|�<��0�u�ˮ�v-�o�Ksz,�h5x�c ������i�Y���T!j=���j��u]��ӳ4ܦF�Ûe��Y;1�M{E�uDN�gU�g�ʕ���VD%��F�j���2f٫I���j �͏��<nv�37�fH2��;(smu�p(i�LԻ�j���%�'G}������-��N�l#��1[v+m՝�k]4Vc��*�=���I2Y�0�*[Cu�f�h&��4�ѧ��H�P�d��9S�|���t���X��v�q�bª�l�����T�
�$^�i��B�����n���~6��ͪ+t߶)8kf�r�f����h)
ʹ�9V#��g�uI-���%�Q@��x^���i�A��yU��B�\��66r�܂X-X]"h��@ ��kC��Է�&'��ˡ�a����n�8�%�\\���_:���I
��{�jb��;�V���@d���F�"�`X|i��aֆiu��,Y���8IM#u�m�(�H39��B"oj��i�"�f�|��k�t��i��m�dy-P�h��]�P�����	@�nglЀ��b��΃q��P�9>�{p����S���A�N(wgn��!Y|*��wL�/C9�m�ű���f;�nLz0��[��;G�k�!Aհ�&X�ă(�}lR9�_1}(�%e��geRU��ئ����]��9��Z��47CWY��ĐH�r��cIqz:Ї�N��ƥ�� #�����{�^�+�BIU�j�<do�/*�����qm0��/��q=I���[V��\�u�Q���ovn;UTx7	��Ks9�#�&��ݫw�,�#�_I�X��ʡ�����v�	�
�j�.��j�U#�4F��P�s%^�f�[aI�J@�RԆ�,��y�((�lj�)pan`3z�)���\{A�P^��ܗĒ<S�Ǯ��q��wK�,%X�����->��t���՝�Q�(j�n����]xZ�����X[Fe�;�S{I)	����u:i�;�7	���(b��B�f�i��$����K�q�4MMzv�{��W�qN�{���:of�l�U�"ކu�;%)��:v}H�rn�N�ه}���XK{��j�F;s��%@�`�B!R %@�AC�L�P�Ө�)`��ۉ��t��j||��}�
Z*i �ry&��SrE�:\�{;�4�ܢK��EOŧ\�X�'��c5��lUbo7-�r�S�(�:�gd�@A%�TS�킪��<��|��X�M��yÞ<�6˂
n<�4��$:���s 6�1�i5����s���6學���4P'����[s�"�2�����w���Py��u�#UI�5�JDspg�&ٹpy��7�r�r�q1Tk��;���G��)<�6Yv�"��N��˗0�h˱6�f��4�3����y<� ��nl5Dp"��<�P؏��dēI-�cDlDTY�*(��k�t�5���ks'#˓���l4��8�B������R"�N����'�o�r9!���9�<�G��h�1�(+Z8K��N �y����9c���F�<-r14q�����c�����lZ��y|;�Q\�ey�s��S�.sSE���X�8��bLG��y�ThyV��1A�5�8`�6��	�:/6�"*����%�i�9+��F���
�u��AZǜ�)���FJ�I��F����gE��^F����Z'E#I�CAAEm�^?�t|++iG�Ǽlp[(+X�3��Ճ�c�"�nUq�0��y�WR�RO��p�\�d���d�'3Mr�����{���U�79��E�@	B@�A2��O���ߟ����>77kY�9�އls�R�$n��$��/�\��N��c��a�=B��Z5��c~�[�ys}��=�1���G[�T1|�3M���pS�	�&+���C��(�I�wqe�Ճ��c�o;��3�B;`]�-�����`s�����-�B)���ۀ�C$TmLD=�]�ed�q4x	���X`N���M�����.l� p��d?����$l5^5<��C�}\,�v��b�\��)�A�F@v�o�i���{dS�{b8*#�����asT�$�c:��r�6W�R���r���0�T ����;�FlS+�b�����)/W���k��i���=�ݴ�#�T�#��"��VzPN6{L!�V�K*H�3��H.×��ΌT�\û���5|	�<5���!T!�#�,����A�[ތfa:�F�+�I�0�8d�B�a;���ʒ,U�w�^j��vS�����="r1��#�>ʎ8@8����%:o^��*XN�De-1�=x(�s�;ΆΰB���.2q����k���_�:A�Ð�v�n"���
�{=3&�ߑ���*�)�ܼ��8R�W���V�h��ӵd<溃�Ԓ�D7'��V��f!����[͔KPa=���q��뭫��U^�i���Zel;�����꼧����K�Y5�z�e"�G��`;3e�wx��[������@�(% P ��"�
,*�B�@��y���v{PnJ�z��n���b��_�I�y"h����H܁AƑ	��0��+�&zޮ���B	�~�B��uCHV���'��ɶE�y�i���nD⟔|�S�
O��@B��F����޵�7(�w^���ю��Q��J���
����Y�E�ҒƑچ	��V�>8�Xk�ܺ��K���:��.�[�Լ�E�B�x8ⴕI�)gO2�S�4�}`*�y�-OS��J���W�����5�օ�����^8��/ҹ�(%퀿(mj[(����������bKP�;��q#���p؜��fY>ܢ���]�P-�s���ֵ\D*�%�;}݋�֨fv�F����?@���}"L�w�p;���w�냵��7�uc3��H���Ax����Kԍ&�$�a��u�f]�����<V��.��� Օ~�]j`��g��r���dǭ��a�2,�� ��P�H�e�N��U�:�{a^Z���N����p޲
�c2�[�o��G��[�K�xf��X/@r�F��q�� ޏ7���0��� ��`6�7 ����(��O��>�-�X�*�_+>ύ������)�o�oK�U���S�(��t��o�>^��K���Vcx��Ce�T)ef�x̧�۵�l&\�0�]]û�Zq��gV�ؖb������<�������վ$()BdQ��Q��� ��i@�@�@!�~���m_���tS<`�a�"�h���=�r}T�ڔ�A�1�{ʺ�ע<ͣ�#��굽����:fۼՕU�g��&��X��8�+��KsP��Rn����6Խ��K+T�l�i{�M/�E��&��?�VQ�WDx<�Aq%����x�����^)�I�������L����s�s��`��	*��ʅ����~����&�(�<�����B��!�Q�)�f��p�Dp��e�R��^��2S�bYX�ʒT�p��_ì����n�GG{�K��	NU�`��k�"�w=.C��ihvQ��vEL/ڋ���p�T�P�_��dۖ �kR��+z�əl����A������0��>� �P��{
7���@�n�^�E�气 ��5����W������ۼ;��Ļ�Xt��#�<��s9�rbS��T����~%Q� �^>l$�Bz��=��{܀%�۠��]퐌j��a8;#/�ֲ~��~�0�ɽ	���J��Y����{U0¼�yJx��ڰ#�|n�k���GH`�à<#�ȇmt�o���,�K-y^�ݽ���$=��{�`j�]"�YKu�)G��䤬��F�v���&\���fa뺓UKK�J���X�]u�e<��;s���3s�Pa�sY��������:�|v;̲�.�����7���V8���:L92��>���*4�*���Ȕ�-"DH	B���()B�0�	B�?����Iwwn�j瓱M�x4�i����֓�^�r:����c@ņv<}���?_�%B'�G[1B�s�R6asP_u���y6�d�l��)��^=%z/�06�>�R���:�;&�F!y9s �鉩54֧�n���{��&$͗���t�A�����;���	��m��K�%t��̳���ޫ�B�*k"Y���-M(d�l�Н�Y�F׺��=BW�wK��6�N+"��m�uwJ(�wY��xi���sKI
Lde9�U>>��lz�ˣqNE�Ȩ1�Ը.���Lڑ�Z�`�BF}��l�zǭ�D�"����<�t^}�o����ࣽ{�h��Vem�^�az�*+��Bk�d5Z3H�(�0�ј��[�z-�d<��[z�n��96���;���
�B���� �&���s N(ʌ8H�2�J�Mw����{gNU�=L�!���]�_j\�b�r&��6�V��!Aڎz�)�v/	�x��L�$�5�ȶ���1S�Ad�*L͝�&�����ܾ_1�x�ނn@���}���@�F����4�㘤�?����'/���e��b�q��ޗQ�/�/�g���ݵ��jG�z� \�^�nvϸ˦���-PX�2]�g����n���l����,ӥ��IIu�aj�|z��OD�����⽙���g:=Pxv�tځ[��1�	h�ި
�[ز�����w%"$�/��6
e�����ު��
��TI	J�A$+H�,
�4�� �QB+H�
�
�2ЈR^�f�7�<�3}+S���/v�"/����������1���y�CE�3 �y�x�}�����lfO5��a�~U��6ʆʾ�Q�|�ݗ���ˤb���R	S���;\�����*<t��Vc��uĆvZ���]�	$��F�=�إ�-��e��s*{���'�C#\$X�E�}�d�P�<EÜXu=�=w��ΞL^)L�.�h��l�5�v	�\���M�*�g�T���n�ql�ѽ�0��A^�������a��=S���%�_'ۆ�� Ė^/�^�OO����%�ÏPI�W�\��Wr�'gNV�N�b}.0>��lZ@����̟3צ�m{���`���
$@:�7<�xX��W[;=�}��1�c W�B,pTJ.���B�[W0,�xfH�{��+�������?��5rG�����k Lq �/^�x5�.���h�q� D�N��S����3j�Ut3���kkM��K7r����	�]�aN+ﷺ��֧�Q��؄�CX�
��ۻV�h蠔)�cy�js��y��IXkNPq�a梮Pj	�z͜eX��|�b��ߏ�����i$�z��6�Ekl��1~�7ޯe��6�I�l�/'�r�;5��g55B!���f��_u��j{ݒ�B��g[z���OwN�^EL4�ؿx���_j1�������We�A��d�(k��'jRj���8 ��?�>�U| �T0�P��AL��4*��)- �дP�2�P�C(� � I*�(4L�
O�^|s�}�������/"�-��Ǳ�dc�6{L���xa���S*IV3Ҏ��65�ͧ�mT^\dѪ���/�C�g c����B�x����k�_�ּ7b���
O��i�fE�E��;-��۷g�[/Y�ƭ��un��zD&�P`f	��c*�����~X�r�x?F��'9wV�����5*�ҩ'~��1��?�2(��t`5��փ�~�p3e�q�/8�ywz��f�rvB�u@�LR�t�Rt��H�8^���H܀�3cX�!?7��0Sr��L[��λ{���	�\C{0�sס�&m�E�1��!iy^=5�^w�~y��f��h+�l=�5��~���y�=�@���C����Լ�FL�;�4�U�<�Y�E�ҒƂ;P�3��p"}dDtB�^@����6���@�l�0r�1 �OR�k�в^{V�����<ʯ��[OdǸ%${�uV]�Mw�Q�/ ��+�
�G�+8P��j��f������s�&�s�#K˦�_*<9�7�q�I�KU�>�BN�W�>�(AUg�����9��e��E����ye��?��h�6,!͸��Z���.'��v�"��D��gc��lY����*�&�g y_c�v��s* i��hug�y���	���N�浄xl����s-=��=��϶�C������3�L���*�^G�����e�
��� �4���A@�ą �H��4�R!BHIP�J#$R�O�}�����������߿_=;�18�#ӴMKsQ�^�/a�s>D�c����D(yK@?HB�*�N|k/������F�#�6݅bK׉�c�@����D[��^F���\Cz��n�%�Vu���}�AYu�y�����t��e�t�_��Tyv�W���+���+�}t��b���ST����c�V#���3'S�T^=����s!��}�U�B�#B|��xfW�z��]�\<�]���8�|嗆�\:ז{!0�Xr�L]�^�TcWX��%��jR���e��=ټy8ԭKD^�g_gWt��������/P��3�Bll坼���$v�[��w%va�{��{w�B��2*��B�ߥ��f3���V����xk���I|�0�f!�(��yn�t^�Xd1)��%0���(,:&E>Eۭ}Ǆ��|w�Hqlp��Q��C�V(Q*�HyB`Yf
(hN^��'��he��,��)��&��qA����w�.���%Z��fv����:�͓�8�	r�v4�T;(��~ɢ�t�1�d]yd��=~�Oս�|�a�B}`'ל{��d�k�W�j��lN�e]� �q�Æw�R��i���m�ܦùLQ�`Ϊ��$P��<䴛KX�n�KK��*�K�yܷR\Öp+=2,0Vu��&�.{ws|�Dx�-G&\|���߾o������������P��!@�ei@`�JB�(�)E�Q��Y��7���s�]�Zk^s��=y�^C��x ��Y�!�t8-�;
8e;�O��^�V�(���ڲ���İ�1�d�5�{#��:�$�[
���B�fm�1%��,Qӵ�m�q���ѩ�y�S�n��En���;�sj�u�8��WC1OSߎ�J
�8+#,�0��X�6'��udtp��35���#Uor� �!�լ(���`%���W^z�m�~!d�$ ^a?�<��#q^z�ֶ5s���N^Z}������]
S Jx�}&=~���i�,Ƽb�;��j�S0��m�Zߛ2�ꎜ�\-C�m���>�v/�3'��'rI�no��/@ %����� ������B×�=�Q��'਎��Ϋ�ծ�͐���vq������H�Cz �zd(�����_mv'in�aQ�w�~^ؖxBKHC!4�w�I����{87�kN�f��])���n>��fx閿{iB"��k���v5 �z�ܰ�3�PS�x< A��Bg��s�S�����7���X�8v҉���Z��3nt�����5�\_*�D�D���%"�/�v =���C�|�����~�w?\$f�yk�`�0�,�9�����Z [%.��p�]G5al�܂�j׮���$H�*-W���N%|�T��v
�J�z�6 ):�����ccb����Nm\R;瓉�x9�y�fd��𞀝�����(�6��p�H�P�_���)@H�PH,�J#0ЃCBR!R����9����?>{�ߏǞ}Z��}[��,1s�^��%6Y2�&��'�J3��D����{ǌz��ϙ��Ƶ��k�����Aе�%����<�V�"�UsW��	P	xd�-a#4��)Rk;��h�8�������%�t?JƠ�.�@�+��MW��~��Tn ���^��E2ۥ	j�����3�]1ڷ{��KS?\c'ȸu��m�%,���.�_Aw;��O��w�^�~���׹��9���:��a�D��������0��@s�3&���0ZS�ä�O��2�ni�Y�ڡ����A����K���uf�{h�=�>O��q�<X<���7՚���q�VM7^�k[���\P�4��s�|Hdk���~-I�.��%�ǞZc����S��� szdJs[�t�]=���%9k��&ެ+����طvm��@����[<"L)�^���'�@q�D<���'�y2mz�G��\i#S�[�����e����^�m����+2���6o��}7��>మ���4^��>H�4#hv�N��@��7�݁�uც��M�y��PJ�9�<I�R�v}��r�VR��A{���>�m�n��+R��w< ��7؇�3����C3Ta]
����s��k����~�H����R�y݁��
��'lG_�*�q̧&D��������@�\���OB�g��>�}��>���
� P�0�H"RH���[}���^u�+�z�V�z9�p�,O�B�&S]z`8}K|.`Y��uosE�,�gh�^f4j[��R�/#4����ZY�H��I�^���l�w����L@�M10��7�9,�T�4f���^_f�)�_�ٖ[�#;��jM�Ģ6�w�½h4K.�ʭ�o�}�vs�C7�nՖ����`���~穸�������]� �����g��U~���|k����y��&���'�uK��q�p��"1�3r�9m��N5�@��YRF��u��=v�D��og�c����e�ߪ* ���Rǃ�B�b0/��k�Xր���F��=�-9-��WcZ�Y�V83���ܧ)0���8��o\B{aє �����P�Q�.ޯ[��㮽k�;�z�.��I��2hӊQӌ'ݑm
�aZޑB^1��(C�C)�|4��T~��2~�Q�~v����=J�,c1C�J}	Ml����:^����7dxBF5Gpnl��g�s;a��X!�L	��	e]�������Ͳ.�q��K���x�W=yߙ���=�O�����x�z����ϯ���������>���~�׽��V��{�v0��s�}�]�m��^�],�[�muB�)fق��Dnb�'�39��p��[�oW@�#���������@����t!�z�@�0^����@1W����3�:�2�Q�i�u��ݷ�d���E���ax�m�;�N����Дzh���Ք`��)E�=☾��z�^�F�t�w,�oN�kU<N�\���;n�ӟ2Z�]�]	O{��J������-�qn�czÚ1��g�թ�&���n˾o�b�v����Қ]��8����抏6����ɧ��\����Z���8�k2:٦��Ay7�=֘�m` ��i7�*p���L;c �7P�Sz0f`����=H5�o9;(f���O)��;�4%��r[D��K+%�
D�{f������������D��xu4�j�5��<�Ѽ��7�Ò8�wس(�1���e��v����cn�ӜѺ#1S��u�m4yKכK�\U���C?R�O,����F�]^1�Q��d��j�w�Ca>��^×�@u�w�F�����BJ	���[��]u��@▛�#9��<������&�ޤ��ɴ��H���b,v�}������3Gtg4���kQ��K]3l'2d���-�wΎ�Yr	�1l*-6�Nv�Gy��(��aݏe�����M���f+����(yT�
�W���`A=�ܜr��)q��=���%HLU�[7{F১9F3C����gU�㧲��<X�8�(�1#؞V��[����;N4jY�3�_��K�Z�x|��6�Ϊ̂o-���jX���_>|��1���-��}b�<j�4��1�
t��w�r�}Ku�wX�PY�]�Zj�j�E�eݼ��6�e��ě�@K�:�L��3��lܴ�cAo]��j+R-�$��Gq�,]�.U���H�6'�,�KҨY���W���X�ZM�Pqղ��_74���5���VI7�*T}]�R���S����Xֵ2-$0b�Pعc7'cو�}��wB��P�L�,٤��y:���[�r�9�A�`�Wx����u�(�9i����
�N����h�b�|J�v�u(U�"m,�i0 Lr+�[Z���#����J^��~n*�ܓ:ޙ�
[�[�&X�]
jTҸ�屇���rڵ(b��y�B�H(����ƭ�y�iΈ�koxYckTf�+C&�S�.�r���]xT�k��Cr�z�`���-;�ʶa����1�����V�'t�(F�k~B����Λ�[Z�h�d��u����g�
Q�:�ҒzAA���Z��VQw�m��0�pioX�B�JK���u�X���&3��<�(C�o��w�W�!�Z��1�oq��mq<�oKu����^�%�=KbE�{�,�v4tV���`���9�v�k��or��3I]���f;�@��=�=^�����Th�-EMW�����9�9E,�\��xk�I|^p<�TUb��J���J�� �E��E�<����K�Ǔ��E�X|��T��AMPQDPU͡&�B���9m�(�U�r��i�9�rib��AȠ��(("<ǜ1<ڒ�h��%S8"����*و�0RPm��8��A\�ACQ�qEѭE�Q46yb"����F٢�Z����bf" �Jb��(X��o6��HT�O#UG 154�LR2r9�-�%#Q�MS�Ĵ�MQM�r�CF��Ti�p����ST�LE�r�Ql�>x�X���P���y9������%3' �EMs6u5EDAMsf�V�	��ij�F���S$I�h�����' 4R�RSs��$IT4�ASBUMU���wc���zt��^l,�'%�1gs��$�
�3F�-af�Ȯ���#�w����Q����Vh���x|������|��kV�큄��!�y�C�A~ΣB�L'�J�9P��% 4;P�6܂��k��6�ݻZ��!;�!��)7L@-��^u�uo�$닿���,��UV�^
�}�ƀ�|�F�es��ft�Wyq��yů�pZw�[��Lj`kd��6,&����]]��L,���_om�n�(���'S�a���>f���t�`���3��Zb�х��a�n�눐�YҴf˜��Kl<d���@ӴMKsQ�^��g2dK���D&�5A�����t]M��n���e�n/��6.ܢ�.�����x�h?��K����ޛ&�+,���y�v_u^v�@����_W�nq���;̋/�	�@A���iD[(ԡ��u�R��1m��������`�/	g��A];�be�����U���� �U��܅j̋7p��V�j� *�j�S�罆m�8G0�`u�&.�ت�j��Sz�^�Ԥ-|���*	�x�n;�FoR�ڀ�t+�q�����N��Q��j��~��`u�����^��$�o7��-��Q���71aW4���>l�ȍ9��{�k�yc�t��:�ő�/�rR��τ��5�CUG�; e�x��^�c3nvЦظ�b)�W��;j�@�\�֩/3^N�7�Z�8(����ژ�pv_frp��]��� � ��߾����+�>�s��+�3w��7�<$��2*�hR�C����L�>[ռ��Ol�(�Bx�I|���Ҙ��f��1;�N�-W�e�9�?+<����),:JEo�g0�ӣ��u��O�����.κ�Tq�Lv�o������B�o���鐇<���	�5��I�/���
d��ß���Q�;b�d����������֖ s&����b��2��#اa��y.�hF�Y��Ow;��]Im�W1b.�����NW3|<�U�	i�-(f�~���`;�;
60�wqOK���9
Fض�3uD�����y�(Gg�9�29I尭|A�	(i�� ��O���4ħ�RXg��<�(����wyݲE!�R���;�U����q�R��t�����6H��P]�v��6QU�9�;z�'���Z�eV�z߭I�a@���`%��ׂ��A˖n熅͚(U�0_��S̨���~ɛ7�osp-�@C�>�ó+y�ٶ�ot�Oަ�ϧ_����cF,3��^�ȴ.����\u�X��B�f�Y{.��O�!�'rQ~��'�^�h<|�;��v�-�|ᵻq/��KyՊ�to�;Z��6kޤWu5)[��{�EW3�QJ(�������]hV�׼d�`c�c��Ρ�|#ح+5D鰉�u�� ��}����Q�\� ��M[���9������nw`�|�_���$���ae��gh�x��B]��M���`3�)�I�*����9��x����77�b�^��9aC��Ĉ�6^�ڌ�K8�s�8��tnؽNʙ�QP������`T�;O>�H؊oC,xg���B��[D>2O^5�{�z�� �V�F�cn%��ۉ�F=<�%s��(�p�׳i�s�ǡ�u�=b9��	�FFNq��Y���B���u�z�^�^�[�H�*����k֦�&���Y�����WI�\<�1�7(ld�ʪ"{�wP@]:�%D�clN�zGr�	�5.�/�`�z3����&�DC�vZZ3�f���d���7��ղ�����~��&%�{�Fi�%)�����F�=CS�2w���V@�<�W(���-���5R!�1���_�S��ħ[�o�ܧ�T�眴/�ޝ�᭪ʢ��s{'���k�� ��t��a�2ۇ`����Z�E])ጙ遲ou^�`�:��U��1\�`�)Pe�XsX&0�>G�e��@A�"mLpm��߱5[l�o4ۚ#6�wr���:�f�M��	�O�)�.O#�F&p��`9�4[�
5���~>�dLVf�*xi{���E�z��V<�^�C����]��C���4�p�!z�z���;v�25�r����k0�;+�5�|૕�x.�㽶�8Q�:�L�cP�/�ۤ�
�K�_.JB��'���C$Wlj��X���|>��(S��6�xd��ղ2�3�\�/4H��~���Ri!��E�n�"s�j�Aqg�[F�;7/N�C<�]xDz��N3�<�dS3�mv;�'-~Zd�ի��}���T�'9�K�yX/���j�vjBY���@jD��L�^�u�=�\��`'Ӭ��>��=��!����.�$��^�����UB��U�0W�B�58���9�Ǻ��^���:*oO�s4�Gov.`����h/��^	12��XXQ�~�5�[w0,�g(gL����Siz��w��Ԋ��M�6]�����`:"��E<"]�?bǞ�k�umf?3L߽�vr0
F_W��]kM�`��pwI.�����˴�}kOC�m��CdS�F��UÜ�Iy]ʷ0RAl ��垌���ɶ�j*� ��T �3��Ų#+��V��k����پ�9���zw�X�#�����&��U�j��X�'�j���׆d\K郑���;Nu�`���ʋ�Lu�dG�� A@���Bb;��aF��}�~X�߱�~�_�=G�#:MG:~KuC���}|Y�U��F1��D�j�B�eNʦฏgG�R;�f5#��-�T�JoR����ӱǩ�TD�6Q��t(�\�/c���=ט���	��ސ�S���R+zl�����F�G��b�+�MvHk��7:���>���^���]��rT)X�I�)�\[gT\:�\c<zD�(2.��N�N�p��!�u��,*�y�ǚ�?G1Oa�Jua#BՁ*��G����	�d[B��k�	K;$6������x�ȞPdñ�k�ۺe0�ˢ��3PM�Z�Rz	%@��g����
��>վ���f�54(َl20G�]hv����ߢ���{~�j�%=�d] �4��Kφ����$�������%C��n�P���r����Cw>	y/��hQ���
9�[�\��~JKLt��wR�<�V����0�)!ޥ�|���Xq!�5T(��:�%��'S�v�5�g��zw7/9����[)m�a �}j���\0g!Y� ,�CW��1f��d{��=B���:z��w�S��`�i8^��Z��{��?j�K c!��J���0*X4br����gQ�;^����b����,��ԫ�:T��b[�Șf��j[��8�\�r|z�CȐ`>M�be��jΌ<�sh+`����0̹��f���L(\
&�� L�˱�ƺ���~p�����F��|s�>2�Y�������%����$�/p+M����ἧy�յ��v����4ޕ3z����۞�m��o�^ɱ�8��[�,0��Oh����P(Wp�Q ^�
�[yr�Y�og�%9�:��C��7U��p�P�2LZ��2����	�w_����(|<<<<�2����n���@��^D<��훜dsz��fE�+�A4��@A�Ñ�fyڞ	�e~��w��d���P��Uķk�m�pB,��̔��T^?}J�c�]����cѨ�#��Q�CUK���;��ؕy�\m�j1p�0VR�(��jԖ�gͩ��T짮�4ͻMnE�0�ɰk3�n�j��0C*�t)o���p�7��M�T9����M����q�K��T�g3�W]G^�`/��6�o-h�	�v'�g���#��lʡK��a�Pp�!W��Xn���>{�rkS����.^P����=C�5�<������Ғ�5BJ��l�>���z��g�k�1�v��j.�[!��>T� ��Ə/�� �I�/����PJ���s5�zZj�'��힩ˡU�|��z	����b��(��*�a��+�h�a�mJ.�����1���w:=���ܟ��E�PƀQ������y)/�2h�xhq��}��'|+g�S�Ǳ��j:Q�}�_���m#.��-��% 5�T?5�]�ݰ|��G��z��E|j�?}��˦e�d������chr�jEw�yR�S�f߸�r��=vV�
]ެF�Le��k�������YD4�RW�b��Ż�}6{kj�)�+�t��La�LѨ��D��oC�����Ej�m���Rf=�(]S�ت)e�C�Wui��7`3E"i�{�^����f��=������0v�Q��6dF^�T�O��3Ro�R�wL ��쌂2<��'UȌ-�S �;�ts���F������L���-~J	{��+�i'j�	���E
�6�ƛۮ�L"oe���v^H�X|$򏘯t���I�����&}:�	�i�Y�V��w-ʷ�V�v���%�d�!�y�߄�'���nA/����NHppGj���d2h�6k&	ݾ��(��ƠlCל׺)�,+��p����f�Y��ϸ_�� к>�b�C�i�g~��䔝mݫt:��R�O����k��A<���w�^��I�Ƣ��h��1���W���wx�`�.�f��S�U�B��K�y�i���o��ׂKSH��3��4����5�Փo�s���}^���OV^-�QTͷ�Pc^�6�2F�=�Z~�o
�E;�nn��\�/)������^,����a�������歺T�J��T�W�?q�l�L�����8°��J���~k����rέ��>��
H"[���!�V�"�UsP~�/��bY[�H�0	��^,���
,��YA� 9���Ɓ{�z�a�;q^�����}z7;-=�,���m,�AfC8R��V�"��X�lo���YvY�+&���8�F���I.>�v�[7���09��7�W�Ժ̝�*���wmi�D�v�M��r�j��S]׎�����{��٢N�;�y���">5k�:y��B���Q���|GG�F�����9w*�AS���I�ů[z������]��T�cA%I����<����y��a)fژ��{%�(�4tEj�1+s_U��.�Z��� s���)R�,9�&
u=�O�x�R}��?�zx�_�����D*�P��M��CZ�Z���0�㐛���L��F-���^\�|:���	�����ˌ���o�Y����-S/C����^��~Um�O��bj�/��,��eOs�R*KᚚFb=�.y'c��~��s(��,z[i�:�@�\�9_de[]�u$�Lz*�{����,[�[x���M����3�����wU6e
��q���;k��ͯ��h��g�J`h'�`;^(��MP(���̃����}e��ـ,���$����D
���x4tOd~9M�>���_3� ��������i�!��&+����-�BC�beg�(ȡ�L8}Kk���[�m�
��=[���Kֆ*�Gq��6nh�P&Y�-�˸8��<����%�!��W�ק�D�l7L�)��۹��8��mZT�ݬ`��j��-?�;�pw5 : 냇�:hOR�ׯ�UK�����]�k���Or��sΖ���|,�Ǽ6�󷗙V�sB�9�M�FH5�O�S�iN���np1c��#Y}�HSvn�J���>�|>���R�ݡ_��|���osj���uú}̳B(wI.�
��A���j�g֟y��4ί���V��c��ۨK��qh�o{�mO~���u�k�֭0�qi�71U2H�3��X��(�D&�YG;k�j{��+�Z���1Q�r���RE	��M�E[V�#<����'�\�lEֻ?wN��^���C[P����c�VT\:�W!���฽����dՓ�.E@��e�j$m�2�uٯ��!�:��lb4)X�I�5.�ƯuEê��H�ޅEצv�}-�Oc:�U�4n;u=�fg`�Jnj~��=��N�#B�)�Bp<�#)I|�����@�F׌�W[��Цz�Hp��2��.�4��.��J�,c1W���"dp�67�������SJQ��;v�Y����W���-��j{*d���3l��c�s�\^Gt��U�xn1u���t�u�䰀�BŎu�t�Br���У�S	㒹��.Qz�b�-���U͋��f���t���M/��j� ����&��Ѯ�L���u����y��t�?0�xc4���h��vu�q�Em��vиa��r�r�R���we�=:f��	V5]�x���V}'&�k9�]��ݙB���x$�ě�V����A��&� _p��bZ�Z��@��$�u�=9Z��2 �YoD��[���a�$w�>�8����g7�z���n������ϬK�s���p�ksX�a1����X���nj�*���8������~��~J	{kU�OX�nj=�ᄄX4�x;:���b��=B*�=��ܞ`�]���R�L5�J�SlN?s�F MI��^��g&;��ǧ�5".v�d��¨��YXxZ��5�<G[�.a��͗m�v� �E�f<�<ze�A���$��s�ț���}��qX�J���1��(���DMǢ�m��f=������ ��o�P�O�r��ތ�v�jvTD[*Q6�ʽ����`L�"ˉ��I�UE��X݌n݃!���y���)�l��NҬuƣ7�`�C���I�5>S�uC���� �����au��_"wk���b�U_���ɾRK��ܹ��#!k�(A���+@*��z�b��;��������eZ��RV����el����Nr N=�%	ږ��D��&BeBѭ�Z|�yB�ǧu�k�=��Ӆ�F����M+�{��-q<�"}�^���y���Jb�|L9*L)�IP����^�G�������}�^�w�}}x��������������������߮�<O7��U
��DP��Þ<��LU��N�IAi�]����<ҵ�9ufM���zۄ���NP�[M"��],hJY��ph�"k�ao�k�>�7��Fs.��i̧���x%�]�-���{�]�:�ȵM%�(
W�i�{@jxV���y��.XeE�k)����68ҽv�r�����fP룠T�{`���(��vu���ՈL�+>*����A6��cCy��̔"�3t����Ś�ge�����:
DǊ�c�N�����\��;�Y�ei�!�˩s�a�MU������$V13�*�$���0�Dغ���\�a^v���9�=��W�;�
�����/q�rz��ő,�ڰ��/�e�9F�r�TD�x��	f��r:2�)��U�g17x^��#�Ί�gbD�}�q�z�k�fC�&%S���-Qkh�1���q�la����8�É:���NÙn�@�4iRy�2�d����v�;�)�S7*)m��h�	��̻�t�7��H{�:�+8�\M�w_R�A��g�a�ӺmK4�;t��"�V�*�YB�0�����ɣR��I�j��M��;M��9:���XYҝ)��>٘��\�2]<O1�Ӄp��T(�76:{�ʡ⎛�WMgc��u�K�J���]�j��!�9�}]����p�&���m�+Z�)a�ܽT&����h	��������nN����ݙ�Z���
U�&����TK}�������u,�T�j��w�j�Q�Fn���u��lix9ӊf��2J4]D�`'>G^�ֹ���7�8(F%�ʺ3�
�����:���(��u[	9�Џ-U��EVGK�T�JP��ܻp���X��_8/s�BT���oZ��r��hYh�� Gٵ������%֩Zm�ŵ2��Zl�tz.3JPXy,�yp�m���{����Ǳ`�u��qc�/���\'7�ҍ�w&x,�-H�o�]fn&�˦�[]��{��4
�N�;C�:�I*1C
S4[��̽T����`n��q�ݵ|t�w��9��X�Q���55�:�6�weҸ�f���U�ݑ[0���dÃ*��e`Km��@���K�R�iI4�Wp�a�6�Q��Pٱq4l�}����Y�0���Jԯ�hR����u\b�P��EAQ�@�JK����1?����<�ֺ�6+im-��EyU�
��G_*��y�����Q_<����9oc|>����tX�L�S$9X��Zi饥kT��N���ru��1nWY:�δմ���J�]�aL�:�{�;-�ك��ƅt��Ѵr�Y�va��c�'c5�<'P4GE��^bU�±t�ܘ�O,Y�8��
&�ak����r���Mh��֛���Ot'kХAD)��7@PERn�/l���A�ˤ<h�T tҠ�y��p���r��68�31LQHD	M�T�\�^ƪ��PP%%R%;���Q5L�T�	1T4E(S��Mm��)y��""*�mD<�`�
J�G 9P�T1@UD�-4��d�)�(�b"��(J��D�G6ZinY���jbb�����*"(�f��f.`̱�b�R��%��j)��$��"5��b(ZB��(j����U<�5H��Z�P�U�?����Z*$�&��HR�qPP�QM&�n�R�@hH�)h((F���*�5��34č��a��"f�������*�*"����4f"h���
jh�一���+�%R�QIDHS\�T�M%5MR5MEA��<��yx�v�E�:��w��.�TH�%���A�JeR~�.�%0őΔNF��N��z��į.q�%d��
�d�Z�`�(]Kկ�3&{�{�����	��-2ưUϾ�����C�hO�>W�	��1�7ƽ���bYU��U'���ד���������,s�+�w0����H0͒"�C)���!O��0��tQt�텵�3�ڢ���������]�i�Su5�^��)i�%�Ù4c�?`�9�c��eD�Y�`{��������ά����h�t�-W�Δ4J���'�Ut){�?˩h깪�P����m����s������i�`���YΪº�K sH/N3vC�B9�̘��VF�9��/;��~��dvg���2kXP'�s�J	{�T��n���銅�ɬ�����Yq�{l���e�P����(Xb��?5t�.�<v�U&6�:�lgӮK�^b}ȧ�ߔ#�
Q����T��*��&
�χ�����P�U���uLO�U��f�O�.�\�#=7H�`��ή�E����v��'$${8I��i­B��?�ܯ]�P	��1؞ݩ��";������U���q���n����"*����Y���`ǅ=0׏r~���>c>�%
��!�R���x'Rں���	�H�[��"��W�Z��+�E�*	�zpu1��N'�}��DT�4���z�~�Am탴��zk/�Ynuӗxt����'{I&���|ȼ7T�B�����>;5����%u��8>����Nn�y{^�]>��ӻ�����U�B�).��^ͧ�xmhg�X�ih���sg��mN�ε��0b�Pci��zཋi�U3m�2�QL%�!ϳg�=[�E��KSD�Z6w�f��B�0�CC�y��OT��	F��'���p�A��Z3I��.�����UWJ��JB��}�o^K�m]��&�f�;�Hyղ������'	�d^�d�d�"���u�s��ն!)Qk����d�U��	8�@�������`1�vI�a8ț�$�y'w�N�.��O9��)�$�5���j|��U��`[H���h	��Lp��7UC���s��������-Y%��)?1I���"��,9����#ϲ��	�|�]�	^��O�ս�aCjI���TCq�M��'�,�H�t$�H�0���ũ�qy��f�Y�e��v����10�B��y/�%e��c�gy�������-��e�tw='�q���3�{jp����ӿ�v��wo�>g`��(y��D;�S"u�	��]=W~v��I�Z�&ޛ����7Cc�����[!
!X���a��V�t(f�;�'�i<�Ѹ�dב(��5��L9s��3��F�H"eep����3��01�īU:O�3���t,���㑩;Uj� �y}W�L�;�E��ծghKH=�3�<��p̅k΋�j�~��MM�סs����:�?$N@�	hY�6�z�m|��hZ�Xv���k�h�}V�3�(��Ռm�����UsH/��!ݳ��(XXS���՚�"�^���؞���0�s��(����0$88J�;�-3��!�]z`Q��&��:����G�P�{jAdl���;�D�����@��I�^����n�-�&�U���V`x���MB�;�C$:-��0S�S���=�ٖhGt��*m�j�#.��Ԝ�CK]�.�/[���{/�yW<r"��@�B1�=ű/b���ך�zճ	]��] �-l�)��l�n�kkV�j�t,�2��-��4�Ճ'��	<��=0��ż���T Bz׊o%F��N�\f��	n��p�Y�A�֠2���
�7���"q�T���M�>�z4�/T��;u=Õ���[N��:輧Db4)\t�dvTQ�R�W�Ί� ��h���d\��<�,vW'�@ȼUx�<�\�]��.�HY)��?Ad���%:�$hZ�)8��^�a@�cE���ow�ڧ���"Ĳ9a��]߶��fR7�oI�}���g��Ý�(��DŮ�q��7UsY:���f��pM};�xT�W
���g|��;;,@z���.�Hx9��n�l�~��
S6m������1��@eŃ��n�E9�(Kq��m��>����:v�ȡ_&v�>�:gn]�kâuL�p��nq"�����g�k�x�d���n�Y�����4!�A~�&���ʽ�j�\�%=X&m��1��ZVp�5~8��o���=�Q�F�ꨛD�X�2k�����/)��ȓ��I�Q�\��w�t/c����׵�t�o^�:�z^�)�-�dG&�wMR�Tn>ߐ������T%�]PF��evilʉ�{ʲ�U�����֮����=΢������}njp��
�A
�5qѝ�Z~�:<�Xr��9�{�Kj���f��:��\���W�B�/s�,�/�>���&#�ݶ�	�Z�y�{���2־ИfY7��5����6�ֽ�a�v�5-�R[ç|�_}�8�[s��N՚rFwOj�C���P0Aam��6��u���;��PF$�x�f:�L˱M�Ι�8k	kܺ����8��2�QME�G��᭙��Uz'���{f�ާa2,�P�Hxuť�<�:�����]�`eIK�hzn�tM�2����	��Yq"3%'�UE��n����z��IWl��N4��{��=o>�>µ�_:,��݂޸�7?i����tx�T�	٠�޼Ti���6�:�=�L_y�����|G�cU�X�.b���d�:b��ފv�KndY�u�[Ʒy���nk0��
]�_8Y�ʬ�@��|a���B�aD��Z��\G0����o��[v��7����ݿ4KG��	Ҩo#^in���g�)�, Xt�O��h��Ꮾ�����9��z��	U-m]�B�tg��t-]
EI��ma�l*�-��3�Bkr%uM���.���C?g��?�G�p�������!)�ɐ�P�hR{�r����z�=[�T�������U�s;2d4(-!�<z��L
 ��CQ���	Lm�JuiI`��R)x]�Y�Q�}��7�s��vr�ye&bW�`�(j��`�yo�ӻ2K�b[��_ݣN�:k4H��z{���eQaA�/�S����� �i.#�Wд���?eN�m�T:ՊPů.���If9��E�L��`�gok%���ei���L��̚_(�{���L�O=�(�¥��]��Q�Ԅ�k��R�]/@�O̓�$ҡ��8���a\��B�g�v͋���o{�U��{����
ZTħ4:��&��k<ـ�W/Adw:�R;����Ӈ�pඊQ�ߝ�>&��o����(��9p�m.��E�����OJ׿b ��ו�3��l^>>��۳1DY,$z�?��nur7��+m�#���u�"��/�o떕Ȯ�3�q��_~^���6��޽q����M�0ڳ�fR�TȔ5��ƀٶ޷�\���O��p��̗O�&y��^;���]���;%*rZ�:�F*Pf'3
�	U���}��0�M����>}���X膄'vmt�Ͷ�}�GJ�>s~Oow�gӯ�D˼w�7\�\v�Pww�2�r͛�"�CG8f�	��>�5�W�WP	�Qڳ�ع�zF�Vڊ'������Z���Lߧ�	Ʀ��X�c]���L�;M��6�5ҩ�ڊn�%Ne��/G7y�)Q`�'��	�&���o�؊���x�!��c�쀪��=)�e�ݮ{ծ��}e����k�U�{����p���^�<�zj
��>�4�nb�š^y� ��4�FS���}C�J#:1�{�4ͷ�2��6�5$r��l�sC��_c�%aq�������y)H�x[Xm/b.==BUc�N�z{���L Ɉ�f��Hȱ/jc��N:�;�zi�c1���o�-��
>���\H$=�]#B�m~���9��������
��+�^oR��u�M2�J�]��{��r���& k s�D����ƀGCf�Fz���	_^or�t�'��.��	�]"�$�57Gd�6=C�q ���	K6�����+%n�NC��-�����o:X�OW<2\��;2����'�ލ�/��a,^��e���`a"O�n�)�rc��k'0��EP��f�ȃW�ĳj��!u�;��z����9��˘�X�Wj%����
��̚�*�OE�;�܊�[�o���Ycv�מ�gޥ.�M��q3�j�v/)�I��Ș��"2|�A��t��n���FpŘ����y��0Ct�J�y�@?��NBn������)	=iR:��`�h���+�Y|3Nn�t3�����00Y�8�xc�[]4�c�ʹ���/4�F���%��F�L�M7�A}�w�w��p�t�c��b��~4&D��݃����wJ�(-�ʻ�̟��:��RC�$������;�U�H���,#��^�k�L#j�ۆ��Mm�ֺcg74�u�˘$ĦZ���WG��sI~����!ۧs��C�>zH�˼�.[�ؐ���$��]�]�ݺZ��W�#<l���^��a@� �/<���>�Q9��`�L�{�1�N��shQ,��T�b��7?x�Dש��,ŤWa�x��.Z)�è��]M�p+:�Kj�ݺ�;������tŶӞ��̳B;��nS��A�T;Lj��|��FD5գ��x����o["���3�#G������WXݬi�	fb�w���=�4����T����}ʩ)�wFI�A���s����3�e��8E����5�j���c�X�o�uv�'�0��;�\w���H5b�^��}(M����x�&^3e�������ҥ��ޣ���sx>���Ī��ST�&"k\KI�v�>��7N�o�
�{_�'��,��e�;NP�`\脞ELf=��L�ci��-A�IV��.�5��z
��2F,'��hH�3��omr�i�6��%�T��F�]!�e�U۽U�{2ws��ֶ�sΜƆZ�	�N�b4)B�	m�2�>j#�ŀ��^_Q���8.�!y~�e�M��+���	����d���	�{a:��Kj=*�qw8ñ�f�<��t-���ݾ�[�h�֑�8�r�ۗn>��v�)�{���LU��E'�I�KEw��1-��I���N���]+�W�ȁt�
�>~�����!����&
z�e�n����E�u��oY��sٜ(��'r'��b���zZ�Cw=z^S�uo&�Zi1����W��������"�x�XJK�a�H1t�(F�����"Z���ΰ�Ik߳1�F��N�?��^5c�=����^�<lt?�0�te�������:s8��I>��~�pp�-hLe>8hZ�u�Y~��iA/maTs	=bu���D����=�j�~=M��׽@�8㛋;�ێ���wU�γyr����H�ȕA� ����=-2�᮶��R�b�_���t����{���3	��n���1$w�;�DN�U�a���W@-��N��Z�V��J�U1�2㷸����q��0�d��S�P���̭�����({8QH�����\�5F�;<�nɽ��Z�R�m?Mk�0�;@���@��:��wSJGF�f��\�
�.�<)��>!���,h���:�	g7.8�	D����c��e�ۓU:�4fݾ�쨈���q�þ�;�@���W���_Pٹ�G7��@�e��5ST�횢��CoH�#e�ͼ�C"L�O���Ui %eyU��S������e6��b�L&�����듛��
Q��}*�!��y��c��7C�:�{�,,2N6��3��|����{޵u���e����52���c ��H�V�k�#��	1P�^ئ~���`t�͆�J$�i����	���iw�a����KsP~"Se��	��"S���g�ј�.'j�%�t���[��l��Ŵ�8��S!#��Cv(�nBp��%%�f٦����*ˏI9x&�w�^��J�n�]'����c�pU0��G(�,h��^�锝	�������w��V���n��E1�y%I��Ds���O�_ZAvl�D&������%?������'|��7����5��,�����ӗ��\�
ȱ7_�5��Wiv,��j�Td7CZu�z�Pd���oش�m9�W���%.���<��z6��۴��
�ő����b�'^^�C�ݾ��֨��ۋ&�w��Ua�V�z̴���SW}��f�w���Es��E��T����NO���sǝ�!p͍"8Bn}:�:0'�{s�evrl�BZХ�(�*.�⮗��i��r�|@F�9j�]��{�ͻ���v>0�z�8��z�ƶQB3�?X��uJ`X���%Q�����x+��sӦ#��ۇ�-kZ�{�U|(�m��d!�)���������Ńj�[+2kXP'�sߒ�^��?2��I�.+bv�7�W4�ӛ=YZ���`�2F �Oc5"k�|i�c�+�3�ҩ1 '�O���&]35�T4�+�]�ݫկ|��.�fTb�o��Lg�`<�z!�[υ�S�~�fHf�Z��
�ٳw�ͽۙ�y��~,�^q	h�:"ص�!��D��XF���DJ�/�D�����~;=}��Ú�_����Pݬ`�=�Hz�ON�e�h��4�.����R�1�:s��H;��}�B�e�{nסj�%�f�i��L�^��èt��>�ٴ��O`ճ*�.�p�mٵ�p�n�gT#ZZ}�Ƴ��ʩ��н�iR�m�2���&�$r�� g���?�����^��������������{���w�����zy����[���X�}Q։׷��aB��l�m����c����/\�T�J丸���qG�o}�-�㲽�ə5�楧C7
���}��������J�ZkI��c<33Z�ձ|.�s��j)������ܯ�f�ޮ�ѵV��m텛
5������q��e�2h�V��*���.���1�N˼���(�/^ޘ͢�1�NZ�y^1Y8��S�K�pu:(�&�����CQ{�Uu4ܑv�I�)��,�J��&���7���Tod)���/2�mX��i�t�GiN���UG����T�� .�����ِ�*���b���*���1�Ґ��YK����FP3�Kk�d𳆻5�:�z�!Zs~S(�63��A�f�+������`�5�l��oo#��ҧbNZ�{�/D���3�$:����#1�X
��nb�e!��+���v%�OA��{Jy9dخ�5X�E���s���;/)�����Y�����&(��=V���Q��Z���N �%Јg>ʎI��P�zL��#;��os�D��˗�w�1�:(����1�nM(t�Oe�-2��mZX�
#$.^�.gdA�>߲���V���-�&Е.�Qf�]����%k<���W%��;8����x !���n*�W2�f�EZnmL��l����[�!J;��F��q+�<��l��AQ�)W�:ҷ�&��8�,ai����
�H;���ʲpPD��R��ȕYa�4g�%��H�NR��������f��\���N��~ �s�Ɯ�O|��/�xp���s�,c����Uf:ܐ��;�ȕՍ%Zst�5�N��,
|stB-����ct��:�r]���C���ē7����vɾ�7�h��<��)GFeE�4���Y��8����;u�S�]��/X��ƟeqUs�89�Y�õ3DYE��K(f'k"�޲��i�°e3&�1d��v�����>g�V�u��C�fG�z�K�M���b��&ޞ(#&x�m��(irkue�0�=��+����1UE�lN��i悞���vh�iRv��G;�e��].3��5nZ�e��9���ZvB<��iZT�m|�R�	�(�b�諳vɧ��Ǔ{[J��/.����4��_�O����G*pzU�V��=4��+O�5�؍�$*Ʊ7��oNCU��u��A�{�sܼ�ͷBt�=�Ѭ��V貟��b�]�pҾ�&)�p,���r���24b3�L�sr�VQ#�^�;p*��{�ޔW��k����z]qJ�N���-crBx�46�닇]F�Κ,�D�k��[a�WM�V-5Vc��_]і[zaXO=!��L6u�1R3�&qWɟ�K|�h��h�B#����
3eL�y�Qᚒe��s�"�/6�(�٥���d��S��p�9��Ǎ5KA$��44�P�D�%PP�$�UUIT��SAJPD�P�Q-D4P�A0�Q4��V�IAS%;f"��b�)h
��Zb�*����*�*��˪H����h�!"�"a����� ���
�;��D�LQ%-I3M)W6��C�B����j��(�9�& ���j��*���V������((v�QTE%4-45EIF�T@QE5EQQD�PDiMSM Rґ!�扪��H�������LB!AM5KB}��M!Tp�JEDF�D�Q%�hZB�()� �(��h�����CK�Z)ZJ���K�KlE%4ST�E$lm��RTQ)/��<��r�=y�3l<H��/�Wp�s|Y`��)E7cC#�t�t)�o�B�妔���m�������=����A���6r��/�ޭ�W�E;�amV����J�`�kϰw)��2�&l�I�f��R3��ͳ�]η]	*q�x�f=[ռ'�p1��/K�D,���,d-�X?+�α�.��~��Ng��=/)y���*U&��i`$��X�Ξ���$( ��e	�� SlCH���R��;���F�y@3I�>1)��t�eI*Lh��eu�+����C�*�2���^��������3r���NK�SfS��)?1I����-�Ú�Lav���z�=�r��z0��:��,G�Ϣ9�Lpm��<ԞΩ���BmNK�|A@�s��j�8¶M����ݻ[+X/W@}�l��5������]4�c9W5��ҋ��F����zTڞ�[ӽ�ܧ�R���/�tQ��C+�b���9T*F��C�����%�O���=.���.b�{V��J:M�_���U#+���7�hXCj���ڙ6�ϋ[�`�r��D���;�����8�$���Yk���� �sH/���!۵�5{C�9�����ds":b���z#Ϸjɮ��ov���w.%�,8h�ZQ� VP���f߉�ľ �|=�Ӷ�xq����w�ۦ"�	��"��Փ��������u��xl�o-={	ƕ��l"��,�#�)"����Si"�7���C�NY�qx���O}�>��غ�bT#�v�N�3L(��{]{��~=X|x�&�
��)�f�\.��ޜ�б�vDdm��j:��ڑ�ǺCs�;��Q3Eځ2�ZG.�N����,+��*��]���f`�_�%�.��4.<:N�b�)��z�}F���:�@��A���x
�h5x��qm������h���E;�d#5��Ⱦz�����cH�	}�Y��=����7��nm��&q��l�*�W(�)?�5��A�(j�IG�n�y7=�*o3[n��ve�Q�>��a�еY$f���@ʛ�7���("�I}�nP��2�B�u�_�g�w�����MC&=�!��/)��hR�T�S.�4���i��N*�P���>/��^��3!Cydt�S�����v�>�X�s�I��bS����#J�qw���FXZj�'��u��Ŭ��6-����!�'��2��v�׽=�.�Re���_�ȮvU��>K,p�rϿF��3������{ɑT��|�����rƆ�T2���Fa����=�Q�e��3c^�C�nkP�T[�Y����6�nºLkb j�b�79_�0wg�}��ઓ��n��=O�;%t6�9�r�$�8�\����`ļ�lsn),G���-�B�y��gu��"��=ɿE6>�"�=Cv�H���&����Zr3eg�յw����swx��f�������PJ��6��WE$�^,w��"�S������9ծ�q5R���{���f���V���������\�&wq�r�a�7��Ҽ��`Ko=CdiH��6�m�[��Nr4�s�8�v8��U���U��j��G4^�4���R?{rç�5�+4�Ͱ����_ZT�Ldnu68�F��zW=�����Q�$��֠9�ߣ[���4ݶ�����z��.��x�p�`=�ȇf7Y<�6��@�~�ױ�����ݴi��Ǿ�����k�}�%�Vp���v�n�����Q�h�����|Sn�&�♜���uw&l�@{�e�㸄��I��6Q�j9z�-:����t
�9��K�2�n��q��VμH��6�&]��i�O�23�`L�"ˇ�Iۖ)��ʙ�Qz�g�8aE��X���D۟����%ʨ�2R�4���֮��}hg�b9�� =S�d.�����Y����Hh�W��T�u�S�M-CR�����t��͊a�1P��?�e��B�IX��f��'��w�X�y�ٚD�{sj�wV�PX@�����hV��p�F�̳z�U�����wQ��ćk�G�`�-�Ԗ[�_<*#\�:�6�e��[�v����j�����{�C��_���9)O4��W�¤%��e�G80�2W;R�Gq�/��L�ѧ�T&���m�)��3(�j����J��[�z���x�Ɔ�:1���Z��#T���ا�������_�Ac۰�P����39�Ef�	T���Z�X��^I�CǊ!�$�����~7��.��N�����e��zaar�c�~/`.�e^IRaO�؄��C�6�k'�|GZ�Xv�O'��kk�:����~�d)���Ӧ�5(���KL��������e��2EFv�U�~�Q�	EMt��{ݸ6C�b�s�R����8����凹i޷�Y��A�A[ǵ��̎&+˜�'v���`���,�`���x.kjy�5?j�d�2�F���w:��{,�zh�ԯ�Z�9�Z�é����Ǩ�{���sL�R�BA9##&��;��t���t'+����l�3܋���C�t�����>��}�f���k���-�/��_J�ҩ�ة�l�{�]��v�,/k��u��z�y�3�N�f@X���]�VkT�<��~/���R���܆�QXGjۿ�9�X]��P��銶�y���N�f�@�v�nX�/s��|��f�J��B�em
��{��v�|���(�^!��T�tKBf�r���3�=�1{�ik�g�暹�X5����V��� ��w�]���{j�JJ�<zZ|;�����h�a�p�e�;˼��1_~�	�m�R���*��3H�ف�ƹ�TKzC�ɶǺ	Hpx���-�#b*��M3�d"����Ϋա�!���cϝQx�[y���ff��è���r��'ױiw.�ui�u�+�yTs�P���X�ii(�4�F���s��[N����B���&5n,�SO��r��]
�<{b�H�tSǟk���.��EǦ=2��s�^�DJl��f����=]�9�Kkix�D��z3���=S�L��%t��d67�/���8�̹�54*6m`;��ح���\W��d]#��T*�v>5{gO"�u�N�����t[��{+�>�}�0�)4�%d�z�$��%:���eI*Mmb;$H싇\�����&9�T��b����W�Z9h��x������@q�t�TTXsQ1���#$�u��,�����ӌ����G��DsmLw�l��_�D3�r�:&-9Y�R9� ޏW������e~�����_=yw�-�r0����{Z�X�ES�{�#ۇ8@q൳���5�*T��-�ڦ(S��ߵ�?h7U��C���dDC�Ǹ*�'.��,ꨡƝ�
�ԆZ7�f�+K/^�j�x&ix�����.'�tw���L�]<�5���oPr��(a���2�gb3s-}]4�yʅQ�\�'G\wr����G�7�{��u�t��0�#�N��!���.��9��k�1�t��*�M�6a�&��<yƧjCz�qaoN'�W>��^طvlip�}aDo=v.��l��ڎ�QY�{��uK_�Z�lXu�e�OG����SFO��_M�h�q� _���s��]׹��2���z�^Q��3�����-?M0�D�LW1n�-�c �޲/߼����ȷ7s�?T�`�+�"�C�v�^��S��h�&l��کR���#=�������<���f�h.�^��|���+�P��^�~5�k2>}Y>�v�;��n���USOH���XF�:��P==ЌV}�~�O���k��ol��UϪ�&ٻ�n��o2�hÍw�g;�h��� �pd�W(5$d4��m�{�=�'�z�`E�I��邓b�����4��wt��%E[W���ֱ��=Y����#X�_���R�q�6��g��s�����,c��ڹ� *Ro�˂�P�0m�q^V�,��n~�l�݌�|e�o�Gs����>uS�gX�}5�lu}�9���O)��IG aP����1)�� �m��V^�b�&�s0H#)i����bѼ��f|A]#�\z��u\�8���P��2凖��OR)h����*�?��Qt��~�ݬ@e�vyv��q�W�`�Ǫ:Pe�dϥ1�(Х
K	m�=�����R�ǚ�����sQgZ!7�t)@Lo;N��[�_�2/nbS�H�U
Rq}3P�.�d��Q�[B��􆶤�C)ۗn"��Hҩ2�0�b.4*6�n��=�j�{��26+W��L�Lp�IQf��?T�#_��2�v�����<�%t�[6��η6]b����W�-/B�Ǧ��$��u*`=�@��=�t&���U%=�q�ז�0���\���(��('dvt��	2�v��1�B�n.�����5i�Y�M�O Z)Լ�T:��;Q*y���cI]k	���<c����f-�o�0���|����:)�������"��bN��zW=������9��z��_fޫ�p��Łk�D^����+#��既����3�%�*��2���`��)��5�h����vJ5��ƛ������������t^�9��0k	��a7^X�=�ǩ�Quӵ�����9�ax.ȯ�+A ������s�cW���s`��u4𫊕�5b�#z��{`�ꔩP���5n���(�OK
y�q�q#��@ê�=�<�074�s�;K�0���>�_�w�Ә�ٲ+��ibR�e�0�o��+�J��U��U��n,&�q�OY��\wv��ڡ���2$�-�tg/��{�B�@��^a�=����dZ1��vFT��:�ww��R���ݐ�?'6��#��*9`S��p~�0=�\|�����S��u�ʋ/mgc@̎!��	r�9�M�ۦ��#^Y��߈4o]�K�X�֕Y��N ���p�]�c�T	5�R��4�^���Z�
����{Ռ7^;�?H�-tb�1�^h��ӛ���yg��XPZT��%�j1��ږ;��f)�ɐ�U�B���g��~U���z����o���X�P��$[&�`DDΫ�^�S�A�	Me��S(nL̰�s�������)LW�"�]���1�k�:y��}cXN�>C�$�;���m1�o6k7�W���.�1�d���Tp&�؆��	�G+��d�+#��Ӊg)���3�Ser�ة4�j9�tRt��] �ʖ��jV�j�w�1�Kl���9�fEV�X{�`�Ȃ�@`�An��B��pmFˢb��ZPX�\�#�~�*��{<|�oq6���D�b���*��3B���`Yz��DWj3P]{����jt���`I��NP]M�P��g++��+f�fy��QX�,�Qj�*�4���Qzf2�ǆ�G���o[��.X��cz�94gs;�7� �F�����7A�K����ӏ�|���z����w��b9��sm�[B�Re���R����� �:LZb�
��ݥYH[*zp���#X)a����zb[̉e��l;�J�h��#f:���;Q��yu��r%�\/�<�_B5jWAY,`��T|ѯ�񖉺Q~���{�kK*T�ky�en��W��O����u���,�9�r�5 ��,c	��#��dz��]���«{�n�n���JC1�;'����`��0� ��g����u�v�kü�NeF'�0�(KU�yx��g��6���D��=��b�N����;H�C׆��<���i/���툁S�,U�g����k���'On�g���X1� C��~�s��{;��2��,:���[Ӯ�d��me����Y�k��Vn/�6
��,~�ơ�~>�������J��Y���e�.8��n����}}]ʘc/Zeg�.6s��=����{�zj�l��NO�GJqZ���E{�V���L��ܾ�[��FHd֞��l=�V�o����<��r,D�� ���x�b�ܱD�V��4X�M�y�@?Feʏ?+:�{�u�S�f":��2���q'Z�V�%��[$w�y
�t!م���<�h���I]lS�\8�������,��0F�6%�����9ܭ;\�C���a"�XM����нnt����=��������W5�A8�bY���+�
O����l��S��"h�vҨ��j�ˬ�ě�Y.�(L[ v4�'�O=y�$���IԨ֘rJ魯��"Gd\:;Y͌na�������wo���y`�>�3;`nʇ`��W�@�WI;LR�)PJ����"3;���:�UY8�4�ul��l:ض���	����=��JT_C0<��-�<��'L�M+1ʘr�Oh�ou�!��������w8~����Q�50G8�C�+z��M7g)��N�7�|�c.�z��j���e�~��ʒRF��#Å1pB�P�1--�/r���]�x�B5���2v��ه�y	���S�����So��"
cH��aD?S��������n�fˎM�2�K�#�E-1%�}e�NǤ��i~�����!�ga�$zxtRೖn2����}n/R�ϒ/U��I�����W��1\��{�tɔ�Y��9�7wuuf�Hp��r�,p�o|��T��ݙ�~s���ǢK�f,@�}^�_���^>���������������_=>>�9s�n_��5�l���Ϙ�}R1�F�Z׮�
��^]p�WV���g?K�Ͳ��[��2�)*���R���Xv�IrWm,̱��b�Ռκ�v���	}��i̡�_tj�X��u���V�lN)����b�4���S=�2�%��gV���q��[;�LP/-&�=o�g��7�e� $;���X�+�=��AU�Q��"b���f!tӵx�_;�U���yc�4�n�	��y'vu�$����z.��j����M*n8�7�k,��}�;�_hg����4z�����k^�Ws%�R �1cn7��YD��l���N>x]եQBĒ�R��oXuy��rۣԾb���im�d�c�����X��S)k_d���ޭ��ɬ�\�*���ܥ%��H���2�`��/]W"<��B�T�Q�l�&u���I�^�v�
�Hx�ӧ��fᷴ1��D�A���;3.bY)���ZB��Wj=�!AY;��C��f��^'Y����s��$l�tE�0'*N��Jlzi����Z�����b������Z�l�1�*]���Jh�B�_`M������</
Z����l�ӨZ��eի��r��� ���;�����G1-����%���5��7ɓ�c���q�kͦV߶H�jM`�7�;����ƒ3��u�<_��7�ꩺ�u���]����*��18���7�W�ݭ]�n�F^W��Axr����|���Q�k^]��ڎk�@�
�É5L��f9�nN��Y�V+��s��A[6�����l�ywRJ�9�X+G��&�<w������S��$6znuа1�u&X�8pI��M��$p�q��tY���L����gz���#�كT�A{O�����٩�k�z�黢�>-���
�rLv�]���<^�і.'�77�x�2����#\���CI����n����{.exr^�Y�7B&pٕ2bojW4�R���ʢ2�D�O�O�㋭�5�;�j��:�EܾWYN:k3tH�X�+X���&j:}��un����o����}׈k��
�4���bU��Q5��uPU�!n�S��)2�ޫL�4S���[o�j.
Z�w��Ys;�Mm�#M�2;�u���-��\  ����$�Ү��N�����)�*��&�K�:h�u�w���A����[�p�԰<��͓3�X;�+����M��u<��R�sT�b�ڃ���G�SR7Eu����7.�S!줵��
it�����ګ�R�r�e��,NJ*���t����n)��}�G��]�x����JJy��H��W�e����/��
�ryNP�b:,Y�� 
Jk�q(�Ws�|z�W�a�7[e&���4��F�4� �!`FT�ѱW:�R�a�Q��$�6LM�{Ai�Mp�T�$�~D���A��I�^�9TT1�(�"4��,�
�s#a-G,ѡR�����B��z <$���[%�,AT�QIMCM1QLQ-@PKV٪ij �ZZF!�f������
j ����H�H���H�h"F!(������X�
J
B*F�Z
�bJ
&
j��&���fi���*�*�� b���Zb�h�$��4QM%U!A@D!DT�U,T�LRSEU4$EQ�&�V�����$)*�I"�(h��"��j�

��)J�q5CKC�h��4mj���IE"QKr0�TS�V���"�J��(�(�uAAC�1Th�CQKE%!T�RE��l��<s�}>}����^�~4�M�Xy�sл)tb�Q3]���eD�v>�m�gHE����r�kd��:�q���lo�& �C�ЃP�$�M���ݻ�H����x?R�%m���B8(y���Q1m�����f�o�"�Z�֮����;�ˌ�I�l��=sͼ��X2�5B-�zc'[�Uϩ�X�6��ޮM4N�����Xʔo}1b�mH�0=q�؄�ʱJO�X~�P���s|�^O]����f�9Iz`���*�9m��|n�'�j��$k��;\?S	���3p��hi��=z����B��\L<k��3�͐�_��Z�dE�B��J��{'q�6@�Z���s��t_�9>XS2.fv܁^�۴�ڟ�2/~s�ZF���a�m]���ڵ�yn�ڵ��ߢ�!�Ы���� �؆Gn]�5�@��T�:QpӚi�e�wV���Ͷ�)�D�A��<�v��1�8�!�~��G<���p��a;��Wmw�����Cs��U<^��S"�<1�^�#r'����R_:��2�������KQ~̐�����-j�УcG%s�W�˔]',J�P�BxI|XMR �?/����թ���}V~�8;v)��K� `v�.�7_0����4o΅Ц�}�����,����	���ܛS�e��6(>PG�N�%:U�$�nH�Z)L��Ջ.��Uw�A�ھ��| �7�C�U���Yg"NL�"�T���zmG<�#���sT��>�ٓh'�d닰J�ΞeVְ����E���'sx��w��A�,Mr:a:5�	��3)�4-_�I�	�\���֪9�����Zkg��x�Myh�ɧ6:�R�Yj@(!��J�o
�y�{�Y\�5v�@�~��gڦy�vvnB��޼��"�{KkP�{�F-A����k	�a�7^K��d�(��fPч��r����nޭ���LJ$�x�f:��f
����g�Z�$�a�
�"�x�U�a+��.�������R݉u;�fM������}�˴��f��E<7V@fp0'��V&�I;��z����e��\v�x�^=���Ɯ�D<5_A.UF���B5�\m�j�L\=��x�b�=���YۦY�B�k�w4��OW�*Zڀҧ�k�A�WA�:�R�Be�����g�0���}S��g�8��c���q�1F2V'jXOq�+�	��;\�3���l��ή�#qВ��ј�-��i�����'�1 �:�W���ҧ�����,��F3Kh�.���7��)+$g��CB������q�m�iB�d޺}Q*��5��(�F�SA�vi�x
|Mء�-�ٜfNv �ޫsKm��':)ä{�\����/+R寘�{|��/x�Y7�r��̣7�ls����{~I�i�Ғ�N�q����7��:�(,IP�6s�+�+�@#҈|C�
�!���˲�\�.2+j�/&q�Y�"t��ɔ�c�E�.�eI*L(�p�Q	�����2�ψ���51�Y����p��C4�7ҝ�wEL-�]ctS*M��0mx�/�bW'˶�~4طkN�d0T3��cC��gs�R�4���@��b��ZQ ���T?4F��E��4���ƽ��ڋ���d/�?y�����C�l<'[1�9�v��d�2�dk)f�p�̗@w�j�+�f�wt�u�!8�_1��A] �pvF@#��+e"O�:��m�Ȗ]`��:ܮ������R�tq�x���}�����{�j���m\
ьh9�k����/u_����&�F������d�/l�@�j}�gӯ����&����(�q�;Uu+.����V���n͞\�Υغ��C6K[=p�^}��A�.g}�1��wЌ��M*�OS�ջ4|�R!m�\]e��0�ν��o�z����1��s��wùs#�T5�����׼~�����M;��
����ʓ��0S@nZvS�;�upQ~w,����w�X�l����=��|�7:���[�
��T�sXj֦&����n�#kwm�k��ni܈�gv�C��/r���b�q*ȪGCn�z�˨/�F~F�y�M������O���t��'�:����}���a�h��,:�WA	7륵����S��|��/Q�N�)�Y�X�ii ��ӛw^�{̋iԕ3u��.���՚���f�3Z��M��$܇�����l�K���a�y��Lg�D`}�]G]=f\��V�m����^��9���ÈC]�$gWtfP�W��@?~�ʥԥb�RZ=�6��#XN�����׭t�C%V���x��Ĳ/i�W)P�
;��<��������I}�|���m^@\:��N׬S)�P�i$�<���L�ۘ���L$S*%Iy��^�Ej	��뼳��p���1%f3/B�z�>��w��T���i.!��1@����4�srN>�-�=Z����9��<��B=Ȅ�Bc�l��#=F;TCp9�^�q���'���p������k̤sO����M0�p��"�a(֘r9ó�׽��n��wkV��(�$�ڼ��&��HLe�%����"}Q.� dS;x!�6�:�����c�P	SF�չ��*�*�v6�*�F-Q|3`�\�'p�ry	R��w�;�[qs[;�f8b6�ͼ�:\��G�����T�
M���y�ˆ���u':Uh��D�|�W۽���0�ށ`�P(��Jf�#���V>���t�q��ҥ�7���wO�q�^���ypB�|?}="�WI�k���I� ���Ҩ� j���{��]�9���LlUh�W�,�9eM
���]�$L+����:��$��Ϭ�����fu�}�����;iNNÕc,�t�i�L�B�s&�[KץؾH�46�l�������3
&o�F�v3L�{�9Ս�w=��}X���Hv&W���0}垪��+����s����4s=Z[7c:�uw&leJ�@<��/l�;"]������s��-�: ��d*P3rH�/�|��=��x�/�˵%!�^��㝟'���>����mR��0"����L�Q5��Q���>�1L�{C��C��)�Rr���ٶ\���K��0�w���4�d����l�PW[�^��zap;��i�T$�׆OV�K.�{�_{"�����ӺӋIK1x�v�H��|1�)������<f��z���]�d�eV�G��Ң���yƇӸ�:O^U���9��W|�������{g�!ހ�ȸt�������C�&E��Jt��w��G?A��N�AN棆�	�4.�I+	��vM7�|�K�jY�%)���v_}�t��4�r!p������¬Ϝ�};u\�e�#�����lVӼ:wI�0^R�m+��q��˹��+:��k��*^ɒR"tG;�����9�_�/��o�k��E�t����(� ��.����4��H�KY�=���˞�Ǎn�E"܃�X��=x$M
�|��O/ِ  Dc;%��#���ZUL������ܢ��x\�G�q�Ԥ-/�z{�R�����Ϟ�=�e'��������Y������>7Hג�:]'n��a�4F^l��������C	0q5L�� �eP��
���4�vA�]\����q��k�j���`a0z�0N×H�Ÿeh0r�?�i=԰��:sQ����s��}�h�3�ٷ�al1Pp�&��ԍ�L<��;7�6d��rl����{�|�W���8� �l:�ݘƄ�Ԛ����2�At*���{%���'��&I$�>�t[xϺ��C?��u�X㦍t�R'�l韫�����;@̶��9$q- �ח�d o���_{�����v�KU����gs����{���)NS�V��8,bĲ�͕������}�������S����#¨U_R�xy-*�+/�Ř4���$K��xҋ&���u8�+�9&(�3ӅɽX�O�.a�z���ڔ��6����I�y�?x�_G�7?f�Fa!�WO�r�7�M7����c1�n�
<���ru���c�l3��@�w&�39qR1"�
	yzW���>e�fy���t�vl��sO��:�����X�FD{UI��4KNW���5\o�+7�f�FMz	�n榜Ϫ��7�0��/o��ct�?�o޴���Ğ{��Syy�GO�A4	�UO�r6�@�ht�1N�����Z�l�a��b��HIdq���������s<m���L6I�)Æ�}�������~�- di4Q�m�os7t�볫��4f9���Ӊ�78����#{dΒq>�[�^5�\�^�>f輞�-}ь���ٺ�1����k��aJ<��p�b�{'���x?BG����C��pR��yȤ.GPl��k�����ކ�-�xlS�+��?�kJl�"���ۗ�Foq��6ّ���᧝Y3h�*%3.nu
������2��&f�S��&���F �%� lx���IP�,�.Nѫ��B9����8�.���6\���K��d�����n6��]0`���-����3�ۓ���vs0�Wu��?����&��O0�~�O��`G9c�1談n�<�f��]�ۢ6;��0zK��<gh�W��P}���,s.��[l�������{���y���G�����d��(&6p���S�����U�cb��۬hJ�v����%C5�e���A �l���f�1��8wv���ԅE>��g��
���J�M��p.臑�ǲ�����P7b&�#}�]�`�-��o�.�%�X��5R5鞞��-â���WsY�Z��ގ�N�2M%Ii����P5acc��V��l���{a�Ȟ����2x{}rG�̸�6(2
��L�>2z�kۻ��w�[�)C�ݺf����
3�W���ϵ[�r�U��A�f�-�9��0�R#H�n;HmH߬?I'�	%Y�����U�����fmjT�1��!V��X5�KJ1Khf��)����}t� A[L���a¶��@��K�v�=R��л���I,<s����J��)����T��vի6賋m�,b�O�ΗM�.w��bE��t	2���m;8����2�"�΅qfC�m���4��-��*�`�M
D�R	UWi!����&vl�9�`C���:��w�� �:��Kj��h��q���9".q�0�G>^�v���0��2ُ�H!p17���pdm�N�dԙ�1Z�����yج��\T2��-/���v�B�r7�����b��mS����{��$��3E�t�u�f�]�c�`����ǺCء�񴍅��(X��/o��=��~���_#��S��&hҀj�}��<���(e5L�u�w{���-��>�ѕ��c��5i$Ɍ#��v��P�{Rot���͝[[^��}>z�x��Y.ei��K��Tci�1��A��Ι�����(�g��,�g9�`NΫ��Vp�9d��W~�����w=�y�L�^^7@� ��)4 �Q��1�q)�����)ثJ]�59��梉��\n�{����ȍ�DF�n[K�����B@oO���T�%�b��zw6M5n	�7�s�՗���5ɞ��Ե�{c�>c4�ܦD�z�a��r"�����#n�P�?]����2s�2L�m]��t)���Qb���f1Ϻ�Ӹ���Wux�w.١���9�)��P���q��c�8���C�;;�ezw�Tɫ����EX,�W�*��RDE�d�V�zZ���*	�\D����xWG�
�T&{٦�b簬�_��4T-�G+�z�޷w
n�"�n���
g!\X�^�
Ѭ���B�Q�
=~�;�]� I|����rs��jߍK��۽V���٧��t)��H@�^�]����0�Y��+��N�f�aݚ��äi%�=����p�VdH�!r �l�$�lp�k�-�Lz*���Vn�N�os�E_��JD����Ndf8@��K�m�G�+c��r�m��et
2T�Y� u�G����Ԗ������;	k(ɼ��;���w�x{ɯ=��7֫��3���b�7(�]�K�
u�|���kڌwV���Y)�v2�YT��>9�Uܹ,�R�0̈́Q�4��E�5^#�]YTfX8{`�@1@5������9 ��������^�o�������������������������������ϱ��Z�EϬ��3d��Fi���t�fk��oT7{����n9��o$�g��e.�|���iJ�v�HܱTR�+�Z��$l����L����7���W\���N�,�o��Ò!Om��n����EFuMշYY�ۢ�*��H纘x�9�[�ˣ�*P('7�e�=㛒L�<���O�ЕD�P֋��ۓ�ut����T�r��V1r�NN��s�'�q���um�-S������-
�W�C1�&J��]`�PYZ���m�%��1�9m^)�"V��r�h�fbm*�[}U]�u�QMc�
*�\-���Ixk������=�����u�#Hm���68U�]Gxx������C�2��\RZ��0�����-���>�#v��B.��:e)f��Ph΃�nF�.3h]���-�G3������0RG���m�@�����A2x�p���ݹ���RE���+t۾4���7��կP�W>I�E�nW7���Y��3;qO�>���g_�I��SB�Р9�Ъ�����haĈ��q���d�QzVU��l| �Ż\۳W�BQ�Ϋ�mSL8����X10r��ܧ�b��"��ơ1:2��^\���W��k�E�e����*������QY&w�FR91���w(��r�N3B�xѾ�O	��)`�ۓ�p̛�j�A9XX�Nu�Jr=A���]��+��"5�i�c8�);6Bk�����X��VQ�d|9ۀ= ����������#�����Ч;&F3��(�8�X��+dJ�fӓ�� �ڴJ���GD��b��ZI�:����ð��X��IngJ�(�tvU:nv>��n�n�C*��R������[XW4H�x��:u�5���%<�)u�j����{4-9�� �o��ri:���W���$泅�kep
�.`w�����:����롲=��[n�O�1r*KXYwT�e��ڨ��ޭ�q`���nJ��|��!�Y��s6rK�ݬ˝/g��Zr��9����n5�%�f�y��[��S4�63��J�{*ª� �:�ycE6�UkJ>Seq�)7�R�/�T��Ps�I��l^-�LY�_-��;,G7��t�'�KN��h��iRJ�S����!�ޮ�lE�)7]˒��A��9yɮWe¨Ŭ"��n7-��u�UN�R�e�N�u�LyW�!EQ;�CgFw���f���&G��p�ւzd����*Y2�cz-�]��:�s	H.ƓW7=�U���t�+�W��`�۷����l�fs
�L�6ˉ�	��B��vl�6�W^r�0�u�ٵ�$�ᘈ����őS6W�z�qMϮ5'�D).ӓ�)s̓5-�sZ�)��L��bk���*e�n]ۜSs�Ō�]6��U�y��������QKM%%����* ������@EE�>܇�Cl.d�)���h������"hh�-h����,CIH%USF 4��ӣAA@��1Tֳ4SEDMi4L�DQlj�""����sf���*(�����*����d��KTPέ�����l�1A4IZ�[f�����-UEQ����("(��9�4�ĴHG�4R�ruwj9��*�(*���cQSQĔ%Fڈ��`�JR�H�B$�*(�Jv�A��h5MP�ETQ!A���w���wߟ�Էk5O�=B_"�+��ZNf.��������f;�Xe7"*�[n�0��.7}/#3l�}��]�c����sކ$g��>x$����3��|į��,?�a�+����5���M�ޫO��{/�s9@�d��>�(�Ԩ2��l�x����f�_ೣ������2���$כ��ϻt�M��j�֎Q7&t5���YOg�v�^d���b��Iʑ#M����{՞c���|���5��V,���nf�`�P����� l��^�G�/Ȉ�|K��w�q)�y)�lz<��N���m����6�2�r���M�t���Ċ��\=B':9��=c?e8|�I��>5�#C� �ߴM�"��U���q.��:f麔]�;��3�A�͓�ѣl��*�hʨF���D��V�7 ,��P�"C�l�5d2�9�k��^�K� �:�O%BUO�s��@�� u�ܭ�/q�z�?D��\1Gm�X��>�0��gĒ����о�������0���r�Dŧ��c@ܨ��G�*�iύ�gT���o.��/H���&g2�8�N�H;�M���*c1HS}�,h���f�2�X����:�!�oW6{�r�j�|p��TLpY�*檜��ZGk/HZ��'������J�F���jS�6	W�Xo�<%���wn��b����`������m��j8��R Yۺ����3)u���oU��6�j�G���Dl�9t��&������:�����w];Pw�7�����9�S��~a]��5������O�w�_�~���2��}3��FfzzH�wg��I��4l3�7��7����#������tC��7��ꧺH+�"jT�L����g|��pF{��3���v'���TP�Uжy��;��=��@���9�?;U��0ו-&�]b�lte@ga���+��z�~��p�Iq=@���)��iJg,c�����}��7�D�P��-
���Yf��,���A �Wս��s�P`���h�) b��Cj`΅�V�鼣~�qwD=��\��ּ�r	��쵨q����� S���c�N�Hצzy�ޏ?��M�H�;�`�����7/K2�ܲr�w	/�PW��7VL�l0�����^���x;.�'�A�^�����z�����5��Ji�%� TǺ1�]��ͺ���3�)u��v73;a-����y�J��^(j#�X��k���H���v�i�&�Ѻ��0jŁ�T,W�����kj���!�z}�Q�+�l��|��6m,�����r0$�,�Ҿ�v���Y�fs�J�����D,�J
iA�z�ٓsNk�%���#v��g^����իʲgF�V�(ג2�B3'n�[���v�Ɏ�ξ��ٹ�W>!������S����Géq�t^%R�����T��v�]s�w��bO��]9�O� �y���
r[T��Y&����F��k������}��u��܀�u�Fc�ۄ�B�ýݎV�\�"a85&��x��H�~?y{��Y+�Xo^��=����[NF��;�n�n��l����T�����Y�>�qI��K�v>a��AДȃ�NJ� =����X���_7�3�F?�:\�{��*B�oi�KVH�a(�T�e�v��zz�E�Q�a(��썽�]z�}[��Ͼ{<|�|c�]��~�q�7p��"��!�`���HǝZ��l�9��V*m�X�R[u_9��/����U� ��k(tWGv٤���]�����IQ�6���{:�^Ds�j��E���@�㪀��яR}$���e�S+���XP�L2�p}���efq݃Y\>�U��!�dP~�h@YZsb]E�T��{���n�%y��'g������E�G������s��to\-4���ީ�~�R�%�zX�C: `�gI۝�C��λ��6{4���͘�8TxfYy�$IDG�K�y��9�z+/3bol���x:8�9���I��T�]P�i�#�eg�R�/4�{u#U��܈i�-���*�f��Y۰�H��ƪ�bf�P��ҕ���
H�[���a_:�~�c]}�s*�zf%��!���`�]���j�}�{H�	GbD��L�χw/OYb{�:�wDY�*�]�K��z���k����P9�0j�8q�K���ZH��O�l��N�o䐷!(��{�WMM��̣�G}�#�_ٺ�y�x7|���*R&Cml5;��p�~oo�ؕ>D*1�Mc�F6޺���J�Y�q���ۛ�o/m��<(h�Dц���%�u�$����
֬�y������F��C`�u+-I�跍n'xѼ3�sav2���J���8^5�4�_v��-ܲ�d�h��@�=d��Yۖ��XJ�v'��%Q�\l6�!i}����/e�������D޾�ӡ�)����1��I���>7H�\|kϥ�KI~|�w��lȈ6��Wn׷X���,2���B]�9�Uܹ,�S���l���0�Ec^w8��Tt�q�����
��[g=H���W�m�t�Y�T1�W}�*�v2��ut��:��o�s�n10T/^C,�ʁ����6B�;��;�լE���$wF�i�G=��(|�]���.����;u��ti�1V�/yW��$��Lv	�4����gȡM:����aC�;J|W�,q������8\�${���č �Z4MiQ+j/%�ƃ��*��g]�WN��LyZ���f��v��Eq����jmU>�uEE፭����
6�L��C?�_@%{�539qR1"��}�p3����@��Vom�k�WA;'IY/{�Eb#"�vn]\�k�鱶���U��)�Ԇi�����H����M���%P㮱�|�2���2���{S�X*a	�[4$�2���)[H�,N�t����_|�\�r���h��z�q��w��'bޫ��l��Q.w�,�M`��X�D��-[���o������DIW�U�F���Tә�[:�E�=�%pL3���&gw�N�.Vy
��d1���h�I�S�>�φ�(��LX��k	��ٽ!R�YalF���һ�`e�-�Q�IT�ȓ��7QLw�M�����עu��*Wlp�-�eq�c�FWt����S7|���evao%�k5J;pY>��:M���ئ}a1O4��}�[��ݛ��ibEr~�g����W��l;�>�����V�����\���]�wlʲLH7�$� ] ���j�`8��$�:g�����%ov��M�F��C��H���T�tȹ�O�7�GR=����2�4b�����!�G�ڨPWo_��=�vy�e�t���#�ϧ���,\W��g	L�ʅWR�M(ԩ�e��='H=�;%:���*i��Vѕ2La�K�k
���VJ��g�3�{7P[t7��]MU&�H��8��]؉�Se��r.�Veó/awq�g*VZ��)�7/0�Us�款���چi��K7�P�A�TCC;ā�Y"�gw���!bY�c�9�0�a|�n#���ò{�e�h�4+������^��5A�ݜ�Q��
��%�3�,�q!�O\����:
-�|3o���YOy�ݢ��S��gG�=º�H�d��r��F9��;20�=��ف��R��(r5�l�cb��l��c�R6ZVɓvë�dԱ����9{��z��w'��oI.�����G�Y��nq�!�c+)�t���	���R�������R(��Pdz����\ӗ��=��y�3��(v��
�3�m:�T-��
&�rF�E�����i��͝��D��ʻ�NU[85ӑS���w�v.�ԍ�%�In���3�%��T���������̷P_�;#ݔ�@���a��l{)�O�y�-�fe�w�5<<Whl]W�O]��{���O�7��Nl��x�p�B��H��=�v�Y��Wݴ�N�{ONw�&����
�B
��Bt4����Z�rW^��q6m΅u�əC�	Y�p�ʌё4f�Dj뫉��JT�$ҹ�M
8,�e���/b���a�y�S�u��|��1L�m\�QAj_l��o��.P��6��񕦃9���T���\��=VV'9����6�� 
�顳Ro�oZ؞���K�B�x.��[\�f�.6��,5�;/N���a���9�Ok�O��T��M@T�t���	�Ӿ�n�ˌ����Oe�n�~�C�PF����Y^���=E�mx���;��������	�� O���u��7����?b4 'l���.�wN���u�-��ݚ������g$c(X¨r �������̞��[��q�zV�1�k��|]�����t�6�)$�g��d3��p_!���}�ӿ�?�	�_^�D��	z������w�`�_���W\�y��wʷ��E�{��UO�̸�H���T�������)�d�kDN��M��.r���8k`�	�����=B2+RW~�#��R�����L�gMMlfa����O/?J�u9�p�w ��t���K!�f��~4�~Y�y×�.\�(�WMY�v���A��R({��]r��#�ɪ��dy�~"���>)�ˣȍ]=Wd���L�&���o��p)(#,����t>S�6�.��6+�ϲΣϣ�������k����X�;�h�J�����V:�؜'p���c�/�4�b��'�4�������А��"pM�>4�x���k(��7�ݲ|ܸ�].H�I���r�vfH�I3!긵33Dt<qDa����E���rE��6vک��0�3�l �ݦ�s}����m���B�/g���j{��{�J=�mJB��'��*2�|uU^c7m{��N>a��	t� ��u����	]�-��7H�]��q���V늖�8�3����^;�v��>&��`t��=�A8s������(�5%�����ȡrHw�]��-	�-}c,f�vt�b��i:�ɩ��{^���W}�˪n�{d�'h�J�q�}M����x9���~��x���1�G=�$�tHd�'J)�-x�d���� l1�Cp-ޯ?������I]� `�<���e
;�B�U��v��R�n���j_��"����,no��3����Q��JU�_ke�����>���8��)��dn�X1�j�<{��J��c\�(��p���]rד�gl�G!mZ�	*�����w�ך��}�זQ�L�$%��߻\ۗ�և�}�2�y%���ok�bhvS�]�L!�b=��̶��=ȑı�n�w���Vܫ,���e[��̼��(�F��:}i���,�IH٫����$>
���&��7�Qvg8=��4���~.��^��8;����S1�2�V<��Ӓ�-�)��on�r�A�Tq��Z���y޵YV�#e�!T����i��!���u�^��a���;�XN�mU܃�v�Tә�g@٭6�-06*�]��N�}���=��#;O; �Ѝ�T$�݆�^�,w��k9A��m�����#y�&:؈��>����d�w�U�[���DVv=Y{��γ�*�[^�
:�G��o@ݞ�%�i[Rʻ�d�j_{�;z{�ۦ�=},�a���Tj���4'�;�/o�����޿oY��������}}}x����������w�7�i:�3�1-����X6qҴ�!�bk�8�LE-.��ީ�������/�9�����k���պr �
��VV�e;̞�iϢk����*&��+����Z9��!7��|�,�5�Z��;�/h�Y�����K&�Q�!M\�kxv�*�c�m�1B�R4Q���V�F����)I{����VQ!ɎͧV2��r�D��th�v��yef�
��u���+E�'RɃQ!���La�Boz�d,�Zv�����O� A��G�b����}���;UvʄY�\�/��WiM�kn;P����AA���Jz�)�ZM�F���.P����ǍrW�bWe��l��\��]0��2i�2�H��|��]3Gn_j��wFb��Y'��w����R�TeM��ّ��6k*��j���_�{X�"�c7p�B�-�Z����e*n�z����k�rF�3]d�;�F���"؝;p2r>߻�!eXں:h�����"3�ѓwCk0�[ȫ6�J�CE�+�ۭ'/"b[ٽ))*K.82��Mw ������|6�f��[�.��Phs(��Wݶ���*K�7�W���{�.�Sk�%i�z�6hA\��F����u��K1W�Ǻ�1k�{��-�@�3�{�S��e�{���d���Zt��/ ��a�Iսki�e1����9�=p�W.Fu��D����v�N��Q�H�ҕǶ(��*�5�>V$�q�fl<����B���6�Nd�ΐc�&"�k�����x;)�,��-�wJyA={N�A�����R����X��HWF�u9t �H�PіEM�I�U2��V��e��̅f���U͙��(�J��ޫ��P�m*8 ��1z�x��If8���������(����6�r�*.�E�$�M����Ŭ���J�tޫLͶ�]-���� F��4�M>��[xjq��EX�1'=���@�ib��Z�}V�,ǌ�4j�t^-���^a*��	�;thnU�LN�3OS�����6��m���i�|<,X]s/�V���۞��{)^*Wb�n�
�"�X+�o�o;��4�Q�]���mV3��M͝u���8�]Fm'v�v,�kf��u��G&`5�5�=4q�q֊�zKwV�[юm?��6�ۭFm]:圆,�0^����U�l1\`޻��doT������u.PSzvY�J^M�vg)ٽf� :��e2�C�i��ԅ�Ve�G ��f;����=��W���v��8�S�c�5����a�E��)�vT1���K
Q�0��2��ov�|5���Ha�G�R���t�O7�Jh��#O�k�G�.�Bqmnŷ�N����[����78���Vom�kǍ��ʇp�J���@ҙ]"�W�9��d���@H����#��`�g�;,�<EM����0ՎY-i샅�z��DS��sHoi�5�2Uĥd#49@�'M+�3�M��V^�j0���څ��:E�d��,
�B��%��@A�-#P��q��%�7@P�:f�zx�f|~}<bb|�MM|Ά�(�!�����f���4�CJQ@D�1t��i Uli)���15E!E4�:tD�V܎I3KC\!��MLE1IUITQKDA�(b��E1&��4����e)iJ���Ӫ�Cڊ �۔\�ӌf�AT����m�
(u�tmh�Pъ��lPR�������A5&���6uQl�i��&*��E�V����[P���N�أ�x�7�|g�Q��������=u�s� ���s�5��@m%pv#>K���=�l>��^���-����wNi��k���q����$Q��	W�+���]�:}����+Ƹ�e+���1�����V�3C��*�ީ
���yݯ^�l�I���T��ڤQ�yѤ���5,(n3��=>��랫��왵�Uf�����~�G39;݊�6��H��
�`]�����G��6�Jv�f�����t]@3T���2��ds���S�OA�'0n�D��};�/Moen��)��3��>٘
ⰾN�<[�@�R�|6��6�w�翶6b�����N4g�����7��P��e��kv'Ʈ���������N������JG²']�؄h���Ed�d�W-��7�Ƹ���e��wJ�*��O��]ҝ��h[V��~��=^۵V�Q�n�����y��\ޑ2�P����Bk���J�8�3mO��l7t���Ѫ��{w7�*^"�=�ȃzhE�i!^�X:	�J�v�p�K����YɁpۤx8|���n�h�3��T��V�n(\�C��/������
WIv��Ʃ��v�-���l��+Z�rG����i�S���9��6���(K��wM�����]|39m�JKH�ȝ9[I�����3ʰ�Z�-A�э;����QB����[�=땲ځT2���]�[��L�õ�,st���]w=�B��^�Hׇ"���nغ|ڑ͛�,�2�+�)��s{�wz�v�O$��)��:���p�~
2�V\�u�:B��^�Y���i����x�m�>'�P'�c�ۄ�!h|,Z��Le����]��'�R`������&�+�-�s���*�n�0�kB5�Q���˨z��w%�>�];==��xz�lO��3^JO�_��zT�N��;��l��ߋr1)���/��,�lF)������wy*{�&T�52��i=�6�em��{�$7��FZm��4�ti��i�/�׿��:�s��>3������7�h|`o�o�����Y�g��[�=�϶3�u랽�����Kŀc���wې��e}c
8������?%�l�l~�ɇ.2�\�\����G�v	���Ւ�.���Ŋ�����@V���λˀ�4%u��P��ŏ���N��x�/��:zMF���'�xgr����k��G�	��
$\�ڍ�n��$׶�
"�,��*�����Z��O+r�ɷ���99���w�jr����{�K`:(�����C�T�͑�geu��۴+�x�[O�U��\3,��1"AD@����t[���L	z���ݥ׭��N�qn�����Q-꺯f\_":�|A�
��w����/�7
����;Y[ƕסV�>��H���j�͞|y�Ie�7ec�fT<6������C�|��+Ɛz}s��.�8+�囅*G����:*,=�0Ej͞ݡӣs����.yI۾�M<R�p������$��(Zg�*�t��ݠE��RF����C�j�-N庿{��w�3Vc;�H���UU�螾ˀ�a@��ȑ`n�F�ܑV�$N����ϫ��s�Nn~��7��Q��^#�����v����c�\��q���-/��7-�\ZWNﾖ����=�[9��_�%��vB��3�|�Q��>7H����Z�Aʚ�h��K�	�����?d�UA�B������W�F��UA��~gå�ͱ�4n��N��7�q���rM�l��i��]o-�����ƺa��Y�K� ��Z���%l��)�݆K-F�Q�Ǌv�ͤj��#X���S�+��<�lڦ�7�=r0��]~j��h~Yz��3�U	�d�e*�؃���,MM�v0b�{o�i3^
�d��K�`�f�a������R�g_�q3!f���[����d�t����j��=M��nF��	�W+��f�;�^�r�LurU�ԍ'���'�6Gi�i��g�kK��T�b�� ����������(��Y���\e�k�ɟH�`����qE@�;�7z�N�}U�0�4���9������fY���$O�I[�2�S|�����Y	�\��i�^�-I_��=���0��r���R�6+�vdڷ��|��7�Gw&���/��r	WvyN���∪��|ד�>nF��h�()�*S�)�3^J��;�B��'.�P��1�m4�{��r�N��ڨ��!Vw$�Z2�F��܏TӚ�G�ت9���^���p�x�o��\�۳��ܠ�PMKNm���ٴ��Y)�T:�35ufg*y:��\�oEr�h�Zx�w+�o��ԑ��Y�ݕmǖ1g*שd6j2;��Q�k�˷��kDΕF\���J(4��i	;�-���63��,��%h.�ff��t%3�Rgθ@���\9��#^'��ISmR=�ьZ.�/�,ú��#��b's��zRW��[�[Z�/Z	���z�w�w��g_��������[S�u��
��7g��l�8͝ʫ�Wu�oc��l�5�[�t���݂}��A�dƭ��4�rp�͜d��X̣Xv��gv��tz��H������m�8�����`�{a�\�Ls��>Ž1�ӄ\�41�%���:$�&�a[��!���ڶ�=��d�p��u�H8���B5��86.���^,���O���vsf��.B���zz�N0j�X�ހõL�}F��>,��;D���)7"rP�לf���&&IQ�`�m�5ſ���H#�d@W��N�=@�J"�^�5���5u�Wp�4av�8:�?���Gt��66q-ѧ������(���j�s�w])ã��Z�a4����Brȏ��C9Zһ��H�@b���Q<��;�e�CK��Y�-�v��+��*�q��>�P���,��	�8(l�}9���n�cz�����H����T�y�j�v'�gkM�ś�ˈva�X�LMËK�J��4����~���H�㧛�I��OӐ΃���ty�%FO�S�Q܏��͘� ����n��*ОE����Sߍ��΂�fl<��lՙ�b�͓�fT�_^��W!�8�T�ƌ`��m~�O��q��}Ć�m�xh�1�:7 �/o�5��AM($�+���<ctcQMWzsM�]�T���b6�
�`��ܜr��:5���4�Y��E����սY���o�ݷr�s�k�_�ȩ�H��b�,];]<D������<���f3C�}{���Gj�ISuuK�^��#���bh'�@���_\��/ݬ�,-�%a�q��&A<��	�!�m�@ ���k��W4q��{v���h1�vˁ m�*��\�[g>OlzTz���D�Y"&6����w��~յ�C[G+�Gl��=B������H�]�c����䠻󝵔v�o�H��|	q��e�}����W�ob������V{s5Tb!�
�W�ǹHj�yX�7->�U]��m>��0��6�n�B��x�Gf��I�&Y�nM�cQ�W=�7(���5,ж��в6w/��q#���c��iG.���~vqOW����v�X!��о��x�F)�5���]�w��L'��۹�f���׼��2:�>y�͏p�`Q}�f�tq띫�է%_a/��������T@�5�z�v������~�jͮó�u%KM|w�:_��n�����*�$�Y3�^H��i��s:���e��l)�����|���P���= ��y�=$w �[<tQ��1��T�ثyʯN�R�8��_�3,���H�Q᧛��/�{,��wǙ�}�g��_H��I��d�M�Ve��H�� �T�ط�~{�w��mom���X+��g���
��U=S6z�dT����fj�۠|5�����L���!���'�ߪ%��W�7��(�]!�[�uh��7�n�f��<L�Y�4;����4�4��G��}���}�\��Fr]~1�e�?wC���'@���AM<�w2
��Y<+��I�ʰ��(��y�^6�xv��vެ��r���d���t��
���j,yrgf���&*&��� ky��<\�\r���%�j���
΄�ST���=Y���W6^��l���<}��F�J��R�j�-nS��ftn[Bl��K6(�,�bjp$!�6ۄxV��t7$U���V�:z=.�	楞fU�0��������D��p�C�2��#`m�U�^\�G�q��y���6m��\�v�vWc�g%�;	r�~�B�fz�|�P8�
7!�]UNr��޽�}�d��θ0�(g��#�9�u��ި��t��&}��̢E�grzs4����ٓd�K;�ҭ��������Ü0S���u<�V�oI'��T⵵��H=�k��R�*��l���9��� p-�p'����fƭ���)��85X��Ҋm�@�gs��p��p5�c,>J�UB�ei�����������݋�D�'}F�d�b�n]��SJ��m��콡�i[��3��E�`<*4i_�\������_~]RO�{��n���hw(���X��H_�R���hnC� ��O���P�l�Ι�R5�]j,Q^�E":��wۑ�tjQ��	�+k���� l��yU�gg�{�U�n,�Gb�x��m÷��M�&�Na���*Xٴ���'�;�#匔N�Qγ��n;����4� �Bh"�&T*����ed�!,α��Ń��^\�5�a7礧f�����:�%��N�f�Y��;�s��c��hdHy4��@OE<�wQ"�ro�w=�v[S��b�vvk+r��V��f*F�%�)Em5\��~;,�R�7r�h�E������B���)s�I���u�zMA땷t�����7D\�|�1i��Vr���8G�aظr�>�8f`�ܕ�WX�����۩���=�w�j��5
��	@�b �3�)+a-����&��z����N��q�A��C]9�y��qL��_���UŻ*&8mK�5�U������z��;��K;w��X��HA�pU"5n�����6DTMN��U�����3��u���V*�=����ko����W��}I�sM�s���Ohr�/W��Uaɟw.�x����Z�������c$�l�߆YK����rЪ�\62��� ��l��:���&�}|�������o���@ȧ��'{�;�Wf�ұ�砡���9�B����|��[͙	�ڤ'W�C���u��x`͸�Z�C}�UF�YX�]�ިl�me��S��N1���,90f(ceO�6�y���Dԩ�:d[Ijk�l���f��u>O�j%>������\���+(w7��L2[m{�**9c���"M!�13�hL��`>٘
�V��G�`k������Vw�;{�!�nO�F����������<=��ī� ٘c�NY�磛�$�<�|y$��ò�תx��W�F�U�8���~;���y�2l������Ǌ�"�YJv)�C2ѐr��z�«s�>���w
!��jeJ��Ԑ�+��2���4�6՘MM7OQ�3*����}��GK?�+�`����dׄ\d�D,%)�5�c2wA�j��Q'����\��~��B:�[j�m�
U4]�;9�V����z�u�ɨ%�2v�F�u5l�@)���V�pޡ��z}~�/w����=��w����{���w�����{�������V+��r�[��zN�)��I���!�����ذ�k޾�2I��b���Q�����j	:vS��,7�[���7 �{v��lt1܆�X�'ww:�~:�h
F�&;�,�Kg&�wG��<�������GQ{�S�N����;�ݺh��& ����u���P���[n���`]��g
N�!�[��m�$J@�>N�^�(��";�d��EH�Vmԭ�գL�t\�U�m}jJl�t�����5��j�+;� �>�k{a��|�<�}Wa����=>�׷k���Rܣ'g��j�,a�h�FЊ�XX��y��e���*����{k4����m�XuN�ڗ@�sp����˔�����95c���4��u���0-��tM�RV�na4�^�jjE�5�V+W]יgZ�#+�r�b�+$ـ��nL����Z����J!n,Ҵ�`�un\^ZZ��P�Vd9�HH��Ar��x��d����N(�)�/WYł�V�O4c#�� #6d��6.��og%|ʐ�Ԝ��2�ͽs];�B�dhùD5C��|�F�Ԝ��{�LF㵲�%�m��q����P��F��Iә��qakmβbs��K��Y8�h�U'ImRPZ=+���y��ݴ�o:����$����ͳ�xd��K)f(��ܱ�Y�>��&�G�谕6�\��Ʀ���z6�j�'�A���
	�k� uD����qުa�gLc6���)u����vֲ���'K�=��g�7�w�>wfh���vk;�n�q��4��]�uZ��8D�o�h�yI(�t��Vެ жK�5�,L6t)����0MWK��ݩ+i�,Y/�YJ���۩wd��d�P��r7�����p��.�:�Sв�}����y���Oy�������2���l�*�HIT0�'x��ir�+��n�l�k�%=-��F�c.�J��.[|�r	��)��!��y�P���C���*��F���k1n��ޡ<�T)�⋺�)��,}��Z�ۀ���m�����I/h����̧�=m`�pu�D�P��b�3j�\�j�5��v<R'8
��j�2�(����%�'W./��kTz�I[0�`��Ռ�Clh���z֭��vm���t~ݦC�!ֺ�,��
�Qeɧy�Ww�C[�m�TC�օ�����CtS{���ܖ���E�������76�hsR<[)����j�8P�2���5�k�:�6��ӗʗh��X�Q�r�;�ZF�ˤ6:�B�έ�C=1���%v�M<A�h���ZPݨ�ˇW:ܐk���aȖ+xT������B'�E+�KE��z*��EW�t�	�1s���5��/�!���IkJ���݇��$Ҙj�������̚U��5Ȳo.��\����EΫ�:X��>�ر���0U�#X�k:�̔Q�ڭAD[`ֳj�ns4AU�lh���j���V��Ql�F���Ͷh"5�Sh��s���0Z�ih*��5��j�V-���d֨��VыX)t�/-ͩ�i*�mm��m44��ZM�5����Q���ѭ���K�
�4��9T\�K8��m���ڍ�����4��i�Nѵ#W�95;6jŜ�4cbڴ���U���
h��v4P���r*.I�*�))�V�0QjɌF-�"-����s6���#m�f~�/����P)�]�%���=�Vu �5��z�?�×����yh����v�S%��w���x0�~�7�I)��E������^�?q>AD-�J�IO?\uө��ǝ �cy2���j�6���}%��k�t��7�W�PI��	�,������������	��1����עt�q���6�S@�\�Z��3�VϺ�U�h��v�xb[���d7�����T� ��G`�S#�lOZFi.��h�=�[ݵ#e��`���U�:8<�� 猁�Di��::껕yJ��xgٖ:����G�a�Hw˿d�Z�3��6:��g�^q(�u���S��6F[<_f���oj(Ki�;�2v�lo�|Â�~��s�����)��ݺ'H���ǋd$H; ��;g�1���9�X���e��j���-?�p�'����Î�M����_��a�Ih��"�L��LGa�7T{[�v�<,���6*ѱ�c2�ϻ��Wx��G2���P!	b����]�[(%�3n�2Ȍ��2,y��59�b6���ǽVk�_M�n\�ԣC�{>g#�=�L��W�C2���!ޏw.Yxx��ԣX�=�������7���g;�u=E��}��7y5!�кν�M�W��-�|4w�`2��{�4&j�e��H����'�M;�Q�����X���>�J�u��-�%=�Dmʁ�ɑ���6*���/�Op2(�U�4���b� ��_��p�;],B3�s���j����z�
��K�:����T�fOM>�j�c��G������1}�.e�A| m��Ic	PH�$�>ZܧT�ReBg8D��oE͌�ݴ��)��/XqQ��[��$l7$U�J�$O{}l�e�r�><L����uel�N�q�d+���8����/�oITJ�w�b_������׃�j��|h?OK�
�෡pY��|�*��Թ\f��eKed��뜼�mt����Ot���z�z�i���\ ?-�r�S��W��Ȏ���5�{�$�%��T� oc�,2�O��f������d����y�Uc3^����ՠ�2v��[o��5뾛G��2v�B��=���w>=V���"��J淭��i�Q���/��7�_-���#\z���/�����N�waj�0�CU��J:�����٧��,Ac��Y�DF#F��qHR&�M�;o3O(���_��k���1�)�~���C�Q��跡��V�N�Fߠ�_��Øm].[ڑ�����==ѳ�O���Va��!�E�+���[���Hj�U<e�@Jؼ�N�&I%5/(�|z���Փ�o��
�T�=��E�
�d�#��wM���tL̨�WK8�>�fb� 9J��f�.��p��@B�l0��t�Q[��Q�U!��;���7{���B��ٴK�V�$i��/mO�)�kC����A.:�4�rn���ϻ�������R0�]kS���)u���3��n{����R����O��0f_��j2 �׻�Uh�R��gj��%�&s�F�$��ۖl[�o�K׬��p;&ؑz���� ��h�p�7#���7כ�V��ڼ�/�s��}V��)���v1x[��	,��^B����2�T���0��yݜ2l��-�@}f�9���r�1�I�Xn)����<�3G��+���:6���׌:*�Hg�3��#z�w˄��VIU�u���F�V�̤�=\}$Ut�W��R���ڌ]{.\ó��%��+�cz�|[_�_=��~~�u�=ԛ�����\��p�ՆzI'����k�S����譡<u�1T��,Sq�}ݝj�{Xѝ�r�H�Ļ j� ,���Ŷ��&Ce�mX;��W��O)��[*��kb{��H���#��70��W,�zD�6���0������6�'$���J1�W�	ݓk��� �&�FS����]l�"H9C��>�� Fʝ���ܗRDԩw�&X[6��k�6��͓YZ,���s^>�X�qa�o�2�/�St-�9�g4D��>�Nz�h��z�i�W�~G�_�����3�Ǝg��ٸ��a|dŏ=5�f�{vΜN�n�V�S'����I�fM�`�!^3�a�hmP�v0���]��oƷ0�Ҳe���H�H1���I��~��΃���:�͏tq���7��hW2���R��tC��⨄"Ւ�lS�3�����lδ�]G4*�A�3/�ވ�Yo��C��z-�Θ��άV�u�}w�W;��5�����b�b�fo ��ھ�G�1��Lw/���TH�U)ndT:�N��7���vki�[���ē��:e&cI�K�&_C�UDHي���c<�փ9����Bsu����}��j�W�f �>��ۏiHH�Cx�Iu��mGXzij�|M4s3������c,�łZ�Q/Ox�V�A!Fu��CO~j|���o���0��h��D����t� ܁��ߧ��`���������?�Nc�3�#	�Ѝ����M[��
��v�o�[�67]��D�OW\v`mf�]XE��m�ztؒ�P	%T�q�u#K�7���M�y�̅2���4�;M>F�Z;�$9q4��K�����"�-�dC>�w�ٻ���$$�8�p��S��� �&W"�ag>H��f�-�R��x�{�kgͱ���F��-vzz���S�����%.l<{�wI�S۳���,�I������k#6��q�Db����&.ο�l?�2?K(�K�sq����4��^9[=L+ўb#c�o0(؍����~�Y�͝GN�.�7S9A�����F���uL�iby���v�w�,ҧ�W��Xa��p�m�oږ���\�uouR�mƬ���-ʵ��YieoT�f����P���(&�inXy:]ʹ���P�kg��gT��"�TN������#�k#��/�h{��{{ ^�h6������s����ӽ��;������
��d���-���v��yO����֪�{r���D�t�v�Z�-�v}�tx����)�;�"Kc��l����t���g����'"���2�Z7�;�e���D������͘�k��t�d�;]�D�j�[��@Q�H��jf�5��x3��k����ӱ9�?9�oӸVI�V�}��`��=T�L��\ҍ<lNlM:���{����4t�	� Օ��h�1�oX��3��q�KK�EK^Ks�Y�Sϸ��w����P�]!���M��R\��'��i��K!{ϯ���DW>����oHt��\6�e�6������.I�)��Ͷs�A�2�,���׼��\�$d�
:�Eo^�$G$Rn��=�]Jv������;ΎS^�t�ZN�����r�:Wmm�^�\z�v,�s�e�x�of���Mɬ����N�JRJ*�ᒷ��G��l����Wb����S'#[�ҙ��7�O|3Wa�Z���="��b��s(+�3�pnS�*օ P��5�Qfv�e�������̮������؞�{fWa}rS��݇Z��j��	������_/�zz@a�	���+t9�����!<p�6�w�o:�7�J��%]#A.�:]O��}��7�$>��B��:]��V枙���s�s�pw�+Sܤ��ೠa���(�T�z���s�X�	ژH���4`���_V�=Ԭ*��6Ѷ"��[�oY���6�^��	�A��:�����i?NQ����Cv����\l�çv��.�v�l��v	@��h�&H욧\�T��ƥ�Z;o�wEa������;j����F�M�7��Ic��	��T.楦���͈�	��ɜ��3t��"(��=�p1Y�HIh̉M�j0KSd֝����ًKfq�4`�q�S�<4�i�ԁ�U�H��_n��+�$]I�Yr#Ŷ[�����{{�1�e��ױo`T2��#b>����R�y��������M<|�rBe���VM�眮Y��Y���mޢ����"�eh��y��nv7��P��0�9t��}s\�G�rgd��~iV��M�6E[��쮡3>�Xy-�(*SXWcH�ߎm��?Z��<Q������w^ѻ��è3��>=���rJ�h�\����읢Kd��=yW{F��H���׶Y7.H�ڜa;Kb�E�:A�L�[Lp�Ξ�X��۹��?O��e��� u�6��K��-9�j��_k�z#;���z�;&I%P~���u>�pE@tVО
����TZ�믷%��?w4�֎�%XF�V�*Vv�u�-�� �y�5��al�Og3����"iG:U��1�f�uV�2'�FGkmuq���wE���-�:&���DwV��Vqڠ	F�F�=�*׽�
�Ld�͋�8��ݭ�1�Ƙ�`S�q�[е���r]A"jn���׫�'^�^��O��i'��y�;�9�b3�q�ԫ�O��[h���m�C6M٭zl2g�3wo����e�oe�}�7����͚�6��m�Y$�;%[�8ڪږW56�	k�P�{]�߻��L\p���\注˵90�q�7(ѵ�^�ĭ�+���Ԟ�]R][�Suo1Ď�w���}GJ���F#Ǩ@��s>�g!W�v� *�����U'9�����"���3�;;�{v�n�g���!Y��a���8ǹ���g� �xE?q �������v)��SMRyn�Ne�����*ˢz�o(��{�!�x�x�BG"�+)FN]'���#:Nh�ܳ��Ӯ��9kݓ`��Ƣ�r�i-��x��a�s��_��־�=G鯩�#��;�7�(E�O����ڻcҥ��Z\�[��B��Hw�[��sB�UA���xF�W�=��31WyՃU�f�d����a���Ti:������M[; �"g.i��&y�6A����[%�^X�[J#�ń���j�]T��]XҟIGdC�U6�9W�ۚlU��7)�˷'�=>�ܸכd�ˏ_/z���sf#���|1�|�A�`�4\�m΃TX��L�G;��7eC�dʽȄ����s�3����Лe�TD��Y�p��f<A��8��dc4t�ޤA+Q��Q� ���+6�A3qi�仒�ېP}��p�U��Y����N:�����2�����ȩ�O�J�&� ��vF�&%�7Xw���vkj-�[�ޘ��z��߷ż��y���՝��G��dI��H��x.�����o``�ELFl��DX��M9K/U�od�wr7�f�(5Y�c� ��
&�;&��՚�x���݌���:9uQ�ROt�;h-���n����j���V��jզ����.�u��}��T{��D��&:|ٞ�Ǐ=���`{���Ź�B#�CO����G�F�e� ����`�{����{�d�5�m�^��^��=�i�F��t����̲�;�č��ʟ�6z� �q�������Տ�3��o�����ů=�詼�ܽ���E�E�и�λUM[�W�vn$�t<ܙ��j�@�|sϿ�������
G�� 
��TP_���#�YE���������?'7�BQ�VdY�f�`Y�fE�FB�eY�f�FdY�fQ�B�eY�fQ�V`Y�fE�a�fE�`Y�f &�`Y	VeY�fE�`Y�f�ef`Y�fU�dY�fE�`Y�d$Y�fE�e�fE�e�a��f�dY�f�d�f�I�fE�V`Y�f�dY�fQ��fE�`Y�f�V`Y�fE����|ED�a&�F`Y�fU�`Y�fQ�`Y�fA� �`Y�fQ� �|���f�V`Y�f�F`Y�a�	�fE�F``Y�f�`Y�a�dY�f�aY�f�`Y�a�Y�fQ�dY�f�`Y�fE�&Q�dY�fU�d�f�F�dY�f� �e�fE�FVdY� !�D!��¨�0�UEQQE2#����&UX` d e eUa� !�U�UVUXt� UXeUa� !� !�U�UVUXeUa�U�!ર� ʪ�
���0�C ��"�å����Ȱ�����0ȰȰ�0����x#���*̋0,���#0,ʜe�0���1��>~�����ڂ�(��3 D�����w���~�����������>#�������?����t����Sg����<�_?��G翐� ��������J ���HU U����A� d����K�i�0��և�b���?O���~4I���)�����>�~��?@�v+�2��("4��L�L��$��*�*
B($�� �(��J��@����
B(��� @��
�@��P
 �Q@|��a���x~��E T�J� �A/�}������
�o�����?�� ��������������>��~$~�?�����?ԟ��~b��C���S���~���P_�Q U��?y����_̑A_?0��c(�
�`@g�D���/��'��X ��7~��=|1 �
 
���~g�C���x(�*�����`>�O�����w�?q}��?������ߴ�_O�����Q U�@y�_��C�)2�����������A�����I���_�����~�ޙ���?_��~��9=��`� ��0~OǊ ������������O��PVI��w�$e���v` �������V�ϻ�$��Ti���j
)J�b*� 6�$��ET"(�M�R�jIDm��Z�H�f�Ui�J�*�m��ZE$��1$��[[�[���f�Z�h�a�2խA�3TZ��(�fM����M��!��V�+e��f6��F�$�Y�ִ�Ukcmm���V,b��t3kYY�3YTe�U+)�H�U�l�e��M�1fL��fҚ���f�#-�������-�̆ʳa%��"���hQeM�V��]�T��m��  x��6�JY�p�]��Zv���QEh����JPP��p�*�4�]7R����h�FՆ�իvV�A�(f�5F����
�`�-v�Y��J�H�Y�[J�n�   �>���444444=�>�꾅c"��7�w��lP�B�b��|>���ܤ�Vi֒�h|7*V�1Ls�i:`Շe\:B�n���ƔֵM�9ӫJ�ݸ�j��l�C-��mZ�R��   9�hP��L��iBƺ�6�����n���͍Y�i�e��J�Έ�J�Lf�+J��uӚ�Š��%B�IY���IP�έ&��6U�jVj�ج0���  �eB�V�7*��6M�F�mN��AgYͶ�:{�ڶ��P(Ea�R�b�sp6�nS���J�'ynP��sT֘�*[l�+1�[V��|   ��@�=�Wj�*�����v��Z�e0ꪀ�;����6��jCۇF���:.��q�@%W% ���2Y�)�kF�w�  �r�VL�gUUq;���@gC�(9��Z�V��Ȫ�[ ���n�"�U'wGEk;�( Wd9ekU�3imV�c���Z�o   ,��E��g ���P)�͸:�@������ݷ� �m����4��� 6��� Μd  ���e�d�7[a����m��O� �� �uW����С��q�x @{��=(A���@Q�<��J���m�N�m%��ж� 7Ew��q�hT�ƭ6��ͬ́���  ��@���p �{�Ί hkz��� 8������� ݋�� �Ew����
��� �Z=�켻��z�F)i$̖ͬ�l�Y��  ;��z :o3�ZhG/\  ����QA�yq���1����l9�k�� ;��{@/w��  y����@��"���ʥR4#MhE=�	)*�� hh���L����@ O��%F# 	��@eIQF� 	2���U(  �5O���?��p?��O�
��s�dз�ŷ���\����U���gj{`��G�����_]���`cm�l�cc�� �6���1��C cg`��Ǟ=���u�><~��VB��?t�� H���Fʚc�@��x��`A��vH�:�e:h�K�f��J�6�v���XtVE��$�{��G"�6�x�\��%�*D�`�����j�
fi�N�X�5aлCYvH�ޱ �^m�b��J�{�o��`�AX�&#�ym�m�w[wn����)��;�Kd�I�C�G�	*iY�op��t�q@�5��9��̶��M�R��)���^���6v��@���G��@!��t�G,p��ձ�u0�̺Պ�	�B;j跺7/&�ͭ�������h5�6�̀�\SV���X�/r#8�k�����%���:��$%k�9vVj\9�zպsd@�5i��p[�����z�4.���bt�:t��x5�U�;�F��uc{n��Aw��[�VAJ�
�M�m�H��N�]a����n�
�EȋO-e�t�&k�Z�2v=�O,�vulsU�B��U�%�ό��JR��3Mj��w �*�鬸�B������S{��XxfnsS���x����Na!�[�'hnI+k�pA��)�E�qL@?=��wj7B�(Y̼
;�Wz���h�R���Γ�S[�kׇ4��2��i�Fu�P�m�h��r���;�jQ�0TC,	1HM5�Vm�:Zu,�L٩V�|�+ 9=``��,t�i;�27� ����a��ËY�����<9Ƿ4KU���CZ�n,`҂�Z,�j��	5!<��Y�Y�:EX�v��2d�^�7w����h��]�%'�,f]�cci��0	-CK�&�T -����H�^�Mdb�����D�74Y�Ei��Ϛ�)ɋ�J�Xa9P�R�f �-7����U���3+l��Fm���uq( Koiު�6��*8�M��We+u���NE�M˕z)�72���^�����2�Q��ٽq�,P��R��QAK6~J�;�/��(�gn���eTL�:M�OMk2�㳔��b�a���R�/M`PI�&�	�Q@��{`X3^����
Q=�2�)���a[&����SV�T��ff���4D��v� �R��J�GK��,��u�1��`J7-Ŷ	�"��v�SיmPǪ�[���޽����U�Klw�C4]���\��V�T����d�q�P��п��4���=\���	i��/�'�h��̋^7�h �'v�-���>yWsP�pk�� �$� +h��J
�cTa�!H�&񋥒���ω�H�ĪnWZ��Lݺa�A���mo��J�BZ�鵲���gJ�{�[���DjѶ�w��J�֪�Ae��7Z0�n�ؑI
�L�L�y�r%�(�[����S6w��&�,��h���H.��tU�	i;��(���2��i	`�b�,4�9�hm�Ow0<W�|�lӁK/t�FI��;H��6��-=Vm��S�Ya�F� hV�3'0�<p�����(0��%�tP1Ja����D���ɿb8)m[X�fJ�+tc�w"a���jݶ�XF9F�wt�b��X,T�����7u*�Ol�ZS�y{f� ��u*�Y����A�&nn*��/v[�R�v0I2�PQ�4�>��.��w[gv�i�6l�Z�T�T`�uq�x�٩7D m*J�÷k�w���y[�f�Xhژ.�EN�����qݚ-����0F��J�۔�REBӭ�z��an��f,0ܠ�iGX���X`����Pf"�XVr)��ڂ�ڀ5�c�"��j��an��l��t밚�n�2���� 	�J^ǿf�2�zw/f��c34�;FNN�=��yZ`1"+4�� �X6�^e1���m��Vg�d���Ќ��@4�ӭ���`T��f���2�Z3�jcZ��եW�Ihڔ����-f��wVd,Zɘ��K*��R�*nі)8��"�>�����Z&ŷn��P*Ke%2�y�j�7n���@LD,3W0)�0L� E�d�K4I�%�ݻ��V�0/7h�I���o\��Y�Q�����S�$���;xq�j��b�� �DRj]���yod���%�e�2�G�M*$�F��n�" Ɠ5�n�+F�Uzc�6������!*�ݯ��G� �s{��P� ��(Q�@��l{�R�i��l�`?�[S�l�I<.�br�w�+����!ljW�j!����&�ɫ��<��j	!��w�MR�i�3Y��(]��������uTnDsE�^`��S��U�7%�{�s�a̎��8�&�6����)*)�W����L�ͷSj�n��4�X.X�����^�.U�V��9��2��zm[�Se�H1�r�]b�c�b�bKt�O�_J�UX�c��^b�9Iɵg-h��diX��6~ƥ���j�%���=
$)�=gа��'<	Fv��T:ǟ>����51��Hi��<��s�xD��I˰Z2LM�˴�/��!�zY���5��KnX�<n^�$Cn!Z��U��Cu� 3a�
����T����r7�+P��[�-�
z%(�Q�;�{x���d�6u �'E]e���hͰ��t�rD��\ґѕm� ��V�r+��c��[h׉���]�9q��+
�)'V���E�H�/&ɛ5'�F�r!N�,rlnX;;���jն�5V+e-��e%(�j�u\����^���V����t�QJa�)�+M�efYhej,[��F�}i� "����r�.���6f�%r"�Z�Ғ����ᩔ���N6F�-ˋ ���Cnʶs&u>##��R
��[j�I�F��y������d�I�+�n�9!���L��"NK�vP��ܽ��.��R�L�J8J�	�n�oT�y�E�.G��Y9�%)
c!��77m��jasv�mժe݋��cD��8�kA�9����4��6�m
4��L�H�
����v�)Y�/60�cU��ڻ%��3����q�6a4���B���9��Ƅ�{�-��]
�"9�H���*�[�``��Z����VՌYJ�ŗLP�v�ڲ1�JJ��3	CtWb�X,�n�R��E���j¤4Kh�z*Zk0���1�]�Z���f=�LI�q�7J����M��Z���꒔KF hbg�Qf�^�fA)͠,^n&���l�,�YdPi�z����s^A���-gV��O/x�Ɲ���#ZE�)���J�7+(X�K��Ǉu�YJ����R: �%���V�������%TCj�eJ�0�*,b2s�Vd���$�s�j��Jv)^bBU8f%�U�7��Q�;C2�$�t���j�B�BY[2:*�ꗭ��n1�W�&i,�(���hv�G�j(ܓ$��w�
yw�!+�s9��[Y�:��D�`�)���U�f�C\@^	��x̨�ـ+G��SSR,���ei�2���5+q��on`�L�6aHT��Uz,�P�����KpRE��)eJ�
��qe�M�9le�i���Lَ�F7��t�HT�o"kE�HV� ��Mtj4�T��l�&h���ˢ$�+R�  �S�*nG1�9�6cX�k�$m�q2!~���"���w.�&Hte�N��GX���O���r��K1�΍������ס����g-�t�b �b�j�����%@��j�zU���m�cǖ�|*MAgk^lR8I4��͚*��qMMh�t(�V凶uhJ�hDz���U��A�5htL������Qk9�\9����K�B�&��y#20�K"�-��& bۭ�ٱ4����8�|ʬ�����5,��	O�DUIp��m,cKuq���L���ZѪ��3A�fm�`P*�.�j��#��A���Fjf\r�F�IV�xC�+P=�'疰���=Ê����lj* |`8Պթ��FM����F��P��e\x4�ڰ��$Rl�����,٭{����9I�Vq��5%�n�ܬr�u��4E��f:w�&�K���u`��P���P��BYih�.I%e׷s%���ت�x(/�L'���[<�ܝ��Z����EZ�Ӳ��N�,<�Tk!ǋݺ�@f"j:�5�%�j�H�)�a5�B"�sU\v��]G�m)xYr��F�܄={pRw�f�� ��	]˚�&	�&���G�ScNo1�[z�R!{��`d��
ѭ����blF��U�\�`.�LǘT��ըf�x,�s0� �_��KV�^�A�w]XT��Pͫ�"Ĳ>�c4�35b;A�%���#��{OdԛC���H��O2޸,7�j��;p��7q#f�r�ɛ�"�+
%զ��t�M�R�6���V��u�(� ~jO��g/E�Qh��x��0K�Gi�z�M�X�pa�	q˔�
��TV�+H���e��r[�V��f�j� J����&�w�`��yZA�d/��t�^`�MYsHLԎT�`ID�w�͛�X��DQ� �p�I)��qivn��cK�5Ib�;��I��
� ��X�TV��U/^K��Ʊ�D9��bجn�Ė�b���H�gIu���)b
�w�CX�C4�9)Ն�	�Y
��qU�@f�f��yB�� ��D+Bsact�T�S��]m$����Yqi')G{s7EmА��A��eK۷>ծl�͕�YC ���C��Kk)��X
��2P�h�4���� �K(Pˁ� �n�5e�̒��,mۑ��C�w�1�bfպÕ5H���ۊ��Pj�x~T�@��OZ))���̭R�6�j��r��S�-R2\M34���ٴ��+��Ie}�� s��&�3���Ǩ9��w��T�Ns@��H�p�~����J8Fs���F�ԑ�v�(�w��Ub�r�7.��E\�ݰP���4�Q�")��a m��Zr*�3@`N�(�!���@�{���'�K+* ���o>��)M��pU��҅���E��$�f��(7�x�W[��u�����-�v�νx�`ͳ��f1��&�S.5��xѻmS_M�fɱVÉԨ�دJ9��%��Ar�1���BLG�m����r��٦�;v�z�p�G�oF7>�5V�.Q��2�4e+��M八&+t�����,��|��]4�bQ��*N��-*f����;)�����:CKR�r��l,-#!?8�7N`�e*��)I�U��F\Ȯ��E�V��z[�����.���֊t�b�4̅�i,۬��X�j �L;�n�2[���n�%�a���֖�Zx��=Q�&�hD�bZ�ȑ��,N�ѐ��E�ڬi���e�#yA�!��m�R�ʎ�I������(�D�iJd7[In*	e,ݽqK6c*a�v]�`j�n�	=�����5	����I�k"YD��kd��G(����E�%�Yf�f�z�Z��ݕ�䅭M���V ��T���ocm�j<9����9Xf"��b���Z��nhZ 7i���5�Z��m�73MmE �֦�4U�ˢ����J�n���,�l!dQd��l	����H��U*�X�m�{��A1V�*Ij-&��R�TE��L�ie�<�]�07��:� fYĔTN;!n�y�ᦴ�r�Y�*:r�̓q���MJ�FKLK���Z�)ZoV⠖�'��)�隱&By�jLཏy�1wֺoװa5]��N5L9�RS��[��CMKK�67%�yg �s2�4�Y�C���̷t�ޜF��~����6��h`�=ǔ��%��J�G��Yz�E�+��mӫ�񛗺S���� �إZ86����
n�6U�@��񕈚݇6Y��t��R+q�pи,VJj���9�+^JL��m-�6DƁ�u1�vzs@)�l�Ci�l��}̭=��J��b<ɯ�p�2���`�X�S36��IЕi��ܻ�X@��e�Z����1vYh�C �"��Ӻ5q��zw�IE���wB��Z�L��4�V�:�\��T�!M�[L\��$�U��t&B�A7tl��)�v��n�17ldRU�a�7U� � Z.�&L�j�A�(�T6tiB�Ʃ���Z�4(��V�xF��f��-��k5c�zq�X%���4u� �J�;�I��"}3h�@+��WC_�MW�b�����i�l�Зb<(T��fe��m��i��M���j��.*J�+sP�����,e���[�h�4fB�4WZ�d�Ʃ4dkt+�"45��Rd%gq��1�t��#5փ��YOtݴeP��d"����k���7�Su^��D`G���ǐ��s'fMGA��bf>j^O#MK�3o1,��j ��e7�TlQ��`��`ř�mf�3i�Y&���;ZU�.��)y.^�8��M��Sj�.�A7��
��3V�ې[��"`��.��~,�N�U��P)���@�%m݃��NλU�^c[)�`7���Y� 'V���N��u����؞���"�I�NQ*ц;ff�w�7+��ܳ�H/V$���f퉒�|��^AL`�T��o/Vh.�)��7ar`5Ɩ����MVф��RV��o`̢�o���ŀn�2n��P��DE{�m�-7j�)ܼ8�ӌ���	\�t� �#w�����;�JU�f�Ԏ���񣕱3sad]CW�Y*:;W7[KH���=�j2��w{Xڂ�&��x����˩�Bb��[���R)R��i�����RP�W�>�t[����fr�%w0��-I��K��O|����z_4|��*ַ�X.����l\�n������.�����O�i���
so��r�W��/@}N�1���j<�aC�+3�a�l_�R<ǔbi2�t`^�s�m��4$g�)�B�p���'���|"·���މç�b�����ۗk�,w::�%�C�9��{o'g8pm�y	��E2nj<�]oݱ1�
��gv�@%rP���(1������؅�ЌA��ɮ�,]ɵx�Wmݦ4�û7fmdWGp�|�G���+�N!��'�t����Y�uuҬ���q�mH���4u��<:{�mv�U[j�s�@��)�gG!,vc��	K���VPV��4*T�o|�X����<�J�#ķ����<�?b�^�贍>��C�*5{v�
�ՓJ#5�Ps{v����j��!�W7��M$�3]�U
|�o]Gp��b��r�h��ܘOIAR��#�Ľ�mK�Bj��t��4�`��/�����z�Ć=�j�Q6��Y�.�'@A�Opi����?2�E>Y����񮙒<���a���v�W��\�x���w��F矖,k`��e>O�{��6P=�HE5`��z��7|��{c�u�k������f)��ȇs�k�d�ާ���|P1�#��|��[�/M���r�.'a���A\���M��$�H�5v!p�K��բ�޳c�_g z'���YP�M�����Ci��Gm��uΥ��cr{@]o^��\z/�&�vk�{2Ӹt��oV۽G+Z����t�޻`�}l;�>�s��s�D�]�)VǛ�0sWX9��/M������~�ߙW�>=j�>��2ֺ��ٶ��r�]�x�Bv�=��T����o#�ri��2Z����v1�r�5:u0�2>�ށ���y�O.�������L��4����~�z��ͻi��ua�{6>/Gy�D�¦��?�,��Fm��`�i��l�߭��'7١�l��iX����IW˰u�d���BZ�;6"�p;{��q1���_ Mmh�]�ӣ�C����k(���x��Mϖe��e�rR��I�o�Y�WH��'�A����YpZ�w��L>�Ŵ�-�;�m��DwG�F��4�O\��q�w��N����7{����铕����\_��Ҝ	�o��3 ���c���I(�q|u�17V��;a����(���>Z�]u���lKub����W������ڳ�D�d�M��r���.5w�X�àk�����hgr�=-�Vw�{PM���B"�E�iU���YD5�ލ�G�T��eƦ	�R����ZՍ���7n�ژ�k<���=.�7�b?�,��q�c>28�W��Vxf�
�.�=����S��=��7�rG[#y�{�R�/y��vg��Re7�yr9d�gxܶ�}J{բ�U;����j6=�hmu�ר'B���������u�p3b�<�b��r�O0�Y�k��Թ��{}@��03��(���C�ht��AV��Yg�'Aе��xq2��n��{{��*�+N^n��7J^,����ܕ��{?чp4$]�@$���>Kr��H��-.��"O'�{��V<^q�٦AW�17P�'v!Y�����	�܂nk�������@� 5��^�����r���]��7�=';x%L�=�����9.�-H&�iJ��I��|��t����Q�uK��$���<j�Y��ɱZV(f��t6�m��0��{fj��/^_H�C ��s&�Z��t8�`r�m�7��u�{^츊���B�*�U^d���t"�%����M�y �ۮ9>�t���)��,֌[c��w�0�-��ݨBh���"�$kIY�]l�{���vM��W*!�qרv���w�<k��ge�Xl������z6���k�d�3k�jҴk��_{�볠T����p�X9D�fe�bOeV�!yws�>�z���o��v
��Sڷ�{׍|iWP�Fo'|������O;-=��k�_Cy���Gz��#��u
3�ՙi����#�K��ܱ�@>ܜ4�8q�Y�^��iu�K8��1ܥ��0���_���Bve�{!c�M�.�؜�P��E�����(�5�0����^����l����=l�s;�F�E����n�vx����tSCZerlQ���$n���+�fY���!�:q�r�O�=�0A��a����fy
��9L�$>��t�:)�Ջ�k(e�̮�֛�,f��^b�,i_*}1��,��g�e���m=;F^��urUu��L`rc�\PhÛ�S�HP:T�wT�<r�~^ͅ�j���L�{tJ�Y��\N����v2�Z���}�v���D�Q5��(�\B����ԭ���F��oVJ)6��\t^��}�*̕�"���V��=ͪ.�	�Ɋ`w]�~�}kO��*�7{�v>'����_�L�W�.l���ա���ѵkM����,�Xw��Ks���`&�y���'t?�<L��2�:}f��=s]Gҕ��ɩw��� �]Ǔ�ed�ݝ�*�����3/�;�a�L�Of�RK'�9>�é��n�GK�{S�V�'����nn��i�.�*��F�T3�_��,Ը���ekw��\Z�5����Y&�;�o�ɓ��]�ކ�$�#8NT����ǚ2��V>��e�O$�f�.��JW��6��
u��S�^r�����oV�b��N�0׵�%��Z�S�0L�[,��y��X�oZ� ��p4C���n�yky�l,�:�ۧ1s;g\�4BJs�[��+���!��5-��;����pK�s�=y�XoAsn�2�>���<;lSG��.�K��m�a��p%v��gva�}���9������J�ƮEf,Έ�:c#2��{�����N�wW z��b7��+�Qݡ��5,�������OK�������a��ݎݽ�T��ɭ��{E4�Lx6�-G�X�0wo8�ˍ怪��Ig�;��f��T	�Х�S7�U���Ż{|G
u�����_L�Ew	����M!����R�����JNٹ5F����<+VB
T�^���ߪ�X&��x)�3^��M	������8VA����qL�-E�[6)i.s1]����v�1�/G��&���^�TS�h��%ya��d5�֫e=�]�X-��e�D�����v�Fas�*u@�����9��{�\*�A�����\ws�׽#�d�Gi�'s6�����E���l�=���\}��η�ʲ�m2U�3>{�.����b\S��5Te`͸�E|W�Q�lgϓ�39��/����N��U�lY/7D9	A_Z��m;vI�i@�E�:ᩪs�<W�pL�pIN[6�0�$����l6�h���&�c8���M۴��y�[M�:��&���w0��e��J�	ef�QJ��D�&Wm���� 鏰�5t�q��o�^B9S�v�]�X8�2��Y��[N�yy	I���4b����n��|0�4O[��&f�u�<��5��IO&�"%����ҧY������@q�3K����5��w������Jl~=��f�Ի�t��(�5�m�{΁
�B�cs���f��僙s��i������}���2��C�h��ޅ���4^�nh��˲�O����g��ýJ����UG�k��n3VAҳ�n��)w�=�AC����J7���#l0vqӤ�=�KC�sDS��.�Ɏe�)qа'V�����O>����>x�2�U�yY�d��)Z	��{���Օ|�^��'�8B�s��=�n�j�V��$G�k��͔Q޸kg���NUi���c�@:��3e��G>K�|F�����w���ܼ����Բt,�
�n�9�f�N��2Z̵T#P�	����*A�<rgPa����s��s�S4�)퍆�'
�Y��A�W\"7Fق=�L�K�����m�Mҕ���p��l+-�ӭ��*�rϸxz�,@��c������ڣ�6�F��moU��JR�;z�`���`��8���Ӻ��=�j��U��_	���p��\\��P��Wcc��o���!];�f���H��9,�l����o��g 
�21-�ޞ�U�ʦ��/W��O��!��')�H�W:�K��Ss�qFƝ}�>�t���^~ou�>޼�Js��ү�I&I�;s������B���T�6����=�'�B4a:�?N.����
�:� m�5=��5̽���i�8k.�5]�13� mE��:�դ;���A8�S3R��`�r=|��ԭݨ���2�}L� �fe�-��·�7�q��j5}l�̫N�e��\h�^a��t2��.��<���TTɡz򵪍'��~���8o>��ּ���[{y��݇�Tvj��y��pE�sW��V����읲�`G-�)��iݛ�"k�{B�m�-��{%,���B���)�x!���
��n�� �x����ۡ�a�FC��8<	J�O���9��/�]^�2���3�(D-M�4�y�F���*�w��j��l�{� #)\˕u6�v� �(�ou��x��� Ŷ���]��FC�]���w�1$M�[]x]���hA�6iO�g!�к�.�Ǽ��pٱ��[��q�	���]k�w-�g�Hi&9��.��%J\��D�+������-�Yh���6aO��m�x���#��LN�{f�����FJ$B����ja㢎[�ƭ>#��݌BE��|fY\	��d( T�����eh������7���Ƴ7��$z�<$�8��c�AT�'����V��cHg\�ƺ��v�>}��j���pw�I
������ۧx����J�F\��
8�1�>��p�w�æ�A��,{�=�ge����T;�,D�k �>|s�mp���e��4#�m؛�v`@�������'g�,{|qQ�I����37�u���]����U�78V�v	�(%\��y���-v֢�ɤ��t(�,\'�V\K,�:#{-�\>�����`L�L���K���35�l�.�x#��n5ӽ�с�y��\�V�I�
l5��t���c>�<"ٺ��	��yў�8ڭN�؁��h+pgᔷ��RwR��a��򯷯�>gur�;HkV�]h`���l3��2��H� Ń�a��t{��Q�)E��ӂ�(w�n=-�C3S�ص���䷼����R5�Qy�vv�le�6*]�3-|PM>uv���)E�>˜��_!��+����b��I�]��WV���V�&�>�v�^
l�ǳ=�����rJ�+eA�mJK%����:�pn����.�n̊�g�wժҡQ-�1P7�r�������).ǥ�f$�#τO�|���o�BDPwtH�F�T��P"�=��m�J��0�vT�̿���k+B��YCR�����7`��
zS����YH����	���2�+�
�v�X
]i���X�ς+�ʧ�j-yMrS`y�6�^���,�$�v���錫�r�;{���tF�a��K����q�B�j�L����Ԭ����\1���y3��6�����1��F��;���*����K���*wq��VWpk*�E{��vӼk�C�@��bھy]���[ZPX�a+�a�ۤ�hڜ�Tg�sف��[/��+i4`Ng��d��7�-�Y98��kM^N���|j�4����G)����f(�c�h�Bf�
	nb[�̵�xΚY�uo�o @>���b�w�͹�L��J�`X-�+y#��]�;^�;N񦽙z0�u�ޛ�����m�<�
��3s-�c{`B%�)��Q� ��^��#�9�=[��5�rxj�i����Q��p���p+>^ŷX����xܵ�:��<<,�&j�Bu����N�w[��}�Cw�iZ��U�b�F]j�#�#}�8�;Իge��q��qm�'D� ���9M{X=�̸�i��"� B�E�)��f�#�e;��k�d(]*������- 	��HCb|��8�X�8�<��Uc�K����]G�򦳥u��g;������Z@�/��g e��\gq��̺�s��)e�./kP�V�Nj�B=Q��"ua4�yƃ�h]xR �����d�[[�~�q��m��]@�f��V�u��]��tX���+�����Ͱ�+&�?^C9ѣ9E��CI��lŘ��%/���Ǫ��g8�N�㷌�<4��Wyn��"W�6�~����6�2�obv^ݛC�$�B������E���
X&/d�3m����W���[f�Z��S4���Y:9�O���l�����W%m��HB�p�������o{��-�x_JG�2�w[�&�u�n�5�N�;l�n!sn�3Ě�Eo�etu/x�_.��zg.:H�|Ǥȉ���#EWzՋFT8���QaY��`��tO�C��8:����@�}�D�3KQ��m"�KOW,�ݬw`��%�{�-��_���ɨp�[��j�Y(D���n^?�A\ �kT�A[�{%d��pZԧ5|�\��H'7�(��?I�I)=�q����ǻ��>���ߎ�_�_r��[��/��Q�\Q⅍Ŕ:�2\���*nQ�����"��s=�Sr��%��r>�Ժ�6��Z����ǝݖw��W�R��+x��������%��o�g{{U��{��d�^β�P��n[�Sh����J0+�v�e-uYD|�G��*%�ޙm�˒�]��mv�m��M6�'��|���F�Jq*Կ� =�{��π xx{���9��L�Ri�|�s^Q�;�։�dfZ{��2��N���emv(�
ae=�H����=�M��D�0� [|9=9n���1.�S7v[�]/=ɫSed`(�!��I�\�̤`6"!.�>�la�Ktõ��Ek�pr�e��V�R<�m����v�����n��b���� ��ݑ:ވ��Jx�a���jز�LF>f�Մ�ݙ��0n�W*(ئ���hU��O��R�	ң�.�LYO��k�Pd�z.94Z�W��fo��]ٻ���l��%{�#%�Ϟ�9gnEE��3,r\��s��� wszSX�ɔ-n>�)�|dc1j)�[��eM4��!N�7��a��Z��	4��\��x��/���/e\U�+��]�F=F�-m����	궮 :� ICS�x�:��]G����uk�ێ���?��;�ӛ�ٗw��u� ��-Q��1�6��ےh�s��r�u�f�hC�{��!�wqY�l�:�=F׀���R�^735	�g)ޭ���ֳD���;<Z���yC�e�<8U��Y-%�����`��(��]5�ݾ�7�D�����)����3pbfX�'S9��vlԎ����9��ͧh
N��&���2�h��8zC��P�@ou�n����s'���OP�e�<-��wmLq�Z��F�'��#�n ���w{w������W{��x�~
�"H`��zBR3Y����%+��O�:̗3rt�8[�;�����m �cy6�u��z%�;W7;�⻿��#3V��ak�:��Pb���6i�|�:�V�fm叙��;1.*���<���nE�*���5;D���Z��8%wK���!q<�a�2e��u���-V�GB���/����l���-�5���K�We^��w�glw��� ��B��P���SΡ�A��*�q˞g1Z�#nXP��\ޡ�v&j�{8n�1\� �]ǑԲ�ޯ	(u��w6\�޷�/}�73\���T�]�a�V.�s��t�5�'nd^��dyB#o�2�3�_�s2��#�؈Co�w�p8��(�qۧ+vo1�Eue6ML�uψ� �1,�|�`�)�T���d���ҥ��i��f��
/�ӖBY� E�y�7}YE��S�-���᯹��Xa�׾нJpG�����i�c�����B�rvb�{ύ;V~���w֐�T�WF'����V�s��������&u�i3�n�_�j�?"��P���Ζ��M7���{kl��yRwI�6G���9D�P�fVa�zT\�\��6O5�&#�7nc�^XL9�\-��L̩WG��oS��]7���C5��5b��5�%=K/�d*�:�*U�,Wmh,Cy�Rd�Glf� ��-z�h�����WtQq,`�0�[UܪƪH�齵X�'em[��mY�|��Ԏ)m8���sA��w��#�c3'˸���FN��˫�x0aƒ�y�z�n{�Ύ�$>I�S0I�t�i����[n�w^�cEl��xO��V,\����q��- ��.��!,�a�l�ޭVB	���eA-!��O+�b�u��pľt�.�ʋ1�bKp{݈Y������Y흃6����^a��:n���ٗ�����E�Ӿ2f��hq��h-Ή;���I�N��ڄ�[�0���|��b��-rs�;f�<\ն��kI���3�M�,��S!�����d㢄�"�'��!r��t��(��wJN�\���w%�M��?�#��c Q��O��8LnjKe�y�W�H�)��c�oE�m��I���FS���d��Rsj�C������e,��/�������j8��<cwY�Z$�tw �d-T�����R��ʉM� �m���tZ;�6���y�g�K$��*enۺ�r��R \�
V����J\ͧ��Im�x`�
������!l�g�e@̼/�W6���K a��¸u�5���"/+GUq��Z��F"U>]��,�v�N�ރ�\'5�e���κ��뻀��d/t���ëH��Έ�f���f�[I�������.tjn�2�����d�v	�ٵ@�Z��T��ew6U���y���mM�7))�i�z�|2g�1eΧ���,: ��G�����󵆶�35Ö4�����p`�(L�@���
 oq'��K��������.��=e�)�o7��M.|n��#Kg3���&h�~#\Zf7�Ho�I�iZl�nL:�zZt�ZZMk9n����}H魷��y����Y#4a?q8Äm�%�{�΄�(�w���|0d�NQpv�(^H4��F	��۪�� ieg�K�0o����Ō�b�����o�������x���K�r��c϶�Z����0+�jA�hOjn�Y\�\�.}o����(�c�)qyĘ��LK]�T�B�=�<���R��gm��<GRw�l�vqHm�M'��i]m;� E�k��Ր���i8�8ep,��qLJ��g"��;����+N��hM���+�G��h���{p���]o��?!�a���eZ�cɺ� Y�p5��|D����9ϭ�����RO�:?��D૷z�5u*�4WFF{[b�,݋�P*ِ����;��Y苞(�3%�<�!����!�ۍ�6ɗ���b���uΩλ��+��mC�Ri���w�Fl�v�96յUg�ʎ�5NF-��W�D�,e��Vk�,'�"��[���P}�����ꇎ�M^�N��O͍��]ǚw5m�x~��]+P�ͱ9W��`�ﰮ�Q�x�s w1t-^t~�A��3Hg���a)N�c*��5ղ�x'!1��(�$}d���((�e�;�)M�)��-����"���u(t4V�x{:Q���q�U��7����B�pj5���Q���	�C�ϗ�clr�?��/ {���j����������c�]��9jQkU���#�O����W������,�onAW�DN��T(ګ��};�:�u�mō����W!��	�`�]�b<UCl��	���`�vu��c<)-�
�ӹTt{'M���D���Y�,��}��ebS)[�sI4d�c89��%���dS�Y��6�ɜ���m!�W�P�4�+tN�p�;�k�Rơڟ5����'�j������5�E��o�>�&q�	�Փ�;.�J�υ	ʠ5�|1�EDuz�X4�,�;ۭE*ۧ������	��p�uo�;k��o��]�(vY&16��xם탶׷� ����ҟU�臃���n��Xr�̵�t�x�36�b�c�����Ƨb�����;�!�v���$j3Є�a�
�N�_"�6�a�
�E��1�}W���N���r�f�6"�����tb�f��)Z=�^�
��8�A��`�1����ƌ���_h*�M���h�h��e���=蹞�g����%�ښ{fT=�ǟe��n�u�-�#���.�9��yH��u۝Ո="��ܻت��N�h���1n�}�� ��V��l�.�=�c�,��z-�nӭ8n��Ճfec��ulV,����4�Q.w���78a�?4b�W����i�+��U;{��-���s0��җQ��v#g2k^8զ�e��]����X6.�L��b�,�`h���%$N���rJKN�a\�ɴy��m�7��m+i�־�s�tvtM5���Օ���n��ۆ�jɶy윯8ξ���O6A�jtm�3e�P�ӣg��w��A���߷6p4���!7f�;P_/T=x6�\5f,˚[��6;�x�VB�j^"c�55u��t��G/f��l��-�G��pTNpw_<[rk��xq*$�t王�����z�������2`}���cqM����j����qRB�G�	ZژmZ��F,�,�T̔����,�����.g����Z�}��N�㣍�U�!�/Dt#�Aʛ#9z�����q7��ֺ�9�&��pc&n���p���6��P{A�{�F9��m�1x??SE���F�Ո�p:�����RbB�@�-U8ϯ���ק s;Ɓ�A�vMȻ(���yj�0��
������W!S@܎�z6{"6;����YK����J���>���|�K��̔�t�u�j'��z��ˮf�p�[*�8�k�ɣkNR=˘����8��a�> �(������4�o��i��<�p���qeY�3kaP:v�72��]rK��Nw9R�Ή���G�v`��W��GB��]�|�D�un%O(J��1;qi�4����^��R�@��i&������S&6���7ӏ����M��:={e�A���3�&\���������Cf�o��y`�Q=�XE�b�c�(MQ�KN'(�q��Y��5�G)�4�iЫ��5&k������:3t>w�V���Cܷ1���L]����9K[,�$�]��g���a�j�d[�w�ࡳG+oX�+)��q\ �9����\�+��Aa�=������C������}���e�3[� ��Κ.��'ІՇH��=�#�Np���:e��ە����tNW4e\���w.L�K�kS0�J�pu ��շ��'nȞ�E��rw&h�m�91S��۾)�pd�z��Nl���Rmmr�	����g��s��n��iw^u��$��U2{羬b���o�z�mT�p٠�|�W�Iƒ���j���$��I� S ���H�=�\8d�/xͤ- �IL�O��NtxƙO(ֹ//v�mm��gW��l��F�:�y��=��&�l��7x�sy��R� �n�f�s�����A�>:��
���&w�/l����U�k�>'/�s����9b^�f�f2��mEl=�/E���0gL�7]�����SK3]� �|�|qJ�n���7	��j�4Ǐ�V7K���Wx��=tv�v�{�=}��x)v�p�^����~��q�PշL���x�*�^]Hɐ��ٽ=<@��}l�b�Ɗ��i���Q�߸�^�A��wP�C���l�yL`��ڶ5hy��0���l��s�����@��N<�Dv��=Os��+m�Sn���<�i�8�̂j�:˻�D�S(Ҡ�m
H��Z��v+V3y���;��7H����6&��#Z���F�ۜ�f\׵��xE�FNo:�pjWM�F7m�k�1v�7t(�FP8�y3mݥC�jՎ+�j���S�C��f� ��ux/jB��8 h�xu\6�����VcJ�m�iVϏ7�S��a�wx�K+�@�E�u!��<����B�[�G��\���Ʉ���о����8�jb���/C��Yp�ā���nd�Q2�و}*J3�[���]���*k&���E��=��R;����9�M���T�}VP��\�L����8��6�[�͘:6wU(���vl��Hr�r�3J9ɩ�`A�;��F$z�vA#��ə}z� ӫVwΑ�Nz��.�$�+;6��b���S[1�k�n=7�)xD�/�+i����8����7���N<$(��:y���Ža�
ɭ����%�+�D�Hv��$=)��K�Μ��%�
��^0�Y�;��嫐��$�t����LtT����yE6���w�a��7�i+��>���@����˼���.gt�<��u��;�h�z�0ob��0V�ɘ�%
ƥ��_j�)�(\�F�P���}�kBcnD厅�ʪWa6e�����������W������|ޢ���}�)��t��pK:��=i�MR�oL롬������"]g�2_pa\�L�{�J���P���}�'%+6�h��dn�^p�,�*��-��);.޻�&kUT��A��GnZP)�RZ'��
��б5xI�^,��{�)ǩt<3P��9��=>ܪ��owf���>x���Jbp�i�O]It��w7�ab�kX�.�w�}�o�}��7���ޖ�S7�w9N�A;��;G��}w�S�J�q��l��8���K����m�f��o�h�B�������N�Y�mNW��5��%afml��/���q��)�H;��Zrc��"��N��n4&cc0o�1�Y��f��M����AwΩ7-u��y���wy�p[��/s9gfS�nm���{T�s1��!�|�
e�8���E�<Y0\P��{���A�s�	<�<���}�DkkK������ͺ���A���`ض�y�!�,Q���98�q��&g��;��ux��u�OIM�Z�ORzI&�\ݫMZL���?Iʪ���zn{��o�p�K��6op.�z�LJNr��>�N��*��ۦ�'_�Օ+E� ����B�X/�o]h�J�1�+M��(WqO\Dw����/0�M���Lh�r�<;����K�����
Cb�ݜ��̝/�����[�8�@N:�(��1��Fq˃+�Oj����w槽��KEzQ4����֛�pN;iNK�l���gv��!��v��o&�����޼�9�xWB [�p���:y-C \�:�;UJ1øO6q�t;���2�������{w��A���n����*y{%�\	�:[�v�e�|.=�0&�ﰱ���^�J2�9E�5��c-t�%������l�ɳ��߸u�j���
y�n�.|T3+{��(/�Ə|��Mև�%H-�Ŵ�,�l�B����\�&��>�}�3C{3�S5?t3&��PA�x6'�oƞ'�������������p�k3˷g�t@�û�x��������`{��������A�ⷦ�#�	H@Y�׹��q�'����{2�/ŝ����B�*�-r�r�x4��D���[Y9������헶�_,,�Yg������z�?�sW�;oH�Ў�i�v�|*�6�g���qѨ,9�8�|��(�rS�)�U�z *���͏��Y��v�q�:�u���]E
�,�Ŋ-�C�W���Z��Z�N����s��z]
�]����{�TA����ު�빨V�?n��MĻ8L׷�-�&�m�۬�m�EH5ݗ��4���X��j�y�D�zn�r�X���)�ë�Ә���[L�[f+�2�H���pX�Lۭ��֮���=u�t���5LӥHQ4�.�!Y$:2����t*;�ԛmڣ�'�F҈���@C�+��=�3�*O2%�Ŝ�s��.���ɘ�OW{n��Xɇ�����K�etջ��Yo��K�/����	��+J��C���r.<WG+���
��db9��	
ݯPKK�N��Z��v�Z��T��ժX��5�n�wWQa�6�a���J�����K%��]g�����|I.0w:}��4�Xd��,l{�v�Lx�f��aFSu��:�
թn�{��:�7�&H�����݋=ƫO)���nN#�b������ڠm?�؎	#����'D��po
�d�}�;�w��\���#���&��H�BI(�EML�:d���8���RE��b�j����Q��DVADR-�YGVm"�e%fT	h]�(ENYFf�h'Hq9�KCCe��);�:����9N@�7 ����k")"�V�A55#M:�幹e��DT�PU45(H5J�
����,j̹*E�ǖZ&�%Kǈ�ЊE
�ÇQ����P��%B�H�V��)��/8\FPI�h��Ud�W
�2MB4�ki��'\�r���\�"�$čVU*� ��Q$���-XJ$V������k���bFfVTRy�
9�Ǉ&E��
ªL9jH�(��4
 (B���8 9�PUx��Bc�`wh��t��Zg��KW	�-���{����ԧ��iI:��"��b���S��~����Βf���8J�FYg�#��ͳ\-:�+E=޹S{Y�����wg˟f�w��8=�Ҙt6����r�ۄB����9�{�]�6��d4d~('r��u���=��D:7E��On������k�j?�i:}fl=sm�F7:5�1�����
���LNF��bz�c4�"���D��������l��j/!�@���r�Z�|����m8��`q��JÁ�����v>3������Wi+��P;Q�"L���ԫ��w�
�e��X�3���q��v��3�䇼��ֈr�.+����u�hOt�b�'U�Ϯ'�������Q	���crb�[<���t�*�p���b���1�{�^3U���"�N��>�!�!1�ʂ���ui��=כ�y�yE��kj�d\�N6���K�〓��.|=��SK�8�u�(��껓����.�^%Qё/ֶ�Ie��>q��(�3��n
.��<���q<=����Dy4Ԋ��\@Sw��WWR�m���k���C�T�Q�V�)�c���i��^���{ޣ�zC��]"7�6n�*�S����SkFNѡ���m��Z�ձ���}܈�!{�vK��{���4�ϯ����zduz�v��>c���睺�ӗ�]�ts���3�.B���(��b7�ne��3N�[U�l�Z���pF2b�+\�xq��Z룣<����;��q7��:n%�<�*7Y.�$ �{����7x]>�E�d����6X������FE$ը���$_��C%���NjNf�|��n���=w���ƶ��quG	v?3>eqھ����6�ʃ$[�p�D�uQ���'87��Rλ�~�w�v�X����w����Q�v,o�37Wi��ַc(=���-��77�r�aaL�<n��]W�b檲J�U�P�¬xA�v����A�8ܚ�w��;z��}�2������|ɧ��N�YG@����Wr����@*w��zR|�umL�g!S�$nl�w�n%/lr�Q�'����*͞Kq�^g</���S�o��ID�A���#]Hzkĸ�9c��3ʼ4r�g��8��LfB2��>��i���;9~~wSjY;�d,4J�^���^e2{"B����`��6�JI�!\��0��Y�E���}>��@
ǗЕ��*@��f�:<��j^z�u9�s��
�/�GQV�K�l�ܙ�f<�����+��^)���Hzx�	�˹؁�i���,��W}�l��K��l,�ܾ�g'�W�*�6�S��N����?:����ދ��<N	�Iu�V:���lU^�~=W��ӣʱ����c�wz��t�q��>�����°_�~�aE�:$�I�N�?�X9�_y�5�-L���I�Q�$fd��k���C/�)��~��%r�����a ��\vDF�ʺkn��e�h]��s;Y Wu,�\���n�zư�F`.!��6�>�)�g�A݁ưGH�ڶ���N�����I^���HU�3dt�:u�c����i�5����t2��d�

װ��Sk�WN��D��I�	�Vb5�S�Ca�9O��}��yF߷��:wn�{�+O��z�|��舄Fzx��`ߠ�/���z+�"J����2rCr{������pT<� ��"89�T�*+�R6	3�.Jӑ��9aث̜�"�D<��]̚�#vƗ[�a9�3L���DW��&7��љSƮj�,�)>��,j��ݭ�10�zE�����F>3$hI;2m�Z�0��I�(��m��Zw�����b�c�M�|"t�7�^\[BݺP�n�^κ�W	fԥBzL��ro�\�<��@Y96���)k3ռqwe��>{�3}�5�<ķCS�ˡF��b���-p(�� ��ۊ��,s��v�6�z���h��ɼ����΅�^Y�V%����d(���(�N�b�3f�r�$�7�O*�]�U�TRy���S0Z�߭eHj��� j�EN[��eŀ�S�`-u�nvd��{��;*��g���0��S�F�?��7B�.�.�щ# \g�e3�]N���y��uu>���'�T����;a���`<TDV��٧CЪ��X�N�������\_\���&��IT �[��(�2�~��g�5~�Vq�@�#"�98rU%���������e���U��/_Z�n5���ˈV#h8	e�A�&V
���c�ޢ/�n��,T���:%Gu�<����Yqb�v�P�f;�z#����3��u��	��"�L�l<��ܹ��MvkB:拲 �G��TV�	M-�>�
�UӤ��F�{�Hq��!�=C�Vi�ɷC�ƕ]zl�����.K4�U�0��B��{=�v%��R��yJ��ٷ�u��1N'S뛷��:����;M��S�W�Ow j#��C�xS�Wq�[n���zn��5x�cH��Q����^<��U{.����l��}��H>*��d���-����d�5�Ewp�<$�X�>VM"�%|�×��=�q����1����uAl���@:?oW�u��jv�M���9x޳�ݛ�]���|V��ֻ<����NѰp�0�Q�Zs5㩋�uhͅ3�=�f!�>�͈J�˒��l�y�m��hFa�:;�=���T�轖����z�faQRLf\q�xeH^�؛����G/Ʌ��&V�â��j]N'-Yf [%s5�*�	�|r��nY�δ;;�ow�Q��^J�E'aɫ�\D�u(v+0���>�9*d�ˈǊ��jl��5ZAWR�d��<�花�r�dtU������1Of�P;�	�ԝ���3�w{���^��3;����ؼ����?�Ľ��э���;�l=�pR����^l	���!W���L�Ӊc����=�E���On�����!��.;d�W���\�HW&v2_q�׉!�OKf�_���Ɋ�V�����v3MDMA\=����F��[�����M��t�1S�}Q,�r�i�P�k���Vu8�g�����Wȋ�S���:�����ʻٗ׾
�9ꢫ��^�����E�¬p��Aw��k��}��6<���%;���c�׼�$��9M�o��gW9S7SoPa��
�J��E3�e�7��wq�ne�9����m�R��S`My��ꐚd��I�TJS��W��ޡ�����,w���=��ŭ�F�A�!�u��:��|���58������C�{�_@��\��-.�s��!�[�crb����}�9������+{��Ȭ���o�O�ݱ���'|�����@|vQ���y�2�뭘�\��U�cO�^;	�r�8�V�B�6H�8	8�����K�xo��Y ���UI�� �Ș�����,�,i�<�
6��7�����Lͬ˫�3t����7���L�v��^r�"���<�a�����-����Ғt�ov����/����˻�J]9�TZ룣5~�3�\j�6^����٭7�{ǫ9�ٞ·�}P�«H��aa4���P��5�t�DdW�j�`r�3o�Qq��(v�-��D�}��c�4AduxA�F�9�M���^�N��'��K^��2P|ф0��}N
�C����3�������#��;Qc|q�;�í�u������^���ԃ�S&��7Q�L��IM��P�]}�2מ��4)eZ]��vܭR�]��,dK�q�L��;;�.VG��[��Rmʼ�y�ӭ�z ��t�W`��%�Z�^���P�.`۷���@%�oi#��x�:qs֘���A7�^8's��1��6�dI��\^�Y^��u-'�Tf8�������\Vx�=+��-���3\������j1����Oo����v�Q�v?N��Ď�@��"�[�$f��nXJ�`���q��m=������M�fhb6��Rū��,�/�Q;�g�Fa<�{�xX7+rp��:�����+y�
b���Oh�	�4�r�+��9���R%�&�'2|Uu�G��(����]�v�
����E��vp>�W�̒�Ñ,M����met^t�B�'�	V`��S�FǺ��{����E���hl�}��š���ɠ��/�לr���Λ��`^�$H'��vR㍬v���g	�����U깬#N�<��F�pl9��a9L���l)Ƒ�C�0,=��h�*�x{��O���@خ+|%d�i�iozx}+=N�fx��v�V`SZϤ�[A�[͹ۖ�}7��!�tV���$3���ZΊ�
��E���D`�0�6C���~�MZ��%�ثl���(�xoI��BS��s*�5����4�^����r^�{ϱ�f�},�Ӗ��r��ڞ���~�U�ֹd6��on�7��g]%�c4[�M�ks���ca�����ins/�C�24��^¯�����}W>�ZK�����e~d�xkV�ߠ�zs4�{޻��qNw>as�&I�l/}�޸�*"��u�N��8ҡ����
��=��L�m�|���U^��to��U4s�g`6p��m�{��(�TwT�l�=��,T��nh�KR�Tk�f�zԺ����
!D��j�|�EG��o���n��������Õ!��Å�hs�x�5$RIٓ~n@�a+�/��l;�˔�Uu�M�������.ȡ=�2/�)��Y�myuߔruS�LÙL��2�MyX��w�juo"wc�[ʘ4O�
����� ~�:��8}n�!�z�w7�D�d�O���B�y{{�y��N1��ʘ6]f�cHT�:M�`�2�c��+)�~5# dX���no"�쬙z���{m��Tņ�����E��#�_��O��|+�,;�g�,��%w	���;Xx%Ms,�1l�y�~�V�@�#"�98p��`��# �Q�k�أ]��U�`L�uC��v\B�A����p]Jg�O@o��£�*h^��Ğ\ӣ�a��Oc�~��|I��[�i`'��Հ���<��9;2��b�;�^\����\�|d�[��{F��}�~��`($�7�*F��Y���s��xr���Sh,���+p�{[���[�	������}j��nvo
�F�W�`�>�>c�X��ъ�]��@��3�N���.�mT�W̵�o���!��T�Ydr2�(�S=��E�V�]�X#[����!�����|߯�F�&_x�v�^?set,rQ�#ĕ@ρ�>!P�)ʈ��{�>����a���.�]����5L"6��C�`=���w~w�H�F��Q
C�BG��o�3�,�K����v��S2�q�T��31۩��S�T���ï����}e�����;y�ܙ�|�S>�ˁp��[�Ѽ��d`se����t',:�f(2Q��dd�5nd�vw
�Wϵ��l��'Z���8���V�{k�.�
09j�9�F2S��Ȝ��WFlL�3�g_.�k�KFrJ�#�=dd��&�ܮ"lwR�~|�Ëg���%L�z'������?+���x	��E@k�)Ui�q��a�����y��*��/%(����v/j��;�Bu�5×W�_
.#���G�œ�=�b�F�:�;Eq|W:4�qը��,J������3�M|%eu��Tg�w�9���E�:�����׬���ع겫ӛ�Q�����t��K�;zX��񌢬u�/u�P��UřB��X���v��.^m��+�[�c�lE�Z#�I �i�K֥���yԔō�/f�+�w�:�tlFQp6���Ŏ/&r�!��.;d�^u��f�
TmM�J^�C&c���r'�oJf��j�eHxE�b���P�Bv3J�PhޔH��G1d��r�~z���y�-�X>�œ���J"��X`�JÁ����m��3����ĸssC��'���=ƀ�eW+�x7� <3�c�_V�Ib�I��5۳���-P��;���=�����~��kL���� `���iu��!,����ܘGv���ʶ�Vjƪ&�Jv��W.�v*���S~��N���ѕ^�$�ƽ�!��s���#^:��Wu�1��؅�����,c���j�n*��Y��$�	�>�M����G��RգG��#��Ѕ;�K�tיqQ4�[�Ie����5�PQ���/��GA��������x�S6�$6����P^�P�T��n�4��ȿZ�#��1�����P��#cE�U����}��8����b�zLW�<�s����GF:j�a���S�`]}_z���i&j#�CKΝ�k��6������,�p��(���ƶ�h}� iѫ!k�X�[��Wb8���n�Ԏ妋qm�0��v�y��9VY�Eж��З�ɝB�o�9�L�[���J.����ꎖ��
�} )���\ߑ+�z�[�{\��oF�n[ͽB5�еyܐ��8�`J�#�� N�=�� nV��(i���^�}`d-E2�Z~�zO:������G(ڱ�A����X<�V�^iv�m�YƘ�xUKv(e'��|��;7�s�1z�Ԥq#���9Սb_S�s��fŖ��[Z��A�;��4R�{��t֯R����ΫA���Y�7M���iX�d�7:�N�V��Q�}�1?Sg����j���('�~�6#��X���d��ͯ��aGW���}�h�v8pOvԴ��I����1���B�i�P:�\����*�H
j�J}7S<�n�vWu�����������V �^�u�7ol/��v���ּ�n�U����m8đ�D$����Ԏ�f��k7�;�n��y�GE1XH+��V��m�r��5���3-Po�U�8���
A��.�#���e�X�����s�M^6���Y�n}5a>������WB�Xƽ���Eru�sņ�s^s��W���f��-q,̮Gm��p����h�k���C��}m���)p��<�{��Q�I���-̗�b�[�������j���xƗ�Lz��ݙl��:W,4�v.����u1`�F��3t��96�r໅�QԳ���8�Bew4'vlꉇ�w��q��þ�F�,���-b�)яz�1�9O��Ԍ�S�n�` ��:<)�T��<s;s3`/[�X;�9F�2�Gs�W[+;�,)�+��5�.�qq�6c�; ��y��G��X��S{F��o.�=u����b0�Ȼf�Zm,vT�엵zl��MT*$�U�C�U�+<�J�c0^G����uf%��\��Cũ+����RÛeV����~���0�7�TQ_�
�0U�>׈�y���g;�ִ��۾��%k��Վ�V.���r� �R���Y�Іçt��m���g,j��o`��x)��}��Z��b�&��ǌ�Q\*�б��<��!Y	It�(�q��޵����W(��n���^�m����;����&dYi��1`�:N�(�;�5W�YMd�w/K`d����I�;6\��w.X�Ct4Y����%�*�h��h����<���՗�ERyE���y�o�P��{��[�i�7�N����X��d�T��ak7do����%�:>nbrfy��7wM] ZP^X<DȠ=�����=�މ16hBr�S������p6����n�S*Pfľ9�_ʤ�٦��5��QJUy{�l�)��-��W%;�RIv]��� @� 1�$�Yk9R����HL�qL���ʳ)0:��EI-erՙI&����A�*��$�%E�����d�uD:XRa�0�)�R�R�"�'%�P��� �U��+B�H�,Dõ��Qj&���0��2�Y�.GI�EK�(��H�H�p�Q
D��ȫ:h�E�P��$�QB* [��I�m2�\��I!��T ��r��PP���W*��<�j��Q����s���� �.r5,��e�9J%�гbu"�02D�\8l��^V^D,¢5b�%J�
V�D�P��r2*�ʌ@���"��&@TE8˹I�� �%�ˤp��ȉ	"��a�t	8���q9JU�J�-����H�&r�ŉA�˕Br�*��)�v���H�9]�A<�"Ta\��R��h��"��(��{K8�Xrn�{�E�&M�g��l%ӳ}Y��� �69���=�Z�}�5�E&��ty0̾����t�z��U��;����n.�����?�q0�8�BN��o�pr�];��>Q�����ax��m�q�!�?#qS���7�|�������z];H�O<��x�w��D_���j���;��n�w�����������M�	�ۉρ��1����o��?>�����,<���.���y?�����y�t����M��;����������®��[���}[fv����J7� }L>A�y�Ό�������z�۵�z���7�N������ S}BI�o ���1;�|�� x���:v�x��'�+�q��������b#�K��/ٙЩgyo ���Dp�D!�8��`�C��w��=�!�0��?�p=0�of�� ������|q8������7�������/�n'q�wt�|���t�9~v�����d�"�Vn���qC�>���G�=>[��޻��~�to��M��~��6��o�>y�޷���]��~{���״8�_���u�����m�m�N��������ヶw����o�q?R$���1��s�e�C���c�2AO�q0�\)�w�i�{�G�ߞ;�;�����������I�B}v����c�v����O���{ͺ�<r�������\
k�9�}���4b����{v�k����|x��C�1�?8��&��C��n;��'��Np:L*�\,�q�&#��e�?;q��x��;\��>���Sx������ߟ
oP��^u�޽~�N�y�c��"�|yw��[��i�( d(�������;㴛�?����~qҸw��S�|C����{��z��?����&x��q����!�0��uP�7�$� 瑽C�Ǵ��\P<I��N��;=BLg�_�	{�m��B>�DD�|7Kݷ���}���L?�]�N���[�o��'�X��۴���~���Wn�M��7h_o۫N�7���;�>&v���>8���>w�n.�Vm}��(�q�D�:�O���˧>���O��N;|��n�߶��7n���>�O]�"���a���߼���o��Ӥ����;_O�7�<v�qRv�v���c~��Ӯ����ݡ�4'��:����%n;��/TH��^�Y9�4�ڄ{�}~��jtd�)M�;R��/y*ǰ|b�p�k〽�9Ĭ$�f��m��U��؆i��u|ɛ����'/����ɑ���&:Vy��׭ͬ�V��z�3B����:�)�Gw��wW�א���\{�:����:L/�߼=v�F��|��޶��Sx{��޻\�{�t���x��q���`��'�8�'�����0��利s/����.w�x�;���|#G/��𧻓p��y�>1�]�q<�벛��@<C���n�����׽鎁��G��ru�8 g
x���ߑ��'G�p��x��c�/-�.����z�����DH��'��$ߐ�������8�}Bw=I������q7����7O�ݧ};�Ϩ|L=^�y��]۴��/:������w����^[v�&������9�Lqֲ�h�;��G����!�F'q7׏�p|w��0���A�:q��8��@�(�����ˤ���:���o���}9���ny���s��#�=���P��� �\8�����pC��S�s��F?���>���é�X����8���7hO��{�ю�q	����:�1;�x�9m�����qӵF�㗠��i0��G�A����=�ǜ�	��l\�pت�0��Z�ml9ԏ��G��	���* ��P�{�����z���	2���s�=������#�o]�&���;Ƕ:��q:�:N�������;q�q1�H����x��-���q�g��7?��߽�}:N8����uq7��8������9��v���u��A'������;�t�{q7�o���#x��������8���O���OL l9 z�c����G�*�=��V�]�?t �xC; Dy@��G�`��t;x��;O���ǈ]�;��w�6�7��x���z��N�7Ӟ��|wI�����8�>���C��� (���������>�@.k����*�v�~�����v���N�N'��;�[s�5~C����>V籾����z;v����;���1�|O]��;�r�'�g�����Sx��;�޶��z�N|��p�{����s�_��V�-�K��q������yӿ;I��yc��|wN� �M�z�q����N&x��G�?!�OSq���q�y���L��n?�����N�v���η�n&�|���̟���R��\�c������q�g�NL嬧�9��Tỻ
r��,�z�,�HXU�B���Q�͜��۴wLfIR0f>3��溓쏊�(Rn�2ic%: Kg�k�N9)���n�MЂ�R�
�������o�ٲ"��e�Em(u��_`��=�5�����@�I�E�#��{���?�=�.��C��}O���N%q��M�q8��5s�bwhx�'���C�>&x�>[�>�<�	�{���#�`� �U�M+;���)*���Yp��{)ǽ� pN9s����q?���=M/��'=���I���w���>���M�����t�>GI�B��q~s�8��}��,I@�x�GK��ΐ��a���/������#�74>��!>����(����z;C�a����κ���n>�q9���1;����>���>�N������ݡ��?c������b(D���#�{z�D(�C�=������=����ݦ�	��N'����<|v�9�1>�|����Ǵ����w�������iP<��n������y���>;����~��7i&&��7?xF��"$G�#|ǒ�"����}~w��N�4���8�kg�$��;O����;돔s�;q7�O��t�״�]�ռC���y�n���Ӿ;H�u�ξ8\.����$�:q�\���G�!���/v9�'Z��kzM׳���{��1;���u�$?!�q0�������ޡ�w�Wo�r�|����=�|@�'}�#�'on�q�_9�!�i|�����G��P�����#��|G��dW���1,7��w�y����S���;��8H^['����7��x���1���'x�+^�q�'�t��q8㏎�ܺL*좜���&,|�wN��7��Gg�<#��g�[#vdm,�f^koϾ��M�&OC�_��籿!��{(�ۊ��>� I'�ߞ>��÷o��B��=���>��M������]:v�o��8�;�j��Q�C�>c�>{�o�Sr�ޘG�^���ϐ��ݤ	�t{ݕt<{�txLnF�>&|Oy׽c������J�SOn?����($��;=��[}@�'~w���m�t�'�k��_���@ ǽ�(�]n۰iwS��0�����=7����S�����t�Ҹ��'z�W�|�
oS��w�u�bw��|���P�8�g�ߐ�wN��!Ľ�������y�Q�'�LX�}􈈡kM�@��w��^����|M5t���&����}q�{l��:#&���nؽ{0���������(>6�H�Z����r�!%���CN���'�5Dd����ͻܴ���!�t �X�y9���t�$Y�N�4�;)*�������^�<^v
�v���2�{Ot��s���q�ێ�}��:C�����=N�q	��緮ݧN��?w�o���N��F�oP�����Ҹ������7�^F$�{�=M����q��s�����D�;΂�QHy?Fo�3����} .�>������վ~����=&���ҷI�aw���G]�����?��ct���<�ݸ����A��'�ޞ��_]�i7�O�y�[|N+�H�vܨ�ܿ9ܻ�j>Q�#�G�H�G��|�;�j��|o��]�ڣ�=zr�;J���q7����C�nu��8�������u��|O�?����y��ަ��'���>� �+��}�˼��ۿ.�
kSS����  ǽ=�ζ���;q7��=�'N״����t��$���{~<�0t��
_�.HuݺM�q8����p)�O��|�~M����Ӥ��!����_���M]��D��2ﺋ��%��|�G��;�9�;�+��'|��������R�Q�'!s���X����^�集�+B1xn��d�������~�S�m]>'��L��W�R|��ehj�O_��f��"�ك̘28���s��e���8��Z'�Z��ճ��/sq�E^���r�8:�g�7W�UQ�)���������H~�R��"3(!^��Ӊٔ_0<'�,p
�o��"���V�V�[���E�ε��gz8���{t�����vY)X3�;!P����ujC���A�{*�w�yr�FbO�7$�ҹN�[�\��q�r������p���Es��^�`f���I�/D۫��2h����S���Q�&�sp��p2�Ǫ�X��ǁ��s���uf�����q�)�������V�^��~�b2r7��n�u����fС�AyO��s�v��e�5��CاZ�+��� �:�����;p��\Wn�3�I(�D,n��C��+O�<�c���q��o�`�d���K��o���ε���޾�r����:-\��"��k˕�-��Ɵ8�y�Xs8�PQ�Ф2-K}	ڷ�W����h�ئy�j���R��G,t���cOX�8�������)��s�A����@�e�@�a �������GFM_�����ST�ꨮ�8�ڭD���N�,�@�o����i|��Y��\����]��y!o�;�E�)�gA��܃�寉�A�C&�m��[�bh�����b})�e�F{��}L�\�uڌ>����`otP�j�&�u�^C����UJt�@�L�;>=8��f���9EuuR��ykC*�)���ѿ>���{~�&��,�ɣa7Q�L��II�8������̛��z�1��7�z�β�mEF��˯,,�����g̗e�a��8"#���xv:KY���X����3��"6}!uČ�D<9֫I��P��h�8���s����-H�|�:�oU}O`�"3ʻ�N�s�K�X���mo����6�����Og�&ٓ�E:-�[���Q��A6��[�%�P���{ۅ����B��Ժ�h�����i��޽aN�9p�*�9x#�v:�������0���wh/�c��gG�y�'��Ϲ���r*͚�n i��3�HW/�+�hj�1��C�YEp��V^Q��=ީ���l{�_
5�6�};�L��2���߁
�P������dO��Bg��m�%0D:�vb�<�6L8�x&�]��e�1`��Z�C��sE��L�IB�ǈf�:�F��b��	O2�|���Y|F��s���tܝ�E��:�<im���\k�w"����U̸wS:�X�uB�>]���"xm5�=oޟd�UzN˔�[�1��Soe��hi�d͓X2�(	��ѷu<o�ED���ǯXt�3��3�r%T��W3s<ל��g��ڷkO��k��{~���:>t�ϕv�mR�WN�Nk��}ɏl��Z�:Ԟ��j�׫څ�Dt:�a�\�hG��!��i7�y���tt���AX�����&�;P������>;�:Q�ߞ�1��T�iJ<��@i��xouI���WVf<n�n�i
�=��4���I�G��l��d�؋r��*:JF�U�|��i�s��k�RQ�+�$�b��"�:�w;2�&��/�R�-�bݺ
����;��=W�'������ݹ�[�9C����zg�{�N�[ݦ�����vc΍��TL�6��N�2��Y�U��O�l�G�S��Q�G�9(�� +���ѣ0M���r3 �<�����[��Ͳ^k")M�c��*�iq��Z���)E��U;���B�[���zL&�RE$��-�1�|νu,�:[Ț/�ZY<0�r
�
�E��]��}]�}�ozD(�
�F}졦%�5fI��[�9/}ؼ/�X��zڱ�<ڵ�҃c�ā��E����i���Qfnr;����
��c��*`��4��HЧ��&�0o�ݠ�
�h������6n]>p^�4�4ll?v�F�;��3	�.���N0��)\�[.��p�[�X�s\bi�4*�5�U#f��Q�v@�����J��Y;�[j���o�vFC����YM�{S�ǣs׸00:Ͼ�Ϧ�{NDJ�}<ʈW����pq�&T�t��a,�x=�P�w�y���:1^���W�n��F
��SKc�8�aCt_?�m�|>��h��9�;���ו���Ë���|��4�m�,P��QZ�F��>Һt�����,5�4a��
#��M�Bl�/s�.l�����]ey�������)@���M� aMе�Cm#oq�.~$fp]���K����wŽg�]���j�@Nw"K�K��&��O�z�Xv��m�+Ƌ�p���EH�����'W��b���o.>��!FX�Ql7~zT��.���x��>|B�FR<�w/6E\�b��ΗQ:�B*���>j]<8RY~�Q�kC'�'ޔ'� j#�x���;Bn��.|�U$�"�1��yW�mX�2�q��8�9�� m<w1�N��3�2��a=�y��j̝�i.^��.f ��^�G�X������
��Fzl�p�t'Ȗ3::έ����y��|�W�$�c�LB6LHyt�X�!�_�p�)���K�Z�϶�\�m}�j�����F�q�	�t%�^G%�}(-�MEȻM)����+0�����ʮzsy1����0��;e���yF�O�t�N��0���yB���ӃnC���Ύ�r�Ř���h�gvZ��ԕ�."&\F������q�?nF�u6�"xm�쪬
[�h]O��\_)/n�I�a�΢�\���/�ɜ�C���)w(Q�o��ӆc���Y��}�;֍T�|O�c:����Ɋ�V���<pL-��3�;^�>�5�hÌ��U点|2n/]���4�\��� ����fॏ��ݧ��_��)S�EW �Ojz�_ݍd��֠x��Sr�]մkb�^k0�� O6�S�|%�/L�KwF,���{�,�'D;4��3����r�o����ҟA+���𝧢��]Π(6qD��B�1���(��x�r�iDU�X*���b��s�:^fzާ�ĳV�y,6W���|jV]��}\h��U�U
��������>8��A�� dX��0��v%Q��ʩ#خ��o��to\��Or�\I�
9��!&SL
��ӝ��lJ�GG��og���n�r�_�v-����['���hgoިg9no;2��_n����#�4�݅��t��yõ��dX���⭾���d���� �r�c�6�����꽻b2�+2�Qc�AF�QQ4�[�jK/�i�<�
-��.�5C��mȑ����}{7��,� @Xp�����3��ziˎ��X�qC�ƞ�,*�"�a2�+�I9�H|���~���jP�ޣ1
D���ϧ0q�k��������c�/�#�ʇ9�^]�G&�{��ȶWq/]	�މg��DKN�K�z�f�z��]մ&�c�C��,��}6��biG��;���'�.:ۭ������� �#L\��D��;[tp������q�d���$��;ݠ,Y�5��Mk��������w�U�`���5f.J���j2��@�J7��呾����ܚZ+sL֏F�����bs����\�5v�ض�������ne��Ƀ0]+��/���u���i�Cs���_�W�(��9Pd�n���DlXD\BK���r_0Gx��F��N��g>�}���sHN�:�E0CGh���'��MQ�Y)�F����x���:FZ��[�d��Q�+�S��HfZ��۞�ȇ۔��V�����=����s�M���t�b��x�پs�b��!�K�L��*��׬�{9�5/C���ݞf��'�)��������-
���^�U��sT� ����B��W����srp��S�a.��|�f�Gz�z���`�o���{�nA��ܲfx�2-W�nr7ratlQ�e����%;d��H؈�}F9
��];��ʘ�V_��@�;ky�vDede̊5��V1�ڭ6���.��A)�_hy~p��n󠣳���u��ĉ�X��EDB��)'�C�UEyk�!�\D2����V
n��Xw�ü옞���r2r��0,��W ��pik�2G���S	�vz8���E��ܗhDd�����Og�:%t���z���W�{nK�3���/�.���3M:�����je��>�˽9华�EU�r�N�m��i���F�ޞ���YLS3)V�m>oz�OQ�����(3u���Bs�M�I��I��M.ɹ���)h^̔�����w�Dt���Y7ޗt�!>�.�9�q$ch)=�7���T�3{q��3�̙���(���oy,��cK��T�i���n!�F�Չ�&�v��	�s�m�|��4�z6�m���i`�5'ل�}j��*e1$�T��9�g��B��`K�ê`�|栌Uu�F�}��t���ot�R�d��ñ,XꍩK�޷|;�̋\^�W�^�-�LjV�F�2�1����������u����ߛ:�.F;	9���]����+l/����R �vj�4�1�!	��Z�c�@���z�ЦS��[Sͳ���b��[͊�V�d_,�v�;�������k�x� ��p�:�mqn��Y��8d�EN��'٥W)��8܌Lΰ���)ձs�o��ݨ'$���\���2�]D=�� �.��B:��ּ�J�v�����M��z�nly�X3z����n�˷F���4�Ή��sjԑ��(��d�2�mt��h�s�4z�V2�1�3f�}�n�J�e�N'qWd�3(v$���"35��Gs��G}��	zG�o9Kx�]��Uׂ3̟fW+������#�1ݘ0�p2ć|�;��Z�"��z�E��{�����:��'�U]��94�)"�Y{�a�j�6���k���JG���M�0��\MN�{�����o17o�w�A����Q��OϔEU���ɚ�x��{Z-������w��[lt���ݑ���������,y'�*�۝������v��U
�w|�q5�	t��^5�������t�w㻺 #����ȋ]J�	X�]j�QIU�+n�@��2�j��&����m���[�5�#��]Y���MW���\��|�����2 �ӭt8����W|D�^���A�.닅�yXA�@E	a��e��N}�T�cM
��v�/����XXO.���� �C(�w�{�?D	�ޮ\���s5
������:ڧ��[��)S���6��y[�{WkI�E�$�p9��̵|�:��ј�띑�[
x�����{��}۸xr���7WKƾ��;j�+]gg+J������M(�kwVJ�ۚ��o���c؈���U�6��	�؞K����6r����l�{�D����|sv�=��e
���cf}ɯ������Z�I䲝�חo��'�|�rK����0�̼Y�p���Ͷ��"�P���9T���P��Tv��y��i^W=�է�V�I�;�d�L�:}�J9W����Oܭ7�N��7�mt��1�8�i��?������"�Aݲ�˔�	�
es���2#&�,��PSd^2q��Ud�Z�2�A(��eV��-X���S���9B�+���W��PPn<yi\�V�"�YZ����#�QTD�)��rbʨ��h	Q*��K�ʅH�TEA��͔E\�+��<PUU�NiQ��Jak��er�#�1�r(��9�0�M((�+�ɖ���s�Ux�+�A��Y�9DU�w#��pY�"���˸�"I8x�<�!�Qe
�˦s��QU3R�)VQJ�]°��fL����\ΐ�DE��xȮDN-�)W"
��E!#�)v��q�H�+*9E\q�q�*�[�p�r�U�Ъ��˕�p�(����Qr3.\�
eEB�ʈ�(����I�EWr��9�"�.�> W�
�@���Y�����o[�S�O8\�Y�+z��0i��.��V�k�t���na�a���7�$��n�3���.������bm�R�ˈ�ԕ��SZ�Fy$�xʈt�<k���#���N�c�����q��Lm����#Y�9�GA�A�v�Y��ޟD��ZM�y����㸜U��np�\8��!z���`:v:/�NS���G`=�c)�(��*k�@i�|�-�vMa�;s
S�{���2�=��oD�@I�G s;���d�dG9�|�IQc�*�g����On��C,�K�$De@�%��͂��F$�ܛNG@q�%�F�!�˝�W��V�jo�V����X�${b����=*:�!��Yq�E�JҹɇL�$���h[�kRk�l�{�U:§\rO��:������]X�[��.�p��'�&=ꕪʴ��VN����;qf�'."Ms��V������!p;�ś��T�mR�to2�� �z��*�a�Y趪���P�2&��NEE�F�X�e;�]��Se_Aټ�ugOm$3'�"��L��S�C�8�j�N��:-���6E��X:��z9u͇��f`&ct�I�M˦��ȥ��zs�c#ڸ�kV���%����n�S<Vz��+x�z�a�Wd�ɛ�{u���-�b��S��k�Dp[�������*�7����a�9�Wu�.7�K�'���XJØT�f�7�B���{�X��ok^�
O���l�Ν5<�G�c���e�&-�������=س�K#�%̍�l����𡦘�y7>K��K�iy�iT>�;*!��jS̸.�3�q���Y��]<����+�0l1�]u#+�`�<%4�)��8��L{�g��J;�u�'�D7wX���kU|�1�[=���t��5������k�)��eυs\73�=��mc׻;�۸7Udb(�S����鰫+�
%�%Q�>!OC���ۢLF���?������=��ye؞6"�ϑR�K#�QKޙ������)���7:�3�@zj�{+�Ɛ5�d( =.�*����b���x!�i�� m�r��}���-��e��x��S����i�f!L7^�	����\ioWG)t�9���# GT�ul�}�[���F�	Ǖ\f(t�F��I���'�ME�Re�
�my.�
5�ln�656�=I��O�zDp�K�C�xoԾ�Γ�+��A*�O��4���c=��V��믨	��!�����5�z3�ӌK^�r'��R��|=|ō�2�r�m�y�Kv�ƌ��ټ¥�\_
�>}�,���+��;�
����{QLb��hi
���G��<�"��l��g�^�ӬLu�Ě��g�%ڌ��(��K"��B�����  i¥Ә���1�Ѳ}�ܕ2^C��=F}�tEh�r�;>�Mv���9bv*&"a���z�r��Х�6��8�&���(��ix�����'���<�����Ƣb�{��3W
��G����_M���$�b�u�˾Xr����a�a�:7��L��r���^_5� �Qض#'�@Mӌ����)���W��R|��ekWbxƨ�H��r��M��d�\.)��&���j�AS�}^������E^���r�8�N}�7��]�ܶM��Qbz��Mȫ���e��8�2���^����vB��P���F�^z�]���g���p �%~��+<l'��c{*x�2R���|����������xa[ ��=�_�̌�!@�RGaԧ����ЃU���72ބ @\�O��ձ���3��
��H�5��&V���9�ӱ��;	�r�8�U�в�t�5���R7����]����s90�b�Y/�AF�QQ5����g!{�b͡ѣ�?s�M�S�ќ���?%�s�z��N�C&r,cge{�gQ�5�}��5e<f����f�����b��iW��n��>T�<����U�5oe�c�
<�ߔ}n����q|���"á�>��=Ȍ�f�%���$ĝ��G7_�,nTa�F7�x %Vs���hͳ��p�( h�%#gA��Wt�c��3��zh9qё|��E��2�4��ma���#��>��$�{��ޠ�9B�b�<�sP)k����L%9�X� Lf�w=�=s�э���EF�;������ϥ��:H�;��k�œ��⚘�P��w�s&B׽b#"�j�`r�.d2kͺwg�Ʋ��*+w��F7w�3=���ʢ��;W����E�T)��}�����W7���NK�F�5M���]S�G�ϲ�/j�?���%q�{~��
d��&�#�3U"��+�|��qg!/��J�"K
G�6�Ss���έ�Otpv�.W_��&
~x��[��=[�񇸡�)ͮ�� �s����U����)_m
�
���`QO:�C�o֑]��5؉Jۻ\�j�+�;s�N��X5ףh=�f�r[��������qܯ1�u�LTs��+w�T0Ke�Q�"+vGC���`��~�*�rct�{q��F�����]�/��Nę�e�wA�W���S���+\V�ld����$`ՓDs����ә�i]�C��	�K�+�h��d�b�G�r*�32 Lǣf���QY]�p�L&,�yӟr���1�s���t����t�q��TUw��E��������A�T����������=�2������D����\��8\}6���a���Μ�*�'�	���_%���+l�*�ߩ�3}rF��b�.4S̾ח�
�|F�:
)��m��}UM;|���9�I"|OC�"ga�L��~j�H�-u�q��r!��Ӕ�UvcJ�2�>�����_L54�N�>.�"2��>��%�F6��mu�a:����g"��񱯒uy���ť	���j��SZϮ*�	:`�1�r#n�%ybH=�v�K!^�Ԯ:�*.J���h��0�#����x"�B<7��B$�L�(���l��o$=�h3�}�@=}b�Ν��NS㺝(�^�b����O�<��̜����z�f�w��/��B���ӃpsK̉��@-�PI�G<�vg /k ��"��tY���^w[��̞���P� �㢘���f2��#zԺ����
sl��s�`�5�T��9]����o����d&:n3Ҥ8��.;H�;�i�:0�Ƥ���B�[�������vG���'}�$�O^���|��pNgA�0+hK,������p�۫XI��L�p!�d׮�R{ڃ)9�7L�{�y>�M(j���{m�Uͫg�ʐ��˚D�^db����F-a赌��2��$u-��x�C�Ms�g~���xt�>�[w��J�2~} oZ4,V˲�u���-}�CMv��-��u��a,
'M	Li�:$��������vkhxw��O��/|�|��[@���uеK�D�P�9���u7�:�S�*u�HF��;����.,%T�Z�P�[�P�f����wS!y�3�sr,�E�M^�V��P�+)3f�d��l�l��q��	�T�4p5t'_쾎$�������S"*p�/�-�2C'��9k*�߁�l�cH;Xx��e��*1�mW��S�֐z�Q�n�ҿ���;�!�ߑ�r��A/��#`.Cش<�6��u�'��-�r-��~NG�V��t��:�v�W��n��2�`�<%4�+!Ƕ�&=�>Y�\�+M�ږ1�>���C{Je3��t4L_�]�(ز"Ǔ6�(�T�q<Sܛ�`�b佯��e
�vح�����Hq�1�C�n��ڬ���rQ�x��ς3U��3��#�����]ըQ��LE�v%�Kgȩvw�Idn9�xx=���߽,h�L�0ϼ��hC�4�p�]�(3�`ؓ8/ tx�n��5�DE�lV������1X�_;A�����P-��֩�����y�S�Z��[1@��z.52B�q�+H5�)�r���	|�ʀ7��,�i��{PB�4(��+�5�%J&O�.���'�{��X�zݶ�2b���q߽�W�y[V*���l!�i�'7t���rӖ+��9�|���X�_t�Te�&`��4�bJ}3�/�Bⷧ�yS��� ��E��U�Bbk
ݙM��}�Ǖ½;+�k~(>H�|�Ά"#������i^�G�uuA.���)¼��.��G�_��N'�*@q�'A#�=dp����ܮ4�{NW�m^,��x=����c=���3�}C��K�\F�`\D�@��D걗�����"P���2/�{"q~��f��a��������x\D8����/���^D��z�U�f��.�J���^�K�����k`�3���Hؽ5$갰��C�2K�����*��W����j^sc�jO;1z�z�b��B���~+c�'M��^ΟJ*C�918�N@����T���2��w�i_�X��fa�5n�p�j�F��P������/Z��3Wf�-Sۍo��u�n�I�u����Dm�Ν�"#2�����sXo�Ҩ�
����� mo	z\�cDv�n����-Y`ǀ�yJȆ_4��b���r{}�O���;>>�$ƽuY�c�>P�b���Zek:�U�a��Y˒��a�`9M�t)��3��֫}�gG��r;]�-uܾw`5���wu/� ��-h%4�Z���n[�<��FT�N�هS��޹�=�,��Ϯ"0W=��Dߡh��S<2t�갑�\ڈՑ�P��ܘXu���\�8�U��rކ c+<lySDU�i>�{Ȯ�Y��T��֐�ij� �t��8yc�ȱ-S��*��O3����7��8H~��I��ʈ�]A�L�_\��x"��h.V�皒��|�ZUSw�V�f\�������cՉ_�`>.���V�|���c}�~�'������%~x�jze�6��5�e�{��ь�ː�r���{�F��bZLP���MD`�d���t�{��6፮w�����]��b%�(��0!*��A�=F�8�N����5�X�X�w>�q�5j1ˤH�q�ɦ�lE��4,��ME�\�cg>I
�VS�~��v�w_�W�(���T5��t�8��P*#�Pd�Dkp�u��Si��(���1g��7���;�q������Jdѿ&�#��qާ�wV���MP�V\��o0�Gu���.���vcgj�2_K��"eQ�LG�0F�~�4�;գ�kHx���i_�uQb�~~�BcVwIJ�n񶴾�O�#<������M������r���bD89j����=�x{��:�y��:ȲO����T8�u���Km� �ޅ�S�L���f���zcz[��}�D:��� ��1PU�ʳ�p#!h!�ȡ֫I3eCX�:����'կ�;ϩv\�8��}�eY�\����3�eXHW������{i!]�t���n��f]ޗ�!K���^�	���9��^�2�/�!+�.�Y�7M�J�-Ց��g͏��V�����";Q�΃dÁoe>����WE���#dLl��c6�f�D�k/���uH��6��8d�u����9����6wC��>�3�	�Ne�h�q�J�}�Y/ ����%��SKڪl�����O�y�ND2�<MYj�҂�vΨ����������50��GO�":+���\	գv�)��ED��	�j�=����n��7x�R�����j����}b*�p����wI��]��m����M��"�o��>�~ɷ���,J��6���c�r:��}%�� �T5B4o�v�F	J�c��(!��-�j(uL�P»j�;�!���������+"�I��@��'с�-�\{��LB��giѣ�J�ot�a�S����'T�W�={���r����p���v�%���jrS��L)f�k9F�\]��U�0@�99�����������m7�)�'�NqX�}��_X�ӱ�jr�Н(�m�@:�Jd����#�	�{��m��LDaFG��:�6�`>\yoEz����{�g`6s��U�������T��Afx�$�g�_@4I9$�H�>��@�%i��e3q�j]NO'#�8#qs�B��б�G����W�N{�r�$>��R�vudC�����X��F�,Z:��u��9����ٓi��qu)�/YD��w*�����i��ubU�~��E��˖L�8����)�c6��/�;����9�	ˈ�\�#�5�@���v��m�T�6_8G8mF�[������ˀ� ޷�������a�dL)�a9:�(�b��D��;z�l��+aYe*�e4bH���L���� ��k�8��3���v�P�V9 ����m��v_�\"�Vh�!X���`��%; H�}a焩�e��*1��nE�n9����[;�3��W=~�E+ڝ��ĸ[	}��_1�WGՊ�)UV����"aVc�~̠�oӵg�G.@{�5��lĎd�_)�G�w�H(��en�;ՙk\S�U�������w�u�����}��+����@֧��U2���q� dt����k��s�&��l��{3�vJ���8��oi��˾7��~�<N��\��U�jj�K�s�4�b��C ��bpr����}Q�P"ֈxX�P��jT�r�K�[��ܷZ�b� ,��s�-�c�t�w#Ĭ����&�.kB~Mxn��}�[��M��.���3{��c��$<V���T��Za��x�;z��pU/����[�jQ��kd��q֯lK�����wn���=Vby�}}3C�k3�ܱ�f������ͻw��vL�U
��u��Tң{��y�Wl�h�9��)W2V���׉����j��[5�.ǧ����p������D3}����(�tE�p7�M[o���"�2r��}�:٨sPv"��ڔ��^L��N1�璋��{�s�n�h �s�'Ζ]��iX�FY0C��2�ӎ����i^���g�%iAg���
�W7Ӎ��9JV-�69-��+��^�>����ˇ��cz�Vf�ȢW ���D��s�	�N�&�oa����̎ټ&��`>Dm]��p9�9J.�ǵ��@d����<p�t�!��ݣ*ݠ�t�F6��c[q���F��ԓ%39&Ü+p]�vm�o�e�6
R �E(�lH����f�<U!'�l��@꽭Uj�ugNm����:D�{��90&�#{��ޒ��A�n�h ���{+�7Z�+]iѤ3kX�:��k˃#>�{uG�u��s��	���Q{��Г0p�N2Z�@k$����r[x����D=��K�z��y$T�f\:�?�o��u6��/{�b�>��_^���G:�Ap�/�-+n�V�� ���/q��[����|r�8XWI ����i���w��`Tᅻ:���ǌ�o�Of�0�)GYj{�U7����#�]�%���á0�������A|�}Z�;4*`M�Q���]�,�40�����[p-�foR�x�ģ� �؃<�-;@��j��	c�;��)�0�q������Igbw�08vp�V�x#y��soq���6]ީ��H�3#�jצ}V�)9�A��7繂At�ANQ�"c�v�xm�C̻��2�t�q�*B�s)/��sTN�=�!�ZӳS��_�T{w�񕦝` �a;�8>�i�os� ��=�WL��Y]�gC��H2�uD��j)Iڍ���/��y�q����_ol%�8D�f��Y��b��ќ��h�f;���҃3�i�������+���'�<y��xR$���l��[ڔ��	�A��y|x�g�|�!��Rv�;�u1N�:����m�s���O�x�}����Y�V���r����LP��*�@Q	�Q��r̹��
%"�t�G(\
���2(ΐB��
�"��A�EDI%�TUp�Z�(���օr��Њ"�r���p(�2@���FQ�**���U2�.r�.��%��
��HAr���9�"��%\�QW<�9AL����I��9A�uC�T��dEQp�6�UD�QE�T,�8AQ29p�����Q3��r��\�I�\���.*AȤ��L(�	��Ar�2B�;"(����f�Vr���NUs��!*
MK3��&x��r�+�r�p�����E\̉�\�TU�(("9�D�`�p��I&�DQą%�.r"	�TY$Qr;)+�DTȊ(��*��\U��#����G(��;���~��b�<�9ژ�����[J�����vk2z�"d�Grɠ�p�s�y�'f7Q9Ҕ,�l!}�R�Ks
��jƭ_������W�+��7�A��H������[���
��+�u@�<'�/
u�����>�ۙ�L���_�������t�6S;.v13�.��tYd��QZ�Lz���w�wP�H��UP9Ʒ{�Hq����w���+�
%�<ISQ�0L]2���gi+�(z��b��+ �����R��Ƥ�6����z�6��ߙճ���M۴�f��,�����/�*�B����n�VՊ�e��`!�i�� jj�	+�1i�.�'�'�����^��#O�BU�)���z�;;l�-��pU��4y8��g��+	����Bq̳0�(�R`*�`�>���!��+ÌA��
#�f5��~���ٯ���-Yg#)��`T�M2���Ȟ7�
߰;�
�'{��OV�N�9�J!g9����fXg����K@C��(���N��>�����*ɽ�a����g$��+i���!F���p;����q��8���瑚��^� 4���e��y_�s�9�����oP�ߌ�1!-Ʋ`�ػ'7��^��[+�%��;�����Q���N��01,��ሪN�X)rynB�ŏ�w��Mϡ"	�����^+�	N�;�pŁ���������W�[g�^�B��`������9EiZ{yVS��n�g��DxU�c�B�V�p���U.�N�C^L�:D��լ���чz�3��߯�x�nVnmʋD���m�f������k��j&����-X�m����nV�(�VP��\�m
�5�KzܞX6�;:�g�7W��DX�ʝ*E�5�(W��n'g�۹7��������a7����0z�o�A}��KxN��!��-��̂�;���	@p�3��ۮ�x"�jHU@�D�j��U=�Ɏ����<�_��C��m��]Ln�t�+A��������I4\�ƌ��$.;(�U�Y���i�;	�r�8��/�d��H�읽ge����I��%�*��4��� �H���ʞ��,�:��7��)b%oO]��y~Q�۰��^z�E���J����4����T���װ�KZ6��1�3P�O��n͛����r��a�o��kθWJ/h���<���C'}��~�H��VV�A�]
}q�/����g�*��s�{	Y]���~�rc���_]����H�>�=����Y�i�����\:��.#�]MK{NջN:m��h6@�,rb[{8mlݳڃ��W)D\砾��ٍs�3������t���S�"�͝���5~�3�\js�O=v'M��}(�FG�D�#l^VF���Nm�&�m��QtC���im�����×H�`C��Knr#|�ؚGR�6���<2�l�w|�P�u��bg*7E�ھ���P��A���y�>�/ ,o�\�M��(��0L������LK��#|Y���v��gh����{~MH1�%2h�n�nM-��͹�1߻g '{b�yU�Wګ��g�_��6��ֻ��8;��r�om7U[�FՍY��ZC9�%�b%?x�c5]���WJ��
�
�Z�'ِ�U�"���y�֔���Ѹ�j^�Z�4�c]z6��EŬʜ6�N�>s0�웫n�5R]��k�e�v:-�/]!K���^���ݛrE�JD�Y��$7��;�R̫ٮ��K�y׍���'A
"b�1by�l�.>�MW@��WB{�^L���GvU�-���]$1E���&^���Q�� 4cK��JG�z����`y3F-l�S��r�<�F��GN�2zQK.�1��]yt�=�|�z����}x T6ހ��9�=�Or���[,���W�r������.�M���y��n�6u��]�����;6k[����r�P�F�tX�^�_7F�Ӏ�A�9r��������;����:$�j�U���Pnn�� �OB�,���,u��"��^W��W{�R�\�ͥ۵��R�eq\R<��NUz_��E-� �+�T�pikћ���pybT9�����{���_m���aҌ��pmX|�� L	$�+�_�HU��mx�+ꐑו/ܠA?^KAwj���ܺ:��2�*�au]ӥuЈ�>��"���}�,�VV��4���;�@���}б�
n���S����Ga��TK��y
����~��Gq��P���H��ź�7iy�'ˍ�^�$�#�s;�������|�3k��~��������q���1�$譩/��� �GE�`�x��5{����̀�)j;{�d��jg�d�f�=��Ȅi],�[���a�U���|7M��xVvVܸq��#��%=��=�pn
��٢�#B�l�1�����dT���T�d~N��Ҧ�˧]���8�����;����9�9qk�� o�@�^'��n�v��?6h��z�� �%��f8�o�1�U6�^�/��b�K�z8�]-�����/�N)��˦�ߐ��FE�+F�Ê���ގ[g�̂�g�PEص�O�!��Pnۭ���k�|`[�]�t�Μ�F��Q�H��V0�^�P������C7]��wG�	�xo��@}�޷>]��T���x��Lyb��Tí����M�ȼ�NQ��G9��i!h�q�X;�:�)�02�v�g6��0�ʜ�U"r�TL�����U˯j����c��y~�2}�>V:S����|J8���>�5̲bVK7:�Ug��n�uQXy�Wo*��qw���;��s���Z��W��"�G8�ʩ��ڨ�~z�ŀ��_���o��q�
�j�%��;X����˽5:�%c��Ρ��-���O����7ںʝ��=缹���ث~����u8�H���Z�+��^0�c9����+�������S�]��Q��hDAf���Io�����l�R�5b��y�,�S�,��iQX�JSQ���A`�Bc�u��T�h/��,}��1d>��w�{%x_=���Zr��#AS�ހ�[И:ms� o�9S��2�����0��FTf�;��+Ʋ��N��7e>��M[.�n#v�XP�������ırL��:w�l)�CW0T$���x�#��"�P��^�vs�f�u=EX�kw�l��*^�I���w���s��c[P;����s���*_��{��S�*��F7+��$�C܊���,�0��0�ذy�ԭy�d��7�uT�����N��A.i��hx�[6�c�;B:�Wxa��tF��9d�'P����궔Sm{����ܡ�	��;��h�N��Q���Y�:ANM3h�G�zE�:�4���\�o5m������M�v�����+3��VrNN�8_��n�jћY��)k��[{4�'Z��5�L;�Qn����x����T՛��8[��SmmM�l���/g�^���|���NǏTvcI�k<���{�A]���3(�E�?�V�-�QG׏e���.�D.�'�o����=G��5ݭ�R"B�d��*�Ӯ�v���ੱ�7n��ʶ"xr�Ď��G�7�5a�n�O:���N;��u�c�U��sE[�Ci�*�/e��6Z��R�oq�|s�ρ���G�͗&�F�D���2x��H^>��˕�w(�G��*��yKue�	�^��[;�x�S_�^�ϑjd����^�K~�P�7$$�;���R�\*��8��q�Ҟ�t�ڎ�5������U�w�ٲ�z�o4�^,�BNP��_W��	��Tڷ��
ȍ�yϠ�%��,S�ѭ��偍>��A�57.n�w��Z����]b*؍��ʄ��mI��WT�4��m�Sr��V�Q�y/31���ގ�Y�m�7b*����@�t�uJdC�[mbYysO�/V�[��s�,���/�lK��*{z�B[}��yo��q�w�8�����	<�5���9�s���<g(,�0�w���yM뉛�t��q�\�t��+b9�[щ4�e�0��n¤g�Z�t�B�%&����Q8X��^���+nw9��F�.f�M�;�61����bZ�wc+���
���z���7�b��熤�����4�����w���5��b{�h�׵��"-mz��y����2�m˼+;�c��[����f��Ƶ�/9���P׆�\tŮ��T%�	j"/r#�mb�t�^-�[����xc�4����#��rUs��؇"��-��^ߔxgV���8t�T3�=��f_��]���3� ��)ǖ�K�������跅}�ׇ�Rc������V�9u����d��pNp��}	�yT�	��/�]���Mp�Y8�r_x�x9k��:�#67qw׵nҗ�����b˞�5}|&|���R�-�v�b&mo$(�o�z%�e��+>*^E�z�>���to����Y|�K�u���7��n:���.��7/X	��d�+��fU[i޼�W9l[��S���w0w�\�m Ո���.o.��7�Z�ϻM��Z�q��藻�j�9؍�| �$��m R�Ԯt����ի���s�d�5Ϯ6���Y~M>�i턯_ݰ�`�t=��݃�෯���FM�W��:���3>q��5�v%��vc8��S��T)[�
%9�5���}Ma��X����ʤ�+%)��Z����O8��P�ю��$��\X�J�󽴖�$��"��K�GԵ����#��<�lS�rdGIs;�q!*�r���b�d��� @���]h˩oFRM'���D�h�]���#o7����;�<("�̬ۖ�8����/4f�,�r��(Z�Ӝ�rJ=�@�=Գ�c5��z ��Zu��z�n��h����ѻ�U"�J�\�4D
������TVčNuǛ��@dgnVW[̶��oHV;�f��j �3Z�[]�q~���;W�����Q���u�#�t�Cb�}4%nf�|��j�ݝ>�[K��T�Y*Op�C��¸v��6%R��GhA�:��k�O�Mm,ۜ[����f��M��M��h؟k�9F�Z����6����Y���hfN���o5m.�W�N����y�tc�8����U��n�w����2���K��Z������[���a���S�7��@X�NZ�R�f�LQzx���Yg���nM�V��B�8E�rx��,c����Y����Q���Α�qw�܈�M�P�1	�|�pX��c��wf��}\�Gf�~u����~�8�BU=im5n�-����e�x��9��������
w�J��oVu���U�FJqO���n)�X�L���U��W�R�o,6�X�ϭNuWB;۬�Ѳ=o_������.C�v�.vHw%�F�63b�j�lv�r���Q�4vjC%嗨���Y�r�e�Փ�z�d�{�Lr�nk=�K_�3����#G�>�Y�8�����M��kR��
O	2A���`�ͩ�ɏ�]*=�Js�����<�^$[yx��ރj��U�JU�T��}�7������)Ȋ��$�3�DZ�=j�զ�`�>�=�`�py�Զh)O/�C[x���WD�L-��:2�DJ��(�ܥ��r���$(Gv��K�S�9}�ƫ�\)������\��2�|3h,g*]"�����O�G��AP��t��n�5���l�V�k=�m����t�T#`�y��C`��[���̧\bOR���F��&_C�x�[6'ʑ�(�A��s��<3crHV���N�M��˔:O����~��;FĄ��!����(�~��w"�Y�W��>�V��
kW;}��XÚM�n#ˎ��TօJ��'u�xb}�:DZ����R�+)k�s���������Rǣ|�sl<e��()��q���:5�ㅾ�����P�[/;�����B��~پMe���p9ӓ�0�2��۳Z�r�׮�su��jw�<�����C��#�az�hJtQ.�`�L��1��nں#��֝n�`�ɫ��U�i�05�t�.��2�-HG���"�{АŘy�ó�
;������,r�W�:�)�2���4��}:�ݖ� b��=	��K݈xoi`�ю�[>o��&o3����K�:��U�
��슳2���֯f��\A��|z��ѡ�6�E�Xu���p�Ս�C�Џ�ZU���Q]��!H�t���ݣz���fh>�٪�e��p�6葇j`���z�]�����B���d��
jZ8��g���K��K���z32b�B�8 � x���ZʥC��-�N˻��9ך%�:�sd�ŗE�t�YІStv�Z�Ŗ�v�~��tNz�*���{GH�j�c������̾�Ǚ�	�;8�كH7�
U�ʸ��sW/�I�q1�Qz7�j�Y�u�4ޞ�t�o��V�VS�E���-��^�����zĻ�Xˏ3�%�;F��z�n �KLW]yͷ���F�.��{��3�V(+��>�Xce���a������C���2�D�:,�&V�[�kMa�,�1�hY��'Ky����v/C�Ŭ
��ȄhN�7�PB愵Q%�ՙӑ��on�]����CAޒƅ˜����w�U����B?q�ml��iM��1Դ��wh�,G��A/:2����/��{�(�RE��N�Q[���0�n[�ݧ��~�L��vd�Wp��F��.�:)tN��'�Ϧ���m���\l񫖊��fP�bI�(m.�%��h�o�q����)�����C*��g��d0�j��{ٶ��z�д���(<�Y(:;�����|h�mt�"kzz������V ���^�~�B1*8��M���V��'%�ʗTľb�Jh.��b����w��,!N��w(lKw��	���L��8A�M�v��L�5r�*��k�`,��o�͙��S��T<ZLwL�;�"n�N��K��$V�B	�}��6��b�����$+=�^.����C���h����@�ru�z�.SAy�tn�U���X��\}.������x67;��������ɟcz\�I��7�E�9f}���}��a�2�����Ŕh�fY���+�2���Ũd�4��3|��}!���Ӛ������@�aimYp�ů6�yk���S�Ӝ���7�<�mؓU$M<���9J^�-P���d�,����ׯ�w�k]��P�0��L�m9 �a��0�`[���1}R,Y��N�	��܆o��Ξބ8���1u��{�9+*��/�;�DOU՗�}���[:����i;HR='�Q~7�U���쏉��(mj�vQ�vm��o�Se��FL��Z�\�r��3����TBt���PEW"Vң��B��R�B���3���*��Q�jD5*"I.b�\��"$�dV�QDΫQ�AEr�I*�UUEU�Q\.PUh�+�s��fa�&\(�#��DL*�FBUr�ӑ(ęZ��(�YUP�1*".�rHH�E�UEF��vf�DE��.T�J�ʋ2*��"�e�aQ$��(�D�*U\�ʩ%Z!YI!*�Up�FUUE�QQr����.r���UY��(#�ER�s��A�.\㔏TQ�Q]AiAU��:�Uӥj���V�QDPr�9p��2�"�g"9�(��ATT\�J��QU9T�D��Iӕ�J"��.jQs�Ek�;��r�+ȧiEʪ͑E�r"9#��+��P���(��9U*TW"r(#��*;�A�
�U�s��T�ֳ��
 ��>�B����K�Ԇ�����`����jm�֨ȱT���\��`�md|UkT�A����!�]�mu���NL��]������ 5΄��V�ryo�v{/��>���6��7CTfW�c17�L�so�V��ݍ}�+���k��5ݭ��9����֕��A�f9��h�}�[�س��%z^��[���I��n�y��udD�ڮTn�z���w"�g��H%q�Ձ�P[��y�h�yզ]czy*[���w�*�lFϏ1��_W��*��V#[�a��Z�W�(:�w��������S�����#d�G��%*Rz�WT�լ��n�+�_��Z��d���s)��9g ��"�H^ސ
GtL4����Ib/����PR|�V���__,}�Xͯ<g��EB�oa�DĚ��q�n�����)�qm]���_u��a�ש�G��9f@FI��Ӱ5mE[�Vu��@e�q�З�.9*z1&�ka1�Pm� ���==��0 �h"��j+,�_?qiz��{���F��W>pZ^<��R�딽��$�@Um�j�u�X&��5�Vjڒ�[����Z��4��*� � �WU�ț�sv�y�)�}��\-Q�jV&h�!ʼ��<� ���r��h��=�L�	o�.�k��l�t#b����m7=�t�s��{��_L4iHM�{�LrԺP�c��q#���AN��Jܚ{�I�zyzz2G��y�M�5�hr_.0����y65�3u�xbG(��Z�鞻є��<��+�y>0q�jb���V��[akh<`�w9�xn��O��P��Q���?�}�ز���(����nҗ��5��1�eW����̓��\P��'s��-�z����u7�Q+#/�	����y��X�wX}��ё73R戥iT_5���~��
��g��(D�b1�ѧ�7�T��c=�ի�G�k���5��B��ţ�F��.z��hk[q8���1��Ԛ�Ә�^�z����q��l�>�P��k���#Q��(n�B�M35%��eu���*\n8�����Ĵ��]eP�������I�'�7� �pͻ*���1A��2�R�%�(�k�U���=�4g+��"r�l�8*�i�5ծ^)C��h[�)35��K�&m+�,*0�نƫ��闼��"֮m7�e�T�ܾ� ���.=��T��H���rX�_�> 6����hEW�UӶ��[�������m��R�t�n�{���>չLu���]��z��tU*[5�)�z�k����t��R�/f���J�)�Q���{6A@�{��r��N_u���}�0g��]^�s������jͱs�|4�Oy)�-����tڮr��{��Ȭ|D�,�(�&I�^�����!S�	W�`���R�2Ɣ���8��S����J:9��h&�t��FĪQ=H�A�:��sQ�7�:����X�DN�~�{^|��O�׹'M���6']���6b��#t/���%�wV?|8�����O�iW�N��M����f*˵'g"c?a]:�ǭ�m�"��~�yu��R���מS��u�Vⷞ�#Y�Jiw"w���d[�Zu���+#;S��o���*߻�E�[�b���x'� {�U��[r˞W�a虗�[���uO�߻M{7����Q���E���B��d֦�E3(�ޝ����j���y�����*U-1���k_!G�@Z��و��7��Dt�[KdM�#���o�b����һ��nj�u���~W���ֱ�Tp�މ��}u���2vxa�����K]�:����9���Hk��Bߧ�+�6߳؈h�~	��3/�7��Q7�tuF1#�R�U�΍���m(C�\��q���<zG��xD��ъ�~��ARX�Ո���ya���/�Z��]d�
�7l��"�w�DD��0�v�U媕�5���1��6��)�;��[�7��yo���~Q�� �@��1��u�t�\�[P֬�2�H�T�g��sYAs���7b*�{zA@��Dn�9��S�g�ˢ+���m���)��-�Z����ۥ�Ϙ��6�x�;�:Ƌt�$��6��%|��u�'��V1����~g5�Or(��Y�aH����B��cM��q���I3.u��3�;62��V}�<qA����������2��7��==���y�`1�1����n���yj��"n�o<���I%*hS4ء�7�'�1�S�L�,�iźm�=oY��=���zs���#����g­oS���*#�G�gб�}f4D�6����.�鎓���5s��!~ �]�u���Pα�F54%�N�5����;�61�F�ON�*(���Wf��Ib�6}]wr�;�ŉs�~MQ�77�i�r��t��c�:glp�S���1�}���^�T;T%�W����j�[V�C>�!�)/�_E'Wf�Z�w����~��e����:��ׅ�7�::v"�#5��r��ٿwaߜ�]:`\�v�ݥ֖�>&�f�l9���}he[�ތ��H��Gg�g}ؓ���u�'s����r�NNsX�v����gKz1	�]>n{��jw�^�EEmOM;nw�r�c��	�od��uK���X�j��n(%���l�.�L�v����u��f.�;��#dS�*A/h��������j�EUŵT�kw3U�֛}bZ{~S���%!�$����\�eX�a
Z<Z��f��7i���*���YrAޡC�++�FA��Z��	M�ymn����J�\��}@̭���z��R���L�k�`�TvCu�9���#:�XS+���<+m��x8

���Ч6\揼�u��a���v#7Z�� xt��ʷ]�LvO�ֽ�������q�P�!�%�:�T�Ͱ�����v�B75��Z���)��ֻ �3k�"۔�EB�w��hެ�pPY��Ͳ��z���(C�}�k���G�	���oC�y��y��z�q���v��ܣ!:�pq��.��=ܻ��+
Р>,_�+�W~{�w�k�?]�i����'���[����}����ӎ?t�3����I����^u���D�#� ���r�=��\E˅�3��i�Cr�q�ٲ{�Ai��ҸŞ�-ከN�C�dq����4ޭ�yڱr���c5�.�W���9��;^o*����)m�li�0"g;�#7��
�~�y^
���f�^��v����혬��uټ.�)���K^e����u�w�6��J����s�X��R��?r�ݬf
�����o^�����q�mΪrk ���}D�2;�6��ޟn5��`ܞ�r�g��Fk�{��M�Gq!�v���	Qp����+����tm��3�na����S8��_ke�;ADcn�ø��b�wntn�b���&TYV;G���+V���x V,m^ݾvr���u��2�*�Д����6�8O�P�|�\��Fl�6dk!��v����r��-��.�Dk�y+]^�/�Z��.�bM��ݕZ+}Q�W%<�����^��3�|s�}�r<R������z��(sݕ^m�d%|�}`Ky]7��g�
؍�^�c�lC���
=)=[2�t��)�-R����a��7�8�0"c��q�$Nts�r�j �~n9���Eҥ�JS�mb���8��3��:��r]
��C�(~�p��P�]K_K/��,}�7&tBk�U�S�Z�kNqAW�O�zE{Us�&�M��y%�P��kn_\>H��6q%��So(;fB0��0�ؿ���<���wK�hC��������:	��b�N(b�=H�<�F�p�t!\���ћv�lvj-$E�.�d�d�1� :�,�,��im�У��[Q�X����U�`�Jӏ8���NЬX�ᙝj]���4�蕅\��+{��j.��ÚbK��g?��ʮ�S��i�]�$8ٻ.�e� $fvoU��UUL��
䥭����Xijt�ä��rN(6�;�6'�ى��b'zCe��v�R�*X��e��{9�ث��:5i�h&��':;|�g�}��݊[���������{����y�'9��OyNl9���뼅��׹����S�=ڥQR1ƋOf#oJ���N�{\�,�De��
��u�u>��Ɠְ>��?}���ǵ"���?_5����vN�nĜkz��A��P�7mkov�f�]��֕����`��^��w݆�K����X}��ƭz�/T���l�s�g�yE�[[�oV]^�6wNa���׼�=�WS� �/��-_��kya���_>F�F��j�d�]��m�hGQǏ9�t$��m2�j�5��a��ou�u��͘%2�<I}�8Գ7<�� �@�{����%�G���"znh��lvh��uX0]hq>���1]\�{e�u{��ۥkd�j�"r��T�qզ�N_
K���'Y�6���q70�I׽Е��aq�u�[�f��u�l+�=.��� 8$��0��������ߧѼ�(�{��9��MY�����|�ͬ�ό^W���Y׭�v"�/oa@��^�:�uW���1�c��o��<��������3h<g*]*U
{���[-fn,����}��zwh��Դ�3��=Ƞ�9NY�aO�%Uh��B{�I�3m�HTFR�9�,q�����5l��~�<q^nLFhz�3%�����w8�2��ס�#��	[���oF�2��8w�f9WU=���%ogN��'@ڌ�:�ЮA[��y6;V���MQ�wk����V��vs%�v%����������U��U�Ig?D�I�^�{�wH�k"�kyt�n�>U���یОU{]���T&!&��[�P�uz�\i�{N-�iFlk�j�i�]��.['V_L�x�2��r��Ei������&�y�F'y���/���|�,r���v�oP˳f%�ʼi>v��,1�f�����͔��|��(z��"萮�}�Y }��|u!�ayM���&D7ۇ͚lv���1���˗ZU�M���3m@�K�/���u1	E�fj�l�,���u5G{U�3>���6���]
Ή ���O��v��V�J���i�͡߾��$��s���s]	��%>��'�tG>n����5d;;I=�Y�z����vUz�t�L��;[\����-k)58���F����P�+_+��ĵ���]{Z��P�ʫ�y��BmG��X\�����\|��Z������y��M=BZ{~S�J�H[��W�+{��Jx�VVl�II�"N\�������������s��T$7����lA�Xz�qL�sz�\?F^�WN����w�k�kȬ�HL*�G.ý��DV,�k6�Z�����*��]�k���G�	��<g��aby�6DսݾR��1�7��C��
�v#�-负pX�lb�ܤՌ�3���'����F��p�ěj���nsZ����[S�%��G���qH�ܞ�0��c�7o��>T�z�{c�opE��;�y���ή:���!�ف�v�:;�&��n�v	y*�m��D�[�o��})�-����� �_�.�A���.�3�s&��缣2��V����2��VV��lTQ��et�y:'T`��WcC�u�ߝ�pQ,�=�EY=B�Û�K�С��bt�<�+ƶ�(��Ԥ)���3w����)�h%QvSO)�Y��ؽ���Yʗ��KLk>| �ֈ��A3Yr9i2j�Se�o��D�l	�>�^:Kk3r���ToX��_<��N��sp�K[GMl��-�Q�
�#9�6 �[��\�Y	^�}��:�=�b��{"�sh�Ʀ�4
ݨ.��"�k`	pj�Е��MFk�4���K3�J�Y�4C���3��ڼF�
�S֋2�\"�Y1l66���4�0�]��D���W�݋ y[�&KʭT�[��Wy]��C�7G���:\��������]�J�%��J�7m;%޻L���s�CCT��;Y�-ܶz�^Ӹ:�����X��v�V�I�+�1M�U!|P�\@y��K,k�vE��W��e3A�h���R���Tƻ*>�r	T�t�Kύ�h�OѺ������:�ֈ��v����1\P�һ"��\U֫�r��gL��t��aQQ�o.���� �0�=ڙn�<,�5�L��^Z�)�[�.��E�]n�Ġ�������Ն�s���1ۗ��:��Z�8ެv�7���2>;q��ٽD���/?C<��[)����*����t������6Mĳ��)��E��q�'�zڇ*X-�Q�v���./�b��#n]����z� �d��"�t寰��veg�O�0h��:+�ӑj��Uk1m�5�-t���X�9����ڒ����wT��j�q�x졢�30��q�l�s	��E
-�5Z3{�,E����ݘ�P�]#چ��uK}y@֍�@��J�-|�5�\�f�X)�����zvo�.1�=����ѻxl��]X���i�Q�gl�U�r83S"���9��9i^��n��T����<k6�ss�I���B1a�=W4����� x�w�u�o/��f	��T��5sa%�D�t�N���*<����U}<�Ɋt�l9Yd�ͨ-�k���[,��Y���:;m;�	���.��+s��Ӻ*�['F��kW�[�jZT���R���̣c�����t�v4��p���oےu�-9�ҡǥ�Cw%��6C�c��g�׻�|���K��{h����]�1 �6�5�|P�B����q{B�pr�
As��K�i(�u��;6mn��w����b��Q���ς�t�3u����o�)�#}9d �n�<�b��h�~����6iE����\�Q�+�V�u[�Sjey3t�`������D_L�g������>�aԋ�{�\�^g;mOh��ƹ���[ZZP�b\�b Ǡ� �0 @UWg(��a˗
"� �PQyM@��0�Ah�r�TUW'(EE�9�U�#0��"�WdDAL"�A�"��2�p�%bUp�e+@�����9G8\�QEG
Kk
����UY�ʣ�E���9TQQ$�QQDEUȊ��9r���QI�

�EQ¤2+�U�"��UD+XU�QY���*�ʊ��r� �AAr�DNZ�B��!Dr"�*���Ts�Uέ	�d��**�8Q�!�6S�(����9TTTE]��Bt(
*��/�x¸Q�J�jE��v�(+�Ôr:� �GQyhr�IFBV�QATQTDQ".�S�Er�����$]9(,	B�YTG�\�p��(Q�QU�\y���US9
)QrG�#��ʹ̢�ؗK��������f�+3Y`�eV��@v��4���֣�)@����c�⶷���h�M�
'�,E����K��EsF3�M���I�������O(�Bv1��I���fc�im����P��JX�{K���u@,a�y6�yU��P�/+z+��	vt��6��ʥ�WV=���^ջ�R�kx[��W;FV�����Ҝ��f�3����!'5=��ȭG�Z�<Gg����5�>7H�{{��}�Ǽ.��{�Ũ���Z��E�E�7���d��m�:���.�&����Q��W"�f�P}�4��֌����L\���ja	q���ܧ��ݰެ�;�7d�:�)������J-<x��y\6���iEvBX�o���[����k�i2��/;ۮ!
��w�S���qPڥ*ժ�-o/��y~�כOmN#�F�\*�����dKq'��E%�]AR٠�<��[����b��F�"�L�ի�W6��3�0t-
�y^u��PǢ0B�D������
>HM˨�Ȟ�`��O��w�k��4�(�{/e�{d3074�9��1�q<!=��9�S�����s[ [/�tu�ż�⩅���n���s�D̤�{.�o^7����K�y�w��A���7�'���*�N���.��2{='�_;��ji~GI�Gy��f�x�Pr��aO{���dP�n�9wڽ��m;���j����3��yp۶��0���#b��+4B�ĵ\�1����/�>-Sލ���M�;�;p�lO�)�Gj9��C��I��;HN���]v��s�^O�׹'c�bS�8E�������Q�js�lz�g����G���YQ�����5����i�y�k;Q]z2���~�|E�mY�j�L'i�?G9w׵t;��c�����ru5���`R���9c�m�.��Y�m�ۇ�S9Z���.dn�;��C[��׎O-~;=�9�i�����?gU=io�߳�K�	�JTYye]f�RB3F�k��"�󲧛�u�����G�S��8����u�F4L��P';5�ڡ����h���3��T�|f��(�*+f�nk�C(�O�.�屺�l�/�߆�M����m�6:Q7ym���=9:�e*`Xkrp�>蕻�*Ninڏ��c	7cT���4���7�B�D��n��o��CvjvAQU�y?�=�V��]��U�	�U��1����jQj�u�]��w(C�n�u�o��Z���G�zՅ�5s�K��6�J�l�~�n)o7�M5b_>F���a���<E�拞9���;���@�ʽ%�{i�j�b5���7��ݢ�Wvl�80�}ćt^�S�^�*�S�{y���[�Ϛ���c$�Y��r�]q��i\m���ǌ=����lL%ཽ �@�����$��Wb�or����̝�j_e�ֻ��O�^}�1���5U�k��׾���{�TM�
j�j�.�-}̴�9�p�b��r��>F��圂ǖ�,\mZ��PN2MKՖ8�AoF�I�l��p���
}��j�W�׫9�����Σ`��sR�&�7y��\��	�����ONĜV�켣���>�/�(0�Ďq��)�m�ܜ\�lw-��uKg��K�W���yX����}��H�T��3q���M�Zsm���nY"��.���>$w�[휰H�$���aC�%mb�c&��(>���WE0NS�C,Tg���ZNGR�롉'������[���ΒŰﻗq�q�Z�$����.C*�f��߾���z��z\~���c]��׆'�t�-ht�]��Z�Ͱs�р��jb��ի:�ZÚ��#h�k�t5�H�]B3$�Zr*����ԄX墟x�>=��Wz��W����k�~]i'��\b���:#]�mk����7�Q+#/ݨH�|��O��<�b]]J�V�K��C���r1��8̠Uȇʦ�(D�q�O�b�y�q���Z��3N&_`ɚ9��̏{�➸�~�B�o\[C�Xsk=�i�X�aTcqَ̧���g+���x�EbJ��%��z�gYڭ��<���=���i�X]�{�C�ˇi����	���-=�)Π�ʪ؍��ʡ�8�{�w9e�V��Њ��G�����Z�0��OQ��*�����vR�Jr�m#n�!^��	��E)[(�o��٬f��zt��Y�&��F6�?��Iac9���Q��d�V�0��{	���`Jַ9�ô�J�ټiիS2�� ���$��JTX�fw�V�!sR��VAA���79�6$�*�"<��3�e����)}Y���B����4��ە}�U��[��=j���@�ob��]��r����h���㹷מO����[s�@��w��惊-��-v9r͋�}�\٨rj����̹�o�v�'���A�2�)=������̖����U���6�cW�3�Q�ݚ�M�;�n��D�#�9�؏g�m�b���M�"�甯�o���X�{@.p��:N��h؟k"�����<������8T��;��*�d��٫WM-����l�s�^�WUN�x��RޛƐP\k���e��z���٦�y؂�n�g s�������7���=�OA߹��"Ӡ#1}�%de�ڝ��~*^Bz3��4����N��٤��4=�i�Hc�<.��^�����`���6&�X7-�lR޷'V���}`&����	}S֕��n{���fe�*�Ohl��>�T/�Z�����cAn��E�v�5-�/P��������`�]���Y� sj�'�Zf�� S���,dn��oَ�2ģC��9����-M]Yaa�������vg��B�&�{8.�u#C��	�ց�o���3��PK�����v�z���ӎ�^̲���ͼ�Q/y!UF6ڤ�=QiGd%|O�缧9u�X��:Ϊ�ɉ��%.քD^L�zJ�R���+�����h6���� Eպ��7���lvP���K*�����
��)ގa��y�(�ܘy{��q%�RF��Mߢ�J����}	8�!.��K�*}'�v�iR�Ao��k��w���Uu�x./��x+�v~�Ж�}��m�
u#�vۖ���kX=ȯ6�W��daOL%Q���V�T6�J���r��ALɵ��J��m%�_���p�°����/���&1��鯗��p��U�����ן(t}G�p�61�6"�^�:}W�a�J�==��8\v�b=��{�c+���5m�jM&ㄬU��k+`[�֧�F�sR��B���[�����!Y�����������?B/�9l]Ԥq�V�fK�1T�||K�\�¼��Ny�/>�IY�����G1��k�E
α����wq����<�v�	�%F����ҡq�L .�zX���������狽Q�c���=o*�t�,�Z������]�XKô1VÛፎx��.Ɠi�9�Oj�����-�Fb�&�P�[׈�Y��X��JJ���Օ/,rcZ�����ͧH�s�� ��3������G�wJ]he[�ތ��"�����������kg��D���#n��%ceR͛�حv���{Ss����Qt�#���gF��8Y���2�Ug�eKN�4'��N3�Ո:�=�H%q���7�oe�ʴ���騅����d�cn�g�U�ggb69p�ʄ���PZ�X�o"��dt_�+9;�x��w���X����姶�9\T%��>U%'~뢕ѬP\�*���}x�Gd�Z��5�ci�-f��R���wFu�\��m�;��SO�l��L��Dg?t��f��r��Ba`�oVV{d��;䃾sO;�S��Y
R�$���w�E.��JQ%^N|��"7 ஔ�	}2�S~=�%�(�k���l�Y<�i�����ֹՉ����9���k3n��u�W��>	�U.9]�"q
u![l�,VaX�/w�_�﫟u�ebk����(Gs������ZI�׹��w�yx-�x`�s �Xz):��z�Âof�k���oFׂM+��~��%*�.��77�e��2�UizQ�Z��%k���5�Η(��̚�]�ռ
E�P��n���JY��:�_z���o�vy�9ԥt׷⽀��[��F�>Tj�ph&ƻ��9GZ3�l��OY���}��6�=S���h>�\��X-�^o*���\�=0�y�<�@#�e�>}�Z���|��m�W�n������kQ�{���64u�0}�
s��{�m ��+&3:���%�e��5�����X�u�պ�_lw}���s3�+��%�H;޴���(v�Q[�.��/�Um����x_�D3xU�i^$��m��u�y��O�!��m��|k�yk���3�Ҳ1���R��cJc��<m%��,雵�a�P�n�y`%.Й�vٚ�eB;ݺ��=�A��`��2�c��x��u
[���=p1���Ti�ɸ{\R$=�r\����ܭ�,�/5Gz�Ce<ٙ��G)���/;ʦ/9>�܏��睦�_n�=U�g[�1�8�h�5�׏.�[���~��W����o-4�姷�9�YU[�PM��93Kul��\�^RhL��HUӓ�J����k�������i���{�����3tE�^4��������`�q"9���Eҥ��w�����fמq����Y�Y�Sbn��it*�!{T�%�9�o�_O9}֎>تYI��w�z/��>Ւs+�ǘPp_p�#��q^)lP���9u���_8ܛ#�a3Zs��U�sF7)�x��y�۰��aO�JU��>)�Е��`���ӱ�O!:�dѴ�3I��p�ÿ#+�	��8��1�C��[�w�y���{ZS/)��|��8u�����A�5�p5��E��~��+�/��#ۈɋ�T2�י~�糚����_'F�0�~��}o;�<�Ƚ�pV��@�]�A��Y�U|�]Vk�Wn�ͫĺǱd��0O�Ɗ��/����RI�cճa�a�]��P��q
��$ �G�˺��>��Z��8j�S;�;{��.���h�E�>b��f&8��3y�%}��[4�毑���ۂ3:��W�������i�J^�ZÚ���u�n�^N+��n-��*��f�.�Fr��Gy��}�/g��+�p�^ѯ���vGfCI�MI�{�^
�޸��r<T&�(�q��yn)=Y������Br�0T�p���Mw5}uF��fP\��V��Pr�����x�N1Õ��:�cq@%�źO�J���3��
q�K���h�i�긞[�,�Cm�n��t6�j�g����K-4��{�s���F�T�r��Ԅq�+":A�>�΄��ڧ*ժV#[�a�^��;�������^ruu6�qp�x�#�����z��T�QN���@��W��nn�(�L=�q�徊�+��P";�{}�,����ie���Os}���	s����1x�a�2�)�{�����Ƚ������ ����e�fh�.g��&�珲���ʊ�Y�B�4j�+�h
���lcc�P$���F�=���c�	�[�=H3H]�R�
[h��1u�Gjc�tl�9qyn�F&���<�[�5���W.�5� #Cw3�;;8�í#��y:R�ގ�G��A��_
<O�E�7������ðb��������{�հ�~D��fn�LX�ھ$$+�d�Yv\�/DڰCP��KB�Z>�N���Rf-���1a�Τ�5��P��j�r�vs=��.tӚ��`r��{g�Y\�z<f]�^[���3�t��l�+^����w�^��mE�IR�CuEԼ�	���V�,H�L缺˔�F�:,�a9���)��D�X�,�1O��e�`�#ø��h�f�����$B��h��7jhz*�5�{���i��N������;�V��\�ݵmz�V���*�]���]�/ZV�tg��1^���8
�o1�Mr��iN`C6Y\�7�E�ӆ�ռnPg�LP&�ȓ��n򰳝}o��Dg_kK�o���|��!X�F��ZJ�CZHu�����y;^&|Dx_P�D[�nH�f{���S��nA�Y��3i헽���-F�V��������yf��b/����._�Ɵ*�]ư
�f��c�[c�9mF����c�M�)�0W3KkqXWJ��xQ��4敊`Y�/�*�εM*/���*B��\����p�o���FVG{#�l!J��}:��VW���)V*{|��fy�w$Jx0Щ�3l;p_}�]�^��5�52��hp��D2Zm�ownW�wm{s���j[>w����\9�zv����X�!h"����8Ӟ��\v���6r��o��9K{�c���l5i��m�%���3q��޽�j�H�C��)t	�^�:�T*
a��z�Ŋ�.��n���Rz���^���wK	�����������m���j��e ﮶�,3&�')��/6���	9��咆�B3+�N:�us��Ɗ"�*ueI��ڮ���W𖷖YPn����s.�^q��+t��`�z��L\�í#�}R��Ӑ��L��	�M[i�b�oh�t�Թ.=*�T�IWk�Zkܬ�w4�[3=�$sQ�����|j�wnv������#M���c<�BjnlT����&�G��χ�17�K(^��pJ�3�j&��_��1��W��$�~$J��>�ȡ������};{��r�����x�]�8f������;]�1� �d��(�><�ԇj=����B��L��v3}�]���I�}ځo;�J�Se��(ݍ�>"+��p;�M
<�Y�/^Њާ�ݱ�=�ź.�aS8�����d��tO}�����o����w5��%�΄y׿A�|/�^r���i���7P;'��Q���Va}W2�9��0�e���	�����r�]�,v�WU���J2(���U3��(�JV��@��i%�ć"���5 9@TDF�s�W ���jFt���H9UQ�r��!r�dr�q�DQ�:ep�5!�\"M��)�H���9�+�TsZd�ar
�5+��L(9S9qP�98ܴ���TG"9s��WU�.Qs�A�DVBQ�H��,Ҋ�Dr�EVa"(���r�h����RBr�V҂�#���Q+9E�*�J����d�E�\��QZ�J-N�Qʢ$�g9QԊ(�EQ2����T�*��s�(����Eˉ�˔DEEPN�\L .�N�(p�N! 9��r\�QAA�*��"��p"/'��".ʪ�"Q.�$TW=09��QUU�"~����t����Eo-��9�?,vǌ�f����}r�Z����V�n� y�P�sg%]�g�R����r�z����}^��*�ٶ�rC3�no���Qi/3��{�A�q�qS�	S��f�<�3y��->i
�v���漿qJ�ލ����7��G��J���C�� ��<��y�fD^L�����=ɧ���{�p�ޥ��o
(7�IǓ���p1N�N8��!\��̰2����[^\񦤕B���4v���e&��^������k��g]�s��E�Ќ��/3%o��9�r��>��}zs��eƽ^�����)��Oj��f��h�}B3M�5C����������#v7qs��ʗ�ɍi���>�6��n�8̠_�;���fQb���xbk��t���e��>�|�<�c�}m��ޡ�g'y��C�׾�-q��ya����BW:2���/�v·���Ǘ�k6�\mf&�nvr��Ż*�8�sU	sմ�V1{���f��J`���(�X��Y%����z;�{>ɘ�M]�D��c����bj�u�z)�s}K7'QF��O������=׮fgL�ƫk��'�ĩ���	�6@��ϱuz7t�uˢ լ��e�5�x���ò�ƹj\�G�g�h�ː����_N��V{�?v)�x����a��@�U'5�
yѓ�[1��u��?c�z����.*��%�II�L8)܄C��Ml�D�i�lemJ���kq���m�����!��
r�P11êڽ�7K��Ws�J�r�{�_e�Z�f��O��!0�ּ��M���|� $�g�o`%գ��_u�iXg5�'���](�e��3O1މk�+��#��Dl�d�w��U��I��Cu��u,�9����糪+r�l�g��R��sBV�����4�R5�C!�Ы۔4aa~����P�J'�h��F�-������1��]{}"�ȝ���E篻jOI����h������t�E��!ۈj���E)���n�����m6��^����pZÛlFho*���r��>�U�.���Ѷ�u��B��a`���@rU)P��6���+�#:�}JP�e9���7�VU.ؖ:[�U���5����x��/�!C"�4�v��)�1}J3Cr���_"h���N:�.�K��츘�w�����Qhz�<w[�2�����Q�N7�	y�:����N�i�J^�cc���*D*�����C��).�ܪ��3(�ј��oj%de��X��*^E�X�s�~�6j�<V��kډgZZ8ק,8��p��Ⱥ_����-z��!�ۑ��1���8}�)�筘8�7=���jڗ��_S�8a�tJ��MLp���qMs{�v�/�7���;��#d�zR!<��谾;�ڣ<���p㠽�چ����i��Ol)Υ�T�F��*f`.h�u�[u�y����@Ių'�uuMM��e�h6��m��*R!N���w�2%����;�4�z�+gB��5�k��Rlƞ7Y��9��6��K�EB���%	lPϮ��������i/<l����3��;��[�lP�r��
Gy)���Z��0��B��9Գ����k���vl��3�����8/u�w*�b捖��d�63ӬY�V����ӧк�7f>���1���͋�"Չ����TIv`��R�شx��q���핿*������8G;��K'W<����y�nL�域�z�C܊m�l���!��>�]P�j�a�=;�9���/��-P{Ѵ�hy7���j()Q��֮:g��¬l�i�$)X7��$����.魛�{K�:O��I����~F��]���麍����N��:͏U��~9BD�{�"|���>��a�y6���e�����E:��B�������2�=���y)���{E�v����Y�5���S�ܬ]U[��j�'�O}�m�d�?�E��7��)��&�z�%N�n��K�g#���8�ŎoZƨ���ٺ�2�V,��ة���^^���%�3�c�`����}`&���d[���q�^*��gkP7��gj�sQ��Ъ�9(���#�K��t�ٚުγ�%���Ɲ��mV�kyFA���u%u{i�������u��{b��r4����Þ���X/��5w�Qaw��S���h���zײn2
�@����/�v���=�$w���{��huuʳ8qf֝���O�9R���W�U��̜���8�5�p�NǆF6�A��+p�I�ziO�X��ھ;��X�[�5ѳӅnP�wԦ�o���>h��"���z�b69従�[T�_��V#[�a�=���F���۬�3�Z���~��ڜ�b*����(�IK�u�u�Kg4,�ogu��O����^�=8���T)^ޒ�qP�R;TgSЎ�E�B/q���9}�jb��r��TB���2�5���s�sL���ALÄ�؆�ovpRҶsZ�{�M����;���%��&���چF��A֦�/^_�oF�\�o���������ҹ�F<;}7=3�:v��N6�sr�'{�|��O��$�ù�]�����k�7���[����i,�XW.�����v�*�y�W�^�Z�t.�\_s�lk��λ1�7_mz2���)k�Q�m� �0k%b�؋cu�1z�jՆ�m�kh<�;a=ݞ ���>�����پ�o�V刜���aO�Q��9����=�k�^q8OC֒���B�͝��<j��8����*�Ŭ��7�N�����3�I慫Tx�??�|��Vu���kR�ɵf��k0�k��njBf�����������m$0�\�sSB���R��y�8�~�~|c���0�Vp�4a��Nz�>��}W#�8��'Z5Vj��T�q������{�|������eX�1�U潻�j�8>�0�B_/����ҠFJ{�"�{U�UO#����E-��݅F��Mϒ^��x{2P�����JV���g�;�}T���Q磪��q��C�dq��x����u~R�J�V�5¬���T���$験��A��We��*��{_edme-��j-��x}�C/=�;��}�1�U��x%R�������u�lzMnWF�׷����춣��N�����M
��XC�,�8�g���9�e��Q�P@��E�W�^�M׺��}�Ь.||���2��
r�G����r0��Q>ߩݣf�O��2���۬����(�� n��@S ��E�ϧވ�(u��|8z5h3�3�:�'f���!��{���q>/յ��>�"T'I��u�d-/�a�����{�Z�1��``���[�ϋ?�|	��<m�9pK���~{ѮaT���-�u���=����X��ݢ���66j%NH��+�̼u�>��Sl흗�:8͐޸Q�4v�� ھ���r�'A�FSu���<�ͬ�!ɦ���z�����V�~V��w{��i�)�����X���&�S.g���H�J�to�+NU�n�s6�mF�]:�5O��z��>�]���p��ɴ�p/�0?B5�+�t���Q:*�f�υJ��Mu��:-���;���yo 늢�6^�w0��]ɸ�Kdɴ�������9ʼy3k�}���^аXqe۰ֽ�\1�T��km��m-+���wzcе�:7�,����ixg��T����߬��~�}.�\�u+��ZN�3i{n��%O}�1:�g����0�������w��oIx8?{�8m�'v����D��`ӭ��[ U��c�*��&>� �8z�/�N����X��ٶؐK��ܹ~ �C+��I�ȯUaPس���wraDޭ���'y�z�rr�F>�&�Gz��ܞ량Q�2���}T��N|QMu�4Eww��^��\�tɸJy���	�����{�.8ޝ�Iډ�(7T�\Բ�W���}�[���ɋ�Z�.mk��5��yE��М�{�M\=F}�Q�Ej&��fM�o\͟�j�XCUA��(����B�J�(��2�+	ѿ�����ez�1XWIv�l��{
�5�h�{���(]^a-m����<��f�X
����"�W>�{ V���')�b@�"��{�W���,.�S��̟`\	��{6nMG���w@d�,z�Wۺ�7��b�:ck�Hg��g[U0���w�3�.�y���C�1n��L�%�`@�$R����K�V����
�����G�+�(=f�w�^����B|w�T'�_" oQ�P$�ZM��+1}�F��z���w�����s�t�󰏧��놓oH�uHM)����)�䂔�>�V�맻~hk�05�-��!�ӛ�cͧiO��Q{Xn�ß3(�P�);$R�_Mw��^�7=^o���S�����#<ͭ�Q��[�p��%�>d�&��6�EN��wuz`;]Y�s�^�Όq�c���h��Z��^�;�i��Έv�]Ʉ��'��_��B{���nF�.]!ݪ'�3�w�#$���v��;`�0_z�6>�T��l�����Drwr/厃�+ݞ.�쮞�>������X�]� �l�z��[0�o��0�u���>޶4\{o��Fy�C���*=��Oe{��N�5*�8��3n�+��c�Jy_#~5/I�k���q���\�M�M��f��uB�J��dK+65µdQ[G�/�z7@\wC=��ʏTv�����a	m�9I�:���0\�,���m�3q�����A� ���1z"}���pr�F����9u.� �[s,�T�s����`\��c�Jۓ���y]\Ҫ��X�Ҿj�'^�h���F���ȗ���`���yl �M[=�=��+�A��%����}p����e���q��j��^�^/�8/��r!��(���'�C�������[5R���.�9(���6�s,}�L��u��a���=����^�tN��Yd������T��q��"�6hu�����NS;=Hwz�R�;�4���{uU���5���wz���:Iڃ0��3ԅ��qکb�����^�kw�g��{��ޒ��U~�f�p�ǟ�Pm�A��ʲ�/��#����?A}P�(�G��Y1�яk�r�p���g�e�_��n���R�i�jw���<ꑗݰ��� oNI@L��P�5����{<|�=�_��<G_eX�>�o�*�Ӿ���8��;<w#-�#5
dk��<j����j|;U�OnowC޹@�4��}��[��:;H�>�h�sĤ�'��T̎��̃a���g�۳��)�5$�d)!�o���Ju��X]�޲6��a �Qe>d��n>�>�
z�9y�A��l��Z�>��g.�QV��˜�w./)&�T7��2�p�7mGڱ��.�*{c��ǒ�rU�͖<Һ�Pۢ�8��.���7�f�~�`�<y�刟-�3�%����y�w�&��
:�Cz���:+������MFRv��'lǥm:7��5���VC	�܅��刱@�O_<�˿gq�=%?��9
���<v2��~[[Y魄�w�58k�L0Wt���R��=��)���k��;*K�'@9�큥�ddF�T�_t�v���6r|:��Y��Fk]k�c��9����;��K�~����$����Z�E�K���_q~�����A���,�Lk�E��2f�tS���\1T�'��)��m���J�xcܜV����q;���)�lX��X��D�G�S��{ݬ4fx���}G �,�g��H
�}�`��l��7V7cn�T�;4������{�?}�z�g�9�az��(]zk�T�@�@Wb�\Oj�����j�{�Vv�ҝ:����mpι�;Y=��^5gjӪ�qj�K��)ëf�1�7�B5���{3V��D?�KNw"� ע��c���l.�H۹�N�9�A��WF_��q1{S��ž�0�+�veu-���.7v�k���C+�U�et��V_�l�P�A'j&PCΛ�^�r|�u3���f�&�i�\n]��M�!t�]� �/O�&hW:	��#��sKKX@���y���ŝ��yA���A��2:�l["��n�|��a�EOH�(�3AS���k�<�V%ه��ˣ�゗G�<��ۦɽ�S�U�z�"�V���(���M��v�[�w�r_leݑ��j��K,�@���n����g+`�S�m��T�r�&��G6�g'o^TQ��׷����j�-�S�5�e�uf&�F�:�-%�.COH�,fl|��w4N��ao��K�S�w�ΎS��7z$������ w;Kg�ԳnZZ�|���L,�2��J����h�.l���;�J~ʑ3���n*,Ζvd��x��vٷ$)��]׾Ϫ��3�u�.&̝���E�yfU�w VWT"N`�2��n���8��])g����zO-�zu���AF̊�ǽ6�Y�&"�}��c�Z2ROf�����eѮ��A���؄�I�9�}�E�$˝��
w�swO^�QA��Z���]�>3��+���mU`"�%�䱣M	��}��_ �n�i��o6�ǫ�h�xY�΃'fS����,�0��X�A����5^۳�$(�b���ե����Յ,-����K���P�t�)��nz����3.�Cw�{���Z��������93_D�GUa5�Q�$�1�4wO�o4`U�(��:�����{��t�*�v�teE�9t�x.�=w �&�V�EՇ)�G�z�)�/3)N�Q���И79iw$,�+�˰R���7�I$r�
���wCk4����L�ky�8�L8 X	̓������qn��/Pd�;ʅc����\����`i��H�Zzڜ_c������"�ӿvn��M+`�H�kt��Zyۓ9L��>�����P��ݥ��(c4Q�5}�Є?L�'	~�^��lQ�����9"���/w]3�Z�g��X1�u�;sy�G@�x�H��~#�r�#�s�f��qB�G�؀�]�ӦB1\.�;�?{夦2���W�J;v���j��S��>H�{6�a}t�܁,�Je��.����mh��u���\t��%M
dΒS��|ܒ���d*1jy:	�>��J�C�ט��O-6�٢N/�kXc�Dq�3N,v��(U�W��F��R��0k�ȴL�r�:�g.k;_Fr��mq��>�ybbͷ�j�AgM-
�j��� ͔o=�ul��{��8����6�c���hc}��:r7\ˡ����j�٧�*˖��`sx��y��(<={<3|TRLN�rL�B�
S�94َ�TC{�5g&- �'ϖX�l&���{�9EzI�ќvrl���Hf����ovi�w�q�-���,��ۓ�7^w0'N��R	�{l��vqⲇ���ע�LeTB�%E&�&�Y�{.X���������.�)�%G(�#�EQUr��ra��*�#�A �.QE;���X
n�+�r�dEG�J��C�t�;<�D�P���U\���W.YҦW+��ȫ�]��((5�uqwL�9JU���UEPa���*��e�놑�	�BI9XS�\uR�NQL�P�L�e�3��d^��J:���;�F�AAA�+�\eDs0����E(��DA"Tz��:���n�x��1	�q�T(���)����"���Vs\Wq7D�d�&-$�eU.G\�r(�!ʎWq�L�0���VeDE���qfNT%�NRsI�eȪ���8��6��]��j�b��I���V��^��k��v������� Q&�����:�!wƂ���m8����xb��촖v=����?�Ɩj�z�_��O8*�+z}�����v��\-f|ˁ@�.7��e��u�{�=��{��0&_�|�,����t�t�9u����]�9��u㨟;�Tf���i���g�>����:j:� �bKd���}>�C������C�sm��mw��p)W
;��,�������N#%� %Bt���[F�/<:�+�ox��h)cP
�0m���Gy�8�=H��p2nu�_���Q.g��H�[N���*�Y��r�@������7D�.�RZn���1����5(�fS#M�z��u�xo�������.�;Gϥ鿗<�~M]ɿ)L�6��5�����/�x�w�=��w�K�@�3������z<�[>
��xpev�ٴ���������酮%�^r��n�˶1a���s�\�g�k����#>-N�������*^Jt���A߶���%O}�����W*:pu��%b��G�ar�{�&��>'2|Uw�Y����B��o���x����͚���rl�o�c�/�vd���vuC�H���W%.~�i�{e��ge��z�!�:q������V�Q�C�ڃ�8�Jt�fċ�A xr;3�▫����`2��K�]L��y�r�d���.	�jU��q�J��i�#Jz��w:tFX�?܂��=�j�;�Y*2�f/�'1��u�Zoƥ�JU�6�f�Q�`�����4 q{��<���.c�g�Nme��7'h�t{��^5v���BPq5�eּ��	z׺<�۞����
�c�M�<��u	�T��w���_ѝ>����I;o!�7|R��cH.an��������(9'�Fۡ.V����`��,�>�9L��P��q~�)�ā��W��sW�2�tC��~k�	�5ǟ&}ݱ��k�Hg��g`�=��Vn��	w�}^��Y�;�䲆�x�GAr�O��]D�V����N�t��ޚ�޳x��~�ci�7�0���>:ݻ��r~4��FC����Y��h��`�g��{~�wk�h�qO��s�9�|w!:��<u#/�T���d�� �2E�U���ԍ����گ1t�{;�������	�jN�>s9�������ۼ�fr>S$�Q�)����U��k�D8�^�*�sN�y��*6�.�%2��T>d�B5�)M�E�W�J��jq�<�Κ�r䙹�Nw\D��(�>q�g�4m]�l�ڗ�g>�XU���	m��w��s�,�j���}EVWw+� ˶i틲�2��c+��t��7	���ih܍Ҟ��U��z�pu)`�\���C�6/�z�o��_�)Vl���o�Ļu�k�Դ�˝��0�td�TC[B��z�=]O7�q�����8;��X/�-m�fۯ���q���C�}��ȫ�-Mo�RT���ʼ���0�{
q��.5�H5,���[0�K�x��r����cC���N'���Y��ǝ'q�[3�_�]j����q�*��̋��Q;^����wh;�e|��3�֜nI�w�w;���'K햍�o��J�xO��1�NCWQ;=�h����}q��×2�I�Ĳ�����D�gwE)73�IH�#�@q�����3��|�[<�����,%��+|4��x����n2�'={�`����tw����piP}#
�ʘ-*�X>��&{�K�7`';�W�w�SK�g�\��<�R��d�Y�=_:P��e�Adv������_�U!�~�I9�ܪ��*\��Fs��y��f�g�=@�^2�Ŋ�H�]��Mۺ���y߽�Y��6���fj�n���� ��n�z}
��/}�P�U d1��
2�F���ӷϡ��4�%kq��0�R.��Yi��Ӡ���/��r�5���fKP�\k�O����Z��f��CήP2�!�`��cn�5/kѷe'&a��Yyz�[��N8�Wn��F�t�Vr�/�)��e؅�~�q��z�.�%s�ܝ��N'�ՙQN;xy���� ��Ω�S��@�_I@%ٻ{A�}b���՝.��Zɠ��+}qW��q�S����9v��9�f��(�V{zL�/
�|�����/���A���{�q��\5K��/���D3�'a�q9�S�%W�j.��^^��Z\d?L�=$�q�FĞ]4."��9���oY�S"�Ygz���'u��I�gc[/Q8��zG[�����;p&c���[N���v�{��w��d0��8{ut1U~��5q�!Ʈ�J�,~�n<'�k����;��D�����v�X�\��x�Ȣ3Ƚ\C����W��>N@sН�4�|�Ш�~������9������5�j���qRB'9U��Y]�jx�������7�\/$���k����������3��6X<]���cч�v�o���N=�ƅ�	�z�ˈ매��f�f��m���J�xcܜV����q;�^i�`A �m�_��(gn=�L�}>s(:8����]L��m /\1����.���&���k�
��rc��z������t,�\�oM�_�59��|����-.	=s4鹅\���n�P��x�"���(��m�g�x'�]�:�퐝�C�ڂ1��P\�.Y�s�g��o7�z�c2���+��]�m��Q;2��x3��7u�Y�{�/���¿4�<<deyh�����4�ђ�؎�|�,�7�����u���=�p��=�\7Ky*���b�ĥ~23����n�%E^�Χ��B�Ȝ�[]����=�nv���S�r�W�23�t���%|hTߺc�
�3Q�Ֆ��v}G`N�Uƺx}�C/=��>�}MS�e�^�%R��>c�5&g�U������z��X{�
�������R��4+!r��Ϥ���1�gnu��D9�eơ���[���W�<�������qњ�>�ۮ����k��#\�;�������\����`O���>��^�F7�.J5�@ޣ )�R�"��}>�P�Z�:j�;���GW��뫷��ߞ7��M�<w�˘�FJ* C`�#���u����*���X�qq�N�%߷���8?�'hyˮ%� 9�ɶ�`��&�L�������;$L��DMۊ�]^�s��^5����S޸h�Bc7�]nM�n�����J����f��=@�쫺wo)q����o����z��&�&�{��J���sn�~�6Ϟ��[�^��)gB9���J�2�*K�bK��Yz8��C���L3�H{a�}d��a*�xHۄ��
�u�c��|N�=ȍpkh���\�Z
,`X�/w�]�ك�ﷻ�^����*���Gh��^�\���5w'ȦL�����#T=��d»���R{g�z��^���dx���s஧�࿲����Zmu��ruXc�k�tn<��;�iE�=)x�9{״z�u����pߙD�����wS���
�q=�z�w��c�%O}E��-Z�uU�����t��V-�
ީ�̳1�a�7/��Xz;m )Z�
±Xᵕ>�jN��rv���p��n�.��{�SaK'v̇��ʃ�YU�(@E���^w������}ܽ���ր+���E�:���:�}>MV��Y|/������O��^3��)g�/e���&�9�U8��Xm\���ˀ��u)�^�?\&W��\n��C�nN.i-f��y��f��N&X�'��WLnڡ*mk��]0nQe�L�uSWr�p��j׬�ܵ�Zn������� ˈ���OO����}}V*��cG�ä32��J6�1�we�zq/[y����ϙ���P��z�2��{���z�bZ�k�(zg���7�e�U�z�6�T:u��yxpً�c#y����ԛH�[9�����)�vo:�]}�_�_f�` E��.���i���~�ហt�V��y�N��xg��e.�H5�9N 0�����g5�F.%�k�p�5<5^˥C��ү(��,�\�K���ӧ���2߃�{I�#�:W	��:���,�B"�0�\�I�'���z���c񫁯cN���ٻQO�t��<�)�܄놓<u#.RJd��� Jk��c��]U7[:�����}���
e���>+xL{a'iD9������m� ͳ9
d�ZyUjw*�R���ntb�vH��!R^�h<�f����r\Br��|\���׀�z�SS�=��V=��%ć�9=7�q�c�.u��]���wR�k���1�$��+ΰ�����0�7.����m�O�40W���I��'�FH}q?a�-m�g��=5�i]Ua��fV�ǻY��dv��Sp��'n#��X�yR��C|a�}[���_���H�:w���x���Gb]!�h~����UOO���ǝX8o�U����G�'���Aݠ���_��F��=��ϫ���'��f���ǥU<'ܩ�jr!������,��3?Xa���^��ְ�Vj~t�:��O���Xl��'��J�����q�%+��zW�j���v�'��U歭^���+�Bp��ienMh�w�a�uܡp�.��lE�@Z�R��#�S�s���^ᣲj�H�����OLTFZ| ����q�j��;�^����w���2$DR:����Y����M(��=B�e�K��a�Ԫhx��8{Gs�N��7�~��5����f���]��㒀끊�7�s,��O��)�8B�^���Գ5�ߟ_2/VT�,�R���A�./�3�=Na��6hu���K�K���^,�-��:l���p}�SY�-w�Q�:�A�L��s��.�*�G�?,��V��k��mɦ��|�F��;]��c�l�9�Cv�Ӂ�҆(�w��%AE��s�8�Vx@����o-t�u�޻��p���Z�o��!��F:鷝R1��@6J���7�W�к�&�]�l��[u���v�@���.㲬>>���;�Ӿ���8��:�ԏl9�g������T+�^�;׺��Qwiʙ �����G�fΌ�u�ae.,��3��r7��^�`�������b�[�e���L�!�c�fb�N�c��Kz�m��Ë�RM��~U�����W������v��,��Ĭ����@#.OX������(	}_Q��k��*q�D���u�,��Nc���F�ͪ��9*d�|�1��n<B~���D��A~�+g<T?����;��9BiE}�=��f�=�����U�n�fu��`��T�3>̂������C���x1�W��feZ�/ΰZ�<|�7Y*U�s��ba6��Ua܋��J�ںN�=]�o(oYHK�ەEf����]Yn!��-�8�$�����\�>�.�z��m}���&���G���'l/�#4+_�A���¾���ea}�h�;��;�Kxex���i|s��zo�~�^��ޕ�@tT<�b���\G�;�e�oxW�׎v�����h,�xda���W��ꕤ��͔��o��M<1�8�ec븝��3g������/L����� X�?Z99�.?;jr�ŃJ�����(^��*y�}��\Uuz}�s��kn���4��~����Wȋ�S�����2�.2+�Xo�J�}�R�/)�W�{].5�^Kh�u��|���*�[�P�Օ<o�~%+C�^3��2�H�lI�r�^���O������cT4tctG-�nw>�H5�|�B���R6���N��<̷�<u���9���Lﻺ*�[����r�K6�]���]<8�e�c�O��MS�Y|��X�Aٞ�Eס���S>��۝��$�6��B���[�=޺�n��W��>}%���c�μꅖU�韶�=޿\���v��m����p@��<@=�E�L�ۮp���Z�q��;(�9
�j�i��m�����@#y�ذ�m�{�`�K=hsNy*�<C�̓�y��׎Qه�9b�_s?�.Rs�1ne�M�e�Ԓ6B}�r�ۮ�df�(�Nﻶbҍtt$d.�&�|�Ȧ���̫�yJgV���/�o]�F��{%։;k�������/ռO�1D��Dj@�G���J�N`˅~z�s=]"ьM�e�˕��g���V��u�M�w��Ө��d��@K�11��qV��C�j$]�x眉[�юsx�_���0\4ՠ˞%�>��n���q4�\�@!#�d����Pgf�U�r�y��s<�=N�Ⱦ>�n7���]NO|��Ö �Bl��;�g��2��\RG�h���<g.S��!�l�T�q�gh�;�i�\���WrVɣɺ_��=�`}�,W��U�藾Ž��L��8������9�W�Oa�e��+ٴ������'w�=����w�om������a����O���@>qw�m��>7�����e`R^�U��ͤ����-Ll_�zh?n��-������+#]X=oo�^�O��D�Y��P'0¸�S�piV�P�#�NC�v�vOwPH �uZK�����C0�B���Le�d�ِ��?*KL��d��~Y�+�f�x�������u�/�u����B��(Z�$����Q� �*;n�[��i�ʗ;I2����E�>��!�mH��BShK�Y���{�� �uvã��y��nfF�<�xvƺ��[䔥x�R�e<kM��P����ƚsz����Yf{�*`ݺ3���)��c�޶���gkf]Ǻ\ĸQ�3`&<�N|�a�l�(Q���İ(u�7X�mVk�e�#�1զa@bLS<��uq>�w���l���v��W��JAtD��.�u�p�Ϣ蝽w�2�آ�щ?uC�����VE�um �1�L7��YY�(L��qxuy&_��J�����
��r
�V2ܖ���)����]�pu�2�_>|�ry`�ä�b�N�[��XI;u�W�]ևp3����%.�u�ի�t��
��ցn��xv��5����Bgct8�8�����IH�]M\bL����C�Mk	n�y@:�V�`��W�ǵ���.^$�����]F%8�w�ar�����f�$Mi����ӵ���]���v�\Άv��H�[���j�T׃O_f�{�,Y��8�pbk�s�-��S|;����==����i���JW������֨���w6n&T9��&�sU�u�ަ-���;o���U�'����N��ٔ���\V"��;\.,&��TE%��5 ��YXYؠ+oi�x��O5�	c3��͆h�NĦ�[$��ʽ���x3�s0B��դ/��ݘ�b�{�%��r�aG$7[�	ɰ�r(l�?u����1V�=�кͺ�Rƪ�2��gJ��{+R���̣K��7|��������{�`}��b�6�x�N,�)�
p���	�PU�efV���f%ͮ�O�o���}����\��`��~(:s�7��⠡�Po�6�vb���v���oCY�j�a�����O�tP[I�s�u���N��#�`/eg5{�[A�u�]m��X .p���#�X�q�w�a�ח7�~�n慎��O>�ۊjAg�`�*�X��Ёȕle�{��dh��5	��]�8�׆o���Ņ�e$�hv�� ��2�Pv�p��t�wf�%z��D�Ԭ��i%���><����g�[3&�������J	��i�u���m�ҏ{����
+����[W(<녙�xn��J
�F�ơt��bl�*9ji�J���G�|�N������
]�Ş�F�Q氈Dם��,Zv�v1n�enlC�N�9�f ��n�Z��Aj�w�v��t1�&��T�j�G��󨳠r�ʧI�,�dԡA�����nǗ9��}g��u���o���x
�r��C�x��������#��=���,2ö�78/Z+4��%T?]�;�^�����e8���C$�9�����6��.�"��m��kvaQ�7�>y�%��V/O`#s�`����m�6�|*T��e�jxٷ,V˷���s���9x��T�s�2e��/9pT�DHZ*�.ʴJ�g(�\N"�)�uD�.�]3"��s�B�+RI5#V�ˑ:��L��뮹�E�����ۧ�J-�+�y@��Fa�)D㭗(�B*�E$⠜.�r�NEU\(����Q�;M�ҹETT���q��� �eM�F%�s�@B�"*Ht����S+�D�МIĬ (El*�H��/&�2<��MX����qC�*��"r)�I*&�Z��0�,+h	�E$D�(S$X�;+K��ˡ��gH�t�gnrk"e��y"����pW�꓉�(����z��
�4�)Qt��8�`DD8넦RM)7WN
�B.P���(�"y�	�.Ď؎S��9�N�y�n���/w8;�M�+P�I�k�U����z;��͉�&��,�o(��UvwJ��g�2�e����}r�h�>;.�r�H�+�r<����!d�~j���[�oW@}'��I'jg��t?}2�b��	Sp�Յᮘ6�/���0��(<'J��\3u��WN+�:k��e��� �@H/���s�6F�ʮ��r����h��V*��b�h�����-B��p��;pڸz���|.J(i'�@h=Ċ.R��z�%���u�k>ȇ����{��x��_
Վ�'�����u����w���B"�}a@	N��Y�C�މ��y绡������n�{���>;�	�%�؇T�ҙ*k�)����5���N��e�)f��C��0l���P��-�Q������il����6� �>faN{V�q�9Y��^��������e���EJӃ=���mo
��K�ɴ��,��.|�~��[~[q��wx�8��$<��T)W�A�ê^[��*���_r��s���]ɂ��'p�N�׾��~�~��d�[.����ivd�GNǌ-��b�We��e�zkٴ��mDȡk��J����ӂQ*�.�u]���Vx<��^�����GLL"��m
(�7����}i��2�5(q:1з{�F�C��P'
�\�uMI�2�&���V�Q�9�I�T�>��t,�t�Q�q���1;�狌Rq+_�۱[U��#V+���u6��'n9��ו �d�|=0��Na��u�i*�G�昰z�fM��������N��cE�o�ǒ�z}]j�ά7��\o�R=q���Et1Ҽ�*�{S�v���3y��(�ɹ�,Լ'�;e3~��cҪ��X�Ң���{��/O���u�����EI�[�>+7��[��2u���As���^��pKd�*y���T�2�����=�5q�ӟ�ie{�i������oYy��}�ܜ9s,z�::�*]��胒���b��\��	�Y��/����w�ϫ��:u�5q��Q��ӱe��peP3�	%�͵A�C���=>c�D��H�����`��u!���3ާ\yMg�]�nΒv��f��R3�A�D�y½������:|���+?}��X���F8��{ ��A�S���\�k�t��a@{��m�;_:����
φ|(��Y�b~6���\*V��9�jw�c����T����a�>�Y~��dMR�=o��X޼�]�S.O��9�|
G�&���E?�;�>���)����r3C��>�����bsa4=�r�Oc/�v:@�t�ޛ����vR�˘ᝳ"��F:�Ϸ�]\<7 ���Dy�>�|x�����fW!��~���LUt��h-���g$_�y7�{+�_+�u���ë�K-��PZܧ&��g�����f�����d5�C*�@0ҭ�L��q\{�\7ʝ�c��6�>s���C[��T��г�{_s'�]bv����P�J5�$%p6��<�h_ԧY�GaZ޲5j>jWE�wc7C^����s����eD>d�D3Q��TMDq�'A!}�=�T����\��_v����1���uoq���!��G.�Ja�}�~���D���Mi��}&���ןG��N�H�8͸zn<�=	��7������K�3B�����N�sz��b�Q��)�އ�쳳�"�f˞Ҹ�F��>ں����ֺѷ�LV�!=���+*V��r|=b}������z�)�8�,5��X����Le���t�3e3{o�F_�lrqZ�rج�Dj)w�R�nyu�8�8����a��x����z5l�������^>�1��\f'��=~��V֩��4wX�{������1��T������������J�}U�{�8�'\���"�-�.{U�}
��R���>��E�jʞ7g�R�d<0zC	lY� ���#^O��E��@\�@��+��6�S67��"ө����7��q87��[������*�ׅ�q��N�C�v�25pO;A���0�K��x�ތ5+L������6��>z�����zi�N�q�m�h��Q����{u|Ѵ����-u싗V�n��{lj��(�tC�����A�S�w�e��hl�����0�/x)�S�F�=�e�f����Q�f�\���T�s����2�����ST���Y|��m�a�'�[��	�s���&PuC�����Gz�Q����W��>��YZ}�9�?>/�r��y76��yW��y��#ހlT 7��~<@=�E�L��v�_����^S���D�n�n�}�:�����X�N}����z.K41��|!��	_)�F\#����t�cVn�v�v4=�v���������N.bP%�"U�&&y��������ȣC1V��Y��V8Q�o{�`��j��\K���M�۬ߝ���e���2<]Nkp�]���w;��owE2J�:23O�r��K���]NO|���:`~F�+��VM\U��0�ů}y�?!�fW͏D��
���gh�;�i\�P�5w%aL�<��5�=��캫qմ�x��l�L�0�MJaσ��Â����+.�\/G'w��o�k�Z��)W�a�doA�T�$�5fD�us�)���jZ��!�~�[5�j�ht�q\��{K)U��>Z.�x�3탷��B���Qxos�Zt�H���j�����]
v,(���J�"u��� ��p������wc�	ί����ϐ���nv%_�qP4�,�~3g#K'�zau�+������wٴ����#��깸�7=��N�ϩo�щ��+5Ճ���X��%��� ����xدտ�����evr*�[����=_��| ��[����8�e55���ҋ�ʘ�R�ݰd<'��p*b�:}=?b�&�RB���,ԶOxe0Gb�"�sre�y��j�w���gO��+�7�^/s����f��J���;Q��x�ܨ�_�2o�Jy���p�R��3m�^�����[���ǁ��>����v�g��3�\T�鋍�BT�-uaF�`��,�5~�ޯmD�#t��u>��wnt��;|��3���eMDex�>�|&���_U�+ك7��>�G�7��?u!��A�����B��a��F�$�@O��*��r��]1�[�OU�}���w@��{�/�M�y-Z�a�y\'t�Q,�D�3
X��Q����{ilL�/�?Y?x�e�3A�`-}qV���#�|s��M��R2��!� {8��gs]�L~��^�.`��v���}d�y�W�+��Fl�z�k�u�w�h@H�B
�N��w�������������tv���\ƭ�<&<`�}fHmn��������(�5@�8@��9|A��-�BE�:VD|�e ��Dv�M�pR�K���}���\{���wl����:ª���zT.+xL{Rv�d�Ke|^�m��+<�(����g��c�R���Yz��3d���O3pvH-�
���{~�<ͭ�Q�u9)���T]C��S�'afk�z��	�4�$m9/�3�W�J�f���u�k��KM��D?
g�h܇/�mt�i��$���fJe����z4�2O��ځ酰]��J�J^�X������o�>�Y����ۿ=�N�E��A����v���~�K'{�酷sw��vxU1B�d���v��ܣ�n2�7���[�J��Z�3Kά<�46�d_����1�d��5~���{�';:�e��שq��K�p���L߶��*e���LkS�]D��h툲6��1ު���rI��`�ˉ��P\�W� s'��J�_GcW�*k�d���q���9�R8V�q'�5���߆r��~Ӗ�	]�p�K��KGF�3�}E��ܮ�J���+ܪ����f�q�T��wX~j�#���\n���c:�t�Ou��=P�B�_��A�	
��]�=xuNрi���<a༪�	�ˣd��`��rf7��]9q� ��\�vsr��y���h5�f��Ob��2���vX�d&.+�I����Pӗ��5h`�Ś�i��c�]���J�1e�̩�\ۓ���F�X5.�0�-��s�*�޷�gp��ӎ�1�Lp�*C=�t��}N�>��1k�R�$�0��=H"�f ��ԡ�^/_tv^]�
�/?X�x=�%�����v���epQD���'�$�ÞR�+J����z�]zW��q(�+[qJU?�!��r���F_�ݰ�&�<6>�����N.@ɩ<���)�ʰ��![�r븄|��p��;���l��hz���k�mM����gI�0�D�%Z����|:W[��|��F7f��ܗC)��[�]]�զ��zw	�i�N\:�dT)��uI	\@�"d��qJu��Ga>��Vg�zL��>�K�����;�����ϋ�2W���@�V�'�Rw L�;�4=3���O��qˑ]$�f�_�>�)��¸|��.��S%��?#c"(?��,�� �>0Ȑڦ7\`t�i�ū�q��%z�F\�v��m��k�[MUɸ�'@9�����f�F�T�Y�=9S�����o���:;9
����?q����ya�o�8�ѷ�LV�+x'�^�ٮ�dy��<}�����fPŖ ֬�����(ɵ�e`fPW�5�8�J��<mMEeH�f����t6�ݐr�\վad}��~���-Щ��1����W{]M��˗��f7\�-����������v�����C��=���p��{ٽ' �����	b#�?���S}t��>͔�Ƕ��e��d�7.��Ϫ5Iyz��3zj���?�]���~w�n!�F|o�99q2���NqS�8��'��HW*����l�,��N�v;�9�4�ց;�g��X����1q��N��ݿ(D�����ӟE��-V�	����Rq����6"{U�}
��S���u(�jʞ5���v줛�nI���T�>�q���µ@5���7d_�g���(>QN�1�}\5w�F��p4_�b�BϏnf�D�E�%�*���eq�ەQ�����x}�C/=��>�jX��:���髩��qq�����u��6N�9�Iډ�.�^����w���j�R�OC�,�3�.���}�>�>�~�����>e�6
5
��#���t\k�L�s£�}�0 	�u��������<=V��#�9㸜�T�-%�� oT����<��YΟ*0�#P*�n�AZ�-�gup��5hz���	�i6��N.bP%��l$g�6Y{;I�Ə��"��F�C6���������0_;�!���D�L=C��w6�9;�.�D�'.���eev	D{�p/��>z��0���ѵV&�S>&��{V#|���G�ݵ˙6�W)�n�_��ێ�g��v�t,@�ǗAG��5�5�2j��F��������|^�����0_ГV�.x��"\6� ��q(�3�"�����ә�i�t<��;$Oӎ��,zs*9��F��rz!7\�t�Л<�ob>F3��=x���>������R��UǮ�����ZW?T>��L�)�D�8wI諄+�E�_kUٷ�����j���dɨ�zG��σ��Â�-m�^�6��]~�T���q��ص����-ds�0㓊rnK�;m�Y�/�ޖOW�=0��VqS��g��<���^OM�A�f���|�C��ۿ��{���c�_k��ע�^eN��v���4�#7S��w]Q��<�<��NN���@x���D�w�{_�*�i��=�--�G��6E��d��oy<���p���:��L��S̞�� ���E�<뛓�S�����h�5����qv S�{��}�Y��WI�Ŵ�U����*�.��0��?�����gH�z�o�i�+�g�W�u8�������~�9Z:%T�I֗:	h�}1{j��Z���R�����y��)��i��Z�����F�9�KN��Zgo��nP�i�|���'�8o���of݋o�������0t�R���PǶ���7�uy�4X��^����|��k��2xѡ�Q�'@�o������	qoF;��t{�Tm��՘/���o����ڎq��ږ�z��z�����x�7{$�(���\�M��'�)�,��'ni�m��5�U�R�t�{�t�m\=��a��F�$�A��F�sh��z�?h��y��fˎ��N�;~�B�'x9�uk��^O	��n�����H�מ��Dz3����/�^O�˺\s�ɲ^��G���k늷O���)�|w!:᤼s#�ꐒ5���&�kN��఩Y f�G��-փiw0����˄��}��-�/k�yX!;�|s}s��<'�f>5���O��}�$��ȍ$z%:�WR���F��V�̈́�ܝ~�{ig�{�V�]��G�(�6��׀F�#�\��fB�)��s����i�	S㽎Nf�\��i�{7��ٵRa�Iٓpܸ��G��_����=0���]��T<piڃ�x��Wf��/��Lm����rwr-c��m9`N�
�*A��d�L-����+}�not;�q^������z����~�=	U=>�k��\yՃ��U��z�{#��<,�P�ݯ�Qfʄ�=�ᝄ��33m�C$�ž�������i�f���@�pi#�3����V��e�H��<�B�iP�bK�f�6ìV	��]^�uc 'oe�=9N������1�RK�Yע֜�ugM�\s���
7�9��^�ik-z�{��l,�ݠ��\�Ѡ�M�(;��Wه �!|r�����k���>|��ice FcY��;r���xg��<����z���ֳ,-�^�C�-FcŊJTc�X��VN�`��F�:Uޭp�U���x�^L+0�z��)�3��r���*y���'�{c�e�1�vhx]ĩ�U���e:W\��:�V�e�x-�����������7/�����B>��<8o(\M/ebf��-h��2�f���D��t۷�9�Uz��S�"�mb۾mS�F��^��=5N��v:od�����w!`ox7
}!̍J*p����/:���0�]Ь�+�-�dE�,h��[�Z5�U�z��B�a(]0J�OTZ��ޟ�k�n�7d��9FY,OOw����\њv�$�����v�ŨF�wF��0��z�;��Ȅf�k�����%7��X�]>��/�MQծK�;�c!�yd�w���b�:�Q�1p*��3���*�(���Hֳ���.�pKC��뛂�wk��1��|��j�N��Um,a��]pQ���,����د�2"B�V:8�����������N���U����'����M׉�ʏ)J��ݕ"d��V���@8d7O�e���A,m��{�ڹb��8����ީ�//28�F�ǒ�r�#�<�U����q̾<�k#*+�q��C�k�#�����%^�5����l�	ىq�яNI+�΍D��N��aR��4Cɘ,i��8�f_\�4h=����j�iSc:]�z��*�4�Zl��ݼ�i�X.]������!2��y*SL�zN�-MQb�<*�|�r��򆫅�`*>ޭd�)vz$�ܔ����U(���ċ���̘�]w(eF����TT�kj�X�ǻ����D+{s�3Ԇ���Q�)����}�Pd�8Y�����S6I'*e=��n�j�7�1i��	��朙�t��'��-&w�?��9�Hr���h\�:^��(Z�gU�]򍭧�ǖ`gA�siM��Y	��ǝ��`*d7��^��C-�U��������1-J���V�1l
e�L���J��\��"C��Mx={Cڱ������ݯ�{���.h �,�-�w���mK��;Rs�A��1j1w'1.�˫����/I���AXzLA�:�����pwK)�mw ��ъ�N��\���î��%�+v�B	;L&-�\wimp�
�Ҳ9��OlMX5���oW��)��%kW���#à����	�H��G|��.[Hs�)�I(�$�\�I�˃�$�!PqS��n��)P�ո�"����$U�ha
��'���(�5�C��q�E�u\m�$���\%��Q�B��ȓ����i��2Ԫ=D��BM%�n8���Zr β��	]#b1ęBN	%�R!:E2,�M��4���N�LТ5HLTL�W(���jQfDDJ"I!%g,�:W
i%Eŕ�B,%S�T�EE�	U�GN�I�2�$���J*�q��D$�9Z��p��Y��)3V�(��4��VR.���T��<�BeUTqM�ge�j�D�;I!+����~林NV���:���;r))*)�x��t��/j�g��W6�WCC橪X�{���>f��k��q�{�A���wVe���L���?���Y_#~5/IӋ�3�:US�yK�TCWQ;���7�3�1B�����,X��+�zp+��V�5<���9*Gc�Q�e����=��S>�g���TӜ��T������f��N���%�n�Z9���=������s��N;�u;�Y��1�.SE��t��E.���7z�\gz�M�Yd����gJS/��1Fݭ>ˌ��J�Ƨ�p��
ǝ0E�`T�{��3���p}�SY�-w�Q����3	�羚���ڪ��g���V�:��7��
j�Ѕ�x<q-�� <n�,=>�OQ-��V�KʔlVm����,�z�ź�te��uQ,�+[qV�[�̆�F:�y�##��b趮';wկ�r�n�r��TԖ���#ܶ�.�T){���9��~+�Sk,��#&b����^:�-�u��#.+�єH(�Az�@iN��L��q\yoWƭj��v!l����;��ǖaÜV�ϋ��nw�e��J=$�����}4.)N���EO��5뙘�Z��`]��r�:w�ϖƬ>��g�9��(�ea�^-���$ֹ��Z��؟I;|�v;v��).��7r�2�`[ќ�e�V���k�pϷz�Z�gӏ�������6�i�^�}k�2{j�]BF<���ly����ll�%�׽�F�]l!�/���.q���N�	���=~�����GS�2�f��U����8�tz�Qq�8�kк�v�YZ}w"㒦K�r���n<|��A��Q:�o�3�{�~��5�x���Rއ��Y�TT���˞gk��M���jjO}��7��4�#47�w������U/��>�n���rR��ô�6���N�|~��/��^Xx��|p�P��}4@G{��^��~k�m
�w�.^���>�:�d�W�c/����4�T{o��>��~Y���h~Kkk�Ƽ�'�����N�?ךo�|���qg'/�㡋�5l����aU����ݩWq����/u�*y�C��{���ϕ�"��ʝ6�'v������>},,��4tn���ђ�{���D쁼�e0+��/��h+�G����ߵ�g[ZeC���Տ�5�Է�22�2���7�1n)�3m��|6�0��.�7;�n�k���U��i���v�����}\�Q�'K��ў�we��*��UGF9^.1�e����{�!�zvj��w�jMa�u�3S�_��������0G�:]^X�E����4Ng`!����սêl�y:�x�i�&coK+�%�;�c��'�^M��bf�]-���;��Y���S7G �(3���3Qޫn�93%T>B��Ҹe�pnd��;NI�2K���/�A���W��N���}P������E|�U���ޓO��ë�^���n�(��dqۅ�p���/�P@ި2��<@=�Eƻ�̟j�O}��W���nc��S��m���'���\�;p��NK�F��(�}�@�p
[${i0��а{|��=�}����������V�����']���q8n:���d�_qȰ�̀��~y�����dÝ�:7G4���j�ox��V�.x��"[n���q1~a�}vw$��%�}[�:ɚp��#�=���Z}Y�q���*6�u�6���� ǫ*G�zz�g��������`.�A���N��3����pVz��>��ZW?T4��J��xtc�g̬�f��]�oO��h�)5��P���ɓ]0�MJp�9=��#-m�^ͥ�2h:�7qo�߫;�F�F���L{�rnK�;Cw�n4�3㡓����끕�_�/7�5���5>�����i�����I��L/mU�6���F'C\��u`����.,�S����ݿ�*D/-�^+Wbה���ܬ��V�Sk�����tH�z	M):�]u)�h�n�r��t̾.�����Eir��G�}��g�{���-���MsY�q����h���S;�o��B�7�m����B��Ҭa�7:�����������o�vM`
��aĪw���b=�U���]���=�障�'񱸷�~�8��x�{P�+�XlԶOFJ w��
y�7&\Ǟ�&�Gduk�tL���~���{�����Ϥ����/��Fv��)�q�*G��
��iO2�k�wHF�yST�9�����<{�_;���X�9'����v�g���΅u2�b�mP�6�Յ�����R1�ɪu��׶1�.�����z)����5�n�F���є�	=<3c��Nn�_��K��Kx	s����b�s�4{�p��c�ζ�r��c���� �Uq���$�ڞ�s�Lͦ������^��v�{ET������k��m�p�-Ө|.K9���L)�̻�cϹ�¶���:�R�ǠI�&�l��#A�~}�V>��(g'�u?���p�Ԍ�S<c��F{�u�{-��4I��� �!�.%*�o�V���\mo
����|�sKg�P5o7Bf���x��^Iec@��ݷ�q�g>S$��R8vH�N�U�T�83�g�[�c)�{��6����!��p�G��y�m̫i��ř��1Z������2����%�)���}ۻ�d��[g���,}��8�*���-�0���[�o+�&�w�S�X��{��f���7M��{#eG��J=�4G6d�:�X��D��s�>GQ<B6�N�Jm+�T����p:�*T�4.=n�MA��!�5�~Ν�!f���B����L$�-�#Z�>����H�z�!���ƣ���Yk�zWW��ޗ�����f�k���'w"�:�Ӗ������Op�ztW���G�W������.�	�0�)�a�+K�޶4_��ly*��k��'�bp�,�	��#�K�s�M�~�{uX�"�t�r��23&�^��IXO�Gl�n=��ǥU<'�ʘ֧<$x`v�U�{=վ��7{N'�fy��Z�n}�������,���>-w�x���\5��Dv�6{ݵ�~ч{v�P�K������%�|�Q��2ga|Nٗ	�X*~��f�G�si��{`��3��WHh
cr�6�s,D;��z�\n���b�S�������Δ$�0F��핞X�p{wy{��Qq��4��#�yRv({�:L����ϸƆ����Ğ��'A��"Eu���^ �� ��qS9������[����c��7h=>�U��%R;DL����ߴcA�iȵ��������S��*�T�l253:<�q��kΛ�x$�;��t��Nc��_Ƴ�*(���<����9�/����	2���G�t���U�S.�9�N�ca{F�څBT�ź;h�N��>�-��[��s9�B��M9C��y���u�z�v��"���l���O������J�s���9�O�I�5P�a��/x	�{�S���W`�.��7������0n �_eX\|���9u�oӞ�k[�1�>'u{�Wkw��a��F��;��摔H(��z&@-*�`&x^��\{�r���s���t��X��]�5�장���h�s�M�n�q̳#�F�����'�Mt¢Z��]>泺-�8㌰�����[{�/���.q���`��BT'�D�_f�o*(*���=����w�}/k�6\���J�}~�;!�O��_��S%��?B7�O� ����Y�{z|�K;ך��2���ꊝ��>�.[;^�ۅ��\���&��ߓ��v���i��y��ѕ;����?O��.�i:��Q�c�S���"|~G�zXזUi�jć��B��l��fwMy ��T�X�徱|_�}���O�����O��g]-'O�e3y����ET��n���3��rw�k�vk�ǹ��ec븝��v�3�|Y���e�чʟQ�k���|��wu,�4�X���G��OH�i�]y�Y�v���ޣ�M:V	�b�=;�����%��&�5_�]A��X��?#m��K�A�nܳ��{Hv���/�:�oF4c��
G�=ԝ��yg.P!`�Z�p��<�|k~U��m6�z�E���O�v�
�}�c�J�~`�C��{�Ս�՜c����_�I��$;���F���9��{,����	�/�]@>��)�]���J�n;���t����u(�5eO"�ag*��khfھ���L�0�����q��T^T^�cvE����r� ׾�|��s*�G1T���׉\��j�Bqs��5��f��B��/��ʁ(��w�5���ry_z��fg�\��E�e�uۉޗM��e�^�l�P�A'je0T+����}޺�n��E;�Ʌ�M�_�"=��lc���{'����!��y�}kp(r7��GO_�t]�pkT��F��S[�)���W
�T�G-v����a׎�}�S�F�\�k�� o� y�er�~�[�ޓ7��Е\���p���]p�Κ�=sm��N�I�7pp�ΝD�2Q���F��N[���wݻ���'	��z���{�P����FI�C����N�� ���s��;���}��|'�re_���l�1/iѸ�+NV�G2���(�]nM����m�ɨ�Zh��{�1!�Χ�Uִ'M�?{s���5�2 l�Yv�Έ��]I�.�eB{Zo���Jdt��;J6�+�=-�汿���k�'�a�1��9h�ak ��V�?�qb��]�ܒ��r��=i�7��5��3ַn�Ol�v�@�k�T+�t�tT���c�J��W�����ﻥi\�P��ށu�P�t��ѫH�\oO2h��|�P��l��5�L#�<P��9�wS�p\e��*����P�^�lT������*�9�N�Lbq.J���N���Y��f�id�}��ᕁ?CG.�A��y'gC�<�}H��mp~ګ%/.'C\���M�5�fϒ�@����6�^w����QW�moڇ��=�?�YK��u�w=嶀x���J�x�V#ޅ�ct���\��)��9)� 7C{�ۨ�r<�Y9�ax�}P��8D��ށ������u��ϩ�c骐G�UNH;�~����r�g��{r~��h����Iz�+]t��{r�4|v\哽c^/+X�1\�������
M�Ქ�Ff��|�q�:6�I:O�3�\T���T%HT�$���~J�ѕ��o�k���7(�����3ަ���5�n�F��H;FP�moL{|RЧ+!贲�@�a�]��n�U���=���t���p�Ц��~%GI=��f�r��st4���G��>&"}���$�v��1�OX��+���;K{�.w�1H�0�k+>O�����MTl�;���:s���ć���`/-Ye@���Ս)�a��\y6���In��t�����靷4��,��7�R�C�>� "�N���U�^�B�'x=�i���aۇ��p�7n���\���v�s�,�jeDڃ0�L�I���{ވ�P����p���yNS��u�Is]Ӧ���Y�*w�mfg3~r<�T��l�S� ��rD�)V���xuB�kxTe�N�7��g6�ó��wW���f�E���m�xß35
d�+�R7d����]JӃ=�y�)Lp�7L���=�r�wfғȭ%\���׀�Sh�Q�*vn�s���Q�h
�N�3�#�=H�߽{{�x	z�<�zo�Έv�]ɋI;2n�_�F�ѥْ}�N�L-���(E�����7kw�i��J��t�ף6��]w���;���A����v���~����ԇ��\s�M�wCD��l���c��f��z_f����WL%2��)ӈyV'�o�SÐ�X�y֫&�����ws"ڝ'*�L�A̠�
����:p.��gZ������3o7��z1r����;��Ԧ��ħ��;Y�Rϖ,���g��0~�~5�v�_�ib4y��c��H�[�f����t��J��Fy���A��������1���#�Z�-�ƍ��8�0�߄1��7��y{Ycot5gb��K^���u=���q×\� Z̓�Bw���	oz8��G�=�4��˾�z��ޝE!�v3:��3�>�=�[�}'9ƿ�f�l�;�g��j����f��N�������Z:5���{&~��f�s�&���S��;:\v�Jy�
wI��.����ޣ��7e��fP�r=����W��	���vlI;��V�2�6hu�*@�����t��E:����]�l��c���:����L����FU1T��{wHR�//X��kw��c�l��o���z7}Yxba�K����={݃^@�:X�K���]Com\K7
��U�*V��!��2h�a�~�7S�K��\_��q����T��5%?��`�U����+V7�J��#�D.����;��Y>Ei�NF���e�N���2
5�F���@?|ҭ��K�e�ɃO��^�u�p���Û��:v��9Ͷ�|\�p۸���T̊S%���D��D�c�u/�|nm�wCUSA�l�s�3(+[�F�]l!�r��>.w�^|h`��	�#.:���4%4>��~�K�8|:؉�"�8�Q�-l��:��qc����S%�\F)�x <<m���cm���cm�c ck �������1�����m�� 1�����m���cm�s co�01�� ���1����m����������1������ co���~�1����d�Mf��qMf�A@��̟\�%o�y%����H��J�T�PQ
���@�*J*�����%��""!")Q*�H���H�����B��T��R���$B��@(R�EJ���4T"UB U(ٔ�*�T�A�͵Bh�D�{p!U J�)D�UIA ��I"��H�"JR�UERP�RJ��RB�@�HK�5I�%J��T�%@�ґIRL  ,�W�]�J�ݡ]�[\hnU��T-�8�MR��]����u�X�����՘1�kUkNBƊ�Z\�ηUZ&�R�U	�P(�AW�  C{�(
n�[��l�ݔq�m���]�Ѣk�Ǝ�Q@PJ� ��@ =�4   [�{x��F�F���h��@h躎�F�4h���U=j��!�UJ�(��   �wG�mF���)Ԗ�#V�m��C�6CZ�MvQ���*����ڃ��:V��9���ֈ�jkj��%��"���W�   C�B�j�-U��Y��g]�Ѧ���M-��[�lr��Ӹ΅N�-����wd�w;:�;�����jW]��ۮ����T�n�� �
$�T��TJ���   Ǻ��p�]ˮuT�ܮ-X�vQ-��vѷmv�m��tc�t��v��8��it�7Y����;�]�M��ݶ���F�.�ͷsL�F��Mm��*t�T��)ID�T��   {Ԓ�r��ݶ��QM;�4���rt��ݵS��ꃪ4�e�Y��˳�lw9+vˡ�ܪ�N��S��8֪�S�k[mݹ�t�wmD�$�
Q�BP�   #�7��Ww�����m�
\�U�N�uݹ�;J�jfɶqm(1�5ٝmR	��r&�ۮ��Un��%ذv+�K-gpjsw6��l�tUAR�)BEUER)�  �{E�I-W�㻭��ˍU���慭Sgm���l:�s$��Z�v5��gMZ�[��ܖ�R[%����J����C�ݮ�sf��v��U�[h�QP�I4d��B� �����nݻ�4�ۧGM�k�b����]�5l[���n�i���wn�kn��Ԯ��c������5�V�F�S��v��*:�U�-Ĩ�@���*�QA�  =�^�[����qRv��n��N �r�]��u�YmZ���t�sD�WQխ!�v�rۦʒ�Ví�7wv�u���i�lൖ��u5���.��{M&eR���d �{FRT��#@�d��(� )� �*   "���MUE  �&���L���a�&���a�@bDI���	�J��������k~k�0$�	'5��B�$! ����IO�$ I?�	!H��BC����|�|D�3������)-.�3m�m���ˬ���S�؃&"tX�Wv1.�kHH�XvV�lb��c�or��h��ݍ�mG��/]]�u5b
9�h�i����LmS{wQ���X����ڃnUڴ����h��)�:����
����e��ÅF���p�P���[�Wn榮1w���R�Ҵ-��ã�Wiܠ��n=kc 7)en
J��C�U4YU2��R�Ű�:8l���4�4,��5�C���W
�E+��y/�L�F�ŭ�3����oBh=y�wKkt��c��=ۤS��!�F��ɷN�²�ԧ������IbA�G��`�&+R[dlB �Ne��P�&�JM����%ZY� %W���3g]5��5�E�JB�ń٥n�yz	�p0m�"32�c.h)�ca[Osi�;�L����a�y+hL���J��w ��M�PڷAP��5�h�F&��O@��YZ�}4^��!*�)<wz�-G�Ri�"�JV�q:����H��l�4D]��j��wK)i)mh1 �49zQ��5�E�r�;��[#Of̉m�a�@�M	�ael��r�F`��+Ni����K7HT�݈2AZfPz�i`m��%����+&2�!�)���Z��s,�cr�����'N�]fi�Wg���L�T[U�E�l��s6bկm��S����F�jq�nYKN����K��n�I�M�
!�G�f@L��R��U�N���"��Z�ֳ��{k*/�H��dw�[��!�Kd:"�����欢��ƌa�VGZ��:;F�o�1�-'h@���ee�"�ЉW�b��if�eS
�(f&]Lsr���NM��L�٠�%4�˼t2�6��Ab�4����0ٔ�ayV�d��?-�R��qE��`�h�U��
.�=ݬP��\wom�T�h��׃$�51��I����ۖD�,q{�k;lY$�q��Z���"��ֱ���XXl^ܫ��$��	�j����ǆ��F	�l
y��5Y/C?Ln�#aĘ�(�/����tS8�B&�7MQIZ�8w+I^)n��f�#���XwC(���]䧎j�*\��A�^��ե��D{���AeR��R���{�&8���&^�lĝƞf�H�(�HfҺ��u�&���.��S��V餷v��EVʒX�5k>�p�@s	�`�蛭�$fD��EZv[y����3&��vX'��xp �N����e�Q	Kqm��r��S�,��e��@�*t��+"NZ����lA��������J�j��Lb�W@J٧(���Z)��%��ݫܗ`�M�*,�Ŏ�̲	m
�j����@*2b�Z6����M+LB��q���+�&-���V���2,��VԶޅ��ݿ�l(�P��eGd��5ՌXڔ���ܔ�ѐ�9��1U�eT~�գq���4N<r��r�Ĳ��L�.�k2��E�dx��<_0�Yև�;��c��&jY�E����0���o��˧����ȷAM���;H����ieeO����֜�Mk�]be"�6im�$�{o1�p����@T�q5t�Q�v�f�6!��)�S6���7Rȧ�$-�ׯ�N�H �F�
�Ѻ~&&�O��fb�u�(o�@ȝ�T]m]-�)0n�o&�ԍ��Pկ���bM�c�6%Zssi��CC�6n!��X�h����MV��i܆-%���N6l&��р]������U���w��ͻt%T���j�cRf?��B��#�f'��J�Լ2��uN���m�/-�
���2�\�5Lj�z�JQ�j=���V�y��Ь�-j�2墦ݗP&1`ǛV�{�{�è ޵��``V��/ A#�ec�ca0X�t�Ң�!��/6�`P"�+�
Y��4�q
#h�H+ŷr嫣7+h�|�5N^�Ȓ��$�-����C��[&�A�x���Gy�JD㡵CX�i!���`�mީf��v+]J�X��J��,���_�4�[5�cb��ߴJ�WQ�E뫬[D��\����3a��n^х�w�L�OKJ����2�L�E6�|6�T�֡jͳ�*qj�L&���!�CC�01f���V�EVNh�XZ�Mu��`�֧W
f)Dּ�*L���:�5�h��Ể�,����JU�6�U!���1�K�ڙN�*�nd��*��{���q��j�3f�����rm��j���L"�.�uj�cn��Ă���>��XZdR�n�Y�j���$�E�)�)jj���)�o/��0��y��WO�3�Â<�P�Q`�T��<���X�S4�N�7G�P��AA���Xt�3]`�rfPwzh�}�γ1��B�|c�H7LS��Kt�ڇa��"�B���y��klU2�Ӹ7uj����P8-l{m��[Zd��,�{����G6R����#���ɷ,��D�h�uy�(��K���S/t˩܃\�Бh��kt��Ջ�sqR����U�J��;u�B��n�]#�pB�F�n��%�B�ؚ��ΓKu�X��!m��]�	b�A�U�Tj��I۔��f��� �LX����(�J�CХ��s�al"Z&U�6�4n�ݛm�o2�f�s��7Iؕ��5N�bYYuo�[!�ښE���z�m�a���]�� �
0b��n#J���>9J���A�B�ֶq�nLNMQ�7�1�g
�eX��F���c �^<��N�i��hR����,αo[@���b��H^!i��XhM����a����l��%�;�;;�[H��:y���:�7[z�͢�%��ʹk7e��%p��`�f;�r�7t3�X����@]r2���<�0�е�S��-lS��!'�V��f#��˵����iL)Z U�se�^j��N�ꅦ��/+!v,-��sN��BqLn�v��֖�2�ˇ1�Y�j��Jyw��RV���Q=Xq�b�l�^*����l[�!T7+b�[���u��׶)kVVZ'E��
z�n�k¶"<6F���ڗm�٠7Nfq0����`�ߠ�cL'�`��"�,�s.�75�F��%�#d÷371��D� �N��]�Uk��銽��qS �ת]`�@�i�������+�[uGk�7��3�9��n�Fd��(�9G 6�jr֛�+oqRJ�)��c���SF;��Ƶ��+�6��W>I^kZ��Ų�G�[�p��̑L�U�a�I��+�,#��0�QѢ����7�˼I�kq��waB6�v@b(�:IYf���wa�j����n8`2���1e��J�Q�ww�ر뎝�*�X(c�r�w^�4
A+���
�p��`,�1�j��'0���*�5����)��n�Yq�Uv�j�3h��"ҽ�Ю� �б�(�eȕ�0,;�)���=�frTK���j��4���	��[��ضE�j�41�]3kJ�&�{	ve�n;���(fb!<z_�2Y���V�Ź[�Z�*t)L�`�Vô�f9I5'��Q9�v�j�� kE����2]b-��o�{�`�B�r�=3]!6�G��+]=�t��Λ��	�c5�Q�����7�4�S�r�����pkre17��n^0"��j�S�xYw��'��B��t%XB0�V��KwH���f�쐓��ChJ4i��ؙB�����7%����%6��/hJv˫;k`z��=EK��3b�f֝�����_6���F&�v���h���Cu�)��	vtm���WRm��5,u��n���֕�6�V��wn��ކ!�ǈ��M*Z�Q��Kڏ�7�*\�9�S;5a/\���%��mDn�A)��ͺ� �$�� ."��PAa-(����c^K2�kj�=��į���K�NV�8�#�c�Pq`�m��t�Cn�8�(�5��ǰT���k`r��C�����Y�e,O%�Ǣ����!j��5|	zRJ�͹��w�wJKH��mܹX�똖�!x�}t�yD�J�d� n�,3>�?�ҭm�+M7)S]<�7 x�-��[��U���SN`����n�9�{=�͔����˼/E$�M؉屨��x�����\�m16�T�Ѹ�4�mM�y����ZZ#�J��Mn�����Tb�w&�b�e���+���,PB��EbB�\&�`�h������/Hۀî�̃i��.+xjⰍ\�z�3u%k?���u�&������\���H%�HQw�g0�aˉ��[1���P�]�4\�5�cUv~Y����Oef���f�$/e%Pn=)aN`�n�M���5埪],����Ƈ"�w�]�x����7��H�QCI[�K���0��fV<�+ �T�~@ei�����Z�NA� ��ǹ�h9 �iԂ�m,bȺw5��<�{V���,Vճ%�:�Re��m-7P����WN�کNn��o[)L#U{x�i��lْ�K@�}j5����`Y5�(*q�)�e'x�9L�6މI��J�2m�ת�)�F�Z+)�enʈ�ʛ���J�����Qx�WR�-���^�r����"P�Pd[�y���E��l=v�TlDW�dY/��{(�&��޽��&�0��p`xlXG t�VT�&�����\��Z�����r�4E2��X�,rjخ T�&�Ul��j$���V��4�����N�A,޻U�0�2۱76
��KZ�r^d�)��S�+Y*��x"Q�$�Y��2�����L�9I[�����yK��,M`�7��=Wn��j�JkߌHC��8���, �������3k$�@�����-���.�ݗj�+R�%�OY�e�74��CI�𙲝�D�؊����Ɗ!�AÊ�֭�n3x�ƌ��n
-�WB՚{k�+�/�S� XA���KŴ�.��ғ�rU�t���Ș'D[r`����l�B �GAme�{�=i�orf�f��٭ؤ�+�*VS�%��s(�Y������HȔ���y���wI;J�ʎ��&��i[�{JU�W�j�u,/�4�P�&��"��A���Z�����9F�L �x��z�)e�[��u.��Ra�I޹�:-%@�v�X_^ʚ*�ݩCt,t�%��vi+��̤���1b�i�:�G2�2�+�����^땎�Nf�ʁ�Ũ��
OK�YJ��-�͟�
�*��lf���ùSjڶb�����Y˽� �)'��j�&йSf�1���.�W��Nk����,[�m%�GYx0c�%ܢE�M�����֤ճ,�MnPb����Y�ӭV)�Դ�R�۸�C�Um�w!U1@�.n��f�3����Cpi�(X���A / b��Wcwh%�2�.�.8Q���u+7R}���n!� ���L݈P-���ʘP\Cm(�U��Áֱi�QL&P�ol�`����*�)�r���^GB�j�e��r��Ե 9�ـ%�
6��݉�jLeJ��#J��v6�Q�T�X��`��(&N
Ã� ���N\�է��L�o��J�D+�Tl�FAF��ԭ_v�F�P�y�\�T����-+;�wf�gDNm5m�x�6������(�*�33N�LV^V�ul��ʔ�F:@�6��`�Z��4�T�i]��{���5�vV�f;��IGr��`MZ�-f���_K0�m�56bw��µ���G^��Z
����Lm�b���O^]14���N�k̚	D�c[{�Y�n:&�ȋN%O68-nlx/M�2=��-Qїݰ⨦@�ڹy
e��n�qh�b�9� ��6�m�m�.]�FQ*����7{�m\hM/�4�P�D�N��Va���P��̍!�X���WDl(Yj�ʌt����c1@4���yD�0��$%I�.Y��3m��,a�k	�Or����@�E�ǋ,�Y�L(oNo�@L�E[t2��H�Z�`��s�ө��1��� "�Z�����[ێ��^�i�M�J�Sa���`���^�9�F��v5��y
+`b���g@�Rj���Xn���/13[7mO�x_d�m^�˟2Ƥ���ڵ!��I���
��=8���`�]& ����)]7�;��Xrԫ�c�)MNI�k6!�<R���H�lK�	���-��Z	Z�U,Ńln�����ܦ�3�B��yZsD�,`���!Y1[*�6�^��j�نS ә�e����P�X�M҈5u��K�]��]�kY���4Ć�zk֧�S1�rU����7w����7)��ӎ���x�Grm[V1iM3rAtH�bXk$� �a�Ģ��4'��D��Xu�cY��h�o"�aTm�������t��Y.nb��k&*D�H11!���⢆��+Xzu�of��!���N�Z�УtXa��4��uoQt-��IT���ç�[�Qt��F�FXqRYx.B�%���A�����J�����m�+p�t^K4[ci[�[ �e��J�ay62D)	͔$���%Z�vvjˍ�6�I��ܙW�3�lbU��ķU�t���J���1z�]Y�'�s\c0�5ynj1^��3nҖ�(�d:����`��	�e:��z0eͷ�Q����(J�I�>I������2�ݚSE+v)�	��� uX ��^b��(Yy����:�n�з7/0;T���-�a�����iem*�Z63��9���(`�VU�C�JeŸ zm6FYw��t���jm�����T]��̩׊�k�����p���u��oc��i�.�
�J�PA�8w�cƺ�F:}�z;X�T�Lю�NLR�-*��C�p�ټ�����]�(^�ɽ��rӰ3ȷ
Bk�i��\[��&��M\6�-��|�J��W�]c;C;#$�'oAv@{-7*6�a�!ʜu�r��,�)���KF�YB0)���m<���N�E�V⻮t�����f��j��\<�ouh�|��v��Y���8��V�v��G$հ�GaT�s%�����κ�X���aJcc*T|wl����u��0�}�����{�uuۅ�a3L05�v�<f;���[*C%t�u��㽑QEY��{�����;Oo-.&!���Cye�n�$�`n������'hű���Җx�1ܷR��xWA,��C�E��yf��9��7������T�7�7y�y���xd�i'a�P���;9:@_s�T.��y5Bm������>����ܷ8��-��Aʽy���c	�䞪\72�n^U�����:L�i�i}
��L�Nf������y[Nܾ���d���-\n�*1��Wv9֞ɚ��[ԟp�Oz}�B�������d��^&i�:���u���f�����&�u,�4��m;�WSkx<��ut�����/{uC@�pA+$))���V����t�u|����-���H7+��ھr�ϭw�T���Q��0R�7.Ț�0��3��ZTj�0mn��Mnv�EiȸXk��aVR���uq�T��A�&:�ti�4�*�n*�p�SѢ����[��+����v)R*��}�Z1f'��/+>�}�2�f1�ae�l�V7��m��P�\�;�:�f���fc�u�l�w��Ҁ�.����+x'M����1Iz��]���[:�1�m1��ܸ݁;hx�0����m������VG���^�>0�Ʃ���H.�ֻF�1����=e�֨ı�K�g���v�ę����c��v��r+�^���/��"Z�ɫ���]v���/eb��e��I�˛˨2r�#��T�ok�y�N�`X����N�TOO�A{����Vj1���i������@j�;�� а�قGj�������aзth<=���{��2:~��r�ݯ��h�R������X-MT�,�0��x�n5�E<��rJ�ӬE��ɕ������BA�v�\���'J;B����,��ƼҞ���Օlφ�:��Ӵz��W�\+��ͺ �taf��i؇#5;,���OuW+H��{��(>7�Vu@�Kg���ֱ���PfVpO��]8����ס��]#.&�N�Ζ�t�wC{Q�[�v�Ӭ�
��"#*��6`�z�����4��S��<�`�}v<ø�y�,�l�5]+W�
�n������rY�ͬ�u"�Mb��s�����O�GV���8�����Zi���:y2\��OPP��GM.�6��Zo1H�-��H�ee�SXr���]�FZ���fh��o���<�I]�Y�V�>{�1/�f�=X3�S����F20#�)�\�Gv���C����ξ���zec�a����%[�DŚ\��zr�J}]2���0�[[���0�����KK��#[�a��D�L�@8�T�Vo��ڝ�f�s�۽O��1�������3o14�t��V��8o+�:ݳ�X�Q��ۢ��w6�w(�c��kj��H�����w�YS^d��8t�)�uGlm��ë��mvLw5&R]�]^	��b[Ц��/vn���,��rE�ξ��:�8�U���BH-W�yqe�|���+���=B���±�k�A�̗�3������rb�Ũ�S)�%����ݬ��$չaD�(�#4E��/O[Gut�C������:u���	�(�8�,>����}�9�fj�;���Y4؋�ϸ��Z�v+��9>�ڛ-��ZW�-�
��K9��0L鎳l*5�Q�NU�X��ݪ���� �N���v�Mz!gif�q�3�*���wWG
q!prӋg��,�"�r]Ijc'j��!{[�|�����c�ִ��2���75�E�\�Ӑo$s#��H�m��A��wE�(^��n�}��b�����x���\��3E�$e鷕d܊S�"��|���qXN�9����/<����I�n獎Nh�q�Nt�1��s��x�t����N,�=7�Fwn�՜�g�����A��#����Q���t��ke�]�����-�V�8?�:N�-,t,f�_����{9�E�2Һ�c�����r!]6f�}��`�f͏�Tڵx����9w���S�a'+�H1\�z�|9d��Ybݗ����z���0_P0���d�K.��EK�uZm��gM҆�B �/LR�mGϺ�R=qUۢ�'u<6�c�X�b.��蔬u�ʕt:�d�θ6��6�/C���)��N�^�!��u ���T�ehݭ� n �[��Y���z���3�e.��s�tt�w��l��h�@�*1�B ��olˡ�'.���|M�v�X�ŪB��ɝ}�ޔ;'��.ݸ@=ͼH.WV���NX/4s~��9�o&�y*,	1�`G�#ա ���7u��DŹ)%�`X��p�֕wt�m|n�;X�Ϟ񘉆��Bƨ_�˧\�y�ݣ�}W�սGT]]�Zخ�ϊ�_'�w�IHKU%_�n��p�bVHodT��"�h�k�W,����uֶ��ް�����t0`vG'zjl}�=��u��r�#G3No$��6%!����K��Gv�8E�
oy_욫̦�
뾥�+��˙3-ǊbZ�;X���i��D�n�R�͆�UʻcWHeRUh�9w%��$�]����i��0h���h�ͥ�9*���]�
�5�[�+x�/�E�XΏ�:м�re�'״݃�)��-*N��j�����\u9j��*��`ڕ!B�۹��]7�����,'7RY��m�D��p�M���Q=-n�uw�NQ��L�e���3�7 �����jF8wU���]�-��ͽ܋7n����W+���w���c��6�e	N�*�n����]>�e�;��dR��k8��,�qe�ӗ�)&-��Z{����BƖ2�R:�M�	K�Eӻ\r�y �4#�(ۖ�7�8���o�|��S��n�w3�1���+�[r1��p�#7�tp��9�n��˨���0)��;��(���Iuֈ�m�m��Eiƞn;	�J,�(.�.{&��=��:��ތwPπ�;�ksu)q�a�bS:�rm���]��Rg��Ceۉ��?�aD��ۓ:,D��v��C�M���Z8�IL^�d�)��k�a��k���;��"�>XӯZ�0w	s�5���Lu:w�V��4�c��w/��W�
t�ie��r��;!���]�p������CZơ8r�L�·�qIX��J�H)u+���v��g^P���ݠ�����o�����1s�F$���g�c�ڌ8>7Cɼ�M�b���������ڼ�}�=ℕ�2�A�����V�3*줬��o�CNN��:�
ܲښ*!��֖e�.��B�y��H�"�K�!�u&�w;4��L��,e��7�w$�z�����0���ㅇ҉�o�-���s���Hj����9�[���|.�e8w	���4�Ɲ=�mM!�W���N�qD����J=��-wYZ��27oA�yU�ј|��F�O������kF�|�K�M�<*v���}˹\$��3U)�e�^d�/�%�K*�7x�E���Zì��W�Et��I�&�4s�'�tX�C,�rY���wj�u}��ფ��z�ZEֳ,Zv��9�䔖�!��N
�r�ȊV�e�B���C6����e�v;�������ݮr�QJ=���˛��|x:�f�p}SM_^�}�Η��'���t\t$�^�/��SyG���j�E�O�2�J���U�me^r:��m񱠡��,�R|9���ြ9Y]s��mnws'����웑�5��j�.�C��4+�7.��u�e�ۗ9�kkǆv�ƥzxV�tc=Cn�5�na�4EPԘ��N<��(MT�L��L�|�X��ͷ������w��d�+öĦ12[5%�n�q�n;�iFz��榪Q�2����81�9:�k���S%,��Tedl��#	��mh̷oB�^���ok��Z����7z)�����.^�{;k_#K�f��ʔZ�g�v��:%̬P���pX`����usuz�	v~(d�<�b��L�c8��E�{Ij5�i��;��}pP�$"�r�H+�1IAƶ0���eɆص�����t��v���/�m�{���Cx&�����GdJ��&Y!�.�=�v֞��u6�ҫ�*϶��U�\��uǴ�byV띸;*+�,���tE���g�.5������+6�����4\�u��&���Cv��B6U�R�S�[ߕn��:�]�H���@�!���C!��Ls���'��6s��u�A��]�\���L��Xη;��ջ��f��ó])�o�4@P�ս��W��9Gq� ��x�fs]�R�W3x#Ǻt�:�e.6�[+zu7;���/v�v{��S������a�C�)��u&�q��E3y�r�c�Vv�o�u�T�n�[sP� �M#�+[!��������?b�J+X�`�h�6�p��O��@�� ��Y8nM���$24�Ʈk9��V��2������kQ�t��t������6^��ew�-���9D�L9K�P;Y\ �0$�z��\�^���/�m��{���]�Wu��@mGӖ�;0`�D����9X�!M��yA���	N�y`y�SPW�2;��S�r�՝zr�9��\���]{��%�G���O-�-PSq�v����R�HL'�3KUz:�v�N4~<l�&�;\�J���BwPMr�خ7��%sr�w�j�� �zmq�o�V9�\5z(Q���ѶA�[}[�k3S��q��Q�'�f^{r�ݮ�4�W����*������S�~�W>V��&f���k:2�c����(u��֩C��yίq��Ȟ�+1�)�k��g�}3���|K�� "fnq��}��Y�V��:����W���U��:s����;yh��=�ح%�'��v)�V7���Oo-ʹ��m���o>yݤEOo�
ű{��5�+ H��J]L�S�+3.�_V��A��J��O��.F���%E]��+��Ҹ^��w���nX���-2��W����Y
��WTk()���v˝�B\�n��r��(u2��'w�CA�B� s��u-�K{��7mvL�y4�([�Ц˧XɛiC�����%�!�vݚ� |>˺�h��Ff�p�}ˇ�Aj�f�r���e��T����%0�ޡ�+GG� ΋�&�޻mr�0� �`/Vt�놮��4��Y8<�ڇ�t���������b��nd]��tʙ���գae��f�� ,�N+X���CK6I��izˬi=9�]��Dԁ�l��p_l8WnuvFxM��E�\�W��J�r�������8Z������謉���D]�p]�/��2E�u�{��؞�N���oTG;����.�[�X]�#��h�5f��h3K[��p�`88^Wqwhɣц�dй��m�U�V�����4:=�R�M��&J~�$�=���M�T��V����L�y�u�Ho�J3�PF�=�H�>�!���C9o�#�4�l���uw>�cc�WuՉ'HODy%�:a��6q݉��ޮ�nu�}��G=����R5�i��R�
�'Z6���^;V�?�l���C(c�}�[��0����!־��X&w��k�iOZ���j�/�6!��9gTfL"�AVvZ}B�*��'��*�n��*$�X���M�Pt��Qg�9��̗���"���ܸU�}oWR��p�R2n�3gWQ�~�"���IP��mF�WY6z����N�/�5��mZ�[yZP�3�ԦNK��P���{].㻦u:M�[&g<���m�:
Q�9]��G:����u3�!Rs��c��9S�-���C& *�&��͹ڕy�zP֚�/J|RҮa�ښY����s8Nv�j���R�p&zTH�}��5��/��u�S&0��Wo�䲸i��L�2�g=
��N���0&����3�hv�Y9(K�;�*�k
wCiŜ�ҷg�����A�Z��w[�:��h�J�Vʼ�$}&��t5UR�ӽ�3�P`�n��(f�|���t�d�j�T�6���ʋW0��]��D��2��]*z �/8#����f�r��ĺJ�d��ԚE?����o{P���!�/7u(���E(PG�V�i�b��JnJr�V��B��8�]͹E��s^+U2��C��m*N��ۡ{�uV��B�K� ȹ� �s�J}C��z�Ze���Ȼ����oZ�EXN�ĝ�ͪ����s�lL	�fR�2��1��V ޞ��[�.b�$2��Kv�	�3���ќ�#�Z7v��.�a-�y|ճ�Ok��=;+*O�W
�,<wK_sx�_$YI��g�LC&�bmJ���ɽ�r��s�I�ZἈ̚l�#�n�[G����E|�ٻҁ[x��r��;B̸:�4��3i���N�Effk���W�ΉÝ΄gn�����p�Xb��.��û{i�Кi��t\�`��g��=�Gl���(<���.����=c���|gQͬ�]˷��:�r�g2��u�oY��d��m���m��m�e����m�������;�z��4�[�N�k�}�z��H@$$?�B�G�z���߄�v�\�g.y�l[�^Z�(�r�6�^X���ܝ�5����B�rY�K�q
t���X�b:l��t) �h(i�+/��7����R՚��!��u��00F���0v���"U�]_ �]�^-c(l	#KJ��`�ux	K,a��K}��[��!+���JR�+�W�oS����s���4�V��jR�W�1�EۭB�D�T���wb`r]�]:�qEYCx��MԠy�k����Q9ӘKb(rM�1�4Ψ;K�6�Y��u� :�g)�t+(WQnnN�\�ќ$���3�
��*�q�I}6��ep�dއ���j�m4'�/*<�4gX��Lab��ģ���ac��e<S�srVd\(��f�V�e�`>�UҮ���a+�X}��5dw6��2�.�{�3ø�n��������5)v���.���WJ=�	�,�k3����>bNU��X�$6�.�]Z۩Z�aU,^k9�.=�9�Wj	;�$��1k)me1˯��U��;��`����D|�����U����R�Ы
�(��7��J}en[s���5������|�Q�`�5ʇm��S���3`,�wp����mD��B0r�i̮�Zب�#4��v�*�v�0�R��o$6��tEN�{�X5�]Fq�YmG8�g�u1bO�bDfU��;aQ�y�ܥ��j��tK����WX����]�Ù�ۼ�u�n]q�����6�gV�Έ����}��fe�R�N����ɑ`���f�j�U�����rW�I7��iC�+��$�n�N��>Vl�[�p�O	��8[qDڹu�e��v�v�V�\�kO���Ժٻ�tT�\��4DY�Z��e�\ͭS*���Q��3U�V�*��9�Wdk����0+V/�����0��ǽN�� |�]GƆ������y�6%��bƺ9(�m�_+@�2�M�	����8hH
�H�ض:}�ܭ�{���6�{N��T:ti��\�չr#903xd�F��&/;VS��\j����5��HŖ��c�}�wMU�kWӰ��}�x3^�{�8x��n�6q|���+�šB"�^Z��q$�+i��f�<XYK��++C��ڛ�����q�u/�2�}��V�.��eu6��4o����!H:ۉ�7w{v�Vܬ�ʣ��t\�h��G&����ݶ����I���g{����5�p���M����O��X��fm]��-ss�EE ��X
X�`�BܨN�������m�[�3vY� ��È��6k!���%Qޟ�t;�h88�7i�L�܇�qV�f�6���q��[z���*�{v�춺�%g���� z@����n�%��:O��sky��[YW�f�F_Z���T��Dޞ�m���ݖ.̮�y`LVDFc����7M���|Ց�kԜ"�9T�Zg���mR�o�ڭ"��2U��n-�WZ�V:<���,<0������^d�lvMTGJ_v�L�/���pZ��P�n=��"���D7k������S��VM,����5X���E@1�7��boYX�C��|iʷ�l��B��K5��.����]��ŕ�ֆ2,�k�*K����W�C�˻nHM�qrKn������F�.	S���գb�_r�����	t���@r���iἻTp��K��GWN$6�X �F'm�,��W����Cr�G�[[�[�Ky"�_ʛ�
��e�D'0Y4�XTC�2�Ft�&w-�u����F���pK�lc��Ib��e��g;z�R��;��qT.��&��v�X�[��Wi�з�X��d��;-�DH� H��K5#T�	n�9�aۼ��oVc�ai͙Ni�7N������T�gs�f�h�a���ƕ2���]3A�]|E��[s�t��l�PoL�oiS�̉rk�:��\�,�xz�t�m*�m�6�Xb���<LTժ�Gk��u���ݩr�����=/f�.��T�ҭ�����!��Yw]�a������J�2���4�Nd܀�z�;k~Xi�:�!*ĭ��=5 �.����7��<�Yq'��+�E[�U�U��JAuqվ'٬�p��cճ��K)�¡WZ_��8鞮zXX��(��ݥ��J������4���q�o����]%�%%N��Y�*�����i(5�xl� Vk'd��80We��[O�B �)�4�V��$��;ti�j�SDj��W�1ԫ����L�vf�7mJ��-`��i���CPlf�彜�%OC"��v�Фd�)g ur��7(�Ðeݨ��2��a���wQ��G0��ݸ!5���V����dy���Ҹ��G��*k�xl
�t�.�������w
��Ƶ��IS�m�]��L�C\fWw^�5u��z �5R�,�ۗ[�YhR����V��3Z��J�18�L�D��DsQ(��;��7�ecͬݬN˂�p&8���N��n��뀡)�Ͷ��,Ž6`�t�y���S4�m�(S"XH[V+���%-�T�^9��{5I#��)�mkfƨj�qJ���yx����<νȤ�5>�{��5D_nU�<�ɳE]��em�F���k�7���/�Ke�x4h�I7oV2�6�,c;�f��NQ�=;U���49v��\�n��e�]B��Ao eȶ�Qw3_m��C�9�o���u�2��⫐�������Q�ũx�c`\v ��gQ�Ũ�(J��YV���F]�8��L:���i$vݝ�9g`�{���k�Z�$�����Df�3.��y�]u�k�<�j�O��,�= ����+8:WeP��\����P+���<�����`��؊M��nu�堇 鍾+em�fQ��`>�a���nGN�Y e�ݭ���뉕|�0�{��PܤE�]���8��F�v���U�7k����K�p崺%v��H�d	��s�'9MMc���g���/wZ�s����-�N�ߡ=6*֕�- ]��Ui�����-��`=+��6�Dh������{\���ԈF��H��YB�ZB�$�bn��T�y,���I���u�pݬ#�R�����r�)e�2��p�ر�i��w� ��ѝ����BAH�D�*�%��E!dn �K9���Q����ugl ��Q��@�đsp9�IS��,�4VE�⻠��'QwEdu	��J�Xt��r"���Lp��G&hu�ρ������!,��^�c���]+(}֠�jWJ��7Gt���+���
�*KV܃���}Wߌw]g����і�N���uv�ɰ�6��;T	���p��̼BWN����;C���+N�}�f�c{X�s��L��Ӥ�G ��a�r|9��E�Gֵ; l|^���A���1n�jo�8[�v�;��G��̒�jP���s�8"��̭�A%L��\�ݝZ����5 ��&�8o\���#tZ9l�\�y�;M�g9v�qW�e���-[y��]ܹL͋+�u��
�#ij��V�ַj³q[U�i�U�s�)�^�U�;��q�]`�`̵��\](�e��xdM�z���[z�!Bdf��v,Y�!�2km��O���4�X��`S]���ۖ8`Ʈ�]���ɹ���Z��,�dmjJ������@B�'Ќd�]���r�u4�l�ɀ)/s�O� 2ɽz48�@����/��m����o �fI$���F>#5o|ߚ�APv��6��.��4!���kZ8^�"�uPƯm��r��6\�:<Z��L���&�L���C�I���4S�F��$��Ps�6�G�,y{�#�͞w��w����5uد��]���B��BYeT�Y��Ԭ�K��p[���X�Ӗ����/��Ukh��H@:����J�5O9\뒦Z���%��⣩���^3���0&6��ĸ]��v��$�m���ɴX��LF���ܮԖ���;�Ւղ��롩�$#C�t+fl���A�����(���y�����"*��6�5�uN�x�_k��p-q�����h��W<E�ō#G�KO�ܔ��붵�oJܤot�E^9�7�k����ϹQb$��m�y�L���U���'x�叢�p��s{*����y�#��K+���\U�[�yY�%���� ������Z�{2f�:Y��;�����a�֫�4U�j��v�Z���X����$�]Ҥzi�X��U�Yi�Sύ�2����!���E[�U(���#M�<��o0ڋ��1W��W�h��[��kY�:`Z(�D(��B��[����P�������^�mO�((!������s�W�7�e��J���S�5�k����5�{Z�u���P�d��[]ķSt��A��NU�y�i�d_r�
2��Zg�(�_L2Q-�:���	gYj_���e�v��d�j��g���9���*],Z㬖M�q���6t�l���q��;n�����G7(9A�v�F���>����q�&�;JvU�,�鲭Z��
�Q�W&�ݛ��S�6��P��Ν�,3:E��uҬR�N�t+�����ZD����,�+�G��t�s� Ȼ��aN;b]52��v�j[�_A��N��5��b8n�Pn�ʷDHsi���M�
銷+���Ε'lK2�;"��E�o*L4�5��[�w+(�u]�ch�8GN��eة	�����O��#=�W}a���;7�МJ�4���>+�kD]*+#4CJ�!̺Z:�x�Pe�̶�a*c^�zEB2REsW�P\�P�<ÌՊ���̜���bm0n���ҕ0�[c��m��JФj;.n�픷VQ狞��T�-�C۾)Wl�u�`��Q���8�6���ǳ���U*J����+I,ʈ�T���R�t�X�È�b",��!,�َ�<F+G,Bv���s���PR��@�5��G}��/�׽%�n#-�	Y����wc��V�>6N��)u1��2r2�.<� �[N�-�n���ݻ��AL�����G�;���j�� VvN�Cm9p�y�rC8�Wsv9;E-���[�V���t$DwN}G9iј�w ��e@+�|nA��y]W�3�Pr*�:Z��Z����렒�õ���>��XJn6�;[8V:�b��4k�Y��*(��v<�S�V���Ǵ+�f��F�o��.�)u��(�j��v�p	�%��M˛���9��+nb�E�z���=�,�'CI@�e�eu�{�t�7G�i�M��d�v�M�K�1KV�#���X�-+�ݸ���E����;�Y�]O;�c���0PR�k'^���cڼ���֔
�dY��1�)�f�be\v:��ȷ3{o�r��w�U�џo8���#�풷'�u塁h�pɕ�P/7Cz����,�:�)��	�nWm���,�3�z)ݎl,4��-l�{��Jc6&fv�ִ��e[(w ��kT:��qӘ6&�1�(���6ok���ǄĳwWv*�V0*H*���[x��bСyb\���Ź�K����w��1ܡ5[��ح$��OZ����������a��vP�\X�O��;r�Ɔ��K[H"�;Ή�S�o���mf!�G�mu�b�T|����`v%{������mc��z�,L�Ou�C9��ͺ�¢�6��yݤ}ۻ,�e ����c�<tCc��S��޺(j���L�e7Q�Ƴ+��N��3�7�	Yp�r�eq�.[��í��S��eŷV[W;5����09��|�� ��̋GP��CYW�(�<���q�Lbxw
�Iq�L��/�	]�dBwy�O.��ȶ;�[w]�Uw)���XbJ�\��]!-ʫ�qa'ך��y�pt�/��#=\���g�c׍R���S����pu
�R}���'�"��0գp�t�v���Κ�ʖ!9�Lsc�ݻMe�%��t�e�%��Ei�����R��N�R<�Ʊ<G1ؾz%h�����X�[T��*#�h�A�[�]���c!]�%M�DlgS,I��_�P�Po���%C}+#��˫�6�,W}c��gc\�3dh��1.:���>)���R�%�WWV�C{;�|����\����]�;�/D s���J���!��#�Q�n��j=3Jt���5��+S-�[J^�X�巎+c᯹J�3f�w����j��ƪ?���@��ɝ�ݨ��R���2֤JK���F8�|Z5�{�'uɻ��
�-�י��r{CKt���r�D1�/�6TS4j �6�O�ݘڄ�h<jv�i��^rWM�+{�QL�ݘN:J�8g'�Iuk�vp6�Gî������8�*� �Q�9Qs���@��g^_+9�5�J�2����Z�$f�=۵p�+��n�ۍIA4��<+'s��ŤAҷq��ܨpK5Ʒ���wx�ɂ�Ub���Cՠ]6���,��r����p�`K3mK������siAKi�>K9�
�:�F���0���IM�.��+�iJ��*�-U�։�K&�Ҩ���i6k.�O��k*0���GUp��٘��J���Q���q�&���R�׃)�δ���|�k]o&rs�ǥc]� �uR�H� �
��T�՘&P�f|`鸨���EfgK�N\��� ᬧ�s{df��6�Φi�|�fsYa��+G5X�����Z�c(c�9��9�0��*�@�\�;�
'-fSEՇ���ԀSl��k7�	��GH���Nk�P(T�=�����~����p$�	&��s7�y�_X�.��kU�!Y�����A����8˩����O������b8$�]"2��p�iWkHΎ��������1����|���N&�u.�+s^����6.�6}��J]�[E�s� K��S�5�`K���g[��f^d����7 �N�[���*���:n-N�k��-�VJ�gd��ñ	{a���S�����<��ћ��ZF=��;꾵�+/Cs㵱��������17)<��h��L��r:+~KI��2��p��� U���+r��Z����f��Y���]�.Z��m�݊��g��9Z���������t
�7�R�\������n�%S�tn�ʴ�<Uͣ[�\��7�n1�Ӣ��+�p��U�=���[����a�;#����"����H ,i��`���(˭�2^�����j����{�i�f��J����u��()���ʾ1��l�;,(K���	�㣹��N��W)WL�q;Km	[x�ųd1�֦���	|r��|,���uz�}o:��R�+�uvnVF-�K{'i�ڸhzL�S�YKLP!��.���jș��Z��)�E�`�CK��6��XhbQfmS8e�v�vGh���2����؇q=���='mnT��L��l����x�r�s�{6��Z�����o�i��=�5L�Iv�L���}�ݷwx����E��Kj9epj���\���D\j����arʷ̆"�5F�Ze
8�m,j�ڵ�-��X��S)���D���2ȸ�AE�hV�<���#U���6��,Ui\ʦ�4�<��H�DmTJ&d�R�������ڴ��m�.8�|q��m0�51�r��.6��Q�m�-*֍[Dl��U*%�y�yaJ����|��e�I�m����YfQEl,Zո��*c��f�r�x�-[j�o�\(���y��̩Kj)b�s*��e��㖘ƶ��5/���FїQ�V4h����5+�
�.5r֔�*���������e�\Z��֔�3j[-H%��%����m��ci�Q2��\�$j��|��e+�Vg%swG�^-
�p�͠��
=鎝M��T��
LEֲ�TfM������Y���!��9w/��}���놌,~���e�Ǚ�6�&9Q����Y��4p���t��s�H	���]�S�0k�����)O¢N��X��
\���X�: �}y �b-�u�3eI���ջ��>I��ZC��=�����0�b����Tq!P�fVׁ�$q%�Ӎ�tUc �s�ӇV�(X���N����<܌��Q)IV�������},�|�7�稐�X��R�UOZeg�.�,ɞ���Cވq8J�AO	��d�>u�������{ō;�E�v�6�=B�+��ˋ�������G����o���&yV�|󩎱 �pC^��soY�|M;Hnj����ƨ|V��Αް-���<����cO�Oq�c�^�S؝6k݋j`q*�ꎈ�"�,C�P���i�T8,�����ܻ嶅�%4�T�t�v1�z�S��jBu[����[� ���yA�J�{6u�.�/�D>��}�Ƴ����|��C>��/DPVp�L�� Ҝe3,ew�OO{S_h�9��C�׮��[�֩^S�r���jK�f�6���ׂÐex�O5�|��[[�3��<�yNo��A�e[��$��!o0�m�ϫ�ԓ������v�-a �d>��.\%��۬�`�vd��T�$�V��8��q�J�����&t��#��mz����^K�ޣ2͎���c�Ǚ��;�a�L���p��v�?,9������R�+��W�fg���Yh�,$$�&դ+���d3J���}|Vjm���m�k+u��ٗX!�0y�:��V;ZG���5�G�Ö���NOz�3������N./�*ua�Ex#�<u~��	�g�xcQ�#�CE�T""+��uw_���/�Aw����	nj�w"�^G����Ժc�����3�)m����(�:��^��O�w��]�,�fX��Yp�KW�`���3=\���ꐭ5�E+^�n�c�u6O{��u�@B Q���m��}w]����52f�����u��}�$��n4ks�.Y��ֆ���60c�lp�u�Ep�f#�<�.��v���7ґ6�[l���9�eOg��]�30R�����x�J��ލ�N�l�}�
��~~Lps�=����MZ�{��nb��=������A�Rb��^�o����,x̻LV��(���<Ի�fxf��f�:�J��U���]_W�B�\��[����������V�'�������ѕ�'���9fJ�˥�eإrs���B���1�>]x��P��D=�0q]ԙ�=B
��#��͠��4�xL�%!��Sc�>���a�vo/�{y�QM>���A�ʫ_=R����������L�Y�u���$���<����鋬7Ƙ�d/����	�<%v��3麆��å�v����Q��'�y<�Wz��8p�Zw.�U�K�{�ka����LiL;^��OL���]"��svm�n�W���f���),g�/%�Ů�u�0���8s����OV����[պ�[SO�HeoxO`�Y>L8�,�K�I��~`'�� ���=�c�֩y�K��x�e=A���Nf'���i�q���\l�'Y<n��7����vl�+��#U����'��[)T��D����|`�pv�4���Aѡ��K'Eh�;��.�Ff�c�٭��u��"�}iك)t���z�lUQ���ʯ��Լe4P<�v޿�Axl�C�ovm����E	]B
�N��#����u�ښje��f!�s����"~]3=�F������ݶ�bqP:��w��c����c�I�f��D�w�����Q�[��ѣ��4��Է��v(K�p����i�QuG�Sɫ�MhN�]�oAHW}e�׆N�
�BИ5��󂃲h7��Nr�Uټ�����)���p����B����DGV�_!�g�̾��ϯ\����3Z坔�V��[�S������,ޝ���)�;j�뮫=:��|2S�וW�+A�����:c�şd>[�*_{>U�!$�bx5TF��E���N�^9CH�g��ꋫ�~��佰���G�-�$��RW�歯�*��&�}�u�R��ܝ��"�>�_���=��k�/�e�꿤�8g��ML5u{㒃�>��wtW�e�ub��=1�sTϵΤ�oө	<�����#D��J�<>��d���P��|m�g�~���j�@t�{�S���h����>����;�I�<ܚ����A[����;]��^�4}��O��WOOG�aM��A��_��7NzM�<�֫3(�D�r���+q���?fM�z�=J��|y�X58̹�g{�v�d��^�[@��m��p,��Am,�\��
�p�={D\�g�cq�ә��=yI�`WK�z���L�+�Z�s-23cH@���5�B̋����G�oJKFJ�fؐ7���x�L�Ѕ������谞���r��v��nq��*i=�iQ"]v�1�׎�򱫔iǮD��u\��0mF�s.�o^ؾ���E�J����.��!K���c��_�p��������1'��K�I���蟩<ɛ�ᣗ9H�L�sщk��X�Z,
��'��|�7Hy��KSy���r��{��_���o�$����̮N�δ]k��k��=�S��
��u��ދ_F����^f3��E|�%�T�;�w�U�ϗ�t]N�2���do��;��7r�X�ɛ�"��"���F�ꮝu:u`���SvD��իԥ��k���p��q�d^��Q�9WO������T��ױ����V'��j������ur��9̏>�lI]�I�N�T�������˰=%LT{|�_��]7�p�f��v�LR�|ʹ�=�JG޺ͩ��z���쬋D����r��|yS�|\������g�ny���b�`���x�Q�?/E�X�/M3<�'i[�B�W<�Z��6���"|;���x�ݞ�;ћ2�ٍAYE7/��zU�|1ws
��R�6����ۮ���(��ϋfrB1(�R�:�$�.%ccLV]>.�Lx��:�7�:��=��v��}���X���WjN,�7��b�Xḫw���h�o�����kވ=����:�=���&��yx��sʟ����J���N�{�k�����}Z��W�I~ױҞ�w�Ž�����8�-���ǥw�Ɵ�A�����p 3���s�w�l�fɾT��9�J�X�I�z����󽔇,����P� Y��@y��Θ�~�5ë�Q�Y���z'I���[�k��h������<Ĕ�A4U��UYq,V��iҹ_��2�|��?Ro��͆�h�_�d�](���=B��h��Y���c��ժ9����cg�%uF���A�u�u��k��>��g�z�I9�j��kj��
�罳o����';/>���*/���~��ժ�m��Go�����2�\϶O3|yE��>���"��9 gu����g��c+�
�-��v����vc齆^:�~���쏬	/Y�P�*-Xi���Vp���xM�ʇ:e�t0�=���H�ɍ���S���M�?�Zz]�(jx�mc���d���Չ�ڋ	C�&�[�����,�'*C׻,w��7�l���R�έ��s�#7&_]'|�9GϮi}sr���`�����W���^�_��I��,��y�9Z�y9��z�g�n��/�M�g�U��b ��^x����w�ln�p_x�J��Z�z�S�����&��׭�k���4L���񓵮å��8��O{;����W`ކ��}�1�V�ֱnzm�'EzZ�֏���=<���+Թ�Oi\|���F�?o�=B�~�JO=�l��]�:o�.�˳����3"_ֱK]�O}����%����{��i�d�fU�\'�o��o�ۘ���W��H�U��ǀ�l�O���r�a�MzP('6;������K�^�Ŷk��V9|{~�z�:�V�ew�~A����o5&�|������&����$��͛�Y}�m�k�v:OWy�81ſ^Mp�3o��^������,b_�'GQ�@��&7�]u���&�dTo�z��u�ݷ�C%������a'bS�ۙz�.�xO���$ô�HY�n>@��������ZNySf�vWi���ǵ�������C�h���w/�.���o&v���{���c,�.JL����5�HI�(��Ȯ�*�Sr�Ώ��yϞ#�/�W�7^bL����WM�Ϟ�ճ+������[��)��h~��
���Uk<{�G짎{��7��S{/$i�+.�ǔ��n�M�z���R�K�$�V��'�����R��8��N��iu����]q{���*���譎V��>�'j�m�_���3����^��"���J �5TF��ӭ}�����^�a����W"�Ӑ�+V�K;���R����I�GuK]v"߳�7���!�|�(��a�عz�J[_9T����+����T�9�#uK�_����of)���x�{qg*Q�5�l���WR�o-f#)�A�JO��S�ٛ�G�����Ҽy���\�}��:��-�L'�kc�v>�[r�U�ib�>څn����g�37���r
:�ZjS�< K0�/�U0@��M��)V���q��M�MCǲ2�;�ހwh�*���	������k�񶳏Kmߺ�p�u
at۲v����u*�I���ө�/��m��;A �Wt�X.�89P��f�{,gW?����w4�u����$������ʚ����v���XT�����R��p�^���qtw��9|������n�U��^��~��ݥ�b��͹�n� ��2k���;�uN�rN�L��W�Sw�ke�OK����w��*u`V���Җpn���_;�3�c�A�Rc�+ح}��淦˶�`T`��;mu���.n��{=Rl�g>������Yg�y��Gs�8�)�F�~�\ϫkE������n��9��!�ͥ���@]nv�O����%<�ڧ�r���wC�h�Z�#����=�n	�����p�1{�����7��o����T١�@o|i��Kc��x���םӍ��c��1��󰵚�^�/��!v��>�tޕ�,֟������gv|];]^{��Ũ���H�`�=,B�؞��y[��r��g
Ϲ��et�����tXF���Љ]��1E�wnѭ��w}�����i���=�p��R�q[]��1�b����q�9`+���R�L���ٱZ+c���S�n�ӃL�%���Xܫ��ǖ&g	1º��i���F��R�
�������~��ｬ�bJ�ҙ���KY3{����O��^��E󧊏o�yUk-�����#�r�B�^L�{<�z����]�������=�s��G���|��&w������>-=�t�z�x���3���I終:��zr���_�w�e%O]������wn��Ԋ�nj�k؟A�=����k>�u�b�^��m��Dv`�p
N���.���b��MLg��0j�C�[�c��=���H�5KԼ���=&MS�/'�ۿ�t���r�|㸽���	�v�׾\�r�(�}햽;��P�c�V����pn3:�>�tq&3�U�j����ެ�7�L���������}n�ac���W���e:4�#��G�ۏf�4g՘�g���eg�l����Hl�'x��Ԭ�E2Ƴ'���ʡ7~�6�O�l�b�Y�̴
��T�'t����!Y/ ��4�x��Q��ųoS�خLb����J����?b�<��������|M�g4���O'��c��Ueݝ}�]��|s��8;�e;mk%BZV�v�3�V2�����S"�L΋�.�8�^�[�;EmY/_��m�Եc�jqi&T��D�8���״��J|��A��Zlc?Vj�R��
ړ���d���Y�T�Q%��1���R�={����EV5^�k}��y��u^4���&(j���5�7��<&���fu��� f�1��v�XJ�4��ھ����J�1I��k���ج�f����Vw��h�%<��%w���ٻle���uË�ˣ�&3��+ ��2��ln�tq��m�IIs뢂2��כ١e�"�CD9n7�S*������e��	if���lw]�lX��9�s�ks�g+=Qq����i�=�aE��Dn�����_�].{҇lN����)nC��0p�*w�Fh���R�g`V�2n�	�d=\� �%�ں9�� ��{p&5��/�]r�!�4�w�n�X����\��S&�����r��ЧJ1�nE��Ѯ閱N��R3��V�f˝ ʹ���Z��H����kZl������o;����VF��.��py�O,��-E�f���짵��͔�3�	;�Vd��V�'ں�)�m��= �����]O3ǔy��_�����Z�a�/����b���r����$���[�qv�G}_V,�:� �����6�,x���$�W_>������fT��aP�h��n��5�`d��9����#j�롛�n ,B򲷊m��dVcTq����B�P�U�K;ueE�X1ƈ�+Z�r��Z��`�ْWu�_99������w1�z��hN����k��}$"�J�4`�3u/�ԩD�_]���Ԍ�ݡ��%����$D-V�Y�{.����$�����5)^� �Yo룱Y3�*58��v|O.���s�i �Xk�+���/mm4�<>&T7�<��M�x
�D��6���G�Nc��ܴ3���@�$�*T/.G�z}���d�pK�$O��Po��:�n�n��X`����y�I_s��z<;��ڂ�$WE.6�G
�]�][��ąwcf�r�;͚�l�*y�Z��Z�rKl"��j�t�e�Ϻú��ݫ�<M'kvRQ�ݼ�A]��Ʒ��=�#:��`5�j�F�:ji�zV�ڟR[ҥ�taQk�LW0m���Koћ�������R�\c�������r���h�y�M�Zx�-H%{�ROn�7�_(�h�K���Ҳ����y���aYx�Ӹ��m-T��&v�u�\U�a#+C���k���2�I�S	���J����-}������(�h6��iQ�Z�S!�nS)�\h�bV�B�PƥZ[F�,���K��J֩*73�JҖ�S�m�JQ�E\l\Qe�����LF���ʡmHֱ�fc3+X9K�Ln5�5�&R��QK�\��jԥ�.c��*�X�WZ6V�#\f*+is3%��[ke���b\[kLʰ�F�j5m�VԪ���UmZYJ�Kj1-��[V����Zزڢ��-b�YG-��J�-���#F�-�E�TU�Z�X�`ʊQKV��Rҍ��V�j�B�i�lJ��*Q�ҩ`�Z��l�ˎQ-B��[K��iZ�)B��*V�+�+Kjʂ��*+�5��b�2U[V5�֍KV�Z�W)L�F�R�jőD���)kXVQEDjF�1D�-h�)J�mE��آ1������IL����a�3�v��h�vVd����ӗ*'�ɸ��+�f�><ƪ�rVV��;S$j����ݚ�H'.�f�ՅޝMy������<�4��:΃_!��2��;��>�7K:M{�����s��&h��{�f�{�x�x��:�`��B�bI����Vs�{`٫�£��غ���?w������e\w��O4���x^�z�޹�i@�#�U'P~Х;���<�1ge8�E�x�~��<��7�ם�{'��� ���.�U�U���Y�<�SR֤�w{��}�y��{�tpo�MQ\O*��,/e��^&�J���N5U3�_�{װ]j�=��Iz�a}%?#�Xj�*O�&X�z����pn@�nn������W���MS�5o`7�0���ϣ�_��;+�
��b��޿/s����v\�Y�W��� �oө}'�FN�e�,5��A�k͏�w�ŧ>̬��3b���T���z��"ױ�|6=�OE4Rz���m4�{��5���3��6��c�Įuf�^v׎�sZ�F*�j ��OP�c:�vj�a����-�\��N�]*�!;�-�M��:&�6#`蜕�8Uwt�/a,j�w�(�����
��뺤�r����yH�����jk[�W�ӱ _�G�[����k;k2RYϽ)H�9q�]�*��:A7���mQ�j,��Ί#��L��G�v�w���x&�8b�L�������yѱ�A��'f�TI�`X�Υ~s��/ٻ �����1/��3�z��������×�¼��������=�'U���a�4��7� {SV̮�v͐�g�ws�-�PbR��=T�w_;�C���[*/�k�5�j��_1�>��;���#ݞ�no��T�u�:/�渿�����\�rW<�3#�y��楿>Գn|��.�[��P oT
��tk��c�����E����C���,�@|���^�"۹/~a��u,�Bz`�Llp�l��VG��&.�����>�.r�O��$��]E�Xxl�-��;�B�����=�g�-G䯴��0���,�9�dp0�@
㏪���`j)�_I� s�ݶ�9�f�xv�L=N��J.�\��tn�p}o�WV��+��t,̤�Wv_Q�2o1����ר�!�C��^�p�Υ��j�9��b�_V���w@=��{Y����*[W`�$�_�[�G 2���2-��f�����W5��K���}�[���0���C<�Y�N"�O�j��<w&��g��s�rҼyS/|_z^��s��@üV&�C��w�w=e�^چ�mB�Gm��g�~���
�X�ڠ�CT���}��{��Ϻ�W���ͼ^�P~4
��r���3I��n����o�z�R�I+�4�2�ät������Ǖ������'&�T<�#��ә�x����v�X5t��������#�}S'��~μ��s���r΃j�"�2R�>�R�����g��r?/Q[��X)�K�J�}}�5���J6"�A���N�)�ΘbOz	�I��qz�����[�u������;���o�A�u�֋���'����u�Ǽק$������U�L�f�d�4�;��0�5^>����w�^���g�e`U��V��`�8lY�!�2�o�;LK�v�e�_S�_>r�6w($K0�	R�����Y�A�1�w\Ҵ�y}����ڽ��nR��v�%��4�I4���X�;�v����K���{ݽy�ْ��\�w@�η�s��v6gynZ��Ӿ/�J.�N�(�����=�	���� �;���U�}�w���	T��s�^Ļ��O�eo�3T�u;Z�^�E��D��
��.g�����K{+��ۂ?�Yُ����W���{]x���1���:zF����C������6���G��O������a�߰�~d��y8�bu��;��I8��<d���{�^|�o^�k������;
��6����	�6ɣ���I����T�'_�O�`T�d�'��~P�25C��M2|��w�m�d���g&%a���s�;����cI�����]|���n�|�Q���Uw�Q��d*d�+��=d�9�<d�a���%2Nky"����(q�i���Xi��������O�8������\���?~׿�~�;�{����O�?!�۶l*����LO'=ì� �4w���M����0�I�'��^�$�&���W�$��E&�Y:�2é'��~�z���}斻z�e�{��巹6���u|>��c�}�'�8����M2u��a&�������CS�ì�J��~I�OYP�lY=d���I���!댛d�o|�Wo��oޒ+�芝_�������X!�	����CI8����<d��u�m�u�7�$�������I�~9�:�ĨMN��@�&�I�?d�m����X��k��eӾP t�vŁ�d6$���Y�ӯ�k��������V�r�Ml:)!�Zǎ�urO̬~jl�="e׍�˭oR6��y���G>̤���ǒ���\�|cO�u�����]������ǆv�u��u�0��ɋz��R������ng;};B�����6Ԟ2m52�zβi+8�=J�MP�N!<�ء�'Y5��hq��Y�z��I�59�N��'��i���������G~���?�T߿4�?�/�ɿi>Փ����<�+&�$��1'�P����MgO�T�j�Y&�0:��O�R)8�����'�?Wò~�����鿫���_�a�ﲾ��2q���{�8�o̞���u$��3Y%a�!�hm��l8���z�2q*VI�:��C�,'ɯ�q��_���i�0��'3���V'�9���g���'�T�rAd�v�~I:��fN���'̞��d��l��y'N'��IR|��Zed��hu��邲���u^��Q�b��߂G{��e/xv'��Os�6�����~@�'wC��$N���p��	�4}܁�䟙?{�!>f�5�~��|��%I�A��uB���U���[3��[d��?���r/���2m;��~I�y5a�x�:�ϰ:���C�y��������}�I<�3o̟�<d�5���?$��i'�O����B���_�4��ş��O�c��dݓ��%ABw�>B�q����I�Q$�'S��I�p��2u�!�^`~d�O_��9���a9���M0���k�N�L�a����s������k�o��M'̝���|�����3w�+'R�x@�'|�0�d�{��$�<5�C�퓬?}�:�6��ܚd����E��e�̖5`K������wԯﶓ��o	�4ɶ,��p'P��]��8�<�T�&�N0��%d�8��O������O'�Z�|��[�
��L0�p�y���x��y���L�}3�0��0��4��I��p�=@���*2z��w�!�6ɣ���IԜՒ�I?n�d����,�d�'|���C�W�~��׍~�?��+0E��	Z�m�|�Խة�����od:��+�W19�t��٢chb�r&M__^S��58�5�n_Wp�Q��&[���s�F��@|V0�]��>K%o\�C�7)4�stfWg�1vk;���V=�W����|�Sg暴	���2LJ����u�XOG;�I8�����*d��;�!Rz�Ú��IĚ��IY'�Y:�@���L���ÿ�{�u��|��NɦLI����̜d<՚}d���=� m�d���u�bVsxu�c���ԜAHw�~I�OR��)
��N�'�'Y7�����on�z��[�������{�+�I���dX~z���Xq�~}MC���8�y��z�d���=7� m�d�����C�9�:��16s�:��VC]��8ɴ�5��ӽ������� ��������{Һa6���~}I�h�a6Φ��0�	����:����>CL�A��xI�a���SL�h{��s������ߎy��ݽ=d�VC�{���m�O�`m�l�}��	�G�����N%a6�'���8�=J�a�a=��CĜA@�sϾ�U�����ZѴ��o��h�t�o��}���O{	��C���z�$������Nn�~���'Y>v�ӿ��6�o���+'�����Èze���2u+8ϾwB��z��ﶌi�M��HW�f���(z�h(݂�l�J·���I�4��L'X}i�O��'��u�6���o�:�6�����~`x}CiY<I�k,��񓉬��~_��;�:k>ϵ��s��{�I���
I��qC��%`h��a�N%f��a�y�rw�$�Zu����K$��'���q��?f�J��C��߻��_�q��Z�[�߽;�׼:J��N3�)P񓩣)�'�4yC��$�џd8�Ĭ{�"ì�}C��rAd�k�;�	��v���M2}��u�Ng>y�x�~<�5��ӿw��w�VI�t���+�Z|¤�Hm2q*V�LC�bI��d:��l��d�'_�|M�$N���so̜d�'w�f���'ﻧ����*Y�9H���Zrjr�
�[�m���)�B^Dֹ�a�ْ���&l��H����'�V"��{l��t��"��v���Xv�|��4�K���{$�JvgO�X6P�V1ot|���f���qz���������s��<�@ӦOXx��7��3L����!Y'�̲T'���!Rm"��N2u=��>I��3N2�C�N����=@	_�__�}��ù�;<�,�ORO]�d�'�<哉�&�x�]�O��Nyb�8�<�T'��
�Ԭ�2��2|�a8�����8�Vs������F^���T�糧����z����?L�d��m�y�4�����M2m'���:����qC��*T�oVO��~2���|��5��g�#����G5�݋�~}���C���d�>�5�!_Y4���N�N=C��I:�9��2|�����<I�5��N��MN�a:��RVV�wO�����{��gu�?s9o㿒VO?X�O�>d��c	�O�����Y:��=���̞0����&2����:ì��i��AHo��T>I�5;�!Rz����y��Otw��o�������󧬓�Mj������"����I������P�'5CO��d��`z�d����I1�o'X�LO�N�q!�Nk�ߞ{|��s�}��}��gaP�ɴ�t�!Xz�����G߲K��;�"��r��I��k�4��C�_���d�É=�쁴�'X~�3�'�T3�{��q�w�y��������˯�޼����bt��Y>J�����N2m+�y�+Y<�Y�$�'ڲ]XN3����&�A�d�����$�	���=M2u�l����\��}�>������a�OP^��z��}�u�����N��+!����'̛ݓ�� ���Mk6�:ɯa=q�l�O�B~}d�h�8�=eM���u���w���}����{���6�~�8�2m��� �I��`N$����'���ru'Yw�:��&ݤ�9� ��m���VOX������󏎽�V<���ϲ���t�狂Mۅ�eb�e�S�YM�9#���F�^^3B�����L�u�4��g)%�<��߿au}[1�gn��]���{ޫ�\fp�]�r�uӈ�M>��8�|�)��EScn�P8�o]�9�Dm��t�#�tz�����hq������(]}��E��I�*i��Y&l��N��}?}�m2u*~޲�:�G<é��>�u�������N�|�'ud�$���s�~���R�ܟ?ݲ�k����J��@�J���YS>g�gO���jè)'�(q��R�� ��'��XN0��y�_�'X~�a�N{a>��{_�~�M~�c�t�'������|�￼��������5��>Hyl6��l:���>a�N3F\d�C������:�É8��߼�):��h~{�'Xs~��zF���cߧ���:���쯇��Υ}�I��$�������VI�5�2J�䇖�iY6����C�8���Og�O'Ό�!Ĝe`k=�����׆�Z�>k?~��:��S�����}~����8���m����2~�p�2~I�;�XN&�7�a*I�7�2Jń��q
ɴZChq��FI�3�ۿg>�?�߲ny�����AW��_~�_�W�o�!������O�P��2�Os�$���'�s	�|������2��&��%a8�2�PP�O���J�����y��+Ł�>�7	���UK�����}�m�5C�O��_d>d�����O��?�4����)ש4���w$�i�l<O���Xi&��d�C�>���s�<��߾�����k�T'O.�T�eI�@�'Y9�4XN2m�~�ֲN'��C�퓨~�s'RM�a�3�i�Y'?ܞ2|���{�u4ɴ|kx��ʅe��u�f�����t>��`,&�y�d�*I��*O�Y?e'6���N m=����'Y8����B�2i�'LN��i��I8�����
?�Dg����w�+��]������d��>��d���u��?d�+	��E��X���&�=|u�	�!��x�I�O�~;�l�'�9柆7߭f�����5v�G]�x�z#z��Q��R�jO8�Y����I��tQ�e��L�X�1U���zrI�U�����w3�-��tøl��3h�Fpl�ڄ�][��+����C���i,y��(����:�N�_!m��n*�az���U���}��#�{M<��2LJ��7�=I���;��8����r2z����T��xsXx�8�_~�+��svE���=�C��O���7�޿���]����qc?�EHQ�v�䟒{�����;��a>aP�>è,��{�Y>A`h�p=IěeC�y�*OY<�^�$�'ڲWL�������[���t��yX��K?n��9�"�v��v�!���~��i��:����M2q��a&�������C\�d�T&���ԟ$�*�� K��|a�u�߮���������e{��'�vq��O��XO�Y4���OS��~���By5�f�8��,�C��Ay�a'�u����$�?sxu��n���矮��_�H+�545_��ߒ��?�O��s����';�Y���i=jO6�2�z�2i+:�=J�uC�8���ء�'Y4~�$�d�V~ް'u�'SL��}�{��?^k��g��0�W����~�[�v��&��N�xu���n����:�=u�d��L�O��Ĝf��'��'R��'�*{�Ad�l��N��{��"��8ʜ���]���{����Vv&|R�|��^~���|o���ܮ���\;i�N?�O��d�M�2z��u$���d��̇���Y6Èh�!�x����c$�MP�	�k��r���5�N_�s}��|���zɴ�����I�*k�rAd�>�~I:��3'X|��OM��'��5���N0�O�k$�>Hyhm��lRx��d�_�r6�Z��U(���vz��������#��<d�u���'�4{��d��{�����;a1&��@��O̟�xd'��&���B�O��d�>Hs�o��d�7�&ez�_W�����B����2q(�=I�v��<d�:3��q��yCL�d���@�I湛~d���'�`~I�'�{I8�2~��w�s��:�b
��7J��;����4���;t�o�|�6�c����E%]�Å��K��o.��Ļ�����T��������(W�~�ni����f��9��mh@���V�t2R��}����s��6ewmi8��y-Kl��N�-��ϫo��g;���>�ޛ��oo��VL?��a*
'l��h,<-�:��Q$�'S�V[$�<5�̝v�~/0?2q'��{���M���s������U4��AXϊ��J��ԞA�����:O��O�x�^�'ɦN�Ad�C�RT&�x��u+%@�'|�p��d�y5a֤�g��!�v��X�_}�T�U�s��f\����}���~^�2z�{���i'�����4ɶ,�НC�'|��N!�k$�XL�8²|��ɔ�@�'�SD��q�h�~F�:��W��&�L���rnz����Wi4á��8�c>a�����Y'�8����!P��k����M�2N����%J�d��
��� ���_�K���)wt��l~eP�c]9G����b�����L�C��rB�I��y�I�Xx}�:ì'����N �7;܅C����]��=I�,ē�?}������ҿsᒢ���!��}Q�z��~d��fY8��O���Ì�d4�Y<aԞ��@�4��7��$Ĭ>���$�����N �5���'6������4>�$�uPF{�g9��l�}K��������I_�'λdX~}d�k,:�?>��2q��k��Y?$�M��f�8��o�I�:�G>è,��m���΁���N����_���{�O>��gC�6��V���m�SzߒO�=Ւ�a:��XOϩ4�L��l�k���q����m4�ԝI����4����v!��@~����p^>�;���s������q�xq��Y��d۴�v��&�>�k~Bz�״����N&���z�L��$�*zjì8�k��q���E��5�׽��߷�{���>d����'R|�2�g�'�=��u������:��O���w�@�&�m���%d��i=k'�8��YY�'SYg'�S�m�Lןg:��xtsϽ2�.�y�/�o�عB�'�5�^ẽ!Q�4eHQ��JnU⃅�Tӂq�L�i@�y� �À��S��lİR�;ś�TF��&wq���h�ԥ���e�쭶� Ek�&���Sŷq�}CEqy����x����T$`Jo�*�V���h��V���u�c]Xh��Z���8bѷ�fɲ�An�,���0+a���̛o#��L�9��݋u�{ov�i^gP9C �Ȩ���c��8c�K+g[���v�����$�wQ�pz���Bs��G!���ͫ�o/j�K�rUm����kv�=��*�ҡ�_g��^J�cL���L�X-�Bˉ�k���|����.���Ɂ�0,����.��&)�W��˵Hǰ���2�e���]�,{`}\B�Fɱ��^2�u]�����k&L��w*�4"�/��V�OM�j���]k�#mq�	!�d�-�:d)ٮ�I���@�u���䗼��WD���J�U֬�}zܜ�I�z�{p�F��`	��f�ǳ�� ��������?�$�6d�]��m�����%���Z�w��: �I:B�P��
�J7�l���riǦvwhn��R܂����V+]:�Z���φF��s8�.�N���� d����B�U�����/^��Ow:��I�bĄË���%	����S�]�hؙ�hpv֞{��pV(�`�VK݋^�2.�+wf�d���K�޺����l�N�TtJo@�.�p:���m�V�)ʐ_f�/+_S��}n�O���ͬx����U��+�c=�Pꜰ�6�mnԌ���p] �yI�֍kQ7;A�V�ރ��s����P��qr�@��[۷�!�@U�O��wuo�dچ�b��(i����N�}o�_��p���4�Ɲ�:�,��]�۳-���`y�1g:'�:Y%�O���%�;zT�;!J�����R�Pr�۾g#�ګU!�[��J�.��}�$دL��������s�{HN�Ƽ��oSF�e4H?d���z�Ev����j�Wz�s`�@���^Nպz��HX}�n,:�<6�e;ᓄ�^�<�����ab7l��ۭr]�Q>��
�)��C����W��s/2u�)Y��i�봫���a\~�gn�\�;�ә6A�Ky&��M
yoD�\�,�y�>����;Z6�WAgۛ��l}�3����*%)ھn��xݎ�`k��$�-���=G�{q���D\�P�[aRHl�sTq�:��x�L�[�\���b���z��}nK.���]BN�k�*�.��[��ͱk�㻔��ev����4 ���Y�[֪���MX�JJ�R�kJV�+)B��hUǫqh�B5u��>�YWKv��V�r�� �3WXX)E��t�v���B���;�νt'�2s�J�t�(��o�⦳��m�������1@~4+�$��1
6��5��0��J���VV�kZ5T�m-VVF�-)J"*T���b*�miF��h�j6��F�����eW-ĵ�5,�TcV��R���ʈ�-�*��n5UTDD�ڕ
��ih��Z��A���%ke�31��[[Dbʶʥ�����h�l��"5�ʔ�EYm���Z�Ԩ��Q�mZ��m����*�1T���-��UkYX�[le�`�Q���U����b�m��DTEEb���m�Ұ�T�
�qj�
�X�R��\K�Ƞ��(˙���R��`Ĉ�.5E��)���0QEJ�,�Z��Z�EF
f�j�TbZ����T��eU�TQ���R�Veedm(�*�1-b*�Q�Aq�j��ƭY)mJ5�+(�dU-(�DE���-R� �������Q\h,U+TE\�rт�+�hBaj5��:�s˶�{�3��-���ۣεu�4�0�qD�e�@b���Q���T6��e����vp����}��	�'>���`��.��$וC䞠�'���d�Vj�q'P��0�4�u���|��~9��Xm����ߒu�m�Y+&�!�����O���<;Ϝ5��u��~��ߎ�c1���'�6�Ch)'���C�N�`k��E�8���H(Cw'~�N��Y8�a>���'�Ԛ�y'NW��������Lſ�_.��5�����?%d�N��6�2q=�bI�8�yC��$��ϲd�V�y�Xu���~�� �uv���bM�w~<��c������~��������Ї�Hl�D�B����)���$I~<�}�OHy���2S�j�p�����s�ѝn��xS��?�sΖ<�����ZM���)��b�ݩ�yx�/>S���T� ��t��J��_s�㖳z��}��3�����^τ�m�R)a�檏����Kñ��9�י�j��m�:kk��ls>1G�T��IW���TB�<�-�"�����L��J�+��j�n{������G���%ve�w�1%��y��l���5�+Ȫ����a�ռ~Q��s��l�����%9D�l��{ʇG��*ݬ�����P�{:����<�-&��s2��C��;��r['��=a�w[����m7Z){���>ᇗ�b��}�ͬ~Y�0%7��E�*;[���;��i�[�]�	����z�h��ƴ���]:Ao&5���W�UT��^�3����U%q\�����CX����N�zc�ۚ�],�j	/'~�*�f�.�4���y�GY�yz/�+��E�X�Y�	��o�$��:Z�[2R�ޞ�>~�J6�ޓf�oȣ�����d�vǺ�R��˨m���^�����t����w�7w y^�پ6Վ ��fn���R	��7����_�r���qLgy�7ޚv��T{���W-��F�
N	��<«�[]�w��r�|�n����;]�Yў��
����\_�؅�ֹ��e��u������=}ݳt�`��0C?l�m�l���A����CgY/��M~�v^��Եt^�T�aW�H��?W��7���of	��ٕ�t:�V��ۮ_�����'lķ���s�/���\z%O�}��ý������_/�.��jD,��$���s=��IT��؂�#�:����|�F*��/��򛭧hf}�-�|n���	��#M�h�_Gd�g4wpc"u7rit�q��˧pk2�z�PdވT�`��W�#�ڎe�/,��;o��uh��m��;�w���G�X�c����磌���Q����@�����k�Z�Χk�\��E���/A2$��n^s�}�iKT��X2u�oo%;[�f9�@��3�ףr��l׌K3v川��C�����6�)n��f�s8�����Pr=�z�3�3�ӷ��~�渜'�Z�[:⭒j\O*���^���
�wa*��
�{����w�{��=�i�w�&���G^�մ;+�2�-g�D}iX����m�OS�{=��V���9E}ގ�Os�^�X�zm�KN�'�����o��ȩ�����&��njc_��=��	�v�=�8c܄w���v��21i���!m�y�w��GW��N����mIZZ㙋M�C�E�����׵��+�Z�x�Q�.���g�S��V>wF��G��w=O�����F���j�^䗝hyb���%_�gI��>l�Z,9]c7��ֆ�O�Z���M�<����n��4\���o��C+1^ƒ�k`��[�A �]�0�]�6���53�h&��vC�4iQS���VSǹ/���vk���S.v�͡�F�0K._E���s)�Za��q��Wn;�:~���ꪪ��{e�]�������t�c�F����W]mk@��'g�鍒;�Z��8��;X!@3נr��_I�3�xl���~=ח�t��v#������\6 O���t��M��%��iC��g��C^W{Bn]&�RM�Z��¢6�����=��9�}��Oy]����C.,c���l��d��]���C��7:mP�쭗����j����j�X�0�b�jt������跖�)�|���Y����R����~�n��ֲC����s >Y�Q�g�E�.O!n����.u���<�v�}⏳�������Yx���#��*�$����ʢ5�el�1�j��{vM��Y�+˗���}�M!�f�s��&$��@�k;s�#`ƛ�]�7���pd�����qx�w�߻T��j�{���1������͙.zw����f��y���X��al�˱p�]ͳ���w�e���v�]�T�R��W{�ѧ��ҥ��|��ZF����x{W>p�Q������k^�')�s{s!U�8m쩬������E����i���eg3���|�| �N�W��]w�&����*o���ZW�&^�|�����c��w�f�t�r遻�I�3�v�h�V>^��Mvܜ79@%�!�p��$
��5��j�[�'��|:w 9o����;/�aG6��J�M���n��=�x{F�w58������d쿽32zUWap���x��y�b�4�{{)-�<j�n��%y���S �G��8���y{Whڞc���Wr΃j�"�ĸ`:����'IӃ3��zVx�����b�7,=|���FĿ�V�z���j����<ĞϽ��ӷ^Ჴ��M��޺���ė�z��뇫~��Y/�4Ý�;:z�P���G�m{�ݷ=kV�o^)���F�̮N�δX�q9�˭���qE=�/q��s���
>��j/����ӎ��yx��A�j��J�>�T�ee���g3uz�´QV�I��X-U��:�b��W�pn����7���.+����F��E�$���ם�G��K�j������ܹ�r�t�
^�}�Q�ˍunTPq�h;��9����շ@c�������4:osjy���y���_}_Wý���S���j�n��v�tZ�-f���~�m�
D�݁ۭ��D������J1�t��඼���R��GG�hy�u;զs��v��ed��'	a�&����I�{����V9��T�=�Wj���d�� ��-y�{ ��+�v;���Sv�U��ކ�-�*��t�����X��ΞV�^��.�ǣ���������@�����N.�k�	Mߺz�/Kry�du�^���ƻ<���`�|��>5�]�kw��Z��`�E�W\W� |���Z]^���Ԋ�^y.��}������꿗;�A�[ ϵ9��UT����/y�\[}��&e���{�K�<�.�^���@�U��7�0����N3.hgz��>z��^��ǣ{����O 7J��[����&�r��u��$3��~w�Hz����T�+�3 �r�uR��ž�s_1�쩙f���%@Z�@Qe�:���ٹ�]eN�N�0@�T,a��0�.�N����ձ��6k;.�$���M�H��VF@�x�R�����0�}Մv������%��Z��}��}��rJ�ޭK��?g��!&9W\6����N���˛����/	�I�]b���<��5rl�1�����̮N�V֋����%��~^��i]�s��{��.�;izc��E7��
of} z�ٕ�;�y����{���y���׫���Ff̚'r5|z$���ot���'t�L���0�{��K�P���V��GK]N��v�/��3|�O1�~�]��U.m�f&��K�Þ�;\��;
��].��A���vc�"�[�v.���j��y�,ޝ��3b���?olG�k'w�a�d���«7����zzM�7ٽ�T�Wx)&���X;/��֯�Z�Y*�o�[9w����@��wof�5�c��a%?R�:��մ;+�1���X���E�J�1�bw��y=��`ޝK��?Nc������OS�����˽un�V�>V�����At���,�><u��7��)�w���Xv�p|��b��N�7�ۜ�VYV�&��C��r���\F��'���HU�q�:��]���n'1�����-���b����|��[7��9���|�5��o����u�?b���?njc ױ>�S��O{���&#�7�����>��&׳�{�$�C�ژ�쁍^����x�,�ۣ��f�V��M�����{����� _��Q��l!��T�)�Q�]�����@���/W��{�l�}���B����=G�__|�����A�/�v��:�hZ=�<�ft��~4����^g�2���C���)s�����O2���O�n����A/39��I�?��ۖ'Z;�=�VD^u���7.+���֏<�v�S���a]Q4���;y�.�_9щk�r��Wբ�[���.�@�~�O���Oy[^�q{G��c&�[��wkWw�>�wl��C�h������v����u��Sl��{���s��Z����)�9;�P#]J�}���S�v�r���o�>���.]ִ��ta�����,�V���� ��^�Ǯ�Z�T{+�����q����꺞�}��%�sV.	F$9��F��#�	J�Q�c9�u^��_d�@�%Jc�.J�M�Wv��Tw����ս��>���|>L�t��n@�������V��/�E�jO\��@oMBxu��:e��7�����^��jW��{ajL�*[��pI=W����:��o-5n�����}�e^@{��p�����k����rS�Q׽9u�2L��7�}���^�3+6���$K��Tφ�5o`7�H��6ˮ���~Z=�8��f��=mk�'�VT�:=-�'/ӱ�uJ|�iz���5KQ�s��:hx����?y�[�V5�g�=����R{�#i�.~�-w��=:E��K識�}N6������� jB;��c��sv$�Ӫ�{�S���N3/=�6|��׋l׍��p׾�ԙa���E�s��Vz89Hy�̹�7��7���{_�'/!u�-�6�k
�YW��	օ�~�R���:N��~�s��q�mh	�}�yë��h��RU��m��L�3��w�
�Ӽwi��TP{ʎW	����D]I����l�����g;ήK]N3�8���93�C��:��J)Jeb}xD�nZ� (Բ,�o&3/�21�S������K�>���;d.w������]m�^�r;|�:��\�o��ނ\�y|����#��tt��s/}I>k�䥍���W���5��9�,
�.u�^�^���0����õ7��
ofH�}��B�ᴇEF��xjq���^�����g�~XT�.�.�~�'k��9���✓N�T�Jz����[:�[�8�9	���]?}��ʧ���;�>�G�H��)� ��Ō�@��#�Y��ϣ6���|�9Z�U���Oot�.vd^�5�o���oo33R�K�a��_K �����՗��a�U�>��Ӓ�����jny���U�J⭞Y]���v4L�^���'�{vgF�Ng��s�jgc,׽�IOԾ��a���R�����/�y,PÇ�w�눩��&|��_z_OP|�=���{�b�������_'S�Q�^��=����\����f�|�Wu���ʠɝ7ћ�A�0>�=�+���m��e�ಚ׬p{ۨD�Ky҅�N�;]YȻ�kh���?r:U;�{h9[A�8�5��*��]/Sع��`E�J��.�+9�rƉݽ�}�T�,>bl ��&��EQ�������w��m����J�N-K�.1��F�3x%d��������۹�0�7h7�-�N�i)Z����+���߻�tOs��>�3:�匶diLM�0j�crh�Y��حt���q�|:�1��E:s��|.��T�!ބ�U��t�m|w�%� �������^2�&�6�oR���9K�U�k�=�V�Ӥ�ͦw{�;�?�2j�BnH�ǫ�N��Ewa�C"�h��t'���h'5��.m�i��ۼ�A�|��.A�g�t�cs�ol��6������؝�;2լa�Z�!���|�X��s�]ǲn�K�F	��n�^�[ ��S���;vɕv�y�aY3t� �B�>e��\B ��������rp]�(�Q���"K�o7շC�o���_ ���-$�\.:��Z$�r�&�b-j�����p�_h\�E��)�L5��{G��ے�x���Y�gs&X��5��j���2��K�yZ��B��lK�]�6�捺T\���a��к*�	�8� w��Sfr��a7��/R�شK�-��>i����l��6��O�e�Q�U������lrD�/�0p�o�������m[y�׻�w+��H�M��mne5}��EB*$r���,ڋ�R�a��sKcw�"�*�'T=3/x���˦OS�w;&KUf]��aFJnV��Y�g`�hJ�/w�]��i�]chj�u�rG���:�e����f� �!��c���Ǔ��B�د�p�}�v��Xh"�hI�z�oKv���i�ɻ_�ܠ�m]�/�*w|��.���d��0Jؓ�m��v!(�sN�2�5�)k%�,y�P���#2+]��Ec�k��M�],�,�dY�.��|�ָ/�n,$�g��!�]ři.=WH�ǯ��ϴu��w`s*N��k�����q�Ш�L7,<�1ԏx��/ijD��wN��kWtn���yJ��u�?vH�]e=&�.�r�R�v�f��l��f�c�J ����|.�y��U^:^*c�<�⇸3F�`�Xn45�cS�΀vf�ùf����w�
ʰ9�7e�"���_l,�s9Q�E5�B�>���3�%l�;�ޓ.�����qK^Ո��Е��s@||�.<K���yu#(Ry���Gcԡ��`�ިnR	=eK���eayb�]e���i6��ٗ)�pR�VY�͈9h�lm3�o�t�U�w���Lf�B���۩ؘL���d,7�j[]r�)D�q*��;�p�.�ݻ��"��*	me�,b�A�"���Z�V�(µ+V%eE���[mkm���DUjX���"��+F""Q��X�
"�`��*Q����TRڨ����QڱT�QĪ.P�Z(�����DE�J"�*A`���j����W-r؂��V�U�E�ZĈ�UbDTS2��
�-R�"�)S&\Tb*�"�+Tb��F(*�1A�j(��UE�X*�\X��iUX�1DX%�F1J�QPV"[QjڰV
-*�Z��EAFڑ`�1EVF)ki"��Y�UTq�mBڌj�m*�eU������XbD(�D2�DD�,Vڌ�J
���30DUH��E-
#j�EQAQ����Kj��*��**��UUiKZ"+m��kV�UH��1�Z"�¥�X�%����Q����D�,��,Dcb(���QT�ʋT�1R،�R�B�X��(řK�U[e*���#aQE�ؕ��-�F,U���E+Q1��ZX[ATE����p�ݺ��W���j8�7���Ցu:C�4�s��6��K*�	�(�SsK�)�˗ZuL���N�w��������?w�s�R��NN�������j{Og{~�u���|=A���>�{[\���7��Hv�����Vm�"�S���I�r��%xX^��m^6�ۃfe{��U=^L����)���e�Ǐ��ѦiT�R���}e.�y�����n��.�ˈ����������4Sgۏ��f���)�iA��d3�����L�u�����R���f`@��n#�佋��QT��y�=���}zl�@5]u���c�,S�7w�a����^ǧ=��ct��$�l��Ps{0H��\�\���>Wޏ����+=�uح��]�=�{i�e�OQm��HX�_��o����H���T����S��tܦ�|zb�&ibGI�G�3���;��ռia�TN�1�Qs���)��\�#���x�l�X�h�w.%��R�0�RәÈ��3R*��-,�	��k��.��z"����8�YX���>@һY�t.��g�=Y���gu�h���ّ';���We*<t��=��RWV\}�3�UL��e����zocF����]k���}���S����K~h��Y���h�rz�]�>cB.Eu��U���W��F���r{���[�g��}R��J�$���kU�贙�f˜�����ȯ���^�k�����u��hv�ӷ�ݞ䕏Z������B�n%�2{{���,=���8)<��G^�;�:�,���7�~�ݛ3gR���A��>3<�X�����k��~�K��;����nnl�o9~�o^��������غ��S>���If��>��]=Ο.�T�G޽���{]�o�^v��`�j��<��k&�����tO-�ɽEnMS����{6M�.�uXf����{$��3^{��׷`"}�=��^n'r/��#~�3�p]����6Wgg�]���O���z�J_g�bt�;�c���$������W���2��gf1���d�Gq�`j��b����I����E���N���Y[,�q����3���o��rȉ���{�q���g�b�?��lN�2_ ��[w]ۘ{4�k�;i���K��5%%uTc���OCv�����Y�y�����#���qv�����u��:���7K�Og�E�ɦ��x�>6������1��7z����K����m;������I����}�}C�\��]��ժqYӮ�`�*�X�!�Y��V��K���L�i�ʛO�K����uJN�ϔ�h;j��D�w�:u����*o��qj���������;>����Ƚ�y�*�pѹj�t���l�7q��5�������my/���"�*_#�^*�{�k��0�R��I���َ	���T�S��e*<��D���W�D����rj+g��������W�L�z"��=��囒pކ���`JfWy���%�Npn?NGީ���.���?�	����E�N_��L~��Ax۳��a{y��=K����˥�{˝��z�ݕ��$\�����Qm=�%A6]�+������S�ʞK�� v'��SAהEns�Zܮ×���@mckShK"`�w���s��s���]o|�j	�gnW^�J"��������*r�_�����7u�&���Ԣ��Pt���U��Pm�ا�{���o�Ƙ����S��	�U�I�Md���~��B��\}\�4��sR�A��˶��l��w5;���#8��l�CX��|y'�dW)I]���oDa�)7��T�~�k��8�v �}$x�X���9�y�u����׮����N|��bnغ�L����t�KV@�g��}W[b�^����	־:�7K�$���{v�3��»�9�D��y��]^o�q��s>�@ףD�!r���=�_�u�l��;`�����6��S{0H�b�ߝ�#�h�q�5���;XTǞݓ-oy��>�~_�S�����sW�H��u��;j���o
&�<���k�Q�z�9{Qn�o��;>�Z��I��g�q,�ƻW��Jy�[�x�Tc�Vd�B��J"�Y=�ʖ�
��ՁDb��~Ub�Fbͻ����e���k'&H��7�sQ�O�a�������;w��e���b@;O
�mL��f87_K����g;2Ưfuu+(̭��; 2�w<X��S7�8�}d���j�li��;�IM��S5;F���ꪯ���v\�sϭ-��������`���sëܥ�*�@�}��v�Gv�}�� �^�9�xI��ݴ;*����_ٺw�+���8�r�(�"Vt>N��U9:�A�8yu�A<�T��E޿=r���t��0�+9��垔����xp��t&^;�CsT����'���v��ӡq��ʞ�`b�����R�nd����AX6^�C�n=���6���4�v�Q%Fsv��<�9�]��U��ke��D��1aqWx�����P�}�GD\�mr^�ט�׳��I�Aև�d���AZ<`w[r���߂yKèK8;����{D��կ�_]�0��Kg٭��mo��"��w^�=r��k)��(Y�!�4�(�ԣ��}[ajPӊ����]���p��q�8�Xz'㾩7 ~�Ydp�,&&$� ֊�+�ZĎ����j��>�k,*\|N3\\�UR�M2��l�I���4��K<o:�����F�|:S���m��c��{�Y�+NP�z�0pr�K���_@4���o�9��ԷH]|@�7�5G�/�Z��oi��[�9D(^�bx�!4uIݴaS��G[��Y�y6�k31mM�ٷ��i���Px�Vō^����>W�_��M���*�^��$��HT:�k��|˨VF��Cx���>ٔ�j�I�H#�swn��a#Qu��
;Q��]E�*@���0�.�z)�Հ��+�{e�
�H�$}��>��l�&�uĈ�x�H��x,[���7�:X����Ժ<Ԯ���#���;O��ۋ�}3d�����
�j�B���	�E����&�I�kv��T1�p/+���K\�]o�̮�㢤+�(����*^d�9�.y��s;(F*Kޠ�=�g��{�Lz�͓�r��Q'Y%[��Z���J��x//磓p4����8�b�/���܀"��yew��+3���p��f1Y%�w$F�����}�w3�U˺�o�W��k(���}B#�rt�ޙ�z:�#+�UI�Z!��t��H��=Ow&��H�� ��佪��G�L����v3��e�R[��׀�Q>�v�Fs�E��a�z�av�ow�遻��4��
��A6ezSZ.x�5}��vmi�1�	s��c�３��bɗ�;�ð�k�`ꊟ����8�EG����w>,r#*��U
��<�b��r��!�c�ޛה��B�>��e��%VN7iRu
$�z���)��9Z�5<]l��B�G��v�9�X2���$��i��q�ww��}��'��Mɵۥ�z��m`[�R���̭����Ջ�P�K����YqԺJc�]��^=���2�\��K_�[e��N�4��e=3e�LC�8!�W�Gy��<O��NɶjI���o5lꪃxX�����m�0�r�hq?N�{X��(nZ�>�͌������G�y�j(�.�J��S>QPV� c w��!���e�{)Vx��'�\�M=����f�zZ5��T!��;)�(���!#>تx�#��?=�;89�,��b�swb��c�V�LZ=D�v��o�1�y�SO�3�P���Vjųo�kW� �y̪���=K�SE�F�wdP�]B��}|�V���
��}|99�E_W���B�Vlhx5��:�w[]��R~��.�y�с��� 4 �X7)��mm�^F��P�ﺋ�ה��Kw1���^�"���ê(<%тT��~���0�($�ǝ�z������Ck���xf��0m��R(��*$=Y%�|0H���A
�d�;�w��:��v���p�ʱ�}4��3{U������S�Ŀzp�Tb�c���� hUt�@�ΐս�-�u���3z�Wa]�K�{Z�yX� �s{f.D $y�պ��\�[د�}�b=���ݷ������m�������`��˾�{���S��}U�}Y���/9=,���%{��)r�I�X�(O�xό��h���Vٕ����Mm��O8W�=g�ؐ��k�o0�z�t$Z�Q�h{����=
4�g��5w����S�������� =ću�:���l�m��R�?ϥ㩧Fv��%Ngrt�a��'����C�w(!�:�~
��kݿ ��j+[\f&	�ο,k$��8��){C��y�W��]j���`��T�i �&L�[����8���1��״t|��G��`�}�+�Y������3Rjf���ï_���νz57�Ce�S`/����ֱt@�V�9S�[���Ȫ�.!�;����Lj,�����hٸ\a������ځ���>(P�	�G�f%�]b�
���HϽԤ'�}n2��y3��Ĉ��jy�2�Q�9�*�R�2����G3aV�+֊��:��OLmm���-�����ޟ7�MdCh.���ނ��}���ȑ�Hv��tW +Y��O���\I����t宝��Jɛ]�I�{D.ASD�Y/�r}��ڼ+�<�4�]����P�߱Y��r��~����:^D���g�;H����X�#=��3::�]�e��4��|�:܏G��v)��͕�ۨ��2�]�Պ,s�U_}_}$�s�����=�_�u`Ӕ�{�2�VG�H;�_��E���8d��U�F[>�ۀ��md~����U��+m�x)�V8|���\�!S�8��=tp��ß<�@�i1,mq]�3�T�u�M�%�Bh}�B�ttl�ጞ����~8$��]%%`4ōj�{z�>ݦ�_iZ��R���Y	�G.Pu�]��h^Z���|v�L�9���v�HO�w�ߛŗ�Ӭ]xR�r�!b �E����Ĵ�{��i������\�/��[�U��}������F�����|@��#*/���!\�k�����<Γ<(��]�i>Ưp%8u�z��c�_P�ޘ,��*�T��_IV���Z�V��<���wQ��|�^{�M;��|��K<�C����!ľ����f1>��<0��B0?�c�]�ȴ7�҅����7բ��Yd�)�C��Pg���e��pWO���]�A@�V9%+���S�mq�ꓟ	Yk�;J�F1�:Xv�5�{R}�D�T=�d��p��W�.��Ӯv�8�ҫ�Y}��3��lm,�8�6 �7.�Yw�Ş4Ѻ�=Vʘ���[0ҏrk���Z����G[ՈM���8��r�A��t`+�u�7933�ܓ�t��{91�oK)�`_VmZK]�˲���Ŵ�r�߾������%3w�� �,W���@��$�m ����mˤ�P���Л
�]#��6�<��L{]�;��A�5��{�f.���6D��V|�@��$p�F���X���e�_�����}L��&��+��CՀz'㾓r�Y��!)�[�}醌ɒsʿ=ex*��cj2���u�@@��r��׶R�n��a�`\4�����{'9�5f��6D�|$9I*��[�����3���!��"�g2J��YR��A\�����K�z�Qٮ
�T�,QcJ�����0��l1���מ�#jl���[{�~2N֬��`dr2���H���eWM��ad����2���gR��(#6L�����Ӗ</uA��&�u<�aP��B�?0�6���\L*ĝL-q��<�ې/]���f�N�;^!Zk~+сJ� Q�Gh�ye��"�BzN�Y��
/`���5��7s�H��-!����*}�ƛQc����w&�^��WV�'\7�	��Dc��5jͩud,�j���;�l�<
��0»����y�C�iq�*�k���G��;�k�˨"m��ƍEXM���X7{�ǹ��ot��ҥ�!��g��r�;ncL�R�+opXOX��$�bU����/��f��e��:
�b7R��!�yj�7�M�T�M��l����K�k��&���Hu!ʶ�v�ދ��avW[�RL����ğX@�ր���r�o�7���W1ѱ��Z��^qQ�Ѹ�g�GG�>vIf�vH���>C�c�c����ܸA�<��
W���t�n���)Ct�*X��)ۦ��]�U�ӊu&�uK����`�����Wn
c̐s:���%vN�a��4P����7�bk/k2ڬ�v��ܢ�J�ι��7Wb9b��jM�u��pf,ү6I��E��#NM��wO.޵/[Y���vv�t�y���̱eJl�R�.�u�g���j͛�V 0�8k1�s��X��.v��K�˶�v5���FՎ�}�D�c���}5�0>i�fr�Cn��z
By/U���7wv�D�x,��������B����̌��ﴫޝ�l,ُ0p	�v2��1=�X:�7�k�]���Q
�Wv��m�V�������K��t�|�iW7�*Z��u�csN:��-�}�cwB)��®6̢�+��^�[��N=c"�>�v<;�>����e�䅀:ӫ�Sxp���ƪ� ��0kUz�͹�nD�R���࠾���M�c޷�IZ,�r�в�i� � u�k�vqpc_'$�]4�������[���,�n�+3>w�N�UyP�D'CW�<�B�����.W3Μ�0�+Enf��q�Ҫj���3$���}��iH�eN�u�����5�u|��qnif�0�2niK ���l�k�r���^�]JO�un��5c���rX��¦m�f���n�K�4�]}��oh�;��٘���������Ws�)lQu6	�25moS���i_V	�9Y�0��5�vS�,h���a�oG\y��W?��Rx��
�K\Ï7�[0An��3�*�='1֪6���s�[C<��.G�ʑ-�7��r)^����evu��z�4��[��2­��ج��	l/�Wf�[\�<�:���\S$F����k���W�I�uJ��]���2��e^��s��Wj��7�8M�k+lG�!�Pi������ �Rx�p�˔6�G��Y�5�8���Z�"m�'�Is\�[�\�����J��`)�d�"�pe�0�6_-��W)�Ƅ�d�w����-������m��#��v�0���.SR�V��ڹ�����(�� ��>]���fS=�-�]m��RŁV�ˋ�M�,�~�깫��]��k�ŭ�ӣmA��ǚ��h�Xҷ X�s,we(��l��WX
�Y���Tبൣ_gV��s�ܚ�ovH����U�mPTkDE-��\�**"�(ȫUPD�U+TcZ[E�ZU �b(0T���Z�Q�"Ƶ��X#2��p���Ab�E`�hŊ�m��cJ��QkAb"EEDb���TX���P��R�ch��QVڱ�J���R�k+"U"
F+j��"֑Q�,����AŌ��TBڕ,�V(Ʋ�Ehն��֢�c�*EJ�[lAUE��V���UP�AcZ���J�[mZP�1�X�ڭecRPQF!����X(���m�EIP��E�UAQ���J��*�X"����E�*
�F��$AF
,PD`��F֥�F+*TUX���QQQ�\�r�A�DE�Z��h�����U�m
 ��U��
� �V�Um*"��UR�J�E��E�Y`�(��%����X����U�*�,U-*�DUb6ш��1Z��QU���T����(#
T�"ԭ�,QTPm%E`�9e�"1Ģ��V�"�-�,U�X�-�B���1D�P�V����%�V+7�f��v���u�_��ϯ�J'z���_.��� 0�.W ur��/huN��ͻ�8Y�	�����7�\�VT1��������~F0�o���6Hc]�͘1yX~��̭s)}
K�3��Ie��"5�ڃ���ʟ�&����{�?�p쨀�V��̋)�fW�]T�Bӈp�k��r�X���ҧl="��@9���/�p�.�Ϗ*�~N?x�ͽs���X<��E�����ϭ�e��{��K�$+��T��U�d��3kŭ<`(��wxm�cQ���#ih����\�n���)��;�`w)V��ᩤf���n|�mf�Z��r��5*�����o��$�_U��=�-�+Y�7���0�x3)��6)Cb��tL��vѺ}�0�W�z5�w�d�w�[�%�OiR����n��]5�2�]]^��	Crz��=*U�98۾�X�e�a:I1�W,f =��W�lH�L�/�Bn8N��@��tH��r�y��C�v+��N���;n�}f�� �T˹	��bx��OY��s�c�ǦF�c�^63��lft�+�'I��u����v]m����mX�;c�G�QP��=��h��gn���n�񑴛���1F6^슔������7Et�̧�v}�#�s&E�Nz�i�{o;,�i�qi�D�[�C�ip��	�f���8ek��hm��x`�X���uv��n�m�e3ȁܹm���� �:{�nU��u�߾ɹ̪���=K�M���wdP�+�xU�u���8�~��N�M����^oU�b{�v�|g��u,z�9��%�)��:��e��� y��~Sm_��W�{|��gy���+�ua�2���s�y�]P�õ"�uE���JF��n��o��A�f�Id�w��W���!�����:�/�Ɂ�THz�Ie|_���,3�T��b��/�
�C�� �O":�^Z)Y>(O����>��u� ��x�mM^}�����f�	���
C��� �:_p3
/��䃫�챂��B�9xz���{u������ ���ԋ�S�uخ��p������{<�F���E��y����SgR*�B��:��zo������5௘���[^�QZ��[�:��R�yT~��7���ݿQ͂���^���a���Â�;K�2rn�]����q�S��E����'D�\�ZV\�/C��ۭ'��҂��;�m�p�jf�2=.�:+з��ܼY�-^{F�9�Q���c�Ήp��}�[ጓ�wY�j�
h�~"�Eoj�C�Xks�Q��7��e]�����Z�c�p�;���g�B6��V��&2�=N�l��xUIұ�b��!���G�us��]���=���_}��So���j�݋��0U�f�O�`�2���X�t�#+�u ��p����Cb�md4�k}�fk0{�+�ϊ��C�Y#�����z�.��u	�]q���7�w�"ќy�b3���5ͮ�xg�l{�_����*ΐ��X�_P�<h�~�����tH����͛{Լ4��z���,	�d��V�y�딵��=dv��H�����ϣ���mߵ�;�b�~��OL����)2Ӄ���ـAd}���^'"���� @>��ol�����7��U�D@kB�F�8i!�^̚|]��^���s�yd�C/>Sa^.k�u�2bN{��u�U3,����	���r���B�4l��-p�>]���ר�PWc�:yt�q
����1&������2U����r�Uh<�����{{0+oԵ��P�%�v�j]Z�5��2��C�d� ��?n���u�p7�asu�yt'��~;�=��$0s����v��E�����b�P���[�6 �%e*]��npl��w��	����w%l��A2{���[������|����Մ;A��!Z�Q�x�V���\�2tom�cj�0�G��w�Z�&ʭY�q�ҫ�}2��hS���g&���r�:�E��fyk9�O.�T%[�sz�AǗ�������x�o���K^l?϶_P��y��J��R)%[�s��"�kK#c�>��~���j�����|�A���u��Ϸ��'9�B�{1�T�u�xkjyz�w՘�7��9�4�xAP*�̟�|g�qpT�̕7��Uf��t�{$t��5��R_��)�c���w���~k
����0y������x���ÈB�u�|mD�|�����A���6E�\�����F�%C�z�E�񿒐�3��b���^ެ�Ψ�wo���Ő�U�p<�\��.�Mg�e���(7d@��~3�q�kL��-H��#.���-{u�Ec�§��P�ڃ��Q�8�Xޝ}��T���#����z�y�����?c�ď�*�*���îf�wPÞ�U)38��qs#`#=����^o��,�nK]oz�j��E�I12���s��!�|6]B���"2�2��R�?'��I�wnB ���`�(�5�Q�p�]D4�ඃ�չ��R����{����׼����+��Y�P�������XS#@߲V�ρM��SzN����H�떢�/���ٖ�T�ս�[��:<�ʽ�!���~ܙ��J9G�m8W,
�����$��d�,���uq�38Gu�	�Q��<:���:	m�o�� �~�z�����Կ}��>G��C�T"�VN�G����!�ɋt6��G�Ve��{�����^ץ�݌g�>X6��fu/}�<9�(;!�k���,�(u������>�9��zR2�֔��'H��3=]�w0�x
��5�E+ez080��u�n�9�&_g���6
H� ��m[g̞+�9��¡�D��	*�h�R��LJ�x|�:y9eձ��3�<�VG�;K���n86�P��^t�K�_�����GM��P��-������1s@�w�wzϖ>�1ʧ����K����	�ۀoOV�[R�!��	T���ҫ�%���k;���,z��?�esG�)�����qKnr]]ҭv��[\��
Wm��Ŝw�ɳ�����	��K�/�7�һɾ~�j�7������=KǴ�v��V�w��*���q沒���4�y��O�rB�ZI?L��Ng���0bB&+������Ҙv�J~,M�P�L[Z¯+�su<�@��& ��ys�����S9�8�U�s,n�F�޶�ۊ�:��71j'""G��ӹ�˓�(��� �&�l˨:<=J�N�,Y3���:Kf�����������K\���	e���]�p�QN�g<Ǉ|J�����k���Y�]j���#2�֒�1b�Rκf�p����d��}��C�-|�+v�kh�q�t�dV/ȍ����㔒b(���Pc@w�"�Uu�u)��tp��Ue�u���Z�ǿ}Cx�㐈H�>�;_Z��o��Q*x-�	����#Rd;W{Fyl�{�6'�c@�g�R�Q�Y������E1�'�� l3j�LvUZ�<1x Ϛ�?��}ŗ�=X[B��t}O�w�����ms�R�2�(l�5����`��-V{�7ʊ��p�1w�Q������3�<�k�bA9��U�H���D�"�l�����4�����oҰ��\�X�s���}[�xs�x���Is��+*�:�*Q��>{�͍��3!NFiAM�WY�]f��%b��)zzW]7V�����''����ڕ�t�ʙJ��)�Gx≊W�\ѱ�fW��pek�D��y=t�^D��8x����7��A�o(@9١�HIgū����"K������O2�ލG:ΙIK�^�q^��f�#�7i��Ϙ��'��.֕gmN���f�a��;r���Q��'8�ͱ�����@X�!{7�bٴ��S5/ޱ�ۡө3M�Uٮ��N���(r��S�q\�>4�܀�#��g^:ⅳ{ȓ�h�\��Qes�Ϧ#@wO��.d����vg����(�*����*�U(�ד�Bg��|C��3A4z��vJ߸�	�G���mh�7�1�G��.���]/���Ԭ��cDW}���O��]�5��{s�#/��7�T�p��Y��Z|+~)�]k�g&=��Õ ;I�L�u:�6���M���(��K̹{�3��Vb`�v�IY.R�2
�ۗ� ϵ �Ϛ�����,|n�2�ڡ��JO$�#�nz���0U�f�^�%cО8N`7FB7�u� ��I������!��T٭����O'�P�ك�/�T8R��F���砸��{K�H���s׷	󤪒��ۊ�5�/��z���<��Ƕ����S�<Bjä(u���)��
��S������^U�����ޔ�M��^K�er�9��)k9�;*��,�����1��l��@]�hg�!0_Ld�r�M؀�滤n)U%.)�a <;vi�
�=����o� ��"P: �F��z�j�c���̽;�qd�EC(++*߽O��js]J���71d���B��Vq��o_yAܕ�0�l{v��^�Δ���:���v��oF�NBQ����떠�G�7�H�ʘզ�+sz�;]N�	��e�M��]݄��.a:�g]Nȁ����Ө�3���_O��̍���>������a6�	�l�Þ]G�gˣ����������n���4���ßLx��d�'���k>JWx�����vehݧ{'}���d����k�����[*$�aυr�(KO��.���Z��7�ܽr���8�K{����h���{y!:��0vE|@��"���HT]�*��������VU�듛Fy/�suf��3�f�B�=�ʡ,�[��oI�ѭEU��CČ�f���O���o�B5�r��j�;(�s�h��T��)�e0x>�A��(L.�n�YX�g����=�k����AP{Hf�	f3å�di��Aâ�9W[��²U��>巺�����W��/}e��k��ҵ�ǥ���ˏ�G��=7�r����0��=�P��n�ɲgq�=}��W� Ӥ�Mu�t<l%!�����Y����\��E[���u� �:�53+}��dاu�2��#YI��	��Ps2��<O��)I�e�+m��:9��Z��'Kf�|���J��C��aPR�沟t��vA�(��|��K�nT�;@g]�_V�z�*�(w.�9�Yw�9����psA%0r�gOWQm���ջ��LkJf$���,*�L��Vz�u��UP.>��U�:`G����
�p�L��DS��e��ѧ��yJҬ�Q�_f�L׹�6�T����̳bP@\9|y�J��ʩI��S>��Q\�Ά�-˹!��s��6	�.�bC�$��i
v���Y�����G��}sf-~�ʧ8��	G����2����x���\�X.�ҧ��~#��޼��Rzq�X��9{��W�j2�UQ����\�؀�K�A|��<;U.�q2��]��%-�N{do/vU�`k�v)3�>���2LΥ��(?|�P�u�x�8E�/�cHS�}�G���L>�ıu��3O��w���C�ã�=���O��%z08:���g&��F:�d��Oo���aT`��Z��|}�d8�ҷ�P9y~z}%Z��Z<.��A5���ǳѷ8gh�����S	�[�.��S}f�Y1˔-9��Wո=���)N����������	֍�M@T��a����%���Zτ�7�.�m�&ˡG
�y�s�h����6L���k�w��"�H�UG~��8{�j�k;��T���	 ����u�m�Ѓ���tڴ�O/������x.�*�n��*�*����v9���owU�F_N9A���::��9[3��ä=�3���\�w��_yd+���yæ�a9J��v.����;�	�٨�L�s���Y��@吱{q�Z�eǤMU��9�+�*����G}�>��&o���Mf���b\�u`]�@������h�A�����{�ض�2��[����	����v܆v[���o��M�Zz�{���XWg��>�\����`���cJa�u)���J�kt����7�&s�|���,&=),ge%�	sԩS�A�Y�LÂ�
���+�u���W���^���ç�{�8��j{�F�t�m��G�,�Ih�~`'�� M@w/�Cwh���=�9��yXY[}㳠Cx�C���J�(�'a�Վ�S�C�u�MF���n�������X��3� �G�Bf�x�{�(�L"x���~%��t�$�3�ݨ$�Stz��5�|g���}�UD2ns*�沓 �h��y�"(]:*:I1��i�4�a^��ĺ��
3r`������<�k�bA9�ʔ���D�"��S��Hm��嵹L��H*>t�plK6Ց�<���<�&���k�z^y:��w̬c�*����}8���d���94�0�r����*�v����A�ݗ�V�f��T��\�C�E��k-�C.驕��Q�Έ��,��M;I�-ޫ���760z����[+H��^�Z�K:�n�(Uޥ�)����U�Zݮc.�CR����4q=�#4cN�Q�������n��wzY�;��e��BV��=���[٧���i�[]�B�t���+?��2s����m��ýw�CW`]
����]殕��ϝ�@�{���÷Yk������}@fڣMް�W9ח�@��v)�ȣNMQ�m�q���Hú���yW}yE��x��=4oW0C6и��q+��3��hX��M�ܜ��3��%fP�+gҠ�;�q_1yF#�����c�n��U�:�:[���SL��JNB^N��=ky�7;��S	{	Ò���G��sU��YZ��PdI���yuM-�5���&�q��C�T�#��][x	͵�VW:�_D�LS�9�ۗ�W��ۋR�Xw]���6�$�v5���Ko�,c�pkz��L�Ba�ɜx��ЩS;��v�l�i���!<���)�~\��qgb!7k����M�Q��5J���r��zؖ���iۺ=OGV$�{L��>���\#�@ʴ�
�q�-�xF$��|l�=MN�c�ɱ�|5�M/��֩���B٣���"놠ͼ�f�785�B�����U���=T��WeZks��7����-*��S��T]�9��]q��s�`��6�M�[���
�ً��ٷNcjA�b%"�K��Ӎ�����S�˝c/��l��TXk}jVi똺�Y���O8��'iz����΂�t4��z���X�+k�\�6GTR�͸��i=����yJ��Zv��L�ͨm�)�t�n�ͦ���+>�*ħ��vo��4f;�]�����Z��}y�zW_a|Ók��W��тy�n����&^:i<:���CrT��U�v�4����b���n�ט�z�ޙʒ/v��Q;[LT�y[�+�z���<�x>��[�����	;>%J�-�Շ�.e���7��knf�:��'\r���v�s�ы��b��2)��vv-/n��P�t�NX���
a�螩�	ݮ&���dԯ)^j��:�h޼�[�wI����\[�@utJ���w�fWF�Wkv�Y��q@�j'gKU�����(d���n�%]�@���LX/��������V[�v��+A�.�*f$in������k����@�hh8��lw&�]�Ө�6�v6��q �:�9��G+I$}w5u�
�&�|�w,kbȅgUҥp��f:��T����|�^�&5ռi�%Ml�48���5L�gD9WF>�/7�k]�I�+'g���x�V��2s����[A�Ox�u��{��һN\���   �(h�4AV,b(�"0T��J*���[*1-eDh�A`��(+iPU�ҕ��AQ*T�-m�#*(,cW����6�" ����T̸�*�U�U�(��b��DFګm�-QE`���e���F���cE�kV�Q��Ң��DEҪ�j�J��*)*���U+e�U+Tb��5�D�U*���*���T`��-eDQX�X���(�"*��֊�(��(6�EcR�*����0F �"��
�
1AUQA"������K[Q"�ұ-)Z�ł��Q\���QL���%��#iEb�""*�F"��b(*�`�*�TUAE#YF,�"�V
����m����UU�1T�DX����"��֫+,DV3(X�ATEQ�J(��X�T*�ň�cDX�b���6�*������1�����QDU��*"��V�����/�~n����B<1�3�} ���n:�)ʻ�쨦%9Y]r���� ���[:u���'+&i'��������������@S�Ү��U׉��=n`��b��"���K�u9x/ra�+����y�Oe.S!S��7Ipg�[ᒐk��t�m�N�LZÁ��k�orj=x�ë�&�	���e(.�"K�������lz��e�
�}�؍�*k��k�ʵh�Z|4vQ&+$�C�|Z���It��g���7BAՓ3;o�����7���쀽kD�=/W��o�s W�*�@����/�u��]�n;�TA^e�9� ����=>�A�`��B�C!�|��\=E�(*�|ǆ�S�s�ѪX��w]�x��)�j���N�y�<�xY����·�5֙�GR���T�� �&N	��wz��ʆWj��f���UÃ4z嵇m+�"^K�yxG�A\7/�A�a��$=ox^O*�M����{Ig	��ó�*³e��xL8�h7�u���)�& 0H�s4�������r������&�O|�OL�!�����x����-�^�<��W�s���w�\��K�֚7����X�����K�k�Jr�
��v�+��]v߸�܅������p6�=�n�~{��(� ������rh5Ǵr:!�����|/{+x��=K���ț3s�q��Nn�q nd� �A���Z���� �ӧl���{���p�d碔w;���{c��NT����+C�����`輢�-��]ɹ����L^Ę���L�0eOw�2�,�mJ�s����^�ΞF�D�:���6�o����;כ�B�'�"��
	�;>����&� ���)��_��xo�����/,�*H��f�=N��z�F�"�<h�e�]t������{N������p�}��Y��L�wkV��p/`�92�RY̘I.�,X.��5��<�����h�s7�����G���*�SOq�>%�"����a�dS�G�\��J��@qi{&�o��y��#�;�V����R��D�o���X�A���"H�G����I/�'���m)�Ov��
�O^q�C���خ�Q�`�_3��#"�6�B�����~'�K�y�w�]�k��$�٫!�������T%�ĕoI��h��]�y�=f��Ks�蟓���f��k�%���2�Ǒu�=鞇G;xF���=���/ex���!���C�5K9M-)Y�c����+���r���fb�xR�I�P\Pe1ymN�bDSyk�F��"��VO �_��79�4�q86�}�fu��o��lͩ��:>c�R�νU"Y����]N=IoI0s0�:�:��wꪧ�v����gk��5��75uAS�]a� ��Y��̂k��2��LVP0�u$z|���{6G+�������d'&�q�l{���-b5��i].V=.>�f�m�b;�kJ��A���]���[]�8���GDd�3����9^�Ӥ�r�PT�x�1"E�ڻ��v%����7��p�Vӄ����%^ވ=# ��[��5���P�Kv<U���$+���{,�vǊ����낼=��3�PuJq��qV}�������d[Ot�[�ܜT��W� 0)-���=pX�3	_;�aϽ2�R�2��̍	B��7���u��u&v��U�;}� �,�d�<��*���7D:P�CP��kƶ�:������ny-F}�s9��2���x���G��E:�1�O���^��>��4Vf��:�V�}}n��z���B;P���œ��=n����ym���W��`�rt�Vs6��bb�%�<^��cB>X4z�L�/Ց<8)
݊5ф؏<(��<����,��"�㇦�y�nR(Yu�-
�R�!w��n�Ǐ�t:�9���Ԅ:��bPo��x���$��{MKz.��?��^{�Ԑ�D�t�_v�ϱp�P����N���7s&�j	�$.��iW�G+��	P��q��h��� ������j>�X�Me�]/�����!����~�!^!�r�ܙ`p�]U�i4�zg���z���=F.� ��h�{����p�GJ�=>��[�;�W�s<�&֔�c}�s��ڹ^��_��xg��L�U�:뵟ϵ̤M��AKG�����q��;�;ӑǴ%n��k>�dh����#��*��B�g��Re_:�SG�p�x�����;�.>ۃ�,�7��A�R_��ggr7�+�>�j��<�\Lp��#/�
�M�u͞�c�߾�i�je;��>�Uk�UPRy=���������#�<}�0V�{�/�(��ޥԕm��i�ˇ��rʃ݋j`�*�Ǳ������z����g�Z���~����U��*hiX��.	1Y����n'Q��}Z2���lR��X�/zt�5#~�-zwj��+|��
�b[e�+IѐX��Vq�a�t(53%��Uhм��ֽ;ZX�L����T��x��ฺI1@'F /H��Y^�+8�'��1f���WK��n�$rH���u�|ܾ�ugb]�k-������8��\�ڟ�EMr��l۬���ΰc�]ѧ��m���7O3f�o16vV@�ܚ��Iq�'��:�`S3"� 1i���Jr�<g3��O�]|h�]�qa�'���ߥE���V�{|��zz�՟�Vs�3�bz{~��r��%A��:NÉ�Ac�����,Z�-��tsz�l�I�=��x�^H�K(���ϻB��9�u�E
aQ,�U��硫���Y;�-�1��g�[G�.E4��({e�G�s�T�5����Cg��ϚDPs9��=827o#����T�/��6e��E��3�<�k�bA9�ʼ2D�R��z)���-t,t���y��4�@õ�A¾Ϋ}�պaq7�<C�¥���s���ͧ��_j�l�v�1���ྙVj�K,�.�����rU��ϊ�6çZi2�c����8���Z���Hz�t���	�bV��I��K4�qD�+K��c�ă�J��L���s�^��㕞۲c2�<�LV��C�ϊy].x����nW��uqV6x�_��s�_��ve�\� ���� .�"=}��c���޹�����b��B�s�� ��΃�!�����>Fqp��]k���}OI�Ѡ���h~r�+h�҆z�%f�ٔ�rƦ�I��rH���č��-e�Ru��Bo�a��D��f�K�=��c����=�G9Y�ObK�he��͹9a[��g�Sl����Y�����N���b�HHKlk���8eǴ�%�73VuAm���rG�����#^��{���g)~�ؘ'�̕�Y_g�0:�ܾ�ƫ��H�bd�^���֧u=�~��w��4`�-�>���2|�%���u;_��	uꝻ]�+�R���%&�)��5]j�g[c��l���W�!�Ƴ�������D�|�_])�
{���(�6�>�/*{���HwǪ'�QV}.��h��Ks��\���x���8����+3�&�p���@�v	��Ƕ=�_�੅�����Շg������4c��@�K�1��u%���r������Wd�9]F����1�X�%3�'6�����,T'h4	�̥��84�:�����>�AC��xxf����ךOt��y���;}�p�=�E��AN���D�X.��ӿq�Bm���-��y��.�uI�������ơ���ȚO���\'TxR�u��xU�=�1���n2��^����^���i�K�E�.aɂ�A�"�s�L�����t�o����fz���R�`)|`�%���L���Ŧ�q6�m����X�uga�2�1W���[�x�} nG���}��r�ϊ��� �b�]�ד���-u��z;�:��`�Q�0q[�P���6:�*�YFm��NH�ۖ��x��c���O=�������۩��"C�X��S�D�o���W����/]_R+�����z�6�^S����y�:�;ز��-	�a��E|@ʩ�#>��ۉ
�Ovv�w�q�}�����d�������P����3y�g��eVTE����"����#4��{u�-��~�z� E�U�R�P�DA~>yn��C�s��`ވq8�-*�Z��g�#�R�/L]_�!-�<E�z��>T�o��/�����x{b�|(���ys|�#�.ct�4���k��.	���o^z�t��[����Q޸�Bu�Wզ6Wo�u#~�X������mL�Ĩn=Q�d[��'�g*c��4�7R,U������'{͵�3X�b]�|2T�z��%���cS2�âHϦ�;�a��i�ȭ��|+K�����:�L�>DS!�P"�E`�t�j�)�W��=^���nx%k�-W�����Gfk�K��J��D`LL�-�2�T�].�N�/�&�܄0�z`_�E�c|���;�Z�Oi$#��o�����eQE]�t�՜y4\+k��v���+�.w�����&�O;}9vJ/*��x%�hY���{���g����ݢ��b�<��K�}X˗e�ǋ��u'���:���2�VK����ˏe�>�c@�V��q�ﾯM�2���ߜ:ߐ���Ҳ�/��Ç���E�`�!�I12��]��J�Λn�;ڛ��k5�u�n�Ə�#�͂á�fR��⋳]�u8uQ�3�:��r[�)M�왾|�{��� >Ž�%z���Լ1�ϑ�9BNHД��<8�"=�'�M�PV���j����l�d�����~=�[��';U��I�Խ�<9�!A�v(Ph����83�E���/N���z�ɖc0����\&Rھ#8������,�T�x�r���t��s� M�����x�� ���q��U�s7�
C��Y̧�)��w����d���3W)3���G�F�Hp�x"�O�<3�Jg�V���|_f�R$���Pzv����-v�Y�.�fh�쳢K5�/��l�V�*���~~�8:`ُ�I+#�xL��ݒ{{Q�,>9S�o+%�/C�1HI~gI�vt�7��y̻LV�좘���W�x�8ߵ��с	�K�O����_m�\���}96s��f�ϋ��9C�3|�Ի�g�׼�k8nй�v�'��:�a�V��ğ� 
�{�m�'��+z�������hM�u���e=����8|��\��Eܮ��4�̀mɕ��ӗy]�>y��#kDl]Alm�:�p����ï��B�,���~)Nѕ=L`_��K�#xm\���
���W��^��<7���FTݺ�>��^�����+a�y������9����F �Z���6�N�4��W_0�Ѷx]F;b�w䏩Oy�b�����7�����3�|0���,.��u�0�A�8�����~pMzޭו���ϡ�+{�{��-R�t�<N��RLL�倪�Ҁ�F�C�c�{���ط���~|�jF�:�/���ʺ�`�j4�2�����)��P�~~���~�{�K��V��/_2FV�U<r��G�X`�pev��s������tQ�����8��oҗY�T��yiكK�}Fz�{b��&�2��d瞥�e4ve��.��<
���m�a4*Pb�D�=�*U�/���m���yJ׿��s�b�"�,֚���K��d��,�}q���|�
c��]�k�bct�|�eoxŞ!��B���d2/�~}���<;~ɐ`Ϫe(.`D/�G���SE}A��JA��QӝR�j�K�}=�ނ�޺^$��}v���Y��5��5��ӮQ��\�sB�Z�Ș
��ݮ(m�L���hu�Lӭ�W3���;p�Ӯ�jM��L��ǎWe��+FK	w˗�p9s_$)>�t��)$�����藴;�f�hw.;r�����ɞ:d��^�qy�e~�K(�`�	� �.R�d���~&��.fOM��Bl�9�6qY��������Y(3*S�Q&+�hxR����ݮ1h�e!&F���=6p����:x���O`H:���[�}]�a��Z���ʧ/���Dz��ac~�<s7�'��OSCE?|�<���f��YC=�c>��g�p�(*��gaP�v�,�@+�����'?&E{��։��ej�2|���<iԼ��&rԙ�~���U�F{�Z��o��nF���>��a���gD��ִ��i�]i*OfAZ�P��6�'VEL3��@�}6���_��2�S�xn���ףl�VY��D�z�`.�X�և�,����7�e/i����U���X'�����H{O��ك��G��p��h���������e_��y*8tTP[d�y����R����я��~ӂ�S/�4�gf�:k���:mf�Ы��^F]"��R�����ـK�u��Q�3��-�+�^������p�F��s�*X�ӭ�w�Lv��lvڿ��E�ě�lG[<��KJ�APEUJ�����U�;�s��Z�M�>궮;{�}�W[�#�/9����"Ӵ�� Q�J�Y.�L� ���<�\��:W��MewT����'�=��9�H�	/Ხ��м�d��Mt<E^�:��>�0���|�WL@JB�4�ۄ�b����n7IZ�+:�N�� �ɍ��i=�v���Nb��X��GE�_mp:&�d]����< j(t�'bwK%+z�f�Ѵ 
��@��'�HP�(�&��!�#1{р
�S���W&-m"؍�:D�n/�\�:�^b9�{�,t6�=
�C�q3�J�����+��%�M7���=�I���i�n�,�iא+���{�e���ǍNT�T��X��	��J
�:%�G�_V��5Ag}԰�޸f٬�وE��Ԣ�=ئ����AHh6�Ѥ��/&^a<l)(eY��8�x��݃�%��sr��Ec�t�쥐u�h�psոVX�����Z�}�fF�m'����)��w�uL�/P&e[��KKOtm��M��QxjAڷ[�Iq�Jnn���E�[�`(^bYR�<����[:���|S��L�bβ��دh���T��b{��(����)�N�ӆ�Y���tq;9T�=6�r�Y��Q�5�#�g������:�q�ggV�Ŏ�� 5%9�8���r�u=Ւ)%)�V�%��w;�Y��K=��j�y��g�$�7��3";��<��)E�;��^d��Re�w.#����v�b�������	��u*#)��7l����殘�;���o�N�t�X^%�S�s��1��Z2�����]O:���5�O"���A���$�7�.F{�������+r�-�C������T�3ieN�ףG�i�S�,XI:S��w����n�}k9$��qݫ���M[��[�������y�룽=�]���hIގIu� f�YqU1�'�,b�%&Bo6�	�¯_��u�B��oP"�q�ML�ޟ/���3VA�Y�\�X�J��Z��#uQ����@P)�������7´�ŗ"��Bށ�ڮ*I�7����PwP�yg�n�^c�G9U=���$B�hُZ)l툾�5��Ic�!;rv�)�=͵�lA�ֈ�L[f˳t^�zƐYձ�����є9��X"a��������'�a-��EJ­����ؒ�E�-�ҡS���q�G3[�5�7���(��S�����o<��
s������2�o۷O���Y���o8mi��b�0`��銹����g*�nIcRs8����L}̱�'�z�=��1��v�(���:�&�(n�x�P�ٍ�:�87Jm��8��Jt;9߿���}��~���X���QPQE��j���QAiK �Z�R1m�*,EQ��R()Y`��ZQT`������*�Уme���b��KKEUb1r�1ULJ�¨*�l(��2�U���ʢ(�U��b�V���[e`��bUEd�Q��mm�ml[,�QYm�E���[J�.eU\[IFR�5���iR��-���%�X*(����ւ5��+-�+-�"
V���B�E�ج��E��X�1��P���J��%�eb�KJ��$A�E1��.R��e�b�%`��QQ��[E��QJ5ETTX���[PE��j1QE�F��%T��ň�cE=ʨ�cH�E�b�4J �H��Em�U��33*��QcU��m�b��Lr9j���EJ�Ke�������Q�ﹿ�\י��}ѝVÓ��k�u=�}��G�y���V��	S{wZ���LWvoĬ���m�E�:�N\iU�>�'�h�꯾+��N'�ǥ������tK�
|}W-�Ž8��8{/= �s�Ґ3eGj+	����c��;�W���s���9�#�T��_tE�`��4�Mw�9���{b��ړ��S}�)z�By{M�D{7V"�tϔ��q�[��VEX�f���{��Q�OA��4?{�DP�ڊ-�[or�eX��0��ϔ���d9�ላ�R���"*�٦J��h�OK�ο��=Ӓ�W��~��]��l����:Ɋ�>��N���GE\2��,M�: ��eK%���؞pS�o�p����V��/Qاל��>�à�|@ʐ.�2��6_"8�4�����m��PfUX��<W������Ր�z��`���#*�TE�/ƥz��.�k��q�����5�U]:�D���f�X:��ν����s���N{j��
Ź��[퓧zp<��J��3*��g=Ќ��%P���C~�W�ᗋ��2����������S�O��[:*}�}A�!��c'&޳�����2c𕖱���[O��ǚ�%��u~�J��C��oN��/XA�C �Eb��բv�˅v.�|��M��H��Z��Y|���kG�+yP������u��W[������ܣ�b�/6��g0���r(a�|�,7���r������iQ�¦ma�2d̴�]�
��3�gv���pXG�<�/c���@{C��l��tO_q�3���:J��dr��!�f7�#����WC!�o乕�-T��p�7��53+zX~"y�מ��������G|ӗ�b�}XE��6�C�Y�E28��P��{��gl;�����U��h�Z�^���q�s�_�p�g:�~��dptt-��3�H���b�#��PwP�誥yfm�]�f/ T�_y�2�m��g
T�YI���{�,��Z,��$��i
w�'}��8�:X��]�T�_�!�}�ShB�>ȏ��f����̤; i(�5�WS�E��l/k�
/5Re{{�g���^�������3�{R���YKq�ϑ����uB/�DWS'E9��E�qi�㛯3�Ƽ�����l��4�m`/��3�>��򶔉m.�dO
B���#�m�뭅k�y�ue
�Đ�d[�p�KW�g8�� fg��1WT�i������/kul�/��8R T���n��]��s7��){�fO��)�~5����3��`�ۙ#�����;�ܝ»w�7K(�0��z.�C������bD�IRѲY�g�z�b�<a����!n���8&gw0v�vi�7hV��R�|��s9��t!�L�;�X��ܻz�R!�9|�;H�Fmu��5#���{���Hg=����*Iy���~��[�"�8V�����U�;�oȱ[�t3����_��7���*�f�����!<|���bR��ej����??�[oE֨�i\{��wc�z�>���ފ�O�Bӈ1Rg��O��JxNƫ<~}��gfX�>fy�WR�e��9�e��~�j�Nr�]� ;�2�&�<wSw�aj(5�g=ٲ�7վ6m��#�s]1xn��fC�Չ\��L��4glxjo�{�g��3m��}�m�}��8�Տf�ķ�����:�I�7�&������ϚS�u����t�j��}�� �py�o]5����޷y��<~J&�R�V�WP�hq�y��^كf>]��؟U�H���%2����3n�r�+"a���E��`|g�-�������z�v�����د�V`�L@k+�n��Tϸ��/~�*�Y�r�J��0�񵩎F�e��z�����¦��hl����.BF�50�����eQ�Y���g)��ϊ�ŏ<=~�~4��Lm=,�s@���@���"0�Zx�t�䥺.�e�{�����U�Np���3ͿC~�0�y(����}����a^M�|�V�}���V��Avn�C��h�u6twN�o\a;N�_gs[u1RT��[�E̱,�a��1��5�HWvxw��<
�.�[�i�yJ�uQO-�OoKꏇ3��ZƋ���m��[������䈯����d3,X�r.�w<x�)Z��6���(7�2���ʳݦ�j�wvj{&��`~�`x:���PO��Xp��V/�t�[�5�����xu�p�q�3P���j���Q�L��0"8�u�\)�b�j� ��$��13g��V>��������d���D��>��>"�L*"I���|��XĦt̻i���Q�=Y���|zz#�+�VJfT���LVIf��/���$w�%�Q���^�V�=�4������1�J��7�\<��5�@�9�+�S� \ �����,�Z�Kp�o}�E�.'�z����ЅC�Ƈd�����{P�}�ܽ�<p��AWOcF�޾U�oU��pqv>�[��`���bʖ�+[^?LL:ϟ�O�iL��_3������8v;͆w\�8�P��N���.��t��: ��-0���\4��V�}�t��э�iRF�߻򚢵+�:��}�h�3�oO���ggк��н>�7�9�^�R��>�vw)|ٗ�k��8wy*%*�.+Í����(,��껻�k��2�+`uʆ��cz�u:����;,�q�x�0�rY�������>;�c�aj�*R�����!d�_�����ףn�aY��D�zK��Q+8�W�{���j��|k>��UV�u85	�bz}��H{O��̭��fˡZ)qq
��lwGw����Vv_-����V�[��y����P_s�O3q��_�੅ԯo�^����y%��|�XL��C�(m�h�~	J^M�^�PM��dU��<�_�(��Z�9��K�1�k�kE�n��谝 � S�U�]�{N}�7~�}O�@#�z��~WǺ2S��j��^�K�Ϝ��>�(1�Ѧ:�k�9����P$���%�~{!�x����;� ��Ny�}��r�]�9��[�ՑW��%�Q�)С�v��{�^5=8����Kۉg�{=j�uV�C�T1u�\Â`��x��d�&Zw�����BM^����z̯)�I�^�T�j�:Ͼ��b�O�����";ACl�U9��y�R��{�\jߺ����z'�6��~7��o�/����`����Hig?v���N�k�X�S��^/QcKv�ۘ��/>��m5_ze��OjoT�6��C��<��]x߲T���>�m.�Oi�e�`����ܖsD����x�SK��Je'�%��9��"D8j^w<���pYu�w8a�0�u�|c�I���F)\�̺W�7y^ڕ}⬾:�%!�f��x�����#}ܠ���f��>�3������W�	��F?�pu�C]�z"88r�.{�=����W<��G4�.7����ɏXB���	���ǆ����++(e8/B��g�0Qζ^�}�'�y'��s�Ql#����.�z��/l�(�M:/sn�-F�}~K/`����#~�S|oR�}�����!�𲎻�������T5��DO6�Kúg�9^��tP����A&��w�+���)
���x�K�C8Z�+<v�'U�������i����k=����^�k�[;�$.ZF����q�:�@c��/D�+��-�;a���+�TJ�n��e
���r���[u�}�.i{����,�8]Qa11-�1LU��T�0��܄0��7=�� �yɷ��(,k<!���F�}3`�,qh�.�bC�$��i
ef'��e#:n﹫{)�0xf���P���#��s6��v���.�pB�S��
Ū��C�����l,�WJX6~�r���;VaːߒkEh�}�{��\�����Ga�L{��`�:�oM����woz!෌��;�N�1��p�9$�^���NT���:��ǡr����&��\x��V��d7
�8ՙM��WϷ��%�����9�O.!<F ^'6�T��OVU�MN>EЖ}P�D��׈3����ὶ�)Y*�112�&%����˅x]�?���`��1��dO<�"3o.��W��7{V�u����up�R�,[�_�L�1�|Fs�k�fz��S��j��X^/���cw['��g���,) *�y��B�.뙿��Hr�ȳ��e �`ɂO.jv�]�"�=�R��ov1ޱ��т����]��������i���樄f�p��m^湪5�>�����%9r��3�YgF"5�ܫ��l�j�_�}L���R�������%��W$a���=e>��
T�S�}���>���U^K���G�6n��_�v��S�݌�r�5�~��)O[�����eU��J�	<��^��-��,[�vG5�ϒ�=7O|}g�3���1S�2ƬJ�^���3�v*�d��m��07�<߯�OL�4�v�7uX���1K�n� �Z���F�n'S����sֶ�i��a�b
z����r5|�]�{Y�Є|����ߠ>�}]�>�W�1���;�u7�\y�)��]�����P�ǎ�Wp��z�Pδ��S
r�����n��v��}\��:��}�l����V豹��k�nu���~Ko�������k�z�������&˂��/F����h�Ьq:�ߒ�I������������]ܼ���]����>�P�PL�^���2�oLBP� �^����..�LC�ϊ�a�S�K��֮futt��x|��I�'bz{���/�r0]��U��,��}-{)�\��۱�r�!��^-݉��BF�50��@K��g�`�pcڹ�>��A���Mu����E��j��H}4z�����-�4��{bvM��ǲ>����-�Q��y�ó9�B�y���.�
C�m �T���Ⱥ�m����)Z�X��y�?����=4N]�oo�7������n]��� �S�Ү��]bct��:X7*fj�:���µ�G��J;y�N���dS߲d2e(/��G���멃~��b�qui,�7�,�����{7�z�ɺ����:�8.d��Q!��%�|2D'���,�КxvtF�X��2�ɽ��Y�,T.]���U�^{�㕼����)�v�o�K4<)}%�� �T�+�^�4|���BV�?ncΦ{gn��4�E��{O�������7 �t���u���:��5@LӷI�����g�����ڡ����Y����q8���]N�s�@K�I�����"��V�˻z�w/�AdZ��MS��'= �Ck;=i����^����s��-|� ��T�ԁp �d}r��A��בΆ�7���ͨ~�ЅzPdt���f��
ߊ{G�G����z��uO���H�I���.��z/�+l=����\6r����9�k�i���Mu�r�1틠���:����Nv���+��z�'&�a��L1l����Za9��.M�E �</`�tBV͖������>�\+�5 �w�d,�=����WR�����Y��G��������{cRk�<���UV��y��UY��L���Obz}���	�;׈��Pso%�f��a��mf8�2�pU���&����=����<��Ƕ��Py��M�s��&�zYC�Ƈ\%����A]YN�8��=6eTYڕ.�U-�)?�)�9�f罦|ؽ�t�4�葧H�|)��C�AD��x���5���ikpr}싴���'պ�RW�)(��s�G��:hVԦ#��<^z�B�+a�xm�u��< ��^�E.�S�����F����c�=�5�˘��>���7����m\�Ϯ�W{�tͩ29m���-Y����O�*"9�����w#ݕݕh��+%1˦�J♡�%�1fo�dPL��W��N����\�ӹɅά<���a���9��K�2�!���*�/�VEs&����O�v��*�'ϟ�����.��	*ǫ�t��.�W���/WT�x�b"�.aɂ�@<DW�����y���{���Vx�I��ZLl�"���;�t;�˃�%�΢�ghe�{�b9k�%rzY�K����<�/�3���*�����|:'�rcf{Og[�<[��]�����K��*�D8_x����V�!{5d;�h/kB�t�����c0fy����p���hus��'>�21���k�؇�:G��+Nu�}��5���Iu���z.�k�|F{li3�z-|�c�T�u�xkɏ�*jߥ�xE)s���H��(�;�į{��vC�|߉��-�Jq1\�*�z['����'�i�{�piv�BnJmy	�=s��U`���q����ǃ�"�c��]��d���T�1��<�!{@�:�֗q���s	5�������¼mH}_c�c�g�ӄ���Ʀeo� � s��z��k��1��&�hylVs�L��o�*-kv�w3���=�Z�Z��A52<w�!�H2cN{�7�8>�S˚�c"��2J⳦�V��e׻��~g0`��5gk<�s@˥J*:��=��@.���GQ-�1.�]���M���[��m�r�@��`Sq}���{0k.
wu���r����z2��o�y�(U�`���
G���3:P"j����ݦ�ͻ(�X�h/��� �"�$*fe�Z�F �V�$btui*Q��u��v7�ը_��.f�$���ovQU0VN�m7�h��++�5KChS�+|��x��Փ&hr�t���{paz�CϬ�so�B>D}{u�Ea���\���U�]K�HRڄ'��u[��V_0�޵|�zQ��r+��<��ހ^Wf�f��v�'�.�m�YÜ�V;����O���4�L4��D�Ú�ɺ$�<��&ƍj<��:��ݞ��R�D���}g��YF2�f�ٴ��vU�P�m���"������otՌI{�n�#K�Ι��q��(s����Z!l�b������&��[��Fqb�g�U�����ϛ���)c�(�A\kk$:<<x���92j5x12�����@�-�kMֽq��uyzZ���L�iꡮ��jnuk�K1�P��K4��md�r)�С������ANv�|i�(�ބ�P<���R�ٲ��)�/V�͆�r}َduٗ���vc���;�$61+E��K[�S�n�e4�3^�w֖�˧����//*쳝I;�6�uaB����/2�H��n\}�aSr�u���wl��WR�3jޙ.�Ǽeq�0T;���c+��Y@���rw@�-+�|�#J�AlI��q���o����ԯ�y� &���T�X�:��햦	��*�t&n­�;Qq�4��B�r	Tª±t5��:�C����6U���pw)��˨$J ����$���u���,6�d���N[��(�x�h�[Ɵ|���O���m�ĵa&X��d8 �$&]qވ��C]�Pq[�񺉀��egJ,��&W�7xxY�m����D��].ܚ��WEso{xM��Z�S���"���R��|��úf��a�m�{I��9]Bz.�ߞB*��4)^�(�ۮ;�Ž����]ԓ%�����JEjAS[c$��&f� Ц�gW!�e��-��Zy���P������C~I��������ĩ�d7��������OZ�J��<�ǑY�em��l��%��r�g�جɥ�z��|ǸY��y��S�����r7����b�o6�VUZ1�j��&u��NΙ����=��X���C���[��b�,Zr������b��\����Y�nP�������Y*=5���;0,��N��.7:��L>�˚�Z�7ں��*Į��pM�@Vs�g�b��4�+�Z;����k綷n�)�O����\�w&�]˸W]]_��-(�"�c*��9h���%k�_������PU���bR+�\|pb(�H��*�EFڢ�E����H�|KV��TA��PU�,UT��eQ�yJ**���,¥QH��������q��UX��ŷ��*���U
����Z����1jVQUQd�U��lDR�ԧ�ѵE��kZ�"�)FV�Ԃ����1*�X��<�̩dTT���E��ƥEW��mbV����A�QETkH��[#���DQ"�a|�V+1�1�,EQRx�Uc"��e�*�T��#�*�J���KeUQ\�|�e�D��ł���",U�*�1E��1UEb�X�m(�2�墪 �V(�����U��UEDTE�X�i(�DP�-��y�����#�׾ae$U�Ʉ�eEܳt��s��Y�Wp���F�l��\�tN����5݉[}}]�sU�9�	7����7E����9gQ�P����
χ�[�M=��#����>g���{Ϲ��j�O�:�Kߧ� ~��G��bb[f`�c�/���3	�lw��k��{�\8�Ͼo b��`�][)W�V�{�,�d�=@�!$�<��E������dޱ���$*���>g��lB��">�g0l:l�C��㠻5���?r�����?8ߜk���}��Ҩ]��SV�T��O{=K���+�l@TZ-�fW�>�����R�X����#�)��ź�-��ӡ������1�>X4\�z.;��1/X�|�}�^lzM�Ц���
�����]��L�1�|Fs�k񙞮�=����yf=S�:oϒY��}[�i��+� 8R Wo"�#�w�u��W�){�g���!{�p��r��!+|�M?TI���j�`2�jbU+��C��oۆ�u���/b�'g��b�z��]�g���,��B�s1��%�tIf�������`CƦ]ѿg������e�b^K����E�3_e����w��*:L���k����X��j���w�~���]�w�K# n���
�i��U��#it�x���V���w_�:�wa�ݨ��`���<�
��$oc�%앵3���OVRV����8�Ƶն8/}�z��L��SG��e���Z �/��3��O�n%*�m��Yo��ݪ<nV�e�8����}I�	�~��>��8��U�Ϸ���~ UԞ��G�1�4r��[�'6=Y�����dBnY����i��HaL���d>����c��>X�X+��t/u��4�Nd����n��oV��P擇2�P��`.	1Y���V���K������o����>�n��������e���f��Y�1�䱟JK�	c �f�|hl��&ۛ���<4R�^:e�����~.R��=�P��`{���,�4�]�\�vC���@����<� �� Lh	����B�#U3�����ʺ�`�j?�*���-�&�k7�i+���bgȮD�oˮBFl'�K��$��eo�j�Ɲɾ@�I�����¯+��Y;@��Y���mY��S.P��b��d�|lqW���a �ݗ��9�woEõ���5�DP�t4U����Ŏk#�R�~�=��4��R����K�-kYw��Q�<�5S&,�39����|G{�M�\ڑ�t�Kv��2r�<�7N,��┝m�ޤ��0z�R&�l>o]t�cx&��zj=�.��o�u�&�SWe鮰K��}��	[��c��/�u�;6 ,!��ޑe�RVhs�-�T]���Br�=76�׾jD��I}�wL� ��
�" T)�w�"Å�V�X�����܁eo�Az�k�kbx_�\éE)W}0\�������u<���\�>��F�X�U���":s>��9�̘�D��$���	�r`�QNm��㌢�����l���4�e�t-�\�U�fr<r��欔̩O*$�`��
_Ig�yf>w�|^?r��N���y- K��#j&=����
�߱p��a��oe{���-,��U���&l�E���vY&Z�g�8^��Qn|<��Oh�_S8�����!�=M�⭽]5.�Ч���*�3܍@ϩ�94/��Jʊ����&�:׊��E=��+�	X涼�'��9L)��`t�)1���;߻e�97o�{.�b�gD�{=kL�%�9�n��w��O7r{�i-��mM��b�7/�A�a����7��Y(OE+��~ףn�aU�-w�,�W"ծ��^O/{e�j`�����]�u� ��u1��O3�(Hw��l�ݗS���9V=.��_���oCr�����2���-�}�������Py����᪮�Ubnb
�4{�Ż���ի�X��.�T}N���V	%�j�,c���;�����ꆻm8�7�U�:����|�����<;�:�U,a2�L��6�k�`��.^��-������Mh�!9��v	�º�T�L������̝�����b.��G�@�Xt��՛.஭��J��\��2�	��_�d���4*U�����i�HӪ�<+��&�2�Hv|�g�bV�(�����+�~k�����\Z�����72�����+��:�=�7,V���g���]�߯n��r���!��yd�C,��5�����s��7�gsN�M1��c��њM>�;,>ՕG�g��z��2ҡ����#�a�����*Ǿ��+�i�4�V�TX��C�*��]ga�8u��)O¢N��K�t=���|��Y���P�ۚ�5��.Z<�7��Sp�'Z��wR�2��Wz�s٭������i?i��t.�8�ߪ$*�GE�h�;iHi���'2]�tөG��F��[�./��wo�lA,��.�g"=��/H���X��:G��6.;���k�c%����;��zI�����9�K�έ�5o��IC�ʗK��Y��n�c��n����3um^`�����8�dG��=��y���U�C���ǃ�(63[3�v��e@0}�����u��V��[����M�y�J0��\�b����N�ڔ��sQ};8�;�'���ٌP�]x�m-�R�Y�7�S,����M(0	����Eug���}Y�I�ܽF
����X����ʚ��'�	�E����F����]�Ol2z��<>>�ڬ���#��!��^��!yz'D�{����cd4���Ƌ�<�8}����1|�x���(x�R3��b�[N���=�6�`8����ݫb����W�{�[����uj[dS#�P7�(+�[�|#�y��;�{��s��=�uXT�Ĺ�^���==�{r�G,&&%�f"��=F�c�Y��oc�Լt��CK9U�A�3���ƽ��y��{�`��!�Ǽk"�[���g��+�п4�[�J8)�C4��P��G��#���`A�[2��i$oeea��<��iͧ�݁i����3��,iS�m�0�ͽ+j�{��^ƣ>G�B)q/ofc�ߜ����*�#BT:Nк1Aة:�Y3F4�max��h�3�Nv��R7�]~J��Ω�l?I\������{�U���1t����{ ��B\q�o��;���5���w��I�J�3�[��AO�M��ѝ�/����>Э���32�o��W'LY���jC��/u^�3��zbSiT���W�N���f�,ٝQ��x��9t͇����EeP�v(P:��+�<�g�-�!�	���pQ�w��[��������8�ݿ[�N�	�
(=�,B�w�`�#е��}���Rq�(p�{w�;p�XXt�{^���!��OL�n�*T�O��"Ål.��q�4:ȋe�;��}�Պ�.YO�8�9�oLJ\�n$�HO�����2\��0��3��^מ�/9D
�(px^Ԭ�jʜ:�#+7��WϠB�*�"�'�9.d�Q @yK}3}3�;�=v�������r�1�9nx��~w�G�����v� �m1�����{�E�\��6=U���5�	�`��Գy�\���榛�*�]�Ki`�h�wc�!O���-W/�)�/��Ct����;;���N���� �X\b��c�N��L���}�-Ά�g�7.�K> ~=�M�l�����=Ьv%�f%���׶�P�R�$Ľ�'�X�K%�0�A¾jfJ�)}��k��T�J��zJ=G�����ӧXI����2���@C$�Mgc����ZN�e(�K̍�[�����=��㆐KZƩ�o��9�m���.�n@k�g=[л!��n��n�r�9˖��t����Րo�b��h\:ܹH�u����G_��}B�r�suzv�>���?Vf+�e����2p/܄7BF�p��we*��B'pۆ��n��{}��L �&C���<�}O>Q*y��!5�`�<}�԰���k@�{��Y���s�n�v�|.�)�O� �f��x������<�{튪f��D�-��Lm��.qW�z�C��q�n��
�
�|f|�S�M�O<���Gx,��1k��1��§�{�=U�_x߲_ϦX]LO� /�1΁�:�E����v�g��X����L�Y���ax�0��L���)Au0"��80<^U��9{�yf6/hz�;� ��GNg�bS� ����YG�KL@��~���a��v��w�m���g��D�ϗ()]%���ǡ��e����9З}C*K4<(Ǩv��y�{��ݷ��1 �yhײ���{�ך5�W�D��%�X2>��<��V���k� Ox& ��*�����:;�:�u��)�Oh�_3��
��w�����������c�bd2��Ů�x�\ڷ�&�{��)���ymx�w���j�1f��ksތ��#�߮�u�z��96�eR�@��4dS:��l<V�O=䓘57SN��se��{�v�����Ԗ���r	�N�]`m��y�=�]^'����!��d8|;I��E+v��`��+U�.�UnxָX���#7�}�q�'R�)��4p�n!���hbd����t����v���-1�%�8̬Yz�3> 9k�'�L��AޤJ�N̂�7/�A�a��53�%OE+�����T2�1�����e��ӷՈ�d��1r�s��JB2��� g�k��Us�H^��rr�*�y�^�������BP�P��^\]E�)p.[���Nz)A;��J���%Hm�!���v�sʞ���xCvx����_��ٟ%u,.�+��.	�-���"~���s��og��Oz�y�딵�1��vG,'B螠�49�Hq C∓�����/k^]0�7�ն����|�0k�����p����0�@����y%z�lmڮ�=yk{��[ &�]ǝ�.��ӣ���'<�>.P˸�"�]ۂ�u#W7/0�r��-��]Z��ʥE�_[
��XsP�2�v_�|̇4��)��ʸ�>�a9��sDA�//n�<n�ΡJƭo<��z&���o:�S�__$l������x���k4�
9�eQ�v�	�ٙ�B�<`�F��%����M��X�u�y�u���-+�խ�5Kީ���7x:���C�OQ�^k<��iFI�ä[wW�ot���'��-�����DTd�'���k JW/�b����vS�Y1\��u�ɾ����@���71r}=�]<.���QQ���M/��d�R��7᮪��\%U�;��9���g�i�����x�'A��f�vg^v��TD�Av �[��mgo.�5��>����E'.�c���Gԟ`��܌�ʈ�JJ���h֢���"�~y~Y�:�H��pc��'�e���\�}��gz[�3z!��}�ٌV
�.��᭤75J�YC)����5��6I�ʝF���;P-o�d����`��h=�Ǡ{1��M�g����pW���6Xlu����}'hk�z�֣[��>6=�q�u�J��{�kJ��̺QgK+�N�l�-{���A֌��rg+ӃN��Ϭ��t<m)p7LV���9��u2j�L	���w�g������]f��vb�x_�d@�'��B �U�(z"�����+ܸ\�>���` �a���M)�W��=^�ߎ���Բ��e��Ķ��ES�do*Ia����"�����.�|��o�͵�v��j���E���j�oK���-y��uG��M�4�4�b�{nep^)�}��cJ��c�:�ۻ��t���AWm�)�c����w�x�Ts��6`Ѳ��=	�gA[�6J�N1NЌ}B����pp��UJA��V;���n|6{Νx^U��P� ��az}�M�IwNm�ȥ_�>����ZB��s��2���#�p�g3�A}�)�Ax��v2�n�NەvQ���`�r��O�����_R���YKq�ϑ����_uM�}ic����ު�^)�h����tR=n�X�Q�LCt6�w��;�Z@mZ�S�x7�E�qܸ3{3�x}�<"��b�ta8,�=�X�\��2����F�^=�^י/��-r�u�J;���L:*B�C����T�
UT5��M8yrA��3֗]�3sw�^ﺼ�E��re!u]B�$��	*�h�*V�1*������]uC�Q�T��r�~���i~�7�\���yes�0���d����LV�e������k_FV:��E�>��+wz��7�@Tp�6�xd��t���9Y���}��1HI~gI.{2���ʉo7�|�<N��O�xi�*�9o�xem�E֪ʉ�ʫ��)_#�T�k��ѻ�x�����Z���yGa���dt�5��h��&��B�
��cX��:����y�7o���믃�N.�,����+T�8J�,�Rwb�{wv9�����+A׬kǲ�r����>���Xޙ�����8x�v�[X��T���R
�0��WXR�����\i-z���´�ŗ{�8���7�/�����{������I�h�-��8���3U�qTW�{5��xJ�l5���+wEN g+6l)��fk�ٔ�.�j�9m�2���Sh.,��Ⱥ�M�n���_U�i&�W�����9��(i�16��7B]u�B��ŘT{2�$���6��=�6=��]$I�M��u�����[�}�M�orxG-�b$� �[d�d�,��E��a�����T&n���d�w!�s��Jc��VH����_��\n!�y1.2��t�ëO�W�5�{���FP��v�8�x�Zç�󭓑�y}�t}v���uW�2���ޜ��"�qԽ�Բ�Nf��Ko=�D�4�<K�N�S�f�V6QW:d:` ����V��v+��ϕ�R�uȢse<W�nJ�|)qu]@�
�0�y�$�u���Z��s�/�s�kg�hZ5��@�'�_ee�b��J(��wt��gQ
9]sի�̂�������
� �9}��۶���{�8�Ty48�4�ۺ�vrg��=�9�3�2��țg���3v��)j��8)�oWފ�U�n�Z)>�:��X�罭��@��X�IIN�/v��t#J��L���J�㛅'���]��5R�˒�eH�U��I/�l��\�|	u5���|��V�ޝ}&�C�ejT��[��kN]f�He#g@�ul=2����d�����"9e��#����wo6��7/j*���鿅k�wd�&Q3�x�~�W�/E� �-E��Z��P�y�8֮�bY��;�Ѹes���Qw�k���õM�+IM��b�V�'jQ�<nV֑�mX}�j׿5,�]�"��\/!�iݛ�B�q'ݺ7G8�Z���t��װn�鄹]qq�(d�2����%����i���X慸�O[��������0�,MS�3�[ձ �)������s��ު}�[Pd��b�����)i�O��<І6��ƞ�J,�䬣]j��E^�j��w���,��q�Du�	�P�>�������0fh��Iċ�l]�J����.�rX�nĵ[�b�e�������ܝ�uj�`c�I��Z�
�N�z����,��e�h����#+���9�ͷp�;Ar���ؾ�_:r��\gq��S*��.����(�3�[t�ڎ��w�\YHY�w�btRW+N�1�|���rmb�;���B�L�\��Ϗn�5���,�����W]��#ŕ|��3���ԗd�u��vd��>�jX%@S���ά�;�3$���LP�O�
�T(PF[Q̹*(�1"��-*(T(��X��"��
�PF(��-TAP�Q��*1�PQX((���1�EA�`��UƬH��yh�*����xر��"���(�W,��(�$F*�PE�E(�+�Eie���ت!��h��-�,�.e\�E�`������Tb�4P�QV����
,UX���U�
�E�����e�b.e�2�/�3-�b�/�C��s���a�(*�3�̵m��Z�\1Ls#e�emj-��<�%��C)DR�6�X�E��ԩmKE��1A_<�*�R��Z��>\VdE��L|C��\�m�ʭ�*\���PW��I�mZ�n1��Qkm�~�=���|�x���8;��>�T��]G��\p�e�i��-�1��N�6K�������J�KK����Y���f��9<OQ��� ���斷aT�H3kƚЄ�#4ީt���a��!�jĭ~+r0��ݡ,ZH������u益;�vy�g��6Od�6m+uM�m��2xU��cj��]o�YS-z_ �^>pIԫע��q�7��4�� ̧�l�C�G�0�z���c�Xσ�̣{=`p��~��x�eg��+]*W)S�xІ�
��+�u���R��'�J�&Q�1�kY�xs���]�oV2��q$�ҮX
�( �ƀ�>�!I�' �OOt=����?gA������c���ѯC�O��(8�c����x-�	��l'�z]TY'xZ�wC�H�����勳�=�s9Nx]v)�K'E N�3�f�� �������]ң>�4����%�^��9�ց=��Uᓞz�����g���DP�)��
��>�*U���xXh�#�q�����-v�þ]Z��6�s����"~)E�� �0  ��9���q��T�]
�}�X�ϯ)�Q�m�,�|��<C�ax�0��L���`�K�dO^i{�h�`9[R�}�r��Z=�I67��Q�!��A�z(sE
�b�mx4�
ixt���/f߲^8���ۻ9D>���h����P�|㥸������
��u`=$ڸ���<,py��5O��@�ǳ{���7Z;F�xu
�:y�,��;#�>6O�w(K*�V�JA��t�m�N����	��~�	��/��{���=�{���U�$�S��>\��t�eW���G�V欕�2�<��8�W�V<A˜C���S����C�~����]���Yt��^[u��mp���}��@���������{�vtq �_EW���p�r#�eTx���o�QVn}nx��^:�E�!^P|�40����F������;F|�AWK�ᬇ�����ʷn�&ط]>�xdK��)x����z�T��澗���7�k�U3��Sܥ�$�>{'&�uݿD:���K��ze��w�����������G	Ѥ�k�%v��3RL���%OE+��~���,@�yD��>�w��b�p�6Zȕ�C,�S�Oi{�K��U���σQ`�������h���V?�m��7������`����l�g�̸��lU��[�ט2��R���A��
^$K^������G�1����_���0��Y�<ՇJ�Yj͍������KjJ
��zn�%�?]�Z���)��A�Wn^e���^�1r�T�ѽ���l��#��V�ǘ�E�4SW��V�\ݶB�9N�5�mp�������ג�eJx��p�pu�i�ѓ�A�MӁ�6�V��ht\��؝;i]����e9k�o*�"R����:�=2�>��΅� �]tH�����^^�/�zAv�A~y��*u=誥A���K���)pyN{��tE�%vY����{)��qƺ�^߅
76��Ss�=4�2�v��2s�#���Saǁp���O'7��.ߥg���e$ć)Q�V���Ň5a���.���d9���Hfʸ������}��כ�M���XhLDU��i��ܦ�%+��T/�m���t;�>S.U<��$v��gϋ��õ�lj<*�4D,D�ig��:<���ja���^y��A�6mn3��\�>B�a��"� d�v��J��wBR��U���}⅗�V�"���v��m�tǮ%������Ӵ�z`���eV}Q*J/��f�ʫ�HEs㚸`��V�yQ��Z��cZ�g���u�Ʋ��#7�N�!h=��`���Lh׫��)8{Tܖ}���uG���Hl�C���;�{�{s%M��`�t�����f2f�3��A@\~��B��[q�7�|H�|b�EZ�F�����Ug���<xR��^�id�O���T`ّ�اbZ�=ݴ@]�k�逾��yڻ�ji��̷
Ņro�[�^r�r����U9�_?�9��R���-.�y�va���Wi�ȗ�������8u�̗�େ�m6=�\| �����{�^ǃӼ��b����l�iEӉ��D�;��_q�3���4�*��PH�x�JB��c�K8;Ĭ+���u���]���1w����ˮ�Y6\mmO(4�E�7V�5�E28��(Xy��!龧�3��޿1�� ��g5Q��+��ub_���^O��dptt-�c>Fr�"�I�ɰ�o*����K�cj2��;�aϽ2�R�2��\����n��^��t�׼�rM����7
5(	$�L��;����!�}�P��">���l:�J~��u�����í�z��ty��$8���͎�.u�j�������a�l�L�؋����r�${֊GQ�29��Q"+����z�<-�Yl���Ck��{�M����o{�+y���,z�^�����y�2��\�P�Gx(M���T�;�	�E���V��!AաN(S=Z��|�m>�n�����1��2�\�,,Gy�лs�5{�-�L�}��=��+���x�5��o����Yo� )od�F��G��Ź�u���e� +�<9�����SR�wǶ�r�]�̵sh�����7s�>e�f����́�Ւ���S�^c�kd�Q�3I��	̵O-^;�A�y�vշ/9wM-NQ�=T��U�>��\9�H9y~z|$�U��+TĪS�&���=��u���[��l���KE�ֳ�0*����h��d�e�3�YgD�kՌWf���Z��9'K���˺7��	�˕�g���|Fٕ�dϟ@���>YD���_��Q��ߖv�L��GK��	U֍�O�xi�U.U&8'-��[�i�je;��>�ܯ:uؙ��*wN�.�<����������$fW�5�	�&	�mK�#xT���#s���c�n(6��Zn�j�Vϝ�U��c�2����󉇏V��P�v�R�H:�ur7�v��x|�-��chO`KEg����q:���)�k�3)�.P]����޷y��^;��*�J��W��;.��+�b��D��a�t(53%q��X���O`�5]��Y��oy��Mnʰ�J�#f�q$��r�V�@2p.��CbF�eq��]>Q�M�9eI�y�����C$Wt�g��yf����[RY�X�>�`q��T"�.�\����uyK���oR�ʈ��Xq�nu��R�s�]/�&�tA���c��N�fSqE�{�,��ŭ�c�*�0%�;��8h��Wr����8d˹�'�Ř���-�B;�X�ח�qnuu*8uh!�6����1��<�g������>c�{��.��r�M��zeX}E
a|O� �a�E��R�sO l�Bm{ȧ�:^=Z����۾��g���z����_l�5��"�ӡ���gҩR��6����/gy��u6Ώ��v�<�k��9�ʔ��p̪�`ALT�齢��[�_����;������D=}[��[�5���1�;%�:��%e`�.W��0��'3���N+�ǩ��u�Jn���:��H<�:V���Â�L�THz�	,���z���u��kn���լϽ���I9N";�LR���k,_���:`���/���E�l��lj�
h��Z��7l���K>(<N�m�O�}e���yt�pT˸�X�3i��^��M���ua�opw��J�UK��אyhL�#��gMf�P=S-��zt:��;���Ԋ����{���S�] �<5�C�zNF��V�׆�vj�3�Һ�_�ǗK{�}�cv�A匌��%pܾ�Ƿ�r�E��/�Ϧ��oj]0��ΈcX9��pe��l>��M�i
�7&�GyWwݛ;NkO_Z�bw3,�l�eӜD|z����.�G1�m��y����C5�����u��&�����ٽ�䷹J��r�����&���qw�\��%����(fa\�����z�=��;Xf�IjZ��;�5G�6N���'���9�l�X�2
�ܾ�}�|��������������\-;�k��ֽ;�r�~0U�f�Y���倹����g�؀G�}r�[������غ`�`��W�#
����U�BK��a���[P�[�Б��R5,���akjE��u�98ח��yJ���S>�G�_���:�4F�%u@�~U�x��Р�G���]�_�I�</k��lʨ�D6�`w;��K��i�Dpám�:+��k�Mw�����g=9C�ϓHq�Bxi�u7�2�R������zJ\�dpu, ����o��߼��j�3f�ez���=d5}1��.��ӣ��Ny�|2\���`�+N����8�L~�u�4z��F���&҂q48W��]e�5gǔgԻ/�`��c��-B�i�8���f��e�F0X���V9٦J�SXR�X�v�����:�5��8�kY���cy捼�AW}^�b#\2��Do$^�L���&%����5����lot�)�)��8���wX�Y�x��+�~�W�$���C�?���C��QW�����A�qr�S:�J��y�7��FU�7V�[��^��+�S؝q�Nޥ�v���bݭ<1�>�����
Z��w"3m��n8�ݸ�����7��}\�׾}�����\��t�#)�w���"��Q!P_`
�Ӥ�o�z�}��Y����rI�+)
�1c>�}C0��r2�DX�%[�}�-1��װY�E�[��fy�7)��F�)��=鞇j�.�Z�%�}��b����9�xkk��D+��������כ�ZLO�
���>{�P{N{-��̕7�����X�f2|\z��K�C�"��p����{,�X�zQ�[O��ǥ���ʸ�{�k�~��[^.���O��ˢ�.������l��f��9^�Ӥ�pY�	C�Ґ��-Sk9�^��c�wܫs�7]��[�vүA��dاu�����:�	�ϑ�i�U�޺6e��B�u����2׷g�PV:�*zuA�M(�b��ӯ���{r�G��bKk�=X��^跢/���e+��*���w܄0�z`p���K|k�l�I�~K��n��I:B�\��Pg?/=�{�c�'����LL��;�;���i��.�C#�����*��u<F��A7�Q�l�;��>�Ɲ�H
�У��>.q{!���y�{MO��<v����-���Aqo
��`���������p_::����9��l��A��/�ຉ�,R���5)[g!���D��l��¤�DJ�G�J����w>��H�J7^�oj�ۢ��+���S��u4iS�m�0�ͽ�n���#�����w����ή���p�`���T&��c�'E/�[��X\%�b�e�_
��^u@}����;llc���z[kD��|�h�d��.��.���(-up�g��-�o���P�_&{g��J%�y�����xK���0�
��\�,�o"��B�f��w��ړ:�f?7]���]���9�s�.�r�Ļ~=%Z��6�]�T����fǼ]���H�=BaB˨��FU�^YO��0��0Y=��fu��7ق�[��^��46��Z6}5P!�a���%�ps��v`�r�7�]%j�H��n-W��ޔ�����U���T�7�w}|@'�U��L�r��[����|F�U���.
{�N�BR�y�i��ڏj���XU�$��\i�K4ChvS�q��w&ǜm�ԯPlw�{M�/�w����vk���>oi��{%��0�	�*���ʶ|xۜ�]X�ł��R�'Ko��\{��G�AS��T�U�̝�F��wQua�w7��������h��ʷ%�!��4s�*۵+;q��f��� �/�9�]�P���[��#�V�e.�+n�D�DH�.����='8�Һ���;N��	1Y����q:��#��e=96)T���!�aZ��J�w4���4A����֪d�ۭ%bŀ�Xb�u�0�A���:�z}R[ո|�ւo&���S��ޝ����-R�RYFbZ/�$��r��F -�;��r��N�8��u���o������~�!��߃��ϒ��'I�K(v�)�Ϯ]�<�$:�J����,�q��ob��~����{Բ����
2�\�]W�,���fY���+h��]�'��>N��H�����;��~ۿo���*��Ny�^2�+g����"�ӡ�� 'a���y����ﲣ����.E4��)Z���9��U�?쉌ɖ�v�R��>���O��J�@�Pt��*p�c
����Ӕ_]y�W�����r�S߫&A�����ޯc͓f�\ck,J����}�PSF�S����y�t���>����U��,����Ml�sW�jv�6re(.�"Jq�8�b����3:l:��ɯ��j�kE�����n� ���<U�S��	=Z��SN�4qTp̓h��+�n��2Pu 3x��7j܄�����w3�������.<��)r�����:������ò�ׄiZ�_j��gc���b�\O_'�i�X��U{��;�yWP�������p��$e2�]��9o;5��ȫ}�3{8{�\gP߹����������8`1�-��w�}�Ļ�E2�h�y���]����6^�j�8법�竱�"�5gz�[���C����Te��{NLI�����6����3��'�9}�:M�u�Je�u��{Y-Wi[�vq�fp���3P�2�.*�F5��^��fc�kt%�=S��t�ܜ3���D楇��sԭw�'&-�g.wG4c|�p�����j�#,r��s�Bҽ�9P�Mu�m�oj�0��q���|'I�携��Xmk=�{�)>YwP���+��2�J�-[\�R�ݞ
b_G�`�]���y����2��n5��m
�b�ޕ�OoM�R��&�Oj��cq=�{�S�����e����e��][ۓ&��ieW>[Ǯ�:Y�Ig�h孮pk�\��F��'6���ٯ�2�̭o%��֨���غ���V���w2��ݚ�u�^!�6� [�q��	ҵ6�Ӊ�u�[�|�uB��7��Y��`%��Ӯ�2���������d7:�Qٲ���$��3 ��`�CN��qo�0%^M(d(�(�B0�5�F%v��7�����X�w�{(�7Ԝ����GzE��41����]�6JԱ��(d��!��<,u�T�){��	=���)�d��Ԩ�JR��º��S6Е�n��;����jyk{�=RNj��N�V�;��V�=b�\�u0S5sm�7�1�	C��G����|��W�y8���w��b�o�D�5�cx(�v)���H���v�����`u뺶Q�e
�Q�sz���l柺�����P	�����ݝn���dQ/ǭ�4�̋��/^B0�Q��G�[ڃ�&�'t)ҥ�3!���HN:�Vޒ�$�wAWE���|>��9[ר����yuqWYH�)�g]r�^�Fv3F�ԝ�ܣz1v����Ƥ�c�xFW��t�r�ө��Y������Hk��X�^Q[�Q8P�}��胙7
��ݺ�GS*�X���v��
��m�\���e��#]5�]S�b��ʙwҷj-JE�AzTYsm �,(�W�I��2���ue%�악͛o4��H2���)��v�H�wS:֞��jo�V��K��+q��a,�߷r�]��'n�S65O�T�b��W"
��떠�y�q�س�0�	]
�̼�g�Eq�#+HtLġ���p����q�+��g�V(7t��h<]��+YX��3DevB'u.�����9���wڥ�	��Y���i�ݝ�w3{;�����A�U(� ��Ke�Z5��Z�e�,����KkJ1��K�L�U�U����k�pjm�0�
�J*�(�ߜ\e�[Z-H�Z���+D��6��<K�[s0�4DU�-�2�A)*�IYG��*�P�h��P�(��/�UW�_)L���@Eb�f9Z�,�)*�4TƊX\k+Q(�c�\�Fڮe�[Q��x�,ģmYm��EQ�D����P��
ԮcsKk�fQ�-Vب�k�E��j�EaXQ�UJ%DbR�qp����%B�[XFؖĶ�甾R��X�51�R�հm-�%�ko�b�d�����̲�<�g�V-�UeUm�V�-�R֪�h9d�DE%�jR��V�n6Ū�m
B�լ���q)����?}�浼��}�}\��Jr˵��NWSX�)Q����	GA}B,��:*���/��L���5����s�k����b��y�1VV~�%��s�C�ϊV�$�{G�Z��yt�pT˸�e��U�{�cS��q�Y��7�7y��Fj��n��&��-	�gz8^��o(���(�x�/���^v֊K����u���AWH=�`����4he-[^�QZ���Vy�[)D�#1�\#����Y�Z|(��]r���u/���D����L�u:��"]H�6%��+��H136�,��d��/"��>̂�7/�A��p�S0o���X]��t�u=�I�G+�{�)���^R6Z��+�R倹�Oi{�K������1�|�C5�ϟs��o"0B$=��z!���p�Ch[(Y�0��wP_U�]	�~�J�XK�����mWf�E����`����ll<_�a�1e�j΅\>d��[�g���Ӣ��kb�@0��P��n�UȫD�(��)k.b#���XN��u֫�X@d�iy��]C�����ͺ���'4��7�l� ����ˋ_������8qn�rU��c榵R%H��f2�oE6��/ݸ�SfVX�2�гv�)X�V�*�X��a����t��	�ˤ���wS�0�����W؆�*��t��}c������%�If���ȖL�`�GQ�}o�TMP��â�A�B��\������__s��"��;�N���������+���� ]���~��X��.�ث�����^�7�&doVV3>��D����I�8�)�
��,9�q�.��x���~94��?]��fm�u�K�r`���Es&�%�M]���ʀ���O��
R/w�~�b�%-�,�a��[]�Q'[�b#��)r��D��I��>���E�J�X��S��<�y��?uo3Z&�^,��ք�0��"� Hx�jH��.��T�t�������2z�i}P�[������A�o<S܌�Ϫ"�!%[�r4kj���f��ݝ-L�}Z�LByw�/�(�O��4R~�`GՕ�vʹ�<4�ڸg�	-<��;{ˈ�+�τTz�7��L1�[~���}B���s���T������{g�]����� U~a޲��Zǂ����ͥ�ǥ���C����F&6��k�O����7(7R���茛&s;Sɳ�1ލJ��:*��¼mN/�^*��iֲ���u�8Q7uճ:�5h\�pp�[;1��i�X)E��������}Jl�J�r���������Z��U�&u5�tWba�����)eX�x;:�pf��l'|%v�ܲ����.��Fb�ean�-�j�����\:95Ne��:�n�ԇ_2sq:����zD�sv��+pZF���p��u�-���ת�b��̫^�=�8P7\+=��3�Gw4��;�z�z4���nJ�x�:^��dazl�
�k|�5�+F�藬�A^�JT��	��!9�A�3���ƽ��{Ey9�xL����{�k��	K���Y�,HI,M�HS�N����!�v����]X��	���j�S}rA#��ЇPCfR�4�]������wOm��F�ͷ�:�}��n�wH\��N�<�kW^����R�ț>FPv}P�D���N��.��n��d�/xD�u��͝�L-�bWF�քy�M�����I����g�Ю�B�g��'	a;O|1]��g���|�l��輝i��}.�����S�	�
(=�2��t,@t=[5�7�I���uc�`�v�ݮ�~N������dt�TI��V�T�껞q��3��M�m�3�xO���UC�L7�Yu�]ӯb��~��3z`�S�(Z�Π�ٳC�^�:g׸3�|4�Mt���o�e�T�O�Օ���E+�ԡ��i���%y_�����2� �P�7�g6\B�t��ve��WY����{�{���dI��0���:у�G}x��@l�)��v�ꅵ��r
2�EN�$��*����x���t�3~uC*�:�>�r�g����֣�$L��MZ��K�엏{����q��;:WۉJ��FϦ�/3ʥϓ��g� {�c�/w��:�l��6�>�Ui�
�����rl�j��}g��>Ә�P��kiDM)�󜎭}Y�
�Dy�MM7��C��{={n�s�g��6'��!�������7�3�l��)����vr_!�}�:��������)�G��iɲ���Ѻu��c@-_MK����Vx+�E��Ŀ�R���a�C:�r�
L�^��'��M���~�4����k�L�m齯��g�и�I��:0z@�{��B�ٿ<�o��+�{�s/r��Ȍ�J���\�J� i;Ĳ�:E1�q*e܄���Z)=���=�}^�,p�1�����|`�pghQ��<.�Lx�N�@��`�}N�N�0�w�z�H�}�c�>�/�v��({�b��d��X��ޖ�e筑��4)|8VP媭�~���X��,{gS��9�շ[�\��YW�������ۜ:����:��w����}f�:E�wy�V�_u ;�EmG_I�["�o%��g�#]����\���<�O�X�@��Х�_u�f���z��'K#��>{���1܏O�X�CE�[ji��yJצ!����JKxS�Ɋ�S��N<k�o�O��{��m��}|�
w��
���Ӓ�N�Q|;J��K��0ꗪ۸�>�Q�Z��v������z��\/��G�'�4|+������&*��1zzWq֊��?7ϝ�=ݗ��#�l��U4��J����q�&)j\ѱ�fy�g��֤�x��Aw�ڭo������7�=	���Ig�<H>�$��x�r���H:�����Gc�7�b�v0^��A]���k�����_*�@� N$gv+�+��h;���Y��ѿ]��'�0��F�����=����G!����`���<5�S�c�CG���{�L�yJd��wl2u;ͩ�/k2Z��QOv��9�L�?W�Pw���y,��/Rt�)����9��E��׷._�Em���i̻����\�|��v�Rq!�����m���9�(�0z=�*����0U�R�Jǡ���sU�R�� ]�J����|�����j�u[���֎:����Zn�P�M���n+�-��q�q�	� ����O\Ċ��M.�kjں4���/xn��Wf��U!!Φ��%uwh����@�eq'��V���NNy
���)��][aI�oRPԻ��'l)g.7��;>[�kʸ{y�D���z!�i+�B�V|�.��=V�ȝ(��K�u�96b��� �R�|��E('s�On=��_����׈��a�:�̷�$��u�2�^�2��YL-�$�u/��d��*{�eTU��D�<�\��;1�K�8n�/bޤ=ޛ���i�P�Ca_&�yI�q:,p�{02>�A�Z���IK�E��^��=����M��J�F�"��h�tZ5֜���<�������#��;��g�fNL��i�jU�)�ʘ����I<#1Q�J��U��<���Č��*�
n�a�2Z|�_�=�4�d��]`
\�!��EX��$�)�JWx����i��k�v��ٷ�W��`�3��1J~����":+�A}��Hϵ��*�K�ׯ'(�|��z�P�^��
�?z"�g�Z>3�B+�������+�� ��ϔ;bC�|�o1��d�i�>JP�^X����YOr2�Dz����NN�6���`Z ��2��zX��)F�=�vo��9�L8%ө-j֯�ٯ�꒔{��ZM�fJ�ΑV�45�vX�+�.S��� �&�a?+ŋ�'��n�����K�����{:1wRSk�v�$y��Gs�n���ںĜ�/��W=���r(;��/;3�1bUB!�~C֝R>�ظ:�zg������'���ٌW�GoM�,e�^�v��8;���W�e���X9�g�3�,��ۙ�~��P��_o9��+QLR\�6�WWy�|�\��;�^��t�8+�S����Q�96k�*�ܝ�S����ᯒ����d��ú_��Ѥ�]#��p�=���]z�>�{--���`7Z*}��9��Gq*��A鬩��kjyA�����
���U��:WN��{�ǲȯ�X�@ކ���t�}�:��q��qW���OnJ��&tk7��k❽�!	��PL���b*��R�;/�&��Cz`p���-dBOw��6gM�v��C��ҥz�.Z,��$9�I��ZB�k�3��'����$]#Ն���_���u4�g3�!�����x�]����X.�;�z-��~���6���X�a�§V��U��Ϸ�{���tw�4P�uB(�qd���t�ź��{*r^����~�em�%��;4{L]יĞ�`�٣S7��Zd���Yᤋ/Mt��Tn��8�c\�6k5�;�N�}n��8��U7�+>�M��zfDsV��Ӧ؁}��ԏ@GIl_hf�R��Z�5c]/��s��	�l��lt"�7eub����϶ΗՖK��_
�%���������Ւfu/dOHPv�P�~�W	�����i�����s�&�P�oʗqq<T毈�,y�K+`�a��
�Y�V��b�t����smS{7q���z��Q�o�z������cGNk��#�\����{�2�k��G6�Iz_b}��l`��+ah��4��c���s7�%|�B�����:TY�#�{��q�x�}S���ZP{����h
�������T����Xυ!��.�<]y�{��f�-8��_��}�{����߇Ba�j��<�\�������d��=���Sg��w覞��D�,��pW'��T��Ϟ;��hC�x&ث�g��=��z�RU��V�J�\>�rʃ���r�mc���k) �{%�P�N��g#�;5�x�4�ϩ��$��ʴ�]AV�.��ka��u04��3)��6)Cxr��U���~����_1��c/�f=�IѐX�R�:�pt)��+�����tj)���Z��Y��n:K�r��Pͫ5�ecA4*f%J��ۻ1��W$FOzǅ���d�`��%I^E܎^�V8����s୺�޾E�-�D�+�ϩnn�j�C���C��スV_�QC��L㳬ӏ��x+ju��q�ػ���ٟ�~��+J
�U=F�g�h�$�&ܰ�Pu��%��Iz��\�>�H#(c�R��ҍg��o�J��TN�eR��DV��?692z1��;H.'�3c��L�u�^~�d~��5��g)���(S
��v�Zi��B�h�ge޿uaceZh�`���<�{b��웜ʯ}��z��2�+g��Ƒ�������oGK�����@���3����ϭ�4��+^�bA9��T���)}K��u^���X�G�[���R���? �*wF�t7�*�Ln��V1�����C�OP���v9x����L& �Vn1�&R��`D/�G��K�4lW��Rf��4�NR����iڄ��~�_���xzV�=X:YG� �	�>�.����q�9�WIpw��b�E�:췫�|���B�����I��2�<���Y��JK>-]���D�J� <%��[D�F��[��.qXߕ�B}�oU	�a����0u\�q�{�p�H�]�J�f�u���5��x�Т�v�Σ�}2�Y}�1����Y��,ʽ�78��I�(�v��qd����o�<�f�<��qU���I�hΗ^WO]�h�L.@�})g=���:��H����SW:���&rmY��޸��5�W[WU�F�"�lg�,�q%ڏ�)�LCՏ(��>�42G��p���] ǆ�e?�����qM��_K�U/�Z�~��R�j�B�=��׷/����s�R����ל宆s�7����߫�D4hi���\����J���\0����s�2
���0jA�A�勽df����w�����z���qP7J�CW�,�˖�����R���;^ؤN3��Q�m�K��8E�0Wq�z��%&�,V
\]#l���w��XȬ8��G��O0\�k��	�r���n������N���<B���p�|/w#\���on7���N�EW�}v�A�'}Ԡ������D�(������,x���m-��tخ.�����Bv�@��Q!�|�NS��,.k�B}qk��f�Д�)�����or������%����(1� ���Y�O�w�^����Ͼݙԧ|�8��&�z8��F��ѵ�ߙG7~rݿn����\6��߳�$�	'�@�$���$�	'� IKH@��B����$��H@��B���IO��$ I?�H@�xB��$�	%�$ I?HB��@�$����$��$�	'��$ I?�	!I��$���$��b��L����W�WN� � ���fO� Ē����j��D*V�
hҭ�hY��ZefUJ�$M�� ЉMl�hխBi��T���e��#Y$� E�@[m�"�*�%-m�o��ZZ��b5Sai�l�Z�E��m�Z[*��ղK&ڌ�K, �f��X��[&[E��E��c-�����kMU��iS6{��5����h��ʛ3J��-�(�fV�kY�jkZX�I6�iJ������kK���*`�Z�m����mdUd�g��e�k����5���   '^ h=�mqD�U��(h����U�;�hQf�n�F���h*�kY�%JSKv;��a@.�]��R��f�j�k@��f��&�em��  ��e@-I����Ud�t�t�l6�g�W9n��V�5���ҝi�ZFm��S���4(���֖t�Р��ͥU�,��L�k����ͭ�   n�h�@(P��U�(P�@ 
&w�x P
(P�w�/  ��A�{nB�
 �B�z��(t�B���t( 
�hP���xR�[a���]�*Rk;��[j�5��mDU�-�l��b��Y�  ׋�m���n��
���uˀQJ
�u�v�ëag.�4�p�.���`-�ӧ�ղ�BT�l�j�4Қպ:�j�Cln�둦�VZ�8D��%��x  	�����J� �i�YZi������

͵�uF�M5Uܮ�m��bakVڀ�Ci�PӶ�X(l�ή�v�eZ���۸[���B	Cf�[�ӷ� �o6�ڥ���@Puh;�P�V�t45�Z��ҩi-�;u�
�J٦a���:�pQ� ��q�)Zi�GMSV��Mm3
SlmE�  6� 4Pf�ݻ
R�m:���;��P*�ge�P� Z���6��n����Si˅�4,&UmgL�AZ.v�#ưݻ�ifJ�h<  .�m�T(l9�t
�K hwk� �1ZP5�� Q�9P��
�9� ��m� ���B���X�l�K�U��x  u�/cTN���ۊ�w�7� �L

��m��Puӊ :�C��e�
�����
�%I�M�^   ��(� �p cP v�nQ�s�T��`UPvpP(��n �SS0 �. � �ƃ*J�4 2��a%)P  �O�R���0���U�  E<�h4  �PSb�SH�1f)dB 4�gZ��Rx3�l�f&Cr�*@DI��n3��_��t�Z����$�	'�wG���$�$�BC�HIO��$�Ԅ��$I! ����?�����Oʴ�{W_ӕ�0,O�%�P���[���ڸ\���V��,��(�b�Z���e�V�oU�2��*�҈Ҵ`[���46�;ɛl�r�u��YM�7xb��Ç� Ý7�K�8o�J8�s$�m�ZNQ0�U+��o��hw=�*Q���O z��?�LX��.R*�̢^Q,�3,�E�J�v���f!N�kp��FЛd����Q�[>��9b���!�hfS)%������f4���C����.L���O2�('�NV���2 ���p�����N�����/p����ū�6�q����D[d�Pnf���|��!�1�T1�W��Mk�;��"�q"*hk�5cKC�o+t���c71�6�:*�3Y�ZF
r�K]̦�z���X*�`�X���Ն��)�T�X%Y8op�M�eMŹC\A�D�;u6
6��{�f�w&U�"�e	{z
9�P1�f�S�U�Q�����ذ�,e�%8�5D��`U.��5�H¬t��m�	�ʲJ��[��lJu{�[IJ��KQ�d��Y�]���!��*u��G.��ЩJ��yh�����1	 hMn;�0Йr�X��L ��H̻�Z�z�ژu��؃N�1�ƀj��Z�cSC�	F�ٔ,S�'���-�L[@�ӕe���e�������ثk���3���&8i�:�P>� ��P�1hU�2��eJ7Bݍ�hKsG��D4�]{#�P�p������Yu��P����):���U�^Lr3�
"������Sib�XY��h4p�1-2GF�;.�u�؂�g`��iV}���Vfn
�#u4*�:m=����1�PZs��-�ͣf�:c�z�e���n�mj�@c�".%f�Ǒ+bzee�ܫ04���qڒ��hW̭��m8�&���.�3����(�cq/�tyyk���$�5d���Zj�-RM�˩%�l�����҅ͫ8N��=3U�0d��u"ݳhA�[vq�1�&�dҦX�M�-��Vi��j�w,Z�Ff0�-�j�4k�k�e��X��;u������w
��K6��n���>i�m�+Ae��he�-��:@�v���d��\��t$��Q׌��r�oc��+�ee�z��QҶ��3hb-<8�Ms��]��ԁ�'p�\+F�@�2r��Ac*����mLUa�T��-_m:v�9��@hz�olm��pJ��8F��Mͥ�1�x��Ãs4�5�ɴU:LQ6��u2�%�/N�pE�m��R7N�����u���&^,��=��+5��j��}o2^����$K]�H�{{�\��i���wv��#��H-m�aeк��8�ʴ0hRʻ�Ǳ=�)vn��$f*6���˛"8Ԭ������	m�q'��9�Im��K[7%+���N�uI��KZYW���\��8��
A#�a���.b�\:;oS�]��HR!��&��0�bVQZ��!���[�e:�Tq�����罇�Ӕ��g�t�vD�h�Q�L�*i�{gh4ũ:o5�ۜt|w7�=᭟cLL�d��ǌL���Պ!ꕅ�j�QYL�)�H��<��{�Er����"1F-��x�bT�Csr����m�%T��mnaZ1��T
`�u�WKl"�ò
�j����D虸]&���X��Yx���h$3��t"4Nw�
���d�kc�[�k-�ң��f�Q���P%�Z5�n��1]�3j�Xئ�"0R2�aִ��/Y��"�*�]=Xo^`���j2��X�e�����5��-L­j��U'E�gѭ�g1X�)HPX����!;�k�i��E:�n��2D�����9�d�r�Nx��B֚�Rܵ�3����t�a�I�f!4�ѩp�/k-�6��j�[א�(�ծ	5���31U���6��g�	R˔2CR
�aO���P�4sEb��4Ep}ӓY�Q=0՗nGQ��`���۵�Q�U���a=5�Yh�C$���ɶ����b@��d����p���'�����c�v�"v俢�c�Nn��!]�+��Ec�;`��c%2�k����5���vE�$�KXG5��w`s�8��sv ��i2�Q�['D�5�ܥ�W��{͹ز��R�nΙ{{���-��W�ڠ�z�F�
�A�ɡR:&"N�ȝޘ�,�E�p^�N�-�+l��f��!&e� X5��B�&�_Ma�Mg �K��$��Vˑ+n�%WoL���*Z��+`���T
�d��[6���tLpn1�(���4��x]Y�&����w,MZ�j�$�Aom@�ŷ ͼ�f��7�T��9w 5�l���fF��2����e�/��l�ۡ��E�N: XW|'@y�b�Oy�_�[t���#BU���{��["�}{����2X� BKѓ)�y�B7�am�V2cdM%e�a}2RP�m��¤FЩ�@U����X�d�Sq�b+� ܢj�^� ��X��I���R{v��@P�JR���v��d��$P2�K�,����"no6�7ĥ�9hQ7��sdb��p-֠�Β����|��J�dܣA�v���L��g%fpIYj=�0�o磐� ��ڤ���>E�wܖ��q&me=F���V�Uϋٱ;��ώ�,kX�b�>o+.���1���];Ȧ�+SS+>wC7-i�A
3XXn�
��Ix�շ�|nゖI�fd;�ԁ˟*�7D*�Hg�D'�*�<�t]���K�Y��7H�Qi?n#Z.�5L��XU�o/Xy�BZn�#�ۭ���ɱ�W��.�"3E\'f����R���n[���H�u
r^�X��Ǧ+9��iwlʒ�ҫ��!���n �R�&�6XK!�� �Z����r�A���,I�s�/E��0���8�$m�g0\�U�Z��֪Qȣ�Č��5�V�RS��Ƌ6�EB�n6�z�Gh�j���FnX͹���Ɠi*`*�Ν�Kn��xv�u��:�t�8��a۩��h�K`zo\�&Ki �:5�ml7xR�d���y �/PE���U+	�lK�n�n)��T{p�-�:�،@nP����P�s�/�.�؛Bk��{JC��cP�Z�I�*������
tࣗ�6�S�m�I�F�5���Ɔ�����M	U��b�VNLY�DlL�.�6�@�W�Һ -���<�]�����Ą�8�iMaq�x��P�ddb�=�ܑ�J0f�������P-/Őd�h%�jׅ����R��j�j�e��E�(̻A3���gJu�+�����&�<P��w�hX|u��1	s<[t��;C+�I�s#���dl�b-�_aBի�.Vc�.l:�Qt�����]�Ei%�nO�t���є[	�kA����;����	�ē�eYt�o* g4�U7�kY�:ԃ�ꑛ�i���$�SO��3�9ڸC�k�4>ل��6�%&(��n�㺵��ɩe1�p������:��22�.��V�tX	t�-<��"4��bR"a�J�2�QB���в�=�R��i�2�饗{��"�dkscB:��I��b�7[r)*VkU-�m���}���>~x��'#���?8m)a��$k��3Jf�x�U��jA�ii�cIKt�h�o�
��{��FLj�YM�-�.��L�">v)��������4U����P�k)�+N�-1O�e�[Z\%���z�'���E��R��m-7��e��7����[��Y$Z��ˌ�L�ږ(Bs]f�J����Z&I����q�	ON�7�X�c����"s��g	8qZpb? ���w{{�J�{�Y�H�����m4�):�W�k7�������M/+$���;Qr��FH�0�Rz��vU"�`�3�<x�@��tL��1&�N�x�����
�?!�s�o]e��^�(�3#�ފI�OpV<�1R�h|sX�S�XFB�����ՓA�"<]ÑXߊFn����q�&�r^PE�Jm��QiU�1�X�]g��YV1��iIr��L��qVD���62N���V��1�aX&�[Hз�TF��F�bR�M-f���jk9wXt�/,�zVT�T�'34�.S8��6n���	(FԶ6� �5��Y�V��-��+��iܫn쇦�����kq�-��@3/��<�u鷑�i/X@B���(��A�L�I�®\l����݌���L��LE�뷎�T˚V��u�B���[u(�l܍7GmɐP�].�R�f��¤���;�E�����x,}2��."��	i=��Sm1+m�Z��&6��l��٧���e\��ݶ
�,��h[b�s+�&ԭM�u�чA�)ne�(�L�̙��55"�Uj�ӂ`�R���Qۃ31��l�I�مԳ���w��ܥ��I)[�#pP�^*��8�]b���`�ͫ�J-V���6����D��du��`,�(h�$��)`K�H ��th"��6�����7`�;����,J����]f�kth���� �G�Pk|_"7!��;ú�~ԴLG��I2/+�
B�j��|M*Z�w�)"M��c׷�Y��T��+.�f��'d�z�h��s`��K��x�fX�;ɂ�E�6�G0!�-AGYb�)�ŭ$QHd3o
b�Z����W�G�����G5LKl]c:��5�dۃdW���
��5�=1+��2��w5�X�jͫ�a�8�j��L	�&�Y� +1m�s+���;Y�kG�b,�s�J���7�y`,E���.�"�)Pn���yǵ�6�R�!Zv�э��+M�g2jD�� �lQ��+�G�âQW����k��ٳ]�O~�%݈ 9����V�Tj�g]+F�8��c"��R,.�pX�>l%Ssw+1�{Wm��
"�͗vw-]��A�kofVf�2�yWS�5���A�5�nb��-inA�A������a��D�)c+�-�Li9CU�+Z�����Y.���^��4���ʂ�d�^��S��R&a��'���� @�TP[b�֛U�`4�,20\fA��fJ#,�� ,TD4�C!��6����!Ue�7J����/^Q�6�V����JTj�[H���#.dX�'�絥�j��/a�0[�a�-eֱn����Xu���v�<�k]���rԥ)�h��n��,shBՄ��#��Ϯ9�)n��B��vnP�!��dR�yA�y�f-��rkiAՙVB�$ڹ���46Ê�Y6�m��e܆�#vٸjV�ʛC\�+V���B���^Y�ͪe���q����R�D�F���̈́��
צ�`��u����R]YW�[ǄiG�8`�pZ�3+C�%[��*��ݨ�5��Ќn!��Q�hY(�6J-�f�Ђ8�Mȯ^�DIF������t��ęF� L�v���iaM	�Y�h6�±b� ���C2��c.�jP*����:�i�R��hƸ�,r(oq���
���XU�&�V�}E3�n[�8�e�-fS���M�W̵��d�m�V���#%�b��N�T!y�r\+˸�7��LU��Gqԏ��l-3�N��sP�u�T�)R��X)��n���tI�$��kihB��:����.�ٌ�Z"n��o�� ��CKA�4�*'�Z5�k0g�,� w6�nl��ʨq;��|j�a+oA��i��n3��ۈ���f�$��\��H3F��p��� ��g�tv���)3�֛��`����M$�5�ʖ�{��*�m�}����njcs@b�WBҶk��#�~;&��qE�Љf�@9y!'z�C�X�,�QZ
�*�TP�2�G�kH���P����WKm�Gy%�E�Y���]�X��J����[f+ʑ��حK&c��S͐�Wv�I��1�F�:t,��S@	��"τ��p4�4%bκz�'jTvA�K̽	
��9�c�,U��,�T�f��cV���ұd�I�x
x*��4Ԭ���r�(�{��-�n����O�1����V13k��f�BA:��P��t6��V��AV�a�cef���G6o7��, ��{@q��s����A[+4P���r�Ք��R%1ͧ��Ժ��ӊb6�
���Y���wF���i��!��`��]��Gwx��ۑ��Tv+l��T��:�Yy��Ti�xv]���
I	y�	�]�ɦ�:�t֪�����enҡ� ��'��b�K-[�i[�)�R����M��{��-��f��Z��^ 5;��OI]�2ŚFW�R&��3�݁co6'�Y��S��������t鍧�� nKGQl��`u+��H�l��g,"�����o�7)s��.��R��[䔓�%���Yt��i�;�l��K�<�������P��2k�{��0�V%^:+���Y:��,��
ւ�b`JŐ��,��KZkF���rXs~{���û�E8H��!�v��H���S�lTǙM=�WV���1��i
Ifbh����$4��"�c�:�{Y!����r�`���'1+"*N��,^3^]�`h�/"���u�*���h!�3j4f3)�ƥ�����ΔMH3*Y4�Ȫ"ov
�VTT�7��Y0]Jw�S�w�i���R�N���j�1�e�71R����2̖o�[m;⬴��CP)��J(4�"�3o,+���l��vK�űֺ�`��V��m-�v��flL�W�#���W��� �펓�id:���4i���|����]C����z)Φ&�^�`Ylc���05���6Pu�h
�I��d�����K�Lڦ�>��ư=�;x�Y3�-��+��*_�g�M0K��^m4�U!�U��;�΄K��dP}�Ͷ�S�.�z�b�B���֑�7sǰ�(�@�۩�9�n���I��M�.���
�J�y�әu��Ʀ��v�=��p��38����M�8�k(��)Ս�e{O�T��B����X���-cخEzejk)�k4Bx�u��b��XK��:�'b�-k��Da--��E:�(2h��-�8X��'n7ZJ�����M�Z�^YgۣF�@]��k������j�:%ή���g�����U���Uj��ڽ��<���V�P�H��V!QYv�;Giuk҄���B�i�ڷ,���V���S_'/��]�fI9�/b脷''���'�*֏!��BQ�����;�or�0�w�M��y�t�t�:
�$L�e���jE�V�Y�ȞT�Xݸ��w�����@��qB^q�S��O(n��D��z�MԌ]�tl-��ȱ��-�����!�� ���� �p�&����L?:��/fuǧ,9�B��5�����f�t��M�L"%2ogR��#�����5���J�q��ѻg��xqae���x;�^��L!b�r�U�dsc�R�
i؏X�������4旎���8WNBS��:�d�y&�vcp�BGSJ�J����`ݐ�{��:Ձ�)��H����u���+ϲV0+��f��Vr���w��/�	fȥ�q�ڨS]ەJ��h�V���:Ь�ڴ�o;P�;��]�T�rr�����U�m���#i�Τr[�DڊĶ�d�AE�;�u �K��= 7�,B.��~<<^��s�Ȍ����P=z�=���`��I�nsݮ泘���6N�٧;h�w|��2w?͏�}Y����.�|xnvNA����;$g<�nmz��K����)�'�5#�!X�K
��D�U�U9�q֜�MùV^�kbk�{8��oG�P]���j�|]���m�uP��������lyL�x_���>+nl�w�1N����z~��[�Yn5�v��hzf�ұn�{��xRXinn�޶+���i^ۘ�.��:Q;:WbW{/��_�/�׵kuzg�v���O[�J��Օ��4t�܏%љ #h[���k�=���ڹ��'���
8ғ,��F;1�����N� j��,�'�¾��i��s:�5x�ü�*8+ZlS��v��C{x�i�]�|e��&���c7����^�i0���v�9znrκ�bun��91�w4FY���ٻ�w��oS$�a����n���b�F��~A�R趤����*�E�F]��EvźA����S3�E�Y.�^v�0s������w �s�ʾ����Qw�����r����+,V�r�V ��"�9<�Q�!d3[G�,�Ѣu+�eMK���m�ٯ�UQ�^���)�����D��3�d�orǏS�h��{R�]C)����Z¡�����: ���ˇ;邸��	4dW�p����h_5F��t����gn�ڞ�{Y7���yDF�)�@M��I�CR�ɝ��u��c\�JJ-�@o��ޡ�yl]�p.�)������θ)�WfĶ��l�St�]�fu5����  N7R�C��e�sWG�>�(;ِ�o��g|��5W�׶���w*Q�c>g,�m�_j.r�(��n�� {�R �}n:{�w�d�e�p�'zޤj�bV.#}��˩]���o-�z���"��=���o��m>�OW��ۿnƮ�}r�3d���wU�֫b{��+ïr�L�둭d��n�E��g��w(�A��	� ��y��e�,w+/�03�{�0�����O����f<���]p�eN�q��5.�Y��W�濇fi�
J�xoo7��PՔ����h�	�~.=��"QE��GԼ����鄋��O�jp_/QUC5j��KI>�����l��T�e|�Q�<@�Ie]cK���]+��,ĞS��2�g�ii�ډ����e��Ӝ�U鴨|4h?'���M�6�)����|4kewp9΢�/�y����Ǹ4��`Gۗ�:���G�``{��QY]���!�ۍ�n��hki^�U�$�P��Y8	Y%�A�)ô#�M�.O=��kxQѾy/���� 朹p��y8=��yf�+V�!3pv�խ��of嬋SVn�r�A��!��L^����>�z�7�b'��&|X]�</;c#d<\K���&V6^�q9���	'�}wMWʆ%�V�!���<:�A��=���Y]�����ቆ�k��>� �gT�B�����+U��S��8u١���輔ņ�;ݓ���+VM�/X���,o;|���4��6��`N�g��`:`�D�]n�y����u�*@Z}��M�<�
nx'��̻�pSJ��J������h=	6xn (+޼ن�t�l�@fЛ:�r�'�D�Z<om��D�
�n2`�u��(3�k�wgg�I��#AO��<��5��v��n�9ɛUv�t�:�(�����[!	k�ݖ_�Q�x�����[,�>���������C�(�wz�dܗ֯DF3�s���SOV2�y���v4*�H��d��z5�AƳ{�Υ��/@��K}̜�	�f�衇R}Gn3k/kd�]��*Aen���\��*1���`6���<H¡@����0�0̥��T���A�O}�deY"��S��;o�䭏y���*b���^(ivZo��ޜ�p�A�Ŗo����a��u�X��1��Z=�xG�{V���L�����;_p9/B���,w]����l�mn���4�Rd�4Ov>/#�i4Сf;�a���Po>�r�������"C���s�!��X�"l�"1�8=H�l�M%5@cOA��ox�Rؼ�{hZy������px�n���U�kNa���ܚ;djÙ2[k����"z�*��Ƈ���Q.5��{�cS����	\���s�5�Cr"�vC �讕�5W/{�-��
u��ZUO;r�X��s=���-�e���O&7{+Pv�9Kk��.�wC�Pa�{�lڠ��0B;`y�ڹ�-[k1-t�����T9�(��)�x*��6�o�ը{(��7{ʵ���{I��tM�:��5l�I�|��:����&9��{x;��O#z�^T�'�rP��B�i�f�b�:��5�|,�-N:6T��׏�d�w%�7J�2v�N�ݹ��
GB��o��p��u��H񠃶�7�ʙ�wI!��qZ���XMv��:��N��0T�Xd����;<^�a���>��W6�$]���Nl�mV�!?��_\�N��n^3Uk�,�G-	�{�R5�Qc�n�#�E1�9O�'�45��p�-0���)�TAK��K�F@�l��#�@n����Ze���S�^�s��Xۚ�<D�����6�[E����w��΢������5�I��f��P���c`:z��C�*��v�5&V ����r�j�cс`�.�E�E$2�(-��2!��]W/b�:�e͑�V�Xqٛl
*�@���qsp�]irkK��#ǒ�:4/��>o�Zω��T�j��k!���R�n1����{{Ou(�r7�j�{z�94�cc9�(�� sn�lޭ�̄�tk�q]R\��{;�ϼy�����L[$y�Ě6�j�T��}v��}��0М��00����B:b��iܹ­
���"���6r�;��7��y�Y�gM�6��w-������(\�U���d��{�.xxPoi�7Bه�gi0mG<�_t9p�=�#<�D��3�NP���G>�؝�J]���v���=��z�g�>�$à��N�dW��[�x Ev�"�R�c����{ػ^.���s	���:�6���:�
7LR�@��	�֛�9�]=2�������B9ҥJ��9�n405x{I����v:�v=�-���l$���<nT/Psr�݅-_�U*Ow
ҸNw'���t���t�;Gi��p�*��eߒ��xV+E���S�A�i1�v�r^J���1á 4�5�.�a�7_h��xތ�AU�lc.�ň�Z�]g"��u��1'�/�і�J���&�Y�tA�{��&�ْCOo����ZU-3����|;���|F�{&[}�8���$�ǔ&R&��6�=�!�!ǈ�X���*�K':e�2p춁�4r),:Dŋ@Ss�'��$�y1��O%��~��$ֹ��8i�J�\��u�wL�Y��t���k-�Z�ɉ��gM˚��2ws��it�Z����rÙ]���L7�t�g��q
|�`�O��4to��=哚{P���V�H!�6�^�ب����pB.�e!��2�"��,`loS�V2�+6h���>�R�^Ml�T~4Ϋq���`�%'zN�;2�Z�f��̱��9���w�o�y)4�z�3C�S���᝚���X8�j�ʈ�5>Y��'ԕ�K�2"6[W3q.�(:V��Q��V[k������r�K���vf����Gj��Ư�h|n�V|��;�O9�`	peQz�n��F�z��ŒW��5!��Ҳ�g��P�����)���9�׹�;�Z�<F!z��>�f��&����\;rnM�\޼���ç�>�X{�_<5+V��6��h��;�a�Ye2�]�ǁ���~Sg"�����v��݁zw|w���xg���=���F�5֮TTx���ѡ�;���(�Q��.�e!�X嘞U����
�Ǆ�
aXȻa6/W<`f�Cb�<��f�h�9ڛ�n,�z\t_c��������]�=3}�B�]�kZ�d�6�+x�{��+mtt��������&F5
�PK3)���C+h��gv�}�$ү���>�ϫ���9��D[O;��{k���9E�,����#�,t���ckQ�ɳU��rd�Gd �Ѫ��Ǔ�pJX��XKM�]7��W"ni}�KP\O�E���.��-���
c'�s5�$#��G�TȤ+.c���s'r��x�����.�|L�]� ���['e��'�Z�c����e�n;�&gi��L���X<��հ{r��Zx��zf#�z,�o��ۂ���F���!�2��W.�b,��`�x�yi;��9X#��0E�k�q�p�H���$��۟	uۥQ�]�]��*,��0wT*�6��o�$�����;�5r������-���00v�V�3��\p��HܶD�Ẓ������fw3+��6�;�и����Q\�ndv�p��-^��hޮ�=J����ldV�7^jye���ŗIr��3s9CQl^k�8;3�>�Qh,���a=d�oc4�楷.�U��������9ѥϸ��i\sH�Ju��%(U�X++	��"b�Y��d�V�kܨ�u3͌1y���ك8$�N�ۡWX4G���������z��U��L�)�s��A�V���
5t�=�W�4��[���e]t9O�ow1���ۍ�j��B��F�8�K)�B��/o
�p�s6F%
XCemh���<z:��ۓ��3�vc��ܧ�~6�"=u����N�oj2i��1��3�:� Q�9��əj��{��K�
�3��}��*�0)*W^��C��V�g��ث,�&�Lɺ���k�8��1ڻN�A��wo�N�Q�����(�;Bv^�İPɊXs�G*���>��+���s|��7���*@�8S͸vѾ]��Nw�.�Z���3��Vx�"e&h�4����zS�q�M�]J�7٘�ƭZ�2f�miT�i���)�3�-ux*����w�ȴ��� ���o��L3��T��<)�IȎjK��L�I����4���6�)���ŐQd��y�Oi��ix�ѥ�_��|4�����E�1:-5��դ�	F���୽S)K�{Z��F,9�e�Ox<T��J�*���U�X� l\"Q���֎�w|�Z/�="0���'��b��}3Ft��ǰXj!a��?S��!B��ܝ�t�Wg��a�Q_���C.���8��v]#����Xu��:��_&).P�V.{|+8��rQB����a�*�q�͑><W�o_|	�e'�0mk�ґwU�yp��=/5i�����Wy�e/�S��35
U���C{t�Uj�Y
WsM#���o�`|z��m�5��'��u ;+HIw��p��:�-��l�O}�[��٪%ձ���b��ѭz���_N5_G�H��}X���Z���r�y�w.�B��ܨ�Ӑ�SrP��aE�y{��gL�5r<0x�wǴWb�F��9�㕵
e#3�o�ܳ�T�'FS��^~Zv���S�E%���1q�t�V<"�)��ҷ/��T�����蓈�7�0�0�yR@�4NĻNi�s[��Wd,�^ޣ`ڭ"�Z�#�Ow�}�G٨j�x9n>��Z��:�lԍ�x�HTyO�������Mv�iԨ���t�[{J�fSk����L����%��w<[d��8eX���T��t�g�'WM��vqYǱ��]`�>/a=}q蹻�[.��\���\���ץ�����m�]�K���6�}��D��HH IO��c�~h�=?�YI9"�{Eg���w�0����`����y����jظn������2�"����[���ˏ{Z�q%dh�Z�����MJ��G!C:�����q(㨐���dW�}d@I~;�j���F{|t��ށ��{�-������g�^z� Ew�A��ZY�������O�\D��4S3jfL�k+��8Ȧ.;�Na��y���ޑ{�h:F嬳'm]��5foi�K�X*@:}����x i��ɶ�U�����i4!�q��T8�[�3X�Y���i���l"��_nE�GC8<�^:�ؠ1H�w<�����
�M���5�"4��
e��h�>�>�=�[��ŗ�=�Y!ȯ6�{��$f������|�8��u��^ռW��8Z��J��ӢP��] �3�(M7�v3^���xd��9�M�g<"v%Wk���[O�P�`.��'o�����g��g��RGz���Vq����!ҞpǷ���Uo��֌1��\#~w���,U��ҷ�a�TA�P�k�=|��Wk^�5f:�m��mn,��.��.G�w+4�ć)�BT>Aج,(&2����-�fܤ��V=M)���Gy��*"�����S�aJŖ �ݫ�}��aΥ�u��$�lkYs����Ű\�{4�u�&r�o�`�W{5���i���u�8_`|7|=�>�����1�u<��+�=םw���:R|��2�Ǒe:���A�d�q��j�*�f��tP�!Fv���߉"˺KOjv�].��cj�������qC�#㞺M��t�L������Zkp��5��`���[���� 2
���q��
���K;0��D�y�S���ZlI�VPZ7�x�ݦ��n��2��.�z]5w���O8�;4]X!N�11;8%*6¾���#kx,�# >i�� �U�u)����iE<�a���������x�AD ګ��:��[��p����)�X.�+��4Qo���l�m>-.q)��56�J�=���T�)&Ju�T�|���</W��)4_[�ȬT�������q�YM�9��p�p5�n���tV����
��93��cxӜp��ѹ=g���4�%��e&�Q�jr^ec����m8	���w�-�;6��n>���V;r����p78L������d����i��i���m�x2W������ ����.!���^�uMNR�N.�[i@�o�ЗJ�I�m$�g4E^�	;�]<xu[�r&�=�6�$�m�>�5���@�M���t��C�b�b=g�	a<�L���;��"�A����'^s3�13�6��?x��Ni�3��)N�h���p� 	�2���v�6�u�Ku��SVP�A��� ��%�F��:5�qL������J8+��͗��i9�Jm>��^c��S�d�n�J����<ns����t:�Ѹ���1Gw}}����eN���}2``D&x�4:Iս�nv`CyA�J�s�~7�@�݇��.�uZTG:�9�<Y�x-A�!�0�R�Q�S4vE��6>0w^�!���R�v����c�r������"�r���NW�'��S����-f�!FN��#��7'ӊ�wK8.�ʳ{-a"��yB�to�X*<H�V崷: �F��+V�D K`�}ݞ����˞�]�(ϨǀQp���%�H��Vn�;�;y�^�Ya�y�	d�6	��u}�P�0�ܸM؂�����c��r�`��>H��hJ��Q.U�c���{G>��c[��)�֞��i��3]d���p��:B9��c��΀�<�މ��ھ5�]��1e|p*��n���T��kZ��9�| y�btV�`�՝p�a���ن�[�eWkd�x�7g ��
}j�X�!�g��`��}�e��2;à�`��Zy��_GV�����$e+�ƟXh�5��G��Ԋ].�>�WO�r�{�^�����tqe�D�rU�M�fJZ�T�c���(�M�9Yt�ʵ/��򫬒�N��o�eD_oB��T2��I'sNQ�&�$��>�o��^�P E���o��e���>���	ږ-|dt���Gd���+|��Tp��Z������N�&�eVtx�Qy��%�:���T�.���ٞ>#"�ۗ�H}2�Y�p-~{p�El9MSYe=Gh�b�E�8AX��ih.�`�G,��AA��i::���KNm��1�b��.^�va-gb�-�vQ�a�ڤU^ӐV&�o���!�VV�n���e��<�p�;.���,-��O^�F0qJM@%�Ȼn�������\ �f�� ��rҺ:�86�ћ�Q��������U�m��2]+}�.R�f�c��򖌢(���p0��6*�\�B�d�L��N�:.�B�%K��&�K4{ 	�;�#������/B��xXb�a~f��b�upY=)4�2�^ͺ�.t�E=��2��&8�D�8��6 ����6:
T���7sf��TFK��x�:Nޮ�}K���ذ�9�s���*'�J���v	�|�Z�:45�!l:��ndIWC���s']@����O��"K)�;��h���цrȴ�u�v�`eeM�5L#�MNe�SQ��0��ݾ��$es�9��U���FJg#��o_A̝�]�$�]'1��>�o��P�oB>t�1�g	�j�����HW��p-\�LS2N+<��9|W�g7�JF_[W�%�f���G	���-�����EE��1��RسC����|M�6�����.�nRPF≬�v�-W��g%�ns�P�^[jE �|�{Jڀ�[oo���}Ts�p�l��rg�+WV´iGw+U���˴M¶�v9:�3t��l��N=n<+����Q\���,<F��]ˇ���RϚ�
!5�p���|��vN�+7o%�\6(z��R��up�(a%�=χI�wolb�'#B����}=bT�,3*H��	o7K��z�Ar�إδ��o��_q��,�:�Ūa��4!P�������U�8n�w���z&M�+>3�k����[��]F�^wδ��s�oO<����s]4����=O���d������h��b8�ȸ����si&�c���8�2�xC�1#y¦��}�ŨsE������@���3�;6/.��"+	�I���C���Э�hbT���W�լ��ngb-ɾh�)��m��zb��{�-�\g6�b�)�;k^	���.d1�>���վ�t���������o	�7� �;���˝Q���y��@C�3 %4�kƟ2�oe�wj�G2�q�}�N+��g\���>�cV(�q
?gq�����"g��h�A����h=���"�w�wI�w�X�]��Ek:¦4�̩#�����%�}�(p���-V����n���R&*n��2ܗj�c������6Q}��m�K2ﯻ~j�.�Cr�]o8[`uy%�*��|�ُ�A)@��Y��[���K��뢶���Z��۪��R9�ۑj����-����TbC�](����z��Ӈ�%C+{GnT��-���[��&	��F_nkD�Z��]�,^�W�t\�'�O��j�����&�j��'L��B�ӱ �Nh��-X*�ۋd�k���o��W���6T�iQ{��k+,5 ƞ6H�<�,*F�z��n�8��QE�u���%v�աN����:�v�8�".�B۽v��2���YV~v�-��º�.��k�
��ekn�F�:�L##�b�~o�8/~�t4,�X�ƌ���'�@+[4���r�8f!��Yr!w*�U
Z��ګ~|���d`��c1��Ƃ=��j"�NIy��'-�e�|��u�h8\�����2�5G�N�ʁq�9��'�8�7M�˥��[{HK�K0*g��w����M^�;s(�>t��}�ñ��;��{��6��i��C�1��l�pin��IՆ0fÖzf0�y�c8nvj4�*��A� �C�ٔa��t��ٲ�׮� V�U�p5�/���"�/	)�R���[�Q%c<�K��U`Ǩ��W����seE�;Ր��\����My���L��)nvT�}�������)vR-�8�t���i�h8��6aj}m^���4M�gc޾w�vOl�#wّ��^��b�����LΧ������/u�b$8M�8��p�KX(T�6�y��p��ql�M� �gi���ے\|�!">w���yZ��;�`��5Ү� ���t;|S�1e^@���i��JZ�[�Khỹ��X^�\���J�:�V'�v�4R�J����1�&�q��}a�d$:���Y�9�z�u�.K���n��D�K��c���sܸj䐂	h6{/i>�k]3rۭۅ�I%��J7O�S�:jș뉉� �Ł8�f��E����Ov�0�7_c[��R�z�3�=d[������:��8^��J�8f$�lz�歜�AD�k-�'wJ���Ϋ}�+�}z��^���2�6Jx*m� �/��{�����{�n�7:��ļ���Э��8*��=�qY��� ��`���5K�6�)��u���|b-)g��v[�\��&Y|ص���GxS"�j���"X9䏲�c�!�- 	ڳ��]Z�����z����{���ͧ'������E��O(�nݶwM�ַW�q�]i�s`�,.=����b�K�u�y�.!��d�~
�D���� "%��k��XuϺ���3Z�
�!u��Åh���:k�b�u^����fƇ]J$~�{���v�� Z�,i�Tx�#7��&�=Qfn!
��B������X�U�K����}j�Z�F��m�z�$eZ)p�Mn,Mh�ɱ�/h�ŷ'���y�	T̬ ^j㲸bPu�+53v�,�S�$�B�g���}\�M�X!�r�Q*�*�f�s{���`da���{�7�ԥ��Y~�{=���tX�*�7��g�1q����"U�3o�75eU�e�ZT&��d۹([E��N���Z⧞r�X��U~Ӄ�wgX��u���!J��Q^��B��&;Y�s��-�y��%!��;�c��E�eD��ZL��\��p���w���V��^��mm-W|�s�w��\ܫ��Y�s��K�*,�Y�r�om�
�.ד�謞���q��`�zA�}ت�W����e+�f^إv�*����4��ꦭ�Er�K&�D����F���L��)P��<����C����~�ui�+r�Eh�W�`25.�����h��4;7Q�=�9���t)˰T"��X�/{Y��5g|�|�E#��q�Z�6f�P�Ɉ������*�46�6;���Iϰ���x���;"{y^u���#SClN9�����8�k�cm�]�ʙ:.�"��t�-NkU��/vp��3d��V8CP��qc�b�(󧦕����N���D��h�gr޷�;��rbe�K�[pj�{������J�"��l���:��\��		� ��2���2��J�'��5�d��\�P|5��O�^���0��@��ek�1?��)1ۥN�����63��n�!�}�����_�C惱V�R��t�נ2�����[��ED��ޫ��غ���+�>!+��6��	c�kŗV��	nzO/#.�9	�U��zt`L��X�5`OF0;	�(&�b���t�@'з�m�XM'ˮnb��SZ	�'�!6��'>CÌ����x�f���V��菵������]X,�{vR๚)=7��0���c���o���c�v�^��Vư&���M�yL�Q�����,7��W&�w;W!�����a})��!O&wo0!K��Ǉ�NO_h�}���O!���;�gd�5������嚲uV0�*Qm�xD�8S^	pӸ�<A�m�8ݡY�]=5���"��Y�6Q*g$�����S4K��5�ӣSN��oj��7�F��g�Z��� 	�A9�J�d;�%����%༨j�N4��Ler=��j���L��Zz��tO��j��"�o�r�`$��:��zX��q���ZK�z�+�f��Z��A,��[���+-���m�3��k-jp��9�`��]Lh9+
��"�@3i%<�#3���ڈ�p��9����2>�)�qN;6�VM���<.���zj���tE��ܷ���\d���͋��cv�*H����Y��PcTo���	'w�
�
}�v�K�X�"�D�lL���g`�=�sy���y[��2�R�zo7w���L���J7����%���*�-�.]OBɰ=ilٰga���0MY��5��5th��B�d�:m��;� �'(�PRpy;4A=���|v^@���6��+���o,� W�L;o��X g� �!��v�ې]i0���x(�;a���>�,	]Z{C��ozސ����]A)�j�To)̱�1���M�W��C�)N���o	�ڬ���O�4z�F���L\�;Z$5s�8:s�h*����us�k/�I�
F`�c&��3Ndo�&����
��G��wm K���wK�}��d�S3qg@o��v�u����;tb�Pj��l<�.�r��
�\�q|񨣛g�ڏm�)p���Ӣ�p�Ӈ;�m�0�έ��sӅ1
�N�,����݃��)���?�<=��z�����@�\�lQ��.�w>�`ftE4�hq��BW��c��|�d?(G�vqAb�ܵ��A�C�v+��k�M�|�gB{ �W=��R"Ρ�����vR�&I�yٍ�`�ղ��\��ޜ8m"�1��%�t�޸m+�����+Lց�pN�����j�U�=1夜�ZR�=�<��SIcO},5s*慗xz�w�R�+�_A�y0S���j�]�K���%M����A�%�%2��+:J;+��ZfԶ�B��/����,�|�{F�޾ӥ:bK8RB��K'$:�o�,/F�j�Λ)>B��Z�1q3BS�d}<f�B�Ôiu�a"�
�]�--��R�n��Sz{k�PRZ��.0�'rx�:f�U�}�Sݰ�z�L��rM 
�
)�q\�{Ub��{{i��'��ւշ��6f�r��5'�B8s�$�uv#��έ��o���X��m�1d��YFE��ٗA�̸WAR���%�3Ny�r�x��7ɞ���]w}��m5|�hz3�O��@�p��Բ��ď����W���=w�b�f����̧X�[̩+gkh���������G=7vgzKyVs�Ѿ��.�w�P��gr\�;eMa��R\�*�%�1܀ⲭ�ƓA����o3f��Y�n6�ꬮ�Y=hyi�Yti�ۊ��f�S2���?X[@���FբJ�hV��#`��
(DZ�kb���F+B��m��	R�
�*�(***6�Db**,Yl��)h��V��Ъ��-���e�+-�b1cF�E�*�*�сX"�+��"Ŋ��km�*�������R��VDKaQ���E�h��R�*��-�Ԩň�(�1aXV
�b��ŋR�UTEYUcm��V[A0J�UkE�����Z"*��DTV+AB�ب��"EQQX�D`��X�b" ���5��A`�A-*�AUUXVE���*R#Z�"��QE���Ԣ*1ej"�(�[
[DcȌcPX�"J��TPEJ�"�UUUKKZ�*R(�����V*��EPP�F
�b�EV�TDU`�DPkZ�E���a`��R.�1��s�J�iTݹ��B���y��)��TS��&M��/�ʻ��_#[�t|/;-n��gV&� �I�{�ٛ�-�˱�q���~�@O$G�ګ.�H��F��#\։�rp��5T4Te�`���bo��4�Um	h��娵������f�S�Zˆ��{�>W�m�5��F��{zF�E�q#_+����)�KΝo.��|6ZY'�w?���	6�
A���b�#qHu�M���y�3N:��!�K���y5]-w��W*��}����Q�����[�b��Ցli��G�~�V�s�z���41؇W'��k��|݇���s#;��rrJxdH��s�ճ{žx�j[�NJ���6����k�/����b��N���k��ݤ����Hnp^o��}�	Z)VM6c���	�*�X������:�1���W�:�]}9�����q[�]��5��WK��u�J���F)������3`���]�c�^W]<u�z%^]�?����c�Rv�����s��2҂Y�ե�u����ICX�Hc͢3�{�c��w�)Mr�\'G�M��-�&�����G�� �]#��Z,{y�9y��P�M��rE;�H�=kr�iP�����a�.�+HoV�㳽�A�	Q���e��'����]��R���9Sw҃w�MXM۷��U;�❌��P�kw[�:H[�j�r�{��^1=X��@��$b-�馵�\�jǥ�v����H�&_sś�:��ꑁ����(jM�^��}�ՒR������s��b,|�˒��\9�mت�N��t_fz�����o�	a�|"A�ï�r2�t'�tCl���zXH���h���D�*�cA���ian�GT�Z�Y}���+�rJ�hS��U!�3�#��1P�c���3�Ш�~����X�Ղ��:��l蕎F��-���[���vЙ���滟B+�i���F�x�k�g�4L�a�"y���Vpwg`��^=�0N��_�R�	yVT��l�V7��z�Zp��뷑%�mVqiF�S;4��N�Խ�\�����=j���N#�k�E��c3Mf����%�N� ƠՕ�h�+�t�C���I�����6��M�V���Z�Ԇl�g<�fI�N˩M8�&�N"SFh��i��:7��Ŭo(�����]ָ�W�E����1צ�+��np��;��☺�;aKh�ak��+�_�X�#���3�pœ�ܜ�v��v0�vPЇ�V��
����?7���xw�vk�,`Ua���b��Ʉv^�{�h�Y�!Q%�/�`�A��*�\}���of��+�)']hT��UmtuVm��ʣIvBxja�<eߙ�}��*�,f�U��ƶy؛Xf�	˲7�sE]	�}9(Խ�C�l�W��n���;5M�X:����z1,F��6��
T')/�ԕ��m��5z�Bؤ��	�u�����(л�KX�=�ˣ}Cr�68���WE�I�)��0ﰬ�%欉Z���c��Y�8�ջ�d����R��b�)lъ��`J$m�;�cN�*�ʭ��n�ȱ��+�T�{=ζ�Ա�^��}T�|�ӕzDL���6�k���ї	Uq�q	r��;T[�Vm�j	��*�B�V��'�f�}v��٢��AVq%@W���U-��u��F6�d�L��YV��jyv�Gf;���ء��
�s��
�&�v��e��iX�������`b �y��ɞ;E�79眭�5����&]q&��R0lە�]wJ%�М��C��M��b�R���I��Q��jׯ#6�l�:p^t'�A F��Q��+jw�!)��C�ߩ���	��Ȇ�E��n��ծ�R�!���+� f�c@Q�k��g�xg����P��܅98*��uoIx�qa\�c:�n{IL$TP��	�+`DN�,$C�*&(�܅E:�������8����5]Sg�	�2�z!�
�ɢ궏�)g�/�De��*A������g��Zd���]�E����Nz
�F�9�ߢEE�:��^�N	+!A���t,�:��g*;O��Ծ���c�ݻnc>��8p5�7��Ԡ�b���r�m�uz�wq�����v��!�X�%Ɲ�Ϗ�UI�C�v��-��E�4�lj�h̕�i�++��G)�=.��g޵yJ��jFAV9��q�c:з	*���ܯ��#�{�3k�χC}�r��YA�5d���V><eR��=t��s��x�^U ����p����43l`�k��,["�����|95R�x��	Qn�j -7��T���b��G�%pnϦu�/��N�6�Ї������l�![�I�,�=	��Ɨ��3�1/��r���̮��l��� �p!�C�����Z���gr��;�pU�x�aY֕]�^,qv�����g�;3�O��PQP2���k�W��*
,SO��̤������AN��9�(�>�U�xq�h��r�Wε�?�?k���3����8�^���o<�@h^�����V�����z��y��	�(�.d\	�x�d�v�#���t5�9X�S�z;)X�F:�]8�'T��"����X��TE���׬�Sb[9�3�W�ӗ©n�ԣ��=u@�PEN*��L���n3�[�~��e����*A�Q�٩;�ٝ<z]�����(_��B2+�r��_�a�W�A�t��	��Q~�A��p�1&���B�=խ������3��Y�HY.(B���'�1��`[�]�O��������n�M�y�"Z�wX��tw�\��pg��s(�>��U�<�V8��8�#��+�k �-w}�)��Q^�7�ڜ�*�f�E8��'~&\!r�ؙ�9Q�>�(�\c��#*��#����9�;���ٴ�Vz�^G��!��L��ݚ�����P��y�K}�o��f*�A32��l!��@�;Zα�/���d��[۟{%�y��u-�d���:��>b��\���Ha��n�~�h�&���>��z1��ްv٥aa=kw�|��z����R��l��C�6�p�:\�����[���V�p#�ϸ����v���zڂ��������E�C�l1~l��/x2�T�������(�ޚ~��xHq���ݓ슻G"���M�/g�9�����7IJz��Z��w�y���h�"�hh�f	npT��d8%׎� �yh��s���u����6[xn;#��A?MLe�X@��MS�۫��]k�a��q�[�ET�Ź#�����aU15P.^:pe^F��ltc�3�2�&��GTC�B�n����������v�҅CR���X������:����[^�������Ww��͂�V�:Z���˅:��D��ۇ�1NU�Z����-N9�˘�Pm�LB��K	ץD���%�=R*�&�ds�z�9X%�A���׭����O�fo/v{�>�/x$� ($>�3^�3B����t\���/�օ��n�*�+��d�kIW�z|�i��C�/fc���jۧR,@q!zv8��!*�]9N�q�͸V���̏���Sf��)�+�=�Rںm�Z���`���3�u&tT�u��U .�µ��b+�rY��o�Υ`�k۩g�;W�r ͞�����<�tcT*�S�Vp{Q��ʭ��tuel`^� eiJ��l�^��r�)��.�쾮�e=7�q�b�����)��Y.MA�%Q��6z����;o��+24a��$G�͢j�j��g��란j��O̝�����Sj\Q�Ը�����=۞�7�Q�98A�Sy*D�7"�G��e���d+�����:�N㨜]ӊ;��<�U/]*��,h��jFB�ώ��ۖ�LC.�]L6�	���;'4���>�Z�`�
lD��5(G��V)"��
RPXu�����s��O���ﰅ�m����t��s����X��G9��`�eL^��M�,���>�lR���=*3�Q����-�7* �W�~;�Ns��N&)址l4}�4GU�װJ�F
nf7d�ni�����y�*_t��K�p0��S#��{u��l�C���[�"b�^�8�"���Q%�+9��N���0yE���8�g�,�P���bZ�I��ޫޝr/dQ٫n�qy����=�h}��g�C8y�;�?eոQ�>P��+.-�)к##]�x��RR�nP�w0&6����у�(O[K���m���~���e[�� 띆��v�0Kp�=��S���l�{�o-���E\{j���	(>sU.ƚ�j�ܨz����')ܻ�F�+ttǨ�
���ce�rue8�pڌ=��6�!h���U>���}A�A�%���B]t�ԭFu�<��y�p�L�;qo>Pw�=�JN@F}Y��@oU�Kt�\4���*^����/� �R//��d�Xi���hhWX��EA^�?v߶��}g�H�k�'[K8����L<��|�z�:�W	}Y���<g=j�Ȱ�R�zʙ��Df{�qP�r�壚8퐶�yN�K�Sy�N c I�N�I�W�F�r�"�Q�n�AN�eF>��ඁ��0�_:���w��ӚC06\Bv>��ԸpO�x�(�h���L2�r��W����$��aet�`K�1���Fa��Ă�#� !X����J�D	9J<@�j��l;��zrk�O�}����C���ӭ\!Q�W+�ߔՈ�9 ���X)Q+��t<`�D{��<�/]�����pY���s.���P��sO'N
�RpÐ"0s�R}�TM{Ej��ú5����#��9������ys*�P=%�*1�p*m��Kq"��k�N���������A}R���=f��X�r�%\�&wv&�ѯj+�6#zu�q;L���'p����'����^?o�H�ev�'��o�ȴ�4��b�(f�Zyt�=]�T���/����Vh�#�;9uu�Tյj6"ݔw�Xި�/�ź���04`�͜����Xp�ݷ1�Haz\8����jPx1N�p���vH{�x���u={���W7�KƝ��>?I3�����Q���Q���92�ոʸ�\���Z�ϧiO2~���H����.6/:зBD�N���譌MbI�u?>��_����\��^�H	\j�ǎR��=m��:�x薗Wٳ{���5�s_4�-7t�
7
M7H���r5&qIS�l���T�nl��58�8%��U۽�C���0
E9�$�9��-�\9��*8*׈���U:�X�?nU� �+����+yYD12�z���Z�H.U��j�XP�S*5�:��*�&ă����o`�!C���A�q1�TTm���<�ܶ��}j�u�dZ����!�+Jq������<'��@�Q0�0�PQ���v�=�������YO�����fː�=ϯ7��в=_r�Z��i`��"����r�P��%�J:�p����tQ���՞�6��լ��2��2��5iI�	)�݈�-��xpQ�)��;<
��O��Y��E��q��z�݀�d�
���i-ie_��L'6�g)�ˮ�ӂ '@��m���է���q����s˳�������%����t���^��Ll]Z�1�WV�w�o�>�~?w�T�u�K��!*)zuL�t�ʑ5�qz�ѻ��㫫�y�ۈ1[$t?j�p�sÝ��}y�Q�%�_�u|���a��uގn&�?]OTT��^���S �߆��ɟWz\uC�<e�PZ~�W++�yk<mG���vރ=Qӱ�j6h_2*���Ë�Re�f�S�# ?C���{���V˭���Y�[:Q�T���"GET������TTx�`��#nE��l1m�c�D�����*1BZ�U��9�l�W/��8ҕ���,{�}a�Pe~�v�������;��s�E+���x%nM�'jxS�u	�\�^�hا�2o���q�p�E�֪�A{P����^A��ny2:}Ad�꼚�r�ݯ*ǔ��M��
7K0CQ��j�D�|`�s9�,E[�Sc*���T����;Y�m��l���ؚS��HO��{�ZH�fО���;�_QP��0�766��Y�ϭ�!9γ�lrU��UU��5�,EOq<DF���Z��=�$��tY�~:pXM��}�JK{��x�FM9�8�&��QN�԰��L���u.�R�`K�q��}��%����t+�e���j��3ۏwoc�9��)���r���y�\'��ڮpZ2yhLuR>_4�*{�:���Ҿ{�`ֺؗ6�����Nh�x�$�b���tJ:; �H.2�6���g�����/b�y%����Z�pM��[������p+�a����V^.�57��*P�����q[���>y��\���E�PQ9V��"ࡉ�k+vS���t��8�Q�yy�0	!ݐ���#�[�yx���Q<������(�Sυ��ԣO�;Q>K�f���B�H����yGw��IV�P�I��>�����ಱq��p45�J�6�|�6�X�y��Um,���`��+�mK�Bl�F��D�v⫳+Yz���	�q=����s�v-K=�m����R�x-A�Ջ�P ��gxun�U������Q�Iu��<�m�9.�U;F��:8���Zj��u1��h��xo��t Hf��2�|7V{���&*�ruc�ٛK�d��g�(E\�;�Mf���仭b9�Q\�����:m��6V�ʑ�sj=�J�\v��yK���6((����WJ�[ aG����^��M���ΤAի�����U
i�M��~�~�nR�ssy��=�B�v��\:gN9�о�%�c{Q�ۅ�i�$}7ܝے`�K$��r���}�҄ܞ�$���ŦﶝΛ�A�t���'8}������j��<��t��܌Q����m*+4�\m!9����{�h�8��Dv�7��	V����'&N�]���HK�
zӫ'�z�)O�j�q�A�O�+�.O�&!�zn��m�y�~�c����g|�cAX1�)y-��Nb�qx�nn�
N�4	����^O�Y)e����F]�n�M�Bq�veB��,j`6ӛ�����a�X;N�͂�IWR�am�}�˨��N�.�;'w�3I�]A��׊���b�y]��x�o��]N:#ˑ︯-�QT�U���������Ͱ���7+^G��ż՚�p'�������2��g[�/�L���:�{.�`����Yj���2�8̂���T$ Vef�Ƕ�Qyw�6N]E}��ʽEp�u�X��඗�d�<�h`���p���1s�B�+H�L�$mֆy�� �Gu�.-�6�YY��]�o,�j��C��C��,[�T��:۷u��		��qNw��� �����f���9i���E�d��_j،��d�9����u����	��ݸ��Qd�;/$����wYá�$.l�>��٧�낊���ּ,�g��E*�(ȣ��뗗�sY)�f�N��h�$3����fθN�|uU�q.5ō�}���AX�,E6ʂ�DTb�"Eb¥��T���*(�H�A���E"�$b��X��Q���dQP`���"E�����X���"���#`(�B����PDQcj1�*�`�XQD�(�Ŋ)ej�UADV#�1EUYX�k"�QY������"�b��12""��[IAX*�����(�A**��0b")Z�őTb�����DATdQ�,m��"�+b��������$UQ��Qa[b�DQQ���b�(���K"�*"��� ����DV*�
�+��Z؋X"`�Ь�"��(�b*��VȈ�1b�DUF �X#cV"�UcAQ���*�Eb
�X"���dE`���k`�aP����R�DF(���jQG0�� f�����e�_Nll՝��~Ԧ����W�9a�gU��+;s�в*�>��J�ޙ8}��}� ]\Qa-zQ��2�9����Uv^�{����P��@7�Lb,�jf)��(�	ۏ*S��������*���˞2��(�z_S�_*4z�v5]J�=?������3��x��1��n��OF:*"KT��yÐ�C6g6�-���4�_˹љ�����gh��fn˼쎦4q����>Nj��P�^����շN.�\����S��A�{QtstHy�9ŵ���u�Rƺ�"���Ўw�>L�J�sQ�X��6<����XC�f+2ɼ��.�����M�w��T����Ӟ�J�3��V\�y�tT�p$:�=%d�j;�v�s�m�G��~�� c�S&�A�"v��:��R�rt��\9�3w|��&�A0ۭ����̈Og�q�J#!X����A�r�gLC.�k����v��5b��!j�R��-g0r;<!V�9jO���f)�X*�2���izxY3����~>�`x��p��B"��F��^Ȣ7�W��Ԟ�!
����\ 2�0^b]Q=�u�-%�̭Ann1��C�chAVw�A�
�y���g�Y�U��`��i�*�L-VS��7��᱖�u��!��ȃڬ�狶��گ��%��<�������'1S��4�ܺq���A��E/f
��h�)�yY#�d�ue�u���L.�T�����(��9�s������[ �G�3G��k(�o��U^�P�W1�;�n�չӐ�wd��e�*27Ѱ�#�|y"�tR�T�:!?��v;z7O��*�=��=:�mb���t�d�l�qy��!ơ����['���{�6ToM=�6�8��YE���/ʡϨdӒ+(�y�[X%ʯ([N_&\[(ݹeA�		}+�����1�U׽�]%O���$�5"��g�,�EB����`�Q/v�v�:���w8��s��ޫ�r[�
��IUB�U����Y!�j�b�1��,���|�+&ʭ�j$�Q�O��\�X����#E�R��V��Wƺ������nL�{FՖ�v�Ї�D��
��<g���"��R�zʙ�R|�7R�%��V�+��╻[���EſU���▮�ټj���Q�n�wSҴs��Q���v��`"Nv�j�0S5aW����V�
�I}��x:�Zj�/��\���ˡ�\ª��̷���5y��o(*l���s���U�#���׵oo�pU����)�[�D��k)�Ҟ���Mu��S�DD�7��\�!�vVg-�����^���r�C��֨�����6R�l�(�w�9���x��h ��U�۰1H�=u5�^�u:�W�~;d�D���u����|H��MD�(���ōQ]s�#[5�a��x�-�����IS#��R��9�Ds.(�W������[t<`�B9Kn��𽕗̹Y҄��ܰ!@p]빂�����.���|R2�����qh�; �BQ�X�AU`���{;\��Y��"��[��J-ʇ��WPS��<���n��>��.��k1zG�����Z�#���;���l���^+�۶�9�)p�PyGg.q���ځ}�[%��kO�tr��#6�ץ]+�$M͙zk!��cb�m߻qBmd!���CQ�����TV1���u�YJ�u{4m�s@W�dP�-�# ��9�e۲��>�}�U�<�%z��X�hŎm���z��l�]���ur�{��ϥyU��ˊ�k�z���C�K�AѤ̉£1gv�4¶�Ч�Áa�>n�q�^��v��)*p��"=�8PQ�ns:_&�J`�u�Uսm��J�c���X���� �X9��-�\XuC�z�dׂ*��cje?i>��'85�#ym�d��q"�;��'Vb(����7h1h��v��z��Kυ�Obd�H�C<s��}�T�)���9�$ۓE�^�[�|[2�ή�L<%M�}���R<2��-��{]�Pu�c��w50&MW˩u��^�������}1��<���J�� j�U����������ʱ�j��.�[���{�"�ٚG�58�9�
�葢\-���D�:�EA�|g9V9j@I>�B�&�d�~��O���7��K�D=C��=�^�ꁳ�@�AOT�9����ÿ����,�Jf�j.�}���g3+�i��������u���C�.��H��K*.,OWB�.�����K��K#G�T(�FK�v�ہ�P9 �e8�
��}��]��U���IOs�<��b'�s*s;�AdTR��/��O9
*p��O�#���z&��K�(!.'+��,��<�_��w�V7��({f2mϦ��9ʦٿj�q}�;�2��%�	�9Q�c-�8��1��қ1������4p�<55mD]y7��a��s�2�<ݚ��1*��	k��ΖQV�zi�D>@�>2L��W@�**�ł�F܋�[up�\�'?	���6��A�R�}��6�f��A<((�FFCvO�(]��~�-x7xx��E�d�W�Ф�n�@UM{�*�JG��u�{�����gm�3l�몍���͒��7#ń��t`J��Q�lC{���T�o��}���o�ay�Z���r�67n����4J6z�������
ڻ�ԞG�������C{FJ����UQO׍�&��uZ��= �ط�ױx�Ns�J������,R�UcÏ�WG�ڧ}�����*$��D������va�X�������A��������`_{�7�ƣ|���] é�'�MTt�U!
5H�-yӀ]��͋�|F�F}� ��c���Q:B®��B��輆m3؃�Mb~4F�ɩ�u�#�=�6��X>�l��Y�6;&k`�\�J�W��2�}9q�z��
C��˃�b|&�Ҁo�(�8�ۇ�1NU�`�S���'i~�;9'�~�u�_��WfK����α|����WR�s�C��D32��Ά�L2ϰ�����8/]�rCޒ:�n��92f�eF��Op}RW�DLLm���m'Ml��d��WCb�,���t�X��c���׼|5������}p���{���/�P˙3�q��TۑQOkc����w��J��^��;@��K*�v��S�������&U`�Ą`�_4�Z�u.9ƪ�}9Δ�.��N���d�8�߲Oh�!��dC~+�v�L�1��6@�0S�����{���TX�6�D#*��f,b��f��w�����T�n13�v�[�nڨ�_��kmSp����>��b��@��|ޒ�872�����C���-t_-u�Q����>�x/�٥"0�qh�����p,j��2�UM]k��JKUc:�n�~uX"��>�UD�*�(�x�tBy~�/H~M�,f�!�ֵ��o�-�],��9 nu�$� Ԑ��tN)"��
�2����6��{�5l>���K�0���o�<�E1%�j�\`n��^ӃS�Ȥ' i0{�s�y'{�����hg=��+�-�\c��7h�s��ŇN&)址m��=&g(������ϱ�����B#�Fa��#����=�4֎��}���yu�q1+�n�Fp�{��Vbo^�o�����{iTQ8������F��_R�ڋ�N9ۻ��%	���,n���J5C|v�P��8�cˇ���A|b�[X[/Æ�_p�+ǥ37�C�휳�^'���t+� �@�Vu�	��uײ�u�|4IREH�dS=^u+P�Xj���'gOD4�]hv�
V��:k�޻��E��':�N*�騩�B�TJ��FJn����~� 7=	�D�BX��VZ"�M�]�x�g�n���p�5���9kk
]SP�MY��l�[�)�xnxJ�uo]=[m��:��^
/�mu��oI5�*44�tF�eź�k�x�t��̼�[bH��}�]d�����ν]ȝf棽�X]M�ui�Ц����^X�����x&c�)U����p��u��Ƅ�U)����i+ �?��l�"�C�}*:��V9qJ�eL���.u�,A1��kom�sq�{�հ���z��OD��mH�6mʁ~.�XN�Bs�*gOj�y<�\��ՏQ�4����U�V�G¹��/��%����qx��"�����zAdl����FW���ZWxf/� �Q���yr R�����j�k��8=93E�R�'�syf�tW)�Ȩx�nB�@����Ds.(A:A
�3����D9M�bf�����C~
m���~qo�!
�@�f��ˋ�T�\;�@DWML��=X)�ӌ����|y�j�GQ����O�@�E�-ɱ�~�s�����>����i)��_kM��:�{�j�n�Dw�V��t�8g6Nex۠�λnc>�ŉp�<��3r	��n�V޾Ì�r�9�NB�}1�"�ԭ5���V6,fۿ^�!Ƴ��GB���=�(�j�=xm���60��D�7��l֥���5���!V6:���7�A߳�d�cy(ٳiۘ<[��c�~�����\+�:M�}dd"��؜>�6�՞t��=x$i7+�oe�|J޷����Î�����4���N~�����u�R֩��G[��ؕ����C�$T
�J9��}{:��'(t,���D��s��@kl���k��?;ãD�����*�ˉ���}��X�х�m�Y����hT��2zULt�F������eX)�^�j��7���V��J�!ã�B���Q���� +�2��!X΢�X��6H-V&�@�Qp�G\���j{�����76�owd�S�MVy!ȟP_4���ޫr�g�C��P+|��
��dJ��ޘä������U�`m8�'cbC� h	P��=���fyM�mP��m<kcj�޹���u4�8+F�j���{������t4z��5 �
=@�;�eA�_Y���}���}�n�O])������S����4�EB�K��(L�J�a҃��j�����\�=���&:u�8��%[;
����u��P�8OE{�9�jaˌ��9�0���7h�e�~�D(�Q]�=΂��.:�ב���蚋�K���Q��YO��m�*S��E�I���ʅ3��aۈL��=Ш/�o� 5�e	����:_iWh����{�k*YK��f��Q��)�)yLV��B�Gd�⛐����p�ެ;ud �Q,�`���)+8�POj1�GzcyDҪB�G�  �e�o��'y�2�L�ϳ[�x*��.���)��g��\+�%�	�U�Aț�gr�]��h��)�>�Ll���q�B�n�e���_��5�ԬL�N�;�bЊa�]�G(z�U���A�a"��#�-����>:���{�x�7
y�L�Έ窥!��.*�>L�n�
���Cƛ�iW�cޟSXR(2�kDD3�Wj;��YM\p��P_��B^y3�n��;y��h���h�M�nMM�+��s���K֛itT�ɑ�1�W��<����9�0�2:�&��,���n���1����*N�xt����^'ph�XY�a���xO��xzW��.��lXO�����:f6�j�r�� �qQ���a�X�WV;l^{(1�*`��ݢ�f�����X��!�NB��-��)�rL�N}w�cݾzb�e$
����.T���Eۇ�1NT�T�G4��ƶ]]�ci���mM��sV�1�/�x�5Օ9�!�M�.���b��^su���ƪ��HU�/��y�q/j|��;�}����XB}ܳY�n�w�@����W��%������r������w��v-�q u���t���',ܭ��G_Ō�@`ˉ��y���o�wn�rkp���]�#�]�ܢjp�S����9���w���b����/��*H{�G&���9,��hah��xo�+��޾X_S�c�^T^,#��|�[�	KS1��Xi�pjG�{�9/qVt�ռ��+�����s*|Σ�uM��=�}ܙ�P�j�$M�B�ؼ5�K�]���݉�U��P !��Ӳ{�;�̨��NΔ��B�2w$�c2���n�9�ٽR�T	��T�#��cf��軉p܍Q�`p�N4F;z���p떪���W	�<���uX"�L�iT9C��hd+�"`�2���5|��N5y�(�1Kit�WK	ר&��y�u�'�
��'�4N)"��
d�B{�{Uvȭe�v��8�QP�ڮ�q�/�b[UP��ᩣ4�����r)	�`�싾z4��c:�`��7�� ��"��ny�t�^W��u��ݿ0%��wn6ҝ}��<Fma�K<]#�`��:>�=�:#�dv"+f�8=�` u�	�<���v�#��w���N�e0�˅�f[�9yG�F�\�l!���m8/��l쥗������Jb��p�9B���Y������QJ1�|��\����Vzd8<W�.[�g�����y.V܃[V�����1�(��L�5��:��Rx﬘;�B���2Q����d��9b�V!e�`C�T�H����Y��c�3��{w9��ku�`�
�b%���^�hzkC�-��z�Չw�F�7����wXU�"�gg!t�1'Z�Ш��r��:���5�E��uF�s��9��J㑆��wd��!K(��VK;k��j���������r77�ń�U�C��q��vf�:3�dh�����GWZ�+�9m]>�,�z�򕶔A�C�zkM)5�w���]ʻk�="�鄍Xa[�eL�q���J �܎��ܰ4	���r�����T����cG��Xįor�г�s�=���'
}����:)�Whn�ɬ�R����HB�C5�t9�ul�E�W*���!ql��m:}�⇫�Uj�[�����:�N�v�j,q��-gX�KAY�7Ϻ�'ͺݛ/�P´pk��a�h_Jxtƚ����J.WO�o�_#Pɸw)f��^�of�0D!%z��S����\���)�O�"{�k�Ύ�*�y�,�=ח}�c@��Q�H�r�v�9�r��wA/ݧ��\�TV��ѕٱ�������e���j�jڑ��J�^����\��r��L�e�����#}<2{A4�2���Xv�4����)}�7���Qu4y9HY �!TK]z!�zeXO=U�����9���v��`K�r�+{���8v��J��A{�1�L�٨�hѼ�Q:�V:J+��{]�{�ÞҺ�=��cs�I漩�y���vE��+xF��{8�pKC�A��Uⲥ�j���3����ܸ�������ݨ\���^���B� <�Uۖ�u%��߹����*�܃��R���&B&��WZ���ˣ��(\�`���Zv=S\��F����T`ܘ���56��7YA�/ǳc�]�)�z���cİ�Z1��x�"��lc���Jk��9n �G�n�/����G�o�ӷk��g�L�QÀ%�=�4�7��wc,�K|��w�F�׃�<�zt���S��b��Γ���F����:>�����ᨧ�n���S��x#Ժ;jFgEj��x�]��nn����s*�)�37�1i���dpf�-w���y joa��ٵĜt6)',��Mw��p,u,�#��;��S�e���1{��Nɧqmb;���j��z���ڎ�Ə9坷��W���k_V����
�Ԗ�.�W��Վ!�t�i�l�H�7)U�{G���VT��l���8�</ �h��A��˥g�.���Ɲ�w�����k��VE�#TD������""(?�EV"�(�AV*�**���T��
��Y-��",X6�UPF�TX�*��U��Eb�
�QX�V(�m(���V�QEEU�b�Fڊ
����X�b��""�+TZ�b�"�b �hU*���F"�QEbQ������TEAH�5���Q-�E�ڊ��(�0�QDb�X�U�
V�dcZ�1U��+1X6��A��iUl`Ŋ�F1ZʩR�c-(�h�m`��Ub2�*"(� ��*((�6����mTRZUQPF+-*#PV�X�,Eb4h���TTQ��V**�"6آ ����#[�m��V,E��"*}e�H�J(ʔX����"�V(����EPTqF�Y# ����Ab�"�TQPF�ln�ᢰX�(���Dm*$QU0؆)QUEX�375�cV�V�J}�6o�u���;)�_"6��ҴrtGn3��q���lhp����.tbw��y��x�Y`7K]_�=� ڻes4�)t�d�?p�t.��A��j�6+}e߯�q��E�q�E8�	R��9�����[��1q͜
E���q�n�x���\SÅ�_p�-8MU��t�u�5��
V��WAR���:�s�[½�(9ȱ�J�R*��?U��&�9����3��7���t3��N�q�C�����J�8��f^�q<}�䂓hw��bf�HV.?f�'��a��ğ8I����a�Z�B�!R�0�Tx}��T	��U��뾸[���D�v�U}����$iRWz�a�����&�0�d��bgvu�ٰ�w�Ҥ;i����(
)�h?{�i'��&���8�!�q0��L��f�d�>d�{�8��]�׿~޷���ٻ磺)֊L�*Iyr��*��é���3�y�B��*,��XT�C���a�E=�Xa�P�:}�M=L2au=�2�Wl`L�L���~�}�O� 8�G�k��°�
�!�G4�B�̚3� �����E&�2�!�R����&�y�L$��0m��u
�6kؓ,�2�����!���%M��~��y��{���̥z�=�*<* J���8���6L!��`2�0���):�`d�Ţ��aS	��*,�~͆P_�3�`�&P�_�kR|��B���0~a��y:�G�Q1��y��U^�|G��Tt	�d�A`y���]�R({�4�a��a*��ɴ��+�k%E �;E&�:��f�ϙ=���fP*T�5�9�d�
)��y�_t��g+**{�xgc����#�����e<���s�����7�g�wu��LzÚ��R~��)6��ez��!XeP�ݢ�ɔ��9;E���
��?!�S|�]���Ɣ�#�wZ]Ȁ�`ySa\��ux���rsFpaΨ�m�_89ܼp�fq~�3���������)tx6��b@�βr��o|pJ�6�-{���'�HN���y��]��ɷJ፺o��3�v���q��j�k�����o,Vm�~��l0�	���	P�M~�I���L2~/qQC�+��wY&��'q��,<³I�9��6�hVy����*�*��I�a�>E��<&<*1�����Tn�o�Wvk#��q0�����|�E�l2~eC:���A͓F��śN�����i'����&��	Qa�<����e
ɩ�bg�Y>p��P0�.=�뵽]����d���l�G�x�(�C�,S)&S;��&�yHWS44�ڤ�y0�Ƭ�g�8I���E �2߳��*A�����i�����{��Ag���W̕"<�*�~�7���p����2�:<-'�����&s`� e+'�m�d�
p�0VO�31f��m��;a�ՆX~a_2h���6�Y�%}�I�QH,��bL�겡�����������ǷWݓ��2� �	���b�Q���A}/�4�!�~aQCg~�2��0�]r�$�a��,�
��*g��|�d�LلP���I��2�hVy�~ϲB��³�9�g����5���?��>>���������{�U'������,�����!P߽��ɶ3���(Vi���B���H,��1�)�2�wB�b�'Xa���O!Y��>����{����w�{.y�[��(��
�]bN�I�+��g�Y:���(J����}��M (�M��!��AI�}�欟�~�rw�4��b�I������8��)QH)1���>���?c�{�u��ע��B�<Z��ް�oY�>M$u����z�Qd���P�J������H:�̝�?�'�i�V����2Tc�&�$�w#� ��S�9���Z~��z�u�ݓ�:¸a�Q�4�Y�L5��QH.�`a'U��`��B�멿���8�)�Ϲ��l�g�TS����
�g~�4�wa��}��Y��` �<9���&�v}=�}�mb��+��&�Xa?$���R|�fg�s�V0��E�Q�'�����2���ƻ��AIY�~�pÌ.i
�`6�&�y�L!��pL��"����{�Q�"%f"������c��~�۸�lg#0J�TFL��t�GXc�o*��Zr�EvnJX�^�^#�Zg����ۺ����K���Ar�3�.���#ݘ���=�}¯H^2��m���-
>���:�V��}�(��,���gU�T#�%�ov����< ��U�S텎J����l�j�P�A�6s؆��i�a���i'�+5���)�a�R�|�'��͓���9�X�P4��&1E�d�ٯ��<�H,��M������s�g��^�Z���{/�4���:˪OM���w�M?����<�����T��w�C�LVMOw=�m0�=���)Ru0�S=����a�C�+�vj�$Y�&$�_��?~�wX�c������C,&�t�ĝgP���:��CGh$���]�	?$�9�n�:�Xe�l�y�@*����#ޡ��dxtxIG�r�sO磜�n��c�c�l��f�=����l*k�<�R�?��E�aP6}�P�J�8ɏӞ��ԕ�_Y*N!Y�c�>��B����2�0��)2�wi�J�U���_w�����u���^���6�R_�\������f�g��3Ʉ٪Xu0�f��2�Y2k�4���a!������f��M�w���B�|����Aa�j�
�g�*��%6�k���|/��'P����������P4��b�,���|���L$F,2�ڲm��?j�,+b�~��)�I�o���~B���Ğt�|�C{�(L0���{w�����z<���@��o<�+��r�T6��C'רi �̰��:��
����`~�u��36L'�?8I��I�*m�~��!1�c�c�o���#`xD{#���^��s���k�7���?x�;d�a���&R
N�w�(u%�!S������&{�f��3(}9fR
�gC�a ��"���+���P���O>r.�@�`��q���A��y���>��M�Y�c�d�9�����L���O3�}�3�����Xy�>��g��~awd�=�M0�8�a�i�ۤ�Ͱ�a2}E&M�e@@� ������9����hm�^[���������JśN0�J�R|�f��I����k0�u��q>9�
A�O8u���4���S�{؆�g*M{��d�0���	4��d�.��( ǆG�T��q��D]<y�z��w�%`i�}]b����=�)�4����[�V��
������kOq�{'yQ0^��e��M���G���_�Џ���}�.۱�*Ƥ=�{Ve��J=���N��.7���c^N����Rzd�U�Xh-��9�V2`D�+�UU$���w��K�����C��.Ri*)l�`�!Sfh�I�;��)R|�@�~�����d�����P�J�=�<�H9�����9���}�2i!������g�?<�<�f��o���׳�s�q�&!�0��T���s�B�����-dש������.�=�(a%H):�5�s4��^R�a�:�Vu�S	����L�gS��bi������}�k>�?w�s���$NgڇXm|³��bM!ĕ�u����*3L��Rm
�}E���T5���L:�)6g����to�ʓ�T��?w�y�0��������6�޿u���_a�Ĭ2Φ~O}�)��Ͱ�nw��y
�AG�f�u0�,1��X�	��SHJ�WH�d��7�,0�d��$��h�W
<& cH���n�tKW��\���W��H���C�d�0����2�h{N��Ŵ�a��5=����Aga�`<�'䨲o��X��z�i�	�l�Q�a��>L0�l0�*J����V��k|��{�O���n�àxDp=1���$Y���=���8~�ɤ�-�I�w@QO2qÿ{2��T�_Xu�)
É��e�&�L�;�c,�%v�jD@� D���K�O�v��8巫�j���g�?$���fiP��É�Z��g��5��E ��5�3'�@��pg���ae�v�$�i$�S_��2mE&�}�����`��c�=�C�c�>屹Mg������<�C2��4�(z���Jəj���*C�	Y�8��5@�3�a���N��6�ay�C�TRw���y>C�=�3�%bͦ\���8�'S������o�}�=�~�y�g��L (��w�O�2���P�P�l\��
��'nZ�QgY*f�(�2y0�sI���dη��R��l��y<�H)�Φ�\d	��|�
���߹��~Fq����`�O}�I��6g��?Xm*O&��ęg�I\��}�H�0�C��Xy$\ÔY?jì*�&R��f�PPS̚�� ��1y�\o>��}����մ��s��`鵵��)V	䛁��:+OGrX���OPe��z9Y�U�8$I]�.��~�~�L�R�(<ŵ�1������R���g����y�+��m�ǹ�n�&��h�l�A8��j�m�\��I�Rr|��ο�T�!���������$�����1XW̚�2ɳ�be�d��;�lﳒ
AL�}��Hm%����C,?*�a������3(c�,*)���'�:�h�j��0�:�Ϲ��s�=V�/7�F�;����'��(i���%$���~d��5�d�v��4��ؚg=�b���aXVe���5�`:���Jþ�
�6�d�=�L��6�Xl�>�
�L�a�9E�L���ߩ_9�`��u�~���u�ވ
 �
�J��*M��Ƭn�X�{��eiR~��rf�d����e��T�'�?�=�q$QM�8���+&}�M?2TY����4����@���TT宛��U��)Ge��ߐ�,='h��+&�X擉��CFq��O�$�TY��&k�� o&�{�J�����+:�+��?bE ���{�=a�
�[��/�7L^��<�˟l{��4¾��'��C̼I��7�����hgy�Y;��B��g�|ɾ�,?j����dѽ{z��Ѿg$겡䗖}�&XyP��>�v���{�=���������\���AgY�����y�E ��a����aZGVa�Y�HaiP���d��p�E&�*1M��y���$��2���a�����D��d��t��S?Is�����۪����� ��a��g0�<w�5�B��<��:�:�&R4{?�&��
�O��,�2���o4R�%b�� ~J������0�Fi�Xe�O3���Ά��D�G�n�tѺ���y@��=;��O;a�b�S/�*,���@Q|�����H)6�qN�ìϩ
÷�f��u0��;�gq�L�G��`V�E� ��?NjI���g�%�w�"ǆ��T	��>5t�Y�RW~�a����2M=a�0ɹ���ݝd�l<�m���;i߽��(
)�j~���
N;{I�O�z���8�W�&{L��G�U���G}�,�w�^f���{�=��LT��h��VT<��r��*����i ��=���
���a�8�Pÿ���a�E6{ج2�Ԩu��ؚz�d���=�/�~%�C����7��oX��� 1O�����ar�N�B����(��Kz/1']�Y\�'�`R��HF1����5�,F���4���w���a��K~w��1O��_w����B�]�j��$M
�ã2JCOm\ы�B�? <<�g���o�C�J�S�s���q�X�!��a�Va��擈Vu�Y� URu
��"����!�R����d�3�����6�Ʉ:�E���'�{���9��N+BF���嵫~���䃛%Oo��:�a��w��8���6L!����,4¦Xk�\�����Z,�8a�5�E0���ΦaE��s�R
L���9�K�p��_ſ���W엹�"���n��7���u0��x�,�O8I��ײe �:׾��HT��{���~͆����i �
Áۖ�TR
u��èa��ų�Ofé�5fP*T��~OsｿΎ��޽�����;��%@QG��N�H,<~�*O�:��;�L:¾d��g��Y�J�53�C���Rjw��ڲ��5�`ש
�*�z�&0��2ϘL��R�Sq�ު��ڂ9��q��6��x��A��a3�by�@�T35��&���0���:��`j���Vy������aY��s��m&Ь��`����rs0��EG�.>J{�_ǲ�W*��"<��,0�E0��?&=�a�a�a���`VǪ~������&��f,�u�4��cI<�g�Y0���J����h��v�(VMwؙ�O�0�����xͷ����aG�0"=��q&P\!�ئR
L�~��&�}HWe��I��a��a��|�&���2�A`d5�gL�T�����I��z�	S��`8�H,��>��K�w9}��ܾ���=+�%E�鿱�:���i';@Ƭ�ɜ�}/q
����1�y��)��`���$gm��<��Va��|ɯ߻�i�2Ws��̞���c�թ��?o�{�s�~_�&�uYP�<{�}HVV{�,��	�_�i�C,��E��,>aSe��H;��3TY��T���L>O2a�QC�K���&=�{�ù�R���ſZm��c�+����bGT�B���{����ɮ~����L�}��5�B����������O�0�a�a�]� �VT��)�2�wCF,X�)�d�ojc����×;�V~��/��ې��Cv	=L�5������7{("UW�Q�]��Zu��䶊Sf�]��V�x��}r���T�����LY=���n�?*gW.Ս��`��o7o5�c
��� �����qQ���\t�s�v*j���W�U�.��o��:}�/󩔛B�{�g4aS��{2y�N!Xl��C=���8��;�HJ�����fy�H
/�ٰ�i ����!��>e��{�4��R<`8:|G�TT��w��}y��~���0��E ���b��
�̵�@�a����oY�>M$q����4���ɹ�1<��a�6}�d��<����}��@�����C��̕�D@Q�lT�!VM|��b2�������w��|�1�e>dˏ���L��
�MQ�4�Y�f�k'�E �1`a'U����HVto��4�0�a��.�y3�*)Ә�0��j}�(i �é~��߼9�k����7�������O�gT���d8�����g��2�$��$�
�0�9G?`�a�
�4Xu�y
��X�(
�Lk��������\����m�M��4�C���W��C߿}���~�=�w\�O����4é�?3���E �y3ﱤ8�C	�o��4śN����'�I?!Y�P�[2��°��ଟ8I�+4fɎ�d�͆2��'��βT�������N]Vun�=���F_�p6�G�x�Ͻ��OM���{�M?��m ��<���1���P�{�!��+&��L�������*N�
}ڪL<d���b�y%zî}������z�>�=��z�=�?~ǧ��'�oY��T�f��$��%a����S̝p���'��N�����a�
�����S�Ag��Ng �d��,w�2�R �W
�<k�"�/o3��)�OVs���s}ӭ�T:�0�a����f�T�q�0��_�CIv��2�: s�2�W��L~9쁔P�J�71�IRq
�3Y�����G��\{#àEH�&77�-��i�,�����玲TU��H)/��,6���Æ��>g	�j��VL!����)�:���!��H}�\IX�)����pJ�I�+6�k��2 #���T^�wX������Ǟ*|���M�opC�ɇ�|�J凱Ey��8�`�Y<�H-a�>͓l���j�,+b�3~���AfRh�y���������ɿ������F	2W�%���~�?�x��lOQ06u��R����Y��(�3��6���.��곞V��Z������GG�����8Et�J�"�=���y����:�ܹ�����@E.�j	�{�y��l�Ά�pw�S9C� r�2�Ȩ���炍�Y�3����w�y����9�&�@�a�ܧ��&�I2�Hk��g�%~d��wؒ����>C)6e�͇XT�~��gY+2f���?8I���M!Sl�7�[��1�c�b��G*�q������X��}}'���Af��	�l��M�ؙH)<���cHu%�!SG}��CL��齚S�[Q��C����w,v�û�8���},o�����#�K�ޟP��@�A�E�h�Ms5�}{�s�Z	�J�y�|�%�Ձ]j?e+�Ϯ�������W�rGf��6GA��f�ڼ��g*�hū��)�ת{��̾CN�0"SfD�Q��*�C��8n\
l��N%v]VG>kjk���uܬ�z�Ua.V��zB�V�?�#\�v���L����(|��;�e�N(�v'y����	��{��V�Lӵ��-u��HW������²j�����ms7�g��u ��舞���-&\{�>�Sj�`N�tLhmz��nz����{!�淦cy�M9<��:��J&oH�"��\�)	qT��$u��⮍xR��@:"ؐ��q%#�3�*�p�R2t'/[ʌW]�(���*��qzVn\��uV���7a4@qr8+k!u-��,�9�� خxHC�e�$Py5�y\K�^��v�5흱�=�瞨�#,��c�SL��o0u`�Ŏ�8�u�=�#��[�"]{G�o���y�	y����8���y��а���+��� ���K9�ڽ���NB>V!�� ��u���<�TۑP��Ўz���ga �e��d���\�\�����j<ݣ�8xU`$���k��O�����(s��롢��T���rΧ�Fs2��Ķ���#8�Q��R�W +���x�0��*����M��U��/�آg?x=�kb:7���	��lS�r�lEjgҦ��8aPE�W�����8۷N6�6w�uH�
���7�Z���N����Siש4���D�̃RP�N��+_�eٝ��s�%�rKO%�At���7�Kr�P��$��A	ײm8T��G >K}{;w��!��=W��v���b���m�)I�ġ~3�O�h�s��źq1^yg`����T;�����������I���մt7�R�-�D|<*9�{�i���{m}�j���
�n�O�������OѰVы[�b�W�}���s�U�v	˿_R��e��p�Q)���r���������h��"�E���mC�W�M)5����XV��o�4��~�~�bm��C�Bc2�J�m��m�խ��ju�՗}� s�⯴V����f�ɬH�yH�
��m��0�xw�֊b�p�Lul�7��].50ccuЕ7s��+xf3[�h��>�qc,v���nn4��r'T$q��-#��� R�o���*�Q�u^����x� �@��:�'W�{+�h:�#��*�l�eA칳�U&���.,�d�c:���pٯ5c]��8�f�p���@9��s1�u�3�s�
�}J��tn�A}5}Ϊj|�����j�E�X�">�%l�1.��b���Ɗ2�G�g^[Ş�������e �(�!i'�N}EO�6�>�.z��1�'����,�����puڀ���7�3�0w�G4��k�K�.\.xR��]u]�炷�eiEO[<�=��	�P@�[2����T�[@�/J�
`l��"*��.aX;5u��$ۈ1�v㡥�ڝ!)���j�N��M�ŦD��#ҽ8�b5ҧH��v&g���J��1a����X��Vy2��!A>���&pE,�#Pt���*r��r<�y�~L:�u�/AV	��TLW��nB������w=��2�z!�	3�Y����m����%,�}�8Q�6�ェԈ��~�溜^u8�(C�P��5 Z�Շ�����z�<�uy5�w��
å!8���\ZU	��v6����cұqK�Uq��^\T�;�SZ�SS-��%��4S���n��CWp�y���V.���M����wfbT�	peKa.\ú��b6�[=k ��l�������D�i��L�E���ܕ��KR�wl
.Ï�?�=�S�q�K�(5�y��Sz{U�%��e�r5��'ճ�8pΚ�/z�`��N����[h����3vѻ���;�\�j
[��;9�y)#My�·.�΃�b�:�s���:�Z�4:;�{�w�yo֏{�K�ݑΎ����Weί�5��zQ:�I@>�~��T}�k㝹}�4u���Ar(���,Ѽ��m�]��s���io!ԚDw�quv×���j�pV�=��6:��+N�_%��Н\B�ݍ7K<1zc�N�� `=�X1[�qa�i�JT�}�{�}!��lKb�H�+�� �c2/&�Y���"�=�"�C��E�����͙�����AӞ)P���nB����o&>���k�y��$�Ū��'����x1`��-UÛ�q�3���`����ؼ-)�46d�Eg{��y�C`�����\����r�fVS�J�\�J뭡3m�V%:�P�u���Bu��Q�]�i�*"{=<�8�A�x>ln��G������$�n-Ao�R$*���:��2����r�S�}ey�|��v12�]���p;���;�n��h����rrዽ/y�I��<�oJt
���06�����u�|O_l/�`�L���v9�࡭W5C�.u���V�LN櫀x��e��/X�sE��=Z��Wl������6J��q"ӗ�{ֱv�e?�s�rluMW��A℮���x�:^9hgS�*>�Z&Lh�J�����˄��Xi�T d���<P�o%�T��k����$�ڙ-����#�TX��՛3R�uk�u3�f��bݒ�M��-x��,`���M�,���a�Mw��a��@���n�enj��/��O7���v���u,3�G�c��]�
+�ٚ"Pϡ}����HKw�6���O��TS�g�αN�|�_G�!��QL�FqY�u\�2B�/�����n�M�5��>�h�*R�1'Baᅛtj:��][B�[���o�*�s��-̻U�j�����r4Y�Rq6�@U:P�Q���j�;���]�H����Q���̛�밲^U�W���#�����3گ��Z�85�I�n�w�c��Q9�D���򢃩L��'&Q*�Mh^�9����VL�#/7�d2�)����K/�RW+N��ա��|�P����K�pj6k�sr�0����ͩt�]�����vU����܈[�LH�N�-��d�)0U��z�d�.㧟o�����dQ��6*�*�"�"�V �Qb��*��U�S6G��TF1dTb�b��e���Ը�.�TV**����1,�1Jʢ�QKAQE�,�Q\YqJ�E""2�QJ��5%X"1X�(�1���Qb)*� �[J��+iE�"ZQQQE�,ATT�j�2#�"�DUATTDEV*"�*�������X�Q,V ��(���"*�"EQDAQ���TPB(�EV1E��(��QDQR0U"U�
�DR[QT���",T�H���EcEТ�F(�`����PX��Q"�UU��1YQX�X�"*,V
���*����EA`��F
���$Eb �Ȣ�"QTEQ`�F# P��-ۥ��]�yY���x�]�I�N<�6�1��8˯u=��]�f7Pq�*۩�mFHu45r+tM�\h:��j���{��f�͘M�)]���QpJ�5²Qg\�3�'2�4m�P�]�0����"�Q	.C�Uר��J��P�gr���x1J���eAhu���ۊ�]��;)߄Df��ʣ�N�5�!߹��-2�Eƞ��c؞�k�WԾ�a}t}�����RV�}�i�Iz=�	/=�}n�ˏQ�����Ñjp&���9���{5� �[^Ui��6�#1.[۾������utZ�}Q@�Bz2e�;܍À�ךe^ŧ����tґm5]ʐ�<�O����|�
���X'�ܛ\��]O�Cv6H-V �9�E�¦"\[�rY(��}�ݬӐ�3�+g�x�#HP��')"t#}ET���C�S��d��;��*��͔���E�ڬ(v)�����z&����K���⫢H�r���-��k	�B巗�p��8Q���K����o�G[d[���l?]��2���W�QC�v�v.�SۯV���,<��u?<v��s�E�Cr�q�X�nY�}�B�t	9����w�"����م����Z��t0ayE��Ȩ�+�ﶆ��{�B� մ#���ZW9�ܦ+|�[��`��!圙��0I��dn����a.Y��⎃��Ă�7ê�72N��ݼ��x�t�-��;�0~�   �.֦�%%'�^|	���t(�!��%�G)7�l�r}��f�Z�s�n��[���y�U��1��`N��",k���Et>��WN:����L؋ˍS'l��cJGkP���* �!.&����������Dn��5T�;65E8�Ux
�l���t��t�}/J�\�+�~�X&H�C�+����c���7ʓ�p}|�M�PC��:���#���]3S���K��0T��*KipCX����@�E�ktNG�Ɡ�ח��EW���"���6TT&��-�ɭ�W�eS��ڕ��`�U��b�Zɒw>2�3�#b���h�d#.�hK��� �٨xt�^��}4U3Lq�j��״n_;s�<^
�3�����g�������0�����Ϩ-�nj<ͭ�^��|�u�>|{Jء+kʳD���(�T�"����B_�Pb��Wm����8�p���.�����E׵V�E`���*8W�]#c�+�p��;�Iw/?NwE����-��4�(�.hy0�P��n�fHie��
Ɵ�{	>s!����|����V�Vl���%���"����A6c�fb];6����ş;g��]���c�}��U��\���Q^��V�`;9æ��I��ot���w""3���W{��7h�S��Ծd'!�q��=�O�j��G
�[E	�*A����R��g4��>S�t5E�B٘�+X�Re@
����v��LW���	؞��EM�+\+򜤘���FȘb�0E���M[�")O=�#�f�pr;d+��3P��{P�ug�Vޙ���0Dd1R�<���<����B����3��q#}k#A����s���WT�ㅉ����jC��F�v����\�U���9�U�EE��=�~���s1wH����t�^�{2��ᰠ���>�<
�H����O	�6E؎E@�U}/�[��43(۵�bWZ�@�`��j�n}���&E����Jg�6��g��Zu=t��ǆv0��d01C7T���q�)�\9��E&}"�C�5�
�F�BeS�:�Ej��x�VU��	|OEE���)�E�멂���K@�<�I�A�>B}J��{	���oR���o5u���B�XKxg�ʜ�8ˬ��>�@Q��iײsFi�+r3{��W��3�E�lU��z�7Zn_Rz[H��~��k���} #�
�L^��J�ћ���Q���]�
��:��nQb,k�$�Iۙq�l��\%Q�\�#�:	��	b������Vg���U��u�;#�z����Z����꯾ {�79��Ε����:+`P���s��@�v�E�9�"��lO=�ӧT��s�2Nߟ�5����{&~U��·�e����7G�7�EO�.r�xY�Yda���l^��z�o�kB�Lev[���<.}hx�:X��-�N�����qU<�8"�w���y��]�`������%?ne�h�F���+K�k���_V[<y���o#�̝�/���� b6�g������:ν��:���+�h:�Q�UB�=u����ڕ�͖*EF:��|�B�%�j'�!��c�U8Q9ՊqUtu���Hgt~�� ���L���}d�"���U7�S��
5��\��������`���>�/ֲ)D�+i}b����5�ӹ�qxp�55<g5V9i�S�9�>J�����0�5�.d=������X�����F�D�sB�(�/zې�fP�[�S;���ٍrT
RzQ�GC�fTX��*gb�AK��A��]�}�����bͽ�ѠlF_��i��j�c�4+�銍=���gێ鋿y�׼t�◱ztg�=�'c�2��ZN
��]�dZ�I��=�줇1]�AF��9�NB#�]˕]lle�l�ε^�b�7Nwg�E-[��GaSV? =�ǘ��1��1���(����S��	M�9�����]�T��v$*���N)lq��<!�i�����X��� �p��5Es��8v���Z}�3�)e8��j�H��S�&�E�\%�ElR��f�)�W��!�/x�Åpy3��o���亄V� ^���j��:�]��P�o)o�E��R�W��t�Mu8���<xxR�Xy���T�'�&v;�F�;�jΦ6P�0``�^���M�u�9�FezM�eLU��ltour��kb8���XBχ�z�P�߹LJ|<��|)}�Y���9xdo�.b�.����C���3J>/t��d1�2�E��հ/�S�u
�}������m�z��Of]�U���X6/��1�3�p���aȵ9��Q`5n��c��j�3>P5뛙�Ǉ��ߏ�9@���<2�&;1 O�&'�@ʤ�r7���ߙW�`'���ڹ�y.��&�T�S],)s$G����nl���.�!���rl�}*�%'�5��肙��ʼ���wv�Zy���G/ke�5�ȑk\�X�%.5J���[�.��/-<���3�������\$OM� +�����T��է5:�7[��Y���7��`�֥}��#[/-�%��G��8�p�zS�aE��;R�ݣ择��� ���B}B��TN�y4z�f�D�F�ß\�!C��}4�wU[�U��8�
�m��.Y]Q���=�j�v+�2��P�rs�S�������UG��A�/�!A�������B�XC5��}�W�� Ws���"�ܶr����~�AOeENmP���z���������u��T���)����{��ޱPCt�i碡Ȱ�h���y����9�8(Bo���u�A(���Vr�qS��p�}���F�ʦV�^� m�H�M�j����YQB8F�z3��ST�['±w�Qz��Ns����N:ӹ��DR���]��OY�uB���TpMC�Ry	Q4��j�e��fׯk���npj��vr�6�J˩�7v�cE�5�(n�?����G�U+�w�
��+ ��㐰�7΅qlե��'ow�y�7c�2^��+�'f���1�8���U�A�d(�*C�J8��κ��e���YqLv��/,��mȾu0��4�nNMh��Mi� �%"+���7��:�}�J^g:���73RT1(\+�/��\�8ֺ�0�1�t4pWe���0&]ɕ����a�hr��ƻ�mC����ZR�5����8���cJ�� ���Z�䰙h;��^%u�)P4�JF�����:���{J�Vr.��+���� {ȝx����`���2:7j���휋*���7M�/g��٨//ob�4o��Y[��U���i���d�B}Ub��c S�C!��}}T؝�0�������32��|�1����	RXl��A�����PӢ��rL]NE7Q�yT�8���鷺�����Y����]�g�٩��Z���`'QX;G�/|���?�#c�i�k�>���Vt�Wn2+1�a[(���QRӯSA����Y�63ͣ�KkѵP���k�����Ô���@^w]�ty�sQ=�AËE[��-`�I� 7��_�0g�0xr�?!�3�Y�v�ױ�bX/0O0hh�l�L�D�����jܬЈ*Kޒ:�w�/�Gd�%wG��ge�ڝ~�^i��B� =����1�L#|R"oy�Gxb�:*�(���qJ�S1љ���PN�Ǒ�ڡ�ZoZ�v��+���֗P��?��)���u��Ɛ���s!k^�i�Pk׽cy�?_��'�e���tgQQP�PP�B�h�l��G"�tkͪ�HSJ��o� L�B�˰�3J����xW��vìv�л�&�u����٫&tmmM}��?��~|~�xk��^$7x�]��ꝝ��ĉ�ί(b������-e6����_Z��ϫy��,	���w�ʸc��Wc�`K�W�}_{]5g7����R������V;��겄�|(���p*�\�ǛCMn�j�2���������cB�W�ﳗ9!\�>ˇ.f�V�}"��r&�a�9���YJ{\���T��l�U!��*/�)�Eֹ��=��("Z��:�΅T��[N�F���Ә��td>EٯJJ�����s����>�B%��F�9�ë4f/!�1W9�-�*��4��pjK�!
�r�ᜁC�h�_�ڑ~ݣ���������Gc]e+�ӗ+8-����ޯd��#�<�,�#0�W�3��­Թ=�4��~Y�V�M����xDy<��j1á�>�BEl�8=�a�И����.�KNWL�w=��lNmq�e�Y#�����R�ϸ����;���W�:�^ȫ���:�Ϩ`�S8�.CE6�g��u˳<���/�U�cQ�/������g^����س�u3�+o�1��7˶̬�~t5a�=_��Z��%�{汕��O�z��
�)�׬�KpV0����v*mQ@"�S����/�+w��:y���%J�;Y�;]y�]�o�i��z�sq������K����T����'7R�pfo;�6���q�
�&OR<qeY�����T�j���f��N{{c���ÑXwP���Q��J�j���@�g�h@�^�MLu�BW�������������g���s�μfp��}���u.S�mt[��Q�t�~�_Z5�<5���t\^)����b8����'�(i�T��;t�~�]�=-�2��=K�Ј�G��*Q#�MNfv$"Fӷ���b=}!�ە���y;
9�̨�1�ʛX���R��+�J��vM���yD�m�|U�m_�a�1��(���:.BSq`��9���w�1��#���e��c����-�/.b���.6��h�+<A��rTz���X����ˇ���('_��gVcal�3��(��k��k��ygCެTUe, �{t�RTLPt�9
����3��qj�eC�:_.�+����d[�@DR�5$p�VR��E��S�E���I�u8���/�S;oMv�2m�oJ�Po?'WPy�/=*.���׸R��ro�u�И�K>k<yº�߰V�2����N �%)��}a��<��l>S���U�|)V�g�V����i�/\k��Ӡ��+n$9�w��*v!���fǅ��mZ��� �
�Y�x{�}CZ���[o&���'���>]��e���8�o#�����1P^P�G��9�ä�N�SSs]�M')Tx�rB�:����������o?S^4�a�O͖!��v�����հ�d��z��_��9��Fkl_=-Gվ��:=X)��'!3FŌ�b�$��E�MWBj��N�E��a�-TUt�N��os���	��*����xN���L��tL�AOg��޳�����9����:u7��q�IK^���pL@3��T�nl���.�b[$�U�f���ϴ'�'�+�M��5ٕ,��z�]b�U:�XH��|muC�G_M*�hP���L8�+GZ�ʀ��)K�(�'aJ-�:��;h�Mx�`t��xtk��X.R�>����e�G�*���Luʊ�nճ9α��@ =��m�nlKg �^�Q�z����c;wZc:�R�r����<A���T���)����c�CޱP[�sN�g��v��:���k���r�W���;��{���|�@4�ᵜ��T>7��<z:��n�n���J��b��	e��!�U�B�.)zuI0�A"�g�F�j��{+�Q�:��䆹yT"�%gT�zʩ��s�|s;@%ɜ	��/����a|uhd���c���te������z`�Gˎ�k�zҸEY��(K;g�Pg7��^]M2�x��%+��ON7��¿u�H��和�-R_,�@e����V\���sh� �.�K;-��EݾL�v72�;��X��T�O&3�p����t����V!�]��t����vU��k��:���]��>g�K7L���4�N����M�W^3�Sd���>�罞�o�s��jʴ�@�`�`���L��X��tȆ�f�h�����WUQ�^v)'�ϴr�s�T\�Cܙo��A��+]������1��}V��s��Z6;w^�$�Gx��W�#�6T(<:B'���c���%�4���^�q����g7����n5�dt��
Y��D���_K�T/���C�T��[8[�NWΉ�o��Z5�m<!ꧢ۔z���W�ou/=��� ����\8��Ɠ���ܫo^w6岌�%b��͒�f�_C�e.)ǘݰ��YW#R���� ��5��{HC����g�IsD����+8�m��4�&��]�0R��ա��w�l�-Q�Sn���y�/ 2�0���-p�z*BhOo^Yl�o�u8����TE���RWxiCc��*��o�e�J��
͇t�;�ǓΊ]��J�Jl���Λ�$�'�»�a*S�T�|���6Vn�%��+��G��Z㲔`���}�f�ܟ9�s�9�f}Qb'����L��3�uݴ²fȹrO����=�%C�}�q\�<��d�Q���y�*L9R��q��Ŭ���q��rwYB�LsH��/�M�E��7,5´��Cs5�������kML�#���9�i�D���ā�|�n���m�}�U�O#�C���k�荹� ��x�������og1'�1T����ka�Q3�����Xe��!yw9�ߝ�@��Ϧ�:	��R'��7��%��¤��rp��@��z�!=%��w��͉z����0[u��\��S�d�neVi�����]r��y˨H�ܪ33�X��VMw8��3i<��9����dG-69wN;-�LyN�XX�k�.������ùvK���}�(�y<��_� �{a�6���yWZ4/	Y�F���t{���0w|+�����܁i��O,��	y뜵Z���~7�䈣Χ�E��[��oP��[�d���:D��=���08�����*�(��Wê��=|nS�O;�XgR�<�R�<C�f��d��d��b\�vE�����J�/I�V��Cl)��>�z��3t����oB!'�����\Ⓩ�#�eoU��+�i!��n�K���`G{
#.���i��G`�x�[X��Ⱦ���2��ׄ5Queuv�t��;�7��0` `�0�����*��5���*1�"���"(��*$X��PX�
)b��21��b�PQUEEb�Q��UQb�EQTEQPF"��b �����U��`�V1X�`�1E�V11AX���0b���AYZ�VDTDU� ���*���(*"�Pc
Z��mUb��U"-J�TDb��1��F#X�DQX��
�A�UTE��)�b��FDU�Q�����H��"�E�(� � �+��DkDQUb�+b�TTX1QDDb���E�Ŋ��ڰ��� �E"1�TDTDVQPQH�A[lPcl�(�DUEF"(�QQ,Q�*��c#
+A�`��2>�5��y���,|2������x��/uŞ��%��e͓.���+���kA���~�xO.k��fݤ2b7��U����0���[����E/Ʃu}Ԭs��x�GS͌�����U�#y�	?]��m���%���_&}\%±.!͉��F(�>P'f�>��!g�C�08f����]��)j*7?s����P�q�f�jf�Zt�ly�9��\)EF!DV�K��1WZ�v,JPGH�7Rb�b���ǂ�"�Φ-�&��6S
�j����Rxe䓸�p�NQ�=Bŏt���)9ؖ}����Qy��@6�A/obʕ�4�w*xDBii��"�6h�2��}Ub��*rV(d8��|E�-��0�n����Ծ�'�{a֫�.�/�es�
{��uƯ����5��F�/y6OP�G@T����	����(��E��`}6�O��u�E��U��QX+��|�ko�
��4_���}�g�
T�ac�!ޖ6��X��v	�.��l`m�X4�*a�E�4�A|sr�5���^��W�n���V�)�UÄ��<=��cX"Մ�Ǐ��N)�*��<��be�0#�Uz㋝)�����q�aYu�q��U�zwP�Z~��fn�$	���WW�4g<�4Q6�!�5bʘ��{�tv�^_J8�s��u�%�V��I��:Ц9�S6SW}��K��N� p�S��еU3	����z��O�jŵ�Q%�e��0b��*��a��V�ɴ/��D��W��D�ȉ���	�Κ�+����$u��y ��j����J�F�_t65�R�4@��6�I�K�Ԇ"�H�>����>��T.�B��d���kU$�B�"z���SyxDj
�w�Z]C�7O�үA�<����"��k���k/n�S�^���]��)��W�q�5'B�� luUC�
���-�;,wjY}��D]��҃���3���+�mҁue�B�
gr}a�r��p$j�iT@Q^�k��:ފqE����4�T��ػ�Q�E�Tq�����C��}�p:�Iפb�r$��ʷ��w�����:4��MTW��nzxp��}�D>6���@�<�:�2�3�*q%�+l�}�Q�jX'�#gI�.B�1������7�x���DK�UF�gc�5�ge�4�;��*�����*�5'��J���Ĩ}�t͊Rs�(_��S11�Q2�=��^�wv_)N��/�Du�s�����"�{K<]#�`��3��¬k�3k]�${�!B���9�k���$�զ�[��'$1ndH�)D�t�!m]	����õ�6�q�����_d�~~yZ�)�����h��">�/�0uOf[7��νt4  vco/���0�-���yܫa���J�U�A�]۽�U�"�������y�o���'T�O�C�!��|�l����ч�Bb�uz¬�H_�����Z��7�b�'n,�]��_�p����ӎAv��<k�}/}�S'���v+��[�8+��n�vRD,2�*W/lyunf�yG_��n^>.-�)�s�r���OZ��w:u`)6/|��3�z�3�u(�o�&�T'fO@V3�Z�D�=�^j�یs��qp����+�Qa��8�!j��l>��/iB�q�P�j�/x�J��ۯ3}ET�uZt�)���U�f��"�z�@��Kٽ[�.l��ȇx����ؚ�
�P��8� �Bt]8P`YY}'1��ۓt���:���[(��X�5�!���|1�E��l闑=K�ЍPk�K�e����N�f+��=��1 >�ۑ�6�@�]^�)��s��Q~�����].�"���P�neM�V��{��[
�P���>.\('�5�9c��nBSq`CT�N��k�ʘ�ȑ����j�(���C⧈�l]��^����X5$�(_R���V&\<u�!׶}��D2�|eK�MI��dUcLwgSE���C��b���\$�4뷽��K%!ӯ�i�X�}�4R[u3��]�����4f����n�S�F��)�(3����:�q����W��Q�o��u3��M{j���`�����Uaţ�a$��(N��x6-j����� �BP��bf6q]St<`�Dy��7C�py3��E[>el�֩�}+O��Rq�
���9���<
�^�t�ア"ʧ�:SU>/&
��*���+uL���w].
��ɨ����$T\5צ�
PO
�PEu�9�}$�ܜ"z#�[x�c��^��,l{�i�g���,K����ϸ�J�����Z��['�䳎���ѽX�%3Ys���Ϗxn�!�3�ń����V@״vh�<7S�S�Mco$�ғ�1�茇�qɩY9s��օ�Z 3�r-N&��[���;l��%j�벵�L��t�1���*���>V�NK�-�z���Z]\v����Y�K���1wu�5��5r���M_Bj�f�P=3DO���PQBT�6q
�΢�^�b��\D�w0�o5�E]���k)�6r�N8T;'c$u�Š�u���<~_]A����=�Ȓ���I�x�8=��>t�
�*��-Zv)t�ܹ��8��V���E,��^���|�O������W|��v�H�x 3q�3��I�^&L��~81��j��S��]3�^yIV�������f��TD.�\��j�l!qU������r�<Rz���"�؟.d�/��e��l]�G9�\����D���:�b�hB�F���ؠ�Ȓ'�T}jٜ�c���<|1�L��ȷ6%��\�.-!y���/t���fiF|��;)�<�*�����T�g>�_�7=՚EA{#����ƭ��g�|Օ�i��h�,BV	H�T\GOB��55:9IB���*��m��3����>W�m�W!�e8�	P��=STR+d�Ŵi�+�>���/�d4��+s��>���v����QBGh�*��������]�^Γ��+�]{;Ү�k��voڢ�_&}].�qbZ�%�&?p�����z�wxd��_�.�L��Z�=<r�?^����C!��2��R��},D��A���1ƺ�]�^*ϵE.y9
�r�X*!0m��⣳����mȿs��eEBhV���k��Y��I���PMd���8��J�*,o�7��S���>n9�^&z >m����5�y�˥��J�E�'�?y�%e�����ѱO�*����|Kb{GW�s�&��U(�D�Y���zn�({+��D�wJ�M�ن�ګK�q[�����'wuJ����?v��G,�w�Τ�������|/�+�Z�w�Y��93l����{R�jp/N���AGk'rJ�~iiگ���1%G���z^����q�Q�%��.D�x'��y>��6��j�����xPzY7��X�)1H��\%T���:JP��+7\a��Z!C�Av��.��l[|F�C�3Fn'�/x��G
��]'5�g�Io�Bܛ��s1�Lq��DGJrf��	��'"}�Pӵ���/9S߯�+�ҋW?K<�zTv<�<�|tVT�\8LO���D��kZ��ǋ���9઺��f	⠬5�w3S���Șc�W��'��P�D��1������r���R�f�y��5���ۘXO$c����p� 8@ٜ��EJ��T�"�R"H����(���A<���ɢ���q�����~��a�����8��63�;j����J��򝸵ur�7:N�a�cG+��]�}�&veC�3Q���teuU`��CǇJi���̕/.�c��,�@�QZ5�Z\��_Nۥ��\)����6NP�R�H��(�U#��==Vfn�簊����j.k���ߢTs�z����<�u:e��f�V�Ϥ)��r6���3y�����E�X�I@���3���3�6O�`�=���f�0��������9�Ǆ���AJ����L=��X[+�-�W_���:y����tz�T�]ǫ;A]}�U�<A�P�]��۬AVJ��Fz�έ�C�V�����E��[���O�0�>�C!��:TT�v���]X�SJrt��ݍ�!�%�c����B&��T�p�F��7RT�~���0����6��o��*�酭>��xy�j9]��W>�,|m��rp��.��M�,���P��N�fׁ�K�M>l���s�٧��}��źq1O,�~h�fO��ԟh�{�+����n���<���w�U/1�}�lr 撶v�O���d��{��^�tBz��p�#��4�מٞwn�'&��bM��{�x��Ϋ���,C�r)����y��9�(�� <`
��tyC���[��}�C<7����
��V�F{j���Q�/� �@�ν��UB���	��1g�բ{����HSp�	*H�ٓ�t��u�<��y���q�Q`�D��1�ռj�gC�KU�p*���϶H��B���7�UM�:�:f7��ld`YG3q��]�<�C��^gZ�����F�\�8
�i}h�P��Mu	ܨ����fl�\���y�(T�w5�z�\#�����N�=�g
�sb�ݲ'�d:
Nm��ii�o�Op|�h�R?!Z�&�7.P���J]�GE�s����Cb`�+P���S9V�Z�M���Ē8>�"Z֓e�2˚QQ�-��̓��N]���c[�Y0`1ʋ�3���j)B�eL���-NKgL��OD�^��2�f7w3�*��gg=4�� �c�iđx�)6m��^{ޕ���_��3�S�
\ϡд.�������V<��\�W�t8���У=��&RaCT�7u�����v&J#"�&�����}��+�G�zq��oS�j O�R���_���r�2�㭹

������q�R���X���|��EUu, �|�8�[��(::g�t%4ƕ�u��>v�WT���*.e0�tEr�RGQ�r��H\lV",�~�
qJ�;����)>�/�:A�,E�9�C�P��u}�Շ�!:�/���ұ��� ���	n�^%���v�EQ�~�Mn�@7�v���C�^V��-Iʭ��\̛@�^��Mon�d�:�]=��F�f+���(C�ga�L�>y1]:�<�3Ky�)�<}ϼ{�54d�W�dW�N����]���)�F�Z�jDGaȵ8�*+N�����ˍ�ۛ;�p�����l�wl^�vr��mu���Y.�!�"�+�4:���:�]��2$mI/uY����%N%HQg�9�$�z)|R�0�ښ*�xl\7�VЋ��� �o+�}'V��[����WÈq��u�1n˾��&4�U�ʭ�~\M��M���[�yT���F��q1��Y�;�ګ��������_B֎tҜ=3@>�((�L�8z�Κp*OvR�r���U	�H���[!�1�AN�&�@��.-�����H�J�mtMx�#MTx������֩>�k6w���
B�r.��թp3�S�~��i�p�ҋr�FD�G�h���乬8���)O�s��c��$[gzTT_Z�g:�/<������L�sr��.%�Yַ�q�w�c�4J��U�фj���j7���}(���saNǻ8F��Q��9�X�8T0���"�
����!,$"YQq~����T����VMv��*+k�gN��h㖼�5\�S�N��A��x.��H�Q�o�<�d(���=<1��q���4tOBR�Pqu~㡚yy�P-�!*%}Ԭs�!��1�ƺ�v��3��݊#��兑Q^�#���UL�z��_bs�<9���>WD���g�~�<x-�h����8�#��z�!�妋��ɽKuR�,�{�&Y�g-kf����, �S�����Cl#e��#����-�:�W�R��.�Y���>���Mi��5+.����A{Du{[�XĊV�b��lCU����gW���&M�M]-w*�}���b#�����-u�z�������	��y:�(xJVy�S����i3srK�dÛ�7i��X0/����X����A��X/�!s��l��)�t�}Q=���E��<\��zi��T��"�p��#!��>ȫ�r/�%ܸ67M�/<���n׽�.�|BO��c���e��>.��9�9\�����T��Hا�U�-_؞R��Z���W�V��)]�#����Kڼ���fp9�e� |+��Z�RGԢ��žW�s�d�t5T�t^�Cr�S��a������U��QX*���<A���;+��@o�_n�v��C^F��W z�i�'�ɟa����:��j�+�}@Q�`�s<�z���F�u.\)�U�E�nDK��P<����s�8���\�H*G�):��frˠ���^V�ϰP��!��`�0vG9LtչY�B ��F��k��SӼ�Μ[
��qB��kl�@k	[X��<�P�}Ό��Co�ք~�a{��szf�X�]�fF�V2]�WS�b�i=ڑ�ӷ5�TBaʊ�j���g:&�ۃh^`H/)�,��ᷭd��pI\��DB���5�M��Jz7��5��S=a����M��Gd�}5a�zӽ��Z��`���!�F���)Z:y_лN�������'�l�m���������[���>瓯cC;��d�e�|��k��
���s�x������f�3�� C�X����7�6(P�ܲ^vP�Y�cH�tO>��V`��^S�QK����"f��aX^��a�:�7��8���ݛ��Ѷi�~�1��o�v����{��	wր;rC�ӷ:3F�|���S�	�fB��9�n�ف�ԥ]�3��[���7QH��ߍ��R��!{�1��6O8���r�d�ʖ������/��oW�'� [�=Լ�z#�=�I���}�|�PL{X#��j�a��	PD�C)�d̦���V��y�&��okg˪�{�]@!����$v�܅��eAN�f��L��xm*��`�9��8F��؜jJ�;�&��Ǻ,�m�2��rఛ�.V�L��E6��d��*�φ�[*V��#�[M�uK�+tD(��/��5m���u�gD��R���a_������TѓY��ѻ�b_UiG�S�Xp���:f�[gU�������at��4=Z-���R�YBv��7��N�w��ZYyܕ��-U��ޖxP�%wqǶ�M��ɞ���ˌ!�}�o�WP��=r'R�z�>�jԘgC\�c�pɚ�wێX;s�V�۶��j`د��<o��;�sI�����Ѡ��oFl�����pj����]~{�pv�JХn��2� �]�Y勝�B�i��YK�����,�pvQd-ؾ�}��#��
��]���,f2��n�Y��{W��Dz��F��a�_a� =�Q�G!��`h�G��N�����zF�k9�1R^�ˍ�A}���)b�>�&U뼤�`��g9�gP�ƅc�L��5� toRw}�{:�׀�~篁A�����<�Zd�3+�sF��h��K.�f�'t�eh�f�Z��9��_iڙq ���a�JR2v�v����q,�{fQ�:�͜�f��/�>�v�T&w8ӹ�'�dfʭ,��h��\�΢�fgiv�-V]��d��qqW�����M֋�m�j�;$b�l�5g5L+e$Jռ_�>�v-l�OI*��a��.�i�n2�G
�d+f���wV����]�����ӿ��q����^�[�WY������>&$��0���q㤘��vô�==j��&�K�*cZh�t����Cs��q���<�8Cu1���&L��7zh6n#S+e�4�J���ri���6�ZK[1��Rjγ3)|���^wx�N�tW���f�|2"��PE�*����"-�Tc�� �bQUDU���*ŀ�("�AAXȠ�*)�U�QE
�Tb�H�T-(��E� �Q���DUb��*
���Q�(���QZ�E��ccDEDjV %j*0U"�R+�bZQm�-�"�J�X�X�AQ�5,DE��V��D�b�R�ԬU
�T�1U�*�QQA���,Y�#b*J�E��"�*�"(�(+R(�b��Eb1Uej1�)E�DJ�V�"1����jX"�#`�Q����UDTQDPQ[J
��D��*�UEDU����-�]lp�:�'���}�쬠W��M��a��;�u�n3d>�����+��5L�}p���U^<���J�;x�`���^��~#����b�4�8��b���;2�%T)�
U���90��Ml�e9�x�f�K�X�T_�|xs������xxk(t�����X5$<:�yr�/^��<d��#�f��j*�U}/�mҁu`��WL�O�6NP�R�H�)D�ڜxt��n�w��T��GT��O��5+8k��g-rx�����EV:����V%��撩zCu"k�� <J��/�یLB.���)��(�f�_uq����r�B����� Ԑ��'�+�R\�~���"�P�ڛ�o��u�(-v�s:7��B!h�͚�9ײ�'
���������
TJ��7T͊D��/}k�.0��JZm)���r��1��6'9�9q0��@=揶d�ux7�C׻+����$���2���'7ފ��3&�!@�d�����3���������y��r��\U�h�7K2�Nqs9ܯ�7l�~Ì�-�h�?"������X��S���<@l�͗ ��t u�����N����l,��y+��@�l^y��<v�yeq���������.}O����/���Kr��wc#!(6�2GEυ�60�O&l�E}TS�yڕ+�`��>��ݛ��2���9{s�<��?(��ە�䵒�}�F�r�j(%�}�h|���c�u;��qн�^Qרۗ��qnr
ta�lr�����Un�vc�]���a��U^���{`O�AVA�	*H��2z�gR�:�plך���'s��$�{8�ԝل�;D=�/��À�e�yN����(Ss�"��篨��Τ`-E����0�
�s
j�8�'�ޞ�L���	���U�<'�q�B(��I�Z�����U�����*x�{Uc��J���2�]��t��D�Myz�����[�͌UʰĊ��.&�/]�#6mʁe�죁;
�{ezj�k�V�r`,�^��:�f�P�`l�"��j��%cx�(�X�ې��S��x� )}���S��L%]�J�R�A�TG���Lk�f���"5�(��+��L�x�:�]-��Ö�I�:��;�����V ��ʊ�X(��ۡ��C�^���{I�[�-M5�.�q�
�W0�y:pUR��*�o&�����x��ج�E�k%ܹ�_����8!|k����1�8�s؏������{}ȉ��W&�k�H7��ݠ&��V�qU�=�hZ�ÒS;ԯĂ�fv��잶:�N��;�Jgp*q)Fk��ri�b�5٬�br���,��!���07m�YK*�ǻ1'.ؑj���o��!��?Z�cQQ�r
����>N��y�Qp��\)A<+!@*1I�۞7�c�Wez����0e�=Ig�4�^���>�Uψb�ÁO+Da�U�U�p`N(ձ]|���0ߟ?��+Eט��رx,5��1�ر�n�oۥv9����;ѧ�`Gۜ�S)#N�W�4X�.j�ёC�3"�x��Faq�~δ-�J�o��Z�-��|�OLZ�������ޝ3NP�0��N����⪕�	�M���}�:'֗WC��X�R9{��:�C�!@i��ʽ��|��h�9��$G���AG�e����ރb{z�L�=������\�Ԇ#��6H-V&�@t�Ùs��$z�`��qj�ϊ��+y�7�9\�Ր��	�QU7��ˁ�"��b�]��8WL��9�T6'm���Gtmm����?P�Y��OD���ճ9α�� x����u<`rs��g ���xn��}�{�FQ�)W�4ǟ�W��wQ,v��s�G��/e��5b�#��i���38�m[���\��m���N����ZrX�<���
ݼ�#X�Mt�1��(%c �n�jSD֬G�3��6�Tu+r!u�P�=Z!=i���P�'-��s�L5��	�ܙo�*�.,��gp�(@������l�ZG���G)��>�S�K��"��x�t�eE��OW_Y��^ᆼZ=%l��ޓ0����l��a0���E\�YJ(AJ�Ө�G��,.���?7j��Ǆ�L���VIz)���΂���8�g���;7�j9Q<&�Q��ފ�{Z!a+1u�cN�Ku�c�9�U0͍QN/�>��X�%�	��Tb��(�+>���y�e��ժ�ܾ{g�u�z����\�J�	��'LFG��tW%�Ȯ�I��K�J2*��`���RJ�x����� ^v,�r6�X�Sʊ�'��I�DM�y=;��zR�}Y�aR�|��8�{J�!b�v	�E�r/�%ܸ67M�.�B�dm/#ӾE�Nu�u^�ݹ{Q]��F�hߑ3^�>��7$T��d8�v����ʨ�t�z8r���'W�r{0�,l��P[&����A�u\�ht7D�6�(7Vݷ8M�,�Q���Y3�R�U�Qc*�����Ӏ[=y�6:1����D��N5㰨@6��NE��9�Q559���g: �Grj���i����Et3�,�����wɌ:]:_��r��v^�T��tҦ���yj�ӉJ���W8���B��M{����Y�6�VB�����V)�f���	Gz�%V^�s[+Ɯ[{���O�]
�$z3h1J�ȿT�+���f���ڢ�`L��d'!�q�=�D1�+W[��[�6��f�c�V�BlS��B��]�{3�k
��Ǔ���f�S�z�*��ݬ�떪�	�G�b�^�؞�e��0o�_PN^{���1�YWu��e�Ӕ�Tb�b 䵪Hv���a�쐬D����k�ԡ&`����yQ�DM_`��Q�v��*CG
*�{���+��3^��V�R�z2;�����\�����.o&YM.y`�`�7��,k�r*)�t"Y���ٕ8�B�D�HJ��ݸ�����E�q�/��9v�4��9$SdX�Jxj��};n��.��L�O��r��p$Y��7Y�3��r��r��+���ȍ.���5+8q����Y��W7O��g��9;^�K����z�4�4v�p(�*����}��`S���`�!��]�NvAŮUo���0n;=
�D�r Ԕ'�r��h��x���s���M:��G�K��뾃6�Hܾu�MCH��6�h�wf�,��VoA~b3�
����Ȕ�68��D`�B��ӻ�&���[G��#��A��W
bD՝���%�ی:���:�Z���=�a�{��u�i��N$3Sv�M��x�!eN�B"��F�9����p�>	�[F� Y� ��ܗ��j\�X���OS��C�Ǿ�i�xJ��-Ӊ���j��<9�ԝ��J��{;^�9��=2w�=.L�u��T������;a{u�͕�p��ч�^�^��c+�m���;�f9�FK�+ko��b���_R�{�ňv�_�e��dҀ/k��w�<��H��#&J�4�ty}�x���-Z�>��>�qO6��:��ۗ��qn{��,�B��8�k�;r���9�U{&=�0)��zH�	X2}����0m� �3��;�YH�ͺT���Ǯ�c��vj�.̐e�[�t�	����}�xX��GG�ƯO�	��ޙޮo��GG�����c����� �Jː�8����9�.CP\�'u��v�І2�}t�@"���3�Uc�a��
��21�AS�[:e��蝂cK�cj���-��q��EŰ*�����D�/zۑ�\�����GC�[2��>9S��g1d�[3H��˧��ޘ]'qX���%�gh��~@�����Kqp��o���v�1�x�v�_[�
H��"��8�^<��LC5�)��J�\W�q9�S��ժ��k��xV�8$B�A+�5r�k1k��1vsS�����G��
a�V��h`ё�}H��ʈR2'\
衳g���"*���p����Qܱ�R`%&.��̚��/��;���Y\�~�w�6�ALG�zqI1���QNR�5�(�j��*�Z9�}�ڑ�����I��IQ��LR��Xl��+�B���(L��*�p\��0c��I]�x�m�F:�H�uט�5\ù�	�2�a�ʍI%D��M��IS�5�;UP��J�OVE��EKW�Q�����*1�C���'Hl��H���Ӄ�(-iq�p����W���W+�����Ya���<k��-���1r��y:"��U{T�]���:����sP���|)Yx5k��9����g�ۥ|�!�2�};�.��GD<#����B��J�@m��:�/�,/���Z5a�nǮׅ���H���K�15�:��������[8�t0ջޑ�rj8\�3^��a�╯	���*gޣ���=W�ԅ��5��vhS���p-�>n����_B�ڠ�	���e
�wK�<rCޙ�mY�@�[�ohv.�]{F_m(�t�z}2�L,��_��JO��&�@M��<��0�AmLbvGv�˨�%e<8C���9��,��W��gl�|�<F���̩�]�x:,@�E*e��wݰh���05�p����]��D����;8�����u�+����$�7W2���vN�H�J���4G�*����7\�ww�dd����lq�UM�r�gH�*���`'a¿S*1˙��:�]Mn�<䆩���ұ�Ҭ��Қ�|tG<x �[3��� WpîGE���A�-��A�	��5P���b���T��=)�4a�U�w��_��9l�҉�bjw��L]��O�r2�V��Q�^����;�x"�
��"��ă���C�GX�ɿ�E����o�W�iʍ��ݳ��}��rB�Q@eu��$H���K��������bب�5�zC�q=et]X��yy�Q�1��%D�9
"��e�:4�Ǽ��#�]7���ɠ-׉�Ҝ檘gTK�����"%��]`��Nͼ��κ�A�g����B����1�������t�*��ב�ކC��L����Rt�dM���J��2VG"�_B/��<�� d8�RJ��~^d�������x�����Y"��(��mqUgƲ�A�ڛz�Q�w�8u��;�m}1\�,�u�f㬚wZ�AX��������2�<'�u+L�Q�:S��}���M> �o^uՁ�S�q��vv�e���;T���y�����Z�ժ����� ���]/�����~�z'CϑU�x�m*����o�
Nv%�C��캸ѻ�o��Q��E	�= &�C��ض���T�'�V)�59 ����.�������oo���TI��K�=���{.�-���B�/*�j������4Q�TP�s���nΥ}�|�jJ��F�aw-��9W�z}���}���с���u�:��֌ZӗA�D7��V:��5���+h�S����.;�aJoj���z���=�w�7(Ɏy�] >eۨ��;�~��C�í��?�'�b��Nj�0�.1NU�`�B� ^�L�D٪s��vԭJ4-���jq�*��=h�LQ^���4�]�	����$�޸�r��r'ɮ4���R����w�,y�쐬D����k���!��b,��ܰ�F�>�XmƝ����xGEX,��ߛ�P�Z��{]f���8���t���B:�f���VwGY�H_l��.��q�S����/�B9n��&p���_8��M�mZͶN�9�*J��x��V��kc���S[���N��҉G�=�駓G�{E�q����uM���ru-
�Xv�	�:��j�XNl��U�ǽ�\�b��S��V��k�䚎Q7��L��@�q�{�˛���M�5�X� �pd�t��|b���ꝟUf^�}�<
�E؎E@�U}/�E�P.�}
�3�>��9BV��tƎ.x-��-U
�	���ʈ ޗ��t��(�%�9�S��|k��s=�toؠ^�[��y��3���n�QH�EP�Mp ѡ��[J*:�]��1��Cmt;��ܽ���o�v�.���HQ���O:S�	�N��$T�!]U�@n}����z(lqk���#��f�"�^*Đ�5'^�w�tnj���8:�[��3]�B�*n���,�h!��l�qq�o�_�h�bs�ŇN&+�,�~h�fO:��4K��&����輼�R��e���
��.n���CGPd��el�8=�b��"b�E���4Y���j���>��İ��ǡ��}�Ԅ8�ňw�� �w}�ZToQ�kB�_\%��[�{"��D��>����}�`}.)���ľ�9�h~r�V��,|V'���t+� �@�Yװ1:�������A�A$�5"��O@WJg��v
=���k^���K�h,�{��ˬ�E]�ꝍ՚��1w�ٵ������< V]�p�IbQ^��a������t�P�;�w�姂f�I槧ֳVx�d�q�ԏi�\>�p�ʤt!��k��T.oN�,MkI���^/<��|�I�/��d��%�#Z]4$S���>��,7��wV�r��=���-�m���U�24'����{㻺�D���bR�V>Λ,4�&ܩ�238P��I��t�@�L(�-}��&IY����ޑ+�y���E�ϛ�$��r�ۤwIsG}��?��#M������G�ӏ��=��h-��_�{!S�1��V�ǋro<�WFRL�$~��M8��v��6O�Te-ݛn���]�0��9��[S�Q���ԃQKv�ނnT���Z�cq���E�ќ���:j�{�H���<uy�QѹR��L����*�����m�t-���E�΋��ou� ������Tg2:��c.dl��^gCۛV\�_W}:��W��7Q��օ>�o��c"2Iqc�ir�ՔVl�EfI�c�u:�M<��n�0�m\��!w
�^�'Q�r�7plM�ݔ�\�������0���];�}dͣk8G�����)����mBp�����+I�m����;0'�t`�bgiƗ&�vW!�һ��Շ�Ȱg5���$\�j�c	��;5Z�Q!C��Sh�iL�ێ�G.��L�=�m��������:ѥJ�Z�+��P�o��)�m>��;���p�ڹk�&�[���ޒ��t+���վ��j9;UmB�����gwS�D��ɓ~4܂�'e��M��]&j�R�.?�=�	��`��6A�+=�"իq���^Y���m�q��3پ{��nt�*��&�!n��;QSvp�FZZ���nvɟ ��Sc&u�����ؒn^���n��0�_x�����g���\�7C�b����6��0�|^"UEx_|)���/D ��-���;DÛ9���:����v:BӴa�,��L���ڳ�ݽn�mm������X�]A��{�ς��	zw4�9�:�Djl1h󣆈�sN�ibJE���\R�k��e�s�%
�J��;xT�积��� ������C=F��-/�Β6����_<�DΣ��6r.��p@�S���E=5��4mnr��,�`.��5���L���������!���n�����P�ɷ���	�μ��akF����)��Ϥ��>;����_e��?iȠ�����1��>::޹/5|�	�S��	�J��/�7}�A۾\�`R��&��}V��V� =�{>�١ݒ��s��� �Y�w\Çy��j�z+��>�R�ad�j��9%d�Е$�hOjG���4vB�<�lh���Cw��m��䘷d�o߹�~�4��U�F*��L4QX�!l�(�*��kVE��UEU�*�*�U����-�@b"�*�"�TQAUZ����QV�T�DF#mD�¬ElbT�Ѳ��EKE*�-�YiE�*�kEAV+R�[J��JʪȪ
V�(��F*-��6¤��T
�b,UR�m����J�(�`�kP�+
�DkJ-�"�*ڢ�����،A�F�ՖՐD�B��V�V��
)T�TA*�DUA�+��ll�ؤ�KUU��#mQT�,T*+e���a[ ��FQ-�iUFZQѶ�j�+�JRԂ��ib�"(��b����X��VإQ����hJ�dY-**
6�[*����y�/?}���o���5s̋l�b�OxʗT��B��4g�d�c�
�o�ÅLӭ`�x�7H��I:���_cH,��Ԃ��;b}��v�睢���X�Wt����ˡM�X4�(�誝RԮ����75�iQu6:��ꚸ
5���1��X+e��te*�3�4
�O4's�����&�IJ�1��m�'�J�<g�V9�P�k*du�jr[:e��Vm��̚<T����u^�D��l#T�@�Jj�(��[r0lە˫�GvζeFs�1Z�q�Uc%s��V�~]@���ₘ=P�U�p���=
3�;jv�%7"��E3�T(tzyVc��FW
�~�Y�zKFWg�*u���|e"3ˑ�;\> F��{/vF�:Ǭ�ry:+���T<u��($S��7V"v�q"�t&��l
1���"�r������[����^E�kEhW�΄z�/�u=N@��ʍI�*&�Ss�����5�J�Gf�$�b���+ �"ԛ��.1�p&pn��9C%�H��]zLn�9�˶byRx��mDwQ�p���G���9�FezM���m�=��8P��kGe��d�o5.�n�8糟����)��觙�q�G]{Y��w{L��K�C+H]ݛt�4zk��P&��TOϰ,+;Fk^�V�`d=�b�(�c�����iS]�
٣o��,��.�.���$�V��Qܩ��8��[�E�S6����a?��0��Q�Ld�5��^���FF�v���ۥ|�#�_Z),b�硛9�φ6+�s{����d����*�M���𱗶��Ceb]7�2{]f�z�,p��6r-NrEE��w�#���p�f�:�7��qk>��"�����C�����S=��Áa�>w�U�XO����;Ҹ��w�G�iW
U~[|ȋ:N�+�KM�W\ٖ���*���7�B��M��a�\XuC�v9*ڞCk���6$�ot̏}Nu5XHgᇨ��b����Un\�.R����p��Q�z�q�}Zf^c���aT2'mp>�KJ�K�#U-��E��{�c��P��s��3�Ku,�ޤ��U�"�DZ����xW��4OEԠ���цj���j4|�ڃ�T��S�������4�d�Ҝ,'a9��c�CޱP@n��<�p��X,BUB�(1�uAG���76���&:7d.�b\tr�b���O�ΠrA)E(J���Ꙉr�*�l<Œ����2
��<��f�߽V��^N���-��*��l��"�㻾9��50 㳞|B���X4 �E��^�h�摍W:�꒚��j̠;�m��rv�T����5��h�{�:�
�h}}�(ot�2Pxg 0�LЁje�ަ�j�X��,j��N��c�V)�C��㛣�j�r%D�u���jN�v����0�;�Ve��?h����{���������"%Ɖu�d�,�hr��M��}i=�)+�b}�$d�˃G�B��;|ȣk�#׽������w0t�Or���;��[�y�X���,D�D<�@�Q0J�j�2��X��mȈ"+oZ�S0�<vxss��S�2⣚�t��j��SCL9��WBŏz7��Rs�Q>ɴwct\�ﶲ���Ӳ��fЗ���l�=s&	~�4�ʙ9C㒗�Z6)��:�r��m�����L����ψ�'����_f��l����ɷ�6jI��ht5��	��ә�õk����N�Qu8d�+z�,eS��Pb�Ӏ]��ذ�ӹk�)��C���]�x�S�b�XhVƐ6��
�*E��#f���3BS{T\����!9"��f��k������3�K=��"����(M�t��
_��v���S�9ų�9'�$��ꖙq��2��
ӽ�6L���mԺ�g�늍���^��Ŝ×��+����:/E1t�xgn*�Rl�}p��5�왕8c���x���9aao_�w}����.؇���m�G����nj'.��g��գ�<�}�OV��S����+�%І��!:��4}�;��9�!��:"��LT��<w���1J}5j^B �/zH�m�@p:�.�Hٚ6�(C��š챸�����'�LC}[{�=#�1ae>���
婘���M�^�WN��;�Nd�^�t������ݑ+�~$�N�u_)���Ȩ��Њ�~�ٕr�jX��8�;�ѣ�����ɏ޷������,����`y�9��z��_Nۥ��wХ����N���v��:j:�On��PW.�:c�QE��D���X��b��j�r<��7op��k�)Ԯ��O/���Bg�)T9^�A�C!_���Ҋ���n:{__d>�D&�v;�2�����T�Sa:
��lD﹐jHB}'ة.B�1��x��`�J���W�}חޯ���S��=®��Ѩ!:�C���_���Eg���z���l��x��g�l�
�.��_��nF��6'^�A�N&)址e{��K�(���8�噺�8�`ܽ��o�[=�.�*��z����=Q�r���dX(.+-�&�U7�|���[�F;$˜2�Z�X�0Pِ�r�m́B=��o�Y��-me'�+su{���wJ��ЉF���I���_�h��M�ˮ����n�wA�I:�hIǅ�LYt}��n�`0���sѢ:�Ga�6V́bac]CA��+lY����m���kih�hx�8q��gs��s_P�ۭ��;�r�X�L��+P�ը-���k�}\ja��u�q��2�Z�>�kV2��(��^Qٞ�M�N�^�wJ��jo�t,AN���`''$�W��u�@�%I"����
�>�l��3(�����s�rsG��%�Y��V5��~�� 7���r[�
��	T+ZT���T�1���u=;���Ƭ��3�w�z�:Jtښ�
/��y=�P�����-r��39:wb�~�b�^N�f!~� ��Db(_2&�����3�Uc��J���21�AR3k����nc]	l>*�i�~�q4�t2P
:��T�H��nFlە�.�e�Q��,���ږ�R�	lɎ[WR��1+ң�����Å�x�(���;����UC�[������0]si�@W��*l-dP*�=>^�S1�h��Q��4k�WII��q���P��5,V�eu�ܩ����G��p��6�Ǧ�V�����'0]�b�c`����!���2�v�S&`9�0L#b��[Y�9^I����Ws���'f��`�Ş������5�.�<�XfΐVi�%k��i����3;J'd�^X���C����`L�x��Q]�}~�l��6��|��4�l
���T�]=�,Y��X��8��L�:z&+��=
�����'N
�B.�tETjO	Q(�Ugm�`�[�kZ�oD�>�^@�o<�?���\�~�c�OyDyua��4���CF�k��+*���Q�UW��pVGA�ι�9�}�^�6�(��ۜ�>!���p+��wS�Msv��C�녖#L�U{Uq�`P�*t�J����/<dnb##wm����W��>{�ƀNz�Qdb�W�V
���NV��R���WG�$U���y�0��}Y���%��K:tb�|��v�S����j��H�95.A��pt2=*lVS�Pg��R�T^ۭ[���WMc|`�s;�M�*2e;Ñ�p-�>vW�a>Wе��4�=��4D���w�o;!V��޾K���+����yH�QP/�1߶H-V���.-�A��wl�҅ݛי�z�b���q�Kb�Gª6}S���ҩ^�V���t�r�X"�d8Cݕc����w9*c����=��������lL�LB�o+���[������4Fc��6���wE7����P)��X�7\2������XP��T0o�L��Q��D���\Ż�2���ZA]����i�� ���6*Cn�{W�c/m�=7�oN��:}^J���AN��K������c\��4��|�����$�'(Eiל���%Q@^<V�C�ȿ�����kP�:�t�:J�|���ȉ���m�eެ��7�.���?���sjv=��X�>n��<�p��\��P��k�OAc�r�]���
$�C�Ë�55r㣔��G'�a��rA)E(J���꛼й��i���Yً��T��:n�E\�M�cU�+���:
.�S��i��vy�z&�����vrB:�kѻ��q]�}���&�_��e�����M�)���5E8����"%����V'N�rX�r���������5da���cn����,�{T��W\]�D���S�şZ]�Owh�Sk��k�,T%�Rݥ��V8/��Y�����/o���RJp�_(���#�ԅ�1ÕtT?&��3�S
��Ec4�VҮ�bǼ��͑U��ç����B���A��hKN� ��5<����4o���E�։�Q����vR3�]����j�2K�m�r\�! K:����b�º�4�E<��2�sX��[��HgW�]y[����W�X�7|�j�����^�U�B]<�1�`,����v�څ�!�O&��l��Z�o�)~�e7nPjcj�Ʉ)W��:���TT	�jL���[�/���h����ޯ0������!��o�Nl�깞>I0{�����r�'xJ	�`D^Hؘ��)��eR�ƪCr�Sgo!7�lt=@hq��q�����PBX��Y�{�?*t�?���~d���ebOǬ&|[�+�#�p�c{��S�G��>���p4���Bo��@>���E�n�E���u+{�Xj�GE)Ǭjӷ!�t�
��OXG�b�^�H���HC��1)&5tO�s���</��c��]�p�p�ۼ�~r;$+$l�]�q������̪k�5��v�h"�"o[��ńtU���M���
���c���j�n�]H�`�q<vf45�"��[ˮs}��Ub5X$&�z+�z�NU�EE�k�����XOe��r�(uK�x�u�`�5�K��B ��r�a��i�.����OK�.z���tF__��B]q����W[�稜�6�@����
���ΚT��@|7Ʀp�n�Β�/=�n�4/�m1�5{��1a�n��5�/T��-\�c�$�)�t�����
<q�P��Uړ)�9��d\�ނ���n�]Y�7[r�۬j˲����H�����ݡp���/�F_�`[�3�����f�qH�Ysb�e��U�):�0�Op ѡ���**9G�}h���U�HOI�<�!�W��
��(�K@�<�X"yЪ�B}����\᝾M�(��s��^Dz��{n/'�m�sy��^*ğ6�AN���C�sW����r*V=����[��A��Q]z��
�+�'ڬ��|(��m��ps������v�����]C�v-�1s��y���fE��C׻�|7`رSnO�ʁ���;C�!�l���ۜ��ޖHky��Sm���~�N0�*�"���`3�m׬�!5w!�<����۷�����*=���Kr/dQ��D�P��0M)>��r�ƶ
4�__i�ϒ�X1��w��P����E�k6��|\[���yװ1:���^��X$�>��,V��U�j=(��u�F���T��{���O��P�y����_�Kt�R�����5a��6&�i��5ܪ�չJ��}�����ΫN��0 5��!�Z����}d��_�RȤ�8ܝ�Y8ûь�����*gN��N����I'���Ol4��+x�n���S�^�ܦ�,������Y%;G;5Nwݷ�n�ɲ�^��9,�.�
��(z=jU����SwFA�OM*.k����o��,��k&�C�z�2.�s�
�@�;<i�H�>�p�_QS�uM��z9�*du�;�۬�Id��4=�},n����:
uIUp�G�.\��=�WU�x���y�]���9l�C9X*�R��\r��P1*��q�CT|+�%�/��Y�G�
�{�7��ǖ�Y8�&�1JFt�� +��k�C���O���S�Y��������o���<EF�;8��+��	�
+����6pD�h��Bh+`E�.����ºn�Z�=Ԇ�iP��C�B��>�¸<�ЏC�_&\\�a��9Q�:B�f�v<ޛ��M�;.:�c���t����"�����.1�C�P��5�!��S����6�o1�,�Cc�1��4��@�Yu�9�Fezhnoz��ψbu��35'�g�����eo)�A���+H��ҵ~>�j�:�V67K>�rs�z����؎�#_�;_�/�X�=[��٣~�.hW�d`��*FAVNC t5tQ�+62wk��(5>[��ɧtF��W�e��!����Y�OH�]�ڪ���d�",N%�s�N���Q�=��|%5�*X���ho添[�t�>͍��r�Su�hS��S����\[(�fl=.�T@!x���:��ʎ�A7�2�V��j�T���}[F�B h�m![Kxv	s�V�,4N!9W#��{���4[�꼰��>0�8���[�tffo��� m/IE�ԭT�N)��.
=xsr!]�±9O0�y�0�F�~�Owi'٢p�K�b��/r��c9�E�q��i������*[��Ql������@uק����u�D��^�(ܠ���}�vj�1��f�bɛwn����i�VE��M;����`����i�S����`��F��Z2WN橼�t:�!���ty��_u$��<R�*2�^�,��ga�ɴ.�7�~V��+^y۝nh�G8~N�^$���7f��fY����\�لf���u<ۖ�t,M��ce�~p�孏e�'�椰�`�2�C��1�	��t����E�:DwK�5�+�u��i�G3@��n��Ft��SE�y>J�}��=Q�oo���X��d��Xv�0�O���L����c������/b����J21vv��km��|�|�|��r��^�YR�s��M��ﳬv���-$��<��e'���p��B�V���,oi���M�����1��C�v���[���C��B�\�9˥`^f˞�W��=��wa��ss��5�0*��h�b�%ީ��(�h�c�,�ŀk�u���9��kG���"ߜ;2#��+���l�s����x�o�F��<6�R[���7��8��CL��Y��),4S�I��� �4����<�j�Ե��^�<�0W��
0������j�����-��c���H�����p�x��Ln�T9��[,�I�M��5����xU]	Vj�Oa#�
���G�Ǧ���v֩�h�a*攳G}\��RN�=G�W�y�YC��٘�c��� �(�Rۊ�<����S�I��Ð�\���z���sŁ�/:�+xb���u�Cdŧ�WQR�et�\n�b��3�Y6�f���qa���]�pͦ+��7Ԍ��j�j<I�P��e>S�|ݯ����Mo�M���E*�� )����"�m۳b���$������`ո�C=Ǌf�]3�+i^�*�s� {N�}n<{:t�#޳���S�1<GI�����Q{z;���EZ3������}��o�?"�q�i����i�D����{�k�q�O�f�m݋�\���%<\�Ng��8�>8��Z-�o�v}�:і#����W��* |x�"i��������^���{���x��T j�w��*�5����d[����L8�o\�W�Wf�����o���5������JQB��k*6���id�b�X-J�[B�dPP@YR6ʕ����
�+"��T"����X�k+�QQ�D`�J�+��B�E"��@*J¡QE�jV�dZ�VT���
��������*��)U(�B�-,�X���m�0+
�Ь,l���ԍ����m�
��T*��)YJڊ����
��IR�mZ�%IR�P��Kl*
6�h�c[���J�J�ʅDj,ZȂ
Tm�ԨT*�mZ�Jʕ�%J"�B�Z%K�U���
֥B���
�����%eJ¨��BډmPF��,��U~��y��]����.� epX�l{e��CW7�)�Ư+�,��("0�Kqn
׻DɡF@���>˻�(��&�r;#���j�-BJ�lu�������kC���L��ו[?.�s{>Y��)��gT�;��߲�햄�^U ��܍À�ך�*�->Wе��4�=��<m]�c4���<u½�{E�6������.�!�$�g [(�s#�r,n���aƧ+w{a��)��ܝ���1������ �t+�S�K���S�cX"խ��z���o����3Ӄ�u,���Z૳)�g��Mx���>��8W�h	WD�:�EF�F>�'��1�������9��;���.y�;��3�4OD�
{A���[{&n������B���<����}(���saNǸ�������W���P�b�^ӛ������t�1�D���Y�u���^�z��&힎��p<�$��P����g�C��؈Ӹ��w��2�b� ��NH�D]ƢX��Nt]K��^G`��5/*���*脫YJ/���H�uQ���üe28��/�f/x�r7Z���s�~ܞ�g��	���*Z�7q������@nk���J�ґ�R���є2T�5G)�Fv�|�+��E[��5�	�h��N�9vҨ���
��)vh�ې/$=�v���O4�k c�to��b+r�Ad��hn�J��Or�l�5|���$��|���]�8eу�|���(!�f�"�����_2(�k�#��2v�Y�^�؉��^�쥊ꑕ;܌�N���p��N�\)EG�p�%^ᵫ���*3��b{=�j���E�*C�a�**
h3a�����T��A#����oa�P�c����o(3��O�4�\02]�AݢĴ�� �6�Ay{{��~���4O���xoE+�-k�kV��2�N@9#!F����%�=�A�Gfa��>+M����EI9�U�z�.?.(m�>U�*���Y�o��%ژi�.�=�wF�0�E����녙���٢/"G���zr���WT�a��5�����ej��k��[WkQh�|�;7<��W�؟
(p�S��_#}Iq��h+�ݙu�U ����IްQM3�9س�{g�F�Cr�!�������� ����/���9B���RUrLt��X(��<�/���Cc����U6���d$opxXw��Y]��G��J�}��57�UΚ���L��S�o/���Fq�\]k�-Z����eH�^�,+\(ԉ���<�2t��	�y�n��5��owp���6_�B���1��Ʃ����g^�Zf�y�u%X|+�����Z�o���֣��m�b"�&�D	I��s�y���o���l��@O(�����mU�ܪ�}���#��f`Z�	Ǫ'w�-՝,j�@�|��^��5[R�"7�j<�Һ��H��&�u����3��Z��r9!c���*��C��$F�u��7��di�׹�q7�1ѫ��s�MWz_[�6&�����j�QY|k��b`B�n��l�w��uMK����"�\R��hp�F�����0�LMq��ͬzҖ�S��^P��@��;̵�)�ԧ����\�I��j�ukU��:�� ��&��8J��v���[�X-�y[f�틯C�D�zzԢ���Q��
�Æ*s
��Wk�-�w ϻ1
r-.������{������i{V��k�0}vBs
�+(�y��깺�Bn'�Lj��X�Ul�w+�F:۫H㹽)<X9Wt|����GzW�b5�Y���%BbE�3�����y���(�	r��w)�sW�y��6l��y�Պօ���is�us�=���0�>DձbӚg�&��%��;��	��\6�8r�|R����^�ȑ��	W8˺�S�5a �Uk{jm�b�k��Τ�z˶S:�3���!��K���X�ܷغ8/{�:�H��9�j�i��4��[��>s��<��z�[[)i�V(oN����[&нr�)��/�I�7�M-`��W�K^��knIY$�/5�v��U��C�Cr]���R��֦��WV���J�]�j�i\,�ڻ[�I)в-��Z�	�;�=���L��Q�n�[T�;�}Hv^�f�\�mf�����3�ac�:�eX����4��hKGN��d�,U���uv �=�Wk�u`�D'��Y�!c��^��F��1kkz�ns��x衻B�'ы��}|ҵ��}/����
��M��Ż-���������S�h�|����M%�n��b7)��}�W�k���3��6Z8���nme�k��ChX�&��6{��_�-�Km�.[��c5eVJ�v��wW��t����;���������*��f�U@EꞼ���-v��\��'d47]_Sm�t+	}�{��jkn����sV�K"�3�C#W5خ�InOiG9��%c�u;��������O��4�T+�B������*�x�U�z��>=���{��G���i�2R�s�xԦ�4e$rN�44:�p���K����wD��*x6�O�{��9=h>v��Z���;4G�`YCt'0�1��R�[R���qR�L�:���ws�مXMq�����h�1<I.VlU���O\;V�N{��+*��C��,.���~z˰��ս��g�Iex-�֞�^z�<�S��%����Y졕��\��k���٦�e�S�Ӥ���n�M�6�=�}��^��8�Iج���N _-��8���M4�&�Wu`���x��fвǳ�w-c��v�D�ܡ!�RWE�M����bX^[���\u1��?k��s����5m��}4u�Aq�S*��B��1�,���d\VWhyB�5��Ț�o��0��w��Φ�y���X�jH�To:ѕ�]n2u5�9���4���4Vo��۩��Y[1$�}de�.����������}'x���:��4���G�7t�mു�.s\�,S�u�aSw�[y��[%]�O�v�S?uri;�{Ƶ�e؆��\g��l�qH�kY�����>�\�U�T��S�i�+���B�"�ö3��n��wD���#5[Bq#_+����uO�	y|x���Y�j����y_1Ñ;�&��1���H��u�D�7[�Q�oڡ�+L��[̺ݬ�s���\�
�W:�hj��g\����<�#��i���;�GE-~E.��|����3~Pъ���'/�D_������1�T)�g�)��Sjh'�)���k��hu\1tF�I�qn��M3/�:�o���k��{�c��|ۚ��٢8­�8�Ȃ�T�8|-ʽT{�A-�g��i��T_T�>˥��!�Zt���|�sx�����e�i�1 pyX+�m~��4�X�A��a����f�NV溯�O��ݶ�d��z��:�&eCn��Ǩ�/U���]W�,�l��/���n���ᮢ�``��&N.�+u����88��;5�����U�]:�U5�fئ=���P��%�J�>H��P��G���X6�Y�x��}��X����Y]ݙ ����Eu��ӫ���s���^D�(`�-�T.���	dM��o.bo�2�s_c6Q��l&���e�vn�J͍��
t')%��W�����]U�榟,4Ս`���g�(�W��o)��z����V@���[�=I1��B�⯶X�)��k�~{�ŵn��Jo�T�\ѼݾZg�~�3���Q�r}}k��U���-j9暎�/.�5Ì܍���Y�8�9:9���@K	T�X;ܬb����UO��w9�z�F����Bا�[r|�� �/oW�4�vĶF�,G^���M{���8�z毘�Ŵ��D��n�F�p+�(K��?v�T��s��&�#�宗gI/3�5s���e��sbk��^A���^��H�7wjN+���li�Ǧ����(E�[�MP��a�����,�FS�V��V=�=]�l��֏X1�G\��d�������ptu��kfi������A���3�MUU���×���O�(��]�뛻�&l�5�)���vp�2�X�O�yu�@4r�R�	{؂������6{���$@�^d��9�I��zQ��ʓ��tg15��s/\׍�{��8��a41�:���5��������ΔjX��b�5|�(]� ^;F��[9��<&��}��i�E��5}��5�ݳ�|vO�3CC���s
�U�k�o�w ۤL[+Wf^����+,0�i�=�y�2e�\��{�A-�2��E9�t�1]�!�A �(p��|��[+5�ɮ���	Z'wS��T=����篙�J�vkjW?d��Ƣ���-�a��/'}]~͉�Ȳb7��/������Z�x���_RV6i��-/kv�&���=��<�
��՜mƓ�.d��lXn{R��.2��Vu�^��T��u=R�ZQj���W:�lpܿJ�
J4jM�]V5[Xa	�&*�}��ح�(N1iC#Z��1����P\j�zR�;ͽt���;[�d�B����߀� �Q�;ihP�]5t�*)g�v�M`�O:T�l�ʵ��SplZ��bA}l�ai�L��r����F����[So%Njޜ#�L�����.;=��@���
����������L�4!	^Ѻ�ѻ�v+b:r]��nJF4q�L�N�I{�iV ){z�4������c69q����1�����&5�]��Ղ����W:9R�V��:f���)���l"���X-�#W+���G��?K���F��t�[Zh��)�w^wg�(v1P����qI�oTub��j�KB��B��ڛ�e�u	^!^T֍�9К�V(d��׏m�{�ݎqM�y�=�����.l�cWQ~��#i����ኀ�x�*�Mx۴c����u��pr�����q\�Z�	��<є�\絙���Y9��^���'��j�7r/�!Q'v���3�x�洽=�ޝ�>�0,���yo&��ȋ�[zѷ��Y��V���ԃ���¬6���n��٢,��Ef��NTf���nН�<�S�=��
ʣI���X�[���K5=[�:�c���e]Y�Y�%M{Lf��:�)�jt�:[%˱��:�Gp.��g'-B�J�c�,wƠ�SG��a�����5J�L��\�+����S/��Vtm-�gmC��\����͖k�p�2�L.�9�^���O��ܽ�m��M���:�p�S���*����ؖ��7o�a���b��:�vt7и.�:Z���J�ؚ��CK�o�I�l�.��@�6�Z�p��+�
 &��k�=���&��	>"��WF�iI�;|J⭩:��Vɝ�[X���8�8��ۗ��6$:��S��F���hgl�r\P8ԟ|��W���M.�c��]6̻��U�޺���j}s��$b>�qάF�+�mU���V_qOq^��,U��S�kP*�Cl�g�P���Um	�H�|�j�}|Һ��e�t>b7;+;6���e�5B�"�
%P5���"cu����y��:���<�\1�њ�]��O�$C��ʦ��F���]�Cîz�����:mfsw���e�]�\R�N$&���Eu<��`�.���F�]�޼X�ַe|�--|�zН%|�o�QB�+R�\��ճm>�<tF�H�dޫ3�N�}������
`UIP/k�8��_��ĥ]�.�Y���%j5�]<�Dg���薝Bn��)�g,1�#�|͛⭗���
_!�Ww�YS��>�:���pcն� δ*� \��)$h'Q���� �wOSx��n�(����/�u���W{���: ��VuY�����v�'x��5�����=����}&Y���3��9s��l�5�ĳC�F�h�䙝�.��Y��r���X�b�}�٠:n\q�w��$�]kj�����6�U�5wi�!��i�ʑ5��K괴��]Z��ݭ��otb7�{qd;Ç�;�4Ύʯ����7J���e����/�(�\�5�x�w�N\d�iK�p�K�P.��[�3�+)�;���F�wS��-�H��w�+p�J�>cz�lT
c��IV�uw��՝��5vk��9#O>�����ҏ}n�m��ϸ��ⱚ�b�
]�Wg""W7�)����� KP�w�y�� wt����U�sat��}RoU�C�h���U%f��\���zS�6����*�N]G]�0�V�s��������9�x�P�]�"ZC��N��";}ې�~�C�U�3�pL:���>����v�\����䘲#�����������7!�e��E�;�UI�S�c��1�����G�����{���՞��d��0c�p���p�����jp��ul0j{�P5��{e�ѝ5?��<B��-�ptᎮ��eq&�T�]���YFt��]�u�K��<FV�_���s�4��8��{7��X�t.��Fv��ǋ���R'��b�6{PW�Mm����դ�v�1���<���as���i���;���@��H.�����Γj��v��ҎG��8�����6��Z�<�<��y3�
ٸ�X��h2��DW[�G���T�]Ӻ��»os	�C��y��tκ�<]�/y}���M��;���G��oHd\��Vm��5�w�Vm��k]�p��+DiT��|�fT���˞����s�YrgJٻ�@���cD*�NO�̛,ڋ(��a��~*6[.�q����3�\����Η^-�p��*"����)�>�=}���i�l�L>+�|�;sz�h��lY�H�+)ct5ɯ��\ j�6!��<�i������W"�rͅ6��0J~��1��>����"9{��M ����L����� y0sb=.2�h�-]���e��\����$�v�{�1��S޲ǥ�
��Q�-_9G��{��TA���r�L�����L!]�P�w�Pvv�룝��9�~�9���%��#m��V�`�`�������)lQ�R�*T*,X��#F����-V�"%��E
�6Ő����dD�hԥ��dm��m�F��EIF��"�m�B�E�X#J�+D�����(-V�ZEQ��A�c*Vڵ��IYYTA�P-�m�U��0U"���V����QB,� VE(�ZQ
����ik-�*#*��-�V�F5[R�J$X"V�ֲ�ҌDX��k��i
����TB-���*	U��6�Q�(#Z-�J�lJ��QB�Z�%ITV`,� �ֲ�����Qb�d�T�����B�ڂ����"�E���J((�����V��DH�������"1����V�V�(5lQd���Ŋ-�Z֥T���
J��dU���V�X�Ѷ7��]뎷�odr4kj��@�^�i�'�1%�*pyd[��k�',u�aI�d�	:�F���W/y���sv�nWA3���h۾7�[�p�y�4����\�'�u�Ӻ����k��_9�ݓ�v��+f��A߹�y�4�m���*�o�����j;/�Ucz�0�����|[����t�6��W$�{8���=p�"۽�#�O�,��m�b���}c%ژq���M\�7�ӂ=;Vr|�~�б�P5��WK��׽򨗶L���(�"��k6]h�a�v��i��'�s�p6�U��(<��%
r�w�;�w�+/��GS	S{�Cf��`���q�k��zX�h�0)yw���9pk�RU<+��(�&���t��X(��O6����\��3Z����t��n����HH)E�&��U"���~֣�K7n2&R��l�P�-Φ�����oP�5N��P;ܱ�x��R%�)Y�;N�|�B���c�.��,G����=Ũ�#k��Ѯ>a���G�B�UE����������`�w�כ}��4P��F[�T�{;��پr'��|���f!�w��.oA�N��y���*=,�=ۓ֕��k��]�P5l͇H�v�\��Ѝ�ۀ������VЖ��帧�v���p/���<�4qԙ|���y}a��-8��1\�h�2��`�7��ŗ,<������;`j�kh�K�w�6&��q#�,P�I.�����z�9�:m���S\�`k�]i��.P���ȍ��`m��A��ڭ����?`̩��'2ښ7����o�KR���Ͱ�"
��m�2�Zޗ��68c�5m�^U��x��-���اSWnc+��=+8-��Ұ�#�y����zs
�V��a��wXUj�Z����A6�CR��-/Oizrk}�'�`o=9�X��j��oo;oB��*$�Lwv�ݪJ�l���f�#8<���fGbج޴�a�C��]����}y(.�M����)�C�����u�6!���"fŸ�{`೯�Q��&��s�W+^�Y&˩gj���ʸk�4��ՙes��xBx�hD����(�#wb8)��5Vnh�F%����3ϹRt�GVL�m�0eǤr�k �0�a]���i_�<}}�\�:�%�G��[�wC2�`[eO���w.�2���a�O�9h���f�{�4R�L9����E�6u&%�Jru�D�܀�`�$�f����Β��F�/Y�'/��.A��`j{�C�������7�����+�q�x.Qcss��gd�P�ԭ�εq���S�؟w��P\j�JQw�yiه��e�<y�d�����U_�K���c��Hʸ
|��BCK�dUa5-���~�T3���þ��ڵ��歮��՗�=���J�#B
�}]�+n�gv�<��m9������ƨ���+Xh�/����1w-^U��h��e(�dNt$nq��S@�~���T3֚3r4���6�2�V9wOT,lz�]3~��F��k�]�[��Q��o�s&��d��S|��sª�-�Mhc�ur|5�ׇ\1g��;��q��o<���eR*�.�J��-�ݦ������(����Df?���~+zz3��K)�zɑ�{p:uC7B˚���^��y�o���{{�*]{8+�� ~҂�w��-�@�~�����A�p�N���j��=*��f�X�8t�,e��ۗ�.�4rN�44:��f6��~�ϥ��/�[�+�d�o3+z�u�G<`�������ӳG�N����!��FsV��Ivز����*��"���=��>�¯ͮ!�[���i3��[��q�z�Pߥ%�*ǁ{x���F�WG��Yv[{��!щαi��wK3����z�bh+��%��_K[��v�5S�`É�����ٝũ����_��G��f��U�����	МB��o�L�^t(�ͨ����!��8�by=`�M\��Þ��]Cr� ��B"2csI�˽λ�,䫊���6�:�_1�����ջr�]��`���a��v�ꇅ5�gRU���VCq`�rG�ګ�.�갚Dw���o�f]��E��e'SxӍ���_0'DUl5V#{��V�Y}ʬ�S�U�t��7��/�Yp�|�wt��sF��e$�KT�E�G���wƆǶ�8�[�����aJ��5�&����#�!6H���i��b�-jV'�z$��|��/iu���M����i��+3X�7,�8�>�D�K�(�ɍ){DNh�0/���C;c�%����WH��{H|��������G>��+�:/^s7U��qF���ʭby_X�pI��"�AD�1@��Ub7[�&�*2�a�|�m��؎�X҆z�h�KV���ʦ�(�P]��;����lF��-WH�
�gz�1�v���Ʀ��ȍs<8*�h�MU�[�ڸ���r�:�tܛv�h�f��[�p�6���Z9:���T�WM����"���v��'��Ʈ�.���ln����@m��p����H���΋˟^�h{kR�]ʎaWX��a��;;�gݘVN�0���ؚqV�kgRģ��8�6��q����
U�U�ʠi��A�[V�aY��ܱ|9~oJ��>oV�׳W����*���Ջ-<R6v�DC��;o��*��K�f��&˿2������^D�lp��[b�p����[�6�i�.�a��ʅ�]GL�Q �܇�U��x���+{;ڙ��ݛT��Ѣ8Q��}��`����X�]l�E��ΧES���c.p�4�Ҫu	�u�gsJ�ȣ\���{f�r*��ڂF-κ�1S4p�B���|�������Z���٦�X(��s��Gd� �2�B�Z����^�-�h_1 �G�Ā{��Ԥ���ֱI�Φչm���묞궣B��J�pt?5C�S
QGyɾ��`�}m�Q��x�x���,�ct��"ߒ�93.�#��(uw�'^�:R��������\��۫�v�l_j�e�)�"1���TH/o@iL�l��{7����=ۜ�'�<ZWW���y|�]��R
$1T�j��4:��Ƀט�[D�:F.x�k�s�MW	}m�������T���NS����,�W������"�\R�	��4�v#!o-Dg(�龅��ۣ�)XT���g���7����n��)�Ժ���3lb���|-�<�ƚ����Wd�ʆx�����>{Y�ޭ�7ڥ������'vE]kC�B���I��]:e��coK;�](���<�`��2��8)��=g��kv�d��Q�M'[s���<:sAU{cL)|��K�G�Y�6�0c�`�����w��e0�tğ���Y��綇�?�ɴ��w�}�v�%.wv_%^���Z�]����ْ��,�X}�O+M��]Џh�T��˕Ӫ޴e��b��/NMuG(`o[δ�����G�jrh����wk�����Y�^�^Gr)r��B���>��H��ݮ`VR>�K��X�o]4L���L�m���vl,��q�u�d�u)��=�w��<��.4���Mke��N�[�T2UQb8��f���Y�o�^�Zؐ(nT��P���}JO��o:KT�cz�A���o;9�nj��X�jM����d��#��	A�����֦".N#":諻ǐ�8��v��	j8��V!��q�>�oB�U=ܙ�g\e��O��=���֓�uW&����HʱJ����w5b���_-�IP�%�DƮV�k��i����Y�+�y�D��j��}O��ʈ�;Hl뚭qg�b:��۸3����J�jG�������j��n�,ۧ% ���W0���{a�-mA�4D���54�u��j�W�UFү�}o��o�bN=(J��\��A.�F�,n7�Y����[�GF�hb:��-�ЎעY��Hƈ��qk�cTs�ҵ�-�}|4a�(�Sw�P�I�p�gP�:�8b�H�G��Rw[�P�}~�W��5:��{ݯ�'QgЬEΦ�(�hn'�H�n{ǶњM؎�k��$���;�GR��R�N��Cë�5��ઽ�Kǂ�o�&�gc}E��\9
�/Þ^��;���מh�>h䑬���1)�v�v�Bq����/�:�o���}�f�u��--/Oa{Y5�*���h���w9�ncxF`�u�z��_w0�fa�ϩf.zU���l����L��MeC��
�EX�F�y(.�E�Y{��%VK]�F���]�ؚ����z��(;�*��7~�T/���;;-hU�L�^�c���⭎j݀�e�vo%��6(n@oD���H�6pU_H{'{'�#O�8�8�V\e:wX�=9����.�R�ۭ��B�b3��W��j@S]�����2}p#$��\.��k�'��J�_)2WR ��X�vVڝ�T{+FD�)8a��Q����7��0��ɓ��N]���tV��.S�e�/�{���)ri�j��=,VSW]^��'hy?[�`��c��Ñ@��7�:����`��.�m�^˿F¹���\��{�3����7�š$g�ByE�䏕�T��I�o��޺�7XCm��%NN����z����ؖ����[U`��W���"������t�5K��[e�Q�X�hAJ�*�����Lk�~��%��M��nĵqZ{)��J���B�"�Q !|�5��;����^買=��im�v�C=~M�jøv"��S\H��Mv"�x^C���v#ag��=yV��/ÎIt�6z�^�	Ąзp�F��1����ةQE�^�Y�l^��|�����U�mY�\6�{yb�X�{���	ڑt�����ҍN�/�1W�3�����^;f��A��6��݋���i�x����1+yޮjp����{*��h�7}��>[���ɢ{��Tm��/m���0+�'U|�J'u������mJ��ܝYV�����X��t�$��/�R���������+�.Lz��3t���/��匮����I�@9{
ި��试���٢�P��NaWX��a�-�����P���kw��\X����������18P�J��V+*�i�ʹ�5,���ll�v�:�������2����ս��f��pyc*�ۤ�=z5E
�����RW3���MX�A+٦�&˶S!�vn�J�ؑA�mL��v)j�nws�{�X�sՀ��7ԕ�f�x6i�b�&���\��#�wo�{��GY���H�8�t_��7ԛا؅w����J���~x�^q��я#�U)y<63��	A�$�y����U����s{&Y�+��3�N�yʕD������2�6'��%�N�(���غ��ht/�/��_,)��2�:�ܞG1��HX���,�V���&:�v�2X,TV8Xݍwϩ�j����:���Q(b�l_#ۖ���)���볺�f���Ζ�Mm!��^��b��#'ra�HM��2/;��}�:I�7{/N7�������:�+�m;�QHW,�E���ŉ�9�]��b}�wD�I���5�C�K ��o7)'z4�|�d�]_c���y�862���FS�A�ښ��>��y�ʳ���sF�ύ�r�Z�t&�$b�Cif7��(�|Men���tZ���z΅%X�� M�,wf��u�<t�2��A�|���C 9;U�<� ���]Y����([���*�a���c���P�7K��8��RI�ۃ03#�)b�m��;�Y�Kë��ۘʣ�Y	I�uX�Ã�G�.�e���s9�o"^�4�Q���@wK}�\�WX��'�&��4�/����5�f(�O�Nɤ��-�K)�HwٚN���ep���y��C�#�C��S��'�|Š/0��R��4��nܥo��'jc��b�D`
��,]�)���pc��<j�}��s+V��԰C��3��,�T�����w9U뤆k��.�Cx�LEF˔�=YN�ޗ�WF^��"�ڒ�A|T�A�Oov�2?OR|;h�z�/ ���{��l۔��{Ĺ'��e�^zk�y�qh!��ö���I�� �0p�/{�b�/�s�W\�+`��MYx�h�N��'/V'#��1\�ۛ��`��nȠحǚ��L��.��V�-��,��(|��2�����H}|��,Z�̿�Lw��fS18v�A�G�:�u�.X��+�����9����NM���O�Pr��K6?	����`����I��L˝������H����I:r�,T�hJw��ҭõ`%�]壪|���Ń�q�v�\�&��:'�V��Ř�	���#m��N�fŵ�G���(�v��\�3�]+X��Fxj�^���K�O
ѧ����ӽJaEK׽R�P�E����:�S_Ӓ��6vK��@���-O\d�^�'���_�oz��q^XTd�.�tWO�C��[N$:�]	�GIB��:��i���(a���������^yf�����������n��w?��W��[�\VBV����Ȯ|��5g�C�k�<���Cn��ˉ&���&eǮ�`��S����Q<��T�����wwX`+��׋���/��50������}a7�8�C��3�y�<�=�炥S��s�:P�ݠÙ�S�<^%Y#/;7`8��
mJ�ՙ1�[Y;%�IU�����2�E&�����S�o_���3�e��d��r��ԥ�m����{�踲=��f��NmK�)Ɯٔ/�.�d�[�JN�3�	tށ�y��G�V7=� Oy�c���&�Bg��]�_m�:Bs��WwhB���ƛ�ܓ�$���c����s�}�ƍ%Ae�VJ1e���R��Qb��YYZU"V�UJ!Q`�Q���0�(�	P�F���Z"��RF"ƖQR�`��j �UJE�-�"��cJT���`��UjJ�b�E��֢[*(+mPJ�őAA`��Uk)R�0UAUemV4�+
�Z�P`����,PbŬ%IZ�+[,b�EH�B��ȱcj2����+�E"�m+kI	l�"�(��k��TQj��ʈ�ڕR���R�V��,����d�T
�Ԣ��@`�EX��YU��+"%e`�U+iD�m�J�b�U*�)��+�(Ȫ�"�1��T�%�Z�
��V
�-�kV�EQAE�Tb��(�X**EUX�Db��VJ�,QH�[b�UN0Nj:R\mi9����%��K��@�F����w�����K.��_1�4�6�k5R;|�`=�ð^�7�-�WPӟP�-�j�z��ߵs���D��nlMsr�)K��g�`�d��lu�h�K¢��6?x��Eߵ�.�y4H������8d��]�������!�T׸lHю��)9����ѱ���8� u�JX���&�5�r���=E��5W�F��+��]��T�'[���C�nw�����N{ ָ0ޠSs^xw���G3:�u9�_�����g�p��OkȾ�D��_vw ���kK��m�����(�]-���*אپ��Z]U�e��)^|P}�w0�c.��il���&�õ�7Nj�(޷1�+��N��������}c%�5�=e�e2<��.ݙ��kP�Q��{�X�(<�.��7u<��.٦�Ĵ��h������{�%���XZs-c��z�����Ho�!>/�ԧ:�on�%WK:U���܊C��@�5��޴޵k�vz���d��`����{>�&A�l�I��H5"��S�	����WM�_I�wTI/W������bg֍sܺQ�w#4�:63��'Tj0/�ճ`�����׵�|�h�&+E9ܻ Kv�_Tt�cX(����Z��d�����HA��e(u=7��Z�yDN�Ru󘭓,E�^�j����=���&lO{z�(.��ǎ`uu1ɤT��4���X��q�~�mU��UZis�]��m*��g�E	�@��رj}��� � U:̍�]���i����Z��]=��r]e��9�m�f)���8�(l���F�W�9�4� Z&��坻����uBܷ���-(8�!��#qA�5����#��� ��s۽��j�s�|a ^�v#���������InK嫲2{u7ׄ���;ȧ�qOm��Mv!���k��ኦ�<���ة�y�'2v�E~�ɠm��-���ܻ�u��5�����ء
x$�G��gg����5�a1%��J����y��6��=�ޝ�YG���P7�q^�)U탪?8�q�,<�'����������1��Q�)���΍�|Q�q��P�}C�A��ڭa��g.�9;�A�-�duo��Vm�Q��^�rbΩ�1C�J[��lu@�k��=�E_8{7�y��hL�}�����3��i?��y��oW����{~�~mr0�e̛
)[\3u$z�,V۽���
��)T�*�eQ��X�Au�E����`��2�����SJn�"���=X�z!N�W�T�젳�?d�3����7z���\:�Ah\�i4�i��g^h�U�6(nX��*�T"�B=w�q�=���75L%NH�S}�1\�MX������>72]�6�8q�N�5ۅ+1X$����RE�N�]�|��}�5nܽ�6�z�UiM��8��у��F�P���;�H�[U`����H��c��Ȋ��=]��䡬[�Mw놽�r�DUmKD�ܬj����TZ"�5f7jf�֧����|�_����o�R����5[S���CF��ɑ5O��Idh������_2e����HX�R
�bF�E�.:_v>,WuӲ@��=�E��ʏ	����5ڵb�u@i>���S�k��m2-N�`�Hv�aS��^.EZd����Áb��8{*J�Fyl����n�t���-h{�<�s�6�L�|�}/I��N�b���<#2"��ǟI�n���4��h�\�/���ת8��T3���2Շa͉�ʦ�(��N�^�ݤ;���ϛ}�#�S��[�]4m�ކ]�]a8�зb��u4�3��ۊ�u����ݯMn;���׍�cx�c�S6���W��ݧ}r��3�OYE�+zX�S@ ��R���a<��i������d�@�W��q�kal�Ұ��vh�q��T,7Bs
�V:k�ltqv;��TZ+y�V�CXo_�\u��oof���yb����y����8���q\��5�K�50��]��ެ��f��<P�H��Unfe�8���8���R�����>����j�e��|�;7霝��N�9[,����=Ze�U����})p٦�{f��`��d9��Y�i�wJv���^h���)���Q>��R}HI]�'��7�%��
�u�nPJ�� ;e�O��9�G�!�M��\r\����ܳ @��u;�r�г�X�����Dm���NN�����t�л���.�#-��ؕ�'�4���y����c���軆F�ף� ����2�e�7��>\ ͕��.�Ӄ�c}S��\"j݁�z��LO�Pw�ﯭu\��eߦޚ�Z�9d�,i�V�G=j9�^�.�;���A"*�JQ77�%�x��۳9�@�;�WS/�U��S�Dc뒱�+��C
�uy���[d��VX�ā�j<�Һ��//���g�u�����ƆHZ���ҧ�Y��⫍\�j�;cW;Xh�}n���Oy1�������]F�T�z�qe'T�=��Mk�]~Mu��*��Y��OT,lC�U488��i�w=�̜�o��	A�:��&�f���UJ������0��k����ʊ��v�H�w{Et��N���6��[9���<;����R�:�� ���KÕŞ�>���B�:q7���=��miz{Kӓ]Q�s�9y��SA�7���B��I��.��Y�K�N�3�E�IYgv{:�w|�M
��}\��P6�B��P>0����s��QNMX��1��/~�|���(a|��T<UY�uݛɱLW:;�JA���v*�ug&������c���\3��P).�X�ҬVU��_gs�2�����Y���j�����5�R�kg��Cr�V�:yYJ�_\ �:�X�6Src�Y�<�Sר-<�]��������͊8J�NSvO#}IlKml�S�QX{��ڌ�����h���/�R>AE˄bs��SYB���>�Oi��;��2��,��呡N.`t���\����xD:��M]uz,��l�$_e�����%�0�;�ɴWV���E�4�W�sҭ����J�Y��+`6��+�E���\��*��-����mU���VH�{��-#+(��8\@{�۹�F�h���BF4j���F�.���Һ����EKOhI�{�e[�ҕ�Μ��9ث�5�Cd�$F�W�9���V�%��F�m:�Nu#
���}ʬN�Ny�1P������;��B��흉����=l@tھ�)t�ćN3������J̨#�Gs:��Ҧ�Fp}�w$&ȹ��skvõ�o�wN�1̕􄭬p>6Y��QA��4�-��v��
����[v2��X��L�M��]��=��P�}�����Q��=Y�b:)[�P�Zh�h[�v"��SC����X(bQ"GC�
��k)J*:uY��+w�)����Mw��H�S�OA��ka��w�b����ywӀ�[7�[�6�G=��P�~�uȚ��A����\�{��.�0*�v��0�[��\��z|��U�5V�\B���U�Yit�͚cLp�`J�0�Ƿo�(>��� vaG��U#,7w��5��(�c[��Mw���Y�U�2�²��c�%�x���wJ���͡e�ym%]�7�{_L?'c��Yև��'e��?hO�<}8�1W5�)c���j���a��s�����V3bE��K��j��֤5d+��޻�S�m�馯X(���-c��#��\�]~D�R���^=�<ƞ��-)���:��|S��m_0{GN�O-x�Ω�y	VX���^�J�	���X��T�݃]N��vr\�0ΐ3���]"je>�Eb�S%�����K-xD��s{'����-���^^��S���*��u��ֶ�!�o���G�)Ŏ�d�V�w����G���TOF��/Z��5vR��~�PЪX\}T�	J(�'�+j�����Kv3�9w}� ��ߟ}�2�hY�K����~�+���S;R�or�Z��7��d�-��^��e�Ք�|�{�]\��PR�T��[��;EEdE�C,��۹�
�<����i]S��Π��+�$1@��.\Z�6So'�%�����5G���	�D�aۛ��g�q[J�)R��w��e��a,�p�_�Q�~ކ]�\R��Bh[��i���:�N�jX�X3�M<WW�-��{h��-�c�ڐ�U1��u��x�ɭy���Uʱ�ƣ�WT�Ъ�8b��n�^U��x���AЂ$��8�v��s���`c��pߒ;4x��UV�NaW��O*�ׅ��zz���كݗ*�W@��¬6��+j���uE���J��)�J�@y0��@V�w&/E4D��CSi��uf?Wy��b�t�3�kK&f�TW-��fƽZ���KXQsq@��K��C����ۘ����&T[�wZ�P��ѣԻy�}c�I�WjC�����{�t#�p1wAo\cnS<n�:�{y��7r�7���ja�t�{[՚��Ҽ���T�/i�X������J�H��=X�%h�K��,%�-rl�e2�f�k�U�+�f�����������X)М��G�ԕ��m��5cX(��<EVoN=�V�WJ�|ūY�o�^�X]Cr�!�Ɛ��(jH�)��kdV�{�/3�c���3�2V��d���:z�1 �ẏ[75z����T��8���6�%�j8��fX����zPJe��L���s���>X���V�U~/������+PA ��C��H�3��IkR{
�P�U]	l�\�z�J��|����ut4Zp��Lά����ԮQ��ꑍH�"5��Y�Y���2���جfT\�J�Z��H�1\�������"���@R���mUL��sL1"��U�UJG��������Q�&Ď��B�&�Zf�Q��hN�A��xlx2�z�gc�|L��&��!�^�JZ{V����Yŏ%�-�f�a��V�.����[,��I�^�:y]���v��#�A�ev�	�Y��W�;}�1D�YW�-��om�t��n��w��<o�����
jh��b\�u48:��M��y�
չ��[9�;`��T+�ç2��X!�4���9����:���E�ދ!�V�|�>��;b�+�}���;�}��������{{5�	�������0����Mژ���F:�ó��<"�����m��#�S+6�-�
��/�귪�#(��������N2�Ք��}~�Av�m=e�=��L8�x/��4��q��q�����+�)T�71�o�+٦�2���f���[t��1�[֭�)��;=�ֶ(n\���B@/�D��'.;eF�wwT�|�dԿr/�{��~�
/y+���J�#b}�r�Ӻ�\뼥ou�3�A��T-����������[~�4�W���$��!$ I?�!$ I?�BH@�RB����$�؄��$��	!I��IO�!$ I��$��BH@�bB��$�	%!$ I6�$�Ԅ��$��$�	'�!$ I?�	!I��IO�BH@�~!$ I?�b��L���&y��� � ���fO� č��z�T��%T�
$D�iRJJ��H�TU$U@"����
%@
$J%B
*�*)$�J"AQHRQ"��	m� ��IV�������4J�k��h"�P�	5%(�T*�+���$����Ƅ��&�*T��$�j*$&���Bk	R�6k)��	
�&�Hd�VڄF�ֵ�A$V̦a�m���UE"�XE�L���j�i��<  �z�jn�B���ۧm��mܶ�]�wU8�[i:�NCuu�F�M]]�ݛv��u�J�P�v͹UJ����;3�VwCMӻ�f���
֩!(�h�+�  6�t��l�X㹍v�L��:u�]+u#���;�]��7:Vws�[��:v��V�]q�VuC�U����\��e�k�	IZ;��.�ZR�*nv�3a hU��E<   O.ެ�+.�tr��J�]��#�Ѯ���lm)J�U8���v9�em���wu�N��EΦ;�(P�B��^��B�
 �@�
(P
��k�j�j�ٵ+ox  {��B�
(P��/{��А�B��/w�
(P�B�z��B�B�
9��4�۝��ΐ5�����rU[��ۘ�ݵBn��w-sJ��5w7m:k�E�u�J�6�5�QR�U��  #áZ�����n�q�eD����ڝwf�4u\)��V UW]�벪
�p��j(�th���$���:eT��$J�  �P�
�w]u]��tu��7Z�
�3�i :���2��t��hTP9��D��Z㩮գMT�B�tjB��ڒ�� =�o*-hS�5����@�D�-�T�w;g ����e\�U��;W�Ѯ�N9`::�v�ִ �\�m��(�R�]h��  p�m�/����n�*�v]�������J����[c.�N릢��\�u
5������ݫ�v���wcC]aA�:��9s[I$I��mTF��&��  G=R�7�W9-ɬ�n��m�n�Sa�uLܶ�N�n��n�UN�57Ku:붕ۤ�vr�jStw�Jˤ�wI�]���ʖT��wCN�ơ�.�h֤���V��  �z��Usu�:��'YQ��u��km5�b��
�˷[R���nJ�w5�v�Jn����-�Ӛ����ws�ZR�jJ�V�����eIJ� ��$�%F# 	�1��CC�  S�A)U4���@��2UI   �I6U(�0<R�E dd#EE�>qG���*9U%=��~W_����3�\�_���$��S��	!I� ��$ I?�H@�hB���BC��s�������c{���ѷ���Z��v��V��:ʎ�:Mk�nQ����Q�I��de�<	l���3��cj Μ�v����u�Zn1����S��X)��f�����utQq1�"vY����ݽ���-z�]��GZ����OP寜�/	�ǇY�m7)���YmSX l�@��A��Ւ֪P�k�fju+4e2k+2��ۊ�"��S��^�u�M:n}�$Ғe�"&��Z�i�)�9T��x�kMB6]���j� @�Tx)����9f�L�b��P֛���n�elz�C���w��H�cu�i'�m��R�Z�8d6�`]]]�Y(b��E��N��sp�yaH11�ֻ����2�V�u{0ܧj�#6��r�$�ς�7��e���0�� H�'�z�ҵT�V�a��f�2��&�Ne���n�$�Xh��wZ5ܔ��[6n��vjДAK���M���ޓ�;�-hx�g��9&0��bV1�Tqb'0R9Z(�dC�.�n+֖%+IV�6�M�[����9N����T��,���EV*4�2��*��!F/��w-GX��W��BAG2�7NY$�g`
��+r����+orK�5�N+[z���+k6��;qw>�4��;��\�Z5��],��Ƕ��0U�("�IY�qh�&S�V�j���G(LW���4����[V4�4a� �t�IU�$g�oKJY"64�*�Z�IR�:�sE�T������2����[���·�-A�@�nc��ܷ�F>"]�0�z�pU+��ƫ�!�*fֆE[�jʴ�@���r�alܢ��IIB�]EXq�R�[j�z+1�U2�7oV/4ۊU��^P��ܡi-�֪ѹ��V��cw��f�k+m��z�[�nn\{&8[Am��0`sv��مí�je��t�ܥ�ca�M�雲��̣�Ib�k���:V���*΂�6e���nL������d'��%�ܹW��^��z�IYX4�
��aEZ�����PC��!���V�DE�n�RזP��h)���0%kݧI�u��ck
�j���^��T�3����z��nV�A��Y֊1��5�����iTF�f�ݻ���i�8�M����W}�+�qC��N����-	E�j)��R����3t�������Pܥr��͢�V&hӓmZR�U�l�jRJ�:+Z��NJʱG2���B�=i�ieX���Shh�u��Ў�ˬVX���ɍ`�DZ̧Z5b�ped�CHjU��A�S�V�hXq\Uf@*Y�ĐX�
㸚�z�d�h9 OX.��d��\͗G#Y�j�l%��d(�.��9��`m��ݸ��MҰ�5�&�ƕ��V�WF2f�V�u�3df�`�-y��K~�t��i����%l�:�]8æ�U�+�u�V���&ƪ	.}v��nMg�q����Lc���Zj f�
�i�����u��f�d&�����^Ea�e�7�8`�pҼ��D��D���z˙mЭ��oB��W���YX��{�M��ǩ�YWi,&�����&�t���3��ohc+,��c��ĜmSF�t�PN��.bw��B��&�ݴ�]=�5��FѤhV���0!�p��1��&J��>�Z�X�� �bv��lԘ)l���01-���F�QULVv�[�(ѩ�b���̢#�zr*�J�Һ�n�hoY8�iP2l��9{Q#�m��3t4~�)n�!�ur���` un̽��@e�G���d����*��[�U�l���wd� f8�4��X'0+�L�S�@�ǖ�QY��J��pcy6 w[�⺺V�2c�DÁ�jV�ܲ���Y+.,�d�@:�V�i�2Z��Sfܷ-P�ٺX��FtP%���E��B�-v���0�]k�&F'�����f�+�.�!f\���$���4b'Ve-#t$�3�蕶��*Ԫ�w`@��M���$��mj�o(^n�R�e�+�C��+D��e����5�'�p*��i�[`O؄��0:���sCض'O�!!�f�2�4n�E��Kc/���Ɩef�pY�omN�M]��P�p.'��W-0�h�LeZ��`Z�Q�VJ%^���KU��Bw'��w�����l͗!�y���+�H�-nG/13�#���R��ëZ��?���%$V�8�nE�~*ڤ�@� V%���D���,�75Xƀ��{D0�a��q�J�d�u��q�{n]��R� ��4E�eg^7i��Ai��6��Ќ�FQ�C48ĬW�EӭiL/b���W���V䗇ɬ��tL��b� ���V�&�t��׆I�Z��.�,Y���)$ q�;*ΑhH�,�r�ce��,��]YY�L���,�4�N$��ݩj�(���;in����9�KP�ጲ��4��VQ/b,��3.��@[آ+1�zB��NA�c�-��NɳA�,'��p\�2�"�2R�<dS�b�U�$��WQ�G�a�02١!�u{i��Ƿy.��YX�8�ߡp�������J�(�1�;���IT�{ʳQ-�*5&�r��#ؑ�Q]����;�x���2��v�z�8(�e�ͩa�f�B�1a{��i넺�x�T�.1Z冮��vt���M/ܤ#.�2�[inS���W`�YZfVa�,6�wG �2��fL+5hLH|(4.�f��¦�щ�v�'IW���58*Z��T�T���!��Z���$ԁ��uS'%�n��C~�J�SַD
��V�.�ͧnU�{�Z�O�kp"�2��3&]���h�H�o4�%����3(<��������wp��+,�m�pB�ݩ�ʉ�eʆ ��X������اч0�܈�5�� .��i�&E(��a,��f�&��{P3����;I����.�2��Yv6�L�o5�e��d�C�z�"/E�
Јh#n���M����z�(u�R�����!Yj]:��v�ۨ�pЌ�2�ԭ���f��n�k��6�W��ĜS�&a���V,�S� [(T��ZʅYD4,�7PI��X�Ef( f���ر�x�%LV��]k`���{Ch:�Уo��3,Q���vm-mٿ�wj[���Lk T贱m���k˰�;ǗG/C�݈�wRA4[N�i���Ҕ&(*��юd"��]C/��Q[��褮�Ҥ�R�pǎ�^��PV٣.�v�-�ˆPMC��Z�-�osq[�ۍ _��m�jA�-�Cjn�ZEf�/q�C�x���^�����x��0*ӳP뱸`�/7&S��J�^�^��OK���g!
�[@F�$�&� n�Q������	1U�f�749�\�\JUԹ"�Lۨ��RqS˧�T�&]��mЩ����"�饶6&l&/#�֤@��M=�a��n�n�l�e@� Y3 ��k)�h�Հ��gU�h-�A*x���ol<�yJ伹��@�a͍��X+��B��5yF�mѴ�j�/�)sA��rV;�c�D8]RX���ӎ��R��eq�Wn:�2���ʹk�{t��Za���wd��7X�j�Хi�zn�2#b�f�o@�q�̖r賺�)��u0�&��6�d�i����MRen���^�l��:U�R�}&n��O�8h^��W	���z¶�T����+EʚMZ�6�5z��2�m�Y#٘��E��Ő˧YN��[ײ�D���\�2��'T�����Vv��u��ɓZ�MRI�Cv��`�+U=l��r�D,�f�GN�w��Q"��T�;.ᗕ�p;������q]��Z,ԙrR2�n��ڔ&��l�v�bxr�'�d�Vn�����Z65�� ���cc�d*l��>��~s,^g�c�ݯ�p�*�#���Ha[��ئ�2Z{Z�m�R�	��y��5C _Z�d�,�)]�60�R�-��I��ͬ�3^��<b'i�{�h�8Dِ�%��ln�7�U�j�6�#(�{��c��$�bV���F�,�%�A�7*97M)@,[a�ygm��p1B��1<;vR���&�%ڦPdг����fх@��t₞�G���C�e(2�a�mm�kF"���1l��S4hho[a!�R�h�jٳ��u�)�LOl�!x$��q*���i��kF�fCbVc2�S'��@KڼXC���Uvl��v64*f��͹j�mc��]4l2��w����%i�2�4�@�HC0U�m�#eas-�y�)#�c6c#�l0�C���4�y�lBF!¨�|ݛ��	���T^�u�P�JKȷ3�Z�ڔ�����t�Xb��fq"V�D�[wp�S)���ɭ��*�5� ��{b���E����Yܸ�Jq)���2!z�v��0D�pm+cyWY4S�J�nV�)U����e4�:�k";��*�٧>j���/we����E�h��OL��s���5R�[%�r��h����RMf�e��W0�[�mJ���m@q],�X�ϊ'��m]I�*AWYyW[Pj�J��v���N�;jһ��1�T��H�[�F��P�����t/5�R��.@�#���oQ���y��B��G�����{Wo�B��詀��H��:�U�V`8��j�i<��yRLn���'S/lbZɭ�h`���:~��<� �T�7J�z�,=��Kط(ei歫J�,�{-��B�ja���Tn�n���ͽ��5s&�ïCruv,X^���isZ�Y����ͻ�0�2�	�MIZW�Ӷ]�;�c��fV�;�p|ZkQ�)��Js7w��M��$�[��-a�@�f7�@�l�YK*8�'�_A���K+p�nd:� �ЛW�Ipd��V�R�CCw~a����k�h�J;n䆉e�u�U��ķ�J�ctn*�`�L@fJ���;�n��8�R�a1⨴`�,�R	�J�ԉG W�ad�+ˏJ,�����iL�wW�녭�gC�����BC̥�1�C����Z`ڸ6�p�3f�ۅ�[[��Z �͉��\z
�Qj�ɻ�1�#mc�������o)�v�峱�V�d�Ĉ)�ƥ�fP���D��(��貱�����r��
H�6�[����қƙ:�13%fa6��@�C@�u��ow0��#9���jq�	���4�i��#{��#t�34�j�O��[Z�bo"&�h鐡�<��d6j;��YU�z��B�J��Ym[cq�ߎ�Z\q�uRt�(���J���찠{x	���2���؟;Ag��y�P�l�P9R ��KQ�Yׁͽ��y�*fY��6*R������{���zS#��[�m�)�a̘I���[v-h�e$�9,�!fl�&h����-f]&`�J^ſ$#�q@�*�(8m�Z�܎���AYO�n^[Ў�����*
�q*��A�KTN^)�<� �а��.�]+�h;����59k#�.5g�yZ`����5,f7l��,�B�/r�G6�G�hmH	��[<mÛ��b*��b�ot�:쾉��$�Fe\���rJ5�t�Ɉ��2��Y0�6a���SVM+^K���X���v���nRٴ��L��V *�Q�x�/b
$�c��Ec�$��*E�]��,'kE�neS�J��X㊍��P!�2�ad�S�t+ۨq�J�QUv6��P�hedR�xI���D(C��q�:�`�Y���r��[Ah���JR���dw�S̛�0QC1�Y�.��ܲ�Xt�j�%I�WΑ�r2-D�f�)ԏԨU0whD1f7R0R���!8p�zlf��Q���%D��,�*����zQkߣ�D�X�ŭ�Z��sF�{D@��Q��ʖS_=z��oLq;���)�k���H���*9�*� mi�\L�zJ�N��b���Ւ�Xh�W���Ѳ����J8ܸ���pȪ�J��vmh�!��&��b�9C���*h����ZT���x�"���,̼�]-n����T(�O)�`�a6-���e��.�%u,L�w%*�)M�����6���nP�m�˽�/agrN�5��s�DX�j�7�<L�[���,e�㡂�f�������c���$3(�D�2d5�6�b�m"%f=�yqF��mZ�] �*U!�t��rU��Rml��dق^��
{�RF�2�B	`�̡"t�m<m�"1�ӽzwh�6Su �T,;*��S Cn1H,[)95�*-f��7!��h�l�m�@-95f�&\9����dZ%�W�4��$dJ'��Z���Z�3J��MĨ����5,�B��^Dn�Y����Z�+�����z�ݭ�Q֌�M-��Zx��W�fh,��z���f�v�MM<в#8�,3\��cL�!WS����a�����q�d�kuv��7b��K��k�.V��ԍV��U�[O�������d�n�j֣���D&P���B�V�cn�M�!��&+ Z�d[H�BT��H ���($��1�(�=E],��fL�J�Z�Cq0�)�	Ijюv�R37FX�ܭ�պ�ͪ�4[(��Me�(nAR,�+y/M�7�P�gh��ʒ-#jvY��w(9�Y����u] Q��z���(�%��Ɗ$���ù�Р����]�yv��,L9o0\�$%P�i{��[�[�
V�b6�-D��>���I���!�v��z�l�tT����s��2�8�Z]WO�����+��d�0���h$z�h���ne��n���`v�-Z�|bR������ɀ���7��utu�m�[�h hu����9��c/�WB\��G�t�Hxjl<'6{/�\ ��=fW�w'���4�-�q����M$�[�I�.	Ý��(���0LPvX]\5c�L�K�F7�`u��+N[�����i���B�Yމ��nj���Cw3���:ü����Z��LG��ƍ����K)j�h��-.��i�p���u�#������rL�޻q2 �ю��oX�idc.�	���&D�� ����h�B���N�n}4�(�1р���}�u%#��Ώ%��Cݔ�OL��j���e��7�:f�8��4�[��N���Ih*gu�19��)�s.����-s|�k��t�fW���n��VG��ku��V�jvA�
�Ԥ�����I!��m�3Y�i��<��[ռ85�f�E�9s�!$갨Ŵ��ÿ���j���jx7$����'�����|օ��W\T)>ә�� ��h�活����$�Ma�(���*6�
-g}n�s:!�K �?o������c�z2#�������[�;e����3/ݣ�����gf�'%̼�W>y��N)r�)�x�;�:���ю�+�ݻ(8J̻�Y�/#�JRHk���7d��[\w���-���,��VF�a=�mW0;��Z��k
��U7�.t��浲�B�x<808%/$�uc��̡<��t!�.�)��tt����P�������vH���)|��:�S���Y��vDD�er�{u�6����#�d�v�vVq���Zd|A��gkF�Fc9p��D���8�O'46���*%�VV�&�#v�ut��a����o!�{Ff�(��l.��ZcnF�9�(y`�g�ӣ�]A�{����X5�g,1�laj,#44���}�tX�R�$У*��͂�}P��CPJ��N�R���ͧ"�MN�(f���I��|�YQh�|��o)���;f��+.�1SP��9|��]���:k��e��-MwnJI��a�UXC;f�JZ��ma��TL�.�5n֦�m-̀걹M�.�G�K'hp钣�<L\��mƵ`��9�6+�~��P�o��Y2��ضwS�[θD��	[����O���������
�e-�b�V����mYp�7P*5rKt�X���Z��e�]N��ۡ�uJUqRf�jlVA��]�eC��q�}����㸐}�&��]�\	�]Dă��vp}Yn����^XO�!���Α��XgU��E>�xۻ���3�gP⇟7q�L��h�Q���ݫ�ݖ2�Q�a=}��Ӷ��YC����fmуm�Z�Z.�Ww}��;YG�v%W���u�ѓk:�wi/H8�;o���8�u�2��^��]vU��L��l��R�$��tw�53_P�4�,ܴ�>����t�O��k{�fY8����&^w�e��-��XN�R����z;�3�g^�FJ(6e�بc,R�H�6���CZR�{����\����(%_��5g�eѱx���J�����'o�y�\ÄZCU�U��;�"~�M�q��xc��.���5;�ܺ�1�u������9=�[�lߜ�}M���os��I�e0(�՘�__ko$�+s�һ�m�gs~.�n1�v���B�)�]���&� ����3���T��Jq�"kmw4��!qs�}�k���x�3(�+�][KhZYhqcot F^�]�x{��J��pz�ɱe��MZ<��w���I�eص���ז���:�mv�-*�p�@�=�δ��Hm��X����ܹ5�����aخ�ԁs릻R[v2E�T�T�Aͷ�2İH��<��D�8������8�JsF�y{���m�6I�kkC������_/�rK�!Ej�ڕ�f�.a��"]�/��h5���LJ��=�Fc$w���'o�{��]ھA����͈��=)��+;U��	t�-� W�0XuZXؽ&A�F����d<[*��F� �;UJEb�=�\�q�5fŊ:�ePb�'WÆ�	��Pn�c�]ǯK�)yh@�̜�'�X��5؏_>�#GRtZ:�퉜Uە�:��]C�0ϟ5=�{]�M�0p���n��MgC��8�	u�̰��nŶ�J��2�I��*f� �*�
睳H��%ԤF����n�n4F��5L&�^��\U��I�oZ��S�d�j���8�e�O�
4��X�-a`��U���NP�$���m�l
���h|pu*<�ul�ojUt��1�sJ��j�Vw�[�
�E*�f���Ȏ\�rb�����:޵�r\Z-�Y���u�|� k)T[$����"/A圹S���ro.�O�	��gA�V��,�;�R�+�2����1�`�3�4���:�d��s�˧H�8�_n'�$�OL�����Ρ�_��)�n�gM[Y��ȵ9ɐ��7]�"�IU��7��u����mKp8��+�q��帋Sw
ƶ�G�|؈\��g]��Z�� F@���*���՝
:V_N�Ѡ�Q��4�Ɲ������0�8��58�CJ����R��s\cP�W�P=\e��gܳ{��b�F�k�J/�e9>&(�O�H�S��:��kU�S�ywa�ԂS���|گ�Ҭ������%�%;�-y��I��I�'&��ki]�z��N���&h��}�z�v�V�i7t0��mntT�]z�� ȑ�8���"*J��М�t��B�"���W��G#�����q�����L�	���.)(����A�ʎ����ap��n�\���ժ"�����1�h��k��fky�
Z�'7:��3 ���m#RN<����]ݠ�z��H���A�:�n\W�T�g,���0*�����КT�ƌw�r��m[�T�S�nfԼ�S�ef�Ͷ;Sru�ҧv�y�	5�wU�g\�$��]jor���H.f�h�*��3VNT2�{w*8	�[62���jPC6;,�V�ԃ6|��xm)���r���%��q�+�2�d�ɚ�­x����2�|�r� ��0R�J�`�Kl0V�����Yz�[wΡ�nG����}�#�z��}B3:&�Ƞ"��!Ī���䑨L9��9eq ���XZ6�f�V��v�5z��0*̱t�k8�p�x�y��`������}f��tQ�)�֑�<=C.�3p�Uc�V�fA�h���*�jZ��O�e$��3�4wGV���ҕ�8VcZn���(�DziÊ���^��6�8��47E�9���[�Qi	���{܃�9���K`Ljк{�v:��4$�z��^gj��Ϊ����(�Mp�O����VI[O�Cj��(����5�4�b�ׅF5C�h��t��=op��]�l�2���V{ce��9:=5k�O�ʐ���E����Pu�yC��)��&�3K.�6�:�>��A:V���ٕ��e�� !�0�-�?	��&�@�o����Zʉ+�9�kW�M��"qH�r7M�wʋb�����^�Ǐ+j�k2�Ag){�i�,��᧫+��s �̪��h*��d��,p+����Ke��Y�l�'�%t
ar���G�Sr���>�_��?<)q���r�X�8�W9��+��4D�Yײ,Ҳ�ʸ��%�0 �U*[wj]!�k�#n,U}	�������*Aʢ�z��7W�5,Տ�ޭ�X���+�} R[Z�8������Y�[È��骥�>��W�"�َ�r��M����`F��zȝݿ{�H5�wPJm�P����KR�c�#�e��a����{�ܳS'(;Urt��K9䠳8��̋k��=��Vܮ���9��_*����*�שn�#+E��m=i�uv�;o~̚�p�9�SC�0ݓ:��m�B�b�*">�L�=�1:��E�����n���o6�n�MpT�t���0�Jf�\��ͽ�@X&Yuy9�%g���R�Ni�$3#]H>�-�T'�z52�.HPOM�"!��'4�swsŅ͢Xo/�y[vJM�SOE0�I�o�gn�9�+��g�ëkg*��I�[F|"����gs��������hKW��/-¢��.�w*�=H(�w���ީ1YO+r�mm�6�IQm��5�%>�����B8���q�F��vΝ.����sZ��C7�KU}�qxV�a��{Ԏ���+/M��+˓3��p��7$*��}E�6����w�l��k���#�|�d%�֙�G�������*H_L��b��$1V��R�X��h�z3敪�A�.�)�u	��)!fe�Ñ���z���\�}����2��z���ӟh��.�J�4;,������(h�� �X�h��u�fVKG�o��bɗ\�u>�:�|�	|t�.��'[��FC����X�pȉz�e��r��c)�^�c�X	����"4Iд������;-���'eJF����
�ܾ��=�?�f�N�FFnf�ms=¥>y��X��Ơq�۫xEݽ/D�C�B�4(РH��Vn���\����v�_ZY�◕�;U��k�/;msJ�bBFu�wÉ�-��n�w����a����b2qeh������Ȱ#hp-��N���e;hAl۩{�x� W�.<�	��cS�fDpiB�.��]�t;�+�=A`X�c	�*w[Pi��r�]��>r� 	]i^���VWE�лIf!��[8j��a�z(�6���T�r���w3t������:�7�m�Zr�Gʣ�9��-��o�V��Co��ser��5k{v�Q���lt7M�ZZP'�UX��Ī��F�oY�TFJ�4{.�r2w�&z���b�"��[{�b�;+�,�� u�]��q�9�#8p�JJ�9����m��^ ��N=��qE䩠�ne�%s~���h�4��r�5/p
�W��:�ug���7�I|�:�fq<�ޛ]�-v�RG6Q��ҙWM��WmIXz�w�U�Ӗ�nۂ�y�g4���U��ǧh<.�H���t���2��_^=:��Vnxa�pC��^/AaǴ/
y��on�;�9�T�b��w�����gGs��ȨH{/�����*;$��]�>?q�q�R���ȷ�c�I�;�KU}a%��t�:�e�V�q�D��0�T�>��q��C;.%m��Y�'G�=��s��1�$�s�G p���Ok	����5V�W3f63w�ҋ+�=�j�;	���tS	H�WXkm$���R-O8BC�������HԔ3vm�9\��-I\��P���厧H���gH�5s��y���A���jJ�U�T^K��spI4�eB�Ц���Kl%�)n�yc=3�CD��%����5����C��*.���(iΖ)%�O<��^��;��0.�:s+{&(q�r���x,�e5�
��B1�vR+���.�d7/��<��ݏGc�;qJ��"��_ur�O�\�V�
P��#��9k�CXO1��=�]sg����Ii&�'�$F����H�s@��A�DER��p�͋5|8>��::�o;�&xO��K�������,Q�-h��!�X%"�b�b�w֩n�h�V�0�sIE��ޥ�ɖDǳ,
����*�މ��.t����as���w9�!���|�
�̽A������$;���m"�R{%�u,���z�Kg�'��o�C:N�TﱝɟGK6�@��MNv��T�c9ҏ�c�� �*69u���4�n�]�s�\ 5{�]%k���|�D�X<f���Ud��"kO��� Nf�R-����ݢ�2�Ն�@!e�3u� �۾��zu�!�)Ք3�J�9|�5	WׅӁ�q��P��.y]{��Ȣ����Үj໱=�G�lk������E����m�Z�ɝ��$!"3C��Y�;���KH�tV7���	�E��+UI�TǱ9*-�ﶴ�8�U��!�=��:�n��1�J;�&nBʵՃZ���Ka�$�=����	����v\��V�yMŶ6��F[�e
�W�g)�V�:�m��Y ��+K���.8v��U�yv��,\Ͷ���ST����J�}w�ǜ�J���Oh���<���̼�s�7Y2[Ӻ�^����JAU�t,嶃� ]V���T�N(�75���%���1iD>��l.��s�/{n yR��������4��6�c��Zuհ�Lo/[���u�LM]/T� ��Ɩ���4�<\`O����h����6�V�+u|��1s)A�@��عg^,F��`<}<�l�z��j�αF���+!g&o&�N�vg��{�M���ѧ��0�!��v��ץ���6�J��������Z�f��Sӂ�+��䋮�_1ۺ�S���=ɽƛG�oI&[�^N4;3�����b�6n礇�!Ǚ�,%�0�g�����]-�7`��ۆ�l11��ੋ+5�,N^�ȼ($�����]���F��81�s���'�.f���d�yq3;�+�W2�%�Y)�˩�Q��;�7-*�╞�\��k7q-��)�8���oQ���E:&�|]Jm�^S�L�ˬ�%���a>4�ۼ�Eb�/u��&�"N�ڮ���p4-�K�qq�f��ؕZڜ4eaY�/��)083]�{:�H9$[������t)�`�I�-��`��q�Ǔ�u>iyW�צ��\���L\ޭ;�6��2WY�;��ؗG��:�_N�l���X�vݒ����juqޣ�d�r�������ո�.��gK}���� �I��B$�O~�9Δ��.����:)���I�e[̋e-��3*��̷��+Ub�v�j�VǪjyu����O��y�+ڻj!��65�e��7��X��.��+Dq[��%i�G�*�c@�Mf֎���sp,Ъr}���,�
H���I^i�e)�/�voEKp����G^gN�7a���W[S��m�v�6v���%'7�o����x_koas^�1�e�, ����2�?��K���;��j��YJ���;�n�b���q�ܧ�����l�S��J�(@�/Њ>�j�=YZL��'�@|�펹m]���ur�:�fm���8z���'V�XC��+K�Y-�F��p�E*O�H7����Hm`W>�����x�����W��Π�^T��j�1��G�q��|-�h��aǗ]�=1Ny|LȺ��}�G����7凥g�G��+ѽW!��T�hɏ7��:F�l�fVY���<PL��x	��Kq.�m���r�EjI_|:�&b�f��ZX��YYX���ɨ�;ui�hgVR����UaAqrN���1��q����9V�b^F�֬O�H��ه��:�0v�a�ٻjcH7x�q_.��W+b���"��a���y��5�8U�C���EFbM��֚�v�s��^:ڊ�8��9��5.^9���P����:�iZ'NA����_^�VT,Sve��,�*%9�ڊ�ml��*�֠�^55��t4�ڭј焔P^�����Y��}7vP��9�%�O7Y�"�Wn$B��Q�Z~�{���^H��\	]MC��QμY�22� ޗ�^���Z�����0�W<TjKE=�.�Iu�}Wdz�q;�>KZ׬e|�F�l����h9Y�s��4�5�1Ԟ�S��x��i���&��ׅNR�%��m�G��Y$ٽv3I�>�T�N���pdJ�
�ee���$�&�q8\����8�Lи(N��X]�Ho�,�e���`nUһЊ���x�EY[�ۚ�Q�We��-�d�sp����{��oQr��=�xY����!h�J�GZB�i!@q�u;c��
�y�/���բ�]ad
NpU��[B7���*�w1��󛵴B=R�uLbA�V��5��_/�r&��!������/8�<�s���d��ݠ�Q]7QΜ�x�G�Wv��c�-��Y؍�;�l�MBJM���ksVc|J��8;1.�B1���>L��m9�_إm@PP^�G��%�}ƘT7�WwM,+̪|)VJ�#�FDf��wY�̀�dg���C�r���v@�����.��#���뼵390b�H`Ӂ�=բ��=�#�U1����۔ke=�775��\�5��vI�y���m��B�F�R�G8P���U��6�>���O�5w]P���!��5b�畯5Po��bǑ�v.>4c�-�Q鹞�%M	���}���A���{�:1,WD��ū�Rr��ɔ���K+w��!'�������1��ˮ��W
��j��*r ��Qӻ�h��m�ҳ,un,8�8�	[�7IՃ�mk�ۢ�ֶ��gi���u�Hu5��?vۙy����-V�2���y�xB�u ���{c��m�Ư/�T��͂�I�Fw:�]��r���F��j6-��
��Qq��*�޾/i�3W2�*���f���(:�f���Z��j�2��j	dS������1���Wn�1ke^&0v5�+� t���	BSJG���ۺp��$�h&���j�e��9k����A��Z��&��Z�� ��9�'��h��\Tִ���-q��*�45����Х���\�X�l���z�|�]��֥;N9B���i��dm�*	��[�j>��Qbz��؄z���Y�RK6VgXW�e���]xw�ieeq�loa�Ol�HǗniO�������}7�]�f��{���u����B�#*�� e��:��n-�N�U�ؙ�P���J�kyT��mK����e�v���Ѱ�4�f��U�9��V ە��`H�e+�� �*
c����ۂ��s��o��w��S|�t_q��|��RD�TF;� |vVU�v
]��`Y;��{�s���2b��u
�]P4V|��p�� ���7���/VK�,�z��rVneQkR��+U_U�Y��D�C������G0�y3i��CŏQj �v�g�r��:r��Q��U�@G��;�;�l)j��2�-�Y��8;pYkޅ��3zۘV�j��Г
�%��[�[w���]]�ƣ������e`S6Ȅ$}~+�:�Ņ8��*c�`[�rӓ-U��K�{�&!}��>���wa�7�}���ö���4���jt�5�G�UhƱa��b�=���n��[96�$H�����f�l��wh�
WSŴ�Qbv�HiF���M��qyrN#]�e��k�\��R.+k������|�S��T�H_'�g���F������K��N�],Y�K��cx�q�1_E��\S�U�[�eW��*��Xn>�Fo4.B�!��7S��f�-m�������b�<�_dR=�3�&"X�Ҥ�h�)u_.���w�OjP�M<�W_Wi��)�W\��ic��(7�Q2�|�J����J���c��k���r�$:�tr���x�1[�z��7S>m�>Ȼ��Ir��;�cW$�Q���^�5�a�=K��x�^�ת�"aEb����[p̦C�O�,j	+��	�ve�u4�Z	�z�';��º��9Y�ڶ�d˵"�K3it�z1w5�w�j�<�)�)��a���Z����葋�2� /'^<��>2�۩�k���w��A�A�M��GK�++��ӈ�x�U؁����Ԕ�ǭ�t�_ƯZr�w0���ي�ZV��P���(um���N�%�'q@.�u�,���]3j���W]qg[�Ӫ^��7J�[� 4��T��p�x��
�<����$̰�Áh�j ��1�e��\5�}��,�e���=��
2�Z܏�;�Q�{oI4̹�_Uъ0;Y�[���5cK�6�`��1�&��CCz-���<ޞ.���W3P-�o�� ��r��G�\4>Yƍ�v�����4E7�V�bݻ���\x�U�59��|�b�[�u��ɺ�\%wp�����s1��ʎ�jo�^����
4�ə����\�3�M]� U�;�����8pM����Fu���uu����KO�U������ڍV�\9��m��1n��pkw���%Í�-�C�f]bmHs_�]��>w-;�#���r���m��=����mj��@���6x��e��oU������#�`�J��:���!�+C�i��Vb��͚��d�wop��V��ՠ�w5M���W%]�t�w��f�����yɸ�]J㇠6�;��v/4,���[�j�3�kc����[��4o^@��Qr00�؛�*��J#Mw4e�Zf��ǻ���ETi0�h��R<���gT���1F3��l��Ǒ�l�H��Y)[��
=y�k¯��"�"�V�I:�&uȩR)�N����n�L����p@�ݛ�V��p<tP�f�_՗�Ჵv���'�T��f��mL����R�0N��Zp[��A������^��&(L�Ty����^�Ѩ��.�3��\�g@+խtB�����e����+�k��	�j�kX��Iq�;�zL<v��u���)_V���U0"��5��s1P};F���˺p����ٮ�t�yG{�v݋��KvS�%LQ��N�..:(-� �&��7z��5|��)s�q�Y%�_ �H�˸�
и�+���=F�hj��5l��M��D?�#aus$�l�AC^�ϰ8��5�A�w�҄E^�ȬATsҀD6n��{J���=�y�J| E�f�RK��Z��Ms��^��zL�	7��_PY��w��7�����V�A�R�{�ͪ��m�쒳���.=�nw+g9-��o(ɝX۵����4��s��8�r���G4~L��Z�Hb����۶��F�V/7ZT�݅�Qb�a�k����dz��c3�f#n�.��*ydp�ݫ�j�}ȣ�G���p��k���n�B�����++�cCh�	m��*i"�5�86MeW4r5�6�~X���l��RN�[�=�%)����x��:p�Yc\bb��rN(D�B�BR�mq��R��u��I�N۴&����6�1��'=Zڇ�Wc��-�n�o���84)�9:UovƚF��vQv�s)F��r,���;}�%浧-��Ru�2���̱H�p�}K��Т^d.������GY7{�;���/���{\�5XvC�+����=�C������C��%Yuj���g
�^�݌	;#ѳb�bAU����l�MK��JP���[{c�I��ԧMu�9wXB�� v��ɝWg���ΡQ��e+��l��w�l����j\e�3O�Z}յz�&�5�`[s ����CV~b����J!�ݻo���a�Ϩ�]'\�<�� �S&�	����^�`�
�>�4m[y�a������W'�wEj�ɠ��W 7J�S]�Si�y$����s5@�w9gTy�Ʒ�<�;.��)�˽B&�K�����&��	�V�.�72�PQ�k����<Y�26���}�2��6��kP"�d�O)l4�(��X��P������RN&%I����uh�2'AԳX9��:�ϣ���J��>��������EȬE򈞵ux/5�]z���%t�ᥥ;����wSV����in�r��@�3��7U�w�cXe������27U����T	S�~�i�i����r/�R;�l�\I�����X�\Δ0�P����lA<��|��ƽ�"���C7�m��UYF欱ר���"g;r� ��ųέTy٦[h��u{]�oK�
wq������G�3/���3]������X ��c��U"�v����b��j�Յ�.�`� .��m]ؘWqS|M�"��^�e^a�e��N���R�H�!�4J�a����,�E��Jgp�OX�ފ�-��goM�Æ��v�l�뀭#''�E��^�n��b��ջ�S��&^�͔_;Ӕ�K5]脼U5��aoF�]�{wٛƺ�t���jQ-��S�b��]��Z��tp�.���n՝�o�S�8�nd�I��Sq�&�-d��Jn��o#�2��u�]��]2b�հ�Y!���ͬ�Tq����M�]qO4M���PiN<���/)�I쮹���j8�~��	�U���������T�M�8�l�x0D�#�j���\J�ӧɣ3@u�*������*gIُ!����LR��~���h"�}��z�b�4�q"ɂ��=ӻEG�3_oP::�Ҳ�X�mI��E�F���aQ�5��&���b�rtQ��  �#�`�Ԙ�r��VZ��}�8a��pqL4-�Bjc���X޺Z��Z����o"�;�+�E2Vw
wρ��h�{.���@��.��]��ʷ)��s)2�sGo��WC4˘�*H����;��^�mG�ܵU�� -����f�k�G�$==D�a��J�k�֜���^�!�2R�Ϲ��P��fM�w�/���MK�D�a� ��4���G�^D�}Y߹ǩ��M4�i�#;J��@����a���LǥX��X.���p�b�a����:Uo\G"�ŧZg
�w��8�!:�yM�t��#Ґ��(��X&� *L1(ͤr�-��of�V4�[��N�<���p(�^�<]��ݳ�d�5ZƄ�!]�.��\e���HVa�����.\8 �Fq�)�/T���U������n��Kw4;P��+�\�,�ܓ�)�y8��\ZLs,V�����+,�˄�ev8����	cAԮ�[�v�U�h�n�r\k+��őA\�l�xqk��ev������Q���V�ʁ;1a�2��m�n��+��uu�F��YyCu����ա����-[���Ec�����P���m���/�z�Xl��6;���_Vf9
<���mԑ�����z)c�^�P��U��X�37�d�)�y��R`�	HM��!l�w�xYF�=����$�]gBJ��NR{W�����%�[8�>3�q9zq�x�<����l�#���zl{]{���k%�]a��;)}1-,�A�Ԃ����Ͷ��v[�L�h?���8�����ݡ�e%>4��Z�n&v;�M���ְ�	��/,�V��d�kN-C%��q#J8�r�!��,�ާ�GQ�Z��X;c�׭���X�F�v�I���oU�-ge-5F:�N�!JufQ�owݵDvL��gqNk[��a����α��9��)�^��ɐ=R�R1vy��M:�{Oٻ��r�!���x�����p�Hm��n��y��]F4�s3+#y���yw)�9}�zj��lf�g
̫�)[z���2��Ej3�s��lgi�
m�<J�}����/gs�3�"^�F	� 5�GZMKuT1V��-^f�<�VKX5$5�$���D��d���UL��d3WWi#������d�"���������M�R]G{�}���5x��VS��4�p:�N��@m���VI��o�TVٺ-_ikZ�ku���:Cnz�ǫX���	!xk��ҋ�b��Xr���x��[s��[��2�:�2۲-Q�9�����2�����u�"�Q�.lPn̕�+>�Y�����{������X��2���W�\
���,�kB�]�\��}U��W�=�1�ξ�RՑ��;'�}��L�f.�l����Q]q���� s�!��#�gkc��3�4���$�x>r��.<>N��2�Z��XXE�3Kx�-��>K��Jl˳E������a�dL���LV��=�U���VoKJ(����8��Y5u�p�5�(!��JX.2V�v��K)�Uo�;:�5X�,�w������BYF�%�*�ہ_�������U�������h��4����S&/�a���r&��vD��7Jyֻ�^Y��n��Q�J��\��V��;�G˲s����uΡq��x��<sgp�%'C����\�B,i��#�f쵕4�9�V����[m6]p�;�uDm_���Ʊ���R�(e�2y��X�۫�[��Z.���Ώ6�c��b��k�]�P��+VGѥ��9A��Yh\��z�C"�E"�}Q/�(�O�� !#+@��^��r���6�k����-Zvd�SP����r�,�&�Y�`��!��[W�o/t���{e�e)9���(�шӹǤU��-��	|0*�:	���tkH��֩�2�r��9+�C����|tGz`�y��ȩ���+��V�Bm�dJ���w+{̵��7"E�헐U�խ�@�2l�+B�/('��=����g��=[W�9��E��{,�["u}z)<��3��&�d��K��97����L����B��b�dDU����mł��UR�0F0E�	+)X�AEE�R�i`�-���b*�)��
����"[�0EF1X��ڱ�������DdX��,X�-�PE
�(�Tc��,DE�)mPTb�b�TE�����E���TX�A�X�*�1h�QH��*�QIdQE
"�DTAU%j�*�EDETcE���
�cT���¨�c��-l��E���lU"�����kkQX"�TUEb*"1`ň��m�,Q`���QR������Ԣ� ��D��EPF
�m��b�Z*�Zث�U��TQD�D�,g���[Uյ�:.��2�U�c5���*�*y]�]��=C��X8l���tWFC�O���;q�9L%�}�N���'hɼ�L����E��Ƕ�iI0��QU��^ڸ�����Z�_=Y�bX/�d2��v�U���Z��Vhϋ���3@��nR(�xm�۝{[x��Du�<d�bv�c����Ұ�|�c"6K�v2���/
>�]���8��f��*g�JV�N,��q�}P�Z�#S���ӵA�1H�w�"�n�ozl�S ��P��(BM��y���u�\,]��������F,���������leGL�{_.WP(T��l��	�v�}��:��̣��ѽ[h��߄����Z��U������ W:���N��Gp�1^
��a=ˡ����)������e��yD<(j�qDaNf�hS:]E�>J���Q�+ �Ӆ����&tM��<�9c���$W�u	4��S�y6hm�2F�l���3 4N�vg٪�F6��7���v�U9>~��Ȱ3$ef�Ғ�QF�{�r���P49���l)�r��j�\�Ȋ3�N�^J�:��nu�{�Z?��uI]�K�\���[3:>�W�sJ6y�]|o���V@��^�ّ���:a��RՉa�p�w�������x��OeB�Q���@�T:��Dn���t:tK?
�T��e&��ӻz�j�ઈ�2Ϭ�Jâ�d��7[�9�N�@[�8mX'�T���>⥸̓c4�Y��ԝ�V���3�*����7ۗC��g�n~=�-�%�f��f��O=~x8����5��{k0:'(�5ິ���CH|��
����#�we�L����w��_��3�07#�Mw��6�X��"Í=�.���Ѝ�m�ܛ�n�� �w ��Q
$�x�������ج��7F'aF�;�;{)��[k.c1Qfv		�O�_`��	�3a��K��ȵ�	��Q�M%��o��	z���|9����!\$�Lg�tΌV(-ϸ=2�feԢ��ZQ��Dv�>�#�/�mv E0B��|.��!�D�4&eyj�9�L�����/�f
�]��94C���Gm�J2C�}�3M)�PT4	�4z�TQm��]|x����O#�u�)3�Ѿ��9[v#b�x�IgL���f�ID�,o-�%��B<5\X�	{Xk�#���ѫ��IM�t+o����5o:�p� c�s4H��1�� u�\�g�/_��At���q9k7U�6̨���F=���_,)�\��e�C�g�z5���eK�X�c�̼G./<���[}���N��D�k�u�|��Br`�@�f�����W��6��E��v*�u��	0������ >���d>�N�M��������\a�ռ��!�}�����¬�wc��y7��*$W�OlhmX��<F�U�C��o�m���ؒ_%�ʀ���\��'����s�{�Ş{�`�m*�c"H�1����W��4B���F�J��Ǌ-��t����\�ݺ���`=@|݈�a�߁c�>��<.��#�e	�eߨF�쌗Вg�ge|wj��Q����.t�1-+&��924��
��o��_�Ta�����,�<����}2^ŷ,�9�i��Wӫƌ����$8��R�-Ȯ7(R��5^�2��Vi,���6��=4Ȱ�\b���(ZU�7��Vn��9\�/ӭ�X�q�sݽ�0S華�/Z؟��C%�E��s�
UtL�Gn����x����{��;�9v�i�CH�G��5X����N���vdA)	�ᖇ���f㧣�<8$G��n�=�z��J����*ǻI��{���H���1MSj��>w�)�Ζ�V�l�T����9�����r�{�kJ�ˆev����IÄl�޼l�����+�@�����Q�gB�|A~�"�<�=$���=v�g�s��������+����ب�F��ݞ>� �6�g�9[W��N�\�3�׏$�|�{�&<�_�I�ҡJ�4��愻T�ҮM�B��7��sZd��U�bs�Z+l�CN�!~�+��L=-��VؖR���AEҐa�ϙUY�r.f\�ˮ��0��]���p��T���j�\������C�������qۻ�Ԙ�I���X��%�P/EŃ}�Â\������dM:۲9��P:�a�;���I��u���y-�B��B�e�@[S�T9SP�3�D*�wl�73oo�y��DjXeu@~8*Mꤛ�J�R�jjD�����5�_w[+��^�rqy�bG�v�p�UrW榔�q0���r��uWB/w�JP��/bw��K��1�U���N �r�5�،�^��xO��/�h[����F��"��o7r��{8GX�ټR�S��%�D׵�۳C���߼݈bެ��Hz�r܈F+s��Ne]Y~/�q�5J�RvR��M���{^��F�����^z�� *�W�n�A[�����Uv9}�+I��ZFbц��ajkh��{ٗ�E^�W"����kgq�b�JTZ��*1��o,���;D3��Υ�Ȧ�]�7��{l�g���(Q��@�bb���iD۔A��Y�6@��iglez_Vw�mɛ ���Ď��7��f2��u�S#
JC�85�y��p��[W��j�Sራ�~���#�
p���T՚���W�mٔ�����>u�O�r]U�� ���V:���׉n��){��^����9�Ƒf�ZC��5J���d�]�^Д�y:1�y�LgtF���%L���Y���v��-�a-"R��D�J�O�UO��ײ���������B�u��K�1�7���)E��=#h<S��3I��f��J��[?9�8�0����t1}l�>�p���!m+
���Z6NU�I#_eyV�=6��/w��N�x�QsZ.��*O}��S����Ϲ��`�&E�v8����{�v��݉��b �CE&���8�*26�2..�`Q��n7CDV�W[��vO+v�;-.%]�,u,�R�\�r ���n�q�P�c�Ý��h�I��6�.b)L�~W��4.���qp��Ak%��%�)�T�A����4w�.n��W��ܬ��A��^1y$o����xFf!}�)��-�G-�7���5>-��λj��rR)q�2�ut��Q�x{!�/`���!��f%Ӡ��6s��U
[�kagN[�~s�l�d_�����5�}�
�|��Û�Jj7B��F���w�~�臎(j�(�4�V8�)�.��%@�zD)��y���C����ܔ�&�r�/ڝIu	)Bq�r���١��H�y͗Q���f
�sUc_9θ'Kaj�\��̑���J�%N���DP�����\l�<�ۧ�ܱU0��L܇�g�t]E�<�t��p+ۭ��"��󁳸Q������qH���7�4��<7��zTJYXC�VbR��܉r���V\u�~��iH��������X�}�'z����j�s_�׶�҉�pƏ,#k�4��b�o2��1�0����쑵��ѝ�mX��R�gyV�������Zl.���y`�_<�ܔ�%�����;џ/<>�b�ދ�����`��F�I��mߨ��.��d����'�c����ow�f�ܬ�{�\)lL��⯥�1<��fۦ��DYJ7�ӖD�t��{�8��v���b��%t}���v�N.���9î� ����|���o2��Hm��e���nR$��Ն�Q-+v`r��RV)��޿f`��t�r��km��Z��1��_>�znMK�nm����_�4��|7{�X���O0�V����j:v�8�4ؙ��%��U��Ks���-Fd2����y��m"*O�z�����c���,�Ӥq��$�����-Pf�Uq}������gSdv�z����+^�̳�5�T��V�E����������!CA-e�tX���:݂��t"�O�ܹ�T��ޫ�~~�q��;�A�&��M(���v�HR 	H4k�����:���wϲtY=Pŭ�"�:J1���s��b�:�-FaEyA)P2H�1�����63��9����H~�ӝ�4ȸ�P�v�f�s8�ۺa9�p09�BNZ����K�F��Y�dv�a��o�o��A%N!�$hȺf�o%om8��� �;v�E�Bj�[^�D'b,���l�RSU�q5�EP�em98�[�s�`�'�A>}�r��ӑ@����G�
�ڮ���w(p����}zuε�|L��]�Ĳ��VyP������
��|�-b��[��k�%�~�n����ʵ�:2*S+k�c��
0�ݒ��B�*��i�vj��mӜ�L�s^lʋ�d4CB�;��;F��]W99A��[Re]%�	�1���Y�;�߳]��T�)&��YTI��\1�Ky3��ga�r9Cr����򾆶��T����	��}t�2Vń���uĹ@N(ɘ6�,�HqvV�63������N�d:-b�}u��������O��Y74EJ��x�����.�^m㩥���=���K�\F�W����?�MT8����F	UMF8f��m�'y�Y�S�Ϸ�̪Xk|G�����`���)US�K��E^΢��	HM�����0�+= ��u]��e��E�,������/=@���|���Uڼ-0GVuQf��:���w+�aMM���oi:�7��=/�&n^��CRw*�L�9�0Z�o�Uɵ���-�r�n9N�,0�^S<�s��X�P1_s~>=-���ZS��b��S&�A��U��]|�v�ߟ�oA>.�p��׮K�����%�-��H��b�v��d�M"/�&KS:�f�Է�5�L�+|�?M�����;�p�"��NFpȖ��"�1=Ar�ͼ��2w��K�*.�!�D�� L<p@���}5��Ϊ}~Uv�Q����7��*��2��;�|��>_#Ы�����O�}�{�'&���cr<�>�r����,y|G�Z!�l�[CR�ϖ�9ʠ��V�wG/pۧ}��W;Tn��+��o�,��}|C7y�l��lP�%�`w+V���c�o),���Gާ�����tm�I� h��=J��3�~~�Bx(�h�Q�"��S6׶m/>�cegV%�"G��c��Y�L��Չ���F�%��\*�q��=�G���Ju���׼oB��U8	��r�5���a6C�?��|��b���X���}-�֫{uvޕ�먲�d�5�8B���͌R�S<�0D��D־�ذ|�����*�)c@����3�ay����g���ѢP�Nez]ޭ�+��S�.y��ط�]��
I��n��2ɯP��
B��<*.P�[�*���T4�	Hz�\IaaC��ѵ45��}m�B�G��I��rNHg̅�Ux��H�&M;懾	��L^�X�0V.䓚�����r\��^�ק=��N�S�K+H���ƍ
P��6��~z6�"�R�竺�H�K���.B4%L���Y�nv�8\�� GJ*��"��9��`�[����J��M�����]5�~���C<�'a��K�:��w��|����A_U���z��=��{���Ⱥ�b�H�J�:���|�%��C����A��y��R3-��-���9Y��Lg��ʵVZ�"���kK�1Q�<�ʔOM��y\tq=��nZ��tMFq��v��SC*9ݤu��eiܩ�U>�qـ�-lU�n������ǐ�ӽuDq�5)Ҍ�^���>�pΝ!�c��f%�4ߥ��WZ;9�׵��<d��lAjqh���x\���-NXs�[/�.PD��n���{Z� o��g:�eOFa�G�h�݅CE /�=gn�3��|�/��i[�B�O�1ӯ^���Z/�~f�N��u|�_"��@�-� �=�P�o|���f�*��x��D�e�3�᳭ە<�'��d
�\���D��y`N��/6F]hKh�n�ky�K�x"D��݊`r�� ܾ�x↨fH��:�q�N1�B������Lp�y;���/��Se⾺Æ��Tk�\�"7B��%NH�r��١� �'9�P��=b�1%r�/y��@�,�"cw'�%�ȿfH��XWy*wo���!�`���7�⣴󴨗��wGY:X��N��h=� �q%\3���2E\
��w��D�@�����ˠx����1���E�fnI��^�%,�!�Y�(�KK���>V7=a� vV�}�ơ���Y�� M�л��]����;�����y���e�eȾ�h]��[��B�6lˤ�s1��5���tF�^�����\k[��hg�}wC@{���I��Z%�c�|z�Tbi��vSV�����)��F[ԐSȘ��௘��z^ļJ�ڵ��z%�5d��m^��Q�\�qsu4��,����Y�,����m�;@ţ��f�= (�Nx���%�	���U�Y��xї�J+[{]�%G7=�"s'���w��R�X�>�s=�/Ͻ��Ie�U��+;��Oe�����vs=�6��B��3 �7��1;��r�ׯ�(tR�Bd�%d/6U�M�}M#�B��2:�q!2LXq���p�{]��ܡ����[Q�T���/�����˾ST��P���� ���:�8�C	���E�F��<(��ei�!J;[�؜���f�׎�r��Ƙ�Q��2�\g���҃���JN<���՗*Jm��7�)R����
�]�qf^N�����Y�����@M[�J��y�Y�1ٛH�&�;ٗ�q�7�|�Mz�F&��hK:��7Y�P�z�&g]��Vuӎ���y�X]�`�3�n�t�yReY�R�-������� Z�*�!�\N`G��4��f=��9C����w׎
U.�<�P+�q�Ǩ�S����npB�7/�6�Ku����7��/�/v��ZU��QXH'�v�Sl��E����Ы�ԋ���Qs����u6�{}�_�J�2������Y�4��&��.��;��{v�����Ǎ:x��^�ه�E��\F#R�erus6�b����H��N��	�����aT�uq'��̸wn�Q�#�š�8U�K�|�h���._T�ڜ݊#��7r��l�gsx\���vd=�)v�¢�0u-q��u�(�*t8]��{��m��n��r^��Q���Y�2��n�݄5r�q	�w�V���rJ�R�}niJ�����B�WJ=Ϫ�u�v���4ҭOu�m�p��x��F��]��:����">+���m�]Wy�I�mɤq(�.u�9��Nq8a�/���sz²;�չZt"ʖ<�>�@*deb��u��#V��AL�U+n�^9Z���p0�;��F\��m����1�%`�Ϯ��
5�@л�h�K��X�E�g:���8�;�D,���[s��%��P�ա�vh׼xܠ��\1�*�k�D���J��!����l�ѷ��Y-7R��`�N�mB�.Xu�{ԧ]Ɩ�^����v���B%*�QG�va��
�]*�v����2���4�h��Ct3�.��^���5xc$*5{{]�����V�������n�pF��λ{��P��c8�Ydk����R�P[ȟ �������
��"�)wb底�[Y��YYji7��oz�ap��a��0v���"���rd��y�xŎ�P(�UQQPVEb*T�DQ�QHȊDTPUEX�QTDEA*�`�*��2,X������"",��AUPDH�,UEQAYQED#V�� ���F��1Z�EDDATDX"�F*����*#1D������Ub�dTF$UQEDV1���-�(�UUQ1QP`�(),Db
�$Q��%�ETQAQ�,�b�UU��aPUPc�b�,TTR*��ȵ�U��D���-����AX� F������%kX��UTQ���R�"DQP(�FDb�kb!Z�TX֨�*�"�VDER�
*�
�5��R
��PF*$U���3��G!{����U����,��)!��SPӽ���:�J^�*��6�b;�43���8=���G����M�[���,q��Y�ο���[[�J���f�P���ϖ
j*���;�"�Dj#�8iy�} ��PLz\�F�S��oUe��9ͩ:0�A�h{��?d۩���gy�uIO�]��b��/�4�y�QQ�d����ꚯ,Kuc�4�ޒOD|0�|U5b��Ͼ(���U�_���9C]�"RS#��kW�^�J�WM���[U�=�6ICʳ(�^T����>�:2+���L5��Q�m�bi�p1x��k��Y,���:t�n(���AQ�:�ʭ%᾿�O��~@Ҙ�I��n#hn��K(�j���=Jx�'=��i�<�JT4	�5��mxZ�8��B�Ff0�_���R3��A�m���s�7[����q��Zs���B hJA��ۥe�
�ԝ��b
V���=�:S!�:�X:���un+n݊�]vE��L(D��7�2�fȹ}�G�nH�P�Zu�N��Cy�+�C6�qE���Nk\ =�]�MQ�4��5%�5ך�4;����{8��,��/We��k}�+�[��rV��泃�5R�5�.�)ܦ � x��휅��`��G�:�^��rg���̐b�w���T��9=5�$�L�����P�m��y�*�s�j�2�L����<(g��5v����П;���fD{ad�!nM{ "���rh��$�J�C� gb��)�o4��r�$o��ٷ�,T��eſm]β~�*-l��d��.�KZ�ő��������+� �竞�=�@|��D|��h��\p�.9���#�	j
��%��z�h��t�ʞ�	W{@�¼
����*�?��aA�ѵa�O����x��ڗ{M��g�=���!�L��a)`���L��P%9�%X�2j 3�_J�講�M��:�|�]&1C�Rʈ���.��X'��8��~�b��y�c�����j�N�����acy��L�E�:B��5�%8��D�*E�|�b���<�<���/DwUV���U����Ɣ�0�:f�x�|P���,S�y�V;�RrT�׮r���Rabso����i��=� �q��L�t���Щ�G���z��=Șõw~�Kv0@�d�G�7A��5~evOP5'r�J�4��愿�S>�;G���\�ʶk�H�\9X����������e���g$�R*T��Y3�l����f�6����.���V`�%vs�l`F��n׆P�O������Ɇ��;ɡ(e�e�^���{�DJ���w���N}��Ր#�tY��j��"Q��c��*�*p��.+��n�a�e���r
��XXZ�"��Θ�]�:�s �	�o'���'��\���굯n�MC���4�c�,T��ԚDEL���w��s���[ʃ�
�+�{��;O;�n�Q�bܳ�t4��Dдj�<��8����\eg�n����$�� L<`"b�_Mu�3�T�w5��و��/|�m���z��`�I�5�RCKu���Խ���a�y�i��q^���v��K�?:�HhCGǫ��xT���5���*�&�~5^S�t��N�雏ϣLeGL�����',�C�4(���5μ��=�Yz�ia燎�${��D�B;/�?{rF�t����ٱ�X*a��ڠ5�m�#�:�	��Lw�ǰ�t�{G|;~ʾȭ[g���y��)|��/�8��r�0�5ڰ�,�}��mj�4,�C���x>�7qd26zl�d�t�J1�#
�R����͓s��k�)�x�%m{�K�[56�w:��ۻ���DR�lT����Y�%+�"j����ݤ.{���E��^����Cp���)*ް�oi��P��W�8unB�M���씎R@;��za��%N᧸�L5�z�w#��' �$y�X�O�|�^��8`Au�xs�P'!�DWU���䍌L��K�y���ؙ��-�6YR�zN�1=U�xy�7�o�N��N�S��ZG���;\h��WQ�YûlAuꮞ�ϓ��b��hx�Cg[�D!(�����,n��j���EX3<B��u.������zP"�����Q�3�����Ĺ��͌�(�%�}`1����V��'JOCr����#K�	)�Z1;gL8g�|��Ұ�#H�p,�|6��hۼ����B͓��t� �;��/.�)���rg��,9ӭ����^3:�NؿQ�6x9[��v�D��.ԄC�ӵzPd�����o���=��̪����DN���8�ґ��h�wP�u|�X�A����v�8��UγPݡ~�K�>[��ؠ��82��T�s9��g��v�_���8��B�)�Jj ���L��������C���;��5dk$�3ob��T���C�Ս�ܬ�7:�9D���Q�D���#�b�����.{r2�$��u`_^5 �r��2V�oX7��CU�-�=7���+9-@�B�#=`���F7}H�8�r�>�Ֆ�����N���_m��Y�8Wh�*<iۜI��ήM��j�(H�lѻ��\�4%L��TXHeJ�۱ʻp���TTƛ9�n/yԑK����8�� XM�~s$a'��ُ�~�6���U��T00�c�'�.^E��Y���J���9�ܰz�LU8qN�z���
�c3n6��@j��(/��c3�zτ�:-�j�"�[�*�m�US���3�	�p�͢B�������M���5�rR�XC���AD8�"Z^��a�����m�.��z��3�C+#�=U�������?	�?�G��v_�譙�	�lv�ギ�U��NJ!�6��=�KM�z"�!�=`֭��zh3eL3���af�9ͩa���onbj�:o�(S�\��m���&_}u���@F��\t�ϒ����Rr6�nƗ��'":��\e�-P�����m���Iv}�`�|/�\ˁ�GVD���V{�$��t�\�H��C�S�����;����5(��{P���gI(j�������O��:1W�7>�=2�a��l�!�)n�BJ��e������!��ETt4	�&8&e��WGڣM��r2Ȩk��1��Yvh��O6�`)�����F���+�x�� ��Y�mu�)�EF���žw�z}�R�1ފ�y�
x߲����,K�QE��/��)�vS �x�<��Դ�n��I���ѩ`K{�'N��:���Y?���q���'բ����t���Pr�0���}�9�iC𐡀�M�VT��_	ٮ�Қ�[o�`�"��l\u�R�q���d+R$��zfv!߃�I�@o�S>�a�;q�<��R`�S�<����`.�`�"jϧS���=)���N6 <i�x7�3g�3f6�>ǝ�'%��"�Duł�,႗'h�$q�gXnݎ�͍*��{WG�e��Ʀ�!�֋o�T��{�&�[�YY�rU�H�kͺ�]�u,��M��R^�/9(٦�6U��߹��3�΁�i��H�2��&X���Zu�P{�מ+��-�Y�P�&��Ms�O�_�o��Es��me����^A�EʍM�$3�n��Uf�k��vE�N�s�Lk} g�J��|�
�0�X�k�U�|�v:s��ѱ:yԋ#{!�fU�{�%�X�,��fn�S�2V�qs�l�>ŔQy��{h!fYs�:3����ķ�@z�lM�W�,��Y�\BE]o]3�L��+켡���M
�+�X���!H6�|�MO9�N��Φ�]n'�&��P�v7:��t�����L�s�mwڎ��
���^�ۊ�%�����t��-�$z�<{�̜}8���:�>w�S5�3��}����ӛ�����lZ�\Ey�P<1��;��ϯ�h�Tu{|��^�[�շF9M�o�;�����W(Q2�+������b�.@{eY|��� e���	��t�MՄ���&r�;S��|w���]ːH�x��^����Z��N���kͪ�w%ʍ��͖3GQ5����������.�㞊JZ� �A�/�w�<2��'f��z�@��`TR���.���S�}0�e�t
�Ҡ�j����:c�R1�w)��Q2ޮ�kLA,D���Ez�W)�J��E(g���=�!�]b�'��ёf�%M{�y��wNw�v+Ղ	�Q:H-A��{���c�;�X�t�9ө�ªmTO^�	}M.q�mq*������L�A�0I�R�s���v�����B����1��l���K�{�{T&AӍU3�gS��B3�@�\]*3P�N��u��7���L�\,�]:*`[��ȯ6�6g�>d��¸��J�J:�k��<ws�[�Ρ&���Q����ˊ�r6{s=�N���s�2*Շ>�"��2�!�U�U�lu
S"O��5Ӆ�m&f�/C�m>�eB���wL�xy`np�`�u2k-�jf�G@���n�֋;{����8WoM��5�nT���R�Va�O#�{�y�<{��BD��]�DV'�w]�Z��A�ܲMh��s�hs�9��3���ͭ�<y֡���͌c��x5[�������+��'"�)`��O5D׵�F�hd����u�i��wL-�Q���-�����0�8��(�{r���{�,c�q&�)��r��]�٩�ݯV��/.��k�4���G��H�\F���*crM-su�R�ͱ�(�g�����Vr���s`cy�N�':7��h�Y�8�L����#�YWY!���}�Bk�0�;U�!���j������O��]�Bآ b���1�l����g�M�vP+Զ�+�R{g�%UlBT���mg��ڌ�s�:B7����Ƈ�,�ŝN{��X����tVLҋ�
��C<�'a��K�#�u�0'WEe`I�¦s��΍MM������M!Z5��9ՠ�}0�~��3�Ұ�U.ݥ3�S�6N��%��KR��Q$k䴚sP�]T������>�-NXs��e�-�}oL�#R59���5��tw���e��5�k��`}-M�u|߈Tg�W��@|<�4�s*#3I�nͭ��z��#}2�=ݫk"������5]1�=ͪ�(��� AgCהv��7ݝGw�쭑ܨL(����Y��|=�{�훸͸v���j>��L����v����"�(�$ϡ�Q1�t�76z���[7o�K�oM���^�瓨;A�hٝ�FӟC��
T=�JA�`3��z)�Z�3ë32��Y;�L,��u�v�c�Άpt�ݻ�n��n	T��4�;�z�-���Ν��𺚦�C6�P���{��gÕ��Õ����V8�)�%�S:9���ܪYs�y��#�����Z��kO�*r��tDn����o��lk1�W�J�|�T��8�7+����:l��ܟ\�yd����|^7N���Dܱ!}7y�s#�ɨ��h.����� ����2,� ��b�d3��V��U��#/Y���g{��$B>�D?[�8��hh�ѫ.!P1�u c2(�W����f��M,\]%y�pMC���犯F7��o�'�������^'������4�/�O5)�A�g�/4�}��vX�Ug�T3�1:�׊��x�6�#f.Y�-�hc�MglR�bˋ���vfQ��݃�P���mrf�\o���N�U����������  �����1Զ��-h��� �r�9\炲��*�s���,٘� ��n�]*�p���φ=���M)�A���L֝EFK�<�+����t��ē�8*F��R�]NR~@sW�@��$��%�o�gݍ.V����n{�X�eĩ؝�댃����
�Қ�:#�k�����C+�$��n��/^)yB(�+��]�۲�Ǝ�?cX���+W�����G�I�̾��$������>��е2�������sT[�(r���L8t���(��]�4Z�
K�Ii��Uub�;�V�:���{t��釲,�W�����p�z!{���M�^�x�� ��/{ޑ��]p�D�Ƈ��b�Z��S�;����ȓ�ƚQi�؇nI$ �s��z��%Ʋn�.a �9��Q���t��n��d,��s��v)�Uv��K�����\9�z���^$��`D�"�6�0�-j�iFXs��8�\E�������Y�[�V�"T�9�^�0uh�F��H��h��4l�ײ.����R9ę�t�1��|loEkFm��ʽ���@�F�'��y<��s!�� ���
���i���� ��`�42����@忖3w2�֥��_�T��]z5b� 6�R]*\w���m���+��.�;s���e�3���)u��]܁��t),���d�Pm�sbJ]=;�oA�����u�']2Z�+�&v�U��r�,�8�욳O>ܑ�����O��[��F�N�hIy+���q��<w��o�m�|y�c�t�R�m��Z��F�Y�:�Vxf���TBzK���F���ЈH��I�l>
荈��� �s+7B�8�i��P��ۂtZ�e�AP�c�W�i����$oXU��u:��N\�ͬ֬�q�s���șL��3�<c*)pJ�DR��X(�d݅�+�c�D�"���)f(�g>�gh�V���B�2���˸�H��F��<W��� ލ_=���Չ����]n�Ap�,�&-W��F�)��1m�yv��f��1U��z��k�E��J�J^���(��%.�Z�y�T78��"�5�ۖ;4&����A��^]�z��A�3�ex�쬃�w�Jbc㏶i�7�Ƿ���L����N���K߅]���m.���N5��<��K����Ow�(;:�9��e0�ָe[�(<WN�흊Wu�ݙҒ{�` ��yQon���2�	qm���V�1*�M>�،udfnN����1�4���J_\
c�/�q'8�X�i�y��bF�]Xx�9������Μ���|D�K�.PV���;�J8F�ui�T饙uc^!J��R`ۉJ��:��( p��f�x��qPL����]�88H>H���Oc�z�v��ھ�P0Y��u�SZ�Q��,u��������o����϶�ߎ!�6�vٝ��Zd1��<������t��1�w-�e��$Ff���*ُS��[�ːV�C���moEr	�S�Ϧ������Ū���k�x)X�x���C���_�T��'6<���J�_L�T�I��B��HؓX�2��k��/~�Zb�������v��J�glvKܫ�P5/����|�8>��V}q�̽o,�<:X�p#ǡ6�w[[Y�\�5\�['j�E���A&�+y���p�V�$q�;�RՓi;�����{�ums���t��,pVc��jY�Xd���j�~�c��r��Ǘ+��`רc���Uަ�@.�i]��2���(qF��8Ťi:�Ą��{�U�LwD��,+�7;��a�����q�l��e㘡2�����is]{V�����{]�f�vSyJ�j�Վ��]�W�Q"�n�c�DZ�1���.�Ҳ"2|Nŗ�S�8,��N�M� �N�"f=�gZ���B�o�곦���CNe.����F�mk@�ڸ����g�G���	ڻSDΑ�_�Й������W+��+�3OR�V������E�Gz����l�xcuo�cT��
鼚y�Իy�U��B��ܽ5��@����s�3v{ٔ��'�ys��=������1UX*"Ȋ�F(,�R
*�*Kmj�$QQE�T�"F��b*�V"�U��P
�QTDAdb����PU���EPkI
(�$X��J�
��ŐQ`�Um��
��X��F1��TU+UAb�(����*�E��`(�"�
�VT"��V2)"ȱF"�$
�E,PDUPEAdVAH��B-�*J��TPYm�QDTDER#Z����Z���H�Eb��`��P�X"Ȩ��J��QQU�Ōb����"�"�TdDU�Z��"1PTR#,QB"��*�"�*����""���@DDEY��c"�*��P�Ȉ�@X��`��� �Ed�Y"�,����,�*"2ڂ0U� ��"�(�)�����ϧ�������Gl��Ɔh���Ӕ�ѧ*r!����9;�\e�HkU�wy{w�Z��B�R9n{���y�pw7�}�,�c꺋�jD�tɡ΁g��#@�]����Fx!�p%f�����>�Vv�u)�G[fv��o��x���I���� �ȭ�c���N�<,�W7GH�����^ˇr�Yk#�fU�[�%�b�euL�È���iR�A��}c�py]w�Tūj���,������%u�O�������y1])E�`��=��zv3=:l
c����0�,K,�����^7�>^'f._:�CO�ʼ,�Y�K��Υ�ɫZ����(�ﵻ��5�����ٙ�~ꈡ*I}c"�0v�YŜ�ˮ�O�gU��K�5�NYv�|w������\�D�.�Ec���i}�ׇ�`�H�B}!{���y��E�L�7�I-l�����n�5~����B�Oz�J�2�v1ϼI�xF��d�y
�3�Sk���Y��K)��_��*J�@�\E��t�+�a+�{Y��{��3�b�׳ ��>#yH���s�֕i�")C9��[X9�"�z?w�Ra�^�{��+0�WnOT�[y1[�Hյ޾���8
�6�[ݰ�%���f� 7�h�es�㝆�L��m��e�I���Wuv��k���&:Lvo�[�/���&��(�[ܸM'p��jbe��d��nuA���t-�n@�R����x{ޅ��ܷ���Z�v#b�!�B'I�	A���~>Gg�ޛ�Z(�k���K�)�|f��#�/(�s�"kʶ�@��
�C��a(&��xxu
�ϖ����◦A/#�kWb�\&���9M�$�n�[������/EiI�h���_֦���9og�n������	}��H?|�\E�uq��+K�C����N�2,)�u7�&R��&��-X/�^���~j�]�3TPW��wQjq�ܲO4fΗ1�ל�����m��;�e�����x2������`���h�>����#��Qo#X,Vj̔�^!=Q�O�C��?�eU�yZ
��z��g��%ם�.�o��ׯ�������z���Q,(�>J��Qca�z�}�3�0��(�a�R�։���k
�y�)��Q�Mp��b��h����8fĜ���P��#�	b�w����Eܰ!d�%>>*<���@�k�/�V{w��}k�o=�Ʒק5�]�)؍�E��-!���4
�;�v�|3:hs5�Պ�+�u[�Ud1�)'�OfO	��nȚ��&˖�5�5���m�'�X�l�͛��c�bUIN�H�;�]�v�j�屼�ӣB{S�o`1�[]�L�+�b�P�Hw'ط�v�+�g�n܊��آ(E�s�=�{�1^���n�N�k�3�& �u�0	����F�m��7;Q�cb7N�)yq�)�Kٙ�\D���gEx�tVLӌ��a󰝆�Ĺdp��� 7^wuBy0p�{��:�V��#`��r��%\I�R5۪|4ѯ1.	���1|�L���KUg]�f�sՏ�9Lo��{鴵3�H��i ��p]T������>���9a��+�sg�L�1��/��;H�	�Q@�&E�v8�v��ע �aPb��AuwY���"5��ծ���o��`Z�|�y��3�A��~`8��7�;A�hٝ�FӟC�pAJ�H;)�Y.I��su�˫o;��0Y�,H{^[cHV%;J3�g:᳭ۺ7�]v�$�*|R���"rq>g��O6�D�;�ƬT���C;���r�E�s]9Pؽ�+!����=W���z�J{�R)����7k�G�ѵ�y[��i��N[%Qv�$��r��\���v+D
ұ�Y�ۧ��##̑���.��d3GM��[��P�72Q��ZZӸ�1�FN#f�oG����]�N�ea��e<��u=�Z�'o!�&6ô�M�5��*G\xv�GbnLy`��m���j�ؠ�w�Ϊ�E�
Yb՘�J�(�������F٬�x�){}}q����%��z�[O]7�y�{�꯫�� ʾ]�s�븿(����i�hEsV��@�@�	����嘽jb�W��Tu�J�{��	�O����E��]��n�n|�[X	�sGn�X�q
�V���ԡػ��.�b��b��go�"&"1����!��U�F7��`߮���k/��U���h:Z��j	y^Ʃ�$��	��CԣK=_@W���GD�x��uC�af��mH/:�6��3��컦�!X�bgg0�C�x�f{무�.���q�W�>�咦�F�NF�0�y�v[|�!pE��F�V,I�|
�0]u�j"C�U�W�X=',�Zڽ�;sC]�E��mJ;Y���"֧."�QԓЏ�������&M�G�|�9�|�vǫq��1�e���qJ/�U�:t�a�,.��yЛj�9W��������3:񣀩+��+�,��y!�FX�e�|����i��M�P�b5w���x�]^�K{��`�KQ&G==��µcy)���F�y�&��C�+��tlV�ӥ1�T��r�I3�+�Y�Y홄*`5��8�β�23�:.��x��Q��ӹ�}��S�-A�]��
��{uT��N`�}]ík��ۨ�]�����mɶ"�[%58�Э�Q\�Fp���#���k�yg�7������줺���I$i~*�o)�WGN����(�3�-��s��݊nf]���>��0�FjS#�Մ���D�`�!m��Xi�Ҍ�;���A�ų�]TuG/g�{Ws��xMk��tP�Jf
B	��Y�D-ɠ1z�Q��f���o�v[�Q�����6`��'5�`U���9P7Ҷ���N0U�orO6�wG!S/Hf�����R�4tɮt	��h)��%P�'�����R�����N'Yau���
z���f�Օ��Ċ�btK�e�c[VMk�rdif:�9R�Lڻ��ᜆ�n�!zn��ir�i��H�0��������X!�ꙓ~��\��V�jI�N���F����]���E��P�[ﶀ_z�|&WM.�����l�]8�ۺr��s�ײr�}�Z�<Q́��dF���B�3f�T\�{P��%�B�V���b���x���uU=s��8U�[�<q��8e
��U���ʧ��5�ol��'�e�&�ݼ\�ߒug�㧙A���vS6�Ͷ�ܔ�F�;L�x �NV��44���P���7R�E�P�
�^��+�K7gm�
Z;Β�I�s����b�(9�ن�g���|�($�w���,ԑ>����/N��٣ko/GI㫁YKc�B�����<�]��q��uY?^��&�rr3��~��3��0�;����B,�Յ[b&���_4�q����m��������Q4�`�v�݁_�+����f9�R�W��ʙ���>���l��q	Z�k���"����q���t��u���V��Į�k*��ɷ/�\b�b�g}��$��MGIB�o��1+��gK[Y�:Dgv�r�o$7mnc�[�!2�^d���:M",pD�*�h:��/�醇�T^,�Ǉ	8�W�ډs֎O45�t�J6�t4�y,�s�q�s\��Gh(����iC���r�F���0�#uO/@�e�}Fk�"��7�t������p-N
���� �% �K���3{ww6\-\,@{B���W��^m�xⴲ� ���"��:�a)��i��R3������lh�ǐo�*�#��[I���w]�XP�4�I�sF��s�Zk�X���[<a7s���P߼��nI�5[���Z�CT�+��',�����C�������ݷUZ�̆�kQӆު�Fiwo�Ӳ��j�z�"̘7|�V��S�E3�Q뙥���NK��Y���CR�k�c�*�fD+j�1�p_�g�a�i�6ܱh����|����fp�F�ǘ�����0y/��(d�j��Xvw�<=� �u�����/���n����;�5Aoï��U[َ;�˪�;��@�KA�!�Ô�捻��}�J\�YxW=������i l��3#��d_�M���E���)�;{Y���ˎ'j���z�5�7��9��'/����@UWU��R�F�Y���,=^tN]�|m�].�aL�K��,�o=�Ʒק����Fэ"ί*U�2h[�+2SN�q�2&k���c��c���BM7��0J��%L����^7]Q����Q�s�T���6��y�b�Ĵ�c��]"�@�Ed�8���!�vv��<GG���x�ǫ0t���JH�7]�jU\_�5L�H�pR%x�FdL�>�p��׸�__A�Ul�{�u!>�ݎxp�cNm-I��H�ZM�C�
�J,
��;��s�y�&���e�5���?&z3����g����!�Ӷ��D-Pb��_.�M��f��k˽���l3���'���a�[�֎מ+f���G|��PpAH�;�qrw���Jr��W�Q�VyՊ��.�ʳfi߆@t����ռn��Y�,N��T6���s����tjh��G�/k ��Ȼr���Kx��]�@��77y�unr̠�I�.�2sq�{[M9�L����u2��C~ xx	��k�.��"0E�����B�NҌg:�:p�n��s�L�1�HI�@Ψ����|��x�W �.�3m���s�'�|O�����i�|��6ŝa��O!�d��!��u�a������"��#�N΢���[�{?n��,�g�L@�=�HT��vti1
��y�l��h)��q5���c6���4���,��_��$�:��N!�L
��N}��li+|�i�a�$�I��I	/���V�������u�| ���T:������'ٙ*����wz��VwvLO�4�H/R���~��!P4�<2z�#����'�3��&�8������m��#�fHU�ڢ��ެ��Q��铉�����4�:�b�p�gYd��y��H. o��^$��1 ��r���T��-��I�O��H��*A�oԘ���1�d�>�='��2�t��'��9��ZT�c��? i+6þkvxɈ��}�:���g�Y�4����8y���S�1�{�z�YY+���IS�a]�䘓���q�+����}n!�"H�$]������>����Չ��� I���>La�`���f3�g�m �a���6�H�u+?Na�O��&0��rhT���d����i
��s�Ԟ��)s�&�d�1�3�����Lǽ�S��X�q�U��^�o=ώ��I�6���!���凎0Y�+&2��8������T�7�S�$�{���6��J��֌d�+=�=�t�i�<]׽�� �0����ޟ��ƺy��=������n�P��1ԩ����e=d����C�����c�&��?n�"2u�17��F���'�Ię�:�'ݡ��ʫ>�@�3vs�>�'�=�﷞{�?c�I��Ag���������S3�Lv��3����bL~Mۉ%g��hf��Ɉ�o3�����nÈi+%W�n�H)��K8G�>�<�};bjw�����n��6J����%g
�E|�[[Ɓs$E[�Uq�?����
�/G�vytW�%m�3	{u^#z��Q��)*�W1Y��bn��o�/�%J4�N�Ժ0�Lu���ȏt2�j��6B�%Gv&%�8�ʭ��Լܶ�V�| ��gl�|���'�J| ��y���'S�]�
��/9��~C�ć;�:�b�0�1>7@���3~C�'�i��T��0���&3�vM!RW����������a�%V#�;Өp<�T:y�o,�M �_��*k�N3��gp��ܲo]��0*N����O��Ԭ=k�%a�,1�a��1�Ă�dR���D#��G�t {>��u�æ�oٔ���Ь��+��I�O�Y����<@�T����4m����V{߲M8����w��1*q�gu��>d�J�g~ԟ�Ǭ
���
���11�=�cĀH��e����`Jcb���s��}��߽{� �N�a���Aq��$��1�ɻ1����5���u<H,�g<��"�Ԭ=��CO�u&?0�?�$�&;���EIY����.��&$�y����{���;D�ԬR����,��3�>�E� �Y*��d"��%�׎�*��2}�i��mư*N'ɉ��é6���/��:͡�8���u�L�
Ŝa�3�wD4����o���oꮸ��o���,H����dxg�����*E���EaXTǌ��rȦ!RW��e��J�AL����'��j��u��+%@�~�Os'�W'�s�$��{x~{��ߛ������=������=J��3��w��S��A~d����h~N��Ӻ��6��J�0��Leg9g���J���1�VN�M!]�x�d����@�T����t��3/F��tw����@~RO{�%�����m�����R#'����M�z����{���Ă���䟟wt1���t��)��i��'��sY8��m�J�z:����ˊ��v��[��(}�A��#�l�E�G���!ӟ���*E�_9�8ɿ,�& ��Lˤ�w�6��T������AH����D����<��O���4��Y]�*N'ɣ�������s<��߻�����ĕ���Ƴ�T?!�c���|�b�0�t�Ax��1~���H/���:���T�O=�M��*u�O5ܨJ�I\���p<IP�o�u�-�ɤ�?~�{3`�[������'6K�ח `MF�|�
�@���N��g�����\���p�G��t�rz�[��^Rpy�gW2־�����!OK���r%s�=���KsNtV�(�VevGh�x4>�-�Q��E�7�����d�{����z���O-���@K�O�-�=d�O��a��0+��v�����٤5��R��c>a��l��<g��Ax���ɤ�u>C<��i�E������E�{��>��(�[���?J���q_zbJ�����Ĭ���3�뤂��'���f$P8�>M���L���oW���N�? iĜB�2bc���@�
Da����m ��~��5�'�H�<���3kNd�6g*�_nҽ��+=���>�g>�c�AN�9���N� z^�Y�~a���+��Y�1����$��<�4��"��g��V~d���'L�&e��~��<�D�������:����.�?��
���y���뤂���m�oY?r�a�܅|`T�'?w�<C���}�~�i�2��~Lg��,�
ş3V����"��g�1 �j��DA$	݈�87�]��6�{�����aS��w����V=�6����S��$^v���&��i�{d�k���2T��u�R|��S�{��|��hW�=�Xi�k�)G�>g�#��t��c����'����a��q ����14�S�bO���*(o�a��d�+���h*9�	��}i;�;��Az��ɝ�AH�u*xg>ԟ��%a�s2q+�&�$޺���W�zy������_���M!\d��ΰ*
Df�C穉��L.Y8������:�Nr�>�f@]0+<��u
�I�ğ�L��E'�������q=&��׃ a�}�w6UO�y��y��ϿwϾ��t��YR,���*i��.YԞ�@�Vc&e�P4��*VjZ��
��[�N<t�uf2c�'ݦ��S�4���9��N&!ԕ����D}��8��I����L�WG����ܷ�4�B�g{��C�� �a��>�x��1��߳N0�LJ�w;dSV8���M ~J�b��$�Z��~���(�P8��}�>>��>�zx���:>��L{>�ӊ{{���l�~M��z�����zκI�
�Oa��Aa��7�u�ԩ�a������Ă�E4���b�&5"ʃ�h�1�d��-�s�L@�R�W�Y;h!'u��}����#F.ڿ��?��/�m�A^�y\� ��,V(f*"�D�W�J��nb{���$��Yj�D�$l�Ca�C0��CCF�Y$��Y������Y��Ay�N�'�<w9!5���ZWa�۪��(�zֹ~��f�zk��/�2\}2ݬ�n��m#��<�;I��z^J�us��[Af���B=�ԇ�!o���&�Ǣ�H�펽i�K횇eB w().���wu����c��Ķ���f��W}�a�9'V�U��Vw���խ)�OR��bfʎ��a���E_rϣ�3�s��ͮ��*�=�v�5<����/B�\9���2��ۢ9����}Z�y���IEa�R��.�Ns�I�}��<����Kl5睄��� I�d8)�]���^��R���CUnk�'����TǴ�O���6�e�f>Kn](��D
�1,�Ԡ�c��,��]�{���}�ŉ;u�B �3ek>���0���v��AՊ�ʲ��v�F��p�o��;Q�,��A򡻠V'&}]�i�J�Y�X��7<F$�V7��k���N��+�]�\�z�����K*�*��D��6����S��R�u�Lf�u�n���ʞLx���짨l��ƅ���C-Br��Vv�<�6}}�.��g��م��<o�V�u����t���}=]�n�k�'�+�Q�Y��EM�rU��S��j�w̱�i�v;�ݜ'5u���uW$�q�-�ݤ�M9%wv>���L/�����	W.1r����H�â�G��9Oe�\k���J����ۜ.��}H`\k'ߺv�Q��ݘ�T���7^��ڣ*��R��NE�Vqn���.9x�-�Z�3���/��s/�z%XYo�P�L�P��6]B�<�AWZ�����Q�4z��a)Y6��Z�|��(H�^�ۼ���4>�1�Xͩ"�����&��a���t�IǄ�>>�t�q���Y��B9g��Vb��s��.>M�=���˫r��S�N��������J ��Al�w~��+�t^�ʸ2�^��ABz:n^����+����\c����w�P���Q3�>��>���cHod� �:�h�Cok��ٛ������#�96''��l7�)�]��:��+�O ��Ƥ�B�/\��i�4MK�v��$Í�-1jr=�) �2��ګvjJ�< c1癠<؞�[���!W�nQ��3f䕵n�\0�b��Io
�,\��'A'[/�}��yiŖ�cɪ��]4+��`i�F�_{�����K�;3�r�3��`�c�W;��γ�z���	.j"4��n����:��T����+��RZ}�'Ʀ��z �-'&�_�P���A/E4�ەL!�H����΢Ov=(̓���T��+�'B��c��L��gmi��� �O�E��0QYTPE��dUQQE�"�EU"�#D��(���(�"(� �UU��EU��"*�Xb��U"��Q�AdQDPUKlX( ���dP`Ȱb1QE����$X�b�`�E,QQEb"�DV(�ȱT�DVEm�2*����Q�Ŋ,
,PX("E�����k*���REQF���E"��bȊ+�Ŋ
(�1UEUUAE�`���P�((��QR(��b��A����)X�)1UV"���PQ�����ȉQb�EQV�aY
������((*�`�� �+

�`(,PXH��� ���R)E�*$`� 	�W�[�����J��3N�����n��i�Fsz����Q;d�L,-��,��<���p�\�匞����k{6vlB����f�m���H*A~t��k�z�
E���ގ�q�q�������'S��32'�+�'{�6��PR?��5'�S<�Ԏ�x��Ô1�8�����H�A˿����Y��S_]
n�[#�i�Oi1���|��ě��bAzϘoϳ��!���s�c�T��p:�g̗,��2m�Vu���Rz�M�wz�j��P_9����=�D �w>�{3���v�ZVn�ըt�4�\d�tհ���+1�'ɤ>I]���i�2��=��q
����a�������3hbO9��C��n u+
��P}� "o�!=���}�KOֆ�t���$�{�h)��|�]�)������x�XoVq>ݓ�+��ٺi'�~B�~� i��g�S�T��3���Ox�&0<�����$A�D	?/�N���~���Ͼʷ�~��H�����d�JɹϾ��3��+�U �J������$��yhz�"ɬ�M'Y=q��_f�&�Y:���2bN!_P��6�|`R (�N�9ɜ2�~k�8���#�bAz}��;�u�c<��&�:�Mxw\�T��}��
x�M$�c����u1�!�Cĩ�>f�f�Xz�06��Ǭ���'L񞉏i��}�~���H�Y�~� �+6�O=�����;��4��
�r�E:�׎�t�܆��J��^{�����+��^���4��'̘��ʇ��i�i ��Tݫ:����%���dG�3�˺ϻ�z���@l���;�L}a�11+7혁Ĭ+}�~d��Ou�6�o;`c��AH�r��{���P>K���r|�������~O��m����(i'I�=�[�G�X
�"+^}����`Tkٔ1�J�Y�(u+3�bM���̊T:�3��i�E�4{�<��*��f��l�ɜ�M$�Y>�7�u
�_Ͻ�u' <O�w���V���r����B#�����O)�R���f�ΰ4��W��[&��7�2u�1r�gd��1�,t���߰yCi�73�
��B��:�����~R�O~�\��g��ߚ�D�4�^�]�d��;�m尕�+}tFri�zN�9�����b�B�H���Q�o��BV��Mժ�|_�3���Wjމiysu�c�Mnuˏ�c{}ê1�UN���8ݒ��=�#3:Ź��=�X#4�ړޗ^ys��^i�Vo0���  �����s�?����?��扷�!����4��I��Ry��8���r��& u+>Om��~`T�Ot�i������)Ԝx�^d��d�l��=��:��Uv׵��m����i�	S�(��¦'Ɉq%|�u�
>eCG;�ĂΡ�y�E��|���N0��3���c��&%u2�?%aSRى��L@�_7���y����@�#į��qr~�ed�sf��w���~�4�AH�v��퓬�z�_yܒ�wd���=�ܓi+:�Gϰ1��PXs��Lu*Ay�+SL1����Lk"�'�H/�	$�z�9�ovB��wUÙ��w)mޮA� ��#ޓ���Ǩ�#�z��y9�N�R�s^�d��"�g3!�T�'��=;܆�1+��g}��*M�_�ړi��
�v�Ddǩ�>�edm����}�߳o�}�f�~��t��dx&O���Y�I�)�?0������'��y�?%H/s���!�;��ϒc�T9{�@����^�z�d�ҳ����<���Rk���_{���uX}]�\�Fv|��E��ނK>�$H�I����X��_�ա�Sl>a]��t4���ba�린*>eM�a�M�q���6ŝa��N����c1�C���_�8�'�k�e%*Z����̬y��k�G� 2V��ޡ���Ɉ�k���RW��3���*
E�)���h)�8����c6���HO�����偉8θ�߹�ۦAM��;`�IO��϶��+�Y���j*���?a�>D��z���<dR���
���OӺ֥A���T���<egwd��}I��Az�6[֓�*�S?�=t���k �i:����& q+���c���	?��
s�T�H1�U��g��~d�c�z{ܚH��q1���F�>��SI���6�=���g(AJ�O��g��Ag�,��H#�u&>0�f�ޮ�t|>S�Mh��?{N�Q���~@�+=a��`��1�_�ì�y~`V{?s'P�VJ�0ߝ��
E:����Aed����R_���Wl�}I��LLC�ݳX�'=����0�4쇎��{WILv9Q�w�MB��v~٭܆PuS����:~j��+�t�)ܤ�u'�#�+�^���:�]	�)8��s�=���K���V�{�����\�!����o�ǳ��M��%ݪ8��H>L���ځ^ޝ��\{E��{4%�m`�� �� �o�r�;��(�Ȓ<	l�&,������/Xx�3��H/�8�n~�G������4�I��&0�s�:�B��ݲz~�$�"���<AH����=M��m��Y��a�_]9������Ϙ��@D�{�GmǬ
��|������Pw����,���Y�La���UH/�����������4͠�yy���V{�&{w@m6�_��~lC�~q�ҕw�P�������}����&� ��)��Ld��yOY4�ԯ��ZM?0*NxoO��L~@�n�"2u�17��F��~����Aq&��|I�hbC���lb�w�r:����O}��A ��A��|�H,�;;�� ~J����i�>I��~C=<���I�ɹn$P8��3v�j�̘��7���M���_�q%d���m& �S�h��~�uv�꿔tWΚ���B>�<	�ｵ+�'��L8»w��u:��w�M?0*�Ɉz��ćNwZ�B�f�~LO�1��!���o�i �a�xZi4�"�Ļ��i���̘�®ﾒ�+�?W���'�~�(�z���`x�hT7�0�{d�i"���%Mv��c=}3�J���Y7��So'Y��5��!^0*?�Xz�>J���0����bA3Ĉ��B�4]�����׭���4�������i����Y��'�V9a����H.���d����~�4��OΐS���@ĩ�M��ڬ���q+{�I�m���Ԩc������2/o{*>���m�� <A���?26�2�穴���?:I�(c&�\`T�>��M�p�y��<@�+C��i�Τ��'������ܚH�i+>+��|�,���5��W��0���c���G�]"�?2f^�yˤ�
����d"��-<v�YPܶc����L>Cn5�Rq>LO��I��Aoi�i!��N���Y�S3���/�c�r�U׼~�f>����}�!�Av������<J�@��
°��1�"�
����KI��
���l��H,<��%�d�1<������(o�����I��O���h���X�7�$m]���;�����pm6�4��m�;��:"��7����b��fK�4��݀�I��A,�ֳ��MѩrӦVb���QP��c{��L^���`F��'Qՙ5���p�ܝE9R���ئ�e�Y�4��������k���̮�K�OP���d5��%O��`g�8�ý�N������Z6����}��"͡���9a��&2������J��+Ĭ���B�[x�}�4@߳�5�^N^��k�x1� Dhvy̟>3L��Ú������7;����LLz�gs	��2h>�5Si��xs�����1 ���䟟wt1����L
���LO�<LH&�j~��7�SY����p?a|0�(�>�U�Y�L}awB��x���a��@�W�s2o�6Ɉyy���u�2�'{f�u
�����*ANO��D����<>���'5M0�(Isw�>ϑ�\�����go���zȢ@��@���x���5@>I��XO�i����g������N$�I�ϰ�"��o�,�9Ϸ$P?���kX�����������~��d�i���b�r��7t�*짆X~f��
�z�g]���$�7f�5��R��!���S��<M��}�bT:���P$�G���j��z��]v���=ǲm?2q��韹�1�I��`i�+&�'�뤂��O]5�P:�>OB�z鞲VM��4�����I���B��bc���Ia�o���<	� [����ӈX��x:����_�vO�~�����hc=�ܓN�&��4O�:�����'�1į�X��I��S�1 �g���X�Ʈ��%ݟ�1<���i�d̨����I1pr���2u|��Yc�G��V�4��
��֎��㤂���m�oY?r�a�܅|`T�'�{��>I_�ӿjO��1Ɍ�E�!X��jZz�H/x��f��H���Hތ}���xI�� �����O3����%B�����ĕ
���4�y�'SHz�HK�'���O�%@���\u'̯<{��|��hW�=��L
���-�]�M9�]�7���T��A�L4��2gSi�y7a��?'�bO�ǉT8��y��6��������h*��&�J����;��Az����5�A@�T��}�?>3�B>�޿߶��ܔ�$733<��8Ɂ}�R��{6٢%����=	�v�j�kr�#�V����T[!�k���� h� �n��Z�XY6�s���I�ZX�9+�.,��gm!�x���ְ�\Ѿ�y�V�❲��E��j����+V�ĕ���s_)́ΕsO*p���x{å,)ٟ�Q�b?�2���*'�$�Дu��}���a�c�R�k����n���sV>�ʃ{�l��ZS��RQ&O�A�:JuM�g�� ο��]��A.w`r3���&�Ԉ�������I�E�D�j��H���|�v.�E��-{�����x�Qq���:c��	��O%�4m�!�s\�9GN��H�1!�8��,sk��sV.���[\��E9\��AӔ�g��q�QbeF�����Ic S^���1�N�@z�Й{���`C���ic\Gt�*CXa�����7^ő��T9�]�}j^��:��׬�wT���_��V�uWp�W�.��u�E�	��$�2�*��<ڲ۾�ʇ�x����M�������;����2�Xw��vo�E������|���r�U��*a�@�D��*&����7g��6B�9^*E��v�vy��O7w���[��ZCd>�xا1x��K�A�΅�Q~�q����Ezad3P�U�g�$;g��d�H�����	Y"}W�ңn4��8a���g��o�h�\hVew.��Y�!�I�i��L�e.,�K��=��
 J\[�18�ӧ:�mlw�(����<D��l\oɥD��TkHڙ��Z3W1���ׅ�u������2�9AWo�<<<&�r�����߆R*�.���UP�c�Hz�����7�t�ؓ��NQ��-;¥�]�A�r��Z�VU8���^�Dϯ��3
e8R꽉�~ӍmaśTu)�U�4�9�۱m,[�j�+⸏�-"Zf�X�<�� 5�BM7��eK�	������T�1l]v��=���}�e�[�Յ5'P�S"�!�X"ڼ��^İma_i�v��핆ؼ=9�H+�j�Z�O�Z���3�P�����Lͺ�Dt������mzmv)�i֢y�=�YZH���.;�_C]�xv(k^�m-I��H�F� ��F�e(3�d�c�����\���m�[������;�J�[C\�q�m5�B�t�]��<���$^�n:[�ȒK��/�2���p�v{a{��x��"2e���+یi�����ٶ� �ʁ��K�v����m�
�;J1��C8:p�n��0.��b��>�i��e���_*�H�����6�מ��%5(3f�j�\kc:��q�7x��:���+��������bʶ��=�elBD�j�����߻�����rV�3#'�����P�W�b�5�1�:iN�Ol{e��עe'y�����O�c� �Aes�e��z�Q���q�x2��@�qv�}����xx{��E��z�D��FH�����,`y����1��<���k������ƥRFEӚ�]+��&���I	\",Is*r\�.t42$G��ׇ�4�:|k�Sr��]�č�æ�v/f���m1v��gu�xt�(�9�n;�C����R	�;!m�f��w7(n�=oOd��i\\-<Z}��bjo��pjtH���)����ۣW����μ���oy�����⦡t�<^"y,��F��F�e�$�hk�>�k/ʯx�gmnnF\{�ܴ�:im���2�,�U���������vR������ᤃ��ZbŪ�R�k���4���v?	W��������u���j��@��q�]���G'�fs=��T��jȄI�1����gTj�`�ĝ��7@��u.�����:�8��k��4�{�S�S��w�l^��h!�,�[�ׅw\#�E�zuq��Ig�Џ�� '��a�NQD�}��+�l�/�H��Ks��P�qJ/�J��4�6��''S�x0?E*��k��܃��r�l���ż���8�E��n�շ�V�ɛ�+�73����.�`�O�w�ޥvd��`�d�\eNq �;{X!f*���W�$��)�̍��:���XڏY$��&�㙕�N��5�E(5�{��5�m�jV�BA�ݠ�G��R�RF��Y��d_���zm�IH����n�:I����]*݅���#��M���P�AWv?\��ƭ�����=K�x�=���U	/!�qm؆��B�@�A��ߨ����dyw\�a�^��;���h���t��s�۱V��F�*(	1����P�/
5T�Ѷ��������`۾�ec�C."�7N��Mk��Ίk�f
Vd�(�'1N�T�
�w*篷6[�rh�q�}rU�H�h6�yā��9�p����"P�����:^?,Z�TwE׍��̾"�]��䫾�%�P*~�\��p۝��f�^f'�`���$8υy�u�kTU��o��c�\ܲ�1Q�L>�4�]�px�V�*a=�@�Pe�³ژ[ZlT�Ӹ�*ë;����+��!�>�V��$��8��9le�P��`!���!(&Bsf���C�U�8�9Xn�g'�P�[����4u��#oR�Ґ�M�s2��zҼ�����Jݍ�8��|j�������R�V����8�,Ϭ:�NG�ћ7C��؉[��-�(�,��[�jS>V��~u��4���.°i�'��2��鸑��H�2��Fvrã+
�'�����x=�S������hϧf�@��k��4EZU�0sV�,��\DJ�b�ﯧz�����ܛl讨�c'I�b��Tt�r1US�:3�X����� �#����{����m��q�����wdT��y���EA)@M�^���(�F�����5�C��;5q[2	F���6�'�.�)�͠䔶`�w��7p���9���|&�_u>{u��&ov��L�p���z�J�3�愢�N��g�B�y��:\�+Aee���ڊ���f���hM�����U�v�k�RNU2hGIB��7ب�k�&f�1��\�����=�v8��s�Ew�����I�E�D�aV�@���|�:m��|�};fz�W9�8�W����E�s�s���O%�4mځ�>.,��	�o,��I�:Mj��.s�2�2���pA�*붧�<�r��<�p�ݳ�gS��FԮλ
�ve��.�d��_,C)/X@���.��]��!:��~�B��6�<qZ]�up�V�%'ʄT6d��L��Db-���+K���֍k��x�Jj��Wq�4����7f�3I.��Z����^7r-�ٽS��OmK�d�+:lg�v�� �:�u��j;�[���:Mb��l�y��x}3w���+���v@�������ؓk�F�FV�#��gM�I����xJ�f��q�t3\PV���-@N ���<��#^��喸���,-�XGa�yl����_��`�k�pJ�C����s�]k����^��,�Ey�}��s�0D�j��kꍃq�xϣd,�-�����T�_��<,)Pf�>��*M1}w�XNC�11Nb�9�nQ}΅�Q��o�����B����gvV���%�ǫ��ּ�+ذ�G�Z&0�FJC�85�7��8�6$����p�2�xV9u^�[</���6�o���C�<��>T��񿗛�����q�k}zevEe�mm��۾�Ԓݚ���ŉ`8E�KHv��T`<��Bh7��eK�	u^�C�t��u�̾]_��Mg�cu���tTt��S!�}z�U_/c��0ߪ�nW=�����4�c]�qr��������ϭB��]q~5L�H�Q%S4���j��U�eG{��Y��w�Ҋﶾ��K"�	��&��#�i4Wt#>����V�_�)��w��#�Y�H��v,İ�]����	�)E�#i�V(7�妚[S}VD�l��4ժ��3��<V՗�\Cި�U
[d�\Db�,P��"sZ\�u�)Y��R��p��Ǘz$�kF��N����ٰ�mHT��_'כ!�sC�S��ol�i��T<{.c��N#u��I�]K��Y3�ػZz�MT�qQ�|��j���qes���Uf�"��8!���!u���K%u��������	:��ģ��f��� �KS�/�
xv�Y%� �zl�W4���8jc��:r�]A���:�;8�D�J%���U1��J֩5���M�sc�u�:\ҭك5�vx��uN�X��i'�8�Jǝ�g��p�ں��f���&�3���+��-5����΃'"u�)`{�9��b��@j�7 M��N��\��(V������C�%���r��ܭ��,r`6mY���%+H�U��w�M곞9|Qj/�G�Wy�*��̱���R^n�͠�\_G�B�K[���ĈCf��1%\�N��O/{��;�K9���)q�ϐ�Nj��f�u��0���Ѹ�I5ދq뙯�}&��[ɵ��۫�-^n�Z9 ��
��D�!n��9m�r�E��nL.�!cTk��r���B��+�LؤS�x��%��S�{��a�=��h"�t�&�I�M��� ���{By+�O�j�C������ְ�8cH���t����������:V���d�ۍ�5���E�N:�^�s\Ҫ�39�7!w�Kx�<�Q�/��SU�1	�N��Ҥ���o�Gv�Z�D��h�k�F�6\�Y�s��?,���S�X�7k2�Ѵ����rRl���ήv7�*e
��|.� ����E��"�.� �ӱ��/�hh�)H�z��Ψ%��6zvt8v�'Jo˪�������4'*=�:�n��kݪj�zF�n�K��6��Nlk'm֬�w�e��9�����l�;WR��+�w��>�$1s��H+Է������d��Pൽ�'��G�s�N�*�X�{��-v�����B]fDw6Y���;����Bѹ��(�	���]vW]�>�d��̧.�HH/x>��Xء��R���Q �I�J�Top^ia���ɘAo� J�ԝ�љW� �X��:�&V��C'S:4�ϓL���٩8����P[)���s��֦k�u�B�9�NJ{L	q֗b��\EڜS��ki�R�F2oS��{}kZ{�rp��X]2�K�2����V�Ż;�,�9w^��}�5*�����%�#(h�������*5�v�l��hB5���Bmϙ��}��^��e�5.��y�%��wNnj^���CjMĬl3�k;=s���V;vJ;9��o�䬖�t�-[$�O1�y�}����1@Qd�,X���QEP��#�dD"��`�ł�Ad��
E"�XE" ��,a`�IU��UQR�E�X""0R�(�*���@�X"(#����
(��X�Q�X�)b�AT�$��A���
AV,���H�T���X�����E@E��H,Y"�i�TX�PX(�P���b�"�URb��DH�EAH�
ʪ���"�,PX1��D`���b��"(�5���X�d�,��TH(��DUX*��aH�
�+%# (����*(
(��PPR)��TUEH�-�U��,��˕+we��稬G�9�u�ׂet�e��}&���-��ʆe�Qqá��3��Ք�`amA(_#������)�a��TVu�k(�O1��q���t�������W{x][���З9BK{S6S��wg�c��9>v���S���u��᯼wh�'���j2
��ۂk���4���A�t3*`JK�nD��w2�u�<H�2�]m�FT���lϦ�+]��-}"�g)����\)���k�{�i��:����㰣�*j|��]G���U�{MOUFy�Z���T�i�a���''s�4:���If�)���0�ës|O%<��L�L(�&ā��M��z|un��K�ߩiW�p[.߯TG!�i��t��G]x�qV��6��G&L��0����s��%�tg�+~	e[<���-�O#:�(�X�7��}?@�)�douf<j���~o���Ea��IsÎ�K��g�V�$�\�[U�%�B`��K��.����旂i��e�F��:�Q�K��[jq��:��;Q!>�#��7(��	 \�]:��37��P���mN��ە��������w�Q�BpVw&���O<1�ι0� cv��Ɖ�����m��=�9�G]㦅nr���+v�'Xr@8�>QQ��A�b�v��o�'s�lS��m�L��&�QQ��$�����/t�t��	�h[��=�&9[!��ͽ�}�����I��mІ��ù����k`Bt�V9����Z�TI��#��c���J�J�b݀���6�CIߊ��Zt�yems�V�w:ق_�BA״�*�i_�L������{�Ju������as�p��Sۘp��|� [4It�_��Y��w/7j�&{
�������}��o�i�p���1 Rw�X��ֻ�/Y�箒{=Z&j��X��yNi�ӵ!/%���ak�G�҃+w+z�=ĺ7�3����p��17/7�g6�PR�Җ��o/J��k��۷�����m�v1#�9I�3aN9��i]���:��.�R���(ǫ�ok��FO]n?K��U�kH�����D]�r��ߕ<�{Z�{K�=���#�&}��Ѽ�'r����ev��&����Qf�+cI���6�s��G#;®ڀO�.��A�1��A*��-��#ŉ^�v\J�}�w~��9�8OǮc�&��Y[�U�%S^���� sD��ɩř��%��]�)
����Q}w
��Zά[�w�&;���p���
^竞��WHf�?	��ڠ�}}�g�Oe#��qӮ��Ά���Fq3��k�ÎА�\�f�|30B��%Y�/�meg�O;|;�n���s���9[a*z��p���Ǜ8�����S��M[�|�-��\#)��u�B=|�Ў|�L�Xx�[�=]b��|�V��Y~���3k���5k�1rwUt�s�}�8��v��Y��y��Z�9378�i0_u�Ba�J^J�
}�;��E�cSTڷ�������;8��ް��b�0����&ZV)L�SN�okX���/N���:��:|�N�]���ܑ*} �4It��ظw��[�bK��b~Ӻ�Wi�Ǹ��F�o��\��X�$f���F����t�<欜�c�r��;y�|��e��۫���)M6)J���H�k�;*��K$è�wZ��N�ߝ��Y��i���έ�eLZ+k#�,��}ڤpSгefK> .��yӗ�GL�n����c��k�>��N����$,��	������O9�޿P|�w`Q�w<�m������C���נ���RꈕN����,VA~9~���E�®M&k[g-�Ol3���թLDY��"�<�n�\؄�I�A���^��Cs}��s�֔�c/"�nf��WK5�crsJ�s�*;Ek���̥x����ܐ�E����'<�鞮�v�c	�n��8+�9��W�܁�_x����m�^��V�һ%9����ި�l(m��Пkむ�xj�0���:���-��Sr��޲�������0�ӊ�<��_���|��r�4�Y�ԥ\�KW����Or�U�:Vߒ��5ˊ�����ٵZ�ŉ4���Ldٖ��*3D�z��|��vL�N�w�؆�Q9*���M�C����綖�F\�XV<����fG6=W���C;�YQ�kz�o�-e�s�n�Y�5ד�n����,�=+�^��d��J̮�ґ[.r͔c���3��[��*-�����m�T\=QF���-V��0��$�z�/�W��Y��O�D._���-d�q]�.v�b
o�^��WN�ڻ�\�v��=�����zq^�ǚ"�з�=gT��<�l��7x��x��3��0<��6�}�v��K�D��P1ݹr_W�������w��e{���}�v��7v��]��v
��Zt�$J�����rT��r�m��ξ5l��]cd[C&��9��뵼��x�L��"�*�N��\����R�PV`�n�V���1��g$;NtQmq1^D��mW��To�{�u����2
 ��M�v�B}֢�(6�rg+2��ߌ=�=��󝯭FJ
Z;���}��
����Wy���s+����˷��iŴ`s]*;R!k���ʠ���F�3��b]1S��SI&]�sFӃc����|6�uf���s`�	��b�����kX<�s"����H#���E�
��ҋ�hN�~��9��KV��͹ܬhge�wX�r�ښ��Y	J��)aV=v���Ž�4�#��ZOnN�`����'�5�ʊvV!�a��nH;���u��܆~��Z��������������xL(M�|J��8+���n6�m�}��V.���eY[��w�d�����xba�n�Sh@��-��W���}Y��$Dʾ>W�
�=�#�������~iR���!���\���[&�vn[K6r���}@�Bnv��g(bw�*�R��L���u��d�x��ﻩ�V�c͝��$WE��A��zfXb���J��n��MޓϗR��n�����۫= �5
*�/N�U������3�U�<1ײ%P�ObM�M��7�%����\K��quqr�L�k�Ro$�1�^���V �w������CI��Ƕ�g������I�7Kjd����`�|{�	��a�t�E�sy���߃ҷ�\m�*�3���;i"T��N���Ѿ�4J��'t�+��驳~�gKTu�x�*b��=])���ܭ��ӎu���P��;����-^e\��V-��-&Q�.��1��K��d��{ُ'˾��2�QW��G�0Vo���魮�d�5���U�=#_wa̺�q㛌���l��ޕ;�	�7����*��F�~���<��$���)��␟��Ah��k����xywK�����[�ո�y.t9�v�*^JH��g��7��pbq'��k+�,vͽ�ɤ�Ҙ1W����;
09�()L��&ެ�]�`.����wYг��w({-���K��kJ~pĎh�x'8˚�&/�;��N�g[����%c;S�[�R�VZ��z�$�hZL��ۋ��ځs��969�y�L"j��}j:�����2�[����SW9�a�R��A�W���g[�f��4�5�ɚ�H6�f��Ҭ��V��äFf�S~�qr\��)Z��<}��k������k7�P2@�o��ct�zo��N2+�^u�����?���KƵ����y7�H8�M�yۊ�]*�/b���r�}[\�/~��5ƀ�|�yL�Xx�[��tm��.4�a�=�#[����Ԭ�e;�X���{NWG[�_Ϸmgj�#dg�/�P+o[5�N���Kif���0*�[K����'����%
��+������;�����{�1�x�8�=^ۆ����Y�T$p��ř��ϧ�v��Q�x����v����=R��(g���72�b�L�Z���#���5(���}��W��el�K��d]� �0���˒*�EXy�'Cû��Х�FsvWoXZ�T�C���I�]'�ʔ��έN{w���[w�./r��)m&c����Be ��̓�m!�+5�~w�m��Xe�WnP=M���c��tד�oN��)�h��^�Ki��so^*z�L�y�ؠ�{�K��c���m<�4�+	�S[�Fm6�b���;C/ϯ�ri[�������ͱ!p���T��|�\���SQo��9Չ[�0' _l*��i�����E�g@��'�?^F^D�������4d��AM�痞�`f򑼉oP��8����c%�,L�&��G(k���<s�o��r�%}�1}�}�DLǻ����O2ɯU�8�n��K�Y6�S���A+ݫ�{���#)�fl�V��u@В=o��\��u�8�UC�����/Σ��9Cwv����-M��-2�/-^G�ewhނkt���
����W5�y^
m�7���1uU�|���*�
)�40kサ��w����˟vS�l�A�w�:V���dk�un���&+t�4sW�:͂FU_X�c*n��^$��CjX+O_v�U���GJ�J���.(ornL��r���y�'�Iy�'����w����|]��}�όO���7�40�
�;yNi���#
���P\h8���:�� @y�iy�#�\�J�W���{7���:�Г�m���s�*�Uf5T�5mY�gnE];���������`&�k�]���LR$s� �!��G;19*�2��g��L��������k/�R�N���rD��fɖ/i�G���I�K�sEɖ��E����}�I�5��j{=����ɻ��<��&�1��:(����6��U��
1�ns^\6��"jx��i+���7н��]i�%������\JI�ں�
\�˨*FZ�Օ�S��e#��7�Y�Y��Z�[���	<�6���5�7�'1p�Ax���N�5��y��ub瀙*�.9�%�<Rݹ����--���a��i�i�Uk�r��UM�����E/j}!f�bP�Y��5��2����3����j\�s��FJ
ZF�<�jV��une�ڭ���$kC��y}˙�1P���ި���)���i�7.:�6���W�se���b��c�tuM�-�4h�plg�<sC��B�Λ"�n�N��jw{6�����S��J��
8&Ďh�קVbڧ
�*��5�{6������*��.]��j�˫V;�u�L8�t��e���Fwg{�?>b���3jA2������}����:�����d�x�tw��,<e�js�EZ[��M��pc��9����zy���%�}[r=�wT���kE7�*;�����o��6v����V_*���'-9Yj�#+cٶ�
�x#��q���)m���l6�lc];~�<9T�ܾ�ʲG��rI,׮ܹ�7Y��W�������Z3��-ٜ���ץ�[�P�%����vvjK0JH��*n�=����BZ�m��j7�@Y�W(;{��.��(�F*��KXy9q�wF-���EX�E����=y��k��KU�͈�d(�y�c3u�W��	%�o#��q�hN�(��]���1qH\��}���Y���uay��԰\�+tS�)mϗ]���A���1��q�p)��a�]МVȯjQ�� %�TbV�!{�V��+�; �i��Z��gt�{'a�x��YC�)ZpELٵ�h�@DՁ��g�Ԭ��(�ٶ�
���^_+����<������:&$���F4��{g^Iq���M9J�]r��梆��>jWi�q`��7�6*S�m�E1nn���;���CY����	���2���*!�X��7aQ'��]Ί��WR��z�`w5XJw��kqr5�mC���n��d"2E,�W�v"�C�o���qq�����
��ϧ`y�H](�2���u��WN�t��{%*�2S����j�T�^o3�w"Pj��ɝ�h��P8�3X+lm�]K��0�e�(���-��f���V�{T�­�D��!Ƙ����I��[�K%���t*@�Lځ�M�����i�dn7�c�[�kk�[z#���i�=!j���X�Be�x�*d]Kdk��sӡؽx��*�:P��P`[���u���[�t�XSݚ�,
�s��dCY�j;bZ:sf�N.�!+��M�@#ٜ�7W�Z߮��*�m�i�Z�Z�:Y2�3������mx�<�9�Ft�����_�ۉ�ɸw����U�2Hv=7��������X��t��1�᝝`V�D7N���)һs5 ���(���C3lH��������9��+����i�G[b`#�c��X�]�'�3�τ�]�x�2�$WS&�U�$�E��vY�xJ.n�,:�]oh��LWa���C�	���*a������0_ݪȧ�p��i��|�N���X���#��je�^P�/�����h�����������5�sZ�m`�q-��,՟uӻ&���d(��r�d�O&�5{
��G���	@+�x肣���ݝj���ښ$+h䫏]���2�P��bu�r���+_����۟r��9��I"Bʽ�%Z��ī����Q$b(��hڹ��9>ǗƦ);��]8b̂�48�ٽ6��=�zX�;v�=�����v���ۧ�]��P\h*mgnXt��Li��)CQ��V�욵J�&�vGt����Û�>@�N>x�၌�S�J�إ�W����:.ݔ4�ۼ�Ӳ�L���ئ�VF,�Đ���=�Xأ��R=c�޲�=m��,�ażm.Z��f+6!"��W:L0�[�f���u�*2���u�����F�
��V%*��n+w��O��f���ٖc�.r�<N^ro�<㏫�T����E��Y`,����)�ز,c"�� �dU�� ����UTb�Q��V,(�Q"���"�DU�X*�#YR(��"�P+���H�Y%`(,Q`(�D���E�ȰA+B�Y# �T"��O���Q-
��� �aE*"Ƞ�*X�f3"�6E(�L`TPP��Y�`�R(cU�"ɉU��¤Q@X",�1�!2ՐU��cU���,�b"�QT��"��R
�,R)*J�`�%��,��,YRAk�b�XX�TA@DD�X�R�6��[d�(,����l�c�����_��g��^;��R9Ь[*�E�dU|�־�0d��U���7�s97���LSmM|'s���/fLP�� �uo�e����ON����
�!݉79M��0�5y>u��]U����{#j:�{��_�=����Z1J�b݇���چ��!�or�C����z��[�����4L���=0����������d���o7wa'�'�a��R�i��v
�v�.}&����_Ԝ���^�Cp,&��=y|�oV
ھk��g���Ni�ҴΗA�)6<R��<�S���R�H�-�U�w�l+�V!4��y���yNh9�v�%��oA
$ü��ʍCj��K�D�K�ά��}ɥnͦ���ƍ�=YzWK|�s� ԰A�ޘ{x2Ӭ�Aw9����c}���c�*�B�1֭t�R�+����kà�GjD-ɩO(e��ש%3֓01w�,[���|�玾Yڌ&i4lவ%nr!�e�U�k+:�uv0�k#�`��֫'�H^E��P�O�7	a Bt��e���H=�!�o��)��]3�jﬅ��0��6���.�pgK�DgDc�Ʋ��['��:����[�F٧��XRL)��eŕ�਽�s5ժU��TV�r�&z�k+��-����N��jv��{�s��Z/ֆ�<U�L�s�7�ı[V��u��ÎПw��?G�PI8 ��}n�b)�{<�lNY��h�z�:V�/8Z�7َ�o|�㚩�^�CUV�x���S����zZ=C؅�㞎|�L�X��c[�	�^���\���벍�L]K~z�OW���&�! w$�究t�=��U���7�A�L>|���`N��t��$߲W^A�V��9n�wgr-���uS�΀���WoZ�ҬT%��<�-�] ���i�Y2p�͗+��w��1�{���m'`��a��6���WBA�Fˣ��ȣ�Z,Lvu�YERy�5���k���v��u�䜢������|�wB\H`�	�-j�dv=��w`Q�w}��yc�<�F�n�0k��T�\ӓ�R�Z�as,֑0ŭ:�)e�3*m�뮍����.��n\�N]��M�ty��N���b�a)w���s:���;
��v��%N�Iw���zk@�r���#S&Nomc�׊s�C�X�k��N��s�k��}�7Dj=>��Y޾�T94��/[����F<�Jե�\T����$J����b�){B|�v]�{&�����
�`b�����_�tZ�J�o��u5G�g@S�ht�͈Z�^{-bm+�|���S�={��uBb�T�i��ؑ��rpW<s�>��_D�WQu�C���3�9�չ���ά]�g�0��l�45�� ug�?&������O��Wo�c�x+ۍ��ڲr�Ս�}x�qnTkhO5yS��4	L��>ܬ�ʵrP�g#�FX7y^9�mv�*�V'9u��,�%O^�q:c�mwe��δ֡�sg,,81Հ^(�ܞg���_>w
y�XA�NzX+���q�hjw�����6iy<g�G$�w�K��(>��^���˧7)k��R$pc/5߄9J�'�|��ۨ6��9���k|�oR�}N�(��^�6Q��Br�����*56�;҈b������R�2(�w
kBY�$�:�)�7`�J�]�e�D���u��U�j�>	���du͙���
jT"O�h��wzn'�z���}�[FC�Ό�۱��5�5:X���7�����M�ۡs��7��R&�yy��/ٓ��X1��nB�8TwTΥt�b����a6�����'��'2Pݞ�Sn��倃�W����=1��Ԗ)�E�Z��`F�޼�\�[��R�\a_1�t�^Jc|��ҡ0�e� �]�c݋�[p�Z�=8�{� ���٠�;�z!�~H��Ru>�P[#�uF'��`�4+{�>���h��}���)�s^s��(�
����bze���#z�W2��>}2}��j��4��ųkCtq8��09��R���/+��4�̸������*XsՑ%��t$�v��RrpW�<r���˵�)l(+z�{��Up/��g�r��YC9봕MZaEؑ�G(:�]�Qx�'R��'�2�6���*�&���7��R{b�W��ö{��ׄ���l�K�:c͔hI`��q�N/�a�6��/^&�ӿt�Ha�N�7�#��2a��g����4�@3�v��m�>�׬;���DҒpo�u���%p�Ճ���s��;�׫{��r��Κ;��s�J�$$�L׵��o�Ʌo,J��x�.��$�G�>�?��Խ�~�״}�w�����4%�m����O9+)��j:��ì�2�/]ÞW
^,�s�-,v1���Ó���/x��qmV��W�w���� _>'�2�����o��5ӷVx��[��O8�f��m4�A���c��*z�(wa���!#�&�[e�C�6Q���E����'�rfnq֓ ��y��J	b��n��k/xSҴ�Sk�mv�r�98�v���ORD�=�K�^�J�V)L������]IȨ�7-ŒN�a����~/��ӥ��(-�k��_Ԝ���K/6�v+����s��z����iι�I�<�}% �� ^X;Ԗ�2�j����G� v�B�k�V qz�<�m<�.6^��
��^�R��p86�s���8et�>�k ��$+���X�*f�KQ�";�bo�";h�����Mm�ٹ��S�}қ{e�{�qVeB�3f�rͫ�*��C54�*�p���V���xJS���zrI�lz�q)���8��2�e�s�yJ%ͮ�J��V�[KŃ��^�ޯ`]7�
�4��ͭn�ۙƖ�[��ۺ���z&�u�����	�pwh�5k��+-:��T�r���B��ѻ��{��jcۓ�l)�4:Tv�Bܚ���V�Ԓ�-F�Oq@��k*�x>°�o	i#_�%���0�2=�X5跉�bu�{}G^>�z�ޮ���-�e�'_��g�\30O3��fp8���)��,/Q���L{�K�.ν��X���G$�7lK�s5���p��U�D�iߥ������m�*z�k��1��w�n�aVDnEҪh<}i��2�]�����	l�B=|�Ў|�C��m�dcWOm���w�U]��|�J9��g}~.�9=ek�]N�v1A^b�)�=o�n6^�-+[mIZ�f�XIr�����\`��K���K�����[��b��a(�nKA�1fCl�p�!Rә(�_q�N��M��P�:�8�L��N���r�ug�ݺׂ^�聦��OR�Uz'7�m�P��e�EL�ܖ�����w���b����/�3�_a��-Syj݋0]��l��[���t�D�<����\��ዊ�p���a���	B�ߩN���yo�Jm'���oN���R#F��rV�֢	�z�"��#Y�cZ��J������k�>��N�|(29�ʾ�k���\p����}Al���n,���s�쾠�y�?=ک�YAonkF�2��0Bk��h����Al��C�J�^�|��_e<���G��V�NcS8�FT���>���@`N�a.��������{\̮=|�F��G�gB�sĥ��L-s��U����я6���GTŭ���u$�PM��4r��N
�z����57J���_��[?H�e�����-�M^5'�ͣ�(�6���	��8+��\�����˭�7�[\�ܲ��ˇO;ڳ.ioCՉ�<���N/e?Bw+Ľ����\�n�i���K�W�z�X^�<*%|�{+Uь�nɧc��m>m�K�w/('��͆YqIݜ����n����b�9ق)Q����e(�����w;9T��6��k{Yx�sӎw%�,�u��l��T�xu����
��6�6��d·��Vs�e֫ҵ)�����\��p.d������~�q�]��1�q��ۇ�𚺬�OMkgzVԣ�P���89�����/��mx�N��q���;���.�%�绕�u�KS�޳!͋��R�I��q^��t��q���<���K�N5˹B*ߧ�:ȕB�1#�CSi�Z���K�H��]��Vc���U��y���)+�P�����9���z8CU~�lM�o �w2k��� !���zc}��L%S��%�U'�/v�0�"$������O*ycq��%LݩL=:z��S#�!%�S6[ҭwfm�Ӽ��r�=˷��g%�r�eo���-��
B|��� �D��i�姱q�36�u�qz��MӚs��(���FKj��a�F`�l��U:���B�{7��Y3H�p;�GW*��Պ��@�ھ*��J�q��9�(Q��7��	@���m=�K��l8ąT�391qr;�5����dI�[�)�Ҷ�Xj�X�0�fJ�u���f�v�zM�O!��sa�7��QxGU'��[�R�]� ���oar�ZSq�������AIBD�Xs#�͂i>�����ϳrE�������SA$˿8c�7�''m�{xl�i�W�[�euT̻��v�Gne�-�e��x��*��؃��b6���M�y��@תs~�A���_o�|����{/^L�]V5���t��I=��P���)�'��ɚ�I���?_#�B�Sۘ��<}��9����	�>����}�߯>������y��͋{��*��³��'�,��&�z*?^���kB�X��--v1���XrN+5�{z����v:7^[�N~�&����h]^� �ƣ�;��u���c].j��8��PE��y��΋}�'�J��w��bM�Sn�7�b;"�q(���Yc�}��J<����d�����U0�����w~zZ���l�V3r��5=�ߙ����>ܻ0�؛��������>�Q���8.�9^�f:|-b4ơ�f��	���]�0r�k�NJP��a�s3�h]�A�w���ݧ��=�X�����M-���&�ț�@������Y�e��Y�%\��ug?Z��:8~����I|�L%�����Ğ����r<�3���Zɞ�<�^��8�G��v�C��l��m]u��E�̛+/}FoԷK�K�|r]�4�iZgKI�n[6�*ɥ~ٓ$x)/�|�;�ZVf���^K�s�ѱ�����%Pn�;��l�7�N�I��=xh��Uɥnn17/u]�C}���֬���c�I�dj�7+r��O;�r�sM�,U�[HOT���"��|rLwf���8�������7)N��Z����A��[���J#y�+��K�L������
�U���c��2�^��vy�Z��<����w}�z���u�L8�m��5�ɚ�O���3i	�K��Opt�OV"�:GO�I/�bc]�r⭠�Ԭ�r�E�LP�]�sഹ�3|(�v0��.�)nm�H}�x������|yT/x�6�ʻwғ�Z˼xn�>zU��[�pΙV]�	8�=���*-��A����u���0e���R#e`���`̨o%;����:��1�.6�-�P�-$��W�ʸD� o2��Y���e[}.={ �گ8�M
^K<�>4�Y�gb���,���M������k�ܖ6���*��O���Q �HP�J�y|)�9oK�z�ʃ��afQ�U��}-�)r��&LQ+(�����l[[����7��XA��=������R�lik���y\���"�Ή�QE�4TN���-;�,>1Lj�[��F��=h^ѹ�p+Sz��Q�z�j'6�W"rшl�b�?�\����sh[(�{3�u
�J��\�4�\�)c�N�iDvT�B��c�9+,h�S8[Dp�T����R`)�[xe��DJ�x$���}�݀|gN��o3�G,J�ӕ�J�m�2��W����R-c�m=8�
mX��U��p2�zen��MwR҈o�k��U=�w�ٴre;"6��6��[���	a������+�yrY�u(��%��Z;Tܰ����Et�+L���'�[�������^_e�\T���x�=�	�
i���oK�ʉ��L�Z��%�
�.*$�vھ��mM�b��I$:v=�X��6��-�����Sh�P��+�ޘf(�6��gZ7��՞�On&y�K�YN��ٳiS��53����)�P��n$��8�ځ���ޛ�s-�/v�6.rԆ��z���]8����R�ë�v��b���8�)�/{1r�Ȼ�����ۋ��oe���V^�0�49n�[�wnH�6��Y�.����f֞���6�f�`�%�ߜ�Ev�Ք�����S_pZ�� �Sn�n%9,��]*E7��b�N�lom�u�'w�P� 4�ۨvp�#j�y�wg1��u`Q�O6<s5�v6uɋ���}����M踝 i�4T�HR4�Wpiz�z{�������$��qJY����飴K�i5��gkX���H�AΣ���g�3w�z�\3K�޸�v�N7��w�!L�O��+F��mSc���}L�D"��Θ�+̾c�N}[N�F;ѸL1�	G\M��˵���"���<�6�Z��ݼ�LX,���El��[���щ�Um��\L�Ʒg�%�Q9[�-Q�z�m�n8��x;E�s%F��&AC�p��7vG:2k�k�`����Rz��I��(����r=��_=����O�(��|
WnV��Ni�r����qrhm��帑���[n�Z��VF=��漮�>��6�x���{nnEB�IID}R�UrC4�-=DTKVq�d�ܬ����}IMģ衼����j]ݷ�'���z	��$�Y��b�Aej��b�
�IQJ�E+d��,D��e`� �(��,Y*�ek��V)�PR�V,U�Ȩ�XV,�Е%a(��D��*�IRAaZ(�m�k+YT"�`,��E�VV,��+-���
�$�F(�����
b�`��"��B�)R��%H�����XT
�QB[A@����EPXT�VR*[R�!PX�BU`T�Zµ�~�%�?|�ٷ'��2�1�=���E� ��A9�zr�5�+�j��N�A�׋s��5��%;-��nt�y�*G�aW�t\Jڣo�㛐OW��G_uʳ��]=[+m*z�k��1��1���j�q��a��ְ��C����
�^A�q�	��	U�#���vĎ�^���ul���}�V�uYኬ��K��Ps��
b|kf�>X�]p��f�Sr�[}`.�&�3���[%;2�;�$-����C�[�m1_L+���-'�v��j�V)�O��:nh���;|�7�=L���-ݲ����ϋܿ=)���ޜ=�$J���{WMU�ǯ��I�Y��G<.L�.<k����t�}Nz墄D]z^�Gm�&ξ{�M��{Tƈ�hH;Ϯ���{@�]أ�{��۰�����<���R����KD:��!%c� ��k�!�-Lǹ��*�̇_�'��3��q�Լ��q�Q�))Q ��@Jܬ	��%��DK�YCvt��6�dLMWY������%ޓ�>r�=}M)�ƒ�jƝy�J%���)U��Y,.�p�����IC����y�|���
'����]z�e�,�>�wi�.���M�C׺/1�4���,��	 ��1n>.��weNj�rZ�:�ԗF����R�����>ro<��*-΁�R7\�5��ܙֶٺ�ջ��!3L����]�)s0�lsF��������r2�����+��
l�	]�쵕�X�w:��QM�dsBF�9S���Y�w�P﫞��|=�%�}�K��5f\���}x�qB�(�ӷ�L�Vɶ||h����_W�V䀺���B��%Y�����Q�X���$b�CĽ!��������G�h��'��YA+���7;^�g�؅��[le�WGa\�tP��`FO;��Mޡ���<��I�toP�:��ݞ{�ݜo`��~�/C;�2�.���m�o�l_�����u��޿^v�yc�P9#ؓ������_���EҧwE����_�s���}%z�{��765Q"cc��膖ҕX�wa�k/RI�<z�n�%6�?f:|?\k��M-��7�t�Ql6QA����4+��p�R��<�Wm��>��ro0��-@�hVT����[�*��۱�K1^vW%�(>�er2�f��5A8��x��S�q���ל������g���v��OZ�\��9]�;�{���>W0�	��t�W���/w����-�8K�z��o5�B���u}�i����(-�#3�tʿU�]��"�s[���\ҍ�]Wo��py3��惝�i�^~H����>���7�"A���+m����~W��	�a��Y���.2ZQ�%*h4:�C�v���c��K��0>�}��5~p���T����FÝ���K+	�Q��{� F�ۯ��W�s��N���,F��#.���ͻ:d)ۃ
�\sVes�|2��X��Z��]�%SV�Q��M��wu��דa��Ǣk0iT>���ʾ�G���~|���V���AS��]��[�8�n�Pm	�4rgY���s$V��Y�X3c���}p��[��Q���O����ߊ�����w��jx,Ғ�*�jN�(��p�['sǧ$[p���jLC����}�'�(�ή���j���U���vs��}!����>�C���8�
ƕ�pb-ff^��M�`�}Q��*�T�h����s�b:�pξrj"観��mSV!��\A��X\j\�}��[��ߓ�;���Nn�7;ic�6uY����x�Z6�d���'\IA�V���9�@��6��
[e��m��V�����O�7�[毜̪YY��y��ع<v1WX�v$ܪm�JH�Q㸮ջ�|��3�g�w:�d�.;)��ب$��/생�U�����`�٦�S+k{I:��9`.��xؚt��BC߹���K���9.����]�u+�a���� |^��R�Y}�ޝ<��ƈ����3\6oF�R��w˘@�?LsR��T�0%���Ӛ�i�.��͞�ٜ�f���m.��V�Y�Z�t�c�nZL޼��m<�4�i��n
�Or��%loLX������kf����.�}��ri_�>.�q��lDG�iLRn�UZĉR���ڌQ)iV��Jܡ��wB���~x/Uԕ��߲C�P�6]q.!��h�3�*��Rdq�0oWW�ڥ �c��.�ڌh]P�e������ߖ�W�x:h��S�=,�X v4+�Y��'���eX�̜|��`C0�G:������zmsT�/h��U�s]8�y�g:�je���`�u�$r���*-��x�H��5)�e��S��#�9���^�OT�L�y6'�&u��C�9B_h;e�Y�Y��S"�R�KK�TӻY�6�o:��qV�2Bu�ɚ�I��)�u�lg(S�a��%���.igt��bc]��Njz`bޫ����nn��9Te��hɎ��.�V!�z�GJ��T���zS�<�i*}�-�:��l
9�jx���/�f��;�.�gA�==
�p��8J��5oW�Nbk����m���g��%.�-��d���C�P���ph��j����#C�^kS-��_�\��<�/��}�~�&>p���p��]S��b,+�&�zN�z�&�R�8^�������o��2o<�3�u	�J�J����|^凥Ki;=��b�u_��@
�N����!.[�P&���QT��#r�¦��j��;�٫JM��;����dశ��9�c��b;�֜V7ַo�/U��ڤ�8�e����p��<�Ε�o�7[(�W�~Wݸ���S��ͨ2�R-M�u'7���^�eA׳p���ܒs� �2�P{��K+�Rx�=��>�醦�v���/5NS��3��e�^J@�␟���dv=�U���{���1�ʷ.i�ΧZ�qL-��Sԭ=�?7 �K� �}}��O	�̨}�7/�zu�Sբf����x��n�ۙ�j0BPR�6 )�����w(��i�Ǎ������Y�>���{ܳ����eE��W#�L�Y%,9ǣ-�ԫyg`ɹ~�̡���j�^]�4�fc�C\�����npW�4�sQ�����	�����L�w���ק���_A��;�r��Vq��k�󼂙�꤃�=�%��H�3O�#���g��lUS�{,*�׍�*&��յ�d҇�JJ�������2a[�g+�H��y�(����[<��a�{��Mˋo/|�l�Y���D��O3�V����x�;a�-X����yɃ���fc�ܨ*tG]���M�X��H��I��*E
W:S�>���03ra��t�y�:�d�SE�B�o�Ƣ�����H�JmKًE������N�۴al[�NY\�_\F��ΪΜ\�a��5��w�C���~��my<g�A`\t[���iY�����Nt���X��b�s�p�+��ޥ��g�"D;A�*z����^t}�ްVz��b��z1Wy�5�]*wq�=��^��7�=�M����i(��< �;u��^�2ҕF ����c���X��y�c9�98�s����ԑ*|#D�
P{���)N�V���VE�S�e��N�a1��}�A>�a��Լ���2
=%�Jg ��ZQ���\�iB���M��)nU��s�h�7Hb���u�c2l������z��|j��Ɯ^����Ӛs��(�
���x�ޒ���F���{�U�n75W�U𧻓5n~q��7�9�B23	���\�������/T#1�h�y:]��w��uۭ?���Ҽ}��)$�9�]=]lR�L���.�n�Z��=�ч��w<0d�f���ݬ�J�?�n�Pr�{�A��eIw�2g.�R�{K���/�U��w$b�A3Z�����Sh5G#�j�8�(ZzQ�ޘ3
v��g�3�nV��x�N�����X}��}��U�_���d^ͩ~������G����]ݸ/�<b��[�g�&���Ѓ]~]���zpPn:�ihʸO2<�Y��S��J�]�75?=���qB�8�6�o�ZN��W�{_��Q��F$�Yޝ-o9��䵝�1��_t�ֻ)��7�߳��8[[��l�3zq��P];���#��+�"y�K������㧕�R�g����輞>����J�K�g%�/�ݍբnv����!|��s�b��;��<��46�
Y��G5(�v�[�Vz|+��^�=C҇u�t/��ě�ño'�YV�`���m�%k�f��2k��YZHٰ�,R栓�Noa�{v�����y��c
�~�-�m��?�z�-�!!��])9����}�2z�i�S��R����[�}j�x�x}���v�<�����5댔�d/!.��k��x't 8l"͉D��x)U�^*Q�y˞��j�J����g�l�x���i�4�G�;��e��7���ĉ�[#WݏJ��JF���1��eS�l�s�]ħ�]���Y�ڱ~��#P��a��"{sc9n#~��&5+���T�1-}���4�i_�gK��I�,ᦪ�v�޳��:
BN��ϻ�ZV�5�'�O)̮��ɕ]�{S�$kZ�+����y/f�{0��.�}��riXp����E�ݧsr+2�g��V�=��3�k�
U��oU���3ӬcjV�[�}yn�-��=|�E�h���8�Aj�v�Bܚ�D�u��^WY��]1S7]��hZL�&ā�:��9�~顟m�z�ϡ��{ߓ��Z�}�^�}y�X�o}]c+��2����g��ڪ99XRپmb�6���D.̿	Vs9�M.�t��bc]�-��]���uŶ��Mj�5s�ۧ>�s
�Ш����g>����!"�;{�e�n7����4��˲��6r��WE�+ն*qw�y�t�Qٜ3oD�4SF�ת� �8�a/�r��W$C��]��3��+���M��J�:2����%7i��Q�ƺ��%ʇp�e�Y�M�,�{�N�0[י|�����ŴDŀ�$�`t�Ck�;�=.T�ά�w�Vܶ�V�l�e�[�f�1��e���+���~ƺvh�����O>�9��}�g/L��޳��$ri��M��cKU���WuBt߅��9�%���Rqr~�C.4fZ�x���n�4���ֵt���~�iyT�����M4��/�Z�%*���yi�M���{�+�LlL�s5�3��k��Lm	P�v�1��
K(�OǺ��D��Y�ĵU���S/1�zp�~H�w�_�-���*]݌i�-�2z,`KV�V�}�%���R���t���K��dU�|qFZ�U�::b�1sqz�9z�=�3��`�JJTF��YyO�a�wm�������
��[ [�\��kJF��G�gB�s^�)dV�R�֟c��	�T������P]�4L�&�4o=�N `�^��L�c�n6�1%.�7�RV�N�-)�qc���6��+�g$�NW+oA�s��)S�K�0��T+�"��d���Ʈ�.�I�� �뛘;�[�"�uգg1��Y1#l=��3){1a�)5|�k�v�^�U7t��,:����~��,ԑ[�/B�������7}D���w)��^�[�Q?�B��o��o��+[��m���h�9;��@$fԻ]ԻuP7�}	�!�o�4(��+YK��ov��g'H�fQ���B�v��ڭ�12��6`�m��S~(��Gj0�U�I,��430k"Q�o�Rʨ;o����)p���^oo38m�B�[�`�
��k�csL���e���� m�Nu��r�ɯl��Աq��w�*f���jj��|nR�f,w�iZ�#8�չ��<{o����1�LJ���c�@q���X��!iベ����Gݮ�u�}ѩp&��$�v�3T,\(l�H���O���k70a1f5)]ew'RD�D�c��@"����,�����iʰ_;}�֯�9�~�)�`e���Qۣ��;T �f�=Atʺ�Xx46�]Ӿ����iE�;)���c��I�ǐC����+��);���q&\��N�f�[;Mj/ G�^�$v��]��)Y��]�q�M���]tVu9��#{z@X���f�K|�KW��;�f�t�4C�~ռ�B�8r;j�%��7n�d�j1���sK�7uh�V�b�)�=p�Z5��3��:���!tc��V�{��]r���T"��U�ήI�Y��VY���\��'y|lj�OL)�D�������dy�k���{��UfA��޾�J�핛p��m6 �x�(Et�P�}��f���#���gz��Q�c�b�ҷsU*�ܮ�Tz�e "{i�.�h�_=��v�s��Sn��o�^m<U�-VM#�*L�lQ�� ROw�ZIۃ{���2�E����/k�i���̩k�U���],vQ+�L��&Mv�mel�w���[27G���g	��u���v��U���g�v����O�lw���g�.���wwM#*@��u�\�p*U�qכ!�7���ㇹ*��u��ڸ]r�
�+<eQ�+6FoV�2>��8��7u�e�^� bSgG�)ڦ�h!�����aÁ�k�%�uZ�*����Qj�é΍��ο&{9��L����EtԪ����3w�3�!�4��ң���U\v�e�DݨR��>HRi��-�i�#`�=Qe�l�Α�kpN���W�~��||-kƵ%�L�%�i�S�z�5���i۰�M��ͽ�j�m��L�\Nܐ��E[G�&�Wf���f�|E�\��8�� ���A�dm�$8����fV���GK�c��l�oqi����t+$A8L����=Ľ!�OO\����Ԏ�Y�O�#��@$��b�D( ��P���R�X-� P�ed+�"���%A�*��)P��DQ-�������J�Z²,R�V�J"*���aY"�UeAdU�XE��
�$�
� ��[aR
(�d�*Ȱ�TX(XEd��Y"�Ȍ"�
��@m$R�m��j,PXT+XV�YR�d�-���F�@()"�U���(�*�j,�k
�([J�ءPY+����IZֱITKE��F,+X[J0+RT�F(Q%��b¥IZ�k
ֲ-�U��R�eJ�E%k�v���B�.֋�@��AZ���-��a�襭Ave�D��P���Q���cZ-�}.��1�pS�O���r0�������{A���#U-���3��:��QM�eD8��ě8�T��1}GP5��Β__y%/�F��U��1}�-��r_�o`�=�кͅ=��ij������!C�B��Al���0��}�~�VM�p��O^�\P��,7�9}�*�����3ӏ,W+��d�EA�x#׫���R�&�Pՙ^��v������9N���j��iv.�������X�|�B���{~m�o�{c�F�1l��]�V���+n������C�FD���Z���"�V�:�����15a���jQ���.��e9b�wU�zԪ�����F�GV�\�o3�w1�s�z�4�v$&��ߩIt���U�]]�qS��7բ���\^�0��tד�v�����R#D�����"^���Ү�q�:ةYSA���-^��	na�Uk����'^�g2�T��U�Cw�GFo���hVh�T�&8��i� j��_l��}V�q�����;�2�vSr��K��1Д�̝o�w��0u�y��f�}$o,�:d%���'Z�������}�ٶ�4�$�C~�P4�A�wJ3E�8���y���P��������4���Y��+�Ӛs��(��s�L��֢#�w��r�`�J�0�y�W��.\�p���q����T�;7quiS[%���V	V2Yۥ7�G��N��6�n�~�q�$S�UO	�x��I{[��;���nw��ԋ�0�	�Xd,��d2]W�sy�����r{��uCA�d��@�N�9`�W�l��Xh�]�L�e,��;o��^�g����y~�4�3��(��������&��Aɑ��� ͗�q����8î��d�_S�m��H�0��}3/l<���E�?>63ꯌ�]✰�����z�l��1��&��A2�s�lT�FةEDm�d�{a`�V�J�dY�VE�I{˃�Ho���^���qG3U�0�,K,�	���"%�Z��O�jY,2-:�����Z4c72��T�6#՞� +RVi�A[�{��b��=���`�q�'��o��	���ڑ�L�y91���/e;������֕B�R;��i��' ��i�S���������Q.�(*��]��U�檾�}�e��6G�8����' R�L���6�`�ù�����B�����]%PKt~lS\�oخ�xc�33ژ��mE��v�1�`w)��9n�� �:xߓ}tz�0�#V�؞�\ׅ��r�z$Û�����X������W��G1�mj�̀��3	8�J�*���]^qo��Փ��ח7���k���bϼ�4�r|�r�@���z[#��)�$��Xȟ�z��uٙO���4�O<E;hRS��J����(q�S�"+��v*�mځ�Q�XACtK�ʫ��풖$G�����>���:ם�=����͖w���Ì"�:�\�-���	�Ep��{PkTO�"N�)��Ta�`B4�}�i�]��zo��v���t��8�g[Wl��[��N�^�*JO�֞�b��2НR�:�8���[Yu �n:�שpSWc�������]8nu��=��κeҘS�ΚƿU�CR���Dڹë+��h"���$��/�8��2N��5�^�d�^r�^g�����\�s�d6f�ɟ]� �;8�`�Wi���>����]�ns�}R�����QT����Q����a�L@=y�D�j��7M<V,q��Ξ��a����n�-4Ч�ne9�ObɎTY/
T���z�`;6h0K��f��oi�Iδ͌cՅlnE|�&�,���w}�R�s@`�mQ5��6*�[�Rmt���:��ۻamz��g�����+Aob�f�A���%
?GC�8Vr�z��X'�rRi_)����
{=cƚ�i�+�G�V)L>(�|�=6�7X4�]���F�8Ϸ�C�;=����0!��;���Ū����c���x����ʳ}��W�>�W�S��B��E{+b��w�&�����ק ֕��9��(��s���k�V�0m���z&��vP+ՑCA��&@�t�:�n�5��]K�����Z	*����=��'�y��u6�����G
B5`����n,j��B<���n!�!�][сtȬ������՘������uvQB&K=,���h	�қ(�X��9�T8�HG�Jøu���ͺ��m��[���KR��H�ZM�m#k�EI|�i,���9��)Sژ���Rղ�����V��E�v8�Ӷ�{�D,*P(BM��<!��zG%E��52��)w�x��hT�5���U��u,�,,N�1��*gQ���{�Q�zw^8�=��)W6���ʚ2U��a�2mh���^=sJʁ쫒s�w{��2fp9P��Q@�M��s��U8`��O��E��nJ���<V���FA�B{�9���٤�ꖇ�5�Ӽ۶hٝ�F���2Ao|d(�:��Ï���F�<�;݋>U�ūGW'iF3�でt��U���^S┒N�r˘"���y:MC�}u5n�C;��y�J���CfF8�F�m�o�V�P���Ѯ��[��j� ��v�1��~�}l�[�"��&���1i��f�ɛ�P�G_r�Hj�'��^�au*���#2�,���m�%�p�9wo��s�ak���r)�إ�_]�X�]���a�i�q�@'�셶�"@�J�q��ߖV���zHޜ^#3x��o�8������"([�8���O5y�k��
��Vb
!�h"y,�&�{錔^\����<TЫ6�Y��#�|��g��>���<��T^��F׌iYt��<�[N�k3������#������zT�fʘgbol.�6iCʠϊ�s��D{�ܙ��b^�	3�u֟���"��>J*"dr6�n�9�Kr�7xY�q\'w�6v�b��[�a8\6��
{�^���㋦0��le��<S�BE�{v�E�H�9�g�z�����W��:�N'<�(3�5������%'�:F�ືRc��
ކԤ��o�7T�N:�Z�􋬞i��/�s.��p�zdqN���^����`�l��]W&}r�
��@�HP��'Mås¬�^�,�ӎ4sYv-�ú���F$���j���Kt�|;�tb�����1��>3�.��=$���	��g%�:C7�Q%,CA<�J(C���}��$W��]6^��WuPe�8q9��,c�Uy�,ѹ��ベ��?	4*),ܯZʒ�zg73'+v�{�@��uG)�*�()�q���v�IaƚQi��nI$)�Yâ\t��ї��R�`��6
���z��\�l�:�S�����ˍ۱V�]�v"��[��Z���$��e�-�� tt<)C��i��J1��Rq#�fÙ���0v�3z��D���z�Ϻ�X��FM5�V)Cƍ�B����뒯�GTIJÃϲ������،~q O�F�XNj6�{n�#�ہR���N2��XU1�ؔ�`�<3Z޾�B/U�ਞ�&������h�ِв:����̲y�Y��#�*DJ�4 (�X\ٖ�[X�fW���>�'��8+x��f�:�Qv*�i"��I��,ҵ6{���8f-�ǙT�8p}l��A�f�kj�{]�(���c����x���]����7�u���g�ˬÄ���MW���ٌy�,<V��W��ȱ��.lK4Y��&��Aʡ��zkǚŴÛ׶�[�;���.E�o)ʑda���(f^�X>�?t[s�#�y�W�lCQ�	�7����uWo�c�Ld�qR�@�����2ctT��6����G���@�1.1F戗�;�I�Z����)�.���CO�Ĳ��,d*�͚غR\v�&ԍ#���X���o�6{�*������0x�������4�G,�������V)�^��Hi^����dv��\��s�=�Mڹ;�fH֤`�,�n�����~M��y��B���ؔW5���Oޠ�r��y;z�A�[�:o؃����9����t��Lyl��ԝ�P�@dԸu�1�_n�O���͘���TV��Ly
4<���r��+��A��8=3�9�ə�7����\���)bZO8���r�$�U�Xg�\L�}%�-��ޝb����w�)��.�{5�z8ʓb��4��2XTN��H�>�Ӡ���z^:v�8c6Y� �б�����z��!�s[b�G��DԾ5�}�o�s�{L+�!��q�B�j��;:�҆��X1�wub�R�Dޢ��bYJ�MX��nR\�K�P}�g{%=O� �7Eஉt;�U�k����FJ[3��g[���"��.T�đqh�G�a��Қq۽����݋'\�O��� 	9���mQ���F�����T`��.��KK*�5W_�U8���8U��?x��B/
�P����)�=J��6�t�Umyw*�������
﫦1�ȯ6�<)�^��	�E���R��}�Pݍ�;nJ�o�ُ��TsHܺ ��+ir��RBv�R��h',���D\�:�9�[��W Ჟ��uO�eK�qb۞W�~jF�Μ!^���1d"�&8^*�]�.eb�2�G삝�Wk�&���r��+�a���h�g�s��C����'s��OoU�vb[Z�L҉aJ �T,�8<O�W�B�.��>)r�ܷ�*�飁��eh(4���W]���&���$,S�Q%m����E�I��	�p8���;�Ta%x\�/k\u��%�����N���b��y����ֺ1��{�P?��Z�����Z8|伾x�����0s���7�q&�r�.�t-N�m�����F���]P�*gr�NY���Ǩ�"��5��}>�˙1׽O}�P�^���ݫLi��ۑ#k���j)_e�?uv����u�*��om9���7}�㇑�f��r��G@� c��u���9���s��]�y|(%����1m�:�	�Uꧻ�G�M��������)��:�a󰝆�"x����-�g�卢�J�ޝ��bX��pA�*t����S$q��қ(�U�2߻o�WΞM�C޹��E9ڞ��cF!�p�5I	i4SiДo�g��RY��U	�[�3v,qq���Oh��:��C6����Pd_���p�#Gdz6y�e��N;,9ux����W����Zv�w�	`=�f���E8�8~pAn�d��=Rkp��^k��w0�8ŉk�!W'iF3�で7n��V�8c ���|R���x;�/-vݩ�k�&������D5���r�R�\�i�p��g N�GZ7�YG6�U���֓�>̬_C�<Z>�b��;�o�"�u	5�8���r�����v;�=n�M��hg�#	����O�6t�ХW�.��ʇu��	/���o(Pka$w���Z��/}�6�*��<��Z��K���Fr�^�1p4̇N�V��Y�z���h"��YW�|��MDs����X�F�5IS�tގ˥-��͞��n,�\Ԅm�e��J�3����W�Y�Dq��5^��L��()d����<���҂��v9��hToe�a���O�SwJ�.k��]:�H��}���%g.�3b�i���n��L�}3s���%�
�����R�5�XHE����ڮb�.�Wv��51�]�Cr�2:!�hJ�{�wG�m��Cy[Q���Wc�����-B�d���!d9���tGX� c�Ϭ<�4�T�8�7�9t��BԽ�{�n6˯>�j{6��qK�||�\�����3�]�^("�}��J�!u��˯��{U��m�cK��^+>KA��T�L�D��}�<��6����絕� �6�nH+cK6�kZ���+��������$D9UNY���x����=���S�x��'>离�`\LU�.�%�ӄ2�$`h7�+�ͫWWP���Z�S8
����l�t�ja���:<�]���Vx%>#A�w��ĭ�����z_E�Ik�IX�X�q�)�q����O	4�M(���.���&k����>ɶ�$����v�V�S�Li���S�E�uV�gL�E��ج�4��n�,W���]�v,pfP7y�7SlpO~Y��(��}���T�Y��:�c=�&�I)�6vP3���L�\��WSt�o`�z:��azZ�ht�%�7�Vj�1Mٶsl��u��w��6<=H��W�gc�������Ńk�D�DV\"m���<��<4��ӨT�ْ4��m�ƍ�p��L�qvd�e�v��AEEw�ѥ���N_�Т�6�kdo �Q�lWy����0�Cn��\��I���t��
��W3|oU��]	t�x��A	�M����k��b�R�*�.��*� {�E�ղ�����ޜ���:R]i�l��7��;���)�ve񿈄�J��料�h�Yם�_>�n�M�`x�K�6�:�^pӼO�o�8P
�L.0c+M�%5��;�m&����W��d�)�,M�3��ϦOC�zc�u��5�hc�L�͡�#���ź�?N�5�H%a�O��ڶqvK6�r��E��k��L�-[��ef�o�!XUiQZ7��UʮV�.�!nK��uBX�{i]X�!�Ie�љ]}�h�*vYխ$VKT�R����y�����[�͕9�P�<�˅w2.�+zF�r���y�ʰj�M����Ҳ	.�{O���h��28�u�KK�1���`�����-e���|e�o'�a�LY�v��K�%UV��t��Hc�yH`�ml�;H<�F%L���n�:3~��%�,t��P�uL1=�}�\3��^�i�[ƴ�/Y���+��huX��S�h�Z����x�U��A����eoZe�J���)1C��h3�ol.�]���|yk��i��F��|G��U/4f�n4)SA��;r����Á��Ǚ�^M,��n�BFӧ���=Zi�b���pVU�`3X�m��뤨���!����ԉ��FF�{!��ߺ�����\�z�[�`��^CV�FA������ϱ!�����^�R	�Ĥʝéq�=��:j�G�WX� Àh����;�r��i���gq�d�-IC��=ٝl��_��-��j��>p�[ֳL&�;}z��n�;�����P����]��axKY���9��ʹ�fjlS�D��6���y!x5����`ᛥ?R�ۧZ�m�̆����P+��]�0��5�V�,*�	Zؼ�����w$<2��Ԑ׫�TUD���Y���y
�\<{9+|�<�f��M������qK���ʴ�D&ݤ� �Y�jch%)7�f�[��	���Օ���tz��֧�ä��!b��f�q��\�HD�>��;�OžnƠ��tj�q�S5u�x�����u��&]/w�u�� E9�>Y]լ
��f�iޏ���ș�F����oN���*G�S����ܰ����Z�m�	Cdf��޻�Ej��-�C!�3�+t��1���S���E�N�-�*�o����)�_]�ղ.u��� ���N/�b¥�n�Wv�	��}mI�m������6�QA`�TX�Y*F��#j���`�*T*�T�)lQKj�,X�+E�j�+dQ�B�[j��mX((6��!X�!P�Ņe`��� �ѥ"�m�2�(�V��k-*���[mZTV�Q��������jZ��"ū-����ejª�-T�6��[j�e`�[j���D�m�ZE�U� �F��
�(´J��)Zʕ��4��jJ�6�Z�iFګ-*+��V ��c[m,@����l*�(1B�F��AKZ+P**m�aF�J�QaP(��Q���J�[aXV��-kQ*�m�UJ�Uh�V�)m�4Z�,�����|ן�:��~;�Ɉ����1$�w4�Tr�S�j�����W"W;�$+bz�G`�j��j:�9�Psw,��]�"x���3�20���L��ڰ��[�FO$/�|�#��=��Ҍ��~�3�G3�]�����ܺ[ǭDe�?>�CR����E�����J4lU�1z�II��,<"�}U�6%p�XY/���
����֠|�}֡D=+|��C�)�4��έ*��ב�ǈ����ߚUu�ܲw�����ϳ$GJ�W��7������u�,�z&�`Tq���(urs�#���.nY�̶���9&El37�HE��٘��7�J�!�j�5�YH�
�da��72��� ���|g����%�ˊx+*ܪ�+Xƹv��W�2{ d\������2cv���݀3�Ol,��[�e*�p�/�����N�I�ےȌU�+�Z%����d����\�(kb�Iqײ�����k7ۢ�x��&�zC��i��3goͻ��O���B[5Z����J%�)����݃�jqR�Q��u#�:�A5�=������˺��
�K>��˴	�dF�Ok��O$Zī	�{��(���m:rT�|������jfw����n��^^ԇ������{N�� �l�Ÿ��x4�^��eߨi�*W[~ٌW>N ��y�*��m�|s��\�5<,��*���η�j'Z�>�:���7tE�/w��1 ���`uM�r,��f�u���m�3��>�:�5X�7b�3bm�������b&��8ESL�8r�e�o>j�Ds *�s^��r�g��^t�r�Η!��W�c~t�?3O1��O*�=sVG<��q ,�-Z)
�r�M-�+����%q3�$�ŵ�#�/��p^v>�yf޷;iq*�S�ӻq����"��R0Nل��=Ϧϑ��c�/�l��S;��&������,�ge!Ｓ¦��n�
tT�D��'g�9��X�B<o���o�����a���K�^�D�R�S�8gu��uVr���׾�������*�Z�y�B�zOf=͗��܇���`+�����d�5pד����Sc�L53Z��#9z	=�u����gMᦷ*�#��/w��I.�A�NH���K�i=�b/��&�P);=�/Ӡ���I�?�1�PB�ӚK�f��5�8B��wў�,K��D��3G{4�����aSH�e�8[��ѡQ����o�yz͋��rV-�n
��^�����79��$��ʯ^�
�Yu����Z3F�d���YԔ�����T��t=#ç���pq��|��,�l��'��U�֤�M=;ͪ[R+�a�%	����^^��i�����Y�,{�
�=�}���I�$��㑮z�������%�0�|����];EL�<��KE����s����T ��5��HP8G0��=g¢��o��<�<m���m�qֻ���ㅉڡ��r���h���xP�4�k�|+�k���Pr��W2��a��۱�6��7��5��޼uU�Y��y����]Tu��U�cH��Q�++qv��d��7�&C�5�ŭ�L����3ܩ8u��2[�"�$ϼ3�ݭ��S���]�l�����4R\���U�X�V�Ȭd����4#G��;�8D>�T"s�s�Y���JH�뢳�P����o����8צJl�%V,x��U8�W`��8��Ӛ[�ޔH�=���(o/v�Ԛ��$� ��@��6��^���x\���n���?N���s]k�7o��0�أj8��}A�oN�8d��z$p�gѳ�;=mr�Ide�u��F���i��}��^��uǬ=�f���GS�C�pAn��v&���u-ѽ����繯��KA�P��P{�BZ9;J3�g:da���w���3�b$@I4/)��������Ae�2�(��r�v�U����s��u���$أh��g$��8H�b�u��p�v�v���=�N�Bmо�����T�km�-�9m�l]�ݮ9��S-l`V���䭙������M>ފº��!u�zN�7�.��]W|�.�/m���f�8��49c�w.it�cyz+#)�`~�x����w0��'��3*�w1��yg�G�lo�%l_��Iu	4��&
���{��e�76���^��4���0���ۡx: T�m����2��pɛ&��w��`����ީ:�b�Eg�ϜE���X5�j�`������R��iY�o��i�?a�r�Gl㍺�j�S͎&��E\3iӾ85:$Eu���t�M��f獵�c+v
�CT�
6���ڧ4皫k9#�`nC#.#+(>�ʐ���b���<����W��ϧ�o�6M��P��4�S�SRM�v�
��)ZE��6)H��+ϟ�g�$3G�j3ɽ���i�SX�O1�O���u���)-��U�ˣk�	it�'�@sV1@k��@���?�U�²҈׍n����q�~FzX�ݲ�<usW��$�!���T��rf|�Z����](K	��c�m��*���	mC|;|�uB2-k�uq�>g�*����"�_�-�)����ߔ�Ok�/�W=�\@�[�9��`o2�:�b�}�<g#y�5���/����E�V��m��:����ًt7��+����V��ܡM��(��,ef�� 쭾��t�Bs�I�;u� ��nf:,R��_t�Vq�Z�M&��Gt��<�%[|ㅄ�T�<C�S�[�-Fd2TKj�a)ҊN�͈�JXT4s�TwD�痥7ݙKR($�F��-��!]3�<����IN8�>�g�q���+h�Ά���'�֝�@�*_E��#N�b�+V8�S8�wCv#b�:lr�q8�]���L��+{C��-���)��C���zX6VΧ��cV2;dyN�%�$\�y]eYO�ޛGϞk�x�*hUʪ!�I�L�$ C�B�C��i�ZQ����8����]C���(iXs9�mY�����բ��<k|���G�x�/�W��S�3^�}%02GTImK�iā#�42Ӛ��o���E��$��rk�ՋF1�˪�ܼ�e����b,�����J���S��i�d�:�u�����3��W��E�rSw�*���ZY��+�����9K����\ߥ�,�6������E-�#.m�qڝc�a�m��gi�Km�˦�
���+��C���?>7�U|e�2d�P�}]Hu��j'X��M�R�J9r���^��$ȕ�]nez�����]���h�*�
]�񝴲��uu�E���Q�)��yl�m�O�5x;��.V���{�� (��bYwv�g-��-u��)>��n�� �S��Ft|�
-�qa��"ʴ�`�a�Yk|Z<Na������Z��"�{��� �/m�u%Gr9C�SDZS�7�0�(�6�Z���^Β�����/6�)u���=�����qs��g��6�f��۾<sϧ�lz���+�fv����ro�ɀvw��Z�.��+�L.	�-���.hKw��t�M�QڀH`�#Gз��coxtsr�o}jR�T1Uo؃����
9x�7`������u�'a�:���yk�m��7�ɭ�u�R�k���E8���"�.��Ÿ�>�p7�����	&�n�����G�#*n�t֕��1D�>(2IC>��:��^� ���IC��e�
�E%�&�#v���q?<ݱ~��{�}:�H������T���|��pq{X��m�Ә��Hzi��y��&r͗�bܳ��4�Y@:۷<�i�3��\��@�@�3���C����m���.��.VG��*j��҈y胅Swl���q��8)�#	p2	�G��g�C�����Y�󲨪`6��L�w�����0��sk����m_ry,�8jVgt�H�F�,�=LT�%�Qd�.g\tR֤峔y�J�W��]8�.��>�]���y&رk���ZC}\��]&�]E}��n����ܛc�.���2���{H3��ۮ0��)�^�A�@'T�κ˃�hӷΏdq�l����:�R���Ԅr�]F���WuBq��� {����<���Yd͙����Dt���y��vl��ӚJ�f�(aƼD�5������(�����o�N-^x+�T3 �I��v������h[�Q��6-�r}�G�ۂ�����V��3*>k4�����|��P�S�x�^j�#�Y�)���J�Y�
�,Fj�5�w'Y�j���]P�~JC�9�h����:sc6$� ��P��ЉUiC�R�^�>D-�~��hd"f��D�t�C��������?wl���.2����4���}�B(��B2�j�@y�߱I�ܩ8u��3B�#04�{f���u��{�r���Z����J�T0$��HwE�J+ئ�jA���~N�q�UV��M�|�4��U�Js�A�#X8�Z�ΤVh��I�z�����H4��FJ�X���5�qWYgNC�q)��1�m�N����D�c�T
�#��l6~VI48F���+�:d���{�]����ߍ*f)�+�2�.�D�^T�d�
�u�ʽ�F��,��/o.h�pU���<�f��3��v��]�%ٝ{�Q��g	3��u�aS�E���i�:O����RĚ���8H;�C���L��;��]���9\ttϙ��q��h�j�b�������ӵ ��$p�I��ŴH����֭sۍ~�!�x�H*�_�^�目=a��4l=R�����gt��>�!��sڳ����b��k���`�0�(M��?D��zE�3��p4�ݻӎ�m�j��Ղ�I�ݭ�#��+=SpHW;�I8�J�Պ�ѷ�Hf�bB�r��(7/�y�qF��q���O����D"��VlE�x<��vP���<\k�pd=f�� ���I~����[[+hnV=V�"�x>�kb&;c�m�Co�H�k�au�܆j�������9v�g9���k�9������p�)�t�(�9��
��x���|���	�#嘞O���v�5�Y�ƶ{Fe/�9`e
�f���NIN|�.�K�nY��qoE�S<��ɶ;*5-���<������M��w�!8�ˠ���bҺg�����[y~���Nvn\D���������ŋ�����wuL�Ik6�VЋ�:���[M��j�ג�<�_��T�f�|0�G���3{�)��;�}�ʴ���d}��'��Q��X�n S��↜{��۽�ea=�^�9��*[�놎��SVAM��wga�U���߷�o.s� �x��\skH��6)w$�'����Ćh�E����
�R��^�b���uے2�0�k6�{谬V���U���?�9���b _:�1��6�Ww�CyU����!w���۰���[�Du���~��tJ|��vW��7T��I����~ΏXCh!�)���ܗuB�k^�\Er�	ϋ����!�UM�ݍ�c�z{o�^s�&d��}tEb���ޙj3�b���p�/L#N�D���h }���q:�z�?5��S��W�cʕ,�z��/�L=�x�Nx�A>�az�|�<�mf�������t=�J��ED���-�<�*"�f0݈ا���1Q��E���S�i*���C�neS��I�W�K�N�3T�<�\���*�ռ#��ݽ�����p��֟���G�hb]ؑ�
�D�5�rlzA����gT�l<k��1�o�B,9�Qm١���Ư�,�H=H��8ͣ���bD�����b,m]�~�xÁN�Y����#�[]���eN��Wwj�rw8���XeΙWOkTji�4.j���K5f��Yx��[^��z�r^�iIO.�P�]�әNS5�;B���/�����"���kF�Ӧ$��m�Y���s��'�v�����_j�JZ�q<GE�݅w-KWO���r:�M�8��$	����`��-D��m��-�B�%>OȲ��q��5��m�6Er߻m�ͤ��,�M�'��}���~���:�xyO%F����w�!�N�ڸ��l%f��+��q�@���Rx�1:%�3%�o���^�by��䞞�Զ��^�`�
i�XZ���da��7ٗ��O�������=`�9�qH�����z��j����.�qe^�Z���9�h�9*�U��+�R�u��K�
'����M�J�hp�N1�y9�-)���R�����B��5٭���,���ېD����p��X���P�/����s����|x��ز,��zB���X���ty��Ky�d?OI8��EgIpOyl�܉p�B[�,p��}t{.A"�_��V�'�Um��Q�H���\N�I@��b�(�����}0Q��A��3p�o�K�Bk�u��M�ڙ"��'����5�Wq���u �O��o��=�S���j�Ǻ���{Ku
�y��|{�	��k%�A�jC+�_���:��42l�^G�p�;6^)2� �M}��;�	�����Tɝ'D�4�ޣW����Ľp��n�QS2��x�"IY�M�-�H:.�ɏ�a
��ݡ��)]��X^/'B�i�g>{-r��� �m�<mr<ƈL�ouƴ�p���p��Nw�^d�A>�1׷ϙyΣT.BL1Hl���.;Ը��ږ �8��/"6p
[κ�Pj,Sk�m�L��NŅ�z����)���N����vu�j�$���A]xl���;�3��ˬ:�h�X�*$��mm-��~fմK��/q
:�]��ǉr�C ��¦NZC&V�����u����L:���477��0*��8�0�*�w�n�,bj���Tgv�K$�+�v7c���E�z��`���88^�w�tE;���x2/�f�h�n��x�+������HV������wœrwe-�N-?f��oգ6�����έTi2�q��o'CY�4r�3�,!*ݖ{Z9G�������i�	�����[� �6�
�
d��&�e��H`L��8��eཿ�����;�j�@�"�};{����Zn:�s5��E"m�
��죗����ǖ��+ḧw=K���C]v�N�k`Z�i��r��F�� �!8�-u՘U3�i����ʅ���<�atT]�c��:u>�5��d�W���O�I���9���v����_cn�"�����قd�����	��yD����J���	>��5B���U�ҥn��.� [��	A�n��ӵ����]YQ����Y��\��Q	[)#u�����H���Ov����q�3��5ǖ�"����v8/�-������*�Ն�s�Z������Uy;�Tn�[�#U-ͬ�B�l'���+zT��Y������4Q�5k+r�.��r���2�..�x��≂�g�"�c7Ʒ��J<���}B�n�]9`ԭ�n��#l�؂�!��>Q��W����Z��R��op唿a�<y�4"��z�T!WMc&��F�١�z+��(�U��6���m��e�
{C��>^����7{,D�5ޝӬ�{���
�V:�Vk�1�.�'�9��.�J�Z�����j�)��VuDbs_u�U��&h���.R&::�F�&˾[�lӕ�*�L���ee5�����x,9IoR���̰Vv]7O��R����y���;륋�.h���pV$�zT��u9'�t�g���ݩB�H�؞5kX�x�9��ƫY�6�J�F�W:��3�uE�)|�1�2����.PQt��RL���Zp����+3캀�6�ߵ���P:�3�kAzD81I	��یL��=v	�h}|N*�Hp�V��0�uس2�k[S��J��<yX�Kռ�ɪ�Vmk��b?�~���z��X�)R���Ae-R���66��mXҕ�el�+-*
)R�j��,DJ%j-�mm����e���-�*���)Kk,DZ�[Uj��J",EJ���[h�,�*Q��Q-�XV��2""d�QR"+-�P1��+
�AA��YR�J��V��VT*"؊�l�%�b*Ū�ők`�������Q(�T`�"֑H��QB�T�Ub�,�IQT"�(�*RҌZ�ȌYUY(�1�1H��U$AR*�
*�*"�,F"���TZ��0UX,���X�1R5�Vb�`��m�"��XĭUQ�Q�PjX�F,ADUEDEQDR�"
	Z��E�ib��*1EDTED����>���kN�Sʔ�wiX�Τ�����l/��򞫘ҍ%�1x�&c�{�e=�:3��ӧ����lC����L����J
�7�u�XzgLu����P��hV��w*Ϛ[�W;�K��>E\���m���m�n�m�V�n`�V����N��"�"d(���H�?>u���m��s筝�����6��[,�[,��i��Ț�p3�tT����а���I�A���w�>�<��V.����\��G�J!�Mݳ�n��8�GuXc�̵5;:��t�~,J���z�O~t�=���ۮ0��)�Z�6q:��z^���6��
ֳ��d�N���μ�0�t��f�e�DW�^�XWu쀚F���H�df=������٥Ch�L&�n��u/�6�����e��|2��U���4��|^e��7޹��z�T�%�D׵�F�U��<f.B����dM�Wl�����k#�vO'm{��!����b��k�q62QS�fb���
8G;��bFb�<�þ���/6�ݵ�H-�cnp�2��g���(�sE��|pἉ6��r@9!��y{t��H�&���� N`��+��Phf�4�-s��s�������>L���F��vl��:�>�0�ب]Z��8Ѻ�z���mq���<�wH��t+�uAC��9:�e<z�'�n��޽�י9]�G2���R_A9�SA�^9C��6���K���}{w�u�Mt��1�y×U�X��q�o�	��萕�roΜ|N�J^�^c�/�0�<ZD,���P~�@lb�>�T�:�-�f�7\FV�R+3D�.�c���5(��e�[��RT�C<�d]!�Y��|������B�ط~~ի�V��΂�&������556��P���]i#�2�!��!�U���=��zE�y��p�+�ǉ�u`�����T8�B2�V�k�{1���B�p
����d�$�熫&��r��(�c�l
[�����v��t��ϢdNt8��v�/r �j�o).��}��rI:�,��By/H�X�=�0��nt�ʦh�g�Q�'>�^ܵ1�vR�oz<�br��-R�`׌.��P��v�`g:��i�A�w�fF¬v$uTC�M|������C��┒N�N�Պ�ѻ�v���μ��y{I��F{~neљ�a����%B��VF����]��^�*<��ƽ��]�f��^GO�^��L��o3*A�'��o����Ay�7%k�l/JڞXu$�Yư��m���9D{3�Lr��E��-9Q|
�����W .��[�C���v9��*i��:�:e4B�z-+���u�O�N\
��y�6�B�������챸��]J9w�u�L��J|����g�mGNDc�(�'������:�0��X]Ga��:l��}bT��Hh�c�m���(��%�]��z
�}�z�W���5q���OI�D"�Y몘H1�d���v�z1+����i��g+$U�6;��S�D[�8���N��&��3�o��8�nb��by�;��ZEqSP�t^O%�Br�]_�қ��<�s�>����3��&�Qo�C��j�r��jZ���+H�^��>I��>���řK�D�`�OoN�y'}+;�N��]��W,���X[��:@s[�(�@�}�l��{w(g2�x���`N��I�����J�>�/ixn��u�\#a����Q��2���Z��t�nο���|!Ôjۦ��DYJ7�ӖD�����A�r���S\���#󌭏�U(��]@b��_��j3!��Bj��%a�:C0Ĕ����URۯ{y8KJ���D�5�g�V�ºg50�E����x�^O�ٚ��̷����u��m�+)L��8��(ձBҕ1ʴ��v��(�un����Z��ΥƸ�J��Ŷ��:��Ĝ���))��n�@�V��6�]W{{�G���Y�e�ĥtTd��G�nnu��gx�&x���;��9��= pӭy�[�Oh��Y�ᮂ���(�(��#N�b�+V8���Ќ�Y�����	�O^u�5;iq*��(ʆ�٥����D��(+gS��&5dv��S�D��w�*�ڋ_���Æ�MӖDj%�\:{�/�]��a%Er�$x�п�C���sU(^7�ƻي����$�4u7[��0�G͹�Q`7f��U����E�6ꑐ-��R��\�)��1�ǹ��O�ep�v��Aң�K�9P�lg�U�@���LED3@R��w��pZ���������Ժ�+��,���l�RSUS��k��j{h���F���;!��Ф�vWG�%(1������*��d�]eЗ���!��d�.4xּH���:�����X�T-*u�A��X˭��
�da��q^̽��}2~�#���wT����Z,��DT+����ᆯ�ڳS�M�·,�	,b�4]e���%���女��0�ݚ)�¶�r)W,P�I�q�F�7o�$,�,�Bf����r���tvH֕u؂���5�I,��p��N],�\�����Zwr9��tg<����!C�M�E۽�9EPU2ݞ��^�Ť�q�O^�$͊��9��Ԣ3Vf/&��2�[갗�"�\��[��b�J�y.����E|�@s�b�r�8:�����g:�z9�UM�نl����A��
"�U	�����h���Y}ت����.��o�b�3�c�4�M��NYw-�
8x�o��.��A�'�a��>���G|x����R�.��)�����-�<nԄ���̡X٭fl�c��7��!eq�ND&���L�9�2�H�j�H��Q�L�'��]���9ܝC�������!��+5:C�cR�J�Bg��`q�#=S<��Z]�#>�ڬ���:��oV
ڋ<���C�8;N�[��Q��i|2N�"7�_>u���L>:g����}���,�ʳ�|<P���q:h<�D�ڧ|�EJ�H!i�w���ZD�i����}T��Z�͌;�{cʽʚ�q˥� �T��>�5������Ѭ;�U7O��}\ۦ� �K�'�kK�Z�B��'xc�'�k�������r�&��·(2��V��S�r[[%��,�K��TWJ�N�Ts��T�r��ACu텀$��/ 'GV?S��V�7�m�yx	�f[,�����U�3o��S�R.V>O��3��|{*s
�S���=;L�����#�nA�7�eu��m��ٳ
�.T{���8d��흾=8�l��no;~uq���׽�xP��*�}�������m��&zS݌��.ug�1�_���49ל��5�z�vl��Ӛ*R�n�T�!]��Yٳ����~���hמ-����Gt�w��+�_qШ�]����Q��6.�+'ked����3qT�Y�%I��}w�X	�}�1Z�\K�^�D	г*/a�	��Y������P鴶7յ�C����Փf2���g-�pJ�o�Hz�5��O�\UNӼ�P	�jn�W��a;�ݐ1g����w���D�����7<�8�3�\��q���������ڜ�����il_��q�8* 0V�ഡ�U���M˜��q�"�"�oFR��7ˠ��5��n��r�B�u�d"9�""������:����x	��)�nV�-�$�*��ׅuB8GX��:�Y�
*�.����b�H�4�gaW\�=�C��-
�e��Ïb�;�j������VCyv��4�Q$I�l��9TNf���vm]����C��gJW�T's�s�V��6(j8�	�E��j[�ui��D�緘P��AD�`趧'a�e���㩻�p�Aq9��w����t)�*�{��}E��,gj��S�]�N&��:���9���[ �c��Y��[�$z���Oǉ�x�;w%Μ8+���ϫ�N9\���V�3xu��1b�~i�ؐ{�y5�#>qB�4r�zĆgݎ���v{a{���{'�-k�{�i( }�����o��G�(���������� �6�α.N���Άp��E_]��զo�9�$&V���|���,}+�%ZD�:ٿu��G=T&�c�T�̸x��qk����*j^��Ƶ����I�c������O���H�\T��×!t9
.�roFr�S��I�D���1i��l��2F^������ffd��q�.�q�\jw�N&P����,��V�]E�|�(7,�������K�v���I�y>��o�ޓ\>P�>gl�O�uj�<7W�NIź���W�f���4���/���8vͥ\
�b���O%�!8ѹt�zalXJ�{�����\jӔ��>�kg�.�}WӾ���2�#®�:EznF��#�|��j��SA�Ѵ�ڸ��]iM^;J��Q�eo���j�@a�k��	`�|��5U�.��9��pE�sG��͹�x�3�N�]�i����'��h�9	gs�]����sEkW+{ݙ'V_�Y�M�G��s�=�	�q�C���4H��t�sY}��)�6£kQ�y.�/wj�rv6�sp�WZ������ٝX����
�t���7�>S]���qN���:yyz���	9ڡ��-����0D6
�7���`�$�[K4C�Ej����t�F�\O���v@P��7Mŉn�
Q���%��(����5s�c3)G6�>[�䑅��t]T�J�I�Ks�ze�̆J�	�E��#����z�wA&����U$��T4�XtP�$����x)��J]�3�1��Y�=����h�̫s�%�E�d������M)������T�̡V,��J=:V���0Η;3��kh��� D�{�$��\hOh�;I$J��J�N�3T�-B��<����)u��M��h�Wp���.7�۱Vu��	0��L�,Ϩ_ԡ�R�t6�*����rF�ޖ��
;\��X�C6�(�ݚi�k��9�BM����;p�E����^M!������l�dvd���wT��l�0I/���
����,@���Z^=ف[kc_.��L�/��\
������d,��d3a%WP��[�K��q֟W��ː�b�O��zsN�A���0�[���
�ó/.�*&�c;ʹ�=�Y�|߉��;v%6o�='7��w��_��e����հ[2y��[;[ңR#z�Α(���Ne�6E򳵱���+-��ޒ�靦����.ݑ��a�y��G�>�հ'C��/����a��ve3½�u�B9!X�wdX��7�]���'���_7��d�(���d�RL�,�h3e�\n1��|��"��W=z�f�@Cx��+f�\�r�S��3�6VG˧�G��ꯊ��r̮�����^6�5ᮅ��r�S��n:㱜م���+y�Y�d9{a乮P2b\b�nh��k�,���8�6�Z���vmLʴ��C��s�ap�9p�I�w�L�T8�����UM�نl������XYX��$����~ޜDuo�-5��b�7��E�u��	�NYp�qhGL
��yu�/�fZ���>ř��^8	!�*v;�Z�k��K.�9�p�Lr��A�+yyEf��y�l�>G+�<���ȝI�ҡH&@�y�(��*%�Q��I��-�v쪶1�����qt��IQ�5���;�,��/�֔�%�b�TɠPd���s��z����U&�zk�u����W��gӨ3���K��U�[v���$��Q;_"?���1�t6�Oj��p����P�AD!��X��cwK�q�4wS=��w5�^�u4��4�����],ȷ/� /���>m�7:�%a��Hwso�o�����k�k1a�'��7K�f��Lt�'=4`]GyhB�:������hޏv���jJ��,�>���3��ޗ�[�Y�Y�N��y,���n�N��BE�2�p�[�z-�`_���l�ҫ���T9SP�9t���Swl�������٠�T�$:r~>��{�lR���T�~4	A�=JŨEz�N��! ]�Ƞۮ0��)����بZfs.�����q#G�-��R���54�}�P:]��W��U®�3�+�u�(�����S����W�M�R>kI3��7��# �:�`י�f�>�9�+!��^�S�rX�瓁<}�:��޻��k�������Z��b����7v�e�yZ3T����k�������;"9�d��*����&'-sN&�QBt,ʋ��>�TmjsHP�����S�;åC���2.\ٌ�d�[�(��T5ݕ��O٣�?ypaS���5������Z�x�ɰL��#v�WU�u��D��.�7<�8�K��&��N�������6�K&�1��#�:I�8�
��|p�0�^���2���$��_���B��`IO� IO�$ I,	!I� IO�H@��	!I� IO�@�$���$ I?���$��$�	' IKH@�x@�$����$�$�	'��$ I?�	!I� IO�H@�{H@���d�Mf�#m��q~�Ad����v@�����o��*
�QTJ��QE)J��($�B��P��*� *� R�D P(
((PU��($�UU	�T��(�� ��RJ"*�EHJ�%*��U
��U
�R�DP(�PE{�Ԓ�JTE"�B�(!D��D�()RH�UPUTRQD�E�%)"@��"A"��UBI*��D��� �r�mj5�5��U6̚�UR�"���(LCP�j� 6�"�n�B�;b�Q 
D  �P�Tllʊ��@�kDI1�kR�*�m� e��0[[( �� j�UE"��A@8  nh2)d�* VԳR��ƃD5FB�%P�V��-��@��iFU)Tچ�5T@�E(��)PR��  �u���� ��
TT�k ��-�E(��(�t�
��Q�� QEw%��E �Wq@�Q@���;�P
 uJUR$	HX �a@(��5�4���mlm5�mZՕF��,�[X�SX����ʬ`km�@4-T��"�Y�0��UhTQE"�T�B�8  ;.��*�1�jThh�F���lZ*��3��h�3F�@F�4P��Zڲ�L�ɠV�"�`�	�D��R�  �Nւ�l�� �-U����ր�l�R���P6Z�*�C0���K60�!��5��5�����!@�JPn  .ؠ[R�T������٠��U#T�alM��� �mh46�K# jR�`Е[V5e��[e�
�T��!�D�  �
�MjjLh$�KCeU� �F����3@#Y���MjCAb�Vڴfh4h�2T�jd���m�(��R��*��� ��ء��c [4YKVCB�,V�4SE��,�iU�4`ʬVZʶSM�mS3
ڍA�Seވ� 
  D�*R*�@ d h  "���$@�h M2h���SmeM4�      ���T�G�4��h�����L��h��S�iꞧ��#��
m��I��S�F���0�@224���l�bX-B҉�3Y��Ef(S�h�t���n�^V��VQA ]X�Z$�� ]��"�"t � ���Љ�� �-E"�>�&>G�O�p`���@$1�QPa$�0P��* �Q!�.�� �Emuz��r�@���ǯ��� U �꼠KKR�O�m��P���<O�Pʞ��YK��/���_���{�:��4�l�Oq]֬��CY�L��s5H	�*cgv�L��ص�X�NHEI���C"ʊ����䖱SZ�u�e�>�\��7A�w�K"�`8�h&��u��'�w�$$,�7a�����:�éE�©�Ezd���w�7X֥��o��G��;O���:��X$�څĥ^��&�Id:��oNe��V�M�JNԲGH�����&[����휢����C+�m��>�'{M��q���f:$�3N*��B���=�ۢ�q�xo��F����ݬ�ue.%or�qIw�wMYH��++c�?F��ٕ-[t"�gc�"�Q��ś��X�B��@k��m�uӾ�j�DV����x�{ˏ3t��݋�y��:�ȷt4��5]cB�/V�� �*fk�֋��F�_&��X7b�ε�4h�B+k@�?"��VV\��Z���v�|��:��Uۍ$�qs��E*�f��E��*�m�[��i�"�U{��y�.����C��obP)Ta3� @��K�m<�hH�6�8�"i�]�hS��K۵�I�"��S�x�{@V�$��.2�Seq�_]	��/nU�m��q�q�[x(aBi���N���X�Rb^����ch.�C���@H]ҳ
��t�,�3a�,*ua�ġړ�b-gKC��A��=��Iz�nm;��.�&T�Q��W.�%��.�s@��%m�##����,��6����8�J�k[w�*��LRbˆ���w]1���#��ܬ7v7s*��ol���ҕ�[�!U+�����˖k�ۺxv�#`�Y)�'p]8�0��,�\�ҡw[��Vn�m��N�J�J�s������srVc�(�Ɗ�*��ӡ��;(�:M�O@[ut�)v�FPY�]+9y/uT;r����ն�m���v�E��Hl��ut�ih�����ۤ�EY(M;�.�Gh���鶫e:����@�����X7(���mVJf�oѷ�����r����В��9�w�t�eZr�c�q�JOod���V���Rw��e�66��2�4�d�oOhm��e�xp���!顕tqu*�c�vkS���
���hˣH=8�Zt��e��O��W}�+"���OR"�%&d�rD�2Ѩʎ��ٺ#9-8�)#�����!��G&4nݚ�.���r]��*�bSf�̴�f\T�;�:4�V�(������X��,�+�r�hk��c9�*��eo:X�Ϸn��W>n��J��x�(�����rbG)�N�e�M5w�P8ei̎�����@K�cQ4wM;1KX �e�eAbDp��܅��%�6+7�����������{���x�i�z�c���G�VR�:�f�c0�bTَ��J�-�c5���� W�Ky��wWW��O:�rh�Z�yZ0�$^n���dX؛�G
ݏj\��YCu?�	sX���'Vzv]��Af-�'��݇6�eh�K�@�qb�͇���i�QH�{��g]z�6��^<JY���B�������G�@}|	�+�y�0փ�om�:��a?��C1��w�[w|m�Ҵn|��j��h���,��i�B�6Y']���gJ���J�7>[z`*�x
�kX�*�XVe��CVFdx�����i�-�'w��5nnk�ׅ��U�اk*r�i]Y�g�n�>y�k�e��-MS61`mѸCk��U��=ܵf�H�嵡J�ug
����"պ*�a�ҥ��$%�N,͖:6 U+B���n�/�f�v�j;l/�l�U��RD�2��F���k(��j�n����ҥ(R�p�{F��B^V�t�U����T��� 	���� <͙wW��J���uk$�~�n�@�X�HW(&se
�^�,vJZ�,ð]H>d���]��mḍ5�f���tي)t~|�]��h��P�Xx�%��"��(C5-�!n�F��e�w���X�*יw�S��7� ��{DE�ԛ}�G�H��a�v1�`��u�B�*̲�ݙ[���.V��#V\#l/��R9��c �A�כw[�i]���'y����:N_^�/�ؖ�_*B�c�^�IV}x�flm�'V�o/� N<z��cPƫ2�[�)�X�tI���Ĭ:���bGa&1���f��l��k,ˊ��:��J2�i�QCYKuR��6����Z�һZ�Pߵ�+��Ɗ��ħ���N�V]�5������8*f��z�P�f�zk9�:��*ə%�WPb���h��"Y�[j�u����K.^��<�7�wE@u�,�6�md���l�C&1W��1Z����������naM�f�Q.��Ojȩ@����yz���;�5w@R�!ڔw)�
oI!��Q�E��wZ��nă���33USI�Əg0���+(v�C��B�6���ހ�+��nn�Z��mm�E�)˓Mقl��i����.R��°�짆V�jlmfR�j���̷��r�m1B�9r�[���CnnY���ѓw#:�K��3{n�뮒��(e��`�6�$2.�>�_Wh��V��&���?mu��'�>ۑʀ��h��#���^����%� �q���r�J��72�ci�Y�W
6�)+��v~�˰�Y{��5�E�!��n��Rջ���:Ь(2�ڷ���+(�-+0�XP#Ჯ�X�q\N��y��O�[0]�4�]-���B�����w�c�c7��8*�Yc��έw:X�D��Qk��[Cjݣ�B���ãm��/+L4�n��w��R6w9���,5yf\B-��SAn�AW��]�A<�0N���W!fKlm^X�u{Pʸ����j��vJP�.�a.�f�9=�h��V��n���6�wP[��Z�
���j��Z���X�\�6�B�H�(�z>H��//H4� Wi�F�%,�Jޜ�����!gsc�ޛ�S��lF/���X+]�Ȑ`�@�q3�ΊX������+1��l��Q�ٚ~�����oP	��@�(g*�T�]L,K,���H��f弩�Ed�-��b���]╺�kh��)�8˨.�L�4ݓQۥ�V �wC1붶����Zu2�e^⦴fe��Q�XB�iR*��cP@��ՀsE-y������4�xh��m#�A��9�2�K�kiZ�,��Vm�M�E�N�6���Z�d.�V-իdI��s1 kV��cs\&��s$�O7i��쑼��ыj[��1XܣlY.�e�fk��>�0��ki��YX
�k$T��q���ф��a���3X�R�d�ыN�#N�R��j���|U&d�s��	�	�+va�'NB�ccY,�|>\,��\�I}��م�<��w
R)���&'E�f̂���Ѵ�"􍳖��aa��8*�Ħ�"���t�ɕk)�7Cq+݄f�k+�4�]@�-�Q��F؅:A���.��z�s=�vuZL-��k��������\t�j����Zog��i>�C�M��е��]y�QͼzE3V,�Dd�&�Z���C�'a���<�/k���m�YA���0���J���o���t�֢�#���F摗��+X�jxR;T�q�\v�h�-֭8����9Y�[̛z�~�h�VE�-e�)�t��F��R��S	ưdǨ�ɻ6�Y2�
����'�㖰G_�����\.<��+U�dG.�́V	�]u�c���r-�YD�g�x]p��:2n�*n�ۿ��]��b���t�g�WU��h��mb|�h�̔��$��+(,ۛVywt3K6�9wʋm0��^0o�wVؙYOn�g��B��J�5H�z�F&V7�2�m9�)]�e�ՉZN�ٹ�&݋�o
G^��7p��0��f�-1WH:�4$m�T�eL&���v*|Bz��W[le�V5{�D�'�6���V�w�6��idޅ-�ҩ���;@*M�Bj闆��2](�bZ�cv�r+rcA��* ����$s2A�6f�3&�4�Vlʹ�T�G�-j�W�Z�����v��h���d�m^,���7�[VFG+P�vLP��`��pA&Ջb��왢1,����j"�
���6'F��yC��"x�h����czz�X�4�Ɛ6��i�[�5d:�^�MU=#d��V�*���0�$�n:6�g��x�-�e�i���fS!�P�Mk�D�m�۽є�Y D&�^���
ٹFO �#��wNYY,���K��ʽ���YQ0M-z�u��vc̈́e-7�2�ύ�7�cY�˒of��bgi�4��Y�M^�!Zf��P�#�e��-#O�%ꖁ�6a�᫶rl4*��֒2^�(L4%�w4n^ �o-P��7P-eI��5m�-H���,���J7�[��i6n��O��j��[o,�� ]�m�Z��֙����f���֪�3j���0��	nE>wBݬ{�W$x[���I5���J����ym��
�x����u��Z�M��V�e̖�oʲ#ta$�X�-���UQ�����Zȹ�g5�WX�a��/F�N3��5s-�+Y�|i���#��uDq���t��`��"��K̀��XΓF��w��9����ܚ���A$�@�����Ry�z\�.��WB�d�F+��A�1���ē�"�}KA��>�3*��h���w�ZО���b�=�7��X�g6�=NX4��GB��ѹ
��֭��n��(Q9}B���Lf��[v�^5�I��vc�1�,��=A�凵��0KY��ݖ�s5hˈcű���<���VVQ̃Y�:@�Eiֈ{�3���f�-��Ltī�fc��f#0]�K�XL���ݳo%a2�ۺv��8�F�r���DBy�k�����4YZ["�uc!]=�n�:57#�X�6ݱ7[�hQ��_�wT �귔3��o{�F���P����,�㇉u����v�����`c���}A���i<O]u����x
v��(&-Q
ˆ*VPE�k9��3F��ܩyfI֧���e,�&���Ƀ^�I`A]��sjK#%�n��ne8�F����X@�d,{Ѥ����ʛ�m6���[�t�aG�"���)�E��7�-�-��뚷n�Ǚ�H��Km�b����F�4�x����V�4��ɶ�A�c�Do�y�'�$˳�l��B��^�.�h1���-Xj�F[�(d{��%����E�u��P�,ͣO)��];9�Z�jB@F	���ZE�{��tL��4�e�-(�K���`�V弽J�!.��_k�	�����n��ЙJ�)���h;�<��|9r.��7b�l��C�W���	W�朤��hH�ِ|�^'c]�6�� �;F��7lcb�w�\�e�,�4.�
$�A�V� V�㗄�w�\�<˙��i]��6�dBJ˖5�_k���Ku�4ڌ;��ү3TXA�B�kɟik+��v�'��3����	�י���z�[,��w#�G!�En�G74��H�2\�N�x�^7�7t��r��u�]H��z��7X�D6J����Uq[�]B��`ib��Qa�(�Íf���V�|��Z�FeYsM�eX�����kf��ټL�J���xMB�b�7N�5"����`��	�i�5�[v�̤�D]l5qa�FA��56�Rӱ�b��*h�6w��UlQa�-3��ɡI�5��SOu-��+��{6�>�`�;�(�-�jӚ�'%ą��"��+-��.�5��Eh/b�l
��ӊ�y�2�0�fT��w@�q�.�Fɾ�.�TM��:�Wʹ����`V�:e�A��#���޽���+/V]%A��K��f���#�֥Ph���cT*dVM��h�0�YB�*<�kT�u�:�m{`�ȡ2j�e�-enI�Z�����n\����J״燭�n�R�*�����h�A����{��a�Z5��S��=0Sǖ3�r^�(���R�?Gu�dY4B�Qɱ�0i�̉JLYQ!jȘ�9��`+v�CD:�s/TQ3�A�
k���\�6XŉQ���lc7�z����'m`:Y�t-���m�N!��f\��y��׊�9����c�c�G��b����L�w-b��о�Ϭ\J�U*$��Z�v�%�H*��)�ư��'F��n��$l��*M޵�_#@測<����	x�U��Vb0]c��K�B!���2� ���4mix�m�N����X�rWl��p�V���//��!=�l=s/0����d�����)L�� `�e6ν��.��M��w����"�*�����YR�G�uV�
��=Z8�ۼ,l�
R��Uœ�;ƒ1A���J���<੧��w�_4��f��v��X�Us땮$�U��͇"λ:��״g�"��tK�gw�.��C}�.5�%��a(٬��[�$�ֶ��=�G������b��Pt�/�Ce	�mnv�P����6����ƅۤ�t7)�Y3�V���S��=!U�K,ő�1����8�%��^�̥��n�ͷ&�6�'���^Phfr��&���SUx�+����.(f���v���@���(�zDn��'o6ݕ���h�q^��$`�i�v��^���+�}*3�ME\4�.�o����"��o6��#��{��D�W���BZ�GxVLm��Y�>i*}�gvpv4"M1�J��Sn��Zz�vU�ݘ�`]cf�l��@O���uֳ�^��z�W���Ѥ)��	�Ӏp+�+�,܆�\ps�w�F�g	�<�����\u�[ھ�3Jw�M0��<Q�$�jB�ޕ������ӗ�v�g�D�l:`5\-���1�r���z����;q���Сk{"�i��̎���ҝ�4.�N��-B���	u�P�����K���N����K��)#���gH�:�7%����S��`Q����^m��YQ�VqoV4��K6<�T��vvt�:�w�C�
��ݵm�A�ʧ��stt��P����s9�h*�������ǢS��(�Ř���bS�X+ `Uũ��a�
��LS��Sk^li-�I�5���5skB��k-Pi��`�ܱ�̈N!)���ڈ���M��u�{��ŵ��"5P��ZtQ�8���F�;��e�3��l�9b�����Q�LStk�=J�����*p���V���svg6Q��=��Vnd���E�G����
�7J��&ۃe:Y���������� f�l��Y�I���u/�s��{C3]+޾�TE.�Deؕ՛��ݹQJ +(8�[�d{ۓc�;*6Zr��<ι|��\jA6>�1��#P�җ1�v�Q�Z��{��LR�3�X��(���&��+[y!���N�dZ��������]7�s��<GC��®���������,S�Ph�pPԳ�=�ǆ^��ֳ �,�t=����S�.�ƶ��U��W��Z��UJҲ�t��Ս��ĉ��݄�h�/\�Mt'��Of��Lɶ��#<�Lx[[s��BJq�ULVm̠�(�@ӮK��vfeC]��Tf$�Jx�^ͼ��Z�;i��7*MY�jƽs5N�A�)������'d;7�b�O��;���e�KRt��.z!��o�ncЪ�swYh��F^��St\Ds	���+'1 6�U�IiB5����	�Pܙ}P(�-�z*K'��[�0��;����]Vr��)��k�� N��ԇV� ��ZtN���-M�����]���v��F7����l����j�tؿ*��C���^������"����Miת�7d*��{�u�z���1���7[F'����Y�V@�f���('�qh�xq�������,'�O�����:q��}BA(F�W���-�qx�mD���тg+/^�0H@E`�|���޺r��IB�
�n6l ���N�T���z;����]K4SWCi�q�9��D���r����n��B��R�e8�ݓ�Z���n�9��)o�.�k�p־�euǹϔ7D���ۍ�7����p �����c�%�ʦB��7��%�*l�wM�xz��q�&���̆%��}�!�n�Һ����7}x2�:���f���68�s]تn�ְ�i���/�WQ.�T��.�K��_fŷ�ؼ�����z>I�ˌ��gJ���r��}��U��\���P����*�7j�gn��GÅ�����櫤p��s�mNB����]�y�Y�徒-7�}bi��S�ч�=L�;��,I�f �p+{\j�g����i�[5:9��ř"w"�B#+'n�[��2u���E�٠^�Z�B�^���4���s�,�dR���nZ��ExQ�����t�X6Sƹ�����+s�r��\#���K�b�|�}6��f[(���Ra�F%[�]��zӳ�� �"�_l��ն���������l��W�T�U;(V�;BV��I�Ɉ�fԽ��\Y{Q�#�[Ԃ�2�r�h�&���Y�bx�`e��7m;�
/�g �kj�-޸գQ�;q�������.'�eBCˑe^����0!v��D�N>w����iiS���r&H$�x:D��۫�~�S����L�4i(Y�F�N�e�Vw�Mߋ���5ΥӘ/C��E�Ϭq���n�^Эp5�%e����0�5��<��`�3�$�;6a�uP��+���wY��G8����;NF ��嘳\�6=��3۪6��ε+�8�c���H�hF��փ�}᮸���^��h��:J���A�u�lř;i�[�u5��;:�gyҞE{�ě��pC}0�{�gu���ws9d����@:@�;ؤ��lr�4�,޲�4��X�02�5xE�ְ�]�'�v̰�=!�Wľ��A�֭����I*�~Z�u%]��o�q/�Å�gR�9�T��!l��J�ݺ0�7Ԡ���L���d�&oi���B�ʲ��޲�Kh��Ve�p��rm5x�^����s��6Ps��S��wͿ)V||�{/F�b=�y����.��<����KY���H��K4�\�(Y�h�k���W[zP��˕�f�&��wD�+�k{�nSâ�aۆ-�n��G"���ti��Ԭ�7���4���ɝ��Y}�n�-G&LꇹR�Ā�e�x�5Kʕ�*5��]�zK���Dܽ�&\�Udͤ+/m�yص�5c;P��J1��w�]�Q8̚G�L+�:�--������_H�rB!Z6�
�GJ�w�N 77�掻�v��:�MY)bs��>�x,���\�q�ݫP�FU�]꜂��{�΁sV7D�ڌ���d�8�V�B�YE����x�h���̷� -�5][��X���v��B;�M�����
őA���kyYnw}��(�oJݳD��2��9RV|���ޘ�S@��&�uX�:�kfvP�W�=W�j�}����էYɳ4W}��;�����2h5[��k��8q;,0��p®����s��(B�m�pS1�.���ͦ 7��k�su�%�3�䅮|c�іC����	#��,ǎJ�����L�z1�\�u��Y��B�;u���S�����&�`�Zۖ%����өv"�U�� � d,$Nfdb��k��7��r����:��Z��s;"i��`WO�Oi��ʲ�2M�e��n���ǣ��l�ȃ���O8��j�~۩*���u�H6]�i�?�]���J�}HXy�s�ШH�hs��-�:���Ib�,�Em�ռ�4��Ն�i��n��]�g���ŹZ�U�7����NT=��:�`��v=�qS�Dk}�z�΢�	�X�s��݋S�jŖbm!S/2� ;���`(�sv̴��C���X1�;�KkF�遠��~qN-l�1W�&Ӭ@�b���T�e.��=�:�4�Gʅ�uw��l�@�2���Zjլ;@GR�kv:Z�7�vzM.e>��n��i������{LJ|��"�̜�A;X��C�A���޳C9*�[�~�D�ʺ�sa�[._B��Ygb�Z�\L\�]��E��̨#;j��b��";cFtVd*]-���M��hY�X����G{�*�·�pvArZ�.��nAW�O�V6��#�Z%Y�r��nb�����e,�W2�uF=7����
%n��̊f��LvZR��N�!�����Ń�#R�Y��zN�zny��Դ�E}v��P���M��3V�s��Q�W�7�E%��r���uQ��"�'�1R�e~��>پٓR�q�u%�1��Լ�ϨN����N��5���3����5�)d�����!��0�;tΞ[�	�g���ZSİgZ]�+�f�R|���N�;�l�H��>d��ގj�Sg��\��AVЄ�1i-�=�k\����K�[g6�*S��J��ݞW��^�kt� ���Ǉ-���#���,6\��O[۶ɺd���ϴ� ��T=��^����lv��F|�Չi튙a��:�([�N�70�O1�]���9\y�\�w�P�rf�w/��M���"�w9:��Fl�5;t��Xo���@���9�i�󳛽�A��Q2~6�Y#I�b˕+\�k5�7��� �n�����޷g�V�����9�p�e����ၷP�'qf���3j4q�j�Q�ѲT���ٗ!L�ʷ�!X&��>猵�l��S��&��uѲ �DU5�3��Qj��7����x��[�,�����+ئ&�B��ɹ{�\TiV���7�t���8c��:����d�Ni�w3 ��i-z�x#��ې��S�:�Eiw_19qz;1N�� �V��\4�P�SV]*쵒nJQ���9�,L�b	v�kԇ����]t(��/�u���b��Sf�)�O�����I�p��ô6&>9�֠��Wy�� g�2�ڌ����%�,C��¼d�"�S-g*��#.uu�U�����0pױ%.���S�l��ө�0e �����[�<*&&n�oTH��8��]���zR�*w	U��SOe&��̋@�Z �r̾�Y;Vt�0�j�P� r�ˌX~���W�c��o˶X�Wʻ�J�Q���,�xy�a�)cά5iuJU�؁$.��]�pۨ�k��25�gV'�֭����ʊ�ll��W..d]o�]�����K�G����x�VN�����I�8���ܬ�5��݁u���2��!���-��
�w��! ����Pl��mk�Ƣ�6����Cl\X;Vqf�.ǩ��kް�Vl����&AJ���ZV�c�:uE�'��nU�6�[z�d���Z6S\y�EF���?.l�E�>��
�r���;#�M���f�G��7K;_KF����,��Y0mn�j)-�:���Y�h�6��Ch�Q\z]`�gېJzjLa��;n5+�r��g	�h̜�[��#0ޛKj�
o,*����\,��kwYם���MT���7X�<���,���38�"1cWG9C�έN�K��(%����F�ië�SNL�	9�M+���X��+B=�ր�7l��Frh���.�XavY)c���tOx�A<2 u�4&�N;���{]ǰ�f5X��n�gQ��[J*ض`�8�s�Ւub������9�^2�+mͼpܭ�.��M��}�e\޹}y�:��]�v�ns�zR�mN��S
�)��V�s�G3�9r�Y��܊���֗Ǯ2���*#��ծ��u3G���̀�Բ�O�.�S1.���εCf�,�h�Sjt��t�Տ��Ή�ot]��
�m�2a�q�$�Vؔ�c.Uͽ2s|��Ե�L���e�8v2������:�Q�ܣN�h:;��TX�%E��l�ܥ�M7&u��Q
�Pn��[��Pdf��[�}r��U�<�'�Ebh�\���,}��
(d�{kt��uڤ�r�R��.%ܡ��b�͑5S�v�z�r}w�iR
�so9�pN�Ŭ��a�9�|3�sp�[��˕�L��u˳�gc��P O�3�Ʈ����e�vj�K2&[��ƟbJeG����a�p�oT����e���1 �E T����ô(�k5��ή<$�@]���I�[Ϲ�e�˺Yu�+$�삔t$+f� ��n�/o��&amYdpu��HL��N�]��ޤ"��.N�Tl��r��_wR�FT��X�*.��w#�v��0*��]�;}h���+N�D�R6U�����&�N�@�&z0�P1�k�odV̘�f)q9|���q]ʏKޛNr��L�/���+�n�VZ�IΣ�;v�fN�6Npț�$���dyr8�y&%�1���E�|��#��I�!��o�\��]��l�Q'L�S�/gBg7b��i̓��5yg68�"��wq"�)͏i�J/\�K�w��ޔ^�fV�����'�ޡЄεzu��RLW���ٛ�6���@f��}mS�n���W,/�;]����|��1���W�J7�K]�ቪz��(�y�d5��nnK�Ȓ��F3755ow37�\}�ޱ*�0t�J��}B�p���n-b��#
X�)�̮��X���ac]坠z`x2Q5�!�#��|��mF)�pخ�d����3R��`���%�*�NXN &����<�0ǘ�In�����TTc�"	��K� ^���S�0��@�FP��g���LV���^��r�6��Y-�F��M�iܥY��)__R���-�Ֆ��ͫ6���F�\���[�hC����aJ�X;�=}3i���iВuo��w`on�hmnm����g2�uX���ie[VJ=�i7�:��<jѕb�w����.�PoE�nr���N�d4<{2F��Y�N��b��m맒�d�â��0�<wۢ��X.�=�hl�{j4�.��e���d�gu,�N���%m��P�/2;�v���t���Kc�+�`������}�5�!XW���+�
a���X���֥��ھ�b�A���Qn�|̿�\�"�G�Kp]sV5U4;53��9��iSq�7*� �K![(�r��{Zd��M{KA�Vk�Yqv��Z��S[A}��On����y�yc-�۝fɔXx�+�1�8Pי�5�c�$/��ӱ�U}y%;1q�h^��tmp?�Ӓ�oa82��\�`T�r�mF�|:;ϟֻ���L۵w��A.���]"��WV3���V�K�gt:j��q�w0ңU�G)n����vΛ[r�e7��;P�Q;"֋�X�#Ǡ�N�6��b?�-�:��2=|��,��zs��r��A�=˜Ew���غ���6m�{�hN��io�:|�7���rV�L��,[J�8�m�1��M�u�Nb����8��4n��b�$��G��	���d`=�H�3��,��X2�Ș�R���k�)V�*�*e-���ɗ��5�g��[k"�viDfW{�MɕIQ;La"��=Že��ʛð��X����f[A����6nӝͱ��+*�����<]���f�N�¨�����_C��݊��kyKF��@���9!�|����o�-��gp�Vť��i��r%�ئ[F�"st����ƽ���7C5��nMYN÷u�&�4�T���X�u�B�wf`��$p�Y�F��P�g� 4A`��2j��+���v!�{B9H�.A38�:��R|�����a���[�5��#4�L!�K��]+#����b&���.�tgbߥ.2Sn�ǝ6��ivG�P=�ZY�"&!F𠨝�XK7.�%W�P�Zޅ��4�Yn�U�ݘ'P4�YJmf�PK!^�{(�]W63����7R4Zkv�)�;�x��L�j8lW|ej�,!���L�f�6+�/��
�{�ݫ4d�k�̓�-a͘��3NZ|ml�Z�)f5o�i`[}4S�P�x���7�]�о�r�;���4�����>�C�ⱊ���+n�c~̵�j8��i��ZW��0���QR�7�b�-��X����y��z 5^��o4kWi��N�^�aMđz��*SQT�y�kL��vu�t��c�`����#�b�kk!w������W�W��B5X��i|HV��˚�Fl����zi�z)9�&]�J��y��5'�X�4�+T����������)ȧP7ݝ��N����jk�,I`��2XJⲰ�(��]|��*�E�ݼ�-Ӭm�V$�Ứl�(N�z�b\v���E��헠���aD��b;Y���ܤ/nK�$v�l�xfv�A�M	v:y��M*���>�c��b���U�Y�Dܒ��m����Jӎ�Ԭ�6��t���!�&!����!̤�P�l���bՇ��*��J�|���Խʇ�yVu��)������0����S��[��Q�6��2�Wr�\�eМ��V��#{��W˃��b�eE��5����]��wظ̺�*�k�7�E)�P�d^�]Y�i��:㰑n���u��ʓt��F�K��U�{IVc��A�Z)C�:˫�,b��`�x4F�Ms�M�%T`X������x����G^u&`�L�rFE[z�Ai����lm�:Wt�kƪ�.ĥ�Z�gP�����m�̴���t�u�Z䶢f(����Wi�;\����GcX�p�ڲ�h�5ݛ�d��{1� '�}(�F�	v���cz##��G�)WN��O��]�ZO)V6�I��+��y����JsxVF�����sTדT݊C,���ё�I���ўU��WJ^͑�aV��6�^41h��%e�`e8p�]���C��dIpK����n_6 |��Wݠ[��\�Keнtmm�nK����R����H��`@v�:�5��/�ZX^�|j@lR}����ҨKj˺l�r��.��&Q��ȅ����8�-oF��J��;-]*�wcl�ی�L�DVB´x	zgY��*o�tܟ2jWIˌ��=�Mp��@#�^;�Oqm̀�}�;,��&�}
.T�)s���u�-�s>W(��s9<��.e�'�bЭ8�.�\�J)��*Q�;"5�+�&�eM�g5�qn��� 1����t�
���<5�m}��N�y�R�N�v��|l�;I,6f���}�y��2�k���b��t2v}��l5��9h|`F�s�wl|��{Y)J/�)ͦ"�Ym���K뽁%��]u��0�V�ţ!m�r��=D�;B���~=�%�Ԑ�)�,�ڳ��.�9���Lv^Зb�m���;4��V��4�G�XY���D
͒��{me�Ո�ǵ���p2ΪX���5IH��=���nS��US�7M6���7�v#D�!��	�N:YT�%}Vd�'%���v=���th�-F.�:��A,�b�A��ww]sU�(��>�{k��X���r��+��:�ѷg~bH^��]�Zj�\J��"ji[�+]K���r�Jn���Jp�t��d������
�w��D'jf�� �\��-8f�n� �AWYԉ&��w��:wu��l�v�K�M%�ui����U�2����S�hD��
���õtŎ����nm�u�_d%.�����"�Ѡf�E��X$1Ugv:��m�rf\۳y�:h�+V{C�:̓{���f��Q��=H���޵K{Zv
&'3Y�&-xzr ˺7�F���o�VE��7���ٹk���}�(�l�(��6;}���ҧ�/���3V�宰���*���p��#a]�R�T4ؼ����n̢�c�ˑ�0�l=T �R�}8�T���C�����a�0�t�K/e�r��;�
w�k�E]*�iˣ.�U�����a<q@v�x��*�u+��*��Ƥ�x�:�8_ ֮�#�VH2�F�48��t��ͩH�09���6���+n²�/�jr�,��Xw�j!��`���fr66�k�ܼ���(��I٪Ql�7��ú�H�J�:~�4j��;9v�]�qR���TD�!��]hXVq�(X��.�N�ʶiPޛl��fˊ�� UHVC* �Y��]�E�0�^j�U9w��%i-"�9�|������)i��&f>��vE�PG�[ѽ�1�)���#q�Νn�_L��j(=ymˑ�x6Mn�3Y�fW��h��EX���la9���t���p��(I���h���r�i��v�=N9s�UMp�lQ�.pKJ�ǳ)�-�� �Qޱ��kt#����Vn��{����wI���*(k����g:WiB��ߋ�;�'��tp)�1�G]]IN�]v�|A�$n�(��ve��
ڊ��'���3�w�&�g3��1�W�X���m�1�lP0��@��T��D͙���%�0���z���4���OL�N�M�ô��2��_E�	�]":L�J��3���im�#�=U�׼���݁f���[-�bM��ɀ��<� �#��m�9���@DV5��[	"�H�Sc��Lʎ����r]���S슍�)�s�aՆ�}��� �OxW\�DHZ�r�����K�SE�Ǣ�`U�{��\�n��)�c�<��܅P*��]mΕc-�Y�2+�2;�y�a3樋�5��(c����4~p��v�Z�N��aQ�'oYWB�'6����[��&�4hd+ަ�=1��q� ��a�>R��m��<��q�U/	�UAM�6���@:�7L]�H�Wa�(���A��<����`ַw�%]��j����f��ǁV�vJ�Њ�g\�lI�SA���{�`E�`���/-���"k #���_�!wڲ��6�d����9�
�u�,e2[���bd��,��y���d=��V��:��I��,5�^��n��U�9T��Tiv"n�7���;z�P�A��P�0�k6��y�}�M���e[��Q�b«�Ju�_m���xzRJ���.x*��3��H��>eg�Y����f���D(�NԷ+��C%�7v�xӢepX��]N�����Y�H���-5ƵJ��+,p4g7�
;�r�3_N������p
U���֧l p�a^[P?�w���\�IN�/�����2�<���	�]^Ӧ�B��Gr��D�g0K���uƶ@ȱwj�Vk�̝�Nv��&�{�HW1��Y��]A�*��y	��
�gq8��kT�ũ`ژ�_v�p��^v������۴���t-�'���v�A��y	Wn�i�8����ٚ�ɭ��'\������0������7�(��p7�����'����#7옓������vc�[}hSO%�+��g˰���OS*}r.�j9#�jr抻S{6� r@Ҟ�TXھO@�\F����͸�Y��E��e��v�Pr� p�/��8�4��	��ֈ�yCF�G��7]i[��hQ_I���0���8���V[���9�jfc܉U�N���<i�X�!�  ط����l�ӹ�x���lfR�66Ei|�X�{o1�
7�����u���n�J��bZV+��1F���d�BV��Cf��y��q�//���(��K[�ԛ����EU����)�m�w��R 9(+Ph��#�+;7Ӡ�%�عk+�A����!�J����XLLإ�]�v���^�G�
�X��8%�,��'�u�U�*I�J&��X��`A�TY�;��z;D;��Z��26�%]e0�e��s<#t�.ty�=֗�xɻP0_kV_q/hN����:�e�v35B��f�G�$n�ޙ*�q�w�T&�u$����RK��Z�(�V
�}�d-	5�B�A�P�/4qx�_M�ڈ��noZ�GyX�
�G��9B�Jy��M.�;Њb@Q����&�7}�f���]��3��)Ҷ�.g,�0���8k|c�z�D�P�'�O1��;���rc�r/4��Eu���=3iJ������9x���*��ھJ�l!����.�G��BT��S��{�T�˔��'�-��i��ge5ȁ�hn]e��;[��t���4�3�H�E���H�ԬQ�����h\9B���͸��;nd�[r��*���c�F�!��M�*XԱc�\�zK��ݫi>Rʈ�ܺ���$����>��6�a
ԣ��h����5�P���W���}]{�E}(>��-���qGq����J9�ʉ��+�D~�̚�t�����<#W������ދ�#B�8�TV�_>䀵�Ι�*?:��P�:ḑ�r`�{���ϻa�Llo*u�M|�&���7{b��d��C���k�$�S]�to��I0&�'����Z3�y�䮫Yu�]��Gvk���v0��4��]�tP3V\��y��Ǧn똫5}�`�'���`"e�礬���ͥ)�4Ad�U����W�Q���Q8�-I����/fѬB��ת�o6ܲ)O9�rdʱy���lp�!+ޙ��B�N^DW&�]�/�R�lf�:UEë�#�Ր��ژ�GX�gLF��]���F�.�r�<§t�H����4���Ҥ.�hf<�;Ƿ��*�J�4*#K�o�ԣ�Ehs�Q��a�?����;\���,�QfM��3�b�\��^���ڴ4V�yb��z��"^��QPt�oWR3�n��y��R��'7�h��}w�[���j�kN��Z*�
u^�X��yP����݁����|���D�g8Ѥ�)1[�/^�}z����]O��9Y�wՊ�s�E�q�Țᆟk�5�>0�AD@�k�D�Zkwf�S��Is�mGΌ�-Ü2(��\��̔��	�p�m�6�){��-�h��BK���#E�h���Z�s����B�ݖ��iC�e�%3���CV��2�8�R�۽�z�7:�:)Z&	OL�P�����q�En���)�r��ļT�FcKn�љ�p�a>ʍe�����}�%�iG2�D/t�»���6]�̺�*%����7����Xڗ\��Q<�jr�xʋ���Ǡ�9�/17�AE�pLfVW,ML�2�5�-�I���m�P�Y�cv��(�G�i뮵���[�O֐�  �_��K F?/���~8h�d�R��5�ּ����;ց��3v[��j�Ԝ��F-5ud������Q�&�t#G�Y���+�G{P�ɟ��y�,�O�p3Gy��[�3����Xlԕt:�y}jd+ѝ(,�����x�����K�����R�OV���zvH7-�L8�e81F�V!CxQǢE�i_+��#�]�x:���G��3�Z�PY3/��K��]`���3�H�fFt��ú���U����ƞ�f�Q��-�@ݫ�S��eGC|Ot��z�8��n�a�+�H�V�͠*��l1  t�W�n�(���γY5w'Rޮm8퀻8<����ޥN9j�t��:��7���O�Y���%�t���ZROy>��MK��ݳ�6�P�&p��U��ۂ����B�Q4L�:Χ%�ń��y
~{�۾��VA/Ii��K���y;9ݧ��=A�����.o*�!�l��w��`�m]�G�왼�.�V�$�������㻧l�7;�ݐ�F �r��䵜|}h��ԦD��OS����ޙvv�J�&����L�M�M�6(j��S��B]r��W@ڕ%J�9�X�*��(9}{}Xz9GI'�&0��d��P��7и�ݥ+�B�'�֙�z�Z��}n�୳}|�ʅ���F)�屝�.P�(,��I�UD�R��Y�HJ�FLd��m�*����`T]8��XT����QQ����ଋ+%`�H�:h��QA��X��WN���c��4��J娪��UDJʀ
��
�՚"AAdX*��!ufeX(f���E�*��*�Y�іj�cb�`�)�a���YP�LHv�Y�H
:���Y��(:��B��,m��GV��%���"�&�TQ`��4���*�@FA�T���T��ĔV��bT���ɉ�0`��AT�!R�&2�E%VE@F,�lY"�u��H,Q\�%DE� *Z�H{���~�y�t�o��pҢ�R���*a�b_8�'���G�]��T���'�զo�����1^��˭4��[νF5��n�)�s��u��xʲ�L�j�ol�������\͟W��L���-�U��̈́dÁ��2�#~����<��gs�y��x�ݏZ�Z&	5�Q8���p�z��Xk8�TY��PJFB3���A��r�*���0-�K��xy���cdε~���_VF�Y����T�
���0hr)eW�W��Y���J��*��*'R���SӪ��!�6I�	TJ.bć�{�;�v����NWB�/��Ui�y|��#��#wt� lH0���j�(t��D�łޥ#�Q*�{�W�:Pxa����TR��c 1MG��k��_O@�9\*QO�oh�Ӊ�K�u������p�Z0J�����(7��%yǠʣ�~��:��K(]�7
�3` ;��HX\AB}1.zL+��zo�ϯn�u�P��a�ͬ��(�[S/"�9�܄���㪲a���'�%���.���{�x���%��?K������DP%�PE8��*o�P��n����&B��WVv�9�i������][��N:l��5"�q_*=Z�"�H!�w׺�K���6��z��Rƫ�*���"F���w�c����^���QNe����.W��s:-O��W�72N`UD��ϣ�[����!u;Gym���5[^\,�+�U8ܞ=	״1Ra�YD�d����0�AO�=�]��U+cy9:���"�
Β��~��`7$,Ryw�,:;d*E-�ĬUا�Ü]�͍70�*K�u��u(r���'���r�e�������g�iS�L囕ꂯ�tO�UpT*��Ge�Sұר`uMM�G�~V�<],ݟv�v�iԥ�`O���q��#�7���&#B9T�_�G�i�ߔ�p��0�����Sd�0�����F�oj4m���::�4Te:�OL *�|�U���*�#�����5Q�E�~u�~�ާ���i��ò8;�Q�e��=��w�<;�v's�.�V��gCG$�|el½2��K��O+��"-�p#�e����F������i'��.,Ԩvx"oاʢ.a�T����{6\5>���:��q�ת��V���c�GH�=2�^�1�n�pɭ�L:;��,��c���I�~�+�Y�<�݈˦Fr�[��Q�M��}�2�wjb�t3�oN:�b��Wm0���貌���m�5ؾ!w�2���K����Y��vΘ�ѻ�'�?���Li�\M��y(u��rs�\2�� ED��=���Z���$=�WG���&c�[5�[��À�x����'�y�rJ��\ ɱ�m�3ʺ���<�eLY<-R46�ȏ���j#C��.�T[�R��ynn6��3O�
��m����ڗ�.�c��Q�*����s�8�C���,�	{���(���V�)恍�\�l)�Z���
��Y�L��x �w~Y{��K͏,oF���T�p�b�l��&����r�1��U��h�o=Sљ	C6�r�y�v�;���B���B�`�&��3�ٿq�A�l=���UpJ�-�dڦ�T<�V1�#;91|�����u��C%�BF軈,x�P#z�8���U�܎�i��u�b��`D�v͈������W.r�j�mN��D�2����`���e�V�98PJJV��ռ���^0?jЃ�������ƹB�vi��!��Vo@݌��;u�0^R��$���b�q} ъ��v�J�(u�: S���b���W���<�YC��}[�X|t�"�x�V��E��;m�%�Ai}w�\]t��o�i��o�ٽʴ^J�w�$�Ymƍ�;w`�v�Z�wÕ2��ҡ�T24�^��/�dX��r���:�&�L!�r���M���o�];�2��ീ�m���5m����u�C��'BQ�8.�T/T��k/�r��i���3LhޞR�i]��'ox�4�"����9:ˁy҃�ڤ"��P�xe�<ۧ�Q�2:��_O9c9�Ǻ���n�G bߌ\��Q1�.����&��*�i�pb�]!4��+f���Q��4;_+B��,1qd�� !������>ae�EVE�CW�Wb�	ܭ1�9�;ew��m�w���t��G>�����+��%���E&��bck'��������LZ�1^�:'�t�c��I>�NgZе2ϨEԦ�=�
l�׳�����������۫P�*����b�L�=;����(��m�9����Sp��N��s%���Ej�yT��z�b�zQ�����4+	�Up����p�M���^��<fHL�������!�"�ھ��gm����}�1�]�U9��f�ܾV�^�U Wl��� 7~���Շ�z�׆��q6m�̡.�ŕō��"����o;r6���>\���̙�!"l�̝h��6��_d��S��|�k�E^������� ��OL+�A�}߇�M�ގ����+ܣ'��8V���V�����[��Nmh�T'����
�X^Fer����QK�s��ѯ�^��B>�=ў3]n2���4����	�Q�I�OW���M>��R����S�+���:�7#�
�͹���;e৞��k��O3�S��k:t+5�;���{�R5���6/k���d�S�����ʢ:]f��x���΍�J����	�6y��{zgԳ�<��Q>:�T^'Q�ʽҩ4:� q��f(����p�Ig8o�nE7�u�$2j�c��S*'�S|��4#c��1�j��=k��<��Jyx�m7�u��4�P���5L�]��V���M��`kR���I�A�^zm��a7R�hؘ�����w��f����7�;@��؞�t73�e���=��R;�^�N�9:8�����r�7���u�ǹ-5^�%�*�m��侩K�u�W��%v��V�j�_L	m*�a>Jm�&�T�+��5f��+�T�#��ʍH����)mgE	��4-�����J{Ʌ����>*��C����R8t�\�_�z�d�����o��W�'P�en��:R�T�.x��[�'�K�숩���17S��}zdokr�:s<-��n\�J�f�>��I቎c����Ԫu�U�&1<�Yg�-���o��S��ۏ9�u��h���|*���1'�պͻ��5�5�o	QM���\�8]v�k]P��/�'�f����<�ؗ9�}qV��}m�\����Z�%;�h����ȥ�"��Ƙ�?�Pq��][�>�Q=��\'������OG_9��Z��-v�j�]xⓒ��3������5=j:�� d>����o_�����ä/��8}3�rR>�{נ���z[9e*��C�@j��MX
��z�:HmwT�Y.3;�mN�K3�X���h�v=nB�W-y'-d�|��O4���S�����^\�Vvj���� [4�:5j����˩�k6L�Ǹ7��ӝkkb�C���)Ƌ|���@�&��z���H��/{�K��{� �ʋ��zTXy\��Z��:��8S�Qҫ.17�[�QM�x�̵�v�y3膈RΖ�7:�3η��4�oI�8��<�u!<z��L�����lvM8��-�9S[����*.JQ%�*�*����O���ޅ��S����U�4 *ė!SYX�c�`v�P��1��zw5�>s�S|Ĥ���>|�U����u=lh]q\4s밹���Īs�2�$��F�
���Y���\�v��:�m��:'��_��$t�Ƶ&6;��ŋ����pZ����u��4TG,�Q�O��lpK0�s;4Y]�?x-���&�!���`���WS�T�Mä���8dd�}^'Q�|�)z�V�Jª��a�g)���r9<~Q���78n��R�Ҧٴheޕ
W�����g+�.�.�ˏsh�{�Vt	��דL� �jj����t�����X_n��˜jA����Hk(�����J�\�&�����\�й9�XW`wyc+v�o�JS=��6������nٳ��L�Uc�0ߕt�|��ˍ���P���T���O��5��XKk����H�[ۋX3({L�1l�;}�E�n����p�_r�Uyv�uz�m��@̠}5�MV���]q��1��7U�q����x��?�e��ޥ/�DO��/8�7%_*��JoA�pԬ�ڝoka<Ż�ws�̼;���3*1kS:R���/�<���������r��CKt�څ�&��BuM�+3�8y2�\Y֢��:��Qҩ\F����N܆�)q�k�B���g�e����\���Le�Ur�G7�Y���(ȕw<��I˕�L<��@N��ѹP\pS9p��k.;�|��y�6�'�
��p�3I>V�vk�m�v�>�:`�n�z1]M��o\[���G#g0MY9�{=�������+��5����	wE�Enq��ҙL����{�Ů#	ÉU�1�Zd?�˗�pN �����Ecq�|�����*�rҝc��[�V���כF��nχ<��3r�GR�Ƥ���RM��bc~��O��/~��1k��G1�!v�yNF��L���O�Hpj�������x�B��ފ�Y��7U�μ��}��,�rg2Cb_;��;��w�tҭ�X�[MY�� ��]�9ٽ�a�+c�\�*��N,�pQ����)QO$]��%�/�B�>����Mà�	�Cn����TO^+�7���o�9�.aw5{8�'p�!�Î���N��X�amg�t�u�x=�v���ǡ<��]h�@�Q�MCC�?k���G<9Q�m��)L����:�G��{�h��׫��1[~��\�jCg+�j�3j��é'�n����`8�B:#��������-)�
����$�rR���3��1;�^'%���x�a�Q�Yz��-n��s����dy5�L���Y�TK�D[�@.�7"��N��J.�w�n�����U`FS��W|��ڻ��y�b�nK��y�۬Yֺ�Z��;5�lW���$[ǲ;������Y�y���2�NGm�-�<g�%�$K�!��/~�xJ����O+��vy��Tܵ���:��e<m��kA]�~HeY�ڨ�P51FMna�PC��X��l�Y��*�R�rǏ���Oyo�#2��Te\�W��[h
[q��橁y���yx�i=v���+·�72���*��K�F���+tstnr&4v���Z瘺ViR���0��D!!��Cܘ���عº���q����,����Nio�I�X��4�7���jurx+3v�m�~Ρ� ���K⪵�DסT1�8�w�..1c���v��K�Κa���?s$��J�'YS�8]�]�5������~(���U�j�S��P���h¶C��P�d�E�L�h�J��
�y���"�^�Oj�;��ry��Y�a�@�V�`{�ǿ�^����g����;9ب,����v汈�c��,�����M�isWx��Usz���wR�i�1����T�w7�="M��[ڐl����+cC:[x�2�5܊��>Æg(�����*�#�V���WC��\�����*���=n�^���ͥɉ�kS]\��;��QB���۪�\�@  J�����v�dm� w=�����>��1���n�<��v⡟9i�f���%$8ٕ�,=Îf������S��^4v��r:�9P[�u|9a�`,�o��9�,r�F[̺�����= ��iRHW4�4;���º=�}�k��MO�f[�n�B� :wG]dĹ��69��1�^C�jt55˞��L��`1N�����>`ß;�nei�s/��E�@�C :��Q��C���V7R�s��b�7�ޕ���*X�oV~V:pgbtNE1��r[Y< �-�5ƻ(ɽ��^a�*�ol-�ܩ8���c�D��դ�Z�*v;��R�ܰ�)Y�39��F�2�Y��X��HTq�N�Ε�3/\���ѥ�,�x��yH�Z;%�8��:���Sv,�0��O,z��������3�p٠<6(�ĭj\��Qqɷ��=��Tϴmk�ev87
n�4S�W.<wC��Ի/;���h����;��@8��|2;o�U͏4���,b|��-�h����}:�c����@����_�L�P����j��X[�e�]CC�qnS�.�/4Qʾ�R�j�����&��ZS��ܯ�kdB2�	Yз=KsuR���PӚɚ
��w�̛Wy�8�ԵI.�9����\T.��ف�Z}:�u_Wb��M2hԻ���W���^��UkA��(�����Gm��ں=P�0{fQ0�X�:��g���PM=vl:ǻ�_<��wN��g�4t��y�yI��w�6]	Jw��UtC9oC�oD^���U�:�7����M.:C8m��w 0�)�˾�0�#8�dM`�����5y�0�Tb�'\͝l�<�6�8�K�<����+� ��m�ѱ!Gre;�����ջV(VN��i�Xms�6iܿ����#]޿^�R�
��C|4
�[�at��X�!g�8�'��GMWtãqX�L�7����Lz��WGz�7Dz�,	�*o��U��ǶO��[�
�I)���/cB����.��ҋ��Mܮ�Y�I �6��p�4zN�h��Y.0�6nք�enlA2��q��jt�Z��J53'RO�=�/&|�/�]��R���48�'J��\e.�GRޒ8ʜ�I�ovh��C$Q�ds�t-ɀǎB'k���Y�����N�p����d�VLT����m%f��Qa�X�,����ʋ-���1�#E+���( ꒠��i�@��"�@.��@b�)FjTbDE�bLWcR�b��*�"�CH4�D$R�Œ(��&$�I�)��RJ �i�Fi������*�@�+	3,XbERVIRi�jVH��1���-��
Lf c0�
EQ���!�A�EN�e@D����P��b��Q�&!�i���eM3"Ķ�T�,�+�
$��*@��	PD�,�Y�V.1��[��XJ��̲)HV����4���QI�=��:�9�yu��[����fe,MC��÷7Squʸ��9���	Am�ؕkhH�I�q]��y�w=�B��\o�Kms�F^��VX�*�Š:�޹p�Ez5�L't᝷I�27.C#�p�3�Z��m����W.���ߜR�����ℕ������a�F���?I�6� �ʿW���h~�g=�G~K�R��~e�f�2��i���O��p��2�O���ۄ�rV�>�c�x?eJҗ��W��/y�Wژx�gz��7��zf"���-��S\
�h��n���p��O:�L���/y�[�-�=
���o�<�fq�}��v�K���p��⯚��z�)�!<x�D�o����/��\�s��䎦nf���ɋ䨭\�>c�w�³X�����Āo���)�,o^Xѱ0�P� �&.i��]K��̽v��*�f�n�#��[��Я�{O�1+�s����y�J����^��a������l�,�B5�Q��(��J�oL`��V��FW=���F�B��]rf2uj�����u�8��l:�=B����%��8�{u`N��U�وA����������H��Ԙ��u�sƲQNM�	q����L���߫ȇ
5M���:e�K�&��P:h�t��w���r�R�N����*uM�{�^���N�Ym�7���j��Ht�~��SE�ӯ��O��hY����b�<F�畁�Yݏ��=oX��X/0pg.C�R�{���_���������.Ճ�I��a��ך<��V��|����~ٸ��1h��{)¹Ą�ݕ�������ԥ��g}�on-`��{J�/"����u0\�V�K�P۾Qp���2^�Mz9���/aua�0q�s:{lz�e�����xѾ������p��̼;{�_���@�����X����ұǹ�ˬ6�ڝm�;[1j?SIO2�:��ݩ��ZD���c8�r����"zT^7ч�GJ�������r)��&Ø�5G	��3"�o����@�S��cO�L�F�˸;������7ff��-�[�t%G�.V�a/*�=���%��a��7�Q�����"z+���E}���o;�$�g(ޭ�wS����
�'���z�in��̸wu�����ܜ��D����Ao�	�2U�J<�~O&���㑽������.��g��X��k�ڡ1��:t�Q0u1W�U�q���'��&Nn���u*�5_`��	�N�h�T=�r�	��qڈ�ў���M�Xu±�SI���[�ٷ�nK�����Ӫ�'������09Hp1m߆�x��o����)�]&29��3�Y�ZT��M��R.q��;<u]ס=�-�J�f�g,�ˠؔ#���=���;���02�}2�����	��Gx7�0����C�������:��,�_	+fR�N����&1f0�cx"@i�������͉خOj�:
���6� ���TD��7���	�Y
��$��v �9�p���N2S�w�	�a���h� o�T�8�;�P�.�{���8=��Ǯ|�����j#|n���׽���譼_lTz|\u�{�K1�c��\�dl��%�t7�u7��z�ʅ"��C51wE%�5���n�����f[��'K�e��v>��z��=9�W!6���V��wbw�3m����Q�2[����5����r�ڹ妄��<�qrpo�5]r���q�I����q���jN\��!�i�G���ؔ����ؼ�����
�MF�Q����۪�����(\����9���I��r�zo�rWFC�{;��&#\�ҳk\9I,����[�Г�g�;�;%`^���z#���m{�kw��SS�����߰�ˆ���S{^+�.1W2D�q��0�y*)V�L�m���NWz�SȧR���U=���v·���wC���|��N��6V�	P��!|���u'�����Y��neL>��;30/�"^�Iỡ����q�␘�Z�v�R�5���ajt��2�.����������U1Q�o�\:bWP_]�w�N��rg];��y�T���#��Y�Բ�oo"�TV^ƥ�o�}�7�T�,�n��g3�}fP	#�Z_tXn��K�b�U��鲲��[-֓]��L�ùz
 k6N+�X�
�gO(0���;��)G0�з&qge�]��)��6r�����8g��:e�UZ�V��53]�wl6�&�ja�噩�u��
Sp�<1<�	+fR:ʫ��s�� 6�{S��6E���+��o	o����O*�4(��4IZ�{�����^�n㉻]~�6m�����Oi�Ӱ����{��L����b��-���W���� �[u��ᰰw��5P�NUF�8��=5�sզ�y�c���F?t��u�Oj��n7r�|�luI�a��a���5�5����ڿ>����M�;���~��u�,�q��P]%cI߫�j�x��/4�J_��O�%_P��qUf,Ŷ�%B�M�
�ʶ�[��H�Ľ�d�
���\*4s9��NR~�����8�nv*"�FO.*o#{o[k=��d�B����xO�����V� �y?gmg؜e��1�g�.�\*L(;��t�c�ؑj�ڕ1��#R �y#�!���S��3���y��r�-;Zr��wu�����s�V� �L_QL��x��T u:1�R���
Zru�Ĺ�ܻ��.�� [�\_���Td��ҵ\iO.1���M�I6���*7�l�n�uKw�;+��B��-D���_I���矺���/-Y:�������$�ފ�qˡ:y�b|pSV㾞��wq{o�b9�F��a;�i��k���mC�U�OXcbB��L�����3#��u�fz{�^�{��N��yl��7�@��S���j�W6�8�Kr�j����-��t�-�h�r�u�{�'��N;;�;��Xw�>EN�C�Ӣ�1��+x7��b���5���޼@��̌}�ӛ��#�`el�*Gp��}���[��Ƅ�\�3���֞��/3�4�끸�tV�t�z�N�h���+�Y���omu��p�=��Q�	�;�p�DktW]E��}t����S>��X�j!��RV�p'K>�`|�[В���	f�����Il�6��T�����ҕ��It���?��,G�3��*���n&a.79\��#Ւk�`�m��|;������7.�;�����M�%jp�AbKRT������q~oW�/n�����/j룉{�籤J��5��w;Vokݮ&;-1pޮ�__MЭ�B�WU�Mn��;X7_��)U� �����������|LH�6���
F���%F���t���HV8&2[<Te�u��t���޽or��V�kP�����9hpe�|��7<w2VP^����d�t�Sв́�7XVoy%����M�]w��d���%��:��IwT�M!l��-kOsi5qŬz:�p�<��r���P�c��������MѬ۬jY��)=5�+|;6��.��غ٭��.B=�t���'��Ʈ�>wq��o�Oz��*ٛ]F9�̜j�em�7��!C����5�x.��)�-�P�:sz�n,�]�{���WP\Պģ������Ym���2�Mdn�>��{�����tN2��r�[\ܡ�� ��+��P������(�4�Dt��˾Te5S��V�[�1"bY|�jP;ƌ����:$fEd� �q�L�ЧG�'�&5�V��_U����+x6mmc//#Xع�����K1�g
�u	�
��B=�ᯝ,���Z���J��O&��[�%9�j���w����گgW��u�R��hE�훏�Lʾ<)x�O���k@�Ox
�P�d�wN��&5��������=k����&VMk�Z���n-��k���;7���g�\���&�VhZ଺��0q>��-��q��i��z�\s�����vt.��\��w�_�`ʍ�y^>9-_l��6�S�����8����ػ��޲��Zp�u(^ ��|w�(�"Q����C�=m��5M��y��%O�&)�{��kͤ������앁zT�o֫�y'�\o���T�#ym�۞��.��Hd�U�r�Q@���U�>��
a]��iJ�1�Y��|�
_pY�Ll��w���Io ���)t��ޢ�V�^%S����AxB�%ů��t�Q��Ne��ol�e�e�>v��[�l�u��Ű��'1�c��\���.� 8�u�i�ַ�J1��M�)	59�x��U���⳰s��;6�7�v(��B0�0<�IJ@;eo�GYC��?N�����׏φ�V����H�՘��SWY)�c�|;�G\�r�K��]1Kxԧ�Ϲ����l�u����K��Z媐�`1�+������N��&\�9;��@V�E��Q�Z9�v�GDs$��æ%�UZ񢩮�q<��-����]7�໕��noaաP��ד��p���GRQt�&�(�Յ��j�n��J�`��[�c���5!"}�hq�"�C�
�}�9
�~�U�*�_��[c��⡡��l9�p��gG�7c"�U�[��n��)��)Ի�qV�-��F�S�l-S6�������q�����ڝ�f�F��E��Xn��/-�+}fOL��ԍ7�7ze���#5��U���ʜ�q�c�z�V�Y 1*�K�y����rE�x��0!t�Sx2QCeWz
U}����C�����\�Ne�����N0����i�n�-셝@}�:o\��5�(��8�3���[�i�2@�W���˖?p��|��M,�B�Aؽ�sU5���v��aTQr�]����[�^Ñ�^T��I�n�q��U��{�S7��Mt}ku��j��㵰�Υ�P�v߶���e�&�.�b��wR��Z�ŗ��d���؛׭�(��.�̍��k�q�\���ƛɘ�L��:�T_%Y<��+UƔ��:�2�M;�o���0���x�ʃs0pj&+W+����wc&p��u4�劯P�ƹCt����� ��\*-5�����F{��Ъ������O�ೞ���z�-�t��Թ�H�t������u�s�m��>�R�5�]��S�=P��ʧ�DM�j���N�w�Y����
s�y�snoG,���G��7���2��L'�=��
YK`c�
%��[���K(�Ҕp�(d{1����t�O+�NoK�Gtw`�.1���\�Q�q3���6GU�m�6�{���8��9w�����l��k`��[��H�)�WSfoh�M�6���b̓t<���H�g%�U{��J�Y��i��޼�C��"�iR	l��.L��K�b� l�|���7�B2M�G>����#\heƮ��U�ۥw�s��e��ZF��574�7�v�#:�e�]��v��å������>۔:d��v5[�ej�u��u�}j�������<�;�l�#C�[#��wi���5��R��{�v5��$u�wSU�eJ0V���:��!��0�s]��L��j�r��G�'�.�˛2vqZ��Q��0q���K���)f�t�m����k�u�o!!��k�}��V~�)���8b��}�q�G�5,b.e���@2���\R�KkVv�V�]9�wDv*����NƩ]�PHA%Me���>�r��g������	��s�����_$��fȬ7\1��r��e�{�>�a�0b|��p��"u�L��6�\��c��c<r�++��./����U+ �N�6�n�T�֤���tF۾�-�0n�r�ioln�{��!B�۱��-�G`�M�tiڥ[�gm����#Wʸ���)��9L�?'�n�c��+�GG4�},)����)�N7[O8��Vm\}����/߳"��@�1 ;�Vi��C�ͣ�7����5^�'��:-��-��}�q�g���C��(m�e�`��Ž�v5���y�t��}B�gn3�]��w#��U2.�E��J;�@��f�.	p�]|�DJ��ğvgr�:v�X�b4/g��Q����ޕ��`��tU<�HB�O�C�G�w`��`�nɳX��Us�pH�ƾ�3�Q8r�d�whT�eU��gaOU��Ư��NS#�F���u��s<*�ev���ϛ�A.��m�������[Y�I��M+�JM�ٹ���f�b�cq��f�u[��_x0���6n���Ѣ��KvE�cY�� �:�o�[{�b������C0E}u��4�m�[��l]:��|ŵ�X�17���1Sm�v�wY���,��]ƸЗz1�2.����z�`��5��sY[��J�孃&ں����hm��y���v�C6I����t�����m�Ce\�{g��E	w��� �u�sGM��r7G�_��V�i�۔(�̬�y�ڛ�����.U��Ψ�ZJ}Հ'M�,��_=����K����[r�^9\S�z�mJ*VL�#��B�q>I&���4Gr���H�j��Ne�f�fM�o�(��3QTu�������ڰ��T ���ai2�dP�1$P�$+p�V1@PP�,�!�Xb"ͳt���k04�+%h�#�&ZI�S(���.X)3,1��"��H�1[�ưU*V�m�E"��,�VK�Ƣ��nf!�
�H:��I*�%@�B��a+�s)qne�V����-�
1Eq�-u���%�[C3YIP�3$������[)%d�J��ֲc4�Q,�Y1��+SL�3(%e�
�m����e�S,eV�eKl�ʶ�«�Y�u@� . fXV�#�\:n�	�Rt��Hi4�T�b�*A�"��eˎcB����1�$3-�+Ef3I�"�VJ�LCH6�.�˖��2���LH��̴����U���@�#��#�*
A�Z���`�ju�C@�
E5lh"{��<��翥��(G3el����{�-�����A��=2�����6-��8v]�u�n�;��Y哮Q�N���<<U�����bu��+FLb�7�y�_9�s����1�'�+����E��"}�p��|�Y��-U�����١z4��L���wc-�����q�t��`�VA[0*��W�ϭ��]�"��ĕY�Jߟe(�H-��q��ӸG׵����).�L�ǶT������B�^8\�Q;��[z�s��=���+X���,lju�F��Z�?#�;�yv{xw���3�־��w��o�y�z��R�.�''�[�uC3��5�%'%>һ���n;[瘷r�����9�:�����O���p��'%��Fz��ʽҫ/S{�x�G���{m�x�o�r�AoʿB
�:�_'�<���v�H��һybu-����{��tA]�q�M\�J�=v�ׯ��E��X_<��<B����՛۞S�+!��X�ST��e�h�x�F�����];]hnu��U����_͆Feu��e)=����9_���t��W�A8�=���T�n:��!)����el])��U�z�=΃��]�*m!+K�5,�c�;\+��M��;��\=�~M�N�h�؂�B��r&E)��-M�llq��o#z�E������OO7�>�o��m�v������ټ��]6�O)78�GIHHo���}Tc͉������ˇv�^P�^��;�����>�1��*:�u�О�U6{<�>����NiO�Ǘu���M��Ӗ�������kQ5=�P�*���,�[��9C[��<�s�놡��&9�V�J��UW��@��蛬|Ы����	n㘝��OY�yX��x���X֙��Xһg³Y|ܝJ�xs�@�n��%�6;b����+X������k����dfo
�]c�U������6;��I�;��WR��c�=���3�Z��h>��_K�x&;\O�-0�-���w9��Q��؃��G�$��x�1�X@[;�CJco�n�+;�Yr��M4%e]ݪ��v��\�Y����C����Ƴ��ܢQ���!���rb�]�R��s��j��O� �I�6��>:T����;�t�N�d��.�w�UUWG�w�N��|���w`������K]�X��8�W
��W�"4���ON��A뉛��>����м�<B��5p��M�9+���[ξ�v���<�-�*b��J��$kZ[:M��r߭���^A�f����l]��o��c�R�-��6�nz�к�!}W7�qJ�+j)c�6�w���l���_5^��]+U�O/vm�oj ��B;D�e����A0�_�.|�^.��OZ��ׅ"��خ5PNS�~OQ�F�Ϫ�<�=t�]����[ƛ;T6������c��������{KB����c|��1�pY��\���7=�ߑeOKy���U�{\֊�r��ъ�Ls$��Ë⒚��B��g:��M�Y�7��+AVoke����+��j��
�`���.���v9x��*��o�%��5� �R��-i�}�c�X+���㕸y]�����������P�r����W�q�Y�%�3�ok!2�+Fx(�U���ٝSU�ٴ6����t���E��{�Q�����{��3�9��:	^�2}����|��%O�y��b�\ 4Lc�����\9gj�Xδ�����\���6���i[Q�ۚ�d٣c>�B޵�})�)���F�S�o)�W���V����z��z�&#z�!f�X뢺�,7M\U˯[�\�Y=D�Q��ꦵ��z�8}|�����1�l�<9Q�^׃�8�K\�t�k�2Ἃ��i��h��Z�ڣ{[�縯2�O����PG�]�=Z}CO�w,������N����o��P���-��}��;#�U�,L \��a���s-����E�u�ʺUe�&��zf���\�2W6���K}
k�e���kާU�B�ȧ|��^�B��t�L���5q�UV��vg�)�J�z��rodr�Y%�F�u>H�*V*��Pv��r�.A�N�,H�	�(�K�J���o,��sq��Ƞ�5.W|ղe�_	+Nm�|2�W[��x�y��&�ӵ�u}�R��INꊏgL�V�H��o,���d�\��YZf�5��q��}�W�Q�F�߫T��C<��6�(n�@ѱ!�
b
b`r�EK��z^�b�1�++�7.T�O'��v?=�����C|x�B�󚮋�����}�ƥw��Է�zV��
��=Kh��s�k�qv�sؙS��φ1?2���x.��+��-�p��\C����T�}JÍ�[Ɍ��0�h�%�� �'YUZ2cͲ�F�n�~������8o^皞�<��<�p���%쎤wKh7���z�l��F�e�Pip��؝�O�q��jal9]=x�+8��%��e�6��v ��GvS�l-��q�	�8V+5���+��q�����)�R�j��0)4���{\�����\7���8ǵ3�����|*3�� ���ɛCιuf�Gk��L6Z�O�y�γ�Y���A�"��	��1��z�h�}� �7�e!|��y��h<�N�Lt� W���z�n�����\Wkc��G�٩$�/`��3m�u":N�םx���l�,�˜�9���uU��{�F�An�jٙ�K��_���DFG'ټ��f�b�;g�9-�vʬ6�5:ێ���Y��ʨ���r�p~��]T�w��Ôq�����ԺUeL`�ou�Y��9I,R(��|��%"��9��w��X�o9�VxK�|�i�ގ��s����޿9����{��tً��\�-A�qM�+\���}˙��W��j��:���qk.��M�t�XG�������'5[)���N1#�]�QI�s|�!���|s,���-���0���Xo�t}혁�p|#�W@]��b�[ħ���;{'O�X��Pʾ���:4.�:�pU]ׂ�О���U`\

E����ҕ��+{!�Ǝ+du��17Q5=�;l��&ۍ��K��<�UʵM��C�d8�8L��T�+؞V����Ȕk���`�$�c�f�9�C�*S�y�РWM����<d�A�	���Y۠3�
f��gk��ǹ�p�S/
6 �u�>����m�UaY�$"ћY��l��G\�"W� ��� �>��R�;������� �;;��ؿ=���j�4�6E���e��-�1;��C����el��&p����m�;V�/+���ݮ�S6�7��o	qM�ؤ�&�v����2���^pX��]AΒ��[��Z���n-8Z+\d-�}(m�]F��K���3��٣#=���To��/9�sԾ�zz��R��*w_$�Jz�u�E9��+�^B����ݲ�0۸R��%9��8OG�x��JƓ�T%�jy�Nx�<F/_��>9�a�Ga�"�Mo!��5�@֛��:UeƦ���;Եo��K�r��\;�����<ڝş	+yL?��}�\T����o�=M�xFL�����(`�-��ߪ�%Z��97����Bx�S+���GS�ء��m���eOW�5�=W�fةQP���c=|�b���/����g9�ƪ�N Z�NM�W��������0��S������T�,Z�r��}x��B�V���Ϣ��,ù� �p]x��m�f<�]*%����W�v���z��8YR���r�W,�����{�k�ԼǼ���fCi�'򪪾���bM�����#���^@ѱ!��Q�S�]�U����G��ff���=��&�Я�b��������o�ϼ���y�~i? y�����0�ĝD9����B9�dpեo=\)�������[�l�����s{�Х7���pI�����
��އ"��
�/�o��Lcy�do	n��WE§���黱�q�lGK�ӛ��!�Ѣ|Vs��t��Z��᡹k�k�ǀ�~�C�_)/�d��k�F��ò�ܥ�}��&�{�t�]���腆
���Pqa��Ѫ/!;�h��63��c�Jq{�\�\���1�魣uKo6&7-8�oW�>{{5��1[k�*ܧЃ����&Z�e�������/Rjz�����qU�^oǈR��{��q�$�G�R=�1��{ۥ���� ��NE{X�wQ��u�̧���[���3)�u9�M;�^�4��^n���/�Uª�#|[�*�����>��H�_�����ᛠEY�geF�<t`��#��ʎ8����UU}j�\��ɯ�@䭤d�:m)�\׽{������l�iҋ���|&��D�!y�R��o�-����^'��6�7�[���\�5fs׺:n���z�Amq�������yɿ~�y]!T �M�{U���7�<���Ϟ�S{�3:��;��˔�g��_9f����k���oZ{��毋�oB�|�7nƍ�f�0SU\�f]t$<�eI�J�6��1�lh9�'��OA�}S��.}0�Y1�uVTj���<�B�M!01���]��)o�[���2�ȇ�h�Y���֯trC�r�1�0ٞ⪵�.��)�-��͹� ����y��^��?e:�FEg�[���G>�eUh�N�`����g��tg^&3�ZZ�)fC����P�<� �9vU,�����o�o_�Ū�l��`����`��L�>�u��u�]�CX�(#z�#���Κ5f��s������S�H1�QĭW���`IX��8fboق�O�@��~[�Ԙ���ڻ�$ӿ)��tUb�5�u>�=[�c��[(��}�W�U|��y7=�W+���=w�v*#��st�,P�Ȃ�>ke�4����^������rjl|�F�R�l-��q��Ӆb���+�bQ���2���vj��t%����pqD������-�L�<8�iErי��>��ͧ�D�X��9ν�*�ۮ�S;=j����^I�rf�I���޸��S�*�U���9-�v��K5:ێ���i�^�����z��=R7�!ij;L_B�-*^7��+x��o-�O��z)
�Ex��������x�O�%��Z�L���C�(�h��7��tf�f�s��K�xS�m��oB뼅�&*�`(�]7�Q5�&���J������Qr�7�G���vm��'n�hܭ��;�{t�O^0ԛ�p*.J�p��tRzk���u�C�1��z����չ��WWwI���6omk��>����˚E�����Q �9kY��m�5�pğB��\���Gr���������5�L�x,�n����j���bY�Om7�e��Ԥbo@�WAR�9ZH�T��FkJ˷������n�F����E�=��Z�L�Ic�ś�fL����AVki&j^�z�k�" L7t�l�P汪h;��l�W7��Xdp��rꙮ�ޚ�:�\���SC/�ev�K8I�o�m��36#n�oΨ��J�9@��M���ٲ#:�[S.�9B�X�v���!�̶�wghv��s)���띘1_i��e�H\y�T�+�zn���o�kN,�fV�;�8c0����:
�t�*����`���0	�ڕ��T)&&�1�������8�/K��4ޜ3�:!��}�wDNl���/���f։�(��cb�D���B;J1Y{*�"���|#����[Ư��9�f垸f�[�ok(��0�s7����t�YiɮFV��Ll��2X�V�n��4��gV�K7Ld���pe�{�5��`qw NۺQ�J�҃����<�W����V�uj+�Umm1H��kfL���Wy�P���s]m��Z���-�����l+k�ڍQA���f�{2�T�;Y���Ƹ�Ʈ�`ő[Zd0e�V\��:X�}��ҷ�Ca{q���ҧ��g�!�U�{ĭ]��������H]�W�Z���곗�9�a�icJ׹Y����y\l�mZ!bf��pm�ۨ�&�7� VK��h6íN�ſg�E���M35��k�OM�r�e��wV1&���r"�z�fl�19w����fE�ۤ��:4��7�v�e�d���{��1��sk0Z���:��/rQU+u�v5���;�]vR:��O8�Q�n3��\N�/x��k��A��ث����0�Zvb�>�%9��*�	�v�,��w�e��i�2O��#R��G��� �Mn�^��G���H��,��Co���uMEe˵��n����YH�wd�b�M*�![�ܳ?��+�>7��%wȑ���K���q�.��Ɵ+&��[2���b�zC}��6v�9p�ΰ��6�r��n�&�3���*9\Q�Y�'�Q�� &j�7}{4=�l�t+�,i�Π�º賯e���$7&d)��O[xWc�f��N4r��3��|�Va킢�����y��]ڇ˲�uv�4�w��є��kZ�w�j&*&t��}�/��[���W�T�tɈ>��v��}��m��˲l�GnU�Ӱݡ�ʹIJ���:YގE�qm�*Mj�.,$���#�+��u䋍WI�6���`
�sA܅b���� �Ň�I�X�J�Kd���PĐ�L��'ڡ4�]SiY4ä1�&0UKH�Kl��b���T�BT1!�(LAB�L�\d���)��E��'V�T-�UH��)�����`�`�u� ��t�XJ���4���Ҷ!XT�J����&3
����%T���MLDAdU�H�%Lb�"
���u�ǧ5�

)��µ���R�E#h,�-��@Pnb�Z�
�ՐĚq�3Cm1Z�ft�4&��(��za��jW-Z��R����-LzʤFV��:hi�i]Z�j�j��CI�ud��(VM%�+*CL�f�Y�M8��4�9�(��`�E�Vf&�d�j����:[a���q���;9�6N�^���G.�j荋������7��`���޻�oX����.g���`�=�(�&5=_}_U}TjZ�|������tL連��p9��\���&6�y1%��U�q�}=��|����ϯ]�:4.�:bWG]�]{e0)El�W�}�jji�rp+�"��_ќ�z1`��c����ľ*�[�'����]��RN�WM��ϡpn�U���7��&9�V�����6�nz�6Dne���e�0�� N���~�T�{���y�gs5v *�T�6�k�*���ډW��ٴ�y��.+͎�N/�l�bŚsTn;�T�n��)�[tqϠ��un�j&3m���hf�ǳ &{��nV���ꏴÊ��C�����.�-��qKz-�m�s{H\X��7��}~~Q�|�/-X~p����+�-O�KW�*��f�X��U:����>���m5={�-#S��y�x���-�:�ֽۍ���K�ݞ�b^��7���z�;�03j��:C<�B�y������;Ӭ�cC�	�ǒ��<��F�Y�0��&������*�&�f^��Z�[S:�(�N����SC#�ke_2GAz�k��;>����e���Dz"#Ѱ�osn�������U��/ڛ�襻M�ݭ;�w���*��{b޷GAj\L�T^'����R�-��l��WfdQx�EH�����%ù�ʦTI��_%QsϊՁ;~����dd�$�x�ٻ���6��ex��P�q>�˅_5��������k2�ujdr�V�Y��ne?�%109p����G,e�k�Mn����S�z��[P�}S�lH]>t�Wg:��g�.�+�&��t�?�߱:[�e'NkEr���c�Z�~v���
�IKɾ��E5�u�U����Ku�ijOj;M��3��4��T)N'Qu�ᓉ��G��[�sU��7��[��)sP���.��p�2Շ�*��θ�6b�s����.���TKg_`��"���!\f%�]2ek'j�h�e\%��5�k �\Z������ǹqd+5�չ��f��e�W]��*o�+P[OO=wB�F�[Z��.��]3��l:S]O�y�����^���H���5o�[aE�1�-4��](�������Dz;R���������ƥ`XƱ����K�WV�ր�PTO#z���jp�%ne(H,�'��;�G�[u��&�z���M��kD����j�-u��v�^��v�\����|�g@}x���F5�q4�奁�.�ۭ�ژ�{���}�5xw�cL޹Ls���v'�{�Jߑk,�N��[�ȥ��!l	9nL>N�^�7�(f�������y+x�⧓O�$�L��;]�Ws8R/d�l�3�����FOB��9���2U�8�IFO=��v��*������НSL�;�d����Ќηl�̹O�a��`�:��ծCr�������RO�����Y���|�p4lH{>
3m+����L�I��1̿U��y8Ly7
��\>j�}3����NA�
�����[v���ɪ��hV	�#�o}1�-(�]����43�9F�w�n�Հ�W�Z�����7}X��
�/���<�zTh�&�x�y����vsW\��%��/��b���jᾥͽ������v3r��/�UUW��Ӥ��''>�C�B�����z��[���)����05)p��7�����C��|����|^��f�*n<'�給�}��g�ק�u��55�+=�p�A[>�N��"�d�w��D6��.�����o	O�1+*E��lϘڛ�^)n�Yof�"��������\���I�7]C�>��.��Н��Oi�Ӆ`f��El�K *)�cZ8l*�E���U�)6��o#{)��b��2a;�p�kg�����Q]5�*������u���հb���n/�����|�3G��~ǘ���Z���g��U�*�<�k��L7���=�Դq���`n��l�
��yA��5$��d7���R��v#���j���5���̟S��\O�/��U�ڞ���7�Ww���8���D��¡����-EWy�(���o9�+��lTu�y�%�y��g^�0̨hS5p��`���y��y��ΫW{�k
DTevK��23�U�`J��qj�Ek&A�%�98���;4�w(	��ݥE�%�G���{��z��s���{=O�k!��x�ox2q����q���}g�\�Y=a�o���I�'��O\Bx��$�4ɢ�	�I�:ְ� ��/���N�}�����D`��D�b"5'�6���=a�sz�|�0�3�3!�N>2�s��I�5�C�0�S��'l�O�6ʄ���v�dv����sy���m֮h�߹��}�,��93�',���!�'�tw@�N$�������d8�q7l8��C|�
��OP���C�&����	�o����w}k	GVq�#���ҍ���#�C�`��1��/0I�4̓�XMZm�̛eI��i8������l�_`q���:�2I��C�o%@�OXyU�z�ڮs�wa|g������Qcޡ�l8�d���'�G�i;�}�m*I�ݰ�&��O�6�ǧg���=�=^�>��{�"/o��;fx}w�|��������ϳ�IĬ:����LI5����&�R���h,R$�N�2VI���$�V�z��HO�Ǽ�{�c��>�yo�����������Z�@��d:泦I�Vo�<Ad�z<�'�+��B�m+&R$�&��V�L�	��҉�������y����ޡ���0>I��w�'̆{�*q��N��@�:d��{a8�a�����q:��xɉY���l�y���=}��=.�+�?ry�u�}�{���}���&Ӯ��I_���x�;�C�w�M2q���<�̒��OPz�ڒq�������C��öLJ�AϚ�%��� �{��,�#��y{�`x��&���$�'S^�;|I6��d�J���t��'{�q'���(�%Cl���̐;B�N;�����cYy�c]غC!v̛)qjܹSqGF��T��Ò���8����Lm�^zȷ���5�l�����H�o!*�u�]��l;��1k��˨��L���n�Ap�*�4hܴv_0�n�/(��:�+tk���~G�=�{�f�]�{/���{�'��2T�����*M���,2zɫ�mY̓��'����v�0;g̒�N��C�G��hq',�N���fuy��<���^�E�;J��)<C^���@�a�&=���*M�$�,�06���I>`xe'O��hN�L���"��=�;'�z3��9.�]�^^�����oHzɶC��	��6ʝ�I��;��4í�1��݀���&��Rv�P�2eL�I�9��{�>�9�^yϹ���	;d�8}Ld�3l�~�|��z��2q+}�	��zÿ��2z�G7��ԓL<N�x�I��I��E�:K�;�Z7�_<�ʡ�F���-'�H�`�G�F!�RM���wHx�̜N��2^���t�<��8���<��z���}��zÜ�i'i<�S�O2�k͞g�j�����^y�=��ΞBzͲr[�'Gz�8�Vz�q��������Y&�|��X3����d��C���'z����2��<z��O~���[��+��Z���}Ä{�#�z G�H$�c#��OP浒m	Y�d���a�'��&�q7�yd�c���c��h�@�Y�b�[������YG{��t�o�p��Ch��]��>@��6��i<z�Ʌ�d�f���>ABh��M�q+'S��q���vc�c�B�ڞ�\�r��+ކ,D�3�Cԛ~d99�J��'��vsy$2}�h�I8��i=eI�'�'w���8��tZz�l��dۥ{�f^���f/����=�"4G�p�=�M��a�IP�o�2{����a>g�ts��N��dēl8�I�=�'�m�R�
�6�����w����k�i*��@��=����xl�].�V%��fo+��Z7l�;*K93��9N]���@1|�"�vu��84��/�U�Q��jv�MкN���v`�%7yi*U{"�8'$�w.���i>S���T�MO��@���G�3�U_UT��{��_7�i�����|���V��'�>{N�,�Mu���LC>�By>�t�=J�[�'�1��y�4�PR���i9w��tl����{˼�n�$:a�'�|�RN$ѯ̓�d�u�I�':��z�����h����=x��N�́����:�����>���3ѻ?H���/w��ߣ�����������a�)0��R��2jg�'I>t�ԕ��08�����$,��*q��8ù�d�Џ!����P~�w������=�Û���7�����j��
��V2���5y�2O�:׹'�&�q��`xwa�	Y������'<�ϼ�:�u�z�.���OY;d99�P�OX=o�qXtsXv�2N3��d�%ed=`,��I�Xd�&��t�m�ֹ���$�;��q�漾w������w���y���5��<d�*}Շ�6�p���t��N�s �|��{̄Xx�G�öt�q���<d��'^ӌ��oi*DG�f=�"!�v����W�瑛��y��'�s�!�i�l��Ͱ2}�C�)'��3��A@�,<I�OR�����s�t�c��;dǴ%��{�G�p��X���ϫ��ꩭ��۝�'����RC���8�ğ3����gG�'hq:=�!��[�!�N2�:s	��z�;��!���Ƅ=�P�n�[[RYn����k><d�'���]�9l�a<f��|�і&�8���C�8��x�$���߲N�'�f��q'Xs̐���G�OӀ���1��>С(�n#�=�">=�XOY;��$��GWl�l�-'̓��ֲN0���T�2m�S�C�8���yd�a�57���I�|���a�����N�h|�$f��M��MOi~��uط) �,�P�����jS�p(��-z�,�cM�JSa��cJ�f�#���TQ2��Ҁu׋f�A�/1���7�I��z�ZY%�й�=�����ٜY�E������ ww��_;�Ϯ���|�����06��M���\��js�6��x����O\Bz���&2x^a>`��>ABh�<g>Aa�tRm��{���󯳳�ލ}�<���y�{y$퇬�(z�x�<̆�8����0>d�'��y�2��}���G�M�d�O�v�I��d�B���
�=�}�y�]��k:�Ϥ�ORp���̛N��m��`q�$�n�q��Cg<�P6�ߖ�́�	�y�NМ@�['�Y=d�hN!�M��^e�y�G�.�����{�"y"$�o�8��VN���2m��wI6��k��q�����6��w�䬓��Y'{��tɦ@��м�/GV���~��w�w�CHVO�Y�hN!�&�2���l�'an�|ɾ��'̛d����=L��<}I1��$��$g�ӣ��G��P���7Y��}*��B=�����L����'Y=Ab��O=/�VI��&���I�'�:-'̛I��w2����ѿ�=v�:��+殨�(v;���¾�C����'̨o�v��8���<d��H)=eC�a�&��Vh5�'d�u�I�'�|��N���vu�q��1���?;�F��z0{��}�{�G��Y����'�>�$�!��ö
I�����<ݜIRm�
�x��_sL�l��'a6������˧�����ϝwߜ�I+���2M�^{�8����T�'�;I�Y*���o�$���5���?S�J��w�$���IX2z��{��k�׽s��w���RB�N�Oud�J���ݜd�+3��q'���8����0
Ͳx���I�}̝�L���a�%I:�κ;�Y����̻d�-��4���.z�|{#{��n�ɥN!�I��T��Yb��}RfR�s ���Wî�����3GX=N�5'a㕃2r|'�`vt	Z��gj�W@e��?(�ʵ2_:ݽ�aF$��G���d$�܋ϣ��G����,Y<I�ўa&��M> �i8����I+*a�0>Ad��}�8��Nr��'���,"æ�]���[{�3nw�+�"ǣ�=B�����0�Oi�J��"���5z�O���&��ݐ�4���t�ɿp8�I5�;�|�Ĭ�|�u��r��6u�w���{�1'I;eNo���÷�I�:ݝ��l'�X'O��'̓����$5���8��;=�=CL�O���D|#ZL��2f���}�v�ކ=>{��'̨y��&�=��ܲ�z�g>��l��4��O'��'n�2O��q'��Ɍ� ������^T�:��������<f��v���oY��I�߿`q��N��8���<��������$��i�O\a:I;����`���� ҵ�U��z�P��gHm���M��5޲I����N�M��3!Ĝ|d;�08��M���8��sx{�$񓹺M���h�K�Y}�~�����3_G��p�����t�`��=C�O��u;�m'�>g]�O~����|�=̇�8��vs�+i<}C��0�K����[��k:�����5�O�M�d�MBx�2>�Y'�pϲN2Me6��M���i8��t����l��}`���G�cގ�|�cɭ�O�r��"m����VI���:d�N wl��(N3�N��a=I��Iĩ&�vÌ�`uݓ�M�q��ya>d�9�����M��?kì(�O�1􈏢���7��|� |�����LI5>�z�$�
C��q
ɴj�R<��OXu�䞥a6�e��8��������[�;z�	�ǉc�`NA<��;�5�*]�c9!"ч�6�mh����v}dJ^e�]_u�o|3����!<�
��H�w:�Z+���1�����Z�ԙ&6�Z�nMW��tk
`0{�`7�̂Rע�j]*�]�*m!+K��#��G�s������{�������{����=�$�3��q��5�2OR����8������8�d�+�ǡ���D>"#�nO�[
���e�|�N2N�u�|����a��;}N̡8�a��8�q'\� |�2x�g�g�'�:>���N'G���La5����!�":�h���lt����4{��}��CI=d��I<d�Y6�$�VORW�l8�ĝ�J���߻¦�8��7�!�� ���$�<a�5�h,'vp�:����s�=�w����LJ�s�����h�̞�j��$�2tk�'o�&�L�I_X�t�����N!:�xVi'P:��*d���o��d�����Ӽ��9��">Jc�{�Cé�%J�y�>@�6����>d���m�9�u�$�;��v�04wg̒�L���@����ϱ��y�|/{��Ci;`�s�d�d�+=��Rv���öt�7�vɏL'���%I���e���v�3�$�����	�5�	�i��+(}t���v|���~���=��1I5=�;C�N2�s	��6ʝ������{��l�L:�0�N��
N�( z����`O�o�}{�5Ͻ�u���������^p*c'�<gRLd�v��i�g~o�,'�[�!�'�:;��d��s�d�����sy<}I4é�;I�&��d
��Ĝ�ύ������ts����9boVO�z��x�$��]�!�'��<�2ɯ~��:d�w�ڇ8����@�O_P��C�Ozs�x�x��w�ɾ�#ξ��5����&�}���2,>d���d�@+=C�>`��w`x�̜N��I6���z��� �C��{Hl�2d௸h�T��_��35��F�Ԭ�{,a4���`��c�VB��=v��,_)�;K96�_w;�X��%$��:����\��Ea4����{%18��>R���c�,^Rٕ�$�X�*��F�Fmm���IV:�[�32�=�Hĳv�2��No�B���H�)�3��%ܻ�K�L��7tu�͡��B�gZ�kfv���N�A٣B��s��At��*���4qh�fa�-�2���Ҕ��	w�*B��ȳl�t�P�e�34��5u'W1i*t���K��Y�g��V��0�މ	���C�$�fmB�9�I伾j-�ѯFl�A���EQ4�qξBJq�\0�m�*lhXrk�뜮������UҮ�.�\L�'Q�q��u�(u�9�+899���*c����C��Sq�n�^m����K �t�).���eӒ.��9Ǡ�i�����u�K��E��[�=s���p�]c�2�P[��Z�7�����C�L��Z���v":%XF�.HY7ӑr�66zũ��ю�l��ۥ*.g\�6��u*3c�ڕj�4�J�ԾS�u5sd�R���<5ӆ��G5��Ù��Dd!q#)�v;��'m���S\��H��&���:�9��X�J�$;RL$Nh*�ku@�o���]1F����Hw�E�J��D6��y���z4��H��>��ǻ|↷�9���d�h����"�D�b�6s�p�nu�ͅE��Nk�X��w�}L����歷��;lv"�m��	����2ͺ�þŋ��ܚ�fس�a�J��(2��9y�Y�}&��^��l��nĕf�L%��y@UG�;-ڙ�O.�s����c����$1�꒺����,J�<� ����*���U���N�G�X� 9�j�+��W�b^��P�J���v�bƧ��t���x��;{D3��>9z���<>�$h��R�m�Fn�y]��hfT�X!̬7���hA�����e+��-^�>��㭢��v++���ZY��+%	���@'P�ZPŴ�tx�|�W;�N�D�wCKMu����ա먫[G53���Q	���ׁ��F���55�r�yP"��Q;l��S�[�u���E��	0�)�.ru��ܼ�)j� qj����s	nc�f#��1��!ѕ���]��V��ƌ�0��`�]k��!�����
5��e�=܁-l� ���$���N�p倨�N�� qԗi�ج�Hu�f]���N qt�[/7z|�Y� \n6�C�Q�R��`.\Y�����N���ޖb�;-f_�|s�/2fFz����uJ����Z�֫l�`�+!Y�C�L4��cRc�J��+��a�i�2�c�J�H��u��aR��V��bԆ�H��M8�]eQ$Ҧ�4��M0�&�gHt�4�֨�j��QJ�ht0��P1
:I
3:�CC]f"�\�Hc��LI�ul�L��Z�i�M=5
22*çN�X)��[�H=Si*WL�\�`�ZT�D�B��J�m��j9K՚C�hCbe�(�KV,�P�M�42�bۘ�E1�YEAˬ���j9`fl�fe3W�I�įIG���Z�0������������"�*��:�gN3�J�l�Kr�Q�C��"~�c(}��3Q��۽1��˒�7������rkg3_Z=W}'e�Q�����3H�7��=
*V���_�Dz"!Ugr
o�D`�B�ߞ�t��?I�!RVO�
v�I�s>�q�5��u�k�
J���6�d����M��̟8�yz@�M�S�r��n�
3��~yL�^�V3�[g����=�P�CfDz `�>����S����m��ve����m'�w5�1&���PY�6��d:O�P�j���T�bL{<�|�"��=�9�����{�~��]�Ld�*Ns���@ğ3�̬�M��!^Þ�4ϒz�T<��M$M��ۤ�
q��OY�0��єC�m1����A@����H�@W��P��E������8væv���c9>��N2�|O��I��a�6�Y1���8�I���1~}�^ξ޺�t�<\�݊�����C��[�����]2b�~��d���ȍ�=1Kz�\R�);��j�	c`��Sy�e��)�D}!�܂��tl烒4Oq�Ty�c�nB�ˮ�r����]��j	ٍ��,�F��h/��Y\*�p��y�Qa8�p�l�;�מ�[r���viJqO-;����VEEByROOY��&�4`��A�0_���"�Ku̬㻒&��W(�������*9So&��YD�����{���O��g����������_�9w�a��&b7-3|pPP-�(Ek�2������=91p���H����L��|r��T�x��2F4,�Q(Os.�;F�;+�|rP50��t�:V�fm�C�`;\v��a\�ыxb[��5��Ы1���9ނ���O]a'Ng֞ڎ�{�'����F�\μ	�����yԨ��J����u<�Syt��>���F��� vJ�����:�|��=�*9�N}{�0��8���[�h�2ߎ׆t��r��3͍pc�K'a��x�,`�n��8*�;������P����E�4n�B�vi��(-Nj5e�Ӭ2�V�8�������cc����B�
��hg�[����z�곃¶����ֲ�J<��D�U��5I��@�_l��{�.��^��_����K�:GP#bNAv�<E��j��+��V��S,,g��O��gzWfyp>���ȧ���3���n����vp�ތ�A�u��H[�<3r�(�,1gd�T��5+35�ڋRo(C���\*S��^T.5i�ȴ�9��c)�LWH�W�q9Isp�o/r�H���\H���'	C�N��̙�>Գf���f�J�!�Q�	�wat�q�A֞'i��C��.���4;�(vɔ�ۇ��PJ�z�R{�^@z�,{���J�;�y�Zl	�"^kc�����6@0�8E�����v9e
y�=7�m��)�ʋ��l��s[���� �4L�qѱk����d`]��eN��m��`ی�۽��^���l��/�W�UR�9���+�#*�g�7:N�=��p�n`TB q$vt.��Κ�`Y�r�ݭx/t��W{����;AA��,;(!ZU!�N�A��bQ5�:$�T+�U�c���A��Z�p+�W
�0�sC�x�
/6&�@A�s>ab��N��)I�/I�w�_�v���m|u�[踚S�1}m��%�l�9	�E������:mWx�`���x;v ~[$m�����b���\Q�b��I�Q1����a!QJ �xf�3�ܒ�$*�O�v�l���9����"���,^9X~2͊��@׸&�*��i�u�L���#���k�L���6]P���������]����Z�9��,=u#��|����/����}S�.p��is)x>B/c*�1�!�,������i�7�dl�=zg��T��s�1P�����[n�p���QQg8��4#n�g5Gz�C�-S�q�YU��4���.�nX��tƋ��z4������mm�`�Ea�(%�u���k�wb����4r+7c��P�����WR�O
�����Ju�e8�u��}��:�g?�	�y������b#*ܷ&�e�ݺ�Ҁ�J�vh����i��1��B��/e,'��ވ��w�Bb�l���
�0�I@	��0j�"�*���
�HM�z���^�j�!x�R,EGN,�]`I��,P��P�s�=+��N�q�����&L�=�S`\�=�L�YW:��.���r	|!񸂢xT�d�}�-O�'U���� ��.��4s}��n+�r�b��.��ЕZ|N��Q�U���yґUp��M�����"�?d��
�ERTź��n �0�@ O9<	N�]���`�b���K\���Pd���i��׷P�oK\3
�\+�`ڪ�_���,gL�t�r���x�<2���.+����&�A(D��l�26:!O��T_�b�-N�mC����V�,p���`uG���-��|umV�F)�7�ˁ��;=���un������V04k|:�%���6�?������A��|��&�b�N<i���+��*ʀZ둦�<��,9���oҧ�0 C(��/)�U0oH�7)���ɚ����;�B)-e�q��j��aZ#�4)�{����F	��n�$�Xbp��7�Gț �b���V�(;;VP�o��7n������2��������c��d��j�=��*��Aa��2��ҡ��=�.��>lU֓g>]ZwR�P�)�Z{K���@uC�슿'[;1hސ���v�@��Μ�[y�W�7>�o���0�_�1��Y/����	�}9ƇnmH�1�8%#'L��З-�a�fT��s*��VT�1�XD�x��S� ƻ��sm0���6��{гz����\ՃeP<0:�~tꖪ�V9�ȎF���_����A|vT�T�����l��nk[���?1vr�+�h��Gh,<)S87L�ڮ��v�����Q��GJ�&�xc��Je:�r��P�N� ��Q1��JD����h+���цش�7�������\Z�!�A�+6_A��;I��5FW<����>��\�yi���@z��*�Zᮧ==�=�u�~�B�v��\#@�Н�:(lv��SL�#:���baTS�LQs�@\]�m1饽r.���j��W:�| h��{q�&b�pS3[�U��`4���6�)#�E>5
����1YFaQ��,�7n��]뎕��18:	�w���I������{ �eV�u�)u�z�R��Z�_l]�4(3��\�}LRo����Ս[����&��`u�j
����fQ�m��$�T">
�w��jțe�;�̆�Q��W�}��=zywU��n��i���0�\>CG�y�E���/�����Bc�m�ir��Cc��9'���W/M�ȨN�I�,�&��
&�F��`����N��	�C�����ڒ3�p~�L�5$F�Q���<���p���|7Ch{�Y�.y�(s��ǃruB����k�	��ٸゃ�pؔ"�\���]����Ls%\�aU���+�����f����G��ϥ;)@���;p2Ї�`C�B@��e7��U�T�mI���XX6|-ϗGNQW�c��Ob�M�:�ؾ�W׶�Ov�	�70��%:$W�䉌�D�>2�˃�����]�i:gy�w�������Iz�K0�_�H����oyn�C׫�5��~U��yU��Fx�Q����7C$GlI�Pf��Z�u�k���d�{<�Z��Y�W�F��!F���[�fJ�`��I��3j6�4.�ma����e�P����ۧ�o�a���ٞ�\'�"Ɍv�[d1���=39m�] ��L�/;x���V�l8��B���7��7�j&o���RгגǴr�dƦ��z�bt�FfS:����e���S��z�Sv���vP�����=�C2���R��@H��1u���r��/�UWԇ�i�o��YS�G�)��ĺ�O���	�pb���O�N��M�䡩[�ꁀ��jټ�<\�L be�QQ�q7XYyP�է�"Ә�n	�܍
�Z����l*�"�z��rGExp����%y9�1�KY���B�o$f�s�َn��~;^vat뱵A��;N����\3Z9���J�n�j�S������5�c�9�1�S>�u���Ș}��y8��+H�P�s'�r��qf.DR���+3z�B���'xK ��TX�5 >S�8�bQ5t'�͛Y���|�;Tc��%��u��	ޓE��6&�E�ڇU�* �D�Qi�GV��I����Hю���ʅE�j`��l���.d��N@α��E��I�ӱ�L��~*�0-��D��r�6�X`���QQQ���	�O��9��P����݂}[҅�[�#u���ȍ�P�g%����L����}ƒ����MW��U�f�CVɩ}v:Ý�ޜz/ۉ�kǏ�����$H*�k�TPN�p��p�t9�_(w�F�ůP�h��N��=6Ӌ�|�&U�?��ȕ>�ːD���|��Ǖ&Ww[�,�QN5���8g�9�j\��R`�u�%#'�on*�(���e�T�yph�>緕�q�1�s޽�"�vFh�iW��[$sݮ�NPWgLTa����'PB1�zZ����C�V疗N�FG@��������U;;��^b�:cwb����h����Q�F�,�*��E���_��A��Dκp.0��*������3e�`��1����gt��a�M(yuۻ��#�
�0�zJ L	�Qg�WUW��J�������s���CF���;��;e���;��#<TJ�s��q"85r����ܸ�#�v���ɵ(��][����!a���M��8H�a�xT�d�}�b��N�g2:'�m���Woh�1��R��7J�)�f�{0D�빁��� ���V�Y�R6D��S�����8�P�e��肆�T�0槁Ұ��0 �O�T���+xNV�UZH9ՄP0Q�1����.}{~2��K[5���s��n�xUȸp�%a�v6�_��[�f���%����w�l���4~�B�t��6����: L�t�344��;�f�~��X�K5
5�_�r�7�π���f��9rb��¶]�QM��*<��2�T��`;k��|a���}UC�$�8R~��S,l*�By����'Go
�ɧ��u�m��:��WW{�ǟď}�S�>�m�x}�����|#�x5���0�<�rnGs ��������ِ���N�C&+�N2DP�h�9<*\��8���z��=�7RT�H+6��eCۢ�q�F���68j��3�������u0f"��T�=I�f7������b,�\�#������@u>�ȫN�va[#aB�xaA�&�
ތ֌�C��bDd����Ż��p4W�eM�=�m�'X6�jcn[��f^������4�r�^���Lf9��J��eW��*��N�o.ԡc��V�pQ�i�����ь�9SV��^U�R�\��w��S���:/����a���D��xS�xn{��{nX�����ˣ�|#k�5���<#���Q��P.��=
k����)��S��szp0�Ԯ�B��{ę(S��l�z��9�R��WH�a�ᜓU�� �4���<��'
U�F��v��|z-�}Tb�m��Q�p(��1�2\ru�2�8�b�=���q>x:��)\*wn���Q�!�˒s�j ���#�M�-��/BU|b�M�����_`Q��/������Mɼ��Oк|�.P��O��$>([�+zZ1��ðt��PK�)[�y,ؑz�哝J&+�"o����C�-W+ܝr8�m=�&-u\�3���6/D�B}���NT�@8��nE*�`#�sĮ/3i�LR޹JX�N�8�+�7�����.��t.���h��^�)P�ZH������kfB뇝ou�6f���tOocR��î���*6d�=�(zG&v\�w:N�A�Orj�[��A�&��jQ��p�mB�G`t+�����D7�I�qd�5.x!��r2�����N�6/3D�e�RGi�7��T5$F�^�Lm���~���|7���.�6k���bY�1l���s�u�n8��[bP�dȄ��<�gg&&:�i{s���Wofo�D�g�Q�����G^�ϥ
����v�`zP�q�����_gONt|��=:E�n[Vef�g`<:�I�P�ܕ`ų�5���T�9�~�'��]{)�<'I'�C�.���aʔ�zr�|>�J؝d�#va�s��G+���ݚ�Y����U��N�P�7`���]�,q�P��!YnI�,�반�\���W��8a[�Nr<\Aǔ��{=�/��ͨfoG��[:�k;1S.���]]2��k@�������
jE��
��mu�O�Ǳ��i+Wl�X�������M�ڱ}�&�Vm��b��TΔyַ`T�;72ks2�>��ڵS3c��nN��\%=�ڴ��=��2v��94\9Mg7��y��q���1����S�1mٻW�>�=]��d�QX�E��K�5s�� e� �qC��4�*Ò�i��q1���ܗ��� �uv������,�n�FL��N�6��uff�\MӖ��]��L��/.�e��d�Ov�`��`]Ѭ��+�t2Ͳ�o{�*�B*7S���ޥ��]|	�Ml�hȖ��x�eZ̚2-[����9�d��	C>��+���pW��Ui��8�&vz�)��N��2�ՃΥG�Xy9�����e
���]\� h(w��Voeީ*H�%mм��R8T�A{֯vc�;]IKzU��gS�Ã�Ae�j�N�+ı�{L۾����"��W[���;�A���;^ՐÐjŽp�CwJͺ� ���n�&��ΞlL�����i|�rĊ&����f�/va6}�-y�p�
로[e�@��%SA�@,N|�秾�\�Q 3��I9ך�],i��2w^(��@-�D���hĩ �Ak�o�G�&�8/�:���%�)�c���=Ȓ8��;٧t�7�U���2u]Q�.K_ҦĶolQ$I!q]wk)�Y��$ו�u�˅�o!��܋�NS"�ۏ#Y���[��5���ս��+_Sa��h�+��&|����26��Y� o���@qN���Q&���9X4�32����jN�PS�&%�9[;��5C ��C�}���L����8���nIxM��k��r�\1���7	��kދ�$jR�����kt��	�����y�u+�R�xҭ��!TՃ�]�d%�'{~�Us�`/��v���uI�3�mA��m��-Su�R�.R/�I���qD��w�Vk��v�BY� ����+V��W�%�Ԓc�WG�PKs��Lλ��'&_;�IG��:]��9vf8�s����C�s�	�**gA5ݸ�/l��P%�O�\%�4i����>�{+v���%ڮT&��J$�b�_ٵ(.�&@�Ά���� 9�$����Fa��䣸nM��qf�$z�I:�e>_E�sD�X�G3:�ᦱʾ|m�C�|e��
�q�d���u`(iX�t�I��3��j2��R[q/T�1L[`��"
M5PRV�Q�ԧT*Dd�
Tt�,� ,��b�E���kkV"�1%AVE�f���s(,Y��j(cX
�`�������E*���WV
)I*c�2�YI[TXE�h
¡S$�Ȏ3Ya���X�ܦ$ET`��uV��
�L��LuJ%��)�baY�ɡ�+*��� �UV+���-ek���Y+��n�ՐЈ�E���m��%��IR�T"/I4���2����J�ejVУK,E1&Fe��Q���d�`e-Tm���f2�U�s,1����V,2��Xb`�������	��Q�~k����	�����]�X����y��f!�:V�>ѻ&�B/V[���բ��.ܚL;(������tы[.:���������xH���Yȉr�.����O�F
�Y˧f���+�<Ӗ�Qn
E�U����xm!H��S��2��n�n+����qTڅ*�I��$`����Wc3U7�ᬾ��sM-��(�J������gy��9[�<bA�w��+N@x�{T�q(-�(<-�z�+ַ#'�����Ҟ��7�'
3Q�Y����@��(��<���A�'Q���t���<3q;`��ݙ*���
f����<"B !2��������hk�ܿOe8�V�/
��iE�f�ts�J���wr�$tW�a@����ʠ���%�WO�P�gt�>0l�s���D��I�N�<�MBٙ��Y=���ġQF8!��wX��v6�epќx�9��1J�3nt��YN�=��4�H�GB���5}rA�"6S��h�S[��4W�/Ac7���N�+�!�s�ts�3�L)O�;�l\z�e(F�kI�6��r���v�e��
����L�>� Ug��Wڑ�������Y��Ɠ68��e�X�;5ɻ�uŴ��HM���Ȍq�c�h�\k]��L�L�[��s�-\��G��rRz�9:>5U~�]%�00�0�;zM�<ؚ6�W�Us9o��{�vG&�]<��G-�ptv���Ҝ������o��<w�7>]`Qe�sӛ�w{�_��ΈqP
����,Z��%Jfx�|	;}J�H�3v��u�,pqi�@�ƚ����;�����F?��Eo���/��r�'�5��3u]�Cy���`�u%���W\�:�ᢦ&ܠ��*w���W�S��2w[�(;��8�ol�H斶�Od����G���Wݑ�xMG7�g@��U>2P2�"�4�p����u�*:cwm_�m�@�u��c�/5Jb�8�!xY,`!���T�(:ʨ�q�J���06��ۊf=�c9�4uo���4z�{&�Dc��T3d� �	���ȫ���+��
&&gJN�Vj��4G$�8�׍;b�C	�wBFAQ(TK�L�����e�y��(��{��'6��wy�L�:�}�z�?�7	��|-'�߫���-��Ć�Z[==��}x�o_��u�z��+]�'t=7;8X\��:N#1|"Ī�roz�kO�5Rf�*i���d�Kw���7�� ��
�X�ДS�~��꤭�/8�7M��5�!|�D=���|&%7wL��C��D�,������k[vk:��Br�̘C���	�/�ai��D�N�	����NE�U�C3��[�J]�p���D�,E ���A�7��JXp�끿�b� �v:��\;��%�5$�\D��E�����0�״��s�ۃ(N��ų
�Z����#=�Cv� ���YI՛��>�00 ����!<�Ď7=���B7��g#�V4�*��i�S��k6k���f�K��ø=�
�(enV���Oa��V�:���ҿBI�5�n+�um���T��3^�:�%�yP1�6�5�,��z�ۭ������˽D`o��=��{*���r4�yw�G�^�,��q*}qW[����ky��C�`�Ru���@�[�ǭ=���:��q��Ç(�)�������L�]«�U��2���ʩ鎽C���e_�����c�Hx���x�q�|��ʳ޵�R{����7�*N)5�Wp�t�koxc9�Q���Ii��sq-��왞K� V�ۺ�J�RԆ�.��5��j�Zs�w�>�F�Qq�]y�嗹]'0>tp�s�JdVJr+���[~������+���2���ʥ�c+���ٍ4���'����5�5��{�Pz��M�~�Z4\%��h읷::7)�0��E��&Dr2U�T��B���{��:��8iSӐ�6{N[u���"Q��q�Bd�=,C|p��0�{R&������W^�+��OgY��(0ƕ�\0�'l�EG�VѭO�׀g(�Gw�6�9m@s�É�|�.P��O� >('�V��S��I�]5���u����F��f�b`��`5<N�#0��b�r����ܵ�Z.,m��<�}�2�I���P��S��=fQ=��u����6!/�r��k�c��܆��k��{D	e�
��������iu�-�(Ml������_�M�K|�
�Jq.z�g���w|��<� ����%Q�wv��Ȫ�2�.Tn�P�����\C��J�@�r�ߝdT7rI���z%� $ �#�΁Xh[^���h"m�sU�m�]�����'yh��L���˶���i�N<вh*���l���kw�����x��R�L�^6E����W��wE�uuJz���_^���i#�I۟e�#�:���ؾ���/�#P��EOƱI
�f��Z$F��Lk����h�������搷ֺx6��r/oHmX�5,���ʉU�=�=C!�(F��'�a�xIѣ�n������{��v���-W��G\'��}>>vR�����:カzEތ4��A$���g^^�gp� ���=p��`>ڝO�lWx*��yV0_n���%���[ӄ�Nu%7ϧ���e��H������B�;4��;�v.�����<<lH���ㆢ�O%���0�g�1��9�Le]SG���C23��OkI+7���Cs���<u+��������&��m-�܈1�cEY�<sv0Ȍ�Ƈ.���0�3.D����(<���PW�Pxsͺ|Uc:"W]���3�z1d�i�����ԫ�T�EzT�k�y�(>��81}.�z�K$����Z�ףR.:r�8'���t��_�  SyW~��̘\z�e��a��ܿ,�� �r���<�W8�x"��A2�`}*�/ $��[����0\l�-c����KAR�*a�k��}Z L��mnE��f¬�����)��i�ӽ��]rJ�M�)�=�ZM-8�){o��W/�Dz!t�X��9^�Y��bc+����J�Q�.H��q"|z_d��3�Y��H,�疊��?Pԩ�WVbƄr��%��QKj�GOx!�0P�1�^���W��=�cB��n�3�Fs�,<+=2��)�0��ca�V�|�*��8�J�{	^�Ҷ��.l'��}�v��u�0G+w�P���,;(!Zn��H��c�`JHT��KfgIrlIuP�eIC��È��<�ޓE��lM��}�AA���^^�ܽ�h":��1_Q��\M*���U6p�CP��m�N���L��k&^��3�3�q�3Č{�\2�X�:N��⍳VX$����]�����}��7�EC����`A5�O.�Xxck�6�8]�r�:XF��TWUrbosbn���-ڤ��l��3�F4O���U�Q�z�犟o�ș���«��k-)��)dN�A�s�m{��$[ݮ�NPA_Lnɘ�=b6 X7�,�2�2*V��ǥ�"ӝ��]�&_��=\W��������r��m\��v *�p,�tv������C,(!d�Go6�*�f�f�:ۜfޑ�h�]��4���˃��6�g\�8��()���]q�r����d�ds���U%]'��~,�F>���U$o�d(gZЪ���u�9c3�_�����8� �m7�^�ٓ0��7��D�P��y�	DK�̧͜%�쮼�̔T4�9�َ����V5��p�r�oFBRF��0�!�PF���Ȯ�UC��VZ.�T��Q�l�=:���:B��B��v�\tz�K��uv���3:@����r���CG?Z}��>R��L\>	��gI|!񸂢xwF�"wa@=\y�G-�Y�����2&�[\&T��+l��=;dT%i�;C�y�{:b-_-��]`phL*�H�%��(:���T�1p�끲���aF�@m*�䵨w[�  ғ����&'��¿^���n�BczXbمG ��]&n�e�N�lN^��;3p80���<Nze��P�����rr0��߉B��|�"�+�Pipھ-���p��y��1~S�$�=��e�!u�Z;".Y�&������椏W���/hz�s=Q+�|�,/d6���r�_wu�^�(�QyL���1X�Ow���Y�o	��黽���;����-� �"-���Ⱥ;`Te&N#7���W�^�Vs�)R�������.����O[|ؚ��U�Gp�p/����i���c5���d��DT�Ί-�:�(0��mI�Uw88W���0��W����ܐ��#M'�qp�f�K'��4$I�Wޅ*�K�6.[�RE�{�@�-�c��'��^}��]�5]�<+�^���n�bj�����<6��2KF��XSͨp4Tv�d�5�+j�;XĖ>��yS��R�2�P��^4o#x�Q5j�θ5m�	B�ǟ�2����H<G���b�C3��K HsEZ�bǫ�ǂ}�b.y`�@���ߝ9�\�N�:�e�kMf�(����X���z[����ާ�<�6{NE�^��%�� Zj�.�����[��bY��׏3w��6t4n2���+f��u�Y��mJ� �z�ę�l� rא��z�]J��G�b��ϯ���$:��>, ����[Ӟjb`7s��u�2�5��a��'� ���`2Ɂ�x��R�e�%�U��Ny �)$qu\�{Xe|��3�D��h�J�9 (�[�VN���lJ}n�#*w[KE�A�d��e�}k3�wk�Tc6�u��VuZup��#��$/��$��}ܦ�/ZQYKk�LWJ���ӫ{R��B٥r�3"�[�����J
����U\���h^Luz�q0�9�/26���޹�霞N��_o%���G\ek�'��Fho�t+�*��ߴ��U�&�b[�`\��N��m�ԑ5�9�>�.T�8�� ��P��0'���=c�K�Y�^oW�2����ZJz�K�a�Lo0�+=��n�**�$�O^�<r�Q��q�Һ�\^�n��:K�C�ل'�i��RDh���YW=m}jܡ���Wd���\�V/#;���P]������L1���bC��<!F�.B'xT�9*�War�^�g�,9N;`��r����P�Ѻ.�X�{)@��t�_I�iT3�F�n� �u�^�q@��޶�片hK}g>��jsâqG��ȶ��J��U���i�J8}ԉ��:����E>Zw9.��.b~?��tN!J���7�o"~�����i��w�Oq��EƘ�f�� �d<��5�����Km6`�sṺ$˘�EH�M(������LUj��So�=+Eoʖ)�{�{�t�g�F�I.�����?;�S�QV�F���ӑ�l7�s}�Hא�su�q��:X�I�2�R�P��OZ�u(Ƣ�W�_*�����LC��6�uW.��s^������cY}��nci���c4Ɖ���|��7���4�.��K�ru�8�׶��P[�Pxq�O�ۘcO�7��<��nW�{�>���5Tz�uK�*%K&�,�*�i�pc���
���d�Si����hv�r�(�,1gd�X������<Oaae�T.0�FC1\�����r�[�1�d�ƕܣ�\��@��{��\H����%��6�|��֭[��+)g���52���ot�TBک�Qœ�^X�����q�I�5D��)�N��r&Xu
w�R�Lź��o��C��\@�M�U����ݽ��v\����'Fa��2��,0��B�b��
*P�u�r79�dp�OF����\Em9(P��1L:��	ޓE��lM�Ћ�����9���^^��o����G-O���:�e�j`���l[�����m^k@��b��%h1u�ʻ��:#:�P��D�:7\AU\:����8n�6��m��<�l5�àU����i|��շ9���g6d�[\"S8�lQ���:�UN�t��+m��!����,tͨ�Z̳��`x���D]a_G������wO镝���:��wU]��:���uE�
�{���)�����Po���|��]��H���d�«#�/�ձg$AW�%k�W*ܹYl��/�xd�)�g���Ջ�vG��aq���w���.�c fjɥ�N
%�UÌn�N}�b��E���o�f�7hl��c"t<4�.���'�J�n���"%�:�M�rf退�w�̱[���ЉX�H�ۘS�&T�wY��,�F%'�+�-�ω�U���ui��>t���N��Y��қwu+{�Yp�Fޑ��F�ys::}�G=7��F7Af�¥��=]�]w��}{�%I;�Ȅ��L�	ݜ��4����&Kx�� ��*.D]�#y��0)w:����sL���1�7��hCU/�u�I�������Z�Z��V���2�pݍtYvH�g>��r2�h�nA{�[���"v��G�{$�N E�~le��ή4Ӄ�iW'��v&��
�ˬ�R����4D�a^����x��gL0�\�;�͵Ɔ�J9β=�Z�q�:���gp����6�,.�:���K�#�۠20~�d����r;H�}ذ��K�X����J�ݎM�;�8 Lx��w�cZ���:�&�3���]�ϸNF�KN�Ρ� 1�)U����=i��r5�����^���4���<�^	G3G'W&ڬ\�UF�ǢF��|�ܕ��[���4P���/�Rg�u�W��"�p�G�w2��Z�3+UՐ����K�脊�;owƎS7��ɀ^&-��tɈdh����ޛ����i���*�xlgV/�F�e��Q���G2�J��[��j���ZF���+P��������)�^��\���»���!���#�WQY� M�N�*�
�s�4^�elя%n�ocT�m��[��(�dp��8M��gMQn^�nIg��>�r���B[�\����L��L=]LK\*��W�S�hI��%�T;���՗��rF�}
���5��} lh�'�l�%�]�F��
�MͧWgL����gm�ѳ�|�<:�U��vܡ)(����Q8 ��;�/�*L�a�ޝ��Y��ge��B��ZF�.��=�C[��<ĝ�y���\�qb=	\�l���]uLФc.u�����^��jG);T�n����gqW�\9�)5!�N�ێF��4�ܽW|�gHL�/k�W�V��  ����J�qq�br[1�	)��ci���X*�\����Jҹj�1�M7.aa�V
J�l�dr���d�j��T5h*��E�+PQB�V�I�ꖷ+�Db�K��J��5ՓYVe+mS)Q��h��$�,�
ܫSf�kZ��+A���m��&5��sU��j�0��[IQkD��iFDDTƥT31rb�aY�Vڕ���1�V*��P[J"\d�Q2���XUZ(#-��Q�QS��R����Qb�*i�X8�WT��Ĩ�EAn%F�Eը8�"�Քb��mc�X"��54�0�T* �b�"���-��+
��%E���Tj��	-*��"�FT���̡fZE��%Z�Ը��2�Q�EX�i%I-O� (QQ(�㔞��eN]%��ǐ����%�L�T(�u��ǳ�V�D]_N�g�c�]���Z5Ձ�<�QN��}T���?z���U������|#>�y��,ϖ-��J��X�*��T��;4�;=����%�ފ���V�`a5��aN�`xc�/`��%��;.γ���r
�2)�9�Zo��tGfR`�u�'��`^ɒ��a�>�gg�G9b�;Q]�wx_�qt}劉9E���C�3��s�mv�d��=�=	�
�Θ�F��c�1N5ٽH�٘H�>B-�Sf��P+�q���Je��μ�y�7iN��D�j𹥼64�H���Ƣ��<.�B�,������zj}���y����s7�������c��1�R�ɂ��+�*��G�`���+q���*N�k��5��Ce�s���Ѯ'ٷ	�E]!pN��fP�ED�R�˩Y���/b����m��.hK&�
V�d\#��=����bSwt��C�fpة�s���g2��t+nY4v|�[�!�Ko��*|��,;�DN��C��y�n��2,Q�ۭ���f����PثU�ը����ܔv �-/W���c��D��i��7�&m�Xuuo����;�M�L�u�v�9���h��c:���Kz��됁˻8�f�_${�r�Mܧr�k<�pQ��~z=���jo++���X�ڈ�\K��b,W��q�����QIS��v%J�xjk)��
b��Oj�¬�:�{:%��I��a��d�2��a��.�0T�.s��s�B��:�h2�[�z����#���c�p�Y���'=�������[]B�sy�F�,Cz*��Jht\)���XF�I�>����,o��oe��N��ܒm��ݣ�с�c6X��T�6O�N�C&@YD�d����r�b�N/.+{\����Ѥu��B��0��o\��#���#M'�qh�6J�K6M�Ts�թX4��ʟ]x�B}%*4�x�A��Pܱ��{I\��l0�R�H+Wz�)�[;1|E��,v`��Ѿ2�jک��������J��G���z��ޏM��oS,dĆo#x�V��냥m�	���fa���Mr���7:���s�b�9A����J�ho'��ɶtt0Z򣆴���c�.fڻ���>��H�:3���=j%M�y�Y���m�"�b��*�3c�8����
u2{�tP���!.:�}��⊆�f����K�A�"���]hi�ֺˈ�;�̮x=WÕ2���Ջ�=���ۣ5�#7��zUTf'ON3��MϺ
��@ɩ��PZ��Wsؗ8��X��{�{�7�����,&n2��l��S��c�e�ڕ�Y<Oae^Ft���@Tjo���ot?����JK�7�S�W(w)|Z�C��Vl�����є�%D��f�*k+&�,��D���b`�d��<N����G%���Zs���Ӕ�pd)��{���H��D޺�1a�$:1�������A+�͖<bc��L���ޔ����~�,W+��p�0�*#р�ȊB�ei#D��.�E���G�M�W��P���~5&����r��C����"��xL	�rG2����GU�[޽���[���_5#R�9E�PY�Df�0�:Vzy\�7�"���$�N��k�1��w�ed����8px�0W�!�+c�z6a�e���tr�6�e\8���&��h��T�t�n�k�G!h�G���K< ���D�ݶ�lJ�b�.z�t�va����R�n�1d�Z�d}���|�{ Y"Dhg�y}ۆ�WI�:]n�@��t���9�3�\<�)��]�6
sY����P!�O�fl}�>�
�"���J������f>�x��3Q������\��Շ�]��6{��c� ���S�9R�{���Q�.�vR�3+�_YX5�ıAŧ� 6t1Ǖ	�ƹ8z���`>ڝ�â Ժ-:��.��7U֢t�l~�T�l�:zX�����A��Fq!�3<�W�X�S����o4�il腄�#S���%y���5鍎����<)]>�*VzJT�5dkI�訖���4_�'CQ���UB�K{0Ʋ�g-�my����;��n����--
��1A�9F��PIp/�u��qT�WL���e��/Ou����9��L(N0�X��3��cY6TLuz](Qd�Y�U�U �:�g*7��9l%M29b�1,f�L"X���t�,D� Be1QG�q7XXzM^�=<ɐf�rHUe��m'r.��m�ʇ�DKJ�Q�.H�XP=�aOb��2&0X���f���t�%��r4�R޸��O�'s��f%E��n����n���<~ Nf���SW��8Q�`A:+ۛ{X����ZJ���Wd��h�C��i�;h˸����*�˸B���qp�s(�ꇳ{Z��:���v��o�����֚�a������'���7�.��F𺶚.��E��U��aܙA�)�0��c]ei7�*�슄��I���A٫�9.gw���}H�,K�uS�@A�ۃ(o�҂���yk,-��v��lgn�n�^ i�Ŀ����\�y*�S���d�7�#�]d#�p�q����`��Q���zFq9U#�k�})m�¢ɊF	�7:%�*�sٳM���r���W���b�	�E����S *�"6�!�X�?��J�gV�q��w��1�[�G�'�D�Doc�"i�P,�'�r. <1�Y#`!��g<;�<��wo=�K88�r¿GN
f���@v\�D'<�'!���������X�0|[u������;#$��up��L�w��]��"��wt��-!���;���&�L�zs+��"��TѺ2
�8ʽ3�Z�vw������ u.eʼ�"���|Q�=޾ۭ;��EE��^%(s���/�wi��-��ף�mS/Ufz&P�u�^2ox��7s�u�և1��0���P�į/tT2m��}�VVg
t͡�l6r�w�.ފ��G��J4.�w>����T�;�(���yhTT�3~��C�f ��R�%r���IQ0�5��q��_R�ؚ��u�0�	����t�dS�4\��щIW8*�2J F���]�byrN��_�T ����zs\O�m;b(�� �v��(��)��\���$n"�]���>s	�+�5�Z}�~F)�{$-0��M��@(H�������Q��T�D�>�V���t����>S���"�N5i�k�+��ژ̢z .
^�\J��"�AS�p���⃧���gVl�-�~���2��;f��� U�����΅G�Q���OM�>��2��Xu���o�]jpk� ��1�r�-�p��Ls��ץp�6:��VS:ml���C���u�c8���T��sC����Wũʒh!퀆��)k���fޝm�ԕ�����3�R�o
�ۓǡ9�T�q�$��H��D�}c.�m�#0hf�f����b$X�*7���p����S��q�4�q7[�6k����[m��E:m5�>�������#H�Rŕ�Tm �����^��5tt{�u���Y>���0���E�퀻�`����m86#��5�ep��o]ᖣǼ�t�ϥ�e���� n�Q�A�k���xa��}Td�5/+;A��#����]x�b}%�4T���A��P*�1��{K�HCR�ԭ˝�nPIu���0��_A|�@��b�}	�҇?������C fh�x�p���\������γ��H���q�(��__�pt�u�Ǵ��a��ΘW5����1��u�܎�/�Ԟ�ǂVE���������srZ�31n�c/5\h��dG3QJ�.#����iȶ��v^ ����#�[Ί߱�7=�n���ר5��Pph�eOpel¸�2�γ6Pa�]5�W�K�3�u+�Xٛ�K���xeg�:���1���'����;�o�C�\�zL���;NS�k֟e�tl
�W��b`�d�AJ���R�fm��]���vk�|��Y���s��Z 1�h���rb��H(u@bc�O\��d��A���@�#^-��k{���~��);��p�0�+خ�
�$D�CfI%�N3#q�&hT	�]nf%�I#�/�����Y�Y[K�=*`&�5�t�阄9a��
ZXD�t��Ɯշ��,II��z�E���g�����˗D�3�o�m`ΔV���\�5�j�$��ەu���Y۵nj�PY���9�T����3?W�B���5�ʱO�ô&{�]p��\�9���WK�`O9#�(z����z��n�ܻ��Mj;>���}=&7��yΕ�����YܒR�/g2�����x��I�`	80u/b�Dl��&�h��7)�������:�G��>��[��o�^�.�����0L�w[f���"0�u{ 
b��ݧ��
�r�ca rncY=rDm��]LpqF��,�nSw1������I�s�U׫̾�.�a�o��ؠAﭫ3<����v�'B�I�.�*-[�H��ɳ���65A��t�l�:zX���O	��U���(.HN����WJ�m�k-,��M#~ӢdȰ�S���%y䡺q��0��Li;Pr(̈́�sC�@kG����q��1�-`�;5�u����>^G'{)]nWulz��^GZN��
(R����sks2U�`^��{T�W�eq�PxQ�ts#X�{�ܒ��)�Vq�Q����R�ٶ�'8����`�)�6�_aX>�`� 5��o�r�7����ptFJ[�\(�֩Q)n]䰞𣔦wJ�`�_cS�@!(�0�؅�/���b��u���ٺ��)4��_UI�E�w�S<����)��|~��Ю�r�>�=JT�d׬�*��8M
�u�RV�07=L\-�7�(�,1gd騂X� ��b���$lK��[ƹEer���7�rڐӘ�m��{DCJ�Q�䎊�XT�tMu�˪^��;R`j�/�@�G��+��bf���o���� �#)E��zǀud�Tn��u�6�qs��c��D�$C ƇuP�;�(|��R���&�lT;�9���Y���rW����>��
N`�U:0W� ��BcxK ��K`�����=�̖+ڣ�s�:�Ŀ��:f�Ӓ�Řqy��
 9�K�����t������Ӫ�X�5�;%�S�����˖Lb���9��a�w��MWeA*�8�%��nO����,],��'\��fP�'O	٦�J��T8�߰)5W�G1��2EE{{�CMk�S���ō�rB�/V35�=�V��)�i�{G�E��T�*o�5�X신V�7��G���3�}+;ub�8���+jS��2Pi��s\���ǧ[�)q�V@�e[5�[�Gb���Id�$�v�s�?#�����*=Oe��l-����P�r�����i4[���p:X[
pS7pD����)�М�(�F4=�t�����-"�����7w����f&-J'(��\(+�3��s�ol�H斶�f��;�7����R²߃8�ٖ�f�X�V����:��7���UN���ۮE	���>�)%���7w֯�[n�p��1޳�@C0�P"}��*����i����/�E�a��iY�*��6鎗,`+r�$��u�^5�� l�0�J={ciC�׼ѫ�B��u�yUpZatiT�渟f�v�R�NX(H5�tmYF����=N,��X����@:�;��-�}p�=�XH�0�	����3�����V����`���PT��Z�2"a����oԩ���G4�}�sɜ��a}�8�Ws�K'�Q<'�X��UĢX�T���A�Cx�1��b���*L�6g_��l���^2` 9������xLLK��
�����s���������/*{*G�0~`ʱ��;�4��r�\�x�ȷ�LU�Ν7v�뢂�j�|����f[\�{[	��ԇ��A��޴�!۠Wn<d�g��q�W�������_��c]�L;N��P��U����=Ԟ3cmK&PM��k:�m·�N�Nv��}k2��p�V������O�Pǵ�5��
�]�U_v(�8]�4�V龫�8�m)X;R�]Ǆ�eA�Z@M�/WM�M���Y�a΂�dZ[ڵ�u���崎���j��o��o2�ju�G�u.f��IՔ�􉸥�����sU����Q^�&k�]�:���r�e�.���I�Cu�Ӱ���[˺˓}Y�G[��Ab�tMlݛ��C�t��J��|��ĝ�Jz��B���.�V��z�<���)\���.�Wk:�8�h�G6�kW���/�K��ј���\K9TM�(�KKNL)��f�.��sx ˬ��Ҩ�"��Z\����f ���ʚ�UwvJs:ޜ������UT}I*/���y�a�I�_!����F�v���Px`��PN��Z����h��}�-+_Jg k&��e�];��3�Gެ��b:�׎8\�.��˸p��;�]��Y)I]ղ�+��d�*%^
�h��'/��v�̗�td(!��u,C��/����i��g
2^V����o�P����'"]�Q��S;��Ɓ��ѩz{ciY�y�x�3����t�	��on�z�Pw>��f�U;��ͧ�TӇ��U�գ��qv�g'0�&��3�R�a�*���K#���)����WsG�t�%]�	m��T�/��P눁-l8�Oui�d��B�Xt+thwi����S��8H��ga�W	Ŗ�����f(���/r��j�kuu�X�ȧ�Y�8�b4�qEL�"�m�[x����J�1@��e�홖_qX�s�3�'�"eʷ2ogHw�|f�e�iی�F�Q����U)a��X��Wi����m�Q/�n1Lx�JJ���tߺt�s�w���d��:��t+"�/�^j�{]9�r�,�u�X-^���Gx"�A�� ���"m��'�QQk^W\�';әuwM���r����gr�b�{���w����P+U��
�;�c�M-B�G��X]u6����͕�4��Yׂ�m,W�	��]�>��hn��EK]�����!��X�r2�ReT�{(��*u����������� ����� ���E�����[˥A�41�d-�00^��:�t���I7JNL�6aZ$��H����6�7�%)�)��U4�.93qѪ?� x�� D�E�"T���Ֆc(�&8�Z��2ܡUG-E�mcdX��uKHTF�AT�F(����E�骰`��0*�����+EְӚ*�b�%����-FM2�%UQ-�j��f�+�*
.�c���U*��cb�5��H���SL�����AD�e���LfKLp�W-�R*��[�mUQu�Ȯ�I���0Ơ�ETlc�QUc�QaZ�E�r��*�EEe1UUF���`�*�ʪ#AmJ,Qm�Ŋ�(�uB�*����lVZV*�U4�V:J(:���EX[c�Ttܵ��1UHŌQDQQLs��9X�H�)d`�UDPXj�#�&�� ��T�;����P�=�nj=0�p�	O\L�gTb�:��B��Q5�A�׻�Y�L���+g�E9����n�Ou&�6�4GI�ס^[swC�Y�o��Z\1���O����e��6ҧ����I[������©���4:��XJr��C��
����Rz��[���e!�,��a���)b��S�m���~N�E3ta�à�&�=@�g��9��Ato�4`��¥M�Ys��D�����07��A��#L���)��1�e�����¾�ڸ~�ٯi�{	GՇ%�+M�w�A�anS]Y)�\����:���[tR�슴�gf��K�f�%�����1mN�Na�ޛ��=j���At�W���3�T��]^z��\��e�&�U��iuP�'_9+.u�T&��h�uwR���a�^�����6,g��ȱ�v��K{=�Gs1���ԫyNA��\��H�G�UB�����a��r-��x�������P9 ��_g��MV���s�>mu�p��<7����V�-<�f;6a�2�\�]�&аNOe���׽3���Ō�:�d��C��u��K��̈́g[���F�uZ�}���1�\Ƞy��hJyGz�e�ڳ��Pp��Ai*�FMl<V �/�6��L� �Õ��=׸��b�p̵fp'�E�d�����ӌ�9^��ZU/��xGa�0TLuD�P+�҃&��T\���T��$>(c���g���;����k�_�LL@N����
%�*&$�d��<N�)b2�2P���78����YuL�R+�C�]I�d5쑑k��ņ#@��`�U��=&�����L̸�Ξ�q9};�u�S�R޹JXN�8�B��X�R`ds�"|!��8\wby��\ovF���3�V�
�|juˮ,���z\�7�*�Q��AV���ǽ�;3s�9�<�.zO\\�;[,=�"3x:�~�J�@T^󬊉F��ez��
�^��ĉ z`w��+�F���h��f��L�RDh����z-0�s~�%�k�4�T?[Z����=��G�S5,�+��TJݞ��W��]vo�G5��XG��+���Fǳ�+���z�F�:6냪^��Fc>������Iw��1��C�+`En�4�!y�ؑQ�*p��;��1}{i��� �)�^;��������nU҄�U�,8a�Qg*6M�X㔪�`�W^���~(�K^m@F���}W�����$Y�ۏ��P�f�#�&�Qh�>�����O:g4�a�c{NO��@�޳r�Ns����=��f�-�p9��f3�k�ة�~nu9�����F�EZZ/:��i����fr����P:e!tFL�
�:�ᬲT<�7NCS�l<��զɂ�����$/.8��h��2��7�頣�#�]J�f�of���f�M�O��v�.'��Ihp��<�"*��P�,��:IuT�x�	z�{�2�V�A��T_MY�g1��g�l\�W]�p1}.L�Q1�ʁY3�o +Y��s|���K��1�6�C��:!����Q�a���t��_� !2���Y9Ƙoa�KSV�R�Y�U��"�̘\z��i�r6�LeC�"&Wr�d���XQ|.yddܡ�,]++�1H�0���w*4�M-ۥ)�����[�'�
����A��ֈ4*}oye�]���E'�z�pU4;�(vɔ;�7ʥ3�+I����(�'���Ů��k7�F����{�L�Zh�*��
�t`���(N��Owô�4H�0�������yEf�RW�1��+K�պ~Ph��$�5u��u�u莥:�Q�l5��7z�ؑ=�tKׂ	K+4�V��՚.�a\�乺��e�E��S�A$�JY���7��[�>��﨩s�hOi!�~�Q7@4�$��%RtLn�b�<6UU�[z���6z�rδ��\�����.;���(1���T9�)^k�:�o,�2[�Ƽ�A�|�˾�&;W\����ۓ�bWy������� �<��(�fl�fi63;}���z<��������%n(�޷ND�Q��a���E��0[X��{��pC�ֵ(��(,S�� t��!N
f����t{�)0s��3 ?AJł׵��cy��a�6����׆�\Ų�%��W

�L�|�ٰ���ZHR�$�+���xJo�oL�%( ��7�o&cY6c��h�Q��U�eh<��]aӊ�u�y���T���j��<t��ھۭ6��u��P#g](�1xM�&�u*��61ª��2����XiJ��.Wm��%$c��cʸ���{v�y��>��� �6�vZ.����Х��׉;b*�G����Oz	kvx�݃eb����e��&إ��=��W���i��F��˷y�h�*�~6Y��T&c�Ӈ��ky8��G&բ5-�,���0�y1;-e�cN��1}g����7�n7��U��8�݌ܨ�/�����Ko�rn�`��N
�>�' ��p!��d_���n�L_��V��ٮ�O/5�SY[ԋ� w�w��؉Rɢ��-�!���	��*|�-?��ɨ\6J�C�7��{w*�A��Z�='�%�P?�--p���˪ȩQ�1*ր�Б��Ki��U�p^u�� '����<xLzL*�xu�J"eM�;b��c+���
t���0�⫦�Ud!��G9<ML����[;I��B��us��MĎ9.#
HF�l�sC����y��1p�*I�{[|���p�IÑKn���V��,���,f�p'��sF�^����wog��F�7�6��D��03��D��+.p1X��+�oeCۢ�g�s�:n�5[����}[�%L6.��;fR��:�c�GÃC�{��X��U���4t�
���s�V�����c �9�o|�5�SڱeuA}�`�#$�o��5da�����+�ٵ��tQ�S�h�-�\�<�{���b�9�@��a�j��Hk�3)�źs*�l��`��Զ��'8Zm͢��b�V�FJl�{���i��waȳ�*�]�z�;�ǧ�J��K~�l6��N2���s�Q�4T{�o���.��k�m�z�����V:�*s��᜹�Vo4��F#��aj�F3��玘��U�E����nvME��ʣ
��
n.^�mCZ�N�*u.a�Qs�;����������a��rۯT�x�kJ�����pLVp��Ѩ-S%�<X��<7�<�Ȳ�R<�����c�.��U|�?6|5lX���@OYؓ"J���t�TOJ��)�C�ܩ�z���D]mK�{Eu4��Q���JޜJbCw0�i; �����*Y09Oh�-A���P��[z�B�3G6�)'\�D2Oh�]5'�F�LuE*�`�e�e�Gdwf4��t�qpKe�m1��-�~�,'SuTa,b�029�"�����X���A�غ"�x�6/�ռ�B��H՜ju�዗.�c����5���x�W���i�+�$���#�3���&'eIws��{e�$F�s�g�b�zb}2��Q61Gl<��3��WLo=�,���Z�u��I����-�`N�k���.d��{f4��M%��sQ��Yq{L�'�B���A��BkB���N�^Ӭ�/�{+���#����CYk����U��2V,葙�ܟ�[���^M.�����5Q<M3�\@у�*X8kؤ�Q�o,�}��qj�sU��r�� �sњ�u�;&�m���~.�����)�^`5�:�֫r�����BP��r'uA�rnc��Y7c�d�����q l.ԗ!w[���)@���n@zP�|��{6$W<��~�'_�Af@yi�*K~D���P��|����|:Ӄة�p��<r%�62��uME+J����Fpi�	��F�b�f��:!W�dXZ��oA�Y5%���-��B�ڵJw��ή�4��&��<��o�e=LuKX<)���_H.�9��>�qv.l�q����d�ɖ�#��}�U��r�T�V2��_��餺���&���B3v9�f�[�á:�@�VRR��CJ��Z�1�,���*��L��-�\�V�3҇kQ���Ẏ_K�.!��	�KN��X� �z ��q'�Bd���&�cQ@ػe��-<�8�:�,���t��7`l{lLkN[��;�]d��� ��ŀ"�!�r�wɧ�+78�ޘ%d�|�TU}���O�G.�k�D�#�#�%�����*��S�P>���QFE�Vy)��˕����o�Pyq��z->�	��W�	��{DD���.H衙JJ�iu�>)I�#>�!�D�r�' �9��i��[pjU=1~K*7p�*Ȥ�ʺ�1��;u�zU���l�z*c�AbP�A��J�r&Pu�x�B�L�wD �����I�+/n���
�m�
D$����%�!g�t`���PYF�`��Z�nw����\�Ԁ�y���.$���\�yPвtL��vdZ����Ѣ���4^��cjQ����x:=!�r9jR<5��u�u�oh�$���#��X��Y��q}m��%��7'��ro�E����$kϪ��/}4_��@���V�Uw*S3��xUM�J�P�8h��3��fj�D�'��\z�:y�bC��#`!²')���6%�#b;]]�I���2�}b+w�OZT
��۶�r�����eD�b���^�]�B��뽹Ԇ�S�������+_e�`�*wR�iھF������x���[��7غZ}�yS�;L�r�f��K�,cP�E[����y����κG����w�2r�`���{,@�4HX�u5�$�lٽvD?���9�0������z��t�<�Qn9�`���k��p����EgLTa����rp�˙h�
�en؊C�����v4�\�fpꕝȄ��<r�e*ѩ�|8u��9ƽ��d(�HW8�љ��B�5\��
�*���Ҳ��1c��LvEy�`��r`��F:�ëJ�"u=�2�UY}�T;�PrXL�<ʼ��+��
�4�zs\O�S� *�v�o�Z�c��K7�D����ıR�Ê�s�85�q����"���/I�Zj7�e{���^���@�_]�uK��ty}��Z=wJ�j}�B'���AݦܞW�y0�Myl�1k��	���N�|k���z|��@��є�Ga�욀B+��y� kV�xo�?	��Y�:�t |����,��O�gzn��zm��%�,[�pe	�ޖ��aQ�WLUY���� Ӊˇ{Ҷ�l~ysj���j*�95���J�&[;�E����9O�W+h�Ig�Щ�XK|�ex����� ����,+*Q�4 �y�&�z���bw/�Vx߱�X�v�a�D�t�B���}Ҧ�ф�%:=Dm�ۥ5<��5�����@ޥ�w=��jgWY+��qnT�|�R�(��}��M<�=���u,dV�h���=5`3����*��rx�Zuq2he��/2aĽ%B����U\: ը���<0/��yK=u�|�+�H��ʆ ��7�#�����=ׄf�H���J�l]a�;f}K���lpH�p��t]�ιrwruf�IjS��b�ᬤ=q�iq<�{{q\�'&�{ 1׆a	�Z,V"���}�Ⱥ�c�U6k����y��~��J�;+��K1e���Vw�QsV�w1����j�jCi��*��{v5����,2]�B1ҭ.��{s�B>��e2�)�L#6+G0Pb���+��
���&Dr5Ԯ��:zq�l���n����k%Ѷ�Q뷹�q�5Q�w�����
p�H�T�`��]�Sٵ�V3b[�J���z��ֳ�W-�܏�_U �du`�Tz�k^}A����ʾ_s�.����{qS���(�\��x���[�ю���;�t��^%�`"ɋ<����nS���|�2����K阪�U��Ba��E�E��x-"嘱ggQ+2���_Q�/>?]L����.u��tojjO�d�� �7z�1�ǫ3d0*+�Ȏ�a'�R�K_*@�ʚ��y��x�]
�`�v\��8�m�X�n�*�l�R�;�.���_\C$�ߙQ��'JG+@���b�w��`�9w]1*=�-���v�� �B��Ɇ��3X��xM%ws+3r�y�mds%E��p7�R��M_H�9�����J6k0qp��b�J,��s��	m3�������Ǹl ��C1��NQ��:�% DW�)��yOc�ė��uX����F��
�.2Y�����)[\6@���H	�aI�*�Cf��[,�ɷK�������U�b�4sT˽5����܅*Z	�E��)��J�f#Ʋ�9C!�=�w����]*�^<�"���Wh�NPF�dźjЂ�)���x�OvsdMgh�ת6���7�R���>z��ph�� ��՛�rGU��/����l�;*���K��H"�0轒V���4��[ʽ�x��1]�:�M���$����帢�mt��� �^������"+jK�&)5BY�Eo$�4s�%���pG:��y\��1�B%���)B���decׁX�Z��D[��9@�$u^�gL�]�ur�/.���N�}o1ޚ��rB�.n)Oj�C��iK�r�;7v�:v�p{�x���&�����
]v.u��)Zu>�&�{��윬\4,-Ú�
b.�r�&?����䨹ʑ]��5���o�8�c��^���.��2^�5zUީxuVdŜqFäN�/[Y�Ȩ�/��Yf�5��mX�j����n�N��/]�w��mv9Y���
�ЙK�HcP}Վ����68�ų�9IѾw�j�j�+F[�����k/Cw�[�땀͇���vt��
�4��m�,�5f;�n� o(�b-�˶�h�۴f�h��H'*�v��n^$�-�4�t���iGM5�r���U���x��F8��z��-��5ګAm�׼*k��V�v�^�E9}�Ð���O<�m87���%��K�ˋ)��+)a����]N��\��m*S;����)� ��u���x�p�/ORt�	#3�.����]�Ն��M`ٴ�l0�)��F�.8�vW���n��3 �^�RW�A2S��Of�:N��7-���B�E�}kk���+%�����x
�A��5���j0
�+u	�j+d�ճ��h=R�\��[���t��I82n�8��,2)r8�j:E�2�I-��\���ҝÖ���T���N���X��m�
�
)mUk(�[AZآ���UM%E2�"��e��]9m�0QQU�E�R�*�ZT��"�B� �1�QSVŊ�,ujj�
�)CUL˖��
��K�"1q�Ur��UEkB�,rʈ�E5(�u�P�X(�)\C"��AV-lb�E\��TEAHbV

�.�i��Q��MR���(��Kh�DATV*���֑UTQEUP�*1�8ʎk*
b��#"����T
%j#"e�D1�D���b��cC)b1Ab��U����Q�EQb0PP��Hi�LAdWV�y�O}}׿m;=���x��������(��5mł���dŐ7[k
1����R��l������U��������9����I]�)�O99�-����"mu\�1�C�11��\�1��>I��pT�'QY��Ǧ��ȺR�u1�aTa,V+����Mu��h���o��ˊHC诙�Ws�d��5}˪�r��y�\\�*
��2�j;�����`v0�,z|Bge�W:N�l���"E
���^��gV��(��H�@�Ԝuܹ	���.n&'ݪ�5œ�ץ� $p�n}Mx.���5�+�~[/q$_^����.�#@��Lmì����&+���IZC�C(��C�1]G\ pV@O/�15]�	UY���A���ġO<��]�z��Z��G�O����n�nr�Nh���p۵�3�T`�Ru�
�p"��ہ��C�:6͉�*p���'�/���jJ����;�A�P��(�-���v)d�s���K0{N�1�ݽ��M��$w����B�'f��q�
�dXW���a�Y>���f��F�¥�4U��,Zק�'���������H��̻M/6rۢ+h���{��蕡�������;=Y:1�z����ک�<Z��w�<�DV���oS��cx,�!�oE�zfEd���E;u�XdZ|:�`�Xk	OUhg�\K�q�c�Z��O�:;W6#����:�ݪL޾�R\��@|_l幍���h��(\���'�/I�T�t��b�*�2����ӵ��U\w8�3�o�x[r�z*Y�VFO�خB�U	YL{%]a��l�c�Fj֕M�J�\3��ʤ�Q���t���7!;b�b�d�%���S�15���:�J�(L88��w0��=���m�ʈ{DCJ�Q��P-�rK&�t���8�$.&�<��[��HS͉���f����*��ޮ#p�>)�r�'65��~A��@�¢���Ƈt%ù�)�0j�j�J��ue"n9m:���TqIT�a��Dsk�1{���ʬ�9,mfch�X,7�t+<�7
�F����J$�^�N�[��k/�}C����4�$��'f���TA���Tr�E�ϾC�1��3�V(��'rn$���e��]�*����1���i�y��WFޔ�;�u�������Ds��W�k��]��^n�θ���x�{wǔ]��OI3(Q*:��3\2wQzz���=��q���K�{S���,k	�[�3��yzi=ෝJ�ƌy��Aď�����vx��0L�[f,t��ܞ;	��,*�ʀ�t��M��%�{�����}E`�2�b��t�R��/�|	;}J��o��!�0����e��/�{�Oܭa_U�bf�f�3($�o�X�:W+�Da���˔��pro��\�F�l���P�>�X��Ob0��#�l����r�Y��l7|�NF\��j��i�S��Tz��D�����.s�Dq̥�,�@B2r�� ���`�7kJ��S�P89��gs�y�����ص|9�Z6�!���:Y˻�f+v�����Ú��������<0���LvS�4_�vތ�JH�F1>�#���mg.,�gp.cp4$z�"��UpZatiT�渟f�Bv�2�]���|��3[���Y=��<(W��B�\�OJ�o�1����(uZ}�p�>R���"�!"��6�����!1<��3�H�a�
�,���e�����VJ˜듺ӏ��XͶ�N�ǩ{�Q5:M,5���|)Su9,��7+3�߶j�Ji6�h6-��&t9�#�Web��SE�[Ea5�&&�{���P�Zw]w���l���kzQ��J�m(��gB=�L�Gه�YZf�5��q�ؓ����	t�������E�������O	,Luz�q(�"��S���|�"2�o�A2��QIS��z�y�|� o��]#�YЩߴ�E�8�+���h�[Rc\Z��pT��̱1�,1~�aQ˅yl�UY����}�OL{D&:�3�oC�FF��wQ�_��<rkHFo
��G9�Џ����վ������6r�=�\�v^D{ p�૤'ntw\��Q�3����������ã��J�w[�+��coc�]�ՏV��l�e�K�DT�
��yK=qX�wȂ��)����5.��*W�zFeu�q`�lyL�6x�W@lٯid��>���,!^�t_sma1lEv>m3u]� ���;nX��=���7�gdU�:�ً�E�נ�;,�!r����/!險�<=^oH�沽VmSS|�ϊ��k��1��fZsYA]6�{�F�Y��{1JɹN���C؊��0�K����&�:b7)V���z<�u׳kw�ޡ��	)87� :��a6Op��B8�Jpn�2p��o{U+w�o[�t���n�QC39���_:�W�Ж�WDۭ��y��$�Qڻ⨑��A�#yi��i�y�vh]��C�|�wSV�V8l���&k�����{���W���*zaQ8$G#Ҫ���$wsW����3M�j�1���yx3�@��FY�>���
��Gq�֏J2�a��IWJ���Ԉ䊾��,�a�4��C`�'�ܙTLqr�(2V)�ZtK��X�rZxs���@��Jޜ��$7s�'`T��. �d¾"Ui��nz*k��F�n�	~NX���C��p"�9:�q����"agUыF� �Ϸ�l�cY��Mֶ�%g���}tɊ�����~��f���[�"S���i�\���uWњ���=r�������^b��#{��J�}�Q5�!u�η�W��^^������CP��OW�,�F�� U�-�}�	b�="�q�.�WH�h��+׮`:����-V)�`5r���9$�GOY�M(h��R��Q�H��mf�8צ��W\617�� ���J�+�;&���]#�]Q�|.(��A�sH�J1��L`�;g&�a����9�-�j�yѭ��k�=�����#�����es��:ݓ�&�[��������g+zT�ʿwC��MsV)k���\��y=U�oA|6�3x4���8�m��Ev���5�*��P��z��nV��jZ,��u��l�3���q�A@�6%�rW�˃�U�b�S��=jR5�$x�@�)I����JswQ�EI삄��Eoc�Ї�`D��ؑQ�*p�B+��=tM"O6�C�zôz�߬��xt+�1��xk��Y;Σıc�W���TV
ٳ_z�;&pCY#�z��G�ǵ��L���&E�z�\ve�Nć.��N�5�i�n�����[�P�Ճa+ưmUn7�+JP�𭳡*��]<��{]�ݷ���:�!m�O�2��g=ncZYq�3Lh�9D51��� �e@顆-ל����׭�3]*�j��J��Pxq7O��oD�O�Q�Q�]��
k�G��+�zצ�����׬�^L��!:�_K�.�᚝0gd���;��_���ɷ��yB� ,LJ�QE��p0��P�׭>�	�r7|&2�����\�{|6����.�%I
(@>�	�vǟc�%�WM�L�uV����g,�5�kk��X~n��x��Պ���{= �]4��L�mg�ėv�J5�sc�*��6P��D�S�X��̜�Q��yEn8��\5�Z��h�b�t�����p��Vd����C��6���ϡ�Fd6��3���C|���{��ַr�i���ķ{�bP�1���<%ù������fb�M�ڑ��u����&��T;���$��*����*#�5��嘫�+*�R�����,v��\%�Bp�b��'[ �s���:L���̾܉%c�G^a����֎T44��\Ύ�h�8ؚ6�W���Q�Ȅ9�ɠ߱J���^A�3�$5��Lm��f/��:K�Q��i�G��z�ov�C��7��<��m%Wm -��e�K�^�*}L��'o�U�c� 0��QqIP�jZ�oV��q[�hi�uȅl5�g"1�>$�V�5��~S���Â&=���ckq��FJ��^��%��!��z��� 5+�.][}�p�=xB1L�E�iup��
lf�Ã5�I�T�܌[>��I�.�wt�r��+:cd�k&�pB2c*�<6܉�jE�܉�w�ݛ�26�q��3�Z�vw=μ�z:cwm_�m��]:���E��q������%�3ii��A�M��H������q��ط7r�m���n�����h7�PH��1p5#�۔�sr}�ݕ��O�xz�˺�T�{^B�u�v������N`(gl|��7*8�S�s�hL^~-K���^ʨ�}4����XmJ�1��Wm��E�n2������N!�xr� /��.��=>�n���¿iT��k��j����*��V�YQ��8=u��	�w.�B���*\�OJ�npk'�i�@����dn�{N��吪��9!i��\&'ɻ�g<H ��PTO
��d�S�jx<���*�mv��r�U+~�5���s<���d���s��zx����UĪܒ��F)�w�yټ�r¼�7������5<�Xa�*� ��'�t�a���|�p���o/Z�z�Z�u9Xv
�^�Bw���&�]0R��\���נJ�������Ĺ�P�1u��H㓑����"cxU6r;ٶ�g�#�i���R\�y5γ���=��Bv�t\��Q�0��,To
�����é�nSA9��6n�:���]]&�H�6�Έ���������D����C�힒���pi�������r�:P���u���c������M>O\2�7C�i2�ؼ�.�W���W��HC.�p��woM�&l��F��0$�j$���[W]K��ՕJ���]뒖��vЬrke�e�w�������^ږ���i�'U�:k�Y=��T��&K~a���	�������,��'��y*�����q�˵��,��aÕ.����zjWyŕ2���6�{�J6�9)�!��w�p4Wj�M����/i�煍��ܻCY+��W�\R�g�R+�'*�����3
�����,2T<t�nR�8�]��;}�/7k����b3N��oΝ-U�?��ޔ�����N����>�+m-���7
�|}�V6h�0lY��g�����j��>��6����:;���z��o#u�ę���	Ԫc3<�uY����k�W	D�;f"�=J��uZ�x�'vzV�b]����=���	S��	�D���jbCw0��vA/�x����h���1�^�g%����]B��;�G�
������.ݭ��^T/{Etx{ �㉀%��}]��CX�0��N�d�/3�Lz��Hإ,RwQæ�֦�v�z��G9�2�79A�f��'�|^Ƶ��!�g�l��Bf웳�J#w�����
.+,�D�ܥ��?I�������.Yg�L�=� �l��Fl;:m�엸Wm<��r��oWb�f���t�{dQ�6L.s�p��n��U�׮�j��|�ԣ�'I���5>]P�D�vq�}̘�S�Lڝo�����GvEB�=���G9#K��|��	b�=*,'.�WT�`����;������ҳ�3Ю^�Pb�tI����k��A
�у��,0wi�L�u�6y�m���1C�g<ԑG*co��*���$§A���{�])�^L[�W=�3�����	�]m��8(8��nyo�r_��J�#֔:�׼�c-��`fF�7Q���C(�e�;)@���v�g�Ї�v=4$\ژ�{8d�M�WYڦ�����+؃��ag�r��a��lk��Y:��<C���vWj��wS�Ee�Ċ�Ɗ�(2��2dXW���_�ܫ}o��ns�.8K�����:t_�ƓL֋��u�����¦ߜ�ۑf�S�^�;Y�^���%��yF�xy�=鍯4�#p�i��9F�U2�_��J8�7q�??=�Wh�Ӭ���/��e�4Xj�6��8��'�J�vVT!�T�7�b�m��ޏ"�x^Sl�z���q��Y�ŭ�xн].�ֈ��G�ڛ�]����V�%Z�_o2�Ԅu<.*�1`�T,d�*��L���gf�ڜ����e��Mt޽�L��k4P8��;\mÏ�V%[��9��T2�ou�����:��ɚR^ۭ��朏�
��¸��%j����o�aܺ�K����Yp6�Y�yA
/�#��ZB�c�n�2*c�+n����;�p�z�f�Έ��'0����"�F�F��I�]�@�Z�#��]e*��[�r�u�}Q%�S�K���OJDQ��F6ի�pr���:z�ѝNV��p��`�J��ឪ�˙��+�F<ǈM�k��/D��w�&܍t���s�ժ�jܔ�ח3��Y���og+��E�.Mo���(V&'vQ%K��(���\0>6�kyziP+�۹8�7"�Q�#��B��_R�w�9�����־�ս��O;D����Ӽw��������=7��y�l�V��VǡNZ5]}'H��L�٤ZMne�z[/�]�j�o'u�*d�V���2d�d�}�h�m��#�G�zupp�ǳ�(N��97-TК۸��6�c�Ԇ�o�q�jeҮFGuaČ�9S����eU���o:����rN5�5]�MF�t��W�Α>�r�а+Up�@��Wp@R���sqKy+o��l�w;�:�̃�6��R��+�50\͕���E�Ρ�8J�� �g�:�V#�ubY���}Cq ��܍5pB����:G�d��*��Z���v�;yY|V6��@�y�\�Z�3f�Q,u��ګน�r�vќ_nT�}��/�Ff�Jf���j�՛�1ڭ�vя.��,T��RXe�ܟ�g���s�ǺM�?a��kv7�:���L��&�0��Q�f��Z�J�eb1h��g��%��e��^�0t�y��ĳ���w�ek�(�.�vbt�������j�o;�՝6[���Wc\���M���؛��̮��ۈ�qܭ�wi.�\�i$<3Q�د)9���-��)ʴv���S��=�}$�lk�՘�D�Jأս����U�3أ%�+h��gaF�kY��P�ɸ�K�`��4�vr�����.;x2cp�1��1�-Ѣޗ7�U�lPVo�.���G@dm��c�n��lYǻtCk��p��3rC��f:�k:`0��k@Z�'���q���c�TJ�p!��"E��*�
�)Sl���A��MJK)�Ǜ�$`�I��bq���]"�Ɂ.̶/��]̢��+�����zઙ�5�FVN�ƥ�1QV �	"/H�����Z�"!Q�����ej)b���Ab��UY�E�
��VƲ���J�
:���mӉP��`-l�,��MU����jAf&1a��][2ъ*��$)�F�QTt�,�kb$�f"���eK��Me��M!��b��TJ�F�iMS2�T��*Zآ#F#��	�Z�c*�ƥKm�&5աm��I*,���-P[k��֤Y��P�i4�ɫ�
jʠ�Jc�U���ur0�L���N&*UM8���hH��]28QE�,b��EZثuQ��V,q��I1��*6�ڣ***�k32�5�Ʀ�DPQW)dSk,�aR���ĕ����_�]q-��u��H(3�#�2�l��.�* ��������V�ol�p�5S�nQ�j���v����Xw�B+�2��2�ÞM�Ⲣ�R��v�V��GԧK}پX��k���R�C�,��̫��A�'Q����H[�<3q;b�b�V�N�j�Pmf�o&O���L�*(�'
�*���"�9�F��LdX��Wj*v��[�®�"�j�.H�XU ���\`^�g|��
y�3Y/ճ�H�S�cq�]k���u�a�����j*;Ti�;N����\S5����e��_K���f	l�S�N��
�r0�ei<�&ܩ��8��+Mx�%�!-�U��sn+3��BՙB}�%�~(!Zm\������bQ;X�S�rcVw/��rj{^sR���NJf�SB�h�r!�4:f��0	#�mi�U|�����4��1�u�Օ
�&:-L>��ϸ�[��b�:U�ani�(k{k-�{�c��0���F�W�Y��h>x�ٞ/�|	3آ���ۀŐ
�͞wZ��/��2�j�n_��j�שoQ��=�mѤ3v�[�� ��0�IEn����
]�-��ͺ�e��TZ`O�M��9PǷ�\��dy�:���[e�w��V{NX���:�-�!|��r�jEe�Lb���~s����v_U\�Vy��xh�[��b�����lS뮓:`p�I/wkw�5.�YI��	�2��F4O���U�Q�^z�׊���(T���
�N�ظYx�9[�0k�p��~Mg������Od����G���V�ˢ��[�V����j��#��K��#�X�_Di������u�)�7v����n�p�vq��y��u��x��_of��pJ��&uӁ��ʨ�~�e�urƨ�Lh��k�\1������X��v��q	�^��T� �	�Vy�0��ZahR�Q��kV4��Bf�����a9r��ãԸ5��:�I�kG�Գ�r��;���]���*+���c����B��LJn��@�|o�D�Rɢ��u6�d�/��~�p:�Vߪ��̪[|&T�S
My�k��GO@�xIbc�aW���M@�a��UD�<"���K���dTRTÚ�J������ǦÚ����pR��E�=�q��T��T�n�E[{��fNQ�=�*j@q�7�I՜T<��7!�,p'^��ӵ+1�Ϙu>���G�B�c�PoW�ʝ��T�<�����]���zg�1JٌP�ղ�nV���j\�]��ʊ8����s/^��u�	�;"���.}{fP�ޖb��yl�Zj�|Q��R�2�~
C�UE���mu]s5G�MaA�P��2��i��^�ѫ�Az�Ssݼ�����\��b��c��T���,��㋽�3��w齾�⦈���m��̀��v>N�E3ta��I��rDX�����.o
�a��o��2I�C-��U,�
ͨ~�ʆ�tB�n5��I�ut�C�2i�nZ�Ņd�b��0*q�IL�H��I���\.��nS������}��I�NLo����]M��зwv6a�6��g��$FIh߸�xSͨp4Tv�d�c���tmuy�co�׮�ş.L�=�IG/��aΛ&2q�0re@�����^�N�nt�ɨ��������U�ט�trndh�n<"�]MX6�V�����&H�Gc�]ťz�W�ªgq�E$�x�c��9�n�^��/"LT�Ѣ�!2T���x$uE����iʌޘR7Q�(G'���N�X�����Yعu�yN}�VY����V&3,�u)���{T�Ex����7�~��_��}b9h�s��9�s'[�c%e�
H��α�k�v���ˍ܄V-��%rp�FHbj��۰�R����F���8cj%u�O�o�dO���=��8�����T^��˭ ��;�;��, ��oD��Ʀ'���v
U���.�������^Op���Ƨ����H��,FaC�-W+��G�{D,�0��3����+Zm<���`���ڥ\LTAS�oĮ/2��|�5�������֖ݶO�;<�ۓ�RΎ'mI���>�χI+���+��{6Lu���A�.�c�(�YZ��mcR�
Շz���"��xL	�s�4�+�ʆ�������u���R I���+���ˇ6anʢ�*/�Yܒx2t��s¢	��xh��zs�;٥�%�_�|J����-R����mI�r�1��CP�&*:Y!iλ�*0�E˺�ˋ�[����x\@Ә&{��q��(F��'�a�8��_ox��G�}��(�|�_��
��ۭtu���xP��}B�m�z���7�vl9��5�PY3.�ī�V��v�M<i\����ְ�Y�9��j�;���ͮK/��?h��n:�@�Ifn��Iq���Mv��o'�Iه3ywW}jعO�r��$&X���R�e�_7o7v�S+&�\BYѥ2+%9)�{�:wb��SGp�O�K��-�ϲ���D6+�Z�
�f��,�ʈ��R��z����;6�~�ZuW9.��.�'�4����
��Iޞ�#�_+mf����q"�xP�;槸��:.4ƓL�*cTo�c��Vߩ,��<��I{�`��,C�puu+��������%E���inF��5���ꏹ����g�f�+y��y��Ei�1J�j����a�m��.a��]���.���17���3ɏ�hz��W	���d��ɔBu����P��Gg��R��I��9��eI� )����8�\=Gj1��r�Oe8.�e�RnL��������Dn����\��Pl|�>����<�%�5HS'��<��̚i��qX�(�S�Æ�q�]?�T�����|�h�F�;�օ��X�6�h���F_ǜL�����Lź��o��C}�0I蒴��(�7C��t�26P���)��8�fu8��d��<�sQeq���z⧆�]n��˱J�M�YQd۾�qeҌ��Ě��.�x�[�t)�d�׭���g{e�%'Y;x�Ҷ.W1L�4S����X�CE��'MO���}oY�G�0����F��.OpB����Xa'��!�Bu�s�����U�;��w�):A���s�P�Y��cã�4[9���pPci�y��tH8�U�f����Ga9r�%�
�ǫ*���q}m���\
�rx�aT	��L��ܖ�^gh����~;0Ʃ#�6��å��_��5e�L�(��ء��9���<Pqi�i��p0�'�!�Շ�Dc�$V�5�ç+�sݱDZ��'u��n���W��̤��Ny�NB1��mEg�(�z��1>�(Q����f�i*S[�N�$'�3��f��d��=�=	�
�Vt�
ɚ?/`"�ڞ_pY�@��3��td(gW�x%2���:�1����6�F�r�������I��Ѕ�~%��!�����0���U�:iYCK��ڔ6'fq���{��ƛ�����#(ؘf8)(=g�W�Q����)��J��A�L����΍�;����-��΂C�|��������fu�MriR4�[��}IM��,j��_R<N<{��_.u�4L�۱�Kz�{����@���&��ߋ�%�]I�5��i��d|��n89�"�䄱%��{�u�	�.�N��fP�2\�OJ�Dpj��!	�˵�U�G6��!���B��LL&��$��0��¥K%����x�`fìM+5�u�!9a�za����n�>S���k����'h2tU��&�wH?@�no�Ez%O9H���"�As�o%�27ԕ0槁�+:�b� 	z:%7��&�q�ƚ'��R7e�Ir�k�/YϏ��%��K[0����sX��%t�����xRuf�p��``mfK[o�����Z9�K�r��w��*S�ƞo|��qJ������]Wũʒk�l�<0Ƹ[�x6�������u!ͻ�=M�U��v�U(	I��p�F��n�8W$�d����0�sxU<9����$J��M���F�����T /��A�r4�yw�6kK'��J�X��:rN��+�nwod}�G�����v�V�Q�JBܦ=~����΀�}���w�,U�n�J`���-�-�4�X�z�u=�E�͍m�T���se@f��kfNv�&�*U���n�Q�A���i�ݮ�͓-h/f$J�Ӄ�&��J/������w5դ*u�wmlx�@��2�,�r��u9
���R���f4H����q�������j�M�=�m�'X4���>��h1�򏒃o�^/r��*�V:�+ӕJ��`�Q���܎�+����X�7��A)�$�OV�V��Z��X���`<0;~t֪�V;��o΋ڽ���>D�[P��a~f=�-��x������SD5(L��zX��������5](f��B�/f�L����aoL0�t��B��{	\j���n5��=�ڬ� �Ѥ�>N��T���!�B��Jޜjb|��('(ED/#t]��Y=��Fd:44�0�U�߱K���Z�o�:�q���d���V\ɾ�tr�k?h��A	���\LT=d��K^�[�"���[2Љ5ۯ,���h�[�i`%\<����f��Yu-S�瘘Tu�c�l� �ھ���c�J�P+�(A����{psȨw�0'������4pK�����V'R���?k���2Az�<F��u�ZҎ�죙|�"�~�>ު��'X����h�	'��/�t�4�»a�w���Ž97�W*anN��$�@���z���)��{���lS2uq�U��M�%i}!p�sGk�f<^�^�u��ˁ�
��Y�Q&�œ�Ե���J���2m*��y��}�{�F�#EJ�F)!Tl��i���o*c\��=�[D���=e�dS�{0l=������֋����0L�u�o�
�%�@�O.�l��Q�P"�BY�_�,�ܦ�]����W��{���z��w�ݔ�EF�;p3��C�8{~��eaWEٿ!�ғr�$���g^^ǳ���l�xY���u��V[=\3f�t\Pi/{�pu�zp��u7K��ӡ��U���>��\��ei�]��Vet�R�)3{��Z`V�Y��~��i鍎����
@f�)މ�w�}!H�u��㺅(����z�t?9��V���̍T�Lg���g"�ƴ��^�B��<�}u�>�J֨o�J��K��^t��j���L�����n��smJ��S�Yq%�g�KM���[�]�����e]md�c�W2��1�����xf�-N���ಁ�DV�qJVzwW:�	#o.������Ƿ�vز(�{��-'3j ���`�.�܅��N�+j]��k
��������gsr�"R�d ��aޭˑM޷6�]=���;��L(̊�nGyŰ��xI��{|���D�	�LTS��aZ��Lt�ܷ��Dߚb��[�������"ZWr�$tT@,*�>�0&K��sJ�
�Ե�Pk69��ț�WR���'�ᨬUF{�'��8QbP���s�_K3���葜İ𬂃��;�)T�1p�+I���"�����G����`��;�������SFX��MxX�e�Uf�����U��H<�l��%�F2k`,�ɍ6�Of�H�˪�;*J`a�SB�h�[F�Dٶ��ڃ��D�Ξ��ܛ����|�Z��A�z�'�.\�bmL7����ihƼ������ɆW��`c:#<�<��(�fRš�L�)����$�%�d��4�{TS�G96���}�W-:��O.�C�2#\���Y��D찧��(]��%�K�����/
@�cSn������P01J�.]Z�/W����}����?��!�_�?f������$@�L��AT _�$��� rj����3���C�R�����j����C�4��f���Y1��7:Y׆y�qBB=���M$ċHH�_Nr%��%͆�3�B�P���=��
B���@�k�A�i����m��<��� ��$�
XjT7�!���34Y�����C��&p��JN����<���8`s�tu��y� @����̧O�>��x� �0��D���	��:������!�?П�����VO�t?��p>�6� ��Q�8�� ��O���� r����@�Q*q
%��d��6�*5!�T�"O��g�����w�9h��_9�r��f2R#��** ,��E�F��ں;LϯL�z�� aI��V�D�
�O�.y��h&�W^C�.2=@� .ke,A�nl�@x�y���v�ǚ�Ri1��K�*C���������ĸ�<�䬞�׺��)3�0ʪ�^����h*k,qC�	ǒ>�,\y��-��@�%�C˨�|9��x�M�G�ـ�)���wW���m9(� ��a�ä`!��Ω��W ��${C�IȗkDa��`*����}�j��9D�&�v��d3�\<�0*k*���5�D�X��!  q4#l��0lE言,�-I��B&�xYj7yj)���[+RP?| N�>��N��~�	1I�57�Z�4b/�{ʢ� ��Y��;LQ7)�E@��<N�~�"�m{6+��z�c��t3�8��?@�:!@�Xn\ˤc�t�B48�Ӑu8�����ɵK��L��J���st��H�T��Bd�^]�b`��QPe}*�c������2����6!��bv�_��oV$�w (�#��#Y^�y�ڳ��^sS���Ͽ�x�1�#_[��* -�px��W�)�x�\�`A�xI����M�D$��IN�
�r�Ī'^A�� @��h� � �Oo��à� �;Τڐ��0�p�#f�b̋�V�z��:R��֑�� �ID员�Z7��]��BB��L