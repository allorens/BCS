BZh91AY&SY��7�8߀`q���"� ����b                                              �
` ��|��-�� (  �  �   �T�� 
      @        � C}���� T��%ATJJ�PRT�R��U$
�HDJPJ���H�"TPE ��!@ o�JPԔ4�Ԓ�A
Q���|�P��J0�{��W 4���&�ɒ���D�	��U&誩8�c"�w�<   �Ҋ  j���s` �Q*�� wwW�({:J{ 8�� <��*� c��>����>��c��@|    �>JP )���RH)T�@(wq�Q���c]� ����������@x޾>�O�� >Aמ�y 8�{ ����EU� [��� }���   /�>�B��� ����>��E"��n���ۢ@��'���>������(���
wX� �OJ}�y=     ���*��/�H"$�	B��Ri��|�ww �p}��@K����w�P �� OGV�s� ����t��*�� �� ��`8�P ��R������s� ��)�=� �`u���c�` ��y��� ��� w��} �`OG{�x  P ��ʨ�*���)QQUR؅�#� w`:݀�;� ��y��{>�Tr@=�8�^ǽ�<p:E\ ��v  A|�P 1��v9 9���Tx �x����[���� �r%�`�{�F�    ˞} ��RE$J
���EJ��` �@�Cv p�z��x=� ���;�C� �IN�L�n��   <}� ����;�U*���v� ��� =M�UR��� ���H��}        �"`R�M4h     )�)*�4  �  44�j���      l�@)*��h�#&@4�M2bh$�$	J��� ��A�h�A
��~�ML�4�	�h�����i��>߬���}fy���$��	��x�}�/�8}�y�� U��W�A>h������*�}���g�����S��(���U_��W�A��А��TE������~?O���3�������&1�0c0c0c2c8Ɍ�0c8ɌɌ�2cc8ɌɌ�����0c3������������2c0c0c&0c0`�2c60c&0c8��0c8Ɍ����0c&3��c3������ɌcL���2c8���1������0c0c8���Ɍ�2c0c0c160c&3�����ɁD���&0c0c3������g1�`�`�q�g1�1��L`�i�a�`�`�L`�lfa�g1�1�f�	�dC��q�L`P�Q1�Le�A1�1�&1�LaSQ�1�LaC�E1����Q1�L`SD�1�La ���'D�A1�e�1�LaC�N0����
��2)�
c �ȦQ
�0$Ș�&0!��c ��0)��e���c �ʆ8�P��1�eC�A1�Le�T1��S�1�a�D1�a��LdC@�T1�L`CP�T1�`C��D1�eC�1�LdCP�Q1�e\a�L`SD�T1�`�E1�LaCY�q�eD�1�LeC�1�L`C�!�H�(�LaD�Q1�aP�1�LeLa	�Le�1�`SD� q�N62��1�LeT�A1�LdW�1�` �q�eW�@�q�dA�@r�A�q�8�0��U1�dG�q�eaI�`GQ�q�`GA�f1�\a(�`W�Aq�\`Q�ʯE�q�a�1�L`�U1�d�Qq��Q&q�eA� `WA��@� q�d�Dq�\eG0�� d1�\`�P� ȏ�q�`�q��FeS�q�dGA�q�Z�T�1�eS�q�\`N0����dWQ�1�dW�I�q�1�q�1�c1�1�1�1��c'q�q�q���N2c2c&13��ɌLc2�&2c&2c&2c8�0c0c2c&2c�2c.2c0�&0�1�0�0�&0�&0�8�fa�a�La�Ì�Ì�Ɍ8�0L�Ì�ˌ�Ì�3.2c�8Ì�Ã.0�c0c&0c8�8������3���10c2c&3�Ɍ�x�`�q�1�1�d�8�0q�1�1�1�&q�1�1��L`�1x�NO�>���_�������pT�ޣ<������>�]�����k͝�u�{�dz{돟X���t,���@��N�\4�T���B�G�[�w�#iԝ���{������b�_���틄z�r[��扣���:�{\�^�=:4�����U��˴ɗSs�LP��0���?QaP|��Œ>�5�BdD퓵�tꘇh�Vܠ]�ݧ�ǗM��n�o�v�}7pvSx3�[xQ"bS.2��
 QǪ^t���W,���� I�I}٠�����Z���e8���,F�h�u��	��哈���[��Gl�sX8Գy#�&��l��"kth#�L�f⋲#n�X�9��/un�{s���;�;F��=��b��R�w�!��[\�����	b&_��+�!��	��>��BlX����������Yw�5�Y�n�����خ�/�]�lېnm�e�{f ���$���u���*�!�\�Yxw�Gj��n�E�/x�3�dS��hf������ǌr����o�ǁ��$�ָl�J��3��nɹ�L׃�pj)������ۯ���3Eg[����	�f�f�׫~�Wi���z�=Y���Ye@����G0ss��f�ĄW����{&3�i�Ì�%�]�$���^snn��G�y((_�UU9OR�LBL\<��P90�%ۜ$�:n����w���^�. p�Jggn����2�R5F��;zs�IL�n;^��+������Ö�I%oV���g�{�.���n!��&̣��<o=���s�f�60y�ñ������9�{��4�b\<u����ȯ�7w_IU5�q6!U��z��L$�8��4��F*	/L��pw���^��Ƴ���'$M)1��7D�w�n��2��&ԯN�q�e��S�1��������q.5)A���܇�5�]�I�Ƿ���ȧt�x�$�D���;����D5�8�X �xX�m��n�'i�w�I:�9�I6���!�{��^��{����3��:�}ݷ�P�󒙄��9)��4�9��s �׃��>�ӂ���|7�rd�����K��������سZuV;��j(rs5 ]w$Sٽ`�{�F��7�5�{�N�Uh��x���;c�۳
�I�O"���ձwL�Jz�����e1(�d�q�����w.`For\��mv����[�^3��_C�]��0�n�C綻of-or���;B��9ٴNZ^���]��L;ڤ�����7pvkr��i0���J��`Wb��x�o_N��)^K#���C���A�W^iע;����j�h�A;f��_js�t�a�6&V
�1�Ο1�x�߬�N�I���z�>نWu����6�]M�c7�t'𻇞�Y �c�r���2���[�����'GٻgpXdj�rMo"��F�#z���x�%�R}�n4o\�lJ��p`P��gC#� s���������{�b���B��H���s��f�k�;��a�+6��qd��ǭ͉p����8����A�o�(3����Kd,�3}�J��29�d�2=}��R��O���1��.�F4�ׁ5Ϻ>9P��=�Wiz�jD�Ǔ��%�9�е�k��s�+��:��,�됙ڃո�ev��zC�бQ9�fj�We�˻@Z;waLv��%|�ñ�N�2.�˥[��ڷO.COv)U�a���E�� ��3H������D\ܦ��S�,X�ܓ+�Z<�����Y���'�0d����[L�v���#{�]zu�;cqn��.�D���ɳ�ʳ�gT��Ke�]�=٩�SL/{7.��c:J���cŮ�d�H�� ��^�`q�#�S٫c��=:wv�Q��V�Kt�0/�a���qt�C	���P6���K�A�ٺ�n��3��z��S ��K�O4Hk���&v �Ŭ;I�Sh6��\�6sBѬ��.iU�k���{/Cg�V\c�J���N���Q�c��w��DC@h|ηO�����
Ž�}\�K�n����C s���7�\H ͘�Z0��Wc�xs--Lr���(]$4�w��gx�%Ǉ=����:4�zX�3V[-0`�7��c�I8�Β�����+�:��L��*�mC���:vI����/(�'$EX���T��9S=��ݏ&7L2�d�&���Y�Ќ�Dg9�M�.h�;��s
r����2�w@�.鈧o6B�Ǣ=����	��Sx��i˨��(c��.ͧ��vMV`��3�ö�q^��l� U�otȷ��9��;XΪb�e�}����Sq�eglũJ��g>U�p2�\��J�t�H��w�n�nn����Qy�jF�k����k�o����޹͕�{�T�X�	�t�[�>��=`��"��t�ʫ��&��5�p��Qt���U��Ճ�NƐS	�&��^�v��aZ!o��]Gchl_ww\����\g���1�,ꓱ�WE+��˴U>��:J��̘	�,��x&���=͘��V�՛e�՝��H�^�^6�<@�8��ۻ�M{B�X"w`ã����FШ;��2J\�/n��v�{��w�=�����׽Gf�%�i鳝qj�-����ڲC�vw!�܉��Go�ۜűZK{Q���n%Ћ�xD����[�������=�E����*L���Hu�	���}�V	1��R{�{�dw��p$���a�s�0�ygZ���#�5p#M�uL3cz��`��+y�d6�:,ѽ�>�+��5x!����#���nɣ4�/1�D� �:Q���jʙ�5ۼw��hjw�9�H^��h]xpx�!&K���:U���7����'x��s�H<�.Ó��@���Qm�[�F�w��c.ͻyI�1�)�r��f���jg�h����w�Ty�8H�51��+��!j
#^^�����n4�7�W9$U,��ܼp��.4�ëKE�U�V.�j�{�K�G+|�>n��f�K�j��&���!�����v��SC��9	��-c��vA�%�GX�{^vp��:�����\ӹ7C{�q-�ϟi|z��'v>����7a9dv��%�H���V�O>��h�r�
�ntG��9��[ ܃!�e�Nܘ�HWڶnF�����>�R�z��卌KV�:�ӻ�`��yƋ٨H�9�gc��j���x�^�	��P�Q���F��7zsS9����Lӛ_=q�����/jYNn��4�/7�-�w��^ف�VFQ3u&۫� ��!�)90�w�p���"��-�Y��|)V���br=S�w->=���ц͝�~L� %Z�7�Le���.�P��n��vw�9*�W* 0a���@9hI<��P�ƃV�>I㷕�˜�:�Y�]�@Ն߶z�K�2���D���e8�z��9��Yb@��w>�~��������tQ����S��qE�j9���.[r拹gE{Fmû#��=��^�i�G�a�{y�}�^����*�v���`�e\�������o�����S}�|�VA�sO ���D���)��i>��)lI�@���N�� 2n���V�V<պD����{*�Dg7���΄�$�v�9u}��K	��A�n�-���.4��v��j"q��f�nK���v>���,���X����Na��7ۺ�C8	U�fP�zv,Io-�.�m5�Ë��P�i�ۭ5�p���Z�v治��،�����;�q�|9$ٙ;�Ν��G[�k+"%\�W]SsS�_A��ͻ9y[9i���;�q���bſl���@Ot���6 $�:�?���}�x͞;���L{����۔/�ǈ���F���UҴ�hߩ��!=3K�v]�1���u�. �s�r\����5X�����;��-Q�V+r�Agn�s�FD�1�:�|wH�0��.n��X\�V�q^��v-�-�աՏ]NE���wUX�ws|�lS�EC:��t'���8��n�����޼��uv�h��/	s��8?�<Q�b��(�D0l4��"T�Qd�;�@^��3�.7iZ�Q�zoe�.��FG�%ǹ���]K㻌f�����mL���r5�|�hr�z,�'��m� q��#u�,�,�ћ��#c�²�w���E�}���}ر����K���Ɔ��e�I�ܐ-�R��b��z��$�qE0���1(;�r�H$���Ҋ��m�|^&\�&!���w3�ȇi�ѕ�Ք)�<�W�wU�b�ɫ	\w��"��54����}1����K��.��L�4�/ww	4��CGQ�5s�a샇q
JK庀X�-����l��b����B-�;��Y�4��$����7x�=��8�C�����}��$j"��m��D�r�5�/��l��;`	��4r�U7(�.���4��;����I(���AV���g����X��v��3��:������q��w͍��1ٺ�0m{sY#�K�<��;`沪�#�wS����Z˽$�����5j�g`�*DW�4�M;���p*%v�.�Y�5�f���zಫ�n�w�9�g�.$�f8�<Kgl��3R�=�³W�G�.>{�9d�7�Xԙ�����%s��+7�A��nh�uA�M�Ds��S�s����� �t�Jv��#T���ݨT1�C��GD�f^¹ν��Ҩ5�1��ꝭq��N��ډ�NĎ��ý��β��������Ȥ;�5e���r����{�b��tܜ��Dߎ�[p�}d�I��ܘ�6�[�_�h(.�U����[��3�3Wח�1�t:��.v�øi[�u�Rӳ x��]��e���t��Owx5'j|D8[���z)m�fȱ��Р�����	3UyJ���oe�	�,B(���m+Qܨ��6�gd9���d�^v�`��oxm(Mَ�@�Z:��@�h�E�b�J��;�;���ŷ:k�KeN܃m������x�MFL�y�׍-lY������gWdFe��םRO�&)wh�A!hκ�SqNv0K;��7������ݚ�7.Wr����&8���p\��m��ې���w��3�[]�v\X�>.����;B�Z����_wN��\2�
d�5e���m��H��d�:�`�ǚ����DS�WK��yN>I<�kܔ��)��n$6�m���B�_��9�z��r�BA�睵�vr;�g5�ꨪ����{Anq܍\�n]ū�q�8�d�w+�P�p4f��c"��?8*�
Z�%ż6�e=pA~!�E��zN�r���9���򼛆q�����'�{��lY���E���7�`8�M>l�9�/���p��~��\��<���4ܓO�p�ޜM"� �K�0v�c����$s�<�(�S�f�����Š�+�t��m͈;��n桓�.��94��Ǿ�;�h��p�X���7��!��^�N�w5d<��{�B0+U�owI��J� i��|�B�2P�k(���������p�y��������[&���|�L�V�C�dt��%nuz�ܸ������Dξ���.�=�p�,�K�q�:[u�,د'��vh�t������i��ٷsdvp*�J���q-�jl
�*k~�N��g��8Y�r�9{C�
 ��<&�-�3�QeQ��_c�o<]�{�I�P[ټ��d������ݍ��9Y�8�N��)v���i}���PÔ��κ�"���V��+XX{�ר�ֆ{�}z�{7L�$���wC%[�mx�=�_�����̋������p��׮Kj#�%ۄ�<ɯ:�yٿLهB��U�0L*�7uG�]Ys��ڂ����2E�\������X��g���ſ:�*�\Z��o�2����:wPLݗdL���Kdy�}��N3�wa\F�׬�~�N�WK*������{~��A���c^:�KG7���=�(?��查x���D���x���ܺ�`g�]�=�w�|�jcS��˲�YB�v<	{��X_nl��L��ų=9$)U�����3���	��O��n���.ҏ���=}+����a�eM��Bܶ�&~���*� �G�f�w�*����
�&U��c>%���C�Ld����2�W?3L�b�W�`�1�S$�o�V7x�;��)�?��P}�y�OK	t͝,W&�I$���{K�=�	ۧ��/�G���������	_G��^�����}7yq�;©'�&�"��"�߻��t+�?$�9+}&��j���^�o��1��͇6o�:C�w��Gp���V(�q�x~1�����7U^~�'zn��{y{Z���qP��x�Ӟ=�c|Q�_�o�n�P�-�J;N��y���A��"��fn���R2�6�a�ۻL+���;R�ww���[KȟA�%�� T�������韨}L��g�r��n�F~�I��L3��76N���d��:?lޝ�;�����߷G�]�,�;��g7�����=Ȕ�m���X{k�p[�z')'�7t����E����u�>������T����-�w������W����c��X�Y=x{e�e(�'�� �I<��o�~/� =OK��P;��'��� ��C:��k��o$��X�'�k��(��6�Ic�&�|<s�yi����P�Ư�<�m��4���M�I%�F�ϙP�d���f�/��f�6�zX6P'�+�v��������Oi'�@�p��P?��tl�8���|ma W/�  _�U)hJ h�J@)Q(
ED�Th
�@�D�)i@)U�@iD�@hUZPD)U�JDZhDZP
�JiJ)E(UiP)AiP�P
�@@��D�@ZP(V��D���V��ER�F�U�P
P(JQ�@����J@J
EP��)R��P� �R����ZZ R�Q�@�QJB���)U(Z��hE�hT�ZD
��R���[���w.U,I���:�1��U=<��i|�i�ͱ�b���\�Amd��w���|&O�p�!��l�*�<	����1�G]V]��:���Z|�y8�E:�
F$�2c��%��2�q�>B7�'��̾鯒�jy��<L��"Yi@�I!�py<�P�\��w�ǅϞ480فcfI-(�R'��xY�|�z�'Y���|�XK��ό��Ny���S\U�|,'�xWIZ�T��Z�*��|x����O�&2!�̬i��Z(L%�I�
�k1u+����oz���S�{�w�1{&G%��i�ms�Vx���w��O�O03�|��}r��!�����˄�������y�ZC�8���"�} 񑣶d�����N@ �,c�&f�,2V3���b U��I��c�W�0�aaD2)��?��
xraAah���te'���&���&�c�,`���\�h�����2��)-U��6V`y �t�ѽKu���Q�GvҙrͻG�RHB����?���I ��}=|G|>^?��;DD��~����>�?BQ���G����xį+H!f̑	���˫9'������ז���3�x�}}��*i�d�3����rj,�숾��#ԩzw��1��ۛ7��H[���Ww�;0�P�5H8��V��J��WCqb�K[��״�7w�u�l�6��v�$�w�{�.�a�O��Fq�ۃ#�q�!�(Cw7��w������/�us����{'�g{'���rM�~��h���+W*|y��7����b=�ջ'�S�6�n�n����@�ef#k�s �e�+�F���"<=Jrn?��� ΃wR<<4
}�9Ѐ�v���Kv��˞[��ϲ��9Vf�����Ց��8��z�d���L�q������Ӽk������;�{��ı���e�'��d]*'����7��K8��}���� ރKzHknK�Nﺝ�`�^3����\5��n֍���~�}�(�Jr�|�v	Ew��0@4v����c�_�;�غ�٧g�+���w��V"��������,��x`G�Z$�24we(-W��L~����yw,�
5��n�wL����\
���^{2�8ǳ����^�M��s7٥<�i���ylǺ|�I!�����J��ex��W�;&v���[[ccCk���Ӯ�믇]u�u�]u�뮼u�]u�_N�κ뮺믷G]u�ǏN�뮾u�\u�]u�ˮ��N�뮾u�\u�]u�ˮ�뎺뮺�u�u�]u�]u�tu�\u�]u�ˣ��뮺���^:뮺�믷�����x�}��u�_N��뮺���]q�鞞�|3������Ʀ��@<=`y{��!Ec�v�ت�i��;�?D�,y����'�n�-��nn>!'�!K!ݭ��w���G��#a��.]*[�K�WVB���m�+=j�:^s�ʻi�xY���[��޴:NzwOt��}hy����W̅�chxa�Cs�������}���]�(�2%����=�����X��j=��^^2� ���E)�;�3�����{'��p��ټ_n�����O���q�v��_Ws����7G������^
�E����C���!h��ѳ�� ��c��Θ�aN��r��ѯ=G.����rO<��{B�������@R����M��gzd|7H~��%������
;ֽ��^���F�9��v[���.kԮ���A	�g�c}���8C��׎��/��Wl]�x�A�N�@�3��v��6��yx���<�'�#V�,���i[n�� �f��#���j'���ÂT^��/g	\��f��D�8�h�Y�Fb��:������5�[��7d�dŨ��ަ����=�j�:J�=�W~�]��{�u�԰z�B��M����'|c��W�^����8��=Ǵ�s{����3��zqЪ�x�kx@Kc;[[cScc[�뮺뮺�|�뎽:뮾u�^�u�]u�뮺�뮺�Ӯ�믇]u�ǎ�믧]x뮺뮺�u׎�뮺믧]x뮺뮺�u׎�뮺���]q�]u�]u�]|�::뮺���]q�]u�]u�]|�:뮺믗������}��o�]uק]u㮺뮺�힞����u�u�����ƶ�-ό��F �W��S(�B[ϧGF�콢��WL[�ۯ�qKۛ�˃3؏��ov_oL%��~3�4��>d�_?p��L>��ґ��ۨ290���{��1�L#o���uΘ�e/{����M���;�.�1�:��K��3|�������d����֓���-=^o!$��}��f��I�Q�͊��+"������P�Mq�IX�/pӅ�;b\FL/��庇��{��Ѿ߁�,����
x.�跃�􌼞��8��mu����D���k�������{��0��|7U��:��W\]r�7$�ئ�G�=�A.x%)b���x���L�/��=�����޷)ڳowl`��Yឿ}���ynu�4ot��4�M�iDR��>�.��l��3���E��e�|�`�zJ����n��<s$��Aw��Wxd�H$� ��4�Uź����G��+篋��������#A��}�[;�_z-�T���V� y�o����NANʷ��Ԍ{��ү���;�`J{���D��Y�;+Ï+�ͬ�>�c�{�>�25-��H=Ϗ}�zkg��rW-Ǌg�h�& 5w��t��}�{ɱ�rÙ�>�8��2��Y42gho565�5664뮺뮺�tu�]u�]u��:뮺뮺�u�u�]u�_N���]zq�u�]}�:뮺뮺룮�뮺뮺:뮺뮺룮�뮺뮺:뮺���]u��Fu�]u�]u�u�]u�î��Ӯ���]u���c���}��n��N���]uק]u�_ON��u�]zu�_}���z��5�F�(L}J�r��� �&;��nt �_J�2��|��p��cð�~��Ź�վ<�:k�a�}*�ʀ��Z��Ej�a,�B�}T��R���y�s�Vgy��?xv�!��|�����3����yb��>(#w���Mܗ���8{���$���V������3lo�[ȴ3>fg�7���k�`�z�u��h�^YD0O����0�8֓xw-r���'Ċ��Q�9����/e=�U=��}����sy,��w;n6���e#��^Lg��2�'�?����C��c(hg����:���ur/�C7��(R�I����o�	8����*��}$eأ�8NE>\\S���D�fzj�������r�}�}�����*<���y<2D;��� G��!Y�R()=���g�`!,���_�����Y�2�ˌ��ײa���L/;w~3s�w{_م�|=�|� �܁D���?�`��y��ת���>�����>�٧�P�X>���`��UZ�b$g�9}d���7��S+.}�z��7ʡ颮�xY�Ǎ�f�>LY�5x��" �(�N4q�Aɞ=�����NLhz��	P�g�:ƭ��}��,=�E��=�b-M8a���MN8�F]��Q95Vɴܳ:?�/66�y�I5�c��m0��G��d����=s�\�h�z��.ބK�;W\�/g�=~�,�GR�M\
�������f�/6�Ŀwي���,O}��rc�|�����?�V����uzy���I��ޝX��{s_ �����3�}���]�9f�ޜr^�gML��T+��a��=�Dy{fS���wۍM���X�R1��f���A�f�9=����hv-х}�`K��_=�X��Wr9ϧ��4�~�ſ<���~�ً&���n��df<��at3����7��^ND3�S(e�f�pw�j���y5Vq]�=�~��3o=�ս�o��M�����/��>�Em�����ր*Nĉ�w���='��Γ7�ӧ��g;�g����Y���|���v6 �	��RL�'[�Dy��yG<sV�;����Nk���3�T�|wY�<a�o��{�^��D�g��g��O޺wظG��ǯ��zh6���<�����7DY�{D�w�/��i�C�ǘx�^�d)�3rU�r#ə��5T���6g�'��\�B�8~�)n�fϾ��vc"�y�mY�p՛�q�jB��{� :�I�c�;~�_	�"Ѳ_x�6<��ėv�e{�Ӳ���iζ�߳-��~�c��G�<0�����ݚ�Ȼ�?���:���靏[=�0�{ؕ=�xk���R��{��w,��'���Z9��4w�e�={kn���_{�g���"��&�}�(pv � 5�97�!`���> ����=���ɛw���{��)�&u �V�r��_�{�@C��~�4���%3_�%�������׳���D]=�z���'��NK�1I��${�w�@&��ӆ9��tiv'�3-�s�����X��Ŵ��dśd�߁��7/cÔǻOA�A��;�k�"�6�j�T�����T��t=6�s�6x	�αs�:v��s�θ�㝉Oy� x�]��}����|����6q����_6�(�~��65m����{ :��wG�48hXX���C}
c;q,G���xF1�1Pp��v:�/t�<]���n��f�G�ί��Ϯo�D�b!�����Ց�b����>�ׯU�ly�gu� 3">��PK�|3�r�ރ<�9*�R3��r�m �yM�0��;��^͞� ��V <=_#�}�L���t�z���_���Cqe(\����X������?s���a��gM���>{��j�6��8u�� ����Qc��XV���qP���px��r�����Z�\~�����ϗ��xhX��!|k,����ۭ��ݾ�y#�S���-9t��0�����U�H�OA�4j�썶"���[[�o
vvT��e��*`�ۉ����<���=^���d���usV{���͞<�E��yi�벧�����v��i?"\+*�8�b�{�z� |n�#S�L��ѱ��[]���f�����/�E�*QT<Lc�+��;��Q�bqcC�cn�^�t�ݪ��w���yR3�x�(��7����7��\w��/ʷ��ʕD�@Т�F	e���+9��t�gw���S����ޠ��>ӏ�e}��{q�Wr�{3L��|K��/)���YF�˻�<ߙ�v#�_F�8���ܳ�9㝂�k�����O��Wة��-w���Q�wO�g��MSէ��ӳQ�^�gNX�c�'�qv�ӥ��>c[�~�yC�d��hH{ݐb���y�9e�y��ݞY)���y��}Y�:N����ݞ�$^�>��~[,1`�l=.�'� �v^\_ˍ�8�(�Mz!�=Ǧtu�d�UHUt1E8�P�˅uRZ!>� �nvoKm3��3���?Ӻ=��)Ӝ{��&,�f�^�s���y��?i�����?}����{�9��5}�]�7mf��9���/��[�f��mNkz]�}���l {���q{�5��,3.ɀ]xs�%�q9 ��mX��wg����6��Y/������,mʷ�b����ǳ�p$����7�����}P�85����-�'x0E]iC�<<��Bc�WO$��ؼ�c��u�4��XgN�f��kW�����P�>�P��Μ{p������5J��Y�=�9T�5��Ǒy0!����/40[,�r��gL�2>��]��&^�\������<��Q �]^z��3cV���=����o=��~7w�]��>`G\�Ӆ�}�x�n��m��;�*�����������w{���Gf�ۜap����8 G�t˚�)�= qws2j��1���f���;�h+�|�,�ަǚ��U�}ejӖx���7-^�옥1��;�΄����[��b��q�Pϊ�����t������s��|.^Y�G}�<����Iy7b9����9��(�%��n�u�.��{Q�+A���/fgh�o�<^塚$��κ3H���q���_�R7dͶ�y��CG��̝N�+��W(��8�;-��ˇ�^�<�}M�r�[��J�*��ч�g�\�KO��[�"�|�k�ú�f�O�Qg��_�o�� �3U��^���r���#s�|���x��4���=ngȡ��4q��=�n���:�q;��
����~5Q٥f�yX��i�����*g���&�'��m�؁^����y�,��y��:<�JAzz����ڷ���t���<��a�i�˞Y�;hl�Le\ъ��m\��-��R���a�ٺ��1�=��'yo���¹�c���F'�t���=~eh����{�4O43��y����緆�9{v��o�κ �v��W<4���L=��,�ި�T��y�s�3`ˣ۲�M�5�#kW7�}����wP��^V³~['m�9jў}����[=��/(�J=沭Zb�z ��[fW�gU˟�۫�v{�zv��f��~>F�_���n�ض ��cո	��9��L|����x�cq�OY�--��$	Y�=�+�>�蠍h����Ճ��3�ĳ8f�?y�y�ʂwt��' ��pI�����/���<^M�)�/����f���w��8v���8YN���x��5N���}kϛ��M�P�s���v=��l��lʍ�`�w=ނ^�������������u'���n�&=�Ev-���^)B<y�Ԝ��Y����q�����W�~g��'W��Ha����p�?��yo����+���v���E�����뢥�K�W��}E�	h��>��*�^�y.X�R�w�w���j�p��9ӑ1@����i���z�=��9/��n��am�C������l>�e��ғyw�������7��%�l�w��AoIs�R��28#��Ύ�`��9�ۆ�$]e@D9.q1�(��\L>�|v��
Z0w���}��7�ݩ\����ۓ��8n�"Cw����N��Eٷ�D�4=R�����Y��f�Ҟ�tN��f���KS�sR���y�<�,+��ҟx:x��Rb�w�|�X�g����c�;�5��,X1�]���/p��P��P7����Uanώ�=b{Q���^}�E�HS�<l���� w�ۤ3uk��oύz�r����qCJ�y��V����gݼ�&�U!٦ON{�0�[ƿ?v;����h�x�Q��4K=���{�ܜX����T6�����7�wj �o�a����/��G�7<�����x���˱�<����>���`�Ҽ���T,=�5xp�(~��/L�G>�����Gb+_3��?�׼yPo�͌��7�ڻo��Onzc���W�]�`C'��[�g���c�Pcu�c��w|����x�7<�{A��O7z(��ٍ���X~�w�:ޣ����|�qxs~;�S��I�5�}����V�V����!�d��$@X3<c���Ns����?�t�n� jFH���w_��Ԍ=��#��>~�/-> ��V��ᘂ~z�'�}~���]��\�C-��x�ݝ�|=�	��O��* 
�pW���������_�"�����c���	���l���f�WyXLǥ�I��.?���D�'�؅L~1�G) �%�F|Bw����f@�R�`RZ�8��f-�4ɦ#dfZM%^�5\�]c1���&�������C
C2˒�P����]2B'b�KpKB�m�KZ1��&���en�Yk\6�
�b��a,��4m�̈́E;Ii5�[�WL4WA���:�Ȅ�	s�K�[�Ȇn���p����R�� �ve`VYD4ȑy.�[098\�����q�N\��&hѲ�vp��4���e���T�4#M�ЗnEa�{sD��ʝ�q�k/<\`�m�ԩJ�ƴs
0hZLJ�a��2Z����4�2�����6�4�h�i�h3d�Q��K�/2m�,tؘe&���U���L�3tHڿ�|O;��fTš��R�f���ͷ��]�&W]��i(ɍU���dԹ#q�"k�3x�.¼CS7�t�����Hl"˚�-̬�#�m��3L��֤�ґ��ф#,M���ij�4��e��:��3(�M� ��+��O�t��Zu��.*�f4�ݔ��eWFBX�Wfl�Дx�
�!M�K� u]îmlm3��]���4Q��:��Tn��b��P[����Y��[,ū�E1��UT�k���CB8�08f�z�mi,nB�i��Кm�X�j.b$�KT,7]an���5�#휴3�7و��L���(��
�m�fH��=X����S��YM@�pj�i��(q���[[y\�z�a�$ �q�-ʺ/ �ш�e(�D%+����J�ɮj@�PT��[��ڌ�bFP�b�5i7eMl�fm� ��0J�Mj���%) ��=f������Y�LYm�j�(7�Ѝ#�J�ഒ���A��q��rlTvk�֩�m���4�u�͗��KkL���it	��l��(Me��].P��,�t�����)eiU���E�v�F��)�Í���y��F7��cLGL�	�R�[�����qe�JY������x]B�M7�6�[��)ֶ���n,e��Ԋl��V[f� !��#�ClK�-[ŀ��m�s�2�K��+YHs��7K�T��孁m�I�K�b[p��X�Т@�ж��%�m���R����kL,�.`�Y�X�t�v"�eҕx0�K��B#�-"��Xms�J�[P�YLX2�lb���Zbk��JsG"mT
�԰
��5&�H���Rm�^)\���b��p�;i[s�h���]�q5Ĭ4t��m�i��S&pX�ZX�&f1%��ښ�΢��2B���f�m�r�\Cވ����,�ƴ�1�+MH�L�]�s�`7��pEsu�\Jՙ�[E�ݰi��%S�R,��]��&���Pk\2:	yu7�4eibiK,t�%��ຐ3��jk�ңb]�-��u&Yo��������h�2k�ł��k3Z��GaSe����0�̫)�Lf��Ñ�͛f�sif1��A���r����jk�K,`�4��{u1�3-*m�n�u���� �0iE�27G7Ch��s �����-f�U�/)����C����L̝oU���q̮�5��X�0���{�n]1Y`6�mk��Ը��c%G[�v�5`�RYcGA��RZZ�,�{<��Zh��a��ƞ,KZPd�-sFɌ��v�X�j��Yj\TI��Q�-��u��^-�rhKs"B�b2��n���,��������f� �%�LkX�w�)���P ��A���t��Z�Z5y���YrZ,��0[(SM���kt�wm�bZ�V�=�ǯ��G����Xz�q���`�`Må�!*�f�Sh�5��iX�\�Ƶ)k��]0,��cn��u���\�[V��it���4\<�kajVڑ� 8&Ҫ�j�%tBc[\��ѻX�6������-�*�Y0ڈjf��6�\��4إ� ڴ�8��m5SD�T�n���뀰r䎩u�����3^���iB9����J�%�1�+5�h�2h��4��5��1K���CE� :R�`��n�,ԻKK��L^Y�)�^��P���V���z�˭Wc��U�B���$V뛑)l�J
;)�c[h4`CKGZ�V�ɴL���&���p�:�t�E� ;G!nɣ̸a�K�s	664t:��:�j`&h�6%�T�N��[xt%�
�Cؕhg��	��I�h�qء��в�k�u��W�0�jmL�e@m�l4��6�N(�H�)-�!�}q��>_�n&Bd.-1@@�t ]�)+�v��\���G!u�&��3���N�e�����uI�XR�5�A�+��`nƲ����5[�]�`K
V��a#KLi��F"=vh6]#��([5A���$�����ͺ��Gk��Xkk��3M	�yH��kkl*��իI��P��K���s�.��c��mM�Xn,�9ni���U�RA"�e:�*���(֑�F]`�Z��X��3M�@���e+o%��1%.�a��(M,�1a�n�[���]��B2"f��K�cC�M+�b�[�Md�o0�� �m�A��u-�������VR4��kkm�e63m���j�����("�\�J�R:��K5+gQ����@���K�h�-��LX`U�q*̉;Xe-Jvl��1㔲֕X�̴�A�Vf�]]��B�bj�Ÿ�2�Y`GI�T�GVŖ$+hW.�f8%��ͺB6`"�*�.^���o5R��!��Bc]5��.q�6�r�W&#��٩��K+��X�-]Iv�I�4�MU1�U8�%n�*\�����ٶLT6��"K�ctu֚��qk��W�v�k�J׮0�UrLki��fd!a�2Lu�Qf��G8�v�������mt
��������SXL`��vV n���9���E꠴���r��uB[
՚��42I�ip7T��-[o
�����p�k.M-3V�Fl��[��A�����;4�l�8�z������&�f�˝U��wkU&���)i�ic)Y*�jc+e����c b�ٮ�k�V�F�%Ų�u˰m�T����|3J�C
,*�J2òRF[J���ˑDVY��d��J�ҜWf��M��9�ce`ʸ�\i���b;iem��tV�U�P�Jõe�Y�]�9l.�mNYB¶fnN��>v�xH0lƻ4,d-���ܣ�l
2R�%�۩B���b����S�Gru���)!vi0F+��mSVg[� ���Xh��ص�K�K���gb�ۮ.+��B�f��L���m0֤[�5%a�Q!5��[Al��Yq��f�Yr�u.W�m�;g�+"����@���ʹ"�+�ʓe�Qatĵen�و���	iج�$����GeּCL�w.P�P�P4�qt�D�k��]���`}+��X��]eS3IQk,S!�ih���4Zn��:�MZj��kv6�V%�lI�8ū6�]a�P��.j8ju�ΡR::�W9�gM�0M�9*@���Yc9@�׮�4b���`���R7��0�V��Knt�ʫZ����f�5���@�6ju6`2�mvz�l3�Q��rQea2�J��1̳B��6Ƞn*jb�nq�U��jst��$e2c6p�����͆�+P�	i� ��%���vm��c�P!��!���%����]�&e� 9�L��9�[cQa�\9�SK�vL	�m��t���.K������pW%�$`��h-�a��Jd]�Q�-/'5b����5X�1�Ue����Jʑh�Z���P+q)mP-�+���S3LB]�����O _�Y���ᙰaԴۆ7X��Z�m�,�aȲS�],B �/��۱�+�B�A�!�m�e+r�-tն^+sx[�*]���L���b�m�3c��d��ղ�o���Z�e���-q�jŦ�*�$�8�Ka/f9��A��i��6,Ŧ���[�6h�0�k�Ԙ3Xe��.�����G�e��Q��i̱B��j�Vi��Վ-��aA���fl�#+n왐��G���*�Еu �Ή� �q��@��/jZ�h��&-6д�hB�����]R�������u���C� ]�ՙYn`��E;�SX�r0�n�e�XhF�9i��4e���6Di�M,�lЫT�F�8GCٕk�͚�Uhn�G�1%+���-�"�y[eJr�X��;Z�ᚖ��2q�4��M�`L��R�&����
�u�ذ���0��/c'͐��n�2�V�7��h�Rbo;](L�n�3�u1�!ttLՖ��]q)�J�t.��)�Z�5�i��ͩw)Und�­��
uz������ޘ�[P6�V8p�ŰUי�,���ю���A��\usٌ4[s`�8��6�.�2l�J�g+�5ѫ�	��<U��UUUUUX0U-V춃�2�e���6.S;SA[a�.n�/בIe�h~|f}���A�p�g����n� �Ǳ��M�.�f�ы$�R`�����-|�,=�n	�}e#6[�+�p�È��*����dEF/L�V"
��#,-�Tb
����**�U�
Ҳ�,�w9996t����^3��lDV܂��=E`�ATUR(1R2�("���m�����fK5���|===::�u�<:"��5DOkcJ�eF�PUV"���֔_i\J�PB����:�Ǐ�����zzz{�{x��ǌ�;���q���u
GYp�ig��Y-� ��X"B5�%h��&K�BQX
�
��u4l�[dR�AE�h��k�L��
��ڲDH[o- ��V)2�I���6�й�A�t聆��)i�%�����m��.�)�p��J6�Z9ә��Iq��T�F�F��|�呶�Y`fH<HYC�B��p��Qb2�B�3%2���#e�����xyx��g���<í ����(5yˌV+�y���Ԡ���u*"V�����َ(�z��TXV�[!`��ϳ��M骊����]@��e�����R ����J�AZѴ���Y18���J.Qh�Z�-+�zj�eb"ʊ�\����"b����jDj^YEdW-TDbUۂլ(������޹n�m�ؗK��ڙ�Tҹq
���1Q�Ѧе�`hbat�!6,�:�ؠn-r.�֫3�����k��fT�&-,��2M���J�0M���M`A�K���ol&�m���4����#R��]�ietk�l֊)6��Kqr�cN��#��il���i��l�������7�.����%	�͍֖l9d�Sa-��}�{���j;��u�����権%Fe5[�Ű�ij�XX�hE�"h���L4�fj�%�Xɀ	i�5����¸WH�@��r��Jf�K��A�d��1+a����q����Z���m-���+��l���Q��c��P��:%��rsXh�)�-������n�8�PT�)!D�#5+�WcuQt��E�e�[.2�-���W�.���+�ɶ�	u���"j��(�K���:5 �-pI�e-�ڀkb�ʁ��
ѕK5�]1pe�.)F��o���7S�P��$T��������6�mJm�YX�XL)6j�v�J��wFX��)���b�#uk�iV��`�Wl��V<\��,ԗ����X�p��j��mo[4��[�y�4v�bד�Z��,3�a�e�]��̭��iv�eUy��8��䈫�h lQ��h�.q�Q�)(q5�����g%�Z�M�6��Ƽ�T`"ńNx���0C
�H!Ղ����+R�K*,���#c5� �4#.�5��#*hKB����mWT�[��ō���Kr����* sj�SX�.�6�� ��(P�dYfr��e�����E�
���-����S4p]V�2F���D]J�݌���i[��Dnb-�Y�%c���WF�M�n*&s\5\;g	�)�6:�����3��$�q�ƹ��eZS��i-e�j��vcc�-�-���+d[k*EC����,-l@�iW�B%-TA�-ZK�b��HX[^hB<	H�,�h�e%[�	#Ũ�,+PJE�Z��D�IiX�%e�hKX��V�4`Z�F�BZ��Յ Z������/ۮF�J�MK��0��n�����ٳ��ck�n2�����=~{$�|�<�W�k ɿ\����D��ey��h6J�%&�@L�T���6���'<�)^a���m�z~�R��JWӗ�ԭɷ�X7��>���"׮*�1�vv3�q�NYŻQ[�o�y4#*�7!G�j�5���	��@��,܏�����j̹Z�g_1��r��1�\��UN�f�i�(�&��z��y�4Co���(���X>��0�~̒<���ݨ��M2�L����P9^{|EC���V������l��f��D�v�[�4�!oVhm��4���������^ƻ�Mm/n�^C�L�fh��7�>�xf�c�m &U�)��Ucʕo2����J�/��p�$�䍓:Y�4w��p��f��f��.�Y���p.�jG5��l�D�;�"�4 Ή��r�z�u��eg�6��4�U)���,��AC���|�Nf����'����*9��Y���5��zк���RP۫�&Ρ0��C
�fyC��^�ͼ����fk
�&�J���g���a�7<�ԓK6��]�v�)zFg�F\f��ϭ_������V~2[]��Oԃ
]�}���0~S�kr��0G�Ռ��2�Vlgl���cq���*a��p�����-)˄�����:V�����O�'�^�L�2�9Dԑ<��{�#2}9v}��x��ӕ��T*��&�C]���Efޘj�oM4�&��<�;
�v����j�36��ro�|ݫ�+g���{�O�1�,պ;���g�x�a�)z��͝>�l�,�DHw����u��3՚"ש0�M3��c3l�G���\���i�[P���)'8�C����8����YFLٝ�G��1z��a2˴	�\Zѧrdf�M��n`��yVKfh�L�Z��;L�:�v�zv 0���Q��ɴ�	����k*��Z�{p.�����h�t�]��}�}���:镇�=�lf{v!�M^g�7c|�U|F�<T�SU8MT᪐B�uA�y�R۷	<]��״:�ҽjf�r���òޛ ���?]6��~��"�n=��]�x����L��F��S*e3�{]���=�̘*5�"�7^���z�@�,�}=�zg�~�7�뜧����ؔ�|-�k� I�->���\u�����Uc�2�V<��e=Y0�)����e�P�	I�ss�h����C=7�I�H�,�j'�����8U{��V�,��>��&�V=6�F)�w���w�<@|x}��=�fk�1�0�/&+�]C�W��XI� �J�s���i��0&P{v�f����M���7��Z -�45E3�+p*�z�i��P�M�����y��+3!�%���6��%��4�mbu[;Vñ�L��e	������f�?�nh'�C�ƙ�c9L�a*fh��s}:�.1�!�-����Ef����sߧ�,9^�����O����5���ߞ	R�ћ��R*�m	���͍��q����y�=pPzǻ�v��<��P.!A�a���^A�V��)��hW�O�0Mz�<5��<Ƿ �6��=ֳ�{ynw���^��)�<�E����[�X�e��4�L,Jz��p���+��M2M�S3R���2�ţ-Jr�[-vnڈd��$���r����n���.ш�J��\�mZF�Yf(<��;!9JU�4�*\�	�a��XgkA.���B���"��,Ɩ�̰aTJ�Y��C6E���͋���f������1#xh7���Vm1�e�A��H�B����}C��\�lm�MjםDl��cF�����E������i�Vx�����m,���5]��.=��>h���m_�y��\BH	��̼�K�}�Yb����N���w�_w'����-��������ž'��I8��c�*��e�<X���+=��+s��e�d=���
g�	�\{���2�G�=�q4�3�i��df���氙S/��舖{3��z{3t��>9���G��C�����5n�4�y�9�ބӴ�*�y����LDd����p�0(�iз���p`�]f��4����&��q��ݣ����7{]��D3��T˿g�G�=ff=��{�wK+Bʏ\m�a2�4˰y�q��:�? �O�1��p�߃��B�& I£h�yu�އ��1'Owk�o�y��ئ��$�\��T�ɓi#Y��8���0����F���2�r�g$1�]��#�0N�>������`�*����zL���/걒[2#@�����-vB;��j�p�Q� �����}j�;��`ڄ������-:'� Ey��La&-2�X�&I���CĻ�f[���}�Fa�}q�>h�v��md��*�C��x+��S�߿O�Opb�iU�r��X&��s�"G�#q)�Y����1w��ڭ��S�5ͽ�Ȼ�MY�w���5�S�g֪yoS�!���仏FwI��3Q�%�?�s戴�Ռ�T�6s'^m_��޿!mv��#���^T������;�=�qH��~7�G.\�.n�I_k�q��;Yכ(���^��;�I����Q�⁫�dYf�f`��x�����#|֙A�n��U&�ICcg��u{nL 7ɆT����x���0k����w�z�u2�Vs��c|�	�!�PM3mU���q�u����]�fƅ:׹��A-�S)�uM��I��5)��i�]�	4%ե4�Ivt^�F��l��Gk1������ǁ�����m6����s��E�~�`���W�+Щ���.��`e�5�k�4lg�o�3/�-���Vn�sQv2,Y�L�R�!��	��8��dS���.L�i�g��f[xVWZ��+G�/f����Rj�j��g6_�拥=H;n�����qxaB��Q�1��&}Y���mϤ�ň>*�jN�M�sY��㴏}ܳD'=�^�:P����㟦{b�K�~ד4���'����K��˷�v6��ꖖ& �,�c33�3���6���7JOYc�G�\R�v�L*�'�o[^4��O�T��:Rz���~��b��h�nn��$hQ��$Nr-1���jA���ܞ��?=�,Eid*T�����z[r��6�����o�氾���r�i�V������s��&�umj��w���b1o��l�a�9ow�0{\�<^?_�i�O�j}k���٥VmK�{t����{,gɃ�9�����ֿ����M�;�sa��Z�/�~��s/�Z1z�%K�|����8��rӖߖ;��@3��M�KW��TY�/�L�뙆��+�
�W�^y{y!;�+P�y#އ�w{���.r�^=��W��u��~a�asۉf���22}q�;��\6ga��ZA0��C{���n��F{Rx��������ei1�����c�փ����d�b�К�ZfU �Ζ-m�4u!�֦SX�:aD�6�����bZmp(]mf��������۬Z�8)���KIvn��
"�f��f�kYZ����1�������Y�Xh�l
�glcTb�3�G��K5�Ñiu�`��+��j�P��֗:�]*hWme�1�bm�2m��Y����O�2�	���VKu+)����gk�Ra�������-�S)�Iڙ��n�QYc�Z��?��b�	մ�>֯;
���Ϫ���wM{a,��L�F��)ƹ̼|���JfF"#a#�!��1�>R� v�v��tг=f[]w���u�1�����8�*��Q.�������0%C^8�h��{jwۮT��Ǻ��衸��l����� ����⾶{"ż��v	��������A��F������e/M�O���w���A��<�����%�Y�P1�T���F-D��t�P3�c�_{�x%�0�2��Y���y�?���w�5�orb]��;^��+�H2ԡ���;���m=mDE>�*��?����uV��q�C4����x�ds}�����F;�E�xz>�f��J��� }�T�V�OWYu��Sv1�z������aXnq�� ,A�}1^CZi��`���^y�=�+E��Ȭ��F!�BS�̣�^ �įۜ&{�_����YB�;���"����=4�X&'7��Ŷ�;�L���)�SU��N]��m�+v+7�T݌y���Ҁ�ȹx�_{v�yCE��h��%0�#徧�Cq*]��3`�3�5u�Vm2��!��f����V��1Z�-�2�&b�}b%`�9�z�[kr�"�L�@�ƪ�U#�������m���:|�WX��h^�ko�RM�����	�oZ�U^�"�
�Q`3��-ͻ��N�o~T��E��S:��=�7�Z���Y4���)S���Y�bܮ���^�S�A튽k}�3Q�=�[�o��ˉ��^)�����o�ۗ�X�g���ۤz�^�f���kx3��}�����>L' =����кu`�]��v�țg��i��J�+����^��,�6�ɓ�]�wC� ]�ʳ�Fwe��]&���˒'�Z�W>d�zgl=>��S;��������<B��s���wO�ɥʺ�����o���û�>G��7Zf?8��艾��<�ʇ"+l32���|������|����Q�c�l�▄�������I���7˽ò�!��.O��+X�y��wp����4c!��o��~Z�N�k�/r�\z7�7�ҽ_&:�<NwG�9�����6���;�����6�J�H��x�t �����H�1V.~��3�[���y}ɼ��w�5 WM'��/�f���T=�>͵q��9:���K�8���Pt{��|m�a�����{�`^�)��͜�ܸ#�}�sx�꽮 ^�ٳϮ���	
���yo�a��.u7������:d��D�AϷ�<���}��&b�!g`Ԋ{��<��o�eŢĕ˳�gl&���MxX{�V��L���#N^�r��z���VÒ�w}��|�����>����<3;�����<��1�a<g5�8���w�$]P�Y����!����mX�z�U�e�&�[cf8(֊͵t����ȍ/a�ss��*��=8�|>�������Ɩ|F|$UQO[�("�h��5�e�<IS֢�V	o�k �gӏOOo��������{x��u��O�c�
����1TX�j,-��U�U[l�
��B��IF,\T,ɳ''O�����{���<x�=������dOY�1ADb"���Q�Y�Y��V����TX1\�\��Q��E� \��
��,5Tb,�hd�X(���Q�T�1��b��N\N�D�IUX �U�T+a�,9j"�mR�2�(DC���B�]CYm��k*�"�i[hc(��wvf�EMk�-�Z�1�J,SR�A5�Qm8��EQETD��V.%B���R�Z��-Mk�[Q��(
Ke�4q�gIUa��T�f2�
�QX�%AB(�q
�>N2.�J���fP̢��u�
�Ȥ���0&ҰX
�8�WP��v���W`���ű�b�1b�
d��������=ϡ����Q�t�`��0C��T��
�p)����'3��L�&݃�&݃�5NǅW�7�&q噐�n��1aWјLlͳV�A-8!�Pj��� ]�v�ݦ림�:Un��i�`�L����"���i�5Jb ���`�Æ5N�}κ���=�4>w0 m��_�w);��(�Y�K�Xт35׵{h�XGb�e��v�������A�@9m�&uT�85HY������뱏��mp,/�����`���V�؁���!I0v"�݁����$Em�,3���b[i3��{�$�-����PN�@;K&
�Ő �\&^��)|��5�0�7�A(aX�H�;��;�I�����V�d;�Wf4/k{x;jPv,2�pXU;�4ɍ&v�s=Z�� !�k���\���f�@8W ��j��8[׏�������i�Ї)��6��(�b�Q/��1����OO�ǚ��٫FM�}�tvo�F�{<�-]{�����3m�T����ǼG� kňbň����I���:����#�t�
� pEQ`+E�-�` (�z��cгN+W�^-b�@D�p��NX$<n����R��@�b
���J�טA��ri�K��u�U��͜l�L�M��r��z?��9Lu�2!�t��;�{��>>wYw|G����:���O�f�@z�4�m,Z��85I���N��R��䥙��Gu9`N�p��3���b��1�$m�p
�O8sT�hه5R�`��z���9h8,�p«�XU&�|å����wk�=4�>>h�7��l��p���T��5j2a���g������zA�`b]�����N�6�9z��&#�^֝M�})�nm��S�t��L(��p��<�q,�H4�� isT��~��8wC5�pm��wZ��u�~a���ᬘ+��>b���'�Ұ��Z�yQ~�Q��\��=��������Y�;'�>����=�*Ʌ��<y?l�z]�ߜ�=}]�f]��T;��2-{#!)�6�O��A��Y�ʗV5�[T�'�N8�q��Ѝ�Ʒ[�e�#�3�lJ%��Z7�X��)	��C!,��;�S�� X ¡eYSL�L���Wmk`X��X�e �7���lq�p�[�MJ-���6��=J����"�2�@�ִ�
̓!��[�j�;��,%xW�<�aa��@�c7Yu���00۶RZ`qE�ku/8^l�eu]!�O��ߺ��38���n�NLCh���%cTia7j!U�4""g����> n&g�p�ۇj��M?vI�-��||�3PB��~1�����y��;��C��wD(� ిGs�cՀ�0�Z@�(W8{�zQw�L�"���v<�0p|�{]��.SK�c�D����kю͚�x�� ;*��*�giM���P������8��]�}a���,@��v Z��5I�ꝃ�!w��3��o��0��x0��y0�8�];���p�H3��{�$��Ws�vj�X���[bz%T�Jx`�gb�Jb��}� T0�L�j�n݂c�=�^TdH��%tc !�d;�`��>�i5��4�3�&i��!�Ia�p�T����&q!~; ��ש����۩�����,�R���q��3ڴX$d��fۥ�n���I��1��膏�\|�i�M\�>�FEǮ��0�M3b�;)��~��u�C����t���N��i�B�X�!�I�A�;a]�ݐ��ʯ!׈������#g?ë��z�P����u�ry���>��r��i�-�fx�^�BZ��33�~er��}1�� {��.����&��5��`�����f� ���=�sT���0���������<��_i�������t3��ε�Ͻ���`;�UDToq��t�֝�i��N!���8�M���C�dyJ�&��l�YRᱣñ��BU7�v����[�t�\z�p�\E2
e.�s��=ѝa��5�u���ٮT���cv�1o�5ʤ���Kƀ����㑹������by9����'��Q��/1��%��%J% �	hb���J�C�[R0������J�X�b)Un�S͚�!GTg�2�0�	� ����Ӡ����,z�./4��$��L7Ԭ�=��Ї��a��l�ȝ��9�\��]��o����� ��{���6��gt�\z�u���fPpX]+D( ݡ��u��#� �C�A�1Gu ��X��lB
݊�բ3L���b%�r�J�qV���q�[q3�o�?I��՛��ί'�'���z�X��e����x}���!� ,[�f@�A����p����N��ٯ��LXf��v���v��M$��r�<,�����������/�>�ꈸ���O"=���7����O^�Á����:vY�] *�J�2�*�
�sV�3]_����<�z��;�*��Y�i7yL��p�� ��T�Ժ�d��e
كi9pS��Ex �0��6VE6�ns��M�9�u(��T���
x���������,E�b*��Mo�=�K���|���F��e%���+� ՌDr���RBdZf{��s�;�Ng�8�'�c�1#9��Sw�f�Q"'�u7���p�ES�SIWF��h"�;v�/
d׊|��8K���,���RB6�������z&��Y1�ip-� ��X��5H8��]˅{�>�é, f! ���؎�9��"hϮ#r��O�z��
�����u�g�W���w �\�T��pD<^�ۡ�OۛGU�H�>������z�9�Tc�v��sЧ�
�n.���缦{{1�����'��ec*D��JN�M�;��V��AC1Q���s��y˸ʑu���`��Cۇ��T�>��Yy������B8��4ᝍS�cQS+��3��֥ �w��p��W�°P�nq2�16����Qk��h�9���P�b�B�|)qm�pF��x	�O�~����>��˧ᴸ�7��d�X \�>�`��>cT��5H��h�emt<�G�؍�g�^���.��׋��'�-�g7k����v!�*�)�����k�fݪ��"�U�א��z0͌�.����p�Dη��;� N8pDӸ�US��eR��жm/z=X���jA`v\
��cT�Mߍ��Dw�&2��m  @n�b�  ���� �f ��p�ک2P�p�����������k0��;�T~GWA|��K+�A������j�����R|�������d�g�n��O�̽Is�;e�=��2Y�uq���~��`LnE�g�]�WG�&��e���R���S3ׇ4�5�~��N��kZ�&f���$bF$��@���ｷ4�A;Ct�f����c,6�^�4�
�\�	fH,EB�6�gQQ�S2(����P뮊�h�
J� i1�6"k���3�m�ʻR�%q��1nC0v�^E��U.an��Iv�tʏ�Kh�Z�,�Ck)��$��cHۗ��J�J��F\�R�2Ubb�4(���m�&ڤ�I?���?Pv@��pa5,1�{d��%؊�]WkS9#<k��Kz\A�*�A�A��>����F�L�{y��ߣ���Ok6BA�p��w��A�ݜ��Е�"����ف�54V���y�������U�K�{�;D�R�z�9.\�a]N��-A4*����B��i��t�TS��`ޓk+�>m�����b yݜ�'b	�NH4��unVF��m���*�Z��US���bcw���
�oo0pL�Ë�M���A��L��R� �T�
�X >P����C!/C	g$'Iڷ<oyn�z����eqoy �N8sT��S���;3htR��7�VU������߮���Ӳ�����q)�����lvpPty��	����O�Y�O����w�
�g+�Ƭ�ϟ8�ށ�~�$O`�X!�L7��9x�
���
�yT���Juy۾�'�W�=]s���i����~\wƞ��|�wO}8�=0Q��9|�_��g�e���{��ꗑ˼�	5I�8�rR�0o����*�!i���<���:��,T|>�fy������ا�UM\�ȹ�Z`-fl�g{NjpAi�g�9�6Ε�f�Z��t�h >?�����鵣eq�y0v ͼ1�eT�1�Ñ4�8z�n�����u��7��z��wr;�{z�o���z��;1q� �r��3`NE���l};ˌ�ˑ;��#�t���pj�>���>������`z����b��7��ñ�B7N׃��p����?}
J_rw�޾w��m�CM^�@V	��
S��n����v�v�톃X�n������}��A����}�pm� �[�������y���eqG�G6(������x��{ܒ@�����f�>��Dҿg��o��Fk���x������|���jwmg5ݜ�.��92�y�B�8��أv��n�;&�pA�q��V{ہ�@���Y�;�u��O5꧜�>�z���VU�jm�\o�����z��Lo�+�S��)��&.��)ǽy�5�*\�0�.+�rE�
P}Z$=p���LY����ౚA�2��M�.ݝ��ڀD/{rX�|�e&'!xj�cׇy��'#&߆��	��r7ո�۫f�I��A���N�j)ç�|BB�A�"1ÑU�]�y���f�S���^/������8�E��L���L�*�옊��F�$�
���>�'�6��k��em�FR�JF�
`��k�����S"'���pD�2nX��g�o�ř�oo�Gh����ݻ����q�C�2gP�j��A�NFm
��dwkD 3Y�O5f���DK�M�6�n-A�d�p�
��=Ε;Ο#�-�`Bd=���T�Uy؊�n[�tXޓOO\eM���9�����{S�k��b��)����ź�9��?�^eZ�9��9� Z���P�۷�b��7����������Nf�.�2�F���G��]��Xdf����d�C�C�TJ���T�ӗ��gA��aU��z��r��M�V<{��?��˄�|�"0rD"@  �����g5J�2�5Rnk
���%�$kRq�;s������_�l�AۙՏ�1�1b�po���r�<e̢��³�ωN��v�A4�J�J�Z�+�Ű4��LMnԆ�im�C����,�p�U;�N���9}�l��n.6Ɣl���Aƾ��Gbg;�ZS��B�rT��sh���q�yf�`�� ����u�ϻ}&,��{P��v��r�8]�a2���-�vv���p��|�A�ׯ�fo�0{�����nƾ���5�~��?�����Pܛ΃�&Ա�:�T�Ÿ�
	v9��ė4��y�\I�ñ��T��Z���l��{����Cv'#�b����hq{��R��^d*�J���,���C�'�͖����b�Ec��	�5<Ӽ�j�pA�p*�j���0Ɲ7�A���x����?��yt�����Jn���ٓ���f��Ď�q�&��Ͻ컴������pz71��=��O��9|VvX�=���/2A�Ot�Ǔ���]�m]�_�5��5λ�uz�SՏh96�5N�;4����׻4vš����:�`O3�t�>�y�^\S��R}�Mx�USy�t���bvg��?
_>�ZM����0��,V
���Ӝ'W����>�qڟ��ɺ��������=G���a螣ą}7����W������-	�^�U$�>t��xm�:��*��(�Y��M���q�r�&mb�;�=zz,�/p5��˳�cg�9rল��h˷C��,�x#�J���x�-�������q��l�[V����5�+��̏���[�(�O{���j~2���Rg�:�H�]����j�}}Xx�8�����I��\�A<�-5P�m��}��x��6��o}���Pu�\�jo�:c�~(��������L�@�����L'���#޷���t�����i�J�f{i\�}�·�Y�j�_|��{�C�ؐwwK��n5�SvA�ר����������4���W?~����d�aΨ#sz�y{����ف3F��7LI��Y�=}�����$��w�z��<��]��|�����8��]���������ǎ`Gk��|:�,ǽ��%�xxR(r��/ߚ���ɿ9�R�gi�L	���M�b�S�6�2tOx�`Ԩ�ţ!?�@A�O�AXG0���m�eh!��:Yt�� k��i�v�Z�C��T;bԎlR�0�e�ty�5���w��0�PcJ�d��m�d�b���q8ʞ50Cm���(�CSs`�����V.fO8�d\�ɜq���|�_/����������Yӹ���IMG9Ȣ�QH�Z�H�bRb��3,��X��X�Ҫ"1`͜�M��>_/����=���x��w��n-P�)Y����̕YmF6�J��Vj�sv(�e�N�Χ's����{����>����("��O)d��1X*���E"��L�����Q��P�,�DTiQr�z��$Yp�DQ#hW�W��*��6�![hT�J�0�*�"�F(*�T��*�s:$u����Z��De�0��,QETDb*V��!˘�TP����dQ`bT���"[DdcX)��r��CQ��
��EPEDb8ױ+�P�(1�" %,��� ��jJ�0*��-��V'� �ņZ9e"d��������ryL����J�j�E������Yb�d~�O<��m�n�G��VF[nAm�6�)4)�6���p]qM��}��m�س!4f�R�e6��X�ج�� e�g,ҥt%h#�v!cz�XJ"�ڍXa���{Q��R!3v D�͂Q��,M�r���Q�Ṭɥ��l��%�MwC����X��5@ε�����+t5,��bE��12RCX#K��ai1\˗�[��D-%��ja��m�3_1fۙ+(7�X�n)J�����M�f�PVHR�o7b�V�.�5(Ͱ�56�e��bZ�hm ������[�غYT��f�lĺ�"k��Q�X�Y����Yy�bז�n,�u	'4`��$�8N�,ıpy������Ccu՘X�����5e��	yV��e�Y�+�a��Ԃ�s�v����Xб�H5G[���mj�ݮsX�"�j&bۍ���;h7q.��q2Y�N��C\�+l4��e�,5���݆]h��0`��,t�j�u[�Iv�TI�	��Gi�nft���]) �;Ra�^�]+65����hG�c�Xn��A�#B+4��ٕ5!3rB�D�Ke�b�e��CL�6  I��b�A&Gbm�09P�0��3I�*�+*fKs��U%%f����a��6����tY��n�@�lƀ��]ۋ*\� �h�fbhbR5��Q�.���V\X#X3-�e#	p1b��q���9�帽e�k4Y(��Уf� -�	D+J���k�;iN�%M��%j@	y�[p���g��B
���F
�l������/����k^������}f!	�m�V$�m
v�wf���V�� ݄�dE�2�����fХ֯0j3J�Q �U���Ê����i�K/Q�b�t��ark���Lݥַ3R���QF��5ع��vE1�4��k	g��1T��u�9����N2/Eb 
�H	ǋ�N֗+�R�v��U��Y��1�u����d�XA�b�%��]2�e\��^�d�����f�@�-�20\��[;Ff[,�jf�]��4��u�#�s.٘���r�%1@K�ݭA�B�s��kK��VkR�,��E-���U��uk5�l����v�,�Bڙ3tQ�0�
CC���?����O䪊�Q;)���(�&��ųnrf\�,��
�~}�z����<>��y�ݧ"��?�we{s��=U��	�����7���qE�s�����"�ݪ�&.������l�Gagv=��#�ml`�;�
��W	�NAk��lW�a��� �i���U�~�����D|��}�����N�<�="=���1&�y�x>1�����'�a���ь��Oc��S��1���ui�g��q�;���~7us�N�@�y�ǽ�c&=����k<hGc�"���4h�,S�UN��&gѽ[�"��'��	�pU7�m��A)95�#��N]��b�x��;�~
	�˸W�k���c�3X�Z�3]+��cۗDA�͕ۇ��?_?�/K��}q<���H^��]���j�Kbw������eevٳ�y��1�:S=/�3���V���m��VTr{��Fmz�-�s�B1�^�����۵�`۾���'*�Y�2��e]����"30<]�\��Ng��ް�@��#!#O,�`J*�(���dW���>�=}_.
n���c�e�`��!����q��EZ�C&�b�8"���Wn�.���,Z�i��l�Δ�o;57������T��jӑv�=s����F.+b����-�k�<7n���Wo�ݞs^��M�C��7O���z!�U��2�m&v5J�1V�T��@f)��>.�����`�'�}�z򻃩�����h�8�6��R��D!Tc�l,΁7�Yo_|��D �lP�-ź��;BW��]�%U"�ٷk��	�������pMr�\9I�����K+c4���Jo;5q��[B6��r�E8�5I�ER�"�Iݠ�zcS�tD>��e���n��k������T�{x8&�c�|/\��f��;f�`�)��c�%;��]������9�6q$���Nb���Nz�����%�V��[�\�S�)�B3�P�X
>���T2�� ��{K���x�Ȫ\�>[�S.s0��\e�i��$;I!�a�Bx�"��ϋώ�ߕp�73w\6W��}�6����S��B�8~�O���U-C;�X�Ʃ�z�w�3O
�������X �,-���=��O1�"e9̢	b>he�uy�ΏMV�����9��x������ �&�8"�ñ�v~����'��{��x�kn��u��#��չ��nch�r�GU�t�n���3ux,��Y��.#:� �^4�ɂB�y�1���uJ��ᴸ��u���Å�Yo�83I���az�s^A����y}b��V>�b"]ص󷺗{c4���^��6!��1G���Fbgc�sZX��:����:�'	?�r�	�A� �8pj�[��W����R���y�~s!�y��; ���,!���r*ݝ�۳��Az��w��_�'����@��p׋U'>�1{ӡuJ���:��e�.�9�uI�s���>F�|��s�E���ݩ?Ӡ+��$�3��/f�^����:��!�(p�%�s|�[���v^_}i�>y�͙�3��@O��Va��0������E�װ v�	�A�U8r*�|������r��0h��~���1��]�����NA1h��\wҒ:@�Q�l����&Q���6!�%E���kI��GY��-3�,��V)�xKKm �v�1�yU =�.��o�{r*�[ڃ�M��R�A�" ���%��;�h4M����f���L�م�&ڀ1I�k�bb�E�΅�*r�F����c&���^cp�{v{�U����-��'�a����g}���^�f1
�ڸ���c�]m����~�����RpAq��Rs�P7i�ׁa�ٹX3�C�u!L)�L��ck����szUp���������Ʊ"^���fUn�v-t�U/1�'b��
�g3J6}U�	�UQ�ёݡuJ�]h�\ ��9���	.�h������r������i�
��~�!�����rػ��o�Q��%�;�%�pWH8V��+s;�� �� ��1�v������j�� �0�	^�QhA��F�U�d	���k�=�S[�k�P�%�\5�#]n�K�],X�i(�E�.AmӴ&ͩ][;�W.K��2cM��9�+6Ԇ^n.�kW-�nC0MfƄr���街qiM���.�)�:ts� �j663a�C@�+D���A�-m�ͮ�A��h$-�T�l�ښ��ۖ:����q�5����?>��Z~~jsSJjg�H�[����R,�`P���u���3��l�Ld�ݍS��mv�����qy۫���˥'��_�8 ��g`w����U&sT��5+�}T&+ӱd�E�����jXW!w�w�f��u��i�8� �f�9]�ٓ%K�gV����'���1��+��hd�L�S����>����Fs��s�'W>�D�kk�A�p�]�����Z=U�Hxz�8O8v5N�='��d���x�٨�<}I�둱��<�rWɣז���~�yx"���r&�8sT����V���8:�Ǭ���n��/��� ��wb�q�@�p�M&v�vۻ|rt��1�t� �Kæ�8��I�a�-y�b9x�e�+��ѕYb�p�n���/���~�	�N"�� UI�ד�ͥ/}����Փ�up#|��3�ɋ��gf����T勈�Ap�h��H�p��_u����=��耬�z5LO">��=��Ӡ{����V�#�\RE�]�!��?qy}O��O���١�5{81�ob�\(���߮)��� ���FX`U�aT�U]���p��mY�;����������vvLՅ����az��m8��2�5�=2*p�z���5��ܶ{����k1�碧��7��X�P�i���)Q����Ņzꮭ�Lᑱ�ò�r�� L�vz�IM�Q"�xI�@�*�e�w"�chHvXl�e8�@($�5�!�m�"���Ǵ�8L�Q�ײo�=<O�9��uq��NAmXE4%I��(�P�R���=9�������� !B#�ڃ�K+-�8�t7Z��\�4�n�L���������Kd�(8V�� �*�;ub�}�y�g������?C�Ϟ����5vt�B�9���Yh�$oc�0 ��N
�n��؈�J-)�!z�X�Y:$�3�2
qÃ���-���l�}���F�vǡ�ヱ�la��G���l�s:8j��2C����{��o�}���M>��M��E�֋��4�"�1����+�j�`X��L'߀φ &��2�C�0�'� �ܯ}�����^vj��m9p�5I��)b(� 7�vg*�zd��v2p����b�}���dEO4�i4\�[�z��(��Ɩ��$v�ڂV�mYj���ۓ���}��2Ս	���g
;�
dREb�͗ �5�	��@W��SN�)�O�u����l�6�2�nsa�َl���XҎ�&�ٹ�֯hpX:[�����")QC�s�@�s����5q�0=�_Т��2d,�@�N]�5Iۙ6F��B�[�wnu�Q��1p|x���w�^U�k�u�<Ӝ&�gX4BlK	�)�9���Q��P6acIr(ާb	�NA��R��R��N*��ø^	�A�g0��ɽ�8���A��*�Ǽ(]ӈ���GT�*}C-�����vv���~���������mӀ���|�%�������>c_1N����FYqB�� u�y�p���|�W���[�L��s݃�������N�z���IT�դ��B�O�0>��('x2<��E�Q~<��%�˘�^�\��s�M�ri�R3�������4hԇ�.�9����:ǉ�i�p�H9�2��ם��]V�k�a�Ч�r�\���������CV�t͓+3�T&m)��i�䃑��� E�>~��A3��AN�A��T����3X1�&c8V� ������XF�A�bAN4��H8!�C�*�A=�ES�S�=M��R�7�sW����M�b�13�T�CR���b�O����62�C��޷n�S�uD����ƲW=�Fc�u�\Ӝ������ñN�S���$�z��E��"�Uh�Sn��i���%+~��xʌ�Z����5�XO�c�W��δ9� ��p�OI ����T��S�o �0�Aߤ�=�1�;8�����]f=�j�W�i�9��j�gcT��n��^�{T�ZR������4,�%2�&2������f�D��*��~w�]1��Ɑȶ�w�����N5~g#���ûϰ<F��)*vMhj@ Ko&Ԭ�a� $2BR����ON�b�����1��B�'.he��gkJi���5&J���*.��YD"4J�ib6[��˪].Ѻ4�)�&]�,���0&��(K1Kj0�lq�93������H��4�vwU���]�W� ���һK�X�e\C�U�#%�������V�XD%J:����\a�T�٩4sdF˳��"��>�/�~�5'�R`� �v,kqͶ���Xm�Zj�1�^�����g�e��2Ͼ����ke������i�n*7l��&����=���L�������9��{���h�ॷ�mc�N�X���{^O�}�Tf��Ja�D�g�0j�����W�׬\'v���A�Eۇ]�������X�g�n&���t������\Am9b�̪�b��@9i�q��O�%��ߐ�g8pt�p�A������tr&���l�rtm�vßh	�8#ԃ=�"X�S��d*��iQƩ���j瓳ϩ��}�Q�(�2ܠ�A�p�Ѣ�AN�B��zЈO�T��ї~���к�c2�
G��E�r�Jl�����Lѻn���n[������%=�'�8r=n��VC���{ޥ�`������B�y+�j�NA��qT��Q�����^�Oq9��т��?�*������l��o��.��&�U�RV�O<�/�S=r_:��XN�\�\yx����1]�O��,2�eG��r@�n���������ǌ���e� ,��obLEJ�S�0�j��Gp��_Op�5���q;�����S�T�x MRqp#�V�*#I�Y���w�>p-KH�}h�4Y�S�U��9�˜�0�8Y�9��ӻJ�S�����7zU^v�nl��x�{Dr����5�/'bӎ��i�&�0r�,���E8��Q�p,<k���^�v{��.���6h��	��U8��:VD��V��gH����2����ݶ�j�n�l�;� �܄ ���a�uc�.�k�h~��%��d�����G���������������>�V�ek� ���� �8pES�`A�E�/1�|�b���1�դ?]�[۴���*��P,G�q�0ϯ�;�N2xXЦ=0�e ���y�527hx�F��"i����� ò�?dn�����[�7�j�+���/~�%>�0�\�8�j��38eͱC�.�p���~Y�c��{��\n�O���=#��I�a4N��߉Rۏ����/�����=>�%�3n�nj�5�{�����l��pi�ʔ��x����(���ξV������`�O��*qx������G$�(-@�3�G�;HK��B�i�{���r,PmX��IFw���S#�lʗX�E�z�>�{���S5,�����vt2c��=����{=)��e�7��{<Yu������ȠH�=��y��7Ӆ�x���t���{����(hC�k�֣��gg�Ŝ���e�{����9�!�����|sX�"�\#�ɦpQ��I'��Og��	�{��"��	�5kWG�|��߷�T��O�7�l�^W.Yn�T$�/��_�}��Hsvr/�;�w�w���)��j�.��\L��'Rzn̲>�⹾�k]Q�1��"ݾ�!�S�92}�n_<\
����xgMc�qݲ�z^�,�u�ҭ>�/�%b��B�ԁa[}��^HJ�"2��W��6f��wv�x��yɻ���A���y�����!����֍�q��@WH���Ik���Pλ�n�ܘU��GNH��p
����� �j�{�7��;�u�]���!��ž����t��x��o��*��g\����\Ί��̓f��!���QpT_��,��K.���^��MC�DC�����MR�<K��n�-v�(kUY�Q�%�LNuCj^f�ü�'�^��I�X���w��I���-8@9F�n��=aӈ�S걄 �Y
�� ���
��m���*��UC e`�,ƠB���!�8�zu��|�_/�������y���iY=�LeJ��:@�F (RT�"���pg�>������|��n���}��w|�r2u��5LDA/�*�d*
EF
*�e�,U5���A�d�}8�|>�/���{{g���g{(��5!K�/&������(����!29<�$��$9TY<��X���	j�%
��B���QaR,h(�
Jbl��(��2��ZȰeB*ŊAE]IX�X�T�9J����1�(����e��b�����D��5X�Z�c�Ad��(Ov�k�UR)vF�4�W��$��!��*V,�Dr�U�IZ���fڠ�2
�ak	R(�Qb�iD�,F,11"
��U���U[&3-�q*�)0AB,��{�Ta���E����~�6�w���] �Ϝ`�v!�U@pEQd�Ҩ�cv�y�{5�Q���HsZ��,y����{��!�9�R�z��r=���46��p�$���ߙ�0l��(f=���%����lI�ŹA-�6�6v�sw�U�n�nd	��  �r�jص���"��܍$(�L���Z��^62�l�gM���SJ2蚕6��xq��� Lj�K�84h�z��k�����\W7��=�+�(��\8"�ñ��cn��� ��3�j�zD�������Oq���?|�G��"����fϳ��8��^"\C��� ��W�1����Sg����^f�����z�����gՅ�S�H@�I�"�8C�2���d�A�p�:Z�n�먼��sO�Q�����ؤ�"�h�?y��^_e�ê#* 廓̅��#��I�)g��041��tWXi��av���K^��o����A.��{����T���p`�(�A� 0遭���.!ݗ5ہv��R��0R���6�H7��G��O}�m��Ҍ�p���qÚ4^�9{�C;k=�\�;�T�����	�Ғwt�Ү�
��3m3��pˮ�D�et�E�6��B��߼������r2�LER4h�����J�q��^u�1{�oM)Ӟ���$8(�h5I���hnP,nSS\��R֝�!�Y� �+8����;�:�ɨ��ppA��చAȪ�}��u/lia,�'�ӱR��I�j��N凇w���FoL߱HS�rՠ�g��eF���ؖ+ܦ��s���x,>��s��^�v6������\���^�:�p8��z	)�^����WE�k���F�&� ���ѣ�~��1�o�hyB��m�^��OQ�q���p�b�2\�9N�F����~u1(���)�]8W:�UM�`4f,����������@��:����ydC��y�foe���׳lJ������DZ��Z.n#���+�op?����� �0�|�Q)E�����z�|�ضgo�)s)s-m�*6&�P�#Mj8�h�gٹ��e�MFI�+rÛ*	���Rl�J�6	��WM5K1�J�9]���%�"l��.i���g�]i�jJ�6h6:��ۜ�M�8h��0F-�j,��츩�7f���#4 �S��j���"7*͈�b����0;Mf%6�biF!-=Ͼ��~5���ƶ�s��5fV�&W]1p6��&Уj��0�zZ��bpA�D[B�L�ݧ��ǋ͙�!�8Q�d��z�\^T�W�pj�v �;"��5H82�u-���%8}N���������v1��ع�a�=^8���,kSm&M�T�.
�$td�6�q:H.%&�r�"�2�q�AN.r��w���U�3�z��+*9�x8G�S��0N���;��뱣q����e_��b9�w�u�����'6���ksh����<|*3�bn7h8�C��zT.�v"�{���MT�0 ���U&�t��>���5��=;{׶�ع�i����;I�#u�Z�r7k_��v��OZj͝-ԃ�~��m����qv��ҍ�rҒ�3b�BS���8���}����]��85I��f濮2���������;��ݕ&��ہ���۳�2�@]�����,��4�g!��Ճ){I��޶��ov�OۏۋgT-�˟y����;�N�R&,K�y�&�_�C�eH`>A�d � �~ݝ\yA���O�;U�I����]���rA�Y:t�JÝ��u�Y�p�x��3 ��@{�ES�b�N��o
�;�z�\���M�vb�6�x�A2�gcv���^TR%8T��f������}��B�Ä�g �S�G�����A�a��\W��%Ϧ��_�n��fG��RUH�
��CX���c���#%����K��������K�$�=�8�,�>�#|���&�p"�����I�Wf�n+��mv��k��d��d�±q�+��X��]� W�1�����x�w�"�?p�8L�pk����E�S�H�6��z��&�v���fd���f"Ԙ64�,�Y�o����䍗��c�T��`S�?Mgtv���w�ٮ�U�u ��k�*b)��b��v!��1�x�L`�z$�us�&p;6�s�P�wf%��t�nl�:U�og8&ϋ�[�"��B씒�������$�1���Ʃcڭ�!��;��Q��o���Z�6���:��<�����^�R=Hj��K��[�����~���P��3��9ȵ��B܁� �  b���,0���~}���%Ѹ�s�D|�׽:X�x)�=�<�e����`г\�k���؊TC�7����p37y׋�-x���75���-�X1Fm;G�U&gj�h����~/.z��٬�4W/fF�k�J�ػA���F  �9N����>=b�g߿-r�6�㍺�㹹�9kD��e�����Jmf��f�5@��OG޲ߞN}�j�����N�^�L�vJ
�8Q�<��"8�jA�p����U8pES�� �c���1��z؝�L౪vv���ח����^.)�7��#5���.yU�����V�/j�� ����ᘖ5I�څ8��T���b�TS�?$��������~A�5hC;!UB�p��/Z�F`��3��j|������' ��@8��e��{�PW­s@5h9
�Ӿ��v�Yz��G���]{��
�3�y��p繛e��$L�C��v��E]L<�|���}on|���;��T��y�v%��amD��.��c�� ��0>�P!�ԄB�B�a�v&��}�h�\[� ;(�!�-T�؉�\���É^��1��gh��67^v8#3w�x���NFjg&�܂Ʃ_qG(�-��QH�I8��K9�Rw1 �e��Vb.m�R#+�j&�.J�G;O�����|���zb�"�Û����וv]�*�b��s��f���db"��gm�;E۳�9${�r	�N�O,��������49�9��cS�N�_Dd�_q�*��i�X�3��!CΩ�R�e�4S��B��PpE��vpI�v縥ڻx����Ȭ������m�ncx��5�;��R��g�6��0��#���irv� �U �ykʯF.�O�s{8k��Y)dE�
ƈ���CCc��&�� �T���D85J!�zx�x=X��v����{'�|<U�p�| j�vǖ @4\� ��p�uP�G:!y���͞���������{9aN{�L��|�3�KE�)oj'���'n秆�HY}�Qk���m���+����OS�T[�C�&����êS�7�4Y}�!������k�~3`Ű*����Ξ?��BO�����x2�$W:��=YK�T�9ؘ�l��t&n	v�y������ok�0�8���k���8�аLۙqD��ve���5ʎ��%�5�e��kb�.�rK���)GVif�������p:�YM��A�ٹ��ju#��M���D�յQ�,%Xٵ���sY63�Kp�kjj����H��\�jhMt�*v"�J��'����� ���[����h�0c�j���Ī�!6�2D������pX����ES�TC�������w�����\{�2�����ͫWA���}�w�ϥ(�S�0͔E;�CZ�#)8 ���r��FtrJ�ع����~L�v�؃U�Y��;���&e0v�^���]9�!�
�� ݫؚP�rB7�w�;=�g����3���pA9N����"�8j(N0�a �,�K�y�.��g��( �k�N�*���d��I�Wyۉ��'"(G-;pj96��Ac:����-~r`����}C��*i�>�1��^��ˈ�@�9b��zf]e�͎I\�7���~Mv��N�j�5:6�>��
�K	m����_M�qA2��.KTmy�l�e��͛)�G9`]����^�F�>�#)���,05J/.s�޿u�E�f�_^��"��L�n8pG�;�qlE܇.�n�$b�D�~��w�j�z�d'�����=B��C�`a�z��l���K�Ar�;�up*�&zK�WQީ�9�T�&��~�)�f�|��1f�1fb�07d������7�}~���t���i�.�P�T��$���z��	dʱ8��Q*���`Ak��U'"���.B&㧋�/��5ҹ�.����r.�Hs7hS�
�P|v���'�g9�Z �S8f�w-T��g;���_4\FkU���d�4G�	U?y��J�-���N��I�5N9��f��>)�^��rC�U��o�tGM�7x����_�A�@; I�L�E�U#�"�2d�������~����\��c�GMA�WsTM��55�������ŷ�9e�r&����8|ۓQz;}�UώsN�8��!c��t݈
�ҢT��Rg�˛9p��	A�\�n�87�+;)�=s��C�f���������)��[Zb�]�zB���A�"�����n��������a_�.�����A:rEgL���CϽ�b���֦�6�����N�r�FZs�{-:����=���k�&2Yd��h ��W�Ã �,�A,���,�^����:�Q�Ͼ=��۹$ v�85I̱��*�M�OZ�^]�0�M��I�|b�b*�|�q�{z]+���C���kk�kպ'��zQ����؊�g�1" ݻr)�Mn���8�����WB����w�����
��U�3����	bE8x�w�]�u��K����+û��D;"æ]��Չ� �W�����e�=����>����E[�T�f����ýV�n�WN/nt��]ٯ���������Tﻇ�O<��|��k�~���fP���j;gK�r=�w����Fc�"��e�~��|yۼ�Jn��٣/��$�~_bhy�L|�8:�������3�!Uɽ����b����r	�A�ͧ$��5N�� �6��z�Tƭ�T{L� �+\9nΘ�*�k+&w��ýv�n�s� ���~���TV����?L��J�s_eUX��~	 cl܉]#��й�V����?v�����8��~����q���g�>=o�/=�x����0��"���g���#�\��=�F/}��" �p���X��c��0e �̛Q�wz������ky�M�ÐEۇb*�=S�����Y-���w��G9�gy3k��V�Aѩ��ņ�F�b� �q���L(}����be3��L�� *��N����h��1Q|*�1F��&w2W��� �8psPpg��Y>95�a�1˸��l\�f�g,[1ݘ��7��ɞwN&�;uq��\�X�?����d�T�@��{�A�7n��T���y���)���J���yf������M�Í�A�p�U8pY�Rkiev�SJu�o�]cZ���^��O����7�b��U��<RXoD{|�;[.+5 ��+Ă��k�8 �8^�5T���mY��4����z��gG]��+��M�j��Es�T��-T�2�"��.������Q���Ep����Wx����y�t;���$���v��NL9�F�l����}Q����a �2{��*?{R�3���3�;�F����`h�������ݨ�os��kޣ��˛�o�y�� I�nIq�g<��N�*Zn��?wa�C�.�zs�3Ϳr~�a�Q�vK�y�e�ʱgd�)��p����\L�o��/^::y/n�JM�v��M�x��G�F�v����;P�4?�	�{w`�_�n�O>�1��엊�;���w>H��`�9����A{�Jm>�/�Ӭ3
8�ݦWS8�-�s�!��E�}��Q���]�@�*6n��̽;��v���c�L1��]}�7�X��2̤j��w|
��+���+�&Z�N�F�|��ɒ��zs=���Y<:/o�~�4!���zh:]��^�<�xJm4z�| �2�{�ۭwǹ�駻Xt#���]���f��������c����zt��Vo�gy��U��ɔ��/x���_{q�������ޗ��Gzn�{kc�bQ�Ǐs	���-wˏ�{�����H���|��ľ��	ug{�����q��9�xt�,��_g���<S���嬨V�3�ڡeh{��q�qL�]?:)	n�������2.
tc'�j�g���(_,x}���:2#.�/V�b����Ѣ��$8�(�gĀừ=,݈�ۣCk}�iᰤgƻ��ڱ�v��Ȗj�
]�÷c����T�tϥ�G\x1���F���$����%���ľO��L!�Y���ѩ<{����hm��_}��6�
�O^ɥ���P+8�E<1�xr�ₑ��x�3ȱ�C��6��@�$�!�)m��²k!��P�(������eH�3�'S��������}�n�=��{��2�����+�uEL���e�p�ƤĩH*����!e�;{|>�����=���>��)����2!2�xEe¢�Ab�l@����g����������=��=��{쒈��i��b������W-��HPR5HR�,��d4*�\HUb���)r���S�1�ܦ��2�VcU� rݴ{�]��-�Q�11T�,b�,�*°1�W,�q�PR,2����0(�/ ")��*�
z�T��P��T*jLI�Q��2�WC��Hj=R�-�d�q��* �
�(� �)���
�k$���(��VC��)̠���3�5(�<�&��[!��C�"��R������<O�L�Dc1D��2�4�� 0��U`�&�Oz�ÍZ 2�k	��3V+�ˣ�XD��5��#�Ѯ� b�`,.3f�.ȳ���]%�U"[0�Z� �4�8m��9�t�1�*Rm�`ж�0є�A����3�dl�J�h���tNK6 ҭ&8J�-�h$��쭆-uk)�*�ʸ�̝�٥6��n:��,���H��s�-5YR�KuZ(�l[]sq��E�f�f��D��h�Fc�\jC�uD V���e&�escsGuJ�#��v�X9��GPX�lV�k	�cm�+���f���,�ks-��� �bE)���GQ6����Yvf�X�]F���;&j�X�JӃB�6��Zlf���eNoE�]��a=���vK�8� �,4)b�+m�M cqZ�KP�ѣm�L��f.�Hi���hU� X��֖�]	�s�0X��Yf������#
6h���c�K�P�h͆�LdcXh%Cuv��u`�$��tU��\��3Mc�M��ం ۫f�;��A�Ķ�35�`𙒶�-%l39��ֶ���d��[Z�E�`F)ab�m��ءy�2��Ń``�k�6�7)J%	u���յݲ��`�K��(eز��䚵����75��&�b�ch�5��ݩ3����Z��-�a���l�t�6�d��NsRʏ,�!u��іl�׆1[��X��j�QL��tb�d�"β�amcc!���Gu��fM:�aJj-&�[�n�h�ihul!{��l�;u��PZRY��Q�J�[��XP+&m�H�6�X;Pjl��r;ٖԗb��Y��Jg\a\�!-v�F�:�c	�#əep�kp���e�aպ^����V�V�3��wiz�4.���u��d��H�ןYz�8�nͶ$J�e����kV�-� cl� ���K*,�Hi��9�k6�hZܐV	d4��%D�6M��r��K
@���]�Ykci�1͠4iL��2��0Z;�U[���1(.5B��R��m�f��p������ƌqi��3�{K6�����.�&!WK�CZ�,Q�S�����CJ�r��_�)�u-�CaZ�]VѸ5��%c�u��Vjetũ�̷dn��$���+Rb�ݠ����rmGg-�>���9�y����z�Eˇ%��L�O�D.ӐM�r)�0%#\ک6�!d�cI�V��כ��Q|*�p� ͸pj�X��C̃��c�F�`��C��d�0�������g�b��M\����7�����]��X�Z����7i�i��3��v��0wK��$c֠b�c�޹�����zҟg6�v����[�������>]�]8��A̰��ć�ڝ�e�
���.�r;3E��)כ��Qp86q���MF�1
��į�̈���AL�w������$P@�%ƚ�Ƅ�,��j�-�V�D��n��>_�{~L#e��2'}�D８F�Wt����7�8��d���{|R�G&v5��U'��.�ħ�8��>��OTs����wY���OK�9" ]U�{�Ѻ=!�w}�ѯ������M�x$f��?xy�1PG���-š�sdC�:̒�#2��|��ŁXd� 9��|~� ����t��=�bͯ{9��ڱ`A�p�ES��FC�U�n1d;;y�%̠��rS����X�K�S�����]��w6�bo �E��v����[mÃv��n�8�B�'�uO����u0���͝��o�v�L�����7P/;up6��s�={�\{ղo[A�' �z�s!V��.�v ݸpj��{V5�_����Bn�ovVF��Qf׽��hq�A�-��؊�v4���X�W#������n�K�$�l<M6�Ql;J�4�sS�dn� �4��]��{���,��=X�ꓐF2�P=R.s6_bm�EE�:C��~�x��~w����T�8�pERg`j�8 Ѣ�_���|1I��kM�������f�L𮩛�y۫���r��3IU�ȳ.�9��Gu6�X�1�@;]�Y��5N%���a��I3�����:g�\MW�MUWF��F�}̪7���^�@��&�x�'o�Z6�$��G,V��{��6��;�M�:�% ��9�,0C �~=�z�/���=�׽�o���+�cz�v��ݠ�RLC���m���G';�85���"�C	�9�+g�����D��g]��f���<��NAn��[S8�A8@���*�r&��n���xR�u�<+jf�^nj�C�5�85H	�S��Y�$��$�\9I�G9P��G2ڵn�Av�����)��Lܔ�s>���� �١s�#�MS��˕{�]��vc���s���*ve��{ F�v!d_&qJ�v�W���;���3y�Tq�����o칼�-�+����Y�LP2�;r�8"�ب����0�B�D��	�r/SU&j�{b�]���^؍����~�˹깝�3p/;5sL�r�ɪ�� ��H ;B��T��]�A�p��8� �3.U�����ُg6�8�JΗc,^�6����<;�U�W�����^��m��}�j��+��)���}J��~Vw��M�L�O���{=//DJ�Oף�[{�H�#�nC"q)J
���<��?�G�p;������T�OgJtW�W���k��d��|�.x7�1�C����	5H8"�����1{A���g��� �AA&�\Wꮌé�B&lk6 ���ҭA5��>߽�q���"�3��g�T�wL𮙛�y٫��~p������%��ь4
�D�[ݲ��d�qC�@Ozq�֯\�ء�$���oj^�eo{����Ͷ��^ �ES����.^����cz���lg�V�ԝ�-��U/1�T��;����y�l􊹯E���|/�z��g�~��_=�>F�C0�1Aqw�9K��k��ܔ8�2�8b.�U/Gz�kzxT�����@z�2/���L�F���A�8"�8-T��S��T�k|N����>���6��ۯރtg�ͷ�ౣ��1A^<Eyݨ�f}S�����G��U��^�Q;5���n�lU{Z��;WY��Q�6jn2���o�z��~}ؼ
�MjũùĦ�۷�6d�� �i@x�r�au6�2����ަ0�Ie����F	�J�a��mܽn�s6�f�3GMة*f��AՆÚ��6i�Z�\\))��͟���=4��sļ�X[�XͲ⨳6��usM{Q����L�T�����FṋIVX���b�b�:���,�������A,�̅�t��u`�X&����	ta���FRibi�m4�\V1�ת*&�8�S��؎�f���f��%��������hkR6���XM@�g�*%�J�S�-0h�x������O��qkHs��N2k�V�����E�r���\��>ϴ�Aۙn��<h� ��ES�j4`��k��L>�9��d��O-,�Y5�<*{�/g3�W1���+�sT���>�h�#99 ���\��,	1 �4��� ��̮�RK|��}3����ϯ���&mh@�[�D2c2��̨hB��r������5I�ϴ\V�fŸ�ۇ��&m<���.�
+��pFR���Bav���U�l���YU�:&{Ҧ�d��@].,[�T�$�>�ŋ0y����^"���t��֊f�wU�P� Y�+W�GT�ٜ0�+�s6�c��Or�/�e�O8v5JX�i�8��WQ٫�=��g4�:b�vߪI��H�p���؊�dƩx�Ʃ;j+��<4>���W�i�b�k��Í��[��3��j�6ޘ}܂���v��9�M&��p/ߚ~;����R�.��E/{��!�`>X�b��j��;���W��S���������a�8͠N���E�{�v�k�識3�8U�d��ݴ�v�q-�wũQ��5z���=�f]љ�6�����×�r���s~N T��y�^�Z��x�-��v�cLě-"����+�����O��w��E,gsX�k<X��{_!���8�H$>���SD[�yW�D�>��9d��0�4W�Oo���h���M�c׶0l�gn=�^��K�$m�JH��DQ�)�.-\�iI�U��6Q�hܩ��l�t���mf]�E,zb��.�,�9HҢ2z�w���p�����ĝ��]^9�\�]kf��|M�V_0�ﻆNL;{g���Uљ���1�t�g�p�ee+�^��b���;���8]��B�Ñw��s��*Hze���N6��<�OZ)N\`��xzk������o�m�����x��UF��%��<�1Fu��5@W�(� �~��2�w6J��.�������@�����)H�J�{=}:��}�~�q�g�,��0 ՠElvT|`�T��2P-�N��rtvY������L����o����tJ������L޳�x�zL�A�(z���8 ��8�B͑� ݸsF�-�#�I�B�Ê��z��r��*g9��8 ���S��ñNk-YOO�.f��A$)k�{�}%��*ٔ��M���KD2�L	T�ZRl�Ⱥ.D�������-�|�ld�z��MR��rc+=��G��E�����"�GV��}�6\b��=H$�4�A�E���NB|�^�Mf;$Q�������DLL��vj� M��,	*Q�G(!�����=������'e ��L�1h8U&�F�j�o����5�[1O^��T��s�o�p�g�9����mY��8,%��_���#�:Ӑ[ˈp{�kC+��]H�1����.F}��rݠ�\��{Z�Ϗ�w���˫�'�%"ʽN�����|D�Zs^���YHM�����b�2r�*��oT���B�!X�tש:�=C����C�ET����_ώ"{�������(0�e�w}��L�96���wu�}2�3��\  �V�1U�;b��1�G��r�b�}�x. �����փ�0�R�e"���e6��K��a���G�.�76`�:w��|�=~�#�ۀ�v�e�[ׯw�9������Y���9ƈv8'82z`;
��@eN�j���D�Fˑ��9���rc�=��\��E��@��daÃF�v�pv��!���p��țp�f��1B�ÀDR�"-Y��'}�\��>��۟?���y٫��X��Y�ohUI�A�1��r3�����|&`��|��z�gs�:^��m�pN.F�y=�����,G�pŵS�@���T��)9]���7�ig�g�X0����Fx�f�,z8��8a� r�r�ÃF��$��eZ�F���~��Eī�/b�ʎg��O} }8����K�}=�L�w������L���@���-��c���~$���`=�mL�R��6�����O	/t�4����]j��e7Z$M[�kI��P ���D�w�1rut�S3����Y�1�TȔ��5����)�B�7��.Ls��tHQ������f�P�0&ծ;U�c2ZW��P�R*����]R��LGI�<]V�9�V]U{J`Yd�P���KB���ډ�[2�t��jL��Z��ɝ���Fdmn�՘�
�2�,��߿k5I�-uK%�64�l�ײ9�2�R�f�t-�!��쟞���79aT���Ͼ�ffuw�L�^�;5p#4�{��S�5jl�dV��iƲi���=�0�(81H;Z���Z�x��笄�g;���8� ���9 ���������9�nc:�o˳�;i���v���ݕ����so�M���]��J}��7���v�9�AȪL�@qw��^|P���f���m&ӈsc k���[���g�g��'�%zd��vj�lQX��rp����=PrE�3�4�X�'*�A(�A�A��j���{t1/w��#1������z�J&s�m��� ��e�T�ŨS�M���)WU�ioߠ��)Hl�D�-t�W`M�B���4һf���J��%��E� ��g5I�T������l��2fx^&;s�7��
v]9����7�0���fN��̦������b=;J�����C�Yn�n��zY���.�,��C���n�=���?.�Dy�4�u����ey��bE���)��I�7��A �,Ɂ���+��ų��}��^{;�y�D��v������6ݜ�.�^�a�T%��9��V��A�N��T��,�8�:�ʃ��6���2�	�Ӛ�i����p��L��F,�` ��I�w��\�gF4b �'-T���.�{3��3��p�	�z����&y�����˖-Â�j��h�v �8Sz3Ra��c ���Ɏ�釯�����s�2V�W�&���w�mu�����w/ �_������e�70!���pJ��H�iWk�pe��dj����s�m�AN�,��;o�m�_weL'�����q�����}�ڋ��B����D<����P��`���^l���_��M"ڛm;Tغ��ݞ�lO���.�]!���͜|�Cn$��,w&k�,K�������v"� H���:ܑ�#��w5J����K�j�>#��Xs��ׇ#8|}��.��:��4��>=��w�U�����k"Bh=�"w4Y�N�}�7=�!c�gP�B��C��2��q��Q�y�/%ǉ�PC��/���<��I3���C-ٰ�i��*�yI���7�a��e�ɗ�����'��	�9��q��z�<�M���ܴugl6�p���+�N� ��K�;�����|�.��;��=�|�:��S?S|�q˃0�� U,=�g�`�2�<e������`�CI7����W<{�,��xN���L}/���ݦY�;�� {D�(]���< �G�{�z�SeD�X����������=6n�\��K����KLyPO!��k˷ˈeճ�{]�0
bo/N�W�	�<���ۓ~��['���.��v,����|.���C'��|/-���p/܄���j��:������2p�����o��?�C3's��oN)�n��yO{���$d�9��� Z�ћBw�X�}���ٻ5���+����d��Ѷ\2�f��Z�f<`�U@�Q"��e,�˨nw��!����sn�x�ǻüR�f�=�����݀AM�:�Ǘ���q��`x�_��ݞ��[�Ͻ9�ծ��k�T�I�]�Bocᵍ�:Rb��-�ػxK��+���K��s�a���i� ������QnI�����G��["���e��]k���=��i�p,@�Z%H�~�/D�5�[��<��+8	H��T�NL�ɮ�ih���Γ�^L	30�v��Y:��2�QV�DU�R�")U�2�̛=�NNNN?'���u��|��dMU�+>q����3뮊�z�QHU\�ǏOo�����}>_/c��3��g��)��$'9�h2y|^1kU���,E%I[9L�P���q����|>���>�F3��Ͼ(��>~ڢe�fe�0��fe�b�c�@ְ�+RbȪ(*�PD�(���i�'������0 򘂓JɌ֡�
V�cR(6�dm
�-��H���
������DL�Pė�VYX�-+"�k�E�ֱH��a�1ŌG9qXm�%q*)�E���VeR(�b�a��*(��:C�Jȵ���g7HT+%B��-k�Qc���0Pk@Qb�⏡?��%� :����鈡骼���oS>�#ݩ؋�-�����f�W9��r�S�> �S�l�
�����L�0�o�8,l�c���\�{����"�Á�������Xԧi@�!�R��y��0�c�/x��8������𳜴����Ú4\��3:� �i���PC߫�{/ꊥãt�a�,�e��UaVh�3�kmGT��dR���>>�^�{��e�1����-Yz��;�����WL���YSɸ��%N��N��Y�1��v!N�G���o�1��F˱m��wf¾���K��k�"����.�Aذ���?&|��y��^!�2�� ��g��h	Rg�J�)�^��	��z���g8 NZ�\8��T�Ĳ���y��y�FH� �F۸cJ�qs��]��x�1Uy�ܜ�kS�����z�����	,L��O��}q�9٧�|���l����;�o�6w*�������>�p�gY����B��������f���R5|f�s����F=����iD���-4�F��&}����c��Q߷o�+���Mk^s��-x�$��TE�/{oq��<�kԔ�����M��P�&���imфu�Zetp�]�kW*m_�|����c�UJ�Rz��V����bxY�C(�g���y;��%�#��#E؂S�U��F�i�����9�g	���`k�c�wx����^ow'-�l�A�Ů�ve����������:q-�q�� Š��!ɪp�/\�Iu�ܩ�#;՗�3O^��6g`L�.E��U&�Dy�ʩ@#=Y�o���Ekqq�-;|��\*�ݽ=���O8Z�#lNbt�Z����V I��؀�\8"�Â�,�U@�*�J��Dה�-"jo3�����f�-�����5I�LER�����WhU|�N����U�9��v�]�6�9�+��?{����<d�^�QP]�C�s6.$P����d�T�~fT�	��Lb,+1|DKe�"�&�`���Y�;�q���!8�);�g���Z�Ϊ\�`��q�1Lm6q��2��jI��@��գ���Ժ�.�-!
Жf�wer@Ҵ�ٔ�ЩA���R��3h(���V�6�j�5&Z��LYf[��̲�1M269L�)�����ڠun�J٬M�+f�F�(�A��م3L̆qW	s2�ҵql�TԢ���\��q,�{/���}�C�\k��?Pl��F2���2��iu���љ�;�H�j�'�|��y�A�my�.h8�Zřog�ާ�\ٜ)�fUbC���ꓧ�8"�݈5H;� �R�	�N�mR��	1[�W7�m����.�賜�9i��� ���6_"�B���R��:y�x�V�[B�%�S(b�ˍd�v,n��mY��=*
3:���ۇ[��n. ����<C�T�MRr(ӄ����aMČ�B"uÝ:\�d8q~��+;{"m�}5͙�lQ���밦l�'s��6�a��Wj ݐɞՐ�*�
�]tl2����[�w�����g㖀}�j4|AN/XO�gs�m �/[�����t��4�uѱD��d�y�*.n�iv��f�����S�<>D�����,B�d?���ݜat`S�����q
�<�<���9`mqm����M��uN � ��c��͹C��N��l@x�n�
_/M��O/)�����'�&G��ND�� ��3|��(�?^�?w�ܫ���_�l�3�bB���"�� |� � �f,8��t�Y�\8����g������6bo<A�p�����u~ҭnS�9r2�� �	�N�e�����+��ǟ4N?��lm���s��An ��"�1xTh��P��K�@����'�^*��Gj8pz���f��dF���a�����z0)���M�-ccJp���IUqcS��p��Y� �L`E��=ӯѐ���s�ذ�8o����s��#1N�����cjȚy�����]U4�ħ%9qX	�"�$^ �
��l�]�R�[u3�
4ڕ�2k�sb[�O���^�_�D�(��j�85I��p��v���/<و\L5�UY�P�DR�7�UH9I�霘:F��'^@�#iÂI�L=���ǜ�b5������r '9�y�<v5�{���	7{��"n�A�e�7n=y����?n;x>g�}�n)���׾3�Igt�)[�]�\��D�w�>7չڑ�D0{�{x�;���xk��� ��D'���b��[9���93�3>�p�j�S��[�!����pAX���x�2;��s ��~p� V' �T��\*�7�lu���s�b�`�����sF�9����؊�pA�D �8�"�s�:z��;y�R�==O���u���^nb�-v�[c,�S�pj�^-�˘}{^]�����o�$�����6x��j��Ô��h6��4�kyh�b���e�P�'�rܠ���F���T�㯔�{���ђ��,2�����+��:p[y�b/]�iQtH/n��:�F�2��Dmi�-���u8�W
����b&'�ొ`V/0;n4_}��%�+����g�(�q���x���ɲ��db��F�z��b� ���]�w��o/;1p-v��$y���1I�,j�p�N��X���b�DS� ��ݡ׃�w۾�O\K����|b�q�Vן��b>�M�����wr����|E�C钋������<�~�m��G����q��z}W{��yX=lۍ�Y������d6�I�������U&�T�Ꝝ�.��ﰿ�n�1����{x͎�bxn&㘃�[mÃT��T��N��X!R/L��\i.��hiS+un�4z�XU��ɭfڸk*�ae21��$��pv�A�)�
yÂ*�wb*��G��ۻ�~X�fg^� ��˞/q���TA��rM6�R�c!v�M��ޔP�lu�m����0<�=���ToU���de�փ�Z��&�k����Ȩ�kyvs� Cn��jhTPأT�r���^Ǟ�,׌��咧��qp ������.ER* R�*�H#4�f�N��e��Z�w$j�q�z�����e�g8K͈L��Kl��y_'ҝ�'i<2j�Iy7�
�DR��Tz3b��xp�V=]�>���G���pX�NA�p���v �!<lOE �n��9Q�+�͛EG!�}����M`���L������u�w��?-܂8�<��H��	۩�<x�{�}�l�!J��b��}�6����m��z��v -_u��.�k�$�Y����w�#ZF��s���֥�4Gn��]����H慬�i��\�4(��-3"�isl)�,D�m���ԖR���FP��m�k\ڌ��B0�`[n4���SV2ݢ��[��k56vea�4�h�����.��q��6RR�rLL%v�&\JM�c�mŮ�2�	�i�m
q*�̳SiZ;9���3J���qU�h�5����1�Qһ=�+�!EBmM%v�)u.2���u�WX�)D؆V�M��ϸ����~TGpn�;��V�+:;,���H����@E�������.�*�Si> Ѣ�=>?�5F���8.��ƕ:=�y���|G33�1��x��O�̢�D�G��Ll���Ä,�qb*���6l�"��=�(R��;{.�j3���a|�6�gծW�4�.Rv"j��V���&��v��T��U�n"����s�7Sp7�8 ���w��9�DyU��]�pMR��8�w)�9�v$,�ےkǗܿvǷ!,���\�r��s�cT�Ʃ�ڋ'�d�H$ �[�:r�܇'�)(j2�h�f�H\B���4�����u�?|�c�,�>���f�rM���Ω���z;����:BD=��BȋAȜ.�S���(�jK\�#��jB��>)-��A��[쮁]��{��wӐ���C���O�R
��1�Vmő]�j�79��S�K�v��!+>��[�4(���~p<��A���̉���V����~G�:7Scr5�45HLG�dGl* X7���靐�C�P9���A�c���[�>v��{��d{0���1p ���+���'5I�8�
��6�񃈧�g �!�"�ge��j����<o3jj:��=�e�RA�͉:�c��2��Ye(
+�E�!��]�`WG�<��s���wY���r>��y�� ����Uq]|�z��w}I�;����~�~J.��VR�-�.��.4�2���W��V�j�k�;xw?����Ȣ�����Ü�����ؽ��Wa�\evbo4o��3���Acy�rr5I�U;��@^���vĂ6S�kP��3��5[Q���/�E�r�p*�zr�.w�ޙ���3H=�<�� ���M�j��	۴[��u��ܙ���ɩ����M�DX���ëx�l��Nʹlsn{�v,���gwo�M�@���:��d��sIاuy���G�<4�!	cV���p*ׁH
�3��o�����:��Z����MR#�9�]��c.2�1q$�2���Xx!f�rw��NZ�õR-T�*���w�"F7C�����SQƺ���FRFRpA�p�ES����9�=�:$V')�NfA=f�ު��;�1V��`�W�:�����1.�"[��~b	18 ����5I؂R��f��d�n�q�h��^�>�S��^c�F:D�rS�L�T�8 ���w�b�t�#]���A��/w�[=�b�2{1sb�R�o ��K�V>��"�?�6�h�����T�Z�������sO�\Uy�t�M@��Ga�	I��\
�;j��������Ț�ӯ;��9�A��L�?�kJ]�t[�>���Vǀ8����v�ʦ��[n���4w�=�b��7�w_g�������8�Ґ}�VK��>��Anԫ�y�|�U�S�!�ӓ�Mx!����}p;�ϼ�7p�`�}W�p�EW�ڹ}��Kk�o������y������d���\-�ErRv)�5K�/V�_�xUD&"gw�9.29�a#�E[l�cF�Tk.eP��5�s=��;��Ϩ|z� r�8"�8 �]���Y=/G��������L<���1�Ѯ��
c��M �^8�T�9�N�1ʺ#ޕޅ����SJ� ��vQJ����ߑ�Iټ��9�9m�1��S��b��	xq�ḊLQi��6�6��41�B}��4�|�j]�|��=�˘|��\�fS��[�}܉�)ow�.��0/�`YUN�P���AȚT�!S�/݋$��o�q�f�Jń�v#û=U.�� �CX��A�2�@]�v��}w��M�^/=^��ནͻ���X��v�9I؂�N 0ށs���f��ٌÂa�#�uA�}�f��=�=-�Tk;=������k���s�dc}�1�C\���w��Iپ��ٛ��yL�0����w���O��c��kpN��.����g��{ ��'n+ر��vT�^��yz���'������(�:��+���U���P�3�ս��]�2|��ټ�Z��s��G�����0M���.��uzL�ӉS��¬��>#�h�斞Ǿ�s3���C���ܩzaQ���Ľ�w7#����S(�}�c��J���T��<A�U�_c���uƯ���M��zm]Ͻ�ݗN+5��!�v}+d1��ˋF�<�t�V[>cX�6��t�DQξC�jr^�{w���r��z���r�,����5tҘ��s�oyz{���s#/��*���'zI4���>�w��s�ߦ�e{�vMŏ;��wٻy5���K�z=���o�V�'�+��@�ynbUr2�*PAU�5�_n�����rݻ�s�3�"o�Ep�;�n�9��n���$#�h{���"C]�hy���r(8���^�Y�qד��{���WU���{pk�/N�c�"��:l��ĔȽ����t�K���~Wp��D�7�M�=�����c����ӍG��Y;V�>ճhH�4���7{<�w�����x�R\�&��q�g����˝��u��{�P<�¸/G���Q�c½�w-R׃�����������ˍ >X��O���Ō�Y����l����.���"@`1�J��B�"
�'otz/7��F%����$�Xr����}E[�;�y��R�X��O	�T��(%+�"��L�.�����:ۏ��>��˶���h㍵�❧Ʀ�� ��j`�V��к�\�u��7���SX�,���%T*����Րd�ǧ_O�����{|�:����g��� �!�tNq)J
z��g�UW�E"��+eY����������{�ٞ����w�$X(E=J�oX3PX5=f���S>{zzzzz{{}���g���>eBT��R����K!Qb��LB���Wr��
��-DB�����2�1�̺�e�`2,�kI.RB��2!�7i�1��C�L��Z����3�BL`��I�+FK��Y���&1mX^R1���J�Ϙc�d�
�-�2ʈQ��Y[լbB���0�R3���x�/�/�C�e��SDfh��l�U�0	�Yr-�%�qsV�P$\"�-����n�t6�Z�20�.h�3(n��;M2uI��v5��%,Zl�i�uMF��u��B2��7�����-u&�k]�	B�06e�"�fٹ��B��5����e��݂�#�Uim1�M��m�ؼ�+�5/[f��,Թ����Xb:f�;*:mM�E��]V��+�T+���uW�]Z����Zb���58ee%������BZ2��l�je�&�.�e	�ؖ+�z�)v���E���e��ԁh�E��X��,22��f�����D��,�ֽ���t39��0��ųe#@�Zę�	�;c��ڀV��u!$��[�rKfPͥ`�.e�u���6$ ��JV�U�ͫ����6ں!B+*D+Q���؂ibd�k*��ݫj��!�Ʈ�h";��b��se��c��(e����ɝa]��VA�Ѯ�5��;cMם��扖�k��:i� e�.��˝JlRd�12�F��0WH0].�Y��h��2M��FV��]q�-�e���3\ F�^lsb��l��T��b��4؄�[��	t��K�%�[Cm˳\d�J��`�dJʩ�����[W��v�/#	V�	ua�q�f-Ic�
S�	t�� �Z\�j9�ic+a�ft�[�ҽQ�m�l$�4�v�H�����b3G����Pka��&�1#��-���� �@��������&���l�e��6��&��ڕ��PX�&.&�K�M�h�W�Ci�'R�����ιؕ	�5�	��!�s�Q�m�l���޴î���E��,�6��qC]vs���f����:ݚ���@f,tfaT-��b�cZ�.�.v]�ɘA�#��C���T\��"�H�?���Nu��7n�h-v�F,�b������ڍ����T�nnDn�vie�4�������Z�mb���;!�e6���B�E����Q��4̨�X��b9Ԣ�X��lV�m�]�W�p�nZT�L9�m�S6a�.c�0ǩv�WE�c*�%�e��s�EA.Y.YCL���!����Ue5T��]4)��~��?q
��ZJ��K�e��;Fe�]�i��inI�4mfw�~������+�9��Ʃ���˫�Խ�&;1qG�T[�p}���4��=I��U'̅R�����'x��Wk�e㜀~�`�������\{�͓��H8 ָr*�N��G97kx{��Yn(-ڙ����Rs,Q�U{��[�pw�{�{�p���xn�bӈ9i����*�;T��l�ߣ����Bb�c�b"�=S���^�Gv�����bn>��r�vV.�{���`;I���B����A��Mv��<=u�\`4�eu�?�F�q����l�pL��ۇU&�Lw5���)ž�j�����W�k���`�P�i�TԘbiv�+fH-P&v����}�^�<��O7עw�ʪ^�]zú-����\E�e����C��	��p�3N?aH�2\���^twEY��V�:�to�=�J���՟#�z�o����]\	=���+��>X��o}�&-Vߠ��N�Ԓ����6��Cn8���gh�[VN�wE(�3ً�'Ҝ�ݎRy�ۼ��G��&>��z�9�A�H5R©���>!�E�u���w��z�2u�+�5�D�b*�?��k��e�3	�_*jU����N!�8$�=br�I�׸%=�����y��� �8�>O�j�{�m
�wpF�L��%�N���p�U>?������1���rݰzw�����@G��vsT���� .P:T�f�����
�X��t�l"�4.ԠD�B��o6�-Rk��s��������Fz���ƭ. 7hvR�B�쾙S:�hT�Ϩ��8�z��"�Â'�8N�ARCɻ8"礴�Ŝ�:�\�Jh=��zk��9��9�����Z�@V鋃T���e�1�b/ψ�H0�Ipuc��2����Ů��Qcj�v�y��Y�y�=d��A7b�S�12[��M�=&�S�@���۰0���&�����d�d7������_������/�b��d��g����&�^b'����x�K��!i��B� ��;VV�+�^��zTd�m����ɻ������q�V�v��5�r�vp�<NR��>3��Wp�,�fv�����q槅��et�v5H9��k��h����2�@��A�a���.�`�-mź�#`k.m*���↖�F����'�/�pAnW��aT��n�-���'s�e�x:��X7��	�vpj��I�,j�b��x>�ёބF��kPpA�p�]Z�o���2�ͷ��mb�p�ES�޾�����g�
� �Ƶ>�1���r	����]CPɊ�w���{��3</ScpW�9�9�AȪA�������o�<��:��wb.��O���^�=|#0{���le��c^_Ƕ]���WU��Ϙ-P�y&zl�����9���L��_�/r��\y���w��<��ޭt��s����_�����d��ۃ�GR��CƠ O5ˈ �v�͛%̜�5���Vn�B��ڲieF�F�\��O6� ��|l�N�pEW�!��@Y�;���/���C�/�����t�B��]W=�$h�C�)�����m.��4=>�~��;ާk	KsT��Ʃ>��w��;q�ϸ^�"+�#�P�A���(^��]В7Pp<�@ݑ�b=HxX��4���0�G�3��i�t���^�������9���E�n5�3�#%d1v.�1��f�4��Rکǰn'Gq����#�!߶�c������r�ub*�j��/ �RR�C�ٜ�`)��Vj�����,���v�.�}���s����A�A�����P�s�Wppv�pA�p�Ʌ��2
�Â"��ǹ�D;���LBݜ+�h޽�=���zS�����' �T�`n������8�5=L���p�	�ug�>�sZ��d��x#}���_'=kc�<�ό�����}Y��]\B���g�`?o���1�n,L�[Uhm��_$t��&ܬ�~ =	��^��w[6)�`v�\�	Z��ԕe0�Aв�2:�p�T��:0s���]��-��"�!��mnz�U7k��*Sm�.d�ޡ)=�X�J��u��p�àW(��b�Z����S�]x��B��Zk�]�Z<ڕ�y�LK�i1)6��6�T)�aV�m@��n
��f��]l,3k��l6���d��I]Tx����?Yw2�n] �q\��Y6��E����$t�c-1J������!�A�-����@9j�7,�FlB}땏�#k�|c�=��$���A���G��n��Ұ`��S����ߥ��5$�m���NA`v�����9���9�p�\ �^8� �ǆ A�@�e�'u��j9>�Jup̍�鈝��8�w��v�����K�$�=+�G]�{���\[Ҝ[����L�8D��$����<�����*c�A�8;�9����vY���P��.����8&��!�-��:����%�5�1r��b���p ���X�CĲb��*�I;5#�O94]��[��3�w�j�v �v4h�h���U^��$I!{<�F^�X�Z^���)5B<���1,���n�q[Y���t�����ׯ EDzEv�,p���ÑT���*TC��v��w_�>����~7�78U�Z�ɹ�aR��p��q�.0�,c{�ó����F�.J�T�:1+�Y�3�p������0��1����i;%�'_y�Z]D�ཽ�4i�c�=y��g[�ϟ>��؄|�<X|���&~�;.U��_��_��x��{b����@�p�EV��0��ik��<��q��1�P6����#T����k�|����j��)��:G��!����ٲ�n�C7NwzOknzռCO?#���D=]�^������upe8!�d�g�1CJ� ��t�_���d=i�К��� `"1õ���qK����,+9�j�rN8r*�U&����_H��n!���/�\V/�A��1���uIt�F�f5�9�D��5X�1Tq���� ��Na�Zhc^N,j�����[x��9�ϸ^�#}�hx<Bڅ�c�c���Eۇ,.��T����9��� �Mv�@��uk�#z�\b�n��fS�F㳚�}9��^�[9�\�&�^ڀqT�T��T����C�o��9�^Q@���N�:w.���{*�����t�k�^T�����.�x�7V%]M{'ެ"����kǍ��[��n�Ŷ%�~���Y�v�@8��Eۇcv�H*�u$7ghG��t��j�x�O�v]��gZ����/W!��A�,8I��o��k�!"����\�8 ݠ]��"�ԻH|;LG�y�{E�/h��h���bX����;&q��j&�-�,̇x�4�A��4�'$��)�ٙb2�,!H9��9�0�WZX�ܚ8ư3p�þ���`�P|���A��4���{{�=�І������9�(K@�8v"�ݍS��+�A7iŲ0w���L��Y��N'ғ8����_R�r��agKjU�`F�Am�	�(�Sc��X�QWD�2j��U�inj��w51�f�ĿN7��D 5���-�z���ѷ ����N�L�j�xb�g��[������J�z���F8pF�j8|�UO^j�i"LP��T\�ݥ=��������ǪL�Kn��j�6�/E��B��@U[8Նh����s���v�u�wG���M���#����vŵ�(�E���%נ{ff�n�'�&�ƶ��(ƿl������Y<�� }�~�� p��B��Jč<�)80�WBaU�*�Rwqw���}�.Id��z�6���Uo�o�S��gs�⻷j��1]G$��k�MH�t�	c�r�6���iK˔eR]h���k��j��C�?~~��ֵۋ�v��uj7�Om���5*�zL�<$�|�M���Y�R�����yף�<fkF����cB�����+��8���#�a@f;�V;�-��&P�,*��)8�z5���l[��=��)��(	�L��X�혛14�>ֳ�R��,{�����c�Iȱ�Z��5̸��̉����:,�����]rb��`[�P��9|���1��T�VFMw�_vG`�;����;��s�>;��Ǘ�'�;@�ze¡�g�f+�/Q�b=���uS��~�֥:i�͛�ί^��>_�7V�U��љ�=I��ˇ5-۩��`���pA�'~N��{�iO���֑L��Ħ׎��9	Rir3�@����+��5�l�]�TԨ�eKcMvu����sP!��61ڙm�Z#���a^����,�`
M�8v�E�@ѹ����,�n7eTn3JȩM1u�[YI�	Z鞱t]�ZB�.�Z�����WY��\ŭ�cN�)����W�Z�.�u�����ë�f��s�?~ŉ�3k4��p����\�M�Rien6���9�O����C�H�{����o]_O3��Ֆ<w}^��}�r�
�2�L�:�\5ޫut�U��OeK�>+��b*�{@L���A��=͹�/S��0�g�Ϝ��ؤy[�0>F�>{��\7i�)�{ēT�v��ʗ�al�y��WzR�.^n�_�����(\#yܶ0w��>��I�KL�3(�*}�*�"&�dd88F���rgr�?>+���L���+����w�zl79�; Ҥձ�X�� �.,հ�*+]sq��v7k �
n��M��˳���vaV�������%�HJ6T��/b�)4ˈ#�øGd�����=�X�MS��6��T���d���o�_5�N�����>�/;GI���7���������'hM�H#�C C"�K/svj�[3N^~����%/3���0�M3}��{���H-�A��H
�g�MU��r�<B�P�\N����>�[��s;M@,Z17�4��1�W���Ġ?.�j�E�S�5���Dg{/�����Ң�K�^*�n!�Y;L�cW�;�<�Sn��5v��v����r�{{q�u/3��.P�Z��T��_o�o�Az}�g��ڍ���'��v���A3�����2�1��.�e�FW��'I%�
��ooy����-�U/52 ��9Xk*����r�E[��W�iۡ	��5$�FY�4��سf�,�����|=����=gF_�A1�������Z䳂�NW��V��VD_������j�c�ozjC}{#�ɑc���O[�L"x��SWęP��˷'a۞���g�yVk����`��;��ڔ��o1�,♾~�i>�i�&-�q1힙�2��f�i��-~x�a6�x�F���D��7<p�}�u�y�T����d�/q�w\��#7s����w�΋4<��{�gk�;s^�
�8�0k�T+0s�rv�h��޾�F=죵"i�{}l^.��H��`�^��
�r�b�V&{�7�ߓÖ�xt�c��!�K��;ν�_i�zS�X�ݷ�v<�y�%g�m�w���7�:y��Z2�}��?L-��^=�a���ᗖ�9�0,�,�w/��X}����%�TӾ��~��y��p�
s�ӕ�OL��#�!��]�ӾY}�^���E���S!�'�$�Iս������CO_����(��zw��w7��E0?�0�(���r����C�c��z�x��9�1��_S��j.䛹���˗�C��X^�k��Ϧ>��\��Nt��o�}o)�s����=�x�#W�w��O�h���4ϱ�҈��V0B��oۜ�3u�e#|��a����2�KY{}s�w�\]�Yׄ\�6|�=u"��N�؟o��-��ʯ�� �n6�����AW�m��;����ޞ�F	���y�{���otxе�wU^Ó^�`��=�-D%�N�fM{Kݬ��Xv!�2jv�وcĜ`k���Nm��AGl�N<u�]d�F�e��O.�׌��J�Y�y��)�Y�t�0���C3��S2���_3'B�)j�q��R-`]̂���<Hn-:�㏗��������tu�38�=������ֲ�QT�IY�4qi���㏗�������_c��4���| 6�AJ�>C-"�m��D�e�
���\,Y"FdǷ���������������|J���S����)Kq(�d��]��Um�V,Y�N2�n�0h��-�j��$�i1�+E�*TU�fmn4�+m-�-�R�PX�r�Qs,�[H_�TD5�WUR9E�7-��k
�[(�X,ԻB�Y�c-V�Q�D�:B�Q�PU1�;�b
�ƨřj�T��N����"���K�"����\�-��Q`�j��*VAkD*^^:��˴�32cYKU[eT�(��n�7�ʪ��U�(9Kl�v�!�$�7��0A�bC��/}�}���^g���)��L�2�5
qMT���s�Fe�B�M2�D��9[O�Q�r�M(���qOI=?���s?Z�9���|�I�o�>Ԩ��i��#���'��w9e�kae6�����c`�r)2HU���)ij���q6
�TRa�����Vf�B9�[k�O�����:��;�N_�s[��;��gDT��z=�b�5��4Ϙ� ����gVh�E��y�o�d�n	��z�q��_y��M؅V6�7�z��+a���n^�\�L�W��j�H�~�P�C�����{j0�*��)U-���K���*����a2�f������w������lF�{�껟�^���~�#/�O.f���7̮�v�
mN��SX���}ܧ�����1�͟�O3����f��zQ� ק������x��U��&��I?�D��hb�	`j���1k�k���!3>V��=R����yꋵ�9\�5�S ��
��.�vZT�h���T�w:_�X���3lB�r�l���tb�k[	�Y�7�w��#��*e3����9y���q���u����h�d� �a^M�H%��P눤!|��3!��ۙ�˽�;����ꐪ:)�q�A�1�L��-"e	��0����X�u���Iǝ��[�͗�6�%	�f_��ߗ�p�˧���{�L����|��f3���SP)n
���%7��fC�a�PК���g���Ӎ�s1����z����V�.�Rj�od=lG��ފz15�7�+���C�H;�$d�ʗ�_�<�t�3��A��['*ʾ0.ђ�=}�]����x�߆OCouy�����в�la3m6�������h\O5{� rT����7Ǜ%�?�v�0�O��W&l��J���[��8��5�'k(��f�3-2;�.�R�SZ���7Z�QX��	X1r��IQ֐5�ږ;T�-F�J�)f%��\��И(���L�5\ޫ6�����)
M5ZP��a�����%%(1ih;S.oy72gV����d�nChV��IQ�J�*ۥ8�l�X�YҞ,�~����O�3,�W80�3K����2\]r�@�E�A����U?��S���3�}]��u��inzb�+rjFrjd۰R(L��8����l�v���Ы�O��鈈���9|��42h�E��sF�^'=��ɫr[��]�8���J��ގ���#P���/ٹ�!ަs����e4��SRv��7�ʺ��7�O3�+gaT��b��+�=r9͵szy�=E*y�X��r�i��BoJa2=ֺ�^<����_՛�s/�r��Ԁ�@L�^���y��\���@�HT��6���c��#���.���c��֥��Վ ��Y��7�=�v��&{f�ǽ�}Ⱥ����16��5�}"�l�Uy���/�n��'7�='���T/��N�c�Bm�
a�ۭ���^�j��;�j](c}OD�3��,���>Z���~�	��q��&���d���>b"Vʖy����p�l���<߯ec��܎s~L�֮ǆ��z�;x�iڥzfe���jp���'k��蹗� ftJv>�&%�4�Ui^��"�P(�H 3j�(
ܫ���ļ]N�����N�w���k�2��d&P���NUG��:��r�=�<����iN�֚b@�~�仙���]4v;C�IEy5F���^��l\	�� 9Sf[�$[��m6��O~��|��������oz�~��;�!�l�ؒ8@�{�-��p��R�\v�k�r!{D�b+�O�O����=�+�HLoY�y���3��m�	�U,��i����~^���^g,��9OIS�8�;�<���7PaFvo �k���>8������Ȉ��t=B�t0 �^�VQ[^��o�ޞ{S(y��3c[�/h��jg�gc���i�J���н�������z���FP�c�h�-6�ۂƩT�f1�ZQ�F7d
܌|�vQ��"�{����N}i�~�8v�P =�(C�om�e��7=\�SpA�mb#�j��H�J��￞�kF��Er�L*�>�������=��3*EX���h��S�������[��ɮ��,�;�)��_x�sE =H[���-�7����b�U����U�����%%>��}��e�É��]�X�.@� L�i�n�������q2��e�SqxqG]z�xߣ���LI��3b����o���g���^�8�~.z���2�{Xt���^_>"���Y ��q��E����L:}�����,�1j�d�OR��W���?\o��Zyx��u>^���V�0�4��f^aV�k&c��B@Ç�*�Zº�`]Vm�	D��t�F���+E�3a�9��݅Ǟ����fe^LP�ɺ:y>LW3��l^����L���rӅ�ז��{[IQ� �v�[�=���Ӊ���{���=)�ZM3+�*�ӵަ� ����5S�UC��zE�`=���s�3������Lǘ)	��Y�|�����@�6�i���B'n����1]�׉�,��ry����A�*��B��|G��f���]	y�������g�z@�sjeL���>=�[N�D8�g=����=W���z�����S%��[��C@��1�~ݪg�����eyYOP�5��Q1��K�Ht&p��Q|pmxa,�WEk�s���__���+���tm�H�,j)�K�ҡ��p*�AXЁn�a���5���3�[
�@&ۍ7]7G�n�X&-�Uٶ;Y�D��a2]����J鋽,eY^��\�^�ja��KURRm�*���� 	c�]ue&Ҙ͖
@]��AMcn�5�jA�eu4.�Y�\���r)��z��S��?B�lG�Ʊ�4rj�V1�a��f]�s�u�ó�	�T�	��Bp�>e�L���ż�����f�j�U!,@�3���!����q�M��b6��R��U�ޛ��2�V��픭⽷ژ��XŪ�-x�ѹnN�L;��9�T��M�CL�;S(	�2�6�9��f��=�<�D�����%�L����,F�k��՝N�EQ��ҙ�A&�[½�<� 'D��%uM����2��2��Q�U��ax���	������}�_��s)��>�~��B4GL	)�7(�G�5����m��%�BB�@+��܃��q.�&~3��]�4�zM�@ˍ���G��m���(j��E�z��=&%��`u�}S^4�"�w+k-d`Л"����^�}B����~N��Fc#<��S����9��m.�'�����E�L�����m���oU�����r��l���I�W�4�[Ҥwx��E�����GMO����{�Be	�A4���1��4��=�vFj�A�W�3]nߩ�������Z������-�
z�T����Ұ���9Й7O�(��9:9�ݸ6�=HL��A�}�#_<�l��<��!�ѹ�D�Ma�u��J��L�Rm�IJ���-K�VkҶ;ʩ5R��:�].Q9������a0��i��^b����r&7m�Tݠ=��W�����R��Uֻ=:���u}k�����n�bۮ�HL�b�A<�_�>��I����������U�%�2k-�xL^���d�5�r�M;�x���L�&��9�١b�f������νηUee���0�����z�r��7�|!�j^�gI������{������P��8�}���f���Y�Lobr�u��y���1oK�Z@��C�Z8�L+���Pf�!{*�p���^{�*�rC i�2��|V��H���� K�Qݰ;*�ƫ]��Kv�	WC(��5���~����(y��<w^��[uO�;{�^�L�=��x�����]^��������i�Sf8~����v��k��q5�3�u�Wy��y�� �p�t2HT*bk�UL��uT�{˯=�I�
���L71�Cͭw.�ؕ�YS	�7]�|.��*��O�����Cb�3|*���6�Fc���J��ꬬ�ȥ�{fI�o����j�^K�K2��YwL�&W\g�c�YUA�}k+��I�m 1��扖s�Z��U ������>[>j��o�3�ʘ{���>x�5�ӈ
���&�������ϗ�q�U��$�����}��ѹNٹ��	f�v��D.&"lMl���U���� �Y{&a�*=j�Tdf�\�Y^�X�TMw���C��K9��T�T�����r�	�R��O�d�
�jaڇ`�z�E_M)��Z�gT�}M5a�u�Xa�ЙS(L�3g��7׃*���b�yF��ΜSje2�֪p�^�M��wKh�Cԙ1�����<�ͻ�Zɸ���X�V&��$�N5߅�jg/=n+��VkkB���1n�w�R�n/xidê�v��p&� ��5���uy��fl������l�@�n��v<_�Js���}��!�\����-�|��U���i7���ս�ٕ����<�
���YNNY����W�ˌK:�o��ǄG��/��ys^z�'R��~�Z���>��u�[�\�ryf���1�c�]���zyeGc>}���oGh����z����D��᝽���=�ee\>�lW�.��?r�]�K��}�$;lԖ�l�}�:ц A��.��ln�<şn�S/�(}�so�nv��<��.vQ�y�=���q?���AF�B�^�5���2���S�W\]}�Pܽ��Jxm��ye����s���rt��P�f�g'�t>8���N��Z�}Oڭ�w��d�i��<�@�u%ۙR��/�z���O������y�\��ްY�vŃ�����D���/Oq>�T���$�6�/o�nR�b��{�X �vg�����L�
G��+��-Q>�/�.5e���V�z���;9ȄrƷ��9�-��O�ȼ����O7^�;f�V���Ԋ��W=����tG؈2W@	}[�������ܛ��U�Y�S��Wg��@Ӵ=�u{|��-�n(��6uYٍ�>aā�Q��./}K����q������N3<�p��!�ryq��{�� ��>ռO�]���n���x�1-v�o۾��<{eק��2n�y�O{q���A�&�V=�d{�G�Ǳ��j� -��(�/�>;��3p�\E�8��\����x�<�� �����{�1�x���I��O�f�f������1�w��e5k��O�_ �x�v��m��X��u�b��q�y+CS�e9��,���������oY�������F��/�]�a��7��c���x�k{J�H�˃6��$��-��)��4#�P�R��rx�����������?'�gC�}��1%h�s,k(��"���Z�`���ƍ�2͛>�6lٳ���3��c2}���Z5��2�lU�1�TS�1R,��� �Uk*1��&ϧ&�===��l������zv��KDD�ڦ8ɊԨ,P��U51��j��ł�%J-B�AEW1���V(��A�":�m��PH+mb�(�;Lf[e�ژ�e))>�W-QR�gzX�Η
-�r��Q�75Ub0Fڕ7	�*:�E��������ˌX*��)�3��D�"�֫+L��
RƷy��V���*1��QԢ"*�.[Z(�bň��R�YmX�յ��oṮX����F"* ""1�E�(�i�`#Z����Y���=m����c'�������V�dt��ڧZ`�����$�:$�,���V��3Am��0ؐjF-�2�]�%Ԯ��ڢsk+�l�*���P�6�`�r�Sa��6�ҥ��(�ˎ�k1�^l.�� ��rbKH��]�*CYc��k���\�iCV`{`�a�RͨE�E����`Jp�lM5tBڕ��a]�f��+U�Fb��ixM00��$3�d)�[�A#.�&m`HP�ל�[V]Hl��ٷ!@��Ii��e]���׵���V�@��lieQɴh�]B��魖�B�5p����3m�vi��г���bz����t�nb�"�fօ{l���HUt9�H�X��-���Z��x,NΩ�M��IJ5��VD+kbn�@�STz�UԸ�hFh͌e�SL��(�ɂޮ#WYX��Yc��X��)�%ibT�D��{�U����:Yn�#�[�e�CfT^�%�.�p��D�IM54pC�V�LV]��ҀL���b��5���8f�X�i�{yKn��
�������A�j5�ћ8E��K1)j�q/\�5�2���8��K�]F�9����F�=�jD),�6�f��+���ֵ�9r".����a�
�RZi ���(;P��#��ָ�KQVى�Iq],�kh����b0]L�����KU�]���L�4)ps6,4�3���\�,8��S2�öy����"@t��,����4(�5�A��[��`kR�9-�`���Glb�iv����ML6����"�b*��m+��T��c����f�v��K�%�VXڼ$�1�f�tJWZ��-��e���n�LWeA*��4���&@�^��ѹ�b�m�c:5�m�C�����d�����c���vkZk��B7��M��"�j���$B{_��[���̚����]Z��F�Ѝ7$;`^s5�*$���@j�9��K��I�Yqe�T*A�HՅ
↠
c#y��e�v�6stq[�J�ii6����(2�m�L�K��szɐ6���&X�i�ٰ�V<� ���lEf�\���,0E�����д]��Key#Z],m h�L�D��f�%S[���K�_��B�Ю���f[
]W+�Uh�����Y�WL��73�����=�������2�.i��=���>�U#��{�V���=bkw$�ɮ�k�i3���Y���3�L��'�ht�ɭ췚>��c��8��^!?��>�sv�M<�U!�A�GH���r���9VQŏ��:�:50�!2�γ���]�w�|m�?t�C�M�"*檡���ҋ�U�Ɉ�M}�������	��i0��2�����-p7w�h`��V�*�^���ñL�2-S�Q=�o�hx#Q��	r]k�ܵ��U�3�nlѦm�#�(*"�*��4jm��306G-�-o�G��v�JĻײ�؛-��R��j��x�\&F��>�O9�Mz�p�*5uC����V�8�����O[ �/���k�F��)�{�#�̼bx!'q�7W-�xۻ�|�y�v��Q��e�jg�h+"B�)�fK]��SL/z�o��yGG��o1�B�����hL�=1j��X���ή�ޞ�T����/����os�����w^�������5�6�S��p.��V�t��}>ơ�+n�����X��'�6�i�&T�W~�v�� Q(=H�w��Ð65u)��WL:���,�(�+i5y6=����~���O�S*ez*���7��"EN^���r0ڑړe��ƚ�j�)g��QW�n��ʲ�k����q����	���X�0�����Z��*�-37��k���~"6�?���N�����t�=�.�4w{;o��|�������>C�Ny}$��Z�
t��l�އz/;��&79��M2�v�q>q�DIw7Y�Ƭ�f��>��xF��a�����s8L�s.E���=��A���9d�	� �S.6���6���"�P�Y^˰o!����_7�zP�o`٪1��<�(�b��+�����sv\�)v����.m#�GZ�B8�t�0���Y�P��d&m�U&�ʸw�
��˟˳�����/]>m�g�B�k�	�R�M�f?���[L᱂7�/V(9z����3�	�Z�5ҳ�;�;Y�%�B��]xU!2�L��.)v?��W�z�E�w��b=�x
M�<�*�a���/z�*�,��>q��F�M�.^]�b;_������mǽ��(T����m�;�T���r�����V��7��*�]#fj���eU��F�R�;5yYC\\"a�!3�*3�6Ŝ��7Y�j��7�g��U[j�����޾|P=9z���W/Jf�xXx������/_�2F#2gFڶ읍�b�Bˬ5�⮪K�S��Y��IQ�Us �v�[��ɬ���os��9#�2}93���%1�w�$���%���Fn�
���-�˚0�&i�r��X����KbsV��uk�K0�^p;P|�T��JcsrFFϞ�m�x������ӗ�K�L����5�S�^�#�Ώx��C1c�o��{��}�/w�2�yw��d�1��^3��P�p�Jص٪�e��r2cS��e�t�Ax��E��o��*fm��{=��!K�c����7V{45�ڥ~�s���Y�lzc��|�th�޾���a�l�C����#��|�o��v�n����6:�U�"-U���F�3N-�	&
s6�;�gSHgM�]en��jn�]�TEɵ�f8�u�1�l4�/fGlLaK�6�,٨�����J���l��� ��ܐ3j�(�VkL�x��^�l\ҶjQ�K�3)��W�r�])�Mp�)Fͭ���VZ�F�c��<M���e�"�)�lJ�%�d��3Z���s5�]�=����d7Q��і���sr1�Wb14�求ϥ��i���b���j�WQM^���%�,���Z�1s�������x$���=T�T!���P=9{���S�ϧi��ʆp&^a��Z�u�jҌRD;F��t�^�ykG{:��{txT̳���*M����Զӱm�&�a3�:^�;}�`�n�Gx��f�Q]�������aP�X�S�=�n~q�Z<�b�"���C���_{N^ԩkɜ̺>��޿[;]y�U&z@L���/u���ʾ�+U]��Kd�W������M/�^-�>[���!����{K)tb.vv ���\3[�#*���#mx"V4�+&r���'�i̷��j0C��Gw�����qX-C��K�\L�j�HV��
�S�� GT<^Āi=��W	��������o�g	�j���Gh�O9yrΎ��/���e��;������V�Lܽ��e{��h � �4K�
�Ҩk������v��tR���A��$պ"SW/Ji�&T�A�4��Rw+�{if���U��55����z�&�i��Ӟ�K���A���LS8��7E�{;�Et�C�葴��]�R����9�Y6�U2[�%�~�����o_I���)���A�e����Z�d�D�Q!*꒭"��	(.J�d��;3KX�l�UH�IY�E����UxWph�;�i���P�����5w��xʟ~���C��P�Y�U��N
�*�@�i���z�G#Ss�䢻�V!�v����y֌0�W)� Bd� �UVVt�kẖ��ᖮ���|��*-��ay��\l��;�V]� 	̧gIŝw�!��|���1N�z"���k0�(]�[[�K zH��2��bj��HL�����3<_G[vUPxT�����^����j��^��Ɔ����ej���z�����+�tv-����J:��r��S��'q����tۖ�kF�|�P��S���743�A�1l��M��ZP�;�r� ��:m)�o4�>�#�{]ov�,��q���s�K��&۪����g��TxZ��z��{���
�eֿc�w��np�BXWwyY=۞�h�v->��ST��Q
�$��si���{��ģ�l�Q]­R��BeL�\����G8�� Zg�U�[ݹK L�fw5y��}w��
g���@�W��Q^;��hn{݋�kԽ6z��΋��{�����q�"%�����x�r�f�*�ѐS�Ř2m��t"��PO3)$j��)a ���L*Й��y9����,�1AX�����Wz������33̛���*|a�UB�'N���7s���v�t9r�-����uV�#qa�c��3p��k)����*e	�5���q�aE�u���q��˚�c0��nj�X�#笉8����Rn��9��o��$L�p�M֋Lڕ�}�����6ô�k�!T�e0>G<3�3d��`z�:62+�Wy�i��=R �T�R	>���ku��u	�{�4�Ǫ�GA�ެ�x��|"��c�N�<�+ʫY��	��wj�b&奱М�Vw^_��(L�k�.�hzV@ �� 2�u�Ǐ�!G�⠽8��nk%�n���b5z���Ҡ���P�tG�*����F��v�ΔK�B��6p��B}:��8x��,TX��� �Y��-�
�D��<B3ڗz����$1���eel�J�
��]q���f�1�f�<ЫLkluFk�b/3U&t΂�l�I�n��ݣc�Zv��&e�+�iTʴn��h̲��:�CMM)n��t�4L#�: .���������:��]P��Xe�1����ȲZf�ত%�
��C[�Ά��s>~���Dh;Z�֫/.Fk�=H��Qqs*k('&�D}>��o�$���s@T��n�3������Wy�Fx��?�>^v�B�
j�����X�2���
ŭ�6mF�{ז��7oh�uJ��Eck�L7��='�~jd�wn�:�ж:�EX�5����,T�kzP��ڪ��4B�$��x���q�58�ދ~��y��9�>~�x[�D+k�hk�lk�v���m3�����S������K�Iױ��*�L�3�]?��i*Od\�*6�X�w�O�64b�h���V5,����P��Kk�]�+��L+�e�8�3Y��Bb��mD�ϛ5y��U"�N�jgܮa�c@���sK?gz/������C�9����չ7��J���`S�F!��q�Ꝭ��F��'�0����:�vyX���^]�o�w�U�n����L����*eL�U/�JC�z)���,���v��1���Щ^��303��5F�����<��	�*
�Y|��2�Ff�	!�SX�qȷ�wY�)�A����jdq�9[t������	˫x������M�vy��7�sfe>lO��*@#=Os��a
볪�S���P��e�.l��\.�*���)ء
ӏl�(7Z)���2io�����otP8���z7���8vv2�2�쾌��Dm�:W���@�
�U�٘*38zWd̹qv-�aA�aO� ^�2��M2��X���*=�z(��Ȟo.#��r9T�2�Z�+u���3�,'Np�ʻ�]ػγ�m,�{�"��]����9肧�m؈�|5�ሰ�{���5cz9{���V��w�#P:�}�+�\��ftm(�z���]�Vk�3`������8�~�8$tiv#�x�{�s���t�f=�vm�0�;��yE��tW4�9��M�ͽ�������n�� xN�cO��𨾡����ٯ"f3s��wi�?{��,=�O3�(��=�}�g'���پ���'�¢m{�ݽ{!׸wI0�����}����n���J^2Nc�.��W�gW�����Yѱ�{�=�n]pt[��z��g{Ϡ�H��
�o��Rpj�2����<��K�H����<^PNW�_w����I��N����®�s���<�ï����� $���N�;wt�a�x��`z�a�*áy�!e�G�i`Y���ʣq��p�ђ{��=��&g�03�q&�E�`���H )d�O��5�z	0�=��,05=;Ycj��������ד���T/(�.�:����Wt%���<1���<6wa�d�=ק�r���t�x�#�cSy����%�a�;���J/��Y`�F���H�᚟U۳׻�f�Ip��w�yH]���+w|�����Hd��7r

U���xp�0�T���B��֟X�ٓ���raA1%��)�#�&�8��+���3�:�Ѿ�����;G����U�1�/S7&A�lEb�Eb�x���T���)ƪQQ��8�|�����o�~M���gѭjV?Z���X"��
�AH�"��n������fϧS�f͛:�Fy,��L�|}|��X��e�%b(���mAb�h������Kh��(��\��2͟N�&�===����w�H�
*�|�
|�
������b
�8�Z,TS\q`��	kw!�fG���<��W�J��"�0DE�<B�X�,c[T��T]g���ES11U���ѭE��1�Z[j���EZ�`oVL1#��gV�E�,c�Dj4�TT3�౶��
�TEb(�J�-��j9T��0H�EUG��ZV��r�����2�,�ܱz��)�kE�0B�UC.��X�D�.��A��b��F��81�[n�E����fU֕J�b��
֍֏",Q�*e��m4�$�I�߄��]������RoJi�gU� ��kL���F�5��>�&VE���������|5�u�}��9)
��(L��S1�/�թmk\m|��}��f��؄�i�9;���8k {�|�!ʹ�@
!�7iH��Af���r�l$0���H�(hN����k(C�C�x_��6_���;7:��]\@!T�H	�U䵻oީ�}+q^��5G=�\_Y<=�N<�i�f���E�t=��;1�\�T��Bt_FO�t]g8W��+�^���4Ra��Pv"e1i��΢=�S����ka�
C�X�v\k���Φ5I5ܺ�Z����/��L{��O�����G<��U)�q�|Q{�p��JG��n�5o�Q{��y��DdJ{qQ��w��j��&-���]�L�b'ɞsMŏH1�2z"<�ώٿ{�~��{;��61�����嚳o�|[,�g�K᯸p��s `W��.�5�3���k
K.��a�@+GBa���(	���M_`��5^�f�#']�Ly��x��cT�Z)�Rk�uR^��V ;����~s~�w��b�Ji�.⌇�(��Ir��q�A��\[=RHU��]2es�W�T�M��$��bhi�y�����R�-[\;*.��'�݈z�L��"�s�1�M_`2ٚ��U9���Y{c�CҚe5�T��M��uw�b�V��h����ޔޙ�gpfnh*8t�����v�4��w��w��ǹ�^'?W4��!�԰��#۞qv{�Z���g^e&Vz�ļ' �-�� 7TH�R�KQ��[ 8����_c��_-�5�ج�]�LY�[]MWp�6PwZ�F�L�bKBЛ0���w��i�@����f1-�
�nB��\LQ��#�0Yt"��v��we(�,����0�l\�m�]�Bh��Ff�.T�<͜��0�Y��u�vBz=��0���Z�kse��]��*�	Z�s�mt�7mS;�	U���2��S���Oɋ�`�֭ö1��r��5�B��Za�ԋ����_Ͼ��w������ﶗ���7���Fv����{�[z@ޖq؀�^j��"�l�����@nׅU�DTr���f[3�W��)���\�`G�!��~n��P2fI{�b����]��E�������=(L�2��@/u��]z�r}�P7��L�eT�GLVŅ�3��&5��]��?�$^ 2�m�*�UU��3��Hݝ�-��WyU����b�^e�"^�E� d�@&� q�Cy��k�Nƨfg!w-	Ә$b"�]&ӏT�R,P�u�y�_A�΅�*���=,5�&!F��	�2Y��m��㇧���:}�1u{y���]���w�%�����p=����E\��b������C�=ݿ�u��F��ph�{r���q:44��Y
Df9{Pp=I��so���꒸Fvs
��L���U�;�1QV۴#P��2�S4�Y�;_�Ӂ��[���º�+3XT��0�ƪt�:�����آ���C@����&��l��:����-���6�9�[KV
36lw�Wr��5�S'=���<�n��wnV�L�ٝN�;8
�W�L���OWP�7��bܤয়f�y��K�Հ���usb:m�0F��Z�X�-Yt�(F�W�F&i��(Ke�U��e鋫�³6 �w�3� �/(�w&�Be2��쮯_X|P�BN�i�K/E����O��z�0�1��q�&��ϒ�tͻ��Ḫ�a�˟#���P�s�|0sH<��u4��}�����:�eZ�CwדY=��B�r�.�\V��K�X���<V��R�+�8i���Y���SЦ�d_�u:��3�N!�-33��ä�Qz{j���N�J"3��Xw;8�Ba��:~����Sfm��RA��3/�y�Mr�����KIL����oz���tXڭ܄�;���:�A]ۙ5>�����o�+�9�΋�Y�A�4���,"�[�scQT�,��ΉRm1+wd���F �7@�LX�R�T�]�Z2}�3F3����:��!	_�;��a� 7�3`�+�;��V<fC9���Ю���zk��e�Ws¯4� 8�I�#�8?=�S�����
��i���]��9����w�=wy�$�(L��fT��O�Tzc�x����m������^�*=}|�q����������!�)���Rӯ�J'g�E�{��}gV�w�-\��D�g��u����:7��˓��6P�˗��������ƪp2��uOn��^�*/-r���
��2�w)�&qp���gn�UEŠ���ێa���-c�Z(4�j�wb��Ơ��nR��E�7i�}���?����ʭ76�"{��]�uo��\k�|1���ɮu�U!T�<�N掊W�{�z�O\X�m�m���^������\m�����d�y8��eL�5��ղe�#�tv���MצtW6o3U&�L�g�QA+�������gXe��v��1�<;6�"{��]�4bM;�����m����Pi�Ʉʙ���͍��Z�G�fV�f]JУ�]���z�� �G��o�\؉�ȍ�;.�ٽ�݁��C�u��}j៶�γ������������6*��3n�ș>���mN��7x9��fA���7ɇ���BSt�׃^&��.�],�ag��`%�Z�n�qƆ����N��
_|Z9FY���6����ųV~�c��Pr	��z��
ʺj�Hv���m����V�5� ��V��5v�bJ��h�i4�� �3Y�hfճa��+M�U	�.6a��FbQ�����V��h%i`Bmh0%�����m���f��;d�Jl�4L�6��vQ�j�أ23Y�Ciexv��3U���>��������6�:h�����f�GM^�Xի
xχ�L�y�g�C�4v����o��j�D�����/��)����]1�-���<x�Y��b�3:�"{��]���@MEQ���}1n�����; ^���L������
��o��|�n���2�����
q�����+q���*=t�_��ng���JN/bo��������0��g	�
.�MD�j�W.�GэT|'2��!���� �y�(L�������aغ�
�� ���Y��Ǜ���ƗMi�U�c赲��c��i��o\<#	��xEsnIe<����辟vz����~�&/ݓ����5�fVBe&�v����c����}�5N?i�1�%�Ԏ��3��G�R�z�<��cX�znm�G_���v�z�wOo��ە�*a�yU=[��4�eUE^kT�sxUC/�|�؟�ŗ(k��@U)��L�{���׮�	����L����l�mc4��7���Rg�Ni�oX�ڕJgb��mg��עUw3z�,���촊�&����UTL�ǳ�㩵����q����U3�5y�Z����3��b��/�<�A<����`U	\�l�m��`搊K�t����NK@r�I�����șCX�.�cv�c�<���y��w\�*��zZ���W��i���L�P������nyD�v��q�)�j4WG<��_������n'U{��	P6���n�K��}b�R��6Ӑ��t~Բ�����f{F�<qP�鐫�{q� ��� ��.��|�>�J%��z#f/A����a�&
��A�T��NT��R��L����\�W����^	����s�5K�H�u�~ג�w�\�u�I����32���h=}��=?�m��l�ޅս��g�g�zmjז�v���>�rD�>�9ӧpEcg�{��{d�#��M�0��CE7;GkFʺHn��e��xJ!���?z~�_��m9��'���=��&��FMmBA��)��r�IZ��1�S�`��̌�ٗԎt��Ra��c�Խ<3o��䨦Cj|Z6��d=%���7}ԽQ{wQ>�ۖjO���l�}��Ӗ�O/2/ùwZm絎�uw<��45�4��jn	��u^0��������Kˢܜ�P���7�<8x�K,3ܜ�ݽ���������G������IfK��@z�& �BeL�f�\�]&��V���Ź�'ѝw�Z7��.�*�����	��� ���|��_k����-Z�%)u�X�H�u�ܙ!(lb'�H�Yg�'2�6�Nw��"o��ƶ��������N�/zL�l��W5S�R�vP���c'��SN��]�����>MVf��l��U�&26���.-����	�$��뫎��w��s�]-���,�S��aR�	�&P L�ܝnȖ#u3�[�g�ە':h���L셴�g.����ztW!�32�33l w�_aB{�����ˈ\�޵��eL��w�?�����3JL�` fg�� �(�{����@?�

"_�`a�tD!�tr����$!���C@��1(���CCC(��0�J$�"s��d$R��&A!�eRDXB@U�!�$B�pB��ET�8)�� ��q� 3<@�H!�@S������!
+x�*��U� Ua	XBEV�U��C�*������!�B*�*����!"�H��*�! �J
�����! �@�������!
�@���(�!
+J��
8�%EaXBV�� EaQX��%EaAXBAV�U�!EaBP!� B!B��$�B%aBB$ B�H�B!P�!B�BA ha hdB��B!�!�HB!D�!B�HD��x�(<���������J��� 
 �@��kW��~���E�?������P o��?���������|z�~���*�a����g�@Qo�EAD�@���?�|��O�/�O���R� U��}>�?��ć����)�?����@s�~!���W>��"�,��"D"C $	2	"A
B�	"D�C"� �	$�A �@�)�A�!���"@�,�I �B�(H@2���0�2�ʐ�2�2#*D#0��� B0���2��!
J�0����,# B���� ���0��) ��3*BJ2���#*@��,�J00���2����
A�3
�B4ҥ4��@*�?z@��i(@�dD
JU
A.��������؟�DiTE�@)/��?��?���}���>�����������`W���?����>���b~������������_�
 �����O���֞�TW言*��4>��@� ����s�H��� 8��؜������ ���|��'G��> ��PY���C�����*���(>�����>ï^����I���?�=P_/����*����o�<'ڽ}����zO���Ϸ�4{���$����*��^��}�>���������~A�O�>_�� ������@Q~���>_W��� �Z��d�Mfh�U�~�Ad����v@�������B�(
� 
      @A �$��    � @

( UI
7PT P@� PPU
( P*�@ P(
 PHP*�����QE @�xU�U
�RDJ�*�%"���$�(TB�%RT�����(�(����$*�"�T*�� :�:��EI@�@{�Q�gI���reJ��	;�$�Fw�:T�v�(3@��gT�QK��H�n�y� P����� ��=.f��`���PP���$��@

b��h)k��*��B]7�����%E�D��h�C-֤E�4���R��
��}  >�)T@ *) ���J�ݝ>��9t��(���4
]�R=��pIJ��
��TWvrU�I�Ԏf$(�ʪP�(���� 7R��Q}��ΑT��R!p����"n�	f+�w�wJ� wgEa��ۨT�
T� �����RU�T�=�T�t����Pp�TS��݀tq�B�Bl2�n΀ R�"�� }w��wQE�]�UL3d��Tv�Un��s�UWp����]�u*w`�� �
�� ;ԕU��T�T%%=�vp�tj�d�� �q"����Хww!J�n��E*� �����E!J+� p>@# ��
  ;�9 � � �gAT�lr wg@ ��= < �� �P*�!���^ Ǡ�5@݇AF��7R� -� ��4 ������+�G@@� 

��� �v �� 9�"R���݁���� 1ܪ�� m�@��2 � <     5O�A�R� � �ɦ` j��Ȕ�P       =�#$R@ �     l� �R�`	�� �%?R�R��4CL�d@ ���d2�2d��jd�M�SmI��{����v� |a��M�ãti�tn��C/�$������} 	!!>�$� H!��HHK��C$����H׳���Q�#�4�����̐���JC�?ڈBHHOK� �) BHHM!��Z���1��{��n������g�r�^�f'C��ѐ�J�P���u}�}WӅU��k���X�gC��ce�ܱy����4�:b�F��u��*�����Ne@�i��m{X`��9A�r�A*���nbh���a��,i^�ãoF���u�[ͼʖ�Qҭ
Pj��D�6�6�u� �)j��V)#�4�,�f�kgsok��*b�<P�����cm[�Ę��m}�mW�ܯ��v���Y.��Y8i�X.<ʡ�j�6a�KfŚ�;�ڭ�z�of�^<�i�ԧ ��b4���Phf���W�Yz�=BMNZbZ��\�E,�Ut��QBII̵����I*ݨ���̶�����d�n&2���sv���maϧ)(r�Ĉ�1R8^e:�����Y�+7�2\e�N�S�L�m�9����ݏ$*�8�˭V^���8�$A-Dlhr�J8�^Qܸ�axkp$��ţM��гN�Q��)�7)�le^Rď�l8u˃)M�DV4���MWԦ���c���ⷧ3u�ob���	�f�q?�t5��ڒ���]]���J�:�*7f�:u3]+���X�f��yy�"c�`O1�͂��vÐ�N�f��5�p�.�t//]*݊�Vӥ_S�4�<��X2 �4�[YF��^!�n�����fy*�n^^JYR,�b`��ѬkY)�-�P�?Ӻò֓ҏx�X���]�Z�ñJ�Yx�3C	3b>JEJiX��b�̼Ov��udQZ6���47�UK������#!@ᳰ���F�Ua�������Z[w�4l�]�ֱ,c+�ԕT�(�t��Ϯ�/��i��;x31�ĢJ�e�R��N��EH�g
T�T�v������sb��A	)I��Ӥ�G��4��V+:���T-f��P�m5f�;{wL�ão�JV��~�������Gd
){���νW��+0�,Yw�a��l��R4��:r�_��n�j�k+-ޱF=��
���e&f����!,)J��rVb�n�$�f(���cX�����L��n3�eO��X�ee:˫v�ؓ��&X��m�I���Qܣ&�-�U㭪�@��Ɲ!�8p���KIʉ9k7"�[w6��᪣�_яq�u���deD�I��0V����'(�]en=x���d[�B�S	�T��U8�R��3��d4m깃6S�%k",���+4��5Jl�^�V�DJ��
�=��ֲ�e^�[���Y�CL�V�8��iyT������z�;�M"n�]��n�k)��/`�v�VV�����y�Uc�������fgבʵU�)�KM�_1uM��w�^X�h<��+�D�r���2��lB/r�T:�"�Y�.V�wrU��E��T�R^m��]ڒ�n��Ջe�5[
��!Q��-R�[P���a��*ǐbV*}�Lt���t��2�	�t�M29!拘^�Gl,�n�S;T)��^]����r�:u�-�D�Wu�2�V��2�p�I;���{�b�+(� �����f�)�魬����91R�O]}Ys��wYW����5][oVK�X,ؼ7���bQe݉Q����wp�6^$YŦ��l�!-�ӆ�^�����,��Ōޥ��2�U���OMn�%;�n�KʭkJ�B^^�����-ZTIa]�h�D,S߲�qk.��r�����Z��8��7D�v�0�5�[r�feݨ��a��w,�U��e�����݃R��v�o�F��tj��f�v΋X�8�1����H�4������R�)U�&]Bs��8�N	Q
w�Pܲ/o6f�hM
�d�A��%:tԪ@�۔"֠���v���y!:e����I�7'�<,�vubĐN��Lå��Z�%�9U���l+�MyXt����/3tFܻ�D튫W�eʴYF�����T�ǲ�Av�))Z�,)[4+ˉ�&�e�T61w�nv-<J��]]ʻĪ諧3*PW�㒠т�յ����f�т�[ˏ2�Ա֜��ifMw�P��۳D�G�K�r^D�,F�y*)tKҦ��z2��x2]��m�C��L�T�E���^U�W��%,�v��ЭN0컪x�1}����e��J^�b�L���ʦ�`Y{�p^�Svcʡ�ESڣ��w,�w2]���D�%bγOsi�wZ�ڦ�U����de�ު9*0������0ZG��m��N�]]bF�4�J���5^]��*��n��L�&SK4��%ЃR�a���$R��Wi�6���Vn�����aX�bܔj"�9,��Ղ���/�%ean)������mIZ�ݪҖ�ð�T.�^՗����7t\ٴ5��bl�Y���i��Fm��B����
�LJ��pP87ne���-SvՓ-l�n�V�ǔN���@S��6�	8ʖn�u)��
�n5�C��M��!&Ժ��TNI����J΍خ�=�ef[�bG1�:��AK��M�����`��aP��B�ѵ��3�B���vZkn�'���":\cohdKc.U����;q��n%�lMe�r�P���j�6���V�ouಜOD�J��A *�4)�C�$U���2u�(ޅBe���0�jUc��\g�{��7׎*�HC�.�1�G/��ܫYN�s]_Φ:��٘6K���w�����n'%ۙ�.r�r�D���
�tj�Ċ�[H�5&;&�X.,���]n7Z�u�A����r�n۵Dh��6a�g�0Y�/ ��zlS�%�ӒL�Xx� ,#7^G�n�6N2l��`&�ʤ���K����]�����Gtأ��`�0�[�j�ú-�wp�!*M$m*KMQ˴٤n��[��T�B�TM�)�xlPU��T�e���9*�qm5�I{krڍV�m3J���X����^��<�wn&	nT��zY���)h���x�D6,Ս��U���BmQ,<�4[n��&m�An�#���7W(h������pц�+��UB�'u29K芅K�B�Se[n�@H�Mi��	:��p���j����Ԯc͹�]�[��6�j;ڂʇݴ��v�1�a˪�f�cנ��X�r��T���*{n�`�a�{X�"��!��jlF�ڽ���x���N��N�0��H�;BD�J��JUL�f�r���L�x��̗*�K6�5T`�˫�(�we��f�T���]�Rr����4%�ۛ�bt�t�����1�lZ�̫(K"㨮`�m���7����TA�W��j�VF�J�%�y
z����3*�ڙE��X�CW��ۊ5qG��a��pXy��!���[�R0����m�2��N�I�%Q�:�3\T�§���S+V��@c�E�U���2^����͂�KNҔ��Ҹ��F�Y+&ç!ٚr�LD�0��A���5un�o�������Z���M4�@��T�Kd�ˑ��<j�%ಝ	��*��v��1eJ�q�6`ϯT�Ț���n�7vý��?��w5f)9���A��b,%3L��LK����p�	�EJ�UFj��w1AD�w�t��Y�NUPfX�R����S2T��Q�̉
2X5U,U�����7�XTܑqV�h���x�Pg �nn�!�3F�ä�H������*���G�D+7v�4���v��-�B�IRKh�l�akk-ej"�I!yuM���IYxT4�	�Ej��ɛw�X6��O,e-8�.ͷ.���h�Y�+�mm<�a*Y�Z˘�eӔ��b�!�{������h��llWNe8~��F���š���N���W4o&1��Ī�nI��gj�:��I��Un�QuMhuX�ٶ�j��n�'I�Oe�x«%跖�Q��#oD�eZ���(hE`yAN�[L�`�xl�sCn�D�ETD��A"�Q�F�æ�afn[��,Y�h�w#��Ma�4h\��PEUF�:�;u+㘰�`�Ze��b�vА���J�\Z�2�,�q��\��l'���J�;�ee٬ڬ���Lø˒��\�+5�g�ͦ�A��N1wj�XU�|��5q)�T���.�bG.830�V3A�{�,��Wn�+n��m�4�4�j�N@V;�f���[�#���op�5����cS�b�Cm�ͼ���ö��3AAhB��������L:n��b�'� ��`5AnU�=� �6����)U�h�eL�!��w�m)]�H��]�
+%B ַV�n���̲m��U�j��&���/A���٥��n5���a*�ln^=�+�K]ؐm�R��nk�����vv��{v��	1nM�%��mfT�&�O �C"��{���V:&��#E]\o)Ʋ��8���q���t�Q�)�QAf�S�f\R�?�Lj��^c�st�i���cTE���з3�*��P�"��x6A.]RyH�Z0��$�Rf�ʰC�mM���ST��^Y-йiZ� MQ�J����52�II��vE��nl�W��v�+Cǂ�K���r��z�knd�0e7k��wxٷcqn"�է��"Z���ۍ�DU�Ԏ�q������+�����S��nK��)��Q7�b�%��i��[�Z%'x�C��R���*���V]���o�U�nK�p�
-:#NV�5�طyy�	��$��l�6jS�q���M�W*�ʸ��,mj��L�X���.��<�5�mKNee�خ�[��ZKn�8�Mdۆ
�*�ᠶ��șM�����(r(�eU3Nl�ȑ6�B��)Cm�l���VX����5z��]�Wg0��]U2�<�d)��
��7�-�deUeiUR��,���ד�GEie��aRU�uv�r;���환�;�*Z[�(Q���&��7��B�i���-�@��ƪ�sr��R�}o]��*�B�ڦ�ɓ�)�&jD�7�L�!�����Xoe�i-�]P$���5G�x-7����a	Hb2�N
����ܘɒvj���Ai6Υ6���(:�#���j �8��J�ő�vk\S]��ed�a6�u���9u�mY{%��Oa�Y�r��eSV�8AG.P�d1��M�\ܙ���6�݄�'rn4q*�����ɕ�-����7IՑ�kR��e����<�rl,�z�i�Es�UR��0�-����Y��i�Έ�֓�iׂe�(K9�a�@�(��e4�c*@�	�쫵!�I���t��tbU�f^سd�p#�੖bW�
z���wJɤ���aݗ��#�GpGRV�޷a��̳tp��^^�Z�n��s/ld`�k׹�*8��L��U��e8�L��,���B�N�ƌV�E�j]n�j:�J�9��X��]��^����Ի3+fC����EW��ڹ�X�T7Q(m֥N���t�oF�,�f��D�����H̫��K����]]�����6]�5Vޡ��Q�a�Y����6�T�/l��x��p��l�7�J&r�Y((b*ʆ.�`ӗW*�gH���r��pU\�y�
�n�eei��j��,=�ICl]S[.)�eE�#�y�+"B�Ͷ�-S��!eUb��m�řfT��ڻ�1!�����ݦ�6�eRr�1�����wx�b��nd�+1^�ȡ0V�Ul�ڒ裌��˭��Y��rث�%I,os���V�'���Uv0F!�����2���U�̚"m�{{u2Y�3tL7H���n��ï%ʻћEɳk$�Vf���2��A��E�`��viKYշ118����H�-U�*
���=���fu�4��Tk+`ET�ݬ�"F0�UL�c4���w-�%�[vP�1]��\K,�wSFCa��v��e�4�9y+m�6�n��*̪tFF"���T����W&ۘX�c<���&��G1�Z�0���QVވM�*aw��,5[%�S-]7J躖�Z�f7�-$nJ��eZ���E���M�$��jֲ/Ff5VZ�2ܫ�x-a�
�����v����b��������y�r�ѡrޜQ�-T��&=�w"yz��$�$�B�.,u���rl�q���/)0Q�G.�mn,������ֲ�TU�Qn]�eˢC�VY!��R�K�����j�Př����i:�l�7.�e�œEH���0#�tQ��䤊{Uy��k7#�4�6a�U%�R^�����(�`Ub��t��cٌ�$S:*�\���7Vq�	�h=BZu�P4"�V�n����W˖)ZU�I!����d!A�k5ZA�8.�m]	�Z��RU�\m6mT�TV�B��Ȉ�(&���ʻt�V�`of/���������{�BD���j��Q��XY�{s!$�d��dd$�XI� ���, �E�@YUEU�]��EwT]�$�I	! � 	 �\TWwq��qW]GWQP�Ȱ� �I XH
U�]tTu�Ew]WIH $�Y$�,,��d ��H��Q��QWE�t]�q�]GUW]TU�W]E]\wd!!$H �RR@P��HY �H) H�B(I�)$�,���!$	�E�AHBE���Wt]�T]�U�@E�) "� X����}�����Q��W��P$��������y�������C����	�� H}g��?�������I���Pc�K�ʇ.*�����]��q��u�s:����l�V,����_c9T/VΠ^UV��ƬKL
V�%ʨ�'N�Ҩ��T�T_-�ͩ�xKc1n�Wr��w۹�+��F�mS=*Q�ni�U�z� l쭗�ަ�rcvD�i�{v3vՉSk3��u��C�'u�U�emY�+�=�Aoo	���n�6v���C�ِtwB��uu�ķ�%�tH�ҔQ����L�md�w*�P�b���͓9�I��L��f^fi0���9T���n�c��mZ[�v����v��6I[�mF�:`�2�s���ُ�D�ǲ���7nhЪ�u98�YSN�\�J��n6���A�!1A�Ĝ��#vam���Z2����an��)��� �w$`w3�͈fq;+x����0�y�p���Z������yg3�<���	:�x��.є��|���D'B��c##s2,G���K\�U9WU��w_i��d����uq)�H��C���w�w��(�n]�-:nU}�ҍ&*ކ��T�L�ua\�f���nS[ځ���^\���ٟ<#5��]��:1uWA� �o\��T�-��f�ԪG_^�T�|�^�1����7�]�K:q㓶�Ek���b�Am_+�c�S���i&P�֬�G)Nt�O����5�/���5ʨ�ޮ���T쵒ٷ����osP'+�˫�gl���T��*�.ٻ�6���o<�,H��`�෻a�$Z�E>;rnZ�{����n>�f�P�ƫ��Ȳ�^�G�a�($�W���������R�͙ͨo�K�uu�+2�H����7����w��&���Y�}��V��%����p�N���]Q��f����i[,<2��(��1�_`]Qgn��U֋x/2'iӪ?&*��Fg,�ŗ��[��Er���uI��s��|��w-aX��j�q��lK��X�+5-�["�z�)B���gX��mt�R[�n��N��3]ݛ�U�w���-�+��py��
���P�2���Q��C�IMM߸ˎUbJ��"�QfV ��)Y����a�d�XTd�Z٤����!e�
��N-Y�p�J������Œ��.��\�3r�]�q8���]%f�u4�ۏ���ׇm��N�=1�!�jf�˫�|��v9C1�\����/Fb�K:�Qܭ�^���u��X�ͭ-������X��ep��a�+��d-&��5�2%j�5y�Aگ��R1B]'-����k�6Gq���i���oL�uauwv�w�V�we3W�P��q�X�ZR��3h�^��Ke��>���.^U�t�B�;��MuR�;�r�S�V���с̹�0-��]�tS
�.ˡ���W!�������ڠ�cbX�CwC�I�S%e��wu�+[Y�L�{@���V�D)�]�rs���ƪ�ml��^֨���r0Ղ��J鈹����e�:Inp����!��i�j��˺眅�|����{/o�lTn�m�Lr�ww���{�����ӽܝ��/�uu���]H�ۦR�\���M|�eM;��$�Y��op�xv�i��U9|��H�c)A�Ǝ�WR�Ն�l�W}�t��/��Ě�s^��y!#�N����ε5�q�}�x�;S�vW9�i[�g�K��-f^\�\��+��gwv����=��P��t,J��$B؉�Y��ע4���-x��Ht�'!��o�E��M����L��T��պ��.��y^r�������k�����������J��\�Rz�7u�l�R���'I�p\���Ƣ��aaW�]Ü�ͫ���M5ܨ�ଚ�l��V(3�kQR�w6r�Y�2T]M�����Yz&T�._o3S:�+ڹ5�&gcC��ʫt�hѽ�U� XO~��Z睧2�<ڶJ�|��mfk	=�Ӗ��-m���1��k(,I�u\��z��n�!�.�AWZ�:U{T�ȽwP\�E�,=��� �%R�ܽ8&���ھl>2����dv�83�j�I��5;f��%-i����6�_dS�l��(6��ٖ^\ǫ�mj]��ׯ���ط��Oe��l�y1a���&�����R���j�%-��F�/d��jf��3]-��!q����E�ӦjS8�����-D��yz�V`��n9B�LK"��Y3K���FY���p뵉��C�A��.�g>���ΪDF�����K �a�]�t�
h��smݒ�Fe#e�n�Ӳf�R�U&���[Y�I��%5GX�͉eR�a�'T���4�|�N����&�+����eufIt��k~�feAu��yw�8��ҹ��v.*��1Ι�p�gqnm'�REA�e�h�ʷ�p�a�����uָ��3ӳ��V9ޱ��!.��AԹ�aC�p�A���v��ܚX�A���q��C)%��י�Z`7��J*�<W���P�f+KT��"�]g:v�c�u>S�w3���8��ӻiwC��&n�F���m��wW��fV�ʫ�֞�0��z���QI���ʷ9�b�cj�J�m�ӱm���Ut�W�^fR��\��`�RwQ�cF_K�4�ɾ���nW��ф�
��ٹ\NbYGR�T���p��4_ZcNQ�t��aBΰH]��B��w:��o��ܦ:7���+�{�&Ĺi��ۑ\�k|��{�ei:�S���yy̾���tgU��(nX�t�'<Ml�70AF���I!��<�D-c�cu^on�{�M͌600b&�@j��(�ڈ�c))s��U�a���cT�mY�S�Z�[k�q����ħb����ЭGoK��y-��ǳU��eQ����&��)�YN�V�����VI:�}��[�Z�Hpӫ}����f�+X��v�K%��t/3��t2ud�6��Jb����
�ܬ�1��I��N���:n�&�w=�ۖ��]�fӺ�QtiM9�ʗ�g�DL�h<��F7Ϸ�<�̫�|n"/����َ��A���D�S���U��A�\�m��V+�`���_ke7�A|7v�f惫^Tt]�Է�B�+e��'���4�IH΋��ry�*8,˻�t�3[oPZ��cr�T��:3W,;���Rc�Kv�
��V���N���).7G�}w����N��`����J�b~�R��Rn���(Nű4p��B�Ԃ�yPU���oc3ww;�`�ã�Hg%F��tv��	��3yd�V�-5P�j��.��'���ΚUC_$�i���9}bP��5L__$�a�3~5&p��"D1kB"�u˻=w(s��)rSaP\#-��Q]va�2�d���ʧl+�����<��TsV�,czqH�j����'}��'u����"��}����B6�޷�mCqYඔ�I:�ʎY!ۉE�O
<�oE�5�,jhN�ԩ
�=�(��w�c�t�!��G�[��V��P�yw�w�sNna��HB��!ok9��w-��)�#�NI����e�;�핫]x�0��[��siH=�4�ڻ������e��pŹx*�;� uYg���x8�v]
�g5��3sr;U�R�'\�ٽ ��s(]����]����^;/�n�-�<��E���Y�aMx6�ee��7�rHذFvW,;͌9G�S7F%w��K�����i�eb�j��K%#S��(өNUS	3��B�F*�j��M@۞��Jƌ�YO32�gETcvV��b�U&�𠠥Hs]8dU��]\Ԗ�m␤�Sک�3�w%���Vڰ�K�4�}�ǁЋ�w�x��ͮ�<Ǒ,��Ռۻ��O����&�6�}ˉ�!�ԛȶK��.�ѩ�ƍff�Z;�Z`�e��k.�oz�nB���gr�]�����P��FUb�IzM���٫j:�m��86fP���ݨ����oY�'.�Bo0VM��]����e�9��eŹK��Y��0�kZR�ނ�Wr��}�gA���<�-[}Y3R�u������[�R7�k.���Ŏĳ�'t�#r&.����LJ�B[K	�tP��5:P�ɭe�G�Huk�#}��CU��0d�b����kM��4>��WFzƍw�8:�����f�G{�$*�3�KV�}}CH�\����K�΃B��GE��+�ϫ��d�v��|�q	bn2��t�iZ+j�ی�KfnC��V��y���~��{��w��J�J��dK�g$;*�BN�r+�໸�<7��@�^u4)��-^�vV���9)ͽ����oh�Cq�A�g���]��f�=y[j2�>�\��އ#nhWk�Ε�EՌGd���ŕw�,fL����@Qb�r�j�7*�^ՙ�tu�"���ڎ3	x���U��KKA١�B-#;&:���OTfD9�)�eJr5�I.v����Y�9l_G����T�,K{�֫l٭5���ڜ�L�u�vt��Tm�u/q;]W��Y̰�M�qV;� �XF�/���U뱌�)�G	Ҥ�]}��4�{aГtk�Kn��.H�1�([9���i��5�d�"Q�MIz���g-N�i�Bj�X!?T�"u[�4���'���Pҕxi`)�����z�P�Oh@����j����:���-M�)eL쯬[}T�H��r�y���dMj�e��m�6����9eI	͚�7�'S2�d*sQY���0�i�͍��K\�B+��%���x�8������H�:��pӫ+�!w]�d�����/������V�	
%��C�WD+�ż讼o=��%��U嬧W�u���J��5��U���Ɲ0yJ8�$�d���o_>���|&��ը��H����Kb��fSn!�%�f-:B���T�wJ��m��V2i�ԭaw��l�����+��KT��+&���.����ÓNJYch����!�+/"c#FȪ��_	4]��A��M����3E�7WL�"�y���6�ĆG\fh%�ΰM�u�3ۛ��R�X#Uˋ�p�1�v8n��z§�	v�0�&�
�U�j�����J��3Y�6�`Q�4A*�!4���4��N��ҭ. Pm�1�kF�u���4:��Bl��/m=4��J��Y¢T��Tҗ���vA���n���"T��H�*����pgcϢ�!E��T��)�Q�d9F��{��(�Ӎn�(�����X����ӫ�9s���]����?Q�%F�L��qc�w;�����2��q���n�ۥ�e;`��1�ab7;ln]Tr�F��j��'��5��7��JR���Ѯ�$�κ7�=۝b��t�R���ҫ�W �个K��n��'�#,��e��~@��r�A5Y�9�l;���lvg6i4.ثk��W���WQU��E(���Z�$��2N���7�+��T�3��D
T�,HBrq�GUe�TBi�Nټ)�Ӻ�5�"E,��J�Q7�vTp���i�F��3uŋ����iܬ����B����ea/7xN-�۝��Y2=&��3yn7O{YT�*���Mn�N%�l��ON��HYWݣ�f�Ne���{T��j��X���K��x�+{wq�ᳬ�y;�����q��_!�+N3khsͩ�%�|�������M�aܷJe�s����1Sv�;W���2:I�0LiMt��K9���p.[g*M���EaN;ȋ�`U��u�/g%-�F�
�y�h1d�X���kKaFc ��:��m���0%�N1v�(3FV\�L֋�嶚����l���*�>�T�WoPe��l�uJ�*����Ă�ITim|�귔��W}OwN3	��mb)i��
IY��oP��R7SUuݘ����h�f٩�ew&�*�v�;Ǌ�e�t�
��l4�&������`��N�E��m�'�
�B�l�r�V�@��y��d��S�Շ�vN69�'4`}N��_t3!Y�`x��d���|��u���+���.8�;��n��w��A�[��U���5G��*R�;iX�ٗ��fS&a=�Vi�rI��T5�7
xD��*�z�Kp����h�ݲn�wJ�tF�ܕf���U+��0ee��*���Xi����gw(�(����J��R�����mU��-]S#W���V�հ%F�[��m�Zr��r(��Qb���,nwmA@Q�[:v��ZD��\*\��-'�ؽz�L.��V�Yl��++0"U+;V~n���b�Aڵ�Cݱ��-�fX��p�|%,FѬ�uF�s0�ʕ�-d�v�������V(o`?p:,�*�Q+��*�=�6�$�%Jm�PG&f^�η2���sw	��p��j���ct6�p� ���X���pk$�Y�5�[�����!		�,��z$���
���O�)�ϟ^i�s�9�X\�l0�c2v�l���u�b%�m�jA�kf�c606���^[�fb�0ܶ�e�S]]T\Ѥ��`B�2�0���Y��MR��lږ��Ԯ`�鵆�n#e!(u��npX%u�����J�IsGC$s7U��pQ���l���ab`\A�E�7 VY�������PTkG3%se���[���o�����0i�H�V1%��ʑL�b�-���Kqh�t����cZ;J5�bA\32�`��׶#��s�3�cY����-�6t��*��t���%ctkb.fZb<����NHP�e�֋�م�l6!
3u��Us��&�$���2-�sK��ib�-k�>7R��R��956�1��%��e9��Bk��� �/&�X��A��.%
,xp\cMMm4#i#c��m,݌kt�:�tC�0�#\�#(�\�KR�F�[��, �y-0�Q��d�sC
��[�lv���г�]��lT�ssqVB#&�V	�yJ,S8t%����]et6�#C�u���ف��I���8�ׯ����1i��1�oW��o�`T�&pŗmcR݇-����]t�iEVQ��&j�֋V�jj�Տ�K]m�^5��Sk��r	-�J��T"m5oiu�^P+-*�2�Z�V5�A�Ͳ,X�\ �:WkT�,�\i�N4�m!b�b���K���mbU�f�.���`LM0�Sa��u�(3C�
˶�qbq��F���B�WRʱ��ы��aq�B�iY�Ls���U�&�1���J�-�/2�����h���v���`�̹������s�K�58�j�iĤ8n��,H�!��e:��7��m{APچ�n�nq ���qHf�x���Lb�&��#�f,�%��#�f;3 $"k��hB�dw[rmR���6�IX�3A��V��H�V�H�R[yڌ@E��
�ET��q�oR�t0�g:�M`&��Rl�m�[��0�"�����Fcv�#�Oy
[����MH]��2�vL=Um�P�7�#+ؘ��r�36n������BQs��T%����`�45�V���(�[���^B��ԚZ0��+-��(��ES��<_-��iuM	n�X��8���9X�e�8���6��a��i���Ґ��=ke���Pfl�4	A:�Kt������^3	�Y�k؋6͐t�iF��/�a�`�[/YB�H9�És�TL�ҭ*��=�0(���IW]+�Va�M�fK�LX+��drjX�]-ԛip$D���m�`f�c\�-+2D�h���ˆ��EQ�E���*ZЀ�@�4�ڲ��:�W$pF񋬰�ej�K��+2�͉�
��u#6�z��(Z��դ̎ļj�g� ��;��؀�SKvDd��ٵ��!�^	�	yZ�幍���#3�37�֤DH�k՘�Y1+	�b�ԘX�Vb0Wk�+`�4լ-*�Is��(���n���7E��b9ѤM�0��P��k�-�*�͙�f�/9�c:.�fZq���1�W��cGH9l�ܹk
�m�
u�[M�˴�-�K����y�y�&�@f»P�L8DKhS0�e�6�շ[��Β�2�s�Y�K��M�����sm���/lj��ˌ�̤6��Q����llԙy1�R�L�v�8�Ѧ9n�I�+1�]�icu��c�ķ3J��u���#�\��R�� /cWb9�2�v�5q
�&���1\륓�R:�M6�H���T�͙���M�Poa24JZg�ΔB���CW������ .#4ƋfL�a���,Y^`^n�o&�(��h�Ѹ����h�QF��4ΌL�&��a-[��-)dX�F4���b�Q����i�h�˫]V�3�z�tt�����H�JrV�����V9I�s����2�f�v[b���"��
�l�g:3Ɨ �0��oP�M0Ѯ�i���ŌU�:Z�ŕ��eKR4��&�e�f(m��n���h9��3me�WVl3:�j���501n`lh&�1�Y�a�����������#�]lL�ۋ1t�ŭ"$�@qt��ّ�	c&���f#B�k�̢ix�R�h�CK6�̥	�(Z����ݨ����+	����G�����B1�5c\�(���t�{;�B�jŊ�긖Ź���m^�#�%5k(ZJ�4��aah��.��N��V�C66��L=e�HJZ�Lܧ4��q��F6Y����2�2�ͳ�-ّ��]\���嗴�E�Fma�E�R���(ݭ$�@�[s��0p�e��!�իq�,n�K
L��KB�,�a���A�%ı05q�6qU�6�6��F��p�%���&�eU�M�B�T��l�0n��`F���
MZ�Sn�&���V֪ٻkKcU[�F^PE�Q���f9M��ecD�0�7	Zd�4	M�\�4�.��E�V�[��6�1�u_+��A�5�ͥ�
��2�7E��,CY`y�J�{3m�jL]s0e&�vD��U���W$��ې��4P����Xf�Q�4Y�$K�1�R��K���Y`G�"�P�te�ku�H���	1abE��ٗ��ˋi�1��K�3"���MiqU5f�M�f6M��]q��(���0��"WM1����I�X����6n�4��,�*62�Z[�J���6E�stb��WCGQεFk-�&/�V��D��T��U���#�v	����ثB��[3l�t��6jW Uم�"�k�c�vs)M�KK��1q��
k�f��6�%�k
f#�GbD�t�g�$Zj$�5㝄(�t�a�]ե�v�D�2��a�I��X(WT�$èU��F������MjXZM�F��5�N6��W]1s�%48����_5�2��m�y�,�;W$ը��&K�T�a�Fb�t��&���䊗v�y��՛(��]]bnV�6hf��6(&Τ�؄����4lp^ju���[iE&�jL�Ц�SUf��e�����E!��x<q֤i��nYi�XK,Ř�IM���2��+�Wkh��n9
��VO6��hT��"35�2�(�X�me���Y�m2Aeې���[au�F�4�R�V���Q�a�jlJ�q;hՉ�����9T�����m�"'��7�4�,a	6�$v���-V���e�[j�:e1)��4G��ѕJȤuh-�݄P-{bƍ+����pF[a��ͻk���� ��F�p�j+6R���b���*m+ff�t1$4�0	������aR"�K��bƸ#r��L��cq�8ɦ�զκ@U���̍v+�����M*�A�-n˰)���dJ�K�藙�e���]nĖ�_�����b`j�Zݖف��i�lxVfR�.�Y��0X����5�����VҐT5Ʒ��
m���٣c"%��0����3X��%ڳ)N�+`š��h�ѥ�!���y��8/���˶�F�.0 ���Gb������e��,3��`Ƚ�\��˭uⴶ:؍�A�ٽ��Nz�l�f��.2���MFSBb#�Ŗ�cfRh��m�u����[A�t������&�[��z�UD#,Bl\8�Ў�m�hs+#v��m�`,�)tU�#¸X�e�$���7g]͠kK���Z�,)t)V����NlR�Ml���0�	[����-5�	f��"D��5m��m�U�GL�aJ[.G+�S\��U�U�f\�9�5��-�������f���fSulwm�0j=V�X��n+]�gKt�:��`�R
��vNu�l�:�Ƭ\�]��!��\�B��[��#�F�� @-���mN4��Ѥ"kk+����ɫb�hиt[LWK��WЍ�!6b�؅��ܮ��X�j�CX����rmR���G���A�T*���:���[bMC�M��%��e���c��R	�M�k��5�8c���X	�YKku��<B;6lc�qf��Au9�pnnQKs��v[�bM4#
ʚ�8V�hZ�V����fF$�mahښ�����a8e�x#F�lY��۫arQ�0�rXh����D��V��qkG)�M��+��ta��Fe����i�i�]�j�-]��0is7h�c�jg/���x�m2M��!�CB˜V��`�\�&t�R �R-%y�f`��P���5�(*Y���tvNJ�blJr�D���-���ٲ��-L�3a1a�3U�f�6�҈ioa�D���^F����)���mL�0��!4KL�X�躭ضō���9��չ�T5�f�ZQ[+���*��������V=j�r�����m�����
�vM��n�6,3.��9b8h�ʬ����l�kuƄ�Ɂ� �ڬj��m�%s��f����VdAdP�mb��f�f1P�9�Z�µԆ5KkcE4]·�<���9���Y�fj�"1eUDQ�+*�EA.�Kno�z1D/[Ioo{bQ?�w�zRr[b�8��
#����!=˰��֓���ւ(��W�h5��ẅ�8�h:B�j���޴࿚��%���+��mdw'-N\q	�9)Ü��mN�nIN�D��,�b�w��J�Y�%ޙ�t��N�l��a�P'O�hr��-��aKѰ��@-��$=����yg�ը�BI�h��F�d��Yl�N���sK��t���:D�4�:'��[Z����q���g��6�Űj�ٗ��{۾���QIq�k��۳��X[e!g_;�^	ͶN-���{n���y�m��:	���H�1�W�t���)J�}���َ�O�N��?��~|��#�X )-p$&� �٩c�u	��-�Q�Z�b�v5ݣ�e��R27%7
�Ju��\�ۋ��Ҍr�BZ�!vAM��!�s�P�зK���K4ζh��Z͂s�ɩW�3��,�c��عnQЎ�¶~��[MXyk��/d�P �x ��t1�Q���j�"GMfl�A��I�PL뵽��;i�KE�V� �k6p�vM�(�[`F�e�%��l��G7����fc��-Rؖ�6�P!�v�8`͞�P@e�%f��Ը�rd�j��(��|�]����u�N��E��Ԍ��D�Tt�Meܢ�aK�3Yt��	]l5,/W��J:ƌ�Ж���u��e%��s�	�儱��iJ��R� ��n4��!�3BR�͖ͪh6Ƕ�e��K��j��.�kl��r��m��2b�x��\�M�sk�� 2�RS
�U�3[ʹػB��2��Η�z���b���+�Dt�sd��^Y�m�۵�fnʄL8G���b,���88�W
AͰX2�]�L݃7^�y�:�.L�`䥻G���Ғ�A��kfw].�H���5�47lMa U�Sd�뭉k����j8�ע�K�U�ۚX�cSn&�)�%(crh��iI�u��C�Ke[��KYm��F+��sQT��X�(\պ����]��&r���y+2�jY�ԬBidն��iAb*me�8�&5f�L����%l%{)kkm�6.\:�L&A,6)6z�0�Z�"5�]%R.��k���E�ez�kF.�hM�A.k6��5�D����6���Dз���d���vj�%���*�V�&�m�:�n.�s����qX
삄�����KH]�[b� ���cQV�lBX��A��PV�c)e)ZRV S�p�%�+`����),KXR��b�/X��z�-�A��e�#[D�%E#cy�[H��^�6��AK@H�R�J��Q��R	xz��ʹ����*�F���o��	�"�eͦu�K�Q�ԷWaգ�.�U����qF1Kx���7��c֨/���Uqj�m��͞["�Ο��9՛;��^Я���X�"�	�
P�F����L��"���5�-v{M_F:���h
��d�䊔0x�=V!�q@�guXH���|D���nj�'�9z����5y����AaDޱfE@�D?I(e�����T<���<��@��D��7��1A;�#O9t�����ag��CPҁ���e�D
Ib̊���V^��[>�oY���w͎���� $�����;j�V��=D]dn�hlG���ܢ�jj�\l��,̬sR]�� fu}cz�!@�$���u߮k�o{!Qx���׷^�d{/�� 6��2#�!���c_z}�����9Z��&]}#�Ċ�w
�R�vJ�n��fJ�uzOˆ�����M�;r�k�ng�*�O��7��OmE�푧� �_N��B�UC���:���L�B �%�"`@0������~1:��߅�<O��ƅ!�%}"
'Qq�׭�h�G~�!7|�'�=�Z���1��">#�
B��ƾ�a�%��A|��V�����o
t(r�3����b:28�����5��#32Et,��Fq�C<�C��Ǯ��,S6l��50�\��CJ��A<@C'_�&~�go���p{o«���!�Q�.�M��Ap_* � ����H����{ gO�܅޽ɎX�j��s�5�~d"��,P���{��f�_{�=�(�"�$�"D/%M�O,�|��wx�k�������K��<1T�걋,+��P�3nNZ^.�ଢ଼����8�&T��W���X�̎> ��Ղm
"$�0ȾB�4a���B �v,�T&���.E���n����W-��.��n����0A3Ә�#,۝�0�}WL��=Zc�	n������Dޱ|A��Vׅ�̕q;��KU�;&�Qt����ff��9D�������m�y�,����I_H�5�f�z��i9̎>?!�5Yp�Ժ�� � ~?I,X9��|p�T���F��"���"�[��V���2>����\���%�`��l�sޫ �B�����F��L9�����	n۬1K��D��`ȫ�A0��]��̭�9V��ZA���d�_��3k�q.���4� ��R��:�"�8�g�NuJ��L����%�&N��*���.>��<�LeZS�'��[k����7j!tK��=��������`ȫ�0��P�"Y�^�cʾ� �S����t��\�u?}`��~�d�`�%�u�-�35��(�Uw�+飉iX����\�W�V��Q��;6��,u���~z��tB���K��9{{�j���+#�-�[�B��
�	;�� �p���$��3�ڬ�\��0���c����l�<A����F��P3�"2�m����z�Y�_P�"�ř#���!�zOY誓Hފ��t5Zr +��J��� ~���6�a��Gu|6��IB����W����s�eb��2���y�xA5�>1� �
I,�D(�!|d��n.��+H;W\'zN�3&v�̎7T��7PDa���3$n��I4�c�T ����%P�Ӽ���I�t�w��~1����1]�Sy��Ϫ�䍎F�/_mH��7u^��翟X5�T�*���H�%�ab.���[�0���.mUX�$���AX� ��L&j&-�Rk�p��j�U�j��
b���YZ�n�(E�t��\[X��l]l��ِ+l����Ѯ3q�Ѯ��[ C	�u �1�Ѵ%�n�T�L]���l�:вĕc&�R�#,�Q�ۑ��M�f��-��U5ʍ�����>�.�h:Zf�J�&A��[�5#atK�`���]�]��=���E�0�����WgEۡ���V-��\Ěp N�}�IB������Nc	�H0C !�X���������X� �	���EV�W�k�������(�J�$AOze��x�یߵ�����)پ��{�3����-6������Vn�����DaE�{�w��Q\�Z�����\��|�-�_�=B�B��J��DC�2�WnY�l����Y�6m��1�N��G@6D|A��� �B �"z��J4p�R ,�D���]ٷ�W.�vZ匭e�pj�@L�e�~y����C���U�"���{�K�M���+6g�7�B�n� ��P#�|~"Ib��Q�D`�=2?^�X���ea=&g��Ž*�1��3���'���%��
eU��q2�`�iR��6��%~�+�D�a�v:��Z�۱�X h
/�2Jś���=��c
a@�{z��$�_�%������Rl[{�`۷����T}��5�2*DI.���OrѾ�Vj��* ��@�3@�SR��s���<�T��*�&���wj:8�0~-�"��Є"Ib��{�=[f���}��rJ{���xW6�h
����b5Bs���S�P5&T��9�MF᥷D�iCYpe�1l��Z�b�%��}���~�3���̑6���[��V�aX��^#�*�/���o��c����� �a�%}"�=�ű�y����1sh�\�;���E�g�&���Aޠ!���3�Ş�G�!�ř A%zWZ�R�F�����7�����r�j����8M����D�9�{�笠���ޱ^�Ed������{�k��������nei����w\+�������@�*�?X������-x�+�hP"~2Kzxԣ#�U���*׈ ��;�
�z�	�	&_�!@���$�?�؟����_:J1n��;u�r�Aj�����C3�ֹ�j�RPZ D5J�lJ֥j&���kClܽamm�(S'����%�;lY�P?B^��Os�e��ciСZ�ÑG���A�
?I*�!��͠\���,�i��T^��Kv��k�� N� ȼ����,i]m}d E��X �!_b� d�d(UB^�Gިg�c])N{�u<�0i��e_��B�"�X�"���g��W������ř�a�^�৹���n�ܺ8Я���|�Lz�LS=f���w�)�!���bX��*������f���^ͻ�Bؾ��S6�Y�.ړ�����[��ҽ�{�(
d�d��_
G�$�1����ckf�N��Y�y�Z��� G��Y�P?B6��i�8�@����UH��Y5j�+GM�p�Lf�Y�jB�6�&�*J��I ��y�	~B��r* �/���޾;*�"h3�����l⼓.9��`��42~#3$Ī'�m�]���q���xh��ޘ�3;V!�\F31T���΀�P� �gm}"!G�%�y�H�[����/{�e/gv^�k��:zŃ"���"$�cıwY)п
���ՄH��]%�ӼmfEli���̫]U;�g;�d2��eEDa��_�*w]y�����8)���{�cs��4(�"�%YIBv���%�Ҽbջ�h�&��k7�̖�|d(��pKqb�ڌj���N��8ch���1թ��&�W����{|NJHM��7����^OX�Ŕ��V�0�f6�AFnm���������Ι��u��-��U�x�W:��#+F	0�^&����4�']ȨJV���
-qML"�f���c6����-Z��rC�Þ�GCe�ܣpLJ�A��`a��f͛��VlS<�b��J�kdnF�k���e�H�M��^��ʩ��0����~!`�l��:-�k��M��7��M���v�� 6�THa�A�jH=�"0��3��z9픪��մ�x���d��b�E_�I��W�a禽�s�KqǕdk���Dc�|MT�V���) �0��	�=��|=����?x�A�X�dT&�L����K�s'����6���@z/��IW�IB��^l��;;�, �s2D�j��p�=����� �!������	Z���Q��DI.��ȅJ��{����z��)��}�L��+�?MR��u�@����s_Q ��d�����"f[t16�X��U��a�U!a�Ή�gm��|��VO>}e��p�/��S��V�����+K|��ʱ"�C�j��A|F�%Y�=޳눥�	>Y~j{�d�Sqbů�ȝ�����SM��j��y��Xw%^w$lp�����b��|�Y���+:Dڷ��>�0��u9���"�Ο�":�S�*����6���D_ d�d(Vxyy��s�e�e1^Ν��tƟM����P"~�W�&�So�	�{�b����	�)�ѣWu�;Ua:�?U�_�9YsWFgq0<��r��H������e�r�ցc�K�W��"DV5<ݤ���kmZ���"s�/�"�A��,_y��1w��OO����{f����%�!�i1t\+H۫l�Xۃ	ͦ^}��с�՘��w�����(��fk�x��yPi��7Y|��r?;�V?��?$��L�!U�(��	A������W�C^�x;���cm��h
��d�En���9e�f���;ݖ�i���H{A���?��9T���F#�T:�q���f�"�d�c�M����>*C�t�j�i]ܻi�[���G·#8���8"2������g%[��w|v�W3/	˷�&v'�j��L�_D�)���ko'm�&!4��ENn���0�(��R�8�:S�:��Z-ubb�zsq���B��Ndy��ܷ�ݾgMn�0�]<�N��5�	�]��4���	e����;u8���u=�M{�S+ʬݡ9�ݾw����P��1��g�=�瓃]��Sr��Z�v���[�h��n��`�mRU����O^S�a��9j�rU�����/��]��\�QW;r��坏eK�l;yp��+�r��n�4L��#�\w�]%�
��(jk
�Kv�9yCZ��=9��RQX3:��%a�ݭ��t�H�l+w�y-T����O/�ܝ�Y���&UX���/E������v5�7��3��Ҩ��MUܐ'��n���7�\l�Q��sUTCSJkvi	F�<	�ջ��wi=�˕�xĮ{[�Pe�p[�6�]X���;�/�2[�פ��5�:�_Q:�����,j-��Yu�H\Lm�i0��r����6)P�7A�$��D*nI2���n�I_ev7���Y��_q�;���B
��/��-�U�uO���	0��ՙ�cב�������A���Gof�=�]Xr_b�(uL�2;<\��%���+�^���(�� k/ooztqY��S�mKoT������j�6��6gNv6�Nanɷ[dI�1IGY�|��r�6��OYV����)�!����J�(|n���~�ok:�m9gqC�@|Ȋm`��mr$q����9����{���E�^i�m�hk!{a{ۻΧ��$u�ί�����o3��?+��V^^S2=�{YE�>�u��{�L��G��yy����W���nK�՝�&�W����|Ȧ�fc��:��g��bbJRLvԲ����Zr��6⓬�lw���<��l�Ё�m����K�}��x��B+�X���=�#(�(�ܗ_mm�����}5%��q!!��gNw�qͫ	�y�ؾ�EGqG��ӎ'۷��׶t�����ݤ�݇<�ٔ|Ғ����qw|�/��E��T(���`�(�:�K���n��^gx�r���^h��
H)�T�) ��<�a ��9�-&) �S)�TҒs�����X烃�p�E�Q
H-j��Rs�����
�I~!��q���f������Rx�0޵p�&FRA@�&6h�;��GI���AyU�)��7��)�B�9�-0 RAH/*�(X��
�9�C)�XR9E��^�/=��t�Y82
��@
�v����;5��|	�mb��@ktZA����.�) ��9p�5) �s�ZA`C����h/<!*&~�DLI�1d�V�F٦�V���i�e�j1X�Iw����<�O�t��$�)�Z��L����G^Y���Rʨ
AH9*�.H.l�����GT��[O�D �#��'���]��4�T�) �����Aa���贘���Q���iI�9��)!EP��pQ
H-s;�c��_��0w� �H�9�ᄂ�P�yF��X�y��]i�o�q ���) ��)����2�H(wݘH,4�^U@���=V{���s�R��<�ᔂ�H�E�) �ʨ
$��¹�bH,20�r�I�
H'���| ������~��k#g�m��Xχi�Y��	!�[��
!I��p��Xs��a����P9�- ��
H/*��
J�;�����:a�z�a ��ݘH) �U@�TAH5P�9p�@�����z�%y�~�
 P	 �������|뻺�X�7N���1��ޫ�̆A����������'����7�4*�$�t�	ݤ�k3u9�UgګT����Ny|<G���
@�贘B�%2�0)Ĥ�Ü�\����QiB��$�Ü��d�,w]7�7$/��;Ǖ���uʭ�k�����f�`a뫄-	��o{�l�l��{�w�P�7�1�:G�L�5��bʹ����")�*�Z�KM�)Y�Ӹ�I���I �����2�Xe� s�ZAH,�O�|��|�3燚��X�#�O�u�<h��#����Z��F+`w�- �Q
H-yP- ��S���	 ���9FA�$�[H))
a�r�L������������F�
AH.�R	�{|�G��^��O��T%����(�/4ZAH,�2S�!i) �����Aa���Qi/��/��~l6�Y:e<`RĤ�Þyp�AH(yE��
H-��R�
a�r�f2RA@�(��©�\;/�}����}�+^��.�{�|	���"AIHS�W2e��P(;��$#I��)��ˆ���r�H)��}�k̵[��\�/�
C`��
�α�aH�I�) �S)��,�]�b�ϞV�u�|;H,:�,<r�RT�E�B���Q�N-�^`i �g���JH(TC}Q���R�$���.d�) �s�ZA``i �`g���[]�d���M��Qiƻ}Q�f�{?|��-<��YC%:`R$���}yp�AH(��b�R���4F�gɍ���WR
��U�dP�MCUɼ��k2��6����.t������P�Z�Eڐu��U�����x��]Hm�?+
QeK`md��0.��رnJ̒�h�%��ff�c]Jňڐ�vզ�Ҍ�Q�g#U�e�=F[� TطQ�G[�Kr�4al;P���^eշ	4̣�%����zǜ���ᵛ!��x3��*Mn��ZڔUк�b����II�G$K-إ�:�!����31CSF��CZ�T��(�~_�g�߼�3TlQ�,�s]Zb�CRkG,!
򤬪*��q ��a�� ��E�B�\����Ü���%'�� ��	#�O������v���t���^���Rs�3���u��xy֫���.d�) �Q�Y���R�T ��9�\2�\�
@�(���Y�JyUBĔ�X]�|��޵�V�=�a �wE��B�%��P7ߙ3燕��u����)!U@ktZAH)��� ��0�9p�<�Oe�f�&�
;��0���T0������w$���Qi ��P9*�)�9ˆ�:��5���xT�eVgE��v8�|����JuUH)����C) �s�ZM�I��O*�) ��9p�AHu�;�]��<ߛ���R
Axj��R�
a��p�AH$
���	#�O�~or'gk������t�^�) �Ƴp�'�����N�<<�����H,F��T�D�AP��H.F s�ZAH,�%<������s��R��r�H��y�9���t$L��UP@���1��FR��#�O�k@x� �n�H8��^U@R
X�L9�\0̲RAB��(�Aa�=G����_/�烬�����CFTX��]�Q�cL�0��X�;�D���=�):	)
a��p�&FRA@��Y����I�T� ��.H.K;����a�u��h�- �^�����$��T �y�C)�XR~Qi0�$Je<����Ü冣���P9�- �R@��w��ڸqӂ4D��۪al�e�"�IEU���P�taQ˺�)f�;��f١�RZ�֪1��@�\��oY�W��>�s���Xw��g�%$):�	�+|�u���}1��uz�א� ���aI%S�W2e��P+���AH)�T+�9����[�ߘ�d��8�ᄂ����L RAeFJ|���i) ����!���,)���`B�%|~��> ��E�'�|���e���lef�χi���)!R�n�H) ����Rs�3Q��
!�Q���) ��aI&���]�{��2p����S���A``i �����Ü��	�&��_n�*W�s�TG�	�2S��
��w�������9F*�����R���ғ��MG�s1���>1�s%���:�k�|J�h��6��@Cg����Ѝ�"�ɮ�&eH$��"$�)u`�f���d����Bh=F���_O��@�JBy��}E@��)���}މxL=��X��Uae49b@x��m|����^Rf.R��q�F?�zA�c{/]:�uy�5k�!F�_�!�b��2�j��G�6BW��\B�/�IVA���E�}�f̙((�U��vuܜsb���Б�7A̴��)3Wٶ���9�P�3r\�e��Ns.��u�����q���u�LVц4�L�)��� ����{<S[0� _:�4#��y�}ކ81[:!�OՐ��M5���T�F�
B�&IVIB�"V��z����9��[��3w�(����"�H�"�0��T��u�z���D0n�$mV��k)]+(��֭ٵ��b ����ןq�ˀ�!��s1I1i�.��V�*�D1��"y�;;q����G?̑ �B ��s���u8U��8���C;��Ooa�f�gD<C�\C?@3?M��p�cpz!��P ���H��%���^E]^��u���6��6B#g�Y�Q��I(O�s�U��@��:�YI_=�Y�}�e�xA��$J��-�� J��+գ6bf!m,*�p�u��7m4��ވ+.��ʎ���e��������^���XϤZ<N5מY���[���P�"󕎕�~a"_�\��z�qu�[<,�
i�$����:u�<��s��<M�R&DDLB�$���D��R����Sg5��� ����v��LY���r�|~�P9�6z3]�fo8Q��}]J
��#s���� �DI,X ȅ+�Fp�z�����A�__KS����N����3T���F�rm�%�gۘ���@8B��$�A�.R��32ƯN���B�a]|�8Я���d�`�%
#���5�I�_w��2~9� �Eo�N�j��k��!�CʡԌ�۽^���ܾ�t�D����P ���T����54�S��У��y��MN�cO��IqF?fb�Bf����G�q�g�mCi�c벎�!�k;`��FR��f�ݫS,�C��gXEh��t���grr�C+{��}���[ȶZ���\��fK��F¶��-�@:��p�LcH�.\D�i	e]k�pM�e�.��f�/���\��h�7v.������v�t����IZ�Ը�5&�f�R���,Q���qbPv�mUB[�\mu�vyQ�"���*KlEu0�f�5�Ji�C:b5��k�e��[E��ŎUCa����θ��v�����nʒ��cF��P��m�(m)J�S�"�hH9���3��d���]F��CΑݯp��l�]S9 wG�~�$�DB� �+�p��9�u1��#�O$�ꅚ�P�8I�� �(F�_�-�/מ# !���y
 �a�IX"J�oOYYYvJ��N��5����G���� ��/��Ib�2* �ܨ�xڏ���:D��H� gWV�]���b��C��A���_O2!��G)�y�^}Qi������3{���}�쯰n̉�ؼ��D4�8#1�d����"� �!(5+���`���e���&�%[��UDЌ��J$�!pL撻�޾�җ�(�J�$B��ṋ�����[���1�����5�4��3�"�� ��S�
���-�:l碳T�_��:�
�����)�,wNs/�!�3���=��gWU��Ȫ96�+�\��U3cC�|  �c�� A����)��t�Vֈv�W~@9���]=����j>*�DQ���ڤ��� I(�������Y���ة��l������7}H����d���Ԫ���U�f ��M�'��*ьi� �neY�ޓ�n`�*)�"���b̊�?B%�"(�ز�`���;��yz��9�\���4 I+�%}[���.!�)�'9��H �f͛�%ɝ1r���3��6��v
imZL��'��ވ@�Ic�x{*v��������ٽ8� &@��Ȑ�".Ңo{�`]�n��-ħ����F<0���7U��3���_k�����'���ݼ�̷6�!d��dX ��~��-���g�@(4�l_o��Z���ʮ=qq�O;�c�������y���x�-"5D��`,�lN�1&��N����}�}�
��35��6�	�j� A���� s@�0F��PX2�wbd9��e�����<�=���Go<	���6B"�wo�ֱ�=���	&}`��A|�2JÂ�fZ��r]]S��ngƞ �7K�p,�1���̑���y%8��R�>��5��[a�1������5���P(Ҕ[���k��@��dT~�)���T��7��:P]2�	�#���6U�D�6?%X*d���.���G����V���OtC���J� �"o�,�}k(��s�h,�{�v�(E���*�2P]	��J��fMW�I{�]��pli��ʰA�!�~?I,X2/��PT>����g|��_ӫ=���'�o;8.~��8РG���lLys+%�4��&��X[�q���g1����R��7n�a[B�=�"N��>"�]{h�2���y�Wz��u�H3���9x��f����ݖ#TM
�K/��Ș�C�����o�����}"Nd#�F�qq�Y��gܲ_�U��R����U ��g�C�(�	���[hU��3��4+���$� �(Pأ�-�y���3���1���Tݽ
l��_P�D(�D�ř	�"&h˔1kٓ���r\��_���:��+;I�1[Z!�j� ##�9����
yݎ��B��?OJ��2P�?$��3����>X���̓K�l�;��fE@�aI���Շb�=H���ڤ�3y���s��g� �7���v=��Q��P?ou2 !D���x��<���}}���'�k;8C�5p#��́�����TMy/�<��*y�3��(r��Tge>�{j����Xt�u�ƃ�RY����W}*P9�j�Z�J�"�s���|��G��uei��9v���v7�
[j=wՂ3d.�Vn���K�ҝF��s�h����nHYim�]X:�m� ��G�ӽw���:�ZJ�Eb��v.L���G6��7.rE;8C��e�����	Ϙxޢ��7��e�W�#CxZ	t:�^m�U���oi�oq��!+\j�t;�vZچ��fk]���`�����+f'%�%�R����f�6�Z4�k���M��|5�.�
��ռ�3B���]���b���>*'>�0���v΄Z�V�.5z�ѧ���gF���-K�yԍ}�W0�e��&�Q�V۽�ۄ�n�~��5#��}L��w���/s�^RP��gV�DǸ�y*��������t�j̔ev�Ջ��)6�Sn��27uʴІ��e������)����E�
�\�݋:T7�x*�oZsz�;V{�S#�v�&-���hm���I݅�
�E�U;Z�L�1���Ru��ݔ�]�(]��Ɩ૘�+�f��U#tzf�PW-m)�Ra*�R%-�UKb��+45Ng�qpi�c�EJ�B�3��w-uc�7uJ���*;�ž��3Εpʪ{X�V&����<G��g"�ķѶb�B��P��"���}-��ݖ}��;�Sm�JBV��C�tׂ@���;�b�Ȣ����w�=��n��vY^ar�ڛ��'/����\Cۭ;��Om�E�QNW{sz��:+��k���e�lӬ�m^G���|�밻[tq_���8`�;���;(m|�(�VyVw=��������X�>�`��#������.�;�u���~Y���k��~�~�w�^W��_��ק]]e�ۊ�w�+���{h��ue�ͫ��$_��Ѷ�����_�j�8�
H"�2��rQ�n�����.�;���]���.��r.�Οn��{gGprW��t��ʿ>�N̒����˶�D��q�we��'���gQ$cnӎ;���m��k�����-��Ί�)�^z��)8I��;�����Y�SA۷�T]<��B[l0��+ɡ�)L��Kqe:��	L7�H훘K�k]P��bBV�`]���nH�v[nb�V��*ڤ�)Л+��х��ǳ�M)(l���팼;I�h��B��#�e�[�f%��pձ�%Pq�Z���F��f�j�1+J�˨Mv.U钥��"�v�F&��u�@�Ԥ���W9�p�3�x���l�ƙ�����I[�UȬ���_)u�g�4)bSKp	d]�uzmM��3E�5�N�Z�l,))YFUs�p@1�6]�t��`�ɶf���N5qt��WG��d�C,6B����-h�LK�C%������Z%��s����!�mWF����pf��8
���aؘu��Z��[�s����f�-f%��jc��BX�wM�����lYa��[í�����X�G2�HmT�,yb�ǜS,֌�ͱei	�M�Qb�F[HR�.�M�7\��2e���X2�h�4K�h���h�`E��Rh�nZm`[�lcocR`q�)�\::fkR�X.[+v���,�R�J<̶`%�֡16l�u�9n+�\�2�.k%M�f�m2�b&���ʙ�y�5͚CAѶ�� ��Ų{YG0I�[�WSs�ma��k(�J��FZnV�v�nI�g�Je8p��%�@z���j�U�<�hD.H���m0@҃C
V�CGS9��̮nc��vCRXh�*M��\��jร��|7�%�z�x��e��0�� l�${K�j�q64�U�&�X��k��3.�%e�Zk�UZ�Y�!�1��M6,d�m*���h�f̽�X�m�س*�9��hYB�R7[�u��E��d��qm��BͩbS�I��SkBmy�mL������i]�l2���E�Ur��Z��*�Q![X��`�S W	��d?�N�'u��1t%7�pM2K���rM��u�i�8r����� ��k�vL�ۭ��u��al֏d�t�Z�0&��v�\�*�i�#r1s��8f�#%cZ(�KP4��Dٺ�ٔ��iê��q�Wz��i�k�]��"԰#��1�q+B[\�6��U�����n� ���P�*
]d�X�s7��y������~��etP�q[,��I��!��h��-�CA�8r��w�?�	��$>�0�m�B/yb;���y�M/}2�ׂg<�,.u=��$�0ȅ2�@�{����ʲ��&��w�����n�Ӻ�a�,��^|�P��4�I(Y�Q��N�,L�����y��O�����
 �f* ��� �?>�M�]���i���7�+�!G�$�,.~�z�ӂ��i�K�A���q���3�����oa~:D$��dB� ���*�BW��yB�f��X��P����R��@a�<��{���29�aRUK�Q%+WJ�c�n��*g$c��YT&�.�lmQ�-+���ݓ|�πȨ�!ss�\��}�뱍����I�L���#�����B��~���V�UP�Et�����Ǝ�������ũ�c/+�rL����;��nb"N�CmbxQ��؟>֚[y�cF9wU������8}�N��<�>�q�u�ά�`��A2D@��$�GU}���l*^�1w��!;}B��|F�y�A��4������D�tN�»��p�)Ǹ�q������LM�w��Go=�����B4�ޗ�D����®xs>�u����N4+�C�f�M-�w|��Ր{hP"��W� �"7��.Q��	:ŇA�_-���)}�l�w�,Ⱦ��(�mon�z��~��qJ��K4"\@�aqUAˈ�h[��@m��{���J�(Q~��,j�sh�x�n�G��K� ��
i_��X�"�������k>mi��B\���ے�[t<q�D��|d��V�{�9�(e	��X"D X�XPZ�;ҏ�
���c�Ý�uՔr��F���S�j.��\g����CL�5��I����}�Iz���s#��,�F�X2*���D������w/q�;��$A��H̀���l��<i�a�|�1�X#�+�M�t���? ��_ŔA��W�6�_Œq';b!�
��SͿAw9�ܕ����Т	��%aIB�͎8��o��!��6�WM-�E��0GR����.2��,�����F[F%�߿� �ڟ�"������~��\��:��k�����
?!�/�̈QK�A�
"�ڣVU�i��~��/�V.����=
����e)#v���Ʌce��W:񜨂҈?I,Y�}@�iw捛���+�����v�]�m_���
?BrW�%
?D����e"y�j�@��̑:��Kk�g'wi{�����{i�uy�ȳ:�=s25�E�&Ú"�ERMk������c��C�#+6��Y��em�Z��.c��6�p�ab��� �>WC�� x��J�F���V�&���m��AA�9�/�T�����r�H ����?FfH�	�L��D<T���m#�i��l�;v��ݮ��-�YSP�.���W�Hg����Ȩ~0�����w�Σ펻 [~����g�j�q �/�ǻ�� �%
C���+�U�/p��o�qQ���?r����u���Q��� ^u�"�����ƈ�C>/P��1$�H��;|�ʂ�����ז﬍>W��@Cg�$���?3��Ww�p�A�,Y�_P0�.{�]�s��c��߬�
z�iʔ�j�Ao*�؀��?%_�%
"��~�:^�>���q���T.��X*;�2@y����~���
�7�����c��{��L`7�ı}�����!����������:�7�'v�_8�_<�������;�d[�q�NtsM2�m��e۔Vf����Gyc, tsH�,4�v�]������&e)��5�*(�-���j�ưK3f�V�q���Z֡U�9��E�H��E��;v��LP�,�V6]�*-�&$�5�\Kit�vj�(�^������[��Uq�	�) ���˩�R!��f��+��}��Y>a˩\� �T��-$��b�٘��qDD���%��s�N�E�t���Ț�\0�3m�D�Z�g�Γ�������ݡ@�W��%2* �!@��^O���=�ED<Tɼ�߯z��ev@��`�Є������4O��P?D��꿈2P��?I(3��)9Nη��?{��VvĘ�_{�d"�X����K���֓�օ�E�����$f@���f�GD�Z�g�.��:e����?lF�~>�`ȨL!~�X�dZ����WP@B��kW}��>���_<C��~FIV �gh�����a6�[+�Peԥ2[K+���˦3���F�pɕ(I�ĝ�z�wP@�0~9�!�/�9^���baR�"�m�Oul� ��X��*�!$��D(�g������Wž3�r�#��T-�/���C�_�a�u{�j�#3��E'�n5�������P�#|�t������k���ǃ`ͷ�営g� �z�#��k�_n̉/a	� �$��L�#9d�T~�mn����.z���kB� $��H�|D(�0��nU���@��2D����l.=�
��?! C��v]w�a~TA:E�$v9�D? d��g-��xC�}�"~h!�a�3y��ye���An�� �P�D )%�:S�6z�4��+��f�˒\-�0�K�r��J��(2h=��ե�,-�5��O����|&�N�����v��C�"���V���u�A����d����(�Q%Y�����^�#���/���M_��H`T����D�}b��	��������"�P���!@��_/����%}�_�^S�\�!sh�2z�k����m��˙�K�=�T�L×��̈�nc�ߵz�}��"�f׾ٜn�T.�T�}���P�s�l�d��@g��oiI=A���I/��+֣�@�-ذvB �!^l�T�n��m�jzA�����/���Ҁ��2J�A��
l7�r�/w`'�b�@�M�]g�B�R��d C��fE@�#3rͧ�=���[i֛gB&)�e�	ZRى���s���%r]��5l{7��� I+�%>��l���7����-r\A�4�?��,ȨA�"7��Wp��2h`���W�]<�
�wx�ƜB/�2J9���{��@i�	��d(P"~?I,hT�1���K5��kG�Â�x���!�P�"�~�	&X��2Q��f����d�X�n�N�zץ�ZCO�?>ʲ0\������%I�y."�3��ԭ��=���*�S�X�ٔ�_�戦�g�ğ�nf-N|`�#���K���C�~��>ᝃ��?޿�L��$�,Ȯc�gg�f3��@�}Z�u�\�6�5= �sP��*ȑ����p�:~�&urց4.�W��k�6[jy\�!@���k/,2\���	�ξ��+�!G�% ]~֢�����T�EM��-#A�X��Q���!'2 ����yb��{�|�/�>ATpt�on/��DxM�) ������ޢG|��ł�A���$�,�#��G�!���V>|%g�ΐm?}`��
 ���V"D?B7�������d�@���5"��1�఩xM�����:{u�$��ǣO����	&X Ȁ��FIS؈�����&R\h�tTs�wӶ�x	����Т!_���^��s(/U)M2��E�9!9����!��e��Ɖ{Z"�x�t�x����;N������+ْ��ݸf��1cvۨ/#�}��(�x�0$��4�!z�gJ�1��6L�2��oU�������1��RR�+6�1-����4�ۂB�t#t\h�Fde6p���,\t����YT��.�-�-��?�G���ԫ)է]�`De�mN�f  �\�Ef��Ba�!6�#[��w6&j5f�-��&�f���턇$lj��8m���~�����tc�Y�	S]�7^y"�E*Kh�a�ɬ)e~�yP�=���L�![��VO>��gH6���b�=5`��q|�� �%
B�&I_]�G9ڳS|��F�e$S�3��NK��d���Ȕ�r��g���b���!DC�I_X���S�s5W92*��5pwOg ���A���|D(�D���03k�����E�!���� �
ۮU�z1W����M8���n�<�T���5r��=�(
 �d�d(W�C|2(}��}Y,jE9��w��,*^ �g�'�X2/�;��֎��<��y����������P�+��nrt��D̲Ԩ��U1?e�D�1W���a�����N�����wҟ�1���>"Ib�2*�������t���VI�ƅ\��
���j��!�]͇ux2}i�ep��7�j�[��y�ܾ�v���.���"��j�gj�W��\�� r�;����Vk�/fn�y���k`"	�#$��N[����y|<�'�*�"D(���%��̹���]����6�o���T� �(d��"��
I,XNf,���A|��U�$A�ѻ�j�����3���R�q���@@b�o� �D��,ȵ�|ޓ���wgz��*z������<Т_ d�`�ُt���4�l]�Ub�$�YK����`P���fuڕ�cЬ�L�#�D�C���ۨ"0���~��F-��	>�*���&�C�"�g�Q�J�D#q����J�+��}B�wM�I�'\���x~;�����nT��Ͼ��[+髈'�@�%}"�����~q�;keDG��{is<�ue��|����E�.�xl�^.9ƛںVM)��=��șJ�3Aі�d�✥A��c9M�R�_Uhಘp�"H�:�*�O%�r�XF�wN5V�;���ؕnaI-_nYw��B2��
�Ff;m��l�AV��v����n��֒�����񂞴�ٖ-5vo%�rl�8����z)v(of8������k�C���Ճ�5h/�W��F"r��VЗ
T-vo�r�Cq���m7i@��%_u:�,�5�ٷw��--8Q�Uw�S���*�*b����7n�m1v��9tE#�r-F͝&L��
*ǘ{���Epo"}��̩���m��cqb�̋6��1�]Z�����;�s��j���ղ	Z����c���[�GuT��ܖ��M㊧M������M�֚U����=����p�4iPb�t�J��s�ŷ�A��R�З����1oQ��3U����Ø�`҄drf�-A��Tף��TB��s����*�SW��xznl���23HW°���L�0;L��㸗�p�R�D9���FR�[�'v��c�Oy�V��ͩ;*[纶�k.l9�EL���hi�|��ǜ)��}���Y&�r;_r�d\�i���F�h��]&՝8k/m�w;\,wW-슍>�4�[�f�+x&�0�Uh��Zj�[�TY�e���@#�ー����wq'ǝdD$U��w^tP�ͷY�Gtt�<���GE������ݗ�yaq��q�QZ�tv�����yo3�����]ï-�o��m�YgR_�e/�jVv��~Y��^]�y�Q�]�{�Ֆu�\_ͺ$�C����I��)%�Z���	
E�mA������_{vY��Yq�6��w�w�|�.����mv�m�:3�=&��������m~]�Q�_+:�C.�������N��4:!J����ʂ��^j��N�;/m���|��*
�N�!>Vrvu��E�Y=���.�#�Y^vE6诶����wft��ͻ�����g��(S���k��⴯+p����N���w��g?���}�V�n�{/:�n`�k�P?�#$�"D(�QG�;���q~�F�31��}��5�3"�Q�d�!�M_{�⼏z8��@�%�ȅL!%e�ʎ,nPip�ŵ,�u�pO���W|F�|2D}��b4[1Q��|��ߚU��X�;6\�Ƣ�u#�HSUK�nۨ����Z6��@�V]���(u�2*!U=��zt��ԝ �~4X�
±�����BA��� IB��/���J�x�x��
���}c�)��n�$��K�|E�A���W�T뱔@��/��(��#$�%|�6�Wβq38�Ʒ]'����Ғ�A��J�E���M1�|F�`�TA��j��]��9լ��_} ��s��n(2��R�R�q�{�wRϪ'��5,����/a*��$e��d��$�9	.���z!V�esS���x@�5L�_��-�����oti���Qe]� n��-E�~z\-�X��?/�zř����,�,f�a�,#�4!�&�2�SIv���.�ݘ`�����f�ia�9�@#�9���bR\̷0��u�X���ܴm�i�$�ۋVA�P"~"Ib̊�ЄF���^���B�@W��wens�Y{��8��~�f.��n�!O �c�=ؤ�
"��%�Rܮָ�����pڮ��T�A�D���L�a$��Ip��*vN�bA���8��"2�Y�̱<���$3��n��y �V����COܗ�M�`Ȩ�D(�%}"�.�E^]|�a�{k�ky�������Nr�����$C�-_���I0c���+G�p���˜q��y��f)KI��S���˨�w��r�N/cL�	���+(�󅚬7��Bwٺ�C�k挬t��͍q�.%���j�n+,&��nR�a)v�D�#��'e�b:M�Y�(��j����g�#^+���Ԉ�������pJl�C!� ��!f����b�A�lp�Re�. ���rK��]n��aideFf�6ajۜ
�lo1&ݱՐMM��]Hԫ����~�����)`m���E���g�\�ɓ:���K�����%��˾{d��b�#��B@��Ɵ���
n,B�"�&j��Td7�O�� a�3(H'2��W-=���<�}��B�0�tz�
a|�@&�) ��?g^�����6��Z"q�7�ف����M��[�fM�L\��;qǝ �����|�����(�[���l�,�}B�"�ń�M����9��T�"
E^�3��_!Ƕ>@"� X ȅ~���PuZ�}�p�oa�t��M6X���C��RF�¾?I(+��7+EnϾP�Q��(�B���,���æ;sc�����Gp˥�.���w�p�D��/��0�-��^w�I�q�����m��o�]u�#O�^��P�D(��U���n��:��LF敘J��E�ܻ�e'�D��"�e:N��֑Y_a�t�C6f�̨�\�m�YY��BGqZQ�2p�M~���\��t���m>�-zM7� �" l��EF�i@�	�ِ���$��� �d} �S�1܎�D�C�bV.ļ�z)��
�]��"0�fd��ȫ�/��kю���GD+�ڢ,�/3ѭw��c�lK��b�Š�Bi��ϴ��}shP"��U����ʉ�}\���-"69�����Sqa(���<�d"8G*�yXh�smP�5dS.�R�Y�6e���CJZ�nl7l��1b���?��d= fb��_T8���gn��v���dO:���V�;� G㙒'��8~L�9�i�[!��@�a
�O3�}�=Sd�m��
���Q��,�_��C�ҁ�ڲ$B�������d̲��^��_��q�P��꫹_�Fλ	y��X�R"C�:�]E�s��[�Z�Ց��[��|�qM{;��QL�G�?!F�X2*!�b'�퇨Qb���H���Y��~̛�-K�s�"w�t_n�H���%I����������Fv�zOT��羶�|����_V:�ܘA��6(]B�$+6�TV�D3���\�QC�`l1��A)H�(I�W`Kh=��������|�)�ew�#As� \� dRJ%��~ɛRؚ��M��+k�f��3�2��Rm�+�o|�y���w�J�A霯��T���)��:�>ǵ�����W�)��n�>�O��X�強q��"�E��L���� ��j"��Ҩk��]-��=v���Z��U'�XelK�9��2���*�G:ξ��3��!(/z�$������&��$������|ֹ�? ?~RJ/�RO��g�m-�|TdW{7Y=<��r*�� )�f�^��2f��V�j�ݪ�0����4�m��ˑ�Ba�Q���d�[A������������>��o��?}�;��^��m}�z��I ���F�A� �I@ߖ�oo�D�'U�Л�,^��N>+�����$�$��!��5oyߪ�&b���~�=�+��$@I*NC|�uj��,n�|���q�ϛ�o�u?|�/:���k��{���I$� ��rH���F������(�4��Bo�τ���ܧL��njwjTc�Z�Vx 9�`�4�#p�k����	^��ت�f������q�$�w����Q1�9��~�I:{|����h¥ظok!�M�([�5m�<�*����
V!5pB���F���-��n-lFhL�RԹƪ$b���☘�D�1��B͡�7�f�ʶ�:�7�m�J[&����KvAm҅)�L�kԍW"ZU3HBE�Ѯ�^ڸ3�Y^����3��+rK--ZM365��)�X�fҮU��2��?>��JèJ8w:�[��ń!�6�5�]-Dyѵ\��kO�I(	�n��/R鹾U\MZ�Rq�=M��b���C2> ���pr�:<^ =�n=t��;��}��x<_�I}�����.���/{Wّ��̤7Mt�x��<�����Z��xU���W�/�_I(e�^�Y��ϻ����1KԽ/}�.��I�sڇ�8��V���	�!$���V4_��b��6�N�o�d��� tRJ��8.+>�[��7�����p��B���.�ۿ^)|<E�/lh&�s���?K���2~��v/\��ye-��zC��mm��$�W�/f��2v%��w�ߩ��^0�Fb���?gs�y6=����`�V���[v���y�&A�L�����-�����b����z���lm6�Md���~�S5�fR��e�8�y8<{=3�t;��$��K����T��U���s�S����T�X�P�%��|��jI(�^͵�~�L��u^hQ������_	�H����\�砖������g%�����yy��=�"�!|r��Am]
�<,�ɀl�7qr�%�.��R�Ss�ظ���_Oܟ^����9ofz�q�Ы�?}�#�j�卋��$R!$�������m�gDΥ�e���Z�1�|�.6�"�V��-�|:!"I_}$/<v��yA�Zw~��'�O��wB����.��# ��6拷Y��uv���o�.��s�����O���v�荷D���W/?=��H��W�!���p=���"���:����W�u? �w�4^�lR����/�%}"N�����)��Сij�q�{*V���`}�C�����_����<�5V�S��XY�[���]]tS���&�Yuy�g��d��͚�iw���^{�+�(m����t_I$�v�y���������g�oz%}'S�Η$��Wua�]]�{	:��H��+���ELD�U���5;�L��"H�������&bW�v}ھoh�v���K�ݵr��`{��]c��)y^Y�t�����*v�Y��,��L٪��6���7c=�����"%-
�F�D�u�ݾ�I�3�Z�j>  ;��|��2>̏�33�3栍_��'��_vDN�j���܁�����_z������4��!��X̎tu1eƌ�c3cZi��9ĸ�U2�	3.w��{�#3��	���-��j\��ٛ��v"Iz��������t�C2�[�U�1˷a�Mv] �!��Ӽ���X-�>��`�} ^U��a��F����/�
���=��:!$��H��牫�����ߧ��I@�]�f��X�g��ۺSL{W�ἤ�"�I' }�GƋ������ዷ��d����"�I�O,�5o/|��K=1w�1v�Aq�[��.�����͑�5}��������U��E��ԃ5�	�����#��u��w.
\�̼�آ�R�sWƲ��g6.�vQ3�1�3�#�6�,���^�:I�;E�[�I�#v�*�up�eسkn�s������r�q_Q�IrYY��2F�[VZ�Ә�	f7/d��f��� TV|�u�S�&�p�wշpwPS1(q�XJ�L8���2���Wq�Z^����x��O��D}{�"�BoNJ��IRm<7���tM�B�j`41j׉��fP��B�6Wk�Nĭ%�.J��RE����#�q�*���w*G�7�:��rN�gn��ˎ\#�ty�ī�i��3��V�̦74�XeZ��������YM�m���y>�3�^�Y���G\�U!:�
h�;;�c=�����1ۇ�}]�0l��v3
����wUֽ:�9����]R]ʮlVS���i�����]�^�ޣ�N���F���VI�m��ݝ[B��[zxq�u8��+n��+ܧ���2�x]7"�3!�.��M7�W8��I�R$J��h��js2���9u;#uLj��:&�;f+�$+a�g���'�M:Ɉ��
�+9S��m9aɈ,V�E�B��y�v�ط��z��T,����ڎ�wn�ౘ@J�MS�����9ڜAWLq��"��@N�.�*������wM�]��-ˈ:6��ِ]�r�j�����?���^vV؊�(��⸨���:�#�2���K;3�����w�uI܋n��u�ERs�IyqY��n��"8�;�E������O�[�쒊.;�(�:�8:8��igy��yw�ܣ�:�=����D�E	�G]�G_�bqgu�?7y�ܾ�וC�ȏ/{H�,W�w˾�TT����Ȥ�;��L��:������N�y�W�Z���⢉;�W�o�>ێo�qzQ�Yq$�]'�.�;��f�.����}����YB�e��nJ��[����[Kl�ZCf���գ%��+�;�#��FArce��@B�(U���cAh��1������ˍn�9��JY��Z����G4��4ô�UKq��iR�%Gk4�+�����o;��eɳ12k4��c6�:��T\�2�R<��7Q��f��MM�l2�p����A�)m�ͩ��h�JTt��l2�hh��9tQ!%[��)cƔ��� �̺�fXn`�
���]��rؽ�5	VG0�R�f�ڰ6��c]uPP��Ō�l�7m���ʋ,J�!	���h+��f���k3�yd�Ŏ�뮬�)&�-PJ� �\a���l�GfWV4	\�l-R�D׷l�L;T����U���@j�f�,���\���<���]�η)�e�K�=WJ�&΋���hVTD�4%��"�ũu�ټ0�.
]�k���G`�&[��4����h$e�T���\���kq䶕u����{h����.X�]s���x�R7h�ݵtF��a
�6hB�m�h�6�pr���ŷ�m]�7CJ�R��mwY[f�� �$]�.��ͣ��TBb��cq�����d�@դ��-�*Z��Tn+�+� ��e%IR ��W#�IXݳ�\��qF�N��khܔ\aZ��Y�����m���%�LDΪ��Wd�S�5uv�\&����,#I�#�R�8(�,�0��q)���v���YjKڦ�;]aa0GK�]��i��d���Gm"�(�� �9����cs4���$�SܘC��B�q����+�v������M2�XL��6��.5��k--0p�,�n
�L���1CF`e�,ẍ́U�x��n�u�&�Uj���*��Я0���+�ط8�]*9�c7�t�<�;˲�L)F7:\
2m�D��ܚl���M1��Ԯ�Ѕ!Q�Į=y(���3]�Bی�(͓XR�KL��WP�j�d�d��9�oP�f,b9�J�3�G5..ԹQ��f�f!�p���qh�,BgF`��f�əI�K�0�%6��b�b�e�1�*�-�mhXZ]fXr�Ã/�����̥�.e�6�Mg��2�y�ي�̭�_Y�TEZ�H"��g�. 3���G+<�^>�*�N��w������]Ҥ���M��΅�;�E��]��}��}�T�1Z���Cb�E$�&�TT޿P��Ж�����d���}%�$Ϸ�
Y�ݍ�'-��V�>�*�N��x����=��u�S�$�H���綽���:�E�r��h����}&Iw����e�6��HE��Q��@��(3X����hLaҍ!iUf�@ڱ`ݻ�5��E$��_'�J�;����d�"�/sf��)��')%	��w���ӆ�ݚuK3KYAά����W��צy��[�2�sU�:,G��Ә��v6�QQ".��ܢ�ҥ~��m�{�z�����D��ug�x�E$����[��[/�ݠ$BE�����c6�^C���>��lv}v���"J�~����b�ވw�����5hPg��������(WL��wcڀ�&�k��C��S�U��m�?z%����V!�6�r���z���}��)��"֖�[c��j@.��5�fm�4\D]t��{��C�6�Y?�/lWQ���M�k�^���ͯ�R���p�+Jz�X�`���{|;K~��=�7�=r��nk�P�_}�6�A�V�v�dPR:y�L��Y�~z7f�Kݝ�&�
��E�A�����ze,{��\����s�����Ui�e� ��W���K;_W�b���o��eir�v�@�3���N���f��L�9]���/�/��h|��ٮ��^v%h�����qv�v<��>o���ue�9^���Bh1dP���H+��宲�����NH����[��*���uWw^��Z�@e<��o�jY������\�`���m�ͥ�9���v�}t�z=���K<����[���r��g^cT��/�C���m|ڡ�<�+�ٕ�^��
�Û�o��=���k�h[�(_z����K�of��o���s���V����ut+���g��a��i9cg��ė`�x��5��#yv[�Y�nG��^Ѽ�����{TZ���k�~�����/���6�m���/�Z�k��O>��:#���qm ��a�^^p8L��THUVJ4�)0�4fX�I�:����UYJ�ڠ�T�Ȼ��rm��M���w���y-�4|�N���N�Q����6�i���ߔ���<`s��MS1���;^׆Z�s�;G8ǵ�obhg��������:��;�YU~����n^���5�]�&���6�A�{�[��Ay�`6�m������β[�h�R�X�����m|���߻���\���m�~�{^׾���͡�~����r��w=�QB׫��ط��}�����j�ٷLE��Wvv����d4Wk���Cv��vE�9a�ޤ�nhK�#���;�O_[�&8ޱ28Xˤ�7Uc�a��ֶ�$�nҬv+���[lH3\�����Ω�F��4K��m"Ut�v��΂�n����Vgq����Mu�����Y\�.&kh3c�����)s�����.k��A0E��ma�6[��P�m���]h�cQ�e�	�XM��MT�u�˭�9QZ͗�����Ú�R�6�@�5.���
K��,���Ҵ(����b���m}�;/����f��xx���]��e�g����ͦ�*��{���{c7���уχ�J�o�6���l��p��NC��m��d><�s�5O�̌����k���n�.��u�g_�v%�\]�|����pyW��y]�۬/���m�r��6�m �b�y�p~������o��J�o�6��&�n\~��;�/v�7wd'kV���(�]l֌*��r�r�^����-����}�q����}��T�Y�ꮺ�I�mpN���н4�i�ޖ���\4j{�����Nw�.	����4�mD[��̈�|w6�Y���U75^N��W'�b�b ��� :�.�����������h�>h��묩�]ד���6�k������C��
��+%��C�r����7h�a��GW�f�M����nj���w��W���o:K�ι���6�mۺ��j��!W6��4Wa�f��}v�ț@7L�^<Y@߆�$��,�7pM�j7,;(�ɃYv�!�.�a�M�5�ݿ�P�i�߰�s���J�s�����gz�o�{4A�A�^oI���gc���-���g�����o�g�(y�yg�����߼�yJY@��ykNtDb�K�V���b��ȋ�Y�*��XM]'B_)����܂(���T�[	;1��g|>o9<��v�*h�?��F���m�0��sső|��`�L]\<:V;�m|RY�e���f������D{7I�����۶��:��r����ͦ��z�a������ļg�6�Cd��0���%22/�h>yLa.���J��J�7U��C����h��~��}��r�#��!����=�z}W���v]����,z�}�}5�x�gr>+�|_w �=}����k��#B4k��j�w��>_��9�t�õ��¢�m�A�X9�B���p����6�|��������9�0U��8�2e�Yޯ{�Pk��]k�cI�@����QQϮ_��;ic_<�t!���oL솘�r�_]�-�T��� }���}��@6�m�e������v�h����2�d�m����ӾD�=���M���vv*�1k]ZrLH!6�x�)��V��B�uUwN|&/4��yW�Z����.
�pB�ȗ���n@6�X�\WMͬ���kBE���Y�>�s#��ƀmg��gME��S~������۰��^�I�Ǻ�3܏q�Ǔ��;�m۳MT8k9��, �In��?y)]�W��_7R��7����l�S5��N��+�gt����y}��4�6|��#�P5��d�T�}M��X.��@ʝ��U�}f�l�Y���VP����/�G���	U�������n$��|�0 �3�6�[���(��1�R�H�a���[�.������R��c���+3PsF�V�,��`5Du
�X���b��9��] &�c���]�v�G�t�c(�
���[�&�M.�`A��b�IiQ��%m[�֘ԮDu��&7.�m��͆V��o%H7.���T�m�>�=��W��Lk��keҚ4�����`sbWJ
�]Z�UՃ��Uh]�� �!?7�s�!���{K�������(aG�۳��]��qK���˞t;�s�yQ��Z��Z�W��\�ӷw�{���xؗ�����ߓ�l���]��*L���km��ߥ+ɯ�����vm��W�ez��v���nC1RN���:�\�_6����%���4�s��n�Otz��n�@����-�Xޒ��aD��~P��NqJR�n��+�V�ʛX���t�������؀��_7�v�R��䤼]Gڱ;�bR��}Z��n��h�&z���V:�E6]i�e�T�m+�{خbn�
:F�s����fUڦ�.�c\��� ����ŒEHyg\��qb�������j�S�ԗ������sq���{��j|�����s�`h[gR�Y�i�]�����3(fS�75�Z<yw�Z����؋ɥ��v�.�����^�{�556�h6�	��-��ȊJ_�TU�Y<�Y�]�jx��@6�yv�����g��V���]�&��xr���t�Ó-���X2��Bb�����{��Q�y�Scu��V��^�l�ت\�-� m6�l�ޞ�+ͿJ�=���!��*Y*����.���C[}}�?_&�m ۗ�5���-��wP��Z�P�y!B������
�*�=�k��f��L=X/6uV}�B�<�r)��u�m��ɜ�ˮUb�ꐳ���\:V�Fj�
����Ӯ�L����d��2���W�&�f�e[�zę����Wγ�:�E	�*��
s;�i�}�Whw�j��\�K�yP>:wջ-�äU�έ�f��wd=�J��]+ͽ�}9���{����|�4�YW�N�
�V�Q��k˹NQ��8��Z�AY-oJ�E����A�y�XE:mlf�����ZjuΠ�/��ҵ���F��SIk8���7��A�AUt�R�u���Ѫ��,��T�V+�����v,I�j�x9
���on�5 W)趖&BxFu���*rL�3�Z'���Y�����wN��[.�N0�-�Kj�����Q��:�f�+�R����	S��W���I���Zݺ�wHv�(bI��X����fY�k��%E��<�!*oq%y��YW����gK#S��xH�_n�nC7�Cb��S]������;ur�a��Ŕ������S)�[Q��s����P�G%DMLC4���j��@��Cq��soag!�K3��V�ֈ3n��=���� ʂ���
��z�zz��=ȓ�v;؆�}�vT����޻�Dw���;���\%0���B�b`e8t�h�2��5���߃��B���,)�֤w^v�G��U��x����޺�/_��y�����u_,m�l�ʰ��p.;�(�/6םGVS��(��3�/N��:8�ί*�{Y�ǝ�՞֞�7��yw������on��"�+:;��u��Y$y�\s�}�ٝy��t۹;2��Ee�w��J���[���y=���;��wyx�qE��u�ۯ/3o{���N,�:oz��;��Ns��&�YsZ�:�8��H����ēP��N�ä�Y&���N��.ʰ�+#����$�� 	��'&ި��ۺ�P�]��b�꾺�e�܃hd��z�����{^�V��0ޣ�u�<ռ�i�n��͵�&e��������)��Z�}u�i���U�k�̟%T��UW�����M]�żsU�Z�Ը͘X��?�>z�����ޞ���r�Wr�Ot�O�95���C��mЯ*֕9�<@dY��cT�����mw���qw5{M�t.�P�6�m��^���z�Dɔ���ԻΣ�!�6�m�7����¾�C��v��w�y�V�7[�kK�Z�!5:�±IE`��<���։{T[�m�,�ig-��ƫ��s'�2�>^���U��_˙#qnmjq��>����r�m����-��)��iC?f:����4��'m��������$���(��F�i�j7]oW����G��ì��QfE��gQ���y��M�B3���w�ܫ��>fnPEU�m����6J�ޛ2�kt�v��O4�����x��ooj��8;�u��C��V�_E�~�%vu���ok�V��4����N�W ����`6��ϯ������w�G�0��Q�7d���6�_������7���F�ے��]�Z]��]��rm���Sŷ��� 0��TV�if��8�97�!/D��r��g�t�&�sΪ��H�2�+�]�cX��0Nd{�����eJ$%8O�v�A�t!kWk�*�,Ě�T혖�c3�k,q
���5���&� ���֌%���s(K�ז鉨&h����u�vza��a��k�ֺ�^mm�-Be���(�+�ԛ76�[���EAj6�^2M2�*V���kn�@��Ƭ1���3^�f0�s
��iX�gm�M�M�{��~��6�b]�+��tƔHޢu��nvx�#3w6&v��~w�/�W��md�ځ{��3���x}���$D2� �_>_|�m|�"^ڗ�������
{��,e�u|�dM�6簘�&������A�z
��m�n����f���]�����ͷcm�:U��};޿�h}NpGn�p�w��L0��^N�H��C�6�i���))�޺Q��0�{}2�es7�m|2&����>T=<I�^�,ݱ4n��.	R���"k.��1��cA�(�i�"�9�����W���gE��Z��[o�Q���:������BH �p;�r�����U����f-]�t�Ì�	�_L���:z+��4�rCr8]p��h�n�L{Ṣ�>�{r\��L��<��W�����g;Ҵn����	jr��ǵ�1UfE/�,�aG���W;^x�ț_6�m�^�t{�7/D�=�m7oƫ�t�]Ox���ʻ �l�X�m���[����|K�ny�
��g9���+P�_7��X5���������[�#4 �f��LjJ��b�)�hlC`���������[���u���젮���ʺ��h�^f��M_۰��C��Te7S�W�t;*�mLmO}�.�W��iඕ�z�Y��i����1|�V��ɐKj֓���{����O�'��~s�}�Z<�n�Ub��ҖwMү�m��|��npXg^Bp�����r��8{s��j�sn�m�ƛ�Kn55և[�d�?e�u�����x\�3+�n ��m|�婜�I]��Ў�j��?Y�����ھ����Yq�8�K�����~�
R�k�c3���ܔڒ��A]4 hS]q���ԛ��};ף�z�x�ql:��kom�#�$���Wö���vC{��vM�|��5�S|�v���>�"o�����,�`�_T_8�m���zf�.�9��g�����i�@�t3�R�ݔ��_�۷Jz,�콧�W�����Ю�tO��:C�O���,��i.X̲,�>��W3=͵3d���%L��2(�d�`h�+zb{�4�*�]���O����m;���>HEA�ݡ���}3V:=o%�����]��ۦ7��TRݣwErc3pX���1�%�e)��y��d�-e���o�ݓϻ=z�7�������g�쾯}�^���E-�l[ɶ�6����]wwxng5�����^�>z�>���A��gz�s�W�U�ù�m7Nn�˯:岽ٽf�T�>��K��v$v*�N�4y�Η�x��^wC�J�^���8)Y�{dVG�&���f���J����77ֲ��������
k᜾m|ܔ���yj�����^j�cݜ0L8u�(�-a+�ָ=�{�Uq�`�_��z���ft��^��V�t;&����Q�i!jϤMI@,��-��޷E�����f�8�2�A�R`��Fۃ;:�hŬ]4R��alD���%���U҄�(�],f���-n�#������cq��;J�j��:�F�hB&v]H٫�X����%�ݗE�Qj�uj�2M��?Ǚ�5�B�BV�tl؍J�5BR69��!�l3�ڣ�n������T5(�[���-���=e�0O������U�iY��G%Ͻ�O?O�\}w�0Z���u�&BX��![�7�/�9o A�>mV��-��؀|���^�<�<�}w��3��y������>Ƿ�i����+�'bu�÷.�=^���m|�w��S�o���0>Ώ����#%���X���Q��5,�u{y��+�u�v����Ӻ�^�[���@\��n��g����C�j��r��)���9�d]�B�u*�f�kJsS��E��]���Fԋ��>���	>z'�GOW��w�ѝS�m�}�W1�ҭJ���m����ޠ�W8��T=f���I9v���ê���4��L�X�7���ѽQ����[���e�r�.�[OB��;i��Y��3q]���b8��5��){��(UN��ő7�Bb��U_f����۰ܽ���q����Ql��b����w��	��h6�nm��t¢�x�o~mg�5��g��L�z��Z��J�a�������_�o��b�d�t�+��;��PU8g�m}�w"�F�������%H+�L"�����ɍ4F�3)�]�f\m5r����Y2�Y��پ��������{�ub�e���};-w:��y��������T/g?����k=�׺��\�{-tM�q���,���j��w�/-���(gZxɫ�-He)�/FV��T�)�|)�f��G��ȁ��|�����ۜS�˱��t�L�Н+������]�#'w����+�hdn�m6��W�
�=�¢�m��ݍ��-���U T#�4n�����@6�_6�~��V��߮x<k�^�=�+���}�6�J��9��pWW��|U�x4�Z�J����M[��U7)p̀��:ՎKK���|��jm|]�:S�޲���<�|���D�@;���͠�/,�v��}S �C,���X���u��f!�A�:��m�����Z�u�i��n]X��Yw�65��=�랯V :&��:��Z�*U�v �s�����t:�
��>m[�¨��^BP]���U�rh���o���q9�YEu�9p�DUB��WU�z;�L��V:0�U�Y�~]�|��O�c�q������ʹ"Q]���#��im��V�fcxUGÜ]���/���'��׀����Q,�I�KŮh�QV����V�*�]�+�ե�Wy~���5�6�xn9p�~����Cr����gf=|�ͷc��ً��|]j��z�}��*�s���hdA�'�=w[W��G�cZ�6�m���ei[��}���]-����1jm�l��WbY���43��.r�n�vj�Zɢt�}�;mKBr��M����m
�m��&������(L�����}�U�^�WT%!h���S7�pg:%����fԭ�7Z{�Yn���YF�i�Tyf</��$&�fp��pT�"����ɶ�+{���dz�ԗ�*b7u���&��G8�P�z~�0RiC�R�Y�����wK.��.�ZZބ_
k;��ӭШ����Pj�h��sf�X�T9��f��!��T���#�M�A��Jr��e�Ve_1���;P�sD-�y�h(�벍�W�c�v���,X��p�ڰ��(P�M)��^��SVG.�ټ�I����{l�.��rc��2��l$��})ʧJ�2��gE�$.��������ϖ]v]1v���f���oN��P�E!�2�٨��Ħ�Ӄ5.vn�6�l�pvd��6w�ת�RR�v�*�J<��v��\�Ȟ3����d_[۪�)��m����:
d���Sk���t�<��HUܢ�e��������5sy���f�ഭY8�ee��rĩ��5/�[L^�ͪ��w����l�%��}�7F,U\��jR�S��(������D]�!�q�h�û�LŻ���2�'�v�|YJ�d֥�in�":�a駤�0��v�t�'6�c�˘m۳G��Y������Y�����ֈ��͙X����T(˩P)UH�2H���d��`��rS��V��!,Tg�rۚ���ce��ި�hihc�2��6ꑍ�$ĩ�9-5�fqf���T�@ɥ�1كw�=TOؑIKR�\	��`|�ɵe�9Sk/:�q�y���#���.�Wy_{]�.:�۲�.�mSn�㶷HEW������e���W��[��Sj�;��A����Ό��+#�;�;���xi��;�*�l��̞݇zi'm�:3n�s��o��7Yem�[q�n��1}��.5�Gaz�����9.���3�*�|�Z��;.�܈�m��diMj"�w�q�I�ܤH����;�K 쵷ݭ�\u��䕖w��������O��e�#�.�b���h��ËQݪ�W��as
��6���mjg��в���f�H�������P��fל��`!�Į��<[v4�4ڮ��؍�yP�KMURL̜�imѬh԰��Vn��y��5�;�!Q�u��)u�-MBk�	tt7Cc��%�8؃IE�k[!
�4j�ׂ7qK�\���$Â�ڳDai��]c�civ9v�p�̶8�e�L��p�h�t1��]����EH��`ؑf����8V4�MR�k��˅��6��e
�`������9�\�5�kh���gB�[dSh�z�� ��0�J�:˝)P^on{"�!se��&���a�5K�Ф���d.�iFˋ�Zb%"��۩���\b:ev%#Ir�[���2;�w\٭ЄYuTK�Vl�˜�l�4�f��Φ0�fй�QK�i�	�1���$ѕ)��M�
G��E��ԔBglX٬#,�L�1��1.��ól��]�la��WRPf��k5�E�^,�R�VT�b�nfC�~��ig�Z63X�v�n�f!Wb!#�]6�ڗ-�1Y*��u��r�R�^���1�i�sx����,�mQ%�bc�3@�-�ahZ�����,��8����.��Ƶ8�l��M�l��RT15�\�]�p���- �hh�k�M�����h@�Y�L�)%��h�A�fu]�sP�ň�r2�x�b�J�\H��%\�[��ELKj0K5���9�'hɀKe��ҘtR`�d���U^�t���MQQ�e�9�\f��!*�P���e�����Y��n��[e��0D:�Џ�yg�O%V��9ԭ̺ 4�d����3hK�rKn�WPGb�*�	c��jL�a�i��\:�
��V�vWlgf���h�*0���T�3+����;�5���k,e<&ơy�K�4����J�Ð J���s��Z�%z٨ֵ���9��1A�-��+t!���^Vmu��.��.��f�U�.�0-p��GE3)�8z��E�f+��(ѥ��7\�ns��xw.�bhm���5�����c+��'�%<K�m���+�����hhh�рb�U1\��ߟ?B@����F��]":aYhhm�]f�4�BHJD�W?��m݁wvk�>���ǖz��jۮ�㏻{&M��m�B�ؑb^��9�q�g+3N��+i�}V��b�G�7��y��c_۰1\��^���㯵Oz�
��}x�Si�G�OI�uJ}��a�1���z�=v��f_��y��7<��96��h7�������,��{L��ҕ��׫�U��Di�Cvx�?Z.пzl���.��5�!��c�?�O9Ԕ񺥫+��c�n�����6�Q���~޺�#=�üĐvK��~S��������z����w��!�`��Gg5�LZ�V�b�z-e[�N5D�+ܾ�K]��dT�nmHɬ¶���Gm�
C���2��.�ߺ����ṱ�����T�rvW.����M�uJg��ww��K<����V�|�M�׋���U]�G�~ֵ��_3���ׄ��v}�Z���W{������ٜ��A�ܙu����P�f*��]�������画�p-����)���~K���6(�%��)F 'a@F���jE]�B�]!UuE]ט�Z�6����`�l��ĺ�z�sָ����n�͠A�5�h;�:�����־�>��S�=�h��<��S��s��E�.�⬝X�����Z���kv(���������˦.z�md�	���<{��;��]̬9��s%�<A�(�vZ����m�Z���zu�49���Y|;��gMJ�UgKh�hH+�oS2����/�y�tG��+�ĺ�{�ju�Ȏ�s�z��m�m6���QM�j��!s�Sy_�,u^���oo�z����*0�4��sP*�4fv��u ��z�8]��n�f��������f��3�+��qˮ��ͩ[8)M����4M��_ya�>�F�qgv��W�,�:�{�9��ط��u�1�Kq}�M���^�n�Y{�k�=��j�LX �>���_|�ӷW�VҔ?>��ϛl6.�i���G���w�gq�7�̉5�cz�V� Yt�����ӯ��K���؎M6�᯳,�횥�S��d:ԣ�����>_�WD_�m�����������B���x[|��Zۿ��6�{/3����˷����ĳe�v�"V&1ɂ�iv��jb�b�+tJ7y|=�NM����Vwmg��G�k=�1���𧻓�&�͠�Ȭc��ʱ"�v|=�p�L���ً�jod��ïz���	�w �w�}���,�u�z�N�ϑc������6�m7�ʯW�z*\��k�M��V��=��½VG�W�ׯ}��܃k���η�=�i��f
��wxz^g`w]ᘀ�&�׼*��3��3��}N�/L��*�6�����u8ܧV�.�ے
��7�2���XW��!��휖D����.A἖�|?�z� A-v)��`������j��YF�.��ݣA&�\���ۉq�:����)�E��qD�楤MkM����b�ة2�{W0�R$�5s�F�!��ͦL���:jڶ��0�5�3(�aR��F���I
f&�]T�C��5��T.���f�K.�&�,	],e��u����X�LYI�������T�,�ْXf��[���ɑB̺
��4\�l���U�U�o�<��h|��n�SO[]�X���u��[�"IϽ�6݀��"�5�`m�Nom�=�=	�½V��[��A�Y؃�/�m���*��.��CwQ~��y�:����܀m|�n����;�}�������[[����U�[ԻOz�Ve$�=���m ��{.��Fv{t�[��/����Y���Q^�Ι�����E�����9�lvj®�v�g	.J6���J�u���\�h��[^�x�y͚���=���u�����m ���~�vJ�j��_[�$c��3����v�-J�R�s2e���w��ګ"e��^�\��u�t���}��}�:��q�r}^����3��V������v}��9��i�\��~���}�Z�56���NYm`2���Z�q��aK[��xι1�����xz��V-y�רk@6ݶ�k�n4d$�J��F��}�&��]��6��������D�D��$�*���ƈF��b����<����Z�.]����'�g�m|C�z+��z��A��y�K���Ɇ��_Ջ�6�m ��^Z3�Z���Ʃ=���\�U�{ª>}��+�:��[p���OSm���W��xy�m�_h���e�̝arDͺa�L74�,�̶���V.�Y�a�����ַL��;"콤�Ïe.�Ƌ���'?	��Kì�����1��܁v�IP��ݕ��>mN�~�=�~�pp^�@/fNT)����j�ͯ�M�`����MFG(��uWGmown�+��j>�A�~�GOk���8`�Z�6.��5��D�PlÝ�QYv*�Y�Ƹ��M�>����Zz�OW|�qLp��1��থC��!ŵ��y����|y�}j�}s�\ho�۱�8v]���
����w��V�HNC\�� 3#��y2�q��"���}��Յ���	��A�2 ���Ă�u��~�=��`����B����;��=�1��t��c�>���*�72����_�o[�e���w��t���w#*��]�]IR:���id8�ũڴYbo]uB�}�������dU��ED$��\?Z�ܓ����n��z{��C|&=��@Df�ّ_Fb�����v�G�P�����׌F�c�\aap�b�+HdUoa6"����,������Y����!�������mܻ����Gi��%�W��0|w�~2/��_H��9������@�|A�A}�{�b�xy߂��:| �Bs���s���5|�B1}�A:�|AmȐ[�%��]s�r(O(�A=��5n{�C|6�5p��X ��!��Ƚ��T�?]��P=��/��h��^�xm�n�{:>�5��?uP��nr�z�À4���!�"A �Ch mR��3���}ú��S�[9����ڟ�#���_6�Qs��ﺯ�7=76�UOHQ1,�jW>���Ϊ����	S˝*+Tc�����j�h%.T>��l����[o�{�;�c�� �*���L��T���*�Q0��mKi(��:B���#��pZZGGpS$�H��QJ�1na6
�[���Y0�(���Z!i��T��*[�l����v8�2�em����*d���bՉ&���ă1?{��[�逼.c4�%�nL�آ]5\Qu�n�q;Z���MW64�UO�y�����˯����Y�4�7u�t�eK��s��\$&4����������������}�����y�l�,����"�{����zjv�_�) ��6��mI
�fܩ��7@�a|svD�h���߼6��Ώ|A� A���g����q򏽛r/��ڒhGzG�]���V^d>����9��| �R<�D7 ۑ%�@��2�]�gD}�f9��>�� ߳�W���W�H��C���@�,.�o�Zڮ���]�$ �!�mI�!��'ax�L��ǐ���W����V���\}��"~-� ��)�!yp��|��B3͙ l�&uR�쭭��PVk��e��ɓf5���f��A�R?6���;h�^|!�p���k�Q���W[��t~���"@-���uU��dI�=2���梡��&�N�W0آ�e�z�L޺��*`�ԏf"j�a�^3���u��{	�:+������5W���}Ё��	���~ڮɯ#|6)�~z�-�V�u�F�K/���� �����W���Ch/�nF^�z�{���,[��}�չ�z�<հ�8�"Kp���!�2ٿH��3v 栁�k�m����k���g�O�&���G�lBq!y��f����͟����[s�p���P��wlq��o��E=�dς��+�Ʈ {�mI�a�+�/�#�Ͽ�Y�1��B�4��f�ֆo7v7]��K���"���Z2�p7�RA�!��-��Ng??}[��G�����/�ܹ�kфw�	\ ~n��Kp/U*�o�[����� ��磶�.=������@��RA�D7�]��h�R� �!	��r$�"	n 	����]Fj�ཱུd��{N	��ި.�w�2ǻvjث6\���4p\�>U�x�����ҺtI��KW\�k���B�\q��[��uJ�M�tw>�:��+��˛	n��	XM�]1[��P��IF��Q�ך����;$� �`R�������<Wu�jx*�q�Ki��hV�u�D�u#K&�(6!��qK�Rwsw)[�S]b7����s1i��2�M��ne���\�z���x 4�2�kӺ�N�鏅Ŵu��ؑE�xݹEnX�`{w�p:ubu�n�;{E�:-㩛�s:b�;558�P�n�~��;�yjF�ǵw[���U��L�)�j\%Wp���D�ON��r�a�R]mj71T;Vk�WvK�t�[�We6gi�)�nU�v���0�_�f�Vڶ�Z(�ZT+/i��Uvj2X�W�ɀ��n6_l�w���Y�����C5AS��a�h蒥���,GS���1�!.M�p�U���q{�Fkh��J��2 �s6�Ym�M�zd9�$n�T��ܘ�M�&TC9��	K�[��#���J�i!L�rgj�@�H�=�U�ιU��
��;���f~�ɒ+u���6�
dR�[3���pkkzJ�{؛�n�)���e���W8��
ٛӝ��r����,v�9h[���VXR���5<t.�eA�g-&-,�g2j��=E��OAt�K�ȉX!���vn���L��%������Q�n��e�Z�;�\Q�n$\jm��v\E3���nʯ��Ma9N�{Y���߽���E�[`K彻B���mZq�{��gYͩ�ec[��{g�-�Yvtv\�۳�"�2܌�:���u�E�M��ٛk&��ّ�����9��Sc,�����n2��n,X[��nZrC&�v��-���}�ֵ�~�/w�e������Zu�IY���Q-�ț\m��c�w$q ���[4Fe��+n��7<Ž�=1��EIW��*�%9�����$�3�|�=�����bc��j� !��ԐCh/�m=vO�3j}��_[��� �!�#�M�y�?}[��GuǏհ��=��Aѷ�ƞ�Dsas ��Am�m���3�S�/Q�1��ڬGxs)�p����S� ���6�ŷ"�]�d�D���C�.�B�a�kC]6	tZ52���!�>a��.̒"f��Q�~�����"Kp�?���?Wd��&7����ܤ=U{�,��b�y�A��E��/KjW�����K���Ȑ������﮵�����l /�"~-Ƶٹzƃ����}�-��-��p��s�U��Z&�P�*�,c�O/�O� �Z�3��|[r'��"5u���e���u9��,~-�y��*~���LLo���wOO^��3R��cǌͬb��dCW:����[�]ڨn,&*,��Y��rf����N�n�,���X�����'�㽫 ��9���|?��@ �ߐD6�%���A��5�Vk��C�t^�1�﮳m���ƶ>O�?7_Ÿ~����~?��C�ܗ|�f�$!%FA��!�i�2�ֶ�cR���0���{�o�� [jA6�܎���������te��,�����jd�A�����In>@�]���1�f��A\ ޻���'�11�)��Ŷ�^����u��;A��'��~ ����|@mȋݎJ�����y�wTx~7���D���p�m̅y���� oۨ#�T�Ch'��|g��������ڐFF�j������=BN8Dp�-�[�];_-���~
����*%o���\ ���j�-�>e�
|�U�6�k��^۾��/Q2\��x�72[�=O1�Jw��/V��\<�4V�M�9iǣ��c� �
P�^!#+�efR�V�M4.�g@ցl�Rŭ���[�ؖ�	C�-05*�*F�KU�i�T�܋��a-���J�Y�˝�m[[�����H��,�h���ʡ����E�e��r6�%k�J9m�#hE���KB�`6S8:�Nղ�\
P��u�n���Ү�HD�cU��SZ�}C�'����j�3ʅ�����5í&M�h�1�9�/�7�����t��/�m/�͹���~�����u�����Μ�{||zks�lY���� ����� ��[sZ�A�A=��ڭ��\J{������ �;P_����ۋ���W�O�� Av�$��pD�nEW��C�������D��5^�M\A�����Amn
����]��؀�G�r'7c���?	9�ÿWG� ��@>]��IǳE�D�>m܂p�E��k7���/�WfϦw���{����	۵ ����_�nG���kR�IJ2$ IQ�)�L�+h`�[�������]HRh�SQ��E����!��WB�{d�� ?p����/�}>�S��ա�67d�D]�@��������ڟ��z���EW�����v6Ѱ� q�p���(������&���d��SO�>�&w�\��5��Nj̹�� >�?|F4�7���������sS�_G���~���|)(�&�=�r$� M��mO��i�i��13�Y)��Ľ����S�v���m��ł.�P��n��]��q����<�j�zNτ;��	����G���RcAxԐs�D6�%����h�E�W��,^o�s���3�~�njo����_Fo�H-�?7[�r���V{�َ�ɋ*l��9��3,(�F��3��r=�is-ʁL�w��� ��A�_Kh&���0����^�x.�A������8Χ�`������������MT=�NC���f���8or�L����"������/�݀�-���L���>�:3�]�}�H-����-��<��	�2nbog��8;^ru�XD
������Nr�3�ڢX��*g�2
/h��Ov.B�kfȸDҧ�o1��(I[��� �mfh�v�n��W@���f���X ��ې$eN��?Fa��e��>#��S����ގ������<:| �R��hȵ�#n>C3�In�~mȐ[����l�޹V�o��~yLL�����mO�� ��W͵`��]xu�b{��@Ib���ѯ�*��	�sn+CL�j)I��j-����?o�~�e�����|[r'=���o?%�n�WG�njxMf�=GcB~;Ё���� ���>�\T��9�p�ǵ�����Gk��O�[�^>� Mm�#�!�=������|��s�z,O� ۟�������A�g�����<��S�;����/�{���Ch|���2Tzŕ~TA����/�͹����w?B�Z�_����_黍cjgz='CRԧ(x*�Y�T��*J�\9�#E�2�	ܮ��qMl�rq�=��Y�jM�."Sw����5���?���@ۑ?7|Am|�Lb����LJ30V����땼O�V��O�ն��ڂ6�ŷ!GQ$�3�����a�"A@��	L̬b����4?��%���D�L�<ڸw���w��Ї���q�-�����+��y����	��7Ým��/@� ��/�m/�jH���	��w�!��H����ޑ#;yϴ�?%Q�����~̈́9�"~-���B��c����	��m|�E�(��
t���= �U������u��!��m�%�@���%E�齸��Г���M��	^޿2�f��k�5�"5�j��T��8���n-�$7���g�
��O��6�=��DTn���{�9��k����-��kﶣ�׭�U��3K�P�M(n��Tg���V�MR�:��9OY�Q���/sv��գ��S��]f�{f�Q����TҴ
�&���\���H�ar-��K6ɔmڲ��T�)X�K9rUKVԊT��E+�[�v�LS%�)�T�WF��p�a���$D�����X�/kͣ�Gi���M[��Z�3F�YL\L���E�e���������k[�$iŦ���`�3��ї��f&�P2��ۋZ�9�#f6Ό��7��/����#p�З��8b�hJ�kk4 �2���M�+cj�U�O=z�=���I��|�V!��w͞�oqxt�!���fFɝ�� ���}_/�nD���p��+�wA�uײ�xq��������J�w����φ�xH?pz�-��/ڣ
��bz��RAm����܎�dC7���>�Nז7�E(ׯ����8Dk��8��%�D6�C�^^�w��{|���3�ṳ�P#�^nG�Ǯԑ�YqrkO1$=��ǲ$� [�xВ�z+^�n忚�u��+wݎf6��n_���w�P_ڟ��9޿,���K=}�&�C@m��tMPLcbVݍ�V
��QR!( ʘ��;��n/�o ��܉�f�w�Ws�QJ5���x��625=Q���uȐ{�|A ��܉���^�C�r��s�֥T����rꙓp���^FEeS5֝:�^[��]�W�]�+\�Ϣ��Ơ���Ob�R��xx�RC�����w���������z�}#�n��F�����I�'\"mȒ� A-��x��0�{��%nu�*_W����Ӏ��-�����U�q�E+���_6����S�܏#E7�����[�D��u�����;{�^F�O��܉���m����FJ�����9<�H�᷹:|'�ԑ� 7_/�m�{��s#W�{�~�[	��κ��rᕊd�:إ��u�JM�qVDP`��ψ?\ Aퟛ� ��c�{�ׂ�?O�͡@4o��LϺf}mg�CA�߷k�JX_I*Ȝ�6[�+�=�|o�s����uǂ�O5��=��-}"Kp���Ӿ�^*�<8D7�$〾 ��m�����-����a�x%���ՙ�>�+�\�Un6C!��qpT㈦��)eL�
�,-��-�����,��S��z6�#ç�z�Iym�mȐ[��7K�n�'�t�P"���sa|A��1繙�W�����xl߾�Awwһ������w@@���RAm ��G�͛�w���>�M�ϑ��k���p� ���������K����k4��L�2����s��iT�K3�f�Jl/9��9
��~~~G��Y��A|[jH-���ضwzH���^|+��>>��_����D{�_6А[�~n>i@�u���()��o�z�-����{<ڛ��V��.��m��׽cހ�"��@��) �����܈��1��������2S�}��>��_Ÿ@�[�Cn@�⠆[�ގځ�<�_g)����v�N��I~��������'e���}�K	
����^"G$��:U��l\���9Qʪ���\�'�	��Ư�V��u�AW*%X����(exqq��p����6�In|�8�T>E�fvk�^��y���xuO��@4�"��m_��
�ޮ�喲8�Z��u�Zu�XQ�R��Fa�l�Mf�*S9`�pZLA��w�?�R#� �/�m��~��7^FJ���G���@���^��C#<�1��F<�X��0�(<3�&���WO���?1��l����"3�wrx-��ڟ�=�"�6zc���;�I}�p�!�"An �ᣔA^Y�����U�κ���ʽ ��\
-� �Cp;�Wl/)Z��A3��ۑ��=��=&J���G� �q�.�n�:����Tﾽ���ބCm	-�D�m{���9P�TZ�<�b��\�$Fz��O�<u���Cq���# 1����h�`z=F�p�R3UOL-�me�mfX���	�����̼�;Y�K3d;�hkŪ�.S,��Y�en��U�����mWR�J��=��يu���osoxη������&�R������U�_K8��&^(d�˯��U������i��pPŌ
�O�'B����f�p��%���NN��2�;\q��]�n]��8�"Ő�ÿp�ӯw)hWQ��g����`��XJ��9�2;9�Õ�Yi�blK��jW�*���޻]đ]3����}y����n_K�z���mĆ���ز�9��,�*���r�=(���3�,��晤ilpʒn�
&PY������̨œ>�g�����K:�|����}�.�X���,R�`��݈���$7k_i����#cc.�9ݬЉ�w�H�6����է*�Par5�T�W�������i,�'nVn�vD��"0f�\���t5k��+���E��ݫN��GW�?�#��.�-�c2��
8"����Iٷ���1�f��}k;,l��<݁:[w��ob���y�p��rN��o^m�/U�eU}��w*��k�n�sv-{Ō���>��YFsP�̵}��wl����7\�U,6ovj��q�M[�j�vge�!vJ���H]��wJ��㱋t�[a�l�����	�-ɺFq������<�޴��sd��ܑa8.��Oެ$���S���^��u	�&��4��eM�;6��{i=�W����*O{yvwgj�ݩ���W�ky>�ry�D��l@�Km��-���7��E�.���n�k�i(�i��[i۲��n��+��{iO�����v9�;,s��Fs��9L�	�m�ֶ�tL�O��e���98��w��w�ݖ��+m�=l��A=�Aã,�蜥������ۭџ{~_/)���@��_k
{v�m��A[m4���P�j��j���>Y����yk�Y^m�%&��#��4�P�.J�YM��yX��΍��J_kO4qo�X%�! 	-������_Lb�"m��%�⡇JG� ��f�3F�rڑ[`�V-���x4�C3&����5&��*^�4F"�;jm �n��`��%�Z�˵�\�0�g�xx��̈́�	��t�	0lٙ�P��]-Qю�݉B�Z<L��Eљ��*,Ĺ�%��G �r[�,/Y��F8@�� ��A�L:ɬq�՛^ѵE�v�x����Ռ���#X��`
��B-�u�0�,"xZF�۰v�#�kWd-�Fk��V(-n���T@�ݮa�t^&��Sdp�
�]c��2��`�3Ek�5���$�#m�M�bP� �6�vXۣ3Т4w4��$����T�YX�U��D��7n��z骛uCb�5��Y\�mh$�v�g
�Y]�㴫�2ڶ�6�3It��5֠h��m����K��K�j�5�,V���!ZA������YVb��a���BV9��.u�����Lڸ�p��5ZM4X��d�@��k�ZU�eR���ۂmat���EB�M��e�Rk�v��҅b���hSj2���mw#�Ѕrb��Զ��4F	��pE�j��C�-v��	l.��ᶅ�A�\*@��V�ek�e�SkG��h��5������������kHƵ)רE����	����;60�h6���F�+a�X�9�	qr�/Fjxx���+͐��n�ci4��h�eZ�C��\ .I��i�����jv6YC�ǫ]��Yz�6����@��VJͨT]�k��Hs�����hф�s��+��	�e���f�6Nfe�&6�5�%��8�K�H�5к�a�i�%���2��h�0CDv!���8L��E�״�&���F�R���D�ٌ�S-�[�����W*핪�X�lj�]F�.	pɒj��j��s��6�����)�6Gj[Q�(�eζ5j�ܚ�t�Fd�l���f�m�bJ��r��4n�MH�n]�
&�J����].�HCؚ����A�������b�k´�K�Mer��\�� ƓKu[�IK,dj,a(.��"Dl�V[�5f��.v��֙�"7��Q�C����ƫ�����O���?�׊\]�f�ZX��auIE��b~��K��0nk0ڸw����C�d|���In���|��=��WK��Q��^�E���y<��{���
=�Rn!��-�$c/�j�ju�X�ٺ��=�8�^�F��������_��In:�^�5f�q���q�$��9{\\���I��w'��=v�������m���љS�Y�`���Ȑ�@�[�'sٟVE{=J6�9W��񬀁��_�����Ԑ~�A�@�ڐA����#�w�p�z�D���юw�5fw_�G�?<�#_H�[�~n1=8��������&��LD.l��Qau"6���Y]�Q�ԋ�X�Ŧ߳��L�/�d����Cho�t���'xn����Ӯ=��X �h��|~mȐ[�p�'�#=;]29׳�`��#&jn���r�[������u^�[��-�y!���{aK��3�š�*��Sݯ�(����K<=��A�S���ϲ⽞{^��� ��E��]#�@�Fd=Rn n���7~���A�+���:q��!/m�tx�8�}"Kq�����z���{Y�� ��RA���w�v{��Uồ��=v����;�;5�|�|{zD����n!����k���������l�e���"��9Z���@�h [jA��0x��d���<8]�X7uuIQEZTiX8�K��+�K�]�9���1�	��!.��ީ ��@7A|�C�u�������tǈ��;�Y3Ƹ��"Nt  ����%��F��y�	|)�ϧ�����A��=�ޝ���Sổ�>ڥ�o�&N{�`�y�p�����z��q���͟��6�:��M�*Y<V�
���L����9s�4ZU�f�si�EF�S졤H�,5�\�YF��=��w����=9�Vׇ,_U@� ����ԀCp!��-�o�f,�sP_�>_6�Hn��6������Ր�����s�˭��|۹�����m{FW�}>�����w޳�+'�w3�o�'�Ԃ�A|Cq�mȁ��>W��	~�fi�l9�+�K�\�ڴf1�j�P�݋d.	XȄR�e�G|~��E�%�D�!8��fW��x5[^��D�C�w=���b��7v� ����|�RA��Ŏ�`�:����G^���/o9tx�r* ���wRg�|���}��퀁�@�ԀAm1{ۦw�Y�j]�39>{�#|���Z��A�|�r$�P� p3��ϧ��~n�o�j��>�k�r} ���;^ߢwz���0�ʛ�lF�v1�
D�ͫ�f�4̺}ַC�Qǂ�Ň8��Aq�'������@C�m����FyCpm�������H�_�R$b���>�q��] �W���$�{q��?<�t��l'�򒫎qEsí�g(b.�f���!"���̂J�c����A�[jH-���]/x_)ʟ	���!.LzM��`�X�#_�r$�An �}������M�}�'�=�N׃�C���D�@����� �p��A|GR�sRA��n>M�ꜟ-[ީ綻��ˍ�����W����q`�p�6Ў�8�=�y�{r�k�����K��r+�w_�o���U���8��6���>��ý�,�D�/�m�?�A��]��հ�;��Q^���s;^'�H ��@�h [k�m�/�$)�Q��� ��D���!
��*�E�����ا/<c�C�o\��F�cN�̇�+�#����E�z�}>z��3RY��A�5X����B���鰴����1�!�lM��M�ņv�SR�Rj���
l�!cc�mZ<��-jVYH�����
���u����f�l�35�Ό�J1��s�c��\��S�\\��8r�3���6H^5�+� ���#�t�]Rl��u�����P��F�`���Uʳe�w�_~���$�uЛ4��]�fXMkU�#3�;���h$���+��@��_O�����G�]�x]\�۾]8z*%{'�Օ��'��9�G�����An#��zP�g�a5� �=�=힝��r+�w_�	yj@#z!�=b֑�8N�U9y� �{a~�[�����|����n7\�����A5p�m�!��B�j9���Ε������r%�h�����Ҷ��ˣ�����A27\z�G�D��"s ���!���g{1d�w��u>�&�n:�7_��S���q�6�V{�8��G�>�k..�D]�cJ&��hi��������h+)[f��ez\q�B���В�/�%����3���'g��B��P�ӮT��@�r�h"A|�RF�����̵���Lw��z�E�An��2>�������Lܽwo�u�]���S������CkDI��7��R��8�����t|��G�?xE'�mr���@���pi�����h@�G�ܿ�w��E���m��sCv��"%��/�o�a��[���RA�AK�ۑ �D���o� �t���B�p���{O��Q�2�|O��M8�&���xp7�ӿzq}�� �n>m���3.�#�����^9y>�+{�)�-�����\"7܄�[�A���lD^����a��
�P�u-��.U�hم!.5��2�e�3R�A_s�5��� Y�"�R!��޴�p�񬨗��l�w�g���-�u��z������X �[�F_I�N���k`ء/7��z�4el�<�O�����D5���h�*���7�����|�BA3��ϵn*����N�HDNU�1«o�����^{.�1��4O8v���x���a@u&�D��P��L�N9�m�Ѯ4�(�jm2�C܊נӜ[kˣ�M\/�o�D�[��!�2'su�-Qˈ;|^5 [A}��\n��5���-��j~#w�/�~�s�W��?^t�-���n��r'��^
�ʢ�)���y��]7�f-[^g�i�@��"�RAm����7�''�WlA��$�	)Q�H�������VY��Pf\���( �L�I	x:�	w�A���-���_�w��8�חG��^y˽��yq� Cƾn��E�q�T��F��Ϡ_ϻ�f���9fe��ف�Ԃ�A|Ch�"sV}5;"A���;��mȐ[�%���ܟh�K�S~�ޛ�ʍʍ�����1��m��@��A^y�>�J������RA�� �K�ۑ!�豾�w��6�חG��w��}�z0J�J�D��8v��J�GSG���Y����n��Iݫ�Q��n���\jC��f"�e	ي��/�����|�B�n!����z��,�40T������|;�(�����ԐGr/�hV{�{ON��s��Q��5���vૌŬ��f�Xfp�-���K�0f{�8�[E��?���/;�7���Q�����}�ʣUs���S ;�۫���6�?��Z�!�����=��Z(>�o��t��G� ����_7�=�<o�Q_�����͠�m���{�C�e�;��۽4�Y9�p)���]��9Z��܂6����OŸD'qf���[�\����K�����{*7.6�O�W3��ͫ��о/|��������n��fTߎm��W�"n묙�{�L��ڟ.�|A�>[�� ��� }�ܜߢiR>Y�w��T��V���&��M���Y�*On���ZCL٧u�BsBH��iZ_$۾��U���(Z�^
&��5���kN�jd�l1�X5�	C��M-m�S��b��v�B��=C�6v˵i3ԋi��$z��80�'i�i�����eU�)�Z�0�T��a*K����J&��·L�ZӮs����ؚ��5��a]\\��&�����������[� ���Nv�W*8P��E������f�D�]��`MY�L�эc�1�4��l�/���_W@���Ԑ@m�������AJ�s�w��N=��,��b�r�h/�hH-�[���]��v�9Ј'6>����Q{�k���A��� 6�m���OGVX�c" ') �����ۑ"W��I��DH��'o��e�V��tx�!�H8�Kp�!�2:���Hz�z ���7�)!���<!�ǡEn��_^ڒ-��^��bk�8{�=�/���q����r$���ŵg�P�,�_uv���e�*2���ܟ	��@��h"�_Khޚ�-���%�6� �YYA�Q�F�ZrՖ���G�׼��������f!�,�|L�E:�G��N!���!��OǺ�"r$[�����'L����h���ǏԵ���Hgk��Uav����{�̘��	xS�3]crl�7*�$\\�p��Ҝ��n�r�d�2��u���~ ��A>�p��˱z
���]��T��AްI^�^���\�ބ��_@mȐ[����Y�oU�xU����|q���V�߆ܡ�Wm[jA��"B��={�e??*���폓�"~ݻ/��%Hu�^[ �N�E{�=�*��>�G�p�m��	n ��@��WsDg���[���xW.��
�s�tv��ڂ������m��X��RT� �~�߹�k*�n��Q"�l%A���J/���%����et�}�d|���$��p��~��v_���6�5_���������A�#�����n-�$<Y��.fL�\8����'۷bW��鈐�f��}�8Dn�|�M��y�d�ѧz�D����"�_7~�^��9Q�/�AA�"�s���nQq� ��5��vL�V.���^5Tr����a2����58���`:�M$ک�w�
>1$��Mƫݲ�NYۄ��v��Fu���B�"�\�ϑl+r�%��b�]�-Swj�#`�눠����o"��+kl=�j�p.�w�{����ꖯ#gw�1q�r���'VL豐�v���Nٺ��Ң�y]\�{�=���M��	�J���'o�v�^|{:��yf����J��}�\�[�-X�pu9i�`��6i�H}�6���B�TNt7�s��aovO3����Y��oMq]\ܚ���~i�������j�R�j�y�b�b�,*��T�z:�����e��z��ʠ�#0�U_eGo���"-�8�hB��$���ߓצU��nv�\%�:��,OG��N7�1Iч6e��,��j�q�mtފ��R�W���lՋ:��~ȸ��os{v���u�:[s���l��zD�P1x�Q���e�|���	3{ǭ�rLZ�sS{�iR��� �*�B�Q{��Hk�[��x�x*0ފ;67x�f����v�ժ�:�������z�7��\T���Ug0@���:�4�/��Q�������0e50�eMB���T��da�ؗ��y7�N�S��;C�s�޹zi�/g!���j�Yosm��b���e��:n�:�V3�^uw3w��3E&�4��,���f�v��ݛb���o1����$L���k�$����9��{vm������f�s�"����GK�����ND�8�<�o{6����ېs1{k��N�~��q$��/ϝ�ۼ��e:�;
|�~Yy�%�6g��9��� � An��u�&)���v�={x�՜����+ه��3��Y���0���~i�V|͵!�DG�~����8Y��QN\綧�$����ᶨp��g��lw�q���֥|�q�$��p	Qm�)�A]�f�����D}��ﶿ4r��sn���r�V_/8����.D�ݶ�R�;:'��v���vR'Y^�wg>�u �r	��$�I$�	���x+��J�s�w�?�RGln>m��7�*��DZ�1����vȓ�Kp����b�Ƴ'���k���UcԦ���L�1��E��Ch Cw[�)ib&��T�������o��&C���q��8@���[���k��gk�L{ĸ�!��
9[6r�\g J�f�A(�R�r��ݍb�W����d�g �m�������[������C�9�6�q` � �#��|[r$�| �?_�}>�)�>��z��������dc�r��\G8�[S��fr��ր�@ A�k��Y��6�l�����G����F�2%�_'�>C}�$�#�p�m��V��Ɉu�������ƹ{=*�������3�/S���fӂ�Ґ5T�e��b�޻}�5���YX�[�iS>]}ۦ_�g.W�
â�`�b���>^G�}��q��� A�n2*0w?�c Ǹ��}3��߇9���4Ŷ�nG��;�����=sA�5c-s
e�,��6�ґRlh�m�� ʘ�!h�`_o�} o ���-����3վ^�2������Y�ݛu;W�=���[�Cnd�p��V���<d������~A����k��yos×�@�o-H �����ߧi��P��N�D6А[� �Խ�HLTtם�rg¯����H&� ށE��������=饸oݔ�y���@/���"y�Y�z}��ڿ' eG�(v8�ʮ���k������B �܏�p������zA���7�y�w��ƹg�Ž�^@�寤v��!��m��9����8����f<�26�	ж� Ӿ��gq��b�Åԡқ�~��[�Wv$,�j^���u�Q���i#���m6�h��U@c7]�Bl�ٱ�B��J�B��ጱ j:V�:�%�Ԕ��1�5�,em�+nA�i��.�:�6��$%uL:PI��X���h0. �V�9H�Y���n��2i��j��K��˱#�������v�2�M,�j��B�7=]�!p-*C���ԨLv���7@�BY�a�
�b��r�{�}�q��`�C�fbP�wg&���R�e�����h� ��~�������_�~n,�[������L�U���&�2.���{�� ��jA�#@��R�����Q��C��?sr$f���t���ڿK��l|��H��v�i-�y���s����E���]���V��n{���8����<#��7��� 7W͹q��A�el/����س�n���6�υ^1�Ó�j�"2ԟ:>�aV����$���m-�$���vz\ſ��$N�>�xȊݫ���?V� ��-����U���۷���
��D���at
�B(��h����3sl �L�*W�D�Z��o�"�A�R!��tw���-����5�g'b뻺�r���6�In ��#z�|�x�J�#�y~�c��uh��-2ӴD�N��:��ۓ	ˤ�י�D$p��X��Xaɐ�����Vઊ6!e���Ʈю����	��78r~5p � �m5B�ʚ�4pT$t�m��6��������}p='T����6s2^��j�.<&�>M�D�[�?� CndL�cƫ.�7�� �&�E�7�ܻ����ʋ{~�@�o-Iϐ�Psj��u���dIn n(�ۑ%���wa�iuwq�u_	��7<55���/�m��90s�n6�'��D�FQ�22���L�Q�+�:��,c
j�%�G{������Ϭ�9�D7 ۑ#=�gӾ���
[�~�]:л�&j���>���}�[����~-�D.�3L���W�~ �A�wO/G�ʊ{~�_^Z��A�L+�B�����!@����@��p������Wղ��"�ۓo.(ȥw���{,�w�	g*��X�nf���1��WRv8�x��%Q��B�p�fHn�n�*㻘r\�4U�;�55���ڒm�!�#W�*O���ǔ�^XA�A��ʹ$gN���_��A-u��v��.�&�1Ğ�Sb��q�q�ͻ�Kp�ʹ|��֫��o��[����r��߇/| �Z�j���nE"�G}�'��Y��P�%q(�8`Zcua,�m�4�^�1�O�pB����� �}�?g�p�?c�����Ց^��s�S�l��z�p� �cS� ���K�ڒ75���:��] �ȑ��/�b��>��=.<A5�� 7�p�*���I���j#=�O�:���h/�mI6��C�����/&�WF˕��#��^ ����m	�@�[~�~��3h��q� �[�1��ub�Q�q��= �� ��K�g�s�+��2~��7q;SZ3T�[\���Ve��&���۹5�7��U��[�j�<�k��j]t�l�YAo�ӧ����־oP@�mI������dm���_�~���Q}>�k=.<&��O�ŐKp��v��W��_"����0r�:\�����c]·Aɝl���3:6�;��Aڒ����'����F^��7����E�T���/��G��܉����|ڭ�[ٛ�f�w������o��wV*�\c����j� A�A|[i�͢����^$	{�~ ��!��6�e�%����͉U�s��P�k=.<հ�-�D��"	n�-g���^��%d��9��}�$�h/����z��.J�����ӵ�������f^��_fȒ�/�%�@[r$��<�߼ƛ�@{u�>Ɍs��<'��A��ChLVƕk��z�6&aI~�(��7�a���6����٨�L��N�+j���h��vFM֎P����v�Vp۫��H��Ͼ�e��j�jj�CM\&���Ԩ�L8�h����lc1�[�
�-�[�[,�1��p͆��,c�K4��ζgV�vA��7�Ulq�F�E�cX�]V�m�ٹ2DI��3�.���lK�i�Df��xoYY��v�)F���SLݜ�f�Zȭ����bg-�6, 2�[,l��go�I�x�Ja�m������f���s�;� i��6
�Mv��f��;Q���%a�uf��B�� �������m���-wپS
����ӆ�c�'ѯX#���t A��6��� E�_&�^�9��
9v��z��ڼ����䬽�^@�iڐ=� l_kJ3>��$�@�wam��ł-��z����j=���UV��;�5g��M\�o �m}!����o�}Kc�ܹQq����܉������*�n��������Η�:��t��ﲣ> �saۙ��Ck�����A�X&y]��z�yь��Q��/��_ۑ���?>��b���,�K�`����]`�tY�.�c�5�-�
U�ꪖ��~f��#ު�&��#�U�An��{�]OU{���垑��u<f2��{� syH ���mH"��s��6����D\zuLl,*\n�m��yF��g˧�2���q�N�����Q{�Vu$�V:����׷��<<�K�������Yޚ�n����|v�~o�In/|5�����ng�8[A�RAm��L�f�_^�6n=[O�.�#+o×�&��;P��ۑ%��7 o�1UOn��}�>��_��,}�s��a�;���A5pl���=9�h_�� ������ [jH-��!�1q����]H��p�^[���nm�z\x��D7����?7�����_����F�D3cr�p�GP*�ò-�ZMb2Ҧd�2�"&xus7� ��AڐA���^��^��2��9{�#�>ɄbGNZj~#:#5/�m����A-�!MW��s=�$���<�{���U�^�.�<9b���	��;WQ.��jA|F��u��p,��|CnC��QȤGgg��훿�t����I��h��Y���C:��Uh��uي�r���nTiAS�u��7T�m
u(UrK�z��)۬��� �r�[�[��n�����!x��Gl{9I�1�{�\��d����&��z:�����b��K�3zD�[�~n�?7	��ڴf'��y�ez�U_������P<A�@�Ԃm��s���r��y�ߩ�K��u*��h�{<̒�&��ԊccA��b��X�T^O�7ؤ��n�_܉��{'�y�J�u��#�l?9Y�2܉=Ё��"s�[���N'Rĕ;#!1��R#u������>�����n���j�q����|b��?�|�nD�����WJ�n�{�~�R�W��nxvJ�gG͵d7A
u�;�K�KH;���|�C:X�t�N�f���q�9p�#>�o�%=Eu�J(�ɬ�Ʉ-㺶�ʕ��;�eh&r�0����կ҄��Z�s�{�vȃ�����J��u���0A��|Cnd[���m������B�>��t^(����7MIv����!�"dd�l �0$�3$�����X�Zj������ͻ~��;�f����8_���!�>�4,�|~n-�G���;U��8vO�z�dxF	�����#�9���@7�m�u6n'G����>A|G7"Fm1�3����N�Vz\{�	ˏ��Ȓ�y7�o^j߻���$pp(�Ԃ�t�%�d�s�G��E��r�@�n��{PD6�ʹ'��"7ۢ����jq�����t}e�Bߏ���&:�ʝ����W4w���Lv1��R#����ڐA��!��z�XQ�������(�g��΢[���A��A�ȰE���?�?X~����UU_�@HHHKh� $$$'��B�RBɊ?D]OȪ��+u�i���?<ю�@�� ���I'g��e�F1*	��HB�@��=���u=���&C2���?y=�RB�/�z}�ҽ�kٯ?�<|��:��^�9�`l�H��Nb��k��^rY��^��R9,<���w1��������y�z������!�|�HHHO���BB�|!%�a��}!�����]���d���/��a��g����Ϝ���!!!9� ���\���*O2K��	a���j}ҍ��{P3�~�i%�0_m�3���D?q�>�����U1'��$!!!���:������2�JaIb~����Bu��u�Qekֶ�W��ɰ�������x}�HHHOI��J��C�3�=�='�?xLB��>꜆�����:=}�O�vc�C�IG��_���_�G��@HHHL���u���=u��O����f�Q��ٯu\�J��~ﲾ�����!st����=���~�>��o�����>rB�>"y��>�,���s�3�)�HQޡ����=HBHHL���������B'~�uԞ�&8=�~S�̅<2O�h�$	!!4=��1'�K�>��'��HI	��(�6$�����E��]4�������kT}��aU�g&9aA�@����K��}���'�	!		��>�?�H>��{ �0���O����z�N�x��Ot,!��=�銏�>�B��|����'�����@�g��}�����
����Q����Os���QRO������$!!!*O�!��<��������s��{�����P��_p�a��$�Q��(����oʾ~�3�����g_0:���޿���Önu�{�����2B���!���| ߭|�j��P�Χ���Ԟў�o����`����$�o��H!$$$'�ē�"{`O{�O��ɿ���$������|��zh>������R������s�w�P�B}`�ĢO��HO=�s���H�
�p` 