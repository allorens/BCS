BZh91AY&SY��/F��_�`q���b� ����bH�            ��R���A�m�(6em�)@հ�U��BD�B�
RB��"IB%��l-��R�)�5A�e+@�����R���ݦ��CZŮ���ݺ�U�.���L۳v5j�+�tm�6[
��veH�V��ET�٤�ML�P*Xiv� �*�o\�ݔ� C��O@ ����6�[[l�4�;���"�[�t�*���:4������.���h*�l����u���y �D�;�:.�  <  w_g��nҹ����u�����q�7ju�];)m�Ӷ��vK�#6��]uwb�ڝ�AiZN����p��;������;��ʕ6Wl�3� �����-���Ӂ�MH������wm���F�>���t�AKco���ؠ6�p���-�T���9��M�bm�](�}��ݜ��t�W�T�[-��|:u@
Gu�O
Q�Q�ן}�_GL�W�׽�zP���}��D���׷��뢅Ic�֏@{a����*����k�y�(JU#�w�� Բ��Z�qK��V��퓦mF�π@m�h�kR�7l��׺w���ER��=��{U�*ޫ���CE�O{�u�V�>�{|5k*���y�!�>��(��wt�[%���Հ��vm�6��j�> �QBs�����cwM�U�gm��f�k[i���^ڭI�'p�n{����ӻ��{�46Զ�9� ojj�[ü�zzQ�w�}{岥�ў���wj�[[]�z�CYh[T��E�   ٷ��ZiTc��t/V�jS�׽
�չV{�w�Pn�כg��`m.�����]�on^V��{/x��k W�wF���VOp�b�=ɥ�ۑ:��wsvaUV�   !�6��=�t�z�U�^���N���
I{�z�e@(�W{� �+��UO�9v9�:Ǟ�^�(�;������U]Z�N�t�@ʷ�  σ� �ܵ�H��z� �G�NR��u��vv�n:�$nsv��F��s�)�һ�8P�F�]!@WB��Sjm�����&�   .|�	�%@֝�w
R�/z{Ǥ��v�t�n:
�7T��SX�.*�B�'w��{�8�+�j��U&���GY���u���  w|R(��q�UE,Gv����z�P�z�n}��W�|�����u��Pη����.䑦Um��UU>          ��R����` #CL ��S�IJU �10 #L�0�D�b�S�       5O��ED`4��!���##LFS��dJ��2h��4�di�a0����T̚)��4�4�M4a���_����5AE1�ڟ��ׯ�������^�����w�{���/|��{���� U�<�?�U@} ����TW�ߤ� *����@������������O�����j��~�
�������t��d/�>������������G��LØf09��.`s#�\�fS09�2L�as�L��S29�̦e3���f09�̦`3)�L�fS0�fC2��̦ds f09�̦a�3)��f0��̦`s)��Lf0���&e3)�L�fS0��̙�e3	��f2���&a3	�L�f2�f0���&a3#��f0��̆i��e3)�L�fS2��.l�́���2���as#�G2���`s�\��\�29�3 f́�\���2��̎ds���G2�fG0���.ds�\��6e&G09�����G09�̳���S09�̦e3���&29��ds�\��G29��g0����2���as���fS09�̦`s)���f2��̦e3#�L�f2����&e3)�L�f0��̦`33��fS0��̦e3)�Ø&2��̦`s f09�̳&e3���G09�̦e3�	�̆ds)���0���L�e3#�L�f2��̦a�s�\��0���`s0f09��`s#�\�LfG0�I�̦ds fW29��s���fG29�̦ds,��\��29�̦`s)�&2���`s)�L�fS10��̮`s)���S2��09��`s�L�f�2��̦`s	�L�fS0���̦e3	�L��09�36`s)�L�f29�̦`&s)�L�f2��̎a3,��L�fS2��̎a3)�f�fS0��̦g0�a3	�L0���&a3	�L�fS0���3�L�fC0��̦as	�L��f2��̦es f ��`s#�L��09�̳as#���G09�̹�as f2�es#��f09��`s#���12���.es#���G0��ds���G29�̮ds0�G2��̮es���G29�̙��329�̮as#�\��W129�̎ds#���0�ds���0���.d3��29�̮a��	�̎es+�\��W2&l�+�s �`U̢9�G2!�D&U� fU0(�W2�� \�#�Ts ʆa� ��0�ȃ�PsdÅ9�2��V`�9�2��Pʃ� s
�aA̪��2�f�Ƞf\�#�s*�a�9�W0 �W0(� \�.ea@̦a3�0`s��2f09�̎ds+�\��6`f29�̮`��3+���09��.`s�f��09�̮ds+���G4�fG0��̎asf09�̮d��fG0��̎`s�\�L���.ds���09��?�M>z�� Y��O�����iMW��1����=)I��9zTp�y�ۨ3��X��s1��d��B^U��sr����M[z�ln�er�I��lX@4��~��rd6&�P�c*��&�8@Fd�EӨ��7r�nS�
���u�����w@(��X9��� ��O5��5�Mٔ�i�T����e,2�ʂ��c�"b��+�V�3Do�XQd������c%���&Y��X�粌�.�V�	r�Fk['l���ۇ4E�a_����,ܙR[�x`(Zk&U�$C��Z�l��pV	�p���9R^:J�]�B����A*���N�ףU��໼W�!E�k�^Xݙ,;@����׷rl�:�e�T���	 cc�fL�˔�V�0K�Dν�'f�jb���i�7F�;*V���:30)��5"j��2lN����z��uL�4.���j�0�ۈ�ZN��D�Vy�q���� 7���P�x��!��e^�7����î$�ب譽���eY�C��a��{*�d�`�"���$��V$w��!�,T�@͙Z�����@.�2��Ʊ���v���0r�y�r��St�&���.�� �:~��L3N]K7Th�W(�Ci�`e����ӑ���Sciƨ��Deh���V�����[��^lNBi[��D���q�钶u�F�)�7XY�0�n�:0@"��qd��Y���ѹ��
W�r:!fG�kx�%̭(ۦ��{BMW2ě�f��;��o6��^�f�u��`H����n:��ͥH��q9Sq�9�U%%�4X���\�-:�����u���J۪L=�0ڹ.�����P��]b�"� iz�h�Y�H�n�[LeF�uy�V��j�^�5�G������]��2&��f�&K������*���T�	�ė��[�P���ŏa�:��4D���R���	Z-�xU�8�Z]{9F�ȓH���Ѻ:�c�h�B#�lM8�jo�d��t�N;cZ��Rӱ�m����!w7p�	����D��۳��j�1�����m2�7IC����q�,�[�X�j]�1.(�p�c =�+hf��V�5ɴ&����ARQ\V�W3t�16u*
-�㛻1e:r������XV�d*N��a�;ơ�Ͳ^5+�P��,an������x#osÐ�ͻK�4��;��� ����q��2�j[�M��M�̕���N��i�j�P�	$1�����9��ې�	S�/d�ͳw&SXM:�nM�X�Z�v�*�nR���V��V�3�P켼��e<��!ЅX1�<f���N�g�"c.�U�j�oA�>�SXrҩ��70)�V� �5St*5cq�4f\.5Ck3N���e�5Z�R�r�b�l�GI�ejrn�6!��f@�[7���ֈ��bL��1Ӓ ֻѹ�2�t��f�m�MP�gaZ�c,��%!N;���-�{�Z���LH֙Twn�V%ABJ�'��t�7#y�eALP�-�0k�ݲ�h$���᪻'2f\�H��損uPM<.���V��A�ˀI�eјVjrB�\�6�Ql�+n���O.L��x&cv5���UL'��� ݝ/)�^�b�`�^�������
YX�Q.���;'~���7*8�f�:S�!�1޿=}.񓛒��rEV�Z�WpU����[��o:�3Z�! :�!��K�8^�.)��R�{�v%fh
�Zé���-��H+aDE˼�i&m�]^��WsF��κm��#��9tF�,�L<8��a6���u`7�ƽ�1*�i��0V� �w{zC��Pq�����M�����*�.�b[��`c���T�=���z��(�q��)"Y��W�4�.����Nm��`/$�X�-�����:+D)�ze蚎��A��4�0� �y%�
�I�N���=tD۔baр�SXu��ܫ���
�(�#*pYvM51��!�[�R8ƞG	��d:��ZU��At��.��b���ܜx�7Hr�)T�ƕf:6�Cf;���6��[7���o6�١��If��N�q�3Pv�8�)A1F,��tr�z�m��-�*nZW�&+P���pej�r��y�n1(��j���Ӧ�����uo2��"&���Wn}�LB�
.�X�a4/p�r��Q{5%2&��ڀmL�Lغ�j�;͸��03���M�43R���ٔ)����V�,��H�{m�v7S37
ݪ�7[ߝ�/=��s]қb�ɇ#c]�p ��zn��Zm�l)6���|��ؤ��T�B�%BLA��_����9!b�c�dP�����͇�'�D�w��YsF�^�᭸���1/2��u�[��E^�<yTCMɒ%�eH˺z�	��� x��w�^�H���#	�lm�N�v8����n+�#ħ��7t��5V�n�L:r+6���0K5��J0*oc��D�5��CH�/�P��M\ح �Rdb#I�72V�p����+<�(*�W����a���Z%�w^�q�s��VeP�-a33#YFP{���������7-�D뱛�]��o�x�f�Xu��o���5������a( .��P7fPO����(��˵�D�ɮ���SY�`L�j=���ir������Ej��(�#\���׸�\�KdhPxE�L:,�kYݲ#�B���7@���E:�7]�~r�5���Q��Są˵x6����[���2��,�T�g1nG{.!�S�oFsh[�F"�ZTH���֚���m���zCs귋s��I�ԖS����w��6e��ћ2퍫mb���5����XE�!bb�M$6F'5A�t�ݺ���%�ZW��z�PV�T�Ԗ�-f�<a�ۤޘh=�ڨET�z�8�{l�C[&�d1����9D�u�����e^�$�g
�o�r��F��2���Ac\�xn��� �f�.��k.2ha�{2f:�N�]d�D��W+`vN�6%[XYJf%୛Y��2�(�Pð&��ff(h�O�pXU���ͧ�[퓡�CL�Ee�fT{cSf�q5��u7ef��z�l^<�]b�m�šQ5+m���,k5)��i�7� ��4�2���(݉.��X��W6��"�\[+a@�f摄M$"���O`��*��z!�oDdǔM:"f#kpݡ�j�ki��YbA$	/Tz��FLk-�V6��{5���i�F@-�*�17N��Z�Z��r��%pFklblf�<9�jIE�$P��݈M��HS'sVℜ���Dx��p[��šR��[
�P��*�n�"2$j�x�����y.��)��[V�-C��o\ͤ��Љ�E髹�n�[��b�(e����t���W���;N���!b�P[�`*]Ha��S����U�T�Lխ�`I��db�%���⬫���U���Q]�
K
��bo/V���Z�:�l U܌��X��uU�]PsN�1cCȷU
����ܡ��Ǖ�[�oJ� ���m�B�ҭ^-LF3��ۓF�u�i��i��Qn�j��$*��Ŋ�V<O�bh�Y�At�K�L��mʴ2��1PN�f�{L^�~+8#-T���s6�[��&��=;YKeG�5�+J�v�1onX�2AO-"
/PF�1yM�7�JSR�:.���Bf�kl̊�����0i��;�iFw(��iј�k���y��iz�Y̕p��n�vz�$I��޴Ь�.�zt����[Q�����-kU2��r�G`�0�wn����h�h��i���"t�j,�aU�!i^�
p\Z�k�.��*e*�Eޛ��ݢ�Hq��ӱ�j��׶���&o
�S�dd���`�+X^�6�^�I�:��T�u���57�*B�c���D�*��a3,Ӓ�֪.��ܰd9�����sՕ�wN3���0V)�1�n�]�]�@�v�
;��\�BÏt㹞�,V�57J�(D�K���[ `�V�oX�^n:j�iw�{j<Ư&��[z�+D	�s[bv��d�!�{v�əGo/V���C6&fY�a�U70^�l�&��f��-�7%���t�[(�L�x�
V^�� j(��ɍ�&ʹJL���)6Z�Q�) ��T�{��:(`d��1]��ܸ�Ȑ�H2��vUL2�������d5$��[&M96]��fP)��+Phj57L=�i�3Yk�Z�L]Y�t�af'��ݲ�s������ �;x0�1r���5�i�(�x��X'DOcr��.V5A��O2�ԫ��>�m��I�[R� <��AN���-fR�ͱC�BI<�ΌˊS���oeI��4�n=���XZ�i�$*���W�S#ܴ�Ǥ:cK�7fU��&恺62X��R���I�bo`L�ݛ����WHag^�rط�R�m�PPӶ�n���X����v�f<��v�b͊���c
�!��.��ʞZ�-6��.-Q�c�.�*Q�v:�Z`�*�pl��JX��h`fdв��{�COqRF�Yd�����=x�䚋�n1[k*\ySՏ`�0����.�Y�M�˲Zj�
�'�=6�^
b��BoWۈ5��Q�O+�b�/q[��X��a�����lQ˺��6�Q�kww�+s]��F����J�a�]އ��L(h�Z΄Nm��ʧ�c�fA܌����$��m�
�<x�R���5^�~�^�z��w��ŗ�*��V6q������:�E�%�f$���ev���9����׎hM`��^H�n�;f��Zbv����dd�Ncf]9�-��~J���06���W*Y�S]��T�,5��:�L��۬8�v0F�E�3,�������n�lV�60�ہ/<��z�^)	�f�4Z�am�����&`���( ���M,�M��e��P���7��!���C�f�۠�x�PS2))�44Qb6�(��e�{㨹S`�����˱���FJ��vܳVк����xX�($Ve�$w\G\�ԛd�C�Q׍�pԽZZ�v�26���ja{��pcut@[׊k��gov��a��xE�RM�Jˢ�]���1�[�Mx�cn�˭(;�+em�a��;�/q�ȷv]�j	۴v�X1��qX��aGH�ím�%���Ah��3�{��n��m�ͥ�.	����GZ#oRlJA���d�V���uaҭ�V��rG�Q�e A�ڶ5[E��1(�HiS�n5��K�^��T�`���N�_(�4u���ԋ�m��m�3��[]&4di�*��8ܭY�m:ǈ �����c��*�F��i���.�mf��wz�kZ�t�=�%���H^�1휛{{E,��n�	6ӓ5d�շ��TۛX%�n��ׯ!��px�䕢:߆�UD�C�۫�!Ŵ��'��3FԸ�����@�T���Q�̦�J֗�rݥ�q�w�\�t��MF^�De�=��K4��)�(���[��yn^ނ�XP��CJ�zE��KeJ��`�N��D��Xȵ�	J���F\�iz1�b���x��2�����0V-�"�	���52նo-�RܲI��1J.������@�(LV������7F)E�a*E=�qi@c�-K�F5�X�5q�ڕ�z�Td���=���Ԩ��"Ma/(�(Y��ɥڃ�u�YeXd�vltse`�E�����1b؞P�>gt&����
�*��.��'�M\��4�ݸEK˳��b��G�%�Y�]��B��G���`��A����x#S;m���-�'�Ŗ�SDFh�u�07ކ3R��w��^є��pZV�0���Q5�[�d�x�Ub�o1�4�v�]����Swnd��
�-���=�iee=t�����6;WR��:��l,�'�&~R��a���Ȟ�����j02&�_��|n�ZB���3�hTe�'ir��bU�6��by0��K�X��0�u�� ـ��/AJ��cHpg�Q�3e����$u
&�\P]�ܶ8�gi|TM�|LI��"VJ+�����U�ˉ�>.���87M�F�@��9��.����k����^�Q�f�*K�^�ea�.*�Z%���V�s*���V���q.Óqq8�bs�a�Ш܊�V%�&by�U���:��<UVM�PQL�/���8�_��tL�6ʉ�[=�x Y���|Xz'8�;
�L�w��nکv�l�;�E�lv ��W�������P4����w��2$�3x�-��um	@�F"��]��1���6֜������Rr��x:q<]����N-��W�Ҕ?��6���gǙ~�0@�ĳ0ٍ㘘���Tp�r*V�rt�7{]��<\�E!�,�bc�Bf6��Yzm=���;fD���3Z��tL�&ʉTTF�����Ķ��^�"ͧ�F�L�=�hS��і]�/�d2�k!�҂�Eٔ)�C|(��e2|]��x��#�4�b�L⮣�'-z�hr8�)��;�x�M����Gx����+����~0*�b������86��|='���&PD�/mՓƳ<Z*���e����� ��H�AoJA���>�|N�&U���ܧCb���3���bn�'�\eL�D�>�ۋah��E>�,�|M����0tX5[W�`M���SfG�݆i�vq;���ؓWK���4yQ0�|�[�A�4M��A�#��'Ǭ��ع�M���������p:ÉH,7�`�{S�*;<�Q�F����㰸]'[h�w	��D����_��E~�I��@?�������~�7��f~�&������r^T�̬e�P��˨�+����ǋ�wm��o�����C�g����L���K�����C�c�1T�@8�T�r�^m3E���-���´��ښ���)�*ev�͕WS�prnVY�3ƓQ�n�����j�`�E�%�%���\F���u�29���Ⴖs��8�9�r�s#s��l�;�R����n��*�W�}ۼ]��M�2m�\��b}�cϖ�������/4K�0�8s7:̫|�r��3tH�YB�e]�m� ��W7� �T��,�J��r��3:q�1)�.��˩��'������S�4�u�z������m��Si�|' �ѓ:[q�����;u���5���.����b��SNcvd��!x�
=���fMj��#��8㡬d���z3h�=�y�MZ��q�`��kۡՃ��]�N�����D�Z��r���sD�u����������N]�TOwp��R�z�B�P]��eu�:�o�����)0���w]�xp�P���F���SRì9y���Oz��� \u�D}k]�׃$�&#�=��U���c��u
%�j[�	\�&�Lٓ0�2�iH�g<Q�����P��9��)XP�'\�.�&!g^rA��\nl%bh����nI�J��2�gr	<!R���R�{8�'f�X멞��8^]\9�!j�v�p�w�	��-n�`ur�Wt;1�MC˃����3r�Ӷ��k���,#�������V제�elњ5RZ�ɗ!-�l������Zgc2���\�7[�:.��|�q����4��q��Ƀ�OÉ9
&QK%���y
���J���v�LJ��8�A��3qq1���wa��d������x�u���Oh8-&�v(d<��;�vں��I/���Z�ہ5˧83E�,a^v����"�v��=����+��ͳ�uGͥ�1�����hԔ�8�ҝ�R�U�ձt�
�-�ngF�"\�p��@F6Ʈ�%���7
d�r�(2�I	���|�ulf�	��:��H��5|{���b�F���Rج-�o���y`�|�ޅ�G�}�M�Q$L⻩e�{m�l�et�.��\��v��	w�kc#)�0�]�l]5��h�ʋ�e��9�(0���FAǈK�y&p��k�����-�G#r�U��p@��sI-�&̬����F����Y���<�V�X�k��ۻ7h���.x5�J��R��Q�)Dt��8�F����}�8]7]�[�V�KǪ[ù�A���/F�@�@.;��6�N唸e�a4�f\ ۺ�0_#0TQi#��>L�GoykU�� ��6nVR�U�hIh@R�!���@6s��Z���tKIp���.�?**��I��s��[�:x%x�N�^�b��j���WX�{_��[�Oo��Gڄ�i:�Y�-�+)��}i�т	�QL�7�*��`��?|���̛6)�iՂ����{%��.$���x�3�hn)J�ci�;�j�d�.��F�9vmA
h%�<�Yv�X�R�w-��3�m��g<������puY��f��M��"�Ѩ)sBB&��ۂMJ�)��k�H˧W\Ꞇi��r�r����H�5QXٜh��װC/7oQ�"gBKva�U;�4O��������Uɍn��j	�2#�9���l�pu��';^1����gl�!�1�����hvW-���*w4f�tHȑ{ڏ���J��'M�zU��\�����u	C�m��Y	2���x���R�z]V��+���oe��m���w��rV�|ଓ�j�x��㫰�5ʣ[��j�K#ON��wI��{V_����Bl�*�q"��e
�vv���s�p�Ђ�����+�&�:��������G���D��5���;���&Ùz��']�rxqF��������n���fHy-�ӫ�Pu��fL1�2���^\�O�ٺ��i�N�ه�k�ͭ�b$�Y��5�*����Z����5��:+����<�wr�R~ǧq<�Y���^�V�M�S��C%��A�p�GQ{�k:�]��fye��{�PȜ���F�]a�9V��Φ8�Sy:\��.�|�篮���c�y:KKrG�&Y[�r���*�E�Fn�7�ɽBc�����։��ʂ��͗`iG����9n��b^[�	,`��!*�g1��8�9F�fe_p�S�+Z��h'���Ѧ51�U/��K���+0�"h��R,�FÌ�t5�qīcc�L��ۺ�}�כ��[���)D^��Pɡ]^���^5/��1�Ux�=�l<�}ȴ:��N9���2)+�{y8��c����Yҍ��z�=}������M=Ye��9;��ν�����|A%˛ؠ��;�����":q��g\6�,uyyb�l��T�,��9�#�q�;WW�a��,`��������;ə�=�%cDD��,�=�M��A�݋[h7cw/�
mJ��	��2�W��V��>�,��Qf��լ��nζ�y!���{ݽ*U�uqJM;�1:ӏ#�C���a��|��sr�	�]Dq�*�7 (�ɗB�FM\1�\"��ܪ�wA�]LwN�D��`��i�LF�ݙ
�X4���|�8+n���kd����7S�b��I��h��Z�2&ޙ�`�fi�k!�
��W�x�Z��c�m�{�̵=9�҄t��Ï���|�+��"둭��gLS�Q|���oV8���kEvQ��jQ[ �+7q�J',Z���nr�&�H�J�%䬮���$��`����������I��<�#E�2�T�/D7
���;wmڜ[��Y��7�����Q&,!\.疫�U�w�ݦ��â���u��,�V'�v��S�=�H���9}s7�쑱�B���fci���Ow�J��k'J����Q�/�R![+���rv�"�Q�[��r��}���I��0B��NE���l)�ˋ
����4� �nb`�%��/E�����1���Ȳ�&+�;%jW'F"\�5��b1�x ��^�%������xɵ.��y�Ƿ����e8���.��׷$7Y���VՁp��&6��yj��73sw��R:�]���ZK�1�׬k��k�y:�|o6\bp�֝����L��^k;�`������]��4 �&�M�3��z���I��vr�C���E!ƣ�wz��_�yV1�<�o4�^A�K6v��,fCh��I� �),c�s}X�ۏ8�z3a����G�s+l��ۋL��y`��@��5�.C���H�]3A�TX8��LaƓ��/fNv�[�Ft��V�e��wV���BV_�mk/o9���]Ԣ)J�r�M�9Y�c�n�'����d.��S�I��XO&�:�m7�g:�EP��}UMȕMÆ�a:���e��X9�8�//�f��s�G�KT�{�$Іgad0]f�P�XJ��\�vY��bC�]=�h��4���!���{�eŅ�����������)�M�,��k)���　t�6T��eXPf,���Y'<y:u��gK��B��ai�y��yǰj�s�8#���v���;�3mL2�کHŘ���9f�֝�4� ^�8�������9�i���h=o�}l%�(n�ݫ��Т�o%w5��!�իU����ʫ:U�U�b"�u�KV;s�#+0�ǁ��kUZ�@�	�^Ao��Q������\�m�P��K�p=nY��b$�ewgR� �{�V�VC"��ݒ�/IvQ
��ׯl
K��o��F�ʝ��s��^�4\~���n�U�D�e[�!+��q�Z� �f�m�ݵSa�1�p,n_�Lh��+�m��K�dV�KM˱��{"��uu���׮�ac]D;�SR=\�gF��=�Ҁ�;�,Θ3xA[|�m^�3Y/*� �JT��R"�2E�V^gF	�C��ޣ�s��	!5��͒V�E�58���
G3sa�B���_���ߪi��]v��-�9�U3
LN�[�X�
�XY�����jŬ��:i��%d���,��L%���ގ��R��S��{�u���U+)ݜ�)��XT`ԍmi����I�-t�b�X��jWzx޲/�apH�&��*޼���ƺi�s7j^��U�ˌV&��w�����o�9�&������ќ�f԰��\�+�m�Q ھ멎Sd�z�67�c��U�F1�I�",����7�E��>Ɋ۪i7�dRD�1ζ���[���[5���Ϝ]H
���8t#l�4D��j�d�$��0�v�<5m��ح6�Ǧ�kE�����{Jc��q$���o)�-�X���l�g56�J*\,�WI���m�c{E�۸*��� }�T)d�c1�T�v\N쳶�*�:�����v(�f>�������@QyW*	_wv���KB1�[Sy$\Y13R�i�Ɇ��Kh���g16д݅b�p'��ϔM��
��d��$0���^�����f�2+��R�y�a��C�8�*�pΉ�����v��!,�,�$!Hզ��2��⥡hm�J��� �(:�=U3��q�U�FSG-�7��8��ZDn^hV��Y�\/7��rLG�w�qԾ�C��9p�]�}��3�{���=��]�p��h*�s����;�.6KX"��[�
zUi�y���.LԘ���E��Uǋ��=�׻;��oj�,E׉��P'�WmY"Ulo�6{I�u�;е�=�d��Ku�Sl	�;Kx0#31���c������\�}��N�q�(��\�k�%��3VM���sd7������X����Hw%��j�綍c�x�xn�M[�6(������H�>�)Ko�OP.�����s+r
1Й]cz{I�y�7�#r�n"���F��W��*��V���L�v��)M+f��Ta(�
��ڹw�c��A�nw3ע:�FA��ʤ��Z����485��պN,��W�tu�k�-ͤ<���4�]��JԣRv�sް�m)�۴�8�N��fI��pC[�ud��ks����Cp�o�l4���DY���$/����7Y����	y�Ժ�:�vK�5�e����l�8��sn���L;��/n`��5��c����qp�^cKATe�l�b�tj���@��|����+���3i�G�N�lv���W�D*�-m������!�'f:�I x���'��c��IR͠RT��ᒚ�j�a��2�V	݃�.�խ������xWX��T[�v*3P�����4�޸��^Ɓ��%j�=����~�}h]瞉1b�ղ��Z�!�
�{�л�'ݛ(��M���M��͗�q��$���{l-9[�g]�>����Ґ7\�����[����U��j	�#U�4���dہV���z����ڼ��z�r\,� �t���2i�v�F9�[rཽu�j���k+����^��o:�Eɝ�,�x1��6�aM���7����I��{�/2�	�y��g\/y��Oo*d��##�Mm����r���}���.��#s��+A��gu����	8	����9���f��!P�57SNѽ���Z26^�L�����ɘuP)(�r�u��ԇ%���p�wl��Wb<��cm�p�R�o.��0�X;�jK.i����-�Ux#��/z�`�7R�۬��c��֚�1��#꼽�G;���!҅�J��kr6����za�?M�㖖�!^�U<I��C��_����U�Fj����98^aɷ4M�{YnhꉕOm4�F��Aδ����z��j�z����*j�>7��	Y��姉��ɪH���)͖�4�I�F���f]�u�c-�z��h�hb��\zګ�,=��5�����Ց��q^�i��"\�����7CSF��+^k_y�JEµ���TK0� 5e���2��Us����.�P�A�n�-l��m�D]NܙV���+�-��5Y����ʪ�h;���lM��m��m�0t�]��N�M�miN3)�պ#6vM(.�sMMa���ښ���x�N<��� E�{�ê�A�U�}^L�H��~CyϾ	}�q^�{��|�Ϝ�^_%�ϼ�B���ݕ��>s]��`t��U��T�}���� |��|U�s�W�'�9|�~y�������������矜)ZG��oYOP���;}������G�b~H����9ǒ��}�{��/�;�����<E|�g��S� ~�����䇨�{8x��9�q�x׬���>�[{�ߘ����O�>��/���^��}ޥ7�r�s�C�G����SԚ��x{�*W}aK�WÝ�v�>z��j���TDG�q�g��D?��������?����O���"�#��D���C����k��������s׿^�z������$Ÿ��(+�yx/Y9�^/L���qK@���6\u�m��}���u��љ�\�#���8��!� ��e3�E�� }����U�4�����\7.��L��f�唚����U���<s���R�{Ӟ���<y�S5u"��W� �^��ܨ�j)�b�v
�;�v�9ne�I��ΰT��D�Y���V����=���U�i�xٔ/�`�O��RT��O�;�,C_������p>dr,�pٲ.��/)�u�C8� !���̃o({�Ǡ	iw�	��/,v�k/���Q�W�Oz�	�;��mk���$-���Œ*8d�y.�Իc`����2�P�c<9�W�^6.�t(��-i�9�nBYYWag�]B �k���Y�Q��1��i����[yx��T��vj��pPM�X07�΢�n���V��+@R�gm�0WT���[fS�f�X@�����j��j3*�rTZ�$s�ᝤ����D���� *�!�(�#�¬oA]����!.*	��%�$W��}�4�;�Mʪ[���͂ogt"6cy���|�,�%eg%d�dUu{�&a畝���1�l5S¤ܰǪuꍘnl:�q*��s��]�Af��\v Е{�����*��KFtg�{�J��ȞvA6�͏�����>��=z�����?��^�~�_ǯ^�z��ףׯ^�z��ׯG�^�z��ׯ^�z�^�z����׮z��ׯ^��^�z��ׯ_�Y�ׯ^�z�z��ǯ^�z����׮z��ׯ^�޽z��ׯ^�}=z���ׯ^�z�z���ǯ^�x��ׯ^�޽z�^�~=z����ׯ^�z����=z��ׯ��^�|z��ׯ�^�z�����=z��ׯ_�G�^�z��ׯ^�^�z��ׯǯ\��ׯ_�z����׮z��ׯ^��^�z�����=z=z��ׯ^��sׯ^�|||||z���z��ׯ^�~�z��^�z����ׯ^�z��ׯ_o^�ׯ^�z������ׯ^�z����ף��ĺ��ߪ�Q�O��j�؝`5(�{�G|ư\���� VZ��u�������#x���-d�wz�cX��}^q�����I��q�w�/�(��&��J#N�)ۂYHd�xq�d%�H:��{���+�4i������N�\:�lbl���H���q\ⲋ��$ʲ�E��o%ذ�=���ŵ�s꾿U[�dt9v��C����m��z���Jo*\Z��p8��D��)��w���9�ѧWOB.�\y�fJ]��kS{+�GK�-��H�<���`�-�zخ�����/z��w:��'X��C)��;-���ҾQՃVFA�S�3C�W�u��'�lZ�%ug��v�h0|/�1SHs�Z�F(-���d��w�l��V�-��S�p�e�\�V��J�W����;�E!���*@J;+mdk�Ú]����
ש��sBK_�̪���춏\����w��T傖����j�]^+�u�>��]0嚰x�8�ص��N��v�r�gd,B{d (����CE+fL�^�un���)C;����ŝ%z��u�/�2®b�	��Ԥ��ox>��+j��9e�o&��x��*ޔ���n�F�GV�ް���l�,�`,�#9�y�5bL��j�ukG��>y�o/\���]��s�������ׯ_�z����ׯ^�}=z���ׯ^�z�z���ǯ^�z����׮z��ׯ^�޽z��ׯ^�=z����ׯ\��ׯ^�~=z��^�z����׬��ׯ^�z�z���z��ׯ_�G�^�z��ׯ^�^�z��ׯ_�Y�ׯ^�z�z��ǯ^�z���ׯ_O^�sׯ^�z���z��ׯ^�z�z�^�z����ׯ^=z������ׯ_�z��ׯ^�z�z���z��ׯׯ\��ׯ^���z���ׯ^�}=z���ׯ^�|z��ׯ��Y�ׯ_O������ǯ^�z����׮z��ׯ^�z�z�^�z��ׯǯ\��ׯ^���z���ׯ^�}=z����w����>��6i#c�^5����m�-�Oq��T��s77K=�^V�s"{��:�u֛�k��.2gMf���ܫ�W�r�Or�� rjיf�ծ�Mh�v솫/jwS���2����4�U�f�k�[@ܲ%���OG_uf�wҟ�{���x����T�9UP@J'u�LCJ'��
|z��\z�)X;]�'��kH�y�|�y�(�8� 5n��V�-ǫV�t1vM��=6E�Ijv�����R����a2�@�	����9�����"�VV�:W#o�T��Vgj��������w9�f�#hu'�V�U�SB���.-n\!�y�3�{��6�X�\������K˂f�(}����T��bT=dml�k�oO
�C79��bsq�,����VV�����K�es2�֘?|9���KۘFZ}��ХHf,����s2�gb����2Bt̐�,[{ä�o'=���X��b�n�x�dc�$D�b�:;:��q'˘�k�8�7�a*��'�N�-�\��|�ܭ̥T�gU����2�ꁞTl��e�s����\�j��߮�|T�K>����V�}�sN��#�w)�e�8%�B�]-]�fӇM�9U�r�q�6b����F�ٔ�P�}!�]��{�f�����
i��>��VRѳ����S8��"7)������u����bze��dU�ˆ�s�Ū���E�Zqӹ)��ڼ��8+o5F:���6���©ըl	bi�$)���(Y���7x݄i��\�0��6-�&e7�}qTJ�
m�Lk��{�s��k���5ޗ�{GNH��u�s�"�Y��ENs�.b���f*�D�]��f��u%�v-�4J{o������g�r��έ]~�'Bn��(Q���݄���~���s�;.�;0��4�m�qϷx���n�Y����Z���*n�\"�I�-=9���T5J3/J�sHz�Q�D5����hz�)Y����q�Z-C��5��р�eӺ&Tr\���Z�r�Bkp����k���(�=
��r�8�u�]:��8�-ZI9�&V�7������ꪙ>��tr�l����akbG�vη��w��F�Y5X6�TI�����O[W�59�����;�;W�)��'����}�WV�E<Q�GS.���t��o$Ǌm�sv���d�ר+J{�n����8q��E�bM-�9��axr��K0�%�����`���qYd4ekIH�Jb��S	ٴ%o�7�f7�gٴ3O*/�.f@�v;��ʑ��f����@6 2�n���e�廦�;V2�{�G}�-��K����-I����*ժn0�{�3%��f�t�mS���:�r 	?���K��r'%���՘,����zK.��wz�7jb2��)T�R�漭ۗqai턴1z��Y棷؄�km;��Cf�]�P��8erT�௥aȰ_O2��v�k=7�����2K�ܓv9n�RzR*fe��SoP���6�5.��ܧ��}pW��;(�����Dn_
nD8��P ҧ`L�~F�jʻ��N

|�٭�kcrCc�q�rS���7�R*�)��.�u��p�WR���q�i�ћ��0~f�.ZR�pt׻s{�uXY���+ʝaV��Q�w�)9W��z���1o*�c[P�z(�j�ۆ�y�<\��ٷz���F ���wݥlL�i���e֪2���ax6㻷A�V��m5�2��[O&�e�>7����%Ec��4�.������v��9¶S��bغ+tI�7J���[oD��@�ݺf�M��-f��,QUs�gX� X�����X��Koiof\������/ �����Og� ���!`c��*����9�ƘxVic
R�b�јbl�.��/��G�����.��<��|��
��B� g!4xL�P��ALq\>�J����jQ�c�C�$��������
_M��ݵb�)o��3�'|�%F�;&st͍؍n�W��䛡��+�F��V����/\��.4"���S���o.3cEF�	�Y�N�q�(#�;1%;g��g{�11)D��@�G'��b���uS�]��g���1��~��-�^)l��Q�E>|�FS�f+o��'JW��]�⧥�8�Zԣ�ЎB�V��B�ekW��k�����[b�U�5m4C;���ev���h]A���]���A�k2���a��3�5�������c�/:��M��ܕ;t�U��s²c|��2�u�ki��VРt�j�uQR�G����יޛ\2`�)靫��D�o���q�B�Wt�J���5y�=6���VƦ�wJк�ݜ�K���\�:j�N��v��\5�c�L����P&ܒ��l8c}5
�iW��s�b�$��#ӧ$��;ʜ������JD�8�I�y��f�1p�.'|�S�^Զ	\����sYo���_n�\*Ai���T����;Mwݮ��ڝ��$��� Sy��}v�]���톣HN-�p{�	�ʰTڀv�+n+2��L����k�#Q1QC�M:�;Zh��H㗚\cQ���n���{tx����ۥ�y�C%l�������]bBg	��vP��UB�,�
9Ml��c����Y���@Θ��Z�_p}9̃�:��&��z�z�8��}���WX��^��!�L��v���zټ�[4aÒgs<����kip��N�U�ܣ��s#}��+p`�N��x����K��3qd7֡6���c{����6c�m���vvˠfu9ݼ�-�]A&�Z�f�����i�D�ف*	V3 �Pe�:�q��VD�Wš=�']�̼�W��m_�c������e�{�2���kz�G}W4�����d��[���6�>��ʔ�Ih��T@}�2ӊ�a�c�V��;��H;ו�]��jPpM�(�V�V��_:+�Z���~=�G�.�B�1K�t�^�-K�gU��Raᕃ�-f�1�59}���D&��n�֜݁�r�&#O��Mwm��{&nG����wI2�>�gY��i9�ۜ�p`�������p:~��,�9qG($��in-:��j�˼:����;{(Q=2��$�Hn���Sd[���6Ww`ޢ�e�v[��h܂���=ȩ��u�V�ұ�e�超�4���PM�J�)�l��H$���\�֌�����ߗtX�8�.,�K�LKշ��tm*vݍLe蘽O�]b�S�3�i��
7m�롺fU�e�Q��ճ�kw��aɪ��{8&0J���ޮ���z�A�L˺�&�l3��T���fYі�l%#��a�N�\�䏪�^ј3>mR.�T�J�V3M���f%��)N������&�8�Y�볠Hn�6��P;T�&��u��S�s��!�aa�a,�S	�|��s��p��)��},B	(at5���n�fpv�N��:��s�#�%mZh��2�(t�Xv�3��R���c6�j�� X����#��Cʰ�:�/�'\VB}�i�g/[pB4^d�&��W|��&.��ar�3��坋���Q�HtL3�P���9i�z<��	��x��h�R�U24�i̲\VI��\w�C�Г5�b�1�vhÒr�C��4̂Ό��ڈ�"���\�^���cFd����9��^��Iw��Œ�����U��7�`;:��ıwh�wc�;�m���� �ytx��<8�-�.6N�wS�ƙ9]}y�zgc�۩d<��9n�뺛7�Ä��Ck���*��R��3���)�%Crn��3Lf�\�ty+\֮�i.อs%�l�oY}T����]`;\^Zj^���+I��2����}�;4�Ow��Զ��Sr0ɘ�pn�y�dƸp��S��Q!����l���f<<]M�h�uamM���b�.�\ ��e��N�U�B��tF�;�x���(��o��3K':�S7d;Y˳��spT�ӆ�v4�;���"{��w�٭���jʑ�J�e9CC9Ovu�ǫ�Ռw�:��=��; �Yנ?W���dݧcr+̂��:��FN��4�j�wEҜi��n���U{�n�9{7���t�ʏS�C���'p,\p/_id����Ϡ�<�r�3�wd���&���L���.�XiA��rV[u��x���g1�淊A�۾�nt9�u!����x������{���E�5�]����F���U�C�㥃�I#�����#r�F�r3L�v��ckL\�8��)e��.�PP�<���iY��4m΁fU�Q��x�����s<�&��$�Y�|1D�n$;�~�����$�%:�shY��t�J[�w�#5�I�z'f࡜�*39�یoU��Zrn_�a��*C*�pw�q�	�ʯQ�Pl�a]z�?os�zr�yg1��ܸ����Y�N�B`��|9*���xU�{�~�уH�pYD�F�ݝg,�6��^;Xňߪ�Xz��bQ�|�+.���G>�ycc�ݼx"l�x��-uI(�I�x4�,7;�*�@]65U�ٞ�5�]�3��6�C�`�Fk��L�ǳ�Dz2�5ۅ:�%��U�S�$��B�ף`u�)۞�'��kT�̠��w��������r����m�J��T�lw[�-a0�s:���z]W����9놠��:��+-�I?�T�!aQ�
��¸;��#X'>�s���i�VL��W�\e��J����'�L[�φԸ*�$1���U{O'�Zv���b��z+bV�V��`y��������2����<�F��fHΖ��:[yX�D�q�ަ鞇p��J����ڇ����]��&�=x��׮=���u!ڳ� ��t#�u���
�#��^�+h�+�k�p;��M^�)��`5)��3N1�|�0��r _s'��g'+1����Y4e������9�0�C��{d�Uo\��՞�nʡB#$��nb����_Q,^���쉋�D/W�w�u�ݳB��
�C��ُ�h"�5WJ��]��o(Yu��8ڎX��T>�F�!im�4@�P�<����:}�}}��9�t����( *�}����������������Ԯo��������m�ny�y�rD6\D$R
8�)qH���RF�I�������L!��� ��B�(�S!�#�/���`�[�"Q��N�tS!��P�~Nщ� -��d3	(f�Pl��-��J�4�TJ�I���iB���Y� �D6�4U[iF&�����l�!t�l%G�SO�`��RP�i��fB��F�.�h���8�4m��ӂ?��D�`��H��A `SaR��TCL�_��ɢ�r2	A��4���O��;r~~����u�o��^[	k�����Ȟv��v�t������*P��u`ŗ�)��oxn��`4�-���7���Ҥ�2��j�<	8�fұ*\Ø^��*��DڧĽJ�z�w�m��6q�j�ܻ,xvfU�94�Rk��I���C�Fq�qf��+�݊Ǎ�+�m�7Y��[Bl|0ڋ�ne��ٶ��nd23��ǞA;M��X�`�m��o��NrqRas�K9q���d	��1b�� ^0�O��׬e�H��ۧ�l_Q�3�W�g%GMJ|[ ec�v��֎��ԖJux60m9p��Nո�����4n�Dy�Z�C�b+I�H4�3,>Fs�w,Q���0�P�8M�'C��CrIE���ǁq��Q���\Yt�-��i.�͆vf�hl�Q,E/���� ɽ���6rK�.�W���B�n�E6'�waWEֳN�F�WKM 锯c���.+�G�좔f$�Q���W%u-�ҷb��t0#�EcՒ�����nv��}�L��bK�����̀Xc*���F�#]2��a
`����4'^"&�Æ�m��i���ffm�o�k�b�R5H��"@�pb8��#8ZlH�a��H����JFH��>�E�$ ��(�����
��d¢f(��`��,F�i��(E �Ų�f(��,�m�L�CaL�#�}���I�6�K�H4TC���J1)�E��g�܁���%�"8�i�DT���ߓ� ���>m5�F�M�i�\@�_H���D��D�}@���E���h�c�(ĸ�E�H�Q��f(	�F��R�RM W�Fq�/�m�dI/�q�����	0Ag�$�2b�qD��Jm��(�L����*HYd@�� �B6�tESR@�N}!�3 a3t�"JO_l$��Q5�j�0 Qj8�$$* �dF�q�A�(Q)�,�r*T�$�f$m�Td��ed	�u"� S����S���(A��Ċ$��H���:t�40��a�HL�f)->q�#O��$؃ֹ�o8oG�sj��&�@��#�iH�h�O������?_ǯǯY�ׯ^�z���z��ׯ�����_��p|>ڀ�#��<��=Ɨ�RRhѶ�-9�oo��������=z��ׯ^�^�^�z�����������Q��<�"/�9�$���z�TD$ɠ�:LA�Jm�V�����ϐ󘣀�W�'�F�*��4KN���4��4��ɠ�rJ�14���f��<��s̴����pj��3I�9�<�J\��b-j)�{U�.�\�z�9�C����h�Zl�M� 4�y�ݘ��*��I���S^l��s�< �d�i��G�ΌT~ڨ�3�c�.A�y�_0j�QF*��ֶ�lo9�y�rG�*8ZBɠ�Gͪ9���랽^x��m4��G7�jG͵ks|�_=!¹Dj�"�����Nk��.5�$(�A����iHX�6�0!)�[A���Ƞ$��M"��$H��}�.���BM7cK�ky�6-�pvV�2Ex�՜���w6~w�����j�QI"�f`F#�FJB�"6��(6h�Tq�[�4���
DYq�0�	`�cH�#,BXe��&�lD�M��L%
��#A4�a�^k�^F+�r�.s���+~<fc�~r���E9�91�Ĳl(�rM�k�e���
A	�"u6�9M�����Bl߶��O���7�]}�s}�������c&&L{v��^�����g�l
��F��r�#w[��X�+7���"����o:���f�³�N}�����+@��}����z����1Qo���00��BU�w��������ޤ�S���?���l2�y��͌>|�����_���W�����;Ԫ��q��ZϏA9뽋&�A�ͨ긞�����8��ǎ*�^SoQ����j~��u\+iî\ZA�9����8�i۩�z�>+MZjj5tm*�x���vD�|�e$>�ML����y�����[���MT >S���W���}{�L;[�����%�G:�9��]9���Vk������g��7��>�q�����O�<�T���.,�A�t5U�P�i��d��s���˫��]w2ٝcJ�C)����%u0��u��ȝ�[B����QWC{�����T� ���T�<D=ښ��vY�5��}�&◚�M���k�O�t����z��Z�����6t�u����⯷�.΍������ �s���Z�� �����P�����p���in��O0cx;T��W��#!����ǯ�a<ޜd����vZ�nF�uW T�Oa��>F-�9ʂ(�q���߯���$�\�����4�����ݑ��ds��b�e<���צ�����`�o���X�{nI]��\g���"��m���Wǋ�t�һ>�/�,)���z�8���%�+�q)ZǪ�s\p}��&&1Y5���f2�D��h�8gwbs��X���`L�?���RR���LZ�����Gr]�MvZ*�(s�����2/� :��^�}�v��E��l����M6�K{]��vo�w3����Ȳ�,>-P��V�NH�^����ю~�҉�����b��7�r��f*������U ����}�֛T.p��n�u��cxh���-����&��85��e��Dfꠎ�,���|Ο�v��Z.Ж	m�gc�KZ�5�Ӈl]]&��%4��3}&W.�K��eoT��Zz-#N�`�#��?O�Bn�d����xq��� �=�5v�	~��d�j������3����Y��[�Y=D���;>�6o�ȡ��\��Ǎ:v�~�G"jkJD	go��81t"�
��Q0�rxgUE��nw��Y����z쪽���̿�fD%�|8���g��ΐl��K���ƽ�}OI Ξ���g�* {��\�<�,_t�TOqV�;���.��d��^V���]�����=����==�(T8G�QW��El<r9�=|�_w�Q8����G�/g�l�v4X��Ä�N�Y�\M%T�N����v#պ���D���
&~w
���q��L���}M�?eAU��[�J���Yhc�gt�$�����O`��퉻��F�W=e��oڴ5h�tg�4@'�F�z�s�(� �v��bj�ry��X�����3#�i�a���m���B.d;r��J9�N�����α7:�Gi�:��[�;��-M/���Z3�~���^۲���bһ�`��N��]
�[�0*�C~��-�A���-EUֽ+Z��NUZ);�T	ElO���?TK��od&�-��(w�um�g���U��}�y�uP{6B�u�������ۉ�d��j�GD0�L�ީ�=�q��*��9���L��W]i�z���8fm��Z�d�e���NՓ���3�oٲ{F�Eb��%�\X{;��#��x5,��z;����7���T����֢Ϻ_�:�W������(�ڠ�}S����'C���L6��l��\u�Vڸ6��}���ߧq�Y�����SMb��}�;e�&J�ӷ����ݓ��D��������}�M��ڏ���X!�aӼ�h�������o�Ү6w &װ5���W�n��G�^����zf�-L(��#;z{5̂wn�<p�ƌ����*�~�|�^�e������>oX
��~�]}���pk��`oR�=N�r�5��� u�.a�S�n���p��1l�.-��q���{�G��w�m_.��,iK��h���h�}mR�8MvF��-L]�A�`�b������k;�h�H���Ԧ�z�e(�����Z67.ީx��fmg���`�dBM X�\��nŽ0p�,�QT�+@ԷPJe*TMfT��I���Z ���?���*s�B}�+�+���*�9�V����{�+�7:{)Of�n}���87�e�c���S5��E��c�����ם�+z���t��wB��4�z���}���z�|�*'cٽ���Z�u�m����������_(�~���Y�$�+q�� }%��Xy�&�Q����`�o�'�{ۦ��u^�u���n�ɛ��+�������KN@���h��m_���X������B}����;����NQ��4�Q��D�}�Me��l��1ZXČ�:Et�NY8�[�������*���4�� a܉��s�F����� �*�����0J����]�u�ޗx�v�`����|G��G��V�Z=9�lN�ǴE�5n`M�_l5��f
G��,�}�J[ػp��j~�M���5�ٗo�Ge�Es6B30V9~SJ�J�'}%��E����ˌ]�Q�I��Id���¤K�c@<�9��E�P��4�H:��>YP��Eɤ|��S� �γ��ٺ�A ��:��WmM�X�r�b��g<�~��rΤ�3+fΙ��;�����cM�ҍ�.J&�����?lGsw��dWHw�Ñ-��k{�e%�V��)tE(tvc���f1��|�>�\�2o�ښ��[��<��^_[��� }b)�E�������!ow%����=hhE�20�$Ci Sz��gy��ߧ�,�El�W�_�pm���9���R�r��'��EJq}�sd��\�u}L����[�e���97���|�+���W_`����[�c��dc���gin�ey�^?U{ ��'��U��we���77 ��?�DOLCǒ;�u)�^����߁���'*�6�G��銙���~�[��9	!MV*\5�ܦ�1t�?U���O���-�%oW�߸z��z��Y��b�I!��P[�Q���ت���{��avCWQ75�N��ʑ��Ys��V�����t�n(�gt��`�H�eu�0��.䦱���)����V{�=��
��Id[��Ҧ�{�ëD�YL�E�ܥxn#f�L�p%3;E�٤�W6M���e��6���p~ߧ���M�a�pf����W����I���hw�*��y����2s�z�'v���^�F5���p��\|8��	���'�j�zd��i=�UG�����co��X�Ȍ�֥�;�l��1|8݁U�/���^5h�}5�6/.�ge��"�Fuxv[`��	=�f���M�~�y�c��;��zT&��#�
��&>Ί�x2���v}=d���U���nk���_h�mZ;��sf�C[�;"8lS����w���_K���%��m�ZY]��t�4g��`���� 8�vU��R����*��Z���C�/yv澓��z#���0+��d�^z�/f��ޯ��MǺ��h=x:�㜫�	�"cW۝�ϡ��� ��4�������}���Z�J�kڀ"x�L3�EI��,;,. ��`N�9ד������EE����J��Uٍ��t6�kz��I����N1�}X�3E�[pE[�^�=)˰���:��φ!Sҩ��� !��|(��Z��Y��d���n��1h�}-Ѱkz޸���w�hk[�V����YҒ����_6%�챜�7�<�R�B����y�j�/{��.�Fi��"�u�N�:�c�c "o���Eۃ�z�C;������>����~t�~�}d�m���5=�qv����+]n��
�cý����~@���\W���˟?JH,���.�Jn��Fw}3JN��wՕ~�Pc�/h�bx���+���7U]�O�/ ����戉�{c���X}E���Ԙ�o�V��>wy�=�F���O_`y�V��+Y�����we��^z}	��2��.���$����v��4*�@==[p���{u���}��f��}�l�o,�&�+�'����|�!����tWNT#�
�Q�9�%]�b���=�s�#DVT
���}�v�׻]�n����V���c��vM.0U9��7-9������gg�����x�b���ţۗ��w
�`�-wz��B^pô�h6��p���{e���y���]�	ٚ��V�
[�a���=]������� ��5m�,��'-�k�޸�a"����u�N�THCcz�Q�����ڦ�e�䴓�6J�������6�[׳����*{�s��(.o�gS�x�"n����ޥd��y�g����6&f���ӿ;�[�4��U��7Ğ�<n�\�r���sq�}�L������ͷ�k�`6鼭���gm\sŅ8��5�#��	��u�*Z:�6mL�N�we>�a��'c�{A�;e�Dx�L[V�\��|gn��+�텵�q���Q��^� >;��ʓn<��k��Xy���x�e��m�뿪z:ƣ�/���1��F�}��W����#t	�|���wMN�[ݴ�t.z٨����9���D뿄��1_Wk����gB���2�V��n/�N*��(�C���}K�k8�V���ODu��~��v@� �>{�.�����*V�Op���v{fj`�U:���&�OQ�i�zj�j?�� ��8ؓ_y_��� ��<g:7��幒��!9�U[3��cb�S��QHGF�k�+�s�Ռ�h�Y�#sf�W�=���+>�şc�>ttV�_̋(���r�$��\p7/0$w��HJû�̠���S�����e���%͔�d#X].���G�f���ZzU�迧��~EkM-j"n����/͡
���N�z�?}�+.��_�7\���ι�e�y���z�^bN��5P���h�G8q���r���~Ɍ��o��e��Q=˳�b��nx�����>q2���q�$��D8D�kR���wuJ�ϻb����#�+��2�m�e}6#��F�u9�9Nj=�k�h�#�������ȭ��4��m�t����E���1����U�3����0���:�ЯV�.c!����M�jȫ㉢3p�yݷ�V|�?�o�^�_�sa�K���$�d�VV�5T'8���}'ZB^��
���.���hv��1h[��6�����V*a>F��E��G����ut�I�H�(7�!�_�~אs��\t�36yF��L�9%�����kׅ��sU�I�h�U+���J~�����b���H�L��Q�:0\6�)WX��a�X׮�mm۾�V�HQ��O��*�]c}QA�đ�8������c{�Hᕯ����y�:Զf����J�g�˷�Y�]�2>s,dH9�y7E�X��W�j��@O#�ɍ��P��g�m�::/kQx�u6��κ�/�敶G@��Q�l���6��%f	CQoe6�y.��E�X7|�f
\�jݛ���5����z-P"�vws����G�l���W�`�p�d�=��g"�ۡ�͌���λ�lBJ����O�٫u�����	��G%�W\p6�,y(j�x5����9�4���j�����3J&� �_\Q�f>��p�j�BS��e��.��K��G���Nc#yR��Z�@���.�]f���a��v�{��9�yOYA�C1��\�λ��x����<*g5�#�aGu�m�i�7��ge�rSأ9�v��{qj���pjv7�ݲ�m��K��<��;�F�����a�mfU�ޗ�Ngs@�w;Z{x��ް3��at˶uj�̀SX6�zՊ�af��Ub�2֦^j[Gjr�-\��*om�m��x,�8����)�����ǳ��mŨ��(�m:�g^!#�t.��io3�MW#�%K5Ù��[p[7�ٖkJ��Ծ�̃;cS���"M�& M�P�� lU�5� �T�-�"؇*Ĳ��a�5(#,
#L:���)�I	[�B�j�p��{�o+��$i)Fy	��%3��6s*!��U����/���K��8L�'{Y��%9i������a
���\F�<��%�ƶd���
��>nlen��u`�o8�0�}���c2��t��ͼ�����m�t�W��i��+p�����z�1���fWD]Y�Z�!�H��	��X1#�I��,��	V�飀ȯ+O1s̼��@�&N�ݺ���lT�2H�<�Ѵ�y�-�Ʒ��L�����Y��2���^��2���z��������p쳭p�O�u�`<�]t�/n�4V
���o��e��aѱD�����4r0g�&T����:c�g2�:e���Օ��	[�*%�OE��WXAL�*�餶B0�u3YW`��.���Q,f��eܾ�[9G�\����C��ҹ�z]�.mek�o�Uچ�eR���FX���Y�p�z�C6N����՛-�*>�`��H���3�����%$��M�-���E���ȸ�����b�`�zE��[+V�̧3�8���C 9�*�۷�̔���@N�ֵ��|����%;հ�3(��r�w��/���':�Y����XJv#�0�n��qCD�I����t-aj��拂�z�m=}�U���m9��������C;0o'p#Z%?#U^�����[�9�%y��6F9�ֶ�c�p���Հ�m�g8�6GQ�בǀk\g�����_������=�����������Ǐ=�~s쁛����dc��.�66<ߜ�� �p���;	�j���Lw k���dy\+	�4y��Q2>Z��ӱ���_\�g���������z�랽z�����~����?��Ǐ?���#� �Y�#����s�n5sQ���0E��|���h�9���z�&/Q���[՟4U�6�-W�8r<������yss{����=���ߧ�?���\��s9�U�֋�����j�f��iP�� _ H��!��"M��l��b!G�F0;k�g�y�S�"�y��� �~��D��,��ԖC�J!Ӽ�#�7��&�|�r��G�<�m뇖�ϐz�sS�S�}�燉����yc��;gN#E˞c�g�>�=x�X|�%�լQ�^r�[y�\���5l����9&�nc{6���mmV�Q�\��}��ש�8�����gC���d�$Ɍnm�{��:�HƵ*dʹ��mY��;{n���_��x���z��uU���+Cn�_� �c��qZ�ϰ�����Fy���G��s��hz���~ڵS^�&�-j�}>�#d��wB�fÙ#׆�f�����jV[���Q�WZ"K3������1�u�nC�J h�f�X���ɓ=8܎O��.�"��hW�A����H�k-�V��5��G��C��#"'z&&� V�k�,�S���Dl����9��^&E�)%�Ζ��ڇ����fY������>t�b�����
�ك�u���&6�;/[αU�pOB�.C�ns��T�d��%�����ҮD��0��0~@���Pkc�Y�0��d��6_H�a�S�y�����L�=�O S���SiP����aċ�v\��x;���SK��:ċمG7gi�C1d ��`;��=��;�S��Z����*����[@咶���qͶ�z��e�z]�G�3�O�J����ɘ�[�6�Ջ|���8�b�PdO���e-:��W�sFE���bf<�&�C/�ь%:��	r�}o�EwH���E����e�x���N�/2�Y6�3P)�6tȢg(e���
:lS��dX\���>�ܣ��y�`�E^�~�f���s0�U�	=��U&��ݣ����Y��޸^�I2��])�r�7�Ҷ&�ݩ�9���o6x��^�8������㧠������B�`6ǼV�v����q�GW������皻!��j�����B�۴=��gG�u��=8��x�xk��0v��o��$1���/<�1�;V����R��WS�4[!�UR[�(�`!=�>�y���Hq:ŧ��ΰl����z6h^^.#�Ϗ,���(c�E�5H�����M7H��{>h�m���c!�P.��O&|-:j����{^L��ff!�ݻ�]�P���q��J���m7#��?q�a�f@�㺲��w��xC�E����H|d��"wJ����m_(,/���3[r��la�l�x��ZQ�%Q���}��C�� ;�X��/���И��Y��s��a�g�+�/�HM��Oa|�ͽ�z�˄VO3R�2Q�o�3P�G�@Q"u��x>9O�^�ų�@��O�^�.�Se!�́�@�/#[��3���t�dK���w�r�oC	0����
�^����L��.�f�[��ӣ!�ӹK�<ҋc��:�1�2סf})���ĶEu�U�)�z!��ST%t����o��.��k��w�F���^K��SB�Y�`��l�Db�B}�����ʒz�)86%��A��Dz�_r�v��CF�k�0�|���}���"q�L�ٹE�����PDZ�gj^IܡOT$�Y.�ڏG���b,rٷ��2����{Ûџ<��W0�b�E6kF�^\Pg�K�O�PP��:�Ikk��c�Vb����1졷�u�Ey�D+nŵz���y��!�ǃ�m��x�q��ř`�� �����I����2ӹ�=���9�E�o����Ӎ.���ǿ|�����a�a�@ˁ���]�F�Ƞݍ����u�zV2.��H�U�h{0��rTS�T|���7�m�UMV�Ɨ�*��������~��?Q�Y�m���5�/4�+��K� 	d%Ja ��ܟ�*S�O7QR��zsC\lR�;̛E"���U8e�� CU�s�y�,|�\˂iN�I,����O�\|_�<M٨���:�Z�V��?<0�#O��~��l&�j�3��6!:O���+�e����[��2V[잓��C��4<(�D5�0f���<�}N42oW���=M�IX�;=@�o[wi�Q���pG�nS��H���{�&4����!��N��So6�}#��C�*�y�Ձ�p��ܧp��C�f)�(��C<�Q� ��k�0NyO�:�_�A2l|�D-"����h������c�C�!"��^ޒM��[iR�8AYw�^__g{�k�S{��8�X�vf��gE��:!Is�|�e��@��gG���x��۷7���0����b2��3cM�Q���/
�Vr�B����5x�+s]����%�K����?��U�{��q�r����[E�/���UE���7���3�#����S��*�]^�`���-{�^=�O����H�\���e����h�Sz���w�&��>�_�b�VpҌ�{Dq[�o�7�q�p�.�|^*E��3"�����;@�La�T C*���5_�������U�ܩ&v�v�:���S��z�S ���nS��cÚj�����zF�	�A��L��o&Fuӊ�����<�Y����� D����߂��f�8��<��Š+�
��uKW$){]M2���݈z��������,�W�Q"ݛS�8n�Mmb��(	�֣���ɾ���0V���珣�2 lL{���n�F�E�M:�{+YM��!��@@]�s��=5�ZXɝ��(�-a)u��=M!���:c���%:aiT��T�Z�m�9�5��Cl\e�=W%�D�"rvY���|�Mt.<,�p';�<��J\P*8�9�O����R���Ҡ;Leu��6]M��Ӽ����v}���矻������������ϗ�Њ%W'�Q��07�3g���w�a�R�Be����t��4��٤Uz�z�t��V���Xz.Ī��="��}��&+=ʃ�L}�ǯ�=��	3�&3%n*��l�u�є�zܴ��E�HN8T�;�(swu�삖Bՙ��̺M�mQ̙�|~�|�t�٫'�{��SS0$+����~�/ڇP��ߋkǫ*C���?P����!�Ʈ�
f!,4vm(��C�i����~�Pa���Q́4t��>����ȡ�ΔX�
���M��c��_b�rҹD�Zz�����W��m�3ȃ�#co@�������>#�[���;���?/�d�oY*h�=-��B��"�O'0��h��=3�ިZ�C�5�0 H�\F����uI���|7�G�K8h��
B�����T@�Ƒ�=#�6����5�/�$��h*��u�;�$/_v7��r��������#.KT��b�ٲ���Q^l�5�5�H�:�˂���C�,�)m�G�c����&p���'��q���2|�^EfK�����;u��c]�΂�*eF�0-���v�C{�9����"�LB���~������!c����<Yn��ݾѫ�
>��&I���LKb�o	��zw��!��T�{�-W0/�`�8�F�LF©���T����^F���ɳBYT�`��
�1N4��a~nJ�`W��Wz��c��6�Fn�f4�FW�nl��*���Y�ɫ����M*��X�~�S�3x�.���>��&:�S�`u��yc��:kע���,ͧ��j}:�(�G�
��8ޅ�C�hҖv�G�G�r�;E���������hb���$}S�:��n��+������
�g�Glq���0�N�4��}t�YɈ��.�%T�vaw8��x�|lg�:͏A�ң	lO���ҥk�P���^ڐ-��_v!EeqSʷp=#a݀i��[���y���9����[X�������n����zG#�1>oSy7o�u�Y�ۇ�'wuU5�fC�n!�ӹ@�{�1~q��U����U��e��w8�ߠϟ_5yn���W�ղ�g��韵l�>j�]�C�fO�a�.!s�7��(}B&sZ��Y���g�C�n!��'��%�ZFK$�=�)��mz2H�bhz���z�硅����L-ޏ�0z�<�0x�U3�2�'Z�͟]g�	9o���l}w�l�pm5I�'sN���y���ᮟa�ac��0(n�=6?����@�{�F�5Z��1m��ۦ�OEV^l,E30hd��c��\i��Ppݏyq�db��k�E����0[�q�6�K���;9o�z-�\/���}ȝ�Q����*�����;/=_#ն
Q�*e;`���n�6���wg�sxky�	��� ���~62a���l=Ě�Ff����$i�]!�
G����J��k���|��b�+��L�e���]j��L$:B�ˮ[�*c��^9����o&�P�d�X �����|>	���8ڭ��hnvR%7�2�`��2q.�ӪV�ו�Ng������^m@��Ԣ-�_�.#T�xkG���������7�C�pu	��MT����Ù��z��q����^��b�8�,�T���k=0�ty�C��O{"Dd������u��N��h��N-_HюX���2��|%�T[��M��t;��k��A�]����������u�����o�a>y2��e�a2���+,j�aMCLC����Fp3���ͽԇ�����zl�~�����r���3Y�KV� ������\�v����4x*9��o����`���3��F�����i�L��+��7�~�3�yho��)����j�����9�C�nZ��q�f�����?Q��P_�Ɋ�W��h`38�zZ¦ژ��i7az�zm�:��.Yk�P��v�卹3�1C�]<����t�^��\��{���GwN��j�{��Rd<�*��C�[���Eξ���]��~�"��é�$�B{��Nіk9'ynS1����a��7B��y�$j���F�l�L���M�\`wn�����x<��^�����d��0��>&�;��c&-�A��z��LX�mژҀ��Lg 7E�s!��}�Ubf�,|ԯ����޺e�{m��+��0�.���dy�j%��:u��x��/$�P�ن*Me6�7��Ix�L�Q�Q�.�:掓�����|�����������f�LBq1u���*ѻ�2~.8y0���t�T�X0z{�!��UT؛���of~1�D���1���K^z�-S1�ᡕ�S���`�@�΀ތp7lL8ɳ7u;�YmJ��!&���s��*�+�W���z�pA��l�4ɤP6���"
��w,�C�)�����_���|ŏz��`��L/ނ�<����+M�5񑵷xwH����Ql�%�c�<���T�����ؖxsC/������W'e9�%ꕡ��o�D�Zz�lq��h�	�l?���8ߚ�
*q�N����!���U��Eϛ/S�Gڮ/銺�@ǿx��> wu�'s����/E@lX��{��J�5xm	Sn�&*�ۘ��Y��C�3�\�.��4� �54E�yA�PS�OߠE���;�~*����ܸ�F��O����ӻꑥ�_t���SmX�Ĭفw�f�|!�����^-"!M5n�X����j���=:a��& �ݰUc{k�fX�ŵ�n̹��]�M�f��~1߸�T:_F��SQ�9�|:��'6TU4,�yw��=LJ�H��2�{�<i�҂�p�wICԲP���� (p�D���!=��e�Xٱ�7�U�L���Z�q�R7Y�ڇm�śE0�4�s����U&/=-����g=��z��?���v�j����ay> ^G�FuJe��d^��^,�������� .��71�\��Z0!�lya�}�<�����~�ǐa���L,-Y���c>��l����p(��{$�u��s�1k����ndlכ��M�6k��`��as�~3���ͧ��'�O�~!1g�Ȩ��q�Y�}M��@���!>��������Jy�x0i��6"�TK�p9�cN���s+}�dF.E���`D�n�cg��%��*�?X�uHs�T=)�T��EJ�W�\�g5�>�܉��Wݻ`�1pc! ����,i���׺��<�]"b��З�t�".T�e�/f�W���P�{n��m�G�@���1͋��}''�ӄ�.Ë\�ƹtĆO��  |�~@V����&`�7:q;S\�4�r���G'��}fu�:O��-q��M"@����$��������yᙃg�u����!F'�|e>�#[���jơ�=#LVp�2&��]��.:r�+o�>�}:��2q�a���a�����k9�8D���W�o�!�(HH��<V8"W0�ǫ��=�z�ԥ)Kۥ�+;O��uJ^3B�Lj�\��JX�h�����M�1��TÀ��o��H��P����7������M���/z�S9�K�k�p�Y\3�wE��3e.M����K,�:�V������t�u�D����������� ٽ\rq5�跽q�Q�yw�|��v���y��>T%<���ӧ�^[Y���J�V�d����د��MGG�����cJ�i#��'�9ـ��#]�m���BS}�N���廏�o�T���;JK�!�,�,�ǉg��׊�3?Gc�ߌ���ɟV`����RU�T�[�ˋ�ۇr�n�[��`[Ő�C����1���M�L�����VЪ�e�
���֨���r6��|��՗"Uv�Q&�'u.*��^���Ǟ�L��g���s�`Kl��ˁv�֖bFwa�r���"��M�*�({����?�)������'y�!��|��@s*i��|��S*_�YO��f37���:4ݖC��)�4��^/�oPkaY�}n���_�5\|��߅~|!5�����ik �ѷżі�z�=nb��7#zo��;�*�f����ӹj��[�&�a�	ʾ~�j�6���Cєdt?k��=��c(���Bk��0�e�����/ǼH�.�N�/}s׻��"Z��T)��� &L�Gk�����[�ϓ���|��{;���y�y��0j�<p��u��`QGj��D��/�p̫�X����]t;6�Z�y�fVWH#!�ǜֆ�z���W)�P�{bV�p�V�]uD���U���6
ĵm��	UZ"	����l隣N��F��R/(J�%���'pz8 �ضpޜ/KX�/gM�� � ��Q=3{�sb-,����p-��5Y�f�j-�@�Xe��+�Y�b����q�τ9�{�[]X��1$�u�>@��P
�琢/��`c�]h�w��g��D�����h���r�ٯ���yE��^����Å�X����-�;'�K96�T$�7��Y��Y�LL�KU��;F�{/�<�u�jޗJh��7ͩIl�ޕ��&gV��ʔ�;��U�����e�빒��o���Θ�;ÝH\��7��+���8�d�cy��a��ux0F-�	��e<��Q|:[�ͷ���Zn�#��kg��sp�]'�-�gU�Aa��ݢ�3��8d�ϵɃz�:%d�Iꤲ�SX��틬�|/��/����#�~}�2�]n��;��$a�,�_>�ٱ��m�m�T�M��6՗[w7kp�Ν�����e�GF�;��é�b^-�\atUe�j�{�Wj���,��-A��M�tl�¨2�щ��S�,$�,`*m\H�QC~ĳ{�&������D]���0�8`�D$Qˉ�/f�]�,T��;WoU�����1�Q��e緥�pջP�-���$P��C�n
{,6��u8(��$%n�n���N�p�SɺŽ��'dKPe��ͨ�$S�L�d�������<������tcƻo]*������=Cfp휂��=�(�/v殭�hwdRf��:UP����:Tk��,CX�Ǐv�i��O%���΂�Y�4-��m�e��������BI�e<�!{p��	��¼sMU.�C�+V��J.d[��C�u��o'1ükP���q��hU�o0��A��U�﫬����fr�sl1���b��!ƕ�g7�;Á�'�)�s�W}���UWc@$�7�jw�$K�Xˌ���]8����6���9OiMڜ��j���le,�ϝ���e*}�m��4P���c�*��+i��[��������ˮ=T1*�\�c8�ډ]��̓�Ѭ[����olb�B�.�B�ğ0�Ł��fx�Amen��6�.�u�#`��k�uqAg'�*]�b�#�	�3���˹��WX]�(R���x�	z�݅�]2���LӺ�.u@��� ���[���G�?-���Y��Eu�����;���Y5t쇌����	en�{\�
w��Cz_$O&z�����/�m�Ͷe�e�u[x�S�YFjْ�,֝�������5H�����.��Pb:dW�7	u|٢���Ur��j޹�j�[֒/������~=O^�z��ׯ^�}�z�_���}><x�>�~����Q�'#�W�s�!kmJ�x� �0��ں�w�*��զ�����������ׯ^�z��ׯ_o^�ׯ_�������}��φX�#�D� ����%����[�sט���`�������>ch�DD,�*�c�-�*����
�nW��/#�A��p����穦���֊K�xs�������G�`����z湃s<k�la����m;a��z�܃�yͼl�[^EK^��+G/\�	���My�s�4\�*9�G���oQ�A���\�HV/6f*�ysՎ��
��[`�{�*i(�y�sf��+��O9�yc�ѯ|�
�uG����p�xa�{�,y�A �%+4Y1�@�@&�£&cFg�ۜ�j������y뇢�h�_9�[kc[F��#��DB ����(�J���@I���&L�3$&$���/�?8��Y)�L�մQ�*�SQ�[;%�� c��J7o�3���km<����y�`Ů�`��Y��w+&h�㘾l��\i�ۃ�	Oc��''�(	l��F=q�O���@ё�q��F4��Ya�2�/�%TZ�$�$�E�BU]O�Q��6�BD�$���4i�R�P��?�����g�������_��|�~��>���o����Q�[��"ls���O��Z��;�b'�|��lڗ����B����Ui�a�;'Z׎l�]<�s}1���mxJ�皢R��;�m�Hy�Y���l�arCn4c�w�����r�^����G:Di����%���ھ�7���+T^/�QEax�)�g����G�}o�#����X	}�C����}����fΕ��z)��^36�kׄ	���s�u�#�%���a���}l�9��QL��U����<XxGb�l'���`�p%ط���Dn�*�W%��hOC�[�ڨ<lv0"��=���Ik)u�D]�y}�*����Q�}q?>}�H���x�'��ӊ�7(�u����4!��^��ź��m��1W��h�ԗGާ�t%�8����S��v���P�˥�0*L��0��{B/���.�抪��Ž�G���y��ª#k P�R�)� T+|9�3�p&�&KʤNP�XoCUF�Xׁ4r�&�V�3f�;�]ۡu�|����o���̯�ߐ���MM�r�S~���Վl��hj�ҷ�$�?R��<ԂSX��ra��C�u�@/�_Wc��!?.'���R_k��&va~)g\˴���o�Ŧ��N&���%R
`z��GY��[T�0�S�ΚE�gZ���q���	5��r�UA���e܀@��`��vnu-(��:�V_��,4�3y��B�C��Ϫ��X��8�31����Y���<Q_�\����������OY�\�~�,�"lb�m�j��B�d�z����^�@������8!����T�ߺΫ�Y�z����*\���LS.~��t���~�ޠ7j,S����l�e�����{70��57d��<��33�y�9���Js����ju����5)���E��Z�a_��X
1\�E�t=�w��Z��<�)'�m�>����/��Qy��?��x��M�,,��&3������ƺ����;\���;@�q/B��5� ��dA��u��
�S��N�;��##���g��0�3��+��Z�ݢ����8�Jj.ͪC��ހ���������%��OK�^"�m,��ZOt?XǄo/���`��
�H{�<z�6�����s�E��;��>�>�=l���[j�[����9�ح��Zm����{[�y�f���M[�y�\ˋ&��u���p��
��\
��x���X+V_���.��}�:ǡ@����Y��2t���a3�u�y�-ML�^���D�ȗ�!�}i��^J���#�: &��_
���+N|���՛=���s5#���4���B} (��X&��͝R���5�x�セ$���(yH�ֹ��CB(�nEN.ɷ	�1��}���r=?�1�D���D�ؠ���p�0#�WW�*8�������D�C2a�-i�"���#d��O3*�tx0k4��3�³zoU�~�߼����]����>�;� �g�s�x�����"��y�UKĈxe���f�-"���s�7����i�[ʷ⌄��ho
o74���Bm�?NT�D��/�*K೪2?lh�9`�1���%�57��jq�xb�G�:j��àL�-��V�z���״�
�����y��|]Q�(<���0��ʾ'�ߵwN�����������ўd�3x�3�:�&���̱v1mD8��uώ��b7���<�������ܼ�Z��X8��e� ͙�:!2�*��S0��t缞�l%�0��P+k`6�)�`xvq�J�V�FeV�N	#Û�_��`bD��=��,%R��U[q�$ͱ��Nn��4��`�-oל���6����J���ʹ�5�A`#�ut�xǢ��O�~J9�iFx�J9uX�}hy���~d%@~���R2Y��68����^xcv��׈ȍ&|����xL���z��;�F��=�n/�m�����=.���y�l��k�i~9�*����u~��`뗷=��H�A�d�Q��寐�BƩ^�`n�Fy�ˡ3�(?��[�t�`�����x���4��/�i�bz��ң�{�0;����@�jj�Qs���s�����>C�6-��B��ne��� 9Ϊ�u+\oP�)K��4`�135J��*67�NX����'F���V�+�6��QO6e���}��Ϸ���<x�)���߽��}�����743��o����hF��=R�ϬAֻ�bg�C�u؃�#�q;
��<]�]z]1OX�Ry���>|�/v;�G|p����U�ިZ�C�8�����{n�J��o_x|�F�JC����'F�1S�ycd�����0q�0�����+=���Ueܣ������*�ix�;,� f��;9����f�s(z0܌�x��m�tl#(%���g�IA��K��?P�q���Ӂ&p����48�������ަ�к�6v�[�[�G��Tsy����V�}���;g�U�O���y�M*rv^%��)-�.��T�4���鞼9hzq�������c�oC�0���^�m���o	��0�W}FlW�2�x��۶�����N^`is� ��{��1,�RYT��e��"��<70nQ&	�O&�&TT�{+5�!�`9�[nk̡为��/ l����� ��QJ}�5o��Ǹ3=?\�u�}Kk�==��,�v<���-X�!)�`����Q����M�lBbzx[�-��=�,�����Q�Qg�Vk�=bX�Y|=}^ff�9�,���י��t����x�l�z�~��Ċ���y�Z�K%�e�¥]0��En5l@��\6�k`�'	�i��u8��<��Ū�W�gE������?
x���O�{���7��㜳�[�S�s�T։"�J.͔���$N<�����n8������ϹƵ���ǦY�*G��'Gj~bk]��"Da���WL)�	��:�ekxm�/9�N���H�z���=��|_�B�r���7.�莅'1�^�ŭ���w���"GuH��1�X��m��دq����m/p6S��%.�.���[[Z�����W�c��Buױ@�7��\�s�T%�f����c�'�?at@�^$k�ϯ�2
l(x]����,�	�
6xha�ڟi��5��Z��g{ru�=��&y� ��O��瞉���<���Vm�C���DQ,��种cyآ��a���ZN3�{�[P�9�ˡ�`���͆k��(��on�C�O��hǠ9��f���yݛ�����/�m9N���e��o��ѭ�=�㐁��>`9̈���K�ZE{�=G��g�T��P�x��f��oi��?r��[և����)��ܿ��B{��߈�74�?+��w��,�_?��A*(��Fq�R��C�m��yET�Kqq�K4��#���k�5�����zw[�o��*_�Ɩ��l^wsc5�(SJ��ݹ*��e��FiX�ΗPᚾF`�n�m�I� �oEms���I��W۾�@P�𠮐�����~���32:l�r��m��3�5�.�6��z�6z�nwyڧ��� {��o��� C<g�P_��y��_��=���������޶�.�}6S
�ֆP�9B���Ke� ~��}�;2��o�m���"�Rj��N�(�p[B"���~��OL
y`(nG0�3�>�{�Xusr�ɒ�ѻ��d<�n7���ڮb	&�.S����I��}��`���VG����g!1�t:�"e�ihث����G�_��)�q�5�q[�j^;��x�|�v"�|!�q!9f�S�Xӏ��*�t�L^s��ޮC�F�3���ywZ�X�{ٕ��[;/m��[�H�i��^p.�۹v��ڎ��S{y������3E��z}���Y1L��S�H千r��q�DU*�{��B/-�U�t���]c��wv�E���6�~�~@k@��<��S�q~sR��@�h)��N��'PZ��-r<���j�uܵ���gx.���ĳ���Ϣ�Kϭ7���/�ڢ��Q���9�a�JnL������,���E�DO�0�3���|" ���o��ށhȪ�<\Q͘Nv�m���<���i�����^uŜ�4���SMD�DƆ
�	?��H��������F\Q�cﮙ���z�����:<մ���ޏcD�2=ѠyP3J�ϴF�)z�� Q����SB�.0ˋI����f}�7�z-�wEF��h?ƴH�`���pd�v�#`�3y��*��w7�Esx�}W�fp�<������Q����(���*��8�q%؇�۸k�����E,��!{ʏ���M�p���!�!�3�|(>�s:z�1S喍��g&����C���[9{e腴��a1-TL�l�Q� �(K�W@f��ͯQ�MXo��.hK�5E�7�y5k0j��^5�&³�~�I@�(o��Ow� k�;�Q����>�XGv�b�?i���7g^
'��t}�������b �=��/"���;�3�"Ao4�T�ՄR�jAw�νU���-Y3 3���Dz��/!&zz~�����ݑ�.�D�C�CN�!�z�=��{����s�v��zx8�Sn��S��Sx��O�[@�1�?*5)��?~�5�ջ)�������=y������Z	�^��r�����z�b��0J&��4הxqY���Q�f'5��|C��-�b@m���1,��J���Y�.����P����X��Z��z��� ���f����5K��1R͛����Y�e���^�ú!2e�{�b�m�������@��;����B�ƣ*�cZ,,�w�g���G$JPy�?o���Ԧ���m�-N6�4������������wH;o�p�wc[k�	|�r�r�]����\��o�h���8�q�w܆ �_�c�
[�A����Q��Wl�]��qi�w�d��1����� i�!�%�b2tM!���V�A��F�w�~���;��ٷ� �����
�������{;�\�jy����1���`-�x�4��	��k��^�R����<ҙ��PWs;W�c���蹈�����O0����mr�zS�jgއ��:m�[�����	O�'2�,��]8�y������3���I��sX)����k+uTO�I~;�!���ҋ���Mm��7�{� *wJI�D�7-��BƩ^�a��Cut'�`�些	�>�P�5���gjv�{c/,�G�R�[~~�Jk��gM��Y�֐K\|e_!,��$����S���*�����9_E㟕��@����?w����cp:dGV�_�O���S��Ƒ��	~�{ו�K؛8q�$}�8��5�|�A�T, z�ώ�#]����6��}��X�<����:-E*��<݂Ȟ����pa�޵�"�ٚ��ٔ=:��*��wN��CҬ{���>�
;�
����? (r�i��B��/ߘ���~��NG�O��Bٴ��u�{;��SW��7��b�л��"%K4����N��r�����S�v�)���)��Ð�����P9}[�S��ݲ8Q0�'��7�"��#�n҃���w���a[L;�i.��l��SC��1�[���:Cf��9��w-�3$gi�I٘�u"69�pw���*N&�M�-��P�����DG��x��<Q}���|���_w�ܟBkM���L�;�m*B��!�W��1�鵯~�Z@�
_o��H�k��: b��2}&�4�z���򋈉��/B��&w���V6�Um�ݼ�>��܈{�-K�5�]G�a[�� Ŭ�.�g�,�)���X�!�}i#��7��o^f�$�|[&?~��v �~u�M5y#q�O��X��(��x�nư��m=�X"�wue.
-���q��n4<�LS[y�����%F0�Q���R׫�GYѼ�s��9���|��Z��f�ca윗��y�O����'�>>��F͍�v��A���y匼�r���-?r��Һ�e�Oei"C3t�_[{�ӌ&�,xb�f�J�CDiB�s{�f���]��ҥ8˝�k�D�ړΰ1�.Qa� �v�z6�y�[3zټ�v8-���jJ��e%Ծ���_�Qz��SU�w=n\�L��ȧ2=X�M�61���gb��]�ѩق!��!0�F@	=��)8���E�U��@s������Ϯ���7�H�d��	T���hU��"SÏ+��"#��K��ƣ���I� n�O��-�,�C�'{#|�_+䷲;�m&{��w.`�a���)Rج󋥱��/�uX�1L<�V9��nVq�D�i~&�1+�۵���,ŕ��U�#ǲ�i�ؐ���A[(�ͣ�F�:]��B���+m�n����r22�n8�y��h���n���<����ޏ7�� ����7����<%r��V�7U��i��#�Ƈ�KK�%��H����_�uz����CZr�+Çvi�cq�w���W��o^G=<��5%���k�����႑>�����,���8����f�&�bI4.$
�+������PqO�Pׂ�����r��E�7�W<�׷=�K팛־?�������A�e���5��z&?�Fo���.�����?���&��<ڡ�;�<�ܱ=Z�nP`���}��Q���z��ަ���r����u�5������D8���+���ļַ7�B<n�"��~k}Sw�b��R�|��#���XX>`㮞܍ޞf�ϐ<O����E�030�}�����L"�g�6��M�`�M��薪PSϳ t��ii�v��)�C�W�b/��sf:�m9��\�4_��1m�
Ƕ]L}8ޞ��v8�?�1����ں�5��V�a��|��2S�� �yx�^�z�e
��VS������M�|x�3�0�\�u���L�wU+	v��e:���2�WBק���z)��Ĥ{�R9ccL�Tl8j|��Y��ȧML7.�2�[�+d�;�����(���#;c���to�)��;�<����t�1�8�V�αۊ2v����7�	fުl��m�Awfځ�8�CT#��D5w��r:uu��u��n�=R���{v�ؽ�
0�9��)�����㉼n�R����E�E:�o@hPk+s9q,��G��MWbT�"9���yj��R�� �����7rn<�e�;��"�z�]p�\�~�������>�2�f�Vno^`�P�X�"�ƛ����ᘇ�)��\I{Z�<��|_`�t�Ѝ�o�2�O
�q���$��"\��k*�����f����@�Ʈ$��z1��6%��U���Cr�؛��\fMqT9�ֻz��e���֡�k-�Rb���[a������وJ�sЖT�V� �DU����:��U���*���.�\�4D��&��_Ƙ�+�M�'N�gI���an��\��]D��	�S�\E.݅p��q7������L����7�N�ᒏ?��z)�"R��z��X��:�Cgn؛[��9�:����1L(���d[�mu�:��i\)Ƿ���u^Y�5����mUy�%C�S�Q�����wV��3W6�mrް�b�A�{5W��|+3	��˼cr7�r,E��������a8cOzJVeΫ��%l��r��𹺌��-��[O{�`;C�b�[q��z�\ʂ0Uw�[W�#[DTF�˱���;kW3
���˖2kVlV+"�t_7o�����o��qd��������WJ�E�K[%֮��w���fV����,��uIywW;����B�X��8e&eR �n�[W�]h�ɘ��������۬�Qw3}�L̉}\r�Y��湪뗣G$Z:)����m�u�id����x;��v�.���sXyF����pA@�K��XR�l!�]*7��-�{3p���8Y�㢳�C	�X�ý�ҝ���%��6��1�}����o=۩�'�Ҙ\�嬾dSq��{*h�_Ԭ�?㫌�<!�Ϸ̞bИ\��r�ӱ��mE	Yq��f^��Chf�C`�F�+�<��\b��4\VX��Їfu��
1�e�샵�����ܹ�j�b���E��*2�GWL�y�,�9��_�h�����)��Nn���8��O*�L� ���#�U�f�g.����akt:�ܱ�j��%0� 
�4���
��۫�H�	tt����f���5�c�w���X�uXi���@ġY���d��]��+yث��fe��v_%y2�G�C�ē�9�q�r�n�m�E�!� �IkM��Jj%QfVE��]�֘����r�<�8Ecj"�6�V�{��S�-�F�Q�n\������������^�z���ׯ^���z�_�������>E|ޭ�=����[m뜼�9�h"���k��׏��m��8p��}g<~�O����>=z���ǯ^�z�z�랽|O������C���Kc�֣6�⭍�����*#��O6�{���⢢��b�F�Z6��p��i�m~cy����rw��j�-��˕�ڍ�ѣ��ęLa��E�E\bH�	g��1�iŋ���mF��,h�DM�U��sy8��Z�KF[lE��济+cEDDu�y�6��Ej�k��yrţm�4M��sk�f"('z�X�*�8V�lDkc�Em�6{�8%8��0m���ͭb�>���s������Xv�5^�r*j֏->N�q��MskX�kw.��X) �8���f6������(j���.�ڇ�6���"�w
1T�Mv,�֔I�R#b�����L]��˘�\F�2�y�u�c���w����<L��*R=��.�m�#�������4��L�,�ޑ�oԘ_����c0�7˧������B/} �9���z�(�C9y�N�D�&��R9�������]"��iO0��O7W�Jg�����Wv\�2���;?��$�Z���\��o>��'b��ދFEV�����`���r��-Ϊ���Q�N0�,9kT���ͽ��h�3�hu^�����Am�u�Se.zӦ�u�Xu1 ]�\�����w:x���:�z�����A�������%����.ќ�ծ��/][d��L�}
 Ɨ�%�s���g�5�Ơ1�P�#���H�I���U�㞯��ޫ��;�21��~���ۜa6����� HQ������L��g�~6<��=슿�`�Ȭ(ף���U�ք��J���7����
Gb���d\�ظ��$`�8���e���H���c�<ݗ��F�D�{�ы�c^��T�g#v��v-�;aI%f�e���٧3��󅁭y\���n����xXهl4�@}D�?VG�D8����>�_�kԻ����VA�A���eNOpcΥu��|���7è4*1Y��ASl��B�͗v��I�3���wlt�W,5_os�?/��E�}d��V��;�Gҕ�����f*}����b���P]ׂ˯1�R�{u���oGN�;�N�� �//?��Y��<UT���{��{���?��{������z�����X��q�<�+$ٳk�@,�8������{3J�.꼞tls.��m��bYm���EfX�ŵ/DϘ����?��G��5׵)��䫵�32�,�I�4
�`}���0�ú!2��y(�%�SJW6�����rE�'/mv�i����R.�li��@�:�Q��^i�
�U)��*۲ﲕ�6��,�ιC#ɧ��T�l��ڧ���'L���6ӄ���T�q@?��,��T��j�t�N6ȫ4ޖێ�nAB���K�0g�������'֡=�"�ҎoF'6��+Y-�ٵ����� ����:�e�`n>�����������>"6��o��{�ʘ���OF�B����-K���n(^J9�2�X�ꑃ\3nl��y:Դʄ�`]�ކ@T�4�B_�N�"0�5^�Sm��5�W�W���k`��"G;��,����"��*նv�^�v�G� ~��xa�믠̐�	n}mװ"��y���X�4�h�f2��}�H�ʱ4�Kęz���C鵄�{ɚ.f\�A��p ip�K�*����V3͉��	�2�-t+5&Q����������͢YU�}˞!���1��L�2_ͭ
.�:.u�M���������ϟO�U�_�����<P`�{�{jwt�ո�*�RM�o���x�22�6�T�
��,��TL�ս2�Ԥ��Ɠ <Ʉ����~"�[�1^���^��S�F�qm�����0��rn~�l��<(�Ο��n�f�;�F���N���E��~������e4s�O�j�����۸��s��v�+w�2�+ �{���{���e�C��>�o�KL�&�,��4Ʉ�`7+�zR��B���bL�d�g�^�A<�xRί�2��Y�b����|��?36�����c�P�gx�����Q� !����k�5����=��QtT�1zF'���_�v��c}"�)?%��n�5Z�G���{ ��L.�ǁ�{�]+^��� �����M��r����[B��!�-�o:��qV7i�F��� }���a�J�	H�V��o!7�}F'���&�|�S��� -�8��xTwy��RւS��֧�(n�����A�ii��[pk��}����ZNV�jv�������d���wRbo
�`�͝�8�W z;���
oG�2| {#��J��5Ul�ehA���9g�6ix3!�N�>��b��'n�C[����]	l�#a�e�~���γ�8�VH�E���`��N�Mi���uę���;��8l��NF�j�fFm1�u�q/���8�oR����B��wCn����
��@��Z�����8�XHhFM�ﺷ������]���|���{��}�
/���"�ǋ�=�=����n�'�TX�<6�#ս}�>�Z�5�����5�#�2k�C�h�0�f�ܵ�y�D�9�Nz7��X�^ӈkcK�e�d�2X����EɯNe�c�G�{�3���9�Z�b�vk�yp�a��h��BO���|��xdUj�k�gm�i�?x�H���V��M<L��7�ȕw~���h��p$���~�3 |o��0yAh���s1���q��c�ػ'q���a���}�����O�>6<�:XHt�	�A�k��ߒig罫�t����݈s ��}�GL��cˈ�7�,yЏP�$s����5F��u��	oyy���&&&#�wʙ��Sj}������L rZ�b-����yw���s1�'eWЭm�gYӍm�AЛ�`��ǜ���/��َnv,Ȁ1�AWA���:[�0gh�4�w+�yy��U�>T�H���m�5S��2��,a� ɽ\`Kf@*��ap��s�}`B��h���Q�_«�"���zo����{a	E4�}^gM�nJ9y��{]��Ъ��W��M�AS��@�r��$(k�/՛�E����&��+�q1�qe�ٛ��ٲ����w۽�Md'0ٵr��jۮS��t�+q��dH/3:$���j�(���p�n;汏�| ���<'�� 
AG|���������*�1P@�+���;���r�����~vk`.�?'���U<�Q>����׵5/W4"��-1̹�R~�b�@��qw�=�,*�� C#m��E�Þw�66E�C�GB�7�Ɵk:U3Ź���wL���ҧ�+�6��׭fR�X���Y��!�V�}��^��������<��B^��3�!��c���A��~NA7�\��{��9~.��[ԌsF�?��n|���a�PI?���_��@�!�:�������2�H�-��5)���@��d.=}&k]겫��M����`�c�j�@M��m�Az]��|��	6������|�����)�\e���yVʜa &3�?`znz��k�!�z�Q�7�O�t�F�! ��	ñ;bv������ �\W�L=y(�q�T�ZcX�;k��A��3@�.wK� �d�}3X���Se*� ��u��kyH���u�x�
�g�O�A��-E�6�q��`=�V�[�+�]en���`��F�i�\tCcrq��7Cޜ^�L����Dj� Eyf�1W&��_����}5�ub�����R �m1�`í�R�Z�R�^���vF�Ӕq�7x^ 87C��5�����u�iV$oe=��{(��u��\��SU%�I�)x��U9m��y�~|�w��"?���<E'�� �Z�kW`����R'�p�Իs�	��P��@dB~�(7��0��~��f��Z����]wv8C�
gg���JDL���ϲ{�Fp\D�˴��>4��L�e��<�w�D�H�Ho ;��e�ꉩ�k�¾k��1_J{ƌ�_n�	z�oo�=�XU�̏9��������ZAA޺dO�4s�3�
Lg���rz�ږ�=O���+*�T܊�G�DsG(	�5>nF�i1\�c ����&��[>W��7˞6�x�Y��/|��
c{Z�)��0���Y�f��wB�W��_F>y�S��}0�s�bW�(�`���ZD?k�p[=kd�XOt�`�2˝�8�lImkʸޖyK^,�p^�Z�T�Y���}oG�Ih!�kh���GdJPy�?D��&�M�ٺS=c8�i��IuLח5�S����>5x������Tz����ne�p���_����C'����!	av9�xd1~��*W9kz��[�_uD����`���9��z|ɩB��z"hT������x}Vfm�m'�q��5LU�W(���pM��L)�.��Hn�fjV�}%G�r��+H8�f�&r��
ҧ+�;7p���a��p�pu��K�x�2Ô��p����a��̫n�&�Fg�ꛮW��#0g^��������>�� �2��}��<x爂R�R���۱��W�]�����~�n����fwnmiT�3}:���D'X��Ʒq�6�\���O��8^Egw��hu˭ʡ���sO�����Uz^9���*��{�Y�V��k�S-�S	�g���
8%ܶ0P!cT����6�6�A�7W]f�j�B ��_��-��1�J9�~7���s�i$δ��\�,7\�3�^�5�&-)�E�����������b���`��-�g�2�Tm�핆E#�9�_��JRS�>�߽ƾЎ&'/0�|&< '���ǂ֑����������]35�$�Q*m�y�b3��.]��Y9�wԙ8���-��!�ߝb-�s/%ݬ�d)�r���3^�9 b�8���p��K�9S~\ZXu&r|���e�qHw�Zcj!{�*:v�mm��¶�C���w�CØ3a*��jeVe�cH[Hy�u	���k��}��%r�mMl�Z�/�#�y5��B�}F��X���T��S�ކO��I�=x�Kej�v9E�F�/�𰪴�Sל���en���?7:�� KVz`ryP!Ղ�R��f�Z��K&�K*�r2��nf(�������e	�\�ɋ#}�J���a���'�#=�S1����#,C6�k�ʭ���'�HA$HBN>�
�T^�f���%WvgG}��;T�!0V=7SoE��ɷ�4�m���zw������>�����*�;� �������Z��!r�a�� o��c�>w���YB�QN&�������R��a�(Z�P��Yė>v��{�>*E6�oM������k��u1q�)���6�(���wڬ��b��7��p�6s	��b�{V�kW,^�����ό5t�{�C'���ͮYn�Ң����,�R�ԎԵp��s�u)��U�7��a��1�-���֠!�Yx/�mb�p���v�Ⱦ�v�j��+_��y.��������g|�A�a��,z�j���9�~�����.g���H�y�R)����>�L���^s>�Z�vU���J��5�5�q��  @�?S��X��q���ݟS�܇FG�p��OC�A�aX�W�9���g�^�744|��h���J���S�}��iN�`?D�xZ�g�[o�qzzE���M�����\��Z<�͐���b�b���e^�0���f����>�@���Z�����a�fKO�����]�z6��B0-H��'�1�0?�-*����y���Z�!��I!��OMe&��x�U�Ȋ�ѻ�n@��~׊���0H��]�,!��=x��ܜ�P��f�`�R�����ml��b[�����9�*�E�xH<6�Q���8͝�
/�������<
A���&]�����x�T�{g����|�k�%ņ�U�j1О���U-���K�ʊ�gІ�[" �O0�d��g=�LT38W\V�s1z�#�r��8;�*n�g-چ�;���i���w�XP#�섞�Ϛ� ̀�t�l���&R�o�3�4�L�ض^"�o�tF�mK���pKEC��{u���C"�"�����^���̞c�t�O/՘Sw����1!�_�����Khœ�T;hkk��?���)���c�i.�����ۼ��p�G96~��C�z���F%�:ũ|qT-eC	���W��摷�E�E����.�v��ܻ����+gZ���Ot�M��W�Y�Z�J��r������i�q�FdV��o�W)]6�(t˫'���ᚻTƽ>�3���L�=iJ�w��h�*x-��i!
���o}�X��v�����H��F��f�ǧa�nפ�ɐ�4�a���-���)��o���q��U���WmR���{\Tt?8�جva�Λb�6k�AsiH���B(������B��(2y�F~F�6��öUF��%r�_�2���S�"�;Ԝ�!����vPM�qxp��S?q��O���+��vt��9HC5	]������P���O��)�0v�//,R��5���_ҫI/\��>���/Ǯx�O9�?(�ZU�uϫ|���c�>.(.�nj�Id��WѽB6~~����|�_�t�H;7H�B�=�w'P�������}��RX-j�l��i�Är��)p.w6�����mx徍&������8ޑ���g�"�@z�Mn/L[z6�8ƍecg)����M�v�u���|�	��r֮%��=�[�p{���Nh��QP{�0M�U I�q9�gMp��C4ӯ)���<���b}��1}a� ���!F���㼬w1��pN��D ]B՗�ۓ�mT��1r���ώ����ߠr~��+�=���a8�}v�um�R�t�����U{�چXY5S!kA�3l+�袯��חxl���D:JME��aC�s�tH�����<�(�!��1�%m}N%����캘4�H��=9#C�;ܳ:]��/�[�����Ԁ1Mr�F!	�x�M�ި%����0�#j�:j�0�ӛa�J��oef�ne!;�X�r%�5�ϤoP�^��)�1}�i�{��zJ��Dd���@0qP�{ Dp�^�u��4_ok%Jk/r��%ݾ���s�J;���΢Y�w�n��ra����óx�^^�� �i�r������l	)ݷ�������Yt�Ti��D�^ ���K�!g>9�oK���uɻx՚ˏ�N)�{�]�g�ÿ�o�b'$@f}�����I�����[ �nV;�l*m���%�.Թ���aɆ�(g:Nc}���ۦ�¢olD�HJ�T�����i���4�.�]m٩[������6�_1hg_��٫-��I���v�//{;*w%r�����xɖ$c\�:t�<b|��P5�\��x{�1�Y�6��%	[�$��H�C��X>��s6+�ɧ�d�-���՝O�B���K"�m��t�um����9�T�*u�YrJY}BY{ѵ��|^7�ם%�sx�S���Oq��^6V5o�H#`�vm_SQ���S)V} �[�@�D��b�M����
�͗���4�-��9FS�G4\z Tn.�\n��efC0�̤�̓M�D�@�2�*�#J�X��Ǎ�Hڐ<x�SΔ�=���E2���gs2�Z+5�hF N!�\+h^`z����亂hb�nwpOj퍲������ڃ+�]�`��4���6V�weg�C�a���o[�}�=�� q"�8X;�ރ{]W�H����h2�{��2���2�I��v�R��$һ��N�*�h���"�mpt������C}���LZS�j�.���]^<r�kFY�'R�42��/-1B�9�d�c&��ڛ4j��M'��}'L{��>�`��:P��n�m:�HU�:X����X�����P\{�����(��N���(�0搴ݺ�ʺ���}�簓�
��s����ڽ�S^�o2����m���IOMd�/U��t��2P�ֽ���QYq�3����p4���8�cW��7R�w�25*��Ω��k�)i9�/��_
�-g�\-̏���B����(����ޘ�E)W�#6�t��>��/A˭�m�T��]6�v���PocP<�cv��Dә��cr��S���v��S��|gNY|
"kƍ�K���,wvS����{8��;�fe�7�G���1�Qpa;�78�<*�&��A�&�HJۓE���i��i��U9�nU�pf��6��e�V���O:M˝��s[�B��c:u+�pP,giDwP�;���s\��Q+%��.�=j��Q��?���,M�,DN��>�Ep��㩺����/��FfFn�ؼ��|�����Y1��XX��0�{+'	-$�n�S�s�Q�u!M
�w��}��٠�\�s6d����>�������<�Z�M�p����kD��ǮnI�s�����~?^�z��ׯ�^�z����ׯ�>?����x��O�ml�ǽ�F�h���1^sqi�9M�U�~K��5Z�TE�j9�9��������x��ׯ^���z���ׯ^=||O��������o�Q"���ւ�[i�mml�"-%%8��5'I��nUZb(t�գ�xr�M��{˛˜�Ͼ5��mZ���F-��W���E)�ճ�0s����mi5�6���ʮZ���f�b�)�I�4�ŷ8p6ܭ4��s�͆C&Y6OЈ�ƔL�AD@@�I��I�eXJ�X=6ڍ��x�lV-�ִ��U�����F������O<���h5V�ƨ�kLN�˘�s5�lb��f�#��5iכ�4F�^s��ܱ���Nm�	4��~��$�m�	$�,��/�\����(9�%ϖ�<�2��ɪ�[��^O�Ý����#ˑI�CI�[���
f��pS_?�i�M�A��cNS�	�:���ͼ�
Nl���(.�IK��jJ�=[���܎i�s͊�������&#��-��?9�O�����4o6m"	��D��e6A�41�Q��`�
���-@�M3�W�H�ߗ%Wb7�v���+��#�JNӋ�i�m�=yE]p
�e^Sm��q<u�p0�$"駶�㗋lqF�榧�@��BA#�P�\d9
h� a�J�A@IaF�P�I%"�� �

#i�p�ʐ��.2�Q"T��b�&Ti	�<��s�79�������g����<<�������������}����8�l�U�`e��A]-�i�/7#e�ޙ��uY�~@��(��J�y�8M4�A�3�;�S#�/w�{^S�\St�f|�w�V�ݲ��!��vc<�����f�R-�&Ʀ��)�B�z�]0H�����-���\zy�j��*������ �m�v瘿4��S�~�dmO�鯵��^4�QN*-)������ݯ(��=9�O�d�7RR���8v��[M1�O�^���tKf3�.w��UOn��ޅD�o*������_&��A(����Dd�t�P�C�T5���ރ�+����g�C��*A���㣲��[��{%HX���6�N�s@�ŭz���q3n�xwX���r�V؝5��hTr�����Z�̓��`ٶ�Y��k�`�faM!����}���Z��@x�	9�;�s����F���5���ߛ��s��]�P��T�G���Sm^JA�V�V~U���z�k�сM"p'�!�$G��}����R:OD(e0����D!�Y���^f��1H؇l,��l�h����y�@��u��2`�Ұ�P�s�3e�b�:�*������e�q𮒢P�̀��$�q���e����;.�$@ zB�֯�����)�Ιg�C�˻�}�b�'Mڐ�o)������Dl]`�2Mķ�A��)��E�J�[�|��x��(U}z��������ߙ��
��W�kdek���(_)���ӓ�]��;�`k׆$��U��,1BY4�p��O3��&-��y6�ôZ2$[$2/,-����8�Bz�;6��w�)=�#8�kK�칐 D�O�H�Un(�T!���"��0=��^;�RfNZ=y�GǮN�ϳ�Kk[�몭�P�D=�>�W-"��`iy{��o^���oUϥd�`)�{I~���8ξ7��fr�ɻW�n�D*��?X��^��n�b9������Qm�@%ޛ.snE��JS��ܶ���SG�q�kj��H���6�ȣU����*ʭ�x���װ�&'�5����9d��T���@³���P���0�(�y������!�9��D�}Fb�T?uW�A�O����l䍠nE����r�h���X��k�`�pu�b�xb�(��M�=J�8�<��/��Q�vA��	N��V�h"]�9aM/����ޗ-ƷhW={	j/����t�5���밖�`_��Ms��+4n�v��}@Ia�"'r�X��v&�MP��21�Uj�i�9���c [q�H*�'��
[M�s��v��Q�/�V��[�8��AS��yLךD&�N"�m��ǤO^9"3���(�6�}A���ݰ�K��+�4��S_�^ι�����~����� �<s�!i>|��������]B>q��
h���6�f����P���X���7��]q��n`��{����b̼�6:�srx�/#<��ǯ{�����9�)�`�Q����7A�9��Y��pE��}�O���?L�w<����thz��Ҿ�ޘ]*�ȃ�����}.�ؠ7]:�7ɮ'5?d�`��P1�fӒ3�� Ls�9�->c"$l!2z�TJ�myO�cR}C=AZ��,��j'O�?�;�B�`������<�׍q�����UIm��3�	߱.��ɪ�kʭI~� ����OL"8������R��)�!C�����w
�ݗ"{&�^+��~1��s=�}{@���z�������@E[�1��dW鶟1co^���e��(�����ڕa�PC���K;��_�#k��X>��n�2ñx2a�Ht�qF����Q�0��2�5sȭ�����+o�z�67����Qa��8s
���ə6���jg��r=�e�]�G'�u�>c=u,+[5�"�/b��9Ck�Nc�|YU0��>�Vg�m�4#��cE��t]��N�;:|P�����-��y0o�T��{+R��鿓�r�,�}Z����� ��ݎ��뛴l�V��c��7K�OI��Ԗ��7�t�Q��
��� ��	�8�$��Cp��;�w�\�����۞ �9���S D�D
y��{��_?{�|����uN'_��zq�V̰��2���ě�+�L���Y���Y�W}ޕhW��^�n���
��=ˢ�^�5�'ÈA]��������%��Weǔ�Ӭ]Z6�.@�0*�=�=����sP5m40i�֟Pz^@lR�Bi�2t�h��y}/��lM�&k��Iy�y}�h~��~JW=��\���E��Ї=/��P�1�E��u@��x߲��i���,	�՚,-#%���y��-�f6@��%�%�E��(����W~ztcs�y7��:����j�.�Bt�w>������74��N�K�4@WI�����j��n���V:�q��J���#��R���޼9�nx��Ȳ�41�����]�o*�4����Yf�7���OMQ�,���C���΋5z)o�R��Ke�s>���W��Sl��e������c�7h��8���=y�@D,=����
7�����e����[�:�N!L���#->׆|t��>i�N�'asױ�]���==��rrtn��ݳ��/7 �Ȣ^6�%]T/�|�8�9k��̳AÂD��o[;��{4GKM]�f�s ʃnp��1q�W&��qmZq��q����]��a�%��nU�E�v.ۈ�y�<�߾��w��������O��<x�� "U(����o������>~{9�TTVb�Sl�&Ӫ�ɋǦ�'Z�а�ٍ��u�b  ���=��*]���4�hO]0����^k�>qR�T��q����}��^�;�u������=�]�����~�� ɾ��S���1j�OZ��r=9<&�S�a_-Y�Q�ވ=Υ�5H��S���ۏ)���	��X�|��$N)������mգk��7C�����qiu�L� iKT�@]"��СM3z�3�ؽ�l]ʱ��7��oDG�!y�n�v.��Z�lք*����~dx�ê������T�s�S� ݿ��};�.��\\���{s�G]R֤�����e�9�f�6��z@M�m����e�2䫴��f��m�i���ޮ3όJ��l���1l���ѭ��CV�0_���#���u�8g]����dL�:{�5��v��R��y���1Y��={�x�\倎p�y��4x��X����,`�Sy���z�C��������y��=n�G2���@��Ƽ�'�z�:��2���A?o�`ʶ��Wk�LT�&�]�ة�����)l�W��u�[N�A�ce��C%����\a�H�wJJSM����ĳw�)"-_N�}Y�J�0Q��Q���c{k�^fu�%VKg�A��L;��Q�����"�J�Z�mE�:i�ێ�⼥����]�]���+3Gt=/0X���;�pz�م�G'p�������~w�|��</������O9�R0Ȱ@��Ͻ��y�O�s�?���ڑ1��Iy�<󦆆�|薫JF[�g/ϲ��e>]�{pv��6��m���O����s ��|آ��it���*x��@�b���M��7
�X�E�>�sj_�0'����"׍W�����|�3�3�3���¼!��}��m$�k�s[(���9ۘ����`ccI�:��=#h�.R�Y��z�'��+��)]~N��4+`�F� �phA�!vlR+2�*�|�P��	��@�6�Շ�يz���yj�זu.ẖjh��x1v������ʍ��-qQ��y>Mp��D�g��i�����=�:��Y�D@�~~8OU[i��C;ɉ�/��Fo*���Pώ�3�z��>�bY{N�����9M��J����M�r�&�/�+ɠ\��S\�`iy����j�!�(#����D�W�G��|���x��nK$N�S�39��j��}pD�!U�����Iׇ�� �yQ�f���E�b��\�5�/��m�T�=�S�7�캵���a�0{��zz0k�Vҁ`��#b�
��SqCq�٥�J����%����1�xestHv5��^H)=�ӓ\(]X���%b{u�Z̠�u�lU�|�m�߱Ql��W���+.�Y�UyZ�X���%�/s��eeu&�3�ﯜ��/�׎x�x��3�����o0����WH
C��ac���@ɵu��* LM�T/j�cj�c�Ǧ|�l7Q�D���j�����U�3@���§Y��#�'��%C�@�r��9"ڵ�I]s/�+&��C,�O��W�\Hnl�ɤWt�H�Si.���ya��y���#�-=��q0gt������u��y�K��@b�
/���]�]�)�����P��»Ԓ��j�g�y{�_٫��4�Ϙ�
/< �,�O/�V)x�{�~k��XЎQ��̍�W�~E�/J�h�ٳ��N3�կ��qjXH�������.5v�0�ϙ���o!u:�D�N2���t��5Z�s�m%���n�y"�&s�)����p|Sf�z�Yt���#�܃�ށ1�6��,�U1�������t14*�
�/wB!o��5�l"��2��[&�/P�{�6�l�^x�!����+}��]��ij8�ީ��=X	`���>���(�|½֟{T;@��q#s1r�_���?eֱ���1^q�8l٧b��w[�R�K���� m<ȹi͆���<9�w̵�XWH�T �U91�ʜkH.v"�0�Y+D���Z�q���[w��lҴ�5�J�VB�*����#�UL�7W}���^n}����}���	��<��<sƊH$)^z�߿�?y��}s����~���Ֆy�_����V�Wʕ����E��N6�;Mmks����Sc��z���-��_Dy�H�X����w=:�����=����}/��Ğ�i�=�W����]l�V��pႶ
T[chn��
P��7B����N0��Z�<�C������RP�֮�.gl<,l^1���>�u�56�:�Ru�le�9�/FF�Ǝ�����	nt�q�ީ���������z�-N�j�'�P�I��"qS5���ev�f8s��{�؜&����K��1�q��.�d�Ҙ��j��
��/����=����ݶKJ��4C3�Z�.��r�q�'��{j)�k���ן�/��='MW�C���º��{�_�<�9�����/���8�Q��J]���VD;��/��^�	���ǒ�x�"c[��n⼜�A���^���qU�$�dS���-��s�C�b�燪7�ȋx�(rw����}}��m�Tx�ZW>k��8��v<��u�_��"_�Aa��=�۰ua���U�����Ƞ+3jTɅ�c]�����R�]�[�\���>����\M��f�q����r�Εd��4u��$�s�E���<���s�$��*��X��d-�v�}ز3%_#���ot��AiA;q�hT�r���w�f[l]��zb~ߏ��T���IHEE	G�?} ����	�{eX��%$^8$�vV*Y6��(��m�mfe�Sa$u�ߥ���ǆ�׬a%��j*����3ᭃ�[��ɸe{vn/f�,�	�,/ށC�����p�8�<=�}Kٓ�t�>�r�?Y�
E�\��יm����`����Hvt�9��<B�_ȗd���[vz��O��5�����{�Z�4��U�^�'Pfo�s��T�ߐ��G�<��4�Z�.*z'س����Ւ�����lczf�-���>������9�}/��3��x: ��T��D<��E@6$�P�
"ͥf�Y�m��lc ���Ϛ���}_�M��X�U��e2 �����p�9��������Www���KW���Z�%ƵH��3�S
����c��Ț�6���v+��~X"���U�Bݳִ�n������=�^m��%�<�r�s�hP����zbYm�*���H���^���:�y{�$EϠ�n�d̴<�v������Jj[ � �wL�Z��kڈrz��t�^�,�a46�RXh*3�Ǳ��,i�^�	�������$���sPG�ݫ{�{�(�0�+kE����]��׮eJ�6=�nK~�hG�B7�S͏��נW����Eߞ��|�s���I��UI�:[��f\�
���C�n�+׸v�˙X�B�t��#�����g0�]���<�\�j���s���I8��]��~������QSǎx��$�A���}���*���:����z�;I�uM �4���J�z5���ʨ�_�Sg��@�|��;�d�!��}m���|�N�װ�su+_���מB0/��m�]���em�x�-⬩ uhs����D��u%�|L�%N�cގf��27]э�E�ݻJ�+�c��r��K�a1[z�@��P!�]��k�j����-��ж"!Q���n�M]�f�<Ƃ�]�@�yTS��@E���	���:Х�jy�PgvKB�7���ͯ#?�8�c���b�ſW�����/ͅ���lk��T3���O9h��Õs���үdFP5^��릗-~!�^�O�}
%��	�>$��|{5ͩ�m��{����A�a8�Z�C�/y}�f�I~U��D[G=I���p&���˨9r�u�����f�w�ϬAϢ��͊}�^�Ô6��h�	�7�+Χ��>�,'nG،��t����u~��*�3'�՟{2}9Ah�`w������a�%[Hw��b�޶|U���u�s]^=a�g^8��[l&��uuM`x��;i��c����.�w�5��^�]l|�Ug$�.3y�C���e�,m�&��(�2���%�M��u>뼼���q�QɇL'������Kv��x�Ҫ�k+RZvY��uO���]�&3wo�	���*�;9�*�3H�]�g�=�++U��M�%t�0vPA�Y�V�΋v�M�]f�ӕR�ʦĸf��y������'R,�V�%���"�=��԰O��*>xq^������Y���6��v�}�4R�	��f�((fP��C��_KE�5xn�W	;]�����>�@����+]n��gO���nqZ�FYc
Y%�V�s��sI�>�Uk�Wm�4�)
��7Jc�/4d�z&2Iжj�b��`�)�f ��R�7T�5���C6����銆-|�3������ ���\��ٱh��yN!��869���#�!^��ϪC�w�������F%�s�\�,zGL��a���f�s%��[އ�6���M�so�t<9@$�[Xܗ�oym�pvik��^�w4�_p��Ȕmh�3�碌x� �馎���Gy�3'p���fgb�8(1�f���,�s6�X�['IV;�é�&M`�7����RS�9L�Q3�d�����Δ�#����·y�b� xR4WC�uc92��������>�v[�Y��i(�	ge�]>%9xӡ~�Z�� <:���?1f���%�R�R��eMR��-�.t*�x���JqF�m��r	Ŷ�[Ӂm�]u�fF�aj��K����"7�f��YM�t����z#�@�,���v��kp��KPIky����yu�A�[�h�ǯ*�B�hc.�kmd����h�k*�э[�.[Nq㗷�m:�Ob�y�C�
!��#�i�ŝ�'.�&����붴r�n�l��un9�T�*��);�kE��Q;�)�Ril;n֢�7�$�)�}��vw�㮛�{Q�{���<rNnLR�bf�����(�-g,���5i���)�[ܺP���;�-7Y���]ʢ��2S�_�
sp�[��v!���z�P��w��k2sLJ�჻�E01���j�&Һ��|F;�*��}g4L�klmk�Ɨ���V��D��Lrܶ�Yf㕷2ƈl+I�U�#�9rv���t��X/VY�����$��y���f^�S�U��%��FET�q�cld�}�tѼ6�:d���7;Em�&��yԇ(7�s.j�\Ĩ<Ɛ��T�f���=f���Æ���{B8��+D�#oSӋYh#v0E<T��{�9�I����֩�ff��s�M�G�P�����$H�D ��*����)��p�6��W6�S�cZ�A�F���1���uZ����>>�O_o_��ǯ^�z����ׯ�^�z��������9�|"bbh�N��gmh4�v=�5�=����\5E\�`�3�NJ+��x����~��㞽z����ׯ^�=z����������9��(���1���P�sp�ζ1@R�%�,m��LG˗)��T�:�����1E�h�`�.mU�c��'��<�,Gj|�
A����l�G�����'��
���j��h��7�s�O��QMQTZH���b��1��SQ:4U�ft褪h�[$��E4y�Aכ\#mW#�Eȭ���[f��h�v�LҾ���%:�E\C ����&DI���c�<�&��.Z<c�h����UTS��X��EP��kKʃ��
���~��9�P��h�7KG���-\���+cO�q%�P[D��Z�/RxF�sf��O#��kllb��N��
H�����$N�N�F-�ʴr�+��������ɥ�^T�z�>VI߇����{K��({��۔�z��c����U��T������!�,a}￟|�~������'��ej������+�����?9������������ޟ&'(�F|���*���� 荟�Q_;��޳3�G�2��8�?'m5I�cV5q�v�\DH�{OBhT��EȦ�`G�ū��տG(v�3I�]����Cs?��*�-�̶�YB�aU�3__�������'���?T�����۬�'���=���)t7��^�R)��9�zk;U���h���ٺ�8�ݧ/��q��[)8���
X�>a�������J���d&�x�^ժ���?8{S5
n�	��X�^s���K�d�B�f�/�3D�U��C�FH	�t%C���(ZԤ�xʞڲ:h$�����xD���>�L�0Wp�7|�WL.sa�yj�b�y��9j��8�2���TԸ��y�]����D#��c�NS���j��1r�x�'_S�j�g���Zwb�3���,�2O�`^�?�]Չka~xD��U;�E�|��#��ߩ��7�9ѫg;wf��RXe�` ����Ɏc�����dFK3FߚCG�2rТm�&n|�k.C���dՊ�{�(�5P9�I�[5TؔRW�LVF��#��S�Z gT¼��؉$�];�bfYKvv��
x�f`D�ǩk�Sw/	8^|.i��;r̌{00���xf�d��c�Uc(v+&��Uʝ��;�g3�J1v|������������3���)i����`�B�;�)bq[�zɜ3y�oT8>mw)ŐOU��[OH��k�>�_�&%�2��0}ٕOw��zy��'ܐᕺ�q�21P֟>��]�m�~a� �>1Bc� ��0ӵq�\���5�5�~�z���A���>�>���|��W�W#Oͥ���v��l�g3�}�Ul�ŀ����3��u��0�������U4]-��c[O�{S��H6�j����6g�y�D��Kk��}>=�Ƨ(� >{?D̤!�@�Rnb���wEwBfE�{uz��?
T�]�W��O�g��?J��ߢ{����c��?Y�ؼ�f�*�k�W���^Y[�e"�jD�U�)�����%\H�y�x�vTJ^�z�c���^�X
���n�����Ly�
�`�n��mm���V���.�������q�St^�Jɉ<'��h����>�	�4U0U�[j:gͽ0��>D�X� cް�f
��J�a�bo2�哑U�HQ��'za����� �,_�%���%U?���y+y�!���3m����}Bʧ�#��懕s�	�P��[����U�͞<B&d�Ħ�h�\��-�$��6$�r��
�ݝ���&�.i�j��alࢹWo��_;�F,��C���E�Gi�W���|>^��D����?|��������$۫{ct�&�b�U�WF�Wdݜ���v��4�~0��
�P�lu����܄���_�jg������|�g������C썳�Wp�P�U<ܟ sR��˧���Z�(憘؟VE�q��xMu逛y���ze%m�k�a1�ۚ7Mm���El����ڮa`$d���ӈ���:k��|�E�<���==��ww��3Gd�""-:�Q��B��W�����a),$�l�k�>�c3�s= �d�,�ϝs����zi�;6�kߦ`�Լ��<ޑ��OL[��S�M`-ŊU�95�:Z�S�n�x�)-��8mk�ޫb�!F�hu�s���jXaw�����i�=�h�Sɣ�i�`�k�TlN���)#cԻ#��D.u��'_��ԟ�4���Vu���sj��关/q�-F.Z|^�������*s\TϲJ}Zװ��Y~.���j̠*$���Џ}�g4o>�1bx�JSlyM4'�a�ٝ��i�fL����q=R1ϩ�Mϩ:�[���\�oʇ�?KC��81y���o3|�|�}댍������N���$�nQ7"r�*��ST{����ZoT	H"��;�����1Wk}�=B�V�gs�0n��)�̦]<�0��"~8y��Y�(��\{�_P:� ކ�b٢� �l�6�^f�xp�Xr�̽��FڋZ@jr�Y�=*����?�9�9��b�+�����_���������[H��֡.L�Qwvg�d���>3 ���Se(�c����^4
�FwG]o��ߦ~2k�x�"�6Ϡ�����%����R���C�1,��M��+K�7>��rB�$P1���ٱxIX��5CU�j�6�� Y5�WO�~1����|5��!z5��j]}�{(��3,yױ��'IQ}0*�|�l;�jFVL���1�4D�ۺ�ef�0�9�9yb��b\�nx/�	�-��[��f���sg�ӭ��4H>�i\��HV������m%��'���q��������o9s�Y'�Ҡ��sL8v@�B�s�s���	7�$����uvO�~w��R��ͼ0�s{/��ϕrs�U���ޣ.@*~�L�u�'~j�)wP�T���ߙX0�;��S-�-H��R���q)��I��a�`��"L�ث7��k��ŪB��El�/�"}�B�s<�K�kDgM6'Mss�
^J//ж��aΞ�\өO��N0ɮDȃ�`lakz�g�ߘ㞟=�����������;��[$�ۡ��X��n���I��A9�]��睝��i�E�=�M��qi�:�b��+��n��#Y���^��i[�<9:�E�Y�Y+m
�x��1F��f57�b�f�Y۽B��2Z��Ni�Jq�D�K������ ��<�)=���������7s�UD�C���?Е_�9�U ����:��<	��$lyx�Ŝ��,��ߢ�����������������B1*�d���zF���I�����ک���4�ڝ��"p�skb�+fڥ�&1���+�3�P�����K�D����P&����x�Q�O@9r<EM߫�uqo��~��4gc	��5"uA���c|�t�kdݥu�.zbC=����q����.(��T�;I�w�r����9�<"�priuIF���,t�mJ�ju�q��K�����E�C�@}�T.�Ƀ�Pп�*(��i@���A��L`��
Hb�^7����I�ݴX+@�T3�ƙ����|���0�}�-.�`����`����2��6��s��7!`Ht������m)zs�FC���e�=�*�d�NT��W�w�s��3�,YE)��'�O�����+^�P���*�j}X�[�FK��p�䮱����|1{�?0��&��gN�����_Hf��N�y�#zO�iP�a�2�l�\�r酮��rANH2����=�Lf`є]���,���Kfq@M�5�l����v�p��Y��q&�G���&B??+�^���E�v����<e������bZ62l-nK��n5�liJk2h�#�*YH���o�~z���{��><p�8C�G�|��~Th�������OPh�$���!�z��4�t�H�R$wT��Aoi�p(b����f��)v�fo�^��L�ۖĉ�,T8�x���^�l�<.xd��:2���q�M'ܝ��a.Ù�.�~5Ő�d�X�}cE6V�;�����<�1��A�\�^�e�å�����ӽ|�N�]"��9Qa�����lz��c����8;k�����! Gz)еy�'ǖ��=��#�N/;�A��]�,��/�P��>VYj.��1�~��ټ���"V�����[V��^@��#��n���V��:L����1e����^*�%]i���K�5��^7C�
!^\������ �?/g��x�>�yP�C3�zu�uG!�78k�n��_g:I�X'<��Y���)���{�=p�[�E�n�Es���l���=��U�^zVC�?�Th���P����4c#(�]�o��W��m�jCW���*�kt�P�/���a%w�,�b����>��G�l��;yj�_�[-���vF���k���[vr�|e����A��kH_s+pM���P��cc��[���c�[+Su�&�{L�KI�(�q��Z]��]��W�����Kܮ��w������~������B�O�;�W��������M�ج�"up�l�h;�q2VX��mm�s�r��^�c-��j�}Ό�5L{~��郑����c%�&ꅼ����&ptK��gT�ٶ�e͈~��'�v$�s��{k�)�OE����46�S���r����
Jem����i�l;֌a^j�p��������_t�O�T�"MXT�덵etn�ڍ��6���n�o��ZC��q�j�:e�Q�'�ꉚ>�A�, ~1=��OS�'Uһ\���}^J}��G,mɜɊ�a̈��{(K���!p�N���Ҽ��٪A�CT�;�Kq|sR��.TX�_��ig��6_"D�"���o��y��](�u���t1�с�c����Kj���IRd���{��i����=-�(n����J��tsj��1�
���O�*=�dЪ����l�t����JKg�����9r�?n�-��~�;�b8R��վ���X\�~N��|��S8ޑ�*d�E�x�
���5ܔ�n����&s*J����v�^3��~0)�:���Zs�%�<|���������W:f�pF8s�<�dl#XıoU�i��eE]^�Yg�Z�k%�.���u��k.��i�������e�i�Y}���7�{N{�H���Ʈ��x,n,֛�aE�}�yC!�ܩ�w�чH�����<���|��o}��{/��x�p�99)E{ޣw�Q+z������F���bhK�wz�K�;Sǝd����.�����"�td�T��ql�=ع���ư�`q0X��g�ʙk&W������?�@�E�^9���Dp�Cz�
-��v�C;lO���8��v�o��b�'�����޼�C!��t�@�d��3�ɭ��5��M�0@C�lg�����wڭ�;F(�ǹ��3n��q��B͚�LN^i}��-;r^x��g榟E�O9��)�AS�D&�d&T	��#�yCS���b_���@����6�~T�l�c�6��	j��G�S'Q-��X�
�wϪ/e6�a7��`��\Ȏ�;��ӎc��<N���ʡh�^CtX���s���PF.���v!��L��E���k�Qj�!�����d^�d�jY8�F�̘/!��;�5��km�r�f��-��[���^�J����"��e�ה�R��<�[uz��m9�^/kg�{b�F�vc\�il�³p����,��͚��1��pZcBw�O��ޮХ})H�F2l��c�y��� �{�S��°�������
���zn`���%�sښ��?P{��=%+�Jx���g�$o����6_M宮q����}x�����
�����̭�<K�
�o^O.-�~�����"�"=x@o7� ի:�U��T!�4@B����LB|h.��/=ƄZ�oW#"$�K�24�\]I�aw��{^G1qt:6��L����q�ֿ��K�0wt���<���ǧH���\�gB�Y��y�/�����W�A�7n0���+�h B�/B^u�/_��ۙ�ı��gO���j����s��dl�Ԍq�����j�PF��$�"y�66Ȉ�����g�|���[}���'���V��S��}^�!ן�{3Ǘ�]5V'\߯y�g�� �gg�Ds
r�8�wg�/t�oV��
FAOX��p��m�m�^؎/@�6�͗Ϊؚ��UBOnB�%��>���xz�(>��u#�*�R�P:G<;��4�����5#5�p[ �,H�Վ��2z�ήF�W�������Gz�Y=2mkqlv�}�p��ȑ�e5=�m�%�줕0�31U������]p,L�H����(�]�8��N���o��ȬA�n2�iW��ɵ�<̞�1-��YOq>�֮�qdϋ�W�����]GqS�+����8R"�	���5���x�c{��m��b�C�n�8T��w8��6�j.R�#1�D��{U��ww|�D4��֠/k��*����֌�*�3��J�Zr�3��N���yy�W�Y�@�p��N�1�����7&��or`|ﳛ��?����IǎNQ)4f`<���Ժ���v*P��+z���W�Ĳm��ݰ�dL�Sp�������,nBɖ`�둇����̪^|�n5�׶FV�,z�{�z���l�
U�������;P���K'��'a{���e�&�<��2"����H���+	��+�P~�Gˢ9BbP"�iUלcR�Y;҈��ͥ��*�@f�����w����[K���	c?~�h-c��,S�N�yu��g�757��;r������}q�܅o�?���U��eN�cv&��ޘ�Kf�Z6:���ݲ��c�(�#ϭ�Q�!ƻ�>0���d����ץ��獊tW!���ot����Ն	t2�1jH��hLc��k$�v� ��
&|�W��igz�T��UT_b����f^��
ܴY>�9��읁�d�s��&�\�ֺ__Ӂ�_�Dc1ˢ��T�7r�=�0l�ֆ�!�E�0T;�S���1�t�5Z��-��u(a�7�q�˭�&�C�4�G�K�2� ?[�fH���C��/�O��Ӓ�?@��<��lI�9�!qp��=�zD�-`�F�ccl�++~"2�3�cnf��S����ʅ��r���N�K](���Y�Ú]Bn_<Y�a�
쭤��d�����kju��s���c��mF�&�JJcdw�n�fs�w�.�-���n��jX��|s�V�|�\3;���;rQ�ObpK(���o9
�P �Ԏ�����[��f�]����Y#�3u�� Ÿ�S�(%�Q�ܰ�6.K���M�vp��$su6�bƮ96NΦK�5��Wr��J�cPw>�г��S��J����1G^[�s5U��!D>]>\9e��n�|ź�/nqZ��T��	��t��,����8%Y�Sn�ˍq&QV���%!��u��q�#�2�øJr�W�٤���er����37u'��֙f�����t޷�����Q���x^�]�J"$M�إ���f��z�i�!�ʅ[8E�Tɚ k%rrSŷ(Im);^�Z��>r�5��Lk�]�l�M�ťz(�YS���_f����&P�S��Y�*TE��{Yxi��S#�ߢ�k�]�g]-Rv�+w/k6
�뭙��-��PaI� ��Ō�^�F�m*BT���ڪY6�ݭ���P*7�g���]�(c�����u�yA3�q'���Ͷ�8�p��o^�=[֟	X��1.ξ�.�����TTM��m���ٵ�� �oV����Ӽז���&�B�¡�v"���"��aNsk�!�/\P�:
-���;2�K�7�5rn��)]�Dq��7���g�ܽ����}��*�ņ��uŎu��Ź	�-�,�V��s�����t�j*�	ݙHӠ���"��rQ��Ls���{J���;#��1d��{ʉ�<(�C'm�I1����eH/!7:.�q��mE�.�E�Wf����0퇵oz�c!�j&Ze�6�c3��v@�N�]�ys�wf`[��������l37@Hұ!={�v�5�v �hvЍ�VR��)��g9�+bC�
>ݦ�j磨=-�[W4�i���0���ŜD�&�����4Da��GF�Z'���(�V���n�����:�v�I�E����Z]7�&4��Z�n����h멟LS�L�@]��qvO\r�eIi2�&SL�e�4�
y��S��ja���k��8����iX����L�a÷z�!X���z%�\���8��^�X��U]A���=� G_tv9���6b�nLP)���1��P�>��U�c�a�|!��@�.����Ep�pH�Cu�Wjwl��"��LI�a��ٱ�:����|�n�N$�o`�A�ܛyL�	��D��-G6�oR+ů��J"�D$�	��b������(�h��1T����k5͎Z�"(�B�l{x�������z��^�z����ׯ^=z���������������8S�"? �TQ�sTj��Usm�h1���y^B�$��MF���f���>=z����ׯ^�z�z��ǯ^�z������?����o��r7�npkF�Ś��9�V�5��)��NI�+��9P��KQ4DAh��b(B����V�(
+�8��ZJt��[ih��NsEZѭPSH�a4�ѡ�#�1��Zv�6j�@mmi5mO�ˌ�8��ZJ��#���WU���ڪ��T��\ܷ�w��G��ȫ��ĔP�N������mIEZM$IA�]N��)h�cEhti�h(���9hlh�����b�Rh�(���G6��3T�[��ѱ�������'�h��JtU1���N�*H�ZJ�����5Z������9aъ����~ZO#��/!��'�~JE��3_&"��#�GI9���$$�jҌ�!qF�i��S�d�1���5	>}�S��c�Ԇ�Vk[���t��R{Y�Ƶח�5��#��s�SCVbz�vu;����.��2�D�/�Y�C�Ƌ	�S`�f�h��nHԐ�ZA'9`����-8�'�F(�b�a#P��D�	d6��"d�
�(و���)E��PG-�	l�c3��G���ʃ��&Z��������]���뿿R��6S�|G:;�|+'o]WL�!�j�|��D��S\�/�qt����O���g͍�s��� �a�(ufصݽ^��ܠpi��E��/򯼢]Ԙ��z'�G����He��[B�`���k���%��i�8�,G���@�.�jm�*�ᆞ�؆��;��h&���o'��U!���B�x�;�4������d@�[uT8UR����޶���FLI� �0p/vx���Y�!��Ma�"�V�覤L7{�w����]�C��*�J;xeu���wx�m��_U���:p��@ny���u ^1�w�]�eK��Xh��:�����k �*�{I�C����>�خ1���_����򿇋����{��҉�9>Ҟ6���a�y�FV�a���������G,��vևRRX\� 5�較�Oge���1��j��ƃ��n�q���;�����h�����N9�36`��k� �|�����gt��Mj�M2Vqs�b�җ#lǅ0ûvBC�<�4���+�fHP���}���*�����7��	y�����n)��ȫ�\��_�f6L��� '5[	�;t�Nkq�lɢ�8�k��o�<g�'�(��~��~}�I��<#�=�pQ1GK�{�j��J��r��;[4bf�:鲎�s�dBjY"级���Nr5&�}
�;k-"�u)~Ҵ�����Ԑ��(���<=����𿛌�'s/[ҵ�V�@�V��zo ���~j���t&G�z�{���Ḵy����raՆ�a�B�x^�odDjӴ�<�T�F�A��ɵHqÂ�h���\�b���dn��7;2D�����8k���A��9Y-!�k���wQ�e�z�|�1�h�{��h�g����6-`�g��u���O��8۫�R�%��k�AiO����_�)�
�{��.1p>N9���vL�yQTY�N���(��X�u{���R�~nc���]	=��Q;�(j-���TJ�μ�k(��~��_j�F��}� U9�~�,Խ����reY�B�Ӊ��CS\V�_y	ݳv�� �@2�*�Ә.\�ܝԹ���IU���oCMwrGM�[͡Cl��<;9-G��>�c���WB6��rm�H��Tu�BQky�ƥh��C �zc��v�ga�A�v�>���[�>y���}���~9�3ǎy#Cf��)U�ҕ�nS[���p�;�Uo���iKv�q�=S���p�W/��$�J�.�D7���ݜ��8�|w���AY^JR��ݪ+2$^4*�`0�� b���Z��:�����v��B�<�<Jѯ�hJ�u����6}����N�<�QOOy��z�O�9k��J��j��lf�_��)_l0������J�'ޛ-`(����)�z}J:}|��%?�S-���{6�Q�U^M��n��{~��:����}��������͊�پ�-7����۝[��b��J�|����e�fe/̺<�jQ lֶ�s-��5���K�J��r�{_x��/��O�'�g�(3	�}=�����hnW�Y<r� L^_}W=_�8�������'�~���BFFIɻ[b���Ӕ;��ҍ̘{kb8��{7/�9����Akq���lf[�5fHnn-A���X��v`�]��r�iYx��`k?e��]pλ�7�Н����\m��3���]lr����\q�&��u�CLf;.՞���s0>��n�	򽗆NSonsBx�Mx�7yz�O��D�_w�ꉙ���$���������Ͽ���������9����Y-�o<��pY���Tsc�S�W<s��Փ�z��I�j'x�
���o���>�s��G}m����ښfD<O�Q6;˫�%�������E��w�T<\_]�`��f�O&� �uA��픬]Gdx�ƽj�p�n�:Ż�T�z���*'�:��βOU��纶O�o.ρRaZ&���x�(�V�C]�@�9��ڨ����Qc#Ve;�N�b��1.���%S�3��i���B�V������`�"d
7�+�Tf�~�p�YӫzCt%��]�e�6z$U���z����n�r�1�-pB��^�Q���-����s}�!v�_�Z�mգ�{�ϕ}m��l�󙉙���WF����NKWV۷���Ә;Iޮx��6ܒ6�d���^<�7!>t��u���t��|!M��]����w�1�u�����v��z?m�y�hv��#����Ӯ8��P��i���%��WDDj�⮎�K�Rղ�x�X�@[2���O�]����M����.@�u�ڽ��Զ6�4����.�8�������;�r{~z�>t/������,��4��y�>�N7cbg�X���i�R��aTYX�6ۊ��xa� ��������J��w�rXӖ;�O�d>�+5+Q	�����MWEV��havy{S(z�R܎��l�/���[y��?�A�Ɖ�q����8�n�G�ܨ|9�V7K��w��vs@��B�V-;��_�3���&�\�+j�����ݷ�e�=����N�n����� ^C���4@��d�Ȁ�} @*(WE#hT�rxe4��rR�9�ݔ%�=�WGu�k�LV�
�G+�w=�XdD�(OL["��-N�[�3���o#�� �5S��ڙ����|��;�5N �&c-n��fw3��ŏ��'��=j@Ϸ������:}SVvJ4�[U�Mr�J�:��*^�&@�زnCg�N{���*]['�GT�3�����w�j,����8�ՂTz���#-�0ʏwr��:8�T���62
;u���o��=��k�븕m>q��{�~��2��n]圵0�\"�D���ﴀ	�&��cY�����
�ל�
��SW�� �tiX�5h�f�R���}]t��ޠ9d�|�����<s����j�vuoK��S�}wW�死y��j����R��;0x�ӎ�9�{��n�Je�t��(�x�iU_+��c"�9`#wyM�쎧�꾾5�sL��.�Q�^�z�JݰJ�r=�b��T�jG,�;�.Q h�x�ӧZ�פ�oofK�ew����2�ָ������W�=�3�o�����֙sI�'�)#~�0)q��[��R��%]����'���r�;vMw��u޾W`;��شfE��O��-�[�^���:{�-ɋ���Ntx�0���41������T}����v�NM
�6����U�\�n�9Ҭ����fů͈ȁ��rT\؁����&*��wf�����Vh_eK�d7N������nʨqA4t�=���h�f{c��7¾9�B�m��o_�0<V��E�/��[NͻN�*��)�=�:0m�T�h�/{�P��� ���Z��3:RE�&���Sd)��Hv�ǛZ8��$�S��l���֞cð���m_e�Գ����!�H��\ͅN�^9���\��x�jU�����^�8����Ў�%��f8�vp���+��~��z�o�k���r��i��׊q�72���n���]��%=f����[��5��v����>���%��x��p0L�`��D|FHVnGFc�n�c������+*�"��5U��l�^�^*���4}�=O��v�1QOsr�Tf�ى��_�M�UQ#����S�)<:��z����řU�M�g���/O�t�S���F�[~��ʧ�]B��%��u��ݪ�X�x�05�`M�`�>Z��&�0�i���m���I��h��+א�_xģ͔���s��C6��;ͻ�F ���~Q$v��9E��5.w�B���X-��eR�e![�w1���wvf�� �����ޅ��\�u��D�����~��++.��x6c���hn�\�L�5��!�Ex�PN���t��Ϙ����8��w?Q����"�Y�ȩ���K��j�a
H��s:��J7*��ZT"_*!��3�m雨�E��u��~�ȽM��6Fo^�],��Bi[�[����*ȥ�t]i�O*y�ET�.���M5���k�f���wQ�0,�;7���o,�7_����y��|��7�^f�Ԗ�Dvg.��r&|����^&��[.��F��Bā�h���G�%��B���<��C�w���U��n�'>g>М��Y�q/�G�i:H�&�+q�3���%w�w=�C]j�����y��2~��.�ޭ�UW�:3���1)�fF<�fp��\W)Q]�u�d���әmٚ#��\��ng�sFDUx`�vj�Q�zf}V=�Mm��q�cu\�Kg�Y�/k�r�<W+=��EKEm��k��)>q���Wǅ�
�l�8Ӯ�<d5{�7Yj��{�ܝ�;q5��Y>�Њ>
BQs��r�{-e���e3�d�U�+��w5�to*����8�0�R�%\`�}���tk@f�����f��bcM�[l7D��ͽ{����Y�ҭ��)��-Ŗۭ5����37At�ɕ�У����C�_2�"J4�օ?j��6�
��]C�"t]>���.�KJ��.+������43j��Υ����P��S蚳��\��ʞZ	�2�t=ؒ�E�Ua��D�1&ܠL��iN�b?}��>�}??�����������bo���ą�/�y
܏w�Ӣ�F�'8�P�^� l�l���4铷��O8�;���۳���*���
o�^.�t�
]ѢR�b[������!�����_sy 68�W.Bپ��JY���+"�`�w�ot��V˳]��G�-x[W@Gv)�����^�uSoM�7N��<&Ļ	f���j�ͻ�-���>����b-ۛ�Hs��nZ�2�va�̝4bI��b�;^��*N�� ����X��Ĩ_N��#�{�b+5��ފ:�!~� Nk:�y��^��&�8{�t*4��Zf���_Vp5sf���v�lĮ���ts�872�[�3�F�u̾kK��e!��9�K�]"�q�2�fz�0V��e$����'U�,Ihա�e�O�|��S���H��vX�[X���{����ļj�K�ƅ��x�'u���\<"�yVx���8��]ҷ�c��r0�dx�U��j��s�m]���=]�H�fk]�;�]j=��t2޼3V���~ڱG&�4< c��ƅA\��u-"tֹm�'<V*���2�N�˧b��9�k�n��;f�����ml��ޤ��#����Cz=@oy�fZ�a3G)S=]/}�ꚸ�b�/�Q�O�)ԍM�^6v8�T��w8�ᦝ!��bi]Ѣԋ�5!���{f[�>��%���ۥ�N�H���|�tOR,N���^}*�fw�՝w�%�VC�:��9z˼��C��z][]�%��4��:���B�f��ཽg;�#���b]�z�1����}6O7y��՞�՞�|�e[v��a�k��1Q���DT���N�����^��lҾ���&����9fy��͞�����I���͗��2���L
�pzS@�ݐ�	Q��.��M#�Pm�Cʌ\R��縺���V�Ũ�z��AR8�ZMzqOu6�k�wdr8�B�l3��yzB��=���~!�Ĺ�G{pT�ݝ-�+U��⛷Z�k���QSi�����v3�W��}�r���ţ3����G�ݘ�0����Ddg[^� �)�nZe+�:rЧ��C-�H_n� �ˑ�h��3}�lB�����.f�����`��hJ���j /avjf�`�n��a �cTIa1�J�{����"���t�L��%Im�G��� c,{JO�C��W�(��Ʊl٦�׺sY[��a�+����b.�������Kx��e������ՏF���V-"P=��s%p�t���OE5Qn>��A�R��N������v[o���ڏʥ�������ļ=��ܺc��c���
�#��ߺ��r׻��xM��kܰ�0t�wym)tB���hooP�9�MS����{*�ξgS�!9���&�Ӟ��.�2}TlVG"s;a�ղ�޳N;�1��U�]��v�N�n��"��1���Q�w;�k���Y��d�˷RT�FX!޷���Swk��D�<�6�0[��h������n��|U7�ݰ��X�s�`�yc������ös��9T�-'y"3;o���M�cE�����v�MΓ��Wc��2�4�d���=���iV�lg7M9f-RRg.4��eR��IN�z'���2��p�lӣ݅7)�y�˲˙+`�8GhΥ�Dm̙��ĲRubX���%�է�����s�\����6��uGw1B��rS�kYՄ J�6�P
;X����ֲ�T덮�lO]�
n�Fr�ws~�M�;%F����O�K�tJ����G��np�B�B�o?n"v����k��[m�NW����}������j��i�7h���lq[��\��Y�Vt���[�[V�I<m�:��a��;�Nm��`y�� �˼�|{�U�**�KVl:�z����k�zhX[�*�r���^	յ��Cu�[]���Κi[<��Y�������πn�n�Ժ6ҫ0�i�(�U�g��c6P�y���},Q�������t�����2��s�qs/��U(��'��.:w7�]�9K��jR͞
M���9b�)\��k�Xr�NuZO�hzv
sI���9�z��.܌+��7^�*���>Ѹ6��^�	��kAr�z��E��%;L=��Z|1�y��3IU��Wt:�R�iC1Ȝ�m�/bXS$�nE����[�=��@`5�l�m�mKY�/u��u�c`�v���,_5�]���J�w���ŗM�`���*5��;��9be&�T�U�ʒ`R�Ɣ���jgV����kɂW�aR����|V���t��`:V�׭�����AS� :Ir���K4kݱ������-+0����v�V�rh��#.r)�{FӐ����5r,Ä�J]��2���ә!��|
1�.���ݰq�]����ށ��͎37mv�h&Z��m�Nk-�n��;B��o��p����������{|�-*iZj���E��z��F�))[���<|}?_����g�^�z����׮z��ׯ�����_��/�5�D�:��5T��#e�D������@k�9����~?����ׯ^�z���랽z���������~ϘPr&(*���N�֝|�UTU�G)��@[@�M%!W,����h&*�(�O�*()�4r@�Ƣ-�K1�m������%��r�Z<�AIE!T;mj�i�"+�ϐ�O*5�5y�k�EE�4z�c�5A��4RR��:8� ((ր��9!B�<��T�Zm��k����i=I�$�������A\�BQȣO 14��>o|4>��&��Ӡ=ZJ(����:vŰ��u�8��JS����@O6G�|����9ri��)0�z�9<��N�@� i~$
!i��/�Wq>��I�i�[`���R��c{��JmŴ�E"{���k��輛P������r��}��8�������.監B�٠����Śv�͇�ᷙ���F���h��c9��'#�Y��"#��>�Ȱ,wd�f�����K�h���ݸg���YV�ى�ܨ�Nl��MݷY������`�v.�hP	�`����	X{��M����E�^W�z=�}�<��Xd��P�����q{쩻����F���ϾP�e�B�O1|�K0g�44aܝrdi#ܩ4�7f'�mۛXzoDC�a�#�r�T�ILM��eS=h�`�����uU����,�r�O������cP�LwT�Vd$�U�4�*0`��gN�����z��aTf�j�P�"h���nU>sR���H�}��S��NV	��YX5Q���o V�z�ٲ���32^o^j�볩�s�﷜�.�@Mnm[�=	 h%+h3��ڣ2i�����&ė�m��2�7TA5�7Z,4��\�o&p�+E){`.l�j������^����p�F]�"����^�G���f�Qバ���jܻz
�aM9��V"2�D��q�0��MI�p�Q�����6�N�b�N˒�����W�_�|>�LL|k��.�몹�ٽ'%#���T�_���W���Fu�7�[��e�Hk�4�Mj�Þ'R�w��0�i�L�0��[^n������a?R/���y�N`J="����N?d���]�g��j�k\=����,����c`Q5��e�y�A��WM�X�|��<{RX5��ф<+%�î��4f���p�8�uPņ�eOgLE%2aќ�[V齴^	;ŧ�Y���Cu�cFg��Yǣ L� ������;1}>S)=���9�mY����w9�/k��<�G̡\�1�T�'6n���a��x��n:Odu�S�X��օ����1�=n���Ax�+7�8Wz�4i�0c�u�l4B#q���q͘�Y�A�y�Ձ��d��hg��L6�&�a���Ah��`9���f��QQ��κnvn�q�=e�h%���z糥ʏ=����\;��g;�m����ye�E�GG�Y��7��U��˓���hN�tyI���M ގ#�Ƕ+�HaZE.螌N��#��mr�3��B�z���<s��ϵ���p��s�y�ΛӘ'�������d�k	C2\��ļ
MR��o�vE_h4O�쒭�8ө1@x�~�u9l*ltSN�U��7yFԭ��,3/)�1r1[)�+w���#�O�(�lx���
�xL�򌊸��*]SV�0�R��,�ݍƷ�l�3���q]�Gfh^�^�d�ɮạ�%r�Y[ >�o^z)U�N�R�Ѣ��f[���#&d|���>�lз�j�z�?�_O�û�N�֌�g����5�P&��Ga�������s�[h���7=K���Q
��Ӻ��y�,Wwy`g��a-�Տԣ�u��B[b�|y<Q�����Zm�ui��5_BW��y�۷drC��l����Ee�b�ޯ��K�3t	�7���u�:���Z{]��K�݇�fy��q���c�"�������}
4��=�v���MOG��ljp&��f�7�[Ǯ�4љYynm3��-�Wt�(�Ӈ"OuN,����g��zWŜ�B&ZûB�� ��5w���US�Lz��]��.#[/�Ɩވkf���+1��⥰̘���el���;9W��5	�㹸t)F�Y��To�}�����y��?��Ngnr+vĳ������$�j;yI��68²{M�p�b%H�W8����7�_C�_%����+��-��.��#�o���t��ٔn�w^�L��ӧrά�%'H�Bև᷅}E}����l{�<���\��R~�'����v�:	��eP����e��34<^��e��y���M٬� MT��¼kxd��
�,��3�}�������;-=8'���wWG�V&@�� iS���e�[_�����\-�ӷ�(�܁��7^��E��PW���J���5��-���Up�+g��N&��������d��x"*/$>r�)@u������^���O_7ݳ������x���-�e7��	k���?�#��麛��ro�Wd�t����'_��)clһ�Q��'1�-����\�x�[h��Yܲܽ����2)5���SDr�v,)�ԕ�r!�f;ǫN�`=���eVtm f�'RRE[Ô�I�!LP]�����v�yAmc��*K34&���-�N�Ȕ%��7Vx�kX�UD~�����|>@�w�E��+�+??48����ߴk��zV�WH�s@��$tUR�����j����5fϟ9�1�j�j�ww���1��廳��i�r�D�f���1y��^8���sW>g0�]���
���@���a"Jm��)4�6]�g����UD��mI�f�-����tvu����]�S5�^�Q�:�Ά��b|_qY��[=����;o4�E�5H�E�B���19�gfA���D%�[�D�񜰄97>�qY�ݭc�]Uo��-4��^3���9sD�	�5&���Oq�=��X�q*�I��{.kƽ��q)���Ԝỷ����W�Ƥ����F-�{��N�qEdvZ���y	��RH�(����~��*{�1��/��j�������1�O9��뉽��L�[����rQ��t/�
�qW���G�㔪ч�ѱ��I"��F�_m��j0������jh8��t���(h���T5�sn�P�źu։t���䜜�WwOB}w�Squ��np/���ɡ]�zsz ���0��oN��2�Y�_��<}�_����������(e�|~����<L0
a꼍xOt�Q�E����[����r2�w9αoh���^Ս�;ǶZ��׮D�l�yz�2Vܽ��v}�V�y&��ߺ��\ԃ��XM,*�N,w�P[s)2��*�/{�Մ�n=j[�Bw�k_�ǀ�J�)J�NI7h����Һ��\Tr�7ӭ�D�����f*C��/C�Y�;{sͳ�ZT��*؛˱�9{�^���xF�R��՗C#W���s!�qua�,�Z�����PӼ�F�A��.�j*x��qs�$3���K��W��	-5\�ս�e�6(1+yl�N�!Em�<��q�m<b���'�,�}��9��O�\PN���#��œ��ra��Wfգ���sZ��¶��ۛ���'��X�$nk�:f[�:�x5C��Bg��%9�n�l��Ū=���-�jfߦ��+���ˁk��Rk|������V���/����i��c�t�G&E�b��a�[V���#5�7X�E�TTZ��)�!$�݂�悥MՈ9Tje�!�<,��g\<���.��k��Ir���}�^>>>�xF޾�T���۪��Yuy{��-ͣ��	"b���QU�>��	k]dw��ah�c��Ź'&�^���{�篼�����{ �
/��K^c�&Y^��cT����,�W��r ,6���[�Q��K�_m�b�٭�t:Α�}bv˺��p��9�c�T0a�v�=�5���H���l�6���o�0:ޱ������
G�x����r��Kx�kV�;����7x���_+f^�K���|��~��ɾ3�g�8������[��ه�J�@[�|z$�>�mܣ���@�T�C^�3<,#v�x�3��]C\*S�q>�j��@Y����QY>3���;=���������x4U��ɦ(�ޞssۧmA��]��Y�2�4ԼK��t�uWv=[t�˕⽻�0<����K�>�����ݶ��Ou���kj98̚���֧�#��_}�[a}�1��:uզ1��
�!L�֊���&�1�=H��b+oe`���7�8����;���M�ʳ��!ѿ�����8�ԅ��S'��fix�0��'cb�!Δ���)n�UWn-*�o���޼�2�E'�yٲ�8�z<������,�[�ʬ��`�l�Oy���G���s��Wd��yf)��XSBچ����xg}����=�}�.j�ݕ��8R8��>*�_�ǟ&�[��DB׾�ko�ii<�Ȏ�"�h����t�+��y�`�}�Y;��
)���ٽl�ȶg���Ѽ�(���Ľ�N�=��Z�e����[#/ۼ��ɩs�-JG{>�h7#";Q��}03
�.�bT�h��ڍ��qh||�w��<~����ï��~}���v�G<n��5�q���+��y�"�[��`���p������Č�y�Xd�/2���eV���V�e�\s����������\<��R���UXTZ�h�{joC���=�����������&��S8�W>��Ȏ"ĕB�u6�P�D;�P^�.�J�@��&w�*�癉���V��9�Ci�#�3]��Yg
3�P8��ɧo0ȰP��킊e�m�.�ϴW�;F�x ����P�����J�����
�Mnm"�2+2^5yW*��L��@��VڀI�O5����j�Ќ�s��l���f��U�����8�����{2���]!�7��*�3ĳ7ީ����C����>V�kD�3���[g�k�[j�Gx���F�����+�:�d��UC?�u��V[؞{j%�ߕ5��ʘ����;���yp�y%]�8�ot����ߍ�ʳf����Ot��ǫ��6uɺ�7��i]򧩦1�i���]F�S��;)n�f<C���E1;���-�Ե>zGv�ԩ��[�H���zakj)t���U��Y����7|��~Y䕙o4�9-��@xwU���5^��Y��1@�սC ��4t�+TPĶ������f�����+og�3�0Y�>ùF�U�s^�x3<���ɴW�j��D��Gst�Yz��<��x^��^��ZtȈ�Y5�[cvbyv���T�W,�y�E�� o4�c�x/����T��庄��&���{C���u�qڨz�JH�ҭby=ۊ�q;7Cr�]��Ϣů���̇��;���fI���9S�v+y`܊�N�ot=S����ő[�c5i2���x)��� �
٥����w]�[��~�}��~����EU�#��ؾ�*�A�l��UP�zo��}c�ī]'�A�����l��z'�=7s��,��o��H10�a4Gr���ɛ\V���fӵպ{(�,0"=DR/�]מ/Nϭ��0�&j�
#��ȝ��P+������o�:CX��E`��ou孛��pط5�5��C�ۍ�왨O%�"&�k��v�*�Խs�H3Fԋ�ʺ7����pk�@%�,�뼵N�6Z��p3�3zG�r�1k�N��[��5ӹݍ>W���B/c�T��a��iiJ�h�k��,����ɮ��6�w?��Z�:�g�U�n*�x���i4W=qt�+���V'�m�f8n���5N�^���;!� �K��]�{��N���7[G�Dtٓ��<�g�n ��d���恩r�� �(к��DY�!��o���f=�d�3;6��1��6҃'
�����/*�/J��� ]AWZPcI���-%�p�Vs]���L9���Q����!����UϪq��x��x�qLmL��J���4o�Atb�-���.���a#��g;FJ:뒵���z��V�<��^�W���5F�5N���Wi��T)�+<�ͶZ�l��s[0GG,,�U����ʑ����V��Ǜ��qu�-n�*d��/SP��@�V���m�[i)[W"0wi��{�ޅ�0�Ś��{2&�6JY�h�#7^!cvnȪ�"���;��t5-�ɂ!R��ץ\��ʶ0��n�eu�GO%t΀u�S���'	f���%,K�o9�˻�y�թ���N���<�( ؂�E�8-��N)ԯ�[�'�>ɑ��rc�6��>̡�3Y)�:ʔ
J��T6��n~��2�8y��F�"1̪[�]��tr�o1��i�«��Êص:�O7%u�![ư�yqN��8�͵��f�`��mu�-�	�����|VZ��o��E��tsx,�l�AB��b����t��٪��RB^��'KFř�g]�$.b�I�QL��&ܸ���j��זRۡ�s��8 T(Dv�ع}Z@�VT�c[�GN���Z�%,5«,iZwG�]K�>B&��T��#���ifG�d���[�T3�����- }��=�M�7�.�[�V�N:}�;�~�+������	d�V�ܽ0�}�ԹLvsWcons���Ae������K�<�f�z�U�K#�����xc��;4�-ё�]�F�vH������Ӊ�<n�U"!ɯ%�5��5�WOSx&�C*U&D��3�V�&��ks-qrtTy�|%���[Gl8s*�NI�D��5y��0���r�N5�K��nI�r��m�
�z���.�ھ[��{��֌��4=�o%�&�������{;.j�ll�a�LKk��Eֹ]�qڤ��P�\v0���_G,���Ion��GV6����6]*�����hǯOn;��:0�6�v��gy�-�ٔz�������Ό����Ǧ��ei�]�.��Y�Ze%�$ ��u������kn� iF�A:�[R��YF[�7i�$,�,�1�˚�T��z�h��U���f������)2�U�a��J[��,v������;�K���h���a����m�6���N"�A]֕��!�i��iq��0�!��͒<�f0��w!��*�%�:�\��HCS�9�w���ԎgGο�����X&��O�N�l<珗<Wx6�h��eu��J�V�E�=�/{�����/f�l4�	IT�P:t��)ȣ�E!CCT��I���������ׯ^�z����=z�������ǯ�?P?=�%�1lji��,�)�����<�%!�4UǮx�}�޿^��G�^�z��ׯ׬��ׯ_�����i�X��Ub��<�MR<����S��6 �b�((?$�r6�:ġ�f ))��x��d�@9���]Di�9>G c#T�4ST4�P�Q��E#I�f�Q&��
�F�hh�:���i����+Z����hi���!��*���%5Q���<	�T�y�RS�tґ'�<�1C�
Z��V��	�z�:���[�I��&!����#b#�`墱m���<d�lPb
,d�9�"[cIF�45QU�Ic�7�r�[bZ�nd�S�gƑ%��L?2O���	ϓ!�e�A4~� �I��'@�b'>0�_?��MJ�m�I�I�n�po^U9m'[T{-�!x�SMfV��-���e$�f��������M�;�U���`��f���	�c��$H�(@X����
��$1
rA�􁂘NH�D"��Rj'�F)"�%"�
HS("�	P��`�؀��h8a��^yyÞp������p�9�������۳`������,
�Kqla3K���q�YYZ���=�8P��l�2'�=�]>�={-�%�Ȏ�N1)�۫`�̼8w7*��I9\����d�Y��;�C�Xl}�d�P�*j�"�L3��> (��n�P�ľ�N�ڵ�p_y9=��QR̟39^�1�qTײ�T����#���w"�s�6���d�]���g����h2J(���ݍ2#��ʇÒb7@wG���r%,�g�˵�r�ŷj'<�6f����6Ct��G����Y�٣��,��Vl�������^�a��}"��S�{>0o�I������7)���w�����l?[�c/}Ay@��B㵙2C�O]�;�0~�x�ط�<��⭚ �N�b����i��י���޶��/6jXUݫZg��x�Cb�W�V�^�cC�+���gg��Z=F7�銲��r�T��*��\ȎKt2*Ь�U��oHI��I��j
"
�=�i��8DU���54N����܆�mE]k8䥳e���qM#�y"�y�,�5���h�v��^o|���Ŕr�^a��>���=}W��z�+�/�.�R�0�q��[VX]�� V�z6�h}<�wk��W����٥\�(]���2%,�O���_=Ε;�w<���thi�>�QU�H�Kŕۍg��ņsI^�3�	/�=�zEW��vEvr>�p���s˧VP�������KzH����$��2�m-�+�:�gS�z��U��d*ʎ�Ix�Ѫ���zߚ=\{�;�q�:�n]��B��jx�+�oc-�+�N�@�qĨMYl��(G#��Oop뤒�<_���_ ,��vV~�}��)`dW�"��s~Fb���ŧ(vk�S��%c�k[���C��?u����	P>�L�j40	M�v�*r��;�f����+(�>ɝ�4�=�0���0&Uɟ�~�3+��AL#�p��Y<�F���^���C�Z��,x*X
����ߌ��X��na���D�� �V@N�v�IS���A+a�"W<�B����v�;�ar����7p7}�ܼDlR����S3{"�JM�Y�%�߾�>������yY�őa�S��������O��5>�õ���yӢ� ��t�5ǞWv׍z�U�o	�f���335�;�o^N�q���r��up�E����@�6�rNq�yТ�}���?dLb{g����6 �[Y[j�'���+��D?�y�E�����w��,�K�ԁ�ONh������[%�R�s�}��o���������s�O���	nM���X�6�]u69��z����9���;�SdԿ;���Ӣj�<��V�t���~���1q���uI^+�mw�̈>!^��^ L���Q�o��R3�M:�;;�	^���W�a)wZ5�]�U�$U���;ZeNΌ�S�r���!�Z"̇'g���F#�����z��%�9�8�SF�u];�����7S���G[�kl�Hs/>�J{h�T��װ��gٗZ��%��
���V�RSK<x�@���,���ΥsV�*(w4�(vl��΋��"`W#r4��E#��nY3��Ũ<V'��K~�dn��geEs��}O#���w�Ce2�g$�h�^��n�����ڠ�����o?��*g-jT��e��5�K���m����u3����)gK��ؗ�-�:�o����J^EqL��-�mHʘ3����v}��_wyt��s+:Q�7�7{�R�ɲ��u>KubEcNp�l�����K�N����ro�^�"���u���/���}�tٿ����H�������6�f6����Lj���_#C�NW���$�G��7QUmu:���^��h���=Zpl๝w�0�Mß�Tf�{��8�q���Ǯ������2!;�<j%�UߗVP���w~ux��ع�-����edq��3R}�X�޴����g�ў�넮DM��qٝ�Y����z�wl��` Αq��ޗ7��d���&��ɽləAxѢjI�!?�/u��k�!u�)Q79CV5�{4�E[	ȍ����W�34U\�kgS~d�!!3LlM�`g<���k�/wO�k1�UzYx�2�OAz}�Z<T�:��`��b�줟8w�)Թ󬸺���u{�A��д�	�����n3�\8NĎ��k6�Fwk��@��G�y��q�p��[|1������v��gdx��i� ��̠���5���JXf�BuR�h��$��L3&ջ�,ut�&i�g:�����2��ʹ�Y��}�)m�(���[�H����T-֪�Σ��d��Hj̆�n�ގj��/EIՉ���	[�}ŵpԶD�����5޼&kdW^H����Cp�&�Y��:�m��^�w�ٜ��y����ֵ.�)gW���`�m�U���Et����%�.���Ӽ���-���0qW���n@e�%�iB�������ДF������|�Q]�*h��۵��ކ輷JxpM+��<˴9�����Gw�R>�ױ�i'�,�C�	]::��*稀�/��l��RS@d���@|9-�����E<6�Q��ջ�;u�7�'�U�{l:��z�����7{|mʓw�	���j<&�����m߇�I`oy2Ƽ����>�v���T�&BU���/x����ۗ��<���?~g�}�-(;�'\�.�{jv���B0����2G��vq{P7�I��t�|n�Ǚ��ZƦ��l2�y��y��q0�꺈�?����f��}B�aa�<|��]^��Q�E�f�R��¹���%aܑ0x����߻��S_c��p�WX�S�T$	�����S�sf���EW +'�n�b��S��(l�O�6�y�s�֛��:�ð�*��>���Pz|q���p1I�Q�+es�_�u����6t�+;�4���<FSd��ǥWS�=R�*�V����T��j�5�UE����wu���{n�ᩏ�j?��r�Y���a=�w��JXu�:+!�UH�f+��'��7�fU���n3�����m��̚�� x�W�f�g�xs���V��H�Y>�kk��$�C
��@�q*�o:���v�po��zpb�áf �����Z��wd��S9X/l,[���#���4�ӗ"�[��1�h�r�n�`��7���wP)l9�}�ֻ`g1Fs���Z�:��Wk�1�4f�Ԣ9z��o���Yf�ve:�l��f�)��/[�U�PS�2��׽;�ը���t���V�c���d��c�w<AT["���r���v�����utC�!W��3�\(��%S{uwFv��;��.�lǾ��>����s2R��½N�k����Ǹ�IL�/��[��-�j�����z7ZO��u)��SW�g͂Ķ��w��4�����r�elI~Tx��{��l�YiO���oꑸ��������#�I���+�x���\��oU�qYm���ZЧޚ�Ժ��b���bm�Ŝ`��kv�I��}1+�+yy���^��Z��,�θ�p1l�S�BFs�W'b�s�a5��*s2`.�oz|��Ni��s,��ɱ���y[�՚2��}%E?w4ֵ��h����3���{��2G\��g��s��:e�k���kj��f���L�������EW]]϶E��]��|<-��8m��Y��v��B�%�`��*r�8� O�=g�*��.Xc"�Aaϫ�s���&�lh����f��܃�ِ|@���Ȁ�����.�E��~/՞�b}T�键���/�}�QN���EX���������	���zʥX����y �%t/��O�>l��fv���{�G-۽���Y��*�I�]sy"��x,+N,�k-�V	K�?����>���r�~񎎟�\ɑ��]�����WuVq��2�k�2[A}��u�m#�rT��g_�]+�R&�*�UV9]�ǻ����ڲst�~+������*���A^�N��⸶.��lr�V�%�e�۳H��wAD+!ڮ�ܗ��J�����l���3��;��`Ia\��Ǉ�j��t���z;��+�%��P��K�ᮬ�5~���^���Y��x+p'������No6�����C�;�W>�>H�Ɠ������v���H��%j�F֭�͂|��6m�z��P����N�j�y����O�������]�x�F��9���l0�.z+o��"��[H�a�U4�S�l�Y`�����O����<���(��̓��4�i�XmxK�JC��fŜ���c��z4�����	t�v�ٛ�8�ܡl�fN�$�-��s�֢X�3Z;ᗪ�G����c�MC���[|�ָsH�j�F�+.�u{�;C�)����Ŵ�/+"�c�3��N����)UbGE^+����͆�|~�|�7��Q.]%mT�3S�;���g�0mG^FQz�1��xӫ^���Fp�~V>�ˑ�A����߲"�ŕ"���1��d� �&�s����F����,@�I�Ӭ�mݫ�a"&ͽ3V�[���U���w�Բ=�B�_�s8�ϕ���z���Ĝ/�I��ͨ��"T�(%�Z	犔��~9]j����Rԛg�����{�I[�K��!��@u5#WCSz�2�������6��VeQ�E�ps�=�|Z�;�c�ES����RU��68�0�
��Fw"Tt�;��UXN���� ��G���M�fG����G�����esk�v�v�+B3�M��l�WN�KU�qNʛ��̚��*pY�����k�=z��4�"A��|�\��إ����PK�=Z,ߥ�:X��/3��o�t�@�O�N��_��:<�eS� ��%gPx7zF�-<�ɧ&˼��D]!�K�]�Y��!]��甹&`^u٣!���gst��㛐�71����`ӛ��)@���;)2 2�1�ogf����^��ϲ��v`�ݷ�.��9ZV9�L�`��K@eξ��Χ��}��7��U�e,�*u��W�	u	��F#�,�ky�*��N;�q���X�}\P`La�v�6k�h�5� ��jU3���>�J�q�Q��[��L-�Y6����і�	&㱃�Ƅ��Fٟ
�RNKg+n�M�9�I�gg8rު�d��3�d?_	�`[���D�@�Iú٧��-�=���fǰ��M���'��׮:��C�5'!�;�VF�	Zn��~�]���v���������0u��«�Q �d��^z�^Z���P�v������Il]�<�Q�E�P�g���8>3N���w�,_E������W_h�e�:���[Ƌ�r^���95rfty{�'	��s<*Y.V����i���֜),��識�5]N�ܼ;����3���qʬ��)�O��o��x���/�� 9�.����w>��!<�u�tN�+
Y�UN�m�f��N	t�hƨͣX&���4�iTK�����r��F;<�7��c_0靡��x:�Y{F�n�V�zk;��`�7z3�B��	�Q��n���P�Y�ݺ��!lfQ���/Ʀ5\�4&�Y���=e��+��T�A��Αv�oev�'���A.Ҷ�b8!����(.��E�v��>��kpK�d�ӽl���X���c��"ހ��W\��9t'a����w��������]兛9NF #�����owC���΢¾��$Q���z�Ӷ\��9�6�3�@�����%X��X��sL�����H&u���+���AW�����	r^��W5c�,�F��n����]�UaK�� �ۯ�&F���9[���wx�&�1v���4'��B5�|��Fu]Xj�Gy!�t{�d��/f�B�,���-��[Ը[�]h�������F#���4d<���!:ui*�.:k-%�s�ُ>��$��I�p��E�1�6�KKQ�*{	@(T�9�xi��*��N�%����#����l4 <#���8�`̭	0�r��ǵɁ᳣ ���Xܘ$/��n_Bxݩb9/h��Jܱ����\��Ug���f�����z��X�GqK��74&�Fnz�1��˲� �Ldo1�g�.���+���Q�)�j�U&�Pl���Ldc]��s�-���<��)�8q�+%�Ps^c%Ԣ������vl&mfQf�[�o���^���7�Q娛��9C=�)o
�:��X���(W+݃���t[���"�����^�� ��n�*���B�6��J2��X�h��2-�,�_vD;��-��a�5�Oq�w�,��H�n�틢Z�A:wE<;�e��Wp�����Y��Ո �*�+����iJJNg�,���,��ˣ��Su]�U��n�c3 �n��A:���N��qC7aC�2�v�I_9\�sv����,%�eԡ�J
�R����~�ؖZpa3S��\�6��0VĈh�[�!�	�ghKanIJ R�4�ڔ�՝��r�O�ua.ځ��Z���u��!�F,�W�zi�i����kz(X�zwX���T2S�%KH�J�֯�Z�ه>���9��=z��Uh�M`��K���讖�)n�Pt�k"�3�ZY9o�]uݓhm[˽1Q�	$R�Y��VWՔ�xb��:��7�d-Ө�WX4��S7U-�"�ڷ��r��yY�f�(��9����JT�:�'H��K�,����/:f�4B2����]��(�j9������kE���TO�tUCG7;�˸%Aٖf���B��PN��Sn{��hs̲�qm Yl��M����*�V�����9^�={=��(�̑�h�6�UQ� ���j�V��rxCCF�#�ҟ6""�������~�^��G�^�z��ׯ׬��ׯ_����CULMW�4ZOr|�	
�)��`�Ry������������~�������z��ׯ_�G�^�z�������~¢�����9��6 �P�5L[&#)���9M�9�T�I�ZN\�)�Ϝ9�׋�*��E7����ES��QDIE��KLy�ZKIEr�PRPh}˹���z�^IA�y嘉�ZJNY���W��p^`�h6���{�#H��m��>��,m�o8i;'�Z�����/��@Ӂ�tL��5���p"�ܖ�N��MD|�*+O�侱��6C��͍��>�4y6�Uli)��=`<��B#A���Z*��ϻ����Uk�PS]u˓(v<�ƻ�+�h��)�a���*r���t�x�Ŋd������S�Ixډ����y��q7+'f���/�h^��3��Y���f�/����o�V!��f^,����#��'���.�3r[ԟ���1wb�_]�0����55V���t"}�_
�桘�Vץ��8�8h��=��[�V^��]А3��W��)��q9�"�n����{5���/ۯY��cZ��W�ɦa݂*&#3���K!�}���a������Y����I3�)��F@xo�p�+��8tG��|55'�`I�3�&���n[z��{`��\fZTK�9�W�\���� �y����o	���t�g���s����y�� 9�æ뺽�.θ�~&������Ny?P;�>���T\%��0ŧިL��S��h{��J[f���?N�)^���r�:O9e��KJx�e�7����6da����=C�_WE�.�Q3i��J�^.�fN�����������*�y��"V�vD(L��d�n,M�^b3��{��^: �5ؗ�Oj6�d���8v���9�,�?�?b�s�\u�p�5�И"c�0�f����y۳W���>�{���p�mG�Q��-�/�؞+R"o���6��_f�Ad_)��lV���������O�5 w��=`ߘW���U�����Y5��1�Z��:�ò/ǎ�FO�[4T�a�˜����?@Sq ���U}]�*�%%N�kω�����,x���j��?<�� �!H\o�A�{�;�av�Q�����#��2��B����^k8��G�\�R*��s4<�}�U|7�㝐>ņ|+c�k�d���U����,fR@�z%�z�4/��|'#r����@�Gi�����<i�ᩡ��
|��\ܿE�V��pЍ댿[�5G���i'�h��wrG*�<�.�"W;qt�K!�o�|���\�P}o>�(*��� ����F\�ڭ�Ѷ�v��K��"�|J8��mO�k80$!��+zb�=��=T歭�[rK��[ʝ=��w��w\naw�Sy����s+��m8j���Xl�������x�D�����J��f�Nsy��p,��F�nc2
L���!�
ɉ��%X���:���S2�[e�dݚ�$�ҋH"Pȟ}�O��脊��\��w�������<<aTZWRJ`K��\���6W_��E�ΞZ� �Ֆ���q\C�� [<ID�6=�E�n��a�lL.��f#=ϝ8��	�m٨O��'u�V����[�\.�)�`��5Dk����=F|��b�]Ƨ��פxy)���o{���R"���s��;^O����Ŷ��Vl_`��*���z�jɶZv3^/^�&C=z�����=��>*taz���{+,\��s�g�Yn��m�܎ �����w�}�A�M0y����=Xg�]Ί�-���;6��޼���y�#-�T�)����o5�L�7���z��2`<gLn�^o���U��s4YW��
=��9�b��x�`���5cE��8�TZ�\���޽鬙��hx�SM�R�QW��P�0]q&֭��o1,�<��i4.H��#;�xv�����Z�,���~'��iV���~*�ڦ)ԑD�y+�"qF��ﶸ3N4M�[�9�I߫����3(�>ݒu�
u�:���g�(5C-�#u�c�Gn��}PP��������5<�ٮ��0W��� ��wϣ�݄E%<p��7�;�����%��qL��_q����_D�>����{�ψ�qM��_
�+��!Q^%;E5Z˳�;��>bH�f�����'�ݢ7+�R��MZ\�"��v��z� V�Mnx�Ǎ1����"�m�zQ~vvw��L�uʦL{"��ֺbEoS��t��Y�K���,��v]�Y��� �5�ΪY������"��U85mJ�����YP�y&�/�u7-/�ê�en��,�i6�hp�c�x��Fg�.��4z���p�_n��8�t^�"=P�j�^X~������2.k�Dg(���e{�#�٪�|����Q��Q�A�{��an|E²��l����1U���gfL��g��$�0ޣ(��Pg���?	��r��ړ������ ?.s^7��|�f�l��U�������3���{
�{�j��D�Zy��e���YD��[�0\��M��^�����9=7{Տ��];��^�_��
`����YzZd��TЮ�.�2�|L�	�.j�����x2-�*�%��qFHRZ46t���D���圧y�Y��Ž?���9�O�|���߽��/ӾV�v׾������W��X㈄���f
؋jյձ�d[~�y8.�0\�s�˭�[Q��$�ҼO�mMY������T]���N�:��O�|�]=��]�l�L$��LE<��A�g7��ր4ZCzwk���Y�T��v�cT�g��Xlad���{��5{I��'� 3߲�ľ̌��B̙�Um�*�X�x��Q6�1�-n1���tSJ�J�{�Ha�=�S�����nB]�e�Y4io+��wj��i:8�W`���/���N��z}p=f�WJ��6�V��$�ؕ�>W�왞}�6Y�jȝP�^�g�-�F��SZ��y�[����麸��"�9�w�b���u��g�d6�Hl�m�k��v�{�m:���O^]��I�r�;in�~��7��lP��$n3���fޟ�S���]r�{`u@W�j\l��RE�=̓�v���ɞ����X��zm��͜��.暡�*�ݶ�y�㡥�9/�H������˯[*��lb�Äl�U�����oG*����}�I����ɝ��N>/Ga�^^�[���w��e;^~�g�?���+��Ҫ�%���K�����K{��8q|UW���ت^���P�˳�S����\�tcم]�'8��:�>���z�u1)�m���&���S�'��7jvu�\*���YmrϺ��|2��3r�kw��V�V�����^k��ꈋ6= ��
�%����Xp�{2�-�$:o^���8���<igT����֢aY���X'�zg����l�;J�S}�Co\�	:_�5�����oS��T���f�U�Q�@]��љ1<�_T��1���F"<f�B<Y&�c0ʞCY��!��`F[q^��X�M��d�'e�5^�h'���c{b��t���oS�ܱE�j�-��+<�VH�����>����ՙJ�YY��]+�;�#�Un�k7H֫>j\=�sf?^O�%bF�G�a,�R'�w�2��:��28�Y�q�4��7P4r�vN��5���Wq�L��,��xK3V�خ|�	�~�'�⢚��!W(�!x6梱ҕE����,�5u�೛��E�U�qnӫso4�5����Хy�wCǮ`x��s'e�v3�>�������$3KB��ʾ���u�{�f��7p��e�F;�°�q�sV�Q�J����Ug�������l�!����qʖ0ik�]x�V�������9� ���_���
Xt�9\G�"';��V�Ѵ�,Os�㱞5�<��ڮyXc+V�o#��.x���]�^!{��Bق��	���:�M��;@�0�R�H+�w���#��O�x��~��&��nN{5`��U��F�u^�������n����ϔ5Vן�lZ���=��N��;z&�euD��b�@Q8��#����[�����Q��ם�@�c��t��[/�ԉ��riӁ^l9�T۲�b86�mY�6z��9���@cCm;�v��lנ+2,_Zɖy�����*�pv�3KfY�_���Vd����f�@d^ �j��~��K�32.n1��w��,�6���~28�UsO�[�Ζx�j͕,4\�*��NS�w�f��0�Aٲ�x��Ux3�5�"f��O;ctsl8��WS-�A��a6����4p�4���]�KŁp��A�R�]D����e�O���{Q�z1�{5�=��F���h�N�K��R�^�-���i��P����y�T�Pz��8}諻�e�T�_s�}�.f�oP�5�«)��yg!UdJ��.�e�a�2a)�T�	���R���+��k6��Ϊ���|��YO;{��MZV�A��!�����t ���*�uR72O�Ȉ�ݍ���
�����Z�j���ʗ�+�c��փ��*��������6�o��@Y��n�����T��>�����:5xX�Y�z�ӯZ��>w*�{a��MߑVP����'�Ե����Jڟ��rft�n�n��WL��"���i9����W�oRՁw@�(��0f����w2f%>�F3r����ݵ3^��\{cD��ȹ .B�v����^��i�B��i��]4D1Hc��B�Ʀ6tD��'�u��
�y#���Dvl�ftuuT��<�O�C�nz}�� ����4���߮�`ak��Cg�աY�Oo�Z_ٿo���8 B��}[2MQ���Wva�t��@��dM5��u o�tOE��z.]3�	1���-=岦�vUh�z*`��Ԍ�%]�<�@�[���/���G�?�A��y^-޷ܨ��9��ԣ�&���k[%" �3r��;m����sĸ�~^�<��j��N�=1�{��t��3�n�n�]�Guc�L^==F�l��)����A��a�ˋ�5���hq��U�����17S	X0����߈]m��?c���٭6Sh�,~(�yJ�dl�{�F�%�QC�;��|;��vw��=iǊ�
��Kw���q��o3S�E+�W;���&��$ϩ���D�V�Ѻ�7\���q\��Y>?>���O�w���]�����Lr���m]�L�л���}Ƿ�{N��Y�R�K"wVEzջ�S.�����0g��K��t��:��m��6��{�Wq"���ڲm='��{+k\���c���w�n�ku*���;K:�h>�>����U��В���%�gbUfV�ݔ |�}F���,�,+��)�!���`;`I�]�ձ���5|�|��U&�kM�JR��e��_k��휕UsWJ�s�{�_E��S=���i=I�����մ��u��YB�H��v���t[)�S:�ק˷���~�|{^yz�d,Ylþ�Ny�d8��V�\|�qK�7���~�Ѱ��'=O�E�8�3��Q��\���]Wt�LW-�֦ꍛE�Ww=��u_w���YO�t�dB�o�))�Uo��PA}[G�v�oMϖ�����}�7��)Y�!i�P�Bش��7L�nlgq��^-O�v����p�Ī������)l��}MלZ��VVA���م�\��
�>�ُ�+�;�l��w��n]H9�_NmX��}����~�k�.����P3���ާgE�E��z�p29
 e�	P��]�޽�~6D��݋�Y]�_b�]q+�o�=�۶�}v��
�Ţ�X��n %'���i[T��{2�Q�'���w�GS��Ϗ�����<�������?��U��#� ]��DDG�������bT��T�np�A��}�� �A���0Ȅ0���� C °��C�0 C
�(�0�2�!*� Ȅ2�0�2��C(ʰ��C
�(�2�0� C �0�J�ʰ�2����C��°���C���2�0 C*��,0�2��+ C �0�0@2� C�*�ʰ�2�! �0��� C �d0�2�+J��2�0��+�C"ʰ���|� �@!�`@�U�U�P!�a�BU�!�`VV@��@!�aW� C °ʰ�2�2���B0+ Cʰʰ�0�2!@0��C
�*�*��!*�
�(�0�2�2��� B C ʰ�2�0� C�! �0�0� C °Ȅ0+@��2'�
�@�*2��
� �@�
���bC
 @� �8C
 @Ȁ0��(�@ ����� �ʨ��(#���TP�a�!����!�aPBHePB�E@�!�D9�q�Q��Ea��U��HQ��H@��M��0 7� ���2�+ 0
���p��*�ʰ0�*����ʻ � �U�U�U�P!�a�a�a��^���=|����� *$ʠ�B���f�h}�_����@?Po��a�����g��_������O�o��D����/�����!��P U�#�������?؀ ����� �������� z?ڟ�/��p�_�C�q@W���H~c����C�C��	�?���?��o��H�u���bQ@%ET"AT(AP�@�  � a 
 �P �� %��@"�a YP  �  � ! �I $@	� $FP �	Q! 	� $X@P  �T� �eIVD! �%X	VY"U�V�8�E����<?��Q�D�
 �DK�����������
���@���G��
���`������������Ϣ������"=�}OG�'�( *�?�����y���Q E _�!�H~������������yД@^���ʘ?�����|	��0������i�|A�<������?����C�?�ׂ������`>���>�p�������~��������>��( *����G����( *�p�����}C�Re���p� ,S�\�?����>}�>�	>�@W�{
����ɐ?��� ���}_�'�Q�|`��>�@Qu�o�/�O����O��(+$�k%�Ͼ }��0
 ��d��H�w�=)T�)�I"�TW�"	J���)(%"$����IUEPT�UR)* UP(��D��B�)TU�MTQ$�Em�m
m�%lh�J�!U-
��֤��K,�	-�V��Ȧm*`��%SZ��kB%�T���Uַ��RTH�:ԛ5IJ�ET���*)J�k6M����d�j�Z*�ڐ2�H�)f!HQ-cL�� �ѕ5��"��m��$TA��|   㝭�wtw�WV�fXR�[S�n�	��wl�Զ�]�i�6f6b�hVm�ni�˺�kv�ju��W':��M��:�T�M.�\˚�UY��"�CAT����  �>�
(H�
z��
(P�l\�z=�B�tЧy{3ڼ��	&ݵ;��.�Һ�Ym�.�s�]����NU���W���ȥ��ݹ�]�wm��[�X�������m���َ�  ���s�������m�s���wi�ӵ����,���t��-�խ!]Ϋ�2���uV5f+m�i\�Z���]��n鎹i��m\w;m-�Vm�$� [E�h�R
<   Ǣ�f��;��ZhΕխv��v��n*ʹ�U6�gq��U��8�Fn�4k��h�ݭʬ7Z�F��5vٲ�ےJ]�d-�kL��ѡS�  ۽}i6؛Z���N����u-�RV�UFm�l�k��t�-�q���:���M�uj��M�:�,lŻ5��VVvӸ��m6Ҷ�EDP��֔A�ZaG�  g�V��˻*�[U�9wj�M�4��Z�Xۆ7R��T\N��;���Z��5GL�(�mgm�Wmt���7YNԮ�56�j����j����-�(�   ^�@4� f  �rp  ��ۀ GjX � ���
�� - � �1!��UT��w�%U�+Z�)���   X��掀 Z� �d` (�  �  fL  ���@��P�.S@h���� Ң4��D�7�  7� =h0( 2�  �6�  �tp
 c  ��� �s�  hf� ���  ���^�C6զm�i�eI�   >
 ��iX  "�� ˸h V  ��  �Y�@hJ�@ lV  ��@d�E 24 �{FRR�@ ����z�*�<�#����R����L�T�O@h4eE��P  �O��Ѹ��K�^��/#6�vc"h��o��a��xWi��-JڱC���������{�<���lc�{0 �?�lc����1��Cc��0 �>���<�a�q~�O���0���ؠ2O�ӎ��*M�02f��1��*�C�nT�)�F�	�9�1�ԁb�����I�O'fҸ�v���U�i5�n�v���w��q�y��:�S;��5)Z{�q�9��������ˠ2 \ר�,<�h9�VJTA'EKLVh��:e�ebw�Q��2���K�r-���:KtZ:�#k������V�S�6*9W�"�ٹ�ZZ���)t9zs 
�+`Ź�����RiF䱷2�E�E�-b�7-Cp[�`�{LAHGkMRb��lj���N���h�
�c�����ӊ�J�2��
�V���E�6�7�>��37m4`�[�����0m�31<��]Mߕ�,˄��fTS��e���˺�cg�l��B�f�l�6{Ov �a���L`6r�0Xܢ�h��U7����ű���B-Ա���6�SkS%3O:T�<���z�S:ة��0��a�Jjͱ�e,:
"�
2����4����v��Q
-n���HÈ&�ۘ2��x֊�g�Af�T�l�a���D�kW��$�@4�������"�����R�8�t��v-��ܻ:�̓[����YX>�ǉ�_�r�טmB��҃j&��m����H�-��DˈQ�Eͤ�f�d;y4�(ປ�ʒ�F�1@���6���we�׮�T�c7�(;�W�l��YB�jEV۠>j�ەw�&X92��M�Vm���jæp�y).�ӽ�FKH��X#�rI�\m�j�̙�,�@�۳@ͥ%G��֌V�G��y���J�Q�T,���l�j��jV�qMY��g5�6�+�+�>,qc� �����B�X��*��Q��7K���+iZ�ے�	��b�ø�ceU��e2ww1�xdas7]I�#N�[z��)K�mӡ�����Lm�����GMb���oy�9wA��*z���t�������n�K�6՝-��X�
��H�:r�Q�m�Ӥ��wF��[�`t��i�٭Y�+��
y���%�${�{s)�ܠND\f�0a��b!���D��
�LJ.�y��+�%�� �ñ��e���q;����d6�T��j����ք���~3w3`�Xp%� ��F���"�#v��Pk�khI��E(�����`BS�M�6�0��ȑ�l'V�IX� 0V����5R��_f/���f$��zEnKOd�1X�OJ�0eG��n6�.
R#Q�he�(�am0�c]�&�uy4K-޼�`�ՊB����HS*����AeKXR�ϲ��'ര�ͤ�V��S*U#�mm됵�=���-U�V=1K��X�R�P�9#2LH��lm�w��"�P��Y���A�U��Ӕ�MZF<��$�kD)�,4܈��hZq���n���MR�)*ݷx�d��ţ�YAuG��x.3��f��<9�%;$�3/u�w�c`)�RjJ[-[����bN�ܚ��6�KR�nU)�ͨ"�x���z�Z0k��2�1�n�ђ"�uuT�j��pޔ ƷF�Ƿ�Q�A8�g[jl�(�VJ�����4mH^MIi&�R��}J���bH�'4�Y��UCEJ��ѱ)L�括Q)`�e�6µ���ؐ�jiu�Cdh̊+ڊ�L�v��t�ڻ�ps��1�� �]m��A�:?XR�i������r��M{.z-˂ ��tɠ��]fu��u�ă-3:�kj��/@	k0ee�U�+Rж���ǭ*7zStM�z��	e<�(���z���B���Ь�I=��#H�f�������	�PoٺeUՐ�4���@	f]`дd˂����\��M\Em�{OA���5�eMX3R-�9�:�Ru0�*j4p@���&h�",�[{&$�cӒ}��PQɦo�%��a�VV ��C-���2\�3g�U�mѻׄ^l���Wn]��2=�n:{q���-F$��-Y���f8�0��(yj����mln'�U�L�G[y���`L�H���l F:[��;��K���\N�jН���0������R�A,ȵX.��;���#��v�n�W;)n��<c�5�l�Д1���ːmݫxT�����\A#N��S�������"[ړN�S��
eCb�aXR��n�\�-QmB#ݰMh�7k>F�k����x�b[�j^��J��*������Z״`���R��[ۛo֔'+p�1�7!��J�\vZ��J��J��wwa:�`��ZM1�hhAX�Z@7"��
�Ňz֨܍?�C�oY�)�X����L�#4,Z��V�p�[l`��Y͹b�\ݠt��O��6�jV���d�aia��ⱸ���$���Cn�5W���U�Ҩ�G�t�Њ���J(�ȱU��k�$�W�i�v)M�qZ�@�6��b��ܦ�G4�4_�U�Y�v�ȷR�ҥ32�H��(���",3ܛ�"4��
���uѥxu�dC���4։�j�.�LUY7V�VX�o.˦[����/4*�x�'�ER��:z0j�ʵ��4�UVRͥ���i��Sı��5� �F�/wi��t����|�m��q�UcH��|Ei�7��ä<y �V@�Z���(��Ҋ:�0"�V�S�t�=��Ss]65���l�Z�����(&n�.�l�j��1jR��3
knV)u�f�L�K2��be Z��N�F���mG)Թr�m+ڰja4�76�Q���f�d&�mF��]ٽ�hJ�a�����񃴔1Ҫ6U��9��&,�F��zX����P;m�f!�܂R7z�ş["��6Z�t��smf��Sh��6�VnK�u��7O����eM2*C�;�(Ũ��`�>�6�6�D�����By9���y�8iƅe'�Ů�Ʀ�E��qY��Q�7
��ܫ݅)��[r��V�٭,�`��R��%e��w����c�����dmd�^Y�����m�V�9l[��w����B�ѡ`�y-0���S����1���L4��56�]�۶��TY��N��V��"���	��
���5��ܸ͕i0�nM�%ڥ�V��;ݓ.���!�[D�A\�1;�1����NP�Df^ڨ�}�(d�'e{zH�?4�P�M=P�Y��B&��o���𳊃��&�Wj�t2���#�������q�i�����$�H:����K)��Nf�6���!ցg)=���-�b�F[��C�b�иJl³$�����+O�*��nQ��f��y�U���e��
�Y�XP�ݨ���YA�Km�Y��i�T~0����:v��X6�&9��9��F�v=7�)M�F]��
�q���6�3h但����ًEh�FkD��j�K�*m��׿[*�
Xw�I����(�gV;(���Q� �:����RnX'V�(ܣzsi�M��+G
ca��gag-�QsEhq&sa����Yo���0�J����
�KTF�2�i��G���53��x^]J����ۥHZю,Oa�)*t1�^��C/c�.�H&�n���[7)�oqѷu����o�jl\[)�[)�l6��@,���đ,V��k#D�9����Y�M9yV��HZ�t�^�X��*1dHH�H��BG)�	Ee
����'K �Veb���	<�bo e�pQ[{(Ds^B��8�4�6jBkj7.Q��^�sq��6(]��A�����J��"7g&���GC��"�K%�׃f�e]���F�Z�%Y2��j�l!
w��X3ᚑQ�ʽLV@��X�pč��C7(a�#B���,#m�z�8 �o#y�]54l����F,��X��]�04*��S^Z+kC��$s,�{.f	�h(�71֭������n�gQ-&�ϝ��ۻAb�i�B^K�ij���T�|
�ɪ����f�.�ڽi��}��;�*]%P�ř�Z��j�~[OkT���36�wn�b�ԥ�G�ѩq�E�`n�&����j�n��]t�U��i:-��BҀ'z�)VP���Os(\
�ᕭk��>$���N�fE(�7wi��Q4/�D?��Q9)�����*��IS�r�]�8��ߚ�S�P�ЬSz���=�l��r,�iL�ӓH.��ԳK�ѻ�wSw f���ͻ 3�U�]���al:Хe-߶=R�H�CTPMvi�挣��F7�n�(�����8�&�i�o�XE֠&�ekrڵK+$�ɦN�@�v���u��+��j��X���_t!����0�bw���ʼ"��]�֡Җ�����.��Kw�ˉ�+a#=�� BҸ��B:���t�0Y��
�i-�"��̽	qf�5$���l��,چ}wԡ�Y�����	'��2��ҴR����MS�J׷�G ��x�D㊆Z�Ki< єM:���2	�������x�h�.R�N ک��$}xF���	��nc!�4�W2@է&��-]Ʀe!*�����ͧʏ �d �oOcI���ە�_O�ц:
e��9PZ�euv/_]���±VY���.�qeH��m-n<I�f��(V}�FP�N;�)�\�Kǻ�=i!J۵"��{�qǸi����NIYQdP,�L�G/`okww~k>V�F�a��W�j+�"A�]K29d���\`�7B�ӫ�h��B�j4\osXd�%Y-�Kk"����ɫ�-*[��pۦ2��>B�T�x.-�M�.�B��VءY�[6�ZrU�N�Ti�5���[��xvS��m���8s�Xv
m�j�4TX��/�����Ҹ ѻdP/d�+Khn:�1Vދp#��;�a��Y�1寶VB.��c�%Y���3l�tTJ$]a���n3�jI3E<J�i[v��,Ֆ��r�&A�ZB�D&øo`�:�͏0' Z���%n�4�v7l�MÒ�oaҨ�`d������m6�|f�Ρ6�M�J�kV#��E(��8wHDlȵo�^����ԥ��K�Y�H�,�E��M�|6�!�A,M���Jfst�ye�M[4����:jjy�f��V$ٚ�/s���uR�t��-�s]i��B*�lG@h�G/[:�H@zM̦�sM��h�Y1&�Lxv��~iʟ	�I�Cu�R�h22���ǚ�|����(r�T��y�d�ud`#X�MU�a"7rXb�D�c�����a�K�2YB�$�n�3CZ*�RQ��h�
��l�]]\Sn��v�ا���B��Xi]��>5�elU���Ѣ�{{{���H'aæ�+$�����6,�7��2��/vP�Ǐ(��1I���%X��f�(�T�i�A�Gh�8�h8�ÿO�<�{R�I��-|J�m5��M���Vn�n�Xˢ��csD�[Q�2�yQ;-XǪ�"�R��-���m�[ZI�+d�'�1f�4��`�@��[(�rŋ*�ѭ˸k\�*-9w"*���A�:HtҶkZ����7K�	��-Ivwz�^�&mݴ�蠀Ɍ�k6�W�ͧ���dy{�A%(�ڛ�\��n@^Մ�EL���%j��G^8n�����)���El�<!����� (���{[(i�� �Bfe�6��Y��2�̥������]��/~l�����l�(]�e]��E���QGD	fq�
�ˍ+�5�`��=�q��a�nVMM�%͒]ibԬd�K46V*���1Eݗ[M����n�����C������F��M2��&E���sr �&��4qӌ�cS��M �<9����D��*ɭ�v{ 9�b��zFd*�,�w�.���6dB�+�#"yOSr�Zj����a�K&�y6�iV�S2�ѯp7acEkhV��Te�gtC+��m])��ԩ2򞜶Z
���ldzj̠���ٓQn�A����ܵWVM3�^2:OsRK7T/v}��� �	�M���U���2�.ar�86 
BΈ�7�l��n�j����o��t#����YсaQ{�21�ڭ:(bo(�Rf���ϕ8���M�n�T�aG�%\����A����6î�ۨ(�o5�y��bQ�@Z��7�2Y�E�o%��4�P�RV3�P�q虹�UÑ+�[t��	�]'�BOvJʕJ%�Jԥ2�յs]2�l�	�U	ҦM�r,�S����kІ-ћX��˖51�j�m��y��#��u'�M@�N��d;n�ö�t���4۷��63%��m��`�HM��ݵ�#H/v��HZg'���Y[z �;�q/t��$0- �zB�)Ր�/�#q�KZnaZƌ�kXSUomS�"��$���wQLL�`�w��f��3H�H-DUn�� �l��`�JL��m�����࠱�C^D�Q�[�0b�y�gv|7ph���Vð�Sx��RTv����\Մ�!�kdyCH6����R�Ps2KY�Vf�M䒘 �5�2�[)*����n�Y�K&Y�VV�#���c)[�hQ)�d��T	�#�r�3b��M
�FM�t����B���t�J fuҏ��f6�:X�P�*�-	YN�L��їMeE����L,Z�����[�86GH�Te�˼nX�.�g���2�e�Yz��ֹeS�@���B��V$O)��M�B�PB�V�GZ�Os,ܼ2�c��W��cQ�ג�̛�K�]0.^� ��°��M;���pɖ����n�޻�3��Q�L���	oM��+���=h�[�MX��jF.:W�8��ɖ�lWZ�&Շy�v�����#�1��qj����'OT81�bcѤkO�נ�4�
Gj��H�ۊ�U�p�)%2�$X�3����^_��f���`��C���L�W����-U��^�����t�_�tB>Av�چ��\��tf�����w�dU^�+� ^V��Uқp"-�����Jh����搬̿cW4pc
]խ;%X@@e�v��v���M����6��,���oJ�ƶ�:X����h/�����BӦ�Du.Gd�$E⁉���*vy��GOQƁ�1F�;���v7u�1���g3e�]���GSJc���>�\�^�4��r�9u���t'K]�cᛌ�勯9x�����'��-i���2NUc&+�Iw�9��ju��!���p��U��e��@�]���o�wh���������Wd��:����WT�v]X�[� �;���$�9��w�,e�\a���`i�/�Ӭ�b�nM���:z�]�����vW*�9��j�Q��_a�yנ��Q lu��Mj��fn`r�h���͍�kEm�r���'Jc�NG�w�����Bta;4�]��x�a�5Es\�9��{I��p��Q�8W��_K�p�%�;P
yϓ�Ԯ�!8��Vu��y!M*�,���#W�0M��C���z�w8'iX��ܾ�8����k��n���l�mm���{�6�kP=5>3E�s�S���R��n�Ꝝ�'�q���r��+�|���b��A�7J���ؤPB��oFP;w���]��LV�=ֶgz�bf�X��X�]�M<����H^�5a��;�-J���`A�-��M�3�&�I��W�t:殕��Ú�Q�֎|Fm\��vK=0u%J�R��-�u���Ĳ%:�4M�Yʙ�UVp��;oh���(�)� �Ն�$����<��v�7)1��Nc�ޫ��i��1��D�g
�u�mtiycpA'�.�y��8v�X�o7V��Hb�-�K��r������NO2��P��q�Ź���K;�P�Sb@Mb4"�@�l/Qʓ}�N�2�q��GT��ڲ�,�E�B���;T@+N7t:��\"�`��0B���%.�[�d�w%�n�EC��!Lݎ�)i��v`��9�+���&�z�	n��q���!~yNUS�����������m�8mM
���.�¸]c#���6�����a=DDP
'#[�� -t�س�2���WWD��n�u;�;��
8�t�X/
g�֚����	eM�TyCMH+D5}���B�'����oA�Z�vG��;�뱾Q��c�K�ՍP��P�2��wuJ�mӹa�5].��4:P�V�]@�6�	��J�a���G��>��o��.Q�p�2��1��j�״�`4/�enK�A�v����1�sK6󮂼��g3��+`ֲ���+{������T�����ǔҎ�*z%� 0<l/�;ٺ�^���u�~'i�t��Q6qPa�KμV�fmF�j�����r /�qg�2!���Rzڳ.���r9�����f�|�Y��Z{n�euk�ܠin�V�s����{��Qh��K�o��L|l�yǡC] �-�8ev����c�3�w\�7E܂�U��ir���[�G�>f�ZW�c�@N����;��ӡ�`��N]����+v�47���:��^g[��':�um%]*�T�oX�8�C��~�zeK\��j��n��	���47��nE�������H���*&�=w���sv�靾bKQ�
h�Z��[X�]���%n0�=+��DwqC���_pO~ޕe^�u�ui�ؕ��j�p@�;�l]6'W�zq
�oB[��'�Kk�԰i��4�9�cv3��%փ<�l^f��岦��tҝ��&u_}�s.��w\��}��G��-]2(a�d�iw�U��3���J鯭ۮ�̮�����Z-旃	�����ȅJ���Y��U+�#�7�aT�{�yK�Y�gu���t��v���zߊ����m�A�Ru�4��jV#��u�%���U�9��J����L)#��G@Ĕ�Ω��BNԑ�y2��y��m�v֤7���x���q�zz�˚�m�b�Q��E����fR�c�t��)X/p�Jok)����,c��M{�g����j�d���.�c���8�G�~�Z|7������OHgc�g^tu�H=D>[-ʸ&^2y�Q�J��d�n��e��X�i�+�t��l뙔�ʏ����Y3��n3N�f�=x;�=q�cZv��B���]Xż��볩a���<�ӫV,��:�ӆ�͙�.�Q=y{�%[
�>��Ҳ�Դ�^�궥�"v�P�.��CM�m�v�p�|�Nd���V��ؾ�g�1��>}��ip����2oq�4^�f�}��Ak�c�53�X*�v�E
�U�Ԥ�q��owZ9�慵3z��L�`X�xoౌ�i��T�w2X��~�7<s�q�pz���	��Z�9B��Z�8���ԥ��1<9|�*W$�]]�_qo58�L����{K쾴�_TL]B�(��4i�q�6Cܻ���������u�+kr�<œ:[�s��)�ǔE�S��4=��9��~�]���uufk\��]��^���y��fƬ[���Zq
�e�VwJr���җv[ĮvKu���� A�i&�����iSѹ�}� ���,d�ܑ�g��U�ڤ�I6�;�фf�w�yxr�6s����⹛	}x��V9��EN�q�fP��z�/e�7��ͦ�	��3)�yu݅��-�}=W�Fs>w�M��meեj���ۃ�����h�&!�dyJ���B)�:�����U�#r�7r�iޚI�S=�2���tc�L̚t<H��LV��N���nTLcF��%ǫ&!��ř�k[���L*�m)�qX�ѓ*vҽʰ��{�Ж���0��E�=�r�@0{dB��v,���4��_i�Pyw4��E��˽Ȗ�ތc�Z�#��{,���eCb��7*����P��F�c�e�H��A�(;y������ jd��h` m䫟.�.���^���moJڦ�q��ʜ���:Y����I��8�L�a��wB9� ��%w�_Et����a�lňm`�N�a��mh����� l;ǜl3�Ƨ �oiI��&쏶������B�"���O�ʔU�P��({�G��a�uizQ]���[S4�u/�ub\,lÏi>���([���Jwy�襹F��Jk��a٣�KG�՝���/95��8�G��X$Z����5��U���4���G���gI����`�	E��~�
�9%y#7��pm�%�E�͒�^���5�9�A�cz��&kjA-<��ZͲ(�����a��e�Uعm���F�t�݋�Ұg�����Ikp�5�����z�b���fjEjSz�V��z�jػ�S�,�5|�]dr�:�cr���0�u�M�[C*9j�5Rζw+�ٷZː�11CwvD��Q��sB��T��6n�Cr�K��^�F8^U�B�њk:s(��\ﯰm��������o%��f-ĸ���&�����ዶ[���t�ή!i	����.��8W� �i��E����y��qT��ʕ�z�b$(JY���D7���w��4���8,3�y4O�>)	�\�|�^�cc$���+|�B7�eYT�F�ً�U)u��MP�X��.��!�D�EZ�	`f���<��[�é���C���M-z�v 5`l�#sA��u	\��
��ނ�q*34�$����0�ԆMQj��-r�{��<�K{q���1�*:���)F���PL�)���)|y�N`]�^s<�ĩi��zޘ�f�lD�4o�ge� �2�X�h�SWhc3;��i3�QrKP�v��6%{Z�t$m㕝�[c7 �i�	��+��PMj��74b7�V�P�~�ɂ��p��K�n�)0�.�<m�w��wPouj�J�q�:�ݱ�>��F��m��YC���q��j�-�b����%7�!V�i��(yuZm��k X�MXwA�!a�P�:2�c�ե��:*�i�b,��M��\
�̥j�)�_2g殞V|{eJ3&X����d�Lte/9+".�L�J6��"��lU����
�j�n_=�5����#��.�*�u�%m���vu4l靡�0r�k4�2�!ݮ���go)�ԹV�����F������<x�Hk�29�l	q&����3���D�nRx��kV�qt���Sw�˂f����Q�,�����(�;�ބ\�\w�)�FUe��k�E��x�B��i�B5��c]%���m�#n�o]��*��)$U�/:e���K�U��ͳ40�g�^qOZ՚�:��m�BI]�بa�/m ������2��N���H��ģNmJV���V�أ2��n�G��#�<1�{�EH%E.����N���7Z挾�����N�-[�*v{w�o��`�N����,	��-�G4�Prf.��T�?~�S-�)�>���q��`#����#l��,�t1�l;s���t�����f��ʍ���q��3�t��=�7n�=5b\�k麲��b�;¢��O�f�*A�h�9�*��u����DN���82�_�[<`٨�p'zho�����>�bh�$��]G"��5��.il^�A��[cu �9'FDa�� �+�]nT�ͬ�Ev���$���R�A:��7���ڗ%���y�úGN���!5���TX�}�ڧ �\�)f�ă����zH�#��wԀ�*g�h{`H)�W!@�����,r�3��]�h9BI!g!Ž7��r��%�XE��*r<�n�]��	�]8�."�9ܢn�i`f�L�"�D���m]LP��f�Pͭ���@�l�w-�O�n���K0��t�9:�}L��z���K7�+��*ͷzu�>�D'!�����E�kMeɾ�j�1���V�n�&�!h4ŭ:�_׾2缙��p�	��ӱ� [������K^���B�%�0M2�ة�k�do�M.�����*�F4���Ȯ� Z�#G���K8��"�����I��
�KQ�R�^�C&�gnӐb�A]2��\�;Lb�m���S�]*1��0�d�Rg5e�zC�q��m��S���?��<Uk�嗑J�,��ʇknp)�δ�C�tLVkp:����s�M]ua�ڼU�a%��wn�WW��T�mvt �|�:�d+��,`��4oa,"�%A(���:���Ŋ�A�����O&h8|ۘ�X~��KV�-��bX�п��mu�eY�HeNR�����u�nfTS�7d��7&���ڵ�sb�0�n�X-W\�P�?���j����-.��"����܎�kF��k��M���նH���96h�f����{��J�$
ܢ�"�q3&]ok<S꜈���uqh���[�=BVa��K��;a�/�ђ>�	�fuk@aέ��KO#�H5�lk_mh�|@��K���=ۻ2��c0X� �[ѸS�ڰ���*=Z�u�V��Juh�*��t٘t�����S_=dfY�-��Qx�n��Q����3��n�t똫�����On�}d�W�)i,a�I%sjW�r_0��P�%�y��K;�/t���B�Xz�4It�������\�YްԿ��{\*���%�����;�]_2�Go1I��+(7��
�0����8���x����-ܳA`��ࠊ�E87ƕ������m��4�h8w�]�ER�u�#W�r�x��6y�{�W�䱌��85�����E�ͽ�hY+mR�:	��������s2'je�a�7Qb�/=-i��^v����qÈ��V%J֚�(t ��v7t�ws[YiK�zb�f�s�o���^���B�����Y��x� ]e���Uʷx����+�����SJ�b���)(c�
C/�kl�N��>y�'Xȣ
�:���녳�>�D�aײ�����a�F����qa˸pB��b�y۳wT�p�\{�?�d�Y�eA�b��;) ~-h�㣡ƹ���殁�Wq캺�}BU�P*ۆ��]@�ep�"���$��ZW�R#	Y�\�y]�h^�yS�̗�J�Dؕ���BE��}$�T:;3�q��ô���)fsN��L��;˾�z%��f��[R�K��}ǭ!+{Y��\�Y�N=�;�x�<���2,�fm�W�S���kܛY���wKZ����3j�s�iй�dc(�ڵz�x�r�R�� V�Z�V�C ��rM�6��'����K��^0joD5�:��h1b��&e������Hk�ls��<3y�
e�Ջkw��Pn���6�KS8���Ų�]()���-�|ju�^�Q��%���4��Mmj�Tೇx�u�j�����r���!
�:�sMY��|��	��ff�sb6f�3�&�h����['s���S��b���_;���-�E[ �ݫr�9>μ���\���!}���"V�g��Uw��V�-P�e��e$*���ps�h���P3v�*Pf'�H�p��/��^���j�}�-�{aR��1�,�ڲ����{8�ۋ@�K3n�g�j]�%����/0�/Y����ۢ-��D�Z��]vR50\d�N�n��V��������+zm>���$�{��H�kQ��A���h��:��s3��;��HFC�VJ�qL�N�:�.��$�VZ}��ж�J�l��q��£�)Ǿ���!f��h,���o���R�:����˓/���4��̔2uI�V�/;6��':_�*�k{]ҥe3ݡ�취�9�v;q��S�(�'L� ����׳�>y�Pu�x�>�YOs�ԝq�i�h�CH�ۜ��Þ��zR(t����O�l����tRCj��z���뀙7�O�>   }���������-���R�R�;%8�6�"����坴M�k6�A�P�;k�Mv�i\@��o�����1�H�.u�	�{V�;E����4��Ƭ�ˍ���pA��<�� +����5�s]�u�7.�G3��m�{��1�T"��Η�������nȝ� ٙ+��λ��z�w���*���P5����|"�v�淪��.hJ9���u��v�����!�;��j�{{U���$�plΩ��Z�tgm[����9����V.7��\q�L� t	pjPhR�_jw9a��t�LeZ��vVʫ9U�U�a����ԝ�6k���,u� �ܐ��`n�a�7�XFP�F�r���m��8\��]`D���&`��#1��լ�;x��֭�8j�r�_u$F��FV��g���V���z�5�u�������l�s�3���j�X7t`{G�0ܻ����9��"��;��x$��TxeL�GVe��-���KS�AƳ���Y�ߜ|Wt��ww��(������ң%�p���Y�MP�VXMU�IY��>�MK�0-U܃�Ĵh�Xf�wΦ%R�5@Zˮu�<��������锕�.�]��@Ӷ�g_޲�D��DL�8*�p������x�Iޟ�Jh�״�Z�rŷ��8�͸Hm�|�c�%��Tȶ�!:�=4Z����HǨ�/t�ԥ�YxC�LlW�i�Y3P�X�1���ވ�N�y���F����L��+�Zѻ��]�R�7]��G���kv�U2;�4�Kf@l^��E{|��FqJ��A�.�-]b`�:�li}{����ř���^���+��U�5<j���9)!}:[�%l�.q�}r�����w�m���R٪j��-��J�,�d�t�f��[�{qks��٦�t�,��[ V��Yk����Y]!��]ݽ�R}f���k�M� �TԢY�iX��+�<�˔��eqF�t��E��K��\�ne��(_-S*�T+Gŕul(�K��{�{݃�ƺ����
�y�T�	����Z�qr,�|e�i�Eue!�~���ok1�)���\]��O���0;ʝ�s�W7��7Uw�Z��ڼ�hE4�.R��Xrd']cS��_�cxӏL{u�8��k��U�v��4�Ppb}d�7��qU�_u����y�#�8U��J|��������8EG�;�*���W�DF�]�r�1���/q��-Kn�l[3b��V����s%��1bivD!5w������y�.�[��i��J�4�[uYQ]\(�p5�84��w�*��V�@��K26��3�b���%=�^M� ��V�Aف����.U��nhƳ#8��94�w�Scsk���S�rc:�@����h�C���V�-�8�)�#�J=��c�V֎���ü�vu7|r�7�t�gN��2�ɏ��*�t�;;��֬A��o��yJ\	�)�e�Dպ�zx��n^�R�Ň ��P�Ѫ�B�����˫UǊ�l�ue�i]�%�޻z'K��w��o`v%��%LGZ��հ��:p���N:��F�JK�E'�51�1���.�����
%.#9f��ꛖ`���z�;�
�<!P�����J��r���T/�mS�]+����-pҭ����UΘW��^T�"+��/�jط�����#7"ms��׎����:��wK{���؞dK;��x��2�J5���{d��&�u�.�]#Yz]�i��Y���9vr��f0uN4��j���v����]AIE��q�A���t�K�6��������+M͔�U���`�C���1�m��,�(�E�N� ��6�9�q��2^�/�	���|3���,O����������ql;��d�k�k6�s-}��	�����UDV�7��z�!��������V���3��S�Kx�j��r���� �.��{PW3ΞdC�=�n�u+k�fP�Ӹ3D겦Q�,Nm.�� ��Ԡ�Wl�ۂ^��Kǯ� �A�ؔ��r驊���7�l5�k�u����;�˝^������v�����/T�˵��+-�X��d��s�(�w��[�^�m�<>���:�C��
L�˧;��u�@Z]��h���V�uƅ�s
b����o�3������
͎�ĎW�қj�E�-"oW�Md�R�Z�*#��r[B�L��`V��p�S��J�Xr0&��$,3�]�=����Ad���}���'�J.��W�{N��L��� � 58f���EՌ�ǘ;~:o@�T��{Z�����{k"�J�)�O�wL�4 ���Y��T#AE}�u�˭]�����Lr�0w�)�b�W�[/��ȗ*u���pk���γ������p[� 
�k,�P�we
��I�����WK�+�s��A�g�Sh�˖O4{������@�4N�yl
��e�̾�ݐr(�$T.�N�n�4��]s�3����#uUޘ#*P���B��q��ڻM:�XB7H�f�N���RgEp��1J���g�?����VJ�B3-6􄚻��F	5������H�&I��	�
��eܹipW@��(V6��7,9u�������r��	��駴�כ�{�ƕ���VBتVV�G�{(�̫@�=J�h<�:���0��1���"�V��i>�Dc{�Xn��j��s�sv��k�7,�%G����:�N7
b�8dP�r���m[ټ��eb[���Jˡ�*}!i���Z�vU��-�WJ�����QW`��ǻ��y"�tS�G+���P�/���.�7hX-S`�r�OM�eZ喕���r(�o|~�:�������A�P����V!��K���,�4���I�q���`]]uL�@��G��g���:����8M;2��4.��rW,��F�[�g�Tk��Q�F�Vs;��x��l���E�\�r;�S��_!��N���}���NIe&qJ69�NYj�'�:p���_7�uw&V�!�a�M�{�lmB}���7�V�^�Ʃ|S���O�[�r�qӬKP^"��;h���@h���Dͫ�X�0���oԓb�S�Sv��c}]{H+�!,\R5����,T�N;��`3v�IP����Շ�ݐ�oO�et���=�9 a�y���<'Lұ�Ӏ7Web�G�(p��w���9����hJ/)#m�;��I�;a��JK=�����L-�V�'*8n�\�V%ECl-�Id
�h����s���f�{���g��֨^I�f�W�Y�Iۜ��m�h�dK�ko@f�ݸ�̖V��Y��E=����+���3P��FigO�z�y:�,��G�0g��d6���]-�����v��Vƣ��xҘS��,���3��I쥈ɴ*v��v��ڑ&M.��嫫=��V�2Mc��K�͹��T���-��s!~(2g����87�o�J���t1i{�(�V7x*fL7�4o'x�5��13D`��\���L����V����n��]�gғ%7c �o�̽����ح�+���ʵgl/;ķ-�̭���g:�Ч!�hd�7E�yyB��GLo�$�py��Jo[Z�V�	��vӼ���ʯ�(`n���p�NV�e�	@�9�/,Ů�6�Xz��r���Y8�z@��O�L���&�a�l��	���<����(m-6�k��Y)������ �5��\=ѓԫ(M��(@����l����o*�^[oj��I\`ml����7]�":jt�ãyu);�F��,�j[Hب�VY�c�q3��X��>m��8�xv�����Zo3_'W�+��s"�o����Q�q���L�.��d�m�:N�2l�{I�)���3z��l�|2� �+�Go�J��[�d��(�VLo��2}�ܱu��(J擏Y{B�m���pO/�h�@���ށ7�s�ݎ�Q�9g_k��O�)]t��f���!猺�B\t�Z��9oUbl�Q쀿P��`�ju�v����ڪV����e#��q�X��<��v�wջ�|��~��9
FM%!�`�Ćj;z{:5b��aT 
�b�Z`�[�&v��_9i)�֯�laIc�����ge�LO3yd(��L�&ٳ�*�����Юt%lܚ�Ԯ��D��(�[��j䝘6>��2�	4L�a�0��Ѫ�&e=������QCwq����^<k7$$p3Q��|�M�*��$-N�2���m�S��VY��Ԥ�e�[zkE������7�˩2��=u�A�z�ЃA�v;��\Ҳ��OM��7BVՀ�=J5�N]��]�R�c"�Jc2Ms��F���C���ih��;���oq2ܖ�oȮ�w���1�7��R�͢n��w*<ViL=�Hi�4[Ѭ��/;9,��Ȳ�yԩ�ai�i��{��={A�"�VJOp�����S��o��*U��I�����~�d4�Hb6b�52�E���U]�d��}Q��5�"	XG��8�����J'�Fn/�k�hge�+�/
���1˦lC�d��a��$��]����Yp���6lwQ����Y[O�M�9�h����%�Rַ3���[�a�b��hR�]r�ٷ�_s �cn΅������lq����c�`"$�4��J��u��[�p��Z:�3��R�;\���y��(V[�t�o9�=մ�z�2�WK�L��%ԣ��3�wlg��#wC٢���Ʒ���D�C�w��3���@��O'jl�&ۼ����"6y��&���R���b/��-5r1ǉ�Tz�r��O��Aƶfޙ��n�7��sl�;TG~��n���y���>g�\�E���*c8e;05b�7���|���͍&uo9S���z�<�HK�وjK����ؽ���ʼ�tV.�{5�}�����R����Y�� �xd�0�Z;�kU�.�Z���
Sy�\n�̚4��I���ی��b����X�l������f�f����L�T"}>*�o�E֮Դ��bV���٬T���tKa�xn����v��:*;���󕭸�hj̥ekB"�Ն�t���ޮ�%p�J5|�+`��L��K����j�&sz�w�N��VQ������q�	��7�s��ά[mv����L��~��A^ݣX�4�VD�8a(��0�|�2Qغᅾ�\77��Z7���z���c��K+��m�7S'a�0ɛ�5h��j�@�Je�6[�џI�D`��evt�+���]u�r�#��,r(v5��%���5l#���]�o&b��^kn^�:YP�����Q�Fs��� 5�5o�K���>2��
���R�N��Öͤ�,cs[\ZZ�Z�@KD�``הZ7g����T��2���/��t�΃.� OI2�ٟ ��y1m��mM�� *�d���hYX,ժdIx�SM�nʕ�>�n�b�t�n����⺷O\D�o%2	�F�̡�sԪu�yh@2�:|�_<�3�G���B����4	6�U��gT�6[���Lcv�.��R��"�AŲ�V�$�2��s;�^�2�^�(d��sJ�E(J�E��@ξy(�=� �!�ӗM��]�3kw�UK�rBq����g���4��7�h;� ><x����� e�U�H��Wl��k%�Jξ3W��:ڎ�<=F������H[�&<B�\h����(�� o [��aF��u��&����j[iL/]�f��}��vP7�ԯ3'��7`5��i1ݞ*�	�x��ߋ�c���R�x��|��K9��IL�����c}�w�j�ʙhQ$g`��[���3�b�f��p���r"��K�)��+S���҄ۃ]�՘f��_Q\_|��B��,vNK�/��}+J�ٌ��q�@r��t�������}74<9�+bmmi� �H6��W��ӚjY]a����h�����?�q_-�����.^,B�i��Y�Cu��^>�� ^�t�p��>*���rT\[l�ӫ�ڰ��R#<c���ڧmͳW�$^�uhع(��ح&B�h�J��K�Oc���]�Ī��X��t�9�*R۵��0�}���g.q�9�'+5y+�L�-vn�	�)�Rƨ��\�ֶ�\��oZ���l�ݐ<�ຐ�PJ�Yw��eƴ��2��0�É��E�Mb��{��@#�����5�4z����h�q����� �8�X|��������xE�W���H -Sϰ� ��eg`�:��(r�����y��;��3�X�q�a��Y����	��6�;�_'ڰ�v� ���o�n�Z�-����7C#�%�[��^G2�<��P�|���Ȝ�Ln�1VV1J�SƑ�f.�;����e�*RwkH��9Lkq�{��젔�}W�*�Y��np�vS�T��)٫�qo�6GK��{���AJrmty�ܻva6[-L�	�`�S3��gSx�o�1�Ռ�=�X^iԩ��;�g�U��np�2���"���)vw>Ƞ��d!^�L���]�W]Yt��]eX��(@�9�k��E;�d.��C_%s� ��|]��/�K0�--��&p�bS��t*X�ݢ裫�i�3���ۢ k�㚄ʥ�ՋJ4�L�,�G	����V��aF�b�gE�:�N[٥��e\q
����~Af^P��ϸY���3��r��Ư�M�#� ƫQ_2�t5f[fΗ$�ޝ�WIe�뽞@�v�"Mn�g�o0,�<�tIK�rXv*>h�B�]���@V��9�`iy��5�!ü2 �D���<%׼���$�K�|>��}���0߻s�j���E�ڸ\c��������\8���gڷ�`�dk&Fֲ�Y����,�,���1���Ϻ�@U�G�x*�*�lr�T�����}��ut��S6֭#rj�v-�x��z��IɻF�*��+�5���\fޭ �qw� ۃ6U�A��yn&n�ks|�8�l�U��J��n���2�nn���t��"���N]�F�>|9y:���m��6v����b�ѱ@�����ً�����)�ג%�8��l�h'�r��o��ؤ=�z ���.��DM����w��՛.�=�|�ܘD��Ӧ�����R ��ѿ�����e
�h�[�(�&l�|4Y�n�!:�n<�6�q�����'m�n�*h���$��X)����0�2�_���ޥ�6�*�P�(�m���zz���_�жY��K��ۉ�T�(���zЖ��+F�VjH�<��wݫ��RM����;��ٳ���{Z�_`���m�x�J�c��
����l�[<%���ћ�w6D��I�M����ܱ�ȵW6)��tvi*��T74z�E1��g�[�]�K����;��2�c�͸kvCym�#����4f����@W�XqJ��;���l]�wyQ��T��Uo�M� ��u�B��*�+(Vf���V�j=5�t��;�	 I�H� .(�(�������^�Qr�P�hr�PUQ��YD*��b"EB�̪
���r�yK�EQjʻ�k�6��UT�Y�PUEp��q��ԔA�c�(�&I%UȂ�Q12
(��qD�(�E(��q��p�D�XE��')ėe�/-����9�@�t�"����I
�s$"�UUp��f�)��8�
"�+M�!9J�IIeˇ3 �@�TG(���L����EEr��H�8TEU�r�ʯ]"�dDs��.T���!�EL���Z�qT�\��9QTQs�8Ȃ"
%H�f���r(��(�/+(���\8DQ�PA9hQAʓ"(�"���EEr9QZ'/"�R�h	W;+�\�w-	�&e�9��"(�U9h_Fo_޽��������/2�)�|��8nh(�UKw��q{�*���Ό�+��I��N�I��L�b=aV��H=Ӄ���_���ྫྷ���lKC�e�Ÿ�X�ePU��T��m�R�x��^�9�K<���y�i&a�'�z��݊���KE��<�9�Y���u�z��3��C��x�ܞ{-nb��(����.( [��λ��`�
������uk��9�9����b�jؼ��c�g \�X[�6�m��|����Y\_�C1��ȋ����2����#���U��&��`���rk*	�eN��A�+Lϴ�]��wy��n������4�i���5����u�BK5>�n'|fJ|g�g��Ĭ�ǷT����*�H��=���G>:���I|ªf
�9�2��/αׅ*��Cx�w�zh�b=u�F��|v�c�LO����1�o����VN�Ðe��-r���`��.j��)��
ƕ��$�k{)�K�h��>�i4���ϒ�:�&��I�G��l��uohA4�����MN̽>�T=���9C��4�~����X�n/K�FD��H���I�ʻ���P�ŷ�z�K�F�Q��m/�e� ±�'F���X}םQ��)���]g�����r�51s'�FY)�k-��u'z�
����}up�[�4'ƟWJ�L*ނ^�ꉰ`�Sjbn�h*!N�zBѣ镲���)��u��f*�O�4�r���E3�����u�����ے�}�n2�e���+vP�M}y]%^mB(_Vb8����k��ğh���ļU��}y�J�n�y���|�����m|�e���-�k�4�{=ޑo(Y��x��v)ã9�����˪��e�]牁N�U^ā쾋 JE����(I���"�2�v�M��Ј�dl��X��1T��>빇�H��g�>��Z���9`3�bi+/Kܑ��t���Q7��٪X�]��#��ޔ�v� ΀;NO;��4�˦G��I��z;�-�}9��+�:4;$��u}�z]`=��,����8�w�v&u�v�]���������e3)Xz!X��T�8]�aβE�}og��	��֠���~�R{R靱?<ވ/}Y�,��ECK*j�6V�W𯸯mq�z"a��Q�>^�=T&��4��Ԡ�z�:����� ȱ׬���8�;�խ l/ƞ�x�vab�&SR�8ȥ��� ��U�����P�*������-��m�c�MRĞm,'�l�0k�j�o.��і��]�<�+��.�����j���R�X�z:-�r���R��ö��T΍18�t���v��o��Q��\�S�h����2��M4�{7�@x�{d��5R$u�]]�ı�î��ȋ��p��Dm�J���V��ѨU}VUtʴ�ܳ�Ι����۷{��~��a�y
w����X��o���V�yT��z�|�39[F�j�9-��ym�W�����ŠN����5�a�$^��wŏ1%����^�&E'��n�s<��*�]�:�6�o���s^�uj���r�.���<�^�tn5 ~�v���bI��O��J�?�\7׏���W���}�}\תe�
=��c���S��Op�zZ���a�y���K�@��M�u8�m�̭���J��UY��H���n_��Q�=Xd�\��f�Q	܆���xi����$���A5��E����.�7ֳ�bƑv���OB{(Q������"�O=���N�=/'N��U�6]�����1�)�D[2���E�X�5!�*L�+�>�����'�#�W�Z�x92g;���:x��ǵ����JW�'^�@K��
������(�˗^���e%J�&�u�-o�	�����Wn�a�b����Vqi�	��o�e�è;"nfT�k��(j9�Fh��sl�8�ԧ�qc����6��^	c��0���<ۦu�^�Hk	��f�1�����y+_]���^�P�T�] ���f_�p��G��-
u����K���:��TN�Z�m�y�D��Σen*Ye[�~~6�՞�������{�b�
��Y��P�f�[�t�ڕ��EK�P�V�p\jSK�r�*a�����CU�P����{ks�8��=};[i�{	��^��ǚ;"���O�s���ը<ꢷ�V�]^�~�٫2>�k��ф����3m�L��b'u��5e��	�u��z�C�%��ˇ1q��q�e��`�����m���[�5���T��Πsz��m���ui�C�"w��D7��;��K��My��W��'֟����S�}+������U�c�~��e�=p�H�6\����{Ӥ���W�C�Bb����9{��$KڣxD�ݫGus�����^�يWU���r��e}��f���.hܤl����{�&|�q_ު��9TE�H�h�\����A�����7���}]��s���֍�	W	���n���S��_.��iW��K�T:�h=6/h?k�q���C_���]�ߦ�I�Z����}���S^�Х�,��4R@�I�,�f�ֳ�P4�r�������V�k���:Ϋ��.�=e�M9z��d�d�/����r��yBGl|!��y%��sL�*
ƯS'�M�Vp:�`:І5�r�)G��=��o��`S˘�.�>�iv��&Éi����S���C,��۬dUH��ˍa�0���;����9��R/mK$hJ{���g+e�I��k[�w���u<X�}�y_I���3;)�C��Ri�X�P��j'!f�`[3uR2D������܋uh��@�)T=~{�0Ƹ��/)����e�'�-���o�=��O
'��l�%H�-xhP��u`Hq����k��&ߢ=!O�&��*������!b$�����w���}�s�}�r"<�Z;���E�m�r�r8�ͷ�w��.��OE����v���� ^�~g]��+1�8���U)�w�}�kKv�u�p��5a�����_���C��Z�]��9T�?���j������Е�2�x�1�9/���c�����ʼ5��U+�^X����x�o�-��K���L����n�ؠ���:�p�Y�W�\B��	��7-�_��������{�N3���܅��GP�xgn�>з,�M-��4)nKBu*K<ж���A�W�����ݡ]��L��I䭶I��l,��VT����UF�=��A�qݭ�{+f��y�`>�ٲ�݈�:��4X�x��1Ay�]8sΣs&9z�ce$�>�J���w���A��m�ֺ�{ �:��/�s���~:�ތ=Ŝeu۵힮C�W�6?'ׁ|�Czw���t���^��C9a���(�ʁ:c����J�I��L9��p�q{��V'T:w���7m|%V+n��&y�Bl�rدO�����v ��}����C9{��5g��g��J|�b
���0]�z"���6�zI�JV�g]G�6�M�}�ʠ���/�gjr����LN�k�T���!��o�
>�o�o7qgu鲧/�݀�h&�8�͸E���ӓ>ú��Ϻ�*�;A�s����ާ�M��i��_f�K��𻣦�Iq,!���,G~��]M���P�T<��k<��ίn?n˂�%�j�Q}R�F5Q�X��^�S���H�6��Y� N
�����u�}�ɰ6�=���z�d{�F��]h�����P����R��a\ֱ����^]{��\�{����>�S����Ug.�ՔK��D�ݖ4d�>�}ti,�{�W1����
1iA��+���j���-ݧ:�=CdTe��޽i�3R��4�9�T�2���F[�~{�/on�VF�<MMV�ʖ�g��5o�wM�Г���Pb�Jf*oS����:��<6�`땓$P�͚��n�)��^�E�>k>�m��{g�'�a�e�Ŧp��e唓*�5�Dyh�i��un���y&Sj�mw������
NlN�u�w�c��C��<tj�ZP�.�P�:�!�T0��Y`�C��̪�M�q6�`�ۊ�]��=p��*�
�׏����Ju;�}�SޞF��Ns�������b���q���NU��Z�~��ë=�}��F�z�T���S����f��>}��N���p�Ȑ�ya�4��fR���m��Օ>�r�x�]��{ק�͙k{���f�<���Mh����:?
��k�u�3��c�xG��z8C�jtʋ��p��0��a�4���U���x2)1�w�?�u���M͸�G!V[o�R�/�q*۽ܣ�F�hYfǪ�,I� uDm��}�/���j42s�k��0X�h��쮩��x�|�U�Գ�SpMg�	UiW	j�/��չz��Oo^Y��k�	�)mI
慾�q�=�=Y͉�k���}�@M_X>���}�� ۿ����ߩ�^�/��22-걙�
b^��U�2�4o�Q�)E�
������l�7�Kw���.QYGm�If�6Y��=����{½)V�.%o��n<�#���}�����8�nu��E��3]9��٧%�[1]���z��dl�]xM[iwRC+kq'�K�>Y���鋮Wc,�m���rI�%������?gy��/*�D�\�&!��ޠ�@����>{]�5�bN2"��KC�[�{�o�q$tPv�bg���˶��R2/�qm$Ak���']C��[���{��*�,b�bpY	��e�0�E����ij���72�Z�:�q��,���Mk���i����")ٻ�^���웑C�_*��ߏ+���^�Rm��.��V��������C�>������b����>ߗ�ԛ~�.�Ρ����Z������޷�P8<=��r�u쵄��b0p�/c�a��5�Y�\�e����t��W;f����W&�3 {��q�O�����u=�}J�چ��'.uҺ���1��L��peXfA���cϊ��E�"Gsף��X�=��:�����=-R�T%�ᷳ5͚b���@Vm��ƫ9�\S[�w��;ou3�$���s�dob������z�z�T�[�5]��j�>ʵ�Lu??���a
�� 3{���r�Z��잒�p[B\	�ݭ\"Ի;#���t1=���� ��>��E��8�ެ� J�,Xq��*��r{a�[�6�]%<!�zI����5��]M�6�y��K�9,nQΧR�C٤Nqd��EֿUeK$f-9�u62Q9=����Г�؃c�*�]*�!�.���$,��+f�M�C�k��5���!��Cz�9xgQ"XTa�}{�f�X�}����������wv�ic�Qo�����v�|e �����κQ#x��xo��G�MV��Q5�n-BGt�"�/n��w��a�;���϶��2\���&��`P��W7�BBz��\�;7EK���������Ꜹ����}��D���y:&f��9�	��X����Kך�+����0�C�(]����r!C.5�D��c�\Gx�C�7{%;��,�5�7�����D��8�5�G��peB��H�4��v�R��&��PT�]�����/rRI�|�_E[�Eo�;��:
F�_��5�
u�X�ҟ8�:���K���&p�pQ�|�X��X^�y�L4ϵ����W
��5�0�q����Yo$O-��*��C	.w���x�����3^����%��f<�c�M�������/9=3���Ʊ�9P_+y���vG��X��Ղ�yǆ���ݮ^>����9A�*1m����^�xk���J��ZGz�dv�qV�P�ӥ�XS�9�,%�y�Vv��:�B��0g=g�{�q$&��C+V.�����e��k���Λ��$2ܳMCkU�TK���_��%� ����>��� +|���я°A���R}�%�^����IӍ߷�+*:��jf\�c@�p�� ��Ogܶ��>��o�=<ي��������l���Շ�ش��B[~�s��́f��� �ES���_^�Ćmn�~�}�P����!��z�a��e���
��&�77�}��p�	}�\���z]ӭ�r���k#��>��md�XrR���y�0p����s*|�B�ͳ��$��	̉��:�����o~�塆��퉋G[ڥ���E/C����u:��n;��:����k�q��:��'c�X�/�X�N�x�Hr��"�X�u]�~5�eMލ��;G���s�"��6j������(6:s[C<'X\��m�q{�yp�_�p��t�Z�w_^k��H��Q�|������?q�;�Z���$
�y��0�j�.����6|�7��m��Bޑ�n�f�t8�_t�Kڄ;���q��M5�n|| ��W��S͆>�����Q](h�`�h���D�{2�C��X��hi��%�6qo��hk)���N�2V���,�7�y��j��lê��^�Gu����#E"�/e�N�+>o�h� �vs`Zgi���U��,��)`�+x�B�F,d��gv����|���q�u��ؽ��(�sGgR���M#zl�~/+��5��^="b��3��V8D[m���r��4Js�3gH��X�M>ķ`ƻ�郻z��-�ej�*;�iV�����B���/.��SĪGL��m�sw�7���uz1?Ed���)vM�(1�1vc��Ԉ�d�Sӻ\x��Y}Q��k2W!��;9=�t�4�O�Y�T�����\��cGA}U�1����3�}7R�esu���`���f�0��)Y�ȋ�re���N�������P\o��D��ȫ�ؙb��p+��e�V�f��tH�������7Q��Tu���g�Bƫ!��&̕�q�ôp?ͭL�fVҡ�۲�a�	�ϑJ=6�	��F��e�[�i;s�*S��V]��x�4�I[������Nd�#`��h�|�c�Q�X%�m�F�h�L7;
-n=VZd��-V�no<(��FN��	�)$�l��vte�fK�t��J�;ss���[R���Mϲ��zWn���K����q�g��lrQ�km�o�ԊN<s��j=Y�zm";����j�����Sd F-2kh�8s�v@��uڣ�ފ��t˖'A�]Z�a�=}֩;�{0R?"o۹}R�F�Vf�����|ޖ[J�i�%5HvE�`�s.-�4&5�D���iI]<l�ֳ%�C{�Y�J��w6�D���k9�;
'>A�����(JU2�� g�h��ε,��IE��X��ӻ�&�����|m�=L:�4��!=�a���G�����RцI:�g:��n�7�o�V���z��c���b��ԋ�H�3uT�����]����{[��i���<cz�sE[;CS�W���m�VJ±�G�`�Y2}���m��<0Nle��̰��=vH�xrkw���Sg`�`Ֆ�*�SR��z��^J8�ű �A���}��YA�r����ݘ���)��b���brpl�mۓy#�Gp�k��c\ci9�7AM�cyU� �yk$�rW�P#��t��R�0���`v�UJ�U����Qx��|���W<�6�Q�j�$��*�	99��n_Å���B�g���e
�j�y��h9�8���G5�6ҀdaX=���$7M#W	2�,�H��F�띘7���;XB��ݣ�%\ʸ_V�����U�Y��ù�l���o'���{�5��X*�+��ʮ���gc��*��7]�+�2���3a�9���vI�D��bn��M�md�k���e!w�`A�6��J7�4�Z�N�[P�/�Ӳ�:d��2�J0,�Lа����˘���y���Rom�C�0E�F�UV�f�8Q����2nԞY��p߅]߼ٹxUe���ȴ"AH����}�s�_�UNG"�\�*���Er����D�*�N��w(�rr9�9�"'%�NU�j�.y���q�Ã����v9�;���q�Ep��s����QQWe\��"��A\�ʧ
Vi�PQ�����9����1a�w���ҋ:Q��˲)�1=�s�ܴ����S��N�T�Q��	P�"�""���q8�T���D�r������	Tx�w]K*8U�'y\��q��UD�I�r���	�¼y��E�2��H�9Ǖ�+�u����]7Ȫ��w��9S��x8Y��Q:�Q+I�UA;iUw���7)�k�;D���*�/)qMIʹT�Äz�(x�L�	DG(��W"#�� p� �S�K�7Q8R��U9}�����{�1g��Դqb]����ά	.y���MI�N����;f���=s1]Jpg|c|�Qr+��zq]�O��]u��{Ns�6���aT��sdM���M�?w���d?'��z�HI��]�����N!�>F���O�|�|�zL>X�C׻һ�iēמ���o[�d��;65RƖx�1&\�$s������T����Н������N��_�z�?=}�x���:�o*�p/��u���Ǯ	����ӏ�'HN��>!���E;y��������Vݙٽ�X�8���>!�a���P]��7�������q�M�����ĝ��+����Bq�y���lBw���ސ���|p_y̻q�o��n%p.9Н�t{������]�Jy�#UgV��/����x���o��8�	�S{x����o����Uǯ#�u7�N^y뾾@~N!��?�so���:w����i;|��n���M;��rBM>'�?��uF?�n�����-�)�d���Yy������q�v�Wē���p>��7��}C����n!�i���GS�q��8z�m���L/��{�����;���6��d?'��ϝHN����~S�C�v�;C��[����f�Ś7�}�����}T>8��~Ǥ=&�㺮��@��w��?&���n"��H|M~�>���ߐ��ގp�\pq^���ޜO��aw���۩&��S˦�����o�i07gz��gg][���XAm�o3�3�_l�ݚ������C���w���>���{OI�S'���>'�8�_g�:���m����x�M�	8�]���N?8���>�G߄G�W�?��@D�ةaju�;�B-}��]����݆��� ��/��ݸw��P� �����P㏯|O;�����|x��c�}OI�]����!&� ���q�P�}� x���<����>����mQ5ڷN�Nއflv�t����w�ɤ����ޓ~Bz�;s���n |I<���۬�ӏ����N;}x�߹M�'���q�ߜ��<M?���Ǵ���{>A��ޟ��=�������=tb���,�������������3C��|���O�{@�v����n���n?<��i�P�q'���t?���^�wW}M;z�s�zC���}v�����'P���I��x��i`�z!���M� x�������\Ee2�p�Ru��'��v�/gt�
�$�vD���	�WB'0P��R��[J����r��Wl��[zw1���tE���E����g�6Fx#�9]������3S�N��pp$�ϩi�7N��ü��'Z�2�������I���0�� e�#࿾ǎ�I7׊��a8���ޞ'����������}M�8�{�0.���q�����0�~���C��������Ă����G������N��<��<}s�Ӟ�����>&���cӷ�?�u6��V8������c�>��`8�w��O�M�cߜ��;;��9���_ަ�����n�1uEu��G6��߿޿�����8�_��si:��$?Q�ӷ��x�N���v��[��7<I<>X뺇���wP�o�������~A�7=%����3�;N���v�ny<;z6�2��=;݂� Z��zB|v�����G�#�O��m��������_��o=p:�D�ω�;)����s��x��	$={��뿝����>ޓ�aq������>�S���;�~V;��6Y���.�	޷��]�4����i:�����\|����C�5��zM�	��?�wo]�8����N�x���#���I7���q0��ӑ�x�L,㧨:�7;C�����J43muUhz�|<o���︇�q?}��~OI�_����h~O�q���n?�$>&��ށ'S|BO_�{���<I�ӟ�u8�&�?��\q��像��Sq�x�~�]��?��ݎ������������M5��m����)�![~w,C���������C�����7��N8=�~�P?�M�~�ǎ��x�~����ԝ���n���n x�������.̝�­���u�X�k66����������I�?z���M��_xuo����r���;|x�el��	���}OO��ɽ�|���ߑ���\��۟����C�Ѹ������#���w�fk�<�_FG@=�{
�t��o�'�8�$���se뾻�'�~�̧����z���q��}s�>����i޷�'P��~���X��!�\��bM�	�p����ノ�y1�ާ�7:yv��nJXJۅƵ����G��#�?|�D}��s�$|	lL���u=�w?�u�N8��ݽ������{��8�L)����u��8���Ă�wP��= x�o�B�?}D�#�;���WU����ji�L����/�~Ә��}z�㑡����N̬�$����ӆ%��=Z@w�{�͢LQ��~I���9z� ߋq�K�{�AJ���D�N�O8ɢ7�[�s���9Z��x3CE��)��ŀWsS+�����@*�����������w�]8���P��~s�0uӴ���p?%�o�q�z���![}O���pH~q��{������}������u8��m�v��n!3�[�JUm=�5��<�gr�mvhv�|~8���'7��u�q����:W|M}��M�I�!?���>�OH{M&�~�8���;ۏݎ�~I<v�����`S~B~�����������Eˍ�5[qY}��b���A����������z�OG�+����������7�#�P���������?>��x���ϝ7��aT=o?|�='P��>��V8�i���Q�8G�ƨOˤ'�˼׮��;� BHzO�A�)����^�������?;r���z������I�O�<���@�s���u0���P�����~���=�u{�C�|N&�&n���~K3�ɋw��B�#�*��
�7���w��||x�@��oI�8�}�q�Oߐ~q�} N���!���叨u&�������{|pN��׿9����[}w�?~ẛ����]����Sk�gz�]W�8���}3fO������M���L)����'�㏿�sWo�&�}�۩����C���<Iޏq�w��n8��ߓ�ӥw�z�M�$�!?=��������;q�R�tר�랶�4��0v�g6?��n�~��z@��;{<�������?|��OO�����7Y۾G]�Zw�k�ۏ��ޓ
�=!����>r2��@�{��?3���~��ֹK7v������;o��]�������?�q<C�M�q�C�W}C�������@�|�_m�~����,
OJ�S{�?t=;�׫�g��<M:q���>�8��I�P>�0���]ӎd���nv��[����]�����	�x�O^�s~w��0���Q㺇�|N {��ΜTߝ!���s����:�Ă�����[{@��o���S��>�����NҾ�'������sZ=)�N'�fb�lajݲz��]��~ݏ�����&���
��ǎ8���M���:~ _�y��������i���w�*�P�~g���>V_�f�J�)}��-��4�}�����3�ns���Zu��־�n�^�"�Eemۦi2�������{��~^HGPԲ����m��W"0��}H{7r��=�i�d���Ł8����2�%��ҡ����ъ��mo%��{�<;Oj�L�!8}��$!;㰎5���u���xJ���^8�����n�^�T{���������=����BqX�̙w�������J43�C��uC)���c8<}�ރ�7��g���S������ˤ��S�r�(�#�eu�J�k� W��W��\��]�%h��y7'�ZW�K�D��L��/Y<&u�6:��2`U����������{+$`�ޥf��׃��dZ�"�7<���d�X9��0�G�u�O°@���W'������g��u��u)O�q��"ps����E�3��e4�Tμב�6��f��֏Z���`����<N]˲8)\g�C1;�a�^�iU`e�[�����9E�����뼲n���=����^,5��P]f|��[���,+V2W��N�"l�}���/U�cߏ������_S�w�S��Y�l�U��捞����j�yk9C��^ V��ݺ1���;/��b�B��w�4S�}oB�����×^oHp������׳�?OynJ
���tz��+���퍵J�B�����Ϙ�KNW�zN�\��^X�K���أS��,�2��P���i<,��[�Ե[���Ԇs�Eh�ʂ�Y�gt���X�zyp&2�<Us���ɷ������
J|�1�\�4�F��A�茅��3*�(��_$�;��#"���om�]��M�ϛ�8�>y��d���B�Q�ؽqzh1��e�r�2PP�o��7�t3�u���v�7=�GT�4Z/S�]���n
$�<���Oʠ�xl����9a�'�]�I/�ګeד�/p����K=��>��m�`3\ �=[����O��w�};za��*�!;��"{˺o+���
U�`�U��D��β ==�2@����nR����V�ej��+���2�g�޲t��Xnu�xL;J!cb��;�t�����}�awԡ��=h��������*{�����uX��E���lJ#],��B�;�@�~�"u�b�Fl2K,���QY�tjp����fճ�1�^�b-��%�i���uuB�,�5e���2�b��g�+�3*��j�),�__��zwP�6&�*�?��b��!r�Z�w���EZ���(�k:O�U�%Rn��[�u�R��8xޮ9n�(CG�9�yH�4su_�?�U�e�-*y�m�ͽx��Hy����g�U������iWJ�K̾���U5��j_c���y�hΣԩ4d����y �SLǇ�s��e�I�],���u����f�o/3�浺S��V(p�o���\��оޣ>�����z�#�=�/���-Qv�ec0�8��.�={��KM�Ka����CB���=�	�]z�a/�~�x��Μ8������V,w��o��Wnb2��[��R{9�Ww��:Ȓ�B|��=�Tnu#��
Z��P���Y֊�jR�p���q��v!U0��=B�����ӏ���6R+{Q�c�±����E�ly��-���>co��,���-��c�-��~v�>VG�h���{{n��h�Q.̘�n���� �V}�݃�T߆:�T�<�E�^�������Hz�{	�R�ZN�uk&�� R˽P�A`c[)-�C���W�<�pMg�	iWQ.�S��8zoX���muvj��إUJ�hw�*���-,R��wY�^]6R�P?.���z��@��F�;k�V��:c�(%o�A�^�zڞ޷{U����|�\�UҼ�bK�2 }j)7ӆ�Z�x0����;�x���8z���[ĩ$_��v�+�-�]/lKC��h��(�4ѨiF6��]�ݽ:��fT�����75��r�Zz[۽{�i�eHF֊�l�6�bA�=�����(#,�/�����X� ����nٱ����u�湉i[��Xk�K�?(�Y�P�qD2�nM1i�"A��Z/�Л£�t��5�uQp3���T���!���w�K���@d��1�@g{k�փ��/�t��z�� ��CӰ:��{��e�E�:���u�%q|LO�0D�A�h�\�r�3�j�ʫ�X�0�
�UǗ�$z(v��Dب+����߫�
6��\wp�9hqk�6�#R>�Yxo#� yG%w�Y�g�_¾����N���:�[�~~6�՞������ʊ�C'���n��o����
a���m�lg��6@[������tT�/1�JO}��g1��F�Z��q�3�ۋ����ػ����-%�đλ��"ۯ/}8P�=��1"8�����S�}v+O���^�9��n�﯆b��Ro�y>�h;�jR�#�U�X��[��u�j��3ܕ���W�� a��?��V����Ȏu0�'��:w��/jyӼ*��E�G1tי�61���(���"&�ʸE���i��@_b#�5�����1��yc��S�d�\����{'�ﱮ5'l���Mt7CY��W�/�
�$p��o��/'�<7ۦ���A#
diH�=�R��F���t��E�c�͛2�G�$�司��Nx<\�J��z��O��/:�n
Ȳ���J�%����K�v}�B�T	�T�B�Cw��_kK\פ��={��8w0��&m���3Ef�p�ѐ�1���k\p�͋�������/��sTθ�ܯG�'��
��O|�q	�j@���%�A�;p��{��O��7U�*�m�J}z�{X�Ll�RM�Lu�Z�|J�^�R{��<��{ku|OE�X�ʘ��8�^�N�"é���y�"}�u�魑�`��y�'tï`�~d�*��ɴ4��b��θ��JI�����oeqB�VM�W�&+{�k�i�
qbtHđ��-�-ez��VO���Z5��d�1J/h�.}��*���wb,��@lN�~!F�mR��7lӢpzD���MX�
�i��v{��-����z���p��π�^��A��U?yr�D{��*}�-jC�`�O��<j�I�e-���d�Ga��~�V������;�Md��]��\*�����KE���3���yL���wyK�F�Y�Cƀa���YY�
��ޏ�SixU�����kޠ���3ϗ����_�aY���Q�P��_{�[�-j}U��-�K�;��"�~�����0�l�g>�I�+h�‰w2)��J
v���.WLW{"�n.�o�jW=��
�����C���+ut[r��w�9s�����s_V�X�i:�嫫U��ozh�9�ٽ4Pŵir���;T�Ӛ��m%�Sy����� ��|���y�zq�_��ѐر��V<)��X
u�8�=u�|��_�ybME���Ȼ5@��O��^;�/"0���D3�(Cg�B��c%q
��479Gw�5]�:�I�36)wX�<6X#o������bW��7U捜�K�:�Aߺߗ������M߃Yԟl�ڡ$q�mb>���z�;<��5�|�N�X,���V�|��g(���@)�f_.o/љ`B�l�wOGT��d���c{���=��ގk���h��f���R���3���^5������.'�����^�u�5��l��ߺx�xxD5
�eq���{L�X=<e% _5�!�]���ҭ���=�ǉ帠�\��*��z����y�H�����:�/})�1��h�	6��/*�a��'�ۛ�~�Y�����虘���w��ËL���e}ܽ�^����}���B��,���I�^�����S�n�$յ�:�2��I�u�=?���a�I��bͯTL�m��C�5(㥪�sY�2d^պ3G����`�m��r�n��R����W�2���n�'���T���d6�_`��m�,�z8`؃�� CDNq��7�{���7��=���旹�B�ޮF�i�1�gr�냆�z��c-�����:��y�^�e��ml��_P��tmUX7E�l�<mn�+�d��3�6د"ȿ�=tn.�֌G�/�B�R�S�;ǲ�c�i���S͋��c�+��V%�l�Ld��1��l�%�k�eC�[t��d�;�jfxv=���3�Xj�	y�#�2��/�˱f�T�a٦6L�P�,f:������U8��/�y �S#���h���\�V9�ለp��\r�ZP��W���f�=���&�èy/�;�x`>����j���՘��;�������}�u#P��UM��}t�fd�0�҈vO' ߟ�5�t@�c����~ұ_��l�)�<�U΂m�͙4�N�BO+���c�ިV�{2��H��	b��xس�Y�DUk}��>�<o�wg]���h�T1�'@���Z�N���{�[Q��.�`ⶂ*1Zx��k޸w�� ��#�8��J��U@6Q�/ඇ�ٳ���o)�>�U��~٣����LsI��xG�����}��|v�P��UdX�5'Ψ�����~��9�U1Nem��ji�]2�C��+6o�i�A�G]�$}�L��*��"Z�B�s|mӝTj�gv��)������6����H���l'��ɀuCv~{j��4���j�&�5}�J�;r�̦���v,��Me�{/S��3T�0Q��L�3b	�^�RЖC����h �ެm����m�ZQۦ-�u�u�g>s�BQ%Tk0=N����h�|̷�/ �x����cN\��I�R��Hh�6ҹ׃y�J���U��V��N��l!kj�;��ND��nd�{�ZD7p	��8��1ޥ3f��1���/��MQՑ��aM�o��V��j����eu����pS�P�Qj#C�K��	�F
S��*�}�O_VF�D��6�l���N"�r^�̃i�4D�j��gn�4��h�BE�+g���*��8�P"��5���V\��3\�A�L������nj���7��Wu4�L�q�b����e^�����|\��V�Óm4�]�^Yc�:@�H�s�Z#��%X���ǥ�n��Aʎ��B�օ���_upL����wTԂ��6�
{m���20}U�47�����H�c�Y8*�y�!d����]\��M#l�Y��@�^	�v�4Z�7,t3�V��K�P)ف^ړV��C/��RZ�9�Y�먦�qᱹE�hZ�+g	���1^T{��g��]&V�O��ch�#��ȸ�q=�F�=z"����)�Im]���}o�Y4	�ȚɈ�{C��O4�"���m*�[#n��:1�k��m	�Eogf$�Q}��Zx��ٰt�qb�'V��
y�f�^/����c�m�)�`HlG�:,��vb9���Q�]�ZO�z۳�Q��嶓�����ŭ����]8��r�*�>]�����z�����r����3=��5&G��N,��#>��W�0K�<PF��&*�s��a�,^d��
9*=p�"<.��ղ�ݾKw&gH��݁�D]�|���Ě�-�ٮ��t7�Hnh�J��|�
��i򶆬7.���Grg�qe����+���Eݷ�ov��|�
P�ɩz�p�\���fmk�����d�ƹ� Ud-F�Tj�I�̱[����!e��O�G̖���� �/�Մ�q��{�Ȑ����u�(Fa�|�M��xN�*MpĪ�S���U�W�f�;s7#C�IɌ.��F[��E���%o@��z!�Qݷ��q����KV��q��], 5\�K�c�.i{z�N��M@���X�w������\[��d�
�y9��V��T2����=�:�X�ǥ<��ea[����f��{J��d�m>|e+�Li�C0b���YK���h��r�G`�=��
�nĥ�v��?�mLܠK,�R�/%F�ܠ�+SX��=]D�r�b��K.���D�LD���o����/ޫ�4_�~�}9�>;�Q�YyXS""�r�*]e�\Lp�P�\e�	E��* �Bn��ǃ��/^�G�uШ�v�]�\�T��;nR�EqRJ�P��.X�;XT��NV^�˯U����2�A���D{93�Z�^p��h^����"��ByZI��<x��(�d]-�:Ȉ�(<m�npS�^�';qq	2�t��G/QI^D5i$��C���J�q�Z�"�.T�nz�9��-KE)UM)ԅE��U6��9�YS�]c��"�%�G*��K�<d�QD�9Åg�Ed҈����DR.rʹ�iݴN'�N,S
�J7S��s�0�P]��&�#�s�<�ˇ-1���w��9\+JHw�xL��*��VH.����X��2��P  ~tZ!6�� �]� T�|p�]�E���k�]59�b/�v�U��[�C*�?�2l�p;���y��fWLyb���_-�����o����`̸�B���o���!�[N��9��\<3���xq�7X����\��;�Y�#�܅yK�,��'C|u���.�����ԔM�qJ�+�gw�:�x!ݣ=�O��K�<7���ް�Ҹ�v�:evX�iҊ0#�:�%�q��?Nȥ'��$o�������y�+7�DMnO��*��"#���]�(����r�{w��w�_`��B"�M!J���ԡ^��+����OZ���2!��Z���Z��~�,r�����u�3�+�B�CG_���^%Q�j|+��܈"6x��6/f��0�ܻ�G!�^T�Ss�u^�w��u0D��R����P�W6��]�pZG��������������`�Ymc��]fJύ&mw�՜O�՜��"��k�z��|�#�M��*fTo�Fp���o���ܸ�6'Q=Ӫ��8Iwp��x%�@i7��U1Nh���-SΏ}��}��QV�x��𙭟����~�i3�_�ԫ�����;�H���4�c7|M�,^~��>����L/u���^t�*�Wܪ#A�F��9x�Og���:�P����..�U�W2
�<4���+iu]��%k�F�Y6��\���jp��CBo�^^��p=<�_Ti�᪶�kR�����U����ԏ��o���S������ō��0kC�%S+�3X�� �-fg��,�� �Y�ޗD̜���q�ȓ�S�wj�8��_o�+̾C<�V�N���_��NhogC\n #�t���/"��3�"�MpwQ;</Ɛ���"=y�Вj�:-<���=���Mqo���޽/v��(������<C��������3��.�[��Jخ9M����m۵�s��_?{k���j�}���g��u�k�A�eRQ��uݶr��;k�3������M��Z_,/�������9�������=Ι�DԹV�r��]Xq��~���m�s���D� ݁e�V�|���r�:k�=��֎>>�#���5Z�~Kg����<1Pz�[��B�˟�qV�r�.�={ӳ�	�������9e?
�j�Z��ot3�{:�;������SX���[����[�o�ʼ$��_���(sL�	��x��ze_��R�/M�+Q&��ڠ>ȩ0�>*5�WE�)��H��4�C<
����fS�tVDH�����)ўlh��5؈���n���}��[�2B
^�ѳj��:J�h��J̤3]����n�	�ú�k�>����nKۺ{�Y&ʵ�cO�0�ֺ[Zк��!YDl�JqC0����L�T��7���Y�Wr�4.Ŀz�Jv�1����&_d�DyJ:Q�^YH�u^(e�j�k3o�����5�<[>=:��ﮆ�Cx�7��~�,�!0%$���&���Y)}�꿸� �Y�9*�si�6���ɃP��5Y���۷����7��0�����9�Sd��|�3�|�to�^ڴV|��1��"%�ȏ^�Jh3T�:��0���]��o��|`ה�_����40�RجxS�<�����+�=�^Y�`x̄�i84��nֵ��5{��c��Z�S}A@Ɗ�f�p�����e�_/
8x�bۍO�������ZL�R���b~N3�pQ�>;������W�<�mQ
�i��9��}R:圕��VEM�k$��K�M)�`1�g�>��[���	~��������u���hoX�oo��ϣ��ݓ��<�j��|�
<r�_g$4�;Z�2�HǛW1���r�k�{R�>ʝ�6h�\�r9�o _N�^�p��T4��{k��	�����9X�-S,Z��&P�Pm{����wÊ��B��8�p(��83��}�Ӄw|1!r�p��\��U�CG�=�|��J�ڣ�c����������:���y\�b��l��5ӄ��W���gf�$,��]�̬ﯻ!}Bb�6�M�N3��a��RI�����f�m��I1��,��s�y��F% _5�C������������ǌ][��V����3�����[ي#���<~���FX�/���&mW�]I�n�J�P��a��ܮ"���ґv_>�wMo���5���J�=��k��<H�(�β�a���L�*�k��liqy0�i�'X��<g»�E��g��ؑ�}n������uT5Yڥ2�����\�om����L�$����������t�lw/��)���Y���хH��ɟR������Ykz��8��u)���]>Y�s[���:�%m�`�Y��{������Ko}�"5�qA~gy�{t@�դ�jg½p��Hх���Wj�*�xcdʥj#�DZ`⦜�;���t;զ�蹞'[U�"n�����:����!�j�RP񁙻tx�Z�=~���a�7'x�9/�[�.w�\���3Xw�B"������]�Y���� �a�ַH��iڷyr��_�t�<b��q4L�F�hR���ﵗ�����zC�p ���u��(F�
;��ASt�� gUr����Ʉm�\7��ex߃�4~�����:|��Ϲly��6��=���MQ�A��WU6�-V��8��M��;aHi��.�8���w�Ň�2�����y��朋�J��Dc�F��U~ 0�|Wsu�'���t�>�Hw,8tOR�,uR/+vq�����컛٩{-���ҽ-y�Xj����w��uDzσ���^�(k��d�}�{P�-�.b��3�>>�����'g��~�5O�حc�*/�\=�G�����U�	���T1���Mp�i�yYN����f%�hʮj4���;�_Z/1�+�yv_��i��al=�z�M5r�����U��ƧR��k<xA�B%�x���//$c���~RG���y:�cU�5
�ه�(o�y��UsU]�}(��_meM��&�1�.w��������u.�w��=q�C>��|�]E1"d���1Z]�l�_'�F^?YqpU�^�ݝ��w+���N����ayr���b���O���y�{mn{M�,��#HU'\��V��j��Zy��i�ہ�q�:�hfjD����.�Nk���P��
�7.�*��8|��xS���S�Cj$��/�!��*�*�o�¹��&�ާVT�
��Oϋ��XJ+��ŵiŤ�ˤ7�.�u����{\g�&�z��D�VzQ��7�t��D�j��P%�aj�\��P�07LÓaa�[>�~ýn�WՍ$�����_Y�0��,����3y��+$%�%�v(fS�wMm?2[K��ם?�MG���_/˪����.�p�?-��+��q��X{���K�Q��w���`�G���rWf+'��h���l��R~T��,�y��k�ew��ᱶj��nu�ϊB�hB�R�^�EA�/=�F�<Tp歅t�֫}Jo�;�t�xJ�wE�"�b��[�(��E�P������Dm���b�Z���r'u���X�W��,z�36���&�ד���v����ah�ݷc�
@E��E��R�4�MA��E�^�ׅs�ó*��Zx:J�����BxS��=���6�3���Z����B�i=T�h?ۂ�lU�(��������Dz�{����~��u��ѻ����)���f\_o�.?\��y��[*���Ƴ��J�b[�Gϐ��U�wI6����ϵ�v�e9�}������Zm�*S��e�3�����'<�F�����c)�����4�{_V�ҥ>�z�iϤwD?gZ7������,\���}��Q�nٛ�Ժ��E
e%��RoGȳ:���
 �7Ⱥ&�J��c�],�a��KFnK�Y�[J��Yc���(� ���cC�m �|�98P��Ҏҩ�q�Ԙ|�f԰]E5�����^G��K�1S&��P �~���������S�n�_�XM���r�B2ul��qMY��C�k�¹��0�w��v�B8��~�K�S�Q~�l�@鍡�s�!��1�aq�����t2�W�^�-�w{;�=<�VJo��wX��Y� OC��%g\/>����V�y�g�`-��Q�ߓ�|=���p��U��r�2Uz�%������ԟ0�S"����1���:���u�>Xt����g�n�l耯�Q�^�,�1V���q��)����?)����g3���q�*�J���r� :x���4��û\Kޛ�5>�`�yl1!�O��9�ޞׁߘ�
7�#}jӝD�R��^$�`�BR�{��b���(��q�'�X%Pc��Uϕ�(���j4��vt��4�*1�bN�!18J��%�	|^C& �c�u�H�M3k�a���+��N��	�v8N����/�T���g����qJ�Lb���Vjo�-��ͪ�p�	B²��xQ���~��y7�a�ƍ+ִ�ʮ2x��L�3
�c!:�p���u�F��ސZ7�c��iW��V蕾퇜Ԥ��N�_f��l���4�J썡��;ڏ��F�*I]�ݮg&L�-��Ͷ��)[}M,�H���tk�M���B�:���/��1�6�A9vv��d�������S,�3v���ϖ�h�O�З�	~�#�r����W�<�m��i�[�uf:�������s����.� +�9�W�/D�2-�[4|v����zw �lLcu	�G�f��|~�)xn&����#��u/q��{�8o����<ݠ&u�9K�g����3d1�U�
yw��z��X���9�Ҍ�\U
J
FR��Ў�e]�\�������ؠ�T4�ͤ��j'/.�U�mkG=\�8�g���X;S�V��T=���1˽N7ɟ-ձn�5�/��!��_�����m�	��z�ǝ��^�?2��)�0��,��P�ߩ�x�~�@���-��L���5�f��B ��ɘ{y�d�n�}j*.}&;X3n2�׹[-�G�i�Si�ơgݴ��qQ����0�(��@9�.�l�[����y{��VUx��	��'�]`�'a���w�`p�F��qCQ��_m��|߫,F,<�PӦ��-�����K�:�},c%�׌E��(�wۘt�4���D��c���L�k&ԻY�a�tH\�mG�{Ef��}l|��z:�$�1>���g6�k�ѻ���Ï^�*�[ޖ���9t��.��������j�6�����������L���D�E�;w�*��fo7�9v���˪t@~��t@ �2���v��g��a`���-���|tҹ��n��W3e4A��(��g�Q���xd�T��wA��]��c��㴄8x����X�]Vg/ߴo�n����([��!=�e�l�U�^�u�D�W��HW��!�2ox�U�W��G�
�4��Vx��dDȺ���8�q�y�'�l�Ê����KS�-���7�nf]~C'�MA�k@���t�K޸SC�꣓�/�Z�h��C�s���F�^��Y#�3�,{R,��?1C9^�Y�<K<o�'��5����y�s�l��6��)2���1���:}�<#���V�yVqk+޹�(eM}�FD?��0���L&��j%�B�j���4��b����݃�߆;T�Q+�*��SQ'�CK:��˺������z��د��C��݌�|���4!��)M�SY��U�\,ܱ�(�Oz;6q#���S1Un���a=�ͅ���B}�9�g�&!��u���.���_x�a(Ѱ� �k�}�����+~Ci�[�����v���=��Q��嵯!��ʻ����Ew>΂(8��؎��Ҡ�٠�5].���t��-b����r�j.��N���;[��"X�f�םNcz����>�����ǌ�bf8^��OO��{�����Q��a�w ���[w�;�B�4ɦ���OQg�;lq�[J)�:���U��+i�Ȼ��U��(���q����5�~�T}����{˞*�'.<IRH�[�H����th��c%�kBe��{WY�x{w�R./�|�*Q��5(W�״���U�c��'PdC�Q������;����7�G�d��ˎ����
fL�Ĩ\���\��O�p��q����NR�+�=��vn"�����RP�UԴY��!ީ��<�6ǼUMʼ��K�1NxϮ�<}3}���߻ؠ{��
���gP���ZU���<����Q���\69W�(:=_}���õ�U��
�x�;nz7z���m�><V�D�6��7����aY��w/���×u��՚�qN��l��R~v�=�r����-W-g�E��)V�Ո����ph/N��{:�B2�`�}Aq>}(�e��:�����,�񃷨>N�I�w�*h5��5��Bq�J	X�hF�=jحɔ�
���wS��"����e�8ٷ��e�e���n=su����>�vwi�ܫ�_���ۤ8�l�)Z1Й31�zt�@�Z�)�.�wR��y�4��ޛ�������]X�4VJj���<����p�g�]Zf���iP|��r�-kӁ��ٔ����֭��{��>(q�ť�x���.�*h���-���a�x"���V�������k�KuCڴ_CS����e�(����:���k��;O��|b:�X��ef'c�^�Ƕ"w�죓�ڻ�_J嚹ñ%4�GyX����9�ӂs	��D�j���/jK�/�7��YPB6�����������Ք*�&���É�q6N��u�(ż
��<Ю	_n��ZDv��w8;�����^��NO�-EVBS�u�����mNʛY'4�2��oS2����sR�$���K�xe=���<�}�,�I�	�.��]\85�S�D�9� ����i'qax�ä�)LƷ$����6w	�%8\]X56�x2zu�r�l7׵�,��Ұ�:T4�KVsf�kjצ�=r{|�*gv]4�9��JY&��_U�\I�v��v�V�̘��쓒�л�ڌ��m�#�p.`S���Rnb�z�����}�9$��m;��u���8d1fp�쫐_#����u��(۬ˣ g�K��~��\Gu^p���S�	g��H���< ��w�W+Si�ٽp�Vg%�[5�jn��ЭU��1���G^�Ӕ� �-�?!y[�չ6J���9�kՕ�����W7�V�Q�J�uzff�-�Rfm��:ߍ@�er��gڭw׋��%WH�)V�YX
��r�e�v�'�]]Q���m�=+A3wN�2�F]^`,fyZ+#�U�K7�:�Af���e5���7[�վ��;9`P�ڴ*g�MdR�ެ#���Z����z�� ��)��P��{v#=��8v�Q7j���ˋo��o))���V�����XP�����"���g�9T'��-�2u�K�o��788S났����=w�vaZ:�)�(��[�u��AR����ee˭���i�����-��fc�4���r�Ts`��M{2g����S�J�#p՛�̇�!!��Zc��S/�T0\
��9m�o9e���݇k�]=�ki�N�`��V�M혌��r>k���\������T��(���hH�"�7^�jlD]�Oxd[6�ԓVꁡE����yݼ>�H�4� ��b���v_f�kok����zQ�v�y�J�#�6�闱����^�tWϕu��M���đ@�4*��ex���fFH��ӝ���F�"#���:U{��s�{��!)1*�AD����*�z�^�VJ�B2�(�"�;Sv��(d����,\���C'k��Z$��5	/yƋ�5��$�[��B�Ҋ��RaBbAQ��+J;,f�\���R��J�U��)�RHOri�RQ-O]���Y��0ʣB��0��#,q%9�9t�9���B�#��q&�VF(�j�J�JBC*���9ƻ�\�.]�
�x�f�HJ�bU�-��G(��t��r�⭢�EPB,�.r*Ya*��\��:Y��ʎ'NEG"3#H�,%-9nNl�Ys@%��f"*H#B�!Z&Z);W9�YJ����8�UJ�(T����#���yK(��/h^E�[γP�U,�S����]t�X��ON������&��G������>A�7[���#�Wf�f�Ön���?{��7��Y��KUm�Y9��rǉ*���?W�ʇ8����.�۝!�k�qoӦ�r������s�O(���NF�:�%p�,�7���'-�.X��*�N,&�lՁ\�J�s>�ͱ�&�{S~�*X��^CSA���m����/6�,�uSa�>ѥe�(�aK��z�eɁ��*�۹�swe��oݵ�j���.9c�N��Kcɧ�'L�%λ5~���WY�}�Ǘ�i{�uo&&������J�GW��_H��vx��G����}��۶%N�_�!�*v�����=	��x�҃�jv��Od�ul|=!�^)��d�y�+�T�((:�k�**!��
�2��ޑw�è��r�ո�JPW�gs`�޸�Ø񝝉�w�5>i0.O/o��j�&������x�^�=��xҮ'�HF��#�Go�Sṹ���F��{#ZNG����m��Ƙ��9v3�?.}��|P�T�2����`f���鬺=�t��yv�Gb�8:[5V����iT6�K5�C���F�OE����,�3jhYަA�;-v@���tʒ��1�4	m��T�yfҠTv�N��N��������ࡥQcu��+2��D�V���^˙�Wbp�ׁ<AW�K�=�)���q���o��5��%�v�ɅP���tetyv��L5��Ҫ�G=V�=\���p�џ��ڢ������]�s�b���)K��L˕�b����RȺ�|�fP�s�f������͙�B���v��{ۍ�}{|-��)�����,U��#o�J���"�a�:qwfժ���M9�9�e�bj��-n{��\�~��X�v���[�+�"&x�R$��)�H�~�0�������mS�����k������ƍmu=j��l��_I��^�z+�^��,�<���D�%R�GZ���ӻ��@��L��7�A�J�%cլU�<�����ݞ���J6�ȷ1�C�|;�L��;�]�}�x/�AB��S��&�P�����X+�Ƹ�3V`ucD�ܶ��tX���O�(v�D�N���+n�*�bP�f'l�6��7j�,1c�8�o0��[�c{�vE°�%v�֦Y�N��|;��5��XzoF�K������#����h�O����{��X#��5�ek���E��_}U_R{�l�[��>sbY-��r�^�k*���'~�������3�K-{y��Νw���v�g0��i�}�^X�
�ķ���;�9{�఻̼R��[����������Y[9�|�1*��o̳�� [��}��Y��s���~B���6=ӭ�c7�X��d�b-!t�#������G���<�鸨�t,&9��>g�gE����0_v��i��Q3�N�]���nk�w�r�p���z��W=5��h���r��T�{��=�v���9��pyj[^w���%Vw�X�����|�����Cϟm�i�&�1�IV�=eClʟ^Ö�)�|TZ�"�Ϸ�~�_�δ�vLQ��V=��c��"�@���R�P�˻���ڼ���r�U��:�&R����mՙ閖��qq�W˩y�gVl���rUU���{�z��N�i
��:�%	��4p�+.��k�ϻ��](�j殍��R�򽐉�\��������(���u�W]���@Y7�r���%���f�����h}�����p����:�DH�nA������c[�����n��f��Vٯe�g8�H^]G�S[E>�Jܸ��7%��X��My�\%�v�����C�ױ+�����B�=;!�>@Gy�Vs���ܓi9�Խޛ]��S�<'jo�h�r�"���oBw���4O?s�Y=W�j�7�s����62j��[[�Y6�gW:�˺�4ˋ[�Y��/�hW�-֯{�Κ��j���3^|����j�!ܼv�������ǅ5�=Y��Tb��VN��֧�zM�]7�
�Պ{�^n����_�q��,L*n;%��v��j�c�u�l�-f�.�+�&�b�M��6�>n��jm7FZ�iʊp�י��Ӕ��2i�g��Z]� ��ZQ�wqi��OUN�9I�����5��ț��A˃F��"�9�o�G{Lf/N��j�,��M�+�;	�uLs�U\��*��>�2�ř�V�ǡ9��==
�5V9�헗y�;G�T��m�c�:�Ԧ	]nn)sz�`6�@��a�K�J�.۱Cw"b�ͩ����F*����K���ֈ�Mݞ��:�������
�k�+
�'���'[���ל�2\J�E^f���g;��)U}�W�R�H[����E���u���+��N3�ڿ���Jj��Dؕ���&;c|����=)M����
��u;�c�����ug{F*��
��#2%�Nd#D�"ųF���]t%��yWjj���8���턥�Ŧ��Ɍֿ"�>E��R��s ׹�6�W��54�Ϫ���ZԶ���3h�[mDbot�yyw��U��^}�����~�+l�철�Tqv�=Yܥ��_^ѭX����՚۫��=bi�*�+;�W��&�/1���ΙZ3��H�5޹��{���@�ո�Ԯ�r�*�}˛��+B��{�����3�t�>(�J�Ӕ�f�|�U�$�d�ݻ��^�-F��T��KK����
�B���4yI����=4���H�B$�_/��ޗP�^��Wn�us R�|�-������Ǎ\��Yڝ݆0���Ǻ���;]Ww.���%�<� e�7��a��9�󶸟{�2�l��64.�\Ӿ����j��\Nu�f��Tz�䳙trU��K]G�)����~����.F]�������ۡ�q���e�A>
d�:\FSc}�����Rې�ib[u׮�+�`�����-�ObX���}Kԟ?x�׌��]�{�Ub��o������lN�3ô�w�P�ܥ��t����Z���sôMc'�;|�GM�띑��+{��K	�%��T'�P�:=˫�i{h�۫��+��V�U~䫵R~�X�ڰ#�V%x;�_�e�ŏ��o-��&�{4o��b��j��L����2لSfi���%lީ-8ԴSCb��ntdo-)q�r����1`K��C]̣�U�c��IKA�3���V�����^z��FX�sy3sǏ���D�S+��^&��/��ƪm����\[Aq>}舣��1��Y=݉��;�w��m��.{g{˹�WFw|:������t9�&�'!�������{h�]��cxe}킅����;[�5�;�y;KН�Q�����4��~;b*��ebS��F�KmARrV��n!�L�{��_nq��_���kݫ<���W�f�����k!�&�t�o�����/#��mK/%����;A���˷��C����B�T5�9�Y���X�3�7�N��a��~�����*��䥋Hx�co��������g۰�5'>�J�%�U��4�y��#V�Ȍh1inb��D�O�ӈ�3Ai��K;��Pv9��$�m\z�����GY���v�y;k�,J���Zǅ�3@�3L�ea)a3p�q�T�:��&���lZ��Z�$�g�۟RL����F0�Zj4�tJ���6��&f�%��y�pʝ}�/��$�Pv�k�L�Y0;�d���W|�i��&xdw�7�9�	9G��Xꊀ�w����\d;�-��~��]j^�s�ބ�DM.�k}������wWz�_$�9YI�Ś˪�H���/bbm��S��.���P���U�Jּ|Dg�!a�b�t�K��)ꬄAdM�WX곢��w�7�{�=�ѡl��q�ɾ&k�$�e�S%�)�U(צ�[��&�]��.��>�x�����͙G��8zm+��k�͐X�ổo�-��](��8A��)r"Ɓ�Ϯw� {Z���̝���h��aVv���>Տ�ƭG��.v��/4��t61���{p�*��������S3������Uǧ%�Y�9ҙ-cj��h��o(z+�Ozw�����墟o�<玼�3�٥gvw�1т�q۝Yދ�� `C(�j�L��n��w���~�����j��kK���3i�Ⱦ�#a�SK��aK왚�1���c����z��6��j�^}EUճ��j�� =����b ���%�efЖkV2I�̦P�C�qώ.��u.�c��[�w%`9⋻���������#��8k�%�$��wxq���.���1c&�-p�,}�M�d�J�֊9	f�5�4S��Q�/8�R�y�����	+C��^�mG\{��uW��l=Y嚎�Y��6t�Y���Vq�}���0*0����vUx_���U�{������½��TS<�,����n�.(�JJ}��8���PM�� ���J�GW�.N�Ùs���%k;�*ū8:<y�~��h0n)�L���n���I� ������P:;E �������qx�g�>.znqI��`�֑x[�_uֱ�jv'OjWYX�kt⮚֋Ja�ݰ��$הrPŁ��V��;����'�s#�c�%&��ǄZd�5Vr?�~�� ��;f���w��~ �J�8d�A��/�����s����N�������|7�B�F�#n�E�g�W{�y:�G9�9���P���<Xk�x���CٓjOf➱�Dן��QyO�[jev ��v�'Y5N�a@�;���g{��:p����ʞ�gwB�xt���9��Z��w5#[�D|-O(���h��>�mz��ϗ��_(/���:S-�j����Y�u��=,�\�,��z�ŵE.Ҽ2�+��2yެ�S���|��)�CV�Z��&�����]W�z��z�;%��U��<�,�ݔ�T���2����Mk&k)�}f�O��[O�mx\*��|�|V-�Խ@��}�0������-�y�̣��/S����o�����t��9���<���fn�-8���8z��X��B��m`��a�=??16�+�}�\�Mz���H����fXe��~�5�i=ӽY�������*�A�}��/tT@���緋	�ۓB�b�K�S���>��3r��b��ͮ��%[��,�[���x�4/���k��ΈS��d�|vl{�M�}����`w�l�]�k.�f����T[�H�䬑�y;-B�����r�R�m��ś,���q�T�@�k:�)�<���/<J�5�܈�����a��UbE��#M���00��ɽ��u>ǥ[g�O}�+��5�Vzt#�Ɵ����n�l�[ë���DϷ{Z>�iS㛕i�W�1��@���F*΍�f,xzo��t�+3����W��ר�����xb^&&�
^����Xq�L�2O+η�ޞ�_7����Κ_2��U&$��&ݑ�Pm$C����"j�~��������Yp����q�����N��:��C8�e
g}����l�&ƞX�}{ܦ�q.�Ε�9�N���҈i��۞VY��s�q�uA�+x�mA&��~�؂���T��פ�|=Y9�u{�]����@�dᕃ��}}[LL-ǃWWf�
4�Z�^h�IBgf��/�=����A�M���)c]*yu��,��ME����y㪔a��龑}��U,�Ώ����4�P�����D+�!*t�."A�h�5����[����_*�"TxB�Ř���m�g<�]k.�;Cz�]CB�(B�tk����-�Ai:&>�ZV�b�۔�$�0��;�A�Gz��s�Ӡg�ΕyVK�un\遄�ݴyZy�5�P�I1HVG�r�����WU�@�%2fŬ}�ގ��\�ѝz�Ev�,���dӁ�sL����죗��;F�{�]�����%�eK�@�v6�W�X�Ji�őo���zi�Dʾ�`v�FA4D��$*Ed�{�����{WS"�;F>����z�{[Z]��g���z�G9Mз۷4��H��V8�uqb��ڥ��������+�1�5ժSCl^��kbR��ER�����`[�q�/U�$v6����a�T��Z��u3u����V��Af��"�a�Z����窍��R��������ä)'������ �ܳRjo����[	����;X2N����$�b��Z����Z�r�t�
���i&�c��{1��r����v,�~�CI�D�S2eYyLb�[�,j�&K�>�7Gs8uZ�r�4�ķ���ѿ3�O,ʭ��;�	�@�T�.b�M����/����wХ帠�LsX	-4lRqh�]�ٰ��am�����	u�;��R�5Y$҅p����
��
����"����5�3�5	 uե���ݚH�$ �t�ؑL1��ԏZmK3��-�0֎�dKbL�ڠ��R\Zu��!��x�g�\Y�eQ�	6
�����*'��аkr>�X,a#T]ۉ�[��,l|��.׎��`rfp�t����呬]5[���d���[�xҊ���:{S��+���*�G�7F����+���Z���4��s����(�A.�xY"Z(��ԳG��<B��
yK�c�.r��.�N���Q]��	GC��lvn�X�����xj�6�x{�djm�� �-���oDDyG���<�n6P7��2F�>���m���B�Pu�so.�B��*o�un4ᾍ.�m((��|�U@p��R��=�����n�r��|R\�	���St��}�N�����E�$u�h��N�\�L0�l��~�����8�\��%wg�|���X+�
�n��n�RN�Eq� �b�"�X5�5B�$�$!w*d�)�i�+*L�9�>�ӭv�����Gt���<-����u^�b��WG�k,��?n�A�e���uu��Y��؏WZa��F��xT�Ȟ��&_f�Ķl�3���N����t��e��Y���|܍��4��+κ���G1謍)�v_w eĳvfKV��Z��@e�Ϟ�ռ�h�lsO����V��gKA]�(��F	l��n��5]�ʃ��)��̣`��[cu�poGñ!}�m��pᩥ������@j���t*��JB���C��z���?��]�sZ���*��p�KG/P���E�,�Y�����®�
��0��rզ��R���L��q�%�$$��K#v��f
x�'%�"a(F�H�9ĒQ��b��6�UQ$iP�RvY�A+�.�Q�!	,�A�P�.��Ԕ�g)A%H�V����-K+"-@-2��- �)T'+��/y��咪��C��+N�sq�Qb��Q�
�&��iZ���d'(��H�&V��UW"QePr2�(���&���˜ʔ��VD�2�"�a"�D]�<jf��
-.��+5')�����f���Z�R ��ITL�#�D#���JE��'H�IT]P��f�J.gJ�%+dA� r��1JT#��]��ÃihQjEY�U�	�Ϋ�sp�2�������tq]�S��i�,o�����{�ʽ(b<%�j��LI�R��K�N`��}EY���P�u�js�����_��o��:n����$�r΅�O�p�z'�~zR⼯٧���D}��f�b����Y�t��E�X��>�`�?U��츭v�'O=ho���S}����Ydz�l[�-��н�O6y%��mײ���o�bv��6\��}C�!7��ݥԽ����Օ�}�{����d�K�T]�����G���uf�S(z�_�Y�2,j쏸���'�s�Y`�#)N�J,[3U���bmrW�~�J��B�����G�;�Ƿ�����ukK0Ҽ[�<Nn>NYk8i��icA"I�њ��ZSA3PZ^%C�"�Y%y��KUgĮ���������9,�)�b5�TW�؎B�޴�onN����u쎾���������ۻc�u������ئ��h������e�7�k	�>��OZ>�E�Þn��d�{�Ra\S�#�u0+b�fD�N�5�p[an+�5�Tͽ��E�]�����jd���cz�O=T͕�8�ٜ�Ǳ�B1�U�-U��7�%R/~����6�/�L�V8�:掙[}��x7��O���)\�t���#�Jiy��\��%
ӬnN��f���fɴg6w���_��6���x�=���R����wVm��!��2���d�}�w���5|hS���BMV|M���-�o�= �b� �{�3wW�Z�Lb�J�dub=�}��UG�y;wr]�9�U ��8<�I��y��}U8tr�w�A��tl������{�/�io�I."��t�=O�f��A|��O�z�vb�`�x�W��w�����������32.���a��elB���r�ġ��XvW�x��]�D}(����OfܔmOW�--��d��m.�T��g���Ŧ�_�������^aUVl�R[7� ���}��\v�)�صu/oϩ�r�>
缒�/�����8���d�~�ͤ��k��E!��5��j*,�P�-e�lɚP�ף����z;��w�5�B��m*�X���cv��k�.�i�
�`ڟC�.����%�=�<72�s{g<�F��j��D���S���H��6��vD#;x�
��5�%��m�7xr�KV�10/`��)3~®r��v{����m�6 �^q5��Պ@*R��qk��z�Qk���Z4RPM�|�5�[1'�eS������c�vB�e�@�{��۰��R�jZ�[J[#M��7&�"m��V9Q�3-�%_N�(���ת�s~#��#��>=�o����E[�Mg���s��Ǳ/=EF�nÂ��m`��{�*����ol�ܓ>k���k�cDe����A����w;f���,L�Kh ��Ε���ߤ�<p����7�V��/�i�GώP��{����j9��Л��iz7x��W�2S��`=GC�qK=��{ƽޝ~g#�T'�S�:<A�V}�M�!�N�a��i/y�7�D�o��o�s�?W��b����j3��	�UM<Yi�nezy�}������O
iz�s���Ws�5~���<;�	{�2Ջ��bUy?w�!���f�i+y�Ay{唦�moeۜ9Ľ�UN�՞�O<~�ٽpl�g��##ym�J����|��7{T��խJ��~����VK۟��V�6m�L1s4_bY��T�T�GWn)y���e<ݱ�x��Y��T�ۋ1�6�v��S���j��ڎ�L�6�&���j�|���c�ێ�r]��v��:(����=���ۜ6v�-i�������{�oh��q+|E��5lZOB/�bn�9ey�vKUڟU�͞qXM��|{;:�E�f��dGk� ����� ��궼.�Ҋ�;���l���J�lJƌRs[u1L'%6�۞�?45y��m���T?g�7.I撼6��*Y2׭f[�j�-,զ�Ų],8���ŷ3����>Y���n?N��[�maAo�bY������mS��WV�9r�%9�,�����pY�k�TϒQ��i1-TQ}�E4�6�4�R��gggs�M�a�e�ݦØV�3�}��F{o�i�u�c�V�W�X��NϺ��l�e[�$s���wv�}��7 �Ň��^��m���ڷ���o���;���{����̛ύ��
�a�i�Lz��ځXԂ�~>����_sZ���t�a�Z�%zg��!n�x��c�0PQ��25挃�U���7�����9uj5����Fީ1��Y;Z�]vS8O��՞���û�����^�/3iV�L�H�^(���5� �m��n���B�˿��r+������U��9�7V�4�b'^p�"�F��l�M�m����y���V��ڢ{�Q{�T�v�ʍ�2�gR�uz漽\�dL�#�q��������i08ו�dnZ1�A˺r���j1:�rMiV��nh )bGf��i�(�6�nU��O���;~�C\��_/���:]!gX���հV����p�:�(ǇϻƝx.{j��z_by0���^!�o���ދ��[�6���h� 9�z3�k���G���&E����J�/�ә�λZ�a��ى�a)��Z�|���Uu��;^ˋ$�t��oS�}�=ڏ)0y����X��y����ղyz���sW�]�a�p3~B)؏��D^OL�����g���kX������L����ø�p�n�jw���/{�k��f�:v����ͬ�^t��m1��Z��t���c�g�Տo'�6���=�r����rW�{�~�Z���m��9�QI����ۻB�vr?Aw/_G�n^:2��r��V�cy�@p4KB��\P�uү9W�՞m���؜2�.] �AE����6r�6x�2`��]c6��yd@Z{���0ft`���/v]�2�������G|��y>3{ՇI����6dB���ꯪ�mlvvW�ж3>�TؐG--�wn�V�i�Ɋ$	cU�V���n�����s�~��8�����W^X�r�Y ֚�탕�L�X�F��{Y���z�T��U+��y�{�W�G}�K��=�����ڐ��� ��j��[a����[�*�%��nzZ���#��{T����=�q:�̬��֜�fy�ޥ�+�1ԯ�Ч�^��[Lv�ʆ��,c)���Sr5��J�	�~%ɷ+ڟ�І5YF}f���>���mܪ/��<]̩e��Yz��V^/xj�,t���ߊ�j�v�r}�=����&������'竄�d��{մe���s𕃬^7��DKې��@N�=7�5����V�Ԑ��f'�@6בj�L�$^Z��S��-���S3Wt�D�t-���#,]���|��O~*=�󱔻�3Ɣ���]�n�����4Zdk��o�h��g E��|WI�Z�_Q��t��B�8�2��~��h5�~9j_���A}B��7y���,�Sat�JJ��o})S%�F��zˏf`g��]mvv̋��\�'���tw:��u�5[F%I�M�*�+��2�9&Lr���7���A��;��Y�}i�jL>ܰ�RԬՊ�+�a;)S3���dE0w&�����E)y��1X�|��}�fڎ)�صu/m>��n�6��.s?M)t}��~�p9���5c;�L;����!�8qv�B��{s���o��oWy�z�ºk���Z�S4�����+Vf�]93���Þ^
�+!z=�ze��ƙ�N@5Ad�P:��玥uh��收A���X7ge.��xc��[�巼=�{�r|�h:���jV8�U�%�*<$�y�V"r[BJZ\ҡKkK�׉^(��M�Ї� �/�������`�o�駞��7��9H<�f�xˇR�oK�_!��BKr�o�/R�[�+�`�<�b�y����a���� �y[Kù߰�b����w:�r��'����Mb&}��*آk1j&|c�Y�V=�WA�OD���1�����O"EάG9{��*�XŲ6#�uíC�2����^Ǻ�g�B}�0l&�;��(F�J̋+��l�����<�^�4���9�l%Áe�.W�JE��ț��uuI��gpN���g"������N�����x+������d8v�>6������Z��%,1��}۶ӷ�%m�q~s�2�\�(:P��b�U)�V��aj��V�Mz�6�mM�/��mMp��`s�4�$<��y��^�?t#��u��fo"��+|�)�W�ٔ�2��8wl�	�zU�󗏮o:,��J��Ms�=�/�ʳ���Sw�oc^0�Gh����UL�>&-Q'�bkY�9e얫�5qr�yÆO:���J�d��xV�2���0b�-|,ԡ�PS�L�r��党�R�H�X.]-~��;����{8ow��f����G�p����^Am{��}�Tٻ*�ߡG1U"�o���O���,��Ȣ�NrՅ�L��J�ۛZ6F��D��N�VZ^C�M�v�
�dϨZ���g��V��G.U�U'b��&*�ᬙ�����q� �o�hUk�o�N߈���|>�g"{�^y�F���S�f��Kn�7n���s($2a��Մq����q�:>��$�$���۔�<�gP�:��l?�btN�e�� �~[�+h��Z�B�eI�3��CKs��巉&x�	w�w�)F���wz��+8�gI9Y9!�����E�֓;WO\���I�'�5Q��z󷳫��+X�|��I�|xR�ʱ��q�*���f]w�g��:m�����̲�W�Tx�"6��TPV0=�5�i[�L&�2�c6�J�۽��T�Co˥��vv��aW1�J߆t�a�Ä�AxZ5L䚫;7�p�O�V9��5�}�\��y��,�mc��M�6��\M�����I|f��y�v��,J��r�/�v��^�%;o�$hp��+X�t,g�(e��I�����wk<��n�&���9Ҍ'�{q�g�S5p��، �eCKbr�E,��PӶ!���sJ�c�X��faV^�u�f�[F-���h���~��gἶ�]��<��͍�:/WC�3�\5�}�i鹎N	���⩰9�P�+��ח�:q���risپΖ���ǅw� A����G��C�'V+}��7��l�.��c�8:�ޚ73RW��cjH�hf/bn_Ex`VD=MR�2s��Y��S|��<M�Xnp,R��/�{T�;1lx=b��T+u��1U��w����l��fH��)K���u�����ࣙ��*���e��dyWP�S�&B�lї����S8�Fnm�x�`UM�j����N��Ryz����[�*�a�������/y�J�='�=/t���SO���{�+�l��S���}^�7�n]GނS\���^A�r�ϱ+�9e\mx�>�`Vb�g����D]b1MuCR������قv�&���x�bT��^�ޖ(Y"mQ��"옼�����q�56�gωU2E�J[ ��׊u�i�όV�^h5P륽uy⍯5ے.�b�E�o�cg��������9c���=��ü�GsQث��kҰ�$�f�ظ��Ql#��rS���%����}�2�ӯ�Z��nG]ҩ~^�}�j���k��ځP�����U��mn�v|S�59�ڧ{3U���\�����=���R���+�
���(w�?_DM.�k|O_���PR6��+q!���bӤ�Ϋ�j4����
������%ﾛ�:�o���Q�}���K�+p=���k&Ҿ�ְZp̪��N'n�rD;�Zd�T)Q��5��I��{Ir�q[u�3RR�i�g+�m�.fl�O�K��nE(�=�kF`��e�,���I���\���c��:���OJ���rl��|Xz�ٺ�!��<Gga��R�ܳ�k	u��D��s[�.=O%jfnՔ��V��9��D�v�!K����=�9���k��ƯTN��2�����W"b��N,P�z�i�*T�WL8"�յ�s�Ӂ�Ca�!��	yQ���Jz��r=J�X�����qK:��ց�30��sO��2-��I��1W:]������ʱ��V鹙v�B�HA�Ӄ�h�XFŹ7:���ȥ�ֹu��ɜ����t;��ɵg.�u�1&�ԟ5�����K*�w-�����q�wh�:��]�pf���\�r��pD�o���������@dryk�����,�|�s+�]`�qbע]KJ�ʱ�f�����#`�z�}wo�M��Q�|f�2�A��Kͼ�ښE� �Ұ��lY=� �*�0��8�W(�wZ�7�I���hU��i�sgRQ�����;V^L�%n#�5�-�����Õ�(��o|��d���O��[�F�<�X����`�Ǎ*u7N��9kR�Y��Y�TM�xb˥��AX{��iv��;3��J�ٮ�ʟ7�(�<-���zM�����a��*����)���<��
N�7$]�n���s�vM����/8��s�+:��>��t�=��wk��YI`<�޶��RA\���:��(�wV�y���N��v&hL�K���C8�d�<�lo�����juB��dv-C�=/�uӪN��w{g�!�����l	��۠lovܮ�փj�%|�b��F!�<y���kz&�޹rk6ˡÅ��B�;]#���ޒ9U����Y���o��Xt�l7V�Ek�z�]��n��}*�	/H��,cqz���;Cp��m��7L�I\p;�}�3r��)
�-���Ms8���})�Kx#��ں@Uݒv����.p�T�S*V%�ا.W"�����a)�1���Sm�'P�JvY1�¦�k�xp�:��{F�`9��d�]0f�q�3�2��e����$yc�o �E����p�j��7��D��� ���7<�̭h�zm �L�u��D�V=��tfSB����6a��C��W2�Z�}M�u�uٰ;A�9�Q��J4=l�f���Y�u����GV!J�.j��S(���;�˷MR;7u>������̽:chky�KZ�M	v��]k=�,�m�]w�m��`�4��g��5������v����t:�0c�ͺnO��N�v���j�,��O�|����-�Z����k�hE3�bXѥ�`��F����1�I�E��EpSz�����u���j�u�����v�R�K��ef�oz��>
�'�$�#9����siF�ES�J-#(����QTyKǈs5��)��Z
�"�%eR�rQ9<�^1HeEH���(�E5#���$����A0��-C�Z�»�qҨ��+0��+V�d�$,�%�"�i��!*��v���R�%EQ��sju�iha�!x����;���8�Ue�B�TЉDP&�O.q���L���#:��*��$�uR��BM-N�l(�W55�]9I)�Ja8�q�ԃm%M���C��$�I!Y�j�:L-��<HqPD(�H
��WMX�,�I!
���9
�ڗ3;� �uf&J���K�a�5�ٗ!�q�s)VZ�H�E"&�TF��f�.DY�U
�"������1Kf`��,,iUD&����"j�fZ��-g-��C���0�C�G�����9��k���s9�ֱ�G��ϲɬ,��ﯜ���Vv�]5�y��" o���#�j@���rs������}�����]�L�Drr7i[<�%��b�1��m�R��,Zjm?k8���'�O=:6~�9N�S}r��X;��|��B�縯�$Ż~kV�'o0��9ū�O���zy����W�����9æ�а_r������ �닄�r�����ƫY>4�'Pw}`c���w޶V
��Ϗ5��絼���E���/������f�fZ�.Z��-��줦��,Ai��[��%D�	.�Jz��6x���n��Cm���+���W�~�W?Q�HJ7�9��U'+}�S�>�����k�eCU�p��T=��w�{��JD��4�^b-��������yF_��yP�}|�v���Y���'HUr�������U�ZR˒����b�nʟM$�uaw[�}<�<<l��<��ҭ�`y9�d����_G���B��nN	���fXӫvc�1�
�xeݎ��=�N��-����2�Yƍ,��m,��)�#d@n�h?1S��΃�{�i-4��êu��ѱ���PtR��0��cx0
�d��������)����y}��nEӖqJ~����%�����3�	�O�h2�cX�4PU ��<^�����d�U���۽�n�.�פ�
�y�$�	�Ԟ!�,<�z��U�ҼF�V�{�Wk������=�k�̷=�i��\�=�Pa��A�GH��~����A7�Gɓ�Ϣ�G�uu�7��:�L�8>���"jq�bα��/��&C]�O���e�l��K71I��LE��+ϕ؃P���۞z{��n�gLt�f�8Ùc|P��W�۾z�>=H�X�uμ�(ڧڊ�y�ޛ*x��̺���نV���ٿ>P_��������NI�������mez�-'���JT�ܡ*��W�R�c>]��w�;�S�	"�d��G�&\�I��+<B�����G,���){j�ťNG�	���.�⛌����Y��zgQ�;������\[�\pN�|�f�b�}x�G�U�uV&\JGD�#g��? �[X�r�v�q��<���z�{债8*`D��J9P̧���˥���Y����q<��ʙǝ��%w�:�;�\AK+��aTE]6�Y��y��X�M���dqG���ǜ��YCG3F{�0r1�r`j;�q*��fܿ���̳K(�}<Ԣ�׭f}��4��m�p�zkϻ�*�t��TC	ƫ~�h���М��~�p�z|�iu.���`{`�/���]����͜�U�˙1�>A��3^Į��|f�����g۰r��T��jY�Sf��)�U]}���eL{�8ܘ4)��¼�H��G����8+:���u��G��sq��:<��O<�לj\�&��b������K3�1u��;��O��K/Q�f�[�+�i)��rV&T�ƃ���f�`�XK��C��G��W�V�z�t���c8e	�������յ���J�>��&�&�Z�k����ק��]0ݗ+��=�noz�q�[V��L�z��_c���k�b"gl1�x����J����?���H�U얽b��T�J�t��ڬ���xٞ��P�=��%���ׄ�a����>z��ۂZ	e�;1�wnGڥ���yW)
�U��IvC��ucF���9»*u���^ި�e=�v�}ʛ���w-�-�c3km��*o���[�
��C���Y�=N��;�)?R��돍�쫕�?a�)_� ��/25e�7sw�>�^4��ŝx����u&[F-�yaM��o���5}A�'�c����٨y�c)N�FV:<�����
��.x��X�<��ƴ�<�D���o�y�>v3��2C�/5�o5P�� +�J��HoUs�p�$U�꩖��:|��R�0�����ޅ�����5���[2	??6?UO�-�A�]�U��qC�u/oφW�̓��/T#�3�J��%ݤ�r��Ӣ�^A�iױ+���]�B����CJ���y'�d���|3X��s���1Vr�`�t�T�Z)��4�K��ŷ;�g2� bj��2��W�"����U���ɤ�D���Վε�l+��$�j~�������m�Ɵ�}��{q��<�x��x���"1,��2Ӟ�:[&q�����Rh�9�ǁ��rW:����N���S#<� m�f�Kre8���OUj�2�%~H�r	/������e�k�O��oZ�d�8-�W#V*�;d�T�;xW%sr���;�v�W��^]���U���\�a��Q�=�it�|��F�<�&p�Q��z���|��*s	�E��gd�dk�*-'��9����3z]"b���]�f?'�E��ͩ�I�*{re�6��@��+i���YF��e������R��D����'R�xp�]��X4)w� �2�iB��l0�}^|銵ˉ�潽:'�g�h�&��H!M��A�P��w+�)`jW�q���oI<�m��y~I���f���J2����M�9`[�0���Y��(��rO��ַ�+~)3���ٯʃ�+�tz�s�8���mY΂���������}C][�{$w�t����uY:������ٻ���-F��:����?u'}�]�ʯɓþˊ�j����U���X�!'2*�����}��rX�u�l�X��V'b��ܿ���d��=�V/��r��a�11Q�ܾ��7��1��J�>�n�{{�k��w%����3�������kcz��i�4�Np��E�i�������7]��7�[��|����Wn�S0^���K����}�-�
���]��1V�kY��}}j�a�����sĂe��?���LhqB���m�-_=bim2�|U��hM�(��%C�q�e�U����oW��q�,��A����{`�rs�ٶ'c��N�u�䇂I��J��|��x�甚�|MqFTгN�ۛ,�R�m��d���F��Q*���`X�
�>���h2�(�^�`���3@��F_
�e����m�4YZWO��еH�)�ea�sabL���)��A-+Nz���D{�i}���w�3�^��.��{�/�?N�o뒁�M��A�a�V[�rQ���uxW|�n�9���O	�X�;���+�rY�Q�0�����z�i'���9�Y�}\}�7�S���f��+y��ga�ݞT�J~����ghª�IKdV��Q��X���葫�c���Qڏ�s�K�Ĕɷ�����l������۽�^��f�����-:���%�|z��nxEØ;,(H��9�,�D��'��uT����#w�3�KR��S�xq<3{G����"�E�̢�b���@պ�\�>g%c39Չ�gl-2�*�
u�.�&�/��'�`��eL��2W�bQ�V2���`��:f�+8W|�����Qս<^�y�ϖ3�����ح���a���ܔ��c�����ϳ�^��|U�P��Uӽק�-|7x�v��_T�kے�/��]�~*��D�8y*��J"&�	���3���5�ϒ�E�b,L��bo�+��,�v�,�80�ªU��vJ���Y���w�K����N�]��3� �F�GA�����Rv��'6!e�pnu�쬱�pα� -��g|7��j�jŽ(t����$�˃��<jm��5�UBԫ����#!]6ah�IE2I��<m�Zr�U^��E��^[�i��\����9e��B��}S��]=���ѡ��I@qcf��8�7���U䶛9M�X7k�q�όQ}��a8��2�AjՊ�::���z?;�[;��s���+�דL���o�(&-�"�Q�U+hǼ��_�O��ǩ�/�w��W%�%O�SYc3�HaY��6�U�E0X�uΆ?^f8���ze	/�+�K�^̢�����7��l�1*7{k�Lŝ5�wh��0��[jf����nZ"��ڂ�Iw;��lgOu۔�b5+�W����;S	`յb%؟dfS��{.l�C���x�X$�Ĭ�.�t�C�ﾪ��%�FE���v��D�Yؕju"i� ��yn䲄��C�g�c�)������?.��?:үi/V�z}<M.�U���zC�r��^v���#y�C>>��]�^�F=�!R^!�Q{Y�3�ί�ݖ%ow�naKA�B�e�KnSf�d�Ud�W����߱��i�������T�l���1*�]m�M�D�>V�E�(Ŷ�m_O{�XLG��u{��0�x�KR)����1�]���&h�ٶc�9çJ���R�z��=�a1�㈽�Y��;>��;���5�f�E�l9���S�)�/�՝�o�ُW;��wG�-�%�v���Y>��Q�<���]BM��>���t9S�/{Wq�يn�mJx���*�o��\[Ax��|��U.��&uJ������wV��Ǘ�샠�gzf+�AN!�^�*�j8���K�{i��_]Iu�a�9ގ!����/�m	y�W�0�L�5���v7�c޴1���N�Z#vK���גկ��ū�g�����V^+��Gk�R;��lU@$G� �i��u�GA��9�kEnC�n�Gliy��w����Nm	�mj|����g8~�3���ܭ�U�J����k�b�y����w	�uo�O9Y=�]�|.9���m�;&���N��2zV`إw1<����e�:-8{��ϙ6��ɠuW�/�U$Q˔�v��W�:�ɕ���	v��9�3H�a�U��4yG�̫�l����t�Oς�x���ܱ�r���4��έn�`��+¤���^�#�ɠ�߄��}Cycf�@�_I=5��ך�������p��[�ދ�R,u���g_���%�,JK��^�k�j�LIPc���o�T�~�r�z}��n%b�յ�5��������Y��q�}�B���PK�6j�4����A\�+=��a�=�c~���?h�����k����]@�:Qn���"�{�*\�W�͗�
�U�v�э���~�w=�B�sŰ�d�2WS�6��y�!hhA�,�Fy-�I\4e�z�Â\E+v� l)�/��gN��c]J���r�Y�7 ���@�jo�������\��z$'ۖ����.�
r��}��g�=J��W�dԌ�$���=N���zWb��h��^�0%��rt�Q�gw��Vr'h� nCpŹL'��K�G�.^��#�����;�WJ�VS7:�}���0��X��꿄�zk��Ψ�=����L�.���)m���a]k}����{��7i���\[Aqߏ�
��a��.����2T��a����k��M2f���~J-53a�6V`F�T�Pn����GR�~��o��=��銵eؚ�}��=Z�uRj*�Zա>�c'���S(z�b�T�T˴�8�fR9�'$+�i�g���uVՅ�sH[ٯ���i�kϨ'w�<㗛\�b��m/Vɚe�-4�IԮ�[gҖ����Lr�������+׎vYcA"t�-���P�>�uW�ї��Yj.ǖl�!���s~g�mc�L������`V��z����-�#[�>�%�DOd�+7�Z�����^|�*I��4�t��T
rZ��uu.���l���_lM>S[1u���z��=@��h�E�����mr�c4�z6H:�1mb;�աFlb6��`�G��5r� ���}yݿ(TP�g%b�Jz�3����T��F��b21�p}B�ֵ�f!)��oxr�� ��V�u=z����沺F-���l�N6,�����<z��;,/�76�Ʌ[�@�8?%��L�Tr���b�T?f�L@��Նf⮷|�870�iP�B谨�m��jup���������7�z�6[��(��7;�Y�б�0�
@2�M�0�ǣۨ��y�k^���d��렽{�2O^�f�i�"�{��sf��^����W�����5�	;=�=�Xr
9Սu �[��78\!YZ��=��v�`�n�e&B�՜�ڻ�xw1��If˓���kCz��q�f�Ԣ@qG|OG34t�rv6MܾW	u��a���S�;qo$o �}i�I�C0R�N�+�I�]ٻ �w8�fnWIҚZ�:���l��5�	��;M3�NXY�a�+��78ک�Jk8��s.����=R��6�<����4���>ղ��zefK+^u��FɅz�\,�F��ƘV/z%��[xn�M��R �q͠�]�|��(�m�q�.�m�@)� ����D�`˦��gsx��L&6'm$���i�,/M��/���k�b6L]�2^uK�Ů�=R�}X�F�W{/t9%�YO���8����ʴݩQ��Q��*��u֬��I�b�E���|��,o364�5�i�t�^�ok�eߺk���j�7#�XI���euL����YVD�f,�;3mlK��̗��=G��;bM|>=ʙ���f�8��=��+8�9:g:8�lޫ��@ P�Z��D�Ya�<�lr�ͧm3��dt�+xG%�qܵ ne���$ff7�b� �\�N��raf��*,skL}���İ����ε50UT�*ں����:m�<��n� T;،���iع�3h���;�y*�F�m����a7%�Ea�Ьq�/'qV�d����S!w��١�&R,����Җq��0�O�dƙQ'y9���z��Lqj���]�­7�{���p��4�]�.Y|Q����on�5ȉ����igwsv�.
f�6���;�քB`rM k]]�ޚ<���Ff&+�8])*����*'T��=��n��R� @�"�;(h���j�}W`1�6��u%JW�R��d���z�����捖@WO �
Y/�����Tg)���~un�����tɽ>0e���ݗ�ɳ8K���L㋵�ѭTx�s��1��h[�N)J���\քPԝ���}��-�z��+M���A����5jf�Y��9�]�io���30��	��zƺn��[Sm�����_���r�ѷif���)�u�w�Wu�����,U�&��8�J��0G\:lE��Y���jW$�^�YRٕz��l��M��P��u� ���l������THB���*�Vp�)PV`��.����WV�;+�E�U��&A�H�EA� �Յq3�FHQ%mD�$��X�$�[Y5TE��3i,�ZBHr�L��!�T:`f&�����䒘���a�:�8��	�%�'+%29
XiFZT�-.)%TDDp�9\I&TjRq*�NjB&�
���&Y��<�!)YV�4��(�E�"��ҨҊ�r*����)r�/.r�U(�.�f�Z&I�����V!Ȫ�M:j�$0���Tt�Y	(�u�b�4(�����$*�-�O&�q+J��8�hal̊�,�5��"V����F�F�d�¤��	$��&�!LJ����%デ,����
$��PEE���d��jR�E��!"ds�l��4�ea	Y������*b�P��
g���+���ν�[��6�z�8~��l�}����k�,$�8�Y����q$����aas&ՙŎvc��Q����&Yc�4��T��՝s����Cve�#ֲs۽��V��L䚦���9�|c�Y�i�>��OT����¯Ӵ雽V��9x���6��5�T~l�J�X-�Df0O��g_����Z.9�����ONF��\�+N��g����E3�l�t��ߨcxi[#=�pݷ�V$��:[��tUUY�y���Z[q;���w5��N���ޚ��14���2C�j���H��P"-�vNFV����o�y��
q*w�2"1��.�z�)�S�t_��)=w���y<=o��\�n�g���K;�b���l3!CV.i+˦q����^o���,�L}�n6~}��;����"�'6wr�+�:H��O8)�Aq	ܙ�n|1}L��(�a��6Co3����n�r��j��Ӆ
�e��{Az���Y��^)�l� �z���ͽ���D�%�m�v8Y8�71�,-��G��h���i��s�ʯ�hV(w�[(~/} u;��{ea�|��c���p�5���X����
�ۙ:G�ݳy���CkE���n��-͇���-����-V���+#(]�U8,�;�=���#�ܽ���8�{���O�^�s�N
�S{�M��t,wY�g���:�ʀ�/�l�^ً�Pc�6�H�u���}��&Lkv$�ź�b��׽Z$�,ǔ�m�8�\��>�Tʮ#:*�3�+b������j��8����#��.��-�%�Y����[.��&�86�6�[��� �i�gm��/�%�����;���F5tq
�6U�AM�!�
e&]�U���I����Y��{rE����R��p�m�y�e������E4-����cm��P�[�jZ�Ƚ������C�WAAM�Js5ӏ�L{�'���tm�K�������F�ϗ\^���XZsL&���Ł��:f�`���#��%�������;+\+CbHתG6�{;f�QW�i�ܽ)���"Y[����l_�C���3�"3-�	�ݖU�T���\U2�Q{���$s6FO8���wG�*U̩M�_�z�xlT���-�.���ݵ�S�sR�s2X�&�lV���f\j�'<:eՔ]���a�!��u�o2C��Khn|�g���K��U���F���ܙyn�&xT51]/�-��3�2.�z�SF��l��qd)zj_��^�[���ت�j�XKAS�Ƣ���(�͕��ۧ��1
�B*��]l�u�G!�(v!|ۼ��;̧NF6K�V��4"��u�%��wzP-��:����0���ǫ8&/1�_t����0ݕ���&�y̧��86��CFd��cyk�O�֗K��!u!�L��4�<�z�y����0��G1��6�e���`n����^ލq�)�ቮ�{f�28=gJz0Es�Uý_Gn�� ��s���6�y�h�e2	���^�/����o���T�~ N~`]d�\�E���e�vi]z�s�-��*����|{�I"��W�!=��Sf7��t+�qx]�\�=4���9]��٦���zm���m"�{4Sg`�z�Y!�E��rq��Oyq89)Cr�9r�.�w	S
�:��bb_���3ĩ�j���{���� �E�27]�~��7*��I��;���ߛct�1k�$-�,�=���ܧ��j��)�Y��e�Q��WCl�ȉ��1�;����M�c��b�(��{i���>�
���U[��u��n����Ϣs���mc�L�ڼ�[
���-������wY^�mg�J]��I�dD�d�b������[fA&�'fi#_�F�)wǖ]]\�n![:Q�'~�֑a)g��w^W@�W��A�rb��?h4
܉�H)3OVJw��zY~��~Y4=t��ˤ7Tʄ�T������2�����wV�����VT^{��:�5��!m�B�]|$�kb����'{*-�.\=�q��tչNC!�ݠs;��� tzX��L�T���؎�w������]×D!�;v1箕K�.��
���)�
s�q[۪��1������St�8+���jݖ�S��/�����e�:��!��G!M��]mL54��އ'���ݸ�&�H�`�Ƕ_�s��N�SB��j.{�/�N����W�����C�=����V��G��n�v���4zI��X��v��=͙����GK�ř�wO����9�@�r�(t���&����g�ͺ��Ϛ�2٢��*�02����Ml��ɗ���3#����v�5��w���i�wG��2����w*� ��}�"��^\2ּ�Ѯ�ܖ\^V;g=77<?\�X�m�1�3����A�͐���8�l�LP��h]t�s�`OU�n��NAi��YSUݛ����Ý�eSv2Q9���yH"���)���*0�6����SFJ{T�e	����B��FTYY�����>tV��xV3ך�z��Q�z[+9���y^FR��M;�������2^��ps��a���ه코���R�"r�q��vQ}:��K����n�
�������w�gP�ʿz��:�g�T�5�C��~ނ����#/ìM�r�v���N�wtI�g��L�p:/tK�E�ޚ9k���<5W��4��sCtv�ISN��Z�.y}CT���D�}E���D�[����m��~�����wQӕ��3+&��t�0/~��%�%n�� ߦ[�M����q�5�s�{0�����m�Uw���q��w���{f�r���mֹ{d^�,i�+�b�(��~��en
q	�U�'g1��%D�۸le	�/�����8���^��OlL!��.�Jw[�����j8��kZI�� �7 ��q9���)i�ޢBw�lΔE�;:��J\;�'�.�[L����^\�të��¶*I�{��s�߽�py�Z�q�%Ԑkn.d�~큃�T��g자��<$6��6u#l뒬�٣�W��曭��3Dqb�à���3[:�U	�\�p~��Z\ټgs[	�D؈缸ʙKS֑�}��i�s�SL�����{��&7G=3)٤-�d�a4wv��g���i���-|]�2ܶ��rb�頴��?X�V���[9"��o�q�y�]�ې�B��-p��G6�wK:'@���_{�ٌ	�~>�Ӄ�o1���dlH����:�t�SZy�KU�v��/r۪�
c�.�E���~�2]�X��v*y΋h��ʼ�t��'3#�ƳA���_�p基q?W���DHgƳ�S�a���U�vI�neN?bb�(&�W�����_p�<m����M����Y\�f�n��
�v�b��ޫ�I@u�kF�Hv�R��.R4.Q����Jr���t�>�U?��F�Tf�j?N���#��]I��T�fGCV.i)�uV�c�Nؿ��o�>᳈v�f�1��ڝj:��k����pS6N"[%;�5����s������.'ˮ���kb�:*X.�x6��j�nud�J0���;�f���۸�	�^D����	��� �X��;�A���gigx����}ԛ7�Ý���9�]�72����%�_NЦ�����y�U;�i����]�2��3��Gy�bqF>���/�m��K�̐��E����٪e^���Y�C�w�y~&'OZ䄎�y]�k;^�����zc���l�-�*׽�\�-�yT�mӃm3n�սL���xe�+%K��){������dF��m�_���#+����f�/̎� {a�,�K��mǲk����?��vM)����;����Toz���^��U��Dc�-~����
�������E���i�+4�Z��M��w;��
��`�Sm���_V�=�w)OM��6���%�����J��C���F3hLkQ�m�њ%�`�����nf�`��莣���N�OJzIޖ绖LT7L<��c��)�<5��[*��f�����
ِvri�%��a�B��8��SB�+� V2+�[��;MՃ�<!������K�t��g`!Z�`p��}ܩ��)�\�v�<[QvO�:���P"��N��G����d6Ձ;��p�[��ޠ��n���t�S+f��)�!ܭ�i�8��l�˄�B��#-�Zb�Uw2�./���z�BC\����veCʹ�!딿�1����܇���,��l�!6u��¸�(;��1��"�B��-NK���N��=z��6�n��r賅b=>��ow^e��3D?3f���ܳY��U�{n��q�H'���:B�E�cz�r%���=a��K��c��0�a�l���4���X�D�J~�|0�,WC��z%�9V �9�d�����S;�^���M���F�-����ד�)��\D�%;��G=�U8��o9��f--��;tZγ��)��ƣ���:a���k��W��|1���	�2�g�R�u�(OA�٢K��E�_;��A�ڥ8"���P���'�ǲcF�@z�����q��n8�o5n�[wh^w>��grc�
9�z��EpS~]�܅��M�{kHT�n1�Bz�e��;�{��.�w+�YyOz�5_��	���z)�C�W��g�RP���j�T�l��PE2�����oS��Έ~;�nr��H�[\#W]�/$�^�w�u�tJ��y����uҏb�Pt�%\'����ǂ�<�2��A�ӯ5挦e��G��+.i�q;v���G�4�dea�Igo�M�:GE�8Rց�=������n�c;�6��!�.�GJ�z�E�y[/s#�s��55=n7�3n��q�5�q
���s=���)�7*�F��3fr"�J�dr��������ɪ���Ezg]�cHw�k�Nz�eXOCWV=����ZCc*�W��l��x��4Aj�sލ��Oa`�m��i����ߢZ��R�y����quS�:��ȍ�.����Y=G
]�;	Ύ7�צ����P9�TOD~��>���Z�h�����c�]���b"����D�L4v�5Q"�@#P�v�c�]*�z]=W� :B�'��,����s/[W�zӢq�ӽ�7�k�~�(Mn�*S��/��t�N:@w�8�����ͦ�������ղ���4�9��A����zu��N҆�=���W\�0��ͭ�8_��"�s��ol�~�kFh��M�-���%��>c�p� ���J�:_���1U����|�E�;��Ǌg�0���T����`eWӰ1�����0�=���ji,��*(�Nm���3s���ᣭt��j&_8[2��y=o0D�L����2YW�'�ShZ1,7�%�h���_�cɛ�n������\�vM��"<��}n��X���.��E�ZT�k�,oV/��0�>��1�'23VrX5�׏�kk��t�а���c�ŗu��Z��ss5���і�]�5���*#�Ȃ������L�,멼j�$�m��j�<2~��]2��̆	���h_D61�2�5�㩶:Ę���ӥ�m��"۬�zuGh.�"�G;�5�nHE�w>�Rλ��f]�+�p�Ǯ����[
��o�fc/T�r�&nHη�m���9��gC�E{Bw�*���_C=�.��}}-�ƣCp�h��_��:��0,a���-q8��g
����a�)�i;��QJ������Z������̻}&�`�l*����ݘ��n������~��Ui~�և��G��%gg���]1Y��H�����4�e����/�l���S�Eĵ���S*kP���3���c�M��M=k�[ P[uԟ\3�����.�D�u�l�-��*g�ظ��,DZ�%����Sgt���$�e�8ݰ�SG_W=��,p�=
]���GQQW=����f�n��x�ɷz�BNBs����t����ZBw���J�[?d��>W>���昪���ۑ�t?U��h�ݿL������#��l�e3���v����\�����X���$����zvu����oy�}Nڶ����r�X�Ou,��m�_3��]ǳ9��2�I�#��S�*S[G�E&u�5�xn8��^)A�Kf�"�5�ո�vNۼ�Ư����π��vUk7FtDpV������T=��b�^�u�qq��f����C?6�LCBB�!�]m��+g�X��g��&7G:�f�]���X��9��y��p��$>�py�M��de�G�J���)G�#�U�
���fV~;�z�oH�M���<�j�EtJ7����=4�
�K(�ws^]��*�]���"]=�fHu>�����)<�
xA��X��#�����=�r�K��h:�u�����Ylt/1�H֋�wJ߳�	�P�K��)�'��S�O�	�DN~�UL����b摡tE�o�Ɋ����v���������,��'�)�'"{hX0�9�3��y��9�nJw��o���)ζ{����%�K��J'#��-��nl�a+E��Q��us�������	�(� �O\�:�������I����g�}�[X���"�ǝ�Lm�YX���T�Ӵ)�C�*m�~|�=x�˦�&�V�:^�;�U��p3��]��lQ|���L��b�B|�5L���S<���s*g|qy#@O|�W`�gB�=]M�)��k��zO�{X��'c������^L�#�o��!����zdfc)�Mqӣ/?�Wp݋ז%ڂ���ڈ��Z�Q�} tDū3u�l�aA�b4z���LG�6�y�}�Y{G"��V$��IY�G��T���Y��ݧ��2&0�<軲�M� �b��GUGZڂ� f�8�2�,�t�kMug׮���9��X��jI6L�4#�W�V��J�+�4�q�0k��GA<^oY�Ɋ�*ث���m��\�����c��p�V}��J��D+{*�,�u��0j�o�]!&[z�˶�-
�t�A�y��y��
�]]vP�jj{�]�{�@��P��̝�����E9Q���'R$�i�=P˩$�4��K�Rݘ9�KF�{=��^�%�=t�^�Dz�3}}8s�Ԃ���V9hA�yx��Ib�A]bg���6��P��TV���[h���-�ݖ�6B��q/ݺUz]N:[O�(u!�E�vM�����e�6�wbH�a9��$��@rj�Z�0�a���w/��2bx�T:�^�������K�PQ�b�7�w�];����t�\�5r�f:�lp���o�5���/sftm�j0�H�:��N+{�5�nZ�]h̬�����)��c�tP�r��j�<5�{�E�}b,ݸ�.�]�0�/� 9RJ�Ds�Z��3s)����MVԋ�*�wP%��5Ĝ��Z��ղ0�d��*_56�d���E ��8U))�Ĩ������YbgX\���3��+�5w�8��������	��x^n�������#�S���[�Zj�7e��qLZ_h;s�ﳲ]v��-��e�E;����I��Z�G��9y '�-��Y&�1���U��mq6�'�7O\hu�7�8�C�t@ͭ2������v�ܸ�4&�5).�nu��5�ܘu����MضP���]ͼ�U>5�q�v���07�[ǻ��DK|�#����eSU9�������}�\+bŤ�e|��#���\�*;�f�LU�&r9���p�`�Z�Ufۈf������'z6sX͝w6I�;�[�� �<�I˸_Z�5ѭL	�OG+};�'��ӣ�#'o�vg"��u�w>2!m'A��n��>�y�3�-�	 0�oTʙ�b_cOk1��U��u;]��\�%�du��v��W��#Ja�������җ�D�ku�[Jl�94u�R�Fi� o�3��|Id��G��O��gPf㫛�_�T� n��h�z_2k�42����	�qfL}$���Ld���6�p��J��l_��{%���l4������.۝�6��1ʖ�8�4b�܁%��řOA9�|��%�аj�Ù :���[B��Uj��+i^M�7x�����
����OY��:'jU�sG72�#X
�k��p�ɕ+��ĝ�f����s ���ݹkk�v�Q}>�b`Pf8-,��|h<{��-��NQ��u� I	 �$��ȂN2�8C�����Z�(�@V�]$�!i)����BuZj'�8�!��ȪֶY��aU��#��Q�R��P,�AI*hW�*��w9��
�b,�Q����D�����eL��Bܡx���*PN*QjHY\#���(QW#E2�U�h���I˦VdW:�q(##I! ��8��aW9U��Th�����H]�,���	�*�PE�(��-
�����"�5G"�hD""��I�
"4)�\�"+���Uj�q9r�C�"��W"�Tr"��-"V�U�B�8x�D���Z9C�)E���*��NSD+�r�!EEFH��(�dDEEp��W(�xɹk#1+dTȗ�A�o7]mxaɒm�ʩ�:C<�p��!��p�S�J����m#��f��c��YɉS�qaY�a9�[v�I�:|H6�[�2�,�?�Y�cU���C�g�=���pDb��"ՙl[Y�N�B�+����q~܍���ū"�s��L�z`���Bzf���[j�t����N�f]��_Sv�;.%�z��ܶvgS�^���KF��.�bմBA�h��!9&����)O]��gV��n��'��e��*ߝ���[��M��`��\F��s0����w�^�; ��D�(�t�^���Xs�?�fų�:۶���uҩu��,�`���Y�!�lq#2y�D⦜��U؈4�x�6���YS6�6�`���us��˘wU
�2����Ӳv��qu\�;k���ޭ�������,��!j#8t�sK���]�Hz�wDn�W	T2D�7.y4j��4�x�$����[��qv3�/�7�|/�L���P�K���ҁ�~��&�1{�׺h�l����1�m�*[���+�s�f��%�S���<��b�dt��x�w8V���fږ��C)���<
�-�^����'�SoF��l�����i��i���E��X2�d�,��m�cڏ�ۉI{�p8P�H�vCO^Z;A\��l��OYԤĩ <\[w�kxb=u�`�}c{b�-u�ɔ-���w6{��(�J֣��'�7��Q
d�}�Z�un�..���{��U�m��H��Z��܇��{��Fn�C��O��U>����}�Ekt�#*2YX��do&pc�i�p��Y�����{�'����g@)��A�:yƊl�ʇ��{&4m��C�
���W9LV�O4���S��qꌊr�y����K�57�et�h޽����=�s��v9|�����-k/�y�<sdOW�Xaʊm���������pT1	]f�od�V����^o���O= Nm��pnf����=5�b��:T�=��������gt��qwD
�`���m�l�1�v��
�}3n�4�{���3\Bs�
�s������l���M�!b��uwTCu`��%��K��61��~�@'u�薶yJ��Jl�DQC1��{:)n�'r���j�|3�;\s���맧�|L �å��	߶!����*g��بh,ꧣtmT嫭����X��K���"4b�sF<��V=�D(��5�!�!�Z��k7nH�px�ɬ;Y����8E�3���Gp��e�v����3@"���^캇W�;��� �d�g�8�����p�4��k��xp�}�6E��ӼK��[�����kh�Vt��\~�-q��#�����h)1�¤Y��-���w�kLw�Z���x��Dq$���r�u��gV谫u�H1+3k��Vʓ46��0N�ز�s�)�W�Ɔ��3`D��1�tl�X���/�Ф�CS#��S��k�Ȫa�El;M��5�`��f�yfL
^St�m�p�FrE{s�OX�$��'��ݪ���gS�[	m����c��]3����z��6�*Ye5�`eM};[��M�ϏQX�Ϯke�q�U�5��7KI�~O�xj����j���Ge;���':g��~���,��{C��3+�v�i0y���@Gc�f`�����b�q���L����)��^��4d'��L�=~hI1ʓ�;��^�`���M�;�Q����Q9���L���xȰ{�@���L��N�E�gM�U`�9S��Ф��\N��3>tk�{�*���_C=���M��M�4u-����/���EZɣ���z(6�n�Lo�)�}q8���w���|�)��J5�$��{w]������5�b�\�+/�Ol��-�!M� 72݂Z�Jzk��+�q�lO�A��g�� g&1�%�n��XGy��7+���+���˴Is~[/*)L[��-n�,��AA�,j%�ћ��t޶��pY�;xU]��v�Zh�ʴ-#y�F��i��׌�2.���7w�H��L~���i�������I�;[�PЧ:�Z]g'��ذ�;>K�|F���V"�|VL��f�r2�3��!)��Vc7�b���*��[�s��6(l�t�^��Pǘ���1�o�ԟ�*2����Ci�;�ޕ���!�ߤ�+`hCؘ �f��n;���L�)�C����ɵA �lE�l-����~&X��!����x��݉�B�U�zȀ���]�wBNBs-[8Ꙓ�H5��K�h�r��^����kC��o��#��!M��_��f�<�Px]�s���u^S;����!B��
2��x�[�q�KZW2۶��+��;@������=+g�[ �F3��3<e�v��j�b��K�3
$vFO8��.���ٔ��z)��ˣ�?X�o+c$c`\7zr�8�h��D�l<�6��)�^�v'�2��~�c��{�]�� .c��E1�yY��cxW���Թ�'���5"���I�����B���w�-L�?_��w���Q7<�@eV�:�N\;=K���0n�c���L㚸��`3~�Q��W�3#��9��]3���"@�P/F�ڛ�;�9�O��CP�L|�߽)���q��1�{|�%�%;�=Mύ�s���zP0%(b�o=���R�`?�����ߔ���d��̃�l��ّz>,�IB�x>�ne���T�oj�Q�0�n==r���s��AΠ���&��)躺�tE���S%�'l�w��&���1N��5�C۝h�z�7�vZ�wy�>aq]�V�����;��ނ4�t��K���_�3��e0��d����	�X�lP�[)��ՠ��ݨ�����Ckis�UY����w�c��Vڦ���N=rǝ��:�2���C,���Lء��(wg�R���F�9eq}{�iT�K��d�wV�=r_[{D��Y��n���b�!>Y�dg�n�M�[74�3p�0��k:B�b9���͜ep��M�SwZ�{m0�Y.�i�M�p[5�B�3���V]�����͹�����\)</D9��=�ۺF5tqQ��ra�L5i�j�:��f�s�;Վm��u�ޙ�xi���P�OMq	�bUc�F�#7`��DsN�[� ����ՠÝ��NUhn�M"z6]Ҷ����BA�h���%9����\�=r}���Ԫ��YL�kT���$k���f�.�,˫����X�҃��l@z{h=&ú#��5��;i`��t�7`�4��3nѮ�;$�V�������Oj�����_�[ �E4�x`�yN@��P�Y��=td�3{���7o��w��ծ*Y\ʐ�ܥ�'����H]uR��+�y|�錛���ț����/� =����o���'��#+eD<Ӵ�g����9�������i��HiO�պC[�j�ն�us�.�d�7,�7�8kj��������I���Jo��ӹ�m�
���]ʚ�(��ƴ�X��%ܛm�����M���U�������<7K%�H[-���!�R���$=�m��+��*�vO;�̦�oْ�A�9ќ6�+�^I3¡���~1l�1��N�A��ɞ�Ԏ-���g�+�$h�n���`U�}��c���O�b@O,�e�����zW?im�p��)���?e3����"�c��h�nڹ���{EoF������n;�K���n����8���Cقw�L�@�=�m�y�h��L�2�2YX��W���M
��m567�vc���z�o��ʋ���)���P�̻��� �OV3ѐ����h�o]�T�i�m�#��;�Eh�|��T�-EM���]M�Q�4�M��),���R�e���2/���W]�7��q�n'U�a��P�F��x��3�m��7�7�,�*m1"/#b7��f��7Ї7(�
�ӓ��ۼTo���,!؇J��{���)�7/�c!1f�:���)ŵ� 2�Z��ڎm�Ze
S���ͻ�Li���(X	�l�	�v�������1�#2M�s{���uv��n�F�{��n*��8����uqS����ǋ��m��\�V�9^�%�ʕ��d�u�ŉ*��*q���6���[G+�Z��&&�޽�ס�ɇYIv���v�0^���ve�b�o-/�E��%�-�	�M�{.�Ԧ;��zB���t�T �͉kg�JR�4`�Rԯ������JҮ��5�2*�9���W��$Rǎ}ղߺzS��p��tAw틑t�v�*�d6�5�Q�f����G+l��%�vYW�Q"���k�}f�R��g�+|��P�8��>���5}nnm��W3LCܳFN�v��m��I�i��5�9րA]쩇�.��k��_bˉ
�'��R��F�M��_��7A�ңxc�0�81�=coN�*
�聅�oT�=�V�fm��-\]�˦�7d;נ�q}7Mۑ`6J3�+أ�m�Or�f�Nv���~�)�g!�U�ro�
�!�C��b���T��ǯ����m,���02������tպ3�dS'����ZMq|~c/	��̂t;��Q2���d����H"�#��~�Y�2Y���T�s+Nq7WY7}��b�͒ˁ��{�j������ךFE� ����3e�ݝ�W��Ri
����?S5�NE{C`S6���k���(���m�8��h]s7ދ�^x���VP9K?$:��f0=*�8}���|K�fi�<��%BK�2���%SZj����Gۿ]-�gvxt�Y�����1�tc�V%�
�I5%ՠ�R��6�!<4�<B:�LJ��8>O6r�yӱ4���9��o�:��Ü�js4��Ѫʓ�wIe
����ˑ���΅=���`>�o�X���p*k��>tTl'|�aV�C���*DMeܩ��#ztvmh7��F�1�r��}o��`X&�S��N�����W�a�)�i;�����&U3���DeB��ӏ�\��m�!�ְJBۧ������}h�@�s����֙'���g�O6�mv��w�]���������Y/;�)Ҋh��x��d��ܨ}�P2Tb��̼+�G6�k��rʼ���v��ꮮr�Q�����l�Cʯ(��-��O	��mvNѷÃ���?5F�E�s�����$�e�c�#xv�	���AS�w�Pj��_^�ݜY��c�b��m��ܴ)�yj��!7���V�:K� ˋ�([v�|��-Ζe1DM���-���\�u�>�\U�X;.�B��%܍@���>��&#�{�)�n\ql���Pa5�m�`��}�?[>U6:Ci�i�/��u���V�`��o	�%@��~1�Q��n�q#]�5�N�Q�����u]�m*碙��eъa��*p�ҶrDt�MK��STEJ��)ַ����K��^3��;o��c�^p��{
�晃��1;6��0�֦�uk�V.�S�)���0-��K$�W�l�)�_w1u�'`�r�Y9|�w�N��픱�8+�X<�����S'0u=l���Y*i؃H�1t��~�����)��bP�Q���~Q8��vS����R�C�9���t�d�Y�vТ3c{m�tE��7��������v�Py�������
WK�l�g��;�\�0�JnI���}��Kc7J��.���E�>U���\a9	�Dc�f\���d��h�e�)�zNS�����Q��M�Q������c�m�l��c,v�c�
lQ��N�Mu�=��g���[fއ�؝���Su=��� ��!G6��`���g��]0�h�et�s���N
���Ͳ���`�����o�Դ� �޴r��ƪZ7d���_8��X�/��7;^Cik��_��z�g�Oz!{�_6G7���3ϕ{��4T��n��'�K��`�r�2Bm�8�[HO�І^0}l���؎�e�b
�Y�
؄�^G��[gB���4St�W���A���*����bݝ�J�T��Sۍ�w�J���
��8�&%�ow�-��Z+�l�`�0��PWRk"r�nR�1{�B�)w�)�T����w��!�q	��!!תm�hD[�-~���sU^�
u�K�S�ڈn��/x�-T�B�j	�"�����*�թ��K���=�<��R�)������Q��?*ބ[���5:�G�2�`9.Xv�V�W���,c���m�i��ܦ���ި�=�Iݏ9��31܇N��9
�L����T�}�d��U�o:Ɏ��M*�7B�u��{ �t`��Ne�����r�&�L8���a4��nOh�c��=L��n�`�J+":ۙ�����lX��O����0���a�F��ޢ��($�%¾��>�R�>��0}�ɣ.ϗ6#�V[�l�Ԏ9����s�f[<1@��-�o�_�l�
��m���U2�=3q��Ϛ�^�	?\��FUm���V�s4܇��C0[0
���d�����仕�.�e�ʙ!�WB�3h����q��x3��t�o2C��������m�'��OL��vT5������	�Qۧf�I��g�~�w�m��y�U��{%[�>��E�����}���OxgB�ɩ9�]�ssZ�q�L�K�[!������pSt����nی��o'�V�k�S���a7B�~��e��F��ߚ��'��0��dvIuS�n%�ͫ�cFHX�eCo�Yu�3�8�Dh��ΥTnj�I1ڇh�6+g��=F�����m�)�͝�P���׏dƉ�0YC+���?.*Nyu;J�4~b�7�lʺ������HQ��q�����]�N5��Q��gnh��%ū�D�e�4~�{��)����=�av:;I祎
徾�Xŉ����zRTӤ��F��Q��(,Fh��a� �.	]7f�mN�f�n�{�
��d��-r%%=zP��-��iʬ���z<l �6�c>��Dh2i`�__�_c!۾�k,*��ul�����X �ZX��s(N��5�� :�a��c�'��y{���x�Oy�������0q%��&������:b!�*2s{�J�]_['2kOP�Ug1�ݐh]�U�Ŵ��wP�v�\[��_öj�ofY�b�E�xXh���k��}�nXh-]���"�&F�F2nP�I��[@�.��һ}O,��.]P��a���$�`ԯ�ш�_2����&��l�-��嘷"�L�C�]�l�Ҙ�����4"o3z�ŝ��� �3F��ٴ�-n��Ã�6�]%ޚ��dE4ք��D�L� f���z6�t#����S6VZޟu0�i�V&�&9&l�S��v�j&c�S��ZA0F�'��K����2�r#�ۜ��V�(M�	3b&�ؽ��d��%t���<^�.�:�_��,��oJm���re>��o@���}k�Ve�\ԧ��3��ѫkH�;jط�����6{2��R���;��%�8�x�D���99����N�S+4_e�\�{	�yJ�ὒ�z�R��v�#��hB�	��SLe?Tc��PJǗ�0�i�è�=l ؓ1�̦�b��2��<k0�S�T�u�W�E����K��h���
=�z;4DBm�#e�w�^�x+�=�(ҏeMu��E_],�����]�Sp�&X]�V9��J��&2�@� ��W&�7p!�)�m��߱wvs>�W�Ķ�{��mE+q;Ԯ�A��XΉ��A]V7��׻t0#�][�ۤ�����a���s����!�.���!�J��Ζ�KN$�Rp�Z�3��К�qK�Й��(�3HS��I�&!o��>���(;`�5|8��Z��k�qe`��P����e�8⎕�t#����KLoc�y��>W��fWY�,�1⎇|��z����)X�,�.a�S�oV;��e��#��q1]p�1ɉIr�
�B�+�ܭC{i#.����k�5����*�3��,�ڳD�]\"B�� ��Ep�J�-�� �Υ׷j�K�@��wM�NYC����{�V�w_���jTdը��+�=�7Rqɮ���,%}���
E�Sf�4���:��oQ�VIv%�b /�E�81����᠜OH�b�;W�F}O�#M�3�!��w��a����tv�K�Yz����H@�$�B�)�J'T�ʚH\�jh!uW�."���I!˜�Ajr��
��W����p�(��U,(�<�ʅ2��{�8"�
�s��AW,�ׂ�N<{@�QʎA]��yhEUAI%EQUӞ�#�S���DQ�xB�wREs4�I#ZT��9Y��;(�LuӅ;9��TW(�(9Ar/hW
)JCRԊ8D*��*T{H�UZ$E�T����J*����3���B�{�qt��TQG#ŤQQ����G9r8TE�pr%AG�*�#$8�OW����\�r��S
�(���q)'"���A�
�EVHt�Q9G*��F�
��"�q�9�9U-"*��S������8�ʨ�(�-�(��UAv8�T���UÅ$�%p��
��v'/"ʻ�$���r��s��B��s�2""�(����ʸjG.A �I�X���bУ6�b>˻��_�(��bܰJtԮJX�Z�]Ã�0�kfv�S�"L�;M۽���;�@c�I.�m ṛ'6 ��o?6�Su\q�����½���}z��k
��gY���
(�ea�"����{���=���n�7T��6.-��|���
�q�Պ�����[<�R����r���a�m^
�y˻�ӷ��6�f�B�B��'�w�j�����(а%3��|=�*LC驩�8s��[�9�o��wb���#�nv���R
*g]�4�yj�(X	�\�� v�vb��k�C�H��H��=X��^k��T+���
�o�_�)�Bw[q-l�;��JUi��%�_�+nNN�c�h��l#���M$�fZ��v�h>:����r���҉n�.�����9��;���{,�m������r���	��Y-[�ʚQ"�t5n׌yn�U.�#�,l|l�2�ah�5q��%�کn���B�/?�n��Y����n�*F��4�vQ�yyc��V��6p�;��j.�F��B�0�Y^��"To{[8Os�:�l�cm�xd5����Rá������1���e�O���pX"3zn���p��g$g��n����̺N�x�iݜ�=3q�b˫/*1A�L�H�֥9u���x���+8�|.5�ìH&�S�+7�Lf�&?f�4���h�~�3G�� V�� ���)+�mZ�����,��/r��*45��pu�K_]B@o	�>F@��&1}��ʶ�n>	%v��x;���m���Vͧ��8�oD���;=O�1�c�OL�,z�)�����,��s*�����M�?X��gٷ癍��W��c<��헂�d!Et��Q2���FK��x�'�y����	= 9�S�ay��D�&�k����t�d��&�y��A�O8�i��2�:���?V	��q6(R��^[��l]��(<��Q�u���5q��^���3߫OSu�!�ޛ;�hλ�����q������7���z���ƽ���޸���󂽊:+��O��g�3���<��(~��ϏMYs��S�hsaΦ�����c�辘0�'���	�����f���(�1<��1<�N,�������O5F:��Z��������R�� ��v	����!X�;�cU�l;��qX+(\V%����O���v�r�Cq����+��B��๦[/*
r�bZ��F��'�Q�uv;�E-q̩�`�����PɆ)��6�Q���\�<�j!��<�WxUWrJg#Ĝ[�ȸ��z��n��Y�qPlC���TϪI����EG_W<{������k�@���*˳?<Q�t�HW���B<�L��㔆޳F�}n��7�y�����eF4�d�P[V/�@�F��%�L�]���'��+��۱�/FGRb�5���u�*�kx����� С{�7[�2��C�{f����Ρ�a������3��6 [��"������}"��
]�ߦa�(N��Bm��f���K� ݐ2sE�WI5�'��^d���2��9��S�`',-�M�Нm��ܴA�l[��G9���u�΋h���Y���"��B
;ݰUv]�<��QLo�G!^l���nf�h����xӱ9�3�>:��"&��&�_{�z��b`-�K�۹����S<�a҉�Exi�����n�j�;����k�G6�F�1�%<sϒ٤�w�*'��.�wW]2�e�~5r���v׶ng؎��t��9!�iN@��#}�`0ᕵ���w�B~�C���q� ;L��ϳ5[�ն��큳§���^N?U�p��O�"[~32��̎��b摡Sg`Y��j���*�l�-7��LP����t�`���\f��ǜ��#rS�3���v�~�a^W�"Δ�����%W��.%�d�ڹ�h`�eX�=�=��ء�;Yd,!����hZny;��6h�rz�;�ޕ��omc��X�|nX�/��1�c\�=v�r�����x���(}[�N����!Jˮܹ�ES���W�d=�o����VեՇ"��.u��^�)������S.Y6���vT5r��vR5Ⱥ�c̺���n#�d5A�7�v�uw_S���v9��J�}���x]��0ٗ/��]ᤩ�9�Z��]��<zx]e�ᒿ7�.j�DZ�u����5��%�ż���\j�c����52�2=]��p[�����k�dAmc�3�7�7�;�!]	6+��pE=��i�w���eWT5�Ǡ��rۦ{��-�иf��$�5���r��N�5�6u{xӽ wW�3��1�<�q	���)�g�Dc�a]\�w�qS���/Ktw���������L �x�U
�R� = �w�0x)�Ngz���f;�6�s_A��}z�2�����������X�҂�Y���=�=�3B�S�Ѡ�ggfm*�FV�j������� �W���t�^�t�S+l���"����{*�Q�������]=��v���;��F�p-ѓ���]߯ٓ�,�eH~�V�ׂ񓰣x�K6��
�C��#nnC�J����fuC={�-�b�|:��w4�gK�]�7ٓYz`�w��;tE⛮}�fH~��8!�أ8m��{�/,���'S>;U5�[o���a�.�ƣ�/59[|�������40bx��s�u)�v�¦�=�BT��UG^($���<|$��$���VX9���)҄j����8q���nx��v�B��`9Bwj����̦j�w�7W�$�͕� 2�/���`ZMY�@du2��hS�J��^����V��/�������˼���H2-�c��h�e�s�5�>��1�fJ~Z�M��q�w�Uu��_h	�L���d��E����d���y���f�l�m5�`eMy=�����s�3��}���Vr�q�3��*Kװ̄�O��]2��`�z�h.�d�,�.��6��.�t�ufU�T�̹�}3���)��ڷ{3�|�9�A�s�]�k�]��A'����E�XS���9�A{���m��cp'|����>�T�4T��]M�S�M
;fN�K���W�Z:���t_NN87��-q8z�3��*�~�dz���Kh�xYr��g\��t�������C��l�+m2V	�'�ͻ�To�q�3\G�I��u�U>5�F�ޝ�����6z;AhVi��mG7��((��f��x���

��H�e]�/A�,-G��z���7������˶��n���"�WS+n��e��\K[:�::6̜g��9�8�5�r9ߴ�!NCq�%�9RHZ�an��,˫���� �t�Ƴ
�}~�V��Kc�j�n�r�7�q�5�E�(U�xt���������'��W�X�t}�;x���X����A�S��2%S�]��6�XUl�`���)d���V,�1Q�r�-�S �d�gm�x;���zUa�t����	�����7��8�<�Bк�Y5�,�RA3tF��s=?uWU:�ǝ}b���31yg����!�w�i�}�S�]���߲	jݖU�;]��#44!9��Y�p]��mu�-|\�n��̩��G!M��]lEos��pe�Or�ӯѭZ���dCN"�9
��q�����Se�5��!�-ڲp��g$Sb�}��:�'�6$#m�z�Z&����-�TOQ��b�Lc�W�x{����2�*Ye�Xe.ێ�ʚQ0�+p��٧g�9�g���X��yl3#�3����T�>���.�L=�rj�[����y���:�Z�;_dvnK���Z��˄��O={�A�O8�K�q��Ɋ�U�=�.�.�c��wT���fC�U�NE`O�L��zoOcv2|鳔�:��ҵ�s��s{M�h�=�)�yH�t
�=)�'����P��M�;�L�&��[v,��'q��T̍���sFRѭ����n�c�e=Ϯ'z���X��妕J��/�6Wi7�����IX��dH��֝�*�4f໻�$�N85�*�]��W��9d�!�Ӡ�J�0���ú))�jA%��ԣS!�P+82��7V/���C|�:�;���qj6w�:T�-�S��)1�`Ԏ�����r��착uΡ�@=0���Q�ڎ�%+J�e=���[?���w>j�¸�Ό}�ʋ��mAMk�/�3 1�2�Ju��W��D�sv�{�:l�쪎�q�f�k��v�S�ny����R^�v���Ze
�J؞��ک�U�l�A=��ީK*p��\Bs��\�mQ�7�q_\9zefS�؄2{_g�V�8�k_�s_!�e1��~�B����mQ�EX�:*s��[3�$W�@���Y�k�u���'$���Ǯ��B����tw[~����)�Y�
��d'5�����H5]�C���w�Gv�4U�GQ��G��Y]*el����0Ǆ�d4[� �6-������]�Sq�4:�a�*��! �����쁀�˦���QLo�G!Y��̀�Ҷ{�sg[.���`��7��,�'8���x��c�=yN�!j2y��.�wUٖ���碙頴�)�@~�Y�д@eAWd��G32�fC�w�6L���n�n���y�Q�@�].�w:��N����tnOc���1y�������!���Uni�m7��t�	���)�B�&^N�@��~�T����ܴ��:�b2�w&�@���|�rG}حMż�U#'f�M����x�sү�+�!c��yј��&͗M��(����+���؛4f)2��W�u
.��+8ޗ9^.Z��Ne�����G�����~�7�$��7J׆O�KY��X�0���~t��Y��t0�"����\���+|%��9�L��3q�B[��X/鏸m��ϴ���cŌf�8�l��#����q��ڹ��l�_���+g��(�gD���PCV�<n
n�ez2Y]5�hOx"�_&�to�����9ټ�Oy��w�ٮ��U�;�)�ڷǵ۵�j�73t��M��+P�?kI�8�NE�gh�F��sͽ�Rhb�۳ϔת�抛��}>=�_^���K�̐���
���ad�F�������{ �M���S�>���;Ҭw���*[8Kwv+��Uê������$JJɈ��z�.T�J�E�81�lսL�� �k�A�e��n�\C�ÝkkS5�ޅF���:6��--��oݲ�(W��w[m3n��C�G���!!תm��Pd����a�Q̽$b��
H����к[���Pc��H��.�\�=�D$嚌
l�Nwz'Du�ت{���qB}}(�~n/��Η|����@��:0�#Z�V�Z�_Rj��XŽ[���/iA�^�$��j��<�Op�`s�evu7�oX6r׵d���"У�aK��u;[�~�nz����g%�>���E��X����o�e,�u��2u���ޚX�8
z�;,N"�<�/U�}�ٌK�q��m��vo>�Y'F>��u�Kq��	�OI"��d�V�z���ON>���������<+G���[޾�#���_����<$Ыߋ���eJv���FN�6����veC�M�K؄��c�
�"��)�ː��<6�nCǥF��u��h
Ķo<�S-�B�<:�/���:�]�'o��{{)�X�ʉ^0����9p�������m�{�/,��&�u����m����l7z�K�e1��H\��랐d]LqqR�*�0*k�}�8�B���y���Sݼ�s*Q��<�y��~���q�'�]u�����@�;-�L�9��E�9He &^GgI�k�����9���''��g����A�O��e�y�`�z��@�u� ���{p�������Ͳ9�yKu^L��b���ތ�w�'�8=�oRpE���qn���ݼ�s�����tn�nӎP�*�Z����=�:�<�P��>��B,�l�%󳟔
���*r�F�Ql��˘#��$>辜�pne>M��T��X�ʊ��L�[=Ou�#�m�͗�kŢ�:����6OTRԃ�)r�&fs<�zMQw��]w��> n'�e-V���{cu7	N�$d).�Z��yh���n	��0�>���Ю�������Rq���㹭p鰶>n���n�uvW�<o�z���f�p+0�V�����#��8o��Fݳ�R��
.-�ٛw�5F�O`bqBÜ$���Ӻ�8�{Ev��a��ٹG!�а[-e�����s̠�R
%n������td�؃߯G�?$��:���^�XO^���ݯF���ЪK�saKb�i���֒��T�f�2ie��>�p��ۙ.�[���K"'/��Y
R�<�����<����cr`����Dí���{��8_9�㽱�����3�5B��~l�DV�2�h]D���&�x���� mawuۗ�Z�t���
���j��q��9�xջ,�J7�;��(
���1�~&�`�F`_L�b�sţ�VCAu�3`CJ����gO]z���yc;'f���5���aI��Qr�#�[9�e�M�'�;����7Mۑ`64�9!�O0m+�vk2M��O���-{4zb�P����!���2���C?z��*Yc��u^��������}H4�����p)���ǖ2�[��Et��/�/̣%�O[�8�mQqalڗ��ho������ן��x�_��yF�6�hCS�b39v3o�A�ӑ����ne���Q�+T��ӡ�o�g=�V�}%��U�Xyu>d�����%{�}7�������{Qpǭ�K�a:��6e�2��],Y\ɹ����3��1�*;��i�H�Лh��ߖj��;7AO�vw���\���n\@��}gV��ںz�&�I&�3�/K���U=ܝ�(cz��ne�9����G�Vͭ*�Ы
��!��vO*��BK��:r��̲/y�ғ�I<��q<���7w.�2 yRv`{S�Kz�j�u3�xP�����Њ�1>�u�^ѮR�&�t��ͪ1�lbr��͎o92�;1v���)�3z�,m:2����7��:ŉ��`�@����]����B%V�^ jc�g]{�9µ_+i�2�B����7������B�+�jJ��#;�
�����OV�@A�-����J%��j��W'_R�����BM�Zz���V2v����/ ؠb��v%ɻ^7C�৕�1]7O�E�j�_,}W���v�ƅݲF<�A�A�y�_�gGm;�E��{�%u5'.��t�+�V:��Y혴²,Z�����a=�U)Wiv�mL�1�꼥��ufm�xM�wpnӇ�R�Ę�5���%��A�7n�:�)g��~�MU��y	��vy/7W]�FJ�Q���&��Q������{���5�`�nvJ��f��3�[�v��ä�Y���VͰ��I�yu@�MD���Q��Q �L6撲_�l�+5Ӄޫ7#DrĒѳ���҅�M�zo+XhE"�h:�/o��6��oo':�:Qd��1�W�S����X�M5Z�v<�"hYqE7H��p�Xy��4M��o�f�KY���/l\��yY���.�Aʓ���z�O����	kGFe�\�4�wU��u�ZS�9`_5����7��!*B��k���*~ž���-L�CEB����!�^dW�3�2doe�S��{\M��0��7�i8��>�m=昛t6bLގ=�h���M,N_k��γYE'S{�y�p���Ա4+P��݁Ֆ�
�V�����c�h�oB�k��)���IL2�x5̫�.��y�	��Ӆ�,�he�gr]�;w% �*�R��Jت��t/�p(�ᆃ�.��Z�ݬ�QV�{���C�bD�L���7��b���]k�}�w�A*�������6jknʃ�f�gJ�)��+����4�WC]�vf��o�Ebe�d�!�t=X�l���A��e�RbQ�0Ven��-7�PjFQbZ7�@�ʗ�^�.Y@u���@��d+4m�;y�ܫ�1ǋ�qڧ)I�rZ(�l��e�ٵ�X��:�5)ݔ[�z�,�:ӑuZ��"�t���	ԾM47x�٧��^U�bc+�yL0bjEWn�Y�p��u���v�6q�Օ�,*ӕ+U��q2UN�m�1VS��6z���W��-�;v�����]�H ����at�(�#�Q�B#�9DG*��㴜�L�����B ���	Dr��TQʮB��¸\;��H��R�9^0��Q���QU�.UȔ.��PE^��n�*��
�.\��,���9�r*�����Z�K�ʪ��ZEDP(�E�*�r�UTr���NUDADDS.w+(�D\<�H($�DQ�dAAr�\�r)Ɛ�r�rg*dTDDEȪ��2��6s�.W(�#��I$Q�eQʮ�GeTPQTI�s�ÑEUPZ%�;�)�$^� 5*��\�JQ*�����QTQAs�p�ЉRDJ�Tr=t�A*.QQ\�QQAAT�@�TA^�+�TPP^4�r=HA\��U�*"��UT���^$�
��xB�Ш��a��"#����.r�"�U{�I DAQ	"	���#=�ezS�n�X�p�6[HNNcV�F&�E
���=�.\#�y7Ve)ӢH������ˉ���t�4e��;�M�������uc��cy:� ��-F�왘A����%�Z�y/ƞ�N6�7�1m~��֘C-�-�FG=�YQs����#[Bw�=M��D�x��ٍ!R�~�u��ek�k�sZ̦�]�(�q��M����=���X�?^ ��-������^J�W |6Y�
E�����(g�ӄV��l]�$5�+x���6�)�n'z���=9CQ���՛�i�՛����즽�wyj<�����e�E�{&bְJB�c0s-�6uc)ȁU,Mq��`-z`�N{`:|�dz��)�7_T9�we'׾/��ɀK>�h��h��o[[Y��^��t�Tw�[�n�P�����eL���[v������[%�9~�~-|WL;)���2u�E��{;��tJw["��R�yf�⢬C�۽�Ӫ	�`p:
<}���I�9�mN��ۂ�c���=������ן�uQr��NK5l�V9��2�L�#��H}��΃3;l5��9�``��L���zB{�d4[��b�(<.����f����KL�Q���ɜ��������v�U��G.<Ѭ�}t{ٱ�P
#:nR�������������T��쏟�����v�'���O�7'g��+0Q6���b��|z$OZޱ������s���!W�4�;��Tg:�������ڤ��2x'LݐB���n˶�y�%�OCO!a��ȍ��2{D+~�֜��R��;�i��]I���L�f��<ஜwE�2�\tK>4t`J��m3F�kZ�g�o�%�_�~��+g��uLr���Ğx�Kf�[.�P�ws>\��6�ō5��f�	�Η~�l���N�2�?o�� K`X:E6��L�2�=B�]��oI݊����f��i�/��2]��ʐ��9���|��u���x��O�#?a��G�_W5SsC�D�=T��-`0�k�F�Ī���(}�t����4���Y���X�_�R<�q#�8*�s���i��{��u��N�"���t�ئΉq=�PCW���pSt�#)�%���hOm	�2I���S�f�Y&{P�6�;���|�5�ޘ���{m�Z�mc�׳�N=7,y���7�G��>L��b͈9�P9�z[���hSb�|T�0��L����'�8�w������/��P�|�R�ͺ����B�38�\�|��Tʮ#:)�s9B�b�#��/:��ׁ{��T���W�O3d��mҲ��\��[Q`�&;��gh|i���<
FH PB�k��F��ܤ7�2�jG�;��49j�Z(�k��ږ4ө��"w�4c���f�zY������i���ꃪ�)�9�&v�b�tc�=��=s[*g>O����a��yT̢mӃs6�[�ʽqCS5�q��Z��pݭR%����4Z�����	�e7�A[v˼��C�͙�xi�!��Bz��$8��.<uSvČSC	۵/]��<1ֺ��Ytv�f�}M��90�m�iT+�
]�ߚf���B�â�_^�]]u³�բ��g]e����/���;�q���%�뭓����BB��	�l6SO4���'�5��م�6�h;�vK#Q��)�$[.�.�S�����K�2��F^���-�T���lns�:����"�Df_�p��M2��k�Sr�pi���wA�̙T�B�������ܬ��9	�0�Y��<4��n�~`�m��d��	�N;��ӾOrx3U�I}%�-{g%ܮ�w�Ws����6ۦ�o2C������Y<�l�=��N�P�*�����x��׆�\5���&~O�.��:�U1�h�e�yX�9�t킸��0k�����V0����9�K�� �u,J�q�xC�jL�;��pSt��Ѳݵ�k�T�T@�5ۦ૵{�j��hR���AJ��E��7q���/���	���x���3�oa�]�
{|A]�O����u���=R�K�0j}������Y��A�M�oV�R�7��0k�,RV�r�n��9�L�Ilw��:�x�P�0�"vٹ+F-��9�ա��̭ڣ\FBw{��O>���)�5yt��
�/�ͫ�cFT�~ׅ=N��4R���ܛ;��"�Х��5��ȋ��ca;��R�I��{ҜYٕ	'0'�u\���.��6��_�Ʉ6��/�b�.�:����a��E����`*��w���9��~����im-ٷ�ĞkC�'�[E���Z�1��872�'��U�gCW�C���ƛ���/2ƪ��M����~�9�Pƥ��v*m��!`����s6�Q����GG��j��!�p�푼bb.�ܣ�ˮ��l�f]C�m�z�.��u��^��Yy;���6��1< ;��ctX�-��'}]6��׎#o˧�i�]OlM���1��x��"�^�m�w���ü����dEvC-g*I䈞tv1��uus����k��b�gy�/z(oy����	߶/�!�a*g�����Y-[�ʚQ"�t5
4���z��E�ڼ��[%���YR�ǦT���CACm�!�Z�����y��L�^�9zҔo0�2ӈ��gyĿuŶ	��2���r����̞n,��7��!B�U��
��.�N�n�v
���{GW�d�;yqH��zx��@�xf�ʶ��'�����.�pv�Q�C��Ɉ��k�<t�}"[Gf�'֏B���^n�p��Ď�Dg��@��*q�\ʐ�Mɣ�����b(���A���9: -�[�mB��7b%5bF�pw������je=���iv[CJ����Z~�F�D��Oߣb��̾l~��/��s�/�G3j����	�|b@�'���e/�-Lc�W�]3����S=3A�#jq��#n��Fu؃x�Ol���S�'`���ǟQ����fG
e���L�e��x���7GKm�S�ݸλ0a��`���:�\��k̖�����m@�l�\%�T��>�q�s%���:6�fJ�U�|�C&(Q�E����3FB{��u5s:)�'��N��}��Pa�n%��D|����y�!ߙ����岙vT`���n��2Z���`69��b�ΌdYn3�c��yzh�v�Od�;�f�g&:�3����;:�3�a��[�`����d����c(�Օ;5�՗�b�n#=Q��ͳr�{I���"0���.�/��dԐ��u����M<J{�4l��,�ٵ%�#�ʭ�t�^G��^r�Cq���[��|u� ��q��Ku�����)� V~I�OF9Vj7zv����%�6�q�ۄb��(�V'm3%��@�I��;�Lwe�wK��o(���[��rK��=|Fr�u�1��)����	3qm�jv����۔6�bǂ=Yo;��yt�t>��	Ϲj�����I׿�^~���42��Nu1�F��#��T�Nj��|��I��D����{l�WrL� X���֡���wJ.E�Ǥ�<4������t��}R]�wᬳҹ�E嬞�$j7F�ptu�s��W�C�B����i�{��)�j�W���0�%��'��W��w�I�1�����_[vy�z���E��d@}�DŶ�N�46z�����ジ�t�c�\5��_l�n�������4rY���+y���w�r�7;3�۶�M�,��g�&7CI��B�T�s���7*`��]QL�ݴy��֬候4���Y�u���|�[o+g�p�`ʆ6��<�[4���~6�Q8��M�������6���.d�w���w
���M?>_�2C��t�	����+�/����CGNI��7�/��a:g��v�][��u��ĉ�}�b�Y����\w��X	�����scC��&��y�	��@0��H�^]3�ֆL<���V/鏐ۍ��kד�Oo�����k/�����zm��Ĉs��]N�����e�<a�0)7��YT�W{z��8�?oV�JW)��9Bh�L�T,�|���#��}0�ي5�ӥ�,��Q�j�)B]�+OS奡*�������c*���j�dLb�t8X	M��S�ͮ�wx����9�̮��=��	�Q�O�:Yˢ\K.���W0��u�e|�NX�?:�V����?_D����S�Q�Aމ�w�ޔ泲���X�|nX������C�BȞ�¬�@1�ީ�l����a�l�>O�U;�VY�ηN9��T]��1���&�����GS�9 ���|-�B|���SQ�V>�[ϔ�W=z�����B����c:��ů�P�Xk^�l��L�mӃs6�[�ʚ�i���-��rs6���3#j{��;.	�tƊ7��LǍB��.�)��b)��cHyj�!?Q�b������2lXI\Ʃ�<㐷�2������*�)��l�riT)����L�μ�6�?5�N��q��$�l�~m0HSy<�Z�q�Yh��׎#o:]�Yuu�=�8%�z�91}��US��,����5��7�3o>�3�Mc���dK�Bp���*��|yn�5/����810��2jfZ-W�9�8}�q����<E�FSd2�'vYR���mѓ��(����i�8׈[�+����^�i�a��hw��R���۴�W�딧��w���$��6�pz�׮�w�'����,]+�Sj���:ʘ,-k�1p1f��*gB9���VTg@���ݹ�7�35���oW^A�5��6]k�򱙸�|^�[�ܝ7�Z���[��!H|d��'��h/�`=I���p���ކ�ǫ�//���
�C��_u��d���w��iWs��K�#z*y�}�!�m�y��bN�1F{�n�zڍ�k��Æ�ݕA��t��)�g��r�zzzi����;^f�kc³�ɠә��ċ?�,ӽO�;�5�Kd�R�$��_���t���/sGi�����lSt���Qm�����OJj��9�;�9a��'�V��9-��=<��d ��x]��ǰM:�\�-j[����;�y$÷����!��_C)j��apء�]�l�SW�E�|�<�LT=*�.��*2��V)6��_��f�U�4ۯ6Gq���y+��B]�g��.�5��3����4�')�>Wգ~ޖ�)�f�E6vTh�nY!�E�ž�O�q8z�3��A6jR���t�o�s����ϥS=2�(of��%�-۹#D����	hȷ�[ho��x���sA��C��;w��I:�4��lC������ܧ���t�Q���(VO������{TD5��n�khx�_��7�kj��T�U	���.�����f��No7��� +��)Ds�&�ukZ�qu�s��N�
T�qe,�U�:�˛8�)b�
���W�L�F���uFW>�U�rÇc�
˝���
�}f�i9r�7\����v��mY��c44������eXOCWV>�#W���%����˦ۮr*�X��'#M{wvf������ �Zut4��z@�G!���,�ʒE�x�;}���H���M�V�)�5��k�FH!S`���� p�	�|�<;�%�հ�Y.�Fۃ����w8R:xP�٩�^�WSW��@P��$2�!�Y�;E3����E�WZ;�m�J<�N1*U�ChU�/�{'�����\{.����T��Ð>�h.���<��-�S���5�����$�������.�#eCW��)tc��]��,�&�C�gDf��~��s�<#�3��fթ����~ 7{tɑY�tm���m�ybzi:�)�w��L�>=}�ډ��"���.����T�e5�;*��c�t׶S�ɗ��ޑ�Yt;�҉�\0Uw��cQVӻ�h�,R[;�Y�EtAs��)�
��e^��y��Dܲ�;U)�̎˶Z�qAu��z�QT[	l�p�Y���{����� ��t�	��n�\l[�ϰ'|o6����<[���:l���s�9&`������@��X�d�^�5>���W�d*���f�5�	�� NHhK�갴<�s( _	P�־*�Y�%�uWD�黺�\�n��_C��m^�։��`p��`[���/ss��Q�:�M8����2vN���S����O)u�\j,V�8��^�FKT��q�\s�	�t�Z�c)��V,��rc���zޖ{be_C=���M��M͝�ܩ�,gL����Z�Be��v���٪�hi#4sb�|�ه코���T���|Q�Z��gHj��S�`[M95�L�\O+�5�`o3L��jc�.#��(���O��=]���p��k�n���k��J�˫]�+��R�DE��{��G@�A�K�4�S��G9�[T2��=b���x#:��8�.��e�s[D�.��oi��Ɏk�<�Q)�l\�w�2���1^��#;��X�-X��� C�uG4��o�+�`�m�R�wۈ"�;�7B�u��{�R���!�$>�W5��0d��6�������4�u$ٸ���ݐ,J�Tʯç�'���5�o�a����� ���5:r^�t����2�d6ǧ'�5K�|�2�E�d[�)��*)�ۃG?7�m�!�i�B⪺g)����S7*w��n��9�yV��N�/q��ߍ������w���8�� c����ٱ�cm����1�����cm�6����1��Sc���F�1���61�m����1��鱌cm��c�����6��6ѱ�cm�61�m����1��a��cm��c���M�co�lc����1��lc���d�Me�t��ef A@��̟\�$o�7�B����Ƣ���E��H$٤!Tj�P�����T�4j�*����k!F�Z�UJ�	J�MkmP���T�*��l��Kݮ֛R��ȵ�Vmlj��iY&������E�Vc2im����[4֍Z����U�ڴ��-mZ�fY�jƭ�6�m��6��q���e@{s�ٱؙ���մ5�3,�[Yk{��lŬ���5J֥FSk5��T�Ыmf�f������2[S3#}�;mKm�kaf���@�f��X������ִ-��  �}����Bê�z���=몵�ot�C��kX�h�� oO3ίg](����z6��=�����n�Ǒu
���e�1�U�m4�  ��}����V�����WyP��G�r�Ǣ�����C��(�(��/=�Q@QEE����QEQE�{Ǣ�(���u��$P(�J�:޼QEQE���R�-���k(V��j��C/   �� kA}��<ֵ�F<��z�@:�պ�4�ի� 4:�v��F�� :k3�(=�({�Uwo;[Ze���&��ʲ��l�W�  ��l��9m�^7�D�γ]1�ǻ{u7a���=�ݻm�K[y���=N[V����T���3��s�㎛j5��n�^�V�{j�s�����k������ֻu��T�J�mm65�XV���m�   >��lͭ�Ͻ�^�E�U�6��n�n�Eٻj�=o{m�j[tuyo{�w^���w^��t�Vڭ]�g�S�F�������:κ�� w��Z��w�m�uos�zӺK�*j�v�j�l���ش��   6yy}]v�+v����j�C���ڬμ�J�I�wk��ƶ�m��&���ݺ�n�O^��]*�����Q���զv˽�����mS�z���n��N���R%[�7�ڵM6XZmm���V��   �RQ���ܴ�ĺ�׶��v΁�ݸ�k���gN�wzoA驷s5m�^�m�iv�S��{��g���e����ݕ[t�����l��e�+׏m��8]m�٭�[�0ح�[,�گ�  �Z�O����ƛ���ղ��������mm�Z�U{�{lGRl�Ju=��p�oW/Z�j�R����؝�K�������������������+�Ъ�^�e���k+=��k[m"�V>   �����y�W{U�L�)ۖ�[n��:�kWs�۹Y�v��㷱Uv]8o���Mf�5��]��[vn�;���Զ�I�gGۮ��e�����5�n�m5���AQd��vZ�l�  ���(5m�[�z뛷��I����m���M��r{n^�ʵ�w^�{^Zݫ\�s�/y�:Z����x
�����KnD�����Q�;K�����S��)PA���a%)P� E?S�U*I�� )� ���i��T�I����#@i"&ʩ5F '����?�����eg��g��_����oY��eOt�����ߥ��������$�(B���BC�@�$��	!I�HID$ ��O�o���e�s�{��c�+q���e5��kEm�V���܈�`�ʖ�i�x�Ʌ�{p��ąSNz����4�-����u/G��G�7m����6��6;���q�$���1H1������K7qT�zk	�n%�q�Ʒ^��wY�6U�b�(�op�,*���v��۱U-�Œ��55��U!8�j�%їV���:p��?��um�)\�=ڷ��w�m�N
yqYp�4髵d��
�ժ¢#g�� q�Tr]t�h��	�d?��
j�]�יf�m8\�����*]��f
ܷ3[��'�,�{�١���ו[�0\�-a�G�j
j�v�)�	�N��*ׁkc[n�4`7P�֖Q��k�L+T6�A���)+B��5����o0����V�H0V���)ntɏpG��j:�B�A��@GtA8wT5�ѫc#�K�k+p=[cH��/^"1���fR�h�ZeWJ⛢V��
�-�20�k2��ցSc!\��D�^�GY����Xif��Q����V`�(cr����!S�r��$��"��%��*��l%t���F[�:ְi9YY�v
��.��y-T���5Ci��c���b�[&ӭ3Zz�ד^�X���U,�M��U6��b]F����bS��LS�B��^fP8�4���ڀ�fʏj�J-���i;����ЃY���q�7�ٔK�ط�=�0,� �ӊ؉h~�A���VkC�Y8�[M�o�V���V�hXU��e�3^qǁ�U��$4�ƚ��`-ZҨ[Zɐ1�l՜�z����y[�J�4#����M 2j�K��)���1ʗ��6K�Q�Ț8n��k�^�:��۲"=��l�dw�j�K����w�B��kU��O
dST������Tv/5 �n��řa҅ؔ���Dd��[T�`�Yo�F(I�8iIw�^� �u$���?��Q�j9��SY��Zz ��%pf��)��r�VY�z
�q+�J��4�����#%����,��3Hݣ(��fjSQf�2�H2���T��x]e�+m h���F9�۬2�v2�6��W/
�^f�1�2�)қ��uѺ��.��
o$H�Dk"`,���!'���>��n��<ʧ�2�H�8"	�v�I	���-տ��nZ
2^&��kt���)�sC�4���N�l��@E��{��n*�� ��*�r��{��ȊӦ�:��<4�x,��Ӳ"�s���W�o%j�� ���ڱz��ةF �$�=*�47�o�I���E��ь^1���N��,E\Qm\©lH��ne��î�P����I֦BOds^L��n��wGa�m��V��Zn�x�^���Q�*6.�hL�H��X��r�i3os%JFF�S(�&���M�K�8RIC�%���ˇko .58��1v�%��B��Gܸ9M��RKkZ7^k[z��F�jh�v�aXċ��y�ɲ�Ť�$�ݚ�����������M-x@���I��q���ˢt�:��ulbV�Q��4�N�!,֒j,pB�S����ű.n��@t�j�|���1���0��L!�u�d�(Q����-�U�Z�l֪m
���36<,�V�V	��[�9>�yb��N���΁{�B�9�#̌��ښ�k�(�VUKDmG�-��j��1�	�V%�oC���x�@��l�n\Ʋ�+(U�;܌�
�6�1���ouD,�+C��>%f�pHA��U�:7siS���Z�K�K3bE�$YWR�;�P��֨�BT�����b{���)eb�x�8��q�Io�H]��O��ʰm+P�g�k�h�u{4BBd�c�Y�������z���ʵ���i<Q���2fG�J�l�ִ��ڍM ;[6]
ɖ�8��4�V��A�h`+��ٛp̖�T��ی���{`�̥S�z(+R:oBuw�nYu�|��8�63ZM�7�����mi��	������D�uw��M�nZ���aa�N�Q[��X�4��̚�D3�X�M��x���c{���>C0H*���9�v���Ԫ�HGX��(��2���L��YoYk5���ېأ��tmS�&f+ҮEOT�q�V�7u�,SgM�����yXX�14��%�x��2��c��o �61a���8sj�۳u7+u��AUd���`�6��%�'~Ћ���[p���ȳT��,A����-�����4�gJ��R�Ǜ��`�D�C����t|<\-U�u�&����$��-}�ei�q��΍���&�ogJ|�l�eK�BV�Uݡ�(n�,],�f\ư���.(M�W��,� KX2�H,��{)Ź�+�"�셷��,)&�O7֭6�F����ݶD���د\ɉ7W,lIB���[k�T�L�"�n��iN�L2@Ē���kt�-�-�TΊv���u�����V;ϔ�CQ6kF���Te;��r�<��n�틣���`i��ߘp��X��G@p��� ���:±�:�� ����1�vw/��8Sa-W�P;S/u[ă�y����f�4���1찢dGO%S\�G� �
�j�l���w��QX��{R4T��� n���B�RRJ�v�X�Y���n�ߏy!&�_�&׻�g/�Hn��ݣN$%����c~�4��;b�ވI���ê	ڙy��r�� .�ff�ïHL��DV�)^ �j#6|mk�3��l��ö#��&�4�"�������04��#�7}���㵛�=[c`lV�ۋf쩠W�C�K4Zy��)a���Sf�T�6���cmdX�*�h& ų&�{.��2�d�wMmB���t%m�r�y/v5Fإz(0P��@u��gv*ZP�W,������	��ւdSh��c�KB��K���kYYs�9��q�o�-��������h��ԗz��޴�b��Ȭ��>j�]�jou7Lv�Kr�[n��;t�rKq4�E�cwt�Y��Wq��y�},���5���n���F�6�oM{F{�"#�5�o�
�lb�̢jf��ܹ��5z��GV�t�9��&�h'���(ٶn�Q��eݷ�[�&&ᫎ�f6�CB��#ow~!���Xܠ>b/+s7&�4ڴ�*�Y�.�������3*)I�N���S4����`!�:'w/qSu�4�)m��� J�&a�E-z�ĳ32ӶE-�K`��V�uT,X�6�ʶvP�5FS�,]�g#v��P�Dܺ!�vӆjwh��+)-�8�阮�I�L8��ݧ��8�2Z.Q�[�T�E_L�T/��f��[��[hfC���b�)�)HNF�b���E�75j'6�^cO|���a΂1�N@93�wIgщ�m���jWOP�&CK�VKr�e�k��B⹕��Ʉ�lhZ���[��	H��k/mJҲ]��)�@4����@��6�Ɋ���p�S�CtĭN��
��3Y�����7^F�!���d
7z�W&L4�I�7��ɤs:zH̶���chѱG��3"��F��N��Qf�j�I�"�Ō�v���;�����"�z�aB��x�%eMQ9�݃QA(�&���U�w�Ly��)wm8��A4+�5^(�n�����e	2ݺa�up�()�+mnJb��cm�O&Q5�f����C�mEY�:P�Iv����Ť<� �̔�1��%��7�bYT��	���e�T�f!)|6^��v �A|EMoQ����T�X�W9�&	X�%^�I��P��>�2�����*;r��3a�F���3+L���H�`ݫ�!;Z3��o䶃k ܕ���W�²��5��Y�Ii8���Mp8�����F�|���)b,�4�	F�۵�/`AkMM���ĳ��؎	�է����KA'/[�A:�QՂƐ\�t�%<{�euKr32���$�8�����K�5d�O#o�Jc�������5�8eH�=��<M]*CZ3bzV����k��Hf�ء�}�1��}����R.�4�t��k[���ٲ<!��ea�e4L�h�il˰���w,̗;{H3.C1뭫n^�*��wrS��a���+*+����!��tm�{��n�L�"�J�� XɦQ�aAe��'|B10���f�v��;ԭ�@c0Dˢ �r�53�r��h�C���dl�wW�Th��ܱ��"q����B�I�kYN��8;�Z]G����ed�2P�+aíc���7	@Ց���!�	��.�h��-i��"TMI��Mב3u��U��2��PVV]m* ⛱R�S&Lۗ���2,R,�˖.��&D�$!�<d�&1�����w�\��Ŵp��PK�S`��`�hi���w��#L�DZ��d�Z;1)3b�S~%�Q�Vc��T�+����a�ѹIV�w��7@D�P�zFZ�RWWq`�́4��{����J�1fRH�Ab�ݲ16�v/�I�B[d����zwTj��M�Q(P��=��܏3h�t�ܽ1�o�:���o���TYu2�I�Vlwb��hV�Օ4�*���0�7"L�A*�X��]�'T��X��cO���gb�!��#�	Q��T6�e�Fm�f!%��2�ƶU����3"wPX�z���F���`����	�J�� {��h��*�:RU��dϰ���k���=���z�Z�0��[��d�'���6tE6��2��3 yw��m�Aj�t	Č�$ރ�)�WD��m��kq�t(a
�c/���6e�N�^!,G��eC�R�8�Հ��v'�d*a���T4�e*��Y��i�"G"���v�9�j�	���0il���|M�,S�]Rn=�̫ ��a����W�m��-o��̤�R��.-�@�x�5I	�	��I�Yq5:��)ueX'~�`X,V[�3�Y�Y"������R*�´�.���Y.�+c,�(�3�3/qGq��y�HZW�tZ���RIHm�aR^:[�cT&��v��ld��l�j;h�w�e�6 �۲�X^j��5��[J16D7��.�	�j�����.
;��B��_ld4��֪b[�� ��9H�u�����M\*��Vj�����yu�z�A,���P]joq*	�n�6�ԍ)y����Y)2]ͼ��Ѽ_C��lR�f#������"dۧ�f�yR�ݠp�.T!e�ʊ�N��Y���VX��V(`�%� Ld�n3
FՙM��6�n�b���cb��*)���ٮ��Y7r�&մմh��J�+�^m0X�[��ˎDV���f�@���QnJᰱ��yJDb������+H���$%=�Bˤ��8��m�g����{�O�Z?0�[�Kx#"֪ӡ���[�ͭ,�'�1���x>_A/+D.<�n7pV&i Z���2ËmT�`+�XqԆ]L�`n��a�n�D��Q��C��Z.4%[���T:�qZmm%���z�V3����dn=� 4��C�q�AΓh�T��BT��4.��D,573m�9�Ƕ�bj^�����x�1���l]�5�s�Xt��{�Ғ���b�#�oI�d\��;FORP��r�x�#�XIe�Ř��I�6���53�V��.��.�������Q	b�t#[�멠ol�U���m�5�b�����u��-HSۊ݃��h�0�W��H�8��4T��3�^OTɈbG4 a�g�l+ $���y�W�I"�n�vE#W/.��R��{M4^*\,=��.�U���6���hL�h��eJ'J���G�ZĲ聅�\�{Em[��km-C�
�7>sh�.T3o�p�,MT��X�KkNFiͼ�H�X�����i�g��՚�n �a5���d�6J�eW�`%�hRe�H��P�Y��wfJ�C��t �E͹��%��Y��qõ��i�wi��nѭ���"���p2������k���YtnJ|4Wx���e\� x�
7[�����%�Ev�*�w�-�7��훭t�X�ݺ(���F�eAfkaЎ<U��q���eI�1t�6�2�mF��͔�m(��,��D�&�6E8Ub�-�fa#w���
m�:
[qѣ(��q��I�e;wa�b�B��aՂ�Ӑ))U��P٦��T`vv�����HX��*ݪM^
;I���Ͱ�*wr�
� ��e�j!%G�ݒ���.��C0��f6�#1�Vk-9#�y�쬰�L�4�� ǎ���2~(ej���G+&-B��40M4Z ޠt^���r�[�������LA{�ދ�	@V+t����P��*�R�nf�����F�3�A��[-�� �ª#�f��K"a㰓y8�7H�&��_7��������eZk^l���.nw����k����lb��U��Bh��0X�Ł�co+�7bЭ���e�"��n�sMe3m���N�<q�wt�^Zf�?�V�h@GV��.�z[`l\����f2#��^Vmצ�Xԍe�z�7��X��a�����Fș����N������+�ZỢ�fD��V�V��7�'
��U�4*YzN����v�\7pJ��+S C]�ؤXt�[������j'qd���'������UFк�R�up�\L�N�ݐ� ��Q�����%������A�]�ҥ�k��r^�pls�����Ȧ�=��<z�Ú��s���q@̅Z�����U���O�5,�����ǥ�o��b�QRfc�z�|�d�]�'[;z�i
������2�>�)Y��k�Ŏ�ܷ����8���mP��sg%�����^�vEX���}���W��.��#��l0OZ7����=����un��v��v�)��b��}�fǩ��>񾌜���լ��.�����.�����td�Rσ@�k���Q�	z4Ձ���]�u$�;b)�N����WF2^�����5C���gi�n�9ͷ3��]�WAN)� R����r�U7 ҮM���$�xl�h�a�)5��7ޟ	�ж7����.؊�5�.4Gn^t��j�Eo{�ԋ��|�4 \kVʱ���94�y�^��p������~�����8��L\x/�V����H�M����[G-WT/@y� ��}�W.����eF��F�Q$OM��@�"f��d܂��n�V-��]=�e�������k��	���]y1dC��U���T%�͊�MZ�D�:�9%�y�;�¼;5��=�z�A[rǲl�����1�7)MD��p�����ό�{b½��挝���GĜ�dξ�b3m�'�_W�����1��ƳE���LK�啩�S�z���,��rrX;�C�x睨��)M�yB��N�R�C�Ҹ�N�a	�v��cN�ې(�WB�v��g�sA���U�2���|'kCmUĖ�r�폜�+�0U���͂2���Z���G#H\:���yQ��W'�^,��=�f�=�'V������������OÞ#w qp�(��<�t�t.q����MF��l�wZ�q����4�,u�$̨��%&�K���;��p�[]u������F��cj�#��G���(� ���;P�����v����5s)��4_c7n˚DG�se�nw��[W�`[`����X(\Q�$��з �9�w�&D��d����uh��]�)�b�H�y}:�1 ꛯ�u"��ֆo45|)�Ci�9�ƕ/3��I�6��h�jK��!h.���S}S ���5L�hr��%��r�/L�t��Vq�r܍|#�[�2I:����1�p';7B�8���L� Z�|���lU����&=�ޫs���~R�ђ�ׇ=��Э�����,&���E2Vv#΀b�M���4S'2[H�JaP�	C(9s�f�\��^&H�hИ�<R�Ý�ƹW}0�֧�:e���Z�%���7$`�A��x{r�=��ڵ�Y���v���r68�C�ws�0ݰu��%k���|E��WR� �M���:�7)�n'G��և���ݏ�ul,Ŧ�9�=�͢,L-�k���6q�/؍Nb߆Y���iB�K����v��:�59�==�,����Z�R��������x��*�?s7A �Wav�S�U�]@�Ѵ�|y��ZVn��v�w}ˋ���`��d�aGE�3y�9���>����#�m��̓r?�*"�Yt�{�a�.��&7����yQ���Lb�b�75T�=�N=��1�ݯ⠧	�Dy�S��u��Q��L�ލ���e�$=nj����{����\�'K+���AiN�1���m�\{FlՒ>�W�^�>�D�`l��5��\I��G>2AWC)�j͜*X�R��	Us�=�W%pf�M�����i���Q|ۣV@QR�XgU��b"��J�ϗp<
�>'J�,�nv�i���[1S.[D�8p��_Q6ڻ���}�E���E�P���Am�}�y4r;7Ŀ��Wo���7+-��jO4��/��c�m¸�Ö��3�y����:�E�}�6
a�A��o�����Ź��'����Y��5��]���,>�y)Xk)��+ͤ��_;w�Y���\ �{Hc�(Dfq�ܜ���3���	%＝�e���Lحc����cU�5m�  ]vӫ���{���\�VDR�8)���Wgp�^8�Wn�܊��9��#��j���������4QW���v�w��d|}��}����2[��KPnŇK�q��Յ�Ie+)DNf�L}���җKp`��*gS=�h:͂pە�#/5�x���4ܙ�ˊ����SPV������Jj���5�wu^�>�8���.r�w �x��*q-RT�<ئ��ȩ��p��^�F�'��wU��4Z�͜����(���e�L�s޺���rI��,�O����;�.-��;xh��B���:9�wLWGA�I���a�������<�{J�6���s�h}����t'J��9-�1�l �[ e*ˏ��
xN�ǌc��.���]���N�J�u-�*�j���f�ܙڍ��/n�U�O�v>x�1��ӽ�̴�Q2�Ut�)qs�i��|u9��ы��:��3Ӵ�,V�\�@X��mM�6���:�?/�n<$3��5�L��s���.��{�z�nB��7��M�;�ħ.��9���tJ���«[�3��,�e�b�I%I�����T����&M̰�?�'������ǨK륾I��_Qj��O^���{�6GZ]����3(V�v�D��<�3��.v���FH�l�5�w}�^E���8�Qk���@3�I���%EVϽ�����z\�α�'�tbLCǎx��j#f���rY�iu�R��w����|t`�@]�\�5�Ԃ�K�cٜ1�I�!�rʕ�Ǥ���{{=a|E�_4�����J��[��������LY�u{B�y2�������OAR�č/*Fg�~�g��A0)���z('pKvy�']�?.(�K��	f����x�uv`�r�T$k�����d��y=�+o-uU˦ٸq|�Wl'�#��oo{[?v���	Qo��歹�A�!P�\g�T�\E��{n�vh!!Y1x��\Uv3�"�����D��D�� �i5+r/�zo@������	��Q����q�ћ9��
��W�v���ĳ��]6/%�����|Mٜq���Rݔ�^���X��P;���!R�}W;e+s�B���ٻ�@'=;<]�2��ǰ*-'p��Rnk�Gw\E�r�������~Z2fJ�Ӧ"�ϷB'��sLqyu�>X��c��[*��A�'R9�6�s�N72Z�q �V�^����P��� �o��	�n�.��y�NTz��}� �����f�Y��AV
ݵ9(!'D�cb��@��v�rh�p 3{�^%aG��wEM���*43(A��7�.-��oIZ�����]��ɫ�BW]�5g���YN1���u��ZY	�Fw�c,î>A��7�[����.�Rǭ��;��T|����\͊�h�@������&y_c��i�A�����&�9����8�h�o�y(*���lۚZ�P�
�q��l�uw`|9��)��:�9]�,�KdWȫ�ke�S1z�����5����v�C�Fxy��]Ѭh�
.�}��u�Ӭ��o3]���z�~�'��>�]������.R�/�^��3n�G��5�̖G-Yf-nx�8�	���b��n>�*d�]��9�YZܼh㳑��p3�1{��Ӡ[�1���V��	���9�o�V�j&�Ҭ�N*�R�|�T��j�f�h򊐗N���穼�{��(�g��W
}�^v����'@��HTr�;�@E1�;�9\����3b����M��.�X�8 �((.ռLoIa&��y���ok>�!%>�zp\��C{���frY;ҥZ��q��"��z��u���y�z�޻(W�ʾ�i˒�Iz�79HZ��K﹊('1Qv���yک5x܃sٱ��PQ�C6>\��e��������Ku��Fon� $�#}t�]ݴ�[��	���fN_b�y�rY\;�k.�V� ֪=8���u״��v�]h6$ׅ�27����AG.�9�7���[	�|:�H��˱fJ\��:�,ڭ��P�{��樓�ŚtŒ�ߥk��D�-��J*Jt6�����o�T�?������)/����i���.3�N�IXa�\�oz�[q�戡W\xi��u����o��2�T�Qs$���%P�.�b�iFN�_����m�q�$���a��e�t� b�h*]j>mŬ��ǚ������1ɵ�;��� ��Ϩ�<:���憐>z�������<mc7�P4�B���7Êy�w5ō׳�?`�^��J�VWk���X5��X� f�]��gwV�g��Jn�ayP�ͳRlf{eG��v�-#m�����G��M�	���0 ;�9i�4�d��=���}�Mɛ�XL��@��9���I[]J�k�B�}�_&ۃ�.	���b�(��?�
�K���B����y�7��Oq��q�{�ø͍ݐf@��5�3=�$|H=hy��<
� S�֊i��4�;�ܾ�u��������=�Ĵ�{��F��"�>kePr�#��;�G۾�ψ6�9/h����7�a����3�U�B��wI���.ɷW��;嬌�@FḐs:�srqt�������]��΀��.�Y�|��A��}x�5R���{]�X�Wb�7ϻe��,q�A{ވ���jx�^�8�l҂����ݹv}،Z2�fU�4�
��V���Te_:B�ŷ&�%*�+tUc%�2^�u�JY�p0����@+/!"��	-Zgn�NR�5h�W�J�>��сE=P���[ɶ�FG\�Z�ϭ��`��.�Q�%���t�eQ�Xg�'N=U��ru`�����-=П�d���]@�.�;��g)�[ϞV�:p�'J��K�5q�&3S] �.T�b��ǌE7�.L���z��l:�ܨa��-$L���YG�c�6h�k��A<��1�a=��5��&���uS�s�U���Klvp7�k4�r�*,�\PX@bR@�e�<b�ۥ��80����n_q��K����192P��d�'�&���L>0�O>�g9�W���m��ji��U�ݭy͗[����GR�0.���)<}���	�F�đ5��fzv�o-y=o�0}���>�cxQ;p��cp�y5M"��J-�Z1Z�h9p1�����Ѷ�[{�����=�F��L�ܡf�y���4%��yd�k�mgC�thXVA���	�{z��{�b� #�Ky\]	�����z��w�	L�9!٥|�R��]�Qʻ��l�gw+�=B����Yޤp��R	������S���l�Tٞ�� ��)}�9�5�|zڶgt��?��å�|�q��Q��:Rإ��\����3�Nj�K�7šT��.[���ݸw�$l���mC2>y��G}V����ţ�t��)�o^��6}����^��y���0�|�R�@Zu����9��9䙧�s�z�f�%�T�sH�[�TB���o2M���v���(W�䲘�"7���z���}��fr� �g��C��ؽ�z�G��yt¿>��I���9_���g����b���!����w��7��Ky�0�R������f*oGM�E��_!���u�pwr�:{Y0c��ݽu�s]e?]IFaFs���,��]܀���e�U�04���mve)@��{:3�\�1�-ָeK���b�O�(��5�&��Z�3�@t�6����
��O�n��G-6�/zCY��<�����(ʾ\E����0�����ÌWH��k$+��{���7���z��t�
E
nWA=-T̽��U�@�WtxU�sE���e�o�!w������x.��g!'^A�s�`���Yي'���;��f�S]c���%�`PâZ�{ZM
�O����t��
���;�׵i@�zm�
�����8��:��� ׼��|��׷�N�=R��X7�է|0�� �7'$�u]�5���j2�������;}��Ր�;�T�Z��u��eb.T��IV&��K��M�Bĸl誇]Iպ��w���NL�s�2���0_@wlCo���y���죔�So�l���vA@v�%����dYZ�ۢ�MXn���ҽ<����)z8�+�3�;�cނ����f�0�%���#��m�,wh�Q9�nVa<�3F��{b���/�8��>�an�F
-���Xv붆�[�,R��5�no}8F^���&�a>qz�ٌV܇ �;p"��^�nKbE�#^��כ^+65�IwA{y|���;yW�vy��^W!�"��z�e���
В����"���Y�9�}Kq� �8��m�Db{�ѫ�2n�cC�N�� �곭�i>x��u�ZP���M���=|Y0o�	�����Ү�̏���U�t�[l�4c�ڗM�\��#�����Ka㛞�4,����_���U'��"���C~b��; �ᰥc��U����e-c2ѩ9DKBhb�'+:;v���Oo��ͻ( 	�xK]� s��L�`�_n�A���llvS3�fш�1p���+���۷ä�(�x���}�pz��%;���.�l~��i���\�}���e�VK*�󗨷�_���@���;F_���ݧ�\v���ǩ4�����A�����q(C���pnUR�S�MwA�m����+���\��i^��ַ�7����[.�~�{�8H@$$?�C꯾�rv�=E~�~B���Gk,m��#m,��[ܢV;�ܔ䶌� >�(��C4�<7�SVu��wH�����/URC���~���0Cx]^H�.
c�_XdN�R������FÝ��f�l�A�x�Y)E�?u:	�,��8�G�'q{����Q�7x��l�9]��WV��EH���7�	܅>a��Ա��D�<��q��Ջqէ�24,j|�b�M�c)�&�^�(�O����ܯC��AGE��\�r��o��x�Ό|Z�^ۇ;⳹{;s�-�� �:�����4�[���%}2��5'��	����YO�![���&�Fj֙u8|4�}d��Y65�c;gU��6�0H�b�d��혋�[cZ����˨�e�:�_P7g(k�Գ�C~|
E�O���7��-� ZX�i�\�lu<�;�H�z,�j��b]7��T:��:㵗$��GJ�F��ێ��V��w���'S�\`j�{kw'�M�q�{����V���t#�^�~���V�rpSv��wr`"������|�7-s��Up0´<�O���Oj_)\)�1��Z.����Ѿk����.z�v��\g��v�w��W}�9:�OT�hʳB�i��ޱg��lB��]��e`�c&\=$�-�XR���*�w(���� �=V�����ޗ�-J�c�ys)lٔܚ;+��c)�@�(e]�uh�$��8��0щ4j�J�]�a�yN�\�ܜwP�6����;�!.����LH�Y���j����N�j�"f�����h�0ך�7=ݱ}9X#Bҕ��j-�N �PN�e+�h�rTe��n˕{�B�6��zm�mU�r ��O.�왠���cf\�;,�(NF�0J<B�'�A@:�Nr��̝���6u��w ��bx»�6��vQ�4�N��� Z3pvܭ�.�\h.5%c��77�Pw]F��B�CQ�MWaKz�j�x�Lb����h���k�� @F��ݫ8۫aF���#F9v+V�ƅ��M��/g7f
���0PFt8����1��w�p��ҟw;��o�{[�[��5��A4f��|�X��K����=c-�4Zs^�Iz�j}O^kQ��5�)�]�7k����9�73# ����h�6��o;i���ƠJu�;�p�ђ����'=�p��v��V��ޓ�LdXw�����U��u%Л*@ٙ(�3�.CFX�n��~� �d�f�=��n�e�]�`�4,�/��gu;�W�۵X�i�E���m_wSo�����v�7ۺq�e)"�7�n������q�C&��ה�)k�ӳ���9���"KM�{�|:p�ܨQ��w��"�_=%wMѦ���i]�cօ�M�Xi��klεAt(5�'������Q�.�-N��c��UևW-��!y�P��F��<c\�Ţ� 1;U��t��q_0V��{��',��t�ğ.�p��P�]��OC�H�n�.��i��?N�SN�CU�(v�c:q�=_Ge̬y���lji:Z�݈B�=�(H�g\�n��B�٬]�,�vbս��b��H�ў3�g�"R�b��a��������W{��	U�4"䬢��ݔSOZ�b�B�+�l :%V��,T.�=g���H[��������:���/��nz :7t��)�F�&��Ս(�B��(�cҽ���/U{��{��Ua�j�7��g,�ԅ+ !֬�hWyez+T��9��x�mr�Q�cxr�y9;����NR� *zIŘ���h� 4H]	 ���ѫ�Z�3Iv�ܶ�jj�uk%��.�+a�zS���Ǡ bCR��xh��=���hZ�u��v����a�2��Cu[���cQ6���ű���U�����o.N���LcA�U}��߽7h��N|�מa��sgP���^��n��I
�ќv �����r���V��W=Bp�6��t�͡MR�d/0jWlK�UH��k�'a��xH7:��Z�lƗ��X�U}NoX&�� �y�ܾ3��sޙ�jA�)�j`�}�-�n���	5@��ɁJ���M�7!׶���;�q��B�igd/g�
z���E�����q¼_Y9����\\y��y�'~�c�ȸ��M6H%�ε���ri��5��l�<�E���D�zr�wJ4��1-�����kq|�����e�K���(��������a4�GU����JY΋m}x����35X4� ���Ui0�v��=���.�g�} W�}�hE�^�%֚%�+<\��=o�%��.��v�̂q�qk�Q���}��֢�Y���=����4q{auBQ&JlǍ7�}Ε�q���PZo��F�kJz�s�E�J�K��v��(���i�
θ3��\3\��ݲ��	��=�V���h�����
���a��s<i�(կH^2�+��nn0�=�>��n�|FMD�1����꒜<]06�<��Ӛ"cz�3�]�ĺ�����ŕ��"�ck�T��6wd�jS�cP�Aū2WI�������k(-C��/0���4s]��v�\We��#kkD�w�}p�l�<a ��w�V}^9 .��IV�����^�6�����S&�O���5�'g��7��w�=� /���{�u�;{�r�^�N,{+x�:�s �@u���A�W�k[�i~��.�̟�{�/�b�s%��)vN�Y���.��0�� �E�����G]����W��`$��V��ҽ���
rQ4���hG�\|��xܽ���k��h+
pS�'��-�5�K�v�2�3,�t��.�B�	�P���N�!�:��ù��WAvp���k�իd�L�6��J���pt�o ��X�|[VxrH0�;��ޕ
h������o(��f��]�{����i"��^|�2�^Ghw�� m��5#{�L���h�Y�Ú�C1p�W���$�6�G�mU�Z�`�7����Lq�6-оTb�fЇ^Z�̂�6�.ٍ�,e�x�殬��F'K�F����2�l��7������ �b]*��e��^�v���9r��-�Bw�E�D����-�G��#ʚ��]WKT��ԭmZbʦ�XjW6�'gSd~i�¸5=oE�7ܵg�	���ͩ%������ƙ8ܫ�X	�9��'!-)v����A�6��"�W�����6@���7s3���@�k���鮡�]��zU��+m�)��v���~��"����ܖA�2�gB��n��p�h-P�ni;��	Ï)���)�O�.G�ز�
�^�ö�T�k_o-�)�8�����D#oN�Ƶ�o|���YaV0�A�xe��;)p팾h��Mc�� ���9��k�����D�����X��c��pv�D1�K��Lmm��Ѻ{������yFe��������]��G:k�,���6zs�1�	���L��*��;���)S{Mlh���1��IY�T�hV�j���|�u����>V���UK`�ؕ0�+�Q��ej���I��2�s�J��=�����(��C��i:jiZ�U��]ԏ7v���D�g�l�2�U;��@�'+ٶ՞ꊺq^�:_?���u��yĴ���Ɲ}���/l�.����ܑФ67��OW.���$��v*D���d-�gۀ��mWr8��Ŏ��j�ȣzhT���� �Q��I�۾9��D�5$�{{�Ծ�Ý��ᕁ���}j��{ۆ�ǁa��� G���`Gh���nE;�	٭�uo9N���W9��7�{����	�����1	��(G[gUC�ԙ������L1/�_e� s�f{����,3wtX�qN��|;CZ:cB�%M�����o��3u�Ƅ�����B��GG"Ĥ�#-���8k�.��-M�6d�f��D(��Ou�uf�M��9P3it��������������	��U�˒w�W��ˠKt�W���N����ݴ?^�O����ǳ)r�i/�y3uYP�F�]�e�W8Wru�:��s`a��i�"�Rh-<J{Ϻ��P��E��>$.��fHQV�k�51'9v�bJ��i�����ua��k�W��:�"�}��=ɘ:�k�s�`�,x���&���1�xt�=E�<	]a�=�V��;Ѵw��lL��~�k�rV+�\G<�x�*�{W:�d�Q({y�M�`�p�K{qjw����P�������N��<��-j�y�R�s���h̬�Kov�.�8�$L��4�2i�Sz�k�,g|n���:��|�����d��t��ҖJ�yHvթ{��@%˦s}�J ���	O��L�i�����Ւzw[m#��=�7w)�3t)$7��K���t��F�@�7�k4D�t��30իJ�m����o���=Z8��D5�P�^�G-fiU���Xj�N\��*���j�5j��{x���B�-�!�<�:�p��h�Z[�J�_m|8{ٸ��iJ=G|��ow��8�M4�_c�Cz��}t�F���'kc�u�5y,֗3�B1m�U�)S7����k������t�4w7NqC��d>!�4������k�y�7'*n��#���C��彵�Y��u��^��y�	
�t��;�&e�W!z�W�֟�GY��u��Le�z��Q���B#@�3r�k"�t���O�;�)�_g[���lW8�X�hq1�_h��*wI1��#Y��sO�s�;���p�#�FRLG�+�d;��=G�֎�n�yB�����:��b���-L��&X ���+:�t��m-�S�[��<�e���e^�5z���zP������b�ק�����H�����^�F�3LK�~�����8�O!��*�L�Ԉ��Aaͫ�8�*�R0��Y�\
*FC����Z�I$��|���fY�V��1fQ�q�Q�M�B��"�y�Q����f��}�ZSB��L��Y<<-��W�ٜ^�����O��=A�p�
��� 6fL��2�����F�;;��IQK-��a��	3�`�1����ơ��"�̄{B��X���t��^u����iG��$DS��-&t�Y)�R�c��z.��V��ݕ�ç\�8Ɉ/�`��D�s�;�w8��<f�PnJ��ga��-⾭V���L2��A���9�����^��T�2%�V�(��Y��b�^�Ҵ��mhO�Pqފ�{pB��{[k�f���O=�����ֽ�d�hȹ|"�Ba�����;������T�G�Yĝ3U�E���z����9n��u��$��O-��}�a|���N�MΏ.��#�mm�iǹ}�M̆n�_�PG;�%0���u�Y=���J�5���4�$}�"�Hi(�ܬ|��<bVn���1���ݬ*E�&t�c`q�Chv�:3R���=��'fF���[�Щ�nq����q�b�t֫O������u�m�x�+ё��v.��>D�Y�=�ۜ%f�*���#���ҹFfH~��d�ϲ����X�[��]5 �@$M�����)��.�7�����J��0X	�b<ۂ�/���jѩ�ws����g��O$AR�:�5ـ����q�9���ˋ/<�l
Hdɺ��t��VE-3,M�@���m �V��P�4���4jn��ٽ-(��郸]��Y�֎K2�O^ ��L�'�7h�X/�Ɋ%�4��'H��+2��@k*�'�h����P[(s��Kz~թ)�T5�{B�Οb�`���cohY[�[����D�e��ke��k�^R���"P��A�s�|�.��9�e�Kl�d�R%j����y�zHGT�=�N���݀-�+sU1.��t�¦�12F](��ܚ���uې����y]qbYH]�L�g@gʮ��g0:�� _m��в˻=�ۜYNt������]cW��SU�0i�}��F��uh]z2�`\�n������Ȣ8J�����w9��\��UhsX�J�F��ޣP��@�JΔ�3P-��`��9��\Ǩ�E��jugSB�R�p���%��Iț�>��>{ a����V��m�_/������(V��ga%�P���;a���ѦA��fuqi�)e��1�����s����W������k4!"��u��� ��Cz��r�r���:���8��u�qV�sm���KQK�.���ծ�/���?hdH6�\���Ԯ�����G�+z0�ݷ8��y&e�V�s�zQ��PEV�V}�&ih�O�,�^S���9s
,��Q�'Vѽ�8qN��4ǬW4�Բ�K����s�X���=��(+;�U��*�!��^�8���4�鿭Gm��k7�6��]F���Õ%/�s�1̅�G#�|�w��<JpV�n5tn�
6��AI���#i��h׶�R�����~TE�F���ܻ*֍b, 9\�C��h\n%B�;�)CP��0ۦv�u<���+Rjl����QX��BmõsN�iqn����Sޤ��I��Sc���:*�W`F�f�ӡ�S	b@[ŉ����<�v�F���E�윝=�H��Wݎ����@V�u)Q�<���*�M��h��Hn�8�4�wh�WvAB;5k��&���!wJ�m33k+ n�r��1l�\εaX�|�dc>�GVe�X���R�z���[LR?8زt���4[�����=�W�J2d���y������ó!}V��.�7n�.�nm�0 7��q���F췂��s*�B� 4�x��/���vlt�z�;-x�8Й�+.�]�yM��L}\��U���|�&�d��W���ŠCm�:!i�Mф���ⶃ�Z+�U�9�{�IҗH��gyf��.B�Wx���f�z�L>x�Z8��<�xw,.�p���0��lV�;\���I�Z�����gr�жn�}��H;Q[
-��i�/K]��'9�|�n�\LQFP�+hˬ}�f9�MA�I7�m�N�����S��v��%i\��/&vӎ�X�IamC�G�;˅�� �;�z������\$���eC�sh�N5���	��7��K�̴\`a8��V���e��&��-���j�^�x$�R�m���͞�=[3�w��Q�3L�hv8R����e.([m�îΤУ7b���csn��������չ�PQ�g�@�M����fmfh�ǀJ�9E��G{�K�a����,��q���$���X����([������2�;�^Z�5m�B}�Ҿ/��6���Sv�nM8��5�	uj`�ͧM��ܣ��7Fp�� �m�*`#�U*�#�t ;�l��S�+f�
�%�E�G��2��yZ��I�h���o�f.�a�!��q~7HD}�%Sc�|��I��7���U|ꭩ�w��f��-Q�-���K����뷻O�p�y'<�+m��Vk�yU?�4��(�K_�W)b�b�J5�1�m�<C1Z�VT�1)h�A��k`�FE�6.Z�m5KZォiX��e��ATQLJVŊ-i��ZL�-m�V ���j(�P��b����J�E������Y�S��҈��h�k�b�EU�X�P��r�R�r̊`�ڵ�2⣖J����
�DTU����**8���:�*�b���1A��c����
�qa�l����#�j�m�\j��4TJ�Z ���(�*���0�U1̕V�u�9V�XіօѴ�Q�c��X��&��*1MZ���p���S,�V�5
�0�Mq-is�Z�++-D��R�����R��-� ��̷W2Ԩ�Z�RҲ֭�%h[J��X�q-�Y(ѭj-�-��U w��pNT�c���􍋀�&W��Ո�PT�S��l]k�C^��P@�&1�K��ј��֨�g�}��\}�l��O�8{�s�i�li��t�C|��y��۬�i�6nv-�I�K�d��^|=�tC9w���T�я�E����o����7F�oyM�B�*��9˞��L�S�[.��ҵ�SN�ۭ��6jy#�-�޼No��w��R�e��Y�\qW��x`�݃����5g�cދu�G^��w���U1�/x��'±M�����ϺXVp���{=�����W��/>�dϐ�'�b��ʘ�46��:w��a\M:��v�VK��t�n�Zh���|Z�K��l�at	�b6��U�WT��`؍ʶ�M��a�΢���^h��= ��O�y�^�+�{�K���s���=M�coS��n�c�����h��c%Q��`����]�s4�z���ˆ*�3S5�V�Y~{���b�vz	搸�����^M�t��k5�������"=h^���wo������'5����u��.O%�nAa�{��+ݖIƩ��Ό��+�H����ܤ�j[M��.=U��Zf��e�ټ	yt:C�~��C��j<d�;3U�ٷ��R
�	n>ޡ7��7L�^������
���>���6�����J�wUɔ24UP�=���syir̚��@6+(9�ʱ=4��3��H޺S���O!_CS&�g5��n��w_�yBށ��ˬV"گT�-��w�}��5�)�+�{KS�i��=�~Q���y�E�ڤh���Dr�6kY5��u^<�K�v7��l�c�^ĳ�yqrob���G^Y��v{�$��T�Q�=����W�j�B��	���u����̵1��:f�d�t5�HM^=ILߩ�0�R��W8yH���z��
���-U���M�[�w�Z[q��2����*V�X���������W>\��I�sf%�ٕ����I-B�2���3�鷜�j���ic���(౺������Ô�
i���&]±6������-�]���~ȓ���Y9��8��1�Hi��
�|c;�dI�Iw\���y���Φ/&8wK'�_�jt����+��WV˳:��'���Ҭ�r�v%��X�:����vY*I�V�6���h�Iwe	�du��.�i�Ur�]Ej\%�k;�W��3���*Qt��؀ԳG�P7}x-{�B��M��/[��-�n�h��f�x����93�n��y�N^wf>jթU�����^.3��Bz7%
��);<7r��5&N�gm�b
�9O>X�5�˭���yP�n��
�lWn*��,z]���e��1�spto��}�s��Ӣ+��>Y�7��@�he&Z�'{.��
��h<����;=��6���k~���C�&h���}
��L�,J�W�f�Hn��X���w�����X��{�Y��I�Hm���	⨺��Y���XL{Y�z�X�P��/�I�̞��R8�a�/1�T+a�w�&�����oM&z��J���|������N����76�E��E��׈-U���ɣ���KBS�Թ;���11:c6�Y&gJHʂn���v��=lV����K_���ev��E.Bj�}�Y!�pJ��Y��Pni�w��)��ܳU{��L�̻0m�l��,Q�Е�i��W�$������'-xe�����w�h���;��V��k:�V��X�A�����K�����ݡ�EI�!{�`�V��A�G��a��k�V�Qՠ����ɛ���;�fuC�I�=��:���I�8��Zg�+p�YT[1U15{���<f�z�yw�9��A7Z,Jy�)ؗ�.EV�����v�Ξ�������0a:u��9�xgz��s���WC���z�g%���%��3��U��F�8�oE��>��U�r�=�,)�Ѹ0o�ҭ+�V�����S��ȍ%Y�xN��m�-�m,WM�Bx5�s=yˢ����3��+n��&��:�j�������:r��ƃ$���DtP�4��[��Cs6a���+�����1!������r���M]�����7u�޹ؐ�����ʢ�<�K�,U�������
�"��V�e���*���7��ԏ	V��z�=m����Q]X��!�Y��f#u���	��-��VU�}g';���Ԡ�:n�:�����������;~�.��������7e��{�7�U=2�����P��ǁ��V{�,��.�۱���h�-�K:�|�ű@f1�i2�r'N�.b�qW���s8<���u|�9�.(s�b̽����z�ؚ5+9X�x���vd��(;�b�����޾Sr*�E��W;'Ԇ�&{4�7��/�u"�H�f�P��o=�l�F&`N�k�`�
�h'�z��M�Nڳ@�B�;Yz�R�9۹���B��2��hp��
���rln�e�t��g<Rj_�{�-��ֆ�C��21yKc��p�3�w�M��k��xW@��=r?P;�kw��x���1g;��&�g}o�E��������uuS}oZ�KK;�����}]x)�A%[W�N�P��K�[05wsf�^��Q���g�+�,	yTR+�*n����m�sb7��{��>��muG@}N
�!z�8����QL�+!�פ��%��b�J�UW4�y�`ћa���I�Re��w���-�x��矺4"��o}w%�@st{�}D���r�:Z�}۝��ƿTz�g �}�X�c�r�+�WWFB���T2=�kh�ш�`�ʆ律��_R�õ��.���9Y�ז	���Oj��^�=�d��ۡ�t�(Y7�Y�KN�g�h�}Y�=e��T$�{����:a{�YA<2F�Ϛ%7�p��d*Y��o9�lN�^$�S�y<����u��A�w4����B��=�'�v�!7u[&�:7/�}�n߇��.~U�(V_�W[�g*�K^�ynT�D�Jۋ9݅:����%zx>��NL�Z�P�����N�u�罝�;4T�^�qĹ����3gk�ą=�Q����hU�{5#@JN����⪵��J�海������t����J������Cp
L�$B�:����!jŕr��MV�Ja�vGw_�yB�#����q� Sw*-�<�'��{��L��؜��u�ev�]e�Ê���gS���p�۝j�ѳ��<�u���uC{Ի�ð:8���v�͇��R��Z�b�I˲�VO�ʯC�W=[^��ˌI;�}1�v<��h�x��3��B�YI&�ᯯ��KY&�q���;"�5DU��g5�yXj�7�+k#����hg'���I]�$�E\௃�7cW;��tD�yrR�I���_rٺ�iuu�;;)��Խ<�����ĵ��yp��{�͓��^��nI-\���r���Э6H�=;����q��%���T��f�M�ާ����b�ա�����ǔ��n��aS���Pden�)�Нf����>T�|ߔ��L�R�2�eQ�l��y3�U%���מ�q�q~��/'��U��%2��hau:o�\Md�g�TF�W��~D잖o2x���������V�Я�����,7E�"��eT6���nrT��C�����^�Ʌ�*)ᦍ�����!���sYx�8�zߓ��p4np�>��m�{ ܔ(v�#��O4n�+n�A�X�M�k)����_������B��弨B鱴�\���V�f4��Ҷ��.�fM�M�����wd]��Τ�ՔWz��:����5�wˤ�Osm;����ybۛ�9C�;��NL�}@\�w��޾��ױЮ�s�%�L������[�V��W�M��sԴ�LEpٕzП�̆hhm{r.�Z>\�3U�-������#�n�Ag�^[=�6އ���dN�\n�8�`rp����K+ (#��&.�.6�{xw{�\���"���1}�"pż��m�����t�
Z��;_�&��w<��:B�&2��V�og�:J��1>sp�?B��H��W�#"ҷ~m:&��Ԕ*�=�R�ݣCj�Sn u���B��.;$
S��\Uv���y�tɭ���P[�f9�cՏM�c�`cu��_j֥oy�J{��-%�p��Ʋk�O�oݪ����5P��o�z��.a����Em4�4�2ëm�im�L��{�ޝW<�
j�Sh�K�!���6
�S֘D��\,�&[Ժ;���św�K�Ji�M֋��JF|ؗB���\�Y5���e����i�.�dn���|��xs�-�:�i�L���F�oo�µ8����W�ˇ)������f�E�d�+Ě�;�\J�����=t�'Y�Rf�Dn��Sޣ0x��,-��'j�2�_U��<X���4�p����F_l��"�S�z��o�c�N�jV7	%�N%���ث/P��Tb٨�r�tΓ5��<̌Jȏ4������\#��`d���J,��^��`!;X8���6�Ί�b�����;���t6d��!�}g��yҎ�ju���qu^�nWC�j�f]���y���Bu�j�'�|�fM��w��5^�OƃY�<����DZ|���B��h�<�U���[�6}c���۪2��(��W��Q�g3wz�v�cZb��1�އ�+�z�m���<7�B���̭��Y����*���!�\�bg}�ѡ+��v�w'S�S�M�fb�q6��­X�ĢVl���#��Cg�)����Iۿ4ڋt���u������E*z^t��z��t.=C�n�s-5=���Ƴ��N��z|�'a��-:u��y��#�v�~ِ;g���>��h(��N��U���-.VoeXV���xů)l1#��]�f�SZ�U�jdY��;Y�%���j���$,N��5P(ٜ~L�C�H�H��9��^v�x���+$���F��I�Pش�<4�F�)��W�_x*9��� r�0��l>=��j�x=�(�g�7*����k�a:���wycp&;yVBs�s�]�(�<ϸnN��CŠ�D^��;����gu"��jN\�K�ɿPg����ָ��?/��۟>�5f�pඡ��v��殨�m��i�R�2�k�q�Yn�K�;-��Y�&em��YZ��!���<�ReSB���'Һ$Ebu���!�;F�ۃR�f�[�֯0�t�W�Xc��'B�N������{��<[�B<�"����k�����Ac˘TS�A�pe�`5��<'U����z�;K'X�)M\M�kY�ºu=t�\1<^���o������c�Y�9n��1�2異���{�{����q}�����^.�Gޭ�}�v�^)��l暈��	u�w��˼�D����ⴾ{��.��ƅfjf�۟4�T �N��B�n�U���_bcywt�5�踐�U�de!��hM�f�R*u��>ȨZ��>���n�Zj��ջ6�6�جq�u��"��L�}X�V��D!��n�:����Ɠö"�E�gh@�j6�o;����*�l��E��!'�v�
ָ��UG��Dx���.���i(:���zu,m.�1�:;۝��=V�Z ��b��ϭ�L����@�D�CC�#5U��Ff��)�R�B3t��-���yq=�-����=ѳ�o]��LKǠ�쳼N1�alj[ņS�W|	�M��L�be	�H����+9AY�+g�}�WO}VN���FS�}5��w-�b��4o@�qh'�
�d����O��������[��c��!6������oS�Akph2�\er�T0-ոU7����s��K� �D	y��@k�~��-�����U�U�wZ���i������J��2}�qz�����JM��g�]�$��iD�WFqp�f7�ǿX����;��(�duqjWkSu<[ie4v��d��ؓWS�x�@0\�9-W�(�Hc�4�����_�Z1 6"_&N�yL+��<�{+}�i	*�d��w}t��	�t�$=е�8O��xx 7{�X)÷OY�]��/;��R�l�L��8��9/x!2H��n�c<����l,�}c����3�.�L��Dr�b�w5<�W�O���j�����Oݶ&*s��=M���;JoH�՚����%��������޹m�3�gC}��w�ۻ����{�t�Q>S
�]#ww�6�c -S#��c���'84x�S�#��e �a��>C�k�W$�P�6	S��20�є���!�1�y �mb��c��� �����$d�G��"Ms���z�����S��6I�����ޞkR���ǔ)2੮��1:�H!��C3$�V�Ҋk/B���Ҥ7���h�����ڑ[�*���L���rI�����4�^�Kڰ% �a�K�˾y���JȺG����F�2���m�ܼ�)�"�m��ݷ<g������ס��%��{�vb	�CV����-�/�Owщ�������I�V�T�@7��m�r�]3i&�(v���|��#�
n�ǩ�T���;{8��Ŗ����v��a�?Jx pܾ�v��^��^��^[�}_{5�7�&����;�i+Y8l��=vv��U[{Ywd1�ib�Ȗ�m�]{M�:��I�X�yH�}K�"o)�K��9���pj��lS5�
�*1��d�|;a�?���2iU�gq�ϦNf�zq�7kh�h"#��Y/��4";�]�p6�F�I���^��biв2�<�Tw@����Xk���k���4��qg��ӑӹn>X)�|) ��Ӊ���`ԩR���$�S3dt`{��������S���	�H�t�X�Au.��7��w{G�Z�Huւ�H�R���%�*�a<0;˳j���9��a�F����@��A�ZZ��˖W�+mm�
ګ�,�Q�\-kF9n���+UEEJ�ff)R�[Z��Q���*Ѩ�\ĥ��֩��[����e(�F"�D�rbU��Kh�cU��u��h)U�Z�6�mE�h��ʍmmh�Q��:��̬ՖV�eR�r�KaPGW�*,�ړ��
�E-�2�q��b�B���J]$��F("��֚��Kj�%e2��R��`�r��j�-���(.V��j�1�t�0ƌG.&C�"�F��`���-�imk�V�����2)X�-c�mJ���mZ�)mDm[Z�\ʕQAV6�3Z��Z���`�����PZ�ABլD��b�Ub"J1d�[fS�mV��U-*,�̮۫U��""*�Q`����5�Zߞ��Ӊ/ͷl!���&���M��g�+y?5�8W��'S�^��a�r�nX���h�pLp�"��7^P�|T�"�B��#��'T;;R`G~8Z�J��=�!sR�R�{ϐ#����\��n�-֝���d�u���F2�nE���=G/f"w�;�����-ۯb�v�B&�픺8�a� �J/_��.}VT�u�t.���*��ѹ]�����bYָ��{�^�����ىX7:���n�:����]*��+����l.4����kEfD�ښǳ)�\�elu�7�N��._a�V7Cy<~�׃���ł�^�4�[x�^*m޾y��9VT�&�[�Z�-��+(5����F[#�������v��E^����(GҾ�Ճ��hP}�}�ڏE����:���@HL残o�t���dj�>�aP)���5�l���}s�Cg	��k�;�G�K.k�8�JܬT�9��L,)٠���l�[7��eܗs�2f-�yY�oŉ�~���F�U�on��BO�f�Ӓxk@xj�����ԯ�+2�u&ըn�|qlU�+"�ػ"��t�=��|���4=߷q��N��9̘'4�����)�.#;c� 7j(_�;���Ȼ�gxz�jOb]]� ��1�k"h!��G^Pk(�n��x��U��GM�7р�K�Ϊ���3���9����am*�ݚ���6P��̘�����wN{S*�~[����[qCͳ��v��*�)�řU���g:���'�
r�j:�o ���ŉI��{a4�g�fMk(6+t�f%�ϕN5�gnc{���*�&:���v�r�X��4�י<�Ӛ���S��ʇ3`���ҩ��ׂ����z��Ew_���Gپ�wu"�m�� Ν�e����NzƇ�)�<ۨ��i��˻$�w�9	�maZ��:#��Ȕ��n��qOb����_F4?�v��ǭ����-~����}��\KӦo�EϕD��mL-,���р8{��ʯ�uc�[��V�V2V\�8���Y:}9{P���,o\�m5P(6�?:C����	®%�yS5���Z۹@�z��N�<iA&�����N�0�j�ݬ6?�zNIʉ�k�K)�1����P+8ACmK<��|٘y�����;@��|.�r?�H|Ϭ����[�EXH��Ãu&�Πp�A=��=�͊��⧷�۬��^�~���qIG*�C:c���;گJ�]4�{���i���v|�g�V^��ݱU'�:����TnT7��عe�rA��A�D��"��霵nt^�[�˧
EW�U�����_1�P�P�x����T���YOM�e^ݽ�cg�z�Ah��e��<���N'iv\�z!κ�{�3щQ�osq+���6��F�ϟ�!��j��ȵy�n��i�����t���/�j�W/=�w��w�l纓��n^{9�T�����:�mՔ���2�;֤g*�X�R�k=�-���J�ÚO���xG/�����uT�&���s�"��,M�b�jF������N׵����:�����9O]�Ƭ���p��2%�ږ�XL޴pO${]���.���;*�w9�+R̞�x��VPz��A>&� i�-ट�o�N�$��퓌���q��z��n�0j�}����v�1�ڔY�C��$:�6�畠n����<������S�ɯxذ��u�z�M[�e�3��*���m&��t���<u"ͺoP���Qg{��<��L���Ե�� ݨJ�v�f�*�\v�j[����n���W�N�(�݇��=�K�����{�ٮ���vg쟓�C��w��u3���oXN0�5���I�~�,�g���N�i'����<d�}֤� .G��=�p2�8<�����5���}�}yd�6���I���d:��??$�I�����1�O��~aP��E�a:���O�Bh>̜I�=�ម 2 ��\vm
��?/adg~��$�@����$�8�|�oX=��N$��3�X��w�z�̞3h�rN��LC��̄��'�*�8��@'�D����34��}�uYHmU�w��f��?ZN�` zɾ�Bu!���N0�O&�����2C�|�r��+	�<��O��$��b,�;�:����w�׷��oc�s�=.�����RM!�:dm$��g>d��<-'X�ۻ�q�������xj��x���a?0�l�6������>�Y UW�>n亙{BDM<~��?k�|��O�b,��p'䕆��4;�N0��O�a3Z� ~a��'���'�ws�	�C�4�Y0�!��'ƯY'�*wZ�����z���u�y��k^�3�&���i��X��N��&"��C����.���7�dXx�I;����ST�H|�f����
Ϥ>��Y�#չK2���g�7�o}��y�����N�)�$�
��+$�z^a���;�l�hzw�!�J�P氺��d�~Ȱ�z�s�2�>��]G�>���'τ���svĺ��/u矻��I����0�'��$�
��/��$Ru3�d:����~惬��	��<@�-�@������$�'����I���'9�\��=�u�~���i���a6æ���!6r��'Ԟ���i'Qw�$Rq0��wd���s!ԟ��nw�*��D�O��� �V+GCUYF{�7,x��\��)�а�#
�7�o����?#.>ַ*�y��7����U� ���^3�aJ΃��-ɛ޴�Ӣ���W{@����&mIvj�hY���	�����^]��Z�
zOh��Y�`]�Y�.�;/��zչN7��~������&0;�L'Y�	�̰�g��������<�I�u	�o�4��,�{@�'Ru�Bm��}���og��ᧈ�I�+�N��=��1�s���{��t���'!����:��
���0P���<fوOP�Ow�����,�VI��N�qM��O�8|�\xzϽ����k��OG�Mf����v���0�>d<��?0?!��a�{�~d*�j)<a�wX0���m&���i�W|вO�6N�8�{א<Ͻ�G�_I�Iw��NO�W��s�&�4��Ӻ������,��$���8��~d<���C���ﺓ�	�x,!�CS��|��>f��j����=B܂}�q�6N��_9��گ��M��~���7l��g,��v�$���N'��2C���O^�:����q��!�{�I=f0���Y�I�6}��'��!���ԛd���9�����sN�{�߹���=`w�`���5�sRv�'ό�a��P��6�;��u!��=�u�8��'���>g�M3����O�|>p	�=�}϶cX��^⻳���=�߽�=�qP�g䞲z����4o�ԓ�M�rO���7��<N�7�08���<��VC��o��}��G�>��}��>�5t�q���G���=�ڽ$�+��Y'�4����,���'R|��(@����Bq���o�'��$�������`|G��o�xA��ͬ�'���d��xӏ��<I� t�ԜC�Lg_e�:�d�;��$�>�d尚���=jO-���n���`k��z�� g�=�@��>���,/���Ϯ����۞�o{���G�����j@��}�X��xY��m��!ԛd�Y�Y2b��(��I�����MoY��1��ɫ<π�=d�dxs��������Y3�:�"0Y7u1�W]9��bRI�@�̻����:�o-�t,j�Vk�1�(.�<7ݖ���j��1\T�ܣ�*��^"��\�����x<�"ݠt�����һ�nyӃbN��^�q$�kS�9v�	5]�{��[=�?z�d����Fݮʻ�ˍ��4G���{P��2x��ϙ&!Y�C�'��u�z�5̇RzɈ�a�wD*CG,r�8�S��d�l']����
��ڹ9މ�9"�0�2�|�%O�g��LgyBu����ԛa�<��Y����I�
�~�d�wy��'��7�d:��L�5�!�
���d����ށ�tIϵ�S��]��ͮ[#���I�L�0��M���|�3S~�N��Sl:�hq���AC:���	Y*d��h:�$�o���d4�@�&5��o�iߺם�}�~!�
Þ}�l�L�"��N�`z���'�VI+3��Rx�0�&�c'Yԛ=�~I�N#��H��a��E��ϡ\ĩ���(NMR���r���(�x��0*�<t�}�@���>�x�	�M��z��N��`|�����''�o�d�C�M���d�l���O���Iy��?^E������O�Ȁ��st���ߴd��')�C�&��w�Xs�
�gzd���Ou1����M�βO��d�E�}Օ.T�:j�+JŽ�b�M�i��Y:2m'̟Zk��N u?rú��0���$��	���~`~a�i�$��T=w;�
�2s��|��6�Bz�2|g%��ӽ��>�w��;8�m���	���ԟ2v��i?0��M�����O��'���m����}��|�Β{�'���]�&�� ٛ�Rɜ������'��{����P<q&�4o�,��M�����?��N2r���'����=��M���a�}�8������ԇ�?3Hoϟ}2B��EU}��L}�|���#�O���7�`q��=VH|��M�	��d�O��d�5<�ćx�N��q��rgs�q	ԗݿ����:��"��Y>ׅ�#�g(����(G��"b�����eV���h������4е*dq��j���ĝR�tU6���������"qOP����"���F���j�m}}׷j�@�z�f��S.zf�FM���0r��%x=0l��*��tХ5&�6�-jJ�~�d
>DM0���Bu�0��೬���Qd�&O�'~d�Rxe���4]��I��Y>����'Rx��>B"�~�]�(�*��k�}��l|}�'Rv�:�Ę����O�V��,����)>E	��'|��(@�'�f�O�6grO�N3<�w�q����~���]foj��� �G�|:=��>C�q;�!XO�<�^�<f�<;ܓ�6Ɍ���:���{�Y'�;�E'ȡ6[��=�M����6���gmd����#�{�|���,�zβq�3�YgXI�=N}a�:�>9߮�l������2b�]���^��5<�'�a>�{��5	��3)_�;Vr�����/�ϼ����$�!�#�	���Y��t���=g�3�'�O�����I���l��Hy&���OY1ٮ`N$�;U��/��3��X�r��G��#�w�|[	��ޠ|���nj���6��ܐ����p+�I�6� ,:�l��I�0���Y����CI=E!����[�5�?����1rC��	#�}������aud�$�s�,<N0��2�+�&�Xq��Lf��8���:ɦq&����k��%IS��ߧ��	�����_\�-o�� �{�~�t�"=�)��J��&[s�C�L�zԓ��/�)4�a8�e���3�M�Y2C��d�8�x����C�ќ%�+�ț���`���9���L�W��0�����"�x�s�:����d�&[N����a:ɩ~�C�z��xe��<Cԛד�χ��c63y�D��O'���e��;�i�0�M���E���u��w�):�����1��2d�l���X���;�@��&?g�Y`h�H}�|D���-���^�;f�uF�rYW+7��ץ�?~��ՒlO�Q��0�v]'����h��΀_#��-�EwӸ吟TyY�+��K�k5(/���
}��&�j��o�{[]9{Zd[A>/x�����v� ��k���q�3�|���3������7M��w�2OPٯ7�:ΰ������h<�~I�N�|�m����h8��c<�ì<OY�q��'��w�OY
@�4i��1�[��^�����VEw��t;I�zɶz��VC�d����	�M�5�q�S�p:��('��8��M�	�Sgy��'����(�����R2>ȿ��Չ�ku���i!�?3L;��'�B��Ϩ�m�$=9���m��6�5d=a�M��OC}�8�	�^�d�O�:���s$?�ȱÆ��DTT�)���Kk�I|=�;;�h?�:β��!欟w�0�����ɶz��u���z�
��'���)'�7̓��>v{d�'-�li1���f������,�Q���	�伳����'NfI�>d<;��	����:�?&�ѐ>g����d�OQa�R$��[�$�|�%H��������oM�)5kV�߇��$��'�6�`v{��:�Ǭ���u0�p�ϐ�I���?3�&3��ߵ�O�T7�q��;�Oȡ5�3̏2=���;�/%]����e% '�-�z��9��ԓ��Փ�M�`n{C�3�|�}`VC��}��>d��@��:��1�fB|¡��dR}�2�y�}�K�Q��t!�	����*���Y8�����Om'��q�Mo��'��!��	��j��3�fY�C�x����oA�0��`i�@�7ܓ�m�e�~�4|���{睿ĕ��ڊ)'�l>����Ne�̟['���Rm��$���OY0٪N��=`Vq��éܡ�{ϸ�|�d�Y1��5����[G~Ͻ�6���d�LE���VN��:�N��)?5��^ ~a��'ڤ�ԛw/p'���C�6{Hxο|n�C|�/�]e�v��;�mL1{�~T��wޚ�1-��#�A���ɰ�-�QT匇�Ȋ�ڽ�d�s���MOCov��B�Q�}�A7�C&�nin�켽�}}��i����z��!�l{"`�Z�yp���t�yܓ.k~כ��������~fl���wrU��n��}�i��?�ڟ}��̌���'�XNRu'�1g)�V�VI����<$��2�+�&���G�>�꽐<ϼ9�p������2�nA�ƻk^��7�&π��G�>P�O�_��I��MO���N#�d��y�P<d�C]�Hu���5�Մ�&��OXNy��3�G�������f6���� ��I�������<a�M�䟘
V~I�NN}��N#�d�О�;�J��&Z`m�Xy�g�I:�����w}.�����o����Xb~d<N̰?!�=d��M���0�C�O��1���O=�zɤ�E�$�'<�!��&3|�>�x_�s� >E������N�����{�y�`Va�������=g�'ϓ,&��&��d�$����I�u	��&2qO6��:���	� ���>����m>��Z�ϧ�s����ī��ܗˈ��0�aD}�R8�$��w��dĞ��E	������ɶm���1��'�<�d�L���u���n{I�;i���{�jB�or��{O���a�{��=d?����?3L;�'��C��~�Rx��>a�'�����z�����=G��${��}�u���ϱ�����o���05lϩ8��N�l�rC��y�O�ROP��q���!�sR���0��0����E&��!X~C<g�vj���I2�����1��p��~�|<��>��Y&�w�{�;l���N��6��N�m8���q��p�\���	Ԟ�!�?2�s�'�2o��gY'�X
�����H���`.�aJ�bv��c������4����a�)$�&������$��'��N���C�8��M=N�d>Hu//�|��'{�q'�����T@���U��oEɩ�� Ճ�ACsy����V]�����%9��	�]{}�@�����h=vS����(Q��;g��a-w���;�]c�Ĉ�݁�tƔ�����]�^^��k?�]��%:�R��8m�+L�ˎ��p��:�3:K3���̱ևd��<%vr;4��x��Z��f?@D{�}�B`~T&���ԟ2z�(@��[�$�������g��$�����q��<gɳ���d:���?!�OXu�tf{����^�S��_o8��zχzL��i'�V<�
,��w�Y:�!��d�O�=�E�<`{���N06gp�~I8�j��������>F�a���>F���;Ż�^|< �{3���CH�rN!�Lgχ3u����pQd�CS�`�~�]�@�'�I�f�Xi7���7�	��N�����{Uj�sa��*��5ꟼ �q��u�ԓ�|���8�9�0�C�m�d:�l��6s�jC����h��u&�'��h޳�0��O5d��=g�hg���$s�>jL�_jg~���۲��O�t���=g�O�W�������:�l�{�m��<�2I�&"��su%I�k%Ւq�yE��#��ط�ݞY�sP��sF��aSԘ��hc;7���!�4��4È~��ì�M~�d�����oA�Y&;�Y=E���!Ԟ�e�ٮ`��� �S�o�y���+��%�2�<���ޔ������
��ѫ�������d<M'XC�==�1�����%d�����N&�0>>��{�_�sd �_*�J�&�>�cP���>@�9��'̞��&��N%`~Cl��Xq$��]�6�0���x�l�gR{<CGS�${�2�}���=u�o�k�4��6���q�1�\0�k��ʛYW-�\�8����
]�9u���V�}8�E,zi�̗�ր�hf��N�ݼ~�S"���J���u��B��h��Ye��.�ey5�g'�^Ԛ���Jth�|���g����Y$�@���ȰN��Y���=�W`�p����"��L�$xrs���E�<�����=sOV�K��:8�F�"��^�5��E�H�Õ��dj�6+��^u�W,%k�2N�bef���u��:�/�NZ�w1t�Z���Y��Q�F�ݬ����u�-c����}1�Bz��h)r���a�Ů���u�W�V�>�1�0�S�^Z8�d�0bޚ_�J�J���\�l��Ϋ��O��[�F�S@��ƅk�(F�Y���-��$�>�s�VK�9�h�z4���L{���"dWj��e&�%��ts^��c��#ӍtQ�Lve�[A?-������$���fE��E��У�;Yǖ�V�f�Z'���jX�`h�U}�a5�`�˒��TGiI�o7J�7W�r��vs��h�wR��: �%���S{��".�s1[��U�+�a5�Z�S`�:���;w��v'>���uY���=�w�Eѻ��P��jp�L�9�3�9�s��kb�� A�	7r�g9s)��Ke3(kn�oe��3l��]�J~�Qbb��~�ؐ,�oMkwha�w�z�-u�����z��8�Ȩ�G��*���3aC�Y��W�C1��MX��{�v! �w�oW%eCժ�%����L����s2]Z#M �x]'4s�z���$r���a�)=L��C��X�G/7�� ;wd������Cib�@�����3!X�x�H �E�c�4��CL����@��(��@٠��S�*!@\�98b�N�U��t�z`�nP��ss0q�����CW����;A��F�7�f��8x9ڀzK��P����2W*�p��q�$��̊�n�t1KR�!�e����	ɥ�{�f��n��D��ϐovP1쾳O�n�vڋ-��x��B��n!��ʸ�%uwP��6�!i�6�kE��&����0ܯ7F�|J��Z�s��3����j��-�rΊ�#�m��ҽ�7p�i�n��������33�T�锬�zW'Hٚ��͘���	�@^4�s�8��+jz�p
���l˥y_X�pǨ��V�J��~c �9���-]:���	�ۗ�.�ޏy�a򬑪��P�b1��z'0X�GtU��|�9-s�OJ�CHL=UY�t�]��TΎ�(eŹ@��!W1�p�SDB�3��a(Ó:�����o�L�$�-�
�7��⭠��xh�Щ�N��<ɕ2� @���Y��c-􅿱C:,\�/�KE
����C%`���!���fl�4�o"���j�X�-T�w݂���1$�eA�� L8pL��(�=�p����:T�I��j��ͻ�,�ڧ�o/j
4ȶ5�TPiB֪�m�Q�֍�mT��"���&+�J��\am��D�9sT�R���X�6TVح��-��Kh���IR�1h�f`�*�m+VZV����U�5j+iE�pT��Q��[J%����Q*�i[h*�-�F���QjRƥm�h�m����R�.4k��+��&R�J������aR����D�b�Q�kZʣmV�T�**��-U��Z"ն-�m(��j-K�2�lU�e�m��ѪʕV�Ѵ-�cJc�X�6��J���F�(�+J֊�t��ܦe��l[eRҔ���jZ2Ԫ�Q�ERƴU�Q�����-�-�U��h�F�T��UiJ�F����QjQ+Q��ks1�j��mm��T���(�*4�eeYh6�ƩQ[k+(�U�ŶU��WXb�[�����k�����M�xCDAԛ[���LLYn�U0�9z �o����X���Aoaj�7�]F�gd������R�����H�n�@fbE[�N����`7��8�� ,�t62���n����֮�Ws�bo4jF�[����+��ջ6�D�ȸ�^z���+��NB���=3Ll�c�#�����W��wD.ǒ�lU;�x�ܕq^�œyc��'�z�_�vH�C�3�i����v\��5��d������f0�wM�J(:�â�B,�d���x��'2dB���~�r��לz���y���4sy#Gx��T;=[ۣ��tQ��Ep6�����md杷����m��㺰U
������CD�}���N����f�w��N�_WJ{={B���:]m]&�gm�Ɏ�\o�E�FkU�H�Fcr�=�@�Zqo�m�Z��i���y-�����>�q�������u�R�o�z��]�/�=��˯F���y��c#�<O�1b�߭׬���A�1��Zq�{N�rS�Y����]��%��N.ɷ[�ɧ�s�u��GQ��[�ޮ�J��8\��>��w]��8+Bj�"Srs([s!߳�f�Ң׆���4���(Z��gm�����U���*8�.�O|���Ny��뼮����qɘ]4(�*�w/h�o&1s�d���<WX����lȅ���;Ҩ���O'7�q��)ꋊON{.�j}3OD!>AG�0g�<4Ѹ2��^�ڔ�h�^��l����`E����l*�v.�x��p[��3��i]� ��P��5 �홶�%�����u��Ѹ��C}�(e&tu��U��-ۗ�"�7����ɶ<��sns��rL�ɮ]�(H����jFx�deR�:�#��v�yL�bos%4m���e\��!�M�bfFkEP�DY��WM;�j'���e�����ˡ{��c��#�����x�E&�T�n���T��~�س�9�|�twu�mŉdt��6X��Q<���(�;R��~�g��J_=.[���7a^Ɩ�z��uK��n���~0A�#�ɓ˱F��*�ɛ��{���)ۀ,�-~��u;J�.����f�̛4�qY�60�v�#��Ԁ�W�X�Fr�Z([�7S�z���
��Xc���%�����Z�ݣ�:Kk�j�Y\w+
}�1t��������)�o2�љ ��uʧ����]P�=����1}Dѽv+�f��Z�k����,�в6���ҝn�1����۵�ND�qo)�����.��c��,L�~�*��Ib�`o���sK��s̽~Z�����F[��%t^Jڢ��Q�N��o�Z��M�^�Ǐ��/��A���Чп��Ӆdߖ�>�ru]��彙�*����L�5eӬ����c�7�3
L���\���w����D�(������/bi�Pj����q�� ��q�/�ě��~b�"�=����j��u�Ei��Zq��.�*r��rX�v�8��'�!Gf��f�HU[-�'�P��*�p�F_dZ�����خ�yJ*�^��j��.��Y����ܴMh�JC6�'&i���&�YqF�Ȯ鶡��F%6��8�9킼����z�}��5U��U�s�Y��={ui���oK��g�Ckj��ku"ض�5Z�rn�f)2u�}-34��zF3f�k��4�J���t�*�pр����fok��o��(����A{HMBeuf�?����T/8{���?9}C[w��{K췆�42+��V�>0L���s����%N_������?v�"�#��;^[j��ջ6�6�جq�u.zd]�Q�6�5�>�G��ѽt�j=m4奍�H����Z�·e�]6;���˷B�N��"����z1ڴ���й;��*"�\�
�c�oM�t�W+�,
A���:`�B���xB�g[��K:���)DsVOT�FUB�r��^�=��t񠼡��rz��{ޣ�����;���x����)�{�����oԶ��P�?,��r�Y��;xz	��ǀg7O���N�wX�K�5�n���j�K��^CL��ڌB]-��%���SԜF�X�mؗ��ʓ�H�P}-
aq�ٞ᥍��mN��U��Z#��Zr�\H�s�l�+�ld����zX�<�T������������n�u��O	��(�\.�4d0��Hg��ka�6�:�KG{C=�mh�z�i�N�:RpFH�l�mw���թ����u3}`)�S��)�i� ��kFWh鶱�_9W�G" �w�M����`�D���'~��<�����}~L��t�5��"杬2l.aM�C\i+�wk1���d�_��J:q������|�5MgVe��M����O"����i�����^	����;�@���G^T��9�>��^�+��%��^����T�uj��Q@,zhs{�Y��r��ͧ�t-=��j�ӊH���'�6�X�xج���9ʲ�םkwno������y[�"l�c�-�ʮ��"��_�
��{9#BVc��^��^�۳�EVlL�j�9Y�=�^u�@������ᎤC23]��W�,x*�Ɋ�\U�MO*Z�d��.�!c��#�}HtԦ{�.��5�l��/�_C���g�9�r�ܗ��)�}C���\oz��h��X���n���4�Ҝ=���9�oKo��a��|5�#��.�`�8&W{{����e���2�֩������
��-=���s,c�#�:�g���l�X�\i����M�v��Q�Eq%��[�u�{�F�
���]xPGoB&�c��o����^��#IM{w.i�=΃�[[��F���;�xx�u�,L�=l���E��N݆��i��T����[�A����u(/ӓ��oOǲ��5���^���뜭�5P)�MB":�;z{�a53��4	��C���x��[��ʢ�iŸ�n�:T��7YGݚMq�I�����2�Y�CK��9@ʹ����X����)r=j�UP�7y�fk=8(&�JfT�M
��8�.��S�VA�)K��9-��f��)�&=��4�>h��L�zg8N���)�YB��"�S���S�%��a/�.C��tv��sRxi�pd>%�/<xf��1���{���n���j�{.P��خ
/�E.O��e���D�X�����)%�﯌<a�;x6�U�t2���Zf{�N������h�(�ʇ-�5�����yӋ���Y�us�>���P�^6+5#Y��e��yl��U��j�	��>�%;�Χ�5Ǌ�f�=l�����%�Oux�������G<��_x��q���J���;r�
k�_��3��i˰�cc	��MrץY��K��t��w�gr�2F�"R6Y�Х�\Q9��]rވ�u�I�ݘ�XT�C��DZ������{����.�ʧ���ɋ�[�}��8�z+��z��rdRM�bf��x�Jɛ~+$��N��y�5�Iά+�d�G�f�?p/A�^a��Y.[�L�ֳ>���m:'c�n�I9T�	�o�\������m7o(��X�<5��u����L��Hb�v��M�Ev��b����-�Y�f����o�t ����i�P�\�OS�bY��z�Cn��F洱v�]}xv%�jW]�n�4�Bܮ�Q:Z�׳	�Z쌔.'�9����i꨽��0$6̌~���>r���ǔ�V�+�D�;�r��\�W��3X٭�6�j�I�q�)~ᅊ}��]P3�����@���̪�M�l���j���2pPI��A3I�ML�AETL䎰ob3m։f�5(Jz�jb��w����a"�
h�i��=.!K�ۛ�12�I��d�.	v�:V����`��66�/u�ܒ��DR�x�&X�5t*�U��a��w1[x��٥R���R�l�Gk	O�Y�32R�A�G�V�s�Sq�o�SV�_Ws�Eb�!��ԫ��0�C��⩹Z/o�x۶�sˊ4�5H-p�=��c�s�N�a�sU��cEr$%�+n�DCV��������t毓Q3����LoM�"�ӿh�$_)� �e�+
3խnOa7���w$�������"�w"�*r��1�!|�&����R�\�:�\�_-���J�4/�쵕uM��Bo{�嘢�ꛛ�o_*�]ʡ��y%�6&���3k.rdSyW(�8k\����[��V�"C�|�K�A�Ya�gZ�ݛ��¡�mWNL�>��Vä#8G�5s���E�f�#"W3��&���ɥ}���\@�m���Ǯ��fq�c����L��٦�V$f�ڱK�X�+��q㉩��wv�>f����}��k�ܫ-�������|�GV;U씭�Ї��2�<�4+S���>��s�wJ4��R8O��y�"B�>��S��v&��w�Sk�(��U����>�}qy`lp���l��])�|��)���G�K<�݂+�w.��ѱ��5���w�#X�������jM|$W5��c]g(�/����k{Gv�����q�J6�C�6`:�Ed*{�K4`HDg������[u���5?xnv+�s9O�:����~Hi�9{��ʼ{�Y��k�k�Q�{�
��;��_P�*:��Z�*S�
T!�����f��[�ө��傔���y�r���Ku䙭���g�Oj�4a�wݒm��LPaէ�����=.6�s>צzXT
xs��d����yws{��"�L��:*�Xm������J�r�4;c���4��yV�%UF�3���3�h&aMàtO+��(˕c�[�L֗GC;��+Cծ�g�h��>&=���(f��u�6�"V�嬾7���=S��i�������sĝ_{�Z�tG��> A$>C}�����WI�+��9���Z�z��]���/&~���^�������:��\�w<��yu]�^�BE�f����MW��5��yn�k�>�z��,��D���ᜉ�tme{7կ]��:},�f�CMNK�:tg����ӜV�z�c���jn�h*�4`����݄�E�ؐ��!���5�����ڱ�����L��zC/��lš��19Ff�١��M�f�Y�Y�����#����?O,�3�̤�V�&rfUoS��z��_��w (����z��k�s�亼�nͫ�HYA�V�"���V$K�J�kf��R�����WS�g%P�;tߵ%Ԥp����|%<�92^�;P��Lq�=��h������;��<Lz�k��1#�v��˷��Eu���-��󭯞NЅMX���_p\U�Z��6:e�P�!%93�XuY�S4�r�6�e�@��^$�VW����u����Aq���:�'���a1�ke�\���w*�_:�B�;&�t��#!Λʚ�0��ǵ'�9y]��L%�ެ��C�(�/�δȺt�S�$:��5�kM��� 8�T��� (˿n'��n�l���z�d���tQ�:��N,"�O��>)�t����o鋬�p�D{NyS&$wӥИ»��n�C�J�}!vZ��Qo��>Z±��龾*c�nmc�b��:Y�e���8�S���q��2תB�cѮ�CA��N6�wE��i���k����m���T��B��o̪%ϋ.�QT
��v'�D�9���9xS�4 �8�"�]�HB���$��MS���{��oz]Z����(әk4�C7�Z7q��7z�}�߅h�	�,�$�%:��0>x}O�q�dhN6����uݓ��lɵ�&?�[���)�-�7��21��xgHq�K���(N헇�/���phS\�v�eX[�|�.]�Խ@��ٲ���]q�漢�tS��Nh?DY����[���H�D<����־u=����GI�f}Jv�u�5����,0��,S$�9���F���ֈ�;|<��w�׾N�74�ɂ��5�h �3N���;HLD�K�A�z]�	�\��p��[���S^񶲋�L�\4h�1��Y����'���p=�R�����m5�.�;;�L�Ɔ��s�(�=�7z����&k�WS�1lPʺ%��d�]�JVӅ�F=�Ϸ��Guյr�y������Rﲳ�@9�|�h�U|�N�(3�#����>�B0z�J
6:fb� ��5��5�݅҆�Lof���0�pW]�`��I��9;�m	�l�S�V��5�:��|�Mm��qѓ�/�n���李������H�i�N�}�ۍ�s��xn�Be�f�o�.��.�.MЍ��e�{���诠�{;4�|{���a3 ʙ�2�)���}hk��k�]I�P�R��E-�
Ѯg[Z�w5os^�E�g�!X�/�Hl��+��
�YY�m���ح�n�5��Sְ�׳,Ts(�q�t�GrU��R�����Ǳ��� :�+zc��N<���b��j���hf��N��T~L1zTy���94�ScoT�e:�U�O�,���l�]�^�}�9�Y�v��W�k'ƻ��<8�]	�i����:8]Ź���� '��h�-hAwv)n��Y"�ws��u�bVF�Okz�̤̥B�F���Q�M�A��sKx'Ndu�>��v�� ��9���NE5�(i�j�s޻i.	/t�������<�!��8y57B���i���v�s����iY0�㐠m�&���Xu��5��5r��HD%W��9C7�%���of]>�w�u�����X�0��K���Z��ҟ.w�Gu��C+8���	p�/`���Bق���OW¼�<T;Q���?�^�y�r��o2�k����շ�n��E+�_�c��n�R��i�u�����ˬHGk/%4
F�Wh0�S�X �e��pߵ��tQ�h�t3��4�N5N�ĚZMJ������޴��֨�}%nJO�z�;�M�:�<���כיﯞ�Z)RڴE�V#mF�UB�5b�[q�L��q�"#�V�Ձmj�V����!F�"5kJ�Z�kc5�eimmD����`ڶ���-j+
%F-�)mE��VҡJE���mZ��Ҵ���+Q*��Tc�1r�mmmZZ%l%DV��me\����MJ�
)m�J�R��*�ŭH�\���1a��iKlT��X�Q����VVU��R����.%��J��eT�JYKKil��jQ�b�Z�,n�5�1��1T�e�r�E�"���9h�L-A�UV�amQ�(���5JP�6آ���0P�̉�kT�Z-��U��"�)Z-l-��2�TYj��km�+,ciUD�E��6�m�U��
�Qk�`�������Ⱥt�Z�ڢFZV�aF��
�j�-��Z����j��J�J�f�N�C�ED��#�����E%N_T
h��ǻ]c9.���a�\ȹ�r�o���w8�B�
㾙�:Y��q���*��)o�{�� D���l�ync�˨^y�\m(r$.�(*��_ܮ�%�{�!�|�PJy�����e>�N(^�Ծ�(��>��̷G�/`�Kx���I���s*q���785� �Yޝ�|����h�:���Y9T{�oBVf>6�z�y�mfH=�S�=z�>�[~��C�U��e>�`�{���F�W�WT�8b�|O.T/��Vk�{t�O��<�q�oϕars"�N���n0�J�b�MU�C���(l�v S�hNU��Tzb	C���δ�p�t_���;�;p!�N�YC=2����Dm���ETg�\���X^A!M�f0���ű/3�e%8�B"���m��WlX���Sǃ�㦅�S7�1�]�x�]JLh�.V�2��O���K��t��neV4z��텍!�hU��F�bT�UH�ӨP�2F║�]4_��`�ub��`��k��	>����P�}���m�iv*��q�z����W�����d���E�ɬ&��'A�h"���7��������D�򩨂�VJGS��h��i�e�.�̞ ��<|+-���އ�����G�b9:�u�fmrC�Uy�:����X�)�/�����"�9�k�צѲ���뢗1�
P�۠�_q��׆���]g7f{�o�ܔ9�s�B9o諭������knS��,�L}����m��"ÖbF: �C�D��%����_^�,wݛ��gb��kҶs���$���*��J�R��px�}��ߐ���芬�mI��z����e^�8�����,�`���Խ��r`�L�@�oa����֪*����W�����PXX�/<��%�{+>�(J1�BsG̪�ļ��ٻ�嵘��G媌W��,E�-0k{>Z��X6Y�4D�:	yX*�T�H�Wze��_7�7&��ʟF�y�M��^�Q�[�Q��er��H�`�OoH�;���t��;��37��e�<4Z]
\Ɗ����58ei������ʠȡ�T�X��|G;����J^�a\ �=8�\I����`q�M�����DwV-�e5��/�j�<�����t���䂑A��ґ�V�\�n���ǎޟmu��Ҵ�߽�e����l-����9���l�~x'�Z��d��F��_�J.Įx7=����n���m>�S�ͥf���"`��qP��W���r�N���`��� ��qyQۘ6�u9��y�*G��lg,58��q�'R�E��{��Y]�鳙X��yS�Z)녱Q���Ͼ��U�oaf6���c�uK�ˌ��4-��^�.!^�.#7�Y]S�T��^�#ہ�wiMi*�.�v�2a�r*8��mm����|�������>y��~�]�W���<�$��f��<�j8_��j��QX,�yU+�*�t+����u�����r��s3�=%�D���<t���n_��x/g�^yW�,���ƾ�$�.6u!��RB�ZG��\��Kո�a�����W���P�^���'�ʡF����P.-6�F=Z���99oS�8ŏ�|_����O�xO�x��Kt�q�*�J
b�~�T1���f�QȬ�Fk���J�@��v�+��{�+K��KY��³jz�����@���>���n��t�o,kp�%B�Ը���b�Ge���\��P�
{U��4_��Yo�$Chf ����0�Og��XoV:������/�W+%/-aq;o7��~��Z����=K*U����we��!s�f|�Ua�퇃�*�i��og{�ƙ���E�T혮�]V��J�93�&�4��{�!z��Wi���xNί��~93���k���F���;�����y<lbl�6�A�/��d���Oe�*�,�}W2竫5��"���E:���������ڽ��yv��g7�^���#�6r�����{�2��ѳ"����[BP�ᢜdE4gSj��C=Tz���vJ��畷�Z�g�${o1oU�o/�6c������A�k<��k?�
խ�/������c��>� K�{�8r�M�����}C/,lYd���ۼ�o��t=�v�c�g��^j˙�X��3��/�
v~�n�,5��NV���h����$���g��W�yN�d#���'��x(Z%o�(���8�8ϒ�����bG�!���˷^�hS�zy�W��ɷ��9݊����2\YS�H��x�(l���rvq�_�v�æ�8t�_>��1!���w��LďyД.�ѓ(��(O����6�zs��6�!S�)El ��t>R�J��?K�5�BPz�/����kٷ������cI��E��3�k���[+�m!���<y[4��:;��[��_�K�h5���;\a�/ST�-�\�gn�X�u^�9�S�����=&�~����GU5V:�]�����*�S�_{/��[��+�u�(X�8'>�]���fЁ�u�P�55 2���B�{�z��3��x"���ˣ��r�u9����5 <jb��ؒk`�}�ɍ]H�A�(��Fu�[�ъ����<=U6�)���b¤G��D�PV��?n�0C��5���0&=e�L[���H�ۥ|)G���o���qh&j�;��^|���!^|�^r<:�S<.J�T���jx�N�ƣ�lIL��� ����:衵*���U]�W6��u�P`����mp�I�s+� �xn{r��xc�Q���Cy��݂�x�Oh6%�-S�
/��j-��oh��"k1^�u�1]��Q��,��x[�F�&�<�&X�I��IS���iP�Z7=�2��KG�g�x���%��`�R�>���X�6�3-1�x����ar*�"����v�\���z[�L���8���@���xDp	mP���f��"�aw�M�Y8[�ْmz���B��Yj�N�+,5d���z��*6��2;D����h��p�d�}9�5q}ָ��D�� s�5窰�{������B��J�5���z�h���#-��۞��u�γ�F�Q*�����K(�����J��	�Ja��������M�����ϵ�z_U����Cr!#��Yޏ�V�ܗ��"t��H��������.����.v����wv�,�s��D����Tc]ON}uA��>c}��|���s��ԥ�=�ӫ�
�9y����m�U��+v� ��A��@�<����;q�)�3�%U#�c�o}���yV���+�:�8~X%�N�pщ�E�.���g}�K(�!Hr0��]Cla��w��$ǘ3���]	iӟzUq����+"�5�U����s��8�ؕ7�b�Y7,fyS���&�
⹥��m{�W���iL�B\ڇ�t�j�XjP�]8޹�T�˭֧�-ŕ�-��KjL_|�P��z�m�%تk|����"��vվ�5#%K�U)o+S̿.|�&�f�:۫2/��1>�Dk�C,����]���������V���H��d�����T��Y{�����2���_����_өa/㽴-y\��d�9�[�$�����W[jr�ǡx{��/z�J�ӄA�3���WT(�[�k[ȭ��$�w���D7�Z�l�cм���K��=+���Y^Ut�8�k f���fP~�����b�m�e�e%���~_M`�p�8�`���%Ȏ,�K�('��g]��cz�!�ћ���BZd=I�p�ko�z�|�W�H��0X�SW�Jd�\��o/nG8��D��N@��ٖ4U���&Ga�mrL!znJc@����	�bl�a�8�.-��~}5��;�嶵3��r��F�
&�V���Z�IdP��
�����<FQ�`��v���V�'��q&��Y�@���Wu�{��ZR��/βU�׮�w�D2�9��;Z�j�X�xT�^�y3��+5_�a��9"�`E��2�׮��w�h��3A��p���Q�������x\PƼe�[Ӻ�U�F�\���b >�ĵ��tʨ�cP9�ܪ�Q��%�ƭ��e�s#JFB.�+^��_E�T;�U�יݷԼ]��fzo2���|�������V��j\B��ˈ��"ʺU�X����yՏ�]��Sخ8�[��[aP��,���5���
��˒�_\w�.p�fMyV��Q�a�ؽ��I�/�o�__T$aP�g�U(t��WT��l\���싲�+�^���zU^r�&j���MT;ͫ�N]#/<����� �G��
x�J;b��l�Z���]&^=h���欻�t��,����u�C�xE���p���>4�=�����
fޝ��KS��Ga�8)�G���g���s).��T�:Jb>^�T������v���6^`i�AX��z�����I����܂@���;�+eʱ�3T�����ΉVh�<
=$/�Q�7�5-�ͮ&a��ӖH�uj=�S�)T��N�}��^0.2�6������ق�����z����ʩ�I���V�o�	| � {�b�Zڌ���c�]G�B�o����=
�H���2��LOS�YFp@�OZ7骥λ/3[Ck��0�Tf�$%D2��F�Ӝ3^�|,P¸���o���|i;a'�[:�����i`/�zQ�o�G	5*Y�&$KY�1�j���P��c��r+�B�z��0�][�Nt�&.�1.P(Ѕ*����%Gy#����<��^
|Vh�P��7<�����	.�C�1]-�X1;�)���qvn�7Ȣ�>��U��1�y&9߽�=(���'�Ŧ̿zz��U��"B�_ٛ=a�g���l�hD[�M�
ӟCs��_j��
>Y�8t�gV��@�͖X��	85x��^`v��t���}�6�n+޹��-ٽ�����y��R����>�|;����C��n��r�p�GB��մ����[�gy�e9��P�(J�xQ�[Hp#/��~}�!��&}��C����[z�a�����0�J��λ���e �S:l���!�4��t&�S}���r�s3f��X�"!��53��Uq��V����f$2�*��;$�����X�-c�`���+�Qk�J�NL��]5k۱t�^�� ˊ�J��*��v5�&v�j�x�dT�B?Vk�7�b.�^.�Rn�mDp�� ��*o\�5}ڙ�0�i�Vk�u�E�%�[8���I�\�\jP|���:|.�U5�֎���3���H�,>��y	�uj��҄��%SqPĨ^��J���u/�/`���<�*Mp���|+á���&υr5�r��1�����s��y;�i(Ϩo�z�i�G�����t�9-��O,���Q����uz�x�ڛ��@}���r"��21��Tt��.�^�`�:l3�Q��+^��n�Eo�[F8b��d���A���u�}�%G���U��P�2:��Z���9\DG_�Ozͻ������n����H���yB��W?�se����N��˕�Gl�9�ܻ��Mv-0X���R:0�݁��Ұ
��}�
,>�L�j�
������M_&��9��k�c�u��e��f�\�>!v�AWw� ׻ǜJ��`�~>o�Fп�x�xwi/��'��<���LuLV<=S�@y_6(�<H�G�f.�vإj���䇝�1j*��V E�mfU��%�ˣni�8���/x7��[з�ot�a�;GZ�|�$�⤞S�[��Z���'B�n%=�|k�dT@3�*��hӷ��pN�{�k�YW���Pr�2ڧ�um�l��W������W]��e_{��Ny�SC��#��p�dn/r�܊�<�Ł0���b�&iEN����ghg�i[�������,3^�v/>�p�hz�V�Ѿ�]�,���������+%Pi�..��w�G�i|����[�Y�U�g�K8���V���Z㡊������Ċ/�P#�lǵ��Q��'�w��^x��*��i�boa7�v�-	���s�d�*�-6`��פ�:�����E�pp�[<�RP�!���>����PsY�mL��P��9���O<�	Kˉ��8r>��-�<Q{p9���U�]�F�{�粶��\��+�P�j�m��C�T��\ڇ�(��R�9���v*Վ��O�oݩ�~��y�j����İ�}���`k��U��b��ƞ�EJ�{��B�Ek��wݜ�c>�x����������`��R2=������gbc��W9�[wp{f Y�����g�Q��?�������P�	J��?�WL䞰�3V�]�Si����m�tvm�����{z�ЇV�*�iD�t�jY�G2[s������2>�Л�hqن�b\r=�I~�}W�/��؟]�utz!��7��7	Va���wm,i)j<9v')kiy������"r� ��6��k�}��z�P���D5S�"��V0�U�ڻ��ݎ��xkIkZ&{�`���m��<&��sZH�b�V�f�����t�&.61��ʚ0U�N�7Rd;]q�}��9�`}�Դa�A����JL����5�Iދ0oC[���,^�[�E��#W��F�v��s�jQ�V�aIL�z�]8��T	��(Q�`Ѓ'kd�&�3Cj�*�׵"�Պtv�*vy��r���Қ�o��������iWrц�ɼ��s\�i2kx�� �j+�Ʊm�3lA1Y롧3�N�Kzf3t��kf9�`�t����䋜 �����}�z�[}�4M4�j����ښەܙl�)��]�N�aI*i�+��I�kz��;1�b�"?vr�ՠ�y}V����I.֧��V�[�|ۉ���f
�Hhw�#Z"��ܭ�5s4J�%�n1l�aN������s��3Y�A��ǖ]9]�||q��8
qT�"'�Cva�����x�'���O��.EBn�ȏ�/I�m���g�g�#��������f��,��*�t�T����<t$IU����ů-��lj3�z|h�	L�0�ِ�}�(i����-�5R��t�3�
Un�w9e���s�Sx�fS�D�.�$/���R��X<=�\�_e�)%rx5�vq��ZE��k�5kJ���I*��4��#=x�T�u7�!��׭�&����nĮO\� �%0Z���Cdk���C5���!�o6k�R�
Yq��A��&�+�>m{���2�t
cq� �`#�$9�q��{�{��9����WIzP�9)B�^C���OD� ����9xC�D��O�r��Q����@�ط���%���n|�l����rw�Jq���:�ѻ�� ��[x:�L�X7�6��o}�)EV^"����n�3C{f�.�J[29P�7��;�!Y�p�د��Z�P�M�}������6F�#+Tۥ��r]����w'a]omZ��[y�fV��4@�T;7�E(�ې��F0�ra����^�2��u�n.���^iاQ�^�S����9>9�e0�<}�+�Qm.�;pA�$�3a(��@{]`[8�ư\��&Rk������丼J�_Q�,��zn�4:V�=�F:�ܭ�'�M�o�}7��F㇢�@\]%�c�x�k]�y˗Td���� ��ǡ���!y+S�{mR(��X	X��HQ�X�(�A/��]"�g2��]�VNn 3��gkɕ"�ͫ4�s���hCv�	O�,��!9Yvk)o���]�1�7��L�o�=��� `5F��V�&"bVVUm�k���Qf8�J(�mieA��
&8�e��*U)b�\n)\L�qrҵ�[Z"��;k��kX��X�U���Ҩ�Ѣj�m��X���T�%m+R�D��������Ykh�V�X��TYif%̲�aQR�h�q���ґkTH��H���ʩX��,Z�De,�
�Y[%��*���Z"ڍ�ZZ�Lh�*�Uf5������b�RT�eF�ADV
��(�!mjKF�F�UKFڨ(�Z��1m���V҅�Q��	A�F�֌ehʔ�TV�X�D�("[m
Z4
���DB�jFLi�Dm�-iUQb֠�E�1�r��b��[K�$b$[K[K"(��DX����EQKiK
�+�+QE"�������(!i(�KbZUQ��F�UUT�)ZG)X*�����Aڭj1DFڍr�V��-b(T��1E,PV�� P 
_l�2]q�P��ڜOc�m�x2UD��r,�(�-���ugA�{��
��}��Xm7�fjؘ�Y����ewK���Iŭw����es�+b�ҫ����	oG�K�J^��*���G[��r��l	
9yݽv��GPvp�W�^Z�8)����lzUuA�<c4	5�W��M�C;U���좈��yi.�S|%�0��-�>_O���x��P��%�M&D�}�r޼�4�D���nJ��4S��AȽp�ko��������3��|f���g.�[�q��W����>�	�%��
�O�k ��I�46�����n:��N{��]�ؘ��\�H�ڦ�p�.,�Υq'òVj����f�a^Up�X�[kϳ��� �j���}�Z��"�e��I�g�>��
/�լ=�� �R�7�69wW�#��U��荚�M �OGυİ!�ih�>�,��gp+�"��!�{0�n;Զ��㥽�%h�k�of����Y_y��a�z��h�>'�%�^�"ʰ)Wsk�A�ǭ���YY�ΙKl܉�.6dV�O���6"����U��z}˒�ř��[�7�ۣ�9n������ �Q�w�N��WV�7��#�F�!�!ƞ.�]�� X�5��O�v�Y&��L^W�U�s�����^ؤ�!د�n�eL��ǝ��f���B�Qu���g[[j�:��`.r��E�oS[�lvÃT�������ުK��ͷ̛�۽�G�3�~�}����uC�tO_.�Z�1`�q�t7�LwWco5�c����}�Y��5p}/7�ϣ����qU��0р�/�}ZI��D����ޞGR���U�O_N��YM�B�/��ȕ��0dc���;~1Dq�ñ�Q���KX�J�Y��_F�Q�1�f{խg�x��O*��錧�Я����8�Pn7;w؝2}W�{KI���g�	�f��~��6�\i��L�����p�?]U%+>���5�>�Ȁh	�QHL�B����	s����b�+����t���s[��Z�^1q���8��� 5��_0�z|6��]ii��*�T��,�ޑs���O*q$2\=�0�%PS� <h.�ixN.�U(B��f�����fDn��SN��Rrnw��[�.�3����ƛ8�������N+�տM�(�g���Q�o���Γ���Pק o�g�]C���T>�uX����eVs�ak���(Ç*�G=y��H�|�������,�TÀe���k\1`ͼ����8ݺ^���~߆�	u����݀s�?{�x��Q�����W���_!xp/���`\X��Ε:��h����y��oA����Pzu���>�էe�� S�cm<������H�_^/m�U��;9t���T0X߮�>�_���4����i�I��$�3{x��|�\tdj|=ċ~�d*�Ţ�>"ک�O����%���φ^�Y�[5t��Q:�k���}K!�wE;V/�;4���)����P�T��CF:~��gq��?B ή�i��{5��������B]a�4�i;J+E�eS�1B��洄��HeN�k�W19��H�`k�N"�J8���,З���2;�u*FW��p��:�s�=��GEGn�:��t12���!|d*�q�k��ʄ��PЍ�xb��x��1�T)�㻚���13={��e
�(���T��Q�:��ʸ���@Y��✻����0�'���IrU�bf7�U��J´��i�փ��Ǭ�������s�E�գ]�>�)��,�lMd[R�H��ȑ��\:8P��K�s����k7_n�����J�U�.rF�s��_�U�ě:<,P��*���J8P�OU�x����RV��@W�6%�c�t�[����qT�ӒFvN+7��TuS=4^�\ ���W>~o?�$f��{O��kݫ��q{�L�N��;�hN�;��9���FD+=Z��x���-Z�Oy�R�}&)v�
���).�Y+j�y1'f�Nw�� J}�gr޶wp������ER��>٦���\E��T�O�TT#n�X�/�t��}.h-U��uG�)�mW�鯬s�����a$��;ǥ`>e��(����}ö�=�c��&+��m��ܤoەL��I2�-�!1�%OL�~�J�_�y��f��j�J}��"��/C��+�֗��r�<_��Lua��ժI|�E]�sL_e1sT�[��"��({�Y��Nh��i���p��!�{i�e��1��w�Y��J;A�+e��b��{p�~�«��Ȝ"���ֆ�v���J��3Pz�#�P��*�����b7�poTޥ8x����,��W��#�4�Sdp{�����m�g���,�ʕ�O��sFѼ�ϸ���XcMy@Fվ�W�d\�V�+rU����s�wg�H5���.������v�3��^KF��-��k�_N&]����JŌ�S))b�UE��J��ԛ�{\D��u
��ugFze5n��*!X�Q�b�p�>�/ ����z��J���F<�B�Sj�0D_=Ǎ>�)�6Q��7�^C-ADv-�g�g@��@�TL=��>�31�Kw(��:mZU�R�9��{1�����{�����P���)����6u!�
k�WaU���V�ŗ���M���{�"�ӝ�I��ß �wS����G�Xo�`6�Vs|���t1L.M���<m'��u��'NKp��]�}��`ڪ��<`�c_}��}������K�{[��X��[{'�:��S�,Ă�k� ��[�����s���GE�
U�D7�P櫾�����a�㼎�&&6�6m#%ެ��Z�9�W�޳>���Oρ �h[���o^<�5�iq��[B� o�;c�.�-������J�{�ɍ��z�f�0>��{jl��%v �ĴJ�r�X��T~/,�|pˊ�<b���y��拫�yO�֮a����U#�>P�
�M�2�����q����(D�ɗs��r�+�q��r�"�3�)���<x:�����Tb��W/l�{�`�C�y�S��������__��<a��HhY~�e1�~E�������a��� 6e9壨���'�겍��CPy^��	]�y�����	�D^30q��]Zf��
ŋ�!�3Yj���ꀹ{*#`v�k�Q,��qS���Pt�����'��q�k dVI5�0�����tq��&M�����!�%d��z/Fk"~]���{R��m�a��Ы�[��X�>�6e4��7sjܡ���w��iM�f����������W3s=|�ō��T骸TΘb��B�G͊�F8nfη5��M�6����w:��.T&��/i5G܄MC�q��*�Ѵ#��ܰkٲ�8t�c�)Eؕ��왬�v�tb&���rR4�R���8�hu��dPml7�OS�Դ8�������U5T���j�a�����,:��݌�Z�(�&+�á�9ر��c�Lv�lN��N\O	����e�|/�����J[�M1�o��b9��S9>*�S'��J��߈G/�X�(ܦ�rMhw}�e�@�ZVG�(o��?gݛ׎6�;F^�F'Y�P,7�Y,Z(+U��7�ޭ�#tT���l-hq��ì
{�y�K�DWsԩ=q=�E3�!���b���o��W�RAj���Ak�@�(c[��E�p%b�r���k�F2��+��k=�S���Խ>P��ī�+��\vk(��Ьt5����`=3�z�se�+u�{rl��Y�W��Q�48Us	�{�i>��g~V���X��q�Z�y?��ύ���\T,k��O�.��Q����ҁ�k�����^����<Ct=��=m'�t���/�+�.��n���ɳr���9z��s�ʰ�v�����ՑN�ܮւ�T͡�s�Q�L^ 4u*�f,_��ꬌ�X�w�=�٭��4���6�t�p�R���\�\�>�&*��Zq7ʼ�~�u�y�5�on�B���Y_N�W!�k�Z^��_�xR���<!�o#�̝D���y5[2Bu㔡Uj��:+���k'��� w�Ľ�[�u�EX;�IW���o"]��n��+�}�v+)9.Y�ܻ`��t�*�s�c���%����s֝��~��p�2�ٱo*��f:�yR��f�,X���<h��6���J�'��Mu���uC��R�9��8�T���T[<E�x-��IZ|.�W��J��]�Y�T�\�u,g7�~�	c۪�=羾^���λ����i��,��]v(���@������8�E�,��kC��E�K�ކm�h�s�Y�iZ8��tV�zm���/UhT���-�rO%+�tx'����n,��fGc���x'\"�r�x27blo+Fl;�����\�+p���n����kwG _OV�3�n �8%q��C6��WӞ\d:��Y��^}���a��*�;���:u�"Ю4��o�M���[Z�in����*w&^J"����nrb	�L&:�r=-�1T�Ɩ�a�z�|u�{\�K�X�O]0�^m䢮��T��#�� �6wv��+.��]Di�����p��[��1a�6X��>8��p��7�4N��Ҕ��3�M�PP��uх�B!�+����¡І�7�/�ch\�ЎWJ�X$�MPWJKa�.ׂ����w�߮��μ�噙��N^����-�7"/�C>b{�Ć|=]�ĭs��"U�z��u/ʃ��/	��*ߺM4�Z`�0�{�G�������s�xX�|S��+��zUǧ�����[ٛ1=�l�s�)M��~=,��v���D㑑x�E	��8z+->�W6�⼼2���?s�)��nt$#�`oR�V�x�Y��b-=��Kx!���V�Z�}v�gj�z�@λ�.e�EҰϖ�Dw��+�pƫ�u��-�RƲ\
��wB�z��b��=*��D^lw�nE;�u�O���Ґ�l��:�侯-�ڌ5v�g�$�C'K,L�N�U�ǻ�N1��dE�J��U�S�L�=����Q�J�s�{�u�K�=)�8�5r��4'��6^�T�&��æ�OZ��aJ��y�NB�FV�/Rط�l�j!ZS�4(:�hJM��^�ۤe=���Ə�)�i���X�`��EՇ{�n�̱\�d���ںL<M[�y.Z��0\~���!E����1��H>���Q�/kW��D*Ru�[J����eOX��V
[����^������:�(Lc��"�U"��m4�H��̊�T�m�g#N�+a�]�Ry��b�/]`B��.�u:j�
j�;!3�
%Wv{��eЀz��7b��C(�y��"��7�c�U�&Q�V��[�GP�H����8"�^,d����鲪�(um��JX�,�E�r6�P����Έ0���D+dY�X�C�Ԯ��\g��7�d_�X���u�.K���JP����Vo�����Aޗ��I٫e׷b�E=�*�o �DA���,����M��a[�>�_h!r�J��.~a���Jl��N]�qaŨ�t�6!ǫu+ɊU3��mՙ!�c�Q��I#�7�c�v�\�)�3���@�?:�u6d�}z��h�䟍O��ɰ�w�U:f������hSŭ(�n4�tk\�>"k||�e՗�*PĶa��U���Qu���E;�������ݝ�OS��e�6xb�iD.Z����м��E(tlzT�Et49���~����@+�=h�1T����+E��#}֞D��ݓG|ˑ����W����B,W�����pa�R�!q��쏳��Q���C��"�����=�j]G��#�o6�y����.�)ଊ�St5Q9�xz���9�{&W�����揙Zy%��?����%�Y���9Ƙ�^'�M��L%�rͬ
���+��Pqg�e��I�15"�N��<3Zᶶ���Q���*k�ea���Ũ�w�P#�GxQ�r��=�RfP�T'<\�Vu�6gzX!YU��S���ϟ�ҟ�_�7�B�����>�pX�X����4ߎm��3�Ɣ�ᔂ�ݮ�Aco,�ks�ߩ���WPugxO�J���R��	�Y���]Iv;����`��ې|��>Xx�P��|��5t�ca�d\j�b�Qeu�Ӻ�HCo��}��Y9C��W�~z�wT����������p��éԴN>'�����;ϳ����ືscL3�ޜ�^�/KP�x��6C�ʅ4�=
���i�d�F[��^�;��z\^gb�~���fO<�.R,�t�*��qFXڣ��X9^��{|�]mb9&�S�XˆU�*�B:��c�s�W�o^(���2�E#��,�:�{���
�\���pK&���<��F�E�X��
�=�%t�Ln��$�a���@ .���.EW�Y�E�Q�h�<��Mup4ŷ��]�YD撐p���q��띃b�d�������zY����p14�S���Xk�k�:��\/7���T�@�ݝ��<+���9�vtW�����^��u=/��㝎�:��3�YCk�ۜP ��\;F�vP�-nЛ�M��ab�k7ڝŪM�����J۾ݝC��5}6�v��������R􅲵n�ɔ�	P.w�fvg���x][#�\ؾy�p��:�e�+����;���0��;��FV���V"Nus�ȫnZ�t%9O�:���2EЁ��:_2���%�a�}Ɩp��Xܙi�R�a�4a{�oy��kh5Z�XN��*�#oK1���8(v�>9����]q��u`���o�n�h<�w��ñtqgoT,��N�/�	F�qؾ���3��V�]I���J;�����9��\��1fj'f�{�lr�u9;I≲9կnV��"�y\�z�xE���������*�`��r�|���ž�@�g�=����i·:��n����^NY�K_���g7����]L���wm��G/S��v���Ϣ�HQ!M�ux�����ץ����v��;ڰ��L�-:`f�HY���R��1S��V�|R��Y�L�=��Ïz�����GB�I[��m���N|�w.v⭗]��a7(`GݬOc��h�-���q����L+���B}���G�+���ʴ%�m�d��㱱y��٩�Wb�y�5�MV7j&s;�.=En�J��2��S6%����Ǘ� �Ui��`�a]��z&��� g�]w�E����mS����3ճ2눽x�ɱ-�T���Mv�"��	�fP; �ˮh�Un�x(c���%�p��P�|�_oSL����n��ث3��|$���\��ߎo���(��GW.^\ @\���O�f�x���g�t�l@�����.��Q�=b��>�.8q�+�zX�ؑ��O!L>_^Z�"��c�;�,���r���l�#���ў,���^�F&��^��>�z�=<�1���dG;���;�jE䬼����1���4����r��|�<��9��UVl������$F�@eR�
����a���u6�f��6�u��԰dNl�2C3k�]Wg�V��M:�4�Y��Ks3����'��c]��Q�V-�e��i���G	�އ�.��5��c}t��}�d�� ��#�a�y����N�]��8@�]��T�N��M� ���Sw����t-:ݳ����2($_�wq�+�oѝ��ܱL���H�v��Q�Dav�r��Ȫ�k'v�e.{oT�,%og�Hj���uz�A�{��o�ۀ���X�~���n�Z�qf��t�I�	o>ƶʘ����=�+�rd�8���=)��<47��]A��埝f�M����E��y�4���K5�X�j�P���ĉie�DQ`��ZԬ�P��2�� �`(��D�PTUF*j�UQ-�cZ*VJ�R�@P��Q-�`�Ȫ((�)v�4���Eb�Z�DU�ej�(ʔX��Ԣ��[lTY
ZT�E�m��cKK+V"21" �%���Ԭ@D-*�Qb�Is1U2Ѷ��(��UKeb1Y�QQTUUX�1F
�V*�,QPQ-���Q�kDU�)PPR*��(�Ub�EE(�DUb�KlDTjfB�V�X�J"(�
�QE�(�""��b�1ŋ��,V)R4�*��X����m�֭�ETU�
�X9h(���屶��QX"��EQUPm*�ED�(��R1X�
"1b�Z�� ����EUX���F*��(�(����U�����UQb������Tb �b,m(���PA�DE��E��KA��Q*QU��R-k-����V(�(0�|1���g���12m`ﯗ[�=�����W������$Nz�z�M�˓:<�F���޹hs*M<W���/z�\���f��*v��b #��B5.���]W�~�T�����83�ўprN�k���#�G��nwH�z����u-%�etupg�Қ�9>K�_���*!�1�K����A�y�Ns��em���2��(D�	>p���/8��YQ��(q�!�}u���/n��&yx�b(|����>P���]<k�X�{i(�Np���M��m�gdL
����i��-=Vp�Sj�<9C`��$�\���V��Wm%���rXS!�z���z̰�2+*�[���$ <mwObW�vZ�B��0��P��=��l.ޗ�w�(����F�b�~�`uBb�\=��O��)���qvn�s��_�����:�ΙՈ��0��u�Xomg��]J��-�
^,��\�9J�铴T���n��Ԥ��s7�7�����b���u��T�hf�,^�Ix�ZT\��Wv�ԧ��K���^�M��U����^ɣȰ;��^"�b��>�|���}��?�Pi���N&J1c�*{F*4y���eht��E�Wx<æ��ɼ;o42��J˻A9��E�,�,y>��x�G�;��"X�Nr��
�[�ꭕaye���V�X��x\DItR�;��]�WMX��w������ +�x�Ud��Ǽ���T���N�*e�\9�2�֙��*���Y�V�+k�l&���&��.����e��*�OP"�s��X��W�K8�ݢ��]iy�\P|뺧	eX���T��c��o)��nG�GH�W4�
��DW�J8�Y@e>X�#�'�u�,�u7�τu6�rH��͠�|p_�Q�2G�\`+�jp�����!Ї�Yl �h�t��p����"9�b�DP�:��BP4��;e�4-U#~E�)��ҍxu����-�hM:�q���X��n+ˆ�C��D��@b��.�،�M�*Y�}6B��e�5�U�w
{jf�{W3^B�V�f���7��H܈����)8`o��^�`���1C��RH���u¯�r�����^�ު�^r����3�У�u��b���H�j�Ak�u��8<7^ZC��Cሐث�PʑC�*��Yj���Q�W���gm�:��!�d�NKx!��(۸~́]
|u��{�2����FOv
���ϋ+�(��y7+N�k�qnCCm;+d栊]d�����+0�n������\��j�7�7�+q���I%�5�"��l�4E�~�˙�u3q[�:�7�R&z[�k���^(H�B�t�1�fޅ�w�7�hR�t�6Rqbs�y�}�R����
���A��v�.MP˷�M'���F�V�Q7r�4�������Ng2�{������}�1+h�^��<<�W�������
47wz�ʊ?m�|�z�wfo�XS�UѫM*KE�e�;J���_K.�N6O)�+-1���U�� p��'.���a(=�{�~I���[[�8�1!��^(��f�6��8\ei���<>���?uK�=�-�,��*E׆�wa����yl�.W��9�`��!����x�P~S;�ٞ�mY��x���g0k6QQ*���yƗ�l��9�Kܫ�n�wdņ��+|;ٙ�{�qc���m`s�W�`��b�@��
.��4'��9��6v�)���g�JC\ru������Ŧ&�[�Vtd�:h[��;}����+���q�x���v���$����R5F/p��RR�!�)�P�ؾ�Vtg�Q�^�qHۅ�l�(�ށ|C�'�=9�jɛA5�"{��o���B'�z��V��Y�uW��/�CHQ�Ð���x�|Hn;7Z)Y�`�޵�gn*a�1�������W��&�aWY�2d��e�qcsC�[�J��,}TC��u�u䱩��}�2���k�]*��E���M����JK��?�ǯ�
Е`*	a��,�.��-3"��ݜT��T*�v�Ҿ�)���3�T����R74�E���W�?�~�������),E}~b�����9��ˆZ`�I������lq!��0�:v��#W׶���;�/*��~5���;S��T��>ŧ�K���8<T�XK���+�#tc��+o���wԟ�NО��zl�5U��u�\��Uh0d�X��c-�����KJ!rև��/<��2\X�nOyu�UnZ��w����aߌb��H�*���
�|�?b�i��|�/��Y��]��
>��*�[�oJ8d�C���*%W�0T�,�+���S�2�>��p�]x���$�嵗4+�fo��A�|���,�Z��{Sɟ}�J��ǋ�&�)���2WteJz9f���TMsID��:��͛�t6�23fP:21��^�R����6GF�@"I��]��x�z< ���Š�X�G������+ �pya�|+|./E)Y���8�U�q������<������N�[��i��뫎^
�4kք���5ᑥ#����sW�كpգC�"R�(����3pk��,1޻��˞�������9wxX��Uh���Q^8����i��܋��f�/d�����)]���ؾ�}�]D���XR�wL��mډ[����Բ�	[^�H�ݫ�9=Py�ȁ{[��dbS	ֻ��#���9ST;�˱S��r�[����[�oS�Դ?�/�I�ۇ�w6���ײ�V3IO�c燱��/KP��v��C�P����,���z�٢Ϯ���[���K/َ,k�l��E��E��j��S%D0Y��<#�'��n	�8#�J�y^.HY�����k����J'�U�y/�ys�u��.Vq���y�Rvf� ���/��$��ֵ�ƥ�XYS�Ӫ����mй���T�{ӥ�,�gH�{�%��ce�߱���>� �\Xux��$��C:��? ���lp�!���u;�e���x�����z&=]CR�'���C�+K��XP⪞�c���j(��J��o�+Jӡs��>�R�|+�!O�*�Qt;�.�Cu�bqix�m�}j<��}~�H�YaT�q}Y����L~�T�c� ˗�kנ�pd����-�or������O4�˭����%)��"�1�K�Z^���b��c)u+3�WCX�R8�}HQ�N�DwA���q���րs� �`��K�|3�ŉ�l��pף�%���^T�u{�/�Q����\� Y�\mxv���m��=×$��m>Գ���ò�E���}[Cy�>�)+3}ֈ���SP���.a�O^^n3g�

�2�omg�8qק�!�lC��<�X\L^�H�=�4M���8�掕i�D������U瀅Ca��]a����o�������=~��g�#8���u��Γޏ�rֺ�M�j^Y�t�&���ݢ�b/���aӑ����}{,�q2��9�����N�3ٮ��d�j��N�1&0�F����zG�x�i�������V�]�i9�]5x� ��������,��w�Sݨrk�-<&��Ur�
�8�
j�6 ��x$���rj��n���F�+/��8���omcھae��Y����(��K̃�Q��ڲ�E��yQZ���b�cM����_>8�YE�|��7baPx���2ٕ�EB6�J��GF	�v��������)EtXZd4�!0!�V�WJ��[=n̩U�)e�I�hʇ�Pp��8�/s|",h����2-�/��jMo��e�rٝH�L�y�q	HC�nDV?HU�WN]#�9�vT���T$ĕ��S(݂�Zr�0�8VY3|27^���^��.xћ��u8]xME�fkL�ꜷ�3��ul�Ϛ�C_��^��-��T�� ؜�i�)�Z�#�$���u��K:�6c2f�Q��Jj�n��Nm���]�����{�q��^�W����b.V�����G�L3{���3";S1�	��f8wK�b#���8筇��b�����25��'K�I�z��A����d��ypU9<&�2r���7<`�2���<
����!$;r����/�M���*�^�0d�e��cgO��T"��ʇ	!X�B�}�^�Q�)�4z+-V�G�3�X轞1ɯwܝ���!�v��u�^��2�磨����a$��;g���}]��W.��뷽�l$�g�K(��J�L�	����mq�Vy�'��p,�]��br'������In�]-0��D��"�|�i^�K�e�'y[����Y0�w�Nef%�'U���fH��t���5��S�j`��5&�x��XBR�t$qVz��7}g$�x=fEW���e�1s�3�y?L�v��ކ1��)���f=�G(71b|�ƭ�Q�p�����5�ͮ<�UY��E�f�Y2��␂�yd7��d۔�ِz�	R���a���C�\ GW�S1�p�|)_lOs�ڬc0��82��7'^��Y1M���-���=!��f�60�6��W&n$��]�
�/p�+��m�&��زn�����n���#$��tr�j�sJ�����/z��|�Σ*>���6�0�q�"�+ΕYC �GMxE�\m�#��#28�Rd�cK�w�1GJu��г���}�o�]�#��BP��[�\tl`o��ҫ�����<7+r�p���G={�Y�YK`�H��!=��\�.K��B%L����V��MNv�陋s�s�ٕy�^Y���[j!�|��_ݴ��3_b����þ���!W����.ӎw���.�Ҧ��mv[�ѸV����!G������S9q��Y�bf/6�u�ۢk��J.2i$?(G��,�g�]pu6d�r/-R�kB䟍wky
^W���V���֛9�CΘ(��n�\K���+�Fϗ	���7~S��֓ʧB�}b%
Ot�k��Ѽ#Y������Q��p5�%��,j��YY���ﮛ�=4�Y��ߐԼ�ʡ�(J �<	�2�풚U�u%��R�|N�eq���鐳�Mʙ{���w�ub���Qx`L衬�֘P�'L��sI9�hAȽp���ch��2��S�\��d��n��6�I��W9�v�]5�0���<$k���
��7Bs+�<ƗWۙ8ԧ����!���Ѥ�,���q�e��\.���2�Γ��*�����m��N�/>�����/70b����������ż�WԷzo����͙�(�ಅ��ja8`��$�w��I�r"Z2,�ك�J̄����"6�
a��ѣ>��������_���򫅔���(߱M�2�?k�Wo3� &7!��L��W��8c�/e<5@zT:rX���AgT8�V�������4�j]wQņӾQ��t�Xt�W�S��=z.[xs�hs��/�3\�NkΉO)�^u�2Bl�*
�x9�ÿp�'�mI���Ojgڇ�M�U�4N��tz�kp�!���A����|�긄��q�"��S�T��^(���[��r�1��BR�Vӆ�o�1X.�޹���Gz�����ϳ��	粋�%���-Z�zJ1P�g�}�7n��a�q[��n�|�v
����H�_��D#~�8�ƹgV*��Bf׹E�nWmQ�n�tgK�)6U.$<5�i'�%���4�u={65K:�5pFLLu��MjU��<��5��R��|�_�T(�����*Ŧ�\C'W �(g��z����9<�z��_#� y�%]Δ�ji�CfL�G�WZ����^m�~3R�������(xE{vxo��y�dj�eY8�.nA9S�t99��� �f`}�+x̧�U�2�*�b���4�t���ᥥ����U�Q�3qT��a��4}TW%������+2g�]��j��}��}]C��'ύ+��/8��E���B<������)
�{�wI�5��Wk|�Z�S����
�@ԩf!���]��-TlN�Wi�lpεl&m�n��2�T�d�J,`�j��
cj�=����F��x¹��niF�2�JU���u5���䬼c`o�:�V�·�Ћ�+�ґx����F4g�˃/��ۧ�=@��b�����T�n���3�b����x�_��8|�����H���o�5�.�{v�sQ��,�0��5�d3>�.��������pмu�+"m�]����銢Ǝ�?Of��=����g��#>�H��B����x04���-Ϋ��'`���d���K�v9&�
p�&�YT3�X�������S�4��h\<D�w�Ɋ�%θ�aݥ�k�hoh��.����ca�Y�ˋ�+�+�V�t*�(=U�S�'Lm�`ݡzMX���cΠ]Y�Y/�k�QGZ��FȧL7�R�+zYǖ�r�H�c�V�λ���
n*�g��ΐg�*\a�Lg8t�n�l����]Y����.47����ػ���,��T�㓸����i#Lu�l�i;;�0��j�m<y�K�G@�e���Υt�5�$6���C����X�����yCFQxk�s��T�t�Uȣ���8�~��kj�>�xE�~���ǻm��eh�5S*��v�S��|��|<�r�菝��|O����&�l�n]1X8<g��ST�d�`�`^3{�͝`녵���8��\�ae�����6�+�s�\�K2�� B{���%��.�l&'�?48xn���xDbm�W��z��<��M��h�Q*K�ݚ���q���(�/�}�(�<=j�tGnx����zc�1�$}��˺�Ӛ��gn����61
�w�h�v����޷]/�
�s�Zt��C2�Ύ���+x��4p[/���?����; ;����`�̾]q�&���m��x�޺�2)�����A�J����o������[�1<wt�#.�Y8�D�L���H�#��bC�;y���sћ;v<+9=c�����;�f;z��H�y":ɥg���e��5#Nu^��q��m��͊
��)v�M7ʚia��HBS蹍�/�흓B��ӆ�wءt��/�v����񝆾KPH�����:3����������"�۰P���h��6��{س�w�oǴ�+Ȯ^��(l)�FZ�Hv='nc�M��.���J��ؗ=��3��%�6\�WM~.�v_��U��?�m��g�c���\,��U����l4��݁r�!O�U3A#On��v�r�D�t''Vi�O�<�%�!,���.���v+�>;����Ouy^�7�j��b��&��_�ձ���L$tڏ+�nҫpB1|r� �K�F:�ۘ�h�^Qg'T;l>�J���#��M?��+�u��M�T�P�EB*-Z�6��[��L;���f*+-M=�'A�g)kB��0��N��K"Di�Q:���x�#�ގ�諅�ݻàg��kF��D�wt�  ً��;ތg�e�S��0R������<�[��𪎭u(y8�'��e�F3qf��2ܜ"Ԧ�������]��DdMث�5ިTS��]�j�/��Z��Z�NB����w��:_8�i.b�=HX�yL��ƈB���&[�S�GelHR��)6wD��7en�)��&u�Ki >��ؾ��������qXݴxn6*�No��wv�6����}ӘQ7>ꚺ�'�4'r�15(R�OE�ޒ'���G{7����+��a�uo�4m
#G"k˝��s��{W{Uw���"�t�.�D\�H|A��=ab5�M�
����>�.[���&EN<��2>�:"��FR��f�؇t��n���nk�c(z�Tn�r��.���>��}a�+�g�!������A����"�T?%(ш�Q �1�XX1�� Ŋ*
�U�h�#�Q@E�5���T�� ���DUF"8�E��UR�*�LCE��AQ�2�

�b
*�0T���1Ab�"(�QZ�(���-���DDDb"#Ւ����eQ�ZAm(�*���FPV�,DUEU�`��kTDU�Eb���������DE�b�E�Db�m�`�k%ERڠ��QF1U�X1AR�DQm���R*��-h��b(���"V�,��,QV�*PEb����1�UT\��*�Q�(��b�,P[K �+[Q���QE��ZEX��(��b�j)�U-��Z��J(��+m�Ĉ��,Y��EUTA�*�R#�ETJ،KJ"�G,�8"��b������QU�TV
��F
�r���QT*XԣTEE����X�X��FZ+�������k�����{{J���M��2Wp�����:e�h.����)�����4��G�� �U���p�k$E�;ⷞ��
����g;�Hs��t����a�bnfi�yx�.�ʯ�xm��g{9k�P�:lQX"��"��ƀ)�Bq{��Ʀ�t�A����u�b�i�{=6���z�xV�����ťqP�#� �Gj�H�����42W��P��/��i�5[�^�9+i�/\1(B��*�^��|%�򏍬	8p�)�`������/ZW���D;p�����^m�y�U���q�Z��r�Ĭ(��p�q� 7���Y-�n�S<���dm�L��7.^Gb�,�]^��F�E�� c�V�逷.ؽ�.��7��j����lC��7b]3Zf	����qA�缘���Q�qSۦ�Xz$��A�{���7�԰��R<:�>'�
s�� (�ǖc�6��d���qw�/q�=T�`/�l��x�=)-&���L\h]b���hdA%�L^n�Q�)�^uV��2�1�����촸�����3��S����N)�y.�j�u/i�,_�׾����
N��KӚ�ү���g��N�x�Cy���VC~���z���y���׹�Ӌt3�^�G�.�Ggx_$������~3�<��6�~����~F���x�'��Ӥ��;D�T�8��t�=ݦ3S^��:N�o�}U]��*�^"�9C��>y4X͜<P^Ve�d/}�S
�7۴�Z��-� �7����u�ngm�7;(_�L�Ux�orQqj����w�E�:���V �K9�fc�@���$�~[�~^�e\IٍGW��(p��f�*/µf��9�Ua������1��jf�	R���po�x�����w������q��bG:}r��'
%V�[����u讯�f����K��(�\�'��9lr{T���e4-��V��	���!rm��ONX4�o:�7[,lVKՌ�B��`8Dq
C���b��=.h����U�n��R�I����ۜo*���=�6��O���s|�}�J�+A�o�`.�ra�[���,l�K�R��,�\oҦ�<(��\wyuAoz�E��n.a�1�$^��lJ�{�`����ۭo������J{We_���b�<|.���|�;���_��_��.�=��ޯC�u���*\b��� )i��|.A��:��'���q�49��,���~qx��)���XT�4��v���@�9AA�{ca���,nM���j�n��E�Zo�������3�v��B\S�a��m^�]���*����H�����e�(TWM	MH��m�Y�tׯo�F#�f:�%�+
7ۛ�Ln����f��W����ǭ�ꮸ�_:� ˆc|��3hF�ʏ�t+�F���hX:b��=�,x4�{	Ex��S��;����5ݞa�T�Q�(�B8�\������A��/n��Sf��r��ʷ��^TŇ`��ɊK��zS7rm X�̖�ѝB���<>�@OM�������5��`L�CY1��u�8IN/̪��LN���ƧS�϶�k<�op:�Go�R�����ϼG�0f�z��L�(q*�.��w�2qYۙ�.�2O"�	V������P���yU���CLw��L��gS;�jU]z�f���z��f��J��Z/`��^�O)P�p�x�C�Xz�i����'�*��c{�e�5�x<Rp�
Ϝ�G����ӿ��V�������FЎ:-��4j�ܱv���ۄI]��f0T"�k���ʾ�ܝn��k�/����z���땣L����/3��*9�d�P�x�S�t��[0�qE�ݩ��*aP����Q}��o��������wnU�@݃ԯTN�����Z�4!�����J���:d�ug6�;�f�HB�ed���b}�dk�3"IW���������3��v(���T�ǎ"%����y�{Oc��Fy�V�٭�S4>ҍ�e)�,��7ڥ���_�>���L�b\��(�`����
FÅ�sqd\h虵�[�����3�⧡A�fŬ�O6�;PY������Q�g&�������q��u5P|�6��p�Q}j���c�h��0ƺ �^,zUq$�q��צ�������9����OP��#�.n{T^���3Ǚ[8�g�\�}CIk�E�Ap�����|=%��Qg���Yw��\�Tn̸���	��|*9�ǅuJ���0�K=R��V*<>4���6�e�c-���)wp#*t�dU�r�^�v�(�T�H�R�>�*���(�D�N�oW�&�vnN�V��˯mi�hU�(hÅ^�@xr��ȡ�M|���l�g���ZSل�>�
�~X��U�U����c�\�u��"��W/Z-J])����~K*p�L�)-՞��z�{��Ћ�@W��Q�o]%�r2��GQ�Bb�\=��ceՎR��s���:j�/�jz���4X�W�5��u�%�W����;�[�$�؊���F�m�k���[�<|���CS�!���IR��"	�������v��C�ZTc��t�4�M7b:�7���J�M�j�9��c;�hl�;)�ơ#>bN�¬+��a���W�lv:yN�Nk�u[��4�P�"ojv�����U��6�"�w��ް�;KG.6n�ґ��<��̪���c�/�I�c�r�7����kM�F�+'�$��g*�����K�ӷS�4���|*��x���-��T�۸B�fsV/��T�L0w6Qq�,��w�P����<�X�;�W甌h2�e��@����Q��Q��
��[g�FՠF�*`��J#�4���w*��69�h�;��B��־}*sb�����1a�/UX^i}\�G�Ck��Q1J8�YN퍍�shƙ�b���$���267S�t������Wk�|��#K�������o��·w�,k~S��ј��z���_�A������̀�J��Gc�����G�k7�K9�3�ݳ2g�� ��؄=k|;i�͗�P�Ї����}C�->�V�HWip��:Hg7�ދǒ�|��
fz��B�3�oҥ�vyMd3a����t�ȋp�� ���]�Q{����h4�۲F��^����/b��iv��ł�Q�o�2:a��`��Y�
S�D>�1�:7���E�H�/����W��xt�[��+Y��F�&R����#i4c�js����S��(���VWt>O�_������3�;�uIN�2áY��!�u�(&�4�<�W���6����%�s�[����u��L�8�����}����P�ku�X�;��#�,�t!�bՌu"�y>>�aEB�,+�=[0J�}=��n��.���
c�-&�\51p^9�E�%&z�#����{a�	'����A�6g�"�
�)���t��Ch��72�
L�����(-�w���Q��D�Q�0�\���%,M)ֈT:��gi^'����2&�A�RW{k:]j�u�E�F}��93��wT���)؜�Nm�3�U�o�xg���})�o��7VR6)}�����l�@����^�~�uoh`�+�Yq{n���֠��o[��L�W��K�}��Յ��p�8ˇ�lR�8`�͔TX�x]�<�M��\�V����|ޮWI�Ho�v�ݶB�U��a��2�V��k�V�=�U
�7�Q���Q[K��*��Ŭ��%q��$󎂊��W�m]��6&+:0J�:,L�ƭ��n	Y�����u�s�G3;x�951�{�pu�x��
e%9�ᐈ�A���P���sG��t߼4<�1�߆H�q�څv8(�ɏ �9rQݵP�j�z��*��v#-�8��5=ws(�,B�Xo*%#p�jqE���ٙ��Y�7	\Je�`�+��O�^������R,(�y�v��<n\g����x��m���:}W�i�]�.v��۰�H���]�ѻ��p��f�z�����Y�(U��C��(u:��Z��p�B:��@RZ���`*����MF�kfQb\ڇ0��ϭm��*f��x��ȩ��=(��[�1:D�}g�^j�9<7�#�WPL���.k|%-S���+�+�׼�9K3��Y��ak�{�ܖeN�TYs�=�����ۖ���=��G*tܹu��H��2IZ�k5޾wfa�}{�l7=�������G	���p�Y��4먷��X�X�OT]I��7y���
��M�B�U�9KL`��Q�(Ӈ��S~��(�����y>��W_�M�政����颦@8�V���<�2�W%����V:��mȺ7�kgם��v|��)�Eq�"J:Irq`�<��E�����-7Y=�q�X[�Ԟ|�wCÓ��5����1\�>�"�i�(k'��O&x�iX��'~���'/�W�����b�A�^\4Ch5y:+�ePdPͪ@߲1�˰Ӊ�vT����Υ���)�u�D�v���p�q�]�RKOW��O2�,�z��Έ��aU��0N>�'�D����A��~��i�Z�d/�5���\����N�ri{n��s�Ϧ69ty�E9�A�j�`�ŝ��niy˱�3UDA��5f5�ɻ��׹
���4����yW�E��2�ׯ�xk��g.��LWU�o����V��ّΰݩn�b��P���ތ���`��ef�>Z�I��a�өh�7Lxm߅�Obp��X;�����#)Eܮx7!��϶��U�p�*b��D"m]�S�W��k9��=Ud���(�W��+��YV+�X�2��8�)��M�
�/R�b�:�E�Tu�Y������R�|Yk�-5˒���ᑳe�"Ծ�Yp�uC5}9 57ٮuٓg�e��*� Q�Dq�Nhu��}�4�9g{�>�e`����f,�m��I��̃ò^z^K��<DA�}ZI�\n��8�[C����~�����i˽�Z3�k��nl A.P�/T{���*��'��\R��M���4��}]^��⑙{3;��<;�H��xe�ʽ��1���«��O�4&�T�/��Q�ݥW���\����@�.��*��͛�8V�P�����@�Ϝ)pLu*����+���V
J2N�Mފ��2�l��v�U�xɈ��4�\ťY�Eȁ��d���`�Jy���#bOvV+ƽ��y��\iJ�C���ֻz�Rֺ9'�x,y6m��U*ڄ��l�����1��86��INJ�r�3�Z}+w�o���/Ԍц�b�U/����;>��9�y�`�(l�^(d���ݳ�Bc_�bsqZ�h� Leg��_���B���zB��r�Z�:R)�63t�ٞ��$�܋4�}z�]s�
_r���;M��vZ�g�!<�eD���Vq���,Wz㳵|�I�	2'���p{듫��U�]��M�(�<<�ĳ�����5x��vO����U�M��:0�)H���9Չ���"���|b��PY�lSڭ:w:���hP�Tm��ZWF*n�wqy�Y��K�6�C"�$���g*��䕾s�NUH}-J"�;�S
n��)�������կ��T�hf�."�7��N��}����Y�:���M�s:�J.�z��	��:wb��uE�4��T(��L�E�u�#�Vw���[�*�\��E���(�%�N��f��Uay�!�\�G�Cj��*���3���fC�[�<̑��ү�\dln��5+F]Ip�3
R�&Q�2G�p�e�-��Ğ�V�.�%[���f����$�t N��yn�ʅ�=j��p�4��a�F�ٍ�4�gxk�to,�*��$ɺ�#��>@c�����`��	�;0u�S�{ٱ�{������P��6Cn�=���.�*��W�����	�kU�k �/zr��86r�w^�GyCB7]�T1*���6\�+�+.)�u��&7��w�b�/�3�������m#�;6^yX�JBn%C�,Bx�y[գ�6�U��w��ַ��xa#��yx9�
�Il8"��;u��4:j�b��aP�B{U�x����!�Ԕ_�kV���"�x݇,��T�3�؝�awqGA�K�M.s�r]绱��R��+}9��*�ӊ3�d���:��'�@���H	S�(����4sM�-�Ŀ�uf����~se��j'I���w��F��][�P�d�^V]�=9���m#P����hPV<S��3�b�`����Dw��+��>1���.]j��hjU��5�Oy=]�_C�!�(*xNj�J���*C�]]x��ԃQ{��̨����[��Y�eF�٢���,�auAu�$] �=0.��[�_{�XӸ�<�M�=X���a�,�F��j�\In+ٳEcrQ�����S��e8XV�}1k/����֠�w[>�Сu�`kE��vV�[�B�Q�	�A��:x,����=Q}�J������+k�EP��M��V��Z��:Vp�nZ����X���gayd>��U�����l�]S�:�]&Gs6���g�)�uׇ^�����ws`VC������O�Һ��F���."�3�j�&���̧oz�v� |K��\ck�T�W��z�tf��&�쯰Jzd�+��xR��AKw��Uh��pQӂ�0^�s�E	�L���|��2�(�.ͬ�j�;Ot��,���f�9�DZ_�:��s��O��0`𱻕�ś�Nx{��P��u*q�V�Лb�a��&�q�7fc7��p�i[⸕A�J�Mі�'x����	�%���p�v��q�a���s�,�PU�;�P��bCV��nWv;d�[�6�v>�Ff���~�˛�.��]M��0���V0H�xG9�|u� ,��C�ˉ��这��w"1h��̖kZdl5�y�N_!�oo7�D�]��P⛏(��G��ݚެ5�]c�CRJK�H���<P�ia� ���a�V�����Խ�C�9��o�ѷ�/����ܜ�Ct��wf��]L�4`2�N�dѡ]�w��o���Q6He�ʋ�Z�<����0j�J�3��Y;ZP8M�z���)̅1�!�}�=���ZC�6>��n��r�6�����nq�A��`nۙ)�V`CpG�f&kz��Uuf�/Rg�ri|�ņ�ٴ�j�6Uql�ä��F�{��~�4�KY_s#�QX���"L���U�D�)�i�(��'(�R�7��s�iZ߆{�'��S.�ŗ�;&)�J���(�x�To)��\���H�=�cU��-������t����
Zt%@���{ �og6����0�=8(����Dv�V6����}�J��U��3�Ytf;�%B>&�RB�+��k�X1q�{�	�Z]j�����[���V�za@��ǥ�>#J��뽹� W ]���j���ºfk��X�v�9���b�#�Q���8�u_]�7�l�Ef��L`�����I.;ݏS��]K4�9��f{zYzԍ�p�j���Xh=N�f��`"��A��t��Ο��OEQO}�ʰ���kƍ���D�|�xU��m 6��T��C(�|9 B�":�"�2�$hıZ]2V㵼�5&S�ՠC���૦7�\<�[�u���3�mο��@q����<��P�/y�MIՃu9o��r���B�`��Z@u��gR�l�n��-�L��������\7�79�(w.f�e�Kݘ���"�0l��k����ޢ��k//]FP7N/8I�b��S'ѥB� �x���e�����%����)���tk�u���UTEPPEGt�ڠ��(�mF*�j$�X�֪��k*�����m**-�X�
�b1b
���͊���cP�PEPKIUV"
�"��EU1�*�ьkDTQm((��֢�VZ0ERڪ�(�jb�UTb0dXȣ��T+�m�F0b* �"�(���r�r�QAHԱk*+�UVڋYEF,EX�1Q�H��E`���#ADm* �b ���1UUQQc-*(�E2�Zъ,����┢���(U5�����`�dEUU�TUX��J7-AQ�DR(�ETAQ�DE��[��*
��UjQ������
	l,D�ETH#.6"�!��`��TV#Yb�AEEDQ�AVҊ�1UU����"1�R�E����(����
):�aҺ�>f]i�5�3�[aV�\/���jj+s�bvʥ�E��,Ԫ���ˆ~כ���)�N�}�R�����r�so����S�,3�w��Vk�m�e��Z�c�U���^.����EV���{2f�t�{���W�"��l�x�v+9W�Y��n�^���7��:�P����c�N^n۹;W>���RZ���싨�u��7�|�N8E(z��<���|��ŇJ��G�؞4�<�I�u�Η��$g��P�*=.�+3��6�K!!�t2��=��o�ۭ!�X��%�3��=���w9�vp�Uq�R��dYG*�Ϫ��O���\�.K���屧�ߨ���b\��ۭ�R�l:�3����(Թ��x���ख�z��Ҕ4}^B�{�o��]���S�f�>4��5���1����	v*ڮ>0�z�ob�x}����1��ô/g$�[����h�p�18肍bHe��"��#�[Hبy�9�����Ӕ�5���+��4i9�[t�T1iՙ��%�tK�WPG|��AG�Ֆ���21���ʻ��2�};�s)P�U,�e�`6R�$]*fF��(ǖd�u��tS��u�]��ՕDue��;LCm�mf���d�8�Q8�g�"G:���,M�-� {/U�*>��f����[w<	�Aכ�-¬��з���W=MC�L�ٍxUт��{��W�:���ɻ����vM�����KvG�2�ؼ_�!c];6ak'L��xw�Z��xq��,;�N��j,ܘ�Ը�Q�f�y[:��Z�6��RP��3�0w��
ڷl�N,%
�%ϣ�QR�"�ћ�M+�j��Ty���Ud��^d�dDv���-\�ki�U���4ԋ,4`�ǝ�O&}&�VP�W�eӭ���2�D03C���\4'�2�yx�W(g��B*򫁳�Nc�q��;Of�/u�ǘ�q&޷�o�80A=ȃ����X��`n��pہ��{|�z�<���f�z泥�0j�a�T"���V|ͬ�}�Zu�ΰ}{[I��D�M�a@���)<���bF]�/Fn���=�j�(��(����Ul��C��<�hu��vU �yKam���_8��ϓp�5�r���\E{:E�t���m.�^�T���Y��3��;R����7���l%bƛ9��;b��'�x]*Q�N;�f�{,����Y�0��]����9|�um���u��r|Q�ù�GD
�J���"i��U���8���:�l�������z��w�����n��T�G�����Y�lک����j���o����b������
�+˲b��;�/����Q��*n^��O����[�ǸP7��`�6x�{�S)Cx����f�$;�=K��OT�/}w,��^Iur�O���7q^8ה�z�: �,�U�	D�GQ�zl�6�E�m\q��w��hH�1Qq�����[�}��FE�}h��󆾸�EŦ׋�(��R-�FW�ٛ�}J�>��n������}Q�&�"[>P�+R=��9��6����:�{�t���6k� B�K�<����6V����W6DB\�iU��Q;���5�W>��=����9�+�L|�f��U��t��SYR΃���)[o!M�V]���G	1��P�׃�k��oV6�x'T�O
�L�� '��d^��C�H\(������پ0�iW���yPdH
r��b8UiQq�*Q١n�e�^QG1m��7�WI���X�Dq��kU�=�_N.�ׄ�#K��2t��썰+)+n���!]ov�+,WeZ���#�qU��V&��<t���״"-��L�����pl�	'q{�s7��LY���V�ʖ�e�va&�x��t/;jg;^��v��az�r:P=F���C��֌7�
��GC^a��x�8Y�o�z��^0������Z��2�=�76���<s˺s�6������p�>��#�5˸n���|&���]w��G���,k�G�ۤ�F���ˠ����c����f�,�<{�P�j�r�۽{(����Q�B�Ou�muUx�q��ˉ�!�K<��Y��^�Cq�c�S�PO���qPo�;s��������TP(�N�<lj�@oK8��/�c&RSqP��T���5h�enӹa�ѳ��?�i�4��^T�]���cL=3s�A���)�r�k���byS7�27bw�#/���Xap<���>o�P�di��6���դ^51����YGD/���\{���ĥ7�>�B��C�ѵ���Q������ϧ�z���>��vsl�Y3��5$��:�Ѐ���]Pv�.Oz�Hs��̸��#���b�k�W6�'A�|�a3�D�9x:�����ÂR��;�Ni��yn���FN�z�@�N8��no��R;�Q��k�l�l�`���MG����9`��珴��ַ�_ޫ̼Z��<ѭ2-�0�AŪ(�v2�fJ7X�D[;,��	�t�z�$�vB�,�<���eZ���>o(Wx��>��e����k��0�{�.�3(��գ�1M����D"�`(�%ۘx�JΐlN�+�4W�LG��n���a��}�{u�P���S�텙� �%.��y�~��ޗ�Ԃ9�����:�t��Λ�w�V]��1<�s<��L�e��˯��]�k#�����]�^Q�;ӥ�ɬ{�/ash�Օ���V�e�}(��ᠴ:#��+�:��.Z"��Pm�N]�փ��^:���e�r$/�`����9/&�	Ţ�YP�ݯu�^{��Ӭ�с������賖��Xܚ(X8Yu+�[� �;�ɧ^�y�Qv�\q���r�z�h��-�&��߃XC*h�Ĕ�EŪ��K���K����v<�<5Q�~��5{�,3<@#�Y�C��.
�������\8�5ײ�u�7)U]<K��q�#�(���]����\�{���˓�1��S�f���x����{��+���hH:�|Q�Os�8���z��6���|���m���w�ݜTh�,�M�a�e�,�GP�l�d'�<�"���c9��s���!F2�Ь��)ץ�/"\���I���8 �8|9�4�����WZ��d�#æ{���QgÛ䡿e7kL[�[���9t*����XK�4-U#r��<�J6Eb��˦^{ǘ7��l��7�	�QrF��-�뮙f��.j�Gv?�<��py��&@�oH�9��x�����|�VN���{�ڧ���3gk
x���`nq�t��n�����"��w�P��	�<u�]t½ ���8 VsS�Y����[ckf_�.<�����3J��M�-r�J'�b���E	�{�=�n�ɋ��p>�6�8�O�k��U#�����r�<o�$X��e�ru��ٓ��jT�&1A���H�a��p�B�|�V�G��S�����ҼXq±BZ���İ>a�����#of�N�o�l���Y�n��C���#�z{��R��(�[�P�|�z+��m����z[���	0��40ـz�R��K��=+� �x�>eNQ.��gZ�ҧ<кju��w�����oM�|�V++܅\Yx�:`=��Iw��zz#�=&��*{�U�+���0���f���Tb��1\��R!���:�sϽG�����6P�����Si��ȳ8c�9��~�s�-�{*�:fY����Q��v�NjfU�C8V��k����N�-���	{f[X�~<g�,sr�3�;w}�\��!�^�ґ�V1��è�a�V�`]�F��:����u�E����n|�m���ߌ&@V��(��������n�T`[��^.ꐔ�Cp �kqw��հd�W�^�&��p�%�q��ʵ��B����2U�����{�F�S銲 �ٽ'i-L6��^��6�1��p��;��_�6V�ݾ�{*.Na/���G�W���T���I�q�#](�+�p�g��C��͡�a9࡙[7�u{v ��\p�4kք�!d2�t�*�Wi��KP�Pu*�ݤ�U����F�NXRС���:�\`�'�Z���u�8e�<�x�'�Lv)ʯ^<\+oo�fV՛=Ow�K�Ԡ0r�ڣ5���r}Nhu�U�ߵN8�mˈ����؊|����\�+���j89t��e�tAf�`�3�\I�D#��逮ޫ>���􀩧s�"]/V�=��=Z� ;t.����K��m�/ŝ��_�x�og������-�˷��]"$�l#%T2f��;�B�#���F�N]ċ�(��Y��k/cr��ެ3Z�sQ�C�Ү3��R�7~0�+K��BZ�'�w��cX}\����4�^w�4듻}�0U�S��]KI���x�~V��p�)�|eU��l�`+[����K�[`'�wj_{xm���P�&�|��؃Q�c�7�
�#���"��1\�-� �ޮ�1�v3^L?_�wfeN����':_�=�w���'�ң��'�&s��{��vN
��Ќz\*����׈Ӗ�y��1�v�����OŻ;�ǋ��@]�+���2�3NG�`�nM�e	2��M��!������;�~7�pq�	�/���+�!58�n���H�mba���>f���QЉE��\�:E~��a����%c��@J���lG
�+�dm��vhw���a�9�V�.�2���{�B�&�������"���꿦�Y�B��J̈:�&4�`8t��n����幗GeJ9q(Ccb�H���άM�����Zx-o�+E������"��>��t튾�[��N���p�eid�˟_M����>�=�5.3 fjg��X������.��E�X"ڮ�N���.1-��%YMʅ�����,�à���}�b!���l��Gg
�+օ	[�
>���O2�p8�Dh�,�o
 �EN�&ū��bk�sQU|y��#
k�O>u��2�ΨŇ���$t���1��B���y5~�Ͻ�Ym���idb'���)p�F��e����������f��7���uoU�!���9��ܽ��ibU��ᴡ
P�Bҡx6��BP;M9�˅!�৯:w̎G���8}�������S���ݴ�P��y���!��KqM`ͣ�F{6��Z��{e����S���6�n��N�����3�<N��ؖu0����b��0�;������v��g��]&����}�s�)S��Gn���� ���!�R�9�(���N�Y���V��φg��^��+�6�=��~�>�@��o�n�1�調oe��9ʱAŅH�aפ*�H��t��#=
t݂�荆p�Ȯ�ZY�S�t�<yL�s��{�X���*ϟ>�C�j��ǲ�d�#u��DM���d1��h�2�uL��5�`���5R�(|��|z+-Wz[*��Z����Ii6��չ]�!��o��ܜ1ٝfW��R��I����X��e��>0���T'Bdu���� ۲rV;��/w����i8�����8ݧ�{�d�D�}�x/}�YT'5i�4�e��G����)���5w��օ�����_�&�Yc���L��=(T�ǰl)]��{3��y��F��б�^/	Hଜ�]=�����vx�R��4r�̼)�����U�Ķ�ӹj���ݽa��,^yӅ�Cѷ���Î1M�`�ޙ�˚�z��7-7=C�<�N�tk��cT���=g|�׳�xj����)ؗ*��w��r�t7pI�φy��vq�ֺ�a��٨��t���x֍�Fs��q�W���f�5y��l��<�^h��+9|�� �cۗn>�e���;=]w�b^�,�n]HCL�.4+­�O/{��4QJ������s�#2�R@����8u��5=���8E(�ϝ��Q��C��P�MW,����T(��I�wƂ�|}�u5g��]�dqn^,eD%Ҽᐈr��l-�*��v�����Pumx�KNꑿK��dYF��U��<`���~'���_3ٌv^]��[Ii9\�l�֔����c[��|��q|p@xx�u���%t�~~ӫ�<�K՜S�������V%{�#�A��iv/k|p=~���.��z�d��ˬ���v���j�"�n��((aL\�����;eU��ǅML޴j�G�|�EΗ�����0xS����
>���ʺ:,8�P(KP���P�ul�uz�(���T�������|z�{��ز����5*N��ʫ�n��,��F��Z�g:�=�ok�EV�̐W-�vQ��B�7��y��yD�^iL�<'�1`�F��NvS^^_��U��=�` =^��v~��d���?����Q�Ř<(k&0��z}�7^���j�K���|�����ʬ^���Bf������h�&ȍbfNJ����/L��eM�"G.�n��$7;(q�]��1)��l޻gs<D��x%	N�9,S�Q6Kx9HDz�=��$2��f5j}1�/[��]��'a�N���#p0>�4N������։���=n=�r����آDg-V���%�X��^p��F��he�M���1R���j��m��:A�!:�ފst�F�+z��Oz���q����,��D�����5}`����RWF��z����ɨ���$�rzl
�u&�a� #�����fd���7{�/(�&Ufv�����o[�s�v��'�z��9h,z²�JT�sכ�k�����W`�����WQ'�;p8�����x��(>{ͣ�z�)fb��lY�]o]GC����~˅Rp��]��Z��v�5=s��Ҋ@��RT��C���[�{Ҧ�Z��G�M�ٓn6m�867�9�L2x*w��&���]l�e�x�mn]�]ǰ7r��<�{��^ӧ|��Iu��8�m�H�f��ub�743PM�[�Nn)��� W+�<�/xuBԇn���.z�&��'ɝ����;�鼛���NjcUaHt�L����C7��β5,U�L�UW��·.��IFM��v�}(Lٕ��>�(���W,����B8+2EL���@�A\ҧ4p5����Z�� z���yN����U�2���ڛgd�oWZ�3�b���H�5��D���,�i:� �B���؅bs�F�=j��[����ѫ�ݹ�wX&��H�ɾ�j^��Kaeޡ][��^6�;T����(���ޟ5�H+��m���8i�����1g�^��X�#-��;�5�E���xlP�tb���*��p�m2��G��ӅH�r���q�h�O���1yd��.�hJCG�-c�j����D�&]`�C#8j�U�hN� ܺŏ5x�;%冦Q�.���ܚ)m�:w!ON����wU�����c�J$��&�i���T����WK.'�9m\?b���r�����s��Ǫ�t�e�6;Qh��Bw:.�[p=�5�̖J|�KIST�̀	0�nu%D']A��5����Q�ۤH}�`��d+�Q��x�v�$�觮|�X�&7{8��|�Y�i���ن���q#^�Z��As$���R\SQ�N�t��\{��>���k\/���H�m����\t� jr܈^�2�ݘa�B1u��oWn��W3�}6��s`7b��f�Δ���M�b��A��z�h���-�!�:��щ]G��]$-;3��sJ�Gw��������=�_=��E� �ATX���X0b��yaX"���Ub0Ub�b"�+*1��A-%U�l1UUV#U*DE"��DX���UE�5,X�QG�b�,AAAQQ�(�(���PE�(�Ek*(��AQdUb�
���F1F�F�DDb"��V"%J��r�PX���EX�F,Ve��J""�*�"�QQX(�Q�QjQQTTF��X�`��bTA"���Ŋ��R�b�h�U���X��(-��j�`U����-VґQh%��( �((�F"��@DTAU�*�~J�1QQAUTD�bV$J �b�"�b���TQ�
�(�QUPDV1,\B�R�TՔUDQj�Ub����*[*������QQ��b�ՔUb*
����Y�<ֳ���V�[t���� �u����kwf{���kZ0�����]�q���D� V�3A�ܺŧ�`<|�s%��Cz�#�Z3ra�զC����0{�ڌx�˵])�e���R�G�yI�|H$�����s�;B���`mwZ���
�B�uc��K/w�Y>��#W#�;;q\3��)�
���uv[!GP-�(B�YR3�\I����q���D_�}��}X�,c�-���6t�>��Ŏ�BƐ�ۄ\P]c_9wpoNl_��\e����1����H�������W�[��F�q�r���d������L�X�9V-:��6yz	RÑ�3W����FJ��}�onq�x�M���^�xx��Ls|�t��<2ʘ&Kj���<����U,t<s�R�)�P����I�`�E����qȡێ�%m�����W*>���8�j�9F*,�*���C�~��V5�	�Oz�C���=`�/zܙ��)�>�ͼQ�U#/<-M��0�x�����jN�w��8&o7R=��N�eK�7�YՍ\������r|�����m�7�fĳgk#c�~f�Ȭ34�Ut��f�jֿuE¯l��n�x-��Ͷj �����zv��yh8\Dˬ�!�r3B�%�;��L�$pbIԕ�f&�c�8��n�bT|4Ig6�V�e_4���d��l���I��$n5�����źW�EW��[i0t����3&��UC�4s&�%Sf�wi�m����Ah����
k<�-3ю~�;��L����i�Z5�g�Y�z"ggN�%N�����t�^��ϙ����O	��򊰢Э�Z�2z��^f�[]$@.\�)	������	s��)�XL\Ѫ6g���gLDf��\Q��D�W�b���Z_��L�6>$��]EЯ�g��[z����9��dW��w�ws{F5��7|�9�K�+��t�Ҭ�+Ŭ�!���	��o'!�T֏%I����VcǗ���]�p�x�]P��^::<��c�
F�EiP�az�Q�g��跇���кۻ����s][/��0��3`nM1��t�M�`$�,p�C��U���?YS��p�!� fc8n�p�ʔkٲ�6p�MgN�$hV����v*�m�v�j�3:y<7��3����EYv?��#�?�I�6�X�K,�\*w�M�/>�N�*Y���f�o���&�Z�s^c}�x��Щ[�
(������7�$�[�v�
�F����m����4*&)k��������RT�����[�!�g"F���!��k7Vx��s�J�D�*�LP�f�>��VL�U��+�A��69�ӆ-���<����<Ү7窻��`��,�:T����~�L�/lwL��:�H�5y����!d(�nYǒ�,��3~S#v&�JїR\#�Y�iK�tp�V���긱Oc2��noxѹ#
�X�D������<��e�xS��W�#"�xs��Ux����/s�3�k[|p9��������Z�f�#λ7א�ހ�;u����N��7��k�7P�r��F+9�p�U�m+:�-o/f)�t��Jqy;Q3L~�lj�^@��W���|P��v���V���xJ�S���a6W67j�v�q˞͞��;���ό����
��Ta���XMdk�4Gcυq���B���t���|�����}ٟ)�����P��U`>=�U�
�'����(��%�ݏd�U�~�i.:���W�^"�c#�l}Ұ
�j�Q}FYͮΦ�r"��n���$`d��@�+k�c�t*��)cY.C�!}������(\K�_�����M{��]����^5~1Q��k�����˚�ﶖy���
;ӹ�B��=���8�}�������m�N�NA��t9�ꉖ�ʩ���w��z�	����#�a�f|-�I۹Ɏ�z����&�s��HG)�����Ba�+�����@-���pY�w�uOɜ�ÞS��ʲ�,��)%�L�l��Zƺ�_1�ݘ޿[�9{{>7^҄����	I�,�4&��澺�+ə^::�n_�$��Xd�v�7�#=�nϹ�Co���Q� ���3�g�!�o���&�hn��Ku<&��7nr"Ak�"�*���YF�������+B�1���@��|�[��4�=�au��7U�?N&�Q�W�R�������v{����賤pOu)����tϹ�a�Y�\��C&)s(�E�\m�#�\�b���m�*��~
UwF8d��z�e��]���T�T����K��F�ʈ[�;�U���<QhY�u\EP���ȵn��g����-K��C��hc{�Z��o�q��!���1c���u�鯐�K��jbݶ�$ ��S�Sҫﳾ��&W���x�v���������%�s̎�<�"��>��\��T�TSsFxC,��Q�|!�;ex$=Wp�|����U�\�0|���%�w5V{\��fҵ>�Ѕ�Q�t����Gp�ew�dP�#<��튮:Y�6�yӲg� \�ћl�z�Lm��h�ž�R%�g<�켠fͽ�%8�C\���C��`���V,w�Z{���©�2��Y�L^ZԏH���w�.�OM�Ǡr�p,%�{q�٫2-�1"%��%Dw'�r&2�ܡ(,���V&�ֈ:�i�F!��������(jU��Ҫ����R���/)�G���с��<��2�C�0k��"�R�ՍS���^�etL1�z,"�A»��ͻ�EA픒��<b�ޜ5�}_:�r�l�\��3+Y0�!�j|�&�X�;w�ġ��O��Q�����<3Zᶶ񸅊A��MH�ܚ���ÖF�\~��㡎�}�Y��Q��$��ǋ����-���5��_�\�ʔ+҇�5]1�H˗�Cz�JMthb�9��$�Z���>3R*��,N[k�)n�6!�<צM�~�>���𺂅�8 &i+��:�6�+�;�L������S���/Z�����T����+wM�<j԰hNm2M�t�b�Ht��,�ك�v,�����|�V���͠�ŞG���é��:�^����f���磞6O")U;�i���J�<�4y]y+'�/y�*u�ϥ�z:d,��ޫшM	�=��/F�m$N�,9��1���A,�D��^�v󣑺w��$��k��nrqi�N��'��,��5玗�{�Rw0�ן[;gq�Tœ<|px��`�ɷNwc� ���k,�v��.aO�]�*�G&�0�,:��=��Gv�L�	�:�RG�#n�;��mGao�(G:��
pT(#^p�#���K��xmg���pc/n�i�g*��6X�EW���g�j�G�R�õ�+A5��� 㡑ݎ�8�{����.f?uom�v�o��i��7��#����\Up���t��OU.s�5/5��x�T8���+�OS�Gﳘ��'U�(DNG����fk���8/�#L,Q*��X���Z���/��J8k㔡�����.;���*d��(a�$�*�.��s�}��'�~�`tw�e.Z,O���],J�唙�6�����k�14�{�����/ﲳmv�e�\#�:�.IHL��خ�f��F����^�6A¸���a�=�f�W����A�߆χ=8���+�*�Qt(M؇[z�Юb?eB0��Vкg��]���҂�1�]�vV��k�Y��ak��B�Q��Sz!9ܩ��FAf.����Kݸ�˼6���xe�>��5�l���ZS��w��E��<tqu�M�{���DEUD>�l�����m���BБF�wwA܈�zG,4:�構�}�C2e8�P�o�C˙ꝕ���܌�̰ݫ���sbM���K�%Mgw,HWK'��T�o՘�6NH���f�f����Ο-�42��� �V�h�]��"�{���R������ޫV�W��Ն 7�^r��|ە	��w7����/���jǰ�o��d.��E����<��|��YΆ\�a��0�k&��j�����~�Wl���p�)`�@Oj��4� �"�>�QS;�*[u�J�Z�ѹ�`%(�r��U�a��V�͕��ıCh�b���U���"S��g���-Z�_d��>(b��Jj�nĳŚ���N�wD�J��R\q�FX�e˹��3U�(�f{�)�+ԗ����_9��+]yi�Gc��)M�	�f}}�Hm .���7[�q!sR^3���=�:YA�/>t��9�4tka�K�&�<���^B����5;�Knnn��V!�VU_o�G�+��C�g�˭(���l�bgn4؞������vR���򭙗�=vD�]�Դ��!\��+Y��J��$yY�8k���@{����rJW!�,�̙�2+��U�f���;B�<���Ǚ/<�t�+"��qss\��f
=�d-�31��NC`�u�O��>�����R��d��=�P|��X�G���vWZO99��άO 䝛b�_s.��.�Bֶ�㸊�;.�	���%P�R&l�t�,xWWA�D�1�Ҧ՜Q�=�\��o�4��.{=ݤ<�H�ǧ��٦ᜇU���L�K�����<'�A�ш����N�.^cX�����Ud���s� &�#����z{A�n�TQ�����jn�ߢ�H�ٹ���LU��bZcZ=�B��zl��$/�`�]�aR�U~�\���{[��۽��&���Z,u��m���Bq��yN9
�V<XPK\�����SաM�z�VQ���({�+1���%�3@&����o�HP���Lm�=o��c������-��*�X{C�	�nEg��r�X�f���ưyB;^��%)z=�ʽ9Ѫ�Q��U�~[@���͔TX�x]�E�4����n�cnю���>����n�9��eV�9�(�8��!|)HU��P���
���\pԹ_,<M��K7��u=�����N��zg��؞5nIX�DP�@v��z��%ݮ���RF�^:�F���Њϲ����;�uK�q�)ٵ�B8`$�O+k��xf���UG�)�����Tп΂�	��ͨ����Ѥ<e�N6blГDZ;&MLi�5�J�{h�v5�J��Yh��>��:�`f��-`�՗c9:�I>�E:R��d�b]�k���;ޱ}рK�8,L�ƭ�5t�D,�E�*���
�
��\���F�\���r�Ӭ]�����U�B�0�KqX+U�������)e�e8�ov�zs�Y���@��f����PN=��3�E�!|^�i�VJ)yl���$b�k�>�J�a�r���6fÖc# ���(v��:9����;���x��r�Td��rG��h�y�r��9M8J�n3֝Y�t�,����dge���c�L=�6|�rT�}CM�B �avvԸ�������ҫ��R�u<jc��&<�k��Sh�����_ѽQ�hՍ<C,��[堾s�ZO�L��r�]e�^̓P�fkEP>J��5P�.إ������Y�Y�iE�/}��"Od��+����y{��4��W*�[�4��P[�����OM:'%���LQ�K5Wq�����I�.̥��^�U��+�IS�L���U8���鴊{/̊�2�����>�+��{n����4��z�>;][Y��}n�sx��S{���_�	;n�7N_��V�2�����V�˹�R�C�J��PEKb�ͲY�vOL}WVJ�v(
z����8�Rޣ�������Ϋ2�k�qd���|q�����Pp��{7Uo07���+}�GQ鐈��@�J�T�:�Ĕ����@,h_s��,�Մ��gY��l���;V��9,H����������x�����M��Ѐx�i���I=��P��cX���*u�/*�ѡjxз,͖I�fN��e@mk��ü���3�X�W�yN��X�n�U:/dK�OES��6�16���yxt��xx����K��C��^R�zR�����ٗ��/�[�ڛx�B�p$�5鍸�#N�K�F�l�A��,(�����,.�l�]"�z�f����FR�V��~'����u�%P���Q̱�swvє�ַ9��2\Gqn4k�U��>�����qr�W����2��=P)���ۓz�{�0%��-k�������!/�u��2����i=��P�ٻ�T�'���߫5F��?<�}V�òZ�8�4��G���+���.;;q�'�(�i���/U�[�����0�Cb�.�W�V�6x}�]avx��un�+򿾴��m"�`�i�ޝ��r����e4X���s��7�����tbN���|fم��=I��O'u_A>#�<	��b�JIL�r^}��!�i�R�a
Nܣ{>����l>�K�MH�Тs@R��m*� ����Ѝv�d�D$G��]eQ���R���&�쨇2 �ʕ=�ńY��m7�ڲwX>������]Z׵��)Q���{�Zɀs}SjzË%��'+}[x��l��pm�K#R.|�yE�7lL3l�r�dԦ�4zO�������fy���2�&g>t���)�`��z葰k8I=E�T�"R˸	�6���l@F�����𽥍�����hzeUGt��m+���M�$�ur��b�P����z�]i���������e�i�7L�=����V_#cc�5F�pH��%�3C;��}�k��WJ<Χ�k�CG:Q/�o��*&���}��dݙ3��v�M�j82���\L�&�nh#t�����M�g+�."K1��F]�X�F,γ`[RV:�g_a��Z{D	Ym�x
X_@�������92��\�!Ø�r���t��eA�T�R�Wr�`��.�S�E��؉wӷ;�Z�G5n���C7��H�)մ:�m����oQ�2'��E�[KRS���7��}n�����Y���݄�@z�2YI[����m��"�U�P�m��/JbU��y�Yܧ��U��D���UMs)e��2�����#��U��k�)���R�T�l���4�{�Q�U}����2��v�%h�(�v�+��~'w=n������\��KsP�����G�6{��w��j�	87�ux�X��/&��AR�q2�2dvum�{[	�e��hHE����$�qjM3��^�82�ˈ'݌��4tE4�4��_a~}}9+�0Q����X�Up����:� 9-H�q9�=���Uw4��"Հ��{y�}��s~=�EE�0b~qṸu��7��Uǅ�Q�.���x�l����m��J����n�&������v1fۍ��<:>��^����p���s�`gV�����4�1���:���.6*��z�\�8Vi��;2���pk)�8���k�܀�ǔubc)���2\�J1���\ L/�zy�1�K=wR@l�l�j=w��9��\�A	2 n��$ �o�t��k��;�ju��9�s��	�-��x���z�ļ0r�01�;kFYZ��U�\ 2Vm��wo�����W�!w�]>N��bc�k�[vrƗ�Z<�9.�U|��al�z	`�1�>��ob$��f�\)͏fܕ��EN�QQ����Գ��n�;�tL�����G�����UtŲ�{L�y��jﭺ�B=��U'�G/l���vA�8̜-���Qv��4���ySs�Ö-���ux cUF�"���5���mDF"1S)@V((��(��Qb"��3�R�"�(�(�QH��*2���J�*ɍb��TE�(�3M(����`��
��3)U]R�Q`�DTUUST�����h��
�DUkQER�f��&$��#iQ��e
1,S�4X��8�L�E����`����*�T@A����h�J3VJ1X����DT#�"�EER\�EEĪ�A��[D"%a���X��EڱYU5J"�QVj�բ�EQQT�U\J֨���
��Q� #QQcX��Da�R"
*20`��\e�����Ҩ�(�[j*�B�QUkj�*(娰c՘�im������8��!�LB��ܡQP&<���B"�&��k,ioFF����8�!�z��Qj��I�}VK�kb�Ҝ�ܶ���Ѝh�[�"�(�Ut�u>'�\�p�~VL\T4,�5�i����)�i��7{(z|To�P�;�P�&��
��]	��1�b��>U�z:dM��5�d�۱}�ԕgh�z�y���"�� <OG�N.�U'�#�#����8t����s����g�qS���^�P���<+n���@쎋�_Ӌ��M�QYWo����������3�V`7���7�y��aWO��:�):،�t�#�Xb�R����X��(2���L���Z�ݜ9��M�]3ca�28�N�Y{m��ڵ����W�lnony>f��o��؂�!�/��MP#�:���맠�ㅞ��h�ή^>��9V^^	u#���\lMy���aX�5�.V��d F\RvT>�����TGe���
/»��_C.��:E��V��̊o��Q���VD\��|SF�n��]��G�L������t��E��j���f+�ӂ��x�3��F�簕�z��}����(���8DA7��Y��ËoJLth_��O �;��H�rM���K��bfH�Lzc2_?i�_(������}J�h��k�{���5�SK��R��w*\�f�E��w�!��GS}���镥��d�	ŵw:�2k�K�-��X�yG�0�*�=;q���`)���7�:���k���/�}���=�ʇ,79�!����}�=�G��L��ώ٧X����<�^�8�(��H��_	´��Z�y�C�����aV��{m媚�o+[����K�^�Ҹ������
����H�򇗄��;��ܞ���CG��Sb�iV��ł�Q�b��2/ԩp �\͔3��[�}l+��Ǭ�v�]�����C�zF)e��C�-8�;J��򪊄{}�5m�̓�������B8u,KҘĘ�pо2��-��^�;���B�Ztx��o���3�b�8`��@F��:�e�P�eLU�P��n{z�� Q1@��^�!�Kt��>^���,{�?hc �$W@|4�,)/�58�s�q�i�J����t�HN8�P�M�ݭ�Z�	���	*aC�w;��9���|�|x��|��#/�TZM�;W�|`��;w�t�č)aWy���(���.m��uƤ9h�v��y;
x�8��MV���t�o��t�`e)�Kx�P�0en �g���l��m��k����S���ۤ���B���t�z�Ҿ�K�,�-ŀȠ�>nV��%�;��=q�05֗~�uoha��J#_�ƃ5Sn����8QCцm'��,�w���Zu<ۢB�პ��E���v!p�z���9�Z�1�����#��T��gP���8w��5���Sh\ E��`#tUu�f��'�B8x;��J�5}
D���A�w���#Qe�PU��o����󌑸qO�O)�(���x͝�)����u��U���+R�2�!P�B�b�:���:k��p�{dYF�1J�}+7�S܇*�.{JWU����6:�pc��{��]����$��5����ŀ�׆���F"��TF[�t�V�H�Y����^'�jd�c�����xGx�0�J�^wι�}�)jYa�_h�]�ОSQt��S�w}fo�i�Q顮}z�\ƌJ�ʌ۫3b�3Aɡ�UN�_Q��eH[���/$�X�J��:oiר(��J�n0_:�"�:f]�2���
i�J0�����T=]A��*\ì7C}ndwu(i/���n��^�nL�j�n"^WT��3-��ɶݝ� ��WPN���0@a(���nq��+fIik�b�*c�sM9R��j�b��ޢz�R���7[c���9*��]RV�"�p�O�`��Q���{��R�X�G��|-��N�z6���aJN�iU����9��O��D�V�DXV��YJ��b��=*.�^�zuCB��$��=ur��:�c�X�z!H���a�z��뤴`<~1ۜ`���9�a�}���E�,�C$�$��x@�S��*�0Xً�x�5�w��4MH���t��������um>���ZgEd�{P�]�K��<]6���˒(46���[�9 ��TM҉�}ͷJe9s#���@и���,��<��앧�+6|f�U'�޺��h��Y��]��Acu�t�T��p1�����}�.*J\fk�^Ҽ���q��xg��5c�I�*��ߛ��r�Q@g׎l�.Kk�����L�}v#Y����Aꞡ/����[�t�Y���^k!�n�&�OD�Clx�(3�:�M�W�����geq�o�զ��)�n��a�. �Mg��,7Y�<�$�dܧ�kӳ�ظ�Z�f�9fͷ(�}H����T`���Pw�:����kĪ�O�Ҥ���fZ�λC�G{[s��Y;2�Tj�X�ڏ�[ҳ3��Y�N
J��]ڢQ���՛򢛋��ܣw[�|�ߨw�t�fo�Y	ݖy��#�C�ZW-����uK���A-�4�7���w�+OIYе+[���4��q���=~}P}<�,�ƙzgL=TJ*����ݙ9�Ϋw$��ap1c�M��|k��j-z|�>�u<������,�>�/����f�$�0\��|�+��0.�����σmb7�_�~T�ǵf϶s�`
��Nw���i�ڙBF"NO�5p8�T�8o�8�;�|hW�dK��Ƙ����~��9ok��`O�!����ޜ+Q�s��*���1pvb��W�׼8�I껺I�f'��/�<`����^*Y�}6I�ґU�0��c�7��oj�޸����u�)J�,4E�(���)��84�U����j��=ml�r8�q��7���p4{{��Jzy����.�C�E���=�4{����x���j���� Y�}��b�LN�ԃ�3"��[�T����Ng�5�y�l�{����7�U���ީ���l[3���a��~�3��Ӧ�i�2����4Xز�3k#b_����Z�q=Y�h��
ww,x�m�۽S�YW�$��~��>zxW��Q���NX})KQ���;1�P�ij�S�l.��,T�F�}�D��ޫ���JޚJ�75DK��ǭ]>}��G��0o<SGam�/� (�u��u)ӰK�������ӞE�=O�� �!�zՑT��E���+���@���s㊻_q7�y��V���.+���K9��,�p>���'\c%-�,���)��6�^]@�.�c�Wֶ��_U���E?vR�."��,���v��*��6�V�xsNҩ�l�yJ>P���B���\�-Б�:�1��;
W��P��&8�Þ�C`kbA���=xbֺ�2E�Efe�9��� T`z_b�|r��h>�C|��Z�ގ�%|��Պ�����I����=9�<����c���YP��.�C=2Κ�F�x���B=qâ�!�vX����&�}Nx�e��M(BR�Z�\��� ���+�%iΚ���=6B�y �x�5Z�d���VE9=��9�B���H܈d2'�5�=�4�K��T|�KW:0���sQ"�U����z���¬�p�x{1ٙ�^��I���ttX�����":��j��H���x6/k�#z�7��ծRӞ��WC�r���dR�Z�u"���=�+���+ŃV���voo�����eaע���\[z�][�P�m�3Z�E����0%��w���Z�'{y5\yu�	�ޖ�)��f�%��+���w��#��q!0y:�����]���:����.N�ml�z�j>���*�g=�s�,���|`���e���s��ؖ��_��P`�t�mxj.�b���\�B5�5�=�(w�;+�Hu+�ڠ��`�V�}��o�|v��k!�Mh�.e���}z�>����g2u�N���7�mX��q��/&�	E��T'Bx�>o�Z�W�����P����u��+8�,¢�Їu��фl���[2E�N� [Fs*m�Rb��XB'6Y�LYjE���KJ#�ל��7�%�x58]j�q6�æ�[[�X�1����loU�+�� �]��3o9:7��"2�h�EgJ�l���+���]ƜӄPX�v+<�q���V�ݧ]�(>7&n���<��8��,
xj�����dj�J�f�ޜ�7�7u���=~�F���nOL���2mY�VL3Ϝ-�OQѕS�
�����6�����eި|*�[Զ��n��:YD�AP���,N���&Q�VĠ�yq=1T=����:��.�����V����e��]����hS*"�F�AԻ������WtV��^`��M�G�vx� g�ܮZ!4sX݋��I)zք�g{%�s��%*W���R=�96xt�S�;�L��j�VmN�e����f��W+��1�4�=ݚ�=���g^K��+Ou�*�sI�⾩�F��@��Qq�p�����օ��N~��f1���J�����`!�����$EC�X��J����u�U�l�5�*m�9OT�3����-}��ٺ��z�[�
0�5�_B{Q�Q���kX�D�7f�˰���v�z��E�r,�*��]�[/��Tڭv�U��7`�nn�k�p�lօ�:���x!Ҡ���o{�wu(jU�S�D'e���+[�����s:�{Ax��
�
5(�C>C	��"���cD�8�Y��Z�2��D������cԶQ���G�4��\�U�j��P?b�ޕ����ʵ)��n����t#7F�YU����F�,���0x�PP�#�3rb�9¨ub�<�k���ǎ�������믲�p�kPs}�ԳU�,�Zɗ���Ү�в���{/��IXanX�(oE�͋Xq�2�f�+ɐ�ܺ��8�E`Χq&��]a��b��+���8݆TNx�,A�lmvBڞ=C2��yLP��!YS)P��Q��S#7gЎD�#����a?�,X��탻�0�Ae������tG����dFj�f�3����_�r� �v�a��'�T��~�p��:�𺲒��y�~(�
|��d>���������yx�z��	Ŗx`!��Y���;��ج[�0��o��N����zl���xԶ~��;$:qM�a
��䈄,>��O��o48�w��6j91K����޽�Uv؛k���\1��iM��zK˚��ޗK�X�w'�vl;�:lGN
ۇtr2��9��=�8%��=m�����%�xWl�.��>P8ixi��빜�|S��ʲ�!dҕP��t�'��c�z刦��i#�mx�Z�>5Yρ�c/$`���d��z�:�b���j���Ǻ��@�;���7s3Sш���ZK��B��S��j����/�q�f��������jQ��)?|�V�����ّ��}hi�R��!d���py��A=gp��ޞ�y=5�ߝ4���	O Bl��R]z�P�t��ؽ��:�z�A���#�²��զz[v��A�L�0��z������/b�u�e"�����W�2A.��uS��|Gv��(|@.�j8�݉7e��B�6�'��}&��g�#�Rf5IZ��˾)۬�T��Cws3�+3`�5���$��`],oypTk�B/8^}nީkq�u���)��w����]�\灗Е}�M'�Z7ZecbV����}�b�Wkȼ�(E㍼�N$Vڬ�n���0RvM��b��l��Ι�ϻ���g��Ѣ󟣯(M��n�zr�	loq���j+F�S��Օ�r�a����c�lĆ�m��ٻY^�n�eC<�8�/���=��h�k�Ex,y��nm�9C!=w�V�jc�`ƶ��)��:�'x��T��+3R76�<|���������S]yk������ݢT^w��+"��L��h��;^[i'�2x;�˵K/���I^�w>�
X�U��rE1�I�Ď�Ӷ��o�̘]ۚ��s~��m���5�QeL��?�|'Kqx���>w���z(�=�%��^����68��T��Y���f{����ng�}�B��`IO�IO�$ I,	!I��IO�BH@��	!I��IO�!$ I?���$�bB���$��$ I,	!I�BH@�RB������$��$�	'�!$ I?�	!I��B��	!I��(+$�k?[?M`s�0
 ��d��I>sx�R IRH�QJ)%Q��5�� [RBM�YJ�UU%)5Ej��!TT��� QV��*A�P��	SmoF�(�h��U�,����3�\Sd����ʭ)46�k�m)����v����ݣ�Z�e�6�)�����ԭ�[6�PF[��se�P�e��aJY�m�#lkb֢0�J���e��F��X��fXڙ��[3kZ�j�jV�j�Š�ɨ����ٶ-�fٴ1Y�ZkL5��  ���P-�4ݙ@��6JkT���S@4�k-�H��3h)�0�
&٦mfR��V�;f��@��ҩB��:�V�fRw59�mP��   v=�Ƃ��[t��F�V�խ�v��텫�)�m�n�ك�V�(�ۀ-��ػ����SN�piֲ�V����H)ee�kYKj��m��/   �� �B�
(�y�(P�CCB�9{�Т� hP�Zu�P�  �Pg�^�@ �B�
{ڷ��B�
��<f�
 �G��f��W-g\ 
S��u���ѥm�\��3f��-��-��  �ʪW�5��m��r�a��T Ww.�����Қ�Si�wB�t�MWs�*�5��v�I��r��
MM@�m��6�wT�+kU1�2�K�  <=�4��ks���Ҵ�GR�i������ -�ٝ͐nݶ�St��E+��r��բ�S( �M�5r�J
�m��5ZV2]�ڵ���h��e����   9��ZŷA�ZԲu��*Ps\ �*���p������6�s�)�5m*ړ�Zj�wkN�i��n����a���hm�ٶ�
l�d�   �;����֩w2�`[i%'r�@�v�T��˸ +�w+r�,e1���BPέ�u�k[��.� ��j��Vd��%�l#5d�UM�  ^Uz5T])�ٔڜ��;e�j�C��C�h���r��n (F��Ӫ�Zv�j�44�Vu��mVZX`�f����  ;s�R�sk����fWc�`p��C`]v��U٥��t(�kk�W*ڎ78)F�������\�[`Yl�jI�6��ե)�*�T  ۞Z�e5 U[��T��$�J`)E�����(n��].�tj�Gv�p;`�E�m�:҉����@eIT� ��F�Oh�JR�  ��hʤ��OS@4 E?�)�F�0L	����`$�D'�JQ� ������}���j���Z����x����_]���O���V&��� =��z?�|����$�	'�! ����B�� �$��$$ I @$$?~�?��_�7_�Ҷ�� "�/2��N�0nժ�Z��"��!d����V5��=�u��2�Jx㤍��v���\I$���%��ɥ�1]f�w���l^��]�렲�3���Z����J<Ԫ����oyV����I��"(�a������9��_bFc(�3w[D�(����lVⰅ"�3o�tÛ+//6��:Ee+Ö��{(�֝%�X�rn-Ա[�E�%3Z��Tc2%�bF&w	��
�%JZ�ivf��4M���jd�� -���V�Q1���;E0x�$���09WX��[B\X/LH��p�/0�-d���zO�j�;��K�P�[Kh�ʛ@�b�	i�n�i��v6���W ���9N�8��,RD^i9CX�f[9��"�I�:ʱ���|n�F33>��'Od�k3�>ٗv��6�(C�ϐ���ӵ�+(e=ڟl{��0ǲ���YԂ�PԌ�Wi�3iIl3g%�엎Z�@J
����e���H)�$�1��ъ�Ը�h�BT���k�W�ݍ
�9Wi�k�"--2� P*ҧ�[�e$�I�%Y"�h,j�f,yە&Z�RT���lB��2.r;�j�;�^����D^4���hTJ�!,�{�l��˴�(�3������\2�R��啫p�\�>4^���7��mAW���	�c,Gu�}�K�v��0ͥ����N��a���^6�S�7���C+܊��E���x�@#�І��Z&j&�LT�6�=�xe�`�
-��.����s.:�DTs\�l*9aؚԣ��`Y�M��V�\Xˠue�Lre�*�wt)��M���Ľ��k6bXتe�1R��%��kA&�����V�6/9�&�V�8Cv�<KkV�,L�"��������իF��p$RI@�l���Z��	�~ ��6���mc�'o�A�d��.�:;�f�X��l�&���i���!$�$�63hS��l�qk�o�EԬL!�-����v��m�,*��]=T�������㷐ۛ&w�^*��
p"���w$/n�y���KT{(����/.6�'�)j/jșbf��������Y����5E���xi�qw+_�
n��wNX	L�Lw�k1��_ԧB�q+����S�-��ö[ǲ�%[g�Ǖ��J�][K2���M[1ٻZ!�R�I��Y�C�D\��vu�$1�*Xo��W4���ݵ�^��7��)����9{B]�d*�r���@�Ѣ\D*��h]�J�z�ȷi�2�Ĩ����l3if���֜�N�7��!�2�<���hҳv�컡
��n���o5�d�'�bp�%0��A��6�k)�+Mŧ5��i\�"Z)���Q]Q0*� 85��.�&��)����bGvc����aӎ�-'"�9�6�M��^�Ƭ�f �X�eb������d���!
ѡf�����LjF�eK@ۺ��T���N�*H�v
�]@�0���N��m��V��?�5�zU��5��\eK�>V2v޽�7
��X��Ctj�6�F��PX�TVk)J�cSv���J�r0��)c�Upm wP�(�CJ��'��0j`���f�2	��6f�h�k+f]Y+Ӣ��D�V�ѵWn̄�-8ݫL�p$�x��M���S�����D�Xh���Kѹ�+"o2��� k��	;�� �Z�/n#X�Z�9h(N:��1��zj+k.��z�['.� F�N^&#�ѕ��m�,f�F�M�L�h��]��(ދ��b�KΒܼc3-���MB�V�2S�IA���Z�(I-��WwP֧MkY,��F��������ۙ�.�[��vp�͌h.^v�ǋ+n�����G7k	����kͪɨ՘���s�wV��C^��-�	��l��P�Ylw�$�˕ё������M���O`[�QQ��sbj�Y pn�,S��OTb�:�����(��Ū���?����#2���ɔ|�y�3{�V�6ي�{��h�@����4�T�+�l�!:�Ƭ�A�y�̣�f!>�[X��I�F�{f� i	V��*A,Ccc���Xc"N����'F�Uֺg[*�;�^��އr!`�F��3i��Y�ָ������C�"ǳ7�˩į�R���
dBT.a_n�պ(֌��&ai=d41�V�ua7Z�kt��T5f��x�ث����;��pl��bƺ\�3���W�4[D�.�ɇT�l�m5j�Lʈ�.������M����V�z�m�*�ī��T���PUˊ�XA�ёa��5N픶ks+pѸV�ت�]ՋǠɮ�f�/P�S�yr�����AlK
͘�E ۨ���A�,��W�5�&BB�����koDō1�7\�5�P5z-(N�Vi���k	�x�T�i�����H�{N<�妲�"l�M��7tVܨhB�$Q\�V���,�I�X3𳠝���M��
E]�-�{X��cVE����Kڅ�&��U�t5
����mYZQssi
��	a�Lʼ/rۉ�#Bt�[�j���љ��/콚�d�����^��[&ؼSm�[:V�o 8�PCa�c+ ݶw*�M����)�u��,Lkf�`�veّF�G2帥�z��4�]���%��h�\��滿�1+M� �D쨮�+�����ub��5�fE�W�ܷ�"-R�ZĈ�0BH(�؃XS��La�9��9��yN�i�3�.�ݫ�k�{�m��[���ę�	��ύ�*m�z�Kb����v�Z���4����)Pb����C�E���w �����ݏ\�����Y)IB�s��94J�cz����z�f�?��zv�<�̺ʹB�����ɤ+S�Mi�af�X3>A����%���@&���a�U��+S`)l�Pm�j�ׂ�U�9B�<wF� �e����i��DF��(1A��-�ѧsE�ZMi��vu��_�=��_-GoN�GZ����9�,�Qw2�ՠ��#e��/�۹f�Y��f�*Й��	V��`�
�"x�f-hI6'�S@��h���@<;��wO�ƣ��l�Hh./�R����ej�Ԡ)�϶�F��&���M�l��vTRGr��-[5��Z�X���^D켽f��;d�[Y��{����E�򻉻E��Q���l]�J����Jұ����YTL�u
����fj֍@ʩ��(�m՚ڵ���wncŧN
�h�h���[�֍n����+.+�7^"��!�ݙ�����Pgmֲ����a-�Z�T�l�	n4�VX[��Y!L[�r#e�[�Py�S6�;�67kb��ȱ���n�s��'i}6� ���N�-ҪXb�K�3eT�y���Q�͊N^�2��,"�X�N��ԜY������^1K#�p�ݎ�(�MIg��YVZo�)b�Jʰ�b��BYvf�3+j�x��9He�FA��в��D^n�ڶ��
#	r��#r�"/fD��f ^ᬵM��vb�j�ፐ"�@�lQ�ص����$智�������1f��	��Ѽ��eKC����2��`i��J�v���+0ʗ/6 �Tw���G&�Y�^85�t�VԳ(k��V��R4
c`���r��ZB��=G>�,�3�퇖�y�U&ӂ��F�-��w�A�+wQ��WIQ�ʕ�r�"V�
"mmڷV&+��ҕh"H%!#wYy�7j@�$�	��5��R`���[Xh�Q�5��$p�#4�y�aw�Ŝ�3;xnؤ�r�6��nV�g0n��P2�eM#��2�R6�ѓp����
ۡQӘÙAҗfj\�o6Tl �F`"���:��H����h�]�3 ��`Ѥ���q�oqGi�s1�a۲���D���`]�:�Mkf�i��ʽ���\�1Xt�^�p�2V�7������cJTȠ��9y�6��sv���zРD[��d��h.�f�N�N[���Q�z�i�KQ��SvU�m�o[�/.��9��n�2T�D���d#��K,̘���F��+�B���)̨�H$t�*��7 �T��*7!�-�[5P��I��-�M@u��˒&D�s.�6��6i�5��Vǘ5S�hە�B@|���ִ:b�Hj婭��:2S�ի-S����
Z�E�42m]��� cMj	m�@�xr��1*���nVd�u�I'R��g����w� �A�cY%*WeԻ�	�5���[]ެ5��;םÆgB�]Y<h��b�2�Fd�S&�����n��VB�k�2�a���zUm�6���k	Y��%kY�eֻ�� Րֈ�&�f��D����D�����M͏��ނ(��Kx�bR^�l����2�*9P�}��
o�!��(�)ek�e8N��ʊ��XzF4o`��iۨ�q�r�h;j·�*c̘��s/2u�Sp]avV7�0���$�
"-9�D{/!˽�&��RT��� ި�G��u�g�4���V�ͭ��s�5'������H��U�9��j��D0��Ba�iXmL������k�kH�kuly)4	{y����Ja�D(b�-����o
P*�fL��V8�fkNaX�E��5r銘3`�z�i*���iJ�Yh=���p)+t��.�1eŃ�f�SM+�n��K�Jg�Bt^L��m����`�[d���W)��eʼ��&��@�f�����(LD�֤dK�d6�͗����3,���j�V��&�e�6Zy���U�Q�:2��l9Ye���ũH+t�k8��[Ϭ����0�᫱!
��MU�V�f��(�8�`��$��aAe��M�)�5��omԬ�QI���;�.�����z!��M$/U\l`԰���c�V^1�Op��G��c@���V�(�V�u���hu<�y[��k":�VZ��0 �c���*�BC��!��n�g=��ש�˺�����uvP�)��լ�r�F�� �$�t�d��bP��Z��Ҡ,a�1��xth������Q��:d�% ڢ-B�u����a3pQ�)��KH�u�y�C.ŧH4��	�.�8�m��:��[;���D-����	a�y�X���v��v^��v�AU�ͦ�l�A�
hT��00��sM�enk�ut�5E��U�=��W{ga�+$P���-ݘF�+���ܣr��7��5Ō#�P!���B`y�n1YA�vaGk7�=�H-��h�LQ��姀��]����]�K���:�P3C��Ϙ�>�OQ�!�3(��}���ɉb:��e�6m�	��q]7��H�ګ���5�6B��E��R�%�y�ޑͲX��53fM���(r�7�m��F� �9HX����l�h�������2��[��hQ�[�*�Xm��jqE+@y��s�.=.�Kax��E^ggz����2��hTtS%�S��nQ��#�km�Ԥz�����.�:k(,�ۖ���w�(im۬{n��+k.�����
!cF���F�ÚE�a2���{��a�Yz�B��iܚ�5�IM����xn��� ��q�FFt���dٯUFʹq����v�J�g
-�]г���Q}�uʔ$R��bOt�{N��]�I2	 f���أ��[��
�j�[�!57n�m�^,ӎ��U�^;�X�䡃���s\.�L�����ۉ�[�O3*�H��i�9I�\;ZE������a{B��a6iQ:J�μN1��KWt��N�1D��G�Z�&m"3s6�[�QD�;�.�	-���xbU(�`�������n��9�B)�0*uv��A�A�2�kɎRY�k]/�0`Q�F,�U�sB�"V�(f��[�J5b^D�Y��e ^Jͱɳ#�(V��1y�h���ɩ�<2W���j�}*=w�k6^�t����TU���.�+_�k
їeX�&�b6�l��ۥ���D�8�YY�`�x��kmU���Úɻ�ū+,�+n�Ò(W��O%�h��\�Do4A5Yg3 /ܸ�Y�&rJ�ؤ$�y2����nض$(!� ��Sj�c�Fd�������iްUfƽw�fc�4�h�s\*R��f��ZĒy#aԕ�7H�^��F�ݙ�h�$h"�Ӥ�r��fTU&[�� ;��է ��$][B������52��m	W�8(�T[y���lC7-AX{[�m�H�e��#�q��ʻѲM�%�
���]R֯sr�`�OЄj�5j���8�92�7,����0 v���e�K&ռ��U^���R�������Kc_]�l��pT�j����8�ƷI�v˴V�:�XqC��Oj����Ւ��L�n��A4��D⣵�4EbÎg�B�9���u��h�X�&OR��� ���Vp4�8ɣ�L��3*h*���y{CkRp��m�N�XB�v�̏e��h6iTq�Qŷ�v�{Y`/fټ�[Ү��% �OV�B�-���ѩ��g�'�"�7BlŠ�m�&�6��55cA\'!�Q�W�m$3N�M��^I�ZM8/j�cʬ�+-��rBP̲��O]�Cng �F�ʔ�B�1�cE��'N�r��5#�f��Z�u��L
e�Z�$ͬ.�Ƭ�CL�7ṆXjǎU��g��]��._�y��)#�Xh���IFh`Ī��W����s��c� �Y@��F����!���lT�N�#]\�̫�ײ����wI�s�z�����[zY�t��-
HhA���;%�]�%����r:q'v�$�k��Ϙ��ؽ�WHY��^2.����䙓a��:j|��"t9u�c��E<�K8�
jM1�a�V�TJ��U�5i�I��;{9!ͦq��q+Af�Y���z��i��5)ZA5�K�m�5&���0����1S��V��B�p�P��o8V���:��áV���w����x�Y�����}��Kw�b[ܵV	C/s��7*�l-gqm�j����w�c�9n��!Ѧ����p�:��(�t�2��fTƝ90pV)��((Gv����R���қ��e��y(XWͦ�z�^��bYKV� p�	tVr�Y�z֒V��LJ�# ��l��^(b���TG%�V�l.��H��83:�7��V�\o��ը�bQK47����"��2����p����]��ӏ�(�׷�]���S�G��(>t�c�-�����ڷ�t��Z��V�!2����6N��:��/$뛀�S��M�����c�8�#����V�@Uu�Ʈ��7�Y��2Y؜�������͡���^��Wz֟z"�}y1���L���� 0�뢥���}[��ꇖG��e���}�]9��x_��З��^h���}�-]��#Xo7�J��Ќ|�*�˽��T\�S7�w�J\���)�b��Y�}�g���4X]"�]�q����p�L|�4X]\q6�
����B�t�A|+,wuL�� ��V֦��L���ab�H�>���ܾV�eA�l�#���5Y�L8G>rW][War]4;y-% �Z�ʌTʚ+e������y1ɺ��v$�����Z<\��t�f��Z�ޚ��^������	&��j�3oz���
�Ex�_wrÌ,�jsT�c| xn��Ws� Z���=9`B�˭�EA��w�l5�����OZB�βثe�8W5�a�f�������
�#dV�+�ܥ���j��PyZ5^f6;�/�\�}�.����w	]/���qh�ͷ}�ΐ��%T�z`Ykb�Z�d��zӧ����=z	[K4��7[�[�]J� &�ȹR��m��UɆn�ˢ�'�J=�w3�����Ԕ�@A��&XEh:�6'�eM��]��t.kqǝ)�橏KK�K�_��qԉW�F�a��ˊ1؃����-i'C��$ŷ�J\�8�"�Pi�X�s����m����3J�o]n����h1�*��a�c�U�	嵫��:�x���9\o�͓&�f��v���� ��N�Lܬ�Σ]q�����{��[��f`��5G��ht̩l%w�^wm�f��陡͖�q��d8°���އ0Z�ơ����S[o)b��ps>u����!�(dzS�u�J�ǤOo���%M<b�g�>;ti�x3��k�fR����`̣�n(������i���9�f��M�(b,9+b7yO;F.��sۙUc�	���b�����6���5J���}��0��*�e#�޹�wR��'lt��Bi�k���{�����YE@\�׮.۾�
0d=*������*w)t�H��j�����Ų\�s�&�;@����hxz����Y:�Z,�=Ի��ҹ�1�Ӛ����eaӰ�譗Q�qӦI�o2f�υhq���B��M���%�㹲��f�����Z��R;g�-6X��9��}�i�%�A��J�\;�14�A��)Պ�V�ݗ����;B��o:�b[�bz��)e��d���=ڴ�nj�d��w�zuf�Wֈ��/`�2���i�R�\n(�И�(*�{�.4����&��Y��BY��P�~�V�ơȸ�4����8^VfS�؅�t���s������.r9�m���W�h�j�J��t�uZ�jWN�z�N���N�˰�L|���.V{_ֈ�\���c�h�٢��\�U�B�f��ņ �.���_.���4L	�l��E������n-��^r�r���2�� ���x'e:8y���Z�D����|���p釓��
�{� ~8���5	���,P�	󧣂��3nOT�qn�����G�2�Ö��f�Œ)oN�Y\�Ke�v�1ؽ��f3�����)]�����(9�+��.��1j3���>�&���ˑv�;�_m�SHt���Y��Z=�gn�2��y���^��ǀ�IW+��ո�M��6���ɽ��݋�����r�g2JpX���Tk�V=�捳��y������O��@V*V_C�u���:��u���d�s̨�+|z�t�w�����x�4�c�F�:��9�7T���Aɾ��������~Q�MgP�KX%�0*��˷9���n�B]��.Q��M<���Yб�OtoU=	[��˶�8�T�hg�c8+L5�ꢵ�+
��h@:{��u�8#��*�V�ÐXغ��Z�z�4=V�V	�Θ��ÙN=���r�S;JԠ�Y�7�r1r���<�'l�ʽg�f�z�a�#�G�-2Z/��%��N�v�E&Ùk��h ��.OTh��&�̮�/��a�@q�b�m�b��C��e�|��'/u�/.�sC.�$m��F���h�'E¬V��:t��ECFN�-�]/Xsl=��e�O3�O6��@����s����Jwh��6RC�u4 -��#����I.���
��!��I���C���Cݘ��.��Uc_ٍ�Y�0�R={PY��a��R�^J��I�bV�E4����֝;�1DŸ�w�Gl��Ƙ>�,u�����˷ol�Mi�m���S��C]�0X���9�q����F���n�f��T�`�Qܳh�N�����S�)�or��J��a�Sh��ZMY������t���F�=t�&z5��s��sSu��JLw��4K"���(��!�{C���n_]��N(���3(cmI��T��]�G:v�j�%Ȩɤ��m֪�z�^`m��~`Q9�v���@Ӝ`��zpV�J1�i�ʹ��O����ٻy�VI�-;�QſD���/n.O�h�z\�[��Ӎ:��Uʖ��.֞#��T�}�.�]X�
M(_L;�;�*�NN�6���^i0����3��+Ub����h=Ge��Y�YY��.
� ���^��a0�笷(a��(c��l����6��s.�r�|*i0]Fbm��s��Ŗ��\̬IQ������'�o8햶��'wؖ���R�PK�����<{Q"�����g+f���:�H�ԏ��ad��[��Su距/����g`�'v_Մ�M4�#�Q�����~Ѥ�hX��V�e�u� w1&L����SHLmV�q�7FV8�����:�a�!:�f��n
���Mt�>�����	q9��I����as[��H40OY��B�":L��	���2���R�HvF�Jbsj���gFE/@�u�x-��gJ;�]�E�ZW	֩W��n����X���"��Ov�(vo!\���ˬ�؂b�-��J�e`/_dL�Yv�m�%0��OV�G�L+g#��ů6C&�
��g�fjq{u��Y#+��LF�5+�ũ�r\�Z�P*��%aYҒ �h�X̤DY����v�)E�h�ƪV�.���X��<Τ��jR9��1p�t'��������K�vn����,��=�T������޾�f��#j��Y�fI���>x�:Rd��v�Q�z��kst컊f�֎�bR�~����{^-����5���s�18}Y�#Y��K���F+�k��ҚέP�y����W�������rȯD0�H��b��tw)�M���t�>���h����W�Y��.�۳5��:�d�(A�7����ڡ��9&�P�J��om_��sY��v��[��������TH������X#x-�<!�B����p7���ѝ�\��B�Z���S�+''G��)dF�-p_SߘI����LY�z5b6��������ESVŽ
�VM�!��v޲���@l�v�3����P�������klK��h8z;�u[�ٰT,�;m��-�ޗZ�h3aL��v�N��<�S\���O��gVLHj�X��!���vuK�U�7�1^.�ў�ƫ���Qʻee<�8V\І�+�~IR�}�ٺr]��b���в扜B�W�"����ú(ă)��,�+�v��ֲ��u��G�\DZ�C(�w�lx�A}a�;�e�9t�R��w��kkxڃ=���u���#;l�pI�,)�h����*����7If� z���(	7˃�HG�)�*�_��v\|g,i۫z��ZLu؆9���΢�7�-W,{Q�vц��Tt+?.0�Kt�v*��v�`,W��#	�/ON�ԤEM7s��9�j�`@]�<�=)a��v�x�P�ɣ��3��J�i�LO(M�������Dh<v�Գ�?t�}�9cpSQCF�Ó�Ԙ���-�D�v�{HU��o;�:W%��(�]��˱�g
�2��(k�L�҈�w)�8����U��°�v⫉�9����p[�ȕ�E���P�Z� 월k�ǋ��s�b��m=��|y�3	��X:�vY�m&1#(�*b�7�⬳�G@g�J��U����f��C,�=LN���,bW"�Э�/�(�ݦU`���pK�~��ʋ�4^�Xn���16:s��9E��1PMX���1�^s;���f��PT<��[M�;�r�:��j�HbVst�w�#�k]�.A�p��7���6��^/���U��¾����%q�6�Z�0�A.M`�+���ɛqh+�'�Ua�/���(jȚ6UI�@�Ѷ��cq|;hn,G̥N�����Pp��Jr9v;K�/�+ML�w0Y���F�a������S1�������`�u�UT�V��l�����ad=���i���\�DV�6phD�6���t���$;�����20�jH�i�����.����;@��x�6�r�E�����2aܴS�](��	��e�Cε ��
VZ��-��U�L�A7D�f����Y�����n_l���f<�~�<3�9�� )�az��ߑв��s�S2hx���-�K�G;::�^,������m�n�b���C��Y9�g
.>)wز�kG#N�-;U�i)��q���y��E�6j�@�/�L�e�̕F4��+�V8^iDn�Z���U��{�s-�4�M
��QW���n�rZ��<���I�n>(S�6���7d"�Aw�&i��\�u��V`�D��t�ͤ�VK-�é��q�F�굁�k;�շ�Г	ç Doa���`�62�����U��z���ju8�O��ʴ�1̵�[t^e�������T�- Xs�eGS{J�>	��R��4$�v;�fJ���AM�[ru5u�@�C�Fӭ4>�{C�fMgp)������Z�������c�wMv�w8Rcq���[�:���b�I
U�k����{B�s���:�\�t��{�a�t�e���w���m����8��vΐ���/�w���$
��ȷ�sr��z��9�n��0����9#n���������������ЬT%�B�\�C[��+t�IW����^!Ճ�9���fA����OZgz�0;\���J�1k��E��a���jԈ����8͞va�lQ�����.RK!	P��p7��b�Ap��8fq�p��/��KYG��3�r$ո�3|����CG�<K2ܺ�faz0�uǷ1�^���8��if��
��OO��}n�aO�70��|Sjƹ�c9mԖ�w��p�n����u�&�$��S�u��Al�%{���7Ӻ��;���pE鋅��sOiׯ�
r��1��N��:ͦ��}����͙�T��Ur39+���k`���]��LYS�m�1c�8^�;i1Q՜�C+����)*٨>�������uN�k]7�iֱ@�;b	q��,m{v�7������3�r
�o���̎fϦT�Z:���ؚ�����7���\���{��+��X��lH�9i�yt�X�+��v�Β�)趱�rfq��q���-N���Np�x�y�7Η�����e;��%�˧a���ʶ��|c2ed���J�й �t��Y�����J��B-�~x�p
J���	ܗ��ւ����V�}��*5�
I��9��E<ڪ*���v��k_8�j�L?�����γfN�춵o�g1�q�厈CP��	��Ы��0�үP�VXyW]w�s�cq�F[̖��P"�$v �T�|���+��Y`1���X�ZAu�X�`�e���hd��4jMv�we�9[IbɇPk�$ӭ��ǈ���Җ�Z9�oa��۳5��b�]�e�Q����~YN�V���%L�� 2��u�����#b���	�F�]�����bN��J�[eAcm���@<��m�ϱ�B�Bk��xYy��u��E�J��e;����Y��qqe^n��g[R��u��wHʮpiٍ�U�Y��4�Z�.�0�W�P�x�oy���3�[�^�	�ߦ^=)��{��,��8_t��d�-�mq�i���䋧:Ɩ����".���{͡��Y[�ơe�xn�W�2Yˁ�L*�D�q�{�-�K$Nh\���3d{l�:�Z���ʷņ�[ul�hU�D�N^�%�&�����j�7]2;ϸ�J�t��sU��p�ʼ<!�<�k�������H		�$$ I7�_�w�5u�N��*<f][���涬qi�[�1�H�/j&(<�|���G�=��ڥmk{:�8bP=2�����K/�L�v+��Jذ�v��������MX�v�Y P ?�!�V>$�k"c���#��Z�dH�(�AJ�+F�����c�-���XG'^�g%ܫ��ǥ��h5x�+�bAʬ���r����|�s�b�Z��:6�t񬘏nqY�����q�0.�,�}�Ykhh!�S��9�mG�wd&y�P�X�v��%ga-��T�q�cXʷyrs5����a\�1�I���[[N���C�ܻ�H]()M��]6툪^ʱ�A��0�]�V�WAfZ�B�&_[kn��2���Ò*ɷ�b�"���y��,k,����_f.����4���u�MdT�ҙ]�n�'`�= ��ec
�!+j�nP�Aah���Q��;0�Y*�
����]���ɨ��vk�\�Yx1;IpYwZ�R��D�Yo3iZ��!��XB�Y�
4�@~�Q3�����ΗJ�٬�y�c�Ѽ�9&��Qօ�BoQ�:e -�s����敋m��AA-��Lֱȩ�gr�]s����]u]{VeϞ<�RQY+i�e*;O��{vͷn�����e�:uv:ǲJx�v;|�'�8B�|6��������ʹC�gg&�Ő���Y��*S�X0�SD�]i�k�v(��'y��v���r�19���@�Vk�ؔ"�8�#�vL��k����h�~ء����-��T6�L[����1�Z�)�ۥ �^���Z8�]�`�cL��T!�v\����T��㍭���_j��c�#)g!�A��v��4�RC8QQZ4��$��Q���Vv�\��e|/��#k�-W��Q��%�� ڑvW,���!$U[ƚz�P�Y���3���Jĉ�hvqD�X�KX&b���"���Lǝ�T��\��l�{��}nШ`y��o����~Ꝺ6�u�S�ܸ&��^K�T�0���^K4�喠0�ɕ��R�X!�F��	�!�ٕ�;Vcؖ)����|pRuاw�4��ĩb���mу��텼{f��:bc����� �̥��2�P֪�]�b:�N3i].������gjd�5��Gk3ie$�M�"ǉr�X��yk�;����ϯq��ɸe@�n��
	vαY�{��%��c�\�^�֩�'.��lfr|�)n�tаm�r4ch�����b�S�t}W��s�)����i�H�s� Ruδ�嗙��*���)�N��R��b��XRK/b�v�7Q��S-�7��vm�Ej�s���1���7���$�-��Q�vF��%�呌�Ӊ��f�m5�:Uz�5WB��ݧI��4)���Y��ѹ�fM~�BZ+����ֺ�^���r�@`X�d��a��
��͗`^.p�R����rl�q��)Y\�8����͸2���wz�35�47�����;�匾Ր��A\�,��w��aH��2��]cV� r���ѥ�ɇl��q��i�����7
VfU�-��ZZfN���h9��rR����U�G"Ũul��Fh=��B�{lG\��B�Bw���]K=9;�l�['n���s:�V��]˛i�n ֤���$�ѐ�x&&�S'��;,K`��*޹t�VWA%�b�L�3�Wr��aFܒ�{�K�Z(�����n)U��\e��Vo;d�Dwjhs���7��\��yx{)��X�px2�6�\۵�U�3i��YD:��J֎�[Y��[X��-�\�we�CJ7�:�tN���;�	u̹������=xݽ\��6����B�<��Ч6���|sd�L
���'���1s]7�//0��{����r�_Lܺ܎�7Y�r�Ō�o"�b�<��g��n�7�s��Eq�
��u�,��v��W��O����#ӹ-K3[�c!�h�{ �7 ce�N�aǚ�)��0��v�}N���9��:[��mj.��ʼ��:9U;�lwZ�Eq�ם������[\�����δ��9P�y��A٥�X�9CƦ	��b��[��֜��T�N�i�����'�9�Y(����[��
��I�ez�SdHsFX�ґ�*�n14ne;IeB�@�j�2����p�l��^�t-��mŔ5�\k�n���&��T�5�7{
���έv�Zn�:i_+(�ah��3*(�`�vuqUq��*;*�9���%�WY�j.�Y����JV��ܷ�ݽ�Ϳ��g�gj���*Tl!�u���Wn���8)��+�I\�u�����s�������pg����2�Y��v��>{�4]D,kG2�ۉ4O1xؠS�K�Y�XY��:�[��ۊР�d�7r�����{`��n�Ro��y!JX��z�{�j���Pew�x���ft��\U>Bbr�]�y��Y]��bO�U��b�靥�E��)x��n�P��x;'�[:s�uc58`%���MD�*d��Y��f���84�ɔtZ"�3勲�=�R�����-�j��-h���6Z"�g4.!����s[�b۾�hR��DMZ�ݗ�	�$�&u��[��"�auo�PV�R`�q9�dݚ��p�b��;ȴ2]����+��l�2�tM��2%�+p��ݙ���P����iq�˴��(�A���sr�ѣ��zOg�霫�ݮ�둁_9K���p�V�b�3�9]yW/�T���z�X�U�:g>�/t+.�����򏨡��-�X<
��F��_��ZUZ��E��ѕ;6��G+PC6�ۦ��n��9���\}a̼�.^d�E{��ţ�Mn�Ŝ�텆���,�Ü�ve��)��6�=���A��N�ʋ�<�{t>Ook�mXA�8�t{�V�1�W%w���ó�S��U ��c���:z���5(j�eϢWRFXߺ�B��p�P;Yu��~���,u*�.��M쓍f�p�6;. {.���xpcݞ1�h,��On�[pL.�u�烝-��˚��r5�9[���_'�@�)�3�CpfBe`eٷ]t�mKt������E�Pѻ����v������U����덧�zP�pu��)H�#�o$6��m1���S�u��ʅ7/S�X�m�<��4�T���u��:^��(�nh�Mhrb��%��
͆ج�n>y�����2�H��|*��vm������4.i��sǛjѷ.�5�}��E�g���"���{������4[9J�IT��>����+���q�U��lZ!���ڔ���'��ƴ��'
L	X�]�c/P��zkd�P���|��+<�й���cT�.���']���k%\ef{9��Ai�U�M|��˾6k[h�R�d�͡5�S��5T]H��/�fn=��"�м�5&3R��)�h*�I�T0t��ח��H��0�+!K��}q����N+T�- ��;%�)s�����R�bd�(�oGb��p��<u�t|�����D^��k��yR�]��#��:�mi�.C����U�U��f��\]��璋�"�F�YO�u�w�\.���A�6�*r�)U�!@�e�yI��9S�jƺ��oB��å�0��'�y��T���Ϊ��Wbή� ��
D�O����˺n�tG��]�LZ�cO3���(�x�SF_v�w9����ٻ�nK��c���\�pa�M��ᜧ��hoV�.�'�F^����W+��D�5���ҙ��Y���^r���u��B�>	B��8�
-;+5M���&���]�p�O&�Yډ�9):a:2��t#�,b�w�P�ـ�vT5�a�F9�@�&1�vG.�Ei/� N�{;-	�yp+�N�B{L�Β�kl4E��-7}u��&h����8�d���l�Z��t�cv�gn�B�E���5d��:��QS��C��=�GL&	H���ǵ;�J�C4c	d��^�e�zhhU�^��M��爿I\oj�ٻ34� ��c��g�.\��Խ��#ܽ{ɯ��摛���6n�謒I	��w� ���{P���ӣ�ٲD�`>�`i��S=9��}�%�h����k{pf	�8h����'���	/��{�Y����m��Z���hp��X��S����b~��*������2�o\���k�^a\��D�_���Z�\r�X,��G���[��U\��)<,ݰ팫��B�9i�bN�3oX�$	|4"k7�_U��]�J{�} 6N��z��QPY�8�;m�%��C��t{�eCCH�S65g�4�:�K���اhO���:�l,�[�[�!�D�V���OQ�м4!�2��O*vo��r@�`��|���k-�KA�W��E-V;荭�J�13|�N���v
-V�w��n�B��1:!
#���z�.ՙ�6.̖)FE:���ŦY�T_$1b�\\�h��ŕ.���30Y�M���y/dA,�w�4�o9��(q���(<�"^:Nl�78��<e���R�|u9�l8�E�][�h��qZ7�M&�)E���ܔsOg'�CQuǐb��uT�s4�'��^WuQ�x��Έ���w�i��N8��A-�dW]5�$9��73�;�WU��a�i��ݢ��,|%�����ˋ9�3E�(���x�αב�WԻ��` V��qV즬U�ѓ`�.�G�Ta�ڸ�\��uL�s+����5���=�Qs\�]Yve��3/I�F����#k0d1b�͗њْ;��y�]1�SwileEp	;.���0�ׅ
O0ֻ�z�4�ynMܧO��6p����p��b5ݤhl���&kUg����&eE��r���HI& �U:�݌��50n�tvnT	 �{ ͑���6�K����$�b�nm�;T�p�U9,_zc6�.�y����m�vT�AeP�LC�*����P��\���G2e֎H!�c6�3H��`�.��b
��6#wc�r��p����Z�H���g�V��޲�$�H�y����'5�����(��#F�+M������/';|�SK7|�:�^Z��	Q��]���G��32�.�g�FtA�o�|��y�Sh�bG�뗐dZ�[=�����o���|��wଙ�����@�m%��QH"T���ܢ���� m���R���uЩn���ۑ丗9է^; �(`7�:�)Q�m�Z.U�f�.цSQeÐ�CH.�{�c�'� ����]JR�qy�g�E�Ubh�|-U
��n���:��
eO�a{W��P�\I5�X�ԷI��vf������O
hcB�eԼL��<3{�a�����S	�fV���9�U�E痫F2n�Ea��jX���j�
`��b^���9eS���E�&�]hC�qm4���>9x�KҜ�kt�p��p���8�uQ]�;;#�86������t<�8�l�9���ֈ�7Y����ha�i_j��s��́ծ�9��S��PU��%r
�����.���բ�NJb̝&�Y%���ŘPܙ��M�E9��x��gj��Ȭ吥"�^�_b���]���W$r:����X��{]�� ��6�XːT�$@��yW\n�Qr�̎�Q���1T���0r�'hݎ.�hʌ�5�O`�97��aӂ�7���1.�.��GL��J��.�G}����Y(·�%�d�û}��;���k��&v$���2�_�xM�ǩ�jv�Z��gq�Q�}�{�X#oxv
-������r�CUP0����ہF�������/6fZ1���e>R��B�I䐋��1,`q/$�o5�.Z�좟c�M���'кt�0�&�u���!�ג���%Y��f�F��eU�].n���1�Χ��[a��QR��vu���Xw�F�Zm�]�m�7u�B���8gkUtЖ��f�l}:��S��kL�NB8�z��ƪN��&%�9��pڷ�l��;zޗ8��R�-�տ��ΐ:�W`7mV �5t�Q��l���;���)��8�����l�g	S1��������sQ�=4���$BŚ��R8���>t�Jwg��0:�hre3[�ݨ��2�@wTۗ֏el�� VU�Fحι��n\�0ܹ���|N�}��wxC����%ly��]h����;�*}���FXl�I�bP�p^�h��h;��>��[˥��HÙsxZa[W]�V_n��y�l��J��!��
wjl���`��qw�S�Ԯ�{�8C�n-���z�;�]��s��`M�_%��]� ;h6�D9έ�7�mvԭx�&��օ�9�ծҝ�,U�rY�Z��h4��(R�wg}���ƙ�5eNde�x�hˉ����(�du���to5��������kw)F�f�8u&ĵ��)g�t��R���,��|�S�p��B�TM�Ed5؞�+�ŋp�I�wİ
(����-z�:Kl��I"B��v�S�;Z/�eNǟcAK�0V�M��+�`�n[�ܭ!+:��i�?b�N��:;��
���6�� �nLoLw�,j�o%6M�.���ف�T���gsr��d��D���Z�	�q�f`Y� Wn�4�'0�����N;�'��L�{�Qw��c��3S9')(�.m����}�T�8��v]\�hwp�5�Ȫ�aܫv�+��j��r	�	�������aƍ�N�zy�d�*�ݶH�Q=���3_r��9�]��=�w�X�1>ց�s\�4������=�0+2ωƦR���6��7�e��r���"�U��Zwuп��n#�.�&�fi�0���KZ\���v�7A�w<���>�P\�"F>��$8��΢�fv�����2އ��Z��(.��47t]"���"�b���dp,n�a�h�oM1��� �VZ��=�Z������ى��*�M�SV���G����{�bSVu=��jj����A;�Ǆ������m������/4m���ڰ�;\n_8�'�L�y�v�9(��%+/�H$�K�A$��;44�CuQ�Sf��C�z�B�$�P�{!ej4�Vm�}����B�(�9��l��a��YȐ�uJ�n^_'�dc���qϨ�*i����j�X�C�C_fcAX�u&�4����a�K1��Zb/mZ�Y7%�
֚o�N��Os��0�Z��ݧ����40ҭ�ږ�L;;��Ȯ]Hk������7;+p��͹ac��uY�e��&HP��'l��)%����n_8��ٻ��;qp�X�VsYN���c9�tUc[���<� ���z�h�vz��;)��:�!����C
�'u��f@���g��kp�;l�WJ���PJ·�P�,!rmy�|����k��Z��vh���BW�2z���b���{���U��)�4��0B��T��Ib�j�"�4	|��3v�W�[/����Yh۰#�ݱ�K��*�K|�%��8lp�.+�oi໲%eF&z�uKu����z����I>�$Q`�-�ekPm�UZ�+D��RҴT�ѥB�"��4�,�������֥�*�ģE�TV��+FV�*A-�-�cj�+V"�QmiZ�+`�ER�Ȣ��U��h,`�F�YE��Uk���-�Tm����%��5iD����T`Բ�KZR�E�TP��FT��k`֢�ұUJ�QX�URҥ�+bUTZ(�U�E��j҃�[eQ��F��-(�m�J���EmZ0Kj(1�*�K[*�����aP��)iH�cEDeJ�X��+J6����(ʖҢ�����m�"��E��[IDX,��(�l*��
��Z-V���V���*(,)lil�Q,-E�V��-Te��Ҵij�A�mm��R�����T+PkE1Vڠ���Ĭ����+-��V�,����R�,���(�X�QUB����ѥm+lU�",[J2�����-kkDkc*-��UUu��]�a�+���5�F�&K}�T"�5^Pj��X�k8����8d�+�@15��d"��|��.OuuS攣W3S��Q��vOpƻ,�f�)��,h��pU��� o%L7���oy��Z#�(J�V^E�p��ꨭ��=�>����۝q��LR�g�ln��ol�	?a�l��%�J��+��60�#^�c�OtX��ʻa��סH�g�卡�:�E#!@�t��N32E��A�/9ԗ�\LX;�d��e�7� �ཞ\�a�.7%�t��W�@l����+,����&Z�lXkMKq]ʺm���:\F��m�V��uz|�R��@`B4T���b*0��B��]�V�'�ʱ"$Ni�V�r�F��PY���W<.�)<bཬ���@Tz\����Bv�5};��rqY���i"�D�~�.��Ld�x_�:�� �b���Z��x]J�eL�T{a���7��Λ��`��X1m;6��T�Wƭ]e����@1��cD)�(��N>�i�)�G�#�ov8p*�98���s�^4t<20B��V!i�Dc^�s�U�	k���`��8	��H{ڪ���Q(g}^#]\K�c�(��w��.ָ2�w�K���
�JFa��jVƻ+�t�o��R����.�x<�7^�Y84غ�����71�Sy��5�:]倧�l��K5o6�릤w��-��ܫ�dil���wm��v�k�ޜt+�J�GF�p�]We��/ܨa����⎛����M!�� �X���Ӵ��[Fb�#�`=6"Y��^��b�č{�nW�ؼQ��t�߀^%Z����I^�����á
�`�-�2�h�W�;C��^��f8A�ddLѺ<�\�y��kJ̄�u��̼7S�aFĉ�sV��v�¯,V���Ln��t�/���nZS�}���q�>�k���2jğ(]������r�^��ϥ	ݳv���of��$�n(�!�s<"����3P�QL�e*�SȈ��1p��!��x=齬T'�5H-�u�du�jV���hrlO��(-s#�"�Tdu�S�O欵[��FgjԢ��8ͤ"��L�xB~G��|�x�6�i�N�p �N���J�Uf�c�(���b�6W9��t�~W:_��!Q�F[�L�>Q8��}���Ur�Զ�q���q���;�2cQ�G%3�y4P<�4$n ��y��]܅���z@m8��tj;�2�rI*5��Ǵ{����m�d���}m��L���r��L݅�ܾ�:�[�ѩ�`�=�;{��;km*��\��m&a������s���6&�G�7)Nn]�G"�}r�:֎�؏F��ܔa����n:�v���+ Xش��B���2�ܮ|'�u�cKjv���=�]�,X�nrd��+����(�K@g�8�
��/L*Q�������Y}����49�SZ�A2,C�|8��w������7��3���~����Mf�Q���ȼi%b�����T
�8<�ЌܚJoL�����}���9�:��%�!*��U�}6�Z��'j�p�E�K"��Kpkym��<����N^��1\E��/n���k�����"h��X}��ѹ����B��/�'4N����vƊ��*GE�\����^�ȭ%��ᑇED�2"B{N��3�3s�N��j�u�q���I�䫲q�+z� h�E��9�
�m�����N��� ����eaz{f���ne��i:���H{s:������oI��ןӀ+��Y�B�A�ZU�iTj��Ql��<���Q�BgY�<��2�-�f1���f�27.�_		�:��}�a��>��UkR{�oo����Z3����1ә��$�Z��KG�u`���T{`i�Ioh��y�aٻF�"�mj'-�7����Rd�Y��Fd���6��p�8��gVũ�<��c�������q�v�rR�$$1J�3���κz��sk�7�ȺV�~�����T�_��X�Q���2�n��1O���ԕ�Y����޷=��Shf���|�J�*�[���(B�>֦�̈'úu�>	��6��jG�[؛G}kYub��y��v��u�j����l`�ܷ
Q�rS�ޛܮK�"�u@�<��ϵmzQ�f��L�]GS��<0:8��|cB��Ju�c���a���� 58<�Eʢ�=L�=�d:#iCk;�O4�v?o�r�w(�"�:�6i���~�1`������w`��,yTI�Bn�,eje7|�7B��j�����i# ~��P���2ܥ���A��Y�Re��&5»�qA�U���C���Z°���ҳ� t�c�+nX���0�W�����nD_�N�-����y�|�r+�G�0\Iд�1A�N1�LH�m*?�x|�7�?�}���w&׷ѽ�{�˙��d���y���c$�I�1��Vj^W�O�:�{r�*�*���5����< qP4\����czolVb��op���y�����VQ�䕘G��uft�6z��G���"-J}����4�b�q�[�5I�(��܁띭����Xjd�,���0�ǫ3�p�y��g����ϕ��'��-�\���5Â��w��S�+��H�/j%��6��tj�F���#`��}GE���LT�����k;+���rbp���V����c���{2\��qU,R�Z��6��:�ш��.�Ľ{�U��7eBV�g�q~F�b/��Awe]�K���*�^;��bb^+��ڦV�4����S���s��\�E�)��m���z���ƪ��w�ڢ7a�F�7�����<A�;t�*�'�o�Br�t�vag�:B�W�>�}�9�!��m{2ޭ�C ��Vn��Wr���^Á߯L����}C�Us����l\a�F�&�UÂ�  `n������x���p=|+BNl��B1��p�����e��>MS�+9Su<�U�{^;	N��g���c{շ>��{ih�=ث	��d�Wt�k�gp��Mnr,�9RK�Wm�o�{�GK�uj84C�����]^���,g��`'P�#���
vk,��w[ah�!�o!*��{�.��7��L77�4!cY�b�\��/k zۑQ,�Rm
�K®��|���
F%h���y
��/O=�%���iJs+�P���$��9�!v����;�yr��a�ϘnC��Ц��`�d��u�^��w�-v�el���Xh�&���cn�����c�zŞvf���e�IO��h�ܕ�Rr;Ǚ�V����|`��D�t�P�/�\�(Ue���n�,�	gǕ`�����q��ገ=qZ���������N�?�#8�'r�"j�&#A��"�����i\�"C��rS��}�AD��;�,?Urw 9�y���Y���;@�7�R������%3A�@�9�h�c�t�[��B�P�H�o*����d��4/K�4:ᑮ�U%���R͇�8�<Ұ��W-��u_�#�D�p*9�A��Ys�'���5߁�p̞9s:�	n�s�+t荎m��Ǧ��V���L����%���£�����^}�dU9���r>2�(�{}gqp���^[ei�F��B���Q�-�頫�<���'Z=P����6�nN�9���(GK�� ŹͿU��AGN+�E��Bc�&]��K!`���� �{c%��*�S�>�ٹS��}�, �����aB�57�O�
�8Ӵ.ϹB��3o���1�O��ΝW^1��G7���h�\v�sK%�x���U���g-���AF��)�g��}��):���w8��|��θh��n�,�Q:�^�D8/�� %H��y�rn�U"�د�i�+:��d�`���x��ӏp�smG��Nܖ���U�d��������vr�l���������uݵ'sj�G�*�>ŕ��g�s�V5Z��uZ��<J"��PV�G�+�"�W�a���BF�ɼ�n��{u�?j�Δ#�f��[(Ch�!q�Q��Ĳ�M���������;�C�(��0
�_u��%�߫<hU1;L]�e�1p�R2(�|�yף-��yF����}{T�;���9�ikj��\8�/��:q���+���`����t�;���G�L�Ƣ�wYw}1yJ1��������Y��=��,�[2�[���u���H��,;O�-�����Gf�e6�-�1�YD�����p�_�)���)<�*"!��/��	o�[�l��,{�jԶ2{1��j&øNkY�dX�~��Í9uadQئ$�y;�:0`{]�h0��MN�j8Ԥ�(���.�9��j{���z��U���r�.�q����u3:�w쪧%;u��j�s��=�EfJ;�\��ym������������2�����Y8b�N-N��0s�%VH�g�+E���Q��ϐ�2$�A	=���L����ȑ#q�1h����`Q+�u��K��<d�sd�$V��ΡN�fq��&񑜴B9l�q��o��yYBM�x����5ū��˶��r��(&iI��7���̄��u�1j}���Q���f3�Y|2�3�J{��-tx\BmZ�{a�77�
sb���]4��O�F;+��PN�+E���;�b7���3g0ޞ���gw1K�pi��2��U�0h!��%c��6����N��@��b���}�����y�w\�"2��c�گl)u�wyW7�=h���*�VD�P�C���	��6�󽽔w��P���R^FQ�p�g<�TD�I�rpd��J���f��8��]5HEV���}�42s�K��X8gK���nc�Op�)u~n��A�˒��Ä���FeC�T�u^8��*9�;��6v��H�[�k�Sτ��OϽ�b��nP�5�/{���ST�Y�j�F׼UR��N��.Ϻ�8)|Nq��F4hMC���i�l9�8'�W��#��=:0B��P Kr�po�����6>�ڨ�x�G�qw�)	c��61�V�q#Sڄ8MR��m�i�l��3�yk�2�
��E�����Z��Ή�z�7���⧺T����Wh�b_!����b����)��DtYcʢN�|u�����x/j�c������%�}�r�l�(E�"��<��o�=��AEC���{�*�V���iu���q�:��/����.�giQ��)g-�VzQ��h\��m���J��ɴ%��������;�w*dԣ����%6�@���,0b5خ���+���\�^���ͽ�qQ!%\X5�aBc���.���)�T�R��^�S�����R{����b����dw���P;Nk���@,�ڹ3~j�xK�ͼk]�Ov���1�a��/NU��:���Z$Vܱ~��f�LT7j�F]ePaj=�d�y@�>���� 5걕�Z �pv)��W%�C�65�]b�����G�,�v+�
Q�xnո	wgvM�ƭ5��d�Ѧ��b�iWC^���W^�1i���*��w}�)o��fǙ�(g��i��5X��9� �NҾ4Ѱ���8C�r��j���WN�$��Dt����^������Ń'|�h��'�s;�Gg�1��С\��x�;+[QY��u�	�L��Q���l*w5������!���D� nxvTdq7����;�+�E5�D�C�jt��Esh�5��z������i.O��WV(=��ǲ�Z�)8F��U#7�	�n�t�u�C��N���\T|h}��������ܱXއV\kJ�׳�RUH�vŊ��>�\�:����%�5�3(�[��3Ż�9]��A���"�a-�V��j
�//pҝuŽB�h�n� �٢�txo_�F�t!�'{�&�D�o�h�gK΁v���ձy����X|�G�&��έ�Z{���b���	�|�h쏝`!�
��PW�V���5����7�Se�fj{-�QͲ���3
����������̎�Ud�Pۢ=^��8vϚb{�k&?+��#��m𽓳ms�
�(��Q���ѿa�
��+��,�ӘX��
��!\30�e�����b��6��%b�����JR��ًW<.�)<b������@R��s�rb����������4g���P������2���Lp�uc���y)��0�X=jz���rf���S)t�T*��U�O���"3Ɠ�;��&��Z��bʑ���(���ۜsNέ�׊Ip�pp3R^�S@��j)z|w�t�7S6!fD�bd��-�gtM��\j�ԭ]��l��0H�΢ED75d��	mƺ��%%��,{�n�V�v,Lb�;k$�)��^��C�D��(���t��j�x�h����+�6�F���ҧxu�G4B��o*�G�Za����pT�#�%����½����7�$<�"z�@�{\u�u�9�����MS�%�zt[Abt��ok"���wl�#Y��D6�$o�B�X%n9��]X)�r�p�C�ڇ�*	���hg52���mp����p��2osK�r�I�X�����3�2KG�N�ƭ����pbzI"�1=�Q�`�1�V���;F�u��Q�z
ζ����J�S�^_�Nb��0H�_[Wz��������%���'H�d�L��U9��ʐ���ۍ�,&�SA�gZ��)�J��#
�Az�x�<˻.��qL:�����{q�pn� �uJ��Pyٖ�\�l%����@�}��y�yI�9�T���b��kZ��Dw��1�-��0���i�ic�,�����%l�ż��Cɖz���j��Hln}]U�^��/[<x�	E���z{8dzɒ�d%a�g�Q W,V�K%��B���^>xtޭ�v�OcW�I8A�ޛX�K�K���]a���Z��E*7/� �ח2�o$xd��4iS7:Dɴ���X@�@��bȜx���]�&T�u4l��`�C�4��
�`*�>ti����j\��&y���.�C���0�㒹=㵩;&�]ƈ�2r�N��5سՀ�	�L��9��^f�繎�w�'	�h'����cT;Ļ��6�S�7�4����b���4��4��v��pn�z���1vU�al���7�3f7�{�f��� "E�cVB��ta�T�T/��kԭ�"R0��-�w�YNȎ��t�ݧԯ/bsh��*��݇z�D��(>r���g'�?��x�� 1|�"�Q�y�ʄ���$d�/��٨w�'
Ė1fv,�Z8�&,�bf�u��Zl^sc��7+M^'͹�p�=a�b0M�Z3kWJ=��n�b�n�<�fU���v+\}��fN3�Z�j�G��K/��{e�h%�
��ނ��h��5d�k)<O��tKa�dh6�@�\�>z��5�zVǫr�'34l���'70�f�eJ64&�2p��n�"j7:@��X�b��Cm<Vp������k%t'�6��H@�yv
\Yun�RF�x�r/w>�6�Dc����H\7�7-<N'�^�
nv
Q�!e1z��4�p}����"{U��i��I��Z��\�F��a�HnZ�vU{�H���ք&�BJ��Q��z��G��e«��8s�r�3!�w���C�z�^�Z�ѓP\e<2�5j�iV��ʞh�M��h�*U�%�0��)�N�g�*��,U��n�?�ZG5�+h�ʑ�E�Y0Z�W6�1HY�fo�f��q
�}�C�}����JѶ4�E�
�Z(�#��
)+Z��m���V��F�*�m���J�-Z �[U�J�mV���±k*�PZ���0R�B�b��IKE�#Z�@��m����DF�RѶ�QJ�X����"�hV1�FR��aZ%�(��YZ�P[F؋k-aPH�BڲR�)bʵ�h(�V��Q�h�D�DQR��(ȥKR�[XU-�*V�m�F��-�T[T�%U���-m-b���"�k"�UeDcR�Ee@�`�+cK(�R���R,�ZUJ֫+m�Ѭ�KJ%�J�-+R)Z60YEe�+lJ�Ae�m����F*������*"k*���[de�m���Z[jTP���V�������-��[B��QV4B��m������h�Z��mlA���V-�m�j(���V�b�6U�EUm��YE��(�R֩R��Z�kB����-+
�j(����e�AH�**�m���Z����Jے���{X7��(0T���ө\������+�4�ớ��}�c}�����6Z�i�@��#��{
���[������d���>ǞC�E�vCmKGr:h*��`��Bu��\S��c��W{��6�ϴ�
1���p�W��E/Y�TR�i!�ߝp����L7��^	�=��rq��.�~��SJ�I����l��W���E�1'��WuA�>��nN�t��s��J8��r�6��>�֥hds�t�i�G)Up(�����m
�m��ꎟ���6ɤ�<�B�i(K���#~�S��]<�s�W��\V��M��Q�2��3>��:�Jbq�VsVfJ૚K6 �4̍��J��ث�W���7(C�z��j��bWFO76����x�K�u=�R�
�xW
�)�zUcU,|&{�u^�%q�⽿u�(7�H��ҨA�"��fa�C�<�'N#0=�c*!��tQ�L�t�:(p��D�m;�����=�k��������nk�:�^t���z���k�}h
w��`�q�wq���G+�$���G<�h1pz}�_��`�]G�������,�ԅ�w�7��	�eE[2YM������T3�f&�<�iϔ<M􆛻��Z��9+°ƍ5w�'��)W�'�y�t��}�[�M��t�.���|��^���o��4u1բ�C��QRcr	��5�ѽ�\��ճ/+�ު�55Ĕ6ݜn���crqy٩��1���v�T���A��9�c<L���O��&;�~
%��P���R�`�.S�i�Z7�.]����C8e�BU�1U3��N�&Qy�j�|�Ռ��y�y|}���溒�}�K���sb6t^ �F�*�T�ޡ��3@О��=G4bG|����j��$��1���<}�2��a�ep�q�*5ϐ��M^Iނ#J�O9,0�3����G5=��y2#�f�o<�/����]fS4ǽ>����y�?M�]1:�=S����~�ȇ$��Ysb�ԕ���V�ND�^S8�6��izӦ���/��4ɮ��=5�Ծƒ�������uc��i_������)�����t'�-�ҡN�v�k���h��-9<�܊um�����5M������Sl��7/�_����Q����7�N�\�����y�Y��b�;4�L���)���<#G
ү�]G[u��yNI�
./L͜Z���+���3C8�6+��}���	n��r�N7,1~G�p���uAY���.�*c6=PՒ&�l�>�tƸrqWzĒ���Χin^�ޯ:�Ā"f���3���н|UlëhP�1��*��{��$�mn19�,�P�'�Fd�[u,�/�:�;�b�F�eؔ�ɨ�\���;{}�d f�U����R�Zk��)����9���6����EՈ�'Q�k�Bƍ	�zvH�9�z��Z�,���SN���
�^�f���+�(�6qdLS$!�w���Հ1.���֮������u������l\<��4x��4,�3��"�âv��n�dHW�t��y���~�څ`³�
y��2�w7R���a�-����w�E��m�KԳ���<3�΍�(�@�6# 6}�
s�j&ô�A��Y�3@s<֦׽�����ח�ÞҌ=&+��:)`�S0{؀ͻ�H<k�6��{��؜���R/HC��u�f)��%;�f+��b��$�zn�XY~���=�O�	Pb�6X�����i)z���z+�#{2�oT�Զ�	�`�V|p�R�t*���V�bw����w���R�ƭ
����h����sܡ��4����\��$`��L�0F	N@�v���֚B��Ϧ8�_#Ok`�3̫U�eH=��y�eW���5d���K�C)�6��*aH�0.�tʑ�uq]�T���(�cX=�����u�I��k�&�U�O�,��
h^��n��@�6AGC�:v�+�찱�� ݛ���P��qe�Z�J A��Ɵ;6��}^a����ZջUZuH���[?P<�L�)Y7����E��l	���ĐѨ�L���(�Jb�!S�ѭ�`�=�cu�0A�+E�~��so�T�(%�9v�:P���Ӕ8!!77�q����P��<�����j��݂��h���o�^Fo���
��]vx�4�!�{���a�߹�%���*/>��\���V�����U���lX�*+�M@J�:���)�cr0ՅST3�*�`�!(s�ģ�����͂9�
{�PW�z+YȣXP���g���:!%�3��Z���#�a
Á����J'O^*�@�m��=^��(��0b��O�{�9�)Yo6��ؖN�!Y�W��_����]sō2�*�N�/����v���=�m��!Y���J�Py�t��肝e�x��Gz�%=U(�j�n
i�z��]���]^8'L���dZ��3b,j��3
g��u����%<!ȧ�N�Re����}̌܋�9��\�g�lI�MMe�56Ɉ�j�F2���Z�S��Y�|�B3�ܒm�w�e޵1=Z����ٻݷ��X�`ĨU�qN�wV��1>h:a�m�ӧ�����`�3x������Y@�C�
��+�i7�}�}$��X�1v'�ʙ�Fc��U�]ָ!Uokc�:qT�]����'J6�jgi��"yJ\Ur\# �^�j)s��PgK�$Ѕy8ӆ[@C�~#�X����Gޥ�X��o�� H�΢Cf,��8Z���.:b�gE������.�ǜ�@����q2*�z͆�l�>z�,5�7OCF�y�.�-�:�*=(�67a?��L8s�gx��4؜���T�KpR8"Y��'^���oH��f8ux�;�ZĔԑ��5�r����ٴFvC�h��MQrыY���h�Y�63/asU��ǜm]n��188/9Ϳ_���~��
/%q"�������E넵v^��z���y�������Z�Yu]{�A�<~�����a]����I�=Y.D$�NY5ڹrA{��O�������T=J��:}lv�GI�S��h�\v�s��Q�l.��/^���n?J� P}~/{���¶�t�|~���{��l;�%�J#}�PUj�,dL�u�+�Y��wc�Y�
�0x�i�|i:��T�U����r�;�z��ƨ��⏑�=�5m�f��{���run�(Q�m=k0��9�v��/混	T/�k�Ox$�YͶ[��[[oe��!	2v�fv���<D$6NU���1ؕ�M+��`�pQ�f�����輼��̽���F�e����b3=|*.��6��7�_}_v$)�%G�=y��U+"c��ϰΈb�Ţ� ���B���gO�Wx��+7�+*���L6�
�>P��`�ӈ�Tb�ey����r�q�o@n�C�.�ͥ�ml�a;�\'9�:�_����=a�}�w�>dC\���?��ES��s8��X�ƃf��ˆ�eQ����	Cu`��4�
�󸛚��E��n*̩�+���3Z3�]�#?]eH����1p"Cg�38�&E����]}��_���U��9޸����|�#ƮX��b������42���j�}ڜfWr��q����V�?8���^b��fzf}���q�@j������ώlb���q�*�P�i�N�b�I�H�g�u�\��f�&�P5��:~f�C>j߇��]�m�<���ɨ�z	� W_6��wjQ�Z�R�4�vFD��K������:-Z�3�i���u��o�l7��I���<2�F�)�W�4hOg����1����3�[9^���WM��!�7V3+_-���#�Kn|��M�����QW�_;u�]D,�]ԪR7L�b�Ɏ�>���-�a��b�2��j��P3Ш�{t����|��p�J�;����B��۶7�n�.�|jJy�fu��l��t#�I�Q f��y�b��gX�����vi&���� �<'�\�Ǧ�~E���S���p:q���Q�.�?���������\�Z�
��Zu��2�#�T�6ܰ�:uZc�����7:��*����q���վJ��d�צty��� ��U�nc"���=�99�G�9�� �[�6�{)�˧ʒRj�ژ�.�M�!mO�b�!w;�r�N7,00©���#��N�S�:��B08�¼�7x���Lz���vS�6˿.���D���E*;�6��W���S4(rqLw�mS�F�S��`�<y��=Z"�ɳ�"b��tn`^��U)�k5�F����cC˅Q���{|�����p>¶��l0�}ƽA'z8�u�+֧0E����<������J����$��޲Ǖe5�^�$z˜/^w�v1־���ܑ�d���\@2��Q6�9�Pb�a\>6"n{KKe4�ʓ�㧪�JX�i��8'��{~���Y�:��߽�?�w)WW���>l@�:�h�!�ٲx�@�j�w�vLdS�l-%�j��{�\�a��1)�Z�ft�-�S��{Y�/3��8u^Q�:L��Uӻtq �WH&U���u�&�v>�F{4]K�>�DF�1���A�s�3u��b�Qڱ�p���Z �0ҚwI�+��"r������=�Gj����ڞ�78<�'�b���cĝMы�+��|hJ ]�к6q��n�'�n ��ܢ�o-����'��"p���:�E
�]��V�`�x������t���iGUp{S�:��+��W�=�Of��eה�O%�e,TuI_�p�c2)�[�KyqǢ�w�GX�R�&��!긍=��j��U�����)"������у\Or^��#c��X�7��A"�8�ʇ�d�F�e�QВ��.�o��&Q5b���ɗfɻt�,[������*a0jΌ���j���^��PC��*��l�Tɬ�q)���.zJ_;��]{���u��o��x]&��J���O�����.티�GR� �XSӞy�g7�?O�@]p�����7 �q����Z��S��^�_*%P�Ξ�~�,���w7��h����{�ttg��
xp\�f�v7V�c�(J	���Th�:�)YN�e�z%�g�?7��P&�)�uC�Bn��g���8{كۢ=\x p�<����T�6�/z:+���u��2�#�cva�:]t�����뀣(ɬ����08���AnbD�rcfv�����{���]\%�nȇ,�� ���mTN��z=詽g)�7�q�o��7�6���n�f�腆�_S����,o����lH}���ئ�&���{�ڴ9�p�cp�qPo
�ٰ�'��X<(Fn�fQ�[t�1���A�˙0������@��"�+(�q�q�1=CV�ld�Jg���w�C	�gmr�&d�꥗�z��ǔ�Nvj�*Q�\�g�1�����@ɠ���h5G��7�}��%�$h�{�;�X��Ր�\3����C�
hy�j)s��Ct�׾�^��z�F27������ �g�%�Zh8�$O�:�����M�����7�Q�%��	WX���1;���4A�X��bu;���u��(ů�#:/��Tx���S2�Pe2'����k�'L�L�8'M60���f,7iB%���u�Q���qlL-�e�����JÒbC��!zqc�h���x�-h�vk�[�gZs6�7��]�4V��E$�=ƷV;f�
�����p�y^O�I�鰢�%q"��	�aB�[��]Y~'�UvŢ�Ƙ�b;{x�K31��U3Moh��d�ǗKSgN��g ;mWru��0�������*�+�_TÍ�X%׼�u�}����sɕ���k������T�lۘv�с�;��P���=�G�sΗWIkEE#�F͍�x�5�Ю�M�6���)
�Cj���2u���c�ݥA�%��;���oGO�~z����4{`��f�+��p�C�B�|�В1T��� �ꃸǝ��-T���τ�Z�F�m�B�%hVs�N5K��8�y��C���'CF��1��z�ϰ;1"�sSC����Z�"��g�!�҇F5['�ut�]E��������Hȏ���#�(�#���\2���ҍ1����l��.3��W:T(z�̩�w�.�q�O/Pq��hdk�0*��ED3<��t�7�1CQ��ҙ�AqO�f���J�b�-������zyTp�� C�u�
���
2z|2!���pVU�0'�[b���<�n�,Mtw_�ਫ�<\BV�3�FC�_�,sC	`�#]D�ʱ��e��,�.�'������q'ܡ�N��
���|���jM�i�4�yd��@Ĭ�u�?�`���ezϹ�h�~C�1��cY�u'��iE���S}��=��C�3��y+b�~�ie�ϿR���[ɴ�'~�HzoZ�񒾲_iY�%g�����/Sh�5�5�'Y���Xj� ��g��(�q���fٴ1���3O��ޑ<Ǣ@�{ԯJ��Nk��ٜ�ײY3Kс]�̏��ǹ<��"��(�uk�Cs"#:�u����%ei�{`�$��`�Ʃ�M|E���j�'���2,�e�u�T�d����̖X�g6��^d噙�"b�hl���,@���9�"����ͧ���{��|�ڝ!��D^��Q������]��x�Xy���mp�-tN��1\�$��^]G�焊�q� 9{�-���9R󻺇J����/E�&���|�Ɲ]4� ���J{.�Tv��*lI��W#���d���DQ�1���R5-�fir8�uL�ُ#�بjڻ[�Y�э�i�����r��L��)�ܼ4w�t4�|p�}v���\v+ԗ�0���hªкHg<�5�;��uh@��2�u+��g>�F�q��y5�=ݢ�����O.GA��|��^{�i�	�GCe9��E�G��R�<�6k�/��\T�,� ��X��kH�y��ѝOhPAm僽(+��FVI����^��6.�^�4D����,�p�]�I�jA
盠��ٗ�l��U2���bY��Pۋeٗ��]�[�OE�ֈ[\p��T0���=�=�����Z�Ǟ8��V�f�^��>൫{����,�3��}��g�(E�5nn�#[d2Mv"���V�P|�uou�I�s���Z﹔k�L��|X���7��2e 7d�۠�!�����74��u�ޅ63�e���X�ZT�57�qu�fs���T�C�%���!BeGe�| ��id��;�73)io\�j���s�bvŽ3��&;+{����4lk��)�,��g��=�U{�j�Nf<��ۧs/+��Ժ*1���A4S{y���7�j>�e@��9j�rv����Wv
<][b6�.�T�8�A��R|J
��a�(L8���0�����d�w�ʰ�o۽ܼ��A�]�<���nѽ|�&�W�48�`�fg�l���[�S�Go��OIR�
F��Y
�	�]㧂��zJ@�(Ǆ$#����M�",7�)͜�����aL�7��u�i��f�v��e4���PB��`��3Q�ᴰ�5_oݧ�A��mfs�����-d���"����QO0��:�{���QSN��VJ����{���h"���K]��t��"h�ayϕz/Y��F)R���۞�O+�'6�9W�p$3�S��Av����bo{(<�Y˫.I���,�j�KM ����(&Tns���Фç�2�f>����[�ut��t����Nγm���2J���]���tG�^����36�EM�L��H{C�Z{�{	9'L���D����0���}yw�@�P ��'�Z�p��-�]�B���v��v9���n\�\�0�:ЛQ	�wL�+�.h	���WWNޢ�����X���p��D�]����&4�1�ON���s�{t�t�Y\4��
Ngh�������i[b빫 �>��s	��
�;玘p���i �����}s�`�N�A@$�A>��EU2�F�lD�b��Dm����ʋD����T�m�V�l�R��EA�Ȱ��Z4���[b6�A����P�Z��
�
�J��-���[V�QQ[J%e���m�T�����Z��m���l�-(����m���X���ej�Š��h��k@�k
�e���m���T��Ң5��"��֊0�KJ��*Q�T�J*�VEb���[U�*��b��Z4�Q��*�Rؖ�Jԕ���T�AUb���,����[Z�l�(ҕh�TE-)+J�m�F����U���UV�[T�*�KhZQZت�Vڅe�ն��kQ+Kil
�%kF�K�������PZ��+KV���c���lV[`��k����-�Kl���R���+j((�JʣF��6V-e�Ub�4B�J�b�������QZ
�*�cF����֣TF)E�D�IKmB��%�m�	mJ�Z�*����J�������h\�.�ס>O������ӗ`C��ǧ�\����g'I+e��tq������)9o<��R�ט��诽�l��ط��Hu_���$G�I�?�-& (����s&���&$����C����vx�H|Î}a�����%g�7��c&��
bԂ�h7�I��:��O?s'��1����y�Z�m�f}��~g<ozcYQH/{�6��񆝡�w�����/_�0�d�7��3?Y1E7�=CL�LCɺz��ur�'�y�l>aXx�uL@��������*�Ĭ�r�NFU���>���~�#�"c���6���1���ԟ'ω���Ij);�f�c�5��N��)�����`|�7�&����$�t�P6��N��i>B�x����ƾMf��-���yt�J3舑b!�D����q����٤u�G<��|�2T�!S���?3o�y��u'�� ~�aY����|��ag���}���m���ɔXu=f�Ξ�t��e37ۓ�����i>b ��ޑ ��G�a�6�3���.��ɉ�~C÷l�S�����@Qa�5�Co��&$��~�M���9�C����
�#��p�D���yx�X��ë�o�R��~��<�~��������8�QClZ�^��
�gP\f���㴂�f��Sl8ʋ�3L8����1�3�O�:�C��Z�
��Y?w}��7���ۉ=B��l��Þ|~���o����R~�{M�IW�"4G�D)(D|�}=�a�xfa�Ĩ�d޵���d�Vl��I6�z����W�
���k�N�]$�a�'5d�Qg+4��s�����=^��Ͽo��_�j�Me��z�#��B���F���C�9�"�R���x~̛I�+'��s4�b��!����I]3�J3��E��zn�ݜd�<C�)�30+7<��4�d�뤜�s��w���rss&�bƯVu >����d�9~�R?2Wp���*m��g��tO=���4��Y�I-�AOfiE ���|���qCٺLv��1:�'��mĩfa��L@QNm޾��_3��~��l?:M�c�
�W��w��G�8¡�9�y�gY+7�{�s(�~g����(V-@��᧬
�Π��~�C�:��Y���0?&�|ʊO&�c4����|�`)��tn���3se��[ 6dt�@�2T!�e���9�"�f����*�7���aܬ��k��&�Π�5]��c'��D}&^V�sKs�j���:�b���7�n�n9j2���;0�ռD��.��.���D�D+�US߽�G��o>Ч��s蟰G���1?����`q�V|�g9d�OO�"��+9�Û0���:�t�`a��a���봨�a��X,=eU@�]��{�d�&!]'X~M=`���P��M�3�3s9(H�������f錬������+4���T�(m �$��a��1�����gS��~�H�x���Ϲ��I:�d�g�4��%}C�=�|�=#�0=���_9�G��]��4��"!E��MfC���%I��;�O�>q�����N��Y1���0׾{��R1&�zé��퍁���u�C��\Hn��?�6��ȋ�xC=
iȚ:���.���Y���3�N�b���}��6��k�j)^2b�320���Lg���!�J�=?Xm�aP���}HVi��&�wTR=*(px#�2o��_	9ۇ�x���Bx*q�C��Z�'ɴĂ��0���6¢���,�&0���1 �I�=�f�^���O5��Y߬��ɻ1�!Y�hz�$�
��|}�������=�4\�TK��:~�o�V�т#n��Vi�<���QVM�tm��Rb�?wR|�n��x�x�Y4�t���L��2��+乕 �I=q6wX�H>��5��Ï�c֊��(��*����1uҴ^��˼�߻��E�S���$�
���1��J���)��β]��5=d�
,����ͲT�w�tO�4�O;��<a�
�d��;`c?2W�7��}�Dz ��}M���ͮ���{�ç2��~���l6�����Xv�a�Y>jC-���ٌ��&��c8�
���/����by��=a��a���4�2b���XWL���Q�"$G��ba֯���2n�V[w%�q���;�=w�B��=�4Ͱ��2��i:Ũz$��
�g�fI�q��f�u1�QO��3L8��w���A|I���S�G�z�G�(�OĆ"�rD��ŭ���L�欘�����)*��?_����I���i��~a_P�;J�Y�~�4ì�����i�2T�͞]=d�c�|�4���ש�<9OH�{�>��{گr�Ȭ�{Y�u���R��mv�&J��Mp]��Ǜ���/���T�s���{�3
�M��$���:�.��X3���׉0���c�fp���wDi��A��dt���ׄT�M�(2��vs��[�-6�ʞW}�%�n��6Qj�=3��{� 
ߒwl�{������?$���O�PĂ��ݓJʞ������1+>OSӹ�ii�f�<O�1'��T6�>�a�y��06�u�����%H.Ӄ��������殩�������K|�ϐ�m��RvZ�l*|���f�?2W��I�m �׽�~a��Y9�c��rÞ��]�:Ԇ�9�oU�H,60��+8�;�H.�DO��N�{%�}𝭯�R]���D{և��!4n��'���w��̟�RO��j��|��,�d�����O�Y�� ~d?&�f|���8�߮��G-�j�ڋI$���h�X����� �L>LOǈi �C��8͢�0��_�2|��v��7�����;jM��'���c����<=�a��T
��p�&�c
���s����|�q�U�D1{�Dz~�1��1��a�/�N']$i��C�Y��H,�=���s�1!繟 Ua��19�'�HJͧ�w�ڇ�UT���uhc�
�r�E�ḋ�{^o�O���k��{�4�:b�N3�� i+=gC�`hg*�s�2{�q���1<d�ǌ���L<aS�nj�x��Y�'�����Ă�����oXu1=���������n��M��<ߙ����l�!��s{����w�LeT��O���CRq5i����cM}�I��Lg�Ȱ��g��06��z�c��`c�+�$�G��Ǡ�p���`�]}�?-�Y��=zN39�N�ϲi��*(q���$�
��d��M3�0�g2f�bc'y�4�YXb}5a��1 �M����<Ax°�j��2x��t�$@�=� ��M��o���ݙ��_�~7��N$���Y�?>�c���0�q+&��9����XW��C�+:�P�w���&����ɦar��;뙴�Ͳs)�wY��Ab)5U�
���>�Mɟ��{�Ѽ�s����Ͻ��=����!���Z��Vn��0�Aa�i18��z�SL�ez�%v�4�01����ԛ�J�}���LgRx���!S>q��u�i��T���7����������a@~Uu ������ŹS�q!�H�B�^���f�^�Oju��E)F	X2��48!�iT�hr�I8�+����>S�c�QA2g��j��й6���0���]���N��YV
���qGJ�b2��2�D]��_�tU��z�]�;s����z"=��֓ׯߋ��o��P�Ǭ��T��fO+����S��>�.�6y�:�5�M�8�ʀ���a�b�f�߹��$y5�|�T��a�CɊ�4P��=�g�7�jK��~Mb_��q8ϗ)1'�T>N�04��z�����������&��
��<=��z�QC���:H/���:Π�����{h4é�5�}^� G���}3O����>��4������!����I�1�
͟��|�Y��y����O�a��L�l���+���=}@�<�c���M�P�|�Xu���ÈVx�Dlq��C��18z��51Ԫ���t��ݽ�ino-���==�{�U�	���������QH)���^$�ğn�0��?�*���妘5�_��=O�x�����i�OXbO���'����ǈ~a�k�w����}�\��Mn����~��>d�~9CgY?e�!��M$�
�d�ͼ`V0���tg�|���Co̗)Y6�M3�%q�ɉ�p���wf��x����a���PYP.���W���{����߾������H,���z�!���q���q�a�>?Y㤂��$yt��ì+�߹���$�N�&�������J��c�L����J�aSV��c?2TY�~_u>��|��o�ߵ�����Z�]���|�\g�OO7�m���8�"�YSG�q6���1�Wi:�Ax¿��I�6�������w'�
)<>��Ϭ����w��N�^�@�^��>q��ӝ�6�5D`�H�H�@I��2�=�u���v�EY<J�2}0��񓉜���0���~���z��欜j)̛I�9���ɜ�*�������o���~�{��w�o���ܿ�y�t��M�����&���C����d�W�S����ơ���n3�J3��1%E�d�YƤRi
�0�����Xm���PC�
�3J�=��Iϐ��ݛ��}��������%x�i�߼Ф��y�p���0:�r~�y�>AeI�9��H,����L�Ρ�������a�y�Ă��f�hmE�P�U�8ɉ>B��9�u��������ʵ���F����*�g𗅅���K5=ܯ0e;*�ڙa���ע)e�]Cq]�=J�2΁�;�u��͉��M�=o�1���D��=�o]o�U�!�sZ�g�����ԨT4.r [���n�&�V"r�;;8�7=�G��O�����p�!\}"#�����������%g�J�T޹���̕<;�h=VT����6��\gy�g]�c&y�j��R/_�
i��Pğ!]�����Dn6E��3q=���;[w;���A{�2����d����
�ydğ>�I�+��O9��V����gY+�w���VLJ�!��&�x�8���/X��_�ro0?=O�o�KF�:�sd?�v;�3��V~�n<j(��&�C��|`V�Ug|��MI��:�gS�����ҳ����d�+�l�u�m�a���ͲQ�I�y�@Qed�����ז�������I�8Λ�;�!Xi<5��O̝��!���O+�%����Vx�^���g��M�[��u�`m��Xj� ��g��(�q���v�hc4=׺�����{�N�����6�&��zf`jAN��/�h�@Qa��c�u�xσ[͡�
��������������L����=����d�(��eH.'��&����5�q��{϶�#��~�W_j�z����8G�H�}��+�QH.��p����C��0�}I����0�d�7��3?Y1E6eP�9���=CI:�z���ٶ��<C��bg��G�"-�Б�h��}�ZzǬ@ {��N�a��B��l�;���a�/�9���?>�{/�5'��i���}��<I�!�6��H/�]��h1�1��P�&3��I��@�Q�#��je�u�󺯓Ɛ��{DA�e~zr��O�>a�y�M3��g�x~�H
,�&��|�����
���ԟ>?��wa��O_� v��g�J�%�|ֈi��W��s'��R���>��bC�j����c�}E�P���4���򤯇�LE ����!��?!������g�<��Ƥ��?k�� (��w!����z�~�M��%�����P�
�0���?k���?Z�fErX{�J�����x�1{�}B�|���<bԂ��������3��1�=��u����La���g2�u��{���Ʋw\ɧ��& /�w���߯�3�_��z���J׎q��]��U���bEQBƪ���L=����5F��#f�}Ɵu�+�[�s���1�\�*%*�&]eF��Աś�!�����2�u�����q�޻���w�K3��4�k{X��|��I��{9�NSv��B�&c쬬p���)3��+�ٴ���V�q�u�%6�k�}_}U����Cԣ����������O��vLO�(q$�
�~g-��q�a���8��������������i&ЯP�2�%x��1�&r��뤂�/�<d欜h�<ǼG�G�H�>�=����O�@���_>?wzXq��08׻�x�fvɈs(b(+<O���d�N!Y<Nۏ�)+�a��ݓn��
�8�ky�(����Y�J�ho
q�BC�#۹;Y��wA��=�;%_���<d�ˤ��04βW�����EH,��]����M��_���o�����s�ju�!��+9t���S9�1Cl�C�t�퇨bu�K� ��<K�8~́�dWg�kJ?k�L�E;�����8Ɍ�*$�{d�{��Xq�C�<s��βV{|�T�i�3����(V-@�{���*c:����d?3����h~Cѣ�@���#�qdܧ�rT�?3�&0����v�|�~f'��<aXj��c��&2n~��O���Nh���I�+��o�h~aXy���|����=>�YQVN%�y��������<�@,�!qF����~����Xc����d�8�IYY7�O������m'�!�T�hm �$R�;C|�@�Vu=a����M"��Vbo>�w$���� DA"�&+'������f�ԥ������k�4�c
�;?gڒ�(��l�d>ݜd�4��4�2z���,1=d�.���Led��4�^Ҥz�v��LE �x��'Y�9�Ć�CW��4�����y��_|��E��ܬ�+1�!����i���3ù�Cl��"�<d�.}�B��ӌ��hT<a����0�*!��^��d���x�ۯ�W�w�󏁩_��]�Oɋ��`N�3�I_^�H��#�NXh�
!�4<�u�|�LH/{�<a�x�l���YXm1��^K�4�]������ԩ�!�+;��y�1�!Y�hx{f�z�I�?g���o�;�y���{�y�0+0���m;J�Y�l���q�d���i��Rb���q��HT;۶�ɤۤ�;�3�L�'�\ʐY����������<��Ұ�����5�{����Z�?j�h黫\���{n*ko1�M����y�"�5]��]NNA�5�S���+w^���V*�9kVJ�Ro���֓TIk��8{��!��w���I0��_ox{k{s��폟�@�+6�a�PP4�3w��I�
���1�W�m�M04�u���sS�J��͜��I��m���w�tO�i��ü���0��K�C>>���=���w8G�_T���k��{��΅�*Ag��1�S`t5q��wa�u�Oe�|Ԇ�}ef (�x{f3�P���P�T���1>���n~a����'��& l����c�D���M��Ə��d����%?G����q�w��a�
���̞�������T�6§��\OY18Ũ{<�"����q�2�I�q����La�TS�����&0x刊��z�n{�2�])c��%^�٤�+��k$���jɌ�s�CH��Vg��s���O�T��r�}~@��W�P�;J�Y�~�4ì��6S��|�Rc7<�z�c�T1�哯SHl�=�o�������~�'�~d�Y;>��[E �Ğs}�I��1 �<d�a������q�%g��{�M�(�m6s5��~a�8�f!�c����d6��Y����{�D@�ț;�a��6����̞{g������d��i<-a�:��#��x�Y����r&�H,���a�LE�g5�O��S��w3�Z�����oU�@QO@��"�cb�t�O(��SԆ���y�>;*A}a�j�3�`m��LN=d�2�ì+�q���6���+�\�V��{�_?��tyi����^�3:�Ү]���'s��>e�����z�CY�����f��S<�_�pɋ{������`&N�6H6z� 5���:���(h5�3�^zj��� R3���TfRf��Xn!_Sn�����io:�u�X�Q[�+��F�*&?E��"n�
Vk!�g�(<�{�l�v�Z�����쾺b���]�Y.XD$�Q鸩�нnCS={�1�;�ƫ|�D�u\��\{3&�=iޖ���ҽܷ��o/t9��B��M�ʒ��uk��y+.þ��F�v.����{�Km�W��ZU�O#B��'Y���Ɨa��{��w�մ��v_J��{��{���V�Ȫ�����PVW@��"��^�Y�C�hj��#+�3� s:U9"3M�*���d	���3�,�4J�3>�%����B�ɰ���0�u�	�u�%�g4����ʑ]��{= �"�� �TB�Z�3V\# ���<|�.<�V�KXK_C�3C�6"��`�^�}Q%���a��@����x�'�Ńgҧ̺0���Zsv���SClU=X�0Ǹ����	A&41ܲ��J�#yg2���y=�~$e�S�:�t�f�tmJ��z�`���ح�_���Xf.�%�+��]7QK.�2U�*��\���(f�Ċ��DO[5�d��q��xo�;V��LY�80ӊ��Xt8c&��xқ�G���q{�IU�����ʯ5Z(�\�!No/��3/�M��w:�!{; ���f��o(W���!	���aZT���ʣUN6�MǙ�
�F��q��5K/�j��K�f�>�i����^b��hg�:h����� 8m�b#L�_%�I�[�P� \je��]،�	��x��ƽ��zj���:]��:K����>��f:'�u�Cc�C��ή��*n���Zlew*�>�ح��$��Uފ�G_AF[pA�T�:�fe�Q<��*�qll�z�+w�z=聲�w;V�*Q�>��d�Ak}u�b�S��Gf��� �yj�Em�;�ӗT�έ���T���r\	�Y�XWϰ+�-w4:���R�w���et[^�7�b4\��:y�[A�_Q���tQe�:	��;@B-�F(t�Rq�ڟ˭�a�w+X��x���J��`~�V��
ָ�1�s�*"��EC3��������Nz�ĥ�⯹�4898͎���6S��ٸ�a��0������¡��f���C¸���.ޔ�P��lh�s�)��íJ��dƗ������1A%�ۇUѝ��!'��nu��K��X����eY���^��5�
���d8C�*��fd�ʳo\�'5sV�T|0�١��q�Q7�� ����},��b��*{�B��2��\1}c��QlN'�#����szg�#\i��9�r�CaV�K�S�]򺮄(ۼ�^��0�۬�a}۬IP~�ݸ7)��n���S�Á5�t���7��ݜ���[�ʳLw���p�o5�BS�M��ߗ�J�z:^ �GcAܢ��u˔yMA��V���\( �6t�k�
�OW9���J.1<�(�څ5x�1<��G��+oU�Z5����7hC�E��q�*�l�N�U8I�/���`DZ�����Qa�W���ꙇ�{�����ڛ��J+�8h���I;�BOv��s"�&u3Q�*I'F�d��.�R�˖���j*,R~tŎ�2�ߺ�����V�Ō�O�j���w�8h���W�w���>�B֒��y�K_�WS���
Ƴw��U����Dd��E^�E��^^��7���f[3e����=6W��cP;87���Y
(Vu���{1
<�x��[, �c^O#^u��]{��ɰױ���s#���qd�!Q=4��A7)���T�RA��cx��C'f���6���h��:�Na�Ay�S�����!w�@�s�S��W���
�r��F��/ul5��{��q�-��Xa�<#�5$Gt7V�m?2=R��uyJ��\>�۬�S��/y�J��kA�	�>���cF��֍��jX����Ue���y�&���v��a�����AfcT���P�ZS<#B�1�������`<����¶*��Ы�T�b�gw���U,��ef�s�������:�s9>����ŉ��b}��r��U��x�H�0B]��B�B6�[�.��h����^�u�f�j�6���T�$��μ�͜1�v����Z�`Ǯ`�b���Su٪�(�N��.�}պ{(�Q���:n�����N�S���)v��j6��*0�QⲋIJ�mf��rTjSZ��&���gq�=���(�],��F-�E�\+-�R=�n�R�]�
���n�Xu�����DC�
`u�^p��%ӱ�\h2���][�s�Q��]=�c�9(��N7P����MO@l5�������4�$ȏr���a�x3pv�X�yM�O/���3yf��J��&Tm�syݥ�S�2=�|v���.h+Jf����t��R��H���\w������u����*gv�L�ʉ%N�W�5������������|�e�C��d�Y�8���f�:���V���V*�Y�����3�GB���׌���z�c�EDw<Ī�h��;Z�[5�nV�6�v8;�	�c��J��մ�k�.�.Z	�X�]�,7�0+�աʮ�c�!V6n�<³{��8���9Ⱥ�Ԙ�A�0l�6Ī��=D�K�K�κZ��$����ɛ����C'V�L�M������ig�l�up\+�균Ӧ��*�UL�;�����9��f�ЌPwƮ�ݕ���jqD��*��Z�k�R��.-���P=�+����ϙmVk�(���H��b������v��,Lt�9D�h�<�c5����7Ct�4�V��Y�Ln�Fl����c�Hkr�T�c�ō8��4�����Ux�b� �[��̂��<�K��w4��5e��5fu
�r�_
N�a�<�\�.�Ŭ�ꎌ���f�5c�tNj�#\F]�փ�u�3��t��r�Q��ǅ�od~�0�ɴ�����M�aY�!���i�Yd�+�8��u(�m3��!�b)c�/�����ʗ �Y���q���{�Wo�XXS¾j�n��x�� ��Zv�R��!B@]�e�#q������Ǯ�;���q�/LR-�,��6G�	�F��7�6+�۬��D_-twzTRT��'=�;��nkւC��(���y��0Y�+��MGa�a�խ����Tu�FS�%�-,���з(R*h�=p�]����
у;1X���Uل_8!�f��qa�ɤ�v��O2��3f
��-����k.�C�t���e�t��q+�^�e�*�'8�#g)�P�!A����V��{%�$T��c*���9Łd���j�Sm���yN'�N,[	̡��_����0���Z~�c]��_�:J��J����E�:�����l�m��öS��m��'(r"���B�L������x�f9����k|�H1��YyRĳE��ܠ��m���?�L�������o�{��=U>���KITQTm*��Q-b��U���j1��Z���#m�Q�(�
�F�V"ڥF�h��Ҋ��ʂV�[R�%,j�j�����
���E���F�Z���U��1VEEQ�(��������R�Ԣ����h�E"*,���EE�--���Z��D[j���Բ�,e(PTEJª�V�����DJ�%pH(bTfQV��DF%h�."��dbJ�
Aef7�Qj�4Q�b�)V",Rڬ�KkDZѭjX�j)Ej,D��DU+L�Ķ)b"�jU[jU@TPT��d\ʌ��q�ʰ�*�j�+
�b��UTr�U2�ȥ��m����J�D�B�Ȃ(*�cJ�U�Z��QD�J�R��9lX9KXVZ�QQ-�R�e��Zڵ����Qb�YUT��Z"���(ID�R|&�Y{��tg��`�ug�B����W��B���U��e� �a�3i�g%z�������Q9ߣ�����]�%�N>�] �\
�"�w蓴�ߝ��c=Pq���*�b����d�Wy'��f.R�l�;��s^�*dq�wUb/�cQ�E,����R����@g���	�s�g/s��α���>} 7i����b>������׆	H���A���Fޗ�wv��w�[�~S�dT+Tׯi�W�IO�5t-����np��eא�Ws�V����ĵr�w���b��/�)9�^ۗWL�6!�W���;g�k��ݪ�L��A��"��;ȱ���K�8K0�\�g������{}��}��U��Td蝺�	r��1�D���7J��{�] Q�fy��>��l�o�I��V��?�����0K,G�I�U��qx����ʊS�X�o<L�j�u��oVN��z�<%�G=î��DWsH�GNf�N-u��rZ�F.����&��q���1��Þ�2//���qSO����T���Si�Α��4�A�Saj�H�G��������F��b�L�8��(t9Q^2�N�Uog76$�ǆ)u=bC�9�p�_y�m옑{�Z��q���H,ظ:�����F���%Jx��gW�R3b��(9��1J6v��k���s�{9K*��W�gO0�XT�5�.�V>V�璑z�Bʙb=��t�_pZ��Ȳ.��G�#��ݴ6�.Y�P.����L��ã��cW@UÂ���w���^�	u�b#][�����=EƵG�Hm������P�5��/���z�
��	����P�l��g��7f��M�ҕ$���;�w
�T���.�#���i3�D+=
���X�oWaL
⛅t���OO�c�:P��	�]R����xJte�����:�Dz��݂��K�fx{���z�-��#�p=QȀ�	fH��#!\�#T�t@M�`u+�k8ɏ/����>ٱ�$!����r桋��"圂��S�|9�D��t��nC�:l����6�
�~�1nZ㞹>��/~��1	�,���/A���LJ.EtMwZI{e,��\����x�.��yq���@z}1�)��ٰ�G Hȅ΢Ey��%�,��ۍ��7�@�<S�3A[#�2UcdAH{�1��z`�:�^�w�Q��,�X�X]x=�Ya"�/�>��:=A�~ f�g^
Vn���P���'��}Ֆ�6�ض)2��8����3;0��Sh�(�Zݴ��1}�Wt7�C�]���E�6��Y�{B��[r��l��95	X�9N�r�L�Ͱ�#�AR�Voe1*�k�5Ad�\���Yj��m_m��dJ��]]06h����֋6c���G�=���۰�w;0Q�7'�R��5��l�=�f���F���u;V�á���%rӴs��m�8=�zw<���ъR��������|��^��2��Į�l�R8�3}ki%X:t�$V)�+�a3��aZ�dX��Lmº�b���t�3�1N6��\��'۳���a��^��d�'��+J���s��^b��hc�M�C���rUb1wl���/lAHu��������S5�|&/���6�!eupX9�A�y�KU^ʻ���{NW>K{yL�P!1�ap'�Dp(-f}�\�h�����Eo�R^�XS �UO��b����G6U!x�>�b�Rn:!��6C���W�1;H[Д�P�|D=�xq�irخ��{�����ӿ!�l��\����fA8s����;�t,��3E�[�ˢ}�n�(�nq�v�
9�	���a��0�������>�[m�v�3]�k�|�Gn��#*ʢ0Ss遡Y��,<��fAo���	��S�F�{�t����B)�݉���犷⛣s($jf�ۯ;�ƅ�:ۡ�ifҋIz�b�<���f%i��e�8*�i��u�uN��[ĵ^���m��.��;b���j<=D V�sؤ���j:�ʦ2wl��gC�K7�j��=�$��h�l�QVUc�ۅtU�K{ۼcG�V�77�&��{������o+W]KO����
�DC���(ԜпCX)�q��!�1�9���Y7�
'us-t�B���]j󃭜~
Ro}�قŋ�ݫ�і��Ԩk���(����s2G���*��4�)�y�h���߼߂Y��׋�T��C�A�TW��}��=~93�	�]��C����F%ª��TG��]�Ջ|Q��6�g�U)f�O�K��෼а��O��2���ZO�# u�Ȋy6L�#a��A�#b
��30�k{���$oU֊\�؎�b2���0������V^�ϸ`�r�v;]��V:
��ZҬП���ىy3ƃ�c�l�q��5�v@ucԒ�"�`��4��b�XOV���-t̎���`��$p��3�6�3&����LF�Ǒ�4#��(*�ir��8�C�<y�zk� �EE�:B� � *���
����<1eF�H����ڴ!��\�p��ⅻt��*�m�M!w�g���S�����;ϋ��mrԤ+ݫ�UqB6���x�]��Ez��ц_:�٬��n��Į�X��B悗��OYŷc��L�'Ry �$gz����8��Q�շʱR�?��DG��W��4�Qhh��P�<�~���-�j�unf�:!Ţ�"�bq:��z������Y�~���R>�҇@ѡ;y|:�jX^����.�r�pa��hB�X��Dfӌ�KD�]���q&l�˨�k�P�^;)��_B����=��l]y?)����)��,�E����53�W����R�F��Gv �%1bc�Ol�f��Lԋ{���8��%g;����g��ৣ�>���L b�PU�l�D�Va��=��{b��S=4�����B ��zh��"��\��`��fn�O���x�|�aY��w�E�ćS��P&#z@Nӛ�1p��B����A��Sμ,4pz���E_a�A����E#���}���z��e��������W ��{R�SS���</��Bxl"(#�����.u/fW�߭\�����بۗU�U+��.yT\䚁n��{�����bJu�_�N�M�*:�|iR6yV�;l��u���C9�t�\)p�<����K�GOS�C�=�Zmn�1�>�
�v1Wxyn�0��R	��th�
My���!�fJr��U�-[ہ"-؝�Fb�յ�N��6Gu�}Ľv��:��z�ַvÛG���3B�#7��lNj��'�Ok�U1*��,C�����  �0��s��V��U�a��X�/6H��/F�E�v�b�:V��?���J��2��U�CjEmu+�������T�4nD7Z:M��������d\��X�ҝML�0���7�{3b�]а�Hz�Ѷju�(j1�UF��jpn��Y\T���5t9�Oǰ,�/&��į�������ዲ�7�����Q�������4!Jg�ŐͱcV���uĚN�=J�+���v����R4*"�r5a�WW<+���fT�K�s�R9�f����K�0A�A��V3"l��bxީ��u^�	����RȪ�c%dl�輎S��m]�2S�u��Q���q����;�I�m�Q���?<�������cR6�)̍��9^�il��)�^ߩ=���tLAI��1w
�xU�l�u-\v�ץ��N��H=�y6�1x���v�����Ż�W��M@��r *�Y���zP��U�c8�.B`�^��� )Ý��56;���D%<!ܹ�b�^�E�g�'�x��4Fx���v�̤Z�W�J+���uһ3�2n��6�\-��$�H��}�ňOo3��ufWy(���U�B�w6�2@Z�ԋH�͈����:�P��W3a�]����X޵u	a�Z��FwC����
�4}�-��Y�h�z̭��+�hе.K�酃W���ޏz=�JTu���!�1C�61\LF��V9zz�7� �T'8����X�S�f���u��̛<D^\��ΊE�t��3�a�6!�M�"����tXp9F.u&��n��{U�H<��;�e"g�j��턘�^#]\K�=Ư�a>�є���P���(*�<�^�ƪU�ӣd�v�Aق߂���9>K8ؔ�A�,خuVUM.�£�5��ktr��KJMT����>��<�S�i����O�u⍜l�3��9P�޹sJ���걷��{E��<��t�Urы�N�zۼ���f�Q�9�#��V�T��,͛�Z�9��T]d�輞�Eb�B��;q6DZV��s����:b�'B�i�����\��/��}��`5k����O��>�
|�C�v�D:}lv�l���^Y!�[U��#D�%��ݨP�Pv�S�b�	���n8�0����
oh7$I�Ր�w{Yǋ��Y����n�l�Ä�*8�
ٟ`VbE���;��IWυ����c��f�X��S{]#F'��c�ڢ)������ɯ��$�x4�:Y�gyM��ܻ��)��^|8=�ݮ����K��)M�\�켦;U�bwB��0�K��P��^�uQ�nG)gA�-��Y1vHl���L F�cM�u��	�����ވ�z�j+��v������,C�;\/؝>��t�ۧD8�$r&�Έ@�S+M�J˚mq޲���s�iG)�7�gO
�C�N��F�lf���O�l9�`���Q��q������J�j�<�����{d�GEDT��O3��h���5���a��0���&v�̉�]��Og0���z�-����3�Fu�D`���4+9�{�v�3�FC^׈X`�awIv����r\��q|���:R8����xʲN�"���Bgc�M���	��ګ{z�e(�՛Z�rU�ƴ�36#��(����q�"���3٩V@���WEw��^C� �"]�F���T����g�L+��.�}V>���_c$_�UD.�vL���Ӂ�P�g����ҍ����yeA����=�ܫ,V|h�fOUPY�-�w��di��&�����0����ϐ���u�������^L���d�\3Q��n2�A�R�,��m\�h#��\�����tPu�W�T�}>S�N�`�MZ沷�nY����GdvK�4L\c0P�͛MRȕ��W^��n� �v��]q��eݞ����5O��õt]ek�&;�9���Nǋ��I�h����1�f��zk�2��wv�q�k����D��?��	R<-gR��P�8�)��������]7�x�Tl1�i�����JɯEt�P/�|�,�q��\WdV<����U\�Ә�s����rj�v��낛��@����������P�0{��S�Q�^�pp´�� rZ@�=Ȅ�NY��,!n�>1��ɸ䨎�fipx ��:<��!�-L+�1�e�T����\֝���s[�"�!ZU��w	��Pr�Ij� �|i`�Fd؅�^��u���jxP��.徖�?y¢1�^�n���R��Fb,)4����3�-��Ќ�.�K��$�>�s���y|:�����+�Y1�cV�K�����z��5���ѠX���>X:����ʗ�}1���S��c�t�!��hk�ɖ�vP�f0y
��D&:X8�Rp苁8Js�)�¢iН���O9X�W\���.�p𢲲$���,ϓ�����=kh/v.�,WI�}�Lf�vŅǢz��̻kZح��p��i
��1d��'%z��&5��W�uf��I���&�"��9��u�^�[#m�ҷ�s�	1�y{:��Y![�49.˘juƹf�K�^�]�Zv�D���J���́���&H���;7 �톟��!��-2Gpd;�vXd�\jԋ37c�;��V�U���������MY��شV@k�,��+��3R��
��u�騹�:�0'^����+r��4P�2"�k�V���Eu�k�,z}���*�챑�6���x%�cu8o�v�dQ��4��`���Hꌹ��5/+�&�ў��-S!��s�Թ�Ї\Ĩɵ�d=�� �ɭ�U��L�h@�f�������9�e|��\G絰w���]�7_yO�nq.����>�n�'�Ło�w�����OWU�W�}���=������N�!�5�ژ�T�4ny���n!��?'�gxt[b�<*��d���5�V���tqr�P�Ӛx1!77�4ۯ]�9Aq��uMz5dm9��gJe��]��wݡ�޵ܻz`k��CȊn�^������g;�)��p��s�ofK�ܗ�<-��P���f�Z'�L��_\KF�z�r5f�aW 8V5���[U�z�{ ��l�J�A,ƈp+�=L�8�E���<r�T]�B{:�y~��ގ���o�LԁVV^4#v��'����2Ƭ��E��f��c�c-+�S��\@;X���sR��t�A{����CE���$Ѹs	[{:�y�a"��b�z
_W�dO2��q���9�m*�&���<]DK��Q���� ܮ����T�����/D���Lˍ뺨՜�����
�au�4�r�݄�;��g]u�{p �m�r�Ha�E�w�q4�=Q����ј�4�� ��I[�ŰI�:�n�7(�{�.�=xt8�9�[&Ӷ
��/�+��\�����Xt4���sB�%��/iV���$�I����hU���}��6'�ؙ�hܤ�:��]"9Ij�F�**J�v:�)����^F��m[�#6h�]3�:`LG|����ݐ��x�^�v�8��Cʗ
5�qvQޣʢ�{%dٗ�w`ʗ]��<y��[H,��&��=vz����M���S1��30��øX�օB�X�|:��>�� ��MN/z��AZ'�V�ZLF�na;+��V��Q��3\T��-4@�K~d�v�f�2�؆�E0�4�<U��_-l�4|żN�9)w:{3�Mצ�;�;�ɨeLIr�L�9͓y����kE��ۤ)P��T�fXS��G��Ӫ���n8��D�X��L�lC�؎��T��5�Gƴ��;v2?,���[���w�����N?�i�d�%Ŗ���%�&�X��R(\u��[ͽ+x�ŷ���)Xj�+�a\�]��ʖ d�0ȫy�k�U��RJ��Q�\���9�R�#�Q_;� �l�@Y�����]}Pc?XYkj%���6�GW����˺%fe���3Q����<�ec l�%���� �y����zI�dT�o/�,�
wҤ'��@5]�(�G,Eq`��Gx+GW���5C��M{�N���y����&�D��7
���6:�r�.چ��;;`�v�[,'E��1L��/3�ܮ����k��7ۣ�v�m;��Zh�`�D���ʬ�q��R`�гe�9r�%F�]6\>=���>0�+O#S[�:X�|33h��n�\���V��́�G`�M *�q�E�$C �o�=����5ô���LhF�[��	]��a�j�wZ!��K���zp�ڨ�^���D�ƋwD,�] �effN�u�P(�p��0�[��U�-&pİ!U���[w!n����ķ�k�^�a��O���G(2+��Ǥ�tu�ķ})SY�T,��̠�L�e.ͪ��[�*� (X<!�Σ����*�ڼG�u�L*�,�T�3QY��](L��I�� ,eJ�ѭ�-���ꄌ#$��Q�%�Uk(��ֲ�m#[j�Eb5-�Z�Q<L�)+m�aP�Km�cf*[J
��F�6����X�b([b�*�*��X���`[bZР�Z��iZ�j�-�2�j�ձX(��h�Af\���mDb����R�-J�K+e�"�[h��Q�D`��UQ�DA�V5�Zʒ�EEXUJ)j�A�)VҢ�(
e��*ck�8�H����FR�
���Km�e�A[cl--DH���EH�keR�Rҋl��%b-�D*[Q[�m��[E�#b�eEX��G,EDJ�V#�k[,�EQ֨Q
�X�X�q
+�*�X��V�hTXV
�lڵ���)��jJ���X��-����a[mD�Zص�Z�TT��`�VT�F�FSD<I"���o,����	�ovf-�o�j�{������tE�YG�s�֞�����=;�s�+,�ø`�;���{�i�&�A���ي��w��p��X`�nH������;�dT���,�59��ҙZk-}���N+W�1ʭ�+�kͽ���ɀ�ʢ:Ux��W����g�(<��s|�	�[��⻺T��\���8*hw����`5Ր=���@3e�2.�b7��\昿g(�(W���P�y [��xY�W��b�)��.j�/�.Y¦�Wς5k:�$�J�<�7LK��q��&���"}��L��/Od@4�� 1	�2��C�U��l�� 3N�@S��ӻ��a,�t�կ���+�PxhZ}�S5�:,8��$�Y�۴�g�Hñ�'9��ۘ����̓�����^#]\K!��ի}�v:�c�k]�϶��i��6�#�u�~��@����/�7U�Tz��+�i��q�(<%�ƯU�>�םÝ�~���6Eܣ*�nq���.w����o�H߼���~�ߞ��f��Tg�W#�,���*�Ѓ�Ɇ4\�C/����l�ڧz=~n��NC1�T#Z�Ĺ��m�_�[�R���M�
��%d��8U���J���̰����wS�E�����k�Q]wE��<v5�]�u��)wӅ��6+�j^��2"CI���H�L�������n��xtW�����9��v�C}@g$��:D����z=��֎�w��O ���ި=R�i!��W�7���U;�3�i�TnD)с=n^��v��"�o�rS�MO���o�����Q'��wTj�7�+ʭW���Z�p��(����sj�iY�"і���'�o����%�T�Wӗ�Ny�V��\�kb�� i��L�s�[֩�������v0Ɖ�q��3�
�ċE_�hucw��8�a˹Q���Gwxi�ŷ,Ak�
�j�O�R�n����Ț�3�����`]�,�ʹ6c����B��V,]:���:x`�s��u�1�aƼ��O�3��=X��o�I���S�3�tk����5�p:8��n���Ɔ7i;�3��v�)Gm�Em����=3=��R������4`y����E�
�@�1e��Ҩ��\G+C�2��53��������]�W]!�R�;��x� Q��[Aߕ��M�n���Ȉ�8߹���﫞k�|f�z���Ɏ�g����+�`�bU�<���1��"��e�Q�}�T�x6���T6�f���IŊ��͘�}:�X�Z�Y&qk�U�o�����Si=��/�Ix�������`X�z�qє�
6�6���AYUXG9��s�w���2�،/�;F�&����vl9��9��7(�ך���FÊ.�h`���'����Lݼ9�t�e_�R��U_UPp����ʥ�?��(:���jq�]�a\n�b�t	}��g���$#�X�f��[.#���]�]����A?)�zc�A��no-�#�����˚6���^fOfz�g��f��T3�G���!l�{R0Tk�!5�V�:�Ey&�=�s"6M�=H��0@� 壕��w;m$��W��8,^�T�z�`c��ev��,F��؊N�`�MZOe^�g�:]�^�zv%��[9��.�IUh�y^�G�O��:����@wM�z{|��`��::5�2��Q8�K�0��i���8N�*�R�d8Uy�q3'�CPk�i\�,F=�b�+鞾K5�R_\�-�r�i�&�I��6uêB�@죃�	jc����v_�+3>��4� �ӛ���!�*�k��i�(g�K�p�`W�4��3=Qs�����<�NGus\�v�S�O�ԱB�徜nXb�½�
�_��s6�пVf+^�H��;�x�BN�s
��յN-�Vq�"�]��GՎu4&�k;�s�sڻ��^n�ܮ
���>s��7!qv��	-<�|�ka��T�FZ��
S2]+�#�x�G~���Ӓ.V6xva��D}����ڏuvu��"�m���f���	���DG���R�+��Ӕ*��C��铍s���.���x�G�qw��U��֏w&����b����9ޠ�m��6c���TB�g����9�0芉�8i9��
�j�eCx\[��N���p�F��	g�b����+�E_K5���;���z��Sq��u-��6�ޔ�!j����g�%�p��p�7䐬!���c`kǦ�ۆUX�#Q�3:-�j%����.�[�5@9��z(\S�m
�l���s{F.��a	'\²�s8���3c,Zi��D��Xq.^L���[��}����x|�y�C�s�U^�Or���z����T�=��h��<Y1y3�,��N�L��9��Ǉ�`���u�T}��u^	�Ú���Vɫ�:�g��ø��.������.�>�*gd�mRb�9%����j�T��jvS��2���X�Z7~�n�b�:V��Ac܀� � �R��.n���L��/�A�q���E�*w7<�h�6�`t�h�FsO����e��Z6W�����X�Ww�]]Z�A�8l�5�9v�o�w1%ir���9�l���Y�*d�y����¦�TZ�2#���
���寴�\�ͤ�`:�s��[w����ѕ6�]��w4�������o��j�Q]�WY�GE6z�'\�x{�Þ�\խ��]n�~�,��P�#��Fٯ6��nP\cr�4�#k<��eF�F��r�{�KO0��F�����(��0��9��W�����E<�3�Dc0�����5��k&���v�O.fA�}6ŋ�*+�M@J�TWTFK�0d�hC��F������}���h���E3Z+�:կ���y�p��-.�g:���8�m
�k�R�6���ٲ�y��L�9��=k��A`_Wh�`���D�c�uniU�B�$�����S��N��.�X�[^P���b���2:x��Ux�Y�����]p$.�#kh��V��^���߫5ƬK7U�)��+�W�1e�d[j�PX�͗zPzc5��aL��w��<.�,z� fd�xY�X;�:��0��.Y�*h���NȠQ�S�{�������4�'r�DX�޺_`59�y{�H��*����0$���)=Rn�m��������TF}�_6Va��6!fM�6��٬�� �vQ�D�	�u�� �l;N@�u��L�N�1
�Q�Vٛ��^qe^kbM�;�����Li������g��%E+���Ի�tfkp׶�)���n<rk�V�습�y�el����ˑ�ö�ߐ�����+�:,����DB�\��m�n-pĦqG��D/��i=\X8}�&6x�ur��E�q��X���q5p=���^m�͘4+kMmݎ��ሾ�_�P��T���u�nQ�6<PxN��8�;fF�r�%3���G�2�̒��Uu�4��gJgt�C���Q6���3^�fN�Lͥ_��Yܛ���?{����W��a�%���AU�f.�S��n����c��}�^�0�9����wB�Ub��D������i!ߕpu������h��j�϶�p��n̮g��L��))��#B���
�3}h7='����y�h��U�9���t\�L�iߧ;�s��z���,��x�Ù��z*�ۂ�]�[7�U��+zғ]�ֺ��M���:��u��5K��u�ɸ��I�5�^�_A|{"cq���s�`��ۜ�;\����E�������y�LA��ԅF5G��#ғq�����a��v���5�vE��U��!�Jzx^x�s���¹��ӿ!Q�F[�(�R�]oX��`�>їp��^S��Ծ2Bk�Q��b��^U)F0���y�x$AUW��v�3��M��p�ͳ8�y��tH��M�ě7%*�j��k2J\*��������'���X��'|1�t�r$�N�FuA�d�IN=��u��������KeS�O�ڱ�ŌF�*��W��ƣ��vS7���A���m'p�3p!ݝ�x+��绒lw=;��A���C��g���gb��
��	��#B��/ܭe�҇�"���`>9��	��+�ϝY*��X!H�Q;魋�&�d�wB��^B�vU�˦�<��5���^,S���6ǒ��@�6!�>�||��-x-�����,X�3�K�������(�=U}o�J^5ڞ�>�S
�d��t}��g��&�z3�p� |���dF#�̈́��x��3��j�ʃ�y����4oݔ����>+��>^�s�I���D�G� �vg΍��H���|��&<��נ��c���R�"�y�KL
���k�S���D�?t�p�da�t�9F('�Z,.i��b-�'x0=�)��%��>���]�+�ڗᣁ)�x����^���P��d+t�������kup�֬f��e!����~�T�x�)�����<w	*����@����};����ǝ��Z{ԥ$��b������<����g *z\e��zrV��.nA���H���������^� �7��ӵ��îV2`�Oms9�r��`n[�v���=�`q�qt���R��	\K"ʶ(�"�$,�b]��V�謉�������UW�G��>}��6�V]�qނ�ٸjXB�:�a�v�:��.5����@J}���p����!�A��|�&�k��7<����B,!ZU�um�>(c��2oЌH�|i���Ê��r�u)΁�fM�N"��b�!w���-�P�W���7V�x;��WFK�ś������f"}ob������N���:��w\:�Cj�c*��J�q9ӝ�/���։����,���u�OV��6qdE�[5%v[7�1�^�2�* �s�r��Hnp�(X�N��T%��y�<��$-g��~�=�r�â�!9���k������1�K�����y��b�^V@��݂"�[v)	�;���O�ܫc3Ov��U�%0 �6#\�}� �siD�w�_��"`S4zh��S��5�iWRꓼ-���Y=���	����4���1ފ�,F�0�Nl���s{F.��p�u��O��΋0B��t3=1V�A��Vq��0~�7�q_�f?����/�Vo2}���5x! o�=�����fL�C�&nU��4`�9Mm1fy�V�-�תt�/7�`T��aM�&�B����c���,79;�ufK�{	�æS�M�����r&�v,��X�cg��}�`��K�#�f�������\�ݑ�/�f	@�V_��W���xu�W�O�:�{r�*�*����0Z��z��;�j�X���ۡ~���5mV=6�xh�;���4j��+�,s�+�e�h�klu�\:�r�Suk���5��^�j��ͅ9h����I���(�ED��Z;n�ʬ�ތ�h*Hg��!#H�,E��BJ��S�ѭ�G�h�����^ORn^U�"�ؼ�J��n��C���߸�5���9Aq�U1��6���Uv�1�k/{��3w'>��>�b�|%&�G��Y�dN��+�C����S�c=}������<u�i��V�j����Ni�,2�}���ʢ���ѱ�9�j�
�pSQ�j�{��X��_,�q�_-�08�´,N����c�(2�|DN3�
�����R_�p�:ode����w?q����_�&:P��3���oHۢ=\x k������zͣ5l��$�ft��fk��缔q����n#�xC�<X�[^M�,g��`*�*�W�f���*�������%����+��RAr��iu4 7ԑ8�%-��g��/z�.�YWv��1ɒ�,����1������IqXZ��Lwz��z($#��g�W)�+��ud2v� �^˹���� ���I���}B$�6��i��&�	a�������ኖ�����Z��v�SF��{�4:g���@;gչ-��s���<b�^�@��6��5��n�{��@kk��s��5��22�Z.�k��'%3���C	t����0lT�
k3��c{(]N�-!Jx��l��i_t��4�'r�%&��_΢4,4.1���"+�ʀc�/��Wٛ'v���.�伈
hx�\��ӰgK�"�R����@X}�S4��i��O�"�RB���,���H��W/���wM���������΋Hh�F�K���Y��&jsSJ+��rzO��c������E-��P����;~����ݰPί;ɜ��X�q�b�%8+��;Iׅ{����
��>x�!�ߝ��د>���J/�n�j�<D��7[6ȿd�B�!�d���9��59y��=�sq3Ĵ�20޶󒘡8g��soĂ��
-O7��;~鰭*B��ӥ�2��
Xr��{��n�Ց�!�i��p�G	�o����R|�Wt�Ɲ��������=��*i˭�aT:}׈�ư��B�P���G�v�_�{�_h�4Z��.�q��AM�eon�!�Y�a�,�Qӣ���7�e���+�F��ϸhm�!�آ�ڜq�2�C+D�R]zW�U�L�X�u��PX{Q1W/��v�N����і�n��	�7yb��I����mh:EDH���̓<�w�S\sd.�w)]�(��E�
��zr�sU�G[�5i���qH>X��sYja.�]��dEρ�Fun4Lns�f�U��0�f�����]S�ﰃ�^v��/KY��0���=�+���Z/��nS���ӨZ�@vq��G`ȭU���(1X�%p���h���J��8X���v��vήn�E"��jȾ��'���d֘砼��֭�K�!YCf�䝾��Q)�3�����u4:���쪝�3q���܃�7E�gkO�!�t��o\�׍ٽB�M̮zUJ������w���`'�11�<�ȼ"�	AGOk�ovG�T�^��m�1f��o�n�h�dS�Gٳ�Q�5DD9ȕ�i���[[�$tˏkY��n�A�d�UD�v,R(+�Y�b�����r�����ˌ����҇6)��
����U��
`�t�]�v%Zε���]>H�w���K�M��M�	и���!���@��B�콘�r��4JLKd�G\�M�:"蠨�*X��L��|�3ٻ&�#��q,�,�v9j�JJ��W��^��Uv�^�F�(�t�YVOb��+ݺ��(�X�u���d�7�E�w���-1unMX�V�ֲ��g�Y}�*A�W	�Ł��b���ʽ�U��E�g/\P�/$�U�}�.e���[x9��(^i'�͕��fb}N�nօ��k;�S:���n������ZN!b� �՜ҭT��k:ͽ�+���=��A�"�+��w:�»gv>@f-�M�Qc�Z&q�i�Zصq^ږt����jl]vx�O%�[���cz%b��b����/S�3e��^�ys�;m+�n�k8��NĘ��EE�0��r�մ�+����>�7�m<N��sp�y���� 
�@�;K��'S'�w`NU�����r���� �u&w�v���r7n���i<wB�MLCU�ppɖ���q��<;���L��R��7�@��sm�e]%��̪�vU*7�Q\:��EuT���n��㺵9cbL,p���L��7�a�	l���n����ǚZwa`dAֺ
ݡ�mM&��̱/{��,�� 8�n������i�E��2��(��\�L(h��7�Чn�\�d�kfWS�r��#�5����oA�=�q��maqO�5wO.�d#лw$��V�ױ�b��V�K���5�XF������{8^��7�w���E�%*�1z\(uD�B1w�ؔ��e�4M;�'ۀ�-��y�z���-��}�j�p��=������X��p���wK��qh�J֣��!��{�.Ud����"���N�|U�n����v~�M�[j[jR�Ԫ��UEV��(ʖ �kE���1-��)TdD%�[F�Q�Z��k���(�LE(��Pm
2(�a�0�5�aj+aP�,b�UB(�#�EPU��
���4*�j�DU*U@ZԖ�ցR�mj��QQd����5�-�Z�,�jLTUTAV�r�e"�[%ʱL��,TLdm��\R�UZ��ʸ���T�ekk�n(�dĬnSQ�Fc
�eEF�m�*�����2�L1�,�,QQ��.Z�R�� �J�0W�̵�.7����dQ�m(�Eb,-mE���R\�����3)EG-�`�V(�dV���ؠ�������ES-�.Z�m���.Z�,PX�堲9IbD�B��3*�VcEWp�V"�E��(�EQ*U�Qb��b�R1��R�D�q�Ɉ"�f+1kd�e�,��"���*�JS9Hd��/����cM(+��1��ty�ǘ����6�.�����Θ,B��J|�lPZC��S�PN��!�C�mS�9�Uan����cb�-�oL�>����O�f�7����)I�$�[��~�OoY�N�=�41S<Ca���G�B�D���.�-��|����#-9�Eq�a+�������)C����xO��:����tiǳ��7�7V�k�sun��'��.�:���XS9��vܫcQ�>�WE�D8 r&�m�<����|����"��1z]��oi����D^Ό�t:�'~B�^��5ܘ2s	'�4�or�7�
���q�>�^��e3�y�4PR�G�C!�Udv��J��)\����9�U��(�OW�y��f@�r@�6�Dh�wAa�U�lJ5�PĬ��:mlT�Vd�������U�WG��ߦ��T��!��X�:�����O���EW�Z���0�D������9�g	�b��k����Fq�)I��+��,X>T[�̲`�x�l�K<]���T��V�:V�bd^����ݩ�=��\v��>�~}�f�S�~��vib�t,**�1�{nt]��;0�A��n�ʃ�<ΏT=���qNk�sI�=�RxE
1B^�	q9$���I��$�Y	��#�v{@Jx"�k�,�,N|n���:[RjdUd�C3�+s�i��,L�R�%A�M[Rںڹ%C*4��K�4���`�7��a��
]j0V��Q�A�Z��u�k{2o������Ϝ�93"�fɕ�cDj#���Xo�b�y:(+�+IE��o-�)��7�s�X�v�]���mZ沶zph�CM�ϼU���N��:���(V�Qsg���o�N�kZ#(�q�c�گb�Y�W���o��8$p��g�m�&b�D�An'V"Fa�Ъͻ��>�	(/ϩ�SH�8��Pܰ�çO�d:�&��Q�J�OU��=T������K9,�#�i�5��b�1q֩��iW5�u�����v�̛���f*�`�I5�=��=���z�ɱ}S�(V\P�-��,0���z��.���z_��O�P�Ix.�|�/k�FԮ*�T�|o�]�u��"��|>ʧ��w�>F\��:jV8՞6ޒ���#���	��L�}ΠkUѬB�v����j�����C�d\ʞ�����čO�P�	�R]�c��Lp�T�v�0t�=Da��P�z�(��ܢ��3w�;F���;��T�M9�K�,`�;q��p��vm�� P�TSR� %޲���:f��Y�J�5���mrV�\'8{!��(n�y��"����d*���J�h�&@]-{����4�Y�V����$���Z��}Y���B����paQU �Xn��!2Ɨ��%d7v�y�(O9�,B�<tSt�����^3�\"�d������7�l;�s^���K ;��� �����7i:��P�듾Y1�a��&qX�^�5_�E�Y>���@7p��ы��nD^ve�Pje��ws������E���~c��c����(=��O�ټ�";��YQץ�v�w���c�Zk��x�������Uк<'J��
w���z�1�vGuНN�,�8��z]�v�����c�����e�E�s�V�U�l$X�M񫨓)9�4�N�蝡��U�b3~L���)��{x84t>��d��"{�ɠ�[��䘃�[�&V%x&�J*�@h��q$$xK,F�q�k�r~N�F�t����X��NJj&�3�r��ǈ5�����(z�mV�q��@����6�y�^�r���cpԆ3o�	�jy5���#y�W���P�p�U~Ʉ=>�t����~�}�����{��=6���>�����e�c�}�aį^�e_Z��:b�#.�ߗ��+)W��)זr�ư�g6�r:�r�W�B�f'.�f�Ζ��;�����7V���N�dANɏ@�]�BՕ�{C�BVx�LO-�:{lu�M=��j�I^tЍ{:�"x[�Q>�&�%p�+�Z47�x!bչƲּ�
�Iy�[8���hf� �B��+Ggΰ�p�b:e~g����,�� �U�	>�V*���ob�.[����	d<�pw�3ԅ��du�W�@���8�@�a�²��7)�����0�.]j<���V�V�Z_�Ϫ���=��,*+����7�p����,�![3Cu���}B��۠S���-���h�U>��C�wC��!C��ƅ*�k�d�w_C�o��=_���@e�cGx���	)B�0�	�����XZ�P�]��OL)��S�3��F�g*Ț�	��륗A�c�G_(�T�=��q'��oub�@B���jMeP���X.�^[O��Yu�6!e�`b�->��po��&�+�n���i�(2��H]��LJ�g�r������duF\L�^�41�VBxC�ƶ��'�|���� 6��);���!nW���S k�gFߙ��ޜ�4u��B���� ��{�v� #��yƸ��<<|��쿻����|�`�DJ��5��â�Q|i�A](u-�G\��g��u,�pM;7F�����e�Fu��m4�}n=�)���a9>7���*K[G�m����W.�(�l���8!�����8"Y�N�+���������=��^똳Y��Gtb�m%;堞8e�Ͳ/'C��[R�܈4��R�H{���8��c�*�jg�%q�ۣ��N�\C����̼7Ɜ
2
�E�dF��v��aHSU�\�ы/�ނ������b��8,G	�F���n*��u^Vɴ=��Ѓ�E
)*3n��|�׻���]��ܴ{ ��f���a��6!�
�v॑QL��3S��s�\��IXK��g���m�g��,�ν^Ʃq[�wZ�Ģ*8� n�3ݑ����^��a�k�Ɗ�N��%qx��6S/����BU�z-?]c]��ȏT��o�"�`6''v}/����L`�58�4ƪX�]��jb��s���w�+���3ؼ�@箛�D΅���U�Jv�qŹ^s5�;)����68X�d-������*f��4sf(=s�!cU�{E#q=^�c9FU�	�N�P4+;�oe�ޮ�b��W/nR{t�C�b�H޲g/4	��� .�c��f�a�X�V&qt
�y��X4�%���ձ����Y�}�%[�)��8:�Y��0d76Y5��\��WP��O-�&`���)�f�W��ou�p�ܲ�y�*�ws�����*8�����S�ѐ���&�]��!\Q�q75��,̋)���͚D��R�>j�p��V�5�&ø�s��P��O����N��U�ggW@��
�h�r]��m� ;u�W�U�u��������1.D��?�ϺVEW<��5=�(&�}IA�Æe�h�{u�Za@���no-�#���{YsD�㙸�\�$��1��P��>��.��a�N
]�#k�!<d<Iނ6=v9�Y�Z��������P"r늫��aY��;������`������	�N���T�^��3�eoT�@����p+�9^ۈ���xHP2,�M��+Z\b3��R�.{���=Lo����7�W�mL��=��h�y��9d���h��T�O|�ĺ$���}�nC�ȧV����Pj3���U�)���-ӧ�1��:o��;2�,��Q�rX������F��f�71}j����iV5�u�{ν���^D�i�k�23�{��.�&��*�u���}�J[�ᩬ'��\A|�Sss�p=P\��������M�sq�:���ۿ��X��	h�^�c)Y��]�'����j�f���:�|����
��z&m���w6')7�Br���-��I&�$�>Z�.�ʡZ4�T��w��%�P��b�=�ک�
��6��0��Qw-��2�(*_P1��+)�o.7ùb��z���)U�̏T⪔�|n��g��f,�����zUe�22@��q�J�����:4G^*���pw�=��Vk�M���SĎ��zx��⮔��rձ�8^c��pb{��b�*��:�Q
��S��k���DoEF��/��+W�� ��Iί����gn JbĄ����n�Px}؎>
�0�����V2D�־�M3��j�� l�،�[>�S���l;��A����Жѽl5��\gL�n����mP�v`���of+�%���0�Tq��sj�qە@�?x/Na󙢓�����r��~�N��Og^��8Ҩ:*��26�LN�<7bf7��m��$�	n�%{��jW��B���1Փ\�б��*��N��{�k�K��ѥ<����l����֏Z{R+�2�M\5XT߫�h�TH�P��V���Oɯ,��*\u�UVP�Q�ӛ�O@.�8�̈́ٷ���t1�A
�Ք��Z�X�&[Iw�g�_�3�jg���F�eT�e�RK쾵�otX����@Y���Z�ʻ��e���BVn��BL�5�w�������ὑb���gw �Z�X�T��{[��U��)X��OE�<��Z�aݎ���T�s�nw&��k��(�@��ps��!�\i�"��5%1v��G�8;��������5�ڂz�=}ѱެ*���֮9�T^8H����F�mϫa��h�q�]��&�e-���w]M�&�mA�n��j�}� L���0���ΐ��\T|h}��Kef>�6��岺4?4��n)C��
ő�.!ʊ�,UՔѱqc����C��&��,t���[*_o�������
�����p��e~gi��6��Q��~��� F�鸣T-�b��t7�/�(C�l��XH6H�i@�3�V��kո���*rOrJ�y���[��(;� ��,^WW��<X�ɁII�fcQ�4�+1b}�|�Ϲ��u�+�u���Cƙ�S� ���l��\�O�A{Y�4g��+����Ŵ�-� �\z�l�"��k��1Te�)��ʰvA����3M��k:�t�D]�s�vA	���ٜm��D�꾝C�u23��¨m�;U��Ӕ�s�*������ol8c�Z���o��U�޻)D�92�{��W�z��
���՛�]kB&�Zm,���KPDs;��9�ᣮc�KT�ۆ���V�'<��d�|����l7b�dXU�mZ9`9��
]+L���PΝ)%=�ۊ�9����U$k155��D��Ҫ�jN�įY�׊���&��J&{�Gf5I�C��DW��Y�qW����+�_Ŝ`��WH�1j2�`]9Ke���e�Y5���
����Q"�ꍒ��н.	���ꌸ��b�k)V�2�8��ڼx҅]����lת͆�`��P������t�s����ܨ���,|�����ʤ���q1�PWmB�Z���e9�^��t�D3xbA���]�:�S�9�1����N���ߧX;U�9�6�á��0�
��h��4bg&X���b�ђ**�a$��P��;��9�1~/	�y>�QK�c�T�o	�\%�xxE�n�[/uK�GJ�r�����������ECs��d���}h\D��<�_����.��؎;y��w4�U�q�>�py�}���1�dr3Q�U��.��G�B�L��Hp�)�bt��|V��zT��v}e�x?�>�J�ࣜ����:�%���2���г8�`0uh�RҌ#��r^eng6�\�+����G*�U�(-d̠��c����5E�otc�W��7S��p=H����c�<��Y��^6vmd��yχ �:�̽�"�I+dx=�ّ|]�.h,N��JBl�-�B�	�g��� �S��6{v%������������#` �qgD!~�ʸ1C�Ӵ���jaj�0H���;�-��74A}�?'�>>�j�;�NZ*��<����`������+�3��
8鉺����v�������8�X������3~�QH�T�xS;X�z��
�@�iϵ
��F�U�]=v�%��٦/���T�^׈W���X%�z�;��Mm���"�fkz&�eiwSKRF��f����1p"Cf��&øNi�'��v�q���dV�<�hr��鉱��c��!��]�.0���y�UZ}�Ĭ��h���r�.�q�h{S��s�9N�6�Y����Ϲ�FO�7]�N.S�e/o��WU�Şpk��n�gG���v��.zfsw�Y*T�q�8Lu�5��'��d��g.ڑ���|���nW�1Y{W<���r�S`����0t�U�k�!��g�署c�-���Vc��t�u�td��T.�KZ�J�^�udz���԰\2�6Hr�L��Q���"��e���W� 4Uʔ�g6&���^���o��^�6��$�>tS`�5��u��:��Mj#�P��l񷝤^ֺ:��k.�vw2��9`��fc��˷����FE����b�B�Ŵd��va����g��*���m�������f>z]\ήؕ{M�,d�q�u�ξ�v�/���3m�v	
������=w���hV�I���_g-y֞�v�>9�1g�5T�n� a·.a
��HZ˼sA���ԾT�i5{gt>�Ƿ��<�3/Xq[ji����c�+m*E�W�&f�@L7�r���P�Bu/p�7�8]ͫدkzQ�t-�V殠�mt8�XJf������=�_vd���7��9���A�m���"���^Һ�@�']�)�Π���a9��#KF�Yy �+g�b�{Y0�wy-��j9��壮ʩ.r�U�-�$�!iV�*�f�ݚ)�	�����7���1HVf��_�%� ^�bd`C�\oa�1Wr��1,S3^D�m��	�n�j�ɉ�27��m��\H�Cz�ڼZhvd�B��I�:���h��1�}�5��#�/��ޤ'�ம{�mŽsz"N�t{a��g7���9�Ԁq�E%%)T]6��c�^��Q$9�%W=*n,���!�A�����c�.�jsm�ز�'u*�bޤ��yS�G���h��f���\p]�mk�U�֑n'1-��YdMN!�;ʖf�wy�b�����[��yNO7fc���2 |z�ح��%HU���JKu;H�q�m�Hp�W�"\��l�����X�8HZ���ݛF
�V9
:Y�r�����ͭڊe�Fb���h��2e���9��X��K
��6�흘衔��ɪ�<�O5��\1NP�N�gl��t�%d�;����!V�U��pK_o�,�n�Q��ָ�ؤ�\�Ll�Kol���Z��k�\R�w C����F�A�7e��b]�pu:��v��h��fB^�ὺR��wp]f�Yv�+�Cd�-�"���!�0�Ac��3�U��Vƹ'@�ն	�(�ڰQ[�$�
���uk�s/M+=�3z���q����DӋT�?��"�ȳ>u T�o]����H�=�Mr�[�@�_l���Cl�qʈ^%GAk���oe�uw� ��[�}pXZ�Cl�+_����H�ͭ=n+���[��������f�Twna���[�x��o7�����9��V���^9Kr����]���wt��vd���
���Jm<7y�P�̥z�w �sa��M���6-e���*5v�_� �����=�6(1����v�Y����\�Z+��-FCZ���	�`�f�6�ț`2�c�~��Z��}�d��*�cDE�j����b�(���[E��1�j�T\���PFUK�r�YUQ��J�&6Ш��""9f2�akJȨ��T�aTQ��eb0��Qr� ��J�*"��ʹ�Ա�P1�X�̹m���L�̂*��\eeks1R#��(,TY�`��e�`�TdAEH�Km��Z2(������")�T�+m�X����6Օ��lm��H�"��(�ER�X��X�H�Z*U���2*�6�(��F�S)�F*3
UU�UUU1Uj�2��r��j�+H,�`� ��aD��T(�b�Kj�U�����J*����im�%eH���kR8�T���*���F��淟�̚�&K��Hޱ@^W���)��̒Mk��ݗ��7K�Y�Sr����FP@�Lٕ��)�
<m��Jptk�aq^3l��꩟<�{��jw�p�u�֮�rV:W���%C֝i��ɎR���Fgt5X����FZ7Ƒ\懕.�%.�N�r�
Y�@�'���#n'q�>]3���n���5�A��T�WG��ʱ�e����5c�os#q���o�и`)_�����\�U��ODΏ1^��R�����S���F���n�YA(�������.tғW%����`란�D�؅u>�t�م�
��o�<���@V?�y�mI�{{7ڷ�`�n���y��+���\UR��N����mE:����;f�,�[�Y	_dWM�I98ܶ:��j���Du�'���3'�ĭwF���v��M��*p�֮U�{٭(�03�ȡ����=��i�l��*�Lt�{L��R�C�][��-�uD;�'U���7 ӂq�5�Q��b�ۀXvn��4S,W����E�<���e�\�XNg	�W]���N%1cl؋����)��*Pz}�O�<�j��l^����V��R�KØ�kPE���o٘��6Ƌ�]�D�@�Gq�����n�Z��k��W/y[��I����[TM��tWR�o��95	X��JJ�{lK���5�IԮ�;���幰MV$�ۻ�狘��ѫ^bS`Z��wwmƒ�ꂚ5�i�R�<o�����W�"�eWPuZ@��/M�W�����5;�Ta㽹`������]xX#��L>Q���85�$�l������Y9V����̹ ��������ԯyY: �i��X��U���W��؅T�mw<�6�iGUh�;Q���{Z<�L�y��jڬzm�Ѳ��b�J�נ�{V8!��p����$����wi��z���OK��.��Y��j���pX3�9ruw�$�M�����ĪWY	� ���}$$j8�,G��$�-u;��s��ᜍ�b0���Z�rSPK�� �7��zk(
��=h�;-,HM��6�n}Y'Tź��c/r?>d��vm�� \&��܆k�Q��C"�N@�(;0����|5����!�U��n����C�\!��N��r��Xͱb��Ex	��s���~�7���.��v��'����|\a�5��h!XX�>ƴ�ss@��c�(2��z+Y�5�hv��1��8% i�����H���ݪsE��a�쬺���w2��:�!l>�Zl�)o)2�G϶=^� ���\ұ�	��x����s�p�)�+��Ưz�t��#*�z�Τu��Jc��nˡ+��s�]jk-��҃�I��ez����/��ԅ�4N�b�0b�l��ԙ�;���8۸w��d��n1{��]-_7Y��e��g�5�9U�Ş�=���:&������e��,z��9��f8EF�,_��W�a���De��?+�W�O����<�]��}�q��v�����ĳUd��"ٌF��b��'�)�z��@!��=g��w{;��S���!eole2���z��H�u��5z�U`5:ڰ0�<KR�H����;3�^]�/�p:������"��5R�4<�O����g>�>WD���x��U��*m�X��g��<�^͇:�΢ECsK�������GTn^MNs!���Ǽ����4A�X��bu;�
C�U�⮠�z:.�p�]We��/ܨ��D޻웅Ø�v��J�>2Q�u�rh1�0B�3Q��� D�1�x:���4X/DP$<�绗Y�i�DJkf�k��a�t�9�h��N�*0�*6�!�4�=���dLX�̸��Wb�s�o#�f�K��cg���(7�R�kI�=��+&2׫<���[[�*��6.�ȸI��VWZ�+��`����\���р�/�����#t��*|s*�B��#s�ө�� {mAV��t����SV���:DU2�;�lJE$��T�Mw�훈z���#Z�s�~���x�Q���f��"��cy]�U�Z��y��׎�����n+�Ss���>�Hu�Cb�@#� ��˙�b�������b�ܡ)���3j�ܡO��=J��N����6�W�3�)�&ի�mM�d�B�ΗiS�{+ �8��F��LZ�F��0�]<�ν^�j���C�bx�F_nG%��������?A��<}
=�N醙X�)��M�.1��>`B��;�ne4�%76d����HaV���1C�'i�F�jaj�0H���t��l�s��U���G{�cі�{^Q�h�F�3���t�30-���'Q�^;)�ee�/�����i�j�j��7UE868X��U-���a��3��7��0�ճ�FU��)���N�r���X���1�QW�x,�Wc2K�x�~n��X!w�󸛈���j������Yu�75�s�N���u�t/�� ��oD�i�c��!�S��y�ڼ��k��逍��ظ�[�a.�,�{��'j�Zr��싨_T���;�6��auAڶ��	[�b��^Ie���[��fD�u	"��6�:��&[�F��Z�����]ġ�D�i�iP�=�-4]4�[C���oL�|��I�j��9�A��zQ�Z�b�e���$�������0���x��>�bVE���_vk��vs��-����I�IR��3�gQ̉����g�a�
+u
*�׽E��J<��Y�r:x<�.c�ӻ]�s�i�#η]�̮�d�O���Q��C*ϡ���ұ�a�Y���􍆙R�Y7/0��נ��M�dd�ʡ�a��2�x82�.��;Ҫ�;F�v	�[�}VQ���m�>t�X�|���ͩ��^S8>��y)z]j��m�kJ̜��Փ�u��3+����<�ǥZW�\��Uī�z��6�^)A�״�T��4t�Z�"b�C��pj-*�X��Q�x��m�D!~���u<6K���H����kX��gO>�B� *����+��A�L�����u����p�Q���-�*0jkA\:J�!Q�r��U0+�/���8:Z��G���C]���E�j�h�Rr
����t����Лh�-o�74�mS�_�����X�E��MȂu�u�^���6����:���{�>��Zu�Ђ
�f�E���4a�~��Q��E�s'�4��ow�ma�{T�u��O��s���u����3q@��]% �Ư,��Z}ɩ��F@`�H���;%*�I٦3n���nn�.��7h�S��TX[�*�7M���ЬTX��N�Q�mS7��1Tܰ\��w�4�V�
8��J\Û5}�#��C*[7�4,�U��{|-���C��SA_��`��e�n�6�i����8l����Da������6*;�e���E2�y7ku��'**��Z����s��k��q%W	�w[���Ƨ̟f@-�l��Q6�9�)wbv2��R�����=��B�c�ftZ9s�<��:ch�[n���a@8��u�u��vm��x����[&*�r"�!$�b{<�C���Ņ��a�|tg(���H]P�P�f�پjк�&��.RA����x��^�tJR���ub��������33��jw;���4�/ ������Q�$hz�jܡ��sM4�:w�%�eQ#EM�0�Z�d�ƽ���c�9���[Ta�b�N#�.�/+8Jk��U�e&�R��|��ș&�iޕ�Kc�3(;��#Ta���"HBcL��_�����B�q�bP�.�b�|.f��b�e�]B0.Q�S;�ⷹ�_�9$� mV�ydQ���-v��s��Z+pu���^��fg9Í��n�"��&�z���w[��"�̏(4w�aƪG�<���1��:[X;��<�L*��Y�6� �K&Ȇ���y���=�5`�Z^�x�â�V�W�ӎ�{�Bf��#{��	7�\��ͷ'�ۥ��]@�^n@˶k�Q�oO��WA������y�Z���%�,c�)e�[�|��q����|���醙n9�F����+/�JAW-��]��:~��;�]t�֒P�q�9!]���8[�����E#!@��A\C=�c&UtM-Y͜�������щ�Qt��dB�Bh�N���J�p�)�CnH�V��6:KX�j���J�@�}k�즘�e2��?)W��3�8+�W}��̿J���}-ϴ-�8��u��N�D%VQSio`j�(�U8�j.��Bb�C)������3�SXU9��b�����i�@��K�g�,��j��T����&پ�C,*��4b<7��*�u��N	G{{����M$����ܵq��t'0��~l���s���4g^>=���u�(�8�HH&R���Y�ȚO��-�c�����Aϑ53tn�31³_�!MR�!�E��t��Qmҳ������y�G�S�2X�ĮZ���bA˪rz��ӊ'�S�E�w!eb�:�"���eÅ��v��آ�VM"�KA僷g��w/[�γ��nonLZr��]]p���~�.�Ŵ�ͣ[��vz�@�!O��3f�,]�����[ʚ��̫~_<���ي�!�X���ѝ5�e��KR����*M��s-\@��*�.|���/;�I�qu���J=�g����z�a��žҽڇ-y�by�L:����TW���\�4�?rs�iL��xvxiDg�y)|Q=¯W��[eG�㝅>�Z[�G���g�g�?r�-���z��Pj*��O��|Fw���ʂ�M����r.+��.�O�f�*�./�_vJ�P���	�%�oSUеH״�\��:]E��s"�ͫ8���RWC����~2-+��)��vu�M������f�w8�Zۻ�t��e���9�5	S9g�m����{�y�N�|wѯw�rˤ�B���+�[�T��G^��Sk��N�<��t;�M���ܠ�$4��)��ǁ4��N3;k+A�(�ޭҾz�u^j1ܹ�Ƶ�x��q婪�q��)K$V*~�s�u��%�y����$��[^|�י���/\vJ5�O�sI�z�8��u��D����<v!tY���}{^k±qy]���7Gr�G�瑎�Tj�Н��~Q���e����yӽ��K�o��Ss��C�nb�j=��k1�ځ)�.�u����{ne�p���;��~z��Ni���.��f2Sң"7�O)��P�	z�:�rUt���kk6����z��ypg^���E۴�m(8�AyH\#0�Z���+窊���;�fs�X�p06lں��f{$�S�粺a��*��ƻ��V�Tl����
�����C]������(�����{���.���>]�!kq��Ք6z�9�SMu����@��.��q�/̽�\F�r��N/���L�An�k|���K���[��b���}\�']W{ļ��l#Y
H3���0Auz&tzet�Ef>9�n%���۽n�1�7�d��喟j��I-37�o}�61)U64�Jj��E�g��Lz`QH3���W��MVt�[��F�&�W+We�E�4�A+W<2S���-j�;I�Ӹ�S1�͉:�U�>���y�T��f�Ŕw�d�x���}�bV��M)(���|z��GnDOK���joGK�R����Vv�"Mə��C'-Ǟ�I��o��/�W���|��-S����';�프R���Mߣ��|�%��G����lZٛjyZ:�p��y<�z�,�kZP�<�U���z��������+-���M����{��Q�-{��k�^�r��������j��zoS{���J5)4��Ec�'';�k[}���*�Eҟ�����RK(����y�7��D�Ys�:�Z�%�z0k�8����1{7"�Hn�ħMS���m��'bkD�ކ�帀�׃����UFr��շ��@�Oot��Tx��!�̭��'h�1Tw*�&�"5�:��]��{�	�U����q_���}��3&�v4DF��®���7fK=�,F�7�Ti��}�t^+��f܌;GVI�Vv��[�M����6�nX�OM�B�M��2n��ۣ e>����Ö���b�(=�u5*9�b��N����4]�-�Ma��b����/t�,��,FI�nV�L�,�;���Ɏ�Ո��:�\�ԅ�M��׌]�w3�
{����N&��Yef_2�k�bF�33;�O	Z芲�XS^"]X��B��ɒ;3;Ev�b��RzЦ�m���[yw)�23�C���fK���s>�����M<Se�ʿ��hQ*���[��T��svX�ڔD����ub� `�Y��	wؗvK��s�E':(oQ��O6�V0jƍ�yc���-�p.x���M�D򲱗ʮ���GMCΠBf�\�>��L�anB,�{f-�X�t�x��1XK0gAR5ї�kxs�(�Ӑ��zD|�7�Yѐ��	���\M	�-hm�&S,7�L[]���h�}����r����0SѽII�U�2,$x�<A�+����`T{`�#���"��Uzo�,u`9�WzU�]u��K��-Fe[�+���6�cK֍:��`[�{uf��v/\=�������C�՜������Im\����J�a�\�T#D���8��a�3�ϩޅ�R�Ӯ׵{���\S�q�s�Y%u��{>�<�M�L���ۏ�I���ef��!۰f�	��W1@�����'����x���8롙¡��(nt?7Z�HT�u�����Z�ю[���D̷����:�,	:Ɲ}�5%eI3R�g)͋���e��VED��ּ�۾���yBH����{�+��={�|]"���P'/�Mx�໭i�RZ=|��t{���Qe>s�tc�QmƝ���e�v��ܲW�˄�ۺ�ř³*Z��aWAs���k,whX���r���ۼ�utvMh�8�5*�P�6�V>ȅ ��ؾig7wH�(Q���{��IWX/SI>�����-� �ݎ�8� �fӄ��2dF�]�7:�s.Ix���p;y,�yDb/!P�Q�w^��*c��k��vH����t���r�O��K�k��r�вS+�egw���mo��D���\M\D�%d]v��{���t���y�+��Ui$������}J�1.Ѕs�����KA��n�5֛���nǋkiq�jh�.�1.����𻝅�h���^�\u{�v�[ɲ�r�TȄj�)h�7s��r�+�N���Ma��rC�2֜Rf��r�lk��lb�q�ň�g�8�)ip�z�
&�N��ޮy��NTʼ���a�wHK�jKyoj	�0��n�gXG`Lm�a�2X���V��4� �;�:��t+��JS��Q�WO#9�L�8���+�\ʒ�y���uK�w9ߺ��,F�U���t�:���PA�8���+#�ޫh��^������H�Ř4��"U��[���֭V
���L=3�z�Lh�]<�r���x�*�v�i�s.-C/�t��8�ͭ�ŽN�Q|�-j���)��pEAD�D��[�+QQ�J[,b�m�bR���PEP�[l�m����AV(�mE���ⲲT�	e�VT�ciJZ��D[nZ�6��DF)UV�*�R�h��r�jڪ��k[UX��b(��`,�r�(#ZR�QU��Kkd˘R"[%Ee�
�ZE��QDcJ(QjЬ��YAZ�Z*Yk�*����G�\qp���X�R�E`�mh�����Z��3)[Jŉ����c-����h,U-�+J�U�\�[r�Qs.-��U��X�e�AX��Ub�)EchW4Q�EG.`�j2��im�j£J*�6)QD��֪�1lS����P��bQVլJ�h�mE�ԥ�H��+V�ԭ̳1�֫�m���-�T@U~�{Av�'$��í����|DL,��Lys��M��j1��u &��e���3N<�:�սR����o=�}=S1D�i��|�*��|TN�
�l}��\�s��j���g��"�V��{I�7{mX��w+�9m=�8��G�9³]{sj�eax�n͂�gse��h�V�y��Z�~Y�7(�5�<�W�͚�3�p}f:+r5���IM.6s���:�:ݮ�������>똵=�F��9͙%u��n�J�eZ�.=Ӛ&j��Y�՝j-hض��>��:��c̳���gS�uP�����M�]C;Ur�Ѡl��ǧ8�﷗rH/w�Fݸ�S�O�WT6���9�j��~g+9ԱR!��>y�~\�?>������#��� �Q�9�:4w)�^�b��a�tf*ȼ�z���7������v�MZu滝�3ʣ���u]�ә���v�;�����}X���Yp�����鷪�N�x�֡�+`��]��8q���0\Ԙ'L���$�o ګ���o4�W��w���5���x�i�mcҲ�g��3����g�<��'Q�*�����OS|ތ�:��Xˏ(��Q�xњ�,�S9��]�u�7uƺ`��t�蓇q����I����k�Q]�}����n7S7����6�u��-I�|��[~SXU�9��1x�׆-=�W޾�����T�×k����q������K�A���k��nUI�h�Z����[�c]�]��%Mg4���V����i�p��
GS3�γ[�U0��JuE[9�{gq�������Z�,][�m�軔����]��4�8e#�Kq	�(��7G�8;�f��Kp��Lu�u6a���"�]Nr8�+ #�fJ�a,��^X[q ��B#�d�I�e*����p��P�o�8�{zH�Ou6�r�W����t(e,���ey�#kڬ�ֺ0�8�m�n���]�c�2w_�ʕj�3���W�qxD�r��˅z�ǵq���j���o���9�}M>ڙ9���W�k��ɏ{E̯o�ؘ��Aݪ�J���=}G�e*em���P��v]�Y�Cz"J��R��K<ܝ�$Ɩ,���]Թ^b�V��8�E12N���=fUw1{�Ҏi�U�>uw�#e�g�X�F
��Σĸ֞3�eZw��U��K�t+)tj��2�ޑp19�m5Q˕N��J�[}��q�]x�֬�W6�o��N4�:;p�K���>��_.���mjY<Σ���Ϻ�]Ԓ�G�r�&m+����LOoU��p�L��̲Y4�S]�<�u��q�E��a4X1��m,���ջ2��ߟ�z,M�;�7ݶ�\֍N���y��v�U�-%�1cml�*�j���� #qIsݓ�-F�Im�r��Z�+v�T��[܇x�B�Y�zB-�Hm�䞋Qy"�p��[׫r���r�	�{�����\�uٴ4��\5�.}��*�Ǧ-:��Yx��N�(�I˯A�pP�fiy�դ���ӯb9���'��W��+�}��b�UNW�,�¢:�h�9y�޾��g�n��:�gߌ�ۉ���ۘ���҂����`�y/&;:�������w�5���LS�wH�k�c��C��K>qK����W��0d����U�S��uv0�Y
�LL�8ψל����ޤ�	q�{#��Ҷ������� \�J:�28E�8���,d�dr�:�Ju˧w��{ѯTe���Jj>u�k�X�`�fͫ#��h;=31����};��I���
\�����CVS9��db�8U��Ìb�]�6+'�t�;��ݳP9��Z�gձ�^�r���v&�\��D����0=�Ik]������2V>����T�d)y��kx�ݪ�'�j]I\�ުg��spN��)�W�y�/[n�MM��]���0��Κ̼��ˆz�U�
���!��N�o^�Щ��)�b���nX�oW�o��5:3�UP�B��J���7t;�Ƶ7Ӌ/+!�Ժ;9�=��ܮ8�Ƭ�6��y��[3mH�;���-�5�~������lRw�I�9�.��\F+0�*8�Hsn.�]�Ngp{��ݩ�>������c����W��up�O���!�Aaֶ��m��r���GuL({o<��X3NW���;Fa6׽2^R�6��m���T&��'SWwr^���܅:�/�-�ᖬ�L��S��������:��[��y`��Mb�%	�6O9c���=�/��\�S)���4&#���S[���U��$�QooT1SHn�����v7�j�f-�)�,*�9Ƽ�q�ˋ1U̹{�
r�˨Ì�^�[��e$yJK��u��1�c��g����T�w��$�䲃y�d�엘���TJP�.u��j݅#��3�k�u�WנA&R*�̚�oY	m�q��c����s�nl�T5�<��!)c�vWe�=��{5��9����i�=�~{�1𪓍�G�6��ӕ�x6�4���N����>�Y���:TvrS���jmF�@�U��kuùc����w|:'9�$�bp�B�hZΥ_/v؇�b�S�3;�w)'iK��ݸ�k�扚��,�m��:�U�m.��u9gla�{=�R\�n]]>Ԋ�����1i�΅]����s�\ox�T��o�roo�m�v��(Tw�+��ұ����g�q��:�j���� ��)t|s�m���-a���{P
�ˍ^溑����6.:%�����Nޙ��u/lP)`}ѷ����a;��}-��`sԺz[��gG��8D׽%*�o`V+(�f&3�г���0�5�_���v�Z�W_M���V��H}��*[�>���]M��rb5�<10c��.��h\L�J���k�u=Ww(�ݏ�,��k�x/U�pbEI��}j��[����iu���ҫ|��:o��ˣ��Y���9�(�$���TҒ_y�ñ�͹���}7�;�V���kNJ�ӸZ{L��S���4��V����z􄠭Q��}�Ϫ��@�q��]}����N+�O,���[~SG���U�k��+�O}c(�B���#�SėGu�������w��}pi������y�ŉ�\�Bߟ(�tsz��dN��^�ε����3���.�)��:%�����u��g�^�$�����S�4�=9�*�)9���b;U�%XR.�o��r�tց�^gb�+��>=짝CSsn��Qg�&L�WK��}�}�*L��x�����vJ�׹,�"}�4V�|b�%�c�P��05<0] QXE�������R�M~�-y�Ox"[:^�ķQ�mQW����c�:G��k���x\��pm�y��ٓ��+�3Y"�v�5���vj[��׆i�c1�y���W��c]��t��Tb��5���6�d���n��n��͸no6�����T�5yf^elmH+wm�6Z�h�.���U�jqZ��y�R�+�)y��mC|6힥�k���ۭ��F���+�����V�>I���USm$�o�<�D�TL���3V�i4�d����0�B���q�&/�����9qױVNJ4��څW��n�ie�qՌ��p\��󙴯�=7.�ݽR��E{�ݞ����XWϟ5]�-��|/o�Z5XqÖ�n*��j�U�㪎�VOU���f����Z磓O��}jDKIE3�X�F���'���_gs�~;�5-�ۯuk����܇q�GmS+����;�B%t�b����!���`����j�����܋�ε�Ot�7쫚Rz�?>�ܮ�A\]�Ӡ�t���²��Q��>৏Wj��Y����P<�QotX��U���N�4�z�̆ϓ(Ӛc�@�Bf������2_��+�u��ۼᒸM8��Y����a��r뢛�ݑ+✤���w�f�s+�sč#�s��1m�F]�ns��K�',��[�^��늉��)t�/�d*����A��f���Xf#)�
/�d�+;����{�90lQ:�vzP����x߲U���r?��L��P�ҺRh�M���.�"}c��x[�3�Սw ����F�ק�Ј���ٙC7�ȡ��\�uN�/����sQ.a���={4g=X=Q�sC�[�|pf�hw,J_i'�<�@��U���.�O��c�l�4;Q��<�\��rb�L�q�6n��ù�O'霛{c�5o*ع�ی�;/
|;�n�uw���5Z����ݧ�%LN��9{�>�qv��i���!�rwp�U#ʠ�¨��i���}n]���	o��V%]l�~��~��a<�<���cJ�bh�$T.j���٫L����c鎂͵^x��v�����X���q�b����ONc��Χ���d���Of�v��حd����k� y�VNX�����v�eZ[Sq;�]��{u���}�M3'.!�ՊR��o��m���p�S}�i\��n@Lr8D��^�ԒP��v󫥵仕�}Q���J�D��kb����d#Y�qE�4��mN?ZU��^�v�%p�L[Av*�m��t�Y�=3
�z[ǡ=�Z��5��o��]
��;3��{~�~�z���K3G��6v��H��=VnI����0Sځ��5��B]s��Q��]�J���/Z����2�Ts�ǆ�#z]s��J�)P��.��"︬�}�lV[c�VO4��u����k���諩���M�0cCr(x�&gq��X�����}�	�s��VK�\��g]�0n�A�2Q��bs��Y�ݬL�W����q����}�Ksg"����Euhu��Y��X7#���IAl�u'���S{Q��ϣQ��b�>y���gg�}W^�,���S�;����I�'b.r�o;�:t-�Wx5e�N�]8l7i0ٺ7,�9Ec�-wA�w�vF�ST,�<����!��0��}�®��/���a�� �Y�]'�O�\�'L�1�w���,"\�'-	J�@�5L��s�%�)�N޿2;*+���N�T٩�MS�qs:3.�m�5ƥv�W��b���C6�'bmx7�	��U�z��/q��V��ނ=t���� �ٕ�u�Y���N5k�r�[�;4�#�*�5�E��@�&b�6�^�Ew���R��+k����:����p��^�epD"3��-�:ԔV?n!0��+�@�_=�M}���|�V��H̅�=\�l�����.�⣜�SiL_r��z��V9�Dc��<���ri��j��*��c��E͞�{�*vڜ�|�57��3�
�=�R�+q�6zJ�����a��:ճ�e�[�1�����=X��M��<6�')l�s-4�c�ưť��yٴc�(����m��^��g��F�q��[���Yn�~R�/W��+�|k�ls=������*g�Y#;�
庫��b�V2V+���Ӡ��G�RˎN�5��n���<���"w@�P
]n��TQ^M���U�c����N�̆�w١�����N�.�)tf�z������w.-�o	Ό6$X�V[[מ:�N5���/}n���Ƙk#�"�\3v����攭N��{����F!F�8W6B�i�7�[�cRc$�&�Jv��K�W2
۠�p��d,�l�m�� �zö��e!��ҋ����v�`p��'<�*WJܡ���mum�*s���K��n^�N枸�x�{y�Kmgj�����\l*��a���{
�	KN]��E��e����˕�&t�L�QrJ[}e��R���n�KoGT���#KT�~�!�9�d[ڭvIA)9�vm�p	�D��t��isGn`ޫ�y�����k,D�m=F�&���(��]Ӹ���L}��� �Ƽ�,�l'AO�G�T�)�g`��5��v�������z��`�kMvV#3�"��$i���ە�j�-�����N�}wWf4���SbfV��Od�B#9�wz�0wo
H7CG�l<7x����r7ە�+��fh�1�cʸs�m�J�	��kG�8u7�}6����.�0�es�t�W�*�c�7ң��R��v��1�h[�&�홟^�y���E�I��i��rbk-_�QE
/�ݵ�݋�=5Y(A΢];2�W��3BV�w�c�.)Y([�8cv��v+7WEW 94l ���k.Ӱl��AMa�x����ݠVف�oV�zť���ǆ�>�{���{��s�]��M�yJ4<�Wu��-��+���W�os�����9�}$��)�U��6���)�3\��
���v�+Y�b�G%!Q�׮ͼ\�rx�w��][o��G��B�����9�6�r�� 9X3��-or��33'eo�z�����]Q`��S�xX]K2p�?
qf�X�5��^����Ju�x�`�Z7pC.ͭN���V���<�ҽ\z�:��!��`H.�s)CRv�;�j�-t��X�t�j��S2�NЕ^9ݶ�*a݌Xw5á�`|>b�H��Vh螋���k,e܂�'���).�J�*ҕ7�pX��lPj(Ж2�Y׀�}��rL*�r��Z�[f�`ύhC{&�eЈ��k�![B�h3�ٲ����l���Ig���w����c�tQ$q�|7�t��v��p��C"�J'&Hۇ2J���/ f�5�V��JXX�
U�`�3i�V�� +�������9X-���FqvF(�->\��Pa䫖�4 x�dOSG���[���`{���:r��U:��Uچ�Sk�Z(�xP�Q�U�D#Ju������'��mhta޶.͡ƒ4ݴ�K��`�rL6M���U1^:mvdGl|�p,Yf�CM�3 h� �EQ���{K2ت(#kmJ!U��E�,QE�Q��-j\�jVT+m��DKj���U�R�ʕ*K�1R�KVV�j�[`ѕ�ՋJ*5F��*cj%��ږԱFZZ�0rcj��Ɩ-�kj*���[r��¨��lT˖��Y�K[X)iE�� &5q-��k)aX�m�j%�QjZ)TJ�6�UcbUZ��T*V1�m���T[�.s�ie�m�d�V�hT�Q�[[jڥZ�k
�QT+�Z��F�ыkTVR�)q��[�Ҕ��h�QD�UAm���(�J�"�)`����mD(����խ�ҋL��[h �J-R�յ��V�cr�KTkm���[Qj���,b�j��,�F-s0�*�KJ��mmqɅT���KZ�hҩ)jڮ`�q��Q�3��G���c�u=��XL��p�Vq��-.zj���Ț�E4���bޫ�R�魢�"2G#[�#���4��z��ruN%�W?|{�ޝ��{}��Ĺu���jGS�`ק]+N-��#*�i]��^�j�#-ٸ��lK��n�:מ��#�qq�w=�.�Z�{|�g���4gV_����d3V������cz�>�5�3	�g��� �y��z�\��5c&�:�4��.F��=���b꘰�%��6lތǚ��b���~|�lp���O��{��õAq�^�4���!r4�D�e:l�w��Ъ������^\�_U��yc���df׶B��N�1��xaU�M�W4�!k����0��?};��)��9y�U˳�N�sx��Ō|���7mr�T�n�*/����<�f�7����k�ѵ9���-�\]]S���Y�B��^]]��v6����m���WS�Cm�-�ڳxQ��yS�k����B��m��}+�P{
�z]�6�uԹ_��PTnOn�UU��F+:��
WaW�v��a�AW3��T�ù[�7�uZk6NWM�|ACK4�i*֗mQ��L�r2.M�}�X���C���k6�a�6TV`������Cz�2%yq�e����<���Y�oz<lXdK5fr��we;0��V��|�Ă�E�g6�Stäxb�Y��s6��OL\�v�ۯށgB��)Z��ǭd��t����9�e>*������z����+ԩtt�-��f���=�U{��;��|�7�YY�9��;��D�n�2Z�D�	�:{�v/n������Ѿ&������w�B�YA@���b�KҋH�Ko�</:��^3�S��[����j"Su��ୗB�EGl�Z���>K� l1j	������@�U�kW��C�bʣEgB8(����ܷ���m2�eR9�}'=貱t����H]Y�������疾��%y�,��aͯv��äj�4i��u�zj�_�1�M4�����[�d��K���7��^O�u�{��mP*�x���@�ɍ��bܼo�.R�qv�n=.qx��Q��=�3��6׃r{�vصR���f*��C�/��x�w�c[�r&1������:�W�NZ:��N(�����Ѳ�GL�.�tygq�C9<X�`�x��Gu�$�=��Q����Z�#7��⮰^�>�㆝o\�}gI���6O�f���m�d��E၉RInѦ�����=�����}^g+�S{i���ד6r'�����Y�F{��E��·ܻ�6�<�M�3C9mbޢ���5�s�9JҬ�	�n��w���n����B���+4�Q��j&����{�7N&l��D.�y7�k����0��G�o�3z+�-^s�qu�k��f�O0��m����V���޼f���|�˪�z��K��mOVl�r���'�Q;�V��)�V�WOU�.�q��F43���!)@�r��5�l����s��NE㉛j�\޺�ˢ�S�;�h4�5F+1pʘ��q��2j�2�;W[Gò������WL\���+1e��;�VAqZ�Nu�C]���s�m�;�"�	��77LV*��0_m@�U�܅��#�r�^�|�-�j\�u@]�<�v߯�ՁA�g��E��B�y�wq.I�-jc����
�c:L��� �:�ͭ��-U�T��eYJ9|��wز��M�6�RZ�cRC$�Eޙ��z�r(�A��w�n*�Bk}���E(����f>|�76U�]}̘3t�"�t��h}y����� �v���D�Lĳq�^��o)Yj�7�L�o3�BVCj��	Պ�N�;v�R�Ֆ�%m5��%ˠ��#rC��u�9��0c/�:��w:'������a��ͱ*7���s���l�ׄ���f�ǜ�ٌ���[;���"���ڸ��Ǉe���q^�\Է6^�CZ���f7	�"����W�5݇#��P��7ܒ���םA���������fu�q��ԃO`\w�[�)ojuB��zK��f��s�⻌sۏ����0f�;|߼-=�,�UG���WKt2qβ���r��Ջ>j�!Kݸ��6m��uk9�K�����[E 3��j{����)��:��J��)��̶�e�z��WU�eE9@�"���i�6&)0�ҹP���{�[��k�G�OZL$�ʖ"�
��\�+��a3�)
Y˩򰻕�s�����?X1#�<Ify�,�����!�xx�䅛Y�;BV�7=�{*6R�v�6��n�ugV��˷%k$�}���׼,�R�O�y��d�U�c���cxc��)no<�M�/ٴ⸵^�z1\ͥ'�-���ʻ/S�i>�67(�������[�yR��W�¯2Ê�<�F�~���&�Lj��צ�"��+Mr���.C��ԫ���u�My�U�F;�;Z��|���WYEv�-�vݓ�Z�Vk$�%�Lꍼ�ie��C�c�,*�9�J��-]�,f��Užpw
�>t�/�盿:���ǥ˨�
nB��1��-�GI��]{&���<�=CŊ��T������[\�\	��ƻ��ed���|�����k�M������<�ʼ(�;���Գk�ذ�8�ۮ�z�OqȔ�g!H���g^^�{9+/&b�3���P�u�7�n�,'ۨ({�b�Rٯ=��O���~��ׅáq�.���r��;�D[y��RW7+RJ;��F�F�u����m��3P���7w̌�:�UWY�}䎊�^>����z�����p�m̵��n+��鼇>5b�x.r�Ѹ��a�4ὧ���Nr��7t.�Rqh�fe���C3JŹ�,�����b��F�krp�u.���j������Q��3,�K�����r��ܼB�A�34
���Ԭȵtǯ]�����5����ܶw�+�e���0���'�搟���˚�&S*����]݃S�U���P����V¾BӼ��%�9�v��J<V������U�o���Iމ�k��P:�m�1֭o��ж�G4��V8��5���3�t!���׭+=�9�;s�Vg�Y��O=���*i��7��p��+⪡��D�[S��wk˘�<�Tk�k���e7���v�v5g��Z�W6�ج�U0t6��4Oڏ�N�����zQo�j�d��N�~w�q�m��q�:�-�ʭ��a�.�n�0��ΟyӒsU��s�o��P�1��S3{�Xl���u�&�l%�1)ƕ���3���*ۀ���O{�2T�T�>�$̛�6Q��1�U6X'T��}�#2�eO`'Ւ툫N^�m`��%;�~��mnQCod�e���q��b���@R^�
�WՎ���U��}35�9`ɼ���fF�娔��E�,ھ��"�6�̕x3zAEU�֌��$�R���wۡM��D�lt�x�*>��{�G���Z����*Y	ޚ�L����A~��nP��j�Ǟʤs���qO����W#�ի�X�N��2w*P��^��ũ�s��jҁZ�r�r�9�6�M�B*����Mu�Ė�]x\utn7�=�j��3����b��W��Ʃ��m�r���d�]��.qy	<��C��-P:c���Ȕ��-�ѯ�=��8����_��T^��quE�&V�D��s�;N�����F
Y�"u�R٬���K�#�^f�Aw����y�{��)k+��y�Lɔ#R'�I�;��썵9����;��m���u����I!α��MaN���l�>�]=5�{�>�J�L:���ӕ��O��\�j����)-���*ŊrB����r���Z��}��X���Ux����9R��!�R�\e{:5˦._OM�v�uS�~ܮ8��Ɔu�v�)�>��&lA1�'��Hgi�&�ԩI�Ֆ�2����Pn_1�c9G��:sY�Ղs���<Feܦ0���^�t:���Öx`ޝ�a6s#�X�ym��j�ݪwi�Ǽ2̰l�ܵ�o�B���K�]�%�L� �j��7Ԑ�[}���re��c�������]�G�W)Jmfoq�y�}�o���up\�j���8�R;4�S�QiI7�F�B�_9�ng��Un�޽Ֆ��Ι,�
j���ج���v\kѪ�؅a���#�oK���:�v�<L�� ѹ��/�k���}������
��p�|�R���eaYW��n�<�;�����\�˩Թt@U:F��lI�j嫔�m�\t������kb/'�8��f �|�X�Ϝ�4ͽl���p'���m��=�N2���5������;.;{	�nx���n��RO�X���J�Z��F��i�\�]�ފ����v����{_܉��QhK�S�2����c]�d��MT��$t@��]�]�.�6{9cD��s����6��ܗ�NJ�v&׆�23h뺜���v�\AY��g!D��,��:lU�{�lRչ�.���Œ��yz�/\�S��T�>���2��&ViaV��i\��s3:�����s�<'I�b���r�J*	L�����9�g�Fe53�� ���U����"N��k�V���f6oXwN�d���o^��A���<��W7v��ߛ��{��ɜ��/lM�-����3n�i��;X�_%�<ޥ]Ӈ�n�u><���k4�]��{��S�U�3q%(�ᐓU�iU���b���_ݮmٲ6��ۓ�g��Aiog���n��RBb֮�˂�W9�O����I��[�on8�X�CT���JY�s6����[uk�]b|xS��T�e��%nQ�x�,�6��S��V�9a�B�Z�j�j:�2k�\Q���)��}ϝ@���?x�)��{��:4��:�^�18���`)�y���zzV/|����ڬ�ս�u���Q'8(��<��4�y�{F�+�MR���U^�t;����r�쫊��n\���Ȇ��~^��P��1��j�^�oc#]����	N�E:�w�zOy�y��;;g!��KNN�Z������K=�w�kO.i��eC���[��Uxڬ�����D���z�c4:k�w9�7y���c GEmh��yK�I汋b���x����0�:��H*�]��d�Z�LuXV�c� ���x{(�<ޜD�7�c{�	�}W�7C)8�w<Op����9��C��&�e�C>��c)����/��>Ir��u��&�nM�l�[�j�g��{:�j�j�`�{�>�׶�?M���^���9���C�T�l��7���U�ho�q ��b��%�Eh#0�ذ��~�S���t���f��3O,��wi�����'H���(�M���՟D�޸��vK�w���|���p����9�y��q��|��+\Z��u��x�wi޿-�t�}޼�b�R���)r�5���R~��A7k��~���9Y[8;mtʠ*t+^FfSw�z�ܾ�w��$��.��Q���=K����'�׭!|��t�du�WA�j��M�X�����cWSi�Y�x򼧂ێ�T�F+����=�1b��n�٤�J����I��|7v#�ݳJXq�dZ�\*��D�X���=+�y~c;N
m�
�<�����ðZKw0�C�'��N��y�v�M��u�ZCV��i[���LN�|�`�6���-_WH��V���^ń{"�:s\�
w$����<���b�3��og�K'N�s�E@��me]:Xph����k'd��vzHTr�rV�1��3Y�ql�� �� chu��oy�Y�f5�T}��ʊ�*w��V&��+���L�~��0�r���_:�c [��cTj�D�}Ƕ򏤷F��S����)]�=
$�GN�[�pfrb��e���9|�J�����ƗB���IF���&��
1׍$��"����8z_;�wG-+�mL�+B��M[��>�|Eo7,S�Ʊ:X 2-�B�/���X#g����X���(�m�{��;��D�t�u2�"�6x)���p��+3��LY���{�&m�؈Y��p���`���@��z�SUqWk���r���R�,ۧ��R(5W ���\s �w[��|�:��c��Lj����H5C8�._�5�9���P���E�'�v��i��{�q���{rc���H6	��v����h��p��K�K�o;l
,T��5}�|^O%8��X��.��ͯ.��]:U�b	`C2�2g�z�&������tJ�b�)�t�}8��cT�r-U�e�T���G��!��I[F�^
��W���Iu�Ӕ��� ��y	;z���ܰގ��8�3U"Wl��BC��2HE�Y�;Ha�{"�ͪ=#X��]*�ݧ[���rڿ�cg"(Rǩ�H]uK(ǋ1V��_g4�Ȭ�4H����͸/h��[mq-�X� ��nT�T�m���$P���nXp����P�r�:���w�L�|��=m��.�D�VWkX��h�Eu�h��݋;�L��BD�]>��C]�rIo>��.xe�Ǽ�M㷒�نB/���ḩn�l���l���A�NXf/��w�6��������t�vu$�f�ix��g���J��Ib=�)f��y��	/�V���Ƴ=Ũ�!�²Db;5jvSe���ʅ��Y���a��si�G>�QM��>U�=3��5������<?>�S����v��k���T��H��w��7���FOl�������c=k�ZQe#�W��ŗ��5h�5M�ˏ��ඝs<	+��c(�j�
Qt.�Yz���(��ک�J�yaT�m�Ƣ-<��Q�ۦ�N���_� �t��F�ָ��_@��r�Vzα�B�u��֙/ql]^QLV��2|���IU�_�/%�(,�1���]gr��]�0]Jl�Z.=�7)��:f�[`f���K1Y�O0�Z#"N�t�--�r�iDE����Ѣ)PiU���Q�5mjU�bĭKZ�J2���DV��m�P��Z��ƍ��)Z�J�Lp�Q��mQj�J6�+�Dc+(�"��,�ij��ƴJ�m�*��,�T�E��V�k-
T�j[h�m)�X+��ѥV�F6���ڢ̷V�ĭQ%��R�h-d�ZT(�kZᔘ�iik�m�km+U*��r֔*�cklm�%��h�V�"ڃeB�*��F��b��U�+m�eh-j�ŬeT��m��"(�*"#iF+m����V��
Q�F�ը����Tj�F��l���U�
#(�m(*��(���R���Ke�FU�֥U��)F�F"�ickJ��֋m���*6�Kh���صh�U�֋R���R�rʒ���3��n��j����r�%�]��Y�[o6�=M�6+gZ��r�]�=ZC$1fVm>}ي�Ւ�+�q_3;V7����(wn�|[�(w�5	�ע��,1M���x�\��5�_�fߦo��[��Ֆ�'W�-�CF.��v�a[�}[�.JȌ~Ã��!Qw�b�TeF'�������c��0ʝ��vB��#�����tE��j'UW�n;���Q쌵y���uH-��}A���#̂�"y�r��H��{�/�t��z}���JC�;pa!�rd�4҉���P������8�̷�b*�^D?6�Nx뢫�����Bg�y���m(8�g����y����Y�����ɀ��{�q�7�촢B�[����ʟZyQ��O�<�N��ᛊ5&\sڇt�oo�K5�E�AJ/gz��˨�
�2S�^Ҭ1_V���{����N1z���	o��]��~�Г�b��w�����o���r'��t���[�w�_s�w/Y!X� {JBT,�����Y��SZ�3���"x5��+����Q(*;�vҔ݀�gi���;���;q��m��P�;�kq��|_.7�S�@���t�����h�q߅lGQn�fʝ1J`�w�s���>S�y��3���8<�W����F���;��6�&��˵�/4�&��N6ۭ�<������m��{\gX����8v���1�X嵉�.������*�\�K}y&�_:AT#���1�(���J���MyI�:�Ĳ�)Sr��]T�\�\[�z��fj�+�NgF���ŝڑ���e�-b1�JOt^*����S^w���c� u�ͺt^�j�q���&#�*8��qM��U^�n�u^�Ⱦ��V#������-K�ƞ�}��*�(*�y��;��d^+�d��υ�ќ��>��یž��Ǭk���"�j"Su���6��*�$�u��b���hX&x]-��y}��u魱��]5�^Pq�E�I�nQ;3U5��ޞR�/���q5x�'cg���������s�����ʛ�=Rl�"lC���_n5*#��-ʛ�n�2�F��]��<��K�c���k%UC��Mi��$마;G���pٰ�=yL��������)���Dc $��u@����V�-�{j�W]��ہ���Q_vʳA�)�ѰX�ոH��%�����R���n� �:��Eؗ��6�`�c}�uNx�p6����.ft���9�����R�|���s^�q1������I��Ngge��P�ը�P�=��V���W�]�U'y�΢��&<���=8�ݹ�����͔��g�9��t�|��o�.�Xt
�z�/o�7V�cr�+����');���^M<����󎻯NR�2ڸ��6󮩤�!k���ҩ5[���w�/x�u1Y�i@�[������L��Ǿ�l|��^o�d����ڙ�s9��~�mWoI��K�t�mY�� O��7z'�4�g����Ԓr��A�qq�/�������z�;^0M��!	��U:�@��QO��ܣx���К"榞�}�J����u��P1��K=�&m+�OM�U�\��èS��5��̛Ȯ�j�9<�W&ܧ�/���7�!�ml͵u\�K�4�ٲrq�M^��A�8�c��١��S��&�Z2��u���ڵ�(�ై2鸬��b���j�^g�����^�B�^�pB�v�Ö����۸����-]�A`� ���u���V��k��o>U�z1��C;�UJ�k�{�'�������1=�kf
[^�Gn�U�;�O�]��6�M�ѥ$ɋJ2����q��o�z����@��վ,���e��\���_s�CjY�������7�ȶi;��Xg͂�(��(��B+�rf�4S�����W��5q��]��C6��RsJ5�r��(��x.+�W��G��������¯èj�g��{�{^�X�"2o2��z:�T��4^��u��Z��B}�mW=C6��ߩިr�.1�.5D<���[���JG{��~@�.�vl�)cОf���5,�3�L�Vt#�ܓ�n��;�֍�۩��y[n��JV�]=r}�����^%�$�T�swܻ�6�y���J��Y�z��ψ�^Nf)V����K�SDGU�C��bwi<�wT����+ɻ�o��$W�u�.h�"lH�d6�yF*��Y]{5�6O��90w{�RyQ��Uw^�_x�=����%ӠͲ$�y�;ϻY���u�w9��Xަ`�wb��N������k����-^w���5nQ�d�����:qv��oQ����O$\��叼�����:�<���g���^�
��Hd�X!&�|��wv��ö�#j�S�aV��}^�޵�^�^]X�8��z1\Dͥ�;���'���jU��ݖ��i>���P݇H�����J�d��%��o��];Nf�ߦ���3�|�u5�i>Z�_w�X�&�Q���p���j�.�{C�>��!�5�W�`|��{c|���_�z|B�[aT�t)�M��vb�<�,���b�㸘�UX-3�Ka�U��f���Ȯ�z׵�w*g�E�;G���,��N�5q�LS܌ȵ��M<��ᛛA���-��V��:v&)����Uu�I�h�ڸ��Mifr����a͏����P�#w�X�vT�9�ڇO���*�Z���[����[~�����ym��+4D�c s��x��,��!�e^��x�W!WM��o����%�����U�Ww��j#����|���WI�>j���:�ѓ�+�m!�.�o(�t�up|�_��	����:t�.*��V��h΂�	��ų#�MfhN����o_���ߨ���z��cq;�	��&�����Y�����U|�?�~
��F��>�c����i���Op�=���ug��y�JÈ�^@y֜��\to��}�\��}}Q1;wK��V�of��:��Q����=�����r�6�������Ž[ECr-�C��^�d��D��l�t����糳O����v�\i��w��΃7Z�pk	���Q�;�E�{����ys�R�wp�.܅Y��Cr���W��(��7X<�NY�=�wG�}�&�{ה}��\���Wv��<�b<-3Ź�ۺͮ۴�uʍ��CU
zm���ʮ��'=��=^����QMA��x.�G���z�c����/[����þ��ú�=�pWv���SP�׍a����Cc⸙����v V�TI����g{�<�6db*�5����#����4/1n��N*�A8d�q���%̺�H�V�&�����U�)���sޙ^�y�k'ZZ�k�e��UP*��TONv`;;��l�3W ��5�dYJ(��]�m���m��o�3��N&v�-�ȦIv������V�zѮ��UeL��;��&E�,l�sZ�7{���Gu��TB�Yj�����¸o�k��S�U�u��2(��xi�z��L��q��(�=�{��)�$�2�y���ыr����͎yM,哺AU��V��N��˘�o6�J��ކ���;l�{�2-JJ�+J�J�݀q�����һ����F�s��#��<��[��j)��Lw	���oҬd�gB�f��!�f���j��ő�N�ܑ���;~�Kf���5c\݈duײB��N�yJ��z�Ya�ӻ�{��f���r�O�d�����6}0�������-=��n���U��7���{e���S�M]�Kݸn���j�ՀY䃺��l�x�kJ�'w+�z�\-)�[<�㷸�k��{�U]���Y=��(
��a�	����ZTU�t=���Yg>����5��_�w�Y�����SW+�=cv����Q�B�;-��`	MV�A]�\���د/�5b�����ܭ��w��9���2=��u��76�х1U�h���	�p�}JY��Sn������Kk�\�f��P5F�w	����\�w���RQo��3�G|n���}gcy+�U�k�S�����zA�J�����>�Z��q�eC0</_s�_������~ϒ��c(�Q�y
���L��=6�Fvj^�/LMOi�ir���Mu���nS�F���(��<�a�W'��#4H�-�o��m�J���wD^��W�j�Z�c��;4���g��=�����"^{��Þ!���3�K{ ����1��+뒟7ې򣶢�XGN�R&տ`����r���R>�إ1�+]N�˗����P���E���8�PUXDk9r��dZw���c��;��/�F�jq��kdB�哝c�˸���7J�N�Fq��j�_�!�X��_���ٓ2p	�ܩ3�Z�ܯ�W;��w6�6��~CO?�({Ce�V�'9��V�j�p,+����q�;*��V�jw�!m���[V�8��m���Գ/1k/�6�!5�
�T&]��Cs��Wc���KZh�S�֕�.� ��L��QO\��F�67r�f-ԚRY���r�3)��+o\��O�{l<`�����F��
�u\��}؀�YN�ײ��P��f@�(aYy-��6])x{=����H�Z��Mt�t��\���7¬臆��Q<�������^7�m%*8C�!K��F('yZ,+�l��X����)��x0ds}hTһS���T�$E�mL��\{��XA�,W��~fp{l�Ĵ�� ��;�p�=�^p}�&�}��ض�zb�o��ɩ������u��
�g�i1P"Ǝ�]�!�b(��w�T����}VS\��¬��|i9a���S�d�%Gg�Rd�V��+�d6lݴ/�=�U�i�� �qӼ�.�B/�
ү�]G\Cu��)�+�:��x�8�x�[iy��]Y���۶"��k�
�xU�[s1~]1±�^�n��ߕ:!��[ՙ��^R�w�LB��kگQ��P*Ѩwf�Umk<��ѡ7uè�҆���ͬ Z��vv��I�iQ���t8�Ю�gV� ��S�`S/�hX�817�w�3�V8�9D]Yr�!�Xt���]u��--wZ4�x�-𾵚>yRc�~zmj��D�8��ƶa�޺՜�BY&ez����^��]o�y���o��]q[(�\B��b��5��;�������13C�b+?>�qڽ�7�\T�9����KnXp�(~Ʉ<�\�!1���w�pT
�N��*�t9���{e�u�G�\v�X5y* ��\Cw`���,{��bs��Ɩ2�57��:*Icy�4罊��X���fN�Si�e�J��8���	dGr#ǜ)�4襂q����Uw+�{ނm�t�c�6��tP'z@U���ZW�".	'U�3�e#��V�Z��ڱ�G��cJ��ڱʭ{
'0&�X��\�l7u�R�^���p��%�)�Rd1��0�mF_�a١���^�>��ƗO*����G�>�*?-����r�Vǯ��.o���x��H�Q�|i�a���t�~5g�l���[]x]��^�s��j�8�W8�a����Q~�d-�/B߽o�I�*�&
�89�ܚ�Wf!��Sq�i4���xi�q�Y��	��N�F�t�I�ʀ3�`�Y����W��2�\���̉k����}��>�o�c�2�Ӓ�þ�g�Je�ְ�L�۾�_���I��IO�I	O�$ I(B���	O�$$ I?�	!I�䄄	'�I	O�H@�Y!!I����	' �$�	!I�$$ I?�HH@�y!!I��BB��I	O�$$ I?�$$ I=�$��1AY&SYDUE�Y�`P��3'� bLz�����}��T�gm-�����(�l0LiY�ݶj��f��*��v�E����&��P�l��f��n�����[35�*�K&��jm���v�FY*wV�ڱ���֓�k�U��fl�L6�l׸nf��]X+Q�=���ked2�s�6*m6���Z6Vݺ�n��D�4KiSj���{�^�m��ݻ5�g.��Z3�AZk0�Q7X�7]�w]lջk�1]1����ހحl�a9��ӵ�n��0�m���ӫ�SU��3Vt�X���-�m2*�ƒ�Vٴ�
/�  .�mO���n��7uv��NRU�v�r�����"��S��l�\4"*�ή;m�
���w#��*:���ۚt4h��벰:�;-�L��-�Y�  �  �S��5w\����:wn�wtR���6�����wnu�K�:jK8S��ݧvեw-�]m��%։;Fwj;��8��Wk�Ԁ��ϳ��V
���n���  �R�����֠�B��<�m*�T��oN���sc�wi��F���㶭4�tլiӡ�4B����P�C�B�	����
(PnU���
(P���Yi�۔uh�p     �}�(P�
 ��� �(P�=�
(P�
(\��w�4{���,�m��ӌn����G}�v�P��۵�@s�Pf,tu݀{ީo8�%�  >   {��CZkO��#l骺��׋����w:U
:�Z�d�r��4��K5E��X������R�m�55�vm�Ӣ��,��������X5|   ��>�J�6�W;m����WZh��5l4:ö�UUWc��u�vtwujUQњ����mۆ�
*Tv�ܭCj�w+Kn   �   ��65�ő��M�QUJ��B.�)yt���������[���5�.�9�ۥwp1�.ꭷ��݁�m���q���X������W.�   =�_S[�Wd�v㛇K�Թ�kv����ړӮ䑠6���ڴ�����U�ݝeJ�;u�ۍݵ�k*5z9���a���jۦ�\{mi���R[Zq@ �  ���i݌��E��]Νk��*��@n��nk�MV�wr�Wv�t��R�PP7.gt����j:��uZ+Bu�#l�;�mJکu�O���Ն�ۀ  |  z��t)�X�V���wn�d.v�-�k��)J�C�S�@��\�ݛJЭj�w�{��(l�;�k�C��3��+�Uw��j�N�(u���@eIJ� )�IJR   jl��%��42���R�=@ )�
R� d �H���H!�#�??�/������,~�����lن��S��YS	��ݒD� #(�+&8X� �"#ބ	&s{�3��IO �BC� �$����$��$�	#	+﫬v�����N��D'5�#i
=���4�mi�Z4�!ފl���x�`�a��n#��9����X�Tfi�+�b�3��\$=x�a ��w���*`���Er 1� fEh�׃q��eY��/C�	Y�^�D5cv���E�7��Y�1�$��mn��g*��EB挕w��U��.4E��Y�v�j[Ȧ*[�Gu0����j�Vn��Y���E��1[��o׼(�)�H�<V�T�P�=���t��;�����PZu�p�ȠOB�ˆ�F����E1����:�G���f�Z��o����{U��*$�֏v�Ӷꉢ�Ǖ�NR�d�6%��v��p.�P��^<���zΎ���r����&�Y�	�E�f)n��P�!=�GSs]�?!P���d���m�H�76Y9!��1�{p�ߌjc�080nn���u{��ˢ 	������Y�M+�J�O��`��|�`}bn�x���U�"��C�N�=D"7q�eބo+kQ6u�	-�����{��1#� ״�{���"��J>-{�Є.unq���c[���O
4/=hѬ2�yx�*�{������5/{��簽�+�*o��Z�f�/+v��j��Z�KiN�1h���b�*[A�1�&+02����V�M�'�G�^��Tv���,��=F�5�N��çx*��=Y����*����u�Z�$k&�I=��24�y�O8�F��x_�'��\}���_��+�	E��j*�ǖ���u�1G���Ϋڌ�.�-7!b��VĄՒ�+��P�MRզ�Xu�[HK-G�Y��1����U�c]�����TTZc���hMwVnS�@^���wc�(s�t}|{/F��Nl�X�^{��{/'��������톞q*�J����<�]s�XG�6k^�;)�+i*���063�U�iط���J��ܱ��k"z�k;�5)�n��[�!	�[��GX�c5�g7q]�tehop��)#���Bb��7�fIFX�$(6~ca��-��7A���-E�X��k)Y1a�A��n`���1;�ݥ.%� /u��>/�H���L��F���t���'״�5/_���!Y�����{%�6���e��ceI>��v;��V7�1�@�����9��sql���)0
p�$V-C������1RŰ:���)Q�_/ �^�]��l�5�8�`�H�ʰ��N��ĬX�B)V�t�Çf݉�j�&��޸j��W�(#c��D���9�v}���V��+�}�i�����8�߉EVɦ�V�7����-,�)��."�0oܗd�@��o\S�\i6�5V9�C�G �yu�}5a:��|O-Ϛ�>>��n��[�
	��u�-I�5}�fMr[ܬ��J%h��
qY�#Ғ�ʲM7�mV**�����P�il�F���;ڙz%�Ie�4����6M��V�nL#wb������,�I@��/mO�Tr�I��)��n+-A8$g)���s	���k	�~��v�4�*aX�L6��o	��,�*-� .�4ܭ�x�%cm��E�(�K6�*w;�#2�S�Xn˙[� Ϧ�ԙ�M-��L�l�M��AV�r�!�e�׫2�lH+uu5hKK�]�U��Yv�AL�P��S1a[��~pmTZ�jD�n�#[� )	vE咪��n+�m�E1[�XSiW��Q^7s0@��� E�5�KS�j�5��y�TN��H��/q�{��v�+LAV�����Iw���og�O��p]@�`�OBe��<=|U��4^���B��Ř*[�e��*�����E�M��n!�}�����G�����V���-O>�%�����9�Xee�\�gk�Mޕd�7��x�{\�n�����`�%��%���(�cUe)����ڲM1l�4P�Ų-f�bm�������o�b<���f���9��p_&���&*lm+�v�Q�}�]m�ռ#���wLQ���j���84f�L�"B�/p
!�j,Q� ϖۧ����;e�K�a��n��^�ͅxovN��=�ª��Â,��.�U���j����.lj
	���QK(!G~_,(����;3oCR[Z��6ȉ�8xw0d=�8/m#�G|Y�J�W��ߵ���&= �����V�ҔU���b��|!�^�#�`�}���[/i�t�S&� ܥ�Y�І��KS�U�-eP�MS�����^n��q[/�V�>:�EW�@I}���t7R��#���������W��b�@�e�l@�VԢ���"h�T/�;=b�{;Ǯݵv�n�ȕ��%e��-&�Ƒ��w�-�-�e �����L +PcMS�&k�����la�����^�Ů��m�&t��O=P(>����/�~���"�;�A'�j(���L1�*���;h�vLY-qN��B��j��f���������1��Ryo9s��:���amn�V�"�R�.j�iH�v�v�<GK�N[�OG�m�'�pi��v$�=Ⱦ��]Ĭ�J������4���C�%_�IL���+M^L�ض1���w�˅�3:ҹiv���O�!�CT*��ܔ�*�#�{�(u{���E�1sv
f�5��׮���0؁& \M;���)�O�,�b����t�S"�-�J5!�٣%Yj��WeU䂍��y)Pf%�(��[��)=ֲ|弲v�B�~Ua����%����\��B�X�EV�Q|2�j�(�%`�N���%H&L�+.��ېb��.K���ϒۀw� ���SKHT.���^iz�
����5큞�Wf� �Ղ������Ek�b�f�)�!��r�-��ⶎ�4��@+�J��n�cA�
���BjC`���8s�܉~��J��/��P[�#��ssj��+ٍL$^M��fw�� ����ϓ�O{�C��\a����i�E��{�Ui�^�hj�R��˔�1M��B���t]�:�8
����í8�Zʒ�����%K��4iekȵA$��6���n�nܧ��Pޠ���ak��M[�)�CVN��Nk���@0x�������n�z��dAܩy�:������ ���YzŲZ\緷ŊR!w�D�:w��h�BM�րq<��
;�j�h0�o��f8�35����;��6�h��ܙ,_��o0j�9[&�X�=�(6��UIu���ܲ�nVV��V�As@Oצ�
' 
*����������/�X�vr�Cw�%3E��
�jcxiS-�%0�vLb�j%]��÷�o�m��i�ol���c�@f��X��?#9W.���N ��(���63��/aUڀ`ȩ���)M�½t��n��7{G��� �3Bֱ	�)��	�KTh�򈪣q̧5=e�9j�o/L�#��:���I¯�JO�6�r����b(
���z%X�X�3���؎ލ��4����P��L�orc*Ғ�+��%D�lr�̑�N��2�л��6@�R�-��H��n�)��r�/�&�V�^1n�4B�v�	X��Y.Q�-�YF��P�����nm�� T����4�Sl��>:���!J�E5o!��s�Zr3W=ě3Z�K+*�۽>�|����y�����X?`���VK�kC�ZF���r�
����*�U�[�`DcS.�1�.��C �G/`̨�/���N�SM�Gqf-R%{p�[�:֭������ThT�:�5��Zj�ܫ�CmCf�)fX����R,�M�k��%B��9V5ôBe��5n����-5�ȯN7bh���o2�t^��6�gUe�s���CU�f����������0e6Ag	#ra̒:���V�=�駶"S{��𰊁,���{é>�;Ӆ%����CfV$���jx��8�e��e-�^�Y��Q����H�f&������+��aU��Skl�F��O.�(�P�-ڔ�7%�N ~�ց��k�reK]hbT��n�Նn,^e�aT�����Uں;��<��� ��X*ѧ�E��7Q����N]�X*ĺj�]%�^l�MR%��A�f3bӣz��G;#{.V�
�Z�o/,ڀ�?!��Eh�+w�sl��a�.�ڧ�l[�F�8�ٲڭؐV����r�������q1�[�!�s�f�3W��#/
��*�ksm�fZAȣ��� �<]��ݰ�����gMY�`k4�BfnR[7��ԵŊ�;�;���\s>,�	�T���i�^콎JVIyn veּqJ��rټei<p���ԙ���(mM듰g6y��ܐa�`��az� ����
&Ek�̐��ݺřrh�a�0+P��5��4�u�vkl�unRsaΎzx��wˬF�|�5n��+��4�n~��D5��G)ڬ����2��i�wM#r���[�55�h�Cቜ�ňn��:Ў��˼���u�X�7Ze�@(�	E�2��N�vH-�u[yX���5i�lү����<�:���0:cr&}\�s�X���􁥢�7x ù��a���`E��
��=�B+�kQ���
S
�K�H�x��J�,�{ux��4˹�T�\$Aܒ��F�dT� �r��깺��Y���Ͱe1�1��M
��h�ɲ۫'��6W�۟bt��SUƛ}9y��֪ak�%e��yiH5KI'{��r��A	��8b�����h^wmF7V /
� �p��Cji�E�gf��eE���$^�;O`���Tf	F��P�KפyCr0V�y�:M*�,�j�{Qf+́X땎*Uxk4&��f����-�V�zhXʭj�,II��8�.��-ꡘK6�Tԭ9�L�fm��Got���G��@���ܞ��w"X�A�P�������>{B�[%�X��kq-�D
�r�T�v�K&��G��g��<wu�Ӣ��5��Gٯ+N^�MaVj6�k����>�""��͋T�ۃ>�Y%�]�ڏ��`���%1�KAP���-��u����(v���R�����/&df&�hҒ�w ,[�.��+7��`����i-
ō��ZË*J4A����|�V����Bi�,�V<�6��n�������؈��y܀��OiD��#�8�˫���Ӏ`�;���:̢�˴csi��6αA���f��R7���ͫ��\h�p��Wv��RܕO\��P�O7Z#����#jVk�5����l�d�q�!X�0Q���U���j��ZI" u����Q���M$$�<�6�B2Ή��M�0�X��QY{LS0�qV킭'�p��WXD|��{t��Kϱ��&�p㸐)c@�3����w��K-������y���|BR�9F��#�	.���b��yzL�`P���z��tS�-��ƾ$������uz�A�-�x(	R��Y���On<�B�8�5D��O6�֯kn�A���P�qPa����4��E�c�)bI����J�m�
��ue�$R�7wG#����ƻĖc�=|�j�c^�ik���nя��~�p����ۭRMH�hM�7t�Z���]�[5��f\q�^�9���� N��Pm��7�ԭA*�MA]���<5mfK������djZ���fy�^�**�,*2@9�I6ͧ�-��{W�;�JH=���=�v ��+)�U�nS{�sh�JJ�r��Vޫ�&r��=�9�v������
��t��!��ǥY�	��Ɏ�^A��Kp�Coe��N�;n�') K>#���A]�'Zv$�X1�tSܺ�F��C�j)�rP{Z�E������ȕb�M�P�=Ԏ�m�t����򵭺̨D�����K��k)�Խ�Nx��@�邁p:V̵f�dk̵j�h��gϐ�Ng�S�o?%���+8���yB�Gf7~����Q��@ۛ�Cx�nR�,3�a��3VVf�D_|�% @:`4��ĕN����Ņ�^8��<[��i���R;����(�ô�lj{��K�g775��I��m\����7iP5 �Mx�8�3��Q�zS{x�K�{�p����|�ɃJ��-F6�N���]h�d��7�V*�zd�����	�)�O(4�b�ݽ�Cte �28уfֺ	!f�V�2Ԑ�������M�Q�T�bZ��A��jU�wf+g ա�	�Hբ(���� ��7��ͤp�w-�Cf��T���p�\�����)8�2�)c��e��L��7%#I�,��	VSL�T�Y֧ͅYz�A�
�2�&3�x���!���6(�*`�C�7�9h\��i��+M'�+K�6M��̷a4�{qj��x�ݔ�*L��(�f^�!�ŚI��
�P���0�K`R1&�1Ʈ��,g���
���ؾf�SM��9���l�^�W�t4Y���:_��*ʰ�U�Ԍ�R.�p<�e����57�����{���� 7 ƕAI��
�����cJ�E�>��W��|�j��WN(���X�t�t3A��
m�이�:���:T�C�ƔqE`!yc3?���j[���=�O�)p�qM���Ul���@�u:���i�gUֽ�c1�G�5-�b�mde#�2U��T�z����{�s:R�v�[+#��GeV���^��r�$�u�&�y�Ҿ��St��P<Oe,��!W�T�S�T�B�t+#�m�]x�V�nݬ�WO!�r��A�,S��ƭ��\>i�s����ݫ*k�F�d5������� ��Y�gYt�� �ʍMlIb�9JL�J�i����:Cwh�=��M���;�ؤ��D�>
?=���������~�s�
I7�"pg���N�����kM��U��V�L`b���ȅ{}�m@h���@�4�ipt3G`q�8�9�4��6E�\��D$T ���LM����ٷ&X�Ƣ6���F�:hI)�Iα��k ne�Z��,*XQ����f���t�����tϲX�U�sg;���t_<�R�P�<q^xS�G�q�.ϗH�V2�K��S�7Lz��(�z'
Sm�[��^wod�}�,�Rz��Dc��
V~���ŕUoPck�px^z�
]	�7~�K\x��#+V��TR��`#����:[��(e���]��"b�h��-!��t*tӻ�CVa�}��k����n-x���]=�{�kyB�����v].�D-��l��\�X����9W�>��n�]��b'Ph���;7�{[���V:�#V���ñ:���di���ina��JwW�*Do�wa�8QYt��h䤄ԯ[:�J�-�s�w�ܬĕŧ-C{Z��\�H�՚��E��P�����f���"����+���u}I��u�u�--��J:xeC,9�������u�*>$v�բ���^���&�ڠxĞiֲ�^X�b�
���٩��~4� Ø�xoQ����.N2�ݭ6�o�l�{*�.p�)Y�/~,8��o�iaҷ�˾{��t+m�sS���n�v�T7�<��Cw`�b��QYtB��	�iIy��˘{����D�JT�����vZNA�p;,ѮOܽ�F�J��u/����WpZ���ܼ�*^=t�W��4ѻ�3g���B���[�&(h��F����-��Y�=��I�#����-役	���EZ�l�Ӄji��l-	�u�R�Z�F�JD�o��¢���M�B�x�`əG�e�y�y5��ʹd6��[eų��w�]�3�u���L��)��^��OL�m;J>�y�U���
��6 z�ܳ�Y�>��ɕ��j�"^Qג����=��cqlح��j��&t���,�-����5,�ST\ծ�w���b�堛��5�ӾlI�*f�1b�UǖQV�f�G��������z��OM����ŖfF��Pל����;:����r��-d�뱣�Frv2q kt�	���B��ʌQ�����-�)�N�Aϕ�K!d�[�xB���&��T1��$vX�ΰKf�}�-�b9���qY�gC��8P�I*�7y�s�P&g"^Ԏ��Q��)fsٲA[�oL�h>{���v�2��zH��˭�w��!&�.��0�r4a��C���ͻ��`z��@n	,��4�j���Y�����Wx�oXx1Pk�5t9�l�ٶ�;ON�(i5٨v����i	[�ᩇ�����i�j�׵Ƹ��׎��]s��:�Nkuet�����2��vV# $[q�e�X�u���24dZ]�*6u}mI���QC����j��_]�1�:U;OR�jn�Ķ�\3��1v�"�uuq��H&��U {��Z&���
[�N�\�����λS���׊,{x�;B�9��«��XƊ�[x�放(�nTF�=I�*ǃ�������K)|�l_r����,��]%tb��cӼ��T�Âk��!~ٚ�7"��ɚ��m�Ĭ�o����cn��z[wݱwj47%
ް�F�t�λH�lRCP�K���{��0J]�V8T�v,KZ�/�I�y�(t�E��E�	��]���>�O]�t�����Y�Wң�����]����o?#ɧ������d���E�d ��N19�tfֲ/N�+�bN4h	�K�դh����.�Mj�6B;9.wtmr�0�8�f��,�9KW���*�GW|��n%��0�E�'�K�[r����ْt�7a&�U�/l�b9xLp��drJ�I�w�E�k �Jwy���O�D�J�.�5�41wG�{y�!��,��K8�.LJs��H23�������7ooͭ���b���|�.��ۃ4j7Q.�]7�-̼�W-���xH����|$h �	�6��ޖ��?����+����Y^�R�GAg���aK煝Ja�ڎN{��Y�K0�ʾˀ�Rv��جj��j�H�ז�b�l�@������)�.[�������c���ݺ��u�5j[G�#��{z�[�b@��R�f����-iP��v���7r��ɶ�ٻd�@�8n�m�C�u�e�p��ɕ�0�����4�r��cY���Z��n��7��Y��]`��V
Wo�p0��|Ff�g�=˧	ۏ�Z޽��K�s1�](���8GgwZ+o�3 ��Y�i�7�4Xٚ�x>ϻ������\YD�t��V*���n*1��t1�IS��-:�Syt��S$1b�na���&,�&�^@N����gP���ј�V^>@��\]�+�,�9�����/2�ZT��jmL�mye�IjY[�D���%��<���uf�Q��2b���sm���7Ow8���Վ�+��V\��x5��z�C)_ZEln�K���'Y���v&k�<�d�.�3�{1�W�l��VF�A)��L��y���h�gM[��U���,��q��F7u�ԝ�ܱ\��0�W'7M:�S��`h��A�,��T��ݳ�J��z;4^D���u���zѐ�:����9se�F��}�_�c
�(#o��^����V�-OO�uv�G����x瘸�{O�z�OY)�*�X�r�n�K`^���1�����s��K=d�=Xܬc�(`OY��E�����m�*��]g��-��K6�6{QL�$�²E�X6�R7����(S�ۅ�*���ܧ�':]0��Vm.�h,/��n�������w���Kft]�䂚h��c/m�ͷ׼+:6�3��8Q�<	�@����n��XU�}P��{����dc(�=n�`x��D��"�������}��K��m�[2���KU�I�m�f�z�4YᎠ4��V\Y�o!�3��vX(�2ΧUun����dN�	;�yO�e�Oi�"�	nе�,��,��|f�%��+���>[Na\05���9Z %jGYdK6��h�*�[��
��"F��7�n��7a�R3����|M��:d�o��Y��nS�V}F�-c�ɇ.:Z(ŵ2�Ҭ�ݰ���u�H٠z�f��/+��Q�_�gz�A�����B����<q�c��A�����ncQ$Q�V�=كJx�k�0]HŮ��,۠�n*Uc7tV�
3�sn�lN�G-؝oL��8�AٲB��̎,`86��*�uS�B�[�1�l��K���c[��lE�[�/-g�������z2�9�%�΄!
�Z��/���T����q��*[��kg(��-�V
���2h�b�t
v�}q���ň���1f@�m�Z�I���KGW<4�nĪ!+&s7��iBݱ�ޱi�ǜ�6�gv}�����$�Vحھ�ѭ�N;��;r[�"p�2�j�8��Oo^��RgVYz]���9� aO�z
vv3}�>t2Ʀ���+o�(��m��Y�Z�.�cZyf�5Nu3ǵj �i10�%�2�+���E�^��N*�D1VQC3t���u��XR�,�f�	NW&����{gwnQ[ױFYg@rs��!���N��'XCհ�B�g:��e����6	t�6���z6�K��`�8��XL[)����/��²V�O��X�C�]Z���Qݑ�lv��z:�z�M���r��33Uj��[ܣ�v�
z�]kz��c�9�X��[@E������i���qr�K��v�۫��jݑ�rN]��"�P�ȯ��r��e��]uhV4q]��o�ڕ���n�b����$��͞�\V.�s�f�.��{o:��)V�&tZ�t/0,��(�Ug_�{�2->��f���t% 	�,vӏ��4{;��-^V������%\����[5r�0fM]&s6^�\{`77K�s��Jp�/����Zg�1iιYt���	{�<@�ԟVM��.\���vu�o{8��-��/�Irlj�9LZ�1�j,	A)�H�92�dN��d3�p5�2¥��lYX��w�'��'�ݴ�3�6���-���	�����Eح�.��ٚ��DH�A�a�Z��7���7�N���=��,R띯�V�r٪��B*�V��M#'Z��i�L<nQ}��q��c��̋��C����B��U��F�Ij���a
	R�
S�K�!u:�1�'U��6�1n��T��CсK]vP����X���w�+��U��T7Yl�*��z;�v&)y��d�ůj�:'9@�I�ojA�w7U`�V�חOR�"	Y:�hD�&�-��r����k��gX�ٷ����vHf�\���ˮ��N�
}�z���i�����|�a�%�S���V��x�C]j��p���»>{"�Deg��Ă�5�D����sB?!��h��"R�F�	�֙�1�{wn��3in�~�lH�s-���w<�:��e���*x��ֶ[�B��;���X�V6�����<��S7�����
o�M�K`jj{"����ZY���T�b]�z�[0LbЪ;��0nM��u�Zz��D�t�n���P�
�%�愽���]���p-�"���):@�[P��	0��se'Y+�����'��0�t�wga�'
�cFƱu�w�zEW<�M�cT}��S~:p#ˍ�F��=��i#�a�(�]Kࣦ���b1�u0��������o.�]�����M ���\J �m�� k�r���I�8���h��s�j�tb�L��
_eO��%�Z��rJ?SC�S�t��szs��lu�����i�c֭��ٶ7;#V�G=�/)(3�+#h�W������q�R�U�L�.��D�۔'�`�u�P��j;��^���rz�F�q�끫R/f��W�ñ)
�\ '�3s�茡��dv�(YWKz�9t-^⪉+hh1"0̊�s�7���z��`gȿ�u���dڨUP�G�-O����l=d��)�}Ƶܸ���>zV��MY���1j����v�Z{l��G��][��Q���v��E���۳\��'vbۮ�f�nɁ,|2!FY���j��yE���;�JˈEp�@>M������&�����',�Yl�{��펯[����D-�U`��v.2)==��%��wr���p�kXΌ�+L���U���Um��#B�jK���WЋF�u���6�p�ȬGwl�iZ�t�2���'%�ɲ��&6k��ClK�#+U��LRbN�J��&�4�# �E�2�6A[u�"���U�\�Z�g�i��=
��dc��V݄���E�Sb�;ed�okڽ�kܛ&N!����٥B.���5��hb:X8�wh)��U���RjY�yrhM��@m�a�uז���*4��t���6�Z����މ �
_:X����zU�x�n�tIm�2N�%%�b�n}��Yg��Y�kp;��l��,����U�p��S��,��͉s����n�[R��,��M�s%.�Cxr���B�V��ޜ�Dhs�6�}1%�ܛ���~쇇S՝��W��H�������v*)�ka����9t[�z��2��G���Q�B��w�����ώؼUP&/�pc+Hi.u�t:����E�o���N�H�G�f`�)#D��	�M<�8R�iN��{�ܦRc7&pk6%�;���X��}��m�|�F��4+�9M'����Xau�!���^��Y>gP�y��6�;x�.>�Q�>f,Ts�S�|�n#Q��#��zt�.�ޙ;v�I4*�6l����F�Gvn0R��������mo[�SNֽ��9+yd��.�ط��V�xr6F�q-�ޮ�3.m��䮅Eճ�T�KB�u�k���0J���;#�۴*��aL��e��xaRL��XvV�&I4��]�Qc4�\����L>�H����#�1r�Gfg-6�SՎ����F�b|���HQͱ���RG4��Fj�+�Jx��\-�1
;�1�|���S؈�qZ�c_e�壮�+
�Y���abnR❵�8�� ��C��]��q�T��R!�U2��!l�{�e�/WΆ�q�����f^�V(Y60��&��B}�LN��#6,�[H���uEwH����ȓ��F���j�� ��K��9^t�\�"wQK�b�z����m�n���������e5Ïe������v�ȩ�x�n��R0�p��n���8�P���Nw��?M��ת����)x��ػt���t�K�@��V1=��B�EYݶޭ�-������̎:���u�n����ƈ)wN�.���� ��>�yKUkM���X���IԈ��p����xȗh�hog����8�D9b�lvq�#���C�(�KGed��\�f������<������$ I/>��w�|����o]��=�������	1=��]f�ȩ�eh���w�﷮��0�ۥ���]��V�k�6�=����K,Va��{a�+M$y-6�z@΁�\����}p�b�\�w)�h�����ʶ�r��K`x�Cq�E��oZ����[�B�;B���n-�9�MlkZ�]E��,O#�dK�>ʭO���Y3X߃(ҍ��\�V���ށ+M٭����c���Kz��4�X3�<��/������h�^�;���t�u"�6�wo��,�ܭ���v�iOꈟ�c���R�6:�k�lV�Y�ݿm���|�����b*[�����i�4>�6)�;���r��o�[�y��oz�#Z6���ˋ���#�~��uDP�܎�iج�+���	3^��d0�"n�������o�t��<�5i�;o�Ӈ��#V��1�{tRE���F��ʣЃptӰp[�E�ŭPY.�77���e@�lM��ާM�ǅry����舵��I��ܻ��Y���$�!y-8���D�͏|��_:Ǭ�a�|[��٪-,kJ��.����Unp�����8�{h7U�&�57Vܰ�jkeMR�J�ӷk��ȃX���n�����}pч��ʧ�/S�*§�q����� �f�]5L�Υo�Ppӷ�W42��֍C�'8&�w��jI�f+v;����|�vF>��3ib}�&�����WZ�ʊ��z'+((j���åb=�L���b�mk�L�LxX��ե����������]�@GZK�p�'b�t##5��M"{S�O��2�!qY�)���`4��QɎ2._�We����U ��%p���hU�*���q�,귃HܧV$�w�0]#9�V36���3�I��hX��wD��ޥ���G�m�T�e��1�8�6�5��!J1��Yva���#�o�o7����/�\}5l�(|�<��s<����¦L٢-��@�[�c��	3u�$QTֺvpJ�lݪR����1�3U�q9�m&��x��U�P:r��r��յ��F-�� ��,<�q�j�������&<EV2�c���f����6�+tv�x�1L]nKͅ,�%������e�����Ct%�N,�b�s�HdǕ���Q�ݼl��ѵO�I�ʾ���JL�E��F�|���ֿ2rѱ��l��^"�rڜ��&�ɬ�VJ�>�!����r�>��eh�|9��Ă�,�s;wF����Ye:���؂� ��kjP�#��u)[f������7d�p��\��P:^i�lU����
��e�L��?�n��w�X�����Q��k��ԯj-7�#����&�֯w��B*��@��1α��Ҭ��5�2�'Y��MV,ǚv�Od�nGY��V����\�p�3��nf)�ҧX���3=��� �LU�k�x
:*�A�-@�4�e��bL-�ɦʹz��y�(pY��9W*n���w��C@}]GJq2*I�x�����&kK�{�Ֆ�AR��t|��ֻwJݜ��R�d���Zۀ-�+MkΆ0C����`�'��x�څ�*�e��\ڹmR�7�J�#3�����PMgi�p�J��6���^�P���3S�g(M��b��G�vQ]a�����gT���m��u��CBX�+:�xNE;��
�SwH����Tp�֭^�kSB3
qŻ���Z�Hv�/�"��ٸ�_m�����ɈU;>�Rq�DY�L��]!�Xv�b ��p�HU��c��cէN^�y�j�1��8p��k�#s�u�{̞zS��(˥�i�M�v,�*�U�jå�R���z�qv</�S�r��Nž����tne�C	=���8��J˦q���>�ʱ�ı�ϞX�_V@9&bL�\�+��Si����C������D��e@�oIYCz��C��`*m��<���Qk��k�s&ɮ�q��֬������a�Onؙ�-�h�q�MH��L_-�\�ʵ�l��������[�r�@�:Rjz2�fw�.w�6)˸�E^TZ	?,�O$U{HU��+t�cdI�w^s��� M�wZ�w�S��_��^3�Ck����wk��*<�mm��ۉg[��d��$�۽�������29bҪЩ�2`b��w�&oMKkh��,�T'w�i�ʵ)`v ˡ�l��lk���̝<�׏n=G(T[�MSh��j��@���1~X�e)�&A���t6,m�d�N93D�,i��C�ŢnW6U���x��s1ʡa�S�`x���p,�:ty}�$�y���������� f��:�T^�C<v��w+�^�1�5ܱ�-�&8d�p�.n�(Z�Faۮ7���g�o��̑:m;�c��I���l��ּ��l8n���;�%Vݧ�����^͜�o(�tx�!!M��Y-��wW�St�9� �����j0z���;{A��G[l0�lO�V�/0_M�WNE�mH��Vh`��#Hmc�����)�R�{giV�-����U&<���K�!#]���S�˰�n�ۅ�6�.Pv�;��"&VT����f��Q�{���<�rjS����5R�r�ݳG�N%Z��|2��eK���XwƋ��Gnx�)��h-���2.�/O7�M-c��߉�<y��ZT��!�ZS+wp@�;Zn��ݚ��FP��#(gKv�|��5uep<�u��f4��z�6dW��h�ˬܱt.��)i�˭�a}cfQ�}0bH��-ȷ��4�".����ܕo��I�m���K�H��2+�t�ۼ������	�=��
�	��[tGM�۽��Tq,	�&hŷ`۴K^�Iޝ�-.��P$���2λ@0z��;��00#�{x�@ǷƌOc <'jj�y���u7�Ь�VKxrT���Z��&u+[���K�]<��Ub����;��$򩛃�UIm��U�;���T�YT�H�v�2o\K�8�������p7����0�h��N.�P��lU�/,Z8z��S-m���Q&�Pu��z��*�Y�T�h�B�
��*�)��;����]�j3�ۧTD:Y��;1,C�����N�ym�bw
U���'��
wܡ�����#�TT�������^j�=��7$��<!�#Lk�(JՕ<Npܣ %P�N%�v��Z�9{`V훽p`�V�$��׸��2L��[{s� l�!�p:7���P|&U�x��ID(]�qb��3��%\r��"��#]�:doWǳQWnӧ7l��ͻ�ݽ�v<��8��ܫ�� �k�XdX����ժ�]v�9��e�a5	��n0�u-��tn`�i�D��3�1F�+֥l�Nj�9�VpZ��r<��*nq[z��ޱ}��R�bV�ۇ6��U�W�"�l�\�p�`o�����gS0�d7��L;N��٬��btY^�z���aO(,�#s�u1�P��6�j�AS��M7���9sԶ�'�;�ѣ�<��l�	����f�q�v�AGEE�T��X�hrJ��ld���9�5n����9��՝�PU�,���IV��B�Z�I}��C��+"<~`3����YK�r�ڒX�`t�����iP�e�n���1ZB@L��h�u*V�+8��8p�h�G�p�eٴ(��kQ�B�kQ�/K8͟�Z�͊V8!�˷�W��w����{���XҴ�;u2���&�Ԁӻ Г��y�(V�ZD��4w.���I��Gc_Q+Iz�ܺ���}&�82�,��յ�e42��<$d�Y��W;��X��ew�R�p���R�"�n� zyq�[f��P�4 ;�w�V��/(�u�oV	���Aκ:t27�vX��QWH���$*gk������অ�p�Vj�f��2�v�7<$)}w�iZavL��p����~z]s��޲/+Tv�r� ��ɌCC�_p�3Ԕ�88���Y��5��z����CF𫧵��N��:��e�K3V�A�>��t0G�/W\�e�6E-�֞�Nf� �V��{���\�4�
߯.�'���)H@(�M�u��u�m
���O�(^ے�s��RP�O�]ޞ�˚�`�n<��u��7U�X[Zn���^����^=/zToq�!�K>07�p]6vHΚ�.nX�Ip}h�zx�$JÆ�.��]$�fփ��rX��=�ngM�	䠽���{8O�����>�Ν{Br&��cDQ6�'�����q�df����p�y�ڠ�]�ݙ;m�\x)�7z1cKխ-��k�L-��Y�i��q<��UmR�E'LI܋̋
x���qS4L�<Չ��5��$#�YՃbiWXr�	ޛf��Gɧ�`(WH����7��E�g�hS��9S$n���[\��K�ge��^��.s(sy�+ΚNaL�)H���:j�r�N���f���[�m*Ŧ��V�w���5NI��0�u T�騴��q.�U:ܥ�y:i��Z��krRK%պ�#�vA����Η��{Tz�P�J�tE^��}��L<���W�
X7 �<yv#�y��5�m+�*��F����G�����E� ̶����kQ��u�}ڊfmM�:ii �uθ��S{}�H _˸�͵�_��rv�1�޼w%v�ZBq+�]w�^�7vt!ֻ�Bf��F�R�=�� ��3$��i�Kܮ�Ah;V��QG�	�/�ѡ)i	��Y�h=xYS����B�_N����x]vl2z�q��w@d�]�Z�ܗ�=`q��]ݶ�PM_Z-tX������N��x{H'�mrba��5�\�s�pm�"Pe�����f��g/HeZ2$6��C��HP���K��f-ܓ���5�ܼD]����)Y���]vJ^d\k�LrO4:�������tn�>���љFV��u8���V�&U��9W�<���wEFF����.�^�(��ҳ��isqj�
Ɯ�ʁTКu�$�LzM�J]x�Je�]vj�w�t-�j{�a&$�Y3i��X��SS�%��^�Ց�X��s��Y�Ox�����������_ܧ����5�� ���������$p���0�����A��Z�F
�5ӛ� [Z#��*Y��Ѽ�f�,���6zm[��R�El`^CΡ7�vY���Õ拊h�������ѿ˱<���um���^咧	ޢ�86�z��}й8=]�y�(�!���v�	��s�����k�m�8\Tv]^�!��B�\��[&�QÏ3�-���hȨ}c	*�ք�q[��u�A��:q	�Eӫ��b�ℕv�%L)-��Ȧ����[E@��K<nu^tC,:U�yՉ-wx�����(K�5L�����D�UǼ����#Y�����Weʡniˢ>d�\��);�8���zqXT��xPg�hXh�=Ѩ�C���]��E�\)t�Hr���p��7��\Rtw���(q����3����V_mF.A�אJ�|��׆��%
ɹ��2�b&���:�Gr�#m�Q�s�Ŝ�X� ���,����p�wHPn-���k�-��p�x�7|�S�V�e�`�|
[Y�6o��������y�1t3Hj�)�Y�≆0��.���)��4S�[��,4�Zj�,�RK���GD����{���>w�Q�ﲷX&r�63Ғ-Թ��DL�s�"
��f�<��#:���\b���J���1�G�!�8��Pm��f��mP0�W׸35�y^�WV�<���V^�a6�Ji�B�'���ۥDV")>�wnK7�1�dt���Ҧ��H�F���[C�=]7�ʵ��i������h��NU�|w�ޔiV��ȭb��9��5���=�c0�>W��ұ���DZ�ὤ��W�/:�Xq�)N�����8����1;l�uO4�3�+|Yq��m�R�t�Qv��8�*t0D���f��r��;E^������R9q�3n�ޖ�����	F�ֹv�Vh��f�3�%=|�h�AJ��1E��+��bU,C1�Wiuu��I�NQ��lo	��<S6��ʺ(�'m�!��j�N�-��jCt$��`�bN��ǅ�՜S}��VӋ)7�3SΫ*�����qm9˰�/in���c �Jю�f��B��|,#�Ifb�p��Su]@�C:�ۼ���|`L+�Kk�=��̛`�~��b9Nf)i�y����js�U����;
"�W��j,Sc�8�= >ܮñ5"M &f��V��K�!3�"��7.J�v�9oN7Ru.�Gl�uk`��v�2+�:r��H�ɡݻL�WO[b7{F��r�q[g���p��n�<3�-������\�%��&s`Վɹ{�C2k����\����B�%�1,�uI{�4�M>�1�՛�E[�7Q:"1��� t*k�f�{C�M�sh����W��s]��
�܀��Ÿ�I��wVP��U��c:��{Q��6{��iwd�7c��U���mc{�+�r�m�nU� 	nnh�w��֚���RԦ<jK���~Ve�a�6kFn� _	���t�Ie��P��y�ed4��Y��I��Ա\�������Z��ݢl;ٕpR��s`v�pe�f��M5IQ��:>.�U�V���KP"�Д)W�r��93Z L�y&8�#������=�r�h+H]�˖�S�!c+�i^���Ӛ:Y�Lt���˵KV�i%�gF�s��[9H@��L��sxui"_(Z���uּ����6��$Y4F��mo+�Q��� =��{� ��b�����d�k���5���v����g�+g����֫ ��8{����6���_Ӳ�k�M!iZ5�f���S�T�F�m����8G���ԙָ^�5*����5�:��p�5E^��r	&>T��F�q�#�̃zb��@�F0	�C,����t��mU��]`�$+z��-v(��m�^��w�4�@���g;u��j�����sP!)s��̾Ɔ]��3(�Yǅ���>ꛂ�[�,�5�0��E5�����|��E�:��MV4��k���⭰�2.�^���x������[`(X����]`jÛ�N��ū��W��J�D���@�5(V�)����-�;2Xe��K����(�t5o�|�$��pB�u4�Tv
AP�J����j��0�%�++���F]u
�&.���JQ�"���,�-aV�3V��b�$�L��5��է�a����SF�˾����w�5,y��d�<2��i�vH��=CV�����R[քKU�7���9�.0z�j�2:m%o��u�l�j�k�^>L�|�%��,���v���L��6�2����SK�F}gA�AiP-�쒹A��B�-��M�:��5�ю,gw��z��1u��r�q��j�ƹ���֢�7	D�9]��1�j�]@,f���ۦn
f�k�e�5�%sjS�oE5�Cq�]ˑ�5�e
����bC�/l�8�(Q|�fԎ���f]��tM4�=�qQ��#�/9�I�圯�u�4�3[�AC�|;b%���j݉Fck�n�S��$ɴ�NNb�x���}�s�r.�wv��DS�
�%sVdTrܡE����U2�X�
-h���V"�QF"���ATcT�Dm�j-��E1*��be(���($QrԈ�4�TQ�����Qբ�Z�YQTLi��Ib�j�AW5q�ը:�lE�Z������X�*���*���X[P���Y�Kl�Pb(��e���)KKF�iT���Ur�."ʈ�fbj��H��Ymt�e�hi���X��0�b�2��-���L����1Q�W-հQV ��1�+kb��M5��*�b�eh�-A�R�TUA�)R�Z+Z(%B��TA[b�F��f�H墅j
e�QI��TD-b�����DDUQr�3����me�V�((։iF����Ks(V����e1(�iQA�J���e��hV�(k3p2���+c[��%y0t�R�Κq�[�"�Gg"�y�g+�z�@��b�S�����1��I��nT����E��u@�1�F�sA<dˀ����`p�U��i��uKu���ګ&ûe������0Ɠp�(l6�N3�޺�pwe[���g�Y���Fe���a�G5ц�]R5�X�j`�r>�Z�r��;_��*Ʈ�F������r���]�	�+�X�+͎�L:�J��ǧ�Kh���}��<Y���xH�G
��\��ǕRn���Ǖ�$��6�33b�ju��j0]���Ʋqld��yɟrگ$S4д��,��«�"�XB)�D���TKy�jd�R[;S���?J� � N;��K�U�ׂ��.��p�^nx�F-��a;&9����W���4��ǹ���\��1U~:�_V��;�t%�ל�W3jWN{Q]J�u��ʺC],[��'��Ӯ�**�6&y)zlG	�ʅ"��T�Ž��^e��Ql���V:���6����5�E������:�٬Ӑ껣3j��x�`8V*��lـ��.�"�N���.xd/]��K�� `Ř:����ز��4莌�ѷ��ߠ�-���>LߢT����Ue����k��혶�2�����ޝB,�HV��7�[������P,���jKn�R�XL\ᝥ!�(�p�U6b���	$Ը^�mR7���&f�s���t�%���
�>jd�rh�N�b��~ܹ�e�7��ul�O29�AgK��^c˝��ɦ�� ��ǩ�98�9��f{f�M3^_}@O�����fw��n�t�zwg�9�O�Xk�<5<j��0��z�1��m茁�����D�o�G�m+�P^��7��y�F�Uì�#�5�#F@�:)̑«������pv��!T| [��4K0�S�1\ɕpe�2������M>�a��|��Ӟ���qu�W��ᗪ��-�/ß^�h�쨸m� X�옴}���7��7涴E�ʞ7��x�:�{����^<�'o=m�)��:cB%q�R.�##���])�eaМT�������ù��
�:.�~c���6���à������]2�z�U��(鄶d!>�1B��q�}s�s��X�;y*�۬��'�>D��Q�#�/%�p."���(�&�W5'[�\*�K��4�s���p�㧗tQ�j -$)�i�L�d@�l
��.�l$�J9Y�\q��9l0��5]%FwQ:�Yޤ��/AW���UQ�w��DXi�Itr��:.�E׶]�$r{۹�A[8ƕv��/O��cfV�8���y��v��)���yT��9m,F_Q.� ���sq�4]����I�TU�ӊ�y�;���dxw�5���<�9PEE��7��
����R0�
�yIA�t�H�f��{q��7���tu�upw2���^���9-Ҹ��չ0�!f��rE>|�B}]����)�� 8.P� Zk�SwJ��KOsu4��MҪS"��2|��S�!�n*��_J�U���^��.<9�a^za�c���TÜ3 N��Ϟ�ku�.VIȱ�m�@J]��⬱�ukf�#0Z68W���t:�����Hwc������3-����2�򎛼�@Z4 �0��)��?�!㲑���vh��\���:���v���<#қȀ5Wt���+�j��C((��|m�t\P�vr)Nז�^C͂��2]��ؒgLC�-u�R<��/?-�0p�PU�X�����Ýۇ����[ZM�Ǻ2�Gy�̫��T͜����>��+q��W�����]�=S�3[CՁl1�4��DW�g�i9vk�h����L~O"B1l�BR����TdH�ctt��>7[��L��k���sà��/�*mLD'���Mf����zv�mD�Ѓw�yh��"��u��;.g]�M[��.�|�vV��v�^�}v���+�I6ڮ%V�m`]u�+�z*}s��Y��MovQ�*0hgYr-�_ZKת(��J�`�|s�U�`�0d�¿Y�f�J�
��!��t �ug���s��yƉ;R%��_��h����	d����!�:�-�+�ć�}��sw����ҽ�\�`e��<���;�Lګ�o(��ƸYdM��¦g���Z([|#p�bH��.@{5Y|#q�6'2Z6:��c3ϕ�	b:��v��Ų��)T�����9�|��Y܎�.*}�נX�G�͉��\xj��ꍟ`��|1��)uՎ��K��j��N�j��@��8�MR���;R��+t�@��ɏ�g3���,�z���X���r��`$L?GtH�72+r� hd��Ƅ��x��4�C}S�yǲݩ���ڗR��&�j��ג�ȐF�8jC+���Ej�b��YF��Qv�F�&���]���}�Zn�� C i�ˠ���T�B�f���ܩI^>���SקY*���ܠ�;pR���t��8�K��� 5R��
 ��m������b�<�`A<�S[շN�(5uR%n�g	�u�-,��FSF�n3��e^M2%7$��T���+T�eݥ�ج���3k�x�ۨ�����欙6�R�ꕹS��;�Qp79�}�s�X��7)r�0����fn��V���5d˅��2&�/_[���W!��o�Ѩ*�+����f��c*�tDK�A\�+i�Ƀd��uպ	e��3���c6��)]7e�I�����HɆ�K6�]�N4���-|�<Ʌ�f-V�q5����gv��LfXpN#b ��,q6�ٟK�MC4%�ldװ_�G6�'�Q���`�Uy��JM��xB����@�( �����{m0�[@(��ݗ-W{x��U�~�zh��vi-��v�
��x�<��Ǜ�a��컬j&����6\>�x0x��N�yX���L��XO	�X�ltbV%�&���F���ն&��(p�c�W2A��TGJ�,V<�b��pګ
�ɆĵЏ�{�pk<w~O�;gH�C�L�aC.e|n2���6��%��+N�,���B8E#*%�e{����𺽐x���p9ʨ�&, �#�2�$F_uh����P��A�A�bB�����b���HX~��H\yꨆM���� ގ��\<k�m�uv�l�ѧٲ�hԍDjE��=��"�+V����p{%[�*����=1E@cӼD e�dtͨ!h��G���WQ]����ĕF�n�%}�o�nr��z@Nø����R���6�V�G�)b�/�u�m�j�68f�ĹfFb��oJ��f�,�H�]c#<�sE��y�p��a�~�WC��U�9/):K�_it:��cl�9�(ۉ�|k���VF����͂()*MCQ 4oӵ@y^ω�Z�u���ǐ��v�%�ro�DȚ/��>����PzPg���`'sQNjx �f�T�,F*�9�Cz���+�Oڴd����x])�(\>l�66� \J�s0.zuMn�ܺ��
�$H&�-�pDu��*4���D�̙9	:�*}u��lƌ�W����N^>ͩ�tC��>cڧ�s��Vn�O�*�.�Y)���V⃀�t� .j������O�u~H��r1����οm���_��Wz�1�k��FUNr�Ը�)w8��oS�WOa�|f4T=�B�`�������Ŏ�;����*��m���� w{�g)X OV��H�t	��p+f��9A�yuW�;x�r�W�6_ܵ���0+n�;����g\��!�nR�V&��M�[Z"��*x�1��	^��	�s�Y�:�:�\�I���s��t�9�ӭ{�Vk��D%����|��-�A��>h��N<әŕ�2�@�7,rW����+���8��sù%ܰ�Yˈ����k���n�n�g��Z�����7�����i�(���7�6��ٹG�+�?ը*��ZZ��9��H�Ӭ��u&i��C��J�l#��,S��jN/%h��z`�.A�0�,�!��˯n��e�
iz�72DU��\L���9�n*����2a��K$�.��ˀ��`IiOa��&�O`�c�\�Hiߠp6��5�
��T-V��_0G'������R�|`�kt�cY�f��yl��n�y5��?��:,C�l�8ի���J��
�u�j��r�����Ys�p<a����;���"_����r0ջWp��f6��l����W6��YO�#,[�(�0rxAK�w����W:7*a�F���D-ڿ���:�{�eZ�`]�C�#C�z�yLH�;DA�u2&e3�a^�1v㇕0׬�c&gz�ޭ+��T�:� "��(!�ڵ�B���ug�y�*�^����-R��B�I4��7E�����ׁ�� _���2`��Iڰ�D;��z]��#+�}~�&�@R�����^&xC����|�Ǳ�o.��K"\��D.�=���蒃(6�E&�5�SP��ouɌgo������hz�k�^c�%4�΋�[j,;�8e>��R8�<���F�9`Y:�F��EYۼJ�+�b�A��V����J�]۰�-;5��Luy�(ׇ�5N��Yd:�+���ey��LJ�V�֫0��o�{�����S<'b�d�5e�;钦)mS�9�����h��1"���C�x�"p��q3��7��]ܨ�)V�y8+�:n:���D:,(�{G�0��Y��}u�O(l��H�j��@�>��"��s' n�o#"Ԁ��i�>��@�F-�h�*�]�L~y�,�\�uv��NW����_7��Y��FP��f��P#�l�b�u�����Yܲ:�n����|��^��1�p�"���`���D��Gu�Bſ�})�]
9@G��y��q�MɊ�3�ܳ��
;���ʚ�o(���A�-�1�MXT��v��m��ݷf�خ�a�*�f¨ԭ��ن7M��숹�Qr�7�&�)T	=���H`��εUKt���gp�}��Hy���:)ǫ6��@b�Θ�|fʘ1���c�'<��*���y�>�K�)���v}dOW
q�ܔ݊�B��^��~�O���a8\P/LE�(X�xK�'Q�nt*�l��q&�uҨ�9l�+���[32��%ge�����[o^�/�i���-�0�*�.s�Z�^�wy{Da�_J��>����Ӆ.�N�Vr��6MT�j���?ۋ&y�ph�N��p.�R�5��0�Mn?l.�v��i2���@�(Б�c����8K�gV���Vl��Gf������.;�|w^�ܝ�[������Ӣ�Y��ԇDƥU#(�U��ѫ��Ƅ��=&��T�PU��#y�ܹ��MoAy}�Q�{r��n�FD!ԆT���2޲1�<ѭ��U8�;�0+#�oe�k������=T��rق�6��:sB��>]>f����T��yk�0=��j����U��Tx5���Vz��H�wmeN2YP!� l5t䋉���&D,;ӫ�H��N�*p:7X�B��c�Z`3��犚m��P�AlcN��Z��v���+KJ����ػ2��:*}�8�R�Qc�+������x��ꆢx[N���#ب�QA��4�\��ڇ�1�aa�8p&`�m +�Yw�L��j�6�����t}�3v'�Io�%�x+@��A���:!UOV���DmB�"H����8�.�Ĵ ?nM�ne	�U��4!�}Dn磓"����b;oFk<N:���)��fp0�cH��D��y��|�e�b1ǵ������ɱa�UB�Ē]F;œfZH�#pc�=�[���{�H�Av�i*ͧ&�Ȧr�����3os�V�����-�;x�u*�i"�*�����h6��|y���0����GC]+��N��F��7�0�஺��+W:C�]5�*0�j�\̼,e��8O���(�I�v�iۣ���{4Pԗ��f���'���}��$��P�-�N��-AQˌk�U��t�R�a��m�J���iuՖ��"C�O�V���s��.�T\����1LZ��Xv����B���-qY��Sk;A�G��<���
s���b9= a�X&�䥷t��簢������S�Z,������,)ĥ��i�wPD"T��5F�'j��|�`]`�Y�`�n�`�ǱR�4�Ai�l.�^'
��A��nvDZL�D�6 O� ':y�f3��C���窻v���9�s�ؔ3:Y/��B���d�17� -����Sj0�QY�]K�]a�&�����f��1(�u����}���L�+��)9���`�����V��*϶�& ���]���=��%�
�i�5)�"������zX�>��K}aэ
4���MФ���GXҸ�.�t ��ě燉��U�1*��-ĀnEYh��B���:
��Nf+R�]��v]e�kPa�4��)��R˷�Xk��<�Ǽ�/�c%<5��*�d����|��p^GHn���7V�V9١d�Y��^�h<s4��^����eN�z���Xə7���bl4��ցb�59�ɯQ�C�X�Wx�qqO��?&�~���u�g"��;����$=s�扻ч%i���˒c�d��"J�o�����U0�c��_P5�mwwR˻q�wS�F��T�����X�ҷK�Z�l�l;4k&Q����NM<��z���=otgRw[�hT���M�����%���N˾hQJVlv_JA�lCwq��B�y��ycw9�IaL�^ت�v�U~��]]�|���x�1o`
�u)�~��5�b���2$�k�� �f����.�&�G�ff�/�b�@�4E��z�Kr��l��yu��NOn��P�:�a榧����1�+���5�A5+��J#N�U��j<��(�c�<���.�X�c�V$��v]���CUA#�uhk����:R+��مJ8���:�+rڳ\��@r�t��ԑ�v�)L��-_fh�J��B�ַiwaf�� -��V�p)�^�=�`��=31��X�C�Թ�	Y;k�b:Ͳ1�;�Ո�u��SXw�'WT��RgYXqա��U�Xz�ЦG�B �ͭ�����P�*��F��.i����Ϥ��{"}�v�7 ���̠M����H"�n�N�+�k�B���!a!��E4��{�!GAڐ9��>�pCh�s�M��mj�: �2�	!<�/�+.��i3�&F��L��c���v��YS�v���{0jE9�I��&	��VP��,\�4?�X�R31�����p�� {w�W��������F�WKn�"тKY��C��<OI��Xp3���b��4�q�3J畑��H���+ץ����}4��ba}w�L�YY����N�1��EP�z��.�t�h��W7��G��œ�g��W"�u����I�J�1R@F�V.��s5,�$-,��h�<k��C���mҔ9tM�v,Z��:]�l��Ojr� )/Ne���uY�`wR~�+���4�M�;;V]�a��^�q���75<:�3=(���IQق�K�f8�D��TH�R��k@����z�Z�h���
�JŢ��,C<@p�	�Ab�U����*`嫅�JU����E\�*5
#�Ѫ��DPk)R�ҵ�V�QU�6�kQ�##Z�Z���ڣkF����Fѥ�`�RҍR��k*Q�tኖ�j��ۖ�Z��2�+j�U��V�E��J�ڃM&8j4���TZ����F���)��5��8P�-[m,m�U��Kmm���Q
R�h��Kkt���ڥnL�ckB�h�n�X�����iF����VԌ�h�-n��V�)J���4m��F�V�fC-�[m
-V�ڋ2ᒥ�X�m*�3.D�Ze�QpU2�*���Z�ƙh�s-�V�V)iE����ZҊU*��h�h#munR��(��6-SNaJ��ŭAV�kh��(���k�K?��o����\�{3�Ȯ�=.�F/�(R��j��Ôw.�)�]���6���/p�5��<�y�,d�'[խnP��U�r�v	-�W������~���R����t�u���TmA�� �Nwr���С��	�^�0�Cڤ)��;�X��I�Iҹ^������y�+)w���Y4��q)��g�<�;�F������'��K�~� 4� ��e>o��xܭ�E򾚺�zi��.�	� `��c��U�'KT�5��/�򧊑ؠ�Œ�����R��j�ʯ6=)ϱR��q�9(��Y�r�L�y�hY��Mܼ#���߽�ˊ=x7�Y��֨��u3�q��,��&2��/��=wR��]?

`bph�y���M���sR�䯎P���>�d����u�(u�/�ՙ1�Ñg�N��׋R�WV��Csf(8�-�܆�uup<҇��E�)USz�+. i�|5��N��s5oQ2%��ҳK���<�̈́���{��tX�����Pի���A�����	Ҥ�_H�5�fo ]d���Ȳ�TEmhW�Ǯ�pB��P|yV{7�*}T�v�U�Q=Ǉ(��q��+�#��h[T�v&f�G:��v`3o5�LǙĢG9p螞2��� �O#��r0q�Zʩ+B�YrJ�샋FK�p�z��ٻmE	��V��Aw�7 ����N���`�Z]�f+;��H9��nMrq���L��9,u�����k ���s�U��h�J�D��^�}jR��n�kP��E��n���ZH����) 9�u�<��:s��@gn+'���R.�d�1`O��"��D�x���{u���΋E՞甫�Foc�3��󇳯�PئpD�MP�n�@U O��d�zzC=h!���e=�^�Q1!�P������|������[f��hpp=+�`�heL�"S^��c����*��+qOt�է�ۥ8�t>��CI�و>�u
�:d����M��(h����h�Y�4�rM����i�ʼ�K���N�rlM��,t��7�hzb7*�4���C���\:�|6:���~Yջ�^��ɩ�\cI{���戥�i7�Zߝ1����4� b1l�C�a��y;]���z�S��qJ�<|ϡR���P�_@X�W��|������4�}/yH�̀�vP�M��ճB4,�:vN��/�.j;f�3�Q=?{��`��yݰf�ݚ͛��r�_H�z�m+;.�s�9`��+���镘Vm�����t�S�,^&/9z���=�Z�߫RW$8MH�c��j=��iT2��T�'�V���哻kq�Ą�����t�{![���du<���Rݴ6��KBB���	�	��17]w��see�����A�Kz,r0Tq����#YX�3�y�J��~ٰ�5+c4���ܱ唱lN�̣M�&��N;&��D�u|�v�m�;��Y��/�k��b�p�Ή\{=����I�R��3b�͓]�� ���0�}<��̸]�(���j�#v+Y����`�W�r%�O������Zv���fܿ����#�!��Ut~�|�U�N�X'�!�B}��0����q�&�Q=�`�P��{o��l؇��;TE�xd]z����@�z2���
��1���[(�7�fWV��f뭔��0���| Sv�EʪrEĺ��n}����Yj�Sg��su��q����JE�
�^z�b͞�<pJ�� W�2ɸ�@1)ԩ�.��<��u�]x�w���Eʜ�BqN],b�"4@f3ܝ�"T��le�YG\�f��WO^<�FJ�8�?f�Nm�б~��5E�b/T�3^�A׺n��#L9,Iދq֦߲[�{����(���Af�ݣ�g�b�I��F�m���ou5��"Q�64��Ё�upq=ֺ���}��n�(=�6z���sYg�(dW��˒�@iP���-���@v�Z�v�U��-��A�M�7���L����ϛs�]��JJ6���{{^�x8P�
��%z�Uٮ�6�g�h�ƀ�e�5W����[o��ɼ�;Kݪ�S��I�o+��'�_�Q
�ӣ�(N�]�994!@���<�j�����(0��7檘��lD�7��Df����^�)]�ʭ�j�0�g>�d�ӯR��l�nq�M	n�b��欁e���npF뺞<�p�&,:�x�>�o�����BⰐ�'�ҹK�*��k�e����yn܅R�{��\�e���I������S	.�+JB��{����_.޳fWhK���$V�����-��X��LX��%M�T�
��\m��� >;�)�|8_����v*؆��1M��SS\�LT��:��:�e���H_��$i�+ .�`��qR�u1˜���Y[��4r��!�o��X�nH��*P�s���b9�]B�#Ƴ0�-drSD��5�O�c�f@扆!��J^��]��V��IH��� �>�������7�j�_p"6Sܵ��p�W��p��=�s���6�C���*��+�ȫ��P��T�E�?���f��kZ�OO<��fQ��x�Rq���U������apQ}-���]�6�yUh�$���E���z��U��6T4\����!w���D��༂§��(�(���Kg u���L� �Mp��E�k���ܐ �}QR�۠�f
y��)p�U����%k����T��̝Y�;����t�n�ޖd;�G��E��
5�㎈��}�Y�xx[����|�78�
*�(l>��p� T'υdNji.�A�ZsP���3	V���[[��F���C��i�L�4�}�lI?1��_��A:�ߟ�Du��;�O��X&Q��Fk$Wi2g�o==���l�1������g��j��P�I:*�9b�y빝Hʈ�0����\ݥ��h�P*�\v棶h �Cr��^z�(6x������dV�ܪ�$�;������ۨ�l39�,���@OJ�Ą)}��1R����x�[��]�Ua��g��3͎��bB�6�xʫ��kB����k���#���Z�gk/�{ۗw<8]�U}%�tUҸ����2�U̱�6�!a�h�^�5k-���}����OP��Ν'.ԕj�+:j�nQ��;(��':�6�y�a��E���9��+�.U�I��+&�v*��<tB�\�B6%`����
r��9��s��L�F���]����"�V55D:v��WR<n�[�{���*��7s�x+���:0,%x���TB�������<�<����ʇ�S��(laL��w����/���0Hr�( ��U4�ՙʿYԦ�:�s���ntia���}��~��'P��QM۸|.H����;�H<��+��U�WDqJ�6�\	��ݻ�;�/�p���ON�Uj��V'j:��qc�N�%&%��jh�TA�(�쵂���[�0��p z�w�OvPU�7���Ns��#ʯ}\�6�ޥC�K�=�$2��§�g��T&Z���ЬU�#���]v��7��+��ͮ%�1`O��"(��@E�q�����y�MS՞뼽�#�t��m�.z����
�"W*0�����"�C��gs�f��׽!�@յ��oZ���sl�����MFo���F��+�v��b���m��D��դd�ѧ�`5��5 �{_�����S�P�:d���.��bF��hR�S&����7-,��Ir��d8ԥ'�o3ﺖ��N��(*����|�9m'�'�f��z�r�/���oc̕����NE�ޞ{q�-���N��E��O��Ch�u�&'nX�t�^>�H���Sɢ���=lI�1�;�@�v�f��!�<W�d�_���]mXve�d���>SC��OJ�Ӂݷ�i�y���ܳ4:�Y"�n@�6�H�Gt�uN7f��R���^ ֬��D���.��޾:��䱱�U���x���L'N����0eJ�b�2������s���u9��nm���a�sT����3�WCizf���ݳRbU���R�7������c��OX�o}�Ղ3�{驎��Z}��M���W9���U��!:�+�X�ii8�f��x?��%s��~ٰ�5+c26a��m�K�ح��\��5h&�7~����x��h�E���c)%�/����!�*�(d����� q��!����p��7�e9o&�ކ�?�T8�_�q�y/P��j��Au�.8�&;2�uA�7Om��Hp��.���\�C��:�3S�2+r� ��`�9t��\�c�[\�oLi�jB8�7ٙ5؇U��*�Eq����82i��"A=��e` r7;$t��a�&{�n(Ϥћ�ܼ��ҡ��]��AZ�^��p�3[�|��\{��X�Ŏl��*�~��h�����e�<��\�-�p��	�V�G9��:��n����9w��	��>ݡx��B�M=��i�Zn�V��&|t�b}  �3�Y�̏okglJwf�������*��L�@��(��Eŷ�|�Z���]��Vj�):��z9݋��C�#���ʕ�����ep��$�'i��v���8C�[9U��zS0l�`	�6��]*�$<<�D��ͩ �mE�^R��q�cp��|i����>� B�Fˮ����6C,d� -e9"����p]�Y���e���pL���;t�l�_�9�l�ؔ�M�\�'9*hd2�)▹���w�f�QӐY�`�!��:�"�ݜ����������υ�DT�ƣ3(�c�}�}�PtѿUf63ݾS�����P���=�S��l�L���1�bC�>��ےh 甲�_.�����5j�*���d�yX.x�!i:t}�t�WBan��EV��������f��j����y�DW���<pX�<����bi�������ؾ��(�f�
���!�0�y�M�
��z��>�XO n�o|���bsׇ}o.)�Z{����m�(W��ɐ�ǃQҹK�򡊄k�g!���U_g.��z����O�֓P�K8����t�w�6�K��es,qE:^�b;��Vf����S����&�x�Z�"T�m�o�s<��!�ժ�蠪Ƴ�b��z{���*�!���?���+���k�Ѿ#��N��c^m�(کP¥q�f, YH�.�C<$C��/U����H��lOi�,!��Ul��ӂ����9��P�ʁQJ��O�M��Ӕ\Ƚ�ꇊ�b��F���� |.c�0T�;����ը��F���@z��+o�<&�~<��ק,�&���_R�Q���(uZͫ�����Vk�j-͂+�I(�5F�w(��ҮQ	�յ劶�*��t�_�| �^nvz�ˉ�\qƋ�4�w�ʮ���H�C��
�*�)6#Qx{���d����4"7O'o|��OA-�=������~J���2��S�k:}^Y(�t�������Pw�&�n���y�|�7Eɢ�3hwϮ��V j�H�v����6���!�60�%_n����\Z�P;k��Vhp�2Q�����đ����u�,��ߟ�ϩz<,�<=Ս �����ҭp�KĠ�ӣ��`��2�q�B��1L�24M7Qb�I'ED9�r�����Oi�������
�(r�� G�y�tw��>��ԋ{L���fm0��Ǭu�?]�T����9I��g`�>����V+A��ݜ�Pʃ��am醷��]�DZ��ӻv�T�9��#بz�ݠ���&����r���U�����f���W�4�q��s��+gf*��a�5s�zyTv�l�1���(d�V�Nu@�I5��@�%��cF˪��HU�g�� F-�9����
�ĄS�R��E/�H�����f�c�;��C�ĺ7R�#!�'Ҝ���%�.�y�5�YL?�8�|k\˜K���ux���H�Q�R�J�/�q��+����*��X��(�O�7��3]�E]5�r(f����GFDL�7�a(מ*$�����Vԓ�E�׼�[��KgeK[� p��*ab�S;��=.ja�3�Ux�#�. s�����Igo��}�C�����)V`���`��[�{�M�����s�� E�95J�+��.�S�� e m*� tb�r<.���;�V��7^���9&׻�wR��^vrr��q�4����������,��k��)s�U�Ά�^�{`��:�u5�r�"ē϶�&"�3��ژ5Pno�2vH��Yq4ɟc<���N�"��_ҹ��ð̋��M���v�B�I˷b�_!z���DV��p��t٦�M�S^����|:��~�Gx���r��5�����u/fv)��)oFR�F"�4[��(<z:��,��r��r�o������q���� Q���=o�ͳ�}T&Ҳ��SlMָo�����Ы6w��>����S�.��V5�b[�Ž�3b��sc�8\ZՃ��Xw�]���K�\��v^*��cwt4j�RL]�n�-O��)ɫw,m�du�ӕ�l ��<���\��T��Y@1������û����u�Õ�Y5���RXj�}\�v�S�2\�wl]�U�:ד�9�!���UPup���(��#u\�A:h{x�^�����M�Ob㜎'Hr�[ő�m��tZ�JH=�h��sV�y��En�Ӭ��]�:������2�"�
�*�q��<x%rDh��T3*�2�f��V&mhT܆bKx�֝�
Mv�<���oL�ե"���5)u'��u�J�.n�'�;H�\�����6�q��mfy�T�;ĝ�r��u��<��j^�u;x�畅eu��b+Z�m]��k,by۽i]�Իq���:-��
鬍<��=���!��.��uX��޼��ܓC:Ι���<Q��'s�u��R̵�^��q�`����yIe(�23�ذ�#����ѹ�OM��ܝͣ����]���)�dV��
��`m��@�އ�@x.�eK���9gs&�q�^8��S]nj�R�Q�ѓ���AF�4�5/�J�
�4(�U�������=φn�p$s��j�ꥮp�LkW�J����Y�r�L����I�8��n"9:ܩx@�95G��Z�,�j"hS�I���p:�n�*`���� c�[7������[s�[n�MzNho%�t3kR���z0Y}Ãf
�6�oq���x:L���J|��u���$�k�����E�g���-&� ���V�n���.�����%������wP��n��d�(�A'Ҟ��[���#J[�/$�,��Nm����;	�otE�s3o��]��npWL���sXV��4�t*��N�
���c��W�v���U�-�	-():��3 J��*Ӵ��Y��e5v��+Ă� c��=/��/�Q�o1F���ۀ�D-�n�j��<5��)aJ��N��mւ�-5�gg1�P�sU屬�E�=AR$�\�Ÿ���P��+CǙ�v]���N��7+�rT��_<�:�V(��{�U		�d5IcWQ�-7���H�˶�C��u]����~�=y8�Ϟ�����[ö!�LN�f�AYf��uj��e�f�&��͢֍3��z�̣U\2:[����j$�Rn����d	��}~��9�ء|,��3��dS1s�f�OR
d�%
\Ilkq��#��U�9X�y}:�TwE�H��U�7���W[Ѣ�ˁu�ٗ}E;�Lƻq�Y z��������h[�b��e-�f��f����Z�m�f�Ɍ:��d��
D�sV�C�˶�*��D��|Rc/*P��+��[���8A��<��f������$_�[R�md�*1��}�b�L2�ض�U��I`��WMAL�F��%�F��R�2�e+mEkV���\��K�f.�,�J�EUA�b�0e�k(�J�S(���cX��r��Q̪���UQ�㕶�+m�QR���*ʢ�S0�ʋE�T�R�����ܭ��n\�[kj�V���aRԨ��\V,�X[V�Q�**+Pb�m�Zڢi����Ab(��M���)�(��-�U�Qb�UD���-�Ke��Iq�KeJ �,V����X�Q��3Y����F1X�V����Z�"� ������� ��IX�t�qEƋkKi�E&Z�*+(�Xc\E+iE�ʖ�PDb��KhT�%���AUTU�X��"�����:B�r���V��(7��d��<F._K��Q�FNЉ.��E�ݘ���f�[К}���\�G���M:p���sӻxm!B(D���x��=b��N����܁q����6�oP�.��n}��Оb'!��Y�t&D"D���	犬 T2(�)���1~�TI��Z&u�wF�qkpoR��5{1����u
�G��Y��1U йa�As�D�w����~���ZI�%�^��vn�o^݉c	ڍ������J����N��$`�</7cx=�K��cu���V��	�	;�0�rtBة�Xq6{�>�4=1��b�K��)����$�k��}p����$@���<���J)���TN*zX�B�����S�U��+��=��1xb������؞�Y'i���~K�J�W�Yb6V�L�H���T�����4�{xY�ǫJvu�X�b]��u��uh���γR`R0eC5Hz�����Nт�B��>����GMAK�
�'	Ff��˘��LM���3p���q��!�
�����28 d����@!qzhv�V�dl���ܱ
k��;���N׳�[��z�s�[y�GODՒ<�a�Q��`�ٴ�İ�ݷ𼼓��+���W�t�z=�R�����`A�?wJ��vF�sK�+'Ǳ���6����rμq[Ӟ�\2��Ձ��*)�d��[�:G���G�ç� �9(�-�]}����M4У�D����d��K���	'	G���+lR��Y�A&VX^��Wd㯣��Y�q�+�61��)�p"�z�f�YU5��J�kq�k���,��g&�[�ɶVv�"�q��V{]�1�����M53�J�μ�P�^��1D��W}^�i��.�y.�u3��ر�Zw��&?I���dp�d2���߲���WBj/��.u��{����o^�B�O]�\)�*��F�)�!� &�\�S%����]��xn.{\u+��4��w/��ׇ�	�=������z@�1��qp%�2� �sV�w!W;[x�e`�Hs�^&Du5��.\��8�3]�6���B�������5�/e��v�/bi����������.,CP}�)$�zt.�t>���N����!Bf�����n+��ĈTa:�Ɔ%�oF�HU��\��<1�aa�8p&`�Z�X���I4N�͑�8٭<��G�O�מ_�M7���O�TBN���]�U#�2�m{�ހ��.�۸{`�ьZ�����ڐ-7�`��S읫n���8�$[��)�t�G���Ͻ�����npt
O�⫋�7}jTw����d�g�N#t��e�V�r-����n3u	��[u��>r��7�X���{݉��K���Dz#���ϙ�V�*��8յ}ŀ%�f���c!�؉�y�Dk}�!f�6ދ�jZ�{�m��q[|߄\Q�Ƣ0�1M����\
��4�!��@�ojt�Du�=�^c����yI�-uD��r}XP�ia��[W�,�^RL��9]kR䫱��RP���v�窠q�<�J�;�c$ؙ��u��8�g���݋���oɴ��2���fFS]�[�-������
t�B-�'���@JUFb�.y��A_]�~�\<�Ѻ���ʲ	K���8]<"������Ul��8)�5]�ג�:V��y9���fC7���|�nz�J����t��4�J� ,?��(\���'l����E��t�v�l�b�e��#8^�	�RR��8#�ݘ[��|R�P8�4����]t5�pEF�u8w׶�:[y"e���UΏY�R�������ڴS&ƇGWY��w�.�ʬP{M��`��#/�\N�D\���#	��Q�P�f
o/�K��^'�q
�N���򅻺 Q�J60���,d�V�dXSӎ��p�dO��9�wc���&�]�ih7'Ay�V<s��*�J�f�]t�6 E,}�-/�����EJ�_(m��2���j6�<P���\x�NS|��i����ɝ��\�ʺ����{����N�����eT׫��>��P��>TgԼ���F���J"���A�\����Jt�&�Kn�����2d�4���*}tЫ SX�D�R��&\���~��Ș&���
�K����)�u��ԓ/��҄��%��}@O־��deϦ>�<&��L+���O.��7'q>�k������#.�\����9�;8!@,þ3-�a��f���P?j$���t�e��dXb�V oE���;c�4�\��7=�Bs��(x��'<�>�[�Iw����zϑ0��\�
��Qxl7�@�Q��}����+�b��pF��M�s���&z����-�=tn�ϑ��r})ǎ��)����@��E+�t��7�5���V��i��ܩ	�u�� �z��פ�?C�ET�:���; ��H�BUMt�z���qWg�u�y�64:�*bn!���4r��
�O�x���TB������si'S r���k+�W(��7�ɦa���
}i\X�����'p�ߝ]CjJ0����/�lZ��&�	����Hׂ�x~׵��@�<A���j�S[�l)����P�KE��M�J���ƽ�6r.;�9L��ꝣ���-[�&Y怎�e�9�O��ƱЮ�Z��'+��6�*�����*gM�,3{ &��ʀ�����1���DDz=:���ڼ� ��@Viګ���1��H�?�P����R=6��<s��t�g�̎���Ɍ��]��7`��X<@T�
�b���%�G%�H��/���{~wֹK��-@��W��}W���C4�A�]�&{"oМӓ�~�B�bx!��"I�7g�Ýҷ�����f��D��Q��n��=j��1�)�$�����Ww�W�*E��X�Y�U�Gt�F�CK��y�ј�'��1�*���#��fl'��D���7�Q����z�x�&�e0F�ToѴ&x�'�ʀO
� 0$�p��G��ڸ ���RwG�y��kG��x�������P��Η�hKCh	z��Q3M����h�h����Kx�Y�s��W[Lو�s�d���ڧNz+d;(���Y���yT��7*ŷ931!50I�هQ��B�T�8�;(2���n��ۆ]�3'r5o c2g���<΅y���C�tߝI(�M����O:a� /�Պ�ݔNM^լ{�܍�κ女V�'�X{V���6���E���+ۤ6�PWWP��ԟf
���R�@i,Һ��V�r�H&��V��ڵ+��j�\2��\��[��b�����0Ҝ���#r�#"f�gN����՝�"�Vf:6�K��Ǽ�Gͮ�9#�o��a霟ݬN��Yչ3��Lw-5(�`�Y���	h�w,)@
Ý�b���������mmҰ��H�x�c��@�Ų��))zSSb{\�a:v�꽕
d!;V���{����b�3�Я<Hx<�]U��P7.��-���r�pþg*Fb]H4�n��jh��������1��9X�N�=�T��S�_tAX����U���{dBa�\�*V+�ZU^�8A���xh(�e��;O�r�`ש[��n�nX���.�=�@
;v�.`ի��NQ�~�I�&�@S[}L$�v���0E�˴�q��\�{��MY�WP*ο�S�!�4zc}�ґ�9�8�,� lT�!c����ӗ!k˂��y��>��~-1M��k=��ڹ����LW�D���Ҳ�*��3��D]�b/��';WE�����*�L;��cɝ�O �.���2�D2���ĩ3���汧�Z�#�p�s*e�Dz�u����0�kهSu\l�H�ŀwR2)U9#2�p2*��1�Y�����f�����PFg_�?Jo>�d���&r\�j���ަ�i�H�呼j�\���Y-�w�CS��M��)u�����	fq˱�q�����յ;Y�:�� 14�e��$�B�}���ޏj�ɷ�eT�L�QvEz] �W��
����Ĺ��oاC���6�]Ȋ��.}��:�UYn^��EJH��6_�'f{����/r�)$�z���Ԭ,FB6�R
X��8��v�;�Os�z͇�$D��RUǛ�m
�bٓ�]������c�hf0��*(�xo9�[u�L�[�+�G��Pg��c����͌���9p�U���
��Z�{�+^n�7Sո�a�
u�c� k4�G:�8d>�50_���7hm0Gu�H�V����gh�N����#Q��7���U���|�b�}��t���ݽSv�Wf���{R��6N�y+'���x���&���Ȼ��H��8�<��Vi�����k��v�����|�5d�x���c�]_}Q�	��%���{���Aa�P��L�Ă��;��%O�;�i�Cc�1<9�O��LA|;�������,�|��8���I�i�,g���A~N����h)�J~����������d����'R�x�|N{�m'�W�<~ߛ=Lx��,=k�J��{�7�L~M!���x�m'9�jx�_�n �Ь
��jì��=_���>h�fgBL�Ώ����_�P��1&Щ^k]C�<2�P>J�RW��>5̅@�T?!���<`T�B�e<d��`V|{��X��.$�P�q��I����c��#��+v+�&{v&P�"��JY�h��,����_�vJ�79� #�(9�D!��r@�/���ȹۨ�uH�<P�Xi�;ƕ��ݮ�c=$�d��wn�l�<1d�擒�}y�A���ҏIbG3K��R�$j���:���ޛ���]�����g}�~��~k����'ɴ��"Lxʇ�Y6�q������(x� �v}a�m��1���2k��u�x{�4��g��q�xɤ%g������/��
���aXW�����T������	��n �<EF	u�@�+%Cf{��7�!]0���q�C��u=?]>�*��5C�?;H,�1Ru?&2~�}���q1�=C�A}d�14�|aX�o�o#���qv9 ��;�<���G���}�++�u&x��(i"��7�jJ��I��'�HVi�Zb�S���lI��:�ɧ�AO�CY+�XϳL�%��I�<���9�9_}��Kv�.���=	��7��<H.�y��h)�Vw9�}w&2����$����C~oz���P4Z/�|eH�}�8�:�_����i�P�7>���`bN���t&U5�r]�����G�{�'G��ӳ�H�C�u�<�w�'���R���㴂��m��SI����\�6�T8��l�ă��!��&�Pĩ���<f��6�3�l�����\�'?�����@�����j[w��Ty�@���aؘ�vɈ�w9C�4�f�s'P�
½�� �P�y��H,�J��d����+�xo�M���sVOf�71�PXy=���=q ��=��s������qRz�La��'��1��j� �d�f���l+�g�c1��&0�s�d�&�++��)��B��_���x��g��g���+4͇�@�{�6���ɹ���ޣ��u�����Rz�zf��?'��A�%|B��Y==��K�&:}v�^0Oo�z�$�x�q8�@��sn�k6Ρ�h�Ԯ��;��,{A�,�ج��kgwq����(J�P����RWg5�G�O8�s���I��1���_�=�AH�C���g*T����>$��X�a�u4��s���Dǈ��AR�2�6��7�{_³r�d��A�ͧa�xzʂ��P7;�����Lf!���R���c5�}��XjM��I��& s��4ì+��?�qJ�_m���LAH��+�}���#�G�w)��A5[�E��oz������ê$�n��dNN׋�C���.�:���,=��ӧwe9S�&,]��^�u�|���OJ��В��jb�&�����_mn��!b���ą�Ӷ�H��#k��o��.R�*�+u�/�]��T��t�#�DD{�}/3y�Y����"(D!�=S�1���>M!�������PY���z�!�bC��2z��N'������cNkz�$l�o�Av°8��Rm�g�1��:��Y_��}~��Ӡ���'��7t���"�z�EAC��ǩ�& �]����;gY+4�s�&�=J�0�9��?0*O���ߵ�%~`T��E���Xv���3�K�OƯi񁫘��bH�1?{�:4�D�/�u���y E�Xz�8���q�'ShJ�Į����&Ь������>2����A�jI]'�L@�+�y��L��!�i�4�2�'�7�h))����^���.������u�̅7�7ڐY�%N������xn�O}�d�~����eC�},8�yf�9��x���Xy�?$�1���{���Az��1�����E�ֳ�lE�ǽ"<����]@���y�R.��a^:d��3i8�aXW��:���P��Î����O̟&v��ۧ�g��i=<��4���/�qğ3�>��4ʒ�N���{�h��D�/���t����;��9�US=���� �a�<M �aP5��钲��b�'++�~;��OT*M�`/�LAa�T�'�%O�b�S�y�]�`T�?32|��ȇ�Ov�X�?7�b&o令Z��'�".�/ԩ�߰2��1���ǉ�At��w�kt1:�${��
q
ϼ�t����<�~�bJ���8i�������1�D DC>���{dQ;{��9=z��b��L@����I^�1-��+?2f_��{��
E��p�Ă�2w��<��H-x���:�M0ߺ�i�
�ʆ��sF�ԃ�{�����@ �^�r1��sw���iC����1�𡤂񇩳TY�R,5��!���& q+��]!�5���
¡��6��

E73�m�_0+*y5�Cmd�g�O;�4����{�<؏��&>���}\��oN�����+�gM�a�Rq�q���CL��b����i �d�1�>������6aԨ.�T�}g]2VT�ԟ��R�VWs���LIP�k��H/S1�K�e��������ow���?v��\��3�Ϥb�݊&�lN5h
ٽ{T��ʢ�1�;�sB��{���\�]�b9q�]d�)kN	,�Pow.VP������.�9Ý�Mm������HZ滏�q��AQ�w�̊�e�,n�[�k���ϥ��HI=��{����˟��Lf�f�f�*䩯�������Xzn�?�>Lv����AH��W���q�S���4�^!��3T������߶i����`m������<�����]f>ok�*<~��DD�"=�N%q
�I���3i�0�ɭ~��E�P��!�x�Y=7x�C�K���봝B��&eӿ߰��X��5ۤ�Ρ�11&<t�}^y��Z��>�x
)��W�����?;��Ya��4��d���Sg;����@�a�l�i��P�Wgs -I�1w�>CĂ����g�X��i'�]����i8�a���y�&�q
¥���^�w������

N�0>a�<~Ͳm!��Xw>�
ϙ�j��+��y��
ԟ���wVLf$�������bAtɳ~a�}C�����l*���4 ��c���Yǐ~�,{�x����(m䬕4{���8�T*x!P]�Y1��bN��3�}�d�=d�M��ޏY4���S��P�?&?���m"�ɾf�Ƥi���扼K�ջ�ј����CP�@@m'3x�~H������4��Xk����!�
��C���V
L���6�_̞s���*E������͟�W�q�����%��My��}ևFn����c<�w.���"��z�
��gf�	�n$u<�1'箐7<�:`W�>N&�g�:@���q�@�T��}�A�وq�ACO�$�:�y�?'�6�^3���
�����}�fJ����Dxz�I�T��N�u�@�+0�s[���+���
��fE��ǌ�f2bC�����&��O���e|d��4�íI���s�����u�,X}���[��z#��G��G�ɴ�<H/{����x�0<=�;�a�b�+� q�J��:��O>J��d��z�Vx�H��偉��1"����<��d���K���ݼ8�]�~"���z �ϴE<a�����ﻒ��_��f=jAgXh�0׶Lx�H/����>x�C��a4�j
}�`i�Z��\g��R����<B�R����k3��U�&&�3լ�M��b�,�����u7�ۭ��J�,�c$�X�E}�콕�6�r��;��a�0|�sZʫ[-K���I��Ķ��ѣ���͓!g;fܲ�Qw�.%U<�c�DU`�uz�V��v�"6m��e@�K�.�M�]�3'}:ĕ�`�mCY��cJ}t8�.J��p��Sۗ�8��Jk<���7��O�Q<lּs�C�*Kw�p�
6`cv�>��3� ��@+��A%�r��2Ao�T��lv.�_T�ћZАĴ	x1��+��i���5�|ͱ�;�,�Ef�|HrM��ںt\q�/��J�K~R�o����3U����Ζ��5�b������(]s	�ꩡ�`�p|����{�)w��;7�MIN&�pIٳ8\3Q���ܽ�Mԥ&s�-����O�d�%d�ݾ�~��Y�fpRr'����]�)A�s)��U�kw�p�P�YY�=��J��W��@�cv�ܢn�|�3q&ō4��K*�2���8p��xz�2��T,u"���2�޶;p)�u�:#�2�w����7d�������i�#�ܮ�	�<��ʵ7 �p��q�+��i;�2��T�&�0;�	
��5��V���ҳ9������i��u
����9��4�^��j�\���ƻ�=)�b�v�P��m��q�$u݋P7��6�]v�X��p��@�>�!Fl�7P6N��3���'T	uU��b]���c@ P4J=�]w1�ٯ�a�.0�]i��c��_;�pn��J���P����r�g`E�P�
&��!����ɪw<e�Վt'Z:7ٛAAu6a'�%�L��9U�
��b���j��0nI>��%�$*�f��Y�"f��&p|���q�&nP�h�t��Sqx���fo�B�,�>)���	���)xr?9!�+��o����7�����et��L�w7#Y��䨴��3r׉�<��Y[�� M=$��(�h��?ʗ�A���*7dy;��M�(���ѯh��T�:H���{n�sWj�董Z	AtC��dc<HF:�4�0�����S�3�*�39G4Ll�ĺ/GG,e�R�����)�w�6�k(ݝ<'�_���˰@D�x�TN|���s��+��(`O(�kO�-�����M�aY/"��H,�a'`u����[j��c�ճ�G���߁Ht��n�m��=u\@�	�.��Ř�l��^)Q�����Ua��#��9@�����i^D���F]�f%������mfޛ���^Də����@�D�~ ���U�`�Ӳ����I..�D"b�	Y����L'�;�^�n��,rE\�Ӌ��[d�-�[˞H;�Ï 8� + ��D��}�d�EU���j�E��1����,D�YJ���
�i�emb��QEƪ��հ�[��UĪ"�E�W-J�QFE�AUQJ5je0֪c*��P�+U�b�R�l����XUGZZ�h��A������Y�Q�Qb�ĭX��J������h�����Q`��� ���""	Z( �KFZTR5�b��*+[����jUMZ�c\d(���%j*"��UDKI`�b�PQ"(#KA�i�*����#D�Q�J�
 ���ڌb��Ų��r��J�R�Vffb٘�C#1�5��Q�DUVҪZV"�Q�YX�����E(,\���-Lq`�J���X�F�B��J��TD-@h�"�?oڰ�ޤr^����W�}��6O1�Ω��w��N���]t�Ig.��Tv��r�rRֵ��֫����l*�K��G���|��Փ1Ϟ�~�����T=H.��?��?�R,�P�J���bs��b�^�!���x��Y���ފ�PR;�u4��q �~p�4�':I���`Wu=�6�Z���u��w�=�7������R�1�|e&{g�8�$�{OI�N&�!�?!����~Cl�R(n^d:�O�T��;�6�R��O���ޟP1&���1W�
���>�z>��3:v)E��c���w����_�kΘ��P�L���d6��z���=�Wl=�1��I�oҚH,�J��?d:��H/Y����~C_�c�N� ��������=�"(A[���S�������n�t�>�I1%s,R(/��N����O����&������'��=k�'�SI8�z��1������h��MjAg��C]�m�4��Dc�|=#�7��'�B�*h}�Y������o�6�@Z�o��X��>�������1����+�+-��T�����C��*E�ɪu�����&y�����{v�2i'P��z*��DG�G�Ыr�ǘ�o~yﺷ��Rg�=d�Xz�4ΙܓN���x���Aj��PĬk�y�5l�3Hy5���Ԟ\�R��z�0<o4�c:Ԋz��x�L&m���滾]����/�u��oa��g�:}f�1'�_�0Ӗ�Y�n$P�8���L�%C�9�{tx�_���1ݓ�����}���ԛ�g�I�c�n�p�h����5LVb~]�?��ޜ'�����+�'������Vk�d�Ԙ�ԩ������u&0��y����i��H)x��f��N2m��Vxw�
�V�}a�w����x����w��{�_+�5�}�ߙ�L�νߛ�}�[��"�}�jM�� ����5���i'��z�m'�S�� �@Z��18�`V���t��1�ϻ�M�u+���~։� �w�rz��R,4_��w�g��bJ�<a����%Cԗa߶�m
�'�Mj�`T�`~��}�3��+�ɥ`.0+�{�����Ak��4��`f�k@G�|}�!P��>�/n����:3���D��VR���d|<N�//|�j"��u��݇��a�8�)��^ᡒ�E1�F�<�p20���Mo���$5�u�М}�C�Q��;�����Y6���|8B�귀P����/p���<ݥˊ�?�_W��ܞ_sp��j�G�B��H��"1���&��b�5'��֠zԞ�S���&�6����~|@ĜOI�4�L+��g�bE:��ɟ�J�2T8�Oɮ����s�ys��~��g���w�x͡�Y=ew߽����T6�6ϜH,���VV&09���LLa��bs��4��������5��ӓL��& q+%e~gc><�Hi"���M_�wO�����������[���r �Y�>����J�*�z�8�㏉�sܓi>B�a����x�PX}����R>d��c�i�O���>�5<H/��t=U������������rN:g��a���M q+�*~eI�*A��k�>a���"�X|��RW��<5̅@�T?!�S[�`bN�_��a�%����s���.1��H��Dy�7��Co^���Nh������{3���x�Z�7�M?2��V5 ��!�>��ĩ���Y�>O��~�CMa���{���=B���2i�Y����X�P������|�&�Vr�߫I�:�a_m���P�\{���ed�o>��o�B�a�1��欝O]>�*>eM��~v�Y��Ն�'S�c&�9�nx����1�c�{DH�,�����o|�JF��`cX;�3��L@�Θi���gg���(i"��6y�ڒ��Rjg�8�2Vi��������d$��'ɏ�
����������~|H9ّ�\Ov�3��g?b���O�>=�>d�Y1��N�s ���J���}g��O�;C-"���� V���N�_h�6��^��,�B�(�C�<t���`q�:����& q*'��������vs~��q��4�g̚��~3�4�b�����]�vO���I�n�P3�f�u4��Z�\�6�T8��l�ă��!��~����γěCDX��ꟹ����٣�Z�ќW܇����l�g���*OSs�a���L@�Va_ c=�2u��+�ayCR(m���|`VVJ��2z�S�R�<�0�k��Y3>ɧl(]U���>��}C��F��)����;-�;�q����Q�b�ǂ!�~k���z�}��J��1�Z��w�����~]�S�/�ʡr���܋Rǯ�^\��9L9DR���f���y��5.���d�u<���vԏ�
�v֍��]feWY��X4�\;��< V����\[��G��#���y�����?0�a���X���L���`q���4�3��9gSL����$�
�Ay�ݺ=d�"ϙ�z鞲Vi�kn�y�z�]���wռ����Dh��DX���uc�肓�W��ړ�x�`TRW�J��Og�c:�{d�N�o��"�4����7>���S�TG`u���C<����|��]z=����	�p/>��s�u��=B ��ݳB@cxʆ��4�ơ�J��h���R��f�h?'��
����4g�O2�@�q"�'���=�c8�R��P��Ăԛ�b�����B�/���<Y�˟�i��md���z �"!%N��$����w)�*Ҡw��F��Ę����HW�������,5&�y�����9�i�Xo/�
��Èi�a_�͟�1"�D	�	Qj�g.�3\Wgݡ��4z ���?!�g�B�|����4γ�;���1�PY�;��i4��s������1<;�O���0�9��x�]�y��m�
��|�CL4��X�j����x2��la= ���Q�.OY++���4�HT�`}L}N2b
E�Ì�q��OӞa6��T����51��R~g��f�̘�������4�k%x��s��1��.Y1�i �`g�k�w�__}�5�|O��:yI��S�V!�2q��3���mIP8���`i��hVn}d��0��T���0>jq��k�oS����W�3�=M<`T7�p�f2f#��:=y���oO�v�5��" ��&�guR<d��5�'��� ��i�0�8�d���xʇ�/��ځ�%g���iiXo�x���?'����Ă���c�Sn�,��o����}p_m,˼�$���������;/�8��W��6w3i8�aXW��۸

E{a�]�b7f���;`y�������=�ì������$��8��ɦT�S����W��\��Cg7��f�e���Y?&3~So�6�^0��?'�.�TGn0�+8�&;.d��++�o���J�I����O1��>N&}HT۶L@�*z�M�~v�dA�{��>B����u��gj꒏b�u�R� ��y����=�9׽U�i�;3�&���u� _!"�w���;o���q���K�����|,�_!ΦH�LQ3��\��CCsX��'^Zy�mG�FO@M��`�ĶT���U���0e�Ev���A7Z��j9��xwX1�����=�����O,�� �l�&�\���y$k!������L,�3�W�}_UWݺ�y��2~���Ǣ?zLz B"��SF��i���a�����z�]2y���u�1 ��Pq
ϧ��.�5�e���R�y�1��#�"����葃ۢ2�J>+���\�<��Xjz�~����& ~|���^^01-��+?2f_���i �C���u� �L��a��t� �����u4�a�a\`W��7���G�}W�"�j�}�B̬�b���=�IY�,����1S�JH/�=M�8�Xk��=CI��LB�ϴLa�ۤI�*VN������a��Ă�O5̆Шq3�>��v�2��=��/2R�_�=�9�QZ�7�t>B~g�?g�'�b���bMMy����O�4�~���O�C2c!���@R|��� x�P�4�P?{��y�|v���]&2c'���I+?8Τ��{�T%O�Y?:}`V7z�;@���O�i ��P��HV|�{g�P�Si�>��Rc�b��
�jN�_z��뿹ᯣ^�j�ʫɚ��"��@�}��"����"���_��K�(�weq��7_��3�U����
�,�s���jI�����v��WT<�^�Oj���hi_yfJ��yO79xj���6�Y����`�Y���B%g���T^C���r�ֆ2�DR�=��q�5�}Qg��-W���b�-̇κ��v�{.��6"�E30��V5X&�d����碣 y�K����~=yѻB��^T��sO�(
�-�@W)BB��Ԫ�[��D�\����-nچ@��t�f�whl�`>�!l��*�ͰV�h�R�c�o^9º����h�x�\�CJ�Bz�$��3ߣ��{�
qc\���!.()���^-�}�5�D���C��괱αx0���䮍w��PZ$+����h��h����ϖ�OU��p뢙��Z>uH�O	�(v�;/��X��V�}-�z\:�WG���}2"E�q��3=P��QF�ܲ`����z�$�i���
�:��62�sD��Z(k���tǺ�X�<r�1~���Y.q����$��
2�̌�k���]
�C���٘�b�����{]��d!��kґ�l���tr3�_k�g�ݜ#`(���o.a����i��΃��P��NJ��
`>���չ}���8�� ?�h��~Gת�KZ�+���W�I�I�<X� �m�G"�-6�*VI�R<��DD��|���2�s�2�ayG���D�������ڃ�>�۝𗯔�07K���A� '�,�:l1 
�л��������֟�Ç'�`"EB��䣺{V��!�bc�=x)�����Q�h���3U��V
��s�Gg���e��0b�Q�7�!p�����;(n\��(��W�<F�9~\����(9e��ј���v^bj�bHuC�F=R���'9�I���{�r�#C����6E&�@��PXF5�2�[uo��u^0���*�m��o�ak��G��_C������[�j߂Ŝ����\̦"F���r]�7T6����ZM!L�0Fa�9�\�<ٍ��8'c�5��w�6�S�m�W�/��ӑZj��0�r����9W����Ӭ�y�����uDƨ1�y)z�����٪��mjVi-��[nEϞ�SQgz���ե����Q�u�ٱ;e�]�=�"t��l����-������E~Y��:�_tڔV��6el�4��{F���Ӷ���]r��c__ϔ�N�6t�Z���]��W��{+"�T	LG�x���gj��|l*��dp��ޫ�pN��+%�a1{��y�B9���Ui���f!ε��m�$��.Z��܍�}U��G޻V�U�-�g�z��5�'�~ĺ���ݨ���d��%Lia�;�zL�zr���)@;��b59k������ڄ�Cfzk݇9؂\eL�s��]�H���[,V�����0[����g���;�@2���_��4�nhq��,��V�3�cm\��3Y�[|����Owi���H7�:���	9[X*��LUƃg�p�YZ�'oA肞��;�L�ӄjNL��=�{���=yͽ�̳7򚘗<k�y��m`F�Cr:��y�{�!o �G9�d�ݽ�U�n��p/4swM٩R�Q�]Q�S�^��v���̨r@����VZ�W�5��U����'�����q0ezo�d�^�yKU�u�����%x�W8��{��^ՙ�C������Xf�
��9�$&v&�_n��A,�X�%�Y��.��9�U*�!�'�7-�R�k���B��N淤��&����v�Ofr�X��=auy�I�yߗ��֣�kM{�1pL�h��o_��x7�W�>U�����gj��$���c�LX�y�; 1�>_�,�м߼��y[F��"���R�z#b���uƢ_k���v�z;�>{[1��,���� T��򎊬����.'m=�u�%[�]n;��¶5���k���_m��� ����Y[�T�[�y���~wf  �jm,��XClK8���i�]����L���K�&?�V5� �θ��v��A"��`%n�*U6 ��:�[���C��=�\��WV;���2�X=�a�Zm���c߻�Ț�0�ܻ�n���w�x{�������/'����{�|�e.���SgO�u�튵�`���ϗiU{ �O�.6��Y<Ņ:X�����n|݁$�oW��虞�V�{�V�oc��^���]�%bƶ��n�<���N�)�Is͚�w.q�bR*�l�3�#v2S��ǧ����d$�ČVhr�흊���99�'76�n�lդf�m��m4�\�Fڔjߚ�a�Us�>��=�\,���گ5w[�D_a����{�ߴ/v�}�p��4ݚ�R��3����#�x� ����u�";'�&����~�PJ�c;�˫�sq�ۜ�CXu�"6]�]~��5=y5�{6	W��8O�Uűn��]ך�Nt�!��kҡ�9귞ܹ�}�Q���>��s��h�:��T��8�'*9�;Wf|��w]��qu�&z����dٳ:�~�Gv��|����C�H4Y��{�W:xk��)ۥ0�
�ՌcvMv�X�;iv�s.>^�/�mV�FN�_����ǟ�fЕ�j8s$��N���%�;��}�2��	B'-P��Y6���_Q�a���i`t��W��U{'}��}�۟@����6rv˧�@�K��ߍ^*O��,����s�����$��t*&5[ZT�{{-ج����:��x��1�;���N�W���I�{b��:;uk9S�7�vr���j�1��
wF]5.g��i{*���(wq�Ꝉ{)OVN�7���1�k�ct����xr����u�,���9��GUF����꣟#�f���yy.J���ve�65��KzC��6��MeA=q^���\�Ubx;��F�V�qks�������סMr�6Ch2���b��\�:�E���nR�	�w�6�Rowc:�(��w��R���	��f
lm�bk{�/)�a�~��WOj&�u=ن�����{��U����c-w�".3Uf���VR��L���"sn��Ÿ��ܷ3bk���is97M�cp��9i���{8�d����ϒ���%:���Y�G!�ɻ�b�1���G1�aw�= �q��H��`01K�^�Ro�+mW&ɹ�u�>�f���*ջ�c\��n˻Wi��v	�}��5hIPx�ل�g��G���grֹ�yػ��%/�,�+(a�nn쬅s���뛄ٚܩ����<]����^]�U�.%�0:h��|��i-�����hr�j8mX�$�X̗�&*�v�M��tf�q1����ҋ[�q/6j1c�u|/a���z��9�B���%�@���|@���6��o�Zd�T6�Zc!)t�R��R��`��?T���в\��l4#~�'S��!�Q������<D)v���F���.��&���G/����c�T��εR)���8*�oS��\ TB~GvjejȬ��b����f�t�/���	��s6-���B�ܣ%�^XƬno���#�k�BqX�j5n�>�Q�g���s��&ʭ�ٓ%��fߛ���y=�Wʼ�eD3*Nt�����ЃWB��II6E�'�e��[��CeN�7�� B�J�k*<Mr>�uc�\U�=Z��)a�%��w�n˽g1zK�J��z:��p:[e�"SҰ�xE���X݊Pcl�;�ܨ��������|k]Ge�&�=yG�eu'������Ϙm���=d��B�򼸴������K6���7�Æ(Fl$�����������a�y�VUc����-�z�[Ƙ#s֙�
ǹ@�|��<�3W)s���WX!��$�Fi�Q�rei��߮�G��N�sٜ�N��KV��v��]�G+9>upBqv�;gLy۹�ܩ�蘨�++{{.ޞ�6�8樓|�8����<� �g�m<�����K�t��Y�(c��v�;�p���Q���\�Z���J{4�>W���]D��CF�d)�-}j5ό�E):�I�ҴTy|E}���A�+%��A�K�ɤ����9{��K)<YKY黀,.�����kOp\����Dh�[J�كL9op�;�S��X�rJZ�t=s�	�f��j]
�Yʃ��W�-��5`X�N�f��/Lb��H�g��~#K�i�٭�K�)� �M���8�;<�l^ΛW@(o��v��C^�n�KR�l��TRr[��`�V���+K]Rhv����-|&���7md�w�u��M�ʧ����әf�F����b%-�x�7Z���\�7Q�L����aXHܖB�2� ���P9ײ_1f՜����sx���^+�8���A�v��=��+4<�w}p�ǵ}0L���5�8�H]�Y]���\��x;"(h�I�̣K�E�E(OM�ͤ��B���R
u�=�ާ={'{ U���6��8S!��.;���=wOQ�������S��
�5���3=
��¹�>Ӛ\&���B����9I�!]ȯ�
a�����la�qf'[�hr���H�����m���CcJ������)Y�L�4�=%dV)�%�J�JM�H���� ������	��$݋�fK9Vm��e�9� 
��"f�>W�U�Θat�[-l{�e�^Wh�A6PNu��iU^�x���;C�ǈ+vB�,�y�n�T9:"����u������PZ]���"��v��X|�p��>y!����mAy�,��]���:�͈Sz���H���)hN5�Ӄl�l��ܐ��v�枣�
��,�+���A
���{���W�Ѳ:�S�"]m�_JiJ�F��hֺ�<�e������,��?���AR���UTЬ�����aU(ڵ��*�b[DG(X�[E1*�Y���E��H����Qb����,V0Z� ��q0�*�UQ`��-��*���Zښq���TUb�*QFVQQQX�KK�h���YZ���`��`��RTm"�c��������Ʋ��"���E��11��)�"����P��F���kZZ��E�X���2�U�RҊ�+T�Rڱ��a`� �����
���Af5�,X��GZ̋�ZX�QE�TU#�nZ�XTJ�cej([*�QfZ�i���Vi�+�����L��
�-*�0TP��m�QTA�*�6���� �@TEU�0�A`�*�r��QE�UZ"��q��1�&��
ͺ۳��k��^}����4�����e%�ɈJ]��&tN�s�vu��&���2ei嵚"j�J��1�9�?�[z���������K?g���;5kwbv�B��c.!����̿u�5�㍅W���w(��뉞t4#����L��S�4��T9�d
��车ݓ�F=��ɋy��wo���z$c����&�]q����b�j�b��qNrBݻ���J��ſ%X� �:@Ŧ�-w���uz��,��rquuT��D[��&GfE�V��߅)k�W�[[K�##�����67���K"��,��z�ȗT����yM�(�zo�<^]��'�k��dz��3�D����Od�Dp��q>m�2��ci��3�\�nSo���S;��6����+����C�Eݿ&��}��������U
�W�J�R�^Sũ鞪ۜÅ�tO�j?^$�3���]������}������46���*x�}�IߗH�n���l�b`�(;-�P�X��I��΄���1����`��E�1�K�-].�׊�dq��E����.F>1N²�G/y �p�B�X͔�c�=w�޶[�-�&��k�>�[ۉcj��.�*Ex���33�K�y��E��W��*���G��µ�������.��G���mC���3wY�l�W^|�C����9���p�{
,Ѩ4V���ޡ�"�F^�^yϽ5d�V}�mx^�y}�D.���N��21m!���N�ތ�l�x���{b����-�9��eK��ˣNվ9Z�+=���[���rUk�\����Uvj�� ���
��X�5�ק�=�9z���T�����&R�ݎ$j�]����y�s��Z��p�t�Q�+*	��|�$�6��d�؝�T恬E�y'��-InV6���?|]}nuC%���db�G�������rr3n6���5������bi,���&�����0�7؂z]p��
��#j�G1�;���{��ݨ	&�ڳ.��jQ�[�Uc�E��'%v=δ�xT~�x�:̃����\�uk s��	�O��5�!
�5zX�L�W�Z����2�JK'j�T�nV[�{Տ^���yN���3��N���y�p춻ӱ��[p${�)�^L�	K]�gqv��%rGld�v`W&@���X�Ve�s]7�� ��,'W��~r��ON����]��&;��:Z���J�!;d1�0c��+�V����u��$���4T�RF���q<���q��������
�600��1|.k���}��U)�y���ziV���Ź7�VB�a�d�rl��C�Qp��}ª%�%�Udn~;���+��5�w�Q�F¹��
���s��wP���-�΁o/x�jZ]y;�����N���+3@�7,d�(�.U¤��Z�ț�ǩ��n�u��۬�M�غ�3�W���~��[�׀��$V�u�Y���a�6w�T��Cr����<u칕�ߍ^$�AՑy�K��jð�hD�w@�+�V����ңu��*_=���V,o��e�J��3�-��7jn&�:��{c�p{TO�[+��j=8a�s��f��X�S�O�Bm�NeC+�abϘ��_�A#�����^�!�-�����9Y��	��=��`��<���Y��h#���~�ƙ��^%V�e9�|��ڪ���ͺ��V����Nf��kk=;H��b�c�F�A�imE�u��@��u�[��cA�N�R�{SF�0k��m��[&:�֪��C^���mnJS3@�f_��x5�}�U�oc:���ڨ��m���S\��l*mPP�#��(R�G[�;���x�K��]���¤mJ�R�R���Lȇer�eC89���n�[�2�n�P�ˊ����G�J���>�\S,�S�x���x����'����34����o��-�S�1�+5˳)=��^8�x'���eHG�ƙ�&Ǩ,���~�Us�+0u[���2f�uryj��'�S���IN�n��8k.�G%��T���N�:&
���O'��[-�tyY�}�gmtP.;eT����%�Q-[1Pz�|�y買;*�����d*P��S�|F�q
|��w�˨-i%�|K�m�����+-𾊵�7��x�z������Kup�kB�a=$�~b=4P���ܭˀ$7��-��]Y���ףTt�Q��vʖ��_�`�u1��)�C5&��B�G�U�nK��-��ۗެ���?D��vF�f�^YW����U,Yk|�{qV7�=+�-�=Cj�v�Dv�l|�����-wb��+G:s:YX���gS{���zL���l��*�>��O/�B'@���������>a��5��Һ��t�:�ՑY9������O���Ꙅ���8��;�$���^P��x7o�E��rnq]T�����]i�����Q�%l8QC�H�'U�4��E¥�~o3n5����/".�<�R�|�o����N/��a�y./��1
wU���bTi_��Ͼ�$��-Ü�)���-}���pE�v�����㽸���h2a�[�j}���݄[}�%޻��[v`�ة\�,�덣����Y��m�_��<PklG*�-��i�y�s��0�lt�L�'�Iu�"��=پ�|-kT;H�	�x��n^]Ƹ̮w�5�^J�r��t�A��OG�q�����n�r���o����˵y�d��96Ϛ�U�;�X�2��#�+��bt���|k1z��bH�Ukc�ͨ�,�Y��к��u:*\9R���T�Z��e
Ū�H�IT�i^��6�h���V'���=��.���%��T�Z�fV8]�ZHO$���ӻ��Ν���D�B�I��	�U�I�՛K��%�t��hսJd
��%r٢���q髎��4:�r��t�:� ��@^�Pk��;�{��J{n������+"箾�vNG\�c�z9BaT/Cn���4.�hnq4\bMR�;����ǎkڲzB��&ans�y�G��إ�ѵ�K�����\�'^'i�@�̿K�'���vҨ���A���6j,�ğ��r�B�^M�4]W��L�Ԋ�pw1M�����-���)ek�>��K.�tǹ=ԛWԢ*K�.��,9��+'+ة{g�����ȺU�sM�P�>�Sil�o�'���7�v܋ZB���InUP��%�:���k�ʙV�[��=-�d��;˥W�&d����/�dB�x�k'8ڎ������n��Vs�kGM=S����N������p�arW�^�gq�Ga�̍��@K��u�]�^\^5W;4{���e.�ڎ$a�<��1�VF�j���p\B��z���2;�^�R���N�{��ŕt5b��K�v�j}�^a��]�ѧ����s;AR_�uƷ���պm���k��1rQU�D�X&J�NQÚ��sb���z�gpT�!2��t^\����F�vɗu(zUs�a@��HD��A%�����ڔL�ݬ��ߡY�:����#̨U���Q~���%t~p�D��rO4"gft��7�^��~�0�7|m���%X�yߺ �E�����f��˧ #>���j{�%��o��
�0�qT��f�כ�1���%���ʤk��Be1�#!�����Y�n�6�z:��D�7f�J>M؃Ph�c])�v5�O<Es�/n�B�~�ym|��6�d�M��W:9D-
y���[��ɩ����K���'y;����b�Q��o�*w9�·��d�I�.�"^�pب��2:l*���ߠ�͛V2}����N��	��x��{��J��k��ɈMAT��B��M��A>7�!��W�
�^]�a�T�
��J�[���r���}d��91���[%ƽ8Թ�P�jŵX�0z�>�t�
t���7��`�p�dD٘{hcW�jW�Kfg%�{q`��K�A+���sV�����C�`S\4e��%+�,�.��+�zb���	M�]Q�y���{���a����]SCI��W�\�I+�ݬV�ܸ��8��ΠH��7�Z�|���_WԴ�)�3�x,�Bxl��S���\�Q>�lח,|�q�_f&#�;����HC�p-f�<̩���tu�(�^8�\�v_�n_#����S��9ȉ2y"����y�+�9��B��B�i^����r;l��֩��c1�h5��ܖ��;N�w����@v����7���D�U�z��r�ik�¶-���j�rZy�f6�c���q����T*�����չ��5ss��_Y'A�\�ؕ�<��#f�J[��2[��:g�����3�9��V��J����Sꈺ�9��V�3�9���H�]]��p--`�vE�w�Ta���/h4�����ҽ�q$ᬆV�֭�O6�.�]�R�Qz������
�t�m����00�N�Uq���\��7EU�y��I�\9��1pz�f��d�*�y<Z9����TP��­�ﺾMe����+b�=B��1`��u�:���h��͆�j���x^�8;���#� n�&�;�ثbG��{�;#�Zխ\ɽ�n6�I[�{��ڏN���I��r6�h0b�`�6"PԾ���_.�������P��q-�S1�=�=^D��i��+:���G#�W:�Y據����HS�!��	�St�Gb�Wf|�>�F��1!���۠�e,���D�=�x�y�O����ߛ�hT�{��R�G������3=5E�2��m{����p2�b�yi��Pc���n�l�a�E����Q��O?e�h�\�����o1F:��F6�%B��1�m^sb鵘2U�7Ȍ�6����j�,���U�8��S��
1vh�&�3��|��.�������3P��\7����,���I١�+N�=ʜ�!��a���]5�i�4��u\�9��C��oF�,@*�V�-�����I�W]�j:���8�&:'�;��Ώv��M���7�]f�m��ڲU^� S��Jz2����N�;�z>26�%>]���=�ϖ[�foRF���EM��	��3�����(�33LW��`�}=�"m@髖"��
���;q�q��-���_m݃��=�����[yx�u>^��؞�׶���U��1^�ڍr��ܒd�V��uڅڵk�������ř��n\��^�w�DC��lUқ+x�Y�zu�~���
�Ņ��ܜ�f�}к.��V3�4�H�Y�`�=��r���,�&z20�f�s����>.S��K�kz�W�;�l=�G���;���K��)�%�TT50��~jR���>�]���x��8l^�uTLt��b��Q*Y��=��v�L��a�2��q�#C=]5�}�~�sßvOTp݅q0۸�*��+��H��6�3��ZIQ>�v*�Z�i������}�O^esS՞W����t�iؒ�*8C��d����bs2�c�ŀ�buR�8����kyꚙu�tT���`��ŏ�߄o��d���Ψ�mj��|�Ŏ�z�R�4�o'�x����D}P�OeJM�꒟w^r����jȬ�:C��
�u["�[�y��0�R���|��j<��cq�\��>�O��x'��hK:�����0�s�z.ƞVJ�'��/�b�'{�nfj���{�c��3��u>�h���p�Օ<ɎGL*�[��]�9�>�o�[�n�t1j�`6�����10�_}
�!k���ff��]A>�k^��Wo��mp2*7z&�u��%�خ�{���z�z�t]h��	h7dj�z6�Mnn=������_�{|{�2�V��E�K1S���)��W�y��WvG�7sa$���.�V���ӴU�ns׈�C��1�;�uNgqb�{�0�+�mLO�e�j�k@���ʜo�YB2�,��(f<j��I.��!}��3zՊ勏#�'g��WɎFzW��y,�}]2�~�T�v����j���Y&�m�V��V����7����X�VuT � �`a�/3�(�g�1J@��\1.���VIt�=��������x@�[�2Ƨdh��{���0F;����r_X�{D��ie ��ܮ�zU�*nXUiu�c���kWd!����_S�U��}�r�D����_:p��:�ރ�V�����Ҋ�j��/�1#nZ�[�6!�����m�=wA�_S	"�9�q\�O�^d"r2�vs�C���,�@�����X�i�]��`
��x3��l���YJ�}pr���ʺ���}�z#}!��Tc�ԅ��k0���
���gF�1�j��2:A^b�;�ߺjI�@u4�3'�h`�@%�5S�IQ�=��3sU�b���nn���a���*7����+�_�,�f��-]�DާR�}�.�)I����-��|k^<�C�&�+,P��'�e��n��If�8�Juv�s3�S�H��r�m�/Do9����3"O8,����cBw.<��qPB��9��-VPvX53�=��I��8�x+��t�\J[eѺ�6��j ���a�1s����%y.�����byX����l��R��~�[������Apy)N<p�����d�o��];u��;�iڅ���q:�n���S]f���X؏Ekw��.��T�T̰�UD�f��ay6��h����m4`�b SuCe�;N�\R�_n�q�&�_��cP�/3�VVl*obu����qR��aM��S/NDA��E��9.X;�2�{�o����FF&]1��]W�p9l�ع���*H'�J�ɢ["�F�ӾpAkjt��]g܌U��a���̋���jb��˼���u.�݈u.�wd�Kj�v�р���l���ԑ��(�Gyo/f8�g^��RS3:�S+ �,\��<���_�Vd�4��^�`��6�w��]�Km�9�W�|�!�0:�+'��H4[GEL�)L�\,L����$b�M)�Wm&���bT����x/�{Xq�p3��}�.�͐&<q �i��Q��g��vֳFʳK��7jQ#i���O1;��ل��C��Xnn����ݼ�g��o>_!�7o6�'ub�s�&B�4���%-\U���.�%B��K�ڂ̖���k�T�2��E�T�U�0�\
]��O
��QJ
�0�\�2�8�ffG�ŋv����T�f�ۦ\8�Sp���S����R����("E1�Jԭ"_�bE"�*�&f,Y�֪"
��b��j(�X�.Qkm��ʖ�PZ��
&"ō�6EAk%H�*U2�4��,EkEQjV�(���cb���#Y(�騑Q�*"�TUPb����*�Qb��E�*#-(���*�D`��Q�*�У���$QEV(��"" �F"�*(��QUEY*�*���U�Ơ�"1UE��D@Fcb�UDDQV*��)ATQ#X�EU��*�*(�c+�*�� �T*TU*��A���X����
��*�"�1QQ�U��P��DEb�cU�E`�*�����"����Pb��X*����Qb�� �V*�E��
�TQfe0b��A0PDU�$X�EH��0b*(,VEV"��UEDPUb�������Tb��1F,�Er�)#U��2رU�E�m)1�S��"�(����2�ݱ�:��@���v{;
 :i��e^��;mq�Ud�B�V�d��zֵ���&�W��9b)&�f�#�hꌛ�r��`�S{nפ�ͽ'��Vf"dx�*0gס���� E/t"����Mhp�Qw�'A ;���_U�[�q{��~�ı���@��G�n5V���9[<�.�k3o�=�9|O+k��WiV�>�3�ɱ�6�M�[���+�߷b}|)�s������1��U�!�=z���v��Wq&���~���b�Qć���`z�K��'�I�5#�+�^�w|z�}1͠!��ʮRwKq�
�V#=��ڌ{ۤ�����z�������*P���`.4$�;s��ϫ��+�ޕ�Z�ݵ�F8Ɇ黎6�E�%��>�F� v��7��&#�ΐ��_9�w�k�E��+q}K�K�Niy��#��OS���܊B"�5Vo�ueZ�o��v�N�f�^Ʀx:�Ș���/�u�n�#�l#M���V��^yxB��Нa�U{@N+Ʉ�=��}�)잡ɲ�Aؾ��Qߥ/���:��{|{���Z���r�����u!����o/R�>[���c�Bf��Uw-�\'ʜe�|��RIE�/�`4]-���܄��4��U屨�0�_��-�9�n��鹿���C�|&�I�z����y�j�*��"�U�.��o��@s���>���S�MNSVD��L�o�Tn���$+)�B���WY���[Ǜ6=T��-�q
Wo[��0��P��sP�u[����;�~�=�/�H���)ݦ�k�v�J����j!��<�㬭����j��@����1:��q�:�u�7z'���������ب�X�(X�nݻ�+�����~��v#�&���yC���[sy����۟I��Ԋ?+��}�:�\��-��Yqu>u�ӭS.:�ޤ�A�8�
�DR]�<M�H��މ��Юyﾗ�����{�+˼���.D�MI�q��_t�}���˷u$��=�q��@o��wWT�t� ��|�����{<4-�:�锵Fۥ+��Œ�7q�䉔Ԛͪ��'��n �);�w����Cb7�f�fo�S{,f����k����V��<�u,99�.�e�
���8/J:y�]���Tü���}*bq��
ѵ�>��訷+);�Z��"ugK�:��=Ri�0�UV5��L�[�P�z��3ҝ,�G�����u��9������כ7�39[�x9�T;��^��0�*s�02����qX���0m�yl^��Z����6�����;F!|��ER��},��1����&+Z�S�2l�̇���^~�x�����zUDبi=��51*Y�=	T3�΄;N[�ܚE�] �3���%�δ1�ER����;��	�_��b�C�&z�|�ǔ��N�W����S�[�dk��u��S��k���w��6���+o��{^���ƀ�f�G9M^60�;T���]�sܩEUi|��u$�=��{�J��:���;��no<�5:�����r=^��3�r��f���y�\7wM�r�3�^s��"�r�F:����캋<�<}i(�Ĵ\=���N���>w�b�����ޛ�+[؜5�M�.�C&�6��U[����
�ܼS�$�5��Y��X�7'���;��7��:gF�#� ��Y�vÖF��\�P��II��YE��v���%�Z�:)լ�{�.��n�w���H�X�|: �̺	���Vћ��y�Fr�#�+�k���!�D<�LLG7�p�f޼=^Y�W9���$�bp����*ܔ\4;��Y��:pb���'7��Oo��aZ� �bc`9��X��<�mK����.����V��S1�$j��f�{<���{����CԧLu���'z����E�
��������#ߌ�vztx݋��Z�o�g?r]�������Ů�]����S��1��ާ���k:��'��1N-���5k�VL�da
�Dr�Q�.��g[j,vRY�$��Q�)[<�'�(�NE�(��C<9O��:�v��\*�Q-��ϹZ��[�z�;F�Ϲ��>�V����x���H�n&�B2�_I�jF�Ց[������,��W:Ø잨��;��&w5�g���p����sUa��r�����_d�bǪ�:B�k>��Wy�yy���+���U^$�;]�v�����<���r+�N�{*3Io�u��i��<5����{e�7+��/��]N�h�3�'��g��������:��c2RљX��e�*��������1g7��zX;��kET0)p��{s�%K�5�\ɳ���v�nj��~�TO'����P�$8��c>K���3�� ���[2Ӭ��*�ll�}N��?u�~O���p6�e�Ɉ��O�"R�����ˋ���h���}2v�yv{���4K��>	z�.eFM���*)=��"ު�v�S�{Y5	ຏ7�v�ȸ���V�9��z��Ժj˃���U:��x��:�q���>>䶗�n;ф2��oGn���{SK�̠q��f\�OK�I�}G��o�>���M��V2{���j�o8Ճ��!*��TC2���)<j^�G��|.� k�{=��_$��>��j<�.�� ��d�ب���{�)�)Ri���yv^�3��Tq���S�Q�6:���eB�����AL\v�ƫ�LO�G�t^���yF�����d�M����z�K��2&x�B�J���������թg�\4w<φf��+���B���Ħ-��-I�w&5�-0/����l��Yc*�̄�͓bIǉ���3w�qi�l�6�N�R�8�	/��s������8ó�aWu�T�)��'�����K����٨r���OiX�țB������]�9�^/v��j�d�[X�<�+բ�en����^�
�~��-B*=Q|��uQ��7磦Yۄ[�i�N�Ԗ�Uґ�Y���5Q�:b(������Cho�/v.�q=�onֆ�A{�ص�R.p��ۺr�����έm�I¾��:���P,:JǕ���n����(K�d�r���Cca�g
��Tv��c����b�;�HQ��s�[{�	��U�i����؝L)%BZD�B�6��GF�O�X�oto"����>�ce�����n��<Y$�>�qJ-���G��������p艹�����ݧ�b3z$��vʖ��i�U�ޤ�6ʗ)���YI�Tr�`�/rW����6k޳�Q�s1j-�F{w�}���T��0с�z�qϐ��kk�z���#�������E�PM�������j�ڲ��)Los`voS�Z�v]�Z�yE
uCs�M"�@�OгĊ(������Nw�����+��+����݋����y�z��E1�[��G�n�4��s*����rWC��˽D�ǋ;��:�I�
a%�h�3GN�_R[�:���@*�O��l{�+~\CߢW!�K|3��\\j�[\�s��������P�)���gozWf��r���23<���-we�cV��ű��W*��^ҜI����vD&��g��������n�n����u�����򠞸�`�ƻ�R�cl�)\�\����{pU�6��o y�s�n��½��|*"\�����Gͺ�S�ytBW�e�Y4����WCY�����r����\������}Nf�[��;����'�I6&��h����ݚ�J�i�j��9W�h	�V��XZ��넡7;�Y�"��t��mA��ئ�'�����$���[C�Ȃ�A<I���0){*_���	�\JuPb��>��.d�Ηun$�~Ү��Eu���{���&ս�Փ�ks��4��j,�p��n�7���M���f�]n�)�4���<�jI����X΋K�^��u0BS�d��9����a\d7�Y}��n�o�Φɯs�4T��*gu�=���4��Y�py�ܺ	��z��{w|�֣,���zy����K��jK�w<ޔ�	�pz�"^:�+bӝ�U��w���!�ّ��������;;�� &xEU�ۃ�kk'*q1J����UP������%�Y�c��'��!��wo@��N��oug�'+c!��d:y�e>��ͦz��]6o8OOJ���{��>�3�w��w�d*�J�I�{��Fv���91:�u����R�	��p�qp�*�̫�~��kj.:�o%���+��UT���.NW���I���z�Z�E���mxf������N���n�Ϥ�����c8Yp�L���cu�X��
��U=��CޟQ�{/q.�㴅k.��"i��3�ۯY��#�{
Ȥ�Q�TtW�EOv���Z&)<�;���l�˶�W>[�9�9��%pͣQo�`�{�(�׌ӥ���-Ԝ!gzkY�&������2c/�;}pJ5�K�2*ugpd�8��K�@��d��79�!j��]��ɽٽY��*�歔](EٔU���P�^J�*5�&��$�Z6��vp��@�q�o����累4򥋙��"fa���a[�	�U�F[�
��i*-JURUC�o3���>��4�/�.�������u�F�&�}E�Ma/q�b��ߠݺ-�z9>
��O�ИjQp�z rO��r�}ܞp���1�j�@[upԽ���rc�ob�T�J����[�qB��QLM��{��T5}�D��[H��o*3���{"4쫎���L��ڝ��ۃZ��]�y7g��0��Nz��ʙ}�X��j����X��P�z�u��4�U�9S��Q�������y�X�����W
xM"��7X�|:{��ݸ������?u�~O�	�whf\[űLSu���I���}��y� �G��*VK�p���7�I��h�^	y���=[�3Y���چz+'1_b������r�i�P��}5"��1��<I-���%�QF}���T��;�r��V�y'���f����浨n���Z9��5|�w�;#��J�D�u��\��\���M��&��|��%��p�픘�����ˬ��q��ފF�ڌ�<׉ҕ쭴�����^S�+zns�VA�`xk��vWu�����P�W��8� >�ه�6�BUZ�3*�Ob��Խ��{�ڨZ�����qG������t�3���U�P�*����뉉|��=]�3I9�3n��]Ǜ�˦�`��).����oj+�Gd5�e®��˓=��p�3=)�s{Gg��|�7����R����y��9��|zSL���$���V��|�)gk�7"UX������u�����\�{��JV�^h':	r�~��B7�ʉ��k��9��G���y����"�_d��)䓟�=(��\F�\��P�a��8$�[��)�ū�n`�Ϊ���_w)���UqW�8�XU3�zy��驫3ͺ�mo-7q�Ϧ���}�'�GL%3�9E<�oH�j٢��[[��SH��s�mu�bVK��>��4��C�\��57M�j�2�>1����k�:EU Wb�U��J���6�w���%�Ay�f�&�o�p�l1��!:y�F��k�vՃ�GV�
]c�H=�N�^�r���[0��c
�m��Χ���D�WT��Ó�L��0��h�E	G.��ԍv�^m���u�����go8Z��[v�t���Ԏ�Z��Z�T;Nd�bm��������m]�;Sܧ؍�h��*��bd�B�G��U2a�vk훻���y*á���ݶ����$��L[�I�DB{M�S9h�����Y��f7���l�G��dk��O��)첫@�\��;u3GR7*�����Ζ-����9YtS�e]5�F5v��vh�9dw o��*E�M��Q$���]h�E]����nv͎�t�u˽�B֖�Ǧ'�ӽDN�gK������y~�ņ�uk�m���7���g�ZHw5(�v��ڊv��ǔ6WBNc�u�2�N�N:���I��~�G���3IŸr��Up5[�Y�j���w����Ł�W������M����wX�#=o&���[�ٷ�`�76V� �j�tV1�]3͓�B���i���}�E�Ng\�΋xɡ�Fk��46�$�/:�=�GW�㒸U������]p����Ƌ���,m��gm���njE�y�U�*���j�\�Q{�C-B��;T��C�{��w13�J�b�v��Y�KX���X v��x�d%�����f$�b�j����Gb���h���盕*]���8��]Dݤ������'�xF_��5=���G&��@�WӳX�Hbp�q�Y��'Bss�&vj3 M�b����I ��^ԕ�ⶌ�[%�p��j��Hd�FW�v�-	��6�^�Nh<YW"�����zN�����nG�J<��
��L�nx����u2s���Eve�ۓ��u�	]�s@m�4�4И�����9��j�?�"1j&`B�J����S�#Y5�hf�F��u`< 2�.�՟����c�= 0b�r�1���7���V=�3"TĹ9������h�T5k�>7�&.��dM|iEv�H�{ G�=G�Jf@�y9F[�&K��LN`W��F+����z�`���w���(,��=�d�����+�cif��]8` X�4��4�U���7_�'H ^��&<W��R��R �Ӈ���8*@V��.&r�]I".�qs����9�h��ɜ��_�"t�VD���;�&J��L�omS�c�m�ۇw���"�Qb�,TV*���1b�("�EQ��*��QUF��DEAA�*"��"
V�,APQ.R�Ec�,DdA�Q�Q���(��j�UX�DD[j���EV
"V,EDPX0�DLJ�FEU�,����1Ŋ���,E
���DĢ���ȉ�AQTb�(��PdQ�,Q��ATb*�DV6� �Qb���EkX��EJ����UAX�H�E�,PcD��"*�j�"����*"����*(��Eb��(�DS)T"��((����"����b�`��*�QDE��e�Ŋ
DF*DŌPX�dTETPETEDV"�UUV1V,U���Qb���Tc(�UFV[jdU�TUE�DX�X�A�A�TX��TAV(,Qb�A2��(���UH�D��� �1(�Ĉ�2�V)V)Q*F* ��ڮ��������߮��N�d�l�PV���s�F�J�7d���K.�DH�̶��yW]bpr.������|�C�;��{���_g���VM%���_q9Y3N+���u�!J�r��Rr6�e�qZ�ɩ���89��nn�����u��Y��R�)}X�$]=xZ#fy5gkަ���s+�y����=kz��R��L�X�Z�Ԃ�U]K���[@BJO�z�O�i��{�>NT�<�db���N�,v�4vOr������j�p�x2��X��B��ݰWA���յ��ٻ�;bk��.���
��3���զ���x���'E�⽲���5.�)�<�=PO]DJ�W/��iN$��e,���69�\xcN֋͝����@��gՎ��Z�mg����C�JD�'\�\� 3s�A��nC�.qtfmfMv�T㍍��J�l�;΢鮺�<�YǍ����;-F���̵K�W��U�d��[yn?{�X��w�^AB4͊���+�X�[0V.��� g���!�Xr>+�ے�+}鷺d�/
7��Ua`+(p�;����Y�ɏ�qCs{�&v�+5G#�qې�u.C*�c�9h��KQv���-ꇻ��������fo&U�3�����I���\�*�}�a7���Ɋn�zT�MCUc�^��V��*&*7V����]�lw>հrz�ra��mٯ:}u1~���0��:.I�/��Q�cC9]5�ݵu;��m�s�%��j��;OI�4MCHE�yz�W�"e�+o�wj ��v�U�H��p��Sxf�R�[���x34��ۖ��I��ps3%c�V�s���<!W�+��4Y����纡m߅�6n�*k�zb�ww1M�ȜLT(�lp3��sR�_Oe�~���\=ҫޑ�@����b�K�O�<������tJt\N��kTQ1Id8�ک�+y�YבVa���"������u7bU��U�Q���.�A�LN��{�2��߫�����njcw�.�Z9���MFPt��\��*����ܹ9�jb{b�3F�u��R���)/P���]���_m����(Vx���mu������_T�*܀Vc�JA����E\�<���v�OL������Mݫ�ȧ����,��9��ݕ�_U��-e[���ˌ�m��nR�������A|�3�s9���_}:Os����H�Ьpi0g|Mo\Qޯa}�Β�'�	�������'I�̢Hn2k*��!��)P�:{+�M@�s��{B0�*�e��Q�{t����~mk2���8f�#ӱ09\T��GY�6�S�GK��G�+��u=/�Wt�HN�yT[����6��FUz'b�Lfl���x�t�qy�z��Ɋ�Je���@�dӠ��]�;��whQ�n��J���b�e����=V[W�v�r{�-�Lu��ź��p��w{rq��QYԌs���0q^]'�
�Xn�	�=�7�ׯ <�,�yrҴ��㸢阣ѨO$a�w�X��j�!E���P����]WY��V��O�{��z���K�3���OU9�˕�kذٯ$�T���t�j�禱����T�q�LCs�|���$��}���o
�]�X�8��F��U��YΡ�H؅>��F�td��ʁ���7Hb?��9-:��zhe���͢5q�*�&�s��n�����R�fCWFJ���{�!qA1��}�TA�q]]F�d�1rZ켳�kU�t̕����l sk�/ވ����4��R����'�ѥ�|�\�nvi����l����f��Gh��31�s�8��}wslOcy謜�ocT�Q:�׻��=�5��"�_�#��&jE�oK��>��r�1�pü�)^^�5Ք��mw��c�`$�r�zd�܎z��\�Hr�=�W���pVO�%��g`ku�{�Ζf���wí�{�̜���1:��,|To��GT�Q{�_-�L�Q}�o�E]7�&�l�.ս)��n��x�U�)WOFT@��QU�����,�y�g�A����o�m�3��簬�FbQ�`�t� �ܤ��x��L<����^�K�)���o*�cr�����ﱚP�椦��w-���R�/�~�3�ط�9�����q���k���!�Ŝ�V�St�o��F������Ș���5�i�d��f�X�����&���j�F��bk(��z��x2]eŢ�0t�U�g1�qB����1 �gX�T�eu��pA�P�톐��=I�q�#=��СƸ�\Q���PQ��+�/Us���ǉ`�O����7�+2�������5w��5��9��ɩ��E-騉�)�j�t��0o��	�*�ff#}ݛ�}��':��_��Cm��w�©��;A�ܣ�E(=��ۖZ��}�ۨV����4��� �F6%��;��غ�0�3G��f]�r{2WVz{:k-���bU��8t��B��$ϡ��x;}��\̓e�⠗��`�����VF3햸�Y.[g��:�
4��N����q��Rru�5}��Nb����Zzj7��e:�n���R����غzz,�oN/&^m{��׺���C��&������
͸��jS�����W�.>�yQ��U���&�I�[u�vnL|t?�~�7Ĭ��C���|v|�b}���y���Tc��0w_��S2��5{Zn�s�bغ�qE�er�����\�էP��-�
��� :��Գ�Zl<;���֣M�����5�Wm��+��w-�(V&>��W'pW9fk΄̱�)��WC}�����}�~lt;w�%ܙkz�G1d��.זȭk�P�3/�BZ�sv#3g#Z�g.a\�:�U�v�D��;rw8�ՃG����aT�e��3�a)����a��I�$񧽟.��,�Y�3˦�T^��6�ֈbغ��+����e�z{Ot/dK]rK�"�l<P��oR%��+g�����W�RuPA�	o}~w��/d�TzV��|�o ���N#�;�Ǳ�LRkS���%Nz&P�@���-�ۤ�]{�O,�x�8��r�z:|�t�)R!�r!��:�[��M�T��� \���]��wNS�]1�]x��rc[��ݚ�O�и�ݧ�M�G�fgZ���Օ��	*�k��v&��:��s�K�m�����:�gjlU�nga:�gz�wMz]�V�U��X7�N|xOOg
a�5�i!���������2r!��&�iτ�eĬs^ŀϱ>�C�5i�4T���.�6�O(�[���f�=�~���������h騭��0Sou���*e�Q�#�]>]�wK��@� Gj��j-{�v
:�P�p���n֛%ʒ��ѩ�r�j��l`�D��J\�ɲGg�o�3��1�Al���\wNc�������� i��T���-k]:�;�BູR�&�%���}ۨ��u���L#�^[*]����yu�.��e�1o��
�z;!��s�d��
��^�È�q:��l�x�̷�K�e�2(,�q�ܩ���vU\����,��U\����LϹ4��ׇ͈��C� 0�������� �㌜ʆe�FP�q�i�U�ۮs�'6��$X[�oN�6ѫ���V�k���цeu�I�WE*�/��S�U�����ʠ	δӊ�{��z���Ց��x�H�[��Kd�)���t���U���Q/8���{+��H��~u!o}#�	���Ft� ��` l�T���yDk�~T4{���������D���)�����Nr����S�q!��æוy��D9���2��Rpu�(\�]pL;1�G��Jǂ�zvۯpB���n�D�74���\nr�v�ݪ�ky{Y#�E�K6A#"|Oi�>���+bgCF��4����#E��T=�lwC��
0z���u��=Ӈ��oT�jJ�k2y��q_���T�nK8�$����G�eX�@nVsص���{ ,��_L�y	�Q��3��\��н�����	R ���]�|��s����`*5�s��w�K�T�ʕ�P�t�f'Gǿ�e�]MOAx�ˣG)���0�i��en,�1`B>�V���Nڲ�ڜ	{W���&ڷ���[�>�x���'��̽�z>M+R��v����Ā���"*'\H�S9q�0����b��x��g7�g�j�%u����)T2\�_��P�<���X㲼T�:� �b3�s
��o:ozWA�R�򇳯�PئpD��j�o<U`�$�z�$��^p=7֫ǡ��|�^�Do-��[O���f�9���B|A��T*:�~�.�=�N}�u�ߟ4���R�s��w36��u�*	�e��B�U�ѹȺs���!��A��s�J��[T��1#��a񹙉����{ٴ�L�m��k�.w�qE�N���|Շf_���\rc���Jݛw�}���zb����i�𜪦��40C�BM,#�y��~��< � ]q��ֽ�Ɔ�;�{�D�PO}#.�����_+���߲�U(*�1e��_qcL%�J����Ws{�����] ��(A�uQz�G�6���s:�I���|n�y�{�[B(X63�:�:T�{>�JY�R�<(0�LM+�L�U���{dC�$�u��g(��}��~#!����pE*�O=�7��ɇ�����bz�²�m�	��+��c*sx��Z�}:�+RS���j�uɢۢw)|�5��p��+���i�۩[��n�nX��녞�r�%��x`�T66tB�wΐ���V�N:��L��$���0���b��ǆlʀ�����Ct�7.�eu�@������n�)<a�o���iz�:լmN$O��¢5�ۂ��k�a~�,킈�Ƞ��j	+��%~����9�s,�o�1���\M5;ENG<�Nz�
���O.��0�EV��<k0B΂�!��.���!4C/���OI�Ֆ�`1�#�9�L��B�X�Jy�4l`��a�Dil�PX�t�AS.H虈]P\��3��c!yyy��x�i?s�y�q��<w 2��c�s���K���s�)� .(�$�ǆ�;2�6o�-����^|#���z �zhn)�륌��r"�S0��Nz�&.W�.P��ғ�V˩z���7H���C͐���Ї`��a�b*1N5���TP�S$D�ɇ%��8��oŬvM��n[v�{4;J��kM��G���V�a<R�x{��R��o���Cl��L���RD�{��ŷ��f��vt��� ��Ȕ�Hn�8;P5�v�kO	�����%䵪���@���х-4�r�`؂b��ʪ���:�.ƞ�̸�ɜ�!e���/�<r�h���k��[Ρ�ۦ�ub
�4��n;�8T�d���՗�E�o�wv���M�Q�����`�o`|	�d�'YZ!g�c+&�XWU�;�g��n0���F@p� KSh�ULp�}6"i�YM����nP"�N�ɝR*⭼�d�˧�g66EIfOS]+k,�����7/������|�$Fl[۝7gIB���d3*Csu=AWOYtH��-)A!M줥��yP�B5�1����|��`�n��J=4�%���|"�yL�eY=��ה������	h$d��w�Sdի��:=#D4��q�*�'Ҳ|�� >;�-.#�=Ղ����F �w'4i�Ɋ�Zp!�U��t�Y@Hx|���\�UꩌS2��DI�[,X�<��������eu���p\k�ŋ� `��J�e�4 AY��j: e*�9�(ϲ{{^�WF���
pB�P�:�ᣞ�U��6��4�H0|��m���Y]z�Jq�#����Q��E�B�� `ᇥzs����[yq7�sP@1��f�Egd���ĉ���a�Gi��hB����`f��]fZP�xM
��rPq�Y7(�|��̎�N:���i	�����'
7��6Nb"jw!Y{c Ν�z-���!��2�b��{�M3um�>u_|ʕ�����}�У�%3��1Ѩwr\R��0nξ��s5Z*�I��gtT�M{{�E�X#�.�N2y��;;"d��1���f5�^�����L�6#���j7]���I�Em���;��;�e£{���u
�Vr�a�LNZgh�����k��haDI���X��RECm�([罺L}�*�̭L��:�>�ޭѨE\/Qf.K+��A����/]z8/��4����BRKބm��o+���[t��[͡)i�`kG�&�L�.Xŀ�^<欢����>ϲ`��g�ξ�S+n�������w��'DDa�tb�:����nG��P���Fd�7{lJ�都���.\$W?I?\���-7����i��ǲN��,65���楻Ԅ����� ws\��ub�Z��v�xKI���*l��@�<Fb��_m�vD��0���Q�W��+�ڵM����4P�AC1����Pܭ���
�ۂ����'�0��*��%2Q��l����%��y���R&*n�W0F�L�5��_1r[bG�K{)��]u�8���DSp^-��u�JO%K~"u���\����t��5�ڒ�\�a�-�۠��ܳH.��R�	�����Mm����&�C��n�-��%�˝��O5�{�k�x��~�>���Xh���\��1�����xL��9�.�����Z���qU�u��r]���R�h��UUsoh�Y,�;ô�gp��%�9R����R
ޫ,�������߮LW�!�1il�ϻ��j'��`H�� dZw;��뗽�Z�q`YI:���Q�@�,�o"���]����|���U掇� P�Ca*�d�e��nue�R��	9�:�<����K�n�F`�e�m?Z��<Û�3 ���_l��6f��b�I���[F\wM�O�`���4��l�À�s���q�r�>�o[
vU�q�<�8)����u�'$�qT���>��J��1]����yB+)��`ܮ�vt���9�Z�P�V���˗M52i|�4�`Nۧ� ��8WA���D��Q�h�*G���9�b̉����4^u���Nl\�H\ӉM'fJL*[Y�T�����X��d�=�|V�ۆ�zض�Ơ�2�b��]���1Vm-�6�Xʣԛ-��
�qM*ڍ��i�u`Y�fQ��o�8�gn�W!y]/{2�\�^��t2� �#�g]I�n��L���z8˄S�4���.lo��	~��b�yVr
T3�먙s�^��&&��k����ê�EsD]ǲ�6���TZ�JO&��oT�}�ۢ�F��܂��>��O���jwv�$t�*���]�(|�Q�p�	��+�0�jЕ�='c�#��.�Tuv��`��~Z,��_a�l���]�����o��<��ꁻN�Pv�P�D�B4f܀���m=��k���(�T}+��m-u��>.}�*�*�b(�QdC�X,F�U��TQX��E�TV,Uc@kb���V�F#b0�PUAdQ+EV�Z5VVQF
�Q��F� ��La��1Q��,*"�b(������F"��R��(��-�����(���,PX�TQ�,Db
��ؘآ�b��"	-S-Ee�Pr�Q��Q�**�V
,X�V�b��-Q�(������X��Z2V�����$AE�b".P�R�AU�h��"9J�
�+*%b�V,�V1Ub�A(�Ab(� �b�Q�
(#2ՑTF�Dq��)��F"Ȫ"���+��Q��""�X(�b���1X�b""���`�
�����UX�#DV(�,V(�S-DL�������R�X*�+e��(�h�c�ŌV�TUX�"�`�UT~ >�o3�Gq�������ьGѬ5�OW]�͛���8q{Ɨ9J��{5�o"�W�ri&Z���icd���u`X�ŉ����Q<9�F�+����xd����ڼK�;E=��,āMs�]�fHn���^s�040Q����DS^�����P�3ed��P$+���-��R� ��O��`�:��T�A��B�{+��}<bgu!��;��������2tי@�������-ir�߇Du��mجv��0I�M���+�/f��zW:E}��
B����YT�3�fF��N��Did�d�-{>����X|q��pԼݪQpvN�d�o�P: ÷5�4a��-����Z!���˭ʖp�}Z��f�'wb�>�ΐ(��g���Y��>s�H
�д�8^��|�Dך��� b�Z����ī�/ц0B�n�0ߓ�N|�\#m��^ o<hR�;���}��-��G��A�^X8M��G{GU�ql�)���UD�}5�,ׄ��ϩ�C�q��ev�1�([K��mT����PA�c�g��ʕ�P�uF����E@ZJ5玉*���t��鞻�-t'/E�J�Z^�W-�^�2L�eL޹���2�Fa�jJ�����Mv���g��E��/�ƺ���3�ӳ P��x�Fyڄ,�!���-\p��h��p�7�%��7��������x�K9� c�-��ƻ4]��ޜS�Tp�Pڷ��,��/eR�Ѽ,hq&6}m�X�<��uJuu_�n�6��X  �>���p�\��v.��r���:����	��s�9�ؤzn1��P�{�s"&)D��L5�,SFj�r�.�Mq'���Yf* Bg���C����p_�n��� eE�Y�7�Of��4�<���i|��ڥ���
�
 ƪ�vyf�;�@z��naeo�8.e����]W������3�>�����E5}r�3w�L1C5w^��8w�Қ��o���<K��t�Ex�w \D�z��	��_	Sc(��J2rj���mh����	��-r�« �$KS��K�ћ��S����'�-��[��)����+�nq� D�aC��T*�2Y���~��~���`"���״��ͽ�]'��A�W�aȧ:�OJL����t�Sf]9�`�D�Ps�X6����ry{�������ǻ�OՋsj����߶P��ivX�[T��q�Xn�h�u����<�Q�8v���>�p<*Sy��7M�w$Cw��ҥ���4K;Q�Y���Y���Ԗ8�N��k�G�@ae�Ğ-���mu�n�vԳ:�y*�]®���<���YS�)X�	v��S҈�G��̾|�E�Gf�eq<�7;#}�z���p�߽�xg�h�\s'N7f��0���d�y"��"pFV��a]��\f�SEz���U�eޗ�x%��׷~Z!R���K�Qߍ�0P��Vm�"w�!���q��+ΖY�Ov���]R�=r<���G���9RQ��ܯ0��j��]���]��Mﻪp���e��LJWP�鮨��}$~SXU����4,���9=Kt�<	:<�$��0C��6l-J��0�ah��\,�QS���:]:�HKk�T�����jĞ#��@�����)�����	�,X��+�ٕ��>�{W�G�����fʘ�~��%���� a��g���a�C���+0��S_�wnfUve��)_q�R}��\�C͐����n3G��Q ��5`�����Ŕh{
�/���Ed+�a�U��y���y����ؐB��2��d@��/k#�ٔ��ݘ٬s�Q���y��"�D���ald��3K ��\�S.H٘���{��<�D�U�c��y�3�7de�%D��RH��Iً��_��,�[�Zy��(t^U!��);7�*��7@���t��>������W7������j�p�.W>G��z�/����F��c����ld!��3Rե�f�;pг���ڦ��S$,�����b������y�x_A��t�K��=.g��P�G �B-]+�ǆ�J�佃���Z|�@B�"��}�E��3>�,s_�rDU�omAf	�D����e�8ˌ#���3����.0ԇ�q34!�����Y�0v�y֩�G�V�Q��ٛNv����҇)k���H��UCSb��)uMP���ۇ�1�ad�3}��W��A�V���3�m�Y�����0���O�TB��o�k��U�u	얖�X��2��yi�Q��� 3�"Ӫc�>�52Ȋo(���U�@�G�y���wz��z��ű}�!ц���9�W�P`�)�Λt�莓|z!d�()]YΩP&n�4�{[�6��3�A�l�.�#}fptHZX��\��w0�B5�00gm*V7���J3%�
���<��^�a؄�<$Kxϱ/�ؾ���ox+�|��`�v�,��k��sH�v+��!�ʔ>�h���@�k� ywUmp�
��$�E�w�|��7���/zU�� �Mvl6l��Ǖw�������<F��YX��gYPR���1�-�
홖�N�p�m�,�����C1)VET�!�Ƹzb��Iɤ��K�so�!�@jT�,X_b�wvۅ����foh�g��a�Uh��ӂ��1	�2�W�d,����U�λ�6��1W��,F�=ǽ�G1�,C�<��&�'%@��#.���r&rz��k4OX�v4Ҍ[��Xf��s�u�Z,�])*�\����m*�)�@C��MĀѧ}��^8ȯS�K�����X�=�P��EA88TA�A���s�-��� p�:f�wʬ�� 3��K�B����^��zo`��Y/b�>L�ߴ�jw^n�5�WWZ�n�^w��\2�F���J"�/GlϮ�^��l�#���M��US�w���\�/3hv��!�V ��܉�T��4��T�^!�����e�_ ����i|hp�S%�E �7t<�z��iڽ.W���5h�ߋܘ*��-�Bkn�+Ġ��:8�e�@��0�BVU1L�24MD'Qb�K'EC�#�l�l��]��9���,Wǽ���w<b1��P4õ5�AT�WUyب ��Sl��]j�O��lM`���5�{�c!��T4n_@�WwAZ@�#�tN�[�Ï��w����^��|��$���ϖ������1u�n��yw��Xpo,����^�tX�$�*��E�\ԮU����v�z�D������[qGn�A�F�'���j�����r�����[n*�Jٗ�>��O�V� {}�w]+�yf�-RK�.�7݀M�z$���t�V�P�*�k�+3��r�޼�@W�t-,Hx��a�S�W���K(D�s�]��ܟJq�8Jig�� 7��"�g�)�Mh:�m嶩�^mT��O����vPۇդ�Z`:l�%LVz��5�P���^ͭYy�8}r�����]7�r(8�يj66;s��5�E��~�2ONn��j�VOe+/FӘӜ�|�L�[�'A88����č����j��WP����.$)bPS#-�����N��󚗺h���l
��ߓ�"����H��P�K�|���k؝���>*���m]^ki\�"E��P��
�0��r<��ZTWOq)[e�A�'���/n��\�Yt�gQ�qV����W��������i�1�%"�i�>���D�h�F�M�y��ǻ䧾}����uB%���j�?t��?g�ϕ�=�� 8:���d�?>8�&uҳ��2g�[��n�E���� �t�EN����c�gb#,Z9�f�+�3"ս{O>�ŭmA�;B���4�L���g7�dh�`q8s� ��^
$���@��)�;�Ef@�k���+�ZN�seH0���1΀O
� 0$�p��&)��4f��a9�ك~N�.�f�챚�y��*�U�!}e^�
��K5���Smf|72@���"����f񱖩���t\�ԙ�%�^ ��=X=��,����U/*��yU�ڧNr4t����;Ů�t�&��7X�ո�%H:���6S�X+��a�R�M�RT��Ɨe�:K�2/�����u��>�wٮƸ�ݭ �.��H-19꺬1��Dn)� u�v�nNs�ؖ��Xb[���koE^��: �'O7��+� ��V���獟V����y4��|,Ѓե��`X�n]��7쭝�x����(]<�=�DՅ��&NPBLt_&��⨩x�Mp��P��߈����/��,P�_m2�' �fUn�&�x�����b�yh�Y*[�ǁF�%���#K�J���[�[��n��r�W��\*��/bI��uc�(��9���C�Q`,��33���O����\,O�J��#TK���pST�#�U��hG,���V�X��\����ڴ�[��g��5S��9�Ym��$t�su����{��6mGn"yj�(B�����^1;��j���t$T�$�nq���MřwW��1T����]S#��`T�[�d��8�ͩ =Ю�Ҭ����t=���0��sޞF���V���@��p�*ܕJ�i�����n,�>�������:�'�l�C�ܲb�D���dMH��gAFZ���=ig�B�λ�亞��Syƶ,|)��e{�u;��J%LCRX�{+��J1�;-�M��w{6�6z�S�cFd���j����L��ŀ%��"�UI1��R%jYx��ܾ�^�.%�H��OM�A魃띐!LFˮ�=*g=.pPb���;�1�E����:�f�4��+��� "9����ѼS���K��)f��S�w��B�^��w��s��r�>B�u/i��b�(e�)�g�Ps��XQ�.���*΍�%=��.쯽���r�%u(� ��;F�0�¦7vA�8j0� ���M��H�k4��֞�s��+Y���>�3�Ьx�:�A:ty�N�T붢�uk�>ag��˳�V_���K�`�����}6"je�����v����ؕgm�	���~ݗk�v��~ۣ�ޠA���&��;����g:W�?{��lc�
9f��y�����k�)0պ��2SQr'.Ҳ�+-�ϟ[z�;!�c^�cV �B�cG|ӎ��w2\R�/�u���F�m��4��v8	��;ݪ�Tt��G��\�X#_�s�����.�Vj�5�^���)A�L��ni�	��_\��!�8$%sK)b��Kۊ�.{Qq�~��0�b�������&-d#⓬�T��'��4��=�t��v$�,��ŗwc)����{{i@�ˋ���>+|�`�0�	j
�:��A�U���p�R�36T�fnvZ��Js�4f��;�%s<�`\ ��=^K��e 1��/�j�#��C�-���JC�_�Tp�M�m?oq��#��rr�n\�9* _�����y#57��Q�#8^�	�RR�6pG
�څs0��R���;�������1W�'i{eV<P�-�����b��[^G:�6*Wa�ЧŎ<"c���GezS9�WU|\r�{��SjF^Ĝ3Xq�u��y����W�K�P��K%ה�&K�(�c�}�m�}�_�rn6�.x��D�E��oO��Qף�`��Ⴤ,��.f�`Y�i�F�v�c��ѭ��u=����3�Z��,��CKq�8k��|9�D�`b�E�&��vt��o98�l&is�J�5��qØ�w�N7+��.�X�x���Ge�%bَQ��[�N�e=�bi�J��N=����#��6�H-�{���?pp ��肔��r���>7��yxu�#U'�v�f�Ӯ�6��q�҄��%�E��7t=M�TCiueQ��;Z�f�ɒ9#=��5ip4{0M�a���R��Y��sP����$p��n��F�K�����@,�����ps'Y
��8T	�Ҩ)�٠���Q����C�l�{��.��� 9�U�,�MX0�<φ�������UY��u���4g�w��`���u[��]����xn���mi~���4�{�Y���1l^غ�u2��V:�'�o��q�gz�V-�p��*H�zV�3_V��i�߇9ך*��]!U�-�/�y��swKģ�FgL��Hq�x��<=W<4/Y�^)$�3˧�`��c=Y�:����ű���i��19S	y*�e3������ޛ��.$)=���ɉ���=�jk o���VF+�����M3b69Oq�R=7�a�nzW��B��ɢssD,��Z�֊�*��ȡY�vS	�RN)+~���Pf՜�܋�N1�
�t|�V�`���q���������؄p� ,!Ӧ,h{���N�¤*�/�#u���S�C,QB��Vɽ'D ��}��.��L�XD1m�W�������0��{��m,��J�ݺ���P�v�
Mn���K%��4���kѷHG��O����fF�΢q�U�_&CE�ɭ�hN#ZKq�%Ƶ���Z��m'}!<�+�Nǈ��R�,%���q�Ԧ��9Us:JV��C?^Ib�t����f�18p.�)�����!�-]����p�w$�-��q��:q/F��}c�p鵢�R���K6$/UYt���V�r���X��p������<�;��U�9kɕ�a��1J0�ClޅH\�NmSk�q ���4�3Ok�Qd;�W݇�Iw���9zQ���j��(4�7(��"��4���:!tX���-�,l�:\7'���������|�+�b�m�=ԅ;�g$ɖ)���'$�*N�K_�v�92��������ձ����S����Y|���=�y�*k�U�ffl2��IB�`�2��w �3��<�&s�9X��8���1�;;��R�M������t��n܊Wfr�Bx������[�amݍ�r*,���3�*�P<!�n*d�Ҫܓ�U�h�Bb<���`�OXq`�;��5z���p���i�2��\Ϟ|��"[�9Z�*t���`X!ѽO-�
���1�ڌ������N��z�o=�4�Q��Kqى
�I�d��-T�g �H���D<f-�EtJ�1)�k���I�d�C$�m8E�r1`��HY���:��,�^ل�r.)������$���X}�X254�M1z�|qtʎ	._,�x��a�t1�Fp����n��OG�sA��	�L7��Q�l�8�˘4;dҺ��&�2Tt�L�Z�����<B�����A��<O9�L���Iؽ�=��(�
�@<Oa��A�f��4�/���Fdng�H�}QܙMD�!��N�����o����kj�`�:s��t���v�q��R݉�#l<D=�X)��$��+	P��2�r�h���^.B�T�D�����Pa�E'�����JDz��]�.����_K:��Jp���S�i�F�r|���%��@�!��d�
�=)Z�GVU��,�IZ�i�z�TLG���#ŌD��p���X�te�����eˎ8��8��% �Kj@�ԱV���Y��K��eP�B8�-�0�@C�ڱE׳y�l7��DV(���Q1U*(���AQE��j�*�Ŷ��QQ��11b"�+DV*����DDTb,S-� �D`��1A����U娈 ���"6+.�F"�ciX�ƣb����0�(���7-UX�-��Z�.4V(��W)U����QQF"�QDDd`��k*5�`��)�
��(*�(��X��b�i*.�TU`�H�\jĕDU�`���ƵE5QC,��,`���DX�X��Q�b*ŊV�E�E�(�*�Z�UJ��T��QAUQUQb��PX����QDG(U��U"���*
�LJ"#cbDQQ����#�bUiC�e��Kh�@Uխ���Tb�E�1TX�)��EQDE�1��fKZ>������9o�������c;�;���9��2�:�r�2w�:��n�aᵮ�鄓���Ғ��e��ջ��ǫs��nȷ`��D q�C�`T�P�G��(t��JR����s���I��Y{�7����~��c]Q��5HR��U�o���˭�u|���k.�7@�X\x�O\?:���)G��T%/oX�Tj��bˉ &m�B�S�F;+1gD�o�F�㉍�VM#q�<�9`��x�w"���|!��}���e���9�VnD�(9���Ո�=�(n�!�C�?PT�s�« � KS����x�o��k����WU����tU9Zj���La���B�TG,���#�P�Y��]�mƦ^/�֦�=w�t��.�������� ����T�[7�B��p�	�1P��ә��	��/��n�nK���^[�W��%H:�yfJ��S�]
˜�5J��qC���Zt���Xk޷<4r�L�Q3���UG����V5���h`�2��J��JL��E����O���'6,�oH��Q�J��z*�^܎�m�{+��"�NL&�mE2:���kCz��95h��ix�a�g�J�U��Ї+���ōP�i���7�U�q�V��5����&���	}�*�w�1�{�w�W�)F9H�����x@�h�NM�3n�\rĩ��5��I��2�Uc�MD�ٹ.:�Hk�op� keEfB`]t��ח
|�pCΏ%���g:�B����%x#E�vQ�kUp�+"'Y��w������9�3mg:���#� �+�N�R���
��bo�qdg�f��G�[��W�P��ٚ֕W��m�d�;��^��!qCb���ą��[�1�t�rǄ4j��\��wur`ի��NQ���|H5s.U0[K�)Ɵ��w�ꈩ�_�m>΂^>�Yf]ߣk�hٚ�j��5{*>����QyHX%��PTmu�#�j�=��9�C�ꭶ��j�����^n'CY�����<�d�(!t�l���Pƛ���Bv�5wrG�G��='�[0�'i����z��6ܻ26�Xc�)�Qf@�g�٣�x�{�	"�T�h�HLX�f�n�5�Rc�x(�Y���f��绳(�@L�!� O�yr%L� �nv/�8�*�r#~�-l�٩��pzk`ŉ� B��]6zT�K���S�6�}D�3-{��r�F�q�Dz�� "*L)�[��86���:�څTDO��c����r:NMY����g\z�ɹZ�&�>ꧦ�Q_z���/�wȦ��,+3��i/=����1�����M��[�����q^mم-��3_)�.�0��}��1������t��/9e׹�-�h㽮q^�-�C�ܗВ����s�Ӗzq����R�5Z+e��[P(�`�!��f�;�pf���,E��n%�UG=Xi�qx3ϥ̏� � ]{�aIW�ꆴ&��ZM!VdG	N�;"Ф�v�7�J�H2�[]��}����
��\�(_L�6����͵�Vr�l4	Ӛ�TN�1yP�w�4�v1��Χ+'����(��q������Љ�y��M��"7�:2��jn�^f"��j�\e��b5S�;�`g�P`ה��M����Ƭ��F6��\����ϻ_;�j�o���v|r\,O��F%���CE:�O��BӚX��\��ɰ� ��C��d7�c,W�a�-d#⓬	.L�G���eyn+��A���{����I�á���yH;�"�ń"�1D�P0��(~�)]8��FW]���f�a�.�G]�Ѝ�n�E���;�κ�c#�8)	s(Ǫ �P�NE�+s.�SH�彌=PEJ*lO�1B9�;�R8�q�@�AҔ<`^���"���CȽZ��l����geN7c��4۝u �x����4`D^-I:!����A�qƯ�(S=������F�oi��B�zC�j��/&�f=�\�u����)��uoJm��{��������K�[�`��A,�܁�|���=�A�����L�w��]/�+u�����E,E�@��Cw�Bj�e��Z�r��1�y[OR׉c�b�[ً�x�.���U�/ȀNmh��S�y��8لL<+��yƔ�"E�l��i6	�`#�w`��q혟*���8�٬�~�(5�Dz�=(3�<�eOk̹�X1Ȼ��(���I��[��{_	w~����w��TlEj�6�%��n�a�u��5�z����1T;{�=�x89>�!�=ͩ݁��L
�@p�Q�Z��c��ye�Ba���ͮI��񑻓D��ʪ� 08�[�7'n�,|ǹJK\�vjǆ�3���^�Ởsq��}�N�F��=K�Ҵ���jE��, ]CwC�к�6�VU�,%qW�c���1�<�{�ٶ��7�wKB��f��
�fq�Ct�a��N��,��Р�kF^-ƦvW$��2G��8]�4�6���U�5�m󡦝�Zd ��X��G$ob٭\��ܲ�k�;��VNa��L����/�N�Qc�� `Z|�v� 7};׫�k�)/��Y���m�5����OB�k�K��<�ٜ�Js玘�>��xʿ 7����*�ӇYJv��;�i��+c-+���\���:��3@�w�aU���>�缺l�"��\z]�V+h\����n6��� ��תo��x����m���8}�٬���\e��dp�� !A
��B�̈8�V1smt[�x�XO�+r��%��x���0�Ni����U|td@n���,�Ъ�;�����S�<��<�^��2ke�`���\���o���Q��F�L�[wO&��>���x��V��Ƒ#˸� l�uJ����:�����`��[�V)��#8œ��X�F��St�n�OV�tC=HFi���5���T�<%�p��|~��u���м��>T��h��]_U����	��Va����R�Ь *6�Q�w�:�X��5���XSgL���Ɠ��D�Uϓ�hJ�1�)�� ��
_+씃��*��=�3����4�D��!��9KQtƁe��[� �WC3a5�ki��XZ{%�ȼ�z����}H;��
���*,D���@7�`��D	ja���x���,��9���F
4���u`��՞�x���i3�`u҅Q�K4>@��CU_ 2W��������\�M�ri���ͬ�ڱ.�]m���������q��״զl������3An`>�2�Ǔ�a|��ū]@R����k�ڽS����=:����)p�}���ֲz�3%}��ݳ*�6����Θ�&��7�s�G��i��2��$z����W�ez�Ɗ����&z�U
/|k��7ʺֿ9��2��x�4,4���ڭ%H?UW�d�Xx�W[nĳ���{�~��1�iļ����X�t_��t_��R��!�`�K�E�O]�x�U����f��b���ko�.�W��SUۄvb�@P���D�]Q���O6�R�k����<'N�:�eB2�H����RgrH�cԗ:0�M��=�:��� tF�B*��J�F]��-�!-�
���!��Mwu��nB�~��ø0u͂)�2��$g��Skqdr�c\�Œ�cq�+@�"�\9�,3G&8A� ����`W��&�W������{j�.z>�kQ.�8ɬ�L\�z�L������Y�4lBG� �b�!�-�:sљ]?d�K$�tHUf�]��{f#&��"D�1���Hۙp"���A�X@�(CA칷149��{T�*s��Y��:6.hp�BrɊ�����*���_��q���3�u�g�P�gq��"qq�D�#���de�y�{�\T�:H�}فۮ�9��"h�o��**�o}嘨m���}ի)	x�hյ�.�>��k	uwVF�	݋NK�gfܴ�BTSka�6t��W���N_g�C����3Z�bk���T����sݙg2j�]F�����hH�w�Dam1:[vۗfFþ��d
e.��3�k
��!�g�����̃����ȘB&5�C93�ҙ��l [}r4�
��-�Qr�f�<���� ��\٦+�����U<|=���j���K������Y��
k�"����MfU��~����Ӓ/ҩ �!5��6\��7�C��3UQ2�@�d��}Ĥݚ��^��*�*�ܫ!�N��Їp�!Yb7Ѫpn���\_Vr���2\g�:m��tK�H���
K���5���XL�]Dh^�P�
HWV�i<��0��;W�u�.4�:x��e��f�Uz]�=�l���z:3'�۪!�o=Ț"��l^K�[�K�\p�����½m[�>��
�J 1,�UL!���Kˢ"���O��s�[�z�"���F%��
��ʋ(�p"C��p+�(0iO�t�wGz�K���׉�s{�z�v���m�&Fx�lO����$4S�������G��u��>�^)9���n\��^�}���:��%+6����rU�3�{\G1�J�4!��އ{j�s���
VT��Y����>.>1Ō�]�fK�U��\�Z��X�{K�z�Z�*���UZ�o�*p�*��:ĩ�&wp�!ξ�����x$�;8�|c�gt¶��QRo�/9��s3�:��wvp@}=��sal*#ܸ:���t��z�mv��i�YH;Uv�_P�艋�G
��h�
�n�q�&B�lQ����]�T���5Lmѓ�R��܉m�~4�����Y(R��H����X���>˔#Z4:���bD.s�V�X�@��)A��&����1/e�,�R�]gq���	�y)y����"a�\^��5�3_l�~8m�Y����R94�����Vy�#�1>U:='[5�
�` �m�)���b��4�uu*y����N�9� T .,���2� �@����ֶ�gZ:f;��h+���Q��4L���(Ys���T��́p�����
5�㮈�^��B����+V�8���h?G���wr�Ì���S�|&��;�7J�ROM��0g�7YY̳.֋�[�O#�:ɓ	�]2Y�E��7v=M�>�+K��g��?*��0���4�̾y�k+�[}���;N���T����l�h�b��8�ɷ�[�"Ԧ�3M��[C_M �Z� ���ѵκ��u�9�a��/F�t���][u������k�5'����d�ۄ�c�������ˡ2������ӷ�7,4�������ܘ*ٱbǇ�ʹ]APLïq�B�vh0��pmk�(�������|��2�'�$�!��5�|��hgb3eQ*�O�<s�����ۙ�ef��[�w=c��͈c�0���捗]�:A�*�3�tfrEF�8p��[���C��E��W�G���Yaj��M�p����k��ZoΧ�U91!�L�/�WL&s@��T"b;'x�qL�yH+.�o�I��w�3J�2\UW5{eܧ�q���$�[B�{��Ɔ�Yʘњ`�شt��;���	��AI�g���ڰ�vf�{/�UOּ*�K�P�{y_��A�ڔ+��~��L�ޘxe�T ��Nf�i����[�������cQ!M3H ���@�SA�/`�IMŹ��.˺�_3�q��<[�<�N6�� u8�Wp���{H,�����Y����Y�5�::���B�aL�w��e��*��pC�d���UP��F���^h�좰���C����@v'S�(
�|z�)ܢݼ��.���jL��AK���
�c4��E_�j�皑�h�paR��o�(��n����ǻV;Ix�9��j�/4���
t�홷�c�rcu����l��,���!���,O&�)��m
V������{6�I�6��~!�	eHl�4�Nb6�;�����3��ڥdv.��6f5@�v���NY�ޣ�εm��o˥[mW
�[i�w����V��H���POHG��ބ�Z�"��vU���bc/S��'���^^^�ÑX�Q�0��H0�ĉ�s�
l�� ]�(�km]���q'j�
�6�<:1Fϰ���
��f�>@��fC�nc��i<l[�ɢ�=�C�<Q�k�U%x�Ct�`�޾J�F�A�u!��#`cN}Eu��e�臛�^�wuO��=�1�1%Hmx�Ҽ�%z�<x+�P8o�>�2���856�eU�m�\�4� �hzbVxZ�|Ϯ��Ƴ�Hb�܀�;樊��Um��*i�>��%�4�{�r��>uҍ�@���4�1l��t���cq�I�Õ�l�w噀��*����r�/�j\»2�ΕA!��tF�BB�����];?tZ �K �\�[�� �.�DU�32�Ԋc��è�F�Qd>S�B��b�G�bn�&v*�5�5]��[���M�^窳��&���i�!�P��Qz��{y<�2'���.,�Ǣ`ٝ��S�N�WF랁W),�6]29��;�����F��ɤ��o���ő�W��(�J�A�l�E!-�*xuW5osN�*�d�f�Jۮ�&�Om|�]9�)*O�v�v.�\�#�oGMb���*�YL���F��
�XBa�Xu�]�b�[��-���A��Hs4%�T�5`��j��ڜ)#NS��e>�C��8��ҕ�88�"4c��Ot�Tq��m"{וٹ�"���Eʐ�$0�آ��(2��[���㦯���`�=9��:R��]3�3U�nuF��7��W�<<�� � �ɜe����1�����[�T;�U����e԰Ls�1;!(�]��ِQ��Z����M�j*V��
�2�~�{h��&PB�B2���s��Ωi�o�K��v��F��E�U�s/p k�n�,�KZ��F�a��d,�cVV�X �~R���c�l�T7�X\5ki^�]l��iu��V$�s��vjcn��L�����-+�znz�DTԻeWiS����JI��J�q����zYY��Uz�H�A�پc�M���С]M�ґMMp���[mK_j�_]���.T+Z�1������g��|�eMHM�n� �+V�pX��#3Z�:��(�Ş=���0W
�g3.Ʃ��ԫ���*�^s���9�l;8�����S�
|��,RjCE��i�إ-�F�Q7ڮ��G�n�k�v�"R�,L�Ӕ��y�)Bb�\�$��ֶ�
�Ճ�c��hRh��Y��Rl�.ƈ[�ia�����u�ǉQ��$d�6����@"�瀐�4�fA���c3!����,�XnS�����2b�]��#����
�X.J�x����<'ψ	f��ґ����cl�bX�s�� -�W���}��jU	˭/�4�{�&Wq��jc���C�Ō�&1KB�GI~F�Nt���	犧�X��s�̆�M��3�5 Hp�>_T��BS�V������1+�ۮK]�*����X��q�B;�7���\�f��[{o���i1�6�f��9���cbt N��L���mż�u'�uhX�y��L���V[S���V�gJ�b�@�@�d��^���lp93"�æ���F6|�n��W$����)�B��T$�;W
Ka���T1��>{j���ˏ@���mD��.�R�����tPsmG�QEJ�b��(�DO�"�
 ���T�TQZ0+L�Qb�*�V��(���5b�������V("�**+�c���TQTF*�EY��T4�0ƨ�؊1UUrʋQT��Abȩ��Q�
��@b��2+QA@E��
(�QQA`��YAQ�D��QQ"(�#5QTUEADueQUm��h*�
���QV(���H�i4Ɉ��*�MV*���TTDUX��"��4�(��@QAUQ� ���iX��M4]Z�"�Eb�*++cDPU#U�QF1ƈ��Q��U\j*��EQPb��m*#�dV(�����b���m,T*VF"+�(��Eb1�/˺���r�އ�/g#�Ok��
O&$�j=W0�3�'G��g���N�p�2�9j���J�̏f�̔�=�K�E��u�]�'��t�Aܪ��p뢙�I��G�x@B����JX�ZS�w��9;<��
k�{�QE�ɂ�����
�3���ф���|�f�6�1*�jh��s!�=��k�|{LE�7LC<z�Q���H�Tȍ�@W�M�@�it���Yn(����9u��&ku]{k�_��*!��1�QsC��9d�E�JGI�UrRg��'g���g�ݑ� h�3<�bD73va(��<��{�݁�n�C��|R{Z��8��w�G��Cf��h����8ez2&�{0�r����S0s��Ļ:ZF�L�O����9jG���"RU]��_��-�D#�x\�����4!Ll��}��&�em٬�JV�!L��g Pb�]M�z�b���k׊�*^[e�W���_m�zn���{ȋ�hX���.�.ȇ`a��MPns�Ӽ��P$�0Aԇ�@˯*�� tr����u ��x�c:.���(l�%dÒ��m
�b�݄�+B�̕��G�F&z�yc��;��&	���F�^��ژ�WQ��ז����
�1ɿ;ԠV��]�L�D鰭R;��ݔ����X�k��]E�Dpk�`�i���aZ�)��=�-��޺���oH,�l�wn���B�/tT��J�B�L4�9��.M����ͱu8Wyf ��Pt��OM2��t�3p��έ��d�O�����{]�.�7����Nഥ`^z����u��ENVM��{j	�����^�a�~�+��0���y͋�"��#o�"}��;oF�g���b����+�](0F4�eb���.O���f+�����o�"��,@����;2�Խ�������],MD�.�gh�����NV�`�����Y(����F-�VOYB��_N�u*Zх�B�=Z:����b-�g@c����B8E#a�D��J��,P�y7+���F���a� 9S��d�	XX�Su�{K�e�3��_��Qf!#�d�I�p���X��y������̘w ~��zP�\�>��x?�9��/r0Bg���H��2���J
�CY,��r��v��F8������+. �t��,��kv�`$>�r/��1���52.�<��vU���ؽ�~;�6�h�LO�\����V�d�轂��.�ء�X��嶉Uu��7����K�>Kྺ4�m�՚,k��]Cb��#�VauZ}��D���k���=n�pi3Y�d�l�]�w�.�xj�2�i�@���������C�3{l.�9���]���@����8SiXĭ�eq;�m=ԥ;��a\&XŴ�)������ ^�� $ھ���d��l���+9ț�.=ٖ%J�]r��,xX�c���uq�K�qk2�p1PY��v����: �>0x=���'���b�R��y*eާ]�����'��(l>LߥM�^n��LW�B��j� -`��{��s<�C�/��Kg®��E�L�[�Y�˞C z�B�^k����O ��Y7�rc��N��K2�~�a���rj��L&f8�B��%��, [u#���G��;��	������@Ҕ.%�9r�С�pF��cE{
�z�@#Y�Q�a
��LS"�ژ9��xZ�.� 9QF�	�4��"L���fNj�25�u�@g��j�W�,W��>���S)�����1���a�d��Rpה�D��К²F���8��9a>�˶ZZ��V-��?s�=e�<�Q�ǂ����WYu����SX��cn �jA�7J�[�����"&7'Y��t�iܠ��(k��x, G����{���O<M�*�~�3�����FV�yu4�_�c��eHCQ��;�*h�ҫ�L���G��ӷ�Q��!�%(�^�Ӈh�oSt���21
�t;��9���&b�[�[���[�Z����L��_[ڶ;Z��s�����a%�@�趇U�.lR�C�
�_S�B^Hæ;z��N}�Ia
�1���͡3j��X�Rt��
j� ]3�h����ՔBJX��wIE5���wS�C�;܃}x���,�P�9DEE��0ʉ��@����~̔;N�Y�i��ÕBm�l�q��D��>���%;J���sNL_���d��W�3�	9(A���cĞ�G�u�]��{[���~�����*�O�2� 8KE�U��oc�2�nΑ�B또��9�a�����d�<����Zk$DK4��%\�Ԯ���v�\��b١���,C����f����b�� &�8TȪ�t�TIy̫��FqQ�Hq�0ɧT�#3�M٢�O�4���YA�P�U�K&��<V�*�J*R��*���x'����~灊2�{I1W�+]ٺ��<v�p�S�T���o�A�fj��ď�E)@��Os�g�Ż��s�{m�i�CJ���%z�ǂ����%w�%�;�]7g�=C�	�)ŷ��.I�xv�5��yFb�b���;��T�I{Wv�kv>��>ѴV4�}�b� mn�����=����n�������1��mE�R9�<���p��n�ĉy����MR��Cl�v�˞�d$~���)���/�[�Ɲ������VX�[T���ck�^,W��7A��.���J���u�X�iP������P�@����D
F-��J^�����b���	�m��n�t�Iz�~�y�y�+�j�*)��~��R��U��t(��C
5��s�U��W�4��_K����({�/
*��D����R���z0�iN{�����>���v�xso0=�S��"I�cԴ�O<Ӯ���*��x������������l&�6�1�]\�R��tc��95X5�����"�k�q�(�rɂ*�_���Y�+�>�C{QY�Ub�Yy��q�[�Q�Vq�%9|xf��ǳf#&�!�q�*a�B)�p3���6`�p����#�Α�.�p�����ct�i��N������EP��5"I|f��i�ɏ��3���{�](��'�.���k�黳]>��<��y�[��D����V@�<F)�Mp=*�C��t�]�rz�,𑳋���.���&���~=)�#�̭|��^�KN&�:�|�D�9ۜy�9�par�$�J���xfo�z?/�M�Q��j�{�AW�nP5��˅�Uc��.��fVV��v�z�Bo��I)�AeޮaUѡݮbC4v�:��J��k�86�����:ev��lu.�l�(zGs�ֹfg>f��ՔQ� ~�Z�y/"/䪻�x����[C)�.b��i}a
���IK=Z�������� &�rE�PE";kˬ��^
���j�`��#f��� 9�zn�?uQ�b�r���dXo�j
6,-H}$��X�-�0.7��dѹ˝C�]zLV3V����=k���dÒ����4+���B��f6țE�v��c�m��$YW��]��͜	3����e����WL�[��IM�s;�	��m�]�N�]324ɷ�t��yVWY�Xo���P&8��v��v �8wt�@MEۥ���ݢP��dW���̺�Ȱ��b|��f0(��!�n��Ի�1���r0��xv��^^X��'���t��9猔-:��FJ���U8F��>)��� �]Zmh�x6���X!���;iq�B\)\���}Z!��錦����Ğ<��Y�݉I)�������SQ�3������R��qBӷ唃�*�B.8ń"��(�j�@\٣������]v<F�Nޕ�*���_Z�VJ�������psy�oe,�	}دMp�G]�M��}�*���zx�cs{ƤԞP[��y�d���L�vX\�ex�;���8v@s����7���_b�?uNԤ酙պ��Μ���:���������)��T��]�����c"\MK���粧)�E�̰:�O\G^1J!�Z"M���K������Uj򭼫ΣT�Sң�ڦ������{ou1��o��W�@puf�x�j�v<����§v�_�a��9yl�=��&E��#j���끦�nl]Qg�����C�[5�
�` �mQ��ӏ�T��k�@����a�<2���e�� \i�O~ʨ�L2/{�����w7x�f��7�4O9D�vJO�7�66� 4�`��&5#7��x�QuSwG+1 ���΂!�z�Q��<4!y�D�^�&�N@���n\�a�w"t&��i�$l>;������o"�*d�D��y��,�V�)8�9���	OL�i -:��4����P��7�ԣNe�,�W
�*64TaA��� �fG�.���ޱn{5����M
����5��h����0\����ps��C4�xk �Gk���yC��^MT�Z.��K���XE=t�{>��T�J4u�Akb){�>ۙ�'�y/y��%�������ʢ��Ҷ)�kΒM���mG��᝾���vs�j#)ӽ��5�ļk\�B��x��O-Y��ir��L�ӈ.s��S�Q��^o�f�c�ڸu�,6l�þu')�0����ᬫ\jt�W��Xv}��>�{\GJ���AꖲpF�ʞ7��x��FUEvI=����v�^6�cغ�T�f��@�}R"t�>��)3L�3���W�I�kf CrC�"�έ��ٰ̮��5��F^�yu5_�c��T�5���xྐྵ�ʪ��vڃI���#:S9�w cL��R�U�eX':��|��0��bW/
guN���
곉p����+�=��<U���$HR���Uz1�S�M�VI	)�f�3P%�ql�XwH���#y�w!�"�D����
����GY���<3D��[z�^x��$B�e��n��d�,k_Eh/W��c�dĠ�� �T;���s�9�bz���6=ö�l�44z	c	��#}��M�*���A��@�ᆞIʾ��k�j�E:�:�!(owJ��ʼ)���pySr �X�re������4�O�y�#��t7���L�Ã'���z�/�Xt�
�fwJ��u�J��x�iY0*�6m`����'w�����@�eh=rC}9h�˸�8�0�1��<��չ��M�j��mvpUξ�D�P6�d�شså��np9�Df;`������x�hBE��P�[
�u	�Pw\ŋ�@O\�\M�\T6n��U��MfUހ�D	Na��G�NՄ2�_�9�5~���T@A�u
���,U_�᜵bI��n��e��t��,o�eQA����&�4�gk0�)��=�Ɠ8_A�j���/�]T�v0���w�|9u��H�U�6.�X�������i*A׍3�s�p�¶�BVT�o+��d�$W}<:oz�G�ixX�ڥE����]�(_��|��'l�wzD��Rb\t�0�-��R;��}�Ȁ�S0���r�����b[��;���W�fN�$��� ���*��̱(d�àu��*�C��E*f;L3RR�쵩���l����-�7���fZ���T��H�0��SVe�G�59��1�ɝ�=�e�M�I��3����i��vH�F�U
k� �3<=^���j�� ibb!$痧b��Y�N2�z+�:��v�NQ�m�&�)UU_=��p��7v�����)�qƹ�#G�( �zV���r�,�K3 ��h�^�k;�̇��]�8�&o\�#��Bp��-[T���l�\��n$�QcFr����d��jEq�{ԹL{�8��;��1V8NOB�ܯ�5�,��i;Ye���n�����F>�Oì�R�K}C�4*�W��C�3eL\=hE�9����Om%�k׶WWf�>Wd	O�q�܍حf�4�N��L���l�`	��ߟf�'B��ox��P�9*�ݻ�b�ؐ�J� i�@�lM���3ܱ&t�N��M[��1�Z�"�$���EPƱs4a�7H,���:��`BUc���[���K����Nxl�r�*�Fd�. JM�M�j"f!uD3^L�V�ȔoMaA����IU�SR����Ģ�+�R�9=!�ҧ C �j���#I�
���X�=ml/v����K�ޅzfl2z�f�aZ�Ԫ����΂s��42�p(�s��.(�>=4!��c=�;���1n*���Ⱥ/
�l�A���ť�t"���¶�`��(RYtJ&h��)vuk��.Hy���R5!�
�x�UV�	��e�&��]U�v���v"ot�8!��K����p�r��T����Z������̴���
��K�z��؜?�B����$�� �$����$�IO�H@�hB��@�$��	!I��B�� �$��H@�hB��IJ��$��$ I?�	!I��IO��	!I��IO�H@��	!I���$���
�2���r��Y��������>�����q���@          
  P ��)
D�%
�Z�Ѫ)Ca�Q* �<ܨ�
�URJ��
�PR�R���� $��R/ �.ڨ��ى�0Ś��J�1
҅)���� �'Y!E�EV�ZB�a&����U�%UJ��  8�"I#�T�(��)��-d&�T�#D�l�p  �E �Ȣ�8 v�z  q    ��  "ŃC�΂��sawB�UEP, ��S n�l]��ݦ�\w
�&���;���f��q������� 7i�+��*��IUŕ˶V�sp���� �--�.��v)��!R�@Xv����2n���Km+&N�77E�-Qل��Jm��
�T�� �U�d�� ��R٪�J�Z�IT �(���$lMR�-(eV��P@E-QH� '(�
���V�e-����!U�(�<�   �jz�R�J0hd`&##����JRU	���� bhD�hx������=CA�M�!��J�  4     i��&�&	��0`��$�I��������C i�����ݳѾw��xZ�[��u�ׅ�V��p�[`�
�5��I:"���?xQ�A:�DTh̄P+��}?V?S�I�\�PD0#P@&~R���D�.HF!K�F�;m�s�[��q���n�*8J�ZJ�?-r��m�����5�{��Q���O��2���{n��c�iCteìp�:t��r�yh����"��b��eO˽gR]������D�d��'��)�����ɢ@�1�ʹ�v ��qc�����(��W�͕B�#��@?L�|�N ��sq��ڻ�'�q�g�����v��j޻V:K��X�mγqv7�oIN>Si�$k�-��<������7�Me�х��'c�ƞW+���D����wt{�uv��a5jޮ�t�9t>3c��\�.'�wV3�C`W6D�6H*���
G']�@Ȱ��@{�=��)|�1��6]PN�)��sQӖ=�`ї���Y1�:D��O�A[ñ+�uںt�,n��,_r��(�uG��t�Z�v��(��| �j��1�[���e�4�X����y'=�9��������<R �m�F�/,Ŕ�ܖ������h��<+O.I��4q�3KV�v�x۽T��*�j��{;!�K�%����>1����]����Jp���T�zJ姨��ۡ�Դ��7h;�f�q��r6En
��r��w�_]`�Y����ѯY�F��\�|�/�+��!)-�rȻI����ئp�����5�7*}��K053�Ųܸ'G���'��Ú5v&�+@3���uq[�ax����v��z�d�躗��a���U"x��{��#��#T�t\������|v�Sf+0�CN���j��v,����p�γd[vqۈpZto����i�p59�n���û��h�����l	����zi
d��o(Mk9tS���	 ���'f�݁��������wb�D�,��,����V�\^�繽���r�����[^�3Z�Jĥ�!u�8������@A;S�����F�PPeI௖L-�K�N�e؝ҷx8��F3s�f�g�Ⳳ�v���b�@��-%{2�'�b��-h�d1��eBF�O�
��ZI�)�]Tഩ���0�|nl����⏠��Y����I���V���Ӳ���uhjS��(:tp	e�°	�8�]�s��(F��V0�! ft���i�[�r��D;��N��j�Gm�݉+��a�ށ�Û�am�8�MF���=ucI>���xw;���{��Nl���qw��G7���[]췴S��Flyb���!t9o\[��|b�K춮�;������;��&����m���	�r�� ؛�4�j]�X�
3���O#upz����{j"^�l�cY�����E�8��Vѥ��.k���`�sv���Dd�ͦ�`dn��r�7M�&�]vY��<ج}�B�L�ݺ��x��8�5�c�Z������[qī�Gp�A=��dΊ���NX�i(9b�WǕAÃyב�ڞFi:yweuC����~{�4���_^wP'tv淌����T��D�1�Mh�9fK�� i|wS�8k�
ke�lq́�e��	ιy�Wo[�t\т��ջ�D�S21!�_ix6���3�_vG!�� U�Fs9� n��<����Z�rYJf*w_f�ߩ��M ��4��$,x�Jn�p����<��)��e�?\\7s�vF4�J�3�O��
р��5:m��gL��,��~���C8\�ѓ�y�7�#�ph�`�^g4jz��"_�������w�+�f<�{���d��o�JH·雁d�'ę&@6�}6{L�ݮ�Nä���I����
H��c��n�Wi�i��.��W��c(���}7��T�� �ahB=�3h���;z�-�����{kM�㕵�m�;-�5��Eُz�
^���Y�'G���~��c�Z�<�\�Ev��s�w��T;��d�&��#�&��oݦv�ׁ[�+Se�&����\Ɩ���x�rm(���N6م��KH&
3wxd:[<3�p�ob,��Rc�������L����9�d�Ի���u������k�\��g2��" ԟ.U��)�.����u��;V���t��n.V�S�&v�լ4�9��o�k��*�x�8t��u��8#����E��٤�����X�'�V��XV#���N�ŎE��9�rh��)zv�YsP�QuAL�V�K�(7c�S�"�c����U���LT�3(Z�{�i2�>�Q0䚞�^�� 4��3ٻ�z�.e�l
�,�B� _,�
��e�q���Gs�ٚ�n1�[�s�x�wJ3{R7q!j���0J3nN=�%�N�uL�7)Ox<gc�T�E�-(��ER�5�)
�m�,��:-;{�Ò��'�ӓ�]a���!�4�U�e�o�/��3���-E�{��N�B��F�c�s�����S�_;�I�q���������G.�YHbw��f;�α~�"u<��꜂8��С�jY�M:#T��=�mE��,"N2�Ek@���L�/�W4��b*�a����c���w�J͓��D4�J&���y`��˻�����\�Wcʀ�Ǩ�]I�l�I賓-!	3��_&�޴��cp'Z��ɛ��Gq&:��;En�S������9^��;��b�|�N��e�g3��grg8���ܤ����J7[�g��'�/㮰��8*㫪Rۧ:����cO&���In��,l�5@xFV�xv�w��L�wX�פ����K]B0x�ܮ���Vp��WD��:(Ψ"�E�ֽJ�m�ov��}W�g.���{��*�f�<���'B탎1�k+V�p�k�*��[�ŭPЙ�t�� .J=E���F�w�cˡ���rۓqb�Y~ځ��7jĢ��Z ��v��0m�#$��hp��&oP7;��k�=sV%k���hvʟu���f�n�k��X͹u���зv뀘D�(]l��1���d3������;I���-F=bh�.=����rf�Ϋ�c�<5� ��������ܢzΔk9V
aӯ5v1k[5|z� l�vF���߾���V`����=�6$L?��U#�O�?�`���~+���7����ު��+����s"�&:|v}#wO��]����������!�s�I\�1]J�b��l���Xw^���pO�F����휈x��ZPv)�;�,����ܒ�B�ݽ� �B�t{'���T��oA3w*��
��X��3	�p�<�$v.	�<�p�`�+���t]3����f%-�#"�|]d���5�e7�&o(=�z���0�h������`[��aҼ�#��{�q�J����㛇ϊO'��!C����u=����2/<�"�^������g<��>�b1�e�b5�5nݽ~�^�+ɦ��;A�C^;������mڳy嚜��1n�w�dS���u
2]��v`�t8'�)f	o�ح��^�6垛��Y�xONVb�a�LnHV�c������x��qt9d��!].�Ԑ��ĳ��2�����&�� �^,F��g��.�<0d���d�+t0��%Nx��2\��h����H %i.�� �̫����vn���Oq\;,u� ᜊ?���4_���0�:�N䑡7=�E�ݱ
U�*��P�`�%�,�Q��]N��RH,᷹Hȩ����6�V^���p̺�<�`���i=�e>��_�o��2���<�о�7�/s�qLXɑr�E�O��^�*�nx�EUX�����L��3]�c`�M�xbq����{�<3��=�L�����oPŇ���O�@U�E��R*B��0M�*�tzp1�]�'�X��u�(�1F�w\�<;u�{�h��Nw���qSrv����b�ա�j�e�(�g�^��owd�or�Òmܴ�r�4���S��:�,�C뛧�������ۢgd�އ<�lW��\f���5!�%=�^yh:9���w�My����}���l�<��
�ԇ�]uC��Kx�|�d�g�����}qhnN��S�֝ԬZ��2���� n��ۅN\������2�=ۜ�T�P�NsF�6���w�VZ1�α���N[ٻ�r<T���O�&Y�����R��;wG@b�4m�X��4FL���.�R��b�}kul�7̈́�ˍ������믽����'��[81������G�7G���������_aҫ����R[i^����z���^�'^�K�M����f;��b�g7���uxUl�n�jc���)�F݇Øᝆ��Ι�^���Nb�uݼw�ʆ���M�w�����.rl��o .���X��(���i�[��4U�/#�E����2��uK	s��RΌf��nlWݼ���!�"<^�odl�:}�W��s�V����yD�Y���<�~~HOj��t�lR��;'7���5�r��Y�T^��˚�/4%�z�&	$�o�'�xL�'*�,���|�p!c�������V��.ܼ�~��w��ӫ��R���C:e-�c*3[yS��̓z�D�)�	(����6�;{qx���<`�혾
�d�A=r�	J�x�-�F����N��Ǵb��=ڳNu�E�9AKb��9t��OU<�6�^5�\9�����ۃQ�K�>o��b��uL� �)TK!;�,��a�f�4�h/�唧�����+^�NMl4��!�ٛG �'5�u;��� �{�]���w���h~���s�yN��f�%�-8
Ҟ=%��+��sA{'�W�4� �����_m�g�U��77ݩ�GOu���R�]�M�8M�w��Q���g�8t��q������PFxU�tC��'�>}��X�em�R�e[v���B�ʔ�|���u�7���Κ�9
����gt�0�����}�9�{�w"8&�s�{nt9Hհ�=�ٻ�3L�6�2IW�_;p�U|��i�(�t,#2A���"��ν��vSBrK��9M�&Zౖ�R��W1��}�GQh��;���V�;q�[QfU����+O��l���tJ�\ ��h����<��&�nuBb�;��}��{QI�԰ߙo��{�y2��!��#��L��Aa�P0�.�f�L%3!jgIO.�ݽƱ�y�z�y3����]bk�j�*Ub��v��"���ӕu��+:4�^�W9R��5���J�7^0����(��{ #���þ�eJ�Zf��AA�H��7�����T�/��wFw׈��� j�j���pٽ�}�f�b'����+^�Q[nIɨ���W��\��|����%�&'��pD7t9�{��tv�km���]�[����Y6�:�I3�K�e�}�k(��FL�vJ �1�"�� �ύ��+�6�M�]�%���/�ۇ�*�ƞ�;�)-9�P������{�s~��gU��w���گwB�����3�>�����|�6�Oy2��hT�:�Ӹ��U��C�j����wu�	�_{|_*x���Z�1j������'� ��\Ċ�b<]U7�[���-^����st�c.m�뙹�N�r�;��J�)��*�ۜ<�/'<���|�Rr����Χ��M��v�Q��z�#w���Gp�o{��:�a�yy�x���kx��H�P�̑�$��ܒ96 �r3��HJ7"�rG�%$��RXS��gP2Ԋ����2L�܎�qz�n\���t�q���s����4Ĺ��o�NnĊ�sf�^���7��m��Q��!'�c�[��8���)�'wQi�i���ԡ4Fpn��n�<q�����G���������:0�i�W�:IB�0ھ����vu^ER�E{v�
M4j;5��
�T��np"ݹ��[�aΔ��ց��c@��)ê�7����{��sn4\��N��b�;������ԭxh i�;��;�(�������I�ŃLC̏ph��.)��-WQ��LV���0���UsG!5���k���T}�
���{�ҳ�z��7Yn	_{�[�܊��Gx�r�Ԇ�_tְ�4Yd�ed.̃�Y������7�AQ�} u����Z,�)�Y6i��n��u�i�7֧tէ�B�Z�4FF����+�Ʀ�e�ns�	G�]_'�.z+��*Z6w:�L`��Q�FYXGb=̡²�p��G����@���i��r�J����
����L*(*����ui  *=Gq�{z�U����D�֭�)�Y���3uAr{�;E�qm�/#�OHcRAYՃ(�H��]��ȋAߏ�ȇ+�=�4�-�u\�̥��C�JFW*tP��X,��^��6��˨�=ȨI��<}�Op�RS#��N�r�}-�͹�҇r*H!1�X���ɚ�V�#��d�0�<+iMtl���P��<�]��FHA�sç����,���]3Σ��.Q�U�{L%@��`Q�j���'����;��m��Ռ�Is���>�$#���Ҟ�Ijջ��}�S�O��W����M7$h7�o�ý�����h���SV	�7�� 0ո;�����]�1�J}� /Tȁ�'��̈́r���x=��Jضod�j�z%���&Mu�����VFN�j�j]q�u��훬$�ᤘ��ݥG� �R��`��xo^��؆��2l%��ԭɰ�L��rN�ܹ[zP�@2�v\��{��Kлe��-С�%��������/Ij<Ѳ��2J�{r?85G������ŻQ��O��#��v�s7@��f��̒��;::�vK��3q[W��9m<�\���c�/��˚OA>fWY\����9�x��7ɳ�����=x*�'+\u��\w(��	;G�2��'�T��=��37�pX��zu�zJ�e�ve�9b���@|�e]n����Y�͘d{�J��0KJ�w/�9IU�)7�;�3Z��QC��E�.����xؓ�F����z�Lx�?\��4+|]�����Tħu��_	���}��܋�p�Y;�'N&)��ڴ��3^*��H2�R��ER�vi�U��!ue��mw��W�Ad�R�9@l�74rµv;�~�7p�L��� D8��pn��e%���yuʠ9э{�92O%3Ƣ���kX)�^�i���}����vj&¹n�WvNW-LH.Ы��S��*������;�%?S����c�Z�5:��=;c�uo�`�����	�S.���J�qw�$#���QG�ձ�Q�f��&�[���;�V+&9����^~��Vm�ьѰ��B���{scҲ�9�"J� #� �^���'��C�h��s���Ӏ���̦a��GF��jL6��Q5�\����(��z�8Nl�'wn�{�17�U�(�q�Iׇ�J.D���!ۇ�	��=�M:��R��wç)�=�J1�F��Μg«.q1��&��d�4��7V�w�yB���9�<��G�xz�m{/��q�� ��~�El��de]q��T�j��%C��1u��f�R��K�F)�p�}��D��Y�CC�}ι_��\w}���(V,܋��M���
��d�	�K,v��3����F�U��`�n�\�SwN66�ɴ��QϜ�.����3v4NX�Hz�3��\��>�=�����o�[�������}�U��+�����j��3a�Q��j�!Un�Dn�9��ګ�
Uˬ�\�	��[�}m4�<Q^��B-����}�0��#@�j�{�����;@�b���yn��%R���k��cŕu=�'�zWe㎏���Փ@CoBL��/ܢzpq7�$�v9� ��_�f�'�&v�ŅC�)�
^�s�$<��Ӥ-,�~o=���rrA���p��%�툽��i�q#o����9�O�3��˾N_��d�On��_FR睇�s��s�%��Z�����p����sx�u�j9�[;��3gPҝ��v��c�B�E��\��v��r�K������DG-P�I��r���3��n�ya�P�ǜ2�S4����HN�z��4���Oq�-P���w������k��*����7�vb�ղe	�c,o�V�+q����}�1��sfeo֌�E0���8�����������%�������7��&�a���;�7 �&��0� ���V4����ǞOs�j��h
�4�ĬP�So˨7Ǳ�e�|�3��-b�|�]��1��"�:g������'�m|��q���1����w�a���e�Ewa��`�K�}���� ���'���fV�;v�s*����n*ʰUu%6W�_�g3�����t��t����7��d����n,Ky�'}0�v��vq�Vi���EWn#���}�;�꾄Ǎ�8��6yC�(��'��>Ŝ-ʈ�t�3��X�@<H�N�6ש��>�;0�E��{��xp�]p?%{�%�*I�^}�-8�*�r�z6�o��E���m���vя�I��uƍg`�U�UX��g��w�Y��p��#6��c�{�ۚ�=�l%�0�{�����=�4N�jâ��C�9ǟ#���yDM�C��w CB�"��yq����@^jw���nG�Xn�ڈ����M�	ސ�b����M=���X81d�ױ%��g�x�=�;���\������Z�f�mN�9�h�ơ���I�NVL:�]En$yZ�pu��1H��Ɔ�k7�����")�Mw/Y/����/.k�^�/���T��K ���!U��J�B����B]�<����#{��̇�{-M�+#��_2c|���B?{5��K.1�auoR��`^�1�3����bʔB���nB�+��i��9ӹ�[>T~:9�Z`��;y�f^��us���]��O,᤿$���a�����7�nxeτ���s�<aܗ��� �a��Ё�^�����wJY��x8��`�Ǥg����v?��M$ ����j��+�C�`�y�0jͰ�~�p[��:N�_K=�L�L����|��w��N�}��&��Eej���<q��&��F;�l�iF_��+J��Ʌ��n8M�uB�mx�5x�L��[@Z�1r&��x�ZNu*�J7�+̣΢����e.yQ�%��d>��^�ڰ�b�D)*�v�}�U����4"f��.m�)�KC�j>q�C�!�l��5q7-�3֐��F۬v��6��<=��`����ͨ����фv����Ca����^�aQ���O��]�u��-8at�Q�: ��A1�3J(t��j�A��"w��L���{��X���{�������V1�w!>{v�/1M�9�Y �I�0����Q]�-��m�D��u�F��郚�;�Z�ݜ��%�������! ��=����K�ݕV-51r�79��j�o���g_]�����s�e!r�y�a�G3eՍuөuC�C�A0
^�oF��y#�v���]W���<� �W���RdQwާ���/ir�*9z�J���O/�N�p�1�1�;�-�q�R+D�Q9v�\�%��P���&y)&�������`<��*߾z8���+n�W��Ǚ�繬����<=J��++jR����fX��s̦-��J��\@č��5�\��"̶1LE-�[k"��Q���(Qq�8R�Xc���-�
�
i�`�+[
ҵMe���Ѷ��-KDb+RѲ��ٍ���Z�(֊�mX�q���f8V�i[ZTQV���9h�����.	F2�����Tj�l����������4P.4�B�O�����1��r9�D�?�_��V}yY�ӻ�k{�&*>ػm�͜G��6�S�`W���^���R�9����k~>�6�����7�����4��8����3^�s[x��-X����9��rsI�M�zn���+1k�n�JFo5��C7�����=:��ѭ�O_+պ�</��p���ї�0a��^��(^�U�y��W=<�~��$�C{[{�aR��M����D�^�4�3��@���|�i6����&s�N(���9/4��6b�m�{�Ow����=;�wI&�{R�t�e�SF�l�^�j�ߊO����c�2�rivAQ1����Uᨋ�n�Y���9����K�kf1�c�����&�5�3�3$x��h�K/'CA)���qX[2�"�$���5k��am��x*�s�y�@۴�=U�$�3���.�}��[�흥/cj�oj��#�~��u��	[���I���E(ؓ^X�����3s�#4o�K�����C�v;�\ɓ3L�@9�V�{�ʟh�@�Ώ(�n�%ɗ�������ɌΔ�� mOn��w�]	�7�O�7_- +�\�x ���j��繼U>�fiw�H�	muF�;o���`�X��f�*�G�&F���*{�����U~=��<�79�=�.��ެ��ǸELܬ�8�N�ې��y�
LJ�)�����̦r���.�����LXy��?5M�yV^�騾���u�[�^���RWD�\N���$����tpK��黽��,����SP�}%��Z*�'{:��dL�$��	=)M����?.t7ڷ �/������-��]�4-���5�{ϫ6V�gxp��1���Ft)ƍ#F֞a�ێ�
�ۣ6��#;3�ӎh��(w���"�
�����V�nuz�{���խ@<����
bP{���7���yg~�|�����v���6)כLa��R�DI��^��ɻ��g�������� >�(�Y}���[X	˦�C�,�a�L�{ݣ��nd[�s�&�el�dW�	��O���d����&w�q\m�;�w��Wؒ�zL�jƃ�{4:3ke�N��SS����y��҈�y]���v;<�x�mm�N��ώ���`��sC��ov������gf��SL�)u��"�;�|AA�%H]�Qَ�༭���fx9������wL����x�}ػ�%���W�����0����t��^�����t�o|����<)�'pl�t�H]�!����.����dd_����q:�u�v��
u�_S�b����Ԕ#���C�=������	�lxw��x�����Oʠ�ۓ3U��m�P*.�`�y�*�1�2Z̗�
��a���d#���3R�l��b�]=����|4ۂ��S�2�Sَ�n.��p=N�´sM��e��a���盘�7C���ҹd˄���ީ��.��$��o�6�)��#z��Q�Y�3Xw.�B�J��;]�UiU�+p�2q�H�@L��[X��렞��}��⚢x��%����cY��`r,���yI8S��T�ټ��M�)W���YN��.�2�{�S5 ��rMm1�e;j��YY�@�<��ǃ��R�)�ճ4x��UWqr�c���Er�˖�vv��G���)�MT�_<���`&�*����c��q�~tl��;���g�N�N#�^e�4Ṣw+Oa?|�	�Y]ZRPV{�y�A_G��e>F��y���ˤ�5{�"8�%^Q���C.��Ğ�f�����kV9�u�<���V�Z�> ����%�z��+;o�T����^Sv����Q5���E�;AEN�K4�t����df��coi�9���'N��y�辦=5�7j |A�\�P��yb~N�/>(�.������R:M�9kM��g�����S�LF�*�'z�K��{f�%њ�Gz�2����:mЖ�윅7�n�S�鼨S��Ի���ܦ�)�W��#yӲF�syb�_��uk�v̼&��Qۊ��u �C��>&u&<x�2]2�s.8I<#�/b ��{�<�s�<�D�ߺ��l�ܭk.̥����iq�aЍ8�9;��*�����M�s������O!&&u�e3�|���.�;ّ�~���ngg!�ڑљ�*&�f�1Y:��Ǚe�J%����Q	Vx��^�M�-�t�n�ڙs��_!�\����6e�ܩ�#"R+�Be�K�ry��_0G/�00x~���u혴$�3��N�hI\dt�@��"�լ���-M��
m@�9��ʦ��Kʇf7N���M��|8n�cI���N5��������q�mǲ�0�5%�7�����q-��=уfi�G��3eV[�G���z�3��9}���ѫe��.����~X�>�cgP�X�G�	A<�e>�K%o�u{ >��4[g�$o
Y�/1Gܽ2���W����q��dX������b���E~>���c�E�DD+&��6����ٮ�+O���}����KŽ��D߮A̱�5�Za@����pv3��|�{0���qE��J����9���a�n!���FW�Eyv_
��E=�8i���/��>���gu�*�ʎA���9���A��*vX+u��| i��Q��K���ٔT�A���eu�y.f�.�u��⡇0֐�v���*��Fh��.�LG:�0�v������&�,�K�eMA�^,�-dEU��wn���t�4u�;"�A���݊v�k�u�}7K;�����*]���<:n-���KtN�Q�&Je������Ke���8��=pQ���V���5���}��*Q��m��x��Wu3GE��g�/���}9�g˕�I��	Ɲ��"���]ퟤޮ.��6����?/u�a�h@�ӒU�X�f�fe�*]�5�� ��ה�+v�����2�תera�rP�%J�dܱ4|����$:��{6�����7R����&]�N�L�ђ�b�3SЪ�-}6)�1Gv�C]���"
��=�S&��i�F�wc�.��Ǵ\�+`{#��M@��5\��jq�ޑ��=VN\w)8x)
Ku��6�3z3�cq�`����%w�pc��>��Y����̇�g�5���]�����~?�u��V�+hX[m���U���4a��"�pfe�f*+��Ɏ$�8�1Q�02��ƕ���PUJث-�.#YEEJ�+A��*����F�J�8�TF8��FT�4��(V�\���ڵ)mm���6�"���&",Uʵ��ֈ(����kimH�F�1���-�D��"����L�V�j"��)QJ�m�A�UX�R媪�-�U�mb����FZZ��p�q�(�[�Dh���s.%����mjT�+U��E�Yh��j�5�;��߇��~���ni��
,pݴ�R�8�.-���U�X���O��麱���1Xr���Q���U����KffnC�f�_v����]��Г�y1�Uy�G�c�0k�Zϙ�$0��qTS����]5z8���ѡBִSԆ�6��m�
.��G��:���c����Ի�g���[>΅����T������J����b�jOd�P��KU}�v�n���ժ[<uM���-��4���\�M�w�uJ��_s������pZF�Y
���	��L�L��՝U�j�z`�$�w�ӌ��jg��5�}�֫���ճJ>��goz��[���4�^��e$�T���<��%8����'�w�g�NF>��""�	$3��ѬD����`����'��n{��Q�ڙ���1���n"���C����,i�]��:~^b�����zn��E٬��&�/�OyQe��/݊�eio;xhX�RӤ�;����o#pf�>��5.]�C�����{�߳+�9<�L�
Z���f^�
�\CW061�
�sI��I6S�!��wݝ��WW��pn:�r{L$��\8]� %!*9$��W;²�d���н������A�<���v_Z�攞�;�����c���+���rYTb����=���Fs�xOsΖ{9^�V�S�J�|Hm��yR6����;��N&ZW��7���>�Eav��]��Oz��-U��٪�KJ���[8����2�γ����� @����f���FF�T�T\{ݮ#����1�p�*��Qnh��\;�LD����,� ̲��㍔��3�+��|�L� ��=�v�\���kvݡ�W�������ۊur 6���f.�63�
|�<��T.R�C��7^�ku���r��{�Op�dޞ�%�״�Uc�W$�W[莭n�r��l������	�h��=���Y!�� �n4�tso��j�*�v<��XC��DΞ��?U��}8B�N\����o�j,��C��ߨ��Z��+��:���*d����N�����?>�!g ���.�|� U�ϴ�W��!»g-���7�\��!�.��mN�¯�}�zwZ}�r��)LT�z{��WaK�<��Y��+��4��U+:�>sD�خ�������M�Ѳ��=��wj{���\c5��t��������s�;��}�2���"��S��~�df[�9T�-,ݿ5���e��6���p�j�U���0�¶�E0�xWӵ�AB^#�s�g1;rr5*���ì;RvX\������~cN��3�e[�Ffu��ǜ{���NF�WF�]�l>8�.���v��9PW�|�4�^t2�yFY�^�l�cެ7�x5���r�E���j���A��^�W.���@tt�(�`+�S�y�ο$pz��Q^�%��oq��x�Ωe��q�(���-a�a����-ͺ��f�<;�ыռ|�L���i�=�����dU>�V?f6n���:���!k^�[����}�6T�w0p��ǒ6��f$�M��J���^Z���-���j�{ϗ��;���`��ޞ�֊[�25�55j\N[s��aCڎݗl�k���h��*W|�v9w��U�h�P��y�X�\v���n���1s�G�3�'��;�Y��ih�����$}��R��`^c��X
�:�����Z��Wƕ�G�]t�22�3[X�tCam)B�(4Q���T�"�RJ��\��r5P�r�/=�C&��]�����u;�I|F�k$������ �.l�������<� � wG��)+7��
�{}�.��Ի��<|�,l�z�(e�w��(Y"e���DM=��p�v�u�`�^��C�v��zy�O2Ȋ��b�r�I�՜Su=x�jl�v��7�V_��f��:n�y�Y;�q}�*C!vU.����NK];����k�Wh$����?�s(q��'�z����{�M*��������O)��;	�Ib;�u�wǌg7����w��vpo,��	C����I��k6����m+WD�:.OV����o�
P�Q��ef��py����50��>��aN�f>L��⺆��3<J����
�Y�/#H*D��oc�E�#rZ��PG����Ѓ�1/���`�E�gi�Πg�C|֋ƃ�,�K��g��@��wE5g�~�!���A~d��߄�׼�n�/v%bM�t��n\�J�m7�@{���/��L:�<�)�C�;q��I��$�������?@�-QxJ�U+<񼳁T���΄�}�_رo�!}�Rߖ�m~��s�^����7+�wx�l�w<{"�cݕt3,�)O���.rr]�BG�djl˘ᔗ5ӱ'x�
�v�nS���L-�q����&����}����9^9C3�A����"���Ίq빚������}��O�_���:e�t2�	�a׉Aao�y�n��+/�G�������f^��h-8�瑃1�!ҠD��(Zt7(I.�(�N�X��cٶ��	bi���˹�wx�8`�u�Y��:Z.�#P��cf4�gj9DQF�\�8a�]X���Kr�]�
�%����B�W�^�eo�՝Xp�P�_�����Ȱ��Ώ��K��ݏG�B����]��'J91��I�W:Eq����I�śf�tc8�o��X�{�^X50�da�����˭��P�d7��ʻ=��%84O"I�Ú�F�J��ʷ��L�P��dX]v�p�;{w�q��}��D��U9���0@���>z�a�!���ӿWO{���~v�+�v����۫�&��P��d����6x�z{7��nĤ���ݗ*)&s^䛃(V�#ol\�en�ᓽ��ٳc+
>�V]�?@��Q ��ǽ�n��v�˜�U��gAk�c��Jx�^��;�}��+��W9�b�6ȼ�L�[f�k>�p���+�	ǲ]"/#/G����=�X��.Օ��1fc_l�#�X��^�ҎZ`.�W�^�\wdch>��V�ty�ݙ�&[��#�-�f��6�#R��J��'"Ifk��Ҷ@"�L���̫冺��E��t�8	]��)f�	�V���ޛC�~������S�L��e��Z2��mA���1J*���mU�`��B�*�ʪ%�1ʭ�hڬc[E��Q�#b1��R�-��E�[FQQJ�"�Ղ!PUJ-�[ZD�J�*#LlZ�Z�KkR�QI�b�m�UDE"���0��m[cjʕ��-�*��X�[h��-l��J��e�C�IY-IR����RTiV�R��-�Kh+lR-D�,keJ�T�R�E��[j���b**���
��*�V*5�3+��++F�V�J%�`��^e_�Yy��>��������=_�ܳ/������Jr�3�	���&���%�7�����z�l5��ui����
������N�a�9y������5��&�V��ں7��E��K�������w�Q���ߩ�\\n7��㍝��Ŝ2prfk��|icu��E�*���x�[om�m^�<6�e�o��*9V	����p��j]�N��v��p���}�p������B���3�>�s����w��]�6�"�
?�/R;��nn���Nz%�+�5��D2����Y�����v3�ġ2Iψ�f)�Ey?d�f+�p�zg�&�͎�0���yd�P�ֺz�BK��xM�i�y�p{��/�/�_�/�6>&�=9�?GO<����clpgjv\1;�o� ^j��E�ռI��ީ����99S�Ӗ!���G��� �.��{,ʡ���Z���LuN�3[ъ�úy�S��Lwu^�d��'��X����s�mxܻF���@�Ήűl�x�Js�+�k5x����tsO/�.q4^��m�2�u묒\��돣ZɎh�d���}3S`��gq��#���Ɵ
Z��ڇ<0�c�$�Ʈya��8n�sp�d9Ksm�c��a��9�7^bt�T3��]ឱ���kb�Yw��s'��G'���59���_7!*�։{1�f�d]�gݑV�F�RҶb^+��wk@�}����pi��G��^�Uc��ɝ.���Fq$BV�Kr��.y]j��88�%�
�ݔ\�x�0�͐��΄ϸ�h>������75#��1tx�]eȬ.1��fH�&ot�L�$V�Eq�8��g���G�� i����$�Qjz�q]�|�q��p*侓9y�:�}�V`�[Or��q�}"z���|�܆H/2w��ySOBy�q1���U/j�%Gc���-��x�bx�bqy������4V	S�_�o��L�e��ސ:?]�c�yN��j�egq�z��܌=c(3����rA��ݞ��1T�jJ���f,� oD�:��}��5
�Q���巖ŝ�ڢԐ�:����)&��S�k1��jD�Gѷ�Y�r,�Þ�b�]P���"r8Ĕw)>�c;�:���96����!h��R��*��w�%���5�o�{�Ҕ��3���Q N�j���*��;��ۂ���������&��}��<�{Y`���k�=~�����5����`Trd���m�[�\ɞ�7���͙^��BM�t}�����臻�GOIw�V���'������D�����v?���$%H<h���X�ϲ��2d�]���v��[7��w'9.��SI6Mr�v��2>�����ԕ=)<'��@�^[.Ј��:ۼ�kGWh�֫i�?9�9*��Ȯ����I��Qs�SY�OWjO\�d�f�wL��=V�B�u�圖l�R��F�|wjc��q�* x=���\Ք~W�=m.�k+Ǵum`�랇o�l"��f*8���2"%����S��̮��#�z��D~Cp�Zr2Ę]�b��\���#[{ǵ��(�-�J�fJaS�2	C��������d�"d��ﾢJ'���t�g���k�|ٛf��Wg�rWl�{��4�M��	ۮ�#s�}��xU÷�V����̺zk�|��Sة�huK�W��z��:O���n{O�R��[T}M�)>�U�:WVv�Vɉ(����m!��U!p�|����ɡ��hbY;���dI�0���c�&r��J�jN4�/*��l��3F�4���.�%F���'ON�Y]����nq�É���..M>v��/-���wb�BP�dw*s�Jڽ;�-ǒu��P�[�{��=ux�4���&8݈g�VȽ�x9�*Om�Ϊ����F�nִ�����8�q�cȇ����<)�5� p帕G�U���<{�Ė�YkÊ�펧O��w�g���< �q#�l��C}'i�����c�9yE5-D�9��̜If�y���C4��:�DE;��qV-���������e.@�s�C�'�/�t.�|ۤQ�h	Y�5{ck��G�Ғ��\�|_�7��TU!K_�A<��S��+7ni^�����B�Xί�ԍk�Ѕ���v;��K7c�����[�ފ�=L����<T��z��wÑ�ɼ�f=�&���o*Q���g��J���0���di��B6]޾�2g����90��3�r*�5䶗y	��iByG���{�&y��|֔|��
��ۊ�d62�#L1T��wD���Ӿ�p2��O{Nkʷ[���Z���ծy�@s׻����Ņ���珻/���H9N�1��B�fRAo��je����}�UUkHW������V��h4�w���ԣ�(/��My��;^b��P*7o���bk3v��/+��1yt�\bp,�՘;�'��ɪmǫ��ԈY&D�x�m�17������a���U6�F�U^�u�$�+֪��T�F�L��&��
ry*4��c(���$�>S�+W6���ו3w{K�e�l���g,w�my"����S)����wuX����&�s���֪�Q��S����xgd��3т��en-�T���m�on����;nF*�7�Ч)87eX��#�yvz[E�ݦF˄�՜��t���l��a9�Z���t������#�H�gx)�dK��|T�>��q�(ٞ���;��IHff�R�7#��,��O���Y{i���- �݋k������x�-�kZ���N��]_�ajnb��3f�C2v��b�,��wFQ"T��B^���OkU��}����8H�$���e���A��?�)R�3��_IM1�*��u}����0��4��W�D�*{&N���oumfD�7�o��=�CX�g��q��Be�\Âl��k��t�&��Б��97�<��,�S�En���>�0��	�sl�#'QBs��tp��{2��U��/��louސ�cO��I����2��¾�n��ܘ�һ^˔���JY�K&��E��}z٫��"T��I�^�C��w=�x�������A;�g��^�+oX��k!�"�%�"2gvᬏ�0��ql^[���M��[�_7Dl�X��Du�8�y�KI=��ݹI��H�V���+%l���í�c�x=�͂$��N<�^�3���#Y
��U�
�΃P�ʺ��͙��%����D�ER���0EL��m�j���R��AT+Ym)m�j���h��J���Je�b�[ĕYZ�S.Q�kj��S(V��-�mF��k`��ci*�Ljb�[i\l\���Lp���+�®Z��@��Y-�J·)�֕T�j���j�WKF)J�(�V��(e� �%(��T�Z��[@��j�VYV�JR�\V�ԃ�*8U�32
()X?�}�~��������f��=�p��`'S�Ȇ�`tB5�'�_}U_g ����}�6���%��&�~Ms4�WR�cW�D�<�4xPEmux�*�V��F%8��Y���
��7[����d�[�8K�ח.�$ԭ�W��9�|��˼�ǳrc���$m��*؅�呮 �������}��eE�O�:%�\��"�FZ<�v�L��n���y�_����:��u���x��bǍ��]K�i��r�)��Nᔌ�*��=.WJ��rX�γ��t�}�u�tG�#s��W�U�r@��,���/��O)
Ӱw�um�>2��'��:�t){�A�q�u]���`��{�RE �l��}��盢w�w�L�٥O��T�(S�1݉p�"v�;1�ڐ=��W��T��Y|pDs��	�ʶ�VϞB��S�'��ѫ�zꜚ���p9˶�0����w:鬸qcryBB�L2����Z%�9�SH����5�j��6J�9���t�Ӏ�b�eO�l�7i�i����dNu�P�	������S��t��åM�Ui��Y������{޻�M���Q��ݵ8yF��4N&].���1��̘���Q����={�ע�ʣ�E��Ϣ{�xΐ�a��J�=�Y�8�P؛n�8ۣ�n�Z��x"2�z�8ܞT��H��\�,�P�S�����X-�@�k�����J�k�� ����u
���u���)��Yo=v|�՚��GqND�U9��Yg�q���Nz��|c�|w�:����J�"���dt�kJ��Vgue8VYp���r�_�S�Ɵ%Gg,��A<S����>1����W�W���Qg����Bk8������t�.]��'����z>��8��ϖ/��}=@eE�v�+���r߄�x&��3X4�>��%��e:���.Β�ח{Eܾ�>>t��;�3]���0&�5�!�&�*���~`s(C���!�d�a�@�!�OXk�O��}o7��_�i�� ��c �M!�$�[$/��`z��$�������V�~9���}�﷯���*@�q��'�R�֋$�!��Cl�2C;� z�z�:�~I>dS}w~����ߟ�
�������!��'̆���1�d��HIMX���$��߇����=��E���'�9a�9g�ԁ�U!�2k��� � (������}w�~�>���PF+�1s�6M:'B�fR[�;��gCp�˃��>��/i����7������ +o��!����9a:����8�2C�����'��ܤY''|߷}�3{��y��v`|���M�N�o�d�=�u �P����o��T���@�$�������w�����c
��2 3��ȥ�J%�c�N$=a>`}�CL�S���<{o;���Vq�g� VHi��!RdRV��2|�y�!��N 9g��x��:��������soB;��4�����ЛI�a��S�!]�u�� ���v�q��i �g����~��������m���RL��$?2`i�$$��=OP��%���<d�~k��w[�vH~򇌓������u��Hq���'z��)�Eb~a�C�?w�9I6���z�r��!�l����q��z�
sV�=Cԁ�hM�(m���L/��y������0�x�H|��$=�2��a+�I���Y=@4��gy��3y�}P8�w� x��'c=B��HO�?2�7�=Bl'�r�N���������/��_xݷ��$����Z�ވc��B��U4�2%	�5q)��q���[�^4 ��x����}_UW۠�z��Y�:��1	�ClXI'�+$��I(�6��
e���9��������~aąB����Y?v�x��N�WԜf&�*A�@�}���Y4ʞ Vi�
Os}��w�����O��
�k������8¥M}I�N2��y�H,�0�6v������S�4�LĂ��Zx�XjS���������Ĭ>aR
T��M2~eH>�8�H,�E���B��N&'���V��H(~>����?!R��u�߾��~�? VLeH(u%H<�fS�R
CfR
g��8��YXq�`|��L`V�q+��H,�&&�*Ns;{����6��L�2�;��A`m� �,�~@����=�t�R
>�����+'���
���g�B��y������d��Z��� �|���Sh��E��RT*AI���0� ��
���L������&�"��>q��������כH,�%O�4�S�>M�I��T�`cR��� ��11�l������댋x�R
Ow�;ߵ��}��z~�&�+'��I� ����4����ɿ��AO4wY'YR
q�Xx��$O�H)=d��J����{ַ��i�Ƥ��`q�>�H)��N���
���=f�:ʓ�AH,�q ���1dS��&2q�<@�!�&;�i}����}��{���<}#��A���OFxN}���;���A��g+/x'+Uh��\�� �᦮��&k{{���w�>}�`�
A~`V�>@��>|>�� �,5�ݓ�R
N!Xj|�����*AV
�P�a�
��w���7ǁĂ��*d�*ĕ �8Î2u� �l�kXAOP*h��Y�Aa��a��@ח��
K���6�~5��{�v�8��*N�'��;q�Ʋ,R
AI�4�Y<��I�+MH,8��M~�bAa���i �y��2|ʐy��}�w_~��q �$�� ���ú�}LN�q�Jʬ����i�Ă�P>J��]H��c'P���K�����������.$,�{�`d�ʟ���Y4ʜdZ�}��l
����@���8�$�$��RkϿ}�}�����`~j|��C?2�:Ԙ�H/��ì*�&$M}f�H������T�� T=a�~aR<a�Ă� ^s���w���<aY����>@��~ё�������~�L�~��}ҍ^�q;�h\Ǚl��o*#I�.�:O�V���;�xMQ����G�0i���1ݕ�Uf�-�w�^��]�k��v�n�{�
���r���(��h���׽e��M�}י���N���:(�����J�q�i�w2d�I��ی��������5��?&�������S�]�����0�n{�ƪ�16x��C<v�F�Q�P"���DJ'0i#�w�gՐ�d^��a����9�� q�	����l��.B3ohS�F���$��9����z{�����b�r�#=y!}��_VMZ�'��oҥ{v�����t�x��Ȅl�@�{t)P�Q��=�(�VE�!�m�!���陌ⶩ��i���/c�1�(DgB��\	|7����У�Y�7�>�JI����ɯ�8o?{݌�Xc+3����q��y�g�?/�����܃Na��q�KA���x��s�[}��b��T�֚T��:�K��:.q�Kg\)��_U}������������*�H����qvd���\j�nGl#I��>� �p0�<y(���x�l}N�ߛ��P�;�i���R�V�M]&t������ ��jb�8hl��m$�%F�`Gt���%l{^�
"�(%2��������l��6��'jQdiڈ-@FĚv��>�Џ��'ԠS��G���w;����M���6�iSO�Y�|x�1����o���g_(I�Q��E74x��2�H΁ AeOJ7����;z��cHޅP4�ӆ�"�4��pRLF�Pڜ�-���ML�����uu�״T	Ʃq�+_eZtf+��;GG3 �m��y�r�j{w�N���3{{�=�=뼫�埾���6x�:x�}F�YA@�0}Qnks��'�oۺb[�^�����m1��{���uw��A�KNa��q�#
��עnp�a@�
>���%�F��`v��}�(��F��0eǆ��3�9�5xv��!���?�P�FL�{^��]Oy�㶧�i�o��~�C׌�+�Ob]�d'2<E��e�;]��#�T}�{��f�x���Dcr'Dy��x�
F���y����O�adt�q�ƨ�Q�v	FF���Z'������#7n��p6&޻q�+'}�7���Ɉ�
��	����^���>��r�zc��;�gH��q����:e�}�����߱e̳ ��'���a\�Po�F��9�����s��a 	��;ɇ�4n^�t�s'l40�6�Dl��q�H��tt����iGy1޷=ݎ?N菏��N'�NU�B����W4���8�7wdJS�ͻ���Ѫ�ʷ�3��K� {�r��(A%��$Ԯ.�E��+:��s2���p�Cj�P��$���#H��ok+5�:��L�H�3a�,�fq��.��(e�79�4'6]h��jK�;,f�r]+�UabV�Ž�W��Ej�u6�S�Q��v�c����I���|�^���;��a9$0T���E؁��V�Iq
�б�h;J��OR.�sr�"�(e��.�I���4,���������	p��ܰ\�+A�R��$�^K��n�+&��`Vjƈ�p���7�xJI�Z���pN��������25���T<݋���4�f6b�&n��������`�µN]���sm�o`Ehp9�ݲoch�h���m`�݉Wft��"Rt�+���$�t�$���1��D�!T$JSp������+c��Jm�7����s�֯Y�Fɽ��u��T �n﹥�+���>�F�",~>ϼ0���ŋ<L���Ȣ�V)m�R�+F-eb�Vըbc��B�����Y�c�e�)�F���QY��S�V
����(`��2+2�̗2�Q��b���ZUb��F��+nd�`W��2bT�[����a��
���"L��Yre�(�*VV6¸�J[D��J�m[nd�.1b��VLj��YL*��S�
�\,���5"���Z�%q�@�J�O��o�8s،�(ǳ��ŋF�j�r\op1tK7��Ͽy�}�V~�_}���=���ˈÖ��|%�-"\k�e;�#a�#bOv&p�E�����nԲ$�����\q�S!�n�W�w8�x1��E���Iۆ@��k�V�.]�+�v~��`�!��������,�B#�.A�s1��*��(�Ǐ�G�NA����B�R����·�3F>��G�!8;![;�p��C�@s[BF�5�HF���̄lث{]}ځP: ��S�e8�g�fȃ�rXǫ^���#�%!lANXVz몯�V�ŽMS�wfݭ`z���~�I��26Up~�oq'�̝cM=��n9I�Aq�9N��������|x�sy�'>�����@�J�ٟm���d᭍3�i�^OwIYR�4[��U	��᪏F�G��v��Zo�%�#����p�(��pҺ�t`�i��$���G;b��̇ʜ�-ƻc`�q��	�� Õp4�@�},՗��̼M�,��FB,�ܣA��G�@�}\}���oG�n�r�?Ja8��Nh�x�ݏq�9)����=9�0Q��h2B������܎7�(����T-kMe�0|�X@0����c�:��>���~ӊ #w܌2Q��٢!g���fT#U���Cw�k7�*ݪ�v��P��
�[a�N@������b�c�%w6)�u������ﰰ�R�ּGH�cTa�4�F���FE⚖�qDa��64�}SU)DK�$.�Jٷ6��`3㐊>��LI��9AϢ���0�Е�}����#���EGN� ^�U!8��-��"}���3e�L��
�pЈyC<o&�[��;��ĥ��g~<5a��ӄh��4[����w���SC���>�wˮP�}�t��8A0�orф���M�e���]X;;�Cp�/?f�������D8yl��=A�РE��d�v�&�,G~ӎ�Ow�)��p��g��N8s̯���t���������y_{S�i��� ��de>����L�
����oAoF#� ��c��裟����kZ߽��~���'�Γ�0��<���S���_�oPXB��b�:� 9�p�e���h�V��<Q���;4���M�u�S�����߹�o�9_���<Y�{|�e�6BPLb���k����I��se�<E4}f�NE5�q�q@�;������Qf��]�4Q`Q����y�Y<�>�s�4p���M�蒈�6�p]O<D��Ȟs�D��G���4�F�H�2�4��#'d3�qD�2C�>�dipɢt��yz0i�aJ(�	�p�M�C�8��}���{���/� ��`�tF� ���8�f�;�����u,Ч[T]�p���6�gDV髉�Φy�1G?W�W�\���me�xG�F�=(�L��@��8����w�X"o������G�g�����~�9~~_i�T`��U������>�U7�	�g�ݧ��{���>��g;�?�'�c7n߳�+�,��웺7�~�n�v��/*�@�t�f8��tȷw�S��x3s7����>������-~_�_v���q���@،#v��8(;O����l�Ʈ<�t�܎(��ϙ���ۻE&��h!�0Y�C��B5{"TY����X��U�C�5��Ӈ���<y���كk<k�Y!%����e�W'V���&�^3�{ս��f6,��/D�.�oi�{+ds%!�Tb9�'����yp_����׮�m���N];|g���~��VT��x'��Doz���:9A4E��i��2C|�_of[-��R& 9(���3%�5�,���goO��q�8
4`��eL.d�D�Q��Q�Z����6Ӻ�45̋3Gso^;��,|�\w:��1E(F��"-����9��)��j���g��=�B5e)�xh�(��8`�a�\d�K�� I�J�%Ǵ"�Qҍ�0z��K�ur>����/Y�(���q��Om�w����:��Sx񀡙��:knQdi���T����d��:.���t�V���LKSai5�y:}���,���
gp�{.���%zs����S����F�f�L������ ֬�O����q�̉�,׹HGL�M���-���ZA�Ô����4NS�z��a��9���9��N�F�6t��>�M(�qҾ8k�q�Ƭ�b�F��9�}��F���#eA�4�1w#9Y����iڂC"�Y���u��������3�u�=f�.�}�����n�{��=z�H�5�#�C�QG�I�g0t����'1è��9(�@���xd.c��̙�T�[�9�McGB,����:p��ȐY���q�:.xr�0���(��)%����ˁ�g�����^�7���pk�q������7~K ��j���kV�n�(�TPH��}|\���ru��ӌk09?}�}O5�/��#�������.�C��"e���s���XpN��%�\ސL'�%C��T�G���ثr':Dl �[$���=��dBcn�q�L��1�p�3�y��;�k��r�[��XEȐx�<�:}Yq>�]"���֟F�|���OZ��w�g�k�c��O�]���G�"''3������lў�8FT]@��F@�}��ˤ��2x�;+�;ي�����50_��<|�i&��г�T2��h�3��>0��в`���2�L��'B�W��\3�7�D���<s\e\��VNfL	��M`S�T�m�ϝ�Q��l���ק�0�i�ɒ:�B�7����Θ����%Zl�L��gշ>�@�U_W��޵Wv��|���/��)�,�c㲲��4��+�:�"�?D
U���:cI2h�fϸ�GH,WY��w��|��,񩀧�D��N(�:�VD־�>��ӑ*d`<C:K�* 3�M�q#����W�G�>��&2����"tG��ǌ�lf�8����j4��a@Qn}����p1�m����i�_���a�v��lK�9�sޡ��Dc���O� �U�xmÀc�ͩԵW&YyAЈF�Q���t�Ag㐝��է*�'�u�޹M��<7p�����o�+u�2o���ZRd�R��#��w��6�;�^�d�`"�#s�W�8���s�u��}�������ù�z��Zy�o�מ�z1��I��(�G�ĕq�
Q����zw��f�=���(�N��#B�B6vq�N[�����dp�Sf����C��z�da�� �hOi��/��t�����0�B>ɬ�>Q�^N��c���P��7}[BuH��PO��F.%�I�O�(�x�H�H�Ety3�d8�n!�}5�*����#�L���`ٳXX�<G9eHs���cnx/#�?��A����,y����=����S��y���gr!�mی������D�	����̧�����$���B��wn�vnۑ�a���xq��Vc�~�q{̑��v��Cד�gH#W]�:}��1�6｛<���>�ɂ���T>����:�w��tq�5l�WM�.���:a�V�w7���cƾ��������3z�s�tŶ� ��,�O:n^w1HH�mwE��kc���:=�+0)���ځg6�����)���<M�4���f7�}�p]����pшU�K"���� G�����Yݞ�����\5^�:&i�r��.���:��II�ۣ5.�ž}51Rw۾��蹵�SՉ����v�����F�j#ݕ�[j�5঺@��9���A�z�n���j]������1�~g@!��9�^��ʵw�4��lN�!�u���:A��g��T�k틹D2�'�6k��b@�C�����Z2��;�w�l=���r��l��SH�����R�'��*�]}�h
�^��ɾ�П*z�t�i����
!�f7q�j�.Qcf�[��9e�Lu�k��i6��_l�Pvotwqv�
����Q�à��+�:ښ�9�7��μ|����3�X�&=�8VH�ە�)1�FD���"t �%p��vk���}����t����"�)���=]7K��"�_Q-��-��e���-�Zb��ơL�1*W�L��˗0����ȷ(bT����`�D������r̹�+ir�m
�+�Җ���c1&32�FV�,U�q(8�ۙEX[
�T2֥\�(�V���ሺӅ�E.��ZUa�+B��M3uL��f�²���u*e�I�1(�,SMQ��V
��2ЩJPP�]9�Ú~����'H ��J�z_t��Z�\u)wS�֭b[ߟ��$[4r�:C<x؅"~�:�s�n�Ol.��ߏ������ÊO�����Gh4C2Q�	X�vd�[tY������ $6A��\8s���S�I���E�����(����(c��;ň���?����B���쁅裴���͞��Di �kc����_m
q�l��}����I�t�da���l������g��9ۊ�g���r����w��V3�y��-����P��)F�N��dm62��W�+����O�P��H∵��Z�D� \u�'{D�Uk}�^gvwB�Xf��]����p4�LT�աM����6�0nac0���R,�e �s��}Ik'�(]{�g�V�����p�����z�Y�	�~Ȳ���O�R��ٵu��7G2��<R�8tӜt_���С�N����>�x������Z1]S.���P��a���32@���*c�/����[��]�����/ϩ���9����;�i4�h|�)�kT�� �'z�&P�Ycz�$"p|���������vԩ\���a��{��V�+c�au�q0�i��z`�$2�U��	���Dv�9��
y������}�p(fAf �NEѻ����q��`�����P �f��Ye�۾�~Ɋp��k�Q�=�V��
x�V9άzU�旽�{��]Ů�/���ӷS�$����ef���
�����y�l#��\�ѐ�I�2�Hd]���6��+�G�(�F�k8���jş�l/� �䭋^��\�,���}6Q�ȣ��Z�Y�k�V�~�����x3���(yn�5�	�hA���V����hIޏi�{'��:�`�#
�>���}��\B�������n��^Ӽ���ӷ����C�]>fw|��s�x�S�w��z�<V���t��v�l�g�n�Al�G��8E0�O�O��~�c��G������P��=��fi�S�v�D�i�r"�<l����h����j>��N�N(Y�s��ݓ����$Tm�.���賫R�]�Sg�<��+E����Ў����#v�����I�����/�{�������4���J'-��}e︩�<u�i8S�Y��QE�e���Å�ue���{���⌔�6=�&ٙ����p��z�����=O�ۏ}�D�"̝ۑ��Dp/���k�nN��d,g�W��p̤�?UV5����\����3I���J��)ব��&��镐7�������6}��#HV׷�Tr���h�l������aqA�� G�ާ1��PG�{fܱQ�����#�7���2hdYΓ�U���,�q��:�x�#ggې�}$`_�x�{&\M�ҽ�f�||������3�s�,V��&C�ռ#��M��Z0��A�s�\W\8�wb2O�T%�7�;�����~7�L�{����C"�q��q}xz��� ���9 ś0E<�"��R�J'vV6vӎ�\����U�>�х�9���q�7�K#�@	C7�Q��UR�#6�]6���DQ��M�faO�b�S�8}J=�r�;�=J�h<`�������T��.=���8����70��[u+�����-ϳ����h{N`��S\�D�jym��"|H@���Äg ,鱷(��h�LB���x����(���YVD���r,�S�t�i��ݥ�~9��<e�k�����w����y�3�� �bsfTi���N\=O\|!���~�+{�>冝�'ֻ�*Q��Tԩ��ClJ���eA���U|oZם�gۺM�?��x�k6�Ws����1�R�}�6:���_�$�q��,�Q ւ����z��gn�̲6��dX��F�j3�����CQ�`�6%�ej ��Z�Gqӥ��<��=f'����7z��+��n�����L:7�Ir|H�N�Y�+ .LmG��}��XV�j�Av���05�r}B�t�G��n�~��}v�y��|�})���n���w�ə�ۧ�9��LsR��6�]ו�	��`���ig��m�����zg�_���l�.>�4��ϥB$�tہ��^���Ʌ}��8)���z�O��=��#@s��c���q�b��
���8һ��::Ù'u��il�������B>��3�����z/͉R���)���,9����b��ދ�����1���Βx������$4��{
&�.78Bp�6;dK�2}�Qf��0��ɝu��)�;����'��F\�Qg�p���;k;)�I�Ϸ�}[���b�{Yp���&j��$�ͭ�A�xAEJ�d�v`W�,�y�%�˃wJ���xX��pK���+�E��FΑY�^\d��z��=��E�<D(�>1k`w(�����d�v��p��F϶�YF=>�]ΡE��z��^�����v ���#�Qه��r�@=f�ܱ����9����2�2.�u�!�$���c�i*�auɃd��Sp �8��W�ĚQ�������z������ai�h���/�I��<C�_(����6t���	�^�8&f=N��o��u��I�fA���XX��R���}?�����O�Cp�pJ6|L���mm�q\�K�����8���k�z��_Y��r_��}k���t8�!A:gc����p�4����/f�\p�X7�lag��g�9W��_�"���g>���9���|'㛃=O�~[h������i�#g9SӢX�fNϨ�z��!6c�`M�gRfr��7�=>��<�d0:��/�h�ܞ0þ��ȅDhS��.���y>���Wmt�������v�.v�#�Szdg �"��Im������?}U��q~��=�_�z�'�G��~]>�����Q.*�i�=t�����a�3���<Wo��/��Ҏ�/�cK̐�0ҏa���T��
>���EG=���s��>��>����kg�5H�tr�}'������F��ْ����W������[[\��x�׶{�+���Ƨ��q5��|j�e�6f�v�"�tq��]O��@���;�oj�'�Q�D��ƛ�j`UP�8�8j��wy�o�H{A���}����lY�s�B�Z����;{�q����}�C��_p��:�p�3:X�n)���j�S���ߟ�<r×qZ������η}�AI�a�0�*I��v����`[�u�wǌ�;��~� ��ל�~E:��7e󘷗�����$U�=��q4�,�>q��h���##���G��5AWM4� w9ч��aG��+"E̋�m��f�<��<���OyC��:�n}g��=t9NK;P��B��ې���FBsg�a��,�e��b��IWٽC�4���!dwa��n,�sn��NOh�+���P?B�?
<(L�辢��ʏ�(�{Nh�\z�����3�xP�h4���;8�tu���>䬔"3�x8|�a�M����3�i��Z���~�q��o޹��]�|~�<�p)�{���]�L<��y�^���^�n�0E^��.��+�,JV}�(����.Y��V�9@��gQ=F�f4yg$�Vwi+����vMY�!��l��3!x��;sU_m�z�^ɛ99�m�F�\M��A+^���8��U��ө:��`$�nqIX�v����d�����}��}�$,��wء���{���}��j�W|�q��p$�.M�=�o87q���Ok�;��E;�ț�����s���ʫ˹#�"��0�IGo뉶"�nOiLrŗ׵�6��ۑ��hT_Ql��(�1�����ǗWgň�6;��Zz���(M�u�U���K�{J�2BE�#�T�oQ���h!�,����FB7�d���Ȥ���\��n`Fb7������[W��D��A��Oi_8��@�\��G��j��z�I���/d�}킬�p-T+�����("�F��AS��Y�"@�����=�U�CwbyU�yu�����*�9�G@����c�3�h��7����U��T�0B؜��q\����u�ӯn�={��p��J��)��ΩY;��3��
�O7T�'V�]&nZV��Е�H9�����Z����'$6S0��
b� ��m�3Aα�8�K�p�)Ifn��Q���5{Հ��������B:-ܸ�[�� #�>Ďd�J�qr�PD��8����j:�dr��Yn�Q��j6��[b��cS-]0��!���R���lb�-*�+j�*"�˫b�1��R����a�X���ER����́Xc+Q`�i�-)YY)s+%HU�Ӊ���Z֭��y���!	����TK0�TN�d�%w&)�_G$Ϫ���H>�ͺ�]!�r����� I��4��D{A�;��q1j���ʞ�{^��g9m�wxg9��LsW׻�F�Q\泔�i}���#AAǴ�A͌���r�YMaQ�h ��,�d�C\��I��qdn����7
ul�ߛE=:^j�5���Y�]O��7�/l=<{`��8��2Lt{2�3�1�J vE��!P�D�j��f{S�|gLQB=�0g�D�q�|!Y�E����܁���C>���0Y���q�odIY�����˻���>v��~<q���%(?�њ���wIӮ���p�vC�Fe�F�pڏ\��QQ�A�o۞�Ǭw��>C��t4�<%eGN�=ݐk;\OLy���nH��D��<`M�����}��}�~�~��3�_����	�1E�.�YG�GM=���&s^��|Ϳ�m�)��S^��ۚ�n���֌m�,�dQ��|�y(��g&���C�%��/�4a㓋DR�;�����p��T�u��݇�
(��"b�m{O�I91D=�!�J���kr�1Ǎ�2O�Lz�0��8E�LB�r��s@g�LQ��+�#���I�(�l�㺬kY������g\�i�����ӽ�^>g�b�Z���r�~�x���]���f�ҧ]��*)M�f�~��Iҍ��FǠr��ٷO��;��*ȸ�:�"�p����y�
}��xZ�c/��Az��;��ҞY���ܭ&]�2Ӝ]��u��fww~���}k1��9��L�خ�@�'�͋#*���R�*��әC�S�i���ʲǜ8ߍ�׽�w޴����o��x�f{L����=w��a�b<E��LG���	ˌ3} K����֒E�>#��#c̣4#�|����(�������3��I� m͑J���=���e�����9�wB�8ҏ}S��QDz+�k.o[�4��1��%H��D�
iW��}I�5[x-�=�(�� i���V���9]"�UKe�f�P�(��YQ�<lق/�t��ꆞ�}�J�7���VCJ���Cv�-u��]���våQ�-�c\I��ϳ])�z�f܎dW�	��Zю~�����%�Y����H�J>>�#�1�3�>ٸ������|{��e��Ӝ�;�kT5�X����kk�_�͡D2!G>r4��p��l�Ɗ#5�ܙj���J7�)�$a��y�Y��y���ם��x>5�q�o��gT�^��3�O(���񷛔�K�|O��f���1���M�M��=�^�M��:�|i��5�<u�|�ə�wE�
(���=��#>�h���"g����-ayې��ƑdI�%�q�<u��_<��\�}�{ֳ�ݳ^S��j�R'"Hf�l
<�Ūƚ=G��Շeuu��TBQW#��	+�����X��od���_dA�/���47��Yۓ5���{�{Z�2=$I��p"���~"N�VEmw���FG'{t�����1�DۮS__S=�׾�Z��o�}��g�c�f��Նyv�3�WG�1�gý�@�g��p-@E���������8��:�+!�Qc�0y/�R��=��NhD�ש�6�i��r��2�{E7���o;~���<՞&e�fn{OG�����/ϟy������\B���V��L��'����p��m���nr'����x�Е �H��!σq�Jݲ�d�����Q��!T�e��Z<��\#�b�WA�N��AXp/?�$u��/�2��94�&�j�n8��.(�/p�6S�8Ƴ$S�W�S��O]�����4�(ldq��/!�&̮٪���n�So��=��x��/�������ǭ���y�E@�Y���E��6}�F}�$�:�|!gt��la�;`Y6D8ځJ�"x���o���+�&��S�������z�My||��|��ϑTQ��Ǡ��(��6j-ƴ�=*��9@g�1�(�G�la\x��$Y�x�3��I�Ϻzx׶�P�JD��@���n$�OǺ#O����	�ʼ�>D�d�s�͐�x��=s����/�fe�|x���[>�s�1ަ��v��1)��4i�@���+
�0���ʺ�:��&1Ϻ#�^���*�V�3�]VӾ�io���I����n1v��e)��?f�x���К���y���\�0���5�6��|�����Y�z�Z5�b���⨠���am������[��Q�O��?<A��}��(�Lq�Z5��У��+��N��>>oToE,y�f>�n�9�Ѯ��P0L�M��QÎ���g�y>������V������U6��Ot�囌s�];N躪�q�8�ԫ�G�r?�Kvt8
�O�~\��F�{��^g�Su���u�y�S�N�Β�g1����\���%�!�?Q>���O���ӈ�%�2ҟ�����C��],e�C�v�%8�%y�U��t8b�S�qƖy��4�c��c]5Yyђz����De�e)����OmϺ:2�"���T�'��Ɲ�-�Y�\��;�=:z�����*�n�?1駫/�3��g*�5�,'��*L�cl�͞�]���#���]q�o���u.<4>LI\��7��,�b�^g�]���7]��>dwȺ'��S���_��طxX��JlQǇݙn[�) )��rjo;�cހ:�P��'Ej
.��w�{��OOg��dX����U,n��i��b�^�moO����P�&k�(=����<P;�,�������J���9�O����i�jn1��d��YB�T�^L�gcX8�?\�{2�F�,l︢��e�[~�L���Q�詧�e�^b�Jlt��\U8y�j3+�v*iDe[���X�N�e��ؘ�7�u0�#Ɩ<�������E�r�ي�D)1�6�O-J�x��KqwaJ󍱇M�ر���I�ń֎�ݪ�M�0������7h�%y��;ng�Y���T��P�r��fF��+����v؍=��¡n�.���;��	b��]J랹��خ�C��=j���E�ۻp��ה.��z*�Kc76Ln�F�Z�3ی���=V+��5q�*��n�:��S7t���1䎾XV�'���|���V�<n8���ߑw^��e�7������׵ȅ\�*L���A��]����7��o�Z��/n�ʏlv�݇�/�N�Y��ݴ������u���!�|��'b��E�#��0��֐E�u�v���R��Y�	���'t�|�6��z]��bRg8{c�Lyf�����.�:[�%�X����5��u��LO{H�w�h��S�@�*2�/k�5���&���"�2m�
��J��K����f��od�H�鳙Q �(��9��3g�d觊�L�Z�u�南)o
z$�}z���mc���1�{͢{Z�ʏ�j�n::䮛���]d���)N�ٺ�� �O.�`�v�I�6�۾o^��D�����W���n+|��0&%}��`�S���R��C��֘��x7��K�4"�l��ö�[�+{B�n����
].]ѢNԡ>�kr�-{�?��{V?u�Z1��$��<�M:Qv��z7�g#M�e-���HJ��;��F�'��!俋q�>W·d��O@j�t�Z�Sɓ6(bK����P��6U�}��a�)F��̎��+w�j>��X��nJ#�P���.n�gdT�M1khlW5�])�EIm'R���V�p�\�J�{�D��*3nK�a\����/B�3NT�"����]Zj��5�o�vdXG�U��m�P���cY�u�$�U��9q��r���+X,*c0��
 �aS%��%��c�.Z��K�J���Eơ������1�LV�2�)Jl��
+��i�X��4��*��[Eb�KjKh"�-(�F(�bUT\e���B��	���RH����J]����O����z�2ʒW;�i�_xI�*0?�ei�q"Et��O�y�����Y�&�M�"��e��v���������Q�;�FˣϢ7'�j�<z�߃8]�e�����{DzU�r�F׳:��;�l�z�3�'7vyׂHI���~t�ϛ��:���Rgd���Ez;ϜN�7I?\����a�#���wQ��V�f�W���V`ܶ��8cy���cyy�xt�[��%�X�b2���&g�ˆ��{u�	����k��Q���I�"�&��G^N��m%O.!���}�o�wLegv��j�����t�e�K��I�s�Pr���ì%än��qǆ��,m�zW=�]�z�!����1]�O���j��oݳ�m����I�𮋳�#�]�ݤ�w���vW���͠�-hځ��a�P�qR݃6!��~"ciy����s���2��>u��/$������N�ei!��]��[?�h$���VTTUWtb��VV�� ����}*��cw�j��Qv���\3����@���ǽSλͺ,��;��Rm����f���<q�k	С�C��ـ�.�����+ݦ�;�U|GcuX.GN�>U��z&��w���\Q���Aڞ���9q�1���.�R��j=u�C��62�3Wu��]�]��Hcy�����p��ؚ�a��>#ϟ�MD{�=�6v�A/ә[��"�<h�M�0�Ԥ-�߶Ԅ��f6�3:�<yooz����v(�-ˇz�V�v�I��}���u�����tP;F��~rz�t���"���좈�z���>Rd�&o����DMCڍ��Ӯ@�b3/V�./
�T��l����ln4 <G�t��U�nxu�:���`�m�N�ڐJ����V�3�}��ɣ����bN��@��P��\�hM-����n7K�>����O�$��z�ʧtpr��Mz�{Sח���ïFF<���y!�%'�������[[���d\�5>��;l�J�գhoۘ&����F�Бϔz��k|K��λ�����xk��W³�p�p�1�76� u�lO\O����j��mT�,��)y�4½\��W��8����S��<s�h�$�=U��6�ƶ�ܶ�)X�=���2�-4���^��:��n�(�p��#m9�i��[�>J����KA��osoD�|(f��$�:�j
���݃�FS(-��޵"
���V�q�Mۮ7�A@ewjN��*�ݜ%J��a��k^H\���SQ'4j�+����R��vqv��v��~g[ ����bz-�֋�6���i���;`�Ճ�7^o�9]>W�+�"cww����X�v���ͮ�[��;9�p�5tf�lY����*cr�mB�c��oysw�K��S��5�)q��zY~�:�U���n���һ����6�k�]Ě��s�����YI�ҵ��)�u�E���>@r�y���	J�%��~g�c����z%*(�^�{�H�{�L<�!2m��E���Ƹ�G��Ф��خ�v���\��I�J�Y���k+�M ��[2\)o���Ψ����;�7�]�O+�����㉼�l�gj'y��m�x�I�q�t]��1�SO�wuH�Ѝ����;t��p4\ʨ�) _�ûv[9<��R�Q����ŧ���-%'�n�
|�J��u�o_os�Ӊ���>�06#���إÙw���ˤ�G|<�8�u-��D)g��a�w:®��V�!�:�u|�g���S�d9���S|��e>�zt�ʙ�3��n,���i��P��SqK���ia��_>=�ob�~�Q��h2�����ȭ�z��|L��w/���3�^tWǋZ�y��aU��m��ͬn ���������{��'�B:���݄�V4JY�5i͎x	�.so2�J����̱7 ���&oy!hs�V�Q�ڡ��ŀ�%%�˒���#y�Y���w��JJ�ی����o�kD�k\�s.�aȆ!�Emo7��^�QQ^U�ۦ�:NO��/U�sc%�����r�)z{S����?4�Mz�#k0��|�ݫ������jyb٥}��d�j�ɨ�b습�r�b��b���S�W8<�כT�aާ��ҵ4�w{�'��aEm��������=��i��2��S)RJM�p�9F.�%]����yMOV�3R�G��zYK>+K�4��V%�����n��nI��il뉸3H�q�l���j�K�f<�i��Ub���N����S�RL��t9�gjvR{��j
���Qӈ����ΐ�G\�r���d.km�7`�*���	N�5C��Ң�IőQ.]�;$]9�5�K�W��[�.��	�ot�����-�ܪܹ�|g�֐����������{�Y���=z��I�B���|�7�e��ɨ�ȡ}@�~\�����,�	˰7+$�xCsb渭��9�&������b�2���`+�H����b���b,��8d�d���(<��Y�Ҝ��{��	^hu-(Yo�۰k^��lCFw=䀐)����M�M֬�sY����2���T���v���t�=:�+,����@�g鵚dU�� ~���J�9�w�y��Ƴ|��ux�Z����h���<r�2�'�n�Z�v*4�	�
${1�3��Ewy��+_]>7�b�v>�3I��<�b,tԼz0�%��oq�3��7q-��W�\;*����ݦvĬ��%酮v�:Oe�%f�mGi�t�v�RՆL߸>ݛ��d�'��rӫ�^�gm
����9��q\ @��x�]@����V���с���
���	=��[�p8��.vΧS�L)?�L޺�+S�(�����[]d�|�*�H�s�ՙ�T�I��J̖�Pt�7���W�,��t�CE#)u��^�[�hE�5p.���!���-���%n�-t��sr<譾����� TML�M|�<�K55���x�p¸�|zW6�8Z�������ey�i�nJ��@2�L�b}�_s�pL����`��p�R�g��j��^�.��6.����ૠ�0��(1�V��3)�q��C�.\q���K�3,��I�P�Je�Qb$P��*fY�
���\��YY��`���m������b�(��,�·)*T�	P�2e�8����㙎A-"�Ӹ�߲��9�~g�>�v-��8� �T�jrs+��bP�$��M��d�t�JwL��+Q=���v��B���ck,ONԼ�sԤ;�MmS؜E�r����	��ʤ�T�Nךݑ7|#.Zd�>׸.':�N(b�%��V����O'Ӧpj�9���|�K�އ����D]����"��c���`U�}'cm���5�"n�_,���Ž�������D-��Ms�ݩY�t�r�2�,�%�MP��;GWV.��"D���sq�|�4N��I�4��"���aخ�"� \]
��s{I���G�㡻��W��-�\ͨ���=��n���AD<r�{օ�\�)�
�U���,§�F��8{�g17R�j��ЍnEr��<���S����C��J���N��֍���hj�zw>0&��̜��#+j|K>�G*Hq{�DΤl�0,��=1T{8K:Y\�����'�!�/]-�w�XQ��/��1�St���1W�M8燵�ƃ��$���\+� ۡ|��k�X<c9�̐q�%v���9iK>k*:�*�:�qN�GK"�G��[����aҩ��n�Y�8�T\��z(*���L��K����`��T=����wh[���7k݄�op��y�v�>~yN^Rt�*9J�yP��{4p~�Ft*�(�~�4=3���f�����'�i8ӽ���T]&Se����l��Me>;GU�l���Ol�Q�l�(�jZ�$ʩ��H��b��~�LSJ�a�����{���h�.@����3J�>����\��q�f9��%6qr]=S�i����_��+�>���'�+�Am xN��I��R���>�L�^��>~��}�+�x�E�Kf�b<]گZ��`�/S�L宬���k�#)��-�&�o��=ˤ���W�V~�6~|�+�W*��!�m���w^�����I�ǵ��M��H_yT�����s�g[U�e:I��sN��B�pө��!��:�!M����"�\f�NԊ�K�<��s�T���u95�AK����9�wLNgq/���2�U`���x��|K�J�c���n���2�i�����v���밣��j�`/}�S|��I�WV̶��U[��n9¶e���d:����Z�p=CݨeC�3=�V�����7��WEmK���B1Z<nC)�S�}t{g���%���nf��g�`�>�vR��t�ٌRg���4)��{�-Q�������kHl�}X�R��ٹ|�"82�^4��o��/�� �z��/�*t�% �6�gBV�����d3"f(��<%��3<�Mw�V��0�X�x�^7ڥ^�ߊ��A���D̾��5d���gL���X�ھ���hoHxܗ��=�F={�5C2:�L7����܅�h���'�3^\¤�ƻ=-�A�����aX��I��������Y���ߍ`�k-����T2Ϡ�|����.:�YO��,E�+ށޯ'{&7���g�x�g1ͫ�3�d���n!W���q�q���|��[y[s �'Y;0c1l�0+���՛2�y%r�)��Jpo%�����X�F�]g��K@׈��'����ެ�K���q�k
'�3�6�vw�#7}2��Oo�%V�1SJѧ����f5JM�1sO	
�]o��w�t.\ᝨ˿X»yl���Y'B�z���h�y�v�����c'qg�ϧ#9�JO�{��]�o��
f!N<�@E�Jw���g�$�m���_�j&�@�����u�i��v�	��7�j�.B��/m��N!��cw��R�����/d�h����玦+���fYw��F�W�NԮ�oe�h�*T{� I�q�T��u���vc�(R�VTub����V��m�9��d;�3��r��»u��-�宴(�v�N�o]ͻi��u1t���630��_s����:����ܡ�RO2bn��K��.�WB�aY,AI��Y�"�^�G�G��9��|��&������Ɣ����d���s��/�F�a q������s9�-d�G ����>xqI��i�5��x�(���:��h>�O�P�$��zu}�C���o;�F������Վ���ߛT�̷Enr�"�ϟO��7��]Z73��FCx�n��p�7�ȫ{��n&�f�u��o�j�w����w�f�������#kwlmBF@d�UkH�])���se��;�_(8�R��۽l��Α��8���+�W��	���B�2Ķe��<��k_��'x��o�{���G�&^��}}�n�7�'q-�Vrd����dG50B5�%%��%ۃ�Pax�!�ϣx�������t��.�y��{��tac���x��i�PWa79�����f�^
��^��ی������g����U*��YZA�Nauޙ�x#;`Ȯ�`5��<�؂�w	i�Ѝ�<�=ܝ̼٥|K�=�}R��ݵ��0��}N�W&���Cv��o=�S����v���Awh[����A@��tK(��b�>�M�3�q����
��b|�A��=��h����N��^�j<~�L�W�f�p�Xp)��fCqm`δTW/�XnDP�IU�\�9���QwVc�O��>f�cҷ;tu`�г�ɗV֗,I}Vfq��륒gW��]F�J��++�=�/Zߥ��{��~��OX�������s�^ђ\��f|Q��J���p���S��z�_n��t�����QN�؜��tM��Nm=�����fS���ZrS�X�3;z�v�?o��(D{�����!���y��Y-��K:�*�Z6�os�ny�`��:\�[
��[�S=��CM�u3-2��oj���v��}��j]F��gmVM�3u�����N�4�A�eoK6xa�#H{ �x��O�� {Nl�&�b+��a�˖�kX�A��uEb�����n���Բ�c��Wm��9̪r��b7��7��j�z��c���|ӑ��;_s��F���I�M#Nu<��凶�!YE՝����'���Q������tY�{�{!VN�k,�1�3-�W��@5M<����cjr(�0	O��wpN7�)QJ�@'	+gl�!{�_t��99�:�6.�7��O:�}	���[�wst��pI��B���J�yf0̵�-��1�B��e��eʵ+���b�&[�1\T��Ĩ�q�\�XZ�C��VTs+lh\�VJԂ0KKR��"�AEĖ�J0Z��T��+A"���)Fb��1�2�\J�C-TE�UDb�jV�T��̠�J4iim*J� �XTEm(�UE�Tc)J�����1�X,^��]��w����krH37z�'E�u���\3���{@��>���]~]M��4=<[�q�ѕ:�n��d
��ot������jyG�mMܑzYj�5r%�(�������z%��y��a�= ״��4�.��N���V�Ak��������WCP��������L����j)tH�ӓy�)NC��l��4s����x(�kR�� g�e��}a�]�0�=V�r6*i=�bz*W8pP�6�zj7x�9�<r���%�=����W;|y���:�GR�u7@�4�i��!�(�[���������ư�,Gov��TZsT��|�asZ���� �s!Ѷ��f�nrm�B��+`!��{+���Y�v�!�V<X�����j�f[�;UȆ9Ƕ�|qT���oVؽ��5�_^�eI����4�fƥ�as�ot���aї��N���e)��}ݭ���xx���m���A�9�bg�,�+c;Zv�E����W��Q�]&[jlR��Y����?�LO&���Y��6��.�r�e#�����걔����i��5�{lin�xJ����u,�c>Y��K�r��y�j�qY����l[ͻ�X��ό�P��9NŌr{9��4z�Ә�	���\52�*:��dP���l<��7������7��Wd�p��{�TcX!�%5��O=�Uy�+6��K՝^AGum?��t<�]�{E_�X	��xgebCZ�����2.%깣�0nZD�vq��	��dX�=��J9��(-m_i�ܻ�P0�ݛ|�݃#p=�e?�{؟P�P��S���䯩��Y�c�����A`Λ�Q��{����Z�����9J�D[<�c���{)�y=���	#�y�9�d9R��BЇj�S�.�=�\M���ή|�#5�s�7��W�.�/)�U��)�h'�=U8���D˲����<ȀH�ޚh
���\�~�g���H�k��ǘ��ç�=���c�b��6������ڗ��+LH�KǢ���Y�3)n�t�o�.��V��
uKC�]��s F��/[ db<@E%�%�o/��F��ت츃�q$��{ݴsӶ���Wye�D�eF��$����~܅oI�����R:L�v���n�~��4��
#���%�	�����J'g�f�%T�K\uGZ�s�J�� =�4�ιSQR���U���t�z ܀O.�TƯ/� �/In����e�.��x�>u�ʶ9eլ��
)��q�7ѩu��:&~�%O^3���hG��Yy^���������%9\hvt��Qn��2�#���S=��5��*$�'*
���8+{�M\ˋ�׳��#>ͫ����{Y�x� ������K�^�J��쓶a�7��`��Oc�Ɠ{���y���<�غ��{�Y��y�6�Ϫ��o�K��N2�+;�E^�Qьn����{/_�Yx3�!�����YOI�	o<�n�^8��ig8���P��qԸ]�T�|�p�ažY�V�÷]D��9($E����ԝ��W�I�(}u,'i���*W5z�q�������n2�F�;��^�xe-{�TE�̭�<=�J!��y��Ɯ����ӷ��=)��t��[wp;e[��e�j�>�hmHC+kw�����}ӈ>Zw���t�Q��}w8 �.�q����v��U����J��:eE�i�+�#:���z1]���{��C; ëz+�ܵ�l�þZ������<����W37l5�9a[���w-?w�����'���=�[[�u:�ǝ]g*�������4�#�
0kF㧜Ͱ&I3��KgP��D���=ȸ�K(>CC��T��ŗ���ߏ�Zm���}$еe��<�z�jڜ���y�8�'���F��v�A��{s�
���>ĭ��T�"ν�M7Q����Vf)�[:{�L@;Y;$��z�]+g9��f�!1z�����<oEsbof_S0Ҳx�}��c w��!����l&���mD����IyK�yא̉��I�鈬[�N!��.��s�@�_R��C�6�j�a��2s��Y3H�.�<�����1&R�o�g�Ĳ��K+Ɔi�.�ݽ�w�<�Ħ�	�y��Չ��o��K��؉ۋ�z�SN�$T6�-'o{��ӗF+��.�Lr�����9�'�3�g�$�3��d��"����pl���H�ݻ��8����2�>���ɋ�9칈�Qzot�E��/�'ӡl���o�B	t7Z�����G�	�>\DJ��[�U�]�D	t�[�F�3�����~�k��]>���PR�3G7R���5y�\A�.�5� F�f���p����K�b薖c��L�٩o��N��dV��^a�ʜ�R���u�j�#:��
��+���Pws��4i��Ә_���g}�g,��4"�hd�V6���.2E6��g<X��9:�E��Nj���76Z.��M���O{�<��1g���n�t;٭g#���{�>ߪa���̪-MIZ�+Ų��S��Xl�&	Y��3o$A�UX�O��;C˰��t�	��H���G��e�G6�<�������fae��9)��������f����������h	!(�������]P�](-B���!���H 
�y�_	�l��WJ���i��y>sKk��(o���9�{���w���ѿ�/���!d|03ȫ}on�@�r�����ŏh�Ԃ��
����X��������|���K�lp�ԓ媘4S�W��1��� 
�`=s������4��B�R�Z{-�#Q�G�&��g����륐��7 <6�0�.�G���s J�*�/� �k@]�'eǪ� �>��@	!0?�BG�P�l����_Y.go�K�qT�0��fw" ��l��'yn����qv��{ѹ'l��qJ��d��f˕��zއ޲z��}"�ߴ���2��^�\��.��M-��ǘk�P�t��5�l��d	oG��=8s-���"*�V�~O'^�5!з/ɼ�sQ�� !�7�z!�����`�A�$�w^0C�W@�G�G��?�0c�Bs�ewPn������q0*)�U�,iE����!��hЍ��0"�TajHԼ�w��Q���d�jLL�zb�
����i	2��V��P$>*8���a݊��x 
�]�9!�aH��k|'���?�f[M@|L���u�Ѡ�>[�U����AB6�Wџ'�8��O�bS�Qx]��	Q�:;k��Ab<d�}���#�FWΡn�0hi�c�3���d��S�w~Cj��6(�x���AE�q�z@��y�g�V��ć������P�� �WN�J� ���o*���H����Ɂu�$�tچOTuIN�
���z���� HAQ�XʞCCh.��{����\u�����$֐�X8p��Z�fW���Ҕ�dЂ!ĕy�����]��BC���