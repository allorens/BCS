BZh91AY&SY�k��_�py����߰����  a4~�� @WD�  �    :=�C��h �9t�{�T �)T*����I�QT�"�$JDQ((* ��U#IB�� �D <                 ��   ��Y�6�Y�8�w�)���7\o
�G-(��kZ�UVO�H���R犸<�7���d3u�P�����nx^�ow�:ttR�pr(�E�w�Q!�   b��%l��(#�]Q ��q!�x�
�^�Ҋ���hһ�v!��]���� 8�l��q�Pv�+m#��h�sį<zv:t�ܚ �N{�J4tl�齞��W��[^�z�v   2. t ��6�ne���������һ�$=tpC� ��l���n��sF�շZ9��*�r)�� �Q x��  '���NF��v���Z
4G�ۏ%�N�����Ҩ���������5��%s��,�ɭ ;�C`  ����vltwuƹ��v�+m��˻u�烻����8 ;��;��{g�வTl�ht��g���+'N��                   (� ��z�JT�42�1� 42��H$�T`� � ��4�!� HB�P	����h0�L  )��M4�EFC&	�	��M4i�# B�*4&MSڙ��=������jhf�����H
��a�R� �҃ڀm FM0���}��Ϻ$Ѳ�j��ܰ��p��?��W��}E@+�1/���"��r�� ?h��1�E@�T3_�������q��k��������S�TP\��������O��� �����ȟ���7ΰ@E�=�����/��3�����&�+�����[1�����f��n�j���{��Wb����
�P��J�p�m���W�g,��T�~�`��B�W
aH����`�Z-�)څ*�A	�X�	F�CB��N�L�ܡSj���H\#U��i]�St�Q�Q}� ���ʦ�S[�W��m�W-�ʡ�n��1J��NV�1F*T��B�!�!;VS��x�;MX�"H�R�O��"�#���(L�"��8�,�:B�U8��lMS���!i�"yǏh�ԢX��lB9�I��B1�V1J��U�v��5�'���#1ǄxB���B=���[)
Jp!aN ��E1	��B�j�����q��cV�3�B�\F���?w�p!IN-Zy��K�V��5�Q�␨��b�#�)�B��B�j�ǟ+D��I�!Y..)�)D���C�
Jp!a�!��h�q�Ƹ<�]N1Z�T���x���B�j�ǟ+�(�㘶���۵nEf6�����q������s�b��z�;T���^�X���"5j�b���Kb!Ҝb9�b��,���كgCDgWw"��\���K�"ܡQ���8�4�#��+�:�O�Bj�S�Bp�B�Ս�!��\\Fse�B96'k�-G6�`�=����<X��x��P{��N��D-Yͣ�B>F�@�l���h�<-��ͬ�!w���{�� ݵp�k[�g��W���[U�3����7!7!5!)Γ�&p��Mᙱ[�]����Q)�DA��_q��=����A���x�F߶�5�#^uD`Dd�#�
a�sL���Y��m=v�7-�zs�x�G��ا�Y�[�	��{B �kp����1����׵���7ͬ΍���ͺ���Ëb�s�sˍ��s	�N=)H�0'��p���v��K�<�`��oU��lVZy(ZRm��g'���&r���l*�4�}j`LL[B}˸OQ�NiO!I��.5:h���<�Қ~
�Oh]�|y=i��o�OE�7�"y=�SNa?
|BvՉ`��h�!��p�DKs*
m
�Sx-5�#��P���ږ�2�Bѷ�kFދ n�B��W�y��o�t��O�o�yRR��HZ��!�~�Λ�j�J��J�,�-�Jӥ
S��#r�2'��������N��&#؄���x\)�аB�RP�#��
��w��r��<.�){P�����o��O��B�bО-�ke
5+�!3(5=F��r15�ӵ*JO¶&!u	�V#B��\�Ai�Ԧ�T�B���8W�S�B��oD�i�,VR~�b�LB�Z.BoS�(�1
!I�P�K��� X��+����1r�B�&)E4ũؘ�qI�	��O�O�ʠLB��	��,9<V�ii�C��J��(�1�Q)��
�r���@��g'�SԏX��1G+P�Z��)<D�+m&+m��:��<�Rc�\��lL@�ڠ���Vrx��B=M3թ�RWpsr��k})D�Sbb���	�	�}�Z��h\[p�
ӴZjS�&����,�WjsoV{y>B��*&.V&�1��5ȷˆ#���R�!�z��*9�	���ֳ؄C�Q��WN�ST�t�5k�t8P�j���.�(��nxr�T�QE��kh[�{U�'JE���B�C���R�b1��^�s��T�ǟ�T+
m5��U,C�H�Q6�]��4�v�Tz����P���3M��1u������!Jp�[16#[Z��@C����g���"W?��<_=Q���S�Q\ޫ���C�!�|�k��+V�2���b�Q��e^���^������Ρ�OP��C���h�؄c����ۥHQD9B���@�+�b\>MH�М"f�k�!�䡐�"b��a�D;M��!�M��b��B��F��,�H�ЫØb�\�!�2+P�b�C�!�1�,P&��*o�"�b��oU�_�#&�\����C�֥�-RL8Bٸb=Z�Hp��B�B�!�>�!e�4�qP��bF6N���:Md���B�.U]B�!�M�I0���!�Ū��	��K��d��*2!��YD1b�ʁTz5����a�n��b1�["�b�!��^�ЛZ޷�r�"N�~1�D&�0��߱!��bV�f�H���	<~v�(N��P���uC�Dj��n�VZlX���.B��6!d��_9G���@��务M8i�'"BZ%��H�ԑ�ZF�e3���ƺ��t��Ʉ)PD?D��#,X�E�PT8B=��7H��Dt8�O(�"���%h]�]���؇˵ڋ�p��kV˛ǯ2z�{<*�ޞ0�a����bo�Y�-���b�\�"�R�oĿ�#�L<釐��t��ʝ^��c=�g����u�	�#Q���~-��㟎w�҄�Bn��!�"���f��Îm.�q{ʆk5��ǰǰ��	�|�B��qF+�[�S娇�~=� �{S�c2!x��B����QTk�(�k�w�T�[�|,P�[�|�3_+�������v�==я�!��d;R��u�����{��8���5a�kol��l�ס���k��S�����b���(sz �j3�`��^���zzθ�a�<Q�;S�����s�;�������z��wH�4�2��h��ΨmZ5�o[��a���X��=��R�b��snSG��c�b����.<#��I�.D1�q��%ĉ�!y�=�␤��-��8�*)�L���T�G�#y�&�	�j<�
�,B5���w�p!IN,<� ���<x�츴*1��@�Y�WC�G�qhRk�8q�W|��<xZ�'��d�������))�����㕫�\8��T츴*1��@�X�G��B�\YÍR���x��s��S�z�v�m��(U*Έ�+��-� ����9�G�a���R*�B��,E�@�n���,V�")lD:S�G<Z���-ħ�KCf���]ܙR5��ȱWdQu=��!Q��p���������)���6�b�x#��j���i�,�q�Qy)F�Ũ�q�V�m±�{���o-��Ks)�"0���FиM�#b \�X??rѴxYͣ�Y��7�u�7��pg]C�G��W�y
��,hZй�i����m8�p~O���7=��t~��������[~����߱���7}���<�J���Ȉ�" ��1�x�f�i苜Da�=Oq�w�c��θQ!\2�WJ�J�3*�u�!e	�VZ�\�+�ae�g=O�k�jݶ*I}�
�*���˟��b<��g�����}r{�}Z,�>�6�b�_f��# �Ϸ]�'�q=�Qi����aHA���bP�HB���}鵷"X!̙�Db}ɫ�k��bX����z1�O���Qn!
o_�����Ze��1HP%�Ύ5ƭ��q#�y�����ԡ/:ĸ9�ml��M�g�p��)��0ɥO�˟z뼴��&��N�(pc9��[�d��wq"3����KOܙu�Z�뢔���w0%.1+�Wkz���BŸ�n��1ռ����}�:�p��(Z���k^�ĭ�k�N��F<7|�k�qk�R�b����%��:�:�8���'���� B!�=33���cw�[:)���X���T�<��8� X������Lc���\ީ��,t���%�8����{6��,P�}!L:\N���Ϟ����[6a
t�!�j?���x銼!�c;������S�
�jԅ�ϑ9�M��7�qj��C�3ǚ�^;�!IJB�մH�T��)�S1�ZS�Yw6���\u�~�-�T��Υ�b�JD!�[�P�����P��|�L[�k�s�Z�(�Sf������%:U��O,zR�8:�\xuZ�jZ�P���<��ioT���<�q����3ӑ�0e윗e�x>��vxc0�U���井=�<y�1�pu�j8��`_M�NK�� ��@�L0u�w���ry�%�T�7�����fM�)o^c�ys3C�y-�1�*�zg=;���8)*y����@�,[r�:����&��B�\N�9��{�7���iq�z��0R[�kRָ�R5�0�F@8dO�-�Jpٲ�<����%�S�b�	B�Sޭn!Lyu�R���9�ZW�W�iu�q�H�T����Q��y>�ȧ��Ʀ1N<�הּ���/���=��J��Jᶩ��D��5�Y�5�����ˍ�q�fN���oR�����ϋ�Xt_x�K��ߦ�Y4�p�ɥ�����<$�f�8@n^'��iC�^ϔ����R�o�(��~�Q�zn��f����hi�饋m�|4�<ioݟ�.}����r������^99����F��D{rf�7�q��e}H�ɗ�y������P�1N�����_9/#�8|i/8p\�~��ű[�3�5��'�DkT�-�[�z]�l�[z�s�ɹ�����5ձO5�|T�)��>h!O���;٥m��e��4��Fi>ruu�6t�K9��3���kw3]�ֱ�}��OӥO�۳��|��ɳ]��+K�ϯ'Hq����6|i=��u|�\)x������q���^������'ՏK�OI���*p�f��A�4���̉9r�5����[{���R��K�6p�ۑ��7�T��xV�]�I�63ƶl��}�L�TK��'&�oܚO��H�3&� ͚^��4�}�,�C}�L�K�8tH���f��d���XC<�|pل4�K�4�Ovg~@1�JT���JP�ʏfL�]:`���T��X1�5�!�b�	rniŋ̞%�pt^#+'�C\o�r�4��J�%F}4��\S�'��1�8�ې�2yf#Z�cơ��q�7��'iB�<������Z�š�Æ~�f6Q�w��Ό��2!� 뎾u结GEM7��.<뮉p���'ޜb^t�ǆp9�{��z�ã&'���P8��[���GX�M��sz�7;lᲜ9�M�ڍ�w}��-�o���^��p���'�y>���)�ˍ�0��� �6����T����S�(��e:2M�������]m���ӝ܇�ӡ���7�|1:ȇ��{�~�[{�VL=��	uqc�zq�xZ����業��f��8��%�%gFRx}��D�%w�k</��ع����y�8ϻ4����ʇ�w��G�p��tJ���|x�7�җ����n͔�H^�nzG���l����cL<{va���1
Z��e�>q�k�^�JWUyμı��8��iIR���lަ�z����e���������΢��=�y�k��.y28�]M�$���,��d7deQ��dg6P���D<����v��WV��$<޵�"Em>�����ף��L˯ u.5�F���8��^OD:<�Kz>��fK�M�q9�,j*5-r�=S�>C����BRl���0g�`��L�{&���p��N^NF2�IR���JIʜ�M�p��T��!J���'2M�ن��<m�x}���<c��c�w�"��!���s�K���!)�b��[�(qj�F�3��@��$<��S��Fk5�=��@�g!��L��rx��n�e��6>�%�c)BY�)��w�޵.+��H�|�rq�Os�O2�ZԾyO%�T�V��d���
p��Xolf�g83ã�S���������%ϣz��pc���:�C�8�!���R��-�f�p��}��
SIt񋭮����"�&N����g4�!�g�8��G���t��ټٱ�J�`zu���w��:�,qk�C|�L��㮬y��jg�<�d�ۦ��P8�n<��ݠ"5Uv}�N��!����Uь�є�	G�y��QH��uN X�nz�����j�7:��u�1�����<9Ͻsv��ͲZ�oZ��N%. @8|��d7��˯�I28w�����
1ܝ<y>۵��w&��r��f͜J�i�ژ�z�`�O����M�{�i3�0���	ӹe�������y�t��l%F]�����W���ǅ3��0ؗD��{\��n~�����;�3'/�3[>90�g��qm����7�./8CZ�M�n뱃�^M8��ҧ{S�cz��'3ޖX��磾�:ys�� �<��᤼1�L0�ɳS�oy�����Q%c�Fw�ڼ8a�p�r��q�ei)��9#(N�{��ÇJlmb��\�J�Zl��{�f-Sɷ����ļ(�f��6S'�s��A�
p�yW�������m��W\��y�饳����Z^�s�%�k�R�
uC��)
[��%,kX֠yS��%���X�$X�W̝��_'�evj;8�u����^c��7����qHy,[�@�s994޻>���r��B�~*s]�<�j1o�oR��۟�|��[�BC�q�V�ݎ��6�ܒ�?��cK��շN�%�c���ޛl�%�Gf�9��e)lcR�]�Q;�T��u^���޸����c�qjoDz}q�ӏo���c��D�T?��&�����?�'8t$~ڜ���D}_��+_XP����h�O�k[�H��ԟ}��v(�s�by�Z����S��B���wLL�;�$� # � �>a<h����Ԕ��\e	Hd%!���|c�,�H6Я7B��~b�Ũ�7!Ԧ�rN�L��2�t�uƓhF0/F�F4j���!�M[����0��w��YnC�v�
2_x�[CV���J\�s!�p!ķ�ӌƑ�1m�4c���$T�mȍC�F�PT5�E
� ����y)�h�j�w�U�*b�L�%DA��R��Un�L۶�$ݸc �W����ut��T�{���%Di�h�E��-�&�&T
hSp4���N46*�c6����&�UIc	%���@N74�Jj��*iYe�㦵Й��dF��&QD�����l�lIˠ�m"�uW� �	6���b-���*��@�z�7n��ڍ&�̺�M̥��n��^i\'W3܇sGR<�z��)%=1&��r���E4d���зP{b����mg ��;�7s">AM�@��T�{(�@�w>��w �ε䃸7:RY��<�A��L����M�x������N-�r��'PqQB��%��w>l��S�E�`mG=�%��P�jS~`���5��X2��Ƞ�x��@\k���Gb��	�eĹ����8�4Ba!�9��[���+��j�=���\�ް*��7�wSԝ��޳,�������a{�UP뾻2�׼
�k��9�?�����'����}�i�H7�Ѧ�������6�Z������[��  0 �  �� p� �$@ 
 ,@ � 4@   �  p�@�4�`    ( �� ( � �P �  � `A 3  H ` �  Ѐ 0	  ��Oɶ�I*�r(�\*@ �����T�	���D(��5
a#FH�@�7p#�C��Y��J̨Q� ���Z��u9�     �   	  � �` � X �H X  X� H ` � @$ 0 p�40	  � 0	 �� � �`  �&v�( B   @       g��k���&������AĪR�@2�B�:�Q�Ad����(d���B	\�LMy/6����J�b��4 @$ 0@  �$ @� 4@   p�	 Ѐ 0	  � �
 ( �`  ��(@�    F� �   �  �΄   0  � �`  ���d(D��� s��i7�	�ih
�(R�P��1�@w� b/LG*c޺�k{�  � 0	  �   � ( �`        � aÐ 4  @� 4@     ��  ( � "  Ѐ�L�   
 , ,�$ 0 �|���,p�����M4�R��)�r(��2D5
Sĉ��)	J)�H�)���.��F�
2 rud��1u�Y�j\�2L�,����
N�ԡ�>�_�?z�(�����W�w�P�0����ɗ��>C�����iO�"��"8���mHDFQ�GQDym|��2�!�ʝii�4��h������#��(�<����ڑ�GȈ��:�$#JDiDeFQ���#H�4�JF")�mGB"f�"n�"��y�ѷ�G�G�i�ii��ʐ�!�1b#�#��m�^y�yz+jB"2���:��#��h��P�>ChB�j)l7����xȥҪ���5yTdQ�ӒF�Q$v
V0���m������7��$v����Q	��R�k�]O껺�9P~z��QG�*p�F�UYbhi�En�
��B0
��մl�j�V�Eh��J�nǫB5FV�-[��Z�5$&���[a�ZU�Z��j�@18�%��0%�Z��˫���B�i@"�����M�*�*keD*�'F��܄v!�B����r��0�J擣��Cu2�1J�dU�)]v�삀(!�K+p�EL��I!Ql�G�T �]W\��q:�BQ۩]n�_�u��YK\*j� �i�HӪt�w,pV�-$I��D�SM�K�RX�(6ETjU+p���+P�-v��K�Z�G�ث.&KQ"�r��X�,��Y��8ꍃ�RU��c�Y�UeVH;�hP!#��(e�dv�]b�SB��µ:�R �� �$m�څڡʢ�c�(�CcV���y�+CQ[Q��%�B�����V�QYm J�rF٦���Ъ+<��9zn�5	�bQ�hՠ'`8؝���VKTBm
V3L
�
�NUt�^:=I�A�,N0nK]�A	����4�H�P*�d�Cn��;Ly�XV�BB���FAWZu�`V�R�>j��Ah�l����"db�U�Ք�2&�\��J�b|�7��J*��c������$Up���T��,n;S�Ym$m��F�[	#�I%�[I[�2)%uK[�r���	�"�W[,z��� G�1���tR��U)d��4JjI̖�AI�Q��RrQ���"�BT:T��[S��ᧂvL����eN�֤R:�*���u�T2ژݤR���#LV*�qƜcr��+��Z� ���B6�a�Q40���B��J�]�J���R⊫+�Gk���m��2�Z�v�!*��5Y�i,m��m�l��J��c�$-����F;Ql��*��m��
��nꊶGE(!Y��S�C������5+���3D�E��F�2V�- B����YWQD�I؞�a�4�LrJU*V����n�Ӊ���5P�n�M��Y]Ա�uK4GBȝe���rG����.��]-��k���A�I��m1��5�;%n�����|�f�,��
�V"Z�-Lx
@��Ie�E�c���M������@�;���) ꐒ�ܥ�rҺ)D낔BdL�
�	Ia$m�c��QT�F�@j�Չ����%ri·�!ښq�%D�U��6WC�8TMGUAdCvH�n�%R4U�ݥ�R	7j��d��分��V��X���HҏV)\g�XVBD�X�@ake���Sv�+EL�՛��c�S@D�����:���ez
�I����K%MV�I"��A*8��G]�68�J�U��P r��鴣l��Z�m��ȚjV���V�0�p����j��SM��T,��QJ)n��e�N��V��n�q�n����L�M�	TU��U�ji�#��(��X��8�6J��J�U��R���TEmR�T&�bn�O�^����*u�ǣU�����#"�Ț�8!��[T��"��lC��V�Ub�@hV�,Ԅv��S2hNQ94ɦ1��PH�)[��c-�7"��H��M��,�4T�(�5ێZ�WX�A���QU\z�j�i��dV*�lm��lq�[&���D�2j�GIb����Z�L'�Ȅ��"��#�E\��*ER��ӎF�hR4�[
�+MW#դl�@d��Q7R�c��Ee�Z�R�RP ����*��k�zhd�8ےXYSL-(V�L���QZ�eH[�b�`�6j��@�pН��A�KI)[�VXӮ����	W���#m6QZ*Ӓ6�C��n���[J�j�i����*���$,!c�-$ht�����UH�N��W	E]��5R6!��GUVQ�q�Kb�EIj��t���n��H�u�-�Y&�nbq��
HJ;cMG+���,�1�Dh�uԛVQVG(����eEh����SV7(�DA��۲�[�i�J�!lVE
Gl��V�J�j�%U���.�

�l���tܣ��U�i��&츖��,Q�GTsR��
�#ei�EԵ�](�q�ӈ�~(��QW\К��pQV�N�`$v��*�a#"t"m9\���KKcu�Yi%`쉒�*�IQ`ډ���_��	�6У�n�`�j�s5�V�"��&� ��Z��m��+]�V���m�hU�Z+4��r�;]�N�*�d�Ժ�q7b�uB��E++��Z�ziƁ�JnL�cp� �P�ӄ54v�a
GE�E��!�X�Er�*�����T�&;b�2ҫl��M�l+#�N(��$v�v���m�jI(�h��i�@�"�T%"n'��M��٦=U$t)���r�ꖦ�I-���bʌ��1����b�b[,l�hUK ��r
V+H:��M�ծ�cc#�Z��*rA6�����[ �6F��h]�l�k�����_s���`  �������/ ��  � UT}�y/{� �  ����似�� �A��I�I��}��`�0/e�K[Kio��q=U<���<�\E����.7锑��	k*"�tj"����W��q�(�t*�u�����$�T5+$PN!���!���@�Q��dj����ޭ��&�ƲPrd,S�؊������$P�i�m��P�mꌶ�`���\��B������CR�,�`h#j�Tcq�,�:�hIlr��Q6�5XF��q�
6��BTb���[�ʞ���GcAk�tj�["h�+n��lT'#����m-D8�jj+jB�ABhi�Eb��Q��e��j��cNiZ[4�TF�����H��ʢmA2�YE+U٨�t�)`؂T*���Ԏ�"��0j6E$V�V�&�-�j]:��u4��n8��	�+U�H5E[V[(��v�&��Q���e�H�jV�M�%�R��:7m�Q69���jF�ꪲ�Z�Xiб���M�ZzQR��`�lB��88�)]��MY]����6�Zݶ15I��QM� M$�T&�UV����O�����K�V�;�lo�8�*�:\�.����sdy��8R�'0�ܹ�G�/d�r���ӭ^d˼���b隊�O|Ʀu\:������y��mz�0��ʿ�+q�E�F!����#1E��E��1�#���^�Y%+o���N��"6�N69��k`���kx��!�ÛX���^�,V]��X������,�F�h�f�����ۗrV��{�v�㬴���0y�hqM�m���lꭍ��8O6�z6��j�y�x�~�hi�8�ӭ#�~"#��h�(��uƕ�UVYֳ��%�i�` .kz��f��mq%�qR�#a�Vkl}�ڎ]���6t)Pk��[�-~�V����ZV`þN�҉�ZE����d�m*��^�M�Ow{��koImqq��1^�|E��Q3�j��e�E�2������$Z,f�aF�8qDG��q�#�)�on������$Ĵo&� ��Ʈ�	2�V^T���{�bf�o͑lz��Z8�T�<RT�-:;��x�G5��+ˆ��6*�6i��o��rL��kZ�X�Q��$p&(��1iE�D9�tkze*ё4p�^��xb�� 4�V�iU��^׷�J�&�n?31��'��8H9V�t՜����k�g�a��-��i�μ�"#��8���+�񮵚S!��!,�� [^]����]E�qp8�����6:��n�٬�%��4��fLlN.#����a���
(�oe#E�f��6�1r��J�O��`���b7ޜ���ܔ�]��,��ԕ����Z�<*G�������H��u��0�a�i�u��m�ݦ�( �,�
6[�-�DyGR<�q�����"��o{�oy�WV=`�c{�һ:��a0 Ի��=���72s����=՛Rt��Z����#�������Uj���\glu+����k.#��2;Q{Ь2��N�β�n�)�Uw�����)��]Udw7
���4Ү�);Ε�˒�����P����T:��w/;-U���B�K���Y%U��:�-#���iZ�!7r�ךL��;�Q	=>��b9��M��.7�h�h�-�R]7�����-IN�M��,�#el�A�,X3�kh�z7�d8���&rɁ�T��42�h����nju���FΘ"Ifr h��e�3���p��*k8x�jGZu��uh�"<�#��yN������S��f�
<�5� 4���&DR6l���UEa�R1tj׸�v��x�H�yu?�!�C�KH�<.[m��/<��ދ�4�gx����kn��}8���R����ǓkoaQkX�~�06�Ȧ1��4w~����G\7K���4�壍����X{�wZ��N��F��#���<�:�y�:�J�PʱT���N�uQ�Ҷ���sW  ���Zt������ٵq0N z����#]i�K�˶� B�Q{�v�&!�\�Ԙ�\}�e�*�|��nm��/1�n�]S76�����kz-�x�/m{���m���G�ߣ�^9���7����f�8�*T�����>V����ׅyKm��u��yuH��uƝ��{u`�ف �m��[�\2&\�zUQ��@o���<��넳�Ww������#d˓>������j7�snM��P�x��p���/b��9"�8�E�Z�m�����h�kc�T�B6�/2�FF��z��*��/o�F�.���Ѳ.�Q�A���h��n�Y�@�x��p���DyG]#�)�M}Nk)FS�M�[-�-I�an6ѷ��.G��a0����
�R� �u���7�n2oV5n��:ʲ��kf�f���e�]�ި�̭��8N͐��U4�&TT�R�6���w\�YY\���ɽ�����.`�ܧN��.�{�Wi��T�ը�0t{�7���m>آVc�Tڅz�.:��4���O�?���j��[�*��kGCG�ȇ��b����6۠��QBcm��ي���{�:��A�)��.�f�P� @.�9��b�ܛ�m��!�7����Q��m5�k�i=5KC&���-Z7�a�Z"����{��7X:�����f]Hq�������v���=���4�,6�wc���QO)��F��"#��:�yN��Gz�g-)��>�9m��-kK7���8��Eu���|��8[n[sYp��s]�u�4�m���F+Fэ��2(PN�׈6<k���,-�d�)�F�����:�*d�f6�&'\d�U��6���4�VI�h�4il{F���5��S�"fW,���2��3c8a�`�3Cñ�e歛i�U�k�t��V��r�Z�f�ͪ�fך�\[6�/5KTU�ΐ��ޏCX:o�g�L�����h�ȏB>�1�a|"<2�|Y�|3��<|Q���n�E~R?2�uO)�Z2��8�ej��ej���f��l�y][meV�U�ͭ�q���j�E[��^e�R�e�qo��-Kq�Rե�WUK|��jZ�[/��j�M<��2�6�6�#1V�x�m]U�ե�֕eZ�V�ڵ[�ږ�F~[(�V���x���[���m�|�i�<J�C<:��d �1�"c�zQTz���K	x�1�6��͞!���:>�#���ʢ��9�f���m3k�[<Zx|=��?�Hx�l��hf��#ܘ�����OL���=(�if�`ρ�0e��z�*����wg������ަ{�"��ػ�s{7������wN�i�L)�̘��"�jjmO=}N�s�/���tm�w6���}����}Ϩ�������tT��n�yͻ�S��Y�������=�����u��6#S��o{�&��41�t;��wf�1���(���@��.�65˩�Nwq��q�V�L�7�v[ ��Q��o�^��H�Z٭�_w�9�?y�C;�>|}*��W���nf}+�_��$��#����?N��� � L̟7��%��=������G�}� 	���/{�������ۻ�����I&��K����k����%ޮ��ﶒMkZ������<�ϞZ�DG��u�-O4��VqY��BHI0LU{߯y�W����&ӥp���Pt��E�h�����_��S�r>^I�b�V]�Փ�<�uc��|p>��Zz�����Ip��_1#�^�9`ė8{23C�I�(˪�۬�ǎ�]�9�}���6���A�;{0�y ��qc�C����$4t�����h��Ǝ�"7�5A��(a8�N�lEP�PfJr�Av��!�3끃��>;^vT���.����bb����õ�r����V�+M,�B�l��3@Q��|��#��Ǟu�^qKDS�.!j��xb����c�P�G�ǒ74wp�BHbi|OEIpi�5��Xw�Ebt���\��Q��&�c���*��f|ݖ�W+Voz��;N�I�$�/�tA�!�X�ծ]DY�ډa�ۢ������q:����|�ğ!th�q���t�@�լ�"�av൷�n���MUmb^B���W�L �q�:��f�������L#����٘0��󮵧c��U��O;�9a�ҍ�ć���6JvBv|1�I c�t�c�w(��8�N�����DG��u�S�F^i�����ir(3@Q�iƧfVk�-�1ٶ[[��{�M��*G�m��m��H&���^�JSS��/>,�5xDTS��/���3Ut��ř��b���J\��ly�1�9J2�6a�Sy.�G�-���#%���ǼՎ޺�z�-JeoW5�KF�:��z������yQ���^27�VV��旕�k�&����C�7%&1��h��IsX��v��F'��0���xn���$4�y��]�o	��Sh��S]������!�I��L= Ho����`1��é�Ɗ���\�7uTʹZE֑�����
<elb��n3�?T���H�2�ﵚN@諸ô�l�l�y�ȶ<�
z�����I-y	~��'#�^~���5`7i�T.P��!�U�{ã�5>�{�`$�!�E���C��i�X��#Ax�6PZ[��%��c4l�M?>E�8��#�먧�����'pb��ʛ���+SkcM��O00����5���9�#Ip�q�O�����GR��o���h`0�-�-&+����.�̩mӪ����s:Z6$|���4�u��p���S#�X:q>&đ� 7�Ha0�t��цp�+�&-Xwc$�VI"��,��8 ���㙭��y����55�kR���V���!Ӊ�	���m�/�DA�f�B���H<Hy%<�d�:���N࣒2I@���W8�^!��ˁ��xΕ��֏��č��bF�OG�}�z�:`�!�=$Rd�+TUu�-Ɯikmo�"#Ȉ먧�[/:ѴNg,<�v��S3"5E����@�ZS}>�}�K���o37�o�����9�R�A�b�q.���+��g��2O8II�@�L����aRG��e�zi:b��0��a,v�
���ܴ�lH0n<!�/Q���K$��qߙ�Fh}��|m��UR�ڸI��[AԢ�F��4L�0r�ć����㘞�'���ѹJC�F�DQ:q�O$x��K��!�1�Gկv�	{zq��bx�"F#�o��%S����bE��h�4�|e���I	)�״��ҪE��+)@ez�	�A��8�M���#�o��8��"#��;;#ӳ��E;��i�5j��UU�hmJ��G5	!$$����#�i61�����fώ�����i���18qldAJ��l�v��(n
��c���we�U30�U�3E��-���Z9{q5���]$���P���O�c�dQ�B�-]�hg��O��i�d18�N�� ��l'�&�,D� ��k�P���]UF����h��ټ����٢�g4��c �P�K��xI��%8!v���Q�F�!1����ޥk��K�L8A�Hh��C�/R�_)�iƟ�����":�)Ã<p�{~�3��ll��U2���U3r�2tMJ㙢]�.m��m��M	o�a�����rgv}���״���5ӵV�'0�g0X�f�q���:�z�=y^P���uX��gF�\���sђ�\��v�j䘶WTU����B�Ŗ�l����w|�B��?!l�9���N���jwzt$��>����yG6e�=�I�C�>8!���T�7��X��)h�-$4q�l�,3jI�);IN���#H�,�kD��lc;���I���㊚K�C*%�p֒�<V�H�6yh��S�ו+�r���||�6Y�)-��m�a�Ya� �	��=t�ѤD�=3�RA�@���Ӧ�AZ�iHy�*��6��0H!�a����5�3͡��#�)9:`��y:0�)��X��u���܈��V-�Jn��b"7��m��È<�g���C0f
DX�D?4��p�*��<`�a�:�8���o��"#Ȉ먧�R�uq5�S�c܅�ly���mH?Qʄ��@�����q�I�̀�L2�~U*�E�J�h�k�cc��H���6]�:F���Dlڹr��A�+kDR4���I/Ix�:M�9KA���$�,kڧ%"�����60�1����
�:�Z�1�a�DRX�~�����&z��j�z�w��Y��G�A��сiXZ��
b�{&�lKA��+[!�Ǵ��+P6��`��������h�&�������N����E-�������S�4�-~~qDF͝Ã6x���Qy��1�� �U�)��F��*򇐒BH	tK��d܊[(�Bv��o_�8�ۆ���Æ*ٟuH�"/�qao�����{֗�]��K:�#��)0c��+F0q�$�;M||���Oz ٹ�OQJua������y�h�5�[�KH��<�D3�#�X�PהXTu6�J.�ERq6v�i^ʤXX,�����q�N;��_�&���Zd[&�H�m�Kfָ�bhL7�$�d!�o�]V���WG"�'/f�-!�q$��D7�VLl�jDi�~mo�"#Ȉ먧�S�uN��V��L���H�n���1�bM	wH�SJ����{��O�ѴoЉ�#-E�`SF���W��u�q�)|a�5�H40��"5�%�Ү���ӻ��r�9�t:E�1D\#fV-��b��XmR�K��1kJ�a��j� bc���6�O�S籰샤`�W�Ó��N�<p�4Q���$	Ӏ��ӱ�)��u%*3��i3���ϖ*�#RFh5h�u80�Sh�*�ȉ5�D(��[ x��������1��r�(|FZ���;h���v�-
)h�d[C65��>"��|Cc�j�F�O�G�x�~!���Q:x�pͪ�ͪ�^�ًg�3j��R�j�en����SJ�R��⪯T�Ql�	�(�H�#�:-������Ս����Z��d�uQyl�-�Ե#�/�e�l�#+Sʴej��E�h�-��+��lҭV�imZ��mV�R�n��X��Q�*<O��a�>�͟������d���3~n��<<����eV�[+U��lڭ^[6�b�Zq��ʵZ��ٵ[�ڭV��[U���.����f���/�o��Q�?�3ñ�B��.�3�"���UO��e��z[��eKVUj�X�:�YU�9���=��=y�U�ޫ,کlڭ�ꭕ��f�i��TU�ѕ�ˋg��բ���#֯Z�i�B=(��J/@�M�B�У#�<�6��L�b�o��k����5��ћժ�r&�")ּ�G7W��LZVw8?��[M�Q��N*�~�������c6� �����3���';����A�����;E��$��3#w'v:��:�X��o����Rѽs�~w�.�׿}�Y?�s�[�Gܫ,����#��l���'[y���ߢ����[1dlθ�1�d����U�_ֳ���ʗ{쩩�Lz̸�ي�D��Pl(,�d��O#���M�,�9��_��w�>��i�^Gr�+TŒ�`��f-�8ejM;_=��ffrb�tb�Y*#ަ߿ē�N�q�� I��}������������ ���~_}��3?�wwWw}��H g�/��陟������ﾰ	 ��}s3�����ɮ\�y��mkqh�"#���yN�Ю�%�6�nR�U�8���W-��@U!��T��Ց�Q�i�"vZGbl�KJ�1�X�27cdqH�[�����d��Il�"n�lQ�j#m�F� �2�	\!�5+���IbL ��%�����"�#��!#�D�M��#	Z�G4K4Q��ʢ5j�R:ݴ�	�ң�;$���j�5\�֔�m�`��G �21
)��u��;+X���*h ��YIkzmH��MV�z$v(]RU-��������DY-�+�#�,����m����YJ�9-�Q�ܖ9CPU��j�	 X��5*qL-j&��;X8��R���[�Ub�VMX��It]7N9%VYl��+��%Q����Q骪+h�vȄ� ���P�ڗQרX֫r9qP�2���lll��r�������K�LP��KY�ʢ��P�B�Tj7*j��%�l�@���ET�[��+"z���Ա:��RV;G+��Z��a[-j��l��g1�chH�c�����߹�[�7�,�]�U7�^yĚ�@�o���p�gv""ݸ&�+b�)��waS�դ�6�+��y;�*t�Z�4��q�U��5=&�-�9������ۨ�����Mvr�&��ՙz�<=�9�8u��]�ﭜ{��,|���'[���{��/k�5�����4��b�@N<�yZ�;NE#��h�X¢��cc�6�&��Fq4˲ͣ����j�"0�%L,a�Ô}5ϳ�5Y��Z�56�P�'f�bm�)�y��x5'`���t@I�\d��d��$�Xz�G�m-�m���E��DL�'iێ��𘜇)o��q/�k����B�33+ط�5�PŢ�]�aH�p�q1�u�����(0a���#�jIf��ժ��2�/�4��-��8�G��W���������F�å!gǆ1�e�a�OGs�xM��0
GTJKC
�h�1��F��ʑgȈ�CD[L��rN��uv�*��w�D���gB�5	1jO'�&�i�����=I<x��Ζ�H�aC�CFac�#�Q_դ�5�
i��7Hь��iQ�qqf*E�a�1��s��ni�̶�5u�5<m6p�C�b ���:�+"����/[n��-pb�Ao�TUI�')�L[�Gd$���ӉĜ9�i������㍬�h2�l��O�"6����DGQ�Ã6x��xЬ����U�*��6ۍ3H�H�r+�1�cĚ\�9�yU*���F#G�?'
P*T�u��Ψ���6z��+��&�>��Ǩ5 �Hb�10�k����n�i�0�dsX�d8D<�����0�E�4�uR�gX���T�F�Pg��]�e�{�wB����6�����5>����lT�
N�)��i�姥�>&�A��A&A�w����8��y 4��)""�P`\C`����ia�|�5�G�C4E���:�g���wwy�2�M#�")�QJ�	-��|غbL_7�`1�m�ȱ�墈�}TSK�i�[|���ͭ�Ţ<����WP���]O�B:��[o�Q7�ጎ8�0� ƷJ �Ȍ�HI4�L1��_[cp:0�iZ8�(���H�TZimR p`�i=/���d����!Ya��ջ��΋�(��e44�-Y����v���#�8 ��<�QpI�:d� �as2dr���oA�g�-�"u<�(%l�h����B4Z�Px�40��8n}Cc��"�A���+�GF�dl��@���r����d�0��у�$�]��F��'!������l�����(�9 쀙4tX<Ϥ��)�`�/8<DSN8�ƞ~mo�-h�":�yN����V���|�5����+F��u:���CMW�J�+[Vk#����=`�(��{c�%	��}�݄8�������s�]���m�̨�SUs�]��ӻ94̥�9�*������I�Du����lw"���ͣ^J��Bj����K����Z��H���������SkgZ�Uk���Y�jH�wh�4�)�Q��}�N`˚y�2��tB2UkY���Y����g6�W)ʟ9��w�S�=qp�Ow�94�E!�A�pA���4�D�=�{���V4(0�S������m�G�i����9H���RL�-4q��|;oL�Z1|���rۡ�B����c"(���3fd��X� >;ƍ�x��<�)� c���Y�=���"&����!!��\��_���?>g32�|�Q2S|�^����Ql���ϑ�D6G8��=e�.+�I���tb1�#m��De�,
63��,�g����Z<���ǞS�-��u���wI�?�!�̻n�J�Mr�cq�aCE/�}ڰ[QB��]!��gE�%��ϜUUl�#g�����al==�ݻ��-­�--�6���`|��n:>6@��p�<6jP�Xy 珜��3��O���|���8�j�b��T���f�#7E�������(3}~�T�IU�f���_"$Ah�#�#� � ������g�1	}��%�FA�i����.�u���Z�줢��x06Ǻ=4Z���i��"F3��i�ߛ[�Z<���ǞS����Mv-a	p�_���1�4$�7�EQ�;�����LI�ε���0�4b�j���iQ��"8���G#%f�S0:<#0�(X0��K��XD�P�ZCK�"��PA�����կ��T9b�{̐o����oW.��^�CL����K���4/�� !�h�:��a��cnLzC�$��Z454{��0�kJ�e�҃h�Oi>$�a���	̑�0� �QAH��L��š��Ll
�&�.����U$�f!����pQ��5��˷OiD��9"�6h�yk�w^Z�,f�:Y������yG�<�Y�SY��z�kV1G�`�[�Q(�ϙF3,��0�L�U�d�����>���1�DN3㭱�4�B_��@H��U���30�˺˕o-�t�~׼p��!��D�`h%٣I����v�\'�m �]h�٤�ߖ�'�'�63�nH������dr���Y��v�uC��,`�p��I$ 7�f�3{"��D���X0�b[Z�MR-�"&�X���LR�VD1a ��_/�Fـ��D��E�i�gҰ��P���G�>~|�mo�-h�":�yN�׳����LV�٘�&���Z���c#� Û3]�:k5;N�eNK=��gg��l���پ�I`��P�O"��6�̘O-����s�gv<�s��1s ������M3S��Dׇ��f�ɜcmm�ՕP�]n��5����/;�UG�C�l�/e7���.�8)�墑h��6�E0*�FEt�ǒq��0ѸO<��d����}�a������G�f���pax`�,��R�~���iim��R�PA����J��n���n��p���X�- c�1G�5��b1�>��"2���X2S�Da哴��2�ѢO0�	8N�ԙ�>A�\��D���'�Ń����lLn��C_[�
KY�1��K�#�Sln"�P��,hw���404���E�KJ� P4S*�
M�"�E�gK8Y����֏"#���ꪳ��Uk]�P���8�7[�j=��&��:q�q�a��D���F�D4��Ϋ5�)�f"�e�����4h,h,a��RA�*+4��Lh�T�è�ي3
G�O"�X@�������8�ig���nE�%(�ؖ#jh��t��63�e}�"�L0a`�Ѡy�4Z�D��@���8���)�z�kW���OOY�J�MXa"8���-�J�5:�A��f��U�]p�=V&�g>�Y��	�]��L�:N7���%�3[4��H�rs��S�"�ha��t��a�x����o�g�����z�����<?5V�4�6�[6�֖ժ�ųj���o���?!�7�&�`�~M�6�н�'҈�#ӓ0�"#�=#*�c��K|�>[+Sj�Z��-]R��-H�i�QX�eh�ћTR��)o���3�V����=VߙR�*�Ζ�U�ͪ�j�E-�r�VUm3e4�U�m�j���YZ���Q\U��Z�[�8�Wj�Uy��ʭT�b�Z[mZ�V��Y�Y����ʖU��V�ͪ�f���VmX�-��.�Vx������Ɖ��%��,g�GD>���(_�L"��3�"�UW��V���Z�RՕZ�RՎ��el�Q��>�6p����
����x�z[V�i\[6�L�]UEZ�_j��霑�h�Z�ȏB���Z�B=(�(�J�ҋ�E�p�Ny����������4.Qsn��N��&W�/.�������,q���{�/x�ˬ��qۣ(�#�3��l�L�is�E:ؖ�i��eY{�Cº�ٯ��en�F�җjmc�˻�����}Qs������&�S�u����Y.�{����P�=w��V;N��[�9��FU��^b��뛝���t/�S�r{'�;T�Y]�Q��QPb���>��U�y�b���K,��P�?E���7����$ 0}��O�������� � �`}uU��ww_w�P@�몯�www_w�P@������ri�\��K�._<�k[�Z<���ǞS�9UT}�1�chJ}���*���i�W}A!�.�쓳W�eⰴ�0aj��� �4���<���4����CF�ޚ��J3D�����2�d�;#F�ɦ'���,���Qt�;J!���cP�l+����)"���5�OS�N��ci�,�F!p�2�,�Xj,bcH)ET��"
��.ǃg�;N��!�,��/�NO$�#�|TDq��b����Wwwq�tU�Ĩ�1��-�DY�|�A�5ŸRi|��ψ�)QX�*SO�[m�y�?8���y�6t�p�ͭH�e���42�q�2BHIi4q:|DVF���˛�ֶ�H|8&��Ğ� �"2�E�'�i^�ǈ^���B����r)��gv9�,�ųj:���yQ45��4i^:����D�`�H�B'�Z!��"�ac>p�;N=�&$GN�I�)"$>�������ⵥE(�7H�3��B�T2�T�$���V�(�*�5D"�K\cd
`�@�mt�j���P��$�)�&�4���8|W�����fm,c<4�"4k�F���6nH|;1�JyƟ<����ŭo"#��]]B���^�n'���ܺ|���+�T����D^"1��֛i��zM	��{r5Txi��I����.H޸������Y�z�M��ȼ�z�"��*%�Դb݌�����zߚ���]����as��f���vs�-�}�rrt��&o-|�/7�~��]��ڈɖ>�+-VV�]؝�MD�h�x⣑U��Ν�]V��4Ic�E55i�W������!቉�C��Çiۼ6i'Q��WƉ6��x�r3��3�5�pĻh�Kc>XDt�ϑGJ����G|r'Y�"""/��YC�Cl�=&T�����;�F"#����$TXhg�j�*Dt��,�a��xTG��үa�Ct��ג:Apֈ��(�2�����j�U7n<�cU1�JK�"|�c�E���{��4�� ���XR)�1:Gi�w-��>e�\u�����-�խ㇎�6t�p�͚҉�%66�r ���+�!$$��g��#"#(dDhf}���4a�q]����	��@�Y�*
�=�=�%>3333�ea�2f�%ѣT���C(��3�#f�Ǥ�*��R6|���A�9��+8��£�>ѤqidA��i84r�0�ޓ�NF�������G��h7�Ub9�z]����l�MuN�>�4F�{�I�l5�}1�`=�<��q���T �Z>DF#��DZQ�L�e��y��q��խh�:l�����3��o�Se��ʑ�!g��HI	" �^�n9#!ص���~�H�N���:vӉ��b&х"�=��hf���5h�i}E��՘r�P�GQ�<���j�=?����~�帬ɛ����,�v�4��ǰ�~��Ý{}kx2���F�a>:�l:�9H�YSQ0�я�i&����a�0(䓫#��Ҝ�:�÷��tU�{w�`썫���c4�(�f�;Xkht��tQ��^�O��7YVh�Y�9mc2ˌ�֝in<���Z�ht�ӁÃ6k�dXV��/1�e��
h)��H���HI	" �|D��,r�FDb�(34֝��i����1Z�sq��ϋ��o)�h�U�VTַW[����#�@�DKH`�lk���������t�Aѐ�,hg���2�a:�(����UB�(�Y��.6;��]��J����uYs*�/��>T��](*���CC]CGQH�R�ʹ"��3�.ב���*�.�)|ҡ��XR0��X*���4�1����󏟚~G\[�Z�kGQ��)֧�o[Γ��Y}M�[�A��N�&�NO�m��m�4".��ߣ�U�M;�S�fTK'j!��3�$�[yQ����L��I�(R���Q����*:�I+d|�6;e�:�9�9�?{��:ݹ��{���l2����y[�O}�msN����p����󔷱�u9y�d�f��n�\�L�����)YxL(�8�A��Y�E�/�i.�fލ�8���������f�`ʞaC+�xi�X�1�5��xDDmm[{6/6�ix�����e�Wi��<a��ｧ��Mq�xr���˧Ϯ��#cE/���7�&4T�z�x��:�c>0(P��|�o|6���I�	�l{�'3���ǙwWT�Jv�!�n-��C��"U�D��60��D6���"44z3���8R-��!��:ӯθ�����u<�9�.4�$ �ƶ���S)�����l��$���"�D7�EC�����#���m���'H�È���mqw܉�%���y޾�Y�RGC]���8�/�P���m�T�mu���DQ���E����w��ѥ;�ɲ����HcE�J*�\)j�C>G�ЍI���>��;�V3r<�Kl�m������s��Xq�).�k�7�iicGH5j@�D<P�Q*h2sG�F�e*��]��k�������,0��u��|�q����ִZ��x��uv��+�qlқ��,P!.��i��jH�3�y2r�JwW�3ˈ⯛c�	��֍e 1Br6��������̱ma�]ᶟ��24ݴB�Rj�EXP��1�������f]c͔w���<_���h�Ѓ/�mi���4�<b*Z(o�[zp�)mK���c�DO��
��������q�<'[0���M��u����CY�}�<�ݎ��2�6���T�������o�fV�4|�q��ߛq��:��/���Rթ�B<���5s���c&�V��VLze*2���HI	" �)3m���Z3F���!�oKҩ]�(46#�gַh�!l�ͳJ���@t��jՃwG��+��hl�QH�1�P�ˈ���鑺���)�A��7&Ô��8�Fˠ���v��iJ�6l�qP{}r���ǿ�uVs�2�����Y����f���G�v�����6ۓ3af��k>GiGF���6���pa���>g�,����>!����d'����W����~8O����c��BY��O'�����o���=��/m���C0t?B=	�#֣҉�#ҋҎ�}�n�[vC���p���xzԷYZ�['��іU�g[+FmQKT[>RԊ�"ٴfў�ϕ����mMZ��[�ڭV�W�Ų�Z��i�U+KfՋm�U�n�jŪ-�Wj�X��q�lz����;����ģ�|3O��W�[\T[;VUe���j|�mV�ڵ"3jZٴ�TS�g���x��F���m��?F׋!<�"="=0��#�2���
/j=�z[/K�?E�(�����霧6VǱ�p���vx�~�^�ٶٵZ�����ך��ͪ���3�8-��G���M��R�T��j�~R��M��������6�mu���MC�sϷ�0߾2m�/���j��[���цb�s��l��6�������[�ܭu��3�jn#�j��NJ}q���ީ���]y9i��ml;'��9�Jq����9Ӿ�Pѱ��tN��:�O��L�����vz�z#79`�ql\����z�w1<�
#�幚��sV8��錽:H�&�!T8��v��Z���y�����9�ݽLÛYퟝ�鿩|��H,�5 iإ����T��"���d�٫O��V�C�����`��5F��H@�_]W�������� ( � +���wwwg}� X_U}+������@
 ,
����.K�&�R�K�.^mn�խh���N��Vk9���ܱ�%�TLDU��i�h�x$� W'�N�B�6�i�v*��#U�F�S+Ԁ�\q�ꠜ�u�Ф���1٩d�RB�jj(	´릫��ӊG5]�
�W)5B�.��Z���v5G	S���Rڬm1**�ST-��m�GX��ޅX�i��u�:GZm������������4�($),U1�&)l�+��C�iPAS�ȝ��*�n�U��Pv4��JG��8�j��H;*#��n�([[��qب��iY!���e�ԭW�61��m-��)%$ ;-)\��-�le�"��F��ѻ$C�:�Q�rYU���c�D��u�Q&i�K`&�j)*�Yձ9P�ۊUJE-��XV�Sv�:�]cM��T�:˩H7 ��vE��ehn�T�We�nIj�UH�c���j$���+�4��R����4⚬��C7UC��ЬN�$j�#�X*'��Z!Q�����-�F�����	�v�O���m�ޓB��;ݷsPږͫ�߻r>��潛��F�d]Odn��5��k�"�i�j�U�ļޞc��&��+.�K�י�_bys�;���<��������El��m.�y����y���s�sP$`qɉ���Rב��։F��2\�p�(��p�%[�������ҳ��0�a{�5���}rBN!���1l���ib5E2u|Y
V��@c-��0�>��=2�6��B��B���;�tN;���������g��4C
2�b5G������%��0KV�i�!�0�m��Ǜc���񰡞J;�M�~����l�����|�Y���,w|��:��k�36p�<D[ogʴ�����f(�b��|�)w}#��m��ZS�ξu�<��ukZ-g����s�y�S��C0t�A�ol�d�f"M{]���DA�F��ٌ�`�ψi��4��-#Q(f��7�ה����m��a��[E�#��hڥ�R,��1sxx�e���1�*b�_4��!�g��F��_g�:諭�i�U:���C.�I,�E"����Z,����.�(����{"=}��'A�0�mR:������of�������1Mv�G�_)o�|��y��V�ִZ��]S��\�9�󗳽�P����YSݐ�BH�3��q��"��X2[�eQ+h�hfR1h�h�G���%їM��<�,h��ٜ0����6��Y�mF��!b��Tj'?,�H�-p�H7�%Uh����
6|���42҄2����m|,1�1bሴp��
�X��c���[�c$�����m�v�K��U��#�
�	�Z1��l��ѣ���V����攏�|��m~ukZ-kuĸ����!Q_1e�!���@ֲ=k��I	!$D�f�iY��scm2��|G��xiE�2�o�rH��bZG�g8�#F���
�Ee���fQߘ�*C3퍦�q=������ጊ�3#El��063]��[�t�6K���!h�6��9lc�\И�B��Q�s��V1�5f��k�ڣf�#���C6����k�ݤX`Q��Y��>y����V��ַ]:�ow�Se\Ba�"7X|����(&��2���$���"�7�3�����媅�U�<ɜ�&�y��9C�Qs���׽q<Z�콨��Msޞ������w֢��-���msM�w�p���:2�2*�t�h΍ov�ٜ�:�-�n#K�����9\Q�W;eε4�36ޭekU����H��b��J|ރC:&qn�X&3�ʅ篮P�=zM>�4��ãI�d{�Lm����h�\=OqÜ���oj�1�6�f�jכ��H��U������_�GW���,��yXb/ ��'�לG[M\jJٍ��g���6*��P�#jR��; ��������<O}�a�b߳��#�|���ϑ��������Ǐ663C\e5*�oQ��r\�BHIC�?X#�b�~Y��Ē�s��(��(��h�|L5�����1���s��X�8Duc��)���W�:�����*����c����ޭm
�P�ꤖ�tm��:��6Ux��#���@�`ľE��Q�61�X�f�����:aiH�jϰ�_a�\�|6|�|��>y~u�խh���N����Z��j��@QA8�_{�6�m6��y��B"EV*��X5�ֻ�14��yjCj�c8CF!��Z��,�����ϗ{����.3Մ��6����4q|b;��#a�>r�W#^Ͼv��.ֵu���ۘ��<}ߛoRC(���
1��H���Z���i��`����-#e��sȳFϛ�����E�"ѽm�7��
�����3cI�V�hhٙ�=�CGS�|���8���ZΞ<xٰٱ�+Z�yu���*>��$$��f�Q�A�FB��pgWNQd7}�h42�׍��:n��K�eC&I���3�Dl��Ѥ��D8|#���n)�A�1��m|�Y��c���^��[F�Ax.��TUBHB�W2���[Mi�=�&t�RI�#AC(�B6Z����g �f��m�Hoy�"�h ͮ����L���Ph��4Q��<���ukZ-h�]S��}�j��)��$�}�u�%�:�|R��+~�!$$��d��j����[��e�V��yZ&��{���5_zk����93��g�L>TM�a�l�v�|���8G�_�u.Z���w5�Z�yվ)���'�������+_έ��f��Tnۘ��'oWoo1��u|iչܜ��U�7_wJ��b����v�U@MT}�D����[Bg��ޅt����b���gT�ꨪS��s1�9�����b����G���y[D)�;��h(�v�����J��WwoN��Y��M`�l�G0y;��:���N�xA����/XWv�LS���3�����J1�N��٤Z��P����)�5OV�*��#v��D[1t��(gW���7�{HԈ�*��a�(�J[/��mo��n�:�ִZ��]S����T�3F��5��K�5l�Z`�6��3��I	!$D�UR�� 1�y<8�f�e����2�{��^��
�������Oh�� f�8�Fi����+��q7E�=�
z�f�+��nFh��U��"���_g۳+�p.cY�F)�rf h��'�Y̼�:��1񶛸�(�U�&���l�(��<�i,�<�#T&�
gi��qY�u�XY�V����io��Ϛ[JB"#H���:�����GZG�GF�2�R�!qgUQ�4��DqGQ�<�#��<�#��<��<�!�#�Q���HDe�G̢2���<�#���h�6ӭ)�2����jUb#lB�[b��W!B���J�>G�J�iFQ�J����-e��K[+ijZ�p�"�u�\[�yky���-�"8��"#��F�eB�!�&�û|ڣ=e�a>�L�a��������k��Ln��UU��^�=9㒱�X��o�T�F�ۻ�3��f��j�^�o��NFXv⋳�U��p�w�pι�k1��{﷚�g{x�h#�84=�=��3��{F�B�&m�{U���Nk��SZ��UU��r���g:���׉R�.Y�I��d��m�T�v��bz2#����Ъ��,c��Kڥ�׳e�Lw^Dl������d����Y[�y�pH XU�W������} `%U}_Gwwwv�� �P�U�}������ @UW��/r��(\�J�ʗ._.��V��֎��e���o9g9fBH�3�>6a��g����*��Pȅ��E�,\��օє�FZ>>4�T����Z�D���'��R8��*�R��`����6�.��BU�X���
 �C6������'͝aY5NľF��$0��,Lg��i4Zk��IŻ����7-<�<F�#�ǳ���{�M�=�a�e2��qm��Z:�]Z֋Z:�u��r��UPҀQ&>c�%�bf�z�X��BHI	" ƴ`q:`ުS���H��ߎ�gQ�C�����e �����؂�#2��e�s�X���S�Ks&-/Gi��hT�6��/ڴiM��{a>q�)�����Zx���e��iTV3���a�l�42��4軹V�ʭ%�6N*�{���8p�0eu�k���i��qcV�F���i��<��L ƈj7���W�2��A�T�͐��M�>Zߝ~uխh�����Y[_%�w�Sݐ;Z��F]��LXݱ����HI	" �o�O'�ө���l��~Ǝ�N�k��('���r�f��u1�;lJn�R��"�t�'3��ogg$���s)��M��e�,Q�S�X`��@N���nf2��"���1�uNq+�c9�uQ�z�靗uS4ouT�n�^�Ӹ�W���^i�y�2��j�H֮o�E<��FZ/����c���a0���J~��'�η�����3H3y���m���;��3�HE��fȉ�k�"<���[+݄��"6��p5+Rk�:R�~��^������ͣ/�+���bo]ó-)��"�una�r[���%���z�4����yN������h��:�ִY�͛�7������G%ݡ�©�o��$���"�"�.4ysAنF����P|ǰ���Іf�9�"4l�<�QӬ��G���ш�Gb)^��a��|�����m�M5(���E-{�U�[�q���W�ǰ�������;��ܥ�ɜ�@�KW
�/�x��44���G�:4ml>�6�J5Շ0�?bcxL[�G1��=���;�S��F+E|�9�>����6`͙qm��<�V�Z�kG]uN&�����q���(�����To�BHI	"!~�N�_�ضNF��6��\�I�鼼��e:�>x<+����1��LF���a�_�Q���}���ɹ7���n�uMv�~��|�l����f7�ag�Y���g��w��5��Fբh����k��Sc*�_m��6��>zՐc)`|��=�i�a�^�:|Ҟem��?"�~qխh�����Yq��F�&��l�+�p�BH�Y�Ə�cf��Fk�H�,�9oÊ�V��+��gt6qϝ���=YW��2S1���חX=#�x!�j�����䍏ϱ�#^�x�4���(���
�6ut���8:k7$���J��?a�/��e�;֞U���:yAH�F��4uij(�Y�Ӯ>D~u��V��֎��emB/��WʹU��S�rN�p���{�� ����s��BH�sw��{��r,�÷�S�W�{[RB&�v����EU��L���ܹ�ܵj�v�:3+ë��c��2Aε�֗P�EU��$����R�jۼ�ѕz��6�B�	�{�̘Q�=�D��ݙ�nm��ڮJuform�,��h�hރi���t��/��iK������4����A���'J�O#�ƪp>]P8�o:M����>��J�*�T���#���OX@�Z"8�����TR�y�щ��v.�0�=HJC�2ˬ��ck�mT]:�
:�(��d��3GFR��;UY�kXe}-�>e�m:���:��Z�kG]uN��v��*��]:4���$$���"\!H��M/*�A���ChN��χx��d>�5�/	x�b��ff���w%]�ܓ��#�V���l�JSM����c�S�n���,E�Ta�����]�Xb��οXWܺ�X�їY32�R�ᷦc���n���r^׵��]�GU�YG�Yq]G8|4m$�6V䘳Af��J*4��c��ah�#K����1,G�Ό�<Q�Z�~qխh�����Yp�V�,E�֡$$��͊���a���IS�M��"�!��o��5D[1l��#s���жKL�ų��#��p8g����N�;���M�F֋<��?�!�hb<�.ͣ5�M��qb��E��b����*w�;峈
��U���m��cF�lѵ6oՁ��905X���u�eO2�m:���ո����ǎ�6lf�h���6�t�nL��pm���HI	"!:�p��}��F΃,�H�ؓb�1�:�F�ZG~�	>�u�}�޲�zֈubg���~�d�H�ߛm�ف�&w���GQ��|�>�yv��Q5}�T6|���eH����4��4�1���UI�xS��˼Kh� �-�-`3�>)N+��gm�663C(;�m��|��m�GOR��3D���<�+��ϟ�S�DF��u�")"#��"":�u\Ge���!yi�|�#�F�G�uS��#��:��Ȉ�:���"�����":����>E"#�#��8���{��8�攄u�DGQi")#��!�DqDqO��>ieFQ�J�LJ�C�)���Զ����qju��qţ��(E���o��������q[F[S(B�!���m�t����A񬫙�	�]�+�2z��-F5�4d��>�؄Q���Q�N#��Je��[N9ي"'ao���}��r#p�]���FZgJs��/�Ց=>�u>幝k{���E:NL�'�r�����@�]d�:[3n�=�x�U*ƹMJ~��ժZ��-�ۻw�=_=ma]����y���8d��^�ކ�k2U�}]���tu�GFoKd]¥�6�ɯc1���~_	�_0Y�+�fcsRVZi̪
�"���[��O\�u�YΗo����;���  �	*���;����� @$��������߾� 0	 ����wwww��  ������r��(\�J�+._-[�-kE�u�:ˋ��U���YQ�%����Z��d@�"���E[��	��Ӥ�鐮F	wV���	Qn(���E%�����j
�Bi�%�Pd�Z���*W�hn��N"���7N�bz��c�5uY jB˪�c��C��@d��UV�"��N�J�7��hLP�zwU����!�+��*2�F螲;%��vEX�[�m=�4"'(��LU@�"�١�r��A���K^�i�1�uDT���Ul���*�vWF�+*��R�ƆʫduK�J(&�v�9*eU֚u]Y��U��&���@���[H1RD�j�喎9���̮&9b�5j����B��,m��1MY���܅�Ԅ��@�SRI�ꌣU����;#h�A@u�&�����P�ڈuZ���1���Ȉ����V��dc���A\qW[5m��[+(h��m��d@�	����Bj�[B�J8���CQ�V���6��c�fuD
ES*����UEjb����nUmJ��8�n�%@�5J�j�V���Zm��m�5sm��fE�[�`��[^��ڛ������⦪ue�.k/:��$��ˑ�*/!�\�a���e�en,OWW\o���sml��fb2�?m�V�P�O��	��9)�	N���y�n�[��3v�KԺ���Y	�a�yxڱ��6���ఁz����Za��5�D���^k�R���<XE�3�G{�9Ww�fc���x�k��p8U����t.3�`E��aE(����<;�0:4Y#&�,������/�G�sL��g9�oc�u�7�7x���4���6�8��uZc�mƔ�NiM2�m8ӏ��ο:�V�[�N63d4t���"�Q��Iq��]�8!r�����T��F��i�����!j��k,���-x�>�{44l0�H-�G���
����0�4�GgaI�q|���/�����{���E�׼pC��T�@�צ���G�[75�:����6-�M�5ު���g����+]�����h};a�!�E���m���gC~g�F�Wx�e��Q֟�q����֋Z:�u��0�v�ʳY+,6ȹ��HI	"!}�r�G#�-����$r�����{C�yE��˧4��b��������1b�����ͤ�8~4���=&�V_9nܥ�*j��3>RCH�>>;h�#o�����<Sp}DT�kۡ��Xe����}���X�Mh���oR7^b��of�T�)�>8��a�ٷ�/�ӭ#�[��yŭ�lᱛ!��ֳ���w�s,m�z֌6��MQ��ƛi��zMD�	�����f,4��C���#m���.�U_ŒԊ���65��{�i�\|M;��y��jLtCZ�+M>���vq�rr��Q�QH�"�h���٤oK�qy1&w��p%��E{s��r�n���хL�IX3�d�6���(�ц���Z�^8�ae�1<��S���N��^[��yŭ�u���ڼ�&�δ�X��̛�$��&�Z�r;���m6�oI���L�>�kr^i[��-�R��[����uv3OoI�
�z#fc�']��TƑ��̜���"3&�)����>�P��ɵ��R{��͹�� v���J^�,G{֯f��\Q5���]H^���f.i�v:�R-�h�ೈ�F�ʱ��ƸJ@��'J����D:B^<a����M����kqd�B�D=w&����w�{�Y�L�qxk����;��!��Ƣ�7��.&���R�Q���[woZ��K&����|Z�E��<J���̩�[u�i��[��y�g��<t�Ã6CCnji�$v���-eD�Բ�ԭ�<1�;��mI	""k�ՠ��"[(����U\)G�
m�R�r�ֱh���Q���u_h~84,`؆�m���$Q��|���gh�iy�m��V[V��ʋ�#a�P4��P�6~�Q��MR �,qB�E�����5֎.�A�|t��)|�_:���T'C��喸Ck�?#���6Z��@�{���`���N4��GV����kG^yN�h��jE�e��߳��BH�gQ�`4a���N���<q$4t�A�	���gƾ��=ѳ^CD|�|;GC�1��s�T����7W�{���{��n#�N�I�.�"E��������Ag{����dL�S�4��Z=D�-�#��(�L���f.a
Aut��#�;�֯�I�ⱣH�Y[�8ӯ�-խ帴Z�מS��ީY�U�y �TH�2sZ���DCk�,��l� a@��>=x�R6���>:��A���Ꮗ6&[��t83�(:�83�pu@%|Y���l�X����AK��7
uR�#Fɫ�4Dt:�M�H��.--�^�PJ��
4�8�Ͻ�{_�Cng��Ǜ*d�X��9�|ڟ2�<Ө���yn-�ǎ�8pf�h��|î$��>;af9Mj���:��8�
�4���mg�i��i����!�z����������G{&�l;����mлUozh}{$�j�{+:�����e���d�D�T��P���+[뫣/.w���M9Z�m1�9��^<��Q3��2oo�wj�]���g��Q~���F�U[\��onm7����Uʹ	D���F�ǥ��>�����
"���9��6�\�B�=�|;ȫ37��=~W����g��qS1��Upv''���w90����#F�Z*�,t��"ҁ��Cw�+M�M��EԪ������rܓ)3m�����m3k@Z��c�*�Q�7yγ��Uo��4��y��iמ~u�o-n�֎��e�խ�����s�U!L�m����BHI"}�9�6݆���q�-_z�n4pg�R_G�rHyu�����w�
G�aѣoOb�4'|�	�vbjh����h��Pdd>F����)C8�#���rB�o�R�������r˦J�������h��V2����!��L'�A��y�+0���p�i���e��kK��K��q�|�t��;��9�q�̿)��n-��|���E"#�DDye�DGȈ�#Ȉ����h��HB!B6����TiDm�rUuG���yG��y�Q��DR">DmF�i�|��uG��m#�|��>R�F�Du�")�mGDDu��8��|�4�4�#*�X��X���"�l�m��K|�N�㮸�ye�DGȈ�"�kZ�mm�����BBBBB�&���X�����[�ۈ[���ҘM���$F�q�W
�N�b#����5m�[F�o��*:#I�8Kֳ71�+&��Z������,μdF��]vN,s��)�2�z�Z�;ت��8D��uÌ��DD�Ȧ�����{}]��-�#�r��"��l�aor"�o%��ǽ2�V�gk����(S��;5�yr��>U���g����Y[�p� �$ ����k��������HUU_|�wwww��  Ѐ����wwww� B 
���ly�<Ϫ���<��ukyku<t�Ã8M7"��I	!$C�6�!&#H�g�f-UF�����.�m8GDCH�bi�Dy���鹽�aߑ|Y��h�3�.[�ܩ\���:*bw�vH�;���>GC^H�uZ(��4�ih>]߁mW��Q���q�C�G�GWC���1���\S�쪩Vql+�^F�ݮ�������8ӫy��張��Z:��y�+3�W�(pM�n��f	n��Wz���$���#��ocϛ\1���Q��4��7#�19>r�[썦fDeD�{WK�� ��U~�sM���ڰ��H)���)��0�6��1��B4�����;��������
t�S�%T��?�����-��ͅm�c�l�h��ഀ�����h�0�g��5PL�4��y1��T�2��<��<�_���맏6p��)u�E��yv�YL�T�V���dTK�ƛi��zY����O�0�}�w�Y�pw�e�=dY�:����7�:��T��Y�PV��ۍ8��X���;��E8��dk���u�%3e�]�eƻ��AQ>�0���O/2��t�+���v�V�k��:�k7Qu���-[��=ܷs{�q�pǏt��|F<*��u����"�b,��u|z�w�6��m����ͻE�֊�p�Txu�h|m|�G�X�1>E��A�����^^���'[���x:��v��k��>�}�Ԯpl��[Aa��üm���ɵ\ C�c.|�D�"�X����K�\�-� ��jm��y���yn�o-n�֎��e���/�l�Y���̪��1ݬtƙ�^L�^����Dh�����oih�Ό�7���}�A�㍣�ȴ���ꑦN�>DU�����sL��*^+�P�ރ3N2=�z��7+熳E١����qs�/�q�h*ϛm����v>\[zm�[Gi�m-U�ǫ��ǭ7����\i~~Dukykq�u��<��sL浜WtJ9��I	!$F2�h��#J����QhĨ�Km���h��VՑ���$��t6�,-�>�+e��9I?Gc���]M71o����.���#g��Ӡ�\���e&S�H�|Dq�����_!��}��6}#`�e�E}D�������r�(�oeio�G_����-h��)�yUx�6�W�h��*�����$���#<��Q|�)l,Ʊ.#d�"�+h��%ĘA��?���!�d��RI�J�-�XC�hm������ ��c��hi˪�p��o�k�;���Tn1���d��^�.��>;_<�lב�#E'�M�<N���t�@�>F��GU�16�qk�r�/#��p����}M�v�Qh�]
(o��WZF�~Du�o-n"֎��S�fsYl��M�r}��l��X����\m��4"�����{8�m6�oK�}�{���kv�<j���Vj۵k�sjr�ָl��V��Õ��jM�P�^uݪ�.s�"c�O���s��[�__N޼���;!$��F\�ɽ����#��F[�����q���U�6�cUt�/bC{H��4b�w�z�R�7�U�]�����sJYŮ7�y��Ю�m.��Q��:Z6�!o~�$��F��u3`o�W\�W��\Cc��U�ӯ��Z�u��E:|DX��&�F��4�m3i��UQ�S_fU�R�/2�~6�<����������${Yżo��Jm�Uu�i�[����������i���F�	Tܢ�	!$$��H�,��6톹:i]V����m��t�����a̦Z)]G�t�t1f���x�0�Vo����㎃��^i�=�� 6)�E��E����"U??�~�����o2�ޛ�Y�0�ңf#G�MR]
;�l{��FF�ú�l::5�H�i��"��ј`�2�ʨ��D[�����qkG^yO'�����dA鯺�V�UX-�ok8�b�h��/u��M��ґe�H���"#G�>h"1R�a�հz��#�*7L�Ur��:>E����'ܜ�&i��jfe�TEw�cm�!�86�w�D|4��8mh:ѣ�Q 6�H��}�r�F#��}��U[.���߸�.���7�L;��+����-�6�Uƞ|��q���qkG^yO3�j}%A�h��UE˸I	!$F�=�i�Ѱġh����h���9�qM��m�5��|I�JR3�Ʋд]c�R7M:me�4Xџ+4��m�LQ�NW�p���k��>?8��l��T���H���-�>Tm(EGW󎢪�'��<�u�7��k؛>ﵲ*4n7�-��-?b|�ø�+N�˨��|���u�mK6�DDye�DGȈ��Ȉ�6��m2�B�Є#�ei�4�#h����Σ��<����<����l�#(���QH�(G��#�w*��H��8���>G�8��B>DiGYB"��Ȥq�yF��>Sϑ��F����eHLJ�C�bH�Z�-n�O���]q����P��D|���<���k[�q�VʖYe�BYL�{��{w7�g8�,�8���A}��W�=���s�'�%}�^N���][�W��j��7��H���q�ǓC����϶�U�U�WFS����>�j��g��Q��}�x�.6�F��K��'#��8�����v��܇�a�e�,�*��e��LaXe^Nf,���Ҧ�N�tعt��͌S��F;m֫����s��5�[P�#m-������Õ�ښ(�wnv"zmʹ��X����3N���������r\z̺߮r�Nw�_�j�{Xgø����l�m_?��s{kl|�{�3x}E59��L��-��FU��R�W]��4'p}��H��j��o�TeKr���������� � UT}����� � UT|������@  UUQ��wwww�  �UT|�.Mr�+��T��q���qkG^yO8������xJ+jQǫb	FJ�Aƛ���cB*���@�Q��,�FQ�ДTUҩ���%�A�궨tN�b���m�P�q2T�A�m���*Z�Pu��U"���;ev���i�9�(��U�Yט�h��,Q��`�\v���PQ�	%�Cu��XFӢ��$���	�P�RJ�r��PNTHݢ��t	�U-�v�-F���$�p+B���d+@8���z,u ;uU��m�@U;E"�DF�c� I[U��u]�J��t���YeM�*F����j,m7a�G
ޣ5jEpN����(��N'�%*�d���c@�tW]�Sr,�+V�
Y.�4[J尌Bq(F�=(�ac�
�6�Ԗ6屧c��e�ze��Q[v�Z��V�*�c�6�%l��T�EDu�� �0��V��Uc�RYUU�h�6�^�%lQ�@,"��aJQVԲ��%^�Bb$Ԣ�LmEKBj	QW%oChEAl+h"a*	�-C��;\`�rnI�
[G[%MB�S+ې�BH���j���]OMo~s|������qe��k�œko�����$��������}��5��:��Q�y�v]��&B���}�Gk�Y�U�H���V3�;w��}�E��Nw�|Ym���wa9Ï�V�.����[�F��M+�ע�͞m����h5���d�"�ȋG�֎�A�C�����Š�N���Ϧb��˙w9��&�/�7ѳz:����N�h�B8���'��4V+0�f��R(�m	��1��6kH��=w7L�9��r�̢T3i�w�_61�C�1�G���
9Ѱ�Å)���#�����qkG^yO8ӕw�6+�%�'-��rԸ�e�E��Ҋ���䃤� {��&�n8���r�]T�i�1����k��|M��G��#��T�XPR����rBlņ/���~^_-�a�b��E��aYu�fK0�1��&�O��-i���GV�A�o�6�<@kH���4l7����1��UU�~p��4���|��q�kykFִu��7銧�ZKJ�X@ki���G��hſ9��#H�9��AfCaD|��Vt1qZ�g�\Z\6�7SiyZ�q3|eU˾=�Yz���9P�33�W\�QL����qI5�9�#�{nMxK�Z#��U��F����
��m.�X0�g�Ll}�JϤ�L�t:PΚ(�N�~Dq�kykFִu��+]�7�.�k��o6�L��9^�ow�
(��v����e�����N����%��W��RҼ��a2� �1c�3#g�=A��+���F�/:|h�����h��כ�ѽ����<�T#k�.���$,Ô�;��f��i��"�vNME�,<��>(�Xg�E6�L�˸��)�|ӭ#�������מSδ�޽U�ޚ�>Պ�ؙ<5��b�B�ȫ�>b4��o��$T�E�������c�:�G�o9��}���x�El�q�SќȤŦt*�����f�t�7q�ڸ��T����Z��n1;�h�uBȭ�\�i�6�*f�dsY�2T^�qn�ߏT����̻���d�v���Ֆcl|>Qx�8`'�شot�º6����TsC���~����b[��ʒT�N���F=��^FGA��=H�;���u���;g+��9	s1p9��DE*��y��99�t�7�̏3U[/z�˧XH�u�s{ٴ�g��Q@R=�]^-l:-��rO���|l(�͞4�-��G����[�G^yO8����.d�<�s{WY%*�-�h-��/2(��`�p��t�O�!��F5��||xx��6l#��W�Ӓ�FJ�P��iN}z_��<m��|�L�4�k����'����c�8����OH�Pu��a����S���6<���ղ9'�Ҟ���`B�:�3�\��A=;�\�k^Xiix�oh�a���k���്�>5C�h�*i�M���Dqk[�Z-ţ�<��i����ʳ�"��K!$ũ\y˘�� @����:ꪈԧ퇃a凗�\E��xk�xZ���H��6�!�a��ϞH��ם�V������/5u����4�)��,+6Z>�7�Ϫ6��i"S4XE߸��&�F���p>H	��9$��wV�Cg�l�p�z�Kl�"Ls�L5�ܣ_��M�Sh��[�?8�����מS��9��9UwT�h�ޱ���qC���9"��v�v�N�hwxÉo퍽o�ʅBR�+X�]CT�H��:u���$Z�"*�H�t�������?1�_��bi��hѡ|t4�rF��άAJ{�Lp;/^%��L�o�a���_<8<�s�����kh�Zq��E��S���H���������Z:��W�i���h��oh���8L{ B�pB�ޭ�� �q��U=�Y�>����q��v���dVtM������^���d�d���S=�qX���:�"��Nn���/\�u��9�Jrs��V��bn�Z�\�o���x�Wv�JM����1�[�\���wzte�M�l�m�E�3��kx���e��q���5�)�ګt��{�{�ˋ�e8�-��H��̶z��4�,�(p,��V�ڮ����|�����+�~�	���qLF�a�r�QRi�S!@Z��\X�PiPZ"1Q�7մlC8i��u��[�Z�Z�n-y�<l��vF��6�'v����գ��0>�lo���7��xt�,%z䝅-tju=/��Ub�sܒ�Շ�(�J��'��C�!�N��G�n���<�t5��,� ���o�`���?��Wq���Nu<5�^��v�>$u�����BW�q@n��oG	��v�>�zt�=o���x�4˭���Ͷ�6�Jye:�DF�GB"2���:��#��h�6�(�!BDS(�4Ԫ���iDu�]y�yG��x�#��"#Σ�����>DDGȊuHFԈ�"6�D�Te�q#�|�摥�e�D�TDG��P��D|�GDDu�mS��-4�#-2��!1*���E"�E"�y�u疷��P���#h��<��:�6����ie�Xx<63���ͳ��k��+$ʿgk"㻃��ŴN>w-w�
U]w$���wS�{Q�w��ڢ�Q�yw�X�\D�~��bE0�S���c+7����|���Yx�TV��;q9,�Sd��ׇy8��5�;�{���%ϧU`5�(�ⷯU��#���Yw��K�Un��[{헒\O6�׳q�3pV^Ǟ����Ns0_v���*?E��^���W%{|Q�F}��� UUG������@  ����}�����  � UUQ������}�   UT|����<�Ϟyn-�֋mhl���6QV�q��E�x�UJ��A�#ވ��mn���$�_.��g,5ZKk�vu���iyx(�K�Z�Oc�#|$�=P蒪�,��yh5�#��iin��܌M�A��R���Ϣ=B�{�܌c�qZ�-������|��b7�c��iN6��-��-��[�Z,��M�83��9��Q�8��uA��_5�I���tv�EU��O���K�K���rM:R�9�BH��FP�
Vt�g��I|s�y�6�᥮g�6�)��Ӑĸ��G�UH<U�,F�,m�acF�>=�T�>H#e�cN��Xۮ%%:�p�R,(��l��,��q��֋mh��)�Z}�V>�G�"Y0N:�4�q]׾Z����CpB)~� 2�}�Ӑ�\��y�GD��o}5�SknQre�h}`�9�ky�7g2�OwFC��ѫn��[77��:}��W9�d�қ�NeM�vӝ��#98Z�����:�!ex��SFF
�m����p�U>��B�oΊ{[�3NQ�Q�]-���q����gX���u4}��G��`Qf�!���W�9A��R�Ke{�J.��,�d�*>�E��,d�Z�E�Kk��X+��^CP6���K��!����R�����n\�a���Ӡ��=檋n�:���`�&�e�#��<L>ٵߞ��Soʖ�O4���~qh���x��M�83��4؋g��Q�4�"5�=�B�3�x�z  �il[�#�Z4^/�ԓJΣ�ZT�>:���9���+d�M�i{J�>�S>K[4�� ^���6�F��Z&G�U{^����9��$\;imyV�yV����ƈ�d-�Ӧ���R�-QҞ��7
p�h4���C���x�a�M&��]���������H�
i�i���#�GQkE��yи��������'�9%	�keBe3�� .k�����v�:�5h�biԢ+��8�x�_�zN����M�#GXZ�Q�2ƭ���p�r66�JoK��(��;����������:���V�w/���q���ȴ����Ya^G ޏqpдT:^(�Z9�S�\G���}��:�mP���#��4\m�x�m��F�ݕ���:�m��u��n-E�t�G��63f�)*q���WF�Ts'#m��C�ƌFpp4Z>��[Mg�tԓ��W��3�5�e����-E�>�˅9�qi1�g��#渹���,�a��Zm�_.pٞ(�Υ��߯��ݷ{�m;���B�5�-��I�Z�~�6׭^�_�u�a�^i󍣶h�G��#��l[���V ��up��Ɣ6�,!a�(��[���"�l�uN��6�W�o�1Њ���0Њ�K1\P{O� z�[sN��/����������#���51��uN�ӛ�z�n'8���-��0��1��]��Ef����9��u>[y:�ml�#���3����9�̝�&;^�!1o���܋3�&=	Z����ۆ���t���8�@�+4�;(���$��z�)���9��!�#�S�!�f4Op���)m�v��'����'�u�S=|�q�M&|l�O#�G�E+�lu�<���0a�F�_��-a��u��E��m��$z���������9��MT�Cum�"ө1���h�P�i�IJVk/a��<q�<��m<��8���-��y�:�X�Zg:�}��c��x���eF� 
�?i[@o��e��L��5�a���z��~���JZ[
���K��W4����Y�E�������ӈ�-��(~9m�8uh�w��w���GT�E�������w����vI�.�{]�ц6|��I�ml����)t�:�ż�)���N���l����/�u�u�����o�?#��E�p��c6h����Rۢ��U�F���m���M@�D�܆��1�4�ɢ��{UQ�^�OP��Ǵ�<<�#,�G�R4m�kC[��1���������"�μaѺu	�{W��o	m�{sI�=��)����ƚ#kj#�<T�BÇ���:��[F�5���������3�E�#&��ZM��-|�F��3�c�ZSn��N�~Z8�uhx�63f�d4�In�ܷWm�U]�sm��"�j�g�s���:����Mj���`�erT�e���*[��"�F�qiis�i��n5�aH��6yDlkH�D5��R-yC�݋���;ٲT���7�6Cu���5�q:a�x��mF�4�����ͺv|���������}�CI_uUUT� * a�����9�W��͟�����յѢ�0�@�*�S�#��{�&1��:؈rH�+	#� �""b�a
����`�`��B`��&`�&���&	!��B`�&��!�`�f"b��`���B`�f5��a��h&�f	�`	�N8L���C0I�@A$D@A1�D$DI�D��D�DLLDLD,�@DID�D�1�q���� �"$�$��""a�"b"b"H�$��"!f"$�"H"�(f	�&H""H��%��""H��Y�"H��""$�"Yb�"$��"""b""X��""$���SDLDDKD$D,�$ADD�$A1,DIDD@DD�LDA���D�,DI$DK�DD�DIK�D�LI��DHDD�K,ADD�,DKB�đ,DK�$�@8$AD$DDK,K�DD�,AB�D�Kı,A$Aı$DI1$IDD�0�0p�$�����	 	�b ���"b�$���� �"��X$�����$�b"b"s �)����$�H�H�� �H�$�"HX�X��"H�"X$���`��a� �X�� �("& ��������� � �$�`�$����H��X�b"b ��L�q�H��	 � �&"	�"H"$��	��b""b ����& ���!��f(	�$�����He�H$�$�`dFFT�� aHVV������ `BD�� `F� a�0� d`a�� de-gF�0��"� `XD�� a�� dR�`B�� aBP�� ` X eXR ��`aT�� eT `HP��@��HP��H@��HE aT `VU�� ��`d�� a dXR@ dHQ�� XVE�� eFQ��``�dXX��`d��``X�d!X	FF ��@��H	��HD %U��H	��H��H	��7�DAD�@B�@J$@@@J0�)
�Ȅ0,2��0ʄ0,00)�
� �*C+0�CC"C+
J�*C CCC C C
C#!
@����#$2�2��� B�20Ȑ�������) CCC#	!�)
@�ʐ�C+	�22���#
@b`�C$1x`ɬ!�R!��He�Hb�XbC �(�!�d�d�!�� �H`�a�b!�b!H�!�b�!�baH�Xbb�Xb�RHa!�!��!�b��d�!��Xb!H!��!��Xba�RXba�e�Xb!�aH�Xba�e�!��XRd�!�d�d�d�� �)$0C$0C$0C,2C,1
KC,2����
A��2��A$@�A$�IA$���,�L�@30D�DIA0D�	$A$A$�I �$�LA0D$�D@KHd+��H@II@���IIA0$IA03@2A04A0D �@D@3A0D@@A�$II@A�$A0�A0A0I0D�1��2A�d4	AA�DL	@L����@�ILP$�L$�2@D	02@�$$�2AI�`��G$��H�$��H Y��HH d�`����HH  �H Y d��� �H	 ����030�ȷ����03 �03D��A@�D00L3D@�0�!0�4@DA0L0����1���G&��3�e���0NL���}/�¨L(�J  �P<D���P_g������;�����g�O>�޼��������~}���?׍�O�k�?�͟���1�y��|����Oʜt}�O�z>�������l�OՇ����O��g��?����O��/����c������������?�D�z��%TP�,���	����O���#�zɂ�4��	������?�#�~_��Ԁ~?�U ��B����_�*>Ӥ4?�8������~�D60�O�:_���bb~���n����=v�u�	�?�搜o��&���qj�����s��\Ȃ �գJ�ܠ�d�
݀* ���0J�z0 H�J(L�$H�k�o�P�.7_3�L�c_��N��0��������a�hR��P ��B���u� �@D��@��Z�N@~s�t�Y���~��/Ώ��=����F?�G����?�?����5\���
(P�p����_��_ཿ�y�?q���������CݙЏ�?��A��>�a�D���$�����`?g�>��?g��A��K�Ъ� }��b���w�?���ã�����X� Pe��U �?{������s�l��Z��8C���5����xHS��?�~�����uDz:cO۰�D��@*� @�����p��Xl$�D8�3����4�^�q<=o�ΧPl����/��{�(��' ����?����/*�����p'�D������_�?��N}����'���K�O�����_����\O�~���}���
~&�����'�OSoR�(�>��Z�~����o޿�U ����O��;�Z|?�>�ֿ ���[��/��=%p�0~�?ٰ с�v7��.�����$?���P�֐���&���s�.�p�^{��
��)�E���~�M�D�z}�������ߦ�=�~����﴿3�M�p��|=?���ȧ��'�J (�ٔ�}�j�B����	�N�@Q��6�����1y?y�1>��z�8O�~�??bfi#��a������w$S�	N��