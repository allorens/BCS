BZh91AY&SY�sߍ_�`q���#� ����b%�          �                                 %B�B@T�X �I�             @                  �}R�	H!@�����(�DT�I�U$RH�Q)
IHEBH�UT�D�����E!_:Pe��$T���B�A@ �� ������B+�(�͝T�ͅU#=K�QL�=�T娔3ە*f��s�Un���\fz��  	� :��@���I�7ח�kTky}�M�}�����;DtyUѣ�Qs=�B���= ���=��O��]���   :��Я���"T��
I�2�| nܫ���B{q ��� :K��H�Cv��B��:�������P}�Ȣ��!���Х� �( ���Eq��:#��I��>�|� s��`�9 ���t	w۽�: _<�S��1���>{����� 8 P ��D�=�T$�����TJ3i%�O�� �`y������I}�R�8��e��p8�� �g��='��C��7c���y��  ��Ҋ  ��Dvo��<��TW�z�e���i��7��Os�p��rP1>��a�m{� 8   ��T��BB��QJJQER>��s�z�� �v 9nC �Ps����Ծ�����*���#%�   ��RJ ���wwIaʪ, H� ����Ȼ� uΪ!` �s�@47X �  P>�� T�J�UU
�����RE>}*�6$�� �# �rRI�a�v�n�F� s��%����u��
  �  �y y��@'pT����!C � t7`��"�ѻ@3��T;�#���       PS�J���i� ���2`'�Ф�P       �Ѫ�1R�`      l�(Ē�4�4 d�@ $�$	*R       B�����H�LF"mOQ�41�=L�w����3�}� P�� �>��}�=p��=)z���QE{E�HǏΈ���"���� ���� ���~C���?��_���~�������T��*�+��Q�
��o��A���_?����ҡ�0�~V��'�ExȮ2+���"0����Axʮ2 c &0�c�ʧ\a�"��0 c"��.2��� 2"c 2� ��
� ��ʁ���
0�c
2 c 02�ȁ���
���2c"2�c)�Eq�^0���®0(c*2dGS��ˌ�ˍ0�q�xɌ2�.0c!�8�c0�.0��0�.0ˌ�Í�30ˌ8Ì8�0L�ˌ8Ì2�32�!�0ˌ8ɌL�ˌ�Ì0Ƀ!�0�.0�.0����ˌ��c	��ˌq�xÌ0�.0M��˃�2c.2c.2�L8ˌ�ˌ0��0c.2�0ˌ��Ì�0�.2�0Ï0a�ga�^8�xÌ�ˌ2�/��2�.0�.1�e���0Ɍ38�c��0����C��2��)����&0�1��&d�L`�L`�L`�L`Ƙ1�1�1�1�1�d�d�`�`�`�i�q�q�q�q��<2c&2c&2c0�3�q���ɌÌɌ�����Ɍ�Ì�Ɍ���8�gx���Ɍ�Ì3�0�2c0c&0c2c8���ɌÌɌq�d�8������Ì�ˌ���N0c&0�2c0c&0q���Ì��8Ɍ��8�1�q�1�q��&g1�1�1�1�bd�d�`�`�`�L1�1�1�1�1�1���0c&2c&0c0c2c�d�L`�L`�`�q��	�����1�1�1���d�\a�Ld�a�1��1�1�1�1�x�0���ʦ2� �"�"�*�(�2���� 8�0#�"c �q�2)��� 8¦2)�����3*c*�¦2���c*�Ȏ2��"c
���0`SU� �2)���8¦2#��c#0�0��c
���2����*��0�0���2��c(8¦2)����&2�0��.0�� ���2�� ��aG�"c 8Ȧ0)��c 8ʆ0��� �8��2��c 8�&2)�
c(8��0�* 8¦2�"�"�Ȧ0�� �`LdS� �"��2)��� 8�&0�"Ȧ0)��c
��&0���c"�¦0�ʦ0���c"�ʦ0����*�¦2�
��2 c ��2��c 8��0�0�2��c(��2����
8��Ex�*�c2(c*L ��"p&��1�M~����,������,�i��w���;��Մ�ݖ��W��y���0�v`;������^�yq�U��J��
5i�4�,U�VxV�L���.����4&�9)�	;R�(�G����X^�Wj�b��U��:�ܒ�e!IS���J�^@q�ͣp���`Y�J��ϳ�1��]�a���IR���5�*3n�#���U('" h��p�B�6b&2����S+a��j(m���q�w&�*�G�ǖ�v��(j�ɷGlSk^ޗD�]�U��uf�l�7)�ܽ��Գ+m�tMJ�H+-:�im�S7�����b�ùe�k.����bκ&�_�r\��vSN�da���i̧�=���-AM��Luz�VF\�ۺ�R����V,^i[D���
9R���z�3#�w�k6�eJ��ջ���Z(l���kp'5)�n��!n[�SwE����Ûa\͕��u��y��F���Gl�YWg(ͦs&���V1�[Knк��"��F�]$�@�ca�0F�aE��:6l�a���:�zn�`N�B3�4v�]�lj��^m�`����f�mV�Y��8��mY�(i�ngtm�ְ�bۺ�1umJ�K��NLǖ���J԰B�ݽp�([��e��!wS0�:��եA��c��kt�AVb�f܂)tk��4�Crdj�anj�73M����ɲ1
 +����;�ǻ����h�Y��ܕp;S\жk�v��n�`ݘj����oCI+�k7^�Y����31�d;���	�<u�;m�����&̚���;���p�{��f�e�5#mJ���Wbb���o��niT���/�@s&gT��B�j��L��{C4�I�K#x@���e[�7��Z��� N�Պst4�� e+t���7C+jh+ww�Y�fJQm�+U�qJ���~v�E[x�U$1-��Re�]�+@�b�܆弒0ͺo%lJKv�YYm��Rc8
���u��qs\H�oY�n�"�Х��ѱCL�����`�U��EƐ�R
Y͕�Y�c��ò]����(@����̶H�������E�&�5�o	%���5�dE���0�ln�f�ki��Ԭx�f�I2�m�S�5',�7q^]b�H�+)�hj�E3�^����i��8�Sb��e���P��fb���݅��R�d�Ÿ�
��E^n4�%hmjʡ`�m�R��lz�sjF3mi]m�	Tf=�Mf���*�F��k&m�����(̫�.ȩvFk7[C(͔V�.���
�XnnS��eԓl��fe��2=y�.��
���+���*T�4ߖ�O[�n�Vf�������IC3A�¯4H&��F)Kt:w5�ww�6��A@�J�W�/h����0�<�A��bSFӭشmZ���̢/=�4Ƕ˫�׎!�c��f	��L(]�!;�l����$^aI��W��tQn�v�%�q�zE��Nf,
%�
��M��ͧ.���-�B�Ce���:1���%MId7f�-����k	�6�<�׶�F'q��˻���E*�K��8ܭrב�J��X��[y��+�V֒e�Ԏ^�,���5�]Y�m�B�FQgs&ا���J�A IH�Gt��N��Rۂ�.bM��å�]��Т�IY��M9�2ͽ�Ǆ�L�m�J�y��J�*M#su�t���Y �!�������F��=���*���s ����a�Mn���n�&�Ǻqe��f�qek�뼺f��)�x�6c%�����[J��336�(�E9c,�]���(i�͗�71] �Gf��i
�Q%+�[����[v��	�a­�+�T>��N���f�ZsW�W�Jŋ���k��U�v2��{J�A�o+k%���W��ڻ�H�G6ĽۛF]Kt���RU���`��fKg2��~�ja|v+5����h��Z�b�Pd:2�l��v�iܼE�N�"3@�V�e0��4�ލ��B�c����ES��eݲU!xX;�i�Z�ٺ�)����n��YQ1����ۘ�j��30�SE�dm�7uz^�SVZ��[��
���h�DE�±��ÓTJ���� ��2�l֧ �+h�M�f�GNK���x��+	���r^r�7�,��*����w`�z6��<�,h��zƉ�	owc�e���Q���n�3��Z��%�uk����h=`CY�����cK�"3\7@��HVL�Xm0j���ͫ��ҫ������" L�w����;ئ��;��Ё 2�;� �܊�^r͈͂
ů٩V]�֘9���V�� H�M\Mŷ��h����{�l��u�-��A^-Ƭ �9�����!e�t�+]�{y%٭�0��7�m��&�!�(�'*��l��*-���ڬw{Zԭ� ���U�srh�����t/5�@b��Dז��S�(�P[b�,�64��g#� 0SQVT��c hւS�t���
Ɍ�o�pm�7�[�8�;+F�*�	-�����%n�X31��C �9�N��eІ�)�MD�x���2�Y&��B�m�OU��)���4h��[�2��%�',7��U����l2�)EK��nQ�2B*K[w���z�r��'D�{�
7���@,{�+ U��4��:��wwGr��E?XS�KXX�]\�(J)-�XQ*an���u+2',ՉC3hR��{��@�@+5f
�LB��kAO.��F��e�x��Æ�����Ӣ��Y��IFl���S��g-���k��W��=��oM!l�wX����CR���oF�Y7��R2]n���<�)�%<W��wT;�L�,�w��/CړD�W��Զ
�R:Afa���]�+s	�6�hl��h�b��ks�蓁�e�0^l�W�s�:T$��8�R�7�\ͬ�[��k5���у�&]n�K��ݕ��7�Q�#�vkSЅemɑ��w'��Hդ�Rb!N���
�@�[yz����#��n��f���ĢӨfn�଱�n��V���5�f@�᧷ Ǧm;��$VTx���x�������V�%��TLc���WL���R���^�%#jHpf������3��������Zզ�{xN^���aF�o�Z�t�.�e�C^8�z�iZekܽ�
�&��v�RĄ�YY��-ʼ{�k��&k ��h��%{W2��vj��6-Dd��՗�^ҵj�{�1�aD��Ŝ�U���pu��m�`hW���lXݵ�fl�Wot�����AN�K��Ca��T6�QCMX3q�{J�ǹN3�o2�%b���IRZE����{��b햴DT#C��I˕��>5mp��4�Bs2��v6m	L@3���:��i^;����@wX�ŬѰ�6�Z�	
�9�M��-��6��f@�KS���DAy�%e1`��u�m���О�0:�#��-mM���*nfR;�x��-�ѱU�Z�͹#��4�6�i�q���^:�(U�n�9�R]"箘�̣��d� j�Pi<�E�X�`���;w{6�3�U��pG���V����U�"ݧ��e����"��uY���+�V��å���d  �:jn�{�,��{2�b�6�L%�o�nȥ�X�X�����除-5#噮��c2�q���;����.�ܐ�n�˨���t��)Mw��˼˄�g.��VV�+<��.�(�<�������p;����F�H�ҵ>��ٴ��qִ�UaYR^��w�wy�N�wi�n�Yś�u�Z��WC��L����Zкm��� Qҩy���"!���Nl��F�+p��a�胗rP����V"�����E�WY7Kj��u�6��{Y�Kh��$����t�Ű'�/Nё ��(����&БČݺ1[װ",չ�(#`z��3`��,�rn24���B���&1��n��T܉��lU��r<�MB�]
:o5�NX
�jwx�O^�*�̻a�K���;g2�c�M��q�����7zrǵ������[GsX7�-��8]mS�-���IW&^
B�y�H$�3]Kq���K&�hV˖�V�[��8�u������'�̙�Z*lr����+�"7P�I�W��4����]k$�er\��"Fe��	�Kl�����^Ңm��u����l�Uɖv��e��B���E�V7��G���j�`̕�F�,��G
W��K���
�Ěr���fMV��t�4v���5)�劍Cai�Y�bd�M:���"Z�FQx�<d�@P5b�B���Bn���Yvw�VS�bn��*b��6����;Q[ȶ�������׵�̏nCGk�.���F��T�[ ��Y
�L��جm� �T���&кץ+N�ڋRJ�����X
�����0	�E�[�����2��0%�E]WM)WjYT�:ܒ��pl�u0k[0�i&Duz����fIN�qY�.����.Z)kxC�W3+�.�P��x�X�!�l�{r�Wg&����M%��������F�9��:^F��*Б��vEK�IJ1f�vަKW���w���ƪ&�P �z�e�6�Z��56�+wV]��N����J��+,]��R7��+:r��aHK4�0�ѷv#y[�/�J�V<v*������a��6��^��s.��jQ���x�۵�Z0eU�J�n�f]�Ńy��H��A%I7�Xp�V�e�x@��6��/m; K�kApb�sH�O�w��N�F!.ʡW�M� C�Z��AALp�v�t&_��Q��l;�P[B�/�D��I Nju0��b/�VT�mͼюA�o,L��3aY�[�Aj�k	�,�Tz�����8�0l�l/`��gL˿G+d������ɬ��n��B*�r�\X��pې[.�~&���t�T\���%�P;���0lL�A��J�4d+#5�.���U��T �՛~�L+n�J�7)f�d����6�6Ɓ{B��u�
��ŏ$r��g���Tt�k9��[&�!�83j���Żp�f��`ɌJ�M%Z�t3A�r�ߕ��Ct�a�b�Ije^ޭ���e�e��[���n�!Xv�w�VV��^T�voR�
��
�P���f$(^v)�J+�Y�	�c�����j:lI.�5�<#pP��ùv�"�r��'1ݭ��l��L�E��p��(\Qn�7@��t�&x��7�f�<�-�pm�����Mi�m��
�u��2���Ԗ8N�s�h���8��U�m��e�26���X��̭���:"�6�n��֊X��[Ͱ��:�5�H�m�/ol-�yv�����jr苚�R�-8o.����}L��^]]҇��x��Be���y�v��ӘJkP3��R�w6��:D5ut�HV�j��@�Ѹ�g�Sےy���xv����N�<�c0SY�5��,љ�u���`�J�n�V�n�츨kJ��iU�i�շVl��E���&��Z���k�`;-�X׎�z�c&X>GR�n��0���]0*y��)j��N�r�6��
�n^��r�!�TC��h��/F�3%6[�(������p��76���f�WH�I�csٹ�wa�p��*���l���Z�]6�nj+-��/@[4�դ�ɵj�	����K�&e����Y��¡��N�f���Y	]�jʰ���6�B0����2�n�֕6�J̴��C)7H�W~+jyW���|3&0av�R�'�7Ik7ؓ�}g= ի�WA&�[��Ù�.��ȥnD�d�f�h��ʽ+�l ��e�Kw3M^AxdML�]�L����Vw�a�*lc.�[����md8#�N9(0Ѩ4R$�E�������D�ԖF���J��s��v��:�%Ė`�՛t��Ǜ�o2�ʀU<�W hKUz�`J���Q�%a�m��o˶&<�W�]�~Ӡ1���-9�6�Ѣf��������L���˳���+-ے=�3u� 77r=��Y�]�a�F��M8F����Xw��+�{��y�܅�Sy�on�����Ë�7g�L�$�zw���IjZ�хv����,Q
ao;򛧕�g2��+����6���]��D��Y$�O�d�D6I��N��!�d)Z�	a5�IJ����U��q�N�T�d�����)����Z�7�
��8(3l�;�b�W�~���/��� KQD3�S�-�,�2�l�VT���w.��B�]���g��/hop	"h�U��R�VD�N�2��$f���^�������%�d�-�g�0�N쿉E��8]���6o�2�p�1�C�3&/��n~����~�!t%dÄ�p�M�t/���w��o�3xp��4�YA��LdÄ����f�Y��Z�Uj�lJ���;�I$�nZ�2�S��\K�#jlhc	�D*�T�d��EN��	$a�r�Y7B�M��6ID�Y�1�g�]�Q|f�f�R'G�P�I���3�ܔ�av~�0�s%e}�Q�2�Gz_��3bZ��Au�� �>��UJac�i%�-�����b��C��Հ�ZM��K,��)�Ì�[@�,�Y*�4�$��C�]���$T�a�w�N���=�����(]~�p�G�Q/����`����2��L7e�t�I,�{C��hV��62�js��6�d�8rɆ��7�~�E5��=���t��3��KF�D�J?�DbY	��Yp�t��tﰞ�]�� �!��л$��vH�g�>�l���L6
�̢UZ�H�I"�lŷ��u��0��֢���i�:��ũ^�u��"��(�X�'��I��~��N�K��B�����8ϏĤ�o�ɿ�K�Un���)5��0�$ܘ���RD>��P�B�^��D�Yz{	FYl�,�d�(�/��x�-��x�����Ÿw�a��c됆Q*���p��{t������l�����o����p�M����D�`9� ��R"P���@y��J�H"�䂍 �!�(�
�)H"��+�T�҅
J�P% �P���T9#BP�%y 
�P9H+�P�@"�rQ� � 9 4
J�(� PO% y
�H�@�R�J�P -4�%ЈҡH�
RBrS����@
#H���%�H��J�J��H�P��ryR*�y*4(R��!NB4��!@�9 ��<q�~e��B���e:���}}�3J�5���@�J�^U!/�6�9߁vD;����Op`��͡�!<�7!9�t�t��!��y�@���rM���0a�vP��;�ň�O^8 �d���ϓ\x��z��x��Y�,�|�$�=��=Iꛜ�܉��@�����-��|��B�<A�}Ȟd�)��u@z�p��EU�~��}�EDC}lo���������w��~�����g�>�Ә#�+� 2f�#�]Z���MWC0姃1�,!��;X�[s����ۖ�+:.��Z�����nL̳��X�傛.��c��Wl�n�
][d�뫺rW���"wj�M��k/�fE"*�e��^uҽ�V(`CP��^��ش�S-Q}e,1��=kmw�)�Ĳq�+���p�{��<B�tR�n�$lS�P����6n��j�bĂya��9]��<���r��Z��GS�m��Gw�V�"�Lj�|�;��{�ˬF�8jv�kl�y�/�VӴȋr�u��#O��A��7��t�Y�7}�m3�J���Nu٤omXhr������H��f�op��Z�k7t��s蓾�lv�wf�p�|�f��6b��*)�Z�ݸU��Zu���r]��В�[�N��v��������ʘ+���S�Z�2�I����4�qj�.��ͬ�Gm�y�W�:^	�ܾefZ���x�Sλ���E=�[��k��N%ٍwp�]�6�n�Fv��N`K!s���x�ٴ��7�-Y}�|���X���d�-����������2��s���a�r�w�k�hE�Z�H��+\;r��Y�ùZ�������[81����m>��^�=u�s�;|=�����}��n���뮺��:�:�u�]u�_L뮺�����}8�}>�N:뮺�ۣ��뮽:�OO����_/N�뮾u�]zu�^:뮺믗G]u㮺뮺�u�]u�_.���]u�]u��u�]u׷]u�G]u�ˮ�u�]u�^�u�u�]|:뮺�뮺㮺뮽��u�]u�˭�S$�r�t���v|lAA�/j�V34�.J诖h 8BV�`w݇a�}�����%��3!yF��-�f�s�(��F��"ѱ�$s/� ���fu<�Ҭ�=ɩ��:��9ƴ���J��M��,mN(�aU�f�޷��gr���^c�@�5[{�{u���ʺ�z�:`�-up᩻��&
rE��ʡL˕�2�����\��c�-�{q�m�u�s���M�m��	��!Ϻ�6�4�V/�G
���(���oI��­)�܎���"6�������n�q�	�M���v�l�m�Y�����y`�C{B��C��&�8Yz;uJ��胼s+�I��v{��F�ByGw7�&�{��vS[#7��uvP�S�@L���ǂa8�l]U�C�d���RoX�Uw`�S)n`g���k<�f�t([�ۖ��X
"�i��������Ő�n�T�P��UƱ�^&���뻴u'[��m�9]5��ռ�Z�δ4ۣ��S6������!'��8��y��u��y�̼kr�*�C�c+,Mj���=�W���$��ܩ��)a;�fU<罤�M�Ӛ"���h��ݷ״jp�m?^ع�i��+�m�Ѩo2A�V�JkD�FWf���
t�Gb�`�c���oo�^�u�]u㮺뮺��u�]|:뮺��뮺�}>���O����^�N����Y�]u�_.�����|:��u�]u׷]u�]u�]zu�]|:뮸뮺�n���]u�]u��뮺뮺�u�q�]u�^�}::뮺뮎�뮺뮾�g]u�]u�ˮ�u�]u�^�u�u�]|:뮺��Vo�[�]x]PJr��x�$:«T`�-[�m�tr#���Β�1�6�
ä�g���pw��ٺ��'�+}:��:�,=ܳ�\r�hڔC��򳏻6p��{j�R�ث�f�Ð^MCn�m������k�O�A19��NBa��7{v�9I��à,Y�R�,>�+/�h��`�Qv�TؗY�
̶�kp�bJ�d�ɪ�N��W�����uˏ-���y�F�x��g^�W:��M��j�$��ѵ%fZ���w:��9o��:e��ҠE�hWv��(��:�VC.�Պ��XV,E���\:�T����	̽��(�<eH�e���w��CV����O�qQ�.����f��}}�^�rm٭�׃(+�@�f�;���ؒrǽ\v8���u/ޣ  �qEҕ����kyq�N��P��[A�Tn��Fj��N�4f��k�d	��6�Ձ��� ��L��y�VgQ�=���ӋMU��e�	A�h�3{Ng-i�nT��:�i�8��@׸9Q�up����6�}+7%��f�]ׂ���8��Zҭi �s���$ge ��p�2X�U��V1T'*�8j{��b��Ogt��������k���3-C*�[�XT��2Y�)�F����Ԯ�!��m^u�������y�}��w���a�]u�î��N��뮺�ۮ�㮺뎺�}>��C���}:뮾]u㮺뎺뮾�{{��ޟ/�]g]u�]u�ӣ��뮺���^:뮺�n�뎺뮾u�]zu�]u�뮺�Ӯ�믇]u�^�|:뮺�뮺㮺뮽��:뮺뮾�u�]u�]u��]u�^�{=ޞ�/X�gr��ʫY�a������@��]֑�3�^mK�HFk'�{��c��ow�����Ly���%\�f0�N�
+GL�m���=��T����.�삘;w��vЛ�r�l͚,͕�z)���v��X�Xu=�R����h����K�(��:J޻���\F��K3��w[����8S���8v��e�8#�yݓ����JS����ޚ�Ku��!#�۳���Zvm���׮u�z*����P��g^k�v�ǡi��z-4�.�����w��S�f����2fUi閲��c�çzs7���-P�� 'tr�cV�c�~r��]���wK\ͫ�ެV�ى��j���e��+�D�֌u�/m.�Mv�5��c�2-�n��	0�u�^9�uԴn���Hcǈ·��^e_es����G^8�v�r�t�B���6�SҒ���h�D��2�U�,,���P��R��E��M����X�������`�v�R�`n��ճ]�L���lN�#�u):v��{����+��+ښ����v�=o����w 4��Zk�5�G啴�v�U+Œ���toh˓sz+n���q�ޗ���_W�̀���AH���M�c~̲��;�W�oE���{���C@�4$p�82��i����p���ݵ]�*��2������GT"Y���;sM^��Պy0�4��������"��d���n@���;ڣ9%]���"�6vvZ{��9t\z��Jf������s6��.�8ݫ�͚"�����չ�frU�d���厇Z;��雋��9��=�UF-ݦrC�z�ۺ��G{@�9�xzUz������N��4Q�i,���e��	�V���f!�P���j���$��~�0+	,���oo@��ٛ�=�V�m3,{k)T�+Y����	�p�>W�A�ޥ�u�1i	���^�W\�	�A��E{1�	��[Y6��g>'�	rc������
w�n�#�7��"��׶+޺�mo:}���Tq��ߠ�o7*����sR��2�7����'�����Z�b� �N�ٸ,ᵅ���P}�l�cު�;M��l$VY���툪�� P�SOD\�AQ������oS]��`�^�j��i�E���'��4�ΐ��c��+�3��-��>��[t��{����d>��׹�S�=��;�r��0��
�W
�p�]6fR��嵧r�&���3m{nA�:��8q�]t\{J�5�@�f�,:����Z����;J��w�5�C�d!��k��귟��ܐ��7ho0.�a�׃]���]�Ss*���X�~�6��N8`ə��8/z;Jzfy]Q�����u�1��h�7�.�Aunӷ����Pz����z��ָ���7�f$%kq����2��\�:�]Ö4c��:��v�:u��J��ά}�}��%+��״S��ޝ�\�n�tCEcF��7���O{ [u�2�ͬ�.`������ާ�����Ř��ܫ}�l�ed��:���(�Vv����R��ap�a��U� ��}��K��d�sr >�Õ6�pF��#�h�����zz��j�9[v�j�b ��b�˿y$Ջ.���u����Yi����!�c#�kͫ�{�$!��S�.�-(:<++*�u���e/0��4M��n^���7L���&z�㸥��oqV:�w��O��y��.a!�x9Bժ)|�˫��[J��׃��}KŬy�I��U5���^�w�b���x�1ł���T�k8�=�Y�UZ8�S�aU��Wr�-�K��-\M�Y#���mʔ�b�;.�b#xv�ګF&-uI�o�W]>m�楽W�i��T;�@�����ȭ��+)�h�7�s�V���nT[ˮ�R��۫@�K���v���nRU�u*wNKk?&���*6��l��jʳ���K�1��ٖ�a��̮�Zfۛ�/(�����-E�g�z��:1�IP����;�wO�_fU�v�ղ����[X�n���,��3]� �07��R�vz�ιj�{�tr��f��:�"T4yG��5Y���Y��y����S��M�:���'�Mwqޣ�6`}�Y(���<��k����2��`��h=%�zoL+�`&�X��h��{7��`&�d�H��v�5ya0^�e�^�8)�U\s�z�[���{��q3���^�+7Iίx�Qק�����_�VY�mwu���L�{W%��C��p���u�У�e��;7�gb �9�xoI���E3���wQS�{���8,Fw"e�Zz	���)���ʻ�+6T�6�L��r���q8%�Ș.�Z唴\��ܮ�ndX��Փ����1W,뮺�7%7.�
�ǆi�z��BQ�!���ʳ��7{��+8�q'%��z�Ss�r�z�W\��=���sC�����Lz��̚��yG�����8N�c�龧y��\���ia��-:ۣ~�C\����̜��{��7}���ni�����|0����[Z�����Ík��z�;���]JL���i�n���
Gv��5��)g�J��J�����;W��/�b8�5�l��x��bv(u]E�䮅�!t�aWMY�=�4��N�"eе���;L�0���yK�t�W˦�y���C=��x:7��2�F������eb��ڽʢT�\����d"k	S���{[�غܷ(�h��Z3)��LŚ)��f+����Vv̳ۏ�.�[�Z�"��5�w|�ⷊX��U�X~WWO4o1���f��4�;x��{����'y��w7�O���us�.�^�< cS7�X�zdk4l@�*G�Sٕ������*;D��Y��������&45��e�̨���K�j��{`��Hn>���Z,G嫒Ac�i�|��l���Y���H#�5^�3*ш�����*"��f����Vڴw�˧�Ǯ��>�7+�Vk�'��;�H��CZ����"���Pn�61�*�ƻ��K+�����mU�+���,����t$E�rv�d9���V���6�] �-.vE��}�UwV�gl���
��?BL����qc]����޻�O����NA�Q�vj��Yrsyg$3�V�=SuvHv��C�}t�u$W[�����}�}*$�����Ğ+C��z��}Њ�:
��s$�(^n�.e<4��%�t�!�y����l�s��n��]�
FV�o���(�i.��θW&sX�(=��hY2���M�Zm��zo�VmX���E�W~�讬V���ŗ.N�Z�Z:�Qx�ow:�
g0s����c�wD�/�j"��h�Cv��L�::�<�j�����MBĨ3G*�<��,fU�ݒ�d͸.V�g2���� ��]Emje�FSU����Z�4�o˷�@�f��i�|�ve���F��{wi��h ��s�MdZ
cwW��IU�.nL^{m�����zul�[��x�r7c)���Y(u[6�9��^Y�%_i�;����s��� ��66�N��cV��z@ Ou3l�������u�[��N���qq�ȼ(v���s�t���P`�S[�RV�`�@5��ίW`�ctcPW�սy��I,��^�fh������o盷R�伎�ݮ�%C�U?9��\�*��.ue{9O���\oz�^���mM4^.��D�Z9��AײŞâ�l݋��;R=�D�]�Y�/ 4d�%�D8o:��v�f��.���z�"�B)��6�#2���u�����N����g:��3%gU��]�ݺ�%5]A�x��u��:��Y���x�9�{���벆P���/P�z!��<i����s)VB�N�� SSOk��<9]����F��'uDe�`�f�d��0��ڮV����*V\�e�0 ���)�ސb����t��=��Y��rK:nU�r��*v���^���u(%"-�f�ݱo�5T�lg���X��U����DQ(��>��"��� Ch�n�K�:z^�#-n�}1T�"��i�ԍ�c�J�]��ֺ�W�㹙<�|kHz^M8�98�t:���ye�άε-݆�����̵��Ɩ2�봭I�::}�=4���FM�"�����Kk��� ��]!�ŗڟE��h�:�t;|��楧���4 b����u�G�>F�*:�(�n���]����{n3c;]1�x��"�l�M���ѻ�.�{�.gv����j�6^�k3e�B	o��nOvVe蔩�畼SXq�陠�QPnl[ws�5�F�%�}b�w�

]Ҧn���\�^<�����	�M�;Xu��u��͗��f=���oz94=�β�9k���o"AL�Z�r��(*�b��ut���ү솥v�Vf����P�s8K���4{��U����6�|��LIC5���<��]�|8��#��)SZ��4a��uo;[�:,�Y�܇,}�V��k�h�*��Cq�P���j�J���V�v�+�����J�ŝA�Ҹ���0κ��3���/VN��Y6�U���mE]�c.��xu-郞����)��e+kl���z�{���o�,���n����^��)sp�Jj����������=�x{¿xW����_��w�W�U_��_���9�x���+�]�DF�k��E:Z�K��Ѵ`�����uf��2��f��c΄|�[?qͅ�	W�r.��mCq[�4?��o���Ś�E������M�`�0��	�����U`�_��o-��,���`�o�y!rZy���ـ�ڍ�1
M|�x����f�<	�i<s���1�{3��<�U�� xM��i.m.iC ��KagK�-MUa	F��k.�Irz�NJ�J��5YT*�ɝ�-�M(��A���܁5�6�e�����ԊPt.�����V'а3qk�3�:��H8�u���ٔk�ḛ�M�4�u�X9��f	�l\��ƨ�Ѐ�嚭�RJS6�a����I���ڒ�YE����sڒ�i�Kb�.�ĥ �&ٝn��ű�Kh��WU��E��'jX,��p�n�P�-	kG$�k,�h�䫶vU�g@SJӓ0�"Dq��δ����y�� b%����9 �Қ�]b��� Q9�l$�4\%j](`��2��f[SV�.�*��JGTƲ�u�4N��Q�l4�e�![�ó��4�y{,�U��j��X�i���1.��� �cp�l���(�m	s4���� &����Hj[�
��̶�f408��b�X˭��XrjK��B���gR���ц��mٗXm�`$f�ڎ���m�bW@�Z��^���sqDʹ�-�m�*�ݠ��c��)�u �`i�\�X�Miua��We���L1���D���\(٬�ѵ
pu�U�$�v�R�y�8�f�+��b��mZvMJ�H�[��G������L"�vɳ5��5�b�%��	[�����Ś�n�ahF\m6�˔����,xU�v"Yl5AT�Y��X(�<P���[m�M�4966V�-��E�;0qz�����^ i�.���GAѰ����3���X��WL�+��f�3c���c)���glűE0�ٴoL���YPc�1�Z�#u&6��	���T��SGChP�����XM��5�R�,�k�Qq��ZB;��.�̹6�u��R�fj 2�E춐��ګ��M\�f9�fMtהiY�6�!LX���8ɝZ9�و��X�j��j	M�2�L0[����L9%A��ѽ�.լ�i��Z�H�JY*�X�I��턯X�ٚ+��k�6.�:9���(VhJv��,�h��\�	���A\k[cnj���hR���6�(�n�h]2�-��6Y�C�2���*���-F+wlg\搻&�1̇m5�\[Na�%cql	�͜*`ri���M��]��;S�*W��w$.���i��#�V�f0�v�l��&�ca�m��JX�W������)��37[�\:��a�Gvt���LIf�[-cd�S��j^H�8lme��X��Э����Ĳ��]sHkQ�M���ݡ��l)]Z�c� �LP,4���خ�V�@%	������4�R�j�]��KR�u�c]�Dx	1�Sb�j�-�9�9�iCL�8[\��Z:!uh)Mn�1M�6هD(ە�@qR9%�x0��؆lԭ�S���l���e�:�a@a%ׇF��D��ce�mf��"b����
�5n5V��e��ٰ�
5n(Bkf4�d�`Q�L�V�b�T�M7'1a�F���(�7\�)���52�rv��aE�6�\g1��B3X�L����{3%6U���l�1�ZEՊY��4��-.���k�M(hmt#���a�1�jh�ٵ��gK�FL�kر��m�1��30��mh�����%ÚTI[�n"�[\Lwi��4��wh��-�5Un�	��� -�qL�U�U�p��n�CL�`�"�hj@�lP�h�E+�.wQu�J\ۇJ"a�qn�Y��-툄�lp漖潹*,R��5$3R��b$qmU�a
@�V]Q�g5�6�ة6�h�P;l]�b)�Z�B[MH��'n�u�:�h2Sh1�T�)���Pe�b�!��E&�˘b]kF�Ka�)h���+��3IF��W.]1�GZ���SLی��T��yh�3K��J��,����E]� ��ڪ��v��i�33ZmL�-6�fB
Ѱ��ȤSgk6#h+1m�ن��[�l����X޹��pU�M�ua[����]ƙ��������Ձ�3�I���1�BSF�c�71�YUÍm=h'`�"��ڸ��.����a��k��6�b�a-V⁚��b=��N��Jb�2T�B�Һ�l������.�P�c.�cK�*���	4�%J���Bf4tم�u$ �s�f�M�[v�iL�eGs�S�Cl���*iEf�1cRb�:�q#G�673HT�k�3<�^n��^F�Vv�BulD]v,��a	@��^+�K�B#�(\�1�]!n�JT��m�AjE�6H	Y���bX�sR�B���-s6l�ȁTv�n]5�[�C0ȅ�T�]5�+I���1Fk��M�`�l�Lq��!���B��v.f���h�.��܌͈�ɘ�M[1v�{Z4V�AZ�AViVX���4���J�&tIMu�&6%�b�6U��%]f���(��.da6Mmtc47 ĩ�u] 4�hI��[��[�;bl	L`&3��en��mAتUs�b]1��5��bPe��6Ebl�!&b�n��p2ی�y����Fh�M���j�rZE��2����"[Sj�˻\K���X�+�&n�:m�cZR�k%�M����:�C\�u��!e�$��[0�\��1̮�җ�q�2�巰��لIv�Kylɥ�K�Խ��Fݵ-�+4���cYu��Z�ƀ2�8���$B݇���"g8�Y�/�4a2�e�f՚�����"ٛim;A#��u�[�&�]�lqjUBX8�<dw��M,جZҒ�fc�y���m�t�́�l��3�%ctq��ŨF�CMuRٓT��HٓY�Vl�!/j�)]70�i�lҜm�Lq��nf��nII��è�r�U]ڸ&c 볫J��(Ƒ6����]Ga\��5�dYc�WU�5�Ev�#�����ŀ����0j�n�3-����5�r�����I:�a����k���gmN,�ilX����GgEj���[���e���e�R����F�)��\\�1&��2֘�4�t��,�9�ԋb%�dm�c�GB�����4Ýj�F,za����r�ل5�#ne(Я9&�,�Mظ���;)��6�dD���i�ņڈݝ����lZ�$�tלXc�v�ɕ�@.���-bh=u��%e��b��.��m�(��0`�ŭ�@�̪i�+S"V�n���U�:�l�,��a
�ٷF!LJ�,s4�{#�����4��tf7B�[hB 2�15��.�25[��dqWsR�!a��
�bŤ�`A���4cV���5� ̬��Yr�kc6W\���Yfh[e���@6t�\�	�9`��Q�کl���YU��Qa]3�.-�7C^��.�V��H��%�t�s1�L���2�+���]Z�ˊ���R,�Y�4��0p����j�l1R1�沥D��m h[�4���UsEփi4F1�IU,6�b�-��v���Z�]�8�qK���9���U&�^�c^�i*���a���Z^m��f� �)Rh�Lm��e3�ta�2����؊`�%�\[,7��73G��vѨX�m�Rb�YtKWLlfSV�3uH�n�Ylh��#(�ajF���BQ T�R��kY��#���:Y���0�l�+L��vB��Z*<�z['i��)s�ٳ�EmH�ٺ����0ۈB�,�X@�a�i4��p�%&.t���q)q�l�h\��+4 HV��̴֠��fYe`�mrĹN�؄a�u��E)����s1e�9�	���d��Ҵ�.3��5z�v����dŔˡԆ1j�#U5֚�P��L��s�J#�\�)n�nP6���s��s��ͨ�e֗F���@jɰ�������M4��xصfl@�0��$��n� �yҗv�a,m\̋����Ʈv�U#��]��-�7h���2�2A,�dm
��
��YvŁ��.�7.[d��	sp͉e"]X��f���-w8���lfЊ��p�e�eр���4�&�i���:�Q�2�5.U��ٮK��\]��mQnf�Z�W@P���RY��Fc2Ja6�a��@4jG�ݵ��t՗j^,kb6�1p�u�eL�4XY����.��B٥��Z���H�BTk��K�,�:Př��ѷ4��]5խ[��f��f�0i��#^J�h�fcWv#α���(g��0q���ɜ3$`��ݰ���XnG��T,r�-�f�3YWCMjJ@��kD�����5�ب�ŶR�-�j�Y����B�Ɓ�,i��T�����c�G"L�Vc��i��m��F�Vl���3S$&�S�'Y�Äé���&a��nԃr�l�h��Y�[��%�ɩ��GU�E�Id`j�ɣ��l��n��l�!��`��ٵ�5ݜu�a�*̶Vj��K[F-t�i2���PsIfRڗZ�&u/0q��ޏ4,�0ɮ�qsl��|	w��h�3 ��)��Gm�mE@%v���*�	�,���e��4H���Fq}U��)�Gm���%۷%�`f���_~y��<�bDf�x��6��]K���i��`b&��-n;����*a9�pʳR��P�XJ\�M-��`,��\���Q*�3B�y�kЖP��h�ѽ��e	�M�����ZZ�R��k����.̳:�
6�u
WhBQ�14���ʖ���ݣ�.F���K΢�Q�V<�M�l]In�\�����sS1K�0��,m���3��K�
j�qj�-&��*�3���B�P�X$�9�ǖ���8ئ2[�ѹ[����)��,4�(a����	nu�GB�0�u�۷켵PQ=����+�p�TC2�R���7��&��9q��}:�3��z{}>�f͛6lӊ�*<�DE�Z�1��Ah�Z�r���fAc.0r��Ya���Y�'	���{=�6lٳ7�����F���*�6%���ҩ-2���1IR��Jf�O'���Y�g��y<�O�͛6l�p�JԽY+�R�"�h*�ڔQ1�`�A���!�:����Bq`�*΅�5{�`�am�J.ff\B`�/8�b�$N@�!��˓	PIk$p�L�f8d�@-��p�&޲���%Խ:�I�r��ҵ���Y[8#
�TRČ�5�h[\h�akcA1�\�X�"ʙKQ�\rLL�fDs3��2ZF��
a�Ƈ�	5��-�d	<z1$�K�;^�����!"H��Kx����X�rB�y��X��48�J0���!:�%�� ��ebl[�}�l�i��kK��0�9�m̧tw&Kmm2�ۂ{(|ιOE�K�w����ź-��Z�0x�z5�F�<(o�-����B��!���m���ZkQB��\0�L�틣
��\�Htl�,f5���~ljR���m8��Ƀ�bal��b�NZ*��V(�ZYKe�www�ޭZ9�CM� ��J��>j�%�D�AII�����BE�7��k<�X��4Ȼ)�e��赘��BiX;@�xvo2��SR�u�mYU%�ob�lu�B��,�4s�@���x�ٛn��l���N x�عL�h�ms	���FR�&݋P�Z�XL�[������!�H4���ᮎʑ1�##��EvJ:�[��&#�ڹ6�j���1�10ڲ�y|%�S��6���LV��,\��\�m"�aˍj���H��Pꘕ�������`��bL[�U�JM6�A�ݢ�����n�!^�ؚ��К-�[M� ��f�DH�\j���en6��k�B�nK�[ƣ�@�#�Mb՗mդ[5�7m*EaP�4�j��۰��MSR6�f��	�/lݸZ�56qc\=Mm�M93���Pu�����]��3JXg���VY�C"�bW;6�Lű���E��i�h��S\�-W3-�],c���BP֍3��Ͷ�\xy��m�Z�Q������^�-Er7b�[�i�l�LQAl
2�[�\�P6B�@j�S8�����9����5�5kr�"V�g8�.��h\� �tz�XJ8q�iv�L�@���g�nm�հ��Y���muf�5��������8t��F\A�fnƉ�&+4ڐ���V��D�ҋ-����Y���5�^2ee��K��#.���0:j�̌�u��۰�ƍԢB���%^��l�R�n���y����+�7l�Ѹ%�%�3ISfi5�C;Z�	����Q�õ�Ry㫯h�T��bhK�k�i���mD���]&���J�Z�2�q)2�h��.̽ukDYP����kۦ�V�йh�\��vb�d�t���ʔ�%�m��e�]Tƕ�m�X�	x��ŀ !�m���-�.��
A�3�Lڕ�&��b6f%�BY�eбښ�QZ�b�a���Q���*f}wt󻻹e�_:[-���al�R���H�� VE��liK^���U��ҥ^m�J!,b�km��֡%D���эl �D�����)+ac�m�ڱ��%%j��)(R�YB� 4�A�b,j�ʭ# �V�m��Ic*ŭc ��K�j�����@H�`�`)"<*D�� ���
iL%!1lK��$�V�л�mQi�n���*���]28�y"E�8pbk4K��,�S�1���I����kRE�:p��3'n��*���SDЀ�,�����I#���Dx䧨��~���R�����t�l++Ȁ	&_[`"	5��R�|j� �+n"�x
����/�츏Γi�����:$?�r�� ��>�$��h�[p�¾W�W�/�J#�i��.�Ƣ]�������AM~�)��ڸ��ײ ��a4�*����0@���!6�ᕗ	X�-����`�SX*�.�2�8�6�ĦB���}Z_R@6�IC�kߪǀ>_/(�7m��]��N��G���������7E�;��r~Q_jW��efI��@��^�@�b�Hf�l?v��/��-�ݎN�xGT��i�ŭ���𸄥������GF�b/�֕�*�����ZA����A9��O���ho:�������$]��Eف��ۦ��0D�w���ӵ2m��	�I��cĿ��ݶpJ�pTz��zd�.��}i���.��K�|�Ȫ(oڟ���;���ZL��
����t�L�h�~���������9���dT�4�$oq��O��DEنA˽��y6(�**�e�m�A��H�;kX͘�l�2ٙE13�1)�R�B��ϖ{��r� S�:bm�$��^"9�i�S|k1�n�B���?���#�$i�r�VP����*�h�]��;�xg���G�"nK�߲n�V=�5	m3�IӦ���C�Ɂ@y���%_�w>T����&͡�]k���P�n�]���7�o7/���Mf���_M1L�ڷwp��;}�Ep�W;|�U?^P�W�����P N�1�}󻫘�x���,�S�w�oˢ���¦4�
N��A#]�T���lu7�D��gwX>�4�&.��<>�����֎n��{�,X�������s�Nb"e��s>���D�ŉs���-��D�Ҧ���s��ʛ3R�cf�h$XX�[a),��~���7r�Ӯ���w��
����qAEk_|lN�x{�_<�Y@Pɷy1��F��H�.�J�_�-�7�����oX'љ$�۫��̟V��o�|��?x3[�� ���m2.���ǒ32F�B^sL�Yd��ׯ���9~��\N|l
�G�A:%�mQn���l׹6��j��s�1�u�I�v�AͶ*�*��L�|܆����j�>��#3_^�`El__��ڶ]c� �?L/��țY��a�2�48-��c+l���� �mE;���遟_��Ux�F�3�X��FṂ N�Dq��H$�j�y;�e5�^�x�>�}4�k%�٥��h&Ҷ�,-�̀/��ݚ,t���E� ݀� �Rb�y߅Vʽ�"�}��Ͷr��Xɪ��7v2E�@�U�ϨD�l�mwwr�'*��3�-Z�[L1���ݫٍ�D2�A��s��*�k���w`�����&�F�wBP�~�~ V}����^5uy�84�v�A���l�H�h�L����rj��ۊ2� }J*�JwG�Տ�`�Y�T�(ӳt}h� ��4��a�ɀ �e؃W�1���Y�J�j"z��w"!���L�0V�K�0�K����iV4��i����N۽�w��}j���ܟ�j�ѾP�t�}>f��^�tc��*�zǫ����8h�I	2�`.]��'P�ņso9��{\8H$]0s�ك[غh�.Q��f�{n3�nj���SBk-�X�!�a�A+]r�1��5Pv�n9� �b�$�Δ&6��~y<�Xx�Aac\�rd�m:�.�M3��:�Jյ�Eu`�kmWK0VL���."\�ݳ�-�h��b\���wn(T��xŘff-�M�z�]�g�0��`��Zl -Mh�5kID��&�"�<m���s�.T�v�H>���~5l�H$��j��un�j���5����PܝRk���a�L\������XTZB�Y��i`�>@"wu��H�7"#��*!����ze�����	s�j�WS<:b~ T���D��l�|h�rȰ	7���G��u� AI��3�v ��d�m
�._2�ł/u����"5"}��T;V���+���߀�!���"�3�sڨk��h��E5��b���l��`� ռ��}��dldlݼ�[�l�i%�!�*���YBh����i���%��0]\K�֠����AS��$��(O�B/�0f�����<oҮ��(�8խ`�32Kd� ��-6(]M�(�ȡ_}W۰�+��W�?����w�ly<ˬ�[WF��7`��w�3tn{���&��,���4sy��q"���oR��$H����F>>��'6\�'����h�����6��t��˺�Ax��i�Aȑ�1�b	"v��}m0	�`����躔��%ڰiO�Ͱ��SYr��o/My0�C�P� ��^+���C|�.�����X�����d�ǅ'�+��g�%�"Dz٨x��o�	��g��cu�cXݎ{xI��$řKY�aunrJq�6��˄Ԯ�Ge͌(^�����v�;;��	���@��l�(5�;���_��|�_���}�*t�)�T(;/��ݱ
���
5�bf>^���A��N����s�C뜯�*�r��I6�I����n���N����G�������f���f��Ao!k�6r�$I�9O��r��,��xJ!�Mf�k�����7[��0"��v��.�<(Tz�T�5��0��&{�b�T�P}k6f���� �Fy@ְ�3jտ��]@�^���%�����	��6��l�ǒ5�1���٣�[#sW�E�^�$	��rI9��[��}~����]�3�c���*�-;CF5��\�H�մ���X�V�|�'�_������bU}9��$	�Ȉ:������S�Ua����������H�BS�ͫ:��o�u������ �l��k�(I$xO�v���|��ޝ=>�=6q�Ĉ.�I���[ʛ�#�u�	ٕ\3!���n�Mݳ�	'of=8��38NÓ P�d����m��=���t<=��w<H��U��=����<����b1a���;�j�+���|z�]�M�+��=�J,5a�;��b��@4�׸�Nm���Z�&�Z"��{�j�p%WX�X?/�j��/_x*���y�6�g�/>2ה�"]����u~�?|n�<�K[BbH���j%.,$�a�.n[BS.t3�ck��Utx@��`�]A~���W�]�;	�H7�kY�$ۘI���P��,Ƙ��c�5��H����҄Q�d����'�����y)Ȇ�O��A$�����A\6j��H��G�A��UN�p�D�R�6�
�2X���sY�k-��A �:�Xk�6ؑ�- �:���#7���C5�
��H'e� I&v��v> ]�%����$�N�Y��e�~��U}x};{���W5
񓛍�9jR\h�$j��pՏ���V�/sa�]��ۘX�H;��B�pٻX�(�iV��30��v'Ϲ-�)=+k]�Հ����*��T@e�qH��Ak���m���+A5����,
�f�rZ�0[H�7�����]�(&[q���nyCUݤ�ö�5J�5Kh[7VGl �Kq��J���jй*[,k��cX�Mv��Z4�3B�@�4��vH�KT
�`�k-fI�K�R��F�ڦͷ-�	X�{<���$Eͨ���#�]�5\F�:����K��@pCv�4 �
�aVmImf3�f��u��5c��qD�`j����$QI�)n�'!�p�h;1� ���y�� I�vs�Qw�ѕ,�WWB��s�W�{&�_&�-�EԂ��m�ĕB��X�*��	Y�[u@$�gڝ 0d�wՒ�KfǇdp�����gt����D��c���`�I�����*�/�NJ�P$m�955�U��"!�eZ�����V�N����F^�e�r���q<!z�pr�]�Vfs�}!�t �Mۻ��MG.%��'m��H��pI ��/>m�{G����<��t��n��v��v-�m�I��2�U5"har`m�-���;��=�{k��9=��5bIZ��/i��m?�]�6��m1�}��R��NC ��Ҁ��B������Tv��!�ko�*WZ�|�M��P�����^r�g��D=�F�E���LA:�Q�����fl�I$�[y�����멤,�.����4i�Bp�2Tk?� ���O��1���;���-�5z�O� �v�� ��W�6�4���Z���@(S��A"+"=o��Z�Y��5D�	ї�� �t�,pPY����K�~�w���rA �l8�H���p��;��?5�z�yV� u%cP&�l��z�v�GcJ���dd�"�<)|>|=�ص��y��~g����ˣ�_��]�I�����ڏ�uB��m�]8�(�@�I2���T4�_�x�ɶee��
�@�m��A�����coy��+��Ғ������kOCw��"�s���#@��-�5�����w�[��U�L�S$[p�AS4���2
9"e�%>��e��lR�&��umm��c35��A�8+E//2���C-�r�Y�2� �T�.��Q��R��JE�ƞ�F�ç�fcs:���b�c�w5��o,���,p�S�y��5?�կ�Fpe2��-&�pYҋ��3iM�۶��[�����9�i�(k	AX �ovv]��$��b������IA���ڼ�n�M�%u޿(���y|�k�+z*�NJT���n>g�^��zP�Vq��5�an�K5�˵�[��l��u���V���Dn'(�BF�9�Э����zl5�A�0�|��D坡N�%Jۗ�'��nMV�W2�3P�u�FgoQc�&�Wͭ�\����rpQ[ŏ{� ]���Ӳ���Xڋ���K�|ܕ��zu][ǒA<�������� K�f�nR�l��5:�^o^�]�b��0=Č:߷U�3��������x�����vK������k�.Y�8�ZE�O8C�c��jq�R�j72�`o�vc�R'vl�Jb#�ܪ��@���xdy���
S��cn��^��.��h�,-��r�q������a ߘ���]�}Ӯ���u��a7�\��۠��6D���݇��Nn�0m�	�E���� X��򵢕lJ�S '�O.K��Re\�QW��=q94�7cWVGz��3�����gWc~\	Y��O*�.~B�F�s�[�I�<���1"X>�	y�4e؄�2n�]�0���p.Ñ���2��xg)R��2�b��*\��!X�C&w����Eֹy���#����7I���{�23��gs���rlٳg�V��ˀ=5d|Ac*�!��֕v�,�����ʑAL`���};��Y��w:��y>�NM�6l�"�*����%�&�5����T�-d3��U�c�*U�_���},e���Fy<�O�&͛6os�J�EYZ�i[��s.-�#*^�9j�zZ�+h�@PX��-P�+l�c�eI��r�#[��WZھ8&�1���en	X���0�Z�|�j���1��2���[W)ADaiImXc�����Ld���I�u��e0��LS��� �1�k����w3���KL0�AT{6�"�Vª(�hk0EUZ�Je)�i���S��th(�}��Rc+l�G-1PkJ�����2�ˊ�L�Q��j��JU��.2B� u��Te�ލ�Tׇ��a�����<	�r�Y-?y�t��l`VAz��s�	S���g^�׆}���nen��X'� ����oc��*�� i���@@��7���铤+%aD�����}�+ �'L���u����{�r�u$��X�N�u�2t�0���}O*~����7y��=�D�������$��- �����]�����es��bE;/�;��2:@�;����+ �ЏG���s�|)�6nz3tr�����{���H�b�4]EЋh]6%t���q���,�1\5q.����[�z����B������'T��������'Q&��5�XyϷ�N�����XG���R��z����m�ׄ'���u��C�����C��s��C�����X�t�]�:���@����pd+ ���{�}����I��|�����!RE��9��T�'q��T����d�B���秛�{�^�l6�{�D�S�4$x.��	k�Y�e���?~�}�Gi���R~���!Z���=�h�����>���;`VT
��}�s���S�J�~���{��_g���F��9!Ϥy���Dd���Y]��o>���!>d���T�{��t�dJ�{���C�Xw0q���~��G��ٍ��Y�770W��6<s=���6�E3Л���5�nS�k2Qz�
+ ˬgL)y(_n�{Z*>>�v�y���������~�11#�$Y$_��y�y�T�BT���L�1�������`v������� ���]O�ޒ��e���=QQbRs}y�q��|��O���p@�	�� A�|q���Cw�l`��'�5�).��$ř���3V%��J�ev�Q:�@�����t�ĹO���~�8�R�c��f�J�����J{�����#�������;�4S��s���%G�Z`�P�O}��aĕ���z���s]����,{��=��'��^K��.�>=x����������R�,�Ϸ�5�Q%I2���g��!\��������GWz{����Y�ȍ>�؞��۸��a�C������8�VT
�d�����铦AaD������o}���|����R�I9/	��Υ)�#+ĩ�׿�N�S���y�ޖ��;gfA@�#�G�v�#�O��	�%��d�����Ax$*X��q�׀�&W�c�|��}���@랉��є}���CR!����,9�w�.���·�q��0�����:a�%(bC�=�����f0?~���;��翍�(N�����D�p�HR����lؓ���q!ZZs��� ���*q�.X�46�x�p}�&�q=b���3�U���ù�+����_VM�X���V76w�b��J�I���}1@꫺�������� �ϙ��Ǐ�	m%X�m]s/i���$tI�%��ͮ�	j���x�{[vp�ty���-Q�u�F[M�F��	�]i3i��#PZ�WF�e�k��H�R%�e�e]^w�1
���h�Ma�۬#qf�k���&!��7��v��=A�&��Πlтʢ�4Q�֕�]L����3����B�4T#�E:�j\P-�y�o�����XMI�4[q�����Yk�%�8��)����c�e�hef��bΝ�"�L��4�7N��P*��}���L�!D��bJ�WD��>�$y�}��Dx�wd�!P++Ĭ;��:H^��
\�3�� S��G�|&�������9��_O��F��D�h��&2
~��������e�_������">� 2��nayTpxMd;�
IP>��߼ϰsn���w���x��7�ψ;���\����|����C�@�B>�$x0�=]�Y�E��N�x!Ʋ���!�:�65�\���~�*uJ���F[w���'����c�}���:�����L��c%��:���ڗ��l���ߟ}w���%�+����G����w�Ϲ���aA`Q*~��h	�B�����fne/]�;���@� �����wY���w<3�=��btJ���p�I�0+,@�=�����u�@F<G��{��{Ā*�{���w�~|�>z���}5�K^��Ʀi�Fˉ���Dt�kfi�e@��|����AѤ�O]�I�
�g��?:d��X{������,
�!K����AH}}���ϳzÞ��<I,�����:�VAh��7ȉ y�<`nI��vH��!@S��z���8�P�����_�g��6��@3}{�֦��Ư���tcuZ��iS���݄p����m:��=x�w���i�F�����N�>�d<���Ϗ���0w'%(�K�?�Y8�@��ya��~�{���xY�N �$����&vvd
x;��+���r8�X[!e�����09a�ISP�<�n����3�?l'i�����?u�=�+ �� �}�������8ww(��$Q����e���- �ػ!�Q��bH�9�<�	 �+�VƮj���F�0  �N9v�'��sЁ,�4�	����@"{)�|�Z�Uv�7*�/G��Jݧ��$|�@H%����$w���+�c7���FxD��H�A�Ad��Ӱ�\�Q�q�)԰m��8���Z �i[�}����CE� ��x.�W2�$I���ǒ@$�Kۏ<�|��:"���Jc.s����|��rҒI%��V�;(3?��̓@M�'��P_�x%j�v�X�{޸u�� �	"^3�I�3.ǎP@2���:�\C�n�o_��9MY���]�"�̋� ~�O�@�|���I�'b,��Q��ă\�M�o^z����$�*�7�(��� ���Xѝ��]���D�r�C��YUB�P�ꕈҝ�oh�]2$c:-�c?�(3�}������k90V�'���R	�\�ggL�O~5IzUwCn�ܪ��0��W��>^)^����ګ�]�n�lT�< Gv+�}��,T-��!fe�-�(<BA.3�!e\Ocij��ª�j	 e� Iy$�&0�o)�`T�K�BaE��Tbc�`(u$��,\�Β?��m�aP��`��Ԙ��f�Bdi,̥���?~O�.-i�b�$���v��	w�d���T�/J��K�IT�٭�|�pܴ�R[r���������+uȧb��)�I�ǯ%̤er�W���g=�i<��	$�ImNș@$��=��!%�%�o�K�����k���?��o��ؤ��}%l�ęt�*3�	 �	,�Z�sk���,�$��G�!,3�1��ٷ�K�-��H/��u��U���i;�o���]�5�E/r��yI �	ns85ry�(�{ʸ{r�����b�ܳL
���`:p5��Z�dY�N�*�B�R��v/�	'��U�K:���u�ϯ/�^�y����ۮ+����FX�2�2���U�{���.?�_e��dS��T��}2�I�h��I���=�[5�dxE$J��n�i�3���}��Ϟy�Wx��n��f�6�X#huS6�4ɩ���i-���P�	�����C5Et�m�Uױ&RDҳ!�$ϗg4B@g��J� ��wd�L��B=E�����Pm��'G��7z���k�I0�N�h鹎؈����+Km>�RT<�+9����UIU膹�x)��)Fen ~ �h*2�T?3�2I$��Wd R[���S����Q2�I%�ے�	x$�[��	�j;~L�Ô���.��w41�󈧝����I%����Y�٭ ZT�yZ���Z5s�g��Qk�U_U����B ���"�'Ē�3�AZP9Y�y�=d�#ZnZ|�)*�`"$��D��lͧ�Wi����ٴL1�W9���ǥ���6�7Y�n5pV��8������[����3�Y��̢[2�(KIE
���>��D+�Oߺ��Q�0������-їM�Y�\�ml�u�(���X��z�u�bRk!X2�F� 6XR3i��h�l+mh����U��iN�6�MLX4�k�(0@�-�Gk(��hS(:�L�iIM0bm�qXh���TKm�.�`�����f��1�In�M��)�3b%�O&tR4��W��Z E	��K�pV']ɖE(,%lc��ю@��bt�#�<�%�����<�JKI�����Lk�6GM��a�-�t�Fo_��~�I��t]�-1*�7߁�^H���I-��)\�R�}�O}D�������B@~�0=~���-T-����4��ohR�
3����p��jUq'�RH�^3�	 �d�$�u݉��We���!�*�؃��؆� M���АIy.�|�'�����I�*���X��$��=����[�̒�bL�Uh�$��3��Wz�i�j�F��=.E� BI(U
!!�f%�l�>�Q;<�]F�v{��.	z���UhńY��)��C�K&ފ�nx)�fStI��sݺ̆�j�y}䗥��@	 �]q@�J(K3uk���Y�'q��zև0�f+MfW�.CFj�6�˥-6��n�`���Q0`[��6�w��'�!_y�4��H%]ҥy#�R<�*Rc�X�¼��Mܣ�$���e ̼ɜ�	0�	�y�	�32^l�`г����=ҥ0Շk�A7�rZ��Fun�������xeA�y�[�g��ov�ss���}�?@�a�!��S0�9{���� �5��@W�fK��� �I*����P��':�-��gL����؍��`R��	t�DJI$�T�sv�N�Kc� ��^���2�	.��L���"����@IuέM"��ºI�o2��H\�D��)��չ�պ��}G�T'zw�$��d0P�v���"%"W��x���:�
3��a�{X�k��fBD�WVĒe ���Q�A/Okz��	�o�&�1ip�R|����	�D�]V�洠�3B`P�͔�d��գ��S��c7W=RoKDw_;���Ȅ>Wt<B}9�S��oU.��0{�s� q綴c7'v!'	>��E>�I��! �nT�h�>mƛ��7���M K��Ʉ��1�	T_>��n$��e�L�I�i�g�]z5� $�;���
|�%y4��{���_Kʗ���%�����k������`��oV^�x�/�֡O�2�)ѳ:�K���.d﮹�����$@H� � =�Q�I�����>	$�ﵣА�iζ��3�wH4Ϭ����<Y�t��A "w�%%�H�4@I$���&���:
+���̚x2Oaa���^v!�$$������i�6��uŘ���f�HRo0f^K3=�*�\��J��
��A�}/�Yeh�b���8�P�2�B�е��)X%\Va���0r:��G�`��:,U��j��H^H��@���)$79I���D�ɡol���oʃ$�%�-"�q�ޔY��I���'��p�Sjڹ�Z���a$$�^[���� ��^eL��E���G.i3�ϴϪ�G�''�����$�'T
�	u[D H����IA$;s��2i�Q:�	v�?�RIv<r�)���^d��͞UJ)wH�1w�fa
d�A#���f;0*��NB� ����r�6M{��	�����j�����of��VsV\X�[��$��4�4!��V���s����2L`�rܝ�3�I#�=��������IXB�?�2[��y�'�߽�j��N�Һ��'Z�������N�r�3K��$Qv�	$��x�2��3��T�s{��k��0�D�	Re�k����]0Zj"X�df���ol�&��e�h����8�$엜1i�o�}��w3�a+�^�)$Q\�z^R~�茜�t-�r����6  ���j�lk�#�L��
����Ŧ������'{����"	�Sũ��@-3��F�T#i�В����|9�%��?8�oL��t��A��{h�iI `yQ[��B@ 屗}Eir��f���$�k� 'Ҋ$)�&}K#�����T
D�,�F�o<T�� H��̖���N伤�^Ko���L�xf9��>D��iH���ňd���d��ؿBy$�sG�K�\3R1�	/tvȒ&G)ޗ�$�^K�� ��{����u�X�W�s�`��뵽���]��t�c2��a�|{3ks7|MD�m�"�=ݨ�9�7���[��w���ܯBZ���vYM�q +ƨhw��r��-�a�T�$�Ѯ���xr�9��]��;��h��m���X�}��2��ħ��>;ȓ��Q	�DC�,�z��{�oae��X�Ú2bR�vnH����;t2�M�ٷn_�Ϋy�VN��mԜih��w�w��ٽ-�
������f�6�z2��˄��D����nJ��p̔C��g2)Wxs�7��;1�{]�s�.�j��'\Ӫ�i�����t��2��or4^���igKƵ��;Z9|�U��E�����zM��Ğ��2�ɂ:��7L:Z�X�8o��rZ�1bR���9s*�A|��g2��Q�3�xfo|����4,hw�i�s&\�˰�����k��x<���))�
�B��E l�鏩[Σ�b�e��S�R���[��a�Ы;\�VV}ݹ�jj٣���s�b{#�[���]�Dk��ӫ�� �6��6���U�/���(x�x�.�ٓ�ы�݅�Q]s�X�*�(����J�I�3��<Nb㗸#�0m��J�VT�}q֢�,[��ݺ��+�v�j�äX�R�bq��!u�]��!:��]��V��G�R���af�gsw��u�����zR�x[Ŝ���e�wg���v{7�R�u!H`@R���(1��fS��^��=^��i�r�m�Ɯ��˲�n�f���MW�}{'ڋ��������DE��f8��U�Wmi��e��[�VQ��|e�U*6ү,��*��NOg�c,�3���gs��~�M�6l�8���e#h�*��U����x�Z����Z\
��c����>����������u996i�-G���+P�.9��q�Z���,Z�Z#S�sPD�%����_���w,e}��������|���==>�Npj� �[�{�\fX����e�-ZУP�cna[eR��fS2��\(��TF+ZP���XZ4��QkQ��Z�ɅbX֠�K]j�erܶ�3
C*"�meEY�*1Q�Ӭ.qƶZڱ�F%���LE���kj/L��J����(��-[c��bjU�E*��VB[zƖ�^,%
�X�KA�42����5�AJ����F
Z��j�bԪŮ�1$�qEA`�mQV,��V�&�D����q������Y���X����
��ZYEDP�|��wj�mԷnR����P���`�4�R�,n����	�u��`.��s�V�ݘ
$֐��BVg2�6��XѶ&e�`��vn]a\ntr.IM恈���[�jB!-��`Ƃ�4�C#4u��Xh�CQZ�,��0�����V�� �LL�Z�m0���2Qu,ȸ衘�%�.�فMՙ*װ 9��:�k����.��� Z�@N-�m�%�4�Ж�\�4k+a��Z�BZ��sI`u���w ������GV���תb�,0"�sIn1jת@����jf������,�RҵΫ
��+ɜ����E,t9�.Dr^mLjXa3(���I��(��+�nͺ���H�(E/-�[cVdжS+�P�M"�A;l��.��KDGj�j�mt�e	J��m�@[E.�S��X]�����al;T��i��r�t��iMɡ�jCd5��y;e��a��]5��!�2���ڶ�nU)�֥�Xv
Ͷ�em�h�b6�
Sm�[z�bhAѵ�(��۬XL1�a��:��A��6�k�f�s1����`	�lq0fX�CkMMm���M���ʹ�s*�:��Hu&.ꉆ�l��gV+�0��	��gd��U�uC��c�j�J�BU���nc�b�
���tÚiR�t�����M��Qs�[�l��@���Ї0̧R��F�=HY�WK�dU�q �)U(�����XV�c���#f�v���=�����\�JqGB9���4��༶�vF�R�\@���1�$fR� "��e��-6�۰�EjB�jl�j�-�S]A�)����,�.���^�]BV�V�5�h������kq�Dq��h���){Me�(;Sir�s17�esc.ڰ�!.��0��:�3*����a���Ļ2h��A%�Vk�-�\���̬Rm�zަ��7B&. \���u����p�Z�؎��ь���G�'c�0"�����g3��X�v5��m�,��f����h���X4�-�Tb��R��˱Z.n�bŸ��b)!5\���V���aVX�]7
8-�ɰ���9���#uIGJ\h�L?�y�yRX_�Bډ V�ĵ.����,����-U�il*�uՈm*��v&�8�s�Q�ԙ�bl�Ŗ�U�,���cX��ꀡ��]̮�e�7�G.�����ۥQU��f:ܵ��7��+5k���X���å��p���&,]f`�{~��bY�8w,�@��$���	�I>�9�0�H$���y葷��`��V�ޚ��P�̐�Y2�t\qX� �h4�?4z I&�pB�t�5]S��2�I"<���^BD�����Ȕ+8�b[�pA����,�3��@���*�a ��32=���D��]$݅���M��!%�����$�.�g��!�֐�%��'�n#Z�����&eǣ"a �A#����Iolυm��z���3�[�/)#60�dAN
qsD�	e�-��I��bA�l�,��.c��d!eԼ�@$�s ��K˺6U��!�����Ӧq^MQ4RuE:)�*��P"�0n:��Gq��X�ms�,٨�߿E���T�!���bw�-$�ȁ��K"��ꍑ2�3��Oo��ʢe� (%ۭ���jbY�8w%�UW����$�K/�7UѾ�w�����غ�u���\�s0g5K�OzA��*܆A�6^����^���+�v��������i���˿^|�~F!�d��#�gz�����d�f� L$_}"e䵣kN���ЀW%*�vd2M)>kD$;��l���PI�]���憟m'x���Iy+�g$�R��dL��l-E���.(w�����2��b��[�,�RA%�"[�̐LwC�fw4��Q!_��ILC@�yaJ�$S�f���K#2$I|��(��BhkX+�i�Y� }��SQ�&QIa}�yI��{��/d4q&�4Q3>gN���m#��4�1)�0�*�Ý�4ՅX,1L�`n��5�S��t�pK�� ���30J�z'��H�Lԣz\���{��8������T�?�}*T$ޑ� �&�L�@���3䲺�1�/vZ��B%%�$ KK�C�H�xtܛ��W\_��[?��wSS��9,ZJ��J�32�1"$M{Ѹwb!��l�ʹT&�6Tڗ�n�y[���C\��IÙ�L}��m�Nh����F~��8n���L���SI�Q~F�@x���>�FyW��6����?�C�K��K�*�vd�M���ֆ��`[H��N�J��$���I%��%�$�K���q�)*c�	.�q
*�A��
���G���,�~J�i~g�>���W^�%��s"H�����^H���|�7m=ObO߳����!��J�J��7m����滳 �6�m��U3�c���~ߒј?��̟��܁���΀�) ^4@K�ܡ�4qX�����_OH�E �r^BK���f �8�T薏@	%0����U�YP�$$|�HR}�yI$@=�������9;�uQ�i�)J����f�����݉�I ��ƀ!?�	�Jz+N2b�hw�~�4�H�����D�����$��َ�ӗvN�Q$��	gk�5��{�����fqH��LO� �	%�W�I |������J�3m�g����ꝰ�Lf?L������}¶h��u:�*z�����q���h��O}s����w�<>P��dC�H��� x$~IU� <���5+ْp�`"%'�h��C䩆�b;f
=/YW/)$��
�Y��C�UJ��~��Yv��U�E�lQ^���ՄѸ��(F�n�;% �#6������!&E����L;�8`�Wp\^�f���4z� ��d������ܲ�%sp�I0(�Bm�ARF�Z
,����1ItCك��R�%[�m�p��3w!�_4@I�@-�2%�K����U���<����e��18I�
��e����>�R� TB��\d�������/$�W���(����2�CCN)\���3hU�&��s�0%���Z��� ���K�t>�$�Hr}��綞CgΩ#�W�ss,��,��Uf�W��!I($}��bEzZ.�ai�N�3�x�d�\���uH�W�	y{Y�!�P��m�f�_�|�̓���^F�h��h�u�nf�� 6ag7�����R#-o�dX����?{���x�����BC����}�ǽj��v[	WA��.��R�:�[R�Հ6J�g 3`�ͺXZ�!n ��U�tL!X4��eP&`��]��f9���m�����gQ���Z@�b��^�ix@݋���s�sRDȖ]� ��JA�.5�^p��&Չ�-V�&YSe�u�e�����q[�`�� `�4�-�&��"CM䍺�RmV�[1��5�a2�5�GfF��]6�U��Kt�R
�F��5H,҆�6BТ}�6��F��/���[�-'� v3�I�Z6CW���(�M�{��,�9Y-e���z��a&ۚ �I)׎Pf*v�L:vp�������ldO�$�ܮ�[#&��4� ��x�2H������\�׼�̷1�Y����ؒ�)1`�Ld��	t�T�����Vc�&L��� v4{-[��`KY�s�ǵ�T�P�(ޗ����4�S�%8d��[K o�uSN�Ia��7���&�����r��%H�~9���(%�͓B�2���^�.|�Q\�V��K���س"�<�d��p�$�kD ��b�4Ѵ��)A �"�^K�D��]��F�K�X����x-ħ.|_�X�$���۳�8\`�E��v�ѶP���ǿ��*S� ��|
�n��($	q��s) �;��_��;7�l�ǘ��S�ʑ)������IY�2F�3v)����>ˤ�K`�@7�����L�SAC{WۻKr�=���W�n��K��N���[Zl��79J�sH&�T��s��&��cU
�f�ȿX&�> �C��U�!�X`J���O�<�c](�$�	|��^R%x _�&�$��<BQ=,�t��B�;8�L:vtJ�wi�]́	$�H�cD$H<���8sO��)\��GԞ��AH$���4z RsR[�$�?��1It6�(�ճ�����Rӛ�>����32 ��9 �Iyo<�k�%��֋�
H�� q>����@.�u��P�ͤ�
y�TK�X���c��5C�I]��fk9 BIO<�+b�9X�:Ɏ�[���V~��lWH�m�42k)Rb�Y��\��MD�V)*[i�Y�C^�ߗ��[���}����Ȅ)#y� @	$�^�y�2�O���;"n�R��y+@&�K�!p��֛m���uY��u���K���x�9sE��Ӳ�@��4B�3y�K�ʹA2��^X�"s�_�H
�[�:v,��O�O�����R�H��{1�vF�vn�8�"Z�2е/:]`�����U��RL;���E�3�g����W��j/ȶl�AK��@y�C�`D�PH`0			�ﯺ���}����?gD"�3����PzC&r];:UP\jb0�X3�1.7- 	/���0H�s)�ĤJ�����m�ԚF �ǒ�֏BT��Z1$�?����>�VƾJ��{<���;�zߛOb���+�b�餓�s� G�y�̍Կ�%bކ������'U� /G�*���aZi�ͦ��r�؝�B.�un �K�R������]�Y�>�d@+�g09/��A%�z	�[��&c;]��\0s�Y �mF��Q�/;��LK1�/B�xt��3��y�0<Ю��v%�a$C*"̐yGxxً�4��$c�i�m�/*y�e�?M;;��:`��UPJ���(a �=�^|���̔�S���:�@�Vcm$)fDYg0���K3{pC�nN�`���SIC�,ͺ�j�U`�7��z׳�R	/V�B�K1� ��v���xn����PfDu�6J�&�X�^������ozp�Of֌�ŒӇFh�q�uV`��lt��I�b�p��|�'�ȃ 0�
���$��Х���������S.9.���}�VR�����̏��r�a�Y�lAe&�k��G�R����$�|�� ��$�����C�=^��{��:�lU˵��է6�#���\i���&1 �
����L4���I�B������ݎ@���3#��D�	;��i50�Yioh�ɶ"H%���l_�X]�A[L�KA:��{Ĺ���T[j��R���s�)$	v7B�$�K�ns8��컵o����A�[�*Z���1,� �ߕ:�D� $om�	$�Pų��w1�)"O��ܒL%����UuS��wN�;9UT�Ot_A2p�}"���Ql�	$�5|�	/$�Gt�dfh�zh�<A�^�p��8%]d���~T|��'��Bd�f�%�w<��I$�ƈ@�f�F�]������n��uh��s�)� ����|�w^:W/*ێ�*v�k��mf(w`:�)�Na�>��빷D^<��>�~Q�e�PX`Qz" B(He���5�7G\�b��X�6���+��4��(a6ͻK��P�F�	f��ܥ6�;bf��ți��њ��h��l�e�4ʖ�r6�Q�U!z��6�-0��15���JYeX���r�U���`M��m�]���F��80�nen�uH�&p����j�&�u�;�5cCb���q�i�if��9m:�a1Θ��0I[x�M.�K�&`ٜX���ˑ��A˪F�]�bWR����r�'^,J~��fwH���T{�K�r���"K]��<�I$��ޑ$�]�A�/t17�%�ǂG����sL��\��;��I>�'�r ����!m[�;e���� �	#9l�	 ��t���L�Käv眿5 k�+�
X���'b�(U%�M$���eIsq�M��z�A#�R ���I��% 5��8��v,K4
�	~h�i����$'�!  �W"e%䗷��08Sk>G@������3�wf�S�p�;�S$����$�^3�I��>��g�W�p�,x�;�.�FB����H7s������鈬�M2p&���Rg.�8��Z�lV�\K���Qb��p#lG;).�,��,� �e»jr���Р���� D�"�a�Ą�-�x0���kK�K���K�#�zⳐvwL];�UU�m�*���Y�[���@F���o����p:އ�ײ���{Χu'#n��զn����]��7z��uy������g����T�W�@<��d��R��Y��m����y��	����AW� �)�ut�Qf��i���%��u��Jz�h�2>��x	���~8�c�q����=�.D���!W�}/��I�s�/^FD��œ3�W �v��%��YuJ-��Iy ���Q��'�ndA��3$N���*/�?�n0h�F�K�!��i�F��w,K44���I I���n�X�.�B@%渎3)��� Ƞ�;؝P��N{�U�V����G��T^Fn��ky�@�6�Z�k]������dkm%<�������;����]>ʛfc�W>3�I$�Iwdy��2Y���t"̴<3ҊI�x1�^�T�9p���Ā�v�J����=��V�1vk��|��Wf� c�g����h�@A&{ܨ�ʚ�W�[l����vgLJgA4�-t�D$J	 z��H� x0�����Ɏ3ΘQ������F���M,� �`mcVUcʮ �Zz�X [�b�n�6kj�������w�U��6%�;.]�=�#v�֥;;�Hxp�N�@m|��T�/W��E
��3*@�X0�ppt��]Ud^��^�aݥ��s�U���~A��ס]�t^���l�լf3\yh�/CVü݌�ەL����p���зX�>�u�	�h�TRbkc���m.��|��D\�po9ʹ�F)]%�:��ZAC����7}�H�f�{��x+Ua��\_���B��j 1��=�:�3`l���+y�b�+j�����|:챽�$��yX���9��)yO(����-v��ek�3h$T��ۭO/T��FV=^+_}�5N�Z2��"b&1��4�@LL�Y�Je��y��:Sع�\%br�:#W^x'^�(ڒ��wssyf�&�՝t���R�ut�Y>�K� lw.�N�f"�W5X�F�u��pG�3L^vR8d�w��׵��Wuv�f5U�f�R�ɋ�W*�&��WL�a�et7�߾H͝{kvl��	zaY�h�����ͣ7�!�Vڭ��5����${t:���Vo-��"�36+�f��Jo��m41������ݣ%��]EM�Ŏ�0�'+�tp���iΌV�q��pԽSr�X�:�k�g�p
�Ү��J�qH�t�*���Xw{�M�#l��o�α�����4{�6T���UVQ�.5-�[��`�0X�*T{'����<}3��������������:
*|R�DQ�V��"G-zf[�JiD���r�1kc+AX�>�o��>�����q��z|���===��A��*��
�kT�-(���"����1��*��))G9c�������=��_N>�oO����ɝ=X ��q�%+�aRX����حJ�(�T����Z�X[@��jWmq*�e�������7T���1al�"�QS.88ܲ��"��-3*
�R�j�C-@X�(.R�+X8،�QE��ʖш�b=�pESm�X[b̥TĨ�)j*X���EQk`�媢��t55�2�U�w���-�]h���2�b��f5�6��x�`��QPLQ1��"�QEDbQ
�������ja�b����2�l�6�Yq�� �!��9y~PSFH`P�Ad�"��$!>��v�_Ŷ�y����"@.o�@���ԙ���'�N��>��o:bu�-��9�p�	>�p	ԒK��@�v�qmzh#R�|�	&?�Œ~3�Q����E&Y�ݢUQ�,�J!$�����>S�杪f�G���I�$��p	��[�fP�j�e����}il�2�'5݄u��\D!��hhhZ�4�fp�v|��!s��wH�h�Y{��a�I �F��! I �؎3*��k��J�z;� 0�$��8&�m9N���'p�T���� ���p{��t�-���Y��RǶ�� ��8���[#���G'���o�c���ñ/��&k�K�y�T#Ɓ4J|�W�$�b�O��4$�ZS�f Z�P!O�Gc�L�@ �5���dS:	�]��g�b5�կMj@ �-��I#�}� A�*M��r0��o�wr�3>�6a��{�N�e�R�O�}�Y��>�N�R��FM
���bgq���{�;�:jݾ�{�����!�2C��'� @)	 �����^�I6r�y'���O�CI���LW�/VC<�z �$J�����BU�.N�x$9��:�s���u�1��vt��$C")���ڛ�.�F��-ٗ:��Idάǯ_p���A�.�'|��>>��H��+"�HH����
<�B��^� c�ˀw�c�D�*��R� W��l	]��uVH]5fC�����y9	$�缏&BK��$|�BM���ynG�.\���SΓ�vvI�=Q �o@��\�U��$L_��lLF#���H��΁"Q%��0�ES��ܲ/����r��x����I�T��"|���<HR��N=�I��I�]� Hɬ�A�
f�ʬ��b�3��JG��n��d��N#rc�Β�͑2@ ����I�,��םݍ2��4T5h�2�cw9���#�Y�����:uA]�I���-PF�"���6�2�뙎�ߧ�3-��zMI���!��T��������m���]au�Ʀ�JC4�H�,u%�dָ��P�v��Yb�..�[`���=sqA�{8)�5��t�֥�28�F �]vc��XK�A�X�m������lv�a 9c�h4��[r��9�e��m\�Y�[���7+4�XhP�͍k��)ى�Ulq�aZgd�n����UMQNV�lب�mc���Z�1���m�������b"���`�V\e,�٭�f�\2�k,��'p��;�o��)�S�|I۹��RD��9&|��l�Jzm�gF�ȭ���x�G_ɋ�'�����d"Sd�e.i��������_8r�ۋW�>A���9��H$��rr�o4z�\��־����D��[�f�)����y�	 ���ВH$���t�X�q%\�
�^I.l�BWR����'p�U�y��F
���Kf�H%x��I$��v��H�����>��|�
�ӽ��q�9wd���X/9��"s�쀺ErkW�rqs*�<E�����2��29��-&�&A�E+D��jb��dV�WsH�3F@)p�ťl��-�q4�rk0����җ�߯τ�L�?���C��T\> ����4��=�QO6�'�y�͚9�â��<ώ]�G���&��lXͳ��=���,T$Z�e�C���!��7Yگ����ɖ\�z��j������t顉VK���v7=wI�@~d�Byo=�?�$�����s�a��o0
�^�YSo�Q�	9��wD�wEOx�*n�	 �kq�S���m]WV�Q'����p	��� �T]y�npX2	�d��� ������XGqx��u��q���f��|U]��5���/cت�u�{���1�[�R-Ǟ0��.���;�ڳ�7F��&8V9��Y��� �|%�h�^՗�>'ӷ���sN���/ا�_�6�_\ES�BÆvt��x�f1�亯_�"�t�2�O����O����'Č�ȀKfʞ�Hc&�2!O���V\�;c:S��6%��@�^�J�ݨ7KUd0bHF#Gn� �ܺtD��Tc�����@$N�Dx�Ґ�cf(vc��y���/��@s[�;1NRb�<
i�|����T�� \�3nD�O���`�_�7�`�>!jU����;肷��Xv)�]�|r��<y^�#���Ѥ0��
��ڄ�46)1����p��Ŗ�{*�	@����)�l�i�����ُu�N��[W�`�0��϶�m׮���~��z��ԟ �0�C�x2�h@��z��������������Y;�pnh�U��/5`���Z�:ׇ��� ��jنą�뷭Iӱ��5�$X@��HG���M�2@�@�]�ܸ�A'9�=`��7�s'Eg5Z�|L�l@>�}���x�}���@��'���q�Ļ�>-�`��Eұ$
"`�-M6�Z�Dqf��$�8�ϟ���#3���<����T��1�'�oy�F��G����n������M�"�9�t��-QRP����D^��ֺզ���ې/�S��QO<ٲ&�,�>����A�b=�����m���Phc��*P�$+˟��z�S�A���Ȅ��o:i�g��=Y��B7`0$�]<H'�ϱ����!�1A�L%nCU��~�3n��ui��D�C�H��v�+�.I:��Ѯ�9��.0k��e��W+A�AxA��S1 �`d�YEd�z<�>��
����d��@!�l�!$/��<�ﾏ�����U�5xx����e�'�����l���j+ ����@��ߍ�bw?@*He�ZA�k�ѕ���ۦ���W0ͣ��0�\#� �ևKcZ&���Y�I��ۈ'ă��Ă�a?K�y�7j�N�屓RP��\�]���Sl�:�&�-:wGҦWv ���[t�<���p|h�v>��$s6��*�Y�-�s�m�	�S���fp]�j��]Ё����GVL�S������j��y�z}�u��:f`�.�$�C�B��vq��K)���DUtA$��j<A��del�����]yLk�Cc�q(�r�Sy٢A_bxY0w��[����5;�Z��l��%����f�%�f�Q�;�;z����!E���{IE�i�cszh��=�|U����t�4�!W5�K5�2��=y��<z��_"����2#��e B��~C�u�<��	,ŕ��ca�/5��
%��ۊF����#xJ�E)ts��m+iUL���@&�1ҳF
��0�s��i�]]� G�Մ�j��0�Jd��JP�
�Ǝմqt�cJvq5Ö���س^���YA#LSf��i6��������.k)	G�v���leZ�R�M�.e�T���F�#�Yt��F��kcXhf]����V1�&�!6,`7Y���cT��ԍԥ��}�vrI`�Oo��&���0�T	�� �{m�Vӽ�:��E`�H>'�-x�b�2�e��Y���u8��ЯK�V/!��H>�n�����伝?����r�C��M�-:W �~���� _�W� �	��|ލP=Rۢ	�m� ���	ءw\�;3����@�]����Ľ��1M�ֱg�/K�L��#{`�6`ipV3���v� �7zS�3G���
��6#�=�]�U�=�tn����@�V4r�I7ݱ ���h�D��e�<>O�Wy��O��-��A�Ni-��(���0[�i�+�������%`T[(z���K\��b�*�Hp�Y��H9��#<�#�� pv6��D�i���T�ݑ �����]��w&��Vz�a�x�nv[vqo8�0nݝ�	��v���@�!Q��u��`��NQ]ߝ�����(c�[�j�D�:�F~�%en�%<'��/g���@�x2'$80��I@�b�P�H�o��������p���:d	n��9.Y���_*6�-Ι&Jh�n�Z����<D���E{��� A�Έ=��؈7����8,��&p�A�5k���^�w.��H3�o �H,Īـ �@�n��)��wtDx���<�'gvvI�@�2�i�_��M��:1ݭ�u#4��x���'���Q�YC�3"���w)�N�äܡ�lXe6ٖbV��݆f�NlT�&����	Z�Έ�?>��ҝ�1t|�{���#đՑ	 ���<_��;�
�P����A�؏D���R�,����#���S���̭��j̹�q�$	��LG��x�kq��]X���m�L���)rjA��Q��'��ll���RP�5�&���3�V�n��t�?֡��������+U�`�\�ѧlW�����Ԏs�Lr�3�ξ�n߽�j5*�?����HpdHd@��J-(�~<u蠦����GD������^O1p�rɘ�)�U��x|PwR�~ņ0�#�zl>$���9���M�8=�Ķ��� �tE^J�����ᙃ@�(�n���6*�ಅPz럶�&�� x��{"|s{_A�"6�L}w�/�������ttS760D�wSG=R9x ěm��!�,��o��ׯ�C;l����\}}���v�D����{�R7�76Y F�V\��A=��`/��;2b���<�n���a�!�aKgVz�y<X�"[^�H����m�NM�p6r+ }��M�Xp��k�I���x�HͲ�"�� �G7=��x�L��0%�l���H���z��k��
�,���<��;�@GĚ�ǀA<ݰ?!�H���ۑ�@7H\�M�11h�����(\W��/�L�:b��/X�ĝְ��cQ(ⓊN�u��4��Ylr�v��JD�=�x�?���!����4�����?�17?P�Ř�)�A��7�&����&_����l��'kz �9�c�(K[��!������p#�ڍ�4����f) ͷb\Ԇ��EcqŠ�Kw�pmpIg̃@�3Z�_�[�~��$�B�?4AQђ٢�B{UDO�{����(TF�	��˱r�A�΀ ��q���"33i�>$�{�`A �gB�-�=�l�UtE�uavd̝3��--�ĀG6\ �e�,�<ݾ���/ԥ7oH�I�ހ=�G2Mh�]˺y�{)�q�4��9����~�7��d@�$O���L�AǠ�[Z1�h�c� 8l��gD���gd	Cr��MMǳ w7/d����bIB��@�NF�=9��M��Ƕ���R���uk���E�W��r�
ߺ�d�sd;7zQ˝P���M��tΔR�{S�ɚ�Y��]=G9+� ����j�S;7;�>��4v��:2�u�SB<,U�]�S����-��(�ջ�g�HQ����뗝!ImE�kD3�6q��V�:���1o���4>r=�����]��K��4pR����d�X�^C�2��o�x^Wu���F���㈋��u�������:MY/�����Η�яo�G2R;�����iG��ڻgsŧ/��me�[c�WX���%�pl�
�0�5w���)��ӫp�CHi�Z��XU�[]�sii�Įg��",�
ە�R���ۻo�ӝ�N�Z�f��dX]5��7C�z2���.�7���X�i���{�W+�6m˗���A̴��wb9҄���i��������y�K���ӥ����Wu!�C���9��eh�]�1R�tep�b��U��g=K�6�ѽ�M�il����7D\���W�M^�	���
��t�X^�o�<�.�^�
��'u����8��ćf���a�����,Z�Z�XS���*�̡}C-"�� >��p��c��F{74,9T7���v��H�s�֩+�I�/���y�Nm��;�vސ6��GE�K�-s�@{.*Υkc��R�����q�Y����(�Xk���
5����I=n�>�����"(T��b�lN�-�x  (P�V=Yb��STb��ς�W,U�DQUAUb�h�9^G�ӯ<~����q��������tkն�U+F�b�H�ԍd��<J
""�AUqQKV�*�����c�������==��O������������j����h-h���EQ�5�W�\b1�PEZ�19pPc����q�#�;��t�l���}>��������߫�E�8r#''���b����7mDbm�2�h��b"��J,C��*���4
f\P��kYR�J5�����Z�0R���.Z�F
5��ms�f�e�j3�ň��X���ǻV"̲�J��T�,B�1�� *���|�QA���ڲ�O�:�UԨ�1�1�������U�����K�4� $!Ǘ�f�Zݥ�e�(*�PU&�m֪��J*�(¥LL0(��JU�eVq)�\J�Z©u+br�m���e����Z�T\eU+DQE&����se�rz�X�%	{�]bXj���R�V�ة4Z]n4�	M�B�z��� �Aщ�K´P���1e��l�`����ֵ���:9i���n j�1�J���als[MFʔ��d������7�m,Í��y�[��f"���;B撺Yl3L�Xݡ��Ƹ�&��n��:�c�,�u��!1J3[m�a�t"�&�V���󙩋bF�R�6�%a"��#.lm���n̙|wy�y�Hŵ)+�����X�8d�*m-F�b1�����\h���������jе�kB�qF�f`����%)��E�LѸ&�WbinH�a2�fae��R��ԫ�	u3@@v�h��fK���\�Tn�%M��UZ�#%��s�1�z�j��p�X���]�Ź5u��W*�vT�krhS:�s6�00u�0�΋uv�R�)���4:��H�W�K@��Q@j�F��jl�a���6U�ve,.��b%�����+	]��B�hժ�A%�qa�ԥ.�(��qM�;A.Ņr�kim�vi��.��/.)��΍#Q#1k�V!�f���F�+��0�kh�)I�1N�b��L����4�u�L��d��n���u����g�<�E�����(�6Z0�������J	WXk��R!kxM�u�T�7�:�رvH<�XnJ�ݒ��l��34p֔�3\�e���{mA�@4ɥ�P3�M��C��Yam���mvXҌt&�.�n�)U$��fi�rF�Kj���Ih-��W�Y\�-�j�.!˥�S6b�����,�*C"��+�6ق[4��`���b��l>�0S�̆����M[�ل�X�]v$�a��䵚�!���XH�a5�rY���6%�vPۅ���XY���h�e�ű��̺Q��[�Hjf���7c=�ZSe;i��[a3���MΚ^�&�KZe\:5(h�E[v��v���f���J�a�s�-l���;a õ&	���bhitn4k������B�# $`D�@>H,a��I;ި��;3m�te		��ʓ\e#�f�mP��k]D0��V˖VR����XQa���a`@Ͷ�I�5vن�-��J5Hk�Z���Kh-u�V2��f���`��Qr��lz��mCQ�6+]&Em�e��E�)�Q�%Vk4�Tg��f�a��U�&��)-������;IA��T�G7V2�����c\AeRٲiC�7R�hB]�`��+{:.^.�'��]��k��[5�!���.];y;�$*���'1D��ߖ��A׸��	,�_��*��r���-۳�O�[���R�Y�v!�U�n0��Kr�;�@�I�� ��~0@>3���ŧ^�~���ǌt�wg�D��ck�@'��A%XxYu3�׶�y58�<	�F��u9|]�3'�p�*������6�b�C�Hƻ���<˵G��>�Άk�����EU��zDf�k�D�wfy�n�j�P=��^U��³[�ٻ��ظ�H�^(�>9�� �whz�ѓ�[N8wQ�))c	��4�24�����점�h⊒��-�G$��4;X�,���W�� ��0�`1 ߐGٹ���6�_FD�]~� ���g���3W�K�.�@�U�7|�p �6ɯS���uQ.�ڣ8��G���݅h�J���ǷlC��a��O,�uZaxGi�I�~�/t��m����r��_;%�D ($�4�[[ݙ�Kwy��I�	�D" �$� � �B_w���������H'���O�|ȁb���|L�M�n�A͕!��%�'bC�Ϳ19�[��$��щ�n�OPՍ]��V3v(�$���DP�����3�r�Ux�nG�����EByQ�x���݈$���E�jB7ǭ���Queس38D3��U=oD|I��/�Q��ǃ�{N��A m��I<���k��[):L�S�tv	9l��1�L\�H-vnJ�L]��αv"T��*E�ʶ��rZ[|���4p�fG��㽼�H �HtlD���]�vz�R�D�����l\�L�� �]�ݎ�b9����+�I3Y�:B%>tG�b�t�MG!��m�8gd�M H� �|�A&_73�#��8]Hg�g��m ��T;8^�w���q��sx��q��Χ�R��e&K@�f�7��:Ϗ�^|^O[���r�i&����{�~FVF�"J�>>;���7��	���`An�s��g	؆��]�H�\7׬���xo ����@ �6�y�n�;K��z�ʼ�1!�Cs.���%h��A�[��9p���:=�$��}����>8�� �%�yAWvz���ׯ���>�_�K���Q�l��k,d!1��Vi����*����ԁ��翆��2�c����s�x�o�Cy#.��̹me�,5����� �	��x \m�g\�8wfx;Z�m�W��3m�x��Q��������^�}�ă���	J�=	�wG$�#�
%����	9sO �e�H�-�S�S�7`�-[<˹@$u�Hc���;$�h�]�=�n�9�8�U@�I������m�1��&�~�]��Q@��\V��m�M=w��`�vb�s����iT]	�\�X[&�^2�4Υ��Ǉ��9^�7ʿ#$20¡x��믟^;���g���4����b�(����ėxm�@��ǈ��≖k�.V�s�^K#S��6~|�d!]�m�TbCL��c	���f�Lv��XB�!(i�*]-Sޏ�(�z�=���ډL��n�$�܆$����oNՠ�it,:���N�o��z������7���pH��)0Ǥ}��ĎW�@�9C�y��q���<�X�h �{�`/��wrw�=�t�\A<�rħ;��Z�o0�ݺ�H'�ófH��4e��m��A �wv�{���+-%�A�����O��z�f�X�&�^_��_@	3]� �V�sSũ��(_�OօQ���Rh&�$�3��d�2@���e�͏[�`//]ep����@�%�N�������(�;�ث�
�9v���;X��n�U&�n��+���0
��f��G�*ˡ	�k/w��T�l�ı^%�D0��Ja��Đ����x�$`$�����WѸ�L��#��6�%�֭V6�[����:�҃�f�[l�uL%!f�a��NC�i*	,��H&i����vz�%��V�L���W%ҭ�ۯ�f%��4��U&c�쐌׊�V�t�;]���4,a]�����Xi�B��{�X�1��4&c+ m�U���P[n��P�i��e0xt�̬��aN��i�)z�F+Wi���<vā`53Z�RbJٖ�R�k]3]���n�����7��A�$�o� Ī� 5��S�0'ݑ��j�څjb��j� ߊ�c�A!�DRnb�g�����W,�����D���b)��	^�8����B�t/���1I8D;��U/z�� �A�qzE1':����j%��:~VW��x�ߕ?�'��x�D��ЧN� �*�1�X����o����$�V\��FWr׉��;6!6��!K�Gy/em���ɜb�" 2���o-k�q���y�����f�O���`�����~F}���S�Y�*����#�h\5�=�5Ch��p�ն&�X0���,����u3;wI$��wz� �n��B�D����~�ۅ���S�|�� �W����M��Aܤ�h@�kt!7�t:z�驛?��u�kp'Z=5���a��A�G���ې:�:�V���3Ka*��4�S#sl�����`<���H���g�i�U�����|�/��)�Jn��0C��d�g�>�3�p z-��$��$��ᥭ^�$���	q�� ���,K�
A��}9��s�}LC�dA�Q͆ &���rf�K
^}k҉虏C�rB��	9 �<	��-	�����-Pզ�$'� �k�	:��c�N�V��-����XhV�	�d�M���ۊ���� 4B�ei��,��WP��F�R�� V&��	k��	��FL�z���k��> ���ޘ7�����j���8�qm�`�}�Ι8fwI$�*���A �K�Ѩq�6�a�ك�I����GWtA&�ka"몫 �#�G+nv��'�@�E�H7��(�u��I ��\���o�3�_��|�����dU���	L�f�<�m<��q��yYW-����t���2�2˚�]o<��G�!��� +>G���D&�Y��ι�'����>$��
��9���p`�+o�K@�G���
��m��0����|���{N���k� ����!��Ϋ,K� �� ����}�$wN�wE���:�`5欎2�������#v{cl��2���i �n���`�(�֍����˦��l!���
5�V���0[t���S����:g�����Gē��<I#rz���[,��?��*D�|��fD����ӳ ��������������{7�g�:��H$f�D:	-�#��NX��?fTz�9@�f�g&�_�����̜&gI"�*�S�_�R���Q���G^�r�Yo�;��� ���-�Cs��w)?�'�'���[�c4�m�A��x$��B�b#ĂF6��ۮ#�/�9��Xh�}����x�g\���r�f��r�5�%Sf�!th��g����{a�����(�\B�n��@a#��uJE#%�a/뾷�ώ��~�3�3�pj�������1��-�(�Y����A&f����:�Hk��~L��������<Ժ��6�l*2�j&��3��q@u� _ߟ��L�|�>���x@#��zԓ�r���v1>���nyU1 �/" 99��d)��&b]�<	�Ռ|z�)e]�#��_���x�%�F�o(�����N���/�z���N���fp�|h��~�ITPI���Pdj~h�����I�m�b	����S���"\�z�w�k�����\A �O�ۭ���>9�t��΁��\=�h%�uk��ϵ/��d��p�����ok��1M���B긂I�n� �:�� �+{\̞�F%���2�*�"��+1pr�Ρ���4�����yV'�����.>c����ۿ��+�?��?��A%�0d����
��5���%�L�\u����sش�(���BS+Jŭ���g@��ʤ5ɬ��j�j-�3uu�W6����0�N.���f��ڗd�ցk��rS$��p\�JH�[�aqz�cf6���Y�t̹�ڵ�܅RѸm5l!l��m]�@�hjp���#��x�e+	CT��\fl^�홆�q�����72��z�õVZ����4�Pa6���,ĩ"��2�rٮ��ִ�X4G�����Cg��~�\@�3�t��	#�� ��sՍ5�ƶ�1�r�v���$\6Z�󕥉b]�D;<H��$�3��qneYM�b|���L�
	'�}� ܝ�� D���[d*��&bS�x��P�[k�	��0.�h��x���f��&�� (n� �6���	�җɴ�J�trW�|;���U�����$��ЇgU�<+t1�� �����Yp��L�^��v I7]O���Ii���$3����%M��sz��U�q|n`H(v�	�t�/�)-�\��mpui�3X�P��օ9���������t�'�D��i3�g;H�H��o7hFD"����I�݈�VY�nN�wgN�)�`6ׂ=�^#4�gꪦ���da�[�s��!0��cK12�m�ѽ���T0�]�Y��}������{��~"D�H���y���6�tA�G�Ɍ�Լ�#)��������̋�R�̓t��>$먂	&Bx�ݶ�{�S�j�H&�� �/���!�l��N�3�3���S+��g��nX�'ƺ%�Ē5�Q ��/ܶ�g4��=�Q �V^�rgLΙ���{�@�_nU/;���3�b�owr��ݐH�����q ���PY�KS6��_��<��K�{~hT�am�Љ֭�KL�1[Q��1Ũ梌lPpݍa���;���ϗ4�\ �;��"��|O�=-ܠ:;tkv�n5z=D@$���Ǫ����$�hFio(&��q��#�b�z>"�j >�m� ��ђ���)�}�m��r��t�4_d ��*��A����(Z)�oS�שF`�wMT��l�8�%4�\�7`1?h���r%N���j�A���.�p��O3�Ql�F�#���Qd����S�;�ibLT�i�rb�qK�bg�}�7�2�*����Â��f��o��媙���7b�T�=��v��]Lfj��D��W��q�y%ә��s��6{śB��V����\jj�oyh�̩O5�;9�ru��Ao^n�7�G��8r��l�X�Z�:`f�����W�|��&��RevĽ���W�9(�̉�c��k��Q۩!}�j�}�o�^㝷��f��
��������O�2>��/+�d�0ku�!ou���pl;���z���zT����r^[��\6f��;��ؓ��|��QEJ����]�Җ�U��]�gR�~��=�k[t,.rN���w���G�n�jŦ�[��r���a��7�
k�7$�3o�N<ib�3�U�i�m'ne_K1_a���ѩ?^ϻ�1�a>�zk(�R�QV#d�8�����6��n�ło��F��'}Պ���ݹ;}���c�]H�i���sa�eA�ɰ���l������`)�n�v�S�����{2]5�M�<7ŷBMŧ;/�[o_s0Z���Y[�<o����\G3�(��U��3}�gr��u���3x�G�����y��q���2�T�^U�;�I��6��W���U��*S6�;��m�/��I�*��RH,�Ȭ�����zn�|��J�.m���\�;�F"���J؋Z*�Ue1.R���UX���U��R�U��J(̴���u�/�g��������������ڊ(,EVEQ]����,^���X<�t%F�i�3�	��ȏc��ϗ��g����{6}99;�N�&�F��)Z�c��E��Q]|�V9VW�[r������T\V�e�c�*�>^���l��}>�o��������o	���'�\|zf�T]�EKl@V&R��*QU~w33`��Db)�ihbk�����U����X�+:�"���\B�VUL��R&�-���
�*��إcC�*���U��Dˉ�@D��S\��,P`�V[F%(V�lU"�fڄTV1Aq��҈�1Q� ����.ZEUAX�!��-2�X*(х��li�b����n�Wu�Tv�EF�T6�TW��V#^[�R�ò�������5(�Q�Zy�q*#YF*���v�G�Q�(�TTcM�����K@�����z�Ty��/���(&DuޔH`�R���S�@"���I~�G��@ �wB漿7B/�r�hL޼yN���bS�y�{��|v�W��]ՂF�Z�@����;[����������+��N]�p�Â8"�tXf9F��uҥ6̩�6���[��|����svk&b㞨��r�I�]��#k����ƚM�������|O�� �-q�8I�g.�i����^cr!B'Ď��P	� u�Cz<���p��L��Ӱ��~���=>��6��B�����x;�?����qq�1��V�g��$��PH'+z0j[Y˰r�Ӆ�Ƿ2D�k���Oj��I��� I��¯ )c�ߔņc��q��;XF�٥��q�_&@���`���+kB���v����)�hۂ��Rů~dԵL��+��bFK �" T�N�5����}��bY�H:y�� ���Gqu�[m� Ok]&�A>�;� �|{?eո���{��2�
J*E�I�E@�Lj�e�a�m*j��CD����X��m�+���=��J�
vg���TpbI��x'�����؈?n��-۝�[��'{� ���ڙ�1v,�ĹюQܭ;A�[��Đ	���-�{���(�؈\�	�Or�j�'Jp���]�&��=}i�o'	jk�r��k���IM��	3�P�Sl�����'bdĪ��T"��pIήx%���m�������>�el�n�C^dG�;�n��˳��݊�ު5ݏS��A�B�U��\�ǎ�'�wDǠ	�m� �Q�9cXo\O�Zg<3/���˶A��Hl�/�� �h����Y{���Vmiw}:�������Y��_5ϳ�ǻ�q� ��D��I�^����ܹL�2.�s/�lv�႙�+��C�mclA�#7h70��u�n���e)3��f*��s�^��,n�#�6`��� U�κ�K���+J��۫a�4�]�F�r��v�qKIv�Ep�r����]Q5k��,&A
E�[G@v�-�"[��j�ݴ�Z��4L��1)39-�r���\��͓V]�;76]���K+u�4p�җ�b���هM���׈'mvE����:'
`��������"��&7�����}��A��9s<�(��$e��m��',�N�� ���A)�{4�p��qM�<>� ���T7R�3��I�nm�3�2p�����-~�����$GZ���G;fi ����I��� D���᜺%�7�
�u[��Π�a�j,��9�� e���$�Ȗ�9����#�7�'�G�q/�h�m�iIT7Fo�Y P���ػՈ6]Q�y-���[�H$wv�x�>}y_'��)�M����4���Z��)u�k���*�
W@5��"Z�����?=_����gr��3�q�Ƹ���� r:[Y܌����vb��G�����?]i&E�d<
�];	2�47��b�23"�����+7$*�����c΃O����չ�6��5�ͥ�1Xee�q0�Fȃ&ϙ�<@$bD�B$az���/�n�N��ɂf髀���ރ�xFYb��	;;/L���$�|� 'Ɯ���t��� ��Y���O�rY݋'�\L�����l^ ���y�A�z�A3�11�z�ғ͹39l�L�IP	�i� ǐ�5[|S���t薙$S�O���[�t�F���"ݞ|=���i�UfDx���xGc�=Ű�p��8����$	{X�5�]�K��P�J`X^v2�S]�Āe�������mN�wvd��]�[P�M�sǡ/Ov�@.���$�5E'�B<� ���76����9r�ܨ^=}� ��U�����:�]�W��d��'n��x��ݵ, i�˛��v��^���Z��A8Nb��I���DA ��1A}�����\(h��.皶�6ҁM��V,O �z��ˬ�d�M��ԯ0��r����ŕ4��Y��.����DH�"��w���_e����r 9䏏}�V�)�r�$��'���n*�ܨ�y��%�x{�$/x���A3�Q���������8�i6�O ��v/�.�hk��>��Z^��]в&��E���D��H\��<H�m��:����O)�N�˻��&�ԅK��v�6t�j�+b�u�iC %.��w����L�h�n�#|�eDo�'���ul;&�dkO��9��'��eV6�wtK��A�A�,����]����؂�]<@�o($bړ��v����qF��g.Y��L��W���Yp�e�Q�I�N�5d�I>�G�仔���E�p�g/'#�3G0yy �r�� �[�$�5�.s,�����GU�uH�A��*��a{�,�V1U��H��Y��TJ�u�"ks�ԩ�%���7}[��V����%�%,
J
F :��u�A}�|$�p�Iݣ�{ʏ���VS�7N<R�!��#ă2��r��L�ά����f�4��a0�E�6��I�+��Rմ�]Q"�BU�A�c1m�R�Y{��ϛ�#D���9�| �2����'�k�5?D��#�z���2�Ȋ�~A��0���p�-�6:��1<��.�{"%^He3�	��q�no�A��Q�L��������^�sq�H)N!�m�21����	$L�ky�����x��p�Y�9r��Zg�:��R����+�c�>A�� ��Uj1)�f���h�bH����,���^���/�n9Ɉ�;�;1�"�A ���B% ���ި*$ks�e�T�~�l͍��ѫ��	;�q-�Y�����N�UE�SE�	����������CP��g������T6Um��'{_CYkq���D�"D@�O*������3)Z7h����ԕ]��a�z���Wg&4w`�6�eMi+ô�P�m !@]aI��eCA;UdZ�,�8c�ZI���;X��,�I�NG<-��8��b��2��lDٚ�jޱ�q�شQ�B�u�̩3 �t5���YnA�@��m�le��4tH�#4ѷ�a��	�9n�6�e�!ֆM��[(e�)�*W�q�MN�A���B+�z�Z�9D��@���?��d"�wn�#�1'ǯq�>���yD�� ��;w/D�lA"}Yyz�˹.K3�o^�	��_@��w�ڢ��A�w+� �H'�{� Ϣ"�9�̾VO�.')��*�UDA5�8�P ���&fx]uk��o_��	W���x{���N�wt�4
���w���2�WeL��"���H$+���$���MoV6��:�+�+���Y�9��ZP=w��8�X1x��V�`.o�s ����2k�$UN���y��~�l[�C�X�w
�R4Me�$�c�v;R5�li�F���3@(��1fv��)%$�����(8/�Y���uk�@א���>�$MSt!��+�c�bϦ��$��N@B[���IӴ��U0����g��7\!�]��r�"��Ⱥ�-tXk�]�U�N�n���6np�ۭ
���&��αyo0�)s����aJ��}�8{�@�ψ�X�k�/�;ϱ����k��r~�����6�a�M�	0#�dߠfV�1&<�$��YU�I�U�}qW�-܄]�jb� �bZdt�D�5f��>���^�ת	�����D��e�����i� CvEkk�w;�td���H���x�m�+�S���s��(2�uA$�_@oL��������_�������v���v)�-�fձU��llB:E!`�^t4�vj�4��|��E@]ӳ'�;���� �үa�'����@Z��0p�C9,��5dH�l� ����A�"�^rz���F��+�x�A��݊>&�� AMc9�+o�A����!�I�:�*���z�9�H3؇V�d���S���`|�W���S��f��"!��}t��p��4^ͫZ-��7j2���&n��9k�7G*�gǦ����O>}{���{�>=��ﾈ&;jw��`�C�8kj�c�e��*��z���ǒ3}� ���ˉyƍh���5.j#PgI��1�� �g��WDn����b�ր#ͭ2�Ǽ��܈$��tGN�춷�NO���"���ld�3DF�C-\V�=�wR	U�)�KK��[�����Y����i�{�f��[w�'�Q>Y]�R#a����2Y+w���ifdr��Mj�-����2�"��eY�I��Ȃ'��WD�YQ��l7>�ߙ�~%���N��Ӻ��RGm��f����:��A"o6 =��4���8Iىy�]�����Dv�;��t�H��UO��y�,���k`�\cGBA�fu=�o<�T�0KLl��.�;mfгԫN�]1m�HX�5"&�#E�Yg-A�%s��n�}�ؗ>(��&$Zy���]���T�4�!U(u�^�+��Ӹ����U�h��]U�'ę����Qܬ%�O�r��>�?Ja"��n��[�
'f�`KD�fֶU�IXWY���fM�a���X�������I�K�ћ�y q�`A��Q\�5��\�k��� ��E�9����L������N��hA(4�|\]ѩ���˭�x�Sy�(���Yr���]��W�`K��f@�w,�4�؂I��4�	*٪��w��挀I �V8�F�ހ��f�(8/�Y��]�Du� �^��H�*1��{�m�Gc�;��u�T4X����_��pS�%�|x�B�G���x�}��F�����2 �1F�A ��� ��ۛU�Ө���S"$�̙�d>!�tZ"�RN6��SQ�2(�^S��D@��&^�c/"Q�V��R�n���+4b+�� ��{q�+�h��+��P�.��w��;��{|�3k�L�u`[d:��z��ܜ��.��-�|+{��Pq����t��\�	E��p��d��L�CV$���V^���*��08P/��8�)oJs�X!"!c��|5�T�xK{�a�&Ѥz�뜬Guٗ�$8�~ڛ�R{}Ƴ8K/k761�*��=�+*:�g��5�)h�{�5��mJ�fJU�����D���,�1�g.�d�4F�z�����w�ά�0��4�X*qz���7�'c�ZGH���h�<��랣7��:�K�{�f���U���LR!Σy ��I^ͧܺ�]��9ʷi�R���Uz�]8ew�j��i	��ւ��Uf��,�վ�tK̕ʴJث��:wY!�
�C�D��F3H�ĵ�À^��:���9:�@���/�:���5�]̂�]Y�"}2=WJ_"���������A��\���\NN�uWf���4^��L:�EZ��w7uhjGM�إ���ueb�Bޙ|&e���I5�!7v(�(�F���]n�k<ye-�c�lRyg��΍�˳�]�۾�!������z90�r���n�׺����K�,���ua���W7J���V��g/pM!�t���TF�e����'L��81"�������f*!5�}EADDFm�jX�m�TX�E�T�j���T�"d��>^����x���}?���������{$���l<���0�"�Ŋm�����X���.t>�lϗ�=��_O�����{z}�}�UT�EPy��^�H�e**�PX�ł����3������3۬���}>ݛ6l�r}::@N%U��(���蒔j�b�h�QV�")��)����G(QUFT�Q`��b�U�)��Uj���r����Q&�*V�6��PU��\#5���N_���V&�8ёb��E���# FEF"�*
QE�M�KB��!���~�b)լAzb�,TH���cP�X,"��&�9rFb"����`�`��E�$<J��X�UD��U#U@���yjF,�A��SZZ+�O5W��C����F1��	l��#:[b�E��M�4!{�п<����<P�[!��P�٧Ώ 5䅈i���؛j�%�s�E@[+��j�h0Յ$4�1��2YnU�n���I�M�,�S'i�hcD��t�T�6���c��*������Vi0wb�1]��®1����n��F-uڗ#Pxq�6j[��2�C�Av��q���m��@�n�f��MT�Cx��AX�i������hn�(��5�"5iA5׵#,�`ˁV^����.�ı�0�F0/iGGh1M0�vu&�>i����#.��� �G՘�V��DLǷ&��Sjh[AKp�\s���8@%`���4�반܊����`����i�&�L2˝�%�K���h�+2fc���ۀ�Ƥ���M�vl�\�.�m�Yh���m��Ņf�7L�"T�,e\��F�:XS3L�5�
Q%fpTJ[t4����
��[f�y��6Ζ�r��ƓC���Y���(V
�W0I�eD��BU]�WfW1`�5��8v���曬m�/��� ��-����敛JD�����c�\6L�)�BY�����<��ۈ.#�݊�[��1�Ҩ8�İ�y��:�`in˅���9�&�0�5���[un!k[��˪<��ila)`�Sa��խ���uF��
^-��<�Q�v���@�[���M�BMN	6m1B�����F)+X!T6�%n)&�ի�f	ll"ؖ]�)�0�"�c1�m1"[0U����v�VYV���8�"GKi��(1Ж�ۦ�d+ucW�rZ���غZ$!,sJK ��\D@:6G�b6���y�;cMB��f�������JM�U��U�K5�U�JKt5��(��R��d�q�,%�hT��r^!�M�-f�S2� f���3���P�U��]P\cg)%�v��e�N�	X��cL�ƀڒ�Q�#5lq�6�K&�ʹc�Aie��Ii��)�V�s�V�bS`zŸ����-;�1+m.^:�C�Ye.�c1u˽N���y,�.HGK�VS8S\kk`�[�E�-�lv&����%�)M���U.R��e�9���c�/m�����n�si���r���1y��l4R�bkj��@`�u�����Mf�c���[��%,t�4fe��:�&ư�1A�ꌹ��.*�c].�X۲��0q�GK�t���Zu���l و2��en�5�[���J�X�L8!lYD�n:b�j��1��akyvuc�n�훴�HSZ��kWGBe� ��1+7xs�0N�;�~i�nz�A��x���\���S�����	�ʮV��H0K�7U����_�ąɑ���Y3��h�s@3����@,�?|spl���u���m�E��)<3;�ߒ7�� ���:،�桏6���c�J�ւN�sǉ0)O&fA�g�Fr�l��C���7�� ��@�n7�eY�����[t�It�`%%�K8y�긂H��;�����;t���Bg�����D|	��ˤ2��]S�߱)6��teպ+�4fV[��\�A�be,������ū����i���=�f��u��{:������P7�嵖�M���kA ���쎢ͬ����X�k��ٖ�^�II��f�N*]>
]s����,�hX�o��Ǚuw��dnu�9�=��QI,��f��w ����ў[�]\qDA�'�OT��|��|��o��I������X�o]KC�/tt�1r���fED��86���|iRCt8��ئ���?�E�tA5�ܤ\;���w5:b�g� �_[� ���s��H���3�2#Ht�h8��5E��A`�<�;5� �H<f��5Ȣ_'\-�f�q �}����j[� �N�"����RhQ���SL`tLh���
:�Af6p4�2l�9�3�U�~����x3�~���dI'� �	�N�I+����	"߮ ��#ENvbK�����n��&:�Lm�)�{Ȁ	��A��^���ӏϛ'�S�Ɏ��S�w���k��E��0�0g�Zm�C*J���Dn!�ݑ��ծ���˫m����S/9-�+��s�׍.�]7�H
#)�L����>�|C��'�� y����i�� ����%������v`�"�A�]w&�#V�U�ǌm؂I9-ܽ�ъ1�ެQ�(j��A�P#�+�]39p�p�x�j�Zޏ>$�v<��Nݎ���3��q ���j �wgDZ%�9uM�"�x���ds�\��9˪X�1�SA.�Z�����[Z�cD&B%���Af$�g�q���A#a^���H�;s�z�a���&b�7���@>9qxF�u�Pr�Y�̴�Dx��b�pX�e�b	o$}p��@�z� 
�8u�K�u���x�����TwU�1$r5x�~H�cw1��$������;s�<O�6��]�t���Û)X]���z�y�_+��w����'���Q�nm��{��K�ݛo��f[$<m������T�qFL-T��J�BS��{_]<������k{b���bjD�N8x	1,�v��|�L�0rY�S;�Q ��@�O?m��Nt���ӊ��x� ��箋�V^M�'��Ϻ��x���-R��k���6�E��96k�Ss�8��و�^�~?�v)K7����K��7m�/�h�V���k�%n��|�<�JmD�#�b	�5N���`�<
�M]Kdm�����z�V���a�An�G�Odsߌ��wzl;3�P��{XM0���J�$�p� �.w�@��Y��B�u��wX�ʕ-����DnGO��|�zfpC�`^g�%Q!^���n۪�E���'ē���O��l7r������|���O�n��]�t���c]X����U�9B�4�����N�|I�~�$��w(8�.����Uh�ه2��R��R5��gj��Ew7�k�;�6(Crnw�G,��4�y�f�Q��,G{�f�	 ���W��,`��ra�#-�&�5Wj�v
��̲��+,An+�v �j�\&t���,wWYAԹ�F4,�7YY��K����s1(l�c��x��fd�M�i�$�͚��l��Ը�.�<��%͘PR[S]b��Wq��Vݬ�r�� vBb�&[�¼��+n���ɒ�]I2�Y�d�n�M3
�+�#G����b�İڭڼձ�Q\�vy�����b؀ͱ���X�Ě��hfD)�7�Ƀ�gdV�\� ����t7r���E�F{�8���đt�n-t���L�����35���4� ���&�[y	)�r�.xm�pj�x����`���^���!����W��7H��'":y��%��PHӗ���rIb��T�;ȫz��6(�dǠ��
Y��	�톧�^���=�I.Լ��`S�Z�K;��� ��W:�O��k�ԙ�={�6��l��H��x �z�@$olA{���w�>zY|#��t�6�bD%͘��gAkܥ+��\�z�q�����~�|��;~7��ߕ�w�Jn�1 �^Y��7um�I&��A���߅�~7@V=�*�i��2}�5�~&�-�]f���,J��}Ns�ӸnU3�3�Xb�>�چr�z&�Л�ݷ���
�׮��qj�w 3L3���暲��tIZ�y���/�$�5�y������M{��v�t{ꊷދQ�39!�8!�N4�a�&|�v�E� e]� �����D���P��-~؃�nSpL�b�]�H"�ۉ�{��\@x�� �SQ��A�؃�0bUGj�ۍ���ɪ������J� �p� ���D�;�j3!Ki�	
���$�oDH�~���O����K��Rܸv�6̘6�(llc.-bFٱ�-Q�լ���h�X�<���~JS�!�0/2IŶ�cȒU��'���g�wUD�U$5�g��-,��-� ���H��([��N�.d��<B��Mӷ+��K��	� �gDf����m��A�H~��f]��Y�P*��[� �Aƾ���{��H.L��c��C3��O�������J�"f�����λo��2veK�C��F7���^nvv�ۦ��E�]mB��[�7_ $w���M&A'���b��@/#�L����M�n�Jj�f�*��"���I ���O�����1vR�]Y�H��� ��M��bSb� K����$�{l*_D'4ۑ�}�	i�Ă�n F���T�Lk:���%,�C�N�%�l�bRʸm�v�H��-a�Һ+W6飳����~|	^w$�.NC�|H+n�A$��q����X�"�O=�	W��5������;�Q}���gO��n�|�s�(ƹ~�%p$�=���xh4��͟���ݣ��P��BJb!ge�e8�&\6<���u1m���r�`'�H�0Gq];��)�\+de��&���[Q;���Xx5�H���	���ώ��w���q/�v����ɷ�>)�r�|Y�N^��ϑ�O���=#]��x�D��fKo���7k��뾐�2%�T�>	o���@&���x�9��_w�/b��KvBz�])��鿸��;��ͦ��3���pߡ����^�n��	��3�X,����1XKS:KiQ�h��a����_R�|��� {/{��O�-&w���Q&g[��:��y)����FN,bjc�	�z}0I>���}����]ښrc3v��$�'wI��`�]�f��72�d���HKŮ��j.3I���s׷�X�L�<;�O����D���^�[�ߟ7'
����NN��D�=��#b�h+��!���7��uLS>�-�Jʸ$k�q�>��'����]t��õ�ˁ)��� ^D�AfύP�"r�y�I5)ŵ
`�4�>Y>$K�r�@;���$��\�ÆuQ!QƊ7d���u���_�M�!��,�Cw� I~�퍛�E��o7�}��T�QQ�U���vrrT�7{qq�C�t驍ݭ}9G���k=�'ƫy�A~Έ�MO�͆���!�lFz�g�v�,��>��w>�2C��H��XL��A���"����=�xw{5p����.o�]vQ5b����{�a�"$������0����V:�]����U
h`��/-]2��Y�2��4���[��`�&5B���M&ʄ�L-��6�39�TL��Ql�&jK��]tZ��ccS�̹�֖��B��m��d	BQ!I���Yv�r;��&�@���PI�KR����2��u6)ɮ�ef$����M�jc�Bd�t��)�e�D�eT���ha��,5��ģ��Z���̨ǲgf��(�h����kMGmB�;c!�}�&w���\"������L�/:s���c��n���W�1n� O�%^��*@��i�f��y߅����&�zb��؀H���	�� ��޾�,ݒ��[7~����p�*�t��ɸ��H��E�;�Yp��A w�-/4��ڵ�����/��lw,����ތ �x��	��p�`�f�X�6�����3���������t�"��O�cry\��n�]hp܃��k�^�|و<�&��	�n��b����1%P�9by�	��A'��Y�p�dm�X벘���An�ƶ�Ta.6Ь���C�o7I��I�]Q�������Sw!r�U�ޤu�DA&�zrn�v���R"��g�񕯐�)��'R�nt*�m6�w�:�}	��"5gf� gWk����s�M�wB!9ȩwQ!��T0�!b>��4O/>=�I�6�H�N�u�1��̞&��9���?d_O��L� �~h�
m��h���ͶO� �їZ��Q�/��c���'�� NO?'�����!������]c�Y�Xb���� A� ��Y>��o��q0o�4UMtAtgB,���/#�Y��]��4/ ����GG�{Q��x� ��Y��"gD\���_��F/��1�� ��At��������V�V�Җ�2��˭�r0�N���o�yg�砅�< �fq���9}� ��N���6��Z� @=���6�gS�Ӥ��&����O���b���y�L�k�z$�l���u�@�D�Sf\s;�4!;��w����l�t��'/���>�|�
��:���W�"�����MfskpZ�4�&衤H%C�%V�OUw�༧b+m1��.EU�`�J��=�������z��ŮZ"�tT,��O���atE��z�A[��+Η�����N�gf��c~�;zs[t��y��,V3:��,P̼HfyYُ'[�gU�VnU��n'HҴ�<7O�'-T$P�� �ӻh�ۊ�`�7*94"��L\�m �̸&�S4!�7c��Qy�Ul�v]9����zQ�����keø8F����.����8w�Vɢb���`i���U���Ԋ\���f��"�qu��PZCz�d��_>�Agi�ͬ�z�f���z�Ę4W$��>�ѝ������t�i�}�vSݩ�|t2hM����,�7u�v�.�
��LGg:y�ծƞ�l .����Do�'��5���U|B���Rݣ6��j��^\�����I��P���ce`��6ٻ̩R�:�f�]U�B�fp�7%�6�{״�N���e��!�Q6����j �VU���2>�b�gȖn�V��th��z�R]^��m�#���ͽ!p�����*���+�4�oǈS��]����c,�N�$�Σ2ew����}(ff�[<�����-K�~)i��
��.��*�k7F��x7�/ <��S.WG.u���]ن��'��85��ͦ���e�����%r���v����^1�=�x�����UC֫�M�������1��N0�)�Vk�Py`�jwwi�@�y�O����c�|jE��E�}T��N��ǌ9�a��ی:a�t�|�7.��wd*6���%r�DET��$PO9���9DLG���3���oo�ۯ��f͝O�]t�*N�`�{���7�J��ĸ���P��8�UW9�)�7���f{u���/��ٳf͝O�]v�J�(�N�
�U�FЬS�`�0F��`�UL�M�������z{}>�|>�������MEKB��mU��X6�$�@Y��T�R)��+ƱV(�B�.G)�J��p��ih���R��`Q"���	maąENZ)a�l�c����ADDb"����h���k(�9EPh��0R
���J�ED���VcZ��ۂ,X�dPr��(��TR�b(�AۙE���2�ʣ�Qy�1
�(�ۘv&(��D���C��Q���R��	�r��ޚ1CP�_�ƍh��֛h��r������>��X�%�����H$t���� ���L��3;�fx@�Wn�F�����>)�� @�/�� �{�){�e_���'��u���C�����Q �H�>(WS��]��l��z1�A��v��������eT+)�ɤt	e�3Zj������\�c.�-��]���vXJb�޾��b,���/OTѫ��m��I\oD�$Mۓ�͐.��ǈ5Y� >O)�r�3��R�t�H�,�Z�w���z����G��^dG�"c���-��L[�'ê�y1.��A9-�R�=9䊌��8;���r:\�d�@��I�%�s��gN�8y�fy�޶�\��3䊺���I(6�tt�Z}فyl��u0k�nU҆{��V�PH�Tt�у����k!J�,�������t��i�t@v�_O��>5��̜~��?�#���w�0Vq�+?[�"�/���Л5߀�����/��n�NfQ/����c������y�Ns�b=V	o\A>'�b�q)m� �No^7t�IP�P
<���q-�mF�b;d�	�]0�qZ��EuTFn�� ��HS/��3��+�݊Č��P��<���W\G���� _,�$��9D��=���w�,����5Ǝ��	 tvD�D�������L�[���'�r�3��B�`����� �>gf��To�������o$t��y��73��t]�	�e��nz�ղR�kפK�@�|H�m�����X����SG�����������Ѫ[�^J���՚���͑�_
�9淈�I�l�~2N��u%��{R��U�]Ki�aR�F#��^˕E���(]}�����1r�Ze+l�lQ�W�!�W�Y�/�\����'�=_��lCB���E����:�!60X���b��V����]�08�R���5�2�1,���8��t^c�n5:��!1J����h�*Y�k8���]�&�[.�v�D6�\<j�D����]�E�MZ��1�P��f
�D��t :��0-�Y�E�6�K�q��D[iaԷ2�gMm	�c��=v2n6@+�!�C7MX�-e�Hbfi���&���!mٸL��[(�EfW2�i�E��S�7�ǿ�.��e�s�߼
x��/$��B#�zK�M���^��S3	=\�&2�E�rX�� Gt��@�i��k�͊l�K�39@'�sy�_�4�9L�\E��~��ס�9H�I7~'Y�Ꮘ��x���n�geS=�	3*����YZ�Æg�J�E�9�BN%�
~�=~HսI�$;_"	 q�Gc���:��� McŦ�w,��93� �IȾ�F`e�5S�o���v�PAِ �s�йe�H'P����DBr��K�ݥbv*�����y��, ��)_χ��;-Ap���i>@bH3�������q��eh��أĒ/� @��,u����w�8�� O9��f!�L-�.f�TWU3�KZ���sG�os�\f����|������|��Y���Ws�u�t��e��U�X���p���>-��אH$���'�j��D��5ӯj<z*�ዠX��މ�ۈ�@��0���x�b��H���n7����@�d�"� ݞ�8���Z�1:�/�Bk�5����M�$�rߢ<I7-ؚl<8���y��	��S���;��N�@z/�q� �}T�\���.̼������0	��wCss3��{p���;8vL�;,0��b(in��[��άn�!-t��K�&������`�K���I잀��Af�St(�������=��!5=����;3�g	9/�U�o@b��-���=����"F��A�#�����P��)�v�3=�Y�\
�+	r��w�43���A��[�A͎�}ILL�h<C�&5�?P��K��}ka>A%O�5���9yG�g)Ӷun��ڵQ��9�7+Tf��o�w@G�z�V�T(�q ������OX�\1t�]�T�S�qa@��3��w�$��qI9*�Am�CI�aI�\Da��c�Iy���x�d����u�{R��v��<n����ъ�,�� ���ي<F_s�����9��xl[p�%�4زh���H�@����]���.�yp�ۛm�kq�r_���，�G�z���j{�M���	���G��B�趤v�T�n����A�]�>��ھN���%����滘�1#���M�{�:[uG���A �gung>e)�Z����γ=���8)�y�wن�D�I5����5��A����k�e7v��MgDA�,W�1v!�$��e�g�M�O��Kƙ\C�͈>X��x'�e�[�R����l�e�4�v]�p�V�|+���VS"�a��3�qt�=9R�ԩ����� �0��Q��EGP�]�tK���^��$���C�v>�I�W�	
�ǂA�G��z"�v�2Bߑ�|yTA2�H)&@N��p�J� 2�RX\`�ڶ,R�ƴ��Yzn�����9,'P4V*�J�o1�R$�u<�����m�%A'�1���F���8r��"h�ӹ�=�޷4��V�ՙ|k���x���8�O��\���N���%�I'=��s G�����Iɕ�v��t�u�@�M�T�n�˻��K8/��R�����Q�`�|�!��f�G�;+y4Q��/���D1Q�T�Zt��C�2:.	>=+22hJ�୨�D�<פH$�0!+yE�R����!����j�	 �B�iN�%؇f!��D�5�t��d��+�\w�|�0w(�����co�&{���GĎg��O�-��'%�]6�J�P!��IQ�m]��Ckk�q�,\CY�2��x��h�@umu�\�r��x�9��ش�ư)��&e����tp�W32���cЄ��Gu�<AG�I�b\k����ك4���%;8����JșU[G\Ӊ��$��0����4s�Dv&�X��u��f�,�1�\��bK,��s���hQ)n� �v۞6�-�12YM̱��&t.��he\�Y��g�N��;�.��E��ӝq$�{s�-�^�g�+M��>R�~���"��0k���b���Gb��%������22޿<�H�:�"%/��A�V�
�E�kI3H�;8g�'!��� ��n��`K,��mېI'o�� d��	��u9.�`C��U�]��*^,x{X��޸A$�b�A��ʓ��|^Ј1uq
���wIܖp^�����@i����z�g��ڭ.���Ď���@�.�$�Fm�Ak�5�4�1\�8.�,SM�V��Dd��m�)�а�Ml5��Q��ϟ��h3;���m@��Y��ߗ��vtA�����q�
�	-��@���S��p����q8��"��y��J���fB�dT#+6kv������l`�_m��^�(��؃������������3*,b����8ȷ�`xW{����$���m��&�!F�.Н����0��n���~pX;'P*�2�B]� _��>6�bR^�h��$�d��#�v�D|�:�볆p桜D���Q5y����Cʮ�ċ�\g�sz�o1�m�5cU�¼H������Np�?����O���鈮��k�)�j�>�n���y��lA$�=r��g�g���������γ#0��*�A�Q"9F�U���Y��q���ia����I`�>�߾�E��o���אU� �A7�1 ����CPl�q\�p�O���3s&D4A�؈ ؚ������˜n<I>�� ��Ɏ?S�9�����7�l��Jp�2.w�UY�H'�;&��9ػpSl���E�eU���v��l��k<7�����tl�:05H��w=�\6�B���0ӭ����
)����m!�{y_  ߊ��o�#м�^��N�� ���g��y�3~�&K1S�/ �b^8��v[yu�˴�vWI����[	�\�s��w"����3f6�*W\�f���d[���Z��5���o@�m�D�S��x]��^3��]���i�a�L���%�,s�Vŵ̱�Gj�īfI�����ϋV:���Q�I ����	'���:����Y�� ����#[w7��wwI;��4��LC�|~r����k��Y�H�؋��ܠ��J�7ɽ���\+�*��LY�� w�ʷ�A ���h\�ܺ�)[\D-.��PO�&�`N�1p��
�]};�]�d^�.�>�k� ����!��;��q��W]��T�/O�&v�7z&Ŏ᷻��>a�e�>��U�e�=�5쬍͜G!4�:�p�Ç�0�S��h�U"0I��F���Ovc�.'eZ��!��_DG�� ������U�;�ӽ7S9��i�5�[�.�e.)q�	�&�Z�m���D�)uL�95�������ߵb�?�C���h�\>$odG���UcV*�����3v�L�F;�E8v8f�Ϸ�"<G&�/�����x �|H�7��{�"z�lЇ�̅{[M��;����y�k�Ms�r��x$o�˽Lk�3Ae�g�%�WwL@���B��t?�L�aWMU��z�O��Ur���;ב�EoNwtJl�0�4��yB��΂fNg�U��"|g��/�dB�޽���A�$�v�@A$���7�!�l	�	��5�7q*by'�6 3ڻ9V��˚���E]i|�6����W=v]��{7&�7.� ���W[�ǂ�o@Z�Z(�v���adV��N�\�G�oAA1��Q
�]�}w��j�]�}z�m�;Ϯ�Y�y��v�L�NC�Rbw\��\���<9��=���_X.��3�&.˭K�bG9衫�nfri��Q�sk]��9rz�q八 P�ے�B�e+��,�"�5^�V^�s�n.�غ����;�w%@2��;ھ��$��U\����xc�΁x�zo48�R�fL�{+�ۡ�mֳs3+��J` q�J����A��˔� 
��쐮/��ɕ���19vw5�//3,Q���
��O3[��js�o�{Nm��ُo+�fЕƤay�g5%,��A�^��77I�t�]]�G:��;��`����q�I��S��m�X��b%�;{bɬ��(G|�J��DX4Fgufa�L����EN��鱵!ݼ3��=0x���Qy��3o9�#h{*���	2�uć�V>�
���7"��Ҭ��N-__vul��hf��ҕ�w_p,�W[�v���z`S�n�C�gm�\��b�Y���)�����n��Ý�I�kd`�;��S� 3���z�}O�LF�>�&'��Oun�3H���r���2�V�hws�����k�O��e�X�˥Sړ4�"�yS#6��t�_e��د��^�2gm̼�;..��቏n5�%`T��.f�Y�E*J�PV���E#,�$�=>�����g����O�f͛6u8N1gIR�uJEEHt���g�1wlP@P��o���}�>���u�����|>�j������,��g��VI�
��� �d��p�ܸ�u�>�l�>G�ˮ�������o,+�)�c"2Zмn/(����9��Tb,��m�m��T��Q*lʊ�7q�R���D%�t���-K!m���D�P��%��V6��j�� �����Y��J�X��b�>aSQ`�����,R�Ƶjq�R^P��`�Y�RШ��b�n�2�)�q��*1Y*T2�Z�kD��R�#+1�G-)�\a�0�`-�R�n�**�MH��
-���1X�
��A��V4I��F(��̶���i[h[+��ԨJ�Е޻oC�ܮ�|�浨۴�i{j��g1�0�Ƙ��	T�q4�m�0U�[�c5f��Ev�l��IR�)l�ڥ�.�8��� ��4��m���56��t5���bfR]ts4١0)&��]+�m���s����P���B��m��R��"\���6�%\��M����0�a��3�pٻd;2͡�k7h��,ܩ���F�n`705v�m��4shݍu��K�Ћ+�[�"�Z�r�-Pf+!]H�7[��JË�9f,�e�KZB\J���]1 ����F��!�2����Jնٛ�k��-��7H�6�h�30km hҒ����qJ�ы�K�͋K1K����345/
�kbі\4tZ��Y��]t�r�B4����KI���fҹ�a0�ii�7da��p�۵����:-�H��L�VW@����Z$!�ݭ(��e���i0��lWm����+vm�չꚥm+����0�`��ÖX�ɘlM6�Z`�Y���&!�i2f*ѱ�Z3M.����M2S$��K�MF���2���	���ve��a��Eh�j�:\ut�V]�ٍ�Cs2ˋ&X���sm�T�5�("KD�ջh..Z�J�PIt�4
�����Utr���,6;"B�B�j�Ԍke�j[�T��֙eΆ3�)N�8k����k�Х�8L�m�Fh�*Y�� �k�v)���3D2��J���f�b��,�	�]*��`]0Y����V�׎(i�F4MJ;3�Jeu� ��Ѹ�@�D�YR��M��a�[��Z�K�#�m-�հ�P*��p�%��B����C]��Y��P�:�tY��M��yf�Wk��+w+���L�֗7R��v�\%ԕk(C��`Z��e�ᤖ�%ll6Ζ�)sN(�+���k2P�u&���j�̦Z�ˊ����!���:��6(��.�n*���\�@`]R�i,X11��u��Dw@�kjUiFj���#�&��-��KZy�&`����@�V1�%�Gi��hYa�Ci.,�1�'m̽]A�df�ث���\ƒ2�t�ʘ	�(F#*�m�b��`A��P\�]���b2�u-c�LF��.�k�X
��`�¬�5�T.�ŉx�m��ł)k��F�&��.h�!+Vm�Q�z�5/�����a�]t!-��)tfM۔+QYewR��q[��cu��F�M�����h��֓C'f�ss�0،P���Mp,�V������8�ȹ,Jt��ߏ�w�$��< A7�H�l#F�Ϭ��Zo���;��s[l&��ͪ?�^���d�q��z`���l�>3�_DG����G�͈U�̎,򡫉y��\>���wM��t)Һʬ��˿@P��n� �?8:�����l��$��wfG�����i6Il� ���+��SL�f����0���/ �� H�n�g�s��Ώ5�@�d#�K�dK?�@��Ӑ|	 ̬���;Fm��8]+���Լx�:�#��$6�y@=M�3��z�X�,Jб���bcG��ް�V���F�U1
ʒ���qEm$��_gm/�4AIҤ�\��/-�x���:����s��q�'ё[�IWDAգ�V���*�<v�<��t��i�ً.��6ƨ�>dăe*J[k��оT�md�ڎn�uD�ZE�Y4r��e;X8�67r��5H"���F?�H}y�<���g�A�x���}�(¹� ��N|�h�A����{�A>��_�J^-YIg�y|g� G�Wr�m�1݃��t)R�Oߦ=i�
X�8 ��X����A n�C�'MM�n�b,0;U1�v�.vI�Iܖ�T��9�$�?<p���s�����O�[�{��Ta�^c�@��^.��wp��Y\]5m���J��F�V[�ʕ��U�P1��jmmEUZũ�f�u8Y1��̏1$$�� m����8�y�#�+�A*�����L�8p��T&�b�Λ�Ew3�6�� �:Z�z;�" ���T�5m���+;�T��LRb�3㘢�1'�{1�T���S����)u��¸{�L��}g��I�n�P�#��n}Sf�؜D�;�.��[]nQu--��R�h&�N062�WJr�69i4��ᩝ�ă��x�{� E>m%z����v��%��V�Q��y�f�g�^r�a�3��ȀW�&���4�XX�Z�A���t��fv0h$����ވ>�{b=ދWOB�e����6��A9Y� /�Z���O����� �fpA���M3)b��A�6��-����a��
L�����}m���7��SI�<�MVs�$�@/�U]�yߦ���a��s6 ���L�)�9.]L�j�������s�]��;�9!��/&�ހ"+�x�maVhn�r�Է�A#:{X�vE'�UMtD Oy q� �h�8���닖Ʀ�:=}��f��A��B�.d�x��[��Q��'���� ���H$b��� ���oYA��As�6n�UeY,�3p����k�-��t����܅^v�u���PX�!��pXJ�,�ow����qj��t��Æv�+������$��Xz;sr}V+�s�DM��'T�4r)�L8�4��1wN��c�\]5 n�����B#q(&j��&V�!�q����?/���&v0hof���D�=Ǡ�yOs	�2�E�p�� W��܏F��A�Ӷ��\"�f�Y��l�3.�����H$�?D%ɻ�=�@�1q�sU=qT��0&��-$���eު�b ��� �k0w4U���D����!]\�K��,��0IÇy�P�ػ��cY��V�OmP7�$Z��H'�ݐ�r��Ȏq�	)�"��o��N�$�3y�r�(�\8ϐ\ُ�OrZ��:�F��ήx$�+	�9����x�f؊Gݱ�7�0�i�od��X?f݊y��k.�G��;u/,�G,-�vw��U����®7�2N�&�*@�Hw��Ia" �;�8rJ$0�[���JF��z���6��@�a�,� ���^��^,K�YW�+u��`�!�Ωj��w:�\J�]Ύ���@�	��[M��f��%�!v�GZ��Fؚ��6���quDs�[��fb��N�V�CCH
����cm��nŅ��65��iD&�Ο�|�i�7,Ґ)�t4c�D�Y]��:���n���hp�f��B�F���͡��M�1���Յ���s�ۮ�� �߅��U�ۡ�� ��G��h�t%y���w��6TF�/�����V4�K������3�!�@�nc��A>16����-�1A �*� ��؀
��i�R���E���蝋�f��8p�'/ʏgC�M�s�"��E`'C�g�{S۞ �ʶ�	$gv�x���I.�݉v22_��ɼ���B;;�A��	7�yW�a����h&�0�۞\Ig�N3L�u\�ğ����.�tm/�"�� I�~�x�$õ�����)Ӣ�B�kyų\5��Yt-�	Kfѱ�rW@�Ɣ�fg �b��8,vI�t����+�p0i���c�$�Ek�/Ɲ�-��Zy*�wh$oQU���p�]��˘��^ں�����dPem�KD4��ӐC�\9oST����k��g.����3^�/f�k���c�7s;\�������7�H"�: �Ms������K���d㴒5�-���3�!�L����D��O�[����omD����_�1���s��!Æ�8d�B�{U��k}s�I;�� =���:(�YP5$e�ZIw�K���*6DOJ�T��*6NY$O<��%�� [�/���[���|g�B�ZI�$�vw��)�֝rB,��Gi�M�a��r9�KTC~��1��9d��7w�j�$�Ǹ	$�r�R�c�4(� n�x��1�������;�%�:�U�ڧ!�P���f��|���x�<H�m�����3���o���c]��ڢ��[ăr��rz���P�[��_),T�6Vt���d3n��	���k�����\Ii�ҡ,}f��_j瘎0���uک/6mʔ�������H,������3�-�1��\3�C1��Qb��lF�{;O� $�� �F�dJ��$�[U�Aj�� ku30��pC�3��a�U��~[|&��P̼ȀO���B	��=}����zPb�`��,�,Y����Ԇ�uMX$�����ax��1ȣK�'����,0;�vE��Θ��@#ӭ�y��D�dG�t�_��s��� �7T�`��v1�mL�b��4I3뻇���0͵��s�|r��g�)�<I(��+ѽ� �m\�k$nge��ۻ61f0f�Uз!�$�^<
����Z�#�hTӊ<|�lG�a�mcYݒN�>D��y'c���h$6q���//w	#�� H;o�V2���Mk�3����}K!u�i��U��G;�{؂�5=o�wh����z"omEw�^>�Ѩ E3`X����VN�q.�u��*ݘ'\��`WGS�$T��Xj��_�*������]��	'76 m�m�\�.F�y32�tK?j˖�b��k�ID5��,6��*�6�*�I�4��`��3��.ֳo8p�:}�Q����y ������s$k��ݭ'|UwtA1y�����;��bA�J5�FZ䪂�W�sz����� �$A�~��뽻N;s�l��N{�ٓ0N;���I=ok���r�1�&+�D�M��̀�0{"��^c4&�d����@�e9�V���˱���NkO&LBv��Y�$�2���t]��{��V	)��W���S[u�,\l���~���i��@2�.fd���U��������t�9�Q�h�.,Z�b4��&s�����Ó(�����߽���CO�+N��9�i��`��4����^�)�eHv�Dh�v#�3�iYSBJ�M�m	��`�QΎK��v
q��F�/g4��4�g0h�ji����5с1,xBZǭ\˒��M���V	��0B�&��mp�{�.�R�."��n@��$r+����*�
a�5g�v�����0/YY�C)�sC�I��R���-��:뱊0���A�G���Ԥr@��cb\�j�h�!�
�`��
bR�"{{W;2/�tC��6�	��ׂA=��F�Z�ؚ�u��:=5O�;s��7���UPK3��`#ⱶ5!7���WV�}�J�<\@$��q�&���}�6��:��T��a��H
	��� �KZ�I��Z�B�����T٤�k_w��i~0e�s[f�ñh~�}�a�M,�0���H#*_�w{#���GUۑs7D��Ml������>5�$��<{���f�}���؀�H�� ���@Ti^��(K)�~U���Jm2@֊9LBʑl�hM��i����:a.��Ѧi���H�(���}C�o����PH��r�{�M58;]N �)� �7)�&/��c<�/d/[�Ǩ�b�r�^+�/�7e��g\ܛx�Q�E�[�j��M;��A���6����GVkȜ����o�!u�5���1�	 ���P	$wvD�j���:�ճ�Ѫ����8h�N�����㝺�I�43H�ް����$�ƞPH;ݏ��t�hr���ɜ�k�x~��gO��M�l@+�u�j32z�Ƃ��PL���Jd��&�U�눀O�e�s>>�U����f���}{O����tW� j�"*�j�x�z��В��cM�fD,e�lv!�ۜJ٘�=z�� k��#��;׿�e�5�B]��߻�'�/q�A>�舅Ϧ�A���ꧣ �ך��I�����.�,�~�]Ὢ��� �M^t$��;x�7k_c����6��'B��tCB�G�P� �rIf�X���JiuQ�3�˙��#QfUղ&�ۓR�"����F�JsVyV�8+e�M:�,�B'�.��v�m�HWM�\"S���)R8��D�1V���,������qH�f>VS�]��r�T�RG��遖��Ӯ���۷}Z/kwJh������fg�љ�y���!��wu Ma*�!��F��[���<�o7�=m�B��Ysoy�ɟ���4� z��D��yj=p-Q��U�J�7��ᓕ�0�w.0b9b��}���n�w�����f��0�gm�%!����!2\�v����eΕ7��p���X+���f�����VT&�YWG,�b�n/��@��Ǳ,흚�c�m�.C�F����a��՚f䷗�1� ��1�}׷ygʓG�y�Y-<-��AY[YYZ�~}e����^�sU����V�;׌����e6�� wn!rg,9�mod���T�}�t�n�I������TtP.��Vx��}[0��)c7g�������]�;�+�Ϋδ�НY�)�g�p���V�-d�&�b��O+u S8
˲wo�*��d��
��>V븳tv��n�][�+�����E�I]�`��b]��wz���$�Ga�n֬w�jȹ�o�\P!pW�� �X�"�]�їY[w]�l6ܷD�23H�TѴ�Ic�̐a<A����e:�up5tվ5#ҳ*�;A�|y��T�jG�Wx��^ejj�8Q����[�Û��U��U����T��Q��s(W"�A���pE�E�5��Tr��<�3�w6tN�s���lٳf��Y���,U����.�\�1T��R�U`����' ��4{u��#���N�s���lٳf͛�U��҈��V�#Eˉbe�K��(ʑh��-8���[;�K�>�:'S���}6lٳf�C��1�%aQQ�ز*��Jֱa��� ���j¢�jZƖR��b�q�)*k.*�=ˌ����̫���Ũ6��(�T�%dFcv�V�uH�[R���ȯe������ʭB���-��&�*

.[+X6֡Kb��ƍ��P�2��e��ڤX`�(��H1�*-b�S�\3R�e�
�q�b!F,��-Ue�.�m�\j�5�PƦ)m`��x�孥IX��X�Z,��������* ���cB�e���̴\ER��%�`�aX�uB���s�z�6g^ �������L�%�4
������s�<����q �;q��I`���_`�mu�.WOox��cʬ\�L�r靍H3�qd�@]o=I����o���>!l��@gSq��\�Ogjz���ZK�|��lmH��^as������p�2ʶ��JO�wQ)�8wb�>�?x�{��DA� �Kq�j:&E�
j�\e$o2b��L�3�&r�OF5�
�
B�Xfk�s�"�+��D�֞B ;Y��^�X�*O��l���w��!�b���I� Kk�3�e�5O��I,������6���yy|�Hw �E8��
Y�]�ckr���Y~$��D?��M�7�{&0�}~�1����4NYcA�'�0K{�I�-�wq�gT�1�t��]���>�*���/8�D�b���6i-��� �x� �L@��y�L�%�4
�gU� ����5�Vn�Ua�����v��}�ψw�5�"��s���~��H
<<��T��6�X�h��X�L�i�CF� ��,͵�3��k�}{�����]3��x��D |H;�v��"y`����[��N �:�)�kZ)g�&��� �#�;;�8���==��0|O��i� oc�$.]�#�}��&�>�(�mS�(����m�8�I��8m\]ꧬ�A�SN��y��	��6ݜ��!��NL�Wx�=���3V� "I nn��:�,UI��T[x�>��� �q���K�S����>1�L�D��@��zl�L�x+H'���`H���-��E-].�Q�l��kjj�⊨U��X� ���0�����7����hԉ�_\Z�}|� Wsa�`x���t!����\ŷ�*��7N�(7��Eh�ޯ{ߞ��#�KjKJCf�H�8�C��������1.ft0k��D���X���!]�qW;96r�+�4p�ܼ�Ek,nkUXf��$���5-wRQ�)����L��$���[X�%S"�L�(r�vZ�)J��Mrq�y�(�6�u��i���4�e!�$P�^e�1�*S^)Lm�6�Bl;��9���ǗqCC�+s2p�s�Asu�6e��|��hD@��5���Wf�֣�E����Ґ�l��1E[���(s��p�I���ׂI���� �t�Sr���V�m`�L	ۑ$z��m33[�L�љ'}��Y/�m����p��g�A ߐ�ޘ$�7��\h.���Ncb)1g�&��{: �MfC�VW۞�}�W�%��lA$WC����kt�Ĕ�pA��'��	ֈ��y�$�l<A��<�ާ�E�|�	�V�@5�h733�(��B��	 �Kt�z�o_jS�#{Č����Έ�gKp�_��?%_a�������y6�m��ԠhW$�&9�\��$˕)p��+T���Y�)�g�׼�%�	���\_�
n��oKq��[5��Ɲq�_�vdϣ���%�9IrZ������8t�Ғ�_���.�7D��*H����P��S5����D�e�r����}f;�jC�dK�
i���+��d���I>������2��-�xl���-W�{�C2j.�vt_�#9��H��@:��i>�I/7H�VG�H8�������A�Y�_��tӢ�a�H$P������̽KAC;��<�3�������8�5ݱ[����G� ��D��,��N���2_2�	7���˩-��g�/���]<�<H^K7��2a����l�c���R%��!è;0؃����1��]� �aCk&I�`�$&�ìu�;��tDUvj"�]<�	"=��W�$�QAc�S�
#(�>=�ω
��1WV�]���A8��ӽ� �ӝL��z$�O8�I��!yp��T"K�z�zjm�!́���1���z�^+�0�S��Hn�|wF٦
5c�r�Lu�]��GƧE�-�5U)�r���PI^�-�Z;�Ƕ�����
 /}���S�� ��=%ovD�.�Bd�ؖ��̃ז���\�f�����I>$f�DA'��C����<.ӡO��8��{�$�û8O1��H금yi����,��S�z�<o��N���tζ���.�?"�qb
H�Y�l�bJ�,90�\�[(͘^�c�;\`����>���.��x��<A�巚��	>�Ȉݮ�9��k2	$vf�GoY�:�3���"$G��i���;�Ո{��v�4�I���[y��b'��U����Ddr�vtK�I��暈�$$3�燀FGl��*�v���~��ϊ��pY�3�<��tN+����x�7�����n*���FT�TT���r�J�I]�^4EP�1�.�O+)�}�[�;5"7��+6�FYSE5��{Q*���4x{���&���fLJ���� �v<L�B���Z$��I��9��@�P�c�!� t�Iq��vA�v�L�E&����M��g1�D�n�˄�ڨ�Z�jp__Wק��3���6�Ky z�c�A'6[�{��nhm�}x+�"<O���p���"8vgg`fI6zq� D�VO8�w��O����#v_�B���af��,�FX�L�҈��#^�����M�	�M�yQ�ݣU�@`p����~1�b��;�]:H'(
��h�m�n�x���(E��w�6��..��)�a��A��4HC��.@~�W���&�q��
�Dˆ�	�وo%){�^�H��ʥKlB�e�Y#{f�d�/�}�$�9��\	���32�oZD-��z;��Q�������㵕�⮧�X�^+Uӷ1X����^_~榅ڡB��9�&��BJ	n$!\L�EL�c)�Lm�ii7e���b휴h*��G\Ժ�K��+e��n��eIj�Ҥ�Bcv�.�2Q�@MHŎ���`��h�k5�s������j*ïkи��Q�4�֋��h��a��Ѻ4i�v�Ґ��&s�[d�f��%M�t��MB2�H�\�����J"��*Z��C9��Ra�����ΓZd���a5�(k��\它h�I�
��Y�k��;:2$F��y��<�>$f�D��_�d�d�Q	#���T�z��L軳��&�][%��z�{d�e�ň �H����3���~ˬ�e����8�L�ٓ�Gr�!
�A�;��<
�n�@�S��-��/��	'7� ͣLt�w
^��H���&5��U)������ ��� ��8~}B����*=7ɰC-$������H��UD����Y}���7A!Kn( �w}	=�!o?	"9�r���%D�x�wAû�d�y��{YR�C�M^�Ms��`.l`)�`�����!r��&��,���I�ڽq���s��=�rQ�oS�ƻP	=݌��T8C35�H���c��~9E�����4�d���-�P�\�˔��oet5�^��Y����Y�'�YM���8A'�3JcV%]�X]%������ns	3ݎ �ݱ L=�\DG]hg������I��bS:,��<
��v �A긏Ao$v�PתqRx����
K����N��xE��w)غr[� ������Y��#�	�s."������
�a�nA#�n �y�U.��<)5�2�!p�$m�c.3Hd�Oxo:��y\@� ��P
��.<|��Ul+52��
�rCj�<�6��cMcIm&Y��J��G�L%!�Ͻ��~IA3��$	�m��Paz�7��:�b	$x�l<m�^,$!�Yݜ��4o`�S��Ǻ���{�L�m���'Ď͘�g��7r�k�<V��3��=���%�Z�!��~����� ��i���f�Xh�j�<�ȣ���RZ�8��i��b��+�E���7YF�ق����7�w]s+f�.���㨌�J���w��b��I9y �1���j�ۥ�l�t]����^�i�l�y�۔�x�$������v�='�}���+��~؊���Pvr�;�&�;��L���1���4�"c� O�B�ߏ�;� �dUc�݇�tN��)�3 C513��M�h���X�D��Ճ�j֓:����Oq�3�~�
ܺ�<t�3l"7� �p�f�̳R��GFH�y���!�)N3�N��PN UxwU�^V�!�:�S��O�?6��w˺ �q�&WCJ��Ⱦ��;:�yr��䦁Tf����1�a<$��5H�x��syA[� �v8S$��wgG�T��bB�o�̣h��l"���$�ݵ�q��'�o�WH���G`�f/���'��ٻ8��%`;��]��J��/6���˳�|���n��k�Κ^Z%�K���^<H���'��Zwd]�;�N�38��H$:��;�����[`�Ϧ	'��#�|����p"^�J,g��*��B�&�E��,Mf�AD��K, Y�!���w����8N��Mp'���I �o=DW�y����\.��x��ǀcʨ�AJ��\��h�4I:'�N���R�����ǀH#�f= �Q�-��Z8�7���c�ggf('>؞�A��q jg�17�
�g��8F�c�A�/-瘂�!>\];�9)�LO7[ff�sE �g��>7]/�}����5o\��w�=��c�p�I�;�� 
�-�	��	FR�4�]��/t5@���G��=�����������*�����Q�|���n(��DP~�0��� C�΍�H	�@�@B+@��2������ @�0 � 0@ʫJ H@ J2�2��*���4ȫ!**��*� �B��}��"+�(pL��Q9� )��
&gc�C���Q!:�����!*�J�B�0� !*H �(�J�q����PB�B�B�H�B+@�B���*�*�*���*�*�
�pEx!�@�B�H�H+@ Bq�W���+H�H�H+P����"�� !(�!�!"�!*�
�����"�!
�!
�!(�!"�!*�!*��
���@�@�0*�!�!B�@�H�@��� B 1"��0 !"@ B�1*�42���2 ���42*�CC�4 ���Aߘ8w}��D�AFdI���{���y��P}���s���c�y�?���������z0�/��9ϴ�?��>��S���(�������Ј ��G�EQEb��X�P���2�Oԟ�_���?b�UE����|_���'=�����?3���D� s�����p�}�@YQ`!E�EXd��VXEa�VAXeE��V`%���VEfAX	Qd�VdU�AX%E�X!U�e�VBTX`U�TY	E`Ed$�@H!@��$$V@�a	V �%HYP 	F����$eF��%!	@��!��T"V@���"P&�B�A
�@�AR�TV�EhAV�V�V$U�JEZX��hUfAZAY� �bX!U�Y�V!�UY%�d�VYa�VREXa�e�VO�8��EfAX$U័8\��~l>��j*��*�P!B"�""_�����??���AA��>�����?������UW�~������W���ǡ?_i�?x�������?�}h�(�a�!���s�N� TW�EQE~�ԇ�ç����'����
/_P~A�a�������~����=hP��0_��4�0��vS��8ATQZ>��~�/����_�*�+�����p>���o���?i��Zp~�>BO�~`���<QE{}���J*�+��A��;C������Np�~��>�������$��t�������|�zq��_�0>������)�����_��Ƕx� ��W�|}~�~@�b��d�Mg����Qf�A@��̟\�x��
�PP�EDH�U �!U*@	G@ Q@�@U�UR��PUP
PH6ԡD�TP�  �"J�	Tu[f֭3L��AD�I"}2��*�X�j�@�����АQU'FR�lB��PB(��=�                                             IKޯ�F>�V��)�4;ۧ� f =ا&�F��5�����cY��5�x� 3�1���'��
����@�ӓ�����m� ��2e]>
x�z���{X9ڔ�4�y�� y�R��0g�@�w
S�҇"�.����R/yU�J��\   �        ��Yj�X����Ҫ�B�{:^fER�{�� �PUY�BUHSu��s=o\�B��� 	�]y��.`u�'�v�@�7�   &��0C zR�� �;[���j�=�B�z�u^��͇�׀ �ĵ��q��ޝi�국���Ժ��o8��j�%EWmB!/�  �        ��ﰼ۵�UW�d�=����\�Z�.Ѹ :���뷳�����Cj��{l���vQv�\ �����u)�{�z�
քT�   ���>���ܺ��;� t(��)�=����^n�����aJ�� ;f��˦������wm^a��Ms�[O!�ZuԐ+|  �        ���O&�mRs����i�n�����/Jz���>��= ���Η��S�ӷ�ǽ�n��^w��](׼ޢ��7J��R�%8π ��o��-^{Ρ� ۶�����n�j�OW�n�m�uw�7t��D��x ��{��C����S٥yxY�l��bJ��/� �        ��S1�|� ���ͳ˻���p 9Ӷ���ngN6!�94��� ����7a마=�%IR��  �}> }x�.�S� 4t9���\��`�  E�.`둮 z{̼�]Q�S�h)*Pa2 S���@  T�1���  D�*���  ��T�����T�@h2d0�J5)H�����C�� �_��g����_��4��\�^\� IO�Ls�`IL�B!!� IO�H@�XB�		~�?���?^jk�bṻF�˩���܂�&%1�e�N���˴:�n�5V����IK��a9z;&V�]��	הH[��G��EwJ��/N�=�e�*agFK^of�12}Wk_Spq-;�~}[rp�r�{~�3��H�b�m�LzbS�A��_&#fA�vl���������m����`��b�%qoBzfU�����"��^pեM���)פ�~g�I�rĻ�=�WmՋ�ỉX�Z'WȦ��wl\N��,�Q�Bf�jN8��1Y%NR��
殕��ڄe�+L�׋LG���,�8��c��Gh�I:�fr�	#����v
�c��zb�h�s��pu���rup���x�4����_��I�i�-�L�S��GT+4�wp�F��5U>-ϗv�2a�cMa RJ��!���c:��*v@5��d7�(n�$��y�ť�;��c-����h�#��̑�^���0����V�H�o��k1g*l_YQ%��T�2]��V��X#�9�厇�=�~:��oE���+t3:�;�X)r�8���I ���v#��%���]���L�ScrP%��a`�΀N�G��H�KN	�>���xn<Q8 3_r�S(�a�v&�r!f�[nP� EOq�cd��P��������e�!,S�~I��b�dk("��!n�؊�mpX&n��9�l�	֫���؞s�����Ң-��	�.��HlK$�Ż��$=z�~�cJK��ܯoZ^�
�k�0�S�F�dHZxw�ܝ91�6��D[�^�y:H�xk�35]F<B!������|�]Ñ�F�����ִo�c:��(,b�f�gp�����c��U]١-Nw�?o<�kQ��{�]�T
L�/���z�]͝�q��ޅ^�<}Ҧ&��8�$Y��Nk�&�� ޥ��؆�Dn�:�D����NȺ��Ǻ��Yx;q�\����z�i�����L8)��Xe�h��*�'�f��^n��=�h�{sln�"ν��nC�k�fL�6Tn�eH�O��]�M]�
�{�6qf�+c3��,e@gΘ��7S�*`���ݤ�	vD9Y����Y"��n�:�]BB����c�J� ����?T�[ˉ��Q�_�V�V�^��:	R��Gj�Hp�Z���C��Α١N�5�9�cB�ƣ��%9hɋ��Z�pA�D�V�x\�2ὁ��%۲���⻼,�^�p�d��@X��u&�k����p��փ[͝ɬ��W�m$�3�������Vؠ��U�f�Lt�(�-맳Z8�մ!�,�z[{�j��60�(�;��l�Vo˰`���(5���H;{4dI��.���3�9͙�s���'ێ@�]eij^$��M���w�Rhne��o�l'.6]�a�������u����邫r�֚q�à�x����n����ɩ82�+6e�y&,Od!�#��h����ÎkūhI��3K��}����\&'��3,��H��c�о��$Z�>�e�S]��=E�1�m���H���P˔o<�$ߦ,1��8vu�� l���"��o��#v-Yٗuk�w� ��/3��t̍l� �w�Ij�]X��˃�(5�¨nZ���*�a�G�M.�`�Rn)f�`ѭ�M"s1�K2�t�hk7���7�`���se�8,3/��R5��COB����!���Վe�����T�����N:�e.x�X�a�J�NG�^YX�T3p���y�w-��j��&�	oG{z� �B��Zh��;g)Hĉ\b�ƚ��:�l�ּ��K��ymj����^d;Z�)ٚuc�i'U@�j�W���z�J����J����Aܹ�τY��Vѽ>Dv`� �YRҵB�j^}�u".Z�9�h,h2����/0d;��d�Bl������V�Qj�
;*�րlX�"�B�j�y&�ֶV�n]��j}5y�tށ
�m�ш�t�w�36;�l�-}WaKc�(ȵF��F�-�9���6\�^�|8c�mhw�ٍɷ�{�c H5���vݻ��Y�#��&�:3l�b��-�q�9Oz��:�Y5�#��<���I�65�h�����q�C�eg/Uu��R$Z���55:
)��ݚ��U��7N�#Zv� �����LY׶�h�T�ޚaԒ�����S�Z:�|ؼ�*�Z�ψ�T�*��I�-Y�w�1�aR��".���PìDL�V:\�h/�#�s�:������I���9>�'�T:ɚ������4��D��R�s%�I�v�ZrB�B�5R�x�5���jͬm픙��);�"y2� F�e*�k�z����q��G����Y��LuR�5V��}�3P9��pù�5�(`�%�;��P�m�fYN�E�u�`n�R��kn:Z7(/)Qa�c�^�(�u��D�/�lMI{�7_+L7?h�][�f���.`��r+�i�?9C���N�<����������e\�qCL:�0XlV{��D%s�����J���;TDoaNv\����O#x�j�mp�s38�ű-�S�DG��%��Q�%����Ga���en��	��9wKY�U�,�����x�T����.Q;�Z�-0ѻ����B.Z���իpM�F��xD�M&��("��K]й;��Xl�SzH�p���Pۛ���Ӊm��`s*G=��pYb�kvdfCr�Cn��;��L1OA��Z3J��1m��50ǏuR�95:r���M���`�Ɔ�,oGvf-��Ӈ�L���
�v�&��7�D���)}��g��g>X����6��%�i;wQ�Z�w�W���5:z�Dk��v�ٸ4h��Ek�6�/�N��h�LZ�����M=&����w3������޼4n�͸��g!�H$M�'3�����-�3�,Uϋ[�FrU�CQ�tSi�j���șɶX0,�&�A�&�r>ۺxM)�ޡuR�9����,�5�+9�K��4w�t����.��1nr�N��:{`ը���ö�'Yo5zr�a,����v�יy��!*Vv5����ޛx�A�I�f�&��,��c͙	����x<쌓����n�M�{��������?I/l�sf`Y��J#^�k���ɖ2��uVC��D��C5+A�����Ytn[���$���z�"t�ɒr*��G,��1��rA�������p�8�����u��4sG���NF�2�."�F4]3�H�njD��	�䀈�Mli�ȯ��/Ce�wuo�c���ЇHc�j�ap����ڻ���=p��!�4����r-|��fu����fRiXzޕM�
���w>�X�lf���<���_m�V��M�&�LT%��
($G���1׷pky��Ef�H�p��N�Z8c��]JY�d�R�X}{u�<&�i�8sќ5Ņ��M�u�v�:ď���ҫ��H,k��Z��/0l�x܁b��p�5�ql��/"��JժI�`��CF�l���U�w$?5���L���O.�YR+V0��.�ja�@����t�L�xS��rO�os7����:,R{��*wq/w�#�og\	���-m1p,2������pl9sV%f��U�7)�чN�Ѹu��߷IX�jL̵HfM�6lO�{�B�;���VC�i��c�x#���>�D2�m.��Ald�z��Y®�,�́]���]�+c�'���Ȳ���E�BU)t���i�\�h�2RF47E܍�d�$.�Vjb!SN5��<tJz·�A�OU��ǲX �3��),<�Ƀ{�YY/�5�[`�Z��ORnk�0��fe�����6�L�.I�qX�d��!��S���yU�1��C>�+��>�d�xT8t_lZ�ݥm#w��8y]g�G�t��t�ncF�'N:�ou���7�;�#�N٨������[6T�����hv�)=]��:q�;u�K3I�����=����S;�H7�,ӭVw#:���R�NvnQ���h��V��ٵ�'YstZ�-MRR
��j�4s�WV=��.�9�[w)kW�p�6L�\��_p׍q�	o5X�l�-�����]��&dQ���^^��7��]/ܯn3��/��P�79�s�ђF�G!�n}ܥ�ݽ��e�ۦL�	y$ɬ,��S�YaY��c۬y#gce�y�9cp�N���1��� G135Q��7	"V
�	�$I
su���[��ʹ����x\51���U`��^`�tv���O��{�&`�;��9Mof��C�5��fV:r�������6�l��0�5F�^J`@�T�bup����hbvc	ab��tيq�3���cEJܵ�b�WSb!V��#
�DOL�]�W�53����4�y���n��f;th�fv��E��;a���d�]�(F�ۉ0��R�{��٦��\�܉�������*�q�2�fZ��U;f��v~u�F5d!�c}^$�B0bߦц��R�%�J��j�t��SK0�R����t��	3���7K�P�er�0	n�f4oA���t�WV(֤m����̻s�b�j�͇F�S��5K�:5tWl�!W1M]���"Qv]�,4�Z��������먬#WQ��>�u)EO˚�qV3&.KX�*Cv��͚h����n#j-���Lr2�؄s�fr���p,�8k"J���a8�%{d"o��ܛ�����7�E��JJn���H �mJm�
VP$S����̯3�#�|q�#D�n�o&f�#�g�J�2�IEDe���ܑ.9�j8%�TB�,a����= ��.�K +5�EڀT����sA���'��Y��-��I��؅T�WN���K��T���4�V����,�IttB��a
֖'ٹ��!�J�����܆gW:�
���t�g8�Z�	���NӝD�*+_*���I�otuP�9�+����	C$9���l��fc,r�s��M��M�'s�.��ĉd:1�rBr�Eݘ��W6�ѕ��`F�n��tjZ���SP@vm�����i[�3ZD��Q�u("�>&�'�+&�#b=neN�KC1���l���bj�ZK���&�*[LH7L0h��?h�vv��!3�
�z+�B滹4��.2�<����Ĩj�;$�����zU3�)I�|������[��V}�h/veu�H���錾c�j��M��f��tat�}�Nއt)CVrQ��g.W�KΉ;����n9��Ӻ��"H�[
��bW����/]՜yz1�tP�V{��7���B��p��fZ�D��&����xs�N�w�t�.��;'R�(���_<�1E�H9˂��t��Q�p��gt4�i7Z���$�?,�c�e�ėe��M����;��-����`H��mK��y����*;NPy>�x�4n��qN\0XF�x���2a�9+��PN��5�m8u���۷���X�H�ڠ�1m�u����&�R��J�űR��C$��d�����6vd�&��F���:�d��_*�ɩa:�÷/�O�仮E�&�t��Um�-�ba ��K;���ز�	�A:��I��2�b�F[u7M�Oܷ�0;�l�����4ʕlr�eIltN�wsY;�KxM2�腎W2�׃�� K�E�#���9���xC��?>�;��f�q�2�`&A!x	�	���{��@��W�w��i�٩^�m��;���) ��ʸ��~��[�v͌@�ulk��k�+.�Q�Q]*��e*�RD���ť���������3s�p�L�Xc�ח$�3.����cGO3/"�n�znrè��gݮD�or1O(�-�C�q��۳��M�H)�I��Sm�P�i�RFKiel7d[�{�v�+-�����n�tF�׎��������;K-�k�p�Վ��M�c��q��r�?D�����	�^�ysd��Y�L��d<rg˹�Vp��T��{��Q5b+jTٕ��MeT�|�p�FJ�w���,ꐡ�e�18��5L�n�I���v�c��j�x\�]8$So����yR�F1�Ԟ���;J���"}1�n!a�
ib�@k{Yf���rkP��$	�1)�De��[����"��(�aİ��X(ȄXV��GeVg
u��^�eBK׉N�;��Qͭ���م��5�5��A�l��4'���3�I	��mla���^�8�5�XIf��u�X֡��YGv9�UBf��I��	�5�r-�7�o'Ы�u����3�)����`t>9R��(������ku,8���!��ͭ���Q�;�i����,̄>�wVŚe��5v[�8�e�5�E�i t���:+$���\��	��;-Ӄ�� |��oC��
;�T
��,�(�I	�!ë��'Z�[e��vs|�`z֋���2�D�.Jt�H��!caӟ[��`Q6�jOax<�{(��m�t��g�A�yҥ�xo11N����0֓ $NʕuI�� gv��2VŔ�|�K�;H�ۡY.+d}�%+:�y�k�.3���	�
I@P��*BY$ �� �P	),�BA@*��I (@"�	d�B,$ �A@� �$	X�!!E�)�� BVH	,	@�,��H� �	*T��d�T�! )!a �@XI ,E!!H��B��E�!Y!+	 �I"�E�$��a E$�@P�V%d�$�%B� ,"��Da�J�d�@Y�%`��� X@�
�(@�`@��$"�"�)��P�$�� �"�	 �$ �V@�@���P�P	*@I �`	!H�$�	'�	!I�yz�1������ӆO1�\����5m���������Y�3���M1�l�N��5 ʗݙ;��mJ��aq�h��a��s���N��|z�b��W�������K�R����=�m�U���b�ż�p�:�=DКc3���a}|P&�]�W�z���rN(��:ʽ��X{'A:�y�=(�*c8&�x\X�`�`h��ױ͐-{���|Q�&���e��u6;�g���yv׋`I2}�y���>�4?=yǇ�o&�H�v{q�NqE�����셅�zUb��~�U<}�e��3�5`�Q�u޳�QfY;d��� }��+�ƌ�'���|�ut1JCs~�C%���l�{IlN��gS�x&,��s9k�Z�f���1yh�����LjC|8=w�.�c���38��7�������Xנ�Ag��.�U��%��i�X���+^`��GK��׶��F;Ђ{�j
��f�sb������lԳ�� ����2�8V*�W��[�y�;?)'!9ة�jB����-�S�f�]��g
�hf�0dw�.�oC	�/+�\�p�ؖ>��hשBY�wȑ�H_C��ՊÌ�����*��\����ҕ�2�1��i ��`��:���w��3�a8�NL�,��I!�S�B<��M��3U��:���|���R/5N��:��*;\�L�J���D]nǲn�u����%$�>Y�|�K���e�]Oû`����ѷ��� ٥�?1�r.V-��f�a��5��X�&,[�O�'�0���OU=�I�=>d��0�?;ܽ��n�xȦ�LQx�WTxLzn1q喹H���� �S�$���$�F�w
7]��C�/@�g��Vپ]�& �,�7M�2ۗ/�]�4M���p�-��Q���t�X��jӾ����G:*C��H�soq�n+��},$O��3+6k$��@R��6�u�x��2�Z������TtK�ۡ�\��o�7�����5�&����I;��O��Kǹ�̏a���O]��ؗx�cou[Y�V��i�~���Z�ĉ�*��U�Y�V�C��/�n��$�$����ڢ�۴UBA�h]Έ��3(����h�C���E-�`�N�:�*�Y�[��h�$�K��](��wC�Tѓ���hjV6�Mj�{�T�$��(E�����5M=2�C��ᛏi8��st^gL4�Jy�$��@$r�wJ|�Rb-��d*���+	�M����7lThtV�w't�j���0Խ�t3WsVb�+���A��h���w�6�[�W�0���K��R���$�zG��-��w��t�KCh����nh�T�΅�D���P��!h����#�ӽ�:^
L�����ޣǎ1�&+��r��PUN�"��x����z��n��V<IK楧q9,��a/���:$��馗Cx�jf�׹'ěR�.Fn�ıBt��tiktV�qBG{�N%��r��<��Om��DnL��ۄ����6r��(�ڙ��L����/,�=�������J	r]S:��r��g���L>�T�j�"��2i�L�I'�t7U�7hq��ZB��)zo�ȃ\۱�ݧ��)�o���	�����m����n�P��wD�f�rw�|3����y�0˳��R�A`��^�G���Q�ڻ����N������tz��}p71@���p��/�e@tg�8N�N�:��Z�'��=k��-<G^�϶�T�yϱ"bW��9�1N�･V�C�چX�xcޝ�W�U�ܥƧnOH={������-�-�d5 ~>ceLl��n��e�{�Fr����SCj&f�'6�Ptd����	�VQ2��� }�w�q��$�;C17��ݭ���g���e��3l�{.c���nG�����_f����w������!�v��=6�2�X�':�z!鋟W�v0���N���R$>��/��YY��v���+�J��gy:�/!ޮy���oK[Fnt<J�|,\as;�`ᴰ�+���j�y!!�ź*�w$�\�����G9����sx��g�^����/H���MW>]���N&t�;�sÁ8�|_T����oN�ɳ�*��Wn����1�2Q��{^�Z��Єc�5h������w����[{��l�I پ��H���<���k���g^�ֺ��t���c��@�$n�Y
ƹ��,[3l��=�-�l�}�O���Ս�:��S�L��4U���7P�|"r�z�*VL��pۚ�u%݅�)a�W�;#^!ѱ��yռiuҩ�J�l�)�W/=�w�a�2��R�k}��}|�phsCC}��R�=́N+׹�0w3��&�&mAp|��|/	귬�'��>��]*�>_EW��\��)�n�v�Өf�m��/��x�͠�n��<~�/���@*�O^V%	�>3K�U3h�<C�m��/@��Y�NS����ˍ^��kH�c�F�����l7�e�x<c���#����~�}�v�ϳ
P�2b�Ǭ�UW��!���q\>T�=g[7�o�ˌ{��ʁֆ��Ӌ��̹���'��pv��RL�<�jеZ��On��U��1��sg����D���]���&"1�7f�ޞs'^���F%�op�[C~76�l���F�г�{2(�eQA\�q�Ɩ*��V�VZ�o�͔,�|�)�	���bs|yn��x3�ӑ�cRl>�q�%��!����7R�lK��bIԉ�&�kQ���
<WwN15�l�"���Q\c���R'(�����;}�uޭKr`6Sb��ݹ�km8u5%����xulO��n8�v�|_q�`���iXn�w|;Ru�|5����z5%ƅ��ttFv-Ƞ/��|��ᄰ��͔��o�l2n���8��\!�k�)Դ�������\q�z�q���PU-X^�u=�+����ӯ�uø.�3K��v6����x��]�%in��N�	kE�����r,E�+�Ɠ�bݜ��f��K�qHo>��M����#�<����]�gk��0�xֲ+$�����:N�T}(i�:�CyV�u�w��7=�7y冭��l���ؠs݇{צo��6��ď�竾�O�{��sc>
H79����t��շs�U�g�V@mwf�w�排.ٜ�㲣8-����wB_��zᆎǩoM�;�er��d�`����s"�<���(�b8��/���y��v�$Vӽ`E�L��5�2��O��3Ԝ��ޝ���3�r�ށs5��s;f��5\��w�*_��;��I@`�;�Dl�
��Rh�\�F�ý�t�s�X��ڏNo
��]��*#.�{�`�>:�z"å�2j�9�
V]�M�tGx]���/�������)�� ����ٖ��7��|�����C��#{�{���j�B���q/m��<M{ s�<�z��Yh��2�<��g>���^~�[`��7]C��w��_�o{�iA�۞G|�&�]ؼ��~nW'�=�zK|��x����1����ǛY�z�1����#��덌�c�nk�$TyZ������>�Ŭ�9���8�L�{{��n��|��|���WD=��R��}]�Y�U��97�ܕB�12f�/ne���S�7�LZ�{��	^Lܠ��\DV����ʵ�_j�6_.'w�X�ҵ4*,��}��4`�&')������+C���ȓ'gu�-������=�m3=�E�xͣA!o�ՖD��	W"���dZD�Zh+ne���pxu�S��p���S&����w]m�q�Ȯ����f��f����8�s�qDm��u�e�"�Դ��k^�/:�c7�֎O^��/�Rb�Q@�����oY��u�{�y�[h�֖���Wǒv�_SX @ra���@�	��Q�W`3k�-Gfw\�;Sv�y2�D��bN[ŧn��rB5|Hq�^�w�K=����o۬���9��S��aѸN?v-���P3�x����^��b����{��&�GZ��sk,��}�5�*6w�>n%��}t�O.�=���h�EǸw�k�w�s=�G����d�P+N=�0k�*��t����l�8k��D�zzW[�.�r�����U�]�<24�Vf=��n�Zr��xv	�F���E�Gǋ㈯	�'��o����<������5���"6��h���m�b����b�`���Sf��:���Q�l�掴�5�sj�A���G�����k��!VW1z�n�`�ZV>w��<��V�چ�v��c��zM���M�Y�4�}��I�W�7Ft�{B�fB��\B��b�v�;�jM��WPnf�G���kF�:X�	#U�;�v�$�DLч9�7ks����Ô:�gs{h�+|��h���r�/md�_f���,>S��A���Y��s+�-�z2�7QdTw���]u�Y烮&��%����нzL�|ʞ��gU3Wy�G�����Oь�O�B��-�δŇqݞ:��87�o#�k�=F������N��ϴ�k|� ���=�a���,�g=/�z�ٓg�j���p4�](� S�4���s�������l�K}�]��PR���u���o9l�v����Tu�|�����,ߤ����iR6��6�+@��=����\��vy��:���{�|����A�������Y�!8:�XU�db�Ҹ�Ef��S0��x�[J~s2vu�i�]4j�K$���������vCB��[����3�]���9�\���T��h���|�oQ�ܝ��h}�Rh��6%�^��k���^�Z ����s��yn���ީ-���&����Nl	,�2��L�Sw����+]���*P��p.����Y�Qӛ��t�pE,�k�9A�3y��r�L�͝E�#n�,��~�KK�z�Z��5A��͛��mprMA]h�R�fr���I��[��,2�ʰɎup�ڄ�4,r�W>��xt���;W2Ҩ� :'\�B���/��������{s)J�l0.�1W�ZO
m�"#4�>
{#���If߻��1�f���ƈ�v���M�M�5�M쮕ۗ�Cv�&��&�n=�����%"dz;��<�r��P]n\�4ԢE�,���H|��k��n����}��w������=��z�ѱ�牤N���|�u��h+��c;������d�ٜ�p�SQMG5d�Ρ�)�9 ��SaC�bA�AU�W���fY����x+7r�����	�r��w�����A���&����q�R�w�Y��Zn1)��XGM]7���-�
%ւa�R2���b|��p%����nO�xWM�6��TjR���ٽ���Ch��h�����'Y����Y�]���o��Q�ބ��,��D����ͦ��� Nɬ섋xt'����k/H��a�PRx��.�3[w�1���`�ѫ�s/'��o�9cM]L�3
]ĕq���՛���h�yƣу�L����?4��k��g&���C4�-�GwmD�d�N�ƹ�}���2�bw�0�ղ��U���/>:%���tԁ���2�z�3*�e�{ފ��Ѝ��1�}�
&�D�p�݆1%P�7�'�4u�eX�fh%�W[�����&�Ƙ�f=J�{v�����xn8j*�+2��O"4���-)�Հ�"�ҷ���	���Yd�Jf�T���E"킻{�$�W��&o����k����o�Pu�X	������6��n!5d�We�5y�q=�=}�-Rs���� _N��*��*��;VR����s@�jVP�@�eY31<e�wi.�I��6���R�i�`���b��,(�9f�	�{`�=���0�D����WP{����m�Ix�HJ>����`�7s�8 �<!�lg`�Hs�Pչ�\�%;�nޢʹЛYQ�ь�l���4n��������}�{َ���]]�9��W��FtX�<Rz�vwf݋&OWr��y��
r5}��IR�C����m�X*�-_F��4�G�w�5r�������ᆆ��io;�vF-30W07�˺��6l����:�m.�p�Anj�EfJ�G���0_\V����E�xke�8��=\����d= :��l=-��1�O�&�l�p'���]FH��(˩�����r�X��}�C�Q-�5w�Ϣ�\H�kCE�͙����7���8z��h���IԷ�:���4/.a�:��z�g2[��ǶR�̣E8��6_h�f�L4��9�}�.i��S�7���x(�����%X�'�<��ZAF��ը^�9����%�Oi��ڃ�(8�9G!Z��"㭍�)pz��ѫ�j���V*7y�-V��u�u:ʿ�o/y�^���d��c���~C{Y��6C�z�sw���S۽S~�/25Q��Q�J6T�x{H�ɮ�bcf�=��>��|�e���mea��]�]��c���b�=+^�r�(�̧So���S<^�^H=��+�^�g]�Hy̖�{_/ex|YC�+�Vy���U�27l���d�n2������_a�խ��n[ۏe�y�ʝzyi�3ovs����:f��A#�Up�Gd�ds;�{;y!Lg���Ί���.#|D]Pq�
	Enn(ڥV���BYD��PԈ�']dܸ@��u���L(�����G}��/M�����W���H�GNݼ�t������l�F���S��]��X̵��e^����#WA]�<��H��;�����ʖ��ҥ����g M�R���y��Fg�g�oy��\��'H����ݒvYJ��{淼r�|���@�$�I>��JWaj���/E����W,��V\=�)fs��gru���X5V��n!�'v�v�g�q&z��K��vⅸ���m���';m]�����7��⋝����.�T'�Y�M�l[���Z5�����
=�X۶%���֤�dֹ�h���:��V�v�+���9���c=,#�8!ή�>����g�o=Y��۬�{
X��u����κrŒ��'\�q�8�woV<8�)��s;��9v����Η�#��<8���v�u�̀����ir�Vn<����M��8���`u����]��b���؊.xŝ��λsY��l�َ��<����ٽN�q׶��ܭm=���J�aշ�Erl	�����k��m�7��[��+�y�z�|�o<'&M�j��v��؉��SS�n��MՉ;�g{+n��W�t�^���^��k��
u�v� ����Z�`7i�ƼF;��6C�w��/�vժ/ ��tt���\��f��wq��\e�^^5X��lz�h%��&�3ٵpk(���	k��,���8��g>�<���u�s�맷D��[��1Y5GE˷�;��N�1��u���3�m�]J�)��Ye�v(H�Xɸή�ی��V�[�/<�nٵ��v۞�Nu��m�b�v�>s��=�ͱ��]��-Vy�n˩�9q�lr1���-��0q�n܆m{�M��m]�j7��>q�G�B����O!��=���lu�˂ŋ�����]ۤ67F��r�n�]8kBnN��k�8�.�b��6׮�/cn� �n@Ta�v{t�Ӻ�l��c�n�s�k=�ʹ��W��s�OU��b;�y��V���i�(/5��ö�چ���1�I�y��uĽ��ss��a��0��l��G9�r�����WC�չ�}�6�of����{/c-��[��K7,����vky��0m���ɨN��4m,s�iv����|�힑3�z�K۬*s<�7v���bv�q�y*=CaNz��d���׶��y7�ݻs��4�p�q<=^VM���oY�W5��Dq�Ξ���x��]��O��9�/��[��4q�.��x���z�8v�bl^U�_"�{[��]=�pv���Ŷ.6�q�'ml\\�@���F�kn��v�	�b��s6�x�yNW�=�#=u�ݵ��<�����I�l����Gm��B�gS1.���Ƴ�K�\�e8F��\���j�)�R���v�飒C�Έq"�y�񷃤�/�Q/;�\g�>7��9�����4��t��O@j��-��w>7/*{�6�HC��yz���V��q���:g����ȝ�`�V�9��N�]�n�}�fMx]m��S���R�rC��A�9�η�W7hS\���e� W'O$c^Z�8�5���a�����R]�����8�<���&�\*���ڡ�ۮ;v5��]��f�@V�+����k�7S�t��ǛT�\j�vi��u=�ᩗ˹뷺���5�q���S�;�Џg^gɹ�� Y�l=o��ʽ=�c�N����`�G����1�sڊ�2���+g����q���p���ڣc�}���n5#�tmf��Np!��ļ{v�S��9�s�T�n���S�ܜ϶�Wfy�Ŷ���=�<l/G�:� ��|�u�8Q��mu�ص�Aǎ�ؔ9���`��o#��']Sq&��=�]������`C����+��z�Iֳ��#k������z��7>���ŸE�=��c��"ݙ�l����r=-e]��_cg���t�Uyf�88K���\���]��+p�6�)�AŲM�&:H�ۍs#�O6Y"�_���H�b������װM��W\��絸�n9��U��������n#�3�P8����s�9����Kݶi�Ko;����ꈞ*3��só�M��ݼ�8|��r���G]�s�n�w<mw%�8{wQd瘛,c��t�����%�M����6��6;u��u�.J��Kse9�wn8z�d��A��
���Z�s�G&ݹ5�CF�G�����6���v���;���G=�۟;�q�X�2�=*GYs�s�9��<۲sn:ك.�<��-A�8��	�F��ѝ��<�I��R�=�s�=p.�	�٠ݍ�7��KkB8X��k�땎�;v^���Zɺ���@H�ٓ��v�#ұ+�װ��Y;>��u�w<���ܻc��X$�N�����1a�%������㱹�vU��`N�ӊ�q���9������}[ض읜�q�9����hݸ�-�n�m
�������������=z�V����:��#V@�6�۞ݫ�6��/oU��-��<m/�.��I�8����F�P��c�<=����u�q��u�v8�z��r�6�]��u���MvQ��1t�"�{[�&%G���g�^"������օɭ���f�F�ւ98Sg�9S�i�v۶�ô֍�^�d���y��w���f���z6�Ş�[�O��y�m��m�S�]�uu���O'jckr=�f8nVa���n�P���Fu��u�%d�uv��������X�{(s۞r�x�&N�K���;�䲕���0=��a�׺��t�v2�t��Rd�d;��.{kv�݄ƙ�E��8x�6��<�;]`������� �^�-�Sg��t'.�ܛ��v;X�dl�Ӯ�]�c�n�������ws��hj�=��Y�X�ǝ���6JV�K۩�������/��'�l�U�t�h'��3ؗk�/p��`^36ָ9٣=ڷ�gN`:��&ۥ��vY�v�}�5�{
v燷m�N�F�s;��/@���I�g�:7/5�[R�����)�+�wm�6�7t��6�
��r yyܻ�|v�Pݍ�6볶��Ӽ�0�3�1:�mεڃ�l��X�JY.��;�v�g��D�����n�̞^H��Ւ5˱.����]n^۷mv�sN��y㢻KJ��G-��51ֶ���k�/n��\'MtO$�m\v���O�����mujT=,��RCU��g�瞊V�lB��T��l�\ѵ/[:Ʒ�l�W;�ӳ�;���/%IÍ؎���M���bBM�]��8�cM�$gnˣ\�=���w��ꎮq��v8�;#��k�V7N�kZp>dn���.��d\2��FԾ�v8���;9zm�m͌�8�[��^v݉��+u���rX}�������v{\��+������ͺ�Ό�m�9�۶�X7f�v�,i��9b�n%ؓ<˷�Mvt�ݔ�nu����z���s��)�<u�Gm���Od:�ކvx���9����n� ��y�
���Φ{y7���jx��v��������$�<�& ����}ۚ�W���� ӭ���V��u�	a��-��Z�h��Ny�`���b�nzψ�N�ٟ%�7
lj{C�zN���:�r�8컦'=09V.�7;s�JL��I]c�,������rN�Bk�n�:ܢF�eۋi�nB;+�}4wX�(Џ�I���B^�d�=���<��3�/6�Ԥ�w�bȧ�UC�wYF��vH�%�-n}o9p���nM��D�[\p{<�8vĸ�;G����͞yW�n`|q\��v:�nt�׃۪�a�=\x9��<�F�ddM3=�n�۔��ƌ���ܣ��A{s��r�Z��g�W����7i���cq:Q�Y�v���V�<�gbz��lv�ӻ9G��ft)h,C�[=p���\�8��o]Q=s�:���ݰ&��nw�퓲�Q� �<u�۳=ۍ���[��7v��;�ӭ<s����g1��"<�ٜs�<6W��]�x�D�����ZK���C���k�G]��2x��$�pu�T<Cֻ@Yء�+��u�m�Դ��jw��1����e�mp����p��B��XΌr���l�s�pk�`<���c�;�.e��Ѯ{8����\a:�nzj�NR<wn7������n"���8n�χ�5��^�v���d�qsk[�;u�Е;�u��q���M�7����G�5�����$=��x�yƈH9M�^N��j��0x;��]�k'�Q���u�j�Ӝ-: ۓ����{p��C:��n��-<�d�\B�S�n�����Tcu,ON�	^
�r��tn��ks��z'�k�����-���]�c��L��G�b�^8��luqp�{�n5����y�"Z#����Y�m�n[v�d�ó�Y+c�6��{5������y��xD�ٱ�9��R�s��۞#n��赂�ڹ�7��;ۮ4�eќ��kV�qE��m��}�1mv�]vj}!ۂN��W[�s��5ۍ��J�Dch�r�lc��<Ys�Ƴ5#n��rÔ�p�3�ɫ��y���X.����N��tn���Vˇ���݁�qɷ1�z�9z2�OEۍ\��[6V�2,��9�#�n����-���k�����;A�j��\q���nG���c�����͞��&7/u<<��M�4��c�y��X�[{.�ۦ<��m��U;U˵���^OPm,�۩jS�۔r��
m�8�ٜi#��7]pWn��GoZ5hv��	�t�Q]l�q�'in�y.�s{]�����i뭫��9��s{n���hŃm���̇<z���8�I�6�g��6:ݤ]s\�wA�x�m�O��+qs�cm{tc����j�l�ho�E��n��;���jܩ�ͺL�&�t�Ѽ�[�.:䍮�0��L���m���)z��	v���ˎ2=y�:ص&��m�;�cu�rP\��F{j��MAv��\���5�*���5b�H���=t��a{v-|y���uݠ��kNn�;��J��!�q�={Q���e�Ǔ���^Ksm��5OZ��m���z��~�v�XUgma0�V
�I0���6��PPX#TH��ʦґaR����L5,����6�e6�L�(�b��00�ֵ�*)��J�2�$�\�����Ra�AEU0����r�E��D[hd�%H.-m0����B�R�A`(,X�0Ԭ�DB&-`�@�V W	X"�A@Z����-V��!������a�a�q��(e	iX()DȘ`)�ш8���1�
,�BaUSl��J�1���Y+�eH�)T��4�I��Ņe�U��p�!�B�[Fնʕ�T"�(ʕi*��kG	0���qR�I�\�-�Q�i���}}mo�����}��u۠ѻM�s����]af��c#�x7g&��X��4����v�<���M�rwT\�7/Sg�܊16zɓ/ny��y�{h6��\��U�/Z|�]:������mt���46��ִ�\v��8�{Q/�p�����q���۫��p<[������9��4%n��T��a�/�n;s�3�Fv��B띠�v�q�9w;�n&9�a��dh6��@t���n.Ϸ����z�{s���۬zm\n��Y���gn�.�F��Lgt*w[3�,Vn�8�����vz$[�q�w2��*c\��O[`��Ux�۰��c
8v�E㷮:;m۔/:�/�om��Pٮ7qs�\ͽ�鼜���=�@�qa�<�	%i��}��f�]���h��wV]�k�t�A�������V:�Z������i,���.۳η����A��p�A��:�kH��e3�y��,5me8����AY�p�;���T8��i��q�l�.٪�xܞ�5�����iNd��#����nѶ�d���]{s�Oc�n���v+F6 [�[�nA�\�Y�b�]se��ڝl��zݢ�磶m�}��ȴ��q�t����ԡ����m�c���t����{K��ݥYqۭ�^:w*��<��nuӞ\�C�;	�C��7�����`�A:�YA�2c#�'G�;Pl�����`�ʝvNY��#��vpv�����%]� �!ln�PnĽ��;7K޼v�cvN-���J�9cz��!���k�۰Aٯ:�������ݾ��.nL�X�L��f��=��`���W�}���{�㌝OgZ���1v4�\����Ύr��]�n���K��ۓ�*b�F�7<�1������d����n�K��㕫=w��M��=]��k���\��7C��I�{-��Iz��{��[�p��G��ʋ��������r)���x˹˝���ݶq��v�ceù�x{a�m��-WW
1p��R����-���08�[1�Lm�d�;l)����{;8q�d��A����nۃ���W�4���q�\"ھ�l��v����ώ��l=����9A��x�!�c�*7Kkh�m\ZV��7J��v��H��
'���ڢCo���Őo���2��ߗ�}��\�'�:�cc(R�`�&b��菁a�5���������R��w!)΅R!������~w�s�MPU�W۫ܩ
��4 ���y'/Kz����nm�I7�@�+�������^9N)�E��\�]3��(�O����\���(0�]�V�BJ3�"<�S2�E��0�}W26�G&|J�m�I 콟P$�c6t���#�<�ֽ��3I�[��8ɝ3ǣ��Gg��ؼgƷ;I�(��Ro3`鈄���H1�ݘ߈ ��+���l��ks�3�+}�L���F��@�"d`(��g���s�>�c�s�z�f�aծ����b���Lf�;���H��ޮ�:.�Ӯ�t$2����.sN��3g(��vH���~$	/hW�$^�k`5r�j^t�:�	��G!$�O)�?�뀂���i��b�=���N�߰会	�������D�TĤb	T����tT�b�UNh�H�Okd�����ןT�5�����\�� O�=� x��b�5�0|{wn�:sy���UB�'��9 (OsHf:��N�e��n�a��;�su�sیv�3[.��n4��<�Ltv�_+% f&'o�!%�P3�ro��H����I��ȗ1Y0�苊��ɢ	w;��1:�3`�1(ʐb�m�7�A��p�G��+f�_���ͧ�|O�;m�IQ��*N`G�O�h�(̂bٝ�m�M�m���1E�R��:�1���~�ħ��6t��8����=w���9�\r�*���M��ш�r.7gE0�qq�*�`��@u��y+V��:*a�:H'ݓ��$���o���h�$�3!P&dOeH�=�{2��f���v�$y�2�����R&_�	V{F�}�o
S2��%7<����x{���q�z�1��׭�O� �{"�tU~�[������6\������7N�kc�nI�st`�r�cx��%�n꟟ߧ��b�OA��b^0�;����{"��J�m<����߉�#;^�	���&D�@l{4	.m�R"y��or�A�M�	�筐O7�^>���O��sjx��/�>Ǥ$Q�h��O��A$���"�Fb���,�FgV�I��퓶�"��!@��X��㔝�f��GA �=�`�H��B� ��ڬ��̔9�x!+$>y�$�p#c��������G{ޱ
���iu]<7�-��,S�N���ft��ǐ*�������k��U�U1�iG\�k�-s$��O���Ʉ�� ���q&��ۭ�����Lu�0��8uV��u�x��|�['r�T�8;��$!J	"�	Bj�9� W\d7��$wnz���snve۝GnA�������d��1 ���5����2��$��ks�2+bj��q{uu�$����O�^�rT�&�bdP93��'����w�*^Uh$	^�z�	sݭ�B���8�u��`��A	d�"|�6gd�>'�緛$��*��n�,�����	�Ǘ4A�v�*�9����"T9����xn�fP�7��U�hI.{6�$�n����y�����4H�8��Q�>P!��_W6H��t��麪�ˈ.��ɩ{"�'7X`�wn��DWk��͚���'�*�\M��9��o/�0M���=��̐DU��YY9p�
���١5<c��%�\r{�S{��K�{�#7ɖO��b8����`cf���\�m��g=�f��(\�F	6�;qͺ�	*��8i��㎻s�i�R��e ����h��lj�`�7�g�6��雍�ɰ/gÇ�['����vM=lrm�i�dQ�v�.ʛ�����e�d�l�����U�������m��a��GX1�V�6\�����ͫ��픇<�g�L�oh�0s��u��ny�b���{n9AT������rˋ��N�����֞��v�@��x�%����v&Lȁ
����}@���2I�v�bN�*ד��1��|�{�1��d���ă0Jo���Az.��D�v�| �{�|({��!Y�5Ze���u�L�ൔ��8T�o}��@?�u�$�a�J:6#��zo9�I��m�s��$��B$O�
`��N�;�&��Wn��$��u�	WuϠ<���0]�?��h��S� �d�@�O{����]�5�]ľs}��%vn��A;ݭ��]� �{s��Q�7`"�̂!JJ��N��g�$y�u;�������;t��=0�����JI�DF&���es����5�t(Ȥs��J�6��$���n�'.�Y���X�n|g�X��l����g0x��������柋4�2F�1:��z��0z:�GE��ّV�db0����щ#o���C�Z׋:s�j���I��m��[�4A47��ZE���Sux3{�d��)�`����O��nEr�څ�E)��|H��v�$������3�&p4������r� H.7.� �L�]
 ޼�B���ߣ�˝�])��7��ÂeǈȏD3n�	'���?<!Y��T��V����� H�y��#�2��Ͽ���v��ܺ^��^9�j/c�NN{��pcd�4�Ъ݃a!>�|�֬��p��v������@�"��6vɷx�l+ptR��~5{4	��IA3�Ķk��d�a�DzVe\w:H&k6��o�9�<Yp�s2�����Oa�x�Gi�~p�H6���񙺅��n��E��O�讕'd�&�Ǳ��5�[ z����Ggr���~{28���ذ7������G۸���i�+s]'^ڪ�t"U����ս��ׯ9�Μ�$J���S���uuR�B��qgė7S^$���9���5<;'�1C\�� 3�f�i���^�(DϹEu�	=��L���s�VNS�YB�$��a�Gwn6f��8�JD|�ߺ�W��U�+c�ֵ=t;�{Pv��h-��m۱����uԟ�����sۏ����������}L�	�wn6b%WL�b��������{��'��cZL"6*�%@|�o����vAs7��l�;�q�vA�[s��LMl��\��D>�0�Kݵ��@7�{A��D�e��"�;�	9�6�'��s���{}�,1�I�L5ߙ~rvN�˺��f*�0�>w^�'Ě��8^�W���m4ٷ�X�~��Fok�0�����c��љݭ��v�\���+��Z�(�ǉw/f[U>�3�H(�����w��o_6�V�2%JJe�b��y��	�{4Oi��ՙ}�$����'�^�	'Ƶ��1}�6 ,�?���gZ80�q�q��α\q�ul����=����ny8�lf�i������ۇX�dp72��	=����կ�P8��;��M��X�>=������$,FfaG�g/��,\wX4�t����V�	�U�4A��
�VӜwzX�u!�K(����z~�J	"N����	%���*9)�ڸ��]�C	���� ���cv��P�T�T�z��U�c�Ś0���x�*�k�	{�էp��u�B���7/b���1
D�ѫ���H9=����_;Oa��;Z	 ��ɠA$=����W9�S�ɽ��{�mF�ǋs�r7[����f7n���-���6���2;�XW,'�tr�����ïEk|��q��N_�3����f6����8���z9�x6� ^�7YK����r�j{po66팻j���xzĤq�s�a��:9�����f��l趃�ywh�i1Q���k�ӪGr4rA�3�5��nf�ݺ�l�W�W�s��>��=��ǐ�^���|y�j]q'&S
�}[�x��N��n��X��^璶��-=����3;@�i�\�7�����=�ݵ����%�v�e�;B�����dJ���3��	׸�$�n�A!�=l�7����3 ���'ă'��;̜KA#glCW���Zv�������xh���t� �gH�A{�m�	�Rh�
����%0HX���A��z�`$�o[d�(㽫�a:���� �5y4%�m��"��Q*�2&;���]�Fނ#f��	 ���l�H��ȫʜ؋1&�k~1��D��A��	R�*[�5ϵ��|o��?-��sT�3k�M�v��|	���ߌ���;w�׉��!$XŇŤ��"p��r��'����]R�7[��������D�"bE�\���n6A$���[8�<R���ՙ5�'3{�޽d��$��a���ܠ��8���r�N��v:��KA�!f\�<�sz�QG�S�l�\=8Z�d���:������_mȘ\`�;�H�Kxb��' '����������z�'ƸD��Q��R���@�/���!@��L��X`��{LHzq:N�v�;�A�Ͷ�$�s�~;ҕ�FD�I���
`�ۙ�ư��X��s���w=l�L����q�1\:�O[��Q*�3&1�����I%�����?r��П;������$M_M#.���s�HG�s풍��-8Gocv��61�q���t�S���C�b�R�;�X.�B�@L�N���osp����H ;�@�a��Et*�#�]�	����ɬ���DL�P�&&�M��R���{QyLA>�׭�H3o��ĠY�#g�)� ~����}w�,�I��
k��wH?��V�{��E�.�΍��f�j��☓�j�̱��f�s('%#P�x���noz�K)T"�֏*Â����ŝX��Yd�[]//�]�
n��P�ܭq�ܗ�����ݧ���D�\��̦Q�x�#{���B]�~�U�&!zl�B�'���_n��p<Q����m��ۭ|cWlݐ�s��d����=� fo7���%s�GK���Ig2��*��3�>w=;�P}F�>�oFL�F�(�=�z.�:�g�mO��CU��`�\P�2�¼����!�V�1��Q�2�3[����l��1@����(�F�q�=ם���+��%���B��ܙ�%�̪�V�U�,މ��iG5�lI���ǳ&u���2��^)��`�yӺ�N�}7�L��w�\�&�L?EF<v(x.c��ž�}VMݘ�S�Fj�Ű閸�z�r���U�(9�p�0Y>:C��BkS����kXUC�zAelU�f�ǂ8j|\���1��:��ӥ�C�� ��ћ"�^>�����{�DgJOA���W����2����\��Ԭ��Jy2)Po�+,l,��",&� �m�u���V
�����:��~�����}ɰf��v������LH�&��.�2�'�3��KĻ�˜ٗ�=��xa=����e\���zü�"���������O�dY�{6�j:+��W�Sk.
�QYs�*wu��m��@Ӆ�=d�̾׹���:�'��|�L�d]���&�����!�j�T�C�%�
��4��	�d�-�B��3Fʒ�m�V���Y0�.Xr�T+!m"���(c�	�-h(0�`�RG�
�jY��B��b��j��d��X
\\*�IYŘe�+Ra�J�R�Æ1B�%r��Q�j%��k
$S8�6���n08EÁ�q�╬S8��c {�{�6ރ�ۚ��\2H�U�
�T��)YX�Zʊ,P���a0�" "f�Ve8dX��(`�U a+*��	�L5AAUE�Z��(1���P����[Z+l+��,-���z��G�5�`�L��W�
��HP$�3"�G]�t�Qp��c����.�P�A{۬��:�P�7�}�`{�͒;�+�xoe�.���~�{��Bs���"6{�I�Ͷ�� ��D_v��1\r�{"��q���"T��L�*"&9g�c��͹ۨw;t�:�nM�j�;<ni���~~��9��eB�c����I')�� �^��3M�
=���Uo��I��{4	����&j���nhWo���mg
�y�C�I�}>�O���l�R��z���ox�����0��%�p��pI�n6I�[�l�s��9�[�}>�C��ly׾�R�aL�D75ݎ�5U�x��I�ݚ�Aw���;z����&R���<'��+\��kE��.���j�JJ6^w�j7���9��ej�=/�X:�6Պ&A�k����r]q��:��	*o�	��qr$��"ؑ^;��d��ܦf}�Sǔl�~y� �tK�S����@���7M�m�9g8Л�c�흼Y���ǋ�z���nzG�"J񘘛z�yr���3��;.h�yݏ�O�{q�u�h�n�$ju>`�ۦ&L�)�"a�P����{����8����m�WO����~'�ݸ� ����N�wx�ȥ�&��3�&b���l�s;r��AC��%"���6hh�w�n���ۍ��Y䈉�" �Ⱥ���>}p��WA��۴��U��v7e�|	����}�%��i7�15�͒EV��'M��`�pz�N�[|� ���lA���9դ�������q��\rgǴot�]Gy�y��n���hm�ǽ�`���s�[Y�����Rԗ�d��J����~���:�*��\���뎫d�nص��=����3s��6�GV�{u:�1ɛ�WvOm���+n]��
�5(L���p���ƓF"�&N�#$g�=�:7Z�݆v��d�;���q�-�U��ޯ&۱۩�4a��ۈ�nz�7k���=G�ZN���P�g�;�ʜu��M�Q"`�w��q��gGkn��x��ic��܁�<�Wkln��Ÿ �Ghk۲\V-�9�7�+==�?���
����H��f��wwv�'�U��Fc,�� ��H���lNv�H΢��"&&̕�ݹ�2PI�K������Aw�$�V�}@�k��q j�~v���D�,�Sx���w��$�kM|��)P����1�O3Ă@����I&���#cPV��S�L��w_Dz�dЋ���:�zIO���I�}B�H$_gcZsb�n�D�s�������6�E�翜$���n���I���x��6A��׈>$_gcf9��l8zV�6 
}2R0!k����x�!�E]����2���v4��ݑ������2��Q3�؛y]�I5�f� �H����]5	���dl�s~��k_M�-��� 6M�4B�ބ��x�:r��IOάop�O �1��r�"��G���nz_<��B�����4��8;�4����rnr��T���HW�+��E�>a�n�FN�������\�5����)�r(�}ϛ�'%a�(w9��A�Κ ������xYڦ���R`�P���ؓ���tq7ǽ�s��z��~���_�
AC䕅;���Ì80�,aP;�~�F�{�n��-���N)�~2j2�Q���Z�iP)�k�\[�8q�ݜ@�V��y���B��@$ ����#����'���m��?Fi�k�� �m9�y�C��d�Q�߽��8$�.�7~���������.���5b텱�ƣx�a�O>ɇ�{���3��lg$�/������5'c��x�������m�ID*J!X{��G�KR
;�~�g8	X}�~����q���c]oﵨ��iK�m�xY��^�>������D?��$����8�Y�������7'=������bJ�XS�{��a�°�
������I�+%ed�>N���sM�W�U�	 s�(r`1`K�m+�|�P��H(��}�|�-��(�r�Y��]��[���0l+��H���'g�Ow���?:껓�E"��y{}�͗��F�s��Ԟ~r��g��R
x VQ>���r� �P����C�J��3��1}1�33a�Y����eP�Q����8����X�H,;���g+*�Xy߼�g8� �[���
c�c����2��Ú�}�8�W:.|3��.s�\.�e<��}��� VPd����߽֍�%C[;���p�C�%aM��sp�A�aF�}��6�Y82�VW^s�ԛ�P7ǜ>/�ߚ�x����{��z��'e*��rɅ�1���p�Y�z�nkݢM%�����>#>��^�@蕇<�;���cR�=��}�|����l`V��op؁Q�>yѺ����f��ϼ�P�8�Yc%B�w���C�+>׼��%+��˜n��W{��m�ID*N�F|�9﹧�{�z��߹���A@�P({��}���X5�F��kP6Z@����'^�-�S79���^:���"�~�)�`H��,�&����'޲VQ����5�l�
$�T���{ǝ����8à°�*K�ϴq'��ed�����a�;��P�3P�	 2�����8o��!��3��H(�>�F�H[)
���ןy��S`�R}߽�6���l��wr-�z�9���^�˛B�K㙝t��t�'3`t�36����+*lM�%19�kP��^���!~ߧ�������
����h�V�t�0��q��9�1�q�W߽�Z��%�<���G�Ny����Ǯ|� �{;���g8��Z��u�=֠n���������x����\���>>[y�N�hz{X��v�0��n� n�m�ǋpѸ�m*��b��z>��BS3 ��$���ݝ�- �p+�y��H(lVϾ�~|,�#�{&�]W|�#�8�i9���N!Y++%]o��Rm*���y~1�ܔk��8�Ĭ9����(���-77���]U��������-)
�u���@SbJ�YD�����q���J���o�����:�����}吗��>F�\�~TPQ*�°�
��}��%�T�B���}��%eH(�5����Ԃ��Xk���j� �B�;߼�8�����S""& ��� M}}A�y�{�1�>�2�VVJ����d�Q%B��9߻桶�
°�(����G��a1ݳ��g���	>��}�|��ʯy��_�-L�aL̄"� m+w��Aǌ
ԅ-���4o��2�z]gΘ����o{���*P@��<�y�q�d�
�{�|��#��m�홚�b�˓
����n��hdN����٢�\4|8V�a��X�o^�F�E�]���e�Oq�.nb���:�ٟ������D��������b��:���\��=sv�kv\�l�v���r=N��p�қu��s_���}[���q9�K�X{�n��qqne��r���"�Gm�:^cI��5�%]ru�Jk���VwGn�c�oIW.��"y�����q�<,�}wn.S<tr&�r�\{�<�z96мcY��;ۓr;:r�s����Y�Cn�GY۞�YM��m��Kr�#�2i�I�/�ƭ��n��3�m�ͅ�'u�t��O����9�<�C���0�¼��5��0�*%+���4pg+*J�C��l�+Q�p���|�a�
7�]W�i��Ix}��W���M��;2���̕
�SbN�Ͻ���++%fkϳ��~�ߗ�o^�������P�J�Vy�{��ĂÌ*{�|Ѵ����|��YZ+��:�o����U{��Tzu�_Lb�Ɇ�ˣh�X}������Ƥ}�h�A�+c G/��_�A\0�.E;�� H�(��߼�8���d�Q�����pIX_��1����r�n�Xn0���u�����f��!��T�����tpg+*J�{�}�g9�k���j���Ӛ���5�|�zAH6�/3��̓�^�{4�BP&	�N$����8�Y�J�2W���h��P��w{�|��z�Xfo=q�aF%�w�4q'"�����Ԍ 8]��?TșBbA�D�!y����s� ���+�뮻n��.yżv3qu����|��0���8)��Aa�}�h:�Z������7�B�HV�
��wZ���*o����;�8S[��jg+,d�����hpIXS��}ǣ�`��s���q�~��5��
��Ry�7�v���啕f�/�˙���Ԙ35�;���R Gu�t\����UɿH���1�z���i���������D�����o�s����~Xk:���Ă�R�P��}�g
A`pk���Z��i��OٜfK����k���PStzeN(��Z��P;�}�OP++%H/��u�`�P�%B��9��������|�S��}�����(������8!Y+*A|�;�I�������1�Ɇ�˳��Xw��������:��5!m�{�h�)i
�i�����@�be��{�ڇ�y�|d���k�H���
�w�~�ĂÝ�y��T�s��83w
�l+����aRX�Ib����r3���;��_n5{��4�P>ϻ��H,H/w�u���h����n��|�-G���Wq�h����N��\`�;Iբ����c$��y�m�3ͼ��hQ$A�_}��B�*	���>z���h�q�Pd����ѶJ�IP�J���nH,=��Zk�9Ϻ���w�i2'��}�Ă��� �o��Rm*���<��0���8)��Ұke`���<+]ѝ7� }���!RA�[;�w{���
��O;�~�8�Y�J�|5�q�Ng��x�U� o��>f��D�RL%2&��8Ì+߽�Z��%�<�{��3��e@�Tw�㾟��?y\emZ?���"_�a��K8J�^R��a箻+�L�����@k��V�s�f��B�N"�.`w�W�U��SX�qk��5�}��x��+ư(׻��j� �B������P��l�ޟ��&	�fd�	�	!��}�vP�%�F�]w��q������d���5�c%B�������Ì8°��Ibw���#ܲ�_�z�w�x<	�ߪ�ǧ���1�ɇ2���9��<`V�,�}����A�|���\_i�[��\�
�@�ba�;ߵ�pd�Q����8	+��~y��>w�}�������j�amɱ����8�v1GW�k�E�kpq��M�-���_�n�\4��+����9���%�>����m���*���{���0n]�Z��ӕY�v�g�PHx�G��}��͟ �����DL����Dn3���OD
��X��F������y����|�M�T��V�}�w$aP;�~�F�r!Y(2�k�tڞ��o���g�� '�B	K�&b
cb���;��惃��������6�yHT��ιߜ���Z���,+('�w�u3�����
!߻��8�V{ݾ�L�ܖ�sH~|,�#ٓ KC�r��������Ib���jd�*��~��8��+��Z���07�Sx|��'�3l���?��P�C^�u���O�w��m����/N,���1bX(���ߟ���]�k�-���1&WD��_����9�C���Ύ�7-.s������O���4q8�YY+(2W���`(b�mq~����6�V�|��Ì9VT�'~��h�ND+%VJ����0��n��q�7���~~m���ﮟ�^����;R�v�Î� �#�������t�~���?�'�i������y�ߴ0+R�{��Ѿ���l`V���MN]q�_��9�מg��9�~�6�J�2T(�{߹��q%ag���n楣s�R���a�»��i�Ib'�ߎ9�^cÌ>��P�'�*�}�~捠q*A`X�>w9��i �Ne���}��M}^�#ٽ�(�����"F5iĚ�{��ȁYH�YY+���`(i%B�+Ͼ9�{޾y���$F%O���h�ND*Ad�+�;�ɡ*7��1Ne��)��A|>�w@`�����w-w����w����-�*An}�H)�>Dv�{^}{[�K>�6�罧��Ȁ/뽠�G���ë$ɑ�e�a��y���&�*JVw�}���&u���{����`����8��+��F�����m!m�����,��� ޥ{�v���q�+)��7�V#��[k���Y�a����@z�{�dg}ݑ�\\���~"��]��uU.�(�|/'�<��i'���\����GU�A��e���=١�=p�4O�I��l�P�ř�n-�:��P��G=�����;�[�����y����wUF턆zh��9y�4���gX��|u�{]-��G;w�,Ȥ�"q\̖s��\|x}��j�2�p5��|��d"�-�e�����3h#_�4||�١g�L����5ƴ��ݱjh��e0PC�@s0z�hP��Y���7�m�_#��� $o�\Q����Ӫ<�z�;��㋈8��w�0�� �a�a.n9�u��=d�pi��t��vhy�����7=OU�9g]EҜ/aW�m����s�{�����:3�#=�'ׯWo"`��;g�'l�^m]����&:k��U��O��l7TJ�Ŝ��	љ�8�	�H·��s^���ߠq�k}{B׶6]�-]�n���}q��&��3�A�4�^|W�k�b�˗^O��ޜ��x���;���x%BN��E&tl���Ϯj�T=�9��ԭ!�TLMº����[r*k[di[�M;���h�i>g@őOm���$�Mb�]�(&���v���.���{�3W����LuܨNѷ�0{�Y�����H�7\1���z�S�Cyn�T[4Y�d��Ý��G�SW^��X����c��nl~�?%1�-/�FҪ�)*�_Z�E��2��(.P*`b����#-0�V#R�ml�����1�Q�jĪ���0���J�6e1�J*��Z�QEU��[DDTU���"�
����0�L�A��(�Ub���Պ*��д�� �a+�p�e�YZ���2�e�8�V1���Z�h� �U���V%J��b5��rˊ\cA�mQ�X�ˇ��F$kUd��F�-�*�R��EAF2�B��T*�"*����k�& ��Q�*,�[kZ�)m��Œ�E"�*1")R��Y���%Ř���[aJ�`��X�6�Z�j�bT��TDF��8k�p�\1�"�X�����DETB����Q�1�������1FDX�LQ�������J��Z�qklicX��V"(�b�Z�,+PQD[eUS��:�nL��oQ�g��Ϣ�z3����N��g����q�h{Yy���)r��p�W�ۅ�����ˈ��U�n,lp�Ÿލp�2�'�lܹ��e�ӎ@s��sv��N��`�n�9б���rm�9z9��6�"�d�1����r��`��8��U�����[��z��bP�p��
�z�z!��x�zfgj��i6{br��g��`�����;�.;b�Z�	�q/��뛦=[��q�:�ma<�99��v�9a��]����v���c'd�k��k�isq�*3R�`��㣝�B�[���؎����"��'��l�nw�m˰��g.�>Ny���nwI��s�Lf�"�pP�B1Z���g������n��b��;��z��T��n�,���<�gqglS���a���m�u�S�����ɴ�����i�y���i'����>�����@�m囔�;]��V�^3t�M۳��g�k����w	x�j,�ԧ$���xҦac�¶:p�=V�ɸ�oG�7K�B��mֽ��m���Ƹ��ְp��۝���a�Fݸ��]69��=�=.y�cg˲�;+�q�;p�yhݱ�h`�^������y�h�6ڸT-9����m�N�#A��ώ���b�{�ۧ�۲� ����F�Y[�:�m�u���n��ջ�͛]���Cn�|su9�<&�rt;g��m����s8�C��û	�V'�Ç�x�4WK���t�}�xX��5�G�ٖ��Ū�u��1�V�y�	�é�h�]�3���FT��X� �uҋ+�Ȼd�m����3�`g�`����W-�ɍ۲`ض.ͺ�u��Oc��&��u����f��=��5ղ;krݍA ���h�n9��ۗz��dL�3E;�G�.��l>�۝XS;`��یq��zzz�a� e���v|��)������*t�v.�SL�x��Oc��x!�C��p�������w׀��t���l��ܙ�c�������0m����ڎ�&zB���d볔x�p����6��C�n��X8M��<�����'3��*ý����]v�mp�8wA�hղ\��̜s�;C<GP��]pz):7N�v�& �X�Gk�[��1F�=��xЮ�
�Ek���U]6�#��i���t��ݸ^;g[����s�x�����\����=`���z���\+�k�j6���r��zw��p��J�����$��;�'+(�YY+�{��d�Q%B��;߹V�s�������uz���J���;��8VJ��es��0c����Snfe��D�3�ޠ,>��=2Ĝ��O �}t�!iHV�+s���4 T����~纇�J�*�g<��;ݞ�j��q��|u\4g� �e%?�q�y��!�%B���|��4r3�Ĩ}�o<�=�{��w��}>@�J�X���0����,}ە�fπG����30�&&I��k���L�z�{�{���@�4�R�|�M2T��"J��}�|�8À°���?��G���#kj�Ǡ2<,�e~��4%@��dp�(c��MH,3���
ԅ-���h�
<��L��T���4|++*�"�J VQ9�}�P�82T��C���B�G��:s��JB���	��O����w����L'F�nM���pas��v�`�f&'�ý�ȄJ�2D}�x��!�%B������5�pe@�" ���A���|�k�C�s�z}���� �a�;����16:eJA3�����3�dY #����т�J����\M��i4-F嚇�;yZ����T�y�9c�}�v���w-��[���V��w�U�o��|k'Aح�H��xx~���l����D
$�T��￻���V0�(������8�d����_|���}ߙ̚�S�qk�m̶����;�;����h�y�i��H/>�-������
q�+*{�~�P�82VVJ��}�8���>�W̠�������F������s{�\������ ��=����%#*�T>�h�� ������T�G�>����|+�w���3*bbd���`�WםBȲed�����g&�*�ך��|&��V�;���aXPaRT�߼�Gq
�Y++�;�ɨ������w_������/ ���p#�<5����t��^�I&w'&��['=�����������w4@wΐ:�����h8<`PjA@�߼�F�R��H-ם֠)�
�l�����>ߠa�}�=�6Ό� �D<��y��pIXS������ɒ�r��8À¼���4¤�T�g���q�}�����^�G�8�YP,J�O���l��
`V����H]��3�1���:���ۙ��g�|*bltʔ��r6���lI�}�8�R8�]{���%H(Q%`�7�6��;��9�j�d����)1���_p�R��o��ȓ�f����gj$H�w^{�CJ��,�vϦ��Oǲ!����U���l�.q�߿}���w��_��+
0���<Ѵ�B�VVJ���ؓI���t($��%)� !���y]�ϝk%��
ԅ��~�F�
B��[���&�
� VX�w�|�8� ��]��������O:������Lc��I�����# o�{�G��}i&z:#=$D" �o��#���`V�o�@�AԤ-��|��C�<|)��1y�}��$AI8D��dʀ�)��p��/d��C���{vN<ӻ+'������5��79����7�<�G���������4ɤ��IX^��=�8Ñ�a������|�;�¤��{�<�ĜB�Q���+���4	��;���(c.L�ٔĬ5���#���=�k�כ|�������H[)
�o��`i ����|��Cl�%H(2��Wf��Ӏ}S�d�G�{9��8�p�ɜ�w0�
��0�AID+���h�8�P(�}�Ǟk\�;����c>� y�,k��~�����w�y�ǌ
�����)�l�)*�Cy���"�W�v#y� bAH/���B�J�V}�;�q�#
°��w捤��n��}�{���x,��ne]�4D.x1�l�'����0��>/����N:��Ž���2MV(����g'�ֵ�.�<���� :d�2�X��ϳ�5�S���S-�nn�$��m�π@�<�@��(;C�Ug_C�?a��߆i��֠)�
���߹�Cl�*AB�>�w�!ĕ�f���7<M�������u�qHjGs쉜��74�	=J��p�2���~��ѱ��sK��a���g0��HVy�>��g+*J�{��͜@�%>^��s�i�F;f|$<
x#���W�7��C�9qS133�A�����}�h�q������R��w����y"����
�*Aaw�y���aXX w�ߚ6�� �c��o�.y��w��LϽ��@g�(B� D�3SfRu��A������{�(;C� �E |9�#r�V��؊���*X�YS�}��gJ��P�w��G�Jwo��1��5̑/�υ����L���>9B'�����AI�a�9��9Ă�P/���6q�R�u�s�k�1</O}= �R�o[�ڇ�s;��76c�F۸M��{�8���d�׽�MFJ�����~�w��e��;�y���V0�*}�w�$N��}3�P!l?�~���|�r�b�h3�ь-�2�t�1�Mo^3�w��Klu�-�ޙkmY�l��Q��U����qg0U^Pi<��6��G����~�|���A�ѯ<�v�g��^�1����x�Mt�h�g8q�
=݌�!�Xc����q��g�x�\���=�7hM�Gi:�a./n׮'BZl��I����s=6���\��g�"fp9�;���{u�R���k�xMĹ��񵬝�õ�p��.���[���^�{Un�`���S�i����7�ۭ��v2�[vN��E�qA���P��i�R�b�#��9��n�+@��e�09�p���cQ�kE�zm ��~���
5!B�;���F�H[HV�
�ם֠)3�4�yq����@�>���jgJ�2T���Ѵ8$�,��zcfp��1���p����C@¤�T��>��k=��c��c�wGFq �X���������5�Z���05i ����S�ϱ�752g|>�+���P�������9�''y�>���@��%e��5�2(�ȏG�>�o}�2�˭[�C�+
0�(�{�����������̚�oޙ1�e0���i�(�Xk���<�u�q��i��5 �}��wF�H[HV�
���0��@���;�u2�����=��1�<H(��G�>��`�Q&DL2D�>a]��rT���Xw����3�����8�ȭ��W�� �B ���Ő��(Ԃ�ﳘ
A�!ia���u�#y���cII
(��H��p[���Ғ�]���"c�vmxƆ6�ם�a�������.�F��N��~��H,�d���׿g&�*IP�+���w>|���ܭ�2���	d>��G�+%Y(���s�
�t�m��72U.]�@�Jþ�ϵ�85!�l���f˥4i�^��7
,)8 �R�bwB'��aW*%u�<�c����b7q^��%oFdI\T-B.��U�H�̅1��$��=�{���~h��B�B��]~�9����X��?{�q�*AA���n;/�wƟ�.���O�oV�b`����\۸a��W�}���T�
��VW�P��>�>D �DyT�����Y]���,�\����)
��:��6��l�.3%D���)C�E��3hY(��T��g� ��ެ���{��*T($�/5���q��T�>��$nw�J�u�y���&FVJ2��3�5�_��ьs8�����2���5��������@������_$ǟL��m�Zc�kP�H,�=�~wP�8�YFJ��{�tm	+�����u�y/��ܽ��x/D�n\�\-�mm��G��*c�Y��θ�kl&�����z^,�]k����;W}�90�(�H,>�}���d���}ѴD�������|q�����>}��R�!m��s��y�9���K�s�ź���I���tq8 VVJϵﮱ�^.><�-�s�pd�T�������Ì8¤}���i8!Y(�ɝ�gk��g|��y�s'�Tl����mÙeˣh���s�0(ԅ�{߽Ѿ�AQ�����\�����0*߰��K�1=�FZ��g�a��}[f��/oWW�`vsW|{2A@�Y<�Et���j[N��Be����-}�{� �z�O�J�X}�=��m�+(�P��߽��8����l�\�mqbDJ� �3�������]i�TsǾI�*J�a���4pg(ʁA*�{�vq���Z��}߽֠g��Zx�W[����!��}�exY� �Mj��L�&ba%�YG���i�++%~�kF�J���~=xe�߿o�0������p�0��}Ѵ��VJ2��{�jM�@�����ރ�W\IT�PD� D"&ax��b�.�d9���5�����f�3��pV.������_������H�ַ�t0+R��߽Ѵ���+X���w�
l@�u�N�=��������P�8�YY*�߽�ĂÞw��e���\nag��ʠ��#���6�1F��|0�;�4z�$�����h��,�_|�����l�/���;u���q"=��RO����^V���a-��HO�O���tq8 T���_|����*%`�u��O1��}��q��H,<�*J'���4q �q� ���u�6%@����ps-��T�vq�Xw߹��������>y�CR-^��to���!Z0+g�{���*� Gח�xY�;�_/�R܊V�������������˘Di��;�	{�Z��+����P�d�t��Ar�k!���.����|p�m�ߋ�<��$��q���P�|��tq	+
}�^3�.0�L��a]y���aRQ
��Xy����Lw������ߑH(η�`Q����� üߝ�8�0+ߧMeH���ɺ�O�-PJ�ʃT�n%��]7!���ۥI66���yK��]�1Γ����71�g�v�9��}���������oߵ�l�T*J���~wp�F���O|���=��<����q'+%Y++���Z�iP)�zk�Ǡ�m6ibVߜ�F�9��p��u�Ͻ�F�)JB�`W���j�@�P+�~wP�8�Y_y+~��7뺕�Z��@�G���љ�#�&��6Ì+�s�h6¤�B��7�چ�
����zU�|�\�߾�_ u+�X5�]�Z��i��w����8빵��#*Q�������d����Vα�3�� ��}֍�T(����{�q��T�1�{�I�s��g���v뾇̛ed�+�;�jM�P.2t���Ìd�\�8�X{�ѩ
����4o��9�s�s~{�:`W~k�� ����7ߵ����d�Qw��!ĕ�����0�ܼ���.^d~�=@�Q�����	���D&��o��>q�T�;��ӕ���?z��"L��جCa��sz�k}����{��X�>8n09L��!pT���Q�`ݷnm��vn��s��:�%�BnR��nsY�L=���Y�H��?�w}}?U���75A���:筶�]�:��r�紃v��7��^�a��R;v��+p+.��I�q�pE����n�Y�[s�y͞]��A˗��g������a|���t��w))ϵ丱a���fe��F8W<w[ ܜz۝o�E���mKٻ:�i7$�X�B'+��9ݙ.n�j�^��G8;E��?�;���y3�[���?��u�~փq�IP�*��ߝ��q���X%@�>�y��J�l�X�Ș�ߟ�&u��#���u^!�����{��dxce���H�fd��Y ?��F���N���o�T_]$�u:I^6+����E*���=s~�`S�$(�����������'ăq���yS�ꪝ�y��O<|�$���o���,�J�!&:��4v��$K�A�����n�~$�rs����0˷L�l�IFJ���%M
y�� �rw��9f+UVf��>Z޶	�#���d���!s�Uϙ{9o�j����鍰�\h<nD��v6��5ε4g�*�o���|��-cc'�������|H=�LI>�Ρ@���3�bjF���F�9_�t=����x�Ɓ��"��q'�s��H��8�S�(�A�zWW^�*�a�Å�JnY�'J6�v�J�qu�g�oY-��os�S�i8B���1��o-��A>'�}�0O�N}>��8^��Y�{���<[a�i�l�=��}($]��@�/��OU����2;^���`�I��p��������S%}�D.�2�_>��$�<t�O�$]gW�����{���U$8Α6UDeݷ�yfŕ>���I�T��$����ŗ�NCFF��� �r�������`�e���T��(`9��d6�l<(��9ᶺ^R��;��v�r	�=[��i�4�������IP��)A��V��~'���oH�뷬m.n�)�s6oI���� �gH�q%D��HH�M�����5qnO����ڧq�XI �vȢ��m�	�&�:�H�*���{2�	�`B*̯��$�w}o�!
����!M�h��u_޻�:���W�`ʧ�f����U�cn��5t.�WPzA,E>&eym����[�c�{
���Y0�&y���e����m�{h�,+j�7�"lx'Fh�R�]�h��'xn:O�����^�Eܶfs76���ҝ��Abb�M��]*�I�kw3�y�w����I�6�L=CS�_�|zR9$�'��W���Y�ŕ��AR�r��������W˸V�������T�ݹ)����;�"s�n�Ӣsۻ�P?�nһ^�R�o.�񛽕ܙ�)t3OH
d(i��o-�N�P���I�t��_N�J}D����̸[y���F���ɣ��nfL���W���O��rfj���Z�L�.�!�#��#������'��t������PO�V�-b�>EO��$�V(0@�mc�|�-�y�]�����d�oO=����zˠD	��Lb��v���@#�/�!��I�|��xN��K��P[{����Ú=�����.Kvj��b��p�B�}�ᴥ��t���R��BK��-j��1�J+{�bt�[M�3vv�����Ӷ�l]&���Tb���yA���}�oA���Gh�;;l�c���D�X]tZ�n+S�^	�=����j�\3���d{G�N��7�!:�#���O�G�yv�ב]����ó��c&Q��p(�nb+��"���N�&5F.l��Ƚ��3=�����R���F�S��Β|'��J(�F"�<1E�`�҅B�-QTQQ+R�ō�V����(��"�Yc�X�
	iFڌX���ڊ*��V�Ţ�X��U�X1UQTUX���E�P��R�X�"���TQp�"
,TQ�"��V�W�(�UP�b�R�DEE�h,b��Z�X�VV��ԫ��Dm,Ũ��#68�ũnE��qeUE�U�`��1����.(��UR�X��c���U��lUQTū��Q
Եj������)�QL[V2(�)DdPf)U�*\ZZ�QS1J�*6�(�
�Qa��Q��"
��%ja�UZ���E��,�U�*��F�Űb��b�V0�TDT������(�qj1�iTP��h���!T0�RƬ�UKFҴqJ֫�TX[X�Rه
��Dqj�bK�(��\R��"��i-*���TR������(�T�Jൈ��k[*6؎)Y�Xb�-*��DDQ����,A��*���@{�9���{���9�����ZfdJ��Q2��c��]c4��Ƒ}R(�E���=;���������f�k$�� _\e!Y�L�X��辤(S����!F�⽑�/;���������d��c`��Ne�&u�p���n9Kn�̸b�� ��x�Z�qׄa�awF;r�u�cK����7�ϛ��;Wn����T�q>9׶�� ���l�bt�� 5s�����6z��%B*d�
&��c`w��2��\�T>���h?��o�i�Ozm�l�f�ݜ1�T-Jd�DJ�{5��ͺ`�x��hEP��}`1���$�o[d����H�
&f<h��M� ��E� ���~�hz��P��f{�{ٗ|��ۻ.k���VZ�N�x�2����ꮾ��
���3!5��ҵ��I.ʽ��5�ݪv0�U�r%�6t�[\�$��=��_����ߏ�ƹLȕ
d��Ji���ǉ��٢�5��fV\G>��$�tv����d���ƹ^�T�	"�_�˝�9*7lu����]uh6�˳ h�wmغ��;/`tȘ��T�3Uz����f�2|H$egP�f3cgZa^m%��� ���l��7�R�*J�L7�܊#rh!`�GUc�����$�Vt��YWґ٫B�D�L@Q2J�b�n7�I9[�^$��lp7'���\̘�u8�@�߿v�e��	D�xi�8���=���֯`�	���d�V��� s�λ"6\Ś�t������2�X��k��ߜ$���۷�����vౕ����٠A���6t���k!�p����u��ozȦ'y�{�ޓ�މ�����g�^�ީ�c��<�5��:�7}����%��bnc�{��\vؔb	�`�2��@�S�������zv&�7$��v�uϹ:����!;/"�;]9�s���#,4����B�6�İg�qs�n�4�ν���Ÿ�c��A�����8Yjn�{kqX3�Tun���ܛ�S[����79��[m�^^Ӷ���VVkOF�,���y�z$y���U�\d�3��[%�q��wGd��[�M��!�6�����.�6�ϵj:���{�5��ݹ���Σr-�����bL�S&&RS���l�A�͚ ����`�Y��Rw�8N*n�+(w���E{sߕ)��	��[��t���i�{Ԩ���r��"纅x�O���dM����D�M�{���Le��X�����
 ���vI��6�
$�|� ���zh3D���+)�1�{�މ����� {/Zs� 9�� 
�}L�GGv3Mqd�Y0�=��L$�c�3ʡS��S�f�v���A�nj�Ù��]��Mc�j
�$����H�vS��A����礒`HPL%10LDk�����Wu�uYp]�q�2)�M67���r��,�/�����LD����%[�,4J�Y�|�ZI/$��c��8"*���L\�U��� H�^����NѬ�����&�(me�P ��l�{�����[>���ֱt�P=gN��ZQ�R6��ƅ��thJ��ef��Z}Z��ؑ.���w,�Nn�e�� ���t��"Pw�����G6�"���*�zw�[�ӲJ�R
k�)y�K��j�f-��$��o�0w���
��g7h�GQ���Ũ��D�JeTRm-�����k ��U]�D�^1���~���{)ME����Z��(0ɐ�ES�v�A,��G0Է.����X߹��$�"a骰���}4��֝a<�]��Ј{��!$?^����H꼕8��:y k�]���rQ3��7�$�����ؿBmÎ#�����:��:  Y���mmP]�-m�Y�ͺ$�&M_a5\���,ZR������ll�ڤU�C��v� ��r� #1�y��ܥ��ڪ����	NQ���D�ATAC�c�bT"7ס�{��ia��	`g�+��;��(Sk�7܆��5�/M�Θ}[��a�^��=�efՑ|���Z/�,�{��=̤�Η+£m���&������wo~ h���D	��S`��"���Ң�6�{�I�V�;N�	����r��[����3n�3�\v�PW ���P^ݑ��&�S*��h;�t� �����ϔ+���-v�z_9a#��6����ۻ73^W���'�s!`��h,(���u/���:�͸ƞc\����~��ϖ99�Z��|<7���9�4�Aٙ�v�j���Z�y��(�6Ǎ� �{M��aQ�0DLɕ
��k��J����.y�A�{�@�@o>󈈎�zށ7�I���]]����hD�"0f~t���M�3/9��D�w�N���p�"�b�H��<H�I>�so�	NQ�u���j�(l�/\{���QfcA�y^���w^kw� u�e���@����r=���v؋��m���e�{L��7j���]+������v�/���G���a�zg�7֍b��y��Z]0�g�� <�xU�-��i�&d�"$IR)����ŢPK%nTWYU}�P�m������[��waF�j���D�_/R"X�!�{3&��&�<q뇪]��zY7��3�q��h�%%��"�~��ĩ
��]N��0 ;o5݀ ~��s�ۊ��v_�a�W� -�λ��n;��J���Q/�vn7@�w�k����n����n���7J�:}<Ƞ����럳0H��!6��ǫr���j���ny�/��.����ob}��� J��n� �7��nc�)U��
�����Au[�����Y �����}N6�꼩�ym�7>wwh�k�M��*��j�(me�t ��i���n��u��[G��
�뻰> ��cix��x��Aވʭ��ԏJ]EÜ*�v���wO�zp��T�@��u���鑖T�K�g6�]�0�/�SţtPNI��E�3����ZY�����Į�� {���߿�κ3�9�<mWd����7��\[�7Oa;w[�"���9�)��v�'n8-˷���cn,l�n����)pm&�8�y�ۍ��y���%�$�]dի;^�n���pn�L.;Q#��Fs����Rl�٨��n�w��5����.���`�=���CV�K��n�<�*�u�{v���s���Ks��{]u�V��n�l������-�&�C�zՑ�����c͋�����
�{n���{�m@������:�\�mw~�7���'�M�դ� 8�� �����I����##^y���v�*`�2Kj�_�^H]^*���.%US׍��D�[X儉@+��m"�\�!�S�2�ou%�V:��*	�*AD�48��� m�?�D�H�=��3�w�do��x����z��`�"f`��DK��kv���V;����k{I�M_>� z9͌�#8_7Nn�JNU�)vc2 HDǦL*��a�ަ�|��y��{Е74S�8�[� ����" ��ۻ	���^��9��N|�\M���Y�m���64c��N=�E�#�����rO:O���|�Y�>6� ���|�.�ͻ�Rnw�N�;��Q���ߩ=��M$�qtJ$��
I�ʚ�l�J�`�و�ѐ�oLHȚŊSD'�_C4趻1`�z��x��?O2��Mu�/�26�"e�vN�,�s�p5+�:Ϲ<��_�@�8��5�{m�{��n��36��1��}��kg�i�{ݾ��&f!SD�2;-ʹJK�3]�� �wB�Y��p��gv� ����@��3n� w�>���+��֯��'黮�I٢��O'�P5�S`73n�",��c�U}Pl�+�\�B��8 ��RI噺�����}�k���;W��L�:���@ vg]� ���6����^���S�?/��+�ݨ�:p��+����Nݧr�m���\M��q����Z�??w�z��0*I�ܞ/$Nfg6m"W.�X�'o��C��}�g�r<@L�rL�#gTI��1&B��{Y�H���ӫ1����vg]�Z��g��� $�����<��ښs���艁)2*T���n,�#��~ >	�{g >�~�Z���h�F�J�*��QGa&�լ1�@��3&��G*_mۧ0�ghnZX4���4����*�j���{�K�ѿ��3�� ����5�v��LB�*L�N�s\V·z^��&s�O�Mh���lX 
��ش:O"��>�7	=��^�xKԜ��!��n��"ZMh��ؑ^�bJ�m|Kz�&H��lKH$��WĜ;����Ĭ;�لB�d�/�6�Ǆ0���tc��%[�;/.{i��Z�*�o����|�.�B���7��AѾ�T0 ̾�p��uRgGi��yfz��� |do��I��Ё(��2f��w����G{��~�3s�� 7��  ,��d�y��9��6�n��	FF�	�FbL�*�{X)N��4�&F�����@ ���7����63z�M��/�1Oo��)=!�U�F�gz���}�{� ��ێ��#ط&������tü/Ũ"��(g%�0W���z��ў�^j��o;�qa�R�×,�yuAf%X���� ��O�u�/ٮ�fb�P�beRm���� ~���ޗ�T�1|-pG��$�h�;$$�퓛a)Mh�肒�fR�bJ#�a{gӞ�D�[���v8x�#�u;;"���R�~|����+�T��~�8�������6D�����'�oq���� o�i�(�ND)��T@�&i�:�v�X ��A6�3}]� ͛�@4I�;PD�M{d��&v��.;i����%}�Б(��1$�1{թ0 3s�`�H6��{!�wX ��l ��mݤ���&	��!J����J�kF�����O�� >�y�v� ��U�q���{�{M��3R�R��
RF�~h?�$�����-���ٳN���}��5�7h �����?-��^��o��Ma`޺Ƅ���gw>��3i���ȇ���6�_����xj|[;�7�gal�c��������}3xwwm9%8v����wQi�yϲ'��JOVӫΙ��(�U���#$��u4�N�x�v�:�C9�mL2E�Ǽ)���^^u9=�>co)�QJZn�}��%�֍n�s=�\�̄���
RWS�ȽX�&�Cz�`y����]�+�A�Vr���׼r��/�,D��J_q���<gIW]5����랇�������U;>��䙤�Ϋ&0�j�ۢ!ݻ]v'�&�B�}����A3�Rw5 ���k��U��e鴗�t���&�Fӳ ��p{��$��Oj�������%3��a��<o��l�\�����΃����
h��� �U#Q�w�\�`�Q�=R�-^�;�O��=�F7<_�g�v�r�j�C�4�q3��2��qW]�j͝��8ӷX�Οv��t	����w�����#��d���2����'e%Ȼ[�|����R�up��5ۮ�XF��dVWI���R�ׯ���;��vz��~��,o�U����M���h~{���iĝ�b�BLsTN·�-�a�1�6�7v�x�%rL�yN:I|e> ���;n�ʖ������o���w���]�3K�!ۧ�2naڐ!t�6rgPN�Z;�]d���ۙ���J��S�o/%1�ī�9v��JeN���y����d��ts��ת�o��9����w����L����LN���]͸su��&[ӳ�}w�r='�ثe��]��4,b��Ylm�QUX�1*��[H�0AUf(4m)��R�"����UF ����R��5+�LZȌ ����`�UD��H�iX�X**����Ŋ�P��[lQE���DEQV6�+R�TH��6�cR� ��pZb�(�e`��V����X���b�,0�hV�D�1�&�8���iVDU�"����#ADEUX5��R�[jT�$qk-*��qekV�Z�DV%�����Ŋ(��*�B�UU`��ċl�qj���+
��*LZ�K�X�EVڢ�*��QU��ŌL4e��eB��`�1aQ ���-��AjUE�"ֈ�-j��DPQ��(X�m���*�����U�*�Y�* ��\	Q�ңmEUťTb���G�+T��Q`��)Q��
��(��k����X�aR���5*�H1F(��EX���b�D�
,P�U"��eT��
�����������}�!5v��M��r�x[�ywq�H���&rz!���Ć�{l�k����n�[f��.�}�
$i5�7�����;�Ӱ�!��l�nֱk��mr�x���������nN^ښ+��]�!��9ny�k�c��{U�<r�c�8���+Fv��X�ўkc!X��v�s���u�����w7n�6�v.W���Q�<��]�Y3q�i�n��s.���{9�C�X�@*T��5�3"�������pl[���նp&�����<��{6]��Ų�i�q�c�X��V�z.�&��������;�q�Evs�Ћ������l}p��q��v���ͱ'Sz��/T�z��m��]�Z�<}a��랮Ӝ� =4�ځ;�>���z(s���k��xt�:��Gh�����5�88y��\�b��G���$jŜW�=6��PY��=Y���j�a�v��F�uxqtZݺqogd�^toP��1��$�MҢ�ٕ�hݜu6J�!�hz9񮞝ƧJ�.2�Ƹȼ�u����p�awgH6�J�n��=��s���k�ٲu��7gr�h�Y���w�ۉ�\a��`�b�yp�k�T=�a�&Q:��o9^8�v�D�%��6�`�z���q��1^��{=t{��͚�ͽ��ս�y�+�7�M��2%���r�v��U�GN�n7k����a������3��;v��-��������{3�s�w x��{Sѧva�uח'O;3�v���%nX�l]���F<[8w\N5=�-Z%㶱z�7�g��v�Y��u��z�m���0�cJc pr<��j���\���C��z^��˻#rlP���;����}���B`L�gqs���ov�Zk�m��˧]����v�S�Hs�
yݏ}\�}T�_,^,�(�R�N�[۵��N���ڴ�g��qe����lC3��l�v�5���G���Cn��
K�����e��:7�ZL�p�Fj� ������W�]����qI��;�a�vq����s72��u�{hz.�x���թ���'U�un�x]��fƱ�&��q/j�L�e�l7N�cH�C^��gZ���[�sg���Y��\�Ն����u��S�nj�EϬ�d���Xn�U����s'H��b��F�Na_ex'�]��ם33���=i[{i�����^�t��ګt���w=a�^_u����y"8�j.L;u��\��O�Ʃ�>|�o�)��PMD_� ��` g<�v �v:`{��~�+��|wxǽM���y����>�*��
)U��E�6� -�T'k�V� �y�w����o�I\�N-�����f`y"�F�2�Lӧ��o�n��]�~ ���ѥ��`�v�I�K�s`:$�|3ѺJ��2R&=2bb��ޔ�\�{��A�}�Ցҷ0�gS���_A)��j+�n]�	��U�J�R�UR�<�:.����6�e��ש�Ju@%�Ǘv�@|dWcix�"�:i�(����떢
[v�H"p(�&���Ns�q��O ��bݸ�z8�r�s8�Ͷ۵՗���ٻ3T�R���1J����� a��~��I/]gS$Ƒ��U0߇]�m��z%�i�l�9wF�U�Q�Rn�AP�D����°=y1�9F�"�W	��s��m�t;����6]�p�l�f0;e
T�&�(��U�x]���:�e�U!� =�Y-���  ��"!�=�����7�o�]k�ή��	!�0EAS""P2&T:j��7�D��ޚ,$�H[�!q��N�k�Ȯ�5��H�gSaQ�ؑF"P�����k�^�]uD�8�rw)����~~ 	g�|��z�W�bŤ��}�N��"%�	&bT
�a�W0A����DJ��3�*/�� $��ΖIi.̽�$��2�!��:�����n���6	!P�qp��$��Z(Lu�"�YS��:�ȴ|����ݗ\�uv���*�&��=��R$�=#䀘�"v]&K��"�Gkzi���j��"L��!��]��H�OlL�Q��g�7o�����0ve�݀9)�������k��G�D�DĒߑ�h�I z0�N\�����+<��[�������<�':?{��9Kb��Z�����L�sY8�����eY�3!���������A!��o�����ۻ@.w�>�*��Q�P��Q�Ǹ*/H"��(��ޖ� �>��ۻ@ ��]��UϺ��z}���ջM�G�p��R*�:�ݻ�����=P{�,��Ȩ��πKw�� >��m݀���DY��#�ğ
��&<(�J��<074wm�]=����b`���qr��k�?��><݌��Q+g��z�" ��sqh����t�k�M�}G�� �L�m�o�M�F`ȁ2&A��\n��a%�˷�'ћ5A箭0 �g]�DZGEv7��gk�4�w_��4e��bl0�h�i4�6��2;���u�B��GL�vdo� 2�6����}m���rcK�l��3~��w8�ܻ�5�>�A�y�� @q��M�E��{ٖ���v����胤A��zf��=l]�s��j7kk
R���%�ۅk�o���1$z�Н�.X.A�}x�؜�]����������&�s������j}0U)�TK�=��� ?vU}\%U��&*s��:v��"�I_lc~�w<vd�V容��"r�pTS�-vy�w�!�.�n'��h�dT�\����33V�I	�RJ�MO ������@ ��g�^��w��m����Ѫ�"V�]�D�-;X�%�j�	$TPC����iЃ.v���u�y����D�:` _l�) �n�)�:`l����Q�J,�0d@�UJ(l�w����8Ӑ�>K���y�|��@lo����}������j�)����i6�>y��uf9Y��_� ���4�|�:����f^�ՍdfI��1��Rw��Iz��b#Ӏf / H�j�VI$��䃲:����
7G�
ǜ�!��mI �/m�W�5���D�/>\	���7$I�3z>���	�puY�0���r��+I��ڹ&4���J��z����N[��<�&+~��<-N؉&9��С�ջ�c��n����a��;sa���:�|�O���֒�d�f#i�uϷ��ϰV6��×�����Mk�n����ᛕڝ�̏lӶ����(��r�1�X�qɳ�8h{x6r%���u�y�10�[���<8�D���O�v�h�ľ�pm�vS��z͑�`��a���� 񇎳���` ���n�uy	�Q��7 I�Rj�<�)������ �����ܻvru��f���J��h�12R�(�[?*9�� ��m�@�z݅�V�Gե��u>���}���~jJ�%�*�)AB��p{�b�@�_h��f/q���I�/6���H̽���?K}��D'7*���#�^P6F F`*�9�vhD�$~M�D����s�<��~�!�״� Ko��@)��\(��R�D�2�Z]�v��^���a&R�%��^��@ ��m�t{�WY9p��s�4����S���b"E54�� @����P�|[ھ²j�@^�w�D4��7i ���6�!ˌ�\᱿��g8��t txӲG!,;��n�v��2�i-�<�=sֺ^1w�����*�nٶ��ps��,$��n=w�D���t�tDEuzr}{6�=X� �&�E��~RU�"f&L)F
r�ٍ����fm�WǦ��g���TO��`�50���ꅙG*�=�hk�<�X�N�嵯�C��葓�15/v�ua�#��/����e�� �����>!~���\T��}�'ӎ�R�T�NX]��l�I�m�0�$��]h���Ũ"7wm�� ��L��S
iA$Us	�TM�_��R�[�\�3�_.��  �����#��zk[[n�`�3�׸�W�B
O
��y=�����I$�����tiQ��n����m� ��x߈ 1��a����;"*~��o�{��}H8��; M;��X�\���5�=pz������ځ��|����.V�yKy�ͤNyN�$��;\?$�;#�;�^~�� ���sxK��~�M}� ;
Ma�Mf���|�2y�S% �Xs�L �go�T@ ���U�m��Ɓ��2���`�{>� O��X�u\���}�~�/�L��'��,��2ڵՋ��1���r�>;�yb#�y���V_���J�}TV�SUY%�χ��_7���K��v7�����A>�u*���Bb"Z~]��cp���2ewl�"`�?T0�f�_�v{6�k�t��߀�O3[�����4��� �1����f{9ݞڅ���^̪Y��o_���5�C@%}�ۻ���1�~"���dX@����	�!3�K�n<u���g�Ϸ%uח�$������͡4Wh��w>�B$�Oa�K $���l/P�#�*~�舆]��_r�h�Q@I���]� 	��o��κj]��Ȁ��c@|���݀�?{v�FT�R]���C1
=(���%�%�p�R� ���� ���Ϩ�=v��� ���dC�۷v�̓�Q*�L���4*���D���$�㛄In��v�+�ug<��#����غ����֠���-8d��A��g�)O���f�M��^1
��r-��wz`�1W,nTD���5�m|��~
����(�td@2�`$!DKL-��tH��ک;)�AX�g"!��}�w`.�o�dD�읊�{�x_�GE�£v=e�F�����am�������D<�0��7y�EL�(���9(�~s糝� >@��}��5�w���D0��kvӵ�6(�U*��e29��8Qq��2"��tf8%$�=�w` ���d������;�fh�T ���ë�����ev�� ��Jɩ��[� ���wM����]OT3�ҌO��[Kmųi�;&mc�$�q?��I�H�ܴ��u�w#��5��o���>�o@Y���J�"bDN�{���D�>�wG2����.ݩ&Euw]�I"6{u|� ?.�_!yՏ�s�.��A\&�!X3L�S��}@����Զ����;�"M�3d�}���Ek��j#ƙ�������
v�D��{��ۑ�*�@F�sϡ�t��cz������01�+�o��'N./N6�c����;@�/���v����d��qŘ����o���8>�8�'>תH`�U�W�.�]�����l�dt;x�iW����[�r����ڭ�tpv�G�@3�y7��;-����̻7`�R��Ǘ/�=�Ool�G����Wn0��qƶ��;Q��#�=�Ƿ7<6��a��ێ<��9���#}�� ʉ�B�:��]�v�H�ӻ� ��{�����5[8i0�/Տ���uv�C���`���EUZ����$@��#�m�\���~$���Q$�E�� %б|	�0���{�����,Q*�D���6.w��� ݽ�ȃ���6���k$�}�#Y��� �#my�oi�4J
��$6�������GU�)5���Bg.�H$J���d�䗯��ٝ�%F9�|���B�{[L[���©������4��;����gM��^� �;t�I/'���-+�|��!T��3k������-��`�ጛ.�s�Lu2�q����N^'��=�w��л�����n���aP���x� ;�� �|݆��<�os���S���� y�M��z�Dfd T��s����w�#(�?طs+����8QN�b���zegt��ڳ�{p�eND�����A��=�v(C�S+�F�^����?�oj�j�������i$�}�4XI���}vM��\o����^o�B궠�eJ��&C��Ot�%��-�h� ������g�����C@���݄�f�hB3 Ę�4)�3�4������ ���A$-��.wϰ��ygUD�>E�u6�tb�0
��$fC5|��	:wi�t��P��9~� ̷�� k���uQ�{h�D��E"f*R&x�;�u��y�[���)��u�]]��;65M���|~a]�)���/����D0���� mv�4�����y��>!��{��R@ז���@vf�B�U*��T?1v<mR l����tۋ��+ �k�כtI��Cz���Il���MEX��q���|�_J��R�eL���۴� �w�̀USС���JI�w������1*ˣV�i�u�d!VQv�-�)G���-o�Y�Oާ����yB�:��{�QcX��\AT�݌���:���!�gWs���I��xO�Gu��k5�jne������}V���ݛ�J�+U�w�lJ�z�ﴧ�m�T��#�)�54�RR�����X�	�ۡ;�k:��v�ki�s7	���j�<�w�lE1��-�����a (S��o���G����L�MK�5K���� ���v���퉴oP��Y��5ss{��9# e�����86xq#��Βiͣ�v�՝J����Z�����!�n|��\��״�>��"D����P��uodm!7��Nj)S*ku�}C[�P7q����F��t���uʂ���w�p�f�Q�s����9d�8^�7�j�a�х��rC1��N�eZ�ڗU�sP��7YG�blz���͋ӭ��e,��(����`fXT)ꊈa��w���/uv��u�TB�D8r�93���v�i�-��ֻ7!I��]���Ƴpb�@V2�c�W��3�w�o"����׈2uf�FՄڥmN���I�"_f<2mߖ��i�ֵ�N_N*�J����ejeդ�[,�i��������ɺ1c���WN���"�~��ߡ�-�%c�����Y�-���"N@��spM�I-Ml�gi���)�z��2�8�ugOk�)��y���5��c|J���{��������q�'�>$�*Ƞ�تJ!X	h��!DWEUF(��,P(0QPU�d����+�V*�e�Qc[-����V%�b1b��*�X����J�X��T��X��QP�(�T��#J�TE"Kil��Em�DFEA���QDE�*
,Z��EZ�QQ*,TQX��UEC���Q""
���b*[Q�IL5X1* �L5`�0D�H�*
�b�\6*�*T��U����kJ�F�Qm��(��*�X��ֱh�h��EE"%j
�[E1�V
��m���(�֩+l�
԰U,U�cmJ�c ���1Ũ��PZ�b�UKh�*�
�E��"��UY�Z��UX���QPX*�ҫR����6�R��J�Q�b�jET�0*��
�Z�Q�PX�EEEF
�h�X)P��(��b��E�\Ye�ER3TQcQQ���T����ij^�}�:���m<��.� �����O|AJ���U&0�����UV/?�A=��`� Go��� ���DaC}N������Y1@.�v��gvl&	�����@6���~��%�춴�D��	-�λ&�<z��"��	�l��H��ΒQ� �5�q��;�ݪ����s8�^��nwV�4�]�^�HT�S5-���TJ����Wìܻ�@|����|��q�]��r�z�����z��@ ��z����g�L�%"�&��
ۺi�uo��׹��K7՛o� a�]4���m8���3�y4�ޮ�}v��O�
IT�jaP�5�䰒'��D���'st=�uW�I��{O�K�٦J%��*b	�
%��7��詼R$>wM�PIy�u2I,z��.�wJ��������]��/מ�fX�0]X�[�]RV��m�5���������r��O��jit�\z���3,ǔ�<�� r� |�~]����:~�%bd� !2igW��I$���˓t����&LV� ��8�`_{n��	��{���?g����lQ�L"fc����S�l򓗭�	����;�y����>Bq2�W`���� 
{�R&��I����%�/�GU_��rI/��[	!��&���#2No�ٰ��rbj�j����	'�9�@�%�y��?Q=�V[J��{��ޡ���>��L"h�4�t�
$	��d�D����Yk��t㾢ﺛA�+�m���̇>Sd��6�GN蚞~�2h�b{��A%�v���$I�ڪ���p	%*|����#)LD(%�n=�b,;nw�H��zwoc@vn����wk��Ix$��n5�TM�ޓ7٪�=����J��I�i�Г.�r���o=V�	JZ��(��;3�%5��l�'fv$�0;����6;~o�<G�p$[d �v��qd;�lnw\�)»I��ں�۶9��� k��l�43���iT������9wmkW=8����l\wE�����x�Ǜ���q�C�`:b�^\s����n��yM���=�1�[��g��Зz��;�j��1��=����7\��ݴ������֮!u��Dʩ�cY0�Î3��7�f���]db��m;.ݮ�v�/K��q�<��R6^�ra�|bv�zېl�q�k�?>~�|ۍU(�Z~���0>�x�Ȁ]��'7:ݦ�����k� BMOr���ۢDT��QT�G;�n@9�g�32"���ba���.�Ds��9"!�w����}�*�t�ޜ��*�����M��f[� 1�7�W�8���1"�?]�a�$����lD�=�mHW0^�
&�D6]�l�,���{��� @��n� � ��k	 ��m9�q��dDJ��ۻ/�D��52W�?4Vl�!����M��u���k�E�f�m�H��z���:��H>�m6�u�QVW�����?�r�q����Q�X��u��k��c>X1d���c]�;����>/kG@�b�>w��ٴ���~��IWf�t�	�-C�7{�v����em���*�P���I�,��`4��n#`��e�Ň���W��{w���F��'O�=]2B4�k�=B$̘�Tu�����x�Ӛ�N�"�H�(�?��<�s�ZI ��i�ZI}{��H��u�73��S���HTf��D�L�R�IE�}��%�^�4� z�.Y~�eWm�` �i��u�טv�z�*��J)U�O^[��rz���̀�.{��~I���8`|�;����f@@�z��|UyM��a���@�����=ɧ�"F�XX0�3@���M��}���@��iS׽h��?������9ɗ�����W������@@��i�!"�w�=���$��z~l�iH k���"���h=����{���Q��~ }��S�=_B�����gf�ڰ�5{u���ə7*_�H ���o�4 
����DN�i�e�����6��|ISU0L�1�g:i�g;w` y����=�R���6T��cp�����Y<�H��`T��E��������b�����l:���.�2Ľ6����|+�9Îk6�n=��WJϜz�|�SY�g�@#~���)+��6M��u��&bf
2Lf�:�����$tE����͖$�'(��=}���ԉ �V �Nx�]�n�ȁ*d�2&E�z��$��m?)u5�T����y�p� om�ݤI���p�=��Ȃ	��

G�+ۻV�ɹ���{n��y�ys%]e[v+p�����
b&i&���릓" ��d�&�;?3�DˌL�0S�]�^���N�޷��ٟ��l��'�$�nC;m� w[B�I&��fy���I������- {:u�$��o�=z��\����A� �D�Nmֽ��^gN�� 
�w�+��U�\��Ό@ 372�"�ΝmH+�k�SU50Pƃ��S�Nrt��[۝�i ��ƛ&�$���� r�۪�ׯ���]��-��<�+��3#���S�}	�=� �>ļ�����*<|Q[ߊ��O�o�������I��*;J��Ղ+-�ݞUj�a�I��;�m�vM��몉TMM!UTDÊ���b�@e�6ml��+o��]��vM�#=Ѵ�����A�\�ʉ����L,��!<�ՠ��I;ɜ���8��W�<`�z�[l9h�芉2wx��"���L��On[7��]��H >.��8h'�;Zd�LjZ�n��@�:܂�\{@����1I�����_E=�{���~m������X�	 ���l �).�u��ѵn+��N[��i�	/k��HP�J$�������� �ݚ�| 
ڙz&������ N��r@�;�i����	�L*k+�mهv��`[ӞjA ���h �}w�8�J:x��O�vTsbz�yD�T�L��h;��L�;����=����޼�c o^ӈ��V����%��B�Qx���L�i�W�<�ɧZ���Ш:^9>^�PlfOQ]�9�ג��g���������0�U+�O`I��f�'V�lGvg� L��L�"���Y\P]��� �u���qΦ��w=�-��n�ƽfdv�l�n4A�׭���c˵q��9{WD�m6K��<��VϞ����9�L\�c���u��ݝƂ;p��6=�=��5v��c�m3\�ݮvys���5/O�|�n�N��w�5������`ˇ[Wx�벑�S��{�l�;]o�m�7m�o[֮�[�뾭�� �ݷ9ﮧ�ێn5��M�{o���9�\���eᵹL#��Pf���L�fB2L�*{�%����M0��������l�w���m�$D����n�*����UI�e>n05L�[�W����  /w<�
�k�� ��v�5廍M��������j*�2HRd2j������׮�"���0�V�{�� |f�S �}�wa�pꠉ�)M}S�4_+��皽�����X��$���M +:u����]q�#ۙM���mW�� �D�e��ͻ��&s�|��=�'f�Kȋ��h�Z��p�{�݀+:u����������y�Q;y
���8�n�h6��0'g2Y��o[�F�4�GyD��I�J"U"^N��D�_c�� H
έc:�����q��"��6�@���ۈ��uUR�j�
����
�G6!�Z���pL�-�U.�e�H'�V̧��t��GR՝д�8��ш�V���:�K��¬ůu���VD��6�ĕ7l��r�̟�`���n���[RA�q�T�J�{6���YrL	�fb$D��Nv]�@DV��� {���yjo�'�1�o^�݀������=�zcH%E)�B�!�$�٧�7f�o	,$��Z�D�u���>�جOM��Z�� �{�wib�UT�)�k�y�^����@u�z+{�EǷ��m ��wv���gY� ���T����>�����p�<�j;]r��{(ƺc.�ݸ��ݧm�m�)�0bS��ޟL�B�d��s]��"���|Ԃ�m�DC��� ��fr�vD�9ѭ�^��+�&%U!3����]4�^��^���y���"vֱ����!���2=}��vH�5��w��B�,���XO�ϧ� ���$�y<���ΠB���4v�����u_N�3����!�F,�]�[��>�����V�v����3�X݊��.�5xk;��I�n~K��ܾ�� "�~�o�
�G�~Iv�e�0 ʉ���Ό75J�	�D/�@{��Y �]�?�/���=yi�ּ{�u�mI[j`�*�"|�Ȣj�f���D�^ۻB�4��̃k�'s��)�[� ��D���n�]�����#H�'ձ��5��R�qd��\�6�i��.''
.�x��,Q3�n�HTE)�iTK��q�!����L> }}ww�Cn+2/3ҋ�M�!���l=�"���M�UK�y�j�++�x-�˵5��Ӿ� >T��PU�&�~~�:$	�����۞됝ֽ�UMT�I$M8h7��`��}���G����#�����~/�n�6 ��]�}[sUR��()�&5]Cy�|$_=�q�ג�s ��I�~$���X�W�-՞T�F�}�z�]�&>O����u�G�`�ݵ�&���n=�L��F�7ݖ���AwS��,���=ʗ=��d;��s�3?R?��w-����\��0fd)��>˿ZI$��6��ˉ�z�����;o������p��y3ђ�u�0����F5�۴�}7eust�=u�,mѫ��l]��i�n��J�T�⢕�{��Gm�;� ��ZƂ�_�}t�"#��ؽ�����&iTS��s~� �`���G{X/��� ����$�~��ѭ�E$(k�Q�q����	
{,���B���J�3�3mŤ g�w�AEn������� �/r������$"��3(Lʔ�A1,���s؉��}˦{ڀA>���kY�{���w�wJ��¦'������󹙁
D��d�-�O���$�9��@6���'U�+�/_�L�Q���@D���U�����(�8�J�U�M{��](��yyt�L36W��a!��Hp�<���:�5}�پ��ַj�ޠ�u㇥�tb���*.6�s2�$LͬyG᷼�sU&bp������N����q� Xy 
"�� A���u.��'�qf�y�n�'��gv�R���"W�6w��(�d��g�Y��n^�R�h)���/]6fA���#-[�_k�w=�������*���^�[SNT��`]^�\�EΩ�qKp����6��b��@n�[�y�>���U��m�y���z���}'>8�[�9wM�A�����b�t͖[4s99�[��.���E���|9�J��ʂ�u���=�wE8�c����kX8�1@��B��<�^cDZ�TO�5fH�~�VY����{���E��Gd�>CnG�����L�`��Λ�g�7XlD�=��f��2(i���:��:*#����N7��G�D;Q��Y�b�&�YDrӒ��S�Y����zE��I�z�'!�n��%^����,thM�ЖUDph�fm���aM���y}s�fN�z���;���q]�{�t����yLٞ�|6�i���q#�~]�2��&�w+禣Tl���w/-�t�un\��ֶ_R/K��+''^sY����7u}4l�40v�:�5�f$2�G��ع��H���U�^�N�v(�o:�}��V!��[�Cؿ3�2�xFʘ�B5���;���;zB�ڊ���V�d�}�qn�8�ry��r�J~��/��1�YQl�A7�10�{�`]]�TV�ɹo#��	�!yQI!kD,J��Q��-kX�Q�Eb��[L%`J�H��Db���TELZ��lEU���ekkb1E"�ADcX���*U�iPZŕm��
����,F)mQ�X`QUŬp��6T��(�J�["�Ո�����TUV1Qj�b"�UV�T�2E�#b�l�EdZ��"��E�+*Ub�T�a
ȕ
"LRɋQ��Z�(��kU��aZ�Pb¥V
���""�j,(��&�UEYb�H*���#+E��mDb#"
��YY*T+X�R.,�LZ�)mE(�EC��@cX�(*1D�
�j��EXŊ
,X���1*�(m�C	�E�I[iUj"����=�����;Pys�>���vW�G�=��5�v޺g���7g��m�ۤ2u��eq���p�I�ɇ�\ڤ�k��9�S�U��hs���/;��ѷ-잮֔��톺@�v���.��4i.qǩ��z���]�quɭ�ٸ����[��d��h��w�G�9��|������.s�=���n�ŵ6���(oTsձi���g4������K�n/]t�n �t��[<�I��M��Yx�vO\Z�V̥�q�m�k��X+��r-9����\�o^�/gs� q��r1�{1�z�nr��m��sҙ��N��4݃VE�1X烟g���ܜ9vf˭[�N��嗲k�1�^y1J��l�\޸�n�Ȩ���Y�+	���[=al���m�6n�Sn�Xc/b�pݺ87N��prsÃ[=��f.�u�p��tWěrZ���ǲǰ����^��v{'J����jr�\�_������Pqp�e�q�nn��k�tk�˲���I�q���gǳT�H�7�����ۉ#��>���7��OF�wjZ��$x3>�;�zθ����f�]�>^����(vݼ����}[q�ԛ �!�=����M�Z5�<�`Wی�6�gj�ц�}�����umn{<:�w.���q%��g�xǷn�т���c�SZ�>�ԙvT��	�F��mlКrj���\;;<roZ񨎖�a�9���R���g�m��n�=�U9�;:v�� ��X����z�u6�b�\ƹ��)- >�n�ۭ��`�a4��-�3[��U�׳�/�ۃ�Sl�n��E���{/��uG]�#kvȥ�Yk��6��s˛�l�+a��fv�V��B�v�m�F.�u\����wm�H�ܫ=io+�i[�!����t��h�mg� vͲ�ƃ��=�Wi�E���EZ���,�g\��K!�۶̚��϶�a��)>z�G�;m�c����u���k�¶�5S�u�[�3�����zS�ݜs�+���S���ݾ�묾�h��pg�]<�rck`9�;���컶�ۺD���0�G�A6�m��`�[9:ݞm�����s�۝��U�7�ں�H�c�k�n���'fչ6��@�*���ً�t'�=�e�Sg����rA|��=*�Ƕ��G�)Wn6�������;���v��0lݧ{����.v��pu��n�o,v���.4���ۭ�.�u]�m��
�����i�znw���*��d;�k���S�	�?��������y��5ߟ���r��`�[��"!��n�2#޺���}C��fuݠ+vw�As�T@�l�����-ߵ؎t��ސW<^&�מ��� wV�!�����Ƭ�O7G�N�nb�I�Ҷng �A4�%�/K���������j*���N
�9{s�$�NCܬ �۳���:Ɋ�T*��T�c����u;:�O�^ǋ�@`ߦ�^�c��7��y��4�$ݯ0�6ڔ����ff*�e���[��;���+�o��D���o u>�,���r@���˻[1B�k��L(Rf(:��ɌQ�ĝ�e�-�նdյuK�;u������骙SSUQǙ��� �3�� ����
�jc�+����XH��m?B�.� ��D̔$SKg�l��&�����n
�t�c8�6�Q�ح�>�MՎA�VP%N+8��倎A���ڳ�bx7��Y�g��b͎�ce�0��������})��[�:�-+��$�NV��gv�Z��s�:��%A2MJ��Rm{-� DO>�� ���]���ĀO�����+�컴�Ӕ���"�iTO��n��7�U� x��~T��&���$�3�o��>neU��� ����s���QB����#;s6�X|��ROmю���}�z2u����'��l ��J���(�y��
�	 7P�z�����1��qF�������O�����m�o8�0�fL��$���y��	n_c� �c��;[��^��� 3��`:��יwc,a"� ���y�L������e��հ��;s�� �ӭ���F����۪�F�V���UP*N=]��+�A�7|� .~�]�$%��:���P�?g�S!g���=���b�w����+z_�]dgo)���n��.���o��Xf���c4ga�o����� �;�.� >=��m*���TL�UJ+�UI�o]C�E�g9dT�ݫ" =��� ;w)�{p�C��o��:�zy�Od��h`������@|ݔ����Md���m���븈�G�{[�� �i��m���5�������'����`4�<�ίЪ��Y�V�.�c���cFv��zW}~�4j(EUT�'�;/����H=��� 	�Eڂ�ns�ZsRU����N�ܲ���*��T�i�AݷM0
&�Q�j��|� @x��O�	�e�ZQ��:���OKݴ��tL�MPD�DTy���΢!��{O� ���n^K��I$�ݭ�$���Y/��Cr�F"fJ�N�����	�r�7�.�� :<���׵� >��nQ�(<2μ<
��͜ҷ2J�j�l�a<��v&�(�
B�Wo#�2UH����t����(,��Jy�d�;m��^��M��[����q��oev�'��f��-�	e��	-��K}�'�d��36_�v�,'�,�D4/�a ����V��Z�U>��}*c���G $ֺ���0'G/�B()&�^�}�����-h�t�?��d>���| o>�Ȁ�ywhˊ;����Zg��E$���d�4��e2UD���n=�A��Ί�ϵr�O�n�� |�{� ��v,v��eX�"�d��^��L�
p�om�L A��� i4z��Q*��S��7v��C�޼��jy6�icCd�4d?���uvcN	���� =�Ȉ�{�.� ��|���8��/I,9�-��8�(�B��&�=˻ �n���Y:/G��y��>��˻ ��j��zr��ö���rY���oN9���)�3EX;L��䯄��P`I�zֽ��/ay�˶/���W8�2�շ�Y�)�j*Q!*�B���e�T�nD༛�jy��Nܴ+�v޲�:��\.���ϯ��9�ܫc���Ɂ�K�c�����S���n9\����v�m��I���&��i�[>a۞8�A�uҖ�q��uq�����g� �C	L��L��-(�\�&ܛ��ۘN�((�<v�ut�0�l�9��Ii+\v��m8���5L�`�[��6�����lct�
�����vkYnw%
yۻf%��Y���dy��l�u
���&T	RT�eH߀I�����9��ٴ�	/?�u�:X�R�m�(È�=ΜD4�f]�ueD�J�(TLT�3�����s��96�S" �N��$��wN��X����ɛnJ�*���(��}�w�� >7}0�<�C��������u��H gf]� >7[T
u�H����3S���m_�ڧ�|}��� ��r�@�t�Lz���m;ۻ�f�515*f�"c���_6� A��M2E���vПV_ n�����kQ n�6ӟ.Y�Vy���8�99�k=RV7��)9���@
��u����^��k���*9f��"U@�oeڰH xv�a� ]�~p§��o|R����˻	�պ�ܰ�"`LIR	�!�U�o�|r���v��f�B��jh���^�/k#rh(�#�f�tcw�{���>]o��7�V�$v��;�BzqC� 䭑�U���=/�Z@@�N떐 �۷M�D(����9��u�f`^Wb�e�#5�3�,����$���绪��I'S��߄� �ݺq�nJ�*���U12��u�W93S�t�"6��:"��7o� _zF�j����w��$v�a�+�j�
DL��z����wc�����w���}�o\�#w�8�a4��6��S6S��H������nɫqY�ƅ9;p��A���uO��w�#�~a�A50T�MTEC��n7@����^�e݄�
�9��6���Q㻝6�X�W�aD��R�Rm�F�?�f�npZ�K[>�$�D��Y�~$���6��M��gT�@�~�{To?JC�~�0&$�ʐɪ�4I'/���@$�Q�;�Ss�QU����:mn<�6�^�^�3QY�g���ö؎n�Ʋ�OgU�T��Q����"�L �luT�F��a}"���mN�-��1�=uG�=��ԳD�ʇ5�'�ق;9�a�+�̻��Q=�R�"�����i]��:&_kʎQ$�6�" +�̻� ��չQꍝY�	��2ܕUT�E*"e��6�Z^H��6��q�ooU�w���:&���d���XU÷�%1���~��ݹ��̥�ct���\�X�<��k>t���R "�aE�o�|�ec�a�$�� ��� :$�\�k�^욯�f� ���8��o^e��.���*;��a4O}ZTr+�hS�[R��H���ix��@�ez�."����-���i/X��bF<�Ȕ$7���n��@|�LD0��i��f�n�om�C�n��u���}}m?�T���QJlۧ�.�Z�V���{��ńGY��h�]<�m���;��`�"# "�bVn�R�����1
�o�1���}�GW��eL��1��Խ�ɼ����4
����)wp��ę�<ۢk= �g0�/ �h��a�ws����^wt�o���#l�mQ�]6���B����N~>L�Nc$�����l���'�Ԫ�m׳�;q;�a���n�ٮ#����ıUԩQ8r5�m����f�� >�ר"d7��ǘ�vW�%>$T|��aP�eUPQ���;����{�"��C�5C}�Ϭ ���r���^�XK��,5O�u�ۊ�0"A������4s;��"35�LDv��d��r=��<7˸�^`	 ��5�D��Λ@j��jT?
�P�6������_���ߝ�|����}�s���GJ��N�ҠW��UPJ*$���l �3c�Z	�6�i�݂d�t;pI-ns��@�W����b�p�Wt��ڼn�{�q��yw��vo:=2�'��]��f)�j�|x''h����Ju���[�a�&\�L�53��!���^���!��\j�l.�<��l�����q��<�ޕ|��s��[{7(]�;��Ş��n̛�I��S�c���󆽵j��ջ\9����ۃ��ɋ�n�nc]sC�3�ӂC�S�_<�r�Ć�n,}?Z��;JV�gq�Cكy�F�vsx|X�;+j9������Vu�Oמ@���ؓn*$u��-f816�X��f��z�/v�`)ώR�;��㵴�����{7=���.����S2f�DOD�J���:�{K��ws������W�ܙy�tWz`�Gw���$Yn��2�2LCO�2���DoV��9h�<[�* �I�$��?6�h�v�O��-k��P�]534ILӆ�u�"��w��E���w4�vp;v[rA$Ӊ��<]y���]�^X������Uq���o(~�Ԁ@�ӭȀ@.�}wafo��v�sU����/��������(�*�B��u��qbIf,�~���LfV��˼I{P��,3�v� H�3[T��J��=s�ٻ�a#�,H!��|�
 �HH2����M�pl�n���v� cm��j��~~��@�jH3�����h �w���@|�o������!���- ܟ�F��j&��EM@!�G��mP��b�zz��ۡ^�G_)�{TwXc�Q��o�Wpv��2�[[�)]�Ď�0�v�6u��T�=�Y���E��|�qó5Kov�����~ ^]�݁�a�ؔW���>����)3����S$�(����ٙ�v�n��A�	w^�T��:6x���O�� ��H�n�A.~��*j$�&&i�GEv��[\�&" y�n8�[�ZȆ;��Vi�[�N.��݁�e{���L��b`�o�u�sp�Ietkq�����i���ݠ���Ԑ ��N� ��sǌ���(�oH���Ok���َ�]҆qm�v�%��{k�j�̿�����g�ێ�T*O��{v� �36w�H��ӭ?%�foK�T9���$�������~�U$J*���"S}7��r��2�q�U{9�{�� �:�� w�i��H4��8f�8�a�u��Ix��p���QT3��M���zĒe}�}�{���H��ǃɯS����(Ȳ�B��sPg���n��-�=9���WN�H�$s���n?\�~6���è��Qy]"+�Wz<R�>�rh՝��0{2Ig��ӈ��2�U��N����w��ӹ���7t��w1M}�Z��w+9��'�xv�-B�����f��.ўA|^{�uaI7gj�e�<#Xv��_68w]���~=�N��b��Oi�"Z�����w\�>ݓ5�\�z�;Ô���{��@���(�gN���b���'x𥏩�ua\V�弐y�t#�3��x�;0�&�|�:�j�x�ܘ��˸�j��b��oV�;��>�8��S�^&��r�^c��Ҭ�Ǣ�Eݚ	���N�����LChR�m8�G��{�����sK6��K�/vdy�o��G�:I��q�\��pwv`�{���M4u�w[��N�4h�i�B�v	C�I(WN��p����/�����w�oN��s?C�v5�ЧU.�"ɞ���棳��ȉ���Ór��������b���L��4��ر��(<�������p�����U�˵[J�c���\>g0f#G9��T���v��N�J� U��ږJ]٭��+6��w"﯒��pC�<}Nz��f��]G��uݕӏ�H�eʛ�V��SXźM����d���'�qU�)^�N6�c���0�@���VƳ�V¹��ͩ��Yn״�6�++�Z��N���$�pc8j�����1��IzEўdJ� �@U@�dD6������"�X��
�-,cH,�" ��lEPX*X�*�2�Qb�QUPcD,*�%H��AqJV��,E�,P��h)"*E��UB*�F�U�DX�	�a�aX*0[n�T*e���aE�ń�VDd�+Eb�R,*)�ZR��PDQ�F

�
�
����
[WEDAAŬ�@�dRA���QF��`1 X�UZ����b��X�����e��#"ɖ��T����$P��X�������V�������pR�1k$��+"�)�E"�L�&U
1HD@TL%���|�@#wv�H" 9���fn^�Co2�����\qF�@�4N���4I-%�oz�a%��λ�z�N��+^I]��%�
�̃
b�$	��p�u�4������^�q�'w��"����p����mI�`������¬� ��m�Dq��5u�y�]���h�:5�vv=X�%�t���x��i�޿�8�d��6�>��o���0��:�� o����.��=�ú��ަ�@�}:ڐX���J��UJ�I����[�Aڼ�WP��Vf{k���m�k�����wh�*����^d����f߲��bQ4MJ�l6ۨ���v�J��V��L�]��j���;�Q q�����%\MUDEMTtѻyLs�vM��Ώv�J�nPH�;���$���BH��ؤ�qaȀ��5�[�R���5usy�p;����o�p⡇�D�(�K�ޭ�J%��2`��)Z��`�OyE���q��USM
*|4{�v����O�H�ځ����f���N��WϮ�� ���z���?�y8��%Y3`�9��:�u��x#�&�t��-��'�E>��M��
C�&�~�5��O��si����ݨ"}z�6ۣ��K� ��6ۢOL���U�9�oc��l �y7مAS�:��� ۭ�$�};�"A$ڽ��i�,g}�T��q��!U*&��y�iXFfmz!�>�[�ݷ]-  �w]��@|ٛM��~uD�
f�jU(`ٶ���f��.��&�
���Z nf�$���J�cw=%�2v�I����ܻ&�WE���f�"�?*��oĀh�a�*Y���/u�VFikm�D�=f�$G��j��ݎ��'Ν�x�Uu+k� ���G8����K��U9Gqu������.��dޜ <xZxƘ�/�RD�V�N�	��~~�?|gb�eO[��c%�>�b�t�:7��\󭵈۞�#�85�h9�.��n��'��M�ܼ
��=WWct���q����Ǌ�)�Z�{Ym�%/m2\v��G��>l]=*V)E���*�����X����<�h9#\3�>�����e�4l���9Wv����.�=���y�m��7c��;;������`8soHmu���40�k��:mt^�K[���m�6�ti�9y{qug�m����!�R�߿����7C:O"��]�a�f�y�� /�Ӝ��D�=�^;���l��#Ӟj�M�b&f!�,�ث��-Sנ���e��~��"Ϳ8��9�@$�ﳣOr���gz)ę1�`9de\�MP�9��` <n��Ds�y7�^Y���`sw�"nu�a �5�Hh�ZLAH@Bd2
�3/"p��s��w���X ��y�� �Ok��O�y�<��)ūX�Q&�{1 �z��D
�m���t >�v�͏K|e���qy��~p�}��� ����N�x�3�n�GT* ����DF�/�)}e��Z�Ѵ�ɜp�'k�F�舕7}��2
���ck�X�%�����������,���)�/3w�;[��D@g�u��u;d��QyXo,a�c��S'�\�w�'�F��E��x��[]�/��k'�՜wZ�[.3ݓY��T�5Ψ�=^+��F�E[��e�e��Y��J �s�ݹwqgDϽ�0��y�6���@��0P�E���9����ܷj�G":�5M�o���y$Af��'{m�N�ɭ�
aS UD�6��[�Z���bs� ���@UD���m� ^盯������C�������R*)����h �:f�r�V�߱��(���"�@�we�� "�r�FG�4�쀩��n�}��/�;V��R�/pkF9�ݷN�qtq�+jc=e:�Y,�[����|��a�c�������� ��wa����Jw�S�\x�?zy� H�/n��{ܤ��M�ƛc��s�33��������9>�}�ݠ�t� Q9�v���س���|���0�4^(�~��m�U�sD�ҋ��ի��d��S0�$7$���>�O��9�dy�,�N����Ķw_c��� ^tM����-p�{��u]�{�=ӻ1���$J�^����v�6Ч�#j"fj@�&iâ}��M\�4X8����$�k{����	���]Oa9䐫�ۻ�K��f�T�����q\��g�w�A;�B�� :�=�ۢI$*$�N���.�Zz�x7(Rᄖ`L�`s�v�ut�t�/T�2��r�2�ɗtX�S���g
���;#��!IPT��*��q�|�٠ �vr(�JC'�"qzD�� �=���.bd���&)@�=��仧��w�a}}˗� �~�]��^]�؄W�0X��;z��o_"P�㉴q�L⒌�������_�R$����^�aK����'���$���Q��]A1DH�*d�r�Vn�CuG{�N�� �.���Awz��׶��߄�&���(C�鉊e�{�z���-I��{����z������Rb��%�V��j�j{�����!fQ6�'Al��%�4;��a* �'�/�X���6Tz󮟬�}�	S�h {��/��TO���ɓus�~�}���/r�~5��ӌU��K@���^\=���t�t��8'�~�?�7E���o��{w)�����i�@������sZ�lFV��Y%����F��X:,��RT���U�2�$t[S�����_��  �=Z��D޽�� �/^^u�n�;�����j�Ha������X�l�VOW��ŅR��i$�mF�$�On]�K�g���Dą*bJ�F��ѬĴ95����l*z#�ozw�C@ef��E��{OVD�u^�q�ƀ�͖ڑղ�L�SJ�J�+�̷�w`��=�k�2�amb����� >�u�` �n]��D�M�УҠ�sY�U=R�j��n��S�9\#�w)��d���
�F�F�?uB0;�Fg���&p��W]r|p�����h���܏��Q����jNq��;:礮�V�t\���d��t���C;v�`�z��V��q\���FvWr[p�)b�5rwL0�Ӱ��kL��n�M'\e�pQ.����G`2�&36^�m�X^*wN�
�65��-9�N�݋�^��tv7Zh��i��nM��`b�fe���upm϶�w]\7/\�o#P�����n��%�[l6�n��D�=A7[81z��1g�=�G��4��y΍�:3�2" LA�<��G?y��2�q������"+��V^]Ǥo6�A Y�w�ڤ
&�
�2Y�ۚ�$N��fm�T��S�$�&�d�ۢ@�٨��,E�O/O�U�]ѯ&%J"J��(��=}�v�=�k� �"w�����������츿�A���� {��`.�`�)IR�TM N"����ʦ��R 7��ŀ�x��" ��ӯ/mnr��u��"��	 �����18�&d)ST:ae^�~H��mt�}q1(óѱ5,�w�ݠ�״�;=��	�{qܫ���9_��� IO	i�	`�1�z4�8��OZ����v1�.۰���{q�\'ϟ���ڴ�j��+���������� t�� u��+�K֒d�$�^}�|I ��{1
$�=9ӡ�� #j�4|m`�=��]�/ѹy�;,'jjB�&�fe�EgҮ�tj��Ցyhx��ZB��ݪ=��U�ݗ�)$�,n�cF��y;$ �'��ڂ$�=7�����P骝�co1 :{�JEQTUCh�nS�h ���L.ۑ�9��wtG ���> �ۦ��B��E0�g1��i�}��J��KP\��׮����� nB�ט`h�,�D�yB���*b%H���I�ٹ��׼-�gdNm?�nߜ4�A�u����dĽ�����$�5���b���K��1�O6]x7c-v�x8�&.�헹4������1$�(����~�o�)� ;z�$�^��˻I�TF><aJ���(�^D'�5V��ś6n��H�"b2�<y2��d��]{ v�z"�#n�$�B�%��o=��?n��]�232���k�� ���vD�WL�f�X4�'4U�U70�w"�i�����k	�V���5��#�����.�%~�<r��8�Ǥ�T59����;�]Y;�����C���2��{ZꔊJ ����m��u���龞8��$�s4"@5=�6�	�>���ӧ�֣==Oi���;$�(�*��G�^ݫ �{^ ���o{����&��Ш�K�'�H|{�i��ܦ��%�����">�!1�m�=��/Y�ەq5�0�+W/i�盶��n�<��W�ޝ��513M W���6D	��7� �����>�q/��� e�]��� ȡA3T�_�3״�����ܽK��u�k)��{�v]{^a l����K����S�~�~A5SSJ��MS����߬ u�y��1��&�����b7�`d�LH�]{4�@���1(�%(�%�k�f����}�n�]I$�e6�$J�u�2�%,�r���b$FF���UI�tRf�J�Ľ4u�Tj�����2��F��m�tK��`�f�P谩�(�N+&�u�s��v��T�RQ RQ�{�)������,�٫�F�
&��W�vD��٦E �t�L�
�M\DR��t�DT/�n����k �zd#v���+����[�ջ����b�
D��=���&��i�	 �v�8绪��
��s��z���  ���l�r�%UD��f��ikw4I�lM-�9�u�ٰ�*���#;]y�����MR���T�A,&IQ""���{-��H�ކ�� 6����C���S��݈�=���D@v�ԏ��MTʪ�����3�onv*�o���܀
������ဃ��ɾ�K�_{��u���l	�/(���$8a��O�DDf_D�f�\WӴ^�����O�z�$�I�;]6�{�v���S��Oo�=��I��y��i�/��E�-�`퓐̚���.퓓z�&�/|�b�4/�� 4�OcX��Z����[9a��WQ��oB��==�����E�Ï=�`�l*�N�]�|�/xe!ƞ�jv<���}u�����t�C!�p��O��Z��#n�:�^7{پ��(�LuIyG.�T \[�D�w<,k�5}b��S�Ŕ�_j��5tM��F�[�nvP��=�B�y,��9�ٜ��g�#p�·�0�^���ǆ�y�oDm��3ˍ��n*=6�UrϙyNطP�楩�u�q8Q�].T}J߰��N�;�T������q�ӣ~��1�k������}��z#!��v�z���r͞�4?����Ì���d��]����J��#㽘p*S9�m����|��+��d	�!S���<)��'�k+ÆS����}��]���$��|������L
�V��s��7vD&=�U=VDM���yת��e��n��%�r�g�`�����y�����P`�O�0﹯�&�2���o��{7�5'����=�����N���d�>�}�\��ug�x3����ݝ{7A�Ӟ!�(N�����ʂv\x�����'������z��yv��BͰ�Ysx�z;M�k�t�v:GAz�*��F����&�쓊��VsiQ���]�{��^=���Clb��PW���=��o7y<�<�>玍�o����5燙ߺ�w�B�w@�)b�`Ċ�-�"�VB�E
0�VPX�U�ͰqH���P���D���@� �
*��c"Ƞ(T
1���a

,�DAV()dX(
V��DS)+�.RQb�XJ��Y

��e���&�*�)�ҁY�QX)�IU	+AL�PQBa�V,P�[ �²�QVT����Y��1b�	+#DPY�DJ��2��)TEұU`�F(��m-*9aX
(.Q�ͪB(

DSŒ��`�*T*1���E�2���!D��1=�>��W&E�)p�1�R���5�v{v��r�]k8,��k9ܞǄ�9�������,Iڬ�[�۪��\*m��:�77b׎':S���]��m�X�ۍqm�5�s����/TH��͎'{u���]�;h�v�]���ɭٮ9��c�X��xꮕ��u����8��kp]�V݉. �sٻ齻\�Oh�K�u���Ո��<�w["�����	Ͷ<%X��xƂo��n}U�[��&��Q�r�m�n`��9�]�x/nǪs�j툷�����sMq8��j�Cٍ8�rݸE9�^��9V˹m�J����U��=�E�cr���K��YyC�cvv�	�@�w/Vm��n��]�0Wcu;�m5f�z�m�5[�9n*(֮����`�}s��.�Z8���h6��  ��Qs��8;pu����ݪ�Ϸl���qV�q�(�8�A8�Ot�����\����U�{.�7�#g{{vӳ��<v��Z�De�l�u�\F�d�8��wb�y�۪���ކ�mm��9N������e7�Ք�V��<�/���[��YNp#���c�l�6���Z�c'>G�2��=z�yw���7 m�g���������۳n��C���+�!Lۧ;��(mخ�)�hGzwcZٰ�� �q�q�X��۬d�.v��v�m��)��3���n�k�X8�6�.!8w'`G���0;ɺ��ݼ�=:��r�'�j{�7d�뀞<&�v�ͭ����,���[�qBgqg<��[����ʷ2��9:������:fؼKëۛ��Jm�G�z�l�W����e��֭���+�.#Qіh�ΐ�v�c����V'��|��=[=�o+�3\��s�.�i3�y��n/+�[V�{�����8On��z�u"��fk�ɘ����{����{�����5uջqu�v�h�c�s�O`�v㪸�;2�<0�v�ulMnQ�f;qɒ�ܗ�X<�E7F�H8ڷԽ��V㮞�ĵ�Ml^r����r�&�T��^q\P���UӋ�7cgC�Z7��V,����ڲ�-�;����u�fz���K�xPp��9.5ѱ�1��tv�ݫnïcc���%_`�JN�*�������H8ݗ{q��|��c5��m�#Pٻ7u��|I�/R�y[�����Nz��<����.�.a����(*��8������m�
r�H�Y�۱�$A8GZ�LSU�$���sM�������MH UIF��=�q �� z>��wo�\=����Y�xΓ$ ��Λ��OnA2D�IJ�M���ۋAZz�!.vo8�}��@E���Mz>��@�]�W�1�d_P���J��&	�@�s�i�;oq����N������w� ޺o���{�vy�R Ȋ����C�Nm׊��z̙Y���v�ס�L�|ۢ@'����u����$�ݎ!��l�A5"���%U:gn�]�`��}�3U�(����1���p������������<�k����@���n�k�������K��/�n�q;����ԐDJTыv3��*��AV��u6D�w�Ղ�������q�c��#���� e���;�"��LG���$�g����<�tc���=��7�����5��)y�MOn�-e�<��9�O�������貧�z9o�(tÈi�6�O1�n���檔VO�$�z9 �-۾�� :�)�����0$��fy�ojU�@M�sR�S����+����  ��W����̎@$����"unSh���ԓSH*&f�'[�S=�-߽k���<��>n/�	mvy�H"�n����H�J!ǒ�ywhk���P�bj�P��*�)�� ���j�yU^��*�� �m�ݠ�$evS #�n�D_�Q�r���4���V�5<З{Iu���l*s��p����s�6��ƾE#��=�s��h��Kn?�g~��ܬ:�+� �ݺ�D;�t�k�*}U�ku�]� ���lN�f�U0H�NA��M��MIz�W���5�[��i�Hl�P�H�׭�����X)wKl��:*B�	��)T��H7����$��.��X�\Tô�:���i{k��Q�rʧ�T�Q�� y�<����N����tg=�&�)�:�7ßO��]�v'�Ȏ�ڍ꽮 NG\׈ ��|ƅ�h�
S�J��M�>W|8d��V2Lg9�AS~�H +Ѿ]�:�7k���[Y��6�m��$�`�پ�@?����ə��B,�DK�^$�mu0I#��6F��c:�J!�ǈ*bd���"  �9wH<�0�T���W(+����Fw������{r|;t�RehV�x�|w:��	=�yL���;wso�{>�>�M�T؎л̺��)����ѿx�v��e��_� �w����	�x�$�c�m�[�2�p}���J	)��PB�>��|I���~$v.8Bu�qK:F�o2��'ǳo ��֊��Ø[X��^jOK)?(��$��~gĀH�x�'Ğ����
S��4�U
[�Z�]ˉvۺ�F��=Z`͙�O]�CF)��s�r�G4�;ms�eG>�Y���6,M9UR���《�h����v{y�	#7B���*�m�x�I�{"��Ç���u��m�I���`�A�{4����ߎ�o��
�+�F�w9�O':��ٲ�n���X��8�:	��������]�l5���:�͟{u�0	$�=�"�u��t��m��OwV6O��D,@��Rd�o�2�ij��hD963�籒OoVS$��i�N�l-��JAM�-�
A�>����~$����ę:��}(���/6��$��8�CC��2J�30�%��9ύ���b�$���A�9�(��ۜ�+�צ�sX~���`��Ff���Yt y���G_s�y,�����@P���^~�o� ���;�B#J�
�n'�,�{�x^M����:uAzǜ�D�y�X������wsݭ����\�(�w�\9N8����ʺ�B�#��	�d[�؛�9{<�{�{���k�V<M^�����뜓�)8%X��nf��Ϯ�wn�j�A�]�g	�%�պf+�p��8�J��v�9sU�c�9v�q*�=P��x9�uλSy��'���7Wb�g9�j����J�U���8�����G����jɹSVӸ:����6ݦo/oD��9�Oiɺ8������oO=mg9�n-J��u��c�vd���]���v��-]����4ؼ�I
Sd�߄��`d�yĂ}��m�MK�,���Z��>���B{t��,��&�`���������s��E�V�O�NTe�$��� �k�ۣ1�*g�{A<�"
�2D�lŹB�
�� [�4�\�V��@ ?L�@�>��餭�@��-�H6���]�^�:���.�H�޶�'�^V�x;�x12Ar�U{D�3&J(���z絲��.�݀�zH&v3��t��k��{�u ��v;YƄ���:�+��]9݂��s����z-�(���h&������Ø[X��������v��|Of�l�7X;�"�i��1e�D��z���V_$����0T6%�c`��*a14A�P��J�g�܍Яb�]l�#�QZ��1�U��<��{X`��Ҟ��*���0=����-��srov�zF��s�A=z�* �;b���G�Fh{
]b��+�@��8�I_�wM'��ޖi$�F=��nCZՐGf�l	�X�8� ��(��LŹF ��#dg_���F��6H#�e�1����R��@K��n��SÍ��e��7��}( ��eЃ�{&okN#`�1NߟwV6�1�����������P��� a=���m�s�[۞�=�{{I�L�83��5*:�c;8L�f%"��7s�Oă��(2@$OFZ�MZ5��s��x�'������˭��Eff&���d���0ގ�{�Y��>���s��g�]@&��d\��"5���e�H�J�3E9}��@��Պ��H�˜2��i��j��ޗ���]Yg�lXs����~6�3��^bty��=J��7A=�GH9�w1�\������n�y&f%U��s��?	 �,��|\ʒd���̨�OS�.6����v�I=�A�	��u����d�Vʞ�Ѿ�ym�H��s�'�Ė�rU�A��͇�MϷE�t�S0	�m�I3��z�!�kaي��눞��� �W!L�Fb�w��\/'O$uw%:��v6��;����v��z��:53"dɑ�v��d�|gS�/{]3348DI��}S;�o��d�f���µ�%(����e�Ӝ�'e�oqQ��q��7ē;P�O��kd	������X�|�d�2�]�I��(G,v ��s:���"UI���SN�����$�'� H{խ�pU��PIS`�lz_f;2�ɲ��!�!^9+:��Iw���>'ݝZ�t,K\�Ut[�4Nɚ�^)�gq�v0�סVfL��*{R��5�I�"�ذ[b��uY9,���t`�z�H� �T&"��.�1?qc����=�&q���Q���n��n�Oc�����^�$�ݭl�{:���`�Է�����9�ɯ1�X�<u��^ݝ��Z����m��&�]�f"��`���1%�����}��̂I�gV���+89aM�	���`���L#e0�X1��[�)�_��u��t\������I����#]����f!Md1UzI�&QQi���������dZ�)�5��K�l�	�gV��:b�e)�RJ&L����p��>MVj'ǫ�$�Ffֶ	$�<ψ���h�EȒ��h �GS����R�Z�y۷r�T�?S�f�k`��x�֍O+Z���f_��o�f�{���v��em�v�����D�>L�Hٜ�h��<��q�^��Z�����䵕x���ǅ)���=����%,%�I�x�fݹ���{��w��؀��"\�!�U�pZx[C�n���|��x�m&W�i���$���[�.x��Sq��]�^��.�rmn�!��N͎Ǌ�c���vS\]���uĚ����棴pѽ�=�KH6��C��;hfd�gY�ɫ�����P\u��s�x9N�K�U'�.ú��-��-\͋�9�����]c�wQ�"�E$�2�Cٵպ�v�ݝ���������,��3*G��l�N���$�L�<A�
*��Vp��WY��I���~�8��sя�S;�ם��&�AI6X�z~?���h ��oĂL�yB��r�7,�:m��d~�0cA�7�>����I�O*	&����B[�9���H����g��@�5�J*D�
 �`���T��^�8A ���~'ĀH�o"�.���|�sȔ{@g{�*�2٘ND)	%&M=�@I#3�[p{]����A�#��	�'�T��Kޭl�>?��rt5�&a�`�I�	6Z($��u3&c!�ť�knc��c4��O]�Gu/������BlVe��I�Y"	$�V�c~3��N���q�I ���&���̣3
bf'�<݆J�T;��l��Z�	~�i��%?�bet�
Wn����Z��ٻ$�x�;�ii{;�=�q�i<k7��H��2X�Nܑ�[����+EK�l��t��Ujh\��{Ex�)�*M3�o�I�}�͟��j��ل�n��A��*A��{ZiL�} ��UT�*��j��k�{���.���ܮ�H'��Y���| �~,��>|��X���4��?0@9�[L�ؑf;S����:�z(�Hv��@$έo��L��:LD�g������Kuv�ݣ<=T^K�^��и��ɺ�y�����-���~P\:�չ�u|$����[ �;:��Q��;7{�����Ϩ<� P�T��l	}����*�brr��~$�������{��Y��^0#X��2fbbf$P9[v�$ݭ�	���U�Ib�1�%~GLNHl�}*5�0EO���JZCwtŻ��龙�N�5�'��VX�]���#*�ߧ;���9�R��$w����1��gq5�^���Cq�+�IQ�(�Z㝺�kN����f�+���j���mݎ��9��z�����i����rK��k
ۘ�]Fh�+�+��u��L����\8��!6��3z	�ۼ������r[X���t͵l.Ad0P����F]��H������4���{Ŗ���#}�{�rMЛ�E��%U�>�]�7F*W��ҭ�j���(h���.G�v����C%��j^a��on�E݁5���욞ݜ~L����nT���w=����Zt�i揃��ƫ�-iR���3�pԇA���L�◦<Z�����;��G�Ic7.��{��Ѐ�Z�yJ�U�>���<]�i��8�f2X��}���6a�p��E������i�⺲��r�AABo���`�6�K7�3>}*�t���Ͱ�:Z��KΣva���3�"={������N��~��7�p~��+O�@��@��ݮ�+���RdО�:��\b*�u��<~�h|�����|�A�*]�+�ʳ]�t��2���X&\%�V\��R^�oJ�m�����q�C9���GZ�m�}�t[��oQ�U��6���c�vv�S((f�].L.�WOon��/|���C�{ץ���9f_EnI�ڨ�ܯO{��l�c�A���vm�4�u�zj�+z�����
8@0���@��#E��ĊE�H���S�*�\��"�X��4�IQb����`�����ˊL(�b�KZE!PRP�l+E� ,X)�AT���QA`�,UAjF(E"ʁD����	TfZ���B�f���Jȡ�%2*�L*)
��+�aX�CV��ŕЬ��T�0U�

EX
��UH*+!��DdR,`�BV�+YY*
AL0�,E8HVE��&�RV�)H�Y�*)�T�<O������p$��[ �mk~$g^�@Y|s���іiʊ�����a�O����`Բ�88屗}u}��U��=h��L�QU PU^u^�O�=K.��2!v��P�<�#.�d�ͭl�z�]z9lY"{�\A��"v���h3�Ɂ����cq�-�qp�p��1�Bs�x���F6�c�����s"ޝ�_�7����I���`�H'�Q��
�m�Hڙr���fְ��8�bT�"D��@�O*�
�݃;[K!Ŏ.1�d	��V�	���P	�;)E�w�.���z��2�^�d� �r�1�A>8kn�$�[���0�sǾ$}����Yt&�����l��M1����޿��.�E��g�'����$�O*ہ@����ܲ_O-z��t�̒��VR��k/�h^/oR����M�c��t�
x��(i��ݧ_E�`��5��Vq�ò&�v�L��sv���$	�VyO�R[vW��|o��rn/J���1V|H]��5�^�/y�`�8��`���}�,�uZa{�z�[<mw�.��D^y����1s��ߟ�?�e�ԁ=��l�A�Yt$����8����ԢM��Ѡi�����P�X�	H�f�s�>:\ƈ�-�����O��Yq@�K�z� �S;S+K;��Ξq�� �#��'��E��ۤ�z�z%=�n���0��	���H�/8�x������ǚ�Z��uú�\��BH$��|�$�}��:ZX�u�@�/���=�Ǝ&[m,lCW��>$�EZ��T`����A9���M�ֶ
0��Әs�Ic[�8�L{s�Ļ�N������O�ݳ�m38��z������{k�+c�W��i�2�iX25u�8�p�9S�u����=�;3�f��3�P���ݮՅI7\��]���ѳ�l��3ŭ��۬b+�/�slۖ6�����Y�W:����{�q��l���m�����X6�r����W�:��mm���s��^^Rn���6�pV�*�LŹ������Yʝ�yrnwC�]��5'q�:��kG���/&@-�FMaAې�` ��I���3���r��G)sh5o
hs�,�5o_cL��)�%LR��f���ߞ2c狶������{(I$����$}���*(�Z��W'�n@�H��͂b+*
1$ʐ���tK�(.�����ڞ-9�  ��$���m�|nzqp�̸L��vL	R�D�5Ӝ�d�y��2AޡB�D T)W� �/y�d��/�[`:l�<H���l�`?�ﺜsŮ��ޏ��'��[�I��t� ��qX�y��@��u����D��B�RS��N{gp���ev4F^k`�N��lH<m�0`q�F�P<0���/}V�g{�Wn6�h��G����㎳$�[�����n��>��	�b&B�������gĞݭ��'��@2�Y*��ݍ�I����~P�Y� �0F�rH0mX�2R��7~��>�l>Pc�pNC�E��,�"�cg���	�%�a��b8r]��Oo�t�ni"�쾊y��A'��h0H<[�Ab��.cN�"+*
*ș�����wM�dŽ��&1,ێ0&�+j����ݭl	<[ȡ:70��0�ٮ����X��)'ǣ/�0 bo��>}կw��+7����XB�wۤ�O�QcH���l���ѐH9�Z�j*�d�f�4�՝��|@a.�� R�o%CO�I�;x^|�i
m����;�!�,��,��֭Ϸc�m�gںK������D�H0����7�$�f`�����a�p���$�Z��Vڞ�W4L]W6 �i������@`h�RlblO�_��"ge�D�`�.絇�i�P ��Z�$������t�}�6��p��:��!b>� ��$c{*i��
�;�\�j�e~�׋��,�$q��k��{7�J��X�����%��x���f�<{%��K)��C�DT�+mP6������=�D��ZÈƨAQ*DL����l=�O�؊�kĚ8���w���O�f���Ҧ�&�i���s�O���T�
T D�;�� �um0��Et��v��z(NvV�� vn����Taw��@)B����̅.��;�C��ixr��l��$B:z}Јw<O�������)�3'�t���s6��I�u�J���8+`���7�]O��l��a	�Z'5O�e�mܛo��-?|�$E�W0�#�u�I)�M�@�{0܎�h)&&`�����ݻ�C|	�q�"L���٨`NgW6H�u���V �Ig�A" 7���d�h�h^��r���o7]2<[ƂY8;�Gp�:�U�Ed�F��Jج�Rqm���=[�1�1`bdl�r�ˌ>�w^2Pxc`�n��ҹ��TG�e�6LFҡD�2T�S47�q�I��ô�s�h��]�	�M�lE��lA'�ڥ��3�!�\"�m�y����a>�l�ӷ��q��2�l�e��ыu��Y�߽��~������p�&�u��4�K�u�;0E�B_^�	'�u��,TT�� )�3&�x��zH2��9t�K��2�*�l�H��m�	�O(H$TOWjJ��*�.������D��J���a�@8i�I$�5�s{Դ��zI>����x��2Ԕ�A30L�:[0WFC�J�C�H���`�I���{�����SX�Ń�]��;1BK=2���A&�UUC�wU�@@6��~Y}t'�����Ӷ;���liZ��5QU8V�ԝw"*(�yv{��uc��Ox셆a�}�@�߫��W���k���?����wn1]+�a�W�;� �K�R�NƱ�Fu�i긞�8gV��y�wn����֜vmkxwcm�zU�h��x�g��v����%kF������x�"�n�M���M۞[%��qZ�>H6�.�.Ӊ꺳����{a��D�#�<a��+��f��sA�=�r�쫻]6��۶;m���6��]r�k=�y!hƌv�8����D8�{n��nN;̼�e׃�!?����4�<W��������I^�zA���l|�\e�d-yl?���Im�L�JA1-���a��W���\�vu�>'؞�
$_v�d���ј�6f]�κ��**A
b&32�Q��W��s�m���-jl���1�����`����АI��߉��dJEDD��Jq�����dTif"a��UP��|o{���;wm��_r�C"w��}(%��I3%��@*f13�誶I=��O�D�S�r�SP(�}�m�I#�v�7"75m��_��ܙ�h���N�h���Q��vvv�kb����jQm�ZT����]�?�����=���$y�l3�|H��مBo�	���x�?����N*�b)&Rl�L�>�{��G�[�U��dЮkG>��ȗ͠X���ܯd����~���⃮�t�ޱ�W���<���V�sU��:[�R���b	�̜z�)������@U^�� �x���������pp��DȄ�Dߌ�v�^v�2A
�ͥ���a>���$���o��1QR*bQ&T����qz8f�$��ӕ�2	$��oĒx�_\Gu��+Q�盭�}׽�0e"�ġ(��]z�'������A�w$_f���'s� �i�j�1�e�����f;�v�.�ۄ��S��n���(�RLrR�$����AB�bgE�p*"S0�����Kl2	��ݺOTe�!�q���ݨ���7;n��z���K ɐ��[��%OL��q]\�1��|H�ݶ� ���@@&��1H����HDB���.}}����L�$��$��,n��0ĺ
���*�P����ckEu����,L#3I~7,oc�fi�&Y}�ԨU�ʺ6��s���>�{{n�ԞT��^�fD% �#�����Ż�ă�-� �A=P�Q$����l���&{R�i�wo0�* �� ��n^����w�+;]ڳ	YV�d��#�ݮ�F�h�����>�m� |��7E��gs�󘪗���kȭ��f=�8rR�;t��#�������:85GN��4�Xd���Q�ݭ�
=9t�l\��'ǥ=�Hq�J��T�@�ϱuU�⭮�uO������z���H��m��V�tD�x�D��Mp;�؂Y&L�@�c�$_o6�����d!l�]OI'�e>�@>����B'(b��4EMQ���s�웓�w13�bA �W��Gnkl�Ofm�.K��ڣ�0�v������ie�+�Չ�}D��7M�ɹݯ��!3���o���kL����T��x���ܵ3=|�;�S7\�=b�����~�"#��8�2�K~3���`��g]0B'{��JwB�0Iqڨ	yͲA?��hX��SÛ���C�,<,�%�Ji�ܽ��&Ȇ��Y���v�ݵ�5ɺ��>��?~wǈ*b`�*`:�|���������~���/�{�^@�n��H����(*�S1j��[��ǳ���3{���u�����C|v�#���q4��TA�"Z&��zN�i'�ۛt$��f2��l���d�w{[���h�?�9Ye�Ct���������^�I9��L�:\e�+��MH��l��A���%J��b��1�	��q�˫�̅Qܫ��"#P'�7�<���>�x��	!I� IO��$�	'� IJ��$��IO�H@��B���$ I?���$��$�	'��IO�H@�|��$�IM�$�	'��$ I?�	!I�`IO�H@�xB��$ I8��$���e5��·�(5�!�?���}����
���cJ
hP@
�M� �N �"�  Q@�	 )�}P        _  -�>��wwl�;x��5��^��ў;�{�M;���Sw�ֹ^;{�s6ӻ�k&��6Yg�7v�[�  =(��}�=�;��;9�.me�m��}4��:{�x>�Pn8>�͙�x��YR�У�   ��6��[kqwm����qr��K��{���.퍱�k7\�4���  !y/ڶ�9ݣl����h�P䷼�kx��[[ݛ6֭�^�   {��k{v;;��{޻h��wim��\�Zǀ3ʤ�;��w=o1�Muwq�x���nu�Wv�s�    OF��R�  �L� �`�~M2%*�@     5Oƨ�R�       ���J$�(�      ������      �$$dbLE6�&OQ����SmI��������[n�AD
\�ŒǢ*"q��Ѝ��D)��������Y�O�G��6� 1�8D@�@��J���l��FA/E�QUCP;=5U������;�ۤDD
�ו�K5���Tu{r�MBO���=c��Z�,b�lަ���g�j3-Ԡ�3YY2em��+�e]��Ki��/6��P�V�vf��!��%R�0��&ں����!�<�/i�jl��Ÿ�_t�M:�f�/�tAZ�Ϡ�feP�v�6O��^eҡW*�Q�.i��b���S+8,U%X�k�M�!AV��[s��A1��Ж�x	[{��hk� ���YCj�ɹ��T��Z�sC�J�H�Ix�b���7Le�mMu�q�7��C�U��Huk *eIx�Z��4��)sq�R���&��]-Z$��6Ycq9i6\2�ӭ�(5x�L�a��3���n�&\Yt�̺�6�WI�b��/p�	*:�̘���̄�R(�n�hPwr���a���ںm�IE,Ib��.�S�.�;���:zv�DBy��y�f7�4�Hf��?\7Pk�mф�ו���u�P�e���5OyS90���eˋ3��BK���2�Z��u�f	2��!դ�FY�n8�3�2�;Ya���U
�f`�����nc���´$ [�ܷ��H�n�d��3*�Sv��t�*TFI1��ZS�t�̰ʍ��Z�i׶25�c� `��LeFrٳs�����Rj�4f�v��Ss�k(�<�{ח�jQSl�4]���qDȪ.�^X����Sb��g/-�4����Ofȭj�3��sMk��{���(����E7����V��+�/i`���,�t�w�5I�gUz̭P:cV��㧇U����ʌ�"��-�ň\3N��بAgm���%,+q8ݚ�T{ U�#�姘 $�/^�t&�M9ue:;��!r�c>-�v���M�.�,JεW����AoCme��9y��M�y-��
�Rܒ�Q�D5.ô�J�i:8*�GE⠤�m<��f�_ӰāGh��u2�(�,�=0�p�'F��i��܆:٨]2�V�Ò��KJ��9.�J$*ۗ���kN��Z���Ҷ�F�Vb�����DD5r��*β��dL��a�wV�ІR0��hc8�3GwQ�[$�lRU��f�Z��]�cf,�m����64�r)���÷n<�v��d�×e��Y{�i��*m (Ī��u��Ѩwbe�>w(\�EZ��,�i���^��nM6̽���`|�
�s%�Й�7fl��f��^$�c"����T�S��!"I��c$U�����#۲�L��I�Nr�(�,��V��ܗPm�U�����J޽
-��35=X�۔ɩ� �Th�R�����l,�;�Ǖ1�c��0]�d2��Me���v}�r�GIqOwm^�iV���R�$�@�a �QW����.{�M����wӃ�S��c��yҭM��J�{�4�
=�˱
�3���ݣ3,�o{f�UpQ)Y��6�ʀ��U��Bnh���
��ǆ��eS}-��1��u�wX��MXn�#�1襊���K��ih��D]�k=7C�W/�t�Q�%軸��Vt
w�k�)���6�����Ƶ/tV+լٽIcTM����dl�
R��z����B<Xbwen�l�p�D���V�ők-��)�O]L*��Z@Y6d`�[Z�䤠r^�6�5cRJ�aP҅���nˠ.�bZEkFPDc�BCy(V��-bQ�:��j��y�ȯ,�������Rm��wv'kuDei�S%�/6CO:�]�������fV�E�)d�v�$Cm��̶���)�����
�8��	��w�>6�T�GV���GtX�E7��Z�a���iZ�#
��T�" (i�n���l[��wPFL��l*(#>0([u��Pi�C���vd�ɳ���֊�\�KI��	Ex��aS�l(�7���)y��^^�"GV�{�l�4tRX�uY�x�T]���@�r(�*׊k*���orL�Z�l���&��J�����Z�K�E���.�ڰ-1�)E����p}#�S�chd�
:I���/Tu�,`.t,�=�I @AdO�F��TU��,� Ȁ@��	 "�Z�����$�(H ** ���H�"*Z���H �(� �2
-ER������{�:s�]�㮫?x"��[�-{x`E�JDRh���
"���׮�]����y~���n��������B��u�8�d�:�����>�v��}4XD̘�`' �?+{}�s��/K̳t3tݓB��Fe�/��'5vbI���Z�=�%Nmf��5lW.�U幤]�2X�7s_]�GO2��u�r�2���U�k�)ԙ�u�\���m�j��כBX�=4�h�5nf�DL�h���\;oeKW��9�KWc�6D�L3��z��Y@��Q��p��Tr�9��Wm,����^�.�g4wX���\��#�4��Յ�}��:<B���ˇnk�Wo1Ib!�X�E�t��".��R�;�B�o$�+Jt^�e(��ڢU���%����v�7Ov�Ԙ@�s�*�:M��;S�qSn�=j>@
�i���w23�`�[ϯ)F��ٿ��][ǀ�Vt}�WVn)˭������:M���̬֖�	�Ȕd���id�x=�ܧ���7�:�]k��4�ym|�6wr��76��W��j��,��fpO&[�;7.���b��f��4�Vy]8ܶ�lϟ;]{���{�3��]ȎE�RR������T��E�{Üy�w��d�+��9׹��U�𙁐8��,��9"���[y`K)3�\����6���mW�a�]�Z���K��2��S�.�`KF>������;���;.�2�Y��)LtS���R�q1m����㪟V��сR&�]�x�u��8��w;C��J�^v�_w:R����Q��C�&��C^#�QZ�h=ג�Dr'��	��5���*nU����3,J�X�/;Z�`��b���˃���v�d��iU]V�҆H��q}�A08�U^���>I\������ފ���+y�<p�Үwb�L�u����&қ��Aj9N��
wyD+XX۱:��ʋo5�}�4V@���ڽ�k`-�uH��H�}yg�����X��ݧ��+�7>��a)�>N��*p��mgF+�Z�]L��E�)	�̄�7#��h�9�bͶNȩj�o=z�hˆ�䏕�X��P��u�:S�9H�Woh�إ)�Pb�+ΡS+,��K����Ӕ%i�JC���t"�x�udT<�IL\e�麭��;J���%٘K�ɧ��g)���Ź�>��T��ٱH5�y�������eX�tfF��:��`*�b�K���o{�����ۺ����z�ܗ(n��`Q�ȶs%�Yάko6^����7�ӥ��� ����I�ˬt��Ծjk]oZ=�ᓖ����ohx��"��J���ƪe����y�e�\5w�mp=+lާn��K%t��WGV��2��F�:����R�]�o� 5�C��"�4��6�F�d�jrL:	c�J8��r��c��w�+�S�/�بܛ�ڹa��d�&ȉcV��[C�ն+������B�U�&�kF��w�M���s��a=`n ��y���ntO��\]no�.	1,�Q��\���ֻ��NqĚJ���e��8!ht�V�8cl��U�v�q��ń�ͩ�t��jFK����� .�0��onS��,�4g\`��*���#�7W������ǔ�o]fRAa˱Qөj,"􇅘ز:�B���J���ڱٮ��3R�ʻ���z�̜h�{|�LV-}Vvv<Ӕ�Y�cn�;0�"�m�����v)\-b\�3HT!L�fm�\9�X_M����N(8��T��*u��;�Zգwi(3c=��f��mw_n���J���صʳ�Ch|�#@�d��m^�5���R����_r�զ��W��LjV�^RÓgp�o�����e��]��Ӧo}���m8-`7GEչ�le��,�e��쭵}��/q:�����}H�*[ ���[j1��Ŏ�"��Z7A�7��>��5EM�M�]Rf�5����Ⱥi�l�Ȣ&��f�K�5��Y�L*�.+�sK�+��Sց����+'���il��:+ц�J&��c{[F3W��^[���" @��'ކ�]�5T����~*
�y�*�+X���M�v�0�Y�5��* ��6Q$%UZ�S��E��v���[��!�N�M4F�7i>�P@�Ey��u�����]�jF���^����Q/f�ZN�7�W9�e��f�Ť;A㇭�5�=��۫t`��.]��aP����y�瞻t'+h�yv�v�NC<�C��œt7cF���݇�n���uWl�k�	�锶�{@c������kY��Z�ɦk���z�������n���{m�9��͸к(�ڝZp콮��=��:\�z�Rk[]����2mΓ��P!�5�Z�Ukm�v�E�j�H�n:���D�V��c.9� pi�x|p*ӎ��us�CJ��7]��1  �wc���fs�mւ�<I��Ӹ_v��U�V���۱�GI��.�[I�G��7N�����&y�Γn��aBtx�[�זm�sEU� !t�%�e�V�{E×�V��uq�v-�:�Յ=���]�o9�1�����<V�[V�ǭ�g��dD.��`n,Ş�ks�ܻ��]d!7lF�lv�v�ۧ�����n�e�[6�t������ӹ���.��Ig�@����iiɀ{,�ϵ�cj��V�;:�+7eu[�g^�;�;��k�E��͓���-�X���{N�dn���y�9Yw����\��\l�u���#r��a�n������:�uM���k���wN�n^��^�޸�6�.�lt=lѧ��ڵ�e��{G<��:.����6��5#�n��c��������7a�*�g��-�nz�=v5�,ub#�R/<n@u��l/g�b�C�U;<�1v�'�Ol�8��<='#[�
8ݞ�:�����=bG�ul���n�sض.�{l[m�H75m�h��o[]s�t;�4eP:�I�;g\��u�������`mDv����j�Մv����n5\bG<��q�Y�狄6c�m[�ˇ\��Ds����[h�v�n�гYcs:
�6�[q����;ag8���m=�7��+�'<�Pt���ۈ˱�D.����*�km�]4]v�+������K\v;I�oܧKA����n�c��\p,l�֗��Y���)e`�&��fm.�)�:�; s������/8�[Z{c��9�۵�V�4�n���*d;[l݇��s�:ݲ99Ȏ���^C��δ����Cu�t����iָ�jU��g�[͵�N�:�$L�tJ6Z� �,�<ltX0r��'�.�%̐�1���v炎�u\8��^�X0sA�<^�ccD����P��M�6-m������[�͹6�8��݁8�i�>�=X�
c��Z�BB�ڠ��uی=��v��C��ʕ��݌hǷV��uk�4ݹ6;pY-ҙ�g���A�Y
 =�����&��	�1�pB H� m1� ��Ă�$H�C���H@�4�d2.� I�Ā_*�D �p�s��ϸ�}��)�c�W�<q�DG*q�O!r�<� yx���<<I��!>e��t=�����S�G�=ܨw+T�O=u �<�����\_�ֻ�T[)�P�pu֣
�.�K7%��.��A��c]λ
�ۋ3R��<֡�p�+���m��� u۳[�~/�ad�k1�3Гu�<��:Wb\S�'Qu��&�ǣqx��sv⮱]����V9���t�7+��n���v����dw���t�ۮ���ѭ�}[=9wNx�ݶ�����y���[�-���-�՘��#�mz���M��t%�R�:���&���5�tp��!��;p�����Sn���֌ص��a�]�w/m�3�y|�3�h�+�a=�w[</n�����:瑈k��e�.���8���R����d�a���:�oAO%ת�_c?�=?�����m�,u=j}W螲���i��7�(0``����&W�e���U_�z�c Wy�6���^X�x���:EG�:�p�ve�f�0U֟$m6����Yu'�K�J�J'lw�<{�7��}�[X�/בTt��K�*7�^�?Wګ\l��'Pܧ������Fd�s直v��:����}�I�Ϫ�9�s�}��knT�C��dx���i#�6��K)��ʴ��m��3�{QM�E��B� T�{u��A�'%L|1���\�dwL�_e�j=���f��J��^Ϲ9�H^���A��zw�uP�{]�U�T�]xw҃���D��)�>��i��	�dʟ};N��
M��d��B�3N=�����H�T`��6J�fJe4~����ͻ�TI�
�>.*�2����#/1�T������	�>=aش�2�t�v�T�R�e�Hń2�oX깠�S[�Zkt��%�R�B!����^����3Zb�r��,���w����!;h�mYEd�|��"��������X��G�6X��;�͎��#�V�b�e���'Z�|�c�.^{Ϫ�o ���7����>�Jh�C1��uǋ UǙ�rr"�B�t�K�^�Ҏ�����!dպ�j�ͧV�j�<�ɚۮ�����r$Վݺ�`�����e6�V����I�q�HP*�nZ�#��[��ކ��b홂��ꩦ�s�')�0�}&0��͙�˕�;�ĪC"���gׂ�/�i�9�r���ԚY�^ߟVa$p�>�A��N��a>{]�c��F*Yj�s���e�q�V.��n�#=z��p)�߽�{�n�\X�Z\X��--h���e�VyGJ���]�S��i�"��mE[�T���5w���Q�l@$����)�R��zfu��@n�*���S�L�Pr��k~ɇq:�\q�éв�����JD��'}CN 4L[�I/qR;����b��/�(�ސU��Ѱhrf�<��������Px~���[�cݾ�k�?1ZZ�]Z�z�v":��ѕ�	aiH�t=̞�7��}|q�%�?��>�:���s�
�f���]�ܺ�_&��\n�q�e�����
G�<SӉ�o\d� ��$�k\��ܔJ�}���#aK�l-�7�~���hׇ�*L��T�]-Z8��S��_ɲ�nYI�RK)a��d�׉��&�4�Z��D��<�V�g�/�%؏�i ��3�=��q�^0G���eE
тy>���+sYJ�F"�{5�������K��͐�`СA���x���YWѨ�YK�I�#���r�����u���v�c���ۈ;kM���-s�����j�n{n�V�猄���}�2�X���<P�1�(�Qtb(�im;�zy@g����(�W1�2^�dJ��=X��* �1]��\�}]�x��H�?9���H�f��s���L]n,��x��WW�MJ7\5R+������^TЊV��rn��;汷�s X���0 ��S~��h�[��:���s����oT�e��'�=�RH��S����~�U����n�b�읤 9�7T�5�a�՞&5��=�O��5}�g�Ԃ�sa��ϩ�-�� E#�*Jf���S}q4[Ys�V���k��z�Ƃ5�*��R��h�(���Ӕ��qBR�|G�By���X5
5J��+�C��*�5��y}�pr���Փeʛ{�XH���L�ˮ}I���ҲG��DX��C
�g�}8LD�uw�w���KT7�&L�Ӝ���L���R:�]͚�끕�m��I6kC����Ns�۟0�\L2�e;�F��[M��94�A�ͽ����ˠ�l@X+�AP�;
|�ڪ\����i
����f�hoCٜ���� �6I�D���q!�C������3�����{�������PZ���܇�ϞyNܜ�:y�x��Nz}p�<�I � $ @6��܀D��>��zy��'qLx��6D��&"  KN8B!�Rڔ	$�\/�J�|G����%Xkc��>����t��a�ݸ��Z|Zu�ֳ^�3��߻�I� �X�N��;<{`�[U:�0X'��mT���Y<F�E���l�~�2�9���"�9��,�$�g)��tŚ�3�E���������v�g�[��)��:�;,��&��w�ծ�v��7�fPP�[Z�ߓM
��V�Zgs֯<m��ϯ���^e�N_�ϫ0�[�E|F�D,��E����R�;�4�td���1�Q�S&�aȐK0C770D\I���k����&V�4|�F-�]�aoj)�ɼ��P�"C�r����_G��'��FŹ�٬L��6�d��vM��6��ڻJ�[�ݸ3�7�L�F'Í�p�AEeb�H���QX%	'��U�.��}�W(�hO�D7sa4h^����������.��H�1a�E��MW�-4b�>���;��ƕg�x��h�i��Ll���Ѥh�ן{��{��D�D����VI{�����>FC��+9>���]��*�Y!5]u.�k"c� ����O��}�=�qH$}B��"}��^
���y㺯	��8�u�!n�占���7U6W8����oC�b�j�ص��S5�+�ҖR��s0�q�g�E��@�#�i@�7��k�UM]�۞�5k�dB���K��a�s8:�!a�q/B����G��?U� ���W�G�� �_<�M���8��`�8}}�Wi�P|i�nr���"��Z6'H�TC.��x.&c�hЬ�|ԣa��g�8����zb�z�&�仼i�NSZ-��C�{%ZV/��k���w���C����:��ʪ��G��Uhb[7����>?}�6A ����z�
�~���rj#����T�~��(��X����N��y�*zu)�S��v�!z��۾���2��"=�I�ɠ0�e����kF,4N,OzVk_V{����dvE�f���h��3O�lh���b�h&Ѽ�deگ�խ5*�{�������Q�Q�
��Ѷ�	ʴv�r���sε��m-��'N��Z�vw9��cWi�S��;k �5�M�E�YL����!�1��d�Z�g�mA�=����V������sփ�ͭJD�{q�_�eЃu�4M��z��\�qZ��fM�Cﶬ���N��qJ(�]5kE�m��ѻ�s�DI-�Q0#����Joj����d��з"����B��]1�N���61ˀ���|T����9���3�#�#�L�Ntf\�|y��$A��3��1�۶F�Yq)�VUc��Df0�)�g���;fh��ʏM���m�����
��A�6
���Yܹf?I��;>�n��l����I�_S�:x*8h�Ƥ��x�,���D'O��{G���^R�"����9�3�9=�<=�F�~"̉�����?ALE��i�4��~�ک�+Z��m�k���5�f�����Y�РW��(K��?˕,��[q�6���^n�9]�H���¨|�Ն(��J��ߙ�k�|,#�M�#1�
�~ͪW�$��[����R3�H��tL�[WQT��oY��C����[�a���V�-��v�\?\?FPo�� �?x՟�t���e;���&zT�뉷�����ۡ�?z�V?=����&��H���ǖ^�����j�B���oђ*d	�o"U�����	-H����t���(mH��BF�CR$����@�����?h;	�,�=R�ц�7�pj�{�o(-*�__�/w�'���;��.6����5�2��0}���!����>9��-4���3�꺗�l�k�c2���XwhԺ�,;�n�bx��w��!7��x�bгOb��y��앂A!�:["��͊�٨9�O&D֓0�hF�v�E�J򽣱v�a:��s5�y$ȵj�y�T��;]�b���Ū�����,D}� p &ppKOS��)�' "��
�� B�1��#B@�H<���=\p��XC��AD�OB��:< �u�9�y*H��B���BM$,p��Ԝ�G*±�J�zy8.8�y*��� G������'�C���e��~k�ӳ��49v�7\ӡ�Ʒ��v�nF�ЂRj�Y��L�x�Kn�<��r��lr]8Ȍ����1���ڵ�7�vM�[��d�\X���c�Wn�R�4�Z��u�gƮv��F�Ƿo2vzg{v��۰�Y\�v7$)*a���M՗��`�ƭp�^۴�!$:�K�3�綎���퉷K���r�;g��ݐ9kƮ+�dq�D5;v/It�݆���Nv���v3َ;��'n�ղ�&��*�U��Wh�"6 ���ݓ��b�v^�#>l��� wz{V8��e���{��+�opq�*�@+]R���l!(h�o�]9ݹ��GT�;p[v���9?!�|��b��Z�����#�l���lB@ɔ�����h������h���B��q)��,�^D����1���Ϊs�$�ɐO4��I$;����:�<�� /m̑ğ]�C�D�@ùJ�窩�r*�"ޭ~F���vX�rЦo3��5jk��H��^�����j�#4���<\�ܞ��h��ؘ����Ԋ�q�z<��g3Y�C��6S�%�VF}wkb���>9 �mV����8�ڔp��>�e�i�O��_O����֟�P�l�S�'J��JEF
��"�{=)�}տlQ���L�͚����v+pU��fO�(׶4�E�q�V$�v ^�c�U�ko"٣��	,&��+&~� <5��'��ZR%���8$<� ��未F����_Mڟ�-,V�s(ANE���UlVP�4J+$��1����j�_��[i��zwu�Z�|I�g��0���`�����x�d��Ц�I�cx�W�:����t{v����g8�)7�R�A�{&Gz,�S��_�[A&_W�_�5lK��oS�^���k�U�)%�,(�-%�����{j#�fk뙳u�[��2Z�iu���"M� �up��{�5M�y�rx�$�<����F�H�g`IGّL�-]���ճ��Wu�i���Cv�]�ܿt�ZfS�4�E@�f��w�_/�}��U,#������3��9*�K��η���P�\�K�Q�'���]֦V���Qۮ��`�y�ꉊѻkþ����2��$m����hX�}�:��J~��/�@�>&Y���
��l}+��`h�}o4��G��	��.�/{�KR���\�����턒B�[(IS�5�}�e�4}��T��=��nFʏj؊<l����������H8/�=� �J7>4���]�?F�oo߃���muD�g�n�5��ͮ��\�;�s�s+��Wz2�F"V���o%醳�lm6GxlYb�f˯6�<*s#��R�͙Y�˺s�'P���Zȱ�ЗV23�{�V|3�;�1a��-�&���%�ja���1����yȉ%�
&VR�|��S�����>O����{Br�)2�Z�`��ჸ��5�=�ᴥ���{M��z�W�X73|M�\�qU�O~���Ͻ���ٗ��ʶ"��ʈ��(��s�_�.����e�^�]w͈�ȟ(���-K�VP��9�fv�"�:BiB�=��<g0H��=�R�Wj��K�_#:���+��f�tЭ٨χ��z�!)rܸ7<�� ;���EUqb�ڇ�M��;&���[b8ěkn��Eύ���ӓl&k���6�%�í�����/��ׅ㼼۴.s��� �R �R�����W�������k�L���jx��_[�@�ԋ@���xg�6� � ���燇WH�H�@u�!���9��k�M��D[�E���y��I�l%� +"hQ�O��6J���J�t�*�k�y���NbߚxE$q�"L�+���� ������/�G�c�zo�@\������q-�*�z��9��ӎ9 S�6��W0�zP�}_ڹ&R������7�8��o�:g�f#��P5�@����k�k�b��t]��Hoŀ��� �@�wƯ| o�Wx����o�Q/�"Q��@�z ��ڸ�R�/{��JӖ�u���?ߏ�$�K��}��6� �^"H� q\s��5�ж�q�5�00DMb�-�z�D����j�Z�I\��� �(5$C}P6�H'���ӌ�ڱ9�|*���գ:f32� vns��`E+����Πq��'�}kQ�͔0�(�ޗGX<'i��J�����Y�2=����HY��6�-Z�<�/{�q�2�����ȓ�=Օ�iN��r0NhΓgX/��_S�����X۪�F�ά2��!1���O5mI9�k3v��^����X�KM�]�`4j[��R���uNoWE7�ü��7��U�3_cɿG{ P�7$1H�<	�sr���w'��Je8���y���U�=��;�|�� ���'��؊磎=���3��n|�\��Z�y|z�L���"����\{/��c����|��rZI-Rʱk,%HU�R�芆y��!��h�5Ch$�����P7��v��q�F�\P�"�����3j\�M��*����D�P�	��qtJ��T�zE��ؐ��!{�� nZ���~I,�K����o���Y�H�9�M�f��2� _T9�kW��
���M�R�Hm�*��TRA8���g�h+�@�s�7�-� �w���6D�G8�Es���8���
ڃX���H�ڢ�I�MDJ :�!���j�uRq��x������X��-��b��Pyڇ��󩽰�� ޑ��YҮ��@5�[����يё�*:*'X����ޔ�kм�D<R&��\�8�[�� k:�k�j�1�!�)R��%E$m�6��Vhs��W��m�يH�W�}`L�L@(�:�-�'6۝�| [zk�Ͳ&�hE$�Җ���@T�\�
���m|��6ڐm�T�H��� :�2 Ih������%�&�5ْ?����������p�j���,#q-�۶��[�hytz�7f�eL[m�9�i�ܰV���v��ۜA��#%V-D�U�^�_m��qnP8��"�F�c�_{���H$���ؾs�Z�@��.��7�x��%����4�&7�.�f)��q��f���D��@�) ���| �)��$]zԯL�'��ws�.�<�����Z^3���]b�ZXB�R[��g��ְ%��y�T��w�y�z���Wt��3�)���� ,��:�>���V5G�h�ٰ���$�=��ioV�`�7���w�qw{���=s�A߭�v����#ރ��o�����,�S��u��u焼�V�\E��"�{�����Q�ٯ���xk����U�J��s�� jyQ�6�����z��ͣçv�̫��I![+�$�7��ĚɅa��ךO������j��#��k*��+I��HԿhw��W7�ZxC���[�O."h�i]	軼��������S��Jٻ�y(���+Bt[EH�� �JT&R��|���fG��蝎+Q&���a�=�e����"��R�U�ª'o|�'���֊�tW��r����3<̗:�t�c��N	|���� ���)	��S�A��F��g��ĕ��\�é�W]uͺg*�1�n�%ն�B�vs���s���"�k+i�������)��-�pTk���n��d����`�^(b\m��r����K��5���<�졃�ԓ�^�5���p�����Q�DE �VU��{G�۪ꖚ��~/�.y\�Z0ۃ�!�oB9w-��Y���~_/�_������|����l�J��ʃ|B��j�5�wN����G��r�ra�����N�b���*8Q�[�e���Y���GW0�{+����{�YP;�ٔ����av�?gVQ�r��,��EC���<=�]��{��_SQ�F�]a4'���>�v�t�+g{v1�6��L%!D$
�$��������c̖l����勼�uj���{�+��PI㙷j��-5��W ��A���L��]�8�:����R��vn�
FVa�Խ˱v5#H�HP��:�o??a���jC�g/7��o�:�����啒��my��m�l�_���U�?.,�4ٻ�K�
tw�#�dB�������Y��#n�踍�tPB�teoB�i'-�ѫݚ��Sq��w^q�3�,J¤��l��݀��mf�8�dɣ@y�b�qd9�E����9XZ�)�v��rd���7[b��
��]mE�F���5t�9�5G7��m���6�m�WN��NR���ZL���v��{�m�\{�[���uyXo�Ʀ2T�k�*5�)�V� ƻn������s{�����r��$�!�#��N���s����ɫ���/�'������|;�秮/s�q�U�*���PG^8G�sǃ��^x�p�y���n����z8��,���[��+�<��ϗ��l�'��x,��fZ8��ηn������h��k׹�|�~��jKg8��*ö��L�0,��Ӟ;	���r�V�1j�l���H3�ij��;X]�H;Is�q�.-��	�tf7Bn��;/;.�ӛ���E�;��\�l��l�d����;�7�t��y�Rpn�v����~����vI��wn+`��n��2\s��;v��|`!�n˷fS�6����rk�3�
0g:�m���T��u[��N��3;t�s�v�ۮ�1mo����:z�	�[M:4��9�9�m�Z,g��g1�B�Rwo]h֥C�Q�������������gqm3cq���\�ݷvz]:���g�S����1��K�F�{v�����YW�9ۆ�-��(���jQ�����?Zǯ\V=��Fx8�<7Vg�o$a�H�V�[�%��-�{r(�Ճ+ox��>kt1@��O}q�% ��RT!ѻ@7�g�9�^��dު��~^S����6mww^��w�T�� G|��;�*a�Ggb5����>��,��4�4+�du��]`[�G�������ޫ#�JI�3|�������6��eچL�$�Ix{׍)jn_�V9u�I<�^��}��ﺸ/eV}����v�f�Q�Χ6=-�S�v���G^����LWeٝ/�XD�p�#,�.���Ngw��ձ��&��w����^�f�U�b �����$�:zj�������uO��	;7C+�eeE�z�0�iZr��w�U��LtA��b�$3Թ�,q(��j����7�~�r��]�z��˜��#X������#[�&ܷ5(�讋�*��c��lU��k��wZ�U+��D_j�K�Y%؉�u���]B���ﵦ�:�P��B�Jܲ������8���ݭq�s�-��9��͊�ʌ�iO$�n)+Nս��K�M�%�A9�����GV�Տ3;^��a���Z>�B�[-ࡾi�tϠ˒��Tx*��(\��ɜ��ۙ����{������R']o'�g�m�C?S��*FV�P���$ƃ �p�E��z�f���}�^p��yW�}�z:R�~��\��n�C��㨍�{�5ADjZ��b���@MBYa[L@������}o����ٓ]Y,��sF>���Д���@��N�^���9fE�Ӡ���q�̍���������l�!���G߶��ܖ�h<>���R�F��;am��^r���;oǼ��:�}�X�_�[Y,��m��es�q�V%���+SU�s]��ݩ�`㌦)eT��~�;��Qa�'��=��ȉ5�W�!Ec������q}'SnTW���QAܻ��q-�E�Ң7z*���ꫜ��<i�@Kʜ�X����̗6.Q;վ=����O~��9�7vIiS���R������'Y6׮�^��ը�q�lb�_o�n�'��q��]�z^��� ;E�m���Q�UX�~��������ˆ�Ⱦ��� ��xr!%~>��<�$��y��k*YCUr}��+�A�A���:������k�L~��e�W?o�Xu��s�9��)8�[T���n�˯�?��-6��]��v�_ٕA-ޛ�.w����au,�7/8��M��J�����u4T춊)PW)C3��z\�<v��-�g^�4s�@�jۍ=���Y��mWS�bYE ������ւ��M�)S�]�7����x���v忓߭dՏk
��ֵ�k2�.˷� Uu]��t�s�u��2�@}�:��؋�&hKO2Y�6H�v������]2��r����j�u���sy���ۢ���:(Q�!�䌢�)=���A]������������v��l�%pAO9��oH�KE�s��,[|���H�.���Q��Sn�^D������y�^��WG9b_\�>��Ѷ���yXxT��w�|����^N��{��>��x��g��7�c� �Ǟ�wG)σ�9G�]����Q�=��8<c���_��S��<<��r����j�U�O�ԣ�OT:��n���[VUk���yҌ�~��~j�3$UE�OZ��*TGI�V�9�̗x�⭜��㚴�M+"��z�5W��5wť�U�g!�_9�#30�/9T��c%�X�)�w�_���M��T;�T}�a4�~a��Lq�@UeZV�(є9�=�Ë��[�
�ʎʉl&�W6�i�(Hfڥ!����>w���Z��=�:����,|Ž]�̵�%y_oM@���G���%��5����u����X*���#UW��B���n�Okpm:��o\�s�nM���u`a���X*��p�d,�/�߳�'?��CU Q����b�]�5�u���v��B��k%���¨�9�H��=��\|��֣�_�-u�1NҸ�>�]$a�4؄�	�
��Q�7T/Gt1z6�)Y��`��uk�&�����2�߱�`Ҽ�OjB!����o*��}���q�]#��{�#��2�6��H�F찌N�c�5����f�ݽ1*Og9U'K$�L���r��^���;�N�L[�})�]�P�ű5Uo�{�y}@gǞ�,Qٟn�e��_B�ہfO7Q]�1���T�F�Y7A �*T����Tw��U�x�F��[��x):�e�%��A��S��GXd����H�^�Y�W��H�)+u��FA�χ������}T_<��kP��͘�E	m�m�v�3�ܗ����	]k �Ƒ��a���r�Wutʐ����*��|p�G����Z�������uY����w)¤�c	�^ޙ�xp���|�;�,ꂔ����s%Y�޻	�g�݃��{i��;t7i�w��m���n5�����W@hȡ6iYv����X[}�fC�_u�Fuط��3ykؾvX�YG�yť�
�5�{�Ŕj�\Y�y��}��p�q-���{�[�7b��T+�u�v볺WOC(�w�WT,�o1�3rNt�LH�L�A��| w�g��*�G�f���m�kc�5[f��\�����"v[�'�Ga��j`$��Q3$����(��k6	�r��Ԛ�yl
�S�
��~�v��]פr3���.��d���z8���~�g�a�@�s�u�U�!~�Y�P���5��=O� ����v�롼]��Wә�Yy�\�|�,�(}H��B�p|�|m���=7
��U��U<D�b�GR�N�.6�o`�Ͱ��w�|�ֹ�=��.�o���e�QJ�d����������Ͷ���w&���i�Kg�{R9��;�u�ސ�;�;��郮�wB��,�U�s<��P����8_O��5o<�o�]�V���nƑ��{c;2�tZ`-�vK=gOmd���1�a��5Ú/meVVVH\+Y\`�pj;�q��9F)�n�U	������b�2����U�lNM���Lvd�5�k[�F�
���S�:�ss:��k�fJ]�c�#��s;��]ڗ�X&��y ��W�fV��Gu���=W�r�������q�Zf�o�}���曦��@�h�xu��*���/)��xQ��������'z��Wpq� ッ��y���Tx�O(>N�Pw9�Ǟ�<qO�̼!ѧ�0��Or9��P���T�s��;��������Ӓֵ�1��Ԧ:�{A���wѸ�m^a����˷<d{V��j�����e�]z9�,\rv�v�`����lS�mr��!z������h[��)ی�O9�5r�$�h�nf�����1��n.�9����q���N/�+:ܮ0p����tZ9{;�S������ݫ���j�yv�6��Mu�ϩ����Lnk�ݖ�u6��QtX,g���\R���B�,좦g�0��93<g[��B"��X8+X���H@�� �KT	P|�j�,��@��=���DN�u�����G��8�63�Q�����M�1���ٮ�(��h���[��웢ɷv��F�R�䖂�Dq���`�C�����a�;�t,��U��]BP1+�Y$N0�Ō>��ۉ\��Rl��^��sP��%����[�w� �b��@��VV]����t���92�ow�"2�T��GE*�V]ǌn}�[��~=x�����W�U�p�#0�5��Բ��F���0��7j�j³e���g�Gԉ���?Z�4��%I]���:���׺p��ǲc��)�BUHZGG����xv4�Xm�c����2����w����.�����ж�蘊'j	J��ԣ���R�]�|g�!FX�S$'�R�"�+Q����]��w�}v(���>A��$�w��g_u�¬�~���x��p��t����Q�K,#-5噄�ϼ�Z�36t���*��d����n<�6iVwEO�r5�˛�k�^�z��Y����ũ�����T�x\6Yfg�ؙ�e��ݴ�k�s�����;��]�%���:�S�;3�&�[Z��7@�i@+�����)(�:2��lv���a�t�-P4�wW�G�8���^/giڔP�YSG�wd���O�( Z�`�系],�T�*�r+F��I�T���S�ݧ��g��Uk"ܴ(*��d�����Uٕ���p��n�jMT˘�[O4ϝ�ǉE�N
��T� �{m�+'�\�����l�Y�����X[y����KԥmOZ�ZT�~�R]==X�� �p��Jrgkf����_o���Q�_������� L5v`˜fK(���eX��bZ���^����w�P��V���=�H�UP�31d�im�����(�^ȸ��I� ���xȳ�z�d2��y办clmX�s��J��D���e�B�)��}�?�x���d��J���Q�$IR�y�Q޲К��eA��S���O��6�ʷM�twE�g��JU��,]\+��/q,WM�����u�SMVL0_�dx�R�[���uc��r̀��(:sTmNSc�n�7f�:��㮱�]�v\n����ϒ�Q���N
�ID5`�bu�r���]��'�{ը��H���6ȣ\�������2r�U�@/�Ҭ�e��{~�K���2��
��i];-��UK%-3y=��=؈T�w��X�e{���V�K<2�9��{�j�!w=+}Z �$��sR9���m����k.:;{lV]���ˡ;�T|�뎥���6��N�ʕ�`� �����K��� �#��V�-��.<ȼ��3G6���%���jƺ�mD�hhe�]�����6/u��ѝ�J�W�tN^��1Z��-�,]T�R5��v@]kW8vJ̮K2�Ñg�o\�ɺn֩Yi9tn���X�tD����B��7�t�P�s2�_?�U̾��¦�����on�"����=F�w��imtj��FM��˕Cu��rd�.a��ރƷy�����������T���#�c�7P
"q��z9TI����M DK&4	���6�"! �-�64�Г �;�p�}��^|��ܢyP�0�u�tuW'�:��$��@q ���Jkw����ԍ'PL?g�r��-e\���"�v+�G<�b)H V�YYu�c�1��)EtwZV��eس"��s��ќ�M��5��m�6;1D���n��l�e�WMc�xe{vC�Ҽ�6�vv׫L�k�p;hj/f]圸�$��R� ��;��Rs:�(Ş�����%��s�;�`*I<SN^�[,�B�카}��^��;�A�� Q��ϳ,Ö�)�<r�i��c\��Mnz��k>��E+c�����GM��y,vh�]l��h�6�ۻܻ�mŌu�iӄMd���7g�ѻcWKn���*%���V���_�0�{%����ʻ���f����NI��Au=D�nD�V,s1x��̓/G'���!�Du�6&Zok3�V���
!N��J-uT.Y�S�}�&u��ѻ'n�[h���)U.�U
�iN˚ͳ�[f_z%�*�a�T�Q�]u���UGF"���{y;��|���q���"���\5�rTx^D�AW�s��d,��̩w�0ǥs�����e�9�����$YL	���F�Oi�����ӌ�Z6�r�*8{��Ky����o\S[�iJ|�c��ډޝQ�Y�dc�4��ͬp^��.���)��8�.l�S[�9ouP5]'2u�����Zn�7;� 27-:T	�����<���3����6�hf{����k0\Y<�Օ�~�*@�m׼="2��$�u��\/^�A���V㪰�3�wT����6��쳽|�W4���ƃs��n�ít���������Xٞ76�Z���[�!�^�ns��fw6T��aÂ��;u�N�B��eF�(�JaH;�ie����f�dEФ2w�T�2,����j�M�,����H�hʹծRF�kf ������Ue5�ˆ(����'#۹��nUL_Wp��u�ζ��6��P6'��E�;��v����U=֖7!�F�x�����g"۔��6i5j`�H$��-����0�}���{�^�;Y���T�Z��{0C��IݬuS�'���J�G��s�O5%A�|��=�)S�
5�¯�җ:����)վ�DT�
"�[)i�d�3:�-�������0'<�GX|{A��p[�l�]�*�&�+��R՝2U,��~�̼���y̡��a���S���T8�*�����NS���`���p;���j�{&������U�����z��)b���DR��&j�F�t�;HP��֏:�72;�"�J��$V%�b26�:T�f�m6�d�^�W9k�b�FjG�.�b���.��V�;f��L:��W�J�0n�-&)�����l�yup+ᱰa3*�7)�l�zP��s0!���n^������1�:���է��zh���IIZ�&b"Y��tyx�.`��Z�M^�`7��X��u%������+b^�%w��l:�\�x�Z0+xh	/Bn7)E�M���t�6��(�`�e�t]H�yWOn���@6�A�����z$�N�C��8 �6Τ�M�hB&�4����r�"��܀��1`�8��J<������ �O t�<O '<���x�O<�r�''�� ���8��_�ۦv�pcrY���9޽:�����m�[���^����d�����{Wk=]��v��um�y^�,nU��gu�7c��ێ��^Lng���]�0:r�e�yQN�2t\;cY��8m;��!]���t>;�-��\�͢\��`�<�jƹ��.\;�;�q�c.��� hf�(��v�-�I�x�ywmTG)vQ�Kֹ"��N�<�ûs����a������֍�$, Ž[l#p�pv�T��h����]����)Y4���ڎ��h�v xc<'E�8����e]�e:�;�]��ƻ;nv�sM�ѣ����=R���M�%��s]Y��Ƙ;G&θ�wY\���lt�����R�J���{��H}�wM�~m)���Yw�(H��
^a�{�D��W���:v��BW=�SQ_;4�f��D�V�b�}�*3�E�v�(��:��[y����Y��Z)&�)g$8����S�`�	μSEX�SùV>}<R�b��PRCދhԸ��d-�,�������DGYD�<��>g{b�N��{����Ing�mt�*F�P��2�.�z�Y�L��Ҥ/��d��ϢĪ߉�NS[碲}1�ָދ��wUQ�Ш��lQuϴ��ּ����ܴ���6&Zg�=�m'n8D߭�Ҿ�\�o�����AH�A6<'�r�>���+�@4b�W��ԯӄ�j�Vp�wi8kR`�43{�
����V�.^c\��$R~����D
����\��4�#hi�ȍ[�'�j����Q�*��X�,��=�ŮH��t�� �e9ԭ�ͫʚqk[@hМ�ݿ3��:�p�_e�Q��V���;��sh0hB3뛤1�/u_	ut�O�Uvp��4.����W��N�����v�=�;��tY�6�k��M��O��n&)��tc)Ӟ��r5˻\�V�7m�q\�;k�ն�䲽<�d4��mA�)[�Kh���y��/d�q��]�\qd$Tz8Y[��,�0
�L�ln��(�z�>�;3�^��)���3w�zV�SQ+�f|��qfH=r�H����TJ�����W/5��@ۖ�%(尖�8�q���"Ɖ��u�6��S�9Mp�s=wݑF�S(A���MT�3$��8��L�8b϶UOnk[��!{�&,�S&����eL=qZذ&����ޓwk�A��ru5%	��qݛ-�dB�\���!Þ��.3'��+r]Kw�K��O�h�����L�����K��4�H�A������1��<�1�%��/  ��#u�KY]r)�4G8f[R�����`N�ϳϫm���M�������%LRZ���%J�{�>(�}j=��,��u��jl���һ�7]z��j�d�$��י�	ndb�Rh�#�Y�2��	6j��N��ػF6�f�xv�L��nױ�_��06���p��S|q�p�yc��TS�E�:�]n;P�>����q� 7l��I�H��0J�7�@�ճR�^�Y��x�ى���M^s��zZ_6'��@,��)�S�Ip�C� �Ҥ1�`�Zi�. ϐn|<s�<�!{��OY�x:���%�)��-��N2�e�ݲ��lR��9����嗬���,���n�/~��mt��m��lD��_gs%6�Oɭ���B �̂M���}�$�L}a��v �`��Z%�Q�smP� �":-P&�y�٩�V���`�K3�j��R�7Y�5�-cU�ZF�lB+fe=�<CJ��@�
9M�e�^h$L�����H{��sY���3ѣ�OM���v��q<K6��A�*�w���iOZE*ʆpw3�w9P�E'=a��	ہ&�ٙ	Sc�OMJ����'k{Ұ�/����ѽyҶ�R� ���%�s���^lA�q6�kξ�V	O5�wRq�;���ȰA'�Q�i���V5d�E�z�vM®ӵvM�5�����Ru"ֲ�r�r����k���"R�T���M�v/5C9�;<�m�5�X�/�Y���UXw�zmY�K��;�'�"9�V�SM���Z��K�-v�pō��old�LB�����&αWzy3fIGQ)aV��"�{��u.'GO��'4�W�#�� ��x33�]�.�lt/�1�e�O&����j��a� ����x��i��4����Pd�*��m8@@shBi� � Cl@�����![B^��A98y<*�w�8�G�O�9S�(�<��0!ˆ�p�$B!�p$	�\���_ �+��<��PA�!��D)0;�/�T<'��� w���P</ 's���x�r� @��i�<3�m ��Ϸc>�1�a�Wl[���u^��φw��i�����A���a}dp*�C k��W���MD��z}��1�nm�|HZ7�] 0Q�!�^{��қ�$a�IDA6{8=cIȂ4��y�����>o�7��	wu�5��WIyd��;�Ǉ�tED׆<{�a,��B�\�0L�Jorq�]R�4��D��,�W#k�4�u^���~�tԩ��z~���A�3�ЛC�g�W��҈3$��J2ez��"�8�5�0�Ȍ�ۚ��3[��a� n0[?-�^R4f���1l��4A9�Y��͋J�H�|I�5�G\�۝S�������b&���ǫ0��k���3Ż49^7h�J(�ܴ���6&Zsܞ�V�S�(���Uw�[u/V��3��R/��1}>��Rj*禧
�"��2*��m9 ��p�Μ�grux������]7;+՝RY�P��7����w�hז��I���Ecd������'�Ъ�1�Q�n���N��l���,�2��j�:
��6��q��ZE٫��Z���L]�m�Am�ޝ��+u�R��rҫ���l{=5z%����T�#I^��/������6���+\�߳�k�"��+Ҭ�ج^�=�j��k�J+ZqcU�����'�x��R�l=2!o]���b�vܙ��B�!�]�t2�����s=��W�U.��b>ɐ4�J,F�njT�D�i?^R��U���..�g��&�I@r�K{�{ίH��1 �Bׅ �&C��,��N���F�H6��q)@Wk�X��X��NH�q���ܤ�~����ڹ�@V�m�ڴ�hn9���ʻ/كͬ=Z�%�+���"H��u]�� �cܾ+~���	��]'��V�AR��4����zjT�׍m�]���ۋ(޾u��lS'��#��&�̖Nd�}Y�"�$��kjE�<k�g����=>4>��=)���U�@��j�"�>��r��"FV�L=�]:��1@a��~��:.��!���b�[�nb�X�`z݃��a%j�]��dnX���r���<[�CC�\6渮��i��)
�m��Q��:��S�4K��%z��ꜚ�+\>���hKLY�H�IG޻uy�.�@L����!��˭IF�k�@Y�$��G`�M};M�\���5M�� �Ư���PH ��)��{��)#��{�sf�$����cUf`@y�ٱ��MW���>tc<���X!�*C��4=�٩S��N�vU7eLh���OGH/Er��C�
�Uu��b�`2��U�2�4�:�S˲�a$�1DJYm-5�̔�<ԭm���j͔�Ƙx�ϩR~�砎83V�M8�覨F�!�$E��v6f����}�p���*f<|#�d���kw�* �D�K{�2�Ⳬƍ
�w9���>,�v}��k9�b�Dq�D�K)�s�V���`�
���>����T5`��L��d���zͥ*]<�AN���h����{���V'�:��v�B�y}.s~�xMb�Y���J�m������T�L����̎������~nFޓ|V	�� TF���:�y��ȬAb�.ܣ���vi�i�V�B-����3}�֛r�8Kޞ���I�k_<�V��z�m���]�NO�uZb�8h��J���$�jT�����Ȓ�T�$�I>)T���iG�䈈���R��9oG�e��Lj�5��E�>�w>�1��@�_��j�@Ƌ���U
	x@���!��=#|uYZ���P""��'H���һ��^y�Ӑ�m��߭[!�wܖ;�6�;]5�3��f�ٱ���`�hR�x0�o��?zq��_��ϼ��E���  �FD���9��D���� ��낏������z|:�4	G��o��~�}^����F�`Lx� e�h����d	7O��Z_�{�W��B8��= |{}$v�W���y�g��dDD	�'/������!,`Qg�(Ue7f$�M�4X�uV�խ����wN�C���DD@�����>����/������d�u}�9��]����o��Ə����k������#H�����L����:��������K��C�=�g��)�?w��<<�����&�p�}�^��u[��~^ω�tv`��o�3n���d?���g�$?�(�)�#�CԨ(��Y�DD@���6���yQR���}�Ń��h�P'&�d��@�d봒��6'e����iDQpP���;�!���r�p�6�P���4!�������U&�1��X(?iqDD����=��ܝ����3���'[��|O��z�����pw���jX���/L�O\ X������>\ȟj}��-��t4����DDQ���흨2|R��|��6I�D@���3�f͏��O��o'�>.�:=���Ä�Dr-���ҋ��-��y�A��|���Ϙ��~��>߳�Xӿ�c���`��w���������M�{�C�w��T;��^��Š�&���H"���X/�a؃�>o��u����D@���;B�2�]\a�iv"ս,���2�D$��J˞������w$S�	v��