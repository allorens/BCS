BZh91AY&SY��q�eߔpy����߰����  a��1��  
            ��J�J
)P@ E$R������RJBN��"��(*��JJ�@f� *���ps�akrݵۛ������wnӸ�ݍ�x�ɷ�� {���/^��<i�z�R4��t��f��֌���ꞷ�%)(�j*��CF��  � o��8�=���R�z<IU�=��Z����ґ^��xc�"�1=�+�VƮ��%%{������:5[7����@�  +�g=]�׳z˶��s�E-������w=^y/=�wG�xJ1�l못ރ�"��m��v�{���^̻k�]��&	�RD 0�sƽ�OmͪVκ�oz�s��t������#�ʷY�У�wv˶��<N���nJ6ڪ�z=6�b�n�v�(W  �E��Z]k������{ԥ{�k�F��s�={ɯW7M�A�������v�z/z]��TE幯wJ�����k���<cG�                      �  ���J��#�`�F����#@��L��
R�&�2d�@CA��E)&R� 2h      i*�6�mL2L �2F
���D�OA2�0'��D1�m)�zj���J444ɚM��12d?�?���ml��Q-*?�(`�ip�.�R���,2�u'_HBBrR��ffٹ�f1��fٽl�����.8p����clپc�6qϗ�������������������D5�����6i���7>8q�Wyo�Fͳf��\l�-�&sʪ���9�8���ǅ��ݷ̗���nw�o�J��$�S�B��g�x��,���(��&�V�a#$O�0v�`���a# q0�#f�Bu`���?�瞹מ|��s�2�����kpɹ�"�!�3�-�(,fs�`��+܄�iX�q��!�H���h�Į�:�~���\Z����1�L�'�	�z��gS����c�����X�|FA.�Y$K�"��k�̈́�Q
�%&j�T`�aXǓ�<�X2�¶�c"2!2��e�&i�!q�!��0��eC"r�3	�FI���1�ň҅�!��0��m�!&sf��Id1)��f2E.�9��0�PL���j
���\IEj�q&Đ�8q���p�ap�e�,��ED�б$�a2nT-b=���<Z1��b�N�-I1/�1�Bdn�d�>�I�L���8c0�%�dC��X�Be�}�X�0��f1Α��kp��:�J�)�.@���d�UBc��3�]�&2;�)(�[���2c(c݄�����ZH�N�@�|ϘƢ$�(J38�8��}
�1�N4�u������P1�.�󈡌�L�S�c+Y>�h�B�d� �E�0V`�x�f�N�;�>�`?�6-)�
�C)��d@�9HHF��i�|��)&4��")1�S,f�!��ɦE��$�do_2�����Z>����J�Ӽ��E��p�cW	���9\1�]2Q�21�ƒcH�Fjd3YcgK��8�� g'�.Ygc��K�3��c�\c� �"�I����.�d�F2Ɏ����	��A���4It/���}�w����5��c��#&jP@Ғ�5	�z��n�"e1w���)�O	|�i���d:K�'�P�1	�m#p�¢�I�c��$u�������<԰��c,��Lg���C܄�2Jk�1�=Le��	��_1�Bfp���4��q��f�1�
 ��dj�p�ȄǫK�$H�f���*�2�8}1ҩP���1��0��^8��(��2`�b�1��H�1�H���dA!b�3��4g�E��ڑ�}�FH�2�3(g�Hf"�R���0����$d��,e�P�bg:QƩ#�h�P���A#%P�gϔ1�3�eAH`�Y�3�,��њ1��P�崾���eC����(b=LgmDі>ZX�MD�`�	�Þ�e4��!ʆuaC��`�Ta$Rc�1��h�cE�(�����2	-$�bf9P�1�mFö���Q���D��t�e��@���`��Q��j,�hL���&o2�Lk��ؤqq��<��(�l/=ˆ`��}��d�u�c��A�>���z��2P��e�����C4f��1�7��=�3[�q^DL/�q��a|����d������Qe���ǻ	�5F��8��̄Ƿ	�����	p���x�-��u- ���D�1�c$�8Hi|�y��&�%�4���%+.�"�2c��&p��D�`��$�����">`�u�*�j�CHB؅�w�11�Q��\G�P�%�|оc[�g/�0����J��Ԍ���"�3
n"�#�E�r�e��j�8��8�J�c��)3](d7J0��(���CN�H�1�چ#Z�_"Ɍr��V@�c!ʆ1�d�Z!�c!چ2��c�Q��1�m`@�x��16�	n1�3�Xƅ��3r�EФc$d��X�t��i�1�(��aŔ�1:Q�<P�1�ђu&2/bc.�E�MD�AC�d���qc)5]51�f�w��	��Gp�D1�f�ڈ$fl�c��⏛HO�iQ
n�1�g<Qd�G|1�(c���F$�$�c0���є3G��at�����j12�������)���h�� �Oጒ�c(��1��ՑBi��(GCÄ3a��p���I�jaI̲I'~L�$�p��������FJL��,d�Bfo�q�1$�ĳ��}C0��%�L��(f��"-�X�(d�P�(z�f�#e���c�Q�Ƣ������E}�E󸁥bx��ڌ���Ysd�w�2>�Ql��C(��DX�	�FLC؈�8d��k0»�>��}#!�DT)�*T2�t�KH�
bPS�p�Η�k"*S,v�7�U��� ���d9��@��i5`�|��
T��SdC�	�wLC8��c��>\3F;qpŰ�3�����#(w���0�L���_1+�r��mF?��d��>P�(3�	�x�?����i����_�
(f���d֬���C�3��	9��C1�؆&�����k��MG��8�*#1�3;�B2�1��-p����(њ>�3MEAP�} �R?��d��QE?�,e�P�ͨ�7��_3Gԣa����8�}��C��jH�`�p�ɐ?�Hg�v�����c"��c��l,,c���Kq
�B.�;��$����#D>V!�6�X%�Ɖ|`O�2C���-���ԡш��#9���o�QP�he��ϘŃLe�KK;�e=ԬCвT��&K0�����p���A��K4����zqC��'�N9/�M@�
����)3Ne�Y
���(�"��0�H�`�c������ZV)�E�P_̽k ckN9�\<\AF%"J(:_1��
�Z�	$�c��|$�ńģ�����z�c���!q����/aI$�L�����*��T��<r�q�O����o���%}}���~i��UrxR	������s��9�m���ͫ��D�&SY�7S4�*�=�5f���'_q��[���$ow��'	d�����Bw�e�>vܩ���(<��7%�j����>�MY���{y{�a4޼�Ԋob����F�X;�r�ܚ:j����mKX���Ne{f�ǼC9�����M3��Ӊ�˧�6�����30�|�f�sľ�,4�m��[S:��z�E��NTF��>d>����f���(����8{�Y�dO+*�'��.���R�����ʵ��.N��b����d�Z�'&&��f��s;�[Sk��.̜�����w7�r2.�o�:��CoTj���w���Ȅ�mn��"p��ǫ9J���'ם��Y�d%�ʱj�~�N��j�R��'��%��?��.�BK	��CyǒC/{ӟ+�us�4X%f�s�J}l����ʢ5㌯�+ʙO��U}�<�o��{ezt{9`��
�Ζrr#03��KL�n�����"��f�;�����̂���8���Y��L/;�e[��^��k�]�ô���n7ˢÏB�yo9:ZޔZw��>��vs�����:v'd��)�Uuӆ��\��M���s�7=����7�׻N�p�w��W�����5�HW�����a�֮����ݘp�wk�y�w��?P��s��u]�;t����+�U�wuwֳ)�e�	>��3��ݙ��U��3ok#2Й��y��y��[�����j7;r�z�e^'ǳ:0���m*������~��7��E�,���-��nYY]wqYדFG�JI��J�r����^��y�Q}$�Ys��,�T���ɥ�-�O�n�vq�7ff�Y��on8۲ɩo�j]����I,SD-�e�؜�Iunr�Ku>:�S�s�ww����m=�
y�<��׏,ʟ���w};��|���x�F�e���C��f}�w2}��-���ǖ���f+����0�^pN���W7yŨ���fo�M���O!R/���o<�����-�ɋ����/��Nk�7�߻��C���t�SqS0�����r>]3��a{�K�{�����hOBВ�\]&���`�w�&���W���m�<a�.s2�܆<����汏(q��/x�1�.�Ƀ��,µ3yӖ�;�i�ɅϤ�k�˝wK�<����wX�L�ff�p�9�y��=�[����7�64��2�ݽ���Gν}���wr�^�������-,�fM����e����3$��~�+�3��M�3O~|�`�}t�s|����.��`���0��E�p�?�*l�����3�^�n�t��t����ֵ�ǎR�]IS��7�[)m���4{1��{�&z�u��\�\������g/��iy+}�֕�E��陙����6rzs:���-��"m�|{�`���\�����c���4[L����b"��xb�vܯB5%o�9���A�*���勳�[�sO'���oN�����ַǉ� }�$�מ̝��s�tɆ�fM�Ò��8rni����i�=5(�_mJ��M�\Jw�����ɚ�2�W�wwݣ��R�ܞ.��}�_F�'�e᜼���?��/$�?;S)��d�v����v�Ow�g��|3Ϫ_�d��Q�B�|əTw����kћ����1��.ꗧݓ�w�%�gx��d�����~t�w�5N]���=�'(6뉛=�Hf\��7��؇x���I۟]oOor�D�D��+'��$�'z��;"n�x���N��ɞA��aҪ�٣��)V��z������oN�/ӇO���'g�����{c����$ɟ�ƫ�\ӣ��I ss�V�i�l�"iŦ�X3+��hc�o��.:�/='���U�����G�����N��)�-r`��z���B\�$Ú��-ns��7C�$����y!��	'�+����p�`����9�o-8���qPk9w7��R�i�T����J=��\z�j�Eөʸ�Sܔ��^��3�#1��NrvR��f�F�U:rH���ۚ�o�p�d�	(NI��Iܜ�y0~30���՜ݗ(qLG�v�$ܓ;;����V<3UQ�c�9���b�}ɽ���e����*
���M�c�R^_2.\�'�I]�}m^Tm���1��U8�F���as!;72l�J��7+�����WH��y5�qp�Z%�kꙎ��^rǰ���w9���q���'�|U���og�`�۝����#��en��&m@������	�'_���?LÞ�M��mL��!���u�nݖ�{�����.r�)��� �l��n�r�n�]��\��յ�g�:c�2�����m�(�m����ƹ�$��󛜛�����j�s�l�y��=������'��������N�n�����iٽ���*j�=�=^�Q�n"j6��f����ϧ9d/mQ1����nv�5T˄�h���s+H��4��/���!����Ʃʌɕ�FN<�K�h���k����{�;�?L�?la��ޫ�Fm��iw��R�G�&�OyB��s�;ˣi�{�r�=���NC�fd��[bǤQ�gO�f��we�^d���8��S̾O��cZ�K�,�p�$�T_f��fn�}�o6�S��6S��ž�ᡒZ�s2�{�}ex*[��]�;����s;=�Ӗ˓��kwlUӗ̍Qu:�JM8�����[آé�>m��ʺ˫�l�Rj�2�
~�w�{9���3rE��m�k��j���ȭ��iLGwLUĭ:�7�;�T�,�EnN�)���**�3e�'O�-WU̮��]2����y�k�=�;���^J~����wid�^�B�Ur �[�h��S�7�u�[��9�k�0��ˤ��zʞ��}s�,���*T��?I��K�2r5��uܼ�4�}�-p�v9�MK��7m��6���'�u���Y�e���K.gN\�z������Wg��fOݗ�����	�Q�=~{�R�r�Ǹཙ��0�T�oH�n+~�TqG�s��M�s������\���T8�si�������=�y����m��݃͞�Y��\�Q�*�ə��y�{pe%�����o�ș�&g�Y:D�+9*����2�2t�(bOz�Y/�
�*~�+�F�s)������6)�����d�����zd���x<�Vr�M�vow=���s�e��{�˺�ۗ2k�ށ��b���wk*����v�(�EUL���{0���=���ί�`>�	���ʅ����H��	��輻�~ve�M�Gl��zs�ݺ:/������"D���~)���N�î��rw�n�r��(J���$n�Z2bl����".�r^���K�u�˩j��H��6Mu�T�.��ك�[^�b�ne�#9��[�]��F+�i�fes�r�G1�mM�ohJT��a�(]H�K��V�W784�nrm��#��P��"��na���e尘Q�81=�3��7~������R���NF�w7��L��X�ƃ��*d����D��a�vf�)"6�J��6R�&��̾&�V���Oͼ�܌���"޻��kH㟻�o&���f�:h���˥4�e���5�I�}�͕|0�.V���JV�&�����c��I���{ί^}qSL�"��]�x;1P�G�H(ݢ�G2e<�S^X�j�a����*"W\w��{͏Mi���@�b�1j�u� Mj�5�U���\���)~�y�������	���E���|�uJ5à�e���Z���g��,��W�=b�{ j��i�#�Q�h��������%��
T��u��&tR(RC�uZ�p�W�n�J�*tm�K�y\��Iu�����`֗�m�Z:�Ψ_>=����2��e��7Vա�Z��T���x��FXcgb����mR1�i�l���ǝ��30�"�K[�Lɖ���K�;+�{9�a�X�?[[J[/e�kSKnt��#}㘴����6*�n�����{��1���ɳF5�H�����V�q�Y�R≰v��#QOfg�� ��V���H�"-��lG�^�����4*Z�<JX)�寽ŀ�%\��6V+E)����,��̪(D��-?� ���@%Bpp��5�0��u�@;�Yc��� �"�ʦf5��u�vҎ�f���t,ٮ����M��%Wvl�)m�l�V3��Dm2HG���a�x�ڤ�SS4��{C�ތ�Bk70-�;QM�S���:�R���q�zc>DPh`"�A�\^�{�[���ezշy����-��j�:���i��Sͱ;)�*��<�&4ԊJݒ��̼�Z��m>w�
���^TW�'��9_���_a�]h:4v��<\x�yo0m	�b�d
ZA��t�6������R�a0z\N����y��5٨������y"���kkP�ѡA�\A!�.e�e�_K�22yѭ�����_�}��������R[���V�m�������Va��ݻv���p�����s�-��o��������#l%��	����O�%\�����]6۶�7��z�m���6�m�i��xۖ�n�n�m�owv71����m��m��|�m�m�M�-��1��m�6�m���}�{�����>)O���}*�B⪁�����>.-�bm��6�۶ۦۖ�op�m�m>i��i��m�M��{���Z�v�r�m�nm��m��|�m�m�M�-��6ܶ�x�m���6݇���k��m��6�m�i��o[��n�n�m�m�m�m�����m��ܶ��ww[���xۖ�t�n�p�m�cm��-�ݶ�6�v�t�n�m�n������� ������G�m�cm��lm�����xۖ�t�n�n[m�m�m��v���m��4�m�m�m�m�m��m��m�޷��z�6���}�q���Ψ���EPHR�v$��f�V)�/[��o��f�)5M������������?s��=�s�ޞ���8c�$��(e(�# �b$����e���8јp�ƌ�p� f��M�,�p�H�@�1�1� ��I1d�҆1�����8��n��E�t�F���X0`�!1��d�c�6.H��d��`��bc8�gb8f��Fp��b8gh�ƘX�c(de�1�i��0��!�0eddGN�}���ïUW�����.�L9�~�8��W��K�Lh�䘗։�!���|_���د"7@�p�~��<��y
�����ה	��j�Rn��Z�N,f�`��F��fv�h3u����wl�+P��k���,W���e����k�(ʑb�݉55�Qۋ��g`uWi,�L�m6�-K����@uB���z��8��c�XRm%vܨ%ىd8͝x�dii�L�����K�R��l�	h}܋3,-p�ȣ���c��!�u�����i�DHP�
��?�R�W�5�kuŢj���\K�+.`�5���^Ϧܵ9+���ɉʕ��)&p�b�vS��Z�\� E�mv�	Va�.�R��f�bۭR\k�Sh�ik�J~�6'�&����2�e��դ��#5�5ᗩ�5s����S�cmk��Zڽ����h39�4ln�L�ڨ@��hVѺ��fkF�Sfh��}��B�\6Jp���2���LG��Gn\�T!^��?y������ޞ�R���{�����}��}�=J��=�{���www}��||��{������x�睊`�O<��y�]|��a�I'Y�0��~��$jPɪ�����h�{��g�hq��
f�[bB�F�v��:!�O�٘_p^����0=aޞ�+-�4��Y�nR-X	`��'��n��[��H[P�`�2VFW������G��	ѬiJa�2��[�D,C�2�����F��IF�������9�d����S�i�N�RN�Ӊ�uG�G����[���~Z�F��Pu֊����V��A'�޶�i2m;�cC�~O�W[F��a�u�u�ξe�u�XqƜu����$�S�G*�_#lխv��o��Ͷ�tt�����ɕ|����d���5�k��]ܑ$���i>�C����<�P�?L��B	��"�{!OX�.[��b"Nчf;0�2���"���.��H�-��ьc8f��FH�H�8���b�Q)����h��@��|9�g|�LF�/bA�;M�$y�;I�2}\�|��`�����nn�e�wk��1,���3�Ս�~^�u�q'�H�r�$ql:�))l��!�F��V���%0��i0��U���:�ZUD4î8�<㯝i#$c$d�qg�j�$!R���*���:�lӆ`V)��8^���VA�sx����61��F��Ef��Ϡ>u�pO�$���@�p��8�jj �NI@Y��qS��'��]'��uKkmø��26Y����
��6M?)�j��y<�@���C:�e�Qf�p��4��1�2N8�����f���}ec��d����MD�D��Vl��]���%"��s.h�aQ�)VDF�I��'���/�bJ�ĥY�\��m��[��C��j�eZ^ah�[�+$��n��m��U[��j��\(�rG>]�{�保;�gGIFu�,iP�*1��҇"�-JR~Nt��\�R2���W+�0]�}K:�}���C��C ã�q,�"��Q�!�q>�ݫ�&���ȓ�]�]t���!���ilc4���aF��qm>Kq3�W����%��*��}dP�8�3Fi#$c$d�<?��EXͤR��$��6%}%m�Z��l��5�b�K����m�J�F�'��M����N�-w���12��of71���`+e��T2n��l���P�{��Q+�Bzi�4�1�lX��b�s�;k��[l>m��u�_:�#$c$d�qg�qj�A�����J��=Y8�S���蒾q\O&қ�Z�֫g&�ikUK��+�X��`2�,e�����w��E���?;4NwG�?1�ɇ��?C�v�V���s��i{��;?u��kkP����I �3R���,ь���4��1��8ӎ��K�u����-�{ֲ�/C���Ό�&��������6���B�v�.���e��9Hy���w�}�DJ�>�*e)��Uɷ)�ԕ��p��U�{�~s����#F"-�+}���n븦�;T�o&
~��s
4E�p���0d����r����N��K��׏���Zԍ28۩�v'�����\&y�f��=�k�,��V�Fo@�V��J!�WF������,�:W%�}�����q�k`6Rd_�Sq�4Eʇ��{\�ê��F��4nC�y����8�f���fc��ՃU����-�V�O�wx��c�}ڊ�n3�!f)�v���,p�̝Na����Oӝ;��sÐ24�ݺ��5�����j���rH�W���In��dIWn�i�[�\q�u�[�!���qŜ3i)V�jE*Sx�a��q�ta�CM��ɮ�&1�L^<��a�b��N�\u��I"8r�UR)G0�zT���aױ��/vS}9�5��vJ`��/����v��[�{�(�u�����k,��,p�"�l�5+ϹI2o�yu��l�\I�>�#�[�T���{�_���������g�2���Y���:#¡zr���wŦ�����J_G����������/���y~L��'έ����aN�_Sζǜ_��/�8�����K��|���؞_�y�'�//��_�K�xǓ�y�2�>k���_�y���&�/��ȿ0�0�O)䉢i"iKKM<���<�-~ak�_�_��������<��/�ǖ��1i�x�m~O2�&_�~^�?>�����1�?:������:���q'_S���8��������'���V�>n�b����a��R�0�4���</���|����D�M-o0�0Z�Z#�ɗ�c//	��$��R���������k��!�7��Mt���CUE񨰶s)n��#̦W�s˚𪆽U�,Y���2�+�׃�����\M�I�Z�a~�������#Z�<s�����<b��������>��T9<'��:&#�́�g����D"��b���(pb�|����߲v:]N(2�|?�о����o�ۻ���>���_������x���{��wwww{Ǐ��{����������<i�<3`�y��4ˮ��ϟS�I%B8����nY3�[9���O+	I�vD�H�g�r�gv[gU��
VЌCw��U5H=��[����!�`OR"I����z�R.���(G����P62�T�dY�*�aSkv��X|�z�@�4�'����N������-���5�P��O�hݸ�w7��<�	���Ad��		ס��p?})F�O8�A;�,'L�>`vQԥ2�������N��*%:!F=���.�\��C�#R���~[iU]�6��_RQ�JT�e���^y��uמ[�0�L��n���i˞I$�BI> ��y�Z*)�B�-R(��}Y�u��$���J��u�EϷb�sp՚�g ��-L$;�P�d{AJ�,d'�eoz�{�)ne���t�����|������<�f�����4Da/�!��(���J�ܪ�#+��Dz+u�m��:�dvt����%��N2�IVS �[5*����rۇȈ�J���DD����,I������ Q�O�J��9�*��V�0�4���矟�m�N���y��e�[u��jfH��Lf׭"�k�6Y���&n,ug��J�d���ff����U���-}e�;1+��S�ƙ����KX���#l��n-���Z�b=�,cRrM��� BFY���ߋ�b�y+R&�p�ӢgZV�[zWa� �u����_S_�]Q�""����U�o��[�5CԊ�*)��%@�H�2	�M�O�'c�@�F��D@�y��nb28%W�\�!__��ʱ)�"���;IĄ�N���?r�n7��T��8��Ԫ�GR�R�P|�[E_$�����j�jSw�K�s俳[�tg!�d�%��$�8QN�`Q��2T���B �ė�<��z�օk�r��;:��mfý%��ԧǜ����08 ���D���?x���# �2v�ȉ�g:�������M���~u�~u�������<�.�ۯ>o�Z��z���$�(�B�>�����UQ�2�:��K���;�
l	B����2��Jz2��ߊv�qs���L�"I�C$�|A��ܐ�N�`oe<���&�А��嶂��r��ˌ�!3���N7W	m�e��FC��!RA�"'w�xe{�}�ׯhM����[��s����y�hì��A�4Bϥ����-������̌�:`�(���&0P7�L�Y9��1����uA>���K�ĵ��%=H^V~��]UW�J��e��q����t��-�y�]u�^|�nU�U�,���D@�����lz09�	�aa�uDD�İ���lt0�A'�-��B�����@ӒId=��`jE�nI�q0DO�K���00B���R��F��fim2�n��l�Kw�V{��v�����Ry��,��i�'BIz��);ȁD1��w{>n�np��]R�]���bRJ�~r�d؁`����&��a;=��m���"'߬��'J2N�XfD�;,��l��?~���3a��"#$�pIK'FHq�Uţ8��1g�v�>m�������t���y�i�]mןSwR��"��2"N"�D�+h~�� ��ؖ�_���U��'�C`��	D6m�
��^I�(�NWȺ�TjJ�N�C�	�J%C�ѐފ#2{�-?kb�D�(�W]�p��&�7y���x��k
��aY�K:h�L�)�d��5!FI��T��pӂ풖��C��'�	`�xk�<)'�a[U�.�J+��ȼ2��%���LҒ��D����Xw���2��C�Z����g�ѲCa��v����82pd(�l�&>�TU��0�`�>螘�@�8!���A5�IL#��^�`�R���(����8���מ[�0�L��n��|����c����1�VZF�W��zi��q-in�akM6��j��!��M.5�HF��į��o�dmKH���ݜR�K�55ذ��b��u1�	�'`��1��� K���zp��(���ˍ	�*(������]����'�,>L@�g �~I���M�a��@�5RUAB)^BSXЕ�	�@ϥ�C�<��M�!'�&�	� ud�Zۤ��w�f�=l��Èu��LK���$�a!`��@҄�C���[nC� �;�'iO�~��nH�b%E���a��0�D�!1QC�U�"H�S&j#�q*����JCΏ�٣��	�v�=('g>:�{���G>�e��=�9�ƶǫ.&��Nf�32����A,���$���8�O��"��I*ڨ�G�Jcn�O�:����X���x�'�(c0g�&�tn\aqw��UTBy�y�!�C�5�a_���[QH������f#��T�6�����K�/uj�<	I|T����S�!�)a�o�V�4�"D�� ��=�(d<�a�aU**�Ωe���DL��~��S�)m�_wvqᎭ�j�wm�Ή��P���F���`��!�0�J�?gߌ�ɧ�d�0Bz��L�{
)4N�PMI�)繇㯯1��8�T���_V�J���O����~~u��:���y��e�[u��=0���C��Wa���1*T��1w"��LR"EZ">��G�k��(m*�L-MkWѧ�������v���ڒ��JB+�b�޴��L;?�3�K����3�jW��Ny�+^���t��Q3�-��!��!̦	�J!���)d� N��;4v�^ܖ��">��Z�vH�4������CL�g����>"�f��X�BR-��jJ�0�"����2�1�h�OS�[�:���ζӇ^yo<��2뭺���vkw#3y��%$����tn�U	�)�?R�X� �![E#���j��M�"��m����2�(��ݓ%�GP���Mÿ"�?D�s��E�.��W(�"6��7�-&C�tXp<�N��ȑ�^RڧmZ!��~�=X}�(�ƚ!�&�!̟CJC�?�i�_���n;�x������`�r�=;QV�;�K�߃�֔��ߖ�<��õ�p�WJ1�1��ǉ�g���|i^8��|����<�O-�2�zO0�0�O0�x�y�ᇘ�y�������'�b�Й/O�H��<C�ǜ_�_�_ϗ���y�\G�_�痧��c�/̯���`�̿-������~e�������y�y>q�O�K����i��&�[C�NUWJ#��i�}�/�������a��0�Ly�_��\�y��<O�����_�/5������~~u������~a���ח�{俓�!��fB�^ �Йq�h\x�=	���[O.'��=����K������_Oj���콞�6_b�\p�����o-��ixu~&�~*{�'QO�n㒺��]�ܥ�Q����[H��T2�Y�beqE�}�9�'�=��`F�TT�7�����|��Z��5�ñ�q5�kaC[�g�1\���2�
�e`�fRӯ@��K��FO>����ǫ���.o�ҡ����P�۟]�[�^јR�����$����0�l�����k����/�j鵙����\x��$�L�R�]4���פ�=bz[C y�s$[���͗�|ȅ�X*ٗ�.<d� �fM;21����Ϟs���"�ͦf\�d��d�f3��_^�0��._{7J� +��U��@5%�b�w�'6����'ܛcd�͙��J�}�P�>LdS��i�w���<'����cb>ɪ}��L'�@D��{�D�u_H��a�{��1b�;�~�4-iԥ�sh��-�ФQ�F�-���i��3k��L:�ǩ[e��v�YA3P�u	���U\T<�hY���
ƽ�JC""x��E�BG]�nswYEL�@�a�̺ͦ2DRV@֕��е��uPIP��$zi�cXc�]?aa�����cmP�P&�;�;�ү�w�i�S�z;KYy�*]mg�s��G3r{4�ǵ2Z�ٖ�4�2�m���V�>kH���YY`��$�Ex�����������������k����{_www{�M���wwww���m��www{�Q�`��38�x��P�`�I)Z<�S����!
(��H��=��D�K���KWX�c�vRi���z,�'��o^�Q_F�[hV��!��F��q�z'�}uokf��sR�r��@2+ٻgo�Ox�T=�XY0�.�s����� �񎭿�/�5&Np��3�n�|��a�c0�2O�Y�nР��_
Rژ��cC�}��R'�<�O���߫j��Dg96N����o�6}l�i�E��A9��p�K����}�Y�$�~_*�c�#��+�t�6�3N��3U�]�h�ҿ�$�ճ�Y�Y�R�E���6Q�i��A�^3�2��,-�^~~u�[iî���2���n����i�|��I$�q��W��U�v=K���s1����)�� �WK�I"-�͛˻�Wxٳ�`�M�R0��b��VN>��Y��M�N��҇��;,�2��թS�fm�p��#�9�Oƅ�=�өD��k��t��M��~8�r��t���m��u�M4�����n�[��f���D��#+[��>u���p���̼�.�ۯ>p��W�v�S2�ԒI!4d��I"w����a�Ɇ�]=^(��ŵ$l�E�T~�1Y�m����E���y�}[�Ɖ����5㹫U���8�ٹ�J�㸥��8���gg��B�xP�Vw='��eÈ}��w��e4�~��ڧnliNv`p0Ӆ>2�k��0�)�a�ŵV��|p�>+&��$�]����0��~y�~u��:�?<�/0ˮ��ϛa��w#�I$�<����n�b?UaI��{5�6O��Ԕ>�/�˦F�Y���qy��-�{�#��R�Ԗ��K!u\����X����N�p���ˇ>�=���46dcؤ��O����SHx}�p�"����[��8~�a�%O�p2L�2D�e�ʔH���e�n%.?>[�<�?:�Nt�<Q�FX��ML�	T
*���[u���M[6Wm, ^�!��L�v4WB?�CiĞ"R[��k+������o)��Z�m�"�]�',�f54z��Z��k+R�W�?  !'�oB�*�V|�5�2�ԷS��ܹ��Xw��ݞI�΄%0=���:o�wQ�U�t���w2ME;'㩧�g���aϞ�V�-m��>�Tj�b�]0~G;+�4C��|�VM0�-�9XE�Z��S��P���#�.I�Ue��묲��b�R�R�Ҧ�c�[��ݥ�W�+mY>C�}X���<���`�U��M�FԬ����io?8��ζӇ]G�y��u�[?����H�UUQ�a�C��U�*9MS�۲��o�6��;'g���::�ĲW�����3qY�K��!�a7Yw�SUQ���(�Ha��>�dnv&�<�!ԧg���&����߸sy���;o�\�.s0��)�x^C��W��{�_��z����5�&J��9Y|�-���,�y#O��NW�6��m��3����1�x����3Ɯӏb�UQ8v�[�D�r��]��l�Y�B뾓,6h��2�}�֪��~N�T�D�_Ϝ�-𕨲�1 VX�S.^p�r�ۜ�N�aa�p����ܚ'�6j��N}�~�����%�w�TT��%0?Ca�$�a�Q<�r󯅷Xe`�X��9��j�\�-�P����y'Ӿ� �"�S����G��8g�ag�x�G�c0g�g���㗸���XYx0�;%���d��"ϐ�1��./�>����l����2�+uWsC�|�u�a���`���R5N�7r�|сj�a��Y�<�~�%e�~�04������}ĭ�HI�<)����s.f~�y�!�>�a���~��w��3Sn��V3���,�c�(�C,f��ɸ�����.�o�d�&�j@Wޚ�Sǥ�M�G�t�#J�D�g;m#5�,%��޺�e�J6�0qf��v
�٥��ͭYS�ĵ�z�/���C� H8Hi�Khթ�U�'��x��K�[R�Ǘ��M���'�<:�pó�ف�ae�T�I��~d��$�q��,g�(�"طƟ��4��G���U˟Sfm���3��o>>eˏ�GA��Տ�i�܄`��Sֽ���T�"����>f��˻
�ǽ����?���)y���<e�u1��<�S{���m�����ָ���M�������:�Nuy�^e֝mם�S�?�z��Lp�l��;���S����ْ|�]<��?|t�+
xttvR'��>,��;�m�atۮÌǭ�)z�&�����魯Q��wӼ_{Á�K(p:�&BM'����~ĭ�cV�qq3M\n���-�˙�8g��ߋxhw"s�Xp<�����?65��g(��=�*�Oϟ�ǜY�6a�����B��ۋۭ�������3���y��<���~f��w#�0�[^��.�\Oy���y��=�/��cϗ�����:��N<���˾<�����'�/�/�״�k�ˇ�i~OI��ry�0�<�2�'�^e�b��<�\�y���Nby~>>3���>�>�'���S�0i�Q���F���-Dy#w<�-~b����������<�=so1��1i�����<O'�痔�W<�l���y�?:��~y~~{��'W�������q��<�mI�����<�N>y�y}}s��4�ʞOI�����i�㉕���^!�D{aD#�qx���Ǔ(��io-�[�/xVx��ȃ��8B�L�9P�b-X;`n����>B)��T����2%��>\7l�z���v���9i*��S#R��-֯����D^Y;�s��O$���bgI�D��b[����g֭ q���x����r`�Jng�?����{ݿ����{�Ͷ�o�����/6�}�������m�������p�<A�Ox��Y��!�y��u�[u��r��$�!�]}&�݉Q����L�&(їm��&i��%�'��^$�d����?����7)L�J9rۖS���p�}à^p�!ПS*<��p:���	��Y~����[tv��$e�?Q�<��rMV뾒r�$��d�7M0�_8����in��:�ʹ��Qמe�^i��x��~x���UTH�����)�&��}O�R��NӚi�i��#�[R�j�h���Z2��zךi.Nyl~�֜�WWO?P��j�n�:�agZ�"a�)�u�Z~�`?}
���i�~���V[Ma��9�A�s��7�J�9m�G���0�2�xp�p>9��4����e�Y�L���u�1�t�v�?Vml?4��8��Nuy�^e�mח&y�<!r8��(��f?�-�'�(Nz�z%�=P�͹��d>m��Z*�O��I���(�;r����r�Vc�������$N���;���=IVd���/�[󑰘xK�3Gi�q�jM5)1(v������1�'(
}(�� 	4�4mj��4�������lM��KM�h�-C�E��w"p��v�ʶ���2���ID�d�2T0�p��>|m���"��ћ{�^S���i��O$��Y)��0�,����s���RtC%�0�k�m/�`�f6�jX��)����aڷ3gO��~K�j�]y��,���L���Val?8���ʹ��Qמe�^i��y�rK|��bI$�z�i�]��~�@��u\�0��Xl>=�M���S�λ�4�"JH��+,�S�
`�Y�	c>&��.	���_����M)˭���$+e�U����j4k���C�����M�-f��~�^Z���)�klӎ��3�}굒~��5hw�����-��κ���m8u�u�y��u���پ��ql����{UTC�L��M5$r�ҷ]?3�I��i�穆{^ｍsF&/_W�S�ǒR,���壅?Ӏ����-{��7m��1�7wtw0�h��0�އ�b�
OXy��uwWi�d��o	R�~F��!�G��ZR�|vw;.tɿ�~��*�f[���	�h|xk��y�ۭS��q��[.���:�Nuy�^e�[mן6����a?"�4�C���z��=,=�k���|2�?m�Jj�C�k���0p�Y�mu�%��B���,�G�U�l�P8HĚ�ˋص{�p��e�*�t}0���.�ϧ���Ti�XY��T0�b�y��P�4S�l��vt�����C�$�����,�Sx?~�9��i�R3r����$��M���ۯ�<��4�3��xf3Ɲ^������h�4��	mٳ\�l��Ufb��� F���\�h���,[j��JV푣Z��N+�t���Q]�c���{��YMy:���P&Ɣ�%�5�<�G]3�w� !#!��|�UH�&���[��9F�	�|��C�=M��pN����(�l��i��a�Ze�����?\I%J�:��4���>��W��U�UY/�ʬ�H�r>a.�N��2��Yz���Kaf}�����9RksqéK-KrM�dĒ�i�i+�9K!n"M�j��i�>]���y��<�ʹ���2�/:�n����I�V�H��Œ)�L������O�����J�am�0n�m�#-#L����<�l��釱:Ք-)�{��̾����KD�}�?}�Y����f��Ҿ�Y��� �P�,�MX�!��N�����u�ɨ��tƔr�7�&��FE|�gjW��Mk���SO�m��\q��h1�c?x��,��4��{g�U���UD6@NS���8}'�d>�Z�7�"8�-��EX�ȱH1AR�͏����$C��Y�?vI&0���� �9�!~��Li~\3wv�2�G6�ÇT��Ð�iC��'��/C��ڽ�
l�i��u}矻X�c5Yj�B�9$[��һP>0��SLC��E�����i��\a����i��Q�_�^4��p��zw�����e[b�}��<UTA3S��h�8�rND=޷>L�T���i��1��2��M�K4��/��Ǝ�(t&@@Q����~�pY$����K�jr�!�b_�t���RSor��K�\��Ǜ5����1\~�4{=�����f�l�U��;L
JR{�4m���g�p��>gNi�a��e������8�����8��y|{��r�O8����k��y�����X�O/)o.'�/+y�<�1�W�i|O>_�__�_���G��<���:�u~v����1����4�q~<�a~y~O<�<�<�0�'�^�b'�4ǘ_��֞c>c����.q���.2�-�Kyq�����ɴ��j䵦�>��ό)��ʼ0��_L/���<�����<�z�˷��^\y~O�����i�<߱/�y�����=r~~_���?9s����y���֗��_�_�y~�9s�bW���&�I��<�'�{D��b|�<�'���m<���bT�0����0����zG��J8�zRg�r{*�.�R�����*�zf�w�u(:���7U�ZB6��Y���s�p͟��&�wI���Ȧ�w��\s1<���mq�1��vM�	1<�Ր�G����=��ݜ,��)Qŕ˓2��'�س9��&F/�u���ѵ5�Mor�E9'5�B���<�&Vn�b�ND�,s�Tܮ��(X�n��3#����Ǐ�s�y�E�'*!���]3j����&8�b*��1��RJ��p���sw����٤���v�y3%x�*��f�+��]�"Ť�w E�w2ls[o�l�LN��T,�}��r�޸-��ӎ3��Ϧц�+�Ǚ0;��rq��.`�.U-z;�'rZ�xc>�-��Q5�W�G.L��QKopwqe��9�W����$��,V�GK1d����b�����vUr7c��*��?���m��(.�J�djD�۵�)�C��6٪�Mo[��JE�"���a��Ա"�U.1R��Bk[^�kuq��4��%�:� ZRdl�"���tݾ7�5��6SK��fud51u�e�~7M=��#<��ҳM��Ѵ2f���6�Y=��_��MB��)�u�Rd�)1v�2�ŗ\[di��F`q\�#[v<rW@�AjR�0��>�ݿ�������m���ww{��y��v�����z<�o�}������Ǎ(��8�Y��!��G�<3�d�#���Q(��U1$�HY�z����(-�Z�f' �@у�܉mx���=���U\k	�2錱6��us)f6����m�nZ��?h JgY��^U��n�c� ����]Y�*���jB��>�Uv��#�S��7L�|�e˻��v��W�M�Z�-���i�U�L��K��9N�&�m	]E���8f\�����T�V�%,=�O4��
z|d�\��+l����@��ؕ"��?'����t�ی�z��b����Ϫ��K��yy�z��Yy�]|��>i��Q�Xy�^u�[z��O[�E˭I$����S����ߏӹ�)�<^���W�d���1L9r[��i��ѳI�mZFۯն�7\̚���=Wh��!�(�Ʃ��۫3��j/0��HJ��A�Ti-��E��ⱋc5�mΧ穖��!����M�(�N��;��A!�I��~��?S����;[q��m�\~~q��Śb�<x��0f2z��:#�Np��UD9�C٧s9�9���Cס{�I�gA�
���=H�rr��S�||i�K��gd\"w�x�4�btu���~�����wZ~i�wQI�����w�^�|͇!���	��X߆)�à�)��`w?C<�yUa֫��2�����~̝��SN9�0��.3�?Y��!��Ǌ<3a��TOF�ꪢC�y�+Y����%>|ˋ|��>9�{�1��~%JQ�G8ќ�C��l��ti�h�s�����~��˔�2ۈ�-�f^�\]��X�q�mcO�k���=�)���3q����Ӣ"g~�������f��U��ukZ&��saJ;�rM$��(��8�Ɩh1�c$����xt�a<��D�"�*b��
��X�Y,U��,VAV|,	\[V!
f�͙Jss1�#��v��2�S�zmc���n�$�z�����4W�j\�u�A�_� !!��dj�]ohn��m����4��S���鈻W���}�\�-o̙1����)��Q�F����H�e�uo��ߩm��U�q����U�J���}D~|��1��m8��a�|�=y��f-v�s3�d�w�ϳC��<%Ik+,�d��7l֑�_8�/?:㎾i��Q�X~y��m��qZ��V����I$�E�ì���m�[배�!�%C�FS�d:;7�a��hDu�}[m���k�٧�9��3���SN��ȕ��a�ԥf�A��ˎ���+�)�Jٖ���5�]��ʄ�/�0n&�6�*<�Z��L!�L6e��4�9gFtY��)�h�����-���+i��^u�~|�A�C#<Q�2�+■����yC���~�Iy�>�Mӥ�ٷobz�M����DC�[�Yњ�0����p�r�q�㜼��~��"�q�4��DGnkjw��ԧx�,��!L�B�g-0�|�?/�P��{<��4��D�������i�
/���;pB��K
}�e)���m.�h���^n�u�$㔋m�ŘQ�<q��K4�1�3�G�`�<k��R�Q>ĒI?I����
�>����#$oi��R4�,b�W�����������n��չ[in���s��O�9� �����i��F[G������x��ڶX��8�-�!�/NbI�z�-��Z~���I�7O�[8�ϾOʹW�S�S͇bi�Y��a�d�4��U`��i�r��8ӯ2��8���u#<Q�2�-�u4*J �IFbR'$��f�u,m�?�5c��#�=�x��N�S�[n��X"rn�S�%���j!� 
'[��J%�	bhE	)U�� ����ϭ,�V0iƫ�n�݇GC�;:�9Ǣa؇�9��c'�iA*~���"}	J��K�'Ͼb�X�o%a�Ԕ���0�2j�at�-|�>��ii���Q��sO�O{|CJ ��<�<,�C6����]ی��xL��04ƪ���6��MQ���x�
���e��
C8�q�4�A�C#?xf��1&���l�b)�1����$YؖL�L�0��UD�-_�)��=�إq};��3�:��Y�TGr���?~��&&H'��#m�ã�|9��G����!�$���JѤE�Oߤ�.G�=��ғ�2�p7uc�il�tڕ�u���T�[������S�v7k���Z�L��}�6���J�}�D�7R��u�|�V�ߎ<�I�~4���3�13LeF���IE2D0`��iH�Q�0c4��3��4bƌњ3M�4�(���1�f�c$b� ��11�p�Qc�1�@Æb0e�4�#G�>yo-岷V���31�b0`�2qC,����ў<1�<x��hxќp�$f��3Fq#8�
,���$e13k�Lga�Æ4Z�[+t��um��e��ܩ��7Db�"i̖-�0�n߲�)�^�O�|���ϩ�ӹ�Ȟ�{^kJ>�f6/#��Zms�iw�RJ��˝>�]j���®e��:.�ɱI�Ź�38�˖��Z�j��	�	\[��:�l6�JpꉺU0]_,�d9�&alYӕn
�����W�Q���{����W�@���=�5�I���)�][9$V�{q�C��T�Tm������ww{�����wo����{������ww��z|�}ݾ����E�<iG�<q�4�N���ï2����~ĒI���S	L}��6��k9G?8�4�V�`�ԏ�Wi8�W��O��q[�߭C�ޟ�X�&)f��s1����}4}^��U��tS��?L�6N����%F)�za��#'˫O�Ytm����ߤ��	L�W����n�;ԘÍ�r�uT�ks��6��2���?Y��!����<3Y�z�9�J^N[�,ў����C�Q2]N��J��2�a����I����LQ�M/棛4QR	�m�������g��!#8u���0��L��v����u��B#,⟚cze��
�����nn�y=���g!M1�0Ѷ%Hè�&�)�O���F�N�
PaJ{��a�f�[ͼ�/�y�|�㮣������x�s�\�ddU]J)R[�xn�����"[#�^�6�r�+F��*�]v�(���$��x�s��m�ˊv�k#Ii��k�0��v�
��"�ں��텏V����� 	i�i�P���D�L���@�a��Y4x$"�F�JX˔�<���ǐ�>�a���'0D/�ˉ���}_x��c���F���>�0đ�;N�H���&������H�s�&�'��Ķ����r(��pOM�Ç<[!�G�N��Og�V9�-���^Z�/2�-5�`ױ���{;:4�9�)�i�Zj^.��'|�8�̰ӎ8�if�b����0��ƴ�3UU�Q;;=Y�S��Cվ&i����I�ђ+�~n��)����aaN���(u��2S�C�,=:&A�}�Zt5�s3r���5��؇�a�"���ð��Zr�2���8
Y=��zzp�۶��NA��Y)�A�2�?8���b�'�u�^vGb�
�V%�\���\5�=��I8�09��UU�_��lW��p;;0���(ɐ�(3�װ�Ɂ�ղ��C({=��2{�����f��J�1k>t|a�F�p�!�lO=�a�S���nW7O�|j��~qf��-_r;�-q)��hp�<2L�{��i��W)ʯ��%�>]<a�m�Y<1��Ɩh�!���x��i�%�m��n�E=�UQS�QDܟ;�l�i��t��)�rN��`�_ۊL�V$���%.����{OW)gi*�#��%>��K����-�Ub��)hF	U�e����#'�`�mu�ۦ����Z���g_���d��l�˦t�g[L���C���9Xa�M�+[m���O�q���p��'�f�0��Qjg�ә�L�ssp�*�g�ɵ��d���J�\�[}���Q��~O�4g�g;�4=��4��y���>����6���/�=RX�,�5-a�����=�9F��,1z��B>��=���du�*-�� %�uA�e�П�ZgM�e�Y����_��[ħ˥�*G0�:���a�)�)�b����#�����΃�EMM2yt���.fUv��Y*�iG��t��r�L��j��7�$�@��s���v���`T�3"�۸���Vޭ6r�{�˯��ifַ�u���~Ǎ,f�����x��i�|d�����ۢ��������=���G�p��/��)�'>~wGwqМ���Ժa;����Lg9��v��8�-�J�|�t���:�	Ny�4�	LO�����5��
��Z���L$�3��������̳S�st�6|������Sdeb]����嫈���p=�&�g
�֘}O���-�7$�6j��a�oaǆq���h��#<1�x�bqq:��ݒI"f�e���RE�f?	ES�w)�-,��~_�Z�]-��ܯ�f%�ߚ5ո)N�S ����p?Oq�+�W(՘5F�ZgP.%(�q�(���[f�d�c�Ի��^5�)hb�a�r�ik�&�,����tX}p;"0��~�u�˙�CO��]y�&�#���F_:�㍸��?X�#$g�3O�Q�[l��c�ea����@��W��U��O%�Yŗ��a��E��`�����8F���G�+pNq�DZ��40�p���evmZ�C��:8b�.>F^�ѹ0l���`���d4��KV����9� �=���N�f�m+��w3K,��S���f��il��~]�U~��n%�>?R��,2��[�m:�J4��X�13KeC8��QD�2D0`�#,`��,ff���q�,d��і3F`�8�,$���1��c�c$��1�P�X�7\u�t먎��GN�d�F�Dh��ǘG�GV��u�]`�1�E�0`��d���ff�g�3Ǐ�M<#Op�$gњ3Fq�҉,���$c,fg�8�
gA C,C$CI�)2Fq^J<�*9=�����,F�p�����d�F�8��E���V��	�w���\�T���⥘�U��r�!�o{��To�.�MZ��U6�k`z3�d��b��z�o�c�����P�y��J^Y�4�L{ :Жh���#���f���;3���"��I&�XB�'ϑ�s����`�$�2Q��I0���	1���\ù��Y|0i�7��;������Q�ec�k��6��Y^�)�x�G��φޑknGÛ�}��z';�w9��YL�);s6�Q�(J��nd����
�廓1ڮXb#�N��^��v�䵾�Z�}X3V\Cka���	�bL	Zv5&�f&���PB*������E1�Z�+���V��+ɞ͑���ܩ܌��$�)�Z�\��G祳"�ѯ�\\���jݱ�
�ڵ�͕�q��,�\��bCkeИ�����{OE/��K�s��g�N޾�b���iu8�d��޵��m���l
Z4ٻSm�ذ�S5�ܠ����v�*5e������؎6)q>y�,5�Wإ�C[�272�yx`�Y�u�][e5��Tl%lF5�lGP�Vʹn���"zۧ��k`gn���alcL�j& ��$���$�yX��ww���x���m���ww{���M������{����������<a��x��Ǎ,f�����3����+��O��b*��T�	�[t.��\�$�$*3)c��2驫�.CG�C�k}�6�.���|/���Y���}�ю�N����0����X��i�x���b�!��S��6}  ��Xb��p��@�O�������f�:�m�.�)�m����q��ww��G����=%�4uRcKT}��4�N�H'��|#.}�%�頇�v{�ge��O�!����Nآ*������= �s���~�����vڪ>�ϙ$r�W��j3g�8w"S��I��a�Q��b&I���~?3�8�h��Ì8�>yozbZ*���s.� PG�UD0���C�T��E�So�FQƟ*��۪G���߮���T¸f�o���4A���	�p��������O��!�J	)�0�ON<;Cm��Ҍ:�$�����t��C�g�'�}��;3[��뻶�?W�O�i��WȰ��:(s"{%���
[�n3;�?7�� ��ƌf�?3F@�$�N<q�On�"�L	* �$�H��m���|�8��PᏣ���{=0܇#�$�|��2��D��Q����}wL~i�[:u���6��x~�'ގdp�N��VUϩ�$�IO#����*�F�v��H��7_��m9��j��?O�L;�w�e���B|e=O[[I�a���:���~y���'qG8�G���51�
��/���l(g��0���!�a��u!��;<��53�����m<��U����oy�m�ĸ�I�ݞtl,OD�I�M�.\y>m�`�6�#T�G��ɂؐd>9K�X��l)8p�z�g��{K���R�=��g�'�B4�u�Y0)�~7'��0���N�J&J��2�T��[~Z�i��Ϳ:�>3F2N$�<q�O}�F�v�ww�x�I$�UfadDO�ISu	�\:�B5��s�,t����ir8l���X��>$����y�3A��vC����7���x-�;h6�+eU�Uw����nqD��=4�Rŉ.�a��k�M����*��Ow�A'���)���E�r���4�'��ͰƏa)�v�H���g�+��S�)) �&������o��%�xu9Q""aN�y~��L�!ê��OӞ/�ATgN�=<{����˙]��p�33[�a�6y��a�(��9U��~��%u�\��A���?~�<h��8��8�ǧg�~I���5Ȟ����a��JR�Ԕ��a�(���)������B'r���fD�Jעh���N�� �D����;�*�_�k�+xyTq���R�m2m̹oG�R���Ç�<9��/w�79��M0�d��aiH���.�}���GR7	��x���g4f�d�I�vzzvzW�k���zUX�K
�8�1/�--���%��w�����^�i��6���:�}O�F�O�>8�]W�t�]��mq���ZR��W3&Jzd
}��D������7*+�+&����������u>�jK��ӕ�~�h��.��'�O��s2p���L�a�����ag�<i���Fh�IĜQƞ<i�e�7EZ_U���&#ܒIDO��f�J	�.R��m��ӣ�xh��O��h�����E��w#LDt�ƶ�%�k�䅇����;{Q-�ӡ;�L=��2Q�ͺi�������Ӵ/Ř��ã�o�b���}��/�}�xt':p0�
pFFMe-�4o4����R?f�.0��L���1��4c$�N(�O4��"���*}��V�R�S�*x��(�W��(�F"���PϓM����5KS��`Y�-
\���h{����$"�:��u�ݓF�%��	��Qq��4�X��6�ٗ� B[�SĹq��mv�.Z$e"LbMW�S�Z:����Y>=�RӅ�~xQ��f	���a��t��̑2�L*��ݫe��2�b�)������}��m��)�%���Sm#xJ�Qe�O���HhD���웅i�:��if�f�i��GSGn*'%:8~?C�tpF�!��A?�ZYŔi�0�1��h��8��8�Ǎ<d+Y0R�wmu6ښ+O|UX�����a���LK0��O���$�|X���)��&pR�t�4��M�J�S��H�.�L2K[H̗�/�Xg2��&k�쬛c���IҨ�$Q9���H�t��D�Op�]���rQ�t"R@��=9>�];�S��dEkӂp�	��0~8��?c8���0�V2�P2�P�%�1��`�$c ��1�3�����Fh��0f3L$���1�1����X�/�$�0`�!��&4/�c��0`�5��N�e�i�F�yy�x���1�c��Q1�c$d�2�@���<3Ǐ�<i�8g3�iƌќh�0�P�bc4����1�1�k���t�n���֑n�u0��1-��7;rsTw(j�"n���&y|�$9��K�"��_$��n9�1x��o���:q:��͒�Ʌ:J�YlO�,n,�}�<�z�Wqu^[]V��K'{���T8�fO��K_lò����W9��"%�?s����ޣ��������ϻ��{���������{���������}g�<i�3��O1�q'q��wä�K�/�=D(Zif�ȥ�
�tx"z�0�d�>��E�Nm�UF����W�aʌ.!=�G�����8�S�@'!�.�J�;qWt���v|����~�k/�[�kc��ΟZZ��%K�uղ�c�ۦM���.5]��8aDO����0(�����p��ZHZ�JOaf�xf���O�8Ì���2R�	Ieβ�d%b��~�Ub''Gf�$�m�#��)Y�ɺ�FW���-�~��O:�����K$�I��Za���j�[��%F��6�Dm�6�GL�mwrZ^�S�i!�ZGȏ3$u\�1QQ��駂y՟��4�A�?m/�W��j�]|��"�a��i��~�x����8��<x��p~�~S�,q�4d�Y����Cm���9-�>ܿ��f�k��&���[T�f[l����%��Bj��2xpoM�*�mf�S���9k�v[���\|� |!Un&&�N61rDJ�L��(�f��_����,3t�8�OH�$�-��6�`�ܧϩ���d�yO��m�Z�}�FQ�\��b�H�O�e��U����S�RW��meZ">��<�-�~}5��4�B���]�\L��\w��͠�Ç0�<9/�(��~v���'����]L6�-�ۮ:�3ƞ,c$�N(�O4�����=�Ub%����y���o�u�饞�SA0M:7yN����3+���v!��?}�{����+�F�w{{�G_FF������+�l�f��Ѳ\s�RF\b5Ow˽VN�*3)�Č��vҼ_!�âd�0���"`��7���0јX�q��g�<X�IĜQƞ<i�G>�\�sq�Ub!����Ȧ�I��;'rQ:�S�S�ru8N���#�߬�q�K�jb2"�)DٙM�:0�n��i�rh��IЌ*v�a�$�ᆛ�s�j�4�B�������i����dƿI��NSOR-��8ӏ:����'q��?�|}�$�T����ΕV"~;)���E���ߟa>v��qyl~a�s�ԒN�[�6���ͺ�c4��;�r>s��e����em�W��ah�%�~Oo�3-q̟�A��c�����Ѻ�u_//SLS����8x�ĭ���t'!�L��p_wƗ�q�0Î�3ƞ,c$d�Qƞ<i�\|��Pʹ����� $�UdI�/1i)
w�jj�vوF]f���t|:\�
�+�H��ŏkQ�-
ԭ-��/?�h����^���S�-������3n�U��8���e�����Yp��nWS1��v�l��j�Ϡ �ўf��(�ג��	S���mO�S��ϑ�aÿ"=.�K��qj�[O�b��7��x�E�n��pM	�b�P����{���m��H���T�Oο`�׈��y��U��s	�FQ�����-O��	M�׵��K�%�:p��&C�J#9���b�$_q��Y%�h����u�a�\|�Ϟ�ZD�Il�$�Ӹ~�C`}�ѡ�gbB��aHz~���V����])���Ư<�{��N��"`�)�T��-�))��u.�Li�6�>��Ԋ�o&�d��,N��5m��*�&�wvm1-�pt���r	��;B�M�>��c��>,���J�����&)��Ϛ~m��y�]y���2FI�i�ƖgA3�/�W�V"NC��Ө}�}�����F�����?e���i:���UJ}��2딳hגmi_F�3y���6��؛�i�C��O�JxnV�Y�C��⧄�����	�����h�ؽ�=k[;0��D����*����e�6�hu�%��oͿS�n8Ӯ>~y��]y��:2FI�h�3���Ңe$��, �!D���EKj�����z�D}����][�ۑ��K�%JS6�iU�jۉ	��&K�y�y����w��SJ!��3x���t&z��dL������	ѓCf��p�i������Mw{�bh��ɥ9�``��2oB�|��wJ!H����V�<㎸�\i�,e��e�F2 `��E�1�h�Y)&`�h�,c8e�K&���3Fa��Q���3F3I#�A$1�c8��d1�3F`�:��:u�'�i�ǞDxb<@�1�1�c�8d���1d��Jbc0e�ђ��Ǐ<3�8�4�@��3Fq�VH�!�҆2�`�3�e�]��ӭ#���tӬ#���$d���j�TLD�Y���Aw���nwo6"F��v���-��3>� b�[#B�q�#����L]o ��ګ�N���I��}#'R2e�S}c#���r�%(����{��c���a����'��Ak� �y�7V�X�Ō*��먲̌yjjK$3#y�~�٪Y#onf(&�[+[o��jPR�̆;-Ȩ�&Ly����b�k��k�1h�r�S;��������}o�z���ʈ�F��ɞ�2nU����fU/-�2�D����Wj})�=�,���ڟ&\����s�L�X��kߌ�p��c�c����&�D>��O4C� �ٜ�J��Ʋ������Z�Ƈ �`b���.������ϊ��R�۵�͸5���3��3쿙��Ktj]\��5C���y�Xψ;�Ed���'hcf;L\ɉ�{���ţ��p� ���F�mڤ2�0L"�N����몕1+*��D�+�
�EMku�p�	��ˉD�;+�RiO����v��Tn��^���-p�$u�i�^���7[a�Vk+e�[���7h���6���T%��G����������QԼZ�ȞX��L�R�}���Z�QakJ��<���=_{����d)��jn#�T
ff6�ЙY�%mvK0Η$���w��9����cF<�c�M["������wws�o����{޿=���k���{�ǻ������{��=���o���0��<x���Oxd���8ў4��~��b"�ړ��(�������5�+..�ɮ��޵�˸b+m`3IH�1���C���c(lhX��홆l܌�5%Ha�v���~ߠ �M�<K�4�J�)���s���DN�O?+�}(�{�a�CR���_�q��rC�D�賿��#c(�}>�����������ʾ�t��R�C��N�;�����χ��G3Y��N�0�g�S�������`��5s�7n�����fV2�?G�y�A(�,(�}Ƕ�(�~?~8��g��g�<Y�2N(�Oǧfv~Hc$�nB�=�gj�"Sm5�u���G�}3_[.<���	��@��NۣU&añ>�9,=�y
{׹na�"����ӭR�}�Ů͗#U��
���e�'��~s�)痉א�5[���|�>a��ԝO�]:+0�|�ȥ�++���o��q����:�Ϟi�2N(�Fa�cc��?R*e{I*��y����M����W�1�[E��>�]�b�wv�z�:���Z���-��Z������� ��`�E�A�d���9S�+���I��_o�HB�[ޯ��i7O?-�6�me�W�m��KFq�g�V�|�vIt�ѤC��W?4��JzU���<��<p�x�Ş#$�4f7���]�͟�UX��dӳ��!�����<=�Qrt'~�_1�u��+��6�˲�L���}
i�ɟ�2ѿ�w-||�:0�)�L�7^�tv'駧K1�K|8w2O�CO�1��W*�Z"#��Gj���]��?>��?+���]��4�lJn��-6�Fq����Oxd���,јx��|��6Z�K3"�C��%��S˃��p���qZZ�nY������c��x"�-0Z�6�%���UM��ؓVB����f�%���(V�0}˜ �!򸈶�GōF1���������[�w;���=��i��S��D�i�*��R�*!�"��i�"d�G!�v&�&G�!�ah�9�%8��.��>[��u���.ߴ��R}�\��,FU̹h�U��{:<�)��0������$y��D��m��q�uלy��a�q�ζ�Er�?j��d��]4�&	��ޢ�SN#mUi�R���+-a�z�i�>#��(�q��">�?Q"�E�*u��[hbݰ�Y�e �ד��K�ge�8H|���'��V.fk>����1?L�P��Hd2j:{'�-���p����Æ1���x��$d�qf��Ǔ?Q*z��M�K�o��rv{�K�a�����4�;t�U�=k��؝��4��'9<�rtɆ�׺������,7J�.<{dƱ�`�dl����!��xz{շ��.��S�;��Ð�v��dN��5��z�á�L>2(�ɢx�S���z-�:��x\ۈ�1�<��m�O�o6��ߍ8��g�<Q�2N8�Fa�d�NL�i�I�w)��U��qc�Y��-�/��x~�õӜ(���=o�Vh�3jhT�Q.!�a�9�0L0��/������vx'���9x8h�w)�_/!�Od�	L�1��(�K[��bt'Ћ�T�:�)�F%8�Ԭ6��L8�%Wθ�z�r)�\m�̼��^x�3�(��'Y�0���C��4Ό`���[+�޾o���P;�3;F�l�{z�ڴ���f��3oW�Z�\��+�Dй!)q-!����v�I�T��7g@�, ��<�ai~�Cy�����TMo���VԴ�0��a!5l��>�=CҚt0�n�u_܆A¼������#h����Un��8nI��y��"$q��e��BpM���^�ܸ��پC����D�y��gS��������h3CJfFŖ\ܻ���F�F�n��:8w�Ǔ�D�N唲�8[
%}G�L4��4���g�<Q�2O���NN^&FLqUb#�ߗF`��7�\SVzj	��u�d�*$rO��뵊�G+vN$�}�>l�8�Wϩ���}�r�G��kwoI�a���BS�����К'�{}n'�|/�[������+�S0����-8{��X�K��y<�4�O�����`�x'g^<<����F�%5i�O<�뎸�3D`�C(GH��"��Q#8e�!�1�3�`�#8њN��3Fh�/D�e1�r��qc d2	 `�bdg1���1�h�Â�C�GN�d��Dh��ǫ�x�2F1�c8g�$`�!���`�����<x�ǆq�Oi�!�3�4f��L��I#�3
�4��gYc�B��CH�!����V��2����>��D�_�4���|�{��C����|ٹ��<�z�٧�,!�*}}q;��wd��7��t D)�>��6�b�3YyMa�E�Ԑ���q����בL��9�+�vv�h�؜�4��l�!��d�}�qy��ȼqe�xKק�1&.+�;�6ss�弻����z�gy�M������7dCژw���⮖��Qw	��WWEb%4[��o/\_F7.��[ur��I8�׽��_v.VƖ��w���{����{��������{��������{����{wwww���x�ǎ<3ǆ1�x�G��8ӎ�����$��it�'ۯ�����K���}v�e�k��*�ӂ{b	ّ/G�M0Og�>���kX��k�R�\�)f�M4�����\0D ���N�1q�Nó�:�+�l�����.�T�0�6��oǧe]�i����U�n���y�e�^q�y�]|�̼���8�o1��s=�b'�<�ǷR��Ұ{:�GS�==T��"aǅi�tU�*��@�f�(�� ��\BQ�p�7-_a�`t�<���M`���� G��KYC�Zf��o�f��UDx�]Nɇ�r\%��>qN&�vV���ׇ/���[�+N"�b��|��q֟8�κ駏x�#$�8f6�$�J4F��Ծ���%uuJ��zoK~��]�CFdz��Ȫ$�X(���<��[��%�P)28�CD�k��n��Ҟ��b�Լ�[]���"} D��c������|ni^�
�˼�f8��[a���<N��}�lb�D~�Z�S�2�0w�[kJ�8���0�~�?z�� Òh6�;C2��BS�zy�p����XF)h�t{R`eh�wu��I�M��Ω�sv�ء��n��ŷ1�E�'E <O�CD��=QΦ����.SU_6�O:���<p�xc��x�#$�8f<�Xl��v�d��{���+�<`t�w�z�Ub!�,}��t�/�T�Gq#H�T�#�C�Z��d=,7�{�)�B}L��q8���#4�֗�R2�M����s�ͻ����sAS�`�<?a��ꩿ=��U����n������~)؝�Լ�Os��R�j�M��N�a�y�^y�]|�̼���8�o3��Z�N�I$��V���N���c������+4��a��|<�&\��Ύ��x};D�����y��,��vI~�(�ݑKc��߬��iO���V���!U��ԟ��-Ƴ�؜�)�vp�H�6�.]��t��}Uȓ2�e�|���HbQC=��4Q_I$�p����1�x�G�2N8��a�C�=h�K+(�UX��΄����â�8A��2�$G�͂g.b �$5ҽ�ҕ�n4�WkfڻZ������7�r�{䍶�`��È�0Lg��a��iD���xk7W���F�V�;K����>�W�m�-���-��~�RG�qL�ˑa��尝	�̃�#�gk4?8�]q�y�]q��2��<��p�<w�rҾK��*�SQ?L�)�q�5�k]�"��'��}Yw��n4=o�Z2Kf��L�&y��ҍ�-�=�`����BX`�%�[]Xl���>��
j	�F����*�COM�0��iஇ��gf~tcП\��Y6/�����J��{R;/5/s�Q��u��+�m�+�;�R�9mO+O��?�r{�1SgT����r�ʋP�}��;���-s2�ǰ�N���� z1:�R�	�V[*��Z�C)f������F.���M:�İ=���䬲���u�u�_:��y�qŜ3*�����I^I$�����*�l�Lਫ�N�<�t!�O�Nu�4ľ����;;2A�8�>�$Fθ�kv�>�zu�Ũ�	i�2��sh�G�ւ�iu��H�`�������_>�3���ē,�[�����˒d�|�����W�s�"U׻��if�1�����x�'�8��?��F����8�+�4�A`�e{�V���m-����
P�,���Z7�̆��\DU-�ܗ��E��Jw8a��N�����ӵNC���Ci=}�.9�������)�w�ϫw=�
\N��Mf	�[�QӰ>m�O���ܮ�h�}�>�e3��u��}WNܝ�p�=�?~{�t����cr�`��v��q2�-<�:�|��<�0�8�m�%��^>��,!e�D�
�$D Ax),%8P�1��y�'����r�6�KaD�̭�Jo�~�x�GE�R�	=���ʶ���͹i��e�n�nd0��7����'I�p�2�i�Q��q2Gt|��X��u���.R��G�'�0��|��gp?t���g�a;���a�/ޙ����b�[�4�O�n��/?y�տc��iK+�VԪ�4lٳp��o~�o��՝�y�5���x��rrN��1����C�y�M�a�':29�"�k7s���MȈ�"E��-��""�E��;��"4h��DX�E��DE��",D�l��h���&�4["h��4M�!AdH�-�Y,�h�dD[F����������Y,��"�Dkh�dH�dDY���DH�",�!d-""��!d(��dH�h��(�"Ȉ&B�"�4Y�h�։�K$��D��!&��ZM,I����$K$KI���d�di4��m"X�Ki4�H�$�d��M,Kh�m��m$�&�$Ki�2%��[$KibBL�4��-�id�Y&�L�bM,�K$��X�L�ĉm&�$I-�&X��im"[I�iL�Ii�Id�d���K$��2D�I�I-��D�$�I��KI,�BId��ۍ$�D�,�I2�%�H��K$���idY"YL��-$�dY$�"�id�X�Ki&YI$��&�%��$�-��ĉm$�Ki%��d�-�L�H�Id��	m2�Id�i	M-���	d�d�d�Im$�Ki%��4��&[I,�Y"Y&�H�i%���$��Ĵɥ�%�I-�H��4��m,��K�D�$K$H�H�$K&D��D�D�X��L�i4�D�[H�I�IiK!dF �T�p� �F$��$��m$�M,�,�iɓKHK$%����Ki�%��[K$��[%�&Y&�I��%�l�K&M,��I���[Kd�2KĚX��I��	���X�H�im"Y2%��Y&��im"X��bD�Ib[Ki4r�q�%�KKHK$&[HKd���HKi�e���L�%�	m!,L�[%����Ki2D���im,�K$K$�-���BM-�Kd�e��b[EI-6���3I���k#I��m�ۍD�Y3H�ɴ�&i�H�֛h�����m���md�D�Z�H�ɟ�md�&��D@`�bi�D���s��Y!-,�(q�D�"E�"E��7"-D�!h�ˁȋ"E�E�k"Y��6��"�Z,E�4p�E�H��dM�\��Y�""h�dM�q3��dH��h�$[r��DYD""Ȑ��8ȑdMD"Ȉ��\�9C��E���DE�Y��6�-�"Ȉ�",���h�dH����E�p��$H��D�"#Z",�D�h�h�i�""Ȉ�&�"h�D�dD[D�"E�#Z,��4[D�m#X�E�D[D�"E�M�,D�"E��������,��mE�[DѤYE�"Ț,���$Z$Y�m�dH,��"E��4Y	-�Gn3�#[E��b&�h�YF���"dY-�#YD""�$D[D�dhE����",��F�,���,�DD�k2DE�H�dDH���dME��b$YE�i�4H�",��#DY&D�h��dH�DE�!mhH�D�"E�dY,��"��dD[D��QbDE�[B��hD[DF�5#Q˧�h�M""E��DD"!dDY!h��dHY5��h�B$Z$iDE�HYDF�dDY	�!h�D��"� �H[D�h�b-�Y-�h�,�E�#X�E�H�D�h���qύ��"Ȉ�&�""����Ȉ�"-#H���m-�"Ȉ��h����"4Y"Ȉ�&�"ȑb5�H���DE�[E���mE�D[D�b-�h��m"�"-��Yh���mE����"ȑdH�"-#-��DE�m5�"�,�BE�--,��D��$Z",��E�k"h�&�"dM"h��mBȑ���"E�h�dDZ2ȑmD��24�|m�h�b$Y-�H�&�D�"E�de�!h�h��$Z4�h��H�-Ѭ���"�"ȑ����"�"�dZ4�"E�E�E�h",���"E�����D�DE�h���4�""ȑh��$M"Ȑ�D,����"-�h�E��-����m���p��x���y3���f�w�?{�>a�)[0��Ͳ��K7�ǫ/?���wu��ݽ~w�{s�����9G����p�=?ǯy�q����n�៣y;�������{�螏_Lp������_�:vy�/.|���r�9�s����w�v�2�?��ܶt<��������׃���lٿݞ�����7�����.M��c�f`�Ȏ��X͛7���kpo��ۛ��m����'��c���[,�˖ߖg�ng�&�'����֝�>�g����͛4{M��o���>dIY��v�ro^���[������Y�r�|3��鳌�?>v~�9��q��׳�]��ϳ=x�ǫ�{ym�9Κܩh��;o����8�{���qÜ��6fsL3f�pz�f�ˍ����09Xf9Y�l�٢��U�VCG��X3�����ә�7��9�7��7F�k�f�n"Fe1��l�C6�lm���e���9�����i�շv�ξf�~�ȷ˻v{�鷆��ާl9�8p��t}��ط��_;��{>M�'͛6nY�n;���~M������ݿCn������??��n���;�f������߉�|���?��}���C-�{̞^��o��8��ӿ!���������f͛�-�F����6�?a�����{���߰��{�3��m�����I���6l���7�̶����?6���.\�|���y~V�zۦ�ý�����.���c�m���f�ڊ�~&
��v�$��Ob�HB]������7-��~.��Gf�:7&����g᷼�q�c��1�e��&�4���L���!�E�����m�6n6:���%_����,��m�݌ٳ{N_;�oԛh�y�ކ�W�s�Ǹ�����_�7!��z�Y3���g�˂�7ϟ��o��������ۏ�r��8o��S~������f͛7��<�����	����Ӷ��6l���:�s�?�y�m�=y�<�[��&�~F��W؜����M;6ZI�}=}���D�V��1ͯS|w#�Ύ_N9�ϛ�x6�}Y�l�G{����3��uξ,�ܝ͹w�{ή�͛4�r�m��ˮ�p��q����3y��8nA��m|�ѻ��{v����vL{�;us7F�ӽG��ߓ;������e�������f�#��3����i����v�M��f`އ�s���~/�u|�zݜ���������|�Z}y��ܲ4m��c�������"�(Hz�H��