BZh91AY&SY�+'�ߔxyg����ߺ����  aM>    �                =�   4    �    J
    z� �  +@ m8x�O��$�  >�  @� �Yn�8����l����۝�|Zt��v���qG#� 
]����'��d:���݀]�@��3N@ hC@{���x   3 �����E�˳��� w)�;���^���7H��2Ywdt�  4Ǯs<1-��e��z�I
�&���]b��0��r��[�e��]�  �� i=]r�örk�;;����kv6�dd�˝��8�Ssu�휪����94qs�1�-�T�c�N�r�`s�Ui��tn���N� u�    ـ jn�..�N�W'.��t�v��4�kkݕ"Q�����WU�9�ZP+zWsz�Wg;G8�e��;��[�.�.�:�2n��˧�bD�    l��Y��Ѯ���s�U��n 8��m�YwX�t�NN�p��nN�ne@)F;��;��yEy[3M3y��;�C�SoC�����7[��@                       +� 	@a*z��(0&����444�&CM4OЈ�T����4�14dbF� 4�m��RoD� � � 2  	4�BT� `��@ !�4�@����  LF�����=�z���6�UO�MʥT�20 ��A���I����Z����3efY���=���[��m�:99<Xl�vfFe�Ï�O��6ãc���a�c���||�l͇��vm�\�O��?��ߟ×_�p�}=�nk�O
����6fÍ�ǡ��s�\8�S�|�l͇b��n�w�򪪣?|8���8߯�|K��~o�_G������F��<1��i�-�e�d�!�.�c�1�3�&�Όe��e�1�c̔�1�z�c(c&`�1�1X�;T1��c��2X�h��H�0mi�i�b ��8LgF3M��C&1�am!!�c&1�e�c#�1�X�	�gFh��3���@�1�������dLc$��38�3J ��C$C�A�1�gX�0(��`�1���gG�B���1�@Δ>2�3F3K�cC,cʱG�u�c(f�ьgX�2�`��!�e2�1��H��V!���1�u�1��DA�C���c;�,F0c0�QIC$�!�c�:@��2���gG�3gY#�e�ìc4��<��3c4���ɱ��P�,bd�e��|�K ec-�P�a��cd��@�2�1�c�Hь�1�����4b e�ǫFYgM;I�cm!�4r��H��`Έc:�1�3D�!�c�4e1���%�1�1�#(c%���,Lf�1��Ld
e�c�uiC$c,���`�Xǂ�2X�2��)�1��0���Lc�cH�X�w���gMic���I�ȱ�c���e2�1c |��"#��"";i��c'J4|��32^d��cc�K#�c4c��1�f񌁌Lc�^&2�CLe�e��1�c+��eH�+�3Mf�@�1�������P�Y,c0��c���S�3�4�1����#:K�tf���3�cC��!�1���,��@�f1���1���1+0e����2F2a1�c|f�c)�c:2��Ό�1�1��c�o�$cl�(� c�+��c$�=�3=C(c�2�`�.`��c��1�]��]4����� �Č�&�M*
�"��+���Lz������<Z1��P�H�c�Y��c%$�1�fJ��c$z�g�1��PP�3�����1�$��d�ma�*J��3���F1���$�1�ь���gFX�2RGM�I�c:1B`�H�=X1�aC��1����� cꁌc,|c4`��dc�3F!�� eacI���11c�1�Iq�)�c��a�*c�a���ǩ��C�*�c6���z�|(��D�$!�b'���=HGL�&6�4֨�D>�C�"�e�C.֚aM!�fjc$e�����`�1d�U�H5D�A	1�I�GN�eZb1�+���VX�;]ǩ�H�1�x��$���;L��� |cS��H�u �1E'Φa�ґ�0�܆���.1�2KgF2�e�2��h��ddad�2@��0cj�Ί��tv�2FH�f���њ3��e��T2�F�$f��CC��,p�c4Ĭ���Ld����(�����<Lf�	�aC��εa�1���f�>t`��c�i1�c0C�@�6�S�_c�)�c���¡�v��hҲ:Lc$z�,pa��:Vq���X�2�2h�tC�&1�ccŉ���1��L�1�1�f�b�!�1�c�Cɔ�%dgZ�1�e�����1���2�2�QC)�ct���H�*Lc�c��c$d��I����UEUW*��y5�qǌMj!����4��P�1�c�c0x��PƓ�1�ȑ1�t��щ�1�c��H�8Lc�Ld�c�c�t|��c��c��c&13j�,c��1�i`�1������6��1���1���1�c$c&2��3i�H�>��2�0��d��c:h�i#�Z@�1�c4�K4t��ũ�H�f�c5�"D+�1����F2!1�c�#H�E&1�e��4��dbc$c2��c#S"c3���Ft�d�`�e�Ae����aM!���2D32 d��؆1�J2�c�C$c:c,dѦFe�LF��ap29c(�L�-1�cJN����(e�e�0������c)����3M0����1�c��2F2��0c�1��LcΗ�Lc�wS#(|��1�gRf�e�Lc,���,�]c+F����I���hfڒ ��Aq"\���#����gp�!�wH��ΚS(�XΚ�f�QY�H� cS���J$���1�c$|��d�c�b���1ڱ��>a4�@��i#���:<Oi�3Mɱ�t��L ���h�0dh�,��,��D�t��#�#�q��X���# �iC:�H$�Is���!��6��E�,c:=\c0�4�P�gz�F;L�I]:t-��H�����H��I�ѝ�$1� ����d3���1���1�>3���L�x�҆iGK��h��2�Ƭ��$}Le�֌�J+�c�i�:�$c�Όc��1�b�I�1������鰙�>bc$d���N��(c�"�1�)���e��D@�1��$iq�c�m0c(�X�1�����H�*L��d��K4c,d�c$�3!1�iC��`���1��c�CѵB c�f���K�@�S0c gN>1���;L��td����3Hc,��gF1��`�!�����e�`�@�wU��1�4eaьz!�0c�@�:1����1�Ee1�K,cΗ�c�Lb�,dҁ�f��- fd�1��,c��c e��`�>tc3�c+T��c%�e�`�(�1�gF"��!�1�f1�2;CΌ�G�:H�QLcΐ��2FQ��
�Fe��酒�331 L�dJc!�c4�2�$�2H
c�1��J4�t��a&��YE��v�f��aGDQ`Ό���4�hb4�0����C-���霡�!r1�����o�C;�3p��:T:�w�eWJ�'FQgYӣ.�k5�B��$�#K�AVF��M�L�@�Mq�JZa���� �K(�28��!��
a#(�'L�Y��(��Hc$}L���:4��1�c$�����e3��h͵��v� R18I�R:tL����M1�i���,d��21��h��f>JfH��2D>h�t��ȓtf�tv!����3���u2� V��>$��;R26��L,���X���Z�,cR�$��ń���ӧK���(c��350�G�2�8Lc�$�1�C(c(z���	C��Cf�4c&��2��3J;)�1��LeH��2�e�F���1���5�a!�p�ьr��!�#��1���֐P̈́� |�cC%-ԙ�1�L �!��Lc:[\C�-�d�����X��cE�3A�e��eb��1�P+�ũ�ec6WF2F3�fc�1�1���0f��i�&�L����)�k�~�g�m��ſ#������h'�M�i�">����3ɜ}�46hw�ٓ��!����=3�Ws���2i�=����=���^��N����_)�QBf˿�v<���~����|�]0{��,�d�M�d�N������w����z}�O��IZv�$���%�!�qf��N��M��a�p����}4����k<��aI�$܇��Q���ۉ똗��3��3L�?��5l��?n�~�b���g#]���WYrdp���y~�9޿B��5_�՗={�%�3�'�����Ùn��/�읂�d'�X/�t��9�����wu����uwO�v�G�E��is�ys�/[������d�ޖ�K5\�l��1U5�����4�'ztx�\�p����O�����n{<��6���Y�+��џzOr3�R���)��kΫ�
��ž�q���qwh�P1w��������c�ʚQ�n{} ù��H�������>�.fe:`�1\�(H��d�i�{�#�w%�Iܓ$3d�I,��m������9�r`d�L�>͆}�o�9�֓���������ߧe�}������ӽ�h�H{������ϕ��`5Xҹ�r���)�%��{���d"�{�7Gc=hx�eٹ�3�5?�w���S-�7�ܗ:hwv$����w�!��w;�V��4�O�32F��0/���I&rI�L�;	�$�tg�"�QI�3��d�f�<X���8>��*�G�j��R��L�]M�*��o�{�8w6̙ݛ�ٞ�'�_-���f��>wf�I�m�w㡗KG�Q��u{}/��0�4	_��Co� m����U�~�Y������֪}��  ;;(�$ު}�x���{����gv2��Ǹ�r͘5{s{82osI��s��ͻ�<su�L!��r�w�x��^�$秇�7y�VN5x[�0[Wz?�w�u�;.T�����;��I��%gs�\��� 	@�����_�����(�
���R���T��fOL�3�i�L�ܹ��P8�>6{��.�2��Ľ4��F�^��?�}��Wn�O��/o��f����n7�̰D�6������Ȟ�>������y����v`�d�fO��j@��Cr=̤��� ~��/�������?�������5�d�fx� �G��bZ0�����I��pZO�/v�;nfe�1po*�j�3���{����n���Z�>���_��h7{��t���8֯��{�;aᔾ%xN�=�}���}����l��U�~m,-��.��x���?ß����d`Msy[�d�L��t���K��n���n滌�u�Nz���>�:z,��M��f���ެ���s&�;s������{ߗ�ˎ��J�s�006\�(vN;�s6���<jÙ8�ｰ�:�:{�^��s�I�@<��f�U�d�}��)�M��$O�ğ̴�To�ˬ{�ܗ�߀�*���`I{(�<n.4�j԰������3;��7���?ݙ���ˮ-�+�<�fJ�B�Y��;��;���v;n��[�����C�ܤ�{3?�;9�x����O��|`|tx����'��34z~3V�,9;r����gO�36jZр�:_�[|qs��ӛ��������߾�9k�dӟs&��ZrH��G��9�~Y�/��G��yuWgk�<�ڤ�"��.��O��V�y�P�*!�v
q�O?bC��^_����#�}�̻�mĘ�eu��e�z���������n�{zj��f��ܖTe4ɠ$�:��Y�Ou\0���]'p��S3"����L��J���G���*����G3���L�}���~��l=�Q��M��o4�����:�������$�~�0�u6����W1�t���ǂ���*0��ogw����L�TX��y�|��F�c�f�c�gf@�����֞�蝳cۢ�j�e�ߧO������ɲ�K��g�?K���\��%���d&�r���6���-	G�ܰΕi���骽�����O����s��җ|�vd��1c�7(o�ŧ;V1�y���;;h�al��ћޟ���^�ߟڸ��s��vi��������1�I�73ssƞ݉h�l�J��S����`w7� ���g����:.d~={ ��3���I$f�@�Ζf|}Y��.^���_��:w,�l�4.��~������i�>?T�T�������M	4�Gw3���v�۝T����l�.�u=ӷ�V�ts@r�єή���}~w_yϞ����ޫ�����܆g��*�\�}}�d	�ۛS�3��f%���Ʌ�$結)�L�����r]�>.�1��g��I�}��K�҂ٖ���#�Zw��VY%[:�vfó��y��u:��6m臇9 ��\u�3�Ͻ=��,\��L�����nc���@�9��Ӷ�3�N�z��{�_6U�jF��w>���׺?G^xs�};���&��L]������q>r]��:��{)}�d̶v�nKwG0�V�����i�ȳ5�������͓{��N�fzy�߿��z���r<�d�|o�n�خ��5��d�N�)2㵇b�E�����n������f�[�V�V��Qk��w��{ڟ����ņ:�g�5�N��V�؅�by����������8z͑��w��}��2�%�f��z��ڧ�9��|�>r�t ��h��6���@"{n��ٕ�}aެ՛�Ŷ�0'q]���:z��߳��������w��&I���ek�x�l�%�L+�x9�t��G���sC�������������H��w~�*�O�ӊ���ٛU�Un��.%uO��-���,w=��ӳ[�ޜ�ƭ��ߕ��^���yކ�L;i�$;���t�S��\��K�ѝ�������	�)�gew׹e�+22��vE\��)u,�u�X}�B�����Zl3$�|w�Y�Y�O{%��%M��%�G х�I��__�qs���P;ޟ��Y0�~�k�ٻ�.G<�>���wl����� >��%�]����u�{}�]D�qN8��!�f$���גs��wr}܆w���}�vW{S�oI��zN����K��A�e�ps�\��1w�3�.w��dǝ�}.>�l��������0�2fL�����vwH�9�l�0z�K�0;o�Κ��~��/�`����c^��z��!�1L�C�8G�==�N���������}��B���RY�70}}.x�vw����{������<��#�7�ݶ4fjͯ�gs�S;��&�y���w�{K���$���w���H9�>/��gK5]����8;~�'SY��ػ�]w�C~&d��臘-���'�_�q����b���/�f3���ng۲w2^l����?E��V�{�gN��`gcY���7I��M����d����hֱ<�7�0�2��G�[v]���^��>�8[�<}���ޏs �f?u�9-�ٖ����z'�g�|�7���L]�����e�>�tȞ5����x�nYA�YBj�;��:��Y������:O)�c�y��s>�;�����}����\1�d�r;�Ք���nwG"�wҘf1x�Oh�_|g�w����I7]�ϳ�N��#��naY���S�M����:��g{U�K���a���.�~��G1ֲ�?x����zf�MP��<�]��]ح����s⛓��e�w]um��v����	��|x�E��])�RYd_�<���Ե�B�JO]�y;����}y��v�ә'�'�=��X`e��#����MٙV���w�nI���Ӣ�1��{��@��_:b�`���Ɂ�-��d=�[�ܘ.��{N{��R�6o��sJ5��ܚ���L0ˏ)�v��'@vgv�nN�>���O�7�	��՗��K��{����_��s��`ڛO��}ɩ��&Ƴ���m��+�� mmt�d����y�;���r�\�.�|/?.��VOc�y���rܟ���K�&�4���.��\Z�m����+���&�AT����,pƎD唕��ek��9l�����YL*Qd-�C��@��_�ȅ*�0vH���ڦQH�+g�,�`�V^@TB�#VKa#����J7�[��EJ�\���Fڲ8�A�lt��!�vG�,�j�XԌqIULuNTE`ZV����Pv�"jW�
q�T�Ij��ȝe|a["nB��*�( ��E$�P�#����US� �(�v�c�m���K,��%�Ej�J:�m:�
MeiS�wJ�M�\ �mE��Z�r�d�c`�%�q�N�B��rڜ�i�J%"�UI�p�W*�Z%�&DQP�4�V*IZ�� �R*5�$�
6X���[%nB��(�����j��8EhQ��W�ՑG!�r�tD����v�����+�,�U�8�ҋ��$V�ȘVR弳q؛��s�2.�J*�D�	;�0qA��`�eZUQZ��X*�$�JF�6�(��@���n"+(������!\��8#�u�܊*�rRGX7%m[kn�	[�N)c>���:��؇_�d�5+|QZ7KD��_���
�U6������� u����j�j2��-"�UP��
��(�*o��*�l����9�$��Sxܐ!S��d�C��j hn�Zr+����"�r'j+
�J�A,"T�̬M���q��Q��e|��qX�K�ʉ�`B�p�دU�Qj �-q�j!W%#�u��u� u@iجu1W�� ��aD�(��iS��~ګNƣ2�|���6�P����A;(�v�e���2���k-�B�Z�	F�F��&��Kd�4���$�^;i+���9m�Q��8�,bjF��N^ +V � �Eb,I��"����Bm�_-d�%���#V"PR�Q�Ӆj"��*��NX�G,)���4N4�V�p��)EGA7@�b(!W ��
�-*�$>>9"�h�:��re����n�R�Dq�k�6�W �E
��S8ڹ�|���!���(W���&B�kc��V.~ǋ��/o�,�x���/�NBP�q�e�����k��s�E�z�J�૨g�?E�>4g^�9���U��1���.����&pǄ�5?�׆j�O4�H����rJ!�⥑�EA�ۍ ���'��֥U�$�ۤ|���Uثm'NB�Q&�K�9!#e-��j�x�����:&یn.�T�^7`���Go���4�%mȣ�������T��AGj!X�n�h�EJU>�m���v�(R�� ��<�^X��TZ�N:ղ���TU(UȜuG��1�*6�iB�6� 
��m���ɺ�F��,�`j!�wCTI&4JP�ڐ�L���n�#��m�F¡@�QZ�ֲ�f�C�j��
�Ʋ�T�� 'T�(�X��Ug/%����D����Q&�,Qb�Xo��{n�(�����g���.\x��ln�����S����<�?��y���>���G����,Sm[j,p��W�qm�M�jֶ`�s������	s���~o��o?1��o��M���[n[m�m6�m��m��m�-�nm��[n�n[m�m���t�m����۶�m��i���m���t�r�m�m�m�UO��m�ݶ��6��m�m�li��oX�m��s��<ٶ�j6gTf��5V6+67ŶmFd�Q�.	�8�����6�֛֛m��m���t�r�m�i��oX�m��m��m����ݶ屶�m�M�۶ܶۦ�}ci6��m��6�m�p�m�m��U�6�m�i��o��o��M���[n[m�n��.%��@VQ�e3Q�ͫ`8	 m�w��n[m�m6�m�m���M�m�n[m�m��ܶ�vۆ�m�m��cm��m��m�cm��l}m�vۖ�D6ۆ�m�m��cm�������ۖ�n�M��z��m��6�m�p�m���ts�R���E��
�Z,"�d��TZт���+"�J��[j�ib�)���XY�ł+X����&Z�`��/�2ʊj���=�����D������>�w�Fv��r{�ޗ�=�k��;����s����눈�8�hDGDD|�����C��a�Ye������"#�z��!���d�gF1�e�M��2K4b�X�1�b�2Ft��`��4��!�C�1�c��(c�Yьc(cm���DDuDDx���=q�b#�1�B#H��i�1���i���ۮ<B"#H����#�t�1�f�F�a�a�1�1�cc!�eC:2�I�x�����#��F"6���"6���mDD|�D}����(U8�o-�V�0�ak�:��Uj"�I	
EO�TY!̭��B��d����b�����dR�4�8�j�Uѳ��l�R��ԥEk���PLu�hە+�����Y�	��9V�dP�Y"�F㼍���,��3"��Օ>2 P�+k#cP���7]i�b���E\��V6�|yb�cq}.\�F���We���b��*�� �t,nծT�`ԍ)�ŭ�a�6�-M�`��d+��Uc��*
7jti�e��X�p�J��BX!7ln2q�"M7*��Q�T+M��t���Z��銬H�'�p�NY\-L�GG)H�mrآ��,r�[�nQ�T���+AEIE�8 �ڀ	�b����-J�V���X�rR���q��b$u���[c��be�T�D�l� h��X(�K R�;lv��4��A*�m	mn�q����#�#��D3��aclCaU��:)�N0M���j������+��O�8�@�Y�\A]��	�^18Զ	�K �)$㼱�9Z���!��o��IU@�������Stm��(��G�ӌj�Kp��i�J��e��K8Z��DqQ:GF(�#cQt�v�,cm�x�dCV������0Q�[9)#X�y[��&(��0�j(�U�u�⊷,�b�H��|Q �H�h�-v��#V+Pe �45j��(J�j�F�P���~�K�5s��#�8QKF�[8�K-��Pj(۔�TN��--���!"�8�eJ�	�Q�/)+�����i��
��HܑIl@ZU�V1WZ�$���V��NH���'K (�+�+��[c�\ԖB�\mA�����֛�n��q�:r2B�B�[+$rXUG(�#i�-�o*-$��X�b�e�Q�&�"�6���\e	��������G-�I1�f'd�����%uڭ����$MWy��;UV��EkɉKN:�Dq�I�-����ݒ)mvDGh�V���NYZ��8�[eR�hDQ�bn�v�Y"�65�્JK\%o��Q�$U��Y#
R�Q�*۲N"+%*C���	g/#Rq��]QDխ�b" ��!�
�%U�4&�����h�
>8X'$m��]$���tl"��m2��$�NUN'hc��Q�5d�:�k�PI�UDԠ�Eo8�������y����Ng9�����{n��I'{�'3��?����m��$��|��s����+�Wu��괎��QDD|e��D�P�ա���G"*%D!TJ�El��7[�R��E�Q��4�DP��(�ө�	�4K)P>6 t�J�Uc�X�$����*��Gl�X�n�A�]���$ڳ-�h�4ڒdN�[��"�E'��@V��8�⃖H�jVNZr0q�T��u�E��RGd���(�U�Vpn�R�Q�U��*�U�@P�B���:�\�VK(�嶤H:�	l�R��jKF�mY�6�D��U�a+�L���NL-c��t ĸ�_g��z"�՛������q�M]��q�;]�"lCj�E�;�s�x(w�)T�Mon[�L��u�y��~xж�j�*X��[6S���YK�l�����.��rӆ��!�=;�7�a!i �%���$X�dE�Ab
�cQ
#��d��Q'J]PċNH�+�	�r0�&���9[��켢h�x��43���?ʭj���" !�SLq�GGP:A)H�N6��ǈ�	��k~�-�:1:R��E�N���B��$��ޝDQ$���4�x�>z��H���DG�����0�BR���]	������)�q�P�M���4�vp���wZ�et�$�z>k%J���$I����f�y�0���"������[v�O�a�ؚ0��3��l7#1ƫ�taGx�v�#�H�b�Ew��3��RM ���[e�ߛ:��y>	���[S	$My�.1󦉣Jz�[S�t\(�J4�L4fX��i�,c4c�d:Q$�">���)��kS\��|t�_6�"�{x��;���#^�!��۽��%Nw�w�(��F��B���l��Q�>Lj*!X�E'<�nN����C���l�4z���/N=����yU4&A>#PII	���Hdp��b�7)��|5�ݍ0JN|����M�%0�ݬ�G1]��-N�2ja�,�1�af�1�FX�h�1�=8PM�0�Bk
���,3��R�d�͆�҂�p�Ssk��ߛ��Zՙ�3ABG8Դp�Q��9��>{�8+EhA0�\TH�#R\�F�qE�%��הS���0�d߂������Xnlz)�p������8֞<V.c3X��1_�x��?��������]������cN�U�0јaf�1�FX�h�1�|�4�����O���4j�q�k*��ƬI���'��=]C��.�}��%���]�沾G$i��L��&�p�t�㪢QF|g�w���3���*� �MѢ�6�Uj�э�����z[X�7%`9��R�Z����� K�o�?O�}����6�X������9��6������_v5��Y2>� �d���6�0�H�[ڵ$�؂b�g��2A8�YJt�h�ѹ�n�t:)��o����zxjO���S�{��}0���-�8h�C��0�4t�p~�zlѸVxra���AOETh�4%8SFB�ii<���G y8c�똬Veed,�|�[d�����w�~O�W�LK�*�#�YJ�mdm�Ut@�U�˫W�af�`�4e�f�c�,�KQEP����_��
�	15ռ�gK�0�c�&�!��S|\6iVzz��۰�C��t`����@�6Y~VJM'���{<�CqsZ.���f�ۥ�PM>KQ`�,p��D5NKS�Χe�ŭ,$��@!F�z�T�9�Ce<&ϥNy$�,������s>0�k�i��Z�-u�����QQu�z��:���ӏm�H�2 	U5��yw-]WQ�ߴ��m_<�816n<��ᚿ6��>�2l�m9���46��mM�l��ɠ�⤏p��C�jH0�s�! �NW��
��]���x.F4��@zs���,;�Ý6zrτ�Fv}��.q)�0�L'p�;�|S�WR���RJ�����RH�j"J�j֪R�U����U"T�Ҩ���,by�5�>���k�J��z��^��y�Y��5C��0�I���S8l,/`��G��c4Sz|���6k�%:S�	�W����j���UQu�z��:��f�0ПLA��y�Z���~�VQ������|4_oF�Sȫ��\�V����E�q�+����&�j�mp�|�𧆄�Rϊ�Hhg�[��ɿx�D9>�"}���� �Q`��a^�٤Ho��fCd�L������ǅ����j��s��w ��\=�[S�i�w�ƥnU��Fl���4.��F�⻕
$�O,��h�a��y�]G�����u�x��4���i����ŇV�ۧzi�j�a��P}itK���P�`�������<�M�]i��&���n�T�s�)#�i�=��%�Na��&����˲��!j��˗9$嶧�2AQa�D7�m&ds��X�)�9E½uDŢl��$C��"���vBW�dv25���u69j(��r�Ѻ�Ɯ��Dl��X��� H
�!����Q^��yuk��'w�nMo�v͏��!�� ẍ�̈�[["��)�fW;�s�ٹ[!"`�����<�AD���]:)vf"H0������|.�h��L�6e�M>������y���;D�kfᤡBM		jh�Ѩw;��\˯����o�ܼ3l$���&�z'N��ِCB|P�U�W-�14jb]���pJ�h������Y��{��ѹU
	.1GL�*��TqP��[T9I���ϙ���n�ss�|�kʹ�lxɭy�	���-���B��*.��L�::Xh�<i�ag�1��FX�h�4�N���$�X@�RIs�Q����KN� �ޙtD�ݯ��\��p���C����S�]@�$צG��sC..�I��WS��Ss�Ixa����d���%���M+�ȅJ&�Z��;�5>0��dE���3_K��NQ��K�2
q6$Sl�T�����rЂ�	RQ&����m�Bq���Nn�bE��>>�P+�m򪖭[�F�b��<�xjpv=����.͟uxCǦM�Sݮ�GIx��x�l����m���L2oC�����?�ើg��V~VW��j�w�Y_+u�#��<u^i��~c����*�����)��VUq��j�ε�Y��|�٪��f��X�ʬ�eVmU����_2��UeVTec*��*�jƚ���F���ɭu�k�Y�Do��VUV�U��xµ�g�ΫX��j5�U�kLV���5ZiYZ�e֫8��V���Vu�5�V���+U�\V���F�o�g|��Ϋ=Un�\eVUeq�k�W���Uem�kef��i��Vb���[mw��ʬ�<h�c�ҵ��U�5Z��:֕�j�ekj�׎��Tתʹ�ʬ���ek�2��q�����VV��7��<�#q�FG�[��Ui�sU������~g�~c����������V�ֵ֕�4�V��h��tx:�υ��E���?-j�>VV�֫*3��5Z�V��b�[�?�����<����0���7�ZߛV5�~��v�^�o��g�_��m���{�7Wq\9��^[�m�wﾶ�����������-���ﭾ��}���4ҽUTu��QQu�z��:��U�M��q��i}�)m-�I��e��D��"O�� �aKI�ٮۣ�5s5\�:�j"`(Q#-�$P2%��E��-�4$�f�ՠ0`d�HT�_�;D�R�u�2~q
xP�R�S�& ld� c%8Sȓ���u�	��gL,�$Ȑ�C�l��{��/�m��t����N�\SVEl��ϳ)�$���9��T2'R|0d�z9��DI�@��i��Q�4 jxX��5?|k�n��L��D�����@���M$�3�t�P��HS쓂��&�� i�CfP?�Hd��<-����4~=����04A�����4S�
22�(�a�{���ͣ�D��5�Hv0=�(N	(�H����I�S�JN��O�Y���4��M>c�]u�_+����i�8�n5��8e��2O��9�rd�H�
|��R�,$�B� xYFA$9��cȓQ���2a�"D�OA���C�f8�)���Q���I
1�J�8��0���b�w&���ۭk�	�(���I���Il�[;�4�C��LtC��R})� �Ry�ɡ XL���� o�[~4�C��C��M�B�%N���� i$�M�5��U�9��'N%H��ғsE��JG@��'��ha4�����P�"!�p������5��E�a65')s�p�:P���%�QM2|!��A�L���!�0I��8xX`2i��"����V����6���4,&�H)�O�
x0��LlI�m��m�|�^?+�������z��>u����i�8�n	��Y��&�7kv�l�a��|ݗqc�]V�y[[K�C����6����y�4�D�\-r�G\:�{�R��1"��Y���o!	\���}��΋E�8�3�d�N��VYHNʁ��GT�ÑV:'H*�qj�ښ���)!)je���'��Y�/n��z��iwfa���u��7O-����^��uuٽx2/�`۞�n��}�q~�X�n	Ʈ���&<)7�d>��3�Щ_G�I��D][z;:HQ!P���`J"P���Ϝ[����?!�:\'��T��d��Ĕ�bl`r `��a`�	b�����)=��j�7�nB�I�:0(��I���e�� ld�ϥ��hd��O�L�<,``���䀹�t+�Ç��@-�^w�X��N�́.���IDzp�pM��
����60(���[tM���}��̦g��9�$���db`�D@�H`���	FK��-�
|P�xPF��@��!Ӑ��7��.1h���䫊��d��+B���W1�4����	k�)k��rM���;m��z􇑐�ܤ��X@FI�Қ�RlI�ȈóA�F��Პs�n���!�tI�*k	F�Fr��`0�����~u��]G�GX�=Du:�����6a��ѷV(�0��~ ��"�-"e�I� מ��6$��'�M(e�(���DA d�ϫ�
�	��Z\'���!A	���J��'��,�N ϗ h�߻��I�:��M.�ETD���E���A��/5���Bt✈v2�C��͎����t@A�}��d62M�y��k�]C<N���'� �����SQ��OCe�2&��_x�E�N��!�����y��.������v,����UI7�'���~T�75���H�z gGã�g
�螈M�И&Pg�l'.L8!��ZV�D�8��%�O���2 ��)td؛@����Y ���!��DM0C~(��X٢���nے��c�_�������~Eq��]~~Uu���GQ�]qM��q����T�و���r0�t������NJâv{M�&�] u�2��l0�DA�Pd}�$40�N��0�}�nCi?D:����r�7��������Nh`N',�S>0��6e6!p��<MA��6'�y��ZI�)�;ơ		��A2��S|'��6��%WwF1�&~�����6!2F�F��P�2"2L��Æ@�Np��]�b�Ș'��܁��pa���������/GPA���N�2���tK��٢�<}Ҧ��w������ú�X��(���;k/"�<]�&�Y�
pCZ��>����h��£���<|~?��M?Ǐ�U�#��׮���i�8�n5��&�W�}�"��	���C�/��<v"&JXtI��d����&��Æ'����ӸJ!R~ܲ~8X�P@��⯘g��e���h���9e ���+B�5k���롮���D�g��c	��9~���MkT2%�I�3D�����KsC��L8!���0�4$�d�skD@c!�TD7��=�d6��@�)�Et.Ho�`ߖ�x'ę��2 �g�� �i���5C���N�0��ț���]87]��P`�6wk�� �82T6!�@ą"��4$����.V��W��'F�$������}��|!��x���nd8�m��ְ�����Q_?:���]~UTc���|��\V��U/�2����B����Y��M��,Q�\�df"BWk�X��=�N<��7��A�/�b׍E�4gB^'0�e�O�w;�.��CS��S�ǃMUj�`(2�k����9aDq�D�'�o�qA��SN;�		'���#�f�$�u�����o}��OK;��{:n.��S�i���݄��ƋFx������͏fju����?�[�o�״�۽ӱ;0B�w���鰦2�C����P==��O����S�z&��Q��3P�)I�KS����	��IXj!idA��!�2%�œ�Ju&�P�d��SL�:P��=�6X�	ޘ~)�D����ɱ����;�m ����0N�l��@��SBv0��P:���L4�؇����4�3)�ƍ����XO�T'��W=�=�o����z���Nv���雀����� =��OFM{ȿ���_���j�9E����yQ�ט�c1�ĝ����6��|���pd�OE)-)��a�-�AgD��/��-��̖BNE
�Uu��6j6�+�M���414��$�<,�NQ��B�a}�6�B~���x�MGQ����κ�*�:ڽDu����Li�8����ש���E!�0�T0I}�^�\�D��&2t�L�,L!OL)�d��]GC&R��ո#80�B����d0C�)��g�M�C�:f}W��`0���L)�Ę0��YHz2z��D1�Mȁ�C�1Y���"�}��M/���E�60��)��I0`�$�����F��\e9pt��\C�9G9MToq��P@5"Uo�NF�J��>&�� ~�,y�d�I���2s8Um������:��$@��C��}��H��|��FCQ6h��q�hB��W��k]�������F%,���=3<1��W��뮺�ʨ���#��]q[4Ɯq��߬c5�gEA������� hi4aC�����kչ�C�4B��`�Q��h����q%��B�a
2N}�R�^�����IbT�e'F`2KJ$w϶Q��'�ϗ��ѐ�B����G~uu��*H�k�MX�|q����[7���p�a�C�%�H`��0L(P2���L����pNY������D;��j&	a<��R��Se1�d���&tiс�@�XS�UCc&�3�d��FI��I� ��v�7a4	���r�j	�q��QQ$8�~��xXCc����u���U���_�#����+�z��n�u�l�c�l)�QDND?2�5Q8!�	sմ�h�2`�!���u?	&D8�$�͇p��u��n��3V�u�w���lhdq�ԫ���n�fS��'�"'��&��:$���"~���h��r!��l�d�O��-�D����%�!~_�c'�
j'F�hJ�X�A���~09��*�ό˜��?��!�'�3�ãI@�3��Q>�!��Q	A#5���������$c8%I;��[�N��<;�N�	.O�̘�(�s�2��})�A�`�@�a0�dؘ2MTD�
!���~���]|��V��U���[���|������Vi�ooYZ�n�+N���^++���U�U��u�:��5�+�oJ��ek�ej�U�Un�U�z|��g���V*���YZ��񏚭u��V�FEz�|��u�*��b�+�����Z�\׬WY�dj��U����ڥ>*S��������O����YZ��Ϋ+_4�Z��j�*��u��Y^3ǌ�귥V뙪�VUeVb��Y^��3���VV�[kmm�k�VV�YZx�6�+*2��_�V>i�+Zj�\ekMx�ZiY�ek��+\u��MW�ڵZ��Z�u�+:�ۊ���j����Dm��u��ο3��������uU�+*��ec4��~~ ��>$�> �|*���>�1�t�G���:_����+\VV�2����j+=i��5���*�Z�YU�W�u�_�wg��{�ǒ�����7 JK>�W�z���N��X���r��jYJ�tܳ<�&ej������fc�fFs9�-"M�=fa#_����v�b%�x#lPP��~�aX�7��uGNKE�W38К��8���Uy�,�v�Z��S�s+���y�lnĠ�+��V²�ȣ` lq+�i�P�]"l$���⣊!c�"'0aE(�����x���S�D
D�V9�8�r��(!%nBW�eRHJ4'x8q��-�r��@*�0�8ʊ��(q���!I��*�c�lE��R�o�Uo��a,��,g�|t�����:9:H�6�9�r��Ze!JYۓ���D�X��t����V��`����V�,)Qbj&�LPX���YSE9�uD���jd+�M~��di�-�ڬM��&ʫjD��	4�JTX7\�����tU�@��nQ�Ɓ�0��]Q���%��!��u�XӶ	1H�����?�R3*v1����	-R�[D�m��]UG;��]l@��#WrG���Y
�|��`��`�P�Fۨ	\���&�R�8ZKX�)8"���Gpl��i`�l�v��Ne�R��Q7F�U�6�2�*H�m�&I�I�J"4?\O>׹��~=�y�c������ۆ��{���wu~���ۖ���{�}��=��ҫ�TGϝuU^��u��\V�1�8��
��rR�m�V'Rj^Y@v���#��֢ d��q! V�X�@F[e,��+�C����W-R�Y8��j��`���v�k+Lj�Tj�G+�cM> �Z�Kk�Uc��]j'l��ԡH|��cT�T�F���pdb�������7�[m7Y�ӈ����IH��ќn��֜r�q¶���"���p���"N���m5D8�Wh�jYkuIJ!����67)���Ƅ�RX�$�j���j�J�BB����7U��͉�Q�E��o{�<��ϔ�nIe��O�;��\�W�������K�i�s_���s`q�{���.�0؈�M�Rğ|��$<�&�Rl` �"pAB���?	ц�Ʒ~��B�M� ��r2|&	���hh!o��L��ղ<O�"�=�_+�[�t�z0ēΊ|`i7�/�@�Cq>6Xy�Ӣ#>��&�J ���M������Wg�����&��h�큰a;��$?#)�>�#��@ @GM#���wf_%]AE3!#�AI�*��RH/q��#Ľ<���1����=�p���$$�Òl�:� �Xgɹ��e�h����	5ҟ����F�ON�:u�Qꫪ�^��i�1�F͇�,v(������!�l�H�)� �ID��>E�5$�I�����%������d40�s�Z�)n�a�P�0糹 3S�l٨a�hC�(����I�t�o��})��0�@���I�C㞛4w�9��>�,��i<e,(	/��b���^��eb��Ђ�l��\�N	��ϔ�edMkC�>(�Ĩ"|'8���u}�>������A�&�")K�pna��r~)H�z'�&�9V��a�i$ֹ����7�~��c���^�W��ʪ��>UUTEz��׮���c�q�5�֚��آ� y�|f���.��ϳ*��KǜssF%(x$���x/�V�FO�?iv����x���κ�������s?m~x�a�Ŋ6��-B2G»XNYS�X%��ښ81_��EbiDKh�S;�j��:`H��a�ɲBz��zy�~�e��Cg�No�p8�6����Y�����٩ߎ��b�	!.1wp����<Y4#~)�_�T|��"��+�WU�xl��Jlن���gGU*(�	��߾�R�����'@�O����"H���<�6�^$�LVEf���h��Th���Sz[.$��DE0ϺIg�4ʇD�sx���-كҞ��)���nlg��Δ��b<z!(V*ę|�$�@�Rx~���Js���%�x`�8 ��Ϣ����v`$�zS���`�fU�56~==4	ù?L�_��8��ׯΫ�ϝ~~UDWʨ�u�+f�㍼qï�&�����r�dV�[���Ŗ-�t�f��lu����b�9b��#���s.li�^���,`Z�ŃO��l�7�\����X�E�T[`���KS�Gad���|���J�ڭRZ+k"t��[���$$.596t������fu�ߛ��)ۑ~W������ޕMO˸��U��;<fG��w��5c[��J�,Uyb�3�����G�<��dpP>w�:i ��+:[�fDؙ>����_?QV�d����GV�{/<p&P�'�W��A濾M�D����D_:::zy�쨭��������@�7�ލO�ܧ�h6�6	�u�#�&�`(W�ӵ�2H�q�E �vFԠ�M1�0D�?C�#�"}��o���>��W5�W����W_>|�����UN�u�l�q�8k{���Քz�/#;~'d-�b��NW]KW�4;������	=��F�0�~�I��\�O�Ǟ�}�A&�y�V�:�<<�Vޛ6	8Q���rDL�0@�:���F4�$���N���~�������ɹ<��ڿO��o�Vpa�@X�rף632�t�a����B��r{���pL�!�G��<6	7�p�?0�Ml�׏��f40���:t����|��**�+�TU:��ό�͚6l�g�&��(��L�kҷa�l�_�!�I×y�.asР��n��w'M0s�\�t|��/gCe8	;O|���S~x�-�*�i�����̄*��f�G�HF:���������}�ws�<!3̞u4~4	ݯ�]�f�~��8ǌ4����m�mE����<�2��`hHw��M~C��Myp�[P�I�II�����h��}�ڜ;ۦ����G.���LJfIM�����[��S
`$���X
fI���($e��g:�K����ߝ]5��~~x��_���������UN�u�l�8��9���QE"vh�d59�r�<'���������=�z����q�W����B]��Bv��c�*Ir�%̊J��$u��������W���H{>)����hm��H�?|�G�
,�:'�z�,��¹�B���J�A��|�4Ä9��<�g�A�CP>6~��zd��]�`Q2V�h��/��,����[�_��؅"�
�a�r	�Ԕ*���\���4��<3>G�GU]TU#������ŉ����N�wTs���H�s,��<� �cY`(��,�V��LPPu�[:%e�
��K+Y��;X3��wV:;�2���1����9��TڻYjR�	��6�T��&���P�c���Y_$�d䱒	�Ɗ["�n�����*1b���=ڧ{�ڙ"��CX���޶��I��P��j�3g1�GqaVM�`T��������'�n�$��7#����AN���|~5���vhB�},ׁF%:a���r�����h�aE}�B�����2	�	��",gBPI⹶Q<d��xϑ��DDTV<A:Y�0LO�>4L��ɣ��&y��0[��z=�-��H�=#�9���=�3������*V��	��W!�&�~����rf��Vd[]�u�.g,���Z1)���HB�NA�$v����GO|3M>��b?":��ꢩu�l�8�f�����M��B�D0�M�I��]9 �>�|�DNg(�,��<v��u�L�R����(|14?{kZ!� �~:S{E���g�( ��"�3�����?M~��?pi��O'D0�~�/0�5�G.ax���&�Y��xRŹ��]-��Oh`"o��%߿}LnSf3Ʌ&�
	���S>����D�Ý#�
/��̬.����צ�<�FMHHI�va������Y���~eVUeu[�mY�qX�[S+��m���k��u�>x��k�Y^�u]oN��u�>|ʬUg���n�+�Uej+궪��+U�W���ʬ�UZ�VV���<k�֫]ֵָ����k�ޕ��o��Ǖ��ez�V*�Z��ֽek�dj5Zm��_f�Z��+4�kM���V2�Z�W��Z�V�2�3�~s5�����������c*�Z�7��V��u��ʬ��+�n�=z�8�����͵��Vi�kM�u��V�m�j�X��X�_���|�?���k�V�׍t�j���^+wZ�:׫�����j����j���k�պ��Ǖs]c󌍣}q���_����z~e\��^Uek�em���V2�Zⲵ���X#��,LG±£����o�m��֚�j�X�+^6��k��*�+��ڭE{�c+\c+J�l�ώ����|]C�f�$����!8�<@1$�f0�0�݁��YY�8��!��97+1[
1�3��8�Gd�XBTY �`�P3����9��E�#������~m�6��뻫^��M�-���������{��n�o|۟z���!<�U�]|�U�UU�ER8�#li�8ێoMi�?�i��%_L��|y?�u����&�|d�Ŝ"	��=*��nt�P�&�?��������Q&��srD���e����O�ŗ2fr����֝B�T���T���z�QF�,a&�Ć�&&5|����8�M4���i���(Bt��;�P��!G��|��%�����wd��z{����1�L��Q0|g
xl�a�|��:��TDu]TU#�㭱�8�n8^3L��>kMhЈ�fh˔�{�F۳GӧO��i��x��?m����ƚiʏ��55t�]�6�wf��}>��4^|'����罹I�6""nS���mvl�ޏ�rCRY�!CgJ7�G����_F�F,B��V�fT�LY�^�Xt���E�,߹�x��Fo4��>U���~z~��]c��DC
~�fMm��2rj(��6�����=��!�{�r,V>0���4�|4GQQH�|�c�6�8��ǜHJj�\�7pO#�f*ُܶ�5l���4,�[x?mx�"��Z�L�B����_����@n��f�8�Bѩ��n��j+kt�ƀu�� mH�"�i*�W_� @��!?����+��ב�I���3_����͋ҚƮ�mV�wF��ƥ�:�j>�S;l���'u���!gVr��UL#��Mľ�3�"#>���X~����*��iN6���iV�o�6�M4���ko_ ��Y�B9 ��;����Kl��lDL������B��ʞ�NӜ���kT���{ť �˩ބ�,�C81�h�ȼ
r�6v�i���T�_M����SZ��tDbzR�VPC?
v3E1siE���w�e/�m�=q�u�]UDGQQH�|�c�6��g���qm�Z�4�д�R��Y-S��S+(�U���2%ZT���ˊښ��j�U2CJ�Q��&��YJR�V+5b�)8�*$*,2N�Ĺࢂnц���:aÆ�'�3Lb���>�D;0��A��(�j"'��N3�Z6vBBM=�
�[�b#�� ����6�R�p %�F�8��xNU�YU���pI�a]!��k�=�,To=���&���~.�\h�;^�58&8�"b�D�T�Zַ�lMQ?JD ���2>R��4�O
�(��"�U,X�mom32�4�ci�|g +�Y9��壯#��aVbqȩZRr�U^ ��QE�M�3�7�֌im^Ӊ� *�6�)�����VU��X������h�Ġ��U�/,�0�g)�D�)0P9��p�@	�ız@T���3t��{��@����,D���AkRT(%B��L��[��(!�J)�3���xzp�C�����'��>�5C��C�����s2,�eN���R�A�S��F.������4�ߋ
rK$��V���ZxW�o��yչ��ax�F�����˫��m>��?R�=��]h��~|��]UDGQ�ER8�=m�1�q����օ���K��8!M5�O��{���lDޏ��l����[e�w�	��!�%,������#�0e���!D��~��������s9_ͬ����ੂq�:Ւ)UV���gNCA��}�æ���Z&���*"f"�(�$��$�'���(���Ƅ� F�S3$X�8<>8~���~7��)�G�yL�r$3� G��N�>4��>:�?:몪��":��G�d�"�$��8�tY���K��։
��FCg�����af͛���hA�0��!r��D�+�˳�Rs2�և\���N�A�̒��N1J�]�4z-�@�a�@��¸����v�؆�yJo�O�4h��S��T�����3"���?�&��<��Ͽ�G(ڬ�����YW�>t�A@���j��շaɨ"!��&&�ʊ�����]uUUDGQH�8�lcq�8Ǜ����<����q�h�2n1�,m��QJ�+Q�fAL�s�,#j��H��O��+�
�Z�LE(ґ����E���: b�:��v���D�7I�l�^@�!	[��+���*Ց�[}?k�����7�u��S���Id�>�I�9��
6�����]]\�:���D:|h�ٸSzE���lD4|k��ko�񣇓epTM���&�4"�Jo��ߢ�GS���!���].����tP����p�H>����������A�}.1&/ɪ���.�������򊺭�7�4�V��7���f���k�jʂ��4�J��+���H�>u�Ϋ󮺪���#���qq�1�8�}x�ٟ5��i�gO��@���>�s������aE@�;��٦�%W7rS�MC�Q���!�g%D>�}���m����ÆC��z3Bi
w��*��E��X�?Kh�  X�,�[Cj��Q�-cE����)��j���l���O��A���I.TGF3~�5H���M ���$g�e>P�_A>;��tۅ"x���x�
#�.t�M4��ǆk����":��W�cٲ�6[汚�QA��uѽU�+�"L�F�]��X_9�����h��0��i�6l}��4�1U~~~|��cG��a7��U>|���BY�ƒ6�S��#���b��إ����[E�����^_�y��L�!�<Kf�	��99;����9�<7��	�S)O&��O�G��oO!N��'g4==)u��J��؂t�~�Of�&�p�o�^�#�:ꪢ�":��Ҹ�8��c�<������hB�|lד��g��>�p��^�BDM~X��Kl��7�̙*&F�R6�"�O���thn5K��Mo
�f�i�va�qSF�i�������z���6��5��7�y<�?959������Ї;C!�}��3�d��2AG�H.��K�Jb+ƏL;2lJ)ɹ�~�lT��xhD,d��)=D�<�ĒK��x�?z|l�DC�0�U�a��4a��	0gL>>��h�2�1�����4��1��c0��a�X�1���ee�c,cc��0gF1���c$c�0f�P�4�
�@�$cу�C$��a�D|�=q�B�DDq�":�Q�DDDDF���lDDDi���q���c!�1��#�x�+O��ڛt�Ҿm���h���u�u�m�G��:���>UW
���Db"0��#�m�<|�^>W�X�R�H�<G���0`�(`1����1�E+%iƁ�)0U7��Vȟ$i��ȏ�%Dp����G���cq�q���;E�b+dc��pn'T���z,YyZ����a�{�#Y�!H�w	k��qB�[`A�U8v�W��eO���͍�6�I�H�m���1H�I��^�3�o昨0AN�z���b$@�<U7�,i*6O�T�ʭ�8T�`��r�I����7c(�b��HE�H���.���˃�,v��r��vzq�C����±�U��K�t$c��JIʥd�j �o�H�-veY.'�,D �"��eUHG
�L��g)��ۃ�
�-t�U��QJϣ�$3߳.BMaM8J�Q���\��@�2�cCO3�n�({f�۳DU����ǪI�Ev�ٹ�V<��e�1�R�\�UN:�ܘ��T9dr��am�#��*�d���V6�ll��_-��:NYb���F��"�&V��vV �X��Kmm�p�&ܶcq�슫D'Z�5$��u�&��J�DDՊ����Q�@���[H�)�NZ���Tm��pD����E[RU�r�]'-D
&J��țO�� �(	�8�J�$q��ěU���2�VJ��9-�$�XT��v7#���!,����6��*U[��X��l""��b�9\)x�$�ňN�W��[�kt�{�n}뻿_��m�M��mϽww���-��[{�n<���GO0�xg]UTTDGQZW�cb��,K��Ʀ�TE��!S�ҵZ�[#�����*d�r��Z�uR�%(�(�$(F����1H�V�4�p�F�-u��n�+�܃���"#m�j�$�6�&�B6�U��WT�r�'F��-NJJ�\���Eh��Yl⊑�P�e�D��q�WUW��\��ED�N1��\	H�E���d�8T!�؜v�HJ�b�����%㲊8����;F�m��@M֚	i��riO$� ���ޮ�W;��w;��c7=�)w,�F���G[��$pT�����W���Nl�T��zd=�_rs�$��6ޘM��w	L���.�Di��0��,�(0������dT���u��s�O�s� ϖ��0��#}�(�JO��S1�[0�s��ЇǦ�x.n�B��̭sX�V�4��m�����4y�k���f}�csM�=x%+Q�&�S�QU�MD%����A�kd����h����5\"kɥ����	�=0ɭ�o��+���͸��Vշ^>UUTG]UTUDGQU�q���8�t��! Bw

�{�Y�p�������m�ʋ:n'�9��vhC����5��9�O��b���D(����6l��0C����<h�<8 �h�ㆦV~�T%�ߛҍKH�Ѕ��:��rf,�iYTw��{ޚ@�"H;&�.p���)N0�}��ۨ�ГF��
 ��M��R�M��ƚ��޵X�o���QuUUQDUW�c�q���[/��O:y<�;٧�SID�5mC�!�ѝ\'�x|�I4�D�8t��DLL�6���O��鳳�a�DR�������Ub�0N����#��;���܋˫�ʪ�O����N���\��lD�<��S���A�qg,B�w>�DO:2��a䕌��i/�?sy�h� ��uL�!> �@H��X�:i���u�TEUTuU\Gl�)�e6l�PD)gO��Zur�)��B ���0�z|a��R�7Z�u?�Z�:���GZcMGj��R���݄W{k'�x��J3����e7�?9w�8n�ya�y�7*x(4���1%�O
$�-b�ѽ�b'�\��e���.�O��F�=����ߢ�l���8~����:a�`��1���g�na�ϖ�&������ki�g�:xt�=TuuUUUDUV/�,Q4�X�5��P�'=�Rc#�m����V��r��)�[��]B0�
��,T U?�U+���T�Z�,�'�U�F*ݒ�d��lr�ʤ��[
�)*d%��+I�V��? @���u����y"�����lڇZ{��~_�{}���=��L<��S~4�r���}=;���b-S^)qþ�~�g���;o
8|a�cm4`�2k�k�>����dsK}�H�>;C0�,�/�UEQ�|���	$A�$K�>t�e�)��_֦\�|�>	�ʔ6&�b �=����W��еl:��i�<�N�u*<2�;�G#��RM	O��^QD��+Q�b�t#���j������vE�ш��L7WF	>90�M���f�ѣg��\TWU�UQUQ�EU:3�I �� ��n&���Uu�! BQ:!r�(b�y�&t�A��"(�
D2���pѐ��X��)���S�~h��?�����M�c6����W�v5�Ƅ��5��(��<��L��U`���&�l�*�jX��_�b���oEFzo��:(xu�D4wZi�~96M�np�ƈ��5�k��y��sY��xǪ�"+��������"���8��c�矵^-�袂!���8L4x'��9���'�٣�)�D=�Wz����kU458z}�͝Dy���o	�j���5)�̎��dx�Nq��i�*5u6��)D<Ƙl:��=8s��mK"|~6hC�,�'O�7��OY$?u
y�����I|�$����Z��>�ș��a�����hTA�q���*!S.!�0����^���Xl<u�G�]G_�UU]DUW�c�q��ƴ֍4q��S��ø?5m0�|>��Nx�����.��Yŉ�	?�<rZ*��V��_
X��ax�E��m���=4�G�,���(������:!蛟�D��Q��h؃�4�N��4�&j�Υ�q�IeY�,A����-��&���l?n��ds��uz0C�=>�
t��.֘omD�j��"7�X���d1x�x`0���?>|����*��"*��㍱�q�8��u��w7�k\q�c�K�0�ZW�L�3g�[q�����/��)UȮd2�¬B]{��mƉ
�U`�h���c��F*�Bp���'U�YF*�"���i�82F���)lB/� @���=ZVlNW2I�n����VW�]�����i;M�m�$�T��\���+i��VE�O;���3��R\څ2�DO�L�P�&�����}�4s��=U�s1�m��3��,��SI�4$�~���?}5{L������\4ѽ�q����Z��N#~�&�0�����,�sF����V�p�v��Eѡ�dJ���s�����Va�B
&Tbi���^"�����'#c�4 
Һ��A1�����ߓI�v�������!���a��>W��**"�*�"����0�)�e6l���EC��i�A��/�*II��4A���M��N���[Ls&������ۡ���}O��\r��<8ad@�>�����(F��X���?�ߋ�$��q���V@�h��~<��90�g�h�ZhJ!҈�t����Do9B>�PQ��Q�.Yc"bYb��
a��x7׈���z����|���G���Di�z����GQ�c��`�0å�1�1�"#��"8��Q�DDi����f�gF2���h�4�h���4�"#�""6�p�a��:2�0`��C,coDb#H��������DDDF�z�8�ǈDDm��!�G�m�4���V��<t�ңn��͢#��:�ub#�Dq�뮼|��*�ª�#�����"8���|��mz���n4��UiU����C��㈈���;;����M���'�T�������[�������閿ڮ�H�6�x�פ�o���J'{���H���y�y�߾:��O���W�fF�kw�7#��3q�\bBó���R��ܹ�V[[�y9�wZm����f�wq���Rf�w�ǌ�/Z��Ǜ]��m���~n<���~�����ow�ǝ�߽��6�n���5����4�L<h���UQU\Gm�c�1���U�n�PD9���'�Sgob���;��$ ��\�;̰e�b�
x����
�����y%7�Ey�!��!/����c��x2���kr(�Z��̎�]^]�M��"
a�ό�<׹s0��:�f�{��v`�v���g>|�n\>�ǆOxk)q��B!�|hQЉ���&�������-��eiӠ�4�Mi�^�7��1�x�]D|��**"�*�"���8��͔ٳ�PD5:a�o�~��Y����0� �`�
h��{/O�/��a����쌍�R[��ӯ�h��7{��ܧO����hЇ�P�|Y�����m��:�'
���)�����F�"SE=. �G;�ġ���V)�D��\(��5��e�(]!rB� b65}3$��{�G��l@��_ ��.>������3��A3���:r:]x��>m���|�UQQ]UDEUqq�1�8�]��y�x���pL>��.�匰axA�.j�oo��zQ��ܓ1T�fLN	�y�Y�R(F��
���4�|����Z�"���P�9N���aGHe�RY��ѐ��B�m1kd꓿������n|=_Y�d�\����z|���
9K
��c]��*|2ru���y����Y�9����x��'T#���ɤ����t��Q�J~ѣbo��a��4aD5{T��~7)���`"�>��6lQ�e
!���ŷf���(��j����`��ϐ�������D�(��<�(:/�DB����BhѣF�C�S�d�n~��:qb�܋��kX�|@"� �Ti��G]��Z4��+�We����I������83�]��lD?'R`�|�N�\<YeY��><xg�5WUQU\Gm�c�1�?���آ�2&�pf0}hA�w�*%J]<HAf�+&��W/�Q�C����ڹ����6l���h�^)BO��K���4��+��W}�˜�o���g&��1 XE�R
La&��y(����e=�� �M���<�w���!	>$�'�QfxE#v�zԋ�1U�c��cv��	P�(Ӷy<̌����x&	M�g��'��~��8Z�3M<�\Ή�D�?&�?��}(�l��DA�-��N�aɣo�:�Q��EEDUuUQ����f�R�ٳf<��~�y���|PD5���&���-���,!�� ��Vt:���T؈]�g�lw)��ne30�ؘpLh`�)������LB��[ʚ�#�%��%u7��h_(|W��b��8�*K(��13�0�=
!�ra頰>� �
fߚ�h�=<��иhDB��ڠ���}��rb�&��x�Z����^�|��Ϋ�ϕQUU�UTETz��1�q�q�Q[
����U����*bB@����sϏ�U�zh��`o������:A�(�H+�CII��G
�QSV0���%U�V����Z�$�g
`��M���p��o�.\�4R���D�O���`���c?*�M~;�Tѳ�l���~F��zy���M�U�H�����xs����:p�����tlD?o��6~7o�30�4&�p%�b]k��玱�������*�*������\x�1�8�l玵������Z��J�VfUf1\'	�>��~ս����l�Q�B�g--��XX��8�jpuD7t���c��Wm�lhhEjN+c����B c��ߐ HB_��gEZ��'�Vc�帲l(�b��8A���pL�vr�"�ڥkj�g3
*fUI�����7�x���N�#��3��l���31UR�	�����w�L�:�n������F	�L�ᢈ~�w)�~J�݇�L�~JJ;�I"��FIPa���_Q��"aJ$ɳ
lѸ�liOH���}��̬�2��#�Ovz?;�Η^�!�ɓ'���C��g�-k�ֿF��<n�VV$��r"�L�����*|�gNDx����ѳ�J"N��E6r>�l����~|����#�"�������ǌc�6�?oִ֍4i�i������;S4r�"�@��t:���F!��V�H������Jf_0�G7ErMvg�f� ���:t���]-0�?�" �0ȅ��Qp���z�e�hжc���fk0�-R��N&����XG\�7�	���JS�B�&�NO&�`>�>�y�6���7><(��S������a�E8&	�ע���&h�RMG �ü�+��QF���ʨ���ꪪ��=q��6lن��ni�࢑��D��e)��4'�}��.3A�DD�)L����q{�������g�W:q��:x�l��Β�d���$$)�:�;��2U[�/�X��)H9+M���-V�Ƈ�U�Ĭ�� ���gyޥ ��gW���F_�ʪ�԰�旹!D�$���L����5��a��u������v':����F�����SG����ma�f�+0�R���O���"�*������\x�)M�6a���Ί)�98~���J|#W�tD���|-N���3�RZ~��P�<�J����H�
\��H��qQ����0�.3(�=?R�~͉�q3�����������|X�i+Z�fJ)L"~?B��Br�Ǵ���ق	ߖ���Ӝ]I�����R�1TT�0� $B$���L��4�X�����c����d�c��X��bc cc��a4�	����,��ec��1�1�`�31�2���h�i��""#�F#H�"#�Gf����`��1�1��"#�i�DDD|�Dc�DDDDDGȏGq��"#�B"1m���#Ɛ��mP�V�[E|�j��<G��Q��Dz�+���>|�U[*�j�33	1�c:2��(����#�l���V�[W�Tq�#�BDDGDDo޵T�;eƮL�ݵw�83�rW�;�
D�ڱx����]��ZZ0C�X<1F!�"|X�W#P�0EY,&DЖI���������XK#c�`V�o�TZ*ќ1���H�Y#R�9JUX�|�7,�Jr;HH����b*kpXF��Ȉ�|�ebY�����P����V1WYHӊZ�JH����&��m��}:Df��	��ч%h(XY ڝq�U��Y��
Wt��$Q�DF5ٸ�(YڥK&2���9��,`��%�x�PvX�{��]z󙹔���-pؠ�'b�yTr
�n`���;33�R��V5P�+I#���e����(bS�;��J�����6cPU6��w�-�
Sb�%p�FaT�S�ھ�)F&��@ݍ��"��Ռ3�Y%���2I�����2:�vā� ��N�V��D6�$m�X�p^I �V�Y`�J[b#�DBS���6�v�*b�; �u�q���IT-*Q��%��;j8���XӜ�1���8�mQ��,�a]R���])T�h�Gh�cu8��r��R��pm
آ�#hh�'�����p`��h#JR�`'NR�ۊ�����7���-�B�"`7$V��-�%�KT�V����FV�M�aQ8��V�bB�ʬrF���*�\������}��}���������ކ�m�{��������ɶ�������9U_+����"�*������\x�1�8�n4���\�vHfN9b�U�E�Ki�Q:���e�pD1�^11�(����6���8T�AE\��`Ԅ�BH����RUZ�u�,��(��	p ��&�1��1����n�:V!C�D�t2d�5F���dMȚu���lI�R�H��@FA�KU�P��˜ Nj3(�%n6�UH�V[lMc�L��WlP�X�V�X��UH喦��2��!�"d�Y��9bu��"���4����c�Oҟ���뽍6���1_��s��^��:�V#׮E�es���߳�������t'Tb��N̆��K�0���_�]i"�+gK����;Ι��x��ʷC�Yż����լ�#�!��#t��8�x씹�K�W$�}�^MTJ��$�fL́i�����H�xz�\{�y�޳y�־/:��x��G�E�
{����n�f��0E�����d!�����WkM&������sS��J'�<ݼ�����Ϟ��MkU�+��|���"�������ǌcٳf6(�O�2y5dÓfL0&�Q�y�A���శ���П|ع��DJ�+�@`|}�����t���t�R"�����Yf�@h�����|mN���ù���m�N!�[����	��E���q�L��>�����ӛ�ۻ׍��?9>sWM����Ð������t���т	ᇻ�t}��c�]~q����Ȏ�"�������ǌc�6�~כ�>kMi���᳓�`�Y�y֘�n�xvR�m0B���9�Zՙt�gӧD��=�
>>=�B�A-k&&��D�IN7#��x�ƉB[	E\�ʊL��/�I�gOs�OY4|��QBqm���N�O��9:o�����7�dÅ0�����h��VXQ��-�f�x���V�,gL0#����G�:���:������*��1�c�8ۏ��k���E��8{��i�TmiG�[g�L��K�������ӚqbB����Cs�*R��cs��/�|�q�ۙb� ��j��N!4�84�;>��YQ<�ޟbE�8xw���82�O9��b�����HB�4�ύ�,�/�98�5�������6a����d؈&3�<�S��m/�M0)����{�g�{�~b�G]Wϕ������*���1�c�8۟�,��R'��\qz��Hqn7YqbrA8�A�9,#�
�Ga�!ȥ���M�ÕO�++��L��<)�!0E��%+�pj�*F��YjN�G��UP��N�Q���D�]j"���*u�	\��fA��1������EE����]X2ڼ��١`�[Hm4�[mr��0ַ�[��p��j*�����LB�����F"w��D���b�"T��fDg��s),(~Kڔ�h�	6x�i|#J�XLJ�D$����Pw�G7�Ǫ�ǆ��_�k�<|�6Y�f96r����=�̘5�uF��c	lu�o?+--Z��y^uD��A@���	�ׄ��g|�孱�+����G�먪ꪢ���\x�1�8�n5�ܗ<�O/�x�z��E�����:l>:>U�G�9����㇇��o0�;7��/��D9Q}�0����� ����k��؈'%8y��j��0A/�&�OM�=��'�~�g�Y)��&�[�@��D"s��;�D�s�Q&A�/���؈���tȈ֛s5u�5c�����E6rX8IHYA�(��s�"@$��U�ϝW�먊ꪢ��G�J �:t�'O��,A��$�>��[g��彔��õ�n6��ANTԁV�*����.��tRYk�/����$$IQ\���IA\åD��T�^
+,��),�H�MWl�R�m��ֵmo��<:Y����|�7�=�rB�f��.��s� �Ϟ�����Ǖ��t�wJ��Y
���6����6 C��H�l�2�@b��K $�J)#I���(�Z�A��ފ.Rst�i*���v`�����<ɽ�Wu̙�0��ٻ���5��Gc`,��9\�@�ɆZV)��C�f�ʛu䈃O��u��t�|P�n'�K�$��y@��+���[��I��Yn��?q ������v�z����VV�Gt� n�P��ތ�%Z�qN@TI3�pؙv��N����9��(�|���؛�;��^���۶bu��N�P�
%��� �Kݱ��3,JI`����=/b6�k�y�k>�|ק�dY7/	�ccn���6���S�J��AM7�+�ދ���՝�p��-:�30טb��T,_mUb����-r��^�EEDU�ڡOR����4ʉ��q��]%�x��+b�����-S8�Z�����5�
����I�J���0��R��P@���+�.�{ J#�L����$��&3�QJ8�J9]�H�yAgL �g��Ǐ���_��E|�U�:�"�����Q��1�m�_�ۋ)�8S9E�6�η%f�&�����m��RJ��5j�j�j�X,���Sl(���5��-6�%[P�حJکU���-&�(�LԠ��Vl�vr�ja Cʪ�k���o���'��As��2���z~�RT�!QS*����r�,R�㰈
I�ԓ�7l/|�䊕X�k�^>b� F�0D�zy�.���+�QB�rj�����BM(��J:w�9%�پ?�F�Ԫ�Y���Us��r|Qa������&�����Q������{Ǝ6�o��>|��u]UTU|�#�c�q�쫵
+���Y��$�V�T/GSí�
�k)�I�ަ�)hڭ̭�k0R9RvX�IU�Q9��*!ڌǌ�rr��+��q���Br�m9b(�lV�!l���Y,c�����nI#�[,�e���� �u��>������f.��nVl�,Za���$}T�h�Z�v�Y�|�q۫��G�0�ڤKV�%��ƒ@h��kd
2L�sB=��X'��O�O4<�Oý�7��>aJk��Գ�;��tQ>:�:x�99F��0�ι�˘�M��+ P�+��e�}5�^�)�r)��r�c��$���d��)�8�6'����*a�0���F~���#�q>|��u�*�WǍ��q�8��y�kZ4���4�(ߍ���$��H=$B����$�sǂ��By��(>ga%�/ٕ���6w'�4l�r�k�O" ��F(S	3�њ��c�_�M!?{��b2H��A	X�$���H�jqW]�O�a$����^B��'�x߼�uTUR�x`"�\ �'����n�`SE;4qz����FG)+2
4f04f�1�C0c"�i#�Ό��!��3,��Q��e�c,cIc��1�1c�2F1�c$��c4c���h��1�c,c#�H�R#�Gϑ�G�:�ZaDh�1�,c��2J�1�,h�#lb�8�<B"1�6�"8�q���|�!�"1�J�ZUiU�W�1UG������DG����뮺㯕�V+J����#�DxDq�f�Q�$d�2ΔH0b�!��W��U\E+�ЄG���Ӈ���Nè�j�4�(
H�>�����&�w�nų���.���I�i�l��Hm�I�(��R�,֚��[c��[[6�M�n08�_(CC� �	�r����g⼳>m��w!��{������{ͷ�wj��r�{u$�I��{W�s�UU|��ϟ*=G]D|����U�q�
R�6Sf��	熄�[^#��U_/�u�9'��rO�<�{�Y-�s�jE����F=Ÿ&�x�ϡ�/��WR~�)7�<����,ɶJ��C�f*������������jsվ�-�-���:|l�6�2�����t�<A��D̐dDDp�L59���9=�̛7��Iᰳ���<W/�H��Q4�Κ3����>UUEW��8�)M�)��=J�_��*���ו���>����Â���!f�9�_�0��(�RX�QG\��sv�I�׸/��	>���@��R�O�8������#�Dl��M�@�d����2ό�\���fN�FY��QF0�LDo��I�ڟ�=����T�B|��E�r��s�._����܈���SUׂe0���\f6�����׮�|��:�#�UTUz�#�c�q�5��=�֡Ҫ޼���Q�l�Q��4^7�d���{`7�!QڙGyv8�Aƅ���q�d7�ӣ���>4�ح�'a���H�TM0�+]s�morr0E�� �Ϧ�o���Mu\�~o|،o:a��zɝo��Wfl�K8x�U�f�陦�R�ܽ�������2�[�MFg4�ճc�jǫ�Po�?)���K�_��{_H�RF춓��ۛ�l�xY��:a��S�߷{K[0<o3�}It�OϠ��|�9gy}ډ���F�3�->���L0�����ʙ���a�0�)%�X���:u`/�&�%"�T
�T�ԎE
�Z�]D�$f,����b�1{���k���^ǲ�l+��,�f�=|�_>Tqu�*�W�4aJSf�l�UA5>)�a�.��r�p������[R��<�iM��qOQ�d��>Ň�>�g^��C�L��"������*�����j:S;�qfc�`Z{�O0�gA�BB��H�Xw��=�����KxntG�_ɏn�ܕF��6ʈ2(�Z"��1ۑ�ַ��e�OO��0)ؓ<v9�e4h�s�s�����ĒM/c�I<���{��$m���]��xt�����=GϑG]D|�ʨ�⸎4aJSf�n?M�T��E���!�Û_���o7��t~�PقzaC7��73f�P�N`�Y��g#�w�byP�{Tj �r �u$�*	���������G�U�jԎ`��n�j-KW����i�B~M�=?t}����\��R���,��qQ���8>��4�_�10�%L�2�p$á�|tӤ�?:�����G�Q#�*��#�c�qg5������>�Y�_+v�Y��q�v�K�$���Ͼ������|xxj{͍�j��jB��p�a�V�ce�T��)�nf�n5-)��	�A�}	<{O=e�^jT��Pw�A\)�ĝʈ�RXI�' Q��_<@I^'�6Ow	�����̓	@�!N����羕�ψz"4Eg(�d���ZÓg�PNOO2h�����"#�|��qu�*�*���|�UM5�X�~}���#2�d%l�g֕]�D�	G-�_ت��+���r�+��2j�,�����Ebk#rƌ�����p6Nk�p)c+�S���1��E �mN�KP'$�I,��Dڲ��&�O���Ց�ȟ	)$�D7e���� $/��l�!ߌy���E�\Ff+�'2��,ψ�b��G�cw\���n���8l��������G��W7��ڨ0���G����������w�3��,ã�j���D�f�3��^uÝ=�|�N|p��GΒf��Q��d�#����\_��`aB�ZA|:i�s�|�(�ᅜ���p�F�B�N�X���T�9,ev�Il_+>�Q�R�7�	;� �.�{Тu%&0�4�xffa�3�4э�"**��#�c�q��5��`İ��N}�a�p����<�-]�~�%R�"·�u,_�jޯ֝�;���._;�����R��by��t0a���
9'��?X���C��t,��Ǻ3�:�|h,�t�f�����Z������GoaqWʚoE��V���_,I��L0����u���sW�V�>��0�[�Y��M	B�?�Զ�(G�4�o:_L��g�h΍�Q"#��Ҹ�<m�c�0����Y�/t��l���7>20�>�?_3y�o�iU�?�����Ӯ?�PgLk-P��/���U^}����?�<,
}����3n[��[)y�����[q
9�$$��78i&cF*�n�.%���s���y�jB�Ě��#�)Ӻ5C0����?Jᄒt��|���ib�9�SR�R� �x��qc�Y�.��$,0���v��A:SF���<�m��M~EWϟ"<G]D|����Jl�٣
R�6Sg�3��ɿ8��'L��ѣKF�nڧ��|�҇����N$/G\��(���Ǚ'#�1���NJ�#�"ccMDO�����M�4��Wy8�����
3�9[�_���T���[s)O�3�'M��RY�P�ⵧH�%	�p+0��y�|�>E��{�Tczr!�g��h�h�t���|��ѭ��5�|nSGgD��#l~�oƕǊE~D"""f1�0c��c,c����1�c0��,��Y�$c�2��шfdc�1�"#���qu֝u�DGȌDF6��!��1�aђ!��b�1�1�ec#�$c$��fI$�c��1��1�R8㍢4���"#��DDmiQ��#�"4��]z�UUG6�#�DDz���W]u�]z�+J�UTDDu�"#dz�Q�6�EF��X�:Q ���1�2��Dq��R�UX�W�����:��pY�ǻ��Jژe&b���0N�<O2Z?��G���F���i��׃�q32�o����:��45��47��TA2�gc���9�"�|��p@���-[���Q��Ui��Sq�ƣ�If��>g�Ƭj�݄1F)�

AbCn7����m�N�^�8��T�OB2�h8���f �eI�(u��c�e��sP�H��ÅV%	�� ��e�&�-�`�nB&���Dӂv��j�2@hd��ݙf�c�$�O�P���Bpl��,u���2���7�̦���q�Q�YJ��"��F��bm�����*��j�f�+�AT�4/��	Ǻ�1���1�((;�*�ǜ��P����I]u3dN\x܊[�@�1�I��6L�Pa��ӊ���t%������r�(6���̔Q[eb̘�j����B��v9�4�8WeP�w�z,�~�n���ǝ���uv�Ƀ$N�=,�!��o=�r��s�8�J�,�*ed������6�l#�}��7͗�[DWڠFI-jV4 ��
��9�`�(�pnW � ��R�����\���N�btLmZ�*���ݠ�p����^,��p��n�h�+�ي7`���,�e��Q�]$N[��5|��C��+�1�e�R)P�!�D,n��9 �	��i���-�������R��v(GȊ8�hdT�I��cR�r�#Mƫ����"�X�n�R"�6���JQ;�,��X�(ԩ�PƆ�C ~W~��1��o��C��������m������ؒI$��{n��s�j���>|���u�GȈ�*��#�M4�,M����r6&���"��(�(�����H����%��[9S�M�Ы�%T+9R�	�℣���W%��Cj�G+� b������d��rr���%# pAcnD�[N�R�G]�;l�2F�c��6���jBS����e�W���!��L�%�Ȥj�J�#�F�,H O��
P��;U��V�GUj��M֤�͖Y ����@2*�C��F��[�J8����o�l`�v(�X�]r��9�$��j�[>�;�N�~�<�_����B�=���\�>�̍�d�-ˑ�u?6����r=��k���(��E:a�5>���>=ɓF�ډ��X��/�[%�Z���*��~_��a�+9En��A
�0��Q��G���	Oy�O#J,���,�&�B,x�ݞ#�4��|a?������?�?v��>0 ���:|Q ���|�U�+R6�Z���|y#
���F�f��p�;�Nup��ޗD�ފy�i&�#��K,��a��R:�#�DuU�#���1�-�t�Hgq(��
D,�xU�'�p�y�#_t�Ӥ����xF�/��!rbf<#�Q��ep�/|y)�u��R���'!�����:x ��g��eDv�(��٩�R�Q�h�U$EDG+˼�(�������o�zd�.CK~�s�&mo(�D�5rEϹE�0��D���/��������{�=�Q��4f�1�x����EUc�4�xh��Ԧ�U͈��U�}I���#���d�Y�P�t�@���fT��7�F�Q��|�A�3ES���q���Ӆj)�D�+?
��dW*�ҽMy!g�����\�zb&!%��L	,�GN�i��NO�(���w����,�%��hA�ܮwE����"��I��A|�����ګ����ʯ�Q"#���q��1�1#]�u���;�T/�����\r3~OǡG�x���:�:P����I�bC��{��Cm�1�BRT!B&���tF�x��b'��������Y�u�*r�߶�Us���{�o���O��/_jkmb�Β%���~�Msџ��k��w=�Fi&�Ӈv�����b�P��B=8����O!@�:.��2�
4��&���j�S�Ц���4m>a��L5��"9\��@2NQ�
I����6��WU��ϕ^#��>DGQ���M��)M)Ͻ̸���svQ����Vו�U�K�����+T�� `A�٘	�o��U�,B�AW�f5n$�L!r��2҅1G+�Ç�Rۉ��?�l�$�+k���9���ES��R���!QVKYlAH�j�H���b|�-n�e�Dӵ:��6f;��WjUT��TP�ːx2KJ�T'�mNW�@���:(#?��rI��:g�]������v42�248�O����^n����]��	*b��W<tC=$��@O秃;V�0D�3��H �(7��,适��3�P�`.|J�C<H�<O<8{-�ٳGR�N+�>��h�&��F�f�~����������o�?6�Ou�oZ�l���-�����xf�a+��wpriD�"�(��<x�](�<�3>S�A�ϔ�.`�>0�P) ���M>1��ȭ���>DGQUX�M<M5UO��}����i=���P�d�(x4g�}X�j|s�S�SEOǆ�+��xf�S�w�s�Ӿ~˖�4x~�l����@�{�ab�[�fn����Y'���LԾ:}��Nk��sB#&�K��l�=�� �>��0N,*M�� �cLK�O"ᄹ��Ț�����.�IM��x#�fe���]L4ru4�����fW�5晘��|�M-S$J�H�X��a��<Yg�=|��u�z���*�i��SF�~��W�s�UA0���˚�S��K~��uzs��YC��'���th�Ӽ|T��N���m�c�"�c_���c�Zp�r�_+Ԛ����#RT��D!��V5�](�)��-�|t�N�O��#�x�$��b�#9��Hb	5J}��{c��IY6����2�R�B,z'�7��0"}x�+�	.��tFr�o�Y�KД�
4�{E'B���)=�\t9,�\Gvd������Y���y:~Y�rzu��Q=|�Q�u�z���)��M��)M)�)�U�b�,��Ҟ_D𧆍}0�|�&�=�gd����:Y]%�Ev7l��*s%^U�[��Y	D=�����h�o��ӇƊn|Q�����a��|�kpf��x�5dI ��p�J;�<!�T��ܷ�`�=�Ѹ��sѦ�͞Dg<W,ER��G&������&�{�GJ� �\1�#K<t�����ʍ����DGQUX�AT�UT�O�둛㎫�X�RM�D�Ņm�@����6��eKJp���Q��F6g��t͘Y��YuLN(՜�����/�$mcO^��թ�*���;+���Tݑ�VY$�x�F�(��a$����X�+��uW(����8ܐ��*�� 	W��?��
8����w^��t��mbZ��[��I�\�_���\��вV$*�;��j�r4��C�÷g�ӆ�Rt���6�0�76zt�褂�R�(���=</~3�A�ȝ>ӆp��������E�W��J������H/���%�辚
t�-p�)���|����o>��y<9	?!�5�'�ưѨX%
~>o2fҬn�KG�H�H���J����**����脋,�N����u��ֵ�Y�Ǎ>u�=DW�^�Ub:�=DDuU�4��1���$�2�|��1�aA��1"���H!Q΅�(0��)�6ַf�N�;=M�9�K$�x���$�:�aGy�t�������	<e�!~+��G}
Z��d�s�5��^/)⯳g��ֱ-4GO�QTA�ԢBJF��Q���Z��~��uo�Xa�����SO����xڱ��ƞ�눈Ң8�Dx�">G���h1�1���4��1���fa��3X�2F1�1��c�1�DDDq�8��#���D|3M�1��K�1���f�lDF#�q�#��D|��cHBDz���"#�DDx���m�ѤDG�DDx�q��F4�"4��6�C�؇ȏX���1�U�iUUU��Ԅx�DDGQ��뮺�]UU*�j���P�"#�Ό��`C,��t�A�#���<|���#��BQ�UF�}���ƾ���~�o8�F^K�%z��b��]t�x�m����\�9m���I'{�ۮs���RI$���m�s���*��ϟ=|��u�z���"�N4�ǌm�kmkZUA5>9��9��5==98M^�m�X>�=0����y}6{=Ao�6�,̶�oc�M��;ȻQbS�/��(~��D�#��T�+����DTw4a�dC:i| ��҂�}�����4��""8��W�,$ [��0,7�(���($��G�۾"K&,�qϔ'.SY�𧇢`��)�k"�l��z�Mz��_#��_*�u1�f�g��QD�P�ZIT�Pg:�8r&��{6#���TQD����F�0�����Ս��۩���i��be.!E��P�u$39��
O�ZL��:U�$4�g��䯁<�҉>��v�ޥ̷�1���z<4Nl���3R��x�!�p�����{���
"N��IM��$B��/������/����y_>z�U���Zq�,UEB�أC���<�Jܕ[]
������'�,dU�uهt���Ƒ�4W2@PZ&%���(^dj���+�y������&� �f�9�j�6V�*��m�`�H�LRr�nG)ƆD�i��S�+��)Q@q���4Т��]��������<c�TU���ի���q�~�����<��V��.d��n�eP����z�kvp���(�c4~��b��_>m}_�MMM�?+�sέѱ<2p2ph��s��R���yE�S�"�G�3��?Jp�o��u�\F��Ӡ�ڦT���t�77��٠��s�����D�Y���ML6l��O'L�����������hIH;*�%�Zb�^�V��m��''ǥ6a�A<vD�jL��R�!E@iD�� F�Q���0������c����6h�	�]*�'��H��Po �O4�!Q�Y:"}�:�&*�UUm_܋y���Pک#�'�Y�Þ�ja���n�珮x�m8zl'#F �j���,�@>A�<_|1������\��DI��EW:?%%�;��/bT̝9���9�*(D܉�mFX�e�R&���'�vE'��I��>�t���É
y��bd�QF��$�,��؞�:S�����6�C^��L�K$��a�,�ǈ����c�x���GJ$��>��v�I���p���\�Y ����٣s��ᾟ�פ��f�'��̸3��ق����_��[w:�m-�9*$�OX�X��"<R���]��o2�&�_���~�EW�x�+�g��#���(���A��Z �.��$j��ӥx�PQf�y4l�>>���vdL�7��C2�M����?����_>z����Zq��x�oZ�*���^(s�8�I �2�AwŖ�(���E�AtG:d�,^0G��@�*m��CV�GHYA�n�Y�q6�FKS:��j9�/2�;�@I�A^�s�� E�Ш$<V%<��68�M�<A�
=s���Q9�g����Mw�zi��<��35,0���'�%<E�ZU�w��/D��Dag�:��=|��u�z��""�KP�����_bѩ�|��H��E�j����p+�lϪJ�(
��$l�n���c1�=D�䭎Z�1�>���Y4�ş5t�=�bdG$kD	`�g%������ѻUU98�(���V�|��FE@�JE@VbUB�U�6Q�9��#7:�<�߿��m_�������58֝}��99���J�>������:,�ק��y��՚��>���[x��ǆfF����|����Z��+�(��`�'�ic��p0�u-�l��'JJs��+^��[:xxxd>[gc,��
�9�؄A�3���ܹ��9����Jl�y�{J�B�� ��}ދ픫�(,��>ⱝ,�8P��s�{����LG�ޔXr��j�D��eⱎVID�N|p0�����.{
l��)Z+����돕U�篕X���QDzz||'M�0�BUU�R���ل�>�\q��t�d0��:�4N�����*#0���`������\�+i�t���8d�OZzl���+���dDx��� ��Yf|{R��ȵUϡ���TUE\�Д(�Ajn�GeW��uؖ����Q[�](lL�)��i[~/'n��o��By��'�0�<���]����x���>|�]F��Q�#����=i�6�Ƒ��������ւC�y�T?���s�5��>q+��ܦ��PÝ�ٸx!��4WR�'�NY�I�t\�s9ڎ��{|�uy5��,l��$# �#+uRG,%+i�J��
4�Jũ��$���7�N���ʯ������>����G}���ŧI��J:Fi#J:aA�8�3��;0<�֫~����`�(a�dK;��֧�4�Ee�&t�s�:i�_)��+lk��|��U>z��H���DEW�4���x�o���Ҫ��pѷ�l��ú��S?TX��Y� ?�#r!�GV��fl��Lnύ��z2��q�����m��j�G_=w�lB$�B�m+� >���<eW A����D�Eb�(�3#����|��0�̓i/��|���&&	.�2��o�������ǆ=>v�>3��{��|?�ٔҖW�UUUٳ68~��:>ݸ��������L0}�(� BM0���	�m���wPț���J0��# �!���"&��D[E�m4[D�dM����4X���4L���mm�-�"�Y",��8"�X����",DD�dB�D[""Ț",���-���dDDYDE��Ț&�B"ȑ��DDY"�"&�h�m4X����������"Ȉ�-�h�mD[h�mDE�B"-��DE�B"-��[DD-��dD[E�e��D[D�m���Mm��"dDM�"�&E�h�,���h��M""Ȉ�$X�E��������"�",����YD��&��e�B&�h�����h��mmDE��-�h�E�E���&�"h�dH�-��D�dDDYDE�5���-�"�""-�"kmm�m�"-�E�DM"""Ȉ��Y�dDDY�h�mmE�4H������$DD[DE�u�8h���"""Ț",�������h��mmDD�����DD[DDE�DDYm��im"[H�,�"�m-�Ki%��[H�D��!,�&��&�[H�,�"[H�,�X�-�H�I�K$�h�H��H�,�&�c��"Y"M!"D��D�m"D�D��"�bI4�D�d���id�D���E�id��4�[I��Y&�,�"Y$�i$ZI%����%�E��Z��m�Y�dIi"�%�C��ƒZId�4��Y��$Ki4�bD�&�M,I��i�D�H�D��&I�K$H�Y�K$K$�%�	mf�D��Ki2[H�K,�"M�K$K$%��$��4�d��"E�ĉm!"[I���[Y��K%��BZZD8[d��Z$�K5�JZ$�Ie��I-$��,�M,�"Y5��4$�I�id�E�ȴ�Im"[D�ZI$����d֑�Y%���i�d�k4I-"Id�iC�.69d�%�%��ZE���ii�%��ZH��[i�K$�KKe�%!-&�ZM,��4�M$��d�4��%���Ki,�H�Y&�H�[H�Y&�Y"[I-�K,�D���H�I"Yc�3�ZD��4�M$��4�M,�$��,�f�"Y"M,�K$K,�-�KH��K$Y��D��Y$�e��H��I�Ki$Y��K$I-�Ki4�f�D�"D��Ki,��id�D�&��$�k$K$��M"[I���D�m&�,�K�l���q���ckd٭�ƶ[f�M���Fhs�.�I8k46�Cke��M��1���e�[ [&�ō,[2̄�&4&�	�	���-�9��#B�'[��BC�BB�A���
!�m��!d$BC�9M�h-�BB�8��$-	���(r�r�HY�� �%� ���I�hMZi7o�Z��&�[MZi4�Zh�X�q��\Hܶ�Mi��5��D�M&kM&����ђki�&��4ɭ&�k&��&��MZi�,�&�kM	��M4��H�&����h�Mi���Hɦ�h�Mm4�Y4M[FM5�Bk&�D��I���ɓI��ɢki�ki�im4Md�5��k&�M5��FI��I������k&�2�h�&��&�К��4іM[M[M&����k#$�MY5�D��I��#$�ѭ4F�4Mm4F[MD��D�M&���De��MX�&���D�M4d�[M4��M4Mm4M4�ё���i��i�i��4Mb2D�MM5�M5��h�Q��M4Md�5��M4�ё4�[M4�Mm4Mm4�Ml�&��i�ki���4M9�82�hM2i���i��ɡ5�d�M5�M5�К&�4M4e��Mm4&�4M4КYD�ɢki�4Md�Mb2F��hMm4&�5��5�2&�YD""h���i�h�,�D�mE�"&�ŴD[DDE�m�DE��h�,�b�"",���4[D�,�hYLME�"�$M�4I�!h�����"Ȗ��"E�E���Kmd$Z"DE��"Б4$,�m��h�m	DL�>68E�BТE��m!h��5��h�BE�"E�kbдZ�ض��D��E��d-	D�D�֋D�DD�"E�ċ"E�D�""E����"�$YB-��"h�",�DY�E�h�H�h�dZ�HZ$[F�"شH��h�Z&��,��ȱ-E�-��dMD�E�h����D�dMB"���$Y�dDX��"-����h�mm��\m�"�,��h�m[iDE�H�"-�D�mmD�m"&DE��"�&��"h�M�5����h��&�h��mh�,��"Ȉ���[h�дH�""-��E�mв&���dX����&��kml���h�,��mm��h��!"""�m�"-�"Ț&�h� ������3���7>�B��Hz������������
�n��ǖ^�㳛o}soǣ���b������x`�%�w�s����_��t��}ז�K\�5��y�i`�=��]=x���?Qp�D�,�j�K�������]�_���s��<n��z�gG��66f��vޏ���������x?�� �dw���l͇�7m�����M�������o���1��Î�~Y�g���l�����g��x<�C�'G�Ο>���3a{1��~���*:vg/F�M���3����_��mͣNZ�vu��m�g�g_ÛK0�,;�m�6l�iu�^�/Vm8�S3X�ZnZ�>�˷>n�=�v8�Ͷm��q��&a�͘m��9�{8�6�[C3Hlo�6�`e �H�3����
K�ą�3�?�|9��t<{����MѼV��͍BLf�f�c
3e	(Hٶ���3��{}Zn�v3�{�m�m��{�^�i������9�8���s��}X����W+�z}{�-�cfl9g�p;x�m��N�Gg_�k�n�o��7j>�{��߿u�����k7���|������Y;fY�$���x�n<��}>�u~���1�6�������mO���������ή��?f��o=�ٰ潏xٛ���oٶ��������n�w3�<?[���gk���n]rl�ُ���m�M�n=U'�rӖ��-��Y�cm�0�������l&��!��D�6O�B�C�>B�ĞIɚ��#11��ۦr��m����[l͇n����Uy����ٯwM�=cfl>+�?b5��N�1�y��c�����w<�|����-�6x}/W./s|���z[��|��}F�d��p�����^fw�=�3a�q��yF|6�m�~��1�6M��{]�_g�~n�[>?6y?I�y���N��>��v���i�l��?Oi4h���0�d�$���Jd��~�������n����3��n{���n�Ͽ��uv�����}��m�o7js�q�z�ӻ��o��r~,���z���?��ۻs�gon[=�N:�9�6�Ӹ���~��l���DŶ�ﭟg/�rz6�='����ٞw��ݶ�s��w����ݏw�zݮ3��ݝ����ޟVq��4�������ܑN$�J��