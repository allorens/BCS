BZh91AY&SY�m���߀`q����� ����bD��    �}QIP��iE�P͔����UH����m���V��B*�*����[Y���cMĒ6 h���-�-�(0�}ń�����m1hd�Yf�0���e�dV̲`�m�"�ZUm�l��i�[bERf����T15��I6��[�M[�P1����M�k-�4�ZңTekP��,��6f*��i-mV�mM��d�+f�ZSZl�l-e�m���[Q[j6�"k[mVcUf�m-��dV^Nf	���c�  1�_ٻ�J�T�큪�r��u�a*��i]UwW���*�=-��m�� 
]�ΚW]�ekr({*mk`��j�Bi�N  ;��J��-���z�R��F�U�����M���T֖;׼��l��������Z*y׍�kW[�W�����ݺk�^{��\��U�����)]��z}�jڔ	�ͭ����Ҋ�x 
�������˷�z�$�o47�-�RV��<y�M;4��=ν:�yӇ��5���%z�#R��V;�,�����_}��S��U�w��65
��[+Qj���l�QKf�  s��ll�]Ͷ�׫�{e*�hOw��v�lm�e.�o}�)�����i��甪N���O:�5+,��z_{�J����U����ӵ�#�ǽe��髵��|�)־�wawޢ�ؕ��Y0[a��Kk|   n7���ƀk^�k�^6ݲT��tw�ུ6��|�}��햶��>z{��{�jC}�}��}�Kl�����:�Wvv����;��2�m���稠Ew��Ц-�^�V�SF�4�-�h���   ���GI��jϼ�T��-�]mԯgEڷ{G���Ҩ�w���l]��
p�{m������<��J�Y�x{^�R��{�d�*�[���RQ�o�J�Ch�%V��VM����   3v�}�%.�f�{ozm�uS�[B�V����\��]���m-���;�i=�T=���J���y�g���4і�z��m�F��z*�޵ު�Z)����"����L����m��  s�`}ɾ����Eа= �{�۽v�=ޫ�@=j�Ұ�����pz ����G�S�� ���y�q��Piڋ�,�kCZ�`6Y-���  Ϫ �z� �I��<�@oz��t̪����*�w��k�mA�<��z���j�ˡ=�\� =���<�t����6�M6�V�jQ��QC|  ����^��X��ݥ���B�]�d�z4�<��l�{Wz��x���+l8�o^�F����z��u�����  �   j`�*�hQ�4h A�S�R��@ Ѡ   )�1	J�~� �    5S� IT� @    "y j�)�Oʙ�F#C�jRSG�&�E6��H��Q�D�}����>����4��'�9���_/2vߣ�<�bf3u��~ �{�?���~
����P_�
 *���������/����@X?�UU���
�v��?�APE~o����Ʌ?f�afW��?�+�e�����������������	���+�+�/݇��+����+��`=a}aYC�@�������2�������� z��ݐ=_X�W�@�������������+�#�/�/���/����� z�}2z�����������/�!� z��`X���=`���(� ��	� �ّ�C�PC�AC�C�*��*!� 	�*!� �� >� ����������"L���(��&`@=a =`@=e@=`@=aD=d =d=`@? ��������������������"�P��P̪� ��(�������� ����"}2���"zʈ�� �ʂ������=e=eU=dA=a=`Q=eT=e=eE=`_Y@C2"�
)� 	� ��*��")�(��XOYTOXYQC�QS��"zL�� ��">���!�+� z���'���oXC0��!� z����+�~_�� ~�����2�?����������'�	�z�>�����#� ��>�/ݽaL�����{���������j�L'�*eXT�X;��I:���;�/~�r�A
�@P@lҖ�{��a��a�fb�qe$��+C�C�[�a��È� <9i]e1R75�5�����i�v؃��c�Oh���I����G��t�,�taسn0.���!SG^.d� �/u�"��ݽܼ�pVd��0��yZމ{-&��]��jķt�SE�Ke�ҜALvl4�$9c7hӆ[�<6Qr�X�tȜ�Ut��P[��J5VX�VO��%����se���Y�(J%�[�jt�+�M҆c:����<�����^�ݱ)�!��Ԕʧ[B�t7X2\ӵ�]�4<�P��CL�j�T�bb��ucB/P;K^c����"h��D��w��nmT�w��zԭ�1h�Ɔ��0Y�������b:��9�^r�&'L���� ٍ�r�ָ��ѣ,R��Sfm��f�pU���Qb�#�t�b�No�ڰ5���1�6����sFC1�H'���C��
cz�[W�^����]ܫ�Z�S���lv�40j�#=ɒ���J�Ԧ��P<Z���!z%˷�j���f�m�!b-�*��>	R��3.)���nL��2���k]�-�P���ʽ�1��{Y�#�
��f-���yEh��;�C,���A�!-=Ê<�����w��s.1�R�VE�4�dL��p��b�]a�f�6�a�`������S�v��('�σn�����Ǳk��y�Z�u�ψGU��u�,T�ց��{�T�YE`����]�?��l-%w�/�2ޣ�L'ffQ�V��x�z�P���4���rjA��X��ڣMk���ӓn��ֹ<��Z5]��$A���ڶ�Q�B�Vi�#���w3>�bM��S�x���k.=��{1#ZX�{`�8��)c/m����
�;&=��֨��zZw��MR�$��S�+.�K�w�s3Ta�^���j�EGq
Y�hF��{�еl뀧N��w�Y�)�I�FI�U�tUi��C6;��A"�Sl�O]�X��L/q������M�-LV�Р127NǗ�a�d]���^kz��;W�/Vf|ǹ�WNDsP�h�ك�)�����%Y�oz�eb�m�%4�㭢+�ǑSY�65�p�hh"�ܣ���`EB����bэ�Ҋ}���h"�K*�Y3�(����Ď5R�
*�u�����n��N��Xy�C��ư���w'�.ݡa�ۮyc��xo.%��V�c�F\3M�Hf�m]���Ы��w�j��� Q�m��bâ��ƶ�L`�MU�Ә��\�:3eS�D��0-6��B�s�v�r��j�7�hk�*J <;�R1m��1�fekF�RZ��sU��y���;7a���8$'
�hl+�E�:C`��U.^G�m�
�X�z�f��qQ��	�(ĥ��+
�,�2���:XaE�۫є��-.�+�e��S��j#��ũ�b����
�Qe���:�9y![��/),��b���J���@�{0�/`��\:����PB�)ԃ%e��b�_�%\�!y����:�������`���7L=A[�Ok5n���騦m��uvku� �&^ŧJJ�)j6�Bdw�˓jP�+/�t/<�o�xYvTAf�Aߡ���"V�z1[#~o9yBa
}3vkj)l���Z�xR53����J�dŔ�3/s�Mj�Kի�p-ya"� �:���Vj�*��B�%���J��f��+�ؒ�ȕ6�tZ��ɉ��x�W�u��W7e^%�O�uy��a��
���ܰ�����,�w��*k߉sv⩹d�6�ovP�f"�-�V��t/o.��ꛔ��a���:L�E�|y=\v����*n�˫e�vƽ��\�p�4.�%2;#CnҊR�?Tw�[V�f�A�,�Ջi�{*��T�j���li����L�=�[��"��*�sw(P:������Vh����;�OR�p7#{sf9���E�+�4�n�nMh�p'a�,m��T˨�A,��R�?�`�*��%nX�6�U�*�آ�f�Qպ���U3�n�k\�T����+�"7&�xae��$Vk1�c�N-Ţ�8	vYWLV��cwژ6�%��a[����Z�^��@h�O�]B��ٱ�j:���ݽ-�݁a�@,ibs1Աj��#(���ۣB�e>�)�\셛��崓q�`X,�e����}���l桷\h���v�l��#7��n�A#Y
4���UV�!�?�<p�i���MV�,&\ۖ�b���IjX1�%^e���e������bK���'�ө�੆�.�ְ�W����D迱��
���V�n�C��T�kiλ�m�%1O��ˊ$����̚�9���l�l\�Su(�EP�<��Y��H��˺B
�1��-�mI�yi�Z(fn�2J�Q��V��ڤ��zV;�B:�c�>w2�R��]��ӕ�K��ר��Zݽ<�SXֲ/)�e�M�T )8Cɀ�E�

-�j�i�8�e�:�D5���wLrJ��GRT@�H��]ea��7S>K,���x�RÐ�t�v�r˨�
�JS�uP-Z7���9�9�V�Y#�-Qf��i�yq:�AX�@6Z �W�j�@#F��n�@˗�K������$���dӫT`����D�/e�7�2�@6��t.���A�T��b�c�����דNˢKڽ����:��vJv���M��7B��4�[r��('��f�"-���E�5i�ƭ��)���	��N`Ua����.���8B�v[�����]p|��u�)��1f�sIB+Y�� �TAm^Y*�Sl�̦^�v�k���)���h�5a&��
�]�1j�C[�Gr�paL��-���Ŭ!�Z�7�5x0����7�;���Z�vAU+l��ko6�w��ݼ{�;]f��Y��I�[�k`���\�l�n�׬�Q.�������5�/]����=Ѳɩ�K2�{Kr� �LU&V�N�a�kwr6hũE*�EXcx�%e���\i=��Ir+Wg-l�3k0
�KdB����3V�&��X�	~E�=7��3M�X���P�fMF֊���F1�h�F�:0:E���4��{l�i�k�ݴ/>i�-�BZ�dC�Z��+0���4[�g|ﶚ6�"�
SxM�#Ǹ� ��R�:(�5`;*�n��lA��jج��3r"�f,��[�k;�nG�n��b麻z�G�E�VMj�y+k5�b++[X�ؤ�ը>(�Ғ������X��Yo,HZU��0���qQE���P�4������:f����O,����Uf~�1 J�^�N�2\9�5�/s*�{���Ǒe�2ݜ��5���l���m�G��7�,�Sն!I��Ţc%�Z��c�"��n<Â<�^ ��NӴ�S�5Ab�\yEּ�e�����ܪ �b���lG��j���1-�nln�Ӻ��&2��Z��ut��m��Gi!�Ͳ�Պm�!sI�did@���Խ�ϑ/�1	��-�0Dw Է1��-�`c(�6�̭rj�s�Fk0&E�^fҦeg�m\۩Ylc�Mm�����J/8ٻ�0����Gu��b� ��a3���1J��4K�+jC�g	8��b�S�Ԟ�e�{i?���&m2�*�v�L�4_ʮ�L7�n#e�R����(X֤�̅u�G����j��-{x÷vEX9���Lʣ���I!d�T+w�-C��p�7�Vܨ� sፑ{����e�+ٕ�0M�˅ԉ���P�I�v�VX/67�n�T��.}$�^��4-:M;k���ӫO2�[�V�1Hd�!�<׌Q&����x���X�3��h���w�Xi$�R���Σ���Az39���Td�6�Q��.�7��bY�:4��uh-�
��An�y��5Ri��z�t3k%ƂB�I�SK�lG6�	C)cA;��)�F�f����^�j��X�(Fl�P�[0d�����(�SAkiJ͢��nٙE�p� Ú��DU�7*����^�wU,r��u���AꤛZN�4��f޾N
�cY����VY�ux-7X��
V�����VU����'n�[)�w,�|o�5>��Ë�c�?�e����i�-����Yr:̛��V�f�DkkuB��&�Xq��f^f��Z��ej����%��f1����ͩP0���e�=�M��R*�������pCv'un�K�k
�^�t���o)fi+R�M�ͩ��<Z���8"׺t�TB�k�����E��{%�#,��X�3�3~\��>mU�F�Q:��%-�N�R(�n�ъƝ��dT(�4@�6v�Ab����T��]���T��H.��(�A� ʪ�r(Z'^M�a�%�任4�N�4>'r�)>�V$��v��x��̫��e��*�e����#@�B�2qD��Ss/N�u�r�����-�R=t)�L��]�6T��ևug3r���0k�7_��@�m��6�%�2��49�+7J�u�r]�7LI��i���
�j��٨����#r��sT�C:V���{�����&�)D%�CB�%L�dE�0V�(9D�52����E�#0�j�J��wl�{LKu�E6�Sې[6�(��K*�Eb�A��fe��4^2�,��F2�'Q��M-�Ƿ[M�H�	຺���N��m�M�B��ðݰWZj����B�����4`�wx0�[/Y��l�c�dF蝪���X1{��
5��j� Z̨� ��܊]�5j�#K%m��1P[�Z���[�[����*���q�d�i�`����a�,M��:ѡ��]��WQ��F82D����a$2VKSU�����Bĉ�a2��cCK��9W�X&Xf�k��e<0�J���:�K3�����i雳E�z�y@C����lWR�DN�1Qgl�.�b���X��$ǻr�N��I?n���.��1�x"@��|�ȈT[GF�^�k뷅�ԩ77$w����ӵ>�Mʵ���y�Y&;�]l1Y�%-�)�V^�V0]���+��G2"ooPpfͤ)C[��0Tr��4�R�#
���Ęr]f��m�dc��/>�mn)xZ����5�n����`[.���:��Q�40WD6X�wa�h�T$�c��`�t�蘕����0�k[����B�%<Y[�M��sZfī�[bKn�E0dg`��f[�lMNʑn��
7ysDhmf5M���%P;M�p��i�L�cD"�Q��c�-Y(����ޛ�,�$�í��i/S��,CS���N�Vt��1�Z�x齸���eL�6�\%�9���N��r��6�;�A���r���h4�D{vA�� JY���X6Z���d6F��H伫�iO�2�U�����1��"6I�n{2��K�5��Ktj���z.!V��Ǹ��vޠRS��r�N��Bj�pR�P�V�f�E��7vws$�X.&�L����l��o�%���0���r�����J���v-��7d{���	��z��2��jZ���n�P���[mI���opJ�ڎT��Ÿ��*��6�ܵ,�L]A�J*&�wo$���YR�j �[���)Mb��*��&�tat�f7"Me��v�k�`2�F4V�l<M��iu���ݤ�Ъ�TB���-����0M1�Ȳm�$���f`��Aʳ�aZ�4p%LI%`{�TR:�:�V򞫨06�9XY�ëwv2\9%-d9_�x�#_���yxvQ�)�lX��q|e0��g+f�wԶd1�wf������]7��輙�8�ă�� ��ڱ�㙺���l`��(7��0-W6 ��/uqi���ݳ��w�;7ɖ���I��8��wW�V�G�\O�f�t���7w!ӢSۢ�ɰ��BMSUo�jз*�^+�F:j�(���^1��Z+3y�l-QX3Ek�<�r����{xo
D̭T���kt��L�75=�dL<����7))t�8*��pދ.:�f'G�ѱ�f,A�J!
a&��3�ʈ��U��"��b����tjٺ�)�lH���ݤ�VZ�`���k, �Q����(��R�ջnLL��8��1,�-^���=�@�-u�5���n��|֖��[Ce��F�,mkl�&�j��%��H/^�aE=֕����3�`�̕m��ݫ�Y��b��Ӥ�A��H�(���3�nk�������贴���n�lp@S3\���4��e$�,22�ᶜ�A.��:��m�tF���M5M�4+��j��k�� ���^��a�vJ!���ۗ��ʘ�M�X�9Y&ʛ2�a�1=t���̴r�����iKvh�������7l��c�#�G���QM�-i3Xͫr�kf�n2+S�bS�MHh��y4�y��w:�j+�o��ŉ��[���BΔ���ͱ&��WM��*�n;S ��5�sX<PQq&�^ن<�;�,�`�آα0�)�Zյ�����n�V.���9��X�ӭ
���zs��4�n�,DE��`��zt��j�=�vA�+ӹ4���6/�,h���j܁�u�7�I���ڊ
�qe��YŇ�2u1��[�lY��i���/8��rQ*�>��r�)Jr���>��ʳʴ:�І�Eu�h�}c�5(V�ϛ��r�{�G���s\�Z��[�\�1�h+=I����H��~JG��o����+���?b���1(]�+NQ.zϦ%o��*�b�kJ�u����"����䬹[�%!���P�}�d�h�G�����Cl�&�`�4���W�h8.hWo�Bq�q�g6��f���m��XoQM￈�~�A����/�?�ɟ��-f�q�.\�%�0���b�+ U�x]���x%���J"ogJ;*�<8��89}f3�[4���X:o/�s�3�[/��+��
}(�9����'^�ZbD1Ս�.�R��Nt}v��蹓�Ζ����4�d{{mǻJ�v�#�7��V���=̎i��qaϸ��vu8%C���;���:�k�B�f�r��Qܘ���[O5b�L�5�܂˾����;��Ꮄ���k$j�f;���8��P���a�X�����Z���N�|��N�EQ��u�v��|���l����(���Ԑ��]3h���j�7���n�NA*��%q]*-�����2fZ�e�� ]���N�;d�9@�̾]�neKʛ�l��p�Z���i�tr���@	鼰7q��_M�9)��Z�,o\}X2�ًa��!ǘ�Xe�ȭmG��YW�-TjM��1��mB]�33�W�i�=�������'[5�®�k���PN>��5qeO�.ط](i��7`�n󈈭��IF�j��c����7:��!���؅�YE��G3-f����vY�a��0b+�����
�{cu����i?��T�d�

<w-��nI�]j
�r��
��2��B���w
����tң��W�D��%up�N�N�������*-H�'O��,v�	Ah��Hi�T��/9����Ō H�yN\+7R�k;��,v��"���V��0�M�گCy�z�=��8yT&�IU��,A��m��lKyou6�}�Qy�z5n�!��4s�fܻH����9���<]n�2�	�nQ�N���趶u�-�e5�Av�'e	V�ph4&���at\�΄n��s���h�gf��H �R�q\�Z�Q��z�:��>���+��.ũ�7 �|�
W��Rg�C�
��̭�������53X�x��y�=�o�}�� �������-�:,�k4�b���)��h�ݜc�hN�w9���L�g��l��1���:��W2��1.^ �d���V�\�Q��n�a���W��,�J�JZB�����gGuG7�cAAtv��-n��[r���J��}�Tb��Ve��3�;��n�
�>���^ź�{�����j���f�n����"%>�n�NٚԂ�m)��X�;�LIT1�4a�,d�Ӊku��L�n��+5�4f����o�=��\Y�Z��u�C\m�OLzc���i��ua���R��0��/)�*������_G�#�Z� �j�8R�[F�{h�ٯ!,c�Dr�K�S��E�|Xܻflͱ|�A!�juz5+��*�.u�G�a�1��.�I���=�Д�T��4�j\�ӏ+;06p��5�\'m�4�
u��\kᛍ�X��g^�\�E[�(�8̈n�n��5�&���D����Ҹv�t���H��ˏ��P�ĵvV8���+I[��(f��=/s}�Hovƾ�$��EV8�s9
i����c�!��_��aNSf�W�v�ʹ�"L�x7��Os ����۬2�Kx�m��
�m�R�3�9�˾�T�v�j���c�4�X�d��3p����V���o��|��J���!\׽s�;:��J�'GSޢXkG ��U�Ĺ��Ie�d��Z�s^�6��<����t�@eI�����lGi庮B'wN�S�l|�t�����T�Ϸ&'t���x���ɻ)D�Bz��(T�*�XG5�f�t��ys.́Y�������t���	j����cY�w�оFov���J5r��%���I�T�tӍ��޶��p��B*�U��s^�#F�����m����~�)E���}]F�a���C/�4�ߠ:�
8���7q��7�f�]��!�j�<�D���q�e���9{�*������F��-��d�Z�J���b�8�2
l�Y	�h�8֎�ъ�JT����kx�q��V���lқ<XT;T,�J�K��x���n�'PʝZ�����|�d�VrR�+{�L��gu���3�L�9f�=�hm�#���Zn�WL��E��o8�͗mc<����rK|��PjR�"`'��UV�{�e��<�Uՙol�hRo[���6�ٮf0h�7�Ψ勰��W2[�v�7k�h :IG`���[#q�9w_]]�[�7^��)�V��F�hT7�������W��굌����Ug^���*�����a�:r:k9Aw��:�����ԶE],U���*����܄���M�4�%mj�t�+�\�e��&�cB{���S�j�t�,�k7�Z�$�D4B>|�z�]{��ss.��n� q��ǯ,]�a��h��En"ɫ�c�C�*���M�n�T=��[����`*
X�;)�Ӣ�
{��Aw[b��" l�-�vR�`���?��u�K���>�8鍐�/�Ý��\�׋sK��r�]�(ƶ�4��͙�bl�j%d���B���mEO!'�	I�j�{C._wh�:L�/��� ���շ�4�܉s�|o���/���[� dP�e�4�RЦ�V�z{��"U麜a�hf�UlXB�O5�68�tr��Y��q�3)�&�i����=�
�93�j���u�yX�b��WA{�Y����&�&9Uf��,sͬ�X���K��S՘w�\��}oE�g� ��VwQ"������x���Mc��0�ǘ�n^��^ò�m�֍Z}J�ԋ�����a�[q�yL�j����e��&�҈ue5�Hp6s�:΁W2�kZaaw���ZoBeqW�)���uf���.�h?��ѥ���;XR��ܼ��):en�҂hв�<����˵�PcB[�F)H���Mu�a�*i��xwdW�Yj�y��eBK��਴�Ҹ��k:Y�9��q����K>f�H�!���qY��nLmK�u��'�!Kq���@�F��t�]��X�u�EP�U�`��Q\��آ��0�/*}u��T��;V*�9�}t8���LiP��%�Ή����N��-��1V���sJ+�&.g���$��9�؉��Y{�6u�S��f����
��;�B�YD,��r���νH]w�F�6y�{|�<l
Z�K�uB�Xy5�Ц�c�!�F���VHLb@���C�E�SrSX���2�3[:�u��f�u�J�_1�2WD�0-} ��R��=�_'�����iV6wcQ>:�.Vݴ!nS�I�Ӳ8]�X�|(���&Ԑ<KN��̣XiҊ�ұ��c��K�V�y0]���5��o��� ������ԩuOX�ݥ�M]F���<�ḇ���ܶ�×����7-��#�7]�g�6����l/6�9�ٕxu̩�3�^����]6�NL5��k!i��uJ&�m� +�'8:��F��B�˫�6��(, =�jK��� \j8�b!Z�f�rO�c��Sy�E�lo�1��kW�,g��.g��f:h�d�[�Z �P2���k�0�n���K�&������ڰ��I�ySyW}=���-B��[�73tԙfn��o�ڒ���v:�R�1�d�A��l9�WU�^H�#��6��p��(L��2��^��xMXʂ2�GU�bt��bYq�T�eƇP��a6z[��)��
�Ko�����}�%D7/[o�؛2���x�:s�Y�'Rz@���)��;d ?�՗L[&�Rs
�u+����>������aj��X[M���T�uE��_a�����VS�/�ȹ�}JK���5��0놶^Rǵ�Y��@h�ul[T�U*�`�;zd��`{��l�&������.8��{�X��G���F�K��w�Gh��T��f��^mh�~��-C �syOk�n
1nN�Y�%M������p�+�ZйO��V)�⥶qV�U��a���*,'�|]Nͭ����w��n��ƚsm%k��t�_���V�8M{ϺGJN��r��ۻF�k31��!-d����s5���i�+�0Ֆa�{�ż��Y�t�q
���B0X�M����
�RBG�=���ؖ�h��D���М�遚�66�	�3E�T�ģCH�gWk�qv��=�����]��x[`���8;��b�v>�iZ+8�4{��^,��q�)ǐI��o�097@�dʁ枵6����M�o0,��p��E��m7KyJ�y�`'���Wn�v��WL���&�[u!�M ��|G����^�:���xt<?���v�5�gs(ˠ���-=��t�i`��%w(l�_*Mn�E)���C'���⮘�5��v�f�|�4a��f%�����ɩs�Er[��(U�[���:^�2JkM�F+��3B[�[[��j�m����p.�|I����{�XS3'8]��7S2�W�XN�˶�U��3:ә���U��sf _P��9�e�w]Z��kS��>!�Qڈ�_���9Z�!��X���Dc��9��}�{;�Oi�38�c��v���pg/c�e�2Է��;s�︬�� �$䆮;��������E�[��C�l��������'�&t)�[#�Vы&�I3�F�&��:Q7��Slr��lA�v���oB �^�r�L@�ش��)@�v�FL������0r:r��OI�;ef[���&#�j(+�Z�)�=g���%�cOkC.��j��*9��|�b�N�Z"�$�0vK��d�&�n�K�xB2�4o�$(�d+3\�����G[�WFNY%q�gfY����p��R���-�f-��C��� �È���y�e��IÎ5U�4;�*	dw;K!�]\F��U�ǉVʕk(�>=�V��
!\���V�f�6
%s�j*iu�V#����"��z�;���TR͎�S�Y�p;y�w,�ǝ�^�ǲ�av9�FVrXp����E�%���陘k��8���v�Ԯ���]����́����b�|'''��l��Ҳ���}���s�"E��8�{ëP�99sR��;9"���)���U���XA���dTu�h.�RNw;#�r�k]t�n�g�9W����9��f��\�f.m3m؁r=c]���%���5�&6�.T�G^>Cݛ9�"�e�^_)�@Y�m�0��R��c~�o��	]0e�b�b���7��w��0�j�u��6��.�x�2�R�%;���y_��2��B$�fv�%i�ʴ\�OZv/q��G�X7��ܵ&5Y�S��Ӗ��l��6�bBr�%Yj��Z}x88�#9ڲ����W҇�U�d.�s&$�6x�{5A�n�=d��a�Շ��z����̚0����;	@r,�Sz����!]�U\	dQ�v�`�ϫ\�|�����Vq2�[��.�PL�:�������X���08����J�t��`\��l�P�=��e�Mso�r�,v�.t4���������<�-5;��`�I��C�S�"�"���4k++_Q����(ow5֕� ��x2��B�v�r�1����;��qE�SZ�d��R	�X���(�A�,!�/t:i���APؔ��m+�`��ul�umb����d�8��:��y���V�pf�ì�/2�k���h�7Զ�MR�<��l;N��39��؈fc�qFlC]�н�zdw�s���9���R�v�٠�a囼ݒ��'A�VoXfw;o��āB��F��?%�R�X���R�����2Z�K�C{SU�W{�؆}i0ctYH
���R�WniSa꾤v$4-�6]���۸bޛ��m&���z/�R�h�b$q_>{Q��W������O�>�\uZ/lI�]bF�;W{k��o��(����JT+`��ђ�K���R%
��tsg�����+�fv�����Հ���¤�#��'�֑뭖)1�	��.o2���`�@}�<�0�s�i�8�ygJ��{4_sD�;*$�f�[Ն�i�P�l���|�+.�8vI��}��o��;xM����Q��Z��AS��ʽ"�T'1���ʭ�kPpkȨ,;f�\.Q���w�ظ�!�׃�b�Ɖ��{ ��FN�8����m�Ĕ����:�;��}��
������iYB������+���r;��0oEI��˛ŉ��2Ƹi�5h��1�Bq�MS\Lm��V	�,�&��ގ��� �=�5�;�vQ�T$t���"��z�u���3�,I;�C4Xv\��5�%�3����xS�0��
CHZr7��1�s] 0,��d�����U�s�d&�s�{.��]nT]ْ��XfE�� �*�}9��w�P�(P�|�,2���қ�:���G8�]�)��ۊ��eqn96�0=����	SR�SaWb�Y`���xJ�Ջ�,�)�%&�˭Ȩ��+N>��5�p�����yd4@�f(V�e �e�F��R�M��vl�����u;����;�KS㗉ب��f��g-�/�ϻZ�-�&�K"TCpۭ�.�sbFD��I��-E��s;;xs�Q`z���-���>����Ӛ��э��r�d�X��
ȯ:�Tf��&�N�I�4�S*U�����֭w��ӧD������hI%*���*��d�*K��W{zFR�u6d�����T�u�&$�n�;��A��v�d�ӝԍl3xB�J�ґ:�o��b�V�^W3�/�nS�\����L]�e8b���>oy�6��p�L��R'ܮ��uA��b�4Y`� h�H�]e�b���L7ƨ�m�B��t��o]J�`%�"!��B�W�K�v��Ja�v�2�;CFI1}p\	��2��`�R�����ˢ�*�1I(�yvL An��*�I4ca՟��2�<���%���v[��$z�Cq�!�Q����! ���|�cqo�w��}�����������A@?w��_����S��EE�_����f�'��h?�|��@��w���x�.�u��l�ū:0���T:�'M�D���Ƶ�M�i2�&�U�vz���9&�?Z�	��)�KUYb�.�H{�n���ֹ9�3r>�w\�S�n�9��M�9��M�F�y�{��xnc�;��hml(՛;[p�3)�7'����5c.�G�N_\{�@�j��t!��VBSޥ/�[+��/Wvh���(��»T۾嚦���Hb�r˲ѷC�R[�)Ӷl<�����5�m�=��D���� ]�׌�͜--I$��0�|�;fS�F��[
1ޑQ�Ͳ�c��OU�1w/]Yb����ʙۯV��+Z�L	��ee-������֘=��RƓ�+�;��hv3���
��Y��MI��(���%�/�m����Xv�}�ͮF��D-�e���h^i�Q>&��DM�<���kc� 4v*����(1SV.��j�R���Bbz�����J����w��ܱ���\%��6��#\i�����.��jk���2`�X�rח���w���k|)��X��Z�h�ͅ)���4�;Y6��hj���f	טc����i�2p�6U^��:��K.��I��Z�c)p졓.�p��b\�m��ɸS}JĻ�����l�����땶!�نG�1��7-.H����R��i�앃,�[�����@;]��v��lQk:��4�A"*꣮���ڕ�I�ڤ�;u�k�`������f�A�`膅�k��N\���p0y��c�@���P9�p>ˢj(�"�Y�u'w՘]�Q�M��D�#W]�d����-��쾕I@#��{��-PF��}X�A�RN6wR�4���a��ĩ�:眷�ȵ���;*E(�0��Ш���Uo7\49�4:X|���J亵lO�V@ƳM{��4i�&-�f����]eI`Wg�;l죸+WJ��p>/,��1���;��ҳ̓�acs)�S�h�KE�bM�ea'�5ܬ"��fZ��	uc
�� �f�R��z��KV��S�Sh���h�k
��c��9��05�Z��V��J�+�Ś/�y؝w�N�`�}�3��m1�n��m����#f�pĵkt��iB[��M�5ց�G�;N���X�"��(�ܽM�	
��/f�hH[��-��,���fg>��n�w�e-��L�Y��+4w74�H�uGc�r��%Nr_'�6c�7Xb��W�c��wU�e*�ud!���ƪ�a���,T�5�z��f�ג�#�|��{6�"Ŝ�>�)������Jߣ���@V]7R���E�mWY��O�JX�(Dr�����B;��k��ѯL��fU"3��{��"x]*�k:K�֞b�� ����_8���N[��Ty����j��v\л������f�O�K�&�չ�e��@���!�ݘ^,�.�)d�
�
[��G3���"�x�����וEvI��"�����a��U3����L�6������g���<���n�}�]�+S��}h�g�����#�Ҡ]5a�BKv7���Uz���;v�ٮ��k����Gs�Ӣ9M�u`Q�Yb����u$�^�P�Q	�DP��������ԝ`/��)��D�,��4b��	����=7y�#+��5GX7��n�j�Ns�ԘWԹ'[Y-��tR	�p�U�Vu���ڍMd���� ��dZes��)vncf�Q�*�y��1�<u"��%�%N����B��JP�����2n!}��N8;����2�ζ�ʅd�s���ˣ��ս��e�T�W&�0P���]���R�{9�7����v��\@�Bkxܽ�ЮOz����̆+�܁�u�۲���7���z�M����u���3-�0�+U�|��ǂ+U��u��@�1|����*[�I����<�ƥ�k��_4�.�Ȭ�XFq|���i{Ro>�rM�j;���/,���2�,pw�ǥQ���fl̔m���큗��;�}�xO`|�n�ժ�1mt�2�]�p�մ>�O�-�E[Gt_�+�CT�.�o��YT�s`�R�2o��G�W�Xi�|;�|�Ȧ�}���.�c������5����a�Z�׿�i`�㫑��ls�l��ۆ�0n�~��ܸ1n�AF�
v+�"Z�hc�D�Ǵ�����F�h��:�:S[ͫRГ���t��������H6�I��P�h0�6���]2J(�qu1�C>��&�i'ht��̃Q�*�Q//S�+cy7cAۘ�G�`�- ��Q���ܶ��X��4L��5��=�;�s�Y�w����LY8!R�E�0��о/y\o5]���P��Ϭ�p�APq�∺�[�w�}-�*N<�R�µ��N�=����*�4.:� ���zU�8mV�_ne'�!V_m�#���Hmu����^�apwʸPZe;`�oK�l�r��)۽Ek��p���rqwGn5�L�8d�{����a�F��������Qaִ+J�G6�I88�D�*ZUT�Y�W���O�p.�w!��e�z��t�.�M	��(MC�ٻM)Ny5u/�գIΗ��mɶw�5�D4�2������g%i0P�!����B�f[��x�����,]5��w���/^���Gz*��t���9WL�Ý�gX��!me<�8f����Fs���Ug&X������no:Pݨ�'=�?�����Ω�s7����q[l[R=}s�P�X��5ñ\eM�/2Jy6d��;w%�-vs�7�8���BԨ�nn�ܤ욷�3w�m�d���i:q1T�˚�ח�p���r�>a������BT�a�螝v�����G�:�Cч�]\˲;ru���pA��Y��7w�q2y��7��oi�֦���rS�oWo<`+xXR.��s����������cWWk�k1�ʵ����,���V����i�w���	���|�g����g���]	Y�1�h���S���m�&S�2�;�y���k��Xt(�Q�N�	zO6����
�$�T�
Y��2��M���Aخ���Z���Q��
�p�����k7t��BZom;�ej̙����	A�X��p�A�;�BF��c{!�{�{,�k_��8Y�Zt*S���Tڎ:�����IDeb�29�1��<��qUm�(�N9"��g��t�ZbylVUqӢ�zC왴�U��Lhͬ+m��'���.��Voe�#���K�����Uc^nپO3�K�U����OJ��n�)<��3��mkٙ���q��I��HI�ޝ�3�1���h�ԸI�ykcj�ChI���8I��ǜ���첷z�|����D-��w%d�rc�4�s�xnVP�ٛ��;y�h�01��������i��۽5 �6��P���]�3C��AZ�����Q,a6��K;�+�ɠC���n�`���t-����<l��2��GdZ���J��Z�lg*E��>+
���ֲ\���3a�X��M��jJ}�1kRs�PB��� VRb�5.Ջ1�d��[���I�O
5Y�eP9�s,�"�3�;X��s.�'Lj$�j)�01;o�����˵o�a;�Z��Q��n��vGz.��yI����6�ݥK
m�;KgV�<�g�UL�9�*���2Єw&��[�b��Z�n�6��	$8����Q�^^s���Wrv�{++�Y�R�)�}ܻx�\��tx��r�[-�Ķr��S+nP7- ڣ�wݔ"�˃7 7����.��p�e(�X��K/|4⨄x6���=h�+��3x+k���m��:�;���\̘�>WCk�1fVe[�x�Ρ$+T��'��"JI^K���-k��vyԖa[�{�T�U���3KD�	e���[�▀}�pjڼhX���GGp����TY�9F�:��v��Yi�����Tc��h�2��uk����ۉ�]��2w�sPm�g��`���5�|!�=�T�5u�N���Ķ&+��!<y�Ƚ+3��Ba̕�Pb�0k����R)����4�AɎdU����kp��"5)P�FL&�f3cbtzI�si�thV��ǟ2���o���I��P�.ӭn�®��-�T-�{a:�YJn9۽v�[��L��r>nL|�7�L�B�f��ʄ��a�xEg=9�6���wd=k�v�v��\dr�`�w���8�����1"�>f�`;}S�m�������'^���)����̩wόD1R+�2E�e�q��j�/V:L}���f�5w]�na��y�	��7������(�����MCE��~yY��|�l�L�:i �|Xct�Q=������]���.��.;�ZUh���R5��ؘ�:��Ks_�V�aw#�ˌO*��ifQ��إ���,�Q�{E����*���K��h�o8X*c�\�Fhwk+�/��RΏ��9�-޼,���f�#�m�2���=�РJ�hj89�Y�w��Sv�N�ݽ0��֩�����F"���څv	5�O	j��h[O�Q�7����	�o]uN�k�Ɍ�h��9ɺ{-3Zo8��M8h�
�S�Y�����0J@�tC2�Nn�H)�]X��1�l�J���vv ��z�!E�Y��P�N�λ�t�ʳ��JԽ���J�t���Y�L�+A:/U\����H��H\ڶ*�T$���:�;ʲ���[�z��9�P���8��Q�&��u�Y�@a�wjM(���-��rH���t�b�R!�i)S��k���$�1�C�&a�f��5p ������9�&"���y�>���q�2)�svQŜQa�z�R�$�ĭh5EY���>]L�Wٴ�K� ��1�w9}wS��׵�mFi�̃P�	fīug��,�Ӄ�r��;�"zЭ��H_��hg:��R�>�+��6��;��)���le�/x	4
�l���rZFgI�<��/��ǩe�)���q�����,�j���˚�fV[��;���$�l⌳�����U�tK?+͵:�,:�,N�Sv7��cPN3���q��7��Ҥ��ٟf���i��[l뽤�P�+,�ӆ���RrOD�kr��0��%.��i2�4�Kr�<��+h%�c;:�*���F;�EwW+*�-��ٸ��2Joiژ���07J�3F�J��[�d������n�Ը��\ht���S��
sܤ�T-v�M�.�*5��:�n[u.n\��K�aga=;�<ݵ�guD�f[�]�RƝ�*ί�$���s�;Q��Ș��
޽2�7[�X��8�q�G��%:�!��R���St��F���)kS���wd����-,5�����3L��O/��Ji)�}v�AG*�
�� �����x4�Zی��y�����vd̫2V�qi��ݛ�T�r ��>�3�e`�p��P�q�����-l��2���
���j}
����0R2¼
3,*�����	,�'��V6�Q��T����W�f�;:��P�{����or��@7&��E|��=��u���*��sC4su#,8h��[Ѥ3r����d$fT@�1	Yz��v�ʺW��#b"]�

�A7��Ee�#�\k�G�)-CDc�g~"n��n��*?�v�b���4�wwmp0.�����Y�u�j��2�SB�|�#�^f�Ū�a��чo��_�9@���x-S����+�K����[�U����'
h�5���[*� l,ッ�_wX"�7,^D��L2�K{2�kY��An���Մ�eR�O���h����E���3{9����U�L'RP}��)Ea,�m�{����Uʈl��1j�y�����Ky�Q��W0�I��!��X�t�<	_<����ė��A[�3!`��t�S�;5�������Y�T�9�mF�(5����SI޼�.
ǽ0��5Q�{#���ES.�k�w�[�c��L�-�=-S<�f=�����[�*�!�KB/�9ܵJ
-�ڞ������뙌p���3S����u�!�''Yt!ٯD@��2�c�7��7�H
 �w��n���ʏ��U�������:�*f�e��G:M��Ó���y���v�:�˗�k�t��`;I�L3�LSڌ��5ν'�7B��m��sʶ	�pj�kf[A��ˮ�#�f��C�,��_+�K�&�D�Y��tP�\F!N�S7%M|���"C��1�`1V,W6��tv��ђ�������B��:���,.6�J@X�i��f�� ���sOn�ֵ;uƁX�;��H��d��Ȟ%�����.��,o�Qr�����ER���6�Y\��������Y�IQ+���.��֝�ڝ��3ղ�eI���jY��ov�اSz�R��6��KE��%A�G����ɜ/.;��hV��q�[O��Ӛ����SK�ՇJ�s�����-M���J�A�,�"���'C�}#�Ct�`�9^��Y�;�̛ȇyK2P
qD���1����w��;�QXtܽ}�w�V��aK�뢲�;������xm)�!ΓlL��u۳,p�.�*3 �xN����r� �j�)�v�oeͼ+��R�e�`5��^t.q�/ݲ`)n�T;�����?F�du�kY']�v��0] ���/�j=ݏ>{�p�\�쵗�Cޅ^���y0h���	��cY�66�X�I�iw�zD�F�Mg�����+��\'���Β�c4��b���Ye�Y[�,�iPm��wbr/M�_=�����dU�b��-s����=MBi���U��Ѣ�-���}�;w�Ţ�Fb�����Om��[Zg<i�;��Ճ�?s��۪��W�����������ܿ��?��v{�_������������_�3������#����{�(�U���w�*tk�?N]����u ɓ��[�n�v�7p�[f��ܑ���ָ��d�vSɰ^-���`�o��N[w����W��mS����ky�#��^ш��cv�M�$S]�=��k{q���7d5e+�=�jhLn�S��*��� ���V���wU�Ȥ�^�5*}�&�������ͤ�L�-�i�o�]�OOl$n^� ji�FW�%]vо�d��7��B߯:#)�^#�kUܦ����Ξ	d���K}{�s`G��o�K^�� ��q�RwoaB����3���\ĥ���|����3e��睯��i���efգ-ݍWv�@fv'X�2P�h}����ۙPN!:�]-�3��Na��Wb���S�mlY�j�ܺ�[sO)m��A��[����ɂ�4K=Q��ԨRWz�Z�;'��+Hs�	�����;�����)\-��@.N����=Q��.kG��%<k�օ4|�3n���Xu,1���p�Θ�e���G�m,����q�!ɚ;�3M(�\�N����7\6��������ǝ�C�@a���9���O��ݦ����)Xt}J��I	C^z� N�w�v���*��H0�Vh+j[)No���T��.֋y�}/��;���A8k�E�n8p^q���[�b�c ���f�e2�������"	$�JD�wWZe�1&�bJ�n�h��Rh�SC�]���Zz�(gF�1t��ⓢ����m����E'cyj�5yn6&��yr�ij�����Z��m��m�;�<�;:*-:�l��E��5ݖ�MkE9��A�4���Kc]��3�GN"�����hMD�]�ADCEQ�-h|6Zz1[-&cM��Еmm!�N��sGIA@hb:�֓6���R�C���d8��&ŝ�I֫F�#c$A�B��mV��q]wGG��ǐ�a4�:Ѣ��A��vɤht�n�&�D��Z���--E�h�P���y]�R� h�#Tv��;A�1��L]�GC�^v��c;cc�4�Ht��w���D^F���Ӡ79�GT꒚y�Rt4D��4��#6��j�4�/��~���／>�M꼜������;(��u��p�+6�@I���c���뮔���Ҫ9�>��(۝�P�7o�l�/�/p(���z*�9��󂒳������#�z���^�r��O*q��N�=ў��UE=X7���������L�&��_���/f����>��n�Ț��q��ރ����\r����k� �e�OkwX�g"i�٘�Lak�=u����t� �=���پ^�y����m��9�n�89*�16��{FV3��M�^�0�2�9Q5����o�zo�����bboa��V:�u�W�m/o����.|䫙)�#ّ�xo�W�^��b����X���(���<.zc���g%�V��os��=������{m�uV��.�i���=��9囼R�0V�E���ds���=�T��dq�9~s�dSf�&機����r��A�֏1/���͛�w	�z�Q�5�yz^��ڥߊS�fȢ�RȔf�FsP{��h�`{��<HPlK��hhi�C�]�g7�.��@��-�JJ,OGX�]k�ʺ؎[ʞ�ov�3�2���rc�c[���(��"�ʽ©�IJZ��ݺΫ�p�L�uQ�;���k�{2�l�[�\��Y��[�O���n^}o��Iw��Y��F�"��6�G����Ƭ��oގ���:�?�@}k/�(#7+�>��;��(	��[��'�#p���CK�f�nu^!e���A����OzNw�[���}����ʍ���oj��'9F�����Y�VxaO�7�}l��]�V���M� ��f��2��ԟ�OORuSw��~�~}�q���x$-{;!B��Ԟ�ƨ����Uλ �73xyWp��ޭ����ʻ5v1N6�Odլb���"}�>FK���Tb�.�ԉ�~|}^U��2�^�/�9��ŝ�嫪D���qo�6G(��?z?gh�"Ͻ͹�`�b��I�:3N���UO%��0y���u}�v��F�W�{�Nr��<�k���{���+i��uZ��5_>]��y=�XT������1-V-�
�_8r��e�j����_����#Һ��Ǟo�r�W%Hej
�ٺ#�W_c�j�YƩ��co�&Ņ_'���1�P��`�P,x(l@f����c�Ҹa��JWy$�Pv;P��\�a��j���e�x:��l6�SuX�!������h7�xq����e�>_{��j��:��l�CZ���չ�3zp����	�x{)s��`�==�^˪�#~�w��7!r~C;t$�XO��vc=JeU�x<��3�ޒ����������<K�Y���Q���,�v�B�8j��n�x��ͩS����^�2��#T��yz������𦱾͏=� �8~iOG�=�/)��$��К�G�;�{$]_A�4kޝ:��ycd�dw��[�k0��#��uяvM{�����e5�
f�l�G�)��A������\�r�K�>��l��z��n�{���Th�ߋ�6���N��YS��<�������b��04[>O�oɾ���~�:��O�f�}ၘ���;z>�� ��F���b����7�A�Us�n&�:g����ÌL��'/nI�E�5�mr�){s�S�OW���}/���:/h|pP�@+�l���C���+ 2ރc*;X�)�3f,�A����1�H-�� W2���nv�O�zA�SK��Ņ��v�]G��k������Қ"�� �0��j�KE/��FOs�3�K��i�9ة~9�(t��V���v%������X%=�_���;�y1����93��6��y�#��/�*R��-`��gܥfu��mX~� Ǯ3d�����t�vV�g��˙9m�ߍ�b�2G��Z}�}����du�t����1&��E=��q�w*���=ڋ��.�wM���0+�%�����;>�|(f����`���k��fx�d�W?���@s:}�Q·���By�Joj�����?�9��vn'�n��Y�d��x�����xl��׽⇘��Z��8<���󜳍:��,�I�zT�{G�Gk�q��%��=����c�"4�lmm=��!���-��X��k��&缍w�!=�l��������U1��Z̌�1�o�>���8g� 驓cL������x��w�ͷ��y���6M�s��`���*��gu�k�rq���kx�To��W��Q.;��͙5��hN��^�ab�#.P���(��Ѭ/�Z�<Au��!ه�ڶ"������;��;V��N̹���JqY/"y{��w�&��J�&u�Ji����.��)Վ�+Kx��ѻ���� qg��C+g��g���u�����),����nC��w��s�U������ F�.�w�ӆ�d�ܡ�[7���]��|z�{�N�|�^º`0eg�o٦yR��N<��D(9�9��EM�݃ㅺG?�(X&���v�ŕf/��\ޱ���{�{<�}�75y�y1���h�6����A�j�g뽺~��EZT^�8���7�~ù��ja��{����d�x�e�̙m�ؖΜ�b�K����=1�5���[��<�LO<y�W�Q���_?��܍�J��l�B���������IBlz�V�~�b��ʞ6�p@:�����ݔ뛼����s�laf�����љ�A����2Zp/#3������l�����/\��v���RŖxʂ?Oll׽�Kkǳ]_9k��$K�����u�/�?-��MӥG��I��2�:���ؔhBU'EޑU�{w'c���!�-�]���ak����Χ�V�:qC7i��t��M灕-{Y>���Ȇ�^����.��Z��T�g+��i�ՠ�U�t�c�n�Q��2���%�C1Ƕ��6�L�Ĩ������� �����ݽ��[����?EsxE`W]����/ޫ��l��U=�|��}Ry��$�?{^ڻ��;�+��'^gfڔb�Ql�'�%z��m`��������Ec<wNXs����gdt�@ȝe��o��L��;ێmf?maմݤ���y�{]f	ׯ֥/�Y�6_��.��^)F��O����߭znS3hﲞ:��ln���piv���uw�����lݓj��)W���^�2Z۶;�K�zv��4�����4|����.��'��������:�λp�1uo�GU(��QU�'�1�fu��{��A����}�ዩ���Y�S;}�z��uyޟ:����kUBd��^��y�'�^K�WY���(<�<�3���T>�3q�[�9�`���􂷇�����KaM3�F��)�Jl[���|l��J�Ӆ�!�U�K��P��7s�r�f�i�"O~;��@J�i�T����Ǉ޻��s���S�%%��1v^���*�B�A$��qhE7,���|&Q��B|r0i�r�n�*7���Vt���l��P~FK��wk���׸)>uGy{U�>�i9�����6k�]x���"��﫽�߷�u�����Pj��ݵ���^+�3ѿw�$���ʙ<��w��(���fZ���Y�7�������O��=�2ϫ҇E/~s�~����=ސ��-��Z�#bӾ����Wj�����{dr���=�&�JK�E��Oޕ==<6$}����}3�r����s��x������:��X#ڬ�����?$0�8�-��'���ݯ�0v9���ϻ�B�ʸ��ok3�uNٱo���𳽩W/V߆6��*̸�V`�Oi;�v��S��f����zDF��8������\�I�Ş�z'�U��{��]e���7u>r�^{ʖ'�{�U}^�~��f]��0b��lv'���g3��W���_=9R��=�W��5�vV2�&~/;�d��c�^�/���*ّ�ά�qKӏb�cP�hh��IhMJuau��^T-����؋��n�l�!2��,��;2�ee����7�w��6��y�CV+� �z�]]:���1\��b��ӕ;9j�1��Գ0kK�pU�t��<G�ڬ�Q-5��,�ڙ�nu\�^� {��~7ϙ��(�����eI�F"�SfS�ܕ����g�ٯr���j�ו�u�`8����,x�F�g� w?���w7䜵�ѩ�9Sӗ���X�
����m��h�4��"��<��ӻ�x�޸�z(�����=�z����o�/���0(N�$���u�l�y�T1�[�A��L�Y�ޤ�.W�{ ����W?-��61��풻�ϛ���$/��?gMdOU[�ݮH��3Ǿoޝ�������<�uy�]�^�ny�w2�>�2���d�\�[(}��s̓��z3U=�:��̡��2I�1^�{�����Y�E^��NP�������a��Ǟ��y�x��2��Ǜ�˻�VO7�:�w�$�ݍw{9q� �P������A{_%��A����^ɓL=]��y�^~���aRZ|ed�oJ��i2w�v!�P{�F��"u����}j9ǹ�ۗ�È��u�5��`�W�q@��j�l�K�
���Ï �AjX�47��N�I��S�$:v�̚�6����� �eR�I0:�Y�of��O��~���w���&���205�C��{uȓ�M�yS��a�y�;��~����OH��k���(p���c1�&�v�������<��Y�Ӯ6���_+�u���g��6�����y���6��i��^��];1�Ի���fI�ѝ�;k��Y�V5��Pf�����J<�~_9t��޼��K����|�T�nq��#ؽΒ�Ϣ�d\羛�~��~�h�a�ǝ���@92+c�3��&[8�"��T՜��������?Ow��U�^Z�A0sL��3��,	���(�4Pݱ��4�#4��4#ǩ����XTa��u����N�"�ױ���g�̻�%�A�ӕ��^�Ǿ��Y,{��k�3�����z�5��t=��?$�FO|5�Tb��խ^�,u7��?v{���ۆ׺�8�}h27��.��^��/�F�x9��Bl�Ȅ�j�Duf��pw:��+!VvdՠҫgYd3���VW�����^c�xV���a�}���+Ӻ��[x��X62wTnJ�㽶*Ay��$�I�P5��vv���;�\�&`S�Ҽ*�����T����p;�9�O�M��||�U��Ⴙ=�~�)^;<l�=�{P� '*�KԨ���#u��ۃuP��.���"��^ΰ�3�����G��fm?ip���{y���Qyl�-Ԟj�9�Ax߼�J���s%��k��2n��s� 1��7��I��o�j:�$tz�57�m7����έ��n�Q�`vgCO)���y�����[�������3ŌKl���tsܦ��j�P6�_��ƞ�L��U���y�|�51�^�m��ǳdG5��a��׳�|6�n�1�/3����ď��Ox{���O$b���ޫr�8+�=���յ���;G3�Z�4���R?7�r����%l��Y(h!Oz�*��l�nmO��N]/I�S3�IK[�1T�`�w�S�`6�P{����7��ɹ&��u�K*Ǫ*1��3����~����|||}��>�����J�/RĮ��RY�&Pz��R�[�(�D��OoR1ǂ��K��Q���°K:��ޛ���
v/��,�ݎ:��3�29.��	��t�pr2��I`i�$��9MOFE����)�(L(c�˯�|�bn�U�2*M�p�,v�7oC���B�+�0��Gewk�y�ޜ�ք��BeVl3
<�^�u�zNX�(�l���6�Y�vr������F�L����M���bҾ�n�V�( �[�Nui�z�!�_wH�V��t��Y�*Bj0����N�3�<�ѰY�d�{4��W�Gd��^M9�zk\3:�f��Y�+���I��,s29*Qv+G"��f=�լpG�h�u��+�>s�����u��r��Zg;�ͫ����8�14�[qL��L�FMu�b3��S�D.������	����lӗ_+�����4�����p�ùT��]E��AFƸ�\�)CO��5X�g��u���V��d�i-g=�Cq�rń�fi�{�r�1sM���}�|���xFN�5�P:ʐ�b��ێ��\���Ǘ|��N�� F�d&���,i���jg7TǇ^kՃוU�s[�b
unq�̹��I�Uo}��m
�x�
��W�R`ǢN]�}�Mh2�]�T�+u(r���5Y�de-_7�7�mj7��I���H-�b����g���jwf��CoK�Xt0�;�X��gCw@�
::�36����/lH��0�������:r�Jdƣ	�S��b(0I�����ӥh~�謕�Z�Y��P���m��4:�u�H���9(ɳnżF�u�4����m\��s���JU�w�aS��1
Ov���[\�FԦ�{�9��1W�x2;�Vs��A�3#��f��n1S.v32�+ٶ�ѧ݃!TEed���L�)[Ȫ$�Q��E�F�.j^X5+�V�����mV��*��㥊Y��Ź�l��&�dW��9ޱ)E�D�C������F��˫�:�
*ֳn1*�&�i��@sy��Z���%��k�j�n�����Zh��]��<��r�{TlC�x��n��:�4i�x0��#�#M䶏9R��ժ��=��Ȍ�5ֺ�X��{�Z��>}��vvNZ�k��ق�֬�	���=�lu�e�=��'ҹ�������Lμ̐�
LؚB@اִ��x��V� h5�M��6�zp=k>Sx���{>����QZ��흱@WT� q)}�Q�Y��Ө`Ưx[�:c��`��u0q�]����Tj���c+�pZ��(�o���p�]�2p>�	Xn͡9� �h�(���յC_cСn���lI�qM՘4+��hӘ+vR�lG��4w d%������ㆮ��W����͙�m�i�/�-��6�Nő>��T�;d�t��{���}��f�:����r,3�7�Zwׅ�%5����5�-��yn��l��̚�u�7eӣDF��\G8�)�h�F�m���5Db�b6��Ӣ�ƃ� ��cy���m�Z�<�U^m���v
;�yܛ�^X��|�C���j|�(j��y�L�
:�c�˷=;{�m�����,绸<���̇O������Q�m�y5�qDG0u�ݲv��hב��Ww]j(
po�n�m��v���[�7i��ɰb:(���Q(G��m/�3���܄�"(&�DQ���AY(�lk7��m�=�ӝ�'�@y�N*.1��N���8�y>v<��xy�S�מk���q=s�q�gv��b�[���=t[E��;�$�̯�&�a����#�D�����k�iӢ�|��k��n�u�m]�.��cϟ;����4��cwť���h��pq�h�|�^_'ɼ�5�+��kn��2C�c����>xmyq!�u�km�u�����yگ����O� ��ں�8�o�m��<�:<����m=:>v:s�!�Y��xZ����<��ض�6������G坵lG��]��חm�'M��و�$��Th���Р	7_g�=�5J��M�)-�5���� U��zA%[�nS=[]w�-f	{^�[N�|m�<���44ޯ��sѢ��2e��b�{MW���E2.��9������&P��Ll$��b��Xo���0�b+y>^�o`p�v08k�|��^}۶��� ��1̂�D@��M�>�t}�/l����QS-Y�t�*1A,�.*�.#Ȥa���^����WsR�n�h�
�hr�a��'3�v��x�����,^ǲ`�L�Y���.фc�jq�Ϯ�|r�D�^[��oW���w�ڛ�U��q���F2���v.���nb�ݑ|��ʃY�/}��FE0Yg�t!<����Љ�O51�s4�G	�G���Y ����bٖ��+�=L���X-x&�C�k�y�d�A��B�Μ����*3̓RƆ2<u���<�)9�1H���S��]�}5�9���/�)O�'�^>�M�FY�`l�U�\O����:�0f�V�hХ�2���Qi��T/hU�5�q��q��.f�9[��!�osQ�1��Ɂ}�-�=.�k��#ױ@��Ji��EEyDQ}�*�uڰ��1���Oӻl���ꁟ||���!�Wܙ��4o��C+K�yz���.,�31o=�7���W�
=�iΖ�p:������̆.�Ћ�v����8�!6���0�?�<$6��e���w���jļj�e����w|j��=})0���rwӂ<3v���F
X��铚�Pl���E�㙧�2�(�S��W9d���dYS0�MG:
a���p����L�A���*@M�jA��$�XG����* '˽b���f�� ޞ��,����z��j�{2o��w5�xw�qہ?�W��]d�p�����L�^ %�oc?{2�Ɯ��[�gp���c f��rT�m��:,�K#���]���\�����ð�3;}�z�{jFƎs*��f]Uf�w�\�,�����z���#�)�7�����K`_P�Uj��<	x�� ��w��[6cv�R������yO����>����i��vx�m���7���qS4��b�+����tH�vFJf��Kk��1�;Eq�0fAv�c��'���c�d�~�b���E�u���x�:��\éQ|�C�D��ԟ�5E���Q������l5��
j��mU��5Q;5���:���o�a^R�7*�2�V�O�s`�CT��"�0f�P
۳[��Ŋk7�=�҅���`yϬ9�2)�jvq׊,�b���ޏlG����+MMN
K5gk�G�#�*��5�������W<��J�V�*����-��æ�(�CdT,�wr��<�D�^`R	����`��3�]���ˡԫO��ίwkqV�񞪌�z��:��ԥ]8����_^�6һ�޺kJ�YU�r]��I���g[%H�x�9��(�C��qft45L,�(1�k[�8���!�F׹�ܛ�+b�?[�G��Ud"�2c[�vT����Й��E�;$Vh	V��]h���^�������3r�S��܅��Pe᪃��4�j����w&z�3[u�i��^�-R
��-66��>UU[����n�rN�k�m���������\�]���f�\v�[@鍙�qřz�ãȘ�J}�]r�-���:.�&�3��+�A���l�B*���� Eu�V�3up;Rm��LRW(4�)�9�y�Y�ђ̔,>igO�ɋ|��,\0{=@���
���N�����|�|�}�<����U� q�mW0(�e���|͕��yj(��	���>��yI:R�p{8�)����OT������liJ�}��N��qiG0X����^yn=ȃ�������3CSx^��\�0��s�����<=-��i�(1Pm@���r�bNC�ͷJ�n���a%��ǰx�7�z<]�;��zC�&־�\�7��J��3���aU*�b���6�.}[_c�@�O�?�g�'|�G�_z&�3ɓ����Ƃ�ޯ=�Ҙ^�I�]&�e�4��E��iFM��ԍէ{��S8ѽrT��a�V��X�`7C�s�,���li�l�hLPU ���s��R��K��W;��n��8����ZT���^��Tm��w;V4�^�̊K��u[�{~ԫ���:����;��:�μ1ȵ �!
=P	R��=,��v7���G�������cM��W�����R�"���2
D�`�y���C[Cr�#ڢ��;G�)�4S�Fӻ'4 �."d�z��ի�&sUn�����l(l̙+
 ~	B��H��U����aq[Ǯz7�M��ݲ�f�E�dx�@�Rnh���n�)�v�k`�!4H�#��WB���mK�>���&��\e_[�����{L��	�B<R��[d�s�(���l�Sb�Ty���W-#Hhӫx��;P��f)���h�w�5'�7f�!��Iۘ[U�n��N�}�z���f]�����-oL�ǯP�f�s`P��&c���Th��4ܻe	��&E�����''�����%`m5�t�-���%:aeT����[mxr���u�Sd�u��@�����c�Z�_�j���:����4`rܼ3d�0�b��*peG"��8����%����|@��w�FQ~������y3hWZ
XL�-ۜ�D��b�a�Ľ�Ur{
 �G<�p���˙��gD�>Ygq�.��]	�3m�8�v�t�Hz�U����_���jݲM80���}�%�@�,�-�v�e�\΍�O2��2��7��5�˂.�$��mvtS:g_8�\:��o�;�r������A��c[a���t�r�/�z��u��j��M_���{���tָ5/�DFzP;S2/pf�mX)�V�����"I���eu��{+D��x���E�T����4��S����E9|�"�N�ؐ'0�+(!u���۶ن�3M����)(��fķm�#x�;<�����C��o�+�@��l�|	�{z�]�s�ҤcgA���`{k<�^�PyОt?A�T)x����$N����{�FXl�6��q�_Q��)�
ʇ�U�h<�dckP��z��4Pj�\�7�!�Ց>�w!��E�18�o6��R��3����gy�"r�C�s�F�ȏP>c�W�������Ad�p�����z�l��D:~)��< �g�����t����mq�WWU#7���y���V3^Ob�L��͙z�d�@6�j�1�U�k�G$�.�͐�Av����zY�c�t����5�F�9덎��eL���ˤ�@��xۑ���ӻƙ&��|ǟ9R.�d�k�L/ ޡ˲�̻X��ڰkK>��%��0C&X��&�� _r��T�0�e�w��@������_����Ǧv1�D���A��}5�@���r,�j{=�k���ٝO���^�GN�ޢ�*+�3O�p���#s1�i���eQ[��q�A�'V�0p��m��.���X.u�Ԥ�-�����+h�8Q-�vrv��ɢ�.�0RR���/�-��U�ûW�P^��tĜ{�_:/����Z��r�E٪d�9�&
�ō������m�p���1�fey2��lKE������<ÝB.;�%Q��
�O�T������-�r#���#���{6��h�_����C���� �
��x�s�o`?�:���y*-a�T_�����A����"n�v�fslԅ�;�#��u���Tx��'�*x0Zg��(���Z)�w�B���gDli_k��?����G�({�e�49%��#L_l�}�^	��H�s�k1���3��3���tЅ����O�M
}
2X�6'��K/��$v�z��G��'y��VPpmI���te���軓P�3e5�h(�,�\�/�X>�b0�6��X�%A�2���>�/ܥ��m� %�a�Ǣ�:x�� ��N741�ֺC陝|�r�Km�Lrw�E�+D���1^rI���UƉ�3����t{w�_nH��ӽ2Xlb�9J����P��
f;0`�Xl��<��]�<�A�Zk��V�X���6�F������Z�����S?�&���ų���S�Ax16��9]�=�l��Fvezgcc��ϲ�4	�N״��T��}��h���?s��~��r��	�;x�ޕ.� u��wBi�n�Y�)�Ƕ�iǓ��2y��q�m��m����.����?���"��",C��K<ɰ��>J��`���|3~i�)N��ܞ�[G��5خù5Z����q��Ɍ,��^y�j�H0ˢ�S����c1��5KE�#-4J`�.�)����tթ��*v��ɘ3X�Ü�S�P�*[Y&E�jע=oe�Kië���f}u�w���V��ڝ������F��n8�Y�Ҙ'0Ҟt�%rӔڧH�Yp\�M�8��xy����;�׫Ƚ��= +�~�s�̷w�#npn�t(n렸��<���Y"�VT��Bswe�k�4ۙ㘫\brHh�r7d=gP{�-��?�-Q���ʢ�ޛ�brX�4U���]��K�~�0To���Э��W*_�.C.��CG���m��h�[b�b��R��"�i��yy��v��{!�u��zfG\��	�3�_�P���,}���J!��oj���
K���Fv�����#L�c�Wᯣ%(XZY�9� �A66�t����UMչ�o��ס�'��%�0��Vq�$Q�Z���MG|_C='��rA������Db��g�vWV��X]��xϚS�nk��n��zkw
UPk_��Uݥp_�\��P�����)iʥ�e2��v�\*�t�L�`u9��$DK7�*���2�Buk�/��5go�*+5H��s�Xu̮$����	I�so�=��SW��w~���	���s���F�\.���3<T�q���OVc��ZRZ��Q�hnW�/Aj�0Z�ç�@a;�l�A�����.�Q�0���W��K]%���l���_�S�(���}��PôM�20Kg=��i,g�	v�v.��v8+f�B;*tRW{�=�Qy{)a�����s�|?T�Kw���/X���0N�@���ށ�y�#���E�q��Snң&���ϔ�Mܧ�D!�Y���;P*�5˖wY�׷_�z	_f�%	�����n��%{xW�-_��b�Kr�����g��:�xA��: �綾�ѭ_l�'+Ә�a��q|��ۼ�}�4��s�Ê�F��WV�K;M�0��hr&�j�H*��_��(P�.������oȏ�F�s8�+�_��a�6+�-�9U~�͌8�M�ؙ͛b���jR0�/'���߰�?���ڃ�%���VX]��^㩞�{�9R6'���8ʬc)��ط���m��Gj#����}�fIsB�Zs�ݘ2�Pm�f�����kZ���z�ۯ%� _���!8�o�v����HB%]Z�eo6����gg$�R�ҥڶ���)̜�e�S��h�Co��Ё��d�\��gb�N��N�J�J{�%ڼE��m3J�ˢվf�T�pۗ���gQA� ��j��\x�Dv��� ����#-�aCL�e�⪙84����l$���/!��y���l��7OW,�ذ��t!�.�p�ך:J�1~}��?�&y]c�}(���kz:6�!-eV��L���j\�O
�s!�욀�#��d���ć��\Y=<����tZ:.(Vpcą��v�9��"�����K�4�Z�������;k��lK)�櫖�r#|	U�ʈH�d�GOEtL�^�O�?���� ��&�/���k3�l�An�/��������Q�Fz�)q0����a!;�2x�3���X��/̱�m�`5yoRcAa�:�*?>�/�Ltt�n�=�p�m�8՚S���U�\�#ٮX�Z�3R3:ċ�bL0nc1Z��l+���v�9쥚�̠� ��(Ǻ4	�q�8�	�e���=�A���x��w���w"+-�U��iXv��P39��*y�	�����_���,y��T8�"K�ņv
{�u��fv���
;2Qh�c�q
��U�����d��v��L�`1�[h"E�唫�C�p�2�@鋔q��X���eN���}�Ŋ�lo2��)X�(nxT�]ݐR�]r=�Albڧ��w���o�����4zl���#�,w{yq:3vHD�ds�I��:��΀�jޗX%�-�]�.�� �Ty�q��Yr��k�nW������^t���A����iię�U�3��ʥ<>?���7���~"�x{�v5L��H2��܆)f�7��<�n�=zw�^u��4�.z��{��&��l�?@p����Ȭu��fV&>Ҕ/����Q"�زHkF]�D<H�8yCT��4����̑��̪}�ٜ���AJ^<6��k��M!\,YZ[T�bJq����0�E�׏Tv�Y�e�q��Ƕ�r����wk�����!��׻�QH�ފEag�J+MS(S���y;��'[O[OV�mj�����h:�"��n��\�èE����TZ~9�T"�T�Wj��
fZt���9J�s��)c��X��θG���9G@�ʽ�W%%��\c�"v�L�F#�º���lN��\���R������]aq�4H!��Jam/ۓ̻)��&�'{L�ε�Nb�J�s���ء�����X���$�+H���hzԘtw����Fr�u&��h&x;��c|���5	�=���Ǐ��}��@w��x~���~"R~�~������O��~�z�^�����������&��p������C[_�������j٢b|�C�b���u���/�J^T/a�e�ˮ�**�0e�Uw���'�4�-�;�]�9nh���wj2��+,��]Q�ӕ�.[�qHd�BmM��L�Lt���;�)����t�W�ШV���#6��ݼ��yw���x�d���3��u��OX��N��{�}�H8I�[$�:s}wz�x��h1.Y�]ǡ�j��1]hc��M��ZX������Eɮ���8ya&���.�Z���Mkؽ���\�6����$4Ձf
Wx�!�X���]�l<���F̲1lT�Nwg �	7�����pft�!H1b�6Z����+^qvfO���î��R��ɠ�D*f8����^G-�����L0��]Q�k�ʻI�VA�����l�S�u�`I��\�ha9�wV�N�Kku�� ��b��M7SN��=��]�kl�5c!����7���Ӯ�t�VP
|��9��Y�2aj�[w!3�+ܛo�h�cs�R`��.ԝ��e�� �t��c�;���w�fn섎ܕ�
������Wi�#3�J��;�|8/������e���:�LUj�J�j�&��灁Á
��>hv�w>�N�!���h���8Ҙ���{a�x3�	1�v&&�oCѦ��QAe�[6�v�6�6Py�8���PMhӫ{3�;V$�t�ҘN�<M��l#���n���H��oC0�ik�WY�*�5}��ĺ	�nJB�Q{��IM!1~���D���M_SF��m���53�����Dv��#�jNWZ)���=�#�yҊ��mnPc���]p���(��r�I�����SV�E��q�a�n���ʅI�@�n�LB[KZ��W�]h�"���Z�;\����FEv����4L��ݡ�J�F�	?�Eb�s�l�Uy�@��&����i\ƆX[ٸ�5�{ע3���x�j�h����s����p}��8�����/(`�Neoik�Y���$����S�J:;iƅ�%JY)t���m�9u#�7�2�gLPfەm
o�m�or�Oi �閆�o��p[S�(>��$r��5l�}��h��\�̝��� m�a�:�\����J
��ۤ���C�%�쵪�p8a��p�;���4q��`tW�-�ȓ��c��|v���cWw���Zƃ�G81�u4-�	�^1��u=��(Ʈ����ors�����S;�8�n��v�Bҗ
�I�
�N���[�n�8�Nh�=��^Dy��:]��%���:�[0'\����8zԙK �%ʱa��(�Ʃ�@�-�����d�Wĸ��)r��D]8�+kt�oe�(�:UkP��D��˙̽�
���c@Ն)�'LsW�ĚB���<u�8�ޒ'Y��Sǧ`Z]�Lǃ^�U%���8��s���O���Ye!�P�0tV]Fڥװ���ƝwVh���rBJM
(AEF?�A2�@ �U��ă�;j���QUA���^]�j1�kME^v�O�[���-�GC�5�yxGl��yq�61�O��zt8����K���m�V�+���u�O�֨�y!y� 5��퍌������Q=���`�y����F�Z���ݨ,[M���l�4֍&�GES�O#��u�;�"���
������&��F�h��-���4��iƷG˼����F5clh���;a�E�I�y�9�4Sl۴b�]A��-ۣ�0Mh�l�6��W����HDˍ ��T�0�*0Hg�E$v�Έ�����1A��ݍF-���4�AmZ#b�����v84m�m;�v�փ��[���kF����C���F�UlQM[J5�X5��i��1�6�D'X�&����y��iאv�W��^vzt�І&��V>���w�æ�匝1Md��ѭ鋕�h�x5N�1�@�w*���F q�Yr�ne7X���V3�����2���W�U}Pک��A�r�?1����7��Z���Pl�kQ��4�<jWD薾q`�X:�2�u�W<���M�.��(��Zm��Y���ƇX��8Ԍ�b-t��3:��aǳ�iW5q���+����^�`[�3�P�ݣ��%�9��a�T9�9�;��'�i۔2���!d���7���\G|�r5�o�R`�? �z���!�. �ۙ�L0w	�i�1�ռ,'���Ҹ�r�B�ބBw��PLMPg�9߾�D����+���-5�8otF$D����be��A�$�2ڙ�Se�D�-��{8k���B/�bC����F�7��yK�-bn��^���)�9K_�f�"Sb�$��	��N<0��Z�ӕS�7n(��TE��˨T�.b��(.SZ��2��k����ʱ�7v�J|0���V��.b	�hR����fY?"a� �P��PX{�Qڄ�Ͳ�@�-%��]9p�jE�[�.���vy������ja`}D?�BZ�,V�Z|o����O �ј�x8m��
�E����8����w�\vl�U��R�zEwB���I�n>�+�Z��iVj)�l%Gx:���Z����Tɴ�:^�_l���j��e+�ľ}���i��y�v�X�'�Ѽa�ѵ��[Mp&Z����U���y0 �ىI�X���>F|�����լ�c��بbԅhP�}*���՛� v���g�!A��Osf�R�-*�^��9H��ө?�ZW]6Tt]�ΝFK��g1�V�M��2�%ɗ����vE2p%9��;&	�LS�QR�Ph�Z��&������a�Nv�L����z��	x�50qz��#�TP��']��F�����u��hh��� ���k
��H+�KX'B�hwӢ}2e1��u�G�UW���������{k�&Ǎa]و6����l0��\�zنp-�,��|�>�|G�ӑAK�p�nwr�Ւ�brD(
�.8kE��x`amӦI������=�`��oAvF󱑎�G��
�x	�7�O�'��4�\9�-�e�
o�^�ַ��gנj����h#����r0���|����[Z)Iu��32+�oζ��n����{J%�+���9�xn�j9L�'�+K�����ٲ��G�zw�I�o��^�O��{��X���e��o��{���`܌
�`ܢ��{1nY����@P�Y��ʥYc�%�[�E��~�,�Vih�;:��*D2N���yQ�b���>I�k'�S���R���`��g�������[&n7Դe����kU��A�������U�&��:�F*�n������:�.�;���ǎ�9c��,�V+�2�=�"��ﾪ�����a�7�����3���,*��۟�$�8���}�+���xz�n�lм�������$It�o�9W��춥|hm#��b��ԐѰ�^��F���m���U#��L��f�1�T
�Z5�/en��y�B[o�Dې}��f�ҕ�;,�f�[�f����v�q;��ٙT�=ۼn�S���PL��zZ��j��J�Zy�d�1F�Zd��ȠF�2��o��`8#qk���V����|��t�پ����XJ����sT�mW6O(�����yl8ͭ��x���V8�r�~���ҩ�1)�jnS7m�*��z��b�9S�V-�T��P��Gl&~�#DƳ�ٷd�����i�TVCyDR~k��Q���W3�aN�d�*��R�(g��"�1�S�m#�S��m�.=��Y�U���_l���x�}Z!X���D����;<hyrI��h���P��q���L@��S��h9�����ٻ�1+�J~�D{���P[�v��;���txl1�L�y�>�=��-���N�[�Y��Q�))�&�d�X���*Z0�TܛN�:۱z.S�DM2ۥ����ҩL�μ����"aJU�WT��'Rܾ8;2���bIm��t�9��y��W��'��9Fp�;���pS�e-fT��K�̪�z�jؐL������zGf�%�����ԕc_jT[�Ah�-W��B3:�H�v4a���Ƅ@և�!���>`�p��#Z{i���SAwM���t�j8�0��v3�=�d�x��q-W�[e{����ZX��2�"_yf�L� �	���n�����;c�G�t���nk&gK���4�.r)�&4p�Φ�,�K�r���`�q��aQ�w�.q����K��n�[i�u��@���5;M�i@Z����6��ʀ��L�*�3?O��T%<>���]�����.ӓYWux�˩�DG(���5lT!�邍�L��Y��a�6�M".9 �&��r���㍚��M+�E��_�����>�#��>�%Q"�d���ON��$�sv`�4P܊U���%-�'&됖Rx�E�H�ЫZ���%[�C,���B��\&��S�� ����7x�wt��u^��%�8�Z[��o#,��_��n����ד�	jԧ1�h��v���R��{�pZq�U[���yz��M�Jɷ�
�y���(��bUw>���q�x��+)���O�-�!�P���$���J:X�X4����OT 7sy
�[��\�����__T)Q����]/r�l�w��E�oO�4۔ܩM����6�f`o!�:���j�Lce��̺��Tl���RMCz���RʕO��-��\�f��(�5O�<<<��3�Kreׯ�̧����c��9/�u�s��$AM>�0�����/��*����b�+t�򝞗�EȎ݄3.��s��hzX��_�]h�v�VϘ;�n���K�a�AJ����j��=�wv�츸b���$�Qu�'�r1}1���xLwx��ZC��j]�+�,�&��+�}����g|*	�Y�E5�6�Y�M	�0Yb1>�B%�9�3<�	�`���e��w:C&y{FZ#�jL��ޙfw���V�AFidg�=�x᭘�ψ���r���3��!8���6�8�,�w��>	�pp�|�!<hu�H��FE4��������N��R�-�p�]�6��X�W�=�<x.��4�)?`�������s�װu���A`�5���{+_�?n%��&��:z�!C���Q��=L7���������NR��ϗ,��b�X�����}x��;����S�rXs֓:�
a�P����::��.ц�3�B�`�g1�6p��em�Tq��KV:�yW"��{�h�$�2����Z���SJ����3<����-\5�<��N�;�Yy҈
j]�[��
bέ��]���,u��P������e��U�u���\�����םO:.R>9�HhSۅᤩ�rs5����9Y�v3b����Z�25�2�'J��������x�x+��Uw.8��4�aY��S޸���M��Kн���(A��H���8���;�-Fu���Z�����jzE;ڨ�����)��ꕯc:	��y��\���"��ig��|
ãcvf��X^Wp\ڗ#b�,itO�93,���\>��xB��Ai��v�SF�0K��!��_V��y�&�w�/���*܌�/C���"��
LZ(�ӊpp.X���0�H�Odo`3L*�hA�����ț�^=Y�6�ml�{\����d�6oØ,����9]%s^�mtS�!A���i�2Kۙ�]bx�<��O�?
��clOLx�r㔊X{쎁�B_)�m�����D�Ӯ�����%�݅�<�L	�LS��,y<�^JV��Q�ұ�U�I�Hժn0y�㹲��y�+�;��.!1�8-���y�<��dчf�s(�dq���!���_�l�n�(86(q���6Z�蘇H�6���8Ъ�Jn�O�H��en[K��f<�5Ay�/y��W�x���E�0S�Ϟ �=L��{cg���,�X�B�Qg���g5blt]Ğs��B�^�]�ul����D1SEJ�ǎ�Αe]��2���ܠu��v5��VD�v	��Pw�$M��-=��W�U������A7lP��C�Rc9L��2��;f]%�H?�Y�#�����V�l������������ �=�0����+�3:q��FEz��5*e���6n!��1vF��]��d1�}AF-S��OH�D�t�E����ǲ,4�s�-�{�#�9�.Ƈ@f�����}:/�N��uO�M�Uo� ����=�խ@td���Ý����v�9d��1�\T�� Ν�r���ڙ9"�i�Gn-�^)��ZQo�N���1�0< �����'����Fx��'ۯPId��[[�h�2�����Ф<P�K;���49����/]oVlm�D�#ՏÜ�2N�e��.W�^�d��n�=�`�eg����H�i�p��W�Vk���U�T�=aF*��j��\+T�I�5��eB���Hu�O�T�ٯ6,<&}j���i������+��[���nTilC.��5\b;o0��JMc_��d��M2��6=���d�1�6J�>�sf��Za躚:/p�LK.��Rh��;������ds��6�mYX¬�љ.�xQ�W�mL����"z*���r�K�]���	�����z��"U"�ħL,x����i\���:���fM��^]�m�_K�K�нfP�G>�/y����5�/�V�lchVf@w��n�1ۃ(�T =��FN�
}�{0�b�5ۨ����|��$2��H9���#k�7e`�=��.�40E�p���ƭo�3ڭRqU�q��;�&)�o��5��x{ɽ�<�< ��	����&�>(m����h�i�R�BH��Y4��}}��8�RSߔE'�x��F�U�Ü��eX�屸xTs��\�u~)�����i|���ϸtϮW���OCQ�yl�Wmo1�7/��a^[����l�20_���s������n�/��(oC���N��@ԫŤf��v�*�؞�d(�(Q��c���\G|�hLh'��G��Gx�,��鏦}{Z����e�|~��|����t���9��R�3T��Z�W������Q��aՏG,�Y�!�̚ވm�{����і�:cca�O�:p�a3��z�H}�&k��3�j5N�s
Tx��F1���Bmy@D6<=�a0�:	0�v�2;U,cXsp�.'K���.�iRZ"<٦Wt;w��mT
"��/���?`����|��;6�A� �;N��\��U�g��3�k@�)�BE�����n�=��}`��7��z��M�ǣL~�э/�;��^��1C � ��(q�hr��6%fX�TcL�jX�4�lG�)������*r+�T�`�5�rn�=��F0ȢK9�%KlR�DeQ��h�3���4冘֔��۔$;G����yl��A#|��J�J-Z��9o�b�B�	r�@��m��H!D��G[���"��N��W�.[�8�Ěz���N��&�����D��A
~�}}���~D%�ѝ!��B�-�N0�މ��,�(��0ϒ��u�$��ON��$�g7dC@:�\bf�M��y:�S�4���l�Oʳ�Ҙ ���i,�^哂���-���V����nv7��U��r1	�c`�4����n�/�m�^Q\p.�Nlb4-�;�T�Ŗ�V��TGe�?m(�A+��3��#jX?�g<�Bc��m{6x4��9��)EŎ�T��"=E�\i�����dk�oځ�Y4j�cW��Ʃ{g��	<"~~�������t-�;�;O�TY]-�3����d�^�� v�"���/ݡH:����R!�t��Dc�^���CsK���E�C�l*���w��{�P -�48�בm�Q�U�r��T`1�^�P6&s�}a�!��#d��,�Z'�|"���ض~�2�fs��dS_0�f�4'�Q��u�&'���@]1 -����98\>�EߥnT�`�C �	���שy�E�n/���0�[�Pl��Ѩϩdx�.��0f-�r��n`���%��=�"��0%9j���1C��O`��N7<������P��F��g���������ꙺѷ�j�w���k<kd�K�A�j�ƅضKl�m����W�vV��ڟ]�iz�T��h����uP���������3\K�J�-�
-��
�X$�a*�ٛ>8��!��B���ˊ$�������m����F�w����ﾯ����yg?B�Py��ֵi���ŀ�8�[������_�k�����Ǉ��n����Y�yn���n\]Q3�46O��x�����C��'�����C��ivrR��6"��e��w\�; (C5�C�2��hs�=�0�UO;�tt99�Npόt3Ԁ�����mu	nn��H��3�״��>x�\z���6VF�Y���~9T�a�M��mP����#���[.�3���Eפ�/R��)����mL<�{ä�6h�"Z�j�wuV�h��WYRgaN��D���k�%��y��z���Җ�P�ޔ�9���y���p�����Z�]y����@^ܸ.ce��b���:�L�2~F=W1�k�]
GLsvv5����o�����]�7>0s�0ӓ�o�UyF��fB�C��ÎA�1f�,��g�����SŊ��2gs�:�Q�<T���U��Y�7�NK�c����/�T�f�6���V�K�\�HA�ɐ̀_E��s�/ݮq)�Į�l�Μ�zs���0�����_�������~�W�x�x���A�c�w^��n�M?X��J9躺�zC���&�Q-uiڶ���1��vf�h���m��選i㣁�4���*��Wn���ӌ�:2��o@�ʬ����Ω�i��ԯ�́�a#v,o]����}I,�wRc��M�%.ڋ@E�q\��as��BԗAM�H�,�V���b��Ή�3��jݰF��P`��]�
�m9ʛ��WV�CZ|��'���՗@^�gY��ɞ	��4�D��f� v�z�F��\�G�����s�4KV|{'XoV2e	�+�!A�+o_�%�u����M�=�r�:y2l��� <���|��ٿ,�2u��1؆��r����4�=Su-x5w��t�.IbD��U��l�%�u?j���5_ +rz�]"�\捼���ؖ/`����HP^���I�f����n9�b_n��η��ƹ�Z7P0f!�٭u20/&�O�V�X��_N��WD +�DT���Gj�J��dbyoer�Nԫ��͂ͅ恣+���(s�v��k�X�=L���]��45yTnS��+�'({ F�ˠ�ç�W�CU�B����}�&�F�L�R��+XW�W�t{���\b왴,n�Xu9Ԭ�GM���uݐ�.<�Z�Q�����C(�b�*��H����H.[��a��y}XwKԆ,PT��1���v��*��ᣌ�]`�Ṭ�d;��̚�p�x"��D��Bg�+^ �oV�^X�2��=̐����&���o�=�"���p�p�Ć��Ʊoq�=�Ƚ�1�=��k���!θ��t�\��7���G�i��������6��~?�k��a�t"CF�1�3���w�+0����6~�a�(ĕp�o7T�Vm,�Նx��1�7���f��2�j漅s��f��(�J�`� �C$X�6�K���v��GJ��-l��C�nW��պ�:*�!D0�56�/&`���3�m6�%���ٳUt*��8@J�s#��%�{\)2ꩾX�j����2�C �g�	�[�]��<#�gc����ٰ�n��V�qh��ҽv���1ޛr��LY-:Ӥ����B��޼�ɍym�Gz��]��f��Ren���{��$��Rެ]��_K3Q��\/x.p�t\�Ѽ�������J�*#K
P�� '��eg3�_Ѝ�ǽ�f�h��c	(�Vj�t���&�E촯b��+]5jI3�n�(�ެl��
EC��#d.�7.��;�;Ym�����	ںތ�wtv�8$ۺ-���F����Үt�	�e���	��2N�l<t��dv��~g�RU뒚y�b�W��>�:����v�Y���AG����@ܥ;6�Y��,d艨�T��� P:������o[%bf���Ttk�'�.�������Z��=E]o��QW��=6#']D�u�����SQ�֓������ծ��(��t�ZJ-����Z�ƭ`�B�q���MGy��:��F��
:u�g����A��ڡ�j����X�F����:u1Qy��c֭���U�Z&#c�V΃ͪ�)-��o#Mqh��Z��͓��K[{:����N� �v:���T���yy�O]���ͮ�lh��E��i�
�����lywh���`�8%�#�UZ��m������UL�Zi��gTS�s�d�ERRED^�*�̘�����΢����SZ�EM���"��0LG6��s�tF�D5E!U��N��c5Q���;�j�`�Z:4Tm��Z(��6�j��
;� P�|=��x�;�v�ϏB{�V��Y{?���G���Ƅg�h���ڳ)]���]�	���8���|U�5�����_Tݱ�{� ���f�����.4�D#�߄=5�>�����`�^7�~�4�p3	�{QR��{#�N��QXZ�-�2K�d��WYR���T~?T������S���E[q�8Jo��ʩ��F�lB=�ع�]��8����
�Nf��١�hx�8tG�#��j�c�oSUv�N[�я�,Y����K_Qk�J84�Y�k��z~Lheq���U#ߗ�TS#ٶ�*�F)�/�zZ��Śo:hb��z��t��֠Lc9z.��������)�C����{��7�gL���]xώ��Q�dʼh�53��ǉ�k~+�þmx3�H�q߁�j�җq;�9Ʊ](Mfns�B���=K�,#�P��&2���k�v�Ý����j9L�'�
_B.�G��P~�ι��,�gk�=
�i~��?ːp|��I�/��y��Ȍ݂]�˹�`q�j}0ܡ�]L��ۺ�ͩ8�0V��ٞ�8T���ao�O�g�b�;�;��M��@�0����M�r씯͸Yro�5�q�'7���Z��4T���,c˪HmrE����`y+�ϩ���&=�_~�q\����G��Ȩ�B�����9KM���4�]W02�W\O~�X'pz[��-6���AI��Yʳh��_I���������Fj�,7�ݸ	]�S��-ė�{���n��^�����y��̃F6]F��v��ʾ����~��{���<< � �8y'��Z�ߊBKEz�Kp�eP�fqX��j���&�x�`��i��U���7�d���Oܞ�kNt��B̼��ZGGM�ܥ����-��6=���wMK.��m�i�vF�X�-����W��m�\8';���!��vǁΘ�»�S.�
�d\�l�YX��U��q�����v��6gQ~u�t;j�"��-2׏�"�a��)Rc��yN�P*�[��mB�F��x��8�N�<�s��B�w�κ�-Άϭ�7ax�es��4���Y���-M=������t�Mz�����tW��81st��Ǜ_-5�s:����f�p�3�h��bVpݚ��Zf�3�lg�����xm�-��h�:As����V���kwx�G%J:*�
�3��|�V�I��bJ��Z����Q�أAi�!rFq`3q��0v#v�4Tj�.�vh85<=cA�ay�D���ppi�ys��}]>�ILh�Ƹ#��c������g�x�r�MN���c>�p�#�cF=�ޘ�O�L�������'�q��#г���9U/W�9����s8r�����؂_)S��g8	G�j��5���W�v�)�W�.�{ w,k���4��XO�Z��3WS[P�{:��H�8��'�='&�y�(>�=�k��y��+��7����`� ���}��5LlI��k���5��l���Ǩ���<��� x �����o�q�U?��:h|u��p��c��!�
���;�A��V����Cٓ�J]&��V�_��)2���[K�gD���=��^Ϙ��� ��ܶK�*+�r��ȶOW�F��	�C�;uT.�8�o���Ch�e0�ܞQc��O�C�KLI����L���ʥ<>� ��=P��ə[��Ppk���AS4'ouPI�l�� 7lT!�.�(�i�q�H��%R=���ڕnշ7sIQx>ɜx�ښ�b}H�otpe*��`o�o�Q ̍ٔ����%�t�%.�����U#�"XU�0�b^|.ff�D�8�)3wd��d�pQ5�1�['�hZ9�]�֜�	�H?yī�� ;pel"}i���̓ݑ��tV�X��[_l�=d�F��ۅ`Jm�]��b,cz���d���=���_)��q:���r͖�E��wk���X�#��U��a�ƣ\�m�T�4����C?8G&�@S#]L���IT�-#nz�ڔ3�Eu�:���Q_w�y���������\���b�ט7�����?^c�=;w�.�$������CӀub���J��:�6��hf�5�_�d�_��#r�9c��M�F�����T/�]��`�l3%�����;2j�0��o	�Ȼع�����k��{��|�{� 0�- 	J�R���ϟ__/=���_]�a#���:�����7uB����F�[7�vX6=09ߡ���sY�lڥw��i~�Ba�9З��lT��ؤSP�2a��nSB{ �%���m��%�Hmy΋`�;��J�$��M�$�&�&�h�����΋Ч�y�N�|U&�9�9��]���5rZ���R�� ?{h� @+�>�x4jq��w�F�?H\n�ڶ��x)peF�P~�0��ao�LW�<	q�<�<XH�eo$c�RZ��9��%`�ѮȲz��p�d+�(��r��4A�.)���9hw�1�le�Y�c�QJOk[�z�S���rn[`5���2@Ce�#Ϻ�����&��
a-ʗ�&C��ɵ�]�
�0I�vԝv�=5܄/MN0���:��}�V��,��s�g�Qa�+�f�֡Wr�zqE�n)7z��a	�}yg*����aa�$�W¢�H���=e��U�D��n5� �2�p:�NOm��$�QD����C��}T9CI5��PvN S	Z�k�΄C����U�Ŧcz���E��p�_�Mi���pE�띶����2o)!3�1َ^.���vǧ��G��9"^P�{y�t�>a5��q:��CC%͇��`4/s�)#��b˹�0�E�/!�/��륢Έ�W^7��{�������܄4�۸����z�q�=hx�{���<�� <���$���fGn[.��ιiς�\�sY.t�w�l:���� ��� (���^�?E��좲Z�me��sW52*{;��d��V닶[�CU����l�b�]A� X�)�ԭ=��=��B�9�k]:�5-�'�Mc�������b���e�[Q�B��#��PԶE붮lZ&Vgؚ#Q�@K��P͠CH`3@��J_��t|y�R^���窇��[�._@�N6Ol��ѕ�X�)���#Gq�<�t͙O�^��4�W��LS�QR����n�jiˬ!��v�^��PZ��+U&��D�z��Ǽ���.���Zzq^�j��"��.#fF�T8�{���r�fC45���]�k������&`�2����b�VI�z��fd-O����b2�C�@$��ը�q�D���dV�"5tlheq��{ʄ�~^�E�A��:۸�������9.��
\P��������3�,���$6���d9��?N=�C�b%mfl��M*`��]W4�ƻl�5c6�0&1��3����:Y�x��t�ϼ�Ő<c;t�4g�U^��u$b�<T�P_,Uu�D*�v��T�u��]M�V'q��(�wjA�B1)'����-���M��̤��P��2���vQ���x~�T�����@Q(��q�"k�v+��-��� �� �f {���7� oxI�D����+(DL"�#�H��������&C�WP�[��Lf�T�b���C�'��\�5�@�T堿�c�Z�x������6���\N�t�s�0���T6u���e�	���Dn� ?/��TMm|:YS_�6��b��~�c5�!��F?�6k�Ke��]�ͺ��5à�pm���7C~�H)����G<S9`�|���T��&��Pj{������x�GTւ*����	�ڐ[i+�X��ZEPŕ��v�0R������2�����s�O_m\�:�n��{A@�7�&��S�k�ꀏU��v��X�O�]�U,�.c�l�F۲C�]2jqgh��|S12*o9�"���htĖ;�S.�US"�'��++�ujg�{�ʛB|*�9�і~{�K��,?W�@��ڠ��_��Ф_�s�0�UIn���_,�ޭ&�D���U{�(��Z�G����'�8)�\������!�(�ޅŋ���bh�(2��#4�_6�|[��Eq���}�J�	����i��/�9p�	�0�Qq��7׷$⦨����f��R�l��:̮8�H��(uv��˞��b�������^{;0�����ُ}}�y��n���4}c�=�T(){��ĝ��xJ�[�w$�зǸ�>���mJ�[zM^�	�*�p=֣�&�}�ڝIn63Ru�7Y_3{���ʩ�>	�I�G��}���Y��G��Q�T(���V�� �{�f�f x=��;�[L͖┷�)Wg�JuN��m��m�L��t������A~�8jݱ}AM��o�[9uL�Bm������Q@�5c�xo�5A>�`3`�ciR�q��S��Ѽ�b�K�3�0��f�6F�[X�S��Ih�������2]��3��H�Z9'&��m* c �`=��Z�|e��1�;-�iVg;��@�Y��o�3WTT3\fwL�ͽ�q(w�e� �ɈӤ�������_;L2{�>�,�.�04��l'42�k���ZCwV�L5��XXY��,�li��O�X/[G:�h��~~,����C=��N߀�*�H�1<-\d��N��!�yJ��m�Q�Mo���� M�ƙ�T��k0N%��Z\G�?"��k:=���dNmhU�؅RզQ�ח3w;���r��'ڠ��Ce�%m2N)����cP�x�ng6�u⭆�CAs\SD�����A�Y�׷�0E���d�$]3b�!��ӻ�M+'v-�
�J0c� 0~��E|tmu�?�����bxXj��%��1+��������1�
Ư�����O�v9���C�ז>,�;�d��ʹM����O��T&�62L}a�jE[��%`�2������b���vm��C�4�|{�H<��'Gyw��U��uͳwg�(<3^[��p��~O� ���h)i�P(P������R���g�da.!���p(Ux*��v	I�����v��{�#�wh�."��C�Gg?h����H��b���l֫�j���-󤬿�d���]�ӈn�8yPs�Q0���OG��].�	ԩ�7�OH�b�M�*��7������u!�9M�0	�d���*u^�y}ڳ�_�M3w�vB���b�(�/��P<��m�WP����GQu�p���R}���m|�}�3��ΓW���P��{�����mjЗe��2�Fɿ�S���d�gYW�e����>ޘgӭQjZ�o?9��A���Я�{7��*�D��|��v�����7e[L��Z�I�=�B:��\dk�0#N�oKV�r��>��o2��2$Й�����!�>��ܦ��;[?�����r�<�*��Y�׳���jl�TJT"����z�i3ڎ�v�ʭqk�*�t��
g=@�s�ǀa� *�i Z~Re�k�~o?����_�:�������'��y��^s���[�4��I������Ϩy�a���}[��[gE���z'�$RSp_P=�VU���Qw�ۤS	aswA�,�Z�H �[<���J�5j@֘��Sf)��;�z����Фx���k�B���T��f�<����μ���X�|�2�DP�Ϳ���M����0a�3{������1�Y]���!�y�X,�k\�{���ru߬�.�L�c�P�!ѿi�s�hVn�E�֜��Υ��#)���q	�=��:~�t�����<�Ldf䮜�Fn@�Y=��p�h'��6�ܯTy���N�,(�VCK�8��]����^�c�z'L2�E���nV�Z"SP��JfΖ�3��_S��߭���`0��J�tf�M]sS��S����ε��^mO<r�+���S��J˂�e�.�1�@����8�I�|�*���Wu�p�\ҔĖƽ0Y�-�O�Vн�e�eAunB�fC��E��n
�*�xy����uT)�p�[�@��^r��STX�R�N��%xm
���+�g��G|���vo�Mլ���+�c�Z�2_^�7_Ӽ�ԋ���.�ڢm�s�(�D��-NX�,��j��	��6����:k<.���؇(n�	t��>{�LPz�)�����_���T��*����Q܁*��>Yd��Hk�Txz�O��#��ڧ-�(*��?�<��o���.�cb`?VO��{Q�u6�wZLv'on`b��<�d��ݮ9�v&�	� ��-f�d�{MN��]����4�s�P��u�R�ZO���h�d�{:���'YȜ���8V5�j.������bcb��'��YYin�J�g��@%PЉ@�
�"R�y������{�{�`<ܣ:�����X�˶]lz45�$��8:���@Ƅ�s��L�Nl��X�"Nݠ�^"�Η}8)Х��0�oO'�Q��/�O�Zj��x��������'&2��X]���Le�!�g-�O��7%;I��⡝��E��z�UL��^/��Xoivv8bK.K���/pԖ�c�t�xK�b�m�H�ӛJ�3����!t{ρ�<��j�0
�;�g~�'WY\a,��\��(��gt���GM�����j聄?[Y��`[4]��Y�+*��nf�GpLz���xJ+��>��>���1�嵬�1���qw�Zn+�)��tL�����j
�RP���A����\�����^"�5�|Ê�O1a���=����I~`��sߕkX|\o�7s��jhh�QD�s��Ȯ�Fx��:�����Ο�r7"z�³����Ȗ������Bh^�C��:R�i�X�CL��˹�2M�&�=B�y�fc�]�L[���F�唃S�v݋��!-�����k]4c���r���Q�F
��?����z<�>�_�����/7���>�w�wy�� ��W�skI⍮���e�Uc�AZ����e �qt���5b��gsϰ��s��лH-FBAϜ�GKt�I�u/.�/[o�j�����P��6v�ɧi��\� t#�#��-�p��ۄ��hDj^�x�Na�+M��b-=��q��ݵ�ح���v�:usC��"��޼f��jtށ{o��Z��78a����r��,���At\:�YV�΂:+W=ePghN�zig�;xp���ѥ]W���ʵmɡ��P���5��7�<i^^�0]��Qw1m.�Z��(`���3�Y�8]vҀ�g�q��X2p-��O���C�x�u�ӷ!��a<CT5Ó��}Oi�4!w)�6*K4G�'v��K�i��]�3�_���ë"��W����'��7)���U_AXA���Ԭs��2����j*�*�����H5�T,j�.;�["����0\��I��!�k��ao嘲��\�u�d$M�@��n���#z��vڥ�]X\^���v2�7OWS�Վ��7[��T�dP��L�*q����e�-�#/r'n-��R��?�`�j}u��)cJh�.{jb*�TkX*��*�d��"�vD� ��=�L�S�wQ�«6~�)�s��S�a�2����uh(N�8����[K-���5�Y�;1Gf���#�|t҈Vʶz�e��i�J솰ݸ�����y��}o
me$�y)��*�|�y��;�<�W*����Ѣm$�2d�f�
/҆HŴ�^������*�u���Ю��𣔎�*b�k<��c���b��*2F�M�y(X�#��3��2��0�����0��q��5C�.(�=�V�t�s��.�`�&=�1���o���h��l��]��w+���)q̷[���w,��̋U�T�L��2nZ%1�;�mN������{[6�Jl�Y��XB���y�}�YX, ޜ���������l�[SMу� �Lz�	t��eD�u�ڶ�����h��[�.�A����yr�3��2.���/%d �ǂ��R%yM5��ɵ�!,��� ��l��9}�z�mN�[�����B����[PV��aEw���ͻ���J=z��W�&\Z��z�C,V�.�S੪�VbP�|�kQ��3S#7��!+5�c9u�mGd=��/���A������A�|�z�2��g5K�JU��x\w��V�`��IPÜ��9K���4���1"���^w�2������M�լ����7{><3U�n�V��t����U��ZkomF,mt|][��B�I׫2WhӏQJ �S\�nb�j�����&��u���sX�y�8$$c�U�iC��u脫v��9:l-��s���U}J�<1�W2fg��{�����0j^c�	o��6�R�5�X���}Ux�����:��OC9���/�wn��~�km��Z���:)��o��榊�`)ִ�������b��:;�(�UƢ��յ��:q3�Z����w��c������������{wd�-m�툩��U�qOZ���th��PY6�����3ASkS1N��Ӫ��X�Y*f�zq���6p|�{8��m�c�q��c[�"NΊ����QL�n�����$��m:*ּƚ�F��VZ��X�Tb�fu��(�Ŭm�Ѣ����yh��MSm��F����DLkEi�E[ͣ���"�6��f��ƻm��1ͫU�S�S|��N�)���EPEL[h�mu��[�|���E3��5����/��cm�(���`�v����2DA���m�)�#X�lDi�G������k����֝�M4[n��F5�Q[)����ccn��$Q]�s��*tUAm�"�!�$D���&��W����|Ψ�;6U��ݻ�V,�N^�6a���C�c��������J�)A����P����;[���>���պ��P���� �f�o0����}y���b��a�#sZ�@��Q��*�C���6����'t���UL��QM���+pL�,mW17n�`e�Ow�V�)��PE��; ���A ��X{�T��w��	�V:��5�*N �j��Um� ��7Xu�I�E�}�S���c�&*:�b���2q^Y�<\'�<������2yBâ�	ۜ��i�t;�8&5�5����Tս��xTX�8��wg�Q��wM�l����4Ns��� �gP�܁�1�n{|;�>/���$���#e�B�|���Rv}��jǷO��T�X�|KA���n��[�ng]70LeCGQ���(UHg��b3f�{5F���8=ҏ˦pmNuHcc[��E�����آ!{0���L��=�>ys�	����ld6	�شn����i����Y���!�mm��}��Lit���'E��G���	�49�0(HQ��{�́ڨp��M��%��N�۫X�gf��6	;ޓ,ڶ[+��ʂ�Qo5�i���^~��pZ�?��JomK����u6Z�)�/��ݫz���(~�����laOUˇ\�pb+\��,����ǖ�5�
�t+����H�S���,J��K)�����	u��5�2��#��uv��ܟ]t�>�W�|:f3��l��n�2��Z�7��`<<����oxx3xxx3x{՗{��1�l���Xv�Nf��c ���$X*)8|�O\�ZbL�*�3�h@D��E�5��2ϔ��r�t&�2�2}�/#7j������˥0���!�P�0���>�$⸺���|�9�M#�+zJkIɗi�����Ez�(2�e�>�jހ��$��Ҥ��߲�_�������\���6�n�n��"�2E5����yP;�Ǡ/�M4�u�(�����K�k	���ص����U|�l�¨�U��$9Jh���k�$��+�e�	����k޴��ӶW�yG��4�Ԣ���+{sVHSl�y���ɼ�`i؃xrQ���Ndvm)�q��*��Y�+��Qi��"���c�'!ο���1����T�������]-NJk�D��G�yIks7�t�%�5�(|�����r-�uT��jw��Z��>��-*�30�\t�z��qY
0O�����~}}l�$v��nd���оMKF���RK�#L2>���U�)��X�')��H��|d�՛�О�FN:a�|��֌z0��k��JR�΍l����S��A�G����{�\x1��)9Hb�AT;͙pRrScC用���Z��9j�Ѥ3	)��<zs�����b;��ދ��K���;+�����R�|�������}-^�K2!`��]COh��C_g�7���y����4 �P����Ͽ�z{�~_�Ӿ���}�%�>u��wfS�c��P���З���q|�#���%Za�8rD�8��-a=�Mo�L�����c��e�:'��,k�I�-�>� �<'�[o�l�=]H\;�b焄�t/�*ja�3�e�ru6���9,�g�{`x�4 0�$i�Ķ�F�L�
�ګ-�<<��rO���xu��n��y�Ѓ4P��yP��PLSI���)>�s��0�km����͇ڙ�g��.��n\�leC�} w�}�}�އ�b�H*�5z�����C��OB�p%H,�w���`h�DÍ���ۍv�C/��w�@a����n٘1�4"�ME�0c�g]m�8肙lQ7<���0��j���f�i��ٞs ;����.�,]���`�DtK�!]�#E��ڤKZ�w�	�M��N���?B=�Tuw��;�TV�=^^�6".��*��o=��ֺܷ0�*����W-9�,4Yp\�ː�|^�z��8�.���� r����n]n�=�Ʀۘ�4 ��9M}�Ք�n��S�n�[)��o�&�_WE��_����< Q}�
n�w�}��i��̩&�2����kY��2�syLF;��n���n��ӑzV7c�p> @�͇�I��z��ū�r�m�G�Qpe�3m�:e��t�Ptî�WF�o�diŴ(q�v���r�5}|>�[���?9�ZA�H�"�<�{8^��j���W�IXCQ�'v5�oL�-a��/�T��X�~�#hr�2�RuoH����4ww	��#I�ǩ~	��|d3N�]�B.��y�R\�iqԆ�A�k�8:���swߣ̒'�Ǣ��,/��?r�ܠ�<���<�4�Q5)�v��i71��R�}k|Z.�d򅅥�8��$a�$�����Y��cL6�0Ӓ{7����-��\D�=Y�Y��"��0�
2Y,��q��+M娦��~%i�\`�	�\�-T�tNk.ᔽM�*�Jr</�l�gԟtد$�-5A�<C�+�'V�'�ɿzo������[<b^!�_P����'U�L���	���3"�if�t�3��2C*{"W-�9;��qF������s��Z�BEW�.
�~SOw�3ˁҫͯs=�})kٷ���rY+��0�a1]��@bI���}�:�h�7;��r��Zk.9�Ma1paŉ���L�&�3bNTzu�<O����!E�ih��F��Fv�� ���Wdt�A���^eV�l,�I���˚+n��o�1���OzѢ2��;t�Ǆ��,k�l�v2�զ�+����'*���
� c�m3iXnp8��Aa���N̑ʹը��nZ��注+���P�[tY�q�F�WvE]<V^�8;3y�| ��B�4-P,�E PhZsn�$6/Ы����86� X�T����:z��U-���$C�P(zj,�E鋋&���8�^r�Vpw�M�{�d@Zt')`��44T��M��<�����v3� 6Hg)��ʤ��瓵vG)����mԸ-SS4ƀ;�M�~�Jh�űr�iÛ�2֮]�6�&�܉Wjvi���i�ۤ�K�TŶ���AH�Jsf�Z��Wr�O��3L��V7���}����g��oJB4����/hF�(��5�=C���5������}�=ꡣfȎ{M�q�z6TV9��V��,;�<b��2q~V��9_��P�~#HyΥj�_IT��9I��ݚӯl�_X ����&i����uc��m��-b`;Ї�`~c�h��:\*=������Sy��M\ˠ뒮./ΩQO���c��k��d��a��lt�]�d�C���SV=vVӮ��t�'�"B�oM�z����W'�K�O��t[sW���m����L�������9Qk�ġ/�DD&�u2�#qQ>|le*���k���v0A��1�ma�M3�\U�_�T�|Ľ�!�>ݿk�F ���,R�~��e�����1���h#<���y� ���q��@�L3.c�3Dy+Io]f���4q
�șGMX��2oo
1:=�˫��g�u��Q��ٙ0�6�Ys+8T�u�ML0�̢�w���H�#M!4
IW���W37����<{�C�}�/<�^[ZF��[grT[��е^�zXy�|�|e�{�A��̑N�&X�t��0���v�7����\\7�=fQ�ؽ�"}�����0�f�lk�g1��$�U��g���LO���P	�-z�	�b�,�/���`���R�O�T��f������C[�]�]Cz��%���D�5�s�'/�??d�'��7�f�vD-�g��]yGe峉ՐF��@-x�|T�p����tS�4�Y�9=���S\sme��Fk:�z�/L���*�4��WW���w3s5I>�	�N��G�+2�z��%��5���`#�B���f�*;�e �'^\��{uϓQ����D���x���mz+���Ԡd�z8������{ܡ����m�+��G��Ծ���1�7?F=�c�*ְ3�L�z#A�Dګ뫚��=�@���qbR��\Pa���
��k�x�"�J�nxO��@��зb�G=_K@�=���s��I�(נ%9�T�`�^z�r"�ӏ>y�$І��XoT�U����ƨ�U=����).,���{,&4�1\\�b/�����2I�F籛YcG
_I:�U�-��u��j�q�4��<Y���{�����U}�U��	���-��@��^���ԫBr�;����:S"#����,ɶ2�V�VM�9}_U�0��7� x ������7}�Ӭ'��.,DU���ZrpV����si�4y��3�^��O:�&��"�[�1��٩;ƈ�p콗G�yO
�0Qj"��犠y�+�ܮE�YJb9R������I�5r�w�<6`���C�K�2��[�\KwT.*�󶮈Qѣ
���L�ڮ�2����ܦ��Iv��8���h���q��z��
�@g�Cw��ϫjtn"�F�dgc�d�4U}�;��/��Į��I��-y�?�yP�r��˟z
�D�c�}��N��Y��o*�JJ<f�G�O��tM���͐�_��ő���~�Os�v\�-��d��W�5*m��ik��Z���A��=Y�<yW��"~� O��7�&�R�mUK�uf�Yx9
�m�`����?uK~�&jz���˧�g���hK���y��<�]�.������è�C�!3��f��̀2OY��tQ9���m��r��!��Ӌ��~��2�����bj��}�OM!5g�|��&�y�ú
gj6��d\�mF�<�7	�R���S��j����2�H�6\�ޱ��23W���շ �Pڽ��U%�>��Zp�����n�Yt�3z;��(�r.0[�m\�ukS� �$��:Lh+�k��9�'	Z��pF�f;��㩓
5��iN�a���F�l����ͷ�i�?��}�-�������"Z��y�nٴ��d�`��b� �^E��῭YZQ�U����P9.�E��Ih���'��f*)�m�;XK���\��oآ�0�(��.l�>���Y޺���VJī����%��9Nm k4�T�{�C({O%�BYB��*�i�๏l�Xػ`z��tV!Ul]�L��]�j:g�I7��O-y0FΗ�b{]��c�:�I2Z�eNaj[pCM3��:���������$���l\?hp��4V��-}2h���E�
�"o�^=z�e��j�:TT˝�zv&��\�4{�2���j�ǆ!�\�|d3;��K٘Eէ�c��_���%���uZM/BkW�m�3m�N��%��3�K�lo',�0�s�,gzi~S��L�i� Nw6�C�l�T��:8�}=�P}iA��@���O��#�����q���m��mN�5c*ح0�b*L8�ڭa~�d�X6�f�P�V�E`Ha#姬F�q�>�R�po�(˫������uK�*���(NZ�9Oޣ�2�2XN!r���0���l�=�D����m�fC�8i���^�Vs�EDmב���fF)�XVu�}\3$ح����e^7�� ��mZ��I}1P�F�����8N��i�
�(w�u��	��^�j��>������B�zq���v�n(��]��$_|���ۏV8���|xy����{���0�m�-dY��0fh|/𙅇*^F��p���b��J9���5*fF
�_���ŵ�������5X���ܮ�L�H�v)�}X`���t�ʝ������������9q�� �� �5��h��o��h!K5�0��^�'Kש�>��a팃���t@M�'^��wp[0�����E5�=e�Y�O������3�p�����_A��t�Ş-�l#�U�}�
mm^oLU]9�ZN'Z��C[w(��۞�F6�R�,!b�d���`҆@�����M�F�C^dȁ>�}�Y'L2}����ئ�c]RCCl9���\����J�~ػ�j�Yt����E�`����u����8�MjAmJ�M��h�˹�	���b�{&��C�/"�u3���*FD���L�Ʊܥ���4˭E\v%� DQ:��:���v���be�%�'t�7f<L�j&i�70����r�[v!�����5G�榀��݃h�W?#�"��0��2`P�h���l>uA<�Zs�y��l1�i{�����l|86Z���Y�&bӓ��86���¾Єs7��a��-�%6�ӘaE�~^��s�ҿ�����m����JW�^��ɺ.�Y@����j����c2mN���%qu�	i���V�y)���*�{�p־��w���f���Ek�Cۋ[��酮�Į�m�Rq��-�:�ӾB��*�h��Ӄ��"���;��''e	l8bC��IqNiW'�I��k��d�a�M	��:�; ��"�N���	{�j��6�s�
 ��+�V7b��W$e�R�E�{2xm�,��h�q�N�K�(��bSnl���6��4�'�S;����k��֡y�V��Yl����jǷO���tN�;C�k��Êv������0�������}(l7cnhS6�Gmlp{������3*����������ÍW5#%�W�2FƖ-��*4���U��S���7�u�	nz��b#7V�ޞɠ�J��R<���g�>����r��3k�����C��}�_�V;X��w�ѣ�1`&���#�3�9��#��P�^���y�(��[G:�'�ř_uE�+e�]��3?MO��K��uٷ���{�[n�!�Y`�\D�~�N�L'��ؙ��ڎKf6�ɫkj��V7��."�6)�^�Sື��ʸ�ٛ�C�(���& ;`��Ky�������}^�O����z�~�����x���ђ�L-� GN�k��=lv�k���D'_7�~��oܹz2kcY���
�#��l����]t�t�-����/��&U��-�5��n����fSx���ʸ;q��x�l&�c���:�+w�*�cw�P��g�3���6�lhލu���yv��^��X:Ľ���|-��呟A4h���f�p2�Ф��M�8haf�oWIOxN2��ї�M��0.�O�q�1�&̊I�[6ēa�+6�&���+8��c+-��F|w!m��/h�_lwǲD%��䝦�gz�Yn���Ԗo5�A/�̻�Dt�do;��Z��TM@�mE�]o��x�]aInJ{S�'v_S0e��;h�Jz�@��k�H�ȹ+ە�2�J�b6ٗ�Z�WI�1.�1m*� �f�gb:��Q{u��n��������x[O���9v�3G��s(M��,E���:ʉ���NM�%�݅��qR��bi�.M�ڬ����0%�tJ�ܟt�b �Y�q�3��aw`�<9�x`��ڼ��g�Si�1ގ�z�}�:�B���۲�8)a�,Oٞ\���x
�yi���<0���ҰC�u+�{�km�"�6$gWwv�w�C�ԅ;��O���+�ְ��ޜ�U�tEv,9k5�d(�T.����|k�^�����+��;՝,�P8+/�
�w�T�Y���4�RbfZ9�Pz�H\L�'�M��Mj�Zcz�νN���
,PC>*��J�\�z�	Eوُr�4�s	՝�ݐkr~�7�d�鲈Z�kJ�3-x�$dp��f����-nS�x�1�YHp�eg \yZy:+�t0�Su:���r������f�J��IW'`�b�t%V�#a�;�R#}Me!yM�$HJ�s���LH�JN�^_��y�v�f��lQ��Ã��z����;_�&Ak�f�ݝ��cz0l�Ѧ
���DX�j���&s`t��,ݶ���d�/F�n��.��[b&�FP�/�3G7#/��r���	�� $��sO�I�3ۻ��hǠ&ks�n4��U�xvkk,�mFMJ��F���-LНR�M��Y�8&��a�X����?�7�jʑ�=�7|l㓆М��i���r6���x��Q�e+�m];=zy,Ӕ�y��M��-���s�RZf�mƔ�������m��(؆��a������.����Jd1k���@���hZJ�,�g��B����+!]��-=���q��Γ*����1���m
F�Y���}���_�E��#m��,}v��]n��ui챢j͒�?�_T6ka�_e��B��G#��2�m3n�R�8������Q���N�_*��fyj��Y��]��ʘ��κ��	Yd���V������RbPv4o�'vP?e~$/�.Gi�c���71NlF#�**�S�CQ�b���ST�7pj���]��Q5EQL�AmN+�4��TQ3V�ٜj�Ӛ��[co7\I�����n�gTEDQ��<�yۢ��>mĞO�U�g[V���5�-h��ym��ShŬk������M�TTm�v5QI�(�Fn��c�E��N���o-��4TQ�m&��u�����v��ڶH��[m�'v�6�kI�mj5��A��f* �� ��5�kTMh�%N�S�"*>gq��(<�{a��1�TN�TUQb���V��Q3T|ب���3����Gs�V����`�v�鎴EDƱ���mU:
�1EC�ųDIEU�Sv�MU�i��c��E[[j��v11�qǄb|�γS=��kcI��v�|Ɗ;���m���.��A13�1TU�.h�����O��_�_}ߏOO~S�D�u����a=X+�77��XݖS�h98�i^�J��v�+��5�kPo��`�0�0�0�a��3aDX�c��~�2�������
���o���(�[>��t�f�G �m�"��A��Ϊ����S�Y2}���qH���9I4��������"���ۥ���QwgQ��$��t��v>��Ző#Fߺ�O+�^Q������
��#*#�ݮ��FL�ˉ���҈�m�^������Fּ��jDXmJs�'�nb��fU,���d����cʶ퍚�均n�DL�m.C%���X�R��xR��Qe�j�]��kX�;[q�罨 ��YZ�UW^|�I�}�>ݙ�?3�i����pDejU��K.N�i���-�dZYC���GhF�L}������ �d����C�Wrg�x�����#^j��늤_ٜ�A-�*��3���>����D����MS���s����ݞ .�S�޺�j��AF���{��sỜ�W�5����i�\ю��L�O��q,�x�:��)~_>"��&_/��R�|�����b#e=�p�<.Z��\�&v�AFidx��D�����ö�@�:�s�x{��0��H�ǚ�T�� L�����q��-��.���	ɚ��[�c#z�h�&`�s�Y�����F�s�YI�t6���^�,ˋ�%l�n��<r�oEz+�}Z�\�+�De6��E���l�(�!�x#B�k�)QC/����/]�)��=V��[�f�KWWd��gFG����x�k%��y���)�^~bgS��41�Z����+yxxA��'�:�k���<�݋��g*��"��,�����.=�}ڬsP0slqg�w��y�נ�愹x&t���a�v�g�n��&���?�`U_����	����~�P�S7X/]�f����\�Zئ���[�ۻ�����n��C4�M?�&&��a��i8�.�`?���J����Ƕ�4(��nB��p����\[6�I��(�:���5��1p��A�-"�w �9ە�Z�;���-
&`Z�tT ����5�w{�xi5�hDz�P&�,���֚��.`mnj길=��l�	���/�P�j)>�	e
�S�춚ؑ�|Ã���i���S�6&�ڞ��xYrbM�Mp�:}�����Ƚ��I�H��R���v˰�X��Gpk���V"��Q�>;j�'�W�v<�5(��[6g�E{a�'��]֥���W��0��%X���6�-6�b��3g	i�Z�4r0[-p�����f�7�����]0�L�?D���h�Ǻ��F�qg�:��.�Cvd�\��e��V��e�N�R�g/��7��q�
�n��Oyӄ�re�]
���D�ы.�Y�eX
�p���p��
φt�Z���x��[�hᣊ�5
{ܨ��6#c��sNԯ�bt�n�6HXE0R"�? �>Mʿxڮ��(&��?�3��;�fK��ߝ��9Ai�<�t�Y�w3�Д����W�.3}(��{rZ��_��6[��}>�(?����|�&��D�=B0��y���*i��U�D�V2�4�����T,�0�Z�ae/*L��0�P�����k�|�#y�lSHOC����1�nYL�'Vo�W�iT*����L�oN��-Gs���������� ��Aw�y�i��[b�f�&�@�`��"��is/,�:K{{�P�zb�v'Z�~m����Ȫ�<���Ȇ\^�Q�/8�.R�-��v8+f�B>ͥ\+Ǟ���?
=.��@��Q��]���*/��T�Am��܁;�O���8&��p����l�(��*v��th|�f�r�lۦ�����)����j*q�������2�Т���M�"'	�U4��>��{�c��{�J� ��[vlrv.DD�^D�$��>Fhe��SP$d�C�mn��I�75��O)�Zf�#�MF�E��Ə�R0W���R)��gg��6K�ޗw�v��Q/�}c���Mo)�*C�.��>�(�ei�.T��̼�D��������O�u�{X�x�����;jY��"��DF�[�{{�F��;��{-�@$���β���d��	b��69���᷵ʮ�(jϧ^���1��WZ�m�}�U:R��L���!����*u�\&���bl-��"mZ�ʹ
��~խ"���x��U�=ޝ����I�tB���e Χb�r|[o�U�'c�eM1ѹ��V��Q���k=T�Z�wMT��`�O�����e�߄�oT�����n:�:���]f�E��7�o���j�8���י,���b��������P� �Ϭ�/1z�T��Ѻ��cf�U�)��)��?�Jhe-���hS���9c#��FA�	b�U�=�o�{w��)j.!��!�Ǎ"ጩ)Әヰ��ZJV��'�m9��}y�����F��~��ס;��%��k�Ȗ3��Pޛ�^�WW�Q�Duآ[p�24+K�R�Xê�.i��\�fڒx9��}o_�P�@wM�U2�;���W�K�f��?#�i<Ⱦ����җ���c|�a�ݻ�/���\X�Z��b���҄�����B�Tj=skS��
ȸ���\��A�`�1���{�"=�A�������@�CE饀���c�}a��n��<Ǫp<��:>�v�)�*б������<��%S�h�{�+�>�ȕ�/\/��Z�m跲�S|�^�jPM��2�4-)�V���Ȧ�sz^\��;��ހ�	!�hol)(z�Dx̽w�PM�r�^hc�LY��+�j#;��3�"5�^ڻ᛬KL�||)�u����s�7�+��L�� �GW�d���#[�c�[*�����bW��(f'����o���A�>c�J�������|��D���\ǊQ܍�*72�V<��Ƭ���!�焜��(#���>c�k��b@*m8z3u	���͑��:�1B[7���196.%��p�u�^�]5Ǵ;e�U@�gt ��Q��T �#����w�Z��S�y���1KjNNnhǗ��"㓁Bj=�Wl:���W���|�C?VM����/�j7�ݠ}�Sf�8�F�߄H�9�1�<�>{�"�1�R�=ߒsz���s�ϰ���	�\	[.��JZ��&�	eS�q�G�5'�ʆ ~�,9�Poԑ�yo�G���t�K;Pչ���(k�t{a�h�Ei�(�Z��r�]��%N�B�>��\�X/)>9/�8f��h����
A
o#�E��k�P��6����=ء������WMŹ3�4�]�0 ��HZ��z�6pg�B~y�G8G&��v��pD6jS;.OH��P���7�7�{�0�7~�.%�B_g{p�~X@�^![�28�W��\}Gz3[QZQ�M���%�0��A�������6c5�=9y��k�xN�pId1CiF�B�@�����u$��c�f^;��\ą�q�c�u@xMZltN�eY��N4�L�Y���CA��ٳ��"��-��F���ei�?@����Ze�0g��l�ג&�F�u�TY���y�I!qȭ�����Y��~�O����}�=���`t6�+a��}���ڑ<���|�n�j�幌�j+/o�o/&�/D�s�/���K����W�4���H�oAa|��!_�ϼ��/��	�u�X�SU|/zZ�}�dR9*A���j2Բ=O>\�����X�]�X:����9/�{k_��W����L<���1�o���&18�H�Ơ-l1��)��=�lO/D0b�e*����7��(�M��� ��a�w���虡{�.�,v���t�ͽ��S~l�1m7������o>����h��e �7P�-p�ܼ�o';Þ��;E[�K�K,�ҷ�����`�TX���e�Vs�����Ig�u>�Bj�|�P�e��ܟ�SXz.�[�D�"i��g�dɹ�=�dSe�D�mO���P�&O|�EX���2(~ߩ�����RIUK��pcA(A��ת-�ъw���vKÚ��8Z�"�z�1$t	7C^cU?]�{�n?��7���ט�׹�e�������W%��.geb��LB5L!���#F��2w�Oo��8���������;��͡@�;$��A�*Un;R�)�S0$����ʽt�-�r��W-�l�/-����.'�]���'��\m�x�g��
���b�N�Jױ�2��j(��YM歱�p4�e��6˜+��$� d�*�h)�6�:a��*���1u L�b��l�tĦƾ�L��؄�k$V�}�1��>��໬��֣�2i�!t�� ���3�b̬Z�b�L�,�!s��Ȕ�{�7p���r��Ed=!��%�AY;OUbԄ0+a���bg���ǁ��@L�)E�M�uYTb�V�V�������N���%�]S���k�i�td�؏:�e�A�n綄����/���{Cqʋht"ʯ�8*�5'!EJdS�-�:��Mx�ΐM��At4��sD"αF��1�r�k�\���Ò*�ɇr��g���p85'���%��̓{8N���d��9�!4;�Aܭ=����g|U(q����ը�q���@�._\��]G+�eQ�[�2n֝�a����lX`� ���*����:?N�����9]C-)踡j9����5���o*�]Seaμ�J��3�0ނ�0��c,0�}p>�k�d�eN�n~���W]	w�cO���-�4)r�9�1�7��Z�*�/lc��չj����X�&n�;�HH�-o�����9o��ڳ��Ô��<�ko@w9� ��g"Xc�I�mS��CY���%��<�<��㞻��Fq�O���L��z ���[,rwwj=����6:�gQ!��c[�uk>��-Az�G����'Q��=p����Y3c"�5���f��[�K�YS"�m�k@ǻ���2�������K��<�dD�*p�3�&�G^U)���v���A�>������e��Dn��t�;��gjknQA�.���a�fw�SԎ�4�cA��MEfY��Ԙ(z����-�q���=�sI���jhh�QD���$6t��	��:(r���3P���La�/n��mS#eb�)���zN�3BWB�҉ܮ��;�5�m=ܵ��+�s�$؆&�)E	���;r�x�mu%�Tw��'i����v#Qi=�n��z�u�5R̒�=F��g�n����r]���CE��bFch�}WfW�d�L��D!�� )���y�\�i��p�5nU<�a�:��r�-,��.G=�2j�UGf��X��*��٧-���c��42����z&�3qj���n-�Q�:'1�-�`ST5az1���Z^��aeN�nf��;�?6JR���R���oaĩfQ����C�^�W��]���w��;R�˺�U`0���#3r�.�X��b�}3�9:�d{�X��{d�i#�%I8Iу��Cc"o%K��x������n �[���f�]u��yigqq�����=�mL٦�鷓V�pg������Ό�
6-Toqv}��h��=�̞p���)�]�!C��YΊ�qAY�Kiki`V�x����Vø�˕\,[x�R�Y��:��vO!�}뿲���_37���SG/�%o�H��s	��yW�/����"����㚧Ka�+���캫�U�ד�jTx���-��t�8a�dDh~2[a�.��_w9$pImKo�&�%F�g 3 �p��cO?[�1�����6(��nYܵggs;�A`^3�f��)z5��fm?���"�������,`ksp1]�q�(3E�1a����v�Gu�ym٘���O")Ⱥik����P��!�8z�B��z+�(��f�����6�D�)�pPl��������^��x����6���r��Ǉ�y?qb�*���D_yBa����Eó��}�ŤE`��+��
�t�Uʒߨ&���1F ��ʢ_�R�OV'�T_QbT�F[���io���zN/�޹G,}�L�3�m�9RV^�>c�P�E�������Wn�u:�%ߌ�]F69ú�N��;�=QF,f���@��f�v�$
����r����y���8�[�o�2�塮��!#7𒎻��0���gd� ���\��S7:�[�����7ՐM�=X�v��S��iҴY���)�R���b�s;�FW��������{ՂQ�����a�_?0B�p��.YT5[Ќ�Ȳa��#�����犃Z�Ei��PH�����m�6�³^�yEq�-�U����jS|m��̕!F_h�W�ǧ��0�y�� e��S�0�� ɷa���<ÝB.��3��ޑ["��kjTI�΃�ʝp/�.J�+ُ��x����C3�ri�f�ͨN���\��^��~�%9�S4w�����!��Werr����|���x\�.CsMFV�9��e03G�7n��W���s!�c�OD���9���n`s����ju�3�<4'$���c�ߘ��#�d���vD�"�-*�=�*b{,���y�3�7:�Iw�y�,<�O�?Y,bu�]�cA���[�waW��I�S�;�k�|�jY4��Fz�ŕ�pGW@�a��N���a�֕��CtӾj�r�\�0XcF=���pF1�N2�]C���L���L`g/j�n*�uF�yw�9w���ψ<|�a�˻Hu���9� ����V;=ц��e�^2��q��w�8���x��>�O�����7������z��g=��;$�<��sM������.�Q��;��bm9��CN/�c=jE�5[�W�2��}3^rn���ǵ0f�UY��)h��v��ș��xl ]N$���ٳ!0�5��~��=����}KR$m���z�s��Vݻ<2��e�+6�A޹�We:T[E< A&�D��W�^�)�X���s�B��W<��
�J����H�Z�^J�7;w������oAtwE��B�����P�"��G�T嗢J� =b��X��{ǌW�-��:�t���X<b�;k3v�.�jBc�Hi�au��PC�-2?�e3w7y�r@j�vN���i̠d&��*V���U�6ne��!��Ɯ6w9��V�Aϳ��c��lP8�'�p��'e�5ܭ���A��#t�,�,�vN�p��k*�ϐu/�q��TvS��G�ܬ�-	6��.�t��a�x�9��T�$���4���3`���Qw*��[��3��q�V�(�Av�kE�����iZ _#���]kr�+�r�ʽ������N��x�����k�O5櫥	kr�7etST.�E�.�Frb�HF+Z��X��B��ƈN�^���X����3�
\�<9��]:�wO�S��=x�cvJ�WX������l
g�_C��/sw�[�*����+�]�-W1n�N�z��ӻH�K��dGi���\�_w;�N�El��YR� u��NX��>�������eV!�fh���w�wv�Իuˤ]5��ȑ�!8����L�t��df�l������g&~�����x�.��9��^��D�k����Eղ*JK1' �V�S�F�9�޸5�5�EZ�O%g�B��Z�x��s��#*�k�;���l����+�*kޥj��N��c,r�8mb�nS�u{&sEG������Tg�)�O�U��J�'`�]H֯�n����2�ӼzЭ��y#��v�j
������jf��SE��xMF�a�Yuυ�q�\��S]Y���vws�֔Н�DL��.�s�f֓��d7���sr�}B�D^9f����<H��ԪaF�*�g�:a)G�AVb��A13�Bf���l�I��X���cz���&��他#�q�)�36�Ia�م��1�x+�H~��GgoHoTW��GB�7ڣ�{�ZU�
�����JQaѮf�5[�*���f<�4�a���2���*iO}�X(�J�P�E����90wV��[a��[In�x�R4��7�3Q�r���V�J��.�qv����Q��d3���ݭ8hZ�+�5��q�o1�&hF��yPE��s�̖2�,�	Z�qv)o2(s�P�.�{�웧�����4����a��d�'q��2Ȇ�_\��k�'�0m�&�g9�ۑZsgbJ��K���=����˔>��,�Vt2�[l6,�m�c�SwC#�qiH�Vݸ��|�R#q9O~��<Z��pk�}�n���m �2 l�$d�F�(�ʍ�x�#�j�إ�^A壪�fj����1�^w<T�kMj��:���l^mM�4m�#a��SQi�Iq6<�;b���c=i|�j�:ǘ�U�wm�(���D�PDכTM�D�5TΜQڴAQ6�I���D|���-�X�G|���/#F�&�DL��7Y��]�h�t�Z�WY�"��RVԆm���Z*���툍���63N�N�͆��&���t�UPUZ��AG��ã�j�a��$֪&�ٴ����k����yk��V×�U1��8��CN"�,CS�(�mU�X���(�d�b��ֵ�b6~\ݵQl��t���TQU1E�5D4�͢ ��(h�:�ULMh��QMtP�:�1�5��Ng��Ay�(4E��m;kQ��Uhz�
.�iщ�tQ7�|%�c>�w���(���_v�-�Y%���Pt�QW*7��9ru�wK$R*Gd�3N��VM_� ��_�������_�ΑӢ��i�l{(X`�v����|�]��7�a����iE�`�����mwX,�I^� O������쿕yD��	��,���q���?���u�$6EA'����"���P��> Z{���,ڙ��RA��D�>��c]S�<&�K�t,7Y3C�FA�q��W'ٔ�wO���?��U�;�E׵F�o�IqM��ώ���u�l����s��ߐ�yp2�6�AʛaCT,{�A�?Y����$N��X�B[p`�sH��V�a��Vۭ��V�����v����3���5���9t��;� �=��I��-�{YE���4�R�|=�-��kK2Hhj�#vX=9���X/�y��l��X8^Dt�S̷u���#|� MQ���4�e�����?�S5��/A��߈���B���VH!�ð�f1��Mf���Q�혭�I��J�w\U2/#p��O��O�vX۞���.9j�xQ��� ���-�}m�u��O��ӱ�Tћ
e��CȮ�e��0������n�m��k�����ǝ���eRH�V�fl\አ�7n���	9i�۔��^���h���(���X�o���h��+�o�`wb4;���3h�gC�*i�fc��w�S��v�,F�Y��h3�`�1�^�%�A����;DW��<�	l��9��ܧ�A
`���Ն;u�-�74
Q���][m+OzW��������Lg~v�qm����<�p���_0��)���]�c�: �8A��v��y5��P�Sw0e̀k��RG9h���_ݷ���R�`b�t�j;�e�����F&*��wR�kh:|u�����!�(f�}���
�e#S�oW��T�l�s۫n���/�0�S!Z�5
���T����
�P� ��LL.�
��vX4>y�)� Үc��ج؅�E�f���<)���ĕ���p�L�	��P�	�(���|ϠsC�)�ϖ�)���7�;h��Mq�{&n/�oS���Z�������v�#��e	=P	T:#��]�����C�BN ����7u�!MQ7�3aY�wpD3f>�tװ̐�`�E0kͳ���}tq����;�ZVC�Scs�����K�b/y���n,|j��->�X�בR�u��7�m�<�gK5�T>�jA���L8�f��x���ؽ�R5��O��ؘ�/���V�&ӗL�q�Km��j�.�ߩ��S���(w0*��W� lއ�6�å���Hȟ��U�<�wƄY�<��oN[g^fy�4y�q �\�IXu�OW���̼x�Ԯ��0��3⮱F���)�Z����Ƣ�	Lf��WPs��خŽ֏W����������k6:ƪl:q�+��O���K`F1E����>������x������~�{����{�6�>[�o�"V�bn�3"�3��i���]�9�կ�����3+�j����YiS,S��6�B�V0���!��9�kOM��/`^kݼb��ś�RS8�85��u����H��1)�*��r*���;_���xV���'�o��,�����[ϻ�\�љ.�Ѓ�u�-ݺb��\w�Ү'��pj�ђ�BáH�Eۓj��E���|3*����̯�����?�F�-5*_���Pޑ|KЎ*y9
 ��s\�s���U<��~��x�!�c�Ҡ}��`��)/�����W�g��s�r�c v_4�9��
oxY)�.1̖�B���B��h��������<��P�00[�	u��
�.�#�Z�[�,m&4���0�ϕ�j��R4ޭj��c^0���� kG���4Pn����Mb{Y�Ti'�"�4<��Itv��7g�1=�6϶L�ڐZhzA7,�Z��x�3ko���Rk�3�A�i�Ӛ�5Y�P��r���/w�^�/A�M��f�^�0y����`� ������k���{��+�Yɻk񷄉I�M�qj��ۊ��fq>�%z^n��K����I�MA�/��I�.��|33>K+%ڊsSrqL�:qK9R6.��L��[}������!������Ns�d�֖����z��ˣ��<���]�̝�����̘�����������z�	�����n��KX�6��Pl�� �Y�7���zٝۻ�FK���/fQ�pA..�.�"�hue���/&i�o�C�/��ʐ�܋��s��0�paK �#ٽfX�Tb��R���˨�/�������j
�����R�+��.�1٫Ļs�&y�\��k��P�g��pr����}�� �xkǭ?!�7F%�Y�|F..�gAT�Κ�|���+���Y8*�F�[Rw��{���GH����9���jn&��6�k?��A�:bN=�EG�"�S��T,폞Z�}2.��2��P���:o��0Z��C�`�8�I�0��k>}a���oB��[�T�����B�U�𸓬X8�z����Hm	�\\Q��y,�P�9���+A�F�c�˓�G��r�Bx�D�6�%|č�B��s���;
X���ܪ/��?��kC�Gfٱ��#&��Wea���r��*�j���r�e7SC��\��0~疄�\{�p�&���x14�n8K�k):��lg��.]t�.ۏ�V/�<�^"��sl��mvb�J�tY��jv�~�+[���X�a��v1P��Rf�.�i	��ݬ*�yV`��g"�����w�w<�6��n�Nġ8BEm��x�̧��1�8�T�Z�Wv32�v���Ե8Ӟch�*މ�����f����hO~(��@��1��D�@�q���<Ч��ζ�.P$ǚ����g�ї�8?W�jl��g� �I�)�dxԮ��|E�`,��Z]�Hke��MeU����I|)���nr�ð��ޓ���C�13���PhcW���36o�ٕ.�������NJv��$vq"�G	hb���2<}�CUb���^6�㻥e6�B2nkawL^K�a+�f����X���9��Mh�
M|�,=wʄ��!8}n��Y��ޢN���0��k[b�V��=�2ˠ
aʡ	�;�tg�`��Y�Ѿ�x�����=��oadS�hE���̖)��S�U���g�!�T�W<��_�TH��y{2/
R|ܱ��������A��j�c�/Z�څ�>�٩j��z	Ba��C@��I�]K��˛=]9�Z}�����*ʮ���Y\������P��2�b�.*���	�F�+���Ӂ�+�)��i���ąt���Qr���]!�[��)���瓗�����Z%�簸�ǔt7��].M������&/[�u闳@3����5菺�d��F*�0��g|���w�#A��Ι��EK�DmOuu|>��5�r��"*�$�"]-S�ۨ�p=C/0͕r�,�ї�Ț	�Q�*.�V�㓌92Rv�xp���)P�ŏ���x\l��$5O�3�պ��ûi�U�;X��􇡭� �Y�-�F�0�ͬp��E�&��wmok�a�{At���Zh�2w-��� ͜%�A�k����		���m��Y�:,��3Xփ2�����e'X�)�?%��X�g2b�.9j���0П���ɻ'�ڢ6�}][Z�!��t�s�bC��`L�n/�ny�}�J�O�ɏ|�v����	�g�ql��ުi�{n^���c�<�؞EW��qG-W0�⌖K<�y��N(��]'\��)����jH+��5�C\S*��k�P�2��G�gc��N[s^�3�;����@{�QP�Y�q��Hd�Z��:C��v�1	��D�jsu�GNu����T|�Twru�
����ZmSb���.|�L��_��yP�2
�=Mw�P�����{5*�E��4oE[$��Q�p��%.���p�=Mt�]��1�#\�o�<f1,��m�tyk�����?�)���ϐ;��k.+Y�����\`c47)�%�TT��&�^W��x�1o��߰����pLN�7�aM[u6�	:���5���k�-����F�c��-/�V"	�N�/uӑk�5s8�i���y�ٕf�����;�����̃��J��L�0��RK����K���Kc�g���x�-�\��<w��Z&7}5�y�k�{XFfK��v9;���!���c<T��f���zja�7rB����Vl��Ə/;��.!��;��~��, t�ڣ^�1��%6������8�YX'r�o+���8�_��/�"��J)��K��P��%��꣧;��X����s�a�/�X�{� >���t+�v&��)�9RXg�oW�b�t��>c~��x���Mt�q]�P�o��� ���J=V�B�����Wt�L�$��d�8��nbHo]� �w�MRBP��T���-�g�'�w��	��J��~��2b�k�[��۵Y*��`f�l��s&%]��KpԌDk���zα}����G���=�����~�v��P35��ߤ1
faD�k���7z�bl'�F��<6=N�;m�1�Ҹ��<�&8��Z�2�'wT$(��v}���������DD'֯OCk�{vi����7��0&(G<�0Q��=��_NI;���!huXsvVa���`�� u�~_�G����m�w�T�v�p��Y�sF��i��ڰ��1�KY�g~{��B��z�]*�p�-��]\T�{1�P��M0td�������&�mj������Psn��CU��7���#η2Xq^"�tj���#�q�/fbw�2��00E��m2)w�Kb����4m�ܬ�<��ò�i7���W�7�J~�T�+��ǅ��5��>�9�?'�(~}����0��B)����j́'�PM��]��e��4U<����$[>އ:8��|9���?���������%9���{��?a�{m��6ό�ω�ǽ�YT=���U���n��|���H�J`v)����㝁��t�1=u�������O;Lk�q�͠^ �\��.Y	����P���<v�m��v�	�B��mg&�w���곊-�g>��T���囡g�nn�;��]8��U1��i#]�Y�p�5S6#L��-�^�CdT�j����	���۔r6p�Y�LkTOeP�ByH�Jb�۫T�@�k2�<�Q��h�v��ݛ��[:2�R�U�;̯Z���%Pp�T��ԛU� �)���g!��Z�}�ܛ���v�'µkM
�7C�R�;'�YU��e`�W5�AA�U��^�#(�y����Ӗ���=������`-���|�i����r�o�����>��w�C[�Z����������'
��;jd�.���ː^�\ܭ���K�5��I�#���{�x\ܩ[$�%*��W�>�w��ǻ���
6+�������v�`��2>�cR�Mn�n_�L��JhGi*=��(A��m�r�g���H�iW��� ��S>C��0B���q5�ڗK�1v;x��=̜��+{��n`���Q���W^P�qM{����fd�-�$����sC�9v�4��-魘v#��G{�r��%#�Py�����L�~�uW9�ƥ�-!ɋ��3��c�~S�wVX�P-	l��f��z��Dъ��Yt��N:/<N�^/<�����En̥b�z����q�GZʨAﲞ�[��;W�U�<Ƙ�N�aٲ8�8d�of�tq�cΘn_��w������L�����
)��!����!{�ψ�fl��]�.o5�"�y��ɨ������C�Cd��bkWP�J@e!�����O���p��X�5M�\�3՘�c���/��+9�p͜E�Oc�����d�/��X}�~pS��C��[t�8Re�ݕz�v���W�v���Vq�J�*��F�����2g������66f��i��G{ccF��	��gH�
���e]f�x�!��%��j�
(���D�QM4�4�]w+<^3p�hk0,���Qb�&7In�)�9U2���2��b��سj�t��T�WuN�n�<�ȉ�t.�^)���^B$d�J�����=�ҝF��z5!��U譫"s��lr��jĚ�*'dw%���y�N+�Ɠ��E0����k��{P�*�^�b�P*����"�\gN�+�ґ����~h����f%����	ݜ#rs��[��i��-�8�fDe�:���a�9�r9�TE)��rE����1��t�׃f�	U�C�dO���5���l[O�.�
��5�[t�\�_'Y�F����a'���J��n߉[4�mxA���5����(89�"eݔs(��9�*�[��hFn��o��	�U��8��o6�B�c�'ԓ��x호�{�.j��83�O�9�xн���dU��r�P+�*=�Wۧ�3�l�e�3�1�b!n�X,�za��!#BOGg�);�(Z�'�����z���O������������z/�n�s�ͫ�S��*>���顶bܣ9�i�S$��.�tR�9�x��6Afk�o� ���b��V$��^nPB��Dl���BiPn��F��kmյٍ���{��	�+�}W,X�и:�1@[Ҧ9��l���*�Sq
�9��f���{u�&%�Wt]�%�#��=�k,�CdD�ܡ9�,��V6�U(Y��y;rA�kB:�	ټ�hHRxt�椇wU��s�i�I��qnp}v�]D�
y�)P
�#����qR�o�C��N�ܤ�
^��1�9\�w�/3�FWR��.���Y���[�R��*.,�p����t�^��6����ٜ�j��{&\�[4U72��LʽT�=kV:��āHBwq�uR�9���qP�ٙ���tP�W����A�5�Gڻ�V�qv+d�=��co����A��1���r��i�[7z�j�ns��9�f�8�n����T���18�%���E��<�5���سh^vth��;#�%s�&(u������#[H�W؃�v�v��%^�P�F��w��=�n*SvȭE�F�Lc�]09.畃�z."�
v��;��;��ή��CKK#8�QP���?m23*D���l�rpI;׉ue':�J�Hد�;(*�&�։�a�a�֋��M�.�P�ɢ��o4n�d��8�5t:��ֳ�;�����Hrok�ɿ��ɪ�\��^V��,�A��f�B!�.�ωc;��&������%�`�o��R�쒳���A�x1TΞM�����1K��̙VԞm��Е��������b�X�$�~ȗk��ӈV�ڱ{dN<�
��V7l��m̑f��J���+�b��V5Y�ŽDh�ז�B1;�)gUά��ޗ�,\��O��Q�;Da镶#�����,-V�}.s�v;���=�L�� @�ͭj�vĺ���	ZL�y3����v�ٶ1��5j�����,���Y�Čsh��%�K4���ى\����w}:��:Ɋty|\���(̚w�V�\t�����'dNI(y#�3A's��������*���\�qaƋ��K٫>̊��Hw/�	u�]i�*t��#;$�s�_	�l��}���R�_^�da�*p���%u��|�꺾
iz��AnU�Ϥ�����٪̦�)��J0���b���z`3�orL���/Ob��'}�Y|�^Cz�zN�� ѱ:��E1�u���<�J��5�i�,��"4������`���t OFQZw��A�z�]k�!�_U�*igvN����Sgb60^fv-��T����}�RX�n�XO!l�{��U�Ю�޳e��m=�0E-�A�cT]I��/�E'/Oh��V|�.�ɣ�ٔ�c�_���s�4�g�G2
˺J�c���dna�+J�Mf��%��շ�����6���RJV��Ӭm�l.�g3�s��c�GCq�/q����ǗUx���kh@�t�{��u�<	���UJk�	}����&٨���ݚ� ��UbtZ7Xn�^ƪ�T3O�Lu��v;:*#U��"�Q�l�m���9�)��3�+���-��
��Z�D��X���u�y�IGcS��E3Ί*-�Wv�f�jo�1%ڈ�3>X(��&�������(��Wv�X����TPWl�K��P�SHm��Db�O\�lG��"�Z ��"���R3�T�#�L�EQESA4yh��G��U1�4�+�A��#F��� ���i���X�����͊��656<�⠠��bq���+����MG���눪���i���8�;t=Aѣͩ�z���LI���F""{�;cA���:�#��kx�V1/Z(6������ɢ���]:�h>u��;�k���DUPQ��颾N����c�����GX����A�b(����>|�B��X�C�x8K��TH3&�f�t���\��pp�3U��e.�ZD��Ü���=�q��jlӲ��2խY��O\*CLi��~`0�m���x��ѽ��$��������}�eQ'��ե?Ic3�����SumI�p>�ƻqa�8��P,&��t�wd4ʾ7]4�'d��_����Ǳ��!��t�-�\k�/�'SOf���Ꙟ�"ꑙ>lT3�;#��`l7��H�U)h2��ÑVѩ��`.M^DQ�����"��.���D�+2zs��-���2G�E3��O�&�w�ّ\d��L%��<l�"1�M������Q�Lw�!v��q�훘�VF�%����y a�h�m2�t�x�T�٩;��R���v���k���鴂k�]y�*�%�W��\f�h�W�6d=� ܪ^���"��u*܇]S7���.H���JS��ʵ��g�,� U6�t+k�Eۍ
�N=����!����Ut$h'U�^Y��-����G�\[�7<Ԍ]{ْj��#;]A�@U�(�����SF��Ɏ�������Lt6���@4`�u;��G*"���jP�ΰ�n�����o$28_'��JR�v1����~���vΜx=�o��;,<���u�����9���܈KN���O�e.�rU]���e.��ȼ�S�7��h�P��0��OѪg��3�uo�9�'y#~e�z�We�"������M�;��ڜ�~��B���`G�S���O�/y;�BZ#%�\�L\�+ǿ�4F\e����ͯK�V�2�"z}��sӵ��U�]"r;4o4{ݽ�'�*m�WEM�؅�;; C�Kꉻ:#)�Ϳ��{�{Q(�T���h��cp-���3[�G�t4ᛠ��!��5�0�����G�Lѫhs��z���i��h1'Z[���G�����{�,-Ļr�7�A�>�=�s������=�m�tlc�\I=X[0���H�lZ��J����m��n�p�hl{�ꦚfN/w�X��1�3f�����R�bg�|�!(�W��<�֦���K���G���7Ne���1}�B�Wt��`pga�z���vl�5d���w��vh�qm��X�]F��[Etf�R�e��:�Gy�C�j'�کԺ%�nm�)j�mV�C]l��b��/��/��I{�t����+��vN]���`Ax���g�\�]K��gC@� �=����6�VH*١e�<dx5�8��aQ�k���k�K#V񚵽"���!x��˜d*5n�!���66btL�mog>�]o�Cҫ��U�W�J�J�(q[U���������n���A��͵�ҹ`���̬�j] k�=�Hý�0������v��f;s�=� U��T4�\�)��>Rέ�M0����WO8&�i��P��'�z�o*1���sn�r���6�%}�ס��h��wn��|9v�/+v�ȕՔ#�D�O��3�K������-���݂��V���}]ܽD�-�N���č�r� ����/qX0T��6k���]0����r;,��WĽ���f3wSk�L���
	OFZc̑k�����-E>r�"9���U��Vխ
Vd���o=^��6d����76���,�4Uü���U3�j�r�\�1�k��m�`��c�Dkes�5>d���;Ә`Ըs��Y%IUY�tz���ǻUhb�F�;���̎��q�|�G����u˝���P�٣B������1g�}�Qbw��?��^���6n�����#�����Hv>�1ڍd��F�wb��ͻkn"LnU+7I�X8�F��؜��
`�]��˦��������/��5�y'��"g+{)�Ւѐ�A�|Fq��<�����ZC(d�7d��v��4���;����|��*�������\�GH�;\�����뻮���U���ug(iM�R#H�	+,�^�u��N���r�(����m]�"iU]��f���7 #�4���` ���n!4	ي�ț�'�p���-�9�n�Ya�T���-g`,ĶǴ��K�nM�����=}������(ov3�٧�4�z���HE@��ͅq����/kI��uש=^��h+�7L��-�T��J�~B⹩�^�H&���/8o��<`�� �t�L���8��R��r����1 f"͘=��oK�>�@����Ӿ:�2�7��;�Z捳��z 6��|/l�N�f83��4@<�8�D�о `]�:��F�wG�n�=,����;�^��M>�A�Uq��Sۼ�.#���Ii�8��-���q}��k�BS�гc>h����cw7�#��k�Q�0�(����G6��qw4:-op������n�;�:��(#�E�e�7y*&�I�f��p��=	%m^
���o�����Y5�`�n�$a�CM�W
<:�Ǩ�yԵYD�K��ő�Y2�����Z1�(�0G����������j��'�V�mv���a���5kOgr�0!M�Fl�ᷳ�,�t���FUG?!��f��k���Ӷ]�C���ڱ��`q�<{a��ԧ�8��N��b�{2-���FC�f������Z��������;��3�� ��Hc/j�-ς�~7smH�f7�?a�/����R�4����w��9[�p^�Ox�qx]�O����^g�7^F�8�v��
lO>�k��Uv�G�d�\c( ۳��%LM��}Wq���3͸�h�)�x!�J[@��SL�ԿK���"(��MB��w~��ͤĹ�J�y�4�y�yӵ�L�_Q��{g5��[/ s���֯�K6ߙ8O٬(���9=��*�0�kU�6s����\�2up\@�4C�3i�|a�#���5h�8�ޖj�����>x��e0�ɧ��2*��bٸ��e���j��t���=��Kd��Z��K�l�wnU!�M�z���8*�����VOE͈۬|Wo?U��"�vP&֕w8��-0�"�=��? ���h��F7+���ٵ�kb8���b�IW*n|Mڢ� 4�B��G�z[W3��e�aj��u����St�Ex��Y/����Nk������xv]��]`�=���@<o�[�����H�[�&�{��F���v4�Om��l�R�t\�n�{3�}��Y��r��$҄g4LF�)�Q��5�����@�����U��a��e�D>��-�M��v���sB���^H�f|*���RV�ܷiW�>��*1��>i�fE�Xl��۩|�r~�ߪMz�~��}~�s��j�#;$�h���x{G^%F裉��Y܌�F#�#ق�����Rы.�4_n��e�t)�T��Hv���K��<R󖿍$��9�+�M��6��
�̅�����R�U�T�"���+��^)���qʨV1#��!��T���"m6����uu��0n�跷 �^��~�>'y^ٸY�8Z{�mx���͚fuB笇��&R�y�T-��׶�������N��7f�&�;��gy���:��cޑ�O�GD����g�v��G�)�M�a��Ɵ[G�\��Vk�l�N7+rW53��
�)g�۰�% cT�.a�����ݹ=�:#��S��IDd�$l��i��Q�z����P���1���[o[��x�]fN���	�$FJQr��J6��k7!W{d����sŲf^�]zN���Zly3���GbG'(����ͣroQ�y�z)�̦DU���p��%�|�tB��K��$�ntnN�^V��I˛,�$0�]��ʢ��U��\i�����%_h�D��C�ۺ�)�~��-m��~>������o��a��3]��p^��v�f�[���|�*��k6o۝��N.I�y���!X�1/�88�)(��gQ��*٘N۩?l��6������;�Z��Ud�j_�ƅ����)�s�����ʵ��4�!�!G��:I�s��Lӕla�t&��ܢ��Q��Vյ��3���s�wx6�m�;���$���]q�T�<��+`r��Vi6�����n��q+/��V��\`�+�϶�.�|.����P,�:�1W�T�L��y1��.7l��|K�J�2��`^��!�~�7֟��ܪ;�\'Vi<��4�w`���7ȫ��P��u�n�-]�|Łw�e�N���g�]�������F�������X	i���9�ZdI�a�jX2FCwP��g���Zv!WM�$��͕��/1�+�ᇛLL �;�v�>3DxY��O"g/�� �k�殇���Rz�"��|������{6�?L���g�婡�<���u���Y����Y�}�bq<Y���0���% �
�B�d"�kf��fٴ�4ݜ�7x�����k�{Jbk���ؼ3XK�D�t����������Z�**��ʟ�U��8��:X���26�}�J�gn%��zX�ɨ;@6�'���5{'���y�/e�])�'K�̖���l���t[����3�0�r�j3�S����n:�wHm_.m�[�v֜}7w�K�Rpm�:�:�84���c�����y��WT�z��\Bw5p�tUk��z�f�f8<59�jt-�x�� j�ˤ<p���gÔ��ʮ�;�䉸['�H�)]B�䂮���xˤ5�{id�
liݶ�EM��WˆTX��H�����A-(��Y4�畽ȫc2�vz��rfR�kI|!�#��\si�Ӕ/C��&�H����5��Y��x�̉�kԷe��QG$�۞]�r�����v�ƫ�����2��µ{��I��b4�\Da���"�!��u��>,�=z��'O<��[]��V?mI�Fj.^�˒�s�Y��� �C-�b0���-t��]ޯ@�ب�=��sz6�ωm㘯I1i�d{��ͱ��Z��.�%�E ��]A��Zj����*�%�i��- �d��hi�8#�d�
��C=3��	����ӝQ��7l;vTϲV"M�<�sA��<I����V�r�G��VAl�v+����6����u�&�*�nԽ�ܠ��i�*P�Yhf>_�%�3]݇���u�Gڜ�+-j��+��r����r�����6�k�4.�5���s_>�5m�����6I��Pc���v�5������f�f_q��ۑ��^��D>�X1)=�_�u��bz�P޵����9�Lf�>ӆ�<Rd���yKN�m��nz�UxE�ҹF��RS"���KE�{&��lg��=�j�tR��|0����om���ەU����.�'F H��L���
 _C��"�S���U�t�Y��#/o��1��&dWp/>��W9M�oJI|�=�Ʃ���"s��F��a��5b�]��G�3�z{/�"�I�
Β�V��d��b��V@�k0�{���>e}.x\�/�K�G�t��Q�ld\kV�;j�uʲ�[k.��c*��e�+w��W���.v�<��R��ñ+E���hc��[>���pّɽs!��9M�er��n�H��Ǘ�������}>�w��=�^o7�dKٷ�2�a���jN���<W+"�q�O�Ν���V���ِ�+�UV��Y��y���Ͻ��+�[M^V�;�6����^oGjR9�"u�y".j��ms��
Xyb�Af-��j�+8sKյ;��oOU:sv�䋊�j�k�@U���	�N�ck��.c����;Y�����q!�����&�p�[v:eݾpb�>Z�_kJ��`���y:�Lu�����f��z�nc�V��c+P#����\���4��'�R��+w��8[u�����1"�J��+F�86�Wu,���F��K6�0*Fj.��Vvd�to�j�J��+2��$8��Q�+)o%�;�Ը����n��;t+p�^���a�[�-`u�d�'Aѽ6�c@b˝��&����f��k���Cy���Q��b�b��S
���r�T8L� \Wf٥���x��9�$����:�v�a�9V�*�v�a� (�H&��d��"�	��8/�ɚr��Uc&$��{p>B�}x�έ_+	��#�k�z��K1���;�{W���EH��X�iU�+�Q;�ȵָ^ij�,��Vu�\pC%6k�f��>F�̫w���wi8Jќ2Ft��Н�e���:&c1Lb�B�Jo1�+����	|��I�Ә��v�،�v���/��o\@�z�!c�o]�Ǜ�n�d��;X�����+Vc�n�����@�9GI�29�F�����t��}2�X���r�Ö��Xণb��K5��i�M@cS)�:oc�­G;�e�f��=��0�pujޣCiُ�7�W6�zcݦʰ�y�����E���gu͉*�,E}wՌ#oj����*(u���̫C�I�VD��̓)���H\�j)B�l
�[̎�$w�z��9w�Nb��SwX���*�ԭN���N�Z���WW�����Z��0�<�֬�wJ,n�ֆ�/�����K�r	����Y�>r��R:�!��M�D]D��w�hn%��:��gl.����,R��"xNl�\r#��Q�C�m��0��A{�Ggi�T�Awm�(�Y�8��gb%��Φ^�;:2bR<!�8vt(I�� �f�����4�����y�%��w��&h�eKt,�R��ꊅ:��	�@QX�(>W�(blk5n��g'xU�74�"�]�%gf�.Z�}��o=E�ȳ"� ��iA(�+��s�'u)�����\�><1��Ã��<������˹OD��8������;H�s�����h��&�s�եb�p3y�^E��ۭ�D��Ͷ��kq2�.��WH̫�j��#����M2�dU��e*]PK:���qv�s��}M��Q���p�|�ƅ��õu��)-���g^��f0c��	$�b++2�s9q�=xJh�
�P�ze$�$�4I	D��UJ���b�&������T>lFv�I��AAWZ�m�uv(+�y�<E%I�MyMkOgy��A�<�� 5��8���T�h�v�Z4�EEE7Fb��6�'^]�đpF�z(14��Ѫ�yuAC^^A�I[k�*���IQ�TQTg8��v֒��h;[G��^m1���<�Ocˊ���'m�=t�U4S�5vq)1S�WN��
 �+l�G��&�%�u%����:��+F����1I3�o<��(<���@b��וx�%�I��w����i����E��hv1UIQ=�7N#�y���4�%M4S�u̱	Et�(
j���+�DO0h:�mh������ϛ=�S�=Ƙ#e���#AR��F$�+�4���E��LE]�Fh��&������|�۷������P��>���EfB�C�ܷyX���4�W���ºa�)��������#c-L����Z���j���}n��f��IQ�2XO:����v#%S�o���d��K:�"�[��������p�pK!U�ONa�߶�hӕ�Ek̖�/{=�u�U��<��0W��w�qƳ躧��pC�Ot��L�g՛�'aN��j�b�Қ��㍷&)��P�/9C.�Op���fDGj�&v ���*��9��I��H�Uu0�2��R����]��>u��Z./�p\�};��,����,��'dV�?l���Mo׍�p��T#�{ؘ[����Ȁ�ϳ0�ű�w���b��6��gS��b�H螖���a���8d��c�U�$�����=�O���́��mx6��E��T��:��ؤ<d5�O�D:�`�Kvr̒�옛%l{sv����p84��S5�i����M.��ީ��/B'7j���9w�W��.cԯ�֧�q�'�p�MV��J6�#���Z2�Zÿ��acok�G�l���=�"��[O|�W�t�Q]���_�K?>�6T��no�SPd(n��HA�&țp
�ZP�WXd���m��!T%���{)ܔ��bc�=o�	�^�u�^��9 �B��˙�9W�;�~��7d�zUt'T
SS�d��P*�J�ì�̔��|&^�Vu[a��U���0�p�Ƹ�Z�if�S��mK�v_�ޙ����rr0��YD�Rum�̧[��6P���P�Y�q��vԼ4���ʌVg{Y��y��u�i�5r(���vE�9Mr ��3YGLn�]5��f)�'��3摑���:J��a��%uez3�f�r��u<
138�B�W3�r�q�|�u��wJ�`�(ڃ�H�8�
 s���LYL滹�q�I��D2.7m)�_�i�IP+���,����:�K�J��,;QY��݃��Pͭ��hõ}3��eZХ�i���v����j��;�n�_����-�{�͂Chp�.�Gj9G��ŏj0wEEuWH7[��s&.suR��!DdwP��g;�̈́hv�D��o,;{��b�j��r���B�T�v��d(���@��u�Q��'�����Nڼ�j��7�����'�A�P.�c�nRL��9C9���q#j�p�r�CO5͸>�X�k:p�Ӑ�0�4h�����V�[h<Μ��P��{0�{δ����wK/�gK������K�=�ӽ�LI�ƃX^2O�]l��v�{���u3�D@��B�^�卤y��j�㔙��Vބ���yu
���ay�8��u��x���^)&��`ɫ/{�[�HoxՂ�>�<UM��u霡��OM.ȀS��֠=�15�Sw�0�ǧ	y�]�{6�K���`�����V�J�w�}��@�%_�[��'��}�/��,�C�u]�F)��q���^ƹ���z���qL�e�1��j�;c˕�L��0	�Bz����N�3�=�9�-IUj�AWtr�m�.���6�n��k'r-�6w\�M4�2I�wos��u�x�M�W�S�r4U��"w9��tK�MYw�o�a��&���ᷜ���Ί�n�+i�Uԥ��)ۙM��C�/!�A��1k��	35��]�w��i�p��wʷ�m-�t0M�3��{��<�x��� R�d�-��hn�x4�^2K}�4��m���RuG�/�o�������i�T�/��ϰ�+��'ݷ��t栙Z���o7��<�o1sƤy���	3��U��+o,�çm�T���e,煛��ɢ��(��Y.VU��$��|Y���O���g3i׋���}�v�N��#��N��ح��5�`��}����u	�&�l?�L����Xr�SF�w��2�{8��Q�3�u��#څ7O���6�����y���g.�5S�n�A��\q_�n��q�9�>%����-P*����q�;�u���!�ԁo�\�l,�����=�G� 3�~}Vż���E�Lf~���B��Uly�WG�lbͳ�ۣ}�;og1�Ĕ�M��K��P�oob&7�f�&*��3{�̆�N�b�͝^y�7�q��p�A�S\v���WcP;�i��'j�����t�z�S�[���g�.q��{�����_wC����S,q}e�:�Dę�w�Jbw�{"��ˌ���j�6W����(Υs�5cEڧ2�z�h;z��D��*P������y]��ⅹ�wYe���x˧�p������<��ˁ��1@;y�����3���ݓ�6�`*��mZ�Kz�xu��]a���qu0/P�7�:Ge�3n�=C��.AR����E��K������]en�o+ l@r�[;6��l�:�@	�+$Q�)/&����sA�����V����B��)���]k.VS<y�.�p1!��[�H�gu`k!�`2���k��԰϶#�wJ\T-��)��Khj��:��I˜K��dO��'5G%�/�r65��n�ʑ��3���ΧmT�%x�b�8'�M�uٍ�&��u��ױ�;��)�,�mi�����1:h��+	n$�J�6v	�YZ٧)X��sӴ�f<��F�}d�y�R}�\�rJ�#�6�2°,~�gj���u�:tC���K�ʄ�@��<�+�tWr���S8��/^.yqNO>��U��6�l����>}orx��Cy,�r6Bˢ���:tdc��F�u�Y1���;�}�� ��":�d�Ӝ?r�z��S�g��'�[{e����W��G�}���1����7f�����3�AF�����<�����`�h�{
�]��ӂf&�[��vK�9����ҫ��k�+��us�s�g"���9a�@75�g;ȬͭB�� ��ё^A1Nbj�wnM}y�^��4	0�]7�hv�����wP{z�1Ĭ(�sO���s�l5k�v�dϠW��S6�͡���܋��;�1��@��#G.�EU"����d ��Z��u��7n�'�o�wN?��-���L��Q#HY:��4�}���l���sm��:�4�s�lg{��g���_5�#~O��|d'�2<Tt�V�7^DdΫN��RwZ�h��O��CSS���w�%�v��Z��BZa���N��i��ڄ?��
>^[�SF�S�~�I��e눅��K67"�LгZ���9ݗ9A��ɹ�Wʲ�̪	cG��l�q�����N��p)�8�m:�jgf.��۩�%�Q�5�mj-�9���!�k�{α���4��58��-��$u�Ǥ7$����~d	]YQ֢{�9�"�ܪ޼�l!��[�5�<0#U	�|�o�и�����?n$l�T����Us�J�[�Ng�ٰZv�U��}ݙ}��-����4����3ku����jI��+�J\8k�+Ղ�n��Wº(���B���v�#�N4)�x!�*ݸ;8@����r�6��ǻI��N�c�AC\C��V��fV�C�7�K��3:L��H2��Ƒ:�=�;�15�C�O�q�����U��U�~��7<1�=�Xd]�qH����������ö�ȏ��#�u�^��9���ɘ|�O���nf�l֢wU�7�0�m���;��u�}=��(�-�ް@YYW�:ׁp��|�����ue�l�3��m���Ӯ5�v46*{���re8��9Xk�1�34�>+�1�&�O]6��1$��Ǳ���m�h{]U[��y�0;c�)e����p4[<M�TuIA�����8���G^�=��.{Ɯ6k�S��@`��]��#t��R �b6�9�R�Ӗ�r��_k��>;Msc�'~�6Ył�Tz*��a���_��e�ٺ�l�c��ugɁ,�*n�v �?��t���0j:��i����z���9���C�B�$�$�E�c�jn��U@-�x�mMH�@�j��Rݐ׿?h�}�qd*�A;jT�a���J�x��t&�)�w��"��x$%祖|wB��R���(�O*��c�Hb���2��N���@')VaK[�����sk]b{g��p@�|����#R�ۋnv6�&�k�!{8���t��A�퍪�I�+���Y�
�^��3E�����k2��
���p}���?!l���a�2;�v������U�u�r;	9WSd=�v�\���|/f�l�v���;�b������+�l��M�����j���F�U�k��^5!��{A�/Tf[w��M"��KNɦj����m��gu&�)�nԻ�2��jޡ�zӀ�&�Ȁ&*2�n����mՊt_(d��;�JE�縆�izο�չcƎCm�otVkE�)�RWe-��w�wmXH�!M�Fv(wfaW=q>�Y��{���)����fspʆ�ն/s�B`���O���;2:�\�lC^)���2������Y��4x�c&dν�FN�==�Y����؛�@q��FlȀ�͋��[<"�>����ߌ�磬3 ��铎���N�V;G��Q�[�gÒէ ��o��u�Hmvm�+{^3N�jE�]��ꄐ7�K�%��$Kh��G����R��Fn��Ť9�u�1Φ"������D	Go�|�P���攚/�lS�4�t��ӈ�j�w�)0PL��Q���v��Z�
V�����t��v�!�!�x�ȋ*���ׅ���u�����ھ�u�K�-b �I�HZE�N'v<�<WTȖƹy.���f�Z�(E�
#DL��QA$6y
������F�a��
,�w2��R��y�+����
��G�栟����m�˽yKQXgJ���ewnlC��iȚy��j�:�u�A�ؑ�+�4���Y���]���3�Nzc��p�g H=U�V�5hIEὈメ-���w;�.�a�=]�`f�ܻ^���v����^�c:6�j|Kw8?��pK�I����h�7ugN��}�H-6����J���َj,3�zD�!e��`��vD�N��*�N��;��*o87vv�R�N�Ns��[��<FG�
��V�n�ػ_r�&��}y�SY��{~�\��yVϻX��m�x�ʸ��'.Vh���²i�q��'�˶�M�c(`�\_1ˏ���R���s�$��]X�E��3�jYR��{@�&%�}������hb��Z/V`��A$Z�׹�x�3L����u�����1t퍼�ӗt&R��bvZ��G�n���dգ���W��{�BccmL�i��:�V���A������8��u�<N��j��V/:�>�ԨL��6e�jW]����v_�l�@f��Ƒn�-"o�����K�tT'�Ӵ9�STLG�U+�G����חkl�3��c���[�]�#�ݥ]Ӓ�(i�Y4-�t��:���oD.ۃ�}/-�#��`ĳ)կy�n�o���6v�1�U/ �9�cm��@�b
�Z]X�@xĺ�x�N�i;��d�ɹ� �jʡ��ϊ[�M�׾Dd�HY �m��6�庶���
�������;�b�O3��m.�}]|u>�V�#�5�f/\��0�L��硧%�����C=�I*�WW���e�3�S:i�V���{/�ױ�#�^�`Bi���7I��j�Sj��pơ���\�[���P�z|}~^�O�����yy��������۾�O��"�GfGJ�r�Q�t!��-H�T��G��f#b,��&ֵ��󨄧0s�0�V�fWc����Zc_��X ��A\C2��<qS�1'�D�U�n�]w�.��v�_q���X35`k0�e$�b�Y����' �h�t��WnxE�r88t�w/�N,<f�MҦ�V��:���Q�H�\��s�h}H��	�s�u�}v+�1%��Χ|�L�J�X���2��{o^jn��yj�-�ʬe�[��'��f�g&�G��I-���-}��3�C8�>���熶�ͱ��b�tj�1�}{��á�G%��Q�:�����z�=�����*NӍį�r�H�������X�T�N>�o�POh�:ad�V�ep�IL�:(���+����(�{�
B��ڝ¿c�+,7�v3�ƕVG٘��Q�ۍn������/_;��jO���pO!V�qRw��p��t�:HG8w���O ]��X�曋��i��K�ǳhgu	�p��<&����A�_++�S�Z��Z�$��P�:��K"_j��']��(r��iv�!x��V���*�ߛ{N�ݻx�[�]q�����S��&�|����vpG$�%��qgjr�Kz�VvK�b"����n�tA��αZX��ķR��2�ژ�p�0i��g7���{#l*�`�/.�����ʂ'���Й�St��AQ�T��o��_:�5x��k=�����ܫᯤ��@���0Um�t�&�Lm��uk���藪G�����5�d�����At�nn'�]wc�N��7gtJ2ecY2���ǹbJb�7o�e�R�;|�K�V��M�/@�Ow'fGV�d��@>8�b�[�I}&���!���`�RY���Դzgf
^����]h杬#�z	a22���酉�l�^0�p���n�]�ңʹ\Ռ���3���$�C�;�]@˕O�=$��԰L�fC���7����b��C@a��o���\�G(S�#F�$��D[TfȌ�	��\y�wr��}�����e�M9�ݝ�ւ���ږ�!��.��V���u��um�q��� ���;<ɮ(�?L�Za����@�e=���f���h�K�;vA��p��{��W����Te�4Ν1�p��n�(���� l�v���t���c��ۗ����ݸU��Gkqh�By��i\{
�*�t89���h���v$Q��kH���:��F::w�l-���n����;x�݂Si*����j�㵩��Z�Y�W��g3jL��j�B*�K:�$rx���j����azH[O��v���eE,��m�3
�ܴ��\�g�X�g	�u��%X�Bf1�3��p�U�N���xl��`�t&=t�mgu�mcë�>����)m��Mw�wƚ�6��jU30�t�9�p�W:iڅ�	J�٣��=�8��G�&
�&�F�����"�b(�Fo6����6&f����>ML���CGF ��1E��{�E1y��41%��DD4y+aƌ�頢�����4�m�"��q4����
���c�TIE%KE�Zm�F���y��'�ԺPv۱F�"��w���ULU>J[m�f�� �h1�DCEv��M��;�!4HR�0Rc&��$ѣk�����·F�ZSHS��tww�&���NػbJB&�6ɻ/QUu�1)T:4CKM4L�SMhT�ьh���
�q�QU&���:(�;b�(��t�cl�tF֠������TǙ1R�Dhx�u�%�F�����5TM��uZąW@q��**O'I����?_m���N����i�����v塉�ˤy��fQ�����W�(~R�f��R��W�7XB�0�t���I�Wb�o���u9 U]�v�^�o�gӒU�RX�*�����Y9���iD�#�	*���^I�bƐw�ęavX	.�3YF�򷳖���w�
��wl����ÅKU	=��|3J��r%i���YWVW��E��9u��$[ �N�g�}1~��2T��h��r�и�D���^��h9�q�E�㧈|���y�VL�E�<�9!�t��\f�c�iU_�F���/7oFV�V������:�?��v`�}�<�[�Q�N��u�b��P'M�����N��)I飻tM�"�[��އ���j��OI;&[�h=���M?u۾��A2�\�M�"�kʚ��������1V�?t�3I���b�7�};$8�۵ˆ���N����i}h�y��Vx�6��
-��]*�+����B�V)��(w���p�q��o�G�U��~Kk��Ѵ���6���F�3�y;��4k�
^ӬҸ�I;�����ɸa�+ݲb�e>,X�]���h׮����%��hԙ�j�Op��F��r�[�O���
��]wJ*��4����c�R�I�/�opD\�'{,�%ׅ�!;����/�h:?���NT���C8��3@o�)�9��#e5�`�W�;M�i�B=yLgSj�����U	�7W7�1Et\Y�g�zZ*h��ǘ�k?u��(��l��Q��!�CR�H��J���S���Pu�p����l��Q�k$'=X5<v���N1��C����v�6�k��}U33^�]�CR���v��椕Z��j�+���v�e�A�<��jǱ��k7L��K�k'�H��b�i��2k�v��+�����C˳�𔎯+I��;�ܵ����u���7 ��|Z}�����ܧ�����e��!=[G7�Uw�� o����Fٹ����e�H�q����WHA��sCga>)�̲�mݴM����c�뒬��Ʒ��0Y��ǶP�%m~�gsl�ݴ�w.wmP�� �������ǈ���/47��S��0ǲ�d����+�1�q�O��.�+�k��z��;[��>���B�ݒc}{�1���c��Ej�u��C���9����ڎ�2�6m�;[��Z82�	��]k_
W����j�	�k٠.y&��3Z����:M�pfk� ;�8"�<�9U`e�VZ�B���
��(r]�-k"�zҟu�M(��|�56I7q�Z|F]>MiA��P�b:23�yb�I��$B�'�c�`��i+l5w��c��O�+B���ߘ{}"���Y#_V'i�q�|;�9�/c�*_�a�=<��2
n�A���3Y�}���E�^ʃ,ը�~�;��k�^���C���Y��� E�
Xby�sǩ��4U̚���������Mh�)�m�{��с\m�On1���d�G����3��l�B�T���m=����.������Bґ-W�LWF��WHZ�����	��6��;��ڷ�|鳧t<_v��"�9~�i1�6���%m��+lr
=*4׉���v��0����l$�4��s"��x3�&\)�c�T$e_F;�O�a-���ܧ�fx����o:�	�/N���m孇r�DI��u�h�ª�txt%�;%�|�v-�b;~�Rg��5��=i����u&�FH1�f�w��u�0�\����Rސ����o7����IA������\h흆[��"�ƀ��e���u.��PTwj��)߾k��U�E�J���������v�.���ް�����H6B������d��
?��*٭���{��!����L�s0�8�4������d(X��ݞ��y��	(�%���vo,�f�p�'������s�dF�����V�w�HO�y�}G��G��zKDkf�1Hyz�zNg�IudU`��ݻ:`o�D���\S��]�Ӯm����Гg���(;t��v]s�DF�S;r\3��w��CR��S��,#�=�|d�/5a�6!�L��[@�f�e`>�H�ar�fnV��6o'���1ts'swOfft�����i���n�}���d���b.��*P����{Zfb�E�^��.A��q$�n��v:C�	�2�*+���e�)ޝrtu��f���Ud��ב�o��H���i�^�:���m�oj�?j��D3D��k�k�)����@+I�,�89tnh[Mv�/-kX2e1�ur��e֕�R��RO9��D��
us �w"�T����S�T���_{:����^��Cũ%w��8�S���c�;z��f���j2T�W��E���_��y�7�¬a%+f��fp4tt�E�����m�7H)M�3蛣^��[��W�H��Fs]/��*~~�u�(�����2�2T�T���t=:`
�Z�����X�8e񮣍){nK$�qQS 堺St����P�:���D���w���vI�/X#i�o	�ˬ$��v���fU%�x�$a��g:���Nm�U�]��(�;��u���9],K�k���b��R�!���oY}��΋
����F����5.�䒴�wl�+���n0�y;p�ՙf0���7�S}z�� !چ��]|�c����W�t�qn������fJT���_������n�֪��*g+a��S��%3[�K�3U���) xc�<�gvwi�P�%������jޗ(ϧ�zV4�����V�݋���V&���o���I%��x��lu����Hs'f:L+�z[|�G�F�M8��N�\K�*��Ҷ ���^���s�"�	C1�*W��k����~I�^-�`�v�)A���]W���C�r9��v�G��TUy��^�2�[��u�M��ֱ͡ح\ř`������7f�c^d��L�iH��r������&gg��t��s��uq�����0K�n[U�ᦛ6	�󍮑S�OJ� ���{)����>cB|��i,��dX̫/�;���I�^�1��'/ #~�#�:ZA4-�_*H���]�qڮ�e��*7>����Yx�+2"o���n�nO��U>�V ���k���F	��~�,:��b{���n�����ZV"k�.������뇾��؈�l��k֑�4�45c4i���˜��T��M�ͦvo�k:�j�|����Kٽ�^�!<��jn���*%�;	�Ϟ�N-�l��];�'Rf;-R/v.P�q+/�R5jR�W�WuG1�E�e��u��1�M�8צ��ZC�d�yy�V�5��s��x�M���a��xVŌ=i���u
�er���ҽ��`�M?I�M);f]��R�r�l6ە[I�H�3���i⇵S��o6.�4�B�M�	$v-ȷ71�/���ޞ;BZ�<�	�D���M�Bm��ʢx�3w6�5�Gu�Sի�`D��F�f�y}���)˅<�t,���["����k�}R�^�\�>��E���-�������6�!�,L�-5X6��`z�mR���J�&��TG�t�;�{!�%�#"���Z�.DU���V���욭�HK�hY�n�2�V�l�# rU�>,��4r6k��tW�DV��>k���U�s���T��U��H�a�[�eZ+u���D����_g��ޚ�ѷ���I�U��on����%�Ő��Ia��1�Sw���Utx����Fl�(Ȭ���%�t�Z�mȨ�,*�N��=����4Z`�pؔ�o�\��O{��r�1�˪l��ں���Pt�������+���_�z1�e��+��WE5k�;�;
x�T9��m��Ͳ�v��|֟{�`��!�v���v�"��Z�E���`���Y�}Gz3�";���I�ݼ����b=ʓHF�e9��n�����$=F^̴�����L�օ���隆/ٵC�ߺ��嫬y������[d��4�T��N�ť-3����*�g-l��]�Ww�� Ə{��-Z�ڗק%��֪º�?	`&s�Y�n�����ⳁِ�U9:�9D�YնQ�W���U"f>�4I��ܐ31I/�B�b�h��e;-��ڇ*��ڔ.�vgg�y��#�W� } �M����ª/�D
1��Lٛ"�u��vŒ�/�HL�K�B�\�_Vs�=U'����Vޛ�p��N6��^652U, �ʡ���(����}-i_�a��}�-�ȶ�#s|��f��&����2z�,��7j�̉��D��k�KWӪ��"���˕�`rMu�t���{��EI�����]�����g�r�)��Mt^�V֚� U�-^�m�ˉמ�˱%Z���C����Ż*�1�b�:sJ���Nܣ�Y���Z}9��%^��n�"�Ii�ִo!��\5iv�qz���x��u��:��j�˭�����횻g�؆2&��(7ty��F�����y%�a��J��C���B�=HB�WW�;��w����K��r�Fλ�x��:,b�bhl
����d��G\��|��շyjj�mW�|B��MF0�."�.k3%7�cI�n��K��'9����CN�����8�7�+:�_v�ҡ�+s�T��ك2�r��-`�	�i֢�Ժ7	�;ٰ����
/�n�V.$M^�����y��E
0��ul����3�M�2;��0����Z���}s��O����a�uvv��﷮�8�����"xt�669�͙4�08J��TH���N���\{pb�}ۧ����,G�� �:�O=�wn`��dg>���������ɱ��-,��C��+�Y���Ln�7��3HV���W5H������Tq��7\��k�/o�*a�S�3�'��/�Q�:jj汩ڮ�Ev���B�m�����KY��THz���.$5s�Ji����kRӼ"�$��Vbq[������
�F�\.��n�����z�u�=w���o%�l�]�K��7��Vr��Jô�YÌq�H���*鬲�����Dh�9[�� ��Eq&�M�Eŭ������0(��B/��o��3��X���f`�b���2�Z<2�������B����L��9��=-_e����Qo�<�u�N����8��vs/���N�����p`�l����/2-�:nK:��6����ӱaw`bov�
�evr&&Z�ԋl=1�����,�uWJy��<WKrDߋ�ݿ�o��{&rLu�Cq�y�Ӝrb���J����u�#zo��l�fm��������wJ�4�콏��A�J��۳��-��b��8VǝoE>>RS�1��cc�e=E��5�^��ۚ�;#����t(��ώ3?�÷fȅ�>�(��,ȍ��Ҵ��o�	5^���2�Y�z�qm�g7F{}��tYR{�o�8wC�3��Փ���OZ�'�W�sl�3�M˰��i�ekƩΊz����a�|�5���[4�Ttx���݌=��\���8���E�ћ�B�eǟY�O# ��@J
�h��:�ǧ�9�UBW6��st\�w���W�g}<$H�zi��z ��}������IÝO^qO\�{��F�{��ђxX�4#e�-���OU��/���>�7����dQW�QE������**�U@]�|q�����A�°���2�0����0���L L�2,ʳ ��!���/�D#�  �D �UV @�|>�*���� �� �p 2�0 2(2 0�2(2�0(0a�yDEAT .Q �|� 0ʪ�"��.@UXeUa� !�U� �|�� !� !�U�QV@ �E�U�K�a�a�`XeXedY�fQ�;CȰ��ʰ������Ȱ�0,0,:� C�"��(� �(����`��>���x4�  L�*Q���z����}��3_�~��o��1�����f�o/�������	��1?_���}_y��W���������D_��� ���h��?"@���d�����d?� ��A��c�9 7��ޟA����	�����k�{�TYQTIUV�  � 
@ �   � & � 	�  � &@ � �UVI R ��   @X@UVX@P ��  H�$�.P�U�� %$U`d@�U�� &P�Ň����t�UEE�A�@(
R���w�����
���������[� x?���w���;�'�����@��ُ�����g�A ��������Ԋ *��W��~����UEw����!PW�������}p`�� ���?1�����x� *ߢ������ ����>�����C�y��ϧ��?��$������ �����R �����쇁I�����@�}'�`������>�z��I��� �
��T���~ɐ?�x�}A��_�����������>0`�ߞ�"����G������C�O��PVI��b�� ���` �����������Ĩ����I"UR��U%"�R��(TH)B�����$%P�$����@��$R*P%T�R
j#-����YS)-�Y*�mh�6� V!�e�5�mmdm�b�kժ�h�C�m���֤�kT�F�&�T��٫33aX�����+�	RM��Ic4mm�ٔ*T�&��j٬�P�J�mKa��JTZ+J&f(�Ȧ��[)�[mej�3���kU�cmYbV��R�Lқ� 8���d����R��4+iS�ӣn��K�9Ju��ڷv:���t�۩Cv�mNk��ls��J.v˅tSZu�ui�Қ�N\�ٵKj���V4�e�*��UZƴ�i�  �B�
(P�A�����
(P�н�� �(P�CCB��=
(U�{mG����Mʻ�]�9u;R�N�֒umn�(�mݭ�u��wn�m]�M��k���C�l%l�4͊.��6�0��  ]��U�t��6�[v�Tj��e����r�]vT�J�㩷[)]
��u'Fښ���ҪRS���� �B���aֵӨ��Δm�Q��ij�l1cl�*R�5f�� ���B�CH�o{�{v�S������4[t�긪�9���w�f�k����V[���ݪ���F���;��j��%����s�v�[6�f�CU���j�Lٚ��  ��hЯY�������ۅ�nʬ*'T;��k��T+j�ҭ�B��ĸtԫl���ڃ@v�:h��S�����]���fZ�f�[F^   �{Z-5޻9�R���lTt�]�l݌�[�:*2�Ԩ�
�mF��Já�6��j9u[����Zsr�P6��[Z���R�5Ro  ��A*�+��Q�uŶv5��:.�[��@UJj֤�l�목��n� Pt���� ۩� e�f�e�5�0kl�#[mk�  .�  
\s��� ���� `  ;8�  s��5�ݧ ��w  :.��@۹`��m�j`l�Q�V�a-�ʹx  ;� ��\ h �up K��  ���� �n @�� ��� P�m�p h� ���mV٬֚VU&�J�6��Z�  ׃�i@\�  7.�  ݜ4� 5��  �5���vn  ۳��(ـ  ˸� <���R�  E=�	)*Pa2 T����  E?��   �?&�R��L� �I6UH� ��ە�nd�����I(�U(!"e�%Z��
��yXE�f�VT�_g����Os9y�r@������BH�t��!$��@�� ��BC�P�#)�LX�RP���!�X�����¯A���I+��ND!ѤY����Ӂd.����k`�ck�4%�AWv��6�ff�)��Z��I��lZ��h�2]GhVd��U�h"� �ة��հ�/2�4.ٽa9��ך��
j;�(�Z�(o>
4I�iY*�J����k���z�۹�JwL��-Y�]�R��E=c6�t��	W��;)YCF�6aŮ0�&��qL�{4��ab�1�O����eg��{�v�u����3�s-QlJ|ܢb ��n�ʓ�m�ȯ�q�bii��ך*�ʊ��ҸC��ad �$��5Y��ћ�@`O1ИCtC'�[
�Ɗ:ԃǲӢ���p�r�Hi�m	�tJ��͕�޺��s1,ODV��ޭ�(�t��)��Mk^�Lݫ�7��K%I��;�w�-Z��:�k���HlX�0ܼj���W��Lڗ��.��X�TZnݓ6��cRf2+��!�L+
?��h���-���*V�5�o+q䶢��q�[zF�b�,��+tjM�}�Cu��Fi��[;(�1�ض��.�275�[1�"7Bm��n���n=��7@��Z�O5ݿ�1��/�Ӛd�A�!!�i]��wDn5��9G!�t���+v���6��Ȕɲ�L�j'��z��T���0)�[kKׇW�]�+f�ĵ��g`�1�	6PGuݷ���=*j���r]�s 57���}3e �<�۵�ѭ����V�&�P�bV'����ޠ����4�(�Z�(�%(A��I��3d��/U(F���b��/];b�QGa���G�Tt����t/\��s-6͵�H�ʬj͸q��4���ӓy�[�coi���]�	��mDOm�bVV)�WH��Ȱؗ��b�6���;49�!��Z�l-"�b�~��,�F�j8ȡ`�7RԶ,g)�4-V"�^���I�aW�!����s5��kĊ��Q]j�I!f��F�������i���$H��o�ibB�-V�ɒ����d=�Bd�#�DSU��ĥ���R��T�o�Y�.�:��h��_mP�q�*6�WMR[��lJ`��6�5L^���i6��N�r�Z��ئ����3 )���&�3KK6�af��.D/2ِ�g1�(����n��ds�T6��.��5I#��T¨4��(q�$z�ֶ�,:(�Z�%u��{cU-ڑ+Y�Y{y�.7r�DI�i�4�t&�A��.�ڶ[�%nC�L+�J�k���{mb�����Bzk*D��'L�c��T�@��Im�N�	��%Z[q�L�u�r�*#MTZ
�8�	[��(�����)�طt�U���j*�Cs �j+wZ���ڹq9/f��o,	�IY���0�6����-m�FZ u�����"���YD�%]Z�u����b���io��U�{�m"�8����w��f��@5� 1��l�e�F���k`74HJ��أH�|�c ��a�� fiBf�ĳ�͑��X�u��+D���J��6�ڎmZx�+̚���d�����M�Y��S$��v�`b�r= e`�%�m�-M5+q6��i��)���8V�E����7��S�ӧ/�(�^<x^�aB�n���1Qj��
1#4`�H�Mƪ�Bt�-e\V��N�!�6t��7�^�;��cT�q�:��@j�m����2��X̣�Ģc�L��l ^m���Z9�6�\�jm�tGZ���q���he��P%z��h,�P��Z6@m-��+	��� �Sv30�C��RMB��յW�"jf�
��l��(�$YX���kzH�lV�-7�j�����2]\�9�e�bɫ)�T֕Qֶ�;�Bc�C1�1��æ;�kJ�YJ��X{�Î���
Q��Kܰ(m"3�-��x�#E�i8�Jݽq�&�hZ��c�N��ueE�&pe�]�RQ�1�SCmd�6w���n�aT��++*;XrH�����Fp+�I
 �A��{�bX�l��n���v܊���v�U������z6Q�H�Ŋ�����Y�V�I.�����&���+����Md�)e�e�A�L5�EJ�w.��/i!�(�[��B���y�m U���Nd+N�[w�]Y��d4)�3�x�B�k!7��âz~Q@0F����wN<�NQ�w�%\D')l�be�Z�]&&0�������h�f�m�t�k0�<���"I��M��𧁁v3v6��p�Ʌ �cM��Y�ĕ1 e���� z�&H�dî������C5Xl�{a��n8@�ؑv��{Y�p�%��[�r���������h&/oE�7vۻ�եj��٭���%r�˒Sv6Էx�Aq��'
�u�����,��r���&Kvk+rP�A��i'��B�y1O#�oN���eM�� �Zk�bè��\�ì	��;'6E����I�d�tÀ���s�+�!R'c�Ѭ��,�̡{G��T�2�ۼ�q[�hP�y5/�R��@� C�	e�6��ئ %��Q�����f��֜��з�lr��	Q�,6�cb�0�^�g6�
��m��sN۷�St)�[I�����p�E�tNӫӱ��bkT�6��*�qn�i��V�Na̛b�,nT&�Jܥ��@�U��_Z��7Z��j�J�z�B��Մ�S�4����d�Yj�w��Ԣô��R�!� **����֧*	坬[�Gq@b�0��%	��0e��3g]k�GTJ�@��ee^�2�@�`1���B�r��u(�cp�oM�M�4h��rј���*9�9�ܕ��r�s^�O.�_�<�w��PQH8MMZj  p�� �P��-u���h"��
�jA�V(i�Ҙ�=63d'Y+T^�Sj�+[�B��ķz����R�1(Lb�2[孿��{���f��U� ٫�˫�G�ڽ�$��X���,��/m�
�9z�<,"�U
�EH'dl�_e�09q�#W�[V�gEv�t���
���&���=�P9�E,�-����i��-,�]����H;Ge�[� ,ށHe`W�yi����D5��m��q�@n �e;�4u��(�W���)�RqAZ�^*
'�%�w2����!9Zȹ���@;wd�.�*"jB��N�9A"��,Xg*]
zڙFW��+�q�*�N9J��wO5���Ri�xS�u�vm�^�{&�(��eh�H\X^�dφ�]KrFq"3�vn�����Sf&���� �m=n+����^\Xv�y��+F�r���+�)�
��q�9��<�	�d,�emc�*�t��ؤ����\F&&U1����s)�3`�<�H���إ��q8C�X�*8�x�LR�9@fX�.�mdWW��J��<Y�6ѣE�%9���5N�įj�:2��p�]��U���.�W6�F6���.�I��LX/n�b��Ÿ�Ey��6�ݫ	��rbw�Ef�0XB GdnC3��c;p�S.�)��L/���b�ƍ޷d_�͠�+�������;��+��ä�Վuz)�ԗ�mX�gʴ�zE�eI�Z�T�n�iX��f¾Ǝ���+M��3v����m�
$�X�P�n�&䕀�o�7v���Ź�Q��u։�����85�"eD��r�JM��2���%}�h�ܭ:�4�9Eƕ-�g7E��v*0f]C^�#��e�o.��w�U����)��a�4̗���#-JC��d��5�5�:�35�G7�X7�T�2���>b9wk��&T
��)�(Hjk7N��w{a+V�z�kV�������%r� 6�9H��,�+]���OTI^P	нФV�`M̥f+[��UnM��>��ebOe��%Qhՠe�a��|5���͍�`��i��:�UjZ�Y�*�o6d9#?;P`&��n6���R�(9�r�Q��񉸱�rh)G��"Ĵ`��Qvr ��#)k4��#w�`�9XmV4(^�q�� M�Te&v#�.� U+�����Mm�m�/+b��5�ZF���ޜ�4(Y܌'�Ѻ/B	�q�0�m��9[ڛ`6%*@�wb^�����l]C/e���F��Rɋ&��/B;t������m��)VwI�A�_����){�{��Bq=q�MarH� �j���Λ�e`!^L�n��!i�[���P���PEme�$���w���⎶5W	�-�2V1Fn���^�j�+iX�k�REv�U�IY�V̴讬t�5:_g9��m�ә���"��1�r\�j�CV�V#��T�<�#V���7B��lD-i�*�n�o3Fk[�NkY����0�T4ca[�v;u&V��E�I���+r�[/�j���F���`�͍�Dj�XeF��$#,�,hvh�Z�� �m�RV����������R���q<�W �q;]����V���G�6�L�r����!��u%!,@���M�j
�, ˷�rmn�kv=��ˊ۱��7-e-�0AoZ�և3r�m+���-F�,�!�
�ׄ���r� ���ukڇ9;���	-[���m��Ͷ���^YX��26C`��>rS�K~�ä7�ku��OL�Y�)i�pm|%]�2spV^S�w���1�RfDieC1� {V��7y1F�JkbU��Sٔ����Z]��{eX��	kpHZ�%S�*��Z֗�����v�1��e�(�	�e����nk	�$:�ON4YiU�}�T2�J�[Y;��K��/.�g�[� ��`�C)�R��1�ID-��j6��I���d�������8N�ƞڭ�n�3�e�/���$35f)+2i��5�`L��ۈ�yz(�or}+,͗R�Q�ӬQ�I�֭/1+�3l�HF�f�d���4�B�����U�N��Oj�ī����Ɔ��-	�������T�n�;�w)h�l�����t����>�?
��+���L�8\����Q��Ԣ�S����аoZ�e%J�X8v�ib�*ae� h ygY�H��� �@�V�����ZÍ�p��jr��}��dQot���4�nT�0�y8ca��y	i�YPV��u�A��lqU�q+���(�֯׻P�j��-���R����b��
�P�+f.X	�:���E2R
�v�!�n��o�u��D)k�{�f+��1��y],�� ��і��9#��'�)�2��u�u�f���i2 ��f�{�n�i�"��tm#���"��)n�Ad:c"(/.���g�p�p��A�U�O+/R� �7N,iJ[n����n���iÙQ�Ylұ.
�SxpUڇ��*�DWJ�j���
�Qr�Kɺs@F� �[�#+4�JKs+/`M�Yʸ����&�yRf�V2�Ak�Yֶ�ɉ,M�´Y�/qMJ���ym�Źj�t�w&��8/*%��j=�h�b Qksk4:�V��t�R���F�V!�ز���L6Y��i�Qn=b��{�*�t��ᥔ��:F�ׇ(��@�(I�C/mm)N�n�v�L�B��)�zb�Ь�Ւ1��z	�ӵ�b��B���r�<���%,��@�Z��e\�Qd�e-�
�.��J&ځ�ev�(V=9oU$�'��ǘ�^��=*-�E��U�Õu���UH�VYv�X ���M����42Vֽ�$*9FD�m3V�	�dܚ(1�j�M�(�##ȗ�M�f;ӟlɄy�,Ҭ�%`)�LdbR�+p�ux.)���R�r�c	0���X��J!�ĭ�ZS��a�p!�P���ԯT�vkӱ���j�M�n&��V�mf�m䶫��Z�2���{�:R�X��X7FU=J��!��c�$�m�41d����ZΆ��@�kj�i�W%F��Xy{� ��M<wR4&��;uC#v�̄�ٳ*1��źEZeՙyq'�E�&��KlJK-8�Z��R�� �srĸ�tPE㧣	���[- v�bH/������ҵ&S�tHy���%��A�m�'��K��]� �3hi�gN�z!�ܦ4 �qQ7�gTk6i�%�y�ɥ�+)�� Fئ5�9Z� ���%�{{J^*ԓk��Q忳	F�+��k6r���$���`�G5�ػ�3n�{�c�z���M�>ݙ���vݟ��j�ʗ��8TF'����ð��̩�j�DXfCr4"�u�C�pь�[��6��)I�2�V���w6X#&#�e�h��퇈*z��@��Um���P$���:˨j��+n�J����s06D�G�F�ŉS�-J�\�^R'��	��X�Zֈ.Qj�!;���m�q?�9w3�����HIMXI���iѩ����P��e��eGI�c�wE�WS��^�u���:�D
J�e^�l=V�Cd(���%V�wi�H�	�E%�+vK:���qhg+1f�;���,ݚ��kJ����`৺6�y��־��ګ�EPj]�[��X��/je�b��M8s!ǩ'��iU��)
iۅU��R�f�c�k��Y�p ���G/���]L��) ��{�`��h<�jm�Sa\YsC:�'t"����n�U����J�5aX�j�[l:�u海eed�沮�.d�dU�����r�����@�j��� :',7�(�q��ů�k؈cB�W�l���[o�x��F�	h��J�۠2+��V9b[�r�b���xRWR�$8��e�CM{���������|��-�]��aX);T��*����R3�0ۈ�E����ҩ�-��W��[����˗J��fD#yX�B�iv�!�,!��z�2GMO���)�S��nv��R��fsغ���cB�M�gu ����4���	�]��Gإ�vKZ���j�7�/������T�(㘙��eg>�k6�!pB�wUJU��b��]��L���z�m��!k��4$�)m@���M�hb�;���m��B���q����+���fr�`����&h���ZKh9�����A\�҆��/����|�B�y��M֘<^'U�k�u6�V=���z)b>tlMs���r8��mj�:����1W}��^	OKa4*饀
E�����g��Їuʷt+7rrA�R��:6q�#ޕ��;Z����=Ƨ�
�8J�;�d!�2�+�Y����-�c��-�fe��W3�kf	ӟJA\��l���HY����7�zA%s���mY5��5@��[�;�kA�Uc� x��vp/8�.�7O�bJ/()P���o2rD6��������.Z<���9t,����v�K��0������#�F�U�.��r׼�{D�g��;�vo]��7Q��6��ԡ��U��x�1󵫭� ��w
��46qӉ�T�Tל�vNV�����nԲ��oR�.ю
�U+�99�[���$1�֛Î�9C{jV�0��++V�@�f��:�`��K�ޒweu�+��J����6�	�b�PP�S"/��	6�v�yX��8��~���8�@(�q^��+�y�� ��%"D�׫v|*C����w�Ɔ�^��A��R�wNu�H��3��-�(���@��C�HQ���Cc�龹�u���RB������uӝG�'�MplHf�1�ͭp��ܱՊۥ2�����!樬-(H+��T�di�L�ٜ�|un�cqT{��ruö0z�f��:�A���a:������T;s:M����E���O�lҹ`WZО�2�y5��R���ж�#)Ql���]�0�ukz�K�I�8Q�.�r�4����[x
D_;X�y!������
�ƞ�ɯx*�j����H]��A����.L���I���F|�z� G�x��b��v09 �k��֕g���Dن8�ev�ަѿ��NIW	�����|�]\�I:��m�Q���<��V!�q���.����)�`�#i���L|9�ȳ��cz״�U�=�1���SM����I����x�ҥ��l�)���n⇖�vE{�o "���.l�Eh��dC�w��	SF�O���&_[f,RWW+��8yjt�K��Q>Ł�``O���M�x!��a}]�fG;W]�
��&�}�v�iv�`ႍ[����悯\�5��M���hu����"w�C����h[k�{W�"���G���rթF��[e)E[$]t��4^�у����2����C2�묉�ܬ�d���<��V��Х���RM��&�f.��7������ܵl�tW�qT������AQC�_ok��ƃ�������Ҷ���l��1����o�w1�v�D+eK{x��c��x�&J�l���,�{����{��`�wbs��'C�4=ո��P��&+�]�.��1��5\n�i���˓fH9ޝ���p��3Q��늱�jo;�X���_.K"��z���Mǽ{����۰Z��2�ml�Ik�|I����]�^��[%>�����] n�s�t� z��8��r�c����+0�C�/��&͹b�=x�ʘ<p�$�̳8搲�-]�\�k�˄�,d�P�ל���H�%7�(�;#���^�C9�{`��j�6�Λ��慪a�k�`��٬�C�iL4����s�e;���/�LOXzl����:T�^�[��SL7E�d�h���������1���ԖzQ]����Ax��m��%����#%V��N׹E9{�AG��Cb��y��{�ZWI�ذU���2m�*����33&��S+>L�rU���"��]��MɎ���i���n���3�;A����w��%�c�r�c%�cۇ�R�K�_#����!�q���j�=1	�:�˦ܾ�)0֜֝(�lx� )��陵��RZ�hЩ|tf̳Ǧ`-�j�5��',����LݻO����{�p8ܶ����,"�Ϯ�oV�;�=�O��1%4�X���;Ǘաn��MK�Z�=u��9 v	FR��%���&��xħ�h���c9�ވ�f���;��v';H�4s�ì�4�O2�JJܵ��m{���e��UpU��Hz	Y�f~����}����:(����u�k'+�%�L`��	�MKh��N�<�U�V��
%�u��tPE^�U�K�I��`;R�Th7)i(��u�mg�gb�U�We�.7],��\Z$cf剀�Y]�������$z�]�*�;�\�u��ˣǭŗ,�¹��rH�`����eat�tk�Ձ�$f�����n��=�Ն0>�_h\p�"/�L���.j��N�gM� ��V����<VR�m��P�9�t��t��`oy�
���t:[-8���5�뺱V��h�ۖ��إ!a3,ѭ�>��L�MyV�C>�R���cEW���%��@\u��a歾W�`�,'@�z�0/2S�w����L��%�s�7�KD�a發���R��k�3�$4��.�xS�[��޺����!E�����XT�Muji�R�����>�9�ӗ:�j�T�
���I�YP�R���p'.D��:g ��ur+�cwT���
g���&�E�k�����(����Y�m
Zm�*��lIaY���R��FZM4(u�d��ч��U����J|�J2���ʊ*S�mu���/^�KMI
��Q��e�4���g�-/(���\+���J����Zy3T�v�.��kn��~�H�	����K��s�Ƹ03��vn��%�43`aZ-�lؓqꤒ��ݴk<�c�]#�+N[��J���R�W�e��YH�A�+�%mC�u �Z͈s~��l��tޮ͋O������w�j��K��I��pE@�]Ii��&� 6�o�2к=�t>��W#���U�=�Vڵ-�a�\q�Q�ɴ;��\VFN]�9R���鈴Z;�'R��=G)���	y�.N��:�{{f�Pa�a�c�#�իH͂h�Jh��9بćEx4f�9�=��-]g���Z�&ַk�f���G�u#��S[fW)lec�Np�����U�'�9ͣ��e#�Ւ�y_K`�CKX�9��޸h�xD%���gl՚U*�+�$�g�\��ZŃuc\m��~�'/��bR2vZ���©���./�5�k��v`�r���D%K�W�=����E��Q�j���p�oRtej�SL������0,�a�dv��		9���8�a��<W��6>�b�
c��5:���*^S���:�=}�ҷ���OxH����.�v��H�L����n�y꠭vB��vA���?-���a�}y��F�}9\�X�;��!�=���")���\:��%�S�[�gHA�R$�Fly�Pӟm��BQ��be�$���a��l�Y�.^�t�֬���cΙVi8$�,�8,A�[�^�kk�6���jK���o�׍h1_��⦮K�9�Ҕ�<7J-��Ʊ�\~N�j�j��F����9oe喃�5��h����T�7��3�|]��5�6��</���	)�/2`P�Z�x����
W`�3+�(T�`��\�T��BmW��WsY6Y�mI|kh�A�� 7���V�Q'+�r��<*ٖ�2��3=���v=���莿Vm�hRb�pD�_!َ��N֙,b?h�6����a��RamCy���e(��}X��T8��OL���ok"�[>W��.�9�X;�j����
X[ʰ��3 ����8��CkDqk�>��c�v�pn��D>�RkuPͱtûҊ7!��<m5k[�v����8�7{u��=̭>.%��l�X��e�Z#�>A�VM��/镽�*o�x,�c��-�2�#��M�H�b��f�,�8�XsIw�kvu��y-�ȣ�ʷ���a�/�`ܬ�˧z񮡷Z�
�ُ�\�q��푗m��2���tU\U��3U��R�	W�н:�T�L���r}�7S���ܱ��[�gd����Eq��0ұ�>ph;;`�_f�P�g�7-q�-�{������R�뮈"	����u1'd�Q: ���*/x���b6c��	�Ŏ7���N�#���s;C��z�pE�.�WT��+3rqLk��U���ި�V���L��Лû�<%���]Mq ������V�>]���x�R�ʼk�J�Ǵ6}u
�AQH�һ�1�]f���s')�-v9ۮT���V;�[Kr_c4h	BZ��#��kzɕ\���I��r��3���*���Zov�Z]+;lKǹ���[*�������w6e%D��QH{�-�w^a@���R�)��2-)5���:Y\2��J�������:5����(3W���tp��-�hD�X�HK|.v1F��Q��]���{d�/aZD�l�;�dz���f�ͫ�f�#EomJ���e꽻J�N��އ;(��J/(�ם%Z9Q!/�>��9
��Gp�ݽ¡��C�j����[yK�����!�4�M#�>2�����ÑhH-��_<�c
9\N����X{i�Dr�t�6�к+�ku�K2@�"��Y$��;N�t��'ث1�J��v�>0� 7s��������wn]ە���yj̬���]x-�a֭PoƮF�@7F�6;:�����ՙ]0n34�`Ғ��Ƕ�uh����Z�.��;3(8�]Lf8��3u]@Ƚ�q�Ӆ7C^Exv�8T�V�7�8w`WH�5�7Ecwvi�K=]Q��}Y�tp��-�V;E@�p��g[���A4�F�^Lz��9E�/�}�w��>����6�>���݈��4��*�#˳[��J�*S�V�W7�W���s��r� �P�gkY����aM=k_L�^ǃ9���ꖩ�8�ՒRw@znڛd�uaJ��iJyҍ`怃�S>߻z=��>��qI�Vo<��XȔ�:���\�b��3����%4e�;�;z���.�!iE�W%�����N!���<���%��u��_4��f�64d�;mP8�o�C��9��wB�D�ޛ�[;�������m,�>u�j�� 1���{�'r�I\��fX�f��7�S�A���{%�NWPt��[eu[�^u�T�R�e</��f���D��I����ʰ)�f+Bҭu9��g(�xB�R��9��WO��8N6���s�����*�i�ۉ�u;.�l{��S��d+.(A�u�����i̭�ڒ�"��D�{w�۴�Ω�w}�ku���%�p����v�+)Jʝ��Y�6c�s"A_B��v�Q[W`eg)��A�B:,��uH5�e)�-�֎�|R<4���
d3�e��ۼE7�W0.[��E�y�7�����	f��w���:C��!m��K6���Q%1w2�����V�Hf_"�j4Ҧ���lإ}�#��I[��9_u�!غj"��XV��5Ld8-4\$���59-K��V��e���U�3���}���+ϱ�W�W^S�Җ8X�ə��4�hV"�uiѨV�h�T�5��fk��3���z��/#�e�8's����9͗Y:��r�$��q��B��}�6���+15cg+DL#{F�a�Փ����Ԇϝ<[�;�qۥ&V�i-���[b��Յ��	R� 8u�s5{��z�uQ�S�V��K���oQ��&w:�KD��b�+�|3:�⑦�֎n�V�𛕯��%b�C
4�H�]c�4�5���\hԋ�
:��m�5�;����oa�1$���ǵV>ۊmi�[϶���������=�pH�S�܍��V9&�T�T��\;r��\��E�T��r�O0�묹�`�1�e����V+=@�b}a�>@oV�$��Vu1j�͍�F�ܼŐ�-Y��{4�(0h��X���U��as��w����9*�M�e�$	���*��[����;w�$ܟ-R�]��^�jV�Ԑr̕�h3��Eu��$���umk�M��n!ep��~^ܠV^7�0�V���
ur���z��K�6�'w7�t�LZy`�s"פ{2�
j�9J
���PRB
�H��2\�k2RM_b���H7o��p��y���	!G��Uܫ�:�^D�P�K4i\cV�Tn�֞�5q�/�����&3`�x)OwTۊ���&˴٨#m\/fM_Ku�:�j}Z��ގ��rpB��WfC(��,�fty�Z8N�VV��D�ʔ��uk��j�gՆ͎]�S\��_Q6����ү��]).�ޔx��KyL��8d������a�Pob:�K>	q��[knb�&Ho,�N�W`FgZ�Ȃi��BԷ�lGn�+���ܭ����^����r�4j0�CI�B�%F���xð�X��zo���{,%Y��v&��U����}1���#�eԝ�CX�C9GJ��8aӊ���n�6-�\ڙ�.�*Bfޗ|x��Q��X�	���6�_[VX�}�oC̹_)���Sr�ku�R/��n&oS��l�=����L�����+Z��]����*sK�N��V���CO�2�&b=T8���a8bo���[{Ӎ��÷�P=i�ܺy��e����A*=��E��w�*F�wo9�:��4T�˭�	����%�F�E
���-,"�w5-�/w6�ϔݷPرَ�gE ��{M ��ܵ6F�����|v��]r�BgI,�nF)s�uq��3����׊��y���� �qVc�x�Te�;[&��Wc���ï5�Ͽ}��HBI	�BH�~���c��m�k�����\���H ����&���{�%k��X�nhk�z�r�	]1D�H����&�V0�}F,�,�˴�f�4,�h��]�<Y�#!�D���de8�IlZ�,��A������o����˦Za��UV�e�RA��dLS�;Hl�6�Kwt����ae��k�a��p�[V��f��q
}dN̾0|0Zv�����rr����2A�DJ6���������V��A�\��,+�i����[�r_��ۥn8'<噖�a��cj�|ru�|�q_3��zEY]Eh	�/)u)���U�ԛX掕Qh[I�f�qn���;)Aw�E=�o��`�v�Bӏ��mn;�b�@�I�Ӂ��7�Կ��V�#�mc��f�x5
j�ݛ�����]:;܁���3�y.��ȗ�e\'F�"k�u��w�8g-�y����\vEQ�x/x\�zh�cee�*#YNCn *�u��v��q��[*H6ݗCnRZZ�rG�,��a�Z�bfk�j��@�Ϲ�����)ε\C�*2rY�U��;Uz'V��s%j��Ā��RL�:�<�s����*1Gn�O�좠��;v�#�K�q�,fwrG�ˆNܓ&8��&��x��dgCcĠtp�9�&�I��]}�mjS�����'�4H�}�'<�Bo�� ��\sT�����+u�Cj�Q��*1�naڋ�x6�2n�iY�2���S���l�(�C5{������_G8t�w0�Ƶ�W��$Q|�(D�0��E{�)cś�p����iWrd�e��u�@7{��1��@���`�ӻ"��X�4�+�W2����9�g2��������f���)b.�Gt�H����3�A÷�����r�K���t��=R�0_ݙz���Q��v�]V،��>�k��81��2l�R�'�
�qU�]#��_�ga����V\��]��*f21����J��ev��������L=�Y�\�bT8j��-�q��˼�mtxt�8�]��v,e��J���,E���WѪ�x�a�bO�}w��tzM�
� T�MP ���UU��1h���d]*�$lr/�8zZլ�C^�5xOi-kW�������͠�wX��f_&\�d�e��3	�6��a�і\2_h\�j��s�zr��<��i̖�%�l������g"Y k�n���X+���:ى�ԗ
�ܷ�`s"}���"�\�����.%�a�۪է+	w��n7��;I<�m�nd��8�X�.�����T�4�]��F���os(*ԨM������+uh�GDJs�$(���\e�:�f,�(Auy%�C;}"WK�*U��0uM"�H����AS\�@3�S�^�:Qf����,����nkF���ꅭ��*3�	��uuIN�9&�{[ï��'tX�^wɻ9"�V�LОP��z|N7rfЏZ<������K&Yt;�|sF`�*�L�ˬ3�L|ӏz�gN�G��LM� �q�.�@�Y�-�ش�uTAv���N�i�<{�6�Z�nҁ����F7�d	ՙ��+^r=F�%���,�1P��^o�`�2YY���MJ�]"SD7Aea7��h�->�?f�e�j���I;�Ô��}���M�����A�n���Ye�
�l���o���v���c|y��'��A	�`�ي�<KW��XLI��)S�Źz��˫י�q��);�����f�J�.݇�'(}�%�0;u��]�_%�d{u��w#�'S8�5���@�Ksd�t%G ���Tܜ��Pi|R����ƴ]��^S:�NϺss[�qͮ�^ǚJ�ՇVn���ѡ]�}�:�]�m��1ȍ�b�{l�C;�H^!m��ח���jb�VQ[Q`���t=5����eu��- �x����.xv�'**�d�R��9����+&��Yy�1k���jb.�+ ͊���:ȆraN�Ƃ� �,����Q�x:��X��ƍ�<M(�ҳ�͋i�罢e�ӧ�xd/Kؘ
��Z��sM��@'��t�g������9�
�Q�
sT�5��	|���̾���t�ʖ�;���#�GғU�\�]rd̮�����7��ٛ���A*8g&S�u�n�����n���f��f�*Z���xG����i�d�-��8Z�N(���y\��g��N�Y�Z�����8�1�\��p>��2�fS;
0����,�ǣ�ɭ�J-�T�8XԘ��X�Y��m�1�v�w8��R�n�o��RL�s�_MH�`56��p��G^��c��Ӧ�]3�÷-��'=T�Q�\ɡ��dx����Ob�@�81\�Ã)�y���k1����.�`f��#�kyF1F���y����-!�W �NN��i��h�wr�I�&Ђ*a�ʳ�a����;��%�됵�2R�^��Eh�"D.��!$���]r�QJŉA���n@���G7h���hN8�
�5�/�k����w�g}��֝_����d��5ٍ��=�)��X����"��n��&>@b]��s�����u���	��S3Tn�n0�p{�񭶨jh�X�H%�4a��+�=VyE��F!�6>a���»٩��/k^7sp�d�ޣ��������ڠXA��H��1d��Z0M��ƮT��W0^m�������LQ7vSm-4c�����v�K^�U�
D�C3�b]mr��y�E5j����]k��gjV+�N9�c�UƸ�݌��N�����Zh(�-�(�c��57>O�
�we]�?�7��ki�r�./���R��Z��&���͝v*p\����)�n�FJ��|WXU5���m,�v5�\��Ʒ�b��:Z/��s��]���Me�1"�k��Y��"
�پٕ��$ǚՠ�U L?kɩ���;P�]��p�e�$:�8�レ���s	|w�zf�ݰ_G�q[ыE�Z9�H������X����AI��՛Z���A<8��2>v�J'ǯ6�@^�,ܓ�b۬o�<j�*y{���>� e@�Y��e&�N��K���!d_*�-���v�M�Z�%cΏZ53V(��1+ك�f�T��)��B��
X�����h-I̋<t���ك8�{�w�hQfd��crN�1H�yd����gI΄hyU�Ԏky�0�n�g{��u��"㥙V�r����2�!�F�]���gP���|������q9��ju{��c�$e�0�ٻ�;��Xy9�^�1a58��-
X�Dr��c�M���EC�Ԭ�r�y]	������t�D��������F��	Wv��ԏ
��ܑ�Yf��Vg|�]�2�:��&,�j�-��t�]ڰ�v*�):M�;��5���=]��vXk��gYV�B�v��il�˿���}Un����֊�M�w
ѷ��)��	Ϫ$�� `WPfb�*]�8��2�!WvI�*v�,:f�����VDenV$+�[�8ݛ��gU������ �P�b����\��d1;�AKT<��w�u�=$Ԓ��E.�#�*��.���K�wխ�@�@�fCE�F� !�``��w�H٭e��-1[d�'k�/L\d���JXzu�X�;!�� E����m<��z�4%�Cc��E!!v^1��;���;�����y1���l�L�ԭn�ڶx�]�j>
��<C���35A�ihB΂·ج�>v�i��.!wH�4�S���r��0x���Pk&r 9�C(AÆ^d|�;܇�(B�
nv�����8(�f���MŢgt}�t�zz��� �v��TY:;Y�P�xcneE�i�V7m�S�1u�:����5ų����E3:ޛ�(=���+�Qn)mT�I����ov*��\�(޾���R�V����f��>�qSF�q�'6��s0�ʊV�2A�Bff�wI,3f�S0�������kN|9커"��S��٩��Q��n��pg)J���k�����.���;��|� �t��<�&����N��8��9/��;Σ|�VqJ��'r& R�O�*�\���n�s���R���-��Fe�t�Vd����_'B�o�,ښw7q��˦�ue>������j��h��_V�
}׷�6����X:
הv�sUw�E �O��Y��1˙N�Q�����f5]�)�����hڻ��Sb�����Q�/����f⶯��w��,<)H��}u٭�3R��W)�u�[x{�J� �:�1U��P�\����u���/��e]��z�Q��������2f��$�iծ,���w��<6�=�e�h��J]<��N*ed�bv��C�k���:�V殡��C��L���j�|j�2��Q7ObkD���ud��ce�X�N���MOp$s+�z���6s���H@:�K5��%�,X.o=Ź��c�.�qlrTE�@�>GY��'�!mm�x[��:-9*fJF.q&��ɀ3�
�Z�76�U��(ٵ]ݧi�� 9K�H�r�p���;U�r�1�f�͌t/s��p-��J����ɆY���tX;fШ��k��<�{dˤ9���f8�H_Xan�2��z3$ G���Op�c-r�]�[�7ST��y���i����bS,�pmʽ����
��=	>�`��k��{[��4q2NN��1��j]�"ARq��P]�z"���B��YF1�>}���2���o��a���]�EeYޡj#�P�J��ا�	@��{��_fQg+tjh�76Y��AyY�J�o,rVr�m.�#K�L��-]-��Vk \��������֩��[���+IY.�H���f�!|�G1�e����)lc�R�hܲ����B�)���w�뫮�����0.��e"Ti�u0�5bdK]�����lv�aWJ��W/��� Ѩs��MVu�B}W%�YR����siwZ�98d�ڳm�5�t��9I�ɢ���QOu�_D�,a����`�=\j�k��V��ELH1�+{�%�� F���@�v�*yu��+jѲ������YB��5�T�&n6�]���P�N��{��t�y1S#j˒��+#�(h�W�^�d=j�88�oHs%	9%��yK0.�l(�WX��4�>׊�ML���,V���y-����xњOp���4>����T�CA��c�]y��gM`�Ά1*�L�ǷH����ƞ� ��G����`,"���V�����]n!@�-��j�K
�8��I͊��뫨dy%�b��d�hi	[]�7X�km�wN��/v��E��;Q�?�w� ��7q
u|���w`Ùh�ڛ�&��/����b�l�v�_b�
n���!+��,����i�]�N.8���[,��,=�{��,�/����R�q�&$U;�-�3@6��V���zZ7X��mD���2d�I��M��L��h�7z���W8oPp�7�.��'4"�:��V�h�����}��L�m��ۼV�P��0]�A��-�`��*�%���N�a��{�8P���1u�{�Ie�y�gs����L��B��>T���G�[CR�VTtk9+��'��d�t�7�ly�p�me<;yYXg#��b��.��K��P/^ҠU�ˆ�5��f`�̲7"v�%�`�Y̧���D�p:a�W����X��\&�Y;A@ް�Ƭ*2Ʈ�U�`���o{:
��m__|�<�1���.���']i\��tr���Mk��>k
�Zu3�;�	���>�v�Π	m��&����4��d�O��f�+�^LH\݋��w
��p^<��sC���+��&���=����#ݤ�u�]�]��e�0�;|�ۘ�׼�u����u������]2��{U�Lw��C90���S@�G
V;F-��)�����?iձSN��'س�2w��$V/�U�\��J����z�C2�ˈ�A��֫�����<���2��WFʙ{��:z�`�y��ǯ�ڳ���&�2���d:�h��-wp�t�ҕu�A��Y��ٯK�:��A�Ķ��F�o[�\,h�*_hx�N��3F��ͶҘ��;�R��e���V�giÂ7f�)��%p}]�N���;$A/S���*6%[�L:"�`��*w��O"a��ػ#�6�k��"0�B���t,�22+�%m+�M��C#����t���Q�2�G���շ�bky訬�SX�w������Y�.ɉB���2�/o^mt��X�B¾2�:��-.0&�ꀁ|ȓ\+������f�"��"ux�ՠr�*ֵ=�.Վ�l��%VZ������F�.��/\����Q�vx*�һ$�sU��ȍ.�GX��*�����Ѧ�u���TS�,�͡�V�F���p��x�{ϥw�u��q�-X1�B�XzL]8�-�0,�5�u����w��4nR�g>���������e�B�-ÕP˕�,)�.�(�I���r�cU9H�\�'�B�UM}��:1�Y ���fR�=Ѝ�ޚa����X�zƸk(ٹF� &�B��鱍ƪ?�b�z�X�Ln�
�p*�e�eQ�[����.Ծ�5qO�mٴ����86�}[-r��P� ��n��k2��9"K�Pӻr]jЇU�[L4��-"#X:[h�������vl�/xe�ލ]-�4Ub��G��9.�J��x��ipv�M3�1 .�͵C*�d�d�ǥ[k���LhW^��v3V��u��I�z	��\8�ѽ6�l��µ�;�;�.J��,�J\� �-�4�����V��/�}��� .��·�x���UOmn-�����ܦ�w&�E;��޽����2�Q*�w�[���ڊ%����:�[�7u'������V�WG����[0N̕�쮑b�7[]�N�8�ڶ�u:��r�&�i���p=j�)Ϲ����w�n��t`:�1uz�LG��m��cd-h�� f�
��܏`�:+)�I��ZV
��=*�u)`m�,v�.��C���-�����a�e��/!��AC����"�f��n�&�B�Q���r�K�Y{&�Bn���մ�ՙ�����ђ���p�\vƻ2�b�嵥jc��f&FV(�
�)|l����E�j�2;M�4T��	���l�w�2��4��%��e�*�n43��A6r���휇n3ښ��o�5���N��*��zC��2�r��(�o�yb��K\��V/�1x3A�x�o]�U70�߈��t�Yׄ��jj�w����jߙ��Χzʹ��k\��hG���-��DwX�a�n�:\r�n"��Ø�u��Y�؎�/dÉZ��Ѿ�9����e<������h`G*l�hI+�yl��fD�[���i�Z��#tw�
t�Ҵ�8W@��}jkW�]S����ч�[���t"�]+��R3Gby�H�Ϣ�2̾Ҋ�K;��{2Q.�^P�h����T���tƴp��%5h���G1��ӣO߶~���~|���r��1��@PQb�R���m���$�E%T+-�ʅ*��Y"�X.%B�Y�
��DV��1
¢�QKl�+ ��,�Qh�0lQUf!X�bLT��Z���eAjLI��
ֲ�1B�
�Z�YU�X
EXT�aRTU��Rc �r�� ��
�[aQe`�AdS�RDd�33,�5(�B��R,Q@��TZ�(�Ҷ�#PR*�r� �(,�ZQ@X���TU��1��dX)1e�mZ��T+J�`��b0�RV��*�d�T�-j-�P+-�.Z�X�*6�R)R��J��m
�J�V0�6���-PPX���]����ώ"X�!ج7��+'Yp�7h���B(�Qmp��;H��[>��.� ��T�	܉��Sm�:H'*�Y:���uW$���׍X�!ݿ�1�03�ą_�TD�Y�{�ԭ��C�զ�r+��@Qd�uy�ʾ�X�h�����SW��%/�	��3=�N��r����b��y��9/n����I���� ���PC�/+�����
]4)�����Fz��1�)��ϳ��1�ld4��NC�8x@G"$�00��]�sf/5��c\˜y����5
�N�'����;Q�8w��`{q�~�5�h��H�7�Q����՗JڬQ���P��p�b�!���z����Od�B��cfk����˱�w+��O���)^�ʊA���G,�Ȋ��M��-�ٿ��+�<���tɸ[;���@���z��y����f5|0z�p?�'L'�6����W�}_��e1B�r1��'o��u�F٭Т\�����f�c�\#��X���x�&	A�H	���+�&Q�.�&bݛw��*�E��$鹞�o���@��_��jE�C�!���^Q5Ɋ�$y���k7����ϳ<�meذ�-�<�d�����abŘ�h�WX)�z�<1��O\ ��U�>U��q[Y	y��՛��F=�r'�'s����:�񓎮	��k���r�=�������i�Y���X�T�K�k}�s9ս�.�W
��+c;�&+!����7R�����8G��r��5~��uЄl
R��;�&����7�^q�{'d��bLZ�J��sDP�祛�i��\ӝ�`n��{�ӳ�1;��j��s;�Ix$��o�ts#��	�9�8�b>�ȷ�uB���DÎ���n��N��P�)�^q�V�c"���S_�"��x��1�̩��B�g���2�2�<�-��6�@Q~�"�����L��(�C�_³���U��lU����a �S>lY�Xw�C���<�Z���M�M�I?ey5Br���_���@w�/f����=���yb۽��4[��U	S70����S��ЍԓMK%i�1�jj��'��F�J�P��Y%�}=Q�ï����l��M�!LTBj�1_s�}&��	�+�z�b�C����9�Enq��Qs�a\d��Q�t���Xc�L�Rp��7QBB��
�|L^��x�G{�}��9�����4���Ɍ����� W�iM�sq�S��ihӟz�
c����G��uer�� ]��_:J��}�� �Y�cD�[�c��21���e�Y�C�fvX8�+�F��p���3��xٮ2�}�.ge��H�|Q��}ՔQ�{Gk���nK�{�u��63V���H'�b��:�k��<c�o�S��p|%�S����<2��L���b6h�a�3�y+e�tR��_��鞶L�4�=��`������zy���g�>u���ۊ��ƇD���J�:GG�V{-,�Vv�8F���󑒣�Z��a�]_e�7l�I��E��P�+��e?P�㲦�ۊ�<Qθ6�u�skv�L�>��[K����e��l��D�p0����Q��'�Y��p��=X��A.6TV�Ǳxj_�\��M��T��
Z,3����ŧ/�oG �㓒��v���|�+9BxJ<�����T��w�yMʜ���k�׫¥�z����5��0�t�'R����li:����iBbW��2)cNtk�2g���B�,p���n{r�v��T����q8+�v�E��b��Q2m]b�Q�+܅�b�����.gy�<�Z_�.un��f0V�!gތ����x��p��[贔�^�UB�r�&6��g`A���a�����[��p'3p�b9��*/#��=�>y¼ѵ�k��TA�F�ek�2��C.*�r*��w��}���30�a�⋌�J�wi5�4�l]��.�Ϯ$$���+6���8�^s��59�2��uv�],N�T��Rw�B���%Y���/�E\;�a�#u)+�G��ޘ����%�1B0-N���Е6! ����G���n�/����Y{͵��Yc�fNp�Hikc�Ӳp!uu��㕊bRj�}�цm�Jo&��`��(ԏfg� L��h�����WJO}�)�a3�|�e�=��m�s�4c�V�޵J��ޓ�1wwkh�����e����wU�A�U�Sڐ��fMW��dL���
@Q���v�wNTsN�N'#�׵��:�|������
�_�L����K�הl}�B���5�OJyT1�"���xۥ�"��� �9��!�n�@��?a3=Yn�ؠ��5gF6q�yc�5S~�~Fi���ˊ��28|}��1�4��I;p�P�����w5�%|}uO$����q�]�;��u,7�z�W+:4�Q�Z�q��L���1bc���s~�Q:���ET-���Jj��,<.	<��^��(��o�qB��{e�?W�C־�l��\�Z�+ �(� �W�\;ǥ}�2�,η�rI������^�x��nM�����������բ1�ީy����z�
�W�����N2�vnT��ƭr�����*c�Z>���_�m�~P.�YQ#eu9&�Wt�p[1��<t�n;"���8��l�6%z/���w76W�_K��ruE.ZڕD�@�K�UG8��6r4�.9�C�޿��S (��N�y�ϔ� X���{O���N��O�K�X;8GB�S�D�Г��s�<ˈ��	�(B�R� .:�'���bs@-eK�݀M���"��oKÅ�!wi�p�_�NcQ�m�qS��1�˸�W*Lq8�n�b��B(A���[�����P�`[�B�gB���\wM �>֮B��ߑ���n��;gi��#QÙ���vh���b�'���2�lȥմn4��j���h�����i@Ε�$�.���ڜ�����9�P�j������cU�:��h�紘�5y�ø�.�]�-z^᎚~�n�wv�|�@l�D���㍂Je��`���:�~[s���Z�b�b���L�-��"��jtu���\s��F5GKyU��j̭4�Gi�ZI�v���)�b�����\�����W�MX�fv=�%N�`��9k:he�{gLs��c)ܭ��#���'T�UbU��C�x��X�J$y��	������X�d!��Qt�Y�öE����\�CE��w�:�Q]Q�����Y=鈘]�p�A^w.��s�XWOk�-�(�#kx�(=�-%�m����S�{"��|$��#�����4v���8���v��m�xI��9��#�\��>�O9�u�Ҽ����ݮ�����:�cjΧ�C. bȎ�G�NY1h�;�4c�����sݬ��hW��o���B�Sд\K��Q����#ٹc�Ȓ��6]�켒GV����N�SSu�\.�C�}�y�,g��ӷ�<4�7�)�����^��`�ݚw%x��q��zn!��㑯j81(Ŏ�Y �Q; C�� �ÓZV���ݢ�宒ܰ�<����8�ѱ��=��|mU���u��~���Uz2ju7�&ɶ���-�e�7a!�Z�)��#��祛��ϰu��Fn�����������-�ѹ��ӎ����u���/�kvh���	�����\p���q���"k���y+�&�m_K���2�dV��X�Q�@�`}L���bԤ[��מ􆴈�A�������d�����@��o��S�s�Ac����h%V;��ah���t�!��6��ai!_T'�Ys��8�(���Y�<�#�0��M�l��<�ח�n��y
೐T�L�Os�Zk�t��`�+���o�*�j��l�n���J��u4Q���;�+j/- r�$�שכ�ߺu�l��N�μs�������t[$i�N������������%�p�a�@�72���!�zCK��{����{�O��Sͳ«^R�q��(���	ՑhX�T*-)f�?=/�WZ3���"�XnLh�W�r���0��Vޝ�Knn�b�/�E�c�����[����ҊC{����f4Q��R�y�	i�vV7�qe%�����0�&��:�� ��0�D9��M� P��|�Psj�7Kv�f�򳑢C��_V�:u�k�^��+)^�!�ɞ���7���PI6P�L�����*@=]��^3
܀��#f��x�V�\Z�B��p�LU/ yr�� �D~���\)�j�7��v�����u�\A�����p�0���*�X�$Tn�ѽi���ra���A�_e��l�&W�c4�7����e7,Gq�S`��<���\r���N�}��O�0�8��V�py=QA\��ɩ|q|��F��\c)����,'h�g*!1��\Mm��[3�GZ�?��h:�(����D���,����K�	�1WjD�H�u���9+к.H�]!T���k��)Wxy��:>��C�	�![}pc�mx!Ʃ�p�m�v�^���ࢸ6KJ�αacH����ꘞ����U��Zj�oк�+{���N�T�.*�z(vJ�[k���M����ԦС���,��r�ޕ�'bM:���ZMeꮧL�C.�4�ύ���WcP�������vݻگ{Ȅo��S
2S	q1���jr�p�pQ���
�j�����T���M��@��E�������H] �����"�*_[m�N��t��VK��a��Tٸz��_�gJfํ��U�{-.7)D�q;�w>�brǏ�K���(�&�pv^�0�R��Gc���R����<j�{�QW[�<J��y�4�*���l;��i��|��1�S��X�ϸ�p���+�[8�Pjs�# w�]����}�zR��]0G��i�>K�p�^���a��O,G0�-�~ܬS9T�j1�n��kkf{���S���/� -Ğ1Q��f�(N�~�`rB��O.�d�^�הnR���F�cN�钏����x�5fU?*�d�t9Hׄu�A��V�?զ*kOd����唄�ˇJ�ʨ}uM�q`i���������41�*V��ΧV�Y�����	&qq���=q��Xn1�ޛΔ^��"�ͣ��9��5ӳ�]Z@�)%��)�q�t����'k������#��}��Lř���2^�|�"���`F��$0������Yn�v�����m���U����˧G��f�ލ+���v�(⭳8L]k�,ޙp\Ҳ��E�R�'�Cy�"�w�}��Zn��7B��񿲨q`����l���A7�5Mȣc�9��
�HQ߷b�{�]h�}6�'J��*E�B��*���<�,]VE�{w������뜽ޡ�/!�Ѳ]�}����~����ע��h��2V��*�1/(tR����{��Xg�V �f��O5\2�{�Q�ϣ]1�-��r�Et��_�`�o�xT��F����s"���>	s��8+䓸Y:l柘�8�̺B�dq��@f��ýl-W�;�X�׫_�Z��Z]R�6v��p��q���_[�!��rP�0R+:r�\]�v�Φ%=����u��z������_�U�4�5��9�F�q6"��8��&��u�&-�8��LL'WH�����%q��2����X(Ȏ�x z6*��o�sK���˚&��ِEDZ�C����m��f���Р�=kH��߹1c���^�ȕO�A�+2ߖf?f��R��R��(`��De�D@�v:+�-�<����m�h�=Qێ�x�?f&[��)g�*�v�ɜ�g��Juh���{�5��l�D��I�ͅ�5qWB�*��s��!��z�|P���g��h�KR��ru	�����S�y�͙W.l���@�V`vrqnm���]�����pd�&)��Ӽ�ށ�k0s��q�����ƺ��o,�����6z!�������H���J�2�h����<��ŵۼ ǝ$$\�Qq�U�����Ϲ��cTt�{w"ʜ7� �$.1��VO[���ړNiS�7���[]��<����,�������1����W��i�(+���p���KUj�x}��ޯ<kW/
C�:�4��MP�bk#${T'~�z��$������[�M�覧�ug�-N�����f��0�zϺ�o�Cb�yc9T� /�l����JȬ����Z��������o��z)�]&�^�FN�Omc:<��O�F3�r�"r8QS4 ���2r�A���jb�&���;s�aq�P�p�ѷU�<4��
g�u�gٷ�z<�9��)��M\�����IBy_���<��ۖ�EٌN���=y O&+h�����y��],�?Vg��!��x1��C���|�)l���Or�إ?01��c�N>��&U��G�c�[��R����7��k�Iu��_l"%[�-�����w>,�#�5��cƎ���|������u.s�X��0�
J�v��J�>ޒ�W'[��N �h�hf�ᆣZ�e��V�H쪱`}|���f$��r�]���1��˲Eڈ.w�xun|�a��r���lyQ���K�������B�bR���f�n��<�ia7B<�L�,М��3��WD�c��n�$�{qVv�"�J@�{Y+�JF�p��Uy�@52�7҉w[s���ñP�:�\�.P�r�\���WW��f��Cn��y� �Hnj�����/w5Ў�[��>�`�OVn�k��Gэyׯ3�sq��A����r_i=FZ���{�'(�EY��,v�_f�-�Vb�k��3��%�j�qe��y�T�M��<�7� ��	��3��/3���@�,��|�!V�X#�����R�4쇛V����t��h�T,{K(��V�u0ֱ�kŲV� �'fZb�F- �'F�K�U�
�ֱ��-U�dc�e�E:���d�,lx�
Zu�Wsfdy�IʳX�r�1PH�Y�E"�gJk:�ھ���e�r��d9�t��
�[�B���1�ob�LV�*�5{J��
�"�R��qE|�S3*W0,&�󃰹�%�;�����YU8��c3w�v�W��ٻ��n=)v�/��Nj ��Y�l�ؙ�P���a.��.�H8�o[껙O8Hͅc�����9+<��(%v�>晭g�Ua�&�+ڤ�5�;��y�8�̄��<��ݼRI˲:���!f7S:�_a�252�����N��7�T���ΓYn��y��"��y���c�o��˸)�Z3���v�n[�&����i��ө������-k�m�Ȯ�����}2��Q�+��6���okmX�:mb�"��8X��b�A���>a��H�;8����te�����v�t�ы�so�a�S�ћ�5E�N��i���୬��.��e����G��oaRL�!k`�6�Hb��y\/~�/{�c���p}r���_r��X.8�@��æ��{�7�ǅ�G�	�h�[��-U�2!�&�j�C�e.o]�W�{C���-4�A]od0��t艢/fؕM����9���1��em3M��P`X+��9��v�RX6�=r�H.4���[J�o�Ҽ�����"ﳳ$ˍ����R�Vö�+l7��8	���J�V��P�*+�L8��v�~p)��̻*�H�u�?e9�Zy�Â|M��;!�Իr��Kkk����of�gmvޅ�����N��*���
�HP�p��WL��Bt!r����;�s*L�9�Sۚ���'VN�]ou@j���<����]x&�������Ϻ {�IWs95��`�:��Yu��Sӏ����4��vd|x����MkxEq�곽�H޼T�aTȽ|�N��i�H�f���ȩ��g��߽�!����*ȵ����X�J�E&%H�jVT�ȌiAH�4�R�d2�
���XQ+
��m�������*	hCU��AdŴ���	e�5�ֲ�̸�qn5�$"V6�`�bƸ�#��F�`��+��Ȍ��m��!Q�\
Z��E�������-�ڲ��mUCb�����Z��[�jV,
���TcZe�����m����eTX[ab"�IZ��ʮR�J*,-�1�*報�lX[EbV)U��mKVԭ�j*¥1�kj2ҵ�)Z�+aP�B�DU�5����U(«*V�(�TL�&Z�Z��E�V�l������jR+ZQ�R�����QUE�im�*�ekEEb�6��`�(��)��aT��n\I����+D�QTR�%U@������=~��^��s�鏑�5/)r�ǖ$y>|Ck6�DK�D�-�8���j��x�
=�4�T�̮t����nw>�a�J�3��xK��aS�G����,�����3IS��DI׌Ě����q8�n�g�6��]̧��N!������T>aS�{���l>Cs��ϒT%M�o�:�ǉ�LC�'�]�w��^��-�ۓ�b!��"$D�	��E'�Vz�w�z���i��}���|H,�{l1*f*Oɹ�U���q1Ѻ0Ӷf�^!�6ì�1'��1�C��?'�{�ͤI���<�*+:/dz�}~��V�{�b#DA���6��=I�����O�T����OP���^�w����a�f�
�VO�Hc<��HJ��Q�dY1'����*���d����^�{uw���\���E�	�B$z�֠c>I��y?w'm�a�����V��s[����<t��d�4�YYǷ�&�b�Ӷb�����je�Ax�2g����hJ�=燻����cf���vk���C}#���������{����X|�?����i���<�dݦ$x�g9��I���A|�u�����sVL|`T:��g��L11���4γ�����N�o����ѹ��,�"0��"0G�M�������mY�J��6y�����&&��*��j�d4��W��O����R_;�M�ǯ���I��~f*Mϻ�����~k�*9�ׇA�:�aڮ��d��H��\`W[��S|�ĕ������ٯ�H*���ˤ=OPĂ���AgY1��u4��1��y�B��.��kOP*N�Sϻ?X�,K?|�P��^����jek���g�}�}�@�_̝?szm������1�V������l>5CHq��$����H,�O|a��4�U�C�Ğ!R}�xèb�!���� ��#�#2O�B��=����e��g��L}a�b��g_�1����Aj|ɛ~���=J�sZ����V>�!��O\VM̦$�񓩏�� i$�����SĂϙ�5�1��DK᥺/.S���T�����j�&:f?}`c���g���3�11��s"��1?!����<H*��*w����h~���b��Jɸ}|M!�+�zɞk	�4��.Z���bO���P�������O���M�+ߗ������dGs��x_]jU�D����Z?o]�4*��ٙ��o���cL�����58	{���s]�ݣ��%��	��znW6rP��eQ���I|fE�Lv���Ҥ;�]<�w r+��Dv�/uu��Fu���S�7˯[U����/.?D?"�>~t�\��:ɴ�i����C
O8控�:¸��͡�:��I�c�_9���|�CÝ���x�Y<��ɤ1>C���*>~I���sw�Ҹ�}��\�p�@ĕ�;5`z�P��N!�I��N0�׹���>C����O�e�2|�l�s!�d����y�a�&�5��I�M����'��9���ǚ���H����ﾲ)�:�CV�z��c>M&�f�:���Sz���&=a�bx{@�8���p��$����h�:�<K��c'Z�Y+6{܊N2|�G��&�C�y^[�q���7�G�"��ޅ���=���m%}�d��4�Y���N;f$�PĂ$��1R�����g�11RV|Ρ������ �����4u�x�^�~���~�DY��I��kj������@!�{�b�C�+�~a��a�J�C�K���d6��Vy��ԛ�aC���8��Jϙ*T8�W�Xu$5i��c�Wx�3�>La�z�����X��&g�{�����q��������N���������N3�8�C?�XT~x�<=�SI=B����'�4�eNv�I�'���y�'����J�?ya�Y���G�25��y���}��מ�L���|
�����c��~���q��S���͡r������s���R|�O'{�i���!�����x��Y6y��m�tÎ�b�XC�%�g�Z<�$���o�9U�5���#�@��O��I���iN���V���2x�?O�$Rq
��|�O0+>I�]<d�i����kG�K�N�f��T�����G{�O�o��7�5�xg��e��4� Q��:j���Ρ��<�����g)1H>�8��6��J͞{��m����~-��q
��s(ꐩ8�}�0�&��`c;��4�ïΒs��ρ�7Ҫw��39#ވ#�|D���7�&!R��&&�|¸�ڤ�C����W��Ag�����H)��ì��Hc�a�T����x�ԩ?!|��<k&�tD�v^���L���Q���-�Q��-1������0v���l��b�_�'ɫߣa�3���hm֤���Oh_zLܮ�~(��w� }W{i�u��v��$�Kti܃.쉭̟DR�k�
ފ�݉x�݅�M<��M
]8�^캛���x�~�`Y�#
��&s^��IP:��g�&�ed�k�࡬�|�V2�$�����e��������=M$q񇮒w�d��������/���[�x�����:^���{�t���1:��Xx�Ĭ=�4�3�Ԙ��'���g�G{���$����P����<���|�x�f���B�̞���B�g����X'뫬����o4��^��:'o�O<���ϙ/�OΙ�������kϰ��x�^����v����0����i��Cr��A�$C|ﺆ�Hz� |���*$��R��J��g��s}j���ݻ���{ﾑX�"!��1d��3s˦q�������&Z�]!���M3��*>�kG���U@��sI=N�0��q��!�La߼��m �h~��!��H?y��т�5^U����|Y���"���t���8�@�T�N�M&�Y1'����+�
ͅ�'��}�>��m%@��~�m�%E���<�C�o�O���y�I=B��/�l�bÛt�_���5��p��A~a������&$��%q'�P�Ն+'�R~q��y@�g����%g��L4�<I�P��v��
��_Լ���_==�͝d��q��w�z�}��>{�{B3�� }|G����i>B�̞�ͫI��;�����Lk&}M2|j�g/)8�1�AV'����6�^!�1�|�C���6�Y�u秈��p]�:�u]o<�BD1@
t�a�:��bOy���8��!����:��+�7<I�*�k�M�I��`i�����\C�J����I�
�2T���4�:�$���έ
�:�s.�}��}�i~ü�f�`T4�]���6�Y��Zu�C��1�u�
��*����k
�ϻ�ܞ u*Of~��c�&$�yi���^ V��²�~����/�we�h���瞈b8�*J�&?�*,�:O.�q�0�|��I1��Y>e0*g9N�I��bA����N;I�����`
�z�����H/</|Ѵ:��$DCS�>��Є�������u���_�EíӖZڽ�F*@�m���t�0Y?�JlG^�)7��>�7��¡�Sba齤������Tyw�fct�`�S���<�uφb����6�M�A���Z�ltJ�Q;��u7�}�rSv�2/H��?�}�,��t��1C
����}I�1s)���L���1��'H�u�����&�u
�a��~���Rm�gr�2u1�����M?2g,P�3k��X���<c��h���u�N���?{�<>�:�Yzo������ZE�?'�c?'�V)��ϙ��)���$F��
�C�1���C���?f�8���ͼN2bN!_f���7�������ڻ~��Y��#�>��b>����G�����<�1���3Z��2UC̰ĜO�~Lf5�P��?d:ʚH,��0>f���Cy��'YP���ϳ��*�����9ޞ'
;{����Qڜ�#������N!�z��~��0�*�2l9t��T��go}ܕ<CT<P�i�J�*�b��_��&̺V��_���=I��*>!�I?&�G�[N2r�h��#�{~�G�#�#��w��+'���r(i �����u<f'�1��d����Ly���<CĂ����&!�;��1�>��e�R�����v�Rq
�'���0T�O�&�W�?����� ��xG |�T�����ɚ�������/l6s���=H*���a�%z�H>��C�ώ��C�� �L��06���b�*�XT���������^l�����FʦV{�",C�3�M u*O&P_S�>��zЊ�����w��κ�ds���X�f��ﱋ�:�|�gM{8/a�#0��8`�5�@�gB��$?��B��ɥa��ͥ��5�2F쫿�����9H�Ϻ��R�s�y�2��\zU���;+S��K��~��+э��Xb��ϛ�_5u�C��}w'�D�Y�+�tz������Ƃ��HJM(
�^c�.�yS_%a'Kp���'Bn�s�س��n{�v�+3�R��5�\���\:�w�Y��lp����pc�k��vA��6��Ը扴�R)I��i�z�E�^�](B%�4��T�����}�0uь�ے��N�-�n��L�󪢳{lz�wx��r�'�c.�o��0�e���F�����e=�6 �8�@R��ݙX��:ye==�
�H�0�{0���ua�aYl�{����1y��#ג����b֧;UH9[�u����_�K@UM^�kBK*�;����F��J�2�Ҥ�"rp���u��z�rܕ�p��OQ���ҪF|L!��enΈP�֊4~4�Y ~iJag���܏���]�xf_�i��*���"t3���T���~&��y��B�9�n<�>]�ss�KS�Yť����,J6):sp�>C(�e��ر)��e�'�t�ʺ��sE.[��hp�p�4]��ހ"���zI(h�0Pu_�c����ck)��,�:����������\�.J��9��Ky0x�IWi��v���8"�#+xef{���H����S����+%Nnb�g�ʓP}�*I��v�S�ﰾ��Ɍ���׆4�n�uc΢��]U��zo8O��G�:�s�E6�(X�3;��;x�����L�˩�P���{���
rKc�k�N=�x�P;&R7	�s3�[���Œ�-45:��v`}�nR�ic:��Wʒ����G>ݑ�W'f�f>M�Kw�a�(3m���:��֎NF�q���X�9-�ǀ�}�/r���1���D� ��;#�9)c���5�j���y`)�pG7��B �]%��[�+��E���Y��N���;؟��=S�حbb���~�+�!�<�?��p���шk&]���}z #\Q7	�!��j��b���(�<��1(o��eC��lu�3{�˞OS��R��F�|T��l�[4�$~G�{U�P���z`AY��V-B���Z�*9�%e�H��k
���0uHF:��.v��t�\b���o�U{m�<���������R�`�Yr��ϖ(F�QW�W�WO#��K�TF*l�qKG0�/��|qY��7�U���j�~��������՟7	��x�o ��p�R�a��0<�lu;ˬ}�&�WL��åq�y|a%�C7�F:i�b���R>KyL�����,U�u���aM2_����u+�mpgn���t	����I���@@#.~��G�q$�-|��K��-����4�W��?QN��d�V8�n�ѿ��`$ɕ�PP�O��n��њ�9�z���7�b�OK�i��(�r-+�]�7���"V��르^�����°ENz�Ī[����fKE�չӢ��>�ZHBv��ý32�f��yp.��s���e��J�Kw���m�@[)�_B�w]������e�l�)���=����͖�CĮ*��l�sP�s
�tDҪRRJ���Vծ�q��\�__�(dv��f��=�8B��$�s*��9̸�1�r�Ȅ��^����˃/i��3�{��ˋ��}��_/�����$E�IղU�ԞUL�-���'v����\i��6&,}������L-������^Y]���+l�'~�ow�sZ*���I�9��B��g��'�X �����s��������6�3d
���klE᪌�q�w�2Y�>�U�{�J����ԗ��uN�h��U�
�؞��'��4-��i�����q���P���֢���#P6b����j̭>&�{]�����A���K�|�g	�LV?�/f_!�W����U�W��\�|��j�RޞPy��軴V�{�I�4����xGq�+���r��y(����e��6?K�O�Kx-yO\�J�ySR���O�Yp�|=6�C,�}HY�T'������ߞG�C����&�WxVƫ���d��T�V�=�L�}�鄬��d�J��h�3�K4�^��O�����V�y�u}�9��4��������.D@�[L���:�}:��/wk3t��3H�������v��Tj[9�^��垤��ig��'!y����sCwqUjjo6ϚU5Ӡ3���*�\;H==����k�s �Ȭ�ٝ���[D��܁U��;���pگ�0��:�g??��y�+rk*��$8�.j���'���{e�*8Ceqhă�R}p�M��������[�fQH!�u�=�=ʖY{YΩx뭓���}�&�<�8xԯ9�-���
}0Ә�ۙ����=�MS��>F!$�/��+>쭛��@O���Z�a(z��f5��6v6���.^�u\�ب��L��6����h�C��&3裡Έ\c.#����%1���2��K��/۸�ת�W���c��FZ�!�-)�lU50/ƅ9�8+��Z��E��ASh^ztܨ+���i�[,�7� �o�_ZtD��j��]�G���;���W����d�sȺ8�`�Q0�#Ry8s�ʀl�V�η%}�^<��/
�b;�՛�I:�8ݛ�tߙ��L�ӻ���aF5t��Pع�1@3s��胤�2⸽I���m�Kw)c)������l֨R�Q�f։`;�t����YM���&{p�K6��}��d��� �ܮ�:����&rYmB��@���7�b�q(f�fI��<�;��ҵ�b���r
��������t��Csg�
>�ъ��Ѱر΢��;��S�^�߮�.�mBp���-̬[O�F���J�ҷBm9�"w=�[ޱ�������j�Z̔H������׾�l����iC�kN���V��H�xk��b=g�7�
Z�uS�!���A�	�S���mʝ���Q7�9�{�h��G����t�K��Q�uW�}/�Ny�{Y\�^d�wdE���Q�N����阷��/�1���ۧ�C��ǳF�<4����d��(Fa>r{�'��,z��o�� �'����C�6۠�G���b�j��5�&�D�%�h�fHr�xU�"1U�����q�E�R���c��� 8G��r���vj6TDI���睉�g��t������ï�4�<���Sd�D?,8gNz�o:7�]+��՛:��j<΢��-�1��0~�RP,7�y�X�����y��'-J�kzM�Ə��g��sț:��/���0|��$X��aM~���k�>��"n�nO��8t,�����4����ZXن���t��q/��]�RU����A�y�d�m#]�U��M��]3�������Σ�(fj]a�QIG&�5Q�Ka+�E=��� �'E���ɡ����I�g�+3����o˞vＱv��'����Eg�0��A��@Qn�,���WU�P�E���,����m�鴗j7s��|��r|��},w��"�⬠:�ol���i�.y�
|b�c9���owԏ0�b��Vyn|z��2���������8�ҞR�<�����W:���%�K%��1�j&�^T`VX�0��7
zh�T�vx�gJ;/p��0���0<� �����|�;%qۈ���\�Xa��p�� FEE�� ��ۻ������O ���H"~禾��'M��+�?c��
�ߴ�Whe�2��Y����(�.Wf�@�'�c��pt׌�@XlF�:'��p��������a���g0�{9:}��<�R�3�lӞ> �G�k�?Kڿq�Zk�i��-ĩ]�k���j�cџ#��}QsX^�0qH������0_�<�ӂ�i��_�1�D`�a�oQ�u��L����PW�_�T%7�C^/�'3�<�z�������T��D���7G�.�'uEIvވڵ��m\��3��κWӘdR��.��8!Nz�q�(���s��G�\��F��ɭ��ƱI���l�u�2����rN<�����;ξΓ9C���ե�H���<�mv�,���1 ��-��.%��'��biA\8�u8CZ[�9�ˊE��	�kA�]3����(�1d�P��ռ,�RZ�x���y���3X�L���A�t-�j�2����������Բvp�n��V�ÁP���ܾĻ�F!:m��}X�
�&�u&%T�sn]h���w"S��wܶAYê�l�K�}��2²s�KNF�I5�'`�����������ʚ�g�,�n�e8ݝ�������� ���s� or;J�Fl�WA���LFC/Ecg^�;�.vȚ��^��e��0D�6	���4��vZ}K3.G�fn�a��wG2�ֳ���4̺�Z�p���7��N��ټ �=]$=ִ��Ԣ{�Q���#=];����Ȃ��y�큣G�+����1ڈ�h�e^쥳��m�u�3kd�Z 4��ly��PJ��FU�[/���b�= el�:_�BD񦅱��ļ[z^�T8��.��j�v�N6�P��'ە2VV^b�!4�5\�v�%7���3���I�v�=�q���r�f�I�^�G7Iۗ��Z���]�z�b�}e�C�X�*L��k���:�g[�v]�EF�a�L��Au�o(>5�^L�����9��4�=�����M7�p��4a=K�ک���2���.�!*cɘ�fU������.��8f���K��A6o�^²R��;�-���2@��жԸf��
,�Z��v�f��W{.�]��yJg ��]
U�N���*�R_pj^�{�����i�x*]�~�wYԹP�̀�m�3m�<�9�W�,�+/�]�X��I+�gPf�Gx���8�ۥ�q�J]'��+��h;�ˢp�Ã�apC9v��D��f�:�c���( �@�<�V�}Y�E�rVC��N��1p7�C�ع�uE!������l�x�Ոe��du�ON��(Nn�c)��eY�u�ҝ0�;z�Gpthx�/n��<uP5(��\ʈU̖�����͂�WJ8�U��6��[�wW�-�%Hf��U��
��Nvp�
ΪA;�ƕ�wHBZ�Y9D�{]!�6�e��\��It�;�L��)��J��U�5;�V��X�`K>dqK4���Nx
u̜TߊWKD|>7�P�Q;�m�Z���N��3]Ϡ�,oX��SP��Ndx�j#6�+y!���j�����݈�2\�����w0C��hL�;�j�HhU4V^��'6'�[��rНS�\�0i�I�k��n7Ηa�,u��PĔ�h�7�%�,�0uԲ��WS2!+��"�-F�k���մ��[Yq�ʜt�}�D*��:���0�kim�#&��C�^t����̵�cG:Zm{n�����+f�PY�?\ȪT���D-�h�Tm���V�fSmX�jZX�U(�dUXZX5���l����J�4q�+R�YYP��[[Tl�r�ŵeB�J���"ԩjV��1�b�ʕ-�Tbĭ��QR�kA��j
1�R��k[X��cmE�"����m�j)U���Z�D�"T�hR�P�aU�XTQV�֢(�-EX�mYEX�+�p�RekJ�ƴ����E�*�Kmj1
��b������(��QeTb֖�,-��j(���R²��(��U`�+E�����-�(ZU�QTS),F1F%���VQ�h,1�TX��Ң��(+���k�*�+h����QR��QҔV���J�VҬ��U������m[[��߲ɂAu@˨��SK�A����w�t�:b�r��ge�kF���q芴+����N_Y仰铆 ��  �d�)�w{�_����Ƽ��!ƾ#ܺ�p�����BD��lO`Q�*b圠��N���ON�)Wx04�ϼ�q�ޞ9�Vz�ܣ4��1_HR�'2�
�9ו*�XnD���|���˗\vD��q,v�ECwP�uQ�qFJii1���T��ԒL�K��aF�qn�/�#�9��O��I܋~��GyXX�ߟ:/�lQ���*�$���Z�zX-�^𧖽O+/>;��ﶓ7�=n��:S7�h�ȳ���t���
�o�5yL�w��"!���G��8mz���B���6W��*��X�J��Ǖ4�yq��]�/8tg���V���S�|N��=k^HPs���J����ܠȳl]��/�c�w5)���gt������:���/��/A�{NJQ�l��a����]�!�\P���q����hp��ld&����/s��� -Ğ1D��fM��Wc�k,v�>]t��)W\՗ƈ3��K2�ϓ�,��LFۻ��#�8x��,,$����NnfWLO܃���i�/y���7���.�)>��;�����^���v����Q�p⃮�Ȝ�:)gx�ɹJ�{@��o�BIr�C��]y>s�
�t�"m�H�8���L9���U1>����Ҡ���a�.���v#��R���+~���}G�kn�x&y>����ó�����s�F��;���^�����?b���zڲy�-V�{��,�^���X�kE1by[�v�ݕf_!�R�p�P�S5�M���c����]e�ξ̬����,Ĺ9����X�U��ZU���3����(0�Vj���5�wx�Jt��n�+�f�����Ѩ�H��ʡ<�ǚ���_Em��w[�.�LJ�/�;�����\r!���cmU���<7����<;�_T�g�v2�����+�èC,�J�9%5?\F�xn1�#??�g[]i������3��r�3�g�y�Vs>`z=�"��x��1@�I���E�g#O�n�e�sN�Ϻr�*z�_P��fE��X����D�_�m����]C�ͤy�㦘�<lµ<���ָ�!s=�v��Օtn���/�ι��]�ذ)C�O=���o��Jg��7+�I&^<�eO.�5�ЈTT�ށqۘ��`[�t���!�ʡ���=���2n��*�5 �T�P�%����u�����:745C,�.R�F��Fą]����]f�K.��XHwk�[cV�����w	H�ll�\7tf:�rX�PSh���
�:�R�)��ѢѰo�Ds�W/�M�8:yJE����>���䨳Y����ED�V��*g��/��:-W��-)�o�TL��ƅ9΋�c5ą����sX����B'�ŷ�l�9tu�0�آ7����
�ţ>�r��=���(&Y\�t�wnv#&Ԥ��9.w0��H����c�2g)X���J�uD���=h
)�.p�Q^�5��<��k�Ϯs��cL�^�e�y��h���Q�m��=��G�۾R;�`ə��x�}iҜ�*����,���UTN�[�c"9�\p��/�Z(1o���x7Zغu\Ц�l�@��1�ڷ\ �𰬺�@W���-EX�N��js^�n$�p��#�JM�On|����N��	�[�Pخu<�=���pu���.9���~�ۃ��&���s��O�>�_T]�ㄡggb�x�f�Τ���s��`�V\F1y��4c�1�����2����1<�˅i~��\���KXS�
݉�.�Fq��½f��w���À²�H�;��\kLgE��LFL�� ��z���И}{t4kg͉L᜕��`T���+�[������mJ΋�Ic��0p�����e�+��݉�r�^wh�9{ÏQ�[�F�u,p�{̼���>��U�̇��
�j��5cd���v��XN��Ѣ��ۧl~��}���s�OLx���~�!x�� +Z^SY�FΎ�u�z�z|�>47��s�j�+��-Щ{6�i]n*E��D#<<*4�R�ްߚa!%g�+:sDK�ig!�豟b�Q[��>U��j%�܂�?7o!�=����%��m�A��$8��J�X�u�Muܹ�m;���}p��Kt�ϡ�@��,��u� Wͳp�b��$f�m�z���6��H�u4��V�L⹮ .9�'�i\K���AyZg�ހ"���Z�<4|<HU䏄�gf����:g�E���JÐ9��$�|�U/�γRnHP�� ������a3����:��8��[����v�1N3�:PФ�J���������kI;�)�5z�W��$�Q+}Hq�T'`�0�u㴘��4�����]�.L ����nk�[rva��K)���bsE�k�X�9j���.����g�Pm���zô�+B�QG�w���tp���9�6[��!�o���g��%R]�%,u�g��%�7.����(�s�c��GB.y���j
��]�Z���	2a#n��<��,MӗjcD�8���n��f5ٔ:!��f�WvLD���O~�B��k���.w;L�쟘�l�J��}{���9N�'q��N�d���/r�#7�QlvD�~� >�?3�ߤ��A��SVՋY4(/w*Ѧv�8{L��q�a�+h��Z�p�)ė��o�KW�A8�ێ��J���c5��p7y�����{~w=�����?A�56Ҩ���weǄ.'L{�|5������0uHF9��"��YL�,b;ٻd�1z�z��/u�o�;r�6"�n����o�UxpuQ+�+��z:ָ�����9���i�E��E����j:�yI]1��~��`C��UH�i�Z5�ܕ�kԍ�ī����L��Z�\���uE$c>e�T��8U�ClJ1�	�`W���/{S��[i9s'P��{��4����[ۇ�:�/K����M�C�M�Eg��������U�=�L������8�W)���
4/�~��w���q�8.T؂y�Ff�ng���HVqΐز]:�tuE�H�1��7q�֙\�ƌȈYdF�S��W�􊮝��z\�ݢ}��z�/��
;��%NP��k�؅��p�y�~�HC^Q�W�.�=�/]d���,[(����O��ne�.���%����o���,��d�T��f�-��_%��|'$[ִ�=�`��q��	R�v�u�
U�����R���ft�p�́��f������c+�lMW	��+҂r����������zZO�=<7�}�!SWpVtx��)5?nD^&�ϵ�����lok<���;��N�E���W&�)͉�f������2����:�o0��"6�=o����h�����U�0J�ALXRa
MP��S�a�`�:c�Cr���v2��cx��3ڥ��8ƈT�'�웹㾪�#z��R6%��a��a�a���w��r���{aI�.�-Vó��X}3y�}.��75��S#��m����7���&�M�v#�{p5ˎ�&��-�~>��k��^+#;��	��%��dy��[;���Tu�TuX��-NW����#���m-A��NbR�{�P����:DF+��,pWwq�OI�T=}2ެ� b��0�w86Ἶ�QFقR7&,V4��_�Y�����k4�_��T��5��w���M���9�a��ylvD7'֌��1����>O�[yr��z�Y[T��tu�+�2BE�C۸L䦯����q�y�r�U�hd)�"6ԁ=�3�j\���:��{�d;GGq��>{�������8+��;�M���y{B�Q���"�s�G&�r�Ҽ�W� �+5I��F��p�t_�s��pB'�;�Q,���[�c�1��gt}��r�D�\{�����\<E����x���� Ϯ��^焼�ơ4c�;]�,J�O�=�=	a��f�9���1p������[U�Vv�xJ�9j�H��w�9l���Ab�D.m#�J㦘��";�4�����ǽ}t:�jT~��2P���[�C�"a��+�a.��Y��̍�<��kf�n�DhLcz6soKs�Xx�n��jVr{�dԤ;
E�B�z�GC�d�1��� f6\�g�SY�c$��SB: ;(�n�x�%�x�!���TL��Ƅ����Q������{��xq^�p�h��5B`�7�l��]e#�3�dZrD	x�.Uq��N��<7g�}�|$h��z���H��3g�kD�d�uU�B6	 .�,vNK�s�����&�U�4�Y���y���T:���>��߳� b/�5��A���:�^�o8�%zsuOp[��]]�7��8���Q�ad1��U:�	����<t>>��[�3���J�^��po��zk�da��pϑ�mW�}���W�
���z���r��,��{��\��@�BD����&G����î
�Wt%ft,�)W=ޓ�v�'��pV��X�pP���h��G��·�W���Q�����Iuv|���k�ĭNKV�to16{��Vt�f�oMCS'2��rBv��O�$�qM�g���Z�';�y38����L�����W�W��Ў�,n�tAB�Iomlkޯ�j���r�#�}�|��6+���^k��e=��R��C�`���c9�|L��q̺ޚ)׺=/�n��d��c��l��eTO*:���	����1��Mʁ���S|��9��r�n�E����3��Ә�Ǒ8��H�T�
��3��p��a�K�7�h;�XXm�L�u�Ɖޒ�[Q��v���v�f�{��Z=[�i�h��@W���r{�E,���u�C����.�Y�fM'j�գV������3V���B6�am�T����?.�u�5��G�o�c��6���Hl>Wۘ��;��g�Cv�������|��vWU�b�󥇟[
E��j%���خ�	O�
�Yq�E*u�r�@�� a�*��z��
>CZDE{����bڽ�*��t���K�g|�|�'�\M���3���t�1N��Rw�b�m�.6�<|Ѩ� @���K�Ù �wN@!a��&+������t�G���y����Aҗ��Ţ����w�P��{H�H����J�th���P'������J�m«H[�oM*�E�:��h�aɷ����A�V$AL�NÖ5^�c�mq7c�;v]�ذ�o&Т8��_������k�N�Wh��̘!�3��#>�R1�;��{��T8�eĒ�YU��|3��f`Vl�A����}�|�X4��i*�䦬�8����W,l��!����#���at󭖱e���%�sR	���W��,���=��:v~tn�.ɇ���a�Ji�;`��p�k��S8����W��(+?x��_�0Mft���=:z��Xǩ�N6�eR0�Z���'1���;7�h�8�rP�J������+�E�$�p��8a��M�9�)1SA�#0�����j���*��A������>Hu�	��P�x;��n����G-dV�_"=f,V#ß�;=d�m,�ŝu�_�;`�c��㷳"Gh���v�v�[vA��{_8}�x؋�k�Sem��5�����z��+�fX�5ڙ-�n�.�ڭ�Q�?7����҅w1�=����q�=˩�	�[Ȗ�ǲ���U��νt]t�ݖ'0�����
���W��y|cX��F4蚬��P}���^{ks���Q����ĥ񳼴�l����n�D�'R�+R�EV�z�gה�k���Y�͑�����{¶���S�k Lv��7	z���J�]o��y�e�J=����EM�3�(��k�X(�G�p�m����3��BC��T}�}�v\jޞ�-�S��eq{�+��T[ڇq:��%���vu0�A�(��ڡ�8�."_Iv�����) f��}!"���\^��(��?T��rj8�اJ�[5��繱��I��sy�qe���C<�R�:��G����B�ﶓ7�us����4G;��wς�F����
)��+��$#�1ΧI�0ņ\������5�&�3*b�ORS���S��
���Y�U6��(��O��6�q���u��O���)cu�3[ɞy��=:ꌾ���7���8���2�@��:f����5���f��CK[!�x��g�Y^'ϑ�Iq�:!MGu����b��dB��g�v�1�� h�0�7F���M&Q��g��<9�����5;��!3�f[	�E�1%��W�jp�F��wqɸn��ى�g�&8]E���2v�l��Ȏ1��%5��v;�qi���W�-�z��j�\Jj�C8�9c)����"9��P��6X�������ѿ&�V�=���n���:Tq�{quV�9kZ逸w�o:/��g*l��ꥡ�Z{��NN(	j���1\�|e��:�N��8abC�U�2Ú�Y��+���5�<G��*�@��8ާ�o
k�tKBcNtǝD��T�=�Z./����0�����42��y�f���b"�O��И�a��xyນJ��
�r�s<gm���������T��t��x��C�ۇ�*;K'ofN$
�o�t�mu��(�܉,��Q��f���N��Woy����'_���ҹl` ���T��_�D��(�)b�e�m3�zKD����gu�+RT�<�n���m^�s�x8#B�]��ۧ�� L�hv��v�U�+��a�9��Or�	q��rU���os�۷;]p$0��L[l�N�i��:XT�pc�]�˸���f��Í������+�5db���t/��C��%c���.�9-|]ǨS��B:��Ugn]e\�9��؉P�cﮏu��y���Ou����2�pJ�}&^�P�D�ꗽ�`�f��q*����a�J��楺��mJm��R\���ŀ��AY���˽ܝ�����Ak���j�7�ܛ��&|����^�=�U��ڊ9��'��cT�v::�G����Z��)hM�Jb�u��ʟ`�5N �:�$�3�^]1��i�Ww�xѬ`{�n�װ����~�սV���"
�{U�̋�m�e�Q̙���8�@��Q�*M�J��:�gw]�f�t[�Հ��" #q��i��֧n'��,.�u���*�W$�
�8o�M�^]�Q0=���н��I�X!��1^���!B��#���X�T9�M�/��nN}����2%(�.�$��aֵyO��|s/����e��7nN�@[IU���a��yN�H����
ym�%�ڗPܫ����T��7ɔY�z-j�i�RfFʴ���Oq먫c��]$��*�'�{S[�i��v�H	KN��g
Xs�\�њ�J��'gd��y*��hn~t�ڸ�ز�;�.���t�7���.Y:05P�Q��\�0X�uֹ����J��MC���뚇m뭻ڀoQ`9
ձ|T�o���6�諹\
�ڎt�j;g8:S)Z�S{�eϏ,��sX�J��$���Wm:��o(�<H�ܚ����n��{�J���ׯ�'h�[ɋ`Igv^ܕ�1&l1�I���V�X��ΰj<�ֱY���7�!4c�{����@��2�̷�������nw^؉��9�c̺��/Z�w���c�N��n�z-�tA1�1�l�x#�N�:�����/�lZ�&��Ol����A�K��f�I�Ҳhe�-e�0�X��U�YJ�⊪cF"�4`�PUb�Qj��4˙l�R�UKP(�iU��V��eE��*�ʑ��ZUJ2���j��+kYT`�T+6�UYYJ��*4,3,�H�cV�E�cTb��ڰ�C�J
1��%���ZQ�[F[**�� �(
1�-�h����mKR��J%�b�+J�*�ѩVUh���T�ȹ1X�TUXָ�����(�UJ�jưR���T-�+Z"6�U����*3�����FT*����TQ��B���Z�[Z�#Y,�r�8���fR�m��"�V(���2�b�m���TUjV��iYjQE�������F"��m�X���@U v'��3����S��"�1]Z�b�c�ɾ���"�+FT��7�`�-��iJ�������I�o�����!.���������	;�+�S<	�\W��+s&ϕ����9�G�Up�'g��ү/���F�B<�E�l�Jo�lc�:b ����_�熷u�}��!3H�RF�T'��P�32���by��ב13�xTo�Xhfs��>u7�p�����O�J	I#'�',JNf^�4�}#{��H�U���%5_-�a���)��a�U{hdt����1־pN�]I����U��U���(x���K�Pera'�"t���������B7I{9pΒʝe��l�!ŔN�y���B�1��j��q�Z$�d� �g
�wvPKcS�:h���&0�[����?����q�~���4�˱`R������k^�}��ng���\t�"����9�F���F+�&:�A\t��{]"bb���E��$3t�p5˛X��f�Y����������aˋ<k°�ӳ��1y*�{kN�ڶG�������F���ơ���of�n]e uD7�ȫN��0��N�"�/<�r��jR�d��U�����B3/(k�(���Y����Nլ��O����}oQ�[��:�+�p)w�=(�
���U�woj̎�#�4��&T[��%p+!�3��	�.0k�9�gWtD�xj����s�m�.�0mݙ�X�d�&n�4l|�� $�_���^s�M��f��ߚ�۝��iZ]JcE}ʀ�I��z@h��4���=�|r@��kπ�ط�"�����V)�o�E~)ծRI�~=�����K-���2t�"�tǾ�
��,�lw���x�zӥ9�p�5vzU�|�
68XufTU����owu���Ƈ�s���	��_d�s�Ʊ�]��!�c��{T7��8~6b��*�zs�n�F-oI%�U�T)9"��B�U�_]}#V�l4`�=�w�dg&��z��p��1�]gd�.���*�lp����L�?Wyo\���ٳ�>�P�^6�u{�^v<X0�Q��}�f1e��xJ������|a�����\�-gJ����y����P��<N�.*���nL�_�f7	[�Vz����Cғ�y��~��e��d�Y�S�6�K��
�<���#gG
�YU!�N�q��6���h�ovw��N:�6��7
�����0�mT_�h��m!�R`yw��@$z���˿t�[�k]틎��CU��ޘ*h�í��>9� x�	��ĖI���gV�Ȑ��89�6�4a���+bO0�p{����\�����Z�mv(Íw�������ɪ�9���f�Js�ܯFRf�T�r��6��0�7�v��G��}�]Ѣ6%.�IR/�o>Ϻ�� ���:;<�}P>H�9+ݚ)1O��밖z�GQ\	{��s\1���-�=_,��"�S���"c�9S!'Nn �f^l�e@Z�rz��y �xgS/�� ��w>���礱.f#^V��l)���D�����W���k/F�Is8��0x*���*wgĄ���%a�I����.�E��z�mI	����ͭ�]tL���%�ʡph����z���*!�.�����d�-�Ъ�fn'Z�[j].�����9�]m���^G��#Z1��n�e���卓`"X��.���9��:�o)�(8��Dst	���� �|/"�t�c߼B"�.�s���6k�,��7-s����Jt�� gt���:��N وn���vg�rt��L�:+��U�k��v�O����(�C�
ۄ���'zP������}%�g�׮h��5l�.#���p���@0ʇ/ؖ2���@g�ux���S<^��Y��߻�� �h�|��kb�-�%b&��2��o�����JW+�62�ms�51}wQI"�o�Et��;Mc�-+�E�����t[����"�:ps�ȃ��N��d�z�۶��]	zov��xW����\SP<+�V	^�꯾��s�>M{۽a�L\5���Eٟ/+����fe�v��u�.�l���/��02j�1�:�V�a�%_W�r����Ӕ�@r|� �*���%}�<�GJ&���٢�0�葮�G�mSG]�҄�Le��,��#��|zj�1U��?���Usx{�0lN�g;���������\�ML��aaݦef^PK�"�^Te�zx�w�J"���@fuVu�y����B�7�ECwP���tQJiL�������i����5Ƌ��a����r<���.�(�#�O֜�m�!�nDح�%6�0u�y=�YҺ@��#�@ 7�` �.bD�/�X�;��eC��;U�y3ԝEh���vu>\�Z���܅��ё���@�kF5J��I_>U�V~ȅ���g�@O<�N�S-�&�^��r�t�u)�rUL���]�F\�)�5?nE�&'�]Q 릩�����'{]���t��)�b�'V�9T�"�{�5}1͚�ne�ۛ�\���R�R�#�;޲�G�����U���k��ɠ�Ë�JZFЙ�ubn�D�I_�;K����}1^.���5R n�S0��@n��l�j^��	�Ҟu��8��&���'�}:+�;D��2	�؁���&�����L�v��YSfV-�ͮ�� N&d���n�'wM�x�$/8ٶL��������3=�ݺ���ɭ��
n:��\�S�D1V�����H�� �$�ipvȗ{y�oЏ�/|0߸��OzPS��(O'����^F���lO,��7Ξ�Y�ܢ��`�9��b�>Ɇ.��V�g'~҇�f�:�"��Cl�#�����O��}Λ�6����x�+OV��f�	ui��|7|�yJS:�q/E�}9z����TT���Xm��k�^��8�s�(C�V\՞ү��+S���\�ʿg�0�&�]�;>�4�pԾ1j�[y|;!͵��R+���5�	��	��(0�V߻s���U������Xy����P>u7�*��v'��e1��J���Hͭcoo��d^����]z7�O�n�3�Jj��,<7��1�XЧ���=I41Wo��,�>��x,
��؞
���׉�c�1�]�(�&$�\<�E�gG�f�N.s1��؞i��i�Y��iތ�9E���O�d���ԨAwP�!bm#�W4G�I��P{�c��$�&9g��X�A|C�͙r�{�v��y
\WL���ւo!j�x ��:����v��-^jӕ�cvQ�X�e�u8��ˇe�j�\冓�+s��T�k{/�G����ɮ=D�Q���;#f�S�gHvU>W�	闤��|  >璫f�o���#���g4�*���tP�" }/�\��.��X��kC�U�MHM��i�[ذp\~�
u�{\T�k�5�3��q1�S��
�n$�n�z���WRgc��T<�-J�q�Xv�$P�J�E�xP=mހ��y�EE�f8E�S������ێ>�g�5zCB�n���C3���y1|STW�ԁ���u�X�,.#Ϥ��36v��D����r��<E��>fw*�\��N�MP�M�N���s};�o��'C����K��\�nP�,�:+~������ζ3$~��m�q�c;m:;����yk&c4��t����sV��Li�E��!��XY��&1-/nm.ćL;��G:��C��K�U=���7���Cg�#�Y)����2��Oafu�[���6Y�!^�0xSrE��u�U������]�f:p��|�O&�Y;lW)�>����do��ڿ�r1:���THB�f/�_�j놌��+�x;b��skl�h؅�Ȱ��d�r�UJIz����ktsr�f1@�:\w7z;����6�C�.o�]vze�hv����=�E�,L�q���:��O���Y̐�mZk��cY�nV�;��o7�2I��ۤ�VЭ��؆Tv�j�|>��CK2h�}��e�����Hxzs1Sǔ^����WQ����v��ˉ�b��{�o*�`���48˜g��@h9�H�P�&Q�-l�f�'�XxLd쮦�����ݎ��f�iVcf����ׁu|��ս��bc^^A�a��YF�kn7r�V���� cOr5�]�䫫n$v8E�$���ن;'A뚷1Z��Hm��3)8��V�vi\k��q��7NWJF�]5�g�*Գ(v\���^���\|zz��P�rjO��J/�[�	�ܧ(��˕H�B�*���s�/�2�r��L�z�]��4�:�@y���FV9���"����V}��6G�ꅅ݌!=A�bz�t��Ll�7���P�@=�ɮ�]��g-�^^	y`����	�����}��ɞ�=1�&z���^{i���%Fu�B��z��h���s�.��U��v�j��b�{mH���㳪n,h��%H��|�����vƜ����N�U�X��ślt���>��F������м�;)�`��J���w�{�ms��.ј����9X��p�&��C3��1���뾖�諭���g�ٕ��Ȱ}f��/�
bPG<�a`����(�7U{c"om[a,vq-�Z�{Q�A���M�9�덖�x���ٙ�,~�l��0�^���G������oװP�p1*_i�5L헓<���tI�Uˮu>�29��Tf��ߏ��.��S޽���~�E-5Q0�:���O�q���<;�2��mD�,㣊9Y�X�� ��;��{R9<�~����:?o'<y�˒���.�����l������Q�ltUf���y#�[m>���څ5�)���t{4��h=�u�gϺ$� :��u{��U+�o������p�ڄ��\��ur�Y
�abew�{d�-�Ɋ���ˈZ;�>���W��n/!�L:��;�2h�h������Z3~��T���
��.��}�PS��Ss�c��(���z--�03��}�S�;E�]~fi:Q�2�'�*,^3F��&�S����Zմ����lQ�V�B��xs3Pfu	\H�z'Pq1��xH��=�j/~Y%�7ڷ�B����S�����ƻ)}ڔbv�36t���G���N��]�����>�q=�>�4$��F{�N������`x)�N�0z������^�n����)�bk��W�v��W	Z�>���We�
���:���i'�z�;L�Q��I�vWƖ���T8�E3��̆�blZٵۻ
�r��$��cP��w^�y�¾/�n����Q���4�#�\�<Y���<sK��r����5��{�&�UJ2�&r��]�� ���Q�Uy����c5:�Ֆ�8�q��=��x. �L�a)���������8����b��������9힓B��ݝ-
���VVKOTG1�P_`�Ys�V�+cL�36{�s��XؕvD���Nދ����E4�o*�Z[C���$.^�0.�f�M�j&�ۋN!r��M��i����{�r{lk�n��A�T^��JF�v �e��ͭO^J� `X|���/�Y �z�4���%�Oy��_u�B�
�Qڧ�kT�8��Ff�@����W�`~���.]͘jWHB�e��hA�uZ��{���������t�������gRKƻ_Go�=
�
�G�_}��}`>�����쟾K~t�~S���K�~�|$[^�?_Zi���Xq _e@�w��bu*�d��`J�c��-�3T�_`1���g�~��Y�YQ׾��@���(7���H�ە'ΣK� �	V��k�>����:��-����[��hJ�.��.f\*�X�p9,n�WU�⪝�x�]����޸�W�2i�P���BS��#�].f��3��5=W}�۳�)�M�z�\\���8�Qn���T�˰G9���7%�L�$�5�ϭ�XO3�|�]nz���u���݉�,�Q4=?O��Q4��{��7l��k5{͟������Ϛ���
Q�hmd��pp*�h���v���,Q}�i�}x:����u�����Y�g�˞�q�A	�S<�����ʧ=�f{j�"������y��yP0�힡����=��gAZ;�2�̹�5tnh"��rJYo$���>9��k#�/�������7g'���[9�t���U]*z�+2�Go��Z���q��t&�J�!�4`uJi�����ՂV
Ꮷ@i�p��&�bx����˓c��Ƈ4y�f9�8ò��f�����X��e5�R"4��ʳRZ}��n�z�Y�ʫ.���@�� j x_\]Q��W����5ʹ��y�:/���Ջ���7���y�V򳲕��*���l��`�U��aY�|�}0�:��,u��&��-����N�@rw�(]�e�Z�y�hC��f�͊�Ʃt�s/l���δL�;7ST�Q�+�C)0�B�:�j�g۴�މ�B,܄kvX5ʖ䲥���Y��{Mv�(����4v�=�`KoH͉�V�Ȳ�3ź�����)a7C�\;x����n�/Rߜ��3c���R��˥��rT�b��RKY¯�\���T��ە:ff�ʟr��5�>�%��}Nr#;j	��d,қ{��4����皣� �����bX��J�;�<�u�֒�X<��˱p!���*d�L��Մ�zi�v$��<AT��{Φ!�ݼ���eb��vݥ��l5��f��n�)/g|Wlʇ���v�+v<���/B�u\d�/&r8ju�V{Oo������6�6]����x���f�h�K�y����E���I�2��#B��m��6�k-����_A���z�_g�Z�]���v�N�z�r��跘�Zգ�G:dJ�mX/G`ȑ�Z˭��j�>��F� �>y�}�IX"k�ro!b��td��O�;�NIT�;odI"�>
��o��SA�Ž��i�A})���3��΁Ҩw�N���oR��8�٠ƴl�,LJ[4���hc\&b�Y&��]�D`��ٟ$�r���C�Ǜ�V	��x¢W5W�:��C��%�n5��彚��u��-����?�_����������z9��&�/_Nh���bi=T�Y4��E�N���wX��S��۬�Ȅ��%M�l��*�(5t6֗(u	�Ѳ���%jt��N�E*�T���y�g跑n����iW�ݲR�[Q%y2SˮU�['�S*+��	�t�L�:��:��� �\0p��"E:����^�E�X-o"���з:;4L�V�n������gH+84�C�$�}���d���or��8�:���*�&�uN��G���divPN��b��]BwU�!��G-Wjb{Z�
��G�f.Ǳ��O<���x���nXt �r���m�N�z���kY�;0�os��Xt�*0�y&e�W�ځ8�Q��NQ�lΣ�/uM=*�3��c%��;��suR�W7���(ޙƪnp�������1�'�,�1�5�R�PIe����������qk��8t��-����6.�\��ms����˥�ũ��6���%��?��Y�`���/%��cѵ����$eB$������o�����ԍi[iF�lTkDUDm�D���mEDQTkC�0�,�W&C�X�ڶ�����[k�(��A�YU���D�QTU�ڢ�*���3`��b�TEE�J8�`�R�X�˗)X�Th���DTUQV6������T�bX+*����Z��2fbLQAV�R�5���IUr�(��E��ʪ�J�15j��Ub7M0m�aA�Z�ӓE��F�eDE��H����0�b����,E�R�1Ƹ�R�E!�E]R6,�J"e�m�PQ2�X�Q�Dr�m�Qr�b0V�e)��Qh�%] X���2��Z�QTX���h�(��ČX(�J,DAQP�iTC�(��[Tr�)�F�*�b
őT�D���\Ρ-L�j�ʣ�rS�q��y�8aS	vA�`� �����h��v
���u�5���7�X�������/b�1�O[R!~�j\;�H�|]D�1=��W��MjM��vv6в1&�����y>��j��y�a����e��~��el^L\��х5�g,E���{��[Kԥ^����ŷ��W��m*�Q�3�赂f�o;�%H���.��X�kc �U��HT]���u|����<%@�}���s֧[�G8�+�6�%)���}qѷ��Yqɽz���w�.��s��Kݷ+���f3���
�/������Vy;[I��Nc�����%��1Tl�b�����p�o���Moj����y*�1|��k��r���#y��y%��5��nt&���sq��P�FF�H򔸂w6�&�.�<}<�K�o������R����ǻNS���\�7}Ar�� ��Z�ʊ�Fw�R�X�P��ιh�W�4��\7��8Ɋt�3�k�0u��$�O���W�d�Ch;~{��0��h�A�L�+�2h��)���*�j�ɧWe�)�i���iK82�Kz�ډq㝽�M�����j�V���F���k7  ��\⹉�����`f±�EV�-�մ�Rګ��=�}�G���u:�<����xF=�WL���.��)�|��=N�	��V2��UG069���OTc�W��4���Ʀ��3ٗ�)�	<u��泗�ɗ�i�:��|�SqԞD�
���A��l)��3�,z觷K�l��R��Q���}��4��CP�Bu�j#�߄F��ѽ6�]��ʷ}�x�>�GR��!Ym`3�Tr��%oɨQ�)°2�En3���%�~����~�������ڍz�V(��o�IZ�p��;7QAT8���I�ALV�r��`)������>(�BQ}Xf�oq���wx��wj�՞�_s�3�I���KGh\t�uE���Q��d��a̅�ƥqѮ��R�s=�H}]��ˆ�v��-+��s8��:��9hg�5�l�c`���i�.B��}�
�k��m���v;��c��k��d����k���Sp�}vչ�%
�3�����U.�kw\=[�W���^t�]L�r�p�޲������`�f�a����MśӝeMHo�Mo��u��f椻X�mn\����7�%2�vY�(-�j��ٵw(�R���>�+;��'�W#���nn��t_�|��O5���4�t��T^�ey��nvuMsŬ(p�D�Z��y�žq��F8]�	���7���[%��d�&�AV_;DŖ*�����"������o]�I����n#f�7Pv�!�ܸ��k�|g�+��c�����	z�8�s��&��}�įww6;
91bV�\��ǛX�Ƥ�����N\���K+����/�:�WI���S7�vCu�V�����Lr�	ݮ�bb��˴G<��~��)c��lT��O7�띫��p:�9�l���<L�q�ДY����-K���ET�c��"�s�9�:j3^�yQʅ�N�
�*�v]��yq����m�2F���������&|��r�m����~�l����-��s�C ��s�%^qO�����A�w����b�:�J��!A]S�N��K4����e�c���ѫ�f�r�����u�e�2S BY����29�k���{��0�vHݣx�ϵDa'	���Uއ[�6�\��]��Ӎ>�*���;驮f_bd[����pN�Η�0�+���{q�<�֞L���U��Mey����ʶ��k�w����Yk:ȿc���^÷�T��[4Ȧ�.ޝ�iV��p���ڦ��'�*9��/��+��Lܰ�j&ɽ��/���6�b���p�=�C1q�6���<��(/dE��=su��5=X�c������[y�ؼP����y�zM�x�_z����:�+b&�~=��Y:
j?)��y��_x��vlQ)���Y�jz�'���O`�=�j%A�j�,�V�Y|��-��I����9��3dրe�k-��qj������\7�
������8�ܚ�n���n�ܝKeg?��{����Oް9Y��P:7��U'.zea͵��MU=���G��j��I%,��8֪ˌ�s�jeW�9O�����]�sr��[������l�L.wkZ��MC�]p��W�1W��L+�=bm��7޽lE��1�� b�q-�bR*&%�*+x.�V�e��*��19����훁Q��'c�l/��@��sf��d�9n�ӓhz����Ýs�b�'rV[��l�}�p%��A�k�XN�3�ٻ{.券��l^�}�}.xtn�x��~��N��f_��:�m.�)[ϙ�P���]��^����y
3��n'���5�'��^�ci��pʇ�2���cKR��}醻���`����皮f����NYU;o��ks6��4�c4���z��H��g(k>.D� ��;.
��)q^�+��~ڶ����Y����Z��x��ߺ]ã��ٻ:4<�5�V��6��֞V�������S͔���=�����3��^)?[,tHj�t��V�UVZ�uz��U���b�uz�b���x�\5�P��j���FG>E��^]�)���r�b�[���U��f��G�ϐ&����}雽�9^��j�ۅ6����7��0}S�Q��'����E�R�r�L���|s_/Uqo}ǟ���/��Y�5�����5�t�t���Ԙ���"/E>~&���A��8�YY�el�lHf
,'x�ꙏqL{��H�6t��
Jyu�A%�b�e�,+���xe��\�2�n�r�����GW�k���$�֓P������-�a�w؏]�7ܕ���yl�ԣ�����<̑������\��vC{0��/f�0.:7�@�ox�Ly�xc�\���˶�&��Ú�p�97�
m���Z�pJ��y��z��f׷Ŵj��sz�N��e��ҭ��M+�qݷ��j!�q��m�by�T�dd�bn�K�Q��fG.�\��78�'���]��u����6��.=�ϡ���</9FD�D���7�ٗ�y��թ��F{b/�{3bsq��Ҹ'�C��XVT�һj/LW	[����>ʉ��s7F� ��Rw3�b��4�W&Rcg��*_����/�S�_R�s5t���Qr�id�k�=ʎt.�b�P���9��'�=���]���lv�7<�q4��E��f;[䨾]8�!7�)u�V�<W[�vV��W2�*���E���5�3X�b;���!p�g�{Ѭ�PTt7�g}���U*xծ�}ǻ��K]Ł���M��NX�,� I�,�����<�E�%���n�@a��"��tޑ7������f�s�q�Ӟ��Z�m�8�4������s&���;�j�GYBҩ׶���QQ�6f���-�]ίU}���\O)�W0�zD��}��ׇ���U����[����o\��{^R�D����z��q��p�і>8���:��U|�������ڂ`�`}%��x�ħu>V�b^���q��Cp�[��or{(��'X���bG-�]Q;�W�n ���|ب�o-�\�uyT7{�mD�ݞ�,!�es˚�VMs�I���O.:�^��m>����S]�	�}y���M��EF)��_�ߚ�/G��C�N��roݕ��|� o7����a]^�κ��+���L��[�:0j���F�DJ�K�}�b��
޻�&��c�ەe.�,��л�֫�:�щq��Ѱ��h�J���K�f.{��*���4bˌ��g���͔�V'�CO4�2�'.U��񄫌'��v]Tp�sS5��j�܁4�{���+�V�X>�=`{�%���B(t�a���Zx[��9a5���B����e��4�7s4��hzɮVRwe�{5���8�ܼ���O��z\ ���^�쑸�7A�6I6�J�m��yo� r����r�'t�N�.G,@G-���-�Xt��'B���(m>��q�p$���%����}U[uta{�J�^���gBk��Ӹ�q��]��"�
���ˎ]u=�.O"u��Ԥ�p�1<�q���r����IӸeC�S���8F�-��sv�B�wn��q�4�]�GsU��bw���g�<��=!��v:q��Y@=��j�1ڱ�"Z��ܨ5ξ��W�j5h3��%v��^JO���<��#^��r�z���W��~k�Ak*;��c����^����5U�Z#���wk�������S�犻�-��k~�h.;G9���fli(0��ݑ����ڈ�lU�Z-���\ͥ�=�m-}'����O����ث\�SSj�,�W�:1Z�[x���ϥ�����=�y��M���̙���~	��Y���!v�Ź���y��_x���n*X���7�5�Z�VkV
�}��� ��^�*.u���%ki;<�ޖ�hp��K�������
��`?M�2WK��<�d��Al@�9s;'n��j��Vt��t�-�v�}x=�lP5=���]T6��;�=B���Ϋ���qҤ\��꧔6��8��Xh_<C׊�a���fE�tk��&�oq��ܳ4���W9�i%?��ﾲ��ŭZ�[�s��G��u��jѾb�B����������s��y#�z�����og'S��7p��W��ӚN㍄�K`loT����{�"^]gZ��I>��:�=���f�i^��W�2���ەK�%Na�u���[]�&�.b�]�WkZ��ڌ�Ϲ+4+��S�Lu�JzpQ�0T�g|��l
/yϸȍ������/�)�6�[��a�m�)����1�T���7݋U�w>�k��UMɨ�O� +�L:���xԩ����V�ݫ�]�z໅_w ����j�xqc��[�6*j�!����H�|Ъ���֦]B6C�:���.��U��^Wld�u��s�Ky%O%�(V�:��⯻[���)���f�U�vNѺ`��\�M����綪�s��skLwS|�����W�5ކ_��Yͱ<D��^^���k0�ͷX�����V�'SyRN�:פ�P��JDe_@��y�ڇ:mi�!�������'I��|^.w'Z��zv&b�	5���9ev]�PT���:��Ë��榘���R4���vp�
���ވ����n���fnƪ����OQ�/�(�{֪���f���{�T^B�f)�k���y;=�w�d^x.�;���dbuc�rB�dݺ�M�T��&�X�������ܔMŴ8�ܞ�3{~K���s�"�����<�ș/�^�u"�ޒmW���^j�4��S��P=��]<����[�%������y�s-ҿ�5���!���MvM��:j�0*~�ꞝ˥�m9S��>#����Ծ�>t5�b��ɸՖ�@ж�	FN�cA��-se��՝1�����)�YkGL+{54�5�v���%�o4:�ۭuu7gU��v��N��28��Ϯ�.wkGL%�U��M�
s�4��?Vh�wy����q1�R��=5�$|��P��qN�Jbf!�Tkţ'.����;W�y
�݅eO��ڃ	�p1+.��߾�]�P�v��yB����ԣcШ�7~1�}�>ެf5�v�{�C2��M��\��pc��k�C�Zc:a��6�')��fЫG�!H���U�n�铴�n��f���$f)��ڻO���z7�9Y�ϲ��2*���0E�������!]R�<�Y��y�(�,�eN�������W�N�����ٹ�fٟd�	y�@�u��\o�z�/RND-�,q�q���+ZCd����9�dPۢ1��k�ŝ�F�two�-Z[xC�Qd:�s�k���`��3Wj��N���N��w`쨢쬻�n4�*����b��\�{�j=L���M3�R4wTT2�l5�a�J�[̒��bL2��5r��L�d0dN�;�Y��>/�9+���Ϋ��ηOWN�Z���;�A0iXx;6JP��t$�E:�*�����w|`�HG�6��^Ey���s��n��׳:j�z󵦟"��c�������&:�2]����M7X�A����婹}
Sк�h+��I*wa�/�f|��Ewgu�N5��7)��q�����|(��.9t8rv��j\��H;�Jn]u���f��|���U��Y��5]2*}(�읛����ԫs:�G�z�E�#�yEu���i�h��T�T'�X����߶l�Z�u���f�2�øN����<#���Ei�:�����*+�/���S�k���:4^��B"	��n�6�Y��VH�s����`0�ɾ��8�߸�2�@�'$���tDƇç�\k��Mlp��9)i:���K��Vd�O�a�[�&-kN�X��;�;lX562��]��\\jq�����܏�W"`t��ٔ���������#�E%�W,�Ö#�GpO��&J�f��gd���]�J��9�G]!�o,��5�iӝ��c�6ՑE��ԍ���G,�c�F���%����R���*�R�:��=�=�9kY�=�_ܖf��@*�(n�B�vnЗY�@zh�,�YW@�枘�3�oNwop�LԐf\Kp�pmR����J�ko@䐵��y�g!y�	/�.µ3!�0�j��e�;01��޽�ޱT���Z��F)�R�{��3+-� �g�[
n���ّ�0�Vzr3�{X�Z�d�Ƣf��%NU���:{���22I���AM��!�+R9�̓�����
=/�pu��Y=p$ݦ;���?�q�uZʔ)YlL��,��h�V����N��q·sc댘�x��wzB\��6�9�F̭�V)�Kݶ�2-�i�.�<��wi��f��+G	ֶWr��BxZ�8��p毬6����(����6���e��M�j�q1��N{�c�O��z<���d-�����[�ڷh�&K�Q����:L�wx��#8�	oaM^�m�z���;��f���gr�Xc���9M�"����������V�a��u6���P.�P��1�Ԝ�K��*�P ��Qb
�YF�,f6(�E��:M`�TTF+F)�Q6�f%��\J�*���(��V���DTUX"1 ��kUb��"ŗ3j�Ma�,UFj�)4�"E��Ƞ[(*�V"���IPZ�R�)dL˖,mX
�Y+Qڢ(��T�AV#E���b��D����:�u�V
�"����EE�Z���Db��L�Eˬ�0�T�mDPDU�J*��Q����b���mA��"���eQQ@R�-�Q���b9E,�ŕ��TPADE �h�be̵�HbU��bX�Zb��"��Ղ�mDR�D��*�
����L��X�5*i�1c[��1��Ul�Is5�AQX,Әc%V,TV(�HX[,�-*[J�,���=�y}�S����*l}˙*
�O�1�*#YC�հ\Z�6�N�1�q���ǣ{�5�&wd����Zw+J+�D}E4D������I�n-3Ч���G委�i�w��EU˹����yK�ض�<�"�b�!5��{xyS������E:�Sdw[�s��\�]�3��N�Pm�-5�˨�3s�=�;xOD�M=�
	[���y����|5�5��[ϵH|/\7�]�k�;��i�1��{�Z�nڝ�d�~����c'�0/`�|�.WS�v;���y{x��"K��y���x���W���\v�(}1�����{q���%��`c��;��G4�}v�[k���ǅʹo�Ӭ��8�����u��?�N�ԅ��ϔ,��s���˄�����K6`���wW�U�b�̃�慼4��=�&�*5oP��s�gO<:��������\?w��^�����gRס���lL�����[�O{��}��{�� �yq�m������1`�d��F�+Cr�iѻ#�W�|�+˰_['ߜ
��{l۽��}����[�B��!��N	�O���n[�&���oVN�|��h]Z�3�Ri�m�;����c:���W�j�hl��,,���vT�pf��G�2�����j����c���QT��3?G	C�>�*N9��[�����SK��z�.�MG'���1n�c�:S��a+�G)���f�\*-sˈZ;evθ�[�yvꖧ�n;U�_��O���K"M`!%�F{����y�'�noV�^�w*�8z��G9�h;�8O�Zv�rwhw���/��ĳq�;��j
�[�/��I��s��!�L���uCv&���sy�#1��W!+��:��N����e03�ݱ�鏺Y�I�j�/ N[����Ubkm{IWD�⩖(��^�^gU�8�ή{_r�뜄؁���ߚ���^-���B�3���q��tsZ6x�����;U��iKc��:�Wv��ss��8��dG7������������J�"9 .7y,�k�^Rwή�^VJ��jz���B�+�r�v5�h�m��Do�dµ;#����w��+R��p.�(u0Cڬ�"��}�8y]��U:l%L�/�<���ٝ���t*���gǐ\���(�9#:̸bJG��8,�P�݀\�9PEJ���'tK?.��f�[�έ��������@���U���g/o%���K�c�Բ��^�^vk�)��aV��}zy��[����0��:ώ�=Y|q{HSh.����iw��i��+�n�;A��͚��X)��c.-��P����gBh8����[^�ou���1���+���k*�s�H~T%�gV?r�'q��'��@�f´�ni�䪶��n�X��+������c]J�)1|���aK{���f�T9���8m�q�6��gF5�柫����`�ϫ���b�x�Ln{����Ws�Z:~W�4�J��r��?S��;r�J4UlZDl�+��¢���9�\��.w-i�S��W[o�y��*�a�6�URɘx�b��mfM���0�p��V���3�m�>�=N��t�H���k[kޝ�j{��k�%���W<������]����P�A�I�akOwaT��S����>;�fU���3S����7c0��y�#����	]�� >[\�⌜۫K��y��u��ɵAa��Q�v	9=[���i�ΌYҮ۬N��}�Ցx�}_?M��+�\�S���\AK!_���¶x�'�*�o�\�����Ǿ��>���n��-<��p��o)7Q-�dOϘ�+��7�G���B�(v�/�_���zs����wZ�T����j�r�7P����M�T�.��0*;��ާ���l���m�78�dv)�{u4���C.�>�[���Vv�
��1Zz�j�����w�Ԙ�o�՛�K/Nf��iE�w��Z���l6�����W�~�����yy�%xWW��#�k��jN����G.ڈǇn�^AV4�ȋ�Uqѷ�<�)
�nb烢���}S�3��sU����~��*���r�@=����o%UZ/d��N��r��9˯�5��k�;0���!p]Qpttk��i6�%Vgfr*����^���������)����V�sB텋 ��Ř!#���طU;�YTwj�s|��\ fk����_;qvb�����uX���e�L>[��z����3�X��S�x��Q[2�E`�æ��u�!�H���_S5.�n�s���-��9�)�|N�[��KW]8C�qSr�wٿ�|>Xo,9�y�hP����ע�\�Z���M�M'ﾴ�fT��i�󪾆�rP�6�W��	U-Ho�J�����\}��E�k^�%�����VWڌ���j!9r�5��阀���ٗ�:�6��L9t�/R�}/�9<x+j�b��A]���|��Ss8.����cnu��亝�l�sc7�o�ô�B���O![<��4�ٍ����K����j޳7����G*
�b��P�9�2��6{zx��{J���^��$������1����9PuIU	�Q�)�FiO��3�70f��[�@u�+�=�Ps�}y����w��Q���9	 ��*�=0�*��k���m?T>GO�)k���:-�ŽW���Qz�������q=S:+=�x|�(���¯R��f���s/6ra���o�qӊo��G� ܻ�[�nX�%�ʆ=�P8�}Y�%*� ��	�m/FQ!�`��(��u�R�4�{�Z���G�mP;��]�7H��i
��� w�A�e��wy���	��EZ�٥��K�Cj�G%M�-�|��@c�[1L�:�S��;/6�G�@�W%���=��1�b�ǚ>������ߡ���{��|M��j�s��wy�w\�bC5�q�k�I�ϻ�����<�z+�D܎�*mt w�,&�udh��W4�z��{���x,�>:�\ak/��>�����tr��\>e{}���z�I�u
��%�VN����8]��q�9�bf��0����{7�l�{j��u*%.��Y-*޳�s��'��e��wj������tg�S��û-�!���CYٕr;�=�,��ΐ�a�Ֆ�h�1�f��M�Ϻ�n7U㌟��1_&��+�0��N����T	��8+�̾J�_?�y}���M|�S����Z�v&���.�4���̊�H���l����'S��/�ʅɵ��T���q�݇�ۼuGM����~����7�����}��BWd�F'�c�W*����|ƕ�wWVSݣ^0b�fXI#Icr:Ep0ɱ�%���QWi��Ε��{�(�����>~����+���	��Y:��Ab�g�����D�6H�+8���쐱�7��vNU3ٚ��j�P�-|�!�ݽ.�Q>�IR�KM���#��'�8$}�	�w�S��oV_憎m4M3
��r���"���.,;�9�^g1~�Y3��{_Ii�V)��.���X��g'�r���8F��{����h��)v�^z�س �M#8�o�8��&B��?5t�Q���,�-ew_E���V��z/���p#���ozu�w��\��U�����|�*��D��C��i]���Vg����6�b�Խ��=��ק˝��������2!�rw��n�RMLn��D��g�������(�p���}���Bx���a=�}���`��&qO�,a�Ԋ�#�q���39|B��0�;�u��(�S\A.z���~y���ǵ�؍{��4�K��@�}����<tf`�Cg��^�l����짹��Ȧ�!]^��P�b��o�*O���V�A9���d]��E&��-+�w·4��ܨef�P�=,{������jL�4�Y�wy#����=�[aQ�_[5�eG{KI����po)�M1�un;���\έ��o�ˣ614槡j=Zd�/��:��}14��2�������_�a��t���ӣ�*�u�Z��`�&��] 6��꼛x���ʾG�Wkx���B�[����vi\jp�ȍ9���@v�`�ډ=�q4A��bN����5Nl�����kU��:���b���po!�a�M�r	�Yw��#��w�񩾼3�;��is;,�c�+��s�==��u�+�={�]"�
���-ϩ�[�����YwO�լ��3u*T9�T�%��uCx�xi}����)�˥_yͮ!��Cާ��o�֜Ήz/g�%5�_
!��;��K�l\�Ԭ�ݨb�:�j{��W���f1`3�o�r�|�]�@��Zk�|X ��s)sЏ."�+Ɇf��Suy�W���5�2;���mh�^*�u��hŇ��e��:�ʂ�:�z�/'+c��Q})�o	U[��:� �^<�
�9v��]��{��9�z��R������2�N�+�BK<���k��m����7�n���h�|�ŧh��j�.]��(4�c�L���Q�ّ�6BY14DT��nR�o�S�$�+b��V��81���	]�v�#WoG'6�f?�'8GZ�I5�K���]�gn���d�W��䫗2��������{����A7�n-m���b��DY�)�����r&fN��hT������׊{U<y�ErB`�Q*��]�S�.d���*Ĝ3�������k.MvD;z������n���n)-Ǯq�6�]�8���|�,��5���5��vRkx�bv���8��4���[\��.�w��Ԩef�D����Z9S�m4�\wn�X�nEP N�f��H�A^B޽vb��=�F�_%�a*�������ܷ8�5���@�c&gx�#w��Ay���T�X#�XBJ}Bo�|gf��z���绦��\�N���*�݈�V� ��'����d��N�黆�9�&��˽�=�
�&4��<L��C�0��,���e��0b�7k<�����Z�G���ⲹPʈI�MCޅ9
#��Op���.��S�������8}\�uq�_��Z�u^F���刵:amZlе�lǈ-����(�ǹ�R��'0+|�g��<��s6u��\+zQ̷��.�&���t��h����W�.�\���v�z,�����%��T���F��YR�wy[�yE�䥳ure2��ƻ���;���N�*.��[���� �K�ޭ����\�b��9���;os��Ux���3�;��-؅׮sΉ�	{���v�����Z���xr�������-ꨋ��O�������t��SiV�?�U�\s��i���M<l�Gim>߂�B�|����
��f��+��G�]:�Ҟ�������W���^AʹUP�l�3�����Q�B���{�T�Wىu��1�����!=������E|�4���'9��]OJ̶S8�z�'�;Y<�yw�U+��[i�㷵=�����{��5Oq��<�ɿR�/��C�r����7ξ�I��.yM^<˽�{�1鋛�N쾜��A*��P*����˅���q����5x�r:����4��8}��2a�n�YJ�%#a*�3.��yn���;��ײ9�q��0$]��S�Wœ{��r���-��AY�(�����t�ƶؗ	�W:Ѫ"7�9W)]���8�>��YJ�|��PH$.��-6pP��k@ݲ��'
{�=�}�Xr�)�$*�K&�S�+X6�2I�Ec��@g[vD>,��E�j����]|��7{Wg�؞�+ �f܇mI���rcM��)��}k�C�9��8�5�n������@M�u�(�6�ծ�Am�)�45�c��ָ���NA4�w����+����wV�}r��չ�A��h�6�-㏤���
��{ՋxëEq�Oy�6�{�V�\b����ȉX�4iUޱKO$�*Շ�zE
�Ã+��n�/ʦE�bf�Rqaimv��hm�i��N�OV�xo����v\p\��E�K�ga��A�z']a��;�)hNG�]w��ء���}`��~d���d�=��s���w9WS�q�1h�e�u�K�ٸ�hy��Y�a�ozC�y���]N\���Pz�8��a+���!����S��-���DXy6����:l�"�H��b�8��E�؝"�2D�O��i���\�i�Ǫc��뤣�"�S�]k��Oa.�C�Wgv�n�Dْ�{B�a�T&LG7��s�t���s������b�>����A�wq���!�J�Р��Y�6����j�tq�L������^ѳ���h�,0(R����o�~C�c�wN�*��5gđFT�\s�ʘ,m<y��x/R�F�EF�!�����=!�U �ެ���f���8��e��86�8@q�%�M�%�A�s+��Z����h	]���w��3rz�=�Jӎݬ�6�`�H�8�X*Fr�P�"�ŧ�k��P��S#�Z�Z����C�-4�F؛�m�!��[�4��.:��wa��8Ɗ�� �.du��>Y*��G�Lq��'��Ӿ�E˛n"yC�dl�a�ts����֋�j�(r���.��X�֔�u�K`;Րr�
�5�:�X�ko�S�º�|�M�}��Y#���K2�p�Vg>�r�>&0�m|���z�=Y/���=wFK�q��=sW \ɕ2r�0.%��]k�z���B�\X���Wn���9p�����ge ���1j���7l�����6�&F���+v��ʀ��W%['1�����U��K�}>s��w6��g%�1�w�F*�{[�r��b7��wi5MY!ri�n�}�u�qc³I������s����8�߱�Q���%}�� �IⲺ�J�"��׊����j�:�J�3��v1�E5O���Q��䝛��\�F����	����@�*���];YNN�_]/�p-��x﷓�J��j�s�5�}�I����bv��U/D�ԝ��U�+bK�$�;�2���Սu�tK�s�-K�ު+9��ځ��}�k��.��]����S�0�)'#jn`��S֎oi����+�Y��
�R[ɈV}�o�}�?z~X1X�UX(T�c"����V��Ub�ʋ%e�aQ"��(�`PDq*,YW,�꒎���Q�m4�,�"��bʕDELe��m��"
�9eE�"̴`#+%@T
�`��QT���k
�Aab�j�Ŷ�X"1�t��,r�"�MdkZ�V)mT�Vc�[Q�H��TX�UUEuq��X�I\J1`�(���aP�Z�T�Ub�Dd���mb1��KH�*�cm�)X`�RE�G�(���R���YDcWQEQ��ed��8CUPYdX����V
c& �c��6�QRЬ-����+X�m�X���V�A`j�2��TXUJԕ%�U�+ƪLk+��Z����^�5��}���
��n��36�(�{:p/6N�x5�A٧�&�x��qP����c{�I/A�K+�RB�V�%,�$��%BnN(νXQ������%7�T7�8��H�r�|�i����a׵H���kdM�}k����O.�[�x�����掿��V�J(ŗ�N2�WE���o��5��NZ���z����
�}��j�����-Gc����������;��/��4����ɨ��lrʎT.�t���/�O�o�e;ͅ��~��?P�^�(���<��Kj/3�-�Ŏk�\��i�2�,Ot7[e�n��֊�o\�_v5/a"Z��ܯ�s���x��GMY�c��
�R尰�;x�۸�!�Dc����
5������8���޺B��t�{{5�}I��~��}��c�s��{�x����:���M`B���I���N�6��V(�Qs�6�1_]�)��^�g	��R�˯B�����z�����r�nqU�tqF+�ζ�b���=��^�'�3:m��������G�q��:;ޏ�'��ν>+i	�))u��p�궅's�\w� 3��^Ρي��z0��}��0��
�7�e�R�\)�kX���V7�yn��Z��K)5��p�ۘվ��4yk������v�9�q ��<Ϣ��DܛC���{�6��9jaC�lg�͢s�#W�-�{�4�M5���Cx;�2I]ƥA�~�"w{{�
f���'�p�=��+�wy�8J}*�P��\po�T�W�67~��Om���熻a'��e���q^�Ox�]b9G�ev�5[z�o�\W��Ѱ�º��'���4�|��ji^��X���%�," t�t�_(�{}��u�#\����Ϯ��v�7}��=]_�B�[r����³��]p��HV����˙�a� ���쿂���6�u�v2��ѵ�o����;W�B�v&)K<��0�i�[�����>g��ߝ�'f��]ޗ՞$=sʦ�Cu򗐯�T�
-`��c��K�f���s��(���ئ���*����>���#DK�;/�oh�V��f�! >6E�*:�b��6�#��kF�z�K�f��B��HL;3t��kZ{��{��:u�uZ����l��+2e�e����\�k�t/V�a�r�Rp�Q��4EF5�Ed���K�m�q�9�6��v S�;�ŧ�6�ŀ�ju���;��7��m�6kI�`OV���u��s�h)�Zʃ��y��/'10v�D�S|ͭz��`�章؋ex����m�4��;�;Y-߶?�+ �X��b`wR�r����3g�?�^m��sE/����������3h��Ҕ����h�0K6�s�&�k��z�9{T|�k���M_������A�o�}*�-j�0/y�ju�!0���w�J�6������]��y��p�V%E�����ʖkW[
5o;)vO>��շ˔�}5�p��׫y	K�e����b���Y���δ*"�*�e6�8�kۋ��7�
ܻk��
%d�����"���,dj5���_>k-h�V����b�p��-���ά�:��-p�d�M��v|2�Z�C}�v�N����6\���)1���o�q9Q9���[\5⼮��Nq��L�#ju�k�����堖��Yq��Y	�Ί��n}��@��yM�!n�f��e��/�}Ssi=��i-�\s����J���B�<D>��R�_v��:iP��Ň���h�Im�q��sk��ɧH�\��#��f`swS8{aԧg.�E@��,*�qԲ�G%0�t���y�����J�S�.̓�>[#�UMkO�}W�	���	=�o��x��+!\<0��+��A�P�.�M3V�/���3i=��[z�e|��sp��r*��{C$�i(/vR���!ݲ� >�/���z簯�x��;�y�?���[1��ɮ�&��Ѭ��r��4VD�Py�E]��{Z��Ƌ�b��I���t���1�%�n)����f�X��>8��OrqCu��`�)�~����K�;l��}1gx����pDڻ�@M��ק:Ԭ��͸���Yܝ��C���4��6ɯ$r��<�НmiY�����LE�:��uP�����q�)���G�ƽ�wJw��A/.�ݢx�3�N�*Lf�#�^#�h)�YO7�s�1e-V75;j�G����,5�H�ѰN^�x��$:����
wRg�yS�V$.֌4����v
3o2����ݜ���B�@*���O���D���m�ż�9�~Y;��h��CJ�iY��:��^����=i��[o�α��cs�D��[ۣF�Y����k��ɵ�#ޞF�f��Ca��;i����n���.lB�~�z�1Q��H��m�7e�U ��P֭.��J>p�*=n\�����@��.bg<�Z�v�:���`msţ�i�{���^8���*��ʸ��뉭��oi0m�L���d'U�]�ڝD<Jj�+�=��%�_F�$�+%rⳡO;
����v����^s�P6��Βk��=N��/5Q��db��}ɨ7;�j'��אK?G����g55x�v|(��*��mֹr�;쥚�ʝ�gJ����|6xak*-���xs�X�N�aC�B֕;Bsyg^>T'��I�{�r�FCQ�PV��yk�v�ӮYP{
.���Q8�d�F`�i�lj�k1�[n���X�[(��r)7Q s�V�J��{�O�[P�W궞��%�`���Lš6�h\︗�(^�c�ҩ}7{�"$s'0�Mn���)�����d)�p���<��QDp�Nۭ��2�bڔ�t�+]`��j�Ӯr8���-`���4�͓Hٚ��l����5q�2�ދ��X�جQ1�M�qh��٘n��dal�T�֥�
������5`�Kfz�NTb�u�&7�1q��7�Uo.�|�ˏg�C�:8���r����/o�tb\�-4 �	��:�+[U��v�9&x'e{�c>���s/�ОE����\���h�4y��ǥ�j9��K��5���������ݐ;~+�Q_N>k!�LUٙ���XW�fcR�l�XS�m.�oiMv�7���k�,���EtB4�c�f/r�hN=�vQT���qj��̷�k������I:��E��M�X�]S�09p�}u�{q�t&�8��Qn���6���S�4(/g��qP!�����29��\��oJ��E�|�q`%3p��1]�v�b�scn�#W����>=�{s�*���!�E�{�3D�K=t}r⩍�(���rݨ�I�EH)�:�2�鏫0Q]�1�	�J�|x
v��8V[���1�D�c�z:��&�˫�x)vN�n�a�9�+:��]�k��**ux���{��3]*W_���_�5��Z��.̾)�V��Y)R��"���xᘽv9�����+��o!W�=���r�Ʒ���We��X�2��\�$��̬�lm-�_�ڛ���>�k��j�/*<��/�	����.�9��g7;y�b�kS۸M���5N��3uC���6�y߷8|6i֏��ǀ�����9
�P6��z��S��y*��?e<�.�7}����y�V�&}�;��ԩ�_}z���Sn����O�q�ߖ�N�\�hw��m�W,�T�K������>��M����9/���h{^ӓ1�sR���=�t5����|f���ٽ���.�������M�QWT:��y
ƞu�eE��ݦ���MRt��shۍ��eVZMն�1^m7km�����u�j�^1���;��|ii�����\�ޛÄu槼��q���ؖ�4���%5�R�t�>��k�a�X��5j�����N��*�Ȧ�VuBl��k�r�u�QN���-��K�*�1'+D;���ӧ�U!���`ќ.��[SN>Y&�i�
� �y���ݏ���J��n|�7r��:����׫Z��C�������+��S���w��=�>G�o�`�o�Z=�,�����)�z;�����\h�����ȅ�����?_ҕq9�^��F�y�|���ϳp�MJ��}�z��z���B�����~�W�7$(��t��4*
�!xZ>Ʀnp^/z��T���נ��k���E}�J	��������^�Q3���_6HF�����*���Ù�y����%^�ϼ�Gzz����'��<�\=���%ʒ:KEP�sԨç_�,WO�s�ǣ}�ɟ��x��>��qc[�F���+���K�ʏT�o�q/`-F���ួ��qg���h�Ԏ~9*�u�*�J��E�/���q~��'GD?M
~t=�~��TV�|ɽu��y�k}�g���#�2��v���}q��a^z�Mi��]Lxt'b�:�ӹ���p>�Ö�佹���R�{nǆ���1%���;n��̨w�m{��������vp�0��WN�KF���r�;ݐ)]I5k0޸���h��;7r�ա(Ǩ���� ��{��+���B}O�&7+&B)c�Uv_��i
�K�G4wI����-}��Q]9�d��v�P���%I�]]Y�s��n+�rq�vNo�kw�%��¯AEm��7ѣ�mp��]�(����Z���%����2���9/�����}q9�j{���X��(�*5^�.S�pmW�����g<-�<<�P΅���X�VWwW<Qk2�oz��Miw��
�#=6�Xq�灸�V3�޹�=�ꉨ��<b��8=[��﹪��}ly��^��������us�zd_7^d�������#�s�:��O�x���}�o?S��h�
)^H�<������S�L�>����ˣ1�����(z����Zf��^W<5�g}����;�c�ǳj;=;%�鹨@LEw�,r)eTs=5��73�?	N.vթ�^���ߴ�,-������d)�,�D9d}2�%~d9���&'q�����f���Af�����l���#}:+޿_�W2�Q �ٯ�H��Cճ�"��9���M�J�rQ
�����k�ٌ�>ξG~da����-{)���0��]U�s�I���7�ڔ_ީ5艉�w*N�Y�*{�2!u1���b���W3��9�H�jl�1�*�2�Aw�!������Gx���!����N�+����d�հ��ذ��YtV����˗��s;�[v�|���{���^.Ҙ�ؤ���,J�43BIW9�E�J�Xzu�9&T�x,�����(�O]�+�\�ւϝś�	�o� gR-�'㶉���W���������#����>��CY����������}�ZJ���W��$�t�zW��11O�hޗ�ݟQ�F�S<���;�'�7[�C�z�_�C�@yg�ր����M��-�3a��ͨU~���
f�^y�6���ׯQ��j�9vj+���n��	G��G��V�q��7��M��������f��;�W.��w���Kfil�z�o3#��E�\o�i����B9S����^�]B?�����eb�D��W�����Zw����0+yg�<6=��b~S�׼���D��M�׷ë���1�	���-��ڋ��(vzkMƹ}q�l
�[Oď{%�0x�_o�C�Lj�v�s����Go��1����]:�و�,��n�˫x���k���r�j�f9ϰGw�z����󻇝����������{ΐ�~���$�PKvn��λ�y3������Ǻ�m"��^��T[N��{����eƊ��W�����6@�FX�k�DC5��=�zG�=�(*��2�4�tō�,*��$m�i�n=hҬ$���YU.� I�Z�n-u8Q�	�y�:�mv���g*b�n[�z�`E;a�q�4.V\��%��W�)!!��ulyyx)��e<G:�M�c��2C�6C��|�3:��v�r��s�l�j��ʫ��X�9}����H��%����X�+F�[�`�C��2K���4',�Cz�VT7L6J�;�a����.*r��Z5�u��}���E)�-V�����4L��	3X3(V��q���(#�������f��[��ƹ;�s���Ѵ7�F�="�c�y{�#N��4
�H���;� �t��FC/&U�݋�giU���ѹƳ.���d�u"��-�g:"-Ӳv�.�낳�|N �=��t�����]�amj�0T�GC޳�cA��8�-h-�ݎ#�4M<r2�x���՚Z�zkBT�^[	��u����U�б�ab��t@�V6ҹ3�f�t���*|Fm����JX�%�VСNX��ˮKq�����G�����u��j��d��x9̶���:>(�nnX�c��fNڃl�ګp����E֏�Sѹ@���D��(k:b��>�؀��{��W��r�2v�k��[��#GB7)�Ğ��i�]�bm���dLwv����Ů#�-[�K�	�t�{��&�J�r�C��(*��r턹�ʯ�<�_{Hl��`�*[���p��il���Sq�w��:5��̩��2h]4t����γ_Vn��|3M�'g��(�-EB�D��j�N�d��i�F3blrR�v�p��0�q���Pcķ��`�yO���Y��7.>�;wG#z�F�Q�[P�N���V-�N��@�A�3�;���!j��n��ISkO<-��lD��ᝲV ��<Z->_N��(7��	�g��,#hc;���2u`���0�X�Ә���L�ʗD	P0ܥ��&�׽`��W|����0tHܞj����Y*�S�?=��ZU�J"���x 3�R�#H��.����;â"�K>(^�Te��`f��7�%)���ϸ�u�_&v��O`R�bz�!c��tb��jǁ�sGm��N9I�<�h̩ڒ�0
��[�	g�*�F�M7�#�3|.�;̥�ʡ)πF2����p��&�akS8�Rw��p�ȹ>k,���:F��&�G��0�u���Ö�1�e�bu�a��^��E�C�z��F[���
��rս�ҝ�� ![�Yl��@���.�@�{h�cZdk�{u��8Ä�L� �xTGV
)�ٌn�oD�w>���NW�p�I�d�$�O-�"����*�z�x�z�6Q-ŹVnH���c\X�:��A�ۼunN����΅��]pӤ-�orR��f�P�s���� c'ϩ�����ٶ
m�XV�D��У�P+(��+b�+
���V
*�DTU�b�U�Vh�Q��ҤQT+DPF
�W"�J%J�AAc�QT0P4���h�QQEejT�Ҡ��X�J��Q��A���B��k3)12��UdYZ�)���@Y�%Jʂ���R������Q[H��E�d�kI����`e���:H`�"�VE�mA`�R,� �@եci1����
�%G,�Db�b�m�ԊlkR,X�`��Ve�QAI�QUH�X�4��(��SMH�%H�P�&�*���$���R婂�����E%`(*�,D�HT)�����V,XM2�"�AdH"�ԨUf�A[eVc1��c#-� �dF+�r�Ɋ�Lj�V*���(���Ƶ�QW�9^��m�3��JrA�%T�m@v�U�7���XX�jo;�B�6������φ<[�-	�.�Y���9�{�����>�Ys��������x�v=�����}%�d�tק/\{M��gf�ǫ��V���5+�����R=p߭d#>f/=�N{��ߪ�q��E��_��G��u2����|xǺ��ǤWN�Q-�Nk(���_
�����Y�z}�����+^��o#�W�j�ە&:
�, 4}i�§���^�s��&��mf֞S���X/��E}~�"�z��,5=q2�LO�����gn?A������P=ug#SYތ��߮.�o�~;,�S 5�D[�������(z�$o��FD�]�\z�x�8�x�;�>S/M�߅G_���G����~��&���Rnf8gS��/�����'<��ѽ���/k�:�^���R��'b�.�������#��=RK�{³y��{��<&�����7Q���`��O���9�g���Buc��\?9p����b㱾�B�w��[v����z��;R"���d�q͉څ���1_E��M��|��U��S)�����E��)�SG�x�Ҧg䫯�p̮Iu���h�l�j�@�c)jG��Ԟ�[iGl�zm��{�4b� af���2(o�d-6wnup��ܼ��n�]2TU٪j�8�FWbQf	����""9���>�����cVaΖ����tW���c=�Z/�'��Ó���W�U��O��_�k�y��骸S��Fs@�S'��:�>U���ߝ���g�~zѥ��kF��ss蜣��6i��|��Ў��n�9w�į�Ӭ�{�������S��$��q.p�[�U�ZY4��k���¯&uL\Dꠜ�W���s��9����q��\<��(�lk��Y�D��������?BT?�j�|��qo���K=�]<��O;��ϙџG�����+�w����%��w��9+zv��퉔H�;T���G���^������2��h���y%���~�"���w{F�1�g[��T�����6C��x��P��t��¼^�낏�����n�}#8w>�N�U���D�.�P:#޿_�B����Cr ��EzhQn�*)j��<�uf�����v�~�<�f�Q���H���C�3�{�tW��z1̹>���7���hT�w����&���א��g0=�1u{���E(�u�>��Q���iw��"�yT�VQ̟Z���f�='��]/�31���01���s����S|ު��������:0��ي�z�4�1�����|ߵ�[�|�m��xe���z�s��2�'w�8����'n��pT��N`CYalvye�,�\�fH�ޚ��:=��Ϲ�o:�rS%�Ƚ"�7�oR7Ro���1��t�:!zo柯�瞧����/�7��hܽ��aU`�Yټ5{�WE����I�7���ۈ��}y^&&)��:φ�B4��ud��W�3F�:Z�Md��m��|�X��]*N ��\��e�>Go麇�;�g�����r����h��(����n���teeW675"�{���|��zۺ��Zl�y%%��h/�P�#6�Ÿ��}�;�A�����dϾ��6��~�E�s�����]T{a����%�ai��c3a@f�`V�.s�g�z�Z�N�z=�7et�}j����|Q*����������;�Mh��ԕu�9W��c��He��Zz�|+M둾���`u�jy�o=X��{ռo��CW.�����+�]gQ�=Nh��/��JES_d֖0���t�W�ƨ�>�"���;7���y���ۉ�^�gv��=���X)�/	늨~5�鋌����ۨO �;1��o�Q�d���u�:�IM���%M�exu�:�CF{�)��%I%&a�;��S.;jc�]��v v�Fi67@V����'1�TW;M��x��ǥE�ȏc��t'�l�*[�d`���:��⃅�d�5�z���#fIֻb�s���0��s~}�l������0fgA;݅d;�f��'��ؒ�:�r�]L%�NJOw,��h������^���Wg����sj���T����΁ޛ����n�M�mv�B�ǖ����	�W�>�-\Cڱ(�7�q�����H�\r7���z���eK/�}�^<���F��T�z�z��n�"��Qr�M�KgrQ	�ߩ#k�����~�P�cv�wj�W9��}��^����z�&���x�;��x��ح
�U�(g�ԋ�7~�*�٢��pWd�q�sʺ|/DgfAԍ�w�&��LM>�i�%��ϑ�=�Kg���l�,=�(����_S�>�S��^G��@{#r�[�@�L�z�dƾ�	��մoK���=���=��.��Z>�{´_�k��>�=�V���a�)�Q$�,�3a��͢[]6a'���I���aT{��ʄ�z9�͛��@yu�q�gjI������Dς����|"���^��K�?G��u�:���/I����Owc����a�f��1s6kׇ6��"��i�>��J���5��O����a�f֏_�:+N����`r�\xt/W<@���J��>��E$6�˫���m�d���i�P㜞��I�SH�t�^��w����'7��X6�k(�����a�巌�K�$+mM���hjP�N�"��bH4zI�o��j��L=�����X{d�;7��N��Jɺ��K���-X�S�5�+��kB�~�����=�"����y�~˷���|�����Ӝu߳��3u��+:���NX�r�4o��X'tܗ��"����w���s���'����۷6�]�(;��=�˩�Ӟ=���_�Z2>��H^d�v�e�=7�=������z4�l�T�^HL7�;=:)�S1��O��9�OŮ��q�n=�wᜤ���H��a�آ�W��F٣�;jgg׽�0<���L�2]?U����zsޟx�w�>�p�����,�ay�c���0L>�GwR��O�8M�EW5=�I��Pl��n�z�;�����:2=V����;���jc�jq����g$AN*��ZaZ�tj��*�F���&�����篅?:`_����5Ә�K��k/2�fκ1�g���w�+=7 nz	��ʓW�a��{Pz�Y�9��=��U�'Z[�F��U��;��R�����~�d�r�G�R�d�E��P_W��7�xҺ8�t��<�=5���l��wq��~#�<
Q�^�z荷T�I%����,{�ؗ�*<kx��AgM��1�h�:�Z%��I<�䰴���.V���x�,K���^�.7KՋ��m�M�e��C�6Yi���b�6n6����3��G%vqs�6R��_;5f���9�������C�h�F�jN�K&�|ĚcZ6mr�^#���w#L��q߉xi�
�_���sg���N�O��w�D����J+4z`��$��wGC�G�Y�D�`w��W+L��5���@R��v*2���#�*%ΏH�W���OO��N�x\�n[����'ћ>'�rO�뛨򸌭��'äֹ�f�Y�Ǚ�|9z�����f43z=��o+<�7�x=��ՠ�X%a�/�O�:���a�^/�w���1� ]dR���{�^[��(Þ���QjNw��{.�ߘ�s��������mx�I���5(���tUG�KW��F��y� 3�n�J�e�,�������_�$��X��)b����2�%F �~�^�M�����z���>��d�#=:�v����yq�/�9-��~�c���(%�%�1�Z������<?�֖r��A9����߯��{�<W�w���F�Z
w"�T��]׳W�>�8O����=uL	���b�v�_�6�y��g�:2�y��е~Y��,�Ia7�k��z}�j�s�l��϶&Q���7T���y�7)��?>G��,�����g�F�Iw�[j�I6O�Q��+}���g w�S���G] }���6���Z|y"̂����j޷mܭ�1����u�άj���P9-��9uՠ��i�!�Y�hV��(]�:٥����׷y�A��(&�R�dĝp�ɉٰ&�'�"�=��Q-ϟ�`u��A�����Ϝ�S_�w���"p/��ʞ�� �֍�;�_k�G������H�c���ȍv����~��2�܁�7;^�U��0=��6�uD�ow���G���q��E�U�:��sސ�g#}����E��U�/ �gm������n>�Z/9���j�z_�@aa��u?�������/�F��^z���^���B���o#�z�^���$c;蘘��-Y�t�9co��l,�U+��m?L����Rn�v�X^�)��.���|�)�rR������iS�<f}�}ǱcW:�t?3�/��3�� ��^쥸��S�Ҋ�;<8�T�9�(Dϑۉ��ו�ag�������2$]pb���;ܳ�N�1q�UK7��<��;v<3�s����蒎\L��㹻P⽎v��GN�uf�]o��/e�A��&n6���y����O�)To���q/�����L���7�Es�6��z���ʴ;������=����~���8��q�_TV����_Dj}.p��Ti�Y�QW/�~�<�%��&����X���M*�u�܇R�0���ϔ=�W���ы xя7�t	frL+��ռ�K@�cŉX��8v���-CyW�t�9�:�n᮰���%�C7#�,�9��[���/I,�hK�㓍'u���1Yt����p��W�����\���Z�xeg�����<�78�׽~F��z%�ٟ���g��{_ *���F/�wM�x|�*��ɭ,a;�q��5�ٮ��G{�'�C�ʑ�^˵������<�y���Q��R=%��P�j#��:ϲ"���S+��A��|<p��|��_�nU�;���3��χ��1=`��$OMIa�����w��vz���{}�U���pu�7�Wp�ϧ�WȎ>�i���Rؿ_���X��S�Y�r�3�w��9��2|������9��2y��hj7�\yz[/|���w�}įO��,��sAj��>���M���$� ܁�q]t* ��'g>�C�|)�Sfz&w���7����6�K��}xcUU��FP�RP(eLL%Qu�h�f�G�亘y���V��E�1��s�9�������T��P�6�,o��%�W�K�B~�n$(���%�s詏 �~J�-���eH7n���X����M3�s��Y�_ �=�[�@��G�&@|j�&'�}[GVy��~��	2d�U�ՈxV���fI�2��T��9����BFRqi����	f��4q�����f��-ӧl:��}���83w������@ة��}Jv�x���k�ϯH�/.�Xi�oE�>�����x���_�0k���S^7�T��s�!�Q=>o�3a����Sp+�z���Wu��������֞Ҩ�%/�t&3~��6_���.r�<�L����s�?��V.}�_�U�E��mhXu��eD.��By�U��y���:���j܀������9�9yşOG����$�������N����7��3W����_�<2�� H��
����;�� �nWW�͝�Ѿ}�*�_�l鋎B{I90ﲽŋ�٭:��ζ=���{����p�ν�M!��=˩�s�/GdG���_c��r�l��?r���W�/��؝nz�Hl,ޝ����Ѝ��z�M������#�-Z)�Q͉�0���P��;-dѹ��9鮬���~��y��2�y���~�q��K�]�ˎ�p����'QY J�<7(�j�����=����L	�w�W��C�����[�W��6V�ei�*�q�q��=q�p�گnߕ��s���OH�*��T�����7n�{�ԇ�3�to�������]�Q�G�v��f��SK�-��"��A�̾�d�f���y,3G�i-�.)JvNJdt#�9
�f�Pyc#�s������ �'+��,c�;V��r�W9��a��V-h՝Ü�����jMUP�y��Ǚ|/�'��%�bq�����*Y���0&-h��Y�.�g�gѵn��3��%�@�U�5Kea^s���T�}�XŽ�.���z}Or���_��e>=�
@ɇ��C��G�!��{T���X@h����=���yU;]�e����p��G>���/#}`h����@���� y�lL�٫SC+W�ϱ�ǮwK�^�}�>G�DǼj=�*�;Y�9}H��Z w�DLS�r���,>/o���_^V[Ѹ��c[�'�Þ��2��7�Q����>�g�re ��{l��.s��b�U���]�$����ۥ��̏8�
<��۬<�7|é���Kޱ*Ds���Y�w������m�w:>ў�n������|Q���s����5�t�]lz�N��
9C�]��sٻ{z�\�q����^ڱ�gjA��$>9���;���J�����]�X�[�[*�{���<X���UO����C��{ۘ,dC�8+�'N\�gnv�ῳ�P���Ȝ�AFH����pc}V}�q|zs� -W���#ޝe������A���,0=g�����}�ꟿ5.c��N���e��:	�0��fs�&P΄�"��Kp�ö�#���Ӕ�]�H��0etyl�y��e��Z�����\3J}Y	�3kh@�0�%�B�!�7�	�|��O�9�m���ss�`s��[���r��i
�>��c���+�f@�g�� �Mv��� �A���kS;�-�,ee��)h��F�+9d_i�]j%�(�&�x�4D���'��������Es��.��o#��5i�Ҷ:�c��98�Ժu�������ͬ�of5/�S��!�VM s
]��)�v�CnS���E�Y{p���3����N�l�=+�/5�U��R��lrܮ���u�׷#J�g��E^gZ��kN4�-V�nG��;g��Ţ$��v������M��� �X��*DϹ^`T(&�:��W��vE�5�T�"j	���\�m�wE�E���O��qc�,�v�ό�9T^���ZE+��#��m�����eR=wS4�爎KD�j7*Л�1�V^s@W
u���;�\I��.��K�fN�6�m FD:��"ָxu#o���]�T�<ݮłu���$�J����SA�}�J�+��ɘ���p莀
V؏��p�T���Q<"×[ґ�x�=r�3o����En;�x��M�a�I�z��ϖ����$�v��z�0�i��W(g\c+3FR���,�	0��|U�@ѩ��G�m*���Og`٣{{��d�@Zu.6z�䑝i7��[�M�D�%چp���M��U��L��8��MM���R�#��>/iM��ؔG��QT�|ܒ�5�q:`6���L�Ҭ�|���`����Y`�]雐�5���ٹl:��79����ԣfwS���*y�L�if�Y�n�T��^g�S�t�b�uu�v
��K�C-� �5�^��Ы�0C8-��Ia�ݭ\x�fj16������ ��v��b̀�sv�S�ljz�|ѧq={ż��o#W���c��9�DmK����n`r�#��,`ce��lfy)c�RҺ��7X�#�M_8�ꓭ�٘�R�7�ԕ|$�:b��Z���{oC��ـR��rc����@=��cf9�@)]� cQPAW����UŤVedѪ���X[����,ݬSx��e?�<�N�/7��,;ub�	1�i	�ʻ���w�8�����mWh�|{u#֛�	}a�B�n����g���ji�z7����/�(WN
�w��]�f�Ռ"�o��\$5�b��;taw�ٷЈ�vb��v_*���]�ox�NOT�1lQ�u���\m�V���,�7VU�s6��2&NG٫��kէ~������¨'J:Mي�re���1�P�}8�Bۏ�f+�֯�����$�)"~'�*MZ"-J��dE
�dUS-��,̷,Ƣ2�a�
��0�I12ٌ���X��[k��U��+#mVLe\�+%aX��b�Y ����U�@����b�P��h�h�Aeum@�E�咳�c%t±`j�Y*���&�PąEk
��TTE��(()&0��&5%eb�J���J�J�Ad�WT�BTr��XV[V�*�2¢�1`������Wd�B�`5���ŕ�!1W)P�1�01�q�Xel[h)
�-�X
TaR([L`�Q"�V��2�H��
QV(�U 8���2�PU1��VH��Y*,
�*E�EA�DAF$Ʋ"ȫ��*+	G-1
��*E�E ,���G�����r�G�#��t�]�%���g��XSP<��
+z�q`=����Sҡ�I��[Q�qވ�t.�"�[>m2�R�c��o��*ۅy-\ޗ|m���ޯ��\�]�\s7	���eO?,�V詚U����n|D��8���U5��d��b�']��C:����{�qד�k��F�t�Ͻ�]�ь�Q}ܪj�/Gz9m�JG�Ӏ��0&"�X�����W�tG:��ϙ��Q��.=�W���\�k�����7�c��*>0�쉞5'̩�`eO#�o
e�۸~��މ��"M�Ѹ�,��Z�w��=�ף#\KG���ne �V]F�˂x��CM�'��=��[L�Ϥf.�ۆ�u�B{�o��{���E}�_����Pn@���]g·�玾�$�o��^C���7��^�낍CĮ*�׭#��2��D误��E��W��2Q���N��Q;�`T��`�V�FO��,7к���[��JV�@�'���2�����a�8��0�|�h�=y]%�q%#�10�WH��=�x�9Ќ��߭��^�j|��*����^�mR��N�������ʓ`/}{�jW��n$�v��d��ئ�h�k��i�2���^^@t�K���y.��T���'CY9���뱪���H��������!ã���9\U�j���Gm��Q�O��U>�΁g�*U�[$�Q��/��lE�e"�i��s����B�6�.7&J��n=�ֱ�������)�;獌���Ć"#&�6�V5hN�yi'��4����N�ʀtU�CN�+̔<ӫ���Nǜ���A�4����#��nV酞��u����F8� W��z��S���W��5U>7΀����xg�p��Q˙c��ͅ�~�j��-��N;��W����}{q��o2�2!z��'>�T5���G�\��IGű��c��K�l�p��XG�3	E��:Я읭��>霒�lv�\{=:�&��4�{��*|�5���*��y�]ϴ\�GЎ��7.P۝���Ү2|+Mƹ��`u�y�sӌ�D�K6�|�����UӚ�`➊�d����}�<b�	�7'�|�X�3��'<WӮ�אײ�m�U,ś��\�m����f�R��\�U�_�[e��)�K�z���㊥����}~�.����Tx��z*�o5z��޻����������W�\:�Ch�{�(- �ߤ��nj��=1��/���}�c��Ѿ�ϲ:��Ŀu�<]{
������c��R�S�Yx�	H�d'���b����v={��d =M߁��^.��bQ�o������������SyʛOhƙ�Xzt@[3A���]�v
뷻��*Ν����}�&��TS1~�zp7S����aX�����	�)����!Pǥ������7��c��"��b	��ׅ���R�40��`|䠤H�`|��kӠuG:��=9���=��u[�V�f�ӧ�� w��-��Ш��p��q��	�j���a��G_#�bN���WNt�����Gv�F�K���`�]�L7WJ�A+�a�.W�>�������z]y��9^���(y��NDo�w��"��3p��\LL/T]"b�O��-�X0WQ�[���<�_<�+a}>ur|�(��^��#�p@���|�2���dƢ�&=�� �P�w��O��<W�
�鿓����r�Z W�l�y�M��-����p�6�@^�f�:ш֧�^�莫u�t{O��%/��v*6�y��H�D7U���n��RqB�<�U��+7�q�˪�I2�g��7r¼��������4��.�<��ǹz����:<s;�߉�'��0���!�{���N�x�9|Ν���N����#\�z6�����&}���0�:��RyZW���f{�G<����B��R~�l�gב������X/�w����jnC���bU�@�7V���B�SD�h���B�ƽ5��X't��^,�����M�N�~~��ܥ�a�U4�YB���Q���X�FGоZ��O��s����-<yf��v��/�(ͩ�g6聥�]���ϙA6mnj�H^�+�F�S	��]�V�wf�v]u��6
�R�dS)K�Oy%������2�ٍQ��j�9���^��������0JKzg�EAx)u^�e�o-#��/]ǯ&w�p��TO;��O��9��c�q�W�֎���(����ڕ��q��U�BZ�o����+�CQ�)φ|����B�U�h�S����>�O�T�[Ԫ�k2gܳ��z:��"��%���qT�����7(6m�ԏy���F|΃wz_j���.H++М�۞���g�)��U��Юe���pz@�3�9�Q7���!����o�i���z�(:�!|��v���/_�s�Selt�z�Q��g���!������*1_�Xk�O�2-,�Nk�Ϲ>>Xy�G:����n�I���/>�X/��F��zn�:H���2|���^([~Թy�Aݧ�>%���5�y���W[�Ϗ���������Qꜩ;}z�9���clekF��M����"b�=�`{�0�UO�s�^�.s��T܀����K���֫�P�̟I�9�t�\Fz�u���#Y�्�N��[u�s�3���y[�s�ٟv��B��f�D�è�s������ۓሦ�b-�I"�3�̮�9��@��❺[t�������}.����y�C�<�Ʋդ`Yr�+�Ojd
K���y)q��Ӓ�t�c��܏�.�#y��t��zM9�pXꛇc�׬�`v3yA}l�����-F�ܜ�7W���v�y�%?�\���7RMyωZr$���������2|:MDk�j!u���J}8�6D�N���sN��/}���G�\6F9^ɡ�2d��V�����/\en�w�^��������<�X=@ϼ���þ^�-I���@u{ț���b�?`��pgא��ٟ��'�޾ef�e�{K=���ϳ��+c���֤�?T5�բ״V��Y'N̋o�n���oR������(e�m�\FO���`o�ڟ]��+=:�v��\r7x�+��8K>������Z6O��$<>���*�u�Z]���b�ؗ=�#9�_���[�h���=U#{+��=܅zl��]����j�%"Y�{~�`O�=���οNEm�'��~w�D�>\w�V����c��T��\���ի����ό-�Q#�zUSjyaL���;>�;�W&�����7�{�����Ͻ��}Lr�m�TmS�wC���t���0<9��ޭ�K�VO;+ȟ}���낍<�\{>����O���}@h�����r�/�m�dQ������Uu�����'&E�e��@�"7.W�3���(�c�&z�n�벳��R	�J=��8���j���o���M�{�]v6�&��e�k�Zuۭ�A�7�vI���0q��N2b��Wm�e<�}�**{ň]Q�P���xQow�K�Z:e^Q��c�Μ��� �~�z�g����>���Į*�/cgb�L���8&�=�)tR��]B�_og���Y��=�@�9����T+�����ә��ߵ���W[�Ϗ�x�{��X��.��J"�iޮ���{VY�T��rO���baz��3�9�}+N�b�7�CݱN��f(3��d�{���oLz6W[�Ϥ�y�w^���Il驇��W���j��ƹ���92㝜�zjF�ު3��9��'VN���U����N�@����"��is>Gnn���en�\�2|01�yѱ�m�'�=���Y��C�>uR�����:_f�#�IG.e������5g�f�y�^����{���oj�׸���E���̿���9޸j=컏d3�8f손�n�|�ќ7����~�+�RŢ�����X�O��~԰06���=��e}��w�����{��gz+���M��n'҆�Ӵ�a�+���7��鿳��ֹ�}h��-��x�$+��:|sҊ��o��qW�۞0�ñ^,��2�kK3�'\��VD���ª����΍ڏD������ց�&�ք�^*���L�'!���W%ژ1�*"3;�����ϙ���N��
�bT�uga�t�U�[[�t�%he��ΡUs�b�D���;
�4����R$[HL�.y�zx>1-��r����Ϸ����H���=�tu}�;C�<��1q�%"C�{b��F+�+)!M��I$$��Y��s�=��z�S�����9�{�y�exu��CG��P�(Ԗ��g*�Y���WzP��(�0=��\d�[�~*"_�Ǹz}�<y��`.*b�OQg�'��\/#/=����|��<��&"����d�]��^
f_�G�@��n1���9�}�ѝ{�*:���6����g%`�X�D�*��GdW^��D�d��wQ
�+�V߭��x-�.�,���f�ͬtc|���r4�Z�p���E�0[=LL7WJ�A+�a�.W�c��f��I���x�=ԸN��,���S�����7�U�˂+��3p�h����&&�W���`�Փ�0f����+���1(/?Se�*��N�d{��9��<���%�;) =���؍�H���>��}�z�>�Ox�dP��~��Mx���z��H �=�6E}=R����}��V�����=�/�l`W�Du[��Z^�Q�J_�;|�f��?:�佻�p��>��P��J�lM9I	��¡F��SôO�Jmh��������>2��ގ�ZC�����a�ܰ�d&^7���D�o�N��db�q��K//���]ݕ��J9ļ�3�lĦ-��跸եZ�ѫ��l��'��pς�q7,+ͭ�'|f����3��w��d{���L(�vT�����MC17�cS�[�g�C�]��Tp�~>e�ȓ�v�k���N���c\�j����$�̕���wwy�h�:����kݕb�=�.;�{M�h���Cˌ�qb�6kNL��El���N#�Z��&��_q�~�2=��7{��DJ�CF|�kE��nK��P��3��d�yz=2oe��}�t�,�g��Y�����Y�ϵ��Nx߶w�^�
��<�8g���D	�5O�{�1��:�lMy�C
�;ю�=y3�N��U�N}~��~/���i�k��:��j[�ټ�]���p#��
��x0z�ި{�)φC�㊽V=��=9��ţ�+�D�O�h��?��o���c�}�a��s#���Q���;�T���^��(6^�������z�9�х\���䗯N�wGz}��z�Юe�|�]���g�@l�lw�̊܋�}W~����2�yW����6��v�w�R=��k޿dz�D�� 7 `ng��G��Tiw��;+ؼ�dq��>S���0-`^��ʾ)CJ�nҫ�+y�S-��������Z��GB�q�Z"U��0S<ƺ.1~<Gn��9e8oE���\��q�� �(�ʖ�IAK��pU\�	�g��v�	���6K/3H�2��X�r��k���c ..�&������ש#��u ^��F�����O�C�yK��>�||k���x*�1qx�����J}gIc2�C�׮*�]o�{'�K޽ ;�e�w^�8'ʲqn�Pp�d_w�9��lܟD·�����DM9�;��҉xz9���yUxߋg�Y��O��-p볼��EW�~�-�M,�%�1�v�鎿��C���ߵ���,m�v.3�V��x���p�Y��l��G�7����s���ԓQ�>%i#�驇�9����Q�t��-�%��w�-z�g{G-�'������� ����gjA��$1y�P���a��'��Z��[�g���3Q{h �z�9z��';�:���N����o�t�K�r��y�&mӷ�{~�g���6g�i��M�[ Tb�~'=��Q��̉�~Ω���ы���}2H7E{8�F�d��f/�D�W9P�����@3qc+�2k�S��}�o��EQș��n�W���T�+ћ�q�WZ#0��X;���i��������z�n|߯����lT�qyx�\o$a�g�)�R!�$mXǳ:��3:�3D�xj�mnA{6u+��ʔw�Y���^��p�N�;���{A���������0��J	h��T<sW
��k�j�<����c�^�3��_f�r�]p�ƍ�1�j���lq<�[��_����7��#�=���%"Y�{b*�s�,a:�*+n�y9�!t���d�N�;��X�?S���|�8�W�ګW��g�}�2�EN�Sb���/�z!j��Y"�y�
���s���������FF�%����e��}aw�%���gn������!�׼����2n0����_>�,�l���Aܯ���%��ldGNQG�G��k�n��6����Qp�L����:@�KGۏ�
4�+�s�H�zB)���N�Lu�/��!7UYMW.7�k�J��ͧ%��$�a��T>F��2����kؕ�Zv��J�ϧ�f��[�Ug���œ���Ĳ�+�~�"]S��l�LL/���&��Ҵ�B2���fG��`��Z�0�ʧ1�/i�g=S����x�#�ϩqȣ�l���&�?s�ON������^_�^��]��M��ޫ'��������9�=~7x����jg�U��>^���-@w����w{<�v����I�+K�j�8\Bv+��꥗� {������8h�^�(��@TT����~���.����9�({6�`� ���AjLD�V;2���;��u4�g4�j
�tU���u$��?K��w��z�@�uV�%��w9��I��(��a��{�T����yƒ�.���u&�o�]�N��ٸ�T�#9�]��fq-RCfVf�H`9Ŋ�D�c+����6����D���K�Q��[Q�[vh�pь��1]�NK���5�����p���Z��˥�LZӰ�D�ke�Z,w��h2��a�G|�`.�J޷hÒp˳F�X)TEfRjr
�5v޷����Ë�]���\��O[G%�5\OT{Y�_ub͛��ʼ%�ҧ�Z�A|���2p+�+͕��]�֩�9���d�g��s�w0p�}�l���o
e�ߵ%�2<��JQ!��L��q&7l��R��C׶k+�i��t!"�3a�Df	�bY�˥"���A�8I7���zk���1���"�S�i�<�z�ol��s3�4�_m�7�Y����20�t�we��B�ǂ����y��+
����W�%�}��3B�Ӕ��T��X��!ֈ��������fU�A��}����(*�����rj�{��vcN�I���n]��ZS㯲��/%_O�!�5P��ZZ�;wH6��Tj\ ���3�	7���h���8�uWg�-� ��$�eaU%�\��a� ��'Yv�5��A��VA�n+`���k�a̕ˡ
.]���t��dGv�ڹ��7��*\�"�mV[�F�v9e���ڊ���T���QW+�{�&�a���*��Py���U�Rݗ4��E����GS}�ζ	��V_|�G������������9��(2 *���*�G	"c�ИKM�*k�<b�8*�j���z���rwȠ1|�
�v}�qq`m��" �]�a�������VAܬ�]x�s2�~i�j��;�Zn��11�e�Y��y{��<�+Ku�BD5R�SrS{{�֫��`�Z{�bA�wSkfm��*ȸ�2�j�Z���ɗ,\Y����S�(+�h�`����۳!6�ɩ=ك&uf��j)X�pDnj�،(]����[��V�_E7�Bĩ�� �L���!��tLW�yÝ�;��Ʊ��P�b��S�X�@��J 0���V�К-��9�v��㰆����YFiN;t�Yٝ�7�u-=&R@Z�OlC)��VG�%$Ѐ��u��&p��Ui�V4g�>����bYn�2�* �nT�����j�sՀ�z�*���ICvnq[�r��ȸ���ެ�����D��R�kpÙ��,)T$K?'�tuJ�h�|���!�헖����f�{K�y\+�L4q�r��ޡ΂�a3�iV��Ң:VC'v`��D���X�Un��,��܄��Ƶ��s�to'urwH�$p��=*�V�tʽ�sY�ұ�n�b������$����w�i�q�4����4�דk������> �
*��-,c �
E�� ��,D�Y"ʆ2\�(,�U"ŋ�@�VV@EE\q���*��+k+�QjVD�J����DJ�,X�� ��P1�DaR���LH,!Z�(V�E�,�j�1̡��J�IU�T���!X)Q�*�1��
 ����V��# �Z9B���
����TĪō�V ���EFEU�B�IR��f"2"�`�DR
1X�dU�VJ�D1*ATX
)��ƭ��X,E3,1�FcP�TXV�j����%�E�b�d1�ID�`�*�b���*�Y+���,�p�L`9I[JCC~�ܦ�t�ǘ�1ۍ�Y�4��g.��f꾬�6Yy��`���;-U35wyy�p�FœsD�X^�2�����ڲ���Z_�7�����Oz���ۇ��_��ު�s�5��{ۙ�����_��uG_{��=$����=7��_������,{�o��`V+�G�ޭez+,Iɵ�ek59���dk}��;����p��N��l};Le�֕v��Vy����2�W����R5^����{A��޾e�ը�G%Qׯnx�G�u�~�<>�,�u�بӧ=u&��R��_���;#}^�"��:�ז����z���28QJ��@C[��FU�
qF��f})f�Uw����ޙ�}��2)��1��KK�:�=�����%��ם|ie��;J�_���*J"�_!�/Q�Z�uϢ&�5�q��%2���?��q��a[�L��_�Å��l4���4�r={��1R������xStXM߁��˸{V%�~y�/Sf��H�\r��|ƟdǮ0}ig%G�gѻy��ϋ�E�����ar�8X�8�Q
�+�W�eWMo�ߤFe��R3�w�z��Ǜ�R�Ϸ�4�_��<������ut��A+�a�;!� ?���܆^*Xrj>�<]+�F�㧳w:�[j�%�=�U�ɓC����[jͭ� K����ƷNh<�6�ܵۂ���壪�[:���9:Ѹ����M��ʔf��fl*i���p#*r�\��NJژ+�MP��{���� ���X�w�|�®+L��(���g� ����B��Z:`����&/��ɟ2W�=9#��瘽h�	���B5��z[<==5���Ӵ�Y�_ �=�U��L�{�	�p^����eA�����Šc�Ru�ty��
��O�p{�5��U ׾3�^�G��
���v[�y���ۺ��>�C�flp��!۝�x^�Q_"��'b��s��7��<�Ec��׾�����q���3�$��r�z���r¼���3k�ke�3+���2=3S����w��ǖ��Gf=��G�ǹ�d{E�a��2��3�����'t����Zo\�aќ޳J-we��{���?b�c�0W��j=�V*߶Θ���Ih���Cˌ�qa<��T�OޫǗ3W������δBڿzHϽ���Ak�Z-`��q%��O��H��l���'U�:�S>�����]f�U�Ϛ�Y�φ�_������^�z<�R~̣���~+6��K�}2�7G�V+�����Nʞwq����r#�/�vǲ������s`S6���VuL%�:�&��B�N�ʼ�vt�hE�֞����t�2��z~\����Wv�ǻ�y
���h���� r^*4q�t�w�Ƈ��n�)w(��u\i�w;8�u�Z�����^`gita8#Kw_U�-I�\[�"��X�"��t��q��l�(�Ԭ���G�dl�*�ς���1}�{�Iφ�K����|;�cPn��5j{����/��{b|,�>��R7��Q���,���%���qT����w%��۩�ۚ�w=u��9o-��
L��
{O����\ת=�T��C�th����B���&{_�v�xd_MuM���iGۦߣ�����ւ��鋃���=�H���0�5���dmy�i^���Z��c��xs�%��}PS��4�RG=�Ϸ���[��^��W�9^]��v} ��#q�k� &k�sB�����%����C����d_�W��)�W�� n/��F(Y���i�]�����&�g��s�U�"~�=�r~;���q�Tw���Q@)�ܭf�F�Vh��Gw���x�*n@^�=�M<�J�D�4v�n������.V��|6c2����j�fQ�}�U�����F/[91�?z���Ǻ�.��gļ7��qW��CW���O�I3�v]t��ݹ����G�j�o������ߝ�p��c��Ԃ*<�����������c?y��?	�؇�q���;��Xem���T�wm��oJ
�N�<mH��8Kf.�z���~�o�O$h��E��3��0��:�i˭�Tznp��r�7��s�w��{0��SSB"p��#�F�yѮ��G�)�x"ivfe(Z4�OVw3�S�~������� l%~���T|��%�_��b��>���t�gw��ʝ� L��|��`�}xs�K���T+ͪ�z}��y���+w�}��_y�5�����������F&�ü�����ȗ�)b��ۅy>W7�����ү^���N2��z^��>�U1ʱJiY�M�O{Edz�i�h��������է�ҭ,��|��w��ɋ����xڥ?���'rg�m2����Req��N��w�[e�8JD�`���{ŋ�&u�EpH;fs�W	���<��;�>��q�>gC��|��������q���X�{(��}�L����ɧ�˃x��u�e��ϯ�w��u�|{Ձo�Z=�?W�\:�A�����!ԣ\�Ǐ}�n�(���K=�V�&�����q�x�}PQ_<�\{ ?Sg7�W�[�V��z�'�m�U���b�O;d��i�����ޚ'��M
�� ov�>��F�%qE��+���#��	\�썡z�o'�Wwz�zǾݷr.9U:/>�n&��T*�#��,-8�_���q^}��'�\ 6��3&�o�ć��+!����Lgib֧f���礈�-�� d�b�g�i�\�͍2���<i!��f����KƯ����ju�m����C*�T3���zwS7��@��C�킅�yq�nm�M�����5P�8
���b�m��S"���]�7��S�%��?P���n�SʧE�Z=s���&b������V�������g�{|�{����z�+��zb༯zg#�8�{rD<�ID��͛�}y^&+�y�C�Q���Fvn���}�<;���N���k��H�O�����ːEB�� ng��,S�ʇ{���-:�����='���W��|�a�zf|W���\9˱ᐧMw�R�,o�|��ѻ�˺'#�K%���\}�Q�����/����~-�ׂ��G��;��ՍLq���4��6m�+9���s6}�zJ9q2��q;,e�p;ɞ;��t���,
���=1�j|���'ct�w7uu)�(�}�H�[�Q��T�؄|Oi��҆��1�5�a�;�k���aw�a��Fe+>��;q)��W�X���k<{ռ|�TW}�nxŬ�C�*���1�[�[G����/�s�&�Ͼ�]`w���|��W��S�S����*(�E�)����&;�G���&���\[:�P�L�s��P��z���~��ǹב���^��	����?�x#�kz2�~��טd�8%��}��w�y�%�;�#�.���O�W�nuo���,	a�ۧR�ۙm$���l�6��{���CeE��BbTS1�5�3,Y�w����;��u���.<^M �>��}��/�h=�
�7���B��1~GF~R��b+�p�2S.�]���O�"�{��9�}���a��&��b��s��u�rD��p���΁ޙ	n�
�L�{V%��+�B��z�Q�'5��vw <�8�����7+���^VT��#��� 2���Ǚ����v>�r�6����$��W��g�c~+�v<F�߳�E˓�-sکJ�XCpv�O,�������e�:���]�W�e�{�9��5�{2���3p��\D���j<Sd��O�C��W����<�~��T{ԑ�>S^*=+m�� z��PFӯ�r�����k�KDn�PZ��򣞉�5��&&�մoO�{�L<<��h���_�z]��O��S���}ېW��Q�C�{���O����ٛu��
�ղkK��7	u4r	����͑�˯1Jfco�3׹��B��o}��2��Wpϋ�����n&�q�Z�N��F��d�.�=,���Q�S�����i�F��T}1o�7��ǲ>g*p�����$��~�螻�~X�XT&��L�k̿�Z�㘦���4v��*N�m���㮋��30A����\�^� �`�П�������7ֳF�.�TyP���ed��J���9�Hf6�A������tP-�'8�eIm��ؗgwRb���|���͹�5z�����$�cV�XM��yS�m�7�(��}�h
�cǱᾞw��z�5�ʱW���t�x�C�&��Dͥ�+[5���^)^>vp{��޹U���)m[���l�%G�h�+�(w��֋X't��_�<�Q���o��ׇW���������@�����~�q�u�)wθ*�v�v1�����V��=�|v�xa鸢ìWp�fg��|7<��r#���s�/�tӢۏffn�ȗ����8{o�G���+#dID���`L_z��d�s�����U���+�w�w����v��W�ϼ�2���z�Jc69�,��Q���qL
<�&��2O��1�<� ���h#G�-�N��}^���y�z=]�>��}�����ՅQf:�K�4��b��Gg�Ϲ�d��跸�Z�K(�;�ŴGzz�P��Gz%#پ�6����Vzn|no��3s���Wy�N�x^4}b�gdǋu� 4}k�}pUC{����Sg>���3����j�m���󋐏�o���/v} c��L��FF��8KGu	��=��*��W[���\$�fi���y��t&V7zj�=_ ��߫H��xtf{�{���䣼�[�r餵q��/wQ�9�})Z��ڠ�gia���+�x�Bu��o7.k�[t�����5D��}��q��+>��"w�%�ǫ�9�*�y�Mp�&>�rKod�&�Ve��䏨 �	e�]�N��|���Ǫ-QN{N��wJ%��|�.�Ƹ���G�+�}>��n�9�f��R~�$����o�0�ۉ�c��C�ZdWѮwǋZn�*%le����n��?>�f�Bv*2߫��/��C�K8=�C7RO��+D�#�7P��[��W�.0�绣"�}܈�1�m��g�ux:�������##|�r�{&���QO��ܗ�M�2�S��q�7�c�Ks���z��W��7��f����+��b�Qi��u�������}��'��a�*uɟ��^<�~�{QK�k�� ����q����׉Q㬳p��B**}X�S����gZ"��{�kE��'N�L��7;,e���=*�Di`o����]��7ӳn$���OdUV���N��|�6��ͭ������,�5��b����kK���L\N�	�D����$z�\VEy���}B�.����_������{~YE��f���Sb�X������<ۡqMy�0��s�t����vi�8�3��#p�����G�; �*O�R3��{2Q�;tzd}���íMӾ�C|�.�KT���+R�m���b�w��;W�[Ns	���Ѝ�4�I��Y3��v���˗8�TCel9OjK�%���K�T�0�M��*�J޽q�{֝bq���o71t�۩u�zO@�{yƷs1#��>e�W��ژ~�.�Ō<�z;���ޯ�t�Vp̴#;+a�3s�9����/M�>3�p30�DS�"o
�{�>�(��Ty|�����ڣ}`h�V���/f��.��.�J�
��U��4�b�4*t���Z>���Ȗn#���I����y�9��ܭ�>Z/�N�T��3�.�ss�Qj�TAs�r�.��1�{M����v
�B������^T���s�J9�H��=�ECʧE�Z=s����=㣭'�z~�#^ҝ�e`��%�g�ߦUzb��S��}���ې^O��H|qDM�>��VR���އu��y��^R�F�}Ǳ��N��ߪ�s�K��9�t_�\�*�i���Oo���z3ɏn��u�wwFz�MF���m_���W���wr�}� {�˻r-�m�����Z���l��̉,��2�m���sra�f׸�|L�^�?����^�,�S�B�T�����ֶ)����]ǳ�T��%%��~��c/Ӂ�\�t�~;'�:X���U����4�2�=�L��&���٧b���p$�
�)���=����6�}*T�A��kTr	wS��"�9:u	���I�]y
u&/A3��*�c�gh.��P�[X�VrX8b�v��CV�f�n�6 ����rŚ#D �7ig[��c��[սX�d��H��F�o�֎��^�<o�gTM|��t��{D�PӲ��UhW>���x��<��S�'�-�>��W(h��<���ǁ�z������׷<b�	�7%��ʦ0��w��3�ߵW�;[�t�y�cޙ�N�@��ײ�f����^G��>��q�F.3�}�ȼ~~�̮�Wl����פ�UG#Q����&u�em�'�R��;y���Q��?exu��CBV{a�+.�kٖ�b��#��H�5%����`LWz��At-wĿ*�>>�i���R�t6�n��m�����US�N��m����_�(��9U�;�qE�4���L�{V%v��=9RE���[�u�����<��m���sN�<{*Q�|���+����N��t��mǅ蘑T||r=�nψ�D6트��[f2;Щ3�o�i����X}^�Ř-����n�I~n=O�}U�!B����V���}.���t�:�+B�!�����ʙ��l�X�����3p�1�"�;7�=�:n�`������a�j��	H��5���#�%�2�J��]o��_�BH�Ԅ�!$����!$�Y	 BId$�	'�!$I?�	 BI�2@����$��BH�䄐!$�r@����INHIK!$I<IO�!$I?���!$��@�����$��BH�2@���@����PVI��WK�7�@����@���y�d���_��IQ*"!@IBg7kD	Q*RP���U��*AU.�)U*�5Z����pp��-V�iUj���80��W@�]d��mS@����֩[mm[B��(Wn�UZ�f�Sn�����*��C�n��(��(��	m�n�*[Qi��UZ�fjV�-uM��ʱj�M�L����l��Z�$D�&���4�EH[Ɩ�˂j�iYh�`&6�     E=�CIR���M��&4 hE=�	)UOP      0	����L&i��S�A*R�&A�i��F�0	����L&i��MD��ѣI��FLM4y56Ԟߏ����8���섄���B��@����쒤&	@�|  I	��P@��đ�?����?�G��8O�C�HĄ̄�$���4$$=$�A�)$����Wݯ�z�LO�����g���IHv��K�y��>���u���S!��(����������aj88�ݜ?�k_�m*rn��0��X:�oU9Lf�X8�yjP�1�2�������$��Sҧ�l���<��l���X1|v��S�Y�<bY5�4��I1U�5�M��k���Gv����z.�WՇ�e���˷�-r�
U��&U^�w�dލ � �i�D���ۃsm��ȳ
�R��9p��5�oaq�Z18.Y�ɔ���������Y+t�w�ʭ4蠫.n`���OY���	SX �0m����Ygl9V#�䢆nveD*��܋Q�u[̸(�,9m�m�1��[�b#������Fݤ1�ˬK/4��oQ�+u)�]M��/>4ȸ�h[y-��  ���T2 5��VP4P�t�0���q���Ch:,,�kS.��[U�m����M���[J�(�>�òF^��֖�9X��.�kU�i�ih�v�=ւ�Ů�@	��GbW���Zu��pT�����][7,��ihPbK/wR-�.h)ê�4�`]MW�4P��-����Hb9�[��$�akE�5��L��0��Vp�Q��Un�>�5Ĵ�[D ��6��Ѽd�y��N�,f� � �LJ�nPaQ�aܸOr�̅ށ�f�J�j );���JĪ6��6=ٕf�%[GvA�2�+���
ֈs.;�o-�U�a��6��H��P��em���ܫ�E�'m���zt"�(�/0���feF�4b�~��Z4࣌3R���cud���48̡�G@"��A�f�#��[�����3��|ΪVM�j��;[��.��6iMm[A�tf���[tE����E�nR�e���*`U]b�p�ܴ��F��{��1`A)��;w���[.̆�<�(�m���1ib��*��n�+�hSE��I7�`����9i��[QL�y�%^BtM��QM�b������]V�9u��Mq2�҉2^Tɔ�w�n��GY/HJL@�u����ұ{�oX^�R}$^�0�{�ܴ�&e���$nV�轣撬\�J�)��e��or:ǃ(��7�r���H�w��f�YB&�A�-`,���2]�ֺD�<w�c�.�o�A���#�f�"������yw0�MY�v`� �Ĩ�Eh$\i�2�,F���=�<��o4�D"�+�w%��L�a<�h���=�fk��(�����YI&�̒��&T"h%�ՄMne�yJ�ʵPR�m�B��c�@��v*�#Ky�SЊ�cYΎR�3��y�<�����DO�����#(��j$LU{(��8+�\����w��lh72��i�e�ˊ�;fH��Î[��n��<�82t����9ֽSX9(��ݥ��ؗq.+&nM�HB��K,͈+�.[y֝)fHҭɋ��26�@�q�J�8L�E�u��ž�mֽ{';�ںnksS�w�z�Yΰf�K�'���V��^>���fZ�]M��]s��^��{,�2�Ѽ��I-Η��V+;��n�g]X4�үT�	d]�Xգ y[_c]��"H�s����llж̢o%]��tu� �9�,��v�5��?)Y��[��cl��Q�G5�)q�	�8��8;�-v(*,䠎ݵ�vp�%�J��E6e
�.�Β�_h��\׽�]s��j�|��'?���A��tR*(��dLV��t@%]��Grī<�t�҇F���\<����U���m�i,uac�v�>����	�+�Z��XE���X�����#Ⱥ�
���©L�P̽O�ae<�`�0�S&�w���I����-(/��]}t���ȵ��u3\1Z��w�_�oǕU�E	@�]�AͰ��F���&l�P�Ӗ��Q٣K&�>\��Fh,�Sh��n�GXMe��fiSqW|���r��:�]�|�\�̔�Fp�=���Zܤ�ؙx���;U��U���Yׅ�s*=V����w1h����CzN�|�D���	u�LSG�nG���eMě��Wc�x��h�m�g[���[n�̊�����֔n�8�*WVPB�ݱ�L�r�sO.�L]�@z�K�+�C:��շ9��S�x�i�F�tk)�x"9Φı��B�:��8��c�-�f蒬v�Y�LNv���r�Ũ'sG�r@ЌՋwH:}v�����7��#��� R9��1%37�Lf#��v�Ee�����Q�1Q.Ҭ������0���}4n�Ͷ��&��b�^ �)b�j�ʻ�mV���+wq��u��n�aC�{�j�(mr2���/���,˦�P���5%��p�2d�i���^Dh,u�s���Τe�ke�����(%4����Unk=�*�T�����ٙJi^�݁k|lu��º�t.�v��@9Zp��J��\�j����2�-�1a��l#��L�ѶT"�[��9��a�8ߝ���+R��z�֯U��a�X��
n*<*��p�lt�hEAi��'A�*L2��K'd�)���e�1JW95��֍(qܴ�vw�vpŅQl��{P�U�b����,����G�����%uewf�6��F�C��l��>qb2����+�ޛ�Ls���}����y��_��G��BC��	�o�$In�p }��� HH}�3���{���V��~}��U��λN���VVKtAU���=����W.%,�����]��3.H�)!�0��jƊu&ZTemj:���ԎK�q�����oQ�2�FN;E`.ц�ɽ;N!�r�w���JY��g�	,8��֞G�q�Q4�����Q�Kuג�P������������:��Gtp��PS���Yo�Kj�AVY��c(�9�e�"� ��!}r�o��-��S�o���c�! ��GCή��:1Z�M�9w%r�Jm'��c�v���D[��6�����r�IK-.a�ugƥ��T�[�t�3K��ʓ/��
h�B1��e*�l=MI�vu������yNwW,�.}ɍ>{B_?�F�6C7 0��;��T�{L�|p�w-����}�"���U\;D���npK�ڽ|�����֕�M��[�������]����[G�j��Y:����c��\(,7��n��^�n��5��8\��uQ^��eٹt��4R8��%�m�H�37�3OaD�%���[[�$����4Q���U�C����f�@<�^� ��Ά�c����kE	rwKz�ap������:�D�F�� ƒ�͊��U���޻ٜI�|L��B�b5,SԬ������m�n����Zi ��WV��;r�k��;$n�1���N`u7��f�.�Ŝ˴Ծ�%��\��^����8(�˔���CuY��,��MR�j������۲�s6�Xе%IXn]�F�[ǆ�&;6��:L�S���t����Z��2��&�6�V���	� �j&�,����O��8�֩N���ctP/�j#����X�������	
�2`ɫ�ݔ3�_��W�����ZӴ�$ϯ��&p�t8h=��@�U��-��|��Z�=����v͆!�cy�<S�x�kF������^GO�úy��C��r��;Me�"������(�+8�O�޹]m�R�2ཬ�M����e͡j���E[V�{-؋*��,v��\~��>YY*�Z�*�XY�Ō�;����:�e�� m=�y(9F�*c{"6r�Q	α�:]NԆ�[o�	�n|��U{K6�w]'ݮ��bu���#c%����7�	߈��n�����n��--]2������=eL;��x6D���J�{[fT�Yf�C��0��_gd1c�[��/9b�lB� �&�7In�8C�x�Ѡ�ϣ;�ŎS"3�����"�8C���i�q��t�.L�]M6��Ot��$E"����9{�C~�&'艎�{?�Ĳr�E�p��8m�R�N��]A�Âcv�80�h�woo(g*ݖ�v!m71�Zz*�m�^voEƛ+)h�Ͱ�P�l8�^�[*G*ȳ9)`���q�y�Ge�}�1� �]Њ�;���ee3%
�6��z���slpM�|j�]�c�/
�ҹ��O�8kʔ"��{T5��Pӄ��VJ�u*,j��EUS(b
�i(E����R9h��U��+F[DTHź�,PU�E1X��5we�:>֯Yמ�1Y�.�g6!-�Dκ�#}�8��>��Tǅ̏��+�����M������W��p��)�2rP���c^���Z
�7���QwW���r:c�v��s��#8�ߐ�eg�K��hOq̸���d���Z�G��Ɨ@{�;���Cc�fr�����L���t��$��u0ϰ]�r�Y�}� �ۓV8V���w*��݇�J���˩S�� ���igP�-}]G0Z�q��t�����Z8��ĭ����V����͈Ka�xisϾ����t��"�c���!x�q웖�XOG�2�uO_[^g���9F	���1U�K������R�H3h���V�W�zhA�
�i%��ҍHc�|&�Ţ��ؚ���M��P���"�M�s/�šf�C�P�"���y�;�puk[b&N��eL�y��%dG��=Sf���n�������	�!ۘXq�+]#q�g�w�mU�6�,���g�$���Ĥ���gldn[J{\���k��)�@��@>T"�ޑF�}�V�܏�_u�s|�m$4@ߒ]�}�7lS��Q�=�}G~!���f�t"�E6lt�d��X�P7�!9,��F-��	u�P���Za��G��e
���l��WXf'��s�,(.S:^:o��<}|��z�d�X�^>�6�q���i�(���޻eVUFP�&`j7���Ｊ���,�`ȵpω�⣢���ko��Fmv��sφ�\.]=7(���_3TlWU�9L�8T��7� �����;b�U2��<|���T֫�++�Eeծ�=��}���;tP�?s��]c�𗻵�wRIMZ��;�pL�5�^V�Sm*���v}��o�����R��:�e,Q�j��!V�M���C�t}Q��uՁ��xk�^��֡�{W^���Xks�\yv���fv��NΦ�r4<uK/��Z�8�|��,kC���m{��������iF�AK�4v��f��칞���gR��iH�׼���YW�+n���ڠ�jd���4�ɏ��+���=<�D���U~;�>�r�Fv<2��,t���+�:3��	�ɼŗJ&���	�fi�}V�\�@-��:;3=�����ݶ�@�7OٻCt�-ӵ�j�]��P#s�C�-��V��u�V����ECm&�L���
�-a���.Kى*,�;���1�燄�zj��]Ǉ�B��#�`�2In��Q��KQ�@�V�1�4\Xↅ�wJ��0]1ib �ud��,B��Bڰ!X�̲q����Urd��Y��gZ4d�%�Ь��m��iX?�*�Ô��Yo9��i�)�)Zi���EE�*�Jj�bEQE�Rzp�)TRƬ�W@�QAuwQZ�KbS*�ԡ.���H��R��[H�M
�D�P�Jat�`���/��q�ι7�A���'m����{6��mOEGc�7�TM{�m#`���r!\�ڑ��
n��\П ^p:X��o��r��Ec7�-gu]��!wW:r��G)^yO�>�\�V�
��^ui�P%U=�{�5��iϖ1��w��1@)j~.�����Gf�Kf8gGX(��'�W����Z�; ��9�"�b>'GP�zo6�N��u��}�$x[q�m�}Y7sF�n�6m�n�k�J�7�QW�ADT��v�^�0!=%嚹J�_��i�N�6��
�Fwn���N��6���lK���^mxS����߄�+p=U��w���z/���fT���6v�mϣ4�u��YCq�*Dh*4����K<��b�{�Uaw�b��yU|�z�m m�P2�Kd�[ ^9^�Y�M0/��Cil<I3HCl��HWw��!����L��(<I&Y8�zB��՜�jHx��$��$�
!�Hd6�g� q�+^��9�b����P5�s ��FYkz7��9��w��=�{��|� E	� �!l�*�5�����$�$��S u�M3���d�ٚ������@�C)$� ��M2)!�m$U$0��Il$���W5�<Ɖ'XI�e�gY�RC,�� 
C�{��1�Hu$6��	4�2I���!�$;Ǖ�=�HaI鐚d��HzI
�}`�LB)$�O*�
�@���zĐ��$7ڐ8�
a'I�&!{�p�;ú�=�)q�w�&�rj='e8
�_�p:�f����s��._ƾ�Br�֪��E�-�ue��e�s\�F�<������bB��1B�'�Ć��l�X�w#8�n�a]^m�Z[B.9��
7W�k�m�(S]:���z�r�77�S�~�#��[Zz����:�)��qu�:_];<�Hݘ/}�*���z����&�:-=�6ܵ"WU���׹�:��X*k[����6g�K���3Yz�w.�i}��rfߩ��ǌ��!w������n�sa�2��L,�}"�l�pV��S�@|;cjvXvmml����^��_{E�5�.i�^8�]$���c��z׈6��.o��:�f�w�:(���+۶;(R�f��G��h箬�c��h��N����p~���
�]��W����m��ejc�Fz��D�5r��sa�"�qbl�g7􏻮��<�(Ny���6v4~bV���^�<�q� �}��X��)뤌����;n�L�do0x=,_��F����=�/��jyI~�uN�U;Zi�%�����ع�@u���CW�$���p"&�Q��N���sw-�+��1�Qs���&�C�ˇ9P�]}WV���!�FU5��mQ�4�7Yϋי�ӈWaT;Qr1�W�wX�$�yv�׿
�����8�7A�tYu�t�+�#�7l�f��J��X�5��)� Ù,���d�MJDN�r���թ��*n�t�����G��Q��`@L�J�lQyAH�?B�� X(�]�N���3�}^�/�����,b]N��˃M*�*�Y0�-�P,�X�V8hD��X�EYww*�Z2�hK�f0�T�����.a�"-�X�UU
��1Jn��,ŔU�l]!J�zg��w���{7��v��~�y��~��\\�����,G�K�R�n�Y���l%VY�f%��/�*��ӣ����ٵ�1�c6߅cki1�B�H�{��9��.��b��|-Ub��GƦ��j���]A5-ګi�;���S��{P�
�\�#|��@in�?3A�ۉ�Yߢ����5rO=�f;��Vɥ�3�K��~g)Rc��V��̯�B͊��NW�]#4(���cq��m��<�����������z�o�J�"=s��$�;B~L'��
���B�a萑3�I�.$[�s��.�v��F�����bo}�Ʈ)��y�y9��g�'w!1C���u�E��֤�f�ͩ2���������o�j��>��.��2��Z#UV:?xg]�L�CD���i��^R�Vb����q����t+�uv^��ەj�zL���ݝ�qF������F[u���>�"!ge��6�L�9ܐuW��C�V?EV�O۷���%���4<�9�)l��ޘj�(ꣀ �~a�9�<��wW�Ӓ����E�|0gV�kr���	ԄN��;��=$��v�؛-�j�[����>����ጜ�S�N�� 5[{a�1�L�Bݓ���,�j��9j@�Gv����%e���~mň�R�ǯ�-(Ȓ!=Jr��F�r�����He�ʳB�Rwu��&7�=������#����J�-&������$b˛�#�a�7[����S�?p����d�o�i�*��cq47�JcLzE����]�����2-P^��K��Ws$�z-.j�ݙݜ�=ԯfR�DDD.3�ͨ��K��C�2��n�Ve�����RD$�7�j�U�qx;r�^&a�S{��F�.5��s�q�W]q��=]�@��=Ř�c�zkK�8�G�}�r36��G�s߀�����pf"�
��R�SQ|�nԣu�Zv��T��1*����X��1*@e<A"8����/5����]rWE�D�<��۾�ѽa�/-��=�G�|�_w��㇪YN�c�> m�91ԏ$��ܬU��toO��<"�����lly���X��8���p�t���03rܙ܌�2`�N�8qt��B�.&��7��FI���z�o����ۇsws��6���kYD��Ǵ,��_��-� 0Uƈ����gV�.���v4op�jlm�P�8�C0R��4���h�����ebj��9V]��֎Ǩ����G)��Ysw{)_:t���TH�<�ؔw����� ��P�s���la��-J���rҩr<���/����ɗVc�6N�
y��+"]����cTK�Ym[թ6���y�eU&�xn�Z�Ɣ�+&2���ʊr���[T�ʶҒ�*�UtR��Ea*��R�b[
B�V#M����B���Uܦa�F����Z�))��)����U�)�ڴqCe.*�uT±T�iLi
����[j�ZB�5Qj�+�aiO7�p�����_U|c?���M�w~a���ԕz����_�����񚿩^�3�X��:]�.�xp�� ֩�|�s
��@� 
^5�^ÀMY.����I�;;�CZ� �7.�I^Ӹח�9ﾈ�����=SS��ޓt�S��o��ye\e���/�{3�.�ӝ{��[׳c���u�v1S쫄�r����2/�	�ٌC_ �O+���u~���ꨧ�?[ޭ�&�a®�eՊ��T\�rN2!@��c���ٹ�N�V��Ҳ�I{.��X�VwA�B�.���i�Lg��B�����]vG�����H'vs�G�s�}�ѝ���G��5װdB�V߮'��p���o��A�)�p9�fp,���-�6��Mǻ�����H)x��CF��lJ<!�|xm��y*��^�h܍#1���s�ٶ^�^��>�w}[�����ҳ��;5�?���:�px¥�f�/keU���)�Bw}w.�PcJq=t(�n^�\��	^e�B�oC��$��<?*��"��26D��6p2]n��՞�Q��-u��}�UW�϶ம�w�>����i\iɫ�c�^��-���S��+иfP���
���{gnr�O�y$�\� ���S�S���V��m�+r�kq·5�ޤ���a��O��>���ؾ�΄�!�ɺTw�.Na]�sn��zřv����&Ci����^��w�dZe>%1�4V��-��[�×�븃TkU����|���L��4���"�^���3�aM]N����5�J�@�)�.�n�[�X���%��.�U��u��ӹ�} w>kfM���$�3����G��E��i��,Qi��{�h�0۔�8:f��-ܘT���(������hm�`�ī+������ۦ)*�kt^h<M	���m0�aIƒ����;z�����|dQ*�(o����h�鏄�GL7�s �*~S�� �9u���Cܡ$��nU��R��p^��a����#ﯲz<>َ����"�)8���fFzf]��|L�Ķa�hw�ޚ�\�N�֓�����8g/>c����-;��Kf�oyl�V��Y�Km��<���2�Ln�n���*i�x�t�v�z�q2�
L��v����w�ݢ�IC��mԿN�X<I�@�)e0�眢�;`�n�~���z��L9��O�rf%��0�8-3t��U���l=x��;�I�,����6�c�w��Zq�|r�&�_7���(�K�o4i1��;�d�d��3����0����ķ�m��cE7ʖ�O������<g��D��ci�[��KCL0�N8a�Q��g0xKV0'�g52i��p�P }����ͭ�Z� ��}��̹�B�Qż�Tü�����^]	�9%`0�öE��d���̛ʱ`Nm`�d�:nR�+���B��Rq�J˘S/�a��q�E����-;u�+-��A�4ʽ�e�VwV�&	�n���d�ĉ"كef����]�b��I���m������=����f�� S���cotXh*K����үu>Hm����]��U�*����f���)^�*E�G�w.�c*�U9U�m�Ԥ��b+e���p���U)�U��Sm�ڂ-T�hi-)�ZQ������5M-+LqK-�r���-���.��)-�5Ku��F覑J��0�8�qU.ڹ�b�RЪ���M%���^�#p�o]9�/�DG�.�1�>���ʢ�I^Q�k�S�ۄ�S)6����l�w��y\v�N2i������6;O9�͡������7�<f�Z���ί�^���
f�-����\I�u�i��:��ٛ�L�h�qg��&�C0��;���ryTAg��`q��i���i�'ޥO0a�_���ߘ�Q��te��o��rlw�x����K��}���GO+�z=T�a�����3뙔���;R�N�U�.j���a-/]�u�۲��A_y��>�
)�Wn�o�V�4�Iiu���a�{~3���&�9��������F5A�ل��2�T��l�1�;�ܓ,����l�oʬM��ͥ��-4��{�3�q�-�yi�s�XT+b�n�}�}�Aθ��Ђ�hK�F|�x�{�x�0�KB�˞����Q�Ѵ�fV����ˆm���/I�3�+6۔(�M�Yή8g',��3�K��I���kx�n�2�CX�b����Yͼɇ��6�a��Oa���<O.�ٷ�P�����}DR���*����k.ӰUyH��#hI�n��ڿ}U�R����0��z�L�4y�f�,6��zf_IX�^�Z�Teڽ{���r�z�%0�Ʒ�Wh�+�a˴��D@Ω��a�n�Ǻ�0).�p�yF�����w0�u0̦���ß.���0���5�����3�8�Ka�T~kǁ�������&VY{5�s��Ʋ�3]������m��-�Ӧ�x�����|�2i/�E/5-���gq��6�i��Ae2��ӯ7�[\���1�+���<�1�:��sty�w[O�=�L!h�����k�y�����7�8�a���s��/�Ǯ�Go�Q����48�5�,�n�����X���I��}������M{���zh^�Y�����^t��������9���8��x헜Y�w]��C�,f����{��U*j���4Þ�_,��N���k���	(�l�a"�7X��d��awG;S/QW����T�%&�l�{{B�<�����k�;��|��	��.�a���m�'R�NyF�V�Z^�#ꁿU��
���ҧJ]���Ӌ�/2sn`�p[�����Nv|'�@��çi�ML��2�Zt�HSUF:f����Յ�m�
S�����0c��]��Ħm5�9�����AB�:�ך�z΍�M!�4���9��0鈝u�2�Il7�N�^3]���V^2g�5��O��%�S9�ދ�d����`�w^�E�w��{ᮊkiqf��Hn�nz�9��"�X��=1�驏��^MW1]݆�&�E2���k�Mn�9��x�n����l�Pw�a��k����٦�Z)�T��۞XkAa�ۗʽvkw���q%���Q|��oy��SN���)���3s"_+����p ��s���8�C/��'X�Eܑ�3�k
��F-�LQw��o��:Wy�}�}3�釡�Kz���4�M�L��� i���4�i�[�)^q���"b���������^�r��\4��$�X�z��M�ԧI�gz,���j��M��M�����'Y��nUJ�7����x����l��:���i/4AK��o|ƌ�^f�閘C�.��.,
ي����y����3#�)��}�V��MΡ
ce�����Զ�����Kq�v�Y��{��ӎ�Y���YM��._��,��h��s�l�kvn��迺U�e��c=b_���I��_��ef����t��<�@ �-v�Lʝo��nZ)����˞�A�?l�^e�/f��$��\q��66�.qu���.���n�r^�(��ieNWX8�H;Wav0��E��A�zi�Yқuɠ,�hvj�%�V%tf,�{�B�b�N��9إ�w��<���.x�����\0`{��'A��e�GI�֖����]�u��M��h> L^�M9��RɃ���h�w��!���2��ػSx����D3`�b�΄xf����Q�g�����k�tײ��;���B�U�W%]-%���Yl�Tn�3
�R�)���RQWm�T7AL(��R�1cX��na��h�T��qu�8�-EAe%��SL[n��5MJ��S��3	m8e&AqE
[J�1R�B����.�	��;�<<�J����;�I������F��b��}Y��ol������x`S%	5����}���w�����W������J���6�*�XH�����#,���2�uy�Z�|�J�0�E+�^�[:�gu�{�/�c��~H�UDb��bޡN���&����
��ᓍ)۳�˧9���8ѩ��ʙ&����$��]�˨�YΦ���
#�^��.9
Æњ�=�S溻nv��{����cs�"����-�Rg�f�z�4o�s��g;/^fZ�S�c���[s��mW��:�8Աcf���RIt�3J��=f̂���;(�~��l["����:W��� ���_���k���!�ӬW^^�9<y���ʒv��kpg�W��&W�0_��Rj5��Ŭ�r�MþW�k�N�Tn�`�!�L�Sޫ=g$:��[����pTS�m��l�z>��0^׾��y�v��R���ڻ��3&�<�Z�*����'�3t��(1i��;ԩ簪nE���P*�1��-�Z8��wW[��+�7�t�Pb~���4e9W�mV^�����!��Q��|˄�T��y�ϔ���Ą7�%��pn�|S5��@6��x��Z�׳�{D��m��P�Xf��ο ���TYA>�=�閧J���_JF�S���u�r��te��of\�x��M�
�����r7xU����C6+�W+T���ʍ��{�&�7�
c�I�W��9��E-8�vO������B��.���l��ʑ�J"���_�½��ۼ�l�H���F6��� �2�����g��˖��ש�ҧ-�����+ךJ�]t�j���R��V�C'�0�9��S��5h�KY��l��l�P�����}��?�Z��%��Z�k6�yj��T%�!v˴r�J=]�������r�`�f���+�'�-�)M�!�1y�3�i�F0��=S{ݽn��1�q+r�Ĵn�S�菒ܞ�r
Mm�@�0�5�ƥ���f�i�.��sY�\xfY^�˻�`v�x'��t\~y�������Q�����h{�W��ӕc_��ϱ����^}=xb�kC]&�)�['oi�ڢ=��f�|�s���8v�[9l;�N���ި��G�xK��NI���qs��դ���4
,CF���N��ut�J�go·�m��+�@�8�pjX���j�.�YciT�h9����Tɛ�ԭ+s~��6SP	�6����̲�S-�-�p���X�FF�6����5V�d"$PѬ�/˹)��x0;W�<ĐV(@�i$�����Xi#A�fL +�͠�	�*f�ݕ� pj�7�4 ˻���p3yWqt�U�>H�?T��P�)tP���-���Sr҅XZJ�*�R�J�Pi�7E%0�X5R�SUUU"��a�F*��8K�F��D)�
� ,�{�\9���p�r�M�m@�tbpk����~��k�K~[���_�Bķ'=�/��O�jΫ<��B�5�z��iy�bEu��qc�r�c���;��a!q]��$���˯>k����;=�J=��⯨��Y9N?2������ӗi�mw�iG��mD�Y����E�5�H�1<��vS��+s½uy]��{GԦa�LI�륕)�^W
�G�߶�w!�^`lrb�x�}���n���p���Wy�mݐ-v46?ˊ��S�:��o��P�`���|o�K I�����/~o9B�&G�JjE�Y����ڀ�����\�W�,I�E��*<�e�Wl�obb�m7:�N�ﾏ�9��5]����Q�E��E�Q�A�xpcw$�iv���֞EVm����k��*VcL3-pz��қ7D�93�*�P�Z͵N_b�
5��K�7�+z�����2d��SQ-��#�[�棙� WԜד��eZ۩�4'�䣔��	o�gH��1�Wjt��,�p��Io]��<t�w����/�����,ou����\��.8�wdcq<2��V�a��䊶�=n�z>���\���Dvoȁ�"*<3*T]]�c�e�xQ�6��Tk�G���_s��u�܆!"���)�=�Zag$�]�����"�'�d��Go�Ɓ�|�eO!��]�ti_�J��,Vd޼�}x&��� k(�co��T����l5M����#���\Ux�>�&����*i�Ib4ܑ�U鬼�0v��v�Ǽ�v	��쇍53���3ٝ[Sk���D�G0`�w��q�r��+$���d e��D_.�'G�Q��
\|�t���1b�t�̉q�*�L��q[�����2į#�3���<9�@N�r�������ģ���A:�r�M�m�[6�[�ee�vSճ���Ya_jgh�ѽ��!��K���,Lwglglc�r���"����Ğ��f�*ߡRߴ�0�\���	�s��\8��Uz�<Z�v뾞��Y�\�-M*�_>̮s��s{�	�tW��Y��^�ĿJx]��C�V���<������l�\�j�-�P����l=���sÍ8ͺ"����.�6���	٭��z{Լal��B���~4듺���u�f����("`H�5��I�ݝ7�;h�� ���VL�y�@F��">��[.�kBزL/$ёe�6d�z���EY����m[Xr�n�;@1$�Fм-�PeG:��f<�êe͎�e]�6R��	}F�P����qQ�6t2��bK1ٺ�`d�*�B~j:f7k�tZ��})I�v��P\�L����i�^#h
OH^&�U՜�@B�9ʵB�]a� HTt�E s5��Y�j͛�:hQAV��)��2���Im"*"�*#E�UR�EQDUPD2��K��H��T���R�Q�1Z�-�0�(��Ff`  ���.���Fja��f�X�� G'y��m��^X�*_���e���0M�ם�����Ӊ���3K���f�ti���
މ_�I�-�T�V��H��hE�9�����W��a�]gD�>�g\�����6���2�;��(X�{Wx�r*|�4�s1�*��A`n��+9=�$7���#x8���:��G6���Y��F�*۞�l�𬧼�<r���V�^��f�
��t�1M�ӥ[��Or���g1��x��Ez�P�D��k1n�E^ܝʂ�(�-
��!�69nʼ�߬��u�5��WM:���E�ƞak<��2���`�d���M�6�y�r]��ᓸ�\�q�ggyA��.ן��|;0���Y�
񵍸3I��=j��D��Q1�������H�}US���Z��lr�~&)Y��F^ptv#b��[q�^z�̫K���7{��N������۲{�I���V�>˜���5�;QF�#�˝�d�/�O��ð�:����7y��V���3���*�y�A�tYM\�|���9q{�,�uH-[�|W�ϏPM[���{�W�^w��سgZ�"Piv޹RΖ�����ڙ�}��C�*��8ќ�/Ǖ���U�=�L�+�%���Ia�	3�m�2�jB��YVH<10��>M�@���ut�
��q�̔���]�
����|Gq�!�wn���ci��cG���se0�����+�!�gl�+W�^Á�lPO<�z�:=���\���#(Mn޵qn$9���8z�\9���3�Ғ�dge�PM�p\yu���Ec{���a�̙�\�ԓ��u+�2�a��0^��%�!�>�pq�.�ѻ��^��V�s�B|Ȭal�6��k�{ed�<8$�i��2�i�@�]�V�e|%kٮbwc�ſl.�������4k���˽1<l�K�%v��pK��M����C�Һ����r7f-��2�N�p���g�:1X-I�E��h�͒���/b�9��]j�F�t�g���j���C =+��y.ts���|����ɭCVA�Jg�c�Yz���D�����s��e�#Ue?���<�Fi{˅ia.��Z��7ad~�wpp�
�U��U/.l�۽-�hp3/��Y�D�ܳ(z��8C,k�r��@e�w �7YRh7��!Օ�+�n4p��E��U���g�f����g���˹����n���}�:�F�
���B�bס��Z�Y�%��֍��)E�h���F���M��tfR��ec\������X@b��wP���S�t����p�I�`6�6�!�zi���i1J�0�C/y��A��SJ*(U�qU��Q(��IEST�M�A��M%2��(�QV��%�2�aQ���TTh
D� |? ?[�y~"z��I}׸��l[)�;�-P�l�η�rb�mz58�:*Ņ�X;q�ЫS)j�]hZ��*5rt��uc�9Xr�{�V�T���Atmf����%����τ�#��}3<���͵����w�^ݠ��nN�]`�fH�#g6��y#����:q��Z¢F��u����Rŕ���ҵ�?U��W�� ���,������U��yL�ײ���L�j�.̗Z�
��`T�:0^e�D�Ӕ��`�k;�^z����/��❨����G�xX��s.��D��+bt�dt3�����Q׽n)�ҡ6{o��vO�W.�s��k`���6��[ݺ0�y�C��cM�⾏�T����m��G�q��s��ݶ]�l[f<2�R��`�û�b*�)X+
�E�"7Y�L�v%!ȅ��"�V:���_�$1���?1�^�IHbȨp�OW�}�v�)(��q�����f_�`��;����L�&+���,���7�7+�(��+��Ϟ8��ca���i�/�t�Q�:�f��q��̩"��_K�C̾�ײ�x��02���t�J��t:#o*3��,��+s����B>������{pfB
�lmr��a�������t8����\��!O	rt�"�z���^����j.�gֵKW�͛�&פT��i�!��Q��ٛ^B��^ϖЊ�{+@�#�4��~�m��1�GQ�����Z�fj����=�WI�(��)!�M�%x�.^:F��8zn�h�1|2kcqe�xj�0㽫����<�_j���ƭ�^lc�����G�K^�/
���2�?9=+�˼����K7�`�g2�s��p*(��S^��� uSN����,*��`���x��DحJ'/t���ނ4��k)j���_��w��$�vQ��+D�@P�E�Z�P�yɨY�+u<J-��a�3��/�2���ٷ�y��U�'�u:܀m4���-�Y�U�J6ʯ��i�.�.�ּ{���{����#���q͠�&���^w�ʛ2�Y�<�!�����V�Xk}1�gnL����\^�c6������������n��T�����j�}�d�L�V@wF�h��J��v,�̤;��S�b���O��dT�r�P�$�V�sE�u��M9��K����������%��������4�K���(��������J�ֽ���7�^.�U:ӱEJ��݆*^Q.]4I�� x�������tV������Yۈ��������L��UH��|��2>@b�4��9}���g��k�X��]�*�9X{
�"vf�ŭ6�
�N3�Ӗ��7S��)k�[:+�7ys��+�K�Q����[�����6Q��H�l�n�T���Z�w)n�X�ғe�&
�U&EQH���RUP��XŪ
iN1B�*�sn��c�SE��-d�|�u�w��!���;�v��-���PV�*��;�����yɘm�7vs�5f�I�߳�I͔�`������,3ַ5qGw��QwI�i��^[�J~bj���\W���.���:C%7�k�/��5�muo���p�<(�cw�<��xv/�䆅A"c���&��5[�a���nƥ;".�������W8u���S���{P�<��f���Z��ZGҘ���IRwlʝ*>������x��<�s�6��KNV*��sJ����f�[�=O]��񾙘��Jp�:"�tV��Z���3<s�m�]J��w1�5�!�����nm޷��F�-��u&���e>����	�
�#s���K��xn�c�-j��^
��%S�h{��nX��>|�]��ע����vUDt,�H��cE0w|\��zS�}3�N�}�ku��hb�֖�l�ym�˼o�R�+�ae5����^b���}w�{2���QC9�M�L�Z����p�y� O-,T�Y��������A�[Z���o���]is�ȴ���*]�C[�2�U`��A�0��峥� u�+�  ��.�3c�ر]����Of5�{���P��2�k�hP���F����r-�؜ke�-����$�T�K�o��{j�9��)��!���8I(ͪѾ��ϕ�
י{{�-@$��.~zԺء�wO�?!�<!���^���nw�<�uұY}Ѿ�'r�8һ�'�{��i��5k�8�?�+Ox�0��B�靾�̆0����6�OI�e=���Y�r���my�Z�ڮ�����R�9�_]hѱ7PE�,����/&�n�zҞ������j�����4p�<���o%ikm[�EO ^Q+�&vɞ�~�[��G<�Pb�������F��ƫ)bRkko%zU�Ҷ	�>��7���9x$Z{�gNie�җ3��uu�bq���érqً-?t�!��֝��)}�x���E�˥}��ɾ�+Ĩ���S�h�����w��u�w�*�L5���>G�O��>TSJ����U����|��IH~?��	!	S�S�Te`�[�a¦4��q���Όx�	ְ�HB@ �Wf6o�a
����Hl��{��nA�RW��=�[!!	�$_k�}�Ù���z�����O^OίA�?,ϔ��8`���Z�A�W���w��7�
��a��!��c}�������~=��~�q��� ����$		��ȑaRY�����'Ƞ�����~��Q�}�������>���{g̀���!$!!���_����E'��{��%���j}ҍ��O~I]'�d�I_�W�^�3>�������W�;�v�j��$����a$! ���L3��q?e�G!$!!��~���c�Y�,��J6�W���l>&a��O�`�~$!!�CI
>F��|&~'�ǲ~���1
��T�0�܇����$�����O���(������������ﰒ���(=TK��q��'�'��'��Y�b{���P7	��ҿG����>��E�>d�ϲ{���~��k��?Y�Sg���HBC�>�<�~���?��=��L�X������dF}U'�HHf%ϸ$�$?�����'\��O�ԟɎ����6d(����=�!		�qj�	?i.X���8Ok�BHH#&J&f�I�>A��1�z_�A��L�'�w fxK��T��aU'vg&XPy�IHvX}����������$~G���A�O��ɇ�������{��������%�?����>�B��}r}>���zX~�~����_�|}�����HHBC�>��ϼ�?U��?�9����I��5�ǒ�������z�>��{��	%���?O��a��$�Q�����o�_3�$��'����Ώ��O�����_�囝<��o�=�������O��;��_(7���?�	���� �}	��(�ժ���`���C2O��{� �����~DOxI�)�?#�7�>�l �����>�{��DǳA��4ML�:�#;�����&��a>�O�*I�z=���s���H�
!:� 