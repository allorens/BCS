BZh91AY&SYi���_�`q���#� ����bB>�    }T }j��0hf�-h֤U�4IF�2�F��EJ�m�P��Z��ڛkV��l�Cc)�m��ֈ�i�CF�Q[aTd�k�9�%*�&�mj�MFMK*���[f�3kf�[Z��ֳl�i-��f��Y�jٶ���d-)D�)Tml�kM��E�*�Z%����)��3a)(�V����f�V�*�����V��*�j�hfTհ�U��Y�l�Y-�����ـ��j�e���6�hm�Sj	[io9��K6D�H  �ܮ�]�PT�n�v����lЪ25�sj�5)� Z�q��[(݇D���Ƥ�W`�D0��k�n�h�UR�wQsb���D|   m}���w5������Rۭ���^��U��\z7��K�O]�Yl�jl��x��m�+ݽ����v�Ν7<n�ԧ�;[f��+�i��W�n���WE�X[Sckm�mFMi#6T��  .[����Km祝*T��ۦ�z�<�ە*�U�v�{Mv��$�yc�K�m�6��]jjK:�s�f��Tҫޣ�֭���S�&t�evն��[��.�N��M�&խe���ҍ
le7�  ��צ��[����^k%j�*����R�O;������j���]o=J�uܫk<��շ�Weg�G�}|�Uf�<�קK_m���jTem��3��j�����e��J��E����lĄ8  �d���h^}y�}��A֝�]��͘��}9w�/�}>̔�T��=T�n��ɽ�ڍ����R���z��g�9���Wm����S�ց��<��	�^�_"��(�[h���m��l|   M���ֵr��OJh���=�}�����ﴻ�6ԡ����}�����a׫g��W�^�nxM5�k��n{6� ���O{�={j�.�W��;���i�q+R�Ka�kM�6�kI��   9���26���ޕ��u��;���Vʭ�FV�ݲ	{�ޅZn̯/��J�k[���/^�T���'� �b���ִ���ts�+Vfٶ�kA�6j���  �Nz;�����G{;��Uz�gV�����T��q�(wW��Z4m�˚��9���݆��Ǫ��R����m�-�� r=��Ѯ|��(��;�P(0vӓ�v5���QW���=5���P�:��/y8֞���n ttvt�hѻ��ئ�(�l��#fPī� ��}mn�_8�zH��B�րu]ǧzP���F��.:({��P�WJ�n��OA����]�G�     L�)R��L0 zL ���S�h�)*T      O`��U4@C@ T�R�@ �  � O��OUU#M� �    R��4��MLMI��@1=M3)�y'����~�����s����g�;.�O^�잞쏯�����������D U����}�T�UP_� U��?��������T�1V��?Ǒ@_���?����?���=�����?���Ձ��/�#��_��������L��L/�G�#����dL�S�L�e}2>�L���#����a>X���dy����d}0>�_L�=0|2�L��G������d}2>�OvL��� ze}����>�L�'��"� �� |2 �}2 �y�0��L��_L�� �*�� ��Q�9�C�"���W� �W� �W�W�"�ʾ�U}0��TL��@�~�E_�"�ِW��`�0"̀ّW�� }�E� �a=0 �� ~��*zeOL���( zd&UC����ʨzaT=2��UL '�~X}0�>�dT& � ���ʩ̪�aA=0���POL�'�P�"��`D�ȡ0
�UL�'��*	�P�ȢzdA�d�ze=2�2
�C� zdL/��`OL����0� {�� }0��+���#�Ȟ��ze}0��P�dMQ�=0�@���C� {����>�W�*�_fـ������>����za}0��L�����a}0>�_L�'?!�	��}����׷��=T>�:��Ҙ���Ãc?�b���u	Uy�OŵA��^*p<_^���spM��L�O�qk������*|Y5l�2��{�bf�TZ�9^������[Yh�����4	%^�PK"�mmX{���N5�x-���P0�y��m�!�C몒����Lܖ�bէ%Y&a}x*�!l��ц�؏n���+7��6�Ӱc IͩsD��檲�n4�f�&��V
؊����
!�)� F�Jx5&��R��JhZ�su�̘m�^l.���{	���Nk:"VD�{�`���iK��b��*�l���A�(���Q!������2�7�G!OϢ�N�%��+iP�2�i��f4Yzo6>��k�n��	&�`�ܽ�5�A6��&�V)错�&�mm���i��͋l�'5Q,M*fnMf�d����S�qd��VC��顳@ʳY+c����v�A��)@Хu�C^�Xu�ˬ���U�_ۨ�VѲ��F�����Yd�H:��Ք�Q��Q�n �ݎ�$�I^c)��ސR��������U����m�e�u� ��Xe�.%�A��cR��5��(�Л�V�YWr��vp��Z51ceMJ�&��ĪZ�/A�+1�`��7n�x��b�l�t`u�Tf��sǚ��N`.��x,��H��:�=j�Y�Գ��Fn1�dʳ,��#��N��B����L-b���
��H��zeQO��yd�{�#2��YgTWX�⢭�'�:c���d��N()D]:�Y:�k%���J��H�$�(���C	�K5�z�B����Ǭl��ᙅlC�[̔���"�a�� m��A�f�=��n\��.y���v��Vji+2`64T����n�-�D=��%��a�̎cȌ2\�mo�@����AU���j�b<9V�j��I:�kV�>cr�'Y���Xl�۴5h����'
��enQ���4��1��ޝ�u���x����� 
ra�5j�'+ǗX��a�z�ѿ(�h�[�72�[��X�*������e���uYL��1�m���C�'UVG[7���IV;�M�B���vo �v5���H�m˷NQP+kdd�ñ�*���m1��:�٧MI�X�weK�E�����n�Cn�ec��q�5��a{���	5�)V��r���<'Nf����IU���/"a�4��#�7sJ�1��2��lcP�TȫP��@3&i��&����6�.����oV݄)l�����N�T�&��h�)uy��rF��%�׵RU�c0���oH�(�x]��Xu��oS��}5�ǵ�S�0���lІM���=�h��5�"���V�1e�M�j�� �3uF!t� kz�Ң��g(��^V�'Yk�vV��^d�Ve��%	a��ܒ-��[lC���������n�!
v�r�+�l�K��y�Z���z���oN؏i��53%=�)3��v̵GT\9C��yh��[�E���ɪһM=*5��w1
��:.額P�҅�`��<��2�ph���e��S0d!J�l��d*HҘ`�yaն�6906��0�z֊�}�b��-���+a��Z,�)�#��Ɋ$`C`���!�ؘ�AvXU�3�&�+5�v ����@�4Qv�@iP{s�I�_���4B����!�X��ԅ�E�E-��� [n8�m��
�CH��R�PF���,��}�Qj���	n��*:1�@�z�{ˍQ[�n�c�MnVcv�z��c/���V3#���߆	ZB�-�-1�*aֈt�#�N�&ƽ���F��J�q3qn�޲`,y5!{7k����6:�%��/���H>i�ooh�EXY���x[L��ݾ+4�솹%c��/nMXe�u6z�ԣ��ecUg]h�<�@@H �jÈ��ޤr�����dgQ�m$p+�ѣY�4*��klřx6*,13
͊�0̘'a�)'nd��l��5��p�q�*�Tbn�pŅ,(n���+��	賉������ 7�{�2��hR��;IQW����JZ��˲i�M9����6���RU�V�.R·S:�L��j�����'2B�/Lי����t�T,�RǪ�Y��!�U�U�`�GH�	�a���t��W��6�cX������jj��7]3��Zn�'0n�ֆ����M�=T�������L���p�t�y��W�ۮ�X�$R�Y�F�r	�h]hL���iR���R�_^[_���d[��ۦ�v�i�82dr�6�AR�:7(m����kX�ݘ�j��*ec2bWk�X��1ZV�E�D���LT
 �D-i�?��4�nT�%�	R�;��U��2p֕�y%n�Ip��o���:΁m���(P�Zdd双���)�Rv�Cw��MK��$��jn��;eu<]\�6�7��un��"t�	`�]�Bu�˶v�մ$��n��S��^��"�#����ehWZ�t��n�.��*K3� ��+14E�P����c0��m%4���'��(ܟe�wuBPI���.L���u�
v��U6H*�1R�De	y��ź��7u}����Uݭ�4K����x�/���;M��r�ѕ�Ę�����R�{��w��.�����rKn ���T���Mܢ2�����-�)�<<�a�i�΅�A�:�(H06Y������l�\��͊�����⚘�d7�۶�xN@�U�U�/F��Ѝ��iЄ^��oU*hH�ݲ���B���YF=7��:�C��$Ɯ����.�v�S`V�!��[�ri�qsv-K��N����o%��[L�ѧH�`����M�&�ї��Fժh�W{����Yf�>��ہ�kl�����!�����׀��v:	�r���;j쯭��=���U�<�r�mX�kk �6�*�-��/V�`&[�[,m��C�^ʉ��k4���d��dY"�4-�O�J��-l�DH��3���fo�),��%P�JO*�KYv�i��?�H���U�v��\�I�͊z�]�p/���&�;Óm��9�	�ّ�i��໶<o�ԴA��V[���TtI�f
7ZEh!lH}�Y� H��B��r�ibf[�]Y��^�,���W�B�HG4遻u}M��q^�!�5-��Lu�S,�,�����;�E��ˊ�1�gO�������F�n�L �j�����]��5D���IYw�x	[�����ٛ��w�[�����z.ҵ�"���QՊ�������-�[n�M�Z��;!��ܱr��z��)�)I��R�u)���6v�iԸ��"�2J,b�_R�]��*�I��tc)7��2e���f�b��Z�7w�ަ�.q����\��B��*	,bw�*�dKP|/y��������d���y��T��X�uY:���v�G��zE�NLWq�<#��Rl�v�^*LW>5��s�E_oͷ�k��y�P��i��: c�@PZ��HTh�ة6�?�Ħ���r�xV��B,���l����p9�NY��m�<N�*�{��еw���c`L�4)�"(j˖r�bOk5�ߵH[��&fn��s~�����fƇs.��LDYL�x1C\	:�ma�/�0�Dm����f
�e8���L=�T�r���AG]lSa'R��	�u��"e��f �\�i2�S�܁RI�4�Re�L���[�~�䷭7�E�u�������X_q�C�a��䚥k����]H��n�q1�����n��]x�n�i�6�`�Wi�k1��挳W�T�̹��6�8D�]��
lW���	�����kw"��͢b�"΄�5m�z^j� {v- ^��ܙV2��l
$"2<�-hT�����r����p{���H���xl׌�ފ�F+D��Lҳ%n�%}�>���&6��GS.��ЫܰY��u���m=ia&�2��6��Vw4� Ge�a�_�eK5�&�ݟ��M��Oj�g�2��iP��]�ͤ���gz�>`7�ku���,2DY�5��S�2�AuV0=�iEۊ���C&^=%���Ce�Ԭ%kX�1*���\׿4�.���w��t�i�M��fǒ1�f�zq�1���f�f�9 d=[~Wv$ˣ��&�#����IX�	m���l�_E34f}�y����2���@��y��ց��(o�՟Fv�݆�1U��H��x`�]��a��[Ÿkp��9�P7�jF�ɧK)�M>�]x:�f#a'V�kZ��v��G^�x$o#om��ɗ���n޻mf]�%:��V����rR�D�d��t��(�r��2���Y��2�V:6�U�( ۧ��tݠ�{엳@��2��^�� �i�_;sv��
�F�i�	�J���:i���f�8�a�V�ٛIb�B�3(a�����9�-��d��]�R��T�j�,��.�Br��V�zʙ�7��)KUW��hY��_���&��RYq��0*���*M��D���i���;����r��i�Z�0;��;S�3*�);9*��i���	b���A0sd�^ on�SoQ�]^�0�7��Z��6�֩+(9������aݷv����4C�]���ӣH�V�#0��M��O1,��C[cR���LNV����)�Ov�'3i-K�v���NS�n�y��͕����

�rA��P�s�����X�YA�3��̹Dw1��l��k�{
�fɼ��N���f�y��Mcӊ���l�r=�r�4o��V`����R�|%��	�C]^0����ES6�N�&N0-��Q7V%��lH�f�7�j���Y[UvM����t9�
{R)V�7d�*�3����j�m�Kw2y�޽i2)NIcp�f
�L��=�V4�4ؼ��FV����c;7Q�H�ưb�&SC�+cFd6��54�n��3BAZ,7�S,<kO�7�ya���u�b�c٩���0I��W�`��Y��jW�.���oD��t��i��!���t��,m��N��A�N[�H��<�Zm���J����*�c�˻�`��5�.�$�C��/	:]
l�9��C�v@ѬJ�d1�܎��e�osk1Q�K1�GRlL���0^��C�N�����Z/@0^���v��w6�
ʺU$mLxI�kjJ	���i:����ق�AKm�1:{h�5�q
OO-]mWShn�����KFM)�墅pJ9O��0�e�Ô��opBdH6�cq��F�z#����q��Ա�ԍv�n��B�S��I��Xù4PN�#(�݅��,����=ٱ�*�ڟ2�h� As,C�\ݺ(^a܌2q�����YӇ����0��i�7MR�pf���SP����4�
�q���A��HӺ$�����s7��Nm���c��wx鷗�N�:#�>s*=B���Jol��W[�ۂ,��6�Amb�K 8FYYbV��Q�K5f3�*&٬�Ѷ��Tja׸0�v�In��̉�ePn��x�jݩ[����Jf��V�"�~��?��/
��m�uS�H<���Y%Le�7&��+Ry�YT�Wj��s����n�]!�4�l�H0�W2܆���`5��n5Y8C��^���P���Fn��cѺ�sI��X7*��[��N;���in��2]��YR�V���qVI4�Ya�G3Dg������j��9���5�SpGW��i⎦&�-�,�$U����ť�.��Z�| ���«� `j���]⒢���d�'sT��^���a�B����
�'gMA��Q��#��"���H��'�r-��ܻx��(�켣Xx��yx�U�-��C�y�4J32�<����Fa���{����ӑ���iV'��WVqخ $:�i]6>��ո��ۻܳ�nc\Ջ(ؤ�l��aTYX	��=F�M@,<�3u�������م�tră^�	b�^�b�7�(94ԴΜ���8��F�ó(У�1Sf�נ�{�Y�g���׿;;Gt�x4)����E�K켺Be�c��[+��0�֩��v�X��)�7��vD�9��3a�.>,m��q�Ee#���I/��WN*��0�OV�2+����دh[�b��4��	[jJ�f�u��5!{�`t�ʓ1@��)"�yGb�{	&�e��[L#J^��ӴNk���u����� *Gz#�u��n8,1�컌��-X�<,G�[�S�]��xNd�%�;X�6n�z�A��0ܗb��O��ʗV39b�幒R�ڹ$�� )[�+J:�%�����&�)�E��Ì��.����we�>�h���-ř��e�f%�[��
V�'r�VPO�A��X�r�OkJ��l��+^<ؐ��eK�^ʫ2[��hG�K>�d���x~���dU����� ba)�&�jؽ)Eh�Qf:�ᵺeِ�%��*Vdˀ�5j��ar�[2�@hV�l��вT�$H�cR\Z�f�tLzS��e`��IY-ި����0�ذ��o�T�Ǉ$�S:��?����Q�P��P^y!��{7�ê�0X�3�x_pM b1�S�	iA-��}tϹ���yؖ��`|�xñ�	�-j�f�D�c��h�$��Y�&w�� L�˾�p�N�Ƥ�s��՜��&��Ub�#����2	������U�
  ���Š�N�U��B��J�0uZ��,>�V�"��k��H�a�48A# �u��c �6���l	V��x@�,=#R�,����d�d9���b����Ԗ-�F�D�ڍm�Ȃ���s�	�� �b��@�0�¿�h��>�%�������O�Q�O�B��{s�b��$��Ȉs;���٭sJS���d?�t�����W���Z�"�Ւ=����β`�^k���0nl�-7hu���E�`���oc�$4y]t������7*��������d��iM�8Y�iƤ�w`tgP}��9m�XI\����w��P@�{��M���*L����]��oA̳��t��Xs�m�ܹ���]�4s��M(�d"�q.�q���)���.��QF�i��$5oh����[9��Dkr^UƳ'5n���T�"[K�7m*������whc�o�B}���ƜV��S3/y�l��b�}���9M��+̏4C�r)j���ûzr0��t�׋|@�TB:��B>��\���g6�$��Ov�㓥���y�qČ��{�\����{��	W��	D�C�Vn�W�;#���'3r��M�A�%c�*ZJ� �t;�X�rԷ�w8b�qN(qXQ��.��İ���+c�V\�|��Ȱ�`D)w��L�/�԰2��n9�i�Tߌ�Hk�]cr-"���&�2���mR�4V����0��ErH��n�f'��q̷I�֕�M���Ԡ�ʪs|�a���pg"��T74�JO������Ä��Þ�Ӥ�d���t���yuqj��F�81M�wo�i�ޡ�V����c3Qhn@P�&�)8�U�rIV�i��鍯x��O��)���(�$�_o6�j���ɎD�E_5�Jwn�����l������w���j)����ȬmLa�Y>�vhv�vs�T̺���6U��Z�tqtu�M풚7���y���iwг^%���hK�(�vl�Rw�ls[D��s�D��i^㿵ʘ����+���#��Vkd���lb��0�7-g*�sNR	V��R�Y�.})��fѝ��crN��ޘkZ˰��tÌg]շ� yZ��*�/�jw�q���Z������If�ЫgV�#V��^7`������z�\4[���QnFٓz�����U�a�3+t�Ѫ=|�on�8�#����&p謌�wu��ى���[����ӡ������T�̸�.��!�u��R��2LR�޳�Y�my�s�z�s\��|業1�no!�6u�\k�#���w�l[  �"��X�с��\���S��y�0-7dy��+��j���,މWu�t1�sz�g���������1.��F݇�,���-V+�Ӣ{�;iف��Z_��w��n
��,������kC}�ȫi�]�3Z���HJ���H��ݎ^Q�$��hK��g�%�)����[P�S�KI&n���pnZztl�Rݎ�:������BeYt$��ܖ�:N��%f"�#Km�K˾��U��[��kDqyj;eM	���l��V�	��? �i-Xt�9{{���N�C�(�,Ѧ�[��7�K˝8G�Mtt����:a>k:�+�'�
�M������J�z�ה�g�3r��=���3�i��ᢠ��6
u�w�����n�tVcd���Y�{�F�a��*�1�k.���6EY���ۣ߬��y;��@�$����ol��FLRW1�^ҬR�빵�9�*7�t��V'"\ף#wtE��Ѕ.��ܜ��}!�_+�u�U��LyWp��U�ݽ�ǢJ�ЯӉ�We��+��^�D��r_V�����P��Vv܊��{�Yn���,d-C��}w��4%�W8�*�*��KyݶX�j���p ��헗s�kS��<,�z�7�s��G_P��I�&J%9��+�;�-�0������F�n�9Q����v�m����6;�hiZ�#F���m�s<�a6��p9�f��c��뫻	��Nv�:)e���H��n�����r�m�p�^���ͶU�]�xe:-�!R�/$I�g����ZxF�8�/v�Ξqf�$�s��}��*=ޖ�t�e��iݹ�]u�EF�jƦ��z��D��;ͼ#h���#��A"�+w���kRق���ׄ��4dvӒ�����,A�A��HуGWJ�z�7�G���ۻU�Ke=��/����1a,�X+NFE�&�w�s�rX�<n»��+E_[�Ώ*=[�7�l����K�MQ�2��[z Q��yy��}�'dA�5�w�i�Q͂�!'D7��ֹ�=\���pT�1��u�g4)�e��Mw�"�m�Av�R֬��v,�z�"����w�W����M����-|�rÁ��|�V`g�v����u��"��B�4�{"�P��ؤ=!���d���%�6�>�6�`��(��w�����/NU��HX��Y���#h8�ls���hn�mqAqm�*�B�vXY�IVTjw];�ywq\�Q6��N�<v���ū���&��o��Y-�����I��]��ޡTQڵX�	�dE�1���]o+J_�Ҫ���
� ��Җ��<!۟$��w��S��t�݆��r��͐r�X�<�#�}�[��8��UB�4������k�f��9ׅ�d*Pɭd�{��WZ{(Ê!ՠc��+R���)7� �$)}��t��YM�ۤ]�";���G�Ǝ�F��=�2�wk���1���@Ͳ'1�����q;�rDv�x�,n�g5�3L��&�)����-����ZsM�D��.T�����]���3���j�n�*:7��M8oe���G�����~LU��ՄoT�Gs@,�t��3����<)�%�ea��og[�:��2��7J���2%�3��^������uG��|]V�`��%��D�v�U��\���PZ��,����-0ژ�.�|:�<��M<Hh,��s,�u�o0�ӳc/!�y�/�hS�o,b�Y�{��[�y}t�q�î̭,:�+U*熣��Ʃ�w~�kZ���Q�
��}�fd��'�8egs&n��F�����PH�Ļ�{�m#�+����^]�ܴh񅑥�դ�N��KKsj�lY��μ���g��Zۄ��'��M �.�C������i-T��o���7d����P��ۛΙ�F�}i�v��t�t���ʙzVѪ��7t�%hP���+j�]l-=y����	t��`��;�_�/[�z��6U�ef蝳n1�ه�s��&�.��˵O�]G��2`ôA���,�d�
��9b%���JB����RO-����|D�7O{t�DW!u��tt����m��E���i��G#.a�z�����8�'+��\��A[u:rzƩ)������c��{ot�	ԝ�.��Ux|=��æ6�O{=��q���N��諅�@�7{d;��eiYN�m��e�Id�w�J�꺌%4���j��4�w}.�@���źo`�3�os����$ҽ�Sgi������Ǌ.*�e����y���M�лΗ/�nk�����j�ΗV���jm)�v�'7���Z:-�lE�<�^4ẙ����W'�溚]�x��c �qs}X�*˿�S��:Yԯq�a;�J��A�����wW�x��Ô�l��D����tN8O�u��B��}J�N���泶� ���P;-�����+F��y��t�v�[|}�E+ykL!�L��,�N�B�z�v�}9pD��N+���+ͺ]��p�Z\֠۠�(r=ү+y��o(u�l�4�O8��vPO��&�pz��!d��G�!ռ���N=��:��1��儑�.wawqbw��h��;�ѧ��{��^��~CM�I����ԓ4f�ۢ�RY�i8�򽔷�a��L���!���{�B4"'*�kj���p����y�oZK�5�[��7;)��ĤU�������DDG��#W����o�7k�ζ�s��8�n����ow.��Us��n����<Qk��U����Hh��ze��ѥ��F�+��[sn��la�)� 1e�v�tp.�S@:	�DB�eu���J�Ngq�pE�}Jɭ��6��D���d��X��."�M@��Y�2���]{�Wa�ڼ6Q��7T#�����c5wU�ZAȥ�c3BU�N�m٘�F��Y��Ԅf���
�b�f�&�ԗi�u�H��̽�Տo;���C%�sQ�\p�Ʈ�����^���(,�����b]�9ǂ�
ʆ�k��oqMi���/y�0�gQ����9�N��1��Sc4��/���$,�;6�sf�s2�=���dp�S	5�B���/�*܁v[�>g�k�]��6iM�ʓ�p��4��/��[�Rt�ɚԲ�5�iw!��X5@�����Ɂгa+�<Y��3629�s������S:�嵻��1h���:�U"놺):�2�֫t���K	�D9�
dj���c�o�v���J\/u��+�H�&j�؞H���ʽ�+
�̼��"�Eg�2��t��R����uЫ��n������]�t�oF�t$��ýΖ�t��ڟ�i��}�t�-vȺ��h�|���6��U�F��QH�w�GV�)�!V���7r.�+n�"��k.)e�[����ښ�Up�G��ʔU��n��J�w�ǎ�(��by,l�Q��,Ռc*��]x��T:��2���,�V`D�u�57��e�����m�m\ٕ��˽�U�'U�9X���n�]�lg^�'H4	�N�ϸU�J(�gt�������k�I��7zc����.3��-W�`pc��;ȧ՘�����P%�b�o_��s��\¦�e��}p���_��5�3�WU˔�b�)u�2�<��r���o}�\H��f�5§o[|M�������*�  ��������$J�l@x�I�����6��AYcN�wB�A��z�$�Vo�:��m�>��IN�:�4�ƙҥ��3�}�a%p���z^U�b��-]���c0�a��R��{�C!j��!Vp�3��o@��k�0urik~��DԘ�
����n�<�4��7.�͊��tV��f�u��D��L�y\	K���z$ �}}۴��[oué��\�D����Ж���W�nڜ\�V��H�ݡ�M2Hܚ��C|y�@��潑l�B�q�D+���B�N˄n��o����r���S���h1�<8ðbf��|���ܬ-�4��p�i1@X����F�oUby�vHF�a�q7ӊ�]�-�?9ٳ�[��R�!y�˥�m�5t�m97�aǁ|�:=}�m�8�~Y�y@<B$ѩЄc��k�,�N^�:#��3$9�����=�e���:��+6n�Q%܅���OD��lΚ�|����`��%�;�e�mͶ`[V�XܩDK��H�xF�-tH��}BJwàm��Dl�Su)�ŮR�L����jUw�ո`m�'zb�ǉN��G�]�^A.V�OF��{k$�{�_+P�<�ͻSnmG���t���D�@��`y�Զ��8Q5�qn����RW�j��MN�O 7��Nz��^VW�����j��d%=\E��S�3.�:�0r�rl�`��Ҽ�膼`���ʿ]_�#�ufzV\� Q;��W8U��\��,ԝ)n*Z�3�[&�T+���Oٛ�����ӧ�"V��2n8�[��}zḓ�Н���9��Ѝ��ֲ,��3s�vM�	��q���n��
��f�gU����G4�S���:I��Wa`4#�����ؚr��:Z��s-�EE�����Q��e�w!ܹH<ԫO�����o��%9F|�eyE}ys�`�r��n�H�Gt�y�tE���PHr���L-p�䘢����+kQ�q���_`��y<����59�lֶt]�؈ݑ4풖���j�*l�mV�}���V���gL9��	#M�&(��|F<,�t9>]'c�f��M=v;F.�`���p3r��T��MĲ7�F\��bw}�çi���y�ӽ;�m���Q�*��V�Ӌ��:�3� ���Ͳ���ʹg�,	��8k��D���Y��qJ�T޷�-p�󽫱j��h���$í��g2�##�S�m�id�����X�y��u�7��K����ޛt�%��槏t�p�v�a�d��9�b+p��u�6���Z�vØYݴ�E��Zf
�A��$3�ήضh.��<j�q��bf*¯u`ig8�X����s#��nF�@�Z�UrQ�x"��e.�^�j׸�op�}����ʾ��P�u�XM�D�ث̨��*^;)�{�[�T�)�y���Ű3�Q�v��r��]�q�O4��gU�3c�N�1qL�{��'j����5�@���/��d���;y��|S-��,><�����Vy�J�y�ݫ����ǁ����N�6լqRX��n¹�{�7\�#G&��`Գ-O���å�<����Ǜ���AL���z1Ǌ�J2�@��w��r�P��.Ye6�ukXq^��l�uajA�oY2�ݎif,j��_t#&4�[��Ѿ?J|��wQ�cڲ4��d����l��Hx2o���P�\��vP)
�%H��:�b��J�ļ$^\�r�����vcB���ǉj��)��/2�tС��	/w\�U62��Ь��X*-��}�kz>�� �J�r�9c25{�;�r99H/j��綰��+BA<MSȻ�oX� T�C���l�gH�.�_}��}m&�OM���`=�'���>r�tj��(>c�~`��|������t�_h�C�S�M|{{o @1>C�?��A�)/Ȁ!�AT�aCب!��tI^{?�������w��"�}����{�����A|=��~��{����O���4<��Q/p�������J ����h�I��4F���̻����֋��f�yZ8�q�+�c��s��c��u��kV;�7�mχeK�S-��0cx�]W�����,�Cu��o{B
��\�sYZSؚ�o-Ü�� �;|{�3rY ��je����29���vT������]�&w�U,�5��&�g	�D�#O�^eAd_
Z�-���̬��لǝ%�� v2�q�\jL
��s��&����hk��vs����#�R��9�v꘏Ay�=��r1�W�z���O\��ؽ��F�v/�æf� ))�PY������.{f�U�\fMY�%[��1v�m�\0$�4a֬�˥�ko�c\Хa�d�<5����d������m�����k�6Km1FP)�p��s6>�.�L�-GZv��`}��ॕc�g\�D�e�:�%B'|L����9���S�ѽ�F���ی�lK��C%
�ɗ�5�IVj<A`�rh�)��)]���s�BL�F�tҤXs��!jZn�;��tI��5]�74�<���Tƚ��Q���Y�����F�;e,4�WiUs)l��NB�LX�� ��f6��E齼�������p��{�H-vp�t�:��-�O���sb�ބ]�P���Qe�5#Wv�bki]�>�%�#(^��ac��8Qk��e�	23�ǉZ������+��X�YI�e��g7_N��n���5��`��2���"��e���Pv�k�z�P_Ȧ:RT_nu4t�C�hF
o�i���0V��)��"C��R�ŧG�[i4H��+�TjI�bc��/)܇0��ku͑�K�`�\��Z�T˳u$�{Ӱ>��8��Lp���!�M��<]�cU'�IۖC'u�����JBgc���k9�8��Z�z������O\�v�N�7()Vf.�	��]�7�����X}�"���g2�N��:��3��iR��������y�������N�Ќۈc����df��AW��%���ո�9iL���~:�+6��`�{�Z��8�7Y�6Q��U�eTȂ��6o��Էo���L�`��g�4�:�H��HX� V�a���f�-�w��\gsɵ��̶��7�2����Y�C��vuE.��nI�7LTQZ���r���$͒��a51��T��ACZ�<����!�s"uNً�ev�7���ќ�����Lf�t��.����hM[�҇�Y��ڢY�s�Jn��t���/����2�otTp�Ooi�<��Q@0�Ų]vi�Ig��5�5-�JsZ�Z��dh��%�D�39w۪e#v�|�����Cf������v��c��7hJ��&�6(�槽JLֲ�D[SG+��8���0�*�86���W��+�G�U�Ri1���/E��`F�Z!�������ՑB�ƜV�Q\��Z�8�}+��b��sf��,:�~&�xv#�b��E\�^��Xѫ�fXRh���$=tګ�Q��1+�Dt��o~����ꂍuG�4NgH��f]�]|e���n��u֮u�NH��l�#諪t�Z_��Un(茣C-4�q�xi����u\&8L�9����7����*�"�yո1���8Y�����B.ǔp��V�rs�<��h����@�#̘���U�WԲ�����ƂY���7.VB�SI����˾��\��err�$.i&���} ����G+-u�p=��n�%V=�����,�݉1{�S����ʀ�>q�n�`xh�lW{ɒ�{k�ͼp����DKS;�9d��y��[u��͞�J�AvKF#�`4,�V�\�:@�B_�ѷK1"�K$�N\�0���ZP,
G|N�Yg�u�@���k x�p��VP3v���P�����}�.��엝���"���$˂^��jm���L� �:ȝ)W��/(�@��`Zr���kq+h\�����'D%'��[�xE{E��h���<`o#<�]j�Vr���V6���b����l�a��t�Wh;��q^�Ea	CQ����@Cx̫�3�,�yvAl^�P�׵��\�^�-��eŚ���{-���*i���V<E���$�G���J���%>�dkB;Y|M(�� O`N�Ԙ[[��m���dE��.���œ7��ja:D-�{S��^ُn�u�tb����M�VFҲ�tۜ�.�d�lӕsyco��F�j�\�OR:��<��Hh]$n�'����s��uQ�e�t�ki�|���c���ފ[+R�ɢ���ʊl���]�45�e��:	���U��<�8��`�H�}��OO�G��������J��[xBg�N���o:t��K�h��wT�k�$�㶇����6Ƚ:�P�r���U}]������O���J�7˟i}3�n4";@�Ø��0*��s����o�A���<{Z�$Գ]��}��c##;*_�Xa��1�R����3�.�\�b��2클��@h�92�^�̫3b�d�pFqw�X���l�!�5�Y�s����"�k�Q��r٠p��e�f�cKV"j��3�m��VN��7B����<XOm��}R��v����l�,�mpoo�!{���M��P��W63m����]J��
�����N޽d�,�Cn��8ILM��/�XWr�R��t����j⣻-�lan�H�$�L���X�*��<�Xe�J7�!�s�K��f��0��Z�LzIi���5�2bÖ�ß�������|�N���eU� U��_Y5�����k�$c\�k��.�&{eC/������-���QC���<U�ܬ��Ԇ�t�[�F��n��������"u���E�ϫr��8�����WN�k'��z&����(k����J8�F��S�hu�{���FV�0sg��Y��Ω�Р�7vf�6�7��7n�U����L9�[Q��z��/p�،�c	 �k�6��ʬ3N��,&���7�@����ь�p��=5C`�y~�Svw~�[|o�%�dyF���.�X�:�,��kV��Ll��*v�'^&G���^���m�Ȱ�9S*Jˣ�Y󗉹��o32��N��������E�YR��*��uMD���դ�!��Bn��-w+���9n�F���ڗ����̐^i�b'���Z�"�Zom����]�Gt�&Ӥn�W4RΣB���e�UrUƻ0$i��2A�z��;�G��P^ɹ(T;�s�th���jZ=xv�o`2[�����BwDɎ�q���D�Ri�J]L���/�e�� L<��4�e���9�a11��bb�:[N*�xr��I��"��,%�k뛼� �;��׌��ڸ��'Y�a�)[�3����*tZ,�b7����U(:�M���V�E��t��])F��͔RH�7Uޚ�p���6վ5�HT*����'���T��v���ŵ���`�؎lӼ���\�m����	�^ڮ���ts�6�oKB��=�4�_h�΁��k+�p�]!�ʞ��E�k$�sI���[�C�˳���檫���=v�ٕӛpR�1�]9i.�!tk*�n��y��O�%���>OoV��!�1o�_h�C��3J��{��`���2�;5aKXC���ᖊ����@�wB�L,�6U�<��,�v����L�w�;��7�6��)�wj�R����J�;��j�]Ǜ�U�`�04���+~���g�rI�Nl�q��SSL�L�w�譅����ˤV�WsL����W�&�vQ����4���f����ö�unJ�cN݈\���U����^4s�_;}��"2���Xӛ�dd*���T�`���ӷ%I�JB�N㎙)�'�4�N8�g�8 {s�$;5I-�
��	�4�{�$��K�_> � ��_��;q�mi��O�����&�`f
v~�����,�8�K�,��U�vJ�2��p�\֓8d
ح�S��P�� ��U��ܷw����c�k߉fm�-	\�}zФ3����f�����U�c����8�#놑)�t�{�b�p�ޭs��*QNښ�R�=;72ɱ�n2S[�V-�B�8�K�z�����E��DL8*^��A/��Ӏ�����˗zNX߃�*{�㽎=�AT��fJ���Y��2&n�1�O>�j�O4h�S<��4P�F��7��qdt�+. �,x�+z��Wh� �B�+�S(GG��e>�ئ�j4���e.;;�5CVU�)���]��K{CG:������R�����,�Η��]�k��+��:����&����c"R^Ҿ��'vQ�p٘��殯6����G�mB2�b�p�qі�"�����''��6�Y�Ox���w��s*�4�l�Vw(�>����I�&�xv�^�Qi��9ML��$���.�c5�ٴr����q�AT���Rk�Y��������v�r�^.ͧb�p垂p�mT_d������FE�	��~I�g#��{^T{5h\�ݞ2�Y\�9-P[:�x[ʰ�x�R� �E,]�WB7E��5V��-����vfD��IZ��s%1%�j�۳k'Rz��]��t���U�Y��%#�8E�i���͇�"�]��Y,�ݶdf�Wr����*wv �P?�r�`N9K�]��������\j�w(��w}wv���W�[�Z��m����XD�u��;���ǽ#�Y�1��κ�A�3��䄹�d�s&�O���yX.��;2[�o+tվ�����w�}�(ɰo]m�\�q`�G�.�-��iө[/�+�kt�is�'=C4
]a��b���ۦ�4j���0mȧ
D��;[�c��ť� T���uy2B��BN}�ek1+��|���9�Xuԙ��:�J��\���QIrb�O ��z���B�sd�+m��յ�5�9q����>���6ڻ�{()�¿��)7�q���*^q��$����%Hs�b����7��m9�w�@%=X���Y�{p���e���ǈ�d.i����$�����74�m��+�ˬ�L��R�B���uN����Y*�mR�lNuo���m�q��[�m^:m�����;;�|�59t�T���뷊Z����o�ӬR>��9�Gkun���2�Qan��KדZv,��cOr�bsfGmwwY��J�hB�O^�YzoE���#�)�a5l%ݧ��Y�L(���[ǘ�Q�Zi���3Tg+&XoyP���X�1���\�Y�.ã+ql|p"Y�b��t�X�K�Ƀ+n�;�Ͷ�kD����tT��,�a\�ptI�A��Hݼxԩ�\�T��YA��j�v�=ewl�]o���p�"���Y]ar�Y�^W i�Q[�Yb4��꾾5���]7���~�K�XҼ�e�ubU��"�h%3K�%�p���/"��n�nkٶ����G�P=P_os�*$E����87Y��`�v�떗�Vn��et�� V�|ys���|)�Ző�4��y_D�#�8;�pVh��{lq�v���j���mj�8�n�WK�	LG�����5od��e�sFA��XJ+���:�4�Iҷ(�2���v(-Y�ѻ�6�t�C3������Ú����AYc�$EeI��#[�LT���s�j�N�L�xsi5[m%x��sc�s�}��T�����}�}y��3�v�)�i�U�7��݊	�WѺjμ���y�Lhy1����d;nކ2��K�k�bf5�Q{�vڨ+���ӧH���������n��26�}-D��IK%^L����ct\Η`WJ�Q���3��͋��q]�kU�!ե�Y���jK�Vv�����ue��^��S���α|�F~M..�n¤aQw%�h��+��r�\�b��z�L՗vX��@�-�U�g[#��w�&�kd�7A`����a��^KX�X�*����I����2�Y�aO��j�5wt����Ө���.��Mu����{g�����f����Ā� �R�i��n��.Ң��vl�_]�;�Ν3��z*BN)����P��[]AF`�\.L�)��'7>e_V@�����v("�>m&���Z�ܬ3�mk}��s#Yi��q��ZtbTt��$��nkl�-�`�֍c�!�kB�m�˕e���(�pЈ�����p��Am[,.�^9O��ΓM��uW	ur�#ʮ]w.1�E�kv�ʸÄN��Rq�8���9̗6��΍�����4��7�x�,���1*��go���k�i��V�N'�e�5p�M��L��غ���G�(�w�$�����A�V�\�jOU3�G��nP���IP�Z�7���x�aq�*~̌(f��ۅGi��x���!��=��&u�ik,�z&Et�`�0���UmJ�۩˩
"^K�y�¥�*e���"w����l3�$n�YM�2��/�Z�.�YWozll���
6(��D�9��	:���ʆfG9�� �T��+W�^�Ep�ܼ��ױ�)��y� u�
��5�a��\�Ÿ�E9�5u�0��!;��E��.Ms��RtΛ4�P��.m^�r�9��1��k.�Â�iB`�H��Oft\�o�����;}-��YJ�Ֆ����B[g���d����[�ڏx�4���ӄ����>��hd'����-��	���7��mJA�̹K�T�<=�kٽ��I����x����݇"�9��U�&�A�E�JF�Ū�}]��̻:[�9��C([�S�ڬ]��zU�ʲ�.�.XK�:�I��,�:� �_�7"����RV=������� *�tϿ��?�������o��L�O�����>>>>?�����38���q���>|<��wF�-u���[��8��^]h�$m��&FT�R2
(B�*��'�B�Rn&YIG'��`��U?��ն��?�������� �&~�C���m%]aʊ���}��pҸk�	���lD�r�Gd�l_"ʤ���[k�֮�Z�tc����cQd������x�N��F�c��yn�Gr�ڽ����I�5[�S�0 O%ٍT���W�s�u�q��X7\I9{N`���I����>�8f��I�Gom�UÁ8��ڱ�6�&�I�� ������W�;hu
=��8��#��ϨF�ђZX.]@R.�̗���'02��iˀ;�R���3����xY��u*��mDoWu��Y��
C�TGJ�#��Ǚ�o6�ؖN�x��mF�J���\��ɂp�OX���|�����WNr�ũ�e�(@���Y*�n��j���|/�h��Џ'�j�(�h�K%Ha����޳|7*^26<�N'0�V`��%�rpq ��ۙ9n�Y!h:�>�l�ؙ����W��o_u'���+L�]��d�v+8�&�KR��K�(����\L�Y%#\�o$Y
��={�ܻ�Ŗ�]$�Z�՜F֒%�4;�c�d�NH�w-�wp�齧����+%}W��ա�:4�^� ���Ōn_S�����.���ԓb麂��p�:���qK�#����}E���m��)1��#�?Ĉ����IB8D�aAHc14Bh�"()$� �)��D�P �L�"j$cB���[^wm�^yw�E�;�i��W1�4!�*~O��L2�(� Q6�$�$��N~�A������Z��^xn�q���{�F+���SDCC��Sl�{�t�S����-���z�B��(������"
(���:�(
M�;���P�EF&�
Pw`��(���F���:�l�$(b��*�K���� �z�l�q�AьlI�RDPR�:(8������Ѧ��%&�R�[����Q]i)Ѣ��P݃CA��&&#�Sl�q�3h(�z**]E�x��$"���tTVڂ�!����|�8��lݸ�J�������b�(4h��)�]tm��LA��4h�4hi�@m���.���j��Rj����b����t=t/v1=ڃ�)(�@u����ɻw[�ڽ�R
�B쿨��\�՜�'Ay���y/l���7�;���/���@}�1���b�: �Ek�*9��s���%[��-a��%�H8{yP�YT
����P
޼�%q�+4�p���Ќ�z�7�ݓ�e�����詁1&oL������#zZS�\�9y]Q��j�eg��X�ͺ�'���2��q�;�яa+:�\{oc�h���U�u��gu�{���_�\���EG޸���es�����ޞ=@��a�ܦn�g^�Q�����ͻy�D������0k������q{*>�F	�܇6UF|�����d��U4��֏����������{������T�������|�3�Ok=�Ŷ&U姌d4N�����n�9�lg`��֏m���:x�q�y;����c3���D˳�iЯHt�b���`Wq�9T�%��T��A�s<wN[���M�']�FH����A��O��u+יg����9��8~Ú�n���W�}�u|����_���\�i�G{�_h���0�����5Jɼ�ҷ՘h�E�9��th�3���<k��.m���]�o����� d̓���8N�'U��œe�vʋ�t�O��3w��g{#�����.�κ�7�����C��>���~��9�9t�=���4ϘM�q�{-�a��u]�}���&�5��8hB�S!~��ue{���yK��^��e$f�r���ު������g��ED{|i�A]����}Yߵ>eo�"f ��C|�����8��n	S�Փ�,�����}c����
o�gW�����|����!Y��6���k����,��c��˾ڳ�����c�W��x�_#�~�+Z��s��z�wV���z�xڅ���s�Lr�=P޳T>�����E��zB�V�����o��ݢ0Ӷ�p�<�d��t�y'�u}��瘵ߋb��*i��~�>\�q�p��~������w�S9�N�O/k��W�#ک�~Gy_��wn��}b3�V���7�-�x8��{�������Ѽ����R��sW�D�
6�L��#���}il˱�/�r��#���,���S/viv�=E,��v�a*�]�I��V���#|�r�왖䕜7���4'9�P �5�Ѥ3�mlr�;���Su»U��9H��oYe7Y�Vf	�E�֠WwD�h�����������+5�7�+�ʟ>볛�s��Ƙ�f_�h9� ������dA�2��y�}c���S�)��.~�'��������'��@���}�ƶ/d��Je]7�9��U�A8�!^�C]w��}���[~�P�=���z�Y�4��g�}p�?J�%��6oeC^�z=�9_�o���<k|�L��{|�O(u
�N���W��'��w��w<�u�#r�\�O�����{�����;��E��4��CV��_V�4{ۺ}�����9sSu���G�T!��4�j#�������;�k��������s��"����j�N��Y^����u<�o~+��0�؃�i���s����:R�@��[�Tc�vw��o��Md����n�y=��4�[[��@ѝ�bt�9}3����2v�x����h<��s��Ҝص�Ft�b��m�ɮ\�9��0�/0��l�Q�9��B�v}�[|4����F�oJ0N���w�X�m����봣�N�z�^��и��QR�����¶gP�Y1�+:���Y�ɰ7�ʋ��+wg���*C�V��z����{`��`W9]�>q�op3ծvEe[͜h���Ne�o�&x׉ⶭ�a�p�3~f����9��-.wZ,��s��q���o�a���t��~^�S��}����Xs/�K�O�'&����;G<�em^��Hng���ܮ�����[|��o�{%�{M�.�����v�a���ߝ�G���x@�'�9���������<.����旤\��?7Ư���5�����ǧ[Jx��gz��wV�[X�oL�x��ѩ�"<����1~c�J�{s"u��ϟ��]�ޘ~�����>룴	�&���[,�gn�~L�ơ^�r��;]m��Y~��BK��޻�ܠ�Ǝ�h&�Aֶ��|�U[�}P����Y��oȿ}��4�`n���|���^{�O���|�NN����R�g�|���y�
J4Yə
��v�K4^or���)r��'`=�v�N�8\����	������y-�<}:ۥ5D�'r���̎�sI��,���R��HJ*d�;su���y���(#�fJ�J
�f��US�/h)B2�w��M���M즞M\z~?T�!9Ń���gL��|���^T�9�f{d��vL�ݾ�=��暑A��/g��eV.��{�ͽT���K��j�
J{�_H�;v�[�I��3��_�sk)���5~Ϲ�� �%��뽸2a"v�轐�%�q����f�ϰ�t���ϰ�Mtx���j�e����{�=�y�]?]"�{�s&2�v/{Պ��Z��g|��c�TW����Ν�d����#s���}���[c3�z&�56F����
bru-�a���L�x����'��k��a�i�@'ũ��`��ك�j�p�g=�����G%8婗����K��YB�;��½�k_/�n�z��n�������g���Y��.�X�zB�`���к�����>�����]xU=�:��\ó��}����<T��{���v��*�붫���eL������[�X�g7Q��*��^��ku�පлr���n��%#�mc��;��q��Q>��o���}F�8M��S^f����ٻ���w1��>θ�+ew�Gڳ�l�n���N��_Sװǖ6S�P���{�m�gt��־��!>�K��uy�O������[��FW���0`(^��`�̸Ȝ_�S�:�=�5�����~�	=8y������ �R����:�k�b�Lx��[������|q.�*�{�׹<*@��zMh=�{o�z�^��}������~{_M%��,�L���<��]�v%]{��V�uXښ����s)����IAr�zvS�~���6�Q#���ߖy���Y�N��/\��G�jsk!�pЏ��*�3���IJ���.����.���������1'�E�^\�O���=�8�t�5�<F�A8�U�ʋ�>�{{�{����~��#����?<��3ۗ@l{��b��W�b�������Yx��y��'�^z,ST��@*��G�3���]dO#r�L�����ͣV���H+xyA�p� ���̽Z5��䪿h<�n�_h�@�r�Lˀ ���9z�X}�cT�u�B�y.�2��v�`�5��&-P.������K� ��M<� XB�@��ɎI�������U���+��@�=e��εӣf��FD�V�Yަ�� <��C�.{MP����]��g�ї�����:]׫=��Ρ�|��gzE= �u�6٫�/M�^�3]�Ϯ�K�g���xi�t������Y��M�q���ho�oS[��6�G�1T��d7�}�����=3�骧��/{�Rn�D{�Y1c��ӽ^�s<zSV.�xEx=\�Wjwx��*zzy��a=����v�k;Mv�4�����}��<>#ڨ����n��3|C�����"�pt0��!��s=�c�~�+��B�]^P[o���8(���}�����)��E[/شG�3��t�{o>��^�Wi*��<�y�Y��h�/�ب��4k�Nd��m���O��1�����\W����de
��v~���sm#���Q �W917�dǟ�y���O��g����^��AV�ݏ�T�{��oi���4{R�d6���s;Y���)���a��B�A��+.���O)�=u�+w����9-�3��ΰ�sƅ�V�u�挃#�@��Q�ɆEN�EX��M�ҶSʀs2��TuݴV��e�'y;blF-��s�!=�������>�����~��j����w<k������2>�d��9�-�����67��/P����5��R�M�����W�mwS��yP��N�<ɬ��x�r��A6ъ�/�^�d*�7�ku�|���#���npg��I�'����f��x�	ދۣ<��uG~���[��U��������H�K��7�<��p�7Π��,o�&6�)��Z4�������<��1	B��;n�x�FNP&�4�e�w���E�H|�!��;b��=�h(����iVvs�l�';�d�Y��s&���
j��ȳ��ǣ���P�޿`y����
�I�s=}�zM�jdO��h���ݷ�����g�Yʾ���W�JVUtϬ������$I�ak��-���k�cj~�<�x=�Q����?VJl�y����+�Q�>�G0n���zm�F�bL�f�F�5��͚孊èn7��	(�����Taj�ù�{���W)y H�C��g]>�R�y0T�3e#��jX�s��9���������^�ɻF�f�U�WL���G�;ʲ>
+J��8�J���k*{�۾�A�{�?.�,�
��{`~��m��]>�V�o�3�Ixn�\�|������Ǖ��9Z,/�� �7��M?Ez㒲��7F��:�{�Cx��5����}>�[5>s��xް��<s`�k֨U����b�j����R9=�q�1��'��|����Q��۩�?e
B�.���R�t��~r�Iŷ'ye?z��>��޿4��gj�4<~t��7�0��F����&{FW�L">�ٶ%u�;���kQl%�M&��yga��)���3��TVw�]b�=�EǢI��OL�7��.FH�,E�2i��a�σ�C_�U��M���&2�D���X�9�WVg2�t�����4��m� �OnphgF󽊝bd�b;=Ğ�8ԃ�}�Z������x��oW���b�y���o�H{�����ȋn��:�M����ږ�{��WK�/�S���"�9҅p]���9��7C[6aQN~F�ؽ�wgDΥv���Z'��EKM�A�[#VMŕ|w�X���^lwy��vWke���S̎�V�(�0ӱZ��2g]8�s/���h盅4	Gj��If�r�	V�D ��������^�@�T�-Ϸ�n�(�.D0���E�ݬ�9߇�}RM�l�������5k��޸�u���a �0o���&�N.A�s7\j�n�sg"Mt�1w4+��o��|q}�Dkg�P=W��)y�c�ho�u.�6~��uZ�c~�羉�2\Ѱ��^,��f`Q[��uJo;�[��s����ۅ��6�{�E�zP��4��gګكt�U�����ɗ��l�=~���HF�����+��y�z8��2hC�>�I`��	����:������6��FY�_A1^8��5fg%�i�p7<}y��Qv+���u��O���_��]i�n�}��7Vܸ�@k�@�*�BLl���ǋ���|�V������.���`��~ik{��O����c�Ϥ}g��q�\����,�pG>����{}>�o�����}������y��<�`��Çu�x�e�M��v��o6Ѻ�
���h:�Gd��;:�n�ʕ��J��o&�]��U�<�<Ղ�C�z�Ǔ6��\�X50 ��bL7�w^�֝1p�[������(Y��Y2;,`sӼ�QmS��с���+��`�5o��7|��\���mot�{B�Ɛ_c��V�]�gi�{;��� ;3dxQÆ�i�P���9ÏL��rv�-"��f&٤�եr\��#0���E�"���R�0Z̥D�FA����KZ���,�F6�զBM.zZ;Xok��o-������׍V�T�fd���� ��=�� r��<s(i����w�Sn��}��7��P�{�jT���k���;D���U��f�#snܕ�� /�u:3��Y�Ȱ�4��Ed�F~��ޠq�>�����c��5�8L'b��gj��q�����.R�^,�5E��-�6��k�˵���u��rݧ%k$�J�܏��b?M������ [��Z�}��s�ṧ�k3hT��9�-LC�P!yl���`�\��t�g��S"�jcP�� �R�*g֔2�ʻwo4��SI��_G�]��.sH�6X�ӟ�SM
�9�;W�k���:q�ʹy�M%�e�M�y%�=����J��\�%�}��2��Vo�\܂M]�p��i�3��2m/-�hRXm���_�و���~�@N�}e�{�0�-g���N��+(�U�Rk� �j!u���D{�+�g�����\#�y~��/�V������]��Limki���Y��[���fC����F:�Vh�\��3�F���pV�f��;&-[�39�=	L���=��0�R��y+^/�>�"�GZKu|RSk��^�e�2v�7:P��Xո�̾V����}��m�}t�m������S��>SK��D�9Y6�e3�)�P�P#�H�`�6�R��Y¨h��F�&�rpɯ�h���k�N��T���g*��%𺋷u�C:�
��:�jeAZi�>�5B�:�x��΅@�AB�[�o�m��(��R��m����Qs:�AD����D��ql�����cw���
ۉ#�U����T�U\���GX�Σ��[���K��;��J��*�ah�u8���fu]����UO��M�{MA�ag�V���y����:v�p3q幍��u/��s��u����H�Zm��&�N+�@TH�7w*���m՛!D��0fF�}�;�q��M��Gg<=��F�/Z�k�ܜ�V��y^�ͺ�J*;�����U�ukX�.���b����rd�ל� ��u!�'A�(��a���/����c���9���^���ڧ�:�31�vo��z������<r��}�q�Je�p5˳]�kb��	�������`I�Ps�Y�E��It��:=�b��f�c�w-��R�̮Q�-�_N��p2�n�����Hy���6N���ͤ������ϑ�Ѷ���>�ʃ1��/Z7�����>F�m�[D2y�C\lQ����'n���Dl�sѶ������hb���#A���O�0�͢���qy����������G�������c�9�y�g�ۍ'C��y�C���b�<�û˭Elh�h(�g�G^y��ll��t:���=!���������i���#=i�m�ѝ�F3�����#��v�Gws���Uݥ�yǛxOZM��瘈�zk������g�Z.��<�v�Ǒ�w��V���3��q� �����Ɩ�`��Ū)�\vMQvMA�b����m��7����q�g^lQqj�eӤ�O��'�&h��#q�v��=���v0F-G]p4�S^yn��|$�1��[U6�=[j�)v�kF;�cEQv��U�)u�늺ד��UC�t7wQl]���j��nŞ��ku�c]wb�J��#�}3���~��ͬf��.<�~aFB����e��ω�W����9]�B=<6�vZ�ݒ���~�����`��%߄���C�����3��NȰ`��@�5 �(�#�{�%	���۩�:�Y{ϋ"��ሐ3�;n{���<��G��M��z3u	��	>DAe��s׾G=��v[$� �p:G�$J�β�>-3*����v�JPm�R���oz-��9��2�1D���[���f�p?��4�"q}Nه�I��:�X�_=t�Wޠ>bD}�)܉���z�rt�����ɫ*#}�DS�Y3)��|��3����D]�y[�q�.��ۇ�����O������>�,�k�
d|�V̷P2�]�T�<5�8ta��¨�!�����6U�=�'-q���\mn@3��;z������<��P%��J@�{�;����)���,��<b��d��v�y7/�������=C|c���\[�Tu�zO�uP��U�5���z5V�e��{��twW��(A����3��y<gRV�7t/�0�(����� �s�/ə�k����p��3�[[��ʁ������(j��>*��p���b�o�{ΤN��S�n#���|�9}�r ��Eٲ��0��Y������:��.T��1Q���캌���hŜ�a\-]K�i�p�m�ߩ�D{BB�݋�⎳�i=X�l�,ߔ�u+͢�Nͣ+p�#��)ʕ�3��K4�'��Vb�J��#�þ���w}�|b����y�E���Lwxg���[ З�;���?��>��B؁��u��2e����:�����fŅq��;�x���q+��������G���2/+�n�bXgf����P�^ 3�wC%*c�P	��[<О���\�;;��� 4�D�x���WI��"��o�Te#j��6-�Z��u�h��|+�u	��Mw���?�A�=���
(�:��J��X���_A�LD*��=�Q���e�1�o[?����q6��N�jV$�^�ǐ��yw�ɂi`/0�j�A�|}�d'3��ouq|w�\�T�����9�ʶ]��,�����>��s�st@|��(��I���DL���oLL����G�>47bq�L��;>	��g>��Q��6�p�L�m{��	��]"�兩�\������?�d�����.��ȥ���L�ec��1P���fޅ��e�����ޑ,h~���Ϲ��Ή�����Sk�S����jՇ�d���LS�� .{�@=7�^8��V{��� �Tɬٹ,}_���/-׮�I��[��IeȞle�~-�)����tY��K���UXN�����#}oi�cnp���si4K�����z��:�q��%��8���v��ʴw%�c��s9�
��W\��yX\�i&t�=}�I�ɽ;�g�R�B����|�S���(Ɉ;��::�{)xh����r��r�턫uŷ��5b�E��s�d]��^5��C�rH~Bl}1��Ql�r̤M��� [#�����>ߊ�.k���\<hn��'9t����r��}��m�W�-��f0��X�^���
�$z�9�T|���W�bF��R3#��G���L��<���g(m	3}1\��oA7� ���T^�a/w�z�2h�S��ym58�p^��>��TǙ��0�:9��8�Q��H7.ᱻMҕ���I�q�������F�h������2e����$`�-ѭ����>�r�V"$��x��������k+eZ�6�!�ܰL���@�E���
����=�,�[=�/���z.�������(���7k�L)�Dxp�Hؗ`�A��}Nj��Lv�oP$�����C�|nmn�+,|펏�i��}�����DƴL�����^<�g��	Z�=c*�1�&�sQ�7����ƽ|hE���~4yf���p�6k���,S=`y�{T�:�2>�	Bt� ,��������up�dF�^�3�,�e-��X��3������x��W�8;+�ɽ�O[2�Seؙ��u�I��:��ԺNR�[S��Ғ�"���r�v��:jGO�F���|��|o#ߤ�����R�>�����ۜnk9�e�9�`����֏#��`��[�/5,��T�|���3��;����{�Tgx�[I�Ҩ�CNh>S?l��d40�U�ÝMTd�'{�;�,κp��c�_�c�����m� X¦�4�UbY�'K؉���G�V"����hjȫ��X!l��5 Zȱ��s[@�hl��0�:�9	t
./e�ѫ�/�^���Wvܽ^#<�����W��%�Tc��T�)�3��џs�bS�����B������ʍI�gws�a�q��d�x�pQ6,�����<�2k�
_s��_[��'kjnE3�����2��Z��w"pZʈy��}O^��y���!�v�
A�4���.Gi�4ll2 �c"�V��-�5L���۪�V0�TfL
��W��;f	��s�3���wu޻ղ�u���[A�Q/a�NyAa�T�݉U�թ ����w�,)��f�[��Ӡ������e�#��+�&�6G4��+��6�ڗ�JJvO$�zto9�� ߑ�ўw[���Hs�F�)�d����s�\F�̚��#��b����A.�R;\�y]w;�x4}^U��v�{^�4p.�c���1T�il�hæd[w�4��Y��w�(T��i�y�b���w2�h5�[ݫ�i�Z�7߱���H:��]srD�r"^�|�r}pg4Z�9cZys+,x#����"K�D��o�[9���^�2����< �)VՈ���&"oLCn{ۚ��3k��\�*ڟG�xۃ.��c�Y��zx{Bh�~��DƂ�t
��*N_C����V'�2�jQ�hO=�O��*���ݷ�\\�ܥ4e�>f�fq�Kd�ui�?1�Dh~2Ct#BK�>2�����T��n���u"t�'�w��QSװt��_��T-x������9a=vy�_�3]��P�O���̸H�I�*��hD�dckS�_;�=C��x:�tf�,��<c8��{��M.���	+]0���V1y}��!���ӱ��o!�QI���%lb�вoNS�t&�w���q��� �@�2�\��MF1�>�f^]�_���m%(6欴�Dv�l����g5�Kfả��{��0�����p_�,�{�t���E�X�O]/�E\��P�쭚�|�l��^�f[t�ң�z�nv���735��<�P��Q��}����'+��0t�]ykj�b�4�	r��{΂5Q!���!��DE�k��#p�s8��+�F7���(ų�Om�^gr��m�mˍ�����a��:�`Zf�U�Z�W/�u�V�`��p]��x߼/�"Ē��{�& ){��'��M^L�>�x��lD�.p*�0��s�֮�(Gb��m���qM�yn<�+Z���v�FL[O���jG�t������t�3�;ҙ|s\�z�B�n��:�/^͇�U��i���l�x�jCf߱��g	���'�L_:�����Ru������j����� ��Ud�H�[����)�=� [�/�l������;�Oӄ3��f����M��k���������=L̎�5T���hT�'�{��rn������З��B\��&K|d���jD�b~wC�)���f���Q��?=�_*u���Q�1����/�Q����Vqw���19�Iv�[�����ۦ6� &��2C���^	D❬$�_L�	.xAg�4�=��хS]�?w9�|�C��i�8Ȫ�L6�O3��kg�t3\���8�4���=S(�p����&{pQY��S��3�j��Xb��Q���4:˙����*�cP��(I�׮1a��H�>���u�<bH0x�P_W	��s��=ܰ�#vGPc��,3�#�y(��K Ƒ����}�W�.���io��E?@�^r���p�N���}^�;��0����a�љ�uj�)��m���+pq�q�B�2Q�Л��V�-��v1z,kΈr�B��&b�!��<���]�yu���a
�q���v+K-cY�,��ʳ�_e�4^^��`6�����5�bf-�Vr�[%z�-Y����)X%m8��f���ީݢ �(���(��I}ބ�0{�x��7E�������ؚ�=����럁T>3d��V�:�K��_WW{��2vS�b��K�N'��TA����k��jMi�~��Y^g��y"����m��uf,b1��R��/gо>�7.(�QB�ϫ$��W&EG)8|O�7lW�%)z�p�"��;,C���ݡHDn\�Q�r�T@�����#���k��Cx�m�5�Q�*d�O��eIj�;��vgܮY_�tu@=g�=4JN|�I���U�8'�X|q�gz1��\�gM����ta�5�9�ohȗ�u���m�.S8#ٛ�W���X�2Z�ʢڡ�x�33®�jMh�Iט����Ꝙ�g{^��e��%�i|��~a��u�F��8�fۛ��|�WM�%U���jF�3�ΧX�2���S�G,m�L�#�\r�~M�|~�ρ�Jf�nu��[�ܑ[x�f���9��y>Ӧ�[0a1N�`�D7G7:w�f�x� �=�<��T(���;��{i�� ��Ǝ|��'�v8�x�	7j���y�e���X@̇�|n�gg���B\@�.�U5��k�؜;�t3�qޯO5�����1�I��`�Y6上����ORW�h97,|��\�h��n��\4�hN�}0v�x��k[���j��5t�)��K_s9]�Ѻ���V�l��M��H�>�2���a�q��h�3z}o�fٚ�w�	����F�\[[����^q��T�q��j՘�p)���xO§�ftX���7����~�(��A���cCx�X缪G�/]:?@�:�x�R;�OFE��	�|��Ƙ�ڪ_
�蛼���$8~���U�h�6D���郆���,���+���lSM���[a�..�mּA�/>̥����{�����<|�l�9�w�4u0�2"};8^��>�x'[0h9�YM`��Dm�TZ��b�<��9.)��MRPVG��rv��?��H��Xh�~�՛➉��h;��/���fcF�n��.W���`"F	M�i���L>��7$�:��2�]j�ݖX�ǔ7|o!�&��Ō|j�ݩgi�������EZ�ײ`�OG�뮠 �h}͎��d|3(��u��QP|�+3�ApF��Z�CO�;�,O��1�#ʧ��,��lO�c�!n��K�ݭ"�aʈ~h��V-Yk�0�C���C�n9��~�$�*������ۼ��7Ԫ��}`}��<ˋ�z�MY�_�Ikknr�r����*#�M�\�i��_DR�$�2�*�;��^a(�Ulk#U�80�����!JEk����gA%�SZZ�pvHج�s�7hV���l�lČR,�l�5���8�e���č��\��v�%Y��n���7{}��Ò�^
䬾�h������ky���Jw<Cq
.P?GD�
���e���t�ob�cy��$��y�R��й�۽������R�{�xid1��t;a���8�/a�%:aiu�bTKl��|=S���\M���f�<��z�Z+ǹZ�e�o(��xr��M�-!�x�.ʒ����q��?7
�@f���e��#6aY9�L���������о�#Oa���r>Y�b�PJ�Oj ��t䶲�7w��Y�9�]w3[2����_����>E��`��i�*3�	,ob�[�xX��jB���|1�U�v�'uLs#�����;忊+��cA`.���TS�ƀ��mn5������SX�[�7:ruk,<�';�[rԏ3`���j�d�&4#ި46_�3�9ʦX����mI�����sπo)Zy��߾�?5c~�����O��-C����͸ֳ���#'��DT��P��*aY���5��̍�V����A��D�z�=���Y�x����V�f�yoc�9E�|Y��,���F"s�;l3?wa�n�^m�q00�>t0�-|��kZ��̋��,'u+����E�#���
Ú}�I����vh���窼��wȵw���?$0*���$�Y����j��F�?�8��Z'R��dQo�(��m͸�'h�艬m��9o�����\�j]-��-�諭�;���pzy5��;XLl�x�(��L�?<�h�B����l��ex��L�;��݀������.}�6J���~̈́���;֥�����G&6_�R��Y�#�P�i�0N�Xב�� U?����zYM��}甆\k�DV9���≿��c˕"�FH��;� �"^h#sH(|=����b��ӳ���b�9�����!��E�k��"�,�} ]��5�IWzn�]��7j]�q�閉�|4gٞ���9ҙl�ѯ�l�1#7���ߝVE��hhK����Ɲ<�����m`I2��_��aN�EE�'��b���r8f��~�\����˯��ˠS� ~���������w�h�B;^ C�/�|z)ｱ#�f��;�԰ي�A<g����M�(�jހ�0��̼-z�!�����ݖ��&��Y�(�Žˌ��B�k��j������ٯF�6P%m�~����}a��`�����z�i`z
�E�Vg;��=^�SP��e��&��䌜s��z}!cE���gwm��� ���ᾯ?������~�W��<||��o?�����;�x�K>3e��y�F��]:JM{��L�2�5fۖo�jf��M�E�3%f���U!ES��Fw���Za�x�udF�����t����#{��&��D�Ü�5���ǽҗ'@( �m���?;[�����S�u;sSܫ�ξ%S����[�����N:&l��d�[H������]Iz#L_4�<�B=�NH<q$�C�֕15�˷�qJ�ā����;
|��� �y-#���0�����a�P��.=$LoԸ*�v�0�\ޛ!@��Β���K%�ؔ�w
՘�#��".�V*ٽ#\���em��rT���_�������K��<��� o�`��b�b"�c�;�2���t��v�m(Y�7��e���P���ُ;��%��;Ĝ��s6�o+F"��KH��R���Y��#�SP�s�s:��ʽd��fkW�l�2�!�F��Ob�[;�2�f�8��{��Ph�H�-�k`�:W%�q[��
��Ϗ��}�|{Mt�)�ɼN�.�|~�>�;w��L��Ye�zI!o�˄>5�9۫9��kz>Ș��f.�7/l��TZ`q��Auw
���x��.b�˷Wk1+T5��h�{���˔$"�[h;B�/��)�c�2�o�i����54��1BW�O]
ŵ�l�O��8p�f[�
�u��]�&Q� �u�QY�Ӥ�f���.,հ���5ؘxP�E�|½���G^���&9f
��^=��6]b��ٖ��b�J
�k[w���@Z>P0�Y=�#���q��0k�fW6�}�n�r�������a�n�.Bj:���<������򚷆�cBD%���ufN��V�Xݾ����o^�Ċ�$��p�nh����JN����H��Ė֔����9��z7C1�a;��ш�m�l���([s������P��λX�rf ��w� E�E�v)j��j�ks=yf]Dz�R�E�^b��������V��]�H��-٣,�vL���4�C]�t�\��tl��W�+,�+�m���v��F�������-�x.�쩕a�\3.Q�M�ť�pOQT�W��{9!�S���%��/�Ʈ�QF�4iҖ�|f�!��mLZ t����J��f�d��{eg`��gt[�2��4�� ���lŐu�4)A�u�rl1/��R������鯶��YmL�*��2X��9>��`=xmuە0k��W�03Dn�{��
e2�;Hٲ�J�S�Kx��w��c7�
䳆�\�L֗Z)��\�JDM�/o������|�&�2�0�p,4�G��]��+r����D[��k@�k7���nZ�� oWU��NH/J�F�b�YɆ�Su/w���S3�sQ���m��ߖ�U�Vm���W5P�1e"q���1PYF�{���!���w8n*�������V�l�cs��zZ��%��v�@Ay�t��bj�l]!�m ���^
Q���鵏�D��6�����f��4�f��E��@`�A&��UE���QT!��{%uv�t�U���Q2]�m�V�g�ݫZ�.,�]zյkA���.�F#���Xѳ�lѣT�֮,�t;�����ӌ��u�"#�Y�l�cf(�v7ZJ
y�).�6k�u�k��\:(Ӷ(�j�4�4������#A�h�6*�)+C���tW���lV #Z���clb*1��5V�c�A�Tb+ˠ<��Q��Ӎ�-�h��&6(c�wcX��람ETs�Ӯ��[�c�X��:y܅�QF��4i�w������-��:���i���** 6�F���Z��8�`���Tt�gvBD�5T�4�����vZ4��E&�����}�K�|�{]������b~����W�'��^S|���̸���k/n������ܦ�^˙�������}�ɱCt�D4a)�Z�L��];7�Xa*"6aY,�6�f��o9�y�q��U���y���>h��n��$�����Ap��z�]�~%Ra�)�t�kg�t	����Wi��~�M�������R�K�#N3����K���I߸��.g((�-t�ʓU��9�u��{�m�v��-@�<H��H��O�E}E��a�ڬsP0slv �6��e�k2������L��cQ�e��0��#�u0u0�a�N�0~>�FBp�;g�j�}�3{����/��9�Ts�.���j1О��=�|�'^}��D'�\[rz�c��9rY{�-��2L��RFl�y�J��N樃qήK]?s_I�5�T]�Cs���pR�\�8�#Υ踶�p�^)�k�!�:���3P}��S���3��/33�
���!h��V&N;����	D�-�1����3��{΄C׷�~�r%���u��̰�l��@J�:��s�%̗��~��������̚�����awK��c��^<�j�'}��D�R˦��w��z��Un������C���޽6ӍR��$[�j�:Ŷ:@4[ޑA����p~�����_��.`m����-C��X��U����'L�����/�i��]wAѐ�cJ��ۼ�C0�t�̬�s
�˹�M����M�Q��v��=VwN���X:��o���oz���噕r�1�-����fv�ꩊu���|����7����?Ie�H���i�"lb�z��y�<�mt�B��Lg�2=��{�c3Vwf��D4a�z��u��{ޘIՀ�)�?bS�n�̘�~l���
�K��F��Z���;zz�v�KC]:������`I�LS��L��_����/LT��#�*J��/f��K���lb�x�qFpr����5���ky�d���U�-#%�cÖ��>�� ������6�}^ƈ,��&͇^�Z�ɔ��G�gc���w�f>u�A/�яz��?��t�R���+�_"�i��P^{ʄ�~^��l�:KzI�Vcv����騬�/LԗkLvlgfF"&9��̶�{�co�ŗ`�����A���)��{>�Y�l��l߳�o�c��"�/�lx�+�������*�<k��Ϩs�c)�à&��x�ݐz-�>vmՂ{φgF�W���m`�:e fw_5�pu��py�I�`TCv�Q�BKQ�@�򉟶v�o�F�d�w�v�vݮn��x���S�ܤ����s�%���<_��K ��K�3�#�r�⒢rۍ���C�gI>bx]_���A�F�;Y��)c��$���H��_>�kj'Z���Q�g��s�\�Zw
-l��
�I`t��"���\wQ��I2�"��}yzc����{�'���x�}�΢��t*�2���*��d��
ĝ�����{�j�9���xm�y�s	��`T�Yȼ����-m@^�2������|��2Z�r�c��JWETgw���n���T����ʀ[6# sO{���k�f���"!?x|˂���`�~ũ�����������ik�&���1QDQ�K}.�	�]1�o����ȅ:r�����9�<q�@�d�B懲���6̸�yS%%�A�sGL����J�7�����n�i#n��oUh�t:�ׂ�D^�a��iULyΨ����,�3usrmԨӣ�
�fT�x�`�����z`c-|m���Qʑ{s����M݈��62�P56�tlT`ؿ^����5��q�DpQ][��l��i �H��b��� � 9���W��^Qf5U�lɽ��c�����9�?c�.�}`~Z`�uu�}v9S��#|J�N��3��O���m�W�d�@?O�נ�1���w�6�� ��W���#��ݿ�� VN�r�jگ0��OU[��C:A��Q��c|�g��Gh0N�	���z>���Л�r/�11�X`�=�΍ɨ�B���j��u�w͸�7���m��K,O��OFmt���Nm�}W[gv�$F�뜢�V����M��nl��\�\�nMű'��.L�{0ɀ��i��G�bv�ƹXz�[Z��p����9��S�2^�#y&����謹�xxxmf"�*���u�m��Q�k���b�-B�z�Ɉ��-��h��O���ި&�(L�e��G)un
}�&���\�g�Ud����{�(<~��}�;=5��*x/A|�]�1��[��R�eD��`Z���]R[�U��*0�-�r ����c�Ηs�(l��-�]kb}Ҟ,޲�	�ɒ;��@��zX�_S��Q��t�����m_w��������+p�fއ�ny`i��9��T���ߐU�t���KI(�7ɗ���Ҟe������H��۔СW��es���D�m8��X|���v��Q:ј�5�4�Q��I����߲~c���T�}�˛t"��w�fz<�e7�H���S���."9�����1��T��k��1�]��3����j@L����������3��a[�m�=��n~5��I�_Y��f٬�'M�B�df�Ӷ�/cbddx�f�0E�;\�q�wE'\��)9�R)��Js�k{��İcF�V3/��Ɔ�v��	��b[�7~���s�B�\[�U���Zr\ ���*[0Eľ�ۓ,�����l�t��a��M��Z�J�j2e��U�.���s�'�ʯ�1�}0O>=��{35��EJ�"���1��\�zQ�']G{sQsiU�m�\w.�'z':����tX3�ޛ+��KJ�lu��)�w/{��q����;T��x =�xxxH�M���B���c3K�f� c�2�kPK&1��{)�A�1��M>�>м�f�gRWۜ��<^��������9���O�E��yͥ�:Ĭ�'�_Ph�1�e�QG�8TYߨ������YT3�%&ϭE=�N �g=To]?����/ϭ�
;`ߦ;�ma�^u�K�s���"T�zS��,��5T�O6w�[^(8�Q�Jg/~H�e�<�})�+cݶb43F����z�ٹT�����yO��
z���8��%Ra���������ིp���qKG��L���Ӊ�`��e�P��+��������K�v�?T!I�GH�� �h�>A\N�ݝ��f�O� \�Gu�0Y��{�VO��5�;���C�ʹ3��Q�G��)�Y��[���z�!^�הΒ~�z���[�|����!9K�}��fdSG�.��˾���� �_���zo	Qޠ.}�0�2����1�	�� ��9>�G��Ku�
���+��isF�6�ʚ��!������l�9L�B�`aQ���*�A�urZί�s����x��$X;�s㗯�}8�2T���T�,E<;!�|��Qm�r���z�㭔����&z�������v�$Pj8��{��y�c����S�a¡��BV�v�*���tPN�x��ce,Ū8go
���_x�D���Q���c�j����UE}{=�Mˁ�9�P��$���\�	�;�{Q�-�ef��{Rf�����Ј�p2�Q������	�+^�t ��ܦv��k���wܙX�x��'�ߞϰ�?܍������+?S�/�Q*�s�k*tr�|��`hȮ���fc��SWF��ƭ�e͛�XL�8��ճ/	�͏�}b�*-����Z֏���̛L�i�W�ʙ�#��*|��V/^��e�[[1�}w�2.D�����[�ͼ+`6��C�����m.��C-Hf��K�s2��<S.~J=����clOLx��I�2�Ў�N�Z��/7�3��!��\Q���9��A��I�R��e"'\@~�n*8�Q�$��R�y���5�c�Z{)�g��4�&4���y���*�2�r�s	,�9�a�Uk5D�׹m�ǥg0������# �:=�S#�UK��Z������J9�����RΡ�w~��KY~]�ٜ�=ý��\r�a'Z�����Lo�� _=�BG�/]:?N�^?��iq��؋q,W�Ux=�h���r��=<� msyk{]�u�N�d}z2t��]�=u����j��^q2ue_F�[:�����v��IMO�b��c<���4�1�]Nb����+��z��%��{!�P����ٵ�}��_#.�g.�w�{���
��|I�����1��F��Z/�e����>.����ҏz�Ɩ �л���m��\b�s�i��3s �gPc���Msd�	��>P6}_��'|�G��z���f��ծ��Zw��h��4���׾Z�zc�X���*7ި�T�zU	-t�:�=�=4�a��z�fk�/j�"ƌ�߅mFxu>��^�v>|�� =M��H"|T��ѓϮ�D�[q&���H�����~ã�[Y)߱������g��Sr�j��@fި�c��ۣ����X�Pw���9�'W���
'~���� �R��n�h������l�v�?؝ǟ��п��G�\�B�z�T%�ɯ��pQ6,TuaI�@�s�=W���W���7
����e�S���a���4ˬb�oiWt}�Tɱ��;�9���,a��!T<�]Z���\{�$ƒ��	��EG�q�	���e2�	U2.sT�uYX��0��1�e�L����o����}~���Dmz`&�z�5����s�1)�	T��n��M����O���È�(��+k�XօU˱�q;mX9��֭��y�@�1�Z���f���g=��qtb]wI6ov3��M��T����3��S��wø��Ѵ���u59 ���C�����F����*M=��Π�cv7\����G4�*��i�@� ��F��N�e+m�����@nDc�:h	��=X���x���zԸ�iIOn���\���=�����x۹�-�'_���r�B:E�g�	��OCk�<1��W��%�D	��\�DA�Z3�.}C�Tj�&`s�/랬e��#�}�����I1�g����W���T6�
�3ƽ90�u��1����?T��ބ��1��c ���ۆ6�����Pa��Ue��`o�lYz:����:�|b��i7�x�:�}��������������>�=����`�c*nEwk�~�SXUf�.W����9!�{2�Jx���i�O�Դ9m,j��0xn9�ј��Ӂ5<�6y5��@���W�<�ʆ#�ӷ�@3�9���}'�`Õ# D�6�+}���-|5��/�VHS�0}��eŕ��w؆�w�n�d՘��P�}c�;6�iN!�q,Hޛ.��Cy�h� �/���n�T��'��X���ӈӈ���Ύ%�3��Q�h*�s�#C~�PTyQg��t�������3���p�,t@�ByY�SFh�oM2�[�I"��kjd���G���a�$cz�yan^��f�[�{�i�H������ lcy�t��=��!Ø�Ջ,R��խ��*n���}%��u����s�x<���ML�����.cpS�e�H�>�?����֜�Y�4vϸ[1�A�2���Y�D{����ԯ�yj�n��Rq�QX��f��&�TI�&y�b\H�۫�F��̷	�P����>����%/t`b�&��ɳ~o畁lk��#/I�A
�E�>W�dCLſ��EӘb�Lx����wE'\��S��h[u�}ѯ'/9/��8�?8�qF���m�|*T����������xE}���Ş��#s��ZhV�E@t��`�n,�����[j�r^��#Ք�L���d��瀛�D������;m���R9��ݮV�t@ԡ?E����#ԖP�r�?r�x���O�T"�<~��c���^�89���W��(<�h���`]�L�	�ڠ��7^�Gh����|�Z��j<X[9Q語"h��=����.(��R'�o��n�_�˔�^����p9�@�����M���E������h�h��|�b ��!�>��֖���o��s��óc�׭l��SՄ��67����K(� ��8���4d�K���zO�:���q8Ҍ�ozq��~N�\��G�;����.���q�uB8�Ω7GW���9WIP�:l*�%���K7裎�!��-c�X�t/Ob��CuS�+���Xv��N�.w{�����/��/����j��뾄�6���SQ)��]j)k�ǥ�U�u��u�zw�=����-g�.:� ��&��^�_ʼ�<_�����Y��!�9��a��XjQ�uy��=�۽\��j�t+w�G�[<۞��.Ȉ���Κ�XLM|�+���6 _}�{�%#"�������+��`�����ƀ��zs����aze	eG'|��i`G5s
M2�����t�i�k��������<�-�dL4�ܔY�d͏���<��9��k��}=�\��Z�!Z�U�t�]<�~F�{�A�n��׼��u&��I�n}U�5c��'7����\�u�?)��'��g���!�ǔ��09�%3~������W(D�m<<'��7��cF3�7޾/���k�� ���s�B
3r�O���"�ʀ}g��D����T��,`�y^V#>^���w�{��g0��}Ί/�mȭ�X\]�[t!}�
������VG��>���ކ����˿�(5��� �莞js2��	O�61X�{Wr7G�ml�c븦�����G�*r���J`�އ�p5��E�uj��c(��!V^)��J=�)��$�n�\?3�～oG�����z�~�W��<|�|�?���޷���X�>i�~���	��Q@:���5���Dۖ�oH͡/0Y᛹��_M�v�A���GsWr�%�Tބv����ƛżsL��%��(*λp�t�*�e��k�V��גqV6\�+�Y��Y�es��mT�J��W#���G`<��P��jSzo�0��.��e�K�0)�0<j��t{y&���k	�Y�QY����T�4���nk݃n�p��-"S{�n`��F�6��*����8�ݲ���^WBݤ�P{e9�MS=S�E�=���e�Ԓ�VŶ4d6u��b'+���B�H�^�i�}�˿Ļ�G������/��6�s�mD�]�.��WC'�FG>Y��ī`��."*��JJ@ͣ�8�V ��,���{8S#��ۚn��q�2}� N�e���#yV>�o)��*�vMth�#z�f^��ZY��@ɂ���R;��g�U�_�/����^�;�z�U�'�t�����l{����hjtu�v�v�"uo۩9�
$�ݻx\I"/3]�7u}�bo�W0�|4
g2���N6H�XJ�t��r
7ē��z��6g_7-ey}w�� Ե{\B�����ܕ
+�Ւ*�R�wuLk\�<��c��$�o�K���;6�]F�ۼg~�[��4�CM��KJ�o��n�@����x�%�����c�pr&"m���\Ǵ4CJQ|Y���0]��87�׌�u��o������Z�:];�����˩I?c됱s�J�ݗk:�t��p�P<P�d�=ȁf���4�/N�<�B��u�Y��_z߇~g3G���ri�
�;��:�v��#`-�ubNi���}��FAv�v�d ���u��h�{{�j�>���I�s��1��[���w�ǩMZ�M�Y�1RC�]5l��٨�p��()}o;+m^GY�Ag:���wQT�#E�"���8�0�{Wҋ��^�㤱k���G��@�g�]�.����3�.�d\�w+xK�U.K��-U��<�]��i��\��l�	�*�g\�TCh��!	T�`������]�	}O(:�A�|(��n�U؁���S#�R鎮�0P�,Y�t�TbF��gwT7jqZXi=�eRhw't�7^��r�T�*��e���� �)i7�9��9{B���4���o��j|�4���2i�;���D�n4+FrE�d��g��L']�q�by�	'�MU�f�Dt�C#n�i�d��%��<ٽ�N-�)nq�W���G#�B�j��}v�E�Ӻyѵ����m�bT��qt���i�:������]�	��z���v�y=��D1_��5���={C7.�6`�������c��8��[.n��5����k#�r�-��v`c#���X�X���y,�1��K�k�r��k��s��M=;jh���m�z�/��N�gq/^���H���e��K-�Gv�-������"5��;e��wݍD�%Q�M;v訧u�v�kZ6�n�������w<�֭Z*;q�Q@��w���cD��qL�X�GD@h�-m�lQ:[����6-�+��#���b����Pn��;���6�v���P�%Ql:5ѣk8��f�I3���wQ�E�w��1=��Vƪ�؝h�m��E�������/xa�O��*hֺ1����%�-Z�;`�v�+OGW[cQ�nܚ�n���#�K]4���U��������A��5��i1ѧ��D�]&�lmv��v8��-��=c"�ե�lc�$�:v3�A]�QME��6��Sv��<�u��)��+Av�SZd�v��bJ��n�����s�U�KY9��Q�>��}u�h��o�=܊�U�>w�.��~�0����2R��yZ�V����EE˶��j����&��"bO}��m����K�ay#���0��e0�kj��q��Z�ն���uU9;	��	%���gQFX��Lxw��\o����F�_��<���ɖ�*nP���W�兛'm��u�+ƾ֐Lb�"5�C��4C��*=��hVxqT����A,��ӏ�d6iv���s9D�k�1oμ"���Gx߇��*�59�QL����		FD]ء���	��`������n�F:����mjc׋�n3���ƈL��7���,n�}W0:L+k͉b�	&����������~�/	�4<�F}_��w�	#N�n�z��b��ʏ�\VWqTC:"᭻ �U�^~�u����z��i	]&^�BK��z4�jN�1;�tO��Jp O����b��+��cs2���%ۜ��ټD��͇7�n+�Y�k�׹�ok�X���ã����:i��3_-ݪn͹���
=��~\�Ʉ��WU�-�@�S�}�Y%|%}��dsH�f��ʏ<����#�����!�A��Ώ��g����{�:������Մ��3�r��e��I�s�_Ua�\-��4u�O��&Yi��:J:wE�
Ie�ѷ�AΧA�:�r���ݻ�ߌ��>������ps�^�Cn���ʞ{�\�f�����5�܃�f�������f��y2�E���Ah���&�0"�5cH�W1����ѳaw���QW�M,eɫ�M�^��s��H8˶��=m��2}��V*���y�q�Tɯ��/�'0����>bM%�����b<��%�8�*6�f�>��L=���ٮ�r�x�B�ʘed`0��H>��K�a
w�Y��ؘ�;�1T�qY���9=�ܛ�4���Lw7Hi\^��E@;�1E��N{i�mM��ᘰ�L�>rF���c�FL1}�0l{x�/�f)QOs�vԔȚ��i�/Y�+uT����Jc`(Z�Мt3��4��$C-/��ێA}�[?�~�g�L-��M|�;��Bv�{
 �G��^]8/ �1��zc�$��$^��51��X���*O���}\g�Ԅ�caE���FPYkT;n�z^��?t��#���syS*O\��o/LO:j��n��R����϶:|7��
��K@�8{�c�71������MSf)���-��=p(?��#�<��*�k�4�>���3��s}/d���F���!��?:*����¼���L�L�c=����//m3c�����3��UWu�l�KN��s���❷w�1����#k[5�	5k�͓���"az1�������h�|K](�}*Y4��nҎ�>罹h��;�û�h�ԉ�:尲Y���U�d�i���������/�?.�L�g�i$a��?a-a��^������}��(��;c�ܬ\kss�'}3b����f8�W�9��p���sּhy���#�������f	�O�ٿ-�k��������V�<�кn��:]�~�PM��0IS|��f�Y�$� ��o���s�Wԧ����R�!�L�Ԩ�\N��8�ұy��)�69�����T��Q:ј�4ra���KF4�ln��ys�5��ɬhy�k��gs��CyK��"��ՉGc�<��hW��q7+�t��5(Eɇ�]*�Q��O�}��a3!�ϟ�!�ޭw�Y�'��f.2%�WRƤ�,p�Ļ�Xہ�}
����d�d�飇>�)����9�[k�z[�"n��3n��ᏽY��u�X=]_�D؟9#l��u�K��������#x!���ǀÔ[����4/P����nL����1�����m��uz�g��WZ)mNjem����~�"�3���(�n%@�ե�:�+}�%�Ѧ�d�E�>`={�=�C���gi�0n�F������ޏ��+�t�K�1(�Y����e4h���}�S�TcTk5r;�Y��L��oh]�Hb�>��'l�������7��S.�V��e%�����+��S��*����Y�_��~<�{�}}���_o���s�&��yv�7�jܢ�<�=���N�M�n=qSI���9d^YzE���{�>�����ew	H/lj�;�u�d˜�M%���8���zV�۾��vqX�}�H��Nϭ$k��_�e�����E�_GN��J�f�}<Ѝ������-lj] z�-�喝}�'�<��VK8��
�.4"�Z��z�s��q���tj/���hf}��&��ݮ����z����D�1i�6�?v����ɨ	s�k#ؕ�%�ݵ�F�.~hз_N���n�&&{��8���W���B>U��R`���"޻��[N�xǴj�����s3́ -h�3i�7nǳ��q�o�]���5��7tL�,��4N�����d�{_U��mҺ1��\�/OIa"&-����$(ܞ�0���*#�N樃s��&-C��s�F[ʻ֣ט|�aC�;�V'%�z��.�t�Eỗ���'�<��P�	J���0��I���Z�IqST ��TFd�/�C��M�3��Y)��rhF7/}�.��Ӹ��	�����l�4\��7��.���ޢ�w1E��]*�t����t?Co��{~&n`R���_�ç2��%����ѽ"��ww���&�2U*�y�����sWr�M���씈y
%��I(��melVe<�uuXt��������a�O��b�8���EW��� ��=�=�{����+*���Pf
�F\��+l_(���W1=P�����m�&z�K�>f���Z�5Y�c��e�4C���bZYgF��a�O׋(^߁U����ڈ���H|�a|"�}��_Q�2�n���׆\�lM���ۭOW����\�����x�^=k2�߇-�׬:LP�s�����Jкh+�WW���/��u�@���1کC߇L$���)�?bS�G,l��!��d�o����B�����<G�whO������I�jS��U)�����eߪy����K�U��{�NN�&��,~Dg�`��<��]Լ|�yk����O)d*��۹������}�YZk���Ha,���ޮ-�|�����l[��QRy[V���y�ݴ�5{$Ê\MBzY�2�RYy�>����#Whlh`� ��|��	�����tx��H]�q�y���7������W�G5���Mw��Cȃމ����,1�����{9���ak�y�!�#�{U�Q1z�Ʒ&y��dԖ�&�Ψ ���n�7�}u)^���\i��{���(�#M:�Ǵ�MQ#�#��"�h�o.�Eu_iɤ�o6��7g��e�j�AkI���.c��fn�����k݁d��	y��������)[W�j.��!�ʷ�QSK|ѩ��}����������7��f  'gT������l�,�xi�=C���\�CH�������%R����Dg5N��k��&�(ĳ�U�lΑ'�<�����ڎ��/)�Wy.T<߁�Ѵx䱷gc��Dss�8�:T��t_�ꉯ�]�?�5~����g|���&��{�3N�f���I���6%�p��Cb�$M�]Y}��H�l,de�>f���r�pG���뮣s.q_A{v}6�S�9�4^w���n��57jx&+~Ǌd���2�E�	���,q>�ѫ����'f;����y�U�	�3
ldw:���c�f�y�\]��Tɱ��9�7�=�[��vJy^ۮ�vY:4��_����hGD��	�pJ��s�k~�蛌G���~�YQ�wh\M9�6�VQ�lcq/S�oL��ȇ�ן[��,�A��*�{s��K�R[�u:x�N_�.c��7Wv�-k�����1�5�,�[���GN~�Ǩc���ƿK��z��6�i@��[�>W�๻:=ǆ��=<%��zaj�g�A%��F����L�ؓ{�"5ra�D�tmuzv�u���FF8˲���C���J�}����{7**ro�8�����\����cv�b˞�N3-.U���+C�nKNp)����vXEJY}��}�0��M7��ozY�����Mwޖ�h�`���s}wןE��{��}}�>�R�B ����'��%�������ߓE�Dg!��o~j�"���Oj �G��Mm������8B��=Q>"[�}^���|��D�Q�����q��q�gW��6�/�Ll�^sÞ�D����7��j�z����?S�u��������/��嵤�궰;��~��Z2���I����Dz<���ua���R�2�Q1a��A��̪#�x����-��߸Ϻ���H���4�ܡ�-�2=�ݛ����y|Dz��TO�TI�0*�)�����y�����o7P��X9�:�M�c�H�k�%�{�d(�U�כ�Y�9�'�Ś�d�dg�`nkGo�Q�B�'����5g7WU�W}����l��H�TRp��7P��<��Hw���_S�2\e��z����!�5Իy?h���}�޲&�ζ�t`��j5R�}Q:��b�ܻU��,�>��|��_L� [�����+��G����zC3�<:�Rq�Q������/+��n��Sӡfߺ��'|H�.z���B�c����Gk2��gK�·4ۆ�!�>�yC�ޙ��d-{j�ww��D�
�%�f���9��q�m^���T,�2�SGN���u`u&H8lSk�Pu��������WM��$&���d�6�jc�(���><������j��vIo;��Sgk
�Z��ϯ������$Q���}r{�]q������xk`ǣ�C+��g�"Әbo��3�+�S,}�&=��/��S�6��S�;�˛0%���(?=���6J,���7�D�QM���fg*�zYgM���Fv��ۭ«r�?OR�Ģӓ�U��kQ99/^;ˠ��D���hv���jS:�E��I���tk�#�7�����s+�wT=��;�eC	=��������O�;w�ON�ˍw�����$`�L�h�[� ��α�Ϲz��f�+�s��u�{�s+��`�&����[�m�s�G?��}J����y7r�K�&K-c����HP������y�V�Q$y��	��xE}.{�Q�/��\j:���ae	���Y���;:gJ�3�4wP�}�����{��V>5��.�`�{��<5	q�b�='�Ƈbzr�7�T���7���'��d���Rj��X/ʇ����8���3�ϧ�@���:	26�a���ɬui�.����V=�-��ܻ�2Xe3e�{Lب/cK���K�B?�[���n���f+��WW�~�� �k��a�����A`(lo:�S(�����e��WGЭq>�ַ{���zbleio������ή�<\���LO^�,�����kksQt2���awWa��峄�jJ�t�T�Vޝ}�̤�m���>�{�>��?�����BA�d��v&j)+W/��ܲ��s��=�t����T{���n��BY�$�����4=��nO��}}~���pN��ϼ��;1Dln��B��~$\��6V[�޶1ט�;=�2���x�/j�{��5?X����R,�,��᪗�{��Jm!u�.��*�����������3'!�m�xjP��=pڤUDY�b���s���T���C��l�z��7Qp�TQ�C\yⅼ�P߱�L���$>Bpe>'������?�$X����o~���Gǌر�x{K��z��n3�nJ�$KƏޢ���Yxth�b���#�� ��9�;��ǜ<s�U�h�S������ߗͼ�P��w�6���+��B*��6�z��g5[�p��GL��c$ �|d3H�R��fQu�O�l���l�T2#�BF��̷�=�3)��p��.>e|fpTIa�Q\�3]��Ph2�H&�7'�+�:l�]��C;S�.���u��B}�{�څ ��"b�XW�g(�,r��;�a�5|�B]�^��M���`G��M_eq_4X��n�^W�N��cm��x��\wJ��J+�o*��ލ�[�Kz��`X�e�"{�[�/���쵍T�qb)��3��*q^Ne��S�'sv��1��fmqu&-���SE���r�U<\�@�9�7�^$^�~|���� y���x3 <�<<����+���ܾT÷���y��kVV�:����X?=<���$��ح�q����MA�����:�#�yY��ޝOAdw8�),$-k>��\@�Q�:> gx�܌,�����������F&`���y��N�1�C��X�5I��#�,��kq{h.Av�C�mwWE�<�u$��wA�ds	�鯮%��U�C��qC��o^&������P�T�3ڋ�Ga�pݲ���؃5E�G�é��L�-#,+=�զ�1�?[���Lf;ל�k���yӐ�v[}������]B�y2�|��F���+N��þ}��4�O����u��,���T^n�N�6����3m	�t����c��|JME��Át�Ñ���/�I�Y�����rW9�\⢭>Y&}�Ԉ��#<����3`��+hsx9T�qR��쭊��@�7O�]�7 ����ʂWB��^���)��pM�����X����{�#[��Ju
�h7Szc�s)|��S�ܡ��]4ǐ��7�AVl]�U�2�d8>��/���}�w��}�C�����~�,�t'cU*�gg�C�	K��H�v]�.�����.��f��l�[�Bю�������GK��@a�>�N�"/�%�Yc2
��,�*�6���S{G.���QX�[E5v��K͡�l�\$���#�WM�-��y�2F���s��
Ŗ�
��@��2�	ŝ�̼J��2؁���b�bՋmΣA�V]s�i�ĉ�H�ݵ�to0RZ��ìl�e��(f]]��}�3�^�aܑɼ���&�3x��Y�t����,xvW��Vm9�ˮ�1[k�۹
5�ՠӄ�F�1r��lΚ/�U2w�D��Nd}.Fn�RrYo�(����N��`����¬��m��>�y�Z��(�K���(�d��X43�'<=r����V���֧98����l��X�
bA��]��]S뤹���/vՈ�jL�l��,�'Gy��́BM�6e���bׅ�	��0�1;�^_<!1�!Wt0(�ǣIC �r�����^�9ucu��t�';5��ÿ&9�V[�ES�&Mf�v�o�y�á�۹�������'�e[=:w j�;���U���n�]��!�N|��:�|\p�7$�"�lVV�Y�)�^Q٨��-�J�bJ^3�������Bt�ktsC�\ΡVضo&]��{��Z=���((�̨�U��Vq�p-��׫(\���Vt���=2�j�؉�]2��i�Z����]��b�)ɷ�T�+V�76oы��5L� ���j;��y���iw��?i6r�7���A�����H�����(TH闧ro���ΎA�4�:E��)��1'w��܇5E�i[�c90F
<��J,��p�ta�X	�{��i�5)��	�n�����i���ل��v;���}����.l7+kn����W��|��+�d��tS/����ID�1XyF�m_6�֒��`�e��l�Φ�Nڮl��w9�4L5��&^��[�;�NnܲeۭI��M`�e����Y��B$��:v�^R�*���@j��؋����ϲ5;M^�c��c,�l���m���\���J���)��պz.RIG�����MZ��,����Ņs��m'�6�uW���O���5hebyҶ�,kub��&.ޱ�mjYEk[����Ze�VAfΈ��`qХ��ʻ����D�~��d�;rWmt�q�cLַ�۬�}��Z��෸���9A��J�3�
j����{���2�-bH]2���t=��j4�u��
�2�c�QKY@�sk��=�G�e�{*��y����V��Օ�\IO����Ӧ�1o`��2�v�i�wjx�eu
)�e냛��y��bB	h�܋�;a��W"��./�tmu�*������(	�òG�:䋧a�i�l��̄ͬ�I�g�M�V���v)3SqT��c�π�;"4�Yy(�.��=:�E���V���Ϡ�����M���	��v4�vkk��X�n��Si�v{�F���h.؊�F�j�]t[i#�m�[���Jx�'v;�b�ƃlt:4S�D��L�X��Ecd�:�.9�uPF��؊j�n�v�A����T�:��颺*��b��H��;6�4i("�h�OOq�j+����X�f�M#j&��1Q���8�؉g�twmk�t�-�Z��@EA�EUv3;f�U%��I��4�==]h�����κ5RL�l���E�m�a�������ٝ�1S����);`��*64E[m�`��QX�SRiѬu�u&���`�(��EU�[j����*h�ڴ:�=�n�]خ�m�J�lZ1QV�\EltX�J���GL�v���51EETQL��m�=����V�!o�0�׼9���<:�Wb�Ӹy�Ϲ���*�x�V�C^�4[�|��˶\a�ۮıe����<U�*�\{y��n�A?���ycu���#o:+��3U���?h(
��h%V�H?�n�4{�k�w.�x�E�H$�Ֆ��W���G���C����Ex��0��P|{���'�z&���S��L�v=�o=�̩�y'�(��2L0��c��.�����ft�ä�M/�����ۍ��J[95m��2u��Ѩ�������%�Y0��xTq�ur-��p�k����½ز߰�5�ٸ.W�xrn���= �H�Z���3%��	t�=.,q~��Ж��y�؜,������ٜf�X�S��Dw>�dv�yt`�^=��/d8���c'�v�����EmwK������dg����R�jYaEx��层���]��m���E��;�9I̡��}2|�/R�Κ�[�=�ƭ��<_�.�є-W���Uiܕ��Ϛ<G��_گv���v��C,��fC���Ϛy�)���t�[9����'����1�&��Dj�^��ht���\��mPXH��	
0�xc�9�ڨr�Z�!�IU^ܹ�������P-���bw���
f�ш���|6!�:��͐�O����(����	�YOև�^��
W_xt���ǉ�)X�cpY����+s-����3I�9��۽gcݦ�3��fdy6�M�=n�\��.�XŨ�֜}61΋은��[�M�ĳ��uø�&\�SOr;��-uꛙ�$ٍ��\�<�Q�j�kK���u���D�$�433���_7I�[�I�{�*�4�������"Ă���=����.���de@7�BT<�}�1��&�ak���h��e|��f%#u����4�uǧ`��Y�5�K<(�b�W��PJ����Xo��^~�M1�y�_�l\M�F��O��O�,���%����`wj���8���=oF�w�We��T�r��|y�Z��B�T�x���`�9}.�_�D��ݮ��F����I:��ϹnU�o��͐}�Wh����$n��&�[ �tIǥ{�s���^4��!���g��E��{LRsx�Sj*s�V�Cȼh�t_�;Β�@O}�͜
b_���*�Wؚ��N�'��>0X�_L�0l.|	E�'��-V0�&����eי�9M�sr:v��P�X�5�`1�2_aH����Y���vv�⨵�QaDQ|���|ղmȶ�v�9y�P77ӫw5��v;�/[�1rqt\�_�󢝫9N15�,�܌?>�hH�Ǆ�����n�R�����I/��`q!�O�XP�yᠾi�P��|�SWa�/C�.SIt�t����r�np�e�����V,E`9̮ւ2�,f��ϡ�g[�Jo:���mڽ{����+}�އ#3�[e*��ޥ��Hs:�/*S���.��^��'$�X�3��R�ޭ�'��*�m��i]��܃�>�r�r�_��!$H+-���"���K��Rfq�u�z�j߿���bDh=|���/�����������߿��.����'u��>"?>�/��V���q�T	�i��_�?^E��8�ĜE��ӳ��5�^;������ �<2@>g�DQ��J�
e����U��b�pf��\k��8Ʒ�Q�^uD����ʁ~^D-"q����O-��{^���hR�S�<������.i�A3�2�͗�b��z��gp�����Q%w�˛�VLq@��\T���c�����a;��'�>��^�BY8��s|*�5��m���4�
�a�'������'
��3�D�7��<����S���OAu�MF��Dc��n�9�	��l�>Q�6��r��]�=�?��B��7*$�u_!*�¼f*)�c5�ͫC˩ι��6���� w� �N��>����P�jg��&�ba�r]b�|�y�υ��Yq���L�wQY��E�<��1�����w����ýFѰG(=y[���+T��tc�$Gd�ll�L��<�Ѹr���鋸|��B�ٰ�m`�!�!ކi�1N���ZI�|%�o{?{
�d�ܡ�^�x̥2�g}kN�ALwb�UA�Jr��i,��ڳ�`�r����SGfl��B�^�� h�y��8�(\�;��w��P-��;s����^�,������݇�0.d��������HR�B� L���z��ӛ�����u��m�q�d�&�Xs2��%>D�V�˨���RZ����ظ/��L0੎nN�=<�ɏ�|d3Or�^��eX���s��>��9��l��=]`�/��39؊(K�n��� p�I��ܥ����������1�s=J�n�xiZJsoK��B��x�0�=0��	&����L�7P��Jn�0Yp+���"�1�K��)cԄ�����nk��/j��-��5��A�p�{&���H9�?2'G@xg��c�����$��t��S�:x��^�b�Jm��P���;�҂�Bֺ:Wz��ă� 0��3�Ҩ;^��B��ڥ]wݫץ�O2��(z�:�1���C9���=I����i|h�`��l�t���t):�@�7f�"X����[���^�g��b����N*ԞU�wU�4�\_O�^rS~γP�'� wN�^�M��Q��?^��>�b�=���:b�����\��ʥ���7�q�����2�}�������z'�<�J���:��ي"� G��N����O���,^�o���Y�����P��3�憗�@i[xH���8����}]GDZ]�v^���Ԝ�}���Hq����iY�$��^������Fke���K��=W���VN�%�[,�R�%�}���3ewU���� ��^p��o��{>�1NK�1��AQ��]��܆ρBF	*m���)���WL>��3�q���{�(Jw�q�3w���%����L!�h��T����<��\��}Ս;����#�\9
����['o��@�%Ɲey9M'��.�ŵTD��v��ֿg)��ؒ���rEP���,�����|���r�~�h$fM�=�"n
q���6���X�΃=c�.�����
̱^��(�gT���[[+'ͯ�b\bWj$(�����<���E�}~j{v��~�7�����E|��z;��c�b����ȼ�Ԣp�7.�B`&\��4�=!�U�s��K����76^tr���/�{�Cn�]��z�eB��3`���2�%�Q�6��<tX�W�߇v�j�W3�e�qܫ�Ř�E>QE��ˣ�������Q �ט���퍿����o�n��Lk��;��ו�e ;��F���%�f�������)���ǉ26c!1q�]��k�X���J�E�F1��0�z�L�φ����)T2a��AQ��c=O��˶��RN3a��.�Y��g>^�������ƅ������5�qKQ@�e��ؠ�G2�)$x��X�.7�b���;S\�/pНqS}�u*�*Yc:
�׺�v0��!R��'U�T��\QD�ۮbowK�n�M4˾_kX�߼ 37��3�'V��yV�|��Y�.��"��5:6w��mxv����'���P�1������R˹�]����bʄ@��1Ǽr(�9゙ϧ����g%���e�G;��X�����·�杺S^�
�htՄC;��Br�=�`@O���Ҭ0�jT	��#,��u�X��Z��ƿ.w�P�uμ���,�5�s�',9�T�<Eg)�(Sk���2���]�)�vn	jv]��Ϥ�ފ���έ�)թe}�(��~�@��W���}��N�%��<%�\g���2̏�̪��n�h�T������J����h@�����-'>�x���^
Kϟ SO��'�5�\M��Z�|���ey׀қ�C'5�Ƣ]۝�m��*�?OMu�#�3]��v��@Z�x)�f8���^njGru8�3�M��`��:(��մKK3r���[Z�c~��3��w�Vn\_��������H����>L1~���\�x��6u����3��P��7eg�u�h��5�i+0{��|No�L���.}]��w#:���ɵ7m��Cw3�6.�W>w2��Zi>4�
��5w�1�,L|��m�=�պͺwS���r���T��|\�DK��"�L=cF�)T(�j'�'Ҳ�����E���ܥ���`�sK׵��L�KU42���{���30�ګm��S�~��a>$��2�����֦�kh'&1��eS<c�7jC�2Xq�Z�#\N�/eP9��/|�"��^0̄TfDQ|Ԥr--�ֲE���q	�����=��Lᎉ��@�O�F�<�vr�m&�A?�tFy�X�63n<��*�b�uZ�ێ1�SI�`�X��� ��<�с��F��!F�=��M:����ź���'�o�f�y�g�`�7ǉ#I�������5ŗ��~�4�xmk�Ȃ�,dF-7;��[�hOAfϢ���sQ�|g�����:�h��@��|hD;<�w��#���sn�Gd󜷨�hrac�+�Sp9�2jz����v�"�8�+y#)�1��ߠN)~I4'������O�՜�8/7�;<�6����(��b��z�<��Yn�.��_
�5�K����O�3��i}�����8>y��PX^ �2���+��}�������U�;M<z��.4�=�f+H�17�z�A�c�̃�fdԋݞ�1�X~��c����)�\���c�$\���k/s+���:#1�����F�ݤ��Te�����5q�d�JC�[w��������_:kowu�bfn�D7:(i�շv�@K�4�95D2�Π�,��f!|랜6���bȱ�5�uTp�9��;�-���og�L f� 3y�z�k�u2㎷B�o��t���3p�<ڢD<��y�Q�^���]��HC���0��LM��Qӽ�5C��2�2%�t\;򊇆���k��`T�w�@�~���ʨ��g�[x��$O��S0��q�'�nS:��VlsZ!�Mr�A��<��ۛ���g�_�HJ^�zq�ڒ;8�t�����3��֢�c߶A]��=\���69Vb��MbN����|G���Q}�	kı[�i��-nfQ}J<��+f�z��CM�g�e�{l���_H��qi�?�pL�rud�/��i��J�fua<S.<�sow��"����Һ�n?���.5�[Ӧ��7�~x�ʄ^`��?b�+�/!���wV͘t��?V��E�����1��:<��>t������(�&��\^r����p�ٺ�VJ�~��t3Ll?�7j���%���y���r�\|y�%���4�q���%q����g�7�m��=���o8���]��|y�߫�)�:{I�{&
�9�,�H�,oe/�mn$5��R�a��^K Ք~��Y�R�F�<���c3���P¥�5�]3OGR��9:r�졯�UeDE6���N�[�3ϻq\�`�oe:WK���ʹK[����͜�f�e�[��oX�����5��}QWJWu�����?~$��O���\:�h)s�_�ff\������3;*)������ĝV7 JLd@Y�zU651�����̵�gއ��>��5
��a|~~"0��U�>>�<��j0v����5����~{�!s�N���濭7w]#ߺ������0J��j�?�bA�<�G�AaY�}�i�˦=��Uc�.�۝~;��@��w��kΡk����~�=0ʯ��5���4�(\%l����C�b����瀼=���v>�TdW�X>��65Ru�DKE��� +���e��b1��|������ջ�	�:�*Ke���jV4��]2'F�z�p����>�������2�����҃������Q
�X���Hh���S�T1�w[�Xv"�����_`�7X6%���mz�g��d�pN��c�S1�ѓQ#�����C;��H>�k�G��kh�>/rj2w7V��/}�Tɫ8O��'0�ġb�O2m�!���5��»�S-�@�'�{M֢��:�8��-\�tSl���a@�̘/*"N	�]��|pzE��A�%���$��t�no��;��:Cs ��:���+�`~g�+$�uò���>M�X��I:�����靚�T�W�;&��8��y�nW�tƖ�tS�K;�"����#��Yf
ӌ�������q�=U�d<;.���B�igV���I�ol�Y*�������	DP4����>�7����b�uѷ��']0��]'@SM�)I���f���f�n�~�#��N��+by��ID�~�7|�C*�QT�C��\�<�����ֺ9��*V�5�*������x�7\�+Ld%G��puƛW�̪�t�~��-���Nޑ�LP�T�rA.�(��}���#`��zqw�zw���J��|3��C������2C��g�Ɗ��7t0F۞��K>�����#�ar�<��&Bz`0c`#�5�s�2'�hh���b��u��C��,����DyDu��b�z��y�h_w�D~�2FƓ�aW��#��Fyg�T��zG4F����ݖ�<]�����ـ��Q8������I�]i�#J.K	���^�=�-��ʎ|޾��ѽo���6>�����ks]螡����W��Ykh�PL�g���p�ԓry�&��ߐz�Ю������P͇m4�n�;N���ϸ�'�����n��
��{�M��#�]U��+������L�~�^hwڑ��R$Y������6o)f���C���?������^�W����>>o7����1�/]��}��r!���,���h�|�!f��̖4�զ�+L�6.;��S��s�c�|f��Ԍ�{l
���Zt�]�r���8/2rVTj�t��8ٵ�����q+���/V�"n�c-��o(Sn1�L�3m�7��Wg� w�����R��"�u�r�%����`�oc��j�ӦAYa�a�2c
@^h �˕��![Y��Z1��zU �	�H��	�t%�RhQ�W,������WJ�ۢ�٣��=���U��d��Y�������0c��[�5ֹFs�w֛�+�#C��t�p�}�Y�pv��K$����P�D�B�i������gl�L��y�~Q�Z�7�S�ea�а���ʒ
�E�N�b�p]�p�s(49q��n���%�7�bn����#�rE�c�}�˵����J1#w�8tk����d�W�+v��7y� +��(��3�ι�R��i���0�k���w�[e� ��������إdhH�o.�Qm�g-���/�;��w������P����waL����J�Ľ�I@�:`��zOp��sy�A�KJݵk<���Y���GN�.0�) ��Q�k���w\��+������Jl���cchh��Vl���G7u#T&#w�]��e�f��mh��ܹ�C��\GG8����n�
�3 MK��m���#�p�x.nph"�r��c�>���=�-0�^z�"��LS���p����y�d�rVl��==7��n�yQi7�s�ب�<�]�ג+q�'��y��M��U�U]��]���>����\dᥖ��G0 �2R96�L4TK�ŅQY
��.���m���w>�2�m���\�K�g_%�	m���4���$��m1��jѺ����/n�㩾�k�.�F�N���,����h�-ǋ2�`#-;���g����E��0�����N�1b�53:u�r����1AE���\�4u�<4��3J��{/��a	δ%�RL.�|;f�uc���w�Zy}�/&����,c�wi]�.*1�#{,pu?7}np|��Vt��l�iڙYu��$;L�H�����@lf*v��p�dR[͝�8Aô�&�cŷc_hL��WՌw>0l��1%��k��`�7�Sr"����]�>Wd�Ri�o�N��2L��qĩ��7	h^�Ի4滁Z�(��a��W�J%P�uq�sg���e�����"]�"v"��-kl�����%}+D�V��;��5,wL/�HQՔc�#}�^�n�Kuj�b��F ��=��Z�ܮ�=S^nHfY�[[7:L�v]���$��aMӳ/F���_Ĺ���F�5�eo:un����~umđ11�~�h�U�\A�4UEAt�c�h�v0�A�Q�U�����*��y�j����V�:�M�PQ֪�؊���4�h����j*�����j�b�n뱮���v%��:�LS13�MT�&��'���-Q���b*������EF��T`�(���v�Pt�"��ƨ�";��DSTLSDA�b� ��4i����Ǝ�tb&(���������UU�Ľ��A�Z�#�**&)����)�6�h�����7O\1�v�t��B���fj����ݮ�6��V�MqU�Lu݆�u�֒ �&���t3��&٨���b*��#Y6ECI6�QSE@v��tttcjtE�Ӧh����kM�m֊�Ѣ*���Jzu�55QAKT�C��ES0h�L�E��Ѫ**lW����_}�ļ[3�:�N�q�������P�*���>�����*��n�.䋼��X�����~���� ������0��.X�	S�F��|���@&&�1Fo�ʄ�����#������<O��fO7T��DV$;v̶���u��MV�d�3��*�1�|��煮uN�Փ��!���u��z%�j72�C�e�S9/-�[������#�ݮ���񋘀�8��ŗ�x�t�^��ʍ����)9��E6���n�g�߯$�hO�;҉��f����䓾��Q�8t�d[�p&.����QpΣ��Qi�f�֦�k99N��*�]�c�ϭWd��sjܾ��`��\�-}r���D[|��d�T2�盨��~ʍa暐��D��exwsG�U�o�/�Nye�QE��`�5q�2�C�R�X�3����/Uq�DD��K�vT��-ȓ��Hwv�\kd5Y]�E>]�&�}�hvzz.��¼ju�>l��BS۶�M:�L�Ϡ,iD�$�' is�+�s�+�5���Њ�Yx7@�M����,�xCPҨ���g��l���s��Z¿A�]H����^0��{�#K�j�����7��>^�/dg'Bt�"�s=�u;og���A5�Dk��Vo|��%���Շ�/`x_"�[-V޲�q-N<J�>���Sw��䇳X/xSK)�0$�\->
a˅a�&oN�s]##�v��n�Y9wDx�
��(�������ff���
(�������_^z�}�}���<�oP��-8��F�5ygH��&kB�M���A d�9���s����D���S��q��:�8��|�k��`cn�	�a�b�������iQՏ2��;���ͫ����XE���@��f��j�>��L�~c��L�=���f����=g�8�Di9����ъ��K~���s�;�>�D���+��vfD�Xݎ,�w�3���e�����2�΍�3H�t��b���6��Cμ��"�
�l�+)��1�gG���B_i���/�:�	w^�C�*%��RMü�Sp�.ơ��z#�b�U�7XQ$��A��jJb0���f�H탏^��ɶi���P[?G5�_cʙ5����82�ow��L�]��l������K�i�:OM1������1I��O�6�%_s���v"�=�-U���	}�EN�u�����;�E�����b��n�:a'�J|��V/\�#�`mv�ŉ�t����� w�r^�ĳS��H�C.�7�!�{���̢�G�&7>R�Mm���Uۢ�;��͠m�.�V98;�_ی^�P4ެ��S!i�9ʭ�$�pgy��"ۚ%�sYe���C$��K�I��
�̢�����)�2�\y�&���Yұ�m��8�q�t�[���&"�������f�O-U���.W���d�&�!i>=�7�|������ڔ�/��"#z 2��s�*�o�P���\k�����U�!w+��|��^���ln�(1�|��pQ���E�����9�L?d���<$�=�U�3:-Ec�T���tf{��k�g��D�W.���EW�:������_�2X��z�E=�`��6��0���
�g��lp�s�w�͂�����H������,�B��.4����Gs�����scW5���WGi�!�8��hQ�����60fmu΄�isb��H��-�N*�H�c�<%o�CF�^���2�!�˪C�/"���:�^��C���F��A�/�y߅���0��<,�L����P��7�jb֎u;RZ�P�eC�3iy�:����.	�<�#�� ��/_I�1���3R7��g�p��q��'�������i0��P�ӚO����_R�."r
~ƹu%AK�7Q�76�z���lmp����1�ؾ;�m"��D���7(�������"[d6Aa�AQ6�Ιѷ.�OVz��9/l��e����I�l�r&�ud8y�u$�h.=���#��>^/!��
��x���y�N^D�OL���7R�;�է,څ�r���;�v��z,�Ĳ�I��C��Z�����j�Y�a&V9s0�r#���Gֵ&������H��m�#C�F^�N:�B�2Tbkɖ�Ѥ��&b}2��j��� �A�#��G�Hf a���'{�Έ~7i[W��j��\�a��T���>�8^�%�O*8j�<P��k�P��F��#��s�FG��>�Ne��PM�\�D:c��?x__'x3��u[����I��p�Zk�f]j͏m�^�ڄ���۪*4�QVp�55��{����9Y�Ϊ��ֆ��{�������kMS"�R�n#2a�;��ƾ�N�\G(F>?r�^E�o_@w7��E����jm8/�]���9a�*���a��]'��l���SLM�lI*���]�h�7�hm��~���XHM=����.8�*)�:�/�k����k�X�g�?@��4S�n$�w0�����[��<S����v_*v��"�*�:w%��Gk�����CSn�kjsV)vu�04Ix|p����Bi�l�n*-m�)�+ l(�݊,�GǙ���F�+�ک��i�����'{&���.���,��£CEEj޼��略����jK-��kl�F�-���`j���÷o���h.�
j/�*3�yP�_-#����8G�������9�h�:5��x���>�ݘ��{PVjݱ6��h�6#=ڴu2X��I�4
�I2�(���F��pz����Fv�����2搮m�&��1#yrQѼ��Vd�dM�ZI���Sdp]S#��;�>Z{�^�}G�ǿ�����B40���f����X���7޸Sx������ǹ�o�~�FZ��N/y�t|�E5��7ө'ܷ���"{F
�[������v������.dckXхހ'�`��x�Vn��/9�0�:՚n�»��Ȋ�J��-����.1tV;6���iۭ���@�TRp��n�=�S��m�g&�����&�&F��~�&EE9lК�c���h�ݻ��a�;�J�r�a�N9҄��J�_z��X��xn��gu�P��-S�F�N���V��()��TMG���m�:��5�2��1���?[Z����W����nZ�ƈ�T��T���|ǟ<��Q�L.qz��lM	\�����	ִǋ]�2���x�2m������֛��Mi�-�8���3�B�§�Ǟ9!��s�f���~�CH�M��9])��#\�}c�C[���ζN��l�҈��~�6�Uaǘ�i)�0��X�+�۫6x6�إC�:T�{(���[AM��$��C,��r�f�T�[	�&7�䑚��Y఑	4��ؾ�9� ��vv�䨵��TXOE�l%@�o �� ZL�3��O�e�*����2�N��	����Z��n'ʁ8�tE*Z�z�Qt�\n�_��ꊁ�T�@���J��g.����V\C�.�9B���f�Zd���mG��4�g	#��YA�]��eЙQӇmF����u��c���7FS���oxy����1
lp�Oo��a\�o��/���1uϒ�0�O̚}���C9N15���\�u�AkY����̅	��3��wxg����a�q�4�}�Ϣ�R5��E���l�dVq�;#o��}�L�yY���
2Yny��3���kđ��X_>"?��6"���z��0��D�I��.��d�B��x�#�_�Wٳ���5�k
� �����6x�}U���*�eKI�wgC��䢆=���E�8�m�hcRΑR���X�-@��M^r��^�����ް�_`��}yW��g�Q�]��u|c���۬g����c˺
d��}����`����K��S�������LU�lc#/����߁z�r��D��搳�)Dw�b8㚤���j9��:/�9D��l�yS�@�� /����5�X���.���+��O�x�>��N樃�T��?sRkTW�.���bsM���k�7�Nt:wB&��:�2�����.��~���_\�9��3��E���*N�߾�����+ѷ�^̰��:f���P� ��/�i���>#���<�6:ؙn�����ogrlq�3�B�B��۲G�iø�	��"n�5�Ղ���*��+uK�\pP2o��!|���8�nun;c�0�|�����<���s���ƍ]�/r̼�&�Q��s�W):���A�=Z�O�X�m�Z!�OQ:]G��/�y{ �b�#zsRC��1�/��3���w*tr��0w�f�u������1eEl��?X��]�>"e����X>��N	NɜE9fR��,�K1�Z�J�"UL4ĭ�閘�05̡ۈv9�P�d�ښ��!�[}�X��^��|d3Or�\�mۘyZn�Z\���[t�>"�L��݅O�����9��͖�.&q��!�P=��Y�i#��ޏ\�qQ�5ʧ�����Zº`�/1�y:4[�9zb�\�F�	��N��+��Y��s�50���qҙY�P�ݍz�(�\C\"ۿ/�����ǈ2H�i3́����M���a�Svr՟>˾<���.s`T{�8Ь�C�[�	�Y=�1����z`�2I���&�$�~j���>�4���J'�"��c��W�&<�=	����E2���-������\(�O��&�;��`�g\��ok�A�N���{�`�k��!��E�?(�k���i��.�u�Z�9z�S�ʃ����X������<��8�b��%l���mz�d���1>%����y�=������y��JD�,���eΥWP�3����ٻ�w�/"ѷ�����Y3����7����9��μ�u��N|f]sW����� #��Yy��z����g0N�O�L/��M��QtE^	��=���cYR��GW��w9Q���]������Z��g�5�`Cz�pj�2sZr\�&JJ��:q祯��c3"3u��r�^4w� },�;�E���Z�I��w�5�FR�����ꝅ��#V�?�M����S᳻v��5�t�Z�XH��Ր�k���w5�ԯ��V^���Fx��l-�1�Wʩ^֐�q��%CʏMⅅ�ߺ�zL�5vM\##cy�L����	�b�uaD���so��W���)��>��6��q*���l���2��-���b�ض�m��S�f>;�[L9.֠Բ�$錪�8l][4��eW��7�u�犪d\橶����Ow00�uqA�=����*e����+%�j�,�թΆ*�hUy㖦#��\���KwbUm�jN�X�9�^.-�|����ۉU���܄O9r�����݋�Q�y�e������}d�siPm񐒤43��et�H3\ȷZk(��1�o�ɟ:nl̵�wl��N���w�(�z�a�S]6�բ��Xq�\3���׎����8�><,�/��k�y���]��ͺ|^�t�{���F�8� �L���SX�x�}�*���wS�o�'s6HS��K#z}��g�x(����2h:�N�|��"A*�=�b	tY@�sVrZ޲��
p���Opw��62 9wq�0Pg�pTQ�Q3,oZ�{MxX�����a��gc�rN�]�7�6^o�Vl�:{M�v�{`Et�?�yP�j��
�~��r�?1�hW��H6�����L�"�y���V�-p�t��.�[hO�~��.�q�?�;��v ��<��`�_���?�у+_s�����t��b�<jZ�{8C;�xg����������;���Q���L8��l�#׵��\���vc�x��cC�Q|1N��w��@���
ߴY�q���7��u����t���g9X@���u���G\@09��"�7.5��t]�ʖ�����/M¾��
Y!���Փ�r�}͙�0׻Ɲ��A�^+��a����t7w�X��Y�5�z����ց��|0Ӵa���~�����OTX6Oh��V�E)ɝ|wy�2���ң���^�DE|�l|d�o�$��ب���čw��=�|�ԏ�;��ݗ��K�����:
�I�^��Sg�w]n�����WeX���Ŝ5��,��g�3M&M��l�@�!H�E�}��l,����[��d�s��R��d��sL�V�s�Ę钝
�S���k���bvKŚ�;91t�k����en�������׼�#|�Q!��oz �'ք�d� ?NA6.���73+56����[�$-1��v�ף�V=����6�`��(����s�$��]_11�O[]iO��:g��F3����� ��|��S�p��~H�R����Ul1�V�f������Q-:�����ӀgW��W�>�Ϋ�b�z�#����a����$�����odo�X��O���r��et��dO�T^�����h���z�X�>O&m�N_���F���&.:5��(�b`s����l�B^;������$�N�όc�Ն�o����n���)��n�x=����Ni�Hݙ�\���x��VG�R�^��Ϋ�/-�z����"��L0�lyغY���3\k���~����7�������fJ�qui�R����.�>
�<r�
f���x}`�c��
���"2ξq��1�^!����m���N|Ag�"p�F�����q��a�T;���P�c)ށ2Xf�����}>�O�����o������?���eX4�֚�	a��],���+y*}t)��;Ubx�U�H>����Y����Y�b�a׸'W=gGT��l�%�P�܍ז���dٺf6��b��e�4q���U�n)Mg����E��1Y7ݘ�۰r�+{�Z�Pv���􆞍0I�b��ʄ�ǂb�VT�Q�!���I������e���6��ѫ�1PA᫼/i��KE�����#��mi�a���Y���~z�c\�W]�N􂘺U�sB5գ����k�w`����Vk��q�\��J��+�]�b�}��r�e�J8(i�9��-���D�v��
a�fwp5?�}�}����[�!���q�V��U�힦a�b�����>w���B�����f+p�#�W��,�َ�wn��
��v�S˳HJ{���zl&�Ɯ�}Ҷ*h�h[]��_3���p�\����U*��1�rg��U�}�!�c.b�n��U��t��4���v����ӆ�����V,�HZZ8}r'�jCU�f�J�A��Bɭ�[�]�:8��9�կ��e�$u�Ѿ��T��m�_s{"���Z��l��N�xC�u�������)�팶�f����c6B�*G3�u��ucƈ��u������@�o�����ʕ^#�@nq�j����(k�O��=W�_k��ZE�{���S�姠f�$�ܼ������0����[�l�mۦ8�Uq���k��Tn��3
�z�r��'�ij��]r�td�I���-ǽ��9�����9�4�e�.5�ю�4^�Yt$ ]��z����\�v����T_.#�|�n���ܽ�%�Ӹ��`��񾹪ir�:�ݼU9Q'���mt YWj�ׅe����2���h]�;$�]ul2������;�:��Mθ�Y�}Yg�,,[(������`L
��@��N�B�뼧J��GZ�p���p�b�v�܊hʋ\�5�Ś�ZQ�U�Z���
Pe�ܣI+�']+�1�S���������6�TJ�[�چ�m�%z�[�=օ�^\��\�����l�n����a��s�d2_'Z+j��Gz�{
m��7��"*�U�'��;?.��Q9R���e��ųLo����XXj$^���oR�ӷ�2^�1X��wf�9�=b��H�A��0J�a�i��Ϋ6,�}1Va�#n��D{�͚��A�_m۽Zo.R$.�}(-��/�;�1�,v:=�C)��ok�f`i�� �Lms\a������5�F�ވ3Ů���R�1iN�ɕ9]�����Z�w��Y�wJZ��@�d��v�[c�~��̳�H�'^%��EO�W"�oH;T�軷g=�6�Xڡ���J�k�$�M�]y���4�ga�!g	OV�rm=�	�G7��0i+'sz �A�3��=��:�_YY1KR�����W]{ڹ���*�aڴS�pI �|�4R�Q3m����i���(v�k1Z4ک��"(!+E�4TTWA�Thѫj(*��
�U3��jj�������F��QS����j6�]h�(&���&!���b�H��bq���ƱRF�\GF*��U֦��6�F�*
��̝��j�"")�;��nق*+tq��Ѡ�*���b��h�[X(�j����ӭ��Zղ�*�g�*�i�� ��i�j��v����#cE%]֨�&j�(�j��
6�DEtj6�ѫF �`�i����b":h��)� ��t誥b��&J`��H�()�"�����	A5�jj"��(���AU%M���CAMQ3QAMN�j�X:\ALt���mE���4�SEUP�,�R�RE�@U1QAMB�L��A���h�i�l[�$���1��J��ح%$E1RDR_������5�wW�Ȏۯ<ӡ��2Fs[zJ���nZ���sT�ht��6�N�[�Jp��8�˱�C�,��Y���Y�Z��l��(R^wgG�mwo.���yպ�1��X@�-�7mGXR���a2�V��r��b>T9D��	����2k�U����m;k����Z��{{�m��fG:M����������hO\�ﾠ���y��u�!�����N�h��sc������d=�|/9�TG8���j9��|~�bMi�~��Y^f�k{_3)Y�C�:�\�VVmܛ����p�i�d�_s��#��>'�O�:�/_ݎ �/� ����V�˨�Q���)��P��P�/L�~�+�;\�a��bWS/T��a�c!��d?x�R�,p'G��z����R|��U��$�wK�f�ވǊ/B�;9<+�s06j�\t�h�k�0�r���ug����Ͼ(p�K���O���Z��3d#R�_j���\�����^�b���n��m�;����
�ǆ!�\��!��_[Ӷr���|��6it#S��,��Q�T�X�g2c�����磊�qE�������ؒ؞�{��%��i7��XX3	�{QRu��᩺z`��$�ٹ&�=�s^�������C�"{�!�F�6z��6o��Uq�g��<o�׫uV
hu�J�S�}��1-20��T;��1g�fW�9�>�n����{Ҭ��v=U�t��J4Pٙ�]�Y��7i<����0����u$]
5,kKڽ�4��+$Λ�1	�'Q_�>�j�w�2�0�~?kt8�8�яD�	�݆����\��F|����@�8A�g�y��g8LR����!��7A` 	����G�;8ػ�C��-���Q�����N9d\%u6i���F�n��&Q~"3���`�v`́��!���E2���ޢN��O�;�i���a���!/�k>=y���$8w���ă�P8���"�Zo��A�*��}�%s)����j^.�n��1�p"��N^U����_t��0�P�DH�^|ҟT��PU���ٶ�7*ԙw�#1�c9.�cƤIy�@��?m��D�y��I���g�v��D�it5�\@��v�n�.����
`�~7+͡�S�SM	��Ѐs��gB�W��j�����G���
��Y��|j��,�"�tT �i�Kf��ֱ��o��^d���1�|��#G���!]�A���G����%2��|D���Y!6�65��}A}���W��?��٭�^[���}f��q��u��dO�Ot�����E�`T�iU���ևJƚ�������=� ��]��5 �L��Q�ی���NU���y�zzƞ��Y�WW����N��6%�o7\AꬓF�݌Z/#�Q���a�9쵕hV�ugl7),����w�9��c��F��#|�����U����ڤ�!���!w���V	�A@!��Q%�mHr�_���.P/{�L�<���f����,��ʘW���	a{��Z�т^
=�\3�`��ce��A�_wP~�(�y�Jr��J��v{��c~Γ�lL[y���L����^J�2h�m�y�"usdv˷4 �܆@osǯ���q�\P1J�>9�΋��ü���LH�Xݜ>!�MHL�3^���U�)����?�Oͽ@i|�_�"Y_)v�{����Urt�K�z��I����E��4Us�E�nBQ�Z�v�F������>" ���]eQ���Y�Z]��@;�n朻9��蕈߽Ϗ�ׁ��g�n#�9�w�Lh'��P����qbD��gO'\C���z�k-*x�`��Zb�W��|	�֡Ų]�x��2"�?>m�_VI����)�K�b��|S5�yr��6ͮ�}��De	3^�ƥ��P������li���-;��D�?_�\�rwzaT9�T>9�r��\��ּ���{�X�h���@��m��ּd��I���T�7��z\���o1=�;�j%�l�u�[������RU�Z���Av �N���r�H�忬��K���wNn��܈h+Ԯ}i.�]�;�(2�d�c1so%�֩����~���kO^���0 iݮl�cjwT�F��2u���0O�xЈg�`dH緶����'�
;;����n�������6-�r�i�(���8�f��~�T��ْ~�up���x��h�k�|�����\��:���̑g�{��aX����i>A򰱋i3NL�5�q6���sJK<�0�÷G]�{����pW�Rz�K��	_w�ߖ!�J#t!�ʠ�J����H1��S�C�C-��7�l�u@��5�9\)9��\{ؐ��,uYF�i�s4����ۛ~��*���}kʜ[�h���k@��蓏}�Q�����yʅ�XQ��EN7K�*��]��FY.�!��|�h󂢝��L�mdph��0nP��s*��y(����B�Mt�qf�+�x�.`Y윗�A��M<N�b~��Ҟ�xq�����$�=^�}c�9�DbOU{#CTw��A��Gp��!�Ǡv3�80ι�K���-�H��h~��AF�,:�o��۹'vyK+7:]bx�#�Q���q&������{�}Y���z�y(#D���q������d�U�e��l�Y�Da�����_o�U̘9�;�����F��z�7���LW>ۗq���{1K�v�­w7 B��0Sy�n�T,Nev)�?�����IW{��v:�}����»YSc�œw]GilXr�dՋ�Z�λ��1| W�����2�r�4����u�c�4S�V����<#/3�S���Aon�Uʕ����"p��ƣ�����C���K*�@�k�>~����'���ҡ�B!�yӓ��==.��8�%� vz�-�<�i�ŌZq��ֺ܉5X�eՓ˒�1=�z�	��@��$s�6-�c���45P���`cn~E��g�*8������@�`�dC�]��x�u�#b��2b�^�meZz�;}�(���7��v�.���<J��@\
n�BY�4N�|f+MD��J�2��O��<���c͟ջ�O@>u�Up��@P��׹�i];<�\�mQ�u�=�=�a�#��YJQ[�f��������sR2�}�Pܸ��EO�$��urdWܤ㓚��u����){K#"��[,)h��������ɸ�u7��;��(����k������[y�;��׶�?z�Ð����%U�������b�qa��9L���W�
�a���r�(��u�eP�3.#L�fEQ�m���g���(%v�/��!�w5��22��<Ik�#�g�,��:S��Fu,ON��)Pd��r����;c�u�n q��§tc%k�E�k7J_.���u[R��p5�BXݝ�=�Xrc<E��#1r��{%�m�;�4[z4�L4^��/�����wOS?L����ÕP�`�e�L�,��Ekz���w��m�մWчI�(���1
���Y1�4b���;����ɯo�����7Pj�u�<Sw?%��X�1w1���-ꡄ�3�e�=���p�c6ј"�����n�<���y��)��jSr|*S/��>��D���Y={���0ZչCO���t-�Fpt����q��b�(�4e��\��2Y,g�H���Ϭ�UV��eM<�q�f����Ad�?�
�#��A��j=�����V��oF' Z��ƙ�vfM���6��Gk�l�E��"�L�:\A-y�*�#ߗ��tˣ:�{I�C���OI8ݙkf��l��F&;_Z)UM�\c�w�`F�{�>5��`h�ȺA��=r������уq�̴�E��v��7�{��F=I�&��ϫ�'|�꠾�	�<���r�$�{�1{y�ǨWGIn{`�:dl�hw�-�����LXݦ<jD��gR�G�}y�¾��뎎U~Q�!K���Y5	SC�����p�ua�����v��.U���ޓ��C�9E>�ZF�5u�|3]ן����*���t��d���ac�4[N7��w��d�pg2q�c��;�3Z\��#�G�Ik8�ZtB�"ֽx���	�%��u{*�ƻk�̇m���A� oz&.2�+�t����s�I�$��z�壻1��xnA��|F	���c�vg������P�o!(�)m;~{�f�eٯ�x�*�H�ʈ�C%�y��1z�#������}!����/l�37>r�VG5���k�6�/	[�O=#+�.�\����[��\% �ȟ�kF���&�f�,�58܀9[ 4��>��)�{ث�EfX�Y1�@~��X�.��xUB�{}�]'Mf�e-Fz��Ή��'�W�t�e�US"�=�m����`S�\��U�F3{�����uAw��-F|Eɋ���B�dO��{~�/�8�� ܶ׬�6�M�]H��mI~9Vs�YJ�}N0l,��O.���h�	�����&�qa�*)��Q~k]܆Wf�T��C��>��|V�9'�V�?:��t*�z��4ƽ�m�=�X�$�:��o�D�=�����D׷C�e~c�nׇ��|6,�0��fX޵T6�Z���)������;���5x�b�0B���� Cu���g[�n��k�x߽6-�9ޕ�yo�m=qY�o���s��l�~��Ͱ(j$�T�Kdz���L�}y�Jߵu�p'��X�����epO��v�d�٢�����tJ�ԙ}�vP��N������9T��>���,��t(�d�]Z%c��v���I�����y�#��.�+m�\�/P��<�����>��n�<{(ש�T�Lo�'��K�Ǜ�d��c �=Z��ћk������	�00����[^��9|{��s����ƃ��iru�Z1p��v�W5x@���9'�/��͈�Zx6����u\̴c�Й�c5�0���C�:�C�vI�ٸ8Ub�;N6�q:�P~jªل��82��P�e�O����Tf��A)��_��n�+|V��ֻ��~��,v=Z�g����>�9�w�1ќ�~U��55}n�!���3��\B�2�_�ADd��n�,e>[l�:Z̽�1T%K�s���na���z��j+&�2���
.�|�ɯ<Ŏ�ϓ���9���k�m2avx�T�`���H+��-insW�)m�a��,�Ԯ���N��!L9�c�u�i�g��j��.��wO�ίw<CW�A,�T��H��ض��Rw�Z���Y�S������b��c�f-��w�&j�7k��µ�M����P�Ӥ�
�����g�5�׉�z�|�\�]�����G[�Nc�,��jN=��ؘ�������u~%�k������-�6�6���L�rQ@����#LI{���S9��5Dv�Y=kh%���Pl�)�c|B��*�k�{��F=u5�K�`�z�pl��f�M.��ҍ�GSQ��'�Kʉ�oY|]�G�ꓤv&����=;y���u�oW��{�\�����^Π�ȳ�!�}]�N���u!��u��bp�u��2��t��:1>2��;�.9�xʈ܀6c>\�e[����f*��F�Q锄e�z�{_T�q��\�%f=���u����p���s�`�=���k5�C3��J��;^/��t�*!gdq��̄-m�2����w:��P}����G5��3�.E�9˴�������O]����\r�{\�"(hK̪��}oֵz�/!��6|��p��Pg���p���CK���׊�y��O����O*u=�C쵂����F�m�x�=0���A�_i�u�/��� ���8�[��m �5.R$�F�a�+�Q��x��}�������q��6�f�����nΪsA�WV>�Ӓʱ��T7��sd0��h)�.K�K��!���Ռ�z�!4���r/��̗����!��X���5S��ڧ���^jQ�j�xm̓w��Z�R�Wј�況tH�Ҧ�.ǿ<�u�Г/Y�AeO�;�����!��еW3��R��r	�R�Q�&�(ueKW}�/(f���{���ז�z�ˇH���Σ��D���P�S�ɞ#F�ƈ՗�<FT����OL;��>�x�Ʉ�M��i�PF��`L�]p:6kxc�^��J��ĪܮY�7�jC[�)�D����{0�fә�^�O�\�s�ݰJ�F��=nTw���Y�U����͊Z�����us����[�h&�W��WX��9@W�p���)��N��(Xt�m[r�~�����l�b��9�r�RQ����hfW��HX���F�KY��`�[��}�H��2x���\�{=^�W�����}>^�`�{ߏ��߫���Hjs2j#]�'	����W�rpV���i��&5�SBKpoc�x0c=`��%�\��(ӳ�n����K��Z���钷7�#�n_@)����鑃m^��֯�1P3f�8_V�FSuWPP���U�5V�����[�x;hv4^.f�V�B���n��L�%�A0\9[���kVʲua�he���2lp�}��]����V���4!��� �Vի\�sǹÓ���WOv�i�s��`NK;i���k�1��)x�WN#2B,O/i �s���(2e�*��DJ����l(7&�E�^>��azjD�!�}3Q�:�3��U{�U>V����k�;��{Q������Ai��H�fq�%��f>�. �G��/:(͑9��)"�X���)BXf�����u}�ڎ���<)����@rU��Ы��]�Z�	�ty�-/�=�h�d+��Mk�G�t� /�O^^��&��ջ��5�㒑�c�hN�[��A�����������OY��7���
R�swb-os�2mX�J�;��Y\Ol8*�h&�Ǻ�T�:t2uIAnU�7�rr[�9'S���2�)������t��X��Tۥ�h�0���� VZ|� %�{�ծ�o�����M��1���_Vx�d
�]M�r\�G���ʴ4a���[��Ed(��6��es&�JCdy�\1�;�ix�ݜ8N��u��A1���\�\�H�V��S��[����^bH�9W���E�Ȼ�����[\,ڏi�i�r�_H)��w{D�*�L���b]�=�Z��i�S!�ǙG,�rJj��3p��1m��Ep8���ԬͶ�`���h���ʥ2�6�@��!tw�Ċ�q6��F�ȭ�ۚX��\�C�J���1�c��Ԭs Z=gEuui�m����Q�qȮ�vٽ��R��>T��;�����M�0�k�S����On�����7���b��֪�C�[�QPp�)G� ��q�-e6�����.�􌊉��ľ��RS�o����,G��6�7���{�W���P6c��7�_7�s��9bU!�k�v곴�	M�:ȳY֬�j.��A���T��+��HhG���:�j��ǥ�}KVA��V5%�\�:������%�mA�Fb����.9/i�ܾ�K�5e�v(����4"�U�����O����˭1V�b%��oH}MR�䑃��9��[�S0*�QH��쳁��1vV���D�242�e]j�ɿ.�����t��]�֯A`j�2��TۮA�n��U�X�ۚH����U��e�.��R)�WNɛY��j�؉���R�GSq�K���x�����g�}o�5ԾE���\���1���F���D��t�+�_5Nͷ�K�
]}9�m�w}J	k�O0/"�ۗ��X�w��0 G-]٦��x:�8��/5<�B'&(�&Tۋk���GX�j���Ē�I� �����I�A,kEL�ƵQE5QU-Ί6�Q�5��CE$�ADUF�TE&ڊ�	6�PR�S��х�EDQ��h�4��[a�4�`)5�"���	i
J"h���"��ZCE$MLEM@SQPE����PIC#��(�

$���-��Dm�*kF��51D�%��,DE%4�P�QPDPV��l&���������M�F��u����ZH���J5���ѭi���������4��4�S0QE-U5CAAAM0�Q1IU�Z�4�Y�J���bm�$A��ITST4�BU14	Q�4�SMF�C�����vխ-D�PP�,��ff�0w�z��9��|���8��u�����F�A|4�J���2T��{�t��lŝ��p8noSve�r�s�Jt�G�$,>2�F��q�{����r�cϞ�ie���-ܝ%�U�ٮ��?�v�i�߸���R�q��ƚ�����}�k����Ĝm�цS�{V��Z;j�$�^Y(���Z��i������~��uƄ_�J��Q���{��޸�"7��8v>q��e��$%jK��q����Fco��/���D�^����4Ӿ�q7Ɔ����Ż}>�,r��<��e�V�(B�z�Dt�][�;n0YWT�ٺ����3I�	 �����y_1�:&�r�|>ݷhާR:[���*����R)Mz��Tl�>�>f�ҳ}�6�OF�	s��u����V�h�F�2<�p�H{�k�����6��ݍ|��h�]�o�zԝ�fޯ<ŎɈ�PE��i�I�#�^�e���.jq��q�Χ�*�)B��z�G�ժ�*s%;��0��N�g�Ne�\�ƴN8�V�a9�Vc�C��9G��+E����R6�#��^-��^�S�Z,\�2�oK��*�RS�
��D�V���5^�O�Y�#=����we��g)M�nʬZ�Z�&[a�d�D�2��m���8�ATKy�s��t3�T
���U�J�C��M��$<h���:��Y>�j�����򖹽�5s~�2�!��Q���������G�{�ΊaxGw^�w(y��,יlz8lS��ݽ?f���ԗ_�A��VD�D1���!�ێ�����\�m���>��-����	��v�MQ��]�����҃Iw,�N����6F�C�!��=�n��ռ�UG��/L����z���5�Ӟ&v�6X�ٯ���l妻��R��o��f��b��sѱ�hs�,�=}^9ϒ�h9^��F'v��H�xȜ���>an1۔��6n���V�o7i'͹������Y�d��ݬQ�P]zF:1���xuu1Ȫ0�k�@�8ې��*��ik�q�sj_��OuP@�2zw�c�qؖ�����W�ڧt�*z���f�Ԫ�;�Z.Fv������;6nm�=��A5r�'�I&�<=�,�dH8���᳧���8��@09�v��d�����=��>>��(K}�g4��Rܟa���66
�龽�Ɖv7��3oqpe��J3H3&0yA��܏&�2��3ϻ'^3i�p�wF��,[�hFn� "ș��m�ič�u�J��K���
2���!������2��ƛ�ԫ(����+�O!$2R��V�Q�x�+�T~������}&��R8�Soj�;pTLIe�jV�J�
Y;춧�}aw�D�q�F��[bi�xeSlC��r�Zޟ>t��jY Q�jʭ�B�GJ-1�z��'2�jǁVۡi��)�G	ŝCϨ��#�va�h���{�ڇ�ڲa�����lă�R<ِ�{O��_
��`�#ߏ��˩c�=��hd_rc+v��]Y�֢}�},���`���d:)>-��[wϑy���{��x�t�Xnܟq�o�+,���Y�h!7{qh}�>��=���Ⱦ��N~�(�m��{ǜ�eF�(кSƬR���źl��Df#��<�zj��[ky��ݺ�7�={�B�f[���x�\�L�4��4bWCܮCj����p����5��E�������\�yyV��vA�s'$�]�n�՟l�3{;�A��e�y35j����0�
���H�]'\�������R�����Ⱦ40����u��Qv���u=Yݵ]���}��Ꮢ�ڎB��'�;]�ySn�Հ��{0�܌uhoY���3���������q����0U�+����E�a�KU�xh��ѹ[�q;mC�[�6^C���8a�:����̎"��+%��OL��Ҹ�!���t#>�-KQ#|6/��L=Ʒjf FoQ��Z+�.�9ʲ[.�^��JC'�E�~w�����d�W�'���9�Ռd���*j��۹/d�xd�Sk��ϟPk�}����b��� ��l����`��>f�GKG�v�%�4��)�wk/��L�v��~o�jw��5.�R�y��G��w�OPO�ߣv]��R;nҍ�O}�Ҏ����O}O�����/"�"�>�w�Y"
l�d+;M �º|i�/9�F�q~�^�㾵\���S��܁��'�V�3/��?X46Bx��
�̷���X�}�0�|0��F��$#�Rp��`�6���X\��r���[*�=�j-����U�x2jfn��}NTu��V�$v&���X�Y:�T[z4S�b�mVu�y���:㺒�OI;SL��nn_7U;���=��=w~����Ϛ@�?c�)����)�Z�'�^����9>W'�K�o���.;����Vo%D�*�O'V���)�7'K���҇c���:ѳ�v�[������=\����u-V$��2�U�3���|v�&��A��!��}�;��'�q�JQ������]���or�����?���������%�����?�0�ޣ�~�p+پ�-�|6��W�q�yZ�·�^�3�GQ���Z�S��$�P����	��v}�F_s'c
�u��$���2�Ki�T��QD��5|�u�G
�j�#e�X2�ۋds��8X���"�{�h�ʧ-�Z5���Y|)���L?�}Bc���m�/ި|$r�������r���+A���i��o�a�<�p��0Jx�V=|���I�ٕ�y�
���1Lk¦���5���T����o�d{��Y�!�R�n������:���ʎٳ��.
�)��oY�r�;]�B|�Y9����v^5���:�}}D�tݠADgQxr��˴���7��\�+h)Fs�*L�d���>��^9N�e�Ϟ0(���tȫ�%@�8�f�P�N�/��Z܎+�����m?m�7qΗ���;�1�4�sY�/��V4̐l�7��9d0l���(kJ�_,Ǥ�\>���WH���ǳ=�2v���jCu���|�x��K(%���Fh�v��=T��O��C���٭Z[��T.;Y¸��Ժ���wX	V\M�5�j�<Z��,�����e�����ؚ��Y V������M�m��03�nv>d�9-��Rsf1!��%|��f�>�["8lT�f`�&��cB���U�*���n�C�9Ķ����<Vu`F䇞���W�/{]c�s���Q\;g�5M�Ay�6��	wZ��[C]{f��2��AvV$�k�Me��^݇�Jg��b��%\oϨ���ϸ��cޯ�s� k�"�7��d����d�25�c��;D�7WC�u�z�͕�(��rQ����'k*e����/mJIN�(�4���!t�[�:�]Q0���y��"�K�7���w�֣�:쯒ӕ�ھSg!��"f*���x��{���<�]ʺj;��x� @�@����9���E����^�'~s�S��z�{��t�GҬ-�6���C/6�^�&`,3�Y�m�y�z����ɝk8�p��eW�gr����H��~��Š:���U{��7�$:���V�k��ខ�ڣ��i׊.�F:����[FW=�Yn��k��j=99�B�n�:�R�P�
#'HX�;X�N�_Q��@��e�}�ւs/u������9U],�S�|By�����y[�{����Ƃ2a�vC�]uI�v̇�WBWE�/՜Vh�A�+h%s�VJ����f�ӥ߶����6�T�e���5¾��/�����ҎԶ����-۸e��|}��m�q9����c���Ms4
��:�Q=FrX��t3u��ݻ]4Fq�5�Q������Rِ��d-�\��6�ؼ&��u+gO��5=���'-5m�[>A�FM���ah3�T���J�u���tȝ��V޳W�5��y����f$�ގ�*=���imv]�)l����ٜyxEy�f�K�|CJ�\�-��su����k��v���j�ٌ�歰}�wi�"������Gb�]D�����r`��e�0��8*k=vͧ�K�P�j�
���]и�zI;����"`eZ��4SI�0W�3��Mp��B�Dv���iUC���t����T?�u����V�eb�b��[{�.�l�a�Zf �B{s4�"� �]M�ٞ��fZ��V]���mʎ���	>��?���3���F�Jn�`�Z�.Cpڑ3t��v������ߧ���1xO���|ۏq��m1�C���{Ѧ�Mֳ��1沇\��F��fK�s#�,��_/x��Sju�cR�|'"��v��~�8�M��Xȱ]^��n{f[d;����M3���=�k>��Fjx�������o&�)>��*�N�u\v���y{~��[ט�J��@c�hߢk��w���XK�E�Ҧ�׵.�<)�3Q�3(ԕ^�I�U�W�ٹ2f;�{(�bij��X�Q� ̹�q��fպ �D}��S�:s�T�^Mf��Ȍ��XZk^n���*�v(������SV�� !Wr ��e��^�Zu5�ˮup��- y��������:�d��ἕ���Ƚ��Cj�ߕD�M*Z��;�����\TMM��t�?�׹i�w�א�K#�f����+�<p��mS^�=�-��]5�r�%�y���H�\��)]B¼�
��e�%��Cʁw���m��N�)��n�ij�88��H}���r���boV�>M_4U�+���+�/�@�f��;ܡ�M�T�Cõz«y5H���^�n����z�*�C"����ͽ^��]jڍ�bx�h�a�P5K���{^��oZ�$��:H^�I��o��#k(L�׼�}+����t��G���������T��j��ٚNy����<�f�p�m�t�Gn�i��J
�LB�83b�M���I5�x�ň�Z�w�F�>���oX��pE*ڱs�W6�?d���Uq+��h"�!\���� ��c�8#�h�q����C8m|Է�?�a��Hs��.�$��#@U��!�4B���c����#�I��>}+�XigN��]���c�yYr����2�Ԝ���g��d�u�d�M�"���nE��2�e�^'j��Ȯ-݇�mob�p��ۇ�ȭgV4P��TE��lk�wQ��5)��trF��7�g|�<">F�ʇ*�^��|��C
�E����Q�z�KnC�2 m�qbɡې9��_��4��X�K"]�ݛ����c9K����+��e��y��k��TJ򛞹�xD�Y���_�|������M#������+��]f���뻗��9��Gg���k&8�j7v��Qඝ�M:���!�!��˽�l<rxǥb�#��l[m�q]��]���GWͽ[}�n�[Az��s��:g���1�|�6��
�U.�g�P�AM-�������C~�w`w�Vsva�ɒ*��[��Z.IqK7ƄtI�*G�\���1T!�2�v���t��5�Kf�S�V_}zZ5.��:�*]�8˅௙}�qn{�������W�S�U�SC�Y>�W��{���{�ޯO�����{������z|G�sT��cк�|�3]fAG��6<�Z��I�#��^G6&�ֲs [Z�Z�v�tݮ�\�A%L�3�P#'ر���Gl[���j�)�K�x�^�ųxX�ᜑ6$�Φ'wx{8��ol�o�t&�S�e���Peָ�B��Eι�n��$�ҫβJ�`���Ԥ�b%3�0����ň�t�)��Qj�#�z�RBf�G+�z�z�j�;��7�ޑU��E*�ِ�ռ����ջK���}yD���$�e�wG*�u
6�auv7��B�l*���(ճ��d��L�ܙ��r��Q�x�9[WE�WshQ��::�t3�$�G���臗���=��C�ܸ�va��Y]�Knhq��u����n3w����
���s��h\�#/t���&PDZ�.��'&K�m�롘9�D��ӼNV�vI�Ы�ЮC.s�)1�e$B��S��V��%�/^=�`�"�
ޗ����v��좜�[v�#x�.�]
sC�NQ��fmҹf�����Ĵ�tܭ��8{�y6�Ю��1twC@|���7ٖ"���!�gĞ�L��*��}λ�7���+�hi��.�:���a�p;ג����b{SgWT�)��Ҡ;�	-d�c��k���2�pT�jɕ���3�Y�ln��V-�J�K薙W�iZ��w��\�ڰdu���x��X��댡hmm�)��3{�:pʩ0nP�n�=P<���7�\j�&�mbћ����NI۳o8�;�V�.��łn��P(LE�N�-�{�oKRga�����B�)���Wŝ���#MʹO���;7��(��(��+�$���f�8<!]�����pݵkdw7d�,�cTדHܕ�%���|	�ٰV�k���hgPo�0�����뿤K�A���Y�[����]u����j��M��}�d����M�k{Ai�\�`.܍���9�v��7��pa�a�0�,#*�\w;��*�bf!p�ʻ���0&��F�i'��X�ܸ*�(k����g&��`�i�ۧ����j�^�;�y��ҷ���K9-X,�Sr�����Y5��΁]I*����r��hd�Ӫ/��[\��j�dΗ�͍a:P·`05lF��Ѧ~�ۆ�9=7�'u�Ջ$��ZI[����*]ټW����sWN�˻������r�oQx�:OD�c?gS����2�]@]n{ii�sM��)`T�t#�v/�wm2f|mB//�Z�G��蛛.�Ei/,EU�ޜ��U���_V�}O���d_e㺘��*�,����ޅ-�f[�5ase��Rʨ�Y��ae�AT�Zs��%H�__3���晽�m;�mΣ&t
��2�&�olB���'��Z����iS��t�F��p��dIyW�LJ}��j��gf�T�r��qޗ(󙃻y:zQ�*���8�M���?�#-EDQ�M�DE�C�m����1�ДTT�K-��:Zi���E�cKEU%Ui4U�h����V2Q�4h��֔�(�Y��$�h��E[�Ѣ��Z�8��t����[Z&&d �٭1�����L��%��h)MQ�Qh�PDU%F��h1%U��Rlj���Fe)"������ՃAHF��Z�UEP�,E�%RU-4Ѷ-�[�֩����+cQ�`�ӈ"�h��4�R-UQN#KA@T��Ě%QA�h�IDLIUM)��ӧLQF����%% �Q��
Z��Ѡ���(����?\����Z��F�h!�W�-_ES��|9j���wS��t�d]�kT��+�*��*��WSI�Ğ�V�6.�1�8M�ɓ;H}QPͭ����,���ŢB4��Z/������]�5��p	�t�u~1��c�t��uxB.g�ղ�-���W>��k�,������z�R������\�>qn���g��:��.S�sx
w쾄�`,���SUq|��&QّZy�҃�K�c,[K\�l���5pȋ�ǩ�':zi0���] EzN�5rw���V�Erj&7�S^�򸫱��*�k!���\���7�2*c�ȹP_��?%��f�yE�O�8��z𣽾]�lwnf$;h?/m��n��d@Xo0����o_��î�U�tj
�Y{�G��,����9�:���|�`2g��EX����[yc��Q�;W^]^�Ѿ�C�� �Rzu>�lR����D<�b=�Q�yC����{��4�Y�`aݧ�)�A��,���@�N�p��7[eŀ
X���6�s׎��׵�ժO�z���q	��� ��r�x<�Of_P?��`^j�s�DQړ��	/5�R�Y �M�ؙK����	S�VD]
9�/z�X�\�����̛�������ᙍ�������=��jA�#jN��_6.������S�]v+Ǎ����
��͗zP3��W��^�������C9��7����P�W�DTF��)�����W%%~�|f1�Yz��#'wttt\�^[�w��`k��s�H�z�oP�"�g$I�f�l�����O�w���U��s*�T�fK�,4�\�H@���:GV�$���F�J��w����5��q:hY��6��fD�ږ̏9Mr ��2���Rя
��n�"�TwEdH����^e~���eufGnB�������v�lܛ�$eꦯNG7��;�/o�Gu>%�\˷G#�q���	r�\Acn��q2~=�`��N��T��o��=��LI�F�]���s�F:x_0B�$�V�j��Gs3�݃��o2Fįt sUW){�y֙�k >E`�y�q� �Ć������u��{����=?˪;�ׂ?����7Ekq���8���<nOW�YK9��m�6�>�i������Wp�Ͼ�3~���{�����(NrӘo�j�i�GE�0fm&f;�Q8	�Q_e��n��otH_
:�<m�/�z
=��Oq+E'kTq�ꕷ���-�� ̓h���q%[S�d�vom$��nm�F�bt�B�p��T�ʈtTܲ���*�[�c��l*]��7�7�\7���\�״䴎�9^�fA5�ў��a�6s+l�:�zj���R�]ˌ�(VEg)�:�X�9��C�&uҖ��u���.�����Uj����3�S}^�"n�_�x�QI1@����\7k���V4rj�s�e��;�-����WUMna��N�#Lܗ<I�����7G$٨�*��쉧�a�K�KY���1;#֒ס����GT1�qUc�����jm[�t��j�˭�Z�U�Y�ו��$���2���I^+ª��㩼e��6�^�q�G���]�oLdw���7�
��^}�/��JD�%}O~�[*�M.�xY|�!�i��=��֑[m��;�,���MC�3�0�T,��U���3���}�;)���NAS��;�I�{q�;��)RTJ�'��<���t���̢+���xkGS�J�C��'0��DoηX�y��rҒՒ���:�v��nf6fe��8�n<����k1sU]�dY����TyO�G;*��8�Ea�Gw;���EM�yD�+t+;]W���䋗D�û�h�Ï\<��͞^��!�rZ=.�Vv��2���=�����:Z)�Ƞ������>���f	���C�1]s��7|)��L�|�k���=��2r�xn��� �9�;�.��І׳�4dT�!���>`-օ�%�uܭY=z6�S��k����bc�ӓ�rq��췫U��b����N�[oc�6Rp����}Y:�H��=���['�|hm����Y�$��#?w�5Jq���,����k3���|�=����lGF�ݠ�n%3�S����,�|1�<{����n;%i|ŗ-};gXmzx�=�4m�b�0���=�WTs_�5�A�uKn�&���^�3b�%4 ʟh�.WOw��q��~��p�稉�|���9?��8rt΀��E��|2��L�l�Q�=Uh+�W�U��ůŽ���T��X��v9o&�q�&�{�APb�ča��M殎-���e꛻-J�X����X�1-�5A+渾���J����gu:�{� 7<�^ƶA��N�'}TGb��eu�P�?�I9r����ݷ�`�=�}�B9\&J��0�.-Q��f�n9k-a��#�ڱ��mN�"ޫ�"J#�Z>~�þ��Ӻw ���x��.fջ���!���_�b�P`؜�M/>�\��԰���p��ҖZR��]��I;b�E�3d��locv��[ّ7�'Af��E�F�R��s(�T�jȔ�ۭU[06e�Ouj�ל��u�}�w5άG�L��^}{�[�S]q#�������n�(���}���)_l"�[�d;��^e�8TrP��Y�j���}㏷���l]�$;8��+�m��n˞+:�����ڦ�d:��S�Lw]b^��6 ��Z��u���~,ñB�#͏<�S4���٫gD�r*m�v|��fv63����s\�р8u��`n:�^D�Z�ʓ9�f���,�1FDu���������q��F;h���+vi[;蝧^��{]����s�f��=�%�
���yAh�vױ�aZ�:yu�
���F�6v������F[��f���,P��]���mG�g�C���C�	x�+x��'^��JԞ�it�����i���!:��]]�j����3b�\ȗ�adqZ�9Y[��\zvt4`�����.=�挂��v8���u�"���R�Yy6n�E�랑x����#d7-�$X��H/.�a�K�@k��N�jeVŢ�+N^�zjҁ���E��%N�ʝOON��{(��2^�Y�Ȍ7f�ϛU>��s5*Ѱ��
�!E�@*:|��6QM8��>vm�PCgK�D�롺�ꢬ�.�h:����Ӭ���|nvݥʠLX''��جˊ�w:��5��+��P�_�Z�m�S.�����J�I�f�eV�+2���V�d1}4�0SD.���=
�s'��e���q7y�AtoR=�f�7����ِ���3r�2����Ͷ/�sV*���{�@�=C��p=Ov��|�"z��u����mV?[��N{$��|2r����zV�~��Gt�6]$o�ےQ�<���[�m����O���
���l�fp�<h��A��Y�����@4�!�|(X�#Sz�s� \@�7Z1T*���t�TD��t�Xb��$�MQ*ܤ��.�k�'o��ޡ��.D�.Ix�7H�f>���=#�)�E{�+o���﷙u�N��}����`��ɿ���~0����O�q�\lV�T;4��r�[�L�.	jf��q/����x�6�R���g
`��Xp�5��Djy���E^��vU�YQ�'#��<�W@q��u��{X7F�;���*Q�c7�ts;�����s2�ὺ����|��w�<{��yƸ|�إ{[M���{�9�cO@��]�ia��	��R��o�������~��w��W�{��+��Hl��ӗ�^��n�l_G�VH�:�sa4#ˍ���ޚ�'��o�%ps:y?��pz7����r��v^wIE!�!c�%<{�׾r٬��f~�� ��Xe0zA�
�*��3�������&Y�j�����_6����7@�;q���_"|�1U/rf�Ϫ+�c�ִ��z�׃���ۙ�s���+�G$jn��^�{w�t�ǥ��ȷGKT�u�,���ل���V�׊�����h�`Z�:�)v�S��S��v&�n��<%��£���|����i��
]���z,I��uǝ���k,����DVC6�Gv̡FNJ��>���"�W�K����L,Z�g]�1��7�i��|�꡺����j𪩱gM�.��yIB���<K��93F2�^��i�A�s���%"ol�Ws�B:��S�� ���	%��|��J��{�;d�;C��iR4�5�{_W��G�?tE�F�2�S���a��s���~�Y��f�T4��Ʃ��}۴��ܸ7�Sy�A&�AN�r�;���{�}���C�R�c���=�1�[&�j���y�J�V���>YOs���!���Y��J�'FKD7F<��1�]Jz������j�EkKm�� >�o ѡ�e����YUjw����4Ȉ�|��Z��/r��t��yd>�䨁X��V�O6v��ʝ�m�6>��f��������v��9ω����������|+E��l�ؾ�ų��Xc����3���M&����^n|N�P;
]�pu�����m-�S�y���5A[Ǳ�MV�j�ù-�m�%��WII���*�1Nh�i��\J]<��3�&w{%Ay�-=Vy��λ��pF
N�^��x�,V�]��Dd�Z��l��#���W)��
��U���������(���4�$�S���	�_�l@t�e��2.��,��}���Ȁ܁gO�y;PV�>�o�w�Ϛ}��O+t]���W�"�%�Eot�t�D�k����"�b硈f^oQI!�9
[.�e��e�όN�)�l�hj�k�~���!]Hsj�DNi	�r[!Tvj2�KQ�3xCJ��,�����ű��cwD1�:�����s�ἂ���>��V���D5�X&�+ݓY�X=��Us��5�J/^��BY^*R]!W
�u�����&����ޓ���*��d6j~K788ֺ�.�뾉�c��5��Fm�ݹ])6�Qz����ɯ�g����Mj��D\P�m>q�k/ۈ�GVU��r�����6����6g����Cul�{2!��S�ke�t(��N&E���*�u�
���=�O���%iD3V��1��ת[1���^�oIco�*^���i{����H�F�L�DUfVQ�o]�u|lr}��/�j�A&և��6�b=����o;���\�f��ɏ�y�W8�H
�'�u�.�Wd�}4yC���)\�Q`�y���9HA���0�TJ޵t��W�#���Q�'ٮ��O����_�|V���V��ٗ�������F�tMR��'θ�F�Bgc��]Ж_���%S��W�K�D˳�"ŋ�&{wr�[Gc�������d\���:���>3r�{�7$Ɩ#t$��B�d�׵�3�d9����p˺}����bK�ɫl��'m�m��6�����7g4�]r6{&���l�p���sb��6g`j����֞�+bք��v�m{4,@J��1N��V���C3 �Yv]�'Zξ����#��ͫK3!�ۼZADd��k�*u$��\��2��ctS�f��<f�)�-s��Q��S��	����QYuL�Xͽ�0�H79e�D�~���V�|��6�E�:�]2�C�WTT��� �\�'*��j�Sjk�cQ�~ .Qk{��${�>�/O������|��op���І:y�7s�Ȓ�kz=�w�����e�E����2��eab̪�7���4��]��@����fzN
�*�m��K���Aq\���Ԑ$�Y�2���1vĭҼz�dX���v�N��\�
�
�'��X�c6d�0W7J��㲶]�1w�X�m-.k�fG{�*7��j�5�����|��\�u����QY��m+iLKK���p��3�Lg�C;�:���R�����_q�d{r�m�d��{�a�p��X���_};��Zo��[�dtm��٦�3�[��ܫrd'@-OveIt��ne��V뾹Qr}�-D'�$Z���4윷�����z�K�=C����6���hYG]�V�-���d[��:vNb���nL#�hėۻ�i�N�0�J�b<���J�7 �m�,������kA~�!\��.^���B����
�{MU�m� Z���a�(����#r�Xyb�+ݲ���C�o�ڥod_��SnK.��Ky�D��e�m��� {�cq컌K��3�E�XzqoK���f�I���-��u3�}d�m�5�תϛ�!�Z;q��d��Lvp˜�_�\]E�G0H�1�����':�2�[�c.�ti�N�L�Þ����iͧ����qh�ꭖ�v�4qM�T�}Ǔ�;f�c�J��+"�FP}�{ƹ�d-���F<��^�n&���:[��v�M���:ѭ٢hܕ�U�k����Lۙ-���[�KC���ӺK�A4]`�6ؾ����O��ޅ8;dV�tR�Qޮ.�˙]�;f�[�pN�a�550T�e�i�B�����H=��L�*f^&i���b̗�Ld]��Ԡ�[�I��h@��,ī��(�yY���|E�䞾�=d���/��ͻʻ<>��p�k��WWi�Իսx��l���8X�`���/ta����]C��k&7sL��J(�;g�;�]tPT/�e�Ӻ}��������Ħ�ls���Es
��M�5���k�]�n�hט�wd
��홑MH>w0Cp��N�[���0v϶���Hq� a�e%�F��l��x�F�'f��C�ɰ%��� ����	�u̥���[y�gG��H����afh�A��(�ǝ�[Q�5;v(ȶ����|��7��W�����m��\(r⩐6�����wW�n$]\�k��l�[n�j���q��꿌�X2v�z9���M��cN=��Ѯuq�dU;"ñ�	l�`gR�'���޶R�NrغV9!�ʰ�n���wM���-�S��af3��L��ۘ--K��ungwr���&A�m3ߑ6�0)�f�Ϳ���>��=��s�և#uy�;��[���.���4��\*뺾�Bl����ԭ�ͳ�o9B�Y8�N9+t��m��W��xE$�[7��ʤ��õ�'V�$�fܳo2�;��R>��W�HD��IIM,A��"�(H�&6�SKA$�
~�J:�vKBPҕ�Ѡ��i4�c�Mlb���&v�F���ħ@D�WK�IDAIӦI��F;&��C�h(J*��"�۸5�t�Jŭz��]:�CZ�v��݌�#К�mEQ7N�7`�Iմ@���KKEt�hF��٪��݂��Pi4D���1t<F���*��n�P= iu�c�лgF�M&�,Ԕ��-�Ɉ���M wmiN���ԧF�
�5T􁢂�A��������e�"N�%��0QM%A����(b����.��֟7��;����F�_x3�_gCm��3��!h��@�s~�c�+e!?xz�d(d4�����wE����������؛���PI32�k��tq��=�]T�l��Õ����U��\4� AL�˥��y	�i�g�3�у�-��q2�e�����mmq�N�ĖԘ�F2�t{���.ăs���`���LC��,�'��idzW^Tu���0L�6A����?+�oK������]:��5���ſ;=����r]\cwج�R��>sS�~��������~��p~�B�6}=|�sð���&ߪtE��z��wȝ��r��:�-�߅����5 ���1�nf�ٱ�{b���4Q��=ә�Wo;����&�@:��>�oC�C�ڊ���-e/��-�K^[�I|���7�ofX���u���l���i�7�x�CS.43�wUIq�ծ���;c�Z;��́�P����LcM���cN�=��&:�w`���~��=B��/Lwn���q�(z��,��V�b*0fH|��Xi�^�Z�?T��x4EOP��%������LڴuA�p`��3b�6��34.}P�V�ѬMƵ���]�5�Z(��O�ˁM����\W�+ ��n�i��0�I�]�hY�EC�e;�����K-M8���d���C��,���_+������7�t��]M�A��j~�&ݔ��졠�6���jl\�Y��M�5�^���1B�R�r�1W��h��pOv�QR[�T�5�w��b�|�O��YR��S	�y:�5|��s�JØ�o�'=y༫���iF<&z����ϑ�y;1�)�:�q���v�]�N�Ԓ��y!+��Y��Cv�_C�%[u���mo�X�o7t���~Z�>��myx�b���q�mBwu0ꔶ���bpU��ޘ��#q�K[�&ɂ�ȱ[ŤobD2;�{:s�(4�d�m�5�Rj���%Z'�\���jf�k�]���,ћ�k$/z����Y����j�({�-���8�z}�������;�~[ېk6݌MT�ݵNN�wu������⻩"Q�:�dv�[c�Cz��$��Y��0�A�]b����.���$����o&�C"��e��F1l��(�q`;HvN�0�˼_f]�Lƥ��v��Ne斒�����0�z�"�U˦��Q�� L�	��͵2O�ӷ����[s�A��;:_y��M�Wz����%��UB����6�*�AĚ?��YX�Q)D�+�3�;�-c�Z�d>�tؗ����u�*"C��R_�u�"3]����X�.zA[L���pW'܁Ϙ�W-�{ͧ��V�b<X#�z6�@�-�,k��%����Թ=���W"�/\{���h#��o������fl_@�[<�����:�k�\̟X��ٺ�5��}ʆ�7�!�_K�C"�,2"ʱqٽ�6`Ҁ��ݵ7���Cz;���ƓO�[���b���Ep���H˽��cLL�E݁w1�P�Bmm;G�ө-�C�'���C(�nl��,�&/� �����TWO����zByQ�K'+V4Z�{��k�]Y5��{^�@0
:���w�A�7@�\a� �J�$��z��>f-N`N\�l�ׇ�+kٸL�ퟂRU��k�^QjKk��wJ[���eo��Ԟ�{v[��𸚒�Xٕ�2�*+L2���Kk�BU����&�e�����"��M	(V�����S~��t_�?���o|���]��o������H��La�1ܶ�}�3����$Y�朆e'ΗK1�����n*�*����S�\y2�z֯}��>*�'׍*CᖧorY���[���$H�ٌ�΄�`�{}1Esq�O�ᵔ��uT_��K=�MO�d�{�,�r�{��~�0Ӧ�T *�4�M7.4�V�t��uB.d6���3�x������U��k��_]�Q����P�W$��_��qY�y��S��B���<�2�b����os�+=�^�حSZ��u���Yq�/@��EP�E���{� ��y��C�=��F�S; nN�ﳒŚ�c9������3r'b�v�@ߝ�W�^o5y�3��2.Ty�Nݷ�1����>����1�}`�\A��!���2�����72�_x��>3��%�ua��7�����A'�����]���2c�xz�Ҹʩ�#��9]ܡo}C'�i9�⭲|ڻ(.9*��Q��g^��观�CY^�k�^3S��}��ז�f�܆>�J��J�t��w�w\v��	d���ݚ�9C:_^(�A���.S�� ����/��T���T':Y���;�����[٢���=ǥ.wfA5U��t%�n4f�9�{�pi�g5����~Ζ5���n^SN�b�U�%+f�B:D�c8�~�RY㸿U�������@J�E񘛣W|�T��!l�"0���1�	�Tk�RǺ��ٌ#6�N�w��u-�}s�y�*&$�nV[NE��ǎ�v{o��xBC��sVE)w����5�49�.4��g�}A��w5KQ���u���P���;eNw'�c�x�'�K5�^n��%;�,X�n�c��Efm(�c��#�^�Y"��F���Q[S{3sSo� u]�\���_]o�`u.7fȭ�Y�u�M3R���\�>�v�R��Ǚ�P��̻�@CM�(�v�*|L�%��ȍM�׷nv�	�yש�۶�^h���-75��?b�q�dt|�Q�a��;�����!vK?Fc�<I���	l�f1�l�m���Wt}�����2�B��f��1DR7s%Q�O��o�Z�X����-��"a���p��s5���M�D��ib_D��nB����]���J�R	�3�=�J�Q�kr�$���Dd;��`��q���Gw���s�K��wǽ9E�~�u6�ǳ6�k�N�����E-�.�7���χ{y�O�C�\(�l>�Ď묐��h�0��vJ~0{�gV@�͒��~���2Yd��j��Q�� ���"dxn���6�;� ���9M wiʃfK�r�0ɣg5��i��;f�pdƛ8�kO B���Uy����#�1<�4U
n��������fmQTemM�Yx�ȉ�T0eݗ�7x�m%m�8)��e���Ӣ(-wFh��#���SjןN�f�u4�(�~�d% �z3�x�p����V��4�5����_�����m�f����h�u-�r�A3��l��Ӕ3�2��=�W��[𞑨$ ��<ܙы6�]�CΥ�t�z�E�l
[��k֥*���]�xY�J�̬��WR0]��i�j�ڠY"l�!�V�~��묔{��px�1vsʦ���yݳ5��>�f���ȼh�)vO�e��p��i��6���ű�̾6�ǖs)E�4��bM��:c:6�+�΋]lZ����w�(�w�����7{lΘN�j� v0�^P\f��!�][���*v����7���+�#��Tc�e�.�NN����|�A#�g�Y��m��@���C���rF��,3�Xk'�[S�mu<�9��z���䧺T��7����\Y���7���tM��ݮK���<�Ow*#����_8��)׼+�G:��ɟe��'T]�V^l9�A]�Xe�>[o�F�l���ړsW/2��v�z3�s�;�[�o	� ���Ondon���-jm��یea19O[�.g(��4�"3�D(Ȭ�:��`%ϊ�/��
�AH�v׽k���G���>{c̋Wp6��[��H�c��u0�;�=l�?O[3��1o�G���{�^��"�f�+3b�=��3k�m���5Sb�4'�ӈ6�iz�T����v���E�а�YY�)�9�S���PpZ�.�7�@�d��b �I���Ά{�g��{S��T��UJ֐���X��،�����.���˦�y\���4�y%X� �B���w$�F�z#�&:��n���,�^l��k�"�5���/;Sc����VD��8���R�*�C&��]Y̴aL��k��/1�L/n�6㬝ivY����غ����=�������y��Ԑ��Keچ�u;-����Fp��{�(�?u[�!�`�م�UB�ծy��q\�Ү/=���K'k��q��Y�a�3-܌��"��j�VJn��<��S>��@ҙ£4-��M�D�[��1!���C���u]�>����}�5�ozl+��i�x̝���Y��n��]��\o� ̄�ݾ�$�{�k����#q�85N�7q��tVU.��h]c����S�����OlV����a:c�/���]�ճ�M�Q���ƛv�����A�R��(�v�h�-�1Lwc4����~�����M��(y%r���}¶�z8�`3����Z�L�y��,�l��3�~�½�=Bc��/�Ub��޶���'��N��Ð��!Xx�a��ø��G&͐����"5*���ޮ�dF?3��S��ȍǽ�:3��N v���uI����G�j$��޺Ү��r��+�I��S��?�}϶鼥�⣲��]��Je��sb�\��6��n*-E����^�tUxV�ΣC �����`"�u\�oW0�,����:�ksUѡӕ��s�95�����͏?d޿<�Fa�W�x�� �'��ڱ��o�׮�~��z�h�t����3��\2��o�5�Lm����~9�L�"��)@���ﷸ�~����(��s��>3�<�N���uvK5�I����f����n;�	 �Iyt�5ۻ%���hf�v��f���� 6���a�P�љ��H�Q>�b�ϒ�T	�j__3{;1��{��:<��1|�D�H�7�䣥wz�d��丰W#;B�dt�]W�FU��m���ZL��������S|�%ƕ���B
�c������W�JԪ/
ɑj��S.���5 7CI�:�0�Ok23m�8V��,�M{f4�g%|)I6T悳*��y�k��c^����<h�h0�o&�D���ĵ:��XL�b��c��Ĝ��4��;��=�U�bY�y��E�BT���5��-�(q�:���Z_>�ފJauLRցY�h4t<˸�����z�f���h���ݗ؅�N��]�v�f�c�)6�C������8V��9Y�bac;�Q�������L�zU<���ۯ";�j���tv���"�+{|ܗ+/'v�Y��ݖ}�mc�"l��O��[�і�upk�Kf�>�Q�=�i��f~~�뗄c�ЛT�vphyj�dk�;�&׼����YOgD:��EC��{��d3���L��u��=9��e=gI���;���@�*|�Cq�_�He Bޘ����x��m���ǧ[O1ٛ�z8����J̺]}>:��=��g��Z��;�-��ʤfl�R���dF�Ǻ�X��-sY���o�����
����MK�2,��@m,2��$�������)�s׳�nV��b2˫�ʧ�	[ �cw\4�Q�� % P��\��n������ә�Y�{�J
�x��^����ɽ�@}5��B����^���.@2��5�qK/0aݽ��̠�2@� q���Yg���=[��?��^���{��w���� �����/�����?����C��'�x=����8V@� !�a�a�a�eX`e	 �@�V`eY�P�P�@� 0� � � � � ���� �".@a�@0� v� :� ����u�|9 PPP �@@�T �A � �D � � � �D@��!�!�@!�!�@!�@!� !� !� !�  aUa� !�U�@ � �P �UVQ�E� `XeXdXeX`XaX`dY�a�``VJ�`X`XeXe�P!�a�a�a�aVV ��/|��x1�~���TPi� y��&�����?���7���W�g��������@3��'�w������ǟ���?��� ���������QE���
��G��� j~��?�w���� U�����?�����������?�O� ߯��?��o��
�-D��(�4 R�  H ��1  R�0���� J��( I @J��������  @��$As I  A  @B �  @ ��+*�+ B@ ��2��*
�@";�Xo��O�DTQiJ�)����������~A�?@��g���uW��`���C�����O�C?���c���<?'�E ~��!����{�O�T U�P@_����P���"���{�%PW��_�0��{����a��쟀��>���@[��~?���@_����J�������~A���� >�'����h|Q }�0���" *���=���C������L~`X>������>|��>~BO���D U�	�¡��?D��<�� �����~���~���>0`�oD]���}}���?P�~����
�2���\����������>��������QUUQ%)%EHR�UUT�P�E)QB��P�*��UJ�RUT��H��UD�(DD�JT�R��"UT��j�j	P�����TR�������*�%I
"��%RU"��Q"@���
�!!R���J�8�T�R�U"�%IJ%*�)U ��UT��)T�*��R��H�"є�E
R�T%AH����(���TU$�u�  w�SU&��B�h�6�2mmK(�l��F�3J�J٨0��E4U�I���dicUl�+�5��j�1��l5U5l�E�BT�A�  �CC@(�A���B�
(���B�C�С@ �h�ڐu0�4mZ6�[R�R��U*R�[fԊ֒SJ�Pj���QQ����$�*�Q�T-��  eȡ�Z�l���SM$�H�)1�ڛj�M��mU)Fj�[2��U��F�*m�j�Mi��m�B�SmUM�4�5��DT�" �T��\   g:���i�&���V�f��U�5Y�*��̆��4�h��ն�UF�4ckj��E ��e
 M)
*�*�H�	p   3�ي�0� �[lօ( ٥hl��TL� ���	 �c4kP���V��ڪ�*�H
J�h�W   &�Rֱm�4Ih�$�@fX�L���  ��V�f��A�`TZ��$�����YUIUljT()B�.  �
(�iMB@���A[0J� �Tʨ�����j-@�A  e�h�U*�BPKlJ*5�  �,� Z�
 �0  E� @ �L Pl�` h0�@�f �V�*UP�HB��.  �t 5L�@  l�  �ƀj� (+S  ����PC`�A*  �J���lR ��!D��  M�@I�  2�  3#h4 ��@)i� 
���� i`  �� �     E=�b��)F@b�d� b)�IJ��ɀЍ�#��&MLL`���~%*�P6�`&0��4�4�(�M�$d�S'�bhl��jA&��ªP       ��G��NG�������o���]J���8�3��w�y����8���u�y֜���$�oo���s� �����dF�( 
t ��S�@ ��Abv|���c�?̟�C�ê�l
�"�0��Q8F� U!�+�"-�8w_|�kc��Ǘn�QPD\dq�	���!��10�����Yd��c���^zE���.�����j`�����`-&�̊���N����v��j��.���ų]��$l�L$��{��E�x�r���fު��m�+@�U2�j��[�X��4���
CQ�bX����i�J�Ʊ[#XIGXʩ&�5�*f�B�	�VE����-ּ���h�W��n�-��*�!���$Ɂ�cH�y�i	Vu�qɹ��D �c���Q�Fҕ����j�Y�p��L�+�e-�k2aN���
)�9F�mބ��Rr` Mm�ƣ�R�Ŧռ�b�YM��ur#F+qR��6���.C/,�N��P�SS�@�)�l��miN`AE�������LoE�{00°1�91�Hb�$���2=�00�y�pմ�-���am6����h�0��ܬ�r������U���j��J�/a$(a*� f�5��g*�Vj�*�+"�&��׋~��ނQnAaV�f�Y59zA�{Jb��������iޗ�U��gt��AA�޺�K��3��b��ZMn�U)^�@vZ�������̲=��"���ǹm��N�YkeK�T+�Ź.��[ZwU,�FeXU�6�S��I�{n�� ��a��e0o����L6��i�v��m�x�9)Ô�`�
�j�~F����+�ܚ��*^�,�ԛ�B(9�wgF���ۀ��=�B��[2ʺ7B�V-9#b�@V��7�ҹ53b����\ڎ�n�&�7���Ir#NӣJe;�f`���t`���c�Y�wA��ٌI)j����%+vr΍�+)}Ԧ0��v��.S%�1)n �5��W��$ҭ��uc��U�b-����F3[���jz��ģPH���^X�vl�/`�J��4�IV6Jӳ�4�t�{iXۦ�R�U���%-PYG˗��7��9�z�q�l�g
�)�0�^��`E���1v or�R1�˽"�E7V^0V�M�Q��.�KR2��Щ%12����s0�a��R�7r�Vu3W�[{AJ��nX�e�!ii�5�W�e�4�[j��P���l�R#�6�
�������/YN�eb�R�mVnK�M15����h�-|V#ve���z�^$�lq7Z���vJ��J�t��㼳JU���66m��Kanm���ֽZ��ا[,I(���ygcד�t�t{��A��ٍ�m(t����N��9�ֵ�e���2��(k:��K[b	�2(��pS���0܊�[N��ҲT��NA�2�R��5�]�s@7���՜�C3cq�֧2Jp�5�دkQ�֚&�nR02-�*䈜/�7NȜ��8g�]̊��Y��̱-���B=fSL�1�b��VL��c����Mj�w]KWb'��|�!��Ď�T�Nlm��*R��oU=4 l��Q�q�͵vf�PӥM�Ú���!��Ch]֭:t��D�G8ū�,lrX�?\Cj�9�dw+�8�!x-&�nyh�Kl!S1]���V���b��wvwvՈ�1l��	%��ej;4��`?"�/3b�ȭ<���
�v�RMl"�5jf�����g7fZJ[o�x����ά-B��v�ۚ�Ԑ�����Y�ZR���?D��%6Z��k'�^�ּ5e`�H��Jjp�n�v%Su�����X�	ٲN��F�V�E9l�p�n���ܽ9q��n���^�D�+(U��VBu���L��X���ҁZ���:����޴2��K�kn�nU���Nޕ�*�yn�VӇ2A~3%&r<�1�y�h���mL�Fw��-ҙ�a��rj	U��8`3cĨ��tU�@�NV����@^c1bv�*��d�z�-�G(��ӧGTY�d�H-��5Ѡme���1mht'�d *�VYJ�57��m,�%��' ʈlNH\cF��/r�9�����3��2 4Vmj K8����E�X���fV��`����N�\iS-@b�`7=Ilhnj�u^e�	P`��c7w 5h�H��6"b��YЯ����ť�s&��m�h�	R908�Y��v��]��Kk+(���M8�/m���Y�L�K�
�*10������Ս�H�gf��Օyz�ܕ�Ĉ��Xv��p;�2�W��5���B$�7r��t�p�q뺽�ȶ���m$�^��X����)�eAIڪvb+Y*Zbh4��h�f�;V�T��EѽQ�s1���U�{��^*5��Ӧ�� FM߆���֪�D�EVT62��9��4�ѫ��XU-<U���w[gc5�����	6& �5�b����[��)M�l�b����Ck(�����`v���,��-�n��l���m�H��_=ɭ�Ӂ�#�V�,mڧ�!jaE؃6⧗��6�i�X����Q�@o/�q�6���YA���
�ۼv�VR ��Z-QR��X�������b���ڻ��I���5,�-en!��AnJkd�u�6�pb �wWYe�eï���eVe�={P�#��%�n�bÍ���tRЮ��j�0��U�� �C�Ֆ�&�����t���Z��s*���%4$Z.��۷��s��Ϣ�pڨ-`ĪY�\|����1T�OE5�B6�s#5.�b��6P�����tVm�S�B85��Ӗ���A�Vý�vѣKpɈ�hM�`�'l�u�N�	��q�4Oۡ2(���z�L����d,�@^�O�jZ��\{uh�� D�����mr���)�̡Q�F���?�К���	6���%5������m^=�c�ݬ�wR]�q����.����R�m
WR��B���Q�h�`Y�C�V�����@���N۳X��IӢ�RwfH
Ĳ�ӈ4�uܖ�Q̰���X#�1d5F�Ţ���&k��"�^�.�(էq7A*Q�F��]�.��=����[��m�u�ޛ*�6����.��DXZ:��@*'��v����fV�@ 
����X��4��}*Һj���N�+,@�lj��EǠn�Mݚ�[�Y��'�QXI"t���S�/�%,�o���0���J�#Oʇ\ݕ�e!�4���2[��;�]��M�1��-И4��df	Hh�HR�lF���[B��AS��f:�1d"��P6�:�(��6���1I����͘���0DN ������-��v�؇&]��[B�G�J�U���u��x��/��Lm�73V^���oiX�"�W+�5�1�����
`�L�Y���0c���+a2�Za--��#�W���k���!���Rk��0.J��ܰ3�"��b�J��VV�z�br��:B� >)�{�Dh�7r�++�Re�Yx��$��
��z�1mH� ���M�)c�E�ι��"�S��c*�ڏ(��Aa�MF)��wtQ�%���"�����7*k�ؕ�A@Ib��L�L�؂Y݁�B��yN�ڇd�m��kB��YnӸ�я�pjt�$�e�l&��V��
�	LL	"�E�h��0�3ê�N�b�i�2ZZ��lK��8,]I�j�g/q-�0PR�C��M�6U�Z�d9[�|�;n�;0��lBNn�Kr�eX���)]�ܰE%I2��	�Z˩��`�7P��lS��RhA��L�owYHj�Zc2�sP�k]%��!%��n��j�^т�qK��N���ɰ���,_��+&��QoE �`��H@�2n�ۻͤ���@V�t�������j�HFp��f�5�Wz�ܼ�7!�Ulec�-�A$(�Ͱ���f2kDhT�^�p�6����*a(mȨ Y�K*���C�F��;Q��sF��mF�6��/�2�jګ �{�	��H&I�x���L!�f� �4���"zŉ�[m1���ͱ�oT�]�SrVIK�*(��3 	j��$d�*Gu�e,SX�4�����3l�����ò�Ƿ���zYd�XN��M�Ԙ�,u��є���w(]n�)5Yqn�����<Sv�c��E��i��sbґ\�oM����vi�C��F��:��/p`L
�Zn�JHs	��m��+3�T�%\�jf�ҝ.�ƪ&��g[����^:�B�++X�]��!lb�6�YcT��L�th�(!���	��$���v�Ú�֋AV�4H7]��I�m�%�M�+i��n���[N$�,��ӭi	Ֆ��+@PL��%Y�pU��+���(u��t_���3t�R-S)��B�A���4�M0Q(�A�7%X���3/6R�텥((�42�e56��"dcp�Q�b�g+U��r��+u���S(k*�f������Jz�,��V��"b[�+j5�^��=���^7��:���X7vQ�Y2�ym�K:�:��������4*3S��[���t-
Ծ��և�"�V��t�qeԧw�ѻr��"j��Cٌ)��Mj6��b�?aȄv��x�ʒҶ��I�S]��iX�f^!	ì
OB����1��k�ʛx�ec�@�}�����l�5����:2�(Z���+�̛�Y�`����kn ʆ�̢.]�U4*�SMni0Շpݐ��i�	"�Z�љL0-XGZܕ�E&�t��)Xy�ۍPt�֪ZyZs�t�b�{�!�c�S7B�.�O/m��Y1�/���r��,A̡x��Ί~�����)Cp��X�%e2w\7u������5��=[%=��	ڇh@���pP�I�޷�e�gqf�P�E����yNmKu�-Ӛ�T9t�+���c��e�2��F�Pe�#5���$#X��lտ�Į)NJ8j�2w>c
;�\�D�������������q+��u��-���.M�
�]�[{ �Q�բ��pay�P�1�,Z^%��m`�
ҦJ�u�J��] j��
�E�d	B�spL������R��-'i�d�t�On�Z5p:X�mL,��+0��^���(#	�i
���wQP`�������b�A�]M�5U��[a�Mh��m`1eK*�e�QR�VkaR�r�i!�Ĩ��	"�a��_��������S�ƃI�" �v�a�b�fQ��BѲ�*�!8)�(����x�n��4˼&��!�ynTk[Ae������8�ǖ�	QD�M�K�h�����ն�*yw�Hn�����/@�٠�A ��Ƞ�*7G~�p�H�y{J�N؄����3ou�Xb1����3Fu��Īm�Vd�2R�3o.V�zn3�'$U�����ch���!�h&����%X��`�[nT`f1�nC���0ڵ�JWQS5>ъ*�[�e�D]e�J���F�xuM
v�Y7Bֶ!��M��{v��l���ܽV��}h����zD��5#GF#)eл�!NM��^����j�5��i:f���Y�CV� ���L��Oln�0����%�o>qn�MРu�
�4Wkٹo ���ay�5���:a����6�krZ;�t��7%"rٰ��Tec�r��f���f1jS����"SC]�P���[�D�T[$Al�$����ڠjl�V�	���9׵2�e�E�J+�.:tl�A�4�������O� ��8��2kHӂ�m��֮^�It�����daS�+P�Ĝ���V�:
� ��n�֢��a��^�%����Tr����Ĥ��m�U�%v�eU�In��1��&��[�Ժ6֪���ט�6�
r���܇&7��$c_���R�����b��3@�� N�N���]9��������sP1i����޹C+A%�n��	�g*���)P h��E��p��ɮ
ס�OJЭA��&�$��U�qi-n�a���Qn,)�-Rϱޡغ��[���Y.���Wj�D���.U���u����D�J6F��ؾ&�k{A����T�k2�55͗����e��CG�(�'�ki`����VA��p��VBn�V�)K��fk�͗X�#�K���7B:�F�����-p|�f��`ࠛe�N����i��V�� /�P[k,3Lf3X�ڵ	t�i�@-�3H�kNm��m5-��J��t%�ɚQ!��LS%K۹f�^5�Jc�7n=;�\X�kwS�Y�"r��6�n�W �e�M��X�ͽ��%��5�Z� L,YA8�[V$���)��-����j��L�Ad.�=y�(9g(<���0��M���My@�V�*�����Z4��-6 i��	l�`k�o-�����m̙�wM6P�����İ�V�.�ґ�t�-���Θ�b��LB�ޅ��{Z�[ie�0��;��K�WX0F���X����P�+��(u���cX��򣹛�a�5�kA��Y�@kCr=�}&m6 �ۭ�_&v�HD�bӬxN��ua�:���l����B����v�o���	*
g���tց�unEV2�2��Ir1/Y��<��Y�q�:*c�$��1Y�^��mmki�խp�N�cl�11zPq�W�P5�7�Q�)-�R�����*2B��#���b5�����Cڡ��q��m�gq��6�t([��/<a1bxx;U�Į��[�&����
q��]�+�"��Ռ:�`ƪ���M�S+�ڎhml��訋��g�^��A5��}���L�=�.&GoqU�8;���Z�� ){2�T#��t�X�}�i��m�J��qXE,��$��bD�����h�2�#pi��I�{SC&'*�(1QY��woP�F�����1l�Y"�su�6x�p<�,t"�׬�W3�v_X����ݷt^\pv8��תZ�ޭ��@��I��|��w!�����e�(
s��s�&a���;Z6��wnVe�cI���%q�M<��)���t�q�|C=��#�u��"��Y[N�WP�(��n�+�� � �qefha�(L4L���󘔚�e!U��3u����̺�B]D.P��;]���y��F��	�5��6�7�}��O��s���[�W	�'#%�fҷW[�w����wll��nZ��{}W���3x�BjZE_=��y!ġY ��/�g�5����l�z���K���2(N�q`Wf�u�H�v9�|��QW"�׵C,�����)�䬼+�f�� 3* ����D�H�ϯ�J����(ݩ��i�����5,I�t�N��l�	!��1wYڱ��^�1wjd@̼u�*�����
<���Ś>��8ؗW/��\�U���a��y���A�z�#7pI����Wʯ$es��^J���fwVV�$:Y�m>����]���-��r���ed��|M�{8��R+�v]����o{��t�(��i�uz9S�4��N�S��M}c��o�3�eޭ1dʵ&�f1@��M�f}�vë�s]�[�	��pL��6�)N̙��'���_�bS�._l�F������'�9���VSZ'��wX\Y�A� Ӓ�l��D��}P;MwbZ�b+�QM�������j�K�(LnK���&�ܥ��%��9��
�����ٛ�{���!�k��z��u�k��Rݞ�ư[t��p��NHjho�W>8�g@D��d��$`�Xz�.��ҏ
6R�����
��ECY@nB6G-vo$�욧a7}���b�:�W�M�3�,�mrǉL�[����mS˴�`��� )^_k݋2i}B�F^'����mfT�h=�b�)pf��C������h��V�Z����邢d,��*��x��Ʈ�T�\��!�����mt(��y���أ٘#��w����Efq"L%��>����LB�JC�U�JwW01�x�� �:�+��C�'R_*td�K�v�$k_H{9���F��2wţWf��@^�1,p�Xy�J�[�cr��)b�k�p�8U�e��4naJe,�z�U��`1��A;MW7ϳ�ؾ]��>�m&�% ��� A׺ ��x�^99���Q�E�._Z��n�$�ډ�.�|��:	
�si�m]�"��m��a�w�Fi)	����}�*��B��(��Y��ح�ν^��+�]ƽ�Y�q�g�G��P*����V��p��ځF��W�&m3S�*U�]�y6�yŠV�l�j��1J����cE��w�wO����%��ub�ٲg6�5"[�SLVЫ{k*(����G�M��Je��*�N�kNk]!B�IХ����;0����+�,S�uT��`��pB�	N{]�СC1����P���:�QN�n*�������*{(��%�u�ͮ4����Ǆ�381�xA(�	:��c�6�oY���Q\r)�c{��>�Ov)�v_=�`�/�JO�wǘ��'p�+�q�Zmoi���HR�.\����w���&v�?̫�K�\��qZ,���|�5��o�t��'��]���R�bVl��0��C5�Yӟns����	��=I�Ze[�"�B�Kj(:�`��T]=O7Y{�ࡁA������S�ll��L�]��o]�;�v�k��^�B�ͤz�^�|����<
��HWg;�����Ă]��]h(�����n7:u]�<o6��T��|AS�I��p;F	V�����a�\&�rt�.��H����������4�$.������ޙC\A�VU��sTR(j��\ѬxvV�`�������yJ���u�J햒5�9�p6�`{�ҡǋ��˻��(P�r��%м��\a�B�ڍE��!g^�!W;�X�/(���ꂠ����`�E�6��LmL�F:a�8�i�1��y��19v��4��U���y�̕��H�R�����C}�!jx,��Z�ޚ���(�ϓ�{Q�.�B=�Q��)w����`N� 7"�5a�F���p���#]z>��Mq����t]��ڊ�U�c#?D~ef��Q�wu��:�eA�jT#Z�짹V��V[av-5ֲ�<n��Җ�
P]Bã]R�����6T�d'H��N�Bkhᵡ2�V���iNMW4�2G��s��#Kk���:�F+=gvѧ�<=ע77kWQ����K(�cd�J���S�+��Eࣷ{6^m+��5���Ɖ�L��<�<��W��+��{]�40�
�I�<�\*8�V�U�{�#�����w��+�A*��]m��>�*k�@pǇo�`��bP�ohWIC�<�Xs]���I���E����u��);oVܬ9՝9�AQj��/xK�'-\�ݳ��I�;uU��]�q��*�oy4���C.E z�̘#�y�����w��Tս�8* k���gZeh��a�����0W.X+�l�L"��j��	�ӽ��ԗlZ�okVJ�&���mZ�KM�\!u��Euo�����u$�B	����a�0���L������:wb��eTH9ZL�o��:^w�S�XD�!�I��R?h�dw0r���}��0�����}D���6В�v!�]�P'a:�gov��J���]��QU6��Ԅo0(��s��ݻ�U51+��W��>�x�.��P⦣�[����̰a�@��yW]�u��K�,t�����
�������=J�e.T��E�5yj�N��8�Т�E'�S$v��mv�����W}0�25����*ŴƝ�dIպ��r����W��U��+�\=����LuӺ�.u5�+�[����)�(�a��k4Rzm���&!z��$8�5�]_ˑ�D��s�ͷ)��"�=��>�Ku���@�D+��/;�ݔVT��e�̫x�kgPP��k��zq�S��eB�s�P,�O�R-���Z�]g���m��	���v�R��nEǋ\�=u)�pHM��u�&����@gE�q���V/����*n��B��wW,R閲nH��ݑ�G�����J�0�3am	�A�g"[X�5�33,8����s4A��p��\m�$�mټ��4�ʲZɋlo��J�ݲ��hץɔ��{�2�LU�u�5�LWh([�0*�Vb��e'Sr�#o0��G�\��\9����N���z1��:5D1�����2�k(�z�^��J��nXY�X4�Fn��VvQ�o�]r=B���|#`j6������6v��	ցYv��k�z��Q�K��J܈W&��ǎ��˱^7��3\X�I���;�ݟ�N��m��j���D���x���a_H�ub�����Ǥ��fl�Y����)�M�Ľ�Ӭ��(�ƕgbª�j�ڈ&0+��:��ߝb��lrڣl����r�Ӥf�M'pRꅋ����:CF�K �����U���l����]�]��y���������&���+�.�_O�AK�ӾT���z���GNi��SBT��G8�	����(���6n*�:��FeKPՍցB�����X�;�&�j�Ӑ}��V�35������^Jӯ�
�ev���f�a.3J�l�R=��ҳ�ٜ�T���l�غ��[K��C���\.>����r�J�EI�U��H��F�ѐ5K��y�Vѫ��i�Ql���
n����[0i]�FdU�0,���v�I��Ƿ�~S/��t�.㇬�q�gM�G_6"�ٽ�쵶��}IT��F��b�NچE�FT�|3;fN��:u���um�x��PƵ����6�s�nm.�L�9��^�):S`.z�Nʆpx�f�N�7J����,�01�O��9�k�7\ڲۦja^I�d%�8(5B�h��!�`3e,��Yzh �	)`�X}B�W��#K6�A�V�Eg>3k�]����v^�Em�
rꇶ�;R�ʶ��9MŽ:n�v40^ԗ|��$NA+�ZBoT~Ǿ��}��Io�ّ���'��ޣ���ځS�**p��wk�OWc�
���y�hS)�B�fU��A{
ܷX�:n�[w���v���828*��n�#L-��ꕘ��n���À4��M���{'q�Rv;}���z:�G�r�=�j��VG5����\%��wT�H_[W��1\/��[VۇP�TYׇ������,��_�cUMr�¹�	������B3w�\Y��eN��F���Nk���z #�'(�sV��
J��Lꕯ��{5wYڲ���xN4 j\K-���}y�]��
��h
r�Frnw<n�)��2��Zm)�&�+8�P۬�2���ƕC+\Zi%��)�'XO)b<��'u�_��7�'2��O-_U�g(*::`�Q�z�p�G`��"����m�jej9�J	p�T�遝ێNf�����R���R������=���ǝ��u�N��2�1��\5v��.�08�pB�\٫���)u�Ԣ�7%.��^ٓ�GTf�����j�+OK��mfV�Ӓ	��K��ۓi��գ,���U���go[e��lM��v���&d����C5�wR��0����k7j�k�������u�J���g�t�0�Q�YG�R/X��D�[6ɾOX��= �oqPXGX��+8ќ4M�L����p��m�#�ul��nS�q?Eg�n�rf�����	���"n��haYFov�Uv[�����>��0.�5���{�h�|�Wv�m��\������J������ek��*'Tv:���Р�w�W�m���:���:��ݵ|1[-汢M�Yt�;,S�!�1�)�[`X9�=�;�iW\p�� ��[@�d�l'7����x�9�j�y`;��ݫ}e5]�ep� c[�f���igUsT��/"�¨t��QA�6�Nd�D
�Rvn@a�I[����� eʽ2m�'m1k)�<�v�; �윯��}/V�ARG����k.� �u(�����m�P�{���䩭��]���@�	���SPp�⮌m���`m��*[�4=VQcR�"�n�!��iD1�s���:Z��o6�$s+5��ZR��ҍ����� !�s���-nT䤣��6�"f�b�Rb�%m��V�t��w�O1�:�\�y�0��ݢ�C�������֨Q� ���=d<�8,���٩�e��1��r�}��E{��%gLh ";x̦]�9���~��S�J�!G���^ל@�Qy�j�g+�Ŏn��*Ɔ
��k�w��1vE�D:R�I.�EN̨,��[;���9�f�$����1��oFQx�Jm�"�tS����4�ҕ۷W}IҌ�6�#�<��r�ζ���AR�O|\=C�斸tF�h��W�J�o$F��ѩW��J��� D��g��G{]^�ӣʋ��\}|��n���
:�<mlw}��A5�q�Y�V���� ��k�o���0)���3[\��m��L��Զfo�B��j�Q�٥�=�k���yAep�Zv�
yVZw����Y��u *b
����5;�]��r����i8�u��rZ/P�𣧱�D�W�A3�l�W�SW�쒷���A�B	׭�V�{�䲥���7�5��7w��6[�bE�C��^)������R]�D����1o�K�R��*��I�S6��3�i��jU�<w��1���Y��m�(�J�|-R��(��o8L�XA]��Ɏ�I�nY����֭ɖk8�V71�շ[G8���h�D�p�6��nZ&*`�Fe��q���	-v�����y�_[y�q�W����-��c�!��ƢҚ9Άc=C{�Vu%�X�u�~�"���B�=��۝�3�s�N���V���O��84�'v�=�CQ*C��f�Ҟ�vRYw��v���3�S|`Y��v�\Y�2�vT#��^����2��'�N���L�U�t�2��HP]��E�� ���(�Ky<ˆQ�vb�K�3Y���8vPc~%��������d9�t�˫����mqb�c\F�zw�!*4PZ9;,Q�{�@o"�t�N�A
�$e�8�(��cJ� PSڠ�Hż���il�7F�_hk1fl�[�� ���p���UjNe�gǇT���D&�-SPR��ԺXȚ��o����ec>n`ˡ'*�@:0:J�TG3c�bg&~��f��9x�{�읍cy\8d����0��a��N�~� ���S(2�c20"f��ro��'.����v1�4�M4��p ""�ԐR�����.��D@�LN� ��'y&��#=���a���F#�t>�e^0�qư_��n
�I�N�-���Wz+k^v���R�ϝ���t\2n׌6f�p}�O�h�&ƫ��t��fv�{���Q�Ն�-ݎ�����d����h�_L�/Tˢ-*1
T�u0��S��i HE���N�q�������WW5����6���6uoEH,̡��.uNyɥEK�@��qt���̊�n�w2��o\��<��m>�y���ʱZ����
ۼ[sX��yI|�إ�+�yv�A�Ɔּ�VV���uټ�3�m	��h�*�}��+v�De�惲wh�<��:�3Ѽ�@�̫��5��o�ٷM�O�V�X�P��#�m>��ɡ
z�n��:q����t͠(��L����v�z�ƍ �CV��}q�8e]���;Lݣg����N[�G*Ӷ_p�n��\��e�\�:4�7��.�X�v"����"�K�&++eph�,hWH�ݧm[`և��6���vl����9��9O
��c��7�r�M��a�wu��$��S�ۅj[�8{ѫ97��2��A!�Ӗ/o��A���Ø�����eڅK��Ԓh� ��:p���x����s�)�ق�>4���&���Of�����|��򻄡�Ni��sE�ʜR���s&����qi'D�<�PݠqR�2ʖ�K;^5�Y�0]ɌL!8ս��9���jm�F�a��#v9�֕h�/D1[YE<k��s�b����N	ب���/kآ�n�e�9M-B)`����mAg]�-Y}Q��E]�6�a��Y��2港���S��7o�l;tv��YA�nӡ5�e���
r��s������h���Ri\E��Ek\9dJ\}� �ͻUg{�U�Ư9G{�!���^Wos� T�cTEh�!C,bV7�5����GYL_�D+W�\*���Uu��!��+S�Y(Z�3`Z{�#�m��Z{NX���j�c�X���y�*���X;W�|xV�R�i�۵9���W�xy�J��q6/7���5��[��1�ʉ���,U�Am�6��M�6��=�P�)�fP߀��(�&Xܭ�*���b�Н]B0��v��t����:е�؋a,�mǋ�*�2�e�jCEZ��{0�qn�U����4�e��sXfD~�C��^N��8;�]���v,�|x���'Qdoer,N^�'5ķ�떜���2��]̗F�����Y�f��e�.�
PSe��=Kat�b��>��#<�U�-Q,Z���|���Z�M*�������\u���\�Q�U'��|��)ʾg�P�W���d�NE։����x��9�t�%��]�<kgi�z�b]��x�F(�&�]ڵ:E-���3����e��Y��6 8	�gج[9�.�p�p�C9�r��~��1����G����]�y�d�I�Y��t�s�;Z���PѨӠepX��u��PߜT+w��۶���#��7�Ι��k���|3�ɴ)bjKLDI��Ve�vp�u�B�@eԻc1�L�f��t��kh��bVD@9׺�TP�ݏɛj�њ�E��٥�S�k�\loau�ME�ԏ����wn��q����;N�CUʊ�j�3U�{�u��jH�K7M����tn�q��eY��/킔���,�����j��3n�_"��P{Ix�%8����v�B����.���h��)��JJ��jdG��q[�7���Zn�+�� VOj�{]|Ʃ�û"/5����-<�ڻ���Q%]�^��J͛y��5�(`��cdi�Fƻ|�tո2T���ȍ��V�g ������}�ѳدNL�6�.�OV0��NÓi��vc^Z�S��tc�e�[���2�VX|��M�\��ө��qm$������R4w���<ܾ�m��+�]����s�(��'F��+j�`J�#���{W�������}/yv֥W��YǄI�1$���u�b�A;�҂��pB��V+ s�7/��y�d�]�p���h�.���ce�.ج�W��٫,G8μ*���h�]z���w7plkpdm��KX�]!��un�a<�FUԽ37�3�[}Z�WB,���Rˬ]/��+\��oo��ļ#`餹T�Ԇ���d��RujHenJ{Zf��4�Z�A9�f�������׫tp��P2��"Ջq�57����c$>�Չ]SzUƐѧ`����f�	�u�P`��&�SHE-��g���!����s��f��J�hT���ٶ�UY|�՚^]:���U���Yte�Z�tQk��\��fs�',0�3ON��塮$.��{���;zӖ�⋆:�ȳe�*�H@e?�WEt��K��
���c�rv�-�⫌Q�jK�Kb`�_c�uժ����ӈ��_=��+q�NJ6&1�l�~Ou�e��(�]�L���>�j�"1�E,Τ��U�6����kC��!����7�(�MXP!]˧�r����E�(66:v7fsv�gG���w�+�Q�hn���]Jޭ�4;:B/2���2�]��#GK�������4q�yDH��2��a�{�l܊]X��Q<�[YKh��z�u�;��e�6�(�;�l���;�M��@�e�\�ι����um�k2��b����Yy�2�:�kzr}�u�;FVp�;i�P[� ǝ[���Xl�[��su�Z�ذ̃QCT=��\�F�.-�Ŭ���ښ��[}� �~�}�������yU�W[�bsHb�4������-΂7ח
��8Ь����2ִ54پ���4�������C,vjY���pR�3>Fg*�o$n��5�C����~ː���	Q_te�}��ŜV%�x��6(���nh�w��evK�:��]]ºu�w\k_�t�hչ��%*j�XjR۩���j��v��ꇎ+g����Yx���v%�r\r�.
��Θ�`N���SOs��N��k2������
/���<}|�V
�|�g٩W>�8�U��)KtN�Ia�0(�n��ޗP+�L�T�ic�)u��8���Eƣ������u�BIy��{������,ю$s�խ
���N�!�y���g7��9gd$qh���n�7��kmb�/��َ��'iaݛ�Z�`���Ѷ��s4[�Lz� �up�]�G3�b{���]P-��򆵻�B�ǋ�<Y��d�g���=���C�:<�7���+xd׶o"��Jy�ˣ���a<rP����'{�Ρ���ܩ#Y�h���ƮR�)N�`��.�⡙˩�Z��]��֭�j����.�]Ç8�N���q��(9L^���W�Y�U��g]�tl__[�g���]*�xV�6����-Փ�tB�|V8V�7Cv��Z�����}�3A���x����W��vţ��V����S��9��[��Z1�N�s뭛k%��t#+P/������\6ň��ԟC�na}W��f�䔲@�c�ʾ,�%
�J�vkԞӘI��i�m��L*y�N��za����a���*�"9tL�+�o
[u0=�)KѠ��$m�-���/1�,^��z�K����be���ٕ�]*2��p���N�Ud������P�����G9E�|��E�%%��7ڋ�̢)*[G�Y۰�����h&Κz�������:.3�<�ڏ3/6蛣�1��炏n7��	i9��X��5���l��2��+gl,���h�d�gu�+!��K�K���-�@�Et���QqWSQ�Da��_j�{y{�au�l�)΢�h5L�u|�"��L��ՁsR� v�u��Hz��v�Y*i2��b���%�.�}�9jT�0{v�#gf.��>�kqR�����V�'T���쥈*%ܰ����W,
�Xݽ�g�.o�1��5�D{.�iš���M��G���ށ��R5��5�ݽ�P[� *
��V@���ݚ��Xx������*�0����L��\����Vc9��i���|���6r��o�ή�rΧn����/V�ML��>�eO�GMo;�bj�&��$SY1�[c3+��e
R��{��ZG=�{��e��MP�=�6U��va���
z\t�݌�*+�h���.V3�L��B�tl
�b�+w�bɡ����s痷O ك�ވں�B�[�pXou͇�
��2(�n!��o�ז�J.��\~�1�k7uӰx]�E�(ް1�N�s�"�8^.����!��)����\��U��+=:�tb�Yav6��!��A\;j�V٣S���J�B��U���-ڭ�2�r�%f^V����ם�3YgHҀ<z��ܥ)-&�c�<#QHL��n��K�M����\!�]-vu9!5�;�����d�i���jzR�\�
�+�Y��S�2�� ��b��a�Rڨ�5�Ø�3z��@�����aC�'£Wqu�&Hy�lC�}��o�]u9�q����nv����:g�"�i���+�.\��sw�y�9$R���{P��ݍ�E���c�o]#7��y��,ъ�=yV�-'�yP�@�Z���qf��_J��a�b$�AB��*���h]_�d�s�;��b���[���U�5�(ͮ�)���e#��Ŵ�3�hm-��t���Gk{q[�a��W���ԹaM�R��9Ɇ���(r[YiJ֞�C�{��v��:�B_gRl�6F�%��:ߥ��70�$�Ѝ���A�����dj���x����+ʎ}�ݡ������6��q��Mt3k8K�Y���y��\�yМ���F�\��1�BSwv�g>݇v�vf�w�H�ޮ�+w)QS*��]J԰�t�a]ˠ�ͽ�](�+ >Dn��9*u�Z78��ڥ�s������ّ�wRٳHh��Pӱ�Y{-��eU�Z�Y��'���ksp��\xn��j�mS|���r�Eq��z�tz�Z-L�c@�/�C��fӥ(�eM�������d��0�u�)��Nr�fEF�	�"vkx3�&�oP[�G'\Sl)���W*Ӷ�#�Gu-!�yu�J���gX,#x���h��6�ӳ���qz�&�X�5 /��Ɇ��� \�m���:�t�hd�Y���m�K-V�IX�,���B��V�?���2�K���p�M�#��jR��WR9fvq:��7Yd�ǁfT�;v�K�3n��P�i�jfң
���ݴ�z����5�vwç@�:��5��5g0�YVd�)q��ւ�/d��{� rd=J�8���$�z6��S���1v�Ջ�^��q�}Iξ�jP*���C��X��_&;U���Ɗ�+8��4�Y�pj���n�w	w�κ�$�r��-wKc�"�SL����_ܤ3�])>ڽ"�Ŝ򫷛�k}z�MYƯaQd�nYUc2�.�t�<�δ����U��Ӵ�-��G6�a�UPsUu��uw
�"M���h�=�8�uq� �2��������u}k$0�pU��lդ-P���-5z���*ՙe��W�ق�ս�ܯ�`.�W�7k���-���L'p��Q@�%�}������A�d�"̛�勽j|����>wm�ںYPi�����)�	�tp��M�r7��"�u��K���}��%M��$�v���J`wrP�U�lm��I���[��Ru#�9�n��:���E-�S�Y�����钌�r�|:���Y2ܧ�ћu��a͹��9SLL�(.�3��e�Z����+՞����s�`���ń*�l����Ɛ7��e�sh6p��x���U��B��o^�0 [��p�\��ԀF��	��(��gW
0�X�'׽}׭�T�@MnjfT��g��X�+�E��ZRs���UהnP��f��P��aͺj�$e�לK��aއ3��	5��n��$j)���m���e̊���!�]��x������&����h�3$�i�Cn1�!�A؞ǳ���%�t�&0�g��y����-(����R���YZ�|MY��Mb���^\���]n�&���5*-�vJU���zr��=���C�t����H�Q�t�g�I��͕�z��8���	ѝ,_N%�o����>�[��a/���jm��%{��棠I����4,Q�(n��v�N���:���@�\�.�C�[L��tq}v �"T���׃�K����g1S:@�U/buj��0����V�.�~���=�Ƿ�,>8Q��3��T&<�j�n����@�W��V������ϸ�Ml�K�nZ*�#�0���l��l��tr�].�x�cn�-�������hC��������j�B�«f:��g�V����v�4C��b�>�3o���ab�Q��/3�'mc��mš�]�S��Ù9���:>֚�|�N�)�*�1�5��<���M�TS�8e^��XVf��K���IZl%.���f��!�
��n<3����o�+�}�DV]�NC��Dv�0Y�S�����u���7yЭ��g0��Mcv�2�� (�9���EYn�r��ⳟ`���]�'B=��aI��S���&t�����Hm;�}��	֥oL�}�1�jG�ݡ�.厷�H@M�h^ ��x7v�!O����U�H�,��4��z���0;���������p���YІ�\��;tG���;�w:p9��&n!98�:�� �&�f�;E�	�`�DZ=�פo(��H��%A�Ӓ]º��8mi��:�i3)F'@�d+��K��ot�����N�=���_-��l������,4[�*�Nv�W1ҍ
x<_d�z�M�6�.�o�fE�t����[�W[w��e��A_"�WM�8�����6^�]C�i�-�&�/�K��C�c�׺р>&b�S$b���@2Ë�ͭ��,��T-�u��2۸�y�t�=��B&J�o����e��6V���03O���S�]Ye%Ab6�����\�i"b!�O���YVtR��R�U)��8e�����M� ��{��s�m��[枒�@��+#��+ aV)������Psj��c��0���u�Z���S;�5�4f=Z0X��H�a�o7'=��Zr��ȋ�oң����Q̛����w\��W��u���!Z.�$�է�D�\/q%}��T^;{�t���-3���8:�e3��<�j�Ok�,�O��ʝM�,ݼ�]{G�k?ʽ�&���S�Ӽ�R|ZY�B��x撻�%�*�WMf�u`�[�+�S�m�a�!S0p��j�jT��%#��J]Z���:5k�s�I�_[���&�q �cն�)r�����_,��i�(���*$����b��֌UF(.HT
¦f`aY%�R(�XT+YZ�f"�P�2B�g��IX��$�X���aR���oH�*TYk "�d
�Y��C%`,$F(#�깑�]jEA��V��B*��*"�2qiE�B��V-eAETR��s3X�"�ڍ6خI[m@�9��2L�E�H�d�C%�3;Q���u����C+&I�i
�m�X�H6��#"�	����"�aUR�a[h��[rUTDU�
!m*]k" f[E��j�H��%Q��h�eAJȪ�صDd�Q�LŃTm"ʟ�u�V�y�*Z��9�f��F*�J;���5&�//oX�sgV*:u<�fu�v��]ϳw`y̰*Ę�9�Z-u����'�q�������_,~�A룑�fY��
�Vnqu�xP�@T�GG���^�Y����{_n��{M�w�Q�=�+�=�BM�����a�DL�d�9��K��#�b�ж��%U��̤<��8�I_o��ܿ��Xc��o�uQkFҞH��>���z�����|H��?��f�\�+~}cEę���J"4m)x#t.�
���iӪ�̰r�.,ܩ��JE^�)�6���YȌ�f���鼜�������Rң��4s_����@�3�
˫�y�e�M> ]N(˫S�\?S���j���8��^����f�n����y�g9/��lW�O<� _?�:1�|L����o<ђ-+Cn��ɜ��m���/U�J�Q�d閗8��Ώ;�>p�����cP����\=�|��[��S���������N��6��� �g�t��C��r![P�vbZ.8��B�,�����!:l$;��Q�r��nD#p8���X��4��i�?~��y�A�߂n���Wrq��Z���6�|r����я�$[*��=%+M��dV�ٙ��,���qI��W��DD�`��=@�<�`�G��tshl��>����N�34Ͷ�qc��E�4�sr�3���/��`;���\�d�'5��yjKJ�X��*6QS��l�A)�Րi��:�����j�(
�@�q �~��\�u�1�6��@T�k�n�c�LZu�Sŵ�s�tiu;I��w�ߞ�|M�b��5�O�P��Vڱ��h؀ �̍�F�dq֞$}=	!Ɲ�lѼ�K��L{���B�\F62D�B*&!!PM\���L�7`|�AD�PU��zI�������ҽ�Ҭ��陋����ܪ
�����G��.9fX=�@�^��P
\��xP��{E��;z��}��Pt��Sy3x�&H���1��J�t|PPTt�GZ�×���H���go�V"���6>|��%�t�N��&�}I��h{>�>!�����>����9�#%K�|�Pک�y��"N�v�+��+�CE[�X���'�l�k��Wf�*�{���S�c����k��"yP���0GyL��֪��6�%/Q���S#�﫮�f��5՞��3' ��[ʴa8&�dB|�R����IZH�7�Q�aά� R���d=��&?3ڴ�W*6�����=��J�겥Nݲ�*�M�{M��#����s�gb�ty(,u�Zj=.�o���n�Y{��u�m�sl�bt���X{��u���rf��>d9�,�塾9�p5˖�V1�@viAgb�������,ovn,����{QlF�:'��p�Uo$��k+8Dk��=v�uod��4�2��\�j�~�~׵��[��veR�`��:<�'g���ҫM.�1n�����w��K3��}`��� tE67����� �n�;�~�뷋�Z�j�^�m�bQJ*L��,dmWKϺ�.K�M��sO��(��n7�}�1��">�}D��̡k4k��|Y����/�k�]F�:y>���Լ,K�-�Q:|3�[fT�W9���k����L�N�'�T����[_9RV@�,-_rϔ�v�kʯ�R��g�,(���JE��j촴��Xx�h����@����4~rcà��������=R�#Z�)���qeU�ݽ�f4���m�,�+��!�����R����P���ֈ�z���G�(�@�q��
�y�
�Z6�ͫ=~���>DƸY�[��=$�ҝ[SV�)�~|�k���V�NK
���7�qxe�;X�&nK�t"8��f����=-�e+���!���>kve�y���fm�j
����*&�2am���7�?Ns��I���VLt&��T<&��Ո WgBd-��}��jɒMc�J��t٢��boMxv}�}/�����$��{��3�?o�a4���|�3/�[:������7r:�&˯�y�-�,
{4��'uc��jEHqTPyYp�F�p��1WP��)�]NrI�JTI�nW2Μ����u�3EĴW-�3b&Y3C�_�[Da��i7��=�
wCWxoӒ>eJ�R�ݶ����ڲ=\�}�樂��>��\.R^f#^��A�mbϾ���fxq#C��V�74pk��eW�0��N���p�����d��&tm)�ڹ���]�����d�	��d�����yVDQ�s%TGB��BU�	��aY�xi�i�G�{s��ա'o[}
m��sj�N�3���=��LL��U��l�y}<�9HE5��[uO�&u����s��h9�1����nKۤi	Ǡ~�S�w���v�X:R2<qCN1�,ϕ�朞tPRUe_�+����PX4���2�3u�u\lNg�Ҷ�{5J�WUb�nzs�zg=m
� �+ �)�<|���.1hTY�Q�K��-�5/��n�u]�Μ�:f�8)�+\�509ڂ��zŨ�,����z���[j��k;���W-A��,�a���u{�o�
5�r�:Ծ�R�n.��e:�d� q���@��)����\e=���&�X/���U�2�*��IEw!�XR%u�Ƃ�����rH�S˵,�XAl��S<@Ϳ�AZ(1�x S�v�J�srg�@l��I��髂�$ �U�F�d���1��)�!bɵ[U�V0L����%�3{�vF@�;��}k�\�υ�S��o��[�72"�R�x��7;<{�b��B"���G�Ҧpu�D���XWN̈́xJ��)����O:ej;N�we�ؚ/7��)TTˊ��T�����_�<*}��a����)��%�s���,�	�P��{c�������U ���dPf�2��r��"���|̭5c�����qg�����5`��NV��lg�����%{���Y\+�����g�o�l�!E�t�M�p���[�3=\%�x���5�����{w��]h�12luDX�R��>J6m�M�v$��8�lŭS����U�/�Ϳex.V근��U�W;�vW�*h�Kz�0��]�?y�1��θA�xo�²�� +�k��U8����ڬ]�R��1�z��e��MQ��}�8ni����+����_m$h�I����r�(�A���v!2ɛp�%��l�$	�9N�ω�zDp+U2!8m=��c���sN+��줟��a�ٛ��5/���C6B��� v���L���8ЗW!;]��.���#�!�M���t��pg3����d����8��y�<8��Ac�Sʙw^�:�����O�s�,�Ώ?����5~.�(.j���R��)�Å��T�l*����t�;��T��9��~��xh9�&y�eZ\~xt
ۇkZӉu���6oM)|1��"��t��UV������b�O�X�h���c���6�#��oR����)�Q/�o>y���ؗw�鑔���l�QJ�fBdw
�j;�=ec����-��펵1V����-��d�<;c�YU���hea��<�'~����#>q?s���؉.�	�2�F�#q� Ȑ����J�9��M���E�HNK�Bȩ����Bؑ,E}1	EN��o�$;�鯜�NE\�L�<J-�J�85]�d75�3�_!R�M��*b�.���*�������{��sv�bj��)+��
��f�̱||�(����=Sʀ�ʮ�e��H��Bz� ��]��&J��Ӳ��]�2��a���[�%Ժ��]F��ۂ��XĬ�O���J�No��`*J�����U����B����)�;:��{�|�qI��u���.b�<{Jv}wh��@��Q;/8�2�Sс�ȔԞ�]Aj�϶��h�:a�=c{���id��N�хV�>Σ�����j��[YF�\����vU�ʆ�τ��U�x?��xx@�
w%� T���.�i�ڽMwl,p�6N=C�\쉭
]��PR�Q�ڹ���Bu"q'����=���]� [a{��q!\�=�ȣY*fj;�r�Iu&,%�be��cxC�5"�
%.k0���.3�o�݁�s=8��K�~Ҳ������w�h�]Ƃ�Fq��{�rT�z�5��DXu�4��<e|�p���8�\"5���ث���'R4�=�L���Ч�'���k�9�Lt���0#��'g�_>�䲏/ػZ�eD�R�}�(G��}�␺����\~�X �F�A�VvTئ׹�,��rS^f������įL�K�u�\��I�t�m�c�_����۸�u�Ix�l��I?T)_��3%��~ :��k��%��8JԼ,K�/a�a��I���)¡�\�4֪:�'09��n��_�Ds��H�J����펿�T��+�<����c7�|r�t��}k7	5&���4{��>����@�l�(�R��ܢŔ�ڮ�D�p�/��v�{ۉ0E�ǖ��}���Wf��b��`�t!	k��s���Ԍv0
Fa��N�M�zlò�p�I�ҡ����L#(���]��1�ɏnb�}�R��%0��᧹9�ڴL�S=2�	�D�:E�D>ꄅ@w��c�3:�����q�_8l��f$d�{�.q���qύ�R���k�̋ؗ�6-��.\����Ȭ���ldA��w�����ζ��'ц�o��mf(��=0��2�ypV �j��W����xp�ʇE�/x�j�II�~'��7t�����_�΍�8��aߦ��U�qSq���@S��6>RS�bY�}P&�U���.�v�܋��nkq�qK�w������Q�l��a�x�9VxW��~	�JzJ��2�4M.|"q��V³# āb��o�8i��,7�/1�^'æ6``��q1��ĸ+�1s��/c�M'5�q�p��!8:~٤�2��Z<�p��l=�5���V�<���O����^ޤ]ڝ5O�J�.4��{��4�����<+�\�u�ْ�z�w�D1�T���ˣ�^����z���8�aX]� 3����.��K�� W��qQO+�c*h[m�g�a�.V���h�1�샵uw9����çnS��|FL�/Mʨ��m4�e�5�3-qW��U�-Zͭ�V��́XQ�c����[� �L�N��s�e)�{8�z+_�V"�'gD���E��;+:1����@N�}�*rWBo�ˌ5F`�8���)��6a�U�.��+%]���M��K��YSE#�z^�ږĚF�n����]�R*���(�}�֊3�.(9J�*��\�@������ϴ^6;n�֥��2�,�!�n���s�&r(�S�[B�rh8y!�k�T��:��u��#4z��#�ۣi�%<k�~�xR�������??	���� ��lm�k�Y�Xֲ����P���R�_p��9Rg�:
x���W0���M�����9�f���K��-��^iM��>��X��7�ѡT9̍�'����:So`�U遏���D��{�{{������3��;~;�Vhw��R5!K�V$�*~|:G;��Ge���N�L���N���sU��FxUK��˾c~�5����{�B��%�sҞ�;#as�O��D���q���"�d�{�8�Cxe���l�u<�U����(�E��j�U�E�mkW�(��g��^D_u�uGΕkm�R�T=v�>U������۷�
�7�+�n�{X���*��M8�)7Ύ�8�;$W��8%�#YKj��� �M�,��gQ[%��2ک����#{��p�7C4�O��nk�J�,��N��Ğ)%��$�j��y�&�^ލj�_$���0�r�w.����8l��C{@멹{�;��[�vu ��}���*��ߑ���u�!>̇��]h�7Wp��m΋�z�r�����Wj[��Ʋ�8�1N���� �g��/��U��މ���Y�z��tX�]2���l�Z'�����p�O��e��zV.j���o�	]�^����z��Ȇ{Qj]�	q��{/$v���5�o� �\��� �u�����jr���Σ=��f���+��S�ԼM��ٝU�u��Dt�K��R���}'��j�]`rPT:�w��#��}oj-c#xW\��]�׹p����e��xh8�	�w	<ji]:���q�u����#���w�w�Z�B�u0��f��,��u�r����[l#~nt��2�+���3�F^E��簅66u��@����ߕS
�]>O{�r&x*;�{����2!_��Z0�^;��cS����mg���u:D}8��0>�O�p�"c�ұ��~�/'���7bL��=����a��oC�y��a���)tU/��[��!�V��\� >���B�L ���@�*ꀜ�oqР[�=����Kn����H=u��Ky����t���h`E�n���`�z�[}7q�]{��� v�ء+m�R���S��y�]�W,�B�q�o#�1�������ܬ�g.���<�w�I�-�fU��l�SO2��w&��n��42G(�-�h�t��Ҏ�T��=3��y��X�C�v'4�]&�RAL��3�H��j����wQ�I�򅢶���o+21>:K����5�1�|�<t�:�I�4�:
�X.�1�D��y��(�nilB=�6�l�Jd�N9�Y�{ԠCMb�h<��J�����V�}�h��W��1B�u0����;���p�&ۧY�D{w4��z�)=�D|5��-�����:�nx��*��{�ʲ��k��¸��X;�'�]�U7`�9��-���*%�5؈1�fU��j�+�
��{��*b�*�m�v!�I]�l=ﰄ_#[x1��6�ض1m��#x�L�z*�\OHv�D�j^�0er���hި%������J��WJiЭ�Z�ќ9e�˘��<�e�V;!1��>Д������m,�݁��,4����P������DE��s+�=��]oCo�Y�Bڮ�6�u�����hK��t��P�eٝ�`��\x�|'T�H�{X�w�͢��[9r't�yC�z?Oރ�v}R o���X�$ifЅۤ�C�%X.�՗N+7T)D)͸��#�۬}�Gl�Z  $(^�:A�֢ϓӻ}Y�ژ���+	�|�vv�wsI9�	�m$�*vt[��-�gR�̭յ��s��;sf�b��1�Σ�PYE#V��{J6�v(��&�B�u�؍��ݜ}���δM1���d�Ć�����L��]wuvP��yf\�0�n^c ԭ��]��У�L�p�U#` �HX����w[�B��]7b�T����4G]�A�V�Ʊ\����̷�r��`D�,r]Z�hRT�tܡYn@;��YqY�InhM���|��g2El8mu���C*eM-Ƿ�J�WeN�ƭ��sE�>�!N(qcw��V��Ρ�x�i�y�'5Z�J���zd�V	��;o���wwG9I�i���RV(�ghȶF>�Ǵ��ڵ�����ڻV�d���s��;R��֮����:�SM��T�k�#���A�ZX��k�M��!+j]�]R�_�ʣ�򳬜��M�uv�mx��fp5jٵ�XfZ�WZUt:J	������Q�� ��,Z�����י�YQN/+i!�]����M��iggwi���]����oZLen�;�>ip��z`�0�f�&d9��]1���_]v���:�ea}�Sڴ;�����X;lTH��@�x��9�36�î���5�L֍KT�i�PR�
�S3FUd+YD�,FUh��T�u��fI��J�a���X,���J��X���	PR*�]�.e�&jE�TRVAk[
+��edFVE�aYib���)��+ZʨjUDKJ�Zҭ�Y��T
�T��UQR�U�Q��*�"�5*ZYc
�UD�#v��� TX�5�+mT����FB�:�Y2Rұ�(��F�յKB�+"�jR��n�q����Z��ʥl�ꈵ�
«��6�j�e��b R҉UU6�*��-�f���E��l�T2Uh(���u�ZU�Q�7J���,kQ����(\Z�B��jEͶ��D��b&ڰVܓ1`�f�QVӉ�o������^�ﺟ^�'��_}o��1�j+ps��^
^c2�h;�&9J�+���0����w)�S��㣥���~���������Y����	�Y�AT��'Ϭ�*����!�|��S�zÔ��S�9O���C�2��
����9H>�x�={�Vx��d���>��>������0�s����Bor�&#&#f"�2����I�
�̗���<`r�+9>��!���Ag���P��P;�������=��X�����r��~L��fz���v��rAT���e`鉫�~�NC�S��3c�O�\�v���A����<|I�:���r��*gğ��n�v�ed��~ߐ9I���hW�,�g���=J��Q�mL��/�s��
���Ø�#�~����:j=q�kD���䇢���I�x�����|��3����C���>N�$�
��y���|�^g���NӖJ��W�q8IP��2�*K�&g��_S�&��NP<J�8�����=��.���y��σ��fJ���N�=r��=C=0��O��!�J�C�8ӝL�Y�|��I��8H/G�q�I��3:��t�= -C�����p�&`~<�pϙ�=H3S�����,��������DT��c
�'ӊr�)������U��T���0z����=B��%֡�
��+�%�no��/�i���Y���8J�lʓ���p�O����1����q�F�d�<LZ�%��2W0+���*8a�?&C�)3=C�d;N��)R|��^������~��>�ɐ����NЩ�玴�=B��/~l��R|�N����^=�2�oT����㣮7���q׽��A@�\����xr�Rd/'���L�U���x��;I�Xw����I�u8��z���>�	Y�T?'	?!R~B�����;�kf"����P�"L����J>����p��P���pNU����g���t�Z��c���%OǞ�ę���XryzC�̟�����'�W�O�;����%zN���=Ӥ����}I�c�>����>���YVk�8�y��)��0'�������P����>a�2u�h��<C'hv���n�
��
���u�x�I�������VOS!�W�tɿbz�~Iu��L��+>JB~�����'^��o߽��6�qi\@�[q�^�$e5mAyoڢݑ̤���p��qꂅk*wj�4_� m	���V��%-Zv��p�Ƃ����vvQI��xk<op��oZ{���&%��$�ɕ]�Ҕ#��u���*b�{�]�;}xH/S�1�')P���{�d����c�凬+�=�xC�=L���3￸�����~���']��d���{aPY��L�	�{<��י��?w�}zN;I^�,X
sa�$�XT�yB~���;C��NӞ�<d�$�{z��?3���!��/�r�8���q���~㎹���yߜ��3?!��vE2NШqi�O3��99��R�Vq9�N�d�
��@�x��a���)�=a��s�״=I�9K�y���Y�����阊�S��jc��Ю�����A>��I����{�'�i
�	+����{N;z���$��'3P�I��s�R���=OP�0ɐ���3�|�����vr�Xx��9���;C��&}>Zz
5wK��b#�e�}��t���J����S�<I^Ӷ��1�L�C��߹��	>B����Ĝ��!��?Z����+<d�P��\��֞'��v¹�'�8g�<L������6�dg�+o4�bc���C���<���9�����!�z�d���� ��ԛ��2N�����\z��NP������@�=NKL°����X���}Ng�"�+,�Q�<�oW�Hu�w�yj��D^�s�`|Z�����3��!�\�>���9H,�x��'�P��ۄҤ�
�O~�p�Oɐ����9@�+'~���=yI�T/^�^�����>SU��U�A,ԟ�11�L�����a�t2L����p�'�g�J�5��p�2~s:�E'�W�w�>N��$��ۗ�N��	��p~d��|���qI�Rx����:H/�?u�5��|g�ٞ��,]�1sS�O�S1���>C'��qzC��ô��L�H?�ޡ�U�$������$�i�,2OP�t�{�^i
��+Ϟ��Nz�03/�Ԝ2����'��;����|]�]~�����B��J����sRǾ�|�9a�
�tqI�!�f�G�� ��<gA���hd���V3�;N�9�a�XT�p�=Ӕ����������OP�������=�ѝZ�?C{p�8�������8��B�;g�ϕ��S[�`�����ʮL++�xi\ᙀ��#�*�y���Z�W��+�9y��:�n�.׺�c�Z|D��@�[��[Ϗ1/NPެz�U���K�i�l��A��X���3�R��T�w����|�ɽ�T��n��"��P��T6�v̬?�I��'��k������~��v��z��÷��yC2xʬ��c꘎�|{� 5�\g+�]
�};?B�2}ߘ��a��X~��3�v��$�{�H*Β_Ǟ��:C�����7|C'(~IRt'��d��'�'�T��6���
��z��r�`T�1�9>�rL�eN������F�O�6#��˙�%��ǆp�y��`"y�?3����������3=a�v}���;����Uǿ~��~C u<���!��/#@��u]u�t���nS��f
��]�/dv�_���_����*��7��3��ឲ^o�z?S�N-��:�N�%J��^�8:T����w	?'��~a\�������y߿��'I�!v��U!Z*���o;���A\���V��������Jʇ	��Y7ԕ���N,��:L�?�2OP���p������a^�����!�J���w��J�+%y���8����X��G�1�L@#�U�eh�d�����/yu���P�����8�'	�d��~��W���C0�*�r�'o�,� �@�0��2�Y�:�8g�ԙ�_�p�U�!���>Rr�H/����������T�u;7�>�*��;�R�7�H��>�L�Y�;�	;B�l�y�V��+Ͽ~�L���*~���q�8d�8�3�K�'�	����M8���9H/�tj�x�����s�&>����鈯yG��#��=���v�w�����:C����������?}C>����y��|��W��px��OP�~���NU����2�^/������;~xN�h��T��4���AT���}�>�޻����z��o�Ԟ'I�z����x�>9�O��t�Y�~->gz���:��T�2��v��{�8k
��~��d�ԩ?�&|d�>N�3+%W�
�=C��{�����S����\��}����t�	*J�&|d������/�������z��;�<f{`T8g'��礞����>�)=yI��2~��VO�Xq>�z�)��oޮ�Ɉ���1���y]�A��{P��R*Iw$�OPL,��^V'l`ԭ�z�H�1Bmiy��j)\��x)U��bs�t���I(����B;�pެ<#�Η6���ܦd�.o��Y�����bu=���!�r5�:���>���h����+�;�|��H��v�3�b�H*�ӎ�q�'(du3�|ɼ��&��p�'�gO_�8I�<a�מ����&g����&}`T��z���M�8a�9FO�?|����ସ]|�=��~�_/���þ~� �"��y�<s9H/iԴ���>C3����8H,�'=S���H/�����̬��egIݡ�=J��9����xɒ|�}��9����:���{�����s^?}�|d38d�����:C�����_w��8d������R
�ϖ'��f�\Y�XP�7V2�H,�ϸ<g(v���u݆T�2��v�Zp�_XTo�y����{��������sߟ������{��9N�Y2O���3
«���<W�o�r������~����:�l��X��l�^��Z�/q%60���.��"�g�ڹ�~m���I_o��ܺ+�`8nc�z�p�@T�K%�o�w��8ښ��s«�O��߲�AeE��fE5C���3�[���>:��ӣ�F��?���:���S�u�f�J��,u]Y�,���=.
K��j�c�f��{�C^��[���.�����`�u|��3�xZ�7��C�E��j�/:C볚U�s�%�-�_5�f+���#ݴ��K5�<����:1�M(���l����g�������S�e�~c>��*�:�xtK��'�"��\O#|�uv`/�e6�3�v*�!ӛ����A��l\� ��&����h� ��m�{0��zr=7� �jn�(6����A�Cj�'�\�&��	���ʼ�m�v�<ڎ�;��l�Yp�p��LTZa�1�9�[OuwT���]��[�"���(��t���&�?���7"9��G|�9:�!�5Jzy�Q�dII���ڙkf5\(�'h�+K}�E*P\uW�qF�O@=�6�:o�骮g:v}V�Zh?&�:�g��2�%py��S�IxMg���N$eco>ySCg`���y�%
A��Bn�}���ل���+ �/>����!O�>O�jb�z�jKj�\����Q�'*7]��L≝vql9#P�����蔪���ѿ@e��#kiؽQ�˷Ճ�a�u�l�'�9���u�٪��Hl�'n�Ȗ#�B5s+�����vj�Ó�Lp��ǅ����f�r!T6,<��S���y�S*BHRf4@R���(C����y˱���5�!!�4��b���6�X��`l��@'�')*�6;/����ֱ�G+f4$؅��[n{b$)ۂo(B­���>l*��6� ^�k��%�z�v�|�y��}��lfW�������88X!Y���<'|�����8\>}:�j��6⤏N�\+�����v�\�W-�~���+d�>�jƋZ7Le6 �Hc�1e<oxY¤��-k=�n��l9�3���^B��Fv)|;d�"�%�B��R�<9<���cB��6媒خ��<CJۍ�3Y��|y>ϗ� �X����wNE��:���t��{�,5 V�.\�5n'��+��I�;�3�*BY�/眎�9)c��~��Եb�x��2�p��¬��[�೯@�r��ʴa�������E��+~���gZ4���+��+�>X`<�s�J�U�Q;Ǟ03B�`��O�?zl�0V�j6lE��_�@5�.�G�w|���\��b���i�/�k��4�R.��#�w�=Y�3��������5�^��;�c�Y0؆�����x2g�K��*=��?Oy{�ܧ(�#�5m��f�r�B
�Ю�zkgWOs�����:����.Ѯ����"�r\�T��1��.��]kE�v!�J{>��eNč�QتUՁ�t��w=&U������p��$��̌pU,�;;mOwD;�٨X�!�h��ڲ��8����8���ޚsb㎥�M�ޡ͈�6�"A�=�n��g^��:�\�����!���u}}w�a�W�j�e��h)Z[����b-�<K�����D���)����]7��%f�Έ3W/�5.�c�����i3�2c�ږ=}�u�O@�q=�9�-v �u�k[54f$�+õty36l��RIZ�9X���{m����N'\}�rC+dᶮ*\@�\#&:N�ͤ�$�(��4�4p��Yg���� J�3/�j���L�'����QP��Yȅ9;�ttD+�ٗ��c��$����D6Kˬ{*�U�	<���C��� g��?���x�T�] ��xf]a|0Q�����fLÙ��lu��mN�9v6d�_Wxi/a��me��yb.�
�����Gq�s���54�j��.v�t�����M�	@�@/��4���Po���u���N�*G8d]�-���&�l�qu�k�UA����O3!o�q�<+Cĸm�+�'���h˄a�Fˌ�|��dpr�V�����b�n��8}i�֌!�*�6�]`�Ӗ�g�� �.z.Zb���ٿ���2rȊXoH�
��ȫB��Xa���ĵ�2f{�
a��sTN�&�2�}3�7
��}��	��zx�����,$���G.z�������Ʈ�H�/~J�ƵU�2�}���A{���{V9�M�&::�3��&�U���'A�2ھ��|�*yt�8d��_`�p9D9�m��2�D���gQ���eoB���(F;.6�ey�=KA�3� ��0.�Ug�2cyj>
�r<2K�D>�W����5H&"�)=�f�vD��n�補���[
8�\�􆋸3ڱ�Og�o�ȭ�����ܧ��K<���ǰ�9�r2X�wxwf��_/FF��5����)�C�̊� ���3� �^	��G��&��U^�a�D{���m����S�3�Ԧ.z��OU��D�)2T(P�3â� �^��[T&ptķJZ���R�5��$#\lAb�zj�N��`�t��}�����KP�p s�F�x�ѰC���ro?�u�	g�{fM��c��@�@��5������90��Z�8=f|Oi��=����Q.�=R�)�Po2~� �3%��v*n#1��S+���j*Ѿ��!�t=��P�x��h��y.�.t�銒���s�{�
�4��]�?�y�A�k�-��O\fؓ����'�YX�6R�&���٨�f���^�̴6�O�z�+�yyj˪K�`ߦ?��o[������u}�2������P�R��ߑ�����>̆�j�N�f�"�+f�YPb�[�Ӯ��3o;�ݫd�x��c�zi�¹Ί��I��������v���_�LVR��#%?����FJs���h(E-[ώΆ���;T.����$5��1q�3��=����b���79ح�o�����W?﫼�#�o��v
3��BΏ ��V�W����d��l�ׅ�T�<��d�a��Ɔ�����*���G��5�^Fg�֋t����,+.�^�\V�~��3������0���e]_��nf���^���l,��>�o��\� ��ݮ�h.���?o��'<�v������yY������f���nER�e����cmu�|��x^�L���q�bQJ�7#��F�P���Nc�\CT��>��D��2���䠍}��&��f��9�9�.3B�ڢ>��G1{f�N�Bх������|�%�Ұ�j��wwm��3�V����?����KGO{��h>��V�É�#���i��ig�������:c�E6Y�l�� �O����՛8S�X,O�k>�5� D��Kz�(��_;�=x��9��|g�E@
%,��؋��3]����6'.a�x�֥Zq���FȗXo��o�H�}Bz\�;	۬��H�iP��=�	G���c�E����8��躇[e�����m]�Z�G��� ��vQ<�M�;�j$Φ��N�ݝ{��]���7u���T,�&nJ뿐r֊̫�0��p2t��:�+��f˛O�����Ԃ�v�]�aV���Sg��DC�޲q�' �ߢk�5�Kb��ľ���Ι����ԩ�N��&b��9�8LXv\�v�pn~w��݉��2�qL_�	�s��|�(�ݮ�@�ʀ��Q��.8vN���Z��=��]�#���1>�G���ؐ�\`B(ۼ�,|ȵt�Y�%TL�����" /Y�O�&��g�֌)Wm۫�#�Ug��SAOBFD�������k/J˚�����O� YfR;�%R���Wf�Z�ay倧J �[}�7��gn��{q�s��2�XG���4A;�8�/t����}*��d�� K�r�=��uz�� *.@O��p�+�Q��LHo ��٠8?	�{��rܟd8����6��Ox�uG���z������)@���?K��0V��w�H\k���уY�׵7���#c�D���I̢��¶��ߑO�X+:a\��yt��V�e,�*�3��<��w_���~b�����S~}xpD����w������!�l���G����������p�)��5l������+> ep���sG�ڂ�[K�ڻ4`��	�R�E)�HN�3
B�����@C�P�d|�ԼJ�x��cB��AKȹ*V��z{:V!�cܾܦ�wR]��Y&7W[��1�v\`�Cf�8�p���86V:�.5�h��� \Mem�L���
&г^s��kZt.	ܠ��Y�̧uyZ� ���|(<7��1֫��_Gc�`9O늠K�.����Y�e#;��ɲј&B�wi����)���N��w���t�S��U�x�*�9��RN���c��-;xy���%�%���$+���X<��S�a�q�i�/�wK#x���c.'�*��5� �v�/����F�).��r/�X��_*%�O4��0��$�ۡas��5m�G%��Kj���.Q���掉��cɛ#��#�D��3����sĕ��K[�.	�*뻃�6�S����J��vU���"�9�̮�wR6[���Eq�m���Fї����<��Ɯ� �N�z�m
���w�	� n��d�75LLZM殠0A����@�s8W��-p>|�[k)�bVJްa����em$�uqq��d30��h5�ud�uVި���'�+A]@f2�с���c;�c�c*���]�Z�
:*�eqJ��V�]���}���^߭��������oojw�o랫1 P|��N�ء����eb���x��m@y1P09�D,PT�ҭ ��9O����*�N�7�k���^x;R�^ur���N�t� ��o��,���\��Z)ɣ�]���3�
ܩۮ�b_gP��Yګ�w�@�<b��C���t=`����w�be�Z5�K����F�2��y�k0�
�S�YS�/��lsc��{]�k�X���H<Y�OMB��ɾ��A�z�.�B�CgK܎��+1�4�]\-P�-{��S������W�X���R�[,��Q��Ķ�q�G`��1��ˢ�A��奞��cW������L�`��\#�A�WF�H]귚_�ug�` `�u�ئ�w�Js�R�����Q��J�*gQ���V�}ɒT�"(�F�̚PWtU���(�F��]��b�]��z�w{����n�w��Z�9�t���m�����P�A80����)s1oKַ���Zgȹ�(�T+��j�n)U�o`��[�� �k3��(`l�]�R���3u�. ��ɢ(M�ܩYң���r¹�o"�.a2�=�9B4wӸ���T��F�N�}�~�`7�GfL��-$��n��}ݖ���]�ND��.Tv���[�hS��{���� 6�i��.cS.�S�Y:�uk�7���W�۫<�nZ��0��`�c�~��~��?�<�2���e�E
��
¡QEPD-�\������56�Ae��
����"��Q�b��+�����YVҥJ�c�.���ETb ���lUUP�-�����ڻV�-j*䬒�0�5���D��h0VJk�����E��h����-e�*�.h��m������mh*�U`֍j+iAD[f-��5��h�A��r���kTJ�ڸmU���`)3*��j���jcR��R�(V��;[iU��X��µ&J��kmJ�M��ڕ6�P�E�Uu�"�����X�
�Sbk-�05F��6��2V��GZ*,EDTm�2Xԡ\�Q]IWP���p�J��3ZjU��cMr�]�V%Ũ(��%ԭB"j��&�#���۱߬n��
�7�(8�u04�\ �䷱�����Q��c P�#r5�:�{}���T"�s D������}����*�S�O�����j�"���5�|+�u%��5[�	Vk���o�~O�����V�Ԅ��<��Sٲe�˭\�Y�&vFɨ��T���"9�W�$E%d�����e��S�C0�����2�od=a�)�qJ{��l#�G^-g�@Gr�q��?]܃��N� y��]]���Av�\4.0>���1�=���vn����]&J4�)��}-�Y���1�u��5#"&��I�ĖE��1�;�}���_����x�v��n>ysՆ�1�*U��ȿ�*��٬�g۞�zyk�TyX�K��i��Ld8����Ԛ	i�&ؒ6#_��q�B��w�G��Q���M'��U|��.��Kۮ�,�{���7����9��#1�D0;�����z	>�yJ:�~�6��B�u�i�&�AV�/H��q����r5���zW/H� �x#����˔T�yj�����~]��V��|���8B����-�BWt�����̅�G]h����ES��o�~~�lzܣ����;��/r������]g>��&�X�!�MZo*��.���И� �>�n^�7L�`�ZNw-��U�4{d;9�9�֖�Ѽ��7#�GV.ޮ�  ƅ�zq�ܲ��/w25�-�ӥe�Y΍�y�u/��Y9;Uz/Q�DG�DC�w�V�n�M�7�eh��@�<":��{��xP@�s<y���@
K�����oGg�f���zHz���[�r�����vo��-���p�5\F�l*��ZZ{^g0z\���|ޥ۱Ln�������g"�NV'g��үy��hc�m�2�<!V���$gp����OqIҬ!d$P�����&P�>4��LM9���QnQ7������x6]��طn{\�Į��oZ�#ùJO�+<�����5�4��9=��	(s�����f�?r��XHGS�;-,�;��c��S96�;��|�9�O�[o�.�_����v_L�3�_X��*O���z����L)���Ļv�u�n�3����b�x�������^Hx�\��_Z(?%-ϣB�p4Jx؇��6zcf,
�Y��̙Tޒ1v�ՠ��б�F����ѡT9�M���
y�~�淍V�.��=ǘx���X���y�{NO�*�:����8=f�j��ʾ���l>��a��wAw�I�1M��v;�co! ����8�2��U�	������ӹ��1�p�H��I���ٶ�-�����\8�c��7��lU��D�Z��]��Z��on����L��M̽1�؝u��^����}�9�OR�O8����q��ψZ���fU�[7����!��@v�iv��O���s���;떻18��9� �?�bܦj�A���B.fOB{�7������|��}D��g�o/����=O���ZO<T���Ek�9�����o����0�9r9�̕7����/wK��ѡZ=�c�o�:���U���VpL��ϳ�"5��|��'ِ�eK\5�'m���\m�V;1#at�i���ҍ]�TV����)��)�6��Vr!�9s:������<��p2�&���V��o�n�:�}�������� x�������士����Ǣ���c]_�|C�����,�)��o� �]u<�UC�Օ�I:g��8�����~&�2���u��F�i9�q.qJgG�oT���Z�s��3-"�U��A�Q%���P����=htD��=���
vo^�p;�3S�R3Ee��S�
�[/��~����t����5�]�phz����u7��ꍶ�MԘ��}���9nu��;r�������f�޻�Z�x��hϚMӾ_�S��ūͭ/=���51�U�G{$��ޛ��&H�q�P�2��ol}m�(��.�l�"/u��;���(�M�gڤ�b�����7/O_ۄs�Bxzϻ�G�}}����9��kr'B���u�3
�������2�;��/}�>y!���8`��&l>U��y�zc��8?�/��ႴU�R�]@f��D֌%��Z���}5?	Ѩg]_&ҮB4�� �'o���:���OÝ�\�G��:%*�B6 kF�^M?�ȥ�9�J\npWl9�ݤ5�R&��@��Vn�[b��TLBB����7�0�K��3���]��������J.u�}�ޘ �����E֮+W��}6y�m����]AY���;����}ȵ��X�*��3��7j�k�^�h�m"��&�^�{M]�b�y�f/	SG��X�
v�Ձ�uu�|ȶx�C�9��O����ʹK��^G��#Z0�]�n�s����$:��T�pu�YK֑}䫋#��'^�'E�8�ܲhF'_MB6$K��	>�8��++�k�;O����>w�'�pSI�Rfd���p��!9�gj�0Cβ�y����6������΅���mC{u�����,Ly��B�7��t�sk����s�k-۹1�ӗC�`��.�׊]��o�ܫ�F���yͽ��*ȫ���Eg
L�)�P�)����iE��]oa|��k����IGjj��I���yL9ǫ�O�"�f9r�Wy�TIZ���}��}���Rq�E:����)����6z��<.�N�w���.�m�bWlF�:'���P/�Ϩ����;����y,�l5�wn+�>
9S��%�f0�ކ��7�xr+lò ��,@��$z�b�n�(��L^���`��N�J��ʥg!ƝV%�t���gplmуb5�C��2W����Ө��|�wXC�$u*��jg1��W�U��q*Cr��?<�ו��S�T��:�k�V��Dn'�L}��kB�:��� g�֍u��F��Q���qg'n�g�n��3��y��5u��.�s����U�k��=g�8k8�BIF[}��T���:�3m��(;�9��3bvJyp�ۮ=u@����I��@fZ[=��CA#d3\��������N��L�!��}9���:��[��eTЍR�.y�X3�G��T�:�MA\6̼]�ۜ]v���Q�q:����m㣫��#�α��je�+T&o� ��EAw�@�Uvp::#&�}��+u�_^� hu=�z�D��5�˚˨��XfQ�l�d�Cq���pl-���b�zڌl��}vl�ȓ�m[*�}[�>���RQoJ�0x/yw�n�#�s�-+j��������x9��e_+V�T�cq���۽p��?�}�}D{fw7�S�iU9�_��!\|��.��ΒGi����x�_>�H?��xf_�p�b�Ro�W`I�m�Nķ;�oKvb��I��Ȗ�MNL��b��-�22�����孏��:n�<�,�J�ٯ�ޑX�X���_��x:�������a�{�8h,�7��k��ʩw��Β��ɶFA���1zWv��TX��Q4��,�6�FG��)�@^��7huZMg���x�����vF�_VpR�VA�;n�+� &�q�8|"��O(��<���Kk�����-�~*��/f�!~X8�u]�C5pv6�k�F頋Ɗ��ƫ��gW���ٕG���Q[�8G}�3�/�
a�\���ZU���}3�5�,�5��}E��0����4+�q�5]�e��Ƥt����*��x\J��ʿz�31��<�}�����l�t�9��'���<6�{'�̪��+Z�#�yD���twmn"EB�EԲ�ˊ���6�
�ϲ8)z3]$ �sӊ��]�̺\.��>��Q�	�;}�EAs3�3SI6W0����˄vmj�N)>B��ݭ�:'�;{b�SǘdD�@#������P�ך{M3�o�֌9|��u�e�k��mÂK�m�oE�u���Ԡ��{�`]���U�\�"���6-��}�G��X渫t��V�J��_\EX��<.g!�@T鱿�S�6S-��"�%c���~�վes��^
����h*��EK
Zb4)65e<HF�
�ݝWXLS��>��e"�)���L<CmPS�B�>H`�!͘�rq�,��r��P��`��^�3Z6Q�9z�-�W#��h��r|�V��|M1�Ё�jG]q/?V@;Ԩ_{m���$.Kz8z���Pzg��t�f] !���f�au<[�J�hڱ摷��/��i��U� �vh�3�s�'מ6{�
����^��"(
�ɕ�D�AjжXܶ3�6s�6z���}C�pv:c$�Ba_ȼ�ڹ������2�!v���v��U��x��z�g�`t᮪[��W��k�����LK��E�����[� ���ң��aƬ�(���i�\=]�u��\j�"�6�L�����;׻�^�sX��U���0��O-�*N���F�[V�� 0����ɗ�V/=v�I�ꎱQ���w�9���Z܃��:	ԧt�*q���jRN}�����T��۪�79f��1��ɑ�vD���=�:}6���w��w�^�]ͦ��ɔ�j��s$�ח],)X���{ ��)B���T�0l�״�By=V���:ct�N������興^ћ|��� ����3i�ᘞ
��t?�\��1^6Cܷ~7�+��6Ջ�Fm-x���v��k�X]�W��������]l��nߘϥy-�C�	�l�*u�nM��[�k��G>��i�D�2&�F_�^&�+s��;:�Q�*I���kLonn����J���u촸����qw���Z1�L$:1�t®��Ĝ*vej�u��Ѫ��F�����\�.5�&�+��`W6��M�#"-��ʉ�wj�\�X��dgԫX���1�����3Ǣ�<��av�����jE_)�+�G�}ҹlԺIg�'���'E|^,�$k�=�P��u��M#(E��0#z�y�d����n8�2'���F�7֤K�''��*n!;u��e��!!z�\�a<��ͼԒ�ٜ4�?�(wl��j�2+�Ca@y}!my��zF����Z4�4�|���צ���~�Vn�T(K�%�2cA/�w�c@Z/☿�7p:�YS&�lM �����M�[����-��}�Lst�Z�J�9���a����ݺ�\]C�;0Jý[]٬���eAu�-��2��}|�\;����Umj��hY�R�o_nE����v�@7�����oL���DJ`.yƓ�L��8�����G�#����W�@�Z�5�7���=~�.Ә��JïÛ~l���A>���/#�n���M�l�uc�Eሱ�������p8(��ӽK�U�C%�C�
U4 ��#?`,�Gt䥏�:���KU�!�CN�{����ՙS3�)rRW�J�:c�,O�����%%�r,u�E}�@�ޚ�#��ͻ^��ީ��:�=�c�й�[ʷ	����t:bCx��a��1���݃�i�/$�Pt�V��>� �vy�Z�}����ۥQ����Y��6��R�"6��p��Q;=>���E�_
י�S��r�a����:���<l������ϲ�d�L.)�H�T�xp��W�����ct�Å�>����1Od�����-���TM��G{"��}tkB�W��K���i
Ѭx��I��[�[ls<�ob���8e���bī�-�R���"�:���c�9�*9�W�'�n�".���==���6��BL\t�n^v�����N����s"�*Cb������]Y��	<̢ݪ��޶�����(��9Q����jV�W��ء���_ہt�q�F�L"�Ű.<��:|o�X�-Ч�o�+ Z�+�y��.K�����}���G���k�輥3��9#�|�����A��}4�v��I�חs�h �D�D=�UԞh�fZ+n�H���Np2."lu�B�>�	�#a���CMl��X���5t���3c^�U���MYHg��X�e�*��A�0��̍���ITVW[c :��3|�^[�J�ື��Y�ٹѡ���'�q��*�8��Ƽ ���j
�o�� �o�ڽj�Y�f��%��rS����t���Ó�$V_݁��EI�T�3��0�b%��j�y����sY�t@U/�(!�{�}S}��T���v�y��5X�ǃ�7��2�ԋ�`�\�p��[��j5��rٵɱ�A�W�#��;mK�3#�s��8��m);b�G���r�|�GL
ڄ��[��~J"2v���G]h��gY��ؔ�].�J�9褿�b5�O��k)�p��^����S�.��3�P�5O-ޞ���Q�<�Fr]�G�-n!��(۫��[�-�He�f�ލBuуԦN#����ޏ�wO�"�9m4̣����*�A��,����ܮ��K�Ji�Z�R�KcVM�E����t�����9\	��$&7ol�(�Y�tMh�֝d�`�jU�3�����kq]`��$tN����+r�h�s�������{�6�Ӵ�g]�ňZ
D�/xS.�7�����=y|cx)��$8@l%Gu],�z�:�ۻf���t���A�����a�=���VEH��>��/m�$��ʐp�/�X��q�{������#�vnAz͇��=w-y�5��B�uH;*�r��Ge`#�o`����n\746�٧���R�_b\5��J���a�&�.�e�U��9l ��	��ݙ�iv�]�ٻ8-xEo�x�����Sjp�w��(
YȚ:=�DMSks���D�'@�ܺ�K8+qj$��������p��q�s.$��g
"`���C,f�h��Z�)�J�V6C�vt,��/Nr�w?��`�Ư�T�9u��R`��⳻����w��V9��1���6�$z�g̜5k�r
���ё�j�e�,{:�5|EB}��S�ν�af��b<8��U���:G�d̾%\�BĆC�\s�HUG8L�g�[
3���� Æ]�ͩz�����仅$C�`���̪�Vz��w��İ��1��ӄR��Y���T��|kGga��طo��4
��V���,
�[�M�����^�ǯ�W,���.�i�����Z���j�>̱�.�f�@�>6��Yt�SRfF 1�fD%IM�g��=#���[	���X=����xrWiW���ZM���Ü�5��H[��M�<��wk���Öt��O+Մ6f��v�w2n��q�:,m7�H�����D�Ƶ���ʷ3b�W5X�+��}�"��/�{�n�W^�;;W�#���7JR���䳝���M3E�˜�c������w�bg�:ܨ�v&��Xr�4��
ٝs����ov�@VF�.�e�WX&i��No>yx��.�r�N����d�����a	Q��YJ�y�j����.�si\�t�W�)�������%�}I9�<��F��$���G�O&�,(nE��8�R����G)mLzo2�5Rp��K���5�_-� nl;�m��i��F�YG���W-�ś�c>?rI�x�P�@5��S�rؠ1�o�Q<r����wu��v>�i:�U��'-U�8K���'c9f�j�ܽ�����>�u�o��}�1��(ۮ7�6�Hn�-^U�_Xǁ��ؾ�����ts��0��.%�01�;*�|����dΩ�����J�Gx�8$]�2`͗������3@|�PX��mulY*
kUZ��ݳZ*���r�	l+b���j,�n������A+6
��E�]��bł���eb"�u�J�*���hkDKlb��`��\�(�QQV��cb�l�����AR+K��Rڲ��V��U3��V�R�)j�f�\�QUKE���h����A�]�Z��V�Z�F:̘EFkm��Y�EAU�6��.J0EV*�(���u+b1E�X
�0�b�)n�V�6����7\A��E �(2�#AB�KJ���Ԣ����֕�����h(,laUJ�Gl���r��a���-�Q*�[R�Q�u�fE�fJ�+\��V,\�V��[L��Tr���Z�Z�Z�\�T�f�\�9*+��1�kUF�ku2��šm�q�E"�hƉij�VD�Ԩ��(1lT��*�f��������~�;L7|���"nm����s�z��C���?q9\�p���T�M����Q}����#���u7�m�) �	�FA��b� l����vH�^�U�B�𺴫�� /�?I�D���%�ozO\�թ���EŔ���3�9HFn�$��v�T&/�6���/kf�}d���]h8꯺�j���K�F���Żs��-϶r�fN�D	R�Y>��Ӳ�������p� �# �c����8җ�~�M�;�ӗ6�;�@;u1�j��
z��d龗}���,��^��>S�T��Ӳ�T��9am��zaOp�ԦfEm��I�����(��ܐ��0�tL�ۺ��İ��B�p5ORRE$A�O�k D����.Lx�F����v�[��D����!Q�`�Ƽ�k�i�x�渪ӖZr���Z��भ��3C���"+�YJ��� ��h�/D�#Z�8�BtW�}�T��B���-����R�r����;!����S+��uai{Y
�Yݽ.IԶ�{����j��[f���Wınq3x��n�c��Q�2o��$:��E
��Ү瓾�f��)q�@��aPkgA�����U��3Mtk�-�@�m�}�U`M-S-уn�f���6I���	��WM��UVg]!�<]���uJBJ���H���t����*"�e�4n��Ygl4���G�W ���67����]��Է�⼙��s�Q���>�>����n-��¾�W�b^:���v2 �ٯ������b���C���t�X8��s�:��>ge	mQ��C�ي�<c6�W��U�m)�Uq�K�Kw~�F�1�ik![6˪���KҲ2�=7pr!��C>�0���4�����Ϊ+S�^Z����s�O���v�?.yݒ�z�d1U*���,e��q
�S�#�YUX��?�a��e.��;m� =��~}��wS�r޻ߦQ�w8亷]5�/��Z�0�6��N�ߍ�։���;p�ԉ=SCi;Q_�9�09=���d7������_P#]���3��a��=~���^g;�>p��uP8��}5B3K���
{B���OH�-a��;�����su��*� p�W�w�yE�� 8|ȧ�i3
�T%��Sa!lo+����j�K���Z�q�j��ʴ��X��:K�g4���q-y���XU�'��=��ˉ��g���|��>�p���\��jD`-��xOvl�+k��j�ނ%����$P��u��E˧0�ґ!�;2��CN��L03OR�n�NK�ͭ"8V_&;�
���e*��Bh�� ��(�t	���x���=��,�`�N�-��U�g��G�R�襓�6�Y��G�DD}�s���&�S}]5?�m��ѦDΧo!��6����v��AuxQ4�=<�77�e�ާ>��ۆn1dqI�#[�@C�''��*o���B��"�q�:�CL�&�����u\�4�w�4;�k�5�Y��ᐺ!���<UR��P����+%q��o�c�]m

\��)Wh݉	���e1_ɛ�9� �[�����f�#h��d�Y uSʀ�ʮ�s�
sȎf�����o*��n�2k�g��ʻB�{�6���DѬ�q��#"�ؗ&t�t
`��&�U���/E�8X!fe�^�¼/&$�/!��� �&�F��hE�_{�H=�,�)Ӈ�Ϣ�5�g��d��ϰ^*<��C\^����4�PɅ;�r媪BX��P���r�_o*fER#�`��-Y˨�:�_Ra`-_8i���Vd���S�W3M,tă��E���fk*���ׄW/3��5�'ð�V�\��J��^e՚����u���)�������382'J:k^�-g}�Ŧgu��u7�u�ga�+����B�M�+�<���wӷ"�b�:t=J���!�g���JW�y�Jr�}D>c����}v���&�u���^J��t�nB�Iu�{������z<ܲ���ôGM��;�(d�#G��vzZY�Y�
���u/z�C�D̋Ƭ��H�]�Yb��dB"�%���l�PVakT'�ח�W�M�ϩf;��Z�~��e�rq��
����Ϸ�
G��_�F�;ϯ�Y(}\���W<�;��������8�.�US�ߘ��|���MLիkjPr�'��Ż�L����;�S�9ы�醟<�X�Wv>��:����5���[CT(6磦k�+f�os�F�%%�aF�qhmAq�D��P�WJ泊d�G�\�u0�|MT��<�S�H��e��gD�m#x������;M������)e*��\.����=���,�@���p�ȵه�ǟ>�Ϗ+�����{*�"��7u[�K���-���oېo�gVj*+N�Z
�)���Z��򬊄�*`��}�-t��k��7=s�O}#��@b|�=�����0y1� ��9{��]S������X���#R8�H[�P]wE��:��V��˻#4j\�e��ґSX�M$.�&i�����J����_k�+I�2��1�K]ղ���1�q���U��t���RÇ/�}��}Cpƺd�p�=�Ec�W�-�&�|y�xچ�:�Fd5�5p�p�b6���;_�Z㓽/����w�ٲt��:�Uޏ�����R���h�|�%!o�ϖɽ�b���f����⎦�'Zc&���q�y9Wj+Q�q�����=����zo�u��5�ݪ�B��LU��("� WC��ݒ�{�`�mT�'G3��Qŕ�^�5��U�x�����E����Nq±t'����M&�U��߲y��"�>����s���m�җd>l��چ��|�r6r�¥�Zh��"]�d�/�j9<�0r��&��̈́Kz�u�-ֹ_�y�i?E��΃����%mboc+��L�-{'w;ovGzs-9+/�V*�'�A)BQ���'�"8�n'�Ô6�����SiT=9������(�M�|��v���4��J9[�]�2���{�;G��ڨ���Ht�a�n���PwCZn�et�{s�h홏9$�y�W(�Q��"˼ɱ�ڳ�^ 8���g`��v��Ƴ���N�0�����>�9"�en���A���p�+�e�Ʉ�R�F�$��(�����w�	�ry��8g�t�]���J}9�<��h�F�`�&�o8(�SW��o4���]�r��Iuq+�����]��}��Y�?E�~'/[�E��-��ޗ�����.�j����*�7	�pZ��ǒ*���Q�7.�v��&�֊�Z�9eA6�Ŷ����潤V�
N�o)��4^}S�4;q�x�rk�w���U��׻9�a�Z7iP���+����o���f�ٓLF�NtR�>K�`�^QyW��4c^��֤�C+	�N�k�N�+F�r��o,�|c��e�k��\�xH)��_��M�WS|�Z��v0���v��������+Fv�x�`����uoO}��ǵK�y�Mw^��6�t���K�?.�:DRpT
�]�z�OL�� ���%�B�)�!F�N�j�^�{�������,F���Cw���d롣�!b�ww2�,Tn��j���+nQ�7H���gb�t��˜� tK����]��e��D+�+����������:M�LJ3U�䫮5�R�ǿb�7��w%xJ���D\=�c�C6���ចM�^�:[G�~�#�B�G��	oa�*I\��X�IqB��׸��~�P��o�U�C��riθGjӨ�M��Q�N���]w�q��{�{P-aȳl�@�S��Б��5���(��v-l]���v�}Ƣ������[�g'm�&�`��$1[j�Y�MaIT�����y��LE�E�L�-���kjt�tjR�`��Σ���G�+����'÷oS�(����8������ӱ��v��cB
9���G^�Ҟ�p[e���8��R(=��ϡ�zUf��D�Nzef�׎DW`��q(��0�P���RY����-C�.c"�`�_�߆�Ҕڣ�${��A^T1I@�I�m4	�wC(��{��Ե;�)z���-��/C��m�^���	��;a���il$we��V�Y�q�gt��Vr��ޫ��,ժN�.Fk��kd�f2q�p�;��B�����&��fI�<=�j,�>B]6a�Z�������s6r�[�u�'^8�}qˤn=��T_ϧiz<�^pǋrwƙj�l�)����b�|{��{�����YQmN��y������SR^q���VD{</͙���1�F�pyE}k;c��p�1#����$^>,o� ��������=�m��T*�Uedd�Pa\�� ]8�_��������'m�m��c�_���ZDv��	N[ū&��&wf俳��{��g��o�÷��V@ꀷ��z*Y���H����B(��F�ڥ�8'���d&��j����y���B�:��0��8�*���=L�kic�v��Ax�L�|�w�xu��o��'�L��l���{��}���1����߷\�R��Ȅ]ܞEת�����&�}���;��ZuA�|t2%�`߸�m5u��C����k��Rν\\vgS���Y�6AˍN�fZz:�w,�Ք�_j�����m9L��U�t����n��.���(���_}�W��F׭;8�}nյ��DL%_L%Q�}~{��]���6��g\���qM�7�Fy��}��s�	T<��؄�LFB׋��̱#{F,dX��Z�l�X����w����"����]Qn��.ԟ�]�3�gTY3ˣf�Sl>)ݘ֡�u�_C�-���5��E�5�&���vk��+m*�֊�Z����Ϗ0�P��'���˩s|\V[n�������n��u�E}��ŐF���<����VLdS���F���f\G�>������{]�����?q��_f��&�>m:�dÈ��r]��;��@۫zon�Ƿ���j�ޭ�aƽ5���S>S���vt�>g�(�>"1���5�s*$���U��I�i��+��<=���2M}���V+���_ZXv����c��2z!��o��R���Ŗ����F��;�(+��z&8âj<�Z�`����_K�*�Lܙ�7���{���Q*���ׅ��m�I��\y�YZv�L��j��\$�]S��밋���W+��C�aW�1r�}�Cv�[孩㾈̾���Fs�j�J]�	��s��˄�q����M�����1/ys���n���+xی�z	���N�[}�!]LUN������Px�����+�)E����6�d6]�`Ԯw5s�{�ΊeqSvq׋[��U
�D�;-��h��J���z���
�;��G��<_�=򳐝��/],�a*����,��.��XH������J��ƹ�;��mJN�<�Qң�0�����s�q�;�wK/�=�n�9�)�M���^8�·�*-T�A��pw�|Z�[���� ��"�mƧ�
��,;E�{��*0R�VUP��ZZt�\R�6\�ܨ�Gn1ɨ���k���W��VSi5��d����Ԯ3�S&�)�܀�_�/�/0�cH:���v����5���lJ�;��u��U҉�;k���u�cgܽ�|O,��-�$"��	�[�&ي��a;-Wx�[���J�X7�i���q=�V3�&6U�*i�J-�Y�ϯ��+�6��Z�u�c�i�t��u�V��T�������ӽF�bI����ꦈ�[k�;�f���Jat.q;4Ij��}�b�F��q4�4�v��.��3�)m)�t�m��oo�t�6�b�ft��?���f��/f�	nqK�5�mK�d�H�kѠv��\nd�I������U{l��H�9H�wx�Y��R�z.s��+���J1sM(�0Np'K�a$�A}��{g�/�.�溶[�U�ۦ��`!�y�d�*�^���z�Vf���Ѿ���*u�i�y�W�|�b�9�/���-r�p�]�@�i����:�+���ܦ����Q��{]@�P��{�-5o�N�kuTrP�M�t�dl<4�=k�Pv	�Y{�u���b�Ϧ�F}�T�ޱ]F�◦��wr�$�c�FC�^��P3i(���f�V
���]qW8k�v̸8�54G��Oo6#�F��.\���I�q�)�C$��r8ӻ��o��/8Gۊ�eJ
peD�<f�ڹ�AS���2�)r��(wf���Y|T<�)�jY�8�Y�;Î��ӡ�mp@����[���+�^�r��ڏVe���h�5�O��\51}�h�:�d�T�R�Y7�ȧ��Z	b�]�9Z�oC1��g�̻T�v'�(��=!\���KI�-�j�I�R���9�����V�s-J1�o�V;s�Ī���
m5��T���{ם4.�w((�hf�P�w��.7�e垭X�Np}�c�����jw̰��:���u �J\�Qh���
x�m�^���Vvt����(����
�lsGS��m������X��bʰ�bTÖ����[�Ϸ�[�]��+I�J�=	m慊 y��c�D��tr��O:��٬\��,�7;�+�\�@l�ƴJv���.ƞ�^Յ2R���6�!�kf΃�Î���f|�M�2h��Wl��]@gv��;�u49�w\�V��y�ƅ��H���-Y�:�Z�%5D��B�Ur�8�+��m����U<�4�p��U�A��c��/RǢ���[HH���ڂo^���E�Ӫ�;P���iWWU�9�{&�_WF﷛8���5��5|@®@�9��Ѡ��G7ّ̀k��Krb�v.v�z��{ݾo�z���V��8 �H����<��.��TlN�zzn]2���IG�U4��]3F�uΒ��^�Υ9�Ԇ4�_��-,:5�R�ە�z�O��1yK�:�5\A�r�0H)�(�w%d���ְ�hu�c�5��������w���MΚ���t�
���D�u.J��hwd+��NN�E>���y��l9:�^f�}�|tK��fuq��ܾ��}K���[B| 4@�H��F֖V�"�O��l�4U�ۙ���-��eL�ڂ��E����Y(�����DYS::�eei��J�*ԭKm[JűL�Q�CAҖ�m�8Uֶ�@�̕�Q1L�±Q�Pk\�6���m�J:�Z�-��һe�6�#Zj��F��R�ZXZ�TX6�kU(YA�:�p�-�ңkJ��)�]h��n�q��*f��L�ҔF[fp��Qb�K���U�ԥ�[R�ڦm����-���m,��Ml�#J5QmURĩm�)Rڪ�Mv+Z��[-��i�ڨ�6��ն���XR݊���Fͪ�n�����մ�å�U�
�PV�V��ь�R�Ķ�s��mf�!���Tb%�b�j*"�m6�F"�Z�jQKѥ.��U\�)U�kD��Sk�Ķ����J�����DcjZQkciL�ֲ�iZF������Z��i��YQ�m�ƴkS5\�Ukn�S �+�(���b*�JD+QT��
 �m\ww���{οu�2ը;�T�OEA�4\j�Bp�����n�]:q}�F����K����(E�9����>������3I���X��u|=�p���������Qx��w/��pw��qK0w62OM8&s�����V��SЍ�ń���J���nL�~���SFݙ.g��eDz����'��IM�zzW�m2����z�ܭ�����Իi�&�I��܄��/	�t��C���Y�#�R�rN�y<ܥ_X�b�<支�v��\H�_.*f.��������CR:����V�q��1�z�;��3�Ra��9%P,\��$��������*��~���VUk�/z�.����ث}UȭOjpOs\�M��U��کS3�T��a��&5p�1��ިq�gv8�F��-�Ӈݑ��!Rwd���K�>I�pA���Š�Y���櫆��F�pA2s��,�ӯ)S�&g��-�x;�B���{}v`���EJ��R.��.�VH�˱�b;D-�H�J���Lr�l^oW�vz�[�oU5(�Pv2h�w��ޜU��e�c�mf�2��Rf�ņ�rV�u��ݨ���@�	�|�wa��� {��\�.�}���Мv�[����0�Lq���Q%<Ȕv��N�\gn7q)�J�'������`ڥV0����ݸ��5ǠC�(�܉Ow"VWȔ��UPFiǏ�@��N�!�� ���&x.���Ev)�L;�{�Pv'�BM�Ŝ�ŹO �v�7i�����bYہk�7MA�=��
�.�)�Z����_a\#A��x�v�	��{.혞�jɥ�i��Zڭ��٫z9��\q����F|�u3U�d��y"SFe�9���\���������c��;��=8�����ط��	����R�����χ�����4�3⺗�ϩ�Բ����k�^�n��s��#~�m2�q�x��؁o����Y:�T%b�u�
��|z� ���77�R�^]ͭ���v��c�1���<�����]]n��E��>�AR��(|�}��8��B��$�'FS�3�{.�mCb�My{[Q��T�v=�)�dθ�[�N�U�Q�����[������"��Y��T�`�5�q+�}�u壸ũٖ�ʤ�7ܧt�ۋ��qtw�o^
�9ԖM�t]�R^�興L궕�.$����֬�m>�o� ����@ꀻf���v
��[�����+���5�K�G�5���XXVA+���:�C8ݣ�K��C׵�~�V?Q�_���|��ܻ���UTJ�4��غxӧ�Q�p񹆪"v@'�f�e��M�52C����䣳]D����1�\oN�C�V��Y	T�U�>�<����S�S�wy\��s��<�Hz��c��+~}��{��R���L�fDR�X'�;wjM�oc���z�*-���y,�߫�joy#�Jt{C�;��&3���y�m;0�k��vM��A阖��BW�p�lt�˗��"{��E���t�[�N3�q��mCN�T�m\�n+ �ɥ�/�\@}�I�b��z�F�us#A����� ӂ�le�8�� /�cr�,��Y�����|(���%B�\�y;(h%��w�4]bZz�O{R��hl���J���#C���=�s3�]�<k�COb�dۏ���Z#���k[z&>������N�Cw�E��5Û߫ﾪ^�7i�I�S^���h���܀r�b���ߵzkq|�r�7VN�W�����hg�gӲu=���yS�:��-��oM�:�0�v~���#�������'�J(�+;e-�W���f���_�����Q'��:n��u0=��Ҕ�~}�WrS��n�6��4v�ף�3$�Fv�e�E�ocښ�N���nhZa�x5\g�h�f��!�g�޵g!8�����$S�U��V��@�����=�uJ����V2�'�J����yt�[��]���\w�Px%?�Y(V&��>�w����ث;�Ү<z��i�Y��ُ�it�l�;�����t����׽���+9�qouii$���M,qʡ�n����WBXMlL�P��UE�;�ד�V5��Ĕ�"7��3�镟>���X���QȘF��\��6�r�1|fu�{���~��f��͕�o���pQ����L�E$c�Z��������ZDE��/YPo�+k��=޺�9�^�:��~��m7���2K���9os�֬:�c)�C9�v0}V������.U�8:=`����zq�۟��W�{�����`�穗�,��}q���x�cp�����V����>���$o���f�{��;����u{3�e}ņ��bZ|uQ���B떲m��9�ثNL�ܨ��nM���YD�Z���}p�^%d�n!0��Fd�nz�_/���x��j�N[!�����5=�a�P���3��S�8��v�hF�)�J�֮Qɇ�Dy�i�գ��cͮ����Tc\^�[���ܧ��Grk�n�[ܪ[v�y9n4�q����ݪ+㧫~���]|�Xߧ �z�対��[��z�7ǖ��0�u�]c���zc]�N�u��4��Ϸ�����ݡYo�p�氮�t��v����)W�1�b�<��Hr{��f��jz)%���qgz�]�A9�Fx(�������J���Ŵԩځ��f�u�kߋW}�S��Q�W�1u"�
������P�$���2��6ȫNY�ӹθG :�k�g5wf�ƞ���z��+d}��
2;�ud<۾��;�W��^-թGz����2]���a(����>��q|�C	c�W��#��AL3�7�v�|�J9��5��(\`u�;��Z�@.J<ʊZp'�O�Jy�;u|����;�5�G���SN��g�
S�B=.or5O���F�]��4��'!Em���]����F�9��J]p�y��+��52L7ܲN˞l��qP��I����6��uT���MAD��+kwmP3?��p��
����ڽ�5e*�(��b+�}Ey��F��OZ�ԕ��n��3;�!ێ	7W�%�u�Sʹ�̮ɥ��W`(�����k�u}��eaYN���Yጊ��0�&����˙��9F��>���fo��QNH�SpT�`c�L��&���fx�W���ʡI��yosW_.�[���y�5AE��j����]����f��X�@�Kd޷� 7i[�r����<���N�͠���b�c��*�p�'�]'9�
�-�m=������W�b��t���V�¬9Mqؑ��h�"W.��MYhb���w��Wn�U�_����[����R�����՘�^V\`O�q�-�r<�ͳ�>��J��I,�Goi�8c/".�jˌ�7�c����ң����(Y����2(v�����s�8O�&��!Hm+�5U��qv��@Z�{�h����#�*������V��9�-�m�Ou���Φ��ķ):��i.����O<�aKrl�7�,;����EQ�4�'
؜�S��p�8�Y��er�K�q�����@��n��*�����M��k�ȗ.5]8LT_#����>A��V�	�Lb�w6��H+���pp4~�J: "'�f�osQ��ѓ���cc�!'zƧM�v8Q���]<��kÕs�K>�+���$�Ξ[u��%�ȑǖ�KPݽ!�s�o:Js�������̘rnF�.[�P��Va��k�>�ǧ]ƒ*��;�bj�j�
�}Y\!w�e]�XWo�R���9*5��vG;�m�'h��3��-@�g�%��۫�����5�M�������+�K��]��C�vj�c)a�����">n�[r����s.4r,����X�����)b�M��%��J�ȵ�t�&�����O6blw0�t̵�d'qF�_Z�MN��2VM���V-u�6,�\�l�V2:�m��!�6���0MB���庢�Υ�:��W��f��z�t�i�W,�l]��=��ǻ;H�8/��xC�@����Eb�߮�7�Zo>N���ޤc���+w�_D[颰e򖶇E�nV�C���k9��F�s<�PΞ��R��VE�ϧ�������W2Ο�:N�ޝ��,i���t��=[o˩{i�-���k�I�o��/A��ͷM���d����u�u�����i��җc��m��`M^3�Ut�PÒQ��1[�(��5t����ԣh����k6|���6R2Ɛn� 7GU��O��W��u�O�*�n������/��j���{F�����u�t�)��2�N܆7;��S��uqm�������oY��g/��6lU;>Yٕ�p���W!�rL��,�[x�I���rx��<�x�M���v�-�˵t���nOèJX��8�/]]��&ټͰUfsT]������5��xF�P�D�q�$���G\�ݧP��U�f,^ۇ�mp�Y�[��N��z�dL%	G�ݲ����(��M��Z9���v�1���|�t��݊�认 X��kEѫE��Ug��E�]��MY�(��JtQ7+��xd�{�:Pv�k�FtޗRR���z�
�r"�mƧ��J�,>���rq�xv��|;!��3��{o���fz�v�&�ލZ�\:��ˌ�lv�H���[��Z��S�B��ű�(�@���������݂�'ee�lf��r��F;��g��	[}��j��j�aS}��� �<�p��oR�Q�⣎7�5J/�q���NAm>�U�����	���ѵ�G��[��9��k	���^�pK�Ɖ����kNbi];.m�}����1ʣ�#%���7W�L���t�9��;�X]�7R}V;�o7/$�\�Vj�BW�ל��QWZO%-�YV�>�Y/�1B���#;(�6���#��.�n�g�q�<�h�Z���5Ւ5�k��|g+�}��Y�X­���9"�o3/=[�kj�o�ۛ�<)Kϊk���m�o�����b�����䯽�H�|^Җq��m����K|����՚�(����˳;s	��̲Uq�8Gn%�᥷�zjK�m}�Z�Ȏ;y3���WW9�i��l�����Y%c��9M�콆�T&�:�����_���ެy^&M�:��\�4'���X�'d�"�rӲ�gCͯs�+����/}=Ȯ�Z��Q�v>�N�Ƅ3jD��I��l+���ڛ�diq@D�拳�Ք�����KWA��}5�(+I����*4�4\L�%�ȔwS��j��ʊr��:F�N�Ko{��e*����]7�{	���Oa��w����(T�����r�)sxtJ�f�fǋ�� �S,�*��i*�QUY��7��!ԯ[���)�l�ұSIg�G���ǰX�t6��MV�R���5�WC.�Q��ɔC�.����b����i�m;8�1^Uۤ��A
.vV����;WO;T�z��4�]5�^�-��.;\�9fX�EԦ�n���Z�Z�j�M���5|"�igZ����<K;�c᪆��1+Zz�Ҽ��������;M�P}m]:�b쾰�eػ��]V�/:fi�t�Ϲ�d־R�ͻ+O,[r�aЏV�VsA�{�ܖ�P���W3=O�Z{�V�W킙��@3���O_��;��RZ���v�K_p�[9�[(f�\k�s�NQ1�����N >Ka��[z�
�H֪lb7f�U���݉��~�-��bXX���)�쉙-r=���]�vo:�cK��nN�4]GA_T��$�ƽ����H���ru,b�M�}I��h�ê�e�B3�Z�z��.��2؈��}-��]ש�;�oe�k���-�#�Ыt5��GV#�)�k��V�WJ]ZS�[vB�c�W 鷵�O�v�XrԔL�ϚyDd}1��|8���D��"u%B�H}���j벲�f�{"�%�F��)��l
���a��̥ہ�n��[MI�a^NbWh�CT�+Jg�5[���ƅ�ϥ)x� \l�`�o���Y�t�W���V)Ög�7�0��`����C%�?�y������������X��rYdB�^(��o� ����#{
­<�('��o����V�9=�7 ہ+��Ξ��cY�if��U�+�K+�+��\���[���qd'�k�}1�Y�z�V�AںYJ�i�+e�в�y���[}�}�}�;{�tCK#^^⩴�|4�Vk�d�6�:A�+Mv��)_6л ��e��PLt�ɛβ����;��w�Gf,\:�V��{F��muu���n]h�k�n�[���;EZ�J��ò<��*�qd�ə���W1Hv<u�i��!R:�u��\wyN��&�����l�}2�U��zO.]{�}*0__LJ��=�-o}!"�u�tܻe��9�<`6�c%�~�ܨUc9GI�7��
P�r%�7|1t3�t�;s�Is68:�yC������ttE|O`�v-#X)�\�:���Ψ�o��YXQۙO�s�pCy]\-�Wu�����:�r+��]��O^6N+,h�ɴ�\�&h�$���b�z6�����!�k��N�[&�^��3�^,�ʍ�d@�m�u°Ꮉ(z.F��e,��A4�s���yw��-����7�c�ܾ��<�)8fqq��N�-opB��Y�D�δ8|��F��YpnT���Î{����^h�{CK��
�Q�J*��lb�����bjҫ3���m�֭h5���j��Ա԰�(���)lT��ZV��2.���Э(љ���ʖ��i�;5DV�T�V�(�m�5���PW]e0�[bYQV6�WZ��֥�,TQADX����fe����W#v21nB�X��J**$D0��E��%�h�mV*6���6�"kTTA\��A�f�P`"Eh��\�X*��+�u���b[DQUPZ�Db�`�J�Q]h�mU��\�5Gk��EX��ՋXU�¦�K%�j�#m�UE�d��EV-�PQE����R�3PF��"15X��D`ʒ�-�5�e��*�-k5����+&ch��V#��3E-�ړD1�R��jT2X1U����ج��+DUEU��AE��SX}�޷}��W �Ok&'y1_q[t��]>���|]
�r����v�j9�Єa��U� �����Bq+;h�N�����;�ZǿM�.)��rf�����踖yѷ͓֞}�ݺ�XB֝r��u�6��*�w^2���]e��q?��[�=%�Th��q�j3�g8�¢7�ɠ�46������H�&Pq���)dʶ��E�+�}|M\k�M���I:j�RL�.��1Kp������C�Z�T}�F��ci�Y�G�Y����ǆ^<�ΞK�_���e.�a�$�V�@\�j�m�Qn�Kch���B�;����w���f��wG��K�{���ʎ.�ŀ�}�u��yU�Ԁ[Qժ��4�6�.��p����g�H3�"�(�^b﷖e�/����ͣx4��9�m��)s-����+��ń���TV���D��r�A�D{$W,�&�2�0����ݐ����Z�[�^ݙH�X�	�r����p.F�ͻ�zb���]�
0�Z�;nC�ͱ�n`KT?r�T��];��T�)D��*��U��+�\;�&S��S�>SJ�ih�z���Zf���O�]�ҭ>�ͽ��Ck���"ף|����aU�����	��qF|�����9A�o.B�{$���ɽ1U�v��I��L_OA� }=�6�{��$/1�1�צ������<N'Ӝ�է��}0�L%P�C����<�3�1�j����^�|۾�5s���nu���� E|���N,���y�9��θW."�w��qe���y/����j�u�l��F�]��k�$�U��+#X��;���,���0��;�ǰ0�q��3vȑW����0�p)��{4�sME��-uq���G�p~�RG55��4�Ҳ7�T]��L��5��ڢ��XϏy`��qMN��,N�2q]ks����zb3b��+dތN�����ڱ���MK�W�hb�pp�;O�:���F<���e�����hZ���L��q��acO~`�^z�F}�x��:�#�t]+�p8�t��o)F���w��^sõ�z ��eQu�b̢t�|<�sS���!��z����驔�}	�/Guֶ�8���:�7��<�J�+��ew9��opY�Ҭ� ]���H��S��q^�=)I?���N���M�{�x��t��8z��V;�s��K��F���u�{x{a���p�أ���|�o�)�ZwJ����s;�_^ۄ�ەi�g$1�䚗s��}�g']�ͧ�|���{����j���lY��ԯ.qz�ys\��P��du^��d>ߖI9�ަa	SwVe�J�f��'~���Q�]�k�Kt��:�d��&��˺�C���o.]�����o#p��k��y�j�]]��u��6ì��&�q�~���qyF^�����/���Ȏpz��Rv�|ư�a$[�Y�g���^$��'*��yfD��#xQ�g ��^�mC���-���.��������s�/>DR�(��Er����H���v]Od֛{W+H��xtZw;�չK��S�ȉYQņ���.���eF+���AI-�kk+2d8yv$��,��$��i�[8��r��]��E�Ĩ�w`s��Wspr��� 0��ߠ��}�VL|�u����R��晜qf�.�^�Pܛ߫��eWK�69���\Ud# }I�M�ܡ]��ME��Z�f*���HݐK+r.P��r��>*�B&�-�܁ی�q���n�ORSf�������9�|M����:w�L�h=�����I��7�S3��{j�m�kR7oa���qqf��V���;��^��~�8�M���z��3::��r�ޭwڠ�Ҵ��;�X�f�-4@��i5�~1E��:7�;���U�u����ԥ/oϖSo�ڱ5�������Nt3�֜��t>О�0q��=�s�ϕ�4�sR�=iw-L�,in�o\'��g�땺;FZ�4�ܗ�C3Ԯz:
c�7����uI��]q����i��|^qR��A�~��>�T�
�T���.*�qY���m.G�{�k�ܛ��X�nN`�^��4��V�5�G �ֻ���a����i��]�@�@U�R�o���qڈlO�ݺ�*�
�Z4Ӝ6���,�t�1x|������fb���閟5�&!b�wWs��K��v,S�j'�$f��{�Wm52N"�#��f@��zaX"�w��ﾄ�NS������D�f��S�M���j5���D��C����G�B�*ql���:K���uSU_D�u�M�˭��#Q��,&L�=7���0�P�v$Z\a�Ļ5���<�I�H�L���-�J;q��/;zQ1e'����+x��Io�/�mS�p�Iq�Et�:���D��#Z����d�M�YP[i�p�p� �{iɞ�ŮAB�qZ^�)�G�,�e��}
ɠ��;���3��C0`��Qw7|�b}��`��^��f�\*7�N��
�F���Q�]:�˹�FtncY���%!/�e�̀���5��r���6��c[{ϷU�Ӵ�VY��Ҧ�,���dܾ�VcUb�Q�1�Js���:�5������Zϗ�9�����8��e�x�Ҵ�~ �xuDl6�պ�접�(�d�x��g?��}�����x�K�K�Ĥ]t�݋0���s��r�73�F�mp��#��1�Jw�=�@�X]N��S0f�,�ף/����Uj1;jv���"����G�&������PO�Z��O(�}����Y�V�N�}qE���*�#�6*��֜Pl�R����:�u�r�mUqok�V���6����I�L^���+}����lۦ/J���`�{F𥄶�o�'r;H�sl�]d�������}\���o�L.F8'���M�).�R6M�SN���^�q�j��P�K�%d����}�����!�q���l��.7���Ć�N�ZF��rKB��>&�b����On8L�n;�.�yJ�`���K	�r��6�3�6�8����f�V����9��{cVR���Z;����E���Ǜ"�{�ٗ%w��J��3_'�m=���B�v<u����gqjk��W��к��"�m^�ݑ6;�VS�C�Yك1������;��}�n�U=
�[��}��YL(G�ТsxT%�u�Sΰ�H_�r�2���ݤ<�FNݧZ����*w6.՘)a38	�����k���F�:}\�i_s8lG(��2�+�w�z1}oH��a�WvU㖵1����<���t^�62ű֗R&���\B��=��F#7�7X��{;"�`͇�b�_٦�ފ�Ů��[����h�AYG�Y{��4�A�����y]+#��n�ޗ9�m_X<��w�q��k4��,�f�/�j�Yh��, ��{�g#*
�:�熹��)��N8r�Qƛ�U�;�`��M�)ݸ�_L������s�7��'i�[T����qud�՚�oi�y�~�u�W&]x%F�%ϟt�?��@��m�}�5_�J�>�Jo8�M��65m.�\�t�wM��U��߲{(����Ʋi*w:�||M�|�zRޚ-�!W��:U��O�;etʁ��7��͠\���J��(�ܶ���=�M�v-�2�bI��s��@��WӬA�=4�Cƻ��X�GV��},��w]��A)B]=DT�nzJG��j�c������s�}�����B�{)���I;��+�����_�t�:�^�+��7/-�Ȑ4��N�v]��Jk���7S]q� ��5��"�ɣ�\_��lu�C��hЬ�q�|�ȯ�.<����^�w_<�앓��-�Me�겸YM,�E�9���t���&,S":TM�0��%\m9}Qʫ�l�}(���{����oL�};T�����"�V�TS�<�qZ!�@������K�d�����5��CK�z�gX��Ŭ�t���׬�<���B`G��-ȥ�j{��>�t�T����U�RY���oYȖ�d*�)�lE�2�#����x�v���_X�QG����=��由9�l�y
�!bKc��=�5�6G����ƶ
U�?M��x�N�G�x�[�vف�	Ӹ�0S鞾�6�6(Ǘb�Ǹ�/L�����v�K*�mƧ"�W�q����c��Xʉ���G!rܜ�-���8���7�^>9�1��P��+OI��
&r�Q\{�P�D�EP���5�f�|�T���׮*8�B�X�۬��,Y������FYJ�ک����%����?0��⨪ۿC9�'���;."��m`����L$�.�����<���rXS�59�ReZ]݋N�����7b<X�="�r�x3��3�����ΐ׶g��=�n-�q�'���|#�]zO=��p<�/D���4��Ev���˙~b���os�\�hy2n���O�0h�X�y]}�^6�:oo�N��}���-e3�P"����tSV��N+�d_3�k�pOwb��_���s���}i	]I�f)�x�ڝO��D�r����̵��}i�������y��(gE�q�;�o�V����u%*�}�[���WL���w[1�������Q@��=�r!�U�t���}0MA�-�D��.���v�������7oHp7�/:Jx���Ҏ�b�Mtp̀ά�������/mc�ws�9QŻ)��/S�C"��7-�/3�bQ&�w)�6wm��KF�%eA6����d77�v;MXzsv�ln)��������,�<p��	�{Ӽ�·Җ5B%��w���(A�ŗ����ZD��9 ��w0.m�,X�Z�kX%�����r�WWB��d��|�"��G3]�{t�Jw����h��Y}�+�ʒP�J���J�p�8��R�H1.�>�݌ok`Ȕ�(7��N�m[Jr��o���<�Jm¾�b�>�r��w�4���jɔi��~|�|���v���h�ʭ'��=|�Wێ��k�i�M�zK;�ll?�gj��z���d�}�'s�������B G	�O%aOJ0��֭���RS+9(�=�q!Hu	n��i;��}��C{�Q{K����+x�k�=|X�\��m-�o��p?mD��\~�[��ex5j��j��)M��B��l�����k7�x�ؘ����z	�S�x�@��1�U��{F�#
[�6��o�[���cf;"I�Ж2��s��LnJ�\���W����S�)Y���o;�������n��OJ� I�w`Q1Q|���* SPn��X�%v[��^C�]���񼓡,�J�z@ڹ_>þ].xa�Wp�Ǝ�Ĥ9�H�RΌl$X�SƐ����jֽ+B�{�6�3V�]�U����[O��}�;K���է��լ���0d+4�Y���nn忺�tj��R ˬں�]��+o�&T�J��i*`���t���>�ٗ@Mw�Eһ�z���8XVڶ�{8��^+sG/�Y�Kp��C��^��:*��p�pe��f��:�2��tӒ�L��� �:i�����]��4���vvT�7]+�ᦳ[�ܝ�B[�V�&���i}�Y��a��N����C�<f�$�\�q�.ㆴ%¶�w4�]E!���p5�[�u�����J���������&�f�ԦMWr��oX��|P��a�ʺ�k���#K�U�[/"�=��75�&�q=+Db��	MzC;횱�v"**�r6�+�
�7õGDW[�)B�wg�}"H���NY�)SҶ�gi�Fl	Uv��%�l�s���n��#�U>������[w��B� �8��n<7��R�oD3n�����R+�H�TF����֬��V�#.lUpD��R��5;	=����8�븒�m��q��+75P�ŝ�X�Qp�[�qz4�Zl�Z���jt�UN���8�*��(pK�H�n։�L�K���O��������%!6)��;ŽQ��6�C�	�k�����f!��C���㗻�v��W�.��hSg���-Jz�nH*hGݛ҅��zs���&�j�O�Kp9�S.�<9r�-$�t^⦶\	5Yx�T.gX��Ϧ7���c�OY�φF��_(��9�wWx�Q�g��X��lѥ4��=+�ז���9�o Z�P�:�skj���,n�fҢ��Nٛ��Ƌ�o��/9Ϡ4{:t�,�m�k�9��2��d���K�{L������
M��L�5� �$�\FL����6Z��� �G��4U=�M�,�j^�+�J͘��k�-�+[�.�)El[�����«���Nn�
�mk��Hn����[}y٢w̷����rخq�-��t�(8�o q�_Ny�F��7�3��*�ȻH淗nY%�âPئ^[ѕ8���e�K
�����c�!�
�Z�I\��8�V���Ku	]6>`vC1mu�_kT��]a�%1�e$�%H
W�Gf�n�<�z"m�guA�*u;�R���I\8[�3�X6��Y���g������6����*��t��t��ow4�ώ2��%�!3M�>�[�r��X�X8%�!<SJvw�V֮�%��)���,��D�˻�k)N����k�(�r�X{��;I�S_q�f�fp<�Wڸ��jw:B�*'�*�������DD���ȃ#���e�Kg�b7���χ�iFWV�{B�]��}Wt�Y�-+u��L�����Rp�6Ty�U�������}�[3f��X��UI�eb��PTm�� Ȗ�0bԪ��QUUA
�*�S\̪�Eу݊���B�����XeE�*�Qe��[Z��:�A��֢�V ���+	A+Qd����$Lر��6�E6�UUF�����Ĵ�TQ�mAU��
�Zъ(���P*QQ����-��R��҂�PY�YQV$T@UVł
���VATR��Ҋ�֕�EX*�#m��F�,���[J���T*",�,DQTl�ZUm��Ŭ��21�Ă�Q-�ETZ�V,DQ��J�TV*2��1F�(���X�^.������y���NQ��f�nR��r�76��O&�xހ���Zc�[ٸ�mv	n��ݢL��/:a͔k$�<�|�h�ug���jm2o��}9�-Zz�d�U0��?J�s�\�7���WN_\i7�ju���{<��W�|��]
�J(�jl˒�e������F�ȣ�r'�.K�,���ǳ�j0eg�)T��zܓ�!]����_5������z)��NّV�"g�n�����ǵ�P�E|[l>��4�[�Q�]_-
�du���y� ��sMf���_�R���=����S7Cg�<���-V���^ѹʸWY�CuY�C�z��y�o�5<��hˏ�-�r�&<'���#.��sv�]ڞ�Or���q�q��:���UD6�����wW5,�����zSD�a]E�7�o\k���*�;	��Y]7v]��(���-�wZ�/.NXx�)���bQʶ�R��Gv����ڊ�6��b��;u��nۭ��(i�'Q��K�+N�&_=h^4v,�`�`h�	`�{t����8��z�U�r���j�נ�Wr�:�'J*$�KࠤM�yV�������`s��+���䟖�P�H���m�K�0��Wv����ޥ����s��/�8��nW�Оt^�!{K��i�kW�|K~�:����J]�І��z�����P>��m�k|�r�斒OwqD?Q�ڇ{2H�oJ�"��֠�L�t��웮���g/�cqB*�l.q2�SY�w!��S3r����)bU՚���7n>z!c�>�&n9���/�����G�Vr��ܛ�w���Jǥ�-�5B��˽W=��3랄�_OT�ʤX�-���zV�1*�&���|���j�z�-�auLsG")s̉Gv肉z�K�llU�`�s�S��9��K����hLg�]D[��.���f�g]e5Q9��vhnvu&���[�Oac�Rrf���Qیrg��Yz臱;@�㝩E>W�*	��b�P�*t�����Ϡ#����;,��.�e9S���\���.:.4.����BH��]z��6Xz

,f��*��W�<e���;s��n�����m)����f�#c�ss���܆����sr�-tX<�M��Vĉ��󶸾/f27���.��J�wg^*5슍N��W��ϓQ=l:��(m��8scs��Z�����^nl^=�NEF⊎8�5J-��\M��o7�/�|VaY��hۄ��Yˁ�/љ/�9@9j&*C��=��9��{�����[C�������Lk����X� �ks%ƜJ�-��T�%%ﻤ��6��{�}�����%����k�\�Q '��#pM�5Oݛ�r[��ݞ\�y���(t������1���������8uU3~qc픱���{`�n|�J5L*�U6/m��u"����`tq��\�Ts����>�I��i���k��@2n�\A�����Tls ��Z��Z}�{�tW.'iD�uKZ�(�/zv��o ��q0M};�P˭��"5T�
��Wt�lX����!P����n^��U^��z���S��;��s[��v���s=���!癍C&����eK�D�L=ko�P���	��s�\\sx��73@�]H7������$k�c���=��NŤ�.Q<`YW�$�]Vv#`���}���}��-Ra�10~&�UIo���yc�A"��<\d�o8(�&H�����I)귺*R�(��麭�y9�p"���Or%�ܗ�[�L�ϥ�c!��O6���'�*_YL�e��bʿ�Ȋ����B�=aZtӇ��y�a�]�q�`r�v�qJY��_m��ٸ{�65:&´h<$��ˢ�^	�j��$"�fM�/>�gDkhOg�O��;���N3�N$���+�u�AF�ߓ˿����uC��ڨ���<��zH��M�OxI �S;-_����ō�re#+��u"[�Xmit��c�:�������I:���q��rjK�o#��i.j=��l�f�g�z�a�;�j�w6�����(�ݵ��]�i���\����ӴV�B�6g���
��8{pW%v��o��H VCλ{��dc�po,	\�ŻژV����
�$��w۽�v��ɮ��4��ܬ8���/v�HC}�X�Y[0J���{V����Z ���tH���"�_dJq��N8ܓ�O]1�^W�'H�)#^~�t�7����Gh{�Fpv}Tx�����ڀ� c+�_y\�.Go5c3�%!Wd��vi.]��o��XVDI��!@��yF��;��a�Ϩ�O9��WwXz�@m,p�����z�o�;���R�@��Of,v^�>$�3�yF\jKsY����d�S����W�z�dD�J�zb���uuK7[��a��y]Įy���H�E�}%�J���J�E�`C��mS��k3C�j�]Y�K��Of\IuYx��K�3�Q�#U8��g��WF�â��LAGx.�sK��=��؎�2�9ޚ����{�]sYa�u�Q�lt������4��<����3�YZsދˋ�#�>�H;��3�*�h`���쿁�/~�����+����2A��;�L�6�T)Lyc�e�rVhf�u�r�����/�s�B��Z��u����c�ץq٭`V��]t���!f����n����z�WN|�X;:��_u�0ւ:����*���w v��q�I��Ȩ�j�ڿ�����[�3/�����z9�å;��5���-����k���#Վx����_�a�M|Ve�|�z27)c�ĩ�٪cV�[�y�bߩu/5������w(�jv��B�6h�g�d���;���<}�s(������ρT�u�M��ܙXe���'$diz�Og���M�ng��hO/��my�s+�����o+���nj�G9�d3�9�w�NĞ���+Y���w����b�j�c�����p&�i������؋o����]���;4��՗+�M#�ע����~L�������\��n��V"��9��y��S��Ÿ���C�ɴף5]���i�+2�͊�H����l^Q�m�T��2~E�)d��sК���i1Y=�u�ܧ�S��ӣ�?X �އ��U�-VM�a����S�S��H�$�h�4��t�/�Fyg%���l��#b~P$dm�Q�P�e�(tWlU����T����`�\��yM/�1����f�#CK�-(B]��C�晓�Q:J�j���;�:��£�0�D�u�#�\�"%ܔ�A��]��jV�9�/�5h�7�{	��U1_q�/mȥ��ԫ�q�s+&O^g{:�M�k�\D��B��p��E�&go)�"���E��n�3b�/W>�<��>99ƚg1���&� w��`���
��5qׂ��?�1�bB�5l��N��m"�l����Q��6��&�)�d˹]�S�ݼy�������"���ٝꕔ�=�f�8k��Rgr;�Rvr���a�<敉qT����O(���k�Tkg��;�"R�ϗ����)����P��b�繕���>R�{��{ݧ�OP��\%D~����׉On��d���gt�;w�T��)k}i�`Ն9�ˍ)^$�v���'���7�(�Z�q�Ց��b��F�!�}S�v�&��
0�T��\ܴr��98q�c뙖_�� )}�&���`[��t�@I�f߹���(�J�]���8���]��5��跶X������:D�,{�v�e�YmM��xY�&�����}݅��^�{��<��qc�x����o�g������!j���O��bB���Iah����[���Ww���M?gN���`ΰ�ޞ��%bw=�[��#%\o(�b�3'�W�%DJ�z�놆?�z��\x�
���ʾ9����QnR>�=*=~�JBWH��g�R��SP�9n�T�b�E���^��l.��y�Cb=�RX���\�`O���G��@���u�w��b��]s�f�ڗ8��1����3�&2!�q��{�G�Hk~�>���`:+��>^��duL�/Ox���V�~��C�5Hs�z����z�~�^����Ĭ���'֥����O������`�w��G��YCuS��s��Ͱ�a��o�y\��	�[=>�����e�<7"f��9��ˆv�D#��B����s�w�������9KRC�Ȥ\d~�=ܮd�ws��Z,M��7>�R{B�ݸy�����!�+���(���4���y۲Q�dga�6�lۜ2�X�o�V�7Ֆ4��Ty[pu���q��oP#{o.�2�+mu>�\�k;�7]>�Jyr���C�pݨݦ�R��n�6��ǳ*Z��d³�+<���F4���$�iĮI|�V��̶'c�¡�fF��r���S��>��;���~��ّ��x]�L�/��u�Һ��z����GD'\��4zr+�����d��eE�V��p�g�|]ϔ�C�צ���𢡄s<a�7�H�ض�vj(�YDG�؈�s�J�ƶ}v=2yU}W��F�w�Gs/T�*l	?.V�=��2r7ėwӳ��۸~���,徇�݁ܐH?PZϮ�Ӈ��j��
?uZ���ᾜ��\R�˹�������[(ׯ��8������Voւ����S�Ҝ;ǥ[�,n�U��dӉ���9�rx���~�g�+������W�=2���bd(��=�Ȱ�m+�h��-o;؜=�i^����1�llx�`���]7���=2����D�b��^7�s�^�k«[�5;�@T��F_�pr���6"}��N��c�^�v=,L_n��F�ή7�x�}c�͛v. rp`TX�|��4>��
���{:*�N�`w;��/d�A��^��#_	0ۺ��
�P�gk���|�wB(�[BS�y�n�>�Ʀ�gJ7y�n�S3��[/h���3\]��p�b�ط��(S���o&��A�f�� f�j�;��t��cC��gX<;okeFb«+}�
� �슊���@E}l߸L���>�*���aߞn�0a���8�3�#�p�Kad��ɓ�߫��w�4�9Pȸ�ME}l�X���yF�dWj�]	��?�����������h��W�2��3�޺@dEW��
�rr7�����0<�e7z^f{S�P6=t���n,��� ��&mj�=�ᷠJ�6:+�i�(�~W�����?b�{��;��q�7=<*�49��������Fx����p�����0�V���_�{���]�]u��*�K��JԼ�����]7�>�^�}��n
]�O{ֽ�$b7ϲ(������s>��}�O�����F9��>��:,u_���Þ _��;����[��ı蛹��Y�2����K����١	�nO�]�H���묺��:��xu3�˘�����	�/��x����sw�}�jzs���� �˛F^��Zz�V:���e�}�s=e����<��^�G��dt�y�Μ�~���2{(��^~��2��3��;���Z��R{����n��ؒ���ݝx$]��8��J�]��Z�wf���z�n�V����{`��khp�.v���Zx	&V�����\"2 M���^�O.�v���;졍��k˫�H�mv�9oH�)�z���z�З/���O3��9�h&��J�F:;c�s�����pd�j8�E�lЋ�QU��
�A�W	��EHs;"F�:̥�BT�.ڴ&�/w2�Ci-��Mڼ�+R#)�x��'I�Hٓ)ku��i�g|�`�M}�!�G��!p�f.�^�vd�rmAyԣŘ
�|҈��F�����1���VT����<=B��ǝYy�:�s�8�� _M�w4F�hs-�ܜ󷯘mj��::��M��܎�캏:bT�Vdv��l��c/�6,�/8j�&�͹�,*|��f"���y$W)��y���`x�X<�����7�����X��s[tm�]�$^nӖ̭!a';�����d��B.�z�����+��p/��r���7G�^S����Y/��Y�dj�q̴˚�J�m�N�=��7}6��r������_ҷ���$J���g`�/�W!�@��S�{�����cvV���(�׏�+�}d� w\l;A�G�69жuk�3��{���U�Z�ȼ69wJ��
ʼ
�5f��:ñ�>Y����V��+j �ل��	4J��z���IfhaP��C�R��7�4ҥ�u��e\) f�+�)R��6�@�)��N��� ���@���YѼ���k��vd�%�
�5�
�b��]�Y�����!J[x{-V�w1��QT�+7\��2m��	ȩ����K���$`��I �x�Z
WY�ى,��k�+��ES�1�ǖ�9\�M���<�[iR
�,���#1#S��V9)':ݸ��㛵*M_�n��.���<��u&�\�W6Y՚�A�եX����%�(��s⎃)��Ĵ-4ӎ����c]�M��]fӣ�YN����v���;�7A�wz>N�yi|�s���ՔR�f�׺�=�կrZs:'I�P�f!Z���������)r�X�e�z\<���+l�+;��/`i'p٘��ty��|_oYm"fۂ�/V-�lrc
̤c�z�U�XS��~��h��l�n�p}yH78��b��"�t��5`��R%%v���`!qHAM�Hn�$Ծͤ�-J�)j�t��Ǭ�e�mr�o�j\'�o=0����S.�
͙��d��x�+�5L)��2�(n-��-�9l��괎�u��`�c��]%-)�ym�*���t�]�ȗ>�:2��/{BlqR֭��_S��U7���		I2B酻�$v��F_v5I�ݾ*�w�	wvK90KyD8c*�"E�aX�*�!RV�Q�b�A�����Y*���UF,`�(�E+TV"�"��`)��X*"��*���FT*���cV�`���H�H�*-UJ�EDJ���
"#�[(�PU�TU���U�*,P*
�D%J4eQ*��0U�	hPF�X1�(�1U"(� ����,k[h"
��1E��H�"�Q�BQ����"�"�)`�Q��Eb��X�
��J�A"1B�PDAE�eJ�+[`�DH�#�*,-�,EH��*�1aYF,�E1T%��� �EE������up򅆚�#���մаsPn�pK��?�Gb�[;Ost�
_t��qce���F��wW�R8;R�$��w.���~����FF���!�W���K�!�c��2r��h0q������%�wG�%��6�����Eߦj���E�O��ۣ+<��}�!^b3}
���S {=q�3�U=��QbL׶:�����"= �I%��M@	G��nFړxW�MN��9ފ,V�x*3q�}��4��N{�~Ǳ�ߕw�C�[0�v�D�R��CۿG\��d��Pl����Wx���&��=˭H{��	3q�˩�^�YdKU2�.��f��`pmP��Y��U�+~���{�c�����&��}�����۩����
N��
}y������c}���1�W=�|y���=<�p�h��.<����9��ned?vL�c�C>���_[%�����u}R�1rK���yؗyO�M�>�NAv����;�eFo��|뢄z��tS�&�����U�|�f�%�e���oefӟP���H��>J�\��{#�U5�~�~o�"�ѥ��cV�M�1���B���ePDvW\/dm�����^�]��g��g��������2�qF��8}!D�J����%-�2���}t�/���7�7{'�2�_�f�tg�c���:L�ُt�+��)�n/��e9�u���E\i�xq.��Z���/Z�;jH�k��^�	ݧ�Tɚ�o��ԗm*��/#�ܝ�cc]rͺ|��M赵��+���+O`��	���x�<޻���:�w'���h���Eq��g��ɜ���r�zr�>o����hp�s�����셒�No���&��נ�)W����Yӓ��<G��}�N���z��E�WZ8pJ^V�7��2�޿]�^S�s�+G{��Q��W� �\�Jv�>��pq���~Ր��R�藥��9Vz��OwR+<@�=J�A��͂ǧ �F�Yֳ%lp��Nǽ�����7�z}#�jfﳃ�2���B7�VR\Z>��|߀_5�@u��V�o��l�;��zOZ��.U�v$�}=v�[��J��s�[/!�:�up�>ʸsQm�#B�}�p�Ӱ��#��Ɋ�q9��lbL���a�E�w����bvLC�{=:��0�D�W ��,T�Td+S��=����׺������A�B`�a��=��Mt�o׳�:�C�"e�q���i��=Z|�U�����&V�1��/�idVE3������C��츇�/2�7<�t�vb�{�H�>�;(��K^�h$�v��F"$��-�47��N]�e���ɞe�=G�ޏӇ�o��t�֧��G�n	����<�=����w���NE*Iրq��OV*�id�w*�2��ֻ�#&ʞ庯�cDF��TX���\;bC�pJ�9����B�*^��_��^��R�߼/�@��+\O�+� ��/�ˆso�E}m_XϹפ��iΥWA�B~����T�m�t�ۙ��>Է�֭~�nP������9)G^�V�-����ύ�z_�1;>�Ț8F���Y���WvG�����t'�Н�`�[@�Ȋ�'�\�;��{���5<�T)��Y����&�{�j8�}۹��j�'Ơh�~��z�]h,0�S��ps�b3)����Ї,jڌR���}�NY�3��=���>�^����ƬhS�;E�m��g��G�}���;3��|}���g�ީ�V|z���E�M�c�#�l7|FAz�*�Ӧ�8������^�өz�G��ip���~�����#j��>�S<�<��M�/]&;M�G=[�lJ�����x�����2y�#rB@���r.��_ڲ��mW1�Up�b7=$:��)�M���<}|�܂�H��O���K�8`���/�_؂����R��g���D�~����W��xGb�,e����vP�';�5��v�-&��P���m��T�
��6LіQW��̽�q�g��[Eog�ޔny��Ik�2;�}��%:���+���e�]n��d�7��l����s�'*k�����"y^�]!D�K�(��VBG���)GY9(;�C`���z}.�[�?R��ȇS4��]2}Y��3��n��ϣ��[��\���D��ﶮ|FDy�d{b��<@c�/de{}���.�a쉖����u�2MC� e��zd�P�@�(t��v�9W��O�؍�k��xq��q�8�	�ǲ׎>�����xX��è��axb��J���4+��AױN��x��U�b����1=��n�M���d-��9�EB�R)���]]���;HzA�/�}jsog}������w+�?/{Lϻ.6z1߆D�*h���E禢�-���9��}Cu3N�Z�Q!J}5~�g�aU�̬�{�g�  ������P����n�5�U[�M�5C$�V:^�BX.=�{+{��|����<�*���'�-����'1ݘ[��y�9䯥dmw�\GW�
.}�-]����Tg�1��#��]h��O҈���Nw���$����xvW[��ճ����|29��}��l��ǧι�J��n�1BW����v�g%+S;�ݮy�hM4�@C�^�y@�R���]�����n��꘩ټ��DsLN��f��oH0��^�&����w1���`8���9�sM��k��J���/��i޺k�a�[��qIΈ#uU2�sT':r3��y�Fq���|F��x���r7��dG:���2a����w���î\x�nQ�� �'�Z�9�{���-���-�����o�F��bg]���\�L��#�w���>���<q����	�O��=$��S���s��DXS�ՙ��\��zaW�����ʉ�S�s�!��㰿g��o��܄����(����7)ːLƦ2�6d�+������ُ!��Q�T|3�y+~������	��x�w�#���aw��wq����G,���L�WTΜ�s6��Q���Rϗ��oUߘ�� �/��ߐc�d��1Y���6}��oY�~w|#��b�S%e�L�@�������_���jq{����q���J�Ty��݁z8؞���lzuWxd=��L�n�P�^��e��\5�����I�u�=���o
�C�x�;ն�=��3鯟�}�>TyH�*�&RU͆o�&���g�T�r����y@���l?%qF��xlm�~~Ι���쩼wn��*r�.}W�]j}�ts�&�zj^N�Q�}��*ލ:�\�nj���|9��̈́��4���ӽ9fl������ߥ�kBU�ip�qP�e6�Md��ۄ��S��k4}
�wGY�B_+7�] �_EZkt����Țr5��]�7j�=����r3��.P��}�uy�ߢG�;���ex\{!�fxoW�����m̼���k�u��vz��v��xx�yS���V[�������\*o��w�؉E�X.|����=�s�[�����q^~�UIz��0fUGn��
�aG��*�<�ϫ.���6�&��Y����U`9��{ -���.^'����j�П�%��u�9 ��+�E���y��?d����ݗ��)�;\�{G����N�.�#wHND3by�.椽�����]p�g��p�z�Z���~��9�	���im���G���1�p�g !q�NT��𾕀pުs��u9ړ�\S��Йўx�(E���V=�3΋�]���ur���BA{�o��[B{�@�e0�P��.�׻�Y�R/�{>���썪�Q�s�N����rx�>w,w.��#%iꗔ��q"\�p�^��r.�3��9�5�Teu+�G�6:v=�_�1큸G�[/n4S۽ű�ܽ�=�dq}a�; ���U�v�k뢄�IJ��s^�d91Z�>鎎W9=^�D���p���S��z��m����Q�7�o���6��Vʴ�[��(Fd#�W�&$e�F�l@{)�$���ӥĨOYꕤ��v�}�aC�D��t�AYw;�]�x^�'Csv��(m�X]BP��|Fsw��Ȫ����gf�J!�-vה���qn�{��Թ�Te��u.�d̟tE\9���@dh^��D|M���rϳ�����F��'Ԑ��EzI�pOMǽ��Nj��}"[���n�,T�,ի�^Pr������#�<��cK"��~ĆǽR�c~���ۻ���X{"e������"|�������e�Ϊ�`��.N��u?��اJ�ax"�C��v�H��U%����v��{�;��3���TT/^,V��t�R��!���{�c����F�m�U;�Mʫ9C�ǼM���2}��*��~����߀��j��s�w�v�rͰ��X���w�5;'�Vg�g�ǵ��}\x�񒀵�r2*�Gee�9��!f����z��ظ�>�`�|7݋ؽ�g�w�����~����l~���߼�s�n����tm�,B�^�W^<yESlz8&\uǼ̿O6�/�v�$g��E#CAt܈�r�R��}"�͍'F��l磍���k����uz�ͮ�l{_���S���>ۭ"7�d�����W��:����3R��ru�;��WQYy�h+ޖ��l�}�8^Ls�o[ }�V�Y��:��ں#�1��^�W;��Y��j��n,��N3�0�_���آ7���esg:��.Y[��V��G�&K=�;��q�;Dx��9�h�w�*n���g!�|�~ n����ȱ�i��*���ϳ�g�)n?�=��ʾ
An���k��P#c���E��C���l�pϨ{G��]�ۍ���6��2#�L����S`O�mO�!�qw��[�C$D�'!=�'c��B27f�ɾ�~����s��AX�@���1�޿A.�wg~@�dw������>��{uK���iI� �}A�U�p�j,�!��ޯ=�ǂ�	w7������!���c�M��=��.�[�YT�8u3J��ꫨ����n}3��nq]%�ϣ<�&�϶�Q�������?+���@~�I�-�a��F�q���ٷ^���k�6=�gz�NDH�������(ư�b~��o�Ь�����Pez��������$��8g�'�����M| BVlظ ���3M9DΥ|�����a�g�#�2�~US�6�6:b�d�BϪ*�-l߸h�}�+L֟t�몽j�<��ѳ��x����-��闟{�b���~��	��'�S��g��ظ�#����T�7}[�r�	�ZP�)�O�7��۪���ۢ,"1Qလ�Z*��v��z����{�!K`��*؜J��մ �-Q+돫eojJ���κ�������˧X5cT39��œ27:��������}��O��<�g��W�2���g� W��
�ro�>��1��Ϻ@\|pʨX��[�q��=c|.�p�e`�y�ϐuU?1�@_�x�ryd�B��ef��v���Kc�YFVF���G1G��
���.��{�[�~����~y��%�L{�f�H�<J⓬���m�eu�dmwh����s6V�c��\�';c��u��P���B�󗅏c�7��g�=y��x�����z����g��{˦}�ۗ;�B��~j�K�	�.�D����e���h_N|�k�e��b���o�F��Gs�/���z���^�e?z�c���Us�}%|�������7h!�9�j�O��;�����9xM�AU�[#��F�+�ӻ����#~�x#�g�	^|��{���:�i`-��U�*�mdl��S�/�~��琳j����,ٽ��y�7�����21^���t�iH����ӛ��Î�?|jf��52^]�f�Bw(�C#n��{֧��1ӽ��I�k�p�]_���%4�%��v]�a���t�vҳή�e^��R������heY���olJ�͓��j�/f�,Lɋ<f���p�YϺQ�����l���;�[{��
uv��3Mw_)ݶwD�;�g��Iܕ�m(���s7Xn���^�bbG;��N�|=��yN�b8��bH�+��h�Ҽ�WS�q���jf���5�c�nE��>�7����H=��gk�{=��`�1��-��[ȻV"�/ZѠ4=���J/�e��fIr�5�}59�y�C~~�R���7�ys/�H�:��ll%W<��U���^{K�w�� ?��&�E*k=�/u��Y3,Ǖ��T�N���!����[^�^���%;������>�H^�@z/�.<���V���ned?vL�~��/�{Փ5V����x������8])=���¦��]�v8S�ϑ���׻*2<��iQ�̃����/{ț\e���`{@��e�Y���I�c�t���s�J���j�k��/O�	ў�Gr��M��6�Dߥ�DV��{]�cB�>O@g�2~j�P��*�n>K�f|���ϽU^���W���ٹߗMl�C���M�P�v��>^�}sB'=�6��;h�^ht�]��g�.�d�cP���У����O��5��g�~�˿?~R����'L��؊���d���˄��)���ҭ�V)Q9�1����������cF8�:�w�����ռ���q���X��TPG�p=�E���K	V��yM��>�}��V�������T~�,�5Z1 u��wۂ���Gz����V�WE���:��0�}R�U�b��}'A.̶���V�
��	X�:
�c�娎�K1!D��VzT�����33'�emv�A��|'�M<�IAT#����@k���x^
[p��TӖ�Ȯ����ٗy;�V�G7^^B��-�g�Wj��d�&-n��.R�7&5xS�Os*T�n�_Ufp���(S[t�ޕ7en��b��{yQ��0/�3��Uf����;iιׁ��f���GI\��Z�6,u�u˥e���v3���w�/�#��e]dw!�Jǖ�f]�j� 3�mfh�][���K>x�ͫ��-�Ջ��sI��5�6�gw}�u�4��*f��)��N�k���f���0���u|"����o��e����@y�x������H{ܟ &kq��5�8���(a��n�՛ܼ�3k(���;��:�vd�|;恦���1�N�v�0R�7m"���om��܍>#����R$; �9,D�]�v��=�K�ʇ��i���{L.�t��tt8�Ͱy<��_txw��
LJ��kPc�)�W\j���ٸ��ux
Ӌ��Q0�mkM:wHܫ�iS�iL&nl��q��.�����C�ؾ*��A�.�X��ݽ�:�D�UЛ��]|�`����!P�"��H@q^ /
W@�w͋��.���B�MX
�ee����&]�;t��!��~:W�WWJ������1�D��Ԗ�!�xMqW[��"#�j+����{�0�V�t��(��d	��ԩ�����MP6�M�})��y�&�W��5�_a��[�W'\�;כ{��E�pEJb��AйM�ے�t&=�Ӑ���(ԣ�Pj�*7�Ǆ�m���2H�`�_y!JX���l�Gfqo�f"n��{6&LW���#`%'����y�e�;�e�He���Ț�q*���н�8,@���K�H����0��}�H��V@kI�Q�y��Dn����4O=��#�n��J�s�'q[��]=v*j ̸or����lWEY`��#c;o��͢�Y6�.X?��AH<���cc͝G�r�=�Q�wN|�Ă��N�����jVk�E�VB��<�s��}|p�]�+0�2Ѿ��,��=���
0D�����b��)Y*"T(*��$X��*$Y
��ZUYE�ETbZUcA�*�� �,Tb0H(`��m�QP�Q������E�Q��0Qm���Q`,���X����Ŕ@FA`"F"�Vִ(�#B�+UAX��"�)�YZ�eIP�
+UX��
6���,
(�B,"���k(�����
�J��mU�*�!TH�`�����E� ��EX2V�T� 1X��f�)3b,3QAdX�,UX�cQ`�6��,FKj�U-�B,Q���d��3Um�Y
¢ň�jd�u�T.��Ot�f��>��Oi�M�OzK�ӽ�BM���[���)q6�h�s�}8�X�ֻ[y�\�����Wz-r+����(����r������'�0���}~}�vXI�� �W>�vQn�%l���\��&�z+�d,��>�ھ6��Q�Jt�7W;�G'�FC�l;�tH���^P�!E�s�g|��W->�W]�@1�S�9G��mWxʽl�����U�{�5Pb��2�mxz��Gׁz��=�w|�xA�ت"⇘U�nf��7���۸.�������tâ���+�FO�QY�ހ�s�>�{j\���8éwV�>ȫ�6� ̏��tz�7s�s ���}�x��z�m���S�v<pOM����ꮰÉ���e��o��V�[�O�n^*�Uv{)5'�2�T|lG\4/Y� ��26LG�\��߬:�7�k�v��j��!��*�n��ĹZ0�S�idV|m����2�x:�"9�Z��.'�Q]��J�ϡ�dTT/\FZ�>=Ըv�s�z��z����Y��Y�&Ga��i�U�گ}�[2�϶+x��ˆso�E�]c�פ��s�X�k�ʎ�$n��W7$on�U����j�{�)��#'�̠-�6�*�~Pڝ�98�d&�+_d�k�ޱ�ic�l9�k�����	I�S�����-_Yt%5�ԝ�np��э�3%�ZʻF�:vYS.iu��AI��@[坘(]��VP���`T�xu>݇�d�x:6��V9{hl��x�����Bng���3p��jFEW��u�n�Y������ʵv;�;�o��zo���j����g�]]ϥ�'c�h�T��@������|#��X�{Ԕ~�ޥ��2\G\?Ow=;]ׄ���۰�'��dAs�6}���ד�u����㮼f��S�;����]}].}�F��M�^��� �U��0������;��)� �	a2A�;�(}g�=�U/ˆE��V��U����'}D�9��Ȓ��v�W����z��Y����'�c����/��(�l��yU9Έھt��&u�%e�%D�^����\�t	�$�ll�쾔��#>ݚHdPzȻ����mW0�˖&�܄��xo����){�1��w�x��������������JW	
���B�����nsc%����{�J�F���
�\/���нA�;޿J��zH[t�bd.�!�z��˿���.�8�[�{^������M�Q�Y�r�ϼ��<���~4$lx� {=~����%uٽ1���lH�72ۋ��+���;D��/�V�ϯy:�6i$���=Mv���5֟��/�:�k}Q�xs�Ƣ�����;Fq{Pi�f��Q����t;aی)�(��;��Zy�];K��c���9����&���3�0�X����S%��u5"G�Ϙ��n^|yb���،�ރ�����os��U<΢��ztb�p���T=8 4.J�ڱ ����xn���W�5�k"�Sߐ]��0|�Q>�>�z�u��By�v*n۬��**�-�{G ��ݍ9��[<�'u��ֽSގ\�ϧ�=n��G�)�t���d	��~���M�Ϫ�Y��Tfǽ�#k�8��W����z#��'bj���/����'ʦ}�u{3)�ng���"��z+[�7H�����Ŝ_{eNy��1�P���a������/m���S ��\'[���Z~�uϊ�Q�wI�g����dVS�����w��sª���֖��j��P��]u׼���2��������)ձ:���u�#����<�dW_��mwf�M���w�E�u��+=��hv�=�=��K$�z'�����x͍p\�p��Ȯ�{�m��9�|9���9�yh(�v��G�^���m�9�h��Y���)�����O���2����m׬����s�������Zz�k�'Gi�c_^�iY߰̈́��������WO�\���Y;]�]�a-�Z�LT�l�RS<����j�:��N����C�tr����X��\��%�iMU$����h�d��*Uy�tJ:�"�h�̸��1��L�!��o|}l�ZB)�IQK۪L��ڜ�viOdU9�k.�l3�s~��3q�x�
{�{2�;ѵ\�49^�dv���5�z3����t�� �WV��^���=2��
2���3_ay�ڤ�3�,u*�F#�,dw��	�z��7��}�M\���gY^�~��uL�WT�ynf�BlH/��K�{اڅy��Ȯ���Mj�\�[�=ʼF}O}��;A���pL��u5� � g������Gj�=2��W�~wEk���Ӱע����p�������q2� �yv�E��Z���Ū�p�������*��bB�>��Hl?u�����-��~�VCؑ>u`L�5���.i2VI�s8���퉨~	�qG�g=�=�d&��3>q�}7��	�mEfP��;����Nh�T*����Q��!�w�5O�#�q���3��eL�Z�z=T��]��t�<�I�K�>���*�YnNDo�K���¦�9�x�8����;�eG�O�9p�dҴ4�5�^4[�����d�r�v���ѥk�Gz�'Vݹ)Dk��W|��c x_�~�S<;�,�����z��uu�ޚq^�ݛ\���e��D���]i�y���g�� R� �r	ˋ��W���A�nv/
Xa��Z��+R�ӻ[C'�}�@Zu��� r����#k�h_:����/9ʿx�G$=��͕��*��ϚC<�~L~��m?ha�{NE�����`���~!z&}��93�����<��jEz♛��^zw�����S��.��T��뇠�z{�M*����_oY�X���n�g��=���G^L�v�u����N7��r!m�l������ff�~S�:s�}��5txzg�X]zJ>� �����BC�dVۇ�/�E�{8�ũ����dW�d�s����Uި���C�"sc��#!���@T��iR=�S�u��tw�G{VG��x�x���`������ig��H���Y��F�]��6@���;g�vO���3�h�_����pxBފ�.(yYv�j�3�PPd϶v}5��\y�_ϖ��)z#�kT��~Ν��c�g�m���n��:�u`t��E\9�8ئ����׹Y�aQ�^@z8r����n<�c���@|9x؞����P�(�J�ƕ�藭��r�@�E߲���s���qL��T������Me`,>��4����B�V|%�x�'�k�b|-����kM.��4��~��!��rG��^���}�c��,�G���Է���l+ �S���9�m���u�����V�1��7�7����~�PF�Ԍ�Mv�\4/Y�E�[�s=f��������u-�y|+v����z$L�� ˿���e�!����,idVE3��  9ڝ��o�Sw�nT��n݉���ʊ���@T[��ӣԸv�s�{�uG��3#q���y� �U��l����n�(6;+.���V����u�'���k9�6��j�rK�k�'2���?;�w>5�;���xnD���)����v�Z�����o�έX��o��·�G��Ӟ�8�i��]׆G��g�K����f؞�h��%�q0��
������dS�[n+�'�.�Y��2��������j�'Ơh�~��{�]h=xw=�o�(u��{y�.����+�����F�_VG>5[.g��y{���,<�ct���n�l_��Ij[~��ۭ���xE�pȱ�]����_��>�!���^ev���>�����{�Q3���n>H�a�Y������r�l��}��Hg=�]��L�o�r�2gD-�c�������>��5l�md�q6��s�l��!T�Q�̧�aKPd�i�n�A�(<e0:4��B����Rk�O���9������mn���SK^} ��xZ�A��K�j��h���vM�wd��s;�W�y{%�	��������7���#��٤������q�-ɻ޸J�ّl߄����r=L #���kv�x���x�g��r�➗����*��R�J_�͞�;��'ѳ>�Ő����ਜ਼���~�w���F?h�9U��j��Y�-�bw#*����y��@���Ya�կdN�:o%!�~���ϩ!���f�ES���GeFΌ3��x|��T}�����H����+.�h*D>ct9.1�3Y	���@mMغR�Ox��R�{��Ƈ���{���f%�10ڣA��h��xoJ��S�{Hy~$ay�w�5�D�>�g��츩�S�����"/te�"�-���aWt�kM����.��DӖ�IJ�����!k�t��wlT�;�Ȝ�S@�ET�"��Wu`�5~�]�W>�Fw��:}��f��/U�O�_����rW> s�����3�e�p�M$�Ng�{��>�d�9�b}y��=��0����p��V�������z
T�zhA��/Rz�*漏�+bx�Zzh��]��P����,M]�;���3��;��͒EN����⩜���1���;;�����n�+��2C���5�Bf� �u�-�Ud�x^��V�����>�*��DeezV�l���q��U�>�Kwa�o2�Q� \{�(�M����~��x���x=�fEyP��|���(y�^��6���#k��g:�"���8���XN-ϖ��N�.�=\r'�X�q�ϡ>��\��>G�r|�׮U��|%�xS`�
��7�@�nW4�2W��s8��9h�2X�j��&vu��-��A��߮��$�Cu�:˱.E��Tlz9T�<���;<`dk�F�D'fVB��j�~�z�X8?�k��LH�(^�?���_M�����ՙ@�F4zS��C�x��*��=��ǽ�{��R�qQ�	�^�����o���3�؀X�����7��j��ͪ,gZ������^�HHRf)v�����{���N�i7�#���ǰ�x����7�[�:��wmt����|�!��#Y���}����#��^#"��=�m�!l8�b��J˺��J�zbP�;�=��2�X�'��^r�V)���<r}p�u	������~��-���j.Ո�t�}(z�]n;��	�P:Y�/����]��<�=��it4ޥӟn�in�改�3�e�r��#^���j��zD���0�N��mn��lҽ�IM{Q(V�c���W+7��,�;���e����GH�b�i"y$��Zp����G���~�紐�4�i���H{����NG�=�w�W�É�*�
��C$1맳5�O'5:8��ep�oU͏+���=;�P�.
>Ȭ���xo�=�d-~Ι��۩f�u
���n¾�����F|F}P���bj��H~�e��W�#�W~���Fw?,��c���w�O���3�x�dvEe�;��e.<�xtK�&��&o����^Fy	�YmWw�mGoT�ҡ����k����!��[}��פ��:Ep�e[T;�\(�:!W���O�����4Z����ԃV�W>�6�D�33GF}AN��Ok�C����TH���$n�a@y��ʽ"�m����O�U1+���w5:_�,0F�W����7��4gј<��y������dA�s3p�^L�'\��@�aẔЭ���g��S�A�������fQc~Ŏ��������`�z˶ьku�mFG]ٹp77�y�+��zv3�m	��d�>�Z�j���S�7W;�ۑQ����p�ؓg��6odd(�d^�m�P1�&����!q��������|�l�b�Dl�,Jq����L�P�t쵘ȷsr�3g��j�4M�1$�<o)��.�ؼs�i:8��l�+�E���.��X)�^�#�q�뽮�ǋ?��p��������e�C>�u�S��|�ڮc@2�dN������ރ�s�ҭ�߾J�}��5�z�b��~8<!o�H] �"���(L�=2�]�/yp��*+̅�W���{*#��/����=�.v!WK�;)ؿ�2}��u��|�f�}���GO����x{����_�ǹ�_�6:�ԓ��gf���g��������U����.�&��L��E��n���4=���idVE?bC}�3]#4���������}|V/\Ϸ��$L���˴���:��h��S𿱥�X�����T#�����kn�y��=�Uw��,O�v&w�**��[��ӣԸv�s��=�;��6]�y��7��;��8�4=�ꭏ]lJ��ȫ��}A��Yp�m�����uM���z�_.��f�(��>����s��C�_���F����dO�"f���"�AȬ�El��,�wz#ރT����^���������OM�X-�UU��*���:��N:�bn<��>my����~��4+��}Α�����vSʆۃ� �l[j�5ºQ�N����^���3�Rh�R�"��N�Xj�:ݼo�������x��{i!nͧ6�G:�ÃD;X8D�K�Ց���^h�OyhD�;Q��ӠT!��$�1J������w��q��d(.ܢz�+�V�u�� �dW�U��/{;��|�&#��6_/���і{f!O�v� �FJ�-��>�Ȫ.������&e$#8p��o|��{ݱ�5u,��ndY����uHȡ.�G���`k��,��t%�)\�ɕ��i�УQ�I�{P;ݩ�uZ��T����a�HVD(������VJ�����W!M��g=y+zTX��Itt\�"������o�ͷ����$V�kq��qˏ�j�5vu�⨼*�42�����m�V�oD"e<ݬ���[7c
R.�n���[�[<��6����� y��n��Q8`��mݢ�u��s�о��KD����ř��������E�;�|��wRpv����::Ix�v�F_!�.�[��cl��J(;y�Z)\(����2aë�[m����]X��u�������}y��]��(�v�匛��"�b��qڮ���u�mv�F�I��}
7��o>YAA�����m�E[&8n!�S:/6�Z3�7��~��wTp3��gV��Neb4�u�f�U�V^����)�ߡsp�M'R�-e�b�*�D��*�.�'p���KS�z9�彠�O�kQK#�P�2s���3}[t�����\f���6��;.Xj<tY��6;2���;���1-�e��Q̚�)"f	�6�Y��wENƞ�H]<�j��s����X�6j�毹`<:���`�pg����w����f^k�R��Aq��"`���V�ꫧ3&��\�&Gi��k���G[z��ջߗX{��9>�,��Ǿ��ё"�,��EE�L�+��h�)�{��V�%�A����k�v"�}u�{s�F��ut���OS�\Vlܒ�T�X���!�[�F�t涑�;Q�#�P�x1�}p�
�ͮͅEVr�9��vN���s3t��% %K�y���&�qeY��Y�ˠ��)��h��duƯ��T�|u\��W]tN�t��#t��ᭃp���^o]�S�܌Vrݣ�j�e)p��N���!�ի�۲�d��**ұ*5`��n�9wwǷkzպR����W�
}r+V�gu���Wo�
n�n��nt���zX���*�u�&��s��˃��]M#1�꾝X��uM<�vl�k�81]`�'��_.���Y�M��v�w�Ϻ8�ԺC�G8�|�`�w��),����T�W��|i�-[eV�nV�����k�/(%���s�i��P���_Z<�Ԅ@e��fi	������{�(u.����w�_Ԏgu����w&�_��%g;�&얉\~8�ߜ���H�^q*�D�X,QUu!QAbZ,�DAH���&B:�X�
d�+cJ*ڌX*�,��+
ɐ�L�iKj#���M��s\�FH�A��AE�kXVUF�6ʔQMIF#,���ɭ��H��ŅIX�Y]mdY+TH��6�	P�R�*��P�R(�6�X��5**�`�FV�	�f,�XҌsU��֠�$U �`��������dYm�)�Y,Z°Ir6@β�dR)�ŋd��
�!�V1A����XMi,E���FAb�QaR���ь"��X!Z+$Y�.B�b�RE�j[b��6�ر�*;�7��9����ӫ�-� B��T��ے,�r�S,"
{�n�Ԃ;�Մ�W
=�6�]!��h[�����3���SjE��{�=�O���@�����}������𜎨�.�n�=�
�]^W«��)d��͐8g����WS�ȏV˼��Y��d�.�l{_���zf�O����V�� ��H�`�F�����Xg�V�𼥏��֞�k�xs�_�`�9�럽�f1x�	��E�\�29z�*�1ϲ��[5�2(=UNs�����j�ó�qU��>����γ�2׏e�gǭ�	|���l�~�S���B27f�A�"����x7~���d��}2`���TR�)�uQ��UǭX�Ϲ<do�� z�*N{ݎL�HS��G�o3빸��}4��C�S��W���F��y�p�3p�]{G���K���3��c���n`���1~�鴬����z�hأ2]g�=3m�N�QAf��##���^���2<h0����Nu�zz��kK���^}�Z+���2ؒ&J��@T��>g0�wT�M� ������aǃc&Ϫˮ9���VX�/ۏ!�xu����@lLL7�Չ��K�:��2aK6~���tѺ'V�wL>���[�2QW��WV�����k�9~�eg�.#&�{�d'Ν�۩As���ykqv�{}�&�lp��;��m���U����m�(���a�D@ڗtYۂ>��I�هn�As�gR��$t�����SK�'ǻ�}E��s��A�{�Ky�ب���
%��/(��H}��EUg�\��TI҅Slx�ݳJ}p��=;�y^xO������_�r*{�dN*hɗT}ջ#cK��3�=�5~����	ؚ����NC��ޯ<����2����½G�U�����-���z*���VK���bU㾡��z�!�\<k�X3�y�ϐ޹�ں�%�f?s6���o�m��u��S�FVS��[,�o_����
����	n�5���gΣ�F
�/s�'�[Q�j�{�YݏtOWh��?0�	�b��?�v�`٭�~�Y�꺟-�y��(q�Y�l$�ϛװ�cի"s�/^�Mg��W.A�h4;"+��m��7��{�����`����}M��.�y�2au��'ֈՙ8^⚜���ų]�#�G���1/�<�ב��M���Z=n��`�:��d�1�y�~f�yٗp}�eΟj|ߺvUׄzg�o����~���j�ϱ]�[Uޭ�Jay���<F�׼��+t�O���^�'|��$~�Ј�
�n�߉yc����IRg�ŐU�<̶���E��0���+:K��^j�]�Hn�nL��F�9|"��i�3���� �%vΰ·�*s}x6vCO~�n��|�b	�kq�J�h�(/S���]�oks`�&�lp�������t���\���vS~M�+ҭ.�V�����1�O<G���Yo}2J�W����C�s��E%q���L=Ꙥ'�nf��(N)�J])ro��U,�:��J�d琢�N�d�~��O}��:�u�;L��u5 $\�sȰ�h�sw���@g��|}�^�)3��3ފ<8�����{a̖*<�`4,-��rݭWѨدf/%R}�#��Z6 >v:�ǉ
���Hl?u�c�����˜���d5�P|�6��:��;uhYUsqz&Z�&��_�6�)ҿX� ��Ι��b)�ʟ�H��.�}mq�	�C�@M�S�P����txv�~�@z,��c����G��;��&'�{c�\�E{,m}׷2�ϲf�ׂ�24]9���2�
���_�����;�γ����:_�Kدj6=�\ҧ.|~~��πxP�+.޽�ck�hX���yUvl׷�K��|P��^Wҭz�!������^>,mԉ�񙢁��3�=����v�|ҥ�TT�Q� ˻����wO��ݶ�I�za�<gu >)Z4ț,�j�d�>�����l�%����A����}�������C7ǳ�c:��
����<��N�2�G.3d����x��k��ݱJ�G�Rߙ���J�d<�������QQެ��7�2 ӳ"��3=�Y���5m~"w�l���@���+��8o~NxQ�;tG��ל_��p�gѬ�<��/è��s3k���'\�\󮥣�N纞gf����G���<;����F�d,��,���{ՑEߤ�/_���֐��uJ����'�&��37��/B���f�[����جLο��ǐ�Tn�:�us����Yu��d�����{dz[@�lw�� ��24h	�[ �ۙ����#j���#�s����e�c�>�:�2^�~}����_�2)������|!g��T��C�*Ϣ���x��"�.䭉��yu��B�6�
�V�s�~Ξ�Ó��NS�R�Ut�����HwN�kY��Nf��w�Q�L��E\zo�0;��������c���g�~�� ٞ�~�g�̊�v��=��8lL󩞙*�*jVdx4=���,�֐^�J��0\��1틿E�f�/Y�>��g���G�v�=�2ؿ�@rڪ����Hr�o౥�]�=|��XK՗���	�dz�8�ton;������ܬ	�I���H�J�
ǫ(`a�+��� L��Ϙ�ٔ��������#��
b�m��cv�����6��� ��e�.�m-l��V��0�3���6��{���g_a�Q�Ժ��zV��?]�쾛�{v�L�B��h`�lςѻ���2/ֆ�M�:����������o����[�ٕ���x�� 2(4;"�ᝯ���9���G�R�����R�v&�;p��NB~��߇�ύ:3�N\L��R2��w�k�o��ɲ�U�^n�<�B�C��k�C����~���KF9ߛ��!3�1U>�D*�bV��3�%��ow"�t���|,g����r�:7��������@���'�������s��p7Vr������*���x�³=�u�!�nUzW����z�]�ݑ���gǩ��#����&������9�,��1l~�ɴϽ�\1 xez��W[��\����Sޠ�z�ۗ�b��<�o�_��؟ma!��
ՑYϲ����]�>��yU9΍���ϻ�ݧ�y��Xo�D�S��x�]O\�0'�a�Y��A_a�He�fy�}'0�x�%'д{�ܵ: ~ڨ>�굂;���Ǐ����_��S�Sӿ?jQ�ʻ$�g�Q�l,k�t�ӱuI#=|{�v��I��LE��-�=�F�V�b�4�Q���bT��yr�u�fPQ�EG�5��	W)Qp��v:`4^��&��Th��Cfrqfo�gc�8r���0��I߲��&N���r��(p ���sW9�p-%9r�x��	q�ͯ]��e�{#i0��xbX�����{��6��o�Jݱճ�c}��^��9^��?ܞ��s+ �)L�Oޔ!�=J���#ڇ������s���g}z�'�
�{�x����0]0�$L�,�+>���
�=N|�lu9D��S[�՛׎��|U�y5����,,w�诽��l>��t=9 4&&ֲ�ex,��+��VL���5Y�g��o�ӗq�X����;�u��~�<�ݻ7m�B���,(�s�;^�X[��^::<]]�Hs��!�U~	W����k� M}n�2$��D��[Aj�$��#�2���4	�G��TZ7�28?w�z-/�����w3�:�����m��ֶ�Y��03a�l��?u�)/��Pxl��G9��8=��;�����+��m{+=D �{�b�{=��g�{G�������1�[�NJ��g�������|�|Z[�K�~�A(P;�������UQ��*�~����u֏����E1ë������"6�o�r�Ⅲj�#�g�6��V��e �߆�1���Υ�$8&W�e,o�]�F`e�L�n��̜5�a=�\d�zVEck\.��(���n��[#V�O6]��%k�j��5�G|fl�gp�}˨�݆d�M�WT7�V�;���HR��gL��ϣ��z�Ȝ�����ɬO��F4x	hoW\=�~�.d�I��}y������9�*�jg��s+k�i���fNA{�js��ų]�]�2����e����kB�E�v��냪������q�l��e���*���,$��_�j��9��Rgp7�Uzt�s��Vd<���VF�Jc����~��k���t�kUj<�oN����uq�"=��K�
�������̜>�yT�FmQc:���s3�����IZ�|�����Bߨp_=W���an ���߀Mo��Gq{u�eQ#��y���9�+�Yx���!�����5z�FE=�G�U\�!�;�d�����0$��;��u��Y��=���.����~�5+�V��}�;�by����*��!�H��T(��mowmz�VW:��J�N�,���zᫌO[;�m�0�?m����YsZ�fm��������jxs��ޑ'�32�6���3~ѰC�?ɸ���ļ��fye��w�����L�[
�������k-1 F�����!���TB��^cV	y�5>A��JV�t�i�F�C[��i=�
ÝG���]��3y�w��َ�����>:_�=���I)R�zul��o��r���NIi��8�|{�~33ވ��Sx��	A��b�9�*�n�ߤ?�2�^�����{��7r��mZ�P��f�ZEP�J�Uǽ�3x��1"Ֆ�����2�
��]�wGMeOZ���j~]��G�wǲ�Օ���|�~w[>�6�^�P\�1Yp�}}��$m����j���v��Y��+�.�0dW���ҫ��y^���;��� �Չ�2���y�>�k��\g�v+ݾK%�ߺ�9�l�>�"�;q��Y��������ۙ59��C(n#���M�sw��煌�����z2#Y��o]������g�;�?1� ��+/��P�5�����9��֩��wu����y��~z�Z�q�~� ����~���<���H������`����Hb����v�m	�N�AȻS��j�=�Pc�Jt��Jl�������UY������R6��#�r��Ǻ��J b�l�T�w(�9���k��d�Q��u�.$z��F�]N�Q�^c�}�_�=����{�xA� �C�*R��}B��@|�8�{�5	�GRu2��G4>4��k�^�|I�6"z�T]�7���D�,髙R��;��̨���\�[���}6�<G�n�n��P�m��r�$|�z���e	A����@���^�j�XifV.IM��$d���V!3x8��ۨ>�U��Ɵ��aE�A��Ht���l���#̚bYٯ\xʬ;z]�Y^�u
�;i�>мo�pп���{X��;��(��=7��~s��=�Q@��{�w>$O�L��u�X��	Y�����c�Cc5+��~ć�h1�A�y���~{��^�7���Y�u��Lz��L�BbT�]͇^Cb\�b:���7�<,8��EV�ӺW�q^�Չ������C��v�Kڧbg��ʊ��V'b-����Wy��;xB���W�)��b\���Ϻ*��� yZ�V��fV?v�c� �����}�\�J���RY�*v=ޯv$9Ԫ�9O�~�K��;���xnD����jE���g1������M���}���Dx���B�8{���zn�nq��~u3���}=T&�w)]�\�&�J#�{$0=��VK���y������@���i��Z��	vq��g}�X�2	���ZS���뒷���G�Ŀ�>X�.}�X�ެ�q��UM�T��|/IZ(���6:�H=҆Pp�@:*��om�	�=Ȩ�,ޝ��t��锲�RP�kz�:���i݄�S��ћ��d�Q"b)���`��{]���YޥsB5���\&��ďo\&LܷP�&IϩP�*l�r/��|M�>ݎ�7p���b ���)�X�.U���Z����\�{���VE��*�^���9���O-�c�7]��z�)��D��w����T�#.<�1��̞��U8!�L��ys�z�_:|9C�2s�~�R{����I�P�x9���eF;�r�oZ���]��9ns��26�
�7�D��g�؎�?���N}KqOO�F��ǳ��/��Z՗�G�_�M��zR���L՟d<��*��p�2���w��l%9ձw���޾��w�r�랟z�c�YT�S4����f���&��(,ڹDe��l{�I,8I�7q����7�p߼=����Ӱk�!虖���.�j *D����w(���Y�SYk޿4��� ��5�z�ϡYcb<hp����y�^�Ĵ�µc۰����漲��J��Zq~�G�*lo*ٳ4�[����i�W������=���d-�C�qq%zvsrU��.z2��i���v�C����iձ�Yo}y�?��z�?�?�(��3���iZ���	2��"�$��EA}^	.H�".md�"�2�5%�'^$��yl��R�+� q�U�;P�B�X	!BЪ&���k�<�.�km(��̬��&ؤ���F�#(����_e��&a��y>sK��¤P�Ҳ�T��{�Hay����#�pJŊz�8[�d��"�I��s�]zx���@`<DD_�@�PDE���1	+C���Ey�	����=��bO��c��:��2�V�$���*����Q��";=f#@Kqh@]�d��`K$d��mH:�&{)t!���8�،cJ��v�9>���PDX�Ѫ�Rv���� & Qx���B���1X��2��Bm��4�w��yd�0�T��EAu�����4��y����{��H{{e�*}��\�7+���y�����;�x7�d���*�n�]R�py&�����>�.VOt/�h�Y\�u�>�E�;$E�r���vb�)�e�}~����
�"�z�c#�=F�&8�q�D�UӼ��GEQ�Q�EA}���}���LJ��5P<\L�fX}e�ʀ�"-���DD���B>f#�`��"�bF���|�)�RE�10JA�,�J!{���e2����@��Arh�ӿ!w� T+�u��`H����'���>��[�`|MF���rP�^��Yc�t�B7W�>��8��'�C�mJ|w�0
������7u���rG�L��/G�1H�Ae|��c���<̷f}�/^�ؚ����;���Ln-OW9*A��yio�ߞAk�"G�#�������Pn-�c��PD^���`ˬ0��"�O�LH;�	 ٓ��5=m!�&W���
�!�K٘m� @DE�X�`ڃ�<^�c��D^��qM�p���OL��Y�������:<�KM"�>$�۞�s����w$S�	
U���