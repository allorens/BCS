BZh91AY&SY��yߔpy����߰����  aQ��� 
�
      �         ��@�(( B�  R�         �*���(��R�� �$3ׁ4�o�R�ȥEE("$
A���ҥSù�ڏY��;�ħoROV������u�o{�'G��x/�^�ԺӀ���ۆ��P��uTq��8z=��t�����U�#���9�U�Nop�prw����� <  +�{۠(:T��0�}�� =]���d'uU\��;���n���bM�8��V�Ie�  ��͕&@gsҒ�
�.v���=�nڎ�\�zW������ب� ]�J�Vތ�U��J���n�����R���K�q�N�T����/oo��a������%��.�`5�pPޞY<��+*ѻgx��y�9w��۵�U���i�T�z3�tznkw�����I@\�l�@�[ I���y�����{۶3�Eǽn�����5�rw[���)�oVӧ��L˛�צ{�y9y��vvw���yu\�.��7"�^�9G�%�R@�j�&jh2B��*J<��ۊ�u�vo�z�O*�̇��'z�oz���G�۞d$E��ngu�m.w�/=�=qt�޺�/{�'ht�-�^���kͻMswk_:                       Q���4�%O@5IRI��Fi��L@a2i�����iH��Th��0 &M0&�@�Ȥ�Eښhhdd�� #M&�JT�i�d���M2h  �SU�4h� L�hj��<����x��H
�y&��R��&����#@���'��TO�Y�vo�^��<���(���^z���z�wǾ{��i����W�G�x<͇sv���8�������ula��1��{�?�Y�f�����c��o��Ms8:8_�v��P?�F�6f�ۘ�����.*�?���fl:�����nr���3��c�c�ߗ�{�������۷W�����?�qE��g���P��4��J�1t�gO�c8��t��$c��h�ɐ1��8���5DgBfX�����J8����o@�ʤ�X�3k���f1��1!�1�e�cC,E0c�1�1�p�J1�c4�3K�2)3��Ԙ�,c�4cLь��2�c��b=�K�欁�d��g�c"1��1�p�1�f�Zd�Y�1�fBc1��#�1�c$~gc2��X��2�b!���ѝI�@�1� clg��P�31��X1�1�c	�KHc�I�cFJc�%�21�c�`���1�c4m2	�c��c$��g�BzB=����S�V��|����C��L����E��c8���p�d�?T�dc0�X�1��1�3F1�gH�"��1�/1�1��222��4G���qh�x���Ey�#� c)�1���8�1�c%��F3Kј"�0R22�dc�G����fe�3�h�1C�,e3F1�Q���fz�g1`�1��1�2 d��1������!�E����a���f�k2�1�G3�)y�օDE�#N|�e
��1�c3���Lc�1p�1���P��h�1��1�c+1��X!���-Ld�c"�3�P�1�Q����$?1�cظd2���1�|#2�e��1�p�c�3��Ȅ�1�c1�q,c�a�!c#��F�c�;2J!���2����e��e�1�c$vi�%�!�c�1�`�ь��Lc�?3�1��7-��)#��:��"�!�3911��X1�$��1�eZgC,����1�2df���%ƌd���2���H���32��3amA,c7F2F11���cǦ�1��1����c����,c�=�1�I�d�b��c�c@ʄ�`�3<��)���c7�!�c�0d�1��1�gy�@��c4f�?P�W��^&3FX�%�c�;�2�@Ȅ�1�bќ1����@�I�t1��SVV�#4�K��Q2d�=kg�H�&PO$AF����>\O&�
"�@�c��!�c$i1�1�L�2Gɟ�#͕D�#����8c�1�c0^��d�cC�)�2�c5�1��e2G	�cظc(c��1�1���1�c�d&1���>Ld�Y���˱�~e��E��e�1�0c�$c�1�0����a���Q#�`�P�1�fC�#'F2SHc�:Lc�i����s��I����=^�UM$"i1�N��,|���F�8c3�(D����,���5g�"�1��A��ĝ�@1��2�H�{0��~���D&2iX��-1�ˎfNr�-+�I�c��$C��1��4�1�c���&!��3�����\!�j-Ie�0e��P���c$�Le�f f
Fh�w����%�d~���maP�&@�L�9\12�`�����I�f�	�e0�)��R�����1���Q��1�c�g�2
��1���d��d��w�G�T��1�SHю��2AИ�:�V1����0r�c�h�2�P�<L��Ր�Lc$|�i��,�|h��`�392rL��Lc�-�1�S�̈́�ሡ�~f�cؘ�2�ic�g1�eRc�Y�p�#�c$c�Lc�^&1�P�c�2��2�1Rf��HńG؋DGuQH�����q�c��T�m��5Q�iH�"L�P�3�ь`Ǌ3`ƕ�!��1�t��1���1�c$c&1�3Y0���c�Ac�cε�� bc��5c�21�-��1���&H�ь��Fc&1�f4�1�z���C�2�ɒH1�;Lcg?.�1ڡ�c0r���Y#ip�X�&q�p�3�1rf�1�Ԙ��D,�1�Ɍ�F2!1�c��8��R��@�c�@�4c#S#Δ� c�Čf�c8��&��P�3123UR�H��qZ��I�z���5d�1��@��C�Q�;L��c,c0�X`���f���(�2�eJe`�{F!�8V@�;Hc4f�S4��J� z�c,��"�1���E� �4|�� �����1��d�ey�cc�1��LcE��2�1���8^c.F1��0�X�i�c,E4�.����-,eB+a�����ؤ�"��c�l���V1z�#3�7�G���+���� a,�Ke�c%�c(�(�q!�x�c��@�1���d1�1�4��s8��)�jF3��1p�,��h�΅��Fg.'����(�ie���C;�c$ᥤ���ec0eI�	��)�2�P6��.�c���$���i4@��,C��2j�$$~c c��q^i�	�I���XYd��-(c2��3	,~cX��W��1�e�����	I����c4L�m&`�>LeZ,�Lc8|��^Fd�ǋ��+�0c��2�C�0cɐ1��2l�r��FcRi#Й�?rd�2R�y!�f�cc�U&1�e���d!��1������c/�(�1�c�4�2N�@��3Hc��L�F1�)�2D1��1�e�8be���/!�c%�c�ב��c�Y���+��31�e��� ����@��h�2-�L������I�C�N4���=�3�h�$��LLfc:�q"#(c�/���)���d�b��6��p�L�1�e9Z1�`�2FH���q���?2�1�1��L#�K�1�2�[�a`�1���c5�2F2�c��7ȡc+�c�0�P�@�Q����q1�3X�aƜS&�D�32X�!�Y̢�(�2L��c�уD��_�c�9�fI,ќp�9�M��a��~�%�D�2�(��`�5�s4��Y��2��c8b�b�,���4�4f���(�S	2��έ�$e3
f��̒E�'���Fa���u���g���C�f&i��8�2�o�f�ԭ�Y�㰡��4���𡌫H��+Lg�f�H��`�1�H�Gf����f������9��a$�e�I����"գ��,gqi`�$b���h��p��f��,e�(������!�Xʢ
c(mY�h��h�t�Q$bI/2D0x��=T3,���!���5�3�)H�1�#��$ư�;L���4���1�U�ey� `�	�1�渒LP�C�3�;�I�0�X�i#s�0ɐ���Jnj{�v���?��~�3�2h�!%����,��>S7���aNg��e:�ٸ�)基����?�ޞ�J+k7��>���d*�Mb��mf������ �������c��>\����}��;f^w��~������]V�e����;�>�}/�~���_l��Y}�O�����\��d�n�f�n��%�B�mE�i��Q�ϺZ�93�FL��Tە���Wn�ԵOz������W��Y}7����T�}�ҵc�x��Neٛ�V5**e�jm-մ���l&)�S�p�UG�m^L+ĦҎWU����P�rkRɩΔ�HZ�ޯ��^؏��5�li��Yg�<��ʃ���8ڭ���-�ߩ��^�f�D�"��yV��ʼ�Ne]<��bي��Jˋ��4��\vE��UO>RL+���/���Q;+o3yG=sܦk��)ǳU=�����1Z�̫NN(�{rF��w�d*�OTT��mWL�_�zWz��?%3]���{&gn�䉧�ndDƛB��g������Ư�����z��n�Vvz�Dfݙjft��X�-5i,A�T�}��M�D��5�dD�uL�DM~�S���w&be�����J���3Y��ɳ}�<�-����՝�]5s2��Ew49��D�NV~��Y�\nM\�I��}����߻��o��:��O�y�Q~܍���)�:����s9��"�U�_���[z� ��v��!$����}W�}q��W�-��͝s35?E�Og�*ښ��R�vg앫n���a�jәܹ\�/&�Y�nTZQ�ʊK:訣!R��uy.i�]�7�EKY�C;6{v�������_VU䢩gg���5h���Q�B���s��SKelej�N�gu��ޞ��Х`�-_3:�O׿-��fK�Y�\���V�hZ�ft�ʅ�SJ��f�yF��W�:�Q�˲���qQQ)��k��SVʈ�i_]�y�\uLʪ�u�og��U�%���wK����V\BP��]*�az�v�R���P�ނ��l��m�O�{�o���5$�a
rR��o�����'被�	��K�����]-�*�OӅ�WHRʓ����t�v��%��ܫ����N�e$�/�kgk�ws�8.�T�H:�2o������z���4/��cƾ_��}��ڋ[�,����'7w5�*���=1빥�u����WyO�u����v�����:�.�y˪ƑP�)*K؝u좷�^��C�En}Y{�j��A��M�(P�P<=�O�<�<:޸�����$U�)�ԫ�fl��}[x�ylT�˞�jpˍ�X�=�9R��̭��rqz{��;e��o�R�/�-��2o�͟C)�sE�~����q_K�/=;0���+�u�S9���sI%�;'�*n*6~Mٱ��Ү����2 ��qDbR������ ̵�{}j�Z߳y�^˨UTk��z�SN��I�Cȵ]*r��w2M2�q]ђ��u�Vb���F�I;f���+^��ԧ�{x��*vHFQ}u���e+Y��d�k�7�[��D9-R������Q=�j�WD�f��г*�y�3�V�Sa+��IBKg�^���ɛ9�_��yl�u�rR�)㮼�\���W)W*�צcg/���ޔ�,��z��b�UJĵR��6{Q��I�:끫Rtr�ɹsr�d��-C�mMz�%���ͺ�^�T�*��TeD����Q�B���+I%tҵ�k%TJ��;Ϋ=YM.�i+FjsjP8Qn�SU�EUAѵ+������^�M�D�!O�*¼�*�'��;���;{��vN�6Nʤ��j�	؛���Ũ���D�Z������8��=�)R��D�V��ZfmE�Z��K���y���V7�m��� X�)̳,��TZ�5ҡ(�d�����*���y
�t�<z�;Q����]�L��j���޵���w���Jȸ"�\������ʛɮ]���mX���Q1���nb�K��u���͜�j�Vmm��K��'�o.�)�
�/jY��¬ɻ/HU�O�VV���""��Z���J�*�M�9+�6A��L��)߷gkjg5e���K6�z.�ZڟMn�\㦖j��dtTN(뼥9�\[���V��əw=w��ؼ�ڊΝ�aBq�8��m+���:�����\-���"'&Q��R�ߩ�����"j��a�~��ʷ�e:pK���Qm�Fbř7��d-����U�I��װ���r���yUSj󯯔,Aݴ��9�~=��y��ǵ��þ}_1�/*meU]�Ԅ,�߮��el򭤷_ʊ͋E��k.�Va�؇\����Mu��][.�qE�C����BqN�%J�/λ�Oa訕�BP�}Y0�jSsWsK����s��N�X�S����j���V,��͛鬩��vq��Jo.g�]�(���E��i*UTX;�҇oo;X�6������ħ;6�Hh&�8"z����
ե��)꽖��>��UA+2�r[�Zfr6�eU�K��W]���p���UN�wi1_D^�\�S{��YN�M��J�\��J'��l�%WQ����ruK��&Vm�팸��UCr���$�E�VU*�T��l���\�C�"�:kT]�5�*�UbX˥3J�4�=]w�v\����ݔ������f2�5uY��n�z�/���vRX�*_|�R�8�Y�[�%�l�FE��,�+�ʲ��=�Z��"Vl�T�NF�j��(���N�ҙ=
;qns�h�s*'�B���-\�?fOe.��_]}jT��Ϻ�TU��rS�*WЖ���yYi;���."ra�[�3�ݓ�S�J�;s�z͋3I�qU3=��ԮEP�q���).籛-	�,΅Y3�5�M���3[ڷg��ws��KfaGWv���E���)ކ�S�0T�w�h1�'�}�.���ɩ鎙s}9��P�jZ��J����y˞��K�)��-��������Y����n+&q����vfZ����Om�]ӗv�b�ɕ
z�,�i(=7Sʣ
Ջqʌ��5��{w3h�D*�ʫ��Au�S��zk{���ck��Y5y��!ud�s�2��R�2�unoL����ml�"�FvvK�鎺�5n̬ɹ�į���w-B����!(����;'UBnf������У��#��~?���������ރ��R�+�]Ḑ�6��O��=31V���Ǝ�-���}�Z�{-��}9������q�7��$���a��nF�1sK$뫋y)J��q>����*�u׮�;s�f1����ѩ��I녴��u����H�ٻ"�fr�^_+�#aDyMҜ���.W4�u5�]I�E)�-*xO+���"�U�jS�&;�e�}��z���K�Z�u����ʿw	}ImlU��n;��IGo׷���Uv���:�_�߮K�"�W)ʍɒ����U1	D̓
�����%��VT��\}a��#�*=��?/�}Ss�-�k�J�zUe~W�izr&5:�JqF��T�ד�_V̽��Q�͌�yn�dm�Mɕ�Ҝ���j���v�\���6s0��Vz�al�� ����j76�Q}�Bu�Z�A1�wB��H���J*�k睫��>�B_F-�2�����W�MC޼z��5l�̣�"��Q|��i+�3�R�6ֲ䭓z�ol�関b��T��p̺�"��t-�Fi{Y�fU��x��%��~L�3N����V�[R��*�sE�U���W�T�Ծ]�|�|��]#��/!]�	b�6;bڼۊ�b��Ԫo��W�5�5�/���kU��+!z>�ǳQ�j�؋޾���y�Ѵ��U�2I�ٝyS1�-؞�t����nP�g'��^���$O׊�*kmC���)��+Ϻ�ov�q^L��v�u�V�N���vKͰ����f���V��{iE�?�ZU�k���Т~�Ι3!}ҫ{.�ҕ��
.�c&nf�\�|��6�-�~m�c_<>��oy,�n�?�;e��d��p��"��*K)n�5����.���M+/���6��H�Nˉ��X���1���~�_9�-F�[�Q���&��yT�u�n���.�^_<�MV�i�;s3Ң)�t��O*U�d��wv2w���o�LwH�J�%9���RO�\��b���z�'r+��&t�R�>܄�߳��{� ��?闫<���͞���-̪�܆����ͼə����+�y/|��K��χ��M_���-x��:�)�K�'elM��L=�hO��������?�^�u꼽��8㿽ٓ���^�s�w}~G>e1?����_֚��^���˹�[��q�&���Ԅ��B�38�����Xx���=��K���学��+�R�-ɳtgC�ǰ��M��gі�j��,إ��i�]��5���1y�#f��ߞ���m���1M�F�4n�e�H����l�!���*cX�NU�0k�ܻcʂ��-�����p-Z6:^ڸ.3�+�M�=������Ϋ��,Ae.�	z�E[�u��包ι���s��ñ,Ɩ��V��ФM�Xj�B��o��o0K3�����_]��4��-5�uGh��o���kj�g�`)�!Yh�a&"�~� ��_5&ajt!uY�4���Ҥ�M5]�/��nm�X��e�n�\�����Ǽ�e`k"vZ�+3%�h�iV`�-�!��z��u^Xa�����4�T���栀���(X;d�Y��]�k��T��Y,&v�,RAs	e`���[�ÉLSo.�3Mbr$�X#�Z^u�b�4c`�Uԣ�P�����Fŉn*��3,å��2��f2Le�-Wq��w�p��M
���a5R�\�M.��?.��{���<���r�cYxk`JIP��.t�1�����ʋ`�
]��qf�*���]-t�g]4A(��	:RQ����86������X2�R�\Z�؍�0��yE�8ԃN&�N�2g��B��{�����Z�1���et��1ITHZ��`�b��F[��Xj�ԪS^u�ғ:29#(��3��6l'��?�<!<	�ų\iXQа�*�>�蛏)*g4֒�5�LJBj퉖 ��0+��xr����ҏ����d�?���>6y,ܱ�l����5,�i\�KMl�Dfm���cU�x�^ݨ��6bKy��9i�d �\�k=��%�~e3RK3*F1�� {{r�f�9��FZ���[��{�H:�Y766�K�EӬ4v�,�&.���2�iuŒ�h���):8�.�0K6�N/;f�ˀ��Kʉ�tL�F�w�����f%�������GT��8^�&�w�=�$�=�ƶ��c$�<,���D��BP8�ffa�.�6�Yl��G5�
�v�F$,��jRRo^��/�걸�Т-��f����f��U%��!+ȷ[���bd���x��)6�Dc
sq�����"XI��@��fؕ��<a���#d��9��t{Q�p�B�cm�r�;0:�n�ZW�����6i���(�[�V�1!6��悁��f�$ŕ���mS��v���x,��:�j2
m%��0���0�[��>Z���ys��̝�W��jÁ�k$RPv��S����1H����fD�`w�x��H�&<D���fH��G�|t�:���́�D� eNn��L��N��z�5n8]�?C߈����r9���m�3l�///'�ϗVf�������ޮ������{��3�$*I��&$*�+fa VHBL
65mͶ��=��7��wſ��������ܶۦ�vۆ�m�m��cm�޷��m��6۶�6�o[M��|��m��M��|��m���m�m�n:e�m�m�m�m�޶��{T��[m�m�m�m���m��m��|�q>�K�< �{���͕��͜��,�cjl(�&n-�[g8%Lm[c����Fqb��m����/��y�6�m���m�nm�m�m�m�����6�m�i��xۖ�n�n�m�m��m�m�m�M������m��i�����ܶ�v�t�m�m�US��m���m��-��ݶ��z�rx�L{ށxFBIm����Bx�!������#ǡ�yX���ܶ�xۆ�m�m��4�m�m�m�m�m�m�޶�m�����o�m�����m�M���ܶ�vۇM��[n�ۈ��m���6�m���m��UUSnm��m��m����ܶۧ���}���$��(H`���A"Ņd�+�협Il,I�q�2R��1(�ɉ�����͜M-�[K+	5	5j)���ՁdY)��b�YS�)\ۻ�>~~��3a�Q���������������>#��<]^���1c0c�2�1����#��n8�i�i"#����"=DGq�ϛ|�G�c�1�c$c$c�3F1��Di����]DCI�1�c�1gD����8��z�HB��33F1�1�cc�P�1�I$�c8bc�P�1���Q�ֈ�Z�B"�|�=R#h�-�Dm�B"�=Z=DG�����H��DG��)�]u��]G�DC$c0c&b#c�8ѝuG^�q�>6�!#kDz��B3�����y����ԭ(ղ��hY���fW����m�e�LKs����F�FXl�t����[(5/z��t�Y���۝4Xbhnn���*l�ٌ6tpql	�3m�p��Kq5�����l��cj�C�fv���Z8�.؛���A�]��E�69,�Ri[2���MT���0��
sp�l�

F4ٱ�ʡ�o���2^�u��l.�-����ErM��Y@��)q�YkLȲ�kH$�":��f�L˒�Y���+�E�h���,�ѵf>o�-���[���Ue�fg�3t�P��l�Q	r������6$x��nvlk13�SS�k-��y�Λy�cL��Vט.l�uB����˾��<�r5��H۠�\Vc7�}���Y�j�5
��CF���̶USW@̫��!%��lf�H�[*��5l6k3In�;Fr�X�Zm4����V����e� �\h�VR�{L"d��ر��KK���eJ'$a�K�����IHն�0Щ��Ͱ���ʔXN���,@[�%�;ܝM�ՙ&�B7)6A��y��䘚ܣ��ZP�� �p,�yX$�jXc���M�>Ku�z�X�>}(��n���%���z�f�+�����eZ�ڠ�t+y̰��������1�}�Ƞg3d`U���&kr��~\��̢���*��]��Kf�(�i�f%�a�-#�4�Bi�fkje�e�c)�3p[1-e�0+jc�l��'��cf6���s3-��t��k	�Dt%�R[6�Z���v��	f�������f�s~���Ux���ͦ/��n��l4V�\ڣ��k�l�'�6\�;#+�g�hd�]B���O�����f�t�*kL1ֲ�7S[��n�;CE� ��Z;gJ�%�%dm�6�|c�ZKhw�����ݙWRGG�i�k*�P�c:%��Vi���*��U��䚬2J����h��b�{Jͣi%����]v�53I���5�ɰDl�e�lј�ݗ���s7�ٜ͜��3L��	$���~o��m��wS���=�����}�����m���ٽ�x��39�Y�I$�{����<|�c1q���c8c��,�I(����|j���weu�ܑ��ix	���5ce�1��`��km�iX4L;Tz�WJ��x{)���\�fl��M����:�N�Ż
F1B�e	�/�ұdׂ�R�Uu� �
8��k��g��;�'.U�M+���h�7#���r�.66��c`�R�ut[n�h�ܥ��kWQ��1o.�\��� �3���J���FZ�!8VK,,[H��c�5H�ږ������D�ӷ���1�	 �w�-��a0�����h�;��%nW/���^���t����=�����e�'g�>���hxa��50��rbd�O��3�ABZUqf���I��ʉ�ix�E*Z�V�ffΙ�������z~��Oo~��Jj:�r��a���o�
'�)���8���u�|��"#Fa �(��/z��N����A��
Q��I���5��\�w[K)�^�3�� a>XI����#=w40=SSb
��R1b���AL�|�I�N�[y�|�Q;(h�����`l׃��m>v0�����cz�I�]K�\����U�rXp�A�4h�Ѳ}�Q$Ae{PB%�P���X�)J����"Aa�3�i��G]GȎ�"8��SoZz�����$d�C�N�
 H�ٿ0�%.Q���ȑ�ό�rXj(�a�R�QHX]3�{{�"M=0��A�Vl�O|����R�\l���=��2��{��~M��,5��A0��F�%��T�3�ðá��qi��\�44;$���ϗ*D������ߗ��6&�p��o��f*&äJ2�c�/�y��|���8��0c8c��,�J3�eA1⎺����èZ�{�C�ޞ�JPf���E�+���=�J��A{���l��+(J�s$�YAfcc�Be4�7XJ��9�4'd�q�_��A�hٌ���v�>�p�98g�ĭ>��s�_>-�����2���O<��4�gٻ��y)I���O<�3$��uX�x+xl��9C�[[�/t�0��<5|�g��8�|���]GȎ���O��d'f��{}�n6"f��VaM����0Ʒx��>��+1hݦ3��-*��l�t�&ߚ{w�١�+o��fuc^�+G]�Sd�r[q���"��dK|�;��%�H�ˬ]v�'����V�4Ѳ�F�6������y��m1%󯧹Rl�����%�z�fO�}?Sp����E�y�
�+�7P��X��tXP�ZU/p�ԗ>j��������o�(�PIg�0��g�����R۳rB�lC���i��	z���v|aТSL>*��PL�(gܕ�����|Q~gN6}K��o?kN��.|��0�z�!1��`�g&��r|]��>�D��դQc<l%�8�L�4��c�Q�#��#��e6������¬V�Z��b�jjn#KoX��CR@��}UB���ey�Qg��SI|W�=��$^�J	�y��_���i��|�=���~|�G�SQs3=r7��^��`�z\!�!���>r�0U��E<:�XQ�'�/=f��y�7�k�Ze%e��e�6l�0gv��#>��&�~�%
�7�~D�͂�>����Fϧ�X����|g>F	��FR��Q<O��/n%$�Y��f�|���]GȎ���#��֍An�iU')>�_΃Ҝ9!��6�Jj�BN�W�
	���d�x�������͘Ht���w��44�|?A�!t��=1`+�&vd15���e��[1ښ)���E��q>���e��c,`S�~���ɸ%Ӕ֊B�O�5��W��>)��oL���Sp�𧆧�­����z���ڪ�ըӈ�8�8��DGV�>DuDq,�޴���خ8�gUPN�\�y����\�v��(�mi�"+�gO��vY�d�>��������{�����q�t~<)O0��&���aL�a�y�7��D=eQ�0!�3�p��$ �F��g���.��!ީ2�Q��J�f�.&f��x����e���6
E����<6l��+�b�Pf�������$DI��A'���x�#t�Ē��}�p@�q��|�Dun��GQ�L8�Q%�Ib)_\�r�!S���/����xd{m�Kh{u��,�D��M4��1��ˇ��4:�!�\ۡJ�[�p��4S�ї�}�s�a���%e�| I�h�Ʋ�yƶ[af额i�$˴�I�fqx�3�ٝvW�(nK	)�J l��O�MO��!!�;3���^j�3>��'�G����=)�	�����\q>�m��͔6oF�8�(jG�܉�;���G4�+l0�y��94}�m�����ϔ����[My�:����5��۳�F�ġ� 	M��ӈ���yo�նOQ�t�e�n�̦M꨾�9Ao#6y��:�ڷ�?R�6�d�I<�,14;	��O�n&�i?#���g���4����>b":�Q�#�㯝me=h�G���xjblf�3J�"'�|>C!��|�0<���os3&�?`�����s舐�=�>�ї�Ek�n�8��WX�n������!�O�I�K��aD��Q�]�(RWܖ�Yޚ0��4��,�F>������Lyꝷ1�7n:��j�ܱ�K�5��J3���)!���͞���:I'4y5��Ke���3J,����`�;`��^��� ���0�df��sˤ��.�4S�x5�nm\$�o�e���<)|ձ�|�b���^1x�xˬ[�b��5�n�x��F/m/*��Ɨ�m�V8ƭ���0թ�^1����W�u�����y���V1x���^+�f�������~W�u_��Ǭk�b��׌^*��b�N+꺬T"ݪ����/H�F]b��R������������˪�)��aX�c�_��������~^���οj�}W�X�b�X��k�U��F��/�c�^1K��k�׌^"�������Ɨ�4�ұTˬZ|^c���ϋ���K�&�+�V4�+�aO�]1t�V*�x�+m/����/�.1}U��|����1x����1��cJc�1x�G���z�����5�:Ǹ��S�b�b�_1x�+}S�F/ϔ�[juZU��mX�S�1�b�^�o��+-��|����n�Xs���R���a��}����O	[)&�Y���Ж�ï�L�ׯ�N]D�U!��4�ll$�ir���Tb]�̛RT�VB���=Tryy,������J" ��"	ʩ�ቃ�4+��y�O��!�y�^ץ�;�[�p���}����>^Xǩ���n���əC�X�y��(\���]:�䈤DJP�_�/g�����[��33��_�33��&g�k���<�33�̼���'{�Ͼ���+����e�fI��3��������"8��"1��1�1㯝m�4[m��U۾�ٙ����[J#$��� �Hhd0I�!�$����eKJ��\��<,�)�Рq�H���~\4h��I��� RM	��`4O�^nL��ĝN�k��˚�5,��N������8!D��� X�I``4?	�Y4$v���	��~�f=���dd�O�'ߪx�nӳ�0w!]d�5��se�Z�m4���I�<^=��<(�UgZ�W秞�i8h�M�-�u����Sr�l���f�͖D���ۢ,�i����.�՘�o��L4L��8Q<�YNx4��ծI>'��n0�� ���b �=�l�|0��ON�>J00N$�u!��vVۣrw����[o$�c�.�١�-~y�kǋQO<�G�?1��~q�κ�i�Du8�[G�-��6l��m��W���͙lT6k	5��ᘌ�'�T׍�rh���fz: x2�$�d������D�I���d"p��%H�ߟ�~���y�\�65Z
O��%��(�R��-�3&�y	D��ٛ�C��'|8$FI�_)ADd��q�6S�"��(,�Bs��i|WE���a&��M�$1
$�2���&��۶B���)�f�s��Gmр�F��`p�a'��x[�F�u��:#�1��l��F��PГ,EO��gI	�d)��4G69M�9�Lض����2$�,�`�#!�K�$�8�����?9X����	�d���L|R����=P�O?��_��ڕ^zz���~q�����c�b1�|�h�E��M���y����n��O:����~"��y����Y�;������;r�o:�7�|Y����vI�����R����||z��W�~�ě�{{�g���Yl�����D�n+�Obo16�h��h~�tH��=<�j�5���o������� ��)�J�B�����;J�0�gc2��a�����4j�\A�{�ՁAѲ��N��S��M�JI���E ���ὅ�*Y���:t����:!���""���P�! p�fP��LG-���$�y&����$���%�g���ten'����h���&��r��<1�Cex$Y
 `��Y&�В�0�)Z���xp���!�;�ќs��xgd�C�C�d��4���h,�Ϸn�(��d��[K�D�$��rC��l=�a`|zX�I}��f~�<C!��0ub�ȡE	��U���kWz6;�����a�_wi�=V����p��΍'����:'FHlԢ��f�
i��D�妑����؇�SΩ�c��?8�DG]i�q�F8���y��m���~���-c��"��'�2C��0=�������!� VB~�)�-Wb������4R��N%�`��;���ɨ�gg�WK�tl�vC���vLJXS�H0��O�b�����$8$����h؁с��D��#�mԛV��ç'���f��O�~��0ɹd��B��>�<��$��S)�Nmh~O�ܜ(tB ~�߾䩻��I��Jt�X���:>��<P����%{�z����j]M��;��a=r���!�$���$�P�ϗ
0���.Jt�d7JA����n<��xd��Rȇ�4���t�4&�;�i��'R���<����%��Ϟ����v��2;7��I @� ��ksP����V�b�漿(���˳�����q�"#���q�F8���M)jl�M�=���K����(�03�� 0a��ӥ���G�[m�;4x$���P=��	8e�蛄����c���$Cg_ʗ�
Ӈi@F4Rq�l����ƶ�Nt�%��!��h��)�I�I���,�����`�6u�3
�[��Nޘ�r��p����r}��ύ�`��d=}B �a�5&��84��	�0Cާ��	F&ğx44CBD��L�ٰ�M��z�82lB���Wz_����:P�>��&q6τ��4$f��0` �d�L�N-��0ѹ�j�{ϭ���Q(`$�C���!�F�8��n(�+��P������8��":�H��c��6�)M�)�n՞n�iʼΦ���@S&�E��/,6�,A'ђ��q�������{������nȷM����m�vDFxf�Kp,C�<�>w��I�s��j|"	=��l�f���%˒i-G5t�7bh��m٣���w89l�Q�c�ܣ�3�ChhC�G�$V����]�.k�q�r���	A�b$�ɂQj��'9����b|�܆�����_���'�(��K'�-8��0��PC��P'�:Q�(�^<1g�iCj|P"0��a����'���M�<���ml�2"zd�(��:`l{y2�dD�O������pK�^�?(��κ����1u�|�b1�qq�-km��\�E�w�?6�{�^u���K�^k��f�y�f���w�YF^݀�cX
583g2���X겋靦���#���e�ԳB�Ŏ�ˑK��gg�pg+Ͱ���� @�Bw�+>�^5F6���mH�k�D4NFP�Kn�	�m���7�-�̳��fJa����	a?������ÅH��@�¨��,����N�X�l�
�<�־�w!�=�CG�B'����C�!�~�ԇD:t��� ��~��&u|o�D�p)���FN�`"t>���{�l�!�d:2lC����~616��>���<����!4!�H���ɂOF} �B�~7(���8��Mz4FC�5�(����O�zےĚ��D����ɹ�I��C��h}Ϲ��Y���R�{��퐋x�1�F�s��%ci��9㴦��<�NNiRBP?	�����~&�DCB%�'��K$�����(�x��R�U��κ�1��8��ZGȌF8�#o�Rַgc;����*��ٛ�"�yG�ǊZn���x�Έ?ql&���RO�O`��p��B�Z�4Q4 #I�Zg�����
�L��фܣ�p@L��l�z��������\K���pL!����<7�"�6!A'o~���	�5�(���E���&��$����0I��:e���y��ǯ+F�
���-;�Bs�m���>q�n��q�l���'��i`Sl�$ҺXNBx���4!��*P؛�	�@��L���Pˏ�va�@�yd=���d42X���&�
|XOM�I�%�(����`;���R&�o<���:���u�~DG]G͢:����|��-m��L�uW�S5�n��Mr�*��!�2t�I��}�ߍ�M,4x�T�o��ra���D'qw.)�|aᩘt`�r�!��"s�8�	6'ؾ�zg�0�?4ѨJ"n�d�K;��n�w�8MS�8����_���r��p���m�rL"M�k&��Wm��䷚�[m�f�����Ȕϗf�?	�6 ģ�?�!g��CBp`g��~X��W~���)�oT��1�����x	>��D��χ��i�a��.���A�FJ&��o#��������>9�^9�,��%'H�l����p�e�D�3�	�,o��N�����x"0A#O�����	�N6:�.-=0�qg�q�?#�8��Q�>G���3$DY%�d{w�bJ�������(��O�?h���00����s4]fc�)���!
Η�JڴZ�Z���Kl��۔rM��8΅��	�6���Ĉ$����2�)v"m��U����ޖ9�Up�a�"�'��M	�%I�)���0^�v2�ѓȝ��?\J��Y�z�<�	�@��K@L��	3�Ó�aʴEI�0���(�)�����a�&�'"C���Ђt�7�xd=ᓢv��Z+JZۓP��HDt4�0M��&A
z2������@�=���́�~(5��#��Ɗ~��	� �M�K�ق~6 lE8zY�ҟ�,d���+˷#�[���ֱV�涬b���/��+^1x����-���/x�����mX�mx���1�+L^Ʊ���k�W�W����cV��c��b����^�ƱX���Ϛ~~_�~~_���-��V1K�/��u\E�\i�屋Ɨ���b��/
�/���eV٪�qx���+��+���t�ҘV**ؼS�/_��/�^)�{U�k�^1|c�z���W�W�^1xˬ^1x��.��W�c��폚�/�/JҰ�R��U�x�6��U�/�b�W�SJ��_�y�_�_����W������V��/m/�c�k�.1|U�jmxU�x�V1x��.?.#Kj"�.?-�ȭU���^1�=�^-~�x�b���_1x�1n��^E1��c��:��h��i�Q>4zfË^+J�����|�S�\�y]
#"nfgf�.�Dnﶲ-Va�Iv��S��;�Ѥ��}{���P����T��<���#Q<ýn��
��7��-w3.N���a\�=���u�{�@��C��Wʑ�L��\��Wj�yE�U�Nݐ�j�:l�����t���z£;�]
��y�������ݩ:�)n�w���?W�n���MgA��n�ݕ�Wl���q(�����{j�~����WZ��睪EzO�Ͼx{7���M���w��o=��r�~u���>���F��-S��Ft��{�E��s=9�u�,�v��%"������oYf�|b��еK�J{��Ͼxݞo��v������%����k����'�I���Ios�͸�#p'�c����w�;җ�������n�y�i��������'��y��c�(Q���'�V�o7�{/K|��Nn^^mt����*�Z˷�N�n��&{?�.�m���;s9��\���Y�5��ȴ����Z��幬k�Bآ�)B���,r����VT�@�8���cxBy��{f�@��نSY.��U�X�eڪ�Jb�3rB"m�G)�"�I��km4�9�C:��˚	�P\�X�X�7,q��v.�,M�	&�p����U��6�Ĭe��H�q����,�:>kH谍s̖�奿E�
���������\Gh�m��m�R�a/ks&.@ <�y�����@#�}�������o��W�fe�������I$�'}�����3=��ԒN��g�}��=>cc�q�����Q�G�m)km��c��Q!��%ۀ��, �m�Ғ6�t#2��i�8ЇSd�-�\�
����f�(k�u��S�)D�)2�nĢV%5_��1��=7l��0ց�/4�&��a���Luv��ܤ�����5�f2cMeD����GmF.�,#�r��]��iF8��A� �%�
�f6MWe!�L�ZX�X�Y`�TK���F3`��omjF�j�M�K�_�$$'d�&<4�mY#�<]�ڔ2�41�+ͥa\���غ8��$�=�S/n�i�7���~�MDN�a����$���d�ՐD���qu��kFe����'��Da�DdÅ��-��~)d؅��"a���-n{Gp?	����-���%�ZuC�:#w�V�U_�jb�+Ɯ�b�;�mj�ik7��P``���ʞ�CG���m=��04}7f���ę{ |�y�٫�Ӝ���Se�B`2hd�aM_B��ᩆ�<�d�JO�����LG܃�0t��l7]�c����V�.jN�;$�0�֐4e&�,�D؉�Rh�
?EC�����o�Ļ(ȧ�L�ِ��C�g����q������D1G�L�ن�>:�!t(�A�DFO;0�K'S4n1�S"`��~��(I������~,�D���0����&��̹�������<��y���3��|3-r��EM� �A#�Ƅg��a���I���D����Rs�v�̝��������)d(��~+2�{��B�8��7�y|K�ūfL\l�jlܸyRC�y�8b�z�%L�͸@�""~���a�Sbba�	���m��<2��}݆�F!��0N��%'�z0�MҌ���ÔDw�;��lo%�r��ۗt@�O<�蟣'H�lu�:�1u":��h�(�Ad�O��# �J�#b�D�6Sf�#���a�'�
}ɢnRC���͞'D8D�C�F~'��~=ه�tC�Ʌ=�'�0g���������gƸHM�Fo��۸�XJ�B���L�Kn.\#�r��ˠś9'�����p�SF�WA�I��5,��L��2(0�(S�X~����4
xrɼ8�`���y�˛�O=,0���6�8g��!��a�(FJ�=��s*��u��C���!�K��\v0�O9�����x��h��X��8�Du�|��!��>zҖ��[��Ӵ��H�}l��࢑>Oql��M���c����=x �=���ޚ�4Sӆ�tId$���ֶ���b�X*RR1�ʶ�L��,#��X@�Г����o������zr�
0(�2�)����9㼥ޮ�|2x#�- �B�J&�å���N��ƣ���Cy�j�Ǻ��d�?�`�6y
h��~��g~mx|�2̅��0l�:�-T�uU�Q�ժ]�e�O�|0�� ����D�g ��k�Qq��zs�/���a�����5j񊦈�"??:�1u":�b8��������o>K���_�w~>�gm��oNtS���X��[ʷM3�>��]�t�j��V�;��֮�Bg^;�T�c���������&�����v�z��e���xͱn�.����%�'$��l��13b����'		.��Y픧����"� :ۡ�b�eЍ�elH�JX�Vl�Lu-��t��O�a��w��h'����!�O�D�9��2h�}�CEy��G�l���?z�j���y>�<>�K��٣�A���m��Y�C�nC��A7����䠜���h��lO�m���֫F���J)�UR�ϧ��[8!��L�7TkV�j`fc��i��,5��\"��6����A������6 i�w�������{˻�6��(�x��;5Z�G�__�������#??:���8��":�>Du�q=0JSf�81"�Y�O�V�e��F�J������S�[�x��>iw~��G_�߲��t��}z��eySϾS��͖QOY��{��[?	���J�I�=�h�;L������@Nw�~�usF���ɠ���ن͈ �w��0%��|�B;�� ^(|���=�_^H��#nv���b����$�c�����:l���狘Ze{2*�l��;U�M�+M8ᢏD�[�5�p]�~:~�����??1�q�"#���GQGON0JSf�vy�6�E"|la��c�Ĩ�N�t6y
<�Ý��U�,�AM�OPO00Ld���\�TT����A,E�گ�zŃ�>7����
:�hh$l�]�cx9a�/��=bF�YG�s�|�|�+��U��_���_8�T�O�m�n���n�`!���y���h��og�
nzq��C�'tJy�J#O�C�Cg�GC�6p���rI�Y FU���>m�~~Dq�1�Q�#��#���KZ�m~JSW~A7@��sb�DNk�m�;И_8!ш~�p�x=(h	?~�<�y(���0���s(�v�!�!�YTh�q�Fwr�?a�OL�@��"ntA8'�)�G<<��M&��f?V������D��8}��p���Q�Y��Q�.f`яJ|W�8����)��8�Us��u~b���W�|Q<�~�����\o�R�zQ�m�mի�u�mK[�LӞ[��b�s�?9ܵ�ӿ��9屷���V�Lb>G��G~b#��8�����֖�������j�Rh��I�aZ}WK����z�g8�����	�����G��ޝ"���.�K�_iW�/g"X۲B��u�+l�v�c�֤È�!�e�e�v�Y�T���mUn6���qM�3bV��O��	�}2��Ȏ�K��l�sH�%a֠��X��r�-�J�\]R�4ɭ؄�午To�	���}�{2�j���8����4w�)��;�\-T����4�0=g�]a<�y6��t��KO�X�}�bS���Nӎ� ��Da��s��]�[~?)��W��G��t���6`h�!<��~���m�d~Q+�(��U��S���<���'�xO��埉�vҝ�^��d�h�^{���+^Uޘ�x��W�3�)Չ�����P����6x�1���G]DqD1=8h�͖SG�Q��ьx(��Sn��_��:�ϿUz�>)��[|߅��㎟�y�*�ߖ��_���[<Զ�~;�h'?i}��㳇Jh�04	翭������Vҭx���X��o�qJz�����ͫθ�|�N�O'ϰ��^ݙ��2�AM�m2Ё%#6p������������Lh�U�e��~#�}�^O�c\��b���bp�Ly����Ӣy�PN�)�/�3�2�����7�{�z��*��T����f굶/�b��qLi�^ؼe�/�b�±����^զ�^�m�b���\z�b�5���c汋����W��b���/�qx�����5�^:��V=^1x��X���ʺ������5��iUOʕU��E���|�b��li������lk��L��x�1}TS��U�\U�t�U+
�qkb�X�|�W��V"�_8�n����c�cX���ǯZ���Xű��/�V1}c�=������������4�+
�S�^)�����ű��ڼҼ�����Q����j��S
��ߖ�V�^걶�Xˬ_�S�c�կJm����^1x�W���5qQ�x�~j���]V1x��c�ix�V4�VؼqlWX��+�b��g��t'�������|hK��׊i��.��V2�5�/���Q��'���J{�M�3�bs5�1t���>����z*s�!�Pr-)C��B��kbj�藯�����9Q	$/.��;ӷ��e�	��u������-|�U�(V������̯:*D�%j^�&�۝Kh�(��m{k��HN�3Тk�1�ԼgB0��q1%X�"�'���-�}�Λo�6��3>Ͼ�[m�m�͹���3��略�6�|۟�̠0�|Sc��G]DqD1=8h�͔ӡE"�)��xp���ڞ��:t(&�p�-�r~X�p��CA�@��5��n*f*x�á�L6`h�����W��=�����o�␬#�[K�ݜ��6�hCVT"6���/��	�ʽ?>[��?>L���)M[֚z鰾�Q�5��DK��&�~d�/��5`���z�Yxp���|���U�1ꔤ��z�e�}����ַ��D�DD����)�t)�}��Z�E>~|���u�DGQGQG���KZ�moZ�V�Z�b���M�ٳ�\~���Y�1N��DD��0��yN�8a�J!	��)�v0ݖ�f���7]WB��fʚ9�aUe�ϼ�h��"#��^�IO~7�����������ѡ<��5m���t�=�Ͼ�+���v~B"&av�79��|5�����â"]�Y����Ë�6h�b���B"�KY��E�N�jW�?,�DL��p��L�4��<y<�ا�G����G]c��":�!��>z�ֶ�[�~쥒��� �wVUyM�e�A(,�k�e�(M���izO�w�7��#ۉ�����x��wn�`�<Ls�O4f'��{���-�w[� �n��w�,��w����%if�����.�]]��ũpn%�m�\��RU�S\�&nr�3���9�j�	v&��a�vw��%��)|\M��tV(�͙���m	S)��rVƭ��T%M)I�15CU��%��,���*�1O<c��U�JS�b��x�OG�g���[��l��M���}֮\M����v�pV�:Z^Cg�?4`���h����c7�PٞS�s[�7'Ə)<���z�]�n�z��\YF�ʮ�4tO��K��<7��*|S����A{�^+�AB�}��^P@ ������i�k�kh�#k��&��p��ph�t����e�y��d��A~�I�;+�9���#�g�T��)�m�q�����1��":�!��>z�ֶ�[}ծ��v(���}�|[���)���!�Ҳ�ċ�^G K�3�&6���;����W�^�t��U馪��<)e�ט�+�^4ϼ�Mb����[a�g�.���Bİ�z4�)���0��u���,-˒�y���ֵEB��1b�j蝝��e0N��<4h��A�&���^N>���NO��x|z	T�i�:u���T�6Q�y��U��~im+��un�c�":�1��":�!��>z�ֶ�[���ɉ���z(��S����|�Zt�l�	O���WSTɣF~�x�:4J?�����������6hC�;�Z\����3,*|̻��m*d���J�2>*"C���a���!B(�GE��͛�$�2h�)Lyc����D.�0�8t��(�)�K�2��b���t�^:����R���('�yp�⪈�0C���[Sf��E>)����b":�1��":��=6zlх)M�(�g���&�w�EA>��i}�����ѽ�������2�wf����?�d���q�r#��\��+��چa*8�Mj<E��_��bqթ�Z�����J8�8��m��*�p�����JXp��8�.��/�/��0D?O�?¸�s�T��u��m"�M�������̻���ؕ`x"�ÿ���O��+�~u�֔[���s�j��*�I���_�|��oʹ�li���[���~~DG_��1�DuFѷ�.Ygge��Ù<ן��ֲ�~ԝiS��oտ2�<x��;o��}VyqǽbV���i� $ğ}lf���.�H���;�v!u�m�\��vz�3Tٴ}��i���3D&'�lth��Gv��XK-
�B3VK���T��ɂ3��:�`@����[
IX5�mъ��bF��9,��)�1;�ap �[a�5p�K�X�SM\�I��g�}��w���	�0A9��0�����)��`�ԧO�A2w�����>6S����WH�~���O����[n��t��ㇼf�6ܚ<(�!��R�o���sj6tD�=�m�	��ޖӰ�)��KEH�dvp��ðD�|��[~m6�]]S��j�i˥�&�mK���is�Vy	�0��i����"$OL�th�}
y�*�EM>u��E������Du��cb#��b6��ik[m��Ey�2��v\�x(��~���ߋ������*..�A�<�|��ص���w��|�;��)�9���H���&	������3�޿Y��h��C�2�*�~�O�QώCG��vh��C���7���$]X�7�L35v ��GR��R�.F:�t����M�	�
`�&�gb~?=�LD<�(wE��>���B ����U�}�������o�S���[|���":��#���!�m4aJSf�(��؆<u��("�!�8&��˗�y8!�m`�i�U��F��m���Ї�0M���Sҍ�7�Y�颔W�Ka���^]^�֥�~�1�n�7�D���L�PY�(m� �����DYlTP���%�~�(�����E=�=/D�r��N~���ɢ��Qᢟ��؈i:��Y��y~���*��D���<��G|��G�ϝ��ھq�-���8�Du�b1�Dua��f�)Jl�O=C�_�����.�Q+�F�8m�*o5�x(��t���Þln#L���ϼ�Qٲ��o!�m�$�����(��yr�U��
��ƻ-�h��n%50���-U��ܼ��e�1C���Q�6�E[8��J��]V�Q�ʦM,�L��8!Љg�־6��I�gS���V��z`��<_�U;�>���`�a�|�W��$uG>o�\�����W��J8����l�yF��V�)�0C%j�]�>|�-JS>w�{�ߝmӄc�νi"8�#H���""""=R��f�f1�c�a��8�0Æ1�����ffc��qh������6��1��ǭ��DDFЈ�#�GȎ8�#N6�)B"�h��"-G��#�����h�V�4�DDDDDDZ!m�רDE�hB"�Z��Z4�V�>DG�X��ź��T�#�Du�І��""">cu�[u�X�b��1uZ"-�|�#��#���q�>iHA#�2FiC�h�\*gJ������Rk���v�3g{��ɼ�ڸEB=��/�͑K�.=��^}��X�Y�7���x]�\Mʙ����F�$|���#��?wJ��^a񳞘E�]�̬����]Das�1IR���W\��h��GTYt�[��1AH�e%��T����~~�������=ER�� 0�qJ���ț�K��	��.g��|�t��l:��x��)h�j�{��O,����3_kIiFnU����S��7"5�<���7�O|{���;��̥��0��}�����YH{V�f��"m����I��W�ڵ0�GX�W��UidN6d���n���]�]��F������G�?x���0>�<{{�~��BˁV(�-���n��5Q�w]L�e��z�Y�t�;�9͕u�9�|x+�؇f���Q�R��	���F�MS�oE]굊�$�����B������D
oj�뮇�)�-�?�m�H��n�	�l͐G�%�`�rm�Ǝ&�a�TؙK�\�L�j��-sq��b���me�)r���f��,#	ƴ������d.ՙw3h��D�i�V&ni	bպ	,�S�o��D���.x��fl��5��ns�����!
hm�X̞�<S�B��9\F�f3X�l\�[J^F-K*m�#�cK2$�R�f����R6+��gP#5lq��K��5���$hk{��֒����}m��������v������Q�������6���q�����e�$��w�%���~z��c�u�:���c�uch�֖����	�Y�/�i	���*��gi;j�Ȭm9�J�`.�<nv�ܮYK�V���h���oe�Y��f�9�tK4e���k11*�uETh96(���.�c�ͼ5-�t�ي�����m����x�������M���f�W\K�W9�S��f�N�8��c5Z��[�c�e���@afY��,m�&�� @���N�<������L@R�<�X�lFĎ�KY�-��T�t`�.����6v?mlL�:r�s�S��F�)�8l����zhهOĚ6"�������������S*M4AP"L,�{H3��Ȕ��N��������;�4 �d���_a��Cnd�ѩ�R�^���zhA|���8d�_���FA9���o���M��r�#+�&��.[�b���yO���z�/�)j>�+\~u>�ޕ��m������n8�h�c�΢:�1�1DF1�m�KZ�mkg;oJ��EC�K:m#Á�-Fyx�7�U���=}��6Ҋ~[���P�O'q�R�5�C=�+��?G�4�Q��/`�"����my?*��JQ��-�����e(��3�P��*
�\�u�15R�Aif��ñ�!��O��=��e��D:�d�vx|Ţb���z�֣��m?#������⃄)��}�֮�J*t���Ø3�1n�q�]c�b#�1�DcF޴�����uw�j����U�袂 ��Q�>)q��,0@��G�c,�|��'t%fxB�<��<dy�[8�4{�Cz�ob��xl0C��-��e���M5��Ɇ� #�`�ԉ2j�K���U�$��f�y�;=axNL=��	��:8&�~?Kj��/NF{o����J�l}�[U�Q�����Y0S����}��}��ЛOɓ�h竹X��$� T )ڥU|ҏ�Z��%?1�~c�κ����1�u�ѷ�-e6l��v�\�111ࢂ!��n�3(�8d~0�?w_�v#?k�u{p�~9������w����R�.q���D��pJS!`��${cq	�ĵ���=��x��w��p.(�0dT{I��B�?-���
!ħ�X"l�>�̶b}����<��lN!�D��=7 �ߔ[q�0�l�J5*��W�~|�W�[�kR�w���dF��ɪQ��_���ÊJ=��ҧ�z�?sͺ{��~C�-~q�X�κ��b#�1�DceAY�EMq���*	��$!O+�fK���n*�d�ʪI	J@�F��=pm4D���6�_u�2]%�3!�5�{Z�=��6*\�u�e���LW1�SLk�2:ŖWJ��kM��U���FYu��l{�	H���b�\�F[pɛ]�,`KL-���cJ�՘�Pȁ�n����mB������wm)��u6��]yQUS�ĢIK
rrS��� ����)�:���C���~�U?�p�~Ԅ��g ��N|
|hІ��C��)�M�xQ7+ӄ7[�W��~S��O4S�U��Tgy����W7bj[��K���"IU��i�C�0�'�Q���sv�%ih7+qmJ�5$.���xR���]Zw��4xzu��Gc���F1�c����g��R�ٲ�Hࢂ!難�G4>�g����C�>0�q��)k�]]|�-�{���FѤz���gg���lj�{!	�ybH2�"H�N}��Km��1v�U��@�

�(?agڐi!B�ӭ�^��p&6�f��&r��.�7:1@�����qJYh��`��i���jh��o.g���l��m�C�f�GǼ��s�A^�=?�>rB���&�) ��(d���uO�u�|��u��"1�cDF1�m�KZ�mnx���!�\jI]PD=<�pþ�~L��ǳ��D6d���pن��
zSӄ铣ҔA��Ƥ�ɂ���m�fw.:��b&CC/)��Y�6uՖ|��W���G���őTt�C�6S�e9^��f��C�,N�І�a��{7�QF{0 A��f�ʙ��(�jbgK+ƒU�$��H��/���*g�$�@��^$���?���Ϳ4�H����F1�c���6��ik[m�K��UJ��~��u��j�p��1�mEy�x��_IevLĠ���C���S�}=O>S�4e��8�)���SX��N#�<0�����v��C�y�Ӏ�o����p����{�!F
a���͞$�|��%�/�S�4�?*��ۍ�J?=��_��m�~T٘��}�Z�Wp�CF=h��M(�>[�nV]�V���2�D/��)D-�rf.I�F�ۨ����GX�1�F1�mz�ֶ�s�WeW��{�E�k�1;~� 	�8I�9�C��?��o��놱�V�H@�z��	Q��xq����1�a��MQZ�Ϻ�m��Zr�Sa��^����{�������]�N}��R"|t��]�O7��A�KK��wlh2���Yv.�B#ʻ)kKvl�e����7]3�-u�V]ʊ���d��Č��gJ���	IS���o&06�u�dF���k�:Ťv�!)�Il6G�V��i)�Ѕf���eѭm]`O��I�'ߪAޱs�1�����~+Ğ\�W�պ�:��"����{uo-������B���|\�)����xF�!�Ú4h��~�Ԣ��WC�B	��,��D���(ʉB��Y����I^�t6/ğs��'��?z�]U�}Me��[oc��t����]�=u>�|��֎��)��k�\V��?��ja
��U>�D�v	iQd��3N#�c��#���6��iJSf�Uwk8��ˉT8�j#��mX�URH.�i�d�d���	R*��T�UL�eq��QAf�:\:zl�f��KKO}^�(�=�6!�� �G���է����S�ᕬs�Â	���N
YΏz� @��H¼O��6&iU� /�O���4!�)��4���3�(��=I�6�Z�,֠��f9t��6+�q�j��C�����>�Nvj/v7B ��L.�3O�����I"	<l[�f�"�TT|��W+�]_��u���0�����Z"#h��QH���"""��"#�")�D[h���帊DDGȤq�qqh���">F��">D#8b�1�c�1�3K��6�:��Lb""�DDz�G^��GȎ��#�[E�B"�DDG��)�Du�h�E�""""""4��m6��DE�hB"�Z��G�Z)�"4�1Hc�[i�L1���:ӈB�h�c�u�[u�Q�0�1�����DZ#�|�#�������J|Ґ�z�Diq֑�g�ۻ}z������kC���ƚ�$�F~/��Da�b���7�>�f;��A��{����=ϑ�㞜���O|�:>�۾������N��x��s.�~_5_N�lYut�l�[c����0����/.���G���}O����z�~W�ٞO��$��<�>��Xk?(+��b6�nέmU�������o�LQ��]XK���;K|�w��2�=�ߞ��������vJIf���P5����ӝ�Y�#oL}�{���~{zFe�o�<���<�#�lEM+�Յ����y{���ݶ���y��}�}���������������o��g~�O��cc���c�F1�DF1�m�KZ�m�{�V�EC�|����|>�r<Ȝ��xs�9�Dx�-���_ǫQ���UV-^�]����}�ty]��L T���u�Ķ���]��;4vd���L��B���33)q6[���Ԧ�)��6R�dc��'�8t�� Đui�H,�8lH�c�c4������i)[��	-����D5=|�k$��6l�~�nz�]��=6���F#�1�1�Dc�DDcF޴����r�D�O+dҲV ��(��l���V;�'�^��x�X��|���)��)���i��^�Z�*�.a�#K,N^b<��a��h}�|���8�~)�G��`��G���5���_Əߋ:&�*p�QN�)�zd�B����}kS�8Y���y4�F����/����M�KQ�W�	x��/��Ǭ��C�I�;�e�V�Jzx%�}�ѱFcχFo�5W�<¶���q�^��q��DF1�1�DcF޴�����|���[��W^~��Zi���n��:���´k=5eb��]�[1���S�Z�a E6Ҙ�nD]�e�\�[t�.+au*��ge��`���[2�����u��p��'��A��� ��m,���b�˄��^9�\b�Vm��M]qlٙ]�&&8���@��G}z/��D!"=��<�.�ֲ�m���D���Cl�ᩲ��u���ֿK����u�6z�Ky��-H���<ۏ��H��V��j�˂1���FF��ge�>LA��|h
�4�0��M�<?lM�O�>���O1��O7L1$��&+qY�U2�*4�fF�kK�ې���D�ԷK��ڷBzh�SsgO���o����^��Q�q����u�c�ch�֖��ۮ�+�]]�X�DO�dz�;8j='�DMY�u��sY�8p�h�`������3ĵ�_J�UR��|IR`!A�[K�e9� B?zH�3�H_��?�O�hf��F��F�ݧ���5l���d΃1�Xͦ�vk���Ybà71f6&��.�OL?^�o��P�����}��6�a���
 �e)�/��BhJg���XS����7�|�枩�����\q���F1�1�b1����Z��i���t	MKz�^��	�&�oh���R�/]黜�vzSE)��i�V�z��E�^&���; ��٪[4�J]@��=�d$Љ��>Vjht"���b[r�ܙ&QM�¨�����7F/(&�f�EJ=�f���9X�$)A<����O��o���Y�5��A��Ұ������Ig�	�<�����ƹ��)��^��+��� ��d�?4���J!D�0Sd�=�\�b�d�SE98h^��|�m6�����b#�Dcc�#��z��m��<�K�w3�rVK爢��9��Z./
x`Q2"��� g�xx{;?��K!�����3F���A`�F3K�urFM�v�+����oXS����O?(�O�f��U\���Z���/�C�!D�ۻ��k��<P�jO)���.�`�,㐗��^�#�%���{�_��iwq�����x��3
�:rPD�O*?�6kb�`a{=50E)M�o�����M���㭿:�Ȏ1�u�c�b>m�ֵ����_�e�Z�L�����s�q
ͽ��>3��)�[m�憚���R.�zdj�G�.fj���D��R�]�$�J�Ѻ���/an��`%�qiJrg sn���B��~HB|�!�d�*�b�M�����s-�����4�͉vt�F�N�8��%��>�6s��W'N��A��/m�BU_��Q�`�%��~�0:"wKc��n~>�>�v�1�1qQ�a���N��h���Bo���P4o���؝��ٹ! ;>O��i�O����(6��6lj�*�C��#3y�%��<�����YM�y��=R~{�m���sMj���)�"�K|�]|���b#�Dcc�#��z��m����K�"�A9D,)(�l;��;�|��Z�4��xSE"3���(��ZQ^6V������A�/�<6a��kɹ��(�y�p�k�ۘ9k��٪���6�p����`8%:�	��;��^�3��n�ނ�jXa�(ë�G���F޳-��40���J"~�<4S�_���չ�D�_����Jt���Xv}�36``���o�#��P���{�۫��+�emKu��q���b#�Dcc�#��z�)M���&���A��d8~��p�)-]�ךR��R�md�Q��_B���I�Kq�����A�����L/��rJ�M
�6�,]���Ç+c'�B�|&w��q.�$�O�~?i��D�amxl����O���uo�6M��+�FZP��I�(,�/���ȿ ��JB��_~��U[�,�0����}���޶�u�ζ�\q��1�u�c�b>m�ֵ���O����P��+�ۃ��ݛ�0M�f��"�R��յ�OE~�`�w�\)�^�wsG�{q������{�T�ƥ��m�a����L�i�Y�����h���a��S�+?#j�+~6~Ԡ�6��27<�蟍�C�)�'��{�kZ���ie?|����_��߄UU$��E�,��I�����ґ��R�j����m�uo<w�^4꼷��5��q�??1��""6���Dqh����qR#��">mG�|��DDq�>|�8�H�c0c�d�c�bb�c�1�c�`�0ጔG��u��1�|�"=DR8�[D|��"8�h�!1�c�`�1�32FP�1��-�iH��":�DDF�m��T�DZք")�ikDE�=Yh�Ȉ�n�#��c�[cjc�X����DF��DG�u�:믝uc[�DG
DE��GGQDu��Z>iO�E���1�1�X�$g���Y�Sb�W�Ӣ�v�x�Y��٧u����^�6�y�� ���y|r:���{�+����Mq�_�>)���vS�5*������z����Yfm�ndW;W�VMV*�Kn�eF�T�Qw%;���H�=�v���}�y�zc����?;����؝����͠hs��i~}=G��{��i����z�|��gvL�l��L�������S��{��{���'��cR�[�N�x��1�{��+�S���t���]ՙ	RS��U�S�*?�n��,�U"�c�W����Tr�[gNY�ǧ>'A�o��mr�nz�������G�
��>H�.7��y__C��7{�O2���>�g�ӧ{=#��J���Y�k�_�\�9�������h�_:��������{W��u������k��|�=�=魣}=��}/����q������z+��H:#wwv&�b'�3��L�]LUR�^�=rGw;������N����'/.��ʹ�L$
�Jz?g�td�((.��
렋�u�i�q�"�E�WT㭆���s��-e�e�ٻ;�:�ඁ�E�5�p0+٫r�e���["m�5�ei0ս�*���ݐ�t�1��Į�s\۵ ǵ�x�u�3c���2�g<��1We`R��n_�c�� <Ot2�u���mY�o(�6�&u[�W,��l�� Ґ�[�A���k�^�PA#���ř�댲�jɋu��a�)s��C=KR�<4G
w7m���m�}������}�|�m��w��}����ɕ��I9;��>�����:ۮ��b#��1ǧ�)JSf��1f[��s%���p��u\�����p�۶��鳡�PD�K���v%����K���k2�+!��1��e��!�)�1,w&�4gZ�VW�4e!�m��:�4��V���H��fW3`�dQ�ejEѷ%�$�Kԍm#�9e,-ѳ*��[��b�@���A���F�:;FU��릎[H�s�(�:��f��|� t#�j�����E^-Q �'CZԔ�(�R2������0���Y�����h�Nz��il�f����j�i�$�Q�(��0�ř;��NE��7�I��LD���}�"�$�H#����KG�����SG�J�VC��l�N�K���2�ji���C@ͧ��C����xd�z�E���%-̦��ֆ�n��)�uW��w8�M�r'~(ӯN��j�;~~�G�~~K�^��i<��]S~|�?:��6�8��1�u�c�b>m�ֵ�����a=C��R��T
��J
�ue�b(�L����4ni:��<:M�<��񫚶�45��O�?!��x!�|�<��'d�Q��Þy)Z�j��l79�0١����sg�SP�Ô)��v?�Dq�V@�2��DϪD�L*D�HM�l���M�2�1�M�Ҩ�������hi��|f��4��}�}��;(�x鬶�mf��58d��4}�G��f^����~ngN&|���@!i�2��i�c4��u�c�16�kZ�m�<��)Zܽ�(�F��g=�e�8?l�tg�M||_t=?�O%>���(֙��6`hJA3*�C'�d"��� (�|�l�1U3Q�sGl�F�\]��I��^hy?�Ǡ���ޜ����FI
~��w��9���9�Wg��M��x~��}��&�ᑶ�sF�3Bw�ݟ)��Y�}�g�?/��_LX�&��֞^�j�^�ۨ���b6���X�#�#�ޭJSf����bVJ���Yv��𧇢�ZR_D��(S���t��S���Q�e�MJoV�Y]�͕�r�m͵IB�QDȢ�h�Ix��i���g�J���;�������tB����מ��ʏU�x>iO[]��\ V|�?� �}!&�號��jPvg��0�Ś&��0�00�O��M���e<?E�%��I�g�F������(p��'G��:u��>u���u��1�1��#�oV����>WT�j�w��n����"�p_)�	[�������פZj�R�SXct+.<]����β�Rۮ`��H�bنܠK��f[�����"Wf��]�V��҅���� t&�a�F�9�au"@Y�6Rj֑��$��3�֪�����w3������E�K���Ǧ�M`n�m���wG��5�.i�4`��f��C8	TJ!�����{�Ur��p>fOQ>�N�$H�~.�",�=��s�oUj��֟������i��m刱�3P����ң����IN�_�Ç����ksTtjꖗ#�h�@�Q��`a����8���Z�dޔ�����h��A�hf��`�k��Aټ���>F8���Dmu���F1����Zֶ�{�4�]y���X!���!����	���a�������^�1��֋)_�~g�����SK���%�1���|re�~KC, N������g�/x��$��� Ek�K���X@�o虘��iR����w"��2�1MiZi�s�V)�>��LYi�coJ��.j3f�w^�=�!|�8$�h�����e/���f�ݫ�p��>#N�����<��8��1�8�mu�1�F1�#��R��͞�����1&�LΪ�#�������C&����h�G�a�{FY ��{D�JL�_T�L���P��
�=�l�ѿõp�_����Ɠ�����\�Vh�XE��R�8oFM�0D�����Sc'�e63�Gɢ���$6h� z`�����¾k�܇��>3�B	|?}^~3��3ٳ�oK�R���m�:�>u|�?#h먎1�b1�q6�ֵ���9VV,!�SCh����co\UPD�C�	��겉��d�Y�!��(f{��(��H���c(D�Є��mL�ҢQEx��%T�=���N�4L�ñ0)�!)Nx���� p��;��am�S^�k�:v�Δ�R~�wkW����0�g��0��?~˗$=9�N�V�?y�Z6ۯ�+m���UyX�3)U'���ҟ�-�6�4��Ƙ���8�?#�u�G�1X�$�,�����)J��H�c]hWX����ș�v����u�����p�g���������/��C\��y��{����v���O���/cc�M帔����.��43�0�;<Ǉ[l�就"%�h����� $"y�p�8�Ņ�� �6WV'!����l�1���2�a����&��3t�����#{�#��"u)�4�$�3K^�ق~��?n�\ב�	�I=�4	�Cܵ-+�G�6h�I����F���.'��a��>d%�5���lB��40��ɨ?r�31��O�҈'aڞ+��z����g����iPZF�b$l)��ˊ\�O?^->��� XS��[DEn
��f"hϒ���?i��q�G�먎?1�F1�6���,��F�A��E	"������E6�ez�}���W����R��=�u=�<�<�f�:<>/��$�30i�a�8�K � ^�c��//F�ϓ)�by�}�C��}]CA�6YA>�S{Lt��mI��a�2sґ��є�)�S���Ŗzr~0��,��o�cr����p�����:S�W$>���i�įs�[i�؏�.��yk�)E��W�=�:��wϞ��>~c�"#H���Dqm�#H��=Di���D|��G�mh��㏖��8��DD|���R""#�!�c�2�1���c�g"�uH���1���c���>Gu�#��␄")""=DDi���H���"#�������|���Ў"ִ!F�Z"#H������n�":�|��=cc�b4�R���Q�"4�]q����Q��1�1�E�#�F�GE:��\Z-��JB��1�1�p� g��pn��m�GH�JZ�51/Zc�s%u���n),���D�G^FQQ�J^]�JFt�z�#j�)���o`2ꊛ�WSJ�8s1r\��鹌�Yu
}9<����j����ӳ�\�^iT�b5b-I�e�Ko3;��\�+�w���;�-�W�Lȼ��_���3�D}��}ߛm�����w}��1��o_w|}�w��}�m�'{��V��z�lc��8�z�����#�F�ikm�ںUzztК9g��ҧ��z7(Q"y�~��n�[MoU�����=)<[��UuU[6�[Om��y�?�$5WZ��Q��	�`��WX�i�m��o�ɡ�:��_߰�����S<5<�]谍1��m^[5Ull��2�����y^|�x�[+̢��~[��m�g�(��M'��)k��:����mD~q�8�G�먎#�c��fR�0���c�YĐIP�PO���ߺy�M2CR�(���H,4y�Ӏ����/�F�[�{��ھ�Ҽ+K�sS �Uie��za�����mPA�t�>�W.aZ��h��W�6���y�L����V�u�ص���y�75�Қִ2�R�|yKZsj��3���>V|�1B�88�}�|4͢(Sپ/�]�q��?1��Uԣ3pB�|:h�ӆ�sIOθ��uq���:�#���#�ͣm4���o~���W/UX��q6�:i���5�*�v���&c�������,X�G��������敄k�a��b��nP���Kٚ�j&&F�ͮZat%,����z[c��Wt׫�*ʚ8�_�����+>
�LuCQ4$`�@�i���X̲��+`nkdF�nc4��#�Fi��63���qrz&�<:C�(gϣ�y�WZ��u莍�("S�jP`2�z_�TT�)����ئNB���B_�G�L�Q4U�%�pI"?S�g�����<4_���;�s8p���A5�kc����MMϞ3a��!�@V�k'����=��rPnH$ ̅�T.��Ч!ÐMϏJ}έɠ�|��y�x1�j��矵g�c��8�?#�u�G��F1��F�ikm���u�p�6�vRt�'��C��c�UPCr�4Q)�t	��j�Oх�xѥC&���>�:��J~�+�@�Q��J������@�I,I(����e�}��}^��Ze��"�!- �(,դ��`�h��,מ�M_��[gU��t�z]4���iw4&�( ��%�0�L,U�U�
��4���S�f9n"9>=:v�4������#�8�1���8��#��F�ikm���Ő�(���'���Z}�D���A�=T��Ԧ��hΝ:�0܇')}8x~s3�i�H���^��|��w��	a�,���iR�f�N��/t�6=,)�p�JQ��l�[�@y�i�������8�=�/�EYs�OOI�'�*�4�����4e4	G�7Yr��j��ʜ>h� I���Ra5��""f0��}gh�d��c��c~c�8��:�#��b1�m�m����m��̯8��|��PNĹ({ز�4	{,�����K4�����9E��	m�-���HU����@e�Yx���?}����h�h�e���Ng�j�Z�Ehr$�0���g��y- �{���W�2�1�fF�Õ�o�� �|qG���w�?�3)�������p��sj�CF�����{92�l�x]���w�]ߟ�EF1�돜q��:�#���c��m���c;�)���5b�Ɓo/{��|2����jb$8^el����BXT���kDCޞD��.���v�FbԻB�j�˵\;�鬫\@������-��"EX4#K\ �)t��b�eY�NA�t-e"!��!��Ő�0&l�
Lfٵ�ʠ0,  @2)�џ�x�㟗��0�ύ���Ww⽿7�U�<�#�6�۞o�R����F���������<�قy���M���w���L-����`˒(C"��Gʓ�W$3��hp�Y��������}�MvJR^-��Mpɥڹs�'i\�U)RX������~HC��N������ofϏ��,�m�o_��|�F��QDF#ǭ�m4���i�V��uUT62|'M7ȲN������@�rж�T�������B'`���x�4x~��W.fM��Oʽ���4���޵�U�V:c��\ngӅ�8`�<W���}q�ˍU+¶�4J��FT6�ѬEu��w�?��i�'��d���3��)q
��߹�]ի�O'O���Jy����(c��m�[��h������ga�a����u�Du�-�m����mگ�.]�6���@�>$r��5��g%0�:y�J�&���*AU�w��4��������	�?���o�?��IUkn�w�"���])C�-�,ܟa��4�k�a�!�N�z�3)��:	ârp�Ir��K43R�{��f6��ӊ��/�=�N�	�߭�̫�����d����ð����^4���??1��8�iu�Du�Ŷ�����M������YT� SD�%@2�;Ҫ�V�9���mg��������h���s���a���x��y�#�B�V� d����2�}�nl78l�Y�~-��٢�������B���BG�"<#�J�&|q'��-=C�i�U*!L �?`��C�R��>��3J�x|nPO�Jt��qu��@'
h��D7��D�`�%��B�#��e���i�-���]ch�GȈ�":��DD">E""8��HDmDGȎ#��OQ�c��a&3D1�1�c���"#�E"""">u��c��3�!�c0�cƈ�">i��m�q�1z�q�|�Z��E"#��P�1�1�c��I%�P�1�1�e�c�(e�Y#�Җ�E"4�4�DF�F�G���n����ר��DDuh�-c�=c�"4�]q�:뎣lc���"#��DG����#��Gz��n4�!��=Dz��	�K���ژ��^���cʋ���[��wVe��	�*y{��_��M���a��e�,���u��C������f�?����/������|;�#橢\���u�d���d��4>�ȻB������~�J[-���������]:
��4����Q��b���RժL����J[o���W�+~�=�<��n��wT��Ĺ��!_l6�Ǽ�/i��|��ާN���CǙ�j����p�;�I(��I>���X��|c��# �&mގ�iFS�[�e��ӧ�g��p��|_��B�,��=J&�6q{��V-uW5&t��.�JŊ�m�]�Uu� ��j4�������]{7�����дON�^��$%�q����R����I�D=��zK�m��;ӗ�wf��/���y��6_oIO��N���O��oo�X�����׵��~'�=�y�Kc��Vؗ��
�IsT�v���c߇��}��`��+�M�����c1_m�,΍m $�>���רll�m��9Ln���f�\Tnf\S^��V(����/-D(���O����4�m��y�u��v㴺���k���oB�jM��r�a+� �2��\�3Rj��ؚVwN��Ηc9��'M�ļ(�s`��YKe���,aU�m�fʹ��g�`�F l:��MH�[�z�"���Uk.�!�[�pb�Ͷہ붓f��&ʱא�#Q,y�����Ϭr�I}4ɵ����f]YM�
ĥͻE`@f�MY��T���ю�v˂�2&�8Me�Z�$X7l]*��?ǿ������Ͷ�ww�+�����m��ww�+���33�$�w��eo{���c�>q�#H먎"#��1m�m4���v���?}�e���a�n6�3kv]p��vt`�e�U0�i�k���n&#������kj�̢p�Zbڸ�\��k���3�`��n�a0�͝6t�YlU5p
�l�v��d����j�M36�-�Lj��H��\l]R4������A�0��-�E������1%x\��[z�V�R��9+�,m�Й��J�մ��Ai.���zk|R���k�u���$��`8���n���a�&�]�i�ls{��J���Ee�7h`���]s�}��/A�Z%��'{���v|�D�Q$���p��Y�.���&i����H�	�)$SA��?�=�b��/~�m���X�ܔ�gǐ��F�ACy�u��6P_&i?p0�|t����,����ʶ~^X�\dVZ훪�MɹT,9Z��?M�J��D�;����(1G���cWw��:��Ϟ�#���1����":��b�F�ikm��`Lb�w�ȲoJ�#�h�a���ke��<��o�6�:	ϔ������h)��y'���M����)��>
S�V��z�`�����}d�H�W���I�p���B�HQS	[�I�H�9���24,�8so��6���G^'N\�˜�ڪ��<۩�=~��_��9�Y᧾g+�Wv�}�3�|���F8��E���8�����ԧ�z��7�e/6��(��}��G5�T����;���Uc�1��=�=q�1:�(����Ump՚M8l�z~L�}�7d��/;ﲇyj�\\4v�L��@0���v{�������N$|>7����V��/�Y�L��ٯ����~��^Z���{�/Qc	8^K̓�O�q�#��}����/�;�a��J���|�ո�u����G]DqF1��Sսi��E��׵~{���:a��UPD�O�]�p�SE%�U��B����c���������+�ЙI�U�3W4]6�l��������xSE<�|r|!����Fژy�>5�ٳ��o
~�
z~?10�f=or��^I��8��/����<>���y��4?h�x�x.��Zi�ߏ�W�~1�������"-u�Du�6�OV���_�g�D���Β��tu���A��q���>�?}4qs�bn�mޟX�3fI\cF�Vb�V�����b"�ڬ��������|@�.�~�p���m����谞^�ett��6�h���#�l��h�[�R4��m���| 	�];��R�W�.���d���-�Y-M��6�CM睴b^�0���;�T��F�)�(a�"~��p�[0�h��~G����rS����(W_~���������||�gƿ��k������y�.S�6�~^tto�1d�,,���Q2a񚹩�{ĚTJ��������Κ)C��O�Or���i&  "bLCL2����m[���\�d�D��%���р�����;��:^�i���z�;��1�9����q�lq�>q�����":�ch��z��s߯�Z��r���i������vO�*|#��ԛ�9��Ꞿ)���DWX�4���J��DOJzl��#ɰL��kp��u��_Z~����=���m������{-��B�%ٸ�9Cgù6L�k�����<�!�MN�������A�-����V���jR!�	ɲ��333���a�N;��ڛGͺ�|���Z:�>DDu�6�OV���R��ǕF3�U̷D(� g1UN���ǜc64w�����[cgMN<��P3|ĭ��toՔ�>����@��	M��-x���_��+�rR�2lW	��K6.r%�g.?���>K���������w�?>a��Ͻz���V��k���b�A�teMI��7�rp���B��J}Ge=�HpO��A�~
�b�Z~����U��޺����>|��-u"":�ch��z��|$�B�g����b���Txh��Um+z��c�� �H#<y/�AG��f�i��9���p�dM��öE�m����l�J�B"
�UMUG��{����3>����>(���vԵ�����0�4{�A��_�V���������S���Ɯb�={���<���_1=�5v��׫{zi�Mk_�_�ٓ♞��!��3P��>7�y{�Da���s�<`EU�O,�xh�lu�>|�h���c�d&�h�7�o��
��թ>==��}� �qçژİ��H���L�VS��厭�Y1_�&>����5m�dKrd4K°M���fY�[����L�I�&�,V�'�@		q��R񉮖��ZSl5׉����X�2�H�K֮��Ҧgm�&��2v��Κ)ѳ�����D���&�"a��l��t��|��]����a鰧�,�O�&��a'���w��׾��}�Ξ��i��6�Ř��<��3]-���D�Ov���i��>a�҇�`a͜�}-D)�Y��V�- ���^�Hb��,S�����C`��J��'�8�JngG��x|D���L>�Q��6xzq��]F:돟8�Z:�>DDu�6�OV�����y�Yu�ڻ�s�5⪂p�~ÑM�0y��i}Tw~6jh��w>���~�\ˬE+A4N��͓^�����z/~1N��H���P��YL��P���0��M?w���~��Ӧ�!24�4r�����!6f(^Xh�,�+��=�B3��w�+\�Ms<x �v%8t��6zh���0ngL�6v1��_�\G�?"6��Du��""#�B"6���#(`�(d�c0c��1�ec4�M0�h�2�1�c���)�G����:�DDGGE�"8������-�"-�z����E��6��aR��#1���cC�2�1��I$��c(��cX�1���Ye���Z��i��4��F��E��D|��DS���H��DDuh�1
c�1�#��:�8�\u��cz�"#o��"6���qDGi�"�8�-HqZ#�B�h��}�S�U��*Q��5�݊�tby����2�F0��-����ױv�$���(P��:�}���b����"q��b�m[�����/�Ws��	
;pW�ѕ4K}�6w\�7�eg7N�1+�f-z�q�P	d��޸���ܦ���ս���Q��F吧*Oj��Lz=��Ab�*��n'�D�1R)§<G^-����c߷��t2�L?-�^!�t�+n�x�z�4�ž����q)�^�ՓzUuvJ�\�6&qW�]ސ�u�����!j�R�g�F�k��̝ˉ}����m��ﾸ�����>m�������{���ʒI$��s7{߭���]q��1����DcYM0�C*��`�0��W&���ӧF�R����Pg���68���� �x�|�(���Մ4�y&���
�O�uvż��
ݬv��R�X2�X���hp<��w�I�$���{������P<ͮ�Gac��}�u��ihZ��M�ԭ����"	q�_���Zi����q�c�>c��u�|���#��ѣ4}��Ql��Pbs@��	z���l�Y��T�J!d�jktk5�[�*ׂ��>��S�驆~��U�Z��wsQ
=�������+3�@��q�ٿ�m�<����0�4hO����8d��Yt���t:lO���c��A>����C���R�|v!>S�|�Y��;�}��u��㨎8�����Q�"""1����f��������n9�"]Rb>�6Q��]��E�u&���&<Ƶ��v��������n��ot����oRi�/������1�X�����O����؛�.��оYko�Be
��5�5�Ό�w,�[�;lL<]�[v�C84J'� $'04���9�0�ܬK� 2�:�ז��]RRmK`0�1�B���\,\k����w����g�!��㳳�J;Z~�x��[��(��ё!�
�A%��C�߼QD!vxK�F+�>���N���2��='�s�֧��%���Kr$�Fi����	�w5�6�V��^4Q~�4X�N͇���A��Y�%ֳWM[�����E�ű�j�/	fc�Z.��D�����f����Izu�<�z���w�ũ��]�ܷ�����_�q�:�G]GȈ���6��z�OS���|�����.j�R�K{�c�ͪ�Mֺ���T	�f�A^�zY�U*���óZdb�#L4t��<>���ĩW��Cg�7
$�0�eپ~����sM�`�T|=��`}զ�ħf`s�~�\j_R��Wi�� �)O�7��<���0�D��<��������Ff�a��t��?	�:'�g�_�z������KQ�׉i�\�O���f�a��)u"""#��m�M=<�G˙�������y�ֶ%����ܚ���K4p���~�8#4���*��<�=qy�n���kl���O�\,�'�Ʈ���}%5�L���Ζ�G��.n�J�f*UUz��)�����⍑}!V?�ۨzl����u��ci��^�|
|~�V~���� �"�b#�o���߽|�֧����������_.��U�t�U�y�,�m���8��"�Q�"""1���޴�ס&���F�Cl�5A ҵ)'�%�Mo�U�M��Rۍ}|�>|��}��z�k�z�F5��L�[�[���:_�B�z�[&*�"!y�c�6׉?S��50ٱ�C���4j	��M�ُ�t�fNC�ᲆޯ���R<0��b��>S�ⶮ�qӞ{�:ի��������g�h�Z���@���r�����2��&�V�_��y��]�4��8���:�㏘�G]GȎ�"1��SoZi�!�W����4�W����>�bf��9�z.�x/?�o���u��X�~m���Wν�|�t�wi��KZWM�����.BX�{v�jU��+v�+l�ݾ3�<�'E��:�Ӵ���a�| $���� �x*�0�7�-aS��ZR[H.fq	ᶘ��3�4���f�
�d��J3�M;å�8O3�1�Oƽ�U�RɆ�a�����%�����_U�6|%�8tq��(�]�S<�l�$����'����<��=�R9b�Z�	$���8|'&��5C��}^b?C���S�ْ�Dwe(�=�?O�/d��v������ψ�K��t�=�ea��x���0uɬ�����Fs��F���r�D�+k~���uu~Z��z�1��q��D#���GQ��)��4�I�ɤY
��P���G>���9���G�[^"j]���<�:SM�~[�$�ӫ���L��"� �j��xP����o�oŜ�>��'��F���h��p0ߚ��R���iԼ��#�Ju�+ͶQ$�g~J~c'YޤQ�h�~0R��%I1�l���D�.Ԩ�J�ߘ9����f�s�j�f92��'$�G�r�J돖�_�1��|��u�|��"#�e6�����(���&ZX�(���1���ZҊ���F+1+S+B�M���AdE�^�U)�Ri�m�,C�0��Q�J[�->��l�B�ߛ�J�Xj��`��MCsD�����3L&�ݸ��z�%�9I�q�ۃ���f��f�FiJ	aJ�WA,��<(��4���$�|�퉚�0:rQ���4=�ggL4BO�A���ſ9��.�OZv�(��o�=X�">���,,�/@b���/!gt]���f��u��G\q����DF1��m�M=u�������ݣ�֭��wq娜o7��Th��_�.��ϓ�ͼ����כ��g�hp�O����⍳l��I�V�It���v��B�˨MR�[s)y��p�k)�EF�t�*?I�ޢ�J	��%��B$�������V�c���)�*�����<=LYO�{W���ܝ4��Mu}[Zj.��������l8���(3D��J'��������{�K�h��[z�����y����T�K+�UUUf�l͇~�c�m�����_�ܹRx-���&`:l���Y]2f�8$�&���3�,��h�����"kmm&�h�"����e���DD��E�DH�؈�E�b$H���E�dhD��Ț-�mE�mm""�M�5��D�dX�h���[kh��-�""�"&�kmdDDH����39D�m�m�5��&��""h�!D��"�",DE�DH�����dDM�4[DE���4M�dD[D��dD[DDE�M���"�H���DM�dH�,������X�"h��DE��&�DD�dDE�-����E���mD[h�4D[D��"h�KmdDD[D�4Y[h���4H�E�Km4X�DE�DM�-��mE�B,�""-	�E��"ȶ�DE�"ȋm�mDE�DDH��H���mD�"9�sfs�DYDD"�&��km�"",����"�DYD�mDE���mb"-�Ȉ���-��DK$H��I���h�I�K$H��"�m"D�M"Im&�f�"Id��M"K5���4��Y&�K,�$��$�"D�E�l�ZM$��"[H�f�d�bI�m$�5�i4�D�d�Ś$Ki%���E�%�$K$H�Kii,�&��HK$H�[I"X�H�H�-��"D��"Y"[Kk4I"Y"D�d�K5�i4��,�&��9�slrH�H��ĚZM"�d��%���h�,�"ZIi,�H�K$Kid���%�i%�$��4K$H��$��k5�%���D�Y"E��D�Y"D�D�5��E��$����E�KD��ř����E���-��4��K$�k4����,�Kkiĉ4��H�$Y��$Kim&��%��5�I�M"X�"Y��K$�id�D�Mf�D���"[H��,�Ki4��-��%�8[4�ĉbM"Y&�,�HKi4�bD�D��l���I	d�M,�Y��I��ki�XZ"Z[K,-Y�Y"�%��D�H�f��KZD�d����,I��i%���I���Y-$�8[%�%��ZKmd�i%��-���--,���h��%��h�ZI�$��m����I9q�$Z�"ɭ$��Y��ɤZK4��%���D��Z�4�D����I5�ZD��i�4��1l�~�l�e�f[-�[,5�6[&e�͝8�]�\8\2Y,�4�[#e����3[&ml����l�e����mcY�ŶhLhX��!�6hL�٦�d&hLЙ�cBl��bC&�hF����!c!l!fB�bd�kN�q45�md-	�wÍ�kA!@�	6�BB�HP�	6֛I��k#I����4�Mi�k&ݸ��p#&�&��i5�L�4��D�k&�kFD�5��D�Mm5���2Ѧ��D�5��Y4FI�4�Mb5�D��&�Mh�kh�M#Yi��M�M	�4�Zi��Y5��M&�k&�i5�D�M4dMm4M&��i5��Mc���M&������ɢkHȚɦ�Md�4Md�5��Md�4Md�5��4���5��4Md�4Md�5�"i�[MZi���&���$��D�5��Md�4��ɦ��5��h���ki�2Mbi5��ki��5��5�D��D�ki�kFI�4�&��&��&�X�N��Sd��iɢhMd�Mb2&�ki����&�ki��#-��k&��5��kBh���&�4�D��Bk&�����4Mm4M4��D�Mm&��4M[MD�ɢ2&�4�D�M4�i�h��ɦ�k&�kBh��D�FX�""�&��""�14B",�E��",X�n#&�"h�,D�m�&&��4YDD�D�ȶ��b!E��,D��4[DDE��-���&�b-1"h�$["DE�h��YDD��"���,��m[i��"�"",�-E�DYD�qm��h�&��!dH��YDE��h���"�h�$YشH�$H�-lZ$H�H[D�[j$Y$Z$,�kB!F�ؑhH�5��h+f�$Y�D�d8p�q�q��[DE�"�H�ؐ�$Q��-��"E�E�hH��HYD�[e�D���Z%���X��"ȑ4Ym�"-",��"D[k#��D�"E��-�#Y,����f�h�"Bș���E�$Y�D[kD�d&�""���"&�h�d$Mm�DY&�""E�5���D�"ȑ4Ym�,���h��$L���,�E�"Ȉ�mm�-""�4D[[h�"dH��"� ��ǌ�m<g���d��Y
C�!�?�O�^R���fm����S:ż�y{?����w�z�7��g���տ�=��>7������o��:�o5�ۓ����~�ɫ�{����������ӮW����b3�v�ߏ�����x��_����������6뷟��������~�}�l�����!�6��D�����Ϳ%������.��;Y�g}�?�s��OG���_�'W��N������^������IQ�8����~�fz~t���C���':Ϗ;��ߢ�3����t�����n�����=��s��N���{�ۮt�nRj���}����[��5�������f�m�����6����m�f���d����a��m�1��!# I��z@�Ic���!r�~����wu=^;�����l`�6��$(I������f�!�l�&m�s�~���>�7�;�}��{��|����7����x#���g����?�����mW���d�6fÌ�nw;z�ٷ���6�~���>m܏��u���n�<z��f���|[�v!���΍�2���پA�z���K���o���������7�b5���mO���y�~����x�\��m[zXm������~�~�;km��ߛG�Îy'\x�#�[t��S��]�l������0���z--Μ�gB�,��͇F�O��ѹ��n���c��r�D�<,�?��!�I��S�񘘆���ۮs3�۽����l͇u7���|���f��ݻ{���}s�?�}Y齆y����?W���o�x=y��79m�g��zs��o�|g�{�O�ů���?��o�~��z��6l͇����l���m��F�0ٛ�������O����7���7�=�fަz�������;�w�4��-W_�ttn����mѯS}�>���97��x�����5�=�?��s�&�;	�_~�t8p	�Y�oF������IŞ���#z���܇O#[��z7y��o�߻��g~Y��N;�:v���[���fw�y���b�`��Ϸ��9zmܛ=����7l�<��l�=��n<zo���nϏ�k��{����u���x���8c��6x�����O��ܑN$'��G 