BZh91AY&SY���~�߀@q���"� ����bC~�z�   o�       (@      (                 @  l*�JJ�
((%JP%J RB��P���E(*�PJ
	(�"@�U*�J@)U%P
�,u{x���@
�)UJ ���PH� (*�J��( �EPU (Q@Q!J��BU�*QK��H���  �� ʀ 	R� �T5UT
0��@� 9 h +Q+@�� �(
��
�I*�!M/   ��Im��wm��Z6�L��Υ*�ն�ݶ��(K�v��enR�J6�+M���[eR����V��mN�^��S[e*��Þw�f��
[�(
E
)T$�  ��W��[J�nUΚҵFE��u��6��T���f����{ޅK��R�+z���h
�x�w��m�ڦ��g���*Ykxw���R�q�z�m���5���J�U (�R�o  wYޕv�i�m�^{J4�+�^�mjU-��h��J��Ъ�un)��h۪��n�� 5wR��N���[X�N��mV�4�E��F�*���*T@�J
�	R�  !�z�PڶԜ�sJj��\�ݶ��m��wC�)Weiip]յ4�m+t�uKVkMWtZ�R�AQ�Vu�iB��t��ڹ��4�ն�b�% 	 $�E"�  ��eSMi�Η)�m����	���)lv�t�SM-pg�Z�P����ٖ�[U�p�(SV�;(�F�iB�u)UZ�v���h��iU���JP�)J( )J  �,��l5�6�
��F��ewT�h43�7KcM�:��R娭3���PR���#��Q����5j*�#T����w��R�P
�)J
x   �z�(��R����0
3Q�U �Z���f+(J���*�v�nQ*�J�PR��jP]ڪ��% R�(     ؽH��Xzꊦ�U��B���*�J��5T`cU]5Dr�UP��P�@$�i1$wU@ 
UURQPP   ��:iC�V
��]�.��V3RHEX�T�UU+R�Es�Z$kt��TR�*j��ҥO�    �$ j�تT��  44  j�$�*�0  M0 E ��<�����1�ڠ���`���cP�~JJ��      ����=6��  4 z�D�SJb�SL��i�4 CC��~O��E����,m[����I�UR�گ.�T��N�+���������}��}��￰>�}U��m�ڶ��j�����%��(������q�Kyo�T�UEb���?��UUm��+�k���k
׎yuT���A�;�U� ��{���e��3m~3V�V�5�2�����my�]��e[̭���*�f��-o2ڽ��[��y��f��k^e��k^e��m�2��-_Y��k̶��k�[^e��k^f��k^f��6����*�e��U�͵�o2��k^e��U{ͼ͵�k^f��[^f��m�����m�U�/3my�o3ky���V��W�j�6��Z��3[�ڼͫ�ּ�י�y�יmy����y�W��U�Z�̵ͫy�W��y�י���-j�Y����j�ͭ_Y�Z���m��j��6���[[y�Z�̫[y�m[�o3j̭V�6շ��ռʭo3U��kZ�f���5�o2���5���m��UfVռ�Z���V�-j�e���m�o2ն�5��̵Uy�ߌ���f������*֯2�Z�-��2���5Z����mm�m���Z��-����U|孶�5j�3mm^e�k�[m�kU^f�ky��o2�^ej�-�3Z��ט�k̭y�W�Z�+^f��k^ek�ڼ�י��36י���יZ�6י��ʷ��y�k��f��m��k̭y�יmy�[̵��[̯�ּʷ������^�������	)�<���p`�fAY�!s�	�ܗ1�t����=�9��)��V]Kp=*�p��D*�s�Zy�Y�.F�{f�R�⊰<ݜ�[����:w>�,W����������u��W+��j��\#a��&�fZ㨓9ל�=�#+}ѥ�@�WL���z��]��������tw7Q	0;�7/-U��R�ӵ��e�׎3��Uu���of��^w{�\����X:E�]��u��]�3Nm<��U�y��m��^��D&��0��
:`�:E���M�pH�}�N�6�������� ���Ek�B ů�Ň�9���;F��pwoM�b�k��%�U�ـ�ٹ����|oDB���eL��ò��г�{���oN;F*���M�c�{�[7;D!֍�#:�Kf6{��)7s�=&��d0Y��{��L̷g,��<X���&s�^ݳtou�c��+�&
�ɜ
�v`[��i�>]����Q;%/;-�c{^�KG3��c�<����$Cf�'@sbH��g7P�L[3�v��Z�:B�a�H$�]ŲI�=�����{�$�ax���w�%��h��׀�1�+8=o:��S3�����D��-�'oA�{5�f(�R�k��#�6z�����y�	�D�4c�-� �eE����إ��{Onq@�ux��T�n�j�� )]H�h������k;nk>�Zp��d��jI��M��^�r�˒׶�qLV��<�9q���?n���[ޛ���wc�3`��jwm�r��1;9�p��8��4=�׹n�\���뫡BF�f�ǜ�V�t;��ܺ����wE�C��Ep����oc��Ww.�9	�~�5(O���Q�tC��M֌y���F��
��C�u�������E��J�.k:��c&$%�gd0�xyn��
e��|����"cz�Ǟ��80h�g^�\A�����=�=f��ËZ�)v� �W���X��������),�hX2����p`m���m��m�JZ7��h����)9�Em[��z�5	v-s:P��j��X�`e��t�wMXn+;�OM��b!�&�̲pw%���i<�S����{�m��3���F�@-F"2��z��@O���;ͬn ��7�p�S�'�����ץ��S��q�4��w6Z�u��`0��<H���S ��a�w�w���n�:��ŽF[�h�4aap�7�ӝ�HD��SBዧd;�	Y���Qw�-\��u^�e3z���ǻ��ֲmp���ԀG���o�NdzGn���ylk�$�Ջ{9�3�2�<`Ǎ��*s#l<�#�}���t(a�ә�v|�P,x"�`�en���;��RnŜ)Ox52���Ƀ`��5�Z�lM�v�{%����Xq>t�e`���6f9F�ɐY<zLX����5N٢v˴"k1i�U�� �������vl����8��9�;��\,��j[��sxIs���C�f�f���7VY�geĆ<���)�t�{'wQU
���ͪ�c{
�&)�x�Ǡ��,��Z�N�Y��� Z���	���	���y�#H�����ΰ�f�U�8�2vK7
kp�Æ+�Jm�e	^ӄHf����'n���nug�u������D���l�WQ�C��=��9�W��1U�5��0��z�n�0�`��X���� �ի���8s���w�.�)M�#�a�]�P����j,1�kx�"Ʌ��e����Zo5�������)5��ur��L��qY�a�n�)��#%S��qho;sAګ�]�5�z�s��1�򽻤kF���[wu%��Ӱf�7�Y��zAr�W���81V ��w�ݍ���Z�c"�1��;��ݠ����9��a�g2su��qe���w�h��`�v�q�\p0K�F��+���V!��6��r$�p��&��E
�K�k�u�N���3R�N�d��1ڦ4��阃�]Z��v���O������a����&M�f֞���3}כzbWp�go�^�^n	5Pp�)B�Tu���Bw��W��Lp�-�Lm�jS�����_nP2̂�wA�
��/�vJ��6�W�W�4Y��4t:��n4ծ�M�������uq���Y���sD퇚�vls�O��nS;cz��˕��*'*�ы�)�H�\qcӄ��G��#����za���<x�ώ�k�n��=CyA.���}}��·�Y���<�rŋ-�28q���d5�{��1j&[VK�Y8��Q8׍O��w7��V��2�`��F&a��+!�AH8ݹ�}�QGb&�i�?�ި�3p0��0��]���'gza�1�m]��C�����
P���5?R-B`�W�*�ǗmL�k�Z�Rӽ.ᵻ�t�4۝"�/��yH
��:������=� O���J_'��=��P:Ayo[j����Ҏ�=� '�.�4��tnײ���$=8��۸�4h��7@��;bs%qF#��U1��fI�-p�Ge�]J��
�P�ۖ$�ji֛j�Ы��{��b�(SzhB�GvL�qv�.��ާ6���k᝜�ʕ��C5��m8��#
k��-k�|���p���=�@��G�ya�&��⑕����X]��قL�<G4Jܛ�ι�e�&���E�w#���p�}�Bn@�	 �T�x��M��;f�fl���K���-�v�F����3Q&<8*� a��J�)��0��KJ�EHH�5��rD���1G`c�l@��<�L�aN>����x�^YB�(��pY�7��*�5�[zN���A�P<n����MpT�����ykcւ��SPl<���W$�eLE�cR����XR)ZBf�mH��G(+C�s��X���Y��!kC�;�������ã��J���pq�D�/�#���9x�8Y)��nه
(n��SU�����`�]��R�SU4s�ot�^��&,zvf�
�v6����L��ǵ��.��c���Ʌ����[1.�`�v:���U��F"��*�;�5k2b
o0��c�bw��~�~*�����7�b:�f>����z��<ͷ��ZRt���gN1������1��C
���^.ͳ�y��	�Qp[��b�+��[��J�r64��5��|޵QM��:.�6���cPd�椛q':/M$!�/j���u8��7s�	*d���,[ݨXiiopC�mh�uP�_Ϧ<�,G��.�t-��c�7w9۳NN���"ӜN�M�k�<�3ծ�)�q�T���׽�i�x�-�AZ��Nެ����ِge�b;��n�+�R] �m.	����i'c�wu�:������ԍ#�ULRF�V��ƌom;�/j�>���Yx�f��
��Tg���ڒVkmW7����x��]Z�V@�ݠT��e����Tں6�Xf��e��,w`�Q抈>am$��F驕��Nrя��V�no-�8�#�E��#�+���^�vjIB��G.��C��>®��ç"X�ʹaA��_\�p����.�*������N�T�0��L��9�l�B�_o�n�q:���80��5��{pi۸:�i�;����vhс8L]���A������j6�����P����3�A�.,�u��¬���pD��l7��z��0	��k��/�U���BR�Yw�v�Փ�b0�.��ܯ�њ��\�X�m���S�uAMɯ�VL����YP�B��:L��P6֗}ƣ.�h�~����v�����n5�6��ܙ5o�I�ɷܩ�z������{p�|�ʅPq׫��^�{�Շ����ѻ�:L��,�0T� _�i���p��	>h�D���;�w��ٴ=i�[�V.��|�w�����ֶz���׳�f��Mv2{wI��/Ǜx;�,n5�gsa�������h�ٛ���@:,1!ogr�#��� b�MĹ3
�xvmY�Z����ы���J�:G-:9 8���CSo)�"��y�� ��g4v�{{l_M������[!�5l�K8b#U8�s;�Ԁ��^nt��I=3Q٨G�G!R�;�O�׆��͑��%�=�y��rF(���w��D�,LS�XNI�d4� �
���M}�L�s[����:�8��1+����"�i��oaJwn�m* �UČ���eC@чyG8��r�vpUx��8�����(E�k��;X�gVmb�Op�>�&����� �:��k��u��A�7�������NU���@�<j0._�C���,�Q�$P���͹���ߵw� �*�u_�r|0mӋ�#h�����u-BٛB�A�)C-��L�
�11��eE�it��|���ߟA��=ɨ1Iۜ�1���jɒ��-�9E�=h"��I9k�
���/}�V:k8�rld}1�Z-B��u3��i��u�vrO���YD{�\u��ѝ�r�=N\#G>��{Nk�-�|�Ipn���HG����d�XL��7*NG�U�ݐ_�r��h2��!�v5�����L�q��TD���#�q�W;N���!�]}iV���"�jE��u�n�#�V��٧Xͪ��G2����M�J�w|\lX�ncS��+9��:��W���")��3��K�	8�L�����7S���
���&��<�"�v���{V\$Ӡ�n���t;a�q�?��9�Nwt�<8�U*�2v��@��0:5�����Zʮ̷N����\v��~�hm�#�F��d]��f��֮U��\���f��d�ivuTvjk#�v����CY�9cov�$�{��E��Q��u�Ov�r�Ңᎎ ])f��i�=U����r��+۷��>�����*�{���)Kh02�+�ᇎ2&'��p��s��N�ɂ���x&ۇm]9������D�O�"gw��|��2��3uc�Sok���ovmwW)kw��ɐ㫵��A�nٽ�������N�;rvjk9ƕ�E�ہ�f�R�_\����&v���ss�zNwnu2>h�v>�7�&�EP�m��Ez�f��n!���gg<�u��4+_���o,=�0b����y1c	��#�֗�tN�l�4�c�ۼ#f�@��i�X�,�r���K��8��j$1�7'L*%D{�Bp�r��xp`��p�Bz�
�c���o]����Ȏn�5���:�ӈ��֗������N��͜zt8�`Ͳ�����]5��g�SN��V�v�=�<I�S�&\`��V��V�ږ�r��nw��ӝk���ͨk|&]7-�.c<��.�Y�����\��W�h����<�pww4�F�.�N�Ȗ�����f�6��k��A�c���5=<����9�Sd�\�J[ˮw	�ZD�n4݉��M݌���}���Һ��X�	�Q�gq[���T���:��jٳ�r�@�y��y�Z/��@)�l���S�i݆�Z�G���{-w\�#&�ß$��gn�[���;�,�p��Om�*�V�yik"rr^�t�b48n3�ݗGs+\Y��zk@LHXv�=x\��|�3�j�ŋ�y�����Óg]���ȫoGW��V�Ή_g,@8���]�F�gg�؎�0M��q����:ٝ�qaLmBv�������"%��)
���0�L��X���b˥ۼ����X�����e�Oq4H;�Z��wPӪl)X!�{MM��3^;]�KN�*�M��"�����ǆI��c���j���q@t�^὜y3�{�̛����e�m�@x(K�Ӱק�Z�ٵ�2L��i-]���jHOg^�h�KJ�ȀX�h䃴ц��85jY6-Y6��	���d�$$��M9qTu���ŵ.p�+IJ���i�Ҏt���U��hα�%IL�,T.��Hw&�\��{6��A�Z�s��>g	,��]���vG+�:/�M욅��ab�N�{Uh�oy1.���C��6�ߔ[٩���{e�䱝7���Oe�t�L]x �ȃܿU�5$ya�͋�sg`�yC94wz��N,�qt;��I�/d�w��o���˚�(��"3����"�S�w���>o-^(��4��D^���Ss��:�QSzN���ݬ�\׽����S]��N>#*�H(�8�����;	��@��]����\��i*��V�ܸbx�������X�f�0�1
*����s������=M�[.t=�lӃ�P�Y䃼F]�N�,�x+�,�v��4�K�,q���x��;��J2F�S���릝�os��v��\����[n�i;Nvix�F&ؑ�gtnq�nG���{��EC3�P���s.��|x�m��(�L2	So�L�es풗����B��-��of�ۓGN��\���+��[F�DD�ã�/�%�À�p�L��d�zZ�G�/K��}I�.�ަS_�C�3ۗ^�޽f�V�lšJOORQ�G���`Τ�I�{��]�E��&#�����%`������<ѐ�}��;�ӻ3ߒ��#�[&Oi�|��`/2�����G�^f��D3pA�ǡL�{ts:n	���a���CO���4��qp�o���DrZ��"�D"i���5��kE=N��L��z�<iîx�p�k�g��Q>����j>;�t�s�#��n���=��{���yg�����~�<�9 ��͍�o�k��m��m��m�K����Xq���9�Ƿ��y޼{�&�[�ӽ�(4:�E�leq}�N�>B竎U�޾�I�����sck�&c�����v����+�г���z�:��|1PnKwa���sb��dEaڣW�x[� o,�Ǝ#	�[�3�f��p*2��n�n��.c͵�c6�HY8T��KR,CN�s�|:=>��o�'��>�
�@��g^
T=�4�ܶ�ŝT�9�SQK�wJ.�J(8��ӳn��������fΤ�:]+9.����26Ű�f��VCJTө�VU$����������suC�!q��J�[���<�s�I`U�m�)�����!�k6��EͪO�,R��P��51�-�㸻�8�����0�j�O���}��;���^ ���v��?1V͹?�Ӊ8�:���5\�����.%�j���N���p	&F�i�#�K�#���s:d`g9&��y�2�9�x��(���Jv�iI��)�͏yF��}\�| >Y�M^�r:���A<� �Ep�]�wI{��w/�n�7�օ��n�����6qG�p�nO�9A[�-i��*"&���Y�Vj�Ɍj�pRk�j��6���[
e�7�]���}��`(�׻&KGg���;�݀��Z'zy��(�����z[@�(@�{mߤe���g|C�gI�fz����ydf�쁶#q�po*�;��F�'V��;��=�ڙ���+��#Ek����p���N{F=��0����فd��wO{��=W���\-�Cp�w��u��,��o,���.�n�'im��ݯ�[q���o{��S�°-4+�@�F:zN��}��6g7t�܅s�H��ԋ��.�v�<����x<�g�ޯ��l�oX��l�<� 1~|ɕ��@?��������~����a�Q��t��#�{z�7��;ή ;7�RwJD5{j�U(�jVQ��Lpu~Ln�z$Ĕ��"���z�z��.��k�n��t�<��/�P�����,�w�Y�}4F�yoy�^����`���/v��`���xM*�I�n�R��f>mV�Ne7t�Z�V��~̤Y�����,��5��p�>���p{[�mr�i�;|B��^�s�3h@�h��=�b��r���f�>󉇇�l�~���-�',�ސ�nL�~[��k���j�-Z5F�e��ފo	���g*��@k�, fUET������i3'��^B��w�"y�?w�W�
]ݍ�7*ɺ3m�����ܦ�6r�9��3A޳o��-�;�9�zoe0�ٛ4x��R ��zk�ک�C��[�$��1U�e���T�,:Y��A���޹�����fu��W^�j��
����-�@���w8�Re�V���\�#wP���0�n�Н[W�����H�ٞ8�����tp|�:&�껀U���o���f��mR#ٸf7��)��6��o����t�u,�����79��'�t�O�R�z���� ���s�#�}ۚC���`^{xw�lHU1���Ƅ*Uqa���UU&�oX,�rZ���*\<�j������1_�uB������<O��]7���㹲�jo�Ek�B,�bе�b�t3�܃`��y
��=�w�S�U�e�E�:�g�G������6�-��Y�_SǙ��
�pj[WH#���*[���)�:@�[vr�L����u��p��#�"��l�GR��,p烑���=���	�����!�G�F��ˑ��f�i������\�d�_�����`���.&�Fk!�w�i�<���oo�gKv��ܙ^�8w�eS`8]��z0�p�$�_���I�"�L[w�������"�x�wx�nl7��7_^�ɵx�~[��,x�� � nH�s��j�3��Kp�߶��!w�uW��ɀ���>6�;�B�v	�m�|aM�׌��⳩y�;�x��=7�z&�����.�B��E��e�С�"�cn�����S��U�t�W�T�S����k$��uCfXT�~���@Ȁ���G�:��=����ta���޾B��_^��ӾP�wb+���n�������{9>Y��N�#Yr��tk5˩��Q1���kg���Waq���5�����d��/��<eG�\M�!����[�w5�;5���Cò��T/J>�0���o���}�{��������V�#e�p��w8+�M��n�%�8�������'�]�9�a�~�pf�OG�̣V�\�����"����ʞ���,Ơ�A��^.�/vh"YJ4:�b��)��t��y�D�j����Ǜ�|ϗ�$������ ��"ژ�	v'&�q�.`�Pi*�8����V��1�������t¶r����`��YT�����oOnw����lU7���߅!^&eޣ��o:{/g^�r��ɱ��\S���n�����ܦ�QyN�yO;�`�ɒ�!�$)\{��S�S�z���� ����+v@;^N��k�7v�y-ʸ�k�w�hw����wT�T�����]������5�O����s`�����R���a:n&�I	"�(�۝0�"��q\v�Q���`�x�MR��y��}�
�Ɍ��7�O���r����o�Q�&���v��ul��e�n/l�l�(< ��k���	������y�,��\<'{��ƻ�|7�}�ؙ�ƞq�r�{ܜ������>W������}�4/�G���՘�^�E��{�� �^�wI��=�(�sV��H��{ۻ��c�m6yO� WS��u�V���R��ւ�NB{�8�h�ԇ8+Y��"�:E�7bO���\b��Oz�77�9������Ȏ��I_jV��l�!�l�=���R����=R�ͬ�wFl��T�����a��� �k��Z����LZMڅ�B#j�X��~��Чh٦�,���J�sk͐J��3"�wj��x�ݝ5U�w��Gi�����(Z'���x\���Wfl����:�fNZ��kD�f$)i͉�K�2sF�b�&�W�N�A�6��.N����>������kr��	�zMX;��u��_t�xwg7o�M��2�)-�0�W�q��۳��f���-�M<�Ht�;+w�}��D���k3Тk�T�>��c�5���F�ߗxJ��~,�thb����������U}��ÄASo��s�z6��f)�W��23Z����Ѵ썄�jNM�g�s�������o,�۾m���|������Ͱ����;2g\nXn�ڳ��{��NRN�y��Y��7;��y�$�����^� x�75nm8��ό5��$<!���Б�O'��	W��Kkj��l�{�]-n����K�� ��?ku�8��v��V�������f��w�:x�@3WE��<f5f��b�L]��1�;Y���qb�D���ËKU���Kjolӆ�.�뀥�������&g(��V���{�����.�dq�b�o��m�`]����3ځ~��{�{���7�A$C���9����D=J�jbg^�{1������K1"�}��{�#|{�id^i⓵z�g��q��m@��;�N"z��ʢ���9�9ȫl��Ny����ce퓞x��l��c(ъ�{�[�i��B��κ���K����6޸]3��|6�_]�����|,�V��)(���z����ސ��g�^���･�-��]�#�KQ�1k��q���U�)�Ĭ�)���7���`���n�}4��������4p�ȅ��K��U=qL^]�Į���}���������wss�z"�C� gb	z�|�e�=��*������t��:�
�N�;7��x��v"RH�ͦL�*��p���H9u{&��;Ң��!Գ�S��{:�Jz�8Ct�h�GK���m���{<#�aBvLd,2J��	He�������'"��¼��"f^�Nf���}�?qZ������_��3�%���Iz����
�=ǚ7U)r��o��Ï�+}�x�>��5ޑ�F���WG$���.z}9�.({�n�1���&y����ߨ�h�ok��ǩ*$r��X��o/|v>����{Ӿ�(h)-,PWz�0���фIͻ���)��n�,�b���)a�{}�Y�kV]B�A��������n͜j�A�-9�>W��<WI�=֏zľ�çB�՛����ueJslb���Od&Y5KV�("��(��U�Є-�ø����;9{�t9.�;^3��㾐����\<�I��`�0s��[�ے����Q:�~<���ї]ο����=Ma�3�z�����O����t�^�	O��'�w�Jt?��m�����J��T����s�3$���o�f�e�V��s�;�f2��h��Á������<�Xi�.�ڊ��c��=x�^��-�����{M�{9�P��qƍBғ��D���/p�����Sz?
*~лm#��m6�3����ձ�e�s\,����c5��&F�+�+a�տ��1��������%�Ѽ��Y�����[�;��.x1d�{����O�{F�f����.\���$7�(RL/�'b��ͻ�@�ܮ����{r�>�r@Z/���=��_A�On�U��w�>4�L)���`���4BT�!�5j΅�̬y#��V�ֶ��6�.uI$�w�Ɇ(5Y#��-��R9�z�K�"g���vW	�$��,yBy�3��L=�ږ^����Z��i����ޚ���4�r�*��m-�։M0]��OF�Q��9��0a�8����Ԣj��r�-^�d�6T���qܩȨ���SԞ��]���wj���Z9����!l�'v�3����I|}h�q�uW�츻	�s�S���_[���z+��?0hFA�ٖU�n#��
��T\n�Șx��E��1���i�U�{�m�sn���<J���[���|��������u�o[/����k>�kp��.n�o��aS�b3<�t�#7`�o��a��zsؓ�����y4'O�>B��އ �xL���/-Z;_�����J���$�����]"�������53��?Uݑ';*��*1˂Oel�\�~0{%��RK�����$��<��Em=�3(����4-5��g=�A4��;�<�{��pa�r�D�ߘ��V��%�]��|+�0�e�p�"�|���]�U�^Yb��Ƶ�c���:F�F����^)��/���d�]��M������S�9H��bsr!7hlF��2�J�0m�a��`�O'�~���m&M~g�؁�Nd�`?/Pf]�"�7��Ѻ�B2ܝCӢ�"�*sKtR_�^�/���#������춋xK����q�ú��q��V�d�Aͅ����c�|=�qğ�,%���|���|�K	�C�O�/_+�x���Y׈���k*��%�Yvl�_v��3tcB) :t��\;���e�4����T�v�t~Y�|_��O{8�yi�e��g�|����tQa����?"��.LJ��eԴ�f�q�C�����2-�$x���l|zvPe'HO��]�����6=�hB�8�V���I�:�$g(��D��Q�Ve��9���)��b�U�q�O���}NxW���]������FD���}�k0��� t������;��"��A�/h��+=Jo۵�Y��W�����D{Ty.�@77����'x�e>ƫټz"��{5�֊��*��H�{ro���)u0���v���O�YPy�]��W�K�ͭ;�{�^�m9>��;���JZJg�9��"��QKbG=����~���^���^jv6�{��<��M��GC����G}7�ft��ϻ�����Vw�G��H�@q�E�=�t��t��J7��dtWc��>o|����(�Z)��FӖ*�/�����גd�}���p!�ޙ��7�L������Sm����+�oobj��x���7=�g�W�6#���	���4<NUѝ�[��͋�{�V�C�,�Ӈ=.Z&��۞2�y�bEt�A��q��'�3�W�ޔz��2��~��c3M��4r^����n]Z=����Չf�??x�N�$>�-���`V�T�K��H2�E��fȶ=�6�T|�W۽��3�*�O/y�9s��v^�W��H�z-f\�~�2�²��CKwB�FAy!]0�ۅ�4��0Oh�	�b;|����;��k��.ę��J�{�*W�q�ӳ_(�T�@�TjãP+~9{�)��_ُ�F�(&_b�*w�^�t�������0�/a�6�$�Cj�IQ�`�9H��<罅�ٺu�>�0cg�ʭ��!���c��V��rz�8���ݗ�1�.9����|�sV��^��	����Z��[��w��.��lKm�\�4'5�=R������Y6�,H���6�O���K�j�ok'N9���:��Q8����ܧe�=�Hd5y2�z
Ƈ�c���c�!���`M��qkB�����ݽ,o%4_��Ěs�wzў
�bo��4=����gQW�� �
mL�R�E�ٕ�tѥ���@���sJў�<�}ED���.�9�;���ެ[���t��ē��li��N,��e�ck����<������$��/ p�{�o>�zJ��{���p�bo�m���N�=�R��s�)-L=���,��M�����,�>�^���DY�i��4�G����"^�:^�i�����z����'ȏT :��h�#���O���K�k�__}-|7��x�����y���G����R ^�>���(�W�ǭ����s{o�Umm��o�_����\�?>��ǩ���""��������������?��7�J,f�TS�F���:���s�)���'�P�f�Z�Ue�ܯwl��6�����w���g�c9�:/�HI�<����xd�y�@%-�eA�Rn��Ӷ�q{.�ǵ���}�B�)s��#��e��W{�|��������b�1n�h�s�i}o�7@��R�Й�L��f�)b����݇�^/�{C{�=�*s��O�hݙ{��y޹2�[�Mz������O��f���,9�b@�^o�}��pv1������K���Ӹ^��m��{ޙ�����p=����Xb�֓;�j*�nA��>�n;��\��g#��2�I�k�`�Ws@���ǯ)���/F�Po�"��юaʙĽ__)'�yLs��Oi��c�p����W�B1����֐˞�ItT�w]#r�>�om����g�ԗ-�1��=�M����r��+��F�_T��f��M��Yr�(-��3�����>��s�)\s�q��9N+M�'���EN>�>�3LO���X�~��y�l�c���;�7HX�Ee�B�x�ɕ7"�bA�f�EЩ�0�v�Na����EL�W���Z�%��wʘ�d��nt.z��c!t7嵗O9t-
�w�����y��\5-a:g[!��3�+6`#��o���SA������I�]�v����%�z�gw<��5�0����Ӧ�ClQ��N���7
`�j�GI��[����!/E��^�Ӝ����7������������(��R ր�y{��ﯪ]`�?ow.�؎�-۫^�1�o��J�y���e�ͽ��F".��2Z]$lи���-ͧ،��5k{��,�N����ӈn��H)�t�r��%�U_���ea��Bwpu?u���h�#r����xb�o�1���Bc�<���q�\(B���c�ɚ��n�Y"b�N�)wڂ����}�4�_���\����>�/3����is}��9na�.�œ�n���z�ce��-u]�3��v#�IT-iXy�߼s���徛c"ѳ%&���{[���D8b�1��8g�6I�.��}�H�E��{.@�@elP�y�9òm��#y��䱹���/�Y�Um���ri5�F`����"�����,OPןi�Zf5e��h#Y��'�:��8d6c9�a�<��Go��o��|����uo�=�̏�kS�y-�=�5����R�R۳;:��!;�2�̌2V�������GM���/\���zF�o���S�|6�Dz�zP;흞��ݬ������87��^�r��>��/x"�%Nׅ�Ϛ��rj<��c��V����K�{l�Iy	7;hY�V�.�m������go�ȥ��=5��=�����r��}8��:O��؍k��o�|Z���q����vQ��<�\>�����gq���s8ìxcDm�k͹VaL=s
��=K�h*���q�|�EV��������ޓ�냲�tb�aIi�4k9~�sa�P^<#C���dgn����>�i�4��iR�Ñnkn`&̃R�;�$�s��_��t�|H�Ɍ���+��)6>z��Y!�5��݈��NSٺǳ���8B�.�a�[-g��f�k)���{ƙ`�O�4���*V��:L�(5��$ؤ A���*-\*�����Y)ݫ��0ң�j���X-��ѫ�D���ǉ��7$4��4����Pbٱ�8�;�N>>�w|�|������6%�i/Ĳ�4�����o�$G
l�Ra~�w����ilP��װ��A���0��З���l���j�>7m��|-e�>ޚS�x�ؔ6d���rj��LY��`�]�>ݼ��3��E�s_&�!��)������kY���l���j�<��z���u�E�sg_��o��{�2q���9h���gk�&I�}ڝ
�f���1��S2w+�����7��7�f°4�B]EB�W��rjEM�{/6��ض�z��vph�݊�N:��^h͛������w��@�1Wbc���6�������Z��|{9L��:�}ݧd�9�"e�&m��)�m)UX3��&�����.�Љ���O#nQ�-���=�3�}&y	徜� �款�$a���-�V���6t4$,��S^xd�P�f����o�$�4[�y�xs{�!zH=w�"�.���v�Y�.G��Xs�0fw�%�m�0��lÅْ�s�||���U;鹷�GݭO&�M>�y�3{J�b��j�΂�Zu�K^�Z���D�#m҉��*QľAg<<��G4��R��v���3�C�ଁ�y!�����ck�/n��=�E���Jg@]=���W.o=��a�z�̗���Ȝ���y&
������W������Ӥ2��>���C)�m��,�ݽ��zt�n��S�ﯻ�i���I�x�{����t�u0�t��!sT����/=���~�֖@;Z��;�^v��n-�R>��*��_gKՃӖA������%}�w&-�uku�h�J^Sa�58O�x}�Q,^���᷶�c���j�������2a�;|fB�5S[�d�p�J��<�9V{ږ(�W�e�hQZ�J��(Q�����UđN��cy�������>��>Y���!�[K��o$��nL�+�\�ݺ�&�/d�RڰP{j�UM��(��%qo�T�]��:�NI�Lq��|{���s�Ę+�����lWz<\H:�F/�w-�a�t��s�O�V&_^օ���>�wY|D��^����3g�M��<�go+7��p��-b�9&��
������,%&ԓ�T��D�I����pb&�����u���'ګuFp�+c)kȽ�Ss��TA{�W?_)3$1<������Uo�}�yk[�{:�g]�ɱ��w��*�:�gn�A�3E�� u�D7�J6��<*�ϗ��ܾL��;t�Anxl�͒���˕3SrL0�t+6-��Wki6 Huw/\nk^ޒ?x�������ΒC����D��/G�s����x_o�QH�,߹�(�����N���}��ǎ4<�S���p�k�
��<0�vvB�:Ϗ
�v��y��v��m�5��図�'\�UO%U��orS�.���J[��T�+t<�CP�w�0��=��K�12X-��E
X�B(�{�9����J����Yt�j�Qe�+I��6A�d��6�ji��i)��{�x}}�����pS��q�<��f���Q� OHG��n�s�L�ޘ|��g��<�x 4��ֽ�F��W�g&��ݙ�.UͲ3�C�8ݏ���\{ޘ������^�^�3ruS���i�^��Xׁ߇-�=
kY0{�fz3޾Ȳ���b�HɁT^���-F3H��-����վ�I=�1N)�h������I��p,�q�����nB��\E�u���`�dK���˩��5d����l�i�P�r�N��A3iL��D@�]��p�<��������k3��N�*d��b�\Lz�j�d,�ߜ<�R�üV�{�X{��>f5s��3�XO����@�W9xzy�<��t����|W�� g����>�t�p�U�3��˯07ǘ��*�4M�[���H<4�����q}B�yz/[zu����ܩ�JR����b����.Wx��$>��ţ l�c�k�=}-X��mv���s�@re�3����ï^S/�hC�NXF��,�ѻ}�l�>��	^	phN/|}�{�NM*ׅ<)^��}����Z)�;|;]��B�浪n�g��OV-���G�LD�!mY���O,}JE��lX�Ǽ�s~Cv�����v� �<�<�݊�b��:B׶G�t���,X8��ݜw	�B{��DPq��n5��t^΍�a���˺h�e�.�U�
3"�ô�=`�l6���A
܈��"��a�Hu*iۘ;��ὸmי�V���J����I����p�`@礃;'�n����/e����y�ރO��.Oo��эJ�Q�%\53�n1�:�yeV�E�䍽3�n�KK��a��^�ͣ�l~�vM����m�l��vB3`�Ī���E{qo��5)&>�^��:��P���H�,,�9D��9�Ǹ�{P}˭��9�g-M!�g��L��uDp*"-޸��7G���7X��FמfS�^�݋��F�
[�ܞ��,Hw�Zߊ=4�,����>��h���*a�p���/����&�;�l۳�n0\�G�ӕ��ٌ�F�/��yo�B�>�bJ���z�ｎM���x߷�_xi����5^/����j{�P�q��J_�'��d��*�;s��ū��0�=9���œ�G+[<Ny�x��]��/����C����v]�A˨r���Q4lP�Pwx��>��{����]=����L�Сd��-�
�)ժŇD;�3c�8�<{�]{%�='�e-�.�,gV��N����y!�fC��w�����w,Xg���k��<�����|�~9Q���^�9��u�^�Jl�}~�(��Z��Ԍ���u�3׭(�3�Ɲ��~���S�1�z~gJɉ�x2V��cMן�z&.�ل�b�W��;�+ȝE������"cjci�Io=�a�7bV��,��5b�]�J�����=�,.�c�{8�����=Q��7A;^����:�{��_�.����p�w�5Q�>�z�"lS|��w'a�n	�4y��٩������;W�g>@��4r�6=���1$˅��8I�Z�%��=݇Tf�8��{����P�Mj+�AO�rM~�3q&ݧ�E�)�����/1�.�Y��\R}� R�3fOgV��n�>�ФI��06.�N�S��:��H��t�,�_eb�4��xP�kT�.��?��<�w=޷��wsm��(��=�*,�9��F�WC��4ѽ�p7�/O�:r��n�C��م)K�M��2�[!rfkZ̺���c谼�ތ��˴Ar��������O���e�{�r������z_z����ջ�s_Y%R9iE���d=���7
Y��AN�h*&8�[�ù�&���}�};s�t��àږ�����8�;�y�tM���1�^��>Oڨ���ĈI�:"8}�v?��&����!͒�|1!���=�:@u�ҽ�M��Ow�ך�1,���S�r��=�vc�=>�#��,���fmKs`Þ狠AIw@�t�7�+�p�i�n7�����^Ae>v/g�̷�l�����Us����Mg��O��uz�ϴ��x*����է�[k�W=> `�ݾ�A����TжDQ"��Z�����������m&L�ת&�ƤΊ�w���U������P�F)S����}�\�z{��y���L�/��.'�W���z?/\>#�?HI��׆m�-�/��um�~ �S77�U��'���Y��x\1x D�nY(�z�o1�F�w���{��taט-��p���b�r�����U��˫٩�x���ky�*�1�B�N\j�������RQ�ч�߳ڃ�pf�>Q���Q�<(ƈ��$+��� �l���=���9�V, k^�}��,�=6>��֬z���`DM;��ۋ�f�����L�W�嚚���i��܋e���di�����"*�I�5��L�"�S�[^���g�oDeBЌ-��x�nԎ����Ӿ��X�����'^�[�/ P~uYm�y�i-��� ����ݝPf���w4K�4����ų�ݾc�����q��Q�#�u"��4��w�=��gzN94*h6�D\2a����j>j��_T8��&#\#4('f�zkRKEn��5�)�x8�$�f�DݬɑZ��m='L捄wdIə���䪖jg
��켴>8Ś2�ux��|����}�oQp���}���[�N�JD�l�D�Tڈ��]��d6aTe|v#k31��b[�^:�U����::	Wv=�W��SvЈTf-�%Z�t&�	��=ro����`��3ٺ��X��_)p:f�WC�n�D����&�Y�n�Ab����D���;޾`����8�d�2��𡢤�9����1c$4	���4����&��@�e���L��&R��6%ތZb){��!�˅S��S�����������5z���׸�<x���9�I�����sp!��{�mTv�H]>xb��Tnh ���#K��\з��ne]:���];�E�	5/tһ���C~�e�i~��%��Ը��U����� �mCh+ώT��sO������s�-1�Q��LqC�_nÝ�=����*�^���J[����{޻|,��o=�1�M�h��p
�ַFg�|h�+���x=gN)�f�5�g�ћ������)����M0�K|L��(�f
TM�L:Ҏ��k>�ͯY�W�+�~�9	Pe�X|n�
E�ےo�߯l�x_q��4����q:�U.�෶/MyB��ӕ���$h f�8�žy������� q���#�E����e�{H��{Q�%�ݛzzWu.��\֮X���FKx���6�?��X�;��s�L@���.1��0�����}n޺3��Z�[@�.�>/c)�����C��`�֊m��©���`�����o`��׽��[;�뤛�߽�� b�(��{zkY�ԉNčB�c�a�f�m�КԟQGy��i������|1oЎ1�T�8�9���c�^�!0m�_a&Q�o���}عv*=l 鎠4&� ��1J��a8�)�+4G�e�*j�\�9�ta��`�DK���~�ǀ;�|EɆ7�-��Mɰ���&�Դ:�{7yuo����|>����]lA���û���������ͳf͛z�^�_��Ͽq��k��l%�����(@���Ađ!0S	 ia� χ�ʎ'²L`H"�/ E	�su'�O��yQ�`ٽ�����4�aǊEi�dao-�HVQ�ب�4���Tf�i��@�ĖtBW�m:URf�iw��O�_?f���t�n��nK{nX�ͳ���sv_?�z�V�"�8��aQ�ٵq�u�t٬�-NY���Q["����l�c1<�[Ft���A����n������5h������p��U���]�禂Ny^�}�����k��UI��#v5�Wu�l��
�L�;�YG2AA�a��/�c�=HN�/�=%N*��4N���h�'��5oh{��G���x4��2Qh�rl��`�x�mE�Cw8����)Ln��!,Mۉ�Qg�����4��'��u/��cb�������s�s��X�.x�`��ݝ��ޓ=�Jf�����c�e=��%�sV�"��_��w��ߙ�V	�iѝ|.z@;L�ssG*}��v�G���.��]�����Ě���1��/ya���xx������p)���K�ݲɋ���{������2wy���c(����J�	s��bf�Xf���؈��\�G��c�c��u0����ӆ�o��\���|r��NoC�pOLN�>��Gxo�xf�~�]g�gVD��Q��*�C��dX�hļ��^���p�q�Ԋj�Y��]��9ӹ؄���t�7v�\�@��<)�D��HfQ` ��h ?[���6�d�(��1A�ǈq$,����`F�m��4Z!���$0�����0 ~8L1)����pQ�C���	�>�w�{�쯱Ig�|����I3{]�p�"���;�1At�bR��LF���$�n�B��FJ�t�]��\�9��1I�rW:(KM�p���(�R�N�v)�����U˔��s��C����1Lut��s��n1S7wI�9]s������L���+�"i,��q.rs�������C�$�
f,��;���wDE��2�Lȇw	&(�Df����ņ��� ��h"��D�A	��Ԇ ��ŘȬ@,$Ģ5	����Lh҅&�d	%`�b��K2) !��("�$"m&�ř�U|o~���Jp�IL�u�q T�S��q���\��|�Lx��C�A+���rVl��Q-���;�P�{���F���㽵��zxHLf�+E|��_%K�����f�7�U�(��+��n��L��Xw�mblŕ�5/�x��d�Uʬ왂m짊����*�X�R�F��<;Wwv:|:��i�������Qb�����(��:t��q��z���pt�X�V���j��z�k��&wk��;]�BlOp۩c�b�2络O&窯ٜ컒�$!=nR��wWA�2�"�B{��L;�+�E�v����jT.���gY���xm��6�ἡX[�미pڔ9J�4����N[3��5�e��U�g������8*T	f��@�{��¢�5���X+'i�}O�5��O���:�;�۪�����*�(qy`��Q��E}� ȁ���R��	���r�>o+b����V:��r�z�[;���8��>��`�}���p.�θ,�w�P�#nn���<vH�X����<��p��w��B~���x����N�u{��P�n_�U�le�j��@�tnw��۴-��y���Ѩp���M��y�;��کn�1&��۴g'Y5	f��T��Tw8���M��L��LJ�^�:����q���+L��2�Fn��n��S|��,�e��uA�n�ϝ��8;CLOc��ݎ����V.�.EY��[���D�4r����p�~�8�FW��[1�puC����I+�C`^�V6��;-��Q�Š�@i���o��aΰ�$�m�y*^�&���#yu�R�s�s	T�ښ��8K�<:������}��1�+l�۔sXv�;������%Y܀�TS���^w_+��z�7�Y�}6q�o8cͰ2�^o��L��D��w
�cg�SÄ�[�M+m빬��;O�����قVm���Ƞ���5=׺�=��Y-]�tNޞ�J�/y�i>��<=n�|� �"7'����1�����&�沴㐕��<>��E�w8�}�m���[��n���l�\M8����{k)�wBA2���u����巙%��3�#n��(�\>���GI�i҉�$�w�z-@s0� �
� �B�i��Vx�`����:>�2U�
�`�T}�؛O�Iӆ+�f ˁ}2#緳���Օ 4HyM~a{��</��H����Tcq�)]�6�8�n�����Mj�x�����|�9v���p���5U�0��{J��b3�@�%_I���K-f�9�_9�.P�s����u+�cRo�����x��'�U��rr�s����f��\\\Xw"T)�J���^ʺg ?G�.	����b�#jyÕu���w�Y@�i7Z�>{щ8Gs����
V!W��(��s�:�쓡Օ�z���2�#�'+{�����>�m�>B���B��B���KuO18|P�M���չH���T5���jh21�ʲ^J�&h���Xi�}�lv��8��]���)f�`���ݼ/�neE��~�9�w�t�sp,ɛ�@�H�j�#f3�W������+��ym_2[�[�5��$�b��ۇ�+����wF�v�W����0��L�����HΜ���K�T���b�f�!:W02��~�U�H�v�J���?l篿Yz�f�yiC��лJ�8�R*5lmw#�gB��j��ޝbf�TCs7!���ك�r�f�k�L�v��!�M�̔V�ka��L`�������x�!`v樺�G���e�Rz�F�`��am+����y&�B+��������X5M���<g�k!ƮZz[ἱ,�F�9�vm�y+66��r�G�Q�س���g1p��"���0�t���4�J��YY�}��nJ�mn8{0Li����)@�jw�p"��1�mZ0��f��~���X��6y�M�xnt<�l�8p��{���qL�aQ_6�g,Efr��Z>SwHm��-������������j����J��O-���S�p�c�ɭ��5����k�8�g�۰��~;P4��'���Z��QI�[��������O�O��ԝ�4e�ad	/�$_@+F�"VE$���n�]a^u.6��>���}��Ng��߰.�8!���E᜞������������z�����5�<�W�Em��_�N5����lkƹV哩<�d��)<�v�$���� ��g��8���x�Nr��V`o��~9�8NN^�v��}p_NR%��_�Oa���4r{]�Mdv�X�>�4�*h�Y��-IM��JΚ�I�ԭ�j	H��=��ڨ���A�h�Z�#��+���3�D��qÄ[�ձ��T-z�KwLJpMtP���5@����c��2�'��1�QL�Q#�5��F�s$$f�P��LLN�z�-�-L�kGRrXv3�ܽ"4:�8c�Uw�j��1ƪrL�jΦ,���-�*�m,A<3֬}��īq:�Sp"w��iį�앾��v�՜n���3ç�m���++*嚃��iú)��1ï��(�8���)Iy$~Z�b��a���ADj�F��y�d�&%����p���XSû���ՎoI��
n���S��<��|'�m����;���P��N���3��,��=Vt�1��M�QE4�A�q�<N�A����Ja�5���z�QZp�����s�mus�
m�(H5o㚄04K+m��0�3t���e��u,��4�]�N��PĎ{�c��t�~�XX��-Z=�n/}���X6��}�X��րj;��oO.A4{��i�R�8�LFo����(�qL{k��{��rh;�R��������n�O8����yz���[���{w��m�ZTl���}�w�*����͞p�T`��*:�J��8�B
��!t�N]����\�3�u��+���P�<�Ioxf���p��[8`�@@�J�����\��7v�
&6�I����V�o���r?@�
$0�H=S�v���_s�5;���xhU����^CP�k/�m+GC��C��|q �u4uɎKL��!u���tD�o[�e�F�9��β-�X!�TH@φ��ia��W���W��mW'��d.}��V�B�Wș�|2���_�S08:�ኜ����Ɖ�|��ll���K7;AJ��
���}�/���9֫%
==#���cl�<#�Rȱ�Cޝ��[�Tm�3ûs��b�e�˻qE�D���Mf�W9���F��3������F��;p.���! �vx!idA��i�J8t�o���r�2��GQ�r�v�;��㪧b�n4���a�:ڌ!*��ZJv.�Z3���Tv���E�"�����3r5)���pض�2�6�+�U�w����2͑��\ӽ�p���j*M����xʧ���Y�2�]������+�V"��(���vN��0�2Z���aq���JŪ��'�o�B�Ƞw�*Ww)�<�2��}�H�J4�p�Ԣ{� ���v>� �1�<��a:A3P�30��=�AIcxo���P.���s�
m��Xc���U�kr�dJSũA��th��U�(+Ֆ��,|��g.����ww�l��jw�S��h;���������P�"Mr�K-`��3�K��.{��w'jԍ�V�x14���}�PŰU	@��R��)ۆ���E��]��9Ě��e����������������)'R9Y(�N�P��RU�}��Q�S��	��V�ꀸs�_;��C���#��6�,�ƽ�'�.�9�s��ZT��H��mJ�܆u�*`��SB������=&�y}~��v~/�E��eW�Ox����#&��s5V�B��.�
sW׭Գ�n�=�&�Bٺ}���+�ųWo����N��9�T�<C�>���<�|//@�	������P�$6�!I		Ԯ�ʜ׸j˴쉎ѹ_Mv�
%v���UXNذ���mK"��M�7���E���Y̚Ʉ8L�1D���l����"���8--B�B�޶�;�)񻽾�g;{?O[Ͱ�%Y��T8l���U� �7��=t��b�����M��E��X�b�ɕ=q8�ЕN�Ԑ�6�槷l���֛��|��_#ͺ��ɟ��S��;�ǲ8R����Q���7��V��8����_u:<sly=y�s�A8G�G.R�l<��q��R��!\��{����gg[�τ���K�h`�_.�M*N���z��LT�:�(bqE�wo�y�B�Z�e�-ʪ�1uY��V�m���X���#g�l�~� ��J𨡆Ү[�p�m����y�j9�)U���6�*��Í},%t��S�k���G�.p��n�w;t�j�%]$Ud��n�tW,�"�����1����/mC��zr�.q����:��ݚ_�%��1�����Sٜ,�M�y
NE�+L�&��
s4B��+1�!�Qw)��hE��5
�$$����i^���r50]�3c�;z.eQ$�q�}3WesE͌��Y�����<��L	[P5}�����[f���xTj���y��m����jN���u�b����Z�DC������\E �����Z$j���{�dr㏛�����Xx!��7ӓ����/�>C�<h�7��}��+�]��t�5:Gi�����q=�)�*&����8tI���qelwv�J��.˦$J��Eu�ӝG7���f%�!���SH��#��ps�'���z��;�tFiX�om'���[���#9M��#C�ᎄ���f���:��7ԁ����{��
�`%�_ȑ����%X��U'��A5Q�w��Ivg���"u�6�U��K�c<:���x5�Y�^�K�ը9�3���2�"�L!�>lQ�2�[�Q������޾��(�}͏.C�ʍ�TO�/ψ~�={6h�l�/N���}��/z��OQ��*Z0^]N�9&�chcy{f
uG�x����1��:�wwVnkR�9���2���F��)C�����.l�͈�͵�jj���Ԉ�D��v7*C�Q� I�{�"�u���±�s��g���w
��\�O���f�5�ʎ�-T�岨�y�Ni9,�ؚc�n��:�����X^�06�\����Z�e����S`;�\W�fO_���J]b����r������]��+L�"�{���.�}���y�|�������6o0G�{��ꂵW,�
��S��³鳥l�ŋ��l#aT`�����B'�_u�©��F��O�F�/��v5��O���:�ؕ��x~���:�I,�Fam�d��}P�DQ��I�Gv.=��vw��;�M��+Kjk(���=a}lO�H=S�v����9���O��Ų�S�cSky��·<�AđΦ���.�\�WA�x|�#s�F�����}�E9ߑ�`�J�x9#Z�}�~�=��O������^�W����{}�n�Td2����L^I,��
2���V����t��1��b��T�B�EYL�
5�W������֌�ޚDOW聎��O{�Fߓ|tԽ���콖�9z�:��.XPaF�S�+(J�a��h���ǀ-a�x V&�օ.�@����.��$oZ�g�pn���/��E���z�9[���GE:gg�ש��(�㫦+���yW�x��:��sOT9�T�=��j��bi��^x剢V�9��K:2��t��Vڛ�q����9��t���<{<7=�<3�ܒx�g�
=�RG��~o{q�s�g݆%ԟ=�g^ӎϦ�r�êg(u7��Ր�n�>���ۛ��g3}�����]��- ,���Fۘ��+����m|�v����Ïצ��&mߒ���x�Y�@���X�jz�Rr��	�t���>�W�-5qxV��'��![�\_Ys���sWȑt�|Πa����Dr�23t�����e�v��?wk��SV.�Dx�9���c/|�gΩ=;_g�Q�~��<�'����o6��Y$�\G��+�{�ș��E ���2����뽓�t^ʂ7tht&r��מ� �rr{7L<����(�C�xys���r�ӑ�����d���O��}�[�#�K�؄�bo��/�b٘]^֘*mmc�X�F6��d=�&e޹�{�~b3����v�=8����]��!	��P��V	�cߙ!2�ؼ�am}�ڽ�@s�|�,5^������ċ|��ճ�$����)�p�J��'.b�֜Al{�\��qd�5��*��E<eBF�],F�B� ��#�7-�c��(�h�=�Ы_[�l=�;�ۧsv�W��$�N�N��T]�	9AU2�uQ��SW-Yzw|1A� ����ի�t�����y�b%�����5��2�c��Tr����;�:7������~��݇k�Z���3���aܚ�{��|�-���Z=n��<��T�iָv�8�_{�?�U�nw+�	\Mto���^Y��JvM�y�T}fO&�����m�n���4;�T;�q�:�V��v$��V��T�%�Hf��ݪ�)��1�hC�tn0iƕrF���i��u����'PΏ��G����^a�\�x<�o:�^w5|=����=o� �<v�]�8�X���Z�����Y>9D����u��=Mgy<<�5�{�XgN���1�z2�,mS0�ب�-<���sƧ�ўUn]�I����+!\N�f3�*�0�隷�]�[�`9�ZK���SUj6SU	�/D��͆j]u%��~�5�x���}��׳S��Lڻlu�9|x�Uᩇ�=�|ߖ�*#�=��NY�u�c���|�=���bNQ*���#2΂V�6���Th0$�x<�%��}�w=Wd��jr|����<<s��w����Z��b+T�Z�����*Э~�Oc�N��"�r^����5U%R���`����߯�{�������� K2�I�����)DI�Ĕ��&"&"�&IQ�̵&,4��1F"$A�)631�L� وe(bZK$�H�JH%#!J���6"�TDe#S2lII����%�b(�آ�v"����h�.����΄�� �K��@I�d3����LP���.D��h(��qWW.���]��ʹQ������9��uݓ���z�p�pfw\��r��IG�\�wr9��$�NlE��gwM	�˕�w]n���\��۝3wG9H�,k����7Ǘ�>��O�d-���Á�N}��u�'EOpĖ�t�g{Sl�o-Aȑ���3�,;� ������9��֭ټ&bP�=�I�D�M��Z������]�ZJ�-���%�|�Ã�݆/�įY�.�'��Q�C-Q[~���՝�>��ls��C�]/��T�֫�;�lto�\E��P7�`i���y��@;�����zY�`N.����W:�GLzS����\�m.��l����9��ߣ>��Du�>��� AV�_��D�}��-���W�'�תp�Jm���I`$-��-��DwK�@� S���y������X���<��b�ߑ�D(�<��}�T�φ�lҜ��L���u�p��؝=A�}xTd�A�Ǖ�Ӈ��0ꐏ���S����3,�*�+�z��5�rmD��<�r���4ܜ�ίۋ��HP�z�)��-�UV�o;ɬq���l�O�j^|h|CV��{��^�˸o�A�~Cߢ~��� ���_��y\@�cU���ݷ$*�r���ŀy�c F�H���M�R�ʆ�1]4Ep�_�C	̸Q���"#��61N�;��T����ֹ/�C��܁�g1:�ޯJ���(��9�c�����&��^����L dmu\3;gw��>��uS��R�}?1�$g���������9�l�rFȨ.���6����x�g�:���h�r��r��ҕ����>W@�y�K��kJJ�����]����t�����l�xaC�dTC��E+h�T1��L�%���.`�5*��N�
:ɧp�c'[{Z�.N���>�뷥��s��u?�|�P�(c�:E�mE���!f'���pd|a�c!�}]�#��`L��;�i��	��G9w6�u��Uvr51�d`7�|���ck)3���y��9/���j�W��!WC�h��_ec���G�P����K�����nGR����r����u��!�GG�Ra�j�Ox�H���B�j�N(/'6�J��%��c2;���.ܦbF\y�����!F&(1��Xu�}��(����7���υ�
�Lg�\oҡ)��� �݄k��]��c��/ʇ폽���lk�K�!�l.۾.>�����ޑ�����}1&�ꄅP��F{۩�5��}���wQ{&7Ӂ����V2d���g߅'kc�:/6�ǡ*� &{x��C�{�}�j�g��"G�Ƙ��N��u�;��U����
a%rq�I�kxS�n�b�����s%T\�W�ֲ{��χo��Y��U1�Lj�a�?P�X�Ήϕ�@CK-�KWa'�$�搰e.gc�����C�9
��1���z��j�}:]c���{��Q��ϞVœ[R���`�CGx\�v���y#�	�T
��J�#f�Io0�W-��$h��*�[�`�p�ϑl?������ׁÕe�˻$��������(�t�+mĠ�	�7��3n�`˵oi��֪�OI���i.&S^�9g��b'����:{2`�2�۱�ٰ9+�k�f���q�ؠ�(9g-2�ȯ�CA�	kv�S�5nN��Lc7�!U[��7�z������/��/��j�#�YQ�GV�����0q���e���B7�_�U�X�? ������9=��6w�")�<��_û���Π!*��8{�xpV_���[�4j�*S��)���2�u�ks��4}��>�`��%-D��b�g˯� bL�B�Âi�h9��?->���Ą�4����>���y�M��f�ٚ��ڛ�w>���G�1tʑ��!q�ꛊ��o��G���q�6 ͗���<��f]�H�M⁏��,߱�@q�&�R����~�J9ڨ旋�tz�9�8ѱb����l�+'�׿K���6�S���򒑁�0��Jg����>+��m@^Bg<�}!���	��0�<qG��y7�h�o��LY��>|.�"x#�W��aw��{����j��A\�:L0kx&��L�ɯT�r�.`���(�f�P7�F/]Y��5M{Z��η����3�]�}��@�B
�BӤ��ņ�N?*"<�/P�o�푎�a�s20�{�����	ens�J�3���^Z��O���.(��i����2��j�l{���x�P}����EV�|+���
]턏u�����ê�y�Le츥WԝUZ�kهhD-�F-�Q��ڪY0�ӳZ0��{S;G\�e�f�h���w��j����D�/W���W�HN�p=��hm��إ��`J����^V�N�}J����ϸ��k�'�^P�cG�9���j����cY�^���2�]X�@G���\�R���_�	�,�5�$��Ν��F=̸�`%�fuu1��bLt�?q��q󘹉�e��g��%�ʔ�dM��� ؋����/p����Ԍv<��� I3���U��sU���O�4o\�j(���)(�i 8�B�z�7��ٌ4Ÿ�?lƸ"w�H�jF���4ei� ¢�cW^�@��M�ĪI�!ԝ�pUΘh��4^��8v�����#ק��z�����K17���ϧ��Щݺs�=,kNb��@f9B��kw�z�Ր���+����b�5c��^S�\�J_���Y�r`⣒�>��	�	�BP����ˇ8��\)B�@���1o�9��5<585ֹ1�:E��L�ϹA
�U!��'��)��jj�;rx)������5�kg��^H�������<U9���z�3Gܢ.�Q��'�:�ּ\zH82&A����}���]_ǕqM:��G�f���ra$f�����.�݆�ƪ�2C����3N17Tޕ��$�j½9��� J����y{Ҙ�Mɝ�D�1�'(Z�p�7[��Z�R\8DݦL��Y��C��}��>��}��[��}�8b��vD�H��Q��2>�"_I�����(�{�7����`>��7Q�u�.�fka�+����ᆺ;n�u�%�v D��5;#k���F�M�a���!�{�bVr<�	F��Y�&�yWղ�Wf0.����v�s�tr�Q��S˴Z}@T���Fc�v�,��1/��sr�F��_�m);�*�МHP>*o�.��>3���W������,�g_��߄je��+��}k�E��J~K+�/��<���8�b�K*,)���VT�����<0�n�'���b^1>Q��=.N���Zgx�����=�D^o�<����}H#�r�C`�a��Ů��hj}��u�j�۫W{�b��ߙ�> �n.��i�:�b�f�]���{mۂ��@�EC���n��#Ɵ��$�N{ӟ͚X�2g��h���m}d;�@l����H�2�<Ѳ,�z�gz��.���:y���yWF=��i�%�6���I�s
qRHx#����s�cO8.�V[T�ƣ���{��������R���oF�����Vp�\�B���-�//��Mw�Xw�dH�tX�s�B�^�۬�2|�yn���kˬw�K\��ͩ��]U�MN�O%�Q����/h���Y��+MڛZ����A�uv���ޜ�OW���T� �.�9Y#�ԫ��o��>M�z�ubX�,*ݹܙ��m�����h^j5FO���|��׼��o��R�LG�\�f�a4��-ϕU��������klOe��I�>�aC���;��3���]w��:�X�n!e��>��V�E��7*fܨ����Şx`�ή��&kw���o�(|ȣ�]��ni#���8�_Ypx���G����j���r\��del�:}��Q��t���a�j�Z6$�>����X�@Ⱥ�fi�\4�(���-H=ئ�I�St��%7�m�n�b��W�>Ǟ���H: I3b���pa�g�r���<���=�O�v�<}N>qП+[9�����ME��M� ƅ�|_B�@���&&#K3�γ�Q�g#V�tԖ����un>!WC��ѿ����3�'�~����� k-znhV��,��oB�\(5.q�@@l�Y�
�p� V�t���ӊ�'X�>rFˀ=7�ʯ
�Ĺ�h�c]�d{�5LS���WKҶ��CzN3c���*�LbW�y��Yw��w���"|��1�4��Лk���hA��]���K�Ѻoy�v�`9����Y�P(�(gV��̃�U��<Ebr�g��6*~V��:��ӝq\��.M7;���%�8/�Vƒ/r+]<�����Ph%��f��q�[�º�0��9�nC��)�.���M�n=dc�(��.r�L�^\���NA�"���>�������w'r���rs�Va�������f��q�byM��ҡ�ˠ85eI�U獿���Č.�X�����{o�e!!�S���W�9���.l�L�Z_�7 >����95�#�JY+�W����;�Y��4����(?P����D�S�1����� _g���f����%,�F1�EY�s�_^)2/�Î��$T�>��9o��h<�#>}�����郂�n�>�9��^���˫�j)�5�0���y�w#6��9na�ps�U[��&�k���Js�����t"/ĕ�Ne�m{nGK����lS��|�8��@G�!-l�B��&�9���,x��ض�k?{�ԯ�H�[��`͌��0V�Q�S�L�f�_Pa�FC-�h������>Cc��	�q��||T�rқ��a�~S@Ǚ,.�6�1G�±:	<�R�A�@[��.�̼����H�	��)�opgyہdj�f�5�6�("�&�����T�]FϏZ��zx�5kr+j$�y�����t8-VZ-n|5h�k�7AO��u�GE���0�0��k򲮙ٌh���1��T진TAوX�
�KK<�j�]�-���;tZ����8�˻�M��.����x �I�bT���}�����S������r3�h�|9��`!x��Vd�" $t�<���Hq��p{=t�8G�B����:"[�����x{�-�4�:k�A��?h��p%É&��`�g��`ף�v� �m��t����%?됹�(�8Q�[{*$q�:&]��@�
�#�*1"<�o��0��(�ϼ��_-�n��Ow&��%��{��Ӑ�6Z��珲��CT�S�%XV.d�"s�85]��Y�&=����!�΢�UEo"$Ҽ���ϯ�Y���3�w0zpwQk�l"�����ȷ`�j�Oʏ��W�k6:��K7�}�1֏��}��%�@��y�������u�b ���X�l<�f�gP%P�|�u�-�l?���9u�Md��]��G�iI�Vي[oQ!�ϕ0�)��Ɔ�}&��
�*T}��%u��J�{fv���6�z�Uy髟E��ٗ�]/�ekD7�k�x�����;0k���oJ�ٟ��s��~�]C+�J�9)��~6@�Xv�_̃j/v�{��.a�-Ǵ�}9��!���Zw���e����r�|������}�q���Ib�5������py��^s��'���4���%�e�8�N_�s�c���%[D��t�����?� Zpˬ*b��M��n
��%o��]��~]�������7r�������v�u��h��!+��U}�;DN�ی�D���m��tH�ڑ�o��d�$�5�K'	]����m�?\E�Bua��xވ��>��f��^��&u��H���b�B���Jp��ɲ?����j�֫�m�ֹm[UwӾ/��]�pzD G����nۗম��M`olq���2��-Yq��>Z����Ԟ[۔F���n}n�!g��ż��ު�.wMKfk!g�g&|���g�dB�<\I���>�3sL�r����1,I�
}�1X�~���/]k��(Y��ɀ/���|)�l���F�\]p��
|��B�e`Vq���B���9����*��W?n_�l��Py� G���6��x7>P�Za e�A���5��`��Yo���l9n�>������U�w��ôsė�K��۝�F,=ˈ���6+0M������ڙ����{����߉79�{ڌ'���l:9>�����J��޸���D°�D������i�I�U}oF��oPl��7f6{mn���J���bc�M�'aWք�$�
h��NtײC#��� DT����Ke��Q�)�Y�=�<�2&�[�6���x%�����j��6(1a��
8d��_@1{D�>��Ռf"���o�Y�a���q���ܛR���\
�,��֠������_���]�^��������S@�Æ{��ݢ���|{"��5���҄�_y�15��g�㝞b@�2/�t5�[���.�л�w�wa��l��Nj�}�mZ��W��r�-W1Fa�r��yIۭ�{̤��u��Sm���t#��k~ڣm�V�6�lVثEh��hڋb��hD" ~���z�Lf2uz�O��g��yL\Zr�Hn._�7���xw��Awj3��q�:�vgT���3M5�!���
q�({��g6k��5�Ia!v��Ky�G�"��^-쪷h�4-ь�T��������_ξ0E���]�0kw�t��͟�٥9����@�p<g�z��s�F*v�y�[�^��X�%�����l���桩?6�!��;=�U=��b}62vd���N���y��c���s4�-"�i@�[���*�r�иE5�64Wm�i-�����l�eV�+o[{�s��ɸ�ȇ������ȱ�7>UX�?7Q�~J���{(S�:z6�h�y���i�
����4��47�����o��
7��ty;��T�Ԁ�J��*9�mY�k�0�}��{_�l5<�P%��h��s����X�@Ⱥ�ftY��1�]���9Y�[��w���%x��{�IMX�qG@�l�������Q8[r$��L9*����a�Hf1ދS^W��HG�ǲS�c#����Vܘ����ns��C�5�Dݢ{B���/_�����������|�_/���e��(�9���r�q �s��G�o��O���P��A��"�)���B�.6Bǎ��j$���ƩumH�.�El˙ڇ��+�TdD��,��R:#��|�y3EK{�����D}���M�g�ξ��yt���:x�� ��^��i$^���'CV�c[�5����)�����Ɉ8J0�]���3�_o��k�mߏ�6��uo~ë�5��<�d�y)�lK��y|Ҷ{"� ;�{��3�y�f(�:�<:0vx���pێ0���C�㥛�3R[r���a�Ɔ�|5Y�#���=An��g,S��5�S!��U,�2�a��/�L��Vg-��3}���yL%�'�-u��bY���i]ڈ��g�q��x��z,��X=O��nͥp����OB��{t�1.�w�"!�!=��[�yd]5��2?������6Z�o)�w�Q��I6�TT�7x�ڊ�g=�_NO"��@8�S/.Y0���4��g���,vɊSYB/��������g�<jN������kT��Mg��d�8�w�޹�o��y����j g�l��X�wl�^���J<09R�Q����]�0ߎF��>U)��ӄ�xfװ)�Nˠ��QSڈj�Y���y�-�]���λ�'B�ď-���tH/(<�s]㽾�uo��K���؍ {/7o���������G�k��nyZ�L��ݛ��f�C��&E�q;�y�{�/�ŞrG@t�w��d�7^���[�n�>�Ar�B�ow���P�G�^0���7� ��F�����i��˨〲�ʘ�W9t�:ﾳ��t�&�p[�B���W�W��_����4��C:i�v�Ǭ2�w+�k˒��F�K���g��W��Yݰ��ae����.L�佊��閪M�9�Yp�����~�KݼQ)� 9)��kc���Q��n�I�U�~��}EǓ%v���V�� _m"�f���=7���Ug��b�>۳prb��C���NFĐ�
��+�V%�E���a�4˞����2gS��{`_Hyy&]|����;��{wp�g�]�u!ݞ~J��qf�!�'����Xpۧi�b�p�l�M��jmP;��l�7����I��/kӿ菇��Z�><��=�$H��z]�jÁjvݲ&�kY{m�Z.b��Ĵ�y��d0�$	c��&.�<�Q�Y�3v%���q��Vͪg#M���}�_t椬�z6?_6���|L��=f�����F1��~���>�i&>��Vf��$NSsD��Tΰ���i�7]���'"cg�������f�h���͝Z�+�.$��5����#���ZڲDL	�"��RQ���2�/��3���W���m���`�d���������yb[�8p�=;4l�|�m�pKLX���;�c�;^��\
�Y��q��00���k��vl�=�.�YG��'�s}����[��M{����^�E�nU������@>!B@�-⏉J�H5�r����Q��(��s�K�\�W3��]ww]�Q�1�\��w]u�Q��I��v0`�1F����UȮu���d����Z���c��;�f9�hgwX�]uع�L�k�.��uܹgvH(���h��Ts�b,�,U�p�J��\�\�Dk��nF"��\���b9pɈ�nE9�h��I�&��d��sE!$�i˴X�,�FM(�F�D�cM&"�w�r��,Blg�X���d`"H�%S�UZb\��b�|I�I>���C�KZX�dK��.��� �Ƀ�����ַ�_o�����ٯ:y Y^�C\3�������HF����m�f�u,���<��c/���t�Y_<�hn1/��W��7�2!��L.��˳����������	�����mz���ʦ	5f/�F�?2�p+6�&�3!WC�h�������	��
�?y�(:r׽!�[�^�{��q� 2�\��m*{>�X(����-�� =�8���P�c��X�a�Vv�Fcǡ��3+�*Ll`Hp��0�-LH��Ե������o���W�b�ƺ�y3��|�oI�W^^q2{©���
9ahM����B:,Kavv�]/�F�m�{�i��Qנ�!mw�>��!�G@�1��C��teyQ�U��6���P���`����C��<�����Q&����ta�LH�����>���E][���J��)�@����QnVnu���5�ǏO��=9���	����L91�.��~�q��y��y;㕵=p��S�K$}N��Úh��<��;U�.�L7J=z�ύS�w����n�@��m��4!ρ��m"z*h����|br��mL������Lzw#nN	�����yΪ�r���+K9�Q�F�L,��Lg1q�L����M%�����˸ ᭴�N9:�/���p\�2f�x`��6}��fG�����
S�W+GumP1���ug��Q|�޽ۻ��y�5�?KҿSzpC�#�'q�;)(��6D*bMҤ���,�!��Ox�Bܞ�n����/p�@:��b4�����╪�Á�ӑhG| ��G����}��(�'��y���h(L���9/
��Q�S�g�5�P�ÃQvZ9d�5\?U�b����u��\=���.�ɍ7M��.��,y��غ��L��7"v)������6b�݋��x��S��F9�7ҽ��ˌU��8�����m���B���52K]2���4d!��N6W0y�\2�G#��_�A�s�k���5h�k�4�j���d+�y�-�������i��h��r�o}h.t*����(r���g��`׿K��3O�~	�S�o�=W�U�
U>'P��~7#��-Ì>=B�E1�b�	��0�����LF͛ڣ3(q�K�on��r�}�S�'�1���W�s5�
���N}5]�v�s�O]�Ga��WV�ޮ��n��q	�}�|�Z�ϊ��Ӏ���P84�t �TY.�h�ժ(=tվ3Ͷ�Y�n��PB�m5�o�&�x'�a�{]"�F�,.�����(�>��1��*��+�t���У��{��w���N�����u6&��aN7�ϚY�^���~�o/_y��d�%0�)qs�p���.�]����_�?gQ�ˏ����Qef;������2%#"�nr�Ӵ���Ŏ{�o����>gp��95�&����pk�ڄ����s��N��ǫ=|����7=��H�N;�Sj�R�Y �5*�+����ߣ��}� �
��o��3����O�)���J�;�o~�W��g�ٗ���a����<������T.+2��x}��{	q��h.�y!ĻC+��`Zd�m.�P�1�3}��\(2�8�>����O��سl�;(�EP�<�pn�Zf�AE�AE�cIq�>G�T�a���W0Լ����s��=ָ������&w_����&C[�(>kI�I���Ꙇ��b����o&w#cg�����/s��:����]�-D�5-��Z��'��wn��tk��Y���R���5�&*��-R��
x���r�0_��jZ�����ɂ�ܨ�w8}_E)c�>�{��E��b=0 �0����F6,[��c��S�S��\���Bk:͉�ɼ���܃s�|P��5�2O
A�L/�+��x��lG�w>���<��n��*�5�����R�_��xO<3��������2�$N��$Pb�g�����o��YA��+Q-�$w��2oݥ��6�>��:J}snTp;��:��;"Xt'�����>��}��7���K��U�g�.��{����p���3&T�V���.3x����Lxq��f�c����F��R�����H���"�.xY���|�	���6�����}�#���3�{��R�>W�ItP�o��tj�����������߿��ߧ��k����V�=�{���=���rv�v_"��m����;>�!T�?���6�bw�h�����.ŝ���9����X�8L�ay�33e����,�	w���N�ef��{�a�����vJ3.Y�y#w��ȹ'��L茀ȗ�,U��:/��-��B���@w-O|ؤ
[K*7}ȭ$fO;�s�+��;??�UeI�j�hxWE�=���֙�)�qeȋ�������Wc��^�;,�ׁ	Z�	��Ψ��򘽧*B���n.��n������vc	C�Q��n���»=L�� A`3lC���`	��9�s��%7F8��PBL�ڤ4��+�4�_i��9߽gWdz������u�_�P�.��[�s��3�>9Cj���>��á�s8Լ����΢x/@�b�>z�������A�5L9]\5:ۼ��<X�tU�Fؗ3��j%�WK�.��_)$B���/�*�1�sFϴ���z�U�n|U�Z9��Y�klp���r���v��Mg�㤜P�x[y0�&K���M���+\��'_���ܵ+��ϫ�\FU9�hd���21�Y3ہ�HR���fMTQND�ܩ��G�v�s�ުzl�dv=���&)l��Wbߍ����+4Ċ}�&���h=����4�{�������d�V�{M�ˣv�&��֦')�.Ucrq����ܔ"�̠�R���� ���[Tm[Dmk�^����ǯ���\����3WfC�ft�S�i���i!�po0Z��o��V<��5��<��l#X��s�[���q,ǪZ�j�à���E���� �7����Ҷ�nX�s�V���'��"�����z�t*��bG%W3�� u���!f"���u2��^ɧ���n6s_�Y��{E�),�����=z�*$G?�������D��F��C�'��fo���G"(����z�ό�^x��:� �Ы���po��YXc��?k����/��~�֔�B�X:c��0����t��Y�Q�\� ���+c���¼��'�]w��X
�ۻ����*:OR�+N	(�d����kIp�OҵᑀĲlA����Ľ��s��2���,��/���q�*�H��
�9�� [�K���-����˛M��8m��Q<D��O#�� �����[�0s��`v�yTg}�:��tq	0��]�^�}5AŦǢ��ӏ�'��fK���=������0�b`Oք`]�e@�y=�J��%�>K]]kY���hmb��:6v.-�?�k���Ȼ���t��v�'�\�{,B���I4/�]�����^����j��ؐ�`���O{;��N���j����<�.�&���m���-�$�Q�6]E[��Ʉ9�"u���������/o���Ki�S�k�&�^ZM��� HѵX�ڊբ�EU��x��x �S{g�?d���46��S�N@�����8�󮆲�s�?P�X�Ή�����RDZi\�p�y;��Q1�t��LCo�nG�h�j7��=t����1�~.��������U���+Yv[g�G��l�|V��	j)�70��&a�w#nN�~:pT�����7!ՙ�bk�f�4�+Xy��ݮ��gձO�>���&�\#ٮ�8B�rG	��Y}D����Sa��M	�� L�E�D�&"lS������\?<����yzֱ{s��\v}��Ł�-��/K����4y���$g^ɓf�N���U�]�ȧ�3o\�j�9,
���X�m���G�8����ה��n�,��Ɂ53�1"][���r����S���;�K�UNY�2�Z��J��zF�����F�y��'\��l�I���W��8VzԠ�R�Y����AS�F��Ҭcr��A�f�O��=c�o��H�<�/c��O��.��r��R�X��7�^-��`���{tz�Ց�a�5f�	�:e��,Q��~�ݮ4�w;x2��!��/Lۚ���=�HNڸg��j�ϯH�^1�s8�8��#�����G���څ�}G��<}u��G��\U�7�L���:x���6���V�J�A�FϒT������k;4���JtS����g�孬�mh����6�k&���|��w������2ׯ�|5�����`+.##�S�%XV.f�!P��85]�M��?J����R�'�ũ���~Y��@��Ujc�=8<
̨�El{>�ĩ���]M�[mT�;�rs�:��0��F�ǍO���.|)�~��@��ky�+		���[F�,.������vj���J�w!��j4D�j^Ѵ.�._�����v��Ƃ������f�aN7���ϡC�5�1�K��nj����^�-4�M'*B�:E���I5y$^Q�z`<�C�_*��*�-�5��$Ԟ8q��X|	,_0	�d(�$8�)C˭�cAM���z�\2�/�����Yp��vA}UN�{-t�m|B�M��n]��bߺ}�Q�'J-�ZK��}
��'i�22p�wWZ���y�D0���H[�rչZ��}�kyuV��r�V��u����[R���\�ޯ���.h1��B��g���~�M\5/��d,Mc��ՆDnUze��C��:4�w�!��Q�Du�T�9��B!b�j�3z��^[R��3Y<�L}?�zef�ɹ��J���$�����>�����qcSA܏|ƕ\� Ȼ��\YR{c�m����f�Α�TM�S�ԑ�`�Z��lֱfc�͚*D�n\fi�v�2����x_P^�s����t���w�[�d��i:{�K����[��n��w������_~���~e�֍�����V6��ֱ�j5kE��}��������J�ā��(-���Z%A��l8^Yb�,s#5;5']k����cބ�3�y�����,�� �m��7��!q��5����]>}��ч��ٱ�N�U�=��X�Iq��-I2
����yJ��	��C�qNȚ��	���r1��.��l���cW$�nzY�r�����N�g�i�HN���߱ы{��l	&��A�5��L�cdO���߱2k�q�
ruL/NM���q�m��Fs��6k�Zږ'v���^`��,���qi��ޫzɋǠ�*
epd������@�p��7j���"P	
�
����Y

]�bY�wW]����5e8�[��&'̈́?|��U��N�W�[��%����@w-KbH�_�^ـU��>�c�3��:�6P����)����'�M�=ʃ�M-����(�D_�yd'b�L��W����-5��'�ϯ�D������oS��4����Û����Ϟϊ�$L�a�t��ǋPƤ� ��b��`�
���҉Mю!&�����g~��On��̥5���gեZJ:��dA�ISWx���Vw��Z{����7x��Yd~%���7��)�ANi�h���<G�S逄f�y�s�R��<����s�d��Io}����k±�D&�����K��^�rN�ۖ�0#��-�T��1
�~�#�Z0|U�{������Ӿ�w��o̶Ţ�VƢձ��F��cm����@��۝��
�NI�؉��G�o�~�g@�_V}|P��]�3[�s��@��o�6sf��Ϧio��E<otV��oA0��y�W��$&���d!?��1Upr����ۼ���g�tU=�[�g���f����D��ޠ8�U��.k�#M�t�E�/M�8��-ς��+��y����yy�ә~d�;�Q�1�O�jN|k�b62����}dC�+�U9��c����m�;�0p޵�p��w��z�y�
�,�� �j�V����i!�po0Z��{|�9g��Β��|W_eV��;���3��X���^�
� /~�r_��Js�j,j�xlI0+�/�L0�]�gd��b��cH>[e�[y߳�m�5�]���sf(��(c�:E��C{����+,:���ܺ��.��2�Ռ��RY��9[rc_+[9��C�q�ճ$��<������Wb�-�B��!�JX��)N5&{���][�rt>��}~?,�0�pTD��P���G���$��p��
b
ฦ����Y�T��S�~�X(�7!h��_O�ju�|�1bk�%~�y�c���_M�"��mS�������p���w���>S�4���E;O��� �Q�j�F�{.2�9t�)�h����kh;wzQ!�m5(��Nr�r�t��:-�W�V#���u����{R)�f�0g������߮��ڶ(�X�F�mՋmfkZKcU%���R����nn�� �*`�� �&��Qj�]����ۋ=ә ��mP�Һ��]��Go���^����$�7ZY�:�؞Slo8)7����j}��f�:�z���]�������<�W�}�ב���ߠ#>i;��(�Slx[�I�k�]�|�KPS��)x��J<gE��ش�:0�Č�z��|�E�#��55f'>�=�JՍ5\�D��r�Ll�R���/�h+W��7�ׇ��oa9�确���.f���#��|�Ug��ΓU��҃N�����XK�C?!P�fb�f�g���2�?O|]c�nzJ9��}����F���H�|�����ᥗ@����i�-bfC��F �rp8��
#���%h��r���>j�LђR�����n�^��}[�~���W��}�"�*�j��S�����L���B�~~��6��*h8OL��8+�Y�ҩLC��0n�4ʭ{��H�ܶ���ep~>����PCӪEBz�Lj�no�����PP�q���m�}2bL���^>^W������^�_�������@i.�3�$�eԌH�s�/����=�^���ȨeFj��U���g��ͱU�{	�3 C܀�|���{�!���I3����R]\�(�΋i0=�òdjl+{�z���,���ʭ&���[UE^�q=qRa���������)lHST%7UT\\6�5E�hnr�����J�����Ë}7z{���1M�(j.sK�{��o�'d"3��=�/3�gf�ܷq�R�t7r�'xg��z/i�1���װ`p���
c�X�z痧m^�)�n�����UXFoo�O9T���tࡴMӉ�:���U*o*��('X<"��C�Ӽ��`;qwb1��Ou��=� �w_{�X2��Of��Jp6��
�;�J�T#Xay��e)�wazt�b^g;����W�������o�����O?z]�$�x����|fS�̖4��{�ԟ��J8�J	��{��l:�觱'-��>y:���v8��$y��M���%����w�݈�~���ՠ�gb����w��roe���Պz��Uqn�Ԉ���h�Ct<����{�oJvv��i$�d
J�u��[��6J�]�oZ��~�8-� ջ��7�}l[��❽�(�ݕ�;�dc�'μ����o��j=ٰ���
.|`��#FQƟ\[p�N7F�'6��Z������2d���ˌ坸�f������A~�sH!����̪=��U��0�le���;��B�59$�����œ麸��v�E%��MuQc��ˊ阍�ø�`�"�����On��؟�Zhv>�N����#�<=�]~�$��^�K{ٵӯ	f{aVyۣ|�����'.=���l�gd������3�e�g��c�F^]W2���g�;�q�<>g�?���yf���J����r��L��!�QڊL�=��H��^���|�K}�|���7觮/U�]��<0M�~�:�w�gЉ������'���r��Mf�t!��n\B���Z�Y�:��;�UI.38c*�똠{E�=�d6Dpa�����9�q]��7�כV5�#���Y�[�挍����?C�E�dn����S�!�Cr�IL��}sI��-�F]�p���j&`ܨY��<�_����(w3SmI�ZtC{:�U�Տ"���
b����ǃ	U�լ���DSs(��2��]댄XN��>��7Hg;�;F�ge���F��5hk��-���:�����ά��{g:�m�2��>[�w����Y��{��|(R|w����;�n��L�u���{�v�ƍ�۸��{�9�K�Ψſ��tZv$1�e:`Ȝ����I��dJ��Ҋ�T)��$����jfa�VV��^����;`�ܧu��b�S.6��}>)H=��k���p������G�9���C{��=x�J���'��,��L��!��S� Y�|=$�H�G�%��D��%$$�Ğ+�1Ei(*5��J(M�戤��ѵ�捠���)"u�dƈ�Xƨ�6��13c�2�c�h#����Lh�a ��&",B�E�#��$�D�I�Ċ6@Ț��"BLh)"�B4hCu�.j
#�6�(�s��dɨ��A&�"(1XƧ�0��^���u�k����׳`�����!Ͳ���?/
�S�=�f�~mҟO��b֍��A�"�WA�����E~~>=�����֩*Ŷ,��EZ)+b֔�b,m ||�	���6ɺ�msRBDs��0 Tةb Nr�b���/+p,�f�7��S�s���tCU�T=n�j���.ʋz�H�xeH�����9��>.�kpj�V�#t�@�h¿y�T��������Xg�ܾ�A	Ua�b�Z��b�������;���D�~���+g��lM�kf����2S~&}�*|�χCn���	m{X��<-a�B|�g��0�d\���
�n��+��'��(7���zK���+.b45NR
�`�G�k����Ks���1��к,�}����#+A7o�ؠ`J�L`*�IUU�r�ĩ��s>�w:s;<r�j��"xR�੿N��[fND
��&�PHI	�b/��X�l:'�tp�㫎��?=����"$�.��Aک���ᦔ���z���s�ol1��s�vJ�9�{}��X��_E�:���,�4��i�i��L����.?w�;�c\�k7�ۜ�^ަ�| ��� �FD��o`X۠2�gVD�����#]oG���r���dn!��c�� �"
��S�}WI����[Ǯ�ɇ�=xeU�+*qU]V��K��ȏrXZ҉Ex��,\�X��ۚt<Bv��(�Vɫ���2�U�dދ3�hM��5���T-ޘ�W[����b�n0�<Wed�^̮"��1Q�)���ML�>������{� FѶ6�hMh��TU���lUcT�EoR>��Ũ��>TE���]��s=��C��R�L`�FlkI�B�x��]ĝ��Y�>s���1h?�ϸE�J�`4��j&���ä�gW^�z;e�_�RW3B]��QN�3Rk�tL^
�U.��+.h �4�Xҳ����r��j_�3YkՆD����{��Eܼ��3mE����KTU�Q���,��y�W}���m����ږbn\�;�5���tmm��ﶻ%�L�SBD�Q
�=�NfÅ��pb�2,�xj`�������l�ӌ�L�s�=��v��Xc܃��m��!��B�e�]�◢���q�q��:)`Ƨ���cr�S��W�p/�4��PM����F��`��Y��䊖Ym��cxW�+���M�af�N��j�S�z]��cIP��|T=��@��z0^�^K��g��c��ѩ����W�%Rv�z�h.��Nvcm�,U�&��A8��[���b!��X]�C'�\�햬�f�cv'�X��By!@�U�/���5�����ٜ����@J���A5�.�ʶ�sj0�6�)�Ш�o���f(Hc�I�'J.2��/u�γ#�l��V���E8U�֫�؛��?n�Dn]�[2�����܆�ڔ��q���J"�S7'�ܸ�r[5�Y�����TBw��������6�򒱵��mb��؄�QcmQ��A�/o;Gy�f�!qY�dz����q��0���­A74�ڭwV�V=������;j.���w�f���GET1�b�[42�r��K�z�Ll��S��hr�c�9lZ�/��e��m=�E�2-�~�,{��D����<1<�.-9R<9q���^���X-��z
�L�+`כ��s��f0Sȃ���x�~��k�Nu����<v2f���Y%�.d_z�{�1�)b�}z:��	7՟X�Ÿ��툰�[�s��3�>�͚S��U%^��x�e<�P��y���=C�p��ƨ>~����xc�a��]\5:ۼ��/�4-��{Lau�|⦋g���;�`d��}aP��j��{�8�a�iN�r��*�r����t�C���gsЗ�[K�!y%��-���ڞϝw��C12\�rm���V�#�[��3%ٺ5�+�8��>��s�V)N�8��]F�:�U����i!�po2�^��ձ}Ӆ�b�<bު^N�Zd�=�R�l�ōT���r+��sat�53y�D��*C�>ϧ�}�)���{{���7�V���� u�{TO{�h��o�/��O"���-�=�t6\�w(������]���%y\x&�V��=ڛH�eÝ���b��
�L�c����9��FnC�\.�!:?m�SW���{D5_e��oη�X��j(���@ �=��\ޣ�6�}!����R�[y~�YѺ<���t:I�3��
L��E��ʮq�_���g1�y�p'�ة�%ೃ��Ռ��RY��9[rcC�kg7�O.�=u��GM�*�y��p�o{i=AB�y����N���Qf��g���C�pB��Ӡ�v��� �l�)��B�S]W:�]�p��D��zLrL���R�^wH�ڮ��ɸY:h�0����,�O��؝f��W�! ؘ�
-��\3�RZ�����퇱�x�o���X�X�+�ض]�ςW�)5#˅j�of�+3�a�
���L_����Z+�r��Iq����#���1�7__��֕�^�F��7�K:�L���gcq��5#�����lq����zkal�$7�b'��pM_D��^�=g�q�b����Ĺع�| l�]7RL�m����Vz3� �����s��\#��='�/d�ԂI�$���ͫ���]�`��O��D�B����H��3��8��gf�z���U#���J�`�0ڗ�|.�3��^$g�כ���=�8�y���lG\^67��3���ւ�f��K�**���0)I�
�3.)���;����~��L�{�Ow��]�>�˳D,�tH�l\#���)��{X(�Z�;r��)�fk�p|���=�{�'��ѽ}���8�FQ�g��P21�ߣ�ڗ�k�6%G��\F��4���D�`�v�"�8���e�ּp�Q��Q��UU�Zo�o��g���D@mE���hRl]���r��[��M�u���؄�w�,iw1|��ঃ��͌S�3(~�u�U2vn�J��}�y�^p�pk-%�㡨�'��P�I^Vs�"��ڞL^����{K�-����5�d�ENO[6r�ֆ��򨮖$K�bG�ة"	��b��[kpb�,p3�fj3�{mM�v��K�F;T�ދ�������'��)�%�s*NTm��;0㚡���[�V�*פiN�j�����ٗ����3��8���;"k�@�#��	�1!K�F��o+^��+���_�0b�"�ґ��kdy�6�t'INƇ�����1�N��aP�D�A���M�������$b�q�L_y�:��o���TE�>+.`F����DJ�����	Jk
��~��<Hf����\�zM���ؠbUjc>]�sS1�
�V�����\wT��׺��~겣qJ*�d�gr����%~���<D�ك)�W�����W/SX�V��S8��k��E�ں���z2�Z�;�i�z-ᨾ|����q���{#���{V��m����4B�f��c7,K$ǣm�m��C�o�(x/*G7!!Um�"�T8��^> |���OS�b^3?�FP����*m�Ҡe��C^ ����Bo+		NC�4n��.��1$ݨ���:֯��I��)����CPg���AU7r���JL���Q��	���:��	��8QU�ײnOkmx�}��zNT�u�5��+D�x�s�c�D�����z��7��w�c��>,q�҄&��b��d(�$<�C-o@�b������ �1����pwj����<C�Y��\8�iq��8k����ّ�׺w�Nl�X�ؘ�lO`�E���w���Yԏ��	�.��z����*�gƘ�~SV�o�ۀ���n���OGlәƆ.�k#I�=�Fe�#���-	�}s@�9�PBƕ�r�nY�M\5/�k!gɬp7kђJv9�e��������r�O/�����#�T�34e]�,[�X�o�U�\�s��l�t_l�Q+	�����0�:9*2dGLȿ�u�"��a��ˏ�֫s"��8�u�x�ns�H�I~�`/V�Q�҅ΔɃ�r.DЕ�W`�_��DWAϯ���~5��k��(��\В���Ν�u��F^r���C�]�iz�i��ڽY�������t���O]���.m��!�9����[���1'��gIh�X��{U��R8�hGB��V�[.6X�;�O�-���e�	+�w�xP.�E��fV?�� G�@}�O�<"rm��T��59���N�$i��}���*�rL�A�g ~��8�PM��	��#��9�q�:�#Ss�q��N���C��Z�E7��Y��NI��c����v�l"��kw��eς��emU��y��a�R'��L��J&���������!Vsy�_�]������0V�t�W\*���Q~����&� �j���^�|e� U�F�I���?R�
��e�R�d�c�>��r�Qދ
���L�hZE�Z���Ω��U��݀v��uךmwG4�L���2i�Q�=�2%�8��ګ��~"D�K,��O�6�/�K��ܛR��鞹�ީ��3�Yֽ�B�S����m@8߰1�5j�M�\��of��M�֊1p×��T2��^{�C�J�}������9��уA�ݙT=��<~�@q�&�����6i�62g�_��ƛ,�q�h�N�ǡ�'������>y��^��Y���q�]�3[�s��|�o�ױA[z��4�Td7��w�q����\����𫁷T�PCi�A��#���Cn��?@!��c���u���X�K{θ{z��*�����N�2B���G;�8v|�%��h��'�k,9�4�q�ī2��ȴ�!��j���Բ.	'ض��z������v�;z��r*q�aǸr��N�^4uhZ�[ۗu)�����   G������eߙ=��~7o>�tyO�T��ٚ�aZ�^UA�q8h�mŸ������<���C��7M�'w�Ҕ��r<7�8ɐ�/����O��Ñ4a��#��ȇ�y\@cu�E�ڼ�@�}'�5R;o��a�b�� �Şg�0|�jP����i!�po2��WV#����5�b��G��+�N��:gݛ�ʌyS�T�8���S��X,���4$؊��ލ��wϡ]�o;Y�O"���߬�����F�򶦲���U;�t���~�\�+]o��eU�k��H]�b`=@�	jf �^����c!e'��G��sП+[9�c��/B�ji��̝��#���E���	�=lA��jD������=�c :� �=��=Wʽ���O����r�o�n�ͨ�8����Q��AҸ,:i���l�Y�
�p�n���4�l՚n���5s��������}����6Tb� ����F&+�ҋ���]�F_fs�~�U�f?a��g�T ��^3`yxಪ��%q
/��:��&���t�pA���xp��Q�d�Q�={n-�i�M�2m�Db9z�2���"�V9"(F���5��,ȕM��%�$��a���Ĳ�R݃m��S���^=
���J��&�#�U�$�W�5�PaQȑR)�B����&���YV�g���S�`"���]~��xx{�j6��pS}�~��3�r�5��(�7�����F���a��J�/��Ϝ��rrES��:|տ`LGv��R�B�;�n!����&xo>]'�{m�$f�bb{hF&��^�N�U�S�Ӝ�N)�i�[���S`9ɚ���+���R�!�\nӧ�C��rö�r��j��b���K7񇌱�TM�O��U�CK-�`J��&BmB����q��n��I�]��  ��a7-�Ȅ�r��c�|�[O1@���~�+j^KQL6�76�3��yUM�������U�� ��`���Ϊ�r��z:#y	���)��cQ�yƆ�k\���{��c��|qn	
�b=�U�!��s��?)��=lb�2�{�~����Bɨ��{0���q(1�d�{�8R��T�ee�)�*_FC߼�&,j�noK����7�XQ�8͎�Sl,9����>f�=��Ym��f#=4f�NǄS���8��*�X���_j�f�>׶��݂���h����U�8U.%���%d���"Z�'*6�!i�fsT>4b�챜���������rj\U�=7�[~�b�S9�Kp25*��#M�E���fѧP��
(��!�*DA��u9�û7A��;��gE�$58i'�"��T"l>�E�x�}���o�R��E��'Ut��ru����-U��2vF�t�#�m�PǍ���[xlV�zj��| �v�=/�����̻��߆{Fؓ�W��M�@����:i��la���1��6c�qs�/:�{�
��9�6�t�uI�t6�r�{����/``�)����[��;��uY>�s�2"]T㾹���83ɼ@��Y�>�"����1�#CT�S�%XV.f��'���otWBk1aw~x���	�"�
U��71�^�q���(�S�W0zpwQi
�눏�ۄh\�Ӛ�i#oT��}��2�I�a�;�j�j�$5���i��7�u���#;�<!7��,���[�s��������¶�ɨeP��G�;��N�ힻ��OV��cYy��	ˌ�w����s�'Gwjڑ��6�i��N���ie�1��H�!w �V��N�Q�o|:�*;ι�w�Զ���0+ή�!�m�\x���7�/]���r��q�⃶��*���_�ڻϞ���6����0e
q��v<�9���ߑ�t����FF�čS+\�7�;3� �q�����$/�x��G�у,S��+[��|�<��4� W���������g������~�_����{{��8a�����\H�$�Ğ9"@��L}sU���6m��:*��~;�.�M�^n>�<%�s����ěx���Q컏z
�9���8}�}�vo��FS"�ꋷ}�	�ďS���\]&��%�N�,v�PT��h/.B\8�e������V����5�>�u0eU\�N���]fm?�.�RgC�8��L�œsj�m`MA�S�ºt~fb�H�F!/� ���k�H���pE��S=�����9ɛ�WYߴcW��7��Ȇ`^Wӧ?*��0;�k�ֳ��=�ƣ�&O*���SJD�}��WR�3f2��E9�d^�&����������C:�����I=յ�/6\���ͪ��$�sوב��CtS�SUp+�2�Ʃ�)����M%�3��VE��m��y ��Q�N��~��#�-^�w����`�b(�E�DO�U�
慴�){o|�$��署��:�II���[k=0N-�9�wc�ݞr����=����)�^u⻻�0�>��c�>��-��.���ㇵ��2JIǕd�v}o*��3�-���D�|�'J5��
��=�J��(�q@��9��d)���ҭ�T�oF�o���hA�d�Ɋ���a��5a������>�|��#��r= �5�/|�b�dC���E\�r���ۥ�W���=��g�_h�f�$�9� ��w�ǅ��Kn��g����y=PY����y�����0�6���<���^��t	m���c͓�.�{�1�j���ɗڳ�~�2��3k2r6�wy�K,k�3�ȜbҨ�0ȸ��&]Qx�M^�ر� ���ي�h�_[�'����Z`�mLZ��O4F�8,�[����b���f�	N1�6]9���b@вͭw�M����Q|�8!��<N�w�88VOZ+~�0�2��r��^/_�v#����Z�����_t�GU]�y�h�{6�=���z�N��t�X�nۍ��y�*ֹ^��aU$��-^�|�ś.�I��T�j̘�6�k#I�!��"�ݞ�(v����z�&<:0{Y>�j̓gsC���fr��ɭۖ� �{,dB{6.b*�SD����/���7B(FV��E�{p��2��u�@�qY.f�=������8^zo�n6n��&l���b��+O'uOa!�<��Ek̬ͽ�>�.Y|'��J 7sn�=S�VӸ/+�I�֐/����M�L�\�\�yXs��h�r�O�+z��M���Y��Id;���/������Cۼ^�p���L�.��JY8�x0�YJ���6�U�V�N��$ٹ��YwB�DIvk!����nNG�
�Ҫ���<���'E�3��I�[�Db�U+]+��b��;l�;�۱�����XpQ���K�I^�e���=�uA�����e'$�����y9��"Z��{����*'�뺭�i�0���5Cq�@��e�'�,I���Kĝ�${�  �>�,�ZM%3�A�L�llQˈa�(��i6"؈1E�Eˌ��*.�nb�X����J�!�ITI�9�,`��r�36RQ�|7
LzcWBB�v�,TG-sU
.pĕ!PE�5�E$��Źs\鮄��-sr��%��W*3��N\�N�]wk��������A��H��r��[��\ȇwd�w:��\�]�s��;����6���r�k�����[��rM���u��(�ck�~w��9���(�k���!��fw���b~��=ϖ*/��/���T9��^�Y}]�yF���>y�}�<�vo�������(����PÍ	(`i��ა[�x{���պ����bv���wI�9D�Zg_^�i3�$�-��9g�E4��ܮۖ�j���B�#�G^��)Y�)ܳͬ���ҫ��ϮԐ�"�h�P��HB�!b�X�oUc�@�DY��NY��w�<X�Y���Χ|�A��nB9�i����(,8sE�`g��_�מO�7�����z���g����myb�ϵֹ1�7J:S&h:	�[~^�6h6��R�͌�{3Ti����{�<߰n�S�@N�&U��	��?P0��Nw�H��t�n��X뢝
��Y������LY��[��q����?KN����tb���v|�`Kݟ?@�Q��.��sE��{D�M���'L�ҏM���m��3�:��3��ۉǄO	j����Gbs2����SH(�`J���ڧ̞�)�}R���X���M�$)������q��j�/a0ېX����Y����tv�X�t�`ZCXU�8g�R�U����UjP'�0��l���]�*=���&o������į?��dS9\�<)i�R{��� �{q)��(j~�0J ������<6&*n5Z��~�p��v�/�!������ʉ��U5p���؇���%#u��[��aΦ���x-��/���X^#W�줐�.��\f.��\1�y0��S��5�IS��嘋��#׵rȎ3_����O�-���7������9_x���=�
=q���@pu@��}d�G*���b��HX\�P��Fgbh�/�!�3��5�th���}�[��g� ��b?_�8���Ug�9�^*6��]�˭��ux���@�:��GE-M���F,�@o{+>�([��]�3Z�����~��~���?zj&��W��s4S[�'�sf��������	��XC>��1���#>.���-(��
ڬ���1^��;n�l�F1I\���ư�Ϩ�b���#M�>��&��l�����x��Έ<��J�f}[>��@����2e�_M,���

�6,
n�;/��f�^�ŧR{�ޒ|�a��ȿ�����Ue�N�r= �xWF��N���)" ����������<��pu��~�����:<��^�pjpZ��s���o Z4$ծ��b�p���W�v�u�@�Q0��=5ɳ��tx���V��v:N7D���$�q�.�������3�{?_��
E��G�
�㐷�:�[>.��%����&5򵳙���E0���-�V6���L�ʗP$��b��g�����
�yl�~�s�8�i�œ�!�0Y�DMh���:
���1
��x���;/w.��w���kE0a�$�.��*�8s�Y�Q��֫�9�rmJj�Y��)���ʝK4����>Z�P��(H��A�l��hi�����=�c.��9��V8)�҃��?t3>�b��X�>�DM}�
���A�p���ef�5���}
��m"�'��=�R?g9a��TP>0�ՂV���	�&)�a��C����TX��>�S�j-�峾�c����A�^8,��1�\B�	Q��V��f�k�X��T�������+^�����AV�Ծ��r/��+Í�[�Yh�3�By��Q���4�Z"��7~ܷ�Y�c��]]0��K�I�`��)i;�|�/�:;�:1�6$j�!�	���O=	�U�5Vo|�+g8��z�핟�a�I�s
qA��5IȐ�.7f�^l��*8b�9O�Uf�a{%�אs�T..=��E@�*�(CK-�	�ØL�څ3y�#��x�}�̜s�kM��_c�?1󭖪��ӥ�c��ط�<�#>r�IrYtKQM���ͮL��ul�v9װD����L�m�s�0�Dx=V�F������M�ƃ�NF讽�i-�1�����^�1~E��5u��[S���n���3ޙw���]+ޱ[N�P
�d�qd�-�4��7:�݈����hW�vt�PY�15�s%)tkCq	&p�������=�&�̂y���<9w{��cL���x��gH�,�?W��5�M���fm���'=�BP��,H�(B���B/�*�,rǎ��p��61JeXJ��W��r����5GL�z��)���b�)>�a9�B����bƬ����a�j$�}u8��Ӹ�����\3�z#buJ\V')-���&pY�R�[��,p2u[3Q�n�rW����]��ȣ�݌��6�g�vT	"b�"��7�_1t�ف;3��{�����]�F>�f�+�GE���0��)AYЬ獜2�[��ψ��V|,�V���q<9��\�g9v� �i�S�g!��`[�р}^'4W��!ߓt�¡ޙw���z��Á�3�X��0[�����0���4��TE�
˃�R�JQ>B�S�^�Hl�d_?���(.��C��+@�\�r���7���@Ī��U0}%UTNo��z���o'v��$�	΀�=�[	+J����	z�~VE5K�|Cy4��#���4`!ڥ��x�~��� ��1��'$c=&=��P���Ө*��L�%A��� 	��I��m�y ��;������p��	�&s�U-�&����8�&\%gL:>z-`b�M�}�a���Ĺ�{9?S�g�|]�]��x��W����_e�4�o��5��Q>�븼|��vB;�{����������oe�S�3������F�&�i;9}�{����X����n��'�;��O���Xc igѳ�.<Բ�
oPm!�.�4�ƪ!��0o�ì�z�(}�X��6=Ƃ�`.�!纪n����K���O�e�����|sJ;~Y�Εث�T�ɋ��0N�e���������~x1·��n��ʜsf��-��3����~Q���Z�hO�]��ϐ����L[��i�?7n�v�`}�,F���c1.�+"�Q��E-����RND��t)�TS� ��>�JQSW�3��ǑQ�[��Q���9���'���ۥ9��,kO�n#�@|mkC����6�����~�$ζҷ֤��	e��K9����=�Ly mo�R`p�&��
�:t=q�����{��4��M��+�ljxjpk�ra�P�;S&1ȹ-roc���K��'��1,o��\q����=���佃t���5�2�~{��~�c�䉯��$TT�%��c��<M���Ȋ�E��)�n���ǃ�/��a�[�y����]yN�ۓ�.#����z�̙~5s$�b�)h�ۼ{)��$�W���~gG��~����ȥ��`�C�VC3�[@�T\̕G�ߌ�Wl�0D��s*�Ue��8md����-n.��k�G��ɻghQ�~��}s�;׊V�.�3�Й�TsN�iF[K�睈?!�&��w�b��L�l�d5Iㅰ���K�������s�\��O�#���O�* �Z"a�`J�Ma�R-j�P{e�"��6�qڒ}{�9/i���G+����K�P���֏?��A�!���t���XU�;;�S�_W�[%'D�u�^W��>,B>�@���4%!!	,�Q�'�U�'��n�ˎ�fg�3�Xuw�~P�yE��Z���?�XdE�7�{����q4��Bc Zr��U(V��3�U�w����q��G%���npo]�3�yt.�!�~�@q�5�'�X�ݷ��p���uչ�u�Ʋi1�2e��	^L$+�᡼�5ވ��.<����;Av�8��x�U�>=��jyS[����ٿ�6r/&��lϘ�ȫ��Ta����َ��0�ed����QA�F�o���w�<�:U\f�c�;>���W'�)I�k
�ډ�+��p8э}�B�X���{�U��5��5�T��U��� �����F�e>�j]`���)����~�c
��g*^�������B�хw�\d9�<'�1����(����V_;����K7F�&��;�!wYd�h9Bf�O��D��O�>�}�$XQ�\vb)5��)~}s�a7��cq�{|��L�q�S��yqG����{����]���g4��8����}�q�i�2,rǍʙ�)�61`x`��ޜk�W�nv]7a�����><L.��xpG��.Ց��b��w;��ҩ����\��6�.�,�@�]�t'�i�����Ч��#��81I-l�qm����x��}>�MM!��B�nI��>ް�u�jxKV�ζ(_L��6�C@��$���%g�ãL��c#�RY��������՗~^x|��g�o=~o�rj�$MձhXC{��N#k�pu.V�7�%���Y�9c%Ic�x�ks���#h���Y���ea��~6%��AB�y����_ʝY�DE�oa�"O�o1���{�<��0��G<��D5y
��
�1�H�Q�tL� ��5�
11ȂRN���~�{��]i�h���^�8$ϗ���U�Į!BRjG�
�8��#�p��8����J�B<0sYvv�]/�F�m^?�MN��m�n��+�f����>���絵������؞Sn����X�ptC)i5�Bx���ݴY�������r�c���[j���ͳ���N�JR�ə��ws�'W0MBc.o-���u-�Jj*n���f�d11mГT��8�\>�&���{�����˫g�����DЪh˩���o`�������r��\�R���Oa��� ]�/w{��#Wd,���ܨ2K�TELe�Gal<k/h��ʀ*�N�0��at�j!w$fS��}.7)���x������z��Z�Z6k�����Ü�B�&obyQ٣���ǥ�(p�!6�L�붳1��l�����Ïz��U�<�~~�r�>x1��P21�ߣ��\����6'���6�#5�&��n��9ٿD��L1���Jq�p�ꪷ+Sx5�y����[�즜�~å1��T�u-�j�A��c�G_�j&<+��X5\B�T�+v������8�X�Mm�T$�4Fm�Ou=R��S�L���',�AN*5<��Ym�����R��;?���a�up�Ca����x���L��7"v+�$>�(A3�Y�r�Z�����j'�:fq�k��-zj��_u<�>��ۆ!�&H���*N��~<rEPpTѐ,˒�������P�噤��Ob?��zF��@Z͘W�=΀�p+41J	�hP�$18�+8r�E�i�l��4{���<��������k�v� �i�Jt��hyF��}gDɰh@ߧ�)~�+�j��S�l����ww7oOI_���6+X��N]�.g�a4<��������5�W�L
T��@)B���ٚK-OZZ+���;�xL.�톺�e'Y銿��\����×׈�w'cՇwrCsa}@ƄD�Bٹ�D
��^ܭnu��S�3RG}�6�,P�Yj��^(3ɼa��N��D_��1�Η!���
#gy��Z6�OL+��pc����;~����7ly{	U���`�Y^��{��$ou�>�v]C�+c`[	+S�N��A��Xz��d���r�����wըM�n2qn�{i��&��8��#�)]E�¶|j�j}�"�kq��P5S�)xi�%�I��2Sm����օ�����Ibn<�9�;v<\KT.01�Yv'*}A��r*�s~��!��=�5r�Ͼ9�0x�ή�!���b�NF��88����ʕ��"g�5�ţk{ٺ�z������S������pc>5�1�����tk���ao�43�뻸){��:����F�gf���LP����E�>Ϯ�b���F�F8����jܭۀ��cbU�Oo���<�P2���
��.�b�J���Xr�
��4r�h�Nl}|�ۖAѯ�"}�.���#n����=���� �|@�3r�Z��Ʊ4�U8���z!b�}_[Mm�s���|�v)%��_jQ{ۂ���kZ�T��j�q�ro��>#�{�D�ނ��^dUuL:�&�V��r����a�x���O/.��ibD�k�,N���{Ӣ�=�K�ƭ�س��+�Z�)��!<��A�9�K�6s``����{�ɾ<��ɳ&�/�k!y���5��	h��Ø�.��5�B��n���xϥ�1p�Opgo�9��5<59��Z�ƷJs�2c�r&�P�� ���M���G��n�=���v8�l:"�*�+��{Fy/`�<U:�V��&q���S�'�ۊ�}��2�7�/b�.O8Hi#��A]�kg6�8�a�7����}:�%;s���ןRm�g���5}�Ŵ��i!c�n<1�Cf��#k���F�@x�zCoGGk�H��R���^*����z�}�=T� ˗'�ZAG_X�POa�S���=:-T�^baZ�u�W}1v���\����/�ێ�����P>ϊ��p���q��p:Dz­A���S./�owZ˜+�T���ا����#��X`T_��t(�48��b��bW�[42��9M�\<ƇVTT6&϶S"w����>�k}:���>�<��֠��V�D����鸬��1�U�1��hG���W	E���ᩪK���G�����97��~���;�N w������=��g����z�~�_���ٚܺ-�Z�˭-0˭ɸ8^�1[��F�fBkI�lPe`�px�SE�4p����8��N9���O�����ox\��*x�M�ұ�B�5]4a���M�Ն<Ҽm�ud��}����4}��h����_��5ʝ${�G���#���9�v�#��/e�/A���o���K�7~�>�鞑"ڮ����h�S��M�T�h�УS��V�ZgDkXdMm�w%n!:HQ:�0�)�H��5?�-$dW7�i�Ӛ=ٚ�V��A
�ђ��+w!0�ZqDUh+kt��1mS��0��Ɂw8��:������x�=x{0��؝�7��5�ܯ�&=a�7;�}��������	����}��1��<F�wo���z��}����w����qf��O6z��Y�y���9o�=ڍ�s^*�3����f ���;���8��=����7�ݕd��s����i�H��p��P�6�;��LӢ[�Z�u��ĕ�o���fwf���{VY�Nt��R&�*�gg����$��9,^�:�L��In�}B�Jl�JZ��+{�$v���΄ö��,T������5�7��Mh^k�W=�_ ���k�%��h�u_d��m���1�Br<�ۆ`>z6�6k{:��ww��j��iܪ�u9�˲�~�|�u�q��o�n�p=�{!���o,�x�Åe�=��A[Η����ܐo��cf6�K��q�6;;�{~�������Y��|F���l����9��џ|:s���{Pך	���;
�͜Wq1�S��g�o{Dj�.��GdA�Јء���;�U��A9d;-	��}��/�E�����_q��(b�d۽�����1cF(EM��T��)�im�r�[���M�ͦ�<�ɏ�Ź���eF6{�n,z��j[�m����2�sV}�%�y���;k2�V=���D��|������=(����9��vs�d�s�:#!�C�M�wO6b�V�a\��s���g.��n��%v-aOۻ�D�e�3�-�@�Cԟ{H^o�\�+�ī�\'��F=��ށ/=��MmڱF�S�h�ܜa7���b��,��s]���jɵ�=Wo����x.��8Ǿ\?���aԼ��_9�d��[V+��ǜ����}�{҈b"���u���6��M�խQE�j7ާE�}��z���`�k���\4��+�{�=\5oY�iE^;���Z{~9�Q����Vk������)�C����s�1�ƭml[���-�m~���S@���?HO��z���Pn&�F�j�'�*%��n���>��oli6|<����y���+V�J�C��#
cM��*��`.n�cQ�6bD�43EHM嚥�d�[$�v����'.I	��6�ګ}��]�	PGh6�N�q�}��-�X6�:=7��;Hco8.�_�qL�{�ɢn��L,cjv\(�`�ʘk6ka0^���I[@��I��{ x��|HlHc%��r���(�6�\�Ns7C�(�9sG]ur�v�nre��[5��*7wk���EEȮ�S��ܣ��#gqS�r�tb��P[�T&���[��ͱ��v�h��ݎ��X�K�)����cws��W"����Z9�p�IN�q���*9��j6�����g*卹O��M�Ӳ%Ύ]wm��5�U�nt�DEcY�E�ۤ��q2nr�m���sF��m�dc��s�:�F�r�T����չ���sN��sEŧt\J�ܸU��]�cQ��
�������*o��z�?p�!)ۜ�=w:��N��F:u �E+'s
Q�F�l������+N>�4�.��s����=��-���71���-b�6����I�ɭ4.g�6(h���¶��1�z{�Y��B�qt�8���O�7I�J�U�3���F�(�Ԡ	T��9�3Мv[���Lk7(��8Ϥ�5޳� �j	��m�Cv�����ό�K�����O?��,W٤�)o��2u�򵭽d�`����|j�Ks�U�[��`�Z�E*�ߕ4���5&[{qRA��\��}'.�A��#ڪ '��ȿ�c��L۔���	N)����0cp��.��F��?k�8��?{�b�}}{�w��1N���m�.9�|]k�|�JpsQ`��>�1��qvp�_�u�ni#��̆Z1l�H|���]�3U35������l��W}D���[�����TH�깘�F&!��
�rVY��^ڱ���͍�F��H�Q�^.�Nϸ��zv�6�sq��*�=�[2M�� ��a�f�M��ؖ*zqL�mW�����γ��?�_@8!WC����/]:�+������
m�Mx��M�ͮfii��[�l,��P�+3S��{�YǮ�~/���W���F98�%� ʲ�˜i�ž�A��p�\��'ꀕ����	�a�<:���k�su'�Z#/��Th�~�b�{5/Y7(��"���-G2v�Z/S�V��uˮ�S������_T�����GucsB�^@�TP>�
�1�H�P���f�M�]�/i�U(f�y����Y����&��|~�aC���L����y�W�c>J�XJ�H\'�c+�ј=9�6�i��@{�x��̶��-���yt�=�����	��%�#h�o��C,l_�n�������tz���Sdq	P���)KI�L��Yޛ�s�lHג���"5F
ֳGs�/�C�;hF>�Q�{�Cb}7�i�w'�*�|e�F��e�7Qv�7{�UI>�<Z�� ���a��A���E7�j�RhT4��@���%�!�P>W�<+{$j���W%l3���Fz��j��Ӡ��-�m|��}���r���עq\}���zk|��9�B���+��4L��"��n`��8nT�9I���N���}yv�{	,S�U�����cU�Z�c��8��\2�8k�!�n!Ҫcܱ��4'�͌SS�s��.��HV��j��z�>�:��L���r��5_�X9���B�j�nn���\��\������oO�h��`XF*�S��5��*Lc/k=�/&l�P�!2��ʹ�r��#��4�͌
bf+��$j|r�"���*�6���!���4�۽qw3��A=�:-�f�A֚�0L�)�8ƪT��SAn5�S��tDI��WoZ�f���7(ć�X\�ܡ2bL��'b�L�L��c���"��'ba�1wi �q��|��f����O=ϧc���&=tʓ��ې����ؼɌ=o��7�cxW�U��K����G�5�0�^�@��tJ�"uH���*�o��t}H�c�����Q�J����c�Kdp]K��N���yF��E��2x͙��&��w��yaw�<ix@���"C�g�B�׷0��(0y7�j�Z����Ypb�a�y}��U����O�̤}=V.����n&9�k�2f�Y/N�t��A�/b��*�1{��=Ý���������FaL�1^�m+WN�p�`p�)�Sn}{+�� �����y�0�E�v{�IGo��	��a!8t���v�1�S�`J����B�U?9<,�7�v��n-�[Y�l��K̕櫣})���}Hϛ��3�}��`c����4i��8��o�U�3Xi���="R�S��1�Ne����P�K]LCϟ����#"s��u��R���^"�L6f�T��m�H�F��ʋ���yr��٬;Q�]N/%Ⳳ+��(�;��;�}]�_��M�ޔ�	?0*Z��5��EP�,���r)Y��[*�։�3ǻ�٧���a�݇���<�Y��с��>cL��<�3�4���:䆷6�b�3PwM���zX�u�0$�.��Ⱦ˃iq��p����:���������ݭf*kyuB����|�X��GHn
Y���vK��-�Ц�ʥ�uT�<y^6�B�A��x�y �
��ݣ{�1�4�i&p���.�<�4r���C�l/WR�(e�:j�ɕ'��Z3�M\%/�j����#��1�v��e�kN��39�HBaj����*/�5;��I>Za��k��jY��D3�I��a mo�7�In�њ;j��.TEMC}�=�\�;>���yc��jxjs]k�ʄ��jd�9"g�����y�c��B��Sa0#�/��uuY����Klg|S�S�k�e^��2� ü�X���޷0�g_�H���Xm#��o0Am�kg7��d���@�;�	�S�3��RNJ����otT���u=�s�`Kj��Bk6\U$ni��Ǔ�z8꾠�,�&�}�5>�'�_�g]��˧��v�%�5��N=��>{e� >T	?b[�K�E��!����_
o]��h��B�#=����g�}��&�r�*��?y�����"�q͇�A��x�/�:����w$�M��'4{���}�rl�y\6oN�qz�;�+|���QMX�w�y���: �q��L¬E���#ru��-�O��L{��9�'Ы��9�B���>�²a�S
���b���Hy�w�l��f}'Z�^��d���ݗ���%%b��A�$JC��hj�+�l��)1PiЌ�EV��ip���g���c�<t������"8�1{��"ϩ@%�`a�U"xo�\ۮ�dC��{5�F�y��5�w���ǥ9L05�/�K�5B������c�Am\G�؇���.�;��L�=�Ly֦w��s��f�N�ݟ%Zf�v�L�c4JSb���1�z{�Y��B�t�3�ׇ��9�jz�x�r��5׎gcȍƚQ*%6��&9�PLD�;�Bm�����f�ʬ����6x�CuH)]\5:ۼ�����U�F;����ށ�%�3�&����"����?�5{�}��'�b�T��ƪܷ>UV�s�p�Mc����1�O�j^�n2:#齨U|�!����E�C�v�<W�s#��jLͩ)������T��3yMg�%Sxbr�|���0���BxQ�ϯ��9�{�|��_�.9�|]kY�Xn� o/P�\ZA�ᙩ��Eꃭ���T*�86����p��}W�ro�;�����.�^�-��9D�{�c����-���{xw���?{��:ͩTnyD�ۉɵi��a�"���}4��%�~\%�s���-�#���e�ũ�!�&�T�x�J2u�����r;��W�j#h�l/��A��3:,��+:7ʚ�qR2���u9������9��ꗽL�g���c>��L:A�I���%`����c!'�~��߷%Vf(^���.Q��1�I�V�^�ʉ����|�)olAA	0��T��5HN���s��b��-S���g��]�)�{%�}m@�ec��DO�
�v@�K��U�˫ިR�n���M�810a�R���Q���Z5y
���U�`���H! &�oX\4��	K��Hj���;ᢲ&�1�t���aGaV%M��|p^|U�J�q���l�1p��o���ٍ�0:�p��dk�ؔc�U�r�Y�Gl�q��o�dE�6�û	�����z�*�m.f�ri��I�0d�.�'���BMCX;�D2��ڴ^m������w�z���7�w!#�͠��}���V�z�0��8�	0���^���tnr�a�Ŏ��q�ޠq\���H91����!�O�bR��芆�[���w��~�`�b��C��]c���X�X*��Zy��o)n
��W[��1��=�ت5yxk/)�ئr�TD�A�p�#�F��\絾��3$V���r(hm1����ܷ�r%���ivTH�h��1�\��X����g���^�D�c��e�|��L�5	b�k�DM�e�U�u4�=�j`��2fX��r�>x1�y�F|�oч+j^r�1WRb�E,�!��_>�hS��������`�F�p��S��UU�Z���ݧ#�]���f�wt�	QWS�GW4����8Ш�e���5����7�^��_,x��M	�0�d8�v#J�y!��c}>�����9�ϥ1����"9ey���F���=�_d�Ǳ�oB�R�Wx"}ǩ��`��%/�h�3;���1fd1�MJLћr�(��f�n"ѕ����G��M<035[3Q�k�jo[�>k��~L�-�tʓ�pB��A�d��M�[Q�c���͗}X�e�\%Z�ߊx�`�l·��9�螌~��={a�6.8p�f=i�J�j�t���%F��uг�6v}�kߥ��;��)��e8<�Z��<w1�ʕ�>�g��w���0!`o�civ
�k[#�8�F�Ղ�3y�߃U~۟|�Ի�/"��t�bXE6��ǁT7����s4ưMa��	��d��G�vc�=[Q�o���	�5QI�"T�t�]5�5<�'�d�=� ���6J����R{�&�:�A���];������4��xZ��Ǔrk[{�ը6S�4�#\�S|��b�w�˼^Q���mo��A-�����L�9.�{�e���e���0�S���F^^j���n��5;�l�[h�O,����������E��c+�(���.�XU��?*!\5��+�܌����]q�;�^�7�	y��7n���i=i�1ڶ�P�a��#�ȭW�w�eQ�/�y��\꜇�] o��7�-�7�d�ˇ�ڗa����Ѩ����z�.ͳ�ŷ�w@�	jE�[��t^Q���?6�3:����?{-O�88���=Ub}E��՜�g��
ʔ�VD�=�
�L��l4��\�iq�����^L{����5^�mNn6��{��*p͚��ؘ!Nƀ�Z��ӟ!]�1n
�m�3�^���#�o6��$g{��Di�}�-o4���nQ�T��$ǜ�'�.h ��A}�t��)O'hG��Ug����*_���R��B��8���)�nP-Yg�ӆn#�wV�.�ƣz_>����;�b��X�lj�r�tԷ��Y�r`⣒� GN��Y������4�x1��s��u,�^Yb�}��9���������ɍn�����X`r�6�%T�3k�i6��G���hx��PK�7��W�@K6���m�q�85Zb�K&�����wEeJ�����۞���%���O��b�9�}�����f=QՁ�˫����$A��˱�r��O0�2e�U"��ⵕ�wK+i��lxL�!��\t�kgZ��u�����e�X)��tL�׸	�9�Q��z�s����?n*<,��B	�X!�Y��c}R%�����Y�i����o��=y�%�ՙ��Ў�<3�3Ԣ���q�!epA^��{�f���.���(f��4��4�=<3�&����Բ}���t��1�.ۈX�DL%" �!U��N��V�J���ƍCy�Ҳ���d�݉�cU��Q�*��� �S~Ѷ��Hdu�3��pZCY��ٶ��":6�4���~�U�Ϧ��Ih%�������n��48��b�U�^���εzlv�oѵo�	+;��_�z.r�����ϭ֙�?'��G�"�7���j�H��O\�u��rk��S�f�C�./=���߱j�\q��e���ȃ���}��	��8�+���q��	%�s�zp�l׾������-�Akd�y�H�M��Yp�I�kyVr�]���>!��!�?;�;�{"�M(��T	T�B��9�x��G��s{٦�߳��胝</��Z�3���������
�j*]�5�0�~;C�F���A.��;�m'���ۜWvBS��N���&y{�K@����1ە�eH�Tű	h֐�{�����e�cPY73M�u7%-�9xsZ2�ck|�����U��07WN��!�V��;>�v%���65
�6Z�I~��*�T�[��c�B&���j�6�᪷ 7>
�ܭ�c!`�vz60
D㊕[S�����'�*�Y=��}��5��5q�B�D���_rǍϕV9O��X<��0�qk%��O�"k	�}�ޗ9_O\
����mm��X�cT�[΋��|�ݥ��v�Zg�2l��j湻;�VFe�\.����c���H�#��:��Ws���~�<B�7�!��mI�}\A4z�)\���S��3��A�gH��Cp��!f'�#�5���縿OީA�2H���$^����������Yrc_+[9���yw��٘����	}=e��v.r�]��'~�9��Թ�L�]�>�]�N�Y���,�1�OxO�pT��j)3�Έ�]�M��qJ������!F]O��r�K�_X�G�7!o���E�*��$l���np�s1}2�yaV���/`�&'�(��&�MJ�����g����*�Q�����=^G����z���_����z�~�_��.t^����y%�M�vZ���"lVFn����0\ȫ�`6�m[�N\�\�r����^��w�CA�S�۱cK����kz�G��8��zVER���ol�����n�N�����v�ky���TK&̤73̩"uOts��8p�Khh󅇾k���^i.�=�����4md6�md�RF r�bdkE�ᳯ+�t�:έ(w�v-�-rg�2i*�����؇-���ҜW�uOv�M�� �Mt��N�.��'�ı�I��уџ9���,d�Yx�\Æ7!�7�<��B�&�COo������I��z{�m�l������KD푺�gVd���\�u�-N�L;N���B�H�ۥf�<��obT���,�z���^�eZr��k2���h�����4NT&͖�w�;�ӫ������GU}+s��s<9���}��/c�5��kw.Po�h�D_J��4zx���k��9��o`���Зy��.�e*���Nvr*lӭ��YO!�y�A�Ry�X�u'���Y:C�=������Q�DD����u��.X�8,&i�h�ϻ�Cf�ټ�7wn�G��v�L%��c`^�#׌��d��ܯ�S��97��d�z���};T5��%�o*́��wr#T�b^ի2�a&�a,0c>�g�x+G*�;�	;�yX����y�G.\ۯB]Hf��9{5^g�z�F��d1��Qz�n��9��%d.���Vy�.���9NW�{�����G_ ��^>�5x��Z�DD�
]�Ҙ:jp�X����@{9���P�Y���
s���.mq�6�m|���kX����m�y�ܱ�$�O,CsuN�`!���1{�}���K�)-��&L���E�d��v��O}��B⸋Ξ�k�2�<��l���D�緾-�OB�q�
�d=�����{:f��SnE�02����nQn����Ώ��`ʮ���$����ע�sw�z��K�^0y�W���8��}�����'�Y�L�������4�%l�*?}i!p'w�Ս��*4��+U��Ovp�d�8�BԖ�ty�ᮯq49W%����bc�X|}��Z�9��-Gx|8�[l�j�^�|s��� sn/>�������5O��?{�v�S7ؽ���m�k�$����pD �s<��ɋ~1�X��CG]Nc�J��'lT!�lT$~y��T<V�C����cxn�����Ǌ'�[4����.mG������q���$�ʧctWۓ��Qͨ�
�����'�E�;;�!yz�O��ۋ�z[޽#w��L��9�P�rh���0�9���^�*K��&��x�s�����i�����BF�#܁g��3.�d���"Y�;��^�d���o�����voK�F�$&V�/m,�d#��J���Nm˥I��%�Q�ct�������'+����n,Q��nh
�\ƹ��wmk��uەE�5s�s��\��&����]9���\�p�˔�b���wwwt�s��]�E����raW,���������[�(�.��s���N껺�:����TN�N��n�9��\ث�r�&�7(�;�wZ+��s��9�E�Nt��,���n���aE:�N�,cA��ݲ붹c���:��'v��vE���\�]��rtnS�t����6�\�+��T�.r�%�:Ws�;�`���.X���\��wkr�:��EΤW�G����%�E�n�V�۠{�k�f}�pw�����윅f9�>��RB����1�)�6�,Y� �ڢXP��+v^U���S��LFMIx4ȶC�Q ��N��f���d��&u���M�����7[Jx Ņ�l)�r�|z7+o�5;��O;��bUS{���o�`�dxC����h�(��c��j���2���xo;�3s��w7���S-E������Hz��Q���j�'>�^�ϽCb\ٜ��5�=�O��Z��"���Q)#/^Ӑ�K>�9�
�`���a�u���GpÜ�\,	��NGgу�[R�hD=�AW���{<��7�L�<ȫ2=SFa��(#�Ləb���)��=��(�o��a�	���yҵ���[�jy�
`����2�w#bm���q��ĺ�U�I��JH��n��#�5O7�s,�׶�w��`_���7F> X�*[/�ք=��8E��TaX���v}�cp�Y��f�1��}�8��lgIEXJ�ꜙ��@�Ha���PrpY����p�9��d\x��7<��|x���ܴ��K����M<�X���&$�ȝ�bC�RD>��>��m[W׷��s����3�yじ�fj0k�z�F����C�L�,2�R Ѷ���l}
�y<��؟-2�'���g{F͋��� ��r���������w�kVx5�1���_AoaםM���z���s�ҿG�=!y9��=�3��G�t�q���T��������1��� �&v���A��l13J᯦z��F��㽱�hʵv�x-(^�fZl~1��AsJlʥ�1!*פn��@�f�+׹�,9�цvD�Y�W����*���X�##��
��:>�c^�<}!z�ӡ:Jv4<����^�0��J�R�>x�	��
H�mЁ�W�c���B|�`�������o�w�g�I|�n�d^d�/��̗�����0���*±s4T&�
p(MWl��L7-|M�:j"��髥���iL.����UG�![���Z�ӤÆ�w��!�'��[
����u��s��9�d��B�W���&Ѡ���t�i]E��������DO��a&}Y���v�9O���<jD�\��sg!�����Rbn0��3���Y�X��K��j\�L�/rm�y���#��-�z+���6�o��z0��_���}�U���n �>1�϶��]*��w3*z�g�~y����YS�򬉯½,��sL�>�C{}�0G�1�x-���E{��p������=�*��&ɱ��>3��)(�i/�A�*��;��G������|���~��w��=����S
���ޒ/��;U�2��[(���n5��*Lp�N��:("4zC��t����P��+������]m57hH_�#n�3�Y�px�����B�E��Kӯ�O��/eЮ�z�{J�[�0��Qu�k���#&iJԤ����~1���^��ݸ'c8W^�s��4�6i&�$�.੊9Tq�����޺��J<!�߳�nۗম��5������B˷(�e�kT\�5PƦɮܝ�Oҵ�|,˳LG`�-�Վf�V9p�j[k!g�g&
�r� G�ⴱ�������P5�
D����
ynZ<�̌����s�Ǜ��7Jd�<����ך�.T��1�%��`���,6\6��緎]!��y1��<U9��&U�>z�G�ni��h��.M���� U���HБA
���>�]W�v�)^�C��
�s�,vE��jY9�K����T�Όtb���v�t��"2'��麘�qu��K8��e#{�E�Y�yO�}���O���g�*�� �n!`�V���֟X�@]��L�P�hk�����ʏGg�v]��'�Bc�M�$)���	
�UV|�NB��f���9�1�)nd�[�G�u蓲;��<�@�^2��K+��
��Bq!A	,��҆�����a��Jc��BU���L땦�])\]�HDӽ�V�vp�桭�{8��l�3{l��w�꘷)�{C�e��X�K�Q{=��{���E�����^w�,�v�9����ot�����r_uZ����x��<�����:
7R�*�fp�CQ,�쩿Ʈ&���k�1��I�Zgx���G�"���~��_(ƽU��G1�I��/�ךXZ��*B�Ǉ.7榨Z��lU=w����u�es��\z�sHd��`�dBo��������9�͚xq	0��.��T���@Dw4A��D^��9L�'�x4��-.؇������sg6iN�L���®Ϸ��ح�x��8�o��l/1HKIX��p��A����fXm�C�ѱ�g��*�b��8�)@ZV�z����'�L�	9�k�5nbD��E�,i��U�n|����ld,Mc��9O~�gM��q&���]n+P���aLL���kl�V�#�[���ԙ�RS�[�v�}w�]����;T��}Y�N��4���k� �47�@n��tDv���9��^�pjbZ��#/���5���)���~3���jpsQ`��@�hI�v��,T�d_��p���v���3�e�~�Q���1��iMkagYgsf(=E}gH��Cp�㘔G��}_!y��t�`����J�<fl��̍��'ӽ�:��_\i�
�0�	Vĝ�~�!���]&:s�+�"�/'i(��^c�	��B��&�����2�w��� 0E��M4VfOQ�2�q���7&qїX�1E���i�z�}�;p�K'���U�����fu��ooDMA��zV�^��5���a�:��TLs����MG��"m�(hXCӌ��˚�T�l�;%"O�ޮ����g�/��n
z�o���ea��t��G&�q+Cyg��-��0D���,
��9�}R����Q�<��a��TP>�
�1�ok�f_@�x{�y�)!|�Ԟ�)	
(���Qj�S.3�Z���{S�.o����:c��nYu��oN�KNS�tFǅ�5"�B����^��{�ZĶ�ܹ���$G�����"ϫ�눷�iLbw����v.%Q�XZmq	0����(N��S�ϲ�P�̿=T���=H�,mVt�ČR�+(�(ע_��z�Ĺ�g&k�
���O���h���7��M���U���Z� 3ˌ�t�O��+=��Ü�\,L�s�Gg�뜩[�D��ͬ���MyP<&<�a�� ຳ1}0z�3,C��.��ߟ<�瘠_�5�J�^��]��O��z�)gzZ�g�͍�L�v�Fm��S��%ǹf�?-�/,�&e뛚�j.Ѝ
���H�vJ���s�vyF��sp{�y\���/F�TeTk#0�(�]Q����1����n�F�!I�fo���;�E�N�p�:�)�/��B��ZQ����ҿοm���D�ё�1w�:��*�`���,j��T[SS�^�^٨�D�F�0��Q�_^1�ǒm4��ǣ��E�w5���j!ªc���nf��L�=d�=���ƿ��P����+�X��>٨ޡA�+�b�',�AN��Ⱥ��x_����I>B�0�d���nl��j[
h�%���x�	aX� ��#�pR�K;`���}q���3�Q�,�xr���opb߼����U�5�?&~��]@q31P�;��F�x3��^��:�OB�����>k�YcJ����D}�V��@��tOF>(�D�ڗ��hd�[�Z�_������v�v>l��X5����A�f�N��)�5a�0��t��
������+�тepƟ�?�<a@�-������� �}���;́DD�޵[�T�[Ĺ����D^�Ypc45N)��+3Dkް�AJ�d�=:=˴�Q+b����ެG��_Dw��g:|���0>��gWu�V��CbT�M����c0����*�ʪ�q&zm�����ND
��&Ѡ���"�i]E������(�h_���7'��Z�!�M��AM�`��7����z��?M�H3�,ή� G�9������Y��c*�[�����n�8Y�
<�v)6?S��3ޥ�������7���4eㄅ�Ǘ�WΥ��B�>���x�<ȼ/nR� �MM�E��ka=a�1Lȿ��Nt^V���S��`*�D�`f�9�����Ϣ��O�p���G��ޜƁ{�7VT�Ց4�(4Jr,V�����뺍�]��U��b?{#ώ]�ͻ�X�b�d{-�="p�@cn��gVD��6�/A�K����;�����i�.`C9�9^c��&�(x��R�m��ñ��
Q)����5�� �� v�M��,/�:wܦ�FsG�Nq���#��	���MӀ�;O�Vl���Ӝ�&����C�S��OS���3i�[�1aK�,iY�*�n]�5pԿ5��5�tّ���9��>�,�K�%����qUt���D�}Jg����s�5��PI҇ᥐ棟�1���P�h��>'���!���Ӡ�w�[����̌ϵ<59��ɍn�/��3b�eC9�Mݓ�*��Tt�J���$�?f@�D���/m^�Q��{��T�oUd<PVo>ȣ�yា=�;�c��iA7�85���1��.�8/�#���>��5���w5k+=S�%�`~ٵ�8�E�
˂�p��d� '��4{|4@*��:P���v�q��w����}a�x�،�1��ޖv^��A�7�6͚��NQm�/oz�"�l���7\�ۼ��r���8[	�F}e��sx��6(ݜ��4𘡆�LڌSvV�����:=���ў_[1�.NF���Xpb
���N���SVO�W
�W+�^�xv��y�Z�Y����8[�O���g�*��.ۈJp@�*T%os��o��>79|`C>�*o���Rd���`i���*�КHP/~�h��t�����D��ƶM�s}s{)H0Gau��uP{j��:N����('�,�Û��$���O�ԭ��ז�:��U�����D�-��Oȵ_i�k_;�9rU��2o�z�d����0�n��w��H7�N�v�#G>�!�����Fe��od����=f��I���
[��ɮ�u����u��[����!�n/66k˽�y�{zںv8���:���|�������,=��>�O4�݄�Slo��x�\�l� t��mcnۢ���ls�q��s���Ϸl��CV�w��u��u/�5�4�c��F%5sպ��=��$ެ���<ř�sp�r�ػ��j4�8��p��>]��r5��4w㳴:qt�����5�����b�0ױu'�͆��!����Ւ1t���;�0��`�F�F+QR�9g��34�ʋڨD��K��)"��T�R����	�v�'
2���r�+���hp��|�]q��S�����V����咪�	�Gc�<��O��{��2�6@a��S���ƭMi���J���CZ��)�3Km��ޖ�8\�ǜ:����pNMyEEE������<i��a=�Pw�ۿy57�ܫ'���U9��@o����vw��au�����ץ;])nro�?��ӧ�=v@T�b+P�ʞ-�;�U�^���hH�+`���X�'�����hYF�h�PL¯YU1�>k��Z"/�Ё�	���˾�s����!|
���u���D������g}�c��=@:�A��GuM=X+˛���P���G����ނr�x��G����ˆ+/��}1�P�%�'6��bF��<�K�����q�Zy���*�Eݡ�L���y�c�4)���G�t{(�[	�]�N੣5�a�u�}1�*�U�:�mFmaUJ��0�����B��0x��F~����� <A������7Ӟ�L�כ�����H&�����+  5]~X^��͈��v�O��볶�������y�W�}�$�=œ$$��{��st���p�ge�7}W�åҿ.���c���Fi��=+���5/��v��NM�b�� A�wm����]m����V���b,#�ߧ���=��{��0��2�+�q? v��L�컱K�ש�a���}�4�)nT��+bMM@���V�/ȟcLk�Y��y�4g�C��Vp"�y_֫��p��Y���3���ߙ�*���w��˳�U�=B[b�zB�\��.;سU�z�ܯqF[OA�I�O��lF���}(3t<�.q�Z�WNK�Y���^z�V+n�x������\�؅��q����-D3�x%t���}�~�{������(�]���AG�"�:+j�������_���},����*�xJ;�Yx��+����y����ΉN��hMtn,+jS�.j�Bj�r=⭙o{!�� 7�}�_��������_����z�~�w�7q��UDK�n�6E��T�`�a�M�2��9��s��5�q��3�/���;�> b���4����uR��ʒ+0FF[%è�$A�-�����ߙ��j�곙�zW�h8q��^d���>�<ٜ|�Ҍ;j��{�aW
7u���9�����y�og�*��z���F��J��P`��[����A�2��j4�|�haGq�p���jm��VDS�(�C��S�]{���{�(;p	û��h�qgBd���j`��v��k�2��N��r�$�_����x��������*�c2΄rɫ�Ë\��PoC��ǖ7�{���w�̎�s��C���oF�w�Op���Thq������-/zns��Ka���?����V;�<Os�U̽7�@���#��y�Ke��W3��)$���x��gvr]ޯ�wEW���{x�x��߶����� ��!%\7�O����x�X{�}O����L��R��E��rr�U"c_ʦ*���k�{��E�<��-�Sހ����7PX<�A�����Z��][.��ĥ���X�9��iT�GL��-A��uo�e�y�ư���F�/.�9x_���M�ɝ���F�zLG�(���+^��z�m��Vh?yA�*�3��@�!͹��'&�j����	��MM�;�xY���[��q�.�[��"��~���w3�<�3xnz������P�d�a������N�҆�^w&v�,7�o�Vd}%�	�J�=��_��]�_���}P� ŭ�뼉��l�����:=� �^�y:�|�p����~��O����>�s��^�y:��w��4w���GOap�����P�Y�Azn�Rв���qOt�����eS�yҴ�Г���;�qdӼ<��Q�h�FT2�E�
V��74Cr�u:g���m�ﻖqUB��ݵ�F����{����|r�uE��y0&76.�a�q�N�X�j�X)"�!�kO���� �9^�{�S��:���A�\w��OIͨ��*�?:�o�_2�:1pPo輊�a�ݥ2�[�b0��������z�9Z���ܘ��ޙ8��֟g�{��V
�^�.i;Us��6FM-�9��9�kC�K��Z<�pN�xIA���To��1欩�6G��o*/��%�}�]���½�E��Nx�i+'`�S�Mb
,�?�Ł��{�쓯8hoї�/A��Fj�[Ǡ����cl�!W��jU�Q��E�d����5mh{�	Tw�*N�%���r/����;.�r�}{��k����5�n50�{�+������3�c�����4J�y=.N$��v�{u	;����o�<h�g���c�&5�fcc���{u�g������<6a5j��T�ܠ�Ѫڲ�e\:uz����&����+ĸ��zN�+�{��שޟ���Fۦ�� �u��t��+�n�F���lN��wv�NZ�Q��I�d���s\���F��s\�s��[����5p��ngu:�\�\˹+�����K��gq��]4ۦ��n�\���7ww:܉3��It�q����"��Q.��7;�Kn\��1�E���B��
lvh7v�#DT��9wt�AI	�6��\��1Iw��Ӵ�;�W
-�I�;�s;��t庌 ��s%N�Wn�c���w]�P`�1]κ��;�g;)��s;��]'us&��]�\�ss�7wW:���t�K�\�	�rD�C�4���9]#7`uӅ�u��5�WwD;�hAu�2QD�Ԍ�[�9ӻuD��㻤nK$YN�"C$��	���L�]�p�D��H.]���R���0�HؒJ;���s�˸�����b�m{��mݩ�5Qjɼ���e[�������k��9�q*v�ܢP�A�vƗ��'*�ץ�d���
Q�IH�A�J���u}���o_������+��Q�M��S���u~��Y���n��}�s��,�n���~X�T�Q~P��4'��̓{f���Z�yCj)�L*ׯ�_���*��g�J#�R/r{inf�5Y�9�C�F�Ny���4��o
�)�S\Fzì��P����#�[/��%<R�9z.���;��7�����W��:�kP�.;n*gj�xjܿ6֛�+ܻ4������hN���S[G�n��|�+����YB�xeWM��<�������M|fBx��yT<=�'�K�/���(��'$C��]*�ޓ�x����k��=v}���j�h͉am��e6<�<�.�{b�+�T����w�R�xf���o��=�}�c6 �@��v�ʲ�o-2]��ƶƪ�6�E���V�Ц�{�f�)����`{�U�w�p���-�;���L,��wsc:Ĉ�}��3.\��9���<��yC��-�o�@��g�Y�~�Zܳ�Ή�ǭ��t���r>aI��˓·���{��\=�.�;��3/v���/.�3��~m(���u�{�r��p���7{�s�@ϴ����J��eD2�x�Oy�(-B]�a����=3j����kO��`�5,�nq�+-���Ѿ����BP]W�-V���?J.p�[~�}��4�mf��ckO|I��T�]���G�O%��6r\�О�;���Zm����`�J�|��`F�'Bt$y;�{u���w�緥x^v��q���E�|�K/���f_��ؓo�8��>o���_jt���5��N���t?X��d��}�p"��
���{:}�
��2%�D�fu���dLq�4�ez;�󞱥�����:T��pΡODI�a���mj5�V"{j'���|ǝMJ�=����O��z��W�6�61���v�1ƴm�mz����3�94���d����uA�T%krsָx�ݾ�(Ǿ�w=���y)4|�Ġ���Q�o���W���0�	ݵ�U�'��>Qc��91W,(��kN���FO)�Zv�x�-�&�;YAVT3�5#���0^.3rV?��;��tN�a�}<�o����|���Q]?H����g1n�!2N���Lf�K�"�n��sy�}��32/h��w��d�{�E	�l�r�A'sD���=aҪx��21�]�����n�>g�X��gɮ��v6�_Tg�B��ѿ#W���]ݾ'%v��;A�\p[����l2�Zϕ��#�ڹ[���3���|�p9���	`y�"�<�������v� ����Y�O����R(�i�[��7�O�O�ú$P��#wꔞ��)_�4��f��<Q
6V��Kf5�S�]ՙ~$���P�θܞ��h1����;�HN�8�V�yY�byX�]W]����[�ZYЭ^��wo\+���<<�R`�^>�9L{��B�J�a�u�Xx��>������v�5P��������;���y,��aq��m��,�f��Ҍ�~4�l�~��T	�G��&��c�뒺���-6@��S߱=���R��M��7t�yc���sV���z�����xv�ߖtn��J���	@&r?M������q>S;�^����`L��Ã8��5���ٗ4����r��IK�m�s�t�����lD�,����B9���p��n㶅]������m]�3s������<U7�=���+.R�p=�0'I
#hL�jX�M���W�<ǷJH���\���h��SfTH���~�����S��}]����SG#o�K����~G9��{����<���ş-����i��^\�1�0���6*_��v��eN��H&��"���$��Z�k%zc�C\O��u�u#K&�7ZP�M��_,�B�(��zH��y����O�Wv�U�*eײQ�:[�)y��y���<�Dja'hx7�{�v5쳽�}3n]���[�eL{�,�4��3+Ư}���e�|��N�|��]�}[9�Q�'�yqٚ�͵�����}�b�����S�������*��˭����O�fQ��:����>����Ao�����M�P��ٱ�2������x�>�掿��X�v�;��=�k����_	,m� ��A��5��;ؿ�ޖX��o︟���4)��ͫ	��O}Y7��ސ��]9+�M�Vz�ͪ��+�����8�a��R1N�0��w5	��\�b��y�J�h��;��Q��l)�{�;���g�h���z�oՏ{�"�&�vI����Ԡ�o�}3�#g	�w�/!%���D}�T��r�
�ٗ��ꌘ���CK2���\��_�{�X���l����3��p<�����I�xXVˤ9l��+�|�����ޖ�����x�6J�,�P��3������ϊ�ީg��Y���x�Y�⟻��}F���D�����H��V���뷐%'�@R {�⌆�_{��O����b��nI�!$y������ܞ�my`W�y�Ѓ�	�>?N�������J�{�s�d������kI�>Z��
�B��kg֕>�8q�'sLyE�g3�(j� ��߰>�����UG�;�J�Ϯ\ʭ#�\^����<s�W�7"V=��-���H�H0����[�F��2ά8�p%Z��/�=3��TF����7����$(�$��<gN�:��{h'�������huD��h0�	ݵ�tlg�l>i��}W���e
t,OU�ƪ�7w�8����b+UJ��&�h�YV=7�w�}S�p��u�a�0�m����kL�[:�B�Ǒ�uA&�o噈���D]���Ĉ;2��t�oJ�&7]�m�ø�]!Y�J�cl�q�v[�4��2�{����n�zSo�����E{��SM��M�ً�N~�������d����M>�s.��v�p�Gݞ%p;��z�7]�.��pM��ag?[����:�)0{��/Nn�c��ͧ(;�L�I��̞Ϳ�!м�������a���"�i?�aL$����)�I��^txS������J5h���/���:Bb|�`�!�� ����^4�ͬ��q����tmz�=o�c~Zo���2HB`��s9�������)������Lv�*AY滼�A�����i���GG�=��y����s�)�<��//��63�����'��O�q���ܹ�E^XZו�����Wԯ����97��ie�?+���(����mŷ�|��F)xՙJ��-_	�
1��V�S�|���{ATl.��!W��F�:�]�}Tb���6{`]Q8d'�ȩ*��"FTD;��D,wzAһrp��'�1�M�]����NN�0��ys�8����f�YO�P��u{���ʪ����{���T�����8���l����p�U�E�3�ʞf�D��O�\�@Eپ��:ڱ��0C���N��p�[�1���W���x#���;�Oz��_E\]*���.��	�����L ��\�Ղ������E:��E �jJ���&�Q��ދD���x[�\=Q(L�5X���t��4��h;/}t߬�-�i�e�b~�!�4n;��%X�č�0�cY��X�;�4��9��D�l^��1gXW�Z�k��ݎ�!����Lzmp�]��iU��2^����M�^�Z~X�ÿ�ѿ��<G}�r��ar��������5�pr�+�u-��6��K	���I�d;7�B���u�n���O�����=�y%��a�R������-�3H����sS��廑�D,��y�������*�)��Զ#�=�8`k�߰�����dG]�izZ̥���#����g�q�Mp�ܔ]q '��~/Ltq>,����\0�UQ^M�[9pcZQH�%�=i-���h��3zȝ��3���$g���\�- '7k�-��]f\�J�T���il+q���f�UZ�0Vd��Z�$TUaR�.���)Q;B伅�44;@�c5�ʲ�ƚ��l�obϻ����&��u?>a����ԝx���jC���H�.�M�]w��,��J��鱉�X'��)�>�٤ƿ�A� �2���ށH@��Eu��/	Ks9?|�����ӠX�U�Y��s��H9g�Gz�_�<�9�mh�}cyO��'~/������_,�T"���N��!��� w��4$�����i��5>6`�V`w�'f8ټ�S�:�^�E���D��F�x���D�9Z[g�EuH�o�;{�w{6����X���HN�fip�`�/LXaW�� �z9�w�{+z�;^��՚}Zw�&�r�~]��rYA�#����ݪ�޴5{XX���u9���������	�Y���ڪ�e"'���lrׇ�]?+��C{����j;S�o���N׾���u9=8?�"��W����f��9�
' i� 65���e�F��/<�u)r���1N�d����&x�Bʓ{T�)�ׯ��]*��^2�z�0)f=��,�.�n���1��cc	�q-Wmh�p�da׬�'��
u#�����\���}}-#N��_CBn��hx�L����W��r��M�8!nh�S$W���z��pA��e[PN��F�zGk��+��k��No����^D���6[�q��>͎�ʫ���I6�p�������6�QY����/���,?P���]ꗹ+~�~��U��*���F+�;~.���g�=3j�e_����V=�j�¼쬲#pGv��9FI<bS�X�B�.���[y��Z:Z�3au��7q9:uĝ�����!�bH&�R�Yg ��gڙ�������8�*!�[�Fk	�s������\�R������,�����h���(�q�:O_m!���������?w
Y��Ǟ��~�y�QֱE+��vqG�8�g (�z�>6h�9��p1(q��y��a�4��T���QL������!����3����4J��B[����56�k�z���Zy�5�b�Q�TN�3��p���Ǧޜ�Ů͞+��a���QIN��>���	��g� �F��Y��
5�����e�Z�5M��\u��� Awa�_��C����3B�y���5�XnU��,�����syv\ja7{�e��'`^+>*а�;%U�߼4�ֶST:����#Ӌ�n%��c�2~C�M,�GO�I��UX�-�ņ��p�Fn_�G���C����j�U�ˣ��9=�5�T���f�����$����s��M�;+W��;'I=�w\=�Vd��|�u;������hv�!�������UZ�X��4������ϣ}o�y+�1���I�����/���k� �kM˝(<���ݼ����o/%f��0�`���E��\���6�Dy<ǳ��{��s���<�o�� �Ϳ�!�n,����q��Ƹ�]��^!�gɱwR��P��j1[oB�k���-��r}�:1eÁ����&���1A�V:$!�)��|C��:�P��^4����4Ћ;�Ǯ%�h��mA��p��<o�+����h^�_����{�~�W������^�߾3�kcA�
w��{��8vN��%o�I�zj3e:�cgnԘpڒ˻�+P���G�(q���u�]��b�5�bPb��M�mU�f\��l.�":S�.�m���t���3�b2u�
��r����[�VE�۪d`+|��=���v�Aɣޯ��V	�e�`]��Ȳ��M�Sr��yMw���^���m/�ud{�����YD���W77c%�AS.R��si*J�L*�
,L�SR���Pe��e�YO>�U�,��:3+CAkp�w&}教�W";=�|:�	��O&����w}�	�o���;t�V6�;���AҰ���3�ǯH��"�׀�V���{�ɏL�����1OO�`�ӔA���wW��fA4u^�M#zu��j1�`��tе��%)�|��j��NJW�.ʔ��CR+JȔ(K.��ݜ.�����B�Q�P�w�L���8�n�T��$����OG�A^{wC�rC�SKva#�8V�l��r幚^e��)S*�H�N�{�O×?o)���Y��a ٻ��DM��[G�:xt���bΫ�N}��-���&���Bi���{�nE��}������+�+o����'����+���z)y��`
�K3�{�^��WϏ6�� �g-A��oX�!Z��N������w���|�a>n��XY�-:��G��g���9�*#۞�Z�CB:���Mw�롨���CU�^��;�TiST��k�{��Ғc{;��+�˄�pkŚ��{oa��ӽ(;^.����<ㄾ�ݻ���v�C-��y7IFI�^=V���&I�6G���,��+�_>#���nzb�I�{σ���s�p��s���K:���g,O�w� ��q�ט������<M�;�(�3DA����g��=zX�%oGS�����yY��������_�֊XyT^�v�t�����m9�ON\i2�{��y�u��;~z�����w޾Ӕ4)�o��.�ӽRӷ��j����(��_V)V��q��%l�sgr�g[ *��I�@�b샪����K��2�;���Ջ1�ڞ+�^@4�����X�K�N��Cl�����ZD�������59�G��t� B�<xz�:}�+.F*ݡiK�,%DҐ�^V���+s�nwj���mx)�w����ޜ\9����zS>/ĸt����V��.���c>����M��ކ���_[z��ع,��b���$��w�r�p�`x�=�6l��;Ǭ�3�?o:�We���>h��T��N�6�\�>�K��B��zI���8<-�Z=�:���rF��$����z��x��SO�.�D^>^�{1Z�oq�3�K�����C;;+H�d?Zv�|{��6G�[�]`�J'k��dz�OF��u��3N�}�N�܃Fq�����LPt������:϶���u�]�ށf���:r�4n�PG�����#�;��.vQ�ːh��L�wn�(���t���s�����s��6CNK�r�%�q�����;�F��MΈ�ܗ9��!������ɻ������ss.u����;��R��wt�S�w'e��jc��t�p���nQr��]��l��w[�L��wuκW#�����gN$Wwi9\@N�n����;�w.��������w	�wupnr�CL&n��u��Ƈu�2S��PFGwa;���Wu���q�;�����(I���Cb,!�wwR��΃�k�*'wr�� 0�u�Bwk�����Δ��w;�����#Gt��Eݹ�wIw:�Cdƚ�D1$.�@�ˠ,�wt�2';��L؀�] �s�s��N�i9�DJY��r�	w[��D��K���B�suݷ d�&��':�DԦ����9َtH���7��C~;���߻�r���D:�Gљhh��0DNJ.j����z�>2,}���7�Lc�o[��7�.5e=|���H)�g��5N���^���%XN >,R�A#X�b�b.�\���J�hCs��g�{��+�]_@�B��H���{z5(7pN�\�N���>;~�Ӟ.W��XZ����މ��4 q����Vγ}�������*�^�F	����m,�z��~�W�J�m0ǭ���)⺱�����$ym҄u;�^V:���~?b߫��<��얣&K��<���:�p���$밯�}���ih�irBI�ez�=��U�@�P�g=�5�X!DP�w���^ޔ}�Akޤwz誯�U�}л-�e���sA����%��D�%�9%�'=jVT�Źs��d�������G7�_�g�Ҝ�{Ւ�Q�Pa�~��9����;wd�Ι��n�:��W�4������k]=��{�Dz�}��-S�&;���x�N��� �N��߼�]u�A��0�?R��>8�w��},���iLN�k�{��ًy�a��N�*|)Qc�9�������u�Ʊ���G�iO�ar�J08�n�ҍՓV�v��]v�H9��`$Ȫȱ>R}��˦T���j��`�t��#H�e+��A
�ʵN2�T������y����"��j�2I*�C޽$�8@#�_`���2���t��mgɻ?:�G��х���]���'�V,���ɼؑA�C0T���4�t����_a�6��񜓻�$��O ه]bΖ%�]��{A��[iB`T�j8��&{C���P��l�g޿�R���F���ʑ�U�k,�������z=���@���Q��\�[���5��B�d{K����z�fYa�ô�־����Q�9����j��ɾ~�
`{��n�ׇ������g1���T�s4V(K/Óv��i�U�B*��^kM/ZL������G���'���ǒ�8!���R��qI��W˘�į�����+:��}���]� �����ޫ��>�����&�ø�4�iA��F��VM�b��(P�WE�+��!�
z�pg�#�U�#S���[NDF��'F���$�5��a�d��AE��8
�#^bc�$%x�~���˸\(S��E�����������	���ܠyVvT<9++��/7�;V�L�-���pZW���շ"9~J�o���w3X��E�mjy��˜/�ok�����9QFWZr}���TY��ps�:���~B�S���5�M���>i�
��y��/�������U*��fz���u�䤉G{�UpN�w�*�s�u�ͅ�5��h��.�a�If3L��:��-���f�y:��F�8��2�U�9뭿�~X��ysu����u����c���>��l�e\�-�=������^�}+؃��W�w�k��x�%aj�������>��,#A�SCF�B�s�|Mw����!��z��ϓn¢��y�ɠ,x��
��ܻ��D���_����c���*�i�Pe��ͫ2�G��\��ZH���Y��K�>������q���7�����}��Ϲ�+z}�����{�)p����|} �2C�bPFKX����`��������\�ߪ��x/�J�<&��S�ݱq�Ht���%x�9�#LF�"Z��Y�Y����֦��M��7E�{��ݽ^u��3���M����^�1���O.vbm��ź�6\�
wO�LC5mQW���*%��a��P�7��h;
\�J�p
ґE�l�W�>�T	����s�Rn�+�w/ <�R3E�Y�L��[{�_ug�+��
�y"���Qk�X5���<�y4/U��8>���Խ�N=�:�A���Ą`�\����	�w8c�vmd3{�3ZL��/%�ծ{c���3U%[봱:"c�7��׷�F$1y�h${䪏���	a^��X�.�g�J�� ���ŕ��ZH5��VHXM�y�D,;���/sނ/9l�#+�s׮$�U��q���w��{�͊>U���o�i��l�Mrr1�A�\v�378TNk���v�}WFW��J�e�������-wi�V�ٵ�ou/v�m���z�ǆ`�-�b'+���x���v��Eqϫ�C��96�kv�;;rͿ�^O^l_���^��rx3LU����^q}��<v�]ƍ�}�t���]���7��*�vo����!?��p����}&�e�2G��rn��9Lu�ݛ�0%&�]��X�����Bأ܈�33�,�:2E��m��'����������7�{��nv�g����0a*�O�&}���2+��������8�o��=�&b�c<�#���u�G�<��~���C�*S�!
�+�6ʚk>>���٩����ӹg�Y^��rU���
�!'�/��j�8�<m&���Q>��iYE��.��}�+�cз�#j���������%�\
�}��)+=�V%%�>|����s_r�B���RGu����/)�]��Ѥ�e
O��7�)���+们-f�Y{�!�9\*�Z�x�fW�7���qv(�,�j��qgܛ�m,��*�m�c��9���?tg���ou��{�CH�����K�FiV�O�A��]�Tz�ҍ�s�o�$�W����萶�v��ÉC~j'Vף\�{KD���Ѷi�|!��g�D����N�������'���{�H�bA�yW���/�#A�L끈�Dݙ�?�~�����h��r�?'৓��{|S��|Ծ��y�2E�ͳ�>�7������L�=�Z����ߵ�s�ʵ��ZO��׻t*���'���i�f?z�{����8;��X�vo�~�C�vW�IVn�����]�z���(�A4��c�$ߪ%���R[~0��&�'��eTz���jF@��*�K8ߘ�S@f㾬�~�����_��.�[�2�Op#z	��W���W�lp:²��Mt_��w��1���Ʋ�s���OTKe-�<��*�o����]|P|[��Wkϧ����T�a��s���+����ٴs�<;+R��(3���_K	�.�[�v mJ[���$��˶�яN�ډq}+��%0��sh��&���iJ�k��:������2���@>=k��Ğ,	������[A���$��,T��b��Tw}��-���m��YX#��\�%�{��<���W=�]q�<Q�lR�p;���}��X^2��V��X>�d�Q���'�˫.�!v��<<jP�b�͘r�iwx_M�M�l����܏z��8;#7'G,NB����h%�ZW4S��+M]%��V�*�l��M��Y9D����42���*�q�#^dh��(-���x=!���Z���=�-��J3��Q�>覻۽:v�uuٰ{�*�=�V��H9��Eʖ�N("��bZfR�+�@�y���@@f��U�_<V,��3�w�{�o�{�¨IU�~�^��Ch���lRS�'��X��}#��l�o,p�(f�ڇ"6��:��{��`��`�M���pA��}� ���X+���]wF3���-�Ҷ�6���yt-��6����
�5�ďcg�q=74�g �\5�9�){�'�H=���X*��3_.��r����NQ�p�ɢ-j�0�UǷ��^V%f�+�g��h"��د�3E�_r5O�>^<�3y{.i�?T�:�Բ�73|��6L+O��A������|Tea'�����)�	��|D�Yʽ]���}Dc��<+I�Öu4����X3d43�z�æ=!��uOj�~5�-iQ�����.�x��]_u�u��u�f}ݾ�o&�"XF�t�����5"�++��œ"�Ɏ����~ ����;lv�=冚y,�N�� �r�������jB��;v���.�@k���w��
��bX�w�p��6$Ȯ<b���f]'_O�uz�d�&�������*���dۈ���$M�$�%�#S<=Yy��;�g�B诰�_KM�SMc��u>�s����M��Ög3#������Y�i��ԐZBQ񦖃-���i�`G���:7��3o �s�T�Qx��� � ǨIFy�[��[y��[�З�z[>�]�d���z������Ϩ�cVY�-�jfb�����{�\��v��y�s���	<u@3�������X��A1�2�Y�N��Ӥ^_߳|�V{�/۪�@��	��y��}<b�GGg�y�A<�2����>~(�i��X9�}���MD�z����9>�C��7�OG�����HC7��^���Z�h����W�幇�6���'E ����~#�_M��$�@b����:��N�e������:o�V��o�Q?0熨��k�洙�;�Uh�(������w��ch�L�M{,�)�m՛����-^������0{���<�͋5NCr�p�^�������F���>�"�r�ӎv����s,oY���74*MAi�`�K�{��[q/uU�v��U�q̳Z6r���ug+bN��DR�RqX[l��մ�H�932�U���4���M˽��@aU ƪ�nz�� ����B��!�ۨ�½l�L��[��<;���c�Y*b�h0�N��,�tfd]u�����ǩ�i#[w����a���m���G\1�ެ�u|�/��]��${�.�X��ez���M�ĭg�ξ�2��O����ox�Uei�h(A��H���q1��o�Y0���L�I7��߶a���Y�'�Mx�{i� �D����Kv0�+8�T�Q,�e]鳵Ӟ�
eɸ��k�`$�`���rz��?P�����7����B$,uv̫��ަiw���ڱ����Q�$0Ĉ!��{� c���.ʛ��y:�mut}\��g�|�`��vyñ�s\�}� ���ˣ1+ֲ&3��^�\�W}&�r�y�Ƕ�fmk�w�BZʸ�#�����+}�3z�	�r�n��G���ɛ_7� ��+�������I�N�;�G�<��!��U�|�5z$�aYbFI��[�A_�����aʙ�O{��\�������fݛ����Z֞��B����"$E�#z��d�����cb�w2��7�O'Q��F�����H��v��ē�G&�ie�Ю����0�SUG3��6�2�w���������I�ݥcR�����]m�>�k�|}�����]H��Em���? ������x��ү_��I��.��'M�^tO�{XF�}N������LH�l�v�{{>��)���}gka�-�[-� �֒���GVI��KO��]ïN��~�;�'�]����7��(�7�Sٸ�n_�����Y�Gy{�Lj;�@�1�{*ݼ��-�:°V�����c���W�|2�˳/���p�4=S�~��}�R�|<���������+,�q"����I���͛�ƭ��� ��
;(���v6�_K	�da�C����{w��`�^v�`���Vp+�b��y'ٱ"�����R�Ox`=~�7����z}ޯW����{}^�o������׀��-��k��M���1n ��P��w���nl�@~���9(m*�b/jďz΅������ͭ|g&��\�9��6��^����\D��|M¨�+�gw�����=F\8Z+�reƚ��E�Q���ZN3����~I���4f���^z��O���Z���Y⋶r�LQ��a��z�z.Br����V�<���cs3Dj(�q�͙�B�,Tދ���]��~�W�P3���]����J�]�y� �¼��{�ˮ����gؽw�Fw��c�3Ռ>s��8z�����}�7�T���=�Cmg��ům�2X���6{�����/���y%��EǬ�7'h�u�YL�9مW��s�1o��s��g�J�P��o�X�=�$�z�n�tc��ɺ����1��~�4���~�vF\�iÌ������Ǵ�vf��9�m�􇟬a�e�u�)�u��O8~�p}�w���]��.~�!��!�a���_&���e�$�{�I'����q|�k��E{F�
�~>��ǰxܽ���ދ-�}k�W�Z��?.��my"pD�gN��'���>����/��?Vǁ�~�1�.0�Vy�=�3���x�K�fd�oO�����m[z�t�]³�6������Y���dߎOT��|���r������	��U�oq_w�,@M>�r�=����n�oUb�C�ቼ�V�w"�;�x��[��l���v둯F�e� i��ջ�1*�Xk�9�wMFǱ�;e_OG�軔�we�?>�m~{��ݎ�.�;ۊ�8A��*졑��3X��F�^O����ږn/_|�^���k��r���$�1��9qf�{��I�ev�u�`���+n�uX"�J*�]�4ȷ{;P�)Pnʥ�(�q�t�>�����!�{���;�{|y��}g
FN�N�gh�(�.�ر0���z[�f0��c�C�Wd֛��×E\M[G�wx�mR�kD�UI���U�u�j�	o���oԞH�oJ��Ё��e�	�Q�C���^���Y���MK"M"fl��KSp�����gw,J��Wq�dWG;��u.�Bt�fl鹞=c������}wǱ^AB��1�&��NA� ᧘�{z%E>�`N�N^�	��op�ڹ��d�J����z*�D$�����4��*{�1�{����/�z���3�NV#{İݛT�7l��d��K��Nӂ�Wo#vL�(�����S���У%)�ou�=����I�����/R3n���%���ྵ�����+�L}���T���ml�
L>'�G�x��yw�Mpɴ�շBc��l�� �v�Ş^��#�����������I��2
���Y1��FX��=��n�U�5tv��a�>Z����k��x	��%�מ�����3�pyL9S!h`O�B��s�F6FC*RdL)F`�p�$đ(������$�sr��� ���s�A��FC)��B	4����wj��(�wt�u�W:3�;�we�2v���&f9���K��	�&i��I��D@$��b�i1n�,w[���)]�a7.�1>���ȉ"n����2!۴w\��&���L�	\�E$�����!!0���LR%1�781��.v�����3�� ;�����F#� �;0��(��!�#wn#IJ-��Bf���Nn�@(���#Bs�(�H�E� ��(5s��1�hx�I>>�Fd��0gv���Fh�d��׭i@}�'���)�vtHۻ���o+���c0���o�u�~<;w�u*'�p��EZêU6^0�<���Ĥ��/���p��߹H��Զ:����c}ֵ���.���ӿ9�M�|��:͕��Z��Lzk���Ǯ��n.r*+}�q�#!�9��R!^�X\xam� ^2�9�};N��v5�r�v�gms�5��m���	T��S`WY8(�piw����ڬ�1�;{����o�|6�V3��	�2)̯0�V�v�V��5�H��97>�=p����Pm"O�V����X��@��u ����5��]��b��6�n���7z����.;��d�+&��g?@�jO�<��,���'�ٯ OE�u��"S��f�S��;��O�>��-'�)���%G"yv��(D��}\�[�}�M��c�r��S_��[w�M\��%ⶼ%,��CC�h�&�Z�r���V�"�B�&}����ӆ&��DvGk����/x��[<��P8� dE���0��2�()�]�P�AEy���,nV���ݤ#��3�dun�ǧݸ
�y��Ƚ�ըEY-�b��t*�K�S�����ޜ�	�d�o׼�[aHާ8�r"�	��sj"(�]<yߗNIc�#B�C};�g�y����gͅ�Lz����\,W�탰p��{¾ͳ|�U���Чu9�s�G�9��ʁt2�Ƿ��l�5�>�_�_��<}K�>��2�W�ha��L�c6"��i�>8���n�@���}^.�����U�
��.�X7�B�$0�����q´e�u�$��mcla��XF<b>�z�[_8Q-�v�����ˎ�ü��x\��r
�������\B�!
�+�Z[���fզU��N�O��gc�<��7�% �輟#�xx���\�}oS�T�핳�o6$_�z��\wҍD�'���&����� ���d�Z�����������@V��'A;���k�����NH���dw
�0<a�2+����ma�bssk��^w����ώf(��Y*�<��z�@�ށ!5��Q��K���C��H:���=ˆŤ����1t���L5�i��h�{��=��׿~D��eq��Z��'�K����4�M�4�HpazH���J�35�AVX��Bd���7WMV����|.�Dv�y�=���x>t��0�
dy��=}7J`;���:Q�5&h�C�4Y���6#v�4��3����䷶9�������`V/�����:���Vٗ�N�z=�$>��c�<K#ɵ���|�m�k�v�z:k���}��O�5�q���#�.�����Cv=��g2��8$��v'�-�8*��!�q�u�C�ힷQí�^��GO�Ca� �L��3[}�Ӿk(���idy)^�tܛ�L0����*�خ�½^�G(v������s�WiⰄ./{�ɠ:�~	�P7�>���A�s��ݒx��W���[}Ų���� �3��;o%_\�h�x����"�p���\;�.�X}��ӿ�&��������cjM��.�/��V�����5�����H:�K�?7� ��!��2ñΙ��`5�=�������k2�Ȟ�*Vo\v�D�A�&���!
�+�6���/�<C�>���e��U�j˚���ʠS׮���/�z�x�ˊ�y������L}�������������z��{������{q<��;޼�'�rq��}B�xm���x׭�a�����A�:�ɸ��)�;pq5.���_���Ook��	ʥPF�3V�C'�J��~o�W��q�.��2}�|C�Añ����ĥ�S���iºK�����f����nw�l?�~�ɚ�'ם��+�Ի�����C��yZ�SJ�5��3C�*��T���X7�<
,l+�	TVK<���s{���7ܕ�����̼�3I[�W��"�����;��]7�M8&�}ɾϛK.�����e��'f�����ݎLS��K���}��O����#�ߺ|Bױ��I۲m���t���C������^�b'� �=�+z�񱫥-��G�r�ܼ�}|䣛�=�5�hߊ�Ap�=1!�k��OTKo��	
�r��Κ��w�2�տ��"���H�����M���E��N5��=�a8�H^�b�9��:���/ϲ������+Ģ[��Jk7����|��Dtߎn>3�.A5�lJ���u	Ѯ��L�]�n=�t�����xj\��8r���۝� ���=n{���h�^���=��_rĨb�!�nb)�Q�v���=��K�@�fV�YB��3bF7f�����B�P�8���b�)h-ݬb�/4$!=R�d�.�,��5��l�[��Ƹ/r��r�3@��n�`�k5�9@z�~���'_����k�]|�}��X3c�ccS�����7^4��Ny��m�(`��H���v6�{hA��#�%�k�G��}D��q���^H���S^����tڵ�fe� �aw�Y|k�֏	-�ԥ��Jv�}~������8i���n̬3�O�]�'�m�!�*=��z��Q+ω��&c�[f��Qrr��+���	��<A�*���am���s����z���M���n%%�J�V��yl*7ÖO7]lࣖsK�_M�mU��z�}Viѷ��<BKx���E0$�m
��s�_g<�,X%-���=�ۋX�q�~�d6���/�^��@����P��]6s��ggx�yl�U��NĐ6�)�Ƣ�#1f�rr�Ik,�[:�ꅏ7P�W$^�3w��|�^T�������w�
qM݋�qgT¯��~��rc��$�ܝĵF��4�p���K���<����Q�wdD�w8z$�=v��'/���OsL^+�J��!s� Y8��v�6 ��:bO�6p�?�3�6|a;��[�)G+�{�{��.��K�ي��^���_�U�~57�n���W�|��ah�+V�/~��զ�:b�p��t��3��Q�G�tr�K��j���t�9��sy5�����i���9���_��L\}��F4��C1��+�k}��68F�T�BwZʼ����|�UK��w��Y��ڿ=�����!�</���@�Z��e�������3Z�1��/�ם/6J�|����3�����&v8#��r~Y�{CE"}�gs�/#�םy}�z但e�i�`[���[V�Zϕ��v���h^@��,C�nn����1�ԇ]+��+���6ʚk>m�
���O����Q�q���d�C9'�%��M����X�8P��2��-��ͮ��Q���s�c~�#f���?�O���u|{D>��#&sGC�9v/W��Io�v��\��:5}�����K:ܻ��w[��r��ҢiA�8�d�Ѽ�n�9�'L�ͺ���[�i����,<���L�t�&��-�Ux[�d�:�,��6�]J���Z.�IEm��J�QW��5"�G�,Fd�{ҁ�l� }�[�N+��Zz�����oc�K�s���<�.����0��Hf��^��SD���v�x�����a�v��S����>F:��Q�Z�M�}y����oZd����Q�	;eR�X��Z�J��u���<��	�g�l����iS��ֱH%�#:��>X<^<�[���D�ׅ��Ӑv/j3�7�Ԟo^ qw}a�7@H�3ļM��c3���N�����:�-6eG�7/!xz$�����0hb��}|A^�;Q(ߞ$a��?��T;��sE9���8j�4�`�o�߉k/f�tUTݤj�+q{e�v���ċ�&ņ��_�.V�CP�AGr�d�(SV�����p�ܷ|����1GW���fnzcF}�}>��
������Y��+~�
�p��2M,g������o�s?S�wx���b�|rn�LR1}'��J,��B�a�JǕ��KªqLPr�n����ju�<J���E�@y��>>\�uIs��I>r,����{�X�X �����av���K�5�MI�5�W{ϗ��۾���Ł�=co'��4vM����y��]qH� ���j}L_#�`�T_n�x5�x�>�s���n��^��>)T�����3������������^���0� ��:en��l��-�����F+�}����dv��d*��'�@�i�������{$����������i�X̵���Vl�_=u\{'���2����Y��=�;e]j]Vd�f�ѹ�g�����"���z;�a�Q��a��f��fb;5��g�w�{r�o��j܍N(b}7�,\�����5rz;�i�����xU �h��tx82�ΖZ��)�8�f�]���pꨳ�i��=������w��'�����W3F݉'9w�]���sf� �=����;��*m<�����ľ�~C�k �z~ұ�����w�:�LE���w�����AF+SL��b�t�����a��n�~>�����H��_v���u4�	y�>��mm��(`(�{㘷�I�?i:��o��G������^�U�ƴC�"���NqJ��+�H���uÞ����	5,lC7}�l��:�ȶb	�XA��jmnV�����x)؅IĠㇻ%o_�c�KZtzö�.���;c9�������pB6����To������7M=1}Uc	�G�[l�/��ë�:��$,$='E���$ߪ%��|#oQ�2q��C4m�y9xo���ٹ¬��x�_����Ԑ���ڿD�/:�3y{.^Tp���Kj͜����bΰ��i���m��e�(�le�6sc�<7�������S�}�<�~��(>O''\F�DMdNw1�%�h��h���s�co'�xz�
{u�P�^��çY%:U2��xSJ��v��/x��7\��o��c6$PN˪ŏ��n3kV%�W�g}�-�C��I_Kk�8SŁ4���;���]flBq��/����h+��+�$��r�ޙedu�+�ĵ1����)�q�����Ũ��̽~�2gG�1b�@q���3l*eD���j[���;.�,'S�^􋧫�Y�������
*�E�5r
PÏrw4�LMݲ6�J�[�|%ڲ�kH����.�倌���w5F�:!��x���*e�l"��7j������e�k�O����R�W�q�����[u��e��{��/�WJ�1GW.%�*2�W�ߟ���l��	�~r���~S3��l��R�X�vh=!���͎~�=��Ǻ�W�ܲ���^�}���e�-�44ǋ^�^_���7I��_d	�u�ƾ����Q9Y�Q����9vv})3�C�� �')[|�"t���%����C��K��(��+�SG!u�.�����o�'�Vw���PO�}e���d���V��8��S���&s����t��gAqm�R38����ꡃLJy=�֎�C}�U����R�}�E�f/�i���$�4���r}�!G��c};�`����|���.�X{��w_v�����./m_�ʱQ�Ȱ���Z]��l�z@�GZ��+.J"*/鿎��UL��m����W^����o��|kV�6�+fkfV�ՙ[3m�[2�f�Ym�[2�f�el�l�lʩ�Y���ٖ�+fm�6�5S+fmfkfV�5�5S5�+fV̭���m���[,�fV̭���[2�f�e�f�3k,�fkfV̭���[3[3m�[2�Y������[2�2�eT�ٛY��eTͬ�ٟٚ9��6ٕ�+fUL־3n�ʳ-fV�ՙmt��Y�fZ̵�VY[2�f��Y��*���ՙmo]�z�Z����S5UL���mٵU3mU2��fڪe�T�kT�V���|��m�e��3U�f֪f����S5��nmU]��lͶ�{��m�ٖ��UU2�m��U3m�̭U3[m���fm�ٹ]UTͭ�f�m�m�̪�e���m�f�m���fm�ٽz���m�UTͶ�2�m�j�eUS6�lͶ�5�+f�ul�ٕS6ٕ�6�5�*�mfV޻zoUS6ٕ�+fV��̭�[2�f�77V����fV̭���[2�2�eU����J��W_/��u�j�m[Z�km��5�?u�o�s����W�.��f���yr��x~3�c��.'��g�ޓ���M1ц��UTWq�����EV�0*��� y�� �@�M����.�9"����=��y�mf���꿟e��ߺ��w�����t~ܵj�l�Ujf��UYj�M��&�m�[m��USY��e���6�m�kMUST�U*���m�UM�m�ͥURm��MURͶ�2�����[k[�_ޤ�~�����ݯ�ֶ��ֶ�U�*��/��U�������0�xP`3-��UU�n�e��;�x�Nʥg1���}�C��*�����M��Ԗ� W�U�������_蚶խ��־o�otڪ���R�߻�Z���{����z�������iea��L
AUTV8���X��+�\� [m��=��aK\��;��%UTWFA�������1�$X*er��p+�L��\��a���ip%�%��UU�h�X�$��(�@L=���'"�H
�+�j�H1kEEVQ��oƯ�PI������)������g),�8(���1!����$(���RT)@�"U*��U	�DIJ�� DR��P%	Q@DB��BJ�� �	E)R$���{d�����EX�F��HT"ER� `�BR���%UP�Dl���R�U)�������T�T��**��J��!E*�!J�	*%T�B*��R�(���
�B�(%H$��)DJ"�I*�U*�PT�� �*UJ\   M"�*�X���qC\Ȳ�B�㥤;g�;��Ι�G:���wkD��t5�%�m[Un��j;j��N��n�t�p�ݭ����a�PIB����HPJ�  Շ�B�
�
/zV�ѡB������N�E
�:6�E����B�3׵@ov�]-��U���R��S:��̖ݷ,�Wkv�a�ks���W&E�M�[]���H�j�QT�E��  	�%z�J��:u��7N�wv��Wn�V���Z��&�����[�ն�t[r�m:��j�җe����c�u�;n�;���ִ��]�Ƙwj�����URIJ���UD�A�  6��Jh��w]#l�P�F�8
�զղٴ]�������n�6�m"���v��F]����F*��]�a�eN���@�5*	RIUERU�)/  ��/a�K�.K[��%�Z�(]I�j�Dԭ���j���tkSMR�UCMR$5��Zӈ���gT�TH T��$�0�R^  6����5`)Q��m�d;%M��Ϊ�	E ڨj�G �S���j�g'Zꎶ��E2��Zݫ��R�� �UEJ�J�  ݽ��Ah�P�d�)����t*���
uCUr�ֵ�B��Q�VicNӭ�1�
 :�ꪧmR� IPT���  � 	����g@���s�  P�� �# 4�X0 �4�t �3�� 8  �(�$J�AEHQRU^  Ӕ �� kA�8;@ Xt�  #,P� �� 4�3t  7T�� )��u;��  �"(BTR�TRv�TW�  i�= t'E�)���� ڹp  j� wb�e,  S� P� �pl����<���U*�� hh"�ф����# FT��SEQ�� )� ��@  Sh�*��h�A'�R$̪�  ��e�6y��*����SLҶu�t�g0\�U��`�Ol���=���z������V�߻Z��[_���V���j�V���ն�m�Z��[_�������@��!9��M�(�DTI��� ��e���H N�oM1��*M��*�5���qӡe[�M���K����%d�d'1���D[�Z1�(�sE�E휑ԁ���q^�U�LX�i�H/�YH�MV+Y�	-֑0�FJ;IJx�n���&��'�w��l��q*+vR ���R�@�����9�>4��Ў[���n�;H�O,L��71l�.śV��A�h��;�L�֣�kp�D�R��%l\$���q����F����YV��5ǆXd�[f��*�SV�hB��V�,u{��ˬ2��\�� ��Z��*��ȍ-L���'`�N�
��د-�xjgu�m�v�M���7)#bMו�����z��\��2��qa��5r�C,:g_�{����7����$���*�L0Z�t4kCk�,S���v�I1,�!'�Zv�q�(�P:$4��j�-0�j]Ard٪З�fӖ�AĞ���Ź`ZV D� ���'a�2�Z{%]2�=ж,�uiVD��Lb���59��͚�8�tT��Y�X �+$!�o��ό�E��
S�h�%h�X6ۦ1A�$�ȦA�u�e]aأ�ue�Ut��h�  f'y��G�������%�oA���c����)�YJ+�A��C)���J|�g^*7W�����ǹF�eU��1J� ծ��رb� �^�-�@�)�c{X{�����N�q���ITi�@�N�Z��kM*t«K6�)���e��]#�R�k5Ւ�2S�|P��d֪R�
��*	���Š��nʍ�WK��ܱWX��;i�m�ݕ��)32R���^��n��Vdx�6�YO6��
;QdN`85��Q�n1^1B mb׺+K��N��!^�6�U���"�ݺ�Yj�q<�D'-�V.$-j�|.�(�<TeH���d���Ufj�ͽV��q�8i2�n��R��n�AF\L��4V\���,Z��a�e����u��V���O�F��w�0�P�5I1H�
z�f����V�6��g]�����X��+
��©��l�h���Q�0.��Yt��u	ٔ�y�,��I۬u&�v���X���g�l���l�դM���R�R�t�7I�/U��Y��V�"�ilP�&��V5��:U�sNA�!2�C*�shS��Q�Or���5T{k��Wk�s!	)��,D��
Y���(ǩ�Su��aP�*F�2��N�$�X�E�"T�����lM3N��g]`�� �˷���JS@R�!�h��F�=i=��4����(ɳ$;0�Ġ�̀-�{n�6��S܏VJ.�ef])�����6����v��.X�ǘ
�2��w�!�Uf��"� �b2��}sWU��r��D�dh(
��<WWy��F�X�L�y(�,;`y.����哉�Y�!�V��yzj�;��Ťld��&����XWf���wp��8�2��k���r��u	$���ǈ\S�s9��)�C�^�7(��5r���`��yS+�f��++$��M��B�EH0[���.���.�Y��L�A��ja����,"���;�]];d�v�عf�V3N��H���8k37)R�����n9o"������mU�Rl��͉� +J�+�X���&R ��-ո�&"Ҽ����e��4-�W���V1�/f�c�U8E�(6�.M9�M԰be�]���Ib���է��k�h�����$�ѱ[w{W�����(�t�hAP�)��7
9�h�iL��U�L;WG\�/ij���(S���ѩ&h�p�ʚ�{E����k�������5�:�2�Y���q�bۗ��'HD�OJ�;��Á�/6�*�7zF]�J����TI'7f���S�YMRӹ����d�6���hJ���!�V��2�&��rMx�M������l�.Z���r���S-T�*�g �w�ȼ׹x���hf�G[s	;۠����bfko y�ZVUԛ�?9d$X��&��t�VF5��V�[�-#UTEڧN�Ȗ�ll�Xu��{��4r�1�@�T�-1Hm��c��-h�j��wpR4��an��Z��W=&�Ĉ����٩����RàF[�́�5�%�����%��M$�.�A�U2�ʚڽ��9v�n�5�݊�����U�d<唲�$-�{v���ݥW��P��`c*�Ρp�T^�Ѣ��A�PY���k���l,U�A2r�6��[I
�j�j�� �0=�4)n���.�XUt6�vS;�v౨��ij�u����Ӏ<��'��.Պ���8K,ݪ���vHA�[�.Z��$�VB�k�ۢ�:6���B�%���.�4����r��-��9���Okt�C��V�z#0�R�ƅ^�<��q���gk]�[�-2�7�f�N��XV���~2�h걅�#�r^a�mȯ����k&���bhR���Ye� �Y:r�*��qXW�v��Z�f�V�Z�� �w3sf=�Ԇ[ GRV�)7x6\��SW�.]��$�j�+�k[�t+qȝk���Ӹ�7n���d��X�f�&8n��X��7&f��m�Kfa/`D��+���7�<5����(cՋ~�I�c{Z�B�B�G��Ř%bz��5Ѽ�v��o�uL�Ѷ����"I� ��['��ld��0��kKYӛ{T�dE��@�������d��X��V��m[�h�ϐ;$��v(dJ�CU�x I�l�aA6��b�˔3֞��um[�z��$�$@���� �J�n\�
Ǘ�kY���H��öc�O�E�[���r˫���#Inl�/-g�wT�Y��4��Tj|λ�U��ݩ��� xM[
�]7Z3B��u���.�[��[�ݛ��Dc�a���m$də��F�IKp�c2j�P�k%�k33��yE�J�]���[�h�8�n�ڛ�F��1-�*k��h�23,I*j;�`�d`�+E`�:��e؅i��r��55�(3,y3f�
��-�ȝ�+D�Bn5V押J@�c�����7$�y)<pS��i�PI��Ȱe���U�a=�2��\Xʈ�5��wf�x3v򘚝0M��˱+�J�K�]�5���Eۤ��i��{�m1�#��j�\Q�mU��f������!)O�Z��5Wk�7�OeXE�����1���d�R��KR�Y�����4^��#XSzѴ�`
	^e	w�7��F��l^Ie���I
��+2%����j��/:�b���Ʉ��#IA����Gr�U�	*�T� �Jh[cݵ���-�tQ���aohX�$c0��V8b�,�uQ�s�Ӥ܈�����ys6��[�%*1Q��EB�-��-:T�n�փ3XOktm1{�"+��!��؊(�.�ׄ�Zs��x� ȷv��ˈ}
�z�8 T�*���4v�z�f����Pyw)��声eəJ��P�os^B���݉�rR��w���>tE8�V%]�՗r-�%����ŵ��Gh]�h��ֱ/ D+Hy�H���@�svK
��Gq����Y	7���&���36^�挬�K9B�y���)�Ö���'���ٌa�&��BH�n@a�V��a{I��6�L�ӏb�y�`���ik�-*�+;�6Y���: �2����)��k-41"  ��.���{%��)�t�wEX.1,�QJfA1�t��ͬ�t#Ks�t��YI�qKD,�K{kh(ʰ��N1Y��:�wY�r,@#�)\jU�L�1�X�;.���:��c�FC+U�2meS�sH.�ލ���Pa�f������U���klt+e��3n�0��A`�A%l%*L*�PQ,̗yP��g�M`��R;QfL�x�u�=�Af8������,�n�,�k�0QL��[�R�lY��v 7v,X!7�P��D[	9e��̗�57[�2��;V�Q�Wn�� -^D�gLH�ݫ�a�X42Pƕް�<��j���9�<�y*�9��l�L���L��~ە2ҡ�`P��Oic��oR۵�K6�:9,ޢ�� �U���P8*�U���:�M��(c��t���7���`^Cy�d����KN�X6�b��Nh�5���nJ2S�u7"�ӳa��`0uhNc�,�t�,��
�"@�P\�r�;�ٺ�"@�v�n{u���@L �F���+ѹ���W[i���ƀ���v�66����ݽf�Z:�������m�D�b,T#�D,�-^()h��ᨵh�q���6\��ͧ��d�jp*Ow2D֡�LT��Й��E�����T8B�;�Oʓi�,�.e��=��嵩��٨nov��ͻ�&\���N&ڛ�AAS㖕^kt~#�8�-}����X�NkӨe�T)���b��؋��/+�X�tb�W�I�����*��z ^^�%�f�5٠,db��b5�a�F�,��6�{6\s�`m��V_�ڸ$t�����+�,k@4-�3(�{��ܭ��ۇq������Zt��)=KS�^�1����71�L���=Z�q#������JG�۬{WV���{hE��Zl�	��S�["�]��h6Q��T��KN�^��D#9J�����e��2i �B��Z�pm�H��u٣���յ�N�e6v4��w[ 0Ti�(c���2T�$���d8>c�I`e�� 1KU�I��S�I�8Й7efmFDL��N�
fbWmdx���1Gy�VIa�wv^�ݨ7L	m<�X�MK���/e�&8�;��R&���R�q��̛�e`�Mn!��X��n�U�Ż�*|�(�,�ٮV�_��U��ywU�"1en�*�
5f�V�6��%e�M���r�t��F�iQM��AY�"kB�f����S	���-�#-�q�,T��J��4�*��M\�lH[����,�>��29�D�v�XE��5�����Î�Ȯ�w����+[p�.[.,NMѻ�)��ii��,���5���&��p���2ʗ���ʭ%R#$����%* �f���[�깂��JrY�B��2*۔�LW(����xJPYZ�TBXC&�r�ud�,ڣ2��,�O컖b&`&�P�h+�wG
읷H�1��(n��<A]ڜH�i�W�IV�������>v���̅P���\w3)�,4e��J��U�܉�GU!(2����Xख़F�j��գx�pm�V<��-N�V/%����9Z����eEPXǢ|ӀٱZ���;U�۩����Â�'tܖ���B���5��)f�M++Q�l�N���PP�:u5V,aջ́�K\+%۴6�h@Tk$����2Co�ut�觕��ۗy���mݵh��n�7,ԡQ׫j�ҳD�//��l;�\���O\�<1;/2G^��	�����*�@&��l�7Rt�X��mӺQ&�ͣ�V:�p��ч7n�f�n�P�b�w����"#[�N^�M������0�=�� Y�\�wR�.#[T�ʒ�­j�<�Pcj^��W :ŕ��		s5ⷡ�])fYH�v�N�(��i�C�q�#VGucl4@E@fLn'�����=3ZUjt#���Y��:�@�)U�A
.�-z���D�7�d��ʰkA���Z��2�����4�0�+��F/E=�l�D�k�kp�_�c�,:c˕�c)9.�3�ɲ�V����E�́��FGCr���+i,Y����wDJ	(�D*H�q3j@�^ZyQMV�,}�
��3��J&�4�B(��Cp^���e �h��me��K�c��nVnK�Vf�����e���ɰ+۩��S"�e�+.����Ŧ�3r��Ɩ�:B�j��ħ�<���-ɯl	V�AxDE��ʸ����V9�!�V3+X��!u#1
l��c�JL*��e�Ŵ�]��^�ajN��
�,��ޣ�sAv�e��Um�J�+n��5�`�w��v��k]ˬ9c1��ڒ��X(� ����sl�0��-S���;�푙wL�'#W��f:��p�I�Ҹr+�rAi� ��I@앖"�h/���ڠܦ�!�p`�aՊ�n���O���IVE��1B�܋*pJF:��4ƻUu���V�W�VO����Ov��@Yg��OE�J�����B���k"`��of�����jƁOv��)��l�,���]�E-'`Y�#�v�8�܆�(�bU�SI����y�ۇ%LUg��ܫ�����Z~n�ߚy��Re�쵈��P��=�iv�J{HƱ<آ���(黙J���t$jؖ�e���A.Ζ���x�yl��J��^$�ٖ�^�:3$xx%�i��	�L��l0�`� eH��o �9H���wp��xT�/e�Q�3M��W���F�i�R��2mn�����T1���b�{�@kfhf�]b��^��ԇ�&�,�C27�]	ETYs9����ׄ��[U�wJ�5�S��XK��n��h�K�me=h`j��h��.���Q�v�V��P4.nF�M����chK&:V�,�u���#BԆ�+�!VF�P���Zò%��WƱb�.��@�G�U'X�3���,�M�2�v���7@EKH���:F��Řb�IY�9f�Ee�үV۳�2�{y�
��å(���I��(�8i�����  ��j7�Un=ۡn�(2$����wN�:�u���*�'}�l ����i3��G7�K%U؈��Ɛ*
�&w����Iض��U<��qJ]��O��&�&f�ro[�oeMk�a������O��)���Sy���:M�`�/y��̮����� 8�k���`�L����%�q�D
X\���]fsLp홶ų����6S�6��w88�yNV��Ь���-��<�=.��}c�+4o% �k�y
�6/\�:��uȊaMw�,�Q���o�!lY�U���h�H=�uǇ�p��:�\w�j�1U�2c�k~���G/�֙���e	�#���\��m��L�qZ*���o>u����	pv�1���T9��*��L�FŻd��g
�a:��Q!Vd�|,[�C/ns�KI��T�ktNhb؇h�`L��Ƿ�Z�:�|�8L��ޢ�As��rU4F*U�|�΁�.�K�'�t2f�t��yj�6��.;�&�gGM֞K��-��W�6v�uN����Ĳ�Z]�WjW����P��|t�J��p��e]�Ui}�/�u�+���Jg*o:�XI�޼}Wk��'J���6�����*��Z�Vk�1k��͵��S<�]ff��N��T��3�B��κ��;~3��82%-��]{9��h黃(���*�{�(�b�i��o[wϩ>�90�e=�f���(ؤ3~D��;�r��F�j�eZ��T�p�a����]��
���c}�tGU�m]��kH�n[�Һ�rp��Gu��I���XU�',�u���xWc�j�c�Yݱz*��V;K��;�icą���׸�9�FPʜ�.N��1Q��f�1Sǀ��������q�z'b],o$K��vv>}��{�/�lsR}���k�P*����}�����fTN�^B�V4���vF�5P3����9&>��i֗/z4v�9�E�	X��k|H��˸���.�����Ћ^��:�b/�p���U���r1��ø���ǫT�uK�.�פTu�{3�f�YӶ����R7 ���vU�YܛO���r�8�Ob�wy���S� ؏}w�ފپ�Ċ���Xs�`��%��h]�O�W:S\�#��H�#�*��%����N�v��Rg\R�t	�epk]N���"(�*�=Sn�1[�ggh\�d)����eH���w�FŻ2Y�:xbc��{�%��J���x7��nА��}�񎜬Kb�Z�k�9U�*�nS]݉���Q���5oT��@8C�
\1����$�a�@�x~�R�oȆ���[r٫�v�l�]��p��
�b��Ş��6�3UDɥkd�Uy�&��� ������vg�9W&E����A�W�f^1@P����c��.��3J��Wm���Lޘ�)L#Ş���G�r�����
�`\M=8�SA����������h��y{�0Lr�*����'SYQu�q�MJ���ꎰR왃s�9�s86g+�[���fU�3}�-��F��Jvp[��V�55�k����8Uݠ�p4w`�=}�����ƷZ�-�YI�(�]��{�,b���H�ۺ�aS�ox�wl�u멠a��o\��kh�J�F���s�b��.gq��ճ���gGX$'���6�K�9ƲJ����F]c6�s��4; �,�ܼ���Haã����Ä$M�h�����J�A>am ��I��T��)p������{�k;��	㼰�z#��rm�6T�;!�P�/��m�-��etB�9��j��vq\��?Ahf���F��ٽg����j-��F"󮓷5A��_\�]+���ܔ��K5P���սv�\)۳o�6w�/�V&��`v����LZ����L��bU�pu��u5�ts:m�a��GZ��yV�\�1�t�ro�X��4��_���h�<��w[�>���\W-�e(�H�7�)1��}�D��K�d��/��n@�51��1�ǳ�6� �D����<ҤZ��G���wˎ�-v��ۥ��;�-Y�]�k�i�rk-c�O�z�1Ϋjv-���n��a���uI��IC-����$-C����L�[S�%����2��o�ދ)�R���ѼR�0Z�s������rmڻ[�64Nsb�~�������1lM�+t���-�}+�KvH���C�i9��ѹ�v�Ply�(9���Ψݣynok0�6X=a��g�ZU���*R��5}KI}�sx���<����0*\b�f��5H�b�2d)=N̎e��{3��׻�ԝ�W�*�$gneu�#/�"�q=n����N|�;�����%u�[]�ˁ��<���sh_h�_L�{�,��e�'��s� �w>�0�ܴ�'H��	{u��G��cfq�`1��6ؠ_���f��vj�ʶ�K�i����euSM�a��VM���A���!��e�tF���<*n<�>��%�-n�W=�:�#�Ws�M���	��A�B��l� ��9�ڦ���L̬��]�{�R�<I�X�P���+PÇB�&�0or�GsŭX٭bE�e�m��nu�WǮ�1�0e�ܱ����A7o��+
c�kR�B�jT�ă�#�z��N���=&qg�{ػVn�sd�p}
�Gp�}���$l�9���Q���/H=��f��X��7��b��̳W2ւ����c�뫌љ���LlZ �h�#3����m΢�	 &�\9N��c���}+Q�8 �� B���d7�/u��F���5�tp+Ħ��8I�|"��vy���*h�#�t���TC�:��c ^�C'���*J��E���r��-�]]�p����\$g5jl��Ϲ�'/�����^�n��47�Dz�a������7"§0��ǋ,G�U�K�r=��Ѿ�5��VT��g�=X�8{�"y	ޘ�}�B��]�ݡ��X�9C��8�]S�T�P̧5�kJ�@h��e�g�n|s��������fv��!�xD�8��w:س�7��kG%�[�yN��`���}� ��*d9�C�V�]g\ i�r-���)�{��aw'م�M�y���R��w]i�Q�Ar(A"��S����޲�dt8�Ӈi���,�̵LwI��i�7�m[QJrή譅��u�K��Mժ�u%�(eTL�J"���DŦ�l*�ᝒ��Ʈ�+���p���r`ޕ[�:'�^6_k�n<�ַ�l�zu�7s+��"���������w�`Vq��]0[�\oy.H��JVL���Y����oh�%U��n�F�F��`��e�8��Ȁ>�Y\�rK43�aU��Vjq����E,���o��Uާ���1���}L��ڜф�n�B��oS��[|��������x.�J�9���}u���B�����%��v�F{�V�����qh�Κ��ٮ.W��ry��1�T2����.л4��r�ڹ�]�f�Oy��sk�հ���y��K4�!�J�B��m�[����f���͉ͫrq���f5��sY�[�� j4��"��]7����]��nJUx�2Ee�mt�+�|���N2�۬2��z �w@�Aa2�}�JX�8&KY��d�3j�o�n��k��(��\|Ha��;5�ז,]�r�X!���q��v�1Z��lW6i��홚�K�=G�����ɌԸͫ�yQe�V��>\yۥ��ɚ+�*�������SM��]�_@/EܾZP��ܒd�0��D�9��s�D�<_'X5���Կ`�ߗ"	�<�F�����ۃc���Z	��&��t���*��/���c$`�-�#۲ܙ��(��$�n<�6r��y�'��{ �EwWpt���[�s�<��!f�y���{�����=nݣr\�]Az-�U�❴�Kq��s�Z��!�A���֥�-�O���"�Z�G�o�+ٝ�̱��G��{L�v�}�1M��i9�U-��܎�\�uJVҽ�%;4q.x�U�d4��Fj��e�Ӽ]���4�ڼ��ճ�ʆS��]!*P���&CV^�T�Sg}tDL��h���,r��r�����m��;��B~��B���a�6����u�������;k�(bf��8r�]6q��L��5�2�Eq�9Ke=����ʶ�"i'����$�F[y���b���72���Įf��Wj��1�bT1.�[��M�ܱS���c2�ŘmU����5y�ueHM�Y��0�g�����욒�2Q�(��U�kq3������H�w�R<H��b�9����[�q�����A��[cI�!f��]6�A}��lr�;&���aYtU"��8��9Q��X��x�[6���l���M�42�ܓ.�k%m7��M��o���땵�k��K:���a����8	������9$<��Dg,�ܟl��e�K�˽ˌ9�yhd�7�4m	�bg�u�=J��2q&���Q {l.������]+���ٚpMjXU͹W,na8��,����Y�7�紹݇���o8�;����o[���Ǿ��c��ΙB:Ot�9;���em��Ĵ�T�Έ��.F�G����_���^��}�`����@GRS��V�Z�{]}�p�m Qc�01�cf��2A;�L�P�dnn��2�K�>��3����x��m5����y�f뷖s�};+�p�*=42�cu�8h��ݍD�t���%�w��хP$��ѥi�tk��o�uf�}ݼSvл�t��atx���m�Ĺ�Z����m<�ir���zb�9W:]�5�4�-�%�N���lw�N�"pz�F�ŚM<��/���DCs���Tk�剀 �^;|�)���(��7����'V��	V�ƥ��j���aᾄ�������y'FA2�ۈ��e�]�wD:	LtL��^>�JU��C.cج�V�ai]�J�u�Se���)L��ɻ�v�^d	��.�HV\#� U���� Į��k�����,]䮀�X�3�E묗�i��68���V�,:�) 9�*��r���Med���ү_s_o�t�g*��@�;�$��{��fV�/%�9��Y��0W�j�'۪��{P�u��إ��$��Q�Z���C������)���ͭ�BS�}�lKwTٮ�L�mg�Okdu2�T���6�o*��9z/i���%Ph�U(]��:`�#.O����#�{��Z}C;�7uxsL�n��]��-��Y���M�mr��(j��i�i�X��Ϣ� �{���Sb�%���y���,V�=ev�H��k�4�wP)�,��yn�S9���ʌ4�e0R*�t=�3g�1����3��]-�A4����@�M���X�W-k��L�0Lݦ�P�ό�ԍ�Y�}4+,�c�2���S��=�\s���]�m��
��(_v4��fm;,�|9�A����)�A�];0��J��Ć��VG�����\5��C�u��	u9�<���^]��K�g8����F-YhĮ��6�̨|%�n��&�V�a&��<��lxV�E�4S��ٳ���&,GK���;;�������M>�@��؛���s��̼���gw��);�ђ�����\�*���wm��ɍ��N���;)��:�e�-��5�|�8v��9���e]A�}Á�N�q��7H���.�/`�y��{t��W�'�.�d��9:��V8V^i6u����0\h�v�&�ݓj�]����nr�0z�
���YN�el������sN��6�ݙǪA��%��Q٠j��}x	��p/�y���w�ʤ�Y�����y�>yt���0M怤�IA�Zw�S��o�ؓ�+|]� �Vo/i`�z��+�+��A�O�ȀwAk�]ˈݘ� ݞi�^���7�l�ђ-�{RQ�_<|��r<�_[l��+����>���p��u���ˀk�����A�i�=��;����ٓd��ݢ��Z�ӷ�:/73
t(پj����ƹ�ԇ���*L̓��>��Y�+�" G[�eH;�|�<.�ʻ����;bh��oP'��V��*�Ke�M�Tp"��'`�싶��
��}�i�e��2����1����S3iX�ͩ.�^#m���&'8n;���2n�e�:��ݴL�j�>�R������<�^���)K�ܭׇo4���]�f�n��G�J�ܠ�nCL��qƦe���[0.UeiŘ8���U�Y{�<�����ZT���e���'Z0"Ь�+������=�إ�h��f�T:G��$��#JO���j���M�e��JP��ZI���3*Ƒ��*N�����
�Vƫ�Pu��5t�zq��+	��vJ�V�Yc�o�L�.`5����mt�:�g��MѾ��ͦ���25�(�`n�Ω|l���������"�
�Es�h\�ZQ��ʣ���T&֡�w�#� �A.�9�����5}j-�7fC��w�WwA��Жe��]]P$1d��_^M�5;�o�����P�n�]��V�ww�=�k<E�Iέ��[vxj���>�����u��P��	y�M1�K��F�H�u=-�{:�ݭ寯 �P|E���YD�]1��⹩o�S��okѷ�yPgI�Pv�IB�uY����[SHo�ܭdqw��j�%:F_Pz2����\��5�H�]�3P]݉�ֳ9�s�M�K���fu0��0c�iq��D���'4.��97�=c%D+y<���m�h�Sdι[q=W��X���<l�as6�募�nH���=�^�x�TV�^a�3%u�Mj�J��9�.��]J���CYaufV\R���.��G�*�&�1
U)�{�Gfef�\;*.��Z��\��2,�φ�M`��-C������2oWr���z[��_4S�C�5w3Ԕ�ӿߟ��鵭m���f��km�����]�����7�#��XK��@e5G-ee�_�p��W^��a ��g=��k�0wf#�h�����Ϊ�GwN�=6�dͩk���D�m����I僔���(-��Kf�-���@�;�u��AN�e͢�
�7Uu�L��}���_gu(�2�X�г�!��
G��&�&N�G����'➛����	��1j<���a޺�z�(np�z�a�wB���W��JS��cu���qq���,������m+�ύo�(�6�F�u9<u۹�1�Z��������Ի��FwɋQ*x�J�f�wݤ���wwq�X�)a��Wcņ��*�ؤÝM;Ye��ا�m�
5w0�>�N�ܝa�K
��^#��rQ�+e5���RZ0f���jt#0��A���yG)���@�ޢ���VU�_��ޒ�4l����8����7yuZ=�@V��A9�[�e��jU���hS��q��� !�ܫT8$r�)����
R�򽙆�Ӣq�	�aM�!$��`��Τ.��pw�(�wNҧ,���l�p�_�C�f-�U)�7��q�yb��C0Z��8h��-VEB��i����>�or��5���g;��]\#��_m��U� ƅ�]C�[�܄;���v�H��t TgF�YúwGK�g]p�Oy��������:��)�;]�C4^�u�
ԫ�n]�$�-�8�V��0�t;�v��;F%�&��K59�-��]�:QrŖ6��`Qs�;���h*�%�;Tئ[\�v�m�I��m K�1S{���2e�J;*�f�eg��b.Q��t;��iF�*���
�|ຶ���p��h�lޮG����}t�"jYS�V��܎W&����Y[��W�������2:�R��	�#y�T'H�o����\<5��|��\*�n�˰)WsU
����24��O��8�}|N��XOo�-5�GnɅ���ˤ���gwwr堇W���<��ƕ��9��n;=�9��0����wm+���%�iÄՆ������t�.ùRps7�Kލ!�p�p����˪�Pp�յm�Y�,Y�9\r�>��	�Y��vh�� _oθ �[�r�����ڵSR���f�7
ɋ��{��=G.wB��&�n�Tf�{�2��f-krۮ� ۸�ifc#�����kXksW�+s-_vk��0
h)�;�36�]��ڗ�`y}\bN���x)��2M�9�k~K؁
�V���*Z
��Ưm��#gZ;#oE�Tܳ��.�h�7˕�\�v�m�O3��lj�9�ܹ\8�f蛬�cG`QªE��Rb�;@J%�L0����N)�.�"B�Ŋ�ݓ&SC��W`�4����ݛI�E�9��p��Ϩ�P*��5[��I�*,:���(�7�X�F](�xe��Z|n��'WR���֯��Y�{2ݿ�b�d���ɻQ�84s��3Y�{�.���K�1ow
��lk��6�:�����"#�a�U����ܪ�X�6��:�����S::�x��^���v��u gn�' y�FR�:3�~�á7}���>�4hR�7����F
;�0T�sJ�GTkZ۝K+џ:��Nc��X��f�U���t�� U�f�R��y��ݸ+HI8Ợ�ݳ�*^�;1*��Q옭7\�e�����0s���U v�އi��7C�W�T�zր3[��.�5��v�s:�;�[��b�Y�x�w	]w`*N�Ҿ�o8���T�*c��������yV��ӭ<�Ny_T.�q���A\^�c=���)s�yе�Wk=6�U�!},��1��^bZ2U��-<+m����i�+�!YC�o�S��a�U�e��R�8m�K��vZ3{bB�qT�[������n���zo>�]�&e�ΝZ���<� F͝b�ﺋ"�5�k��)�uM��ة^�9VG����!�$�c�[[��%q����9'�p)�az]$�N��@T�;�iu�ՉY}2��	��p���1�=ӐA�@�=�������f��U��\�,�1�3���ˬ�6朡`wuW#�I��y�c�W���#cm�+/��4��_[q�䡦Ձ��"�Rz%6t�f)���x�^Q��]S�|�����r�b��-�p��-sB5]���������'.h$JX&��]O(�O�V-	�IڏLe�:�	ɳ��]�ι;,����eQ���j_%}�ط���bB�uZ�E�RΤkFɨ�Ș݈ep�7Cl��i�U�����y�6�Vg��,e�t�Fh��8�ɰ��Co)�|�p쥷el/N��̅9pEu�M�e%q�;�4w*w'K6����z�v��K-"�L�e��+mn�1]�Ʌu�ʹ\����tW�e�J��f�EɎ�W�,`���&^J�����U®cܳ�IK�1¬w|~�*���񗔖�u��
=%�'����*:bô��|��̈́vp:�b�ֺ odB�T[ ���:����F�\�,3v��F���}�[��O�bd*�v��!��qа)�v�X�T�7P�}��U(5ջĎ�I�7�'gj��o;tK���M+��Ŝ�������������h��ά~�����0��\4c�y��
�
�M���
��i�zӘ��Z�*�®W�+O[�9Li1���^e���g^��m<V��p��<��a�oD�8j�'�I���yZ��]f+]%.�3���`�Gl��]�@ܠ�0,�e�;&��@���nSCZi�t�M((�{�r�4�J��L�W)�4��q[��uL*� �'���t,�y�ZX��G0.H�ٺ�������f��RPS���-a|�|7�ޒF�@�t�۶�c�m�M�0=�g]Nkxܑe$-�ͳv�c�G|���M*K��>t3^n*��hxlm��hw}�VrYw�麾
���7��* $�C��ڳN釴;���w�N�&�d��կ��|���G �B԰��*v��J��>iL���iݘ�,u-#�r�"����\xF��!m"�y�ƶ��\;���Ί37�̀<N޻��VV1`A
瘸l�:n# �y���Zh�G�\5Eu)�ۭ���ֆs�\�Ý���
>����b��@ǭ`ƗY{y��-��V�լSƇr}��n��eُ3&u��^|)����j�>ٽvک�f>n����'&x)Rm�Y�1�N$Ȋ���[h�|�V�P�xz����:���t�oZ��<B�;؝*
�w^vp����)J�r��NKl�5�RM;�j�d��ܹI��&����lv����iEK�x&�aOŷ�3�`��.E
i	k6�;���X��p؝Ad�J��Q��Wjݹ�ˏ*�\�1+t�=2���w��nc�"�{(ƫ�U@2�v�-mm;���R�)\9,�3�x;2�ͫ��)ئV},�W�Эi$s���sWh��zu�ЊwwSͩ���TTv�P�ZW�������7z���ζ��;��fZ�7���ē5�u��xÃ�<��,9\��(�<�9*ER��پ�fKb�Kԓ�kt���c�E]v��4�q:Yuy� w4(k5��:�_4/z�᷋���T"|$�l`�1�εѶ-�9n��>Θ�#E*���y�]�9i<s1��l��[.�%�)��T�	
�v�[{}[�+�ҡt�A�D�k�a����@e��6[�ޮ)�����9�*�+]�wӻ{dܬ�鮜Ƞ>��Jq�8�{�C]�;y�t�Z]WPU� v���=����(!w�ܰ���	�g�v�^*��}j@�m%�4��ipbq�r���5�<�����v��1��h����eM[}{Lv1O+�T�{�y��^]dGpʕc[�<\b�&��ݺ��d�ܼ�-"���!�`���)�j��*	\ӫ�:�k:�2��Hh��;�����wGmf�fv��yB:���ڙR��}QC���� m�s���g&R�k1e+%l�(���x9��]=�n������v����ަ�+b2t��4�h�,����u0C�'�x���.A���p�{������$-j�`��&c.^�#�Ր3�;3kp��Sck�r8'�\�A:�$*�۝�hH�t࡛��v9� i��ڛ�Ω]�7���I;%��W�/h��E>�8	A��j;\/b;�;h�b2e�SK�n��-{׵����^�5z�t��=�|���g'���[�6(�gk��vZxh�����V�6ƉLn:3묪����� >���K��vu,�Rp���MH�fTq|&j���i���2���t+��D�����p�ӡ�N[A��Ơ���;���V숦�0��a���Q�������ݡS9p�s9��J�K�Wn����CY�@&󝅳�#��Syn5�ll7S��ՇmvSb�=bN(�R|���t�wo�x��8Q�XM=7!mv�}Rb�+�3U�ö�mGC4�t�P-\��uی[U|�;�xT�n��6�ΘeY�,�'ֹ�F��@j�톆�ΕY���ΦE���MR�����o��h��a�yW�V�1�O����K3T6rF��]-�՝h����#���e�@f�X9A�+\��Arx��(��+\(쀅 Q9�mu�\�f����r���obkF�3B����ب���^�T�/��y���qN�lf�o��I�ۃ�g���P��xf�g	J���$u�z�s�tS�0�T�rI�
�Me�u�(ۍef��]l�i7�#3SYET*m�3�lo,ң�V7Og�eS��o�3Gk��eLdB1u�Ā��A����3��y��b�,��2����N�{��:kD%�;{��s��Xk
�>�)��呔�r�Z\���r<��`�!�w�]pI�dU�Gh�J������*uvm��U��Q��V!�o2�Hb��!*�^
NЇc�7��Y�r⭖�k�Ts.�z�<��k�,�;CX���ή�A�*(�u��i���i)���������x���tbH�-��x���kl"�Z��0P��
V��}a��0VV��:��T��pk����R���:�ҳ��q9�6V�W��Z'f�b�c�_s�77S�QQgdư�<*��Vf�D��̸� ��-�����ᭌ9��M���u�t�O*�(�N�!l��>�̸��|��P�:��[��ʛ1�{tm�wYǛ��I��dj�b��H	|nCt����՜�z�>#��*C7,}�Xĺ�R��p�:^"��^��sB�T�,ٙ���kI}Xœ�/8.�
%uǮ�K�EU� �������l��t�u)Ía��*��0����rf0�ɪ�J��U�e6�P!�K��u�@R&�(��)З:j���@�pNK:\{m������Q�I�rk��(��9;�<Q*E��,U�u��y`�쮚u�N�&;�z�0�j!{@�[4�\�l�Z]�j��h��D�ck�]y���2u�q�r��Zd�Y���
�XT��3RA�7t����v�r*-s�m7asWu���e���{�Um�ˍ�[�8�F�K"�DU�T�)A�8��y򡀢�ev��F���.S�����7�(j�;�u� cT��.��t)�t%G;.h�ǌsA��e�&�%�I����#&��Ʊ� ��T�ʔ ��c�i#Fo(uȭw�V��v;)��o	G��tNkc�%���S�c",��ޖ@攕�\�)V���2��>����9�,��
�%l�Y�t��R���4�[�s����d��
�����{u���
{π��x\�h��t;J���0oPы O����`��r�KuY.�L���B1�.[� �S���፼J��A��;��:�(� p8	ݺ i��|���rW��iM"���r2P��&������츕X��̪5g9����j��ʲ�ٶ�������99ƅ��v�9�>.���+ҵ�V*7J��c��^�Z37p.I�Iӽ�j��C��[tЮ�B]�Uet����
�Ko)r�ɬCW:S��-�Q�bIW*O�m����r��켹6Ze��ҖnGPP#�iu٬5��kXh(^�n�� 0��aah`���Դ^�Q����	�YHu�3���B�
����kk{��L��֡pr�ޏeiJ�CYc1���cI��Jt��m�6;�$ˡ��mdΰ��+�[+E�tN�,�j﹚&�+�W��s2]��c��#�f��h ����6�V#�\Q�����F��	7'c�E^�G���8$��k���ƻ�����=oRf���`��ءr�Y�EIv��4��9�y�N���-��[b���4��Y���)g�������]�����X)���`C�g3��;�HK���V���&M/�b��]��pj����ˆq�۔%<��S���)��rv�CZ��y�eڎaMQ�p6��x����ݦ�v+���9���:�����8�T$ebj�a*���v���0Z�]|Z�q�S�hlW+��4冊y�N���O0�M�2��ɣۖzL͑�W>w0V'��h��T���������|x=�uv*��"���Üph}$��[H�P�42�`�&��Pu�@GWx���-��{H^�EN����D��2�׼��{ڷ/����*T��hN�#S��t��}wn��X���_R/�@��A=����	TBnY�����ִ�+�˧-��8�c�쭰�E�=�:ѓy���m���ND:��zE�ta�����/(����ɓ|�vU��脨v$\:I�EG]����nj�\{�ι`��w���`��v������wo*�;t�B�B`�ސ�k;p�M<B_8��+������U����F���.ܥz��N"�nr"��������������5+g��j��+���L6��h\k{���
�@�D���S�́}�*Z!⨍d�&-�]։�{q����iur���-�ݲGv��U���(�MS��Wf �N�/{�;t��g5�'�[Εf+x9�ϻ��2��6�)�\��[&�ָ��k'WyA�cw��E�[`�9V�w���p��;<�y���`����)RC���_hu��dZ��,SeCSC�˫<fb�2�u�3�^�u���v)nP�_r�Һ��J�]m����Xt� 8�
����˘���җ4��
:�Sfs���)ͱ��3Ry�c�p�h`��ڻ��ǲӧ�y���
�����ӻ��ы�>+����/4ξ�V���RV1�j�v�c����j[묈t�:���%�ƴYT��*�G�zɸ�"�Eoj25V5���u��1v�\u5Oc�Y.��6.��\J�9v�&��:��󺂇z�%���eM]�nJ���9m��o;vg(�+�4��\��tfʡ]:]m5g��w,,wZu��r��$j�n�-�t�BN�Z��̷tR��+4���sNZ���MY�����aL�J�8���*7���we���sY�T�¬h�[���p�M�f�V�̹ť\��Di�	�Xv���ޭ�j��4�����5���<��{��0T�.�ZsJ�ޝV��/~�[C�@P(li!	&9�0�wu̱��
�Q�˲R��Fh��#Nt��!�:뫺�� ����A.�t�$*N��$%�vAs�;  T�&d��E�q$�I�A�&��20��W-qM�BB(lɢLGwh���
AMp@���60�M����c&�B��S��9�J���2�� ȂL��Ⱥ��`),���`�M�wI#C�w.�26�ėv�DKu�d�˗b$B%%4DE��H�#��@S&2)Q�ƀ؈�F�L�nI�"�6$��Ȕi2�̄�B��p�4ə�1$B������O�����~���e�R�S�����D��9�si>�YZh�S2�RN�b�R�}0v ���F�K=��F��:�ݏsR���c�ۼ�0h����t�,�:�v+�ٮ��h����R���� h�#؝���xs��3���D��|�٫�\_X���6�����:���6��7�)�Ȱ��\V�1�:���~�������"l��J�xV�1p�B���Q�\����>:�o��#����x�;!���������zE�룳S�U�k4�D\44�FP!C�9	`�u|-LWb�5\#��D����[�`q���p0K�G�����V��N�����r� ��8Wu�y����Jc³�T�veQ~`h�\ޭfa�N�.�;��٥Y؄єo۰N߳=����L���{�_@�'s��5&��U�qwq�[&-��9P7{R׹��x�[}ޱ�ш6,OR��dh\�I8]#�,�5��K�\USw�u�t��v�]킹-��W�]�r3�o�� �.7�N�T$t($�	�"P]S(���e�wD,�vB�9�>ζ���;޻|ps�e��#`(��XQd�*��7�{��q>%D<̼Y���`�b�á�wm�V��&c��8.��OQ���#X��s��2�yK>��K���\��V���B�S��1�
r�R�
��z�	��3��|�Xn���w�\�vo�9:A3)�	+y]ˣ$+QOP�{J�|&��QES���Ȼn!�Y��Nχ������:ԝ=`d��2�*J5��w<�q�ɣ�́ٲS���D�F�1^s<��S�(buѱ�ڿ\;�Q���l=v'M��}x�{dI�v�k�����.�؄X���x�"y�Q�]#��hb�Vlrj�'.�"��yG�;�.�=�r�,{h�WP`�^��bem:6:�#՞�~q^֍ݕ�$;R�n��^�fv�y�2K}ƴ���3�gO�9;?I�>j���������x��oR��x�>��ި�Qju%% b�.ƈ�O�B=4J�8�Y�S�|pI�9�.�`ֱڐ���y܇���XX��Df��&��Pu��;�/L��������������uH�E�l*�XLf}�Q�㜽��S�D,���u����8P���q��5���	e�b����6��O���*C�� �gZ���!�ygQ��Y���O	N6��a��Q�b4�,?�Y#BJ�\Nd��l�����QU�I$��aDD��L*!�g�:���(��<�suh*���t����L�
Yuܔ���E}���f
w\U�R����zMYY.��o�xhGZ۹���f�d8z���vӻ�ӛb��hģNL�0>.h̾���5�*���[�(.��L[#U�s,�Ĉ���^�����Iʵզm����ͷ�{���vˣ����+F�3��\K������Df�Tѿl˅�.0��VV��/�9�1|p��-��w�`�#6á� ^��ȻRI�4zPKG��*�v�.�(QxS�Y�d�܉!�u�cK�ˈeal�y
n��E�; �R`�*!X����ٱ�v�ڼe�#b�4�|}�mx�"`���ǯXt�09��mX}�q�P�+DM����~�~#��x6ߢ�I^ ʈ��LŃ�6��K�M�D��\�Ȱ�SD`}'Yq�p��΁Gg5�"����-�.N��A��@)V�d�e`S�OhK��c��wO���ْ�%�L���'��w|���*� 1?>Ӏ���+2H�i�i���sV{�	�q���>�k�6@�7N}���6<۾��� �%q�jR6H� Bg�P���cz���R��s��S{���ћ��$m �[�a9����%�/ |�$��C
��o�T��ɗ�����ڍT.iQ�E��^���a�s�REy��ɿ' k�he��I�(���·����˅̩�N�}�RǞ����ڤ�Q}Y=5�$�8��.CIݤ�+U��]7F/+g���q��e�N��'��tu��U�fe[��9O(��.�(�eeb$
x�����z\J�}3e8��=�n��uw��R�3{�,'��>K^��T�G/a��:uZ�_ʭ��Q�-��5��Q�\w+��3Q	J ��>_�&�G�L[�`9g��7�5�>���Z�׍���!V��ER[�kVz�=u{o�${z���gd�ԟ��V^����LHj�`P���㙿�
�YM22E�Jf�m[��՛e�����7�E�œ/�y#c��9c콎��������G�ҝ������Ù7֕�e���d�׽C��"���m_�j�,W��|���%���/�ܮ�[�v��{�ܙ�7ꆧIq	i��r)�
t��=�M�����}���E)�KA����:.(���⠏`SC�0��
�
�BE#��B�@�k����q.�r	����;�՟C@V�?w�Z�'���bC�5� ���;�
�]��ki��"<-�V��ӨeG{����b�g8�J��B���+<��K3O��O�T�TEⲦ��.�_d�H��z��6�jF_U}�'_ڀ���x�U�Ow�_83F�,��s�Pfq������%�iiL�\�-vw	�q��V�E����:�B�dA�=�=���p/V+%K�{�g���W��u���h<�(�\w�S�u_c/�����w8�7��� �����3���dp�[��c��kywJv���tgB�W�]�	��.�z���.6.U�s*9�.C�ӍɁ�m�+��O�R��4�^d*���
{׎$-����l��vڙ���������%;l�&��p22y�Bu̳1�${�����?jf�>�>����������욋�Pq�����]n`rՖpA�D�ׄ�T%C��{i�M�IJ��U�4	�'p����&l�1Y�\�됅��?W˺�+��V�.[=W��})z�odv� A{*�CV2�����t��g+��k����e%�tn}�BΟ{7�篳�pAf�����>��x�t݅�Pl�:�7[+�GR��D�4�!����޹�E#��{c���{������~��L��z��>Į|k´xm�-}�G�w��凧6�zwWM�ГVO�R7�j�jd="�N�����*���ipl״�FQ
�X��^i2�1�Q����D���Ԣ(n5��:�a��s�����5�K�1��L�]���^,g.���me ��WB����Y�f�	�������r鳹J��j��`8�٬Ŝ���I��bV�c���^b��v/n���g__:�C�0���������G�:3p��h�Xź����`cnA�֏"�*�;�����:�lf��<�^5.��IQ�6�L)
c{z��x8�Ltm�s�u��j�H��L��t�]C�vb�7���k�dY)Y�\O��
��jNҘ�����X��z{;�����b��� }�Z��~�fا��G��o�[��r/p��6eW�Ӳ5�((�Į�a�Κ��M��^on�yq���-(Ya�ȱ/��ڷ�eP0�U��'\��u�c|kÞ�k�b�I�D�6���eu|1���۷�9�_�g�aE�h�
O���}%B���Z��z�o^�q��}~�U��7^0��玻��p�.=��TT�t�,�Y��c�>ԥ
����0đ�LP2����tl`�����ʍ�븛��bt����o��)�?z���qu�G���:�41X�ءɫQ�ˮ��\�7���5��Тw([�z�!ڡ:Adu>H׎ɉ��딏Vr�8֌��V�IH��v���OO
��}��A�����}Ƭ��)֮'��GW����4k|m��9hA1�3��Q�n�{�~��	���2l6�#�C۸�"�2:B=4�Q��<�S����X=���Vb��� vqt��mR^�`��	��I�ܫ�6R�'MDc�
�V-N�}����
7hU��ʉP`c��GC�Gn�5w\�
5�K���(
F��'<��̤.y��Ka�jZ�Ju�&�;�r/�]Y74�r���{�9s;CP|��|���B���D`�>dչPv�w�o��8z.�>ƫ,9���G�{��U�fz����"yN�4nʇ{5/�>�������k�p0�k
`����̃ݦ;8z ݏ����`�0��XG�DEn:q����R�go1=�p���m_���<w,���C+����2	)��!DB�'�
�ޝ�8��!.1Y�E������׾�轜�(QD��U�v�X�wrlu��w����� X�����W�؉�`�<M ��_h�~q��3m��5'#��bIЪ���˾��X[v��%\�C��#�.��N����l��ߝ֡��3���U"�M��-�/�3��A:��V���vD���L�ۏ^��F`r!mP{��tH����W=}=��ʍ�"����O��,�2,􄍅�B]�o:&,K�\�B}'OB �{����N)O������yYA�\�5�
$�i7�G2�!W�zm`�����or�2�c�-�"����ux�T|�0^�vT�;�;����^s�RPF���e�U��O=p����;�|	���}J�Jf2���Dwm�kSH��o���g���>tz-c���_V�-�Hkuo�����q]�Y�{���WW�N-M֭shCY�WG���D�J�b!8� R��j��A��](:��/���,��2G��T��]r8�rg s��m�}a�@2�+��R��H�	��I�h<u];�EwsN��i�LyLߴ�#k����1�D�%lq��o�dW�`a�9�=M�{��TQ��ɬ��<����=!D�z���/z^�Nfz*H�4��&��T�xm&<F �o@�;b�z��դL�B�:��}C"�����C۝w��UCG":f��*r��b�r�o�'��D����S����#$>��~t������^��vx`�ݯ	�oQ��վ������{��ٖ!SԴ@p�4��=�����7�f*�o��# \`Δ̖pV�P�l�*T���u}�	���>�J�\uT��?^
�s]j�6i��*��c�����7��O7�^Y;t�,�&r�-L�"�VT�d�������4�ddW98p��&js�v�Bt�[ul#��wT��`�CS�2��4
�)�=N�=�=5M�0�>U�����/Q^ͷ`�^�a��V��a%��һ���W� ��]Omv�Ku�1���i�8�(,��hr���E/�t��f��
I�b�㽄��V6Y[p��F�
*eL���i^v��v�ٴ����9V�6f�J��ņ����3�U#���P)(>�w��M�G�*��V�̄"�:����taU�jp�JR;�l�r`����	R=&�^��|������ ��>�޿+��6+�O�]�K��W�{"=¯ex��<��Sv���:���;(�;��|B��H��ĳt^�cRU땞�����*��/���8�{g׉�o�`�u֠٨��L�B*0�q�u�y��({q,5k�����֧bIq�x!�i�6��Ozr��� Em�o��A�a�gVJ5��-,]0eFv�*aP��utvJv�	�).F@�6�NX��������D�bM��ֹ�W�N�&����[��peò��k�[�ڢ�Z%[5�z��Waj�i�t&��UrsD���`��D�BNÓ6WZ7�C��\Ë�>��JY-B�霗�éq/Y���l���V�02"@N�������`��R��N�2s((jYh,�*
�W��ê��+��4Pˈ������D��z�-4rn:���1��>�eק�Qx�Q|F��t�s�V�A*j��ٯ �c%W��I���~�~(�����V������o�,	D_��}�{Z��b��۸�g}��y�]�emy��օL�a'�S篫�ï�p�z�n�Z�.������H����m� s��g;�jJ`�Ћ�WE�r�i�~���5�x��0<�]a����b���k´/�\6PY�h�[��$>j�Gީ�v\�ڷ�9��L�ӯw��H�Ӯeo�݂�oO�h�q1rmjIvnVѬ�ul�}��9*A��-�j�.��/�u��K�G���ݜ����=�i@�����f���&�����Ux}�<-���5���V�#�U|�H�P�9^%�hl�grH�m}=^v~�Y.+7*t�d���8#��5'+��Ү��	:;�=�<���k�Qd��-�^z<6�V��i������������*�/p<JF��¯fޣ#�r�� ϰce�ӃO�,���d\�N;'+c��K�<	8�K�T=��jS�K'z�7��j��.¦w���["	����[ボ�V��*���7ǯ�l; 2�&�ǧdw�~`����C˼~����)��[=9봎�����q�d(
���u�se�ו�e8Q�"d��Edή��8#cܫF�W��eF�;�ǀ���`6㹡�ywS��v�����Hm�s,��ҧWh%æ�'*����;jN��q�\�<�2�:e%������:U�䱜ם[���^����\��|*���� ��|8Nx��k�v3���Eb��c;��	���6�������sc�b)���M���\(><���BK��_^�� ��_}@�����uw��y|��[X����5K�5gC):�y�x�V��Rb�1�4�gX�v��1x���T�2l�qn�V��)�'P�'WVU�n�A�^^�S�ރ�wJ!c�6�H�)��XsE��݇�Ov��(߅�\���k"sHvb��V��f��i��V�p����ᬍ���w+|�7Wt.�����QA�b8t��CV���}�T�(�Spv�:������:�G���:����!A��[���ր��|&��or\�>5i>\�C/��6;���hw���xD��/x1#���^70�Y�Vl'tCx��l��՗s�7!w�6Q�u�F��)V2����3�k�������)�WIMu(g�����sA���y?���	�Ǻ��m3���.���j3c"�z�K�<�޴E�34O5:=�Bx ���`���[T����G�<�ʋ|��WWAV�Wu���$ <;0WvP�V�h�K;NGQL)�+�8(��^�^������@�2ʣ���W���tmXȕ=��� ����+z�xsZ���ⴏ>V�'��i^Drw�7Y]O2^��p�L̕)���ߢ����}����Z�"S���H�pv�H��g��nS�3/��2��r$S=���v󝍣��������+�[{��zp!k����f�N �g3X�#s&�1�C�9m��1����'�;���M41��4�nk.��z��&ܭ�R���񟖡���8KX��Ec�z��Ԋ���cYָ�G6�f x�:�J�$#bǋ,�l��a��ض�S�V0`];���8��ZM�so�����i���8]n^Jғ���.��e�g5�Nכ)��z��u٫����R�~�g�b��Q�C��Sf��<T=6�el��$Kc�]��V*3�2 -�y�u�:��Ė���>��k���G��صu*I��)�N�C��[�i�4՛�7nb\�N���p�*�w�eTMҺ�Ǫ�^�"����+�փ�x.�%���So#hM�<���]�}���K�\8��=���-l�S$��]�eI35N�C:L��]�۹��n������I��Ԙt�jY��S�7Rҳ]u۠Z� ��as9[ޒ&��}{I��n�ϔ��7)>]�w&p[�ϫ2��0��-����YJ��d��T@T�uֆ6�@q�q���gm�*u�N3]8���s�4ɭ���g+��p�5�d�E�f�K]W[7�F�QI�]���+N�{p5�d�������[9,��m#���w��#���ŕ�b�F<�9}:��z�P�B���W�`���I�L"$Y0aL�&"$�� 9\D�aI3Q�!�2̆(��F����#F1d�̠�HL�茔D�(JF,.\F3��R�d`̥�RR�54$!I�&RS@LJ ha%��f����7d`�31�J4�M,�ɒ&A+�J2c� ���`�)i )�].�d�D2J!dD$�H��&���1Q$ l6@�1���I���20BI��sp�(��f�1�,�I43D&`�h1b66��@A��)�wt»�L�Q��PZ
>��� �*�N锪�$�ӥ��M���}���e�K���	�8���Q�7�>�����j3���F�.j�,���el5��җ.w3��+��zk���'k��Z����+��x���;�s}|W����m��h��ｷ�x���[п�w޷��W���__�?=�ܫ�r���;=���"+����4DI�+�ݮ���{/���^}��y�����/=�>��k�~����_���ѽ/�;O:�^1��.�|����y��o^u�o[��/ֽ��{^-�~y^���׋�^�����Š������i��&{���"4G�,���ז?W��6���W��m�v����K}W76�����~+�7�=u�+����ݽ*���F���m�|_W��ο��5����{W�n��~|�~�F�dM����5�:��p�"0}"/�o��j����o������W��k��ߞ��ޕ�^�>y����^/�x����o��\�/���w�5��[�\��x~v�/�o�����6�^����zT!�&&���0�{Tx�>#�m�|}������x5=�_�V�o���Uߝ�߾����x���~o��h���|���k��^-�߾�lE}^+���>����k��������~��^5~w������[��DL�0���^���,��]!_[�����W�w_�����ֿ;�C�r���yu�����r����}W��o��?|ץ�+�[~_�����ֹ������{}/�ѿ~}�o]��x��o�ޯCR������2K�:�}�,f^E�*=�n��\�~��_潯K����7��^/�߾y^��}k�w��_�x��ץ������wu|\ߍ��ߊ����ož+��w���ME�����;��u��	�T���[��fA��Q�e�L ��F�����{m�������Z�5�����^��n��~_�^��o����<�-������^փ{޺�W�������z�������מr��x�0�#��>	�u+����^r}���ﵿϋzW+���-���|^-��}��-?��������_˥�v���[s_��y��zo���׋|o-�]����zo��7�ν7���o����� Lx
s(���.�^|�B��O�������z�W��k���y��V��������y�7Ͻ��z������Š�����W�Z~u�o��W���so_���/�ޞ7��~_�[�<m��^��� � >�ܧݣ MȮ��7�1ւ�����ۖ"o��3͕��5ۙ�nG�-I��	�G��k�j��=�,v6�h?@�/���(H6�n, r_ڻ�P��� �f�mr���>�n=���!�{*ݹa'�*�|�G��G-2�Q4��d�2'�,�P�[}��
~��zG��(���E���T
����_[z�oϟ|���o��{o�����y��n_Z�|[��}�ڼo��^/��������o��c��x���Θ�#�$G��菱z�3M�ut�������ޚ��ޗ5~�-����W��yzm��o�ߗ��筷��޿���[�����[|U{��<�|[�o���W�o���(�������	��Dr���N�g�������h���[�\��z�~��W���{�v���湯Wy���[��ޕ����*�����ϟ�~+���}m���/��mʽ.��y����m����7�^��yǦ��|3��|�_�'kq=A^쟵�����ok��]�ֹ�[������/kF������5��[�u_W�z�w��ε�ם��oo��/�^y������[��n����o����|����@��"�!��9E��{�ۊ�����>��7�nk�ݽ�K�����5��^��W?[x��}��k��+������{�ֹ�7��^�v�>/J��76��|x�}m�E~��ϝ^���y��������D1hj���Z׶��o�gQv#���׋�����^�������k�^6����z�ur�����ﾽU�����y��߾}m���~o��_��x�o�z^�x��[�^?<��oJ�><o�:�sn3���)�t(}�ǉ�7P�ǂ�\�������/��V���ݫ�����߾z��F�W�������[ڼj��}����徫���וz��}W����^��5��|��~>-��oJ�w�-x���ǣ2���JS�}�<hFh�� ����������ܫ߯�/So���=�y�+��o��/��6����x��ϾW�]k���>����{oKţ�ߞ_����^+���-�Q���woKO������W����
���3W,o�>A��>�
B������Ͻ�}��zZ7���ϝo�x���}�6�7��7��ߚ�����^7�����\��s�������h��s���ﭿ羵���ͼ�������y�}�|�9�wx���\�6�~c��$zb`}�SM�m�G�������6�:����7��^/���h��_�z��W�Z/~�������k����|�叫���y~*���[w�����6���sy��{���K���Z>D����&�/xԴ����W:17�V^���[���Np�ޡOv� �76M	��|��ezf�dtk���p]�dvR����
ݚa��:����Ֆ�-[����i�¼�;�������	2nn	���5g�wr��nS�:�+�LN"�i�S������6��c�q4G�����r����W��nW������������o����{���s+�x�~��zZ7���������~o~�ކ����￟�}�����<�ן꿯�c��<�&ۗ���1���5���-������������|^~}�o�{Zy߫�M~/m�m�z����6��~��o��;o�xwj�7��`G�i<��o�b����/V�ƪ|�����{^5}��^zo�|^5��_��וz_��<�+���m�_=����ռ}m���Ｔo����޿/�|���Z�5��[�^*���޿x7����>�P&=퉏hau����_FW˸ߟ����������_{�K��[������ߋ�޵���ߗ�������+�~��ޛ�n�����߬o��U��[�ޯ�n󯗿�U��x����~��˖���W��U��HW�ދ��b��Մ(;�w1����ӱ���E�8'r���^��zU�s~5���o��-�\��痦������~��+���|���}W��mʾ?߾}��F���~}�E�{k�\7�߾[��W�⿛翾���>���W���i߇T}�<{`�����+�x�^����{oM�^5�~v��r߯U�b��[��6������<���=����~y���������W�ߊ����m�{o�no]�ߟ��0T�|��.��٘_�Dz�X���>q��{[��ݷ���>��5�߯5�^~��o�o񿗍���x��x׏�����y�}_��i������8p=0�����#����pS{4�O���zq�$T���� 8�u�֌}�W��߾W���o�k��^._~�}������+����K��[��ux�����j�w���ݷ����޺��n�]�Ǧ7��-��������}���>�7���[���=:@��ǽ���,x�@�׋����V����y��5��_��W��|��n5��?�~���ήX�^�>����7��/�^����Ž/wν7��I�H�D0{�%"��>�YMOf��}�f�yh���G�?�ō>���������p��Qo��^+�����{��\���z����W�}^-9�ڿ[�����y�ʽ��{���꽭=u����׵�����.�>��K/0�ȃ?���K�5{�����Jfg��xX؊hOY��""�(%�7u��V�����J�[{p��A�;� �ru�fb��Ď�ڰV.��l���o+��QWp]:��\�c}������'v�c�p9����x56�uB.��M�G9������M{>^�|���5�x������oj��>v��������^����ﭿ���۟�ߞm�{�}no���[��U�{o�>�z�E�[��������ֹ|��V��k���k�f|{#����q��#���}Y���1���x����������ow���~�[�����zZ7߽�˺����+ţ���/�����^7��m��_ͼ�~~�y^�|\����~���ޛr�U�����ob(�@����5W��s՝;=K/�Ҿ?�x������鿛wv�ϯ��<��wu������n�����<��U�y�s|_�y�}[�zZ7��|��k��W�k����z���k��������#D|��\��>��n�M�����������W�s}����o����o����U�ͻ�r�{��=-�\���Ͻ����W��m��Ǎ7+�v������5��W����{�\���0��"4Dh�|r�������(��o?�|o�~������o���ס��s{��y������~_�>�����m���Ͼ�ms\��-������~+���o�z������_�^}��ޗ��-��⯫����d{�� (�������ļ�3����ߝ����7�����]}{[�]��_����o�<k��^/�yW�����_߾���kA���ׯQ_W�Z~_~}�k�>��������Ѽ����������A E��2c�1���z�z��nVw��ߞ��|�ߝx���|�|\�+�ݿ�M�m�}oO�ޗ�Q���!0�ޘ��q�ߞ�>�v\�=���ޮ�r�{2JR��RP��f�5�kL�@]���W��n'f|_0</�B��U��w��~��1��/T�^��:��J|P�,w����{��qW3�-|�����ܘ�7�Gbkn��M��IG�� _�<�vGG��~^z<6տ��h\��8]#� ���v�藆��{i:N�K�}ڥwq�E����[�t���9�c~N�u��͓fp��,Aj*\��+�-�h�q��V����Q�;�G:�'I��������I�ݲ�S��aGj�S����b�Y�&om�lw����b��s�Ź}�5xH.����U}�'%V�d�����<]=84���l6E�J�CM��l��<	9_L�q�"��!˯x�~�g��xk���P�t5Z��9�a��lO:&�W�`:DC:��4p�Z�;��4 #��;�F�ϻت�����=�z�#��:z�K�`�f(��7���F_�Q��I�P@��Dv3��ә����U��.��+��Gh^��ĳ=��	]�zx�9;��K>�"!b�����2
��8m./�v��IL��iJ\S5s��
�g���OR$[#!A�[o��Adu>H��1"Vӣc�s�M�>�Z��Dq��9z~7���F�RRS���@"�鞓8x����>�ۙݕW�di�y���B��*Gi�7�V�����]R*�u%% b�˱zb�:c��)�@%xena�{�Bs��ܢeת���D>���)�sZ�,,�N��\��V�A�n�̄��γ�N�u8�eu9�of`�=LU�e���*��׬�{9�5+1p��ŏ	���O��C���d�՜9-�&i���쮑�ꔮ�
��2������W2�0FL]CY[-Njo����|yel��̝�l�l_Wf�i�$���3�����-v_7�+WU��uv�e�a����	�(Ԭ=��Z.Lu��r�R��`��2�N �m�����Yh[I��Mz&�au���i�wg�}�@ݚ�T�{,w��/μE���r���M���z.��3�;�1�X�7��U=Wڸ��EWY��fJy��퀪I���=}]�:�� Q��Y1�܆�gֲt4��_d�U��B�'���A�[��ʌ�)yRrOw���.�Yd��)���w�~��U�ZLQ�ȓB�.��W^��츽��"�x%���>���W�~V�N��Xl7-���������I%����>�0�|�u��P�^�u�9�̩FQ�n=zå��_ݹv��/f4��N��v�T>��C�i�']�/���BU�gݑ���o:&.\��t��F��[�]$.�Z��WYܤ��.:T�+����} �Q%*�l9��!W�ē� ����u�>�+�T2��룉zA�����'Z@i��xR���k�3g�w���tf{'�I���>5���#��s��ly�}a�@2�+����u��h�[Xhp��:x'�l!IX���g~~�'[}|�%�b��5ү�]��`�̳�����&�L�����X�f��]�y�ޫ0s��2^W<O_]���<�	��/�lǺ2�]���l�N7��w&9��:�7��PO�7����ۡ����0�ޮ�[b~���H{;���ȋB�*\�;�e#q�I��ն��)�"i��`_$��6�B��O�˴MS�h�)T���^8xn�f��+;�O-A��ɿ' k�|�bs�R���i���P���$�G�����mAvA]"��?awTpp�U�'�'w�b�%��kY��g��0�/f� �]�c�U����l�z�!u��}@K��b�T�u��LM����}}�p\��_-��~�+n���g�B�q2�7�Pok�j�p���c���\�#�5�tƄ�XࣶR7�}hxL��2������8Ջ�*"a�a�9�ܼI�\fwi2��b�:�2Kd��f@�|Շ�U&Y9Db:گo��@@vFC���C�ޗ���ee�s�X��K�b^g \��vL�:��!�<�T�s�tG�fH&j;���;]�zhŊ
�7AB�*4z�Á^�U��5	{K�D[Tyf&��魭SR-vnW�eV�b�(k�u�mqb��?w�+_	�F��X��ǕTM�V/9�-��U�g<�3�:5h	b��4
T�vgt��L�ڴ���
jR�S�L#р�]�*K��#m���څ�Y|��8�ʗV��=-�W�������r��v���Z7h�� #�a˾3zCiW�кj�X��\D�Mq[���S��������u��������_�ؕ|�vnpm���`�h���Ww�t�tܱ��*<%��뷙�u2�M�(�}@�O{��#l,�;
͙ߺ���� ��x���9�S�5�m_Jw[t��/i��j��ˎ�`�;N���ݘ�e�)�0)8/u�l�|��7�2vL9ͯE�y�#x�����%;l��ґ@���	Îb/d��E%/2�|:�ڲ��#��k�co�1u[9׆_p�>��.�
0����z#���s�/���}��r4�ի/j�q���=�T��&��q{ԡ޵s�Zu`�#��4�S/{�J8��H���=w=�`dBr�Nנ�-0�FxJ��8�^צ��H��	�Ǆ^�^����X��r�z�7(�"��[������'h�M���� ���m��2���.�W��#b���;����S��*v*=��T./fr�C���j��'��)&�
���ܸ�Ը�=�3�J���C�,4�Z9݂�mf����I��������p��)v|�f��� �*�H*��w0*�^Xx�$��Q�8�G0O�I�VV<����W2��N
S�'1�v�2�u\�vB<q�%�:�[O�RF�7�׸�=]�����S}yMFv���J��u�fײ2��ˮ?���{7�[�o�_��4�FQ8a�Yꜣ��ONXΥ^�`q�uNÁ�\�=�=|jk%.T���H�����o�Y�yS����̠d(����N�/��p
����9�T�!_!��'/�%`���?OS�N��l���[XeC�����tsŢ�'0;��GB��젼����:��o�7I�-�nz��\�(�9^�۩��.Q'MI�h*��J"6D��u�t=l.\J3��vGAg���zv<�Z{a�"�?�o�a4�ONG}]w�4����|9\��6ú�C��C5�Y�kN�XT�*!{n8\xD��#)zw�Tʍ�A���A�@��f�e#�[U��s�����iIҐ\`DӺ^��z�-*��{�71'K���>d/���Cķܲ�୾�р���t<l���+�l�c���I��:o�,�B"��! t�y�Q��q�n�������\\�=}j1ˤH���D�m��;t'H,�������"˱������_j��V��y[We� iX�v��ĨC/]	���w���E�
]n�mk��l70�����a�vZ�j�]�"�ܽ�%�js��},���Q6��Ҫ���Z��֮���I��3R��A�6v��oY��;3t��!��3�7�꯽��_sC]ܓ�r����hȴ�9)%Z
�4�8E��ꮓ5<O��iBWoA�v2��V����9�}�t��T�gh���69>�XmTţ̙<u<��ɳ�?O�����=�Bl镥/^�5�[g毲xK��Wa����I�q��̚��Pv� �MYQ[��H�,�*p�+L�".C�#!@xn3�j��`nʇ{5,r��7�g)�UZ2W[Rn�lr�GVT=��fa�s��@ݚ�MW��'���(z�����Ήr�}���%��Ig����E�Ӄv}>�u1|Q9�B���^�79a�KݍĜMgm4;mɞ�'�舛m<��+��6��^�z*m�b�i���r�K����U�.�ruga�A���ܛ\�ѱ�.�Yd��)��n���f�t8L->��ۏoW�~R��)�4I�$d��VU)����&=�~�(P��r�X)��f��v'���'}N�@G�Y𣥼DtV�����n���T��ǯXt��0M�s3�N�֑���:ɷLh�S�;��t��s����[xժ�Qc��9���Iy@r�pn^��Gi P����m�5/�ҥ����c�K��m��Z�f�w:�v'H+c�t*�G��/�:S,+vq����{j��3-	�R�]��᎔C��WE�;ݠ����:�t&�e���F��;�y��)�(j}Ycc�h�X�kw����Y��8D��v5d�������*�c؃#�F�*DM�̋��`��*t�J:��A��,���V�ث�G��Dͬ��{z�N`=��i�v�is<y�sl����f�YiV��*=���C^��o	c��=����]�%�}�uK	�-]�n�3�Z��ܭ��s؏�U�p5 to���õ��hc�a"Nv#��8�[��.t�6ɫ�s�z.v���j���NC�sYX�F�BլX5]!�>S*�2�sj鋻'�+b�M�A��]uǛĈ
�h�X��[[6�	�j.��f���lF�J
��;��us�	!�}��f��VS�E�4��yqH.3��Cȣ�7ܢ���\s޾�\�����EP�͔�UH�2�:�\��:����n�Y�-�sm*4��8��O���AZ�^������_:2�u�2Zuˊ��)`O7d�&���wJl�ŧ2n6��Յ��*5n��*�56<a�]�,۶��dZ��AR��L������	ǲ��|���/����Y3h��r�s]�8/�
��B�4̻�4�镙�+ J�/�����L(N.�2���q�"ouk �t��ݜ����ӟ���2�l%Ѭ�Cs�������Ҷ��vVbR�\��vЙ��v<]WVWp�Tj|!�Cgrۮx:��I�	*ً.B;���@��J��c���Tg{w�r��X�>��*��r�K�����6�mZ",�n�	�x�f�;�M��O7��.�$�͈��eĉ�y��((oXU����K;J3t�Q��Tu۱;,��r�6լo�Mn;���0��v3��b�A�Ƥ���5�{��� ͓�һ�
������fJx�k��^>5��A�`�V�}���ݹ8<x�Vu�,U���Q5ɵ/+�*���:�U+62�ɝ�w��G1�G��f�-�S[n����y�c
u���I��B��g���q��Y�X����M�T����%��haH)v��N|���Q�4�%u��c�r�AZ&�co����ˤ��we�kJ�r�R�Aq<��bY����z���W�p�T�)�ߛw�!#��<&]�v��T�D�W.�
�[vS[�c���W���B��̓l��W�;�T��:���Z�z�1$��ROӡbK^�^	mG�f]W*�;���Z���Qw�Օ�-��É��J�20b�:�e��mb��Hcv�޾�-�]���R9g{�Ŕ@tĈ�̆t�wNfm�iruީ�6Vuw�\N�Ď�Na��[���
�B�ۘ��6"��d��αPd�F�̨�̚N�lF�,�'9Qd�殖A#i9s9�q�&��)�t��i)�\ф�W(�&�	4i��؄�*�0����b1V �.F��)H�F,&#PX�jH��F�]�	W5�a�&���svcF��vᙨ���� fk&�6gw8�����cfS��,��b7.�J61	03(�]یb�81$�9�fj(�qe;��-&������\�FƓ0�,�v�c �ȢѤ��X���(
"�sZ�ƨ�l{^�ǒf)Ճ^������S�'!}u�P�5qk|n�����'�h�Br�6��w��GZ�o� �=��jo�XݳCJ�}���l����hU�ĝep�$%U�evGK�ޚ��.��ֽk�kb��LZ��Df�l1��I�>��a�A��*T�Q��
'�*�l9���KTcT}<ys��w����?1�y԰%�]���tq6�A��R��2zkH��}���}����Y����vA����FOq{�`g�׫���9�������E��B�%q+7���\f�D�d�j"pv�_�" �7��@OK㱻��Lߴ�#+���	��4�|�h�g^���t�՞~���IY��U�(k��yW���jf��+;�C�9�!���qJ--s{έ�{5:����$�2tY�tdT���c)S�X�W~Q��e'N܍���Le�=��6f��5�����p�v,�:	�g�!�uי�j��mbS�������FC�������'P��	���x�
�ѡN�n��|Fb���A���1sթ�Q����"�9�wiS� ��3mך7�����/b��*"i�0ק��ɡ������pW���uȇ��� j\j񭉉��c���j+F��t����7v��l��Y��/V�
�ËY�Z��r�.j$S�bf�耣w��|ܱ�3b�F��Iop#���L�6��[�+x
�סM؞�P��oeu2�'�������{
d͟��B���$�'�2�T��Q.��v�j��oL�r$,t��gt��J�jU]�f�\-��׍�_8jplˈW�4
�2��:l��<]:�'�J)���
����������ȃ<.��<$��w������Dh�����2kc�U�w�z,U��)�)�CX�AvT�bȈ>>L�ɽe�پ�VH���]����>O�39�-^� �$(��Qm���bntlQ:tq'���u:/9Z��T�(���U�+��d<?gǺ���!�Y+���2�������N�� =�dM'~���G\nn�s�/���#�w��7���J�q�l�;Kd�ζ��_�o.�%���GGT���b��J0���<��Ze2�b#xױutvzS�Ȉ�)\���{ˌ����EM���\����y#�A��b!U#����L!�Ei�7����C)f]���L��k�Y� �ྭZ�{W�%[�٦�"�]����|=U>#NA�^x��030��0�Y��i��m�/�!�.P9:f:�yGN1��u�:�V-\���s�_����l�2�G�n�4�(̾�}��m�lк��c�`b�M�`L�.��(��V.�JnH���7o�����޸���|h+������U�z�#�xxx �u��I¸����?W.�J�#(RX��PEh�r�C�Ϗ���P"d^t�k�P��Z}r����[C`=Om�y�WF�
JPW�vU��+?	�e� ��w��C�딓C��S�Xa��Y\ĺ�tè`�y� �{�Z��_rBa噱 
.����C�wƍп|Kc�Ը����;�3�N��d="�{<9�C�<;�}<������v@ЬT,Y#+�t9���u9G�"x�r��\g�zS*�Kui)\�Bk;�f����R�3�>��mɊ
��]��Wd�U��i��P�����pי�y=�zoef��W�����1����鳹�J�xeWZ��-�2'�(��_�����Ӿ���7��-B���،Ƌ��_��LU�M�o�Ӂ��C��9^��u1��$�#�9�200
�嬙�=0�Zϋ"��G"�Į����Ӟ���l�'ݾ��Ů᪰@�5�M��D�����.�)�M9�";�+�d8�)H�j5�S�Ü�;# te�c���l>f/�y���Y�oTY�}�����V��ݶ¾ݼ�N�<��qϦ�Ц�I�C6�; ��,�[��-s���~�R
��]i���j$ߵ���h�m"��i�2�I��͞Uxo&��"�7�ϭsX٧gP���{�:�7
u2vx���A��$����fn6R>����M׍ [՞���+��MK/ڹ�o�Q��CM>��r$�xDGw���I��=�냺���-�#�R{�E�"��r�{��o��S��^:���}(�FG��,&�R�=f=U�٢�zǝs�I�P�x�:��6�lئڵ��$8��%X�Q9
1� ��h�;$�Wy���u7��{�;���q�5O�{X��z�����+�� �q�<�WI�(�2��K��k5W׭���8���ȫ�H�v���\y=�7�&�<ɒ��1t�ba{3n$����r�N�D�a��k1�mm����'��U�uU�I:�#�$T���ӛ\��1Ġ.��>��fV�U���X�^�a����\=�<4$S��oWMǨ�����:*qXa%P�Z�ѽ�qQC�T�(��|�A�!X�MTd�en�BҮ���Y`��(���:��f/ݟH�u1w�N����U�>�e����G_}`�%x��,��TZ��7p	�]v��r޼��LF�WWL��%�5���[��ue��iE��vL��Uu�*NZ(S�z�kl%�*F��%�S-������F=
�������QSy��Uw�{�����`ks�3�#y̭'�B M�r�u�$L������
��XLV�:g���mUp0(�<�.��f�;#������7�p���Y5�S/����X/�&}�/gw�m��G�y�S�r<t�ċ��4���%���~J��abu�cK��q�6r�A��	�	DCFo���n�Q��V_�����8�P>��7���m�\eS�L}����c\�����{�E�ͺh��ʽ9Qˮ�h�H��t�uL��${�n��M�t��zn�ֳ��1S�&�����4C�l�8�6zzG
'����*�#��E+tT���V{'# ��2}�|����l0]���ƒ��Q���N�#�� q�37{��'9��'���'�@����Vc�QY�$G�׻�{���3p-�VAm��ps�	���ݯ)lx���ӊ����>��q�M a3�(OJ㱻)���$es�to���4�z䋙w��e徔��Q3֧�A��U�A��\��'�R��i����g�d��Z`�P�D�bXz�ޠ��)g+�5�܋Vw-�c`�Pe�Z;]�<�;���;lp��[B��l@��k�r6����n��N5�O5�&�i�kh��r�)'�&��:wɅ�	�ug�L�,9�5�]�⡼/ε9��a�W| ���{�}<U��3�d���U�h[�^��zx�uB���CMv��-�����,]�SW�v�+v�.G�zs�
��H��H��]>TF+��Q:��j�`Y���p��V�ھh�66'�YPo g.�FVK��T�X���.*dLH�u0((��㙷�ù���r3��'E-�.Z�c+B~�3b�F@ȼ�l�����x�y��F���?z�V��,:��7j�=��Ȇ�Ҟ7]�0hg�V<�,8��'��%U7���UI�L��sCj�݊&/;������f��!��r6nR_���ۉy�_1�W�x��ׅ=��>�ف�N W��xPi����T�����u�^�Ep��XxFP���c�]a󃽓S��s�ﶖv7�/o�ݣ��[r���{���O����Yt~�up���ԍ%�K�c8�d;ٙ�����n�n�0>�
1�Y�ߞ����O�$�3�򠠵ż�C�2�m��J�.�͊/O�����a����-/zd^�s�Y;\��o�L����^�Q{n�1���Tk��~ŵ.ۊ�=�x�OJO�4h��/Or�����}ާG�=�O����R��n�\ L�Q��ݘx_@ `��,,Z��5<�/o��k8�Z�[ݺ�ھ3)V�Di�6��s���Sox�b�z��;�Y�����=�9���Qe���D̘ȏ�#�W��ʼUq�r�V&�\wd8�<ܘV�"�����A{5���ꍭ+֐"�`Ɩ\��JU衦S*x"7�{WG�"+qG�+���������M�5��Y�t�y�${�G�$�騿u�72��/��E2�PK6_s�w��мR���Yg ŢU�_�˕)Z��a*�O��4���]8�MTΣ_ ��x��V�7�Ȯ��r8X���ҦK�e�s�(�Ȅ�8�v����yBv\���5c&k�U3��SefT!���K���@
�WZc��*�^'`�}�n�ޡ���co�[5��H:���w��+�~����QT曏my���x
�]��lb]U33��(�r�2|�Mӌ�WR�x����ۿZ�H�ӮeowijJ5|V�:�-��7�f��k&��j��Պ���t��g��Z|Mޮ�n5�Ģf!B)@��vcw5�U�)��tn��LpO{6ӕ5�[K�q�®տ����{ON'd.@x���1F7�|�Z����y�ô�5��:���:圱�t����0m+^/K���X���L�z_q�ݸhηX��0ߌ׶;nV��c��S���4Nv9[g$�t�W>�8�r�<�?��zgs���LIR��ɮ��g-N��Hm	�x�nLq�� � �[�l�L�����#1�;N��l�
U�Ҭ�o�r�M��%� Ϯ"6A�^��;S���HO�ɪ��iWc��ǒ��HF������3�h��.o.�x�DEiY/�<Q�����P�!�m*���]=;p��"�q�9[v.����r�m��{�QBMA`����.��u�"J"�l�MJ�flz��[\�#����Ϥ��$��[s)�g�P<Tl���Σ7�����Uc9�n�h�z2�1�ł�e�弅�;�9'z�i�ү%ǲ�r$�lp07Y�!#]��'}����EB)�������TxW.Ķ�.s��:����'�{�oo]��~�g��D#<bI'�u[=E�B\k%��/>��#%+]��^n����V���D���Knr!ۡ(#�A�G��["�p�hO<�����Ցf���~�3�ʼ�kF�_��RRS��'�q�?uWI�8m^i@����Q��uO�l������WR;Gx�:�כj�ţ̙<u�s.�jƸ��!�]�O��I��ړ�@U.��]��]�K�Z��G!h,�ݹ��N��%G7��)Ä�<�&��������K��c�\�E	�_`�v�ky�\��XXwu���݋<��.�g���]�	u��.���@��޺���s7�gs�jb���<=�z_pM�=R��ϰ�$�U�S�k�1�#�~�	Ŷ��d-45^XXwh�\k�1ud=v­v�,稗���;a;�7�/L��Dp�`�
�GR�$o�eG���&+�izs>��\�~�M�?{m�ϣnj&;�T��D�h3�>��B�WQ��0�4e����& =�����8�e�Fp7\ȾsQ�w���WL�?P�� Z/�i}ST���Y�WY�%��L�d�&D_$�c��Cd۟b�iN���;��ݖ���;���E�`m�	T�l�89U���Y,�hr�����:��3y�=7�-{'���DH�5'��$�('dV�9�}j�H�N���]86�ea��=l��1ޕ�W+��"`����X�0Q���q�W ������dK��Yb�4�עʐ��ob=:\
IRtZ�S�%��~�B4N�I�x��$!�]�u���[n��7�x=�K0N:׎&/���E��SD`}'Î�gU*
�\�hG��B�ȝ�}1ٓ�n/�6;x�^,A>�e�1��SV��0vm���xY[\(��p���K����c�����B��`)�s�F�kz��*H/�>2Fp8�m��㽬y�[J�����8�T��]+K��q�|!�z���B��]�\/�?xx 8���.�.�'�A���:�F'�'�-��R��y���^�c7ΩD��*\g9�����a�;�i��E���C�tx��PF��b�8��ƽC��≱	�9^�W�L����xCݾs�У�9�#�p� ���l�;�ҙ�i�FW���6��I���O?X���v�����s�ix�9$8PӀ̎c���&��F��ZoڝL7����)(��=�x��6��{���2l7 k�hel�2MqD����AvEzWPȼ�OMZcud�U�r�vWZh�E
P������c�3_%(it�=C]������2B�;��0o'S4'c�M����7�	�b럪C���Վ/ÝS�`bu�g������k����J�6{�{ۮ?qS}Y:Nv:��"Ԑ��ѿT��3�3{���A��f߷�p3�h3��lO�s!c���2�DS?���M��a��Y�ҝ��SKY(�2�5a�UI�N
#�&n���9��>�����^���������ȗt�q/3��=��/��
5U��w�,JFE^������[�=���p��h5g�d�l�y	�Z�'��w=�9HV���%ա|�9��/����[�P���)�՜u�]]6[RӾ�.�}�U�U$��x76��w������b����#Skgn䇩��1���6��lms'�Hq)�bO�
����Y���EDM�"��5�S�ە�qӝ2.�Un]�\�a���l���a��yc�������4��جm��g�n��;5Z<�qg�����:�.���Lt�[�'�i�j6e�y�҃��]}cj1���r�Q}J-Y�E��FJw1���i!|�윰�DԋW4�B����UygRP�gf;g��a�(��K�<܇�f�ҺJ�f�jt�:Ew+������O[]V��e���jAL�\�^�YO�\�δ[}z���`�.ws,�u��tM����]����،�/�������"k'�4�D!/L�-��L8a�8�on� (aa]�q��*���9���t�*Z.(�L��Gf�᠃ǫ%jU�Y����=)M���Q��vxs�l����z29X�R��z���f46��[�:޵x�W-tL&��liX\�lAڳ$�#�>��ײ>�ocb����Æ�dV�� �'�Ⱦ|_�+�s9;�{�.��&]�+���1f*��]w>����_-R5�Xp�]a��Ѻ�7mc��m����>O{�t��	T7�əu�y��)ӝ�wb�]����_f��M=�R�{M�}dz&o7�~����k�c�bq.��HoW4�6X�u_,�������]��E79<Q���)���v=���Hs	�&gZN�b�Ռ����M@T5g�W��гG���o��;�\�"��a2m#S\}N����w��+ȲT�/0qWk���7�YQ�奬;�(m$�/�M��۵nL�t��μ�N� ���B0V�⽝D�1x,�$#Gr����t<:^��Oc��b�ӽө%M��vR��5��.���@R��N^���7Z�U���֚�-oRx2���r�c��k��gM���}�`s�>W���ѝA�z�Z/�A�������Y{n��e_f���vK�+f��X{ȕt��w5��ကk�e�r��n��!$C�S�+�)�'�4r�{��T_lQrM}��29+�[�d�u:P��[���N�bs�<�P���v�`�Lv�0[�>ŅA����ƿc�'<���.dJHo9R�/e�k��Dn�CV��q�,���J�1���<s*`��>��FG�AN�����NF�y���f)j	dPݍ���}�v5j����4��.�w/)��v���d�->9zn��t��l�Io��-ԯX����.\��n6RM)8��!}S�UK��w+�v�q3�1�P�à�8t3,&����=t8Q�KW_r�F�v%ڲ;��Ugtt�!�ӈn洲���C/�Ъ�@Q�$�3,F7wF�j.㴖�]�T0���PT��	D�)�D(�L��ADm�4����؃i9nI�wk��2ARM�q�nɄ��F��be]��!��usF2&Ҙ�4�4/nFM&�t�Fйu�͊0A`ш���H�s���%�S0Q�1r�9��$ت"$$�4b��+�QCL Ed'u���X�"(�E��Й�M)�sb���0d�ذh��A%��"�#!���RbJ43fh�hB�#S�׎���n�0]E;�>���]C�է�}}��++�Σ��j��G0GphH��q��Lu�Ͼ��ﾥŵú%�4z0l+{}�*ܗI�+,�l�\+��������O���4�mb^љ�=�9b�^<��W��a�l�S��������"�>L���Oeۓr��׭\�_�t������G��ϋw��ąa�Z��y	�w�K�	{[�'��>�����አ��2���y��bY�z}	K��9�F�h��oz�6�W�l�%گR�}& �l, }O.�m`��8�!"�\o�&�M���ː�盓z�$NDr�`�V>��CE��X���"��u�2.��xWx��#x�����)�dܫ�V��K�&�q�æ���2y7Br�S3�JS`��P��'�ME�֨8�ˇ�9kjVM�x�՛b��*+ЀK���N'�x��s�I��q��}>l�G�r�DgÖ{��W���5�E0���S��>��2^3.#�
02"Bt	Q;B��Mr�}сu�Ge�����Q7�
S�]l�V�����cj����
���xvU����5dB<#�_���4��;5����.1�Mo���ˏ����R�Q����cvE�t�i�vk�Xڹ�K�
��G�C���;HN�N��Ÿ��;���9���^wa;�Cх^5ݛթ�])����L��.u�_�w/k 
�{TC�&`i�����w?��-��Q4�e?z�1����a�[+�G|��[��:�'w��QT曏mZ���,Z͊��a]a��0m�=������b��[7�)3�g��]�^b�P�J����_h:��'9aƝ�*��ME��CJ$ex�}9
�r��&�gR���y;���)<f\���v�$�c�oҔ�:�75�9�pǕ:T��B��W��uN'g6�=d���V�rJ0$4GDM�|��+N�.�;��^�6�v*���>���B��(7
V�ib{ry{dU �\`�5&�Z���T{���b��M�S�P�]8����b�p�Sx6�TbT��3Zh�	6�=^�;!��wؕ�X8�zpi��"��w���6<��٧�!l]Mz�pq��!�u�c|k��|�x��a<�o�s�e�U3�F��ZW���1�FD�ܸ�pM��l; <Ou���}amV3-ύː�22�'��o��K�2�F��ZGZ��_�\{)�P�Q�p1��Ł$-&4�jsh:؇��w@�.[��E�;�֗GEp�lf�=��9�\7`h�Һ-_�����2WLJ]�v�	�7%�Վ|�"9���j�����5��YoN����2���u˳3:�GN���}�X[i*�w:`����c�3xu�6�gԫ��\�f\�)����=�䳖���S೩��	m_���eF�u�M��؝ ���G�!,:H��1�l��qU�Lb���2?3C�27�V��D��ۜ�a�4,��Uk{u�B̙P{2ys����rbgz�떏Vr�8��~	Pri�]���Ȳ��>����^�����=K<�b����ȫ��ѽ�\o�����BC��Ģ�d��K=�ޫ���z�vH'�5	+Ux�f�
9�[g�3�,W!k�]n��쬘�^�n��(�"S�M[�l7{f���7�E̳���R�����`Q��sx�^�c\Qȴf.6��5:�B�u���aﭫ2��9���ʨ�]�J�M���V��..������\t�v�"��������7\ȿs��Ӹ}��	��q]�V�P�1��BQ]�+�������4�x��DpT��Z]{�g˞�v˨C��˶ә��9��m#^��N���Yec�[��͊���̸W�Yd׹Je�:�V�]�V5� �
F�R��z��O_S|rm��cuk�ۮU질����3Y�����h�uՃk���fJsh�u{Q�tGZ����X]�"�d�N�-�zAt}}�f�t{E:2�x=����v��V���+�� T��qNQ;��"�Fv����{�R��p���I	��X�1DlI��J����KG��*�SE�>�4�pBS�"N�V�e�����nE�Q�/�R+)��@�9�`4)I��eDH��(�mW]3��*Q�k�KŜf�zF<O5�D��+ty�Xt�1Ȅv�j��6����OQ�#�́UK%��:Dv]S���8�����t{ס	H��i��D���V���Wa�����}�7�����5��{��>�%�]���ƒ�9�1כ���~��Z}��f�vB�2�%��$p�j��OiY�$G��v�}Z�$q���9��1.mL�x�[W�g�6\e�u ����*d��$�9�0�L��q�͎����FP��轄���*�eR��#`l1�7����?�NIƆR��j��\��
�v�gٳ�t�b�\ifmq���u�Mȴ��I	�FOy9Z��/E{�'�F϶�[�6��R���84��m���p.�4�:��w��UC`r#�j!)@Q��X��@�^']U�O��a/32�k�:F[��=]����
 Д[n���P
�z�o�z�X֭�Nܺ���	YH'u� ��ɞO8'���z�̧�>�o\�N���֧Je�9�a�Ǚ��\��f��
�u���ES
��]���qZƳA�����u�u֊��Vj��<< ��o��$�L-��Oa���wi��Aj�B.=ʂ3�
�>�3�!I㗽���c��=�%�d��;�-��+V���J�^���[0���e����;�v����*b�1�������=��Q
P>1POY�.|:�*��=�(�ِ&���L�V��p�/l3w��R�ޢP����q������CV7��.��n�_k����cܮ�f\B�V-=��]5����� >�h�2峫�=6��8������2���g�}����,[9�z{PX��~E���4��El:P-�l�N���!ụP"i�d�QY���)MB}��
��͇캭�"���w`������^x/����`��p���`�G!Q0��iԽu�����C0��]��]�ĳt^�P)SÞ�9�Fߞх����a�2X"
s�-? ���h��z���k�\D�PBE^*��8)5blL��0�q�gv�f�u������8E/Vo�+����+h;/2�^����J�S�t�l�n��Z�k�Yk�+Y�_�f>��>g�únB�r�m��f_d��|%�ǖ�ͫ�&�.�}�2宷�euL�9ۙ���mgV����h�OcTʠ�V#.C���g q��(qz��ҙ"� qw:��o5M��U�}�V/f�}m�\,�qx����"�6�M�T��H�)�k�c	��'�9׆{�~?Cv���gnv���/ƭz���^��
0����Z%Xf�$*T'�'v&G;��!���Yd�-�}��BQ�]l��S�tb됅���K��+��T��:"��x��E������pe��u����t��m^�S�qͧ�Y����^��1�P���9&nfGs���>�|q�꿛,7�[�^w��%#cp��9;�9��C�1�k2/u��۝Z��=Y��z�D٪���P�
Ќ\6P��:Q�\����7���Q��w@ߪ#Xtj���u�K�I1��9݂��Y���iD��9���'$�x�nf�Y��F�c[�4j#�z�B�T�q���\o`��"�<��a�(�@|Ts�Ιp��V0���Z1X��ekh/�@M�^�#�����g8R�f�gcFnT�e�W{WV1��!춗AS~�`���F��ۨ�����d6LR<������]8܀����%|���y��9�f3����h�LwX��1G�n��y��R̾�x8c�"�'�C�����S�͗�B���}���H���u=kf����b��Ί�c�s���Sޚ����=��Rt[E�0V�꾺Y��H����8�usFr�_�������{}�1_z�(Ԗ�>�;!�CHPQ�J�,�����i�h6E剹�ʕ�ep����ݖ:�����l;�d������2�$C�
�]R!�
R!��6j&��[��I��rR*���u�k$z��є�ep��=(�����!�|T�bH�ͳ����3-��+���=	��5'J�d��PrQRQ�#���$-&�ȓ��V�8��a��3;;���t�
�tl`����!�ʍ�븛��bt�K>�D)��!���_M5��u��󠧑ܚ_7��*��ri8}qEy�����
ct�OJa^��Sj�?A�:!k�K�o��׵���9M�4���
����4�%�!�2e�l�*� �ɡ7�j���x�?sI/��lF���9���V���Ο-��/*u̳�oǶ�$?l���o����['V5=�8�9��Wu[�{*��7Z�����E�̸�zk���gg_B�
���S
9erU�[�z�-�y�<1��4k���ʑ�fY�H.9���Q�t�SOUi�X�^Y�K�k�ϫz�@r�9�5�w0��+��>Ju�R�oWY����\5�}DS�]4�nn�:[愤1\o%h:�N5�\�ri�lR�o�}��_Z>���<�٫����&�2���u^˙��b����˗<�k:e:F2���K���r[�je�8���6���-ټrcw:��R^���	��az���$$�xP�I�T���m���T��n��o�'�%��ݟ."n�Ŵ<r���'e��XU����7���]�Z�i�{��\4��}�H��!o�뷕B9���e��@��+�cv8�Q=[J�s���wcm�����=T�6J��ұ�^�`6��B�����<��lN:-��5��������EGO8��Դ��=�X.o�
�)F֗��mB[�@����]�>��8�)HL+�֟@6�-��W>��=Aв���&�,����-�\;}���b���ܰr�wX����"�E�Ң����v`p?콷�ˬȺ���|����;����/#
�D��Wl��IĪG�9�MΩOku����JE����[�-�Ӗ����\X��s;�v/��- ���M|��������t�0���f<<i�n��֗b��.��SL����5�/:����X�4Ro��p��<3#�td��߼  $�'M>7�D�<ՑJў#���=� �q;ۙ��z����q�e�5�u�Z&zG/�3n��B�L��z:�k��]���bM�*x������Ǜ�i85����\c�:ګ<�گ�Iu�.^N�n��C�Z��S{7��T�ԝMZa،�ʭvbF�����Ũb�*����v��fZ���׷+2��0�Z��`.��란25.7�,���Y����Bm�J��9:��s��^�޹�0�|�d�f���9؞�����������v>�h�z'����	ϝ�+-����v7r��ܥ��v���mf�������]��P9��J���ٵ!B#����m�N��f�08�E6��[zs�|f����m9V`�D����U���K3�X����t�an([e��ʥ���1V�:�|ϙ��=I����M�o+I�������_��'���ۤ[�ӯp�e+��a>�N�3��Ά�qh!��F�d����a��6��<T��2�"�Â�wwB�j��Ǔ*��{ȍG7^�q���2�y�#OL�V&Ӿ�]���)Qw�����d�O�<Q��A��.Qv:�R�c�y`ce�����{`���s����7�k������������t��WEׄ��w�>�����E�@�]��q��8m8�}��P0������@J|h�ݷkK��&��J��;I�Q�mŲ���wapAKb���b;��B1W�=��f6��X�Tξa֤�0�8�*!h+��ly����	8)�
�;REgNz���D���U'�k�5p�C�3j�pJ�d(�z39�����P1�kC��E�JhM�ڿo7���M��`2ƻG�����9�gG�ʗ�ҲTھ�!'r
��q-�՝��mL�����+���9ٷ��w�_0Iǝf$'>�n�ŞKj�s�Rsku;�*W��(Б^>�=���
�o�6���i��Y�iv�����ξ"��[f��r:��z�%�6��2rصn��Q�TiT�Z1��v-w�T���l���\75�t6�5j-�f�x,8v�����J�����q��x���y.�vԱ[T�Kkz��Et����x�=��T������w9 ���Z�u`����v��Y��&�r�vD=��ڡ���}�-��q���c�o��X��8~]�4S�D��s&"IsR�:�.h�����jnWK]���;�Te*h�=+�U1���B���8�Z�b�=M��!�%���,���������Ij)���nu�_8w��,�(G����BT�� �!\�W���]���٦�G�)�]Ah�Cz �O��dt�Դ��p�����uEx`ٯ�hb���\�gI���N<����/����m��o��U3cLv^�����=����0knl81|:k��̶�yS�sT`��1Ӣ���/tS��P�6��	;w��t�{�����wgnP��2.xod˧ۊk�`<��4�]N\� �՘��n]g*�MДdO�W̍������8��+�95j>=X(�w�)0��!�z�8qh,rq�%�[g�v]0x8P�:�!Jp�J�[�X*��/�6�����;_#Ĳ������"�ڂ�h�7.Qp�����i���'DZ�s���n�V�J.��׵-<=F��ǶGw�{˳e��y���&s'��T��K_n*�3�2�|VLZ�y2�Y�?q�ф�>7��y�U��M+�T�����D3��T��B�LWv�}�,k8"�)�W`;3W��&�P���W��ږ!�F�YQ�j�,����ŹVX/3;�����Q���]@ξ����b��5�/빒����vT�G��|�4	�0�;�Y�@-S_S�ܬ;A�
��%W�n�؊���Zjl�z���D�oKt�R�4kv���Wk�.TS�y����+�V͹��xfR��5�ݷI2�NJr��4�v�ʍ]�*��J�K�-���1��u ��{\�vY�+�t�M���k�h��/j�Y9��it��@�n=�귅^T�M�����ǡ�x�r�EX�osGf��y��E�i�W���+I?q��jY���e�b(�=�*ũ���������%���1ض�9(�7P�{��]�ra���[��ʐ����Z��mF�粲T��Q�,��G�;������}�i4ZMhe�X� �����*i�gGMޜ�uN�)�� ����t^낝�P���3�(���Ϸ6��myvEC.����\���{\VC�Pwk��MQ�D����ʾ��+�4�%VQ�X�SQͭ��-ܧ,���{A���ǇY��ec�0 ��30m�,ݜ�y��[�.kR��FZ&w0Մ�I)���ѵi���^l�䝍P[7}�ZPj��&�V��kB���)ˮ�!�����g�n���1Del�h���'01#��C�!F�Q�ٖ'�����?���u�K`1� Q�fd�b(�d��F�F"��wj�K�Ȭ���A� ��kwu&����Gwۜ5��"�1"b�[�#I��Ŋ 9�2m˚I%�4�&$�#EF�.T͌c"��9b��Df!As��������pL�p��r)(Le�9�0n\(��nRI�wsF
4F�p؍7u�0X�:nIa���A#b�#Qs��t�gu�K��cF�&c%��MwnN밹�)4Њd�������TXd ����(��&j#0�,뱓E�\��¹���~{\�S��Ժ\ ��.�s��7��=ǽ�����8��	So`��4�'�R��߳4tGջ}�(�lz��P�����;싛�N����k���̃��-�K���8#���5��O?�S5p��!#-�2���u��6�6m���fW��6�su��f���Z�9X�����ċ��ڤ�X�һ3RxYGhY9o�C���X!�C�Ⱥb��z��Tj2�;�)�	ܖz�\_=���"��{G�A�]=N�b_��ꭈ�n�T'e���W�*[�cg���U�#��r�Gv��C2�u?J���oz�>��
��VԤ�ԪnLR�t���i�0��-4��J�~w�W�[fүEGO�Ϥ����j��5j5����Qx��Ͱ'4}�[Z��Ϋn2��QP���>.3*�I��b r�K�EO�
����ͯrܸ)w\yف=ؠ�,�F����H���`D�PM4�	�1��MN�Z��b�˻�%�!\1%�cOiF#y<G��"����C3��PHI�ϖy����΍#E�u��Xfy]��^��S	W��»����ʹ⮈ܽ���ж�)IMX|�q7�2k�v�Sꃅ��)���&���By��W�yĎs�X.��<H��T�,sE�k�#x�����2���u� |�Թ�S����,��l^����67�֍��_�}c:���6�s�5�>��Xq�?@�� ju����ۆ��Xg��s����#B\:��/]�]�ݤ���~]��c]�YUU��-᪄�t=9��۳}�h�ޓ4����I��w��LU�{Y�ۮ�ba�j�?��O���M����N��l�i�f�\�ᗙ��=^W�V����ؘ�W�}u|.���m'[�C��Km�@�����"{#,g!���z�7=����4��Е1�9t������_�fFe ]��&�*Jqׅ	�I�)�R�mH*��l_5��y�+of%S�b��9B�,�r �W�]��A�XU�޵�=	|�^�5Z�g-j�l�=?yB�%[�o�}V<=��b��#35���q�ȃYl2�P��m�=�p��7z���;4s��c����e��辦�R��K/:%�8��e�.��M�������=.Za��K�)���0��],�`��f�Y�K�<{�s��W5�kv�,�9K���A�CUGgZK�ө
�l�o.:�394��� W)�����Ur�� +�h��\�t��˲�S�CS{�5|�v%��muD
:�����g�0W��^V�1�������[%��O/�5���^P.�;���آ U֌�\��:��c|�|w��^�k��O�����Ѫ����%|�t�Q�������2p�1��JD8 �*5s�G:�1q��ұӛ����WC�
O=HWol㼓��q܊	��(��R�� ��yvf�'�(�p�^q�[�r��Re�}-���͸v�*�29F�t#�AZ�oF`�m:cl-�����v׵2�7�5擃I��E����E��8;*��/|����^�F��<o��ڸ�s��L"��\�v`tZ�;����0���=�Q4�T#S���^eO-}��kە�����g�Ƥs%��x��ǺF�צVEE��fӋȾu��T&�P���Jw�淽�yp �@h��R�du�]������G����Ύ`߅q[��Sn���+g@�:�j\�V�a<�g�h
�E���:Ro1�9�]w��;���=;b���CX�Sr�ݡjwbܱͭS�|���\qʗ�]��+���Žןb��b����o{���=�*�:c>�y=�7�.�sC��Q[����g�����v^�}��*�s-(/�٬vm�9��2���6�k�q7ʕ"󞜺ۜ�;R�6.�pO�[�I�B[{~�ٶ���9B�>�` ť&r�`~����~�8��YjƗK!��l5��}b_>�{=�{�ȕ��sۭ?v�7y�g���]�R��qo/k,=�����jjtIO�e,��Ȩ�qQ��)�|�Ӳ��+��[�^-<��5�"��������Ի���1����)J�Tt��H(I�iIb���뫼r.]�/L��DT�8����q�V�e9F|�)���q	l^��)��f4&���]z���N>��M?vs�m �;��<Ƞ�9NY�#��%!�:(�����̇	��.lZٹ�X�-���ysA���6�[9K�Zx����L�����V(Ros�Z������)�썲�����%qW�Nɇ/��j;+��(���1I���w�7R�tv�Rw����Ӵ�PF\�b��q�K�͗/�r�ݗ��u��Wu�R2����Vv�z��㚶qc0_ _CӪ�G$�;��9��V7��h��}S^i8g���~��6��6fg�7������R�0{B�{w����n����mT�a�����e�rz_r�Sbq�����2�=�Fmg�߱s�Rs�kT�fZ6���Ozչ�ztT�a$��5׽o}���Bv�w��=n��U�u,�w�;�^v����pt�}�R9>�f�E�|.���
���ѩ��V�!�p�t��-�b@�\�)��`�u�������u�8T���,�s�'�s�36�n�M�P�c��>�\ͪMÖ�|[�=,���0d���:w@��oÌ��Buѭ��it�q^���m�T�P�7��L�s�y[����|
�2�ȍ�9yP��k�HIJ�-c�l>�҈5�yU�ČV�%�%����1ܢ3|P0�W�Ԥ�L9�ʖ�I�}r�{�$!+�N1J�k�*-9A#*���8��ʃ�:��z��Y�wp�<�AI9��[��걛�3�.�F�Q���~�P�&K�g���b���lh�sq}vk٨�8\�GcUku֫Ve�1]/��r܈�wI񳖇WV��֘;�+�t��X[ֶ��5��מrؤ��Q��}P��OWY�B:�duE�*�%з
39mmc)���e�5�s��[q��B*��u@��;���|�dnn�9�
 �C�<�`��C�[J�;ո݊�rǗ`2�?iWh�p`*x�Q�}����|y�Н\�ŋ�h�ҿC}�(C�|*�g�L.�֧څ8��q�����ʣ`��ryvV���h�y.s�f^y�pN�uj�=N��l�n���	T�U�1P=���;-Z��y�e�2�|�)l��*sm���eTl��Tз�lc�_��:�u��&�?xNg"x�V>Qn'3)������0�>��٬�"-vJ;*3Aۓ���drELe&%�P��7u��X�s�ؘ��k���že�o��"������id�����M�d^�$e�h�����Ojjeu{�v�YQ�[��ܓל}N���PFN3�;G�ǲwv^�b�5Pv�a�g묎�9���W�qs��.�[vo^zy5O���O0�W��4g4��N��7��LV�eL�uu���J�2���o�Ǚ�]���]��
���+�:Ԏ��
4I]]�R(ν�f���7IFe��P���)�XP�|�*S����]��A�gQ�#�S�p�O(휕�Aޡ:�׶�j�����t������K��Y����}�CY虯)�B�޻w=V����4��E����ضd�8ֺv4��a���|Z{��EFD�뷟�t���R�$�|y��ₜ��7)���ҕM�kc�Y���͵B*;q�u8�-�c*���rbhb7xЍM_��t=-醝��\�/鼕�k��J����!Tz�Q���!-���f[Չ���އo�3#�@-�[����'a�8�Y�aOy)���O��ম���Â!G���pM{�V�=ύ�,gr+����8�.,��tK$�6�O���9�+�oIi����[	�n���4G>�u��Q��{0m�Tk��S�u��A���a[���H���:�����[oNC/���x�^��ٺ�����^f�,�\y�Ao_���+ �_r�vQK2���f���`���CZ�b޷�uk�U\j2�{P��M�|��w�r�`Y�;+:��ܴ�
�KI#�}{G���L��}SM'�lk�pN�1#�5��Pm�-j�V��p�	+g�ln��U��u5i�kͱ��eR�V�%Y��g��{���e�}e����+'?E'����{=z��s�;�=yx^���ݼ��~ۖ�Ռ���_:��Bm�	+#/9=�L]�`�#^w#���8��%�X�Q�>��;�n��e�c���B~�3Ҽ�9Hc;ގ�������z�g�O{�eC�������A�8�����msX�'6�O�X[��no8J��gM휯R�ϒ�pm�wEd7<��*oXwk���a���X��P�������7���I�go� ��;c~q�g��;��t�i}TV�T�-�a���ċ�̜���w3'��3i�AN�6`�����t]-���=���G����#k����Ad���̷�]Z׺Oi|���Ӛ E�n���\RWEt��R��i�:����F�/v��l�c��A|�J����n��:�f b�*��)CخfK�^]��.2`(A����EY�]�tLɈw��?�����ˣ<��=�-�W�j�{�P�ߖ��#�
�w\{�7�Z1gz@b]�gw�s�r�8��O���v�eyq\G/����G�pZ����k���������>�ұ�,�"�H���<Gm	�Yܶ�Vފ�|������fv�o8"�|v�>jᾇc�p��t��1�p���jR�垄�t�6��VV��M�ڿo'CZ-���N��5���#&�DȂz�;4>�.`�����X���sH�b�z[�>����r�����s��<\#��a֏8����n����3�<�ћ�g�߱s�Rs}Ѻ��㱛n�S��닞�:�l3Nbߚʡ����f*���Y�o�:�K\nr��j�-I��N���i�k7�sQY<A�֕��g�;��RŒ�>�g��ɷ.z��y�H�i�S)��z��
t�Ϗ�NO;|��Y-������Vk��yLx�m.�n�\6��C�Pp6���a̧p�J�a
�gL�E�ݽ|gD�0p��ݎ6�w9`�5e0�f��SA�T��S�,�r���G��mq��e_D��X��J(�z���Q)���q�:�{��ھ���6s"P}~���ڤ�_�7�+�zV���Ĩޫ�ƛ�kc"�(u��� s��<˪���*����=Έ���-y���jC�:t?P/>�g(S��<�*��k�HC���؍Sܐ�N�Ӭi�����z�����hPٍ�2OAz�*{�׻tEaW��6�es�����װ��r�7�P(n��t`5#eH��aN�ݱ����U�c�K|h��a�k��gU��BaJ��#|�U�Y~F�tV��g�oV'�e��C�Z�dpx�@����e��]P�-���b��b�l���@��:��qP��kܚV��ws<�A⯡��D�L�t�묺'c5`a�2g�%��J�4'�m_���h�\x���m��Q�(����6X�h���#�l�
t#�A[�S|��
�r������W#����"�Y${B�K ]!�O6�Y��.�
�eq���!�s�q��ű�j��w�묃J� Iݘ��v�@��q�:�%(��[�i*%|	)�LN��Q��%�`Wt���$jVV�|,�X/f;�Y���Y��z�5��[۾�P�"�o59wX����&m@�9�;V.�D�E܉![6WA4��c=��J�����JQ�D;��v�v��hޜ8l~�no�L`�_"��h�h���s�-���t�G�Y��1|ip��Dg,=N����\�H��c{��K����ug��2�!d�"����jek��_U����R`[�eދ唲*'�r���%I�ӓ�����E���'����g#� �S��IjX�5v���]K���q�DF������N�7����C��JU��M�e!ǷB{w}��C�0�+s��oQ*�7�@�Th6�$�V�4ĵS"�*�賙�G��t�W,��^l')��x��N/@W*4���kr��y�{��3ghw�h
���7���'8�Y}�Nr��g��9V���X�.Gf���;�i�3�K�����E��K{.h�SrV$�)X���/�EoF������P����*�˜k�P(Dؾ<�y�=��w2#�d�����!��]>9:�D	�0�)!XHw��}M�;w�Yb��R��r�x~�h�*�X����; ����@U��R�����r�IG�\i�V&�M�8Zӷ[S�7�KOo�+�_qNԝ1T�Fa�q	3��5Z�֚Gn�γ��E�^*��^7F�6Ҵ�\UԈ�:�9`0=��V����	E��}���U�Se�L���1������w��:H���\��+������<�j��l#*�ӏ#e;y]�#Ɨ!��kw(k�ި3z��Jܺǰc����)t�Zb�*.�<�aYJ�hBU���c:V�*��)t"JӶvk8厧�����D�����}óz:{��p���#�7I���f�"!�nC�4WY�N�2����n�����H�(\1b�ð=�q�IVi�ŞUs{��z����t�}c�u-�����ڄ`PPb%F�/P8�Ү*��k/����R�7�6�#�[�9w|�8�u�A+ܾ�NiPN�HK��n�7$R�F���1��$z��0[�Z�#e��,%gV���x�*�x�
�����ͱǆ��t�ޣ��(�݀A�;L�8#�(.�ǘ�����cw���qޡ���x����.r�t�f��Bnnm.�s�)���}�I�m&�͡�AF�X˅��+v��4�*��"�\-�=:錵{����eX��y[��e�G+qL�vʘ�9�2�B���F�
�T�K����BV�&1N+�<4�iQu׻��/�W�����`���:s�Gmwax�6-2��%�Gf��u�5�|�n�P��q��rׯ���o��lbP�sn�4���FK�!wv4d�9�[�a�RK�bFX��p6���$h��wk��͹аRbH��p1�$˻�n�6
.n��76ܤ�DL�wn�����L&wm�\Ƣ.��	$%E�G6w�����)4���(H�w]9�;�'69]��ۜ�b*��N����κ���W,Y.�B�N�E�� �p��*�E����w`�s���.�:t�wr����;��tQ����z�Wf֜��]��]O�"AP�ڱ��R��r�o�]�n��=i�ry��1�����1���g��y��K���w�4���ټ��Yzv&�t��G��m{ަ�#��+"c8d�ܯ�����+d���ڣ�Ѿ��ĝ_�V�I9��L3VЍ��k�u�qΎ�!F*��X�Ϟ�C7���=�Bylm���r��/xbc���ۚ�v��{<��C�Kf<�҇����ډYy�H�|�)������[�"J*ebK�*��T��՛��3(��|�M�T��
/��&a�U�6��=�~ֳ�k[a��U�s�&�d6�[=�浞e�>�v�շ%�7���Nb͜O"&�0�t&��ik�3�0�u۹��X}6q�9���޹�K3�]ւ��~[��Ya����ބ��3���noIgsY��~��ΥK�u�E)9�M�է���i�SY7&��igX��n������^��?^�k㠈��gw_:.�-�Zy����3L}�a��Q�7eAbc��]z�����`_�77v����w3�2E��-��ɾ��z�����1���W��Zo��F�O�%g1�Ɲ�'.ȳ
7H.rr9�ۦ�- |6��Wr][�q-5��Dr,M�ʸZ���a�MS�Ⱥ���՗�B[᧚��{�@��fy��Ub���rp�-��v�m9F|�)�q	l_�W<��tˁ�g+$k���Wm�I��y�z�3�oEl���J�`��Mg/^�Q��!���f'Ά>9\��&��p�#�U(��<uwu�DO�eX}��kt��-��&��X�{CS.���I����� 5淅d˧���rb��)�A��y�6�̱������X�$�m0�hFS�U(.�'"�|�X�&�h�(�"��fuz^e	寳�����s���dK.��IqE��ˮ~��ٔ��ٰc��g���Z�|�Fb�6�����3����mӫnV;T������ذ���j����h�s��>����WS�x�c+����l~I;�a-�h��)z��kz�6E�9C�.�=����1���b:���W��WXǀ�Z1�߶�Z=��&]��M_M��t��k����5{��;q�X(��=�o��J��3U��6�N���sj��(�Pk����TBE3��P�U2�Cz`�͒T��xY�xn�E��k��^u}2�w�F=W��*��9X��u�"Pj����-�����{�g:&j�L,�3#]xUh��bsW�b���y��u�K�~��U��6ީ|��u��;�����{�)/}=7�b>���b��:���x���.�>o���x�����6E��(�,�m@����=ެ���+e,$��p��y�{&��}�����ߞ��8�)J�����A@�N+�R\X�5xO�)"�j����ۜL׋}�!��nʇ޵��W����_]���N���EI����Uߗ�H�HG{�ߋ��f�ȑ#t[��K�5Na���A���\('9�O>{��@c����o��ڄ��ew)՗���y�W'G#teB�.mv��'���M��� ���n<����)f	^��[�V9���i�<��K���a���*9[v�&�wJ�`���쭇5	C.��=����b�`���J|X"r9h��t=��MY��Nތ���0]e�4���xg���YBS�egS��g(vAJ�R�����"�qշYC���ȦD�*�0_U�u�g&�r<j9ʝjЏt6�� rc�]Í��~��@k��:b�ף/�]�W��Ҧ���w��f9�v��'\�0ۮ���k��2�YU����fqW�=��-���������i�:ܤ�/44�5�c{/9ѫ�3U�xYN9!}U��ż�L�LF�M�W�댱���������x7Y�77*no:���I�����90��ػt}+�ś�����̩M�t���Doc�j�[��i[�;�o,�X[��AΩ�F����0���Zχ���g=�@j��œ���ί}�����j�!mo]��Oe�����p}&����Lט9QNq�ȃ9j]��������	��Q u�Ӱ����|TT�UwB;2llm�t%:5�=�a���מrؤ�����Ҽ����7����+�[(o�o��U��Ǽ}��5�Fu��R�7��KT|}~�[-�"�/]���%wZ�7&�"g���k�h���vP��)b�}���"��-�xT}�m�PV��l�,�����էV]Ҳ�
'G#[c����G�'xW���eOvzEV,NC�ngلAe4��bY�xh�GY��Nԝ�%���_�_Ͻ�CO5�!oP��l��ý[�'���QL���{�2�L��d3��؎k����r������uh,cÙ����3����oE;f@E��)Tl��O.ڱ��-���#�o��Sh\�a����vc��|�<�f
u�녹��^��^yG3�(�/z��a�������Sk��lk�f}��H�/�f�73�="���3+c�c3��,�9��5f)�^I�X�f��#k��V�6�b}�՝�=�يo.�N�fuK̩籶7S��X������uG����B��.���Zx̬��cn��q�@��U6��y��[�yĥC`l��j������٢���Y��͟[�t9Fez�D=��V���Y�.>+�)�f�VS�L�{psw��(�ws�'�Y~޿&z/��x�Ѫ6��8�吮��ב���7��Jm�^�k:���o�F)Nܴ�sؘ���½�X��� ����B��"�fđxel�}�]'�)s���;o��w9h��[�CL�BW>���e<N���ﾰѧO�;W �$:�P��s3K�\��Nos|�f�����[�����ٶP�	V����վ�n�^2��y߱4p���bt�KqV�X�z_-f�Gd;Ý<{7V��ʷ7ܹ]���U�.U��E)8����������<w0�Yݍ=u�u��C|�Pم�),�1��c�Rޚ-<�����M\Q��O��ݣ/��R���P���!-���k0[�1>$�	�9��c|��/ɋ�o�ّ�J�{�odW���/�|$w�[���m�f�����lj��Oó���������Ey���9�au�����[]!���,��K��f����c��|�o��ۇa�D�Q�
ˇy̠��9IZhE�䘇r{��]��ymjeכ��I��&ƹ���	�̥盛���p���q�C���_mW �̿e'�{�uM��˴�3������Y+3tU��ऩ��R�l�Y��Mc�t,�y�@em�3����q(-_�.AS�s�97Kkr��}��k��8M`�?a�*���nn��r��8��.x֕���z��&�'N��^���E'r�>f���6�Ld[��ӄ�)��ȭI;'^6s��vbuGO���#3�K�<������/w�{C3��K{ch���I*{o���(�/��[�6������������hu&��l,�k-�e%a̽�om�P�^�j�z�ߠ�����.�lwM��W�k�f�X/���ċ����n2^�����͑n�s��17ޤ��F�AkR�zo�ڎ���*x(�	��
RX:�AI�������ў:w@�V�r���N�5:�W���n8[e�ͷ�橍Pٕ��O#u����佲��G���t�iu��ku��������^5��r;%ߛ�GO���߻��h*c�ܢ:A@��^ڔ�+��u��s��f�\LL���l5���y�)JT�[��Q�#���zG,�'^l�H����bS�^-�\;}��fշA�2��~�c8���V�Z��7�[���-[�����������L<�к�K�j@��u$#��7���,Kvw0�U���7��Sӆ�m�/�	/u��
���r��V'�&��������9<	aȺ��C�^�^��(�L�.[�p��n2�=��{���8��Gz�wu�Ҹw�`�"�l�9f���GHX��<J�!v�!1ӝ_��;ڽ�r�ӕ�WXKB����@)v��'��g܅(�.x��Õ �B6��k�k��y:��]y��v��ݧv�S���v5���N,'F5F/AZ�� ���o�J��U�1r��ȚETl���l#^m�v!eP�f$cg�}���}+ސ3��=>��~OA~�9����[��~��0��2�YT5a�U�5|'jdA�*���}�gw���SH��������I�S/o��9������0�i��:w�+����I��5�Fc���yF^r춝���d�]a���V������l��Ȭ�9�l��!�6p� ��3j�q�\W����z��ա��\�z޿J*�A�S��{i�L�!�
��Ƨy��Voun�)����R)��$�Z�De�x��:�{r�w�h1�Z�U��mF��3�S�4*��2�d���Ϗ�H�h�]p���2����}]˸�n�I�i��i��j�e�}��ĝ:��c}w��8�,<_4�A�`�Ӫ���zs�]:1_����W��z�OB��v��Q����S��݇�ѐ�8AOrǓ'AƵӱ����5����i����������������dY����s���w^+��KtkR{cXko�am<��&9��K�]��mSއ8���x��55��X�[���X�>���웡�*�ux�Q4v�
~�Kcc���-��'���ޭ|�p������X]���;��r��W��S��	����v��[@V�����VK��V�=���3�x4;fB,�AJ�lV����R)��K�Ɍ�����A\�]�i��9M�7Z��"g�l��C�k��=��6:��r���v����V5����j��s���5ى��Ω$t�8>Ԅg�`G[�����j��[CUZ������m���C��%�N�}%��(HI���P��9��*Y����x�9p��m2�%�W06�������Gה�Z�v�kM�+`xT����OWu\x���at���扝���^V�}�ۭ3���z�YՓ9ࠚ�r�:�o��v_j��K:�<foVop�I�R�쪳&�]����o��9��+���P6%Q����cj�o&�X˙�;򖖉�K��w��)�������ӡ��^�����$r>^��7�.��D>F�d���K��9MK���4Y�(9�Ĭ�[���!g_�j��ˍ�vS�n��o��9�S�s�¬-�rM��z_f߃P�	}�v����f�����9���eh��
~��^�‶����}�a�bX���,��s~�6L�=����D.t6���]�BR����ke�^wΕGr��˯���>��&����d��G�v�QE,8W/�S ��qxd��.���v��(�y����:w壢�v��vo��]���T�J�|l\��q��n7�m�Ӕg��wW�=�=_��X��l#i��GBU�.0ͭG�O��ZY�:��֫!j��`����ViaI"9��bQ����#ҥ�BS��0T�b����ƌ� v!J�fyҤq]Y�g<��}�ilo���2,\+um,�����[|5�f�'�n��h:�c��O�;īh=|Rw[*Z��:��9�v�b�������v��SK�e�#i�*�X�����v� b>�G,M=����!�3Feqok=��AE��c9Ũ3��NK$�RL�y�c�Z~�I �"�i^o#��h��>u�����פ&z��`d�3,�v���f*r$����wS"}�q	V�*�T�v���Wxxe��.���Q���$��[x-DV^:�d<�vV��i-�0&�'c�\�n�u�[�P�x8��*p��Y\)��*&t0;�٥���Doe��I)j�XR��}z4�ƚM����]�t,��y1���|����1��w׌'�2����r�*�r�W�LX��vzEwp�m'˫`��h�]`����.ƒ���m�A*�a��63Ū�w`�E���WE�2�� =���Wd,�O�iFtF(��Y�˃�jٝ2�I�t��f�v%�G��H֜�p�|(n��`GRI�7���ӹo;�<2Z�]����N�o�ջwڛ�2���ξ�Qsu9	+7�o<K���[��ܢ�����k$�A�N냀���L�.���v��9p׻ř���C���#Չ�-<GZ��3va�"iԈo�ۘ�+��Z���ui[���}�CKmR��(�vdʲʥ�ڨK�qn$��6�zs4���=�Rn�R���sr�xr���7̪o�D��V�Q��''V3��u�P[8Mb�-�}�}w��JF��w���.�5�p�ǵ<\�O\Õ1q���@:�
�_D�
�{��r'J��
�ܜm���kt�D�&����m:׮���}N�tS�wE&����c�,��xq�ز���'�S޽�P�b�r]�^b�B��9�Ҁ��;C]:������а�MG�+�r7Չ�'�����4�,�r�>\j�Kɍ���VNQ��պ�fn�%����%C|�S��`�(qۍ�e�Kv9�з��ak�ǦOi@�1�Z{���yS]�lP����Z6՗W����:��كw�$���uՠM�[#HZ���tj�f��&P�ٸ�{�����WW;q1T��u͕��nQ[�`�;�ǐ*c�Ԃ�]B���0I�/�g02�jk�J�m����<Z�u}jJ*�mA��jC�zS#\Q�`I�Mh�V0T/.�X�!�YY�&5��l_[��'}{t���7�]��7�Ի+��x�Z��:�-b_5�Bvݝ/h�{���#�h�9�vg'�c��w�X��R}�uD��k��g&f�M��}N�vBaC���Z9��66�pּ�g!]�/n��TP�� c%�㻤��r��ˑ��K��ƹ�F��ۧ"�ur"�GJ1ww+�F�θ�˧*wgr%���Quݍ�����s��;�-�sr�����Ĥ�W.�w]�nW!���\�7Mҷws&�E˗n��7+����ݷM:�k�u�QN�r����D\��v9���mp˺�]rحʙ�;��8��.�"����gv�Ww�uە�.\���9ܹ�:-p�]�nXܧv��l[�wc���:�.n7Js��sIsnk��)�s\�s�Nm�;��r�.�s���.n`�ۻ���wwS�Wu��9r茎l��\��ߝ����~�?�y���q�{�_��Eu`��.R��8x]z����M���1͢���;�o��,�7K[b��m�d�5J7�v3��F{1~㎱���&����gr)����<Gm@���7�vn�����j%������z������J1�>.�ͩЕ��*�tU�˓��6�kyg���L�Ny65қI�Y�������{F���_hu	t����7��}��!��<_
���[}Z���[�pQ`oh�n�5ى�1khFg�yc������.�T˨���K�ع�o�u���{F:<5ټQx"�Ќ�@M�Fsڛ��jRJm]	���K=<��V���y�2��cW��z��4&�~V���D�mD���Jqׅ	�|��e7%��������8��\z�v�[�]S��Z�܈<��N�ᅎ�an+�n.[zW^"n2��fiT�2%ڳ�)Gus�:�N�4'PKa��-�z�k=N�=��C�s�[Y��V-���)r��Ʈ�xk��9J�^!�͹RU�+�D�Xa(�9G3b2�NҎ��n�;!�Z2J�����c]Mt����b|�:���Z 
��$���P��F7�1ƅ[û�����mw%J�M���A>��O���ž�:t ������j�{>�;kA�=�7�d�)o�?���h�{�u�ˢ+3Z��X{h6��7�&:}���~�u�wp��e9ur���[��m���x�_�����Z󍢹z*:{Ϥ�j9��q��ި�p�b�q<u�bS�E���;}�q�Bی�(ς0�G�J&��.U���y>�:��j�N�F����.��W�w�g�<ȯ6�:
�=s�y�k^J��z�6�z�$>�˞w�n����>j�7��msn&Kݤ��1s�^���w��V}�B;�y�m�+\Л]����v��^9�%VD�T�K�OO��;��Xe�j,bvbG(�C�ne�s��"$��'z7f�/yS�N2b��nj]2�0� ��|��E����y��U�I��Sv��s=���wz)9��j�w�ޯ>����Vk5G�5tC�R�`@�鲽vv������(|70e��j�;��+�X�Y�n�|�w��S=�ﴣYX0��O�>X5Ӭ�uN��ޫ�N\�<�1��������fcÝ�1�m��xn�%A�0JxUm>�!}}u���ŧ��;Z:�0�딻{{ �f�rbm�O-����%>S/m�9��sk�V�+@^�=Rن"�����̠_H��nr���$e��)��`�q�wm���SY�"U֨�OqZ��9�es��M�TJ��Z�{qvє�Op�,�E��M�g=5\�^�ʥ�U�:��uѭ���ͩ���Tj���ձ��J([�)��%��f�6�þ_�p0;_a�~p��	f��fw����؝+��^0�=oWҹh�܁Cw����jW%5sJ�ǫ׭�<�������x�u-�Ԟc�dv1眶����Daw}���L��O<�4Tw3Q�+k�o��e��E�jx�d'�Z�¶N1G�=N��������� �-����,�O��i�o�2�E�u�J��Tp�&9n�<gYg� w��{'W<�qN;���7F���u]�7��������r�̄�M$Mk��_�/:%�AK��m�j?�9���ֳ���ðDv�!��ճ��Z���w(��[|�-��NS+���s���pW]�k��BL����,	��G�����{r����늓,=|�̾�a�Q^m�;fB,��C��)Z(^N�X�𣲽:+V��wٔ�}�Z7�%�kɾ�a�1�G�H�Q� �-�1��toV��q��K��7�j���O�M�py�5�3��)|�kb���&�tk�l�un���m��kvj��դ�ba����)�nm:�r�9�o�]O"I��4ӎ���1T���c7u:ܬw�_Es�H�u����H�y޹�p����qh3�]im	���.��r�iN�f�x��&��sꋻ�N�毝f߷Q�u����;p��c}l�I,֩��]��ԙ��h�mE{������;����[U�~W�ޖϩ�A=�ha��U�t�k�H5cK
��9&�6��^����2T�`4�Vw���'�矝�Fo�DK5�9ߧe�uT1:[�a���}bZ}�"n7�ד�S�fb�g���Y��OM��Ot�����a��$+;�8>�n^�=V4�be�����̪2��g�r��nrq�m�Әs�Wm�˅�HWb�Xܦ�m����:*'0��Z�'un ��k�GP�r>ܮ4Ҳ�R��ɧ'8�!�K�LLK�g��#gǁ*ڞ�}vU	J�M크5�z=�E	sWP���]ۥ1��:X�շ�m*Q�9�t���#;���e�(�S��
�:b�z]��fG�KOk��vwm����P�>��+�y�Vkv{�=ւ\���i�&h��>��{�m�o��>F���` ����0Տ���]� ���y��ίb㼚H3z�w!��]�!]�^��OD�8*�����}ܾ9�jy���c�9���lㆢ�[��z�W���1j�덹/\Л]�{�u2���M��3:�'�7g��W��+f�D��:1|�f-mw%D�-�<4�=�ڻ�bM+������[�wl�~]ËlFhk+]�5�[�����?N��ʍZ�䧱Y�}*��������=x�6��ى��s�c3�=��5	���S+E����ƹ㶑T���j��ni.
\U��^�'|Ww��c`�WAE��-�z]1V�mԤo`���ꕜ\M�]f.p�`S���!�𤯣J�3�����_�Yh	@�vtm��p�����`44�V�^�i)�ܫ��m��E�i�e�|�nRv���Z��oל���jM�/5����d�~�o`䓫�,ۉ��m��je7�]m�����T.��uآ�Z�z��Xԕ��E_>�s�=�W�,O���I�^�ު�є���[����\�[f����ge`L��	^�J���u�ū��ZY<�s��ꓺ���j�#+:�\��Á��:g��ʙFoq�d����"�k/��Ya������ꊎ�p��,�'�q@E��۾.gkqF]R؝I��k�Y�yة-Q��|�z��t9�O�u��E��Px8݉�yӋ�)�[�t�9�ͯ[q��.��!��Y�֪ʻ���,�v�{4�����}��u��\G/xn߰T  &P����6Pˍ3e�<�أ�f�:��"�֜���ӷA���U��[8i�u���n�R3E8jme? �d��YCrM}Gf_ڔ�s�\.�Y�^T�,+�@��ì��:���R���0���1m��&����@�q�\7�����2�����fKPwl9�ĕo7�q�}W�5ڛ6�Y���iޫ�k�v�Ў��΄i����[���g�*��n_m���r����t��4��X�DoFH�Ρ܂�$.��y���ywC��9�L>�k�IuM_&i�5�,��b�S{ʝ�`R�9���:���H}�u��+ث:�']x�f�����b�yl�󫇽���b�<M�U[��gyP�[cu:r�r��LsY�u�"u4������q��q�&Zq��3$K+�y�X�N[M�o�9���.	����^������-�vi�+4H��C�](����=>^���S;�~���������e5۪�E휪Ps�R�2{���Z6��鼒�'��=�Ke��_m;���R����$���B�6v>����v+�����;�}z[�a���|Z{��GTu���겧tRē�Ô,)�m]]Gc�)�+���b�Uu�)�ȭ��GGy% ��\D����)��<շ][�H�;A���${Bb�Ო�ͩj��	�r��e�t,r����u1	�`n�2"ܼ�=B'ft�NG+3�*��~(F�l��uQU)Q�o1�������]D�:1%�=gi2�h��� �}��jJ�Ӡ[�^/�����;�e��f8�[́o<�Ouz*:wϧ�<[�fY؟H�O۴�Ds�R�ns��S��}ۍ���}�A�6c>��5�δ_Ӳ��u���Jh��(�UK���78�m�6�#�3���9H�mހͳ9
d�f{���'9�UUi��ُk���˚=υNϰ�k����Q������,����_)�3"��;9B��o1��zN��ytdk��4ӳ�h]{��oR�q��;o��ŵ�̛�����j*�[]��oB�����O����t-Wl��i��v%\�L׳i�Ua���y9
d_l�J���s������r����/��V�OA�A!]+k`�c��H}��e��Ұߌ�y��Gٻ�yݧ"�b-%A�c�O�P���й���k�v��N��1��4C�7�G�xQ��X*�BR�VˬB5gA`n��0�{���w���'-[O��f�S�fT�෉N�lf�곚�F��6WSw��K��
��Ă�����=�3~'x6'|�z7p�]����z��Q+�Gq�Ah�:�1��r�n=����&��9Zf^)�n���G;�ی�`��>�뎔��W�D0��>T����Vb�?(α���qS/�G�2�TG�+���S,��9�{n�,U�k���̟������}ۙ�z����3��J�N�S��;��`�r���g:"��f���B�<���{��j�ꋚ."��P�K��rn+Un1:���L~p�n[;1�(�m��5�̞���i���y�n�$�A�b`��/n��Ͼ�z�U�^���]�v�OA��s�\�xd?Y��;n��}>��'Mqd��d!ʅN�Eg��b~3��<㘫�פ��q'ʷŷ-��h���y�#.R
�ɝ �Q'���wS��^U[�}��[3.Q�j5�O�'������=�����sH�$}�Gޣ��E>Nf|�ݠr!�mh0�2Ǻ��bꍾN�1�>�H�C��&�q�|̉�Q:PE�X�ըM��+e���$�Ȝ��q|:Px��{c�[p��,���% ������s�T*Xi�'���0K�,�Ҳ�v��nTs]�$Δ�2q�������,��_�p�a.�|�ٻ��gEt�%%�A;����
��ի���»�N�.�������L�\�>�,@�x1����Z�r�t��)Y�[m^���/kz09�k:A�Ko�eZ�e6t��a�	���������5�<'Rq��ߕ�l�ܞ~��ޔU,�2���:�|��_'�k��-!��[>�̹�v��q�rr@���v��H��~*�7��7�M��U���k�����0�dK�x��;�{:��|��X��s���zn7/..5:|}� �����/����������{����-�x��=#��t�E�>9�-��c����0|�Y����Y�����ߦ�Fh���}�������6�PU����k�~�@{�\1�*����u�����զ.��i�����Yo�~8c���:XD���������*U ע0����9�LKtW�T8�ʼ%�ZQ7��u��4�!d�������Q/A���;Pq˓�����݈J���V<}{[�;�<��/m�����K����ގؐ�gĜ-�YZ�=O�>�l:&ʍ���z��J�e�,wp�r�{�rX��a�T�z}Z:��ꎔ	(��}��~���ZF\X��­���B77�k��z��WhR�;E�i:�l4:ڬ
���G5�������:���i�&�]��@O��u�V�_]�d�͚�����f�l�=].�a�H[n��UvXKjjŁo]^`�9�����/8�1�%�yR����v��{Kh��𐽭��z�;D,�{�R��T	꼼�|�����^%���j0���F�2K��K�u�[����N�
�݅��1:&Ш�q �4�����F�Sp���v�B�Ţ�u<���#{6�Y�gf�z�uue��z�2�o���R��dn���9cs;�fq�8���&��qp�'Cu��Q`�,��*��-�Q5��;'e��V(m��&�BL�/�я�:�+cM��|��o\Z��n��f��hу�K)����!0��$U��A�IC������n�&u�C�^mۉ=����ƺ*v#i�SJ�G�x%N���R�[5С7']��䍴3ڂ`���妕�u�>Ϯ�I�rO(�/0�Or��p��θ��Ge���"���Z���fU��<mv[�-Y��7�w�m�t�[6巸.�m���]W�՝� "�]r�K�OKQ�wC{ظ5V��j��uWW�o7�K��Q��3S�Ϟ�k��:��k8
e͗�Y�_%�o<C�����-0���oR�Z�^nmO���]�e�+q�I��W@*�T�ϝ�ҳ����}��� 5��o�� k�]Y�X7Y���:��v�
���$X�1���p��Cw�G+c�V��/�r������y�r����y�PbhFY�7>�Q�g[��Em����d��e���:��ŕb���8����"Wc�]�1!Zd�J�n�`9�-�Y��,Ar�{lJ=�����P�}W@wQ�[�e<���+�.���ݰ`��!N�5V��:�'�G�ࣤ�o���[�c)敀���t}��Ψ@ؖ�y�d�Y����'����F�'�n_vU�Trӻ�H�ygQ�j��:��J��7Ul�uQ7M�]��k�}W��Nw�7��C9wg"�|:�t�i�n�p�mhB��lnj��d�jj�z;s��;['iT�K����-�m�baq����q%��c0Sf��B�_!�C��fm�4$��j�ܟU���b�� �j��A��m[3wNG]�o��xv-�'g ���e���Dt�k6<�7|��a]����d����r̓r� ;y�����4�7��
��w����z��]�2��l���/勄
}ڮ�<~�uF1�Ao�Q�t����X��>7�o�u���u-��w^"�1lZp7�[ǻ׻�+ьD�F+L�&:T�D{C��7SE1F��z��Yvͭ��:����*��\�5x[ɠv��v��v�"�|Nɽ�1дz�=1l�vة��+�t��8xwe�3��qF��/���/ʶ�M�f�ǼC32���0�!�Ԅzt�n�`=Ck[[��g�p��0��r@#ޏG���jw\�]݃;��74��Qλ�]+����w]� �r.ss�т�u�b��v�p��f�`�up�M�t�ܩ�;���9r��˕�]�9��-u�I�wn�]wrs���v����lTt+�n;��r��g.�r����ܫ��u�܅�s��\��&(4\��4��r��LG9tL`�Z�l��r�D�����\wUҺW.b�;��D\��]1h��9p�ʹS��������K��ŮW.�㻨آ��nh����ɷ+����r�ݎUs���nC��cs��k�Qr�Ds���r�ɮrr.c���ܻ��:����t˜����n�D��������G��N���ܤnR��f��M=f`��r_:���n-p�4�s��ZBJKF�1[YSK���*tSva��N=���=�_�n�s'�]L��)��Z��<�ea_=���θ˅>E@�x��{�j�~�<�����Yb,΁06x�)���Gԝp��n�E��ӟ7'�����'*:�s�z^F��s�.��q��.��)l�l���@����s�=��<_��s#���}Uiߞ^�N�s����q8mӨ�	G�a*���;Ft�/B5�jG��o#R�:��[���-NfoEz(���mq+�ς&���Z��%L�#��;1%m:3�q��M�]�\]�O\｛��R�Yq�ơ��Ga�L�i�5��)]f6x� �g�\�/
Hu�r����1�C���#�}�9zoSۇ�Wtn>��m��]��?�"�P�ٹK���ʞ-�gnR��;��lyp�:|�Oa�u����ݕ��^\w��N�bq.J��]��c&��q~{#&���1��S�3����zcc��dT�p_�ʴ��� �r�����G��C�����l	ǘ=��2�.����]M����Y��0���r*z�9�H����g� �;|��x�<�����w�O�U���m�L
&��k�e��&��s3�VhT5��`Ur	�FT�vʆ��-���;���^�M��'�	�o���{���k>9aZ��y����y�v�����b�7m5ƇuE)>�}�j5���:bC��YΎ�����;����߫qh_�h>>&�|Uzˣ�]t�uXD�C8����Y�:��V k9/HtSrT;�Xm��啢���9E�
������5=�y�z�.t1}�лEp�>���\���f:�U"w�"�[�l�����C�h��g�p_֤������U5q������vS��t�v5��ʉuJf/�BT�)��K�.<�2�|ܶ{�ѯܨb���ɒ�*�o���g�8��,"�͒Q�~qcjz�ߺ�����F�4k�(/�IG=�c��ʹ�����P�n ϰñrY�����=�dY�IO��C-։-;�6��=����`�{V��Ϳ)���S�G\y��]A_��C��Q���&�=+��9���J�a�Dǡ煵�����8��e��:���{玤mê�=2zt ;��&yց�_lɔ�j�J��É��f���N�+�3���s���mހͳ9�'EA��+���ǨR����xd8�բ��3�8�\c�Q���N_Ϝ���`��̋]���W���pS �!�`Z�S���'޿SE<�e��e�kn\&I�˗�*ddf�Za*���$w6V��3�3��7��P <�Zk��Ub��k�EyV^e�*�8�7��t�
���Ҧ���w��nk��h2�7��ܱQF�"�
�ӑt�79ᜧ?�R�R�U�%.Y�и�*Zo�Դ�s�����;2[.=�����I��Z�w�n�Qr?�$�g���d��"~�d�])��H�q�9��!��:k��fEY��x�Z����.g4�~�b��H�,��0��Na��u�n"�p=ݤ��d調$��v�ܯp\���U.>��3��ï�B���G��}��2=�7//�T��t����*�J=���<ձ�U=S8�G58��~ܭ��}9'/�\;`L�<G��{a��{K��z��3��L�N�d���C��Q2�G[T7�U�ha�r��޿�Q�*����.��D ��&x+ۧf/iPj}�,���r���r��[Q�O>����5���w��Fy����v�2àgJ�.N}Z�#q�Յ�.�"���aҮ�L>��j�D%r${`?��^�ab�5��? zq)qî�WӁfP�b�ˁS��ҽ��
���k+ږ�Y确�H��o���َ�Rt�iD��1�&ꊜ���k��^�w�ۛyJċ���?_r�W�n���u�r��=�75� Լm2.���Ch�y
�Z��8�}>Cff"�޺x^�S&k�Ȃ˦�Qy�祐�*Bu�>��!7&j���s��泋PU�\Yf���륽���;J�N��qr��EO�͚jC�^����|g�TK���x}�Z;致B��G����t Ϥ�_OI>�K�1�{�B�נ��/�q�O�&��!�g��s�n<ݑ�i���(��]5��G���߽���vH���c'�C>�غ�o���z��G�a6۸��]Z��:�Ϸ2.�{E�C��s�C���7���m1%�;Ӭ��:Pw�>�|�؋��Ydh�g��t�*������뛗:N��5��E}��&c�����m:7^��W�\Ƨrs�8W�s��m�sѱs�A��&�`k�7wR���!i���ED�����v�������O�g�5�H�<�m�ѿ�� ��`i�����RO@���A����p���X�系Mu[�|{JӺ{��ˎ�G'w��� ����!���f�~y��3���9]R3�CY=ϰ�r<�(;��1�Ҵ�;����W�*�zc�4�Y�������Q�SAW�g�{#��Z�3��rp�;>8�I��k���Τy���O��Z�W�{�0���vV���V��f������)��?�*�uFQĆ�o:�>F-& �^�o7F�p-z�<2�^�8���q]4^.�NU��͉��-�j�v�N*�����R�r���ŗA���tz��|��n��'�m�V�f��� Q׹�G��*�k���r������b���N��'0W�/�yW�J��4��:Lȯ?Gd�D���y�Y=�/�ޞ���]u>;���哢���M�d����xk�z��]�ܞ�1���:��ͼ�����i��8e+"��Ss�凪)�8�����H�(��>�<�=0���y@��3���z�t�3�������z4�x}�2��=�o�Z�7�}Z:�����N�g���q &�=�7���G�cʦw��R��uboR���k����Qۇ�p��|��N�i��L׽��;W8�츭�A��h΁?�foL�P�S��Su�n[�=��8�N�
5,n} *j�s�FE�^�����Q�@�.��)l�{3�N`S��1;ᠶ�]�ݑ���:��]�����iV�7�ḇN�P% %�	�`�譕��B5�罡D�g�2�`)�;�Ƴl\��_Z-����"nu�;u�s;����G�����=徵�_8\��۰_a�o�9�h�{~K��m��4��VW��)��:�/~;�
�U�Pn�~�h��Q����K�'D�Ք�_E�#����U�&8K=�h�+8�p&�Q��Ɣ*��X�o��y*��Zt����|�p�tz����N�����U4p�םGi��g����Zl(6�;��5Y�
���3�qi�}62�r;�����<*nq��z^��Sۆڪ��S̙7�\/U�/�'��������=}�fF�a��w���X�ؿ}�KN��Bߒw|c؜S�y�z��I�br��������3�h�z��}8�R�ฮU��v�w�w��s�ދ�R�.{�j�3��[;���&�^�>U`��xP�������9��'0¸��=2T�>�δ �vq�����=�Cn����2��<��X�>ܝw2%��9���Yts�J�m�V��Sy�h�^{;�Yѹ�&]��p� ?6��{�r���u�ZS�{��W�}'.��\���'��<�u~p�o�����G�,=����q@h�,.�.�7�S/s�w���͇���nN_��V%�7ݱ��_rFk"�&���N�ⶩ���ڡ*n1:��]0o�:�>����C�/�Svv����,���%/�7{$�<���{u�L���o�J�MƧlh�P���m���	��e/w�sg�}e�5����>F��<k�,��e�̏|vRR��%�����h�Kk���6=
�`33�Oh+�U�-�ٳeq�����B��3�!���y )V#�4t���Οt.��sn��P�=1k(K+�'rć�}X�n��fqY�啡M[c��s�]E:̭�e���"2$�[�v�Ǩ����2�t�ZVz��&v���&�D�(_#����[��~�ݡ�4�p8mR�W�\D��R�$i�W�˚�ڡ���������/���&�[�p��|w!�Ѥ��H�uHM)���)���FO)� e��t�L_=,��&=�ݦcrv���g�[8�km� ͳ*�+��C5K���>��w>�i\�1;��\WS�rJf��ƣ.9��7�r��Y6�}��ԇuS��g�ef>���Đ����wA�És�к��~ޥ��S�Ά��Iْ�xhV�ޢ�_�O��dԼ�X��e)~2ON�@��ہ/�+�]��і��f������>`c���[��s�J=qG���:fۖ�w�C5�H:Y=��o�9�:��a������G��5Ͻ5�~�g���!O��z�ZuO��:�{�.̏}��#ג���f��T*�>u���"i�t��F�>}E�L�'��3�J�S2�R��Ӫ�z���k�I��p��yk4#�6�}�f]x���u�2N�x����\2y�OE)l��v9g���>�H�Ʀ',b�AyC+��%>;wt�!+��[:�9����`^r���vG\�u!�7/pr�ǩd.�(�U6�˭��82�+��(L��'Uů<4R���9�-z��v�i� �	\��U�zI<b�b���WE�VMu;��sz��s�b�'�%b�7�/a-6?���5>%�����qʓ,r�͏g����/�sخ�9"\+���q��N���]C��=�NM�j�����y�Ŋ)�[�+��=2)Cyѭ����u${���A�i�ۙ�P_��}z�%lo��}v�{\�X�~U���;7o2�G�2����D�s�C�!m�7h>8''�
%�J����P;�BI�fo�~���Ì����+��n)=���j�G9N��y�#.R
��l��� >��̗9}�ExE{�j�!�¶��g�~�Ucx�)�C����!�g���ܜ;y�#.�3z��R.2=8i����fZ˩�~�B:T�O:�oᲙC>�ы��z%;HǢ��E��=���뒜6#�����v=Cߢk�<d52tљ��2�#Q�q;ը�8����{#WZ��L�����h���3��t�i+��d
�j�k�N�	��bw�
�tr�+�ozPs�A���~&����C�z\����j�-���Ѝ��Ѡn�x�`��0��N����Z�W��-}�M5���t���s�k��yx#EU�**�:�yK��yYAi��ĭ6x�[c:�2�ur�n��e>�|�LI�vg�㱔�?9�"���_�t�l8"�ՄÛ�0g��@(�.�/A��4cywm	SK2��Ȑ�3_lrj�-��<V�ϯ��?6���q�n#S�cͪ�7��6ݰ4�@YV/_�A����i^���ގYf7g��c>�
t����~G|���m텑����bt��w0sa����7�f<9H�ɧ���I��
?���X:;le�]KIӺS+r��򩧦=�N��������1u����~��?i����g�q�?O�&P�C'��82u~'=Ԁ��ϽyU'�
��;M߫�{�NSJ.�_a���q��c��p��Q9�az��(ud֝�TX%����˾�.ߪu_���Z�������M��*�}'EG��8n,�_
Ϡ��+�wrrl/v���c��l����wb����[�z��c�>��o�F_�r�:j$�(Ǽ6`���W�^�\�\k���I��%���������F9��ۆ�}MS�V����x����Z#���Q��di��#v���S�:���nhNjV��5�ei��(���:�j�s輢d���
=.x��`�5і���f��EF+�g��p���s�k�p9"ʜ~�gVA�뺹�����z�y����z�jݒ��v%r�es�7�ξ
x����5vוW]�v��8��Kx�0����3z/����+���sTw%��K��z��ƎS{њ��B�#�z��I����X��Y�N7�����3
��F�� wTDL��H����3�G^'|4Pc'U���s���{���ξ����Нn�q��N�j��G�����:W������>��x����]K���܌	.��\K�3��m��?;���2�z�����B���z�^k�uM��\V�i��P�Q��������-�@N��ғ5�J'FC��Zߦ����tlk�.
�
���W�z�����ZoSۇ�Wto�y�%� c��*��[
�t���:���y0����tm��+���ชŶ��v���W�	'U�:#�ro�����۹�^�[���^���N#z���/�ޔOG�.�X���>�U����ۗx�k+ɷG�^:�Շ"����J�)Y�k��2�(W?T��D��f9М�
����J�<�O(����4sӸ�����i���hzS�Fr�es�Þ87��#�҉̳0�k��kؘ� ��3��})�|��ۙ��X%�6=�?H���7'��1l��F�vV���Ϥ���%��� nk}ճ@�U���+��NƮ���@�4���o�IW���|`&[�6|)k|�=�-u4JK�lqWst���x�K�K��#��16�R\ky�5X5��F̸3A��¤���x�6@mm�zetu��I�������Ue�����:�]W��T�Q�٠(�>1ޚ֫�&kV���v��D�fT։��Ԓ�>��ܚB:�U�I���+�ڹ�qYٸF7�t�������|.���f�u���(iyW��k�x%²C�:��V��������/����9�l��ř���mlw�j=��]���X�[��ꕭf���"F�ӱ��F�;*X@��D�r�uqXʸ/q�2���<��Km]��(�=F,n�Z�4c]-�r6��u��HR���uL����ӅS�����	X�\��^Iu�-��P�5ji����n2����tfo��2� �a�5{+vQr�j�!wβ�a�Ž�:�ӡ�ֱ��C�{�N+�&uFp���q͹r��rStɛ�B��Q�om�-5��@�o�_*�Y�_d�F��Nk��.�,���d+L������N��i�G[�y�Ď9�ve�����1HiT�;<�]>�����j�`��u�2��ÉZ�:Tn�-��8�2s���C&
Eb��gK#xn&�ı�W�[p���K�Fv��̫��9b�6��o�-�m�]A�v7��	J�u�
��0��{�1Z�u]
z�	�R���G��չev,���޾�C�@#���.������4im�nwT���C��:��x�5|x]X�]i^��r�I��^c����˼�Z��{ع�DX%�	owe�t"��V.cmX�W}������E-W�2���ӭ��.�W-��(��f]�5BV�{��j�c,��;��S:���R�-e���W��Σ՚V�Hb.�U����]� ;,��x�[�!���>��^}�|��"e1د�W	o,S�Ί\� �[{vk�Xu�ڰ`�� ����Y�w[{�dV1��\���}��Ӂ4�q��\$�w٘9�ۡ}� 07�5��(�"j���Q5o�wN���䳢��6�3/B��n��f�ޜ��Y|ڋO0�ѕl��ku�g.�����@�<�2�gj�+\A��"�,`im���'7WZLo^.j��ҕ�Nj���J�S�%u�.!���>W�+�h�[�?���x�+5)����0:r���9�	 [;�74:wP�3;A�х!+�t���i�e�Jj��<i�x�Qb��;���#V�e�7u�^��ٜ��Lv���,>��JGm�ۯi�)s�Z�֣�]����'���z��V	ݘ��]��k��;��$e�X{$٨�fr��mo>�}�+���y�z������!ƻM:zY�kqg\��*p$�dnV�k͜�V�͂�u�Vҍ��q�}[	��wbq솞_S$v<���B��Ϥ�w���7ӸV%�V�����U@P�$�(���;;���c�uȐf��]��P�m����EDk�1s�����w\�tK�;��G9sB7.r�g'nY!$��9�h.WJ���+��ܰrwh�J1@F���u
 �.]ݮi���:msbGu�u�#q�X��ۻ� P�4�.�2��u�r���)ݧ:���MC��CN깊"�l�wTsr1��r6;�;t#�����t�"J:]�nPZ�5;���;�1��+�&�Ą����\��]7]�H�X�a��nh�9�&+�9\�Q˻�����Ү;����ё";���)���Ź�d�ˮ��Ln�%Δ�Q'���X��;-��7n=jwZw5�=�7+��x�3+A�1_}܀؜mf�"�u��Umj���۬��v�*��mN<���_���+]t����mˀ��̰�#�M�r��܋w��S��|��(��q]c��F/s��[�q��N�KØKG�O[��_�j���������y�ea�r�����Ra|	��Û�׵fd�mq���3�2��nH;QP���]3��z��J�MƧlh;>��l+PMx��Y���FF;oQ�	����0�\�5Œz��'�{�ȿ�줧�n�_��:"f���\���{�㏴�hHs����h�C�8z���p�T+�\�j8���!%*�}�1�������2�'�ڌF�뉿���A~��r�K�23a�!5
d��� JM��2.��u������xD8���e��ظ�m�v��9�il���[u�#h�Oj� ��Z'����7��I�,��2�p����F��e3x��m�>�Fӗĳ�3�KF�E��bj<�
^^q�v��� <S�H?�N�����9�k�%\��.�ޥ��S���1���=�ժ}Xj���ӷ�xg��zv�&=�/�I����%��DJ�J^�i9J���s�g��>@�D����2tP����lJS鯹�F�Ú�d!pۣ���y��W�qAWOi�s#�#�,��ܧܮ>g���q"k�+�Yԛ���P� �=��9<(B�`���nx��<0+nZ��;���
�t3� o�}�f��/G���~n����w��PȍyRl�z���	�1��0�}�r��B�KJ��/0�6����cy�>>���3=�w�t�2=�R=d�r���I���V�(��3#<�v{���8�둒^㑝-���VǕU=S9�sS�wPv�ׂ�\�O���{UB7+`����}yA��&W����Ua�y���ʁ^��U&Y>�8���q�Zw�y߷I��uO�U���֖��#�%%�[�����t]�?y^)`u�l�I������'�"�0���V�q}�|+T[�<�41T:P���rn+UW����vS���b��wkԽy�H�x܍�7M��<�xc�}S���$�0���z��۪�s�y��>�q�����]ҙ�q>Ec��^�e���z%���t���A��O��
%E�UB�G��:^ʮb��͎����\W�t�-��f����n%�x}�9N��KΙS(t
'}Jq�2���/�셖f\I�${+��2�^�Ucx�)>���n����3�q�8v��vFV�C��3�j]U��D��&���f�}�֝��U�
�Â����%�)����wmbI��$s�{�u!���%v�G_�A��m:���r�1����?�/��WOh�I�X�2��8�;ֵƺP7�r�]�:pP���obW�5f>��ϯ�!:��3�=2��Ժ"e*�ll�P�Fs������#�m�oo�oq�N��j��{rT�.#y�N�:�d"J��S	_�h��<�h\W*�va�}r3�||��N��k3�/"����YG��q��F@�v�M)d���z��/��7��k��vMPr_lud��Z�ȧ�n;z�p������2���F� ����5҉ڀd-7�����7L�+T��=��#�R9N7n��Om�}��7N�R�00�*��k�H5����^ҟ���t���=�(��v���w]Y����Ҹ��F���ruZ{�N�s��~�:߮��x읧�:���a���33�%��c�d�w�z�ˮ����۲���W�B���=:�Rf��U��F�r�eY��߫�k�lϏ}>șc��
�*}G����糩Q�}�aU�<�3j��������3w\��1��uo�uc7ѵ�b���8x"}�0�_	|P����L� 5�!��=�K��9�ɗ`8��H����u�ǲ�(�9��C;*tݖO����׌�׹����\����,\zb�`l?M���&m����i��+���sj�f�e�t�����,]>��joc��5�M���s�"�]>�ީg��x�]dCv�oyA�{��0���'5�Ĺwn�X6�Mib�:�;Z�Ũ�[�4Q�*�ͩ�Ғ���u���iwb�vE��)��r��u�s��Q�ꑗ��$�E��lJ�(;;���:x�����e�9�&�ۖ%J�Dit��!���ᾙjXމ�h�#�{h��s�]�G+�r�>q����3�O�uC�����u2�Subo�JޟDk����Q�i� S�W��g�=CTe�3�.ϣ�����`t�3qe"��1]k>����������AUU��q5�.�ߔ�v����;qn���ꑅp.J5�A���Kd�l�59�N�,jX�ݞ~�om\\�,8�}lz����n�p��N�N�i(�,�:LL󭣯����H�<�(��2�'��w��4rj�P�����D�� �~wJe��=YثM�O:�2�o��WVѺs���7�7������u��C4���P���k ��nT�q����}7Ը��f�O�}��Uש#�}�+M�{p�ڻ�q�<ɓ6�alh�53e����c�==^���4�>�6�9�W=��-�/ѻKN��B�I�񎄛��"�t��������
�tB��yz����r���ߣr�������s��Z�I�l�xW=2Q�Z{�7`�3F�9"���)u�Z#j=S��k�!���u�Zq���SO�='	�M�?-���_nhέ�79�.�ձ\\R.��y�
����v�;�7^�����]c+����\�I�n���]��d���{�r�pq��]��7C���]X=y^*9��������W���,�����9P�:�[�n�L��)��@
�>�<���3�7\��:��}���?T�_�(��3Ƣ�ҵ�7�܉��g��%L�u2�=�Xcܓ�|�Sr}�1l�Uý�/TŁ�S;��xr�=�u��$���9I��"g�5z�\V��;E@h�̰�9d�<��n�ފ}q��﷖�$�f�)q�uVڱ!�c�I�q�Iډ�	�
�j��_�j�������it���:�;�,^BR��{�����zm�ۅވ3�<6��ȷ$�2��_6������Q������h�#i�Vc��_.�/B�3�h������3�a\�ƾ�,��e�̏�����רo���{�u3�'�+��[u��SG�I����U
��G��� �!v5�&�Aw��ȺẴ������Fq����n%�� �_npa.:���W� {;|�����<4�L�R��6=��FY-�J����&����������OJ��08 �7V���v�c���+܆���g��5�ݬi*.[&��{��MY��Ŵ칓OM�Q�K���.��m�4�����b��/��N��
Dp�ח�z���bH3�����7��F�'iC����9>bw�__���Ʌ�����8eǦI�l��;$�z+�qѼ
eF>5|�����,��̪{`gkkk���zn\�:�`��fEqGd�:�*"T�4=J{gJÜ�B(oH�/����=���R�/(Å��d�|ܸ��FTl�'�'b�,��b�We��e�zi�]h��>J���۾�}4_���~=�n��:
f���w��P��{e��=0�a����e�j�#����!������+%#���r���:��؝g�Ճ�~Y��O�r�y��U�Y����C$���h=�|_�UC�K�2��9�3������g!��j}���z�mge}��
����Y�/\�瓀�ˉ����"�U���O�ʁ^��Re�,���6WXJgN\��]�Oz�D�V�狫=i`��ټ�/�t�c���J�S�e���l��4��	�~l��уc����}��Ӟ�§�-�	(��eW�Δ/�ڧ&uHEj�/oG��Q@�s��)L���dzeU]���a��ci�Vw]�[��Y[��{E�����M�܁^ưٵ�\��铴�}ӻ{i.�����
����8-�;�7��@R<�Wnp|-�ژ��W5�X��z{���thmucx�j��H���`M<pʤ��Hg���z�p}�>�+˲��I�2ƌ�q����c����.gWV��=�r�Ѕ�[���h��n��O�G_�����<�-JU^�ʮMG��q��=Q��|��%��on&��j�s����!a�y�#.R	Nb�輯G���:�mےm����L�2�^�X�>�O�&�����3�q�8v<&�X�)�{gsp9�ȼDS�&��C��tǪ]?JU�ޙL���3�n1up�$`U�f���鹺܊\�}�|q��9��&�'nS2*�]6ja(�#�y�ОS���Ϧ<��٪>��ٶ.\�X�B��,��3���Ǡb�Q<Q;�>�N��}+i�z:,�".�C<g/b׵�˰_fM��	�W!�������2�����}҉�B�]�Wm�{���c�&Mue�n��>���K�˝gkv���=�=��>N@S�7l.��k�H4���M��i�V��J�Ww�. 	�����N��J���t�7���;�>�M��r��n��1��K\��ź���6�v���G�)�Yan�4�G|���ޮh�ė P������審�[ҕ�٪���Z�u�r;��X�Ծ�U���VJC����?�������Wb��6�9E�Uh�\ �{Z�'=M�Jw}3���_	���H�iw
�n^������ZedQ?�?+frß��@�W�;�Y_F��*|O�t����v>��k�"2����so}�f`8�Bڣ�<9�N����5�#��,���2���d�R}'��NgJ��=*:�k1��+^Ȼ��k�s��Cuc7ѵ�b���8o�'2ʯ[��<)ً
�K��)���~��3hy�\}��3#�+N�>�M��<=�VN�����e�V\��v�����q��Q�^Wro�P{�.�B�anȸ���[�z"��c���_v��b�<�ɟ%���U�$f�ě.M�f��iɽ�BQ��J��K���'���)�c�w��W����~@�q�L�T+�������f麱7��oO��ei�����7���c�{�#}E�4�n�ϑP(>������'�����e"�*�g���(q�IU�eکs�2�V�t�hk�Z㏤��7P}�ꑅJ>� w$\��H�y��pcޘ����Vq8��2�[�g[j�E�m��t��㸜6��M#%��	W�t��Ds��U�!���{{ҫ7XO��՗������St6`�+�n�%;�u�;6�qn�v`U6W;V\�	�����\��H�=�f�8���@壻Nu��/����ʜi/[��	O*ef�-�z�Ku�|GS�Pd�ĕ�V�ڜ���fz��O\_=����旹�b�]�95H(r�~fp"[s�o���&�˙�g�=�)�&����+!�H�䉝�tn�Xʸ�ۄ��h�e����Cn��f�_��w1ݵ�j�s��k�)GG�?,D�PfW�Ǣ^�
��W3�}�+M�{p����)�L�2@�r���͋�T�X�.��/�&�a����Cl9�WS��~����I����f�6]��}�+}S~c7�z(�F;�'���9@���囏��3�q���=0��VT�8.+�i;�b���s�Ϧ���X����^���F'#\��Vdؑ��l�3�po�t���Qa��͇a�{E�U��*@Z�a��z��:�.uc4�rtW��G�����Y�k�u=�2�\څq^��qS:��a� �rO�<�Sr|���P�-�� ���K�p٪��/�K��� 4[K��[>y��YP�P�H�ޞG=�;qkb��$_���s��_H^~����1`vh� 6�x8'B�V�9���BT�'V��`���5��rg��,z�Z.�����q�G������j�"�Q8�djN8�p�J���w����������Q� Q�h}yв-�/�;)ǽ�KP�&:���#4s�Ȟ⫨�o�H��c�{'t�2�g@�.M�L�c7�y�7���س~.;�#ފj��7�8��RA�P���]tϻީD�u�
[��O��_g{�2�Kz��p��=���6��ϙ�p.O��=FP �9���zUmH���gp��f]g�⺉w�'�.%�x<�SG��=~u��T���(��D�|4+ܪz:؛����p�3[ZM�s̼�1�=�\Mķ����>;�֍&�x�F�Ω	܆y^�Ot��7y�틮���)��D��4�/��g�ƣy:H��ϴ�r�`-S�G�=��g���e�~�<mp�I\n ��F��2�p�����F�q���>5q����)�;r�w�|r�vX�ZN�3�%z�S2=��31��^*u��=��z����V_���ک���z�J�m껣	�fM�r�kBcٲ�d��(��酷�	~1Q+��=���櫻nf��q�'�0�)C1UX��wt.<�37,������*A����Z��MI�RV��!䗆r=!�R�|_ԧ��ϻ�������T��r�Q���~��R=�Z��g����򲓾��7�Clc6�ܴ�'V9W��SP���;M���'�mL뒱�����W&�+����,�'���/CfWgr�s4Q`\,*\���4)��u��aU�nst8r(��;�Gd9J�^���x�o����94t|�(u�ڻ�����w����E�2�<d�|�������!�������Q+8����|�n<R�W��.���ŮO��{91��V���˴�eJ9��9U�=��4m��؉P�Z�uJ�V�kkAJ�i��F��X��A��7OM�Yz����gQ�����|]��)Moum��Y�+V��.E\x�n��u��mW�M��ck�dL�����ZZ�Z<�m�7���O�^-����^��6�R���9�xs�(�WlD����4m���3�yݒ(,	!t��!\)�@e���G���0*���.�d�P�Цs���v:���֦�)h��'��͈��BX��h��携`������2�-��O$��n�tt: m9�����y!*7��;~Lk/&ɝ2%onQ��_LNb�O�m������A��2�Y�+�wt�GPGb�W�^��/g&����*�@��r�gC�F�s��4	h���nj��'N旛0%;�:�Ch�\����F���$�aό�Y���~�J�����^0��E�����|3>��1��].7���o&f�����Ar���یwn%ǟYm���zet��U�1��1&P�\�r��+t�[u��ť|��C��to��8GRR�]�a�qb8u�� ּ]��q��y4c��Y[���:JU���y�Ý[�=8٫�!s�b*m�f�I؄�5ս�����%�� �2�h��0����f^U��S�5���OX�Oპ�n]� s!-�p]�����Tx �Z��S#.����ɯ��V����V>L#1�ӗ��r�B�P�m��EܗA;�7gh�:l�	�ڶ���q��	��H7l�vb�J)}h�Ho�ƑR�6��0v/��#�`M�f9}a��F��9�S�us*,������Z�A6{�������!���wtd���F�F�G,���י;UlK�dĦ1Á������]�H�Y�!��*Aj8�wn�7>G�9;��6Z��r��hYӰl�ꥨ�%��m@S�Q�0!1:e.���H:k����QS�KCp]s���\I�&���aᲝ��8�'>H�B<`�n�ʚ@c.3h�ŝ�K����7ݸ��A��0���0��O�[���#�RYΜ�T(; �q���a�]��rj���X6V_h(��W(��ϊ��ե����b�QaR��E1����w�w:�[��^Κ�������`9X(<֕���%�R\4��.�c���e��=ӝ��W	{��R�(G7�3/;�6�ge���B@"� ���r�r��I0��@��v뮎u#;�WwE�q:n�\��Nt W8��n��š�܃����I�"nt��\�#64N끧v�75��ƌQd�nnq�e��H�4��$\��.na�b�&L��v�iΙݮ�n��wri�TC��b��3"�+�&�,�3&R�D��).�ss9�;�"N�11w]ݹ1s��!#K��wr$n�WH�ȑw]&2I�C!'qt�\��Ĥ��*A�I��Ӯ�\����	F� ɧq\L�e1��;��,�Hw]��B)��$�J�	0" �!�r��Ds\7w`FALw]�I�A��lHʆ�&!�H$4�(���@
(}�����_q}}MJ[wp�vƽ��֌a�ٽZ���q/2uŋ7%����	��u�N��j��N/��zz�����Nv�:N�%���̨��+���+	���L�R�9US�3��sS�wPuZ��&|�O�"祏vy���rm�=����2O2x�L��|��,�9����g=��W��`���^/�ۍJ�{�GVi�w3�"9�×2����ۧgG�*O�2e��5��j�W斑Z��\xN�=-P���Q�3�}e��e�<\`��ro�3p6m��[޽��Y"q�>h���9`��8t�z��K�{�>���4'r�f����`N��(m���V���S�^�D��K�!{�-�=��r����ӣ�\�>aWA�^���V�ھ���I2��t	��Q�[I���ĳqM��ܵo����|��Zo�R2*��]o�绾c�����|=����k�,JX>�)�Ucx��O�0��Ǹ/��_�A���Zngk�h��(���>���Y�O9�p晚S �Q�G���)�}��L����]<7�q���nLu-���V�ElY}�^��9��n!�q;n���J�50���"d���;���%J˾Q�w�l���Ƨ��[:H�z�A�(�B�����gr��.��1�Yz�Ѡ\����F9C�y:*Wt�6s���Ө�Ǌ����J�;e�V�ʼ�sNV�]Υ�]��m(TY��uv{���� ��*�ޤj���oX�2L�A��Zs;6:���޹q������,�β^�9�Y=B&B��Oa�F��=�F�ON��8���]l��ߣ] ��j�1m����2_���*<|��A��D�72-X�~���ȁs��p��HFp�B�
���?m���`�M�j{ly�WG��
z���*��㌼�\�XSN�sp>��J�_��t
������k�A����@j2�r����������{�nW^�-W�^�pi��z��/&}{(4}(u�2p+��Le�u-'O�e3q�j���P}�6�=�K�fa�jÑr����<��w�M�ϑ����qg'.&X�P2p+���pY���ᧃW�Z��� �J��x6�4�����?0e�#��uc7ѵ�b��S��'��zP�5QyvLǽ��Ͱ���qS�X%���i��i��鳾�\2^y/iE��߀��nV*}��y�?K=.=��ڎ��j�NӐ�.�B��h�S����B��V��ۜQ�\�5�U�u%ȧs��5W�3��iɸ��BQ�Į�{K����2���ᾛ��t��b$=��Hl�hT
n�k���1v��RYĚ�Y��.��:w ^��/@���Wa����w��%l/(�98�*�CS�Y�è�nޕ��6ۜC<�h���o^v�!��@-�|���7(�;�x��ӛ�ҁ����%�Y}V�r��i�ͼ�{o�Y��]���_�X$�(�>�W�T�����7MՉԩ���.C�ڧ�yj�H�m��;o:�o��p�ƺ�@\�fn�Eb��o���
FW�>�P���D�KB\N;���;\s��p�Ǜ�9pꑅp.J5�t;��/�)l��-q*�]�O���=�S2�2S���^'|4z"[V�w��ru�M�<w�˘��d�\@Jxo���T7U7�U{݃ex���kk�n)�2�!�X��`���"�IN����h�D��<�J�;-ϕ�7��q��F�IJ�to�\v��p��h�e����i�`w�W �R��vf�*.C�]93_9�ty�
��������ⰭOnj���㹱¦�gY߭V����֓%�m���b���2k�鯏����_�=��b�b������T;�"Y�{���s�.uF?�+�1�Ĺ6����7������+��xpo�tz������=ۦ�К~%8}L=ʯ7�>�{�N�9Y�U�V6�*(/������`�_c*�U4��1=����k{w��^#-��gm��:�bڊ�]ӥf��4���b�l;e� u
�J�f!I�D��^�i�S��z0T=�ه�û�n]vo�X�ݖ��OfT٭���n�ܣ���yYA������z���w�3�|C�1ҧx��:�s�ր�}lzS�Fs��\懰��訏?T�1Ѽ��e���Y�WKa�3��YU��Ua�����F@rN�r�M��;�ų膕p�6��=�p��E��R�m���1O��ܢxe̿vc��k���T�}�,+��M����j�����uV�[5�����q����nN�rIڙ��L�W�mS���T%N'4���ID������z���Ec�\v���|ܶ{�M\>�i����RAڃ(	�_/��}��O��4U��Fm��9�u��M���p��=���6��ϙ�b����=_@_F<ٞ����E^߰;��̇�N�-��wM�D�ӯ����c�8z���j�B�%�9�;E�/�3��zFXb�3&������Y�TgO�'�[�p�~��r�K�22���n
��t^NXY}�rW	~�;, ;�>*H�J�+��&=��L�o:�(���T]�o�@��z�=���/�q��@�>FQ$�9�#pvH)�
��Ը�����q����MP�aU��;T槷'�z�-W��tN����'|�p|���m����ű�׳��
�q5$Ti8�场ĺ5B�ޝ��ښ��Oy%J� �x2����̳k�hh�±�� I���wԨ��|�y[�r�q@���*�˘���δ�G����'�f/ĿD#XB�S2*#�;4fc��:�
:�sϴ��6�aT���������xZ�e����]ы�N̛N\~F�+e��5���lK�=�ܭT�kѽT;9���=5��Cn5]�!����t�e�sc��X�yRF�'����*��U�k�z<�q��a�WVa�����w[.7/-�s/Obt��;�:o���y������^������s��NT���ɇ��|o�XNDgJf�-[�UT�L�1����Tå��]�;�^˳N?���I���\|W�g�z�M��2Q�6e����c�=�]����,�$���ʷ�`�����~��S�ݮ��1��'��ΎڗGF�iPjkq�״����ywZ���2�|z�N�,S����]q��Y�+��4/���t��S��\J	+������������J�iua`r���%)t��A�i���T񸲉;n�H,vG��;���%��pgՂ��*s���%]%��Ż��z%���1�n��DO�Gs�0��o��Y�:����7+"�IA���ۛd��d��:�]�}X��7I�vJd'���L15�:��kh��m�N�p̌�b���Z�v����̙���2��̉>���r��{o
�p��uMgQciմMGK��{�.�ǌ?��'��s�Ҟ�"��۸�n�ۉ�����9N��H�G�q�J���~���W�|�u� }5%0���R+ت����z[���D�����=���m�uyI�6��>8���ni�2
= q�tDĥZ������S��T���jZ�]��qRз�����C��&�q;n��
d���S	_�6��<�hz����-\���^ƣ)Y�y�h:�Ԍ|��C�9}e�}g+��F@��j�j:Q;�7�*�@k��H�q�ZQذ�0�TgǞM�K�W!�o��\4���̰5�����4��T���3~�T����OM��&`��EJ��>˔�׷n��Om�|ګ���-�
X-7ެ�x��#�쨼c7J�D�����k�,���鳓���<g�az{�V��ܼ��N�MW2,�%�0�٥oz3�o��m�sr��Pu?]�/&}{,#���^�2⺖��t�w��H����:�f.�T��]{b��j�;�S��*�:��{|��g��99s,~�8EO���{
T?�P����~}�n3ي�����p�]��Ҋ����遃�\�U��*�u.J�[�z�3�{��|�g�-�
�����G��fV`��!�u:S�]�N2�뺫I\��"�ջ[ܱ����n.x����&��	ؙ���`�k��SA�����K��ͅ�5.��v�[�3Oĥ��<��CUI���N��C��ܘ����!/�%�^G��L�����,g1�yx�k:8����Nk�Ԫ�����+L���.[9ԫ�i���Q��N��Y�	��5X�Z���q9�#�5g�ֻ�7����݈^�vEǔ��r�0�]pcgw��3#������ӑ!�y��u��'MIl��z�]lӓ�P�w������rY�ٚ���f��}��`J3,���t���s��'��	;_L�!����RR�}j�qMՉ�C��;3i�n���3y}�@�<��HEi�=���θ[�>EX6������8�3�)=��׼��qV܍��4_��������~t��}'�y���ꑅ@�(� ;��#_A�q��k*bk�ڶ�K{d���s�Ύ��;ᠶ�_���N�Ix�'�~t�&�(�{�$�5{R@����&� ���$H��tlWKE��C]�Y1�`'����_�fp"[s�G��Ld˨՞��WN�8	�>Q/�*e����7d��{N�Q\r�7�:ј��]n���rFm�L��X��
�v��ۃ�E֜������4�,��&����Z�y������<g.<«�dx)��-�惗Ľ�b42�S�der�ׯu]9���������(ĭ���T]:��w�
�,����;y�[����^���##"�h��Jm�eέXs��+\q�T���J'E�͞��pVDW���;�a�On��XԢn�ue�KY�ܽ��t�&�m��]��Nr�N�����Mv�~"}l�vHU��=�w�w��dR����m��1��✛��^��F��|t2{`zau��)a�9�ҡ�\#����r����N�v�;�r���>�br5�(�V^W�
���{�s�&}����H�n�=!�ہ;��z��=8�Ԁ��ǕS�Fr�e{�uc4�rt:�P������^t�)���o�����e��
��Xn�S'��@
�rO�<�Sr}�1l���j-�iz��ƻ+��~cߡe1^������=�+�����RwnT��e�x]2wޤ�;��R�sw�{�ot��j�ee|�og��QC:rNŋrI�.�KG���%R�y��s^*�[��Â'4Ǟ�vZ�^6] n<�2����KUxϴ��7�� �@@|PU���y*9���zgu֟]̢����ާlh��t�z�Gn!�p��g�'����=�;�@1l��`�@�E�O�2_]�b�h|�,?�3�+ija!��%	����Ry�׺ ֻ|��,JiǶȬ�gqAAn���v\S�����FqΈJU�zͧO;it�ﭼ2F^��6�����$u������#���V�B�E�Y��֯K�2p B�����P/�`�dYs�ϡm�K���h�Zu�5����|w�θ7
�B�=��Z�k'����(�31�`�ZM���VdQ�n1>���o���_��܈n�i>�������{}�Y#}��ˏX�"�U`�s'���)�r�h7eqy����h���O�l��%����+_d����M�ӓ�\&�@�s�f��+���H��&%:�SҸ��2m��3SR"�d�����.)��}Fۗĳ�s>d�B5�#JfG���Ff9�M���@Ψ}7��w_�Gz�Y����ju!�������&��_�����>���Z���'�G"l�����}��a��������׳i�W~y'wB��t��� ��?`�z��콃��m���H�^~&Xل�Na����a��Z_gu��r�Lls�|}�'A��u`�G�q����<q���exX~}��R��Ù�b�O��S+	ÜS+rձ�UOT�lV������8���Jܸ�uG&\���nj�8pz����oL��~%ٖ#@y��	�IsZP��;�YA\�.�����P��¸_,�kV����~llK��~{���t��l{��y�I�:V�y�RWJ|�f*�_E�lm��j��~@����ًz;�R�x�]v��ebo8q��Z(��gto��CmI|��v�����7����W�>ӱ��3���×���3���?��Z��y$��Gr�W^�Jx]�9�����ʓ,S����\f�>U�b���7e�.�w�@�=5/��O`R��D��Iuʃ+ѥՅﰺ`�8r���l��)�ރ>����2������B��ծJ��;$��F#^3���]S�=w1+~��b��x=�KG=��Z� ����z}Z���X7���y����$��0�L�
ⶐ��Q,�7�KV��!��{�����F���=\'2�#(����e���6OWH�Ԕ���7��[/=��9�?���P��:o�L�g�f���\�q�9�þn���9�f�L��tǋ�.%*�t�s�6w��s73��=݃:�T�}�Lw��HǢ��E���Cn�v�uLȯ�L��f���Eu����z�q�no�]9���A��k;��T������|�q��CDW��AK��WƟȃ7n�~ZK�D�"��S�b�Z�R��8�7U1^iS%�.#x*��{������խ����km����kmڶխ��mm�[o�j�V�����V���ն�m��ն�m��ն�m��m[j�����խ��[j�۵m�[oͫmZ��Vڵ�����km�=[j�����խ��um�[o�-m�[o��Z�ߪ���������)���texe��9,����������0��<�lƅh�h�B�jZ b��D6Ѡm���  AG� ������Y��њȬm���l��L٢�mm�L�5��-�	kl�ʶMY��m�����<�m��lm�Kh��X��X�iJҶ�,3&ʵl�ҭQ��bm�Q��`̨�[,��*盯ha[7x s�5��gvʧ׸ލP��`w;j�5`T�l=�I{m�]G
����A����1l��t�j�� �S�������K�i���G�ǥ R��`t �Q�V�: ^{���M {޸i@!��>���ϩV��n�QX�� .BJ�������5��Vŕ����ֻ�l�=Y�ܳ�s�/'{���#Mf�9�vҦw�=�Fk�}Wu/f��޵[c���^��oOG�FCخ�T�Wo.�޷G���[���a��ם�u���;gJ�Z���k�l)�����ۖ�S�}wy]\gJu�{���uu����u�^���N���k��W^׷�������s��۽�sۺz�����ɵ��{�kY�m�[�:nvWlH����}}�ζ>�;��]=��{�{�Uz���m�k��������܎����kaz׻��ױ�Ok{g������;����˴T�2̯l�Ն�w�{�{�^��۝�xw�=��j�ɺ�wm���^����ޮѕ��ݶr��xW��h�qs��u���V��on�n�n꭭v�܌����Ykn� ��Y��Zu��n���V��9��.q{{׵λj[v;^�޶��s^�{����ڹ9[t�z��w��\����{�u�-��Y�����l�˫�lPπ �W��mW}ۗ7��O&����c�E<��ݱ�k�3n�;vvWq�=6�Z`�몽�:z�ۯ-�n�"ZK�U���퉛Y Fx�}�t1G����J׻�t$f���֮���)����+�u��;�ufOr^�|      ���R�5G�a�  ���%MF ����L�i� )��JS�L� &C&L & 4�S����%4i� F��2b0 ��&5UT�@       �$IL�4�z���6��F��hxFj>o�}�W��>�����Y�=k��>�:�&k\w�ֹ�_J(����]&� �������@ �@M
m�q�7��}����o����̓�?�BT����QDI0���U=�4��+��d�*"q	�~�>��}��#�~������ӰTQ��_:4�h5���0$���?f��L~%�c�É�$5��o���;?-��9�nmpi��_�{�i۫5��n��7*�z���[G2�-�n]�6���ݸ�F��i�V��m�R)�v�Y�a�wU�� Dd6���yi]�e#L�sh�-��\WCܲ��om�U��v�v���AQ8����b�"��&�%;�[�Iv��xQ1-�˘��3������B(Z����M�C�/A����ս͑�W[sP&�
�������H��H�b�;ݴ}J���&�Lս7}eu�AO1�6Sk�C�Hu�]b�f꥘S%^ԭ��AV�D�V�3Tʌ�*��W��VzY٥�-5��E�W{YQClM�2e@��S�y*R��p����mڤ1�̶kV��\����/��b���8lAQA"�[�D*��"��O@�3h�EJ��1�QR����[���i�W�^����,����.�5�FIv���[Ւ@ �t������%�Fe�O���![G>�,��lȎ�B�i�䖲�x���ŻH��;K�6��9>�r��bޒ���˂��[Ts�Z��́V�fTy��5%HZ���ed։�Cӓ-���b�F���=��P�/f��@wY�w�uj���mՊ	����V��7JȚD���`R������hm�z��ބ����1y�aYIk5y�XJ��bMY&���2e�ر ����cu�Z�Y`6����rj��:HX6��9�]� bd߱V��/7Pj6�G���6��f�#��Q���m�H�����I�e�Չ�b��T�U�I���Kj�Qچ���;�6�lf�����y�����\�xR�wz.
 3�����2�TCvԵV�嬄��ZǚI�b[�B��'�T�$ey�d�ð�.�m4.!T�0���y�qh�kdݓ����"1����p��$��.�c�:f,�i <0�Tl�$��H�:�Ur����WX��M+�7y{�%�F�
/$��aӻ5�c�6UH�����7�E�U� �/@�1V'��Wp��W�fҩ��Ak]�z)V��^�f�k0��#�&��X���7A�\M#%X�F���Y¥�h�z�n`�F���@rΉZ���c&G��܃H�9'��jXe�h�.�pkn�ɢ�2���`�6F$ƍ���y#��mš�To �3��.T4���Q;_kHQV��y3."�u��Z��gb// yY�����Gh��j�6��X ��7�7)�*7S$`�ckw�9l��v�v�δ`#i��vQ�MG賉
F�h�J �(f����1j���*?on��l�+>;���X�2�uf^�Zr�Lc�2�J�VM�v�)V;<5�`A[ָ�[��BI�x�ǲ�Y���8���Y�r�z��Bۚt5�ԭ�"y(�5qA�)醦�O��y;ZckD���L�S�+HB�4�ʁ쩛x�$`g%�l	+5yQĤ�y�{�ՙJ|r}v��D* Ӱw���4��r�[�+�Kz�������h��cn֐*eZ�$�p�x+U�K.bLak)��ދC7X����t����̢�����\�,+~��f�Պք?m����v5�2����#�R&+�Z��CF�[Ӂݪ��諳h�ʷhl�T�c�`��V�Z.U�w&�H�>X���*�ky�Յ�@�y<'P9���@ѻ̴;)u��D^h�6��������D�M���*4��l$�X�hU�7[�
:Z��@���0Ywi���kXoBnb��c�q5Β\ޑ�B5hY����ڰu��)��'d�����U^ʚ^'���D]��n�J�r7��aa��|5eq%��7�ɬ�L���kkT��zѵU2͓F�m�w����6�5�E�Ve,apK�pT��X(��qz�`"�Z�v*�=�+R9Gi�B*�ɢ(-�u&f``�@GE�f�rΫx#������4�Td[؞�-��VII�cf`.�(P��꘷]���j����q$(^��jʫO 6��Zw����ƹt�6��^�&��g�h8/4�7]���N*�A��هw*�	WF�E��ͧ��@ێ�D0��jh�C�͌ô�1��WF�5�U�3Sz�#R�UÔ��K֔�e�̐�f�$�E�xe=GB�N��d��0Z�y�*��lF���X]����H����5�vFɣ��Yix�c��iP7.�h2������9u��S��w^�b�&�ک1(^L�ї�w,����V�֘;q���.5��u���&Vj�����n���V�p-"'�^����A=�M;z3⳸"��y�F�U�J*�5S:����L�A��n� ��%X�[��-�V˹��
�t�=+[��he`��z��t�3h��Vbcn5f��Q��˻ߓ�i4&h��ti��;v�����m�CD����7plRnh�+f�7S����� ��N��w.`�駌�t�{F�miOEiK�k:4��0�/z]��خ�����l�ݭ�-raIh&���4G&t�;��Ck0�u��s�G)�I`,�����y�@���e��=�%�!+� �ɣkC���aH����ܨ$�%�V�y2<��fK&�M�tV�:r��֒�BTHh��E�X��i]a��^,���V����*l\Uje�Ԣ�J������TcffY�lB��V� 61��6���)�nk�V��elV�5kp$U7M��X.S�D����cM�fB����A�O���ƴ��wOꛒ諤����R��Ȓ�;��$�'Q�YV^�cb�;W|����w�.���Z��e��wl�z��xo-Drն�U���j!�/6�enb�l�-��c�:��WH���&ݑt�{ �Vؼ"�Z�c�������g�[�E N.�/3���mŷ�m�<B�B+���L�i[�����[^Y�K�icA/��v�H-��E�'i�}x����8���淬��t:���{�,���<�v�
']�>�٤��Gp��t�<�dzV�ʏ��sHk���E-�z���j�U�M	c5��u���5]�'v'�en��f
TKׂ����q<Y�gh�m3�Zu�ʽK
5�q�W$w]�KHĻ��Ks]v�W�`ͫk71W6�1&��%�tݥ1b���k�^VQ�uhb�bTT���7e؈ltp��X���@,Aϱ<	B�Pam�ĕ��[4���ki����7��-f5 �F�Ԉ�J��*
�F%�̓0j�e�� �y��3I��QI�1�5�
��6]*�����I�5k,��F�f�ŒN}ʙO�Ue4)]r�Wr9Wz���K6f$(�f�vt*{	�/K����[ EV��Q�7�]�a^�y�mɲ�ڽк�'(���	a�mu�K��o��®�X�Z(�-�4�u���B�����w���ɩ�����9�)2�
��k�h�2fB���*�m-y�NcF���Rb�&ɥu)m�z�
{�X�K`֌`5������;�q��VU��H�AS:m]E��fB�Z^���ص�h��6�	'%� n�2M�.�+U��K�P)
6��S�*ɥ@���(��*�ꛗ�5�*���OM��t�ߙ9v�B2H�E,ɆX������R	i�Ix*�_M���Ӣ�:�e��P��/U��re%��M���Lॕ.�n����hU�Gp���V�Vs�s�&�qe�j��X�]s-n�ĕ��r�b��Q�����2իK��Xv*�}�aT�v�e�7De�+^�*�G��I*�,P�.n�͍ջv�yH����w�sv� j��I�v�cG6�tu��4J���.BΞ�h�ݢC\-j��v�U�*�^�#V��aMn�XX1e3Y����� �B� 6�M@榶�BAG�;�Vnێ�U�ԏu��F�R�Qz5K��]ȝز�z��j���;����q������7kokŖ�����@ذ�����ʍ&4�h^ ^�]n6�T��
�˄Z���ԦVR@1W��b���V�קNW��h���1@�4Ф��CE�P9����Q�.R�V��&�a�S7��f�U����?��8�(�ʔaH�[�Ӫ���é5r�y��T����Ÿ Ugw%h(��fk�'��&��(��[���72���Z�j�=�V76��E�؎�RB`�1��@��l�T
B��9�
�����6�N�FT���ڼZJ�UtAZ�"�8���ݒh� �e^)<r�ą�b,�b�޼�:��v_0wqXF��\^:Ie
w�j,v��pUL�F�T��n�]�9�g���o.ݼ(�%"��Hi9��t���kc�H��t5���A�)��-�)��y)�b�,��pjє�H��bRm��a�F��i*�dq�8�<�ɻ�ނV/����ݺ;�Pyiyh�oIʘc�wf�D.>�7�k����6����zA-M+�ר{f��!�n�^��nf�&�I��i��vZ�T�e�cn��ҔF��B����t��N���^�cҳ<ɑ����x*"{	�g�?~c����g�}�u��)��`��?������b}W���=��3h#����Q�@                                                                                                                                                        �                           �I/2��1l���ю������شn�9A�u@&,���eAjVt�`��.�x������0m��6�"|�,}ܩ�ܴ\4�,��2h�Y�0�F����w˄S*�k(�M�4��[�\���5W6�R����j��ǲ��!{=^i��{���7 t�)Y�gll���SS�a�6�Ey�ܢ���� 8lWRK�)��*'#���[ЧƂ��K$u|:T��4\������Yw�-�,pJ>)�|@ �1���N�G"t�߱L���0�B��|q)j����n-��s3@=�q�î��si�(u�$��`���ٶܒ��3�=���W!S���g�r�}�L
���ō�����S��B�G�x%���gu�<KIW<�q1W����t����L��������{��lx�vK׋��YA<� sC�O�R(�e)�X�ޚ�k�ypHU.�a"n�r,��7�1����t���mC H�2f��v��Z�Pi�w�U��6��$r�v��X-Q�<9W�r��u:un�Nu�Ĩ�_I5���u�D/w��&�Kt�1�
�8�6OTz���ݦ��m���ɱ�"��E0�{J����-#��4�6摺q]>���<V����՝t����=����+D�[�,�+UK��bZ��èS�)XGe�`7�^�r�;�w���i[0rӒ�T��	i�^�4+·�5q��Ӌ�v�8��;�.�����1��f^�U���'MQ��-n��>�Rڄ�&�K��՝��h�I�2��Y�lC��B�-j8I���s�j�Z�ɠ�Y\D��if�h�����m��~����ƞ�(V�������9�;���a�ջ��Bg���:�Xn�5� .��}X��Ӂ;|����D�|��p�/qh���B�n�VMޖp���rr��Ryw��l����P{k>����r�k0a����yGL����qjV%���|C.�����$�#b�IP���׵}��$n㩩n�G`Ϋ�}w�#]���%@�O�.�C5ζ*�kv�[S4�ԫ�����hYy��|����D���ՆWִZ
��r�:�<�G�j�rN�gQ�Li�Qm�\��2�+���ۈ��Y.�K��P�]�����K���D����T�li��3�hO�Z��m�#p�"m���kQ�֠9yҴgE�{h! 
����!vD��,��[dQ�E+���kI�l�yV��(k��L��٥��Y�o,�C%a���ԕ�Z�-6�vDr�S�4�ΘZKr��mI]F��e�n�1�ŝ�V���=��ң�o;��7*@r<�pI�ݎlT��r��D�z2�|���杠.���n8�m��;�M[yB�[�]�[	ٳ�.;tĻo@nm��r�7��o�]r9+�*�Ba��,_(�����:�*�˜�Aq��h�shPŭ^:��2��фX\ō�+.�o7D����q�`>��ˬ��.Ժ9�c�h:U|�y ���t#T7 5/�Y2N��t�*Q�a���,��q��ͤ�K��`�r9�"��w�����R�0m�|�����w=�)F�Ӛ����b�Y5>�!j��q�p��XVT�]V�36����+�Pq�BH��޾��V�U��u�4m5wx-ô�Q�}���փ����/a�s���r��^�8�+y.�P��̔�UIu��sYa�Հ�t�7� �����5�l�0_�4��Lezm���/������z�hq�/i��塕�!׹n�hX�|q�r�@ZHg׎*7��pc]ܞWc/@q��J%eE׀�=ܱ]�]���6�mL�K
zJ^�n�j9zq긥[�b�+6����-�]����r
m�R��r�Y��Q���Q�F��5e���Y�ʰ�`��p蔬Yz���]���q�;B���n�@��"�Z,^��^�Q�԰��筝]Zl�{ad6��ĕ��n�;�vp1��F,^�����B�}���!��E�>�.񘌬0mt<��nrw����7�����.&��h����+�kdt�j���GBN���P4�9B�9���K�������Ӯ�Jծ�u��O�Ͳg��G�sxN8��2�h]�=�,�]r>�D�"��� ���ZɝL�!m�n3�fLR#�wk�#�Ί�ý`*ۜ�y�ErFH�yu�{5���L�F��,ڛKQ�2�i��S�
�]�R�`S�\���h5�"Z�Wc��-�:�d��f9�=��ܭ�v�����hdj�諠i����
ҬT��e����ˏyc;+�sa�3k�4
�d���Y&m�٣N�F��mV�$�Z�w�bqՂ��>��Ԃ�S��f�,B�5��J}>��i�@T���f\݅�S�Xg(�Q���c��P��^�[�/O 鍣��t;��Âb�ķb���J�j��]Ԏ��o�uu���D�;�1Ң��8�$䄫o1�&���9Xs/�Դ�&*��d����A�6�Z�hU��R̊�F�0�� bn;p�k����ec�L����3c�q���
��y}5�(�*T�]�L�.��G�[ .�p�͍�H1	Kw�hP���������6Q/�ڻ�Z7bI���^�rɖ�5�)o^�+��I��A��� ׻t�ZJy]L@�[q��j���ɴ�zm"�����H;v�·)�Si^����՝K��V8��Q��NZ���]E��tC���W5����0@�GP�b��*�
�)�i^���y���ڈ�cn���X�������.;<{k��8�Y�{q��+�\�i�X_)
o�'�e�����'6��ϖo�eB�sq�b�|���q����mQQ-�Rŧ��u$��a��:��|E�ә� V'�m�8�^�J��$�S��>�{�t���1j�Z�r�`�������{)�x�m0k,%0�3��µ�,_x{��IS�q!�̫�s��;�Z�0P,ɋ����(��F�C�Nbt�.팅�
��bqK$�I��Vp��wN�s3�E�x+5d,�-li�V��Pe����6u�B�7]k�3!���2�F��hs"� k��-l�6�i6�m�N��D�U�p6�H�R���8�ǐ���#�v�y�
�b����)�Н������ۻ���U���-$����4�쭻�5E�M��E3Y-�lM/oE-���<)�.i8H�_��-I�2�o�T���q�������հ��S���������S���srx�(�[@ʔ�@Z#��+�j�S�t����IסM�ص���챐U����J�8]���a���9
5�;���Ѽ�Z��I���R�5�œ-�}�򱯓�z(��x�x�A��1��5��b����PH���h\\*�jG����Ӝ�Lj�^a��y����RO���oF�6nɝ�+G	mi�g������QR����yfe,�A�ý^�C"�la���;,����'�]F��)�uי*��ie+�ܺ�Ĭ=Z1�#؎��NE���l�xh�[�W��ͦ�f. ��]��hP �:�8��!�պ}"�A=\��9�UڮCt..��Yl�2��
`���!�����Ü0�Cˢ��"�!F�Q����v�s�nЍoU��jUi�}�@��^�7Y�Gĸ�:��#���PU�t��L���,̥0�L�5�Q�QTx�,]t_\TB�67�*��Zໞ�k@ݎ+�(Q%�O���ջ>��=B�D�Զb��h�w�t٠'kN��K�����`.�R�n�h���&l��2����=�_�-P.+��z�:���6WdhG��.���j��.�จPG%ׯ�^���QC}��QT̍����n.W�B�PdKC�Ӗt+/W[x!
v#��N�@���C�fbw$G\�r���7*Zy7e#QLIGl\]Т��;�":�^[D��u!Qv�\B�;�-����/���oQ����,�ø������Z)�R����-���'(�u:T�T/0cN���;=�0	4��Kl�[���dSo���=;(#X�p�Ow�TN o.�չh�W8�:Vo�����׊�O^�<j�
bRw�V��#̝�WF�\�K+Z�k(�uo)P��������s]�0Ik�\q�R�l�%�Wt���̩{��^:��u1��� �nG*���t��JR�}CU�J�f�JǼ�X�&�u�l�F4�Xk%��'G����j���R� -��viX��z�x�SAU�3�m)�+>�E����bn��orf(��Nv�7��Jf��#]� /����`��z&$�5˖��,�����KA�8b��h�	��aV�{�Dʝ��������	����d����7�S ��������B�^� @�`���!aך�.��A|���vJ!�����0� �ǲ�{b����    � ��           ��������j��gz������?G�QDM|$q���q@��4��j���/���]�F���+�4>�7H��j�����j�ƅr��U��=�F��,�nf�lI�6�9Wv� y�y�n=y��0L1�@�	�8J� ���b�{�R�;i�7TA�N�!�ݓLV,K��pVғ�y�6v�T3�nք�=����T�n�WK�0՝k��n�<l���Ge�;���A�cX�Jb���b�����է��-��,��BX�ν�N�M\V��t��֓C����0�pЇ|45�N��Rn�R�>�b�v^ØAW��N�9��5��MVR˩)TJ�e�s8�b^���¢��M�ʜ���W�j��n�m�����F� 7o:��zɺ3wd���`9�>�r��[՗�O�vv��d,p,d�l����Yt�|9"l��(sY�T� �kV�ެ�W�ۛGU�f�$�{W�|�HطZK�o�$&�Q�'5�3b9�����-\L��ҐՀ�^��Ր>"���u�YQE�8�۟�p8�R��+�����K��DY��/*Ei�:�ڥl�����P��	��س�y+	1m������jXj"d�}�Am�8�9�bJ���p���S)��w&g8m`C,,��)���(����m��ݲ�#B*yxd�..�a�qYcw�����\F��ǎ�n]�ID��^�h&�ɵr�͎�v�a��i�Q���V�=��B%�$���g�%��T���t�L����*�4�T��@�L-��/��" 7p���b�[٩i��c��/�	���Ӭ���K�b�������s7)�X*Y*���`hw�˦��Cy�n�;R���F�\�R�%��=Cu$�{�Mb�-41fm03G2hF󈎞	���C{�Z�E�1Ee��,}��ջr���nM<5�	���E0YXpV��*Y]v����@�%��zʦ��wk�m���ZbDq)�z@����[YkNV�n8V����K�:�K��)ә��5LP�^H�R��0��|��D�)7º���Hޠ�Wx�GJ��cE�qi��(�s�,��y�Bx�߉��:k�^`,���nmZ��mU�k�Q��;��_SF:�+��w�X����YńU�z:�# ゲ��@]�%�2�����tR�e/����)g\��wOq|�f,�7�J
�y��f���2��WJ��9p��CI�E���/���՝Yo#�����6�u�)5|G^�Gl0層��`Q���uɱ�eu�jH�����|�b�]!�s�`�@p��k�n�Ʈ�b�Zw�t����Q�.�|�ު ��QL�r=�5m��f�B�ֺۨ6�c�A����V��
�/Gl:6�-,�] +(�,ӡ��T�0� Ӆ\�t�u���.��̭t�R�9��C`�W+f�3�`S*��1sLwn6p���3;���>|�^�F��̷֕�t����o�UeBT�}I2m�u0־�F���m;j�}F�n�o��Ȋ�]�s���U�Vn��f�x	�Q�����c ����b���4���Y��������8��N�]AM���H��2�W�Rp`m��x�KI��g�Հ/U�R�+T��6�BtZ�%��:�b� y��0���5�F���Ŋv�e���$�1Τ���@L�c/inV�W�`�@�-����tz,Lk�s	�U���xb��iP���?�����	�ƥ����@���h�m��RЃ�38�ڎ+�n�E�VV�C��Ė�G3l���"�X���x^�[��:��?7Pit�U�q�v%nr������Y�oK��Ӓ┢β�3�QN-Wv+��`�5��KR��r9�����9!�fݭ�ՙV�7�V:��F�h�N:�|ER��&v\ifD��ȍ䗛��v�i��"k�]S �=y��,�����n����� 3h�i�*{��G�u5�U̝y�*�p��E�J9�8�\�zJ�Q[���z�R�<�h�0
+c���}Ke���oS����2uR5�uՇ�fj��r�]X}C�gthVj�V��/�j�Wg��z�}�$6B8�
�AT<7�a-��b�WI�v�f��J�6�Nr�T2�mn����f��ˬ��ԃT5:�ٸ���a�f��μ]�#y2r�V��Rc�Xp%�+�osĨ;�[�[H��$��u��d})�	�.*P�����!��e�l=��6�^��1
Xu1�ht@ԝ%�bVbE�%�cԝLZ��䤺��wY�s3�b�*��.3*��S6N�\��\���Ϡ�^�RÆ��n�tu�V4z�T���C/�����҂
š�C,��4S�|���P֜�`]��yW�f"S�F�9B�s��ً3��g�Mu�oX�N�k���.U���Zؖ��}άt�k�,�uv��"��K��hx��)���
_t%5���%�*y�â�F�30�hGX�����ju�:Q��W=,��вV1���ɉ����k_J�W��T��I���^��:�g2��+���~y`��pf�gJ#���,�Љ�-�(!q&��j���OTc���B�b�F]�<�cf�<L�Q^�휙x�Yy"�(s/s�T��E	Ϙ�MV���!�m�騰J,sWv.�Y��Oga�e�'�c���/�j��B�F�uO�@����
��5C�aі5�j�I����w`D5b�D�wa[�Mͬ};^�n��c��"�n�5}H�j���{0�҂7���+TrE���-]��&-Ok�.qv�vn-�6����Q�-:U��9�u�7�(vW������Kv �ړ�.N<�/Mgwv�A�L�G<�Y����bl�`�ʑ�o�s7\�%u�
;Z�B�)^=��2��Oc�D}{�e���P����i��*��Q�\#t����D��>x(�,�v��X�̨m,�7O���q/�,ۧ[�>�xL����:��G*U�p|�������Z���������<$;����/����.P{|�)wn6��Ȕ�jb|t=�z:%J��Z�)�j��k3��ZQ\����1�g�VR��2Ӿ�+뼔�k�5�.ұ�cvk7�i��5z��ò�IA��^K�Mb+�fh��f�E��uX[QmdӇʖ�^� j=�[��)����:J�7^:<Vy��!i��#�y]�.�P(�{,�$Τ!if��y��V�' �i�8�2^��ǯ������`툔MB���Q�)'i�����2ٺ9K3V�)�1Ѵ���M>��,�3���U�"�i�trP��^�)����ӡ+du�������vu,��X�˫�A"b:�Y�j���j�Ve���&��ؼ��0��.�
P��&�4�ͥ�RVi���s�e%�4��K�����w��i͈J��X0��gR�k)
Ob=\��zgC,fMI[�����p�}�.�'t�A�<4	,�WkӦt^��Zܤ�[��i\4��x�TڶO`�x�+�q�]�Ik
m��V�6�rx�Y��վ�����VM��4Jh>�5�`��_6�7ԩeR�۟_tuu�5X7��bYG_��Yl�#�LK^ ���J��] -GBJ0]�(�*���]l�W��;/�-Y���Ҳp��_[m\3n�d�nH�R�j�Mܪ���f�
�	P�h��&h���ރ��>y$��]*<��|���e��l)򚊒n�.�4H9V��m]lb�
]�"�$�is6�9�̜�Y(��tJ�����4`�ّ`���K�hpt�u⭮�}	����2��d�C#�*h���M�g�_f�lKm^RՅz�Ck�7mtB���rK�X<��շh+��p[��TEd%��s�_���M�K�ernsU��b���,��	n�Z�e�V|��j��GL��)16чL;ǳ�-9w��6��Y�/4n�Mϲ��f�����7��Z�]6��O��PL���v����K��l"�M�'�;7�R���r����`�R�vB�V�K�u�,����O%��u�����މg��r^`_,��uxY�14#E�[E�h�yb��c�fS�fc�r�5-˒��4nb��d�1�r��B0��M1�atOf7k�wP���n����m`$t��gi�wV�p��������;U,����]F�sT��H�}��i-U��:$��1l��|:��p7��EX9���ը��
�hd7����5�!�o�g$�����W	��F�&���2U��9�+E�v2��r������_���`]��&�GH��i�Ú�V���Z2��d��6бh'�u^��(�72�	MYj�g#e⤆��G��Uգl�ʃ�!��OB�*͚�V�ߥ��fP�|�u���ꬻ
;/�:��0h�ˣ\�a����@�V6�!��(k,�:�^ʴ��N5�6��`��s ٣�bK���Ӹ��+ҟqH�W���R�u͊tC���S4nC$Xn͎���ٹ�]���rݛ�eY�}��6�tэ뻨o�@uz3j�p�fiߜ�'@iETc��VƱvU;k���l�{�S-�y��m�w�u���<�o�?%Q�j�Hn�(D���;U9>�EL{�~���?�               �ݟwG*S�.��*�
ט%aºn��f6V6�vh>Ù:����q�
܉P����MC�݉d�:L�ҁr��ٻm��}&����}�4�w:�$�hu�]
��;�g��oG#��\�� �6;I%IaP��V�M�����{E��UKx)�,w\�m�S��*�iޜq�[��1�
\���mW���ݕsJ�x�<�b����k#ɭ���j�:�f*�u����6��V�b6��a�L���>лhm�[�F�c8�*=z)�94�.Y]ILn��gmqέU��N����}��h!-v3K�q^�}[ݵ�L�%�Ua���.�����n�~��*fe� 癩j,�5xo(���JT:��x3o�[�aܤqd\��;��t��C�+U�]#��`�컏_C�C��1���7�u㨦�f!r�.�Rl
��dW
�#�@� I	#�~�a�^��Ʈ�!�ʝ� )
��B��JG �ZB�8 0��� � �!������/,�j{�7�Ȣ�{�2((ucYQAHQL�U&FMPUQE&ف�&�0�"� ȈJS�sX94�a;f�L�j�BP�W6QTU)M�j�̌s,F�*�Rꥊ�J���J)hZX9�d�I�!�P�L��cV��}e�M.�!)
�$�,��#��IKݑK2dCH�%!��HVG�鉟��C�{��3���[����Еfڊ���B^����s��sGDiv��6�oF�o��KN3��'��?��Ɂz<��ۡT~,��sW�.�-
d���D��X~�ؑ͑^�3F���|�7�ԓ�˞K@�i����{����AD�z}~�i��+�d���+ޚ�߭L��<�@V���[F���)�}���&א*�5y�|��� ~5ϯY319�ܘ�C\��t��h��}+7׾GC󺉲���2Ak�6>\��O��}Xt'�5sف��5YM��yN77�ַ��c{W�q����ǎ��廩M��8�u,n�yRu�αj��E��%��]��&^L��mD�n��d\F'9�y.n�i~��y��A�}_��o%���f�t÷ۯV���4�Q��h�Xf��vQ`�ី=�<�w��Z�E&:��|�h�{�;��2��](u�$\٫�j�syᕐ�3A��)��eaM��b��C4���:�(s|��c�s��ɟ��92턵۟����	8�.�_���� �������JN&�[u�K]!i������OU��W+���c3wםqA˂/N}��b�?9���_rG������ '����)�{mr���G��{K��K�:rQ���Y����E������;ދO��]��D;,�n�ކ���,�wuo�7���P๞%dIή�o�����MeL����l7��
�՞�����������z��O����=h����W��^���/G��蕈����γR�;��Av�b�ƢƆu�� դo{q��k����i�\:9b�4c�o;�Jv�U";��Q��s;���P�K[�/�MV��e��ba��Un�\�4�疛W�ÓJ�y���{���	�[�f`���|��lpf�wZ��}�{܂�Ғ��a��^U��]�R�^��9��uW��^w�S�dvN?h�泄���n则^�V�
�Snh~���4�]T��Wq{X�𷇼l�K����t���e�{UiKW�XVs�w4�����i�vmvJ,�*��a;b�[Y{�k�*�~��'Z���W�@�ʺ��o�޾fU8�O9�uށҔ�i��u�:Ū�7Z��qw���	�+ح�i�������m����;}��̣YWQZoj
����S*��`�9mX�}٪�xf�h��[�;v��%�6FZܜ	�}�V��J�� ���&�̲f���Sq�������,KfR�U˷o�Vn��k�{���j�T��LIɔ��;*��	{S�Pz�1�p��;fD�BK�*��g#aޓ�{�s�;�7�.ָ�������c�.�ڒ��H-�w�S��e�ԕ�˜nw�ܥ��iH��x	�rc���o��0O�;{S[W��y�k�l]��QY>�B|��W���<Y�X�ay�F<��e<W4���5pW>��=��뽅EE�*ߢVM`6��l���
�ɜV�.z�|���e��~������]����h��o�y�':�B����R����d����N��2�җ�P����8�[�6'���Dl�[�ia��:�����N��4��M�*�st+�|n*�����옵R<�y����<=�_qrtt��32m�zNwN)��^&��R�4o�í��[����:[},�:��˦�yq���A����M�6�یR�:3��Vġ�{�^ȉ}w��~�>�f���}���㽦�X{�]��k����y��~�ßPC���j��R׋n�9�q��얲{�b3)�K�ϰ{q�]x��=.��K��B����0;#�c{S�܇[�2��A}�X�̊5����H�]ߦ�3}(��=��d�73�u���;��%�t;��]oW�Ob��l8���ӵ/�2Y8An �n�^�����QZ����K�g5r������LQ��*�V���b=
<�+��E��$ҲDU�z�i��Q���ڷ��w�F�}1"s�RN�*��v�[RH[�ً�I$wGD��o�{Q	{S��1ea}	�dH�S�bq�c�S[��k������oc��	���V]ʩ��7��[���b���ב^T`��Bu��8yU]�L�{5'y�7~�[>��G�oլ�NoZ�9�/�/_,�\�w�{6�^̞����C��c֫���i�-�M�z��.�u�VU��:�"骋����]�a�w��u*X���n�R�����&+��E�r��s��F�Ԕ��K���ÙX,C��2�z1�Zum��z4������'3����}ͿmK�3��?��D`��3�<N�*�zE(������n��>��u.r��j�i������	-�!ʨ�f;�wN/_V��xop\[���9.�v;��T��qrcq9<ғ9o��e�v�����T��l^�̺U�xQթv���kg�y2�.g�Ps�(�__At��5��ڄ�=�u�2.Ox�Y%t;�ɮ��q���>U�6<�8�u���A���������|b[�Kn�������[(3�����:	�r-�VO(ez���w<�w�#o"���m�P�Trse���G2#�&��7v��N�qc�w����
���Jg6��sLw��ũ�[���w�1ϫݳ�{�	�`�<�2�R���NxjhWzm���W�7Ltt䛱L�%��e��-l}c���AN��X���+O�=9=��>V�mIC;:�����.�1`��qt�M�B ��mx�i1_�#\p����8��p��.�A�-��ĥf0�5ӴM��ԑ��^��1%�Y�Y���s���I�\s���%����Ns����۫T6]ˀ��\����|����V^ �h����fK�y��Q}P:��Zj��]��i��ۀw|��}�����dY��K�{/h�NA�tL2�2����^�Ntf�g����eD�ɾ��Bç3�j����AP�3�j���:sb�u푽�D��z=��ʛo���Nse(�U��;�T�Q�U�Oy� ҉�j��v�3�"���a��ͮ�`���޳����ŧZ�3v[#���d�}�(��wC_���M�zp��7��7�-�աzp'p;Z%�"�G;E�(e^v6î�;"ֽ��%ju身lK�nE�5vc<�\����XwZ��ngb �zr���t��^��m�T�6D�J������>;��>]�}�+86��Տ��:�jz�{�<���%[����Pg�ޝ�ݚѯ_ݨ��Q��!�vy��u/m��.G���j�լ�������p�u�N9fU��|p����&��*�P�����������{�#�Vw8�����HW�t�����o�|6��z{�/&���d��n��
f��, ON���Ի�o.��5����A��y�&��`Xn)=�{�|��W9�z�5�D׮<�~�3����o���*/0[7�'����s^��۱����PU�j�eb Z|m٨t��R<����QJ�>C�o39���ut !�9�Ŗ���n[�*�p�À��S��Gҕ���|�r�OT�d��������2-���@֭��X��ԭ÷�3q��^zW��}l���2ܖ�bZ��1h��T˝�=�`9�l��{����i[���f��QQ͹�N��M��M�>6]s����?]n_���i<nL������,���H�U��KD�s:�ט���7|C1^udg{�R��n��sӭ�<���{�7�o$�|�b�w�/w���/Ӝw�:�����8V÷�7J*�)q噃/�5����fOSʩҙ�s�Z��.���� �X�g���aq����@�?�γ��n�<?�B�~��*�`Hv�x��F��cXژ�9�3DǠj���K�rح��-i�e��`�������֊Bp1о�{%!�#��朋0���ԅ�8嵶�4�w'ߢW՗���kZ�&��֜�8� ��3�*�B�KM�i��4�r�]Y���9�u��P7eJ���*ȶ�T%�Qqvn�4�yM)��
���ˈR�Ҙ��)Rr�`�P�Ck6��h
�wR��"BCQW�����z)����wjo�!KF�\h�+�4=TAU��AR^dt�%��:���e;62�dXPM=2�iQwm�$l4�Q{&ֻ�/�&��V8���;��&u�{�sՕc��	�h@���â�.o2�;p����]���%��[z�Y
�``m.�軝d&6�����.��	uor�3�7+���B��e�Z�ÐҺ)ȃ�Q�}�%eu���.CU.�b��Xi��n�u���cpu~���	k����Q�e��j���f��Biܸ��"�ӧz8�Kz9���)޺��+����^������               ��޾�K�/��q�X��)ho4tVT1���S�N�f��()N���Sz�N4v����gAG
骇g�VR�l���M�&�u�P�N� =�`WE� S��+ȯ�]1������hB78�X����$*�mZ҇�F��z�1��L3(�Y�W�����`��0�)��!m�	��{K���Xķ<�P �9��3b&��#4��yw&�L�ێ��5`F؏�-������i`�̲�]��h�m[A������6no�N��m��f�����{k)H��C�ɣ�=97�7�>��w����.K[��Y�[�Z�X�S��$6ؠ��v2�b����b���F�;2N��W��
�|����pBf�$��T�a$:ȭP�����j�y��;�f	�սu,��R��g�A���=���60D��zWF��Q$y  $��������ER�IE)W�m�F�("�������(h�MCk���2Z�i)D��r�(J

�dd-B�eITd&@����H�fb���4�CJ�P�N�#S!J���PP�!M��IE SK@Āq�U��@P��-%)q��̆E!B�$B{BR���
R�	u�o�v;����#�xu����-r���\N���fvK�	���y6ΣR�W\'7�"����z���ُ�:��%;y<����yN��HZ~cj��F������;��<�����a�3W����]��߯Ng�e}��+S��G�ے���^δ�+��z���5{�0�n�!�ǚ�C�V[�`���н�{�ܖB{!n9���k����v�� �c�����ELb��\��ȓdo�e�\��Nuu?W���ͽ�]�|�u�h�3�F�ҨW'C����������ù7������fǇ�^Ԗf���\GR�t�f��=K��Ĕ��[^Wej�hT'���w=*2��yV���^�q����!�͝ˊ��V���et���^)K�|,�Mӵ�N^�ES��L8ָ�c5�?��~��q��W�x��1�m��%���[���D-ژ��ת=56��G#�58Ԙ����X��K�������_��R�2/U��Ҡ�Y��u��U�yz+�����}�6�\T�h���������&��u�{��=.���f^�sG�ѣ.1o���Z�#�ۃ��(�����ظ��&{ܟ��N��_���w��=�����[�E*�r/���?U����د�5�{������
5�[��m��g�z�5�ꈕ�����;�~��Y�`�R��D�~����[�?���'���:�Yz�r2���N�������ԭ]WZ�ޟ�([���J�KY��}�C�No��_��B�>U3�S��+����~���������dyqZ^ĐR��0f�J��`\��������`�B5��*9:�T㱌�w�iw*�*�I|����\>�]�4K[���G�}G���wk_e~��^�=p�̉΄�䶡U+�ɫƌ� ����u�#ޫj�yH������L�ܬ��mU�=�Ӧ��Z=U���E���>��mo�W�LU��'�����r�~���!�<��h�M�^�f�����K��3ko���"��}�o��qd=���Lͧ���a����Zo]�Ԕ�SW9�y���g���!���ETs2Ї�~)��@�N����F�m�>������Ɋ{��a�� uׇ�ԟ�~�D_IOމ\�"��O�Ч���M%Tr{���	j㷽ђӁ_����������R'F�1��`+�L�ln�U��Lj>�r����cE�5������;�j�I��C��͋L�Ս�μ���i�(X��D�$TQgыp��Y�5(��?�W���:,C}}��7��_uj���~�מ�oZM���z�J���޵"٭��.I�;���k={y.m�ES�ua�앿b+�%^�]s���^9��d;�pq~�S�J�����#ٛ��z �E��+n�s��G���B����������{go���:2�|\+eL�uJ�Z�U���g��"������~Pﻍ����K��u���|C%[���=Jkl�!���=��Ǿ{�u޻ߏz�P��Sӌ��׸=��q���	׺�}��|Й2�y���]��K��oօ�B��][��sɿnN���[���~�����[K��]|���5��.�yǸ>��r��~��a�r %��mq��a��}���?�l
K�ڢ������_�T�J�>��{�l8������:���`�}�7���|���4������ĺ����β�����8�}[l�;:��@�ol��3_�3E7}v�+�tΗSk2�Ѡ�^���w��O4�#&��w'Wm;	I��h���<N���Pш�����H��������ߏ:��m�u
uVH�`��k1�W�����5)Ի{��K���pw>ƥw���_!y�ك?6���|6_�FO�t�����g��&�]��`�d������ǸB�>�J�nt����`=���m�����߿UU��x��4,��_����OǾ�̽\H��z;��]���/�k8������S��Cc1�<�`<����}���㞼��7ۯy��=���#�C�=;�˘^�����,W˙y;��V�G�J� ��!LC��&`�����0u�����'��ri�m ywr�!��ܾ�ħr�&��ġ�X�2;qh�{���8�m#�&�bҝI���Ѷ����y��5���G��^a�6w��6�������Kܾ�̩ˬ���w6�;�����y.�bP�:��/;�z۟wߎ��m����K��/p�<0^��6w��W��%��S����8��G�ˉ!�|�R��;
U�S_������c'�~��DP�Й̴��K���z���Fyv���^�g|S�a�w0nW��'��~�qN;=��~�;���똃�z�H�0y/�x��{b��aܙ/q��k�^���{���Ol�9v�+yNs�y�Þ}�=���<8�:��x�䌑��1Jy=u�w��� y�o���]u�I��!K�K��s�*~����6�V�|{���s9y��*��֥��0�jGK]i��Vs��-A��m��7&'��S�3=�@��c!Ŗ�lꂓ�ѫSF�y�Xs�����J�ݕ����jv�7��9�~��=�r�.�|w�W��� (�Oe�W~1�'p�sޒ��|��<�!�X��{�.J�m�/���瑜y��q�^u���yԧ���om�!��)��y+��h�+y��N}�;���;��	���o��#�J�~�ފ�V���67W����|K�y���Oev����|��d{����iM�v��8��\�c�|����{/��{�g�m��Xu�k�9�3���ݸ�^��|\������B������]�qH��⚔�c}�I�{ o9���ɶ��o�߿{�o%�2S�07��|����_^w�aM����^�o1�d6��=��pN�v�!;��]��_ ����;�ظ���ν�oT:�ް�v��ì:����Gr�/�0�!�/=�|��|�4m�o>�Sԯ���y�;��nx�~u��ל��Bqħr�>���lu�s�!�{/��=��B�/��{���[h_d6���v��u!(O�ݮ}�򷯙k���U^��K��u�������`�'��<���X��+ܝGr�q#�8��0��/p�U���E}��gy����[hy��6c��}���ຐ��^��x6��@��N��2Cx{��|�yN����0������f���\��g�d���>��GУ�ݴ��'�P����FJ�f�<��z�Oe�S�0;��}����S�m�0�ï;�N���G�k����4�m�Qۻe�{ɻ���٪��+��y���	�V���­���]��z$����;�*א�hR��q��ݦi?Z�����ѐ�0���e�iL��:뿐��@)k�ߎ��;���_���'�w���5��T��>A��C���r�h�y���|�h��}�����}����{�����s�>���j��_aԇ�=����w��C�;�)�=��/�Rw/qΌF�
L�P�����"�}�6����s���U�z��������u�{���H�w� j^:���6:�K��s�r_c%���^��x�G=�m����������v�C�N�5�	[�k|{����8����6��'��]h��]�7�R�z����-���nl��5�v�=s�~�߽Ò�!�>�Ծ�F�؏R��/�w	[��o���� �W�2D��%p��}���n,U�����~E~�?}���~ڏ�.H�-/��p��=b��m��{��qO`w����7;�J1�%;��ݎ;��k��߮7�n:��s�R��w���4�I̻o�in���������cX	��m�)ܦ�y�<{�U�b��g�������S*��?~��������.����}���8;�=��v9�@˳��\� 9���C�1:���7�5G�=�Ǿ���{�m��{������N�!v��=<��(GX����w�!�_e�yx��w��K�8�/q�W!���[{�ew��w�~������!�s	չ�{&����Wy��!�rS~�e��`7�ｴ/�o�ݐ��Z�y��_�ט@"���M!�!�E�'��Yyy���'�G9���+ߟ�.����iRlg���qT�#��/ofҊ�mxOV��w���8���@{�o�\s�u�|���eT@���|�ι�G�����9ʛ���˿�0y/�o�#ܞI�y�8�e�G~��ܾK��<���|�a��~}��=ｳo�C�h��lSx�lǩ�d=��۝����Cܾ�G2=�����a���9=�\w��m���ˮ��Wˉ~:��W�5����d��`��љܯP|F�by������u���b�?}�~�t�0��;��-�ϛ����s�︇R::�Y�̽���Z�y��18��4y�w���d�ƥ�	�?W
������e����rN��������)���^����z̕�_|��x�u��9���N�;��}���O'~����՛m�=�����1:���M���^���aL���z�R�����K�4��b��L)������#⇍�������#�|�x�ъ�'��@��u/��� mq&Hw#�wyd�ǐ<+z�US�L}��*��<�K���v��Ƽ\�������t� ���7�#����{d�����O����ɬ�� {���^ch^5�{ϙ���ߜuϾ�A�����u�����C��9/.�%�ն؏p���^�����|{��M��=��ּ�~y�7�˜�[�׽yϧP'��%��}`=��m�I���\���X��o�l��y��k}�Sh2�G�7=�<���O��k�U�����j�.��(rf���`��;���^T��78��nFY�p�17,YKT�=z�p�ʓ��|���@;�)�ڸ�|�oG��zNlI�Z����篐����
H���g<q�^y߽��d��J�5)��>i(=��w��	��/�a�_$�4� y�֖�����[�0=Jw���y��(����c��������ɏ��ѓ�!Aǘ>��qK��^��C����2e�lW�{�-�|��G�t����.����?ن�_>����߰SQ���<u�q@������1ܾF@��;��>�A�̺8�\B���κ���y��9��m�мG�<�Hzf'r��0�@�7�B˼�uu��A��� q=G��ɿ�C�}����:ͽ�8��y����i}<�\B�q�Œ<ǰ�Hq��+�d�	���N���^ �_d߽���?d�??��v$�|k���ݻ^9N�[����d\bstEF"�^/n��؞�^�+��׫ٓ��"tf��c
�`7ީ�ޗ{�z���蝨�(vq�kW���+-�zI���R��r?fV�m�)�ڳ����N�1�p���Mk�'Qn��bvF��ˉ�\���7�g$���a����){��.��EMK%��f4�x7
�菇�����4_�?F����Tx�Ug�2��gJI��q�UȘ{8�]󹱷��|���D)A
D 
Th�B�hF�)ZR��(i)("
@��#*Ogt���F��g���Y�;Q&�l�/�wwx��n���9��<�~�k��G��	4�����~�P|�}�L�쥵�\8���[�x4\o^1�O�?܋�,*f�Us��6���4�q~[��p��Z�!|{�,�^G�z`����[�\�|W�ݖ�s��Z&�w����ro�؂�V���߸�EZ�]d��ͳI��3(���"��7t�ޣS�������l]�.bK��K�K���t�x�y�ws��N=^�_���[���磓޸������X�n��+�����7�(���S�`�N<7�����˚]����;�0!T�{�aM֫0'�ݍ��t�5���$���~|#c�%��ͳ��FS\V���4��q��.|2go^-N�P-'j�M��!�$�ٱ{oE�z��n����`\��[�T�ڋ�ŨA�����z�2JB��R!nb6����u)�Eմ\͢W\9��|�ka���-\��tErS�p]�אU�2R��]k/��ɷSw��RBC%n[ۈ���5����<`���h94zp���U0�Z�x��'�+ꈣ�,��u�]\�W�c&�w���y�Pܙy��R�
����m��JU��̺8	�uf�*���Ɏ���o���ճ*�Y�L�Ǯ���/"u̮/�Z�S(�7yv_]�8�"����]w��t�P*0��cHD���ڐ�ݖ������t�Waڌ^��ؼy�7O�HΔ�-�	�����;�a0._T�S�nU��FQ�[�u"�ȭ�Sɤ0W㟦9�{�           $�I$T���:dyב��!	É�;e<��VՁ["���{�8bl�i�Wq�y��W���m�g
�]���xN�U���Gf�r�e7Gtk�tN�[M���a`E�nCT[x��)���/Oc#c�_��ʹK�n�f>(,K�uޞ��=��M#��Yy����kW@]�8��e7�͉DkP��VB�)�q�ޫ��yy)���G��,��ו�;��*�Y��w�Gj5�_����5dT]C�.��L��;(l��zئ�$����J�=�Y�HJ]�m�R�ӷO�t�lu�{���l%�����;zKH�����nV��S--ż"hc/,�|��I/]vb笖��PҰC�kڻEַ��
�lC�wi�:���k��]��kM޹��hA>r��=�<%d;�[MEj@ofŲ��T��w����1nd���1a��IL��&d+�<�	!r?�������~��R�ږ�6��	B�P��9)M!��1�J��6�|� 6��%�=�ri��(��KCIZ�"�
���Z�)5�4$M->�c ET#�.�� h
@9�B��()�('%���L���iJP�*��Z����y�i"
���!h
����J��DOz箻�☙}~e�Ң�
��Wa�0��N�S3��^�N����*Ī.Oea:�E����}_UW�Ig3��ߏH��sןr���To矰u����_��ݯղ�g��Xr��ܑƧ�sw�o_�j�Ol��+��T��+�{�:��s��K�ϩ9�h����6ym[S��ӵ�rV4��WTL8L�f�{�,���#{;�0���3$Q�4���Qc����(��Y�W=���f,�����Ư1\w��Iu<��2�Ϝ��|�zS9��e{����*���*�d�h�|�fz����]�mŮ.=��T?Ȳ�(���\��݇0N>g:5o��j�N�^՞/f:;0�Z�ʛ�/rg�����R���J��W��R�d�(yµ���s6���F��9u&����D�{���e�<y���'6��֦�z�wMͯ5
:�ŋ:�d���D�����!�VO�d�F�`��q=�^nU�}���W�W`��S#��'h����q��}mlP���J��䞻��z3e�.vܧ�m��suyC�PQ�����F��oB��y�PO���ʧ;�~4�ysV��r��PO���S��17��M}i��xj���ElJo�h�y�n��~�S�H��f!}Vu�Lu]�������WP���Gg'7���,�O�ɳK�Zp�>��T��\�(�E'7�t;\e�c\\`n�V'��;�$ջ]S���u��i�u�a-�o��r��:���j9IDg����TJ��HV��Ɨ�33�f[{M{y|7�l��]+��DO�⤐콖��>��,����BXΐ�/*Ceǰ<���-U����C��j�{�����,I'{�YՋ�w����#Jw[���Y����.�a��*�':e�L��\K����������}�xn���=��W��p|�P1��ޓ]�\�ɳ����)Nó��Fr����7�' ��b�K��[s�8�I�B��wV:Ζ+	�yNK4���϶�̿�
���:��-uuS}��ֳk�L��K&[^����	ڂ赒t:��Y\��4��)���x�eJ�o9�W1��'h�J�̮u��Q�ɬ�w��}}�_]��{Q4�7&Qj��b����	�vW��+*���)������+lȤ�gy[~;}�_u�d��3�z���i�:qusSҪ�y��ޫ{�k��)�U��P�k"nT:j���O{jr�؞��K����x1�&�7;1���+U�m¤n?��n	��rc��`���!���,�jA�O��"ޞδ�Q+Gw^k�X=Ѩ��}_}UU��=s�;Z���SݣJS�lfO<�N�L\�?(�����6�}�Śߍo�:�c��4 �Z2jmgsN��C�
����ĭ�^tvJ�����;;�1��ξ�J��gG�&���p�;<����'8�u�"�K��&9�.�\�X���W�I&�g0�XpҌ^�e+�=m�p{�5Pu[���z�������Q��@�iJgf�A틽�Ck��;�_C{��Ȳʂ�}Jx�Q���k���^q^�¨}�yj����_�kJ7���8q��!I�z� ��r,��x��|�xI�.�P�Y�y\7�,�O��W��z63��Wj���"����OK+_���6�;&gn�+$ET�M�����72��-	:�l]�T�8rp6�n��}}�ol�ڹ����*k���l�[^QvV�����4�<oI�yX���\!3Ք�}�0,[�Y�V�sm�g��ݕ�o����&�$5�����٦
�|)V[�ֳ���'�f�\i�uz�E����**м��6��Vߓ}!�������^��!9N|��S�g{s�����k��\��	�|�o'����w�ձ�����7:EЦώ8���1�;{:���������h����.ƫ�aBf{�_� yes��ޑ#�/C���p��(�x>�J��5e�f�9�v��h^o7�S�}Xkմ�/Mi.�������L>���P��'���#L�Qx�n��n"�ۃ�����'K$L���Fnv��$W,gb��m�����Sbk����{m�͡�f� �U9��^񏜝��着��M��o�'�Q�W"�QƵK�8k��|}�wo��c�v��K}}���4:�����O��/oSM��n�se�"��FT̨*B���{�����I�J^�+é�u�V��&U�f�2�F�v�:8_#�)u��?K]�m� qOd�1��ݥْ�3�k/ޫ`�����L�|i��g�o��ʆ�ܜ�#�7k�Q[L(v��V���ih�)�7���\]R��O[�����*ߢL����u����c���ٲ��h�V�]���*�׫Gq���jt��#�k���;����6�}b�p�(�����77Ry�/eN�%-���"7����ʔ�;Zܮ�����01�μM�^Q����e���WR�lcWz�@��DGНx��:�����g\$�ے���wE')AL�Y>��f�H���}p��W��A��'�ц?k�������3�^�)�/D�=h�-�]Z�}Y+�l��RUˮ�f�#�L�W�����j\%;Q:���W;Q5������[�_t��1p^S��TF�Ƕ�>�S�����[O�k��c�}=r��z��QV�(? �|�Fh�[jw��A�ٚ��;�e�L�G\�u��K6�N�
V��s�p?}�}�ʵ@�E��J����\���3q&)��y���>��c��N���H�o�C�t9��ֈQ�>th ��}�N�c��D���6��b K�n����x:M�RQ�(USm�6n�zV���(��&��6�F�m�NL��GEi�܊~��ꯔ$�=�ݴ��V���{u�.�5����kg_�g�ìW���!��Y쳮��/IS��8Piv��X��OU�½̕�?I���퇃�=GD�{��P��>���"�Uw�9O��Ԩ�2ܮ���ǩVF.���9.n�i\y:�{���G^hz��m��3�Q�r�Gj��ů7��>�IP��>J���̞�q'?5B�}f%Qo{7c�W�uϥ�Ҵ����g��X�=���-n	��:���^X��p���$dO9�y|�w�&���SR]|�?\K���)y�ݤ��,Խ-�PVxO�r1���,L��)�-ھP-��X��V�������r.��֕�G
WD�^c�N.v+�+8�9�\�d<X���ƨǙ�ھ��*=�R�W�ӔÉ�\\W�}_|�6{�y�Y�>���#�Iۻ�{d��ߏ����D�)⚋�M������AAS-{��F��Ē�]&�����F�5]X6�N���w��I^��X�Wqr�
~2�I���mc��N4�u����8��/���ge��/MG*���f��W�oo�d�߳�o4TZ���:z*�|7�Y��ޜy���es��ٍ��y_fOS�_D��^���)dҜӄ�k������^�V�{V�+R���T�I�������h���G*���a���T�D_��
�ќ���w�'_,���-a�gH׿htU
q���CK�O��:������pd�FVTOӷT���W]���`9gR1�Z��R�H:�\Y�e�w�4�ʱ4��|U(�:� ����QO����{����g~F���U|���t��9�L����Mέ�б�<�ѥ����|�Ȩ�b�Ax�W	�{_9赓�PV����E�I	���fu���f_�r;��O;�F,�U�R:�U:O���i=�CE�s]���:�:j�^�F���r�2'}�3�l���P�Os�Z�����rx5�Q{�V���]��e��ͬ���B���̩uD.���u���Q��UTr����򭆒q׽H[���c�y�b�q���He�N�u�4�a�G����=���w��j��d7>����=�k��X��Tz���_���<�
��+u:�B^�ف��c���#:����EB�uf�k��N�o#�K�;��)A0�� X�j�y�xf��;��q��Vh�-�q�8�i')���;��$:8tN�ۓ�%���32�Ъ�$;e����o����f���%ga]�;K�L�
��\�wYd��
ZP4����\���ͷ1���/��>A-
�ٳG�,�����mk�GT�N��-�K�7�=�ts|�+�8��q��bV%� �%�'{��T��������v�Z"+B����^1+өA��㻶�Ѳ��u�'��T'��b��Kv�d��%|kEt?����2���lޣ��%��|)�@�["�NX���}��j�7����4���u�ږu��-�u� ��d"\��FZ�θ�H���|^�iP�����Z���V��c�^��9��.u��E�:�i��ݏ��7�����n��,c�E���i��!�(P�ш��Uºɾx����j'=<�               27g��U#VQ>݃ѽ�:eu��_$���7۴���:���|�ص\��-�P���Һ��hn�I��P�����r�7�4-�vFÓ���r��c'u���hm!����j������HDd�_2#�r^�v�"!g�E�tt����7aMx�(��d�,���@�t�t�Hq��[w�v�)s��m�aIEwL����d�E�dW��l���T�3ȋL�0C'1l��k�b���譁TXD`�N}��%�22�$�,Ò�Q�j[��ׂ�����%��.4ɶ/�ZM�ks'�(��/gМ�%H���o^<3@�-s�VM��c�|�U����,�ɏO@��0���hW)� w�>��B�c(����9��t�v'v�:�=֛v&��>��ʅ�r�m��77b�r��S�����Ê橙Po^"$+"R���NIM���H��=9��L�}3L���W���`�QP;T�����A��fR4+f6c�eAa��(�d�@�7�$�6�D�#0,�	� \��ְ�)�/e�%�m+Z�� i�F��2rn�L5��K�9)��BYbf�
jZU���ʮ�T���*�L�岟qcx8mj�SufKn)yɵN�WF+ڱvb���I�Ku�\��_}U�����R{3��sz���)��G'4�o ͭ�3q^gFW��s��:���j'j�e<k�z��OZ�ޣ���ܭ^���ut�u����}�F��F����ә��>ۿAO�Ϫ�z=�^���rrҎ���S��,73�[rN}�)?z%s�v�̽�~y.F2�Z�\�����PU���E�+k3�|��9d;n���1�x�N�
��V��έ5�~�Ƽr|k%.����i�j67�l�kS�"���)ƪ]�\���S��{�Z��7;���6�_��p������>�s�FŹ*/0Z�XO,u-)5V�.����ר%`'jϳ�QA��V�쮞��A[%Zu��zqg`RiJ�J]O2,��:N;�	t+5�bڝ�������.�^�-��w,ěj4�}U��<{���C[3O�gP4hFqJ��r�����To^1�O�r%S;S��b��ުV9������y����6b�%w0���Y%z|?Vs�������TS���6}�sp���Ie��z��}ܗ{�8��"'�o���_{�N`�y��7&���7p[���!2�On;lf�E��_W���a��ꚋ��U�d���2o;�^�;<�Ё&�I�V�ܟN�%�r�'�BU�BQ�˼�g��D�s䷛��<�W�̞�*J�l������q#�"���Jq�=W�sHG��1��B��IG	M�#��	�I��Y �QS��u=}�S[jo| ��r�o���H�я1?L�V��ұ���Wv���{��#���{蕮p�B�rֹ������k�������wCF�MX�q��J��}ٳ>�}{wf��޳Sy{�2Cy�Қ��������e	�.���B���H��1ιtX�w�� ���yi�_z��xq6���>��L��u�	&��M<F�G����8_L{b��z���~��C�B�{��Y�註偵>T�Wr.*�&�~�ݒ-d�8�����+T9	�v��%n�6��˗�O ǭ*�p���˧n�L�)uTB�B�`���m���T��Ҫ��SY�N*����g���{�|�7+/�m�󼨔3��^=���*�aIh&:Z�`�#�דt���IXP{[�*M}������w{�():���r�LEd�]�Z�]ՙ����˂m2��	
�[s�rO�1����#k�r\:ʼ�����'4[d�y�<���w��Z�Ûַ���qѫ���5��I�ؼ^'�������e�퇒o�ԭ�s�^Z�Zߦ)�[k�oǽ$ԧ�&uL�\�.ejn����}�.�^�oI]~���uo�G��S=[%3�[�7�כ�;��wf�d���Ϯ��rm �{�^��^䢉���Y��.��$%>N�f߳3UQ��QU����F�U�PR:Ѱ�_'lq�d,�7�L��\�0��F���Ԯ!]���ɵ�����ڥ�y�t"�_VV���}Q�)l��n�ɈдK���wP��#�M�����ۻ���l�c�i���k��<����["b�*�M ���œ���S�Y�Q�
U�G}yR%�U�0����}�2Lɽ����8��D�5	�N�;�*ˮ*�iz�Z͞�Z�P%�{��D�� 5��������
O�����j����+��6���k��qIyܙ��&Su�*��K�of?�Q��Q��Qj������&��tǱ�����Cq��-�x��fj�M��8 ���qo*�)ػ�6��lTY�������u�ոY7�{x5�9�{��!��m�j�6�p��)�A꺎�kգ��M��&�]S(8
���H7����I��e��ܕ��]RrJ䑚[�����񌭹ҙ�W_��Wu��h������뽗oEXV���ۊ����>�����+�"�՝3t{#bV������R7�^��$w��s�0�LȻ�o^�î�	�f
��Q�u̬���q���">���?N��~:k�������3�8���u4#R.����'Go+�:��w���Җx�q�d�}��o��d_K���\�^�n�Y:�q�N�k�����Kn��`(����[�2��T����O���A7�]���&�zF;�F�77��h��?�����ȸ��.g�g�߯%���ck;)�M��^�s,��P;Eѕ4�z�X��)�ۨ�Z�yk�Qdr���}#��_$�J��5��T�/o<9U��GeW�i��t�gc[3M�`K���K�W�[P��;ʲ����~��${pn�F�ݩ�%V����gs����kWN��F��g1�Ѣ_M�!*en>ҍ���8��打 ΈZf)Ճ.����g�����bB�m���jTEF�ﾯ��᱿O]�ԗ$�'��q�zs��{��_+�{@D�y�C�w%�xO�̣�ʮ�|��m<}J�]&9�M�g�%Y�-9�dr\ݏ�yϕ�ȪR�/s{���#�H��_՛��ŏU�Y&�wB��[�\>�Ϯ�e�	�����5�b�onO��������°�q3�I8I�Q/����Ƶ�1���f����P���sM�r�q��J���KA����*Y����n��嚼�������rd}9�u��� �7u��:]���:L�%z}���Gq�OO��k�*:���9{۳�Fx�%��T+_��dYUgDܫXK���H��s=�uwe�p�81��V]E�e�yZ�Fh������5(d������Ka�P���8k��s��֫��ֳ.��#��Lm\��JĪeirG?W�UG���Ny���UlDx:<��M0F����"���0f�v��w���h�{��IW�Ld~����X���v~C�BAtz��d{&{}�=�Y�ċδ��f��Ɠ�~�@}f"`�	��37y��|Ejҍ�eVP�>�<~j�T��u�ω��7���-7�0Se�Nw�U�Tc�9�����<<+�B���6?_�xվɽ�gܢC"��7���ӹ*����ȼ=�U�(�<A���s�t�l���3G��eAO�BMњ�VG<��ɋ�3���������6@Қ�D�贼]�]�y}>��6�<��$�M/{Y]%�C0�h��>(��˿��O��7\ٕ=1$�{�.��z��-����S��Ƶsu!qa.#�"4���J6*���޴j�B7�hՂ�μ`��%%�	���v����Yz�G�}|�K�G�o�#$�7$T�Q�����2�0�#)5Ҥs��}M�{�̫�����87�_RKq��yS�c�^���J�]V.:g�r�'ѓ��1�#/�7M����f�8�E8�<��	i��������G�̥�ܿ90������!��j��A��btM;.�"��#�nv�Ǹ��S��"[�a�yd=$BgϜ=7ж	ME��9PhYw�N	������V�-_�<�[���x ����y��pp�0�o�Ey�=�`O���W)p�آB�u,K�֨5�W����YQ+��������"�
�}@�x���ܻ�>,�<KC8y���_�96Uu�̓t+\t�X`��\@�g0���<bͨp�(~�x�{S�w1�߮v$�~�~��PoʪI��dH���W(f�.v�+����;���Hg�D#:6��� ��\����̛e�1��d���v�{5JQ��i=���o���-��lk�F�ө�{L���i0��ܜW7K$Νi͒R̬�H��r�h-VTO�4^,w���=�
j7?}U)�/�{�k�^ٞ��b�_�#	�B��ayq謢z_x~��+"������)�]�u�OGދ~�W�W���3l�1PTj
�g�o�xb*'&����x`�Ƙ�X�TPy��[�W:�B�o���{g"d�mK�c���w ϴ(���{_��v^ۮu�}���Y��*^���U~FVp�Q�M�2��*���]�?(C�]N
��9�;��ޙa����G��C�XkL�l�!��׾v�,�����]ž�؂=�� ��X�Ը�Ǧ �̷�P��Y�_/]���nN���U�>	�2�h�F�`�X�rĴ�[�C{Fz��J^���x&���*����K�qX��+4��<�Q�ނ7��u�`p��q�~^>�]�P�::8L�����-��K�=H�U㚭{=閕[F�jܬ�9|�;p��'6�K��҇,�I�(��o���F�D����s�U�T"��+>����M���Yo#7�P�l� Z8�2����լYZ�P�7ª���V��*�V�V����8�:�`�v�*u�lK�3�m��0�a5�[�#ʹ���V��;/%E��T��غ�c�N ��N#u��b�M?lO!㳕����-��8�=���hך0R-��,;q���:E�QU�k��]K�tz���k��Ef��⅝0�cm:2��p�T���q/v:ә@Bu*��'�Z�t�]p�(Q�W�B��#��(�6�vbc�^�.�޸b���{�B�knVQ䚈.��{��L2��f�r��K:պ͙r��t�
�i���$� '&jQ��J��y+�롛0�sR�Z���u�P�еEKKS����q��ǋ�JS#��]͞��O��7M^�9,v�쫨e@���͆�`�               ͝�o/j�f4�\����� iV^|vٓy0���`_=3dm�֥\��a*OYԩ�ط,Rˎ�V+�����^�C��]-�r��P��-Bn�It�Ӄ���P@n��S�αy�끛gz�cB�.��9�ń���ܮy�W*�Y�'&>���]ڜT(�<Z9\�'&���a�WY�w��pf�l.�L3
磘�VY'���Bڻ�j��A>q�ian��vRU(��y>٩�>j�O�$u�j��Kgk0ʳ�^���6�G�mo$���N;��e0���;cd�����B(���y)�آK%R��2����'9]����a1�׊�	hդ�:��β�d:���V��u��n<G����E{��o
���[�u���ĥ�	�ͬz���[�1|zSs.�$j��/#�1WV$T�����9kU�)�Pd����ỐKY���ξ�͙# ����"N%�HRД4�A�A�G��-NK��.���(�#y'Rj2��X�d�NF@a)KJ4��$L�+@�P�#��944��J���rG' ��j��*�(r0�ZӓՕ��#*L�S##�ȡ���A�eHd&Ag�?E���s-ֿrxamֹx9O���L��p±�w �xܔU��u�����W�����}0�����.��ظ�a%"���s1E�a3to�х؞r��ގ��DH�@�=��:~7�N���5�=��3e��&���iO�5����ԕ)�x�Aֿ�V��c<�ի;�>�[��2Wo��ph@
���@`c^<�����y����*�VƝ�`��zI����ICƶJF�1<���V�_��Cr8_�*��{ʦ_����:Ί�bP?�^��h����>�xU�Hj0{�W���Y]o�&���O}�O��j֘���[����) ���J������;��Y'��%�úW�"Z��Q����ɽsw����@|B	�$���[�uk�H�Q����Y��{i��n(�R"�ؗ�B��xڼ��)��IA���|���:�ﯺ�gj�c8f�ѫ����������xNU��^��Bn�`Qc���(�"&���R��ɉ�._�[�|.�Ҩ^Y��u��n"b:. Tᕩ)�;�+�"t�O*�U,�Y�֯�wF$����Ga,12-��1QP��J�K
{�~��b���]NL2�s#X��SE�$�-�EI]w�:��b�.�0(j>7^����p�o;�>�sf�f�==�Yf� ��]z�}~�2,�: ~�Z�\x�ễg�=7��9�Գ�Z�$��G|������+8\^�&�Eۧ�7��~�r�A��\ۮ����(y�^U�.�Zh�kC��YX��^��f�U�=U���^ :�Dc��N��6j]j�_.b�8C2w�a�v̜�����������G�%W_��k*�<�f�ۑ�m���F��pU�<��F�Ƽ0mo_��xy�i.�C���Gvֽ��b��yM,��2�\W�
�x��n�τE��7���*�������G�*�S��y�ڼ�&�#���C��{���'��u�7��"�"T�^A�lrT����FgTP
aU򗓖=�r�$��hlЁ����v�a�;g�.>�z{�%~x/��S68:<�5t�p�� ��'S|�� �x�_t���S�V�ɸ~t5T�+��T�������{N'MxK̓ܧަ�S_u�۩�q�`�7lP@�t(�R���s@5�+5��y�@�9��D���Z��`�=P��̮h�;WD��Wm�;�*}�P�N��u������>��(=~@h�i{+�4zQ�&d�B�#�S�p���jϮ"���᧳k�?v���3���2I��<�7ir'L����-
��Y�L�v_��Y�Z�8�g���y����mW�D^�G�r��K�?�PB�
��8���gAW�j����)�ΕDI4����y��g
�5�u���o�g(4�xׅ���(%��(��KR���Z0{T�L[��� uf�G+vRW*!��3�TcǬݺ�	�E�Z�����xn+�< "����rK��FD�w�ԂḦ/�3]	�Ѣ��̦[[�/p�ˈ����$��o;��y�uƟ� �d��{���)V��Kͱ^+��g�c�Ji���WJ�� �8f�<b���f�����=}��Jp�):�(�U=Z�$f���jW����Y���y��w��=�~�@C����x2�X�'u3�Z����̝�D8#��/��P��:�/�<O��?YUn���AYҢYB�os��Z<ߺK��ʘ/ѨV5]����CZ4m�Z����G�J~��׳e�C�E���R{���)˛N�&�Y=���U}}�Pw�W�56�h��s#�3�Y�i�GL�o��;ŉ�:���#�V{nn䍿q��>:t�(Ġ�#ZSA����0?2�|�r7Z->�wu�0��A�2�ZdV�/�>�!�Ї}kG��l�hۘ�ٍn��API[X��_�(�B	��h��aEj�Hi���fv��l�*(�r+X�mn5�*����!"������;m�緢�@jŘtQ��Q����.;�����SX<+�Q�+~ԈXa>�ޏ�#(��S?Ϻ�wg���j���7�_�{�ֳ�C(1Q��?F�ݫ��b��}K+�)���d������>��âdV) ������/w�z>�B��C�n �C�׏�<�]��Q�e$˨�KW,��Zװ���4,o��n��pUqQ%WB֗�g�/���WL���3u.��"9�0� �躦���_ '7�UdٻIf�zG)���=&6��	����!�J�⏆�F��#a�R�s;�#����H�e�E��,,z�� 8xL8|�_a�]��Y�y{$��V� �3�}^�{̇W�^���ϥ���f�[�8�+:�)���A8�|��������E�p]O/~��Y�S|�&�c�-��{���t���Ӗ<��c&-��ǳ�((�U�̠�R3؟���wM�'�,
a�tQ%��;,ވT�f��}z�
�=���D�Q�܃O�G�^f�u�7�����9���*����Zb_dY����!56��z�j�{�'GZF�����h�XeG�3�@n��W�Խn��U�7g��=]ŉ���Cń�!1Bui�����ӳ
��1�+��U2R�i;͔�2.&/-��u(�"�H;]%�:���0,�h��|�����1���������
�;\@1")P�]AQ:=�����n�{�"*�Vn)kc+��e
W�_[�wQWD��F�-�͑bro��} �
5�5�W�������K��uyI+ix����X�A�{/�C5(�_b_i�ƅjŬ:js�iĸ��t�eK���O�&�Q���.�I��G|��ң@�5�iU�ƺ�y��Z�,�q�[7�3%��*����P�8���L�5th"wn��A��Q{��Xq�W��3���*_7�����F�YU(��W�w\��
�۹4>�f]�X�S�V�UϠ� 5+�j)h�0n��+Q��yM��9�����'{��O��+��e_0�\I�揺�2ڴ6���1V�`P�
���[¼�p�vr�`�ӿ.���7�/|����흸~��C��g ���	i���C�Uq�L�[��j�WZ�����m�j��Ν�툎u�|]Y��੥��஧X��TǄ��چ�4�{�&�\.�x!�S0�K����Ƽ �tJ��x�w���v��jE^i���ˢnKt��P���cvs��f��W�p�4�S�塘n��;5t,��߹N`_W.a�rKN��j�^FӖzѥ�oQ�pK�3)[�%��ů�?y��S䈅����\ęEb�yn��"'_��W=�:S|$�QCK�<aą���V���>,��V6`YeЛ}�0��""4s2����r�l�흩�[|hӬu�]Ң���Ίe���a�3X�_4ic��48s�5q鏱D�A�A�Aw�v���~���!%E�q�\%�X�S�۹�(}��r4��
�W�tV;���.����zk�&.�����!=�H��щS�Xn�`�I�#�S��v;��2�bDzu��E:T�4I��-�\<�hU՝�ꃫΝ;�f��Q��2�lJ���*$*,K(�͡i���d���z�h�M��u���D�@`������Hb�9�s����G��B�W-5ˏ�WJ�� �zT5���u��6������GM�-�@�X�`�\��(u�l�VC�1;=��XO"�:t!�K�8�i�Z�.��Q�;ь��B	hU�8�z�Ls$��p�Kh4�.����vx���S��.6�<nr�m�^�mʝ�$���WJ��u!���оlCz4o�.��X҅�#e�V	9vw�����ʐ���d��H������z�r=�z��H�2Z�^���s�2v�����tܾ�Ar��?%>����=�9������-󓿟Tey2痰0���w��ش��+���v!G�����K�9O?{v]ؕ~�Ơ�^���:Y�i���8gx�3~��깛�Da����a��"H�%�*�Z�SO�n'^�Չ�C����MDW/Ԏ�+OD������C)
^Gjf8�.�޼��ϵ+�g���)��Z�'��>2�n��^�����w�APx�0��?o�9Ժ�ؤ*]V���0(�Q˷5��o|qሱn]{Q�t< A�V�h�8)�K��#5�y����):���Mc�\�����n�{2���y7j̖Z BN�u<��t=c�hR �wp^l����4^׭ww�`e{�+G$�3��QL!�á�|���~4����}҄f�[��z��8P<i�%U�=��;�p�ɪ	�i�'�΁ +3�΢}�w��iq�[6�v�Լ��l��Eލ5�x��N�Bm��=��k?��~��+�b���j�t?����N�T��E��U�!�G�O��Z��q��>���X�y�79pZx|�z߼qб㮖�������n�nw��������q������Td�;!ߕx>,\x�����wgOI�K� Vw�_�*ipb���*�|����^h��k��.��7��̲��4����L"�~cA���A��f�~�Z�Z5m��z7=�XN
^�ʶ@�P�}pe��+n��|��P/h�'��K����i�Ѣ�5aQ,�Uǂ��G[���L��/n���w�a/��%�vS�W���P8k0*$ l>&���9.�^\�M�?�K�d�^����(�Nt�����Åu��&e�>�Z.I�QQ��-LU�3������H�t��\*}_��n�=��Gs�(~d4^G�y��b���s[�׏��m���4�f;%�]����õ��#iP��M%Qb�P�͂v(�S^�\l���R��ǎn�s���%�+|��\�+'%�]4/%.�V,��ĬJ�2\�!{������~0��ux�2�%�}�� 튃�z9E>eV�f� �	vl["�dy:v��+c��#5g�ӷP�nTX �؛�/@X*�ɡ�*̙gDޘ[]ֺgȗ*ܾ�\�͊pՈ\eK�Mn�f�J;�(V�@:�va�wbT�!ܱ�ys�	�UZYB����GI��/є!X_A��=�<S��x��>��^�'4�J����w'[���gu2�|@�q��㭭ř�l��*�z�:ۊiu�ڧ�Z��pH�^�;%�Ho����Of�6/�mE��cU�v3���bn�R�1Z&��j�d���&j!I��J�]�D�H,�\�"՝U���
�)#w/��鉼��lm�WT{���             I$�I��E1�a;5�BZޢ��)�M�ZC�Mm���x�GmTI�����
�v�k�n������=��R��].��ԹcH-S�f�x,+�]f�\6��b�*ѝ]�	W�S�l3��	�S.k;��Euج���Ζ9q�G,�u��l<7�&� M.��)��F�Jѵe/-�2�U6��Iecjf`$��p��ZMG�W7�5O��΂��-��u?��4������(�iKz�t�{�:�ej����a��K"PM�;O$9[�N��c��1A�:���u��3֥I�u}�A�:��_e�9C4�!G��ۺ��s�����n�;��ЗFf��	�Bv-W}h�t�k�b�zYsHGRO"����N���d(��8=6��i��k���f�j���796[��W<�҆vwD]#�4���5r����d*�ܙ #�� ��!���?LDA?}���CP�"P��Rc!���Xdj
 ʚ�jZ5���-fP��Lfa�ـ�NKCHS���$ȣ*(�','�Ѩ�%Ȥ�2��0�(�h��,k#3(2��+m�lM[`�F4fPd�O���̪rL�lƲ-��^ㆣ0��0��+�3302lr3)�(��33#3'#&rr#,�,�b�(�r���p��0 ���A�
�#�ͻp��upr���.=
�L��1�����T�؊f⮘0th!�����q���}_t��{ހ���.�Qv�/���B�V��4�YJ��cQzxq~-Ov�ۚ�u�g���I}�
���7VtA�X���L�~f9�'fu53��C�����i,䎟��Ec�+7T��褝�n^6=Z�g*P�Q�R�2+hr'�{e��u�������^�&l�@t�}.�W�F�HHR+���e��\~�|o�~�ܢ�삮����U��jL��p���
��^���4���Y^��	�=�ܮ7���l\By�%�n�#����I��Y�YZ'�G�T�MexةVkG��;��j�jd�w_=kǭe���)jTD'V��̯]&_z�/0�ns�	^�<GANf���P����^Pl~��>K��wTQ�G(��E���� �V3�XZ��!.����>@�݉f;��Zͪ�B"����0��e�Y����Q)J`���(��8I��k]	F�=s�ͭ����~��n$��H�������Q�)�U8�< �)|�,(��q���/E��f�A����Q�~��Ҿ��
��Vw��vkj82���DJH�Tle�XhyC/ψʏ�^ӕ���v{���魁�Y�7dz�p�w>.rե���C/�M��B�gH���l���u	j� ��_�ֹ�b�G�{u�F���5���I]��zt��wKL��u]i���\�iĘ|&U$K�ʉ��:�RV��oTt��;ޘ�f�ג�`���ִI��t�<��R��f^�d��飾LZ���)��iA.��!���U���<�}��}C��#0���-A��S��^u\ d��z��j	����r�u�𻦅�s�V�"��s�+������������7�E�� F��jF�� 7ei-!y$;}�6�]^����&b���oYҸ�LX@��TXegV�JB�J�8y�ȩ�H*�3O�m�=�jb�sJghW�r�!ԙ�&�F���Y;<��V���b�:��H![ϧ�����tR�DY>�����,�U��eQ5�kBv�aq���{=�;ؠ�8��޿�����޿3fTWV�&�����H��nc��C�?)ތW�ᡳ��0y���Jt}�LS�W�[ҷj�����@��4���W��z���I��2G��T�ޛ�խ��ey��ELl�0��0Θ���m��!{=\t�Y�|mS�rz���X۟m}�a�m�Za���M���
���G1h[�[�7n�����վ
�J5z�< j�G`�Ti!��]`3ޭ�&�Ufb�P�Qv�m����P��H�U���� ��w���F��wws=#�,�B�Z*q��*��}4СWC��1	c6���'W�5C�f�Ă�A9��d����[Щ3n�Nj�=8�W���-�m�ņTyu��dN�^ev�/�i�J�!���JA_����������[�s�y���Ϫ��e��<���iS>`b�ջ�˭
��'&�S�M�z���\W�uwp���Ȳ��Å^�J�x��Sp�#7d�=�Mu1��R0���;��Q5���+��ٚ���@Z�z{�*��6�:�؀���Z|��ߍ^��f��wI6�B���J�~����jF�=z��T��}�S>�l�왱p˷F�Yء�.?l�!\|tz�T\�����~�[3�����K�� ���ad[BΙJ�d�<w�G�!�ʍ���Í�Uۦ�h�����ff1�)���C/3]��p?�~��G�����ݽk�K�x��r�.$��h0�}�<�W�Y1��(�yHX�EOUf;�M�D�VY���T|X���t�Q���~wmV,Ŝ�U�C� Q����Xł^'���YĦ��`�5M�%���K�i���"����s�ZϊI���=�{lm��\���x����1?{5���Gi���erW�,�I<|<=b��]1:a�м�d��VH�P!�}�۪�5�%CYQꝚ�zg�g���y�k��wox4������~T��Rf��4c�¶�����)[�c3�ozH��h1/�=oE*~]f��<^����Ӗ��z�^��Z��o��w^��������1p�w��Z�7�6�5k�}1=<�A���K
��r��B'��2,�åo���Zf�q����.|mÅ�ċ�i%3�:is�4�g)/,{�������B0���*�*P�ؕQ�R�2)md�J�hNaw�w�`��ƪ��AZ����·���:u[���,�&���zrk#I~�S��b����Tܼ�����e��j�|;���=�d�
**U����pS"�A,���<���o+p���e�,�J
�OV�^�IP]�{.��1��9/v�2ƞ�K�����n�
X�T�<�~������b����[�F��G��q�L�b�Y�$�*��q��ܝ����y�) =���i���!�4y Y���C��t�ٛ\(���q�Ry�Y��jLR�VU��%�sٙ}|�[9ݺ���|U�-q�C����i���#�Q�L�;�)9�o�g����xY�b�Q���Nac����`���g�\Л��Dz��N��6�����ˉuz��lUK���Y���W���St8ϒ:D�����nV\e߫�u�0�[09������޽t�-j��0�<t�@�-�U�7%�lb��2u�WK��JjƠ��}�E䕿���!O�Q�f9���{g�v��WY�����Eǩ3�:��$Ĭ=pK��x�Z�u����E��ջ\��
�ށ5}���B�&�&���o�����錒���E�X1�M�`�r	����(�Xݫ9oxZ��=��9Q�z�w�97�7�Q-�AW����<]#V��G�-�EF��Z$ս���s���V�wh`c��y��5�\.�B�^҂\_b��6��)�Ξzɱ ^��j�� ��E�������\�yE�H����1���>Ny�/ŔD��e4C�qa�B�����s���c[s�͗.���`�|)
C0��иߍY�R�$*�*檓rq�D�1��*��>��� �~�@�b��,Z��[���7vL}���S��?[3���_��/NEuuH�`��AȨ/^o��)�vU�w<oL�͈+�N����5j7\����Z��D�jdCCƼ(��@�y���I�N�&�Q��͚�G^��x�z����$a��bL�[�b���"�!��Ֆ�Cڶ�`��ˌ�$V��u�kU\ed8����R����i����(jX��hf�6��X�gG.�f�E%�e�^<�J��y��QC����gq��C]�3'v.��=�n7?UJ�$�����TK>@�C�^W��yW��o概�WY����4;a�/��C�%��*^U:�F��Z� ���T�M�˩����'�2a��QEۭF
��!r�H�Xa<0{v��~\mߤ�V���v�U�MZj
�~���\��T�T(V�������|O�,��،S�Cfz1�&<a�`���~xvO]��r�{'v��g�/�#,n�����eC�W�
�A*�e�^�%��f��c��-�W�i��b�3j�����*���NI��%��,5_������G�D1T�-�*|���k�-��L5<(#^��zy+�kR��.�b�;�w������G�M^E	�z�/L_yg��*�h�
���Wnt���r=.v�)�f i�9�V_[��N�h ��]%�:AU뾽j�COE�����~���J*)�ux�&'�Fᷔ��KF�ӕ�2%��[k8i6�G;�ķ�Tf��~��`�>7/��՟ݝm���:����Sj�U֥p�Uѿ�U U�/ *��
D����b��y��\���|�z:m���oD~����,:Wʒ�K�?!�؋LK쉻�Oݻ�� kK���n{%w���0��fgW�D�2�p`�K���Q�FtF����ڛt�֊d� a5�+ʛ�q��7�y�#̨À_����i�o�֊�4��P�02@�m��a:���o��%^T�3���/
�9CZ�.mm1J�.��������"��i�!�O��-BZ�nN��󓟢[��F�ٙ�p��=
Z�#@X7E������:�O�AL¶��=|�^�nR��k�Y�%�[���oECA�6�� �d����&�G���g� 91��[W;��
W|�	t�:����w��8��)x&�L�@�Q.Bl�|V�ܗx���yM��,���Gb��oz�o�R���pޭ�;1ߥS�>��\�*(�I<掚s�4����N�0�Juy��QH�^�<W�<0�y(9����)u��7}$��r>.�Z�*Ă�U0h���O��ʧ=f����i���0�](���dxkG�j������R藨��-*w�}"U��ط^+��J��]iB:�W�ǅbUl�#ޮ�6zs�	���
bņ+*��g��: D׃��}�N�t.nt�G�u�������sؾ#�f���@箱��Of���&Ł�\�&&G<���R��`��5T��Ds˲��Q��)1���zC����<���S�8�r��0��K�����]Iq~�L���Y�"y�Ub��W��>|�*ӁV�S���*���g���#�ɨS�ǁ��]�	�4�2��k�Z��GzD�I�%�]佣A��f2g±'��j����F�X�4�X���9�{a
;Id�p��A�3��r�<tN�.���
*��m��aY΄����Uo�\�0�0��ǵYaCH��wF�gDg$Ϳ�U�W�b��6�t>�1�4H��p*8�C3,m;
�EpПB�)���׃�6Y��^fs+n޻�P���Q����i	ܩwuo"�ٷYk�`n$;q�{y��Y�t�S�a�-���hn^��MleL*��l�� 0�Ag_*��V�*Oz��+eF���
S9_��uA��5���%<,78:N��.���X�x��;ۄ�%*�ƞ@s��.ͩh�$��ֵ��I�Vi�TtS�
���;��y��(��Fwj��a�O8�[a���wE��"H�W�F� _0C���f��O�]��'����E��Y}��@�>� ��[��kU�Է+z��۹��           I#m�ۓ���1���ڏnּ�@�[�Η��0r�fZN�� �6d�X��n"F\A�{�����c��Yġ��VR��d�]�0�\뤹�����E-(�]�|E*����wԯ�bt���˗�w-�B���dMj>�ЍJ[[�Q��X̏�(E�PWVX�F�htu��q����Ur�b�:Q�+��v��0��n2LЪ[�Ob!�ME@Q .�2k��2�Rњl�x���W 4ɴ�fIָ��=�_�V��=U2��T迈���9i�3�1F���Kflm�&��ܖB���L�B����nrԈ/: t��F�W
]�R�t�V����5���uF��Ժ"�X�jF��ɞ%�SH��S�ulv� ��7�ǵ�ۊű�Y�gT	�������5h���PP:�r�8bh���v�3�R�i�jɟX�� 8�s��lل�r�� #��"ʋ������ّE�Uf`��ޜ��9K��M&Ed�Τ�a��e��d`f�fXEq�U9eAE��U�Zl�+3��,5dQ�kQ�1b�3��DT6��;�V��&-`e�a�kF���(�lj�s���hĊ#YY�j�-�mdS�Y�c��0�hʹ��u���eNѣX�4h�#���ֵAQQU|�T`��p*�pѱ��qV�ˠ����+�O)i�3��Ƴ�q�FQ�!J�;���/��M��}y��u��4||+�"�K������<���k-�K�TO��ٻ�.�8eAj�`U����@ׂ�kgQ��́4�j�<Q�{�sM2r_�G�{)h4�����ñ ~��dZ�/j�糺TؼM<$h��ǆ���\�4���ç��n���M�~�@����]#V�*�$V邤t�Q$�S-��v�=7�2ppS~��h�x@hו�h)}{J	֗3��"�Yy�{ӟ�g�Q,xI��}���69}Z�U3�T �B��|��A��TM{���x}��L颈�H�G��4*��.*�≖��$�u8o$�u����rz�?φ)�������Ɗ�:��kp�����xE�D��j�lW0E��_�� K����Q5�&�Wk�My�2p��j�d�p ��^�Srm�i���=�馷�įW�55��KӸ��>a�f���sN�k���z�9G9
s7��Y�m�ܕ��cG*�u�������~fT/NTWH"`�t��ޒs�z��2����;�+L�͇p�:>��)�s��[��<��c��4��^�g?x�py�\89�V=�P�^^-�ޯ���������R�0��H"kE/�J��Īg|e�gF��E(~oy���-�MB٨8����[F0�s��=��%;$���a�!��P�[��*�[�U�eaح�=���kf���3���S�U�n�!�!J5���'���a��r��{��~T�yڃ�|)�&��}V�����Z��ilS���^RY�ApV�j�KlJ\�0�C�P���)�2L��w��oL�v�Ԏ����5����i�@3���x��7��v��0�vB�ѭǶV"�S���F�}��g6�y�P�����7K���֪��[\鞎�� �˽�i-���z�i*�:�N`�K)���}P���s�u~�oh+w6vԽ�YC� p~�Xk
�j�pRW:䖯�x�[�ov�:�hy.39���x�ҩ�_b#ЁHX���h�V�quѦv�{��i^5��(#]Aӗ����*+�������V��L��\�"r�}K�Lc(0��Ph���^�=\t/���YO U.��HN�^Osn\�Q����E�,Þ�ݞ��>ґ�q�f�[�$��{�!{�Ǿ�o)o�^]�V�Ii�E��7j����b���gM��f5�p�e3~.���Eb�A׌+C�+Y�'s=���Cvk�.�`�B%�D���9�I���>*�<���a^�r��p6����u�)���^�Et�����,�&���Yef�^ޚ����zϼH�PF`�}�LU᥶
9C,�{�?6t���חVCS)�RF�8�ȱ����z���ӂ���h�"�le��j��Men9,����p��ֲjB��˳$Xo��3�'1�_Cw��O�S�g&������K��k�י��r����*�Q�lh}.����C���h� ��Κ��%�W����*�:�����6yW��V��]>���S���7�V�N�g[���7�!i�
��(���*���h���%� �)r{�%ئ+�gչu�p��,*U�$��X�1S�u�i�G�U^���ό��\aFn1�u!:�&�e��C�W2iTlx�29�xW_biY>/��
�2E���K��D����&l��KP�.�V�W�4������䍴�X�}�=�wS�$����W�!��T����y�m7�i��s��~�� tQχ60�Y�����=� �W(�[�������w�AQ'����° ٲ�r/DH���)������|N,2�*���h���������u�d�#-=��Ƣ4ڈ;`RQUˑ�j=�N�89���o�m���E�۔(��JYG�WA�v�WN��̪��;��l�r`���?hwq�� N/a�b�����^��`˃żɮV��7���8U�OK�Uqq���������Z��*�%���uf6�,�ޤ�:=5�r��Pc�5���*�o��:A�/ͿN�wv��b����b�mi���^;�(����k0�SR��z�xW *���U�41�i����ZX|��<��ٚ=�B�*��F��Ȏtx"kM>e��w��W-�vK�}x�~�c��f�B���tN��h|�D��#��$��ld�I
�A�>�q�\v�<6��t��LK0�U$<zzt���zm��i� �$U�����dt����s���݇I	8�%G�������Z�^�^��O����h�/�T��n:�MfD�㩓�cM=�˿���I\�JW�VŅc_/!��Ȓ�,�٬�ʾ�f�Y�U�XkkS�P�i8Jd({�%��d�r"�۹|����g�];�>�r�W�ApڬBj_"�k��^|+وz�cVzf�q�'�NH����H��h�`ڼɔ�;Õ���[�e�T���H�������WZ�)�u���
��;k��!�f߮n�o�?Rh��0������(�����>�O5�Z��}�������^��x2�c���'�ؾې�S��.�>�r��u��:Z�K2 !�����Ec��ٿ�AY:睍�ay:�7�oEu�����R��@�BҸ1h�i���W�9��G���ٝC��_������
��#�֊^�T������s��[}ͺ �ҶT�͚��Z���WM��K�.v<Q.��=���c�-=`���Э͍�j���9�`5Y(խo  m��x��	�G&v^��}݄�uۘ���O-=�� �;w�LU�#i-ln�f�*MA�r�����&25a�: �{����aQ��w�6�9���~\T���c�'~������F�ZU_)�YT>Z�&q��h�l�A�w�Q@�'�O������e\G��~�Q�M��ˮ|�Q�V���q9��ӻ>��0AXQ$f��ʕyS\OY�]������N��u�K����\�K�c��>5�G�S��iu�
�"ʫ��m��[�{�X���?�C�G�o[���"�T p�5)�I�=��(����{y��}�'#K�Db�s2UT6;���͞"� �����J��Ei�	%�����égڏ��1�vLK�k�}s3;��'�=Cq��[�V��-+��R��k�AH����%�C��Z��uǂh��X�yU�S�ȥ�\����!e�2�x���׼z)��
D�����P�����2��o>����Sr����U�Q𤺝a�R�w5T3�VS�e����\³��td��J6��ބ�V�n��Y�-�-)�9��rpv�jm�ċm��|�����.Yc�W�@��VcV)F�\�~ AiB9�%�͗��3�_K��3���KC�� �$�٣A/�� F�N����h{e�Hh�
�3]�{i��>P`N�����^{w�����*P�R$o��GN�̰/�z�n�֥t�+ou��~͓�!�āe��∡�iQa�s�]��b���uǖo<Xzbv���a_�̧w�+� ��ut�^٧F_�Teי�*�.ob{�4#3��~�iқ=B��QΈ�� �^OB�z��(R {Oc~�;M,
�\=���.[�5�#�b>%�¸`�4���I�*zd�'k@�hxE��L��:+�y�/�X �b��==���/�X��,Ձ������,�
�$6"J������^/�7r��k[[�ٽ6�G��.JDv��*��B������iN�XZ����.�P���temL��fAW�4�y�5!zԥc.Bͥ�4Q|܎~6&����&���S�.�8�x\$���\ {)p�Nn3�;��{�-pKt(zڴ3��4*��r*�G��;�B�W��տ��R{�9%{���k˯�V2��t(����\	���m��K*t�|(p�cԶ[�j|_�Vx��'\y�IE�I�$o������H!N���]{ٔ�8�����g�K�lBp�-�w��;۱Y���q[JLu��6T����to��!L^�-�T,�{�=�6M��`3��E1B�NCG��K��u}<�Ez�_�ut��l�d�y�.�tz�}w(Sο��Nw��t�	�4��
����Ā�>�kUF����x�d����+U�i,A䁣ɮk�n��y��ߍr�[
"l�C~�h��Ha��k����}wp��J�jX��c��65b�q�t������F6m�lK&Z��N�Τf��*.���9�w�rti���-^`�nz��Y(�C�
!Gr'�������E��W����{���A;�i�_nkKAIԹpK�Qo!=Ǯ'���	�>�1����T�9V|���u֘r�th����\���d`BN�;�z=��	��Bg>�J���^Ţ��X�r��z=�S &�\&]��BPי�t�^�O=����ʴs�/�9 khk$B=��:��w�x|*�� �F�qH�c�{g:�!F��)�R����>�5��:2�����ZOz&aL�2s	���q�\6v�3�DQ�ǁ�h��B�����߽���y2�J�N�B�_��T6?E�X_���D���_���W�����1�!ÑCҽvR�,WOg�uC���(����?f��9jP���j�����x�퍛�ĺ��?m��?����I�Vb�/�z'� �g����i�ʇ�Zz4�n��+4ԀJj[˻:9L�C��:�dn�S�}1h�9���k��WƭZN	)�oJ� �3o
7Kn�7�dP���\�[��S�,���S1�6�j7e�b���q���B�.���!)i�5v{����������J��q���hF�1;��ߙ�bF�N�'u唟dwfS}����VJ�z5C�ΜmRͶ@��@h!$�X;y��(n⦈��я���w��RPNt�zw]�g�Pl�D˧}]K�� �B6�*�KT��.S�5�4+[b�Kr�4,�%퉩$թteJ�&��q�ݓuma�Mkw%*��k!��HÕ��#5c���uw�J��G��TU:r����Ys���yci_9��U��V$�aZ����b�窢+f�[W��V���K����kH
�c	u
b����B�*��;�h���*npX!K���=]Xs�8n#~��W��               ����d9��/7 Hҗ�A��ž�GM�Yى�wsZ
�D+N᳕�E\����v����	�	f@%�ɍ.�S�w��������&ҊTs�����l�� ��o0�|/�t契��1�*,��%�[���r��+Y��ؐ�h�y�G <8�įaԺ����U)��p�:�$L�>�Չb�M9s����0WSt7;�_
"��4�Sum���¸
rv_/�E� ��h�"��7,s85�3e�Uk��rث��s�%��ʙSF;�v�����>���]s�ᠿ��2��-��;�(���F0�j���kh�+��.�L����9�
ڝ��̢ mV�t0���V��%f��Ѷ�SG��^
�g)]���lb	4]J��,�#�/�j:�%�#h�E9�X�٭�i�}�!�.骂��v!.�Ĥ�h<<��Gfv�vAܫg����6��~�i�h��,�0��Yd�F��f9�DLNM�u���4R�T�CKY�I�9UF���00�PIPQf%.T�Fe�YNf�ё����-A�bPD�CG��%��\��#SEST&Y ]ᑬ�(3�C-Y\��\������5:%"b6�
H�ԅ�SY�#,�*�,���dQjL*B�����	Jh
'V�,̓�r�eUfPd�IBPSu��E1U4�QUg�ǝ�9gh�s�θh��c�y�N��\�Ъ�eX�[c�G��Wc{����K;��:Z��s�_��oj�5�Xt�#�q��6t�o��
_q�Yٛ����i�l���Px����x�8Mh�������9Lm�7Ѹ�@��w�l�j�x�2���xi[F0�\`˪��C���c�Ö>W4m�6���^U.�W�`�@�?zQO������lu�R:=|��
UW�{�v�m�Ƙ�9p!t��-<#��󳷹Ӥgڵ,����Z��Z��*�k��v�sd�����L�W�h��!�L5�X��q.4-B����St2�s"����
�AE��<*����$@�+��?����p- ����������}A.�4A��p�*
����;�G�عh�}箦7�g�K�c��19�\lg31�p�d�H�'��`^Ê�ߓ��:%Ҡ�Mr�&;z���F��8395X��؁Y�UԍsJ�	MG�g�/���YZ������W�\��.1�+s�Ҫ�Z��C�y��{&3�n��e�[WȒ��~�R��򃉾�t�J��[�&ܝ�ݜ3�hi?*�Q��Yf��g������˩
e�Bjw�tUFJ���/!_E~T8��ii�&r��Kn�ei���"��ɻ�_϶��/`o|�5�R��	���*������\3�{S����u�������]&����5��
����0��Q��ٽT�>�G�į]}�ܪ�5��dH��A^&�41�
m*~�{}��p�T�/6ତxH
g¹�罞ҧ]>(i�<��ړgw]եg
0.ze��7�5�0N��h��]j��]z'%.n�2�l�3e�L-)E�}KM����>�0A�#`lK��ޞ�~Gj�Mͪ��I�B�n��<�#y{|���H;S�.���&��Jk���A�E*9�Ѡ�_\WDoIn��t}��$���Ea�:����y��4��ZR���X�U����f@3�e�1ofj�MF��n�qOޮyu�n�gßy�w\��}��Ȋ�a�^	�U+�/{�V���Iӏ��z�+A��R�0�m@�XT�؏�'�A����i����GH^1u�!G��"��K���:�ʞ+ʮ��Iu���t��I�]���q�?Y�F��֏(x�%M��]C;��-:�A_�zOt�U���HhR��'��t����sEj�<UY�ޜ6*}=�dI�V[���!�G��Iϼ�Rf�U�ٮ7���^._ou(ϷޡFZ���E�!�4��_�t(��~�/���o��{�f���J����G�f�b� `u��p�~(�������\�=�lz�̦��WP�ث\u&+\3�0x�KR��=��>�Ÿҩ~�c~YCz�{��Hw5����uAN xWJk����} w#��9g �Ѹ+,@���喌|�m���+���{ʝ���ǔI4���#(���P��$v�ɯP��;��M�d<t��j����/�{.��?$bi��J��LB����B����5����t�\�W{KÞ�i*� �m��ntgC����X�>&����Z�U����5�*�Og�5���1��Eֱ}��o]֎,]\2�hR���� � h����]�8䴖q��So%|#'�Z��$�ov�y/����#¬���	�A�(gc���X̔h֤B���4UE���s�:ϕ)>U�k}i�N��2r�Gx���\���ۣ1:��Z�zxhp�_�p����0p�Z5uƧ��Y�@�I�vtv��B�I
��Pk�^f@��uK�e�~�ge"�{�v��bCPv��� =��_��>v��Yk8*��-M�]��g�{�Ӳ��<�K�G�Υ�=Č�T W-C֚4�:)��ŧ�%#���4�je�wR�:{uL���,β�s�0�
ǖR�\R�Gv�-ΓH*k��D���Y���N����Z���\�uǝL�e�U[q]k\��o�b]���ѽ�����dA_�@t�1k��u�C!��c�jM�)��gu,/�D���m
4Fw=��خ(���C�1[���ޓא>h�˯c�/��X��P���b�,V���Mޚ�^����H���+d�����)zՆƏ3<X�$���߶(:;�y1�0�m�깋�w��aҸ�����p7�+��qb�r��I���
����������M�=�aѿJ�+Ҳ�x��������>٨������}�+��P��9���m#�m]<t�ޝ��q���Ӑ��#9fC~�P^0*���V��MfOU�&�j�g��hXP��e/f��_�UZ]��jq� �#g�R�%���.N����l�Pp����*ޞ�~���6�g�� ��:����nǼ��Y�m�1y�iA*I�1��;KH��6m���,�Rr9H4/����f�T[df�ʵ��L���ɪ�fv�.?=�_$;�?o<�#<Ib���8��~�k�ث��7��u;9*\���x�R���>;����*�o�־��N��n7���L_p��	A�Ga�sU��e���4���W~b}D�Ι%xAohf#�-1��s1A#9*���׳ʑg˲L���E��9�|]UШ���I/@����v���O�J������S�44*_����*X�P��Lݫ=�J�>?�u��:.Y�Ky���\�YP�s�/�>D�`��\�۵D��=���T�|_���x*��5�Sb�s�� S���w {�ޭ�_�*�T�7P�~��tN�*�V)Tk��k)��tLL~��7��5Rn_�e�C�ê�D�mP�轆�C^%x��z@���d�©�ks�����X�6ߊ�peC�gS�����زu�f��F$:���v`����/~n��j�EH�6��$�!��:��{��y��F�#Uh�l��ڐ��mf=Cwu$̩?���T�2T�6<8L5l~����Z>Lִ��<�bT�l(��ԡ�o�G܇<{��V�q<]���z�X|=LSʠ�� �tL��LK��k���Oqpf*C)Ļ�{��~�G���/	wd�߳�º�z�*���4����"!�Gó_1�y���#����:Sg��]zy��)Lz�eB��ZO�n�����O�l�xʂ��q�e�t��m@�[	�41!�d�fo�7EX��y��e�9�CC���
3u���!7`K�>Uy���JH��uB���;cY����x����R��A�y��ۛݳ���u��$�)(��ǅ*����\��z'3��5p��iIR��8�N��6j^���;u�5�l��:�]��d`��kڴR�Z<�q�+Y��Z�(N���X��YqEӋ���ɷ�'K2vԀ#)v��9���=��r��&7����{���ͼ*"�O��9�q���ج_���h���)UcU�j���D�����ᙙ��R{�ܭ��r��P�B�q*��C�XC�㬽;g�*d�}��+��z�T^"CO��k��Z��Y<�8d��u{Q�;�ݝ��'=�Z��y~zv,0�8{
r���g� t�EŹ��YUCDSUJ�`�*SQ}C�f���&:!�p�S�͏n�*C��>� �]o�ْ�TZ��^*rcu��^s�;���A=/��0.�C[�Y\xW +��7HU#�ٿg��`��]����N�k��"4�0p��4xtWӽ�� W�Ű�3O��*��t��b�gA����~�C�E};v/^.P%�b�G5�[怤�F��:Gx��EU�vi�U��tؼ>�*y��.�������`�FQ�R��J���9��aD��J9j�۩�v6Q��Ss;��#{�y��6�0��cPj/6P�./x_���cg_�<�D���bM��R�){@�,�x�"�!��w��w����+��WB�� 
%^ 7�0z�2< ueC^���3��?tUf�DAࡑ{��u��-S[�S*�Y�y��F����.���e� ~�!��ł8h���*�y�&g{���oX��U}q�X���p}�q~T�$�9���9g�5��|=^���YC���5��Cu[C֬����Kb��R,3�Fz��{�N���D��-5ۊO���.�`�����w[��͒�z2E80�C�5��߈ z�/��-;�4Q�by�W�OW,�,*8��'�&��E'��ژ������0L{]=8,,�;�6r"O8/f8�8Oc���%�o�Y�T��p��^ڝi��Ȯ�h�R��7B5�/l���T:�U�s��3B�ja�fXGMX��o�:F�u�S� �9O:�vܬ�X���!���TM��{J�-1PJ��Wq����KN<��5N��3L;������
��:��xM�aѻt�gV�twg�X�z���^��^��̆����2�U(U���]ߊ���<<HB��GG��Ԫ
W�{PMV�S�KSrz��m�I~9J}�$�Z����-2�υ1�yV;\+kl!"l����z~Ylo���?r�!x.I��X��q.��9�#��W�j�m���9Ǩ�<K��%����۱�����5)���^�I��D�_/���c���zT�\fMzjI�;�.�ϟ���]������]yUY���J�.���%5*���:�dޏ)��FH�0�ե�b�V$�@�z7p
��Mo��OH�=^��:�iexVk�J�L;6;L�q�e!Ay�~��� �u�(^^��˭����/��^���^3KO��m{��:�,�]�x�(���]��T�Q�����ڱ���;	�{��Zq��Řҥ�w+Y��2rP������o�j��u�.��(H�;�se�����E&6�RZ����V����|�){F�����3o�F�̽�©�J�6ہ�
3Sp�.�r��A3;^Lm��bl�t.�i��.�XW;��ˁQ���=�R0��b�i	�E�벗h�������W�O�V���#����iA�g"g9�Y����ƌw�w�8�4�x ��(��s9	,��  �4s&N����Y��ٱU�t*3��䚾J7-=�}[�2>2�����[��Y�4��=zx����4Www
E�U_��~����Y�t�S�ʜ�0�� ��C�3�7�6*��A˂�����V�df������2���(s���:ұe��ɳi��e�j��Wl�;�l���V��܄�               7P��De��n>X4���N%BWp�]��]ӹIt�4�h�ʻm\b��c��fK$,���Z"�*�����h���mXP�{K��1�MmZKH�ҊF����xO�m&q����捉.=Y6.��`[���=��Y}Ӛld����f&t܊���0��,e�t��x�Ž��@�W�%�BL���ݔ`s�gX�ک���	�G�ID��Wswz��o9�5uH�^6��)��x�aW�-�Ҏ��Y�q� :�RvժT�oIr��#	J��Z���r�>�J�3F
�e:�I����{��)�>M�̈?g 2����h��i��U�\<t�B��Ck��� t��mĤ�u�Zҍ�h�`���3��X{���To�$�cr�F��q'Br��XΕeQĻ4
��Pb�wYl)5סٻ�36Sp=O�|R_JˋK�k�h���v 'J&ܧ�';﮺�z�]�AMVT����E14PR�R3AC�"����*B�l0�����u��(��*��(*$��JI�(* �*M�"&$���
�2KY�DA�,��U u&T�LIV�r���
i���(`�)�i(h*���
)"����"����
�����������#���ALM5E�R�sdR-%)o�91 QLH�1I@SCHR��M�̭
SAML�1?G�?D�����=N�ꆱ���c�����C5���F�6���������!)���5.?�F���x����f��C�u��5�^)�2��.�+0:�(i|(�MY���xquU�}'2���P��l������^�.���\6<�f���Tzv�b�Z�͋�.ܼ*��X�Q��f�i�4fkG�OI��Դ���h\b���O6�V�{����0�T�d����<ə^��âpy�x'�;0wx|*a��O-�/B�>��oc�	����B&Y�G��:��]�Fq�g�9��v�E~��0e��Wj�=8I'M%�u��������>�9��걺��=��A�����[}�꠩@4i'ڴR�\}ub��}�\���c�=����a�Ҵ�����ȑ�
Ӷrt�xТ��L�UX��I��q�dj�͵`׎�q�A6������KZ4n%uw-Jĉ��2M ��t�]2��WIɸڴ�oY�퓌�ݧ(/��b�3���޷���5�y�u5,d�.N��3zy�ϣ<O�IA^V�O�ҦE�oF��J&�~�v����N��5������$���-|CK��,��m'���h
�d��������m_���7�-ݯݾ��xZ��J��Uk��!U��?\%����P�,d��]ċ�Uc&��-sB���W���i��7��ǹ����,�=(��<e��^�C�1�˥�)���
)zs�y�Q�z�yO������P���WG�f�b�Bd�/����7&I�}ȑ�S/��P���([\�B�.:�j�y`�co�2��9�y4ф�UZ��值T���د�F��Nf��<5E����rXE��V�[��WH�]T�Ox���%V��h�V��͞��u��J�S���9^>�_9�x1D�U������O��n�]W�*��8��������cc�B�bd
�-��Eͥ���1�ϥ�I���J���Zlw2jl��2���#kf k�8w0�0k8$�@x/{e�'�Z��Q��-�+����7�^~U���t)�v�+v�u8.�hR�ƽ��ӹ%��S� ����}��
��������:�j�wu]���$�<q yz�	n)��A;�i�_nkKA�r����$���ֱ��@��C%�HU�kK}2��`B߈�3�%���=���k}� x����K��Z�95V�0����{P��G�y�=������KT�KZ$��4-%�0y%����À�����{�4nd)�����D�O��Wĕ ��;e����t�ݷhT���jU����Q]fE����\~'O�.��,�� +�P���y[��w�J,�����/ʀS�Y���k�����^�Z�����6�h��@�;7�x��g�K�)4E���j�6?E���y�5���C����v5��j�STR�B65(�y�80-����o'ym���X�n��Ι�	[�9V���p�s4���.U�̃��s���xm��zi����1��珅֐ �l��:�x����+6�Gﭿg(̙�bz'x)�8}3�_н9QnV2Ƀ+��B
F�h�F�W�O
�0�2!^��o�n�b���G�նj�n�9�S㇕F�W�L�j�V���"\o�^��R׉%?E�[L~U��b��`�{�We>K�����^��/��m�������P�/��m��[@5��==۽���643�[_Fz��%�Vd.���ӵ�,	u�Ks�Sz{ze�3��&0T=�h��~lu�PR��Ob��.�h���#����'DW����Р�� �vt��kOg��is��L���H�	���>	�3��\*�yWWF��
���Z���&�ԕ�K�{���].�઴�x1��Aб�v#h��iXy��F����X��m&4b٣i���Z�����JlR��.rv�Vu��;v0r�rc��}m�,m�c�/\��-lQ�vt�������Γ'n~���=���nH_/�x�O>|<���&]@�C w�y���#�	q�N��;�؎� ���D�qR����-������a\����� RV��^ƶ�"LZ�A��Ͳ=��7�v`�}�GK��:��>U�^e�%u�>7���e"����P�N�5[?W���>S���[k�TW�y}[Zn�D�2����0h�;C�L�:z��+�	P������z��
~��s�.�5��E�D��
Zea�f�3b�˃��~��Q�R�g����~\�P�*�!�����rf�
�s���B%�N���o��t����E�<N���p�Sp���6z�C$�$͙[s<�*٣��2y��sX�x:o��t��}X����~Tڀ	���`�]�b����$FfV*E��/۫|��x�Ԉ;x��:�7��:���v�|�Mۨf�v;�N��{��A	/]vwQ��M�#��=�$�����~P��.��&��{���3�B�6�0�)éw���S1�G��3�N��&I��'3o��;�狄Z�9P#�a�ZK����o�`�������睔n��=�eF�k��0Y���K����h�<��Ϫ/ָ��97K����gX�p^�n��S>�ޞ���7�S��ޝ�,�$����ʛzN��`erٱ=�`;޴�q�fU{u�b�ln�!��U��v��u�D�ycp��>x}uV��������w���ӝp�V%<S��@��K#��㣓�[|f�a0�]tP�R���A�;7:�����-�굼_�����p쉖7o�k�WMB��=��
l��ӷu���Pb�ޕ֋�WsEn=�xn&G:�G����G�������?|�jq�j�VSƣ�7��o)a�V�����d��z̓&�&=�_�Gq��W����ѣc�y���V����迚��s� ���s�`�v�$`�9�\���Y�^-�܏z{�m��sy�~3i�O�d*�ɿ���:޾���~	�b�j���%�����]e^��͞sz�<<�ו�m{��o-���Y��,�8mt�ӷ������_!����»��z�������|�3��[tp4w���OÕ;��0`�Yv/��~oӽW����e�eZ�����
B�^WDtС^<&��ٺ��c�(ثjM6)ѭ�4�go����v#��s1��rh����mN�@�ZP��us!���%8U�1���Yc����-3�?{(�|rx�X�r\u0��g�����@k������x�Z�8E���X��-�3=P[�Q_j�P��#��`EDs�'i�7~�ڋ��O{��W�q�7\o�YJs5*uܲ���{n^�{;��>��_�0����:�ך����]����;��H�=e���B�m�x��:�2H�'���X���Ш��>�u��uG�g��x���E�"j3�%��\+�u�̞���@�"�x��r:��M��Sя��\s��6�g�Բ
�������7>��i��:HƲ�Ī-�vi���ؐ��;-�2�W����lT�CsO�k7^M,1���u�N\̵�9Tl��)`8B�&=���v��Jۦ:�[S{F����Mo155Ә�)�ӫ�9G�Zǝ7ѿ������s�mҿ5�wѿ�1�����ZfP:]�2j(_�%���mt���|�=�'L�O�6++ەSf�i׀{����+2o!0���#w�Ѭ}��%e+�G)v+e�����%�l�~��Z�UHjݿ�(|ĽUY76<�p�*�l���H={^4�{�����{SF�a�^R�g����lg���^�I�y@2����:|�:�M�M�哚]uM-}*��g�����}H�C���,�P�6K�xs��KU�x��*�VfOyn��^^��]G'5cxf��fOl>f�^�<��}�e��>PbD\kA[�A̴��ZE���Ƴ�@��Pu�2�WВ_xW��+��Io&[P2�����0�yQ�"�B��}c���n���n
͕6P�_(���|➽�����ե��k�&�b�ʍ��[���6o/92�e����ڕ��Fq\���B|nj����i?�N��~��ǉW�N7�V�^���J�u2�������E�9��S��##���\�۬w�u83k�B��*_:r bu���4wc��=�#�^�/9T���.J�� ��}��>N
��9�V��[�tF�#�B��P�ǆ��G�_����*�ۚ����}J����d^`��m�^�s�R�[[��+1�z�3��!�hqMH{}S�GF 2��Qq�rUۮ����{kU��X`�Z������~���w7q-L9D�H]q�u��ږL�y啶��S,лWN�"���0𶙛1�lB��r��}A��5E Fnn�tMD┳7e��\�1�m.e�T��dY�1�h���[�d-��ʲ�)�h5�,*��{��Ų[u�`�0qዀ�OK:o�e#y;{a��4А;w��w�2vousw%��M�N*��o( W\ެ�VC��B1B�n��4;Q���0=D��?n^�$Cש��m@)�^}�9��n�jYd�Q�F��P�?��������3lP����K$jnW;i^˼G �tmc��+F�d��ܒ���p"�Ư, �
gnܼ��j�[��j��j6��(D��:����4K���I�JfǝO���*�es�ڵkZ�� s��Ρ̫z+)����Ov��T����#s(,R7F��\���w4)@��<9^k���F�2��>��,�y.�L�����X��
�Nι�ێ�s7e�OvQ�'APg!�M0�m|]u�                 f�w�%*W�%���-n;��e�^��]wf%�-f͜��R�u��ݿ�OB2MÐ	��\�/|yC�j"�7wut���;5Z
Y�
f\%� �v4�rn�x�f�Ԧ���u��hH�-��x����U�ڲ.V�aA��ү�k��ܦ͛aCi�k�%;�]��)q%��>�׷a�v����	4@���n֫Yڲ�o�h�`v����ws�Ğ��0��^ `��hT�h]-[���+�P�UM�D�s��bݸS�^kǳ����c���KKB�����<�TU;Ҏ�ռyY�fRj-+�{��,>��%�A�i�1�0�b�6,�9H�j��է¨i e���@�Q��r���rdji�R�����! NĺS��l��ͻ���{�	�p��"��"?ц�ާ�mzo���G�V҂�ƕ�Co�Fj�jp�ZA��p[�)�4�N+���몦����� ��hh��3 8��5%>C��Rǘ--	E4:����2\�*T�Ba:� �i2L��*�)(
�@Ԛ���Y�4-!��EBR��� �h���<�>Z��\�ZH�9�®$�^l���)
WP�B4/ꪠ3SV;Ժ�9aru�+D96��ׁo*!�ÁG0jDU͹W1Q�R�n��mF��L>�1�ݛW�i�{|��K �y��򭈹����F8䓶{t�{��z����4�Xq�z��F�ڰ�����U�U�\�`s��B}[n���՜�F[�6��O���*��m�rsP�l�Ǽ��^��{o[E�xp���Au�6�❔�׽x�	 �����Um��gx�.�+�^ï磽B�9�x��Z����ޗ~���e]T�z�գW� w�v+�|��e�U8w�<��v4���b!�Gэ�	m]�w��g�W7y�{���M�%b��mT��n�V8�u�J���Q���Mg�M�2������L�e*U���ѻ{f�ͥ���
Ҷ^�蘥Z�yG��̶���+���L��.�cF=3�>��&�]�rb����2]6W��OLCK�j����"��������3�vi���k̫��kڈ�]�ݤg���<Z�7�����	u�_�:�E_<���'���g�H������N:�ι�F�3�g�V传�<��M��o-re�4c���r˰U���3`�����G	��{�j�ӯ�ڟ(��_ŅL��q|��]��Y�^q�.�3p�FyV����.�x�<��{��ܢ�x���J*�?*}G`���x'y����-���B����0��#����_�i7)�%%�R��Y͉�	o����[�I忏G�v�]�2�Kw�^��q93/3K�'��']�!��" ��s�� �V/�Md�p��{n�a@�+����z�
���˦����]#ܙ��9�nu�����ev̝��\]��U*Ӯ=�fWQ��ݪ�,� ��y7�����ܜ��rEG�zf�<s����,re����{a�Y�6#��9�[�\+�u�2^�Ug6�fM��9��C�䧱�տs��$�H����sX>o�s���
�;��,S�]�O&���'"=���*������/|}�l}���כ���[[��\�!L�E}<�9���~ȭ�����|�9}Q��|r�����l^��K�B���������V�{�塏��ȸVT|�U˘ÎF�I铄��n�x�?f��:?܏e��\�j<��}�E�S9�9[ɤ���]�ʳy����]��1ܽ�$P��^=�M�YV���h��n��Ķb�g^R��uC�����\·��7j+�јVЕ�sx����ݞ�1�»&ڭtGܶ8��^x.�C�����ꦮ_C�3�U];u�6z� ����W��U\���AI�Ҫٴ�ʱ���z�`T���Njt�78�=�\۫�5�)d���󸦰����u����Eۯ߲�9���6��2y��������4�4����E���j�O{ݰ��Zq�N�mzhO�K
���Ow���*ؖ{� x]�ZM�ʼ�{�S~ͨ����q8S^��	���u[^>ev��ng\%�7<M�=���Nf�Ge�K�y.�6#�&�޼��E��ۧNN��bBdg{�x�<���w0��B����2�(�7���]��D^x��0冲�|Ӵ�
�W}��}��]=�w<E�@�ů��#�J�R<kT��c�&fgF�{m�jSHf1~�!;$L���L����e^�vW��c�UQ,�Op�i�ₑֆ27��vvN�y��}��B'�_����n��^qt}��\ů�̦�6�����V"����ѭK�W-��g����+H��z 2��Qqw����~(���t�o�c�F~l�>�F������hIt��O'��?Z��b� �Us�׶�x�ܖ���⾏������v+���Sܧ]�L���;X�]��X�B+��r����^��U����	˚y�O�E^�k}�8oz��Wɺ���e7s���Bj=x&������^�-�Jɴ(��^s�Y�>�W�<Tܮ�g�n<�0AkD�M4G�i���`��Ӝ;8�yQ�s��M�1�ƚ���(�B�N}W�#�zOA���у,f��5�$��"��-CZ1*�O�|7�ǂ��mRF&��AN�
�GCS�\��%F�>+�N��p�ǜ���{rU?*���u��tz)W¸��=/�\%��L��t�代��m�ZjI=�]5��-�j���$�#�zE/nk����:�d�i���ס�t�y�W�\5]W�����A�*�Ezy�}���Ϩ+Ut���$�{�˿�Ʈ�;lV:�l�G��xG��b��/��O3�b�����̠Sx��*��~r�a>���Y�6f;]]�N�ڟ(��\�f�Ԯ�=����S���j��=���]���^��u��$�z2�T)~k���ʹ�7YVY��~��tq��kd��;�q���*Rkvv�=ܱ�[�Df.��]���k�֣�%��;}��E����^	�m.���:��ҎdϽ�϶PN��%*Tf��Wrwr��n�c�R��몊�_�mݪ����w\��ܛv36k^2r�VПd�z+(�3���Uɸ���,u�y̝���3UnfJo$�S��kѯW^7�y��+�i��9�!�ݯ��G��*6������ڽ���g:�J���ƕǓ%��\���ް+����5���]���_�o�=��ux��	��\�k}>ډ�|�&����5��7�e�*	{:�{�k�Q�N��ι���\{U[�~j&��Z��������Z��{�7;��E����!��-��2d����(���P�V�i��#Y�U�r�������	E�"�,��B}���*���AA��y00��'K6ܢ��d3f���֔Ӛ]�^�TM�y�(;ykp�z�%�8�Jm>��9Tz��g�zֱVW����s^�%n=�2�D`��<��O�y
��m��&w�C�����蛞�m�U���2����tv��#O�9���r�^�/e��z��ظk�l��E��4'�p�=�,��׌�Uu�ϳ|J��1�L�=�Z�!9�]uM,��Uv���a_oo��7�s۪����$�Y�Xu��w�T�������!��ڬ�Ϸή��99���3ko.1iu�E�v�[+&u���q֪�<d^�}ή��I�U�n����#�����wӕn�ɣ�,�9�
y�Mj��Y���K�`�޳��ޖNܳo�+Ż���i#e_����I��otwKm.
?�$1��y��v!�2jR���kR	��m���<�7����h�o3��^��ܸH�]�p>7�5���'�az�>_WL�'?^����Zޏ��?��\��c��mdқY�<�nYǣ3�c���\��4���' ~T�~������������)56Q����� {�/xq��.�����]�)��5]:��r��}7{�fH�f3���O���Wk/wVo��zW������Yu��:�zI�ԚD[���\s�(�\oMx����w�A��\���5	�G���}D�v�Gޝ��DOu_z�UM��}vje�Aró�;M�h��k�ϓ���c.�U%�Eְ窝,�{)�k.�y�݆��}�-�7,�+^�d&�Z����.]]�[(���I���>�8;qbon��5�^�%���03�g�oe��� Q3{�M`��u#�<�hk`���+�^�:���}�Ds��B}չ��a���p��*i�m�OZ&���WeC�ox�dA���^,^x�CU;*'F�������Y�4�o'3�bL�k���{.�g�89|�hK
��kbTy7*����b��+��ڧ>�*�'��==u�:��~15��_'�U�[y֓��[��חy>��W6;��(�ns��\bt���d��=Q��ފ�L�;�MϱuD�/ݑ�Ӄ��Mq�TaKMƛΚj���.{�*3�Ƿ3����TZ�>ϫ �=��oO�˭w{A�ke'��U�ٳ?z�r�*����������T�QC�%���%�����TQ��j`����0�/��'�d��=�SF�bkGZu�pl�&��A�Ӱ����xGq�X���
�m�
�h�Q@�P" D�=����A��nbbF��'�Ħ|`�������9|�q�qs����ڔQDŎ�W2=�E��m����S��O�6��3�<��}{i�œ[�)���<���_�����~c�Z4���;��� *"�O?��|���{�� !y@� DO�TEDO����Rb��������������ˀ%?������A��O�?��}��O����TQ��u?\�}'�q,D'����?BH��tlBr�x�[��K�?��sR��m�3�5²o��G���$�|�I��H��G�C�o��Ҋ(��O>���F��ۂ#eQa��'�l�v��J�8���>F�f�A��?�\�	�<	���l|�*(��^���0�������}&� ~�̣���j��~������� �������!����������ѵ�ޜ��G�3���&���φ�������O����}遼`��1�<4>	�br���y�����>�ܟ���滣���'���|�_
����w�Zr}'ࢊ"}}��]}��$����ף��:���oJa9���U$�'�E?�?��;s�$�O�Лv�H�|l/_�GF������hTD�8��AI>	�E������� Dės �yT���8]�����h�I8�Y��ʏ�#)�x���BK�'o o��Ӥ���`��TQ�A�����z����(����~�����`���Ё����� �<�����?��~jh�p}K�m��~������C�|�d��Q��J���������Q�?��|_�L����N���(�&/�q��ӣ�������>a�b~?���)���t|����>)� t�ʄ� ���cAi_��>D&���@�O�������'�w�_��:�r=��2�}����ED�������	��:����,��nI��)�}�|�h���d�I�a���}]���軪}���H��'���?WO�&����;���_���7��}�0Q��>���������<&��	���oο-!�����%1����O���Gߛ���w$S�		�i1 