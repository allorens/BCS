BZh91AY&SYz���߀`q���#� ����b �    `                                     P   �  (       (   (   �      � 
    (    ��H �"R*�TU ��T �J��Q"�%"
I@ I �T$�S�$�E �"���& 
(�n)JHR��P�Ut y�P�n�P���7XtDY��'t���tS�ʨd
w]�B�\�w@�E��Eb�� ���Q�Z$��ʽ����)>��̪UIUǼJ��/iT�mcj��)U��"W��yd �=� M����@d d9 �P @}�� T��*
�U�EQ@�S��  �� �����(�uD�� �@�t+�� <�'@	�xP/ =7X��8�� P  �  s� ��w� <{���� ����{������f� �Ǫ*< T ��:� .�� � 4 (>   ;�� �����I!k � 6�� 7X@9 1�{� /w����l�/@;�������y�.�
 dr��`�   h�   p>� |�v 9p褬 �� �@n��v 90t��G ��� � ��@  � �=�R� 	**����| mc��� dd �@ -��@d�:C���:�� �`   �  {@� �JX �@����� 3u*�p �@70�� ��  @_  �*U�@����HA�lx���� �s� �ꪩ8 �@7`� �n��"L 28�r� (� �   y:�à	å%p��7`t@1� 9�Q%\ Dr �`: �� �      S�JR��ha4�@f�i���"��	)*� i� �   D�2�T�OUOH � 4   l�@)JF�0L2h�a�@��JJ�OT��bd2`��L4�� ґ�4���4ad�B}�/�����K��yq@vO�9]xA�o�w}�s��À�� �(�
��*|�Q_�U���?��G������9?����|�?�
����r��vUAE~��L�D��((+�������_�� �,���dّ�Ȉ��*~,*�L�����*~L(&� �E�DFd@tʊi���QL �2"�A� ��AL.� ^X 0*L"�4��dM2��L��P�0�L��"i�4Țe0n�a2'�	�x�'��7�!�"x��2&�SL)�D�l.�0�̡�� �4�n��t�:d]0� ��,����������������c�L.�CL�� �+�WL/��fL��0�`2�at��;m2�evet���#�L��CL�L�]2:awet���+�L/i��+�L��XL.�0�at��!�L��0�dydt���#� �0:a2�at���4�$�i�@�t�*i��
��PCL�,��2�e 4���":dQ4Ȉi� �*�PCL��L*�T2����
!�L���P0�aP4� x��i�eCL ��0"`P4 i� � ��TL"�L �(��CL���M0�eP4ʠi��
l aT2 �0��=�&N�׃�@��[��/Y?S�g��E�U��\�i/{�G{��ĭ �M�IM�ws�R�m���W{�Wq��C��B�V�cw/�:�Eh�>���u�8'6b�8�����cb�E�R��u���k.�@W/k&�Y׬�����;���U����P�H�԰��6���R�֎ʇ&�x�Cw�����f��;DZ�iA���ٙ0j�@0��F�:��.G�7�e΅�#�ak^u����'�wM�U��&N��K���9��l�-�ϊ��F�!`ƭ'���\G��{�v��]XNL}�	^��Z�{��/���M����*C���!�i�3�	o��a��	�8�DFk�.+��
�Q����AF�[r�T�x:܍��q�㽄�D:nLM�k�ػ��9y�<��g�kO;��რ�׽F�۳����4���%���M)�=f� 4�c\�2�����)�����{���;�qc�J\�[����x<�F'.���uA���BТ �����xt�~���"�ˋc(�ńZXرi��nދ`�X���)�G>�w(��c�:��]�R�{�pL =V��ai�r	���Iy6%�;IX��e��7�t�5�`���|�=L��)��.�"��7��j�.~�����M��1�&��.hܷ{L� ��W�q�GY`�/kF�m���8�)B޳�B kgVǦ�r��'�n_�,�-����{9NӖC��0wJs���.wu��e�]�-4(����	��:M���t�Io�J桮Y�5��s��p�}��^���o=�G8{n� ����3R����8�o=m���e:�l���Ì7��qv�BM�%H6���U��{�a���`�b��n�p�sZ��w��~/����wu3$oP53f��w��0ݘ͏b�a�ns����X�jǗrJ�7���3:��VH�-bVgM�`��c�ZZ8@2J�k��YQ��S��/;���b�иlu���d�8�S@+�-�-�f��C�f٢��y`�U�o��9�74�Ԗ�� g%��rx_���'-j�J��p��~������vj/4��ob��ɕP��^��GX�4�fvꌦ[��˭9L���z;]F#~ߦP���$*�D�CgMɶV��Y
�L�gv����i�����v��55h��N��jY��vv���1�FL�3��%&�H��CKx�V<�	�2�ɋC΂�un��4�2���G��W)�\a��ddl�ȹ�{�:a�0)�S`���\Oi䓙	�[f�_�C"�z���[��u�-sph�8�����x���y��t(�Z�0[���]� ����.���9ɔۮsnd
$�,w��EÚճm7Łp�	�K՝�xv=�]v�!߻'����ʩ��D�k��,�e:�F���i��i!�wPΘ���)7�ݎRk�wI�۴l����B���<3
��zF������,1Q�d�ݰ��x�h<�UE�������͈OT���ۛ�ܣ6�R�Q)��ߴ��|��z����]y�nvq&>ȣ��	��-�3�1��.z��b�
Ju��� �"+Op/��<����p���ep�;��/�@�4���!Y�2ع�n��[ܣh̹Ni���#P�Λ4�lY�gG����Ɛ �Vt��nc�)����%����&.|q����%}�GExY����p�ZH�k�F¥�!�>]^��f���\�o%�N����뉚�<��:� U	���n"����X�A�=���#]rlrؘ-��_�`�ʄ�yRf��2�,'���U7Ǹj�Z��M�\6�8��xV����sx�;�]Y.���p�N��qݛ��q�7n+�5l�B�ض�
�O�[9��"S��%�״��&�"��}� �f����f��7F�Gu]CE�7ZE$�SB��X�&MfZx
G9I�{� �&��+H�l��p�,��@�+B�LF����6��6�@�9:L���Pc�OgP(��|y�ǒ[/w	����[�p��ś�4� h�#/����	@3{9v����ΈÌ�(v���p���Ի���	 ��Szg�8I=��Wȍ,G7F�ޭX��ٷ�����ލ+8u��h�1���q���0�Ӽ�ϖ��8��閍�Z^��w��l&j����n7�Ni'�]�lM1>F%��Θ6[�N}�ۧ�p���M
��8}w$�nP���K�-��!�����f��v�����&��_>N�G90u�Y�1�l�/ F攷X[m�Y��F(�g����҆9ף�n�X��W�k鄝ׇ:�S�]��s�t�iְ�v��݇V-���8�N߈�{5�%]죗E��6.<T���T�w������c�9����>�y����1�k6������E�,hیҾ��R7�=5��l,>8�����!a���� ry8�wJ:n�x�{����9χ
�ʙ��������;�i19[h���uz��X�yiԬ��/��ɨqx=�9�5����[L͜L�a����}�����t�"<5�����C��N�j�;f��M�O}���p�)r$�v�#; � �t�Ì�W{:k�tKE6:Q���ͳ��k9t�{�|�v�}���;s�����)Z�q��a�I�n#�A�X�&O�ya]��`\��/n9�8��"�'p��4e�igiz�ǋu;��ޝ�v���/u}���4M K؟��S鳆8OvV�A� ��A���&��Qb�yP�Ɍ��8���|����$��Ԧ��^p�����f�Br,�Z���F��V���r�{�	�Y����ya}˝����R6�/��f�Ԙ�U�t�5Ll��;����FV�*o�����$׻7/9U%���y��VyY�]ʽ�n'�	ӣy��:�A8�6rfś 0bٹrYz�i��f�}P�LGt�_�G0˻�7eL�0cPn�<��\6t��QmZ�`�<7�&,��q-ųT��vj(�$��`�`��Q*�N"�;��Y%�}c�M`��v����߹f�1��ñ���a�#N����n��oVH�<'r�p�u��>�i`��(#j���xz���:�#)����6���`�ww�r�'e)b;^L�&��L����|�h5f��ҙ��!׈-�uW��FG�W�TE�i`B�烏��9l$���uO.���=��Z۽�ݏ��%��憁ѩ�yV,|�m�ۮu�_
V�9�mJ��dy�K�p/(Я�ga�):��~���{刌(�O��|d�&,|>�c@�9"�m<W<�3�&��o�N�}v
��j�^hO+P�N8�N|)ś�G�S����BWyK�{7�1���aZ�p����E��4T��,��V&s�pї9�b���Q4���iǺ��BhŃgn��8��_k�a�{dC��u�2��+6����-��FV(�nL� /��D J���AW؟e�Mgb�6���wsr�z#��%c�&�V[.<@��g7f%/-|d����y.��"���t��c��רl���k�[��Ĭ��аoXSͮ,���ݚ����p��f�I���ۺ#ܹ{[��_��:���"&�Q�@��7��r��cL�n�6=�7��W�_]���	u��'�z������y�����$�6���ym�0�k��Sw���qR����D�g0��sC��7��(��Z�n�򙒑&H�J�����v\a�V�v�|�$�2��~;{
4�d&ۈX���&  �3�N��p�^� '�p��p�����1�1�ؖ�3{6�쫠R�5���Ljea;�&\A�W��̅���W-,�Ep=�V�N�3Ywq)ni�Φ�oe��q��ѷ��<�q
����p��c�:�I�S�$y�O�!�n��'` Ǻ�Z�Ud�]�F�yq��N��1�P4Eb��s��s��݋��	���u�3M����4��/�	�x�;�E�jų�����)�.�	]{9����/��Fm�����v��Ř��/�,����ɶmFc�j���v�g
au�Û��c��,E�wg'ژ���;Q� ��w�V+	J6sf�W� 4��M	��|�ۅ��N����j�?/^͏�ǖ�:w)ے>�guݣ�99���p�#7ot�R�-�u�a��'5�7O��J�
�@�7#��ZD����oL�0��=����hQ�0Z�sۗN�LYн�)=ygqKs��t5���=��ۛ�ts>��;͊�A��>=�MUŰnh�D�H���ֹtC8��C�����k,):�8��©��%C�����A�:�[Җ1�ج\r�x0�Q+�i5��s�7TZ�p3V���ͣ�LYt�f�z'	k����
o�r�ړ�X��cIh�!��=n�܍%��V/qP���뒺0�A��HR���C�E9f�Ȝ��7�3�owl�/�-�[I���W4d�����HV��9���H���5�jH��]5w,�I:Βls"WI�Ơ�y��k;���n�5<��Ktt��7l� ���Q��9�b]���u�n,��T�^�Q�8ȕݵ��N��wj��zC��uj�!u,�Y���j�0��`<)�Gn�c"�X�9v�ۡm�	ōwYf���aWeUr���F�n	��٫L��e����.`�vg1ϒꔩ�֬��.�W��˲�ع�p�U�tD�;�Pq�	Jc#p�[Κ�8�{c�m��<��u�;�&���k���&Ѱk*�}yj �Hww�.t-�3e�v�:�v�[����������J^M�
9oM�7Qc�sw!�LX���1��:��J��c���To7 ��Q�F�5�@|���8
����,|h಍���`��ۏVo�pLg^������f��6�D��Clz�fӁ�	�ĬC�	�d��N|ڊ[;=r��I,֞2��X�_u9�����7��ȗ%�e�<nn�)��[�jxZlD� ��Y������1���|X���tvn�+��R�Gcم��*����Z`�;s�7��o �0]��d�rGI�N�3��t��ﶳ��1��;G6d���@���
����	�݉�n��6w;ؗk��|�:aFʡ�6&�I���[�l>S	��ц
�FO=� �ڲS�\�U8z˓��s�*�\.�(�l�aLk<�M�ۉ�&�7n#�v���׆��� 3���]{�2���7:F�7��d�p_��u�7��ǮmGB%�Z�4SE|2Jv��y#ǨӰ�t�CbF��z��pl���;B��6�p�XD�����P�� Z7pA_m��Dü�Y�^����k�p�/@9^c�}���p(2UTڬ�9�n�V�}Iر`�oE�ft�C�.���p�k���֋*!�״�@��?��t��uF�Xb��\|�z�R�Q�mc;7�sW�tє�p��ܹ�p���}�TnW���r|������l�ߦ����R*�#v9p�X��T���H�(0R���jf�b���M�bS:gQ��C�yó�`sf�&^c�:�g�DE3�[h0�ڭ��
ú{��)	�3w�qA�<�F�Z���ݪ�M���R�ɻr�z@*+*X�.��Y�|2�nt�1�}y��ʖ<�wF�1��<��[�I/C`>|��.�������Q�r8(�34��B냹�U
z~��2��U�y���v����Cn+Y��oIս�H��|�n�C��VE�@�< ��5��k���^��\�'I��T�:;'b�1hŶ���]�-����sZ��cW��ʛ����h�������v�!�ˠ�;v�9����k��U7��.?i���&�0�pf���7�f��ˉޯtm�4Y��s��z���i <;�(����-�ݝ�a�UݼC�rf��ᛤ��mu��y��f�@ħ׬%"l*�8䰜:��!n���jǉk{N֬�U٠4q7�wgI��7�莄{w�֜8xv�f�t�=��0���{sq���/Y�7NѠ��a�j��s���q�ϸ�V��}�0wn���/j��G{��I�]B�E<�lɚ�D�tp��Λ�a��qq�����{��i���]rlγue�|8N�ξ2��+���F;w��8��5l�rn����sY����ƞ��{,TL&�l��Ӑp�$���8\��L�slՏddqP2S+7p�j�+;�1Ǒ�؜��G^���ʯA.��v a�W�,�pF.dr�3�E��m�,�L\ֱ��PkhJ�x�F�q���cxۃ�%�|W}F��إ��p����.��GkMIVgr&@\�vv�����-9ٹ8�;M�������	�k����hNB�Ĭ@��7�e��0���	�do���X=��Yt�Y>��:��.������Y�O�v����W�o��xg��{V���5��o��"7J]aJ���IX1����f3a�(���x�OԃV�J�_�)�d��Z�*T�yI��E7Ĳi$�K&��I�Yv��S����©�|�Ө����̧�ZFĳ�S%�����N3���n��t�T(�
�'�|oIFzf��;�i��e?��-�`�g��<l'N���X��3�X�l��Y:R=�R�V�K���"��pL4&B�06�� c$й�e���0�=��G���;}�i�7����>�iO�C T�2P�T)(r$��D��U)C%Ar �C!G%�Q�D(E(A � � �UG%�J��D�JQ@��G%�B�hT2�!A�%�)@�L�
V�%P2(P ��U�V�ZPE�Eh��A���2 �ZPF�Eh)EJ�E��iT�B��L��T
Dh��G$Q�A�R�Q�QiDiP�J��B�) hTC  �R�@�Q� )D�i�rU�R��J�D ���'�{�}�-��(Ch.qx�����4&�u�'�4��(o�{�=Af�o0m�#�om)��x[ط���<E ٍ��[��-	�q~�E�>g�}��������?��4� ��o��~�����B��)�?bTL�,���Z���P�{����~�p��=�̈́�-�}ґQ��=7�ݹ�l���7�Ɲ�.Ql\t��1��U�T"n�x�]^���p��k�L��:���Oz���>Y�Vl���n��Cد�l��gpp��(�C��y^���2W�W�ݢ*��v������R�..��o�>�=�
y���3�Uѝ��4GӸ$lb���{ύ3�p��)׷�F��.ަ��h~;�-��=��=zg{����ou�]�P�uC�~^�H�i����v�//�G'�C���+���Y�SQ}�/t�t.�xA�8�a~iE��c��cX�۳�=x�~���Q������Z���n�vm���q/�Sڽ�酏sM�V��K��{KR��6Ê]�]�}�6]{��V�4�؛��]ӗd#�fy�y�����&�<�����"���{�/k� G��!{��.��r9;K;;�q��������;w�����W���;(1_7���C1a��C-��3مūa�8�SSf0M�����ڮ$���Q����s��	��]��]=�*�R����؏�䗊�x����Y�;ݝ<f3�o�f��fq^]�O,��.c�=Ҋ]�xl9�8�m�=aX�]_����SN����4o�>�b�~�g�߬�#�����y��X}��\9�h��;C����a��qU��S�� ��B,�Oކ��w;=��o�{�ջ+������=��?w�xw�p��xrһ�n�}����t�����K��[��x�3�y�M�Z.�4������}懘��^�s+������:�W��ޝ��6�%ǒw�#�r��������1I6�xa6G3����nZ�������(k5s�/=������\ؔ>�K�$"��kK�z�J�����P3�m�s��\�u����ƌ��b�4��N���cY�sƱ�_Q���{8A�;�.��϶�L��OE�}�О�<���4{u�x�{�^{�NZS>����j���?a�N���ۛhӞ�Ρ<�����z����7��U�{��]ڋ��=��7=�Rr��#������{�O��7��}�$y��}3�<6���w{y���	�Q�ל���=��\���P�A�ɾ��Om]]ԣ2�,���}���g��>��N+[��\|���JP������n�7W2t��I��i�Gy�)��ox �uoQH��Dv�9k� ��q��yF�f��<�vN�i�j\^�z�����#	��%UDk�����މ������J��>׻�F�G8Na�h���7��$�	��'���C�Ѣ�ы�&1"�u+��zC�O��>�b��w��yh��svm֢ds�~w�nü���3��N�0e7�@7�>��i��>���3~�ya>�x]'�|���������(���sCZߥ����t�~VZ����H���,c�ac6gh�ƫ��噷�{���kY���O ��������uLԻ޿nے>��˽��݆�����g��v��!I�ƴ���\M�ol|�2td����54�i!
}��o���x���{�C�l�J���'��x���	a�)�Ʋ}�6+r�HT]ὓ�2_>#��}��<ץ�{�bґ�w�g�씌��Y��#yV1���ܞ�iX c{��2n�4�]�`�ܳs��g�'o�f��}=@�7f�)]>^~�{�Ubw-���Ǽ:�^���]�ܛ���jVE���\��Wf��='���x0����K��o#� #�f�6f�ٳ8��qto%zWްgn\�L�� �E�>&o(�Y&�h�'<<�s�X5.�9��0M�� 垎�������>�U/��>�^�2�������M�Kzx{�;�o�ֽS�"V
���Z�aX�M�������$��Ԕ+�/X�+���:8�����V�׼@0��W�j�M�}p��� c�ۜ��*͞��p�rw���i^ں{��{�\��7�\�(�:��z��Kk�n*���;KӜ<�^��o;����P�c��/�R��|�^�ߘ��ˍcN����Y��⏞n��_1{$t�ux��"��"~���{�����1�3��'Э�'��*���t�������{�����[=�0q}����<�2��O���'D�b>��xN��pe��O�%5�e��ۡm=���.;{ɵ�.��ϗ��ל��q�>&/x��'�x����v�����|1|<f�c�'��lf֯"�V.l�����aO��=F��ޜ;^x-��� �A��OO=������Gz��)��u�\}Ќ���yM�g+��qM�)��@xW������8�����KN��[�f���;�xz}=�����=�G�F�yo�����c�}���^~�!���'��^����ܧqӸ}�ׄW�ܟ�!;���,�������{���e��rsq�$��z<XWu��DrQ3G�Ut�L��{m~����|��n�`C�������+v�����va�<ԓ~��rp,kx�wͻ۾��YZ^S;݆{=�&*	P'Q���^*
$��v���n{s�{��B"^�JF��֌N�Uˡ�ve���_N�*D������TF\�M���Gx��Z ���(�}�;�`*M|'y.��}�5��u�j��G��ײ�s��KV%�>���s!xogt�t{˕Y}����!2���a��E�݇�Tj�{1�`�fԳNzʆ��k�^�4v�]{L|j����.�q�����)^Z��~#�����v�V���p�����T��7,�lW���Ƿ��A6�=qo/;������}������2k���	��׆�q
Tgx��A'ۑ9���o��>;|g�3B>�ڽ�b=m�����t�T�ۛ������s��_v�����҆�s����V�{׻E�g�����n��ǎӔm�>��O^����ݑy$�D^ˇ;�:��G�ծnv���L��j����&yf�8���e�pO�ǽ�v����>�ǧ_1U��������y���H�}<��b$f�"�'���j��#�Q���佃f�d�*4�g{}F��i~��on�ð�۳4��7ӻJ�û���C2��}����_pd��w#�)����9ЕI�7����}��=�ĽZ�u���s�=������_n"GOXn�y*�Ҋ_��z@3ڽ5t������ 7,9=�}oL�ִN��ݸ{�AOh;�<a�n�t�5˯#[��������{�99�:�����g��R0tg=3G �$VX�����n%)�-�!��ȼV{��;�w��ps��d�f��Q ��	�23{����p���z�q�3�����p��g:�4t����'Ak��J�}�1�?!�=�+�|�8 Λ��m+ٽ��s����2����v�yx��ZL����Gl�>�i������n����Gyy��K-�{�y�e�U�/\�|N��S��Yxg��������Nx�[�#��]�k*�}�y�t�@���{���s�m�vE�l�N�ש�~,Ξ��F�a��_r���Ԩ_�(o��ƙ�}���zE��!�
���q��+��vi��{8v���w��ǯ��z�T��{A9fv�ڗ�Da����ѱ�����כ�"�s�_AR�t�F�y^�޺}�]����v����wi��9��ڼ���/K�<ԥ��9���A����o�]�9ף�VTٹ�x�h��v9Iy��#��6?ke|����w��q���?i�.���,�|���Y�Г�y����+|�9��w�f��������pt��9��e��=����1�_b~�� x�7/o��oo��찃��Gy�[j����g�O<�� u����,���d5�&zk����\�ymk�D^�����8Q�/�`7�w����L��}�p�=�=����m�Q���Nlf��T�7�E��e��Y���׽���d���a'!�PҾ�)�m��r�MP����K9u���nx�(�#��i���k�al��ឋ�^���F@y"xU�Xt�e7��D�yc���<���ﳔ���z%������/9�d��߬V��}���{|ׯ�'�ﵭ��}�������7Z��*gj{OX�p�w�l�b�)�"A�<�?xE��'=�{�|tM/��p�}��n8+�9�ѰҌ���Pqy�q+���;����\>W��o{��M��ڷعGȈ�	��pp]8Y^]Ч�&��j&umM��ty�7�wޏ�-3�L��o��\hQ�a��4�at�V}z#��<ۙ-n�����i�h>��h"{N<���:q���}�ɚB�[/���^����<9���+M��n�������o�.����}��^;۝ٺŖd�g�>�!a�-� �s�|�k�༺g���^Au��L�ɯ>�.����L�:�J6_#3�;Ţ0�}z��3�M+/�����ě>���!�}��5�����j�:��]�\����7u>R�Ke��l����[��xW�,���Vo��V<���R�g</;�r���:Bĉ���i�{��?z,;��s�z���8S��ήKx�qI�p�9WC�C·��|��]G|���v!�f��+�b���w�m[��Àq�~����A�f�A�0`~�Q�V3N3,̉�9�0E�]Xː��B^бxqw��W�<�۳�ǵ�&��	��ؽ�w��qM��>��Y;4����i�̥�C���z����8ћc's�̺���R|���Y���.�̆lYȾ��7�vyO]�S�����O��T�>����"�e��ǆ3�����������vI��t�����RN��ۧ��Z��~ak`b���0�Q����Y1P�n[�◧Ns/<���Տ�G�=EԪ��{�!�ő��E�0��MW�MתU����1�fV�����U�n�&�
 �G����wX}זਊE��÷qj��'�d�����{��T(��\�hEٱ��I��_k��ig^OH֟zAxQ���*��g��ʋ�{�H�Ӽ��v�狣�'�?i3�k9�����4l>���ނ�V��/{ ѫ�ֆA��!U��b��ИP��c`4#>�vq6FT�yo��rQ^�Qs���(��%~[���.�U�v��E͂�D[��b0i��8�9�gj���� ��`��n����M�Ş�$�Gy�z�y�E4f�����y�,p���}��ۮ����:#����RY$�L�&m��Lw�)z�r���4�nI�6������!�ۺ���7����s�[���#�3���T���Y�x��f���ݼ�=4�Sɧ0����{tn T�oѡ�`=ݻ�}&o�xg������/T9yX�٫�>������q���nߏ�>ɉov���ݮ�o��(���n�8y�0��\�{�.i�}��Oa�����ꆆn�f�{���/p�o�S���g&�2���j.�����x헜��.�{�^��"�p��+�zZ�^�ۀ�n��m�s��A}��]�M���7֠^��DZN���>�$���7=��''�b�b�Bc�}��§Q�W�ͭ��/H
��=�N�K:'ʜwuQ�H.=o�awS	w�AuM9���z��h�^�e�7:w�q�;�� �Q�2����N�=�b�}���E�OZ(�~��-�����EC;�K���P���ݮ��N(y�Q�`@�g�ɒg޾`�@�g�w����1z�o��lo���^�wv凗_Zx���;{��ཱི��w�ؙ�E����"d9�ۋ�=[�7s�<�}�Vn.�bȢ]��g���p3�8�W|]��y3����F��:���7���M6װ{�O���p�����L�Mۢoa����r���]h���MC)z��.P�ka�(F�=����d��=�1�u��<���n����ިun{�uݧ=��`�Eq���'?e���v�y@�I�����\�h�_xݻ;�8�C�����N�\�r��[]��g�R*7�;F�5<>,\݀�w��2����}�)�PƳO�}ۚ�R�/ � ��:����
8Vo�[T��}!?^"_n�N��r௵2C9�˽�VL�8"���ǻ�}׷~��o��:=7ݒ%�}��c7jOG��1��t�	� �/��tpX�G�4ǽ���G�`c5�뫓n!��q������9hf:ڮJ��\s�T�<n�k�Џ�7={��0�{-���|Z[ؐ�f����"s��o"��kԞ�|=/pS�'������	5��"�i��x�=� �޹�0�"ٵ��zs�����ϳ��Kv/j~8 A�����<�a{K0,����i����{���؆��3�:#��Wm:g��܋���g{��yy���9�F+�����@kw���^��m	w�ڥ%�Nz�k�f,o<���>2��Ν�pΛ͹��p��|��~��	{ޛ�3��/p�^�{F�����U��s����JU�M�d��y�]��L����K��t��e���8>��W�Z���{E��䞐��F�/qS�x�Y9�]�=��\����u����=�6��:1���u�G������Ӹ�|�1az�+ʕۨI����Ǐ(!����5_�S��O����]æg��w�ޮE|�	^�ެ��{�efu�oN�]gð;�w����ĽFv�5�_l���Sk.{�^��wa�G��4ozL��Y�~!jȦ>����ťv��xe��4p�=��۲���.�#p;�������w���ǩt�����Y�"���l~8�g�Ҽ�Z��&zO�f�X���Jr��X���������=�=��{�@�׷������|����W�?s��38?X�������۷n��S����_-g���Z\̦�O��|���'��۵mk!��s�ɸ��h?u�����2J����X6���#�Z|㽊��\5ή���g��ua�QE�X�ͳ��D^�ۛu����u'����My5��^7d��v&q��qċN�L�����[vn�{����0
�f��u	�m�h}�Λ�l�/B�q��iۄs$Oc����XV�KJ�L����Iq4�%�lVbR�[��l�&V�`���O=�V��Բ@z<�q]�k�@���8�$��Lpo�n�=�Ԭ�[q����=����"�N�kEiK�ۮ�N�������\hܬr��� Q9�l$�4\%j](`��2��f[SV�.�*���cs�p��u���:���m,s�g�K:C�s^�5�j�ր�"�W�z�P��Zc�̀m��Q�le�	H��D����M��m R�ZD�5
-�Fl�[z�Q�1f,e։e�f,95%��!x@�3�A�X���(S�v�[�:�\N8�r�����<j�����Y�bls�\�����3��i�Sv�A���6�ڱ��0b�g�V���K��<���n����;��vU-��j�6��̜7>�N؂�SdK��y����c�Փ��E��ۧ��[]<�P��܀9��yN]s��`�+t���B��سXB��-������r�Vն�����n�K-��*��#���`�Ǌ�@�\���oB�V+��uO2�I���%�7A���ņ�)�;+�g��q���i�iv��X�+B��V�Vls61,h�M��:�S�.�ئ���l�J��hKq�Z�#u&6��	��ҙh�M�B[@Ҽoc�Wmwa�.2�[�բ���<c�����N5قm$gd�0.1T�,r�M^r�*�M�#�&��M��sx$�E��;�8�\�j��գ����P�|�ёJ[ngc8����=��e8顃(y�gp�2�t+�õ%uk���fP��7l��W�v̔b7n��f�����ݙS��GZ�����c���s��z�������
�4�	���/<�9x��fs���xN�-rⰻ]�'
��X��<M�i��v9ۡr�ϴ͕�єy"J����j1S��m[�v�V˞g�e���	[.��/ia��B[ ܷ'mza	���QR;�z��H�n�v�]�ѯVvx�=�V��Dq^R��W&u\k�[���=�R���q��ctW��1�pd�cd�����I2��Ogq��w3V�wr�m�8�F=���75����ǋu�h�i����-0BYtieu�v�g��Nlp�. bi�z�f	JfhgkNe���B`7���v�o)#�j���;]F��sƺ`�f���H���m��t��4t=:<P�Q�G�v�0�jIfy�ɐ�����e8f�ݥk��dx�y1���ōt�Y���K���H�an��u,��\D��:1�U��[��q��;[h�����z�w=�����yw%���Bh����p��c��Tח���ȝ[�
4h҄"��j�^��X�cp����³�u7'0l2�i,A�R�2��M�uuĝ]ٝ���c*Wo���(m�Y�� �Wi���0�[eg����v�S��r���TQ�k:��Ø�p���7]Gv�C���|�-�3,,	�o(�)1mᙻ8�����M��ݞbm�\D&f�g���ї�͡�K�4��V�!����[\L7��77l���s�yb�Qh6��<G:^K������ͻ�'I���ĨA�Ū�pc���9Hv;&Z�M��2�E�]u0�8�T	 ��n�S��ŷI6�!�g׬YyuwRa!�K-��8��c���@���V�%��Z�,��h��@yS.��#v��pś`�^K&�H̖kJ:cD��1�R����i��g�J�yK�y��a4	-��)h�E��Ɠq�;g��
۹e���u��ѕ�$ ��i��͈����b5��ɹ1\\�{��K��{-A�t���<��ss��ڍ!-6�f@�Z6SS�V�C�N�
�7m�n�ӝ�ۛ����n��C N��u��[&mH7���Wcd���(rθ<#'c�o�#���!������RH��y�Td�ٱ4��6nHe��&Y��'9�y1�H�.�Lj�&�W�ǥ�����áv;k�Մ��O�&�q�ʆ�CE0��4�2��Y��M6�R�m�4И��X�P�q���Mv�P�Yy��i�LL��cÂ`V�Byɡ�P�G5`��1�ͣ̚�l��1�mv5#t�8޳�rl[c<L��!7��b"�e�,Jl+�^4���0T��Z6�Y���8����B#��Z�ԛ`��i %[��i�,�� ���43��]��콮�\��,7A��	i�����N��fk��M�`�ivf8��[]ۦ�X���+�X��y��.�<������4Y�n5*b֌f.B͒ۆ/,Ť�b+4�,m����T��q:$��Y��ڒ�+��y�j������p����g���Xv��/@�YX���ۺ��)�"s�V�mH���u�Wq�YáI�����p�6oW:�A&*M5-Й@��N���������B�3��6	�;p;���]R��2����g��ʺ�Kwk�v�OY��Ev�gВͻi�i
k�q�c�����ֱ���\¼M6𕭼Jʎ���T�JA�d���nK�1�գ��j�{:�22]�͈r��ފ/
�f�Y�C�#� Iu��Tm�R�#fb�0̕hA%h��a�x���ە�q��l)x��pmqլ�����x�5���7Iv��g�e�|�v�e�ۅ:��m���;���c���<�[��l�n�.;q2�.��,v.�i�	��.*���q3�%��F˓���xN��\dHMp܇F�;\�[ͮ�X �=��8(ۚҏ<�n�[��u�s�Aϝe�=�,s��1�]�	�6np������^<����]�������1��w+VLg�s���u�ΰ�L��i�z�˝&���@��x�宨��c	7����[C�:�����굞m��bYr3YM��mDn��'��A�
�W�綂��6�p^y�e-jm�mkvD����������p���rA��99�P7%�K-qw+Bb�3ʆ[��,؈-�E[�`�t���s\Fخ�]���'��9��l�r8��N�����͐F沒� W��XW&�����,p�)��6�]i�u�cst:z˹��Jkc1�V�m���ݑפ�"l�+<s���	��`]�۩[���vȅm�,�ݛ�F�}����Y�uUqR���e��Q�	n���u��uk�C�ܪ�;ìڛh��'��۰��m��)�UbE��K�м��]�b���ѯJ [/9J��3⎙rʕ9�#�F�Ң��a6�v��
�bŤ�`A�r�c7և���rAsu�v�ۚ����isy���=X6ݶ�t\��mSu��35*�j9MgqO<k�&�s�+
�֌."Y�RVF�!nI�h�\S��kK.�Ú�O%t�u�M�x㇝�r���-�=�G��!v9e{6��
�Ϻ8�v��u�s�<:�kr��Vǁ�b��v�k5Tا`�9��R�]�7����{Rֻczl��t5��G���f�-�n;i��Wj0Y`ʤ����ˋn�#���żi팜Uw&.��X�4�66�ncW������=p�	�Eqj9�ݺ�n.�������Kf�#��f�[	����f:!],^�n؎�j��z�>J�aRh7Z�5����4XƳjF�e�`����e��ɍ}�������K-�Ǣ�)fn�k-̺�ţ�
"�i�xqV���\\�m�{��s���z��"��XͰk6*�0lI`4���l�!n�ZJ�u����a@�|n���٥=E�Z۱�Oc�1����c�ўne�NienN�Ɂ�i�\S����ܹ��5��rq�����/j.����H�Aɻqx�S�����|l1�gM�*�xm��pZ�(j��&Li�-he�KLl������=n�<�����%݈�r\ڽ�.ݢ΃"�]nRo6�H$F�f��R�e��E�e��'vް�<r��p�ڰs��훎T��Г	���r�%�n0��=�r=9m(\�9�|]r2u�=��r�t*��'�4v=e^���U9��1!Tύ�Sp'0ٹl�[w&O$f�r���@!͝n/<�l�%�ysc6�US+��R����va�r�\6�)�ˁ��d.Wr�:3U�����3�9�+��m�mZ�n�e�n��A�v���-��rQ�/a![g��֎����ݮ��[��x�k����ɓW�l���e�.rv::������MX�̥��P��fbԵ�jF��Q�bl��D�l�Cm+4fҳ�b�1n�f�����n+�y{h��R̹�X���󥕥+����y�E���,j�퓞��'8gs�L�QƐ�$w*�ئe�4�!�Z0=�Xpa7Z�8�X�ʻ��<N�}8�Y�� �:�݃�'R�N�s����]`��nx���	p�[I�.%���e4	㭺��j���O��-��qPX\u����Ûu:�	M\&nJ������Eٻ8�f��f���k���75�_Uc�K
&��^�ۺ�pq�a��"Ѷ��F8om�vΡ�{;#{8��PT)�l0�լ3���,yF��n�'4ږf�h�\沰���=q��O|��^��+��f��	��Gǳ�6�"�u�D��^84�ꎅ�t�z����8�l0����ӲYM������*b�v2�7[�nΚ���X�,��8�Лe`m]u�6oKe�΅�d�3�{��W�y�ڬ�5��&���֜V�-��&Շ#�dHU�^Y�ln[v=�׵VnVy�u啞Q�ս��m��tI�֝�z��Դ�6���k�{k�����/;��on�mf[ۻ;��gRjFw��m�����ZF&Fam�C��ڎ�;4sv��5�n�+��̛ZYm�դ��B.����H�6��T[["f�[��)%�7�!h�ax��!o'�ͱ�����;k��ټ�mZr2kfӲ;�#����^cI�%�9�\�ۋ%���YP�Y"���K[Z����X,a��g3e�VZ6��:��Y�;:�����Ή��G�u,�A#a/B�	o$:7��r�� ��e�kjmy[۰쵷dTsk����S94Q3�XN9�f(���o�{�aV��J�D��1�iHǘ�4a����z�ɧ��8�ħ�o��n�:h��P^�v���`{k�v3��tfsk-+�n��2��E!���Цb㙹띴�s=��w<a^�+���ظ�n���M���)�����+�%����E��=��1:�f)NN�R���C�X�!��������x�;4���x�`.�	n�������U��V�q�n��@�̈ghv��ܴ�ڝ�pz/j���G�8�5b]6��]-�(�n�I���ڕ,��U�,a[,uqlj�]��|�X��&����ʇjT�Pܠ�mm4�x-To�\��0D�.�J�-�,H�Ҥb�	�lܲ]7�e���c��,���΋��o-���O�:z.�]69��ϳ <�3��2èٍ�i;	�+itr���Fiaa�ٳ�����շiܩ�᥷]Cun� a��]���ms�<��u@QIj�3-�],c��
��q��1W�4�m�2|�����MkNt�:�`9�w�[AX�1l��jn\>m�И���N�>�#�m�c�;�fS;�n2�r3v�JF�B�6�!A��h����jf����j�0k.��+�B7!��Ŗ^`ML�h��1yݐpJ&^�ǚm\�G�^�:��p �`1t'79T㐎�!M�g���l����ɮygqr�v��i tl ���bۭ�Mr=(ռ��xa��6��d�	K��%�9�i<�.�d$�X�чkk�n���tdN7<ຳ:{8g���.㊻��y��Jv��p>v��nO[q��]+.�И3a5�CJ�e�������R<�;^�'�����8W��Ru��s���4�{b�-�5�%s���v�pm۠I�橱u���-�H����nr����[�ͮo���L�|n-qL���껦�iHF3ѱ��{]�3��m������j��׮ً4a,%,_zz�������{���{1 r�6Ǭ ��ab�R׬ᠲ�4�IR�T���JZZŠ��H#-��IQ(�ԥ��
�K����*���嶄�F65��@��9�RP�N�	Ia^1m���Q��m
�8�R6�J�BKV-k@��J�KF�6*^a,��"�#K
�[-+
��,l�ѵ	H��g�����l�/�w��eN<�2��A�y"F58pbk1h�ɋ[���c6�@�˘m��$V�+
;���]o�+F�uˏ�W�#7f �G�����ֳ"ٜO��TE[��e2�'A�t����E�L���Dm�]�m��w1 ���O��sOO������d��TV��F?���LXlk�A�/5z�b�38ex�h�����1)��<c="	#k%�yX��ֆ2�}�WA������ܸ4�*���/3$ �'.�\r�'P�m�7C3��C�l�U�.�$v��,Ͷ�l}��E�M���E��	�V���N���3�D�
�QX�`]���/7�/o��X>���;?���� �Ǐ>��}OB�E�d�݀9L|΃���;t^3���^���H7�t�����tR{�p�E���bͻ�S�ܚ�sDͫ��s�����,�n�'�S;�e��ǈ'v���l1F�7�Y}����Z�.�Ӡ��'��]l� d��?�=���
Hi�u��'���`C�/ۧ�K^82��̃��3���>ȝmvm�� '��ڡ �ܼ o���e�b�C$U�я=���-��gg	�	�P/SO>��Y��r
��;�?^�	��?��@;�1mlà�TE�ש�L��]�`ͭ�vҥD��p�6桥��؎솭�d����N�I71Y!L��X���M�� ����srb�>c�jn/-�� �Ή���_�Q��I B�C̽��?�&�RаUz.��O�7%�A��H����l�ogMB[L��v;9	�� ��<	 �\��O��z�������~�95�����1��'f��D���J��4�W�����ŷ����?N3e�v4ۇ����ݚᛎ{��s��~6~�$�l�N�L�ʴ�v哦b�v�Lm�d�!�+�|D���U�H$k�j��a���Ucf^�BS/[u�A��8�o �.�a�]�p��^`��;v�	$��Ǡ�;V�8�Τ�/��ߙ�|��9�
�n,�Y]^{��OF݂�[�j�T"���ղ�}��W��٦(''|M^z'Ē��A$��ժ嘊lƦ׼S���H7Y1Z�B8���X���bU�y�\�|M%��ۆ����}�� �v�B��9>�N4�'�~��0� �؂�����l?�af@b�(K�i�k,���^H����{V�'���������N�_s;kܛN�Ya9���t��A#]�ЀH9�������?��{}5޻_��*�R��t���g<��@Mh??���h��� �J��3Q����p˛D����k%��c+lh�U�"��m���wr��3i����S�A$m�V��r�-52 	�ȂN:�P	��ܼx�=�o�^�1>�� x��sHE�uhZB�b��SX`�,-��-��\:6mL�i�	J(������ː�ɀoDH4�n<�͹x0. k�7u6�����|O�;U���KP	a²߰~r�3i��ӷ۞}���j�`��E�V� ��ܸ��!屻�^_�*�R��?n��h�V?�g��x�D�Kǉ�%��]^Dn�$S�����t�Ui0e;���S��cv�m��O-.�d�����0�w%��ȝ�4�5��M��!�x��ʩ�8)�Θ���q�	;W1�7�"6��k6�*���e츂|wrb=��L�0V�K�0�K��k<��\$��V
Q�j7d�n����Aޝ���MEZ����g�/l7=����[h)����ވz�x����m��:���s�mn���s5f(��p�H�`�p"z��8h�p�7���������'�v�,��Ċ�[�ge&�4�V;��p�H�X���%���`�&�v�rm)�x�<K	��B4Q��seɒ=�ŔÈV�V9��ׂˀ�p]N��mu���;r g^N�=oZ�������k�N���Zރ��=��q�Yr��k��M�<�0��[v�lq�"v�h2Y�����Q����R�����Q�Q�J�F]4�@��ix$M{5LA��L����
vCf�	��x�[i*��\������\zZS:-��5٫$N��ǉ'�7& iZ�RN��V7�����	,԰�X���T� w& ����5���,�6H�ܗ�J>���	{PHGY�ӆ �Ŷ�.���u.,{��ٛ1��z}*��g�K"p���� ��HBI,X
�D���k��h��E5��b�ĝ۷��Aj�\A>ק�625��+.�#eI((�$�92���+�=�<�癠v�";{N.)ד�\Ifd���b��w�&!;�|�x$��sI������xx�4�w]�FfK�l�h�wt���.�&�:��� ݒ�w)�6K�y}kk�ƈ��qE�PYN�����;��w@�I��ï������UY�����p�vex�!�ĂIw1'Čz}1�Nl�Ko�{f�|����!�[� X��l`^�LCD����sO$�+r\AǦ���X:?bIb��7�F���W�{�+�.���� Hط����ޫ���F����u�/J	�3��/�Ė|l� 6�^/��d6�b<I#_�	;�/ ��:�[Z�5��緍���&qk�s�Q:�1��Cn؁qCЎ4���KC0pJ@�ni�Ļ��p]���ܸ�I���D�7n^�R-N�6cv<}��f<Hzc�Ń�gA�$���j�4i��{���2&`�5��>$ۗ�H5�x�Ym��cFe9O��gwL���f�THWO0������$}��֧݌мwz���zmZ{�Eof�Ѷ�����g+RD�Ѓ��K'/jRʸ���d�m��k;{�q影N�WW� �}|"}(�ח����^�\���r`4�zŻ2�s��^��7a��f�\A�+{��B���/����:?bIb� P�[�$�ݘ>�hOz1����7x�f�PO�5W/�wrcж�L��ߔe�͉����Q�Pv��d`�.ǮwE��01�&�"Pr�\�������\�z��>���������0 �?~�l~B��b�k�����+6^<HS������vN�C�U� ��O&[j��Ŭ�|I ��|_�x�|Z)� g{V�DkR�^X�3"�3�d��<y�"<�;wq� �i�Q�L��F���J�A3�/I�ڏA�6P6��p���F�Ys�Ө�6ϕ珣^<A'ٗq�2�����b��fvyM/xlt7��o����ʁΌ�~�v�k�h\��{x�&x���{�i��Y�\w��`�y�^�y�u�=�%/��sk�%g�(}��e�<ހ�2��
f�5�b�L"���������f�/�����`�S��=���j�5M�Wk2�,���i��j;Vwz�"�f,E&��b��|�V}n�;R@�19o�n��H1��G��K,�4�6ٯ�nm��	7[Q�%�A!fZ�w�<	��r_�!7�Vb��}>��Z �}w�9Z�N[.���x�H0Ғ]��:I�����pW��K2X���sZ"��٠��� �r�b�5j�^��fE8d�'`�<u�������`W�A;-��Iv�楯"��ftA{��2�@��p��� �*�����e�Nϔ��>Dn5z͹x>���@���#WS��jx�u��»�{�������Wyw9J9�??B6x��{u��oz�m:}OM^^��]����]��v�t<�ZVn��U(�UVAka6tb
cm`�m3Z9)ogM
��8-�hnA�"�vB���]�pm�� ه�v��.��ձ\ڍ�8���\�R1�"[.礘,�Z٣Fݽi3�����J�S&�����ٰ��Ǩ:��t�N<�ݵ�rh�౮�b�
Vtr�f��2��m���<�rGE6�m��J1=w\�N��{��^.�v�
U��W+O[<����Èڳ�]���GM�E�qp6�l)3�-���85�������&d3�'u���N���dY��׏��|�����u�A8�/�O$�{���\�*��	 s�x���ߺ��,�~����w�Ԡ���;;3x� �-�c��H�����ҫpi�U�$el�-�� [�`Dj!L]���3�G��!���	 �\�x�F^��FCV0�'�K�d��Ι2v"���x��wL��7s-mhv�-@$����I �~�?r�ӯ-'A���� 5U���$VR�jGA�Q&�]nƭ���J6�{�z��S�Y�3r�5h�UG��EVˈ$���������Y�o�Y�&�ܼx�f6�_�C�8� �`1y��1���E�+��a�����ޛ�5G%�����=�<���pN���pe�3��=@ՄE[ouQ�F(�N�-grZf[4"I&�%�oj��y�3�ɗ�@�w���BKBD��@���	߫c �&�˘%�/2w�Y�I ���6�c�-H@Dk3��d���m�5_m�2I<m�$M�Ǳ��^g�v�/Nq7S�a�-�@-ҀO�W|3���:�*6|�2�O�A��q ��O�6���xn��bz_����u�턃�ض�YK�N�l֒��m�.�r���o߷�ա���gA���x�$_�8�1 ��O�f��C�l{mX�Kӂ�m�	�Ɂ�A+b�33�I�@ܖ��|���^F�A'�/�m�bb�Le��Rշ:��#r^I��m�,Pp䡮�B&���������q����__W��|�_\�uq_s)@�K�7���K���;|=�/�B��ɨ�d����d�hlyg.�=���{{�-����:�bp��Wn]=6�ku��g�c�=���9�,��:�f�:�E����������}�����t�f�Y^_�����(x=:��&�N��.�^L�@���Ń6{1���j�~�]��ok0��^����5U�6 L��e�����3J�@z����S��P-���kg@���\�͙ý���ms�Z��^�z���2 =�N���e�ۻ�6븵�.��ksv`�c���qwI�a�y��|}ݡ���9�k�g	�ّ����y}�*�S��/�Β��dg&����Z�uW� �y�t/nwq�k�:�V��\�9�9�������0����	"{o�l��L��>SW,Y�v��\�Re��u"����P���;��o9�T�^��Rxl֮��� �� :����I(vM��U2���fwl�Ǵ��w��ti��⎧�2�yU�@�c/��ob@8�/j�MX�y�cw.���.��|����K��C���o��Ww���ޝ�1�_����=��7G����_h�5��QI���D�q����C"�{4d����:�2E}�3�頍�����_��x? ��}�1�iK}tםT���� ��^���1�9�C����Y�S�68sVr졾�DL�ݱ&�a7�~f�ނBy�}�������H���黎b
�M"�U���vK�g�nxm��MRq�7Rc��b|6�k�֓�ӛ�9�L�a�� x������d�����V[ۻҼ���y�G��Ji���t���m����dv����Q�\�F�@����㈭����Y��M���[��g�W�m��o����ua��K��],D��i:������hk6������{z_n�9�-Ա����L)`^�	�a���XZ�qH<:�n:��ͲP�u�1Ω�/�R(��w�+�l�{B�b#ݬQ�6:�Kkk�-���Hd��x71��Ic\v<���Ɍ�!V-�-�65�dsg�^��/_{��C쵨���R��X�v+�]��zc.5��B�m�x��X	cI�!1r�[%��X	z��+2�V'K{�|.{��s|�:7�'^۽g��6�{u��],����r�Z,r�Fm�1�$�U�N�:��l���'XE�3y�|�<�nu�f��nD�xr�sfv�Y�o-"}���vf۫*-�bw�M��f���털�w�Ol���Lþ�۩%)J�Sq�<�� �^���ͥ�;��(��!x"�@�� �
͞|��T�`O��mζ�9��2\�rL�>�H�>�'���|�����v������rR��2:�;{/1�&y��ّ��gU%7���ޞ<���Or���	�k:��<��a�%�dZ@�E	�����C�Jy 2N��x��$���=}Q���?Fʹ�t��ʻ׾s4n;R2�غZh��E�bٚ��wZ�c�+4�@Q�ԝ�ܷϯ���p������h}$��y�r�̹JRk�o�3��!������BrY u�\m�Cw:��>�$L�8�+����P Utd"$ �^�r�$�t�ȟH ��} ���#�=�ص��9\q����	�aI����91�;C��	kz�y`�L��ͻ��g�����mD�S�4$x-|��1NŜ ��Vt�)z}��{��̕���@��* ��<�� �PB�׍!o�x&�������u�5��ːd�	k�z���:�mYǛņ��oAď1��!����N���[Ϣ!��O��.d����p�;JR	u߽q�'%��Y)��~���p�����l��̙�����9��'Ss"��!Dk
�N(S=	�;-#Z&�=Ƴ%��̻�F�ҝ߷a^��]�2?XW(�^-��4�4��x�XME@�"AȄ#���,�Θ����C�Oy߭��� 2R�;���Iy�Fu����}{�W<Z��Rv�S��R��:��8 b�����7[�:��y��C`�&w!2pĹ���i[6��������O> :p�箘�~�>�}�>;lm�o�	�d�s����Ja��	�z�~.HL���������9 �${t��ʉ� 9�"gb�y$�Ȁ�}�@@�]�<�	#Ȁ?)�;3�6�޷�z��L�;�o`哙p ���c��ٟ�g�t�@�>A�FBc�z�a9�R��ÿ{��%+�<�y�7�c#�	�ہ�E� �@F��b�v!:t�O��$�5�^O���N@d.G�����y�%�0�$۞�%L���^#�G�}��:��J�rC2;�w�/,s	�|k��1Nřّd�DxP(�v��x)�[=���s��9�n��m߽�ĥrBd`Hdc�mޱc���������s�Ta�C sv��y�}�G�V����>Mee�y8vH8��>@>�峁̜ˁBd']y��<������/n+&Wv�>�$xNF<�|@�%0�5���C�qJ�L��]wǼD� ���N6�������bJ�;�ä��i>aԯ�����Z1�z��"٥Q�_��Բ�.�{=�u0�ޖ�6l> ������/�1��4J�rں���,���rv�xm�����x�햭�O^���Yz�\[�դ�m:)���;�f��[1�&)��f`�(˨�n�K��+�uy�i1Ӫ�&G���h��nmd%�+\�:���^4��]�/��z��A�Z�z�Y�/X��㨯GS.,
�I��g������p/4:�	���IGS^6�)�"�	y�:�۳�{]���G�f�T��[�1T�)���Y�I���q>V�ڴ��oI�Ηs�O�N�u�w���K�d9����9)C����9u΍w�x�B]�ָ�^B������o���Y�΀�'���s���ͳ��_�~��}�){�ߪj3�A��`�iJ=�͸��9���S':n:�|}�@G�DZ��c�Uf��Ș��Dy��l`Yك����!����~����ԻA�������Ǥ9��#�G�s�{���)��G^s߼JP��)Iֻ�q9y�)J�M�@�"|�D "�\�I;!ܹ� � ��|os&/�TXO��z\�}���e����R�g]y�<�C �"<�|���>�sD>>�\j�o�JC���kp9#�L���3<���r���Vt�)z}��{��̕���D���ʈ>�&�f��l-���>�(��k��9I�`2N���p9-�">�#���D��U����wW�>����J��WR�+u�m��޸���� ��,6�`��2�Q�������p��i�;JQ�q�zI̸d�'\���y�>�'�"+ީ�<$�<5e�s��m��㾥<s7���9�+L��ɸ�DIȄ��s3.�)��tϽw��@d�,κ���^��.�wgxK�ȺpD<A&���i��{v��ȍ�-���Uʴ��ƈVn��8B�]�h6�[I0-�K�p�g�r�_��)I����x��2R�'/� ��@D ���|4�㩷�pY�N �$���t����)�R#�D'={��Nm�0s�0K���.XL��$26���6��3�=���C' 2r=�\y��)A�C���\q$��|)�Z�N��;�E�zH��������� ��}�O�cvG�I^�C�2C#!36�]��'-��Y(�C��ǅ�b��}::��E����#� \=�1|!z8lYb���;��|#��}k�'����J=�{j9g�@���|ȄF�V��|G�E��1$�2d�Ny��y�jOr��#���@�"<@
�fsy�V�1�f]���>8tؙ��l���8�� �mN5�1�mv��GR{����,��gO�I=�n��9�����C!-k]�]0�bBda!��^m׸�1�!�{���S����\����<=�1O���Ȁ����>�>��ko��3��8����2=�=��^`�sF�w��{��6���D�!�������BrY	�ö)�a�Ǹ���&T�1����t�P��}�H�+"t2���(��!x"�u�DH |���:��IrLa�	�m�{�)��uB1 ֥|-[מ�r�1���}X����Y��H~s
˾���/��ܝ||��8�R�G�o�pa�P�ꕈҝ�oh���w���#�P�2\��Z�%(I����3����Y�΄����$��l�旤)Ώ��U��^�$x���d���!����׸�1�!����7�<�]�'6*j�y�����k��=<���w����33vԯ�ެ�R�)ֳ�`s'2�K�'�Ϟp�O�饍��vӋ
��I�Dx��'!d&6Jfa�z��%+���  kM�9| �(�J�Lz��G6���sm�^4��n4�7e���;Uˈ9��3�Jf��/51I�]�s|������x�y`2p��2\�u�ڎIy�rR�[s߼���&C���y���糆�|(�[q�"QI#�O�D����Ej)ػ� �Zݮ=�.e��+�3��5C?Q�<�O�RI �ۭ�2�Ir��rd$�D���2Y���N[����\V�x��܄�Ĺ����eٙ%Fs�a If����n�}Б'r�!-3}1�f��Xjg;(��n�uU���爈��e�%�u	��������	 ��SǏ���<Ôl��\=�JL��B1V�Y�Ly�d	�r��q���t�n�寮�|�z��-x�ӻ��^�8W���e�Xjșטq��B�86�F�|<��{�	'c6	Hw��́d��ȧAD��e�$�7�O2�y�Y�c�2��[���H��ݒґ).Χ�LF�
�k>����5�" �]t��jkn�0�a��0gl�9��������*ff�?~�m�I�� ���bI3����)��ViX�)wnH�E��k�i	 "�m�):,C����I}}|��N.Ӯ.Z�v�G��I9*�R$���J(�"���!�w���f���'q��b��C1hg�]ƺI$�d�̢Io�{���$*�:գ($�]-�-!%��	nO<�@b��7�9LK�];0�hcu�O;YtIc���@��.�א)"R����x�q\�b���(�ꖐ�>�c����E<�5亮�e/$��ΉZP3�z�6Y0kM�O�I �\�̢Hg:�^ �[3i����`꺦C%*_%�y�d��+o� ��r{7K��]�H�~e'כ��N��t�8α�edd@j�2�lʸ�,%([�)�,�_���O��Zh1Y�f3m�_[��nRw!�6�5uO{;utc��k���cx����]e3l��@��&o
ޗ!v�F�8��s���l8��!+�����,���;��ق3�Vn5��/Y�z���&�Dm-��܆�nưS�� ���r��l���z�T�	.��g�n��vu��`�S�7��z<]�z��xv�.{)�uqmZ����+k�%���m+�l�`3]I�:mn(���(`���~�pw!�w�t]��xSQ~��%�<�̢RK��D�Y=���GlR{�'��sGN�@��Ɂ����n�ҷ����@���
RQvT�eͪ�5�R��t�@$�Fc�2�]�� �q�n-،�W&�.��mJ,.�'%�p�<��})����R�I)��gfw
�t�>��K�њ��[�̒혓2�F�8�'gL����v�\����ۧ�R�>	$�]�L�%
�3!"vq������Lk���i�DZ9�o8b�8>���ͽ�����+�n�>c�o�ۺ̆��ԗ���@I���>�W�]8�*@K߽�y�~?��Zy��Dٔv�J�4f�!5[��م�1V�M5�`�#W����~gnŚ$�Nw�5�4Iy*�}�+�"����R��7��-���;�}(��\F�����3�X�d'��I����8����*ST�p�SR�!;Vg��5�m���*�ݘ:G�j��M��4>�lc��^��i��T�!���b���J ��]�F��y��[�HRIP�fGw=ڍ���ML'`�;:!�����
W�A.�ǉI�S���=�"$���o�A%�W�e]7�$�A��d]!���%;vkJ��-Q�e�D��̀� ��̐�މ2��H���ܒ�1��x$�<ř���:�'gL����/um�JI$\���P��:�r"���+���^���2I/gVĒd$�7V��o+z��	�D,š�1�%�Gn�l�;s�,(ؔq�;g�����A�;snŃ3��"dR7�o8b�8��c7W=R� �׉I.�f(.zי	4eQj� �j�L�l�1�	���	3�������p��5A.���H%�ܷ,�M��^4�R��25���	$���	���p�&�RUGe,����2�&rK�$�f6��%$ήy�J	�Ș�m�xc��r>oO����wGv�w��r����@�}�Z�wz��{�[s�h�:l��c�w~�7�_����o�l���𽯢L�$�I}�kϥ!@GSS��'�j�J����O{]6��J'y�R^I�Al�<�I$���&ý�!ࢲ��w�d��k6Y:I�p�<Ą��^D�A.֍��O�Q9��Y����HV�D�d$�K�d�<�Q^H�4r�+S\#v���C�P�����@���7O].��rtX�Y��U�Q�#Rn����m3��#��t��4�v�� ��F���J@�����AOS"'j�D���މ_����9]/>��!��Y��`�X����P	M)�\�-����	$��\�̮�0e�O�k̩�RLs:rgW4��~�}TX�%2���$$�W��y�	X���J	!\$��d���t$�]���QI �9A�&8$s/2`��e<��l)��30��A#���:<����1A$�+�b<UT�۹Ǜ&��Q��N�sp]�,�c"Xn��^�K���\2�k��}��e���Ӊ�:�u��,��������O��9�N[���m`�߽�x|ג^J&m�ϲ2�����;�A��%\���Iy/��C�q�X��y=V��I$�qL��K��H>I��u�;k6CR�I��t��&��eŃB�1����fS����Ė1�Y�]�q�I�&.Hr�:{�(��L����ҒA%�o��'히�5�r�7S]ғ]s̠
E����8N��	�L�9U�����w�n-/}oBR	�[�)��Ij���B4�����QB�nq��OuF�����җSd�J	Fs��� 	r؋��5����f	 �^�H�$)�����>!��1	8�D�E;.k�fx���$��l�iI �KT�K�I%���c&�:ɐ�	w=J�)';$�b0p�c%�gE��H$o:�}*��*#�A%�~�@$ϱNt�����3]����p:q��q��|}{����=�@�l�܂P�4<��Rd�{�
_v��Lyf�P�Q�'��������D-����s0M��{ݦ�}�+�gE;��W���دBZ���vYM�X�=�ZTo�#�{�]�F{#�%��_�UMɦ����oB!��[�=ZZ���U�U���p�O��,^=�$޴���!�>jR���R ��w�3��]ق&\�K.-�n�&+�Ͻ�{�|�E4�u��1`Tn�{���>^��d�<>����ōl���^����um�۽K׷�}�V�|s�������ik$�����O�w��|R�2�}�; ^y����$���=������}�d�2�3�ل+�m�1�o�/��=j�]��r��W���O)ǵ��q�����/<�"z_X6p|��=�9��ռ�t=�=��k�zw�o�o�q/f�7Wo�Â&>d�s��,�Ҷ�T.���{T�wcp���t���V����>��-���[�>^Y������pO�8�)es��z�u�9c�>
��0���RP�XL�B&�C��U��e�1M�ל�gw }� �z1��%r�{��`�v�Y�ϝ޷y۫�U�q[�g���G.�^=�S�A�seg�sK����xɸ&ٰ��Wg��=l�.����dׇM��<&?M��{������-���.���D1/ Zc�y�{.N��,�*���2��n�y=������f�$�e��;�'����H\cg<>���߆��6��z�x坥���4�fکJ���g`m�R+ȸH"0=�ĩy0j���u?�����Ȉ��,�|ڌذ<�#Cf�G�k�}��o�Tl�V���m�[�"������޾�ͣ�wa�l;��1e;�c����� �"(���a,JY
A�{��כ�ϝ�{nma3I��e%��c$�l�g\��G;��ݞw�Ohӷ(��ƙ^w�{�[v,�x�{^�����n&�Yͬ��Ҷ����[MU�����:Ȭ����s2�-�1��<�^��l���N������3v͏�{Z�4'}����<���dt�e�y�Q���s[��,�y��K��7��K�e����������^�R�j����k;5+jɵ�]��T�6[vظ�,8�k�L��qIkb
;[�]�����Jy�1���/{�6�����k{�=;V�$�[�y}}���AĶ�[m.۶���KW'����-�Ds�(Ue��t10Wri��jݣ���YRX�6���Y�k�恈�U�ĴIeƲ��lq���(cK�23GY�8�M�8�U�Ȧ����w�(j�X`����Z�/G\:[��1�q��Bg��GgF���ƃ��
>��fG�c�2�Z�Z92���DN-�m�%�4��w+ �NG���s��m�1�[6�5f,%�ɷ,�,��Ԥ)-T�#�s)t!r�꘠Kg9�撦R���&�WYEhu̳!wGO6\���--ƞ���5=]��n�=9��(�v��%n��k�3B\����Gj�Rk�n9�2D	HE/.,���Ն�&����]7P�M#�'k�Q5�D�Z";QWn�p�6�.�T����щGU��[E�f���퍜�̮!;z*�מq-��1wb�jnM���R!�l������6�lq��pU֣/=2��`$�c�l�֠&��k��C\�ѽs��^F� �R�K�� H!ڲ˖�[)vۊ��u�D�Ǝ�
=j�1Ov�u�$Ŷv�N:��΍z̐�hh��0z_7Ph��u�v����n��Ƶ֍a�qd�0����u��E�I��=1uUn�뎞s�$sn�p���^n�X�p:g+���v�#�BU��e�M�s�� VJ��hHnҥ\�%#&)�V<�J®ݥ��Ȩ��Є�����ً���'�cg3'g��v��Yg��c
�P0Tlv�\m:��M�m\v-Ϯ|���3G�Бۡ��Y�RZu�t#�*�K؍Զȶ�vM�XR�\B��(�1�汆֖�fx���玺8�^v���uZ8��L<����4!��5�۰N��t�{��Ȗ��,&36.�	�z�)XX��* '���{lٱ!�ġ{Me���u��4��]t�2V
��]I�\�㞎;=�%��$��ڝ6Y����Ou���,�b`�&)��m/N��:g��{p�ʉ\�c������	چ�qc��΢�۱��Y�5�Iٮ��MՒ\���{�M����ո��B��6�\��C���C�<��M�8:Ύ��2ZK��M��<x��%*��j$%n�/cb��	�sc��r`U�n�ĨNu�ƥ��ttZ$�&z;��z��tf�,�fML�V6��W7T�ˤeI�]4��<Y�:�	D�mpn�1�F�f����Mbe�6��(#���V�Q�����?���mR>'����.'�RD�r�Ș(��H.���z,��X���T�r�N���ə!��e�$.K*�vf`�.�bBO��>��{Y�[�}�����A$>\��/!"R]}O�H�u�9���;��|�p�Ι�	�URӗs0��I�ǐ%��	'|-���n���	/$�(͗��+�s�<�K�oHI�r\�q,O4�F�����u-;�	$�G����I��>�/�f7�DϹnT���E�!�;"
.qB�ש{��RA*혐e�D��#�\��A�\��D����&R^]Ѳ �V]7[=f�]0�v	��&p��t�[\���ծ��y�r����
;�4�u��'|���_�5������L�X�IƎy�JI��!(g���Oo��ʢe�$J	vƼ�^��j`K;1p�K��%][ I�#�}�h
2&"[���Tܶ�w	n�PZ%��żnf֩q	�H:���[��9f����MFX1�츺�Wd�7g2�,;���4�ނ\����<>�3�E�D�$�d|�L�_}"e䵢�N����%rP¬'ff�I�%'�יH$�]��> J	 �K���������I/%}�(���l�����X�gL_ɃUP�U�K�I�}�_r�2&-��JA$[��&RA ��d=fc�:��x�HV�Jc%�JT��\�L|�f%�y-{��e%�Vc��&����,]�9f��}��)���dL������|���wPƐ�Ě0�b<Ν:w`�E��\"��<�F�l����/2�!��,�V��~}�/�ϙ,�p���	l]<�) �	WF��A$K��K�w{/|2��S�(�'�3u�ȟJJ1B<C`�İf3 '3�.g�ep�wݖ�Ǳ(��tl��H%��a��æ���8x:����JU=Mw Kt,����7���	$��s�N$M �nوx4[�a�%(ʹa�z��m��]��^r�����rR�,�2��y�V4�ɳ]I�����V��	?�xfNS�^I${#`L��Gܟ퇔���a�XN���I�%'�ז��rE=},�J�*$�$�����I%��� ��l:N ,�,C�\DLʪ��1E���d�&�a%f�Ŵz�N��L�vվ�/���! �V�6^BK����tW��4yiHwwY�����.8:-�]�8���)�����L���O���H�y��@�&��pI%e��$�K˟��B@nX��Z8��n���y="e��r^BK�����\$�PJ�i��IT-ohH�\���Q>2�H$�'�K�7v<�E%��[�;NN�]Tg�v�R �gE�f���ݙ��7�/�� J$�	MEi�yqH�����i$��'퇔�I7v<�Ww�n�:N��:!@����<�e-��؉*�R@%F+"}	��+ɺ��|�I�����)Xfm�,�Թ�S��%]�O�k"��{�Q���c$�T��̜U��ٹ��?/����{�Q�-����)y�ǵ0�"�E|�������E�B�K�]%��]����"R��y��D���*a���֘���f��R�	/%Oz�(�����Q۽�*���}��v��tK7a�a��4����u5�q)�.Fi��B:�`���_>،�e�1�_pZ^�f($z�})y$Cz#L�<������ej>J�����x)gw)�ќG~�F����Y~�������Ą�o۷1L���� ���y��	 �F��J���M_qx	g}|	!���l.�AE�N(Uy.����*�}���[Q	���,q����w�>I �	_F<�)$��4̠Q���gpɘ�b�	�����`Ku���f��=�O���%gDi��H$�s.�s�y�=o�@���~y�s	ޟ�^�nJ+t�X���*�~�)%���H���7�g�� ���H+��R%Kڟ�\�<����`� kwkD(*�[�)[�T�=[�u޵ܚs��]y7�J^�� ,H����VA�c�y2=�1O�ؽY�;`��<<>>��< ��CJwrQk�������s��{l�m+Y� ͭ��x�0��\��k�Q�b.��Xl�� �õ�@����6gGL�M.ڗ�-����U��Y2l�xے#�k���^y2d���N�8n�Y��4���iL�cyãx�F�B�h���Vd�C=`�<�O5�&٬b��0K��,՛��X�2�]fV�j�tCh`,ȍ�b��e�R��&u�&�+�q1�/\ms��ۛ�L�0��tr����3?�/q��~�x2�	n�l���'K�C�N����C�OR9��O<�QI%Z��e+��!����`���E��I��`b0�FMD>gי�B���I$�ne�.L���o�&�e���O��WbKp�� �L@���C^KJ	/f;"a$���h�Z�̙ޥ� Tż�{Z%O�\��^RS�`�m)����\�ߒ��{މ,*8߳4�3F�ʉG���{��K�H$�Mݯ�"�#X�Cv�Y wy�2�R��y�݋2%��c�pBD����*�u�ǲ4ᔫ�iA �HR��yE7�0I�����ɀ�G;h�����B���yM;����)��q�f���(�e@�YD
���vvD��wr���}�*����(�KL^C�>E$�wc�/�4�絳{c/�*w�R%��v^BH
����2g�� ����%	�e�Ow%�C�a}��wf��~����jgd�youk�G��ئ�n�gN��S�2�8�řy!�<��;�OZ�ɛ"���� |�c_��a$�e��(y&��y�6�'�1��P�T� ȫ��!�����.�1˹�I$<�n�y��I(����%��%Vy$��'����	/$�|��C5%�QE�&!�.v��Z�{[x�Y2ӛ�>���A m�y&BK�y�Tk\/��^���^RGc��S�%'8��=�m$�U�;!�9z���Y�$�eT��J�Mw��H.�R%lUG#c��&;R�_<����m�l-^f0f�)�'dw0tqL8^q��nc@+�"�Ry����m���o�8'3[2!�-y� JH����uL��m�#��������D�n�y�o�V��#�$
%�0�����Ga���5sE��c|�Ȕ�ceg���%��\����9���dNwk�IBZ�rgN�3�	yy�J���J%�e�T�I��+َ��7P��wT��1j�����s��Ȃ3��ޏ(���ׄȶ�3J��5�/M��=�vB�}p�Yo�[y�x�3<=�U�Ah���/��b ��(����Ȕ����3����$Z�������h鈉�v�D����% �@%�1�d$J�n�m�uo?VrM#\��Q��>���K}i&)��\K�K_�JI �T�'Β��Ƈ8H�)��^Y��3�B>H���D������3�{j5���hU�vh�GcQZc;������i9ީ�v��ѷ�5�2b�DML��f)'�p� �������
W�A%���ғ̷LU�TO-w+̧�e ��"R
-@\���1%�̀�WtˤdϾ��"�_gd=�OH$��F !�H��։&"��N`�U:�)Utӳ�gpΘ;9UT����<���@$�K{��n3��R���H�dF�W�Z��
R^��[��.����QI\ƺ|۪֭�Q�3p�$�z׳�	/S���3/�I���ze�E���f.$�K+{��ܑ[�r{���a𨫹DLs��t^���ۋ�;g
�v��+���7Uf��L�4�>����(Ī� "R�V����8̥5��&r];:b�@���q�s��I"�l����#�ۺ�埅DRk'^O�d�y�� ��$��^e��_,������}��b?tZl��mc*b� ��3����6�(^i`��m@ɹ��Z�O����ҴѪq��.�{��,�3#�y�dI%���BL�жYioC怟f(�"QA$>�Ʉ�?dѣ�����՗-���910��i	�U3��R�A �>?J�C3��}�x$�ڻT��-wp�9HX���1%����D�$$Z�e �JC��zM�z���<���e&��H	z����ػ�郳�UIT���'ajbt%Y�) I��Iy$�;g�#3G3�Cm�	!yd$��*�7'.0g�/�Q��y���).�ؐf��n�dK�vK��ؒ} �H$�z�(���� J��e]�oJ5��)��
Won!����r��)���ndե��uf��4��M���^>��݇��C�Bm#���ν������W��f����*�]'I;����m�%~L�yvn-�a��)�3A:;B�&l۴�.���6X@��Bnr�j�n�V�3H�:�/q��i���b8�ۇ:��o<ձ��[k�k��G؄�Ӥ�C��۴ڷY�g�YV%�S�Q��[��������1�㫠�A-�,���N�iz$�&��qj�����e
��
��n��i�kv�s�1l��ǘɂ㛋s&���)vͱӈ�i�g�vZ^��%4�њ����Ͽ����"�e�t��T�) �%�1��I$��l�'n����_1z7f$ςH�k�x4s�[�h�N�2q`�ȸ����!mY�;e�⼒	$�VcĄ�I-��*`Y�#�F=�Y]�$�,K)�1I9,�P�J�m�Q$�Nă($��Ӝ�Z1,Qxl$|�@ u�̢�;Ӱ$J@(���˱bK1�	��tf,C,��1�	g�^e H�+$L�����tIx)�^6zE�c�-����v��8�%�N&�U�a�	�y�BJ\���n��U�2Jr%�d*�0L����e#�}�n��.`�,�h����[1�"�`�lZ,v"wE�uրC��*�7Bv�a,�<����h�qw��-�Ǒ(���>�R�I%��d%���"�hܜKz���QA$�"4̥��A��1t�C��TD��2��j�5n�n{+��8G,
%VI�g��:}ߗg�����p\^�q�x��|�{٪D�֟g�_����پ��X����ow���"{�� 	J ���[����33��\q�səKݿLI��K9J��]4TYۼ|��z�$�R.�$�^B\��*PI$}[�!$�	^�r�d7q�ť�=�up�Io���$��<Iz�p[Spb�1t��.¶��%�_�Y]J90H���Q���Cs&$ςI#{<�!GF ���p��萇��G"�Hht8W��R�&f��#lQw�W� �{��2%{��$�>E�-�i�ye�3�9���ퟻ}�ޘ�2��7P�If����Q��j�ֳmJV&m�z�l������u�6���	U��^H�ْ�!$�!%ݍ �I{�.��$��Z�Q%{w�$ϐ	{=�.rr��p��{�D���6���+X�[5���RI+�f$ϒ�31���2�$��x�͕5�W�vR���Aٝ1)�`�.�tּ�b�	J흸�3+�8>;�����������ϧ���d�1�b5�
5��9�ݘ�ɣ�7m���}s��G>ٌ �a�wL,�c��LLe-�v��������>����������������^o���-]����^�'.�Fd�z0a�h����w���C��7��vo�ξCs�7�кռ�k{�v/Y}Ńy����>��}�^��'����������ط�W��| �����_
G��,�T�����<����yh[�j�KNi�x�J��,�mM�e�D�o���p�s�ų���-F���xzc��wP����ޙپ��v
��w��䦃䯔�;x]����mW�6�g��߼6M6�_���]۔����p��-�͓{ ����Z��^����C]Qjѷb���nM�C�Ѵ����(w�Y2�}�3�����6;������+�v;�9N�n��`���W�G���㼼L��ퟀ�����q�����l�xt	�}� t�o`��v�b�Uo�˪g�v�ҝΚ�a{&v>�%;�/&�ѽ��9�{w�#ǃ\1VO���(N���?[�T��r�p�k!Sۃ�O����4��wP�}����{��z9��2�&HJ�e�l�ۗBD���������߿��<��t���ܧo��S�|�鷰����Z[����|���"��.�������)ޚ�e�'�K�t�>KN9ޯ�����#N �n$w�a��sϸxg�>�7����c�#�_���7��|�~Wp���b.{~���(�K�NQ	�3 sZ쏤��������y���??o2�Zݍ彬�L�!�,�(����3��I;��|�m�1SkKm!�۷8���C��k��,GgVd�wgm�
K��2�6[nm�Z-�͊tW����Y��]�l��y�v�j��K�,[d���-���Vw�{g�){df��.�D˲�����N:����6�^�zy��4ۻ)������i^��pqOi�f]����kDq��Ֆڜ�I ���ض�Y�e��vk/2:"2�:�0�H����^jw�'�Yf���;��o4�̭n���9���g^d��A�&`�����5�TᶈI�J�[y�/n�yz��,�J8;̯i���`���&�`�66ˁ��r�J�5���ffaߞ��7&e`(���R7LU��'�N�]��f�n[��s��$�tED�$��cީ$��#c�D���w��I1�e%76-����Y&.�\��Wϖ�RI%}��<_j���ג^짩D�d��1�e$�F��Ղ�tN���A&q�{Gy��tt�T�x�:btPmv�-����;E��&���;8gt�,� ��sN�d�$A(Y��%@+�#ʯ5�f�C�7�eJI#�Z�B�r�9v�;����O>ς�����n�S\"N$��q�BI$����Q�ֹ��Cr���%��jr�ؗs���涜֐% �!.}|�)$���<k��N����-���E��>������"��vUK�q�#���MZK�_6ʙD���?F ��zbI��i�DD�u;h���pEA}�&t�%�v�F�N���3.�/	��ݹ�Vᓆ�A|��rZ^�.��WsY6�q��  |}� 	@�
� 4|<��I���"Vf��l�&�N TR]��*PI$}w��JV�a[��)1l��d�:$̤J\�dJ$�7:bL�:G�pu�.�f"s��.Ν�$���$f�>(��ʞ&크M��f�)/[�Y�ߩ���زA���<]ř�����W�b|�(
Θ�>K#��Y� �x0I���>쉔��d�!6���P%��P�o$�ӫ4胗1Yѻ��vRI%Oy	�$�v�I���(Q�JJ�r�%�Ȕ�aO:O�v�;��&c�OU���$�2�οN95\U���$m��H�ICs�&B!*L��rȿ����(��4x;�<y�C�D�����$�!{�e$���U
6�W��$���D5���dS:��)�UlQ$�I��ϼ���>���7'S$��dL��	/u�D�I��g)��=ٻݍ2��4T5k���;�������x�+�/�+�9�{��0o��iNNǛ���TW�4禔��j[����Z/��wI����@O����*t����o�ձ��4��(���F8l&-��ۉ�;m�����q���@���qњ� 4�I5�%�Kt��8���ⵣ<h;=p�.�ɥ,%kA�X�l�����7iڷ���{�7��B�Zb]�6ְ3�T��1ڹ�&�3s��4ܬ4��E�͊D,.5�v�*p�Qv�ݻ�uW��sUC���k<c��z-�7���Z�����́�"�@���.%�l�e,�ٰH�jH�e4	Z�2������ �&Ц�N�j�#�)"kg�	$�m|�2Kzm�gW�
��%��x3��mmv,��d�;�b�U�Z�K�NL��ᯜ9NmŃ+� R̞�2�	$���e7�y���\/��]�A+��Qkp\2�W��]6�3�K� lm�>��H$⃙�bۜ��wѤ�(��|�>^H�n|�2�T�c�����N���T��h���f�R[y�A,�k�d�I/6�b�d$u����hꈾW<����D���˻$�O-!T�j�!�	s�쀧�o&ő<�'!�K'�HH���0ȔIK_#����H�:�P�R�L��&�)AWg�#M��מ�� �p)	�LF���0!�� �J>95؃��&t���i�dI<��dJ^H�ᯑ�e)a�鞏[���T�I.~�0g�4j!2���N%��u���J	?�C�+�mZ͓��=������6�ỻN���.ܾ�f�;"Y}��傟#%eOck�gk�>��\]�@�1I�`5��8LA��Ͻ�>��"� R
R R#��-) �
� ���mO��I��~0L����>o)�P	fT;�+m�A��a$::O;N��݊�TUř��A*|~1>I$�&ή<�Aշw���I%��|%K�#��R��)��`�"�M(�ח�ݖڋ"�g0&��)e6!:�39��Mm��(��$�l/Iy%��x9+.Iۆ���b��~��IU�Z�]s)X�_ER��������� $��O0N�ކ��SJ6BWP�b@I$��ƙ�W�B��$ϒ[�GI��W"��N%eȤv�Δ�qjD@�N�Z�{�ۇ�%���;�u�.�ӯ:x�V̈$�\��bRC�![�g�;iHR��s;1�����"	&U>�2�v ��9I��`�E���H$��X���W}Y�$JA%����2�	+ި�) �1:��x���%#�1[�M��e��m�ɉ	���) �>�W9;�Ha3T*M;�	�k?:ta�v�!Γ��|���]g��{*�	@����)�l�i����osWr�M+A�oc��a���_����w����7߽u����'Ā� ҪСB	H�B��J |m���V��fQA%}Q&|����œ� �.�܃vk���� �un������%�[nZRD��<e#�Ϧw��n3���Uo6�ϥ����sL�%��]��y��I%�φ}+$�t�dWu��Y�x�R^I_mD�	v��ȏK9�Y���@����I)���C��א/a�u(����6kt=�ĸ�.��,��؊J�߂���,��;8��%T��W�H���	��C��Lϒ��s9s���8]/��@ߪbn&���IH�-Sf����I���l�S�Mm�4��HoeD�	 Ruti�(��	�,��gH���+}){�oHN�E�v`�Tx�y��OU����^J����߽�p��$�Y�O�I�Ѧe!4b>M�ܦ�P#�$�3��}}@�#��AI+�׉I$�K�]fRI%�����|�EcS	>��ت_��9����]d�����p��6��y#�O?-|91�\���3��[��B ��-�#~x6��l�[�Ƽ7>@��@��� �l$�'�M��y;g$�%���u�Y�H�T�(�v����f��ztp  ��������!pw��?}OD[}ScZmJh�˄�[pi@�aCt�l�f��v���ʐ)�V�oO=}��#Kj��r��y���A,�~2% %k��	<���M�n��.�����=f���$ձ�}*�����vt��<�3-��4��;	�yi�m��I����4��$o0ng�S�E%�I�ooV�;t*���I/n��fp]�����_�/K0J<�Cf�J�Iy&i��;U�o�c9�x�$��̑"Q^I.w�R%/s]viN��:!��/��yn�'�����S�a$�u�	��A%���g��}�r���.O����K)���1_q(��]�o;2�QI5�̆��L�:)�Rj�5M�1z�6aΤ�j��2�I$����Ov�����:�z��&�!E����U�!�����I)���=��anb�V���L�o{R����}�Z��~�um���*�*�!�8�pwnM�y����[�8�ot�����]�W�x�x�j�e�K���ڸC
�� `5	��(�f �pV�� M�s6�ļ���r�m�M�M,,���&�lݥ��m����c`�6�]9lS=�]c��q�I��+���tiD1�,k������"���͎
���B�ڠu�>��J�Wi�Q`e�̼%M��Ɔ�ģ1�n�v3F=�b� Cu�����̀Rb8f��LY��%��~N��%�g'���܈2�J����$�]�Q&BW��o�"�w���b�ʑ>�P	/*��R��#���1f,If2[��	�%��qu�)��H���S)$���	2�F��Q����r3�G�2��9$�����i*��4��K�)�|�($�������I���}��HomD�Il؛�t���p���7�ڜ͑x�a#X��ŵ���n�(�Ksj$�)��ݷC6�[���_1t�kf��n��ff�����-�יI����`A�X"td��2	/M�r�	 ��ډ2D�~m�yg
�I��~S���>��#�E�ve��pS�B�{;J"��)z����&0�l�����~�K
}�b�\�4�=$�5ʎ�H���	��I{�vD�K}w���t�`@��㔉E����L��r��r����w&D�黑2��#ۛ��\[�"L�gn��c'��c;Uc�i�'�n�;N���%A6g<U`�+4����gh5,Y���ji�?��:�|L���������|}��{��ﱥ$��϶�I2AwӲ �	��%���R%!�>��$��I�5W�gc��"RYӐ$J^Iy)��z���W�$J�ډ2�(.��)\B�<���3�UA)�ν�5!h�.���RIU�<JIG��%�}"e$�s�r��L����k��$�	+O��vwgd��<����dg���g�i[�*�$����K�zD�($���)��˜;��]FJ�lr�����:A��������玲li�+>�NI���."L�,�b��/Jvd���8b���q8��I$ONt	�(�%���g�GM�zu3�A�o7�$�D�+���C/I(�r�ً�f�'�ތYMb���}E��r��	�$�K�;�&|��̏G>&BV)��Ce�C_���Il]�L���)�M
��W"D�H%Oϲ�fd�����A�A�	
6k�Yᩅ��S�U��-.4��������}����/�g�Ny���lK�d�8�"=s��tj�>���i�@( <����n��31�:���Ey$?ц}*d�w,���@i������pe*��Y����5D��+�#�H%{��{NK�^[�n��N%�̀S1��	��
C`pH,��4����B�I+엉I�q�m��~}��S�)2�^Yq`�oz�H����<L>5V֋t�Sl����*h�J�\g�Kf�m��C X;A�=z����$67��8��e�݇�R�I^��K�Rս����o��{�"QA$�"4Ȕ�6�fL]3�UA?N<�I ����Q [[:��h��R	�?F��EΘ�!)�34Q��p�ջ��p�+�c��;�hbv��Ԥ����x��	 ��}�UqvA%��ц	�]�1$�|��� �D��"s˚�� ����h�T��F����\=�R��J�%��H�����~���qpK�}��W�#�n��""��i����.�y�@�Lk�:U��K%���p�A�$���/���tݓ���K����4��Ylr�v����x>T)P�ͯ���;��>.Ns3��p�Y��)��>���D��O��%t�M���~���$�}Q�I�$��bL��^\���=+��s;�D? \1H�,'b\��	q,�7PD\�ie�ʪvcBa�r񨫬�������� ��fA��)�~�&���nK��$��f���)4��6�P�ƍ7r�`�,헃!$(<>�	���v.饤)k�iRI��b��nx��ȉ��
W�I.혒L���g4�$�ɫn�B"NK^Y�Kg�K�&d����z����$D�ƟJA$�:�MsD5��d$��bI3���Hݍd�c�wN��쇺�zh�N�������7D�J�ȵ�橐��f����4�kb�B��NI
�}�!%��u3�Y�H�phQ�j��&��Lvl�摥�$�M�J�$�7Z�yy�3-q��\������3�=��:t���?�����ڟu�w�
�{N��6��V�{Cg��ֻ�یk_{=�V�Hzuq�\�C���	;�3�z_L;�Wd�`�����勴�n��L�#�z��}z����|Gv�!a����g>c���:������y�|7ta��b/�w����9���K5A���ɾj�yvo�yH�L��ۭ��c�<pћ�ەM2;�P�<�����x���î�'q�h�����y2���O���ǯ�D̞>}=^4�3�r�-�r�/�Eɪ������Cc�������w�ý�7�SHn�Z�|������?#�d珷����U�޻�K3Oq�_e{�v*�Y>��Oy]�Q��,#�[c�WX���%�pl��ی��"^��gޤp\��3w�}|��[�\��/.��$$ҁ}��s;�>{���m�u�����r�{{��fұo���	�p��3�
�����mۼ[�����s=СӜq�w�A�V�i>�޺o�	����>�\&i��ڡCƯ���w�śK�����C�G���R����mh��p�ᜃ����y1v{��z	�^�F�|z��o�	�Lu���BF-�1WS�xhk��ů;�����p�޶{�}��[�������S4��'��6�#��MI�r̛�ayT�h5ɶD�^�������dQWN�6����׻��)���=���&�_?dK��8�w�=���l����f��f�tRH���ٯz,�{2
�����YzGW��~��kn�խ\G�v�d�0��?�����6�l��@�y�9$ۭ��N(�j��&���6���f�a�f���H�\ۡ��;"�T�C��$C7/2��D��f�M��A:�3ͷi�.E8�L���=�t�u�:On�,�;�8�����'';mKm'��$s������΂ ڍ�[^g���ge�lL��I��6ȇE���E���3G��ם�{���'N93�"���&��ې�<��r�ם�xtB:F�)� 0r�Im��	��9�k���\^Bf�j׷�ח�NS��/}���{և{v�⃻۶�O0�^֥m��-嗝��e�A�ib�^ݎW�R�g����9v��3���9N�����(�2,	ȃ�c�O;kIݚq*!��ʋm�h�n����-��3������6x��cx���pLrn���\W{k�ۍ�x�D��o* ��8q�^q�mֲrV�ٞAvnNb;S�q���?�j�Y�$��%D��F�EAul�bM�q��M.��]����,�	��c������˓jL6H�MllХ� �.;�x���y��v[�tv�s��	#���&�/h�r�s9�N@ܘod+w�4|�3�;��e��-�D�671�8l\�{q$���,��M��H5�ij˨�P�l�׮0�M�3��Q�����Ζ É�rS��wEhy��,�,�ԧ=���e���#;��
�ԫ6)�4�(�0����we�=0u�E���8��ع��yp��Lm��FjA�0NkA��B]��&�8ݺژ�N'-F����Lr籂�pu�$#��"e�R�
�/D\�Xe{�{^'� B�2�Đ���=k�8X;[�Ԫ��v.�s;'9����K�u�On]�v6@�j���/�.���`��ُ,uq�	tŅnFe�n`N,d�.�:ۚ��q���\c��r+X��=�z�e,aa�tջ7� �ݩ��h��x�=�V�[K� �,��J0�L�l��v§�
�����~'�^�MG#�S'6Z0���V32��2�5;Ù��F�7�Փ�{i��t����R�x�;�sqz5�,i���ss�ZƵ�s�.om�O��6���4��uA��v]�.!.vێ6�]4v^,��\ݠ�"���0�c%b�%�T�����c�;Y��Zm��`2�;p�n��;n�7-�}O 6��Y��t뷹2�G]X��9Q��27c��f�V�m�,�t��|)�3��z뱞!�cnH����S0-�ؗǉ����h���P��5�%�L�qQ�:�a*���g���&n�0s1n��
H�a��{m��"Y�[���a������F�s�q����Z�ێn�Ji�F�ab�ij=�+s-�RXo�lo��4N�J��J��|��=��K�k��gk�"�V�؇�3��ݞ�T�^�c�ݎ�b�hΩ�pp6�x�5zU�Z+,�.1�K�Z���F��� J�]l����f�.v���Ŵ�҃����W	��.�����l][=q'-'`ڹ���������(�up'��ձ����S��mV���"��.�u�a(;p\]���i8��3�2j�+��4f�gۣ�����j���mj�0�n�w�JN��s߿��x~'1D�˿E�-s,�I]s�I"WGF�$շ{j�m��hf�3ʪBI$�n0Ȕ��Ҡ�8N�4�J��eJ�@^��,��gevE�I$��mƙ&RK��� �%[��Tu�Jw��������',���;���)܎2%����J	$�Jܸ�l����y�̕]Ƙ&@Iyt�i�)�[�]�3'�v!�]ډ]�׏ya�����I&||2�It�r��K�/^�L��}�����FT��Y��h.��ݙ�ZB]m-)$[�f�HPa�rY6�N
ܩ!$G��T�Q^Kqt�JK�[ж֖��މ�[�M���b���m�1M�y��\�s`�E�0�a��c��s������ҳ�����w"e$���n�(�f��[�ZRE�ۑ}5v��9"}(��U��ϓ�x72p��Ii�ܦ匄���dى��p���v�Q�@�e�:0�~^o{&��L�I�$%��h�އH����U�����J�{���KOꃻN��p�(9��"��/| �������}w��o4>j�e$��L���T)E���zΑ��̩��Ig	؆�&%�p��	U���H$����חQ���5(�Ѽ�)l?j�J($��t�JHPxp���0p�饧�o�D�����'ih�H$���2Ғ	 ��d^�{�zԄl�R�}�E�^b�����?z��JΙ��IU[�O	��@��x<�����S)$��-!$��n�2����~_~_���F�	[�Y�"pZ��I���f4g���3M�"uM]ċý~�l~��ٝ����i����Q�.�E$�S�)��T��]�v�[�D��)!��u1pX:HpjP��ԉI'섧����!�*CJI%V�����]O��Q%0.�֖�ߓ�y��g�H3L����|����l�"R	$�����<F�u@p�����nM�%��΀eo��~&�s͍�qO]s�W�sI��=��ۛ����J�m����Ɔ�o2Nh^S�����> �O�  �x��5ʪ�D���2��Iy}/����L)��!�'b��Ji�}Z�������H�U\Hp)%���S!7�\�ػ��s���a��Sd�HKC�,\�N坚B�|�R^K��$4��ZS�ܶ%$ׯҤ$�^
1�T�)$;�(*��TF}3���JL
✦H��ݨ��yX�'n�v�j��y��G9����;q�����fp�d�=�1��!#~L)��S)��5��(�����Z�ß�ee[��H(��S) jң�Q`�û3��=l�����5|��;�<`I��n��	 �߱O���]�,�I\'���Ɯ	.��Q���xU*�Pd$M;v�JI%Z_��N��&��%�S^��H�b�JA=ǘ�&p��$�4�觉�7E���y'�R%�B���H���$y�ld1��*;�i�~xU��A�s||�s�1�Wd�֒qQO���{ə�l���Z��;�`���EEs����uC�S����'����L��F��hR�Bao3��L��J[\�3���TLK}���J��x���xn�Ef�Cq�T�䌪w�S(����d$�{{��>�����Wfk���1�!��` ��� y�l�n�;�C�.���g�������j+��}���<�I/%�ےRH$�oLI�����1.��[Y��z��K�k�j�J����S38D^f��c̄�Mqv��9C�y��L�k��P	.w�S $J��$���������王W)��ȳ��Դ�fV�J&٧����%$�	d@T�����6��%*w�S(�@v�ęI{+,$��2 ��B�W=Z{%�Ra-�bq*���II,���L��5��:�q�6�Y4Au<�)�nL�ŝ�Ii��t�>	L[g)��ͯ�`/\PK��P)�tdI���IF�q�S�<�5u>e�b�[}�Y�.��Wj��!�6h�w==��y��Y���@�K���v�e�VK�k��]~�̓s�Lد
�e���`�~������@L�BL��G�1��*���`��L��f�i֭��m&�tY2���ئ8܍zJ�z]���ɶ3Hl�4t�gg�X�1!š¥���k� g�d3C��X���	��s�UX鸼��S^+�[Så���*�<�v����|e�5���(�P���V�II��n����y�5]�q�fH���u��P�MR�Y�	{ů�c�c/|�|�)k�v��t7m7)�;���c��&�m=VM���%'p�~j��r��7���l�D��<JD�$���e+��l݌q��6��{�>�I^̇�R��nb�L��%���ߒ�(��u����"[�����HV���I�^�&R���%v[¹K�*�K1I8D:.^���7L�A"c9��z��Dײ������%�S弴sʬ�D�v���^U�!#T��vLS8!ӹ����T��,�����%��]/$�^{�$�e#���+K��؄�`�&CKE�JK�Ya,pC�DphQ��r��IT����w-l�q�����n�i	$���>�I=�dJ5�N�V�e[k�H�\`a�;�.��ز!Di8� ����G;W#�8f�����	�����/��~s�fv,�H3wya۩�H$��4�t	�H$�28̥b����2Ꟈk��Ȁ�I����'��S7�D�1 J�d�L�~�$��ƻ����ML���J���#Vp�v�usy����AmԀ�EK��u���� X,6{=���Y3��nCY��W��������x�'�� $���X�$"in����7�χlI/NG�$H�c�`��9ɺ6:䑂^; ΂g�#�j�nD�z1��$z���<4�����A{���F7�uibX�pR9y�FFt�]T�o�=�L�fD�A��� H���F�4���=^�$�ML�]����g$g&�u��� �t�H7qC^�ٮ�H����F�� �H��Z��m�8m��<�����`c����c���>���gn���{0Z�r&4�Q�/ߟ=�}��8=�ɚ�I�&���"I#j7�K���>(ڼo;dO�-��O��t��3�I �*�U�L�M8�GXq�9���'ē�φ	��ޙ��W���zη����j����O��ջt"ElgD�I��E�TX��W;q��N��]5��v��N���,p��O�gb�y�T�>�uƨ������<�x�E;~6�����m�ۯ���`��&I��\\���.9�ǉ�>\o�7�%�r�vp����kS4�y*� �e��$A"�w�A ��uԺ"Z ���<HO�VX��@�/��v7���[3���fAԐ��T�`$MFl��'����6r|�زnp�C3�哢V��v-��f{vP�䊌SK���1i�n!���Y<��K�s�,�t�;�=���A��	$-��هql�s��y� �	����Y>��Ν��Y�����Ȑn7;[E��	�����O���3�@#m�d�;���n-A�ݞ�ɬ�k#g����ft�!�Ux)��B��$���}��N^�E{r:|'�.��c"���+�;���h����nm��{���:�I$����|H$sv@�D�������8�!��	zV�q�D����]y�d����Ћ�#����N��CÇW��G0T�.���ʳ-H%�Kˉ�|HA$�A0�|\yם��Og\󗛐���'
d���O�ml�#�͢��R�U�H�驒A �����6�y�~��dd'��lF��vw�oI3���-�F���ݵ����4.�Ͽ��+�q���7;"A%��d7�"u۱Ai~��s�c�ͤn���'Ǽ_ob��:]9gr]�8��=�z�)eW�F�b=���<CewD��G3v(���z���r{�1���Vϵ;���(2p�H3�W�@ۮ��O-�vF�������0$�f�����]�pY��Hz�~����w����ɒ �[�b	����,.YRަtu��w��IƩfZ�]:I��� �9�056��w�H�깒I�n� �:��@���k���(Ġ�UyN}�i����+��n�)�A3�;7M㛧;`E��˫�5�:;[*U6/9��R��d�<|A ޷��e���_~���d�Ҹ��2����t�'���{tk��a�,�����v����smTp����)��S�Cl���ݺm���lob�&�Y�#�0bc���=tTc�ڶX����r�	�ŏru��gǁI7.Ⱦ+����z��1[�%��	ۡQ8۱N\�ї���!�]��oS���\�9�yM�۲��<`⓯�u|����f���8z�	k^�gg�Q�/[���x�_#L���;f{/w���[����:�-����$��#�	#��fA�.K��cT�1���a��N�]̂	����ibX�pQ9x�Ft�� �ݷ��Xò��~�A$�6b�I��t̒n��Xz,8.�ԕ�B�.���)�8���l1"��LI �Yn�##��^�q1N��W�Co!���晐NVO�Yݙ��)�*gM�Ǝa4;��ձ�j�dH!�:���c�m��|XeԠ���,�d�&r�y�@鍹Ikθ�ǽ����t��y��M�3��z�JΊY�:���!"�.�"�?����e���u����a�����	i5ù{�_���.�$�h"V?0&s�c�	}� �mף"T�q���<I5[�2	�7M��N��g
$����O���!A��3N�_��K?���"��#&��}���Ar�V�^��ý����4�S�+�̆���B�tS��@�||A L�3$��^��뽪+Zֹ�_�\��a���W�E�(�;�9�bY�^)���[�	� �칒	fBD�m�S��W�|M��L�B��H�VD�`��Jd�&A�U��Վݏ�|k�&$�*�ng�����|叢�Vɻ�{�nd��ܙ�3�,�8�o)3=�*V�6P���$�L\�F�vL��H^�̂	�l����4��oH���[���Fk���`���уO]a$i�-�̎���v���4��~�}�ni�:�v���fA��"O��=-���ѭ�!����S2	�Wn�O�꘶�dC�I?�dĭ�bOV�3�r�Q��W�s �	��g(�ތ����)z����f��.]"��@�/;d	\gz�ڦ����g�{{t������_���/�$�f�EyXDc"x�$�D3wn��}���K����j�w�څ���Ѿ�|;��mZ�sf������u�`ٶ�����g�{G�Iw7't�h�뱌�3G�K������j+�rg`=�Dr�3���v%W����%�S��}��"���<{����n��_{�������iR<��Ϯ�Y���,N��P�_�k�l�n=�噴!
��q��h�A����!Xi{��{��gx]�XK�����x��{�S���0���{���yx7�z��x��~�ނ
|�+�|_vNp�p	�ϖ�+ߴY�*�}�����?l��,l�=@�+�W���}���[5�N�k}�<��N4����c꧹��z� �Q��Q��k��l2/5�]�g����a��{��CUj�H}�b>Pt=F_l\��,�Cۚ0���*GZ�\��3����X�!%���S�:;u���o'��{}����z��SZ��X6�*{ug:B=G��b�4�v�����=�����V�޲p�~��>9�_o��Ş��4#&�e)t���=;�)�ƭ����_Q֗��adpg��o`L��l��N��؀��mSS���oh[ͩ=�^���=�iZ�G{<�b ���t>�����f�:����{�S�qy�M��~<��ǋx��=����I�x�W�7���!-X��g{�U/"�9��e�5?�r��������^����^��wm�Q9�woq���"Y3����+�˭�I��͈�+,b���v�ǵ���>`�h���>��I�� �s[C�H{g�=,I�'#�]����il�A��*kd�4����,�й����D��]��;>������j��n�J/n��{��m�;���bG�{Y/k\y��E����^׽ǽ�w��m'#�ڼ�|Iq��!$2�6�D9�yZ"ZafYd� ����/��-.���҃��"�j����9%�yz8N����z#��=��ւ�93r����#MHNrG�.��C���'�$��mg8�#��-$�ms��P;�ŶGr8�vNq=��ו�m���{��ρbo�i�H�$��d8BD��I}�8�6�rq��J����xNe�\NU��,�;C�8D9�}�'��9Nr���ߣW�Q�'�	^2��fûBϔ�u�3��S���fuNй�G�I&�+c<E{���+nzewtOo�%�;DL�tO�qn郧rS&q2{D �z��$sx��n^B��$�7r��oL�d]E�PO��u�f˺8tP-�`f��Ľ���0��j��i�&Ѱt��&���|}��6&t��0.9�.=5�	5+z��q}"��e��4�n���v�}�׫�O���S��r��;5�2H2��(Tn��'�����x�	Q�/�Sw��L��Ӱ���n��b��0.�؆�1+6<�ę��Ie����(c)z�f~΢A>�n��r�zD��2��]��(;8S>=�y�׭�G�tG��I>��ِ	'�s�ǵ5솨=��MJi�;a�_\����H���iDQG�{���dQ������ys�������0���(y"f1�c��� �|������ĳ��I����T�$��}q��V����l@o��k� �\oL�I���=���+h�k"�X2rᘧgd����7A���J
���dvv�6m1lH�}����)˳�)��@�v�81$�FdI �Gv�@)��27S�ΰin� ��$���ڙ�1v,���!�5§
��4�6�uPb	�'6/fKx����c��S�D�]j�O��'	:,��!�M{j�H�%�y��H9P#B�Cb: �}\9��"A'�m�d�2n	ݘd�CL����
�ͫ� �utI$���< A휜>oel�f��2g��c2��]��(;�K�&wm��uV�1�Xj�P�=7[�Ky �zc��j�}�3�,k����l��k�m��NA��^h���:b����?�����ߦ+N��)����Y�����hzsbv[Y"~���Ì��9|<K���t�3����ۓ�������:��:k��v�8x��c�V�s���zč�W�l����	0@�D�*�\k���ԍXЉ��[���vrZ�L��i���[7ȺƉ�,��I����;s�T�x���.
E�k
6��^����n��!/j23c��#]���>Y�Y�����MHBٲj�K�J��)pa�;m*m�y|!s������E���`6��T�>��?�CJ�5�Ȯ���{F�v�own��7��ʙ$㻑 A�WDu�	�;����=i�J|�9��!��;6��� E+1�l��ZsGy!qa�3�2p��������4��c���j����	���DN�=��{�!:)8g.�3�軚̙U�_���p7�� q�$ތ��g(g|I�����<ɴ3; ]ݙ�Tf��$���3�+Pm���[8��`	�<���W��1�_�B	�;!�i.�1�q�uؖ��㵷f�.�����گ������ar���G7��|k�#�Hn�d����~hr3*�ru���z<E>=�'��ZB	�pY��Ȏ�ِI���hoeV�Vic���+=f�{�B#Jޡh7!�.��.�����������g^@��~꼷����G}����\����~���A ���D��d��d��x���
����;�`�3����v�D�]���	��8�ÄW�=Q�^H�h0I#�zfA>ʌ-��œ�f��Ѽw@����@:�'."�>$\GTψ>=�iaּ���W&r<`�ӊ�/MN�����D��fj,��������ȷg��D�u� �U�S ��\xGk�3<�p��;��8wA��wV�ô<ru��NMS���E5G�lvJ2�����<��.�̃@��4�`1��ى���s�����q?*���ّ5.����.Sr�>=[p ������f����WoC�B�v�f$|{��@%�9��Y�b^�9ʽkP	�EU��p�"�'/3�Ƚ�'�Wm�|H>�oW>Ɨ|P�:�CEOw<շ���&�]�i��cV2֤�1��ߧ���:�����v�0y���j�1:i�h[UɟL�=�N}X���$}x���<�>?}�U�)�wN�&gb�'�喢�-�W}~�.�A {��� ��:b˅�����θ�HwZ[�ӂ��`\S�Tf_`A��.�"oq��\�`L�eL��H|��<H�n��:�Ã���'t���ݝ"�5�6��ۨ�1܄e���<�u�����ۖ�x>��gA'%� K@�S�S$ݸ�I�n� �DE�i6F��bǾ�����8˃�;�]�:���zY\�~� �A��x�zb���ق���v_>�.a��\�r�':�|zV\ ��O�I�N���� �|�\��u�=�䋂�X9x�NGd�x����M�$ʨ�	;+y@$�2��t����x���fm#���:�r����D6�S>���
��a{�,�V1U��l�����%�� ��5o[��۸�䋈Q/L���{����|F�,��I����G_�P[#{+����5�$4��x�ʮP	9[��>fQ᭹�G��y�=Oկ��M����n��cbjZ��T�	�H:�n8�8��:ʹwq������E�����<^6�<D��1=���L��{Oe\��>ǄH�m�&���t2�X��Ge��n������W�L����N�o@�ӹ9ŷA��U���;3�A�Ӡ� ���`L�nD�_�ʱ{��lk��en�D�v��GToL�jD�if,�f�|s�ۇ��Mc�W��ĂF�_H�H7�uV�JyY�3��fxP	���A� X9~�ߩ�zd�7."ܘ����"+X�$N�t�'�7�p{�-��2�*s��k�m��uO-8�{'�`]V�vq��gw�w;�6/}��jw�m|ɍ��p���ܓ�6�32��jv���U*�ʭ��$ࡓ�{���ؙ� Y�)�t��8^���v�qn��ӈ��Y3���G����1�;v}�c��ڔ7mf����v�#Ϋ�R����]<��-�km��B6k��.�b���k�q���I����W 9�[A7;\�|�t�{H`�.��I+��4e���JJ�����
�+�K�7kv�m�nw���:��\����[��:��k2�n�s�a0�f`�u�uV]U�dX����>�b�d�Ma:]�;b6�;�xF,��b�gc�P�y�>=q�	^���<�ZUv���x���$Te�r�ܗ%��6�D����@�����kF��u���� ��}�,�3j�k���`�e�a\�Ii�����A���y33��+_�Sz���O���d��\Aǚe�ٝ����y[�;Qj�ݓ)uvTɾ�E�^Ǥ/+"$���M{�sC��W:8nn��'6�Sif,�fŠU�}�"H���C��2�,�ǣ��}�w� �.�`@$����z���/qpw]�֥�HP,��8n��G���M/X��;�ѡ�l�=�3���ۦ�%8.���A� ȹxչ2$gV@��I�l�1\�ю5�>����I>;�� ��~�S.$��̞�Q|}狱�#��1�����9�9f_�Ѥs�o���M�=����8��X�W2˞���̾	&^R���yo0�)s�����3�$�OutAt�|���S#3��ES��.\;�Y��.Cv��eoCJy(F3YUƉ���)�ϲo"�>�l�"�#Pb� �bL�����(��et����Lyz�V(� ���Ֆ�A�m��[��@4�趜e�ٝ����yY�Đgc�$���u�t3� M�t$\��Iˍ��!i�6vz��Y�_pv��+1�ؤd��9U��	Խ]˻;�B�tt�.̩=��}��R۱����[��U��MtoLzB��FK�1�K,��+= �2[9@$dW_��E��Nt�p�&gjk^I=���k��g�ʩ$�sk��k��fA�$̝�@�U
���|H>�n!�}4���nk�.��Kૺ17	��vv����4\���n፳�t�{����;�#��ܲ�p�=��M��Z:�য�@�v! ���D�=^{�n$1-DmS�Y2�s�����ė�Ss�"H뾞���מh���{P�F�3����-U�>'ăy}{n����H�kD(�7�rd�@;��#����f��>v#u��.�9.ٺ�)͈�v�p�sX�d�(�u�/J��M�`j˿y��]��݁�]���� 0>;w���(�,���)P��{w-ٲ�*�z$�ؙm,̉,]�d�&�5t�[�#��.�(v�U�ĐH��ɒI=���@>�������b9Ψ?�|z��A� ��xYs2�m�� ��K�^N������ ���}CM{}l�8d�ĸ�إ�_;m��'Dv�9��{q$�H&�� �@�S����l�h�B�4�LΧ�Mᇙ��&	i��v��:0�;mfгԫN�]1m�HX�5"&�#E�Yg-A�%FV�:�g����̙���.郳���<�A�ڈ$I������U�h�=U��|I���>���6_{��1�Sh�s�L
w(����x�\�'�u˵�SJ$WY�6Ɉ�4�q�$�^�\���LA]�ww2O���O�����"�P"ס��d�	����q;Iݝ݂	ܺ�4�|\]P�G/j����x�Ux�#S�4��2���tK�C5���e��%���4�؂I���;�X��/a;�Eǫ��(	{1�5=�A#b��(8/�:3�Y�"�ej���'�Z�DyQ���V�Od�����T4X���{��fA�fd]�9P��:�r'������F����Ȃ���GgOH�=����=�>�;�����:��<�]��h��=�����N�6��'��lS7TKq�^�ؽ��7�k���4q�_TU�i}�q����w�2�w�?�j/_8���̙쫚�g͒�31d��^FM���u��R��D����S/Y��}�"O�;�Gݰx��w]�y��緀�U���>�Ȟy5zbK}����{��g|���~~���%�/k��PtIǋX6ʖw#|}�x��[��[���>�O*-�01,�቎��;
W���#c�]<�#ҋ:�R'�Ձ/9��M|[N�T���i�'a�>þs��O=k�7G�����;����-��ރ-}��D!�g����r�Yj>|�����}�վ�	�2�2f矏��M�j/;���N�o�ud��8GN\������W�}��N/v���ۯ��\	�=S��="O�oa |�?yϰ��]'�X��w���;7,���C4�6��	f�9��v/{|�l{�o�;�u����hǊ��{��Y�jxpVp;>ܼgXϞ5�;�v���	�7='�����!�����:Ao�"��i���xx�ӽ2�d��f�Oop��1�a�O{��簧,�}�#(��,]�6?iM�X:�����C|6��c����h�&�={X�&����Ae�`{ɽ���ǣ�O��o_��r��7���~ֱ��fn���'wM�.������:9m��F+��Y�\��]+g�S����o���;X8���Ce���8���ϻ}�^�#�0g]�{���;��f5񵩽�T��u�>�/o�
��5����әnC�{d9B"+�D�0��������C�8����ۭ�98=�=�-�Vې������9.Hs�� ��X>��X8��y�QtH��죩|�@r9RI�'���3On�s��8 �Hr���g�����.��{n>��;;f=��G�Ӻ��ÛY|��p�;ΰ�����^e�J88�vs��#�z��rU|�����������A�Qm�n�S�r)�3�)/�r��d�A��$�)*&"���j]ЙgA$wiiR^ZH�%�B�yՑ�ۇ R�3�(����H'��q��l�����mÜT�{�� ����ն�8L��m�RG�7�t����g2x�!�խ�[#`���pUpv�3��
ݤ�ˠ�î1�<�׃3��)�v�WM�۠3v9*���{Cy����i��p�
td�@y�Q�+�-��4`���b�-��\j���sgk4]Zr�%���j�H��<m����M�I]s)�Ќ��^����:��?#�v
�O�( �r�[ݹ9�ۉ���'�n8��+:�s��ܞ#�7d �s�9�#��p�^H��=���lݛv��]`���u\�����l�gs�Ͷ� I)�MgV8-��Af���h9�.3�N+�v����6ϣ�ʒ�9n�[��>�B>�+�lL���M�m0dҩ�Ys� "o'd��њ���w��m�k��k:^�/=Wbh���k]�������&�����X�l��r���ۺ�]6�ض����l#�x���l����$����Ob0�ۜ�
���!B��d�&E�׶m��MF��cb��tvwG<9�Unk�Zx��n.n5����g�l>޶��ɸG���En��H����tv5�R�V�t�=͒�}��wM��wϋy�H�qb:��+��c��Pq��f`m��Y,�]1��
R��۱�͍�LÞ�mV��P��vyx#O1���l�[JA&F��W�[�����㱎�Э@sj+�h�n��\U�6��V����BMiԐ#f�˂�3x�)խ�M�D�v:;Y�:�;`d�Ȍ�-� �ؖ\���=fm������`��<`�V�Jn]1]G�M6D,5�2�GR��j�3�(��8�,`���N��}�6����-��ݺ{z�M�v�rP�l��p�x���DwP��̨�y����K,(%�q"؉I�5_PM�G^ԁ���=Ü%ؚ�Rbɭ&��4�v㶪�&g���^����] .İ%f�1�4q1���	u1�D���+�8���m�����V�C]a��7�r�(j,�խ�$X^u@4��Pz�v�-q�+ƛ.�@'f��h�k��Jsn�5�Y��JZl�5E^YM���GS<Wk�7	�܅y^3id�8}���]!.ޞ�_�����g�	 �Лg�Dϭv��F��!̎샃�d���sq�\ҕ[I�-έ�=s�/0#ėn|����yị/!Lö卑�Z'����e��������1k�=���>Ѵ����v1kV������v�,�l�	[/>��8�k�����q�Lw�p�v`��wd��������f��=��̬�M�X�v; @&�W0����\���E�P/��ّ��k:<���;/0|I�� ϊ�]9��aQ�n�g'p>�{�wgd��]��s;������W@�Och��!��d�v�'f�w:z'ć���3"Y2x��Y��-;.hf�x��$[��'ě��[���i��~N.�h'cn�(9/�:2�Y�$�r{ F��m��i��`���<H'�'&A>�s����F�x��~������3A0ͷU)qn��`牧R;���RcB�;<�66e�����>ϵY�VN����G��OnND�|n7��o-7X�c�m�kvzD�&��md��̝�̂��>�F�[�iz%$:n/w�����ڻ��j�,��|c>C�x��V�n�����d���s�t������r��{�f�Of�L�&8��6��A=�92	"����d˟���bͩ��}����v`�dT��Tz�Ft@>2�<�7D
�͊k띙�.;����vgd�"�܇�.g{��]<&�k�I���D�H�Y����5��ϵ�>9p,ŊA�̞$���� ����#�s`PyO����>'�#r= ���ڕ�H0��Wdɉ���/h2� �V8�ї5���Y�;E����m�xk�h73���L�����JK��N���� �r7 >$��J~4�(�����C���38!3�%L�9Q�&���AS4󔘽��\P ��{<H'��4�=Z�^{k�8��g�����c��r�2w�2gT$�3�	����<��n�&EF�)Y,�m<��~��/-o���ug�{}�֭�>ܕ�n��[����n�ʭ�E���&ao�S6C��y���A6�� �o�6����f	fEL�]����s�R���v �NKw/GloN)�Y��F�����n�s���������&%f��ToD���x��l��CX���	�9֣Ă}�� �Ή|V`¶�Ѻ�9d�jɝ�$d�jX��c:�eݜXy�v'l��3� s��+�.�Y�$�?�<
�[{�GB��1$���&�cy�q�&rA�ڈơ^��	Aˢt�<�M�L����r������3�}p��@z3�A �����*��Al���fg&r䩓��!� �E�I"�3���U�K�Rm���;c:g��&����r�3�˙<�*���b�`�u\�����ޙ1���<�Ɏ��v�T��N�X͞��}ջ2�!��'�|O�]9ڸ���(��7�g,닳��C)��ѪQZ�oߝ�bŉ���2��A6��C�f	fEL����$�o#��B��Y�6�V;N(4yF�O����}�1�������C���5�ܦ��sutr�ӻ�DӗoFi8��58�ۓr��H�5��pvr�8!�}�id@b{��_bH ;#�<m��K���J�o��zl8׳2H���`������L�tA-��s	l��G��'�b{�#��ɑ �������Ձٞ��K	Cc��+��]��z�
�ޑ �{c`A��#HT��y�꬘Y�A��ؒ	܎�5Q��g&r��^���:v�,��̉��}|�	�=��.���<T���S �eM�A���S�vys'^�D�ކ�����,�O����$M��@ �69A���4]�۹hT\�L,�OsJ�
����'�m��40d'7`�6�+��]�����\�}�h�����o6�ݭoVk�`N��:g6���p�D��4ݻQx�ǫ\�Xu�i�5����������wJL�i�T��њb�:ǰL�$T[GK�ܝ�'	G�]���na��6B;�F북عN2�8��p���f��:��;��:���ަ@��eT(�֫�m�'\F����K��ѷM�l�G{�N㹣{sKY'jݡ�q�uQ��ݝc�c7T�p��س�D�g�n�k�D9"m�	v,&�-��E�.�/����r��	,ȯ��ڹ����l�;=�cjz��kj./đ��r-t�L��b��!�o_�fj�+��@�I5ϰN��B )�k�.yi�w�Ċa*8/�w�񞭈 ��Я!�o_�t#�y��	>�l��]7|I^w$�N�P��������͊=�1�$��PH'�e�*�ٵ�ػ�$��v��Y;�9pT�/a�><�y	]�>����t�F�L@$�ת	�s�l�/q:�".��V���Ðڱ���Qlı�gAkk\a+�a���b�#rs���:��!�wH;:~s��=|3ʥ7G��H�����뤓sz�Dz<f9@$S�bo9vw$dT϶��g�<}�q����{Q�%]b>�9�g gʛA���֚r�Z�ʦtfu+^�ݛ/P.}5i\5)�{�Of�L���{�+s��y���s�������?�ƿ�!���> ������53���Ţ��9E�L��L���%v�>N��$�H0��uL���~ �6b�I!�{fM0�n	���.� �Ol�{ݔ*���$�j!��ݙ$z߱s���K<��~0OF֒W��ݙ����l�'�v>;��v�4�Y���ތL��L�A�� �yl�1o�j4�Rgv.�`�Ʃ�kCc`��ql�R	R̓6Z9řMPf�3k���UZ�JN��\�����$�Ϸ� �g�$��D�Uv���|�Ó�d@'���A#*9���tBwu.d����S�f�뫆zGēo��$��u��=5,��rn�8	Q��.��̊��e��P$�q��A$�#�&@��d����ն�~Q;n�"_�"���q٨����w�ͥ�j=nG����K�mw���w#�+!/���Qr�+uC���YQ=g�&�{"A�gG��ȵ<���C��	�U���M���ʥ�����I ����s��ٌnyB;+k	>���O0�lE��:,]�A�� ��m��cp���v۱��	U]s$�
�ȀI��`QS�u<Ъi%�
Oқ0��\C;X�Ä���::�w�cO�Sl�X;3�Jvt��a%yܒY;�:7&#�>$�́����<q�Xl�*��j_��A�݁L�Z�JN����%�y�\������+�s�(�5Oф�HW�	�z�K�	�z{9F^�W���h�I�u���>~�NK�e8�\p�5V	�/�vS|k�b�[�	�f�g/es��g��'Ă������<O��5��S��
dT��雩[N�ǤO�x�oG�4�ٝ������\�̫����>�.��=rU���X���U�xٚ�|Ȝ7��Y�ԛr�@�h��x#��23�~��n��ңx�@zÁ�����a���C�pTH3<�Dx���IM]M/M.q`j��A#��L	�vwL��Gx�jiɍ�XL;�$�)��w.c6�1��� <���FB^4,Q�Y���-�|�^ߍcH����Q��A�{l�A�;�S�kMt���°*g��� �%��ǉ��P�W��C'b�T2��d�j�DS��	��`n��@0�d�e��{�MV��g�L�P*��D�}� H.ҧ��2y-�1ϖO�"]���KnwL��2vX�	�t���l��sL��c�]p���$De����K�gtl�j,��xP%����T���t�����gknd�	/y�#��9��l�i�:>7Z�|Z�z$H/��#޻MO��{�w�a���[:׻bآ�5_T�f�ӕ�#$:M��*���77��:�j���^�� �#���A!IX��j~XB��@�g/v��Wc]��se�թ浑nP뱭E�����+�A�Ӎn��Ї��nX-rV�'��ẞ�.�]�b�n8�Q�;1e��Vb'�[�v9��u�¥�A�,6�L�����5���<��]�s�z�P#����#�L���FGj������xՎ�t\�\ڎ��.sή���8O7	�՞nٷ��k�^㮫�bzz�h��6�Tc�5v��Gbh;����^]l�<}~�q��;��v
��2�Tx�ӷ� �@$tgDӋ��o7o�v�,���	�\���,"�哳��5��l,ɑ�K���[��d�A�Ώ�u�������ǲT�6*��y������OL�	=���Z�y�۬�[J�@&���A>$��OukA)���`���s�q�r����ʊ�����OKg,k�Y�������$,��<�ñ/�Ni�CQ�ʁ�ʥoKvj�Wk���wcu+G3�L��;�� H�m��b�ͻF;��a=����ܔqm��ۤ�2]� �.�mWe�*\kL�M9��5f��.�����:N�I�]�5�>�����|:[9
����u�Ȋ��M�l#$�3hfv���S&eo/x3�x���@����ٹ�AÌ
ۚ[W"sR�K�y?BY�Ni�ױ /�k{���^�u$�l��bE��k=s�����u�/	]Y;-��ǒL�M�3�~��V<����y�&۝�d�8v.�2����l�c�u��aJ̨��w��$jFڶ ���	���rd����d���]��1NW���x� ��Y�A�\oOa�<FU�`�uwC]Ћ'��%#�Y͏���$�����`�x;�\�ǉ�� Hq�"W<�[�F�	s7��t�Ŝ3�\�a���h��[q�=�u�cf��\̺*����t���1�r\0:s�6�p�I���0@2�d��N���6Fֿ�S���~1�W��.�8H'%�F�WL���ޜg�׷d��T4�@$�d���u�t� �W֋^\�;�4!;�a��%�go3�!�L�3��� ��$h���|}~�g����y��?����4�+��Rə�K�m�gj�wja����6���̖�"�C`��wWn{��T;���-C�u�i�~ٺ*f�y\]�D2??w�����(�G��e�{�8���k�!�\\� ��9�w����_wn&�z�mKN4��|��n�o�o�v]������5��k�/\y޽uf�׺�R�x�k܄�S��z���ܝ�^u���
��(�Ny�{�t[;�S����-햁��s��:�Y3���ǨϪ��{��{�s^z\��8&��b{�N�T�	�d�4xjLx�2oɝƎ{���Y��:jgx�9�z8z����S7�J�{����t�%�h͈�p���|o���������7��
�ys`��{����g&����h[�o�����Yz�����wP8wۺ�j��;� rC����f��N�˺b��k����:z�Q!�Ky�{77ٰ�t	F����k�rc��4 ����_�ut�V�K}w���+�4w���#!n{;�s<�/j���c~H�)˔[�9�ݹ2;|�w=������:ƴv�ϱ����E����!��ã��4on\c���"��6�n�7oP��p
���g	n3��#����I�}���o�����x����^\�>Z�>t���S�?]��9�E�׉'���.{���o�����m�G��8C��/��|HפyS�4��� �g���������EL�Sp�S����0�E	ヸg_� ���Hs�~4�٘fF0��1�s���oy���g���%���E�����m���qGFbNArr]#�m�~[RD�˼��{cmΟ���EYn�ܳ�w�GϽ��M�q�'��δ�kI�ۻ8��[�n�<��B��L쳢7:(���/�Rp�DY���C���k.�mq�Z�qـ\[�x�2��4���q΄�tQqu�� �8�#��RW���:����ۯ���I��A�۳����q�D�9%�t�����++�^�AՒm����2� ��>�W���v��wg�h�#���+��D^���rp���t%�m֯;�#��J̢N����;�:ĺ/�u���|�L����6��N:��w�E�y�i�tf���jB�֔^�m�d+gg��KA"�LGdwL�MLJf�%�pᙞdy��c-�#���d �$uE�ɿ �S���Kbe_���$��h^8b�}�P�Ω�I9=�jWS��]�oq��'Ǯ;bLx�m���oOG�����y�~���J��֚X5�:��]fH1�BPus]˴���YA��~���B��SdW�g<H:�}I\oD�$4��:Y�_�x��z̑!�X�9p�?�5&�F��G�E��[.�ѷO�x�p�E=�L�`��8���^�L.��6O��F�ĺ.ࠜ�oOKOE�I'#9��pw5]�9S-�P/�A$\o<d���)��:v!�����u�m.�&�	&^�O�GtA�-���ݘ��LWS��](g���m��E��	�Z��Kݔi2M��^�~6{oq��\aq\�T6u����ӻUN-��>ˣ��<a�)��4*<_32gĊٚL���d�&g�T��A� �yg�=�r������I ����:[9@-�Ʈ�n�k�H� ��:fI"�9�<���p;l�8un�԰�C��D�x�Mjv݊�������i,Hp�`�{1�'� �@$l�r�dt@<���WE��A�� �g� ��Ř�"�A�U��s�,����5��,�	�� H-���1�����Qk��9Wu��LΚCO�|��[��A�|���j�f{ j�����	-|�h$]��K��
	�i����W�i��Vq{4�}�$d�j�A#�g�ؽ8F?5׉1q�%���d��Kę���'�w�bM9�1�����a�=1]	${e�_�'[g�O��vY��KL2�4���r����ev���1�2�㙶���^�c �5��o�P9J������m�b���5J�D0J��K=�4�NC5$	`��;7�hvC���c�$�U�Zd�`Z&��ι���GsA��a=�m���9{�q��|��;Lo=w8�
����4\,ɵ�;l[���.+v�.�:|R^{Dkvnn�k[�ر�$�SCn����Eź��n+n���Ԓ��8_\�{Z���D��y�#+�,ix��q\��uLJ�=vI�d�^Wv�Oj�zD;:���X��T��s�+��]XJ�[j?������_�X�w%ó���^1�ăҳ�H���Q6���z�L�@ ���P	C��Ĺ,QN^c�f0�i843j�1�p	�Y�>;��H2��2�Qcr�����k�B�fg �gf*P�3�1�W��I7���������$̫��guL����Æ�viM%�9�N%�
}�m#�䁈[�Ē}[�3$�	��>�{�\�B�$��oב8�ໂ�9-US=s>$rs�Ѻ;���#���x�3�fD�A���l��D�����抃��!�p��s���sM��	��杳/kIe�g�"��x�3;�Ò���J܀���ē�|n{��U%N������@���ɑ"�̱����Pvy�� �c߇���������xv�W�*�7�8Xr�ڵ/_����T����yo�{|�3��ō�`�\�����V�g�E���ڊ�A��@ ����ä��=Դ����b�(��މ��ɐI ��0��f0����d�/{&D��ވ!��E��������؞�k����Z�'[%��)��*�y KV�G�&��M��::�4vD�}C��rჹ��DX1}Q� ����j��3�/]�	 �]\��'�-֠�ܪ���'�����MӚ<$9�,h�.�z��g '[��B��㶞�؄�.�n �,�NK@�ڮ�I�A>�n�/��0Cc�V�����Au� ��cpt���NK���]���!�-���=�I>$��]	 ��hG�!���'j�3�T���DK��,�]9Oh��	�f�޼��~ILL�h<C�&5�8I�}YI�'?��Hj�����y�s��"k�}��g���O�gc܋�`7˵���.��՘��k���@Net@'�u��7S�4]��T�VÈD5�s<����n��$����2���0��"0�k6�$��@��<M2fK�vd�|b�Bھ��k}bl�ы*ؘ��|c˓V���1&e���|O#�t7X�]FM�K4eu�`��71��j#��^�K�&Lř���|�ˆ�;��������PI>��ʾ趤r�T�m�0�}'�-ڠ]�����
�mWd��������T=�I-������TH$k��ލ�S�������c�C����
�4��$��ځ$<OYg�M'z�sA%�����w:*dԇ�+�.Sw!<IɎ��c�짞 ��qA]���$�ok�{k����\F8I�g����Ӿ���7~��M_�j����3�۾ˈ�Ҙ| V���X�t�a�ԩ����� �]�m� &2���C�\��z�
n��$�v\C�V>�H=��A �[�Q$�M�\Gm^���F����yk�2��b�U���4�YqJFP���ֶ;!f�Y�L�m�|��K�VK�vd��ک�į ��j$�|oz���lnj�3oR�J� ��TI5���k���3��F:z=�1���,�� O�/�D�}�	�qt�m�.�i;��\��ೂ��-{1��&|H$�u�N̪ev�-�˅��ʙ �H7�p ��r�	wr��g��"V�@�=�.x�r�$A9�q$�\�(�n���a�����D�Z.Y3��@���zVdd�%��@���D�=ԉ�}�e_(�/z�F�w]��|�{TPI�x�Jv.�&lI�L��!�����l�@_�K D�����N#��n
�#��0�g���N�����-k�/���WB��'��J^6�����vwm6B	]t%%�B�V1�Uv�� �>%�^XӔ�k�LV�X�m1�uqX���G��8[���T�"ęr۷n��D�Ӌ������дe[)�t������o�2ܻ6��O/k�᪫bsc/�N���݌�*l �9�Ŷ���� B8,F8��%�� |�g�÷	�9��W�j����<��ؽv�z�G7>3��xj�� ���%3n��%عH�('~�ۙ� ����	'�-|�����:k\�z����+v`C�
�,\���@;N%�	���Ek�{��$�O�gLA>'�-ؼw���l��vH���K]�0;�p�"+�:p�@&�wG�Y^��M�=�� I's�� l�b�	��Pr\&pX�z*�]�w�کS�^�#��H'%��^�{q��v���A���*��Y�'rY�x"Vvx4���H8�Sw����l�WE�a�#�: G��u� �Fk�L��k"���E��~��B�U�g�
�G��].�*���;.�-%��b�*M����S�߷��ŗZ�Y��������W��&����c:d��gv���~�*�= �F�n(�$
��:.Y�2��̂ x���[]\��Qx낳!v�@2�G�!�rV��2�7W�ĭ�U�#cز��n�"��E^N�DW|��_� z��[rmC7��=��{��7�}r�j	��A&�!F�.Н���"lh)Pb�fv*d�(� ���H�H��,��;w	'�-��y��d쭆K]��p�a�(y/�sW���Cʮ�ċ�6z�7���3=ύ�WbբxW���g��lI��fp����U����ޘ���Ƹ�y��D�ݲ�	��ْA �t����ﾟ���Λ��?#0��R�$2�膇[��tܮ�
dmm�pg�T�ŷ?�ϭ���QM���%f����	�$}��C�i!�6H��n8H'��q ����X��CD�����+S���ӗ8�ȒO���L�(�u8��1�����l�oY)�tȸ)y���$�ɇ�@�;��pSl���E�eU���v��cȬv����	�!�Yܜk��/vni�l������Y��7Fr̧w��Y4�3&�Mv�Y�ϋ�$�m͙�$o�#м��
T�tS;� �(�zWׅ�ĥSI%�;"A>'��!��N�v���y�Q���b�G���� �*�R�;;�EC�Q"(��@��]��g���ȷ`�2q��H�� �@�n�D��C���,�lAe�I'b]]�E��ۛ����]�e�n)��tamVŉ���_�����tɜ37pꝹ�I �lD	�ݨdc�׍j�T�t�#�"�����$��w�h�♆%��K�;���6�鈲	#sb vWj�AxL�w'�Z�|MK�6]\�L�w�U]1� �@�W�@6����z��pN^D@ ���PH��p왋��w����|�P�:3[l��A�K_(�}�{���gl���Jw����2{�G���=��0G�q�rL�w0s��ve��!����}��̹ǳ&�������&��COP'����-�ĪE��	3�irb��y�2$��UՂr�b<	�>�;� ��dO�V���ޛ�����N��)�S��S&a���3�Z���9��#ڢ˛�݊� ���gVO^�����nN��h~/�n ɜ�|O�{&|o�+�s�9`��M�� l��A2�c��&p�p�>�깟ɻ\�r�0�f� �-M�A �~�!��À��n�N�7I;����xc:ÐI��ؒA&�P��Lk�3Ae�g�$�� �T�]!�%�	�Τd�L�5E/�
�w,��y2I���]?Y�|>:K�<��0Xvt2pJ�>�����!i-�y��䃶H�l�H���y����88�\pt���{t��뺾_/�����
���dw8c�%xNǚ��^*�\��v���%�I��5p���{N����zA��s��Ӽ|6	ހ��8a%�����X\;<�c')����Ag5��h�`�gN�l����[�h7��hW+���{%���]O<��q�`��Sh��������;Go���y۾>���p���g�7��{�Ѷ����+�����U��+�lgv��B<�ɻ��W�v�l	���5�:w<�|��;���gx��ppgӣ��Y�vy3;���]��>�V�\ԏl)����QXC������G<3�������^�=�nL�W�ȟc���&o3��;�b�>X
�;Ӽ�x�׳7��|�g����k9-�����b W-�\��!���s6� �Y���|W��,�����Oo����:�a���tgB�+j�N�9��z���z<�j�s���&x��*�/�9&m}'��x\�2KO �
o��{f�x4�I/��S��0���%�\����v�y�vz�>z����9xM.L?)�ޤM��F{�m1Ih�{�i�	������!�t�b�Q�#�e­����◤KG��>�d���>�X4�}�wPnE�٥YN�A������H����;6d
�ܽ�Qg^u����\`��N��l�Ϸ�Ld�^�f@��'�?.�o����������� ��/_��ؼ�]0����.���guX��<4�&�^��05�+G�5�~ɷ'�r��{|�C
��}��(;F�'�JA�i��x��S/�F�,Q�  H�q�����I9vYvpT�IOoO#�/<�:;˼�����+۷Zv!Qߚ΋���q��u���E�]��+�N#��e��G^Y�wy՝��y��{��ާ����۬�fC�;�ռ�?-W��kj˶��qZ�&k��SnL�,�����#;������Yy�e���}�_�v�w[n�N��ݝ�E-��g6IɃiJK��������Y�rGY�ZG�Ԗvٴql�-�,���⣻�y��i�;��Ց�v7�׶��3Ȣ���r�����7�p�&Vyzyya'eD��N���Cμ��Z��Gg��8+/.Kʊ;m֕�(V6���w��Giw�=�'���m����5�j۲���Ő�_���_��k|`�]Ku��cf+�uΜT�+=5԰)l�ڥ�.�8���&X�ɇ6P��������]�)/2�̤���i�B`RMi�WR"�Y����[c����`�i@�]�\tf;ci��M;��Ϋt"h��2�,έ�f���/�s磰Q��C*[p=d��'����;�a�8J�j X�K�W�YYf�^:���:��V�FU�(Y��6j�҄i���dWyz�Vx1��q����� �g���`9u�����G;�<Nb��� �M8����/<�'n�xGma�����X�oN�X����qJ�ы���"R�P6F,:��3i��K�B��Fa�,OV����Ƒ+\�X�/Dj��y�[b����q�r=��ˮ�^����2����Һa�����3��ݲk��p��c��W��%yr��wn����*R=	=á��-ٗ^������]�x����3e5���J��n]�S���������b�{<Js΢M5m2�iaf�&�E�s3,�j�X���d��"m�(a�&�0tQֈ���t���k+.�b5�,qw2V�7\��G���T!gq�rg�w8�����"R)T-�CJV
�K�I�-W]u�jc��M��q��^5��P��������5شl��zL�5���<0�I��N�)�1��]
XC�M��[���CF�n��&����������W$��{/�G��xݮK�ڝY�p���nI�Z�Tq���M�:1����;lm�����C�6t@9��YRP5 m���^��ccӅ����4vX�K��ް�qh�\v�*٬�Д�Жv ����MI�hq�]=\�u�q��60�F�ۥK�=��U�����Ke7�v��	�c�7����b�XBՕ�14i�d��#��v�d�@qm�ͻ45UIӎ������N]7�݆�����z�Ô 	��)Uj�Wfc���B5�����5�m �,"Шm%ł��;D��k3^T����1-��9R�K�M踪{#P�Rh9}A�k]6���Xm�fev[nK�|��#�&�"�JX^ۢ��
�lW獨< ֱ��tEtp��,T�M6��5�T�5j0��f��-̢��X=��ت0r����X_��{�g�F�uЇ�坢�u�!.	��N;7=]v�bz	�ƶ����M���.ѳ����^�2vw$����+�gE�L�?~x֪�|IތȐ&���6�u�G�˫h� u� +�zwvt���:hz/я��n�q��{a�ʲ���r�rg���ވ�y�
kY�<Y�C_��ͭ\>����;��!�L��\��A��x �.���D;C1r�qJA tfO���n��;���ix���*�KB��f26'���tDx�F�_&�|2/��#�s p����0(�:���p|H�fG�@��7�����vjb|	#�b< �Ci����,gt7]��~c�3���n�oEφ
�����)WZڡ8�h�m%��6]����}|���E��;��[�8���@'���u��JG�}ss$�|v�"ƫR�]�D3��T�P�}�Λ���11e�&��5I��ʕc�olo��8��cKn�i����,��i��<�i=��N����pk ۉ�V0j�f��z��oy�	�$
���A�7� �<��������S�:�wIX�gwvL��C绂D��h$�O6�Ψ����$�]� G��/*��Յ$�f���+թ��`Y5��n��I=-\��vLH'H��� LE�j� ��s�fI�Iܖ�%v�|I��ؐN�r|��Tu��^'�-���w��\�a�ߠo�Z�i�WM�Snn��C�i���[/��=Q����qӒK,w0���S���K�W�7W0 �@9+2<�	���T�-�{�g�<@�NJ�PJ��cl��&N	p��T�f̂;"+;���L�v��6Z�����v�5lZꋂ�x�L];3���y��3�>=�9I>�	7Z�c��;إ.���W�t�q�`2�������K���ȏ��J~�ӛy<�wv]݌��ܢ*�Z[q�*�ML�4`ler���lr�kvjz<H9+q@��Ӓ%�ͤ�k�;�A�;R���N7q�1t��,�7�Q0�FwN̂A ��^蠸4���J?�L��wv0g�N�E̟��D����м�~�o�ңĂn�zD�I��zk.q�!����l���/��^��ԁM
t���	��&lv�-�NЖ\Z�b�������&-�G��%nG�j�z$��x��T�L�?U�9�É��N̓N_����.�G�WL ��5����]��;��r�&I� ��D_��8��՚�\�5CnE�x�tv���N	p�3�� O�vC�$�z����q��m$����$�z����p�Βr��
TF�ob�����;q �|Nk�@$5Ms{���M�(3 Ո.zf��5���{�)^T�f^<zQp���/^Y� �k5�xhN���wܹd�]����Emт�[�h�F�ߍ�K�gwH8giP������g9�<�ܩ���w:.D��Z�	:�������a���|�n?_\�����I�u��!O�v����U�/V�̶˄l���z����r٣�,c�}��W[��� A ��|r�(cA�]��>'ݏ�E���Ȃ9���`("�d����qU��Lu��lQ�����s�)���ʻ�Ȫx����b�KI+���t�d��	�NC�E
�x㹣�<H$�F@�!W\�)�Xk,�N	p�ș��ʂU�#p!vIk���k'� �wvܻ�\�5�#�fJ~����U�Nř�f�d�2a� �f\I:�ܝ��힍��\�O�㕍��ޭ�,��8�n��}�l�}֜��M��dkV1�iʂ*p}�k�ؾ�����;�k�_|֓��k��?/r�/�,�~������;�l`>�Kv\]�H�0�P[��8�y��G��[N�ypBޤh��l١���ͥx�F�p/�9J9M�Xm��t����{$�����Q����s���tw����R��pL��f��{ E�q�fyC��69_XNq�m���CI�f��
�选��0�pl��q�8Ӓ��$elv��x�����c�ae���:j�n����2�8Y����eN�j�������Q-t��nj��^v�LȠj��]�� �]�P� �\Ǡ�d�t$��ձ'{M�mDg`��qd�UV4�K'%jN�8gv0k�WNfL���L�՘�e��"$%]sAwul���^�gu�#-t��.{�fmE\ ��L����rI���E�b��	����/�U\��H�zٟ)��-$��ñ.�d��x	fvuWI��9w��$�z�����,�j׋�7��n�-���'b;̃u]�|I�>;o�^#3pV��r�� �*��dI�~�x���������?tֱ=�����z!hDn4�e:��WVV����K2�i^fc-����|�f�'`�� �x���I�+"A$�/_�x����-��Z	5��E�6ǋ��$���R_nb���ڲ�����dPd�rܓ�"L�ug��s��>j5ڷ>�g��[׈��ݴ��+�-9��ϐ���r�����>h` ge�̒H7�� �W�ϙ�|�ɢ:q�I�
�v`����Ft�Ȑ��9�� ��T첄dDu[�Q$��z�����yK�8h�`�r�z�|k�5}u1�(����#�-\��(�T�Oѳ>$c��ZIw�b]��9Q� �˥f(k��[f��@�y��A�$�:N�W(���s�%���ʒL�%H3���9���"./�͡�u�n��j�g7'6[�V%ׁQ&����'b;�zg;�I'�:2 �	�r�R�c�4(�]� ��F�y�l3Svt�v���S0�E>��d�|��i>���$l�r�Aw��r����}�v����̐v.С싃�G���P	>�OUpܓ�r��%����Λ��ɵ��n�ڤ ;��[$�W[/7n�$���%';&6��5 ���͛�9�On���>'��v���~B��ҝ�'��fF��ɞY��;b7(���� �� �F�mM3U�H�[U�Aj�� ku33^!�4όJ݆�WmD�������^D@7+m$f�T��繷A��RΔ���3�ι#�v��uX$����YhJu�ŊV�K�.�:1������"�{��LA��l� |H�쩟������J�r���l0L���ɐv.�8w�U=q� ���gq���&�� ��S�� ���X×D݂���qm������n��ř×�ݠUҶ��$�^\H� �����x��=	�<F�M8���ۙ�!fɶ#Y݂Iا��NSq�slVկ~Kƌ]ÒI��3�A �G8��Ƒ�;g��˪�ex˝���c���V~ǩ��+�o�3z��C�rUI�݅����i\7�K�[�]^��p�,Q��1-y��# %�:V�f`��!�������.㞯MS���Te^ӾG�<H��� �ssng�ۑ���˕������?ch.�֙%"&,�p�	
|v�^���B�J���l,n�����K��4�M�=}rE��ĐI쎈=��A�k'��d�q��ݻs$�P�%��3�E���9�#,.J�,�{���[�w�<��nӎ���w|�)�k[2f	�;���݌$��I;W	�!�b���1���I팏A��	��3��;�v��d�,��V���{#^>�4�d�"����K׀��'.M����yP��d��A�S���z�-�pX�陒@"�:#ǩ����zF\����̀|w?J�3����~�>��گ���O`���0��L!ͻ������2`����ʊU4�1)�K�b���,���n������|o.��8&^���H�=lq;�r�px�Du�[WoV��إ�ݛ7.��0sɺ띘���6��nx���ɔZ�ij.��@A`MHG�%�z���k��`n�fͶ6�p	�L��=��^ގOH�v��%��u�cn0��Ǳ�UlU7U�����5g�lj����f�+6�T�v��+^��`$C�X.^���8v���S����[�.�ݡ���:A9��K�f/�tC��6�d�I��x$:���B��XrnI�̞��O��s�S�dyx�;��T�����}P��Rz
�����O�'ױ� ��-��7PQmq���6$,�j	×L����3����K]zCA{�
�j�㪕Sv�$�����~0e�s[f�8r���w`݂�
0���H>����˞KV:��s7��	����\��v� �cL"	=}��{��Y�������]	�z_���r7�]ٵH��P�[r\3K�dS�vLY���r���"�t�M��-6q�k��],��1���!~)3�t}p��Z�PH��r�R�
�u4���u8�ԧT M�B��&/��c<�5	>�|U6ɡ�a�=�M��xx�t�˳Jçd�v�<�w���n��_~���g�n��~����9m7����yY�O�>�{������`�f(�$��˙3�x�M47iDu����]Q���:Ap�Ue]�^���}�� ���B�.���6`$�8��	{��I��K1�]�t�8�3�M{���>,���I��Xx��v�-FfO]>���P	�;�h�ɜ&r�<ϟ�vg���ٓ F5�)��ٳ�w����LMwmĀI>=�1u;zDH��b8n���\�ǌ�)�ʄۄ��=��r��uÎ�\�� ���ɝ�.Y�'�����㷹p$�O�:bܽ�y<&���T�`z�n$ޣ�ngfيv�|�A����N�3��Mf�ȒN�K�&�3e�3�����pQ�,v1��Qf#�=��=s:t���;���ǧ���?������-�IMN�3Fc4>6:�iɶ�ƈ���Nݴ���;}�9,���s�4gG�8��eB4����r}�^��Fzw,𛲎�w���7}�&����1�{�$2�s]{�9�曖�k:��������I%�
�����{�o6����̈́�*m�A[��}���D��m�_hЄ;�o$�������0O|�S
��B.�|����i�X�wI�������������rg+�wc��qI�&�%�}n<���E|\�V��7��q{{�칳ޛ'9�"��%da
�;"��z�q�a�^�My�>^��7.
o����=���ug���xm>��M�3�����n�sӷ��D�Ȼ������K���`�FFLX��B��
�u�����]�y��%]4R�3Ӑ�=��A�h������I��o�5]�T��M/y�u��5i�w����.�ph���s���y�:�������s�O�za�:�ח+GR�^=���M�k{���l�{˸��(����a��0��S�H\F3����J;����<z���z�G�߱>S=�;�<�{n!��4���#�=��n��� �4�����q����7꽭g�Qx{�� ���Q�-_|��|vL����w}sh:{��t�ۻ�	"����v2�Ξ7|t��z��#����p�.sy�д�XO�"9��铇f�#ޖAI��r
��ˋ^-k�$\f�0���O�y?��I�$:-������v���ox�K=9)�f��i\uy��������q白�w��e��me�q�u��w'yGv�\/n�����4��7��#�q��l���ӛ^ڒ�+�{^]�{ԗgY��;. ��γ�2�:9��Al�sn���qљq��^�Ώՙ۔�\�^غ;m�֭���w��gQrVol���i�м���I:{ޢ�m�gvq���/{'�^V�=�ft�2��{�.��鲼��;�;"^Z�����EޓZ=��Ӑ��Fe��[�:��u��oj
ҋ�l��;f��ו����[Ey���: ���M��8�������5y�z[o";����[����E�g{h�-�]��H���/..�\<ޢ�'���}A �tD|R�K�C�!�[���W���̴����0�A [���If%�_����`�]=��K�UL��\L�rv3 �m�H=��m��^����9��}��$㗲�<v��Ǌf���9s��zK<h�ۅI��〳����}�����/I<�����1]���S&p�܄��9��$��9�|H;R�`���![�U}�00���lv��:x�сZ
�Okhd(ņz��D`$o�^>$u4��v�.���'nT���͓~lgvv�s�X�L➆$�m{z������=���z�b<F�O(&:���ܔC��)���vl�U�\NN��$�wD�S�$��˟z��~�5����4NY��������ǘ�{�I�=>��x���pJ.r['�d��Pq�؈Q ���*Y�R���6j^w�>7O� ��̆`�����L��`1W^�I�<�+7K*����e�8�}�ӈA gv\�x���}��|���|��fl�2�����:zp���8���k��A6�9ř�����~O�*��C������qN@bA��ẽI`c�� 7���N �:�)�kZ)g��O2�n̂|(yOl�gq��y&z{7"`�H�4���q&�$]w����I�gF2o��)i���)�OJȀğ�ˁ �]hp�Ⱥ�OY@�Q��D�v\ω͓~lgvrYyu'�3�;��C���{~�J�j�$�77nD�A���7Rt)��O���ǉ�FG;��p�E8��ڹ^3�MgD��B�y����0V�H��`H����|H;�/�5�uF[7��ڄ�8��c��,�'�cU��;2´c檳`���ƍ�R'ulK[clcJD��/�͔+�_�B��=ܥ�v���e���ԯ��r�<$�uIX�᭹��6_C`Y��OM��%GĘ���F��Rv9���̓�:��k&l�P����C�D�Uǆ��+3�b#R�u%��#Gcr���vN�]p0�Ʀ94w!�k��Y��rg�	!V5�I{@��J�<�e��g]�=XD�����Ì;ѓ��P�e!6�p�G���ͤ���VXVj�f�x�J��Y�[&�kcz�5M������lP��5y��T�f�?}�A��C�����tI ���I$�H��9��=m�ߛ�\e���~0H'�ۗ2#ʆ�35;$�L�f|g:��wacn���s �+��dH=�1���+�C���Rb���<
�}3 �OfK��W۞�}�d}u�s$����[m�5�fb]2p�d�hg�Z0���O]��L��ĂA��1 �=/�֊)���}��3 �I�733�)&xu'b2H9R�g�޶sޞQIM���#nfO�:`G����O����iF�w���ݮ>}��i״�Fq8.2�,rz�)�{�[s2��
l�j�X�����3LK�K>��&�_�n��'���*��j����!�&d��S���4,��(�rZ�����<�Yg�:ZR\��jb��Iû�f��pe+4�3����Mg%>[��O{=�5^�GL���?3�f�ȗ�����"I�$�wt�x���I��	m��d�&��r��̚�����̙θ�E������I��Iy�F�t�H��f="zz= m\���2g���d�K\l��h��%�8�$��[�n@$�_8���L�}��w�T H,�Qkv�.��gb�̘܇�M��v�Pr�'u�6�g<A��q$�ٓ ����	�I#��A�wd��9y��ve6!�3�Wh��	����vUd��2��gCd�छ��7�؂>3ӯ �;{.$��].�6��<ɶ|q .��"�mN�,S�I�<*�ד ��^oa��j�˯A���	$f�\�o.ՠʄIz�S�MA�g�l���i�c+^	$���M���Hn�Zs��^=�ѯP9�w��s>���n�-[�|htQ��iB5�UJi��if�Y�.�Rw�3XP&�4�--B�︐H웁 ���q$�P�L�[$�1vtfA���zx�Z�kĞwǂI�#6��|H$�t�V�ا��t J��u�c[��p��O1��>$��������=|wI91�$e�\ω���j�l�1����{��8Fm�W��Z�s�Yw4*r���A7�;�g�����������ǉ��^\O�$�{f wv̠�q��$�ٛs ��f�I��.�b4����E��=�e�Y�̨�I#�{f xlE=)�F����F?'�g@�vI �G٫��&�a��lw���S�'ǻ:�IntǠ��2A�;�;��>1��WDW	Uױ �I�1�R�}늼���]�:����c�g���QH��0yod��n1��r�}�Ǌ�ql~�n5H���;�]��,@-�.y��a����3z��Tv̒�t&`�̓.Ό�sm�{%�٧:�@���s$�{vW�<v���(.t��|����.���#���B�6kU��a�<��r%]�]KgG�ɓ�K3U���	1p������28�fLz$�Kq��Ot�aTsSl�]s�>'���t����H���9v��N4G� �P����1u��1@O��1ĂGT�!���9f��hz��q&w��D���pA>3��`�H��bN*�Q�o��{'���P�c��R�grgd�	��GU�;O73���|���o�@'۽�:��\t+1�^�a��A"��$!�Y�r�4
�Z�����}��>(5dU@n� �k��|O����+�M�
ɗA\��l.�2bg�T�g%�����S�h�Θ��};����-�7�~K�BD��2=��y�۩�ˮn{lc��U׹��<�g�_�<��*��B���a�%��&t��L1���j��ץbNm<�2�M�U���H�E��t�G+a-l�&�ivКXM�k.�9Wnϕt�[�!�]]<�۷;�9荮�ۚ��1⭋��a���z9+B���t&�����h�iM!�%Ѻj���֐�B¯N髞�p;�Ȇz;Vw1 Ob�����`��<�mg=��׶p;T��:�4�=�Y���8�؞{v����YA��Pt.%?t��|�T~���ю3�o�����I ��ӓ'l�`��'� ��DH���)��;��p��O��͙ ��y=ӝ��JUe�L �)����9E����;5��n�h���v��Gs`"T1�z~���J�Z����P��� �FoNL��f�)��0���s=���ӛ�f�@*��y��gbAb����f�3k)�yV��J	��ÔY�$�q2��g��dV��w��/j2�s]7LoHR݊  ���$�l@�<�$۩��ǫ�~���_�bi��L�G�Q�B��R��Ĭ�j�"#��h�͍�nj�o�^���O���h?�u�[��$��\�	$�]�"x�aʯV5ڀH=�=��8C35�&b��щ3�o ���(���=f���N�[�\Jb]�����rx�MB��<�p��<9jߘ�Y���[����Q%�اt4���6�͵3��-�0�:��� H���	��؁ ���ۈ���޵���;��JgE���<
�*�ِO��"=w�Qws��'��[���q�$�w� z1��$�N�:r^$���kmU�ȒA �Έ��n��jY�-�eG=^L�CoQ�#K��jP����i�\ ͘{�q�C'z{�yݐ}*���܈����Z�VGlŽ��~V�\n���9�{(����}鮱`�]f��픙f��{�~����JCO�7�^�~�A5�� �|H�n��Paz�7��G\UL�H��؈9,Ik�w`䦐�19OQ��'vS+�ؼ}�>'Ď͈�g��5��k�<V��;ّ�Hk!�jwNŋ��3�9�I<�2O��qW5��EW��E`|ƺ�����U�m,��0+=�M�&Pg1Nj���HOq��^\/0g!:����Gzr��ܚ8����aN�j�� ǒ';f F��5�ӄv'���ټ̦
�eӴM�OM�ǉ'���`�]�т.7��,��L?lEk��(;9O�pļ	�w1�$�=yQ ���e4Hy=Q �z~>��ʙ/9�Y�(���|8X4;��j�^�:�suONP,[h3\&,�WQfxМ���S������CC@QǞ9��K�l"7��LO�l�\�5/��	<��`�=�)�:vp�PN UxwU��'C��X�a޽��|l0I�.�z�'��?4�.��9ձ}Y�#ce����9)�LO7N_La ed�%�ɮ@'Ɵ���޸�J�&�.�QvtfA��,H[�,b��eDF�aN��L�I=�{Ÿ�q���;�Cf_�:�1����;��'��Ϸ�
��ϚE�t�e�K���3Z]#�������痷d�����HUYd�O�5�ǉ�ӻ"��w'������	��ˈ�i�3�$lV��s�I�.�z�� ����R��+��%�r]�0w.�����tn��ʼQGnk��ؖZF�ZP1���}����I�:p�3��2�  O]�D�A �om�_�y���\.��x��ʉ���L����҆Qȑ��s[)����um؈$��TH$ݵ�N�կoO0�{7d��z���;;8f('^؞��(��Sv�9X�
�d��ܼ��|�� d\�>\];�%<ɉ��l��Nh����D��|r��	�^���j޸==��&{�1�p�I�3�(�8�Ti��A#�� %Kp�H���{�����޷x5�[�����w��>��1��� Q{�����@�
����������&��8�����ʋ"����,��� ��0���
���
`劈!�� ��9`�`�9� `C ��p;�n0�� C� �0� C !��0ȈC��(�2 ��Ȯ `ȀC(���+�ʋ������*,2*� �0�ȈC����20*�m ��������ʋ��*,2��*,2"�
,0��*,0��*,0"�ʋ��ʋ����0�̨�,0
��0��*,0"�
,0
�
,0������ʋ��ʋ�l¡� �2��(,2��q��:�9�?h�
!B�����3O��?z��0�������f��?���q������v�?2f}���y�˟�|_�*
+�����?J��+�{`TV ?�����>@���I���I�7�C������p���wCd�����~w��������>�
ϭ�PU ��$D�@�	�@��@�A	eE��VBXe�TZTX%�a��Qd%E��P�Q�V�@��Qh�I#������w������(��4 ߨ�����~����������}��w�3���*
+�~8��Q��;67�O��a������)����}@�(���~�}�� "��J((���!����}_�vnl�

���v�H(��@b}?b`=ׁ�?q����r��-�76�^�9���PQZ>G�}��/����}��(��O��]��Ϟ��po߁����$���:EAEy{?#��@�(���ϻ�8
O����hI�0?A��g���N�	:��
������}?Hn���?���>_�|/Ԫ�
��y`��eUW��V��>��>����
�2��f�jB� ���9�>� �`    >�                            �  � �(d�M(� )��� 44Ҕ��V���4�AE
h�
 REUQJ(�4H(   �|                       @               @       �L IʀY���9Uѧ �  H4 u�94*# �� p �Qf��  S�  ���z�@ � 	 2 �T�]i\�IE(N� hR�"�1٥P�T�3J�ТI�73TUR����U�  �       R�J��:�
�s�j�6�U�*�T�P��� �*B�����Rr�T�i"�hP��j�J�T�� ���P��JC�8K` Q/   ���b   Hz ���t.` ���C!C&�0�@� ��Z U�   �        `,�� �@d� e� qT�j�Zڷ0���˙��� ܪ(�δ����PZ 	<   q��=b�-�Mik�q"��;+F��
�J��m���p 3J�Y�����b�ڥ�ӥ-2��kA��@  �        =�Re��cF�]֦���ꔹk�'Z� ����m�8���U8�u�3���� ]C�W6���\�U�f f  �O�W0�c�m�8 �m5���f���w+kNwq�6Z��*I� :�]�fu�յͻi��9�v�-ʶVjPQB�x  x         ��xrӌh[���W6���9��(� b���؝����QP�`�p�0u�� w]���;�(顢Jh2�  �K�hlsn�����R�k�봢��W6���22 uӀ4(dn�Jr ���ه �Sɠ)*B4��E?	��)P  ���a4��M0=��F�RP# #T��i2�J�40�I1JH�������٘bg��07���}���0���:O�>�IO`N��$ I6 �	!I��IO�H@� B!!������o�8��Y��������n��;�+�n����ow����281P?v;&^k^B�X�����s�V���6>�(ۚ4�,�܇V]��ۏ��98\�&���q��1$�Ǥ�6����䜤���'Z7P�n��sP]ͮ�p`%��؀&���ػ7�T�^��53�߮s4��L!t�4]�`�-���;R*M��z�"㏧�0c�G.�r�:��X�Y�@3nC�f�i�;D;���h�c5B#�����&Ezt�Y��k+5d�o�r����B�{�czs���W�d|w�SpG�T
*wd��G{'8�>�����8/zD��}��9�ҋ�ַٯ9�rõn-ӭ/�����7���ٹq��
������D=ٯ�C��ef�8@ȎV��86v����w4��r9cٝ��&<���˷��_w�}w'U���;����H9F�X��nL��*�'٦-�Y�y�\ЦH�2�v^!�x�V��O�6���7n^���@�>z�⠫�!l˛@Sx���e���߻8X����X�1�sw �*DR�gHx�I=s�4vZRDgkqs|C��ә���>��R�$چ���[�pc��6�h\���1讵�@�Ǩns�8�[��c�6kYj�P(B��t�Qv�/B��)�p��3\�z�8�+h���z��GNN$��!�5P{�0n���8̱&�����ڻ�cX���;
]����	k�ίd��5���uDM�`8S�ޛuj|�X9�B�]4��-=ݺn�f=�#x]ɝ�*SaWgˎ�|sQKr7����N3����q;�0B{���<�k�,vu7U�D��枕9:����㛼�ݘޚrS���h�÷�7D8{�F%�n����J��S�Şő�<Yk
/
9��r<�=bOC�{Z����܇u�0�,(�L�Y�eE.$�#��{s�3��f�����݉���5��b���v����ݱ5��M�4u˷����q��o{���rs4���J#PSh8v<���Xћ���.>l�9Lo�K&��dQ�	̬]�Fm�"(⛝��St��:�J*��R���:��W�RzЯqwY���Ё��ʊ�ƍ�n������F��Eƌ�¾V%E�&�o�L���F�a���u�y �4�,aa0}�w��c��۲Tyj��y.�ν��ܺ��\5r��x�%{�����ׅ��af�����TFE�eY�����ט��b�O�7��.��0��.W\�֍ΚCQ�nӝ��kTa�=���+[�D�E�gf�X
�2ȩ
�4��d꾄H���9��CL<�5��������n�0X[�vֵv������u��O��.
��n^���y�4:w^��A�m���4�ϔ�IfĄ��Y٠�FL�p'Dg;tf�ۚ���>#���q=�h�F��8p=�O�3]�ٴ%U�%5�nQky�Z�9�N�2m7j���N�M�M��[ݔ��cxwƦ�;u�n�p8�w�]����u�0�#�"�t�Nusp�5�ۺ�я_2q�;��b8[ȰvK�nR��)B���X+f;ݴ\��6ӽDN�;��FI���82䀋�u�%#sV*��c����ӂ;ځ�i�vrӜ;-�0YȞ�o;I�w�}��Lܛ4��-9�h���Q9��
�����2Ó��jxT]v[�����]X�s�@M���[0g'�jgr��b{s��5�(1�ڀ�j�N��6Ķ(�}1Y�g-�2�k���b2����7���hT����r�����sR�(��\��^�:\��c\L�FtեՑm��[W��pŀ���4C3Z#���i���L
�	zkvS#��w�\닦��4k���T������On�@oFn����扣d|�)z>��l�;��DN�Nhܛ��S���H>{q��F�ou�?.��f�����W(�,�DS��c���h���ϭ�J��T��:-C'�񧱱'Q9����li7
�fum���p��󷰃�}&W=�ax��ur8���0��w4��X^�FL�컅]�&��vf�U8�Ui�CcN�]�0�$��u�q���y;6kta]4&EÝ'�g#pCۖ���:C�����-�����Ⱦd�k͵����ÏMH�q�{����Ӭn��Ed�^�t��<yGn�}n��y����MiˑP�bɈ���}_&�ΏNuy1�ȷ3����vT�7��ea�swav�q�1��-ˀ@������D��V�Jd��n�޴c=!f䚚��~J�x�vb|�'G^�2:��T8Ó&nU�f�#VI�ӲQ�z�2��B��\�e�]�h��z��)=:�L�8�Pn��t*0��w�1L%���doZUσS�a�*J�E��f�w�ʛ��a�����+�ò�u�N�́2q7X�L4t�1#t�(G�b]�!͙�U�t=�=�4j�#�{{y�tt܊ l�Ε�޻o5{yv��3��27Y7��!�P�����o� #5nǋ9���Ӡɒ�z�3�X�̚�v��Gզ��P/R�v��4'�ݽ7�3I�O��ɩ��-����t�a��D;.�c�y �ūJ�D�5�ِ�s��@��wgY�;���uUdH�<��8�����4�Np���m~���b7�L�hq�5��t4*�P�N��`�]�ن$RboqK3P�����_Ps�wV�W^�ѡ��,�Ѯ�ŵ�u���ڲc�1ڸ
E=�%��j���2p�2�
��W��nN���3;�	���)��`B���]�c�*t�B�d]��D�I���f��=�V���K�Xr6y�(#8�#�,VN�=�M�z�'��z�Kk����#�bv�2og9��=D5zQn���m�<�}8a�*� `x]r:�H��n��p�q{�� ��.m΁�	خ�0oE2Nm��`Ѱ.<g}f.|���r\9�n�N�sH��<�1�ƞkOg=�;� Z٭�������M�I�d�b�*�wt��V��S������(kw����q9;h�O)�F����0rh*�r"�]���*�3�hgNţX��9c�~�P�`Ti6�ѧaܛ5>mëB��x4�q]�n@d����@��:�n��{�B�T���;F��A �
�����+)eҸ���N6�%��ի�L��LX�[C��;�������Y&Xu��'b���¢9\"gN�7;/>�go�Vޝ�Η7p���& kr����\J<u>.�k�3e�� ������j��6; �R��q��7㳾:7���\'*�IY�0�Z7��?n���ʳ��}5D6Jђr��G+0#»�v롤���i��aD������p���ضd9`��C9�v�@<�0�1�����lڕ���En;um��|��sד��M"K��V=](��jQݴov����ܑ�t��:�����K�׆ŋwZꘞ�������d�VP�ŻF8Ʃ����\�����8r6顢�S��G=�7Or�i����\+ 6b�����(휟4X7��_�[՛������g,���KI����m����J��w[�tr�ܶ��'<4ސn��:�v<G�8�������V>v�׆�Bl��3�G,ս�&_��V<������rm�z4k$��e�+�l��|3�� 8�Ʀ���ʽ=9g
����N8^��UG0�y�NAftx����;�`Հiͧ�9@�r��Ŗv��]4ם��-�z�^8^�z�䯛	ˏ��N7�Ӌ
��]����jc��^$C��i[Ö�/��2���"˶3i�w�]��n�rD�;�i��u<dl/�k�a�u_1�ـ�9�� ����|Cޚ:ay!;�F���Rx��C��K�S-ǋ�:u1��
�mن�z��S����fr�L�{9���ã���o�)b��k��}����r��y;��e8�vG��dl�d�{�8�8r�0k�7����U�kۄP*����+A	��'d�+9zl�@jz;�l��y�y����2.[��ʞ�Xg��i��t#��;��3s��ƞ5�d��ў�b�������-T|�����+��\����x�u]�p�<��aST�\�i���kj�Vk�8%<�<O*#l���"tʠ��G^�d�1˺3g=�S�`o�����5u���.��E���t���D��3��NZ��I���]��n跃�&��M�@�'F���*n�m�Ը�P9�F�1vmܚ1��3���A��4�C# �	�XyJ\Z;IOf(ix9>��%b��M<q��VUFE`�qD��`[c�Y���4��,h��,:)���7�s��s�蜖�Y�\�ѧ�ީ�[�=���fn�Q��`��w�=s{6����ۃ:-ɝV�{� �$��N����P�u���Xy�x\�nv�xNn�]��R�w'����rHَ.�����76p�it��DȔBI�Ɩo\Zq-��7P��GH�4��	��´�(�Y��36�)��P�I��;n1�+�iG�y�^�4��|��ʺ<���ɛ�`�e�Ǧ$�f�3�*q̮!�����d������n�ÂaJ�T�������8�Г�|����sA����~��Mu�HR{�Ѭ>y�"��eAj�ގsa��,����/h��j�%���<�^*����q�2Ei�	�&����n�m0djc�|�u�;)G��"�����v��Q͜z�c.����4�D������SBs�{9����(!��g`�ڳ���S��z�� ���fn���Ǡ��XU#[�ݭr��{�Q��)ε�Az��>�q�%�I).7x�-�����Z�6��9�$=����ߡ��"mv>�9�s�������H�%�*0h+{R7.�"Mq$n�7y+2�����[A�i�ǻ�k��#�-�E]0s5NX�7��3���	]v%Y*j��峁Xwo*��pL�Vu�N���P�Mm	���X�U杉"ɢSx}�p�<�u:��mWpd:�`U��[Fg<�3�E@�"�t]F����f	�"9:m��N������.�]���k���Yˈw������L���HԔ�sz���;��m��6�����&�����}����e�gd�Vsif�;4NJ��v"���f͘^���N����� ��q�kưc-W �G��įL����������i|�շqr�V�ܶ]��qv戦���7���-�nX�b�O1�6�;����wA��,�>�'7.s��1*8���f��`�HFo}��1��v��:�)�DB�~��V	��:�Z�).���p�݃��4�G6�ƨ�&R�M��$n"6X��&�ґ�P��t�w��w]��ɻۏ{p��z���\�/��z�+٬�z�}���]���Ǻ�۽=� 9�?jIu~�F�h�͎v�Ii�Y؏��l���s��䈬-��ٮ�:Sܹv��d�J�Fe{ܳ�;Un�8��\c�]�"%=B����ݠ��޲��a5Dy��f�]���﮲���u^I����zV�#fj}����>ܸ��sN�ۍ��n����h��Uż֡�>�oe�à�g`@׏R ]CDx�Y���ݹb'����p��e-��r�����v641M{�l*�
��&	��n��	��Q$N<�So�q��i`��z\d�9�/\�2��h��u�۝����1_��'�x��#@��Ǽ�t�Fp��	"�nuǽ[�/l3����4h�R���r�'*������<��A�Gt����,/sowmfܟ,�8�\�:1���[˰m�(���´6�x1��;�Pd�)���o��=۽��HD�`8VwK����[�	}�ph�mX�[�0�!K7��D\\޷B��a��%�w���L���֫�=nvq2=r6�/�3[��Z�y�'4e����\ۆ������o�n{��i�U�*&�n�Љ�Ê&d&�Dcźx�X7�n>а�o.�S�Vr\�Mguc�b���w_I�B{.՚x�G2����iJ2;iCxV{T���Û�=㐞ʄ����yĶ�n����n9Ӱk���ݜX3�z��ހJ�꛽��xw(ٗ�9��|ZkF�$gL���/x���G�O}�J�wsȣ‎k�Փ�k�؜9�qU���ok�P4cA�Ɲx���H��C ��J�f�]V���`NkA'3p\@o]�w����R�;D]��yI�k��I�jݹ�U�F��1:�םH����J˱�ǹ�4/PS�o#x�k�.�0������;�\���97!�yY�*kfҲ̽x%���.�w��}E٢WZ�KC8��`m�ol��$)v��w>om���a�o+[�SY$��ϐ���f�C�.k�Ħ�ŉ�&Jo�C��R�Ol��*6E5�~\Vp��S���.��y�y���scb����Թ��
��{O�A�c���3�by�mdɻ��xs�h�ƺA���5�Ӟ���n�&�6����3O�A�l��Ft�^� | �� ���.�q���E�(Ln� Z�Fd���{��[�O�\�_������Y!	'��J��@�H
B,	!� �!d�X��$ ��	IE� X��RH@�@�HV@ AI �@�"�RBE!$H�@�!HBd�
HAaX*��
I�J�E�$�$�*V@�I���� �@�H�H@��@"� �*@��!P��AdVI
��V�aE� T!d$"�H(@BJ�	RE� ���B) H�HB���$�YT@Y	"�	%I$�RI*@!! �@�!R 
@YI**I	��XP�*@I ��@$$?� I��@�������������C�Gqyz<����H��w���v-�y�f.���S���ea��(u�G��}��s���:<��]�Ÿ�b3�^�qu�Dނ��iT�q9���Y����La�/�<��_q�÷�CP\̛���7j��Fl��oT�=�f�;�^<��^j's�3�| ���?\�Of�&��&���	Ù�mk���F�S�|�1��L?�{�<���X�.��xL`n��Mw�LW�:#�NH���!��p��[���)-m�P,��o>M�ǎ�[�yy
bE�7�4܋�>:�Ũ�T���/��\Nx������8����=��������w�K�vv䙵�`�4G�勱�l1��결��@z2�Xڍ�5��xg��/*��a���;��rުj���̽�$M�nم��u���Y��*W�k�6^H�x�'e�ų7T��^��f�����2�em�D��̊�6nӌH�H�&�.����1�r��3Ɏݤ}���u﮽����{��(v9|O(Y��f��;[&Ѓem��m)�j�D�VŖn�dY5"�x��Xy;`a��	��qo��ז�D��M��+�78��7�,��@U�eLV��t�F�ƆjUx�嗂�L�{5�D c:��Sz�Rs�Ӏ'��7=H��/�da:J��Ҕ�k���;^���N�� ttP�����sf��/o���]��~��}�AcM��<n:�'ڼ�}���xMu��^g�Lrn�מ��bK
��P�M;T�Ԝ�d�it	�gJ*{����Ju;�=�=�?k��4kl�^����뷄ղYR`�=����	�{���v{��aȻ����I�D=��o�Û��+<��,��h>^�
7ox�"al�U�*n�g��L����Ú�|��|3��F���]�a��uo��'�W��&�>�K;xiH��5��挹���		�0[V0�(㵞��<t����Ϣ�˽��+���*���2��,�ĶC�L��Gm�޾���WO{U�O��j������$��M���'u�r��k�T���j�&_w<��V!�'dUe���UŜ����� �ٻ�����܀C�ՙ��Q��5�l��:nh��o����2t��7��7:��h�V�i1kbzB�J�F���t���g�>FS�B�����g����[����;�������|ﺮ<�v*9��V՝q2|iEP>�q�s�e�F��s������ B�n��_�ڽ�b�g���t�Oc��pjۇtZ�����f�%����ܻ��/.S���5�~��r��;�4Nv�󇑷��zxo8R�l��Z�웣��������6n����ժ��vYt{L�[���571�w�B��h��6$B��``E�ݾ���C������/��AG�䟎�Ń��f���v�z�9=HNwio<7ި}IU>�Ｒ�1̓h��\?Y�\eC�6�7Ir;�ֻ�y��O�_/u�<�q�?"-���Ƚ�F#�h���P�O.|�~k����)�1�ͧt��z�����}t�
��g�A�c8�tg� c�~w$ݯ=���r�S�=usY�\��M2�<0el��{K�������%n�Űv�n�՝zfN-9|w��g�W�o;jGa�L�w�[�sTk����p��О��_m��<&H稂�|G`�ssی�S�ޕ���X�������5?���P#�����à%���A�y��#���4�ԯ?-�[�ݺ����!��6�`[����Ӻ��.�����s����^�uz`��<�X>x6F�-y0����[8�;F.�fG6k�T<:$<�m�9�uOMO��=�	��z�{C��_4ɒ|w�^���ūش\�繦���.�8�CVE�����V-�z��w��y�<��JL"��{�|ȧ�Þ�kM���1�$��{E=�W>������������=Y:��Ȃ��==����=.��o���W�s��xl�邠\�J�l=��^���OW�\�>9�����ٹ��G{Y�y#�I=&�Ww�Y���O���O6�bm�̻'#js�o	X��u�����˼e�k����2���&��ʃ���{|8z�Nm�҅{-iJ(3Gp)�z�k��o_<�3V��_a�\=j2*2�؅�;iޓ66Ѻ������*<����[�	=t��{us�5�^�k���Z�ܘ�%�X<q��E,] ���w2�f�������/6U�̂���u�?TsL�y�����%�&DM��Y]tI���6k�����Ќۣ�.�^�nt-V�c�f �o�'�=�=@����E!]Z5.����y�ױ�Ȳx���Y���+)޳���.�VNܓ�$��̇sC4��V	i>���g�z�;�ʐ��������p�����n����@D�UG��V�٬�T��[���h�nAG!#:�9)-�����W�s��#���z�#��?u��ŭ�_��N�aFC��pEE�m���ͽf��3i�|�/ts����O�xu�U���A��u�x�8�~�|w��z�>{~��ʷ������/4�>�n���v��V����'N/gt��o��|��-ݏf�� O܍Ɍ��=�ٻ���Su��V?=;9�5���E��9��o�]ɚu����3}������s�z;ⷦ���(���qRc��8�JM�(�ҭ��������zN���@ѭn�˛�
2��J����T(Ў��t�0p��Oo�;?ob0��{����mc��[�!G��!bm�h��r�x.��/ MY�w-���fAj�+�w���k���U�V���{��u�'���ܡ{&���^oM]���, {�lɞ�7��un?g}|ѥ�b	��4'��M��gq����wn*�F�{9�el�}��=����U�*Q�n���+��ztbw���!)�%���zk�#�0���lJQ짰������x�����b�W8�
9�ٻ|&⫎�:Nچ�mOh��X�#�NO��.�7�:�{�q��/������"u���\��7'������x�Z{���Nf����f�$��x�3ց:]�Ր�d	�ȳ�*��ScLA�b�m��k�߹��G�����8��f�}L�k�xc�vn{�Q�P����{|�KN�$;��ԯ��٣�Op����b	�����	�`��۹I��ƺ���\yX��~ׁ�z�����;i�����VQR������g�pՁ�\�t:6��P���hv�'��$�5���𝞆xrn�W��������M��wN-��S�B{='B�������7����+�������CX��X]sB&V�79E��7����z� � ���%����.z������e�� o�zo|}�~^y:Vp��ⷵ�$��b�s���s����L����az���,C��׎��^���v��0�����\z�Ѭ睲;Nz�|�|���R�����(���5��]'��5^�㌦��վc��n��j�Jǧw"�m��[��ͨv��畝�g= ���������!��,��w���?�UϤcU�x�){�N�Uu�����p�#�&q�ww�wW�hU���+m<��bwc!Ǟ�W8�R��_�9�TtZ� �Ʈ�%�c��&y�qr�T���wYWѫ�j/+GB�m���R���m�>��*w�����du�d��Z*��^�O�i�LA[����#�}r`�����I��c��=x�ɤW ӂ!��r<pg��]�쭨hX�F�����W���7S�ˇ{#�L��#�eء�E8.@1��f���������QZ�}-׈槕ᎋ�j�����]��svof��}���q����$[os ݔm��JoV�S��і�@@��ɭ��F��%q\P3��<�=���e��7�c�<����p�M�{�� C��j�x�X��x�����"�򘯾^S�e���%�! �EA�W!��)��/nNW��V���u8=�����:�@I�ww|+�k���{'��R{�f��&�#˰�b���g���H��m�^W���4���ߏ]��z<�7��龅{�_;,����#��\W.�s�x�n{G��x���"�幩����qS3&���ph�s`�D�'Fj^��P^����r�m3ͫǻ/��j��y��(8x�Y˟zK��7=ǯ�4����)���]�Ř4���Cu��I�;����H{{��%�v��lǞ�N#�P��1>�(t���n��}���I&���5��=1�R�r�?H��`�~V��|��|]�G��eJ��c���d@ñ�|��^i��4nL��)�{6<��%�f� ��˽�[ �=��N\*�����M��פj��w&��~,��}`�2nY�R��c���_,��x��z�ݧ�|���6�^����Ǚb�Y��/D��)��&/^�i����ؼR��FY#E����C�c�n��se<#�G}�y�^���Ժ�$}��|��y���`��Q��F*�f�U,�������`N�88O�������8�q]���G���Q�r>��u��za���4o��o�s�Q������
�u���������Ş�n�J}�w��NO�}����Ɵr'dq�w���ߙC))ɦ,���P+A�4uU�"�*8�=���Ѷ�k�x��U1V�4���׭����x�o{�l$���1�'�|�]����堟K�,�l�ʁ��7���
��{O*sS�۝�=s��<��\�F�=�(��+���3DY}��%�nnPE�D=�Z�pN�M��ݹ7���ԉx��&���q�<yi׏���H�<'/q��oQ�o!;<~.Q�吱=�J�����<v�)��ۢz�VI�B������ޢ�P+y�Yۮ�=u�'��O@�����7}:מ˾i]�N{4�-f?Ov�%?%���X6��b7F�3Ƣ7K�g���$ϻ᣽�ׅ���t^}Q�=���ZќE��\������|������ �ׅ;U�x�wn	;W
QK���N��7� ��}Iun�����sa��m�/���ݽ���}�֋J��*M��{c*����Np�Old��U���8եz�vU���گm6z/c1�ԡ�ɕ(d���V�y}�\;�Ż1�3^�{_p�*�A��;�`^~��6q�s{y��{܍�%��H�3rIܡT�
��Ey����������Z�ޓB9�f�w�e���v�gp��e��V]j�)�a��;<��G����Z�g�n�j/h�Z��T4��9N�X2.f�#F(�}�����]ܕ
'Bk�B����=@�{eJRfT���ڲva)�_�}�9[�to��hk�����D��Mq�w���R
ũv�^����ݛ����G�d3�Kˋg�hNV��]�B��Ko��6|��#�ϳdt��{�8n�w)�q��/G�M�A��^
S���|��G�4ⲒV��i~�(��(X��w+a͒�;�=�xx��{�4 �¦��dAF�y�|��J��(��z`��3��S(�����e��f綮����Ѳkر�Q��x�S�^>�$ �Nm{V�FzW��;5d���W�r�F��&T͓�ٻݩ�e2��=�76�=���������{�{'bt�:ݍ�8*�r7f=@��3C%{�{(�1e��'i���4��t#��oao�[Y0U�(��p���:f}���*53��'���z{�7���x`�p���:��
n=]��j���w��5g��c�kH�����~��Ǝ[�5?����0���ٷ٧S�,D Xo��R�ڑ�n[�!wp�H��`������^ض�t{!hl�-8�=r�Ӯ	�2DжI��h�<��m���b��wOXȚ{�y���\R���'M��Ը�dM@�#'D��A�Gr��\^����jV!�-�[4q�$���$��W;��Vf��{�3ýu����M|�1�h�߫:�;R]弻���+F�xxe�:G�u���!0aW8mn�poj�g�'��=���X��,��B=�Fh ��D��ʞ�=���k�-Ky�pi[�p�#^�<ɑB�E�2����3�;ޯ}�r�h0Sn���{�y�{9o�6g-��8�����{��]ZÕ�{qc���,8$�GTv�gb���14�\ܷY��J�{<H�=����
��O����/*m��7n)}���/`��懻<�`�q�����51�x�Q��ޣ��h[�o��sQ�V�ar�J�� �"��n�{xW��n�AsH+m�gZ�-ZG��;����9��΅� ���ٰ#��kz�Z��Lw�	�ۮՏ*KsԿa��Q{�{v��������|Lrr��jl�zRcũ��^�4nw�ՙ�ܯ�%���/�M�w�=��l�=zz%�S�Ak��b����v�<kou��0Eg�gP�&^%���+L��v�S�'������'��|3��s��w�d�5�����W��u��X�ge��=7;��=V���-@9�������w<1g��G��|��J�:v��+����qm���V�Zw�����.�ί��x<�Z}4�^�G�7��=k�Y�G�g���[�Hsi�U�ёb㏏�E�}Q�BQ��n�^���gJ��K(��|�[�#�28�\�!u�|�q���j+utV���a�K��n�ݜz�[�V��C� �q�[��a3T���W��5����ȭs�%D�w���CVYu{z�u���=�:w�8�^{)&��g�"��f�b��H��F�2�P�:��()��p8Y2%�q�z�UT��#6B�ɪ����� �������{������iױƮ�y��ۢ�L�OU�t�umiy������̘�C�$�彡�n�����ѹ�/onxz�� 0Lm��xq�������|�KJ�c=�>�:�o"���*޹��t�c�=RS]YZ��6�h.{!s�l�6t�c%���G�9�nøs�
�]��m ��}�M�ב�˥#��]:��CW>�9�֕��9*U��eF�����gq�L�&�2Ǫ�X^b��l^^�G�L��K�<�\�c��<Z���hQ���-�S�EF�ɞ�"�:�.N�{��dK��j�T��<�d������n�l�k�����6D1�n��m�Zon�6�I��W\�F�sӴ�fџn}<Bv�'���n��V���;]�܃��@{K�ny͔�W��V:`�sd�t�wUA)=���eM�sF�6v�&���շa���n�f�q���kpO0�[��#�CP<Vn�p��sp<�w3귞+�6�+���9���Y�c�aș���ήتݸ���g�n�=�u��aK[����u��NX�S�d뗮1����Ǉ�9��s;�yG.�<���(�Η�#��<8���v�qz3 :;ttfu�ʠU����� 8�����[�wi�:��sv/m�X��i6"��1���9�nk3�m���1��睹}[��z���mw#��d��8s%p���ۍբ�6 ��T�Q{5�[�nA�<��կ<�]+�];׳n]r����ɻc�[C�nָ{;;
i��wbz��Ğ����ۧ��n]��
���v�nvL)���܃��g':�c�v����q�r<��s��sq��ӷj�u�g�Z��Omో��sب�gw�^����U������А�{ �6���ڸ��5����ݐ�"˻��<��8�0��=O7+��u�sn�����9G�V�z�+&��A.�ɝ�{�Ź<��u���;&y��.h-
>���9�XH�[1�WU��ح�rx{u�훮��=�c=Ԝ��C���'n�s�:<�ٌ�tx$���%hy��v캝ӄ�;�+�myq�Ovݹ�����x��ݤ�'p��
=!h��v����]����pByt��7eV���!��6��rۜj�D�������Y�H6}u9{v��O� =vy�i�wS�h���c�tc�w����m��:���m��&+��ӎŹ^}x�ѧ�ӸP\��Xv�[P�vծc����&��{m��{&�v݌<��M��=Q�hU��p�ή$����\��ۙ����N�K������m�n=`��̳:8 ��nl��s��q�=Bv��9�j�紸.ڳ�HR�'��zD���n'��7v���;�n=W�٤��9����r����"��{W[��4��iݫ���]������ˁ�Dq�q�ǵŞ*�hH��o����v�ri[,���4u�pՌG\�d^%�λm�G];�=�g��.6�q�'mv.�4�����m�;sɄ�Ԏnۃj�y�|�#��ۢ3u�^�g��.|�ų��pn�:��!�6�8�����:��w��N�7)k��遫�oON݅��\)�R���k�BHw:!Ċy�������KϏG��+퍙�'1�q�s�D��u�lΐ���ų���=�lN$!gC��]�Z��8�OVu���鼺� ��R�u+ѷOq�s��d��=;n����{R�$9۳۰\���p�8Hl�rb�q�����ѯ-����ܞ��n/W-l��n�ʜ��d��n�mu��K��ۮ;v5�n��ێ�6��u�a�W���ɮ��N�7ڦ8:�U���L�c��L��u�n�S:��=�rv��\nOa{:�80��>LÈu ,�6v:9W��Lb�	�4���h�g���y����̻i���c]w;�z��r���j�m���c�;[�H���=�p.p!��ļm��<�����\�ŕ,[�om��[v��񮛳=;�mTs�S����Ƹ��5�|�.�EF���kb�8Y�궧n=��69Cy��:ꛉ7!Ƀ��g<v�ǵ����\��e�A��9���t�3�8[�2on����=��c��-�������k*�;�8DA��)�^!�88n���]���e�J�!͹Jx ��&֓Gf޸�㥲�\�D��7��j�<�Gc�ē���W\���;�v�w!W�/��m�Ƿ��w���ćm�Ї	q�1�Y��4�m%������K�"x��k����6�vm�K��q�J�������ݮa�ۺ�'<�i�uݮ�U^^s�s�d���6��n��%j�'7N��]c[6�#ŀ7e�jLu��v��yq����l�ʝv��\q�lp�á��ϝ�grU��3^G�H�.wnw'!��<�'1�㭘r���*CVh��#N����l�cqK����K��N�	�٠��{Z��hDH��i�X쓷e�=OZɺ���A#�fNxN�ې�t�J�^�r�d�\d��u˜v˶9f`��׷c���e1e�g�����;��d9:�X���V�F�ͬulm���[d�n�q�s����\�ѻq�[��v��d.^#>���G��u�(µە�u�li��j��n���%�� =�Q�8�^�]q6��q������>7lvG�n��uG�ۗ]�c��u��X*��m.�g��ugҚ�u�Y�҈z0;��+q��x�tb��K��Z&��:wz(5��N���Nu���n۞��n:�e� n�ͻq��^��u�������O�q\m�e��v�����T9�j�쉳���w0𝇐�\%S��C�!+$�Oi�\���q�;V5���眶9ɓ���6�9,�E$m�c�n���S�n���S��ۨ�d;��.{kv���'a,e<Wg�q�F����z����ByH6�)nr��.�t#չ75�c��q�F�]:�]�pm�;ٱ�;������޷>�X���;U۝ƙmĽ��\�=��β����Y[�kf�xv%�/p���+@��wf��ӘCnܛn���nwnW���aM�n۠��!���l�J�t$��y8��ڕ<�Ӝ����;n�&�Μ���A\��J�`Z�2Qəu��jhqQ[�����񜉈���nu��Xcg��ƲQדgvN�g����n�t���y���W�(�.Ļ��f2Zܽ�n�niǣ�WfiP�v��ӊck�mU��p�n^��'MtJO�uט�
}�ø��	��n��I�v�����F�ݮh���N�V��5���;us�;=s��kϖ�s؎���On���`ѻs�.�t���۲�×,K�w�۪:�
❎5J8���uoF����y�v�V�9v.{"ᗈ$mK�w�;F;8�v��;�1��؞�+u���,���Bv�^ݻ=�q@�ޮz�Y�Xy�"����k�{Z��ق����<�s�I�eۇn&�:q݄�nu�뱎@�9�v���k=��퓣ܞ�u��\ru�9����n� ��{mN�d�Bv���^OL{S��6ks6�OQ����$�<�&6��i�nk/U㛶*F�י/K��w\@�q�4�]��<ϰT�;���������Q�p��v����:�r猧e�X��s���۱�JL���.a#e��9'v�5�7i��Y�m�S��Giw/M�#�4#�	뱦��VK�koCȬ�<Ҷ�ԥ�7���
{���!��+�w�Y��˄��ܛ)��޶����d��\Gd�8��gۆ�fn`}]ywc���H�x=��a�=\psøyU7l;##�3�\m�v�cFr�qe\َ�g,u��x�x����v�5<F7�%�n;<U��ɻ��۱�۫N��*8�h,�FI-�v�z�.8	�3V��q;�tO\�$�;�m�p�0��x���Q� �u��nc�v7`;lpl swm�ǫTO�`�;Y��=�\�� �+��ɍ�Clsh��A����5��=����d�RKpu�T=c�u��{T;�I�u�6��g�����3�4���=��g�gev�W�.z+s�����.D�����nN�1Ď畇jN�s��H�\��nzj�NR<{w`����y��s��]`"�u��2u�qsgw�9�%ܺ��hS�*n1�'�%�u��^�;^�N4Blk/g�bwd7lg���ݲ����V)�y@ۢ��[����u]:�]&�Gl.!^"ۨ�-l(Ѻ^��<ގ�z��os��K�z��
Q��yz�@�d.�1�ne�����u�Mk��Ҏ{��b!�&�+�\���n7m�qr�r�N��z����z��狙#vu�pn��um-�#۰�PM\����ݺ��eќ��un7Z��n�c�v��)�J(v�Mu�����ڕ؍�q��q�<Ys�ƴ���	rÔ�
��dՎ�=nj��ggpoMŰ��u\�Z���wlݸ���^��=S���5r5+f��&F�ћ�{C�����ƺ�����ɳ�:q�:�!�z絎��m�W]fl��g�&��<<��M�4��n�ͮ�koe�t�s�q0U���ƻd�� ��fZ��6�U����vK�����:�n������91��mV�a*H�iꊳuƤ--�
Y��k���9�f���N��nװ�m�F,l�{2��T6��p�N9�V��v�����)�t�]ؤ�8��5ۣ���b�I�v9�y���<gX<��Qٴ��k�@^b-��=k��<c��<Y��n9x�F-�srsۜ�GGC�1jL;Xͼ;�cuq�5=uў��U5k��)6�.�i{r��ܗ뮛c�nţ�7�λ���i��gv7IV�bd;n8�j99�����v�����nm��c����R]-��\]�C��/IZ[R�UjV��+�PQc+aP*#
���H�cc8�0�V-�,j�eD��
���*���U�*��ʕ1�5�b�c�Q���cQ�6�Vb�%b�4QA��TkX��Ym*F�+Y��ܰ��i)�C��a�4E#h��U1&!��Fi�ܸ�ѵ�T�T�-��
��0�`�(�����e̦1c�Ub�m���-+Q��B�J5��
�eA�K[A�+QTP����+kB�J��Ը�LlDEB��j�3EQ9k
ZcS-��b V��D��CI1iX(6��L`,�X��r�E�әJ���MaU�+1UR�-�RТ0�X��r�XV6�cW-B��F�H���l���(��J��iV��X�2�QF��8����. TQ��mZ[*T���(���%kB��Rط�Q�wm�c<w=���_�S)��I�g0�Dew��g���ݷ8�h�kOm��"P��X���wk�n4%��.9a���;��>�n�mɵ��{D�5���?��M��'R:ڭ���Ү��7F+��8]��q��i�ɶ7v�zyN+g�$��rwT\�7�����"�4g��;/k]`�Ϝ��snr�x�<u\r��͵щ�Ʌ����m�O��K���Zu��v����lGK�.�/3�r�H�j纻��s�#�W�G]����OC�9�v^r�۝�9�'��0��F���qG]q�.��^;vl������:�g���t4�ܼ�:Cms�n.�v�7T���9���#��u{��ݍ�$vcnk.�F�֫�ʝ���U�<��NnϮ�g��]�^l�e=�TW.���sۦ��z����C�c9pp��/�q����`A{��ې^P��u�;\ͽ��� =a�=�@����y8Jӹ�0�q�͞��{l�ά���v�'n������V:�Z�Ϯ�K����I���[b۳ηq*�q4��z�y�kZFN�	�����a�YG��ţ�.�Vc�; <=tv:l2�����m����f����M��	l�댴�:uH�e�v�v�؜��]u��'c�n'��Z1�9	�ݯ�c��W,�f�ڝl��zݢg����}���l�K�@s��67@u��a�r�O;��W���[;��"�;u�w'nnU}�R���sˑ�vڇ��-�v� vM�x�Py�۱�ٓ��1ڃg���=N��X2�k�,�^���ּ=����:7Yމz�K�t�M�����iaz��v���pmֽ��vk�v����[���6^[v�ώY���v[r��þm�?3����]�j.b�i�b�N�s���"WmZ��.�v#��r]h�f[gp�i����;����n��nFk=	�T��Ϯ�U��WjL��nK�����ݓ�v�y_�r�s�P��G���;;�<��7p�w*{"vpeݶq��lcg�1s�ܴm��j�WE��K3)T�m�!l�`��Lr�c��ɍ�g�aN��{r��	���v{��n۷��ġV��U��2�."�Jո.R����F�V��7�9C!��m��m��0{m�M�`��6C���9�Ns�>�(�O�C`���Z�y2I5u�"�k��|M�U���[;���H��6	��&����|z�*Q�VnJ�A����A>ܾ�O�;�>�(*KsweM��4Υ~ƑI��
����$�w�I$�yJ�w�ط:��'���TH#��jA+��A�aCb|oWdq#9�$�ٹ�	�ZĒO������ި�P�M���9 ���h��$��ڡT"�Fu��X�����@�N��$�7�T2�ܜ�� ��b<���7\�ms�Ͱ�dI�=s��Ȯ��x�v��-��ձLD �Ce���̪�α��og��²�-�#�_MA�\�q_x����)ɂo�$}�.EI�B���aU�`��wP³_���*tѺt����G}x���F�kB;��i�F�M�LS<��R����v�˕fwscgu��fGA#�d��$���� ��Z��Y=QNo��6`�$���b�=YN|As'��>#�Z�ɢzUqt�������Py+�4�pʈ*j'o�'�VtKJŨ��� �	���O�7:�}\݃8����A�|�}�!,%!����Р|{�:h��T���5U"I'��v��{7?l��%�O<	�I3X���q,,�.�>��s�۴��Ӭ��ی1������������C��|؀�gx�s�@'���ٯO���0D]kg{%��������v|`���A����$w^�W���8UL��3;4���|����>'ݛ�T	>��ط?���1z�a���%9�Y  u����j��yo��ɹ/���{}Q���kw�:R��cA�WbX�W����BY����2�rf<�/+���ٹN�����F�*!����)�ӌc�����H���v	ۂ��Cl(P��X��d�d
k3� ���H7��TH$�V�^�U��a��V��ٝ�$TJ��M��UW�@�*�ρ۔zz�n��ꚪ ����>$�Z�[�0�K�g�J�e����՚��GvMӸ���kےw07F	r�cp6�j�q\5.�E!��=�v��ݳD�Zě�Po'f��L��O���T	��
�d6P*�1��A&�"3�
��	c�sT@$�ݵ@�?I��6L��r�u�j�d�nw��J�[e�_���� �J�FhJ�wٽ��#�{j�uV�$Fj*��l��k�w;Ѽ&�K+���emȐH3]].92D��^�dFJ������c�:���^Nd���UNV�.;:<�>��q��W#m���k�Z۽*\z&)(�yQԻb�+��Q!��kI6�j�>�N�%(�xQM����l��G�]�����,]�6�n��vz����D��UWJ�F���-� 5�p[A"Aum�h�2�y$wnz���W;2��ۑ���߇��+������^$���$�H���,�	�s0Q����}Ӗ����B�4�E!���g�Q#������^��'ĒV\�|��Mvz� ���s{@��tPch6P*�gc�|O����|6j;7�u�ˬ�@$��$5=�D=:��BE6�:����72�$t�;�|
��>$��{&�'�s�f����^"k9�
�H�(�bQ������OU�q��b����S�B�>���5^�����wN2f�/�0;G��Vي���
b�?vݮ�9����ى��׽�������Y�K�;�Cg�_A�>=;�o�%���tC$�ۅ �bQ�p\1�[�kp;��z��۳x5�5�`�n������v��ug�.���O�'W+(P����6u�������\dt��5�`^�(�['����s���ɶ����6�m)�zޮ��ϫ��h�Y�*��.Lv�l�`�G[%C���Uy��Y�r���L�oh�0;�\5��qQj��<�T��IN8��3{nYqv������Hûn�'����~~;�Zb!Co�3����͚$�;w:���S9�ctP1�n|A.�zECU��p��U^���|V�!d>��V�>�]��׈=��TFd���Wyb\�9�V"��Pb߯�����D��t)ZQѭ7�`c�̪$��Ϊ�<+�V8Ba@�c�7��uՎ9=UB��'ݽ�T	Ou��n�鑕�ϳk�E���C�A�
n=�9�|O��[��W�m��G���گ	۝^�g��1[o.�K�;��&D8��D)%Ys�b{c�ln��kA�ej.N�6���~~����I��A1xx�vU
{��(�=�"ẢG:�Q2�񝻺�$����@��k`�$K��B����N1 �<Li��l������9*	dn���wume�=p#��y�����"�bF����9!\���A��ަ�d�O����Sy�}�I�����rA3�N"�4#7�bs7IT;c4�l7UW�@��=��Jr�_݌��$��Ϊ$�^���>��DX�Pbؓx磕h���$�˚$޶$L^�T᩾�r�⻘�0�zExE����5��m��I ����'`jkX�Vnj�kĒ_V�H�{]U�}�7�n�F]??~b6Q._Gr���ώs Yϱ�\��a�ccngr�i:����C�`����c�;�r�|�� �|HW��G*��l���;5�I%��iS �J	b ��Tj�*����$�Յn\�}�#�>%��'ī��<ZB�K��|+&��&���2�A4�B�L��$�AY��@�&i�һ��u_QQ��6�ًɻ$�{j!�S�����ԩs�ꃍ��{�*Z�B�g���j�_G��+���4�ZЧ��u��r�� ��u"�-��M&�pT���؅�b-jn��I�]]TA��Y�^t�X�ݛ�|I��rO��-!��6$�9�	=��#��TM�ǌYw]TH'ݻ�Tg�bbLEW�䓍�W��c�a�kS�G�;Z�l�6�[Q�۷e4�0Ha��#�_&�� oǾ�r	$���h�}���Fy���<~�z>��'�`^�x�O��A`[�v�Q>*S������i�DUueQ$��Ϊ ��r���BM9�;�xf .J "	�uF��������O�h�yH�19��ݬ`$���O���ڢs�O$u�8Yh��x�~hC��W�wu17uTI �ol�>$�W8��D�Wq]d�@���@���l��P�n8=��{z��r��^���r�����)w/mT{f�xN�����������|��T3#,4�m�&�uvU	3��I�/��f_t0A��dP��mP ���9=y[R�_�<(δpdC�����Nu��2������g�t�\��'f���o����!�:���\�UI��٠��k�I]���wԞ�mQ>7��4J�Ȫb-�P"Q��bM\wX3VSQq]�H>��T	�3���FN�<;�4��a�l�!��cg�g �3|���\R�I�j�m\^>�q�4���$���$��*
� �H�uF��B���уц��P�L�Ϥ>���8�Ċ��'C�Q0�H�ਆ�K�� �	c�T�zyVEM��$A��s�	!V�U�U�ngf� ڎ��Խ��m����X+ycwqa�-�]P�Q�a�d�*��b*^n��pn���oh���Fo^=�'U���ӯ�L�W A��tc;�ӵkXQ7mLޘG�o3����m�⋳�)��F��mŀ��e.Z�f%����!팻j���uv�Ħ�㺍ƍ��}��`{ r&�Y���m�ݠ���#Z���܍�ʩ�ɸ�v�n�ۢgR�q�w1>�>p{I��{LR�`㓛ka[uĜ�L"��H�و��.�͎����y+`$g�Q�)�a�����=������\�\4�'����<a-۷�`��"a8�(q�7��,4�m�+�#kr�L��$*v�lݐc�B�۪'ă3��n��L*�bؓX���2�������h�y����fw��AU�U@�i�:b������� �
[,`$��H!��ɾtH�޽��\�9�z��H+P�mCPA�p`��w��r*����!�ӟAguUH��No%��Y�o�!^/g���!�6R-��UוD�{��^3��ñg5I���I*�2������^2�A��edu����0�"GU�n�����r��y�������kv}�7�l2!�1��lq �κ�$�ٽ�F�8mv�	N�A+3���b�|�0�6l4��?Y���~��ge��K/MȔ�Hǡa&����n��ܗg.�oe�	�}}������,_m��q�n4C�r����t��N§���ĀO�
�n�ĀO�w�����yP��1{	�Z�^���y�P$1�o���{��hH�Ե5Ìk�>וT'�{f�Z9%`bi0�f��;Y�ᨭ�6?� �`�/w��%���4���>�N˺�!b[P�a�PH޻ڠH$��rlA-�D�jMc�^=��5�Hs|䱗����;�X�����_ �xQ�S5�v�7nz��8N6���T�b�ҡW1����NN�^:�'xU[�Df��A;�� ܂V8��S9A켪�}�ݵ@��(�������Kw�H��w�]m�U	�>��ڢA ��r �v)��&� 7��:P���[.,8�s��D��H';/�4�qۡr�Z�w7�$�����<�b]�Yҙ}�d;{&^3J�n���9$M�`jӌ����������q���V=Ҳ�����'�zA�n�JO���{�`�ujԻ7�oD��Gz{����|Ο9@5ﻷ^�۞�,P��O���[S�n ����X����pX��o]ד���aͲ�˜r���M�zjj� `^��L�L'83�Ƽ�[��X������ܚ�D����s�m�shz=�i_|n��a˞>����C�.z���#�2z�4���8�
�7�����������w�w}y���]~[�7=�Ӗ����꟯�������:}�|���}�_-#�W.��ع�^����؉I0�lx��'�p��˅��e���=��X�p��V�2v��{�;v��7���zw����r��So������pҮv.����`�_QFnn��˔���u��Uއ��a��;A���N���W���7���>dJ�wh���bӫj��r��-�3}�)����A�jc }�����`G�k���޾�uJG�7�c~�M� �N�� ��&B�9��=���m~��eNO}�_w�^�
�����O��1Z�T~����`�΋sT;�W�����n��e�j+2=�_�F���a�5|�K7��S|GHu=0�q���w�����y	e��t#��]{Q	~�X�l<�s`��vP���e���2�I�r�`ue��MCx��]\<��嘉FvuW�`l��{\;yg�/c���}q�Y˜�q��Gw��EKhT��@��S�&#�dҤ�+e�5q5J0�R�T-��m�Q�������j�+�T*Db�`�!m��A�#R�Z�Z±f2�%X[B�`��@�%�E�B���*��+j�1�Z���J�L�TB����R�ŗ,[�Z
VҔE�r��إt�ʉR)mQ-���b����X��˂�UT���`�V屆R���e�4\d�[mm�c�F"�Vŋ��dW��
*��������)m�ڕ+e��R���F*[E�b,��DTbj�T]%Lk!�8����R(�*-Z��Tq�E���E��WȨ�KB�B�E���kR��5�am����Xy��T	$��rn���$1�oՑ�=�Tl+���]ȠA5�$Uwee��+��_k0	���B��+��2����9��*�U��wբl���9���۪$�zk�IUݔ:�{�K}�6���1����b2&�*"-�c=��f��Լ�ӑGS�&�W��sU���;��s�P���뾪$��\�H*��hǮ�3�7��벨�|zk\�Dg@�Y ��4چ�5�
V���z���g�-w�ɮ~�O���Auo�*��dE^��yD��n!D4�z�Ē
�۪$����ֽʜꈺ�A���w]L���͖[M���������Y+��K��>$
�˪nol�L�k����㸕k^��X){�߳�n�l+O�=/��ٮx��LzWL�BAFE������h^Tr��>��L��i�$��rOP6�1pI�a�'Ƴk*�۝4���8�y����%f��x�yz��h�e꜇��R.O�����6�r�:Bt������%�/%����+ع��C(8m�Ig���pT�㝔�U��z��ss�l�ѽUd�Cb���J�ڪ �Q����L7
	�׹T	�YM�������o��W�UD��n�uQ ��%��ʳ{l<��P��.I8s��WeQ$�nt���;g!�R�T����	 ���۹�0'�~H�pb!�)�v���67x��˪�Κ�7�j"�+$/j����C�!s���9��I3;�|ky����P�ӭ��W�'ss��$�3|�����ա�i8b3�ɝ��4)ۜ����!����Vj0��HCE̸�IW٘��،)T�����2b٫�ShY�@�a=.��3�q�]������'8t)�qV z�;nfݸ�Lv�\�ڹNl���έ��ug{t�#�c�%�vN�q��Jۗy�����B`/^�	Omli4b(�5�#=.���k�v1��d��3=� �S\;����c�S�hç�x�f�7k���=G��B�{u�}��v��YQ�uی���tp�m�r�]g��R�ku�w$��\�V���,[��v��vnӋs�4�X)�<���sA1��	�>���{�:h���I�!��U(d!;��^$��Ϊ$FE_��	�T
�kv��4��I�ٜ��\���w{:��A��~�m�ۘ�,.���%��20�(&'z�*�$��W9 �ԠVpĲ ��nx�H۝U�I3u�I���AB;	8A$�����c�r"���ʝ��J�Κ$�L�t�� ����Mh��Aۑ��3ݓ7T6#iD��^nPڟu�I��:�����
�2	U�^�g+����B��<H�Ҳ.*
��Z�>����Ճ)��v�դ7Xi���康cO=�D4��o��ۇ�q��{Ēg�\�A ���ꉅ�p�MnN^�ꪯI�3��I��	�l�L1&�����)*�6�DD��C�E(����p��"�#��1���y
��c^��$�jt�@�w�!�[�E�@��Rq��M,9�'��+�̟�A�3�H�I
���Q�N�)[��DNg����F8A�p�*�Y�ĒWӵ^3Y�hn���|fs���{=B���0�(&'�׹S�g#�6�����h$.�ʠO���L8������0�ws���C�p��%���܂OצA�f}n+�'���7ĉo�	Us�(����@�r����yn��L�	�Pna5a����o�/2�}�Ϝ�����unQ�p����~��? �p�����$�AY��DGf�U ]_(�Q�*w\�I
�v��B�3�\7	�0U �o�Q��3Wg;]�U��^$���$��;sd�E�͍�ߍ2���$�U����4	$�9�}p����5aqWS'b�oY�q�^<��6Q�%:o/o�Y�Q�(Q����/J�Ş�0(T>��^�d�U�A�߶��`�W���p�qTr����]�X�����+����H��T	!�s*�;E��UOeQ%���-�PLH�{U�H���r��`B�`��UuCă�ݲ(]�9�5CBޫ�aQG�9��&YpJ�{/\>$�\��n<F�ŵp�Y�z�nk�$�A��P�MG�-�5u�Ds7�hO�w�"AkMp*P���?Q��m��u ��%B�~�߽��:����~v�3R�ְ��g!Xq�yϼ�Ì*J Dz�����=:�y�O��H�*|��xu�+ư(�����PHx�]{[2�u7o8Q����Î� �v3��l�i�+�Y 9�E
Ag����������D�
���_>�ϯ�n{�8��aXV%����Τ��������op��㌠C-Ab( ��Ϳ�@���h�����q�����9Ґ�R��~}�����T�~����~�&��m���1;9 �*�6��A.��@�g�3�0>8?~�ܗn�Ɵ��u��4cqMɉ˚�>�z٬�+�5��@����*{��u�+
gǴ���\6ڈ�#����2�G�#��|#7�H��>��<;?F��Dx ������P:��Z��w��op9i������6|=ΰ(gvx���'>:�i���gt��0�]�;�@��8��cq�R�h#�����-��� ���}�v�Ԃ�Y�d���� ��IX!��^|,|J����"z���o��:��VJ��FW|���N	P(���*��@�� #�W_l�`���<;wE�Aϸ;�g�tY 2�����BҐ�`W|����*T
�&~���gY+(�P�����}ﭏ���M�H���#�=���:���+0�?w��9T�!RQ
�<����βVT���y����ϼ<H,��F��op9i��g���,����v4��f��@z���{�~�3?{�����YY+���{���%B��3��wp��
°�(Gwg�,�]��8������z�>�>�����ND�q~���Q��a�6(Jü��6z��HR�>���l�i����_�15�H.��{�@S�,@��g��wp�:�R
����:���|Y=�I��R>�E�X�UZ&rL��2MF�"UA�[A�j����4v�L��j��v��=t��?���yjW�FFM	�N\�Ø֋��/�}:��\5SZ�Z5�n��Q�]zh�c�bq�S�󞎹�s�%�{U�`����֎�K�.�&4�vn��nu���|[gϧ�-��v��7e������"��i�1���u��J��늜�p�cX����0�m�UĻۆ���Y��xY����\�㣑7t��:㱨��7G&�n��Gk���dź65��+�tc��6�u���)�V6��Kq�H\gp���IӚ5��۫m�^,c<��ml�Z2�肍�u�/�����5Fg��+߿�oa�aRT*JV���ѝd��J�C�}���t#�Y�f�a\���|o>��J�m!m�}���H/n?w5�R�kM�yI�'�~�͝N���Vfo����^�����g�O^�]��J��*$�)�����R�����q'B>���>���Цr���vg��w�>�D��o�/�e�k�p�D�9�����z����=���$�B������|~�!\P��b&�w|#<@T��&~���gFJ�2T(����H��<�����T4B@��!��GÑ�s�oa�ㆹ�Ӻ��O� ��;�vtgY+*J�~���p�b"<	��5�L���6�|P��ϱO����p/	�ޟ6�Eyޝ�&����Y�N��=��Τu�������{82T5��w]���<H,75�s��XtaXQ�ID��}��;� ��ߦ}���*�|�E�:�Jp��m��;q�z{w����KVz�u�]�n�78��������娺�SF|)�7�l>z��R
�{���!l�+Fo�w�r�@�}~�����f&��<�:βVX�P>���l�V^|���L�mDW��>�nL�G��H��u�$��7M��2����7z2�L@����0$t�7�1�2�tXW1��ˠ���ݻX��Gt{w�����Q�?�������|��s��3��@���߿�u �Z��~��rZA�x$���ų[|"+�7��AA����Z�sZk��4�I�߽����
��R�;��p*IP�+������'��.[V�w;Ï�|�Dy>�϶u'D+%eH/�w��N%@��ߥ*��t,�,��}���{����XjB�~����ii
�i�;�9N T��>��7�]��G��{�����d�T>�<�gR�k���j���k35y
Ì+�~�{0�(�ID+���l�gY?m�ۛ�}��q �y�;��:�X�_��7���l)B�>��7��
�����/��_�9x�b:W��\v��E��ݚ�H1�<�6vf�������]%�&�M3����I�{�ݝN�T������{8�P�*IXY����C��o�^뻿:�}>�!Ě����:��VJʐ_y�7�8%@��_w?\�Z�h�
����� �Q�阼� }��ȭ)
�[l������
�|��}��dx�>� :tk���}󜑤 �#���)j��d�M�\�:ì+��y��T���V��vE�Y��>D �D�Y�9���n[ʮTԬ�تzpG��D��o�k�F>�7��U���w^.���3�>��gX{�V9o�h���K�0�5o������		�s�@�J���k�;����m!m�~���ïX�q���� �&(¯ ȯ���CF���wy��5t���d��%}�������RT���}��C�:°��Ib{��#��*ӝ5���xG�#����Ͻ�T��·/����k�P;��~��`V�(Z�{��8�|���������Co�y����R
p+���nH,��P���l�����}�����aL�!�����R:���lk�Sg��݌Q\Sƺ�]f�ܛ�?������֎�Y�W�V0�9��'�(�a�����:ʁR�Y�����tB>�{ib��L���ٟA!��a���7=`V����35��k5����M���l�v VVJ�nl��s���s��}�O�����%H(Q%as����u ��
�����$�B�X�������ه7�s~��{�D ������Z�ќ�ÿs���
5!m���H=�*A_]w�]o�wy�~���J�=��7����������H���|ߊZ�Al$T2�W��>�ńb�����|��#��,B���|�p�'YP(%@����@蕁Z��w��op;����ke��X��6��}s�AF+�e�=xd(ȫ�ת�:b�
�S�c�=�~���ҳ������t�sxa��ز�?Mg� @�?R����:��ZK��g٪-\֚��'�w���:�@����2W�w���^u�_|�\zN!ԕ�?w�=�:ñ�aA�IA>��>�ԝ�VJ��������Ĩ_Z�y���s�K8��"�1�y@��3sd��c�9�]����5������d*u����ޭ�Yfb��_����a���Z���y�}��)JB�`V����s�( D;?|s���3��	< ��=�p�?����D?{�l�IXY�gT4B@��&��
��F�>����
�\���e�c������8��e@�*����@�T���]~���KH)j[�u�������n��yz�4�M�É�E���ϤY� ��d���׽�{��ĕ
$�=�[߷��o�髿�8�|3���}�$�B�J2��߷�8���}�N�6�b(<	��@�7��upv���������vs�!m!RMyϹ�
ANeL�Ͽng����כּ�Q���Q�� _ٛ"�G��U�U��1�Uni��C�;W����I�
���y���u�d�Mw�=�����A*���xu�Vk�u�=��p��JB���nz��$���}/GX3?Xj���Z�6�عFMpѼ;����);���csԇvf�UZO͡w�Ȣ{J�}���f��$�ΫjsM��F+�y��m��p�D�=ݎ���@�;fht�T���K=$���'K�6�;�Em��u^~�����u�?{,����ή�̡�<l�w{�{i	�DԸ�n�e���cC���f#쩉}+�76;�HЦ�\�)p�^X���հx�w�0��w����!T��pq������Gp��J�э~�N���Or[jsAP��Я%����#0.E�/{��4��]��Ɵ��3�~z9ꜣ��*�>�؜��_?,��:�a���/r���}�-�{v�2��݋tL>X��<^�]�����ōq�	ˁ�=ɖݕ~A�X�s}nM�a��J@�<x�}����K�&@L{u���Lr�ֱ>�z��=zb�P�r{֎�$*�w�y^q�+М�n�yc�Q��gཝ�E�M����֗{:��{o�;i����|�-~��7�^}H���ӷ��:�,��g������Rb�gM��4��ӎ�l�/�B{:�¹d�N�\�ܩ�9^�A�����[�}�����;<��{SxL;����@��Y��n�BS7w�۔XP4�{g[���w�Jk�\�n�oW}ަ�纰���<��x+��+n���,�XB�K�a�D�nt]��p���\'���d�iQ��p�)|z����yڼ���zj�۽���[2pZ�T7>���u��O��{����j��,*�_�e��3���UPDGL�Q���R�Z�"�
��&
�kc��"�5�スL�Q�j�6����s1IX��&�(��֕���2�[F"(��AAVDEU[K"12���(����.
��J�ڱ"�Kl[J�"TĬR�ƓME���ELf��-�9kV1e�S�U`��V%j.[���]R�a���mQ�X�Jc���F$kUd��Z�D���%KP�+Tc+(��R�����QeE�1H�J���B�Z�AJ�",Y+DPAQ��jV8�dB����,�r�6�������EJ(6� ��QE�cS�6��(�m-�EU������UU�E�-"�,U2�*(*����VF"֫��ƔH��m*�E�Z���b��l��"�a�󞙣5V��76z�exRq;�zM��8�wX�)��nZ����G\�i�f����۬����n6���)r����!��ܥ���V�q����i69���g��q�����Q������o;r�.0['�|��/gOm6��Le�Gp���ō�8�ѣ��^��͛�;n6n�{N�W��8�a�v�JPu=��`::���б���ɷ����[�۸��2n����cv�OV���8���;!Y5�n�w=K�ؔ:�5��F^�wA� ���tw[3��iI�[����g���m��������&ľ��n��G.'�盱�����v�s��n�u�8״Еc�t�o8ɐB��uۮѡ�;��ЬM�G;n�9�^wu��Dn��(�'�ޝ۝�l�r��볗q��'<�\�m��d���8��]Z�(w!����]�:gwN�)�7b�wm���ꗳmѥ������4����)���W=I�;5�N���6��8�&�L�]ܦ�g�ܜv�y�Y�3�٭��� i
���î�7:��3�t������W\���$���V�ȼ��nx�^4�c���V�A�xOU���n޼�f��/�  y�v������;���-�۝����n�n���$��
�1���u���8�����^1�h`�^�����sp���ٸ^��.],�s���x�x�1���n,Wn�s7nʐ�h�r���d������h裵/F��l��<n*u�y�	�s����y��	����qp�p�Sp
�n+y8b�����E��v�#xnMx��6e�x�VSs���mW�N�m:�ƀ�g;9Ȇ�ph6��Ն^U�'Eͷ���gx�vvv��X�&��0l[gɹˬWGGo^Mћ����̓[�M][#���-�ZA�qV���w�kI��b��!��r��f��{s�
gm8ѻpvs��ֻc��V�v{p�$��%gn'q��J&^�ӎ�.�����S�5�H7��v����Fb�]�۶���:�`^�&�mɚ��5dݺ�7.��كmǜ�`��GL/B�����:�{|p�bS �����}��q��7�+g��՞�W�ldT];�;:��[�y��p�=��\�=�s'�nγ=o!T�]pz);];I�t��=c]�n�x���1��f��8 �s�v�v1�nt�ۉx����Cv�z������u�v�U�� �0�k��Gob�T���*v��㚯����w�5E�����O�'�}�gS�����W^s���%B�*IXg�{�p��+~�����������/�C�0O|�l�N���+%]~���U��EpMD� �B���T�� X6|�:r��:�g�d��!�HV�+u�>� )����$wݓ�g�}�|�}�@��c��; ��sg�}V���WR��֭��+
���{0�%�3�=����H	  DK:�g��]R�q `"���Ϸ�
A�H[,3���,������m�&�%��
"�G��>�d:��o}��oW�}g�Dx}w2(�R
�+
�~�:à°�|^#�{�G�t}����d�hG�>�e}����T�}�N��4ѳI�w�߶X�-����9Ґ�|�Ѫu4t�h�� �VOmW�$W�(�YS?~����td�
!����d#��P�ϟbL(9�Aa�HPWl��<Z@6�Y�۝�L'F�nM�z�\�۬��B��}�-��6c�#���ɐ|¤�T�B��}����N�� .��Y _�G�m��������3�x5�[�����K��߷���Jƶ����^�^#�f}�,� |�>�>�m�e�2�Q�B�K�Ҙ�e���7����{H�8-{ʮ�Ԯ�m�����
���}�\g���5�?u�׍��BHI�������d�Q%B�+��}����+T�Gӽ�E�� #�/#���m��F{\��N%@�<���宜���p�D�9�?{���jB���߶q ��������������*Q��{���������D=ߞ���tIXS�͝�WE:֭��++�����v��WM�w����#̀��'�s;d_��JFT
D�{�~���R
x9L�_n�[�^G�>����G���M�h&�m6�.+�YG��Ϥ�u��VVJ�����d�k[���8t�C�$�?}��w0�

���{߶u'P�����߷�8%@���t�>���K��d4��@��(��w'���xN���4I3��Pemn�O�?�}���]Ƶ��=4��Vsϼ�tz��Ԃ���w��HZR �����@S�=����>�y��5��ng�%H(Q��߶u��)����q�E�ӮC�:+�}�{0�*&y���7�=��s�����gFu���%@��{߸u�V�`V��߷���m
ìn���룟,_x_m}>s��"��[��j�[sCm�'{߼�gR
AgY+�y��H(pIX2Mu��U�������N>�zZ��=����-;F��ژ9��9�F>�9ډOUϫx��D���C˝����v�S��K�U��XC-n���{�� %9�|��aXV�����:�d��������E���a$�E� :��>��6�������^z��H[@����9�B�B��[�{��q8 T����~���X�<�������?�7��{���'O4w32�d6$�y�c ��{��ą�ܶ��<�����_��߸u �;��y�~��JB��=��ۇ^�wy�s������7?6���B�uhy%���#56C���C����-�!�Yg4���چ�.;�q=[����v VQ���W�w�d�AB��.}�}�:ñ�a�}��O����Ot�&	���gRu
�FVJ�?w�I�N ^�~د�CZt:8i�+������G�\���Q����w��g?����`V����H)�@�3���Ă�P�{��㻭}��>ϝH���#��|�`QXH��u�g�XW�|�A�H)*�}�}��u H���}�t����� �!5�Z������H[a�}�w�u�=֪�ۚn�m8	9�۲,�Y?'��C��H�&����T(���߹�!�V� Q����h��,���U�X�V.\��]�S�۞�4�p���r�Ǜ�L=�7�|z��؆=4�׵s�&�l)9���N��z�_�x|�?�VK_���{��*9����3�2�u�:�Xo_y�a��������EZ	�WD��t�P���9N T��<�ng`�R
�ޯ�Y��>�!O{l;�9B��\��vk�3ŷk�R�ϲ�g>ni�z��r�8�|6��A�p������Gj�{���B��|�:�%e@�H}�_P� �G�oγ1l<��,����ZA���3���ǣ��}���nj`��dX#�ןH�,���G����mB�f23�'s�dQ��D�
$�.w�y�u�XVT���G�����fl�۝�7�8%@��_���CZt:8i �����(ԅ����l�JB�HV��]f^����c���� ���eL��}�u�++%B�{��gP�G���wJ�-�^|,�#{�2=c�!�z�/���<	�@G�;>�gc:�R
��϶q�R���g�t�G�/�`'��!������Rۯ�̾kU-�hm�������q<��d��|�{9*y�������8~&��J�~taXQ�IS�=��:��VJ��Y]���ܜ�P9߹��(��,"��1ss�'nTMN�7��yC�jXw�5MPlo+��oi�7v�.a�;��+���ض�ב��L]ؗ��~���=�t��@PF\��˵��[5؁�ѯs�Q�`,rn�Y}tc�5w�;y�-�-t���s��B�GW:G��k�m��\lX���IsƋX�Q��Bu!���%�ƺ�����KM�8�3�//Y���N.9��DQ����ݟ���vw;��<&�\�nx�ӻ3�]�+�.���n^��/��\��m����-�ݯ,���n��c[v�q�j��anJ8��FnZ����NT��'o6yl�n�+@��ݷQ ��sG�!�a��q�Q ~!
�{�ã����}��l�ii
с[���� ��4�ܹϼ~�� Y���:βVX�P>��}��u%ag��<3��m\���cF�����>�"#������聚���>��A@�*����`��Fo>����$x�#l����e�������"�Ԟ�f!�چ�1��I�{��N�
�2VX�]��w��%H)��/=��5�~����7�=a�°�
���s�H,������}���*x����M\4�^!���Ͼ����t��G�H����9�B�B��]���� �+*g�s�ì�O���oٝ��A@��o�8�Xw^�W���n�����<���80�%B�Ϸ�:β:ο_;���Ϸ������o���R�+R����H<)K�{�u�a�����o��~�v���c�.��$n6
X�;mvD�����cMm;�w4�?���?�nj9���i�N}��l�AgFJ��]��w���
$�T��{���8ì�n�Ϸ'z2~����Et�Ȳ=`������y��P8s��z6�\�R��@�Jßy�70;��7���ѷ���Ev.!��2�ۉ��z��W\�gE4	%qƧ�H=��E��;����T�q0���j5�0���N2�Y�L�h���n������ ����vs�����`W}��{���Q3���gFJ�P|�<����w�k�>��G�>��h�	H��^Cq�w���p�B��V�{�g�}�� " [aa��%�NO�0�u+�����{����e!l����|,��"�s��L�mC��Q^Ȳ=՗�#���in�}�>�}�G�������
	*V�{�q�F��*J�}�~�ԍ�?h����w߹�x����Y_9��ܜ�P/�_M���\4�Ĭ;���ã��H�O�H�C�|`��8�*}���+{���@S� ���w�ۇY������� k��E,�|;�&�ko��߳���ٜq\n�kr��희h�]��eLt�6�Ze�T"��o��m&���х}��oa�%�T��>ߞ��gY(ʐP.y�p�D�����{���9�`y��op��H[a���7��
���/�ʍW49n�m8	;�����YY+5������'�6�s���*%B�%as�>�����=�߶q'D+%ed����{��-��M���D �p|
���q�V����q�ѩh����x$�E ��τ_���gc�Ap�'���Ϥ�+�};f���æ7?*7���D�|ݣ�;��زa�,.C;ҎG� �]���/l~n{���	#����*Q��s��ì��YY*C?���gP�J��ݜ7��)P�j| �\�� 8���9EGVV��Rm
��Xk���gFu���%@Ͼ��@�J��`V��op>+�=;;�/m���d!����N}��f�|(\�-L�mC��Q^Ȳ=u]��N�VQ���W^�����P�������?{�k�x��V矻�!�aR
J������;��eH.���ܜJ@?gof��>ρ	�ne6�z!f��X�=��z���k�6���:��
�G��o����oM�����;���ã����{���gJB��[�?}�@S�!�#_�D��� 4�������>�>L�
���߶u�+�����C�.�5��Xu�|����r0�'��~�������z�����l�Τ
��y��8�Ԭ�~~�{����x'w�.���Q=����q���n��j��O�O�~�͝N� ��W~~�{���%B��/>��	�7�s������>H,=�*J'��߶u �teH.����'�Z����a�7�(Y Y�W�{ �N���'>>�(Z<��vs�������}�@S�J VTϹ�ۇY����^m����r�4�̝�GF/'�	=��J�<�(Y�	}2��|7�g�^w�z1�;J���*k�C��v��Wg������v�/� I�A��D7��~��:$�/��?5�\�1њ��0�
��Ì*J!RX�a�����}�Q�!W���\砏@N��DA`u�
5�����R)l3�}��,ߏ�G"˭c~f�~�r��i-BEBv�aΈ�K�κnCs���Jˍ�v�\�E��/bNF��GZpچ!Ä��d|G���E��e++%y�}��2T,IP�+3�}�!�V;�zy�~��?	���vu'D+%���������Ĩ�_�����u����8%a�w���(�
����3�	��$U�<�h��>��8�R�VT�\����>�>G�D���}�ܴ4NfG0�|/�љ�.b���g��7{0�%�>�<�p�A@� O}���7}���� ��| ��k�9�����-��\��ïA�T�#�$�a4`��E뿾�A���%�u�}�>��"<	s�2(�Ȁ�*Aa~�?{�u�c
*J���"��Ӗ��m%?-��G������]�������|[sE�3R��H,=��O��(�@��U���lNf��`V���� )9+����gY+(�P�����u%a۞q�}��:̏���%��~��`��2�I
�=��X��2�ۖd��{��9���u���f������ڍ������x�a�߇���fyIE����,p݃�y֍�=�у]��u4[���QS4�N���j��{;�u��r�N�:���lV)5�;t�)�K�|~V��n�Pu���\��ܒ��u�����о�\ҋ�۪4�v���oa���x�8"����mu�Ÿ����.�j\��{=v�<Oa|o7c\���D=�6���̻s��p�:x���ۨ�oj���&�n�v�Wi����Kջ��v.6s�$�=f�x��8;S������cn\ѧ��a�F�=�{F%B��V�Ͼ��u���X%@�����dd#�9�}����_@oh�'�A}���p<��iaa���é�r�ɗ�p[l��d]5�#A "<	������'��{>�����IR�\��C�:¤�3Ͻ�gR'FVOOM�������������?A*��s/覰tp�"V�~�a���cR�3��}���-
B�`����)��e�;�g� ��H� �����ۇY�J��P�5��l�����>�?7X���Mg!�a_=͙ѫ��<��=dG� #��{�
D�����@�J��`(��L������|>�ܘq�������5m�5��yiĜ�y���
�2VVJ��}������u�]w��"�D����9�!�V0�,O���l�Ad�+%e{�=��$XO�������.F�2-�B��-1�.6Þ7"V�;œخu�!��N������)�4�֒���}����͇G����{�}�gi
сZ���N�+��3[����n'�s�w�u��D<ן}��tIXS�^�^ѕ��u��++�������f�N�������{�Kwe�4l5�x�)��˼:��s���N�W<w�������o���9)�i����%Un�Լ`���x  ���=����3��e@�*�k߿�u �:5�c^��w�
A�H\ߟ�W�:s3���������U=]	��P��N��{���O
�J�^��w�����DG��}�p�f����4����0�+
����H,�Y++�9��'�S�~��[�.�5��u��SY-���Y���I '���g;)e!Z������ �"e�s��������z���]~�L�}�@@�;��,ߕ`�paL@@�q#z��$��shV��Q}sLR.x��2����YZ�|D�M�nuD�z����	R9� ��$���a�a��9�ҩE[��۶�H�5�����U����7��`�`r�ӽ�T>'Ʋ���=�1�q��پ$F�ڢ|I��bD^�ԓ%�	��� �eeQ��ƞ��ovLվ��I��� �bw��	�2�.�M.��A<#q�PgŻ� �A����|Pڽ��)�#����R��7���M�>�>��@y�\�}����'p��KuY�-��w�_d�Y��
����b�z�zmo�Uܑ�b���Ԃ5
���X�ɂ�z�;���o�g-�	O����NQk>�����_�3�L����v�{|S�Պ�!���g'�������v�]r}�ZK�"������9�f�:$��Ū�U����.,/��ŭ��yd�^�*�a����"PoH{�xo�ޗ׶��@-��wg}�X�Po�s+}�fP�i��ʺ��4���T�6�r��fC��d^�t{�jG����ъ]vI��}����W�>x�H�|����4��?(�X�o��F_��I�(b���|���P��n�]���{�����n�ѭ`"��״�
��}���@#ͯW��\Iҽ���N��������Ļ�o��j�	����rzG��g����H����J�� ��^�9-�:�\N�����=69{�8{��7�s�7;�7v�f���S_��Fo�Om��������'����-�Ѵ���j~�#�-~~�m7��A�Bya������9���茞׵���8����+lI4�E�3P'f`��AL��5��V\]����{/�Xp���-^��u���O� 8�n=�^S6^i����������E��{aY��A��
���4��,I�8kwۙ�r&l�(��k����ݍ��d����r���;�{������,6��
~aU�ե���ɑ��J
9j���+Z���2ҥk*%JDQ��1J�6��-(�Q�r���ŕ����+j�*�Eb�1e�UEUX��Z(�cq*(���꒢���j�QAUEc�,U�#�`���k�������EmEh,b��[����ڈ5*�K�F�̵բ�M��A2��LA2�2ʢ.5TjX,kʡ�L��r�UTc1�����U���UL�p�TB�-Z����".e0�)�EF2(��DdPL�TT	R̫%1�R�
��J6��+C����A���(�Z�ʊ��kE��YR�i��cAn�Ŋ�T�U�*UAJʪȪ��b�j"FҨ�mh�Q&P�)�X",U-J�A�Q�WQAX�[1�UH�#�h�X�
1X"��e�QX�QT�H�QEm(��TWT+�UE����ƣJ��c+mb��q��ji�iD�"*����+�0F1PX�����������յ�?D��^&b�2�j5��꺲K��LeTA�X�I"�o�������]q�ht�Q ��9� N�LD�B�������	6��k��ˣ|���iv7 N7�$��7�(�y�TG0Ne�˛��A!A^%CA��{nGO�vq�K].:��8ywF;t�֗b����~�����,^վ�؝��A8�z��b�^�ܐ�����7�(��u��H�d�P�k{*�IY5�&(��4�=�+��#;��I�ګy�d��{{���ܜI0Є�"��Օ�(���@�O�zЉ���۵/�#"s��$�guP$z���f""���LGVZ �����>'ǣ{��"�����L�GM�Z�*�W�5.m�ժ�5�L[[;f=��e��n�*�[�x��:�b&bI�ȝ��N�����:έ�U)+��L�� {}��ٕ^3�<SM��6a��׾��������'ٍV32p�GMe�Icw�Q��O���??�}����d�=�4�:��%F펻y�(�VCiEؐ4��t)�����~�/A͢������|O���M	�VȐr��wj��6v#�]WTH'�{������D�SUx��1'#�s5@�O����^ ��V� �Y��\��As�M����k�*�I&����D�3#A�w�Lm�ͷ5Ud��ު� ���$����"B!�B��VV{oygAB/�9��4H'�v��I�D�VJ��:��݌:	뺨�X��Ʌf""��$\OuU�e���Gn���� ��9O�'����bպ�9:n��O��D�7�S�[�t��=�#'c�t��bgFM�p���(ms�Ĝ��8�TE�U(��B��&��VO�� xzi�-�h�����H��tm�s�����i�#�(m퓮�=;[��wt[=X�w����<บ&���ϓ��ՎT��lm�'2�s5���.�x�db�sѱ��cs�VƓ,�0�=��`z�ܻ�s�rn0�Q곺��y7@�m��^Ӷ��=ѕ��EE�p/3R�n"����g�Oo<�K��n��Ύ��{U�]��A�.nGg�vy�<��GW8�A��B��v��u���n�M6ڄن�{�˪ڠI �V� ��Ot�;4mf�;�)�V��� �V�"j�6�0��LIu]�D�a٣�j7-C��rF�"�vD��O�'��������I��3Ñ�Ӄ��o $z2���L�t�u�f�fX$[8�A���Dm��40�j�wei�+��&���9�����A������3KM�d�ۮA��1	�,�Nh�<����M b9��D"B��	&�{��9�4c�U;��o�R��@�E�2XIÂb ���kn:��C�\n�>E=4��R�G��NY�ߟ����g<t3�� ��q;�(��|2;z����q���� A ��ݪ ����	�h�eCE����� ��S��LoG	�u�-Q[
T��`I�
,f]�3�]��o�ค{q�S��"��!=�C"��/7E�BR�s�N|����b��Ϊ$}���TIe'��Ĭ7%�:�K�!�BBi��U]�(�r;�h�O,[��76���E��M�FGoP����&�0�������/G�T��$�Tn�W���ơ������wake�pXMC�5ݔ(d��u�
ʎL�H9�4	"�u�;GXN�GN��Ԉ��ʼ��'\�r��7P�u^J��G�O&ӥ�9t�ܔL�x�d�b.";�J� �n�S�S������|Ed� ���һ�Su��o��$�wuW�D^�"0` ؄��s�A6����h����A>���I��rA:���	��:��$
���	�aCe6���=8 ���$��I��8t
�/��f,�7M��cek��^ٗ�=�z�	���ǹ�6maDB�@/m�M�G���>�ky;��W4�4=j32�p�&�Q#����O{;�I��@�A��rL�]n &�DC1 ����NI驛z$�R�$�O��H$�u	ΰ��NY4;o'*�L��H�E�1����rH!t�ɀEln�+��E���$�k���[=�G��&ל�^���j"B0��I�M]��v�t�v���<v�n�����4��u���Ͽ�ke�pXMC�M�eQ>$�� �A[=�@�/���#0ӛ�$�kg�"�R���؇S��稙�c\�qluC�
2g	�[; ���Ag�Spz;+�p��3��n

K{lI ��u
Ǣ�cw]�zs�F.Q	lz0 ��~��>��r`�^6�M��ۚ��7)�GM?O�gVMx���������Gil�+cr�`�i��w��v��iͬZ&\�w4�N}{�t����Ƹ�P��8������W}h�(��e��Nb3��Aa�yy?{�  ,|�w� �:z�B-�C1&�o�A���A1�NL�m)`�&-��E���G���Q�0�Y����U<R+��ٜ�9,�8��J�����M�Aqr̜f8"�I@c�����)0a����׎|	$��[TI9�!�9q1�<�����A$E�e
1���P(��j���'���s��s.�A"/+*�$��ު ��Ў���o-�!WJPu�"�
u@λ�|I׻�D�{����]�%F�E�I*��$�}�T	���FD�#��AIo��̺����4����H���@�H5s���rE��墤"vz��=�l8mۈmU��$�kg\�z�Ԛ�;t��D���ι�|N��U H�W<�baY���VoC�����x^�K���T�tHS|��)�KQ��6����P��s�7@���N��絇�s��x����}�i����n���r��x�Ȥ"X��p��|\$�	��]���l�T�2?����m�[�-��'ou�r/k��Xݰ��&-�6��\�mō�����)pm&�o<��9�	��]��%�$�]d�.����Xm�n$\v�F+)���87vz�M�;5�@�npl{l���^q�	��ny�v��:S�EV�I��ׇ�`��=����^&[�Ff�8a�����M"����5�[ڭ1�n�:'�Y�ӄ�Kxqc�<����Cb��ݱt���dځ����~��5�A~5�T@$}��(W\�I©R���z���$�ut��T��	���ֽ�^��d����g��{�z�@5u�H �]�3WE*��$�C�($aBa5D�fUH5��A$F��Lf�܎v8���^$�W\����m�lD:��2,M�YO{z"�iy�sD�	���%wV��Dq���i�жLNM���DǛ����O�_V��K��p��7TA�r�[=�F�g�ܫ��ZN(H�PKm�v���5m���64c�M�{��dg�5y{q������m���C��u�\�Яkk\��A!t��%^Xz$��bt���� ���$��\��0Y���)��]��t9剪D'D_E�4�҄.�N�g�����~�0��lu����F����<����F�.zC�|�պN/9!�� 7�>��2�H'ą���A�Mo�{wG�{I��+)3	�a��nݼ ���hQ�&��$Q�|��1c�����A˭r ��T>/�x&�8PE�e=�~�oz�T���Fc�I�*�2�Y�=H3��6Ğ�$��2��!�!��ݜ�$�����0����xOVT��Bʽ�'Čݞ� ���N��qR�mF�{m]m�g���ø����������z����'"	pQA�¯��y�PAF[���t�;g��sÐ:���o7ƹ���[���(��M�x瓟��`1[�0�8砐H%]fРs�zk��	wMҪ<��E�4�lO8(6&a0���Vl�  ���Q4�3qt�HȖ���Ψ���(B)��f�;��tR��F�E�ƕ����#ln�PMe�D��Z��a�d:���އ.Gx����sퟦ�1c�e&a�&n����\�V�/�����z�$�힯P9u�,nf��:�k׽]�(7,���!0��>��ʢI.��&��
ꁾ�٢���I9u�|Lf�yyв�$I�l���8���p2�A��d �um���/J:�:p����a�r:�?���w���tC�/vrh|wvzEH��� �TӅ�w�
��;g*�O�:z��xL�cͲ���gw3.z�od�Q$�͞��$�k+�cؗA8��廴F�+`��\2Þ�]8�k\�I;��j������^$j뜂&�s�2Zp�Ժw*%�̛�devt�>$@��� ���g����k{w&�
&�Y�j�]a�˳*�ڮk����C������}����z�;����Q�h$n�3Tp1{TF���J����|5PVRf�وu@�^9�>_ml�O!���`��.x�A��r �-�ڠ]�:9j!\h�Iح�m8콥{gӞ���f�;=�������ȧj��/g�S�>{�U�I�5��H%oV�=
4��0�*��`�Ml�Dg��D�%3�s̡DK�����rt�	��$�B9}KF�䉭��'��&CcͲ���I%_V�H�QY�K��p��W8�	wV� ME�+`��.a�k����hڛm^?�-ρ$��]T	'9�S��Z�x&oq� ͚�Bp�$�et�$�>飢^;��%Ipt��t�$�몁'5�M\OCo��<���W�������w)�Ǯ�,ҩ��<�b�U�H�q�ܣ�'�&�k;[t����^�d9A��p?u��jfb�M��5��4`�ydw�X����j�n�|JҔ�L��?�݅j�v�HJvA���v�{�[��8A�Z2t���	]+.n�[H�^�4���E���v���}n,���Ķ�g�G?u��K��̾/���rpW؉�!͗}�,��y!)>>�����D7��e���!�c�;��?x+E�	��xN��
���r��z����̈́ ���g�7Z{�v�zi4b{d�-�]e��F��b�9'/�CR� ���z�`�1�W��j�x�py]��{^C����wNܸ<.���l����q�>�33��y.�#w��/ZvǑ���'�v�cTw���4��o`��:yo���=����&��.�N���zE���wz-�ś1{ѻ������&�����}�2�|/���/��t�g�nҋ�jplɂ^��"ri�N���q'�����8�$PK>X-]���8(���3At �m<E��,5#��m�q�|��������<�7OR�՝�q*��h�gL�.�q�'c
�=���Ѽ�V�[�"���l��SN�?����l�d�/�=(�\����{��9��Ӱw����G��r���Ğ������a�����F�ӞN�tF2�ddtm��ȼ^Ku[�O��3j�\��{Q-���ف�ZtR[Z4��M��w�et����ޘq[���N����J�V��;�ħw�}% O��'��%EUc ���am"���`X��5JA�F"���Em�Q�*�A-�1DU`��ʢ���m�e��b(����Q�TQT�
$U�+�`��"*��"X���R"��+kb"*��ң"3I� �0Uc��
��E�)TQq��D��ek*+����cL`�*V(��&5�PqVDEb���ib�b�*1UIm�m�R���XZU��
��EkKV�(������b�R�b�UUT��&"uj���%aQEI�V��*,W�+mX*�`�����JZk�FW�)�*�@�DYe�q�eE�-eE�"։��ƣ+r�`士*�H娫Ī:� ��*�$ESVb+��E����L�Ҫ���jҌ�1Db��W-�j�%*,T��*:j�[L��Q�Q�����V\j���R� R��؊�"�"9h���%q�`��[1�LQAV��?���3m�[���[yg\�&�[n9#��5X�9�<��� �)ַp�f�<L��N�7
N�O]�,�O>�*�X8�=Z���{<�<�����[���kl&w!��μHk���'k���9v�E�g\���/��D�&���r6���gqt)Y\C[�ٮ�=�lZ�=e��+�v��m�����u-n;ry{jh��p���(�[�k�����g=���G�lqv9{����^�݌�ug�jV�oc�k��s�z�rn.�nn�d�ױsò���]�5<l;;��{]�Y4��� �6� *ql�㙑`�q�n./Y��n�Oj�;.�`7g��t���pqv�r�jN�6
��$����D�nL��\g�kg�K����U��\TOc�g�c[����v����O$Sz
we�Xh��*ᆁt�nm���6f7r��@zi͵�H�3�mv�E+���h{xt�:��v��:݆��l�v��;L�=��;���z\9�%q���өB�sǫ3��Z�GXxc��ѻ^]����u��z���ɹ7�N��Qh�ʁ�4mۦ������rsΧ�q�Ү���q�yP�u@�v!����J����b�Otv�6͓������
�Y����c�M��`�\;;���tr��`��3��;q��7o"\A��۴m���=�;J3��{=t{��͚��.��0m�D�5�Bn������u��u������ewm��X��<��*��_2�x{���۸�xu����OF��1�u����cp�';S���l]���F<[8w\HE��!fx��c�i{[gj�'�u��s{�3�;��c r>�S��ܻ�=�s��l��Þ2���C�=�[���3��u�=lO��nK��:���r!P�a�\炞wc�%>)�|�x��qJ�:Aon׶[Xlҵ�N4YK3�m�d���7Y&��;�t�Gv���LBt�l���7�ZL�p�Fj� ������7π�b��ce�9{A��7u�"Ep�RqA�ld�קl0��4���cnf�Pn�.����_4�1�S����Mպy�v�ك����c�	/j�L�e�l7N�cge:��j�n�̯�����իu�S�]��T�ۚ��>3�4Ol�,7uڦ��ku̜h��k1o�~
��
뵤uΙ�uێzҶ���d<v����=ڭPuk�3�7S���6�^_uݠ��$G�D�v�m���[OlU_������*�:��$��kj�$���}���Y:(̧$U�d�$��
�ba�__eQ]2�,�|�I+���Ă@�{�D+S%Dӗ"�G<$E�SHE6p"W��{�Gĝ׽4I'�sU�ɕv���_1��V��
�9�U�^!��1��AH0��j��oov�x��TH$�縪�x���g���l�^�� ,O5��k��A'nu�9�npW8$윜��@�{�@E���+��J ��rw�w����a( �(,a���;��<��ݧ�r�q��g�y��k��O�����9�I'1ǣ+��I��Mx�I>���k#��2�xdW]Q��Ux��#i �14��A�y-��0�u�U*��99�}�������J=���!G�A�"|�8������NW���Y�Z��hAE�D�-ڗ�:����}�_z� ��>��@��9���&g(l�c�ڌ����pT�r��*����9$�o��v+q֒�}�@�	 ��91�R���8k�;g&.#s*wz;E���� ���$��يɸ�&�OU琓�H�e���+��f��|bj�W�T	�w<�$���B餆\Mll���1���[��թ�7	;�V�(Lu�"�q ]�<%�D(pﻡF�"6{��x��r	!uv�S-�׹rr��ޝ�:����0 1!�LI���H���L���P7�[�4Is�I �-�ڢL��T�z��A/x�����&W�m���ջB�&u�g�!�Ud	��7d@�4�[w����ig#elE?OC�<�ހ�����ym���96d��F����P/n�i��{�{6���A ���|A�!u}�@�^�
�bE�__e[Ub�"��"���rO�>U]�@�@�{Ԑ���Y��|z��#���H&�C�5�U���O�Z�e���W���O�+v���Fkޡ������H��o�k:�Mk���ݷ����Cý�oX���zg�����0(�e�q�x�J�����g=꣊��	lT��9�A*�����Z��6�k��
ɋ7u�?Fl7���x�I]��(�3��Q>\�J���::��f�E�pˈbJ��	��dW��t� �I�{3�4�s�fG� gd�P1�j!ZK� 6I�5㛘�z��!��vt�$;vv��E_[�s�7���Տ�z�%忭�5�K��T��n8@fK���j��L�T�{�h�H|���UP=GY�P�*zv:��v�n��Dkb��|<��쩹�I�5��@1�ڇ/~̪�Mg���X��mQ��y�#wgdP$��\�[vY���]lQ�-]B��l��I�S�-s�`wbBC94s.�rȩ���]�9�G����� ��\xq�>A �����I5|�[[�UqZ5\�$B�� ����'ۏ!)�0T"�p��[���s��Zr�e�X���^��Q$����3p���25���r�v-r�8,0�l:�u}@N�VI�3�,�2�r H7�=4H$����L��P 8.��$���s̨;"�H+;6hH>��ω$l���"��Hw����Q
,���I�Tsr2Q$��Zpf���v�"�gP�E_EH@����2t0�V��qJ6ܗ�Uzsgq�����9�X�#�iA~����Ys-�FTV��N�7�wzL���<�>b���v�p��[;+���{� ��!C��H�z�i�:��q�[[��Lq�݆��b�un����}#���BƯnε�n$��kIZ7&�1�%��69�
�nwa��l�grk^{vN..�w��z��ў�(���u8�٬a����ɒޞ�x�10�1���<8�D����h�mvX����6��l��'4<]`0��w[��������j�D&��3�	6JC��MN��טA;=�;x6�N�:j3��-���xC��т����TI �lT��ْ���x�\չ9=8	VlT�di[�AC`�Gd^O����봜Pkjg	�W�"I ���3�|`q3�+��ۼ�"��%>�
�Y-����đs�2A9ھghT_>	�r$���3�E��(�DAa��a�k����hͰzÐ��tĒH����wrz���}j"��t<s�L�ȸP 80؈�$��L�z�vDMFʺ�}��9q����>���>�On�U K97Q��+�N1��8��&��4��K��;q.�����KuG�Xq&?<���Q�$C
&|�^9 ���ϤH���&��ͫȜ�2EӟA99�$�5�0�&��̪'�5�a��ɊQQ�Ĉgp�Z�B3[hc	�.����.�^[٧psV�no8�@Pܪv�7{�͉{��T�&kJ�pU�G�xx�u� �W]��>!n��� G8�Z�wV�[� Q5J
�i�Gg��h}�m2"#��B�{��9 ��m  �o��-��N�
�X-�%/9�x+��O�"�e�-� ��o�C�OJ=:��=�q�ǒA�]Q5��
(ȥT��C�s0 ������+�2���]�����69�v@�:�u�Am�=�3ñ����G���J�� 7=�(<����'S��\tm����h�����`'�b�Ns�M$M����I��+��'�}1�~���� G��7bw���+�(~0��1yP�IC��跆�̙�|� |�=�=5�E$�\��ɎȻ�t��,�T	�����o�@�_�� p���ܮΎ*�Y7�����+Utۋ������.oBݣ�mr�'��=0�"Z-�+��t�u,����}�/wk��L��;�W����߻���:/��d{"�H���0�7����a��%�	���-wk	&��H����^H�ݝU:��Ɇ���y��w_���4����T��g��A,��K8����eR��sz�!�>=�>dC@%��m��<挣����#�O1��#=�sq��9%�7:�ȝ�q�3����������~�͢���T>���0n\�r wkq'aE(���T�dDe�6�y�Ǧ`AUM&���� 	��u��e5/=x�""��p���m��ql��z
:�M	ި�Q^h��O$�o�s2 ��]��I��B�៽��~�� ���q���6�Q;�L�P��4�i	�굓�RMN���l��]��>�s���S뼥<�f�?xy����=�������h��Z�.�g{'��x{*'�uO�{�w{&L5��z�O=�l�6��a�� �2O�W�k�I���b*JI�cGVy�"߿[L�mFŏ���z�~̷��l ���m2"wv`}�w�b<`6�%�>Q�0=.�6��G]��u�:��WN�"�9:���~��ƌWj*����S����i�|kz톹3�E�O��ǫ��D0�fݰ>���ń 6K6�6��N��xE*����" =�Ͱ��m2��%뾯h��=S
�I���ͤ��ev�L> '��^���R\�eǀ�9���𶷛a~�%��D��1T�n[3{�s^9�-"z�&�)$�I{�$ג^U}n�%���cۺ�פ�陜I�;!2ABCZ���U
H$Mg[�J���l��e�D����Y]��dDC�ʷ�k�g���u%���H�0��&r�A�{����
�EH�Z'�lJ1BgE��As��z���-�s������ݟ��(/�3>����m�XXA��=������i�v ]�R��g���f��=�o=�u���01�+���N����N�я"�;@�/hGE�����2L���@{v��w�v����#�N}�P�l�\�q�.�]��.w����w���z�ӷ=����s�s ;{U���ݒ���YS�pl��&�\����,ҹ�Ǘ/�`��v훭�>�N��hˬ�n�q��c�q��,������Y�>]��ϱZ䦘ICpY����L@%CA�x��q��B��[`�e�h:��ꚭ�x�^"�&����@|.��p��蛘D��	�٨����B�1G��&muu�{�>=��� !�z�D0� ӣnofr��ZHky�!�Xp�f�y��� {��ȃ��O�L��T�������>~Ϋ`9��Ϫ`A5P��M�}��ވ:&g�.ʋH�S˙4%z��h�A%���T]97��^ ��L+�鉗�d��i6��4����U����t9j��(�x��>�l A��v�3�^�o����[��n��;v�ndɳ���9���O�����sҘw���?����n���
�|.��p�)���D��v��E].�{�W�6� @���'ejl@& 0��t�c��I)�/��[��kt�
�4�s�qMܬw1�LT,5���xܾ����w>��<�դ=����pe�k�ʓ�\.���< ���{&��]�=��`�)�j�/}?uQ4�wi���s;�HnM�(��a4ኊJry�&�Y=�B�) �ҕ=�E��������C@�{��%nSI�ن��&���}yy)�����4� ��]��=ꥮ�����%���:��zg*`PL��T��~`�!u{m�L;j��9�W �`ռ�)�f�;�;����+��t\ƪ�]d��w^��/=Kp��%5�=�l���b@lU_Ͽ��_܆���4���ޫ��{��L> �o;i�{x������I#��m }������4��R���C�.��i2#��UD�̟>�� _���/m�U"��N_Y3a�fw��6v��o��JeLf׼�L �m��D ҸQ4�{hX�Q�+u�u����x$ΰSV���#%8� {;]����{r�%���zor�Ƚaf��s��n��Sܷ�wp��o$��v�ܺg%��9/���e�r%���G�	���9i�t~U'�Mλ��%��>�ԣ�'���yi�w�c�� ��^T�z�)���޾v-c���Y�eI�3�(	�O�K��mr�l�lP�tW^��徐�8���
o��`qG�ďj��ۥ�;���c�L���Q2wC����y��f���~c7S�^��(6vرv�� ��t���X���n-o��6s#I���#��ћ<��Q��iJ�b��>z=/xu��~!��*daA�n��Q��6'r�lz������Qϫ�<����Cz�{ӻdp]@�h���(-;��ly���0��Ҁm	�;e�G3u/?x�����N�_<�,�-G��B�A�>Y2ۣ����	?	��sKF*����P���`�ϻ�6uk8�)�YX��x�1	�2.��F�ï3�8�*�|ŜJ��f(0
�ֈ��o��ݨ��}Y�8�)8b��o��Zź�w�W7wC���g�����K~�kߩ�U�&>X�g��3�G�JE����^�t��M�6�o��s�}�{���GN��`���pŽu3�eޥ^�e'�V��r坐Xw�6Y�����nBgIf2�3c܎��r"[ɚ������S�����޺��_�ޯf�XL�����6<�̼�ya�U2"�"��b�(�`%���
"�؈���,X��2,�cQQV$TE���PR �ЬbYX"
[QE�����Y��īm�,�V"6���U�F҈,���bQF�\j���*-�	l��Ȫ�1e��X",U�*,D�(�PV*(��IU�Vֶj��AS)X���B��j��1Qc(�,���խ�Mi�Vb�eEX�+*�iA[eVګPTUMP�AQ�[lEij�*�ȉY*)m��#)-�DV(��IX[J�Z�,PX�5��ҥ@�1�)5J��EU�Qk]Z*�j�*ȳV�4�E��TQ��e��T�(�l��lR�ł5�E`�ֈ���Z����E����$uj,+1E��
�`ą�]Ye�"�(T`�*6�AdX��*6�I~�N����D~~����H/m�o��Y6AJ��*�_�����UVl<����`� Gm부 ��N�:9󦸳�t�s��H9ܪ����1�PR�*��D6\nsj� ��M1wz�L[�Y��0����d �y��W�1�wL嚈4�&b ��^v���mѯe��nwV!�.ۯjM�S�߼��v�Wg�m� ���v |��nT;&#���ell�o5�@ ��zݕ�%��x_�<�M~�BI�ͼ���tO;��Հ z9���o:�D4�g��i�ڮ�}�u{�4��R���C�l_�� ��[Y[����]�o� ����̈���V�6��o���@P�Rޜ���.�0�"��d�A%��I���˱���x��?��.� �o�=�棢��g���u�3@ӽ8���=��SK��z��MܣY�.��v,��ve�{��'�*sj�I��\��0�HBlR`���L A����<���d�!�c��"�u\D03{�3>A�Ӿk��������]������ե6Q4��n�v�)���'/[���������������B"�F��٭�""-��� ��ٙ�pm�R��V]�\k��$ה��	!C�qF���"�Hc����b[2'������������i�ݙ�@��g�I�j�y�wА���L8!CA,��I����n0 �ٝ{xc�˄c��@ �u6�ٽٙ���ނk��C���Tn����F�ل�A���`����fb���ۻ��q�h�I�|��ɿB$�E����#�'m�����ly���ۇ�	۽�����ۓ��*���=U8%[��dک�����n���L^�*�vf���s����n[���\��yV�b����x	�eD2�Cl7=��|t�nk�O[�:+u��n��N,��gt���%ǔ��ö{W];v�!#���qqѹ�m\9�n�J�P��z���8{kZ�����]�.;��kh�n<v<��.뎂y�
˺����Y����g�택\����f��А���K�W$��t1�lm��5���_]z���W<2��cY0��v�o���z|,\�
v�i۳v��\�.�m�<��ul�ß/v��޶�'�?���}�B&)�_%;:��K�foe]�Ps��y6�잻��uq�v��0���D��
(�D6�y<܀\t{陙m׷��0����f ��{5��o�����e='h_H�L!
!���PT����I,����I7�,�i�緼y��`�8��� �;�ّ�9��r��	�L(��M&�ٮ�._�z���_c� >@.}Zƒ$uc���Nvx�$�>��&�;�UD�2W�;h�l���@��6Fv��&�����.�����޽�� {�u���|���6�j�S*�~Ȇ=�j�m�Kb�1R8���	�8����O�Y3��&��@p��;�oŒ!���+�]�]tqGnN�R }금]�^ǉ�{��{�1 7si���1W�IU�5J��:�z�JZ�gK�P}>U���c��}�A���Fj��.���f���ƿo|l�4l{����<���������}Y����` >�fۆ �ͦ�@�t��LC�$e�׸��uy4�"�-�|d��� ���s$\���*�ٞ� �i�C}z�^�/����lU){}u��=]y��aIC�긆�
��\0>;_fi����:�����Sh��@� �@���{/��D��y�F�NY�#i�O��K��Ʉ����٘����5=�s���2�$�[0��6���z���m^ct<v8�F�!iz�r�ngpM�)4`��:�*���H$��ש/$M��UXJ��V�'�;y=���}X�K��l&�C�A�cF��3>��6�[�ίL��\��H �J���4 7_fDDj����W�On)V���ISU0)��4�t� {��� )�θ���*�{�-�]#��ɲybg��.)5���%��oov�N�P�D@15&��͓�d�Ƥ[��<ہ�Z�0[�F^e� �v'� LeR�� ��y_:�(%m}TM��*v�K�E�؃E�GK{��/	�����\�
I"V��]�a#9ѳМ�H���&���uIW�pBe��\mu`�I3�5�	`C�ɯES��� ���p� onvf&s�f��]DAd�\��P���5lvHq�����s�huk��˙*���+p��+��K搂T0�P�|���@R$��{` �cg���B�?L�o�]I����w���xf
M���͘��	$e�Yw{*�W���u�D��{��F �N����p[p��ϊut������� �D�\�m���S  *��TWC�Vod��{Ѩnwe�6K�s�j�$5�T'ɸn�I�f�����Gy;�_���p�'�]�I �^�$�8� �#/m��U�2��;</`\n%6؁�F�ɞ@�yP�����)�7�>�=طW#���т�ī������M�Q��i&���|�'�I���.ɽ�S�l�jb?GNz	$�V��zB{>�y�g�P��dFWt�� W?90��t�Kg��x��� �4[ �Y�na���zfcvz���>�c�ŷf�������!�l&���ۗF�^I���z>*��p�go���<�Է��dF 
ޝnC���@�"��D�m��� Ή��ugQ��z�>����4�W?Sa�IO�cՋ/�o|�]�Og|I�y˅��/
)���{O]� ��Qi ڙ6�&�:�s���"wg[�\�M���U�RSP�����S�/1�H�ޝ��+U�@ ���g���~�#c����Dj:�������MMT�J&�?��Λ {���*Զ���v��Y[_W���Z�N"gs��H'�:�+��Η���۸�@خO=\^�v[�����Ck"����w�y�����b��p&&�/mY��M�v#�0�fdB�����aB��	l��>,��!�8�ŕ��]��� �>ݻ��x�C�u�s��.ylo5������ƃrYMz���1˵q��9x5D�m6K��!v�[>z:�lvz�S<��1��ֶ��4ۇ&Y�����؃�i��v�;<���R���ٻu;wYޭ�q�ֲeú����M<i|8;g��p:x�j����w�i]��wU�n5�Rm�7��&Ž��h��<���ϗ��6Q��~���R@�]SQ0��[����nSL _�ogf`}3\���'���nH�Y�M��ig.6�8�آ��U	%S�W�=djY�3{9��q/'��~�+�S��sd����lQ9[/$'w���$�s�q�<޶�N� �oe7�f�y��ӎ
f
L(P��g<�j2��u�L���D�M0� ��y�@ ��N���|�Nj�ĐNn�W�P�����d�N�.�ͻ�H��5�G7�o���.h��@+��p���7�"�ӭ��s��/:9�GDy"�D�}	6XQ�����s*�l/6���d�5s��`L�??��~���g�,��[\�G��� ��ukG^�yپv�D;~��f�cqQoSm�10�3�MtuT"j{`�x�����N۳kΡ~\N���;&��S���~�F|���6�}�Gm>��<jAl�=�&�{[��r�����[�u~I� ?w~��+�;T!Eʈ(��w�qgj(6ET�M&˭�f, ����H ���G�kɳ�wc���30+�;"&^��A��<o�O���m�M�9���l�y��7
� ��uz���7�Pd$��u�ߒ�bl��I��n��k�6����q��e�2/�ܣ٘�/����
�η$ I�c�JXcs�:;iB� ��A$[r�����n��q�#錺�v;pnŷe��q[9�[���u���d�O	ݫ��D�$�f�		 ����
�b:�tF��oD�t�rixj�&���Q1N�/��;�O����=Z�ٜ� vֱ��Iy>�tI��sf���7�VH/^e��n����%DT�L6�}<�`y�6�/U�.6�����3�T���wnI��7��-w6��sU����:�%�Y&!� �wU�\VE���EU�"r�t͈wW꛻���D�:��A�E~~� ���4
Z���^R����l�$C�o����rDD�����@gwfdS�W�yDEe�J;#*�*��S� ��6$���%��ZQ7tV>�����
���?�@�i�����oǲ7~}��ߑ�[���F��^]�q�C�j��cci��.''Nx��.��~��v�]��Q�Q.��|�� �i� ������$��[�a��H@�I/���IRk٩}_LR�U,h��nf �m=�5��ӷ� |ʳ�n���ui�nb�^�]M�u�K�B|ۆ�DM8h/_������� ��e�<��#�ʽX?o�g� 
��l @��v]�Hh��Pہ	��`љ���!wg*Y�w��E���l���wy� z�u����3a��'m�̄z�^mb[p�f�<����^N�b]��]�ܽ1��5Ŷ	�gz�*;�q.[�+n^�����y�tۙh�dwc?$��c�I
����z��M6�]�ى` ogm��#Y��],x��}n;��n#��[��Dݷ�mhdf� �(2��E���Y�q�+������͜m�[�6�[MW�߿��g�ʯ�����Gww�` ���լb!��݋�:��$����@��q�X0 �0˦w*.pBI%Ի
��S�p{�9�W��f` $z�u�$-k�']y��nڐRc٨���
B����{q�$ z�v܀Dn��Ew���"7�n��1���mHm/�*�UEDM8a|�|�T�.���@]��@ +v��"�ӗk�� �6l$�ξ˲o�&��6�Bm�a��~�1H�t��~�G;�F����[��+vu��Ӎ�+���������N���g�5Րj�),r��:f'oN�ƌ�+(�N޳╒�j�[��Q���<9��������+,s�0n\���.���Jr�IW`��f�zcbws��q�77ro���qoD^݉{��e�����D5���n[��y}��_vo�����m3v����*l�01M�Z^Я����5�7�g��Y����n
E�)����^���6���g��w6���w��P�r�٬��Ƀ�sWü���{� z�N�y�?E���,Y��K�g_r�y\�a�����C�S	;�t�n8�
f�U~a0aم�3>~��-���H���ȑ}�8�	���?h��8�y��N���'-_J77�ns�<�l�7�m����{`��A���FzC��z��\ץP{ݼ/A���~՝��GY���C ���ziu>v_zF�b��v��z.����ɷS�)3������<��.ڠ�̰���n����w�Ak�ו����/�d�o�b+��9�;sE���'e�i�1�X���[�JC�|�����6ܯ���0���.X��D��76&�^�W*œ<�wөi���i��,^�6��p:�;<�9�7 y��矜�n�!��yQ�O圼<�S�ޢ��,x����ݿ���A~��ƫUL��_WHޞ����>ܞ2�}i�,ʼ���o��I�8g=�1|���G��qx�6���\ ��8V{;_�g��������'HO�j�:g��t	<Ew�{�{�0�H�UWo�#��*��w��<��o#�i����vA��M>�g�Td�Ҵ�(���kF,X(�"�1EPE*1AE"�����4�D�F,QV

��4�D�[`X�b5���QEX����*��mR�Q�6��YQUE��T���e�����P4�EAUrю4m*DV
���X�-EX�,Y-���"�AU���UAR*ʘ�"�]%U�X�\�c*��*TZ�DĹj1��M3dLe&��,�U��Zʣ
�UYm
Ec�c1X*�(����,EPD�CIX���dX(��-J�sc1��E���X��X�*fX
�+b���ժ���EX,EDU��k,PEQdPUP]!Rڥq0DU�Qb�
((j���%��
i	QdX�I��V����T,Ms�6�53��Z�x;�g�g�t����H�r$u�b�c�k==��A�+��M��U/oP���溴�ۮ�Wx
�r�=s{x�٤x.��A�g�{s�n�g�m�;r�N��l�2���4;;���I����v�Us�n󻶋���z6当���T�vv�] )nؚ윙6�t)My�����]c�����!d�5�;7I�����t{&Gj�?���d:_Z���9L ҳ�8�7lb���J��v��i�p��9��m��\�]�׋.�C���'�v�ojB/Bmm���òt��V��C]��#]���\���,-�۶�M�^��ln�d��#�7ջv2�;h���Jg���mZ2�`͑q�A��#��U^��w'y�]j�ru�c�^ɮƗ�LA�[�-�K��A�"���Rώ4V;��z��Ŏ���l݀ε�2�-�\7n�ӭ�\���-���k<��1��[�XB�x�9-��&;,{\�u�/g�t��lsuچ���ʿ�������۸�n���zh�q�e�m˫%ƺj����*@�b�U��qy�I����w<>����Ŭ��G��3�#�u�=r4���K��>^��m��;vݼ��=|�8N��%a�mrn-՞W�+ی�6vv��a��-�9���[x�n܆�o(l�$��`w�v�Ժ\V�1٩��l�=Z�.ʒ�l�n����l�5m]��(�l��Q۰Ȝ�kr)p�r�3��v����<�ݝ;vy i��+��'�GSkb�\ƹ��)2{z�u���]�ն�kq�j�{^���:�M�ɻb'.��z��E��픻�3:����ys��ͳǶ�����B�v��AO:��*{;��pGnU�vP��t�9��&��z��sp�q�k���|��f�Ŭg�g\��Km��lɮ��n�� x�q\��l8�V�:/�X�Ʊ6�2�uٲb��������V�㝱]��ҝp����|���C�$[�ڼa�*�Ӯ���x;f�8����Ge������\��q�܆u�h�X1VM�oOVJ3�s��㛷;'Y7�ں�Ѳ�J�^�����V�ۈ:ܣr���ً�t�{8��M�3��s�1�v�=�Ƿ;�<p�������C�<�=��cf��s�m�\��\ۻ[��t�cJ�sn�9�z��UѶ�L�]!��7��M�s��:��r�OS���O����!���^�`�[�x*�ܻ�I$�ceh$���$޷z����ٞo� "�gm�'������R���M�)3"�o�ޝ��{��57�E��~�@ +�����w��RZ7���T�ժ��s�;��d���U�4�6� ]��0> �W���Q�y�Ҭ��$�I<[��^O�.��[KZ��BL@j�yofm�����j�ś�� n��0�D�c@ ���n�=�iפݚ�&��TO�x,�A��+pBw�VDI�߬��.�W��僘���lP��$�g�ww�0<�b�gOL�(����:�����\>-՜v����f��[��È�ʆލ�=�M�\2��Y�A��+�8܈ ���y�{gc�*�/nb �����g�T�D���
V�C��f,�td+���լ�i��=G�s���4ǀ�|c�w�o�zO
'f�D�w������\�5c]@1I���wZ�L?���k�~i$�H=ה����*�'lu�/+si],�r���K�*
��U&�{6[N@��ݕb�$�곦�[قI���*�䐾�˻	�
1��#	Cĺq^S}���d�KGP�I/$�w��N5�W���K~�*	%?+"'��̰�$Bp`5J���۱iy"rz6hB�K:fH\�nZY[nM$����vI6OF�WW7��[��9e�(aP�%0Љխ�u^�v<�n5�
t󇓔�q;�!�c��[1����m�P
zIy8�
D��;���  �}ZȂ	=��7�Vu6�"_~��v{6h�m$d��bC'��!B�Bq�bI~y��$����� WF�B),Q'F�ދ}M�8��l �QU']���� �7m��#�}����a8����ha�,��2��o�,H���St]�A���婆/{��t��c��=���Ԙ�,�l�eX�6bf�5J#��S�g��I{���� ����@���.b�"�Q_ERm�]9rdV�HD]�y�� �w\PI$��R�qd��-����)�I:+_��N/�PPG	�\4{��N�+�)�6�b��5����g�,���""3��{[V@|���-�+��[����~���O�J�x��[�h�I��\B�ku��X:�a�Ųk�gs�?�����4kn̄Qg����`|Aq۶Ց 
��h%�j]�}������q���ҍ��M�a@)Ѡ��[�) �Qx߫ރ7��` ��ۮ�� /�ӈ4�5�A�������ĴT���D�"f���.;9�D4��` b~���7ך��@ �qۭ�|��C�k�Sh�a�)��N�Y<9��eWQ�Y���VD/��p��{�f>��.F���q���e����{�$����Oo#�Ա1gz�Og���A�{�%��q _j�'���	\w��wi8�^#ڻv�w�6j ~,wY �W�\��B�[Ieι4��[���XV����"���]D4/�`IW�]w~KN�P�m]��.��*�J����� �Z��mL	������yr��K�r�^�<�z	��0��G���J�����"RH^mu�$����U�Pg��QI%7\��Rw\6�$�e"�#�ە�+#m{}����7�nȃ���p� ,�>���-w�V��^.+a����}^ݸE4�$ApL'}ȳ�~&�_<X �h�늉���ݕ��_u�$�H^u�݄�\���D$��h�������W���H���""n�f` ;u��v�|�W�:nI͌�뺛����B��UAI������ 8��b�tW]��	��\D4Y����> |n��{<�o7^���K:[��� Z,��}�1�i�]v�4��q����9���3u�^:��8�1ׇ�q�j�ţl���*��������^��Z�L;]u̗U�E�|��]uOV�Nɹv�<Q�><���A�-�B��������3�r���u�6p��1��ǎW�|N�nu�]s�[����g&[�t��:rϘ|��"=n�5�\x�z��`�V��{�}�����i�qۍWm�e�ۄN�H1�x���4lOl#�8�R�J�������]�T�����u���zm��^aQ�S�k����;��x��4���5�csɧ�6W:��~�������#����__��ג's�ʣi ^��ڂy�����z��t�!�3�����=�����I1St�3|�����*oǯޭL� ���dF ���j�&%��A��n��' �'9�e!&a�}��������4 \(��=��؎�?>�Ā@-��f` ���P-�֪E%��"�0�~��ŏ�Y�~��  �N����{��r���$�Nw����>l�ZkLL[��3�T  �nSL�٢�ݡ>��j{o33>�㵿����N#�&0p�X���\!�Se �b�R�n[VRs�g� *�x�q{h5�������'aAUT������H ~;na� ��[�;=m��T�
��~�π zn��/�{'�"�2�g��B�w4�X#��$_O�[ ��F㐢鎶�����vvB�#b����k%C�$�Gf�ju��N(��kX�*NM�u��^�*�J�>m��'����$_{)�@��y�Ӝ������x�8�	@pB�K)nU4�D�m�$�C5߰o���I�X�j��I)�D�)9�(Ґ�$T�6�5��L���FѝmQ$��e�h 3������X�n���Fю�J�T�J
A$U�Az�M��{�07c{�k�O�TA�%�9�X��t�"!����1e��	{��~.?�r����uR[&��]dC�{��g����:���� �3��~���"\����|�@�]6�Y��f`FB��?
]���* @|_k��o� ��LU*�컴���<�:�ڥy~J��_y���>�o{3� 5<�o(���''�F�y�+�*�B���Rl=��q����	 �~Y99�*�]��EE��[]=he(���j�4��S��(}�һ�xf�2w6�m���V�2�#+w��19DT�5I�Q7	mo�Z�w��*Ff��[Ǿ�5�w�{�b;�{��>g������@ ����.��=0�{c��x�ٕq�K7�٘ �����T[^���'0���&#��E�'"��_{s�Ƕ��I���Q��ʸ�h;{9� !��=�=@�_�������ώ+���&�e.�\�H��3'n���@��>%-΄Σ��~�?[Y ����{\Ȁ=���Db��\��}�S��Mb��tI�����oE̝��Bi��Y�S˲�4�[�k+/#b�6/���g~��>��� ^�������dEm�~&t�t�a�R��B�TRo��gf,��{nb!����s���ۜ��G���o �v��>�\4��(����Sa�ܧ�7�Ȭi�Ul�>�>y� v똆�k��qv�E	�#l��3���y�vv��DM�vb��ĝ��윥��[F�f���W�ǣ���p��	��d�����F�١vO$�+r��A��L\D��3P�e��s ���i���o�2�nv��@|7kj���a.#"�_\ENn�-$`ˆ`�'�nޮ���xv�z�J�F�{;pm�v�3�[��|��w��*e
��S�#_v�@|���>�n(6�i�i�MV[�f �;��C�^X�E��I����s�I=�Y�[����|� �d���m9$�]7|ya��Eu���	h�g��*j*f&j*-���o� �~�M0@J옾E�����/}���ڢs����b�JR��i^vy��׿ �l}n��	�;q�<��'���GJ�*�N�iP+��i�P"bJU���ަ�����kh{��I�/�D1�:m $��?~��lg=�k�,�l����q�����L��������[��1���'nI�K�����.�3�ְ�Ww�i��z��f/fȝt��0��ui��X�Qj�Gh�qG58��j;�ś�26�:�;t<��v��s�뺽��y�Wvns��'cЂgr�Mٓ��SaƦL]i�wV���ݮ����ۂ�ܘ�&��54;c=3�C�S�_+w/\Ho��Į7cl'�-�l�1�y�s:�n݆��c�x�c���:��jνOמ@㳗ڨ���ϋ1���[��l�-��ɲ�\�͂�x�8�r���m+����{7=��9(�"Ҍ�w���
�e ���U�U��� �>��7#�����cm_L�	݊���6b0Y��?��{�>X�[�p�����@ 6�@����A�k���Y�����$]534I34��7" ����#\GD[�T��> 3�RDA$��{�p��3ɰ�0�E8�q�콉��{��yC��@ �s��@ ;ϻ2#;m�?v�sU����/��9����bP)B�TR�n>˻I$�b͚�T��4Z��\�YD�lf��a�{����{[T=�[� ����̑����H`�!D@A ��!n����v�s\&����l���~�?1���c�RX���0�\����` w�m�
�M�1x���˪h��kz���2OdD�&a5 �L��� tW��P����zl����e�,T���]0��ʺo���<�ďb4ȗ[�m��e�v�_#�˞X��/�4x���w�^��՞��*���>�����h�%�us)m)ua�2v2l�`�6?��{�0#�n����>��EOf��a��2��.��� .׽�� �}�<����E�p ��!�o�8�Q�~n8�[�dC��NT�-ד���I'U}wi/p�#�.�C,�x.����I5�ΩZ�;:xm�D���� o�u���>}Ww�D����m�˞�]Q�w5nn۵�S\��m�J-���\- Yp�@���sܷ���1\�ng� |���R |�����O�ג��׻٘� ;�:ڐ��TAACN
W�˾rk�[W=i�e[~s�o��"��dC@�Sk���L�ilQ��3�]�n_�^2Mh1f"�h:e��N!���ڸ _c�=���o\��߅�NYH�\��������r��%M
�v��X6�� ���,�
P=�
�&�U�>�����T;˅�ӦL��� Rm�����t�`ڽ��+;yF�a97;���,��!��H�I7w���5�w�/wy(�����zreNm��wR������!#�i���;�u�Q;9o�{y�s��n/Lw���ܞ�Ʉ^=�t�k(n�S�W�a��v�]��ɹ#tͫ�i�5(�',�"݇���$Eݺ�ڲ��oc1�uo�o�j;�{�����/�'8qPi��Mɍ���]���M�M����C���)Pd�]:��_��v�G�#�6��պ�Խ��<�o��on�8\˨
���s���{����.u�_r�˞�'M4yt�83۴���I�=}j��W����Db���<
O����K��D��.ǹ�f-궐׳Q�����^G��
v�u�:�=�/�ıۃ��L�l��>�>�ƕ�c�l�9���f��/]T�o���ؤ���hW&�|�c��	�P��z�ʏ{p��%�9�T��.�5J���{��`�w�w ﯒��z�{���@X�8WP��ٵ�_�n���s�QtW��u~k��lN�_�	�OA��U>w�+Ц�e�u����p`���{f�+cT�n�z'�)ݯi��U^������ws�&W�s��˓N��w��k�AO���}�e�m+\�z������V5{R���(+`�4��"^>�
׽���U��ǚ�{<�M�9�<��S`���XȌ��3�ATPQB�ePDYib0²,� ��QTdZ�Kb�R#�[j((bDb�V�%`��cUեaYA`�ī��h)"+2ʪ����`�PQZш��8¡�`��eB�+��.��Ņk�WJ�H&����C(T��Ҥ����$r��E������2mfeLk1������Z�d1��Z��%d�D1���+q�D$�AT\j8[��u�X���P]e�SIP�+QH��PF
�ڰU��rB��,��
,2�J�VH�P�Df8�c*"�e��T�&��B���2�����|祴���AgS`Qq�مU�Qh���f�[a0b�I%�<����p����f���J��O}��o���<Pb���D"�	�nS`[���+{|���7��3��}n�|+s��>z�����k�}�O���9���8�D���ۋ=����q�5�vv=X�������8��W��?uf�J55ſm6��u6D /W��3�/<Wn�x��F��6� >E{:�@^�# �Pl4�W���]K�H���^ǹ��ux�  >���4�W��1�Um���g�<�վ^�ꀁD�ҁ6̝nb���� 'a���#;Pt���Iy"��&�"�C2w��� d��`\B$�l���ݼt�Na9��w���]η"�w�z�Mgc�<�2� ї�L�RDΩ5��oE��=�u�UPk�����03�,��ݕoR7��S�˹r�'���&�5�ySQv��"��6�����U�E
*le�s0 �m[H*��*k���ٮ��Nl� {��3  �v�\�0q�0�T��2��U��X����3��A�<d�Ӝf$�Ja�c��i��a�j�����ި^I�v��� �3�m��o����w���$Dg��f��{Q5�d&jjgS`���x�*}�u�Y��n�̈�>:��B@j�7�t�s�T��8g�P��RT��ٹ��İD{�ڸ�Ax�ꍸ���<� %����H��ӄ����� �L&��"���':\ݟ{�V ^�cq� >�{m�C!��Wu��e�9{�%����ܻ&�< ����mf�÷�9>$ '�^�v݉w��>��X��f`Dy�6>��Gz��Wb���{B	�N��4�������fuîyD�������ԟWĭ,ϙ�φ���e�>[;}M�16���s���l�a40�Ʈ�\��-�OR����u���E�]�W�d:�ɹyy��F_^O pkt
�ݭ��۞�	�q���/dwe꺻�L�C��6�<U���V�^�[g�K�$v��G��>l]2�b�_�v�wW��<[c�pq�x���w
��=x����hϷ�9Wv��t��{[�<�<��ݎ��cuOm�m3�m��xlݙ�l���f�N�]s�cWc�쉣ѧm��ۊ��y4�x��s�?j��Æ�8-D�'W�w�K�/%ٷV�� _>u�?�R���L�����I�G��{0��hRm�BI��ʅ��.��t�̥w�N몏�[��p��9�jH������d�Vg�e�&�}��M�$�����r ��:�s�.�Zܛ�_�sy�"o�)��>s���\�L�)A�[AN�]�<3o���w�p�6�D�ڶ��c ;{���饞v��u��8oup	�A�`�Xl���`y���Ȁ�;���E��"x}y�w��0��6۽����dZ⪞ښ�2�1AD4�A(�4��"��q�ۣGYp�ֺ��.L����أxj����97�ESUDN�$y����z��� �޻�K9�8 �y��+���$I3����%E�J�U5D���:�|�`|=�!��nK��;�owB_�
�-d�sg*�i��=��<k����:�N�g�ʙ��Q���".K)`F�1q��u�o���� �H/ݕp����̈���g2��
n����.h��n
S3W���L �3w9���"9�j�\ݠ�q� �E�r�DD{u�d�юt����� ��]g=�[q%e4��&k��&�Iz��$�m���9�}��>��k��9]3 �UR*Sh珳0�g��mN78�:�=Û@fw��_ �[����#;q�./T_YIřT8-�F<��6�۞�{)s��5��mն�uq�+jc>�K*��������TUU [��_�~}�0��n"#x�yË5�ӈ��	g��f֯���"����M�={�l ��G�g�.������� ���m $⢹����rot��0�6�����8-D�����D���ےI��)�s<b%D
S;M���=ۢ���ac���}��=�w������������|R��K��v�{s�;swX�^��DW�{3 @|_nS`}�LmDL�D���a/�׆���Ē]��w�n[��"��Z�귒G�]�m��%�&"NJf���8�A�_�U���=14�1˲���� �}M��"������dTg-��b���y���We��x�(�^��^��]�d˺�E�Km~���b#��x%��<��S��I$����$���oQ9�������i���@�ȩ&�b&i@���m\4�'f�ލ���ow�����m�C��]6��F�9�w^=_��tF3q!�-0V��w��	}����[��{L���DDx{\�M)�D�)�n	�bM6TSg_�q76u�a��πA��U� ��n���w[�B����fU�i�پ�5��5m�?kS}���+pMZ�f:�r��{�@��v��ohѲ�6�.뺞ӽ0s�ANn�&��B5L"N	�ﶹ���Ӹ����;���w�w*�#P�o�� �{��<��W�`��Ƞ�@��c��I4�e'8��얁y�2.{��L���8g�>����A5U���7� ����dA�����%�C!ۆ�d���u��I!�7�꼑�r��!Yn�4��e�$vL�3|�⪷!��_ �>^yۇ�D����6�=�˭�އ2�*I�R��	�}�i0�";w��� �Y=V�*Z=��q� }ή""+���wa$!�(���pʊ�n�Ϳjuc���p*P�=���!�=��vM�$��]h�TܵP�aԗ�v�J���bp�)˥�]�F�H �{V��-�]�}�㴦����n �����/���#_�<����;Z>wU<��Oi�xGN�M��jeȅ7�w#c�b,�M�ޓ�n'���L'�z���!a~�O�ʜ#et��|n{Mw���p,����P化M�h����rι�+�չ)]��PO��x�{�Ns�լ�9�[�ۙ�8�^}�pS��-�RŌjN����Ӱ��v��Љ��`�u�k�(�;���w@�6�e�c3e�;u��O;�'`W͝����A�v';����@ɯ��z�� �֬�+����۞���]Cp�p����[^).�1�l6�cf�:�5ˤ�]��vK�=pX��G��4��1�#<�??�{~s��+Ӳ5���?�`�A���ϰ���qw�W�ُ',��Sh �{ٙ�Yw�����P�4_m���;[3o�h�[�� ���fb��{V�"=�k�]n!>|I��� "Yn�<V��1` _�մ��1=;Qw�F�V�����f  E��l�Ƣ�LBp (a!D�����i ��� ^ۈ��E��]O��,�+r���2HV�mݤ��'"m8`�����@$��G����yy=j�3;��D��l ��`��N]����M{�i �a7� 	�4R<=<�e�����wgs���۰ױ���k������f�]SUY\���f` >ٵm� /���#c.zf9��o� �6�@%�[H��`$\ ?�]��>Ϯ�z�݉��S�4')v@�N��5�B
��@s&jvN���$�r�R�<���/o�zbۻV�-�uCwǆ�����x�+^y޾� ���}�V�)'y�Ӡ�zr�� K��ƌ@-�5U�}���/��  �ld�c�}}��z�� ��r�@"|?CV, 0�Ʋ鿥cPJ�r����^k� �@+�e�` �w;3���?ɳD��G��ل��Ôl�E�C	
''��$�]�}T\1���c"�/�i �/=�m	۹ِ[�}�����'.`TcPX!�H�%�\c�;P�3u�����<)v7l�ɠ�������dUU3Q2ަ� ��6 ���]�#�`���g��ؒL�#5�氓��X"�Z��^��<a�zek��VS��� �e\D0;w;3�Q%]Ue3�Ʋ������&����
��*ᠽ~��G�s�,"��mƶꇅם�yכ��7���_9�}T���l;�-��ܳ�~�<L��S�td
�*q<�+�'�ơ��Qo�Dr ��N"�}��٘�=�X���P�5J{q��]=\�>�t��ڸa,����}�O���K��v���h,wn��$��)t�Zb�6�|�1` �ڶ�O���7�{�Ѷ�ê�����o>A|_f��[�rL��[Y�����R��?v������ܫ��ɇIZ������xݳ�UW��_�\�14�g$��q�����+�m�	��f�Lc�Ne[ ^����,P�"D����2�כM���Q���_�rk{;k� @.�������ڶ� �'YoJ�Q޺z�R_tU"j��UT���w^��� /�j� ��	��ĩ���[{ ۝��ٮBO��G�K	H0J �Z�"���w�.�"7޶�r����p� �s���K�!�\�����q�P�y����4[�v�.B�h���`�37��y����=#| ��W�YKJ�h�Ǔ<r�Dhd#:kd�	/Cλ�Kh��,D��	*�e���C@�k�YYSlI�>�oݳ}wa"L��"�INtrF��f�)�O�	 ,b�Cƃ+U�랃���k �t&�m�Nۖ\��;u�q�r�Ͼ߿��@ e�Y۶~� ���a'	?�':��y-��7}u�s}�vD�"�:�@<\74J���4�6��\D'�.Ϳ�UN��0D��ကD�S�H�%;s����w��2a0�Y�L�)����ͦ�H"/�[�� Nk��Mn��:����8@)��T�%)�RLE��xSgm$����rIY�<��K� ]w�� 9��� �=��P����T^_�=���#j���%���B �~���W��~�[]t��f[��!��6 ;+z��\�b�]n8�������Φ�ŪХ�)��5�4gbŽ����eLC�?�P=Dͦf�cG�O>�v5�Q�.n.�]�Z��	��Q���`�>oG�T�.O��}�d����e������J׽�ջye�˸IV�����t%�vڳ7�0-�T,�q-V��l����P�B���u��C�:j��ۺ�}��'�d��P�.fo��խ�Hg�u��ns�w�R�!��%B��.�cz�{e��~a��}�k�)�K����Y��=U��ȟ�Ď͊]��f2 n
��٤�.n[�Bn5�p{w�/��^�7G�`����2#���t���,;������R��n�g�����6X�+�N]Þ?n�OC`cTKxjأ���8N�ZE��؈{9�/ga�s���Ӓ�J����nޝ��t�уսQ����7VisB�}Q���a�g[�+wFv��=�&�u�b��3��$�,�zP�d�5���$�2�){"����p-n��Ǿh���޾^�{u�0h���@=ݘi)�u�1���j^�{�^2`:��e���J��a��p
�M9ͥ����a��uݵ�V�̗�@��fj�@'h�t���{;�@�g����Bޔ�c�Vp�%�pn�|g��;��½�$�w}�/D�Wj�UC�ps'R��-^�8�B�2rg����2�M��{��r��y�3y�����~}�o��=���C�֮1������2���p{i{�i�E
�=�l�:��5wE��I�ߑ�����T(�E��($1��1�d0aYX,+����A]2���(Ȣ*tɉ�E\IX�ZU"Ȳ�P��-�([j@PQ`e�TAV�b�@XV���Z��(�SL1ӧ2��X�5�	Y\J����UT4�Qi*#V�-d.P+1�cJX(J T��U�i4�IuE��I&8��- �
����*�T�c+��X�.\�k,&���[ee�aY����`�5�H�����"�E��µ�:��4UZʕ����EBVLˎaQ�0��T�e�eT!YY*DSY��\�a��ki��Ȗ���������b�N&[*6�F��(���q�;p{??�������ōv�̤^|�μ���uu���-;0[V�%vf�qn�>���ն�ݭ��sv�S��:��v��vr� z��!,{v�\�p���@�Бv2�s�=�'<�74�\��[Ac��Vح�mmSX��M��q�Zt�݈7^,�t�g����ݲ��q�-�&�f�UmgK\#� �[�{wh3ǵva�Ѹ�س�շ�3�ۦ�m�c�ZN��sWJ������F%��Z��uP� ��v-7�k�����]M��ш�����c���
��S�d���M!pW/����&�ӊ��ۘ���ڇ�w3�ǁ���Om��b-������Ӛk�8�Z!�cN7\�nq�닅L6�Wl�c�eɉ�Z.{]��c�W3[�x�/.�4��<';f�ܽ]�j�����#v78�8�W=s�fj�`r�TQ���]8� �u����.�sq+	�m&Pr��Qs��4v���876N�	��n�]Y��mF0�tQ�q���⮓���\����U�7��7�#������j�;pk[h���-���#n2!�[ӻ�r<�n�ڃt[{�nJ��r����e7��)ϲ�Ώ�/��غ�n0#���`��sm�u����\ʼЧ=�8��V�nK<����l�t��mں�;qv7[h�9K��q�u!��C
#cBtn�u�a��n5��n�,qs��۵n7R���3������v�qjmr\N�ݹ}�P��u�˻zh��`�W,'�[���]pǄ�{G3��wj��Hø�!fws�M[����\�ú�����N��6��^[87n�gw1��4�Ν��0�a/=]`9��[��\����%�9�+���c�;YxC�6�����c/Iή�6��u�/Y��^�ڷ/v��������t��E,&���d�nf�`=��T��b۶k��W][�^v�hŮ��'�nn*��ZvC'7�N͉��*7<rd��1ְs�P�P;�V���4��u�՘�h5֞����<�&��^��lH��7.�n5J��������5j��=���=h�k��d�ִ�Vz�8�]�����=vbbY�xPp����lkpv��z�Vݗ^��Uu�{��RX�7=�1�H8ݗ{z;� �������ٻ7s����^���b��`�Y��q�]6��Ƞ�\6:�j��=����h�G;�
F�;v6H�6p��a����mٷ5_�w���R�TP%Q��羧��t�  ]罙�w��m*'�U_{4�ݦ�@�H}�M���~&H�QJ�6S��q��!7>��zaê�@C�u`I��{�w��NEG솠=5���74J�D�3Ha�ަ��y�� �Z�����i�q���V�|��05�D��j�P�'ەu&?^�^��@ �ܫ��@oV�ݤJ\�5G�,�fI]�:&��;�2a��8��t��r�֗�A.{�i*�ԭ�8o��΍��Osf�$J��vM�y�9��G��;2s�c�l����'[�=�m�	���燷d��&G@�Jj�ƣȄPo���=�m� {Ϲ��� ���[��٨�b�\B���$���'`��,D�I(M�=5�y$Ñt��6�s�LNz-��o��Ԩ=�3�a潿A�F���o=����k�}ڴA�����
d�}bRn��po�b���MMp����ڝZy��q�/����f` [�o��lTFG��x{/���C�5�HJ�(�R�M�s�� ��[ �y0��ۘt$�I�%�q�@}�8�!U4����	�z�(��Kyw��{�?x n�7������� }�O�N�F��Q- ���@+5�Dza5R�v�+;�� ���6S[����芩��@};o�1 �#�ަ�@nS�����r���]�������c���B^�+q]�k�G[��v�8Sbw�Lk�\R�}�����e�����o� :��m  >ܫ�����-=�����]�v%ys�uI-p-F�A[@�\	��\��M/Z3���+����`  �k}n@ ۔�B�S����;{<�3�$5��A���D�Ch�N!��?nSI� '_M�`���'������Ǫ}#Y~��٣�7ꙇ�O��=�^v�}�68(Fu��A�}�����8��w���`B^Y���8Sګ�D�ϱ���nS�c�9�$��JU)�S��Z��]�c@{����>'�;p� [�ݘ���e�݈�M{)�8���Al()�	
����k�wu�]�ʡ�W��+�}5yn !���� 7��wimӫ��]�%@PB0���8vom/)}r�b�8�e�
�G=�7������~v��!TTQ��j����� �oeU�xT�e�yowobo�'�Ή4����M�$��)D� ���UN�����D�g�F���V���O�v���.���3������Eku��ڳ����KM"�p �+�	�$}����p�#���b���`=�V�A�o���F-qF⩉(�$�G=�6���	��i�� ��u?� >.��fb�y�̒�u*m���I;]!~2^�٦���䟩�e��+�,SY'4���uE�����EK6,=��gs�rn��<�w��x'P��L�Ӟ$x�aB\
1=��� y���V�/�C�2��h";{�� 9��h��us;�Xϰ��nz��s�D�Nu�ݵ.���S��=V:�e �p����?-�DL��)�/��t�| ~��<� ��m���}�j4���h @ww{3 �Er�'�3���ЈJn�%��� 2	�� �{٘�A�vڒ��Q
$/�]}�(o�2�&0��%��ώ���` �N��A �G2��_R�3�pDf�y���'[�[r��TTASR4��O��ٯU��f��$��Ё0��~�H��4�K�B�}�s0����$����o㙾mQ�˳�==��פ���6�{[� �7���8��,�p{ �2��PF�T>��L޸і+Ibci����#dE�s�I)���E\���S�_n�̉�o^1��Jn��F&//."���o�ߟ?�X���9�RK���ۋ����(��	�d[�؛�9{=�Oe�/|�c��f�Of�\n�7Z�s�s�P
��s�ݭ�|��l9ݻE�s���g	Spst�W���qGi]`z�է.U뇎1���X��X��`�C�ι�jo6�C��S���Ws��+��g�-�W�m2�����)ҏG�pt�:��pukv����^^��NS�t����rqAr�U�ۮޮz�k{Z�s��T�;2q���.�Bqs�l5bz�a���oϼ�1�~
+6��NR�iy$ I�����FD��j�S���ĀH��6�<㌇2�T�U �=�?���զ����� �\$��ȹD�i�|���k��ow��8�RyMT*��h�����q� ��F7�{��q� > �~�c �"~��"���x�8RxR��`]՛yu��U1�U�$�SsM���ǌh �oy���]h~^���fk����*�d4`���w�+"8H����9�����{>���-�}���H;���s荞׮v�T��#yM�+8���CGw`��m�ɹ�{uA�Np)�G��h"� ��f�]����8�8�r >����<�sٛ�c}�o��9�h?t�r|?����g�*bSh����` ���3����3�������^͹��t�K�!��!#�}�}<kio��5y{{e'���zN��sq��#u:�uY���W)���| 	�� -���"""	�:#Oh]��|�� �:#��H�K$&�����;���g���J�t������8��@�o{3 �3���h�lG��%�g}Fy�;� ]^�$@����� �f��Ww_)\iG���H�9���=4AR���2�����z-�S�rk�a�x*��E�I̺�a�����H"��|ڣ�Z�Mϧ��=����(�,k�)�OOsnb��sμS�}��&Z���Q�~�?��z�]0|ߡy��?�A�oy��>_N��@?�f��ȿ�wKmI�oo{3 �Ob�&�� ��q\=�PL����~�s���'1�w������7DS/U��s�Ol����D�o�N�-�ͅ=��X"/��ڠH�o=3ڧ]ئ.�������cG�(!ՋO���ߊ��.�e��a���E�@���3�s��������Ϯ;g�$Ɣ�^az���þ ;w���E�Lf��h@�-[ef�}V}��4�ʚ :���b ���r�D���N/A������>�f�3)9DǾ&�P��z�����Ki�q~�uf_V͸� ��f`D��TA䗔�EUBQ���k�[=�\DA���h&�}�����ܽ�N����s�;��c��n^�/;gf�*T̔�QY|w_�3 ��ͷD@����ir騩�:�S���9�٘� ���A�ܧ2���&��&�?��O��&��_��ǳ����o�>��s��	�[r@����w�5�u���~-��,�Rl���j���^�9"*b}��)[�Χ� ���@�F>�����
	�T�LJo�K�̛l�VA�hZӘ��z�u��~�c��{�"�}7YІ����ksGr�U�;�v�)����)���d��/����2�6q㣚�GF�K�6��pbK�g=��-�D�Y�A��H��@Ғ*���n���� ;����_���z�q��H���r� ����ovY+�����f�`Q�0Փ\ǱcO`����k@11�ι6��������f;�i5��=�TD�Ki9 %����(�=��E�iQ G���RI�;4B*Q3JDS����C�u�Of绽^�����,}M��{�0 ��mJ��L�w�A�)����&�R�i����s|��<�M�W-���|� ���RA�o��0��ѥ+[I�&�Q�/�ܲnb=����ݰ>۞n@w��1 |f�����q�؈�]l�rE�x(ah4h;��AIi�lgߤ���5��[�cA,��fg�|/���H3��p��Lv�4��P�Yqn���D��U�"_�M�&V�lϳ�z;�7���}�[�Q,�I><��v�OD=�4ѺQ���2��%p8�'H&6�K���\)���˨��v燛��x�:�^չ�m��Ve�8�1j�m>!�L<>�x�6ʨn֝7n�sD�r�`ָ�-�s�*���q�.ۯK��kz!��N͎���E���\=���uę'�J%Gh7�g,�4�r��<�fd�gO>s՗/ϲ=l�\��;.Ͳ�v�û��Ŵ����6.VώI������c�8wZ�����UmV������56�o�AГ* ��b�-ˌ��I-��y��6� X_��b�,ߋ�N���{{�ϾD�G�1�iDMC�z����W35QK�/���O���]�ݙ� �/�����z��G�g}��o9{>�1I�=T�D�)N�7�ݘ���6� =Ǯ��C{ӫ��7����wvdF �5�@�ܨs!��l���0)�kcMf��a ����>X �{5�C���{��vK�,�q%~��w|I���d�� MUCe�o��Ȉ�{-���e��wI�ʃ�?{31 �E�g6�� ���%��K��(nΤ!I*H���e�5�Ϩs��3\Z^�ۘ�;��Gܽf��?;}��S)B�&���X |�j� �f쿃��^o�Jy���@ ����i7;���XI�O �]b�*Sb�}���=�����
2��G��,�v��Q>;�^���&����~���e���/]y����8�~�^������ ���D0}-� Jz�X�juR�u���!�
��Bj ��g��@ ��v?�A�y{��sfdH�}�"�[V@�����)#ojA(��;h�vy��;�S�� ��m�a�	?K����ova}Wޣ�V�:�H�~�՛b�1ʪI�U*	�����?��	���wSJk"{G���O���:` ����!�����]��\�Ud[1����ı'lRc���[<�E�p+��R�8��v�m��f����ڗ���d�(4
m�~â���'� 糍Ȁ���ݙ�Ei{Y�茒��n�5������
`�
R�H���q�y�b��g���Āc��D0;�ݙ� l��8�����Y��EL����M+h7r|܀ ������tמ}y\e>���ޠ�җu�hf�_y{��{y�ڠg<|�H���o���<_�AJtӽ�p���Ǯoww��3}s3UN7��f�m�9dJ��������O2Xj35W<^8`��輼�d�M��w:��qGM�G�^�4zNY!>(�m���gP��fEH��FL�(F��g���t��[��/@F��;'x0����_r�xӻ&&�Jǽ�X�ާ���f#�9�����KXi���27&)�5>~��wxSnwڥM�;�:B�vn,�>~�;�o�
]���5,w.�O�#�h�c
�(懱���a�i�*�?)�Q��q6�r�7��Ѻ4�'uE�Zj����q�wZ�&���:�Ȕť��S��s��i�u�%��a��V���6�ּ<���Q�WNiň���n��IH)uݜ�s�-g�F���4:�����ة�ے�v�CТ&�eV���#r�=NO�s>��M�ƻ�v��@��q |U��[b]�]�� �T���܅j��Pǋv&�V�c��]b�[�&	��)�Ԙ��9�]ӓ�]-�W-����=��q��;Q6;�̹��Fo�AU�^#e��3�n��!����{T'=����u+�`���@Y=8O9�9��۽;TK�!2]Z=�z���_N����i�/�\/�^�{��.�����w�s��o��yM�8�>3}�犗�g��(������X���w����������wZ��7"�3����ڒT�i7��v�/nIdAm|{�z#���=��G�|��F�YR��%�[X��X�D������-���B����Z�F���(�Vi�E�U+--d[���I�kR��,Pm��ȥ�%�B���VKJQr�1F(�Z�-l*F5�X�
��B�إk%R��X�(�m�B�J�����R�((,km�e��Ub�*-J�
�(E�m����
�b�V)-(�TM0�[C�d�M%�ɕ��T�-BȪ�PMP�ZVQFAA�&&&*,YXV����T�m
��1J�keJ�J������j�T*B��)UYUR��d*,�Jʕ��PR�%U-�ԉ"���FV�+JX5(�Um�ư��m-jZ�[D�+#JV���)*��[A���dc��*Q�jT*�B�Y(��.7V��J#mT�F���ny������� �c�ADD��� �.�Xx͝�!*k֠4��O4�@ �wsq�G3}s
���fvVwd��4@.ˌ�B��B"	�d��ߑ�~�� s7��TIS�t�a����-�V�!���ݙ�|��6�͑�쮈-�m��T�&Yl���0o!�[�;Og�)m��{!ۡ9�h�z�y����߳����SMlp[���@����9�9��O_vR�W���dDC�w��0���u4J������m�mPh�/��vVEE���c�ڄI�owfb�f�� ��	��y��}5� 4�ݡA��)M���������a�#s��R�R��g� ����GC�[Vy?�Z���f�ji[k�)�~�\�9qK'���=��D��C yӏۓU;ӹ3�<m���<c���ӑ��2�j�W�P�a�����s����9�[�׬��J����|�>xјοvH�F�9ƞIMe���$�{�AP颣����@|�8ܨ�y�F��<|���f` #������� ��H�ʳ���5]�~ޔ�pn�L/u\Vψˊy��wB"/<ݓ�1s��6�0_kE�!��s<��]�I �����!�NX�������fل��=c<���a� ������H"�5M�2�o{[�>����  ��9u(1\͗>��om�:n��R��	����o���g��=0�6h���h�ڲ�t�jA8;�(>��
R�o{6>�*�;�q{��Aѷ�Ղ ���a,����a�5s��{;+���l/`�h�)4�y���VD~���X?]D�J��=����Y��O�}��D03��3H�6�oz����gB�K�\cd���}��t�eܔ�G�N�}7�ۚsO�l1��y��/��M1�z,a��T����k;>���Hl�`Dc��l�7�������3e���N���=�
�&�u�v�ۂ6:�;��x���v�EuKݹ끷,m�M�\-t�W6[�����r��Zv�9�=����r����W�:Lv�ټLz�������@ۜV�J�͝ח������;p���蹋�{ս���.6mm�D58����g"; �r�-I���3���a���g��\��n���Z�g�y}��k�(�Z�����6O�)DT�W|T{�ڰ��iȀ@f�nf %�d2��sGG�΢ {Ӎ�:� C`��M-�ݻ��*cr���yOk�~�߬ ��2!���n���O�.�N�9�v,�4ԡW���� 3��y��A��^�dPHe��wSH�ΜnH>f�u݀��H�S��	�٪��V*����۷]{-�]l� ��ّ v�_O�x�NZ4X���v�"&Q]�$��& MyS��Z%%�/e���������N\F�{M� ���vf ��^�*K,qr��@����DG�E���z�ws������m�����fI��[Y�7��Y#x�C
���銡P�I%�wmQ&�\���2X-l��Y��������۲l<�<�%��`�l��aK�������1A��.�omK5��j�ǻ�/���vi�ي�(���«o�����E�٭�KXiΕ��S� �wkx���A�B��NH�bw�8{k@��T�DT���� |��3��� Vɽ�q*�WS�;�>��s3�Fw�=1a�����8&'�M_���n���7�D	x��L"��-߻_��5�:�dDR{~��@-�GL�*eB)D�T6�:7�n� ���j-^Ju��4�u߉?����ğ�'љ�� :[ruO���r�����;�壞���{Onk<,,��ܻ�n��}���{\]�1s=vA����ߏ퓱ͩ�}��o��G�3��`y���=8��Ӫ��y��Ā������T�*Pت�Y�*�Nk��`�x�5��"#a��0�󥶤�b�����rf���U��0p+�0Vz& S�T{5� ���������9�<��>�ǎzB�nN^�76z��t�7\}�{�Eq^<�oO5�8�g��{�94X�؉m���4\v�3��^�|�y�Q<�l�-�)L������w�gY��G�IQu�R�D��M��o�����*QQQ�͉y��0����O�qa�^�aN 7|��	��� t�/ 򻇷�X��1 ��ʑ@�;7:�~��5g7: D�0v�i���TN��Ӽ�:�t�9�l�b\�OOta<�@Ê��b9�� �0�<�ې�s6�
$�ٹ�@�����Y��g/�h@�v5���UEm�P$s�Y�4^#.ŵ@$M�U
ws��7X�b�&C�n&ٶH�|������>��w_H�	 �Y�qoak���uP�ww:h5�
�P�z& Ux���ȷ�pȽ���F��D�y��Dx�e����瘜cQ��-lNt�)�7P7�;q��Qǚw�Λ&���+#!�J�Ƈ�c ǧ�݅@���j�#2���Pޔ���	��r��O���s��jo���յT9ݝT ��k �u�������ι����#j}���GX쩳<�r�F,=e�D�hG9�P�L�l���Κ�3YO���]B��*�$�nu
�9b"X)���ِx�܆A��ЙXo��N{u=�A$��Ϊ�k$0L�D���r�L␣2g�\��-%
4Tף����5�$��ޕg��x	$^�uQ ���S��A(*!��󦕮�:�c)�޻���I"�V��7�S;r�9Ŷ,��=�D�8 �,�`��A���$��UQ��v��u�Z�}(I����C�_E�u��s`ns�uV�312𭍖v��8�I3f��{,E�k�pI���:1%X�4��DT�oq�ٌz�ƪa�y·_mg�@��&
��h���b!���sq�N8�]YWJ���F����n�5,SZ�-"mzZz{6�>멐n������������k[ûnHw�^6^����q��Xݬnh:I'=/v7#K����E-��ݗ8�܍-��bˊ�O,g\��N'����w΀��~i"X�y�t\k5�en�\[����.U�Wk��s�ݱ�n�bj�=K��FG$2�x ��lӌY�rrBl����n@��^�i���������"P�A7�r���5�>`�&���<�te����ܡ^$f��228��h8�"����&��d��Py O�}�ͱ��w���u��D����gTv�e8��Y=S�H�;b"X!8��6�5Y!�L�mר�L�+UD���{'M^gN�O�6k�X ����.�r�a�TD4�0�g��^$�ؾ]��>'���]z�7w:����ֆC�Uq\���&�̍�t	P�0߯��Q$��t׌@<��-V`���	$M�]P�;7:���Ք8t�̖"y�A�#	DL���פ�v�v�-����nݭlZ^cv4,�z����%�[6��0w�C ���GĂ@���
C�X؝ҍdϟ��.h�{aJ�(j0��ܪ ��*�P�u�������֢ן�D�ڗw��Mb�z��^�\2\���5�Eu�]��1�@���.��B���%����.3a͘��ω��۪�;7:�q�u��5�G�v�c;J"�؅#���4���H�w��7�f;V{ ��z@ �����T,ĵ��Zh����U���p�pt����g�v�I nvuW�$�Kv�D�Q^�ݓ �h�%���� ɘ���O���d����1
��b�c�� �nt�#�e�j�c���B��"YnE��6v�&�ݲ�ū��A4�+T�	J���������|o��0a��5}5T|O��gH�:VZT��\�Μ4������H��`�,!*�c�'����S��.���#�s�� Ҳ���:�J'b{n��G:�%C�.}�[�DҲ�A�l��	�һ&�)#�u8��:��Ӗ��E�J�FA�v�,���B�eS����wP֣"3p�X/U佭YU2�����@Oi�P��� 7��$' ��j���R�'��l�� I ���I'�}�S�jVC}�zz'Y"g��WAك�"�q �,�I�Ϊ	]����q��v��ޡ���ڊ}�y�������� �Fn���]�S�b�^n65�El۳�.���%�l��kR^�!�Z~ųޙ 8�j������vܫ�mk�O�5["O�t��D�7����G�d����A����oĂ��S�H'�{�U�|M��D;]��]�g
V+f�4c�$M��z� �Z��Q\�5T��I'�Z��@>��UP'��T�D �7sݹ��s�ݠ��iP� �+�A>&z��^�h�Ż����}ba�2�T����~��U]~���m��}ݪy�i������.��q��}�&7��h��L�J�]^��^.3u�yUچ��S������ê����|o/zh�psw����2�$O�GJ�A"n���ު.�1:-����[��a��ur��ɲ!��goG+�n�͆��q�L�?����׷bh%6�T�W|I�Ϊ@'��^�{;xwH��������H����)���1�
m����MoU=���X�%���q��}=�U@��ޑ@��9=[�梬"όX��D��7����z� �_t���܌������O$5�UD�{�(d�F�%c,��*�eƅ]�dXMi �:�I޽�H�Q�<����[�n͓ ��A%���@;�����>�FH[ٗ
c�N�2f�|O��?y�(�湟���$��H@��$ I?�H@�P$�	'�$ I?�	!I��B����$��$ I?���$��	!I� IO@�$�	!I�	!I� IO�H@��B��@�$����$�@IN�$ I?�1AY&SY��& ��_�rY��=�ݐ?���`s_>��U 

�HAI�wt((��PH�x}J�PT�UJQ)AC��/�����JE�q�G���gH��r%J�����R��Q�ԑJǽ�T��z��BR�Ӿ/���� -ۇ�AC�7B�T�� ���J����E��gW��y��W�$@s�EwB��FAJũ*9s�;��IC6HI=��P)x�V��B��T�+�z��ŪW�T\��D�    '�)T0CF ���LE?F*�M4� &F   F&�i��R52$	�0C 0a	��*�4�J4hdd�4  � z@�)�       � �#@�)�Sjz�S�hl)����t�v��[�nj����%B�������~�E����O��g�~T��P�#�1�� j�@(���@.��D0:|sU����||'N����C�l�k�cwIQ������4Q	��+ߏ�#�rل�E��
2�N��E�J���;X�/"2
.��lɦ)�+Ts�,۞)����h��/Ԣ�ٜ4\�1q�0�j�&U�X7wRN�b���v�c��Aj�m=�!æD����ۭsoQ��&<ɹ6X��LE��jE�jE��"�%�t�wy��CY��i��v�e�M^���<A\62�;ub���sQDd����l4 ��"=��Ģ��!Zo.���=�X#M�-!��f�(Mz�9��]^�u7d�10�`_[cֆmݸT�2�D��5�0v��1�m��/R��o(�ŖmfeP.a������%<�q�.���R���mV�d�b4�����b�qz�M�9V���1:Y��TVm9t�����`�-�l�2�2�4�ɛ�����2��P�	1Z�j��N��oU79ⰼ���Sa4mم,��/fX��9*+�����H�"��;X���e	r�Я"wA;L'u{�m]l��D�z\yi�V��ɘ����Y6/ؼ���i^�8�P��2=�>ya�g-���X�� �t��osTך��n�6�}�<� ��Ӷ���lmSo��Ϯ����[GF ����Bc��[R�m�֖e��WD�VX\#��LeM;򭈂���&�����
�,zD�J-Jz�T�YÕn:���X(�ע՛lm ӹ��N��wS@!��٩A]fL۫[-�]�{)5Y�
�4e�P��57kN4�@�n�����7$G6�Zc�h������Y�eV�Y��aJ�W��8�0�ItU(��(֖�+l��ڛt�wV`�S���"�72�
��e��x��Ո%�Qf�c5Q]h�E}���� o	VJ���S3d	�8�iF���ɡ2���`o%�	袍d�I���l�tnnW���t5G&v'n�J�Rf�̍2����RE�d�e;�@��n���j�`�kQEcni�+*2]`*
#b��ɕ�[��Pu�����W̳�M�
MV�]��$�+F���cE1L
z�+4lnعl�2�.F-��9�LL����I��46��f��yn�̺D�l�7(	�rGdIx�
�)�(���K1�P���'�Y{�
�o"h,�w��$����v���*��xF��u3Ԗ���u%[��p��	UQ̐�ڧ2�e�J���t*@��Pu��T��ޔ6�,���N����t�W)��	�-FM�i�@@���U�D^�����ڱS2���ݢ��3�t��{I�X�ԛ�h<sɗ�/Um�5,�U0ݵ.d4P.����$�,�rj��߫`�r��[�0Sԥ�+f�(k��3Csr������h�����e�L܇��\F+�G�'rMc�T�(-U���8!��F�࿴>g���z�k�aG)6�H2�GG"�:P@OtD*
�"�P�H*� �H���P@��
H���2"�Q�*��	"�� ��U*�ޏg�A�xvW������@kt�ض�D�md@�&���� ���2:��Y�~4�&��Z�Yt�~W/�0���&��@���^!N��|0T1��vX�Yj�쩭p/d��I��V�9*dY���G�ܩ����Yr���r���.ˮ�X&�@HMe���S���q��|�Һ��%��g@��2n�K�eţ>٤]�|�3s����G���{ZX�bB�`4��m�����'me�dmf��.�s��ܠo�:�Ck�]>�^&©|M�Т��6�Q�X����a�uc��C� ��E ��m�g\ͧ�;!{�_vv�嶋z@�0;,>v�g#���m�[��nt�q��U���A�u�E7I�V3�o\=8C҅�[�0٠�.����/������V��VN�.�:�̳�5J%�Y�5����=�咙�u3wLw�ZeX,l��IV�F�g��_����ؖ�"[}b�A���sl	1%!e�	!{⤃W2!�f�v�}J�d�ƺ]g�h[/7࠴V���O�J��&$l)o�����@�v��o,�AV.����+�͡�þ!�,Ӵ��n-��Ή�N��:u�9��s0e����]+���S>廈���1H�:�k^V�Ӕ_IgMTo"tv4��]w��Q��MH�[��3Tuz�UN�sTl:^kɅ��`�g��T�dCFͭy;�kq�-	��Εϲ�`������/��L["�يQ��,�nZt`������jY�Y*��DμY�<��r�rOD8����T�GC��E��Od�u-�����K�1J��̣�@��Ȝ��OF�q���Q��%f6knf�u���z�`��܄B(�/d�{���yY��V�T+��]�4;�]��^��D>Cy�8i�K���7ER�Wֹ�\����<��JQ�^dM�ʠ�r�I���R�x�!m]��EJfJ�3�KuS.��ʘ����'��V԰Z�bۍ��Bj×]�'��2��-�Pk|����xtY��q�눊�:t͊��W.�e�����I;fra�*.��Z��U��Pw�i�eX�DټҨ/{�\�R��I���*�'X��Sӣ6���m��ݺ#fu1k5�k�{'u�Rl��jTw�[q�6iK�s`"��x�B�*MR��*F�Պrw]@d��I:κ9��?�KF�p9����޽���x����50\�,�t�Ķ�F����n�g3Yk=��u�sm�]BH"l�;ʬuح(�c�;1���]��N]�����9���R��a�����-r��ւ��h�4��H���,�}�u�����e��ʎ���-��O(]ˢ��`��_[�����z�&�������S>��@LRjۼX�<�`�ט��@�b������]�9����m|�li~CЈH�}h]�gK���=�����OZ���vAkf֮ni6A��(�7jVV6ֺT���W(jqrkD���U�]�a�0����Bf��.��Q���¨]�/Ufзa�kU�l��Λ$Y���q�*��]��x�-H��5b]H�͈ʔe%.�n3u\�P�ю7l��k��n��U���eXT�bf!���]�Ў���T6`�jf�L �biU
�]90����;Ut"��hF�ɲ��]��k�2�T5f�rkdrV&3��,��ōOg��F�����J�u�H�)TҺ��:���
,F��;��֗L@�8���WhL��]5�+��8�+5e���Ar�f��ԡ�9ucc��f�>V�խ�.g��9�����u�X���[v_Mr�m��,yܢ1.��h��{Kl۞�]��r�X�ìDT���s�i����غ���N�>]�	���;N+.�I��낎7g�ηf�gX��[(�������R�L���.�[u�9���E�������m�M�;Q�"�JG$�Z�CM�,��B�cn�L�%��V��c��A��q��0� ۨ�l4(("K��n�.r�Y�{Tx3�#�m����7B�e���*��6�*AҍH��n�G.�WX�<hCd�����5��vT�0ڣe(Xh�fl�*�km�]4]v�+������K\v;I�oܧKA����n�c��\p,l�֗��Y���)e`�&��fm.�)�:�; s������/8�[Z{c��9�۵�V�4�n���*4#�n�fĸio4��J�R���h3;�&�Ѝs���-����$�ٖg���kW����o6�];\�����V܃���UR�u����F�틷Is$&�a��#,��M�T�m�:��g�����/+�7E�kA(������1�̻�e��X�B��.���Ռ0�1kM���$*�������,r�:��Z�M�^��9�;[�6t�tblv��[�3��
��ݭ�L�\�==�3������b �Y���$Jv��� ;@�u��u$�N��h�ph@��r'Dש^z%��������}s�^�{�߱�|�gʵ��4���nɮ([�1b��舵�sv��g ���V9���t�7+��n��֩mS��J�X%�T��s�x ���>�����<]n�zN�ԉl��vL�-ǖ��ϖ���rlζ�kz��Z���)uF�fn����:8`{��li[��-x����9�-�j]�w/m�3�y|�3�h�+�a=���=r��],��qq%�(�uu	� ���
)tu�W%׮f��w�?s���j�1 %�$����ދNA�����[�ߧ<֑"^��F,_�XU{�b�q���
��s���ku�T��L,��1R�[d�"�wf� �!��T�yQ�mFQ��ѵ�n���5ύ���G���R9;\�^kN�^��6 ���~kZq&"4�o�2�;[�Z�b�����RE��3�]P*N�aS5}����cN:-��;�ҤFwmTC{�L�����Qb�Qb���{NRJ�jX���P#�Wǣy�m�0���X�����4b�93+��0D��!0�6`2����"��[*�٤B�fm�J������w/���Oh�!_5�9��$��;yR~�b���Bۣ�ڎi`l�c5vI��{�x^ݾ�f�Ń��@TU�D��0R收������"]<+n�v׫;�҅���(���Y~��#H��bĮ������Ѣ
qF[�0��<�!��hY��S1^�\��+�m��ۛtkQt���C�m�Kȸe( �R����j��V�av�ܻ��8SI&�C����[!H��nn�a�"��^�l��@�J�+H�;4��������Rh��~�9x �0Y�m YƓ�,�%C��s0!�Zbh���y]�"�&�P�0�V����
���ƄP���y�4.oz��oF�]�����֖7�#�`�v��֋
EB�׽jn�y�Ds����)�K��.7E
`
�d�i�*-�gnp@��G�36�o\=kM�J�k��],Z&-8�.g=w���0L���լ���~�7��x]�眜�aD�EE��IpZpLV&X�����,�.�ji�I���� K�a��["�߶�1����������~�\0\i�orb��`���̰N�ώ"��o@0��=5�e��⺠���^���͘��"�OF��"��f��RF�0`4�E4^fwT!�����k�����=��e�a ��N[��e�"gg�rch�?<ۛ5kR2(��q6�/޻�l��$b�q�{�Ԣ�^]B�X������4y΍�\Wha�#,X�V�猄���}�2�X�՚X��l@c�;;g��Ϸ��H��[5.,^���H���
�8&*"f����{r�+��8�4�F��m�da�TE�B��T�#x�r��W/�!yʴm��%0Km-���8 �x��;�x��{�^��{��RU��x9: #���q�^�mIF�"�Ab�i �cu�5�'I��kٖ��,E��c�,�Œ2�R��pYp��&�������B7v������}<6��q#X��5��P��ĺG����׻�}Y�o�n�|�3||�rŖ���#�LR(�t��ݻ��F�Y7�:�d٥ep�I��+�ۻ˭K�-�.sŊ�Q�i�FP�����bvs5d�%�ۻ��֭͗cse;t��ş�� 8�ZZ�fә�XDeT�56\I+:�\�}]\�W;3�ż�<��n"B�uQ�OrG#sȽ�qy8_���c�^T*�b�^}Lz�N��+�y��n���Ck1�BS�
@:a1�	�r�$�2���s#��;W��,�:,��Q�3~��Ä��m�(x��+�T"�%8&�7xI�snB,]/�+E�w:F#DΫj}}���i^J����^kWQ�$D���)oI����N*$�J?E�"`o}�0����0�'�73e`CA�i?�� ���/���mu��B<�E�ն�z+��ܩ\#¨i9qC;^�^�ָkq�9,Xw�q�&�3�,�4�mY|⣳=���	����f�ϣ�l�4����h.z�j�*]nkv��<�:�3��*-خ�rX��WA�g�e��{���h��D��}��K�]Q��GY�J��nf&G�}wJ��M�=˕������usK�%=�8=����LX��@�n��	.��S�IUy�cx���
��C��]B�3�K�(�p�$�5���c���l�*AO��i�s�����H����rӃ%B���#amt�T٤i���\A�u�i2�4ZpKI��{6lpA��n��g���pY#�&-q%6F9ޘTD��'��6t�cr��r\�b(z�}��__�>C�"E�]L�<���H��&�E,"��mwx����k��	Bp�]���"��F\�`E׽��'�qD;i�ݹ.���������*���S8LY���/�?�7�}�j�.'V��9��?�����~�f�ũ�c"Ĭ����Qs.j��7U>���/C*o�D`�z�xp\��l��1��Z��]��&vnh!�w��ma�XȒ,Oy*�l~U��#P-*��X���{�?:b.��=�z%9[�O&��F�$8a���Z�n6���s��mr-h9�	[����gmcV�sA�8M�i�&�7�>D�#I���bG����.���pJȢ6����.W�Uג�A�f	��ٚmҕ&7��fu�w�q�8E�ɕR��%�|(��M������:H* �$F�ۂ(G����ˌ1J�faɾ����"��
P���]�-8C>=U���(Z}ʞ#^UF��"�J9^�^�F7���P%�o��uB(*��M$��8��|�FRJDH�9�BtF��2�4���ł�2w���b}�&��&c�����'���LX=�ߜ��u|���i�X��ڞ#�p�Y,�E#�w�(��L�i���w;�E*��J����1�e"8&`��5��՗�Rh�J��"ȱO���r�N�|"�ËV�7]I�|��n�l[_W�P�;���߹xI���0��sth9�.��u���� 0ov��4S��<h��r�h�kL��Оj���|�
c���;��d��H�ߪ�Eײ��KF�+\9iQ���B���_������?�ܜs��3z_l��:N�m���H:�Ѥ�p2s!Rq.��i����+�)K����Gw�!����Y@V��{){:�gb�;�����e�]hT���ma��C����uX[�k��H�ӧ$�D^���4�NW��E+{ �p�%���y<������+ҝ	�K����	��TxO@J������}����A8�B���BM'pw/Rr!�
�ty("������|p��B���OH�������|��&,*Y��X�ړ��;���m$]n�F�k���e�l�<˗XĲl�w;��0�km�&��K���nX꺆Xj.��n���q7a���k��GN0l��v�ag� r׍\Wb��d�jv�^�8�ŉv^��V�{f�#cq	,���6[i(�#�4��e%W2��(+�svnX�V[b�v^�#>l��� wݬvHm�lcl�t�|<xJ��\�-ԭї`���Q�`e�5��'齯�>8CvZ�FvN����J��_>�/����>?4%e���X�IG��r�YW:F��5|ȕ�����a�ʱ`�Tg]���s�r8%*��)[W��$V>��u���"�Q8g:��� ��{��Ɂ�?uН�|�r�J�V��B^>�F�)��{��B��#��<E��M4J�U�ZYi�m|��w��	�&�(Ro�y�J��mt�lZ�ָ�d)�p�8e�՝����F�/bL��2���e6-��in9���v��C�"_c7�EU�۰(��i�,��K\x���+cra�+@\fʤ`�������0=���*�0!��V����#�12��&����"H�*^Ԕ�o}JH��e�\`�Xn�:��DF�fxuK�ٕ��Wz�W�ើN��Ĕ,R/�J�/��2Ң!1R~G	�)�ӂZL��l�a0F75��&{α�֕	=qD��ǖ���Z�t�(�f.]�����Ib�h�$P�T[g}��RG���V
�[������=F]+�m�∈8w���q��l����Z��:��8�ͧJ�2���Z�
�4.��f�m�"�y������`,�b�W���E�zE�w��m�u��T�sM&���ܤ>wA)uܮ���ȥd⁉�*-��i�ю��������0�W��JTK�#>�DG��*$�i��T��������~��[i
��BVZ�k��o+�����3��dö�<ޙ�9S�!.����s��p�j,�ވ��}��9�!'�7��0B͈�:bU�(�������ӣ(����1Q���y�ƕ��j� �tgyJ�[��B�����N��+�+yd�+{�U�UP[��Ҳe�2������������2�t�{&�z�q����<�M �{�+��r��a��(d�J��>Yn7U�yaۭWN2q���7�{����Tw	�jf�Ќnƭ�f��л&T�QEr�v4�(���E���,�0Zl������!x}2[�����UO_9S��L��t�8T����,�R)*�-CG,��p�y�۽�Gaʉ�Kzf����_خ���?Xd^U_w}�E{������ݒ{?/�����ɣ����i%DDp�KX�l���%AH�jT��xJ��U�KK^�q��h�m�"^ ���x��� k�)�g|�H�x�Q`8ێ5Ҳ��Tz�s1$�(IYH�%���;�#�uZ�Lt�vT([ģ��d�BF__Yl�:u�|�]��V9�s�fВb˵	i_u*�6��zԜn	���6v|�VuV�S2$�2�bp�iK]���R��y����y`�R[�]w�޿�V�S50���������X�.��9�]�Nk� ���OhҞ�� ��C�<�N⹹�s�;��)�㪽)�|pw�집�>B| s^x�Jx��E���1���^�iJqkOB�=W A�N��\x88TO'����-ק�<�P�W�5��X�5�, k}�I1�����qq�L㖚_��� ��;YX�b��C�F�w�]P'U@�j��s�>y � ���	"$ޑ4Ÿ�6�`�g8��
���i-�)V��DM4�c\�5�q��� � j*k�@��q� iH����%��gY6��}t��7�l��Il롊� P8A�"	|�^X@�DskYX�Z �����]�ܶe�Z䴹z���}x���Z�P�@7��q��4�Ӎu��A�A���EJ�m*���ײf kƺc��ЊH�m�a// ������� kKq����b��h���`�D�N1�4��A��`5��D��1 6���;��Ң�����(Q
�Oĵ.��R�r���Mٰ�S�k�mZb�[�e�BÚ�-&�YS]33D�SsJ��{�|���I)!G�#�֎,�`�H$���W���@�$S]���L�6�B�
�����4�f)���|	�8�QD7��RA/� �cn1���no�/�5�V��j^`�*jVY8�YdS)m�u�C�L���el��iL�9���DE�`��6f������
��3rV�r=<�aȐbd�;�9a�NM�}�۽b��_�L�T0�c�j\gMt❀���
�v���:�����E�#V�2���)�_}j�u�lm:���% 9�%�%���3�!YT��W�oN��b�*(_��U�QF�yzuJ;gr��A(\j��j�_z=�k���* ��Ȫ�p*�m3�_}��n�}���T�m���y%4^��1He@���j���:.ԛ���F !��+�����/���F{���N�k�3������7F�sn�ʮLm۶��um�м��,=\�=��66"�/��g��Z��m�2��:h�;�s�if�񀝠�Ӈ�C�.!��H��3x��p������=��癭���]ˇ��D�Q�G���h�W��e��4	��M-��=5�!
�"�zv��y�j��������`���w��Ԇ-���+ɽn����H]�\ԋ�\�˹�,3�>����ߘ�{�R����T��[6��̓r��\ ۬������jf���k&!0����+K�y���9u4u[�l��I��W���>��D9��_g�'C�9��J� S��}��t�2���JN����]{⎀I�#��ӡ`s���Ʃ6��2ZS�P������]�ܚ4�Dj�-sя�걶�[;V]��'s�H����pbʺKN�\��AE�[��D��`HJ'vr�o��^8�fVS������l�����N�f��s������u���n,)R��5u�)�q��=�LU�����ovr��򶆘�B��IH�L����Ч�>��<��^=oYx�h���-��m�)�xW�P놽\�7y�|�����^3�����yzP���x8㤨��<p���wp+��/=�}�g��[n��K�NI��7�v��M���G�!�]�aH0�-�s�`�͖hݵ 3\ǜ2�K�g�4�f4�bFF(i��mzk��+f !������1�cu��,��Q�:7Y��A�r2m��j�v�HmGU���a�3�IԳH�3I�K����&q)�y�Ξ��u��N�1�lUT�q���҃[��6)i;���kR�Ǩ���li`K�g���A�K�C6)�hƲ�/e9���+Wme_$�nj3[yh�����o?;��?�[���������:��o����i ̬�r�c�����-[	���[}������uF:o��2&�@���lek֣興�X�_�VF�y+���Jg�BYP�ܥ��<K$�l�8(�d��N�gn�!Û<��x�
I�>"zط�7k���O����#���yLF��-w�>:q�̼RI�" ���X,��h�Z���g�ܽ��ЀX�Kp�����������i�c����+�|���Igp���z"#�u;lV�ySB�Fm��8I�I�[O~��\l0�gw��WP-�P���z'ry^%�B����*��f�z��j�eDk�&uy��St���*����C�\:�Wv��s�Z�n��xpF�b���.�S�-XmM�Wg��2kr��������4�P����*�8�"D��骱�32��}}W�U�4�U�c�gb�)��}������}���^��7�@�`X�4R�Q�_z"~����V�̧o5^��kŁ�9m�+W+���-CX7	&���[=Ieo�`�]q���t~^�١�ߌ���i+����?O�����7->�'�̗���̠�V`��[a"�]��d�:ܻ�B9U>�"S��Q��H^\�#�Y�W�C�N��r*��ۋi������u���g�uc��,�L%�gn�'�6n�陜B�d����b����
�������/&� �$��L٫|�O���w�z��0Bi=�n�K]����mrV�~E�|O;J�P�h��9ۊ@v��
�X� �0��{��;x"�{�f�����ua ��]�s�Q&pDR�9�̌Q"j0�<pR��o�w�Rq�$F���	)�'m�h�/'�1��ټ�����}�4F���_:���3~��d,hu�p�
�bɓ"��IL*@����{US�|'0�?-f���bQP�T���2Ȫ�u�R;�>\:�S�*Y��Nɚ+]^�ҭ��W��^|C���B�ws{��>u�o�9���#�t��u*C�^��QQ좝��ɶӻl}w'G-����`J�A���7���)s�|�;�t��f�����;�5�d�U��vҌ�	�b�BP��a/S��m"S��p�����m:�RA���q5�<r3{���	H[�%!	����l@@�g����<)�w(��n�)!�i���!F}����ߕkf�~eE��˚����K`��0ٚ`5$�8E�)���z���w£"��;\�Pu��')SWܼ��ǉ]^�W�����R�}�G�N}����ȘRn{���d�m�����ٽ���:��݊�c�QCʸt+��R��q��l�U]&��ʑb�;�Aoi-�8������=i�;/3��#k�\cW_���3��Z��FUNK�Ձ��wd4�Ý��g_?���_�`�!��;�M�,�2bjVmv�1	X^}�z��m@Dt�p��&jj����NM�}כ�XP�U���;P�*'4���������j�#��5��󯁟��q�B�x��DZ�(b;��J�דRq��h���"�!�-=��ч�E�����m��DӍy{�W��]�{���Ҧf��{�}��y5O���������.�0n��	Q$�{ۜ;��T0�v�Te�b��w&�sŚ�y���b��5yG�l���r�㲒�J ��=�VU��V���<
5C��m�o�;�tp����w��wn,���{��*@��j�P�BVm���Af�D�F�ysHI'˖>��+���OO_(OY�5Tm)��ˬ��Y���ΐs.��*ic2"�Ն� ᥠ�sqQi+���I^%=Ϊlee�"E�;�X&���]&�{�;�ɚ�B�0̚"�
%����΅"%�E����=<+�nm^�S�UKԕ����س� "D��͌
�j̚�{0F�B
�s+�~e0P�o{�OE�Jn�{�γ/��<�wH����J�ِ�����6��b��S��EW��Hީ�H@RJw�NPpy�J	����4]7�o�x�t+g{�d���e%}�|6�Ub�.�ո%zxm��u����ͧ]��%�E!V*�K �P�%4��oqFБ�[��v*�����d�s3d�-�y;��,�H�Ƕ�ڸ:�̗ȸ����5|xV�>�1�oT�{�1�c��Bp�I-������k����6f6'�k�n�9(����&7�Vnq�Q�T�Z�P��zRR�p���\���z�1Y�w��j@eg+�a�W�������F�gc�Z�-�Z�޾��:wt�mu��]X�� �� ������� ����_5�889���qk�ԁ	' u�B5�������� !
pR$��=�<Ġ�p�Op*��x����|?/��R�	B��g����ծX�������٤�K&%��*�\e�1	s�i��&��uM�M�	�s-��-c�`3Ķ5Dl�������ݫ���j�yv�6��Mu�ϩ����Lnk�ݖ�u6��QtX,g���\R���B�,좦g�0��93<g[��E#���uJ�E�.v\�����V-�J�E�5)�kj�is�l\cV�����ņk[��f���bڥ�K�3�t�ј�GU�L&���I��p���w��Ŭt�%xfJ�LY�9�e�r�Y�' A=�|����ܠ��%,m���h5���Ib��t��_W	�s�>�>o��eC�s�2o�_O�L"lXb�;k�U�L���5tp��h4Qa��޾�d��3�)o1p�뗣�Y����Q��j,�f�3T��wm��32�z~�z��B�-�3z������"�w׺z,B��4�a�(�ou4�*	����8k�����ͩ�� 8��9���2��u�&�_Q�ci�d��ࢋ!�i<��Z�vg����4��"o��I��X���S�}��(k*E��D'>���³���$P��/��` �i2�^F	p�Х��%[��:�\�5#!��$���.6�uհ���	=�7�(ڰ���3��wj,DfL.��3��B77���!!�wK���0´h�
���L5�����v���%x{��;v���G�;�W�Wu�����X(�;׬mã��xp�+΋�әu�fDdՌ��B-�Qi.�;H�Ζ�>�h�v����V��P3]�Z��şn��t�RF��&�jH�쩘B3��'�16p�`(h@NK7����`�#7�n���.�!�U�inmQ�I�R����-}MT���Wx��)��qu�Yrv,z��%3�8��)���}W�{��uU��3���a8�-���Z<}�YMnm�W�灸|�#-�W���h��qp�Mơwǟc҆����(M�t1	�I�U����(�Z�oSf���0��T�5c�����+����hB�,�Ƽ��]`��>B�{�'�A1�o�zv2 $����I80T&�M'������<���ݳ�]�ig
ܸD�1��ӮKy=7բ�3���'"���Q���)bd�Q]�7H)!�b��`l�Ç��o�w��1�.�<(Z�tcZ;ӻq���+Y���(S�\JUaZ�|Fj�.��aI㸔�Z��.�Hˍ��ݷ���"�����r̽�w+Ns��ȳ�`�i��bhU���*��{[с}W���l����<�XSiǭ,�������d����E���8�������J�}zet8W ,T��c�Z !�@���c�6�@@����Bp	pB�B���� q%�d p-$-���J4�!�M$N �4-�g2���B��uw�附)撵�����w� ������q�9�/r㺻A�hF����nՊ�j�"�g@��W�d�r&N,�q�u˶���6��x{nZ���i��n�����.�nc�Nz�b~r�hYK���b�Z�1���\+�y�F��Qu@i�׆�C*׺�*�a�He��d�	�Q`6���̉���b�"M�uuJ&�VT�웳�̻dv�)�^�u��">����{q+���Vz5*v!���Qqbd�u�D!�06v;���`8';���P�{g��ղj��(���(mP���٭l�&fVwy��>�p�����6f�Æ���vv��x"%���ۭ>
7�"�?Qj��SR���Ƕ|�w��?j��\熐g�;�C��6.]�X�P
	�`����c��T�=w #<��� ox�D��u��g�>��y�e�c�i�����_qiOj9�="&�7k!��`�ZK��o�&�z���n�q.��Vﰈ�)���M��w�:G:b�A����z�.�v��j�ˍ��jI!�\6\/$�p��smU��LŻb����9{&gseN���;���+�f���ww�-r��������X�KnToV�ST.^r}�MB�<_t���q}�fb�T���Z�&B*i�_wA�^�v��ݾ�D�*o��#��7���9�n��Fq~�2��*ȥ�-���ai��PE�H�A�ݻֲܶu!1�)D������fv��zX�h�Ꜿm�fEwu^�T��c5�Z1V>إf�9E�SI�n��#D)dN~����_�7^Zұ��b#I]{���"�'/�$*� ��;$~�f9�s�GNd�pRT�
N��[!��d4�oo{k�Ի��|��;�/I�u�ҮA�ܱG��V�'�Goys�ZLY��~��v<��s�cb��U�j��g�푺������C[���������:�8kV���ݘ���1��2V�7q/[�ѬNKq	���v�wP1�h�f�c�����ڇ���f���-�l:�\�z�0��LWVwo�6��2=7q麮�AV�9�k,����ry��X � @  ��!�IP��B�����d��,�,B!K-,
D� �B@�J^J@��Z^;�ؘ  ��pB@���$ �K���>_g��`�et�ن;Vz���^�8S*���u�p�t6af���/2ܶ�MٴK��,��MX�<۫[R��{b���iJ �6qF�tk�Qn�M+��l˻j�9K���^����w]���۟Mǭp/׵Dd�>�n�!`�-��a�˃����G4n�'��խ��Jɥ��ݞ�v�vnq��aI��+l�k*�(Vș�"��wx�2m�.����N4��%�k3ml� �`h���h�h4���?!ͮ�=uwKɝ|fx�
��{ت�"��}�lU�9�ڣ1wd)p�p�	��{:�1LU�EP�ޙ�ԣ���E��r`OP��"�}V�.�;�<H�B-�1(Gl�	�
�O�^X���&��[�S�Yo�7��*]�#.v�1LW���yl�m��H[�u��v5�w�U��ۻX��%[�'~PXI��𜑊3��ǧt����ߕ���Z$�6�^E���%w�ɉi�fQ6H��)�6NW���Sb5l�s d)	�)>��=w{*.ˮ̒ڱ+��33���/?)頏��+ކ[#܉c�d���	F�$��q�T�@!�Ђ�%.��:Y\��\1x*b�{a�t���ќ�W����@d'6�RNM��ᤶ[��S}�Vx��Z��j�K�e;�Yx�3�y�^g2�Q��:V�,a��"�]]�g����sn�o"�EA�5�J붍e�ɂ��}�I���^ݠ�?828��O$���Y�wu�m̼�`���wov�y�.�p9dH�#	7زu�`R�S���}��,g7Z��TC���������I��L�T ����B���7}]/v2�ȉ�O��)x�� L�Q	��ۛGjv�R
�42J�!�P�.q�g�p�0M�v��SyQvw��ʦ��5�8�ї�ψ�x���[_1Nv��ӳ{L���4'pVZˋѺ�e�f�ya�)Gk�q�az���M�gi`�g��V���rڄ@p�eE�Y+3;�ϣ�Y����͟�#s��
76٫�g6�*��a���3~|� ��ǹ`D��
}�Ӱ�`η�va'}+#oq
��L�z�v�v9��9\�
�C��a�]h0��od�XuW�X#*�cb�I��m%�[W۬��{�LȽ������J���D�������xu�\�����%����A�9�W2�>
]�ti�x��Y� u۔�{{�"���p)�X����n)�M�Bî�7wCvݠ�(Y�-�ً��������a��m�amHIs����׃���J�ò�Q_+�M�Y�hUH��*L���}�*�H��Y�o/*:#�]���)�I� @�$$�1F�$� c�!�%!���� ��bpH��'���8< ��y9���v H@�B Mi�%��'L]·jĹד���B� �&i�EÆ&[��۳�©��<��Qa��f\��:]}q"�uԙ��rs�vԢU��t3�Rws�/+2��B9d�c�X*H�)�(���ǣ*k�gw���q�>a4W�jX^n�zd����o�a��㐪���yrh_����6~W[m�l�"k�ͼz��^���{\s<[�CC��q�s�S���84����(F�NQ����.�W9��-��<y]�/���/��y�7"ǡ֎y�°�p�`2�����n�Ay>��3�]q���٬��#]nډ��j��ǘͮ�F�����W�䃐�0�p�*z����D�{�(@�@����j�V�Eޏn�LL3�F�o���2�u�+���_{���Ve�
��2Ǝ>.�l��"�[��6"'��P��#�s�pV��H�[`:{{U����b�(��Ң(^���'��;�4ЁS�,<�͖z��F�dvc�ӭ�}i����e�9����F���X�*-�ʄ�J����#��$7qnD�I!��1u�f�Ĕ	�8�%�m���H�`���a�v���<���FF{���4��/��Z\�t��2FE���r����%�6wDUOޣu�0�C�^����IZ�-�h���,�&\�b�����CW��aHL��RH�
�y�ݐD|,D0��ȱI�T��x-	i���\%v��z%dU����{ۯVw�%�Xc^��Pe��)"��O�+���<��uV��*�h�j���W�K�h�:�m�U���^l`b(�5/X��g���͒snV��p]����+޻�0p��n,Sn.S�|.*x�E[�%��d422�)&���ڄ<�p�GSXFw��A�<��an's�~���]��D�U��_�W�
�yQ��ff<t�=r�����M�%�3��P��ٜ�E!q.B4b�����8pM���F� @�YR=t���z��Tj0TH���Y��U{mY�i|����̻M^��� �AX��\�SYwp�U
��&3L.�F� p�8���Q>&1����M��*����;����<ǘ`��"�7U3LKH�i�r]/_�ZQ �����������8E�LT��=�i�cj-1
!!�S�{����a$;(�RI$�|�PJ<Q@@~��d@@xoG�e�*���kJ�E�>}=.c%���ܸ?��_BȈ��"�4ŀ�09D=4��o�vG�����N������2r������^����pm�x��U��e�c�ckӭ�O�9Ԡ�5ƭ��Ě��AK0X8�æ4o���	��|��_s>�p� ?�Aʨ ?�;�)lw�俒vPv����>i��G�����o�y{y�(� :� zW�g�� ���l	�������t��M��+���{�W��B8��<�|:��u���g�,3V� �ߖK"6����t��[$%�""�(T{���p�3H��,V9֑j���0hf�������s
�3�N:β��y��t��<)�.��	}�}J����#������?��B4(=�;�,�A�Ny�O�;������}���UY�h
t��.�>�c�I��\�^��P��$<�������<Q�{H��|=c#��NXMup�bC�ҍ�d{hy���Y���0�_��EJ^��&�GSC@����" 9��B0~cf�頟�����(phAz���`o�ض��ͪT)!�a�,�sG�F�*�m`��
��� ;6ga�y�/Zv"/�w���I��t��}����ߨ��nu���RXǿ�9^����@�:������q"|S�!�:Rߏ_#@�������z��uN�>	TR�>�5I�D��ϱ��?��}��?���n�	���0��n��hG"�(��Qr�e��pq�>6g�����\��kcGmè�?c�������n�ӳ�%��u̦�<�
!ѳϨ�T:H�N��^���|��8�$�0_A�J\�}��C�go1@{G��N����,���C�fZ]H�4���[S�	��?���<u:?�.�p�!��'�