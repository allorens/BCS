BZh91AY&SYBJ��6_�@q����� ����bB^�           �(�  @M�@�4� �@    )�@�   4���rٻs�1:�U2lf�ֲQT����hPJ�KfQ E��6EV����&�f�) Q�ZM���%� ��Yh`k)U*�%"EU%*M���3`4J͡+k26�&��BVl���թ� Y�J̬�̶�&�R��Fئ��m��W+L�Zl�p  .Dx��[� wj٫J��[2�km�����f�(�Sl���҇U���7[UV��gE;[l�iӥGkJ��Ŷ��j��TkMcZ��j�  ǀP Ճme����r���ta�  ��z(�i�z�׳��x  識��  �;��JP{`)�r:Pi���Z�*�$��Aj}��m�fV� d�� P�,:���up)� �yX �z��y�lm�+�S�:P���t�إ_:w��{�|��Ol}����

 o{�RA�*�U*�JU� f���R�/>w��U�>>����A��}ϥ>�U�{ ojP���8z[z�(w=/� �����#�t$�I����K� 4޾վ�B���O�[m֔�k	�4|  l���CA������  祎��#��@'��k���z�OJ���� �i{�n�� n�\�(>�z�U*�M��£"�Ux  <E�+_o��J /</w��*��҅(=׮{ءM({׳�S���7{e�=SAE�M�E A�׸Sւ����֚�y�|ɛmhҫ@Ѷ�f�m�   �� ��Ӕ�=4oy��Mm����҃[{�xt�nۇv;�i��J:��p��T{���� v��ր��( �'�Ai�$�α���3�  ۷� \p ���� �рth'Lt 4� (��� ���CgZ� �N  6���i��ʭX+E[ff�|   �v�: WX CX �0 0`�nh:}�� Ӏ 3;m�(4s ���T�͵,Ͳ��)��P��  \� P��� ݲ�����a� �q� q�W ���  -���{� ���       ��2��P    E=��R��@ 4     �~JJ� ѡ�@C@4  �?�)F      �~@'���F� h     ����Dd�zjhʞ$�'��4�oHɓ�������L�C?�&O�6+?%��p�^uV��om�~�a�m[,/Ss�w�� {�� <YP@EO� @U�/����p U���>���1��{����J�� `�z���'�PW���,	S��@W������������8ʟ��|�9���	���`Ol��0'Y������`��	��(u�:�`��X�/X���A�*u�:�=`��YO�@���z�=e,+�T�+�N��YG�	��*u�:ʝaz�u�3u�:��`N��XC���G���P� xe�X���@�+嗬!��(u�:���@� u�:ǆ@�u��)�@�u�:�YS���S2��:��`�Y�!� �{a�XC�� �u�:�a�YC�!�:�'Y��P�(u�:a�'Yl�YC0'YC����u�:ʝd>X@���z�>G����/���A:Ƚa^��P=��P��a��Ys#�P}�(u�� �XQN���aE:�
u�T�
����A�
��T��'Y ���dQ:�"u�D�	�TC�:Ȫu�� ��D���S�"'YN���d:ȫ�¯YN� =`E|0
�XAO, ��TS���D� � /XE�
�`:�"u�T� ��T��XOl ��̂�YAN��eQ:��u�T� )� ��Y��dfD�"u�:��eN��YS�!�L�XC�	�P�*u�:�a��XC�ˀ:�d��@�(u�:�a�X~�XC�����a�'YG�>��X�	�=�`�$�������?l��m�i�UH�PW�n�sQB���A
v<6�����Ra{f�g�\a����x
Z����.��ݝ�M����74�/1慙��p���753�5��9��N�V�@�B\��[��Gp2�m:�
�>R�[ۥsxL��ɦ-����9��lM=��ۚ;!-$p�M�3L�2@��8��XX�۰��2nC�f��W��_+l���-$N�.Y�=;^L�֓0	����7�3�p�ɳ�8tv�{u����S:ߨ�hSw�,9�J=��i3I�F�X����w5t9����w��ᧈ�Xx��� ��Ղ�[�F�0��Fr�xi�A�U�� ЯA�S(ͯ����0��� <�U�S#�˱��[�.w��"%�^Y�1t��7_ŵ5�Wx�]�H��7坆�+D�fosɶ4	CD��n����;_S������k�w��[1VE�B�k>�y��&��oLޘF\"�Dy�5�.��y����.�1z)�v�l"ٹ�ol-�͇s�i@o4%1�{d�0S��g�5�;{t����f�o@�Ѻw�F�M�T��U�2go;�A��C��v��wp�����sݤ�2�1΂[]zm����*!$ ��S�߃B�I��2�=l�8 ɽ� �f��6�·���j�z0�ؠ:�9l�KW;���oڔ�5KݢR�+ۼ����b�YBh�n���GN��'��v䳛���t��1�����4)��J�:�K8�wJ���� t�L�ֳ�[�ZP5��ɓ ��Ls�M[�A�fK�N�j>Zdh�8�#���B3��٢b� [���.�{�\b]@Ҏ-�s|����R؛5t/��{u�{��/�������۲�r�X���0�}kܚ��8�V�24�.�b�TP���1n7�����UܻZJ����|���*7tm��#ٵ��Y��R�x�iؖ��<��K��r�x����FU�5�FM�5b��Ӻ���=
�ݢ�}�wP5���n��tպQ�͞�c��L�l�.�C3�S��w�[��+f�0���p�ww-D��w
{�VA�݃Ih#���@����k��٥���nU��j��w\흘�sN��[x)��V3ؘ]���Z�V�v��Ž�L�(�uHq���X�2�/�� �s6>գ[�*�w+�/Q�.���ˢJn�;�@T��F��S~�Ws�j[��A��$����B�ۊz}	�����2�9[��N#'&�� WB�˦����2�ɼ,!p��v��1�0qF94����,�ˣF�E�S�).5��e.-R�n�>���2E�*��c^�Z��A �f\�ݤ��&u
�q+Hj����[�Zm8��t�c�ǲ�wG:#��uˠ��pÚ��:���:0��c])��%��RS"�)�v�t�A�-デo���� ��LK�p٦=�9�֤���M-_��j�96�"GP��%+@��N3HRe��DZc�����G� b��j���`��)	��|���U��(��@�j���k���R����5N\a�pz�R��^����u���+���R��Nk�6̹��uf���oH.Ԃѹ�ve����ُ�Օ�a�gf2� ��;�H���N�w� �p�iw���7t�5X�0L�uh��2�"O�p�C�ۼzq'+ҷh}SGn-�	�3�Ot]\7&v�U� �<�yY�QŇ܆Y�wOc;�[H����U�����]ګ-���lN��ދ8�� S��x���j4��������x �/���f�# ��r��d�7�v���U;{1��5M3{�ʰ:�C��L��e��r�����s���۽�k-�Y��|n���RL-�4�$���^M�7sx�!j�)��$0�a�8��:�#�.�X������ik��c���@]�*�>KuGrõ��2���d�#wȥ���ۓf�ն�J�N5���V�v��c�w�m��"ދ8��cN�F[�ޫ���e5���i����=�(��y^���b=���|�^1u׉ )S��|{N�n�Cz��H�v��\�]�j���-C;Y�&����8 ˥�'_E���}J$\���Dr��ݠn��lo�¦Et�ʪ;�)jc� ��rK-��8	�Z��&EvQ:��[/p7�00- v�>B)�
���m����;*��Z�8I�ǽ7n`�9hX�I���cV��p�r����t�j�{��SF����rݫ�rO�@^纴�#� jk�ԋ�ڱ����vO�;(��*	�c�/=�
h�f���,��A�wu�amѪ��$.�D%5�ey;�������T���ޞ���@�_�,=�q4�>��������'����G�LL�ݍ�Fqv���>)]c{e���Wj��t���n���w^��˃v�Kz���sN�����rkJ��؞:���IҎC��Aw
WY�y�5�V�H��
󆃻�"�r>�r�;��m��ΈkƦEә��]^���^ZA��a:��ڞQH�=A��M6qW�Wp&ݒ��霏3OeJ���f�751y�ol`��iXİ�Jӟf	ѡu`�5{`����8�|��8"w6��a螮�8����Ws�,NY�nr�Ӯ�ۧ\���:�ٺ����A�<n�Gi�b��<�W+��yȣ��gU�7�[���޶����v�D�S.��=Q�5G`vS)�7�^
saM�8MCp����`K!�o\�R鯞oq�$�l�Uf���_N=~���b�8.��Y�:�K�޺p�_Jވ��A���Օb�'<���m�Q�5�Kce�.�]��<�Z0f=81^��'C�]��۽PPy�t�E$�=����i��i���ע��c��5i=�j4 E����7�6d�vr�D��!STz�7�=xT�9:��(5r��o&�E�-ڹWY�zf�8E\�nI�/nm�'t�\{�).8ܡq:[�|l枯GۄӼ6���L=�
���kA۽74�k�����3�8[�$�����b�,�c��
l"��E��f��r����×.�j���)���e�s��޽ ���|��x��r��n�����ܫ����@�ΰr�`hmo_�دQ�?�2nErX�P�&S��'����sb[��v��]�'�t�䤽�Ϟ%W^%t1��g|��ۤ\�nȷ�Y2p]fA�����"�#�b&S�dǭ3v�f0����u���I�/qI]����7��q���C΁�Ov'�u�$[���T������ko�o0�G��h|-^Շl��X{���_ݫp����3�J�Cp6�`4�=��렱R��Ι_e�J�2�Xp�
�q��o;��$�9a�k�Nt<�A�ς�ն~,�uc@�]cP	<ź蠯����4'v��vؖqO���npG�M�!j���\;��G&1���.c\��k�T�"3�jR>u�b"��T܁��Ã�hJ��y�6�C����x���������H�D�R�v9+XE]�J�Xp�4r�}�*��@�,`�5�\�ب��i|��WL�9O+����Z�g;�Ǹ$���.�7�p���{E���7L�b�e�Μ�Q�Sw�*߻$D��:L|u���l�8��]�iyۥP\�-{��o��J-��.�	Ӑ�вN��
��]B�+
<ubN�Q�|�]�uD�<&v�r�c��WF��RGugl8�f�b�u����!���1!�%���h�)P|������]v����:ɬ΀Z��2�Ӡ-�h[pǦn��XtT���Sc��X*j�w#+C�wF�^a�^��g��.BP��vB�Oy�ɂ�rb�t�p��xܹ�q��m�u��z��XA`�9;�J�Y�#9�^ W#�H�ѿ5����Ba��\��W42��I.ܴO���灬v]1��]UWWWwwJP�B����N>�4��+{v�BG�/�wwIuu��,I��d��+��J|�?��Bs_p�ʙ��>��kzo#�
�|μ;B!�<�K�6ܔ=��w\+�CFߜ0�i�KLf�.�a	zlK��VG+��'FfBfv-�۹p�h@I�
���e��Md׼rl�M�Y�!Y�L�{ enQ�:��<w�]�7�^��ɝ���VЖ%�س[x)ejw �#hI��ot�CKt-���Z0aʥ�&�|;p�f�BBى|`�k�AȈ��/n�Ba��T;V����#��k�`w,$kYt�-��'6��hY8@\�J{�:����jX�U�RQ�e��2Pq]�F�H$�1�On��԰{��Y=~6�Vu�ƈ�oWw
�D\�ތgR]�h���pNPs&G�;��\)v�xf𚙽��Pg-�5Q�Z�R��}L-�g�"�*,�p�&5����lv\b0M�Ui�{t0&�]��	Zbs�睉��^��ɻ�:�\x���͇�[@9�{C�BF#�%��%��8�f�X�C.��^VqB��-$ŵ%<;��	x��o���_3��՚L���3K�s�۩�;��L���.˽	`�f\�'Zik�g�7%�'��T�MQ��o^�(wb�1���XB����-�@Xr��z�I{�:5�<ٷ6��,�kJ���'b���flu)���o�z�y��77N�z���w�*m��.�Om�"���¶��5R�L!w�z)NG�J�����Heҍu�Z�O���jq�9r��8oD�ZAPvʸ++���:��d��
'K����9��j�1�ޢ;2lL�0�X�d8�l�q��/G�<G�]תx1	n���<���䬖�Y��������4��,�ԄGW	��a����_91�c��q��js�ov��r\��4��-X�eo�	��lY�ɪ�S�!!�P��`��L�3b�R��c��=�HT7u�;4s��[�1����ϯ�"��oc���%��vm<�t)�m5��P�5��ˈ�p�͖ٸ�k��B�L�M����˹�������핃i��M%�X��M#���N��CD��77�H��i��`�(�L^�f
��h��ʏ`��"���[Zb��;�'��S2�>t-/DxSt
^'��@�K������#jdM����b"���)���#q�,o.���Ni�_�qT4��d�z�6�uN�r���@9�Ͷ�Wo���f��bF����2y�?��c ֯�bۻ�Eo^[ʎ�C��Y�_P�Z�����5��ͽ0ʠ�5
�e�/>�7NC�^�ڭ�Bz���y�oQ�b�YC� �yW�|xi�����0�@�
�>��z��[��D��m��eՋ�ZH���7y.���i���=]��j:�Y~����L�H�o=�e]u�����uj��*p�ѫ���No�n	��=àܷsC��F>��2)nYxciA���s�.�� �ػH�����w��d��{�D���m�aAj��ӉꙢ��1M[,�k�H�E��H��xvo��y.�"�-N���D:��X��IԛۚEK,��٫B�s+ٷ��T��ov��V�ɭ���2�\�8�����l�λɈ��v��e��'�Mʸ#��h��F������$tW1��J�/g.\;T���}!�����o`lAhB3Ϣj���i'�JmsV�V��h���i�Sjb�n�l���q���h�������j�0k�`u�N����Y�t�i��k"Z�Ԃ;��3��_]ʓ�񮱔+O��W^3��8�M�g(v���r�c�h$�´L��m����=�zW%��f�7's�������K3��q>�l.�تݶo�Jtp=7xʖ�'&.�w�nՓ�*�NGJ���.��\�>i���{�^p � f�����݊BS����[Y�S1E� "�n7�{�x�R�7QWj׺Ì�o�����q[Ӻ�]�j2��R�kpZ�~7!j��R��o��g��⻫E���ܓ��nv�;L��:>|��1����˘��=o�F���%���b��;w'[2���i�O�f�zבM*�6=���Q� ���]Ё���'P׋��{�j�y,!������N�/N:ZM �9�u� ۳w!���;���.q>�{|�YdhQ�brˬ��@�S�!�ʌB5f(����=Y��c�3&��^dk<��5��id��1�QtX���7&t���HD�t��]�;�H-�$m�W�]�o�-�A�V�F�L�^�f�@Ge�˦9�h]vo�p
B����{�gn�s;��,�WY���<0f�j�e=���5v���:]�1�U���Xu��(܈�#E���/̙�i=�����J�O"��R�J��\�Გ����<gx�ɤ��e)N�Q��*�i]uRS��t)�)JU��l*Ę��:!��*����� vE�4"9��@�d)ai	*�p�gnWiZ�[k3��J!-E+��<��4D����a>��z'�:o[�Pw��k<U�BU��l�����!W\1�� �d��63ev)J�U��D�Ki@&R�b�Z8�Zל�}�jX�.;��I�d䕖�;��HB�`��l��"0HF�)��0�x���`WŹ��>a�:�OC��)�����m��-�u���qC���}�oo��_z��xO�`���CG�7���<Wn�u�ȭ�r���vCWK1θ�V��
qc˓Q�Z�/�l��-ָܜ�p���ڲj��iȅ�Ki�L��wJm�ݚ_<���ȥqJ#V���_]�
�=�׳��k�X-g]=ه܎m((%��8��M��F��~�vAS,l9�@%�SH4]��n��{w�Q��<{��G��
TԎw3v�;�N�ʯ�؟�5S�`��`�s��v�T�1���J�{�&u����.���ELg�!�*r���u�2T_J iY�+����4��UX��e���Xcauz�[�a���]���Vuc_$R!��v;��U>�g
b*�ϸ�ړ��`�Pޭv5J�=�r%�[�ּf혆X��.�KAn��R�K�B\[6�� �d���4
���o�ݾ�$^�;�_�	PlB,�\q�ȊJ΃�tK��v\W��
%/��|C��� ����qWlt^���Oc�C�h�_�u���R������,��z���ދ�z�a�J�rj������y�/���Z�.��u�0�|��%^T3U��^�\WS"R�wm�,L�6r���IcH]]F�b V��Ղ�;ck_Lu���8�HQ/v�r
�#�݌��o���yKP�Z��\�����c�gW�̗��P[�<�ʱ\��v��ݘY��5��1)�읺�\�'�R��P���A��q�k���8�v�S���w7ͪ��8q���+"�q�5�t�s{�P�l+�n��} Ҡ�EuN
�f}��R�L$jegW.�������l:�;jڻBȾ�:GUw�Iu]1[/4�7�OK��orۍa�L���7o8�*m��wl�36m.B���㓛��>��B~��"�7JA��<G �;���G����C`bc�^>T���j��V�:/q)g7��o,�eM�g��c�v=曣Q�z8gY��$���6\�p<���g��3f\��fpeV� [ 	56�����R�b%��3����n{|9��n
M���*�v�rm�{��!��}��z�߹�^��5I��:S�X�b�s2g$(�щ-xànb���Pny�Ph���k�U;�n�;��5ޗ�!d-�>���o��5�P�n�{�%o���Et����}���;5��hl�|��0`�f95nU	se�=\�V�@N�^]�,�x�ʝ�-p�t_D��Q)8�����ʫx�;�'ѥ3� VA��wa>�T�Jg��saZ;��;r�<$��;ذij͈���0F�Wǝs�Βٽ�j�#�U`j�Yk��d�]W����yWi.ՕeܽIc�T&p�kG7ln�wA��F��o�[M�e��b����
"[+3M3B�j�U�};�����x=sm�%�%�Oڼ�A�ū`�Gd�bZ�tN�Gjѭ��[lL>)F�e%�����G�Ҩ����CթQ��p�k��&#�����Iѷ��3�vJ<&�灿�/�ɚ9I83�+3�m��k]���h�0�S&�渨�Y3����owG$ە�v�i�gWVHh3Ls���Y"ž1׽��ĽH�=@�|״��H�J�J}Ġ��7�{�hY���T�n^fN �Sܡ17aOkl��U�|5���������`��i���Tn�����r��:[:(B��I8��;5f����x��t��#r��u���t���Rb�a#)RǷP�}�EN����u���.���}�ʎ���b���EL��Fc	�\[���CTq5�{d��.����5�S��P3I��Sh�+'�rJ>0xk�b���+u!�b���BtQ�i�u��vG]��esɇq=!S��p`�u�&䛩>�!�pZ��as^�a����F�-�;��&L[����:Sl��������8Ա�����cHX�f��4���zE����t��4|����"��	�B���lފ�2i��yZ�=���r����^��j�rp�w�Pc9Ֆ�R��ѧJ@�N����iEa����+8�vAމ��5e��������f��L���ݱ3	������ܜ�V�)l�F[�ćE��@ѣT w&��#k�ǵ{j��77����A�(.�\Ck+Ga���Gi]���S��#7b��Z�x����Kl��,�k;�N�s\����C��z{�U��f��2��}ѝ�_&k�z�	pm!j_[�@�R�xn9<0͉��qܳa�x6�����Y����r?A1��ޔz����H�Ĳz���g�V��@f��wv�'��\)^d
k�C-�.��n��c����*m������N����no����s=�BG����Xj��uH�hIxw(㉙����.����"�"]����S��@)d')�i��5�=o[�{�-{�{½��~�@��C��W�`q6&�4��
�m�o9��4�܃�Ua�I�8�Y�V�`M�T=��3���(:euvms�P�m�2�T9*v�lP3e���Du�d'�v�Ք����7Dw�Ĺ�}�bX���z�?R9�os�&vղ��+�A=��8m��9����ic;�δ�Ԕ+���ov�[rcDЊnPv�n�N%�f���������˫��4mgVôl�Y\f֮�#b���8{���mO��e�-nX7�Z���i̩�>;���.�気m��:�(j��S�rǃE�?;��r��gŬ�����W�<�M��S��+N]�����Cʵ�:��I�֥[�;wR陕}����n�.�dH����I���y�� D��ަnJ�+�:]	9СSEa���z��N
YV������Z�6�YS��lie�n��h�R2�N��X���Q\���Bz��MX��}�h#�ԺY���f�C��ծ-���o����^]Et��X1�H��_}`�P�wE��^�Ê�Ɉjc�±����"��a�+���3���,Ÿ��ǉ5�>f${:�ݘ+9�r���0r�;���9i(�{��9�aw��Ko��#ʹ�Q&jX�/�-�f�rӷ�C�(b�YXd����P�ac'f�6ޥ&�㴲]�F���mu��܎�!	s7d����hom�}L��h�|!r�.�ɵ9�U���t���hH;�c��5���BWٙ�WJJ��3S��2�4���n�B��;n�ER�y�<�(���Nң;�T�[5�Ƿ�ͼ1���C�^��x�4s��AÅܦxR�A��V3[Z�.�ţ��TQL�b�gQԇ(�V�x�W�k������xՍ#�|F*�o:buo�>k����U���W|&lE�D"��>x���9��TD�ɛ۷qذ(�ӮS����7/V��ܠVg	9e`{�o
�ý>�.�;V��7b�o|�1�L�WyO]Gg�j�Rj�|�+^����VC�݁���{�dyuYΪ��g_uT�)���2q%mmK�^�*�*�ٵ�pG�bʈ�Z�����ۥW6+]��}\,U�����ol�n��X�E|ys��Qβ8�҄s0�s��H��E��e܇I՗�D^�l�pA�6
�`̥�P��cǯ���D�b'�O�v�O�,�
��`�6�%κ��fM�7�30�5ץ*��Z#��2n&B�;˕�t���)�7)0:����4���%$��%��a�,N��$�lik�{��.��z�cʘ.���L�6�)�^�bo]z��^��>Ĳ�2x��n=�Z�;�{�����g���Ga�.=�E��1�y�Ge����@����-�v���KT�n���sb.cYͶ�{����}��ޗ_| 2�����I
�cDo.�VRB�4�ǻ�b�V��u�0��uVۿ�hѺ�9�m"�ON�Ĩ<�Ձ;yR��ؗV%�����i����Js)~vļ�{꺤�Lɍc繷w(���K�RY*�S��"�t����E�3��]	
��e��i�b�*���OJzy+�����sQ/�@���,�Ɇ���X��0t7R| ;;�]e5�P���SV�* ;���k�`�5�6���33�+sA���7d�i}3�0���[g`ﭲ]�%�����]q�X�n_r��d��0ֻ&���5̫�uq�c��0�kJwm��3Vl���͜�.��8��+U�3Zq�iq������h�2A�Qסک�{(�0����S�^J7�L���9�Κ:��qR�Y�t]8�-��f�xP�wItՙq���kr�`�r�?�B�sX�+]��{f,��'�Ӱ佥��&2K�9طK�������l�8J�k@���x{����6�솀�I%��T�F���UB�0�4������ntgM���̌U>ئ�[�9��&���p=�[Q��of��f��[�$l�����+*D���Ns��z�۠&t7]1^�l�k�gI��n�	��+�.���>�r)�a�؆���<�7�m�e(>�a�[�n$��,��(,�7�{��[������/c�%�o^W���Z��u�F�)	�ml(T�mS��'�{�����5|<%�{
�.�X�w=J�Erv:�r/`�-S}2��V���xi���kp/�]�z����,�&ۉ�횷.F�x���O���F�~S}�S�},���û{�z��a�yH;���\�`XT��V�*ù��}�" �]��.�͞�O}~���Nl�͠��pv��^��6a}�Ԧ��B��e�w���8N�����xh�eୖ�7������
ܝZ�6���P�eB�yC{_�S!iS$$��w'I�L�C{¾;|����df%�Q�y��x�j7/qWf�Q�]B����U]���.R���yq����m��|S��$��u�f�Ɏ����9�:�V�V�J�]�]��7Vz��	�� ;��Z#0��2v�/6�3������R	������D��� ���O3B�^�t���Y�ƺ�q�
iumLG��8�Tù�l�N� ��������C��Y.v.�6�k���=�Մ��pax���sX�J���7�]�=��M���ܮWB�������LG�jQc��Wx�t�d�N��޾��n�[�sT[�EeB�K��l��v��AW���:�k�@u�8����$O
��ی�2��;؆n����ʥ�������_�a�'��7�f�m��΍o3$��e��I�v��q�Vt�,�\����ٜR���L�V�Qm�k ٗ�}e탭`���^1C_}T��;�}�T�s4����pᙻZ�j��isK=�Ps�+W.�[�p��̔0�� B���I6���J�'B�|b�9�6�]OX�2���o?S�� ���^<-����C�#Y��7]��Ǣ.��J�r,U#�b�n���0�[N��Քe��U���3��/nuP�м�XyJ��A��>B��bD�.��\��0�6�F�S��R��.���e'W��;H�՘�����B�>�b{(���v�&]�<����S��!��w9� r�lb��:B�����Jw�u	;�nn+���]ީ��+���Wh���۝*��_9���.Y��q���T+xM�/a^*��Iu�O>v���U6y�;�;�gS��x���:�Э]"��6U�n:x�qSu�4.ݐ���!��"Oo�r�X�kA��L���;dЙ�xC���<i�hk�vJ�/(i�Φ.�q�K�pS�v�|���ƕ�����a�IZj#O4���mf|�`�v��oMb��팈��cy�S�h������N�o�xeE�����^���7�h�7{����v�a�3!��������U�[={Ӥ���z��%�n��Tr\{�B3��d�ë[�]�\~��8&vx,�������w/-���E�8��CX�>kf]�����CS߃u}�5��^�7O7��$�+I���6uo���>y1#���Y�H�SΜ�=����OO乸|����P�_,�כS�[ {s"+fe�G�uF���Y�����W.�P�����C�p�q�͍��+���SN�2�,�E���8���aV\�Zȭ�5��ܡ�PJ(�k�P4��p�=��jj�Z��@ũbb���r���`�����ɃT�y�M��m�`^���<�.�YI�n�.�`���V7v7!��9�䕬���-9d�E$�;�X.vl<o:���Δ�+��D�Q:"շ�Gv<�V;�k�E���dT��k��Ѕ��G�}5�O�ENz��2����t� "eE�y��L��
��5&�]q�%��W��!��ZiȻ<�}���*3����i���)����e�;���`t7��Q��+��M���I%��%	�P��S)�θ!�_\�9��p���of���c�#��2�r��^�a�kz�qY�H]�A�yU���U��Q�Z��*x]HSz��\\�C��ڔ�Y���ˡ\8�5*�ʉ�VK��8��1� �#���KV8�P�Fsy�Uj�-�%������o3�H/L���6N�G$8yI$�.��m���y���.�,>����2k��r��r��wC��j�9�:���֓
���Zb�6��hM������w眤{y��K�C��8���0hC��;���_q��|A�B��=�|�ݶW�~y��9�r�����'Ğ ;�O;x����CǮ����hC�'�_� ��ܴt����o����{�C�?�""����?�����������>?�����AE��������?G�}�������>0+��Z�b��=xA�-�l^�"c:5�K]�d��v/vx�������p�=����;J/�i9C㻔3�n���0��9Cl�W'm�U|��O��<��L��F�k7�AV��]�D���H�T���K��`��ҏ"J�q��	B�(��z�&S�vTtX\�.t�%��7��g��e��wUT���E���˒}/� j5��2Ja	��l�]]��X�n��K�bڪ��r�����d��Sˋwk8Db�Fv�Ҟ��<f������F�uE}82f�:�Ӂ��������4�ΉTx�ūl�/=���}&V��e&ݔ,��䭊�\y�Iْ�}qS�ǚz(�p��m����G�9ݥ�7Pf�{�zZ�S�ґ�����$&��pLu�r��9�
����k}}���f.�%���z e)m��p����bmT�O�Z��^M�)�X7o�n&�Noמ��}z�kޥYQ�bɞ�q�33]������]����C0�n^K-��Ki���{v���t��#{��,�0����Gu���詈�r�c�<z����b���W�ܺ�{����A����w�ö���̗�����,�-��ɷ�~�����Ԕ��y�b�v� Z۾6j#$��PVWr������w@b������d�E]\��/25my/y�w'��Y�}V9�G��KB�|�{�-�=q��η^Ǟ�>-%jͭ�M\�Y�++��段J�m�v�"z�ڳݓ2h�8h�wZc�:QZ*)�ӿ;�gH+b6�ý���q��j��h�+�[�7�:��bV���iO��	������!m^<V�3���*�t�b!)i�D��o�7��쑲O�I�ɧ�{���<O=g����^+�:��u�pO�y<P��{����*��L��C�V�jK#G����<����6b@�#�b/��o�Z�hܹ����B�L�7hw���r!���ݚ8{���WB1��oi�H���q&����Z���^9��P\��v�	w���e��9ؖ�$;&�
����W,=p9ۀU6;��<V�p�u����z99���v���l�����8�����j�,p��cƯ�p����т9Bh��]��	E�B��VP$K�Ä�=�̾Ew���݊g<�u�g�(hRi����P���L�+
�$S�!p#�N֪&�Ig�\�K^F�.O�!�oFg������sR���kG:L�Y{o�r݆<��[�C,�k��Qīt7s(�u5=k���znƺ�����<E�
��oD �8����p�u_�N��(�&Զ
����X*=t��摔�'qO�u�N��O碝�~6a��wJ�f�]�K$ՌhXTn����'JB,�!F��� �fx4@������,��F�1|�K���2x��L��"��ܚ�α�k�J���I�,538(��<F��\��՛J
�>�X���Ө��-Ըe�;+s:��<{s�����G�z{sƫ�y2!��/Ď��l���5.B��Ji0��8此ڂ��eW ��㜹R#��q?7����gбsz�8ꚼ�"�1�p�&��4����1�b�{�ȑܙ�'s��v3N- �I��7,��s����[���ˤM��u��P�%R��j(W�N�z�ݺ�!�F�y��7�4h�lz~���C�}�����g%���G�;P�ѫH�yάe,�k��ûz�<�K�q?q�B��ڮ��1)�}�³C�x\˛^4;�v���u�Y"�oW XK��g��ݴo]�;U�Zy�걭ӞV������S��k����V`���71�4�J����ʅ�8�d1�9�͛�í�xf�.�=�fS��G��
9vd�2�]�)z���b>�+���xvuj�rż!2���Z���o����^!��7-ˮ��q���z2#L���z��|Ѧ��soe��;������2 ^ɉ2����&��1)���q3݃As}�k��s�h5�"aRΠX/tl#�����&g�t��&�m�����������~2bM@��NQ3 �O	s�-��T�ax�����]��)A�K���s�PZ�p.8����(ٺ%%�3�=���%�c陼:�烖S��a˝����q�Օn�QnJ�[;$7犿x���������]eڥ��3s��s��˭�۽�:߄g�񶇄�s����ݽb��=�
}�!Nok�zn�`O^3w�"{�x��⡜/��ѧ���Qy��4�!�H�����
�����?qPŋ���^��p��I�X��)��sVf c%���tk�w�MC�\7�x't��Yvtm��)�HQ��WP��9rU��2��Ƌ�4lG�ƈ��Ⱦ�f����A���{Oک���'<�5J~��=��M|�\v�%[���rg9���N����^r0���$|����r]��O�z3�����w�v��,a��7�[�<S�D��E���w7��� .,w�;��?꽽)��e���+�]�]�S��\�2�<1"2�)^�r��9���b��ۅ�Q�?�vA������F��\���^y�\-��׻q�J��㏋�{���Xl��hB@��4U���r%0\{KS��e6BԺ3w�v^#�"�:!���-1�wx9����NzR�T��F(�b�"M�6��k��y90���#�l�l�3���:tl���N�(�։۰潮�GL�I�k<���y���&�C�,Y�=�rk=�p[L�=�S�Ff_:�q�����k�U��fLӎ�q?m�w����_uM
����v捜^�u(\O�ݬ%�&h9�ܰ���*��k@�m�{�Zk��D���Scτ��5�\�^�zsm�L�yM����ܧj4�e���t6�3cF�h^�d��x1�}���ڊ��V��d�q�5��D�8�I:&cR]vN�م�+iG���ݚN/ �է��!�^��ힳگ��Pg#�D���K�N�ǚ�;.�ϑ�gQϚ�ͷݴ����m�,˘���4���Svf]q��y�" GZ>�"z_
9����M�Ķv{��D�s��^�,Y@����gd�a����^�Fwiᖯk4��[m6�q�����c*�]��+;��Z�4q�
�u��*��}��3���%ܣg5�̆���xE�Gm.�6��5E�q�o�[��ςW&����x�yq�
ʀR�� W8�nGy��x���G���.\�I�s�*C_W��ѻ�d6��{��I�0{���t��h�֪�2�l��n�^��>���:S��䜴ޅʕ�v��Ce仔�����X�Y/�w��S}�M��e���q˕?+�J�j�gQ����
��}��#N��q:��4Q�rd��}�Jܳ�U>�;��ʵd�'  �Q����8��8�oݙ�>M�/��-�U�A]�<����m��byYԄ����G6�q�:�֬����v@�J���1	&�T/H�ڔ��5�ݻ��-*�o:��ᦑ�w���%�yï����\4�ސ,}2(�o�g2���}�;�	3x^������r���Dd!9��4;.���"e8:Z�L��z�[`�.$I�\�����*��l��7�r���V��ձDgH�kM�<�F-�gp-<�A��v��[m�S����ǻ��|�zڶ�+��Z.}Yn�|in���V���Gj�
:�wZ�2���.�|���ҹz8��͋X�"�N�R���VjȅÌ�Q��gڮ�,���޺�כ[�Î�uEs6��j�x���k�e�ks	��B�z.]T�W ��a�a��d��w\�]b�d��ў��ST�F��.�!5oo�}K
(��)�6ɧHf��9�!�V���'S����w��}�����a�Ͳ��V���^$��MԪ�\0�rܥ��;��`��}
V@�h{Y�������䕶=V]�U��*\���d�E ���,���ՀS����lQbh����v ���)�H�2������S����sg{|<�/)�L��5�	�IzxI�&��5.�N��_�2��BU���I!�݃�Ѿxϳ���A��7E���_H��B?jȽ���}�t۳��7�E�sX��b(��Q�QP���e������uuTq��X9���믭�MYQte��Wv��/�'Z;Oa5P1KX�z���"�XF���wCfZ�x�)�}�J���ޱy��3�����˞o����<��z_/�ތj��J_%���C&
���.�ز���,fhڄ��b�����9�U�ѫ�.�ܧI)v��^r��yw���C�F�Xu�A�B#!�5�آPK��	v�j$ �c�����O-BVJ8��=�.���b�#�����~�y���۴����t���j�Y�2�lW��#��N��B0�x�#,v�R:��٥��-	|���?9�$�j^��鲮ŀVq*�p��"��7��\�'�/s���:��X������f�k��4����G����kK��ә��I��%*�)絶Uk�z�vc���X&���}B0��F}IIc���V�iԿ�8���Ε�4n˕���,�1�&Q:F΢��]�D�B�c�X1��\(|�oI�)1���D|ދ�s��rY¹fhP��O76!��n���Y���m�-(t��[c'V_J��e��λ�K��uwHҷy���|��B�ޚ���D�4�!u�ִ�t���yV��gX͚J��}�f���kM��v��IgN�w>ι�tu+��^�����=�+���獇�1��,F7�x���odM}�g�c���=�"�O����)�y�k�d}��5�P�ni�\�U��7���
�L;'��k;�WP��6��:)���d��T��ti��j`�3��q��O�L�!Eݳc�E�<)˥��8�Ɣ/�e�"RE�w{ίi'��]�ݾ�7_dN�d����'�0<t���B!��ה_I��z}�IXvd(g��q�]���Hf���c9�[7����8&�q�+��Wl\Z��5�Z�(��ʮ�����M��b�1�̞��������	�Ѽ��]ZH�u�Չz�MxFx�*۟kŭ�yM�����W@ڸ>�ӤĐ�����Bʠ�NL`�{ݜN�y����}V�{��0i:*�)�ٌ��z7� ��_@˽oh���v�Y^�� ���=���s�#Ўٽv�}#;��P�af�5���z<�^tn���.�e��FO'Yu�y�BЍ��{�2�X!JYH �D+~U.�XN��\F�QS��E-}��s�� �.T�����v�L׷(��)�Z��Ç+wk��;*S�<�H�\&FG������
O�p�vJ��-<��R�LK��lWT�_Mr�*����s�Ե�5����T �scm���J���jK_��=Bɽiج��Գq]�}bjxR���� �5 } �yՋ'�?{��no��ׯ}Xʱ]�G��8���LI�(�0��}�����Z�n��)�P�$)q��v<ۨ�t�����@���=��,��7�IRs�y'CLk!��ʽ���M��ni�;�1���?lȡ���y-}o�z��*�(3��9�������W�V.�l�Ѯ�z��0�+�wq}Q{��H��+�DL8V���YΛӮ�Fr���F��9��·�Z�N�����3�Ԩ���dT��7��� ��w�u�Px-�o�8(ΟN��KT��\3&�oa�d�o{=��[�Q�dw����=�bW�9[����U���\�Q�,(g*��#��$��M������c$�gx�M���	�Aخ�q6ا�W$�7�i����G��Ms7"�#��]ޜ���t����h��9�1�f��k���̝˱1%�L�>�M)��U�P�c����G��>ǫ�G�C��,����e:9���J� �Ѳ�Z����*�����_n�Ώ���Wq��@e&$a}`�~�4m�PL��\����j��g;�ǳ��3˖�5�q�����=�=Hbn��f�q�u�c�Ö;;q���-dU��{��T�Fx�H3NӶ�������2�k]�b����Lq^��r�9}��.���,w)���{X�[^����{�+��{����@(��K�8��]�l���K�ӱ͕���=��{���j��y�ݗ�Π8��MsS��af�$�F���lSc���g�^�;�#����׎Xw}y^΋�w���z��h�\b�]!atn��V�'���`����<������%0���r�!:Y4�k:u:��]'E]��x�$�%}���`���-���$��ݚ��A�a�_S��,q�6��U�t���ػ���D�F����(\ڏ�0ľ���$,,{=�zbktz��eV[[�|g���8^3p��t՘-}�;�{iI���>�λ�/x�ľ����&�׹�#��?cg��@ �= �q{'�����F@2OF<�{����Ҫ�wf��*Y�<�^��{}f�r�Z�3���pu�w~�����=o��5��5���#��s�&qݜo"{Q��-N7><F���x��^h�QIbS\��{����=�5˗i��5��!��UpU^Ùs�6��8P�6d�L��^߷+�0��D�b�������,�:���L˕t���_>B0�_`R�g�o������ U��������_�����?s��?����g��}��o�����}>o������߀��_��s��26��~�4� ��Q�-��A�
� �`���	�6s��"�*��#�H���$���H�a�"�m��MCmBR�?�=�������GW��i�{�>xj�*�����Qxu�+��RY]��A!*E�u�Cl5V)��Lr!OIkw�z���5����f�2*�{����]IԽ?H8��:]�f�X�\��y#���zgc��h굽�)I�'n�$7��J�R��N�z�F'�8�*�
n������p��Es4l�ov$�������W���!�ü�^]3��Xz���+l}3c/�NŌ�Ȩ�N�=(��T+�iX���+�@��K疳��e?k��=ډ�5_!�e�ٞ���+ecE͘��{']�P:�Mw�I�54�y����G���&���{|�onH'K��ē���܅�|F_Pe�G���\�a��D��({м��03Qp.?S�>Qw?Q��ҙ���WU�ChD���)�3o��St*y���z2-¨+z������4�(���>���6�Hv��b/YD��c�Z�s������jJ�X}4\���ݙ'zb�.�\s)�Q;;�I����蛸��ˈ�g��m��mp���9��7�������(��:�j��<xY2���n0;��#��o0M��h.��WH\׊�&���Fw�r��zx���|����I�'��>b{��q��b7%w<W�6���u�P��igQ�e����F̃\��79���H&Ix�I�[3�SE�!d7-�A8�
4-��T���I&	@��I3��Pm4 K�)XQS�O�JD�m��E>P7
3�b���@�J#�BI2A&8!
�12NG�R��D����d QI�ZN(�MȐn(&bO�V\�M�H�AE$�i2(��,�g��<p�ڹr����-��$������������6t�DUI�F��SI��ĕT4��i]	AKQCl:�)	&�J&�j��bkMRb
JH���j�5�4:J����$))j�b���*i��*�4����ӋZ�D֨qU�ikMSE-$JD�5QE%��@REZQ)UPSSQQ���1-cf��i����u��&%6ƀ�

H�����]$�IlB�Z��9�<�CJ^�h��ij���&j��䋥"b�QK@SMPQN�U�UMAN�UR�i4�!I��S�ξ|��|��˞��H�G_2X�_J�;A�.�����O><��#���u���+@�]���Ȉ�ut�޶�j��ϮPO(k��)��jeaO$E�Ʉ�!&2����0R�Đ�I >�?BaRft�F�@bH�Ah%q0D���窟J���$�V��&�h����rQt��t瀕�s{X���{U?{��U���n�i��t��Y��u_Y��w(�^�"ȸ"��"�#�5�xϜ��7���Xg3Nꚞ��[8�Oċ�#����������[��D�U����ڽ\���ֹz��Od�WHj�3���;���h5�i��R޽W���z�o�VMS�G=Lg���m��s�#kG����_9���(ܶ�Ը�<	�熷��{���~�tլ������P�h���w�k�O��2mc�zNݩ=0��nf�6}�!���AC��wa�s��7�u}>_I=H�x��=�#�O6s���T��WO�xM��B�����,q_L8�.|+6�tŶ/�������8��G��*H��2a@kwO[7e��a�Ģ�>$��g���}�#�w8�BR7[&"/V;3/$��:#�.�BD�U�6e�Y\;2�ZR�v�]H$xkM^J�BTЯ$�ϻ	�/�J9����p��u:��1t��M�H�o�k&[z$�7�����Ru,R�L�n+�)R��������=cg���N�/��dTgSڹ�/�ʺX��G��^���u�&Ȝ����p�ė��N;}FR3]����r�V}2����%��7!^G}��Y\�Շ^}�{��+�K��A���pi�#������c�Å�=��C��㉺�le��2	�i��֏�x�����Q�IJ�fo����mnכK�1G��<[x����Z_���K/��\��r�$>�owӡ�ޱR�e�O�����oۀ�����Z�&Et_{i����>�g�A�q���6���<�1�ܛ�(��h^3횂:|�F�*%[ө�$�'�ϧ���=u���hT��䌾�K�s�'���4�6����M��u\;���||�5J�]WZ~�py�h]�h�2[{����
��\_��nz�\�X;^�I��Ɲnd�+����3� ����sY����%xf� o :��d9ê�<�]�Q���	��-L���U��ov�y�5�KH=ZD�/���b
��M���0�Y��d��nw%w[񧿫vWڡ����^�j{|���y��0b��s�������
��{�=���7�A�ͫӕC��H����=��+n�D���Ӈ3�Y����.�����n�)/ې�$��'C!�OOD�sd�a���"Nˋ��1���|7��v��r���ei{�I�"w�
;<�����'�8��6�o��8{�_yՑT8lW���w�Cqu������=s�ҪLf:�~�V�T���V�����.!6n	Mxb�<SܭH��RF���也*��].L��h���1nWx�`3��!@��N�d��]p����M����:�R���������W�4C�ꙟJ����'KԳ���?�z��3r��d��R��mX�vٗ��]c�
nǼ�Wr뺃�@_�v���mg�m]�0j(��8ZVNT�\&m w��l4@y�Fc|��v�3v�u�9�+�MqS�ߡ��4;�SNy�4��o���w�y��
�*�m���uM�(���i�x�N�1���Q!n���ڽ��3��o�Z���7�>�{�3a��M�p�f*��#��'m���E�?H����ޘ}.���ȋ��ٓXs#h�ۭ.NKq��<,��oA�;U{4�E[8���"*�y6�c������zpE�M����G�X�}�I;��'���:�P6�������9	��q�3�v�5�9^�z�N������$�q�	��:"�4A�{�9;y���Re�/l��Z����~�O�������|۹�1Y'�l���T��'��nȈ9"7������r��h�w]�s|87�f�j�+�t��<x�x>[\0��Ý�K�ɳU��v�uyK���O	�ݧ=o����&�E��_JL��~sw�{ՠ�ݦ�5�^'��d���7���q�w�^�m�KM�E�%��>���������"�g��6��,rsfT����~�4"�c���ͮ= �J�>7����ѳS�}Ӕ��_<�]J4���L��ΎVO�A��uM�L�¸�6�r���^}8t��f���u��-ՠ�{�j
��TXÈ���-�1n���ǝ�ܘ�J�fJ�vАqQQ��Q�o�7hoJ�����c�̛�B�Kʸ��ڏ��AV��G_��n�T]��(|���6�kҝmk~�$�\p�;��%��6��ep���|����K�niWu�p���5瓷m'H;$_;�	8 ws@���]0X�ǅsW~�IW\�����"W��bKݛ�����������(����<i��׽��7i=%���uC�>����\T�<r�|A�Q�4Oc�+p�Q����n��y[���;�������Ѽ`}$�ΓB��mF�VW�^�#��=��c��zP�"�	[�6΍ ��hƝ�gDe�I���M`<�'��8�]���FV����.c��m����$�ĵDM��y��YT�+ݘ��'S����u�2��~�����c�f���"H�k�c�$�2xߵ���}����pK�EǟA��{_�L1�r�h�܈��X�|���nhN��Ut�;�����z�w�_Hh��\YTg9@�>C�p�q��۔��/%���;����p_	oY��c��Y�
�twjV�e�l��+q<�й;Q��
�G�� �r�n��M�p>ND6Y=���gy��O��='��{.�V�xq����sZcIi��t|�	؀8�u����v���[��g�~��>���Sݳ� ��������ݔ�{�먙D�<�·��H�����M;��'k9p#�[]hg����^O�U��F�Ϗ<7�!�v��L�G-gC��Y�~����N�z0����;,t��Á8���V_[��%I��X�:F���홾�|��A���ѓ2����sX�T
�`?�U�,\�om|�p�H�i�3��N�]��;}��x1�ǰJ�~�e������o`nx��'w���T��z��P�k�Mer��k���)�]���y��A�J���K���+np��{�]�T�f\T�8��|A�4g����"�٧e�d�:�K���p��l}գ�졸������7x� ���Mc\���&����MSQ
n�:�c[�SuPK�~�����������w5ֵ��w�k��r�i鵏9�;w�ܥ~I$��B��ڪ��Խ�\���$a��<���� ����!��-\�n��ܝ���u�.�ccm̽g�9�=�zP7/���j�A�u�8����=8�}ۄN�_�ez���H�v�	gfV�f�m���V�����&W�b� ��������½�q��ߋ��|j/W�7���vG�=�˖4���$�<Gd��:�[-t�F����*�zx�8�P�ek�P�qu?Vz���>�����u���y�yדf��o�_V{����kN%�E��Տz���y�z�V�f�E�;�S������ǻ����{�E���R�{�x<ʞ����|C�"�PT�g||���{��v/L;�$�=�9K�6����/lߵ��g��#YW�fo�d0Гv7��\�vэzp�s�p�͒	�QR{�`^K��	LJs>�4���a���Iw�������T�xׂ��~e�C��]O*��m�1]+��_QST����\�X�N~g���.[��I��]K��_��A�.�?�*%�Mvn�E�D� ƠrU��t�ݽ�n���F��$I��.�QX�+�t������m	��=*��I􌐕K|-���^u��{d҆۩��oT�$O�;����촜�m`��}���ƹۜ��5�q7�1�5aM��%��s%u֫��ȩ���$�IˎK�d�~�do�}*�ڂ������xb���!�\�PIج���W\"w{D�DL�SUS�3T{���q�}��@������c��!V<����}4�/R_��|o���ۉÙ�wE�5�@��i�f��KX�������'�;�Z�y�'���[ϼ�����2	�nګ4�"���j��w9^��M�b����J�\2��̎�[x�i�l���Uw#f�Ϫ���o�O���s�.����ƫ>�R��y��Mx&�=D��ګ��nh.�"��v��p��<x����9���/V����z{X>�)�|��F�c}^�,>�q��R�v	^bS�����L��ݹ�<��_yz�c�Z]�@�k�~���&��v��G���7ٞg1�*��>���fT�p���q�Իޥ�`O���vi��G�&��o�,֘A�ߩ�_j��T���X�^�d����*�YI�����9�<��^�6���C��w����5���ߚ��5b\6��Գ���6 ��aϴ]I\`yWWqI�t/��u6���,�N�aDY&(�1���=�.��[\0����_���w��d�ڞ��OaӚ����P~��=7�̕G�*�M�=�_eJUO��(�/�]zwMo�/��K»�(���t�ms����c�FO��m3TM�RەwY��of�ҽ[�z��k�*�I�����I^��x�����u�nq�ֺ���R^�W�<@X<�Y[_;bMn�����%đ�d;�r5eP|��a����;v����Û�|�~��wqoX��!WC���Ϩln����A$F�hb���s:0�h��옙�#)�U�Mb��cS�r����.��:�I��OҵUw�4x�b��W�����G@�%6��R��,��ī;4��r��}F�׉�i��fz�m�Ds��4��^��f)2)�!�l���,��&P��,��ѳ�Γ��=&��og��
��7l�{Y�.jik��H+�呦;�G�>����6��D�\��㱒�o-��Zg��&[��+��2$	l��^��a��(6L�R�tC"y�v{��U:A�'C}���x�^�kYf����>�*\�ʆ�Ԑl����N��Gl|��:�� m��H&��LЇl��#�qr�g�{W9P]ƒ�7�����WvJ���f����3���el�[��7�eZ��O���L��@m�.lf8����N��M���,��E�;��u7^|=[,�<Z\�G��w����힖�%�"����">��E���\��+L?���&�̛;d�O�}��^�6[�nj��7[Ɲ,��Y�*60w�!�~��o̝���I�O<�վnf��g����K�Y���8�G_���8h���g�X�XaO�6@ɜ5��h99ݦ�q�3�-/�3}5`���z��1^�>c~ hҸo0�y�c.Y�����s��'�X���d?
��"�d�oF��;�7X�tg��88z�Os�ވ�uin6��λP�h(-X��8H�m���]����q��@���z}��?��x��������g�������}~oXF��S.������Z$�J�Vg�����4��̎�A��Z��^
[F1�x�i!u�1�����zM��Ns�y�9A%�WD��el���7�m�AU�GG����N�z@-W�{<
E���e�->����5b�ҽ��^p�\aم��;����_��A��fgH�ĉ�M�Z�<X�d7�,Y��8��v"O��h<h�\/w�)�L�R�EM����~g�Ł!�=�9b�sB휂-���#L�9�kA����zv��=�,� š�8M�]��^����a.���y�yr�(��!�9��,��|��ӺŨ�<���z�o`�%5�9X ��k��N�Vt����C{�nr�����}I�����|��bm�of�_Y\ɾ�܅��ۡ'�Z7�S�)�%�7��c���p�:��J&����w&>��ֱ%��D��&�|�!���zy��iٌ�*N�9�{mKKKr�����Ȧl�U��M�1#�&��glQ��{x���U��h*n�)6���]����l�!0�b�JR���u6�):��ꌍ�u<�y��I��2��k�'�,�+[j�˷J�&��ܾAլ��ȊU���^�S�<�jg\E8��$��;wt�45�@�܊V���4`�ﵼ��x�nMa��'�͕s�٫��H*˖�]���n�U��c�d$���+�8�tQsB)�ʟ-����cÝ@��ߊ��y	˃Ef�}Y��K�5bN��ﱝ������{����}7�f��%��ő���Cѷ1��4�~V{ˡ�ߧ<Qj�@��^��I�{��q�yA�Pp��O�0m����4�wst����8��2Y��5�=���95�?yHp�H��R���|�S3����!k��S���̧���Q��"$����˖�a���Ow���6m�W�P4�j뒳��_ʇ��h!�e��Ό�rQ�t�<��;}�Z�M��t�7��)�.a;��6�������p�i)�W^��C����7XU�hGw��1a5]��	֛e��4_	����f���O�$��&��w;�� �R���N��9[y�y{����
8R�O�J+�1��6#E#��7vǁel<h��V^�h����z޼�\�g�Vq������6�m��@6�w�8� ތ�)93F�2t�ٻR�V_=�ė	pC�-�� ��t��7޾���� ��ݹF�~�C蓱���� XÝ��=[ɢ���ѧ"���hFaP���w��Sl�l�#ǇǆK	�V)�
�,Z�ݠ�)����B�UI�y�xv�v-����S�=PYhя�ݱ]�2�}D\�.�o|7����\W�f�[��� �)����&į�xvo|���w��@oe˺�m4e������ߏ_�|�}8}�PST�4�QE�GɱIKAF�%-Q�%$@LĚM5@QUI��M0L΍5C�BTDE�ƀ�j ��Y������������������
V����*� �!�hh(i�*��
ZV�"���d���l�7.�ֹ6�C\�i�q4Q�`�*�,m:�gI,SkA���\��5��5ʹj`�I���L�&�39$�Ma��M�I��Y'T�g�ɸ�hgh��A��-���s�1M�Y�l�hkSS���hy����ʹ��S6�+S�*�O"��X��Uhq���F��O9�&s$Aˎ�S��Z�h9&���m�9̧$l�O2s���ۜy�A�ص���ρ��|�m<�mi�1��%,���B7ML���]j��'(�Ǳ%Z(ێfU�\O~�_VFZu�3�R-��F׾ߩ����!�s8���� yA�^���q��F�cn�$>�hON�<_Cz��6"����,��I�i�K��/�;�hE��	�C�"�:����M���lǰ�4���A+��!c��p��I��$Ǹ�^�����6��xS�;z֖��Nn�}<���5%LۆeJ)�`8Bqk�%�W7���B�p�NC����N��-�Ò�o��m�]��~5'�}���͓�8����r1�6�QH����(�s�1l4�ǫz���-��xA@����D_�һd�D�U9\�2�ۄp�����=�#4����#��s�;y4�=0���$>Q%ٱ�41y������z���M&T�=�	rO=?D�U�b):�g��I����<���Ǯ�f�&�i�n�d`��Y�,�SȾ�o=�a��Q�����r�[ȥAm�F�)�by(�˵Oy���^~L ��
<���mLpm��iNqD19	�^�(���̤�9��}�댢ۛ�j�vC��^�qK׳DM߿@�;#�ߖ��Bl����;&��g*���/�<����ꭄ�!�{�FF��x��nU�u�&����3#��z���k�;�s�;y���$(�5o.U���U�[�e�\Ԡ4x�ҏ�J#+x����w� {��DF��]>�V;���f��粕:�镛����9�v�1��;vvV�B�?f?I�n��K�t��I�wk��(��5��.?q���w���r���>���7�`-�S߶=���W��~�ɪP�O�T����t~���1�o(�{`����g '�s�uC�&��+S����L
g������z��Es�����}�qG��zؚz��k��tld!��=	�r�mgՆ�pm9�a^��;h��b�-�h/a�Üv�m��}�K]����jY���>3����8��ԍd����N���.��]� q���i��w����n�����o��%�q�5�&
u�*q��lu�5&Y��g��yf_,5�0X�V&�)@,�����ު�6���`�~+vyIO�ۊY�7�/w&�XgOe��\yo��A����X5��¨f͗_d)��IX��6��yo���l`�Q�oL�pz�#�*(j�'�:�'����V3ю�ơ�j�3:
���?+�/䠳�t���<����b�ėw`zu�=9���2Ǳ�):�1��qi��S�M����=y�^tF��຋�o8���f��O/
2��KsU��s�����WV�܋����FҹӅk��3i�®�u�tv�$$�2	�������3���P[N�K�U�BOR�if^��v�ݳf�����|�a�YJd��:�W�%n;M/�?��@t��y%�o�7�k�L�uNj@��@�󷰛k��z�Y�H����	�r�	�$hZ�*��[{��&�o��b�u�:�0T�h5���<~��xլ��Fb�i�.r�{�]��\��T_c�;C{�K��μ���krD���y�����s��	eC��0О��Vյ� Du-礔�l��@��!o<��t�"x�X�����r�R����[��D_4eF_V�m�B+p����L*�J疯Z�I��RXבڈ�	D�{�Z� �� ??W>lP����F�ֺt6��Ay�f���J�¿k���������Zx�_�@=*5�|�2㷺�#��652���dRJ%k����{*	{k� s	hN�/*�q
���-Hw�����3�`����6��m{��jy'��<O`����n�;�+Vd�}��W�����CƠ[x�j��.�8!0���~��vI��K0'r�xEbLφ�G+˭��X�8�;$e�u�q�v��-�sW��TI�bhY�O����y}��}��kި=�u}_p����?_8������0k�TR�j�M�c�1�����,I��=��_-��{G3b���:�Z=@иA���ӭ-������U:������� ��.ءU�؎�(E�n�kK�P��۱�|=��kJ�OP�Yvb�C�2	A(�2\�]���e�sq,u�5�`0&P�. n�Ch���"*��D�n�7�����_�cFdrW�Az*�!\�_[I��P�� #�m��5I�:5�Y�5�X$ˉS�W�2�Һp�鱬q�^���T�Z������٤��O+��ׯ���´�0��S<��%6��~l�8�v����l�s7	�0hФ�E����q%���7$v�����t5��i��Ђ�i�q$>P�		��x��Q�܄&-昔���SJm���2��
���B*��l�=}Ǆ���C�`!:A��!<�4սyܬr��P�g{��D����	r�ĲN�7E2J|i0��og@���O\�����&�0V���ݹA��fG����ZL6�l��{E�}�]0�#R���eAi�n��r����L��n�G��Ί]w�S60
,Al�� �4(��$ڝ���_X���L?0	�8p/n�,��3WQ635�ک�?�y�1i�ƶ����8��a9B��ˁB�w9��C��o7�o]])&v��[B�*m�&�7U�#��:)x��7�`���*�7&��><�_����'�)�R��Ǵ]`�w�ev�Y���W_+��d�%'*��Ъ����=ũ-���Rl��ys���#5��;}֮Ay��{�*����{�ݹ�v�1��  �+�b7*][!�Z\=�>B5��?�Ý~ىmZ:����	V��zO�@8T���L��Y�_�zT�a}u$�tY��t@�0��dd�;���J��?f�Q�³��aGk{��L����<�������fy��31a�v2`3?�h�^G	����H���jv�&�˹˲�U���r�*�f���_��zH~,�|LP���ź����x9o	0�촫��v��zvk����j3\��q��Fi�!�����z��yh�������Kqٔ�B�v�4�go ��KH��Z@��I�uE����CZFnf���ë�]+ܤ��4)�\>wcY{Ku��-V�.�8Y_���_��qx��N[��jlԕ3i�A�{��FI���m\5qw:ڶ�r��l�=�V�ht�vx����,:/1q��^UX���P�E�	l��*�e����=��
��Z2'�Fq��|��[�{lw������M0�� �@����f��{��sK3Q�Hprgy�zN(Q,��Ji��(�7m�����R��.1������~��_�w� ���-t^�H#�o�.Ӓ����&���MWu�L?L�`��+����Yϥ�M'�U�\�؅�E�=%n����e���+���#/k��D}�_KA���!�;m�S��N\;0��T��}�>���&�r�񎵻ϽP6�gf~����񞥥�R���vl��	��� ��O8�	�~1�г�ȶT�Mmb:癱�7�u۞�������7Og�%٭�� ͪa3},�O�d�q=�i'b�hNO7�����8�6#������o;U�`��R�1��"�@A�:[hLpm�{<�Qs�!�d3Ҩqms_^��g2���SWg����^K�B�f������-��0Q��^��c��+���^w��g��3No�L]�Mq��5��	�Ͱ�L/%��t�9�D?�X�]���~]��\�1�JCL�y:���Ku��TV�c���׈ɷ��z<je�(�wf�� �"�@xzql���A�s�jsM6��u�\��BՅ�ux�e�~����5�@ףp8�r�	�5�����1D2)�渨:�3��-���鳞��:}���GP�I87��i�{�y�v��sQ~�y7g&TT��mM��!�9PT}�,��&T&~��[�ޠ�O��-���� �]�XfI�={i�{�����?
��P�)i�}�D�GE�6D�N�uN6ۜ���2����綷￿o�fß˯~�5w'��S���h�{��3EVUl���{�%�=n_���z��N{��Q��:����}�2�c��[V�<�wW�70�'�_���y�
�8��5Yƫ2�su��^�ueZ�ib�S���־��U������ "P�N<{�����{����<|��s�|�M�Q4���؇�#��gA��h�ְ����~͂�x<�~�}�
O«'�_��
��Ɵތ���}|+3�q����[���ɢj !��z͛e�)�>zw�X03��`%G=w�ѓ��	�mT^��zf�w\�V{�A	���g��=�T	eA.�g� v>5eEÚ��A��!���d %��wFk+j�$"q���v�^�XϮ�Ź� ���tF#B�ʢ�d� \N^Эӌ��}J.�/4�U��
1�x�	��]za'`$^�7	�����	�{��#>��l�hQ0���V�����r�ql�+�f�Od[
�N7���i鄃��M�k��f���Θn�R�7�H[��K�%͐��"���<�סĚ�ũ�-��n@��i�'� �y�,��Z����Svb��:Z��0�JOEE2.�8�9��zk���3�kj?�ןC����8~DN�5��!\��m�ʅgl��%s�P�r���),�#�;���X4(+w�������/���s��j��q�Dd��R�׭7�p�l9���%QaV���3t�Xo���B��8��H���VڋG[J�f��"����iϰ������5�;,��h�9�Ci���C[��ʩ͓��b�̈I�ݼ�X��^o.���Y�c��o]̣�)V4�J��vÏ�u�[ھ|�3e�ڛSq^��DQuҌ������]���i���������{���ｺTZ�❟H`�,y�q�X�����4-Z�k��_�s�PK�r����̧�Z:pL%=rJ����#�5!�bՄ����������m@	��;h�森�#���WVΔ��
2�'W��r��zw�6����B����;xɁ.��ƈL <F���9.�:��,��������iWMp��:��N��u�2�>:"�׺���k˼xL��ݡ>7�L=�l���XsC�pj�Tݨ#N�3"�x�� ��$������!�:��[��J�R���ys�Q�~u�{(��E��_�c��-��Ar��F��n6�5t�æ�{�������f5��/o
���#����Sઌ`+�NT��{J����aV�D���÷�n��Od��f')S�b���{��������C�\8�v��q��ږ��%0|�&M�$�݌%�F�<7:��� y��Ȯ��{i����vH�	N$�ʘS��^!�v)���;���7q��Z#�xp���r�x��~*Kx&���л���V�PmbP�,�M��1�Bp+���E�������WsQ[��S�|!��kY�(�\�TN�#�y0f�*�d�5�K���U��]��u��KWo[b^���:��hӦY"(�Y2��{�]�\h<>P�����7�v���m�ԡ�G��h�ݰ��@q8x��'��ev����Z��`D�s��{���ݜ]��CW1a3�̤�
�-�����ߩ�@.�/��w0�ZbA�lo]�,�\�=�MC�f�b��9۫�Xg:�A�c@��h�#�(�ah�]9O����yt�� u ��7q�"�_��9����Oa 쐨f֟A���`&�4(��P�⮗�j ��n�Ab�. e��ң����>\[�sP���0r���[�ji:�3�T�Ԣ�`K��ը�s/�vj�&.M��C��UV>��c!�N=#�C�G0���0e�׵4ڬo]��M�S��jCa�}�b��q�VW;n�p�����()�^�_�\d�}��] =>ØO����L�L��cү}{W2��+W�KX����S��N��5x�K1�a��p�^�`<h�\�U�t)�9P��x=M���]OC�5�!�d_I/����!�@�b���b���z%�>�f�}�S��K������@���}�i��Q���dn��۹��Z�&����q�ؚ�qJ��id��M�Sh"6]B��ĕ#�e��dB�ڮ��Vw������іe�O�KI]��<�?�07*��.�VU�=JE�nh���q�M��#�#6�/^�P;r#g32�7Ch�6��T������FE�h�/Xds����d�ؼ��uݕ�$'W-ݍ����K#���"�n��7�oL��I��{��C)~̶ɽʎ�����E�3����AKuˋ���5B�������3�)z�T�r�?w�Y�~�N��k.�ws����^mGke�����NPz͜OX�o
�H�x����Eǧ�]&��o�â��c �f��zB�W���րJPd֌J~Tx�0�ј�oV�^�������%���#��繥����n"�tǱ�
�5�^~����=���+�i5�>ņ�Y_�
V�z�:��_�Lr+Hwk�t

'����0R/��+�Ğ~1)�|�R�i�7�8�\
4��G\� �6�ד�}��%f>����@�f�}�f���7���K0S���R�4��ߦӕ��*����4��wQ���s3����Z��S�0���TG�d��@A���?�E�sQ{��t�.�(�rpG4Pb3_�2�k��S�����i�K=��l��h�#�N�K.{� Ss{j���TS�KI�s��]▤6	x�21���?y>;���"�t�~��F���_~f���M��-��(SkA��Rb�+6�OH�T#�[_t$���o7J}�Y�� �v�x}r,t�������~ǯ����?c��������{}>>>�_�����6e�1��,7��+&�=����٠�)�D7�!�;-��D��B�F;4��Z�u6f�L��ˊ���7e4
6T��ծ���<%��pFyG��8��JJ�i�M���. d�����9��݌��[�xk��$=�)�j�gPٮpεr]����[���I��3�͝�^J-��M���b�߮kV?	�J����P��}���)�'M���� �ƅj;�̶{C��{��W�M7���x�����RB�k�?lP���ym����ڰ�^��Z��K`(c�Ꮍn����s�7\��J	�Hy�.yF�+i	ֱ7W��k����X�LV�d�:M����y�W�q&�x��z���D���!���)me�Į���dz=�y�ÒVZw��u;����y��.�Nd��.|������ur���s�R�c�]�*Ȩ�R�]��]'�D���34|^���vE=��~�z�4W��>)k���ؾ,�QL9owm�d6GFz�8�4tNgGV���p6�����ض'�`G5u�'}��d��`�E��L{f{�����~i�?_g��&<ވ�۬\�<,�n�Q�/
�
��3k�I��R�^^���G`&A�������Z����oV��0����(���ۍ�<�9��/�Ud�I��;-1G|��j�v��,z�y]ǚ(��۹��,�aͥz��w����o��k��N�V�t�l��9:v�O�77� H]s�6_���&���K{�L��ߓ']M�������'�<+���.��WU�w`�����x,yc尺����۾�/�`,s�S~���&�.`M�-A&:�{�0Ǆb��ز�CH�LY���[���r�^9*5w�Y��}ގ��C�f *�mq4(h�� ���z���l�[-F�^��V�X��̧n��Z��S)+®��!\۫l1�?[�P�ޱ}2�(ͭ(�U噊�vP"[������[AlMG���2;w�X�i�ȫ��N��-�(M�{N�ܹ�0���2�&�����f�.9��������܈����&{�� �J�0�%e	x��]�G��oS�9V:�����ǫCE�o �o�ٖziΉ�d�q�tc�tu`�}�}��8r�7��o$��hL)3�J�Ƭ�5-�u��t:;�x��B���
�f�q~甅b��63&y�����ͶC���.�n���H�Ļaw�NŤG�n��gLxfj{�]���M�6⮼�Zdt�Օ$v0AF���靖��&7�����!�6�"�͠���|�K=ZY��N[��$Y+8��T�*���n\�:�gM�}B�K66�QlM�N��v6w��]S�C1��Զ��w�$��A臹yW�=��On�M��4��}tx�z`S9_�"}/4�6��U�������w�	��h~�~3;��k_��ճ����M'��]4֓Z9/'Z)��H��+O6ykF&��H:M�#�
*��)
����LԺHEB��5sk�T�h�)i^N�@i���l�&�\�@r�P�Ul��l�DAHҔD�E6JF���!j��KCli��5��)�8��+�4�9�UQ%&��u@i5MQ%IG�LKHP1�@^0���(��)
R��Z����$
Қ"b
J�h���(��
i���_#���_%/�����$�F@Q|D�3��� �l�J�x���K
�Y�յ�56��:�ţgc&����iuj�C�,��"�Z��ba';����y۝,|�)M%
q��a�!M�b���B#`��)B�,B�`��������=�<<<�����o��ql�WV**�,00�-�z� ����c�-�C��YOޔ��/�^��Wy��_p?�uv���޻Ub�,ބ*�\�X���XO�_tgՆ��@9��4��@��`;���W���(cR�S�!oa�@׆xBgh� �"ac��ԍd�oP~y;��P�f��q�O�Y;�����e�)�Y�9�I�_�)�lwЃ�C@.9�&u��NxoH�D5�B/0��]���<�u3Li����1�&]�����m��ȧx	A�Ų.��šɉێ�W����׻���Ƭ0�q@Y�5�Pj(�f͗_d)��IX�~�U���۳����J���^��b�]NH=`NE[W(!>��� �z�	eA.�g�c����xm�C�zJv�C;��mm�*&L6��pP2|,D󌩉�i���3�v�A������F�+�����=s���if��m:�^����� �����'l��p��M�^~��=�b%:o\W�l9@ס�k��Ø�Bu*��a��Y>�x_��a����ƿ~F���l'������G�mz�f~NPg'�x�&��>*o������4�ׁ��;�&Q�J׌��wl�%�͞�n�/'g�,���>�K�򦦈�9���.c$旌\�$���9���3ج��߷�l]�G0�D�6��j"2:�k����� ���y��+�E*!�����-�Z��"hӅ�;�0��<��0�'�W� ����zn�\u��m��Z�)���<��S�*m���09����=5ʒ�J
�z�g�;%�ǾK��k��hk熂�Nϓ
Ge0�p�啫���n||��hj'q,WU\�h�]"n�l�MT`X���"d^��� ٬�f���d�,(]<�eN����T[�کLZ�tt�9"���r�������0rŦ�ƺ�sm�^�(���9���_BOlE_�v%2�9z�5K\îD[!�a�O��f���9ͩf[]�XsQԨ[ZSDft�R�]
�y�]NJ�I�`9�ǠYr�Ɂ�8!0�#m����d�L�wtn�(�k�]���8V&n�g!��J/�����G�g�ŕ��}�y�#Da}Y�'���l�y�k�GtOKrr��⠶�ާa����{�|	I@A�vÂ-�<S����;�^�!���N��{�ʛG!h���	�(��E��_�c|/ ����At���4���M��l�}�Q�x�"���Z�
��Vm�p��Ȫ3lY�	��X�~�D$K�Ni��-�7��o��G꽖3����W�]N��Ms�q"�r���p��Dp#w8�Jug$�WqH����U��;�wاd����
�4�S{�2ٛ�Ӂ�l����{�� {������0 y��^T� n^aμ���9�K�����U���ʖ��ޥ!s�� ʭ]7���YHB����n��B�q���?XئxAll坃� �q��NԷ5?)��<L�U:���k"�lG�N�OnP�������,xs����c�V�pc@�A��l��W��B|��t ��\c34�s��7�gEH���ǯk�<'�ZĢBa�������Mˬ�U6stϠ��ah nGt�N��d�8�,��&�\��s)���֑2XV�S*�i�òpRf.��۩�F�58�$��~ǒ醄jQu��L��MCu�r�q��P�˙�gf�����mt9h���4���`��"I�P�O��]/i�?7%�ڸL�;騵�=��(^(��V�\<P|�^d�����^ͷe�	���	�d�2�l���r�f��tD�M�m�	�̡J�/K s����#Xt��=í~����`L��F��C�A�4�er���K�J׿%���'��u	�TB��c���t����������pv7S44l�_TEΏF<V�lF�fյr�Gj�
��� �/�UGx��o�����Yǻ�<>%�[�M�z�$w�����:�
{k���.��%���޳w��ϣ�F�u�O5ے�~�*���㓊~�6�a������xx �ڹ(t�ޱ3W?�wM�0�1L�/�r^�W=�2Z�d�*
,3�.����  w����L���wd�����C�u�s����d3l��Q~�^=$=-��D��N��-]b�s�x��-f.��?n�ph��xܺ�l hu�$D������ƃ������Hz���e��{�U��
�_;n�Omb�cR�S�
��sCbY��G4���@i��=uE���oP֜�4�4���veL;C8�D �� ���<�}y6_�)3cT*�����R��U>���,V�ߠ���Q�6c��{8�Z�R��8�5y#�6->���P������8���Ǘ�6,6:�;}Qԃ�aܥEzt�)�є5���(�0�ј�oV�ʭbL43j��]�E����T�G�-�ې8=��'�A8oP�2�=�?Mr�L��v,49YM^Ed�x���b;�]Mtq�pP:|2%;6P�L�� ��<��S�����E0
��ɭ�^�I����J���Ŭ��R��u��@0�m#Д�l?Y|ޗi�*�$vQ���'*��"�`�mqr�f�����y�l@4�ޠ�EJ�'���E��s�*��qt���؃"���>�.ߛ��czC�5u��׽�lQ�0]�X�K����uлx�n*���|���>�vpoL�*uMYd�J�q�s�sݳns��e��u| ���������(Ҵ�Ҁ�>�w�[^����y�j1�@:k�o
��'�-�tZ���8^ޣϡ3� !� �M�&86ȝ���)�Z+�"!M;wV9�|Z��p�Z�.��Y~!@%����bXa��{`l0Q�>�#�N�2���{�決D����5����T�Uk]��^jԍ>�C�;��!���R<�E1�;�ܙ����.eX�w!�f�����F��cB	�kX�x�Ǭ�>�S,�\�"vk �K�ի:]Wd��n�$��?��D��X:�����mC#�V������j+��<��іא����QԀm�z�ˁ�P΀�`������r����OC��M�i'�s4�۴g�S[z���^�H�����x����/��B9AP4Gpyx؉��v`k$F��w7���'�]��Վ�'�d�ni��I�_�)��ȗx�!�E�4�&u~�m�1]q�u���+H��z�;7b//?g��5_zs��V�6s��g5��ڏVȤ��ϐ�aW[2 ڵ��T�J-z��º�b��b����2j*��Q�+6(��jyR^����^*��������\z���}&��!��lcg:#z�޻��\��)kt�̘GR`��nd���غD��x��KA~sK��[��=�{�r�'7h�P�ٲW
O/���6hpx�s�7���[����3����d�+[�vC�7��������7��
���̩�r��y�>c�
7#M�ȫjT�Z��A=��&zǽ�`�?V�&=շڸ������V����{��r,D󌇎v�.�d���T��S��Х)N��;��6P��>�q�q����x��q�6����� ��A�k�0���3p����	�r�cK]5��|[Va���="�*��]�M��vE�*����zA�" �؆W[,��k��*���5_(eƕ&X@LU�y��䉠_���[�	��A�v!?Nf��v���+�^L6! ��K�5}^;uI��Ͳ.�q��[�#h{��R\W)� ��ӄ4nO�v�^WG���E�C�c�^��sSƅi0�9+�Z�\��iIb��0Оً�=S���y��K��*��0��rl�� ���ίƲ��d�6bUE�z�O1��Z�e3���6�ݪ��:�Wa�������k��?1��Z`��6:�su�B�xX�l-w�4(>�2Ü'���{W�����=8+	t�#��� F�4����f[^�Ø���[��O��F�Ǌ��\'�% |/���5��/��ٹCњg��5z�ݥiQ}*�N)�|���,=ɽ�+�3��~�L�*�|5<�=�|��8Μ���g�j�=B��E��$|�~���-�;�zg�VWVK�LU�(�{���>u�^�<{޹�}��
�*���}w�cH�q������:N���KsQ�^��W���>a=�7���NI����^�g]Ig���iڹ�{��);�XW��.�8˱ׯf]��-�tg/>ה��@���D�53<�g�Z���$c`�nq���v���tC�J�öx��e^�xb:�c�;������,!d�"�,q"3%'�U�m~݌k�&��M�z/^J�!^�k��5G4�ra�`���L�#,��Y1��[�#�G��)Ĉ��/b�1��&��!k�A���j~�z�	"�PZm��%�%G\={za�e�^�����p��?�|�����v���{P� �G6�++�T��k���`�hФ�%vP��u������Ё�i8�!�@�b����2F�m�=��z�n���ƲP���e�Rv���S�[�l�*ո���(����֥ۡ�M����p�<�"����k���2���Y'X�ʐL&�����M>{3����8�m�f�r�s��A�GcH�W�]�(�ao�/��(���`�����XԚ�*��V��䬋gD뼋h��{\����S��;�	����X�9�Y����k�f�ެf��p`LQ�M�����s-	�74D��R��l��偘Ml\׳=��uhx��y�ۜ'%'\UGk
ʫ��uvh{�����f P��@�J(
"A�����V.���^+��fo�p��0͑�+�Jcs�����B��v�?�P8|���\Z~b�V��IlR��	�[bJz2a���XG�̛Z�#[�mMV���	�+!�VC(O�1�#+Z�kp}���%	9��w=,��Z\=�!�!�@�p�_�bZ�I+������ؾ�E��Z�[k�8�ҵ��+����댝���]�k�0�yE$�L��umD�Q�Zr=��z�˰eRb��_7ܧӯ@��c��A��g�3O���P�p�cZ��~��C�p���5�Y;	�����~]⾏�w�mx��HD[yn�f��q��ڞ�7cKh���Nؽq.�� ��q#�*l��Fk���3�X��{���Š����ĕ�n�d�k��FbvUލ����D�̙dzT-�Qx���6���n��$��Ҹ�|~B?�s�7�N�a�U��D�w>��O���5�,G4���4�FS���s�C�z�EN�}ɥ��څ_+l$�6 �PeB��ԑ�Y�����P"��0��a�{�g
�A���N�U�٭�茑���4_�J����^�R��q��,�[�������l^���,��ˎhQc� ȌM�Ե��>�7=���-b�X��L7�Ch����z9h����ҼJ}"��#w���w�f1�|z��Ǟy�|��|�׍���
� P@%4���ϯ[ϯ�ao	�h���w�"j�XB��`z��W���M��R��ND�aG�1��[��:�RU���bh�9�l%��á!ç��s���R�z��A8�G�L��p��!M\";.�7bRe��Ӯ�c�Ӓ�?��H��E��`�_	v/J/�bi�|"S��S%C�m�O'����ɟ�ONb�,��s�A�.WG��ki���k�c�H��`�vI���4��ݐ�'K��˾�˟"�I~�Ȯ�v�j���y�XE����D&�w#�K��f��A��yi܊<��x��C�&R�TZ~XH%��܌�����'`����T$��
R+D���޵51H�������Zn��~Sn�B��Pk�	Sl�r��iș�����+�t!�*T(��X���t����FM�؟�埣`l�I��9q��ǰ��+�:��d���*",'�"��.�yoa�I(�è��:���7>��Q\�L�/�����Iꍤ��*�?�P�k����d�!LZD>���t�C8Ў�)8$~^�B�����z�c�O=(-ᨐ�.6�؟�k���F�P'�v��p�
���ׅ�&n��-�/���|C�0��V�Lo@.�c[	Ѯ�Z-��8��Rˤ$���i�/�\�e������:�~ս�VR��ӵ�K����=;o]�P�s�{S���<?7�<0�h�JP�R��O\��ﮂ�l;;�p��k�	��F���Ai���lmH�J��A��N�Tζ��m�]�D!�k]��b�_��:"��<�����(8����DL$�"���S�>�f�㴔�CW>�U�K4��<�4se�C����U�mG��IFz��/B[�*;����/�u��\���b���A�0�&*�+��"�!�-�<���'j`���hFI�l%��S�:�!'�|Ǧ3r�9mZ�����	�8�Z��t�n=��I�P��y�z��+/머[W ���.�`��v����v����2ǾQI�ֻ3�Q�	����w�<��,)�\[g�T\:��|�� (2�p�;g�e����)��4WN�LWQO|2�B�X�$�dRS<\S�S�Ы�8މF4�t���2���)$��	��{���Yz�n?3 ؔCoI���0�S�D�78]�)ᅍ�F2�1����[2+�$7G;r�o�����egUCIʔ���8Ⱥ�7 ��F��vng�������x��}=z�}��o�������������~�rpW����5ȭ�wא��p�A�v+O/�����]����RL��������X���ҹ�Kz�u7Cj��N��R��W-�ۧ]��3z�:���r�G���hѮe=Y�1$6�*��~�ڵ��:y�4�Z.��V�.���u@,"�<�
nO�3H�Z�[�1;l⛼���ð]j�dD�ۭ�nH�,�t�59��9��l�}�т˚ا�c�����ÞO6�!�)Z�M�����8%X�\��D�؍f�p\�^�B3;���F�����+��zN�=Z�'g�%y\��@�y���\P)�c�mݙ��>\G�L��(T<��g/����"v�WaHi,���8�d}t��KR�g�#K��[YV��׃��v�o������2�{���γG%��|��3h䦰���s&LM�Ր�P�C�)Mͳs��y�K�<!���nu�(n�NOcz8$����΃��R�+-��.6C7�/]Ԥ��C�z����e<ޙ)�4����p��'�|��[챢�{�;T�Z��\5������)�M.����]@��_a`�� ��}s(����l�f^o:0���I�n��B%\�0wq�t:��0&���1	e�-��.�2͛=��T�=>v��;	�F��5�!���e2ܻ�1;�a��rh�Fl���X}ݓ]^^�P%�\D�K1����hL� �l&�xJUA�{��FR����܂�����s�C��+D��n�e:��R�.��.�W��b6����{�ن�L��]~ L9��ћ˄ڰ&Ta�\�yJk�������R�}�	ȫ�Q��%�ν�(Ew�;�[.��8�+&�&���k�������|}q��m%0����Ӄ9�qr�4թ�����f׭j/>�x1�N�Zo�����f��$k/����5*�o��,ջɊ��]�u=reԳ���ɪn��,=hur�&��O�v�h���w9�{f�[s}�W�=3oC����;^N���y�x��������ofnU��3i�ק����:�D����e�L:�kq^��T:f�;J�yI�q)���Dx�x�&��ѥ�I�9xvI�[���c��k�a}-�*�c��eHEf�ҝ�[V�m����7�mnhW�z��cq���2��2M���.��̾W��-r���%JT�B��[�a��A��0���M��˚��������Ӹ�`h�vv��%����E|s��hW�۸1���OU}�b�7¥7I�G��@��n�]�r��j7�6 ۩LR�db��n�*�����l���
�2��U����÷��%������9P��@q���w?z_WY$�ɶ�a�,�}2\�	p���Z\��İ;��I�̸̃� 3�f���R�������z>5�}|�$�j����("j�(&��������(*�&�ɡ���
��"��"������ (h&4���h"j��(*$�)R
�h��6�R�$|m%U#T��@QM�4-%0:/9�4���h1RPS3�C��XԱ%R�PV�%P�9zےh��r�h�
<��j6����h�%�4��ڨ�2s���I��l��j�'���ڊ)M.�1;e�����SZm�*�i5���ͧAI��qh
�#��ǟ��D&��Һ.��w�͌�O\�{��a��gά.�S����v!�&IΆ��j��ǫ5l���nG���J��}U���- P%*��*9���:ROU��V���\�П�Ol�&�%s�P�r�ͥ%�;0����=ޕ#5\�I�s�ಜ�K��jP^/���"n/^��Ve7�2u��*�
����1�q=IZ�3)�jK�L5�B��j��A��i��O�����T�^�4-'��;�lS<�tb̫l~�"sS��^�zUzy��6��{�#�0p�39��9��f[�Y0�F��;+/:1��ڬ�v��w�P��+~/�Z�w�3hw�>�+�|���"O���(�	�]�G9���������x�M̷ca����S�Q���.�a���&e�N�}�����ϵD�A�_�ox�*�����hZ�8�\�yO�:*1���;̋!⻤���O#.��);���eKd�E��d��UO��@vC��3B-8�̔����^�E�Z��^��v�D�x���M���q��t��#1p�)�L Xt�O��h���O��L�JB]7|*�N�M�\Ӌ�b*�V�&��zӌ.@�66)�<�&Ɯ�C��i���HS�}����	�~���f�xxq2H���S�E�KqR뙻�R]Jt���ݺ�Ih'_��Ӳ
}cJ�7ł�zi+�WU��U4MW�~"�S~�O.u��;잽���p�AEi���ƭ6������q��bH���އ�n����B-*��JP-�< f �G�a(U��loΨM�;�HL���vP�ј��V�����t�pO>fA�T�Fo��X�r�v��K�nB�^;^�Ӹg������ħV��	�T.����CV↨Zĥ�WWE��f���4twk�@�״T���{a�Ot�N��K$�s�.H�`����ж�sM�mF��
�Jm3!�r�8�r�^�v4�U��.��%�f9\�L��7��DN#WO�Zfc�T�VA�A�Ý��z8Bn�&n��6,��P�U��b	�ƣ5�E��\���S�̊�Ƽ�z��k���찏ty��֑#[�bK������Oۓ�J'�i}�q���2�Z��3*Gs��@�����a�����vb}��$3.����T�b-euW5��V��ҵ��G��+�񞺄�*!v���s
�>��粭�/j7J3�v��lt�2a��н�&�$'����ӯ@��j;��hņv;�\��ӫ����&�f^# =�\�!�'�w/ِ�����|���!�qh��b�|�����AM������j-��W,����=|3���U����tn�%��Nm�c�˨`L�\8ѻ�՗�'�%�5�1�;}�7���8��J�[�1)�Gs�Uth���w
����t��ݧz��0V�#b�ɓ���`�ǒu��1&�z�=��������R�4��R	�yVǉvn��E��#T�(��&t����vvRb]��, h|.&%M��{�H��wk;Ot�L���y��-],�8�;�O���T:��,�� ����Ai��I�uE�����#D��V�j$W�6��ڈ�͗�Cu�i\�0�J�~ߧ�
}y/��Zfj�;�0�Bi���D��ME��1:�V�w?�e�)S6��(2��6���^͜OX�o
�H�x��Ky����Idl����QQ�"�j����^�B^�  ɫ֌�{Q�a@�NC�M<d�Yq6b�cԭ͵=-���Aq�`�an��{]���\��㓯K�t�%��i5�MGw?D���S�١z��+,Z��M+JAq��]�(_�J`�g	H9=�O�馛^J��W��(�B�����l���j؊�涱s�O�p���a��}	I;B>���?A�<Ъ{C�Š�����V/+���b�t��W4	\���5х��<�>a�B= 9�h	��V�����D��27ֵ�`��E׹)�������'�C)�./#�f�p����>�x
�n��;��&����������>U`pv�<�l۾�\-� ���-+��h������5^XLb=�ϗ������+D�S���l�#p��d�Z=��=	�=��цD6�LZ�AlʴN����q���y3&I�O[�r���믪��
�(��i{���{���N�Es*����lĲ =����8��e�����
���$;�<:0�'}���׶]c�zf����wfN�uP�sbL�cB	�kX�2m��O���6
���u%Y���e�$P��.+�2 hM�ͮ���������Q)�P/�^�����w,��zb|�m�J��mz��K����`j �:T����D_+����F׳��d���ò."�r�y�E�I�n�Eso���-^�;��x���X�P�,ݩ[9w��߶��=Fz���u��h?:Զ�P�4]�q�b�8�wtE��x86D��!�E�6R��B���Uq�%CW0tm�{jq��`ޟ@�R�6�A�n)�A�܌�O��=sͼ���T:s*�"�_su6"��!�-�<�G���6��$P�2j*��gY�6w��{赻'��N�)g�Cʒz9���(Y�����=�Q���O�ga�-@�S����`a�wAe��ۼ���b�_e;k�`�<<��O�d<s��.�d���~�c��zo,��#�ݬw�Mo�<�n���z=y�*�nS[�e�:'R�oCf�}�}���>'G$/�f��G;0'w��\�n�!R�ڰ3)J sǂ��4gǵ�۰FIB��T��,� �7`�D"d�NV��N[q��]�g�}�HHRL��->{���rh�i������Q�%��ۋnQp�1��-�����S�H��n��n]d;8n��U��ʎEZ-���$����u��W�TS���;���祀�7�H��!�"u
vh�m�0��u�kOCi���)qN�7mD6wQ�ȳ��|��Qr{dr:p�|���C�ǘ�«u�6�%����,�@��z�u@�5�j{*Jz��m�u���g��گC�gF=-^cR��ڽ6�\2�d�L�6�`�,�˨	�B���&@��-j�'����Ttb�+�*/=�����c�(H����������{�+�~5�,�d�%IaN�9I#�<�
4��<���N���Zhr��W��ȐV�(Lv`ka�=.�sD��J���0oN��8[��.�R�����cJr�l��%�;�8a^�fp��4�|NB2C�(ݫ�}4�5�����L���ҵX�4f�z���B��yX+�a���>uOe��R"f�Q�5§B�	�1>��������,(]�ñ��f]�h�>�(�.����	���^%OB���V=P1w�B/�g�p{�1��zU��%��d�*���鷟��,g�+ͥ�`��0e�}��bUe;T�[�]bS�L�)F���v'�6�~��b!���2��*8�����o��y�v�p]�|4m��S�u�7��(�R)�^5�+u�&6���N����|x3�o7�3 ���{�f�0��x�+A�Ի���-yS�
���V��v�C�;��J#��m��zoZD3��K=r�� ��r�>�	��s�W�)�%'���{k��cH��C�_9��G9�J�g�E�6Gh��������7nZ����S��C��~B;�^WT��]���¢��~��imqC=��s޻36�1�Z������H��M˛袣��3�&lB�[Zѷ+���NGR֭����֠�	M�9HL��K�~��[�*�~�ec�g�-�;^y���;-Z��Dr��|ǂ���C$�5?!)���)�PX&0��vl�*�j�P�_��rZx�\ϝ�\uګ!���8֌r��L�c@#�ϻ�s����`��ʒ4�N�V4���7FfB[����J;�j�-2<���ʥx�Ƒ*���ϻ"���E��WfD��\ǳ�;e�a�%����-^w����N͍�2��Ln`Su�'N҇�p싈;I��Aغ]%_��PX�����_��'�kg�?����\�ݩ^_�¾z}}.�_1�y�A�����y��6Prk���7%�vP���d�U}��
h�������x�h?p	��B��N��T����e@6��\�I}.v9��Q)ফ��y�1ؤ��&'r���Ճ�`��<��Z�Wxo���g�T�@�K54�7����_ �go�m)n��3<�S|�eEI�����&F륐9����F��:<�/�-*DM�����'��-פ:��e���I���8��������שG1��m΋`�>�1���]���F����-xE�A�=S�1~d2a�q�^��V�Lo�<u>�)���r����SmΗ��[���f֍!�Ԇv�p̸d���:�^�'a��n�;mgJ���x���8��w]ݩP�P���C�������~�ƀ��s�z��_�.Y}��t�~=�o����fS�~l�#Pʋ%)E�ʇ�b�I����=^����xg� ���2O��z�T^=����i�p���e�z�6ׄ�ZM3M_��su!�q��y6�r�Pt�Ub8�O�	�18��sq֠q��^N�6h��F�UT�y�ۓ6�'QV�W�PeB��i�e���P�RQ]��W�w+�K/�3k;/��".=$R���ӱ^�w)�A�R��Q�aB�Lc��gn�[l>Q�u��X���n�r�(#K���yv�"�b�jЂq������}��׾��i��X�uq�q��_")Hl�^�4``]��Z�3V�>���G��@u �u�b^*L�J%���]��U����ظ ���g|�=��Ξٔ��S���Q2{D�Җ�%e�+\��u�]'R����:��}�ky������꿫�J� ���`�!+������X���Dv>5{gO"���	K&%ٲ0U��v��<.:�Z|h��㴲-a}EH��	Mmq�8��m~� Ǚ6c����}}	
��W�Ob�)��OMV�oI�]y�Rr���)P[E�1��1v��氀-� �z���]N�?-ss�_=(lR�b�ԟ�D7����Z~XH%�./#���0�����+:�R��o{���kC�.'f%��uķnr�k����r4�8�U�X��z��ȭ�:��i�r/;�;y%��!���i���<�2)��4ՀwJO�c�o7J|fg�7qץLGe�f�v��sT��\[�sQ��� x.�!-O�~���hv������+�1u�9>���ƅ���{[����+Z���GP�n����h~)�?��|֜�5��hgz��[�nI��}v����Ӷ�\u4h��y���Ƈ�����и�X??��9�@�����5O���[��P��=!�ő��`���z�h��E��9է�I��{�>�B:���b��<��J���Do������K7N3����S͓��7)m]��xޥdVz̜Ҿ��Wrtx�`����WG��E|i��Ǟ�{V�o�J�v'	��u��R��Õ.fX9�"��tG�NowS[��_�Uuu���}PQA,4L���|}RT;�ŭ���NluN6ۭ���T��>�h76k��~�db�mW�ڏ2ա
J|gl��k�B���g�!0���I�j==�v+�H8�0�&��X5��ҽu�V��WN�rz�3I{���!Ej��c��ߖ5���\���Vڜ���㰂{��½���ɶ����4��9�����[�fT\9��̂qu�%�C�;.�d��fAjyj܌Qg��f�Zے�_��hR�*�
j�q��.P��3Ĉ-�����N�]lk54�MJ�Kц�L��M�N`�9w���H����qvt�	�hUӍ��e�k��gV4A��/z3[,�F�L4�R�� /1W�"�ג�@؎�/A�-�H�9��L�M%���Ol�B�cO��O��~�˻COeIOW�3l���9�Z���8���	u�2��m��^�M++���v����zW�����x�sgi0���\���V��;=����^k'�m�J�^�{�b ��/���~+ʺ�r��pW����W/�|E�ڱ����)�^���C���oY�*����5����K/o�w�n�@vҽ�9R��[�1��b����o���Ѿ���CaZ-�}+�������y"�EX ���Ne;���
;ՖB��qݥG����  �O�BICCH�s߮���ǿ��޾~����}v~>��դO+���ܭ�
OB�01����Tu��1g�����mL��w��Ԇ�bV�W�'�u(r������ v��WFsFG��k�p�õ/�f^i�#7U�D�����xԳa�Û��@�O�Z��0�;\j[��/���s&D��R#�qE�YX�f�OdvU6[M�j-z)��!�%��V��%�s��Y�Aܢ�LIv����btE��E�@�y���'�E�`�>�,��
yI��$��y�F��k����oR!�;�QC�A!�(6Kup�FV�d묌��[�O������Je�̔�e��7c|/ ��ۀ�]f0چ�ݦ\e��y��M���&���N�L\:��L�`~!�a~�����eyH�Ω����qO�J�ݣ���­s[gP�+U"V��p��l2�*�ئxBcO�L�meƼ޹܄�7F$�j���g�l�s7	�G*	�#"S�]�.�zw^��V�ȥeWW�ƞ�>U�;�z̈́��N�P�D���#�O5 ���V^%:J�B*�؍��^ �^�/g��������ޯw��������w������/{3������������+Ӓ�!��Ӣ�Q�U�u�.2i��6�Hf�ƮӾ�E�F��>�!ǲ�D�9h]�3j� ���v%�vxV�hҠ�I�)\��(K�}*Cٴ�Y�n����in��2e����,��9�8�v.aq}�S7\N��6��@r}[�.��We�tԾ�{�җ��J�v���r-A*�;xe����z�r΅N��st�{*�.��d.<�.\�[%ls�]苺�\��W3GC_��eBpo(�o��˼w�+:���	��d!�-��m�m������0�kΩ ��e�/g��z�ht�M`�k���t�=��� �8A�d�F�XX�E�jQz3��nX�/+�r����Z�0p������T�̺T�"q�U��rv�7չZ��o#�+�����w}x�>���4�wޠG���[I�]�+�t�+��qᓋm���ʱW���ZGR.�RB����x߼��"�d�W�]��=���Se4��:��Q	�xs�Zi���T��c�/J�E�u=|2ռ�oc��&� �-��-˦�늍��ୡ�E�N���T�߆�D�܂�rd���V �[��z��(�O��^��c�N����x�h�~#�05�!3ۜq١o�x�m+��:����*g#P��_]�--���&)��I�-���n��%�J-!��s�C�w��x��[��,~AA���<t^�(B@����m}=wګ�K�o�����{}{��ARuN�<�<���\V�^��B˵��*nI]��s>BW��n��P��l�[��%	}Ө��^���[��F]P!=쥉Z<����z�zM�+7X��es׶��8�{&��{4I�A��e�: �Oˬ]�ў��T�+������%���Nw���Ґ2�}�7��y�g+�|��8�N�$�ͫ�B�(�8Fu[���м�墺~c��Y�n�̽�Ov��i@8V�D��3
�G;+�V�Sٽ�c��ȹ�������c�����<uP�,s����Z�.*��q��k[;�|�j���)����y���PR����Q�m�9kc��}+�vg`=�c¹j��l'c˸��dy�﬚�ȳ}�K7(�Qܛ�Ug�12<I�RM��y��=-^�_W�{s�Q�/:7f�!�A���GH�ce_3 ��H�ya.�U}e|��FH5�v�ck�qL��R�ND��C�,���Jo(��%�kWB9��ƽ�,�%���^��Ǽ�7����7��l�b� ��{!T)ks�;��0�#XA��}���X�Qj�u2^;��}6骋�2���:���Ee���	\�1�x�\������DPQ����>[�Kv��tӾ`�0�C���`9�c`�2��s�l���NpUo�ڻ����`�d��	K�mb�m�Ӥ"~%9W5�:�F�**�mk�0p�rt�/#DE/69*B��ZZ��U\6�A��T[D�x�3���֊]&��ɣF��vqnq��vΪ�#h��F���0rN;Z�)�h�����k��)�6�El�Q�[a�1h4Ө$*�h���j��hѭ�b��(�E-�N'EUʄ�s&��3͓0m�A;�f�AT$��RQDlj���IF1�"�
����@jm%;h6`��'E��5O6i��A���Zy��T���<�s5��,E�PӤՍ� $���rIc���DG�!
� ��3��7�W���>�q��%�/6(��ia�#��{w��:��|�ޢ��|$��\u}�j��������h"\"Ed�$��㜏�湵�ѹ�8xΏ�O���~�Gקpy������XٜIe�߲^%�k�zC�h�(>W�	�v4'���锝g�ĲN�7E2�K��(gy��O���\we���WsZt��&� �\�.Cwc@������EL"��Yn���g��"�}(�*�)�����1Լi uh�	¸&{&="��+���������خ槫;)rT��Z�O�a(�62��P������W�:mg��ܮ��1Q7�|��jb�0&ܯOM�M^�YB�Reȵ�f�*�Adi���PO����ώ�n_�����d��s\�^O���W����TZ�X��XW��Z�WzK���(�u,�C��?O�g�k�����U��Ӥ0e�`=E�C�9i0͸�/zm��ʤ��x�}��}:�L�5���y1��UE娎��,ڽq>���l|�.	�gЧVyX���n�'k�s�/����^���[�p��ăg`m�6:���H^�����&%�89a��J�/{Q��gH����h�Y��f�S�!�0vZ��z%�xA��# ��hoƓt�W�)��?g�ZD=�N|��$�KK��`תC�n�8���mh��ޤ����2�|�S����s��>�с��.��{�'.S��{N���S?���m�r\B�Z}�)�$ �Q8�0�#鈼��+�G��]�����r���|˓�S��B6v{�Ƨ2�z���t> tNo�%o
�4��#CZss�L�������|�Sy6�r�PgT��~hl�c�gQ׻x�WWʶ`�ሳ�쾪����DSf���o�ʭM�M^~�
�͛j�*�gt�X��A;g����,/�d��hu�>��IS8�(ǟwq��5.�.��8��lAq��,�ox�yN�1j�F���%=$`�as+�_�EzqW5?B	�Q,��8�Jw2�����
;�7)]E���������Sۼ��-D�f�	�����Q��9�/0��#�q�~�ADJs`.�L��I��G\�6=C�@0�m0��m�pd�o+�p]��,�ʎ��;���ƕ&|b����oH�AmĽ��>G�e��@A�Ck���t�;�������`Vܦe7�����0�Bn��Qi�c)��#�#4���+�{K��F�7�7��,`Paq� C��Hىe�~�ɦ��5�vvQy�R5�9O���h�Pr����34�og���ݡ흇�`P>���;�|�s��s�rO�[=A U����#&�k�=��)^�_��݄�'m��G$���{l���CZ��:�x��O��_��y�|B��]r9����p�0�u6�@�kd������HZzK�B��j�;�"��{1�vr�Ɓ�s`�{���nfJ��
��˻�{cgF���o[���S�
�h�V����������������7���e�(t[�2�t0gA��y��!�]�uCs��84-Q)�ei��)m���z����Nn�^J<[���U�%���GP�{Q�.*<!�t�N�k{�gtS,�l���E���HA='\r	��
��;h��e��c���w��}�;F��X��H3��헎T�˭�uHLM�P~s�dA1<�@�.Ťq������O�ȗ~M��[e�%�I���`�;h��B&sc�q����� ̳L�]�yڼ�� �ȿ�E�5'egcvj�6]��9�	�T�\�w�fh!��[�U`O��v��ء ��Z�W(4P�ZmܵP���e�:U��u�ٶ5�,�)��)��4?ߔ{��VE�2�x�6{� �X�coc:3�^���F���c��Kmz��/�N����}����("�Iq�&'��F�i-��N�Ǭ�X�!	�p��s5�lb�����bUˮ-��\�:��g��[��3ZɈ[�c$sl��ҡ�Iv�m�ˎmd�]'��%:��Je'��l$ȶ�э��W�0[���6[�t�^��$ٹ������[K�n�J�,NX!�NL�*�sL:/w�#��	��5r�P-�秛�j�<��
�{Ծ���ǫ�|~Y�NV'χ\9N>������3�:k�+݇ ��-[k�<����<�1�:M�퀔�v�}U��-_�RM�=��D>�5��Cg� 醑�F�,�x	��9�Rt��!�K��w��6�殲1B���JF4Ð_���n!��P�;*Jz�3l����'��8�D��KCӘ�G�VD�$��(+0Å�0�7s�B~�Ol�©�J�g'0Q���5V�J���y�x�LQق5�H�܅�~Aaߋ=`D{˥O&f�Q/|�GA5�څ�
{����0�j���k)W0-r��ۇ�|C�t�}ni�	����H�Rj��չ��c�^�
`;��QNW���Y~��S��ПH��4�ro�5�Y�C�#�ԫ��w���i�p�_W�����,9�� ��5��ݣ7�j[��@��3�T3Q�z��D����x�n�!اDwK7Iܢ1%ی;}&e�B`$^���(����cSASb�[?<�yw�!H��ݡ=�Ȩ�D��v�^;���M��b{�)�>�#v�C 8��CP�lh���Z��(E�d��]S�Vouᯀ��������� ��C�����/���Ӟ���aշ����7�O���X���nI؊�r�3ז��v��=��(�[�s��8��0��)ēY�����Zеd�W�炵���w�7	{���e��N^c�7�+����o:��)X߰�1�V>�9�Ή�-x3�|�`��s��������W#^i��[����tS>,(���]��4:Սaf��ŗ����H��r�R�եHZ��eB�Ф��p��l:�)�{bY�M�-�����{����^GLp��/C�.�vq�F�73r���,U�B�ܮ�g�u�`V���Vqx��̓��g\?
6ŗ���LD���CK�*��%2��)�PX&>�U^x�n���nY7nW^��Uk�Z�&e+I�E9{�[C���F�ߍ6O�<�����=��
��O���T�a�j��ru�~���s���		��G�L��,?ճ�z=���,_2�^W�_�"�S-g�;�Pʌu?�$�*0pN���`3���+"X��1=w}��]�w�É�3��Z�O�iAcAt�~dC���}"6��CM�|.���fk�i�oZ�g�t6XVԆ��sbzq�j�r��*��Q��eH�~Y�KӇ�; 8�]��35Y*x���c� :Nk�ji��d�2J1�v��\���{���u,�q�l�1�gU�mB��s��Z.48|���R���J(Ձ�MW�8	L]�ݽ��J�c�R�;"j����-m�I{~�r�/����VN���Ը�#�RSۗ0�˄�*����"sk]��Jf��g0��1���0gbӅt�S��G��}����������f����$�7{�6�f�z�3l�K�/Xj:��\��;���T���\��,ƌXgd\3p.4B/0��Nç�ݐͲ/��!�r
:���F��}���y�㎂Mv��zN��-C�C��tK�y,#���_=���ݤLcj���6�;��`����`����8#@�i�K���EC�{"Y�--!���3�����"L�W�k�]Q��鑍�73M_Ia��P�%��]�3��	A���i/�o��e	;��}F����j�k���ʷ&l�nY�������
9A�fͧ{�����I�Ηh��o2�p�e�W��w�8?����Eǧ�Uc�N�zGq�L���ɭ��5�ı�%������m�,`���Ve'�>��?1�`p��6=��� �1W5?B	��G!�ie��ک�}�2�1�@�4��Mw����趄�o��$*$�6W�7�A
���
bTT��eAEY8���%:N��:!t�e@�������Cϑp迬���%,��q��=媦K�����{"a����E�7F���I�>�t���K7�C"�5p]"g</�9�f(AÃ����LrsѪ�e7�=��,4�Z9L�
d+�͡�h�t�n˷��.� �{�׫��>@Y�aͱ-u� Dr���zɾ���!��=�>˒���V~��d�I���4�㘤�g<�T�}E�1����~��au%�E�u�һ��L��P>i�)���/d�:�ۦ�u�-?,��7������Z5˚�/+:��,7��\:�vbX�؞ɦ��8�r<�Z��a��v����J�vG'ǻ�z/D;��u����gal!��<���:�¹Չ2)�z	�k�wJO��|�o�2���>�'�ob�|��~�1�!9_s���5�W��  �^|!�]��n}��B�.��f/�35��M����rv=:�W1m����!�A���Пܜ���i�#{��=��I&�maw=N��OO�˺�*�I86��;���uƀ��Ƈ����re04Gk��Ӱ��W��.��.*5����X��A�4"��.�aض��q'DYz�o:!���
�6ҍ�".�t!�XQ����uN6۝��fY��y�-(�P�6�5F]���O�/H�U���OY�T]'߇AI1���~��DX񬽊��ϫ�v��$U�A�w�{��By���eJ~�.�9cGg�në���ծdյ��E��W��>������U�:��Z���{�)�Nh�+��+Fq������*���<��*X���N��A��x�ףN��-�F�W��wưp@�(;s㖾�nͥ����K��j��ꩦvuOJY����ׅ6Y�cW��I1c�d���F�0����P���L��ee��Ƀ���A{b\�z.!�	uc=�|jQp����'Iq�&$�-�;�NG]u�ѳ}k�:�{�p����Ek�s2d_(����Хr�����'�T\:��g�[�r�{LD��՗ѽv������󲾖b; �6�Bd��ħI�UI8��t�	�hM�S��L��^mtu�ٶ�\kH�9A��3[,�s�=�>�v�p�V74�Z{H����pY�E�k�/]w����/�T���O�}�'�!��~�0��YWa�i�eIOW�m�uZ2K���r[ov�H�'Gf��r��z�B�=�5�ޑ>𓶘\��r����=SX��+A�y剨�R���D�����RD�,��,;�m�耏���TW:�s�!@��Vv���j�CJ�Z���c7J���L]�<@�@����-<k��;�ɹK&ҳS�x�Ol���	��UL�c���Z�⠗��Q�$�	����:�-<��t�Nj�~;K,n�zV��]�ܩ��ewӽۭ�K�sn�s�-R՝T�]�2��M��¹]L���յf���Rσ��Tn�E�<����^�%�1^������ݶ���2EZ�2m��O�R`��J4�o�J(�7c�둾0�N�1�0M��}��Q��q'��ъ�����!�n��a�@�T��5�~a�v���^��sr�g����X�&��tk��X�
�R�]����R�@۔XP&$�W�˱׺��ڥZ�h\=���?�`vv��,�STI���"���d��b�ާa�e�iG�Ofs�6xa�D���hi$˴��-�{�mᎸf�1���@��I��Qx��D�o�r;^�omEB/U2�ҐylN�rW!
�#^in���`�x �������n&�qqAف�9��5����TcW\�K[V�!k�A�xZ��7^����.B���Ea��*
�s��]����ƴÈ.�峍�������Bu��HL�֍
O~��B�Ӻ��T9��,�3���oco/_���I�����b��8Hu�x��Q͡�	L���S��RX&1mZA��{w�[����BGNc�m�'����[@N�|����D��ק�e'YT���wZ"�Z"r�#��|�`1��E7QF�
�|��s	���>yq%��c�`��G{�tCM�i��=�Ι�0�+�Ȏ�3��J��8{��&zm�MIH37okĆ��=�ӱ���i�H�v��2���R���ic�P�7��~2;\��gp��q���"D��#�8�وN_.�7!�>��F#.s�T��Gp��H+ׂAN����Ԕ�%-'c�^������Rt�)�]!�ʖ���1�噃k�p���3cH�u@]<���ǥ-�K�P�~�(➗�j-?5����Zy0����<�#�찏v�cH�X�0��n7�Vc�8��(Be]SE��L��0��vJ�/i����C��8���"��Ư6�	�3��Z뷝�h�DS�(���[SM���E���J��x���`�%��)?3&K{U�W�������ʯ��!dÐ^�����!�q�^��+2�1����F�K���<H{�w�\����cq����O�g!F��æ�k��>��wO�7d3m���5��;n���(�zu薁�@��W�D[��s�]�,#C�q"%M��<#�����?��H}?��)�~�v��`�~�U�,xA��#<�Z�-.���D��ZX�*�{i��(�v^�t�C�:�}d_����P֑���l�yrXrU!����ȼ�O����<9�/�fpu���{�4΁�-�:l���f=�7&m�)S6�A���	���<5��?˟O��������}��O���z�~�����ϰ�ŀ���u���B�f
.�@�`͓�P�!�`{��$�e��&Z���	�����������R���mn�J2�~��a���a�i����x��Ӧ���ҼХ�˳R,J{�V�׽w
�L�-���.��nø�uz�l��4Q��^h3yW&/�(}u�y!-�דuڞ7����q��X��K1c�;�Q�y�D%�sÍ
[ �Ĭ�m!�~o]]5�.ȉ�J�^6�]��#�:��WFOyk�T�1tOqtã�]�88��o����&��ւ���@Pt�-Yp�z�`~�;����cI�����]9�e �K݋��ݬ�ؚ�:T�ZN�>4\��+�{��txsqA������"ņ�|�ɝO8��ȗ9����"������2A��;���5�G���yw��kA;Û�S�i�_(ۧ���p���{Q�c�����f��1���r���Y�/c7Vx�ۂR�g�*�3$�KˊҶ��%抝۹1�t�����L:_[ �(C�����c��.3)rJ�my�C)!���s�͘�Y��w4e�V�\z���=�n�<3rx�g��J\:����6���z��r\������Y�f��pA�Ў�IǦf��U���"�������\�UϯQ���t�F��}��:#�.O]�������nL|h���tx�ynk����![-�'F�*C�Me��p=z�@�';o��ؗc�l��ۈ�+�d�I����5����״�N�8�>��7��`�C1��~%;�楶s���.������Uw�5S��[oD�y9�Vtp�H�ݲ��}�i3�^�wG��{�'l���l4Oe��DՄA�W�h�^%�'Q:8n����z�D�y��V��i��,����:4|��c|��vn���9fD��;%k�xyWƠt�.��	LŅI;�����q;�X��q����U \.�Xm�W���ֽ����i}z����=,����{���d�/rI/9E7����>�<&	]�F-p�t��a����K��g�`t#�n�C���9�f�ݧJ3��\�C��uA�.yHF��=W?���|�����=����ӌ�OF��`�M��=lc{}����J"����%ҹ�t)�سz�D�r��MKHs�bOYR`�З7Y�p��r�Kyԍ���xV�]qe�9v\��r������(�Y��ٻ�Xf�.����N�v�m%�N����0�hE-@���x��	�&^��H������n��>��u���w����9���64U�����ɔ&(��&���\���]���,��	�t���Wuܦ[�\���"��k���k݋��G=E�<�=�b@W\.�N�v��,TPB�ct.0Y��[���7'2�G8����1���ʆ�J��ML����.t�9�ks�7�j�x�5͢�lU��*�
�mN�y!Hh�����4MU��%%j�ATQ��SUT\ܹ|sO
�3�b(�<���E<ښ�"+��)�Z�9h�-�TUS\�b�xx�(����ʶ��"�\ы���i�[N����X��5����xǆ��͙��4k\�6�sm�s�'��6΍"��5����Q:�q�T�r�\��9�n[E\�%�6"��x���.bֱ�Us��gsh�nUsk1��[���c�[[��W���"�k��pۖ�Em��71[�͵4S�<����h�8�Ʀ
��M0DISlb�4EIm�<�sns�\�s���k-��6�ns�1��9����7���lF��k&�b���2P�Q��M[X���q[`&*�����QC���DQM�V� ����MA3El�X����������zx�o<6�D�mౕ�RwN��5��N��8����b�0�M�V���
ww:r/��ҥ�)U��9�ys�~km�ޭ�t�w��ڽa�w��u��`�kϳ��M����o�	��p�P��Ӽ�<�`�Fc��o��
N��	~]���\ܵ�����(p����ai�8W-��Q,��4��U-\";�e5?R��H_x���NP�d3U�6E�l���s�Cu�8-R���o�I�}1�l.�L�i5��\���FFC��G�@0�m]L�q�M�!ä�j�����'Ь*�%�1Ѓ��m`s���Il���х�ϴ4�D
�C���a�~�{.����"m0�l��5'�uL5ϝ6��Qi�g�)���9�5�k��sK_U��J�/U�|��-���=1�Blp�����.ѝ��ߵ��Z��a�,QkP=u���^n״4��ơ�'���6~蔈х�u���%�9�B���ˇ�+Ʒf�z������������y�S�52͛^�wc��AC�q��~�u?*�uA嬚����KZOve��(��PO�^���]~����_A����+���_��y��4;�9�*��"߳bNV��NF�$K�$�[�w�X
���T �zq,���{g���v*p=av���P=�V�QL���Yv��oAa���+m,�;��1��b��X��srjK2Q�Xt�rA�|�� �{�$��jL�����5�jd6��i�����.]�6r�vi'ә�8��5b����+	�z��]�["��}=hX�˅Ag�X�ԍbl��w��W�ӵ�T�&��;���_��d3��M��'R�*ˁ	`!
^1���T�m��7����4�t�v��� �8���@ɵ���7 ��'eO����)i�l����I�=!���������u��Ƒ��St�wh�m5��|�3��x���J�����γ�͛e^�i�S�$ŏ1�`�$s"ė�W`wA`͙�eu�e#|�U��Za��]��	d�M���Ƭ��sn� �]�������-�/f��#����W;/ �q��2=y�e�~��Z�B�),%�\[p�뜗��ݡ��!U�9�֙{
�F�7TƗi��b'ݒ����&I�9�N�2)*��]��gy�,��qMLwswC{CE%%�F�4���@�!�5l�G}Θn�R�qx	���"�D�e0g�wk>�.��B�t�|���<A~ǡ.B{�L3���ʎ�8�ݕ=�T��=���)_�d�,1�]��s��2Y3}�U2�s��E�s��g����R��?s/�z�E��8��y�GjW&�gW�ے�@]rJ�n�H�j[���me���eˇ0S���KN����{�+�ήs]��H�8���ok��������,3�m�ߎ������c�Y[�՚� ��b������w�5ʒ�HAY��@ׁ�T"��T�P�{M֗C]�gfM��Q|5Z��JO-j�'�	Ϗ�?mA�$L�X�8v�!3�"n/w�����Kg�:���b6�	�j���qvJ���c7J����}j�+]��+�q�U�Tg��P�9�o������d&U�!6��4-2��;���{�PK�X����sY{�kk5����~y-��m+u���3=�	�@t��s��c|;h�棩P)�'��Fƥ��9x�j��r���.��+S�Ղ�vD��ȅ�����v;�����E�bK�SE2�K{����F>�ݰQ�Ls�G�rs�q��Š J�^@���¶nq���v�9|5P�W���Pz���H\�Pi�e�N�U��6�ƀ�π���e��d��+-#�i�XU�Q���y\���2����i��<�z�/I\�(r5�q����	��V����N�~���O6��rVJ����������������Хa*:��zq���C��I\��B���u����uc�s�l����re7���F@P⾡�)�o6���dz��z%�ۢ�d���;��Ľ_+ͬ��l:M�L�誐�6�a�Ɔ�5p�)�%�+d��ʖ32޴�i����u���	5��(��*:�i��\0=rJ�v�_��:���y�lJ��&H��Ҷq���n`6�3tI�F)	�
��ش�(���!��l�I%����^ӫLZ�Pf��xyY�/z�HM�x��;�P~BS+/�)��L^X�9�:s���d��p�g�B�GNb�[�9Y�_D��&�ʘ'�_G����^U5ƪ���yZՠ�Է���C�k�4�S�_8��s	���>y3d�&�����i����n����\�QAN�E'L,#R���]=�A�����"�*0pN00Er`���ZDlOY!��۰+nS2�����v�8�8���='��JK���.5�BR��^f�}����v��ja����0�&5��[�0��v*��Q��lR���@�<�0����8)�|���Pl�.M@qa�ް�ǘ2��SM���E���	V��OJ׿�����%3[V��YT.e�NW���� �a?�H�_������/zm��ʤ�zI�����V>G_;N��N�q���,ƼXgb\3P�`<�wh���;��a�[	F�'	܍�Y	FEj��X��M�r�p�������7�wݱu�k��*�WLQ�52;=Ǹ��oV�3��ig����;@� l��)Ҷ�܇j�l�PQ�����d���t�,�5�Pcv�����Q{8���@�8��lu��Iz��;Iy����C��x�����&�v�=�d��&�59�<wթ��׽��Azn��r����c�����ڔk��g;���oFUV��z��`�c"6L=�O@�^=��ޏP֯fѦi��,:�WAP]�4?�&��Rkyn��l��u{�h������J�c���Oz����F�nL�jJY�� ��l]Ļ=�<yڤ�,��v�-���^ǫx5�Q����,9.���S6�.�^�"\c.�ŮFi�S\���8N"��=�{��+�FRk�=�&?�l"�`��<���G:oM���W�9��*%�{�Fi��4��#��s�:y�iD�@�'���":��qy������{�=�XtH�;�y��$�N]�?&��ʊ4���z��y0�����s��&˝��]�ķJ['��ܓ�1��E��#�L8�)?y�Rr��E*h��z0���Ύ��͊�U�hb-������@r �И��"�y�9���tڪr��(�
.��|��R�N`¸d'[��b�{۞�A��ܨ�-D������MײuI�u;|^ߓFg]n��W�.(��EZ(z��`��k��BMe��T��I^�4!7waqעhkO=��$�N'���Zs�9�RwZ=�̵�t�{FJ�Aށ��w:�v�1��q�$�Y�;���f�H�w��vC�2!x�q|�Od���8k����6�ک�f�Q%�����Ix71��������z%#Qjd.�k����X�u�dS�q"vV�*���n.�jv�)I��b2m��)�l��i�Y}ฆ�!��|:�y~op�/�TRԤ힘5/X�����j��M��+O�[���u�W�Ө4z���.g7��	�s��4KL���6�Z62Ys�;��ƥ���i'���i�qh���3t���1�P/a��G���O��K)�p�gh�����6�k�l���(h�n`�r��㿋��[{���sk�I�P�b���s����/���)��N6ۜ����,�4Wt�v*�$�kÂ��~�V�q�v�[�_�I���RL`�}�<!�����b�端v��貺�g]8Ԧ�)�CO-��75y+��Fu�6)��gO>�{C/�H�)"8`v���% �e�����y�C��/4�{L �Z��A��ʒ��r�om�ʋ�5p� �Y�'&/��.R�B�t��"�WWJ��W������b(	(�hA���L�i����������,�wWj����pa��P���_�8���>"�TP8k��Ly����_t�J�Ae����smp ��5�s��Z�s^��SvD?��1�W�}�pao�f4+.7�1)�Q�`Tdz��B��<�[妅(RXKjܜjQp�%��<�9ǩ�Ӹ�+���3�p�ޏ\)f����=;,�'�SsS�&I���i:Ĳ��2��RʹqM	�b��_V�g��T���E��8���@ĳ�AňrO�e��H�醑�J�,�&+_�I��kKD�G{#:���B1�͐P��/N�o'ېaa�^t!�˭/�g�
u���Z��9��k���X׵���[�H%6Ⱥ,㛀{�F���r'����z����{�Oԋ�}�Z�]uTg]_&܎n�Ɠ
9�[�j�'�),i�a>��D��<dKQ��'�����E���b�N�����B͹��.�	TXU��c6)V�-r��9���o3j�xq���$�<z�#�k:�ֹv G��ƺ�G��=F��j�u*�u��Z�◥'��	��Нk֩�M��gB��~�r��Pk[/�?�_~�c<�Cj��h��:��S�ֿv���$��sS�`�4�BzZ���0�x��u8XP�y��:a^x��79.�:��9�~�{h�߈����m��ʂ����2��ѫ�.�I�?c�r��\�S,���ޤ�ۅnT/����jgW+wӀ�b��z\���
=�'��-� zh�T=�O�oN�OU�����ԟ.@�xQ��sA�$G;�/Z�=Pp��k)���1-�N�n�����'+�q�y���ߒ�k���m�����������hy���_l����mqw��]�m�G��(%��$=� ��>�1Jݗ���؛xc[��e�0��wm�e���b�j�:�O~�R*��u�^>�5���/@%r��ךn2�5t�ê�E3��%�ۚ�e4�m��K�3kǜ C�q"3&��_N�ʖ��j2�A���$������c�9Q�uOi�{��b+T��
)�M����`\��<�1���mn�Jl�R*�
O���+F�en��Txm�ܼ�
͝׬z���S�;@@Ŵ��K䉀��_W�i�y�?!)���_�}X�k��F��:�Ȭo,/�)�j��w���z��xOm��!Ŵ'H>T�����B�6��c�WO\'�_/.3) �ĲN����gΦ����]�5Z���=䈆`�Fo١���Wep6�'���KOCj��bi�/h�ϻ"���E�x�T�P�_��hw��G$O3��3z�8���q��)��E�-�遬o��:ҙ�Q㊺^����֔4�L?5'�>a�r]��ܯ?#���OYmէ�eU������"��q�z�r)sw�M�7�*P6���lC�xS[�����Zj�#�TbZ5],�޸�kR�4$�Ѥ�{;}z�W{��'�B�޵h�T���*9��RQ���k���b�^���KT��/#Y�$J��>�o����{jh��3�a7"��F^��9�J����1�<eة����r���Ɩ��@p���c�:�Cji�X���Ҝa���v��Z�C��>%�����t)F�����vB�`�C�0�������dd�>�E2%�a���(�3۩ﵦ�V1^/
�R�F>�3�GrY����A��;�@Q���
ug�U:�|��/+�e^c��z�����g�s�-��1G�(>�gƺ�GӜI��/v���U���C�=��N�ǰ:�5��ŽA���0v�rC︴$q4� �o���T?l�'D�p�؝��/�smy�KMp�L�9hd4dkL=�O]@E���7�kNnf���Ò�o�Iw&�6*��+��n˿Z�_�LL�P�>������΄l�^�����3mȩf�eHC�uO��p�f0-X��2���D����7ύ4�s�S�`qm�Eǧ��7�\�W��y]E�c��{-h�A�Z1)�Q�a^=��U��B�$���2`p���x+���yD5K'ޑSm^�����h�]Kw9�ث�����![�}�v|tٲh�=	�U{	�����쵨��}ymh��/`�x�]�f�ئ�3�^_���Ov��*���p����&�s�����U�8�/NRsi�/h����F9�L���-O,�����g��ڜ�	�r�d��F&�D�I��;��t���E�(.*��Zm(?-�f��L&o��$vI���'�)��˼Q���=���=���{�[��`�41�Rg��אT3cL,�Ba7��{�L8�;��N��9Z�$��H�����S
�2cf�^��F�i�סA��f��B<�?6�f�y����`�gZ�qms����Jv}
.��e6�r��k�׀OD�f����-��ZQ��7c��+�vJ=g~�6��b�^�������]�p�p~[�(% �Cג��MbC��b,(�c`t�B�H����B�ԌZ�Y�mk������2��o�kP�c6R~k��y�J} �����'f�
�q�w���/ߑ��f���Sam}�C�?Wj�j�Q)�W���U��O����}�A��ᬃz3q��\ų��[����Ш�G��F;�ŜhGVI��B�R��^&+��~�q)���eT�鐩�F��C�B^��"��	�D��66��5��7�?<��uSI1E���.Ÿ �^�w���}=~�o����}��O������|�~ͼ��;����4���c��T1�뀡�EI��h���kE�uk���ҳ�%�@F-��'W玍�4L=�q��L-���}���Â��ҧ�&K���Al�	��,��-��iR�l�_s���᰷��r«NSatu5�,ɑsX��iq�D7��ӄ�0]���gf����Rj_9�=��|G�=�����Z�-���Ɉ�� ��1'���p�.z'�Hz�� Iu�����Z�e~��w��UJ�+���(
P��򺂥�:�h,mi�Y)�ꊙ|{)�=���3w�Z�3.��&)�PA:�b��haߪ��w�/)ȋ����S�OCWwS��+����&A�2J����g�&&\�S���ѳ��]�����?���#0���"�ZC{��>JΗ�m�h�T7n�du��!
���`��hcή9�FB��:F���Cbї��;��f�%M�/8�M[Pi�|�5.5|��X�n&GT��� Sޜ�5л�Oy��qnf���$̴��Y�|wG T=���nԧOy��щ��|9KY��v�\�g�Q��]2����%vײ�w�M/c{ɂV�P�怶y]��6b�'J��;X`�c;;�t���<��{���M�@�*,���H�r��a&f:ԍӋ^�`�N���3��"���޾�R��_N��kG�e�1�l�uJ���(�b�n�1y���m3ښXL��+V��p��[��N��b��JD��� an����i���:��ּԦU�%�8@�����W7v�n�
��N�E%B�&��en+��Cgae���JT
�eZ�k��GBmSi�U��x0n�w����ף�3�r��ێ����VmY<�A��$n?�ӧ��d�Y/���N�W]@�W&{����r8���7KͫNk͜w	���;S0�	f<�'������6_{z��`kէI�.[��]0Q�N�����5\�XٺOvQ��!��$����Mt-���e܏19m���j�"�c(���:��&x}8��-K���x����'�]X��2�#����c��l��uyʜ��QZ.��qc���ԇ/�;�F��q��%�큱bW��R�W�سm�u�C�[�#�Aҥ]DjW5r9��o7�i�{iq��\�X�֬F	l����ď �@l.�i^��(���ո����̳��t��Vд@턵^�����M�wN����4��S�M��N�3˻�]�/L~�|+v�o
"�R7�ݮ���r*����d*`�κ��kS
�������4w��ڲﻪu)�C�=��>ۙ�Ԓ%�Tx��)S���C�i�����z�X����yB�j����У]���<ov��t-`y�c��i7�g^��pU��j\jgI!�i��wF��`�"*�"�0fڂ������j)�cALQS�3�8����	)�e�h��"N(��+X�t`��s���S��TDD1���Dlf�����*�uET�ED��E.٪

��b�����6���x���5F�R[b����4�QTS4�.)������vĒkKET�SUSTU%UE:�"61%UETն"�j�b
��� �*��l�SLQ1sDTVQ35��[mD�MDPh�DPPDN�+lPEQMQST�m`���*��*�"�("j�Fb$�b&�ӋFb�H��DTLS1Q�b�������(���IERSET[`����K`�N�f ""4�lo9US5kK5�LR@TATQ[i�"�
(�f"(�9f��#m��%�ɇ5D�ULQTZ�ECT�ETTI?`�=��-{���܄4�4A%��'Ǻg��D;kF��tH!�D�����т��{2��+k���z%�WNsn���>���N������d��}e�*|�-�KA��"��'�&�0�	�'�7����y|p?i쭫����.����mௗ�R���l/�-�&u}S���=�>��4����5����G;6<�PE�G���mD׍CT�5��9��l�w������N2/�W>��7x�۪�ŝ��Ej�CYr� ��@�:ϛ�r��y���0R7C�{���a�k32zJl��ʋ��������5�A	���	ͨ�.�g�=���^��KGj�T�8Te^;�����`Є�B_\t<k�Y5�\���A�89E'V��Ҩ����8˹�,�2l���Yq�ծEj�{/���!7���]	�����Y�O�%75?Bd���u�Hдq�O��Y@�uNhЮ{��]�Pf�H�m
�q�!>5�,�@�rH�l;�0�ҥ2婠K���py�XX�i�|�w�8���i���w�xa;�!#}B~��G<����d�%�F���]�N�M����ƥ+n
�/���P8�{�F׶k�|��G�+0p��C��ϒI�8E�5�ҽ�Ǯ����	�B�l����-V�Ry���4��-BD�܅�PXv>C���y�H3U�S<~�^6�n)��*��[|E���n�7J�v�rF��6����NP��o��&��L6����\6�r�
 �#�XK�{'@�4!f���
!�Ƭކ�@�"k��ۛZ�]�{�z�;a���������Y�˴�M�����]~��I�%�/�~ƷqlK�ʊ.�Iȡf�8��E�Z��3t�Z��hw�A-Rm�̟3]���X׼,jhyj�0u>r�#���uH�����t�q���{*	{k���f(t�G?���}>�򎺼�PJ?�	=���A�g�f<� >�5�,�h�&�u*��ֺ�q�.�(��utC�&n�j���QU,Z����Ɂ���x�	��>16�s�쓫�n����b�k��]]4�Wj�^1�.�^�L˴�ϫ�������<Ěy"�,#М���b��˰�=5h=��7j�4�#2,�Wt�C�	@A�v�pE��xc����X.	Z����z�����>�c{�'�zǦ�؏{��Zt��|��N�{�.N�d�B�w9�y�!S>�$�����ħʨƮ�9R���*B׿a�U��Jң�&���j�Y��#��l�n9_S�S�6)���Ʊ�c�C��i[8�X��nj���/���u���|�٨!Z��P�w�<�Q�c�;��*�iYF�Y_��IeL����CH�S̼��nCۆ����ef`Wy����m�Q`uk��2�����P��e@��r�lV���W_�,����^�d�ِ���V�Ʒ(L+y�V�H���:���S�{?��Z�����d-�ѡ���\�u���S�U]r�n��뚪k�zn��ٟ��4���"{��w�ħ�I`��B�F�c�m�kE��(�BYl,Ɂ��'5��tK�]�w9��u�@�z�3):�^%�u��)�$i0����!>k�G�f���V���Y����Xg<1k����B�e�J��Y�ʖ���^��-��[�].�ѥH��̞~�{�.��"u	���_l�(qTqWKը��֔4�L?7b�a��v�lOG̲I>��*�Y������������L��u�r���˛Q��B9!�����E��\[��u���9��ǻ !എ��؂z�f$�ު��s�B�k� ��6jj5c��n���������}u	����������&����GS22`����||x�^��v��w�kihz��:�lq�N�x��c��A��d�f�\<����2�緂���ǽ*7�y�Y��Bkٰ���-��}>U�,v��}�
��}�>��KxU��l�2���A΅���DJ�Ocj3\�h9�������- ���i�/����>W�ߺ&���=��Io=�M��[I��	�^���SW[Э]��������T�"B�3N˸Zx9��-Tz�!�\�5���_heN�5�v1�}����~��@ULS:�]7cvh�U��N0�]n���n��N�o��i�ڷ�lZjfJ̲�p&�9�{z*:�U�+S>���C���!��x���	����=��{;�1�,�4�}%�P�WA�F�Ww�NGeY�p�
ɲ�ͼ4��=�MHw���F�ӫ�T�K��6��K6&�f]�e(���&���i�����kW�����6�i�`"��`p����:ª�	]p��vdaM��;*��z��%6%2b�4�ģ a�y��>w�yXũ?��f}D8E�K_�t=�⹚Ǭ�B�e�7!D:[��f#sW����M2��$f�X�i5�Gb�\����1"�Њ����f��;��8wc�t
Q<�ƥzK�|$!#�O=y�%:O�"S��S*Mmb:��kz}�8�߮V��N��-��A6�#zY������*ʖ`��L8��Fi'�1Iͮi�Hθ�ӹ��n:k���.�Zýn���O����¸��Bm�1��og���T�H9	�]�R��0�m._C�إ�z��]���L�"�����#4�s�VG����kÐ֙��>���u�d�R��xCΚ��८�KR��)<���i�&�r�ćyBF���6H.��{��j/��H�xM_B7�Z��<
v�;w��/-�s�|}=��b�ݔX�v���9�Z��h���{Z�,he�Ǘ���H�i��rn����xr�/�od�E�g��hdd��^�؈� u>�7���\>^�L����K���ځ1����x�0uw{0ъ���h�UO�Q{�NH��M[]�Jo&�8��R�A��l��n���a�p�6��m��������d����-�P펓��&��4-XQ)�?���-{���駎@���;G����`��z{}z8U��8g�M�"�OS�����?���N
n�a���v���4���wL�7Ќ��r���uK�X]�	�x&Q��(![��HL��P~yp�^K�E�qYQ��1��"+4+�ti���|� ���~T9Y_��I��X�o����~g�zz���!���kX*~N]���{D0*��L>r��`�?J3�ڮSj=_l��y�>��·g���e��y;Ä���y<�׹{��H��C�� 1n+��FC^D�΁l�����K1w�_j\\��ݕ0�pZ]ڵ�7#��9mCL$�kt�P%�]6Ϧ;M����~�S�٤1�(f[
u��=F�%	x"Z!G#�Y��|�/�h�2���+��O�Oq֌�(/T�S���jU�K�<�3��z 0e��`�4ý���M�A�$�ħ[���2��t)-]#߫���mK�Y}�	�/���@����/���/#:���I���澢� a����6:ѣB�4b���8�l�h��� 6��Fk�q����#�R ��p�u�1�$�{�ז��[��{yӒ��sjl��3�n���V��Ҹ7�K���������
w�'�9��7�
w�]�5�n=��o`���] �D9��r���:��d�o]'�0�`��#�7 �b���)=�Ч^������q�́��"'�pG=r��\��v�a�܄+��+Ȫv�r�5c�_�����{�F׺k�$�*hA��Ρ#_).y;N=���SF��C@�*�2�/U
V7�ŦbrW<�z��OiAc^\jHO�ѹ�V�U�*v�7*cuN�oF�ML` ����&\���ܜ�k�qv	TXU��c6)V��^�Xsx��ϋ�(�4v�6R�4�z�^b��CjF���hZ�R��ҵ�%���ĵ�SӑS���,�������U�����(xls��8|O7�,�n�j�Ԩ/ͤ$�MS��1�Lr�󖺜�@���=Lx����T<��=+��H����M�X��d�����^	͜�[w1°�&q���;/q�c�D̉��q������=s˼��_53]��l�[k#}�����~G��9��*�ΰ~lԔ7��!�q2�'[H׊xn���s�����?�Ut���V����xp�4� w'~c�mۣ^��ի{0a���x����6��I݆���ラ��0lО\�um�J�	WID���!Y�D�'�u�K8�"��]gV��`�gmu��g�&�$�l��îP�L���w���{
o=�0Y\ۻ�v�~�DG�@{t_GT^=���Ɛ/ ����y�%r�g͢�-�*ɱv^�b���Y/0�Y�kA�q1w4^�U{ra��(��b�j���w�KI4�Y�q�wꦅ�s*����5���S�iv]�t�r�ږ�Bk��=L��^��4�FZ��H�u'���|����2��_��f�Cq���>�nqBgUwv���}g���>���EU۹�eL�:�$Fy��GL	�R�7s����5��o�`�|�wL R�^��L�O^~���u#pm�:���[b;�t�*�~�߹o��.�r��c���7����c�����4e���jUʺ���Xv�rcN��-8�<mlO��ԑ��xjvǴ��{G
��>��7�e]�R�-6��!�l�Tm�VrʢQ��e�F�Cy��l��v�\�z|mt�i�E�7��kz�>���*<}u)����1��H�[<��`�%���ѩ#�a9�j��V��]�"0H����Nmԋ���������i�������-p�3���o�����U�'�NY|ݑH{N�(ּ&f���N��af�ѝt8��]<ƍ�������:{�vE�}�vg齾�n�g�o6�����H�������ww��r8ÌE��\�˩�Q�j�N��h׺��Ô7��v��Pm�����T�.��ϋoW]�RX�Z+��#��}߽�Q� k*Lq��Sj�a�z�Uv?��Sw�FCh��-g6�/q�>Ϻl�q#@���a-u={5P5��Ʀ��y~Ca��8�/���鼣y�WDD��=ݎ�zS�V�E��Y�V��\��S��k�B5R4�OV�\�N�W�3�2��dƖi��G6A4�u�fҹe{,�ńZ�6�n�L�
j�̪��u�zK��j�Ae"��J�֏]�K� ��_){51�L�r�� ������ ���ځT�JI]�N��G94i�T5�ӝ�i������"�A]7��b��mH�9$�+�@g�Z���Ea�Ź@��ўUm�s���2d�c�17�we��&��e�Y-��s�4��$�)�5qw�,ܣG��K��	7�-E�fB$ɼշh�

T�r�Y-��}��`�&ˬ�ۑ$�8+gk��_)R�Nt57�	q�{�Gb,k�{��vxʛ��-�}���������Q85N�<{�RV�ˬj�up��Q��I�8�a�q*��2ُm,��/W�^�j�Z��W2�޺�y\8G-�A*<m��Y����w7@-���'�<m�@�����4%>zOU,�M�%��v9f��f�Ǚ���-:۪�,׶�NV}�4ٕ'f{�ލTiɺ�K��n�AF`^�0g���'}X�n�s�l��k�l�!�w>p�tv`�4��\[Vo��T��葍�C�\��kl�"�m��p#���هs,'cl���{���ݺ���k�u��TgB/4��������9��:��s�+��r�z1M�CFG<��Sݎ�C�v�[T�Z<�Q��1�@����<��U�'j�	��is;���2��"C�<5" i�Yj��ng�����[��v�kZ���Ub���œ*I�
/����T��=��������@�R���Q�j�.]�����;�*�n�h�,�_Rp]�F���f��Ԋ����mn��Y<�dl��n������j���1G�����ݥ���/C3:��OKt�a4��.�C��)I�*�j�Y��!-�g|���v�u5� ��U*"������� Ȣ�P_����3�Nkޯݹ�Ju�g��mӈ��SpW^����pYh�bot��W$d�IȞ��c#K��<F\�;�sT�]��x�g@��REϡ!���܁MRMV6F閗M���ߺ_�U���8x�O��T�j@ܷS�̑tB܅{m����K����xU��I��%c�R\ty��CU9̴�t�-p����{�\�~�OVsI�i�p�8�*MY�nJ����Sෞ}����}9�W)f`��;'8΂s/�@=��#�xW��J�]J��%�'yҟC�g����)�v��<L;�5����uZv ����]Wr�x��(J݈M+��Rʝ�Ze��`�a��\0��2{Uv�T�d���� ��h�x�=��w����{}��!���z�^>c����&|a�o�n8�Y\)�!���K5��׉tz����g��K����t旘^V��Vt�)&�O/#}>zM�c;|4u`��{�_;�e��+���g�yJ)�QC��&.ٮdu��N��8 |%ߩ�}������*hs��\U6�o6L��M��bP`i'AwM+�	�:��=�GD�Z���wF�S�Ao
ܝg�U�@m���o�{�iZ�nWT��Cy����9-T�"��֙@��xX���9�m<��[��եXo��:�n՝��>�Ml����Tם������~I����|%�����h�q0�s�=|8��c�{�]����4�/Y���v
ۧ�C��������5o�p���ӡ�9�L[yg�rW|0�H㴬=簰xvѰKo�S� ����e	�����w`n+�r'dhWV��1Q�c�MJ�Y�	92*�X�v���׋3z;��R�� �W_���-��IڹKf�}/7u��2�mL�c�P��ڵ�S���n�(��(��W�Z�
E>���8s���n]�z�*����������r��rr�yN�rçv�����FΞ��L�ɰ�}։���v�p��8<%`E�k;�®��7����Rh��������j�l"h��Ŗn���}��^
��֐�}��Ye)ee	w;�V�%�£�pUvop�V����0�B3
�nʕ"�������.υ_%pItՖ�㊻��XE�j2
�V�����	��:���N�ɾ(�()�W�{cRI[O=���Y���e,����,��Җ�4�Ҹ����<Gj�F����ŝ�b��<�R�&!j������n�B�l7ۻ��F0������{���R��ce�㈎�{w8*f�c��>rx#�*Z�r��(r�iK%J7J�k�s���͋�B� �r��u_]"6Ƈ:Wv�L,�7=��w����	F��rr���l2�r��Ә�IޥmR��t���m��wP�[��:�v�N�*vV�F^��jG��y�ĭ�e�n\�֓�_(��x\�eY��e��zG�!�L�l�ge���̨K�9�:@���_����O�����W�lw��7ȳ�z;~��Iqe��I�s���tᨾ�Bh����K� �=ۥ�})�Rq�wȘ-_-B� d�-�Օ�뽩|�#��sWh���y���6[��=ҹ9��%c�.9\�����/���_.��S�F6�����ɺ*�_3lY�>�^L������[!�6�v�v�u�uY¯�3w�c�]L)�CoB�8���,�l�	�����'e�H=&�1y�I��Q��0z*������$�o���x���^��M����uشb����َ\L����.7�N;���܋��wU���$�UUG�5v��TTA5MDV�DRU	��.έ9�+X�� ɳME2�4h���h��`ڭ��������3D�ss�����E���ƧN
X����g&�L���IIW6��u�(��(���iJ6�hѤ��cl�QLV�Uö��֔���LQ����h�UEU��X*��֋eѡѣMU4F΂�6�Y�)��`�m�m�r�Ţ���DMD5��F�(tb+���bآ-��m��}�9�6�QICQ5MP�FN���@��LT�8�i�UU�PE�KA5ST��Q%IQ�Rb�QS�`�1[b�)�)�����٦Ӫ*����*�RUQ6�TV	���1i5[d���J-�1��kED[�
j��5Q1IQLU��m%D;˟���_�z@����چ�[���MS�\Y5��	�R�yR�F�Tr�T�N�1^��2N�.� ƽ�*�rz�uM��A���u-�5��������:�=c}�+�7�8�\��#��␮�toJ8��7����d=ѽ�Λ�3�Cp,��&/�n�R�3�wq�����A��yQ2G7�&#�WN�s���h���Bm�p������|�ټ*��ve���	ǉ8��tTy~����⍱�r���e�u�G�^@zJ}�W]y���w��y3�Z��2FUR�f챙P�)��!�b�V������츩�[�g��iv}Z0��mr@�;�<,� f�dә|��-�%`���z2:i����/6�3�cK5v�)����'n�T�y�ճ�nM˞�*B*j�f>��n5.���j�I�"��n��P&�:���fly�����d��dA����R;�%~.�,���<U����o)dq���A#x:�t,fs�{И_z-V�
�(W3nM�]bGX�%���]���!����nm�>HwM�Gμ�ff��O1�ʘ�}������ųW��-���i;��cIg�5�WV�p���r�W��$�e4���9$y#���$X��q}R���
o�@��#(��*|��Fev�DEp[twv;�^��Mh0>�Ay��{�t�skc=���WNe���;t��m���VI�2T�kly��_H`�<�tlF��i�cJ��N��(�̌�4�G����� ��	�wP8��Lg7���on����*�5E�ǃ?U��z�-ל_�*R���d��X����S�x��w��2.�$<F̵��I����jqR�ds���v�Lt��#�6ǆ�D����[LTH�N���Kek�:/���H�c�z�g����M9m���Wj��G���N�m�u�"�ݘRC�:��i!���e�w~j��ݱ�*N8"���"3[�3�k�y}�d3��"� ~IWM��z�"cDULod����c�׍�_	�Y~A,�l�ԭ�c��D �������y�g�� �J���ͫ��Sۃzc�ٵ���'�u��Y�ssv����I���s+|j;$	w8G7-P-�����ʄ����R���V���e�����CGX�g�B��f��a+���h::=U�G� u�7���V4�#�Ņ�����{^��2ܩ�=���jV>J����+OQ�*����J�:ӛJn�l4�7�;�Z�p�<e�5R���D�6ʤ��E�j!^�Ƞ�R�OR�{2}sNf���=�K��/wx;[��;�!lƐ{KR�m@��)J�$�SЅ��j�i1:���L�a݋���jR��@.9ȩ�T���;HmH׹�� �H|�3M*�x?\�<㌞O��Χ��ǝ!�NX�?t$�8�~�������_"��O��H�r�'rCf>�y-�Z����T��GGW);�}KS���Jf�T�[-��_'�T���\�����9�^7�9	����uK�uG��̛�:���w�]�˱����k�3z��_��z̳&�*�--YV����|&}�'�z9Q���P�Jin�T���e��%�����6T�u��[���QAM��N��Z�WP/�k�uW���>;͂"j�W�²:��5��d�h���u��6�9�,�MP�2^��i�Άvl
��n��׏QK�ڻ�F�b�Qu������.�HM*=�e['J	���s�l��^�����psou�R��Cewu�:�!�ͫo\|%�G'��N�'{3��|*�\� |��0=/��Y~�:�wl���m߮x�������m��2Gm��P:G4�	��u�$�F��Y���qOfmt�C�ni���Q%��讞�1��1/�� ��l�Te^�!��w;R�Cϻ�		y�r�U�ngE���A\�f;*�fK?K�]�F�o*��w��#�T��	���ٴ�r�⎟dz3{)|h{����j;�Z71�_�r�-�Z��� �P�%����4��&�-ͼ�cyRf%�F&q�����!e�@F.B�s���lœG|甯9�#�����y���0���(;����"��koq�Ll�E茫�GD��yi��P(�rMP��ۛ�!P�ȑnH[��Bsz�*�T���z0�!Ky�:9�IX�!.2+e��ϳ F_��t�uX�N���ƈ����ᳬQ(�G�Wo�ڝ��1�S�d\��MBo	�m@�(��ת>����<���Y���s/���B�yR����sQ���2M��y[�xGtl��|T�D���|�s�:����9۲�� ǲԚţ�J�2���JV�읞���״b��O1�||B��9�u�\g�����4�*�H��j��k�`]p��y<�,�`�KT�<��I�؄�nY��\�wʖF8c��#�WsuD��ݭ�*�8#6<o���ݦ�W�׉�rT��OY�.���X�o>� �4�W@doKu��oh�r7���(�
�c�!��u��ǲ+i'x�ůi�����a�F�!�|�&�P��G_K�*n�>>F����{��$�x1��t۞�C��VҊ|��-I�wx�Th�»�>&�lޓ{��=�m��0H�Ĵ��_�ؠ��#��6���Dl���9�!hϪXZ�����s�x^"Eq�F���+�������������_��j�f��g��<�P�rb�.*@Ċ���iW�����@�t�k�#��c+�MX�hed�A�ڣe��>;��o���V:1Av���|[QQ-�f��J�-���)�i�[{q�����4mQ�q���r�esz���侍"z� �%�'n�v��Jf�Ov]���mr��gmX�\�Vs��Sr;)�z���[M��϶Y
�A��O	�q�|��w��sќ����U� ���eg�Wd����˫g��v�bM��H�*��0�<	��w/S�&uB4O%P��ګ��(�hE�՜���c���z���9EpB6�����;Ǌ��]��Zb��Y�٩��A;c;�Ɗ�mO�
+�F��H�){�P9-���c���5��e�L5�
p!ۂ��d^��8������7t�	�Y�k�c�3Nj^���/���m�»�)�ldAO�|J��Tq;p/Mn<֮6�:Z�"O��G9�{ZA��XP��S�WNe
��0�Ҽ�W5֧J~�4�K�������Δ��҉��J�qt1z��}�b:���Ŭi�s���*gF�
��7:N�[#��r���/�؁�w�����{b��c�K��"5����& ����w�,��n�UZC�����v��u�+.�
�4���0Ӓg��F���Xf�Vo�k��n!��k�3��ג8�rTu�D�S��(�`�p�S
��\Q�ג�ɰ�j�k{Qa�0�6i��Ԇ�l���T�[y�&��.��U��;7��>�G��B\����%��b��3���}��/�tM�U|vq������f��Ĩf�ǻ,�q"����7[�l�g1�Z;)��:�j!�+��%]7�lgV��A�n硟f_�������D%u�<�{�h����Ndd��耂v�E2�����a���އ��ի� T\�)x?��;ƒ���͕�L�Er�K�=�\ՔVF�p�9מ��_n�.2F�W�AM(3�z�ٕ꺷,�/kM3M���[��=�0uB�v�]��ny����IO�+��F�q��ojjU>�2	b*�7��b�mP���"�g�4u�����6"���W�Ӯ�����}B��85H�瘺��z���)5�����ݼ}�&I��{�c�n��Z�7���>V}�*��̈́S��t�F������k��K9���sR+�����\���Ưc���U�����ݷ0Y��L1g�5d0�_�ۗy��
��:�P��]�x�Y����S�t-<�B���|��-˞LwX
�3�����fKǂ�N'm��<��S�~�h)ZA�9���T���-�
��jy'p�$�o��q�(���&���z�#䉐{�2ڕ��CR�U܍��SPõ�c��6 rvF��?);�&껒����J5'�yT�h��mM//c`�ʆG���r@͇	=�7RafJ�/�k�{�cdbB"�
-�n�ݨ	��}#|A�؍F���dYG�n�4�.x�kfGv3�^�[1{�t��=A�z'�6�`_, �[Q|���pѡj}��WS+�M�lh�f�)$� tQ��8�{/�����m���P�'a�k�Dķ�����P.:���g�P~��"����Gs:.p<���ƛI�P��zf��(�B��ޠ
�W
�[�-��i��~�yu8R�(t�����"*��*���Z���:yO�ǯ�/�kL��{)�]��c�@t�������l���8(An��Ҩ�Q&�ܚ1��X)�j+.��}�*'����H{",|����w�f�{;�s�	+j��#L�wJ�\^����tGX�e��;6��	rn{�/g\^�ٷ��-1�Z�krs��T�eF{�%~�jD��&p7 X���i[��j5��~Ac�t������	��}dӯڧ|w2}�O�g@�("�BB+xl̅�5]��7#�_Y�$��"�9&�>Z��n�vdH���JY�4��*Y�CU^��iP���}v8���I.l��l��5S���ք��+q�4,��c����h06ԫ���+L.'])[ϧc�3�M�#�u1�u;T�H~0������!t��W��U,]3J�������OU�F�#����:^�`���e�yF0};ճ%9���[���r��=:�����)�-oݞވ�F�t�}�Fl��`]s����eLs����Gycs=�n��֖�q�@�N���P�|�ޖ�v�p�pF��S�^����;:w���u"�b�c'�6@�8M8C���}Q?������n���%_\-"x�L�w�!Vh%�����f�r��(���-����3{�a:x����/Sh������2susn��<�?mb���c��=��|��9׉���нzM@��4:%��3Z�\�"�Nv�S��&q|��*tiA��k#0ej�&H�8�a/}��F�r���cb�4)�Q�����#����*7���n̶�7{��I���\Ǖe�@����y]���L�Y����& ������W��������WMeߤrm��Nc�$��V���/,�见��;����w&��t�.*�0�UL�ڨZf��s4�#h�)Y�K���e�9�l���=E�����Cn&�j �u�D��� ��$�\!u���SNf��
`_�=�h��C6����s��m�DG�ap��{T#@��T"����m����|Ws,�q͹5ovǂ�P��W#o�В���l�x��W.�uT�,�g��Li��8�P�-�pP+�F��V�%ClQ2�{׌�k��s��� ������Pd�S�p�vO�VȽ�'߽�����C�������{���o��������^�S��gm6��ȚKP6�(������Л<�.]1Pe5V{]�n�xq��LLW�Ue����:[��6r�j�Ej���VE��i��3mb�V<qrt�lP`�Bcm\�/%<�eh�D�<�;+��vJ\��2�^j�7M��Y����^c����.[l�y{�ߝ��T8TLhx9J(I�]\`W38KǹvKw�թ<]�',���懲8F��q[0y�E-��`�/��{�"���O�T�	��t�_Eo�<&l/uvZ�%�f�2t�.D? ���↞{�u�#��]�����0w�/{x��V�.�W�D�M���*���u�D�rl<���[���wX�!q�y��ŷGY�w�;ܱta]R�SH����[t	ԷR�WY+!�W�y�Ӹ��7S��5v���wq�VN�U�m{�Y6U��C���m�P�PP�h7g��`
�<Т��:^0�ȣē�I�Q�Ŝ���+1�)K�+"Λa6�ܮ΄�8�K���/0���>@��)m[TS����c2"�U��D�;E�ɲe���Jd�u�Ś���ZuL��.7��p[R*³�O�(�#H����e�,03���d͏�q�ѳ�͘Ů���6�k��>ëB� ]o��m%ɼ���s\�zM� �k�Il�ҲY������RmٙӀ���G����3Jl��\9�{�׺'j/rPui��'U�q��l����[q�ś�ݻ2����r]��ڰ��{����� �F�T��.�fA�D3�d��,w	�dj����r몖�L�0�#.�4��=0���|�=��}��L���t���49�aT�Β��y7)p��j�C�vخ�٫���(��F����j��:�:�o^���&h��t���;��9����Յ2+ހ�T��:��e�V�}��Y���٪sMo�D}�o�/��ڒ�?Ot�uxm�a���9�2z�r"+����[�+6zd�urUz�p�w�R��2�]����xv�����<���i���]�4�]�H��A�8po]^��1!.�C@��<��R��B���;=	D�$Qi�sz�U�bL��)e.G�/z���]��	�<�6�.j�2�ݖ t4N���\��ܮ�F�M�S����em�C%?]c���J̆<^7(���Iv5�ɗ�t��R��=�6*�+��o�Λ[�۔��L��CO����yY�n�N��{9�K<���m��ϣ	$��j;����v��o����u$�Yݏ�]چ�7fxr6��oηL�x����}�-*�tY�8�֧�t��byѩR�#��f�}��E�	�
"F��������D&���y��Aw8�!��2a�� ���*|�S���<�Qgd%�&4��ׇ����j���ý�R�����t�G��e���2�ss���ݚ����qL�E�D�4&��ESAi�T�SA�b(�*������KMRm����f��N�S��A����:��(]���Ul�5��m�U55ZME4��N�j$�Z�6ɝ���E.�R5L�1h��j�M �ֶMl`4�(�!�(����������Z(bZh)�hj)���1:4PSl�%Rv`��i#m�U{ښ &墩)��*����� ������kHb��Ѡ���h"��CD�T�R$i�(�b*��i���h5����T��i)4�4�U4TMDQJui)(�((��)�i*�AHQ�SHU,LE����3Z6�L���1��hi��� �&'H:��dh�"G���|~���BKP�M"K��'Ÿ~[(3{������;ۯ���9F��>(���jr%s�)N�gR��H.�gR��0Ykl��^`����$�Ci6SJ"�LD�%� Aē%�E"���e�{Z8nf�3�gLG��VQ2��#���w�7̈*v���E�+Y�U�[k����VUqF&�s��6��L��!��N�f~~�>��4�͵I̙6��|�ԫ��mMEJ�qyޥ��[{T�\�j���ֻB�ª��|6F��p�.�۠s�����H;b!��"�3Ӈ�hnu�!�1��>��ϣ�%�͈�Y"��7���2�ngI�.T�`o8]�Gh�Kp_OPmf�;�`%�Y��K5���ɶ�-�W׊�����9��l��h�g�TE?O������+7�C�v�>�Q��ͧ��A��ܻ���ȶ
�Z���Y�c�[��u���,a��J���Fj���3Z�-&�#�i"�5���-��ͧ���,��;��'����L�ܟ����;����AH�����{*�},k��QA�B��ο)�N�/�Җ6�x�Ƶ~�d���������+7�5�����z�]J��`s��u������VÁo��tO�/\���M�n��R�;W/�9���Xb#%��í#]3b����L:[bG���6�
���Ӕn=�7M,��;�mi�&�yK����b!���W1�#˵H{[!����IOl�#C6o7M�
�(�Vq�m��R[8�_��y���Çb��jGz��D�6[C���ֿgQ�y�vqU�䊚~�t�t��E�B����Ri̱i�2b/�<��j��B�N�����=�[1���[���rᛮ���Y�e硲r:F_<�T�Ȳ�Y��;O�.*���;�E��/Y翳���U��5-��/Q�=|�@�[=E#]˱���E��[93�٦�d�
�$Ø�:��8�&�)Y��S[q+��,����u�+�MBϪ�?��1��pQ�����+���mpv�CoM�]�ϫ[�^�>��ܡ[!�����p]~�j5�����p�#{���f+WwnAƝ��#��I�4��;fGPc������Bq�|��g�f���0Y�jE��)�����C�Z߷S�Zy`�k�.J�N�R����s])��w֐Iz�e'���>5�EＺ�j�Δ���Wu��U�e��Cy����]щܓ!�M�\sU�O�ś��hڱ׸�KW��ԣ7(��	�m�x)nsr��V�]�r
_O����t��D��S��g�+)gS=�{�;s[�r��~e��"�������q�)���喨t[�w��}ܛ{!Q�%�`@�{�bWSyU�˽$v�dH�j��i�Zjr�-�Vg3v��V�#��@�z��=��Z�������q�/~hƃǛ6�z�#�*�i=qQ.dagA\xX�� ,�Z/��r�䞷�<M^��W`�$�7�v��w3�^�����#�����/ML��5\u�az0�;'�MI.�xI"��I��n[����7�3�#�+����k��]y���m�6�7a#̒K��T��[ka��֖��X09O�����=�����nڅ�Šu�U�W])[ϼ]��/^���idf�p�ʘ!��$����!tW��U��iR]���Ɔ�8D��T)7�M��Q/^��c?^�]Ȝ{�6/k���;���=�yE<7��v���Ń�V��0�]_S�;:�$���z�޷�[�M�뱚sh�Àԗ�D�/��{ɹ(�ivm��s*�іTu��8��tЙ��|⽩��-ƭ�5�nX���rੲN��a��e3��09�oWL���v�pٜޖ��ʹ���C�jA$�P�� ���Kl��t�'�[Mx��7�2�:�z�-]Yͽd:s�t�+���nu����Ä����u�gP�M��7�|�:i�f��5�*:����(j�����	���|Ȣ�@h�Y���Z�S�R���|e�3V�$�Ż$���+�mk6��\�qT�/e�F�p��R���w���7B���'���T�N� g��3�6*5��}i��0S���w�ּ��܏^!�����@�����_	�M`�wri��tS��g���	5�1�+,-�a�;(fx��Ά�*���)n$�+�u���W���8B�#��խ0�1��&3B��ڧ�q��1�÷�B��iP�eT.�;w54�j�=>�{{���^hW�L�vP'O���{�Z���<cO����@�woZ�?��l(*���aW_x���K�B�w��$Ul�u������I�9gsjܼ�p�/l.c]K��u�:vz�{�r��C^�o$+%�ǰ�v��c�t���)���k�e�Ҷ�ξ�:���}JL��]�O�b��r
}�'�u�P�r��!7�&�I͐�A�x
�i# r��|dwJJ��K`�w9����V�a���ݕ���=9���l�ӝ�T%lpS�p���<��w�O�l�S��z��Hodo��Y�8�+�����R�,����%p�CVp��7s��D�>^?��$���V�+����v��a]�����b�x�Ƃݻ9���LVus�"��Ux�b�ϼwM��Lv3��bfL:��{���斫���ť#fJ�GJn�8;�҉��z`^J}�v��ܪV�'�S4o�!� ��F����Zal�|9[�v��z�@�I u��\��욑O�3���d\>ّ�$^�����/�468�R�hly�~p��5Z���m�����Hj��wFaD��8��n>ok/-!f���w���)�!��G�li>�����oY�$�-��e�Ҙw����`/`n�z�ר)a�ڤ�/�7���o'*�6Q�X�D�=���D�o	�v��&G�9���=z|��õ�N�X�ȧ�y*S��Bc����<�N��h�<��h�ݾ����ڝj:$�:{���(��?c�yt+������C3XwCKU-�v����;}��y|"kyu�	�Z=WJv)��d69d�ȿοo
G�n�+ٔ��,@�a�����=����\��	����#3�j��WMU*����#Vcn�׉!�ϡF����hЋ��5���!\'qLYh�T����e�3��51/f�ͣ��B��D�R��[P+�%΍�z{�T�������6��y1��X���ԁV� �p��U�ჱuzFS<����t���Ggi㶼8�E=��uө��[$�q��:zSD�\{������p�2'<��ץO%a�q�y$��:�C`�6�-Jm�1��tOhe<����A�͎���T��r��Vk��G���'�}�ó?9{&?܌~��������.}���d��lв��G�_b_(51�+sm��.�LL͆;uJ�U��]�1ƴ�u���L�;��ǖ���嫹���]�@�o)^K��6�+%^۩���M��?���5=˖��*�%*���� R�mtXoI��MǸ���k�kr��ge�����[�}!m��ۮ�����+�=���+�����a|��7�:�G5�&�rR)n�E�����K�����~����[�0r7���q����x+����,
{&X֌���~}�"s6H'�P���#6G;��ow�B�~�_Yl%	��$z��x���F[z���z���ݲ1��v̎��:Ǵs>�2�AϊQ��x�pѷ�E$z��G�_H��·��Ih��FGg�λC�jȞ�[Ը��w���z�B��	k͓��1�d<��`�4�G�,��v�:��Sw\�.����Dl���GW�Bp�dצj�2��#���*��a�q���Z��r�x��V�}�{	�%ꧪf�><ޤ��eK�ݑ7����M�v�j�q�7�j�GW\xTK���W �s�!nQ}YfpŽ9�m�V��Ӹw4<W�[�7@q&A��^uQۼ�M<M3�y9>>y���न(��J�ʺ	L�jڱ^�h��2�i�8��u�p��NDx�[�IY��tK�%	�}�1��.UF:zU���vʀc���V����x1�)k܁>��	�w����~r��R��ŗ{l�G1(`�1�C�C��c!��T����ƪW���tj��%e�*	.x�>Z��u#�3�Q�����m�Ў������ �b6�u��ΒV�*@K����z�U�,b��������l�I���C����f_��*�<�7�t�6��gk
_"m�з3Md���%�#�=�s���$�S����(T;�,�*�Q$k��n�of�J8�l�k�Y�{b
� ���OG�T��%�f<IIUk��-��t�m�#6��]�\�P��{��2��T�v;�2���Ԙ��{VP��J���`o-۵�����&�ִ��Y1�E���!Ř�u���ݓ���Ѳ;��st3�Ӎ��5t��ݢCE�8[=�<UܳN�$�"G�L�,w��Yʣ�6׳�]�M	�T��Ȅ�,�xTk'}��'2�=�xG���)������_D���C�P2�18D�ߚ�i��vӞ��D����[Ժa.�d�7J�^�1��j)��Z��ei�rTT.��f��7��H���G_�m��碻�U��.�^����������z��9_W�|��a"E�6�gN�v�7]Y)I�ms�tڑ;������៸��)��o�Ր�7�,��S횺��n?(/�z*����6l�i׺ �;>&��ɴ^Z��O�tx �]��w�2��#g*��<� ����7��!�JV%��/-M�9�l���U"�Ɗ�v�}�&:c�h��:��j/��B�R2(����[wQ.S��*����y��e�%���1MϜ�vػCrS���J��U4?j�c"��g���j��!��m�(~�;�2|ҏW#�m����%���Y�:zw�=L��|�P�6!�3Y�Z���|�Nv�����ElpS�w����
���H`���n�^QG/^� U"��Tz|��}�xm� ��eջ��~O�g'�CM�Ϛ�M!����r�����Nj����!�}�	�<�a[aw�r�ݼ�bp����ڮ��FDv��N�ndw.�q<�;���i�����s:�Ҙw��yv�Ū��G��ԥ�~�$�ow�3:��j��D�Ĝ�)������{m�|a=�5{��g[<�܎������4��7u��٣�|fZg"��Hyb�E냃5��i8_N���ގ{3=:x���{�iZ�M���r7��B;��+�f���0ϣ��3�@GO��tI�䴢f!�ݦ�x���sDl�p��.�0�]��#;#rw �T-�χ7�dv0��+�l�hOW���l�1���9����3�'ץ�|/��Y6xMf��us�8󈤛2{�g�_t��d;�.��f�u)f�t�'�{5��n����m�a)��4qcO4v
:��c!�hWD�]6��$֍��ގe�ճj�:jW�p���V��-t�E��=X�
�ew�������<���� ;��
���2��܋�jHO��2	��q�f�i����k�j+f�����]�a���,����d��f�P�Wo����X����p�{m�qۼ�Wv�i��E��.�ַj��ac.��5O����M�2�&y�F�z���8;������������}C�����{���w�����x����W��ٳ���=�n����D����P�4²ʼ���-��0��������1��۷��+^��<�'�e���UE�4�#�]F��K䵠������B��32�=��H������=�׽��4<�rzr��r��Ź.M�r칛��\7+����c�佁kw��}�,{�a~]��ǖ�]��,㐩�5*�b�쥣!�����Cb������L�.��;m���2L������9�KsP�����Y���u�7���'�>W��Omm1�s�7�m�쮂�{�1A��� �t�蕘�*�!˹˹c{Ns�8������	}z9e�b �})�+��ĺ�YY�!���܈҃��WJ<���B'
�۵�����lZ'��q�'�yg�g5�sޗ�*�R���ַovYǙ>�_0�l��!�K�C��,����Yxƽ�1vP����`#�D���z��k~�R�H�I�t�i��������R�"�����[s��}n{|Z�����n-���\y%���_����w��2u����<�4 P�
���u�	ǣ���"xr�����:<F�5�1c6/�����xe�M�^l��8Y����U�\�@q�7OQ�݇/���FEXh�`�Z�I}�ھ(�Ut	L�/(����|��1�I��HS۞SՏ�����enU(�;�i�1y�A����'z�:,�R�6ٺR���OD6����=''����Vr�d�D��l�)Ӆ�K�n3��<�]�V%q���o��@uL�j��A;f���ևm�F�ie6�2���.l>�QiP���%�&��Fʐ�+y������X�nݱ�pD�tiF�]�:�Tʭw٫����z�(�����ӄz���^Ks��_ f�	�����6nW_�^�yF��>�J[���oe5�֍�W�ͅ���TZ�l�R�!FVϰ�y�V��{YR&��v������v�vA�"�I����R���u�)]��>��]K.]�Oؒ�d|��YϬQ��R�X���!d�&C�:�Y;�$l%8ʹ+�>k9ͷ���7�U��e�H^ǃJ3zlM��˃���'���Ծ���+Y~(0��î4d�l O\U�1��g]��Si$�̵zșk��h���8T��e��8e������K�=���>LK�L�򠴝���ʈ�㋦���9#}K�7I��g����LO;�=�2�=n�g�<kT��hn.e����+���QT� �ŭ��m�׬�YjFc��]����ٕ{i��qC��ҽ����xV�w��X�mf1Qv�3�u��m9��H�o;tVs( �5��1`�#q����k�)��߷u"�aj�^]�ںUm��cѬ����5�W{���+.��s����|��s�펞a����#׈���N��}Τ����߿~�����nd<�W��QU)5#�KTQTZ�UIH5[e�#0�Z�y�TE��QU���(
���D�IJU-P��KD�Nڀ�ZZB����"��
֖ )�(���h���
m�,�TT�ƀ�t�H��Q�Ji�@j���
GN�����mKT[!�H���h�����Z�4eء���:)�"�JY�I�
Zm�C���]	�]�F�@R�Q�7��MD�rMFΔ��(�m��hY�*�C���@���@kTU��.*tb�����2HTmI�)t�"��lQIE63F�*"d����
cM%QAlb��)(�*� �
J��g�������7�|{��u۝�F ���ǜ�����J�H�4t���d��8��KF��{V�ב��J�hS#�d=��=��z'
���7ws?w�'�TEU�u�S�̀E�A�+��ছ�y�����=�8��];��JVܸ�ד �]@���6�c�]@v���7v��2�"�O@��v��i>��KyMr���-Y����vؕ�2Q�C��t�G�s�%�ձ�G\���Zآ��K��)v�z�g�S��| ��q��)�?�6@�dY�3�B8Ѡ����U�	�g�Fot>���*T�����y�f��z;0nG���'Z�mllN��֛�G��^K��A��2F�m��`7��sv#��'�H���� 5�UU����-�o���C���=��}=��P>|�ZA���x��M�X��
�����9Qh�`w�r�� ���h�y�<+du1�[
�!�i���F]���qx(��W�*ѿf��!����y���6�ǂ�6vFd	��佺�6ey����WH�Z��-�9ʑ���=�����{ڊ�q�^��h��d�[�� H|ƾ{}��$v�:}j�Rk噂�.N�:���b�)^ۻ��m\�Q۫�N�g%.;�	u ��sOJ�RvT�F���d�q��֪�s#�z�DFݣ77�qh��/�2�Z|�m3nʄ�	##�j��#²zu[��g�J�z�l�ȥ��S���6�35q�m�Y�y�u�H2j�A.Ɠ�Ok �Ü�8a�\\L������!��S���
�&���Tw3�^���=�rJ�A�Tըג#�ſh>B������+/	REK�5A���:	� Ul�mֶkҫ����{���(]�6ۄ��t�󤕷K&������+:,�w6�|��"�k����p��:\�m��*��G\�^<ޕ�KL��g��O��2��;: �'���z(0�@�n�Eq��ؕ!��(	��ET7���W�Y\�̈́	��{��<&^�0�l��\0X�j���&��p~c1ْ.Db��-����~=�귏+]�����>L&�H#6<m���nxC<��\��xY�9:x�.)�y}�-�-zyH@a뷲g�[c��vEϳǂV���oCe#��=�ヱ�|'�~"���$$���N�1�#Rse��/�ԥ���gN��r��R�.�<i���1yN�[���fHW���)ka�/�X}�WY�)����W<��#��wR�+@���Ǻ���doKu�5���H���oc��a3yUF@WXyw��i?NV�����C��ШL�r -�4.f���d0�l��P2���f�Z��&H�-���㊝��������x��/����3��,����M�;��tԟ�Uhf��/$�h�<0��p���7:ВLpN�?`�g�,�%{5uѝב�2+*�n�=Ap�s�D�v�&��<�o-OE<���H%V�~���W_�F��jT��^'�qxTKW����b]m"����0-�F��v��/=�����x����s�ȁ�B�<��FS��l�۹���[��+�T����[��s��*�ɉ�rDyvػCrV��'�vS���Uճ�\�`��ܬ�O�s���8��#)�F�o��JK<��iw�S��QaW�K�#g�w���Fr�<�Zڬ��u�;���'���]�OM;x�7O�Z��)���{b6���ʀ��F1�5�-�WK[�����	@RV&k���
� ��&[/.��,&d�on�4�57AJ鏗m�`�m�ÔU���yq�=�.M�aoQ�����u؀�; �?P~���:�������TT�U�un�2�{��^��MW�#z�V�*��*B����<]�6���]B��k��t۽B���z��ؤ�0WbskcL�H$L�q~�f �m���]��|�SsEOe�&9y�쇠c"7�6�g+����G�k�����}k�V�f�g�c�Q���q~��3Ƃ�Q!�T���m^&��+e��h�"sՇ�&\ݯ'�*���_��@#�x8�j����ͤ]n����ȭa�++C��m=[j�Q�����g���#���,�������	��i������槪���[R���mX�,~��t�B,���P�
���];��s�e��;�8���~�u�����v�|�5Z�Q��tÿ�j5�yJ��⮐��=�JОE��^�9=���Z���<��]Щ�BqS��e��)�r�ph֮����ϕ��B����e�ÏJ�#���'A4{�Ɯp��Gg+J���}:]έڽ�߯_��p�g���ɞ۵�<-���Np¦��X�*\Ru�}a���)^�6z8��۸2�h���H��IZ]�Ѹ�k-Ǹ�o2���&�~��7"��R+�$�ZQ�)��k�`53�Yw��ە8j�`n����
�����k�q�5����;5tS�Lz�x�i��9>� ��C{2ni��`��Bx���MK:�3��ޞi{�l�Ǝ�9$�ueP��v��[��[@2���EM?/"���{��]ìh8NHn$�<D�T
*�?Tuө��������*ܪW�%۲�r:&����;�%mˍ{^L�˨��f;�@�Br�SRҫ��Sз�! �.~b��Wd��T�*\�̛�5���2-���}f�w[p�ʕ4ּ����#zveuz:竱L���RP9��u�ųQ"�^&9��\�]�յǴf��:�#fu?,MK\D䒸d@��z��{Z}����2T�����|���q��Q�#GO�����k����.]U?K��<�Ɇ����vh1
�gWٌf~4χ��oY�ѯ��6մt;H0k�j���N*���d���_A�6�@�*则�3�cįu<֔��2�w�egq�b6���N��*t;W�Z$7���9&;�������z*�}[\{��`vH�A�����uB�P�Xe�8��sf'z���oGH'�n�(� _eW��l���t��=A��Z��z��׷�h|,_rM��P�
�����8�i���>�n3�Ih:(�l�ќ^3f�-kG�k3��B�<#>ثF�w�wp��N����k��~���ׯ��ee�c�CE����5�4&j�.�G-��w2���^�S�ً�=���X'{�VI���t5�`bU=S6{�T�;0�:�u��V�X�����%מ}񋊉s# �Ý�0^�\VJ�i��aWhq�&�A9z�ч���$d�I�:��ϳ(u[��rl�`�Z��z������^3IG1�+H���JK�/	$S�!��+ʖ�lq�&5&�a��:X�gy�H	��\�
�p�mǺwa#c$�7J�o��VC���dh�w���v��I���&(W(|��
�do���zכ��u0D\E��<�E|ن/nT��z�z;|BBxˌ�E��Bsw�.��#����t]Mz�ƪ�ԣ*F
\�aհq��ڻ�.�d�:x��wF�n���''L[v7�5���p�^��(,�V��9`��C��~��2<�t�l{lʡ|[�
�3���k���=MJx��U�n���p6N�{)���e��}�W�]����9ߺ�Ői��R�R�����P��#���`�V�n�eT�X&�M�^��驊ή|�8��u^Ǖ��Jݓ{����a^#6%ƺ�fr	�D�����7(��i�A��=�(q�r����ng�f[�s���wjӶ�y�tp��Й�`8��Egr�u#I�r�FOthn޾�Mn�N7n��^�bM*�.�f�^Y����H[�d���XZz�1�aX��S�n�8����ƫY�x̿���aײ*߳N���v���E���̥��f�D33���܈�%�^_}Ր΁�,�zJ<(�}�w;�q�t��y�zм$D���h�<�o-O�)�a��p�:�#6ʔL^<	͓u���QqB��7���,]�;ჴ�HoBO������l�^\Ki0|�ߣ͇s67�(6��{����u,y�p@*a�4a=��¼�±���s�K\�n��n�w7��W=x�k5mϞU�Ý|��bօ�	5��8��T�{�l9+%)���c'�qS�R�(#J��[M����Oa����}��k\��p��\>�xR�YB2;HU��V�.�#f�2/����7����4D�:�k��nM�"�aغ[�R5B/%��h3Qˑ�k��Ns�P��T�w#i��W�uǊ#$Jp"�Ry��#L�FN���Duf��x=Gd��?WHk�[^pE@�����e���yql���8�IxޒU�H��_om��<�t�a���1��a�]�i��ީTq<i{��.�H���Q����k�!�Y��f�;MTń}X���dBꍾ��*�(���~;���aȮ}|rŔ��{{*<1��r�8[�6gUGJ��C�-������76ଶ�sqp��j2\I޵��~�6
pD����R\T��㆕Z��l�Z>���"�� 6���#��z0K�3�9��]Fff\��.�|����u�x�`{�����]�e���7c炣��?iI�e֜��v��wmW����m<<uZ��$/:��!uV���I,2085r]��c�x.�7�m)��;_L5w����L����:A���ͣ��q�̈�YM9s��Q���{��F_ξ����� �m�v���Pg�o�uř�E0B=ٸO�e��p���m�vZy��<Xƞ/��^�].���t���g�*�������H�]�5�yF�舱��y��'�h��Z���v��X�0��a�!3�*�+�X؄��U��;"�$6�$�%5�[ڔ����|{�t=��>���n�@�.(+���P�dЋ��D,yj�봟4�vg����FWޟo�uZ=w���2( �M�i9^�+�ڟC��_Z�ffS�ܮ6� ����AT
��#)�Fx�܍WޅW��"E�NE�� �Tj�������l"�����iF����U⊪��G]:ӹ�l;%u�V'����j�mZ�(q����Ӂ���)\O����Q�(���ۚ�}e�����1�?]��y�3��Wg�d� "ʈ:Z�]A�c��и��/��A3��{~�;�xhD�'N3�� �Ю-�m((�k�T�i
1Nƌ�}G0*Fy��S#[ǧu'���.wA���P�ɖ1�K7�]^�oIҦ�����-��"���܃��n���J��K��[s����^_n*�x拍�;�v�?�&.�[�����^��������9�݈�7lz뷆�6�C2�Ib�]� ��[\!�`��26g_ʧ�������P����y��[��I�Mގ��@���a���C���2����L,��0j^�t�;G���,S�h�U�^ռ?��?j!� ��M�4�mu�V���Z�
�{�z�_eW탼�{k�u���.P�{G߶f��7z�8g��%+à��_Df�������`���
�����Л ���6�(���T�b���;����Uy⶯/iP"�vtd�;��9e���O�5��v�D�߳/����P��UVU�4F�ո�F�#}G�� ^џvۗ�`�z��_����}�w���|=� U��TE���y��D��@D]�p8p���|O���U��0,ȳ� L0,��"�+!
�2�ȳ*̣2,ȳ(̫!̋0,��
�+0,�3 �H�(�#0,��*� L00,�0,�� ̫2�³*�+!� L0,���(�2�32,�3 *�+02,ʳ(̋!((�00,ʳ̫02���2,ʳ� L�2�ȳ"�+!̋2�ʳ̣0�ʳ̋��<���i�fQ�dY�f�`e�a�A�^2&� /%P80��Q� �C  C*�*
���
�C�C �C
 C �C( C �C
�C*�C" x�� �Cx�U�( C
�(��0 0 2��ʪ��r�0��ʪ� C  C*� ��0�2����  C( C*�*�0�0 �+0,����0,ʳ"�0,³ "�+0/0�x�2���� L0,ʳç �̋2���� L0��� �|G��||�����EQU&T@�?��n�������~��g��������?����������pǳ���Sg����<}���~H���~'�����<����}$�*����D�������i�����?�( ��7��;���~$��>�|���������~����AE�Uf@	A�P(EeUhY %UbEV �� $!Ud`@ RVP� $UXB@ �IUYFP �d RUV@�P�  A8����?��ܟꈊ"�"-@+B��@�������������`~'���y�
�߃��~�~��?���O������X�/I��O�
 *�և�'��ǣ��OP ��� *����C��C��=���@}�Ό��*�?w�����|��^��|������p x o�����r��x��@_�=��6���c������ϼ<z�p>����pp|�E ~?i��?��A@_����~(y
O�zy����`����~���>=����?��( ��>*f~_��L����?W���^�I�������|0`�<�@UA^_�����<���C�'��PVI��q ـ��` ����������ϰj��% �T")AE*JR��;�D����-�
�Pو$iCJ5�mUBH�*��M2�U*J��J���ikYh1)�����]�'��$�[4c6���C��j�oY�Q�6�6٢ҴI��������l-be��b��bU�UU�����*�+�WݝV�e}��Smݮ�͖��&m�Ѥ��6��Q��V�d���YB�Sd�FY֦�մɍ���Q��-jF�ѭ��P��mSU�Y��ͭf�  ��;�گ�nݳ=OJ�붦�=��6ƃO:���n��=w^��n������Ý�z����6���^��{֞�ޡvu�G�w�']+����E��e���d�Ԋڴ�j�V�Z��4�|  f�CC�hP�����B��� 4/�S��C�CB�
>�����lhR��޾�:ݩ]���w���uӥ��qզ�v���YԡԚ�v���v��ޅ�3�y{�[�*�K�wdi&��6�2��  �׍�;��z6��үaB[��:n���b����sZ�9]���Oc.әѥ�u���r��{���<�at���V���{hrμ��i޽δ�����{���o:��J�F��Vd���#l� 㽼��텰���ww�W{�4+�7������{�ZV��e���sqv�\���kt�{jz��F�ve���{öJ��j&U&ƫ���ӡ�f�N�[z����Ql�mm�m�� ����O=�4�՝Z�їU���
�-�
ي�u���v�j�M� L��w�7r��CA[�P+LPu�6�6(�f�I�ET5��   ��֕M�����C�U]iwwiݭ;��f칺º���k��:�h���u��h읶�]sۻB�D�m���%Z���Kͼ  �FZ���op���y�V�QJ��]��t��nsG(6����MQT��P{�� 駽뽭��(
u`� :�Z�+L��ƫX *��o�  ����p+����< �� ����p �����ӠSۀ@9��@ R��+MR��ݳ�@�����[IU[UK5MV�h+�  t��@�y�4��  �n� Q�q�( {� n�.r��  ;�`�(�x��[ުހ�4���ѭ Z�5�Yf� O�  s��
Py�` ��  ���N� ���  )�{� =]��  �3� �{��= 置� > �~@e)R�h0�Oi���F�di�M���%*H=@ �!��*   � 5J� �@OT���U$  1?������������l?�O�63+6g��!�8tL�Yg�F�b+%nA�<=�x{ۗ_����z�j����������[mZ�ݭ��m�筶�m����[_�������]�H)���$���qMю�÷6ɩ,e�É^n�DlG6��33v$���sZ�V]��/%Ӂc��7P��w[����wr3(�BgE5t*cq@�p�ڸ6�"�bݳ6�GK�����^X5*bjn�nD"Y+]Mb��)X^7q�qhrR.�WKv�O����y>��rm�C>ܛ���ch��E �eK����I�c�uZo1�%G���B�d&�t�mXu{���T�4ܕ�]cJ���#Iۥ��X�,<B40`�3h����fUŹ(V�fٷ���jɸ����X��E4ս�eLJ�Ѻ�a�DK��i��1�بF�Z�.��GH%���YXnaT��Ei��)b�&� pEBӤJ�j�Jj�SI����n���q��"b�8�%�v�fmf�tB�+Kb�y�uzF)����D�ɵ�b��67J�j3�]e�l:ىl�oN��t���!�T��n��F���ڠ/Ի�
c̖jQA-6�Ϛ�m��KX当��v�"�\:JT�X��U��ț��2�m��KV���/B�*^G��Y��
:�V�5����p�`��N�^�.���vɳ�-T�y�	���,�q:� ��&x��Q2�Qʶڭ��Lj��J��r�
�7�d��A@3��`��V-�#rVT6��;{�V�m�V����햓����g#��OM�Y:�P�.)P�M�Bo������ou-m��G#f3M��Y`�na{��p�>������,*1�	̳N�g��T-�L�%n�Q�iZ�T��4HJ�Ɣ�r�;�b��}be�"T1��#�5�R��c&�FR����mA�@Yy>��FHՅٵ���� u�S�g�V��$��Mj�"DZ�%��j����r^��j��)��>QV3PiV��_ۊ�u$ܩi��ޗ�-y&V$Ћq��wN%Y[0�����ƈ�E�XQ��s%d'EYx+��4Ͱ �Ux�(Got3a��p�&j�M�#�`�;.�H�ܴ����ѣ��떄� ��l��@E��[6`��m7Y$��Ԃ�n�Օ.�̦D2��&���4��w��Ri�*�2J�+qa��ޛ4����C,۴1���EX�r�[J���f����Y�Ill���n��E왖C���XyLn�X��l(�S.�F%E��kƑZ���D���˫��a�j�f�j�6�GLZ���Tv��U�ʅ�B��W%��%���8��-]�6VC&mF�x��]]��0�FU�zS��l�2�.��[H�wU���#.ǂ��^P�"�'�^�����4�S�X�($�J��	����&��<E
s��4�K�2�HT�~5��Pn�KM��`3��I�2��A�Qk���V�T�h��[X�v��+R�L�n�m�ۏwn�#�hm�[O#��h�%�u�F%�ŗu���^�p)�5��ϱ�O�G{515T���nV�٩�#�Lj��v����IE��`����4�iRA�-&�s�u,h�*��	�4���le�u�{+���yX�\_	�5ԧOS�{�)��e�ϚicE��]�	/$xo]�e�72��cq����f'��=Cn-��a�������ѥȆ1n��޼�y6�3B�<�˭�����֞���AF��3�h��Px�aʅ`1h����c� �ّ��;@(�;j��"Hr]���b˴�۫��.,�JM�J�fZ�~k��߷r��LU�T�ձָ2��ң�H	�t涷]a�ZԱkq�)j��cuD�e`U�$*Va���5ʔn��i�U�m^���`�Q�\��������Y)���+��w���l]m�+�V乙O]��6�%I�;�=.��*�I����m�%�;�f�3T$nА���a+��r����E�Ĕ��+D���tv2�l+�r�Wrl�&�� �'+v����L�����A]:�Y���&�&� ��t7u�mj��ɡ���J�@D��ó�F�X[�����`�fI!�V]���U�r�Pͣ+E[Hl��,�%͡�v.Ԓ�آq���A������f�2C9u��ڳ�a�鍩���Fi�Mj��.��R���<ʒ&�!�i���a�!�˕(PT��:���K���u��$�0އx��n�p)��Kn�����F�S��9�c�-�n��X�I�5��v�v��2��U�ã<�N!�F�
��p'+f���i���YxM��eL
'J�2
�@�K�oG �ܮwP���^v�ʤ�o1&���7��.J��^0M��y�"�8��z�MI�U��A�h6�
�F�9SYhe��fe��j�Yi�X����qQ�󻥚�	��,�19��
�fT��T�i��al�����mm'V��Pb��2�vp��ԽD�x��b�ʀ�pv���QҰ�r� �"�ݑ�%Y�W�Y,ǈ�ՆL��d�U�F��Wm�r$(�&�`<5��8^�V�.G�j�G�Q�v-�3o 7ML�Ljd(�2kO�&kh��浰�D�R��R���ɒ�
�"޴�kcFԵc,��z�ps: �2�Q�:�򜭕���S.e<M��:K^H�R�ۗ��m뚍;i�*�n���3���){X[�ͬU�d�)]�0���}Y��[hJkK	˟9L�eEt�[��5������K��(
f��la'5�݊;u�k��6���N]����kڐD����[�	�M�%��B*�8V�b&�Mњ&U�PV<����!�oeF]����Z�P�)R{F\�
�%�h���zw%�{.$�E�)[x��`Y[�]�WAMa�["�zJ"���B[1#D�wB ��N=���ʓu�/$e�����{�N�k[�(*�77S8,�FԀ�׬��K$�b�2��q����+2)���kF�f'Z4��]3wx�i�jg��*�`��JC4mj%�wK����a�բ��BD!�-�Y�C#�d��0���{�^�gLW%�Ժ�>�4�]-�"/�0]:��[�E�
�܇�1�JzLx���2�
�̼v0nTߴ
L�i�>*<���m+6(����l��Zp�I�y&D4@�Kq�n��ǡ1�21{IF�#aj�Ef�D֪s2^�@̊���qH�;7z(5�ړa�RB���7SoQ�X��d�)Zեm�rm��aw%N��)^f��\̹�ܽrS#�[V�7���[�OJ1-K[R-��L�+-+�u�˩��y5����с�@��ɬ���w�b�ŀ�c,�hT��0Xf�v.�.�x�.*ծ��B�E݋���i�ЩTgs�N����n��<Cbt�Ҧ��"�pL�L�Z�\I�ˬ��N����Vg��V�f)F��Yg0�w��ԨSh�y�94@@��w��bGfh�oJ�EX�����[(�{"�"�J$��tm��e���c9n�J�|�j[V�;�1اx+\H�w�L�b��Z1�^V�9�^Kme#�M��u�L�2��)D;���a�T��:�cDz幙�%U���]�h�"�(���6�8S4FR�e��St�j�Hf�m�o(���4�Z.maL�Ԥ���ӄݬ*F���!u���y���A\�F�wv�x�6�/�Y��O
����*X������߬
ªp���6�A��p��I>�>w�w1]�q᫢�o!ѳ(jٖ�k�Ym�Pڵ�������7�2�BӺ��76�x'Ɲ�	�	ujyD�4�D+�w"��$b3ա����ݱ�Ċl/U���V��ף����lJ�������HM%�Sb2̘.��l��,@R�R����a�VD��,�|��erw�9n�"K��m��X�bzn,y`�{&M�g%l:�,yxwB:�{v����n!S.��n��&��Yz��
C�w,Cp��M��7�R�2�nJ�_�
�~���!`2i1�j�!�#٘�ۻ����'%��.d �ŷx0ZU�I��FQDm��|�yɢ��W�¬���u���ä�p��[@e] �56�W$p;�,h��Sm��(V�ud�q"�s�6���֯���:�j�[ܤ��\Z�(/n�ƦZ�j��T�o-�j�*��R���Y���s#���u��&��?Mq�#j���OUbvIǺLQ�o/t}.
Uj�\t�$�M�t3L�cq���@l'q�60DIn���unG�)f8��iҗ�
��� d�����gcpU��;HQ����Z-ÿ32����fM���j�T>���5�ٕ��m�L�1�wY��jo���7"B��@���j�An���)L�j킷`���cJ��	��hU�F�O���`�ݠw37� [���s`B�(��]�*�(�B��U�r��2m�&Yp�.���u�w7�̩N:�,ϕ�1��w4�X�b�*���U�ɠE���B��X���aȲ���e]��j�F��Xuf����qi�t��'�����%.�,�����n�V'�	7,@]�t�#�f'Mc6R'Um�F��������,ؖwql��BE\sYɔXҔ�X�҈������P��q�HaWp�� �t�t���WSy{7�h��Ah欴�ܹB��&��rkr�x�Ѝ�#V�z�ӪS�r�#�%�2|Y�t�9>�6�˲��X�:�,�ա��	9�� ˂��4��k�+iX�.�]��d�A!�f�A2��CM�y���P�G����M���m���Xr�a�:�칚)�V�AX3�y�����-�=�k��$0+.Gt�(љJ�egңJ�p�r�h$�ִJ��(�����nʄN�MH�8E�kb�Q!=&�,����8�H���B%��,De���kn�qYa�Ô7$��ݴ�2��/M���z䊕 wU�߭��Y�] lVL�d��3DE��6Ĵ�\��`V�o�-�,��6ɲ6��f�$)IA�Gn���-Ge���8��(=����1)�i�ݘ)m��-+6n���a�����'DS�U(�GI����M��	ӗR�hס�%�"�~��5Qn��P�B�����q;��4}>Q�Z���Z��� 6hX�#6kKec�q�5��ܠ-9�%Y�[��/�Oip114n��&����6A�����a�m�;���3D����)��[%Q;�u���E]�����U���-c��/�d�"�g!�{��k�8 OA�(,+`�R���g�3�IK��T���Z+���K�[ݚ�I��A�r�ʖ���\ۭ���ܒ������Sa����[b��0<�t��%�P�n90!Z�֚q�QY�LZ ��R�b�1c�����,�jLW.���d�Bb�yi�X�ܹM���,n������-.9]T>*���|y��i�j�Qõ����p+��oU���o>čU��c\�q��u�uelR�K��f'�ZCT�)P�B`项�J�U$]
s*٩�e#SҤB[�����dT��U�hflX��N�-��$QH��NLu�&`�%m��{�3�Ik�s7f���t���(-�U �X2J��9g���/J
���S6�LP�q�b��10�(�@ɊC��5�yhл��c,Y%J���x�޻�aEv�+oi�̈��ᱍU���E��\��x*�Cv7"��ե�~[���2!��֋%�#E]a�0TC����J�f�V�7yx�"���R�2�c&I��F�T�6�2�ɫK��[�RR/j+7d�Yq�)�̉��:hbȮ�9��oc�-^m�u��ڢe�O�4�6dyWIY�R�^�]Fj:w,�[Q
�N��e�*Ske��\j�Z��Lm:��T�t��%7ncsksj�2�n0Iz�͘q1@]wܚ��Q�fL�n0M!f��p�.�vEFnL
K�h�����*��&�za�6���n25*� ��0K5��Vu��#1:��5t����Q�l����  5H��Z�X�d6M��@&��;�n�[t��� ѷZ�Q�p�*���p��L+F`.�6]G��͡Z�w��<ef�s�!hěE��ն��X&���d�y�NH5��b��&�tޖ�Sf���*)��mb�
$�����r�6�ڂLL��s]7�#w*�ܼ�,����(J�GK2@�ۥ��L�0<R�	ģ�YW�P�����gĩN��v�KÉ��b�J�m�5흼X��XN���I�icn-d��Ѽ$俷̒�y���Z�b��M%*<��7�}�ۻ�``^�t�-6٧C`���m$rl����4/�8ڵX�Of6�P.�%J^6��)<۩g5�r��Y�V�2v��mX����%�Cr�#�U�ȩU�ܽ�ʷ��v��/r�K�&	��� ��QX�Om�F�M2�
Y�DX���e�j�'!MG�5�a���N�F������F��r�t��V� 2�eR5�U�����^���k���*Q#�B]��CG��e�H;@����fʧ�I��^$���]���sm 4ַB�ì�Ð���ɕ-I����1}�Ip�ge:V�R-�{nޅ5�q&�����'n|��Ơt�q�^�cGdT$�);�7e�IYf�.P���Ts(�R�F����H��=����P9�[v �cS�YY2Y���)m�u�v�6�h���_+/4�AxFU�
k��=*Jn,Nd��A&�b���b����5�L� ��Z�m�VQ���圫Ѷ0���7-7�m�y�h�%�o*�!�eE`:;/�{Ww��CN�I#��V�J&^[b��M�TEC.��ր۷Q�R"��i����z�T��R�N^$ዋ���JO\a^�	�Pk�m&��r姰\�+�L���u��
�]yn��^�,���Wx�PȺ*:VQT{B���L���]\�aNc�g3ɱʳ��ev��M4,cr�^+ci|��)�0;@u-'4H�s�[ۦ�.1Z�ݎ$��D6@�Z�E���墛����쒋�v賬T/��������]`��J��>�-)1�.B����nR���1T��u�[x�#���p{�w�*9#����amC2(ka�AKn��ܡ�uI�w:�ib;T����rF�[�	�ֳ�L���H)�/��H6�I*p˱L0n������_���f�rm˃���ֽ4���J�qwK��������-jFr�x��qS)R2��zfO �_P�L��M$�::]h6��`���G�G�{�� `�3+gM��u /�4���1O���{�����c�!��m��ҋ�1LȷVf�ۓ�w"�G��<��[��i���7vs�k���U��X�W�ow:6���;Y�@��9�΀���B����)���X�2�KT��ۦjqp+GhM�����r�4����7K�����F�$_���nh�Gr��ۥJ(��)��i���[��s�vx��x0[���^v���k��r�S�?����%ZDuo�O]�mQM���coos��eޭ�*uq��[�H�Cuk@7��grn�,~C��Y�'�YD���L3����]�-�R�5�^��͛:늾�վ�ok��Eǳ۟d��������SEm�JOm�slE��TTc��gmV��p��R�y��#D����0LMv�Gz����S�(^U��eщ^X]S��U������9�*]nN5�Z���X%�[ ��V{4��U"�5��qVM�쨾Yjp]��,��c�JJg[���؎f����r�b��"�Ffs����T��TVMѶ��,͓9���v�t'C���r�D��S附V�B��wGU;T�����.�x-�e)XErz�k���+��q)�k=q��Ñ_vb ���q�����`�w�Ym��C�]�z��42�i�h�%�[f�[�Iv$�/�����떵okb�H����q����K���'U4x�[�2�bE�k̕��V&���HK�U|�h���S6�[�sM�q�قeK��M ��XK�m���+�0d�7�lc��:k��l����-oZ�HK<�WԲN��y��a��f�M29^��<��ֲ�_Ku�X��+�qrTy	ŵ���1�bC�B[}Sr�w�0������WV���<݃��][�]:����ض�J�y�������v�M\�/��f�ڟb��p��9a&,���Q���:h��,���v���<-�9b��>t�BՒ�J#�2��䙽2�w�����!��;k5b�ZX�Һp�q�C'9f�h�u-�݁*�{BT�:�}�Dq�o���)6��2�����	�v7��*^��F�ػO����J)��x�J@�g���^�7�#!::�AGY:��F���y9X"M���[v[�f����m�uz��@��oyp�-���k��Tk` /y�=s�j�ȤΫr��c_���[�܃E�.�C;����#
vw�=j�D�`o���t�
j8�3q���/���l�Y���YsN�F,�3�`�i��9�2�l�rֱN��x*,��q*ܡ��V����ĤhT�Zr.��,����df����.�K\n�O��D1�-UZ�}�Gss�
e+s`ӻ�+�v�p��j��ᔩ.���l�J�U��Kk��Hl�F��YE^$��?��ξ�s�W�C��"9�X�kp��c"���,�eĻt�.-C��z��R���0릑,�T�a�ⳬ�5��LW��wIV��:���rN�Sr ��iK�{���*�ưX����e3BN�m7Wˤ�ׯ{fQ0|��] �x(���Ѯ˘���w3FۈJ�0��%��C:������u�T�Z��e�B��w�@�7Rz�(_(x��הt�;X��+m�5��d�F�9*�/�ܜ���d�O�w_�Sz�U��F1Φ6��l'2&3��0������X�Z����H�S�}�#��˵|��W����Wvb��$���^�R-��X������L�u���խ^��-��=�����{w���z���g����������m�Y)��� :Ս���zK��Q4�hW*�c(����(�u��D>�ZOWpoi���*��9��bՄ�82�t��MTzh���*��:Y�5oq�#��:d�-��5�*�� sX��[Yy5GC�dv�M[��|�m�C&Э�R�]�J5���qj�s9�=�r�T%#�,VXKIP�I�֝S�>�A��%L<����	��8�P��Vp�Z��/5*� �I�y�w��'=�v��M5�rnaX,ڢT������i;��6kښ�튋޼e�)�*�r˭&�7�k�ڄl59W�֌ ���mp"	�f)�ʕ�}��R��2���V&4�M4�0e'/��n��z�o��ٰ+2�����������+��2�egYЇu�����7�Ƕ�▄�t@/b��݀�ydGbGN��$�/���fG4I���Z�[ۣ[�ejh�Vu��
�k�.�o��容n�evdTw9�;0�q
r���CM�P��w�Wu�ue�c6�ՍG�{%�*W\�(,c6���Y����o[K���m�g՛IkŻv�'uź �,������>W���,�5�4�.�,�]����n3%;w�l����D����&d͝�tҬ�N��kx�x{e�[s':5@��S���,j�hi��f�Œ�0�ŗ��^�\��S�0v��\#@S4�{:Ί
�F��n�&T�Q��]�I����P����"ȁ����NݪY���Z����q}9�E�5E�B��|�MMh�.�� ���̂|y��$��i{��iB],�oP�������}�q�&9ǰ�IQ�;��s6�f�[�)X�4긍%�bq���$�����)X9($�ՙ	�۳�%&~9���]�>���+UA�yZM�$)R=�a�cT�'qU�+%'�4�}rR��G ��MmY�{��ܡ�]&Daj�vE�͜�9׶����(�l;���F��=:0cXgSV��YE�Ď�ɯM��5̗M���l�y/Y�	z�l��1�Mq�"����W��δ��@g^��Y�TkM��̓�B�<1�zhp�z6��'�;%�7(��&a�P�����(m(�s�+B�k�%���ޡ�8�8��&�2>�����Dt</�ѽ�J�k2�:c6��J�� �V)!��/+��;� ��1�ӴH�����-��;uM`����En��{%*N�`�:t�r�����xl��K��Y�b�G�ސ���NW�rfe�;��Q�jť�Y%5���z1�F�|����_ 9�dt�P�����5u,�w�Rۅ=qؓ&Wj��;��m3��s.��[���Gch�����e�Uӫ���-�H�#yOsX�v�Ҕ��vNX"kr��X�w��F�*���;0�Y��]|R3u3��(�K�J�M�wsZ�B�堡���.�n>�v�*�g:m
�<}7�O��踈/nS��T�0}n�^޾�����āS9�q�z#tw1��O��{��	bW7�%{#%�[�T�s!\+):[y��N���}LZ����x��q6�d�;:G�Y#�f�[��_u�z�s��u��@Ԭʸ3dd���YrX�{�=�Z���LJ���3����U�v���'���Ɠ�V�����V����C�,����i��Qgmq��8�
�vm �R�'>h���,$z$�YW�L^G�z�o]ܢt��L�`seL���d�GZ�Q���>ڃ���.�`���õt�����\�JW��˃��q��K��Id}}hVJޫA�Y�o�KQze��J+�ı]��7�s�\.Vڗ�KH9+C�x�z_<�r6��v�Q�)���N
�qg,+��(R�_[����M��aV>�E�Lu�2t1#���a��*����%�(�c�:�c�e�����v��E�$�5	Yz�*!*����se`��e�tM��.ܒK���w%�A����̽%����ت�pPg���r��1ґuK�^j��5�Vwj��Eۮ��.u	�ٗj��
���s*ĕ̓�[���]�ԣ������Z�2�lx��q+�h69�"NX�<kj`��q�-0*�.ʬR��cu}�~�#��ΊAw�Gje�1�os�|Ѡ�X4�I�g��xw�#��[��Vv�<�����.P.�ʛx�Gi$;ԯ���N�EIX��W����>M��SZ��O�z�M�Q�j����\�7Q�3z��ZL9�p�t�b��DJ�lX���[�*%�ƫ��8�A�t�ݔ`�aՕ��ك�{msS�c|�G�_��c+n��S:ӵ��H�Qt��I��z���l	&e(�'Q�]%�)m��a������wa���\`�:��8
����[Wr`�7����.�v���5��zd���V��Q������۳R\/ �!�[%���n;R�C[u*mu���Q� �mퟝ_4�a|��� �Vm��*_�Sq�r]t<oF+(���K��n�e���+�-nIN�C��re�נl��� J�o\�@���°IM�_lՙ&;�vVL��_j�JV��n4��%Ԭ�39'�u$��*�0u��gRl����J�/�:��m��f��Jh	�P�]t:���
�:�e��C�{��X����ȑn�Q�Fb:��*�&ՙ4�))��*bdŬ.Ȃ�^Nior�f�}�f����CN����O���{݀S��ΰ�v�v_q��֘�g�wӦ�
�Bj]qb���m�j�\�ae+��Ou#OC�
�j�A:V�B��<���5y2B��~����z�{�6:��m*k��8:9HD�x
V��1�������"�j�S��q|�׬d��l�^'�[v҃2��8}����ݞ6<U1Kqt���s%e����K���6�M�e�j���b�\���@���A�uBk��㮁0nv}��<��x(��YawtӺk2�.���>�ʕ�B9լ)j�R��X���ǟ z���K�v��$�oH�R˄+�r�ź²aKm��x���:3�}@f;V�3�m�r �D�T��Y�g�}l���T� iaGU���:��3�t���¡�5z�g���hh�#�g5t�]���4��ϺsWr�G�9֍�f�vT3���8�2nH��W�X���
�vc����X��}���/8�g*���\�|h��̡@(�D��d>6��ӳN�"|и�׃qB+��Xo�S�h�(C �z�z"x�#t�9|�Ҹ��+����R�C.�c��<ݐ��m�	����*�8	�5���P:⬘��g�b�˶���=�
)��ۡ3_�'R4�JL��Ejuc�ڸ\�ڊ��+�{6L.#�6��K�2�*�	�]E*yk�l��Cn�R��MaJ��{�r��M�D]s�֤c�:0`c��
-�v��+a�y����kj�kS�.Ը��U�C�
�v4^�x�e��N&V�'S��p5W}�J�l��7~�j�M�}��k�f㥵��N�7\��S���,��s2��;7���ųUճM�i�6`��:\�c��^S�t8�-#�A�H�mK���6R�%Է4�n�d�l˻R)Y�}#w�����ݭ�3�,�{jfEJ��+��Vp��&`�C�\	j]����OnNA��䃏Ij�����s{���u�[(�]α�[�q�:��׺؃��r�_A��`��6���V�n�"A�J6�텚�\�l�[�]9�.��Zmt�:v<[��sU�dI.eK���	C�J<(P�{ɗ��W]�ϏJ�ԝ�M�t:e+��p�.ؘFQ+����g7�aG�:v�އ{���ig_l�H�7�]����͸ȰpI�j��ܙ��-��t�!T�V�ݒB#���,�9���P
� �9[Ĳ��eMέ�;�YW�N��ի��U�_l�EC�]nݴ�S�KV��������^������i�]��[O����3��6e��\iF�p�:g�2��棰7�$�b��������JR���,�Q�l;���@/M�!f�xJ��
V�]�v�۫�9h��)e,�x���EK�u]X!TR�7�7�/�7�D���ڛ�-NN"Vmv1-V5�W�c�}W�aak�]�S��r�`r��ƍ���n����a�h���K͇W+�b"�w�=�BS8�>�P�K#��Lf�v���k"���v���db�+GVY��89	kM�������c�;��c�Nt��Utm�{�6m���G"[������(#ά�k�O�vi��'ώ�(�0(4V>8�L�[[�WU�"�f,tju92�����k3�ҭߺlM^�tsM��4��]�"�=��]�.''��y�$ٮ�s9�E(Υ;]ڌU���j'ԋ|��\JW{@�x3-b�����
]�Dw>�hb��ar��
y��ju���4���xz��1Ӹ@�ؐMm���c���b��PM�O;�OJ��q[�X�
�ùj�^��[�C�ZLx� ��)^�ȣKjh�t�̣\��
��֣t����g�k[����5��͙A�+��`n�|��.�i�[���ێ���hp�Ȅ״i�*kOX�&�����H�$�Tu�)�*�u��c��u��+�@�q�6�H�`M����+��Dr�K��h���ZB��<ɰ�N@�/fX���qd��VVk'��y�����߿�5�����쭶�m�߮��ƕ�k�������t�>��/����Ε�Jo�G����e�kHG�巬\�%�kU�lF���AYJ��ǯY�w�E���	��,�M���kͦ�Qj��n+�[���o��:�Xռ�̅���ȳ��'B�.J@' ��#�s1�y����٬j4q�� ACXG�,�A��*rZ+��2�6ZZ�Z�T7��t���S�Cq����V.ܷ�ʛ�ғwE�����s��9N9B.�2�)�>��[�-�g%]n|)�Q��ӣWv`;(�Y��8���.�ob��8Η��1��s��{�7ML�jc���$��R�:;��X#H'���A1Qb�Czd\��3����Ӱϛ:飐�+�M��{'!�,WAf�G&��@M̩@��l�A=M���ĺ��]wA���)�G�jʹXn�MBtI�6�Vv]�܀l�m��2�����4srh��
r��r�M��*;o��o���/:,9y���	wz��S+	����	����i���Ip%�r�2�
N�;|w��;*���V0mM;E��e�܋��\��-e��52A+��]�-�]v��r�\��6��X�U`�)ʨ'�P�jT��[B�Q�M+��Rsz�~�ށ��ɼ�jl3B�8���oRR��^쁘^��U��J�&uu^�t�Vqx��uK��ɻ��_:�l=�9��KIRJ}n�zF�Iyy�����<�d�ؑf^Ժ�,�mX7���r\��ۻ�o��j�5�ڲe�xu�E<B��V��g�s��MYz�>#0����~�-�q;����=q,N	k���H����f�EDh����f`���	P��-��)l3�VꄁN���ڰ�D��ʋ8Z��5Jf��K���� �sX�RbI�L�J�c�Ʒ�ge��Vq;�.�ZJ���j�qZ S�m>��]_mE>Kc�7�����3�Å+����-���૽�.�Tٍ�����\���*Z�\��[�Z@�ڨ�o@	���������f��t���2<Z(mL��k%��qڵYld*�y�K&1$���\��,��r ̜�rk[`�b`GK�`�]��8�_t=>}���#'\h�n]e�)�e�Ro;�I�T2��m@���OH�U$"��/q��uiV񛧧;�5�G�6W[�*-e^��Z%]�I�� ���D�����CX���
Tt��)e��wR	�MY���{�@{�
��X�>�&=FSa�j�`��؅����;�H��2�J�8�ږ�us�~�P������6+��uҧK�	��Z�벥i�ދE�� ڇ�nΟ��egqԣ�]�u;��x�J���h�+X�Y"����i��{��};(�h�J7�
��hz^�F7OeK������oF��؝��t$��`q�]�R3����s�`�L�qxs B�o�v�=�a���QP6J��N) ;����*X���Z�l{j�*Ņ������k�!Q0���zh��>��B�G��5έp���h.���ihz+#Q)1� �ȓ��Fl����NNj�h֑CM�.��s��r��g^�� �9p2�հI�sigc8���`�nT����u$��pd����Z+3֋�+ t"�9���I�n�v�`�%lUgti�O�p.v}jګ�;��(*��6�q���b���r�=`�r�˹�I�iWU�e�`u���@�����U�2O����4[YI�G�����Z���jc�]��Hj�7,��£C�J�U�s��	��[��ג�c��M`���*�X�K�m���}}[����4NWYꆐ�g`�ء�8�cj|GmoWT�z�໅��kŅYj�ƪ���֤�|M��K�s�� ,�*=y�-P'�a��:��g��w(^Lݺ��Z�B���f���Y�e�$��U�*ri�+NJ=q�6GtN�8(�$����L�8]#FdE'Z�{[Ӹ�?cfp�8H{��u;���] �TYi�Bn�v�p�*z(�]�:m��co,�Qs�ܑ&<|���\��X#3�mK;{��S�4r�b��TQ�E�����Ymj)s�Oq!�e�ìI*�R�8�E֬��a�b�ہ�f��ܾ �-,7�݊%�����<z;-S�F��9�k�Y�Qji+��.��(�:o.�R�X��Lт��(tև�^�v�Y�,�����wS�*]+��'l0>ư�r�ZE	
�����1����5\�Ð�[�ee����fb	S�s uZ�9ˈ��u�I%d�BW7�{��6l��en��c+�ha�O���F��d�n�ĺ�}�����ݍir`]6�Mr���ĭ:}�i[cpE����h_#R_nQ註2�){�{�����'k���J��X���R�h�gu��NLʚH{��H��I�����n�`�u�z+;�t��Ŋ�i.�tVj�I�2d�\�-*)d]���0.��r�v�>yʱ:4i�8�a6	�r�:��B�^�c����
F�b�۹k�4��Cb"�����@ ��Y�;�fJ�W·e�z4�YPL�� �Ҕ�taN���ս��Q��+e�	ɭ�J�44��>J��%}2^eM�ū�4�-n��S�9���q�X�Ƒ�֠�m�yo 8Bp�W�_��(����N�l�A|�_sMu�����:l��y�;1���'z�l�<٥�GL�*���Q����:�鸉��S+���ųA�'�t!�jFz��X2�gG��&��J�\;lZz�iا�X7&���i���b�U�#L��Jfβ�&vm&�c�%]���Y�5��,�O8�BC��dk���I0,�Û�."�����j���u�,2/kZ>6�>K{��s��{�5��Y�Ep�EV ]&����<V��}��Mm�	SVR%��Y�gT)hVo��Z싱�l�ǒ��j�4�<�������Bл�G�*-�ajO��sθ��컾B��y�b&SdX�XHh����z��c&�2��˴�{ʓ�$�����r��J�鹂g�_��jٷq�gm�Ohe��Ԩb`�ͱ8�i���έ�������7�Sje<fk�h�����5vм�TȵX�ޫ����8E�F�x\��u9e��CX�:�^f�|ܭ�2�V�.L�3�Gu���=7Sg%�%R�j	:�7��0��#�θru���-\�@���GP@h�6+����a v��7%Wǝ7z\���`�A���t~�3lӧ�oܩQ���i${���&���Z0܌)�t��#'סa��Μ�eϤc,O�`�q��5��#�]+8�v�ኀb��[u��d����H��������^f%E�uu���*s;��SE�fR��%����-_"�qǻU���ژ���Ҧu_	Z�|�^ ]l��-�wt]���^#G����*�v�}�v�\ݗ�c�d�{�n�V�^�:u濛Z�,���ˀ�.�[4Aׂ:���1#���ĝ���(n����vu�┾�V���8��o���M>B�Y�����ќ�87�w��YT������R�żh@���{�L1I��Q6��mr� ��!`�=ӠU���ө�	C-h��x)w�]`JM:Y�*G*�NV��ǧ��V��Ɉ�ޚ�,1��7-�p����3AWż%km���h�ΰ\C�nvTU�͕���� )�{$4�j�o��{���aK��^3փ��3[u�n����@ꅓc!}2�$bU*T�~ܼ�)��V3gЄq������[N�r�4�0sE��@:�eR���:KMH�u��f���w&���:�.�}C����q7�U�G�t�#8�,�K���j�d��J|�X��� 4>�n�V)���H�'����sf�omD�M�TZKYx��R�M��}o\B��L�;e4Ə���|2*��!=�Įx�@ҝB��j_u�7.*�^U�k&J\yr�,΀����Z�t/�*Z�k�J����{5���7��<��N�|f�s]S)j�z��:���E�oP[n�@��nk��K�m�tF4@�}-�Xv��M
��f#6>��5���I��o`1�X�elyݮΩ8Z�V�����{+�{�;���HZ��J�9�ݩC7���k&���b}s�;������{mˬ���'�W�-$�f�{�]-)�N-Q݁n��|�k�HR�L��.�e5*B��r�C�w-wV٦޲�}r�^�Z��%��٩1���$S��n/��'d�?\�(���دh���U�3djV�.]:om�$�!EӮ
��EHK��h�(j��A���J�K��@k�H�[CT[��ޓ�#�R�ٕ۴��6���n�
1'�����X��B�����T� twv��b[�]� Dpj�n��
��h�褢��e:zxQ���S�s��3�C���Rh��t��.&,lC�{gM ���6�0k���e�2�v��3���Շ1
|�ۋ좵ܵrΊZ��v������;r���5S����@>S��,n]l�A���-��]hͭ}�K2<��hK���TGmv�5�b'�t����`Z�o�5r�+|��.�E[�WC�V��g��H����e^�ܥ��Qٺ�Q>}W�%*�@@���f�pN��x��U�0(&���ɱ�,��Uc�\�w
���@��*�����yJ���:l�j��siRS��v[�C5�*���둨4�7�Ш�v
�����T�Vh:|/�c.
l3bWjښ�{�Q�t��ޱ`	ծV�c��J`T�q;}3J��6l����6i
�T�2�X�QUJ�ҡ�[-�����*,2��r^�Y^%;L8�^�|ݪep͡[�4��o���c��0VhF�<�;��}\�{՘�:ŧhl�QYQ�js�������L�l������ڼ��)�)$DTi�7�B�!r����9�G�w:f�(�lp��y�����r:�s�YMօwd�:���虜�|��L�NKF�U"k:�eЛ	�gdǕi݌}���W�
��%���	�x�1rŽ�ۨa����e��h���Y�J�a]fU�8�^*��L�<[r�ܺ��K̴i>O'�s���o��H�]�^���Bk��N��ӫ{�]_����(����**�^!\",�N�Ie28:x�BP�R���2��7��;cg*;R��]*Аu��%o+�:���)��4u��MǮ�#��>�J��Q��x��΋���q�S�������5�� U���*���Wj���vv�ڻs��J7��v1R<�<!k����6��lb�
�m�������wJ�X�T���:��쿣9�̚�e�W�S��_4�>|��[��X�Q�&J��]9��X����b���X�p˺���,/�f�3�7�Y��ӡ��t����N3M�t ��b�q�J�xw����\�`\2�G�څ�jN��R�Y���{��.�|[S+E(�ʻ��ȥ�]�[��s�����n�d��Z"ʹ�!�;QS�s!��;��݅س8�P�e��m�\��q&��3/��1�i�4�Ԥ9]����W��	�L�]���YB�;-�Gy�z�R�f�F�8�)c`���?�p�2�I�����j����=4������xJ��cjR�c�|�Wn��ay:V��O���ÌRe�;�Үh�6�Z��V��+�v�Kpt��9R���lm9*Kf�J��w��]�P�G��)��@e�gC�n��+��D���}�4�֙��pCzBF��&U�
��e0��:����譵��x5l�o5^WgC�`@��+�����$��. Űr�Kb��=�'�5�zVRT1�ںW�wmc7��q�df")h�{o�m\����I�[b����^#;fӨ�@�Y�l�TB�g6��xU�z�L�9�Ij��W�ڶ���H���9�9��e�HұF̂!Z托�)�+V�W�/1�f�S3�����6��{%���.��oXX+);��/���H^�����p5
ٗ0ҭ��[���[W���U�<�������Mԛ�n��gA��H$N��k��$3�M�C(�R�<[wոC\j�Pk#8F]����r ̦�cԞ�	��n�КiM3���t�ud�b3���+�Θ�/���)re'6	U��jޖ���QkC��ܡ�W���b�ٶ�dj�k
V=ԩ����ޅ�b�LU��]�]�܍�ư�����|���{3��F��tx�Ѫ���uT#%���뭽&I1Ůء&كD���䦴$���V��_7Lɦ���l�z�E��&~ͦH�|wu��pY���h_��])��2mL �|]����L����˗F)�HPkV=�\2_��]D�4�WGS�*�c1{jQ5<���u�⏈˰���Vf�l�R��2��Ҭہ�7�ƚ���sD�6���bH�Bb�K�"a��oc�*Rk5v'9V>n���H��u��Z�.�����E�m���HJ�jR�%�^fj}j$���ڣeV.��r�XH�id�#��o��ѼG|���Z8M��]{sgd�\(��֩�{�95���M���Ѥ�u�އq���
O$�Ti�D �p�1��'����*&���]ɹ���L����k9�(l;ɸիL==ۏ�.���}S6T�(�x���Zʔ��K޵\�S����e�p���u��9[��u�|���n)7�>d��C�+���e j\���4T�k7�ˌ�tUܦV�O3t����*���Z��cc;������ݕp�vr�n�Yx䠻�܁���ﾪ�����������oo��L�̎���Vj�41��u���;aatvjt�Nq�X�(6h<���B�9l:��T�6���Gk�����U�J�+�����.���G�.�Vy�]��&A�zXG:�E��V��v-�;�}�I�&���j�co���Mv^=�%x�s'bAR�6�c�il��Q�/1�v��?<ǪUޤ�����n3Dz�T��m�����V�v}1���+�<�,��գ�p�a#�!e���1M�v0ܻQ��Ֆ���=�����=m��-�:S�^�����;��b�d��ZC��:𪩌B>���mm��zr����2���2N#/���(�%�͸w��a�S_���a�~��n��hv�ۡ��r�2V�s��e �
�'.Nq����U�/���qBpY�u�	c^�����ǜ���V%m>a.RQ*Q����殶2bZ6�q��m�d�� U@7"s�0{"�s�"�� -܅�N�,�HAՆ��^�&����e��%nd|p��t+�!��P�:�me]��F&�֬�J���υ�!+`�Ay_2���]��ór�۲�t#��
Ca�Βs�	sm��={���cs;60������Z�ՄD����������Ŏ�.�+�9��Hz`��y����w�jwAw�V!=zK�����3K��b5����yԢ�\��3��#|�{�ߟ�����������ޔ�L���6E4j2F4QPh�3!6��#F���Z�&�MA���D���D�fZ ��Ib�c	�[�HP
)0�D24F(�4RM1����Ihؒ-�$j-%�	��F-�р�&�f���+DT1��	F���"I��@M�5�HT	���Z5��3(�h��"�C)cF�V@�H�HأX
��(�$X�(�Ѣ�EJfdر������!G� �W�}@}B����NN��,8�I����7�ԝ�#��u�=��t``Uv��n9%�],�͝u��W�=����I��:<��i�!e_��,��F�_�{�#\%�q֊4������n�{ץ�B�e]L��}&�]��#�OG�ǀN����cZ��7���Oq�.;b�)w��z�mcݭ�s�roy�`��V�6Շ�,�5 Tmp�1}��o�]	ӝV�v�p8:�>
��gYiۿ�0���4�h�Y�t{.��4�ea�j#\=b\n+�Z�3
�)%���P�@��\n5��C�wFK�G�����
�[��W{�Ο��^]��&�;����n�**��EOP_�a�1|�1����x�x.0����]��3SC�r��v�t����:�T"r��i��w'0M�kD�Y׎Lk�}t��yڑ�;2��^J�b�Kݭ!�V���Q�2WO�ȇ�}�p�V�P����aj���t��-د�bi�$b�����Ţ0p���'q.�v4�ׅ�K�u�^f(�y\^>�s$��:��V��C/����{Q�}�*�#���'�T"�*m`!��Xj�U׷0��={u�SGA-��^�EbM��l��2M���b��ÈZ�U�3��3ne�6M�Ӂ��@0rð��cM���)��	Ì��o-��ZC�&ґx�$���;���;�a�,Wm�fO���φ���ٷ�[Sk�[}1���d�/�%��ƍ�w��=��Ǡ�x`厗�9z�X�+�0�(� �B���N+ek��.��z��82 ٍ�EFL�S����:��>���p졸�wo]��,����`�!�.��T�ΞDA/�`F�8H���d���#Q�UA7�V�|[�L[1aSt��ho�g�!׋���3n&�c��>���F�d�4'Wqڱ�^q>��Eג�rV�6�t#���N�N^��k�/�`��S����;Ř�G��v�9��}Ҹ�{�.�mH�����:��Ϛn�E,�dѸm���j�G�L�ʁa�v;�~�����l���!^�[�A��r�*V-ØZk�W�!'v�c��3�盬�Z^f���Gj:1�N)C=W�{=���J��Co������١���O�3�΂0�]|6��
�fǎ�4}������4�����c�W�*c��,`9�HѸ��e�Fs�뙎fE���:��/��)E蝎j�_�뫕^Ť�AF�t���2vю��O{�U�q+V[�=���_��<2:|�(jA0b_Q<q�}J=1��i���hw&Z�١km����������S�*ED�Pv�G��_�zv�����}ekB$u�|E��(Z�S��.h�n�p/u�8�h��'�i�T[�r�G�\�زN�r+�!��2�V׾�s��v�/"�i��`�K���[����W������}3J�Ny�w�Vte%���1�_͸u&�U����D�D��T����U1��L��\=��y��r�"L6�|�K��!��^�=b[�e+
Ӑ����2�م{;)ʺ	�2�;`&��k2�F$�폯�p�ϋmT=�g��1Pdc~�*���>�j�A#Ğ~+"����Hn��!:��aE.�0\s�hƲ,�C��p�j���ӛ�/���
��p.K5��&a����ZM�9���}£뉹n�U/�;s�ođ+/g����8�}"�5�o��O,�?1�|R�A\^/���5�.5�Ԡ�]��Նwsi�=w�s7�.pG"�̓�۾�r!L���ƥ#d���=+��tk�^�m�S��-Wf��ѝ�[,��O�ѸNc�1p�m�����&'��(�5ף&�ڬ8�,�ɾ�g�Q�C�,;�/�V�Nd5xT���'f��1������9����F�C-�Wq�C��w\��s�b彶�Gyu�Ǧ�T*�Ӧ����lH��g��p�;��:Zsh�e�*�P��17���-[/���lS����[5	��[��UܰejX��':�7C`�J������L-�[��N���s�`�:���FKn�'��Xz(�z��7�!��_pP���h��Cr�&����ugM�����յ�%�Q�������!�*��/]�n����K�u���_�]k����}edm۝[��$K�0�]�)��8���Uҩ��Me��W<�	}lk9E�"�����\g���%��ۧ:P5�<��H�.b=d~8;7��?�ޔ��R*�3���SHd�$��?�M&Y;F5mWۮf��o������Pgy���z���]6��׋aߨ���Y���H���)��l����F/M���1�aj2|�ܺGwg%��o�̳s�1�.*e����ϴ���K������N[=���9��E���Ȱ���2�;�4ii~D@h�����^��MD���]�b;!��F�0���@-��|#c��J�JY�_��֏��ó�i�D���
�2�v�g���>"C�љ^��	Vq8y�9I�j{��]Wlho%�PD���X�^��]Ǯ#���	���br�t�'i��q�V��C�9�����8�V7�Q4�n.�F��"&�`+��9�%��0א�p?/tk2Gj�n�v����>�-譒��g�Jb�6��H���Q��+A��iD���WwV�ɕ�;2^�Ǽ�-��6̳�����:R/c���U�<�\�	����9�rmE�de�^O��AJ"�y��w?��SitݠS]9g�hƳ�����m��oJE�!�18�Q���F�O��=S�8r��7n��ք����B��un}�>?f��a�ڲ�-���J���72Խ�e���qr{$��L�WV#B��W+�V���kW!�����橒�,o��N6��=OdJAu C��`/i�rD��z�Ֆsӈ1�y�EDjyl6���0�������qT���a�0�-1���_E�e�NP��y�\Y�
����k}Q�Z�7����v딄����U���~~��Xz]�k�h��B_�]�:5�L��s�y]��6M��)L�ӯ��3L4���۴&��r��#P�W�K������B��z���l@��CGY��GƄ�d��S��k!�uN��s��Cua>~�m-�6�k�|����V����>N���P/�H`t�<7�^`x^�/�&dtB���q���J��/R����e�e7�WZK3Qᚪm�v��Pї�[i>�ڷY�fl�PP �ɯ>R�"�6����E*g]Lto��"�e�-�O)�36�vH�p��o�]���w����y41�vJXzh�V��^0�EW�����aN��$"��"�3��R�s��ٺ׋Op?1>'E*,O� %�j��R$U��S�[���A8U�<|]\�B)ĺC���;n��kr 8��y�u*�!4ݻ�[sK Sb�vSZ�r�{�Z?0�Cd��ڹ��h���p���{#�<a�y�*�������*ܞmOu`Ph�١4���9�e����O:� )� �<k�  '%䖆��6��ێU�L���ٛg����E����i�r4���W�aU�(��@�ȗ'�U7רqSO� c�"�fRS��������m_�졭��<��(H�s)��xd�J�V��Oެ4<WЊ(�5)�3t�=�_M�4Trj���"bUO,��Jqd�9��$�o1\C�t�Adh�w�_dG�c���ֽV��n�y�6z��i���l�	� [�9�%U$S����#�D?]Q�x�S�YŹ1M�u3=}*ێz;	�/����5Q"�Y<ɢې5�2q�$�l�;5'�Pb�
��t�9)��n�ʰ� ��ոi�u;Hu�[�ٷxzIF�P��5�p��=p�U�ge64�yO�qQ;����:U���.qO�k���X��[�[N0��&��"�oso1	ʹk�G���J.Y#��+=s����FSjTw�̗���Ɩ���e=5���bN�ϟO�M}nT��Q�/J�u8M����
\����T���ݣPO�`U��	��|<�Ѓ������s��-s��{x,UT�<��P�M�k{*v�#%.,3��P+�"쎰%�ICˏ�� +q�1p����s��4A\&o�CX��N�^X��l��G��m
��\Ne:̂�}>T��'�;�F: �J�}n�1%T%u�=j�	�/^b�>���lVDl�N�ג�3⑧�����W��!�:Z�#͡j��C6�'�ɯ����w�e��u/MI�H�`@�П�1��)�*���nMdH�)����<�������eY�岥��8���D����U��Du�8��.r[ �:+CJ=�&c�n)LP:�1�k�HfA`#�ڸ}�g��s)(�Yt7;�����a�Je@=	�*��N�K�޸��x`���^�R��!ΐ���R'Y/w��nP�2er�R:G�`����5���}�N���W�:Ѵ�u����=��&�k���\��Ho�+��NM �&�E[�b���o�V+�
U�̲��>���3A�������k|�L��i;WD��S�k�]�Xy+l��F���R����iR�Ck[����_S�>�p����sV�,ޤ�w������s�H�e#٧}�y�	��7�pY�H�1�(q�t���]�03M��Hh+)�$�j2L��M�g ���\���F�p
�'�׌��@�<"QV6�����ި����a8
S7�����}n����b���%�5�T)�H�F�Ls����F7�F�:�J�nc����+M�ju!ךؔD�|�ɡ���ȱ#��I{aYK����:�ݲk/@�#�`�+�,d⧦�f�U_!����q��e�M�m4N𫉡����6��������Ct���??��a��!�}�lh���7�ULFN�*J���\�Y7�_�4������j��ՊP�1P,o�̺�Q{�Wu@��}�2Mr�}%Fk�Q�����w�����/I��u��j���{�.�|X6c ;3T\�D������Rtn��ޏ���Qp�b-�P�T�e��F5mW���]
L�
��a�K���=���'-{�8��8.���`+�5Es��>�t��<#3[�F/�6����1l�o��i����h��Q�\��o��=�Fu-��.O���e�����bӘ�hJ���Ͳ@��V��.�d�t�Lk��.F���%�8�q�5Oo��_No*�y";�f�^��Z�,:ȕ�z�8;^�����MBk�H)��(�7��Ռ��I�.B<����4��
�������~pzl��XV�Z�'��g�{�Æ�}�B�[����iHn�g����v#�!��F}�&�*��'�ľ]^d�[�j"偮��kʖFע��>�Ğ�W���t�)�=��	�����!��"�����ך&�l�����21*��D�t�I
a��0�@v0׹k6�^�$~ɏ��td��{%��eL1�r�#j-�#/�4��)�EJ�́�&���HJ{��^�T$�h=�p�o�WȔ��7�#�9����ۇT̊�2Q;��su���>�pR�q��@����D/���b��Ln#,;/��ϩ�Ֆr h���:�
xT�n���X�p�BcJ�x	o�{W�t95r��_�ԃ�j�1pT�_sT�wKv���떖F�������9�E`c�)}��C��c�J2��++֎�-�tiOv��XC���*��w9ܱX;�F hq�KB�ó�Z�;0}�g�ڨڗ9��i|Y40���ӣ�be�k�-��eL��I�xb:�F��\�H�w\ty%��7»ݙJ)���Z�w�7ҙ���̳�Y\23Cl��)圢����R�d���.��+�N���d��G���&�4ܲ-�Q�݄��ղ�Ra�oZ��X�\���#aT�͊��m�'w�s�����ꄬ=.�5´]|5З�z:���N`���t�^q]O���[.;m�֦a醜N��9��W����l�iD�\�'{8�w���|}<U!ޡ��G�����gS�q��˨b��Q��l��jO�TH]�^0�d�Yk�h	��Э��|��Z�@x8k�����F+N��l�l��f	��թ׽Sk���x\oeO�,����!i�5���JC�;���+�=$�\x^?N�d��~~-y������C.�p�:�^�C�#���;pF
�x�`d���n���Nt����k�wƮ���n,z%�6M(xu��*��we�'�����ڜ�OlVߦ�C��5��<�e�z~Ci�\!h���� ba��xFdu�-W)��8+L��H�-��r)�����]�y��Td��T|�����s�ktf�ҧ��������2ZH���u��p�ڿ���7��G�P�7�C�g6x^�+�Y�����Yq�ԩ�6LX�r���O�Y5�*[��]���ܙ ֚q��Zc%)wIu7��+C�����rXW؄U�U�4�t�ot��LC&2��`�\!du3v�'^uqʴ����ϛŋ��+��Eu,ۆ�d�a�sv�/����6{C���R����P��=[S/��dGV��Jqj�T���C�/�����듸G�W7�u"j-ܣ�S�ۏ~���(0��*ak{_����v�خ�v��b�f�c�5�RrM���t[�LT���g�X�%:�N��k��_1N;�P�DE���k���P�r:6KnT�/�6����[�e���
��)�n���cpHơC�:�\��d�������@.��ћx0f���R�9�8�$Y��G0�)³��\�^���b��E
���Cxt,��C�
��[���,������h'n���"�]�
I.���]�G;m������!������S�٥Њ�A$E5�XyW�uf�Z[�ү������s�O�a]@w0��7(��)l#�7(�T6�pŚ�`�y@��U�JqQ^��LA]�
�3�j�-�=7�r�]�|��ʗ�j���PW�,��/�kmu3��-�����kn��4�,����$�&�)��^�\�=�3��%�F�@iD`�|󍫝6`NVt��/��W`4��Z��צ�/Rp�����ϱ%��������K�tu[aҡ��ù�!�7ELZ:�Ӽ�Y�tE7:)�cvK�2��W2���U�uuټ�km����AIV�ڽ��N�-\*j��yo%>�Z&���A2D�E�1�ɺP:.��yS���&WÞ(�dH�@ڮ���ʶz�oO���V��δ�-���ٛ\�"�h0�V��:������|�P32���G^����E�;�w�W>�������P�|�]H07�U��x�he[�OK�|7�G(�q�K��읥h���V0ӡ�W��$u+30��I����nD;������A���l� �A�%;0RW7��Jk+af��l�ޮq"��S��\z�c���|�a�w�%���*��wJ��'2���k�P�&ɖ��"�T#TY.���]�����9�6���S�]��ʍ��\�2�W*Q�r���R=ac� ������V�����P�Qj��青��x9gT����w6����18���<�,Q�U}#F����L�˽z�a������輩 ���qtX:�]�J��9�>���7i$1P��=Y[o���oegA���%��H�t�Ɗ)L���l?6}�C�e��p�7g
+�%p������(�)(�vz.]�t�(�@�&�k�%���/�L�HX���������и�RH]���ǩ���A3��ێ��Ԩ�p�w�HH㰡��eK��K�te�"W�����_�������ߖ��M�"1hj1b
f�1�1�,͂��E��э�IL�d�Dh4�HD!32�6fLh�I$�0`Ę��5	
,F ��!L�f%3F�b�C�!�c`6LA$�P%�54�"���H�B��b4a$MK0D�4!H�6RƂ`RXf��XL@��0C%%��LI�4� �F�� ��HSSBQ�Sl�eA21�Аm�1A�c3�0�l� lbLW����~9���n0���cgX`�M�b��rE�N��]O9�nM����K効5��P�$)W��m�{m����c�������?�zZ7�����z+Š�^�^"�{W�z���v�������?ͼ^-/{o^�ߊ�_��-�^�w޷���y_�O�6���?}�ܫ��!?O�1c�>������k�s&.]�?<y��W�����o�<��W?ͼ^{��կM�ۻ���W���Z7��y�y���������ϝ^?<���םk�ϝ������[����zo��^/j�}����� >����fF+U�����>�Q���^+���������c����ߟ>��~7���o�}��ž���w���|�ʋ+�7��_�ϝoJ�+�x��Ǎ;xۖ�������~���1U��,�Rhg���j~�A��p?P|W�x��~/~}�W���m�~׿�}o�V�_�~��_�zW5~_?����^/��~�|���k���������W6������^-�z���i�m�^�?�}""��{����#�s��<g+�"q��{�y����6�=7�ݷ�x5>ׯ�V������߽��޼���<k��~����h���|���k��^-��^�"��J�~��|������|����������}�${ �����Yzr�Ŀ�����{�}�й�u}���zZ~���x7�nU�������6������������_���y�K|W>���޿=]�ֹ����??6�������{��o��|x��>���X�#��2��_5Q�q�ly�������[wεϿ�/�������u�okƼ_��w�W���Z�wx�k�^->u�_�zX��ͼW�y��s6�;+��ߛ�o���������Qo�!����1�>�s�g�˰�{�����y��>�үO�ƍ��{��ߍ�o��^o��Z����o��ߋ�~+��������7�x�+����痥�|W�x���+��o��_����o�^��_:�PPt"L <5��O}A^M��ϟ����-�_m���z>v��x��b�����^��>z�~*��_���k�ߍ�5���?�oM���德��+�{Ư�߯�zo��Z7��ߝ}V>�H}T�͓�H�m�H���߳b������lEz_���^j���77�w�-��o������7Ͻ��z����~-����_�x������_�{mͽo��/K�����ۿo�-�^�6�x/^v�
��Q�Q���ޕпu+i�(����5�rr<���#���:��vwU�dy�4��:I��Su��˭I5AM�V��}[����Ϩ�qw,�c�<��\-�c�9�D���R�j�A�5�ز��C��wb�p�:9��rzƎ�ÏC$g�PTQ.���J�.�����QH{�|c�#�G��z�ץ�����ߝ������}����o������n�~�>����^/�/�>���}_Z�|^���_�E71���j���urǋ�oV�}�������8�m��i=j�Ǉ��}��#��E�6-��^�˛��6��߿���=���ߕzkr�{��o�����/�{[��k�Z+�o����/m���������=�n�K��!�X��D�� �b�o�r�����+��⹼U�s\���y{{m��+�����^��{^5�{������o��������^�y���s~���{���W����x�|������~߿�T�.j��Dp�������0����G߯w���������_��^>+Ŋ*"��m��zZ|����>-��6�x��<�������[��_<�~-��5����xD�I}�q�(��ػ�i�}�����������ۚ�����_��oo�����/Ž���x�����s�����ε��7ί^�o�_���w[��=]��ܴW�ξ|��o�n��t�E��>��pY��r+՚�Ĕ{�=��~�����Ѽ^��}����W��^�}�ޟ��|�}�z��叫�o?���W��o���_�~���������^~��[���u�zm�ϝoj�����_>"� ���">�d[�N��'o�di�;�]�Ҧ����p��#�NhG��H������皽7�}o���ߪ�x�o�{�����[�^5{�>��oj徫���^U����^/W��<����~o��/���-��疼so���}/�������>x�������{���^����_{��~7�nU������۟���+�}���o������7����|�^��7վk�~�����Z=���_W�^?��Ͼ[Ң"8G�}g��?|9��tG��uY�_�����w����x�����{�o�;o=��7w�-��˻y��������m��m��z��_�����W��ך-�\�6���?}_�E�+��ϟ}m��:�G��{ğy����}�^dW�ߐ7��7���y���x��wu�<_o��=7�nZ?=���u~7���W��ޛ������Ѿ/m�ח�_�x�_���ս?��W�~׿�5��W,}^����_W7��/�2�������R_�Ω����Ε$�n��C�B�m�+�Vs��
Z���5&�7�f�I�V�yf�
�H��&b�&ħ�5�������%�m�J殹G�e�
��=xuqTQH��d�KH. �!�-j:75I`��݇�N�K�}����}[�/-�'���ߟ�������U���ǟ�ok���˛��*��x��}�4o�ܯ�������~_�^-�x�W�_��~��oj��/�ο��/ţ|~�v�o����oغ���h�">�k}�+y?q�tخ���ׯ�����[�^/�Ͽ����U�s_��׭x��ͼ[����<���������~+����_����ܷ����m�s~�������v����y��߯����1��{p�88�A��k�����_��^5}�=y龵�^5�ڼ_�:��W������_�O�����^��|}[���/?ߝ��v�{����+�V���}��_�x���~u�����w���W�LR}��_O�z�z��v�����ߞ}��o�s�_n���5�ߞ���o���Z������o���J��޼���ۻ�������7��*����K|���}m�u����U��Wּ^�ם��Z7��_~��+EW
�+�����=��O��=ݜ;���[�5�W�l�����}��zU�s~�]�o�o��_�zm��sQ�޻|W�;<����W��mʽ��4nm��}���5��Ͼ[�>����ؽ�#�������mfJ�{�\ߊ�_o;ҿ��x�_�;ڿ��7�x��~���r���b��[��{m�W���~u�K��o�����Z�o�^���V�W-=���>���0}����R�]*$����V�lS� ���s|o�ϾW�ܮ�����Qo��x�޻_����\�߽��zk���m�﷍��x�ߚ�-�^]���^->v�??�^��>-��o����W�>�>����FV�����"�k2�-S������Š���6���������o�k��^�r������ͽ-�\�o�:���[����o��W��76���K�\�wu~�_��|@��to[6X�xc���X��v}�����[}������7�}k���>}�o��hޗ�}�\��ڼU�y����V綿���|��׮�����~����7�~�z�~v��Ž/��^��n���DH�>�	F#�k:y��q�3sћ]�˄���-���zhѹo���z[���k�\?�y�E����_���V��ֹ���z����W�}^-?�;����x��_�}yW���s_�~��_�O]o����b��>��U!F���|?$]Ӧ7�Y� t�#���	�v僆*2p�a�(�NT�30�0S���QX=�3=N�&f:��O��	f�xf2��M��9��,����J�i�]�s�b�f7��C@�i�&H�oa��
�#E�O'<Id�4Nw����3NI�2ￕ_W�w�F�mW?��B"��H��i��E���~w_��oʽz�ϝ��s��ߛ|_�o���o�yoK}W}��7�Qo��{�����U�:�/���V��kǾ���
^=q��(�P╃/�덺��{���z}ޖ�bz����i���������W�v��-�����z���W�G����}�zW��~~����{m�ߍ�_�~W⯋����<�oM�o���_}b(�@�F��h�~Q^�X[��<�+��������ݼo�n��������Z7�n�|���cxۅ{k���W��Q�ε��5��y��o���o��痶��_�xׯ�k����������1G�m��cՈ`���O���b��_�z��{�����Ϫ=��s��w��_�>��o��Ϳ�>���~��~6��u}<hѹ^�}�-�x�kڿ.����x�7�-���s�#,Ǉ�"8Dp�}�p<�1�u��GO����߿�[�[��o�y���V�������o�~-=��k�Ͼ��~���W��}_�s\��x��ץr��������V�W-�����ͽ/M��
�.�{|Dc�G�D17�����6���<��[�5���u����]�ֿo����oo���~U�5�x���ﯪ�Z �!�T��?E/ު��#j3J�6y�o�+U*������)ۮ86M��>�'/:���Ce�1
%Σ��ڙr��6�XY�ĸ�c��UW���#u�
��
���J����b�ZfB����S�3f��'�!���Έo�0��ڑ{�|q��Ou W��:K��'�Gv�31��[cs,��f}o[Q��a`Z�ǈ̂���	������C.�q'K���?��7��M�	�%G��w�s�g��.�����7���8�W�
�w*��(�W�cI,d���(Y�����6�����ҭ�ӻ�pɒvN���W��ܶejs,u��sA���k�����:R!.�Pؙ|��(9�}�˺V�R���>��"!���nuV�O�wp����#O�,�w������X�J����'Z\�p��8U��;��*�ڌ�t�\�F�F�֥o�2z^�����\ "����^ᤴ��Ʈn���*c�A��H�l͍��ֶ��n�5���r�i�r4��g�::d1[�.��q�HU���[u�0����S�����N�pȖ��p졦`�6�'�1lp�h#�����)i/׻Ai�L�q�i��	�^S�.�t�6����i&_�ؼ��vh9����Ɇ"�'b!�Z�Q�P�l} ����T^H�st����k��^*��hh����٨�N�ɤ�p/� ЄX
eI�(��5��ә�K�/ƷP�2�nϨ�r
��J�G'��jdt,�dѸM���5d�q��J��o�ۮ�eˇ���;�[��4q��tG׭eD
��S�Gv�>?94�@8��+����ئ�v�]J'Wr��&QB �.a�����<63�V���١���O�1s��+�"Z�esZ}i�T��N19Tf����S9.�P��j��}��I��9Z����3)>��0r��]���;2J}CTVX\���e���u)�Y]�L��,�#�u�V+n'v%��!Ho6]�÷{�F��qcഩ4<ڟ������ʵ����,O����dJ�ad�P{��:����'�����@�s^��y1����<��Հ֜�/��񧾴&���O&��{�⍌�����@�z����GSO��$ �2/�T�lϹ�ߤ��m?"�y��G�|LivV��l��/`V��ӟ,Zv�u ��<#��Y3�s/r�yƺ>�SyV�yn��Y&��]������pz��l�]c�T�-������u�������T�_gD�5��^�>p�Cz���v�"����PB��=�fT�qJb��N������,v�s|j���@UI�%�.f�*ߊ�}>0�id��� F�1X��4=��%�w�GJ�0|	ƣ'C�}�w��R*C^�:�˕s�>�m�� %:NA1̬�k�$m�W����ތ�Ǖ��n.W�=�.[�b�.��݆�Nx����'U�N� q�T<>?U��ǎ�[Rb؆�vA��e���Dk5��}\�$C6!���Vۭ�ࢪ�"z���\ZV�4s����:M�`y�/5��r�}��P"םw�\��
�ob[��|^A2lI{fT$��hT�&�<�eg�rs�i	�{��>2���^��/�E���_6v�e;bF�B�n�8u4\����2�N}�f�i�+f�
9�<�4��Х.�q%^��ﾈ�����[�
ӂ+��H�ݏ�Jf�4�1�ϭѿ����Ù�KȄk@�Sh�p#R0���&�-�����逸^�B<��P!W�0����oS���
��;4m9��1=�V�s�֮�;�N������1}��Mj�3]{�t>Cz�T��?K_I��}z�~��k�u}�<�{꜠�6>��4���c���_�n����7U-p���lh_&/6��E����C*�N��:��!�_�
����mX�8�>�ls6wj�YM�����xҹ�v��A�)�n#vձ�&K�o����]A�]U�臇�f�<́���μ��q�1���%����YU�[�\<U5̲w�1������[��EY����h��w\�x(S�mi�(��n)���I�82��}9�(zj��r�`���g�A[�0'��x4O��2�����5�6��W�H��n�Zx_�/
Ԥ"�9��4��
�P�4�V��Tv�z�wbk�ۊt����q��2�ـ5������g�ԗb�Zk�����#ԛю��:�ˊ�\Sh�زl죒VT���w�D�5�r,��	�]����R�d���Q͎�;��yQ,��M�J�(뛶����ŗ4Vv�i��k:��{]O�(u�D��%��������/d�6��v�I�eAwc��"���?}��_}�S��O�A�Z=��x���w��h��%�� B3��*��&�շ��Q��e3)Q䔞씢l�-�r��9��{�#mU|�I=} �RP m���~W��r���]uꂣߢ;i�MTJ��c��a���	���{iD�#a�+ʛ7����{�8"��"e*�Ti����o]<4�Idޔ�9��ۘ�������H���5%��=����=�\���5��
r��|~�����E��̉:h�u�m��t��a;��J���p�#�A*��
a���"Ꝯ����ݾ�C�J?;���L�oF�;���+v~i�"^3,rX�A�� �Zo��qHu��F����F�6my{7R�D{�|�_MUѱ���e���9V���4�����Ulm�q�R�u��c_���6�c	ǪL�g��i�>�zgo�E�B��}[��xz]�\+G��C��防�N���Lw�j�Z��.�>`0؞�?0*p�?z�����h=�U0�=�]#k�%,�Ӥ��=�u�����fl;�}z+�O/G0�S�2=�R�bQ��(N����/1k)vf�����wq�7�f��^���TxCW�Z���Qh:
��z�ܸ�wN�#r�<��ޛ�Ӳ�e�*ݸ�e�ɛ�/u�[֣����}��W�G�i��='�tA��^<M`�(b��k��,���@WѸ�C�wAg�I�XB�2�3�q�:Ɗї����x�ƀ�|n�]
��	;P�W�P�|�3"	-�#7-������AI|=L������w���6�x	6�}�?�U�bx�)*P��.V^�:�5��1`���"��%=���\����*.�K�8d#�����'�9�Αuۺ����8*P<}U7������p|»u	r�1�9Z:�&'���s.5G�j��~�<��+"���.5��Z��@HК�J���!��4���θB�	�RW�[�b���ε�ΐx�� !$��#9e#����s�n�4[<0\G-v��r4�b p7Rr)91�=lK�9����¥"a� n��8Wi"�R�S���熎���a7=�B����>��Ně��;����x�	g� #|D��1sκ��Lp{��F!���x����tﻝ�FL!�ݱ��Dų4ۭ�㸚0Y���A�"em:1�\�;eZ�k�b=�WX���wV�ͭSu1��\2�m��t�^���n䩴��G9
��
��U�w5� rkQ�������FJ[	S�՛�@2�5��g<��uf��yeq*ݫ�史]ֱ����R]̃�&���XΞ��Պ{�wh�}�G�������4�p^f�CW�Ѩ�J�ɨM��`FEq�L�*|5q>Pc����*�S�N���\�%dz�g���x"�����U"�O2h�ɺ�C5B��Y&y�q��:����-=j��b�C_+�~Us��9Yu�Ug8�}��������չP���[b1hsQ���!(��%N��Շ��7ƀ�Z��AVtk�:٘���Y/ڰ�_�~p��0��l��Tm ��BY��F/�~��
�f΄L��t��Һ�Os_ �1Dd�e�����6� �fY�e��b?a�C����ӗ�O 	m���=Ʋ�1� �xה[�T>�ѳ��XL��C [j���H��O��))��k��Z�:g����]���,wa��"2�v���oT[��F�b7�.�O3̭�_!��1�n������:�r��CI�1�w�p��$ר��%�[JEQ�	1i�ܴ�`�`2��r�R�}�`٩J��qì{����V���H(B3�����=Jb���폮5ä'���B�9^�
�|{�n�DD!����7P��؝B�*�IY
1.�.[n8�*���6v
�S��j��>C�ڌ�%��ɞ������Sc[��Nv�L��J�c�]�����B��@������v���tg=�wNT���mL���HT.�f�b���k:n��[|�MvU#�&l92�d���&�VNg���(���
ܓ(� ��+l�
��Ӈʚ/g� V�=����7�:���<��H�wDguL]��!��� ���� R��h�q�����]�1�Ԁn'�u��Tm�L�h�o ��kZz�w��z4�;��q�~+m-�9��F�f��"Q��s.�۬:�Q�K���0�K�-�	�r�T�@���Fkq"�f��;y�у��*�t�`Cv���Ts7{�V-ִ�Y�%G���aםn�i}��+�;9�`hp��d�gt��L8�pI�mL�{���ڳIXM�S2d��4��-ϖ��
���n���Ct�;(+I�g,Y�HzC���F���򚷰�j�1���l�+�qN��W�D$ř/%I�/n�!��.�U��I��b�Ϸ㮭ME�����X�L�(�ȹJ�d9�ܖ�+�'lJ��8BefMA��MK��dÛB;�|��[{J��ˬ�6���nr�[��8�r�6Rb2������[1�ϭ�y�*fA#��0��Tcq2hv���I7��bx;R((#l��r�P*�%XN,�Q�������d��aC��G�Ud�]V6�`T�7��qS��ͮyk��ʐ丘yzH\pSz��Y�P�Y���R�i�(�����w|������6��eJ�t8��P:^��F�}%vcWb�GW��u���-)�ʎl���ɉ��ofѬ+y�\�;�2�S�F��m	�j�ҬS�0�8<�v��yjQSV��5�ݔ:�Tt_�!�S��4RY."�?��;H�*�V���]_ngdqAZഁA�T�%�fM0[�B�*��g[�y,Ho�	�@@�ܼ=e��:j0�;�5or!$",V��K�p��v�^%*W�ܦ�!�f�Εi������۽\�5�E�v�N��}V6�{)Q4҂&��,�:Zu<5��$N9��Bݎ[̴v^S�G)S�WB-{��Io`�[#�|��ɕn��qMǅb`>�=����UiY�V�XUb��o�q�]77��Vic�zqR��f�)Mo ���,�2���yw��.&Y ��odW���t3��GL�P�1eթ��3f����v���9ڝ�ͭ�2��4)b�aI@G"Sd��͑*��(cw/�4��	��.�=�p��<�'��ŪSim�-���@�[��Z�r7��;��$\�t���z�����6�^�_a6�:�.��;�[���I���+�Ж�*G�L�@�3;�ۆ[�R<��8�N�	#w�c�<i'C3"�M$���d�ys.�U8�e��_]��%bi�1�#�P(II�1F�0D"&���$UHѨ���Xؠ�c ��2�ƈ؂����b���$��TP�"�A$lĤP�P&�db����ĄQ&4fE�F���f�X�!1�F`�!�M��M�
�iM�2#$���͉����D�2)B��bf�Dd�P��]�$w]���3ss'7$��p�(Dhn�"9r��(�Hƈ�&�]�d�fi;�a̄��d�(!����z�\�Nqְ��Snvm+��WM���R}.�Z����-��T�#:iW����6���޵����s�W��q��:��������;�$�Ƭ]��Խ6�ꡝ��*<I�W ����R��[��~�A�v��N7�ש�L�{�zl�����SF2#\�;nc�¥L-%���P*
U���Õz+/�����S�O�6�Ĕ�8R�������09��#�� 4�a�����܆�j�,i]��#4�i^�kt�\���76�n���2�I\b�{X��E4%�Y]����ɀZX����F��Ύ&/~����'1�d�%��v�{�3+u!ϚY����� /�P�QJ����C�j�.�oy���
��;4h�7�p���<�w�J�=��S�T���C��Y�K����=�Zʖ�)����������~s��� �ٖܰ$�6>�ו ��'����������Rn�%�fiT�qu\3xXa�K�Sp��f�/���Uw��UZڱK�x��7�f]p��X�$�K"z-k��[���`��ѿ�vձ�zMD5_.7����{�"����0���'�Yرپ��N����v���MTąR*�K����ҳ�U�]�h�P
୾�����Ѣۼ�;��)'S���m����'x���Y�̀ =��B�]tXu&r�)�	�e���������)�Zֱ�2)jwrǍ9���������t�m��U��u\uM��D�'��@/W5p�T�2��1�����u�l��S/"[W|��"%�X�m���p��1��3�%I��R�>��ٔ���1�S,�t����M;�fWe��6ҹU3�Z���6��t١���V1	{G%���TY]XY]|h�W���)�Ǖ����r�J;�az���>�g3N�c\n�Z>����m)�l��r�v5�3s+r�z�Z3b�[�����o�n�znntu��ƣ�$�3���<y�ˠ�\<����+Ny��O����-Sßs��m�c��{�#mU}ΨLu�?�{ٗJ]�f߫�f׵W9��s"�r*�mX�2���X�,��;NBrm}m�9�f�٠$E�Э�N�wW �!���'h��Z����B:��_b���)�f3�&��Y5b�����d'�@]��뇵��Wﱽ(>H�|��Ƣ#=T�:���a�|~ڎ}l!w�'	�4��3r�=���ڀ�Y�0�c&D�`�����.�'5t:�C��U��b}g'4��d��$��n�ǳ���F�Nz1<�yf���j��kleՅ�3�v�,�Tp;�j��Y���"�G;6T�C7�.�vC�E��)p��=��Ь���+������	\f�S[���n�f��
��ٲ�kod(��#ﾏ��n5-gK�Qw�4~�7S�G5L���^E�uD�N�#��������l{;[��ϭ�8:1E
���Q�屍��61�L�0�G*Ň��1���姢>����4���\�k.V,\6��RBu6i���͇�� 9��䂨uݘ`B��i9Պ�F�;}���ѷk�@U;Bv^���W3[���HvFk�-���Tqq�o�:*X��w�
TX�*p�r9�q��>�B���ΤF�Yd:�p��7�[N3������9����;i�9�
�[�^�W{n��W����xQ���'8�D��y8�T�e���H�p�;�[�l�E*�t���p���vY)\��!\'�s"h��7�*z�]*Xr��Bd|���!�qN���i���}K�m�2�q'I���Bc'R��D���P����&/�@�#_F%w8�zt|µ���1����&,f̑\��+yU���j:	8�ȅ��#�J\C��@��B�J����t\F�e,ێ��	T�e�	��u
�O57��F�80�x�MC��J�� 6r�ծ�r�K�%���o�&����6��YN�n���	���ӄ7���6t�u�,%܍�Y���f�ȣARo2��n]M��W�47�eG��d f��"@j�ҹ�E_ﾈ���^�O �>C�����_t8I(���}e#��ڬg*���,��;}}��1�j"���R��������?eGL1
$�z �dX�𨀴��u;���۽P�f�͹�-��X�p����nxn']���q<Ag��G4���p�@-s�V���T�w�F�ݖ���	#�z&�wh��5han�1lńMCn����Dc��#I
Tj�F2�b�P}m�s	f�qJ[=y��+Z5�ÓЛ��,�W���"��~�O�tbбy���"&�Q���<���:�Ⱥ�+���Q"�O2h�&�y����9���V.h�$>*�'�EVu3��?�^�?|><b�Y�P騪����z���ZbWF%���iY��}�x����@f�w]��]Aʍzm��b�ݔ��C
]�ev�o'b��ڼ~���du��4�������a�Y���̃�pn��CÀ���c�t'�%��z�UHe����fY�g>l�
��7�/,��ӗ�O 	m���C�٘v=7���+��K����9��z���|�����a]z%�ˌ� ��Z�9ŧ��y��u	��܏M����O�0:��6�U����+h;[����m�i�ɛ!�/��u8�9}���},˴�rp����5U��JW\s���}�y�z���=���L��t���jȾ���G��IW�~E��ł��x|b��oOw{���#<_��S�:hN�Ę��K,��)��n�c��������\�U��s�I˾�&�#��Z�!x���	dr%��DO�������\C=f��x�*|�_5y�M����\�_?|j�����U>Dep
�Ҏx�LƸ�R��u:c�z6�Û����y�Q���q	���g��P�'��A��,�l?����0����jB��7����C�yMϵ�ì�gU*���|�PS��N�P�v�vX��7����O�&�[��AWO��7\!7�T����O�H�p�8�ұ�A1t,�W������\����{Z�l�ߤ��5��ܜ�W��l㜬�Z�,NO-t=\�{(n��p�H�gŮ�^$D|v�j�94�,a�E��ry9��&�/���!a.�=�A�EF#֯	(i{��k��*�A�/�B����������އO�+짎C��%L]}K%C҆���]׮�K�̅���ɾ�N'���f�M
��������iC��z�ڼn�c@uI@%�����l�v�Gvm�e�a��Ȍj�qg>� 9;�e;�ۙuv�e\pV���#�1IX?}�}�UT��ז�;P��������$bvQ24�:�/�������Y��o5WԺyy�I.\�IMgK�B���㛻�h��e���Q��T,��"��B�>���.pE�Ӑ��ӆ,�<���W
w9���+%�S,GD-t�,P8u9��u"0 6����*^o7z�k=~��j{��cNeu�_1<%%�}}b��5�~�%S7���j����4$ ��!+H�`����,�A�'h��q�鹜4�d�Z���V��P/N?7��UDl�G��`�'c��V|"�ǅDr��.�Ꭸ%�'��Ϛ�=j\hU�[=)�	�=]�{(�����έ6��I��S�:�z���zlb��g�*��q��&8$��!��sF�OW�;V���|������K�Q�����0h�3�B�g�݄9�8�Z�o+�崧z�#��n�Gb-ތ�q0�cQmϺɓq�I���'��h�<Ǹ&�J�U�1����.�Y�/O�Z��9�f6��M�ꑷ
��Pϡ�~�^�2�]c�&j�dqd9���]�c/b_fդ;jVq8���L�.(Ž����nT%�O��X"놼�]hܽ
��'����}=㮥Iժ�h7��9N�Yލ�� ǷO9�j�8�ק*G��^���4L=G����
k�܌s�'�}_}��8�/U�8��S��GB.4�E_�j��Ȥ���L��n
�c��@��n��]Փ)ض�231���A]�A�`�.�]2�|4��f����dJvٌ�oJF&hv��Hb����:�$����\T1�<����$u꘡�ސ��2���:�����j�"�7-�۠��l2���pb�����#���i�:<��k���ؼX� ���v��+��w!�~�橒�`kȢ# ������-9�Dˇ9����r��:�����1�k6��O-���1��健�sC`<?	�dǊ����ޯ5�ߢz�Y����~,�4��z��J��맴�X��c��c�ݗc��o����~�$�F4�x�
�}F��/�ҷ��0�T�3}���S0���q\ʱ]�	#En^\Jg��J����@`������
����#��^�M\Os�j�m>���s�ֵ�����;ǲ���i��+���#u���^��Rv�isçx�������e2�SH��r��Ŋ�9>�׀��9U�̀�D!��:���m�����%���v$$���G�a�{�ŝ�����bG/�v�W��7O\�C&T�QK�\���"��	��
�Zic�����=�vDjWO�#E��;��,��_}�}Q�X���2$4�3#��T�ޣ���w���6�x	6�}������ٌn_"ۥ=<:���_��E�ćW�So�¥���g��ZC�G>�w����9=I����3��ai�1�8�T.�.��0��BFzZ��Vo1+�&y,�[ѽ"~�	5�à��I@���Ƽ.��<_�4&�+|s��_!�۬T"@P+5lR��u5QA�6ʿ��Y�� 1?��eX����*e6�_�gb�2S�u�NL�a�[��9Y��#Og�؇1¹�h� �~(U�]���Orݮ+E3���۴}�J�{~�f󎥽�ۿ���7>n���z�'���~�`qU��GI��<�#��m��=ړ���{��r9��,_p���5\��T���"b�f,"i�Z�Q:`�@���#6\Ԏ���o1*�q{[F�g����1ZѨĦ���p-�`E��:g�L�k�%�����/]nΖ����A��{&�jP�rMn�Ӽ�|ި��uE�n��Y�V���Uq]D���=CE�C���q���n4(`���2%M�۪�*)�F�a��mF���u����r_��sA�>���v��l,��*�u�Yk�Hvb�Y��p֥v�K���Y��<�9�^z6���^%�}�nuJW���r�r�Q_�ﾯ���{��wF3��?�S���c�(,��?Te-�+>:��q�N�7Ɯy�c�.�.��� |n}�d;@�ǌ�iXn��"����X9�a��Q֫I���A�Rs���v�vP�Wk�ZY��P���'O�3�΂0�|����a�t��xx��~��u��/�:.��M楎���FO�V��a���u�뙋�sC4�k���*�E�<�%�*p�E�]�;��0[�'�Q��5�\O�X���#ou��;���}�H]ֿ"�y��Y`v/.)xx�7/��ˬ�'���Tu/���W��.�%�O2�z����Y|c4A��Dn�o)����檣��7%����LL��ЖG"^����D��Ϻ��pkŀ����;-�Z��=��SW�٫ҡ�Fă��<+�RQ���q�S�Q��s/;�S������Ч��,v��p�>3��B�p��=�p
����R�
ۿ:y��s:{ݶzG'�%lM�V����c;��(�#�9�c���@����<�R��ӊ･c��ق�"*ͦ��:���,D��rW)24��ec���e���A5���t�s��S EI�\0p1'V���3q��.�%�x�4.��;�]�6�h��;��f�F�a������^�](�<��˖�o������޴�T��u���!qx��ã�-�p|wa����F9�6�RJd��V�X\32f��΀$���ݦ��� Fi_b�_W'I������Vm��Z�Գ9��L暨Q�ВB�H�����D����+Wi������C������Z+�����S4����P�P����_�Ɔ�R���5ʼ�h�����i��C
X�I�鍚��m�����a�����#]�Q��ْs�<N�����U}��w9{����q�õ��+��7��k������{͡��rS��.�y`�����1��]($>�棧Bŝ~(��[���מ}�lh�Y,r�b9k��qb�ð��Y��r���qɩ�pOIG��tu;n������J/qt��
��6���>~zM5_.:�`����p�W�a��]�@�����:�\� ƿ�� ��'�ïM��+Y<l�Z���ҧYd�)@�,Q�,�z�q��~Ӂ�Ō��h@�"�w��t��������*��͙@+�5A��x�7,�*�V���݅iS���1�m����%i)U��Q@ŵ<�v�Q��q��)�.���N��mCK�]�y�rq煩j�y�ʳ���r�u��><��B�ʞ]��[���5��D�۽�}G2�삀�ė����7b�ͺ�܃-#�	���_2�lo+v5��rq�-n�f�E*�h�PG{)�Y�n����څ�7���6���ksN���ngb�V���c�p�9���:��\�Zn��1!�a�0�w��dPB�8�q�����dV�ľ[h��/�.���ӫ0E}��-�|�)��t��=oX+kk�����n.��0u��e^hk�]�y�Y�J���^,���Ӻ41;�!��	��utղ���I��!
Y�G�/��,j�I�-c9��&���;sK�R�TW��b0�apX�ie+nY���+r\®`��<�۝���9L�.��F-8]�ڃ"Ml�޴�P6��㗛��l՗�MܩgMPj���-�{A0�ٰ�1n�����ח�1��Q��[���;� ��%��2֛(�Nr�aޙvaFb�8�����2���iJ��IgK��U�`N�c��(P�T�ZpbS*�Y|U�]6����m�%�hⱹ5����R ��r��]�a�0BFqS69e�5ی�i]]a*Y��f�39X�l"�����[D(��e]�@IX7���)��rd�t�n_P�ˈ��s;�n��I�j��sl��c��87Jr�*ύN�@��,pu*;���䵩5��Hs.�Ƿ���h���P���en7F��[3�N3/�0�A��|�ˬ��ݏt��6:	Q�Lʂ����L#���ΧS6���訄��Wl�>M���OH!Q�w���K�5�5뺚YY&(��{��"��<C֥�|Y�[�b��n����Wu>�l5A��������ǝ|�9oY5�ي�,��.�u):��ח�h\�b_:�ܕ)pM<��ڛ�uݛ��_'������2lԎZ!�^`���y�q�[6Y-�Aȵc�gG+B&�	9Z5�*i1@�-l�0o��[�a���)�2��˺��f�����0�#pN���i�B�v<�y:��<�*QZ�ʂ���w�#t=��K��#{�>ba܏j��,�7dS�+p�x>�Ժ6�r}��֫����p�\f�38d��V���(�h&BP��M�"�2���u.`"�p�m��\�$cp�둂�C0^9��Pɲ�KF!G��L��]�[�]��}�)�]��Rf=��f ��i�3 ����V���S�-^Z�cx헽;��Bf��g&���e�w�ܑ`��:��M��V�.S�իK�
ŧ�.qn*|4Km�
Ėh��~,�����-�B�vL��kF+���a�ٽؕ&�Q��S��Ѯ��2L-�Ehڗ|@�} ��#L`d�(" #D�wpt$)�����Έw`P�F��2$���Ȏn&	�hB32HW."�M���(�$"��8���\��Ww\܌P�H���!w]��!�;�BDf]�K����Za���:���r�ݹ	��q»����˹v͝��\�.�0��9��9�;r�%"��)��N���Fu��Ȓ.t�F7w]ݒi�& �l���S�K�v��Eww���t��ܲY�I��pwpA"��ۻ����t��dE�w\:\�F;��2�1�9��wqC�u�¢w��Z�U.��w�����{�������M�Fq5d_�� ������}:ĵW�wbbz���X���Z}2�������_z��<���$��=2����yƥi�t��R��8xsK.C���J�.����d���K�o�����p�����:�� �q���R�Ř6`����77/�n�*i�(Е:^ns!��f��ݺ}�����ʗמ`v�{����+Z%�Fy�Y��7�a��V��3�C�mQ���˸�n���J]���!��r��z�m���d*~9�=q��\�U�g�Prt� �yCQ�)l��=���X�=�Sv�^�+��}O>8)��]����
B�����k�	w?��J��ƶ�]\;"S��S�p��7N��`�;P�<�&�qp�cTru����J5*��@�"bO>�\���a�v'kx.�8$ӭ�iZ��?Km�gŵgƀ|OJ��*�Γ�W#�A*��,�}g��[�x�Sׂ����-�R�Z�C韷��K`�1��# N`���̀d-1,!�N�㋩�����;�%��ڭӑ�m^m���1�6���d*����X�g��;��hٞ�G{o����.P,��tH�z_X�L�Z�'63E,*�K��fA�"��mp�rl�]K��vb�Էj�%�P�4�[�&�c�Rܟt��w%F��F�;GA �IӋMɮ
2���d���JfaNhp�$�&�m�bI�[�~������Q^��-M��fM���e����/��2�.
�[�oL�� <�����J�"���{�=^͡�;�y������,o@��T�1��WR�x���\)�zbh1KmE�L\L��wQ�g"�N4���]<9Ƙ,�<MA\=�9Ҹ��ΆN\gR�[7G��Gc�]y�m-�ʨB��{"���;�cj�t�0`5��i�'jb��B���f{_�
`L[v���+N��;����ݭ��m��^���W�	�U�Z�7UQ{%A��<������gb��m��T���ʥ��6�Ց�e���/�ǇT�=� z�&��
l֘p
5�]�ϸ�zs�?0�CfKTƊ�xrz�վ=u���SW����4��t� �G]uM.5���~��hMF�o�s���w��9��E����R��K֮8L�����fll�~���X�E7_��Q�J���O�on�g��]�y��TA�~�s\+��<_҈��$:ԧ�oܪ��l���+�����j"Z)CI������F��Xo�39�k�G�ʺ]���b�,��B>����Yy�ԖtϜ���݊�w ��L�t���kuc����etC}����:ք�2�m�妶U�$�������7���J�2#�:C�MW���m��4��ZkЙ��#��;�а��P=Hɾ��O�y��V�#�e;��r��pF��MZ�D�C�Cn�x�) �5���*z�-��{YQ�e�F'蕴��t�z�W�(֍F\%P��n���0��c f���}�츼g��B�Ea�|��3������Dk7'�F���e��v? C�<��ޮ;��g�w(����pՒUE\u:8��<�;Ң�~
Q��Vs��}�阽��]��>X���9�I�r�n���zV(	��t��
�R��4�dzvd\��9��V�ʪ�p������!ƺVy|1W��î�\88�2����0�e0b���.ેFid����_ *7C����7\�s2/��~<t����F����_�y����x�Ń�>�!pI|N�0�!z���\j�����]�h�����R�~.��(H��S�'f
����|���
��d�Ĳɑ�s/pS�8�����/��ⱕX��3�Z��3b;K�'7.��JkW�t֕-�c�f*���
����ੱ��ŀHU���e$ؾְQ���:pT�B9*�\q�T������Ʋ�u�Wue�'T+j��j��o4֩/�2�keO�ui�����{�׵�R�ZFU!���#��$�Q0s	h���^��������^�Lwog$��z��	�s�m���Qp��V}M��f/Ox�$�z�Y�1���O���+�W��)y{%�u%H}��X�6�a�g��1P*�Ę�! }��!=���'��?,;ZDOMd�.s���F�P�+j�˾5��V4Y�D����l-�{��:��C�I�9!R��>�N3���'��D�q�ʺ|wa����c�����������5;�;A��,{:L�� F&��Aj�qx@�җu}\�$p���s������h �����/؄lX��'t����_��w��Qt:7D]�u�X�z_���`�I�:����������&{��r�$:�CJ��U=c^K�x �_�&'��?m�+�Eg>X�ݙi�b��G4�Ѵ�#]�Q�_l� W�Q=_���f*%uF��o[t��ӥ�щ]�qc��Ѫ��.wt/�X
e���꧖��֯U��`�%e<����G�b��4�&:
Y0�W��'83Z�B���c+s��^�q��Z:�\-��#�����k�u���1"+_s�=�Ľ%ñ3�(ܛQ��=N+�m'ǰ/�f�@ՙ\�^-�r�է�]隲nR�F�O`��J����p�����NC�_W�}���d���N%.?;gѷ,B��cY,\r�b����x���,/���R��}A^��-�M����:��W�2"�F��ݾ�0L���U�㪦hU@�X���B�F蝆��W��e�uҁ�">��r���;�:{�
��ȭe��c�.k�&�*&�oIu3f��K��a�3X'��q.�_GIy��\ǢϫR�;��ʽ���`�9&�mk�+Q�x�=�<#u:�c��:j1�Wt
������iװ�:Ê���ȷZ��J��G�.�,�.��C�"���e:���]s(Ѐ#6ɒ/췼��-�=\�=py]�/���W׺حϙn�f��C.1�m��鹹����k�ݜ�a�'T��f%<\�$�~��Z�h��7��x2"p��
[�`v��lhjG<���~��+�87����U���#�*��k�����o��Ē�q��2F_K���bqr}��R���ˉ���*P�^d*R����]t���ڛz�X6,�i�)�!��^�;P�͡n�)�dL�Wm�A2ˊvլ��R<��*�-�f/sBp����j�+�.��D�v��;&�)w�Թ�9�@��gs��8-]�#AU�SjY8:�F�k�2�V5#9q�Fퟞ��pÀ�y1��%�DG���\��cu±r1�&��l4���ې��ʌ�$x��^��_�ڢ�ZO�{�}zO��o+���+E���S�a[VYρ�LOѐ�Ua�2`T?+�·�zmr4��7��\�Cd��)���\�!����S%�2�בD`�uD����y����8�����k�yZO�3r�;��Hm^m���1�6����@B�����\��/�rC�#���Bc�~��f��0�6��ǠRe+4�:��Q�΀tl�x��e7ʧ���Yv.�k3����ױ���j�}ƙ���%<j7+�^i�W��L͗�r���wn9,���OL_re��"���N�n⳾0��=�,�×�f�&
�2��ӷ2�/W77����9_r�T>L����E�����໗d���n�|�*Sw쓽Y[�&y�D�۽7�I8y���&�D�zd�xΔZ���^����-�m��/�\҂`�5{HS�"ʋd)�<�D����ky�׃�^N$�s��z4G*��ؐ��\���AlBޝ��r���TG�e��n"2�ǳR����.�;9�+WK���z��
���p&��C��d�2�.X���}��M7�꥙�u��q��z">��y��e<���w�Z	X<�KꍥWؕ+�-�8j�6��n��TY�~����{3�i��yc�NQ�5~p����k$ ���FX�C����O;z����S�ѩ�-��6���r� w3P5%p���sPr�`�{0�x��싞.k/�����)P����
���Qߛ�I�0�m�..���|�x�ho���܈otT<gi�2�]�X�=}�VT�>eCV����٨�mnG��\v�4�7��3hT6�3����j �SO cV���6q�+�"^����W��kG*�5�&�;e�7�oa�/{���	��U�<��ҙ�a�5���S���C����������C����Ѩ��.9lj���tC�a�*|��Eg���Ϳw���@%`c��u,�2�su�\9_[P6��_g�k����P��U�C}^\E("���Rn��r�b�˛�vs�3T�sU��6{��!Zx�P���\���=kf^�3ۘM]s�4*۸-ҫ�����G���[C7��1���9�
�"��r�:4��;oD���VZ�3Y4�R��V�N���ޓ�q��ܒݝ�z�{���cZe�n�a4+�˝F�c��R�k�}�F7�U
��!v9����l�@>g�_(7��n�	�g8�|�/8�o���Y��*��nM��h��ٞ�Ōѯ�$�Z�'����\�i�����#p�{^�56�n�2���
�{��!�PU�@;�.z�T5z\,��i�ӨP<�ބt�	�ɹ����N[O�j���.�P~�
f��!���<s<e�
\4w�Gv6��{y�(7���q	�����jh��/����7�5w�6�.����*�̖��{�o\5��8[_6��/ܨ!���J��g��lZ�s�9Tv�֜��-鯊O/�5ٮ3k��q�d��ܧg+�ΰX��9Ȟ��[~I�z@�b��������XV�r�m��	V8
�m�T�Q��*M ���!�KEi\�!�\sy4���[����'#��w�ö��H�a��1v��q"O\���:�r��2u���`�$�H�x��Ũ6�Z|��F�7T���
k���6fi��X`����11+t2�y;]��ͱ�嵽:�@�Nٳ^]E��h��^.��W�G7]/���ck����BǏ����������ݞ���� +�ͪgê�ܥCA)���˷r'���+�j�Si�|�S�ݠ��,���G"aR�l�ԎЋ�6>;�iŻ�rY��Rp�N9��	�MDsLM|��v�Dƻ#����ky��W�k���9���a�ܧ��T�ԝM,p��p6�9�V�"cX�{!=���'vEK����c�j'��S1y�~K�|���ؽ^ǵ��G��+�V\q��F�g��Ⱥ
7�	��]������W�E���|���{�p����@ˉVv57*vF��ֽ���c2�.�{M�P����b/�1r�{4�q����\���8��ͬގ{��~���4&��{8��撌��\e���k�4�Ls��Bi�p齸�Ҟ�����	�VU�OZ��%��ڵ==��p���R���P�Zm��.{Cٌ��e�M�욌9�X�$��՟{<�+�Gٻ{�N�<�]��㵉V�ԩXseo�A7ζg���P���e�ޚ�{#�[d%f�C~y�2t�ͤ3���;�	e�Gyn����c+
�\�.la��9�G	U�{��Ϊust�6�̦�Fw��'��}��pݫk9��zݩ+kj���A��p�^8[M����y7v^�*�(voo)�9�g �|�l���貖�)<�e�}��5��Vw�l)�����V�Hw�|�`��b�4��!mo�����K���f�%�ս��U�'���*}����>ﻤ��q�5�gNu�s���S�z�����۰�R�g0TCl�/�ʾ����h�E�H\�=L���j��'��?�O���_���As9���<������y+f�Z+$�����s|��y=h��o�y�����r%; 0#�n�5{[�cx��x����U����v�O#��?jx�SQ)��q���YNN���2�W��.�=�v��b���/>��4���sŚH1^���8�Z�zߍ��Yꐰ��D�p������3��#n�h��MG�V�J)�b����.�H��� ����v�ol���)}�����$ǧ%V��K�ݹ8޵�����L�(І����e�mS�Bt���s�G��� ڛ ����Y��,�{]��e��듘��6�;ݒ����5�,זo�2�qئ���j�!�)r��N/���(��׈�8�IwMӗpXw�'!f�=Α���w2(�2�FM�<�\]��j��jK��A��W
�dL�`���O��=Z5+�Ώ"Z�QC�;�9�@�ڹJƃ�1��aI�ʽ��_%G�r��x�;.�ڡAPz��W�����D��kA֭ZM�M��.;�B��eB�lv4��M��V�A{����U�9y��wNV�*��<tm��
V���R��Y:��W]t�w��;�u�j^jv,ݬ�1�]Y���� MXY{͛ ���[�4�����i��t��yڛ��/�QÝsT\I��NG~UW���b�:ыj�I���qta*���${��mB���ݺ������vs0t����qI���{���syѕ��Bl�*�znƸn��aS���-�\'b��Ҩ���;3 69��,z�q��L�7ڈ:M��{����I&�|���{�w���%�������Ty]� ��&b�29xv�N�Nw�X�r���Q��q�7xM�d�MQWo:��s-��x윴.�]���������I��):N�Ӻ߀�9A鲌6lV�r;e`wf��.GG�ݧ4B�sG�[�5Y�ב�Ж7r%��J}W|��/Jy|)�W�ŗ�=�RUq�&�싴;y�3�V�[6gRB\������f�h�[%���5Ν �7@��Z�������X�Y]�ݪ��v.��� v�&֞�%����<�{���%۔�=Z����.����冷��(7��Mm�fA�!{��}n����(㼧7�g40ֹ
��C�@)u���:�����s���ҫ�j���6Vn8�I�4f�.�I���^�!�iaR#A��&�Yc��;�$tn�܂4@#ݼ<�;�x1�;8AO������Q4S'Z5�*�`�P��[u�n��*ߗLn��s�;)�a��$lQ�A�o	Ff�r( �:�"K|.��^2%h޽T�M�n��/b���1^���5���1Wo,�Y҈&�c�6�>�qV��c�u��u�#j�[Y��T�r�*��A83S�m�iF�U��YV�s*V�,u���)vP�2@i�����ވ����b�-ⳑS:J��{5���td'_�k1�F��ɣ6�STި�u[z�f��7��C���k����	s�a�ԝ4d�W��ʶ`s]���[�Y��|&�B��q|[�!�h��H`�p��n�/noem�e7�v5��Q�XByv��[��T���F�,�un����ݴ1�툔d,��D�v�<��6�eJ�U���ԓ��>LM�d�]�F�':�� `��Gwi�E��c��!�7N����u�uܐ�wnWs�$��u����s�v]��v\���wH�J:\ú�i0�w]�wW��H�ݢ��\�G]J����ws�t�ȹS��ۙ�;r
,cS��v���P�#��W\�:������Wf9q�j��wn�ٜ�&��3;���'u���M��t�����8�̛��r�����R����.��t���s��v��7w].˺������]˦n�된�'u˻����G�h(�@��ѐ3��j����}�h1��nr�ec��.�o�&0YqJ�{���N��;<c����x2_���Z�r��C�oLsWKE/��^�sq�f�Q�6�U��.��f#F�a^��[� �4s��敡�o(e��L��x����yݕg+��
��F8��Q,���{O���wn��L�M�齿�v�Y�w�g\�f�e����⦆�;r�OOVӄ�L�q���7��m�ľ|~�g0	�at���1��%�D�Wk(?eXp_�R2��2?���~�W��gfq��x�9oGH�q�1���m���1NQ�4=9�=޸뢪%*!��޸�8&Sδ���}�(kn1����-�iP����*�j����a2'P|���ݒ��\\�9[Z�\f��r��_
������3I�Fs�ʤ�9��8v�h�Tb}�[J�;չ�{���;P噄Bӊ��Z����3Or3�������眎*���Ҹ�v͡P��ڙ��Xy�nGP������~�r�Q=�ܩ""ÑyE]�_�v���˛�9�B�<T��Sd�c�X4 �Ⱦq�B3@f�=�*�Fs�XKjƞ��]eN6݄�̾��_m��D�੹M��;*�B[zt�=j�T�<.k����ާNJN^!�hG���c���j��N����9�M�q7�&iND�']���Jz��Z�J�C�bZ�ۉ���9g}���}�b�cJ�ַ��͗	�ی}��k�&9�kk���OfVR�7��<���ּ�w�ʹ�;M:��N��Z��E�jʭxn�5��k�f)�6��n���x����;/�^ѷ��nV;�R�����R�|���4����]���S̑�GpS)��ʈ���^g8��|�>S/Q�����f޽�Ǝ����u�%=�3D�2����h�}%1�l_$*:Zlc�]0�S��9��zi�u'r�gk����}HvP7�%�TN�kC��[X�'g�;(��3�9�Vds�z1缾�<գ�]�~uV8<�#(J��ammh��i�)�kU�\�"د��Yp�}q��VW5����YB}���h�3l1�So'`�;�T:�ɤ��m�{��K9�S���x��ηΰ����o9���5a�B����U�^;{n���m���eٌdu��u϶ Ĝљ0�bE��oQwH*��rS�XWc�b�G5�
5��������]䌎�wJQ�j9̇ݾ��<�����\5��mCi����P�`t�G7a��[����l�f/�߫B�uK��%�4Ryq��qy�8�B���lkǉZ�W�ŋ�� �A�_��h��V�k1����ž���ۍ�ʸe��9%�]ӯ	�)X~�\`��W��BEe���	��0�9�2�V�Ëf�%�F���&�]���C�P���t4���jt�ʡ;��5CT��A��_wRUF\6��&�;�m�p�D�*Bz���\��~���L�J8.��6[����ok[.�o�k�bSq���^�nZ�؎n���1�*��j��4�OՐ{�_v�O#��"��'�{�X�M6�msʯ��狾|%=�Um����O���n*�'�습v{fﶷ+"��Z��^;�l��Ԝ¸O �o���6�U�%��!'*�~����9��r�����7�Y�¹ӓ�v����u�a@SR*�5.(�V)u�l�`�{lW�J��ox�Y�;*�#<.���{�j�<)2�5��Ӝ3X�f��f^t����3C��wb�`�;�v����Zܖ$]���b�65'Xt��m�2fv-iP��ͧH�w�er=��nr�����(Z�}�ݣN�棷)���6�)���z�ᵽsެ�9�]�Wz�\�v8�ݵ�{�Z�C.'[.��M�t��J��OUgaڦ;���ccL�<�A����7���7�.���`ltZ���o��|������tw5��vj��(���=�T�\RT�Kyc��,����F�"�z]��H�\H��������=#ƲD�ݴ�^�s	��P�Վ�nU�.5#�Z�C���T'����j"����5���s�����o)�Y�
��QyI9FQ
c��W�Ef���㗛�a�/�|�g��pL�&[Mu�SJýK!��P�;NY�D.!,/��[�A�6��sv\O.{����s����p͠��r'�T���u|��}�Y��׾�N��I�[��j3kv�����k�df9�_<4:�����P��D/oo{Z^ʞC�G�#��F��Ҳ�%M컭(�:�E�N$f�$��v�餮��6�=j�d�`��l����u��\��X#b���$G>x�x��ڝ��X;��m���+\�}����h��gb9�-�#�J��0��0�R��r$ep
�T��Ns��Yѩ㿛U5�,p�PЎ��.'u>x��A�h�W��G��W���U��SqǙDۡ�ӻ���ݷ��6�o%s�u�t�	9}o�o�E_gU��s�������K�֬��sfg%(�Ch�NF�Ѧ��� �~�)XF޿Ri��v�z��y�m;�2�qo7[����9��e�L����o�=�\�t������*OC����&z&źon%v����d���+q�]=�ҵMp����	p5�K���	_ѦZ�-��I��m�7[Q��o���n������PՕ�&]���U��<���ɐ�N������gT��ب���iu�-=�{�(w 7 ��+���뢮��$X��@4�F(ܳ�9�X�^��%�ݠ)ͮw��ð!KF(wQw��rDa��CFn��98�i�B��i�;3-��i�iƆ;��J�����v�z�nf��o#a��s���`���svn�12|�d�\��O$��ԛ{���c��9`��P��O�A�w3^k���k=S��r?o)�W�Ҿ��e�,k�\f�f��_@����ɚ�x^�����S��\��@����[J��ky��3���x��2��ƓA�T����.H5�だ��k���r�X��}ɥ�;��Cqut�?n���Մ:em�����=_�C@Z��yv���u����,=��le�w�$}h,�=���㔹�*�Ty�h��k5�n*�~�S^�S���������Je��&�MƴdF�"y����Sن��r���x0�(b�����V��u��m���W���F���U_|���CV��^�bP%�E�[IO���_Z�ֹ�=�UF�eK8-�����������^����e�;�S/Qo_.u�Sڑ��Uݎ��Y��LǱ7L�z݇�0�<y^��^˗�i��w,v�mI�ב7�H6g%y�6^MG$PŉP����]��[�ΩI�x�owht0�)�c/�-fJҕ�J5Մ`ؐ���G�n��3�ܷ+��w�mֹN�y�h����N����b?��Z�;�n|���i�on������-|J����/s����5BmZ{��qJ�W�Q���D�&�5�n�b���FW�5��6��_f���7(��`U�I}GLSź1��^m�kU��\6�^��D[���o�Z{pof";l�Rg�����=�1p2�GM�᫋�D�N�]�Q)Q��c����i����U�fne�/������c��pv�'�)%�
躖��I��ƻ>��8��װ�y�U2���B�����%������;����u�o��|p� �9��ʰJ;xmGK2�S�S��KF����u��*�׀���zo��s�5���~�5�3�*{�D.��JUA��MDO.�������ݮ�i��c-��r�GП9��|��G"aRH�Πu��#/;ư3T�Zf"w��[B���4�ޥ�t��fIՖ_c았�yↂ���v�/mu:=�h�I� x�#rf;~�3�+;�ַQ�,��E�;QДsM<�{��%�}B鎐�%+�w�k
COE��M��V�w�s�����)>�̥ |�Y2�Y�wm_��j52������bi7и�Dtw���z��ۋ�9A�d�	cݗ�8����j5U���M,p��p6��*��P�8��-zd9*9'"��EB�]�A;y����%پpy>�1,��a��SNԩ-�틖!�{�7��6����I�ߴ��Ϧ��_x%�r�ar0'�u�uϫ���7�g:�^�F���E܏b6s OxtWTRSO9KCm�9�ldK���޸�{��g*9������S:�X2��ef�ޝqj�����TualsM�齹]�p���;�z�"��=�Ҟl�N~�3�a�����5q�Ҽ-���5������������[��2�^��M�δ?AJ~�ٵNU�T�Kyqᬿ���;*rm�R�AM>��*f��Ψ���?@|�K���)i�)<�r`�����$1�5
��ݷ�n�Y�/D�WK�I��F	�V]p㻸�c���r��������,�:�.ݸ5>�d{�0wk(�Z�k�hԮỺ��Q�fm`#s�IB�m։0���_!|EI�g[OE���mޘ����%�ڒ��Әz����}����sjd��6���P�>���P�o��`��'��O�Q�d\�	rp���8ͫleC�e����K
Z4S`f��t���QuO#O5�vj�bx��ক�z�c[gj�(�1�o2�u;�g~Uˍw����ݓ���[���k�|Ն�;�f�V�D�0<���>���*CĞ�w��ǰh�}eu���SSk����������i�l��|0�tpe��H�a�	��D�m�rV�\Nsڼյ���M�}�5�)y6���B��L�NF�屩
��xD�|/���׳R��L��'��ej�:<��2���r�i�q�Ts�u�H��1T�˂�U#1ot�v���=���
e��7�k���6�Y���3* ���ۣ�A���ܝc/9��[N�S)��:���u�q�z�ʳ�X�(3_�@�U��J��c�6��f�α��L�u(�Ӕ�4(4��eLΉp�vqXn��F�m��Lj��[C��Н]/+s����qo:���Ǩ5�r�P����G;:��qcf*J�<�˚�v\��.\/zӮ{Ž�򮨟G�L7�����ꉹ��K��TO��2�6Λһ;�)�T�O�Lɚ���J'O<e�j��uTK���P���e��ب�I�ܽ�+�)a���˫�����f���dRd�yT��J
ĥ-��3p�<��O�A��������-=�7�Q�O 6`�0*�)8ZcbaۺU�wGs�X���	7����-����Y����^i�w��d��\zl�ꎼ/��;{X�%�5�ˎX�dk�מ/>�� �+��d�2'B ���~ѧ�����b�JK2ި������w�q��_<g[q���{`�ٲ�S!:\`�c�:Vj��(������+�w�{�ڜʻ��y��蓐���j���<�V*�^��8��Nx�/A�<Q����o'�]��˄�2�����2���X�5opE�5����ۭլ.�U㬑r۩*6Pl���ʮ��ʉ�'Vw3&n(�+Ӯ둑Y��c@/�/�]]�)%��P��U����ɚf�u�s:��ck"��h����b@Ax,iD��mk���'6��6���X��%ƅ9��H}'����o��3�{א7۰�e	���]�����G�ӵp�TH^��,V�Fk����2 �p�7].�F����Y� ����	��C/��)�E���e�vv|�Ixw������0 r��'(JTW7��tC[A�6.MK���#�a��$�˓�{x�V��wf+���������O��ͬ4�mG(����/��g)�9�
��u���G/�5R����U��Z\�B�q�✚�F������`
�f�Jb;5����(��t�*�6�����&�}� �2�k��ٔZ���z6E�0����4�ƌ�Y)79��'�P	C+�����S24�<�}S��Ƶ��&Z�lt����V��Kh9����cZUL�'c���]`ᤩ� jK����i�¹���Sl�bK���5|f��;�-mB�<ʾ4�-�wk�.��� �W,+Gs�����z��hcP2��YV
���g[�چ�SsdŮĲ�ܮW3��'B�5��&F2��/�33]�52��.�6�tWW^1�W�89͕��Y9�I7X�/f$һ+m9�O1n^�Տ5��Xg>�p��)�jw`��7��Bt:��9���us�
tΣ̬��yˎ"����X����]��)h0��}�µ�����붐o#$��&�m[��cR���tSC���Dի�ĉ�ؼ
T����1w!a�D0�R�]�hY�4�����k)����0b)�&;t�jFb����Ӡ��6��Ι�I����2��k\�o�KbNW9l�A��bo����uJ{{��`���YsC�AX0>�:�A�*�.��n�#'n��p�UALm�ᛕ�
n=�	��_�ɷ{���?9�r^��v���ogR��^�������݃�M���u`I��g_u�e�@��轹�Pn���Ɓ�ǹ��$���uY�1�\�Nķ��-71M-�]��.u( �`�Iv1V&� �mm���o1Bڱ�Qo ��%�mDH}�+r��"��V2M����C"d���٩��	�!6��@û{vH���a�S2�e�Z�R�B���3&�)�4p*>�V���Nj��QZ*f\!#�(��]q����7�L�s�q
��ɥ�Z�T�6ݎ`Lj�i'H�/��. �J�ڕ�ٷ)�Fei ��k�}֝=�1V:?`ݗ���(�Ƶ���
-���/(���f�ڛͩM�)9s�7���8�lVPu�2��T�d�1`��Sc�����3 =	�f�:������z�����?�t���s��u��N;�\�Jw]]�'nr�n����� �C�vs��L�K�u�rC��19w��r���]7]w]��waNq��u�K�K��Ww3�;�f]ӣ����G&D�B��˸�l��)����� �.�s�.��9��]�fD��۲"�n]E�a39�vb8�����7s\��%wwu�r����a�N����7wM�����Bn��8�:]�wv\��陗8��9Ҋ%Νv�6����@��َ\�wc';N��˥$����!t��7 ��IwnFNGI�҈"w]�gN�7v���]+�e7]��Ά.���N滓]�twuۭӻ���ۤ]����ݻ��f�]qˑ�B�T֝n4�L�jOXs�>�6uR�S����� =�&��jWw=�"ݣ�C���6P�!83��n�F T����Sת��r��7�i�����n5�#7Q���C�����d�C�i��$�k�Hi�����y�;7�u��Ú��m7�Z��k#*�-����{�*n��߭�~�}ş+IOO�w�����k��r�(ٍN�u�.j�+��`�w)4Jp�̨;�1{�	X2��Q?F[�je�9�|ֲ��u�wVG�f�_\��L�ꉖ����{{m�!1�T_$���Ð��枵zI/՞M��~L�>���?P��XL˞�� FsxaJ:����Ʉ�E�P�or)��/�m�LE휨��ǜ]C�ܞ�]�����x���z����H�+�p�\&�\���7��{)����A�=�Vv��f:��GO~{��L�{zᬼp�����6�\ln�\u¥[A��2^��~�0��+���oMAIǾ�핞����]�k0E��o:�J�����S����nNZ鳼�#n�2,W�k�2�q)KW@.�;�PO��UE�U�6���b^��kj��&�3k�6��(	��m� \�77������u�B�<ﮚ�[��f��eg&��a(ޜ��\��3hf۝�ޡ�����C�V��ͼG�	��O5�gZz_ž�=Y�n�o��
���T�"Nf8�-1�Q@+��)������J��;˭֛d�������I��n���[�g0T6�)�3�"T	J��O�[��-�g
ָ��E��"�}���s�5	��a�#�0�	�G`ss#�a	c3�ގ�9�S�Ģ�vI��/�2����bjq���vCmЯj�;�F��r=��Ĥ���;=����{W�jڈ�V�u4�m���M�ev��vB��
U�C\:-n}3���f/>oȮ=�s<㏅&$���^
�oy�r�ߪ����r���N�=�r�~�:&��Sƅ���3�{�N�9���i�\�o{ٮQ�����ֶ&�;��*%����]��ps	ŷϡL�`�Z�f�{�4s#�̨*���Z3Ղ�W� �����9��b�U=�.,��B���}wesR�1�L±r�N�d�y�~�\Sf���⅌b��%��pC��#9 ��{{	�2�i�ը"�F��������ha(pk�3YO7��T��].ڔ�mEݭ����q¥t��#�,j#��.;���)��i�n�ۉ]�'�����u�����a����V?`}_Fӄ�4�W��E�k/���|�C��w:�z\ף��,�����*��=�2�JS�Kyx��5�r΍[S9�ʧΛ��c%�]�����@t����zG��fl ������%ϸM�?�C[q���8�B��P���Д*�OYBI��u������4��Ѩ)�XV�r�ڋleC�g�D�7~��Jz��J!y,+��U�~�s̄w�woҸ�,g0T6���Y�DuӍ\�B��<�}�����뚝\�n��ڎ|��o��ml�.���~{I5ԐJO׈z����5{rV����W��kE�}S�0Ә��[��;�#�{E�޲'��l:n�3��ڮQ)��в��A4t }�v��ǵԨR�ffVі+dW�X�^^3��~�f�*�#�W&�v����fZ�11�+�X����Y<��&��1�B[�;���>d�p�tr���!�[M#�����S��:��B�O��stm��bCp<�*v��[���8;�*�X�ak아���Slr�Oz�{Խ,r�#|2P{�G���*����Iuȭ_���ٮM�S�6�'Y��']p�Ú�P-��D��+��|��DM�(����+�O:C��V{�nO>�2����#<�)鋓/87�i�:}�O��E�=�̦6��np���ﳜO�m;�2��]p�n޽�ز�=�
��������w�;k�'5k=^�������/~�E��٦��'pgio�~9͟��}�gj��
�j؟OTm(J��W�����{	�e��*M�����g���X֎4e�σ�[�X<�#(J��VmzӛU/q�:�.m8E��p�\co�O;�{b)�j=��_��x6=��t�d7�oI��j躞TkR{q�ۈ�^r΃iT
1�>�� �0��]��y�9����r�n[���X�f�ͧ�~�I�r�?;��h�Z��m��o+=B:�X�C{ֲ�#�]p�JY�@����s/r��1�3@���\)�NR�|š��z�@yFۇ�u�Ջ.�]S��-c�b�����D4x�Z`�L��?w��~�8������%���FM��+��/k�5�����\��b�⤃迷�m�Ti�!�O��i_�ޭo0n�03��ei,����"7���]�S�ҕ��Ŋ?.���0��wn\�Q)^`���o.�`��z�Tk��A�͉�B/a�q�����J�zjaS�|���Uʣ(����7��.1�q�
���6q�\�Sb.#2@��y�S{���j��ou�m��Y�Jn1�3u����Z����b���^s��zVA=�q�;ɝ�P�ډ�\-p�ځ��UF�7XqWm+�;�#w����ؔ������`Ǚ�Y��)|�ƾQ���{�C�}�(�	(��Sl��$Gީ:U[�*�I�[Q�|�fy^���	Ԏ_I�FL���<��L�e��v=���V{�`��Ϝ���O�a�Y���6�}-62^�mf��g�|��|Dܰ��c���9����$��In�	J2��`b�#��._3ܖ��i�Wh�ja�xܕ.��w-�	����,�2^�r���֦w���t�.�}&��sjJyڵ��3b4�k��8��t�d�!]�71���6��p�m%�wz݄�p��)�u,])R�)�.}��_}�7����_f�Λ�9T��<����N��a��0n�'��?��Tm8*�:W��V�M�R��7��y��*�Ԕ�W�#O:x��wk�P�R�����ލ�j�8[M��k�����&���5�U?�����P`.�����t]D���)<����_F̩�81��]K��%VL�)y�jͅ��B���~��L��垠C �S������lI�ԧ�65�x�{�Lc-��,��'T���=����r��q��e���4�֤��p�ڇl�!O�)P�11��t�ĝF��J�iS��.{�"�>9���ɾ�At3��\u#�(�,���X��k��I6�u�Az�orsytje�7�5�4�|��v�|�b���Se���wK�,̑�1��T�{�D�=����v�䚵]=]tа+O{�8*p��!��*�h��=\(�Y}��i�v�_�?P��`1�/��Nx٨7m"-�����W�TS�T�R�6�YJ[��R[`�IGMnmiX�r��T�+����R��
�:���s:K�H֎rP\HW
�\�����lOO)�5��f���֯%fS�{&w[�e/ӭ�0�S�!q�ۦ���ϛ������n�x��4�l�p��6�^sʨ��7>�|�ᘪ&���!f�P��,.B�8n��m8N�d�i�����^�o�������ɥwNܾ܊��+�&��7�{䭾|�L�c"^��o6����Vr�5����7��W�k���tۓ������G4ؿ�7��v�=���s:j՜�݅���=k��7,,�<�2�Vz�A_.�m�Ws���E�^��̗������Fd��e����#�Hf��*$����3���^���Tn&�ji��:c�(!�W�{���E�m�rc6�`
,7�I�}�tme�p��8[O;)ZU���wϤ���B4F�c��@��?4two��+�Y<��{������T����^��C���WZ�Ml�"S�[Ac)�/qzC� �>�A��v+�c&Z-��U��Jq�2�3�������������0bTIs�m���ۺ��E�Yݎ�j0uj�ؑ�x����������-LԔ�v\�aZjihH[�-��6���S�7xZ� �/d2�tE27�)�n�}<���G���s�u�Ұ�U��*!�v��*��4c �\��Ӯ.H/녲4��N�{�����+Sj�7��6��ڶ��$�K^���#yY�y�����/a�h�=)4g����:�f����Si��N�N`֎T��r �h��P�=�|�}-���N��`RW)╮����&�icSQ	��#3쉈��+rv}�-YG+fb�m�?yK�1Ur��b���떸sO�8o*���:~����.Iӓ�q>�c���]������\|\�-����f��ѓ0ˌ��.�F����,��g�`f
�Ȓ���Q1m;S-����n���0�kc���j�[������G�|;cV���L[s�C;�/����{�l����H�������W�~�b(���Cѽ{������Yt�|&��=<
�%�9`�PW/8��g��� w�G��</�LKVͼ����Q��	�j�Wlp�ڭ���皋�{ǽYG�vv�m���(!��C�x	�K`���)3��j���[��s�������=���V����wj(�:���?OM�m���w��rP�y���%�q����u��[w���RS�Kv�����Z{q��u�g��ٖ3l#:r��<��U��M����Gy<��T[���-�6�
{2t;j�{nl��)��Lqs	8��F�8{��:-颓ˎX�k�·��zyn){:Z9�*�$'�}�`�-9�C5}��7��[Z�7/;��C	�x���J3��GH<m����������FÙR��_���]���x���sy��\3hSoa�9U�j�dc�=�����Ǭ�P�i��!�2�l�B|�|�/��*��Cg�\���ۍ�P�S�� �1q���\�[.Vn��ܷS}�}S\����/l�K�/�CT+5S7q����e�����~��A��r�҇f�������6�kw%�n�DH�ْw�(�[�^�컽2ۓ���/���.2���g�x���40��Nxi�hҶzpuft�[2[���v�|�+o	�&c�u-ͥ���[��wj��ڵ���j���ռ��g{����^������Pdε׏v��D�t�5B����z;yVb?U�CY;�w�%<Wwr�ֵ��i��Bӧ��7���dAy����<omPo��oب^�&�j���u���}jl$�Fz�]~�M�t݉�*��G�P�*-[�g��c~�z�_=xi��4�L$���M������|�=������w�	��\�h�=:��w8=p��
��-�i����V��,鈽��y�y�R6�� ��7؞r����Jڍ��Q�+�ب�e�&�_��	���rP=���r{�MӀ&�����Hg�l������W�oz�s���=�v|9{6�fd�;1y&���T$-@n�ai.�t]Kzh���#���]��͎S>�g���w���1�d� Pߞ��#���<���y܀
���c��c���}�s��m;�n7�m��r��}�����LfC�h���Q���ޠ�K��$���uM[M��a�/����W8�.b�o�L�Jq�j�Ȼ���v�ZS��.&Fo���zܭ@�m	��|#J����Db!K���BV��yX^u�b{Ί�ՅfNE�z4uصQ 0��r��$B��f�D�,r��C�v�J0�ki�ɐn^o�a��E�h����kU�9Bu����0��]��3�[>;A�CtS���ILj��[̶�dk�}���X� 7��=֧gݏq�Sĉ�����j��X!e����	]���}�zľO*f�f֖m@]\�%>�:�R���Pբ�m�]7w�{��}9@w���Rqv�	5���uD��P��+6'M��wfS�rɬX�v���[�|Zj1:U�IΗ����ΰ����5^d��.��8�L����f�\*�wiBB�;�a�����4���g���B��n�\�;9j�3�]�E��x�|�*�+�o�GRrغ�H�^�t�q$�V9"(b���f=
5F����<ky2�Y`B��{L=]k����Mбn�^���tδ�.�̥�[�D�T䭴Z�X���9C=4�%��]��e�������M�:��Y��y^:���H���(�9�w���(�-hP��o�X�>:��}+�t�F\�ή2 �sM�F�tAIAn� ([�[{]�QT�xu�4&e����
b%c�q!f��\��Kg��N�x(���t�����>��W�c�ET��uJ�lI��@3*c��W�l��52�J����ŢCR��y��i����]N��37{&��@��p:�� �Ӳq>v�Ӏ�dd��¹`�SyY�<��8��ʭ�+�5��<��f<�q�@4�ZRP�5���(���Zó��ӛ.��Y����q`���S��4VWpRH��x����'`̳'��dP��$�U�˷wt��t34�����˶!�"���G'���ݼ�9����Y�J�����ȇK�=yX,'5�B�ӌ^o2h6�Ҋ:rb�uɜy��/V�t ��f�5wV�V��P��;:���i���yG��_gעVS�t�9M�xk�����ˮ�9�W8�9�I���Q�),��+��6�wwg��w9b�甋����B�K2�ڔ�k��"K�^p��!�W��w�*�͍���_�l�fس4SBq�2���@{����ΧO"�g�W�V�y0���N��:%�P�3� )M��X^�l.�H��2m������u��+����{�@ɹ�/<ź��,�_��1�bw½2�i��a�ʸA7C�;V�|[�B,r�s��s���t�޽�4c*�����u1yE`�f�,cQ�e)x9H��T�g"}�w��ݜ����.�JIyk:��Wk�¶k��c�08rwo��p��7W퐛����wV�Ku��s�yZ�ɚ���ܢ��|���k���ڵe���.��-u�y%.���g�I����j�
�Oƅ
�����v��]�7u�79��H���������Թ�wsE&R;u�n[��s��.�ws�s�˖3r뻜���$����.� ����+�F��]r�+�������G.�L$��Ye�]�.BCF�u���r��wn����t�v�u˝�)����st�뻔����"����8���.�˜.`bA�F"�s��i�@nni��u&�!JAB���wBaL�vD��BQ˖s�-�ƹE]�N��#&ň77(�w6�L"�3&��$��.QRFL����+�\�1���&�79ݸ�F9�,�7s�� Y ��Ѯr.dL@�Ls�y������E���q�B�!��H���n�Q��.s�3�O�WV����w��r��^^��.�j
�o�:\#��JT��A\�r�]��u�.��Ҹ�,�������ʂ�|�A�l�C]p�~Ez^;�m.��>9���o�����D�ʣ�cT�Y;9�->�̡�/T�ۛ�kS-��ߣ�a7�9�(Μ�ac��.�0���9�f���2�'9�^nLFs�p���������G�BԳ��i�%{��?[������۫"�7��c��8��o����o�}k\9��C9���B���T3��&W_*���#-��}��B��Ύ��Je����C���r�tU�{�jl֚�mG�D"��s��x��[��z�U�G)�l�{��j5��eYˌù��]0��Wl�jb����fd�j�����__&*9���齹]���y1�rU�np˄�
q[e�R��A��dm(QXf����"�xn��yW�)��:�r�7��,V�[�,���v���E��CM@�aEl$h;��ũ�ѬL-������0�_�^�����]�8&S�z��[��jk�<��t�إ�H��C;��gLZ7/䃌Z�=���(�ːU�2GӜVq���v�q��ˈ�d��~�	�ek�1j�@�>�.������[�Po��(k/���F�0�US�4:���$�צ����N�Y%�S��Q�-�I���p��c��:��P(w|� �r�ќ�7��������Q�+����q)��*{�8ͨ��T9S
���y�x�xm$jո|������cGuo�sk9�\Ҹ�_��
��ܘ?k�w77Eи������9���4[7����-iʈ�ڰ��.Z[ք0���UD�����ig'�y�����]�q��F�ztf9N�zOT�Y��+v\Bz��e�;�r& w�H<���V�\��R��ۭ{w)J�Q�Ga�q�u�j��cSPۍh�dOѱ�nT}
�mc`4�����n�Hv[���{��g\ru�\9�hm7�Vz��>�G�p'�D|� �v�{��k�,�X�c�$�D�m�mm�&n��dA(�ڮ���H�#�%���Ybx�ř�֕J��vQ뒕�Y�v����jk�>چ�>�x%K{�ā2e�X��):���1�����8yM�{��̾��qk�("Z��7)��g��w�Ny�|��1�O�y��sY���<�b�&�2��a-K����z_q	�v�>���������
e�p���팃TjDM�4�>��E2o�f�x6��ν�-�V}�C+5�oB�UsZ��nyt���%��Wz>��&k��h��}p�f�؊.�X�!�Y�9�3g2�6�J��K��M�-�jƴvK���Ĭb��a@%�t����=�����J�Ku᫴�눖���jʦm�9v��V���j��
z����}��D�l�I��~^�C��ƫ�qh�6�Cw(��_̦�����9�r��A�.{��:�zj ����G�R�r����[�jL0�������r��sҲ���<�Ȭ����5��@o�t�*��Ub���p�Nr$�c�����n��׬��B���A�D�-{n�-�8���Þ�i��:�	�"Yܢ:�����*Y�ŕ2���m��X�����9��s��[�����y�'�k��kH���{}8�Lm���Co:cZ RK"�V���۝��ޛP�i�����&R��S��x��tmd
[�{�c3ZsQ��<�N��B�{٘Dl�=�0��ו���6{��`o;(g����I�>9Ϝ�o���x�ȘT�� �b/F��f=�V�R��.bj���[Q���gys_&�]�s���0��AF {�Fg�k������C����7W�jڍUj�I�D,p���t��uy��{�6�����=�eؾ�9���Ş��Jyvo�Y��<�oYɴ1�g{��7+����%͖�	[�K�[�*�G7ԕ�{�p"kb�k��O{3��:'Jk3�K��p��Y7�	����Ъ�cR�B͎��j���c"^��mo_ݛr.�Py_xi	��iW,~��Ѿ�����Z�z�߰��	��r����7�p�eW��OP懱�}��Lc�Mxr�	��٤}P�؝+�0�*>�e�m�ľz�(��Ex1Z���沐�M�)	7�no��^���E�j�H�D�D������Ӝ��B���Y-#�U;�z�tH��M��OU�@�u̷y}��.���֮u��L�oM&u�g�s%3Pve�����F��w��Y�ێ�����Lz2�Xf܄�V��v�ʷ`l�$3����w��QY�+|�@�s���j�,�/F�jf���r�IP`>U�Ԥ�I}������rf$	V�{�j{�лc����9JR��A�?��J\���Es�Q$���d�¦������ې�ͨ��S�f
{�����ṹ˦!�h}mhS�?��y��b�ނ�Wޥ��
��v��3�faء]�*�e6Ķ�)r21���s_D���_c�������㕊���X´�x/�=[!�'���43a�kn/`1�i�^�����������"�^걞����.N��JS��N��?r0
��ܳ|�#5n�lO+r:�%��[X��i��mƻF�=��P}��G��$��eCv����bR��)�w��x�ڧ<^�^�a��"�E����6�m7�Ϸ���$�m�	�]�7��BXW�&�ߺz�hZB<�kؕڬ9^�+q3���uÈ0V1#(!V�X5y)�,7���h����l�d����ع����1�M��$�޻�p��B��)��ιL;��jK�ޡ��L�����b����
��<�m�Q�I�)��8�]�{6�#u�fVjw�'Ub�q6iUOg�fS|l�@��;\v[�p�y�/����S3�]�ӞsVU��]���r�t%os&�ł�e?�r���>�*&/�f�&źoK����L������1�����-�Bn}aC��Q�&��
���]�jF�㕶�h��O�n=���ѫ>��vK���*Â���FP��==�'��YU�o:�.m6[��1�Yq���i����:y�E�]T2hJ1y[��[j���'ѩ{o\5�]�׹ţd?Y���N����z���u�9��1i���-�}���e�,q��r5����I��a�dv�����$���ִV�k3�w�#�-�p�܆�D�{��z�s���ⶆw8x���{5���#��M!E�AP��X�]�0���@C	��;�L�8��;��r��n+$uD�Q6
zN9P����99O32vޅV��s��wI5in�Z���Y4u`7�"}ŗ U�(,*ӂԝ�l��!�e˺����үT�6�
K��C{թ���
��I�ܼ��5Y�<���1��φ����.ڽ��scfL��g�����.�8�ۚ��2���W_��]�C]�{%�T�rXR�^�ھ�$�h�秼�1T�᧍���k�Fu��j0/��^!}��闇|/J�'�.9�L�Q)��x��p歡���k��)�����H�y�j��(����͍�ꕧE�����Gu1�ڬ�yd>����z�y��6��T=aF^TḄx��c��;��e{��.�ȍV���~��̤ ��.�ﯯL���gᚶ&�j­>&@k��}�������P� ?Ll�D��r={Z�-lm&G�U)�.�1l�6��y��q�rO]ωCo闄�Y�k�#�O���3�u���*X}�)G�|=z}^%2�}���z��7�#�hp�:6ܒz�P��.^�eX9�:ww�R���1�����<���9�/
����ȯ;�v�4�a�} l=�y�
<�-��M��2U�;��u<��f�ǅY�Pa���jE�����]p8���e��:-�՜�qY,d�[����%��u�lq��%N�*��v�U�ظ�B�ެ��=�r�XZێ�Ș֒�"Y�'��.���W������{��X��x�̩f[�����w������=q�;�u]���Z_d��/+�|���_�\�5ǉ.��~"EF̤�!z�'��{��Eķ�џ/my��G���"d�9���&���k�s�'M¯T;�rY�D@�3���o�W��&5���o����O�.����yؽ\+7�x�+�����oޒ7��%�\�Ȁ���H����lt�}�Q���q�]]�^�Q���>�?���?[g�8��`�kA�{נ_ޜ�I-�ԶG��{.��U���|����
�:�<;~}�Fc��G���O�����h�$d"�K���O���a�7!{7��'<:��6�i�	S�|�R=q����/��7������|�q�Q�X䱿��t����D���p��*���D�m���^�{�ƨ�wx�o�t.���-B����ϝ��>���<�5������#���CW�^t�!�R�||�+��}���:9�W�����n���wݥ�!�F��7��ՋY�"�''�n;�G2C�M��h�xN���^��I�b��`-�����L��*u7�U�j��9x骛gU@v�"�TJ�	�貊n�i� �Y��9Y"y�#h�����S叮�8og�Q�-���O���s`���9k)	�oA �W����=��n�+'AΚ�5�'J�C�lvYتt�IdmȺ+3�9T�{����~���y�sS���\k١����o����ߡT^)&�ōxZ�=��ކ�k����>�*g�Oٕ��ǜ�~>%�zy����*�5��3�פ�܄���M(vzT�{*���s>��&x;�Tt\T�S���K�k��|z��=�SW��Q��7g���o�Z��;x�?-?Q�w�.*���	K�5�A���A��>�.1ǩ�����w�M��N� �y̕3�*�s�S���O��$����U�%�!x{Հ{o�����u�k�ힶ�b�ۥ���]?[���;�)3Œz@(1���m)l�yw�9`�:��V�~+ij�U�=�O�oN}�H��� �ߵT����0�%T) yIׁ.����J R�ja��(Y�uE�r�ϩ�\M�>��C7⴯��:z�=�#|e�؇2* E_����TN�$��Ct���^΃�ϼX݆g��֩�/�ف��l�L�_}��%�P��/�a"e����?#�G�S�u?ImM�N��o�χ�7��u�/+�`{ʏ���2_����~�G�� ��OQKq�6����w*�p�`�Y��!�Z1h��£�\�]���b eO1
�ڞe1M�뾾Y6�j��$//M��	��N��)Fșy��x�����-ڦx����<B���ԓI������3s�^�a���,��"8z1���R��ya*���)������o����r<.=�wB�}�а��{:W_�Dﴞ�3<��n4��z����TT��ӟV����޸|zڞ�y7b�S����z�.��9��+�����8�!���aO���������f�0~"�J�
c�aþ�J��f����onB~�E��Qy�;y�X��f��x�9,*�G��;U珌^)������pۊ�\O��_ݶ�=����3�?E/�޻��������ٜ?�EE��|UEG����Y����(*�::�r��.|Nb���,���?g�؊�s+=걼���{�hz������f����~�1us>?�d�٘�P�"��VMi��@yg�i�Q������
���ʱoh�@�Gw}Ī2ޛ�:c����!jڞ7|JVf��T;�U#}n�o#�P�;���y��f����z�o�G2��w,>�\�D�p��R6��x�I^4eT9��P�c��*��:�=�uV�&�n���>�iϷ�<^����S��^�9\�6J�R�'�&X���
0}GM�y��n�f�;����S0	}:~nW���.zX�w����%y�%��x鮆*�� [�>r���8ma�g�C�\�7b�2Z�8&���$b,�ٝ:�;2�g�p��RX�Q���y��*�9g;1��J��b�.��g�خ%5�.V�nN�K�n�*�Ab��+XĔ�c���>Ck���(�7�Y�V��E۱3T���X�q�h)M�pDK�����b��97ڬ�A��2�K]�NH,�$�وJ\�T�:�_7i\�;�gwuC����kD|\r���kzXJ���� �3w�q<�ʚ�v�i!O�iN'¯suQ�o/��Ǟ��L�Ư#�߷/i�Hz��o��N�T�f�#�sWv\pGR�(\}�z�O��W(2D�D����w�2^������,���#qA�j+{HNtM �m�-�KG\�+`�yϫ&�<2���r�F�tDܣq>��ʹ��ͦ�uJ7x*�Gd\��V�\��"�0r�tˬb��W'��k�s���!Y����/m�^�F�k�]E�b�\�'�7 [:f��ȉpo���F�4^�ݘ�R�t�]Kdq�r�6�}� U,x^w���:҃9d�Uq�n��� c����;�X=�l�Z�חzv�j��B�/�f��U�q�wR��mF:G'n�|��^rG�EN:h���۔rӧ�HlJ@��1�5�&Kc+6�4���t�V^j�i�竛�ՁJ����v�W��c�%]����w�:�m��\�a�@��
���╧��@WU���2��Wus4
�3^�\��:~|���k$�v�չ�@�,�*�m��5�13�CхV���j^L͚4j}�rt�7���m�w�`e�k���g�l����i����VJ&l���ɻ��2�V.��v�3A�rѼ��Ev�fy���߱�Aԕ_:o!��Q]Δ�u#Ʋ�7���v�[r��4,�}�O�l��� ��ꆞ��n�IR�/�=aj4���kR��Ҿ�Ev`A�4n��}�c�ܷغ�eb4�<srI��:*��[HV	-P���"^�8x]k
��4.�2���t�y��ˎ]n`����%wwl�ƵF�ɔ��7.�Vswc�㸑���=�Z.��6�.���fCe:���ťe�ò�5:/�,�V:�<y]�O��r_T�X��,[g����M������ٺ����c݁Tܶ��JM�|���N�;������W�'r|9]�*�H��+v��pVMW@���b��.��_T]XJU�:9�.w�NZq�6uj},FsZ�'v[��ܸz�=1S�I�kz5�¶�Z$�;j��(�lf}�ȧ�8��u���O'��7�b1l��ѕ*��d�[�� `��s#C:��y̖TNp�d��:��j�#܂R�����d���]s��gC(�Իc"���6�e����o�Y�T�%�9s�A%%T�+}� ���T��KL{]Y�7�U  ��*��(�B�D'8���"d��C1��$F#Q�k����wn��LS#1����k�q�.�rL���JdC(�[�4d:��h�4���wvwt�P2Q�7J�2)�Ahر$�cF�9��Ԗ5�Y��d��'N� �AI&���dт,d(�,��26�Eӗn�B�,)��"$4ɛ�����FfGN�,j.�@Qw]BF��6�(��r�Gw7@�B��;�JCl�$�5�k���VJlP�r�h��t�3��;�s�#wrE�!�lX��b�%��I���+�$L�n\�4�ܗwR��k��1n��1�A&�)�*Lh�ە�E�TF��HDIA���t��U
� ��1���ve9��S��ي�`�u�L-�+�RXҷ77Xެ[�J�&R�L���]��%�MGv�1��5�.�6'�N���8iw�/�~���R��ubo��q���|C;�ꅬ�2� ��]+�d��K�[c���� �GO�g�l��]w�W�HM��ֆ��=��v;�4��pw���7z�_��9�� ��_�'ƣ��ޣ �H��^s��q�ւ�;c�iƚ߭��Ԡ���F��u��Z�~���U�`�s�D��12�]F�Z>�f�]��d�li#c~jϧ�Y���٠�� �Y/�3��~������w�3�]B
��F���MO'�kd'��K�3��v9pю6ϡ�ƣo��~�p��@�<k��3ZD;�&Qd��2�l������Q\���s	{�z!�o����7��q�y�QOex�>���j�q�L�0�L�#Z}^�v�R7+�{����N���E�Z��/#���w��Uq���^�q�p\{׶M��oL_�������}Re�G�%T�򸁵���O��T���=q�w���,�}���}J%���9���'R�d{��}��X�yS����ۃ0�@��ⲽ�K�1S e�W�D�����ɺ�v!al-{!.�W�:���j���k��`Oc��B֕^�B{~���5ٯ%�WK�|ɩ���:c���F�j�2E�=�,�o_N#�5]��8r���7\���"�K�K+o�u(�����[¥�ف�����n$s�=`�Ɍ���/��q��R��T��R�ݳ0��*�qYU�I~%I��&6��K|��P�y���Srr�j�ϡ�H,��.5N���(m���_A��W���vmH��x��N�ya�+���r:e�w���n�����ǼT�Tf�+�Μ���$�Z��y��ѹ��ol��f~۔��E��B}:�4�>�y�/K���:��ߊ�&�шF���/���3y�o��H�?E��}_@L�b�R�Ws,�Subo��ÆGz=LnF��=>��:�����tR�d���U��xñr|iU`@H����B��O�+��."[��V;<�#�NN�f����z�y �}�A��F^!n�C�%��D*3�뉾�^/u��Ek̪��%��޺�앶����'���y��^G�ޮM�{�G\z���2\�Ȁ���"~�끉yz�[��٫}��a�^^f�|n5�Q���/���>�����`7�-̒Ѹ5-��
�N&s"�k{�S ��
�m&xv�K��#1����n�ȟ�L��3Z4��"j[�'�[X*�u�S�(c�����}�i��/* ]���p��#�G���՗Z�.:TVD��sg�u���Ta<9��^,Ē��O,lB2�̨S�e�ڹ���ZI����2v�%�K'�w����AlHv�hh�i&�^��ڀ��2���v}f<�M���Л���p�>7�R=�*�0��>~�@�mk�S7��X��R7����\�&�E��&\	xb���������\��0ߪ����/xQ�� �]ڨ�'<:��� ���,\w��>%hɇ�'t¿�պn��尕�p�F�l>�x��]{he[C�?Uy�ޡ�K>�^���j»�����8���v��VW�i3�˳ws�:�o[�v�zt�<�3�J�S2���5t����{�.!\䜾������o�d���$��^�����uV����(�>�ؼ�=�&W�'"����������o&tQ]%Ҭ�GX��)�}�KS�ӿ�.D%���Tt\T����,�ׁ�/S��>����j�pzțv=�>�j�hū�g�gĥfX��3�o�A����a��}^_������F1u�Un϶WqY�Z�i�� U����I��WK�
︺��_5���������l4�Z�~�Po��(-�o���1�*''���\�Pd��a��>U�i��\�o�s�ܞUxaY��6ɉ�0�8�B�m>��`۵짥v��J>��B�qAu���AVsd�M!���Eg.��!B�%v���$�͕v�����%֧]�j]� �p�:�a���!�l�>o.Y0L�	]�bTA���E�IGO_%ErR{�W�l��������~Ӌ�<�7��q�U#m�0� %R����%������c��V��{A@�/���r9�?+����"��G�'O\g�dm��f��,�>�0�����`|��K�
S�x2�8fy�j�E��0={Izgt�{���Ͻ~�'��;�C��G�fO��l�'�)��)�����z���u��2�����h�{lV��/�F9�}�Ϊ���W	����AH�GkА�z����U�ثF����;��}^��
���e��|��P���L�g���C7�ԃ�Y=@�|n(�����Y�U,��u�m�Qf�ߨ�x6�j֏==�Ѷ}?{m���]�{�տ_�������ڐiO�T����S�s`W��y�r��,���)���;���%>��YP��WC�P�����yt4<����E���z��M�����=4�?@���YLl�����_��۸�:���?E/�޻�����?�:1l�W����hϹQ�ɔ}����L�U����9'F�U�w"5Ss���̯[\�=Wd�k����{s��J�vt�<�Ct��@�����a�"-���A}L��մ�l:u)Ը�Ns�P���@]>�fj�YŔ���Ƿ s�ԓ2�(k&-�c�Y����ovPĖһ�<�Gl�����Ηeb�4�u��m���5��F�]� 5��&�v��W�1�s:vd���.�kM�K�<�4����#|��'i���p�f������AK��\w���?u!z�����)\����C��U#����l�"�SC��wعU������Fx��_��<�+և�dD�p��R6��x�I^5UCծ��\�=y�9%��]S��>�s�'�S�����8�eg���:�윮
��T��Od�u*�e����1]++�\�|���Q�Krº�񔦄�U�>���>�Hg�ڮa�e�=^C{6�3�܌�
>��uP�f㌶X�}u�9�W�HMϽhh������=3K�5{z"�7xg��1Y�7ﲫ���ʀZd��E�L�9����Ç�}�lzlW��3��z��7��"M�F���o羸�7��D�2Y�@���E.�vMzu>?ndc�N���3�x�U�$�Td�Eۤ<}�D�>����\���g�*��Č���&D'ꪐfH]��޹�o0��<������m_��?z�>�� 7��5�S�rf������[�C
�Կ&���4�r��"�����#A����=+�+�a�:]&G2v!�w��ݬ G��ީ�WW�.b�,ӳ,f�Fs�Ŭ���p���R�{Ae�"'X�눊�����}ˤ���9�����J7DV�bf�M])gs��7(H�br�9��Z*�)���J_�������������@w��=s'p�9� ���F�|���v}rpu����V��V����|n9��<o�h��D���=.��=��L��؍ػ�w�h��8m�J��F·'�pu9�u���ǯ��G�s�7w-���Rf��FΏv�BQ��Jh�u�Q^�U���̠P�гj��z:�w5[ KOeW^t
��=亲��^c��_3;Լ^|�V;�}�.6�X����^d~�u(����FJn��ŧ��C=8Oz� +=�dZ�M�u1�g�t��^�B�N�눹�(m��í����}���&����5~���`׹�����z}^&ӗ��ؿ\{�ey\og��B��$����|�nItF;��U��*W�<N���Jb�З:�4�>�q���������^w�F�O��;�g�\����aXe�� �|e� �X��K�!fT�q�X�����w�����v�Z`K$��{�J�X�^�;��g<aع(��J�,	�R$V̤�!z�'�^�;�J����ߗ�w=��)Ze
j=�(8����z�L�y���9qVgr-glkE>.p�Uz㰂mR殞��tU[��u�a�ۺW ���Ru[���(o�Z���;�l*��=N�m����l(���.L�G�M*���y�94����ڮ`$���^-�2	ׅ5�ē�Y����xE��m��R�˘}�H�Ua���q7�+��x��38�0����9R��&�mTO�_� ϑ��p�sޒ7�,J$�p��������8�G�MG�ֽ�L�耥��bc��cZ~��Nq����փq�z��=9�,�Z/s���TU�歡=��^�dzt��"b_W�J�#�a㏌�z�����>D��s��>f�x��,�������*;��q#��R	�����>��u��Ȅ��~������߬����T}���s������f�b�5u�L�d�Š��}dH	�VBƾ�]��c�9��b�9�0��%4��yb�w]܎�����\/f����Ĩ���]^��j����u��#ٺr�uU�<��?^߆|�U�rz��,�^���j»�����gv��w�=��Fۏ-�\;��IxN}�|�m:�N����y�sS����k��j�$�멇Kk-����F��=�ϩ�|zp;�ʭ7S>D��3���<�L�N}N|�����,^�F�����|njb�N�I�M�ʫ��4Cy�>��N���F)nVJy�E�����IP�=-�r6U^�)F�����*�0!�Z���隫�g^
W��H�*�{b�z�FU�*d��_v�$�%�w6KV�_WP�Z��,s��n	��:����P��<�Q\�#OH�9c��g_��~��y_	��*]R�yN��KK��/������c2�������t�[�s=��j����B���S��AZ\P���}n�/8��<�>�2[�ULT3�}9��f�����{�^�=�s�R�F����K*e#qwQ*���(�r)��v�V������^���O����D{�Ǹ���W�P�$�3�*����VǠڛW���{z�{ˎ�]����TOKw�8�#�{7��q�U#m�0��l�J@R��gh����q���e�=�\��ϟU�F}�>�w���['�tF{�L�ڏL��'0���j�s����} ɸO�=�\��ưu�R>��l���6|N�}�[�2<M]������^P��7ﲫL�$���DĞfED�g!G���m��[)��苆�w�x�B˻Qޥr'3�9��[�,FyӐ�qM�Hw�-�'���Fp��}ʘ�Vͻmx����S��UnF��U/:�>���b� ����2v`�zh�D�=�ÕP.!����)���#���0[�Ե"#!W���C+`����ӫ�I~0��4e���̾f����o�ٍ�������U�=�u5m)έ�P!�cY[��͝Ɠ�v�${������m�mhӹ���F�g"cn�&����T�*��(��[�z;�-9ܯP�z�����w�~���{o��sTS�P���d3�b㽵 ��|J��Yt^G�[�~���+���~�E�����ā}&y�kV׺{�h��P�q����{�8<��ݲ�ӛ�ªN��8�������^�c/�JR*}���/��m��d:�����R�}�=�<������3����%�~�?�5��@����W����j���ک�Q��Ꭹ�<�tw��x��vd\w���g���;i��k��oC`�Wa�	�,]d֛�t��`e1�!��{Թk͍�6d{�o���]{ǲ)���Y.R��Z?&���1���G�0E��z�1�����e���t�a�K�x�W��"��)���W��}^�<8���]�#n"�x��W��D�>�)M��k{�R�7�Q�F�ϠK7����>�i�������S�W�xv}9\�d�+�0�����𝹺��<T�	=艞G:�u2��+��z��|���}ޑ���o�3��^gt4$(�5���J�~�_�ѿ���F���'�x��l��>����	Q>����[E^^��vM�]���-�����
���`s�uv���a�|p�'Û[�����ś��f+I�NX���P,�O��{5�H_utW�j೙�D�r&`;�c��tɂ�]S�K�\K��7�����ʮm�-��n�jR��:���G;�����or�|�D$�ڪ�K9
	W�@?x��G��3�\k����b�&p�L�*�b�p��!������w��BÿO��QfG�:H����4'S�������"x�^��;��׼��8\'�lzQ>~3��q�z���뉨�3�p����"��o��F>�4ȼû��T�^�>�s�z��{���f�[U�*�HxO��ցP�R��=��ǲ&%x{$-�Q�
O�8+��9-���K���Q�yUQ��^&��ޠ;��n�ny�>��t���꩓�Szh���u+N��}~����;ۇ���ȇފ�(��1#K=>��3�>�k��l�+L�>%W�2a�Z�O��n���<��G��u�~����,��z#����w�����p�*p�!��S�HW������/ʷn��3[B���]!��mSe֣)�2��V;�w�����b,��a���P��i\�?>Ŕ2���ء��?�i~�fi� �^vE©M��wQ��t�ϗ�п�N����ġ��F�w2 (���^*��PP�bnvh��N�����X�]�g'i�U}�h��i�ӷ�8�[��Piu_TJ0�W`� ��pa.�����T���1�����ۛ'��BZ����b��+Bqm�0���za���]vLW��f�/�ܸ���mݮ)�u�-Iѻ�� ż���,����X���Γ�s[社\xaM�X����E��[��b���*�N  �i�X�����܏ (v�����s-]�v�\1q�q� SR)dʌm�L�FD,��uW-�c;vY锜8�cm�pա�ܧc !*V��7)���H�\��Lw9O�XM���AJ��b��GĜ����;0�E�'a(^��J����sS�Y� �;��˽�c7A0��ѦNZ�qq݄!O�Q��@^�`��'�.�қ6����B%^2�vHsn��[r')��N�����
��V��gDB�7��n��n�+�F�#�J4���B�0XT�1eR�dR�F���囨�neGPV���tvИ�*���;�oE-��M��<��%o�)&�-8h\�u�M�	�ْ��=�.��1J����!�ovb3�biE3gp�t�;.F�P��s�k$�[��5�R�e>�zU�
�u�l�T�8ӈ�QQ��F��E���e������u�6O+JkI*/o�h}Drm�t�}%���Q0�Ԯ���E^lY�ͽ=����kl��ǫii"��%Ci�BK�ç�'.�1R*����BQ;chs�;yM'h�����`ݮå&���, r�;Je��b��/5�>MA�XY����Ǥv�{����7E�#X|���������
�d���ȴ��%Ԅ�kd�w��)��8��D�i����q�x�v ���g3�u{��ы���(>(�y�Ζ��[g�l17&��llE�gH��C�,�Cd��i�Z�B�J�c�����Wu6���t�R����l���㕼��u�*���H����J���{�\��4���0N�[����	�&lV���WTk�K�ۈ�7x��
5�:�A��f�`$��4a�T=B��bO)�K]��w��Ar�2��/(ƶ�=��T��x���upe�6� 9Y��Z9Sr-2��i�!�� �>���e�K2�|z�[@����#%��\��vEA�gRnU�;Q������d��hm��on���*�o;Y�.�μٍs}��p���(�q�
�q���ڟH�x�;�.e�fVu�]W��� S�B��K���Գצ�uS��;���x��ێ��i��C.��c�i�}C��וqk�]N�,�ѕ����	�W�/��LPe�Aaq]�fN��9W�Pl�Sg`��1�WVbB��#�oS�w,i�,��+#˧kP�x|�]e�-\�Z|:�Jb�+��6v�K����/&N׭��gfwe� j��
$��c �n\�f9٘�4Bk��7v���wBd�Ј��Np��"9�	S�t��q�[�0�3d�۔�QP��Ōbv���c �C+��昒`��)$�.ca3-��w[�-�;����1ʻ4F�v�g+�"�� ]��N����rwY"�B�Cn�c	.r,"#0,��7h����$Ys� �N�	0��Ȁ��%wn��.�\�������gwwQ�ؓI�B9rI1BGu̢��l $Pc�,&��d
0X��\��;��iKL�s��Ɛ9ۺ���ۻrwn�%˳�HᨰEGwF��Q���4A�&�����wlw]Di��A�ˎ�b.m�\�a]}uWW@��5�#ـշJԫ�,�R�7 �j��zC#�YɺnN���>::�^R*t��[�0:����<h���#na}9��|?��C^�U\o�P<�tϠ;���7	���m���*|�3z=�������5�uw;^��&�Gc�Z�?HIØKa�~�0m9���_�����+=C������P�
:���w9�Nu�iO�k��;e|hSF�)�?�X��K�eK7MՉ����n�w��^Bv��m�y�9u5P��s��.J5���`@H���))�^�����dmG�!Ϯ��o:싟! ������+�#�����t�Q,�"�A�ps����ёՙ�s˲�Ӌ��w��򸛟yb��_G�\8������U14�K� �5��4�P���⛍�]�=�=>��nϼ^�5��F��?[g�8��O���{נ\zs�N�jg�]_�ohhV���B[��^D�?�^�BFO�!WJ�<;~
_������~��|��~���;q��u��yN٥�D��:�Y#ȳ�Ff=�X*%�xи�t��%O��?T�{ʪ�fx��ՙ
N����J�H��)����F�Y�Pd��}b}�*Z�џV����c��x����� �n�@�Z�M��k5Y�]aٷ��m�'�mCQ��f�÷�#Kn���$J��`��)�	v/�?sC�V ��b�����9�FKQ�W�]�"�94�c�7y��o��OM�뽆�����sjݷ���:�����u�t��a��^�6�9ʦ�y��ֲvK��֯�Oz��Hu>�`��٢������*�L>��aw�^��Ȕ~��
�x�*U,-ټ�C����oo���8��<ido��o�V�ȼ�d���gz�rn�|헾���C�R��qS+IӨ����!��i2�yV��V��:��4:�r�2U��D7"��b�o3_ag�����EN�����d����./:�(u4�|Nק�Y���v:x�as����˨z�ث�c�''N��,d�I��R�yN��KK�p�O����J~駞�7�{s�M��2�Ϟ��y�wb�F3�gN��>WX�x�u3�o�A����a�}�¯��W���$�wo>������?W�VEz�}�
�#���Y'd��2WK�����k����{���w��w{�*��D����,G����ћ�3���\{�Ǹ�ӓ�\��B,���84R>IO��ԏr���Σ�Ѫ��/�˸�����n%����^��=�o��ڦFtC�a�d����T�V�z�*�߸qs�s�(	��x�-����r9��&��z�!��ZTG�'O_��Y��"_�o�{�`��x�f��B����U-����^�ȱ��o	s�Ҵ�hv�9S��b�2�խn9R����%͇p�'���Eu%�V�D/Z�C��̸_�oB4�Ps�ŋ��sbd}m���M����}c�x¸�h�Be�
�6鬴Ԍ)������Hz���ɐ|z �툟Q-���1C3�޵H,���l�A�u�}q/��J@#ף��J�W*�%�����U^2*�eI�㤎�+�h_ԝ/`�y�o���6=�4��|=w�%�ܾK�A�pC�}�Ϗ��K^5�ۨ��e��0�b{T��Q�-l�V�^pʒ`VָSr�u_���=��u#�����>'��|���*>~ːQd��2���V��~�9=���I��Gx��������y�QO}@:���}��X��ԃP�ĩ��wn��>rWt.
}�#��R��q�/��ԥ��y	��}��o=um{r�\g�˹l����^��r�ꙗ�K9((ӡ�Օ���<{��ܥQ�:����Ox���%r�"�7��N������ߍ��G����g��i��*r���J�����<�<;k���X�WA��v��m���w�2�x��ޫ���aF�T�A���a�"��Y5�K�<���H̥�W����D'�~23��~=u��(n�~�B�mO��R�3=0�{T�~r��ɟ{j�2З3���!y:�5�ѴH�<�� p;�����o�	�	��Ү���UwV|)nZ9٨9z��<��qa�lM��ɛ������f��������[I�ҵAc�O�^��-ퟺ�l�f�����Ӓ^*���;��Ìt�RlC1���?�j7�1T!_�|�����^Y^�<;'+�DtƆ�ּI��~;7�X'����S/nL�/����[#T�6�_�Pv4�?aϷ�<^����S��^�NWW�Z�����7�w)�W���I�(��C�[��eԳt�X�n��w�x�9��C=[�������꼊���S^�����P �Pe�0���-�2!��x�W�HMϽhh��y��]
��f,���dI�n�7#O^?\��0�e( %Q@1��I�+�u��W�"����/tIS4��+ʌ�!`��A�u���=���7�TM3%�D@n�O��WQ����z���^�<��Ë��o�Z�����a���z�_�'c�3�!��L{D�x&_�V^�v'}Z���=}[F�S=y����y����W�7ޤ�#Ƽ �g�ց_;�&n�ܺ��/B���w6�N���r>)V���q>Og"jn_�h��O����{>�����F��P�����gӛqO���{�y�YY2k�1��G'ã��ߪV�Z��/#���w��Uq�~[�u9o�^E�d�z�j���7N�
��&��\����M����k�\ՙ��U�>�վX�J�t�,0�����2_�Pî9��֛�^�ðlY�ٮ'K��Q�|ɰ�4;��WS�p����U��U�{\�q�WϭgI�JШ��9�b��������N������G�L5ckC��iЩ���Ly�GL-�d?XZ�+�c+��?W�C�H�Jqޫ��u�<ʜ7���E�|!fկ���{s7�J�S^̛Տ\ҵ��A�Bw�F�W��|���ԼZ���=��B��eN�0��_��4��#�4x�ؽ<���/�]U��g�J�> v&�U)�8�WN|ۤ|�օ��vOvC#Q6������S�'c~	m�:��K��:��:O�a�~&ץ����q���q��kn�Ne�8ޏj�=	��!�s�|.�I=S(z�L�w3�1��K��������/Mܹd�8ׇx�J�֛�y�.��=�Q��$�2��|�R�x���{�n�N��G�j���^�Z�D�CBP����=~��dA��b�H���`@H��2��!r	Wk�j{,��ݒ�~�{�q/޽��י[ޡ��=���r�Q,�=��8�G�������WwW�hu���̴}�Lj+_�������o��p�sޒ7��LMC�.v}~�)��H���o����T��V.ܴ;���h+���O�V�e$�.��`*��N}t͈IŖf_U.G���]��4/����u�J����PEuM·���e|̝��͏��z9h=�5[q�#b����b�ǉ��#��������F| ��D$L�W������5����O��p}9��:}��߽��0]�1j+��]h����lo�o!��>��'ȉ-�Ď���
��T�����#Q�ʽE|�>D���v�GH�P�8�]t����=(��k@���"���3����Y�X�q���\�R<�\�w��s/"���X8��y��f����{����2J���O��kk�k�q����H��h������ݞ�����U��M�{��\|��,w�d���d���a{\�y��Lx������1��?��q����m��d'U�rz��,�^��&�X�/��w�{Ъ�nnb�j����9��gǺ��%#�3�'Nj��vۿ_W�?�?~�����ߩys�ox��;^��`񷿼ɝ��?����Ӷ��˝�ʭ7�+ģ����<��e���̢�to/m\W��J���{ѷ����i�KE�y;ixc	A���t_�ӡ�9�,q�߁�����L�>��u/v����W����v|�Q��ӿYd�\c(���L��!�F��A�YLI�}����5m�Vj6��5�=SU�� ��}g�Nһ\�
�7ڡ#/2R��v6A����+�I����	ac��W�^�Y�P�������Mm�� p�&%�%��V�G`��K�ك&�+Y|�f����5�T�/�� ��7'ϭ�^\q�=�Hm�X^�}^_���1��^�S�C���KOz�$��J�qz8��>erߢ2�����Q�n����﫞X��Ͻz27�>gr7�����q6x.�rQ�Y%"�o��^EO�.96jG�\�}�]G_�sM��.�|n����W���HO���m��}{��4zG*����S�gĕ��}��{��x�p��r9��&�޴�9��'O>�b}g��n��lV2/ѓ^3NdT �ؗDLKu��/ŌL�#z� ��~��M�q5�ٙWIɏ>ű�VP�~�Q9����q=��K5�a��#$�)�qI���f|=]^����:�{:���v�2}"��z�ȃ�+>9��K������2������=�*_W����aM{#13(.� 9R�컛�y���;��q�+�μO���&n4
���K'����t�� .=y��o��S�G�艵[�t��������^
=�WF�{�տ_���r�w�d�||��f�i}|늗D���g�)V齹||��/����4�U�>��7�z��}�8�F��ti�}kD�h�L���ob�v�VX��+�%v(��u�
�o*���v��ϕAA�RLQF�䡬ϯ������5�S t�s��g�As]���U��q�p�u;��Z�B�=J���4m�}��ǳ��g2y�<zo %E2�wEɭ��P�;���i_����t>���ۊT��9��o��ǳ�S^�Qf�(��ˉ���j�>���qĪ���z����3��'��:�T�iW�wT�5��d�y�g�f1��z#�O��v�\������w�����ӼY9�C���
��n�,ύ�*������Ԇ[��`[t���:`��^��t�q��.#V���R�3��@��C�&}�2vw�B7�����H��~�Ȏ5B�nȼR����W��}^�<;'+��c�\�꺊���ɫn���$���0~Aؒ������cuA�~��߷�<^����S>sṷ�ܣyy���z�E4������OOTD��yS-ς��f[������#����>������V��sw���G��`O�J��-�1��x�{ԄĈ�S�t�&n���Y��W
���|����x�:�޸;z��qD����� ���E���C۾������+�^�?[dK�3���c���'�����z�k�d������&2>�S���E[>%��|�{��^��n����Z%���m.�R7!R����KpgLU$}$s�u�ޮ�Hs�&1�X{��@��
�Sb8��ǆ�Q�c�M�O�<�G�*>���oۣ�J��>V]n�q�L�y[+#���N�4Z��bV��BξZT���G�ԥ��bc�ֲGO����R'��'���p�\)i|�P�ڢ�J	wlykv>_(X~�RA}>��R���z��߼�F�ͫ���ԁ����Lր��iy�=t�ك#;OA8��������<�5�=�����K�q��q�j���{+�ѭ`��1h��Tk��Ui�+��T*Y2k�飒�\NqR��}^������I^����˟T��]���`�z���z\�����3�㏉U&�����>Ӣպ�{9�7^�������UW��V<�^Y����w���u`���l��Xݳ0�P'4���{o�$l�=ޏN�y�J�=� *7��U��g_�x�^��#��RW2/!K'v���]�u�ȳs�oOo�|%���Ss8jR���4׀��-T�亘ų�Cn�Y�h{�E�ױs~�%��h]��{���L�d�_U��p�=]C����<>~&����h6p<�zWV���I�vk��rS�٘��Y#��ȓ%��%���L_�n�����z|8B�;es�8\��Z[{a�*�u�M�U}����p,�>Y�v;219����b�V�T�Vh�j�(��J�y0�䩸h���ʺm�]�n�r��D�oD���p�9 v7F	��\���Ӧv�1A�(<������18�ME.ܕ��v)�:Ϣ�����=�s���+�
h��)�!�.����3�&(w�2�������}޿ޏS��ίy�{��xñrQ�GĔ�H�8B�\��t�
 e5���:�}���N�'���$\��ѐ���WzF_{i	�p��;%�D@�΅.Y�lT��f��eΓ�L�bcQ_}���n}�ay^G�ޮM�Du��&Ϸ�����W���Ư�|����_��;�����h�3Q��kF���6Y��x���.��Nuv��?tfw����϶�~�?}��f�L��28�_��:T�����#Q���Q-=���2ce�[�7�\�y����zKp�#<�LH�Ω)��u`�s�4.���iKә��g����}��9����Eߤo��wF���~.�$X��~�����A�B�Ȕ�+"��8*�q�/F���������c�9��c����:��ޟ z׳E���mH5>%F}~:b���9{�g|�_q��T��\��[	_���꼎D>�Y��x�d�Ws"��ѕ�q�O�m��h%�`�{W$oO�M2�	�GNR�P��B�)Ò%��.dÝ x{R�sf�bF�"�@��G�g��̆��v.��d<+tgź�u�o5]J���++L;�έ��53@��b�`j���R�v&���؛PK�W>�,��V�N��u�;J��+F��
�H���IPK�1���V�
LV����j�';V^o4Wј��4[@����(v���G�w�>+U�jR6�t�m-uy/)E��ArSH�V�mS�M���k�ɝu�-}l��ql�����>��iV�W���ڎ���,�MH�W[�}�Sh��2Aⴍ����IZTW�]��m��
q++`��Hs�$�Z� �W�hd��`*�6%<�+4��yn\«�#B�������ݶ�A�-P����ɺ��Ej��m��3~G3w&'6n�ke +B���l�0��(Wn[�[�eiK�%���Dƍ��N���,/8�;�vۥ���۟�s2-��X�at�0�z6�N܏����7yGm��z�D���tݺEIg58VQoe����ܹ�ǵ��gR{od���Չ�b�%i5��+I<�λ�܊8�/�/(
\Y8T��������fr���8nM�ʲ릐���<�`}���r�N��@�,�ۇI[�͗WP|0��e�R�(��yi� Q�OPr�N��".]�7Q製%�b�T��i�x��PKj����<����@N=շ�hl�P8��E�W��⩱l�B�gv=�/7��(Zk�.�RpԵQa�kc������k�0J�$gf�ܴ��+/��r�;��]�DK���wF��=[o���B�*)�c��'w2뷣�KaEe�;S*��4�V+a{�ifPwKY�n��g��!��VꠧS�;�ɽp��c��������jWD����-���y�L�$�`'���rS#.'���+1Yw6,��A�^����o�և�jӈ�(%==����q�#6=�fR�q��3�����ל�t�\R�B�D#p�"�����n9�� ��13���f��';����q֣ս�K��1�ra�6nՇQ`<��gH�蔷:�7s����:���)��6S�:tF/�%l���]��<���h����nln�p}e���v��z�+��dJ��ԟ��Q�0�V� /q���&cmv�dt"�%������f�[$Cӭ�LV[��fy8,a�Fڅ�#��;�J�u���"�Y��;�Z�]���Y�tU��M`F��R��e�Z�u+�,��jC ��/Db5���F=2��M�)8t������47���N�O/�Нhds$��@�'\�%�#{�M�E�D��S):��;q8^�O1&ލP�z�؛��2���D��򥺲t�X��r��ծ�ډǼ39Q���;�	�N���ƥ�+�ȥ��Fm;7�H;!�hNz��ݝB�>IIDQ�ҔF/��QN]�.\�I*��2��AQ��r�II��D�ѵ" �c&�b)wp��B#b��E�`ѓL��A1\�$w]F4�V�r�0jP�1PJl���%�b�FH�L��\M�j��h؍�j�fLlG9�Jh�X���6CcE�$�j
,&�[\�BŹnX�
��-�F�d�.�&���cJT�ts"��F��E�Lܷw]3 �DPF-$�����X�`��)�+%�4���D�زi'u���Hذ��������(����H���`5����DFHܢ�Rh��FܮT�]
��g�A�yK9�:9xv��)\��kns�.���8	��W,Ӣw�#�"S"QjX�'m���]��%�K]�kU����~ *����e{�e$n�}����/����c��q+��o������$��+��{[�J��?\}�h�j�8r�~��Y��Κ���x�lˁX��=��i����������Dz2���gՆ���9bw��i��мN%��t%S�:/�C�sfX	E\�.��<����ݯ:6���)��u�ϩ���8�����TY?u��
��)}���S��5�oʹj��7I^����O����q�c_��<�ԇ� �q��2�E�v|P����Q�ă{�|P���T�#+��WIe�Y��^��3�}@>����q����rQFV��OF��훫�C���/�f:�{���e�yw�u�uĖ��z�y�f��|o�j��ra犜>Ѱ�!N���l���@椰&u�o��^D>��E?+����#��x�.��m�!�YTgb�l���٨?gwd���~*@iAfx���az%��o��7Y�GZ�;��u7FkO�e/U��*�Y�F<}������n=�\Ozg�C$��L7p:�������I���-���{,�Trm����9e� T�ǵ�k�4��5w�Op�����׼eMBl��Ϭ�ˢnu]*;�yG��'�w�L�����l�9É��@:z�\�RL9xnVv�y,p�ĩeXȧ�znC�U��9��թ�mvʱ#�Ivr�H$�������������>��>J�.��F�:r�M�Hw�xS�.{wx�z��Yf�&�~��ɕ'�G��>}7�s�w�H�_G���\B����f�@�~ːQd�mOK�4��o$y����B��=�>U�s��l��T=:��ǽ�WF���u?_���g*�g�ó�T���Ϥ<Ox��a�:�;E����7�m���O�h�C�P�ٱX�|�\s���J��A��t<�ɜ���A�aX������ۊT��9��n;m�yp�d�.��௜__%ـ�Ly��I�ު���߯xߍ�8P��͙��CgC�����ү�������}fp��d�C=`z=�<�L�_��N���ޫ���am�N��N���yP'Ȱ]Rq��"����Fd��]���q�r�F�`Wؽo�F|���G�������Hjɞ=|J_+q�{z�oػ9L��}��UC��Uq��T�q��vE����+��+և�d�p^�7ꓭv�+g=3J�e�zɣ����~2�fA]!ԕ���LBf�[�����*7�<^����S*�!���~�֒#�W��gt5�)x�:�# �5_��4GEM��(����X���ú��{k	$�Z�D��<X-�K��X+o��o�o�vl���V���ըL��oN�Ւ�Ǌ���3ї\��S#��wp�q5O:��J��[�rv8���{��ɘ�'�����V��`����b�C�����]L��MՉ�n����sO��r﯇���SwO�9��W� �2��Q�P@�,	
W���e��|��yx^JKb��{Z�ȹ��z�ё�o����z�=냷�f��ʀZd�H��,���p]m����/w%z���C��}�l_S�=��&����7���P̖i���'���8O=7�\��Lz'�]F�g�/��ƣZ�-?;c�H�dx�O���=~���}�',��su����LѲ���u:7JZ=y��y���m_��?z�>�� 7ޏbnO�����!;��:���=u�f�K'�%2�^�
��^=e"���T?{��q-d�"�7��v��Q>�&����D2�uP�ċ���btqp�C�����ӡk���zzG��`��L+�j�)�q��W�>�W��z\��^پ>�8n8��C&�Z��N��=w�1�$o��^�XO���'Hz�n�xg�זF>��{�0u��xzEp�>'1�����*�ЍW�<���19�.�йb�� ���N�
;��\�r����tXҼ��B�蒼�7*cB��e��f�c6�����̎�U��RЂ�L�%�y��$E����b���aҬ���̕�]�Y�v�]ڛ����%�hH������chU�Ѫ� ��+�s>�fT{Լ^B�X�9��V��^���)�u��W���|<?h	خ��U
�*��/Į�4���"�JnN;��Ӑۤ6�u�g�}�s�����^����>��d�����L,�U#q].�Ι�q���mz_��5�:bzq{՘�Y�e�ϡ�Ey�od-�+:rN��rIꉔ=�rO��}��K��~�6u���/A�ݟ�ޔ���ܠߐ<�3�|�>�S�Q�Pg8�=�Q�rA�2���XȩT�W���P3��\3�1^[VW7;Ձzh���6߯Æ}ޏS����{Σھ�9��%�|ITe�߲0qaÑ���}�<���s/�9���O�+��/�oף!{k̮�;���u�\�M���oBFnO������~�0�IJ�M�t�e�Q��F�+����X���{}����{�GW
<���LY��n��z��2d�k� ���&[�������C5��F��?[dx�x��a�R�]���`w_�%Wd�p>ԯ��S�3_9�Z6j[7�� �J�J�<;B��o�U�j���\~�?mZ8��:����'��.���n�4��/h/e�)붱D�z��w��|^e1��K��B\�wq[宖Z�hݣ��@Gl���}8�"�t��F�|<�C����W55	��w%�*�_,�
�{9˴�-���Z�|S���#��c��U~���9 5L��qgT��|5T_�[�V:\n�t��~�
^���K�a����Gy�]фߨ�~.�3Q�]>�$�"��0���p�������j��G�y�<��h�>�������wx�o�t-�:��ޟ z�{4X��ԃ]>%zٱN���O���S~��W�[�Q|}���r��9L�>}�4�7׀�~ڱ��/�br�=Yו�/��&��?zY;@��l��;��#qS/Iӑ�_�����"U{�^��ә��bjs޹{Fz<�ҧ$o��vZw9'/���n �2}:�eW��^%%��^w���,(����V�-���zy��;�X�|�������:K�]S�:$�SS~�ں�g�V_w�����g��oާ��}S�Q��s�F/ngYd�\c+�g��Y��HA�w\��V���a�ⳋ�#O�����5�}��+ԇ� �q���\k�Y'^�}�Uc):ͽ�&+��:�qS+���D������FF�'��F��}q���9���W��w�^W\��nmoqV�c)�p�����R��aՙ�}���Xg*D� �����X��. �Gi��*ك7:�wƴ�a��wWη�pV�n@�h�6���8b.�Ǻ��%<�@��{��������=u��,�9)ݵ�օ*^mC���+�������F�F�̿��@K�0�L�Q��O.�|n"����qzG���@zn���z��ƽgz�TǪ+��]MzE�2���6O��<�������x�����S��RGT�	��^ꍯWGr�ND�t�D��N��}�,����zB�L���iO��2�E��*]�;�ɯ[kד>B��_�c����s	���q=~��Nd�J���2"J�
|l�2Zȼ�[��k`6�*.��W�fX���\����~dyY��L�%�F�t�'�'�L��]`��cٞ��	Χ�&l�}Y)��G*c��y܏�y]�^s�|��|�!���~ːk�u]�����D�.��W>�v��ʊ�պgK��ͨzu{)�G�����P���i�X�-���sb���Hq�T+�_d�>�(�Q �|F�~�V��/�����on|����~#4EB ��������Fq��}�Aֲ�o���3�,h䰯�:�W��R���Ͼ��s��=�/ ~5���]�!��?}����Ox��T��׼n<m��#㳷�L�~��·'$�w�z�#������%��^����xjk٠��~V���09X�i;ܾl�J��o!=Qu0�
�"b��I߹��^
Y����4CC�Ł�{V,��'^�b9!�6X��lĮݩ��	6�)𙶁ђ)�Y�u������ܐ^��&�Ǘ��6䏱��[sm�9rp����vWzuxc�~�>�g�顛���{o*t�Ȳwo�0�w�GOVB������>�6=]5���Y����?�o��r=u�ϩ��!���[S�}=��*�e��Z��s�'���vzc��R7�_��L�][�/���^Y�C×��1�����}۫��.�J��z1�H��sĞ5%xѕP�(ϑ��Y�����2Yq�0�x��ؠ���N��v����ȉ��%R�	=Q2����C���n|��=MՉ8�Խ>׳�����r�~Z}��|w�3�ΨZ��.�P@�2���x��l��˚��K������OvJ�Y�W�LMĿZ�S�#�u�0�䲠 ���7�3;�M�{�����hS+��|�Z���3�^�ZdO�팃��c�ޮ�oｾ��7�TM}�gg�7��ش��>���g��������������kZ�.�2�H�x�{ӠF[�u'��m#���Bu��6g&z	Ď���7JZ=y���y���������圯��.�[�Y�x����fS������E�<�	��F8�=Ж'wq\��AA]�1��k*����z�:��ą��;cz��$Z{���F�����Fb�_���L����s�Y7T1�Yѳ�+�P�}� �֠5n�m}����Ka��,�[����]�p�)���y )z����f�O��Fe��8*_V������R/J�~ۏu}������iĞ�=�|�=�h�?z��124i��:C:�����|�J�98���1��5(�1�ћ��w����>~���O�h�>�W��g��=�VQ��3e}�Ī0��6�5���/�4�.�z��ӃЯ���wW��۽	זF>��{�z��^��*p��Y;�ю���������G���)� Oa���\l׫A��U�[�W��|��{Լ^B�X�=�2v�����ԪO�yL���<N�1�p�Q묪�T��+4� bn��U)�9�5tͶ2�nb&ƾ��̜�+�Nw���ϯ�S�z���(m̼ ����T��K��r:g�ƟW���ћ�����['�/�������y�>U�����7'E2I��eT@���|�.:�	s>�����Լ)g�:�.}���W������+>�;�m��L�;eq�h��)�!�.&��c�jDyj���gQ����,ʟ����?_��G����Pg��w�o�Q0;� w�'�HyZ��P���I�&��9��Y����Jo��D�=1�[�&�]B[|jE��(�n(�r�0V���rݞ~�Q�N�co�׻�Ɂ�������׌��D&.Yu�WU��55T@s��6�1|�0�w`��qw1V��n�nSn�=I���qL��iH���3���$VL��:��/����"�^��3��w��'M�u8{'{�ӵ?h�7��t��pr|d��ʠ�t	��\M���{��r7��&��X�D��{ޝO�Q�>�R��U��+ﲩ��s%� 9��"e��x������5�Q�	��;�>C��f�Gz^H�NG��NA�s��"���*ZD�4e6h�0��RqJ�<:~"�s�)���z��Q�\_��_����㞙��' �sl�_"�H&�V
�s�4'�CwUܣb��>s�׮��!����ީ��y]ы�M���~�@�11��t��P�'�>	�:���-���T�Q-ɏM�ތ��׸�F�1����~��p��O�|�^�.;�RY��$ڒ��a�Ҿ>�Q;b��wLz�n��r��jW�����1:�#��CƖ��&��+G�n�8l>���������3*FZ�'``���ݨs��z�^��#T��~��Ľ���p5�&6�exW��F}�>���;z�8_��$��O�ӷ^��eW%x�z6e�߾����V;Ыr�O�_���B��+����^�
��Z�B�V�/n��;�+:]v�@���N�:��o�һ����'��S2L��P��C���1g���{�̸�d��X���9��b��Y��vM�yK�DaB��@Y<c�ԭ��+'�3��,�Ciz����~�O2��y�r���tU��ߗ��ۙc* L�R}'G��p�wj}}]�e�vj�u!��J}�zg�z�O���K��/�^�즮;���a}�����)\c9�8��]Ո�E�7��Qh<��S8��������O����q�cq��ⲽH{��9�\�7��;�X��Պm�ik�I�C4ϊ�\T��hmUD��K,B�����O���P�޶=�ު������C\%�Sc<.J5�<I�1���}FXJ�D��{Q%*xy���u��7��x�+��ZUd�����F���K� )����ׁ�[-C������%��lyFԌX}w��[���<��;���t��dmǦ��H,�B�G�Anx�2�X���;�<*$��Uw�h�My��E��0={Izgt���q=z��C$���j uX�W����|&-T+��is=�C�I���f|=o����^3�+>9��K���Q�D�#,u}�/
ȥo0��G���po�	�1Q/iѺ�k��C�j�1m�H�j�w|��w���~���5�խ��Z�j����[mZ�뭶�m�[mZ�ֶڵ����ڵ���[mZ�ֶڵ���[mZ�����m����V�����V��5�խ�km�[o�[mZ��[mZ��[mZ��[mZ��[mZ��[mZ��[mZ�V�V�������)��%� ��,�0(���1"��� IQT�J��"R�����
�)����RU)
R�D!$J��EU"��J@ 	B�R��������$JTUB���QP�Uk(�0B��T$"��DDR�F�lҩR(�*BU$U(���T5�gJUE"� �EQu�*�"P�F�R��B�%D�
J�E
[b)EQUB���D��@$�R��BZ�*��E\  ���V�e, Z0֥�([h*J��m�j��5��`��U��QURچ�Z�*L���j�)�$���T
�h�
��x  �@+j׭*�Q�	U٫BԬ�<��4]ͷE(��1�:4P( ���EQF���lp ���t0�ѣE(
3��h�F�[�!*���* �F�8 f�����EP(��D5�-L�*������h�����0�i��f�
+6�k�f�*�Qj�TB���!"�(x �(�WCF�6�P	�j6�5��UUPU�b�j��ڲUJэeZ��(���T2,�M� ֖Ji��)R*D����� ���U��{�]B��US2�@j�	����Ӻ�
2�IH�`u���K:�W`bƊkM���&�4(i1[c�j��"�5*R�TTRH*�  ��h�SZ6��@��Q���Q�hvCV��FS(�N�ZE۝�M�hi34mIl�l�Ѣ��b�GaB���D+f��Ī)Q"� )$���x   -sFF�Ddb�J�����cm�-�j��jR�X����lJ��6Uam��J��Z�����@�6fͱZ�����JAJ�*%��J�   ���4)&�(Ԫm��&���.l���Y�t�N�5R�� ��T�i���X4�Z�kMh��6!�6ȨC �C�]�8H�Q! HH�K^   �����A��t1�ڴJ�L+V�A�������lд�j�kA�Y�kEjڕ5��CS�D�Td	�DB���)RRUTk�   �VT��ٯm�l��F(UJ�3L��kj�-�T��T�� 5Nȭ�ֆ��`�҅����SS��*�e4(^ j����JT @��a%(�L&@���MOHњ� )� �*   "���OU #@))�*���C�#�$B9�+(��`�f&��	��׾F�{�_{���������
�� ���S�Q�D� * � (��?�浬��f��c�g�t�:Y�iX�w,b�{�R�"2����m�L�W���۽W	�#�f��NV�LJ�i���77��؀o ?diGgM$��$�6:w���LE��l�GS�t��-1&a,��d��`�$�5�6�@V�+kFm�Y@�[�݂�`r�e�,��S4������7�ŉ"�H���M��u������ ��]=n���TZj�7��n�˳W�d�2���e��Z
��/�VfnV�V͸����9;K�+ �BR���F]]�pM�NB�[_n�Y��-�3�NyE��6 2ص��<�dMtl����`��Wr�t�6�T��".��D
-F\3�B�ؒf��VF�]P���"7��wB�]bb��0�q���p'w��i�^
J��4������ڽU�+k��2���IX�V&ܴ��ݤ�yU�M&1Q��\ʸ�bR^���k_M\.,#���YW����#X�wͨlU��Q6�KN�͢����r_=w�hM�n-1�����Vj� ť��f�Bv]
��wkZ�n�����C%�^�NK:�Na43�30���llŬ$۩u�KB��lFM��#,� ޥPb@e�+s���=вZ�I��jY�����H{u�F������E$����9)TET��"�%���򴺟IN�υ'u5TS�(ш�����U���ڢ��ըn�ۭ�3X��â�:�+A%]��՚#�ŀ:i�Um�j�%��EI[bQ`�ً#��&J����Qi"��Kn˧rn�,�U$.�r�ʷ�[瓟�
�(�����y���-E�����[Ms^GV�Dڒ�sKv݋hr�!��S����R�p�zud�5���]��zޙG6�eӠ����i� W���V6��g"x�5���&O����{��n`�ƥ�̠�˙��4,��4P�B���U�l1��� �w��͟Z��R=Dr!�i�FQ�h��fX��`�әuw�2� �C;���	Z������m�m��ܭ��y̛����S	nMW2�VJ�at�Ÿ��m�S�)��'�	��k�v�!CG.Ҳ7��o�5��ֺ5���[h�,c���@n����5��D�RQ�vF
���aSZ�Fh]H�͍��G���Y���2/`J�r�M�r��	nL�WC["U��n�hđYXK��v�f��ت��rT(n`�H/$�B�b��5��i�;/@H8�1<��e�x�chG�5��|��Y�n��q깩��gVlDַ���V`p)��Y2;[���"��T��&�H�������趥;"��4k�%n�椵�b�Kq��pbV�p,B�ytRZ��v�c(}r�e�:��oGt��5-l-D����w1]U�0V�aJ?]^V4L����Ѻ�� 
?�:�e[j�H1m-;�,��2��(+`ܦ�%�;���c/k&�Y�t�
�V݈Pυŀ%{NP� P����+�T//�mJҢ��=���Kk�IT����;���T#�&V���(�(=VD���,�QT��בܕ���`'f�8\"�+�D�m�W��{I��	J�C��x������(��J���F�+D�f�*��lJ�n�j�#6-�*�C��=�MimT�X�B���ml�h�C<���K�J�2��n�Kiá&bI����uMxi4�A��Fo-UJ �ec͘�@cW7,T�F�Cm�E����)��z;�-a��]eX�ZD�l��5MWx�:��^@�۳n��d�%�e���^���?�n�.ٵyٗ�)Vݥ�p �"j��3C(ѵea��a蒸�:��EZ��[x���"�(FX�B�-!Y��c(�7b�L�MS����V0�v'�^�z���Yyc	��)Z)��J�ڽ�tF	f��m�kN�r٭�2"��̠��Ю�KFS��U�nXMg�+e]����,Pl�$��ny%�3�u�7(���^C.ٚ@^X�mn5v�mGX�(���A�a��f�	v��òDВ5�����aLYu�bă���`wR�v�m0�[g.65��S4\8���АӶ���K^.�7Ebm�V]⥚�0@v��Y�m�aV嬐�X�/`XpR���ݸi V�qH��!�[��r�-X���T�����P�Ød��Cj �
ac[J��efԚ�#$wn4�	�o,�6VȵD�����C%��B���㙺d����b�7F`[{p�J��6��{S��L�)�Q�N��r�����Mvh�4���ܽɆ�Tר���D�Ub\;�*	cv�����9���wL�д�寂zٸ��-������-cOTV��D�D���߲,�eTȒ3iZ��vv�[�����4�ڱYUw0��ĺ�n�V��'�4p@�-��d+�V]w�͝&[�Ͷf��l67�
%�nŃ��X�b2��mL�V*F�^�v�z�Ej�b5$��OFϵ�J�Lͬ��*N��r�T��H���x�%��r�HŚ�&8&)��N����(�r��:�!t@b��Yi�9p�[x��EdF2��[�#^�Q�)��ɣ��{.֡iP± ���
��e;�%r��ǆTP�X�I��l�V�LH�W`4thǙJ�K�n�;eR��XCI �
�j÷���f9�J"�����GJ�`��$���T��L�V�i�qA�E[��"K�]��Ld�K�WQb:�K7 ���I0ؼ�Zt�\W6�
��$LJ�&�ͼ�b���-K���mZ��Y���,���&��*V譈S��yz&��ѐ7�mZ�JXjXϭjPn�rd[vQ+@42��q<�L��.Kw����]��R)�b,v"���yX�eӱ�Kq&��ܬHY���J"��˥�!`e"T�6j҂����P�ͺ�X�R���!򁭑kcI��旮�i�5�.櫒����Ě��J�v�ֻ��ٌ���F����+o�P�F��9�A�!)Ca�%�͘XL�I�h��E�[�)�7,���hb�d�0�m�tVSk��x����T���Ȱ�{[�V�9���+Fd����J5W�����.��3-f=o-:"�5.��OD����Y.�;�VƀYYX����7-c�Ks�E�mnS�Q�U��X��q%��uʁ_؍�+n�E�(��h;e���I�0�:��[�U�# �mXi<0H�`5+/i0q`�r�3%#v�ДW��n��T�i6������b��I�]M	��M��t66�/�#�kn1@غ�*e #��N�Z��B����T>8.I�f@�`�r����pZ2ځ_-��f��,6�G,�X�Z��驆,Ҿ��ں 9���Cf�Js�V�bP����%��y�2f͢�KT4�TݘlM�Z��O���&nMg���R5tIo,34l��(�*���K	бwNm^pe:7*��&���=�5�2���R���*5r�[Aj,�"E�,\G�ɫ5���-e�`5>+PX�(	%n8I`��iF ��#N��.�A�Ćc0\��Xmn��Q�E���M�7�㖪���=f���m^��B�=�،eǛ�1�T���LP[��Z:�Aj��#+p`P��Jx
Ů��!%=�w�)J�Hh�v ��Kk2�[NQ�9��F5i���NSs%�A9�wFCϢ��ˣ��m!N9�X��]a-��A��l-VpSE'��ܭyBɡ�M��kk�m���w��(�v�Xq�MMڤ�7w���9P\�
kv����2l)��� �ޣB�=�7!��Bp��k5=�훁-yf<�I�p^mxeT�Z��7GiM�Ɇ�J���r&����<���\Or++Idؔ.�)ch����M;yB�IFH(0�MH�H�7�[9Bɭ��dn9��Q�1:4U�-���h`c2��h��JZ�7�.Q14D�2�:�/VL��#N��2�7˘���3)l�)�]Z���V5ͅ'f哛�E*N��P�p2�J��jU-��jd8�2�++E�(�G�*��0b��7�cٳ	ݡ��k\+d�E=��c�E�� m*�i�h�����Kp���M-`$�4=5�P�G;��;�oq�x���5V�1�MD��V:w��Ĭ���з�B�q���%�[�9a�`l�m2c���6m�)G-V+oZx>Ԧ��5�\q��3�B�l{@nfJ�7�����x��5sUm(@���Bc*`vv'Y{l��2'y!Z%mcxk"�ɚ�d�Y���%��m�	��̍V�$f�\��`W7j�r���%C��]˘
�%Vf}�w)-�9��F���#Xyy�$���+�[�bP���a-806�]f�wh�i-$�܆Bq�VeA2����7F�9���� 2��ʼWC�Mn�X�U޸�c���S[Ԛ�[��n���Yu�j�L���F,��+2u� P�k�&�
�IFk1�Z�4��m�%��-9>�p%�+����uj�=e��Y��*6��l`�h'�W�[��oC���V�j[��]ec���u�%NE3#������\��B)��k�N��\�cj�`��a���3
9�$���l��˧v�:^36j�VV�f=�ddomֆD��j˫��)]V�P/pBH�8iE��	�FH���+-��r�����˳t���I)r���r�aQ8Y��6�<�n�M��!M{cȓ��ԓ`WZl�u��@��e��v���򍴁Ͳc�R�ȱÆRC,ᰋ�@-��0�nR̒��(J��)���e�v�چ�`�bPutc߭�ۛk5�
U	T�܃v�tQ�a�K-U�b_�2S� ��(�WYMI�N�a3��4���S%]�=u��F�mُS�H��ϛ-�)LT.)�Ǖ��6��ڻ����0[sYıCh�`�(�"u:�*����VLV=&��ֈ�Y@�ITI��kPL���n��QP��[�0 ��q4�^&�l��S�i�j�ј�-#kU+�	�Um�]�R�Oi�wF�5$n����x�6&p�/j`2$�d��q�1�+譿��1��4j�ӬpK0�Ӡ���d�;��Zc�(�
pݽ�Q�WJ�m��"���-��37-�O�ٗeU�L4&��f��b����͠4��T˖�[��{����ѵ�L�"��ؼ&�,��M�V0�Q�����Z1��noN�[��Q� ��[6�;M� �¡VV�Z�عb��G�����]+���\�qV�m@�<&��;Ux�-l��qFՍ�Z%m%1�+6��+u;���j1��Z[����yFؕ��#SD�z&��0�nhJ]��J���FJ
I��Ҏ�O�y[�L	9�,L�7�	qh�Xq̗�,%cŃ^5�����h�3n�`��-�Z�į�u�w�mpй{���u��_�SWN�d���Jq&Z&٪�WZ��IMH�7L�A�f��"Jbkf��2%q��j�x�h)�	N���Ǆ=7�:���ۊ�i��Ҍ�6ڹ�����z�O\�l��C�
�6M+�s౥Fka��v^���֛����e��Y��\!�|6�_K�kb��H)Q�Y���WPpA��jS�~˳J�)b��m����y*l�a�(�9,�W���F�k��i,vd�[x.�&���o�P=�������x�+L�
ƼF��aT>�&V�Ӹ�����E1��(m�~����-Y�R���f��bb"�Xp������赚�jz���[w��J�7�U��*��>�&��Ȭ���yz�e2�(aux�Q�09[>��8��f�Y7q���MM!B�k��.�U� �a'
7.�ڔ��ޢ2,l\+54��Hi��%����JwV��ne����,qC�	vٖ���C��	ѡ���[�����Ջuj��"�@�2*f���7*�b*5�daZ�W��ci��-e�ib���4�$��S(�-�2�,ù�9��4e�[(2q� �T�KJ��Q�>;�V�JA�	���au>�$��u�1e�B���[˩�)<C^��E�5Ea �c��B��ٙ[R�[���cM�`�J�k��J��y�h���� z܋�hw�އi����z� `�&������T8��eT�+�N���@fRݍ����)R9�E�[7V<	��gH�m�9�m܆Z���fR��j�*��^�Y���FU���m��9�Q[�6���eݕ0حWPf8⸑˵�"e�w�5퍺�`�D(��HJEV��zUK�ټƮT9�Ÿ�[B�MU��E1�m�n���"i$���%aP�gpH�lܻ(զFi�~L��5e��I$�ت��	t�iU(
Rn��Ѯ_H�ɕ�c4Mqǧi�!��U�Ԋ�u�?J��F������[�	aS�ۭ�i��n�k	ų6��Jl;���˕0,L���e�X�S�X��Q����n61�X0�[�SWC+m�/�S�/FbE���������X�A�*�5
4u˙G2��1
����tdp�5P:�;y�(ށ�Z]�m�b�%,b�x)0�Q��E�u��Ѥn�8�Ӷ,2F�:H�	a��3E��/e�cgi�)��N�nhB�Zǫc£0o/뭬��o\�S9�En�vj�É��WKfY̭�Q��ږ�&5�m�17Z�GAk:BD�@�h�5�`/.k�FZa�ff�z�g��!$�= fM���hԭ�5B���93@fޤZyN�A[��n8���A��Y;׉ci�a�Ks�wy3}����[�b�7+�FNf�.�@����^l�!]�`��</�֥,l�{-[\���C8�C��\�\��"K���Сw���M�Y�hWN�8b�PS�(W^��@,���Tr���A���b�8}����7�e�#t*�4u%a��Rŷ��L�w#�T�,x9��]��jT�����V�;ɼ|-�BU�>���άl�rJf�b�(��X�u/HNm��<34P	R�걪#�H���v���`������	�:n=�7��!�t]����aI^��9]j���V.�-ه�0�{�j��L���*�:�Y[k(�(�|�����m�|��s��v�λ�&e�((� �����t��:�OZ�QlT��n����]h�ᕂ�%3O^Ǭ%ʹ�yQ�"v�A�,�N��h[���d�n�7$���l�3e�&��,d�m.���-�w��{��x��(:��鍰QX��3i�<���-�MD�r�,%X�pfv�k>:��yZ���w�G��d��S������߹�����CP��x^��c�$���n�m��P!�� ��e�b�u���a�B��hC���+f��Cb,ߧ`�'�r��(=� ��o:c���X[�̣)�%h�|��@����X���4U�]�x�R���0s�A���0��`!��UF�h�������]"*ڻ��v^i�2�S���o ��cK��'n-a�����'��i�o3	:��B�>���ۉ��/j"8=���b�{V�� Q�wV�.��o���Y��[�+�3�ƖO�-d�`���,�X�Ag�����G�l:C�z�����x�9`�n2�Y���"j��euv�E:T֩���Ǧ:�+�9���=Y��F1�eJ��J��_dM��(W*5u!V�NN>�8�k�v��r��,vC�͉�������J�B�.�wi��t�u� 5>R�tU�;��6�Nބ����|"rA��>]�(u�g�t�oI�i�N�U����W�y�jȹ�ҋ7��f���|e,���(�؁���;�}���w��
���qJ���۰:�*���K�03y+,��]��g��1���v����k+���d��lג��+��g	�y�]��Q�n�k��oVY�6%�+%I��pebD&d�t�Q}���#%�SF錆^`C�k�/���Ź��_̛��$�̚Nv�]v�<#SR�yD�J���"��s��N�Z���
Y']��J
�24�c���g��&��3�4up��`��F���BQ�el@���e�5:��Й
}�v�zPt-���i�c��l�U;�M����OǷ+n�L�Χ5�\�d�}ƈ瑼g����J���:,��5}Dٶn��v���T��	��
�O�@[mK.n��N�-�\��G�ͤ��ɂ�"lJ96\�[�9qum��r�G��y�Qgww��l�W[:��kO<;FAd7LRw�J�紺����
9�,vMg�Ve�YW�O|)��+C̻i�u6�˄��]h660ϥeG�*eJs(�wB�@0��sv�Z?v�̃�\Sk�A�t��b�p��3��j*�	�W6�r����7K�[�t�ٜ)����2�Nŗ�0���{�y���'�4�د^�9Y��r�N��)]f����H�#bg0��f���[x��I[��kZa���VMtoUM���^�=�΅�b�������J�.[v��@Iώ�ս��+^Puz�ڂR�H�S�JI�)vM`�Y�V[y�Bs
�p�u��ˀ�b����[��ۯ��X5�N�J��N�L�O�9=�����nu.��m5�h�xN�w�Io{O�ݤ���8�S�ʗ����J��>�u�4�1��2Ԏ�w���ז��E)#����am�wy.ݮ�ᓄ��3Ua4S��	t�?8�:۽*��|��db�n,��cc���ʖ����i��^��)u�K�Fb��T�[fS�����9��ϵ��	).����ǟQ�u��x�}Z�۾�<�7�t��O*v�s���n��#��j�@�
ǃh��FGQe4Gv/�{�4C��w]{ßk�u������7�����v^"�>�T�t�Vs��6(��{�<u��r�e��3�����O���y{�u)�:�T��y.�]u���y�,2]_1Hv��HB���3�sn��֥��rjn���?kQ�H��DE��γ�F��qh�#�_u���x������v�����y��66�}%�y�3>�y���ok.V��'�L�,m+Wv�C�u/.ե)R���}�m'v���ئo`��cgd�w����E��X�*�K��J�:S��o�l��F"�*�B�8G���Vӏ�F��@N(ohw�P�Y�
,R������Ǉ�(�UĖ��vu��Q��.��nq�%'7#g+y�\+5��6�K*@ȼ�#�D&�8'O�~�o�dɰ�,���\W�ڔ��u��ʜoVs��j#�{.�ݣX�Zh��iK43es5Se���\�I�0Λh�XlZ��6�톖5wy��W�Sa���~���j��ؤm����w;�Ih^>��V+bC�����Il;�Ѐ:M�R��Z:��RҸ��G�Q�.J.=��2���;*�96���l���Q7��Hp(��cY�{�l�ܶ�az�k�kL�n�*��_:��Xr�$�N5!���ʴ���܃gw�h�oi�<���H9X�ˮC ���������`��ꙃ,Na�w&Z5��l�9�vN�ōm��<��Ŗs�)�i���`�4D���q����w�'j\0*�3ڎ�V�p�\13ɜ���[#Ԯ�kwm-Y\� ���o�	���}���%;��ؤ�Ԗ����s�Yx�gu���X�M�w�ԃl�� ��},c+�>�Ӎ,�w,*�GH�[�yBT�jPGe��\Ǭ�fb#��Í#���+��Y�[7�[1Z��2M�d��u4k�m�cC�*
�]������&4"��٧(,W��S�E�Y�+3��ݑ�[Qӎ�]�.� &�%�����M�7-�k�a�4{l}(b�U�c�[�H◺�6�1����|��7���P�u�U�t��ӵL?���\-��X��l��x��R:�ǎ���6t��\�|!�\Đ"�fC��(֠.�f��o{rF���v,�u2��5��s�V�z�P�#�o3������G�ہ]z���t�m�)ݕ�墲D��18ᗌ�;{�B�R�ht�â�UгSh��w�O.��q7�gIZ{mIB�C�~��r�P<�E�,k�@�zL@+6��}9.��ξv�f��b�;gx�N�V�[ۃ1hMe�}vv�G�^w�][�)��v9'��!n�P�j�������Ù�����hst$��o��CB�Ǫ�Z墀�͍���H�تmme�Ί�A�Y�îq�e$b���6Po����Fu��r+Y�F��w��M��)�q�7o��ε3e�u��&�m��U� *&�Ta	1�ٸb��k��͛p����:�\�������-��VvVY-3�V0�>�:�[�u�jǊd��m��c~}]�ox��s��U��p�"e^���[6���.���Lo{�k!	/�1.�ΛN�l.$�}��|LX���M;��4%l��Lr�m_�Y{��ѻ���'�6i�/n$�B�B���Km�چس���Q�����z^���b���:�oַ�֦.���L�K��^�\���q��\��ѓ �n���R
OR��p�О���y�X�眺|�w�@�o%#���ޤ��5R�5Q���W��ʓiV�;}xq.��>~\�bʅ^W)g�����X��_hyϓ����1P�­� ��������e��!�3������NU�bt��{�J�˷�e�Y���P�7b�� ��@�:酙�O�q��>��ز�n�S�	�ǎ��s+v+޽��3�s˕/v�Sc���K�%J&8SX�G�4��}�����Y�9I��qJ}[K���+���&�V�����s7�?G�J��f։AG�i��䣶���L}��ƪTEԊhN3;;��4�oìu]��XBW�k��^�k�8�����f�[I���c���5J�0�o�2\�[׃��O�g;mt�=��jvts�:	�a!2wG�MdC:,�g�����Wö��F�k�A%�++�H��a�Y�^n1+^Wg��_^V�B�L	RӮ�lBT������*�ݤ���ӒNEgkע�AoJW&L܂`���g	լ��иem%�)D6�.R֣%���۩�xZ�c�-ή��0c4�U_��f��+٫3:�����c�N_u��\:��ͮO�� ����
qQ�|���|.X����s}O�pFq7sV<�(TΦ� v�De άżx�9�ʸ���$����%�X#F=���|��i*Z�0ދ��dĲ��+��n^c�����{8���1T��M�H<ԙ�]͂�lʻǈ`{�-�]n\��c��r�1j��v��3�Y�B�H��t	�W�ټ+6�
�Ifar�G��U�6�F��,�Ȳ�]r��Z�CŅ�n��O�����O�.�q�e�P������ա��[sub��p���P�K�wA���Dn���e�Z�i�cy�د�2n؂�~��;�
~Gs���L� �ռ�	�9��:�+%��.��lQV�S��n[[��[��/h#��a���U9�n��e]�nES�Y��t�7�^�f�0`f��q�ʾ����0���@ik��E�M#����l��{g�|����YqA��4�������WrU�u̢O`}ۭ������x�8Mmd'��9�4��@������l���,�4���ܬ��lV9*&���hS�Y�I�np�M�����h�|ч }���#�I�]���J�K���ե�w<w9|���{>'hďa\���9�a���d�^�G����vறC��yY]����D�vɀ�C�</^	�!9-�G�AY/z�����ރ����Hv���yzbˇJ�<4��z��eP����g��5t�z����k�ee#��{R���ZYwV.�r�Pbj�ᴓݼwy�)y�uEs����j$��2-�a���!o5�;sV�B]}�u�ks���Ѹ�,��a�W5$�+<#��R���[ˋ�����r��ΐ�ڑbmrkZ�ֻ�˺�E'A�@I��P�TQ�S=;{p]B#�ȫ�	yOO��u�c�Z'{z���R�-�W�b$ooU!��K�u}Z���[���)U�gW�ݷ�6R5*Ƥ�����[)�L=;�+3��MVjvB��4�w)�⡩��T�vȎ�_�^�wTk0rM�nH��M�N��m.�8�b.0o]l��c����C����(�g{D�N�����ܵ���Nq�z����W/� ^Z��u�z��� ��h�{ה�����b�ͲƷ������C�,`��X�]�Q�W6(h�,ɒ��Rds2�rγdRgk�-m�S��W���R����6]bR�ZQ<��ƺ'>�6MO�b5ǐ�3�%RWW� Q�S^��g�R6]q��e٬�;���sF�MꎷH����ؖ�gV۵��Nm<���z�6Fi�1�場
%����{{�Kz�aX&�Ҿ�'z(n�$#s��G�r򺼊�Y��yF��{�Ƌo8vVvΆ_p��t�s[S ��C��eY�IJr�bq���+��'���2�$;4���k5d�����J̈���Sn��q`;H��p]Y���,�Wo��c���ul���6� ��a�L5��-{j�<�mlˎ.��-]�tCh���L����,�Z��;@.�&>�b�7����*0�om�|���lpu(H�*N������U�{��6^�gt	{��\��qC#wi�sf�|�U���0GI_V�g�Մ�C�<����*W��'�c�Cv�֛�c����(k��H���7�k5t�C�"t��\����\��eɍ�����	������/�t��-�o�2�����u�.!ܨK� �V̥�k����V��hȞj4^q�<_xp��Dt��J�w�y�z�_2s�v�.��3���Pݸr�Kb�0�vaLa���̩�!��t�&�]-�"q�و�@a˼S��9�T}�t��v){�dT��u���.���D�m6�v�5ta�*�3�5���M���O��<x`��C-�~�`�c�F��!1��[�YZML֒@�ú��5����B�9%�9�ݾD�s�3��]d�.W[F	K��F�_U�Xຐ��H,�VҢ�Q��_^��85Mw��vT�pb��.�؈��]����Sxi�܁/���U��+W��&�2�|����:���hm�ݷ�ݜc9+���&����|�S���\�s{�B����v��һ�� ���Qe*�9�m�&S�;���$���X}��\]O�t ��|����'6eh�fp\v�����ĦJ��1��9�9��*2kz��9:��՜7O��Y�t���\�=ED��p�M<�3�,�b���Zݗ�.�_q5o{'n��G��� �In7t��$�+�Q�"�e;!��!��+Z�pZH���	�i�C�4k�AOb���-R����|Y�E�-��ɶ��\�����v��;*��R��a<�CJ�>J1��ෲ>̴�2�n� r)��w��w������ve�A*�y�V�[T��!-}y$���Q�:B�VJ�9_i�HR><��X��5�O�����Z�u����&�"�ͩO�PL�njGV�2���R�Q�
_^!��j�������֦����m�4�����@���Q�* �����5і� ����/g�Ω�J޲J���[�k�y!]	HT��/�W�t�lJoޕ9:��0	ۙ�[��em���wk������O��7I]�&L}�l�k�J6%����v��r�#���rؔ�)L��J��+�h*���! $��\����u�{hW�RU�@Rh`d�u�ǻt(t7`�ʚփ�8���<;/���0lb�c��H�����}�+� a��Y��V�!}@-,}�]K���IF��^�-����<�s��A���>�	��]N�+ۖ�&0��ٯ6��ޤ�<����L[�cڷH�R/Y�^�5ܐ�U�� @[dSכ��Ȯ̡ҏ�V�r�&(��#1�4�Ŵ&ˣ�\�[�_YI�fӻziLK�}������;;+'S��03*-WNjW9NWإ���@��uz���g�.U�h �N!�*�� a�����/`��2�� V�}�S$�i�@���;,�0�n�ޝ#��ι �苤4Qv�R'V@��l������'�lZ;�˥�m�v`:r�ڈś"��v�:��7�h���_+��n�Ԉj��@=:��Bο�$����]��̻�])��*h+��N���0Z*���S�y����QV���njXA�+e_&.S"R��@,>�N��o�c�$ؾq<��v�:����)f��%n�*�&�s�:�n��1@֪,]�KF;E�1�K1��M��,�N:ueM�N��٭���-�p'��������j�k\��˽�hb�!黎��ׂ5��U��		�n�C'`��a[,ې2�Z����tf�#M�B����OZ��m��)�J���M�c䞪�K�[�9�R�Ю�c��-W)u'R2��b��əYn���8�h�hS�d�̘ir�Z�헭[�+2*���.�+)S5�Ɔ������Ũ|bق����e.tV�/c2���UK�*���)���*��D��-�T�r�es�s���դ-{��+&3�;�h�����*Vg[ܚ��׀Eo�ڱ���]ɫN�h���y���yO�h+-�	%6f��D����ɝ��oV��n�+�޽�[�n>$s�Sr�u�S��T|� @:��0�.ࣙ��]M��W����%�lwZ�{����(�-�O�rQl�����xح����¥�ø�4�4ؤM
�E{��soqm]���}��ж���kl��D�m� �W�͸B�`�j��W,�Q��=��1Q���{ן+dAϚ8EV�L[�K8�©�u/.Vm�w���x  _�ˮh�/
/p��n|�/��MW�h0o2�eWNNu<%��d*H��&��4��y��ռ{�7(r�sn�m�9K'Y������m%Q�vu��8�k�qy�Vnm؛��o`m���8b�p�Ksi�80Nj	ZA�wlf��b�p�
s;�5�٪S�nѠ�F�h�vZ���k>��������t�UZ�������t]0��_��[��� ��A+���4�zMw
��1����=ֆ���JT��=|a�ڦ9�� �L�@.d/����a`7C+�l�5����r�V6���ng�D��L���QRvL���ӿ����]1N�Ie�h߁��P��t�C��u;��0������p�!��7���V���|��"�3E�q�F���I���9X���b�#s]B��`��Ǐ>���A;�/�S�<��a
7-��R����vຉؽ��1N�k��ե+(�����ae��-��L�z@x(��kuojûi�D�WEf��p�D��ܣ����W@��,��23O7�RꛗkiT9H.n���«f��C�Wp��Iټ�;��Ѿǳ*<���
.��*��	�H��¡:�+0�ƈ�J'�L�<!IY} ����'_c��]E�ݢ�]Ю�v�b{C��̓����kW?p����{M�uJ�l�]8��nW?���V�ю�n�Xܺ�HDN �E.oU�\�¬��īw�^�ZC8(-:@����i��ȋ�a�i?�ф��%����D�劍t��e�
��G��goD��*�x��Z]f�XVV���z��>��&�6�K�^.T�X����"�Ճ#ͨ�u���k����0L���	{nv|��Qw�D;���ډ�m����.��OUo��[��䫠z-b�]�tڸN�C4Z�!�ҫ���]���yK�֥Y�rKH�Q�a�[�%a����ӝ�qQ[�����ZN�N3Ԉ� Xn_�YwI<hղ(����
�_N�w�u�A�F�)-[J��k��7��uVRG�B�u��"�E]Ҁ���v���v��q.ũqFl���j�3:�Sh��7��[�c�Ԯ����_-FK��e�Ж�G+��^[�^���v(+�p�<�HJ��q����tkn�ëql��L��@4)��ݽv�ZՀk}r�^�������\y4V�/�>���U�cZ/�2�T%��l�[r���,��<�v>+���:4��y��hCN�-=�JX���U��RDb8�eo�d=�t*T
�k�;��2ҢV*=ǮL�y���A��R|6�T�T��� ����nt���5WQ��2�V<�i3ۍp�f�5�k��υMڟlv$wʄcLwHJ��sш^�;��r�݆pdt��J�F�"o����4��V<�J� ��ʩdo�Igs�b��왊��qLB����K��8�-��k�RVs�Q|F�!��H�[�_e8h�zzi:����5m�rU�c���H�C��T�wлg���'e��]]��-�k2�B����i� T��l�?��%rd�þ��`��@Do#cj养7��wWK�]҉�	���H�M���:uɽ@;��t� ���[�E�������5����ow�u(3���W!ۆl�E�),��-eѶ�-��{�[<t�J}0[��W�۠��[��z� �,`i�O5����YN��H� �d�㊴c&�U�z�ơ�l�\FWW:�rk������^�s��ԍ�
����X����$��ԟ=�9}Bh2�b8.
e�ͻxMZ���N�鵥�6�u<��PWu0��S�,6�f:p;��ַ*�&ur.ev��sݑn���vi�VD���;���Yt���U��}�@	��6[Wu�HW\�b��Д����҆H8s��Eg�̴��H�wۄs�'y3@���x�f%�MF�TԶ7L\�5-�T�-�ꕢ�u�^��� ��I�@���֋�/z�u�C����*>�+,�J��4���S��L[ɽ��lqm���nL�U�^�zUJs�LR�amt�M,T*������`�f�m^ڭ�8]�m�9[\�9E�m�\�r���{8T�"�Kd�׭���f�N����eڑ�W�h>t	�3��3�����N���+�D5\��f���n�Tevrszk�.�;�ͬ�{N��
a���a�MP��(�Sar���F�Vt������x���SB��k��rD�u���/h�7�R��s4<ֈ��s��X(7��^���I]+��7��]"�cD�zGl�&*�Z9*�ی��$)�"���4��.��[���8`��me$}�1q�r��j���v(Zv6��"U.����.ʮ˛���@U�/J�Dg�f=޾��\�ɓ��S�z�)���E��
��W�Kiػ2�?�ä�o�P��i�U�i�����YI��Z�.��)8�K���d:����PƝ�pފҲH�}mva�5�n�B�f�h���M�Dh�7m�E�K�pb*ê���ٝC(;&������̏4�#��՜5��m��ۉ;��T���&��Q�J�E�O0wv�ӛ�M�J_K�͆�f�l��7��McV�-uŊ/��SA��n����JL��_ho�u��ӝ��L�{�����/a�2���e�PNIq�"�F�ӹxxef�*��u���v����N�J�[�0��<��T�b���L,>N�uv+��J �(�
�ˠ�\tղoK�)��h(�%n`��U� H\���[AoJԲmU��V/w�N�Nw;�+ԩ�X����˽��	����r 3jk\<�G#PF��n7�����Nq�ES��q�F�s{鵌��(�M�t�nL�kC��k"\J�6�(��!Жv���]�u�I���)'�U��a�喭�}ݜ_sh�����a��f�1��a(o+�"����QnU�F�S�#����Y�;'e��۠�ɚ00����|��.��4ƃ=���LHO�۽K'1�"����l]E��L3Fl��Ŏ��m���B�XlY@渫E�R�<t9R�\v*���W:�Yx��ƝIϭ+(�r���2�oI���h�.�\�'�MIn�J�;�H��%��`Z�鍽Z�V[&��:����ĘTn�	Z�H���om��P�]r�}�S��se�Ul��j8ų�JE&8P��\(�=�qT5;�|����J��%��6p�j�]�F+��@U�mrW��h���4)[���&�b��G&����5;+��*��o!�0�����u��k?_W+`�P�t�x��.����*+xgҥdzC�ޏ��G0P�Q����:D)�/dt�'D�g��I�JX5��}���@:t�ң��i㢹W��ɺm�(�����J���P�����T�Y(�H�7�0PĊ��A��ůwg:�W��������]XK�V1���tuc�8��P>��
ɜ�Ze���uu���:3�3Un��	�^� �{E�ǩ���;2��(Q���FͶ�ʏf�����"���gCE�; �v1�ϜC2C٣:olK3x��+V�i�\���Q��V4k4�i徻�;3��I3���;Si�en�����܂��w��	v^!��Iզ�j������!�1�ZN��T<�����vi^l}2��%��0𕰽7W%�n��][�]m��H8"�6�f����R�c���c�mm�ss^��E�BO���]��,�hiSLI�E��QT��5y��Pl��ᾅ�%s�ڐ�]���/i�K�)_V��Pj0ܳ����g)���ۋ"+Y���3���k���M��ZU��L�C䂴�U�®�%i���7G9R������->�E�v��6[st�Ҁ��-����ɬj�!����R��1�i6�q�:ok�Q̅���X�WC3�M£)���	5Vf�J��[�V4[���[o(�*v_j]in��*K�S/��J=��C,V.\���ͮ�<�ZAO�kAXǛt�qΊ�[BC�Zז� �����}��S�%��Ie��Y�F��6��H�d��u�����:����� ˭���:�1�O#}	�����[�����1o*@nL��VSF���4;�8�*�+Lp3�T���R�u�j@��V�1��(Z���)�{�C����S��j�@J�+~w�qIf(slQK��(�(��9.(��o�<���8B,Ԧ>���7aS�n�ϲ�HU��w�G̾� ���Ѭǎ�1��M�|#�ǐ���^���Je���E��
Z�o��^���R�Q%��C�u[΍t�AЄ���H�uv�/�Pg`�֨�c��Npڬ���ZR�
V_L(]N;��;�Zx�C��Y���Ie����q�����V5ո����Y�Q[C>j��z�3J�HU�#�qX9�}�ѻ�2e�����5����1�k�șH����-�jWn8:���y�q�"U��t	) ��k6���*����B�}Q�I�_
�\]u��R�[P&�}���^� G,Zк��6�L-��j�ue-�Q����ldS���c�Z���έ1^^bV鏺��ah��C6�*;�@a�KyLx��gew�����b��s��+��$�@�m�N��Z/�wE3{�Q���pT��ie��:<���6�KE1j���CE��`SsR�WZ�[ji�f�yV�!t�s��)�T(��*	p43f���S����הx6��*k�*��q�;�g�I�}yK6�r�6��ά��'�����2G���V���)]l�x��݊�Hnm)VR��P����'V�3$�#[�+(����Ck2��{��D�5R
�tr�X �>����4��:tx>o/����Qe�ŰTe<y��pX��5�0�
4��./����4�7�/�+��6���[��SM+����w/2�6ʣKL��>�2ãZ�F"gƲ�.]�X0=�02���Ͱ�u��o�k7�a"�Y9��!p���t�Bv2.P���4�V���#�*4eb�/FI�^��1��f��5�S$cGsE�	
͖�p�S{tu��)�hF�k��)Kh������JF�
�a�.!ݛ&t�����e v"ct�:<@�j�֢lĆ�L�Xv�j�2�i̠#���O4&�NvpF\YBE�����5��ZW'��6Ă��z����F*Y�q�P��C�K��mjF�j7vDi�Y#�N�V�E0	_9��ЀWC�w�ѩ�XwG��]؋Q�#�zb(r��%���f:�Hjf�(-̄�Mز�0')+j�Ʈ���H/�Z�T���me�⬘��*����1˜�Go1��˂b�v��or�� he�A�ŧB�SOO;8w��,����@��?kB�)zP����	nX���fGa�Y��SptE`h#ɹ)RY4u��Wv��g�--���y�􆣡ηat���gU=��ݢ����ޘ�Q�ԶD�R�xN�m�/�UW�}_U}���C�������5O��s��WgVĞ� �²��q�d�L���'K�Y�.cQ�����V���h94�H�_��N��3��������r���i�ᒎ�����=gQ睔0c}���g5%��9���v���J���ϵrB��_�ڝ5�Y����{-��9�z~x���(f��}m��:I�Ĺ��c�i�*ˢ�����F��5�&(wNpv�o+=�p1n�����`���v���u��e��#H��+���]���ݛ�2ڝL4���q��mk����mqK8�@S�φ��=�_[���᷃HN��EG��2u�7v�^ÔV.=�X*�.�#6��rB�0�%oZܡ��ح}���v��6^��È�JB#��mB�G��Z��)@�f��iU��-�[�:8���j_\��ZW��ൢ/��n>�.J�w���t8�Ldλ���;�SR���׸�\�S� X�`�Y��ƻX"��G��b�q�+��'7w�5Vs5���cJ���;�Rp��L �-�2�tPce��CkjZ@a;[��dz��2T9�)ܴ.w1��`�
���_G�ʙɎ�d#Fm�]ʘ$J�:Jȁ۸�K�yFq�N�,ax���/��|nQ)�{9�rb����+�Go��w(.�^�8D��y9��=�Q�k��܆]	�b�gr�fj95
�W��˼d�t��X�"��� ��PL�TT�,�D�5	EUP����4QT=Y5AE$UEU�IUEE!�A@��@L0�UJRR��ET�D�4fT�AI���MT�5UHP�KE4RMIBRD�IACUML�ET�S4U�J��QD��DA��-I2�I@QDIDU��	%�ED���E$4L�AMA�PAU--RP�EQQ4�1	UD4QCIE.Bd��UMSIEU�KK�cD�QM44���a�@�QE90��PQT��D4�aMTUIA4%4��ВUICI��P���þ�<��tWW"�d��m�t̬c( ��y�5�h]h�VT�n��B>����4��8�r+_Jƺ��T+�V��b{������f�}cP1��a��]1:&t�Z�c43I h��%�.�d�T��H�UV�珤ƫ3ݶpe�W�|�,��~��������P�a	疉��t����S�n���=��o��h;�l���B}����o]e�\*���
v�Q�9�n,�ۂ�ծcNT�Y>���+�-��߼��蹮"���I�Ƭ�VX6�"�X1��/O>E{��:�۾��n��^b���:���ϴ���gG�=� 4�մT	M^�XQ�iG|���f� �XaՂ<'M�m�,�/�ua���0Qβ������X��
�N���������cK>��E�C��w6�϶�#](�-��ǳ독ԕb�������5�}�z��\<�����̒���;���x�^�kÄ���j�w��AO=0&��C1��G�6�YA߼�u���>��=C����YC�38���WO$kY�zd�zU���4V�t�Z%@|=k6�2����Nm+>sU�MJ"�ezƿ$0�1�:�M�s9�u2��8)L&<:�+A���]�2�ӷ�&ց�N�
FgJ2�[�)M1�����X�]��pr��e�	6����mkƚ��!u�g]�*��[Jg��K-T5����)�۾������.��]�숩�zy�>�VZ<K*�Um���q�1C�sQ+�Y����T=�G���9�����ֹ����`����+q���h��q�`U�`��:������E5V?�{rG��l;��>8�7����d�A����v�Z�E� �.$3F;��t�o�>���<n�f�	�gP�B�{�Ať�s��k؄.�DH�%���(��]�O�S���r��:KoE�sﲹ'y-��>O/�WLӟ5ç�$��~���X!�:��}�wE��nL{�:��{�I�pP�z�ηJ�zK��IC�����|�L\|dW��ˇ{��職w����L��^S��p�d���P����v/w*�1��Y�X���ȃ���������K?,�6={w���q�yvaxR>,�ċ;�ǯ:��@�o���~sư��iW��UY��8����x���d4Z��Z�~�ѳ��j��M���w��+��:��9]:t�͎���t���
J��O�V7.���K�gQ>�-:��ҵ��z��̡rF�h�{.8�B;@�{;���"n��`��ͨV����B�#S&IY��ޤ*{�v�3�u�u<]���v9LS���`�\/4^N�4��G�S,�4fbݫ]��P]�������p��wc�t��PWɍ�v������R�F�gWb� �u�G�CL�s	^u	�u�;�©�p�׍5�	�=7Mnw��՚�.�˪��~��(q�Z�<vԋ�o����^3��Μ�������r��0��Z�O|^�S��n�O��I_����.:�K��P�Fx��F��w1i��������9Ϸ�u�7����QZ�W�+�&:RXϧ�xa.AB����3����������CΟ\��q��k=�-w5xơ��Xdy����Y�p.9�KG������e�^5�~m����d�
��G�3����v�͍k 6�w�P:�/%"���qw����޻0'�7<�9t��������:�zQ2zv3��fN5ܲa�����!⻷^�Z(�8����^��:Y)S3�Z�9sW�S���Y4�׼�������H�m�BW����}�ڸ9�@�x��xP�����8)����ïD�D��0����Z+���YnI���;����װ�&��H�_��8��o+>�3ڧ�zVu�9f��bG�<e
�L��LI
9Z���P|E�z�s�1ab�B��X�+���*.��7��;�W^8��wy%�m�&\�x��H�E@�,��Ԕ�d�]W@�^��]���ٷ����U�/+C�,= ��������b��,=��R���/�d�7��=�'v��8R�ԦB&����ߍw醑�ғJ��du+3�3b�/��	���R�S��ri�eI=�zwVޕnL�ǎ|�Z�5L
2�U�JE�(��ڦ|�I�/�{sim���9l�]���ޗI_�CȮ�8�4��=�I2����a���~��!���e;��)g[��sٖ'ϦV1�\	�w��yV&׽upb������g�@�/|�5[�I�Zb�mpܭ�<�����(��q�8f'�S,ybY�)�{'L>�g��e�
�V��*�LY�kƖ�
ߊd�Z�s�1���:L��))�t�?>an���=�k}r:ηr��w��K?Vd`�ζ���=	�Zg%׾PfA3Y�j�4��q�����W�0o��ZV2s��9;�Tf�]��e|�`3�9�$�yds����f���{�ᗨ�=��$��30S��x�oW�A��^:��K��}�h��w\���%=���b4�­h4��Hχ���K�XNv���q^��3�VZ���r�����\�v��.�����ӑ��b��+<V�w����P!ú7{]�ͭ��<?p(��}�Zŕ�G��B���`WI��w[��D��.;�GT�Uڒ��J���Jv]Y��t>Q>
�Q���}�j�3�ʁ���nPbqZJ��c�y�0��Bw��������1P���w���w�|�?t�A���^�<Oc��{��k.tz�+�w���;��q����_?W�\�Nֽ�{bS�nî��Ol�v���/�s�s��v�?o������qe�ޝf{|ߜ~�˗�}3��~tB��s�:V�k�����+s{�z&�;-�s^�|g��i߽������.�A�k<it�=ͫ���[Y��#yJ�Z��]c�}��؝ǂ*�I+GK��0J��=}H�]o���}��H���7#ʢ��*}}�T��dy1n�aɻ��rї�|r���Iz����0�P��'����q�ot��{X[Y�Ӻ�6!�j�s����{W��mկ���s��Lt�[���c��뙽8Ã����U�*Mz�ӷ��[���q�fz����6{a^�jG{J�v��.ͼ+�3�t�k��?y巑O��]����igY���#�E�>�u��9��c�-�ir�W[�d�����~�>;��ع�gA=ұLj��P�/�����N�vƓ4D(w�xP��_��U�X���ǕA꿚��JN��i\�Mwp@o������)�*�|���R.�^���g��o_�Ƞ��@����X����{�	���KZ�/]��^�ᵓc�����v�[���^��odֳ�bRw���@w����3W�__
��v�sm�	��N�s�Ǿ��ͭU/pu���:(���k5�+b�m��p-�86s㛙A�6���Ft�� ��.O\^�n}X᣸���^�`%��1�/�+�޹��xD��ic ��;��NV��ӣ����4w��N�}R�hN�u�[���o�Û��R�=^1���'�%��GG0r���K�ey�S��W���4+q�8�����W��t�(J!���U"��S]���N}��d��o�S�}��}�y���fg��uI[R��xۡ	�����N,{�"�ٟ.� ��'�]0}�k�*���	%�傶����֚��7r�W;�%��/#{ބF���i��R����i�+���1�H�}�VEZy�f��{&���*.��آ�������wc���k����b&`H].����I��YP.��W���D��D5�ڬ��C��=��|���܌=����b���ߟ���:�ӛ�V�;ǎ'U�Ok7Tx<�]�jXs#���{�;�;����k:w
�G6�T������=�mV>�<����b[q] N�=��o�>o�����b3����8�D��3�{]s	��ܧ?wuXj9�{�o�����Ў0��6��ԾÎ�ў����Q�Xyܑ�u��>��_Wמܞ�ۃ>ײ��hs��1���͓N�\�O-���~���/v�p�l{'��\��G/s�3dɺ�1�?��f�џ5�ч����x$�s�f�#W�Lxgl�>�r�r���{dyG+),���VlO��T}�y�_��2��j~4-�����cO���w-u��YQs>
o����ϖ�[���}Q�v�v��:�*��Hy�c�Y/]'pc�s���N>��w�������
t��tq����N�t���]e>~��*��[:�9IZ�h�^�ް���{�fQuu�0`pR�e�x�p�SV��Ӥ6|���V4�W�r�)�a8�:�7uZ��R�m��|��$�.�:G3ԝ��.ι�0�����euvGݡ�3OVs}Ӆ�J�JuŶw�I��z	2k�7�N=Ҏ���M{3���U���g���+�mMM����y���8;����'e�q�#)�C��N�>�;]ǭ��[��:�^PJu<z��$Op'�;0wv�mmcֽ�;������5�\��r��?�t~C�]����1���v�w����w�%mp�.����+Y�K�R{�b�e#�u�
�\�d�
�cgr����K�>�����lL�����{)d�i��`���&�r��ݝ����#�0��� wN�	kI���J�W,���jݓ�.�i(�rx��|�C�J�Q_���W�Ae̢L�m�G�$�3�F���Fmg�ڣ��i^<�{��w+\���QlE�&����ٕ��c��eb��|��'��n�O8�9oݏWW}OW����(ej�Oh� ��F_�P�}]��xa�C�.�BLgb��1u��O�%�a�*,�A�ly֑�HjD�e#Lm#֘��/xR�k�vH�!�{rq�Z,
*�.�]��n�:%� L�h�ީV����t��-�
�jr�	F��]˻�?r�^�x�k��P�m%o���w�����cz�bƽ[�z�/}����m�N_�8��29��~���}^�}+�?T�x�c%�h���^�½����z��,���{q��ƌ��i���{�����!��j��5z����ټnXNt����~��]����Z��{ۼ9��2��K	�_�-w�A�͜bL��P�6����=}������N�qן�x��gh}�v��ﵿ|�;+�6w���*�v6���W+�Δ�oo5]{z�H_J;�D-��r��_S��G�,��Kp�}���.�m��[��{�^|&G��L��tB�s�C�S�P����Ot�%�{��c���9��>�;�d���d��`t����Af�"sg��&'�{�a�ñ	����N��ǂ*�I+GK��'f7:|�W,�\ ܉=PBmTYQBL�=�������aV�Ul��D0.�r��xv�5�s�U%�끡�?�����\�Y��bY��04cNB���΁���堭��7CR�)M�R��z�<bS����h��. ;;G^���zw���o�/��U����]�d�6bs��=�������������S��kbO_����'.|��pnW_ۄ���Jo��<��z�Lވ���lݡy�=&����*��k�M�ǝ'���4L�����U���&���U����lkܟ�y��>{��Μ,9�Nt_z�:Ϳ}
��R;�o���ǪZ�I�P�|ֵ�]���e�ly�r[�ߜ�����yk��n���A��f
'0ƽ'w�=~;�6�o�dY4G/s�3y���y��|C��7�����s2V�/<m�޳�5π�Ō�p�8\��t{��=A��z����½'��Ul�p+7_l5�˼���_V��́��s�!��w��~(�d��yc�O����W���%�鎡|�������ᠪ'ۻ��������s��ӏ������>.��s�s���}�ʎ3V�y����}��v�a�:Na�}�A9��13J�F�Bc�_K�BKtM��:��*묭��{�y�����d ��V�]���!B��Ss�P
yۻ��˦*h97P�j�Pͣ�k��o]�p�]����,U��l̤����q�R;���H�kl��R��nvV�ɋ!�wt���)����r����E|J�,�=��)6k���yl,�q*�2�>ѣQ�_ׯI�3�d�=�b<$��v�ת�ʲ�����`]�����e���R�.��I}�7l>m-��U�U��f��b��L\,Nmq�1J���\ǛB�[�v�_�������R����֋�a&2��+:+i:��7a���Saͼ�73OoEb�>yÁ�P�zx�;�M�,\'�9����[]�$�4��e���)hx��	(fV԰�֥PW]�JȥqS\%p�W��0*Y/m�U��e��V6�e\����_b���R��+�Un�C�{Bu��9܆�q�-��L>U�p]�g}�q\&��~Ⱥm��q���+&g@�&��Āe�b�g���r�ÚV:�G �!l��i|���l-�ӽ�ִ3�"��BE�T�p��t��J�Scr�������o)�w0�;����Ou2��w�!Pu����xBpui�M�@�Yk�����I:�� K�4%�^K��L�����+e��;v-nR��fpJ���t�䴷`��ȅ�u��}��E��"!
�ȍm��-���@�Ɂ����|��%��k��+�
T6/:��6���Z�9�W�Yb��
7�^o%�R�ι��ג1��q�or�d��'L�5�P"�xr���25�=����V�	ݧ5.��=�����p���$��%+X��=��6H�A������f�o�B���]�(U�7�hdT+�£�m���g���t]w��랸Oc;�s!��W �L�fV�:֡�p��Z��أ�{�5w�p]x�Ȗ��H%쒞u��XE2%�΅�8e�戱�f�Ҵ719C5�wZnGq���i�ⷵM�*��Ku��&�C��2<%�W6��ݮL]��"ĬS`V�ʕ�/-�-Z��9%H��u��>ѽ���ǰ7WA
�Gd̘w>U˪gRF�����Z�K%��Y[���2����P��T��*t#w��e����A�w�d���O�-�a�2��hR��k�e������n�A�G���MaTխ;,�T���i�Lйc\Ĺ5&U�]0�Υ��o0�}�5�YW��H�YPt�b�'M��mփ.n�5m��󧘸�����8f%i�!W��%h�W��GZ�:�i[E1���q�.�5qN|�z�����˺�v��֋�]��
�yLgoE*hnvʚyf)ڹVo'ĥN�Ygj�̴��+�!�a7�N{��ihݵݓc�uj��K�d3څ���W�c������={�ꨒ����(��
i)�iJj����)Z
B�*�

��!�j�����0��Z"J������	�*�� �Zh�����)�i�����"Jb���	
ZJX��
32��
,̂��)�����j�b)hJ������� hJ0���������*X�(���	���Ɉ���(���(*�2���� ����0
&���)���L����$J��s0���j� �b"
�"�)*��*�"(����3*&���&J�I�j
*3
��(������ *����2�+3b22�������"ih"*�����(���h2
1�02)�ɂJJ"#κ5�s�_>�Ԛ��<���'�;��!��Y��`j���>��)'�Y׻�!���%�j�٭��y�N�`v�s1� �ƌ�z�5������N&����󣣋�:���n�����U��d���:��N~���xl�7����t�"!�[��]ݛ��U�e��c�wW�����^f�T������}X&u��]v��h�������^[t_�(wu����O]�5��9�^��C���Ֆf�9���]^��o����>�y�s����Q��=w���7�z�RƧG�����z�*�����*;'Y���ʺh^߱���6��C���F�;����IlXp=g���v4L�����:as�;���\�gf��}s�F���q���zs����R�3��Iqu��g�Ie��+�2X˔/=������e�p�8�s�螯hp#�F��5���6y�V�P��-оۓ�nu��~��r��g��8s'|߈꽵NU��n�q��Pu�޻�5k�GO(W���~昷$����[�/�T�7��mܖ���!�N���U�>R�)vn/�0�<����b�K���.V�t�Sw�Sg��}�({���;�[����l=_E]3������qΏHt^;8E=�sZkW$��(�<k��{�3I}˸�Q�_�9����:�|�\t/�1c;d�����MF��z��\���O9 ��w=9���fֻ�ڠs�Ey���us��u��<�oމ��NN�tv�3�ӽ�8����2�M2�*��;>�}�4��q��W�SW��Cc��tϋ���s��Y��#���g��&&w؊��|�/�r)�O&�{��L��쪇�h^|B�Q����9�������������U��%O�ڜ����'����0kk�`��חoqwgA�w�5�(r�C�����|yE�g�c'/��)���/\��pnk��3��~vB�ϼ��/y;�l��0���jL{�����sj�s���V�L�,?;%}��Ӫ���|�}~Ƴ#�v�]�s���I�#�
��pV�M�0JvJ�`8�qC_P��4�bC� J+�vrZ��BVfV�њ�w ���:�������,S��Ζ_��r��:b�8�{6b��n��׮QT�w:[���mf+�X���R�DŲoS�vpLL융��<��-��S;���ٺ�P��u.@��_?5�o�UJv���2����>������pz��w�����<��\����"}v}�N�By֒�''��</9�*�18��JΈZX7�rM�>�cv����v���t�Ԏ����L��ޗ�U����e��\�����pF1U��v�WG��Gʜ��ǫ�}kj�Y��q��������{�=׿mw��_�+~��WÕ�o�@�D}�0���o's&���z'�s��r��G��?F��|l��;h/j��5�ԇ�-m�u-���g��*������N\;9�۾�X���y�^m�}�{�>N��C���f�7�8�i����He�[˶6��oO:�G��|y2vuA�͜bL��Tɲ+��'���̈́u{5��zN�����:;GŊ;��w�������{�9���f]���%�؂�#�,zm�/�`p��x�g����9{�m��Z���[ub٢��/�R�K�/x��-ɉ_R������3z������Ƭu�V�<OB��ͻe��=���*2jZ�gT�r�q�w�����0;k�Vw�+����W�GY��g��l����/�Yֈ�7�u��t/��Y��7��y�λ�m)�}���_>���t׏���o����4��F�Ţ�^�ɼ�އR����9�;��/��gx	���d��dx��N���~���{.b(��Ok��^q�z�y�}w��$�%�-�v�ޜ�^V�s��u9�0���,��ʺ{@f��ﵗw��/�2<���z��O<TU\��e��1wm����z==�����|�^~�仔���a�]�����z�~��J�2N����Ͼ�����~��gӷϿ#�?���hd����������>�	Cܻ���w'��z\���O�Z^w�d��w�bu.�?]�;�p��<߿���V=�^�����i��P�>e2�w��R�����AHto���>�A��4%����+�|��.]���#�伎�br����￺�ܳMw�_�7]��|�Z�g������!��~��|{��R�
�x/�r�ގAH��Ò�2����w��w�i%�^�{װ������Z��wR�\�����}�̕�Z_��������}���:���}���^M��Z_`伂�}�B� �9�<��}����仌����%����;��}!��6�����(~h�
C2V�Ln�|s�[��#�\5b��
�
�sM֎��Vu��0f���H2�a��a��A��r��1����z3��d�^y����������WK�󐧯�A)��]K��dP�e�{��,��V�
J��,�������}+7:W<�]�����u/����C�_c�X���z����>u��y��A�w/�i}�r�2{���yZޞGR�Og>��w{#��}���<�w�]��z�~��g�{��|�}����/%|�5֗%�C��?Y�w=�#������&G�`n
WC��A�y/Ghh��?"0l�>�}��5�z�i,�~���>��ٮ�_d��r��G�=����_�w{���'�����y&��X���]�F�ԯ�r:?`n
G��u��~!��{�\��u]<�5��ď�����ߺR��?o�9}�-��>�/���֕��^�֗r?GZ�K��	��'%����C�9.�Xj_��z��T�����y�����:Ys��lԯw}��_�$:<ރ���p=�)K�7��}{���sH}n���֑��/\�I�������	ۘ� ��B?
�s��~������[��n����z��Wp�?u��~��ӯ��w����r�^y�������^��]��r���۾h]�R����|>�~=�p�9�|E�_�Y�I��������)?9�nC���;��>�Ws���K��KxH�{�~��|�����Od?s����?=����+�nVN̛�u_���}��ex�ނ����C�P>ۇ%�d��;���ш�_c�^�9js��7&���>�J�nk��#�?o��U�����.�}����G̀?k��?d�M=��<����)]���Z\���7&K�d����%���Gr����{jK�;7�2���?~���?Η�����2�7�a�}G������9+�g3G�w��J��;�)�<��a�^C�����]>���~���X���y���)�<�����fy�Ѳ�G}�S�]����In��8&L���P�9Zr"I�Y�8moR�.�>�&��=��R\x���T���51�ѽ뱜��d����s�S��)	z�ib�F�K�.ǉ������ؖ��z�Iך�q�c��u�O��;/�_W��}X�=�����Y���}�����[��:=�%u'��h䜑��?��'����ܾ�OO7�2!�o�?�w_w���]�{���|@���_��R�{3ӱ�����Q�}Ǹ�M��:�Ow��'!�ߴ��Լ��ߵ�]FI��z9+����w	Ѿi���d���	C�?�:�����|� o�9���q'����z�o�\����ZN���sX�J�yw�Ի���z<�K�;����Ի��=ޅ�I׻��)\��{��~��O�?~�HG�߯��$Oِz*t6ﯯ>�]��׾��>������ם�r�e�w�G��z��`nG��u�'RnG�_h�:���{��R��z�}��?�~�?����7h٦��j��{�^wןlԽ�Jp��rr_oa�{����}߿��C��,�����b>܇���;��2?brM��:��~�pP�����Yy��o����w~���>�_u���}��8k�OP�A����w�#��4n^K��|�C�.u������K�M���N��y�w+����	}�<�~���\�'8���8|g]��(?C�;�IC�FO��w �u���y'y��K��{��=�/�^iw+�Ӯ��/$?��K��F�O'����w��kλ�����^�kg������}d�@2#��P}/ђ���仌����(A��ϱ^I�oG%��?K�>�����o�.�w=k�.I�{��h��|�����w�?{�o�p7.��xk���22�}>�7�~���M˸��7��似��9�)y;Ǟ�?�������.��^^��~:�f��~��Ϻ�[�o�=����prWqοirO�?���y'�0O`�]�FH����O�_�������S�ރ�w// ��iJF�ח��/P��a�w�u��w��Q�?�0�}s�����j��M?wx�")ٽ�]7�z̙��^�2�C��f��{&���Sy���Ό^+zCޔi�mʾǦ����b��O3õ�p���ɼ� �oA�ar�`�7y�0r�.YYV����IIi�St��G�rom����߾������ޓ��;�����~����G��.���_#���� �}���wy��;��ѣ��P}:���������7�� C��������U�r���wa~��%�/7潾��z��b�9/P�|s�#��.�ƕ��K�P:Oq�����u�}&��0��#ν�}Kﾇ���;���t�!�����(��{�K��=���^��?h�^�~��r^�����~��_�@����z
p~����]{��%�2_Ɛ������?�λGT��;Ƿ�y��T��]G��{�G�tw�	���O�i�Ww �\��<��|���O$;w�'�}�����=��w��y�!�?#����wL�����zOve���D9.��2��_�ѩ�8u�y/ ��L�/�6y�?+��?sO$��a�w	�����`���G������ǽ���e�!:7�w�ޫ�R������4��]�~��=�������w)��w��.���C��I�~�!u9�ߺy4���������S�ّ*�B_��~d⟾���%�d>�JRy.�a��v}ޗ;�w�˸y�7+��tw�Ի���w���ɸ|}�H{K�;=�~?�7�����.�k���;_洞�ϻ�����������2N�愤�_�u�%y/I�z\������y/QѬM��r:��w#��GR�M����#��3_��}��{�k����������=�����R>�^oO!��A�4����_|����u���_|���}��Ӭ��z��c��w��4��Lg~*��6 �����jOdxu��R�/o�h`�A]���w$���r:��y�y�%6�����{���y'���K����}���C�*��WeM�΅M����7!���냦���A���ߓ+��,��U�f:������k�٦�vDcU4�M�u�����+9����6�.�EmGʛ
b���pSǂ��9�u<E�չ�V����N��z{�hɃz�D;�UU_}�����߳_l���F���X���~z��i]~��}/ ����������ZGrrN�oG#�I�}����#۾hܼ�w��ך]��zy�������u��u޼���K�C�������%<�K����~�#�X������A�y	�ؔ;�q�����5���䝙��~b<��Շ�����w�p������5���zߛ��y}/��Z]���]hra)<��rr5�}'�w=k5+���br
G����Mù�7�C�y��sJR�Ou՛��}Շ���9ߙ�������5u+�9�hm��=��Y��zy֓%}���irOa?f'���
O�`���w=�R?C������+�ѯ���s�׼�9����u�mg�����~�p~���x����_|	 n��^�K�z����o����d���y�!}��&���>�%���0O`ܼ����np�����k7���}�>��������u���[�r_|�;sz�ܿ^A���r_�zy揭�ܽK���<��ܝG|�H�K��rGpoX��}K��{����5ֳ��W��ͽ����~ aQ��!��iM��=�+�p;ޓr��S�9�r��I�a�^�|7��\��~��X����'Q�;Ҝ��zyނ���ۙ��͕ۘs��|`{���" }�Z�>D}��?��}%��~�w/���t�+���S/e�{�;��;y�GRrW}�4���=���4����
m��o�U�~��+=?>;1���}DGۈ~���#!x{�C��9/�X;��y~�������z����O�w�2ܽA��~��rM���.���Y�\���������wk]���5/sBp=�IA�}����hA��G�^I����d�/�ش�w�~���_/�_�9.�?�����ܞ{���y/pg�{�>��?o�C7Աn�~$~ut���:�Uz������ S�������^�x��]rn��,}a�:x�O���Ť��Hc��c^�
�L�� ��̮���}RD;�_�G=uo"ܝϳ�|:jg���>�(�r��Om1-튋���`�R��Q3���������~���WQ�u�C���ގ���N���ܾ�I��4%���Z?J�N����ܮ�}���C ܯ��O��S7�����F�l���o�v쀮�o��>d}�}�����pv{��#��^�G �r;���)w�p�g ��%����+�~��.]���G��yy~�޹޵�+vq8fjs������W����_ߩ
�S�w���_��>��=���߻о��:Ow��R>�כ��w��4���r��!����z��|��i����M���[^�h����B?
_w��'�>G�����}���]���Z_`伂�=�B� ����:��{|ގK�����������-n�aiݮ�k7�Na�u�歹���y�z�:������K��X����GF�䯑���C���K�)|;�K����߽h��3x�?J��ϯ��83��O�V�O�Q��W/���L7/%߸>sK�_.�u��z����C��Z�|���:u��~�#�7+���A�y/`���Gz�?o��߲W�����?�}�}���[C�]�ۛ��wy#�=������K�.�u��=���NK�7Jy�q�ԯ�r5�~�>}p���0���>���g~��2��y������9�JR�No_B�O�ޞI��w/�ϭ+���s�.�~��u��}����仚و{%�k=���������{̵�}��_ ���ԯ�oA�w!כ�w�y���Ҕ�����}{����!��{���֑��/G:�d�����.C�&���Y��{'����ҵ������ ����tK��ъ������+�־�r]�J[��]���>=��}���/R���/�������\����`ou�p/����2���*��KO��t���Da�jV~��F����M��=�;]�~�~�+�g��8�3�]-ɏym�G�yφF:�,BѨ�tg�8ob��]��p�Q1RE�s��
Y][�'e�R��u�Ǟ���ﾯ���ώ��������?�>D@����@�y'�0ø~��`�C���b}��������쥼�z�����y/�=��[��>��矵a�z[���s�o��������_��q����^�ނ������({��%�d��X���	��~���w;�zMɫ��ߏ�������c�?~{��d�ok����^����������>懓ԿM=��<���z
Wpo�.FH��%�2_M`�����b;��=��ƈ����@3v�7����n�f7>���{��~�䎧ro�u'%w�3G�w��撃���N��r%��z?J��ޗ#!t���~����}�������Պg�x�������u�x����wy�2�=I��䮣$�����?�����;����4���)���&C�?����.��������C&��ϸ��*ɿ�;Xǳ�ir�%�G��y'��S�]���^��>��>�����k��������)\��y�7�z��|��c�C�H����^��+��]Y�����q�G�{�.�|��ZN�%�:�'%{����:�r���G��{�rx{ސ�z�s]���������G��_�uп�����->�#ޘ�-����?�{.�$���%�{߿�ܽ>w�˸}��٬G��z��`nG��t��ԛ��}���^C�|{��W�~ vX�� ~?��߭n<_����7��5����r�2S��h;���{�7�=��z~����!���K�]�F�nC��k����9&�����  ���˝C����}���>������#�?A���rz���oG%߸�o�ѹy.�a��C�.�w��{����Rn5�y?���e/��ﴄG�����w_���?�U�n�ż_T ��A���Oi��Z��+6*�;2Ƅ������ǚ5+�%]�.ˈr�qIK#t��������3uܹOWU�~�`lsQ��[�.��li�]�Nf��TđT�a>�dky�5)�r����s�ДV9�i`�ɻ�t�x�J���l���6�7����*�:#Jࡽ�����=R�.`;ف��. �b���ԙ":7M��tNr��t� W m�X4��ˆ*�w���o*��X�vq�N�x57I��C�`S�F<6���s>30U�˦�hEK�[�K޳B����kU�M��M���)����k�����E���Q���	@�������4�˹���'��f$!��[��JJ#w�^FX`(�UD+hD�2qJDf�A�wBP�|
��ֶ	�A�;�Yɪ0L��A�K)5X���WrH�uLO�-���߯_�Zd���u��NoV��vL�9���:�IKܔp<)
[��[�e�'�3wx�.���[r�{l2��Q���m�����AMG��>����N5*^�N�B��'fu!j�>̤�Cb+r�����Y�ʙ��`�&�Z��yW�"W{#��vWf�[NF-vC��-��`[����o�����j���8ڑ 0-�*�H��R�.�����[ܱw5��B쬮��7�e��_8G]zӵ3&&�d�>��9'u���[�k6<Ė-أb�Rw�V��>�U�)[D]�^�sH�j�^�5���Rn8��+Cj6�����&�fݍ�R����]�oPٛ<�*s�#�#_:t�-\Yb�ʶ(���.�:�s{� �맕���|�t��u-z�<_mV�^Dx���
+:��xn�����tc���8`yv��t2�i��Ƭ弖'����a7��dF��-Nr�99�L�Ɩa(�b�)\�{r:ˡ��E��o��CL����w��t����7}��l���U&��0���Y�y3^�}��J{RX�dd��a糥���{܀���(^��f�}��s\�@��X:��Zͮh�˱��0S�����^bdV�ӷ:V�J��WeTWX�q=�r��E�>U����x(�Zlܲ�m��ǎDѝ��Cլ6�0��1^����(<8�o�H�|��wW8�.2^h7��šT �M�ۣ�*����*��V\/8��5�m��|y�^�0�*�ꦴ�}K�b=<*����ÁC��ds�8�N��)�$ʷyǁ�l�ggz��c�,S�J�lUc��f`�kYeţ��'݇p�2ԉ�ځ�T3�������{0���B�[�yB��1�'	�*-��
6��}�Y�ԯ��l�7�VK������/uon��-Fc Q��\x��,ϛ]���R�˛4�'h7VT��£��es���	���[��Y�,	<���B�S4t
�]��JҚ�%����9��E�3���7�����F>ڎ�b�Xު>����h��h�2
����,�)��(32����������H��������*h���2������&J*���$�*�
(((�Z�**(������2"j���b

�*����
�iJ����� 
��
))"*j*��(�1`�)�&�

Z
�%����h�*�h�����
���JH*�*���B�� ���r�*���`��&�&�*&�&��
����������0f&	���>������y�z���O��&N�8����gs�3c���kݫ�W�H�u�6;"S+s�Y{E�4,�9�N����~������~���?s����&����uA�>�@t��IC�����7�w �[���G�_a�~���3�������.�|��Z\����=���;����ֽ�}��wvw������z�yߞqOgR��jW�9=~��
G�uA�������&��d�w�	@r�7��b���7�������+��?�K��z�ޏ�g�M��7��>�zqo��#�����H�d�C��X'�~����_`��F�~�5��r�2C���i9// ��R��~�zy�#�^o ��^�����x~>����|��}�����⻷7և%}����{)�a�2�I�0O`伎���~�q����/�N��r]��w��w.�����n��^��Y}���_�������?}���9�������h:#x����t/��隅��f�o���.�m��]�'<�$�ɝn����uބ�t�R|	6�-���ۥFGLs��I�J��e{~�_V	��L�/8h=3��\Wm���������}��q۱��3�.8Wf�h��ۘ"7�t�Q�rV{.7� ]�d�7g�Ԧ�o�F]1���$p�4h�0"T��1�
��s�ܮX���S�r��G��eV��''��</+��i�W=X�7k�3M�;�G��������63n���>���g��}���!׃S�җ/r��u� ��lL������_n-�,��[sm��B�0�yY�+R�I{{�p����X�5ml-9/���5�����n�OW�R�'h�a��] n�^t�!Lo�x��y�g#���گ����������x�X?��4�c��;;��O=�����=�57ڷ���
{�.z�q����Μl9�N�hz�/����.��u���J�sɼ®�޽��r[ߥ�ߜg%�{C��ٲ����ޢO��W?M��◓��$���oL��=�ik���i���7���|-�w�����TW{t�it������t5{(�:�Vњ��s�N\ϏN�{G�OO���Λ7k��+g���N6�V���ټnZs��*��͓��u39�o˳�׶ӛa�KVv����v�˨:��7�$������H$�{X�;;�����%�h�����5q>�R�'�]��&�~�c;2_�.5�>�ex�ןL���%��Do��*�a7��ql�/7Im�u�v�?o���:{��	���λ���㭢��2S��TBm�\�[�ƌwW�F����A[�h����S����Zɉ�fӼ����WDQ8ʗz��ݻ����6*J��N}akȥ�Ӈ����-=���o�ڷ�#����+!�}W���F����u}��/�\8��|�\�߾����U���R���e�'�hwP��7=�ǝ��-��ޙ/�\�m?&_�ޛ훯�Q�淇�����h&����ٱ<�wzoݛ����T�������G�����,��et˳-]��՜�..n��fi8����t�N�]1o��V��:�&ܺ�8u��Z*<��y^�z�r�}�}Ux�w�����d�,|�zltt�vv4L.�>;~��X�ܗ7=��ǲ�\���k�7�psCcӾ��{}�t;/[���1�<��:��Y�s/j���6����k�o�3y1���o�cK��7����[}'�&����2�_����cߝ�/py�Ny��W����BWkOk�	+a�t?�	�}��m�t�P<���ק����m��\��q�I����i�^�i�a
� �]�/U(Ǔ�e9oM���Y�i�W\]�6���%�!�|w�η���� ��Q�b��3�65����_N�bU�٨��pZ�����p6�nN�gO<������a@3*b�=�u�+L��N��-*���{[��]My�}���}�ِ�{���Ǟ����{݀Vs���������C���xqf�^�R��#�]N����N>��[�Gs���^��;��Â%����E��o�~r��=�`�&v��'<�8��,�󫵆+�D���o�J�c�>�8(���{��56x�^�����C����g1�ԩ���v����a�腰�_|jyl���<�[��Y������/\u^�/����hx �5�k�ψ{�bx���MA�:�����VyU�K�@$��%�_��앬��U�OnU�y[�N��ǻܴQh��\���o{#�<p/�beKxJ�b�Om��X�+�t��yj�����U�~ݤ�/+��r[�3��7MV�8|�]���O�3�9>����v�w���*ro��Dk�Q�-�zmS���B�Zxk�un��dT�I5*���tK5حX珄<+w95>3�뮗&��b�	������ di�%��m��в��3�bR��W"ٻru�ӝ��F]�;�NU��l�\�����AD5�j�M���j�rѧ�9�߫�����$��Rz������l�i�]���;�U�x�nm��^�p�{�2�ͷG/w�����^���_�����+ts���϶=�����/�B�i[/��v�C�sYS�{Y2n�=���X�-�a?zo�	���Iowocb�A�9��p�Y�{��=��\Ù�?/T���ޙb��TIƈK���*SU������d�zw����~~4c�3�:��e?`I�w�]4�qW>[R�Ju�LV��l�bG:w���sg�j��[r���w4�>Vz�3�u;	kQw�\ٱ�$�z	���Y^$t���L �_�P��#��Y������Z\�����t~���X#�[/%k��'���5��b�����/��h��,P<�ξ��O�WM���f9ʘ��p�g��;v}�闓:��u�vF�>9!���V���kܲ�L��eM�Z�/���;���:;��V�;`�=�M�Y��=�_^m���d@DTwv*P�`����e�����z��̥�C�Ae�XEK},����3���ɻ9޷S�
[�dr�4d&�q22�0�{��o/}����z{g�]/υ��ry{��I璯;"��$��.V�07D���Z��/T��=��c؊1M�b������v���Q�U�Ϝ���}+���ɇcq�֧5�*�w���ʺj��'�������¸Xj��_�>�g�#�~��b��;�v�h�^߽�GW��/��&�������[{3_y�z5�)O�:��ރΔ�6�G�_���Oמ��$�6���J''�nU����U�����s���N}�m}����;���y6(n���TT��s]��+]l���w��\6�/�����3y1��9�`vl�x쪓�E,�U1<}�W�н��pg޽�g�nX	���7�G;}o۽�n+��_t�3=pk7=��`/u�]�@\�1ᝮ�r�r�|zw�e��=ԵҒs���x��%�x�����V�hp�86l}���)$����-�R�-Wʕ��;P�[U��GۯW}��;�}���hh���t��/�vY����x��m���L�'1���L<��@l=D�<,��ᝫ���F��
�d.�8��k��L�E\��_u_|�>�q	���Ʉ*��ʻ���������Y�'y����=�	�7���gh��.�a-�Pu��̴AP���]�dq5��ǯ ��2l{x�u�gk�Gh��@�v�ۅ�w�^G���çoZȷ�ߞ9��$��|&oc��m��ˠ��i-���w^���|*J�����x���\�Os�ɑ��λ׵~;���Ls�v�3�"ㄹ�C��'m�@c�����I��K�G�b�����]�Lv�R��>ˡ�j�O���؝��v^�}*㹺����7�jI���Ov�)8(��]�{k�]�o��=�b��ٹ��k.룭��(�j��޻�o�����ELXpv��m�.����r�e���\X�*�/�ⷝ��=޾ٯ�`ވ���KbÁ��3�;�vv4L��A.����$�i��Ͻu�}y��{j1�8޸9�\ǧ>�6����3xG/$Uj�}�v;�;l3� {:��S$o��ֶ����v�s�y+��Uͻ�4I}9���c��Vlý2�(�4�"ޛ�&�3;zQը�'h�[kI�N񸮯{m��'Ƿ�&+�t�Er�د�=�:=��,��������oF���e�>��go.�^S��sm�~�5��q�ɏJ�.��;���͏�B���#�j�+tw����_m��ײ��W��R��'��q��V=O�ߚ��V�{ń��t����&v�t��~ڵX�#��v��E�~��=�Gԙ�+7�S8��ƭ�wX<}�57W���f�J�g
�p�7��:`.?`�o{���f���/S�z�5[so����Z��{+�[l�2	QΘ�߾�}�-��;�5�y�O�S3��Μs_n8��]k�7�o�	U�o�;z�/�����Kq�`^-H�tYp]��zZ�_WZ����s�ٴoe�t��[��^��e�w�����e	D/��>#�q|�M����u�~^U�f��n<��ޮO���}X&u�x;!k0���=��ޡ��u�z�nVV�os*��bBW�}n�]pXlI�n�����Fì�j���e�i�E��������2uz���G�y�A5��c����-��j�o�ؾ�s#)���3\Ɖs�8�7-��l&��v����ʼ������ow9E{;�n~�5��fW�I/�K���ӲP�x��Φ�{z���;ǹ�7[Ԡ�[3���ږ��*~Ϝ�ܛs*[�i�_��Y�.�H���ͬ�ר��~����$��ذ�z#9���UV)X�(��!%nL�:��^l������9����c��Q�7���y�,�^l�={�o�������m:+�C�ӽ�{yj���,�����w/::�񶁟vt6#ǧ�{~��~Ú�g��{,e��������sfz8M{����u�/s�?ps�ٗ��5�[2�]����
퐊5���ɩ-kk�xL{�fۖr��ǹ������0�qN�(\���O���`��S���B����p�SOH�w�ϰ�o=S�:n�C$Ca�\�G��jl4ϖ���TV�����&�:g���unT��Z��-f_W��Ո��0����Ô��,sčdb�25�lJغ3��ziQ��?f��y�==ຮ��y.MC���ws�Os��e!��ܱ���)v�k����=�P��E�gj�w��2��(����2$d�-mΛ�M���ߪ�������t�����k��ghv�����WX\ٱ�$����s��b�n�]�y'Ӟ����Ǧu�;_:;_,Pd��]�Y2\���}��};G);�^�����v^8���v���b�<��&;�|�D�zx��v�~�����?{�痓$˗կ�����'F�l�v>Bw7���z��֬�p\���)<�U�`�^��K��2]���V�^VƗOyٗ�o���2`�4�u'��7�qۿ���+q����F�5�ު��ܶc]�φ���l��ׁ=�t���<#.�{b5��#�}{瞭��ʪ�sX=��F=N����&R{��Qм(�rx�����[�,.�����;��§ыp==x;�}��\ߩ��C�pR�F�Sb��������;�5�7��}�qrߏA����Î�=p}��.�w�Ϋb��26�)�1ڭ�|]�w��@���f��s�ڱ;��.K�M1�U<��
�f.]d�۵.Pݢ�-6��t��9��]�A�(�î>[z�P5��C�X�]ޝFklv42�[�k t*��|�s���)b�w���EڤҜ��K�;@a�-Vձg���A��2D�aMW�^cn���ԧ�ё����{��V���Z�9j� ��t�7 H���`n,�1۠�������=@[����}XC��o&�]+}�y�Nc��NR=JC`-�b��r�l��"oBwz���Իj7(VYx�\;]ܹԵB��V��l�+�����  i�r��3�����m�����O�,,�3F�%W����G`��;V�8`8g}�����֭��*�`��K|��-m�1���N�����A�X�m��1M	�Ay��`;YZ��(哎hM����'҃�C])\oA���������U]�fJ�i�K ��%,N���K�j��B�8�����ɜ�pI9
ZAѣ����v{]{{xZ��*XMh+wkX�V�f�%f'��4�Kt��L�˂س�Њ�ym��	A1�L��d-�uҝ�r����g����Ïi��v�Ra�ƅ�������oc��N��IU�V�Y�T�ʇ`-+z��Z��ԭ�]�mɉ���v�TJ��ۇ�B���F �j#A�Z�q��ҭ�����4�J|˹�9�ᣝ%�;���k��<��W������w�d^�� m'Y�h�uv/z�_S�5um'Y'�;~y��K��7�vX<$Ɩ�zZD:��W�UY�>���ʄYhY	���^��V�M�B-��X�!t��ϵ!�֌'�@���%�����'Do�$�i�gt<옣*XҲ�Z]u�t+��4eu�ci�@s	�����cѦ"�q�Xn��@L�,Մ�A�h�5�eU8�N�i�yS�5�ۗZ,��U��[,W]��gRw֬��'a��t88��ˋ:��V��̂��1;�R��-_^���J���pN��ӷ����ӱ�s��R�����\k�&�<.(r�J߳ƵN�|��U`���/��E����r���RKK���
Vs9q57�4���\-���fV�Jֻ����꺝f�殷:�碳���c�Pf=�O����zڶ7>�s��F�7�s�c,|�mt|��
�놧Vc��[{K��,�:�V�C�W.�ղi ��&�.W��S)���3;6m�� �-�W��b��e�,ۥz�X�U���gs�LZT��GMvրyt�Y�TL�.��L;�K��o�G[���fV�F�I�QN��r9�i,[ƺ�����n�5�g:��}o�W�Շ���q&�td��P����q�˒�Cz������/��מu��1DSTRRQDAT$TQCDT�a��SS���UT!ITP�PAa��EEM4�U%L�5MRT�%Q���4UEUA@T�UE)AS%5%����1��
����&"��ek+$*�����
J��'0r��*�3������2�30�
30,���
��),�& �:��Ĝ���3,"���2�*�������l#*�Ȥ�0��1ֲj`�%�E��U97!��:�L'psL��͎�o�U���;�c���[�����q���v��@�<D��d}�N��/���}�|f/t�{�b+���VOFf��ߥ���q����=�~�'���u�#�:�f�qO]��5���}��}����r��8��s�帳�A?U\�~��s'Tk���������+����[Fk�6ܴ�������iҢZ�������̓�Ǿ��qa�ƙ�q�l!Z7�8
Fk�+����L�y�"�s<�4����j����S��]A˄���i4}W�7Eo������bP�6`/{�=3�Y֎�Ŋc��7�������';�0B�a�\N��\��%�z�����}r�Ӣ;j������;����%o�̲�|�!�W��t~�����u��yr��w�YC�W��^�=�:sӳ��>���0�M���J����nnv:���gk��9���2�N��N
o���5�]�A����WOk6'�vv��)Е��<y�h��ݠ&�s�y��;;���$��G�K�%+��в���yW�O-z�xn(��d���wn��v$��m��K��ۑNHӌ�<��yh��J<|Űj�vn#ϴ����)�mJ�Cꝵ�ε6��P2��-��k��+�W��.��些~�^��r��:K�K��'����Ɠ�WOsoc�n1Yg�{����x���st���'ȁ"�-��$��u-�2��O}^n�o���G1�Js��7y{n��z#�c��Ka��s�{���ߡ��g��R^F�|�vwh~>�t�8=r������3���Ƹc�7�y٩�h��n���|���'���R6^�4x���f����ޢ�������y.�ڭ>\�/D�F��\�z��(?J2�=~G������ީ��O�hI�s�xt=˻�|�_����y=��	+V˰��rW�^��S�/��;q�l��{�3m�	��	��z8�����f�x�>S�>*{La�u��.΃����1���ܴ�@��{ܯ����3n�;�x]%7}Rd���Uϒ�V�|��$3 ����q�\�����g�z�(��MX��i׳>-�Ϩؾ���;n�E���*H3�Q�h&D��ʹI�Z����%yhT��ow��EK\�R76M�-1p��}��MI^5n���7�/�H �h�jQ�f��׍���7��I���9����}�j����ų����_�����{�͛��$݂?�v��9��B��=���һ��'�X��צ[����n_�s������{�6��ӱ�ot����\���U�79���_J!��.���쭓�,��㴭Q}�˻�\��7�}2_^}3��~�_k0�}�����F�]�+w�������&�
^v|ԿI+D��L��P�{��
(]?K�����*�9Y5t�<�]�j[�?c��9=�*}3��Qm?a�$ٳ^@�u�+e���R��އ�]�lF�IRSC���ĝ��nt���;��u�f熎�R��Iy~��{�oD{�8�W�c$L��ە^��X=��`�o�L����~��]6/=1���"��}U�O3'.z�t^����=/����'��-�}zq�~�;��~5>ꝿy�*�&s��_��^��W2�`�H��k�0=���%� ��t-7������lxN�_	t�2<���Mܷ������[ׇ��&̛|�9�N��!���)�.�T��h���5ݼw�*�v�e� ����+�ϴ�?UU}_R]9�w�d}���W�z��9{��3c&M�G�c�}c�xӰ�^��V�E����OIӫcI�oM�	H���99~�??G����9�{G�*�w7c:띗�7P-�wƸmh�^ppߛ�ʛ���q�v���̤�:�g���K��2�k5N,r�]\�Gh�u�<���+��s����]��&�؟Ggd��+:<d<��ة]asf�a8N�G�q���b*������m�f|�Ҏ��GG3��r��9��c�����9��_V��{��w����v[��	�h:!}�X�yϷ�����O���k���Pt�N~�qs��]�r<�}Z�:�c�ψ�ҧ�Vds���ǲ�3��-׼����)<�J��e{d����VP�Jҹ��- (�j��:� f��R{�by�k}��|�ǂ*��{�ns��n��P:�M��p���S��_-�j�;�j��bs�)�����ejI���U��-���ʕ
�{K������'���@N&�8��B��@�|7�)�Z3{��T��%�cY��b\h�v��9/5�<�Γ�5�P=߾���.7�yǑu.�Z�ƽ��z�^�Ru��te��b3�f
)W�~��}�}^�U��h���|���x��Q�=�uoS5��0��oq�s�*�o���m{���龃�Ժ��k�}�g�Ȑ��uHe�n�uW���y��T�s�����a�zz5��U���눮n���>��tl2em^T}����M�����c��{A{�nzg���4y��<������qо�cղ�ۖ��3�]�t��ε<���!+��֛5�k)+�az]���}l!Z#���m���7�+��ѵ}�wm��k:�=�G������wv�XS�a
���zͅc���߽���L�7��a�gG':`.?dӛu�gG�~��Kg�4C/]�wI�,mZ�u�/V��WWy��x�����zg\���|X����eQ��V�G�a8EЭ�1��+n���i��F_
ѠP2����{��l
����a�f_Mt���E:����[�����|��s+D��F�����7���nq�fZP�����FZ���|�FEC���o�����C����f��W�',VԿ�6o�<s|6	Bf󼙽��%�~�X,2{�}��K��9^�͑>�8+㳬!΅�;��=�ޛ�8�q��#���wR~۹z�gN�(u�����!үy;���W��rz3v�=n�G�O&�c���^��k�+���W/��9�B;�Ms��;L��u*W�KB��);A��t�Ox��n�:y&��x������x��D[`x�)�y`:�f?|��S�҃��������v�˳�C�F�}1>�%�o�~O���$��w=W+��嚰����9��ΦEX�1��-j��t�˸{�z�yK���[}�/���#f������\.]�X�CiB���\࠸zX�l9X֥ݑ�>Ѽ�}�I�m�:�W��f��=+�^t|�\LpT���>��8��X%��a:yR�R7��Y^u^�� 9{��n����	���k^	�&	��Ӽ4׏��χ�n��2M��X�f%x^������9��F��ԫ��ml�G��u �o�Q bKh�����1LV%�a"�(���{oD�'V<�{/�}��U�n�p�F�:#k[��w�ל�>3i���W}*J]ʸ��c�ø��Ur���T�_W�}Y�9��{O7����m��OqW��_og����tՖ�E{Rƫbz	9}��vg1U��W)����b��z'���F�������Ƭ�[jv�W�j�r�ۑ�yv�ׇ�K����M&GE)��|����yv]�!ث7�]���s�8������oݪ�J�7}UP��Kю�&��
�J1\S����=��]�qT��c�m{���r�T�%�����\^�e��D�l����l�e�=��r�{���_,�}
O�}�
��%�b1�o*m�wA.I�a-j`�\]���3�����z��>�2�^�浀�S���������ya�����KH�T��� 5�\�?eeOi�]�ŞW�R{��S: O�<�%X��~����g����'��e�OD�;�_{'�s����G���jZ���2:�pjc*,1����jr��(V-��.�p��<*a�h�uvc��9~A�Oۙ���ꤠ�J�㵛�!z�5luTW����x��/r����+�/I�Hn��g�������ꦶ�*חnU]��:���a�]��U��]�t�RU�6:o�T{�	��H�`Η}���(H�t�m�c��q+��Nd�݋�)[GPsuo5S���V��
��?+o.�`�׺�ً��wE��;?}�}�S-IS��yg��I*���J."���;k؛�QYcz]%mCX�1��˞�λ{C\����G?y]ת�}F`Cx���U�8�৕�R�{�h^V{�΃ܮ-�TE��٭~/�iI�=}��{����^�| ��?�'^�lٮ�����L�|*}E=��O)Xt�ߕ3�I�Ļ�E�:]�wF���D�������s]xK�o]%xd�.�q��>}�|�`Z�K]֡>�0q�ܮ��,lY����yo�GY��^�@�Z@`�2n(��ec�q]^�wv�'��ꚸN��:�qg�vYNf��^��w�s�=��ͧ��S%�Ε�2�dQ�Z��%a�V�
��/x���U|�L���9O�msc6�u�c�֞p�-�3�ƫ�׈�*+��M�h�`��H��"O����$�t�����d⷟y��C�&�:#5�dʆ+��(C�u'b�uR�Yi5�n�{�]5���i�A�	v��4l����>5ɔ�X�h񰙨��K	�T��nt�J���h��y��O������;x�%
o�5]�I�6����ߥ��f�DS��^.�T�M�SS9[غ�ژ�n��x3���Q6�����[�E󵵥�׈U�����Q=.�����P���4wF���/'ul)��.���&2�m���W�W�5C%{��5M
�sb�7��~7u���,�S����rz��r�C�(�ގk�<sZG'�kN�'>���ڳF ��ki���&� �y�i�8I�=��%B�5<�:��tWf��K�\w�<� o�Ē��AAB/yPe����3�R^_��J+՟IS��w�����?^g�j�ms��xP��e��t�J��<�7����2��=����s��w�ݛ����;��:J^GP��(GђiVp[f|�h�߂��a�q<״я���3c��̷���G|��Ur&>G��PuD3vAފ�H�Y�.�C��:������[��yڧ:df}�0R�� 4a���
z�J'Ɗ0��Y�O-,�s�N�h��JrXR��E8W���O�����[Ciw�%�,,�ΘN��p��5r-�����-�ֲ<\�ù����eCy�̆o��x�>�"����i1�^��l�<;J�+����ܿU#���
���MyX3ˆT8*���{O��l��vF�N��5����y|L�C�d���AI<�(vq�g�>`%� �X!^b]9�+;���w:�鏲��!��nva�K����0eoNCk;�16�čA������2����Oq��夒�z��B4Q�ɬG���| K�iܝ0�꯾�Kܧ{ՏS��~��Ǡc�/��1��|-"�&G���P�|t���MX�NPP8v�ok7/�E�_H=\ka��O���:��W�l�Ď�R�+��ѿnKMvm$4O>���	�Y �Ւ��g
w9C���k�e�yYh��3S�	]n`j⠍�����m.�x���P��io���l�a�rmBZ�A��5ݣ�>vk��\���vs�ל��<T�q֒L������[�g��6Q�����p�,p�dv.C7�FL��^�Z��;��zw�z͇2�C�t���qo�3Q�)�~@��ޮ����<�̪��l�
7p���$~�z�8]���(v���D�+���)�c:�)���p(�==y�=W���Sn��ye�5�E�cNo蹟:t!f�+��u�g��r�7�<qTP��r���b=41^3�S���_(����.�=d�(�/�t��;���r�8��ԗ�nI�;��{�T�ٷ�kI��y�a�ȃ����8)�0�̻0�~4��ܞ�{ޡ��d��6�Ҹ%$+���ZƝ��z6�#:ƪ���D���Y��Ysv�:��v����t=�(���to�wA���y�
��A�t���}��PVԷ�M��U抖���>�y �ܫՃ�;����Y:�%���H�h5Y����,���;���M�t]:�
��܀G��`�"C�����g�k2����Cm�������aiwK�[��]ter<7x��	�]pM蜏@O��s�J�y�y����%�7=�0T֝ozN���N�\��ܬ���q����N�h22�(���u�{±LjFXf�FNc-���G�l��*>�J�G 㼳`c�[���"��ý��yNj��;��b���X��8z���Ñ޵j9��`!^��k5�&[�؆`4&r�Q-�
761!�m��x�L#����vLto�F+	f�������6��cT��O#U+�ʀ3:ӗ��ʅ�p[���:ږE��0�J)�m�!��_ .�u���	��M�fy�v�5;b�겺d1i��m�9�O��yɝ���.��uc�8�t�]�����Woq�8[-I-��|�s���#;�/�D����zaO����}K�#����Q�r��$,���)��&VWM�nX��\H�JwqM��d$��LP[�c�gy�ե��4J�P\�A�o�U�hkb�֚|F7�g���"��ݻ�r�g1�h�_v<�31�\��G�����u�4uΐ��9ewr��9 �vn�jX�v^P�#<�	E$��ܲ�Z��إ��-G��Qy�Z��{7�S�+�a,`B������	���nù��R�b�_X!ېew�Co'9V;&�{)�ߊ�8�b3+5-�qp���98�i���&*3>�2ɇp��X�G:mv�b��W;nt�۷�7����5I�Egd��1��YRu��|��UN�u��J�e|��%������V֑�×y�W5�Z�t��>�K�O�.x/���� �0�Etm@b+����R�ދq�1���HN�*I�W�௙���c���b��	H�D1��m�6�	�i+]��y�C�ܶ+��}���Cv�v�W]�I����iur!��Ŕ����ey0�q6{�;R�b�\;_Ko��Os=�0\�tPL�x� �K[H�p��=*wȱ��=YϤ��w9J�v1@�}��%��\ے(��:΄sufq9Xd�>}G,��\�c�g�=�a���,�v;T�w�e:]C\�M�c��U�2�wZӭ�!��c(��ˤ�1�x.�� K�	�A�ǭ����1���^�e�r�mp��_fؤ�oʵ��59J٣�XMh�?$0Pf��R�d���<v%t�=ثp.M7ͺ۠+�ɛ��7��F�C�&�R��ǹL}-�S#�Y����Z�i\*��8���O0�vڽ�04��� �"�=�N����0r��"��1̰������Ă��22���̪��C��I�f`ًYa6��9�Y��eXe���ff�5�fYY�EQFY6cce�FcfQ��Rd�Q���fNc�N��TeDfdF����ff8�c��$FXFdF4�fQfYc��՘�ưĳY�����3
�2�*++0̈��2,�j����kV��� ��2��&3,��d�,��21���r���s�Q��fe����f9`Vfe��feYfe�XLU6eFSf�V���̲�3(�r�0(� �h|@ @T�!;]
��KP��ႝIi.�=/]���˷�6IV�aT������Y�e����oe��]%\x���Y�-����&�����f���:�� X7�͞	};ưA�Y�n�=�0�7i�[W�ޭw��nnuc�Ą�~�@���|���٪����.pP]�c���Q�+s=���+��ɥ�<�nm��,SC��@�/��1�S����s���X=�zY�g��6��;��.M�I1�+�9[˦���h�#xd��X/�1���'�Z"����ތA~��w���N+:o�̎�y��|�d��b%f�O��=��.wg��P������S��Y�|��Qf�32��Z}�螬�����>P(՚�I����9s��_�ZL�W�/���-5��qX�;!�r�����q�
�<}�O�1�d�{�3�0)jyU��$��,�`c�I�D�VDb�NB`.[=^!a��&�=����6(m��T��/%��e�*���e�R${e	�zQ2�K�[��i2����M��uw� t:,98֛�hm�Dx�	j\��)�QV�K��8g��:�@qG���tp��/G�W6�R�p���P�vg��N��-�L�F�r�^J�я.ƕn�Y��1�î�A=��[��bs�3}��u��j�\�7�3�����@RÔ30E�˾q���P���p���Xd�zs;�������{�9t�޺_�h�������zPv�	��T��H`ݸ<(S��$��uz�����_�*<,�1��^S�=�uc�7`��Y��g&Q0�h��'����Q�����ϻ��*��Pqd�A�ަx��0k�R��?�_�ISzeæ`P�n:�e��'H�󾨧_���Ϙ�}Y���W�q�9����x���.�S=� [�ny�S�N���&����Y$��GY�/-�%DZ3ǭ������J�P�ɿ{[�G�$�U��w���H�o�җ���a��Z,�#s�E�]y�
YK�l{Õ=��\ڑ����7�E@���4K��z"q��zא|����Ȅ6��:�>�|����P�\��C��2"��~n�(���<G����t��z�b�^� ��e���Sob23�G'��҃����ɹ�nWb��nXذE�9M.�޹z����޾�%�|I��ُĿ{�I�\��cP���9��q`۰��)���B����Ax]��|1K�g�+�h��Y����G��C�������>ԮhB��h�4dZ�]�v��.S���7�L���}b*�c��U�]�:wh���N'Բ���wj���K�j��ݩ�lt';��R�tڝ��}T#��s:�X�dY��+�p�-+J�vM_
����$ߝ3�b/{;-]���쑻/s9����x�O�K�F|]
�KKFٙU�X�`��GG��Kǹ�;�o��y�����.��gDf��j
�j�~Թ6UC�:��T�����t�o��y)�+On�&?��i�r��Q�)�v�A@I�]�o���甧�=#Iw�Ht��Oo���/'�0�A��8T�W��^OZ<nY�i\`�ޓ��E�1.�v�����4 �˞[�u��)�I��}��X&��R�֟��04׸������nR�҉X��5�P_W�P� ��ڞ.k���p��RcҼ(�]K�����m֡F}�]�>����s�ZWN�����D[�E����P��vHN�����ήu���9Ʃ�D����夆�����wp����7�뇼�'���^Ύ#W���Y����M�]�XP�S�!��&��<��������q�c�|��J
�Ǽ"lnj�f�}�Q�|�ߩŬR�2W���6K�w�����K��50Ǫ�� �c�,��ʟK��:⋚-Z���ふ*lZ���SV�2qОuowJ�b���?�����W�od^ű��>�<}NTW�Z���:S#3z`�or6"��`8)�XK'ME�6kW��;G���9o�� 8����=���w�xk��0k�9,య�c2��О۵vs���i$�����OMw����T8֏e3y�̆h�]�l�"�������t����E�Ͻ!X�lu��+w�2���0��_�f,���K��E��ף\��ұ��{|��~m�#d�p����|�d��OR򿼼�şR�,�^����X+�&Ef�~�������n[/9�pGC��|���d뇼+֏��Eb�����g�_M�~����}&�"W�0����fX�s�>	�3U�vV��-6��b�����l��{��#pR��/8�(�tb�����6�ϓ��1�;&`����r9n�d�X���'K��\cX*�K��6�o��� �z�'<�*_�ˣ�#;�}�L���e��[Ǉ��u�c�ѯ��,Y\\Y�̼wf�P�C쾛ZqK5�x�|��%O�;j��d��0Y�.$��p���W�K�څY��@U�\}w�6մ��S*���L��V�,6��鷀� [��֐�򽙛*�i�J��c���;J��;�ʾ�imВWm��/Ah�j_P�k�۳!̣�E��p��P�����d���?�Ö�z���!���䡰��x(S2�ҙ�p�#�[V��n��'��Ѹ6�<prqa����<'�ȠGb��K��L�UU�kX�ό��5w?%6N�)�
�ݵ��ݩ8Tk��2+�pL�w��(D��մ���A�;Sۺ��������a�cӭ�ᲓY�آⶇ3U�3���cc���Β߽{��9��m��P����],\C,��U��uyґ.���w_c�Z�Ye{0Z���G���Ȗe\o���l�H��)��R���gڇZ���o�
����OwA�^ޓ���SX|�v\�9�ڮ8��=���Qyr&w��^4K�`��a�5����f'�~S=wu�㫇x&%E6�i�<�
{)������t��k��oy�[���i�\�,`ܶf|�Vt��q�8=(o�}x���;m���Y���az7�=�Xq�;��y"K��c���� �6)�L�S��O�q=Y����c�0�x@�UV�{���������I��L�*}DF�,�����QPR۞�B��B����V{޳���Y�m)g�Y�3[3kG�x�w���(8���ݐV�MY�Q��{Z2�d�r��ÁMx�<�������Q���nzf�h�E9��v�'~����}{'��W��UĚ�Ѓ�Q?���r���[���r�l��ȝ�i����=ʿ1�Q>�6(oRk��M���4�Mꄛ΢[+<��� ��2s�W����=�b�<軋���!�T�/%��_��U��v^
w"G>�ByNc���F�ٯy*��&n�.��{sVf�����Ij\��L\^.��d���crG�o���U�fG�E|G�5ؠ�׼���<��JԴ�I=��5�[�e����L�V��ے��с���͌��2�w:���0p���E�סּ�� <4+n��ӟ�a$���XB��f�3�S<f}�`��A�EB��J���eç4e��]Y�Y�b�o{��6��� �F��Q+��R�����E��t���Pfs&6��[û%�8������ߝ&"�RCi�4�
�[�tp��lM�(���.��}��N�p6�?G��o�Q�ܪ`�4�����z�e�B�yT���'�_O}v���~�y���q�{��Y+�/y��:s,��{gI-�z��w�k�������#Δ�[<ݪ�-�L�6)J�`�l�(r6�.y��Y3�JQ�w]�C��l�-�}�8�����v�e�O!�����Mm��;���ˊU�Rە��R>�Ͼ�����o�y~���%XLƉ�)�lt�}`<��� ������yY+ڕ�Ǽr�=EC(�=�B�c9m�Z�:f�����<DK�s��ŕ�_Ek]���^�un砜�:�Z1` ��+h�Mu�g!K�6(a���-�����v�:x��\ŭ����K���u>�Z�a{�����Rܕ:�5�@�݇S��}��Y����v^WSa?)���1�!�Ӕ`���i�xϗ,�9����FU��cΙ��Pi��-��j��6�`����.5}Ce���"�_ԽjeV�e0j�S��>=-]T�zo{�&���3ؖm|��>���i��ֵ�*�]-B�^4�6�"��9��]����c��om1qԼ�f{��&\��"�{}�ύF�e#ҩ>(D=ղ��>�~���ȸ�+���L�W<g>Յ��H��,�ʝ�q3�OZ<s��1���;{}����٢oR�g����-�:�fME�i��j'<�/}�xTOM%O�uc�^_�z���Ŝytw�3"u���/9��5ìuu��z^r� ����^{Z���;��m��oJ���}�\rgmס���������Q�"g��
�Y�	�6�3������ۗ�6�a �9-g3P��A�r���ݏ;[�V.��woW����z����v�����T6�@�J%�*��e�j�ظ�ڊT>i���$���	洛{��j{�qk���)���?x��0 ���s�ZWN�w�p���#B���D�f���;��9�s��|�+�+r��5v��(h�6�B.`��Hf�R��d�i��ɿk���y�Z��
w5�y^Ԍ2&z	V�.���gTC6;	��EO"�{\TE]/^t��Ɵ��R3ԗ�Ӟ���˅I��H��?����O�h�d�4G���܁�J�2wssw��N�(��ZY�������=/"��]�f�c���
��3�|��d�AP+��=O���g}�wa<`�;�>T�,N�p�qpu/$��m�=@�c���z����Yk��Jw���A�|4��<���{�+}n���9��化���M�s�zdD��:��:��kC����x�^��=��2���ڞJ�2�֍�J��pSttU�M�_���p��R8�g���������\�;�0S��t;�c���ܝp��z��`�n��i����m9��-;hP�w@��.�PΧ_�����c��fϛz�iY��U�f��a׃���Ӯ��z�X�SAy�m��{ҭ=�[k�w�����l�#���,G���J��(��B{�;̙E�d��� h,�1J�Ƭ9�{̗�.Qq������Hh#�A���-?��2������X�{+m��#B�c��ަ}�%��|��;А~I4UxQ�5�sTK��J&�P�	��JO����j�ѩb�l���/z��z�ff�N�F���Ϫ�K���ۭ��9��b�<�Z�f���=Y��F�.�<���;��E�f�ۻF�ޤ_ǋ�j�_��۷�&T"���y�--u��7��{�θ��o0?og�zz��X=i�C�@����e�
fXηJY�XW�w�ʓy�,mf��`��g���H��𞙜s�z�ٰGr�*$�x<G�?-���ԟi�}�:q��Q{)3�zR�/�n�~��;��"�G��p�OY"��H�=�y�R��S��ٖǱj���.�v/wT�������Q��dA�����xg�w�?Un5�kk�{x��r}�1��!���</��˃�Y���Ù�0RV�2*��`������
�ڭs.��7;�}�����O�<��+�>�1�
�σ�~�;+Uk>��0��d!��|�ԑ�5�a�˫��W.�f,z0��+��m����'U�ȩ�ݮw�"��:�a���d`��P��{Erc"��t�M妮��"g���7�N���TtR�]w8�SЯ���2P��W[Y��5de�(�KA�&5W9�XZT���O�������Խҏ+r���)�Cڅ�C<��WR&l�ntݿW�[�|�5�s��GP������I�zW��8�M�kE���G��ԋ��\��5_��x(�KYZ�.�^��n�d�X�/�ЉW�YfW�X�ױ�c���yY�B��+�:�H�}Y�+H�P��0n[3;����z;�o�X�s�;�����E�2��g���V^
���2O�
/E��G�I��T\�v�z=�뺛ƍ�V]�./�n�q�͊�Rj`��m`��3�&��s�-������Z����y.����A��p���cܰ�!�*��Iy(l-�^R�/ �vZu"G���JO�q���)��߅��D�Ӽ�zP���i�f��
��.�[ʮ,[�t��Pp�b��z�y�S�bvD=�G���<��,>��<��JԴ�IJ��uX���X�nl]C�=ӟ�Lm� �C���f�7sW�S�=�uc�Xn?xK�9d��pOY0��܏�/�w�R�oUf�uW+��Vv�+CUw|�B;���Fl��]Wn隋�;	.�]���enj��K��W*��֙b���{��w+�e�ʷ�ZV��P���.#VB��J�����M�F"-�<��p �sk8U�r� �)|/S;�	\7��6�/���5!I�s]'W:�s��]Ɨ�������ҧ׷|OKYf��g�dP+��F�&�m�e��}��	2Q�ޤQ����utG9��eL��w�< ����*wm�o ju<�W&�<��2)����bt��m�R�.�1�9�	]0�^g՜5�۪���]S')u�W#��.N�u�b�0K0���{*-u��Q�uӸ��wƷ;���v�nW)I:5�L�{�U�Uۙ�c�3(�H4��(�u�%J��%��׏��okUڊ�s������'E֮Ǔ7"t�`.U��Hr������
�u�"�,�V
b8��6�b�{��9�Cp^k��ޝͦ����'J�r��
Y+��m�<ޜO\�^ֆV�t����z���]�����y��)>�������b�4��W[�@kl�F������!PR���{�bv�[�=s�vjF�2�������6�h13�̍;vw8[�M�Y!��g2y44����n�1��EvSY���uZ����ݣTi�'	
)�2�����V�W2`�z�9ƇOI����W��9J��\˕�Ɨe���y� _dD�:Sxo�]GÃ���ȡV����(���9.����׽^�n��\�c5ZYG5�&��2������&S���s+ju(^�$��ܥ��i�kv�\�]9���){�����jgaŴ�WF�ݠ9����v���0< ؛ʻ�p�)S�8��V!;�Q��YDw>!R@�}��9�Z�K��C�Õ����u:M�6��vV��(�8:�g-o�d*] ���J�W$��}3���vm]<Uk��-p��G7��â�6Y j��{�t��`3�����i�͇s7�B��B��Sd����nR��j�Y_-Z�l�ʸ�*��f��ˁ�G���ΎV�x�-��T�_�D�(�|F_P�DEt��=����^��h�I��Y�2���l�I*.s�h9��*�
�t�Eg���e^�7:�h��k p"�Uu��ݾ�ͤ�Bn�S�j�c�]�j�vgV_�IS-l�pup�[R�$!�Z�g�gl�(�u��^�|�m1 �/=XS�]{kq��fNrjz՟�{�ЙN
{A�vǈ��׎\C���B�y���;u*��'*�
�i`i��`4�e�	�»��4ؗ(�P�YĬ����u������y�).����L�)�i锢�)j���6����}�;�r&��2��m�F���Ѫ%�B�ۍ����Nʷ�u�X�,ܐ>��J6��V�@��]w��gf��$��ժ��ˇL�)��1�(��L�h�e��*��"*�r�1Ī�	3,�+*�#"�33+�"����l+	���#Y�Y�e`YVa�YE%�E4e�f�Q�a��h�0`��p��
��b,��2(l�ʪj��#2����2����\��
ḭ5��:��0�"�q)����̣#0r�2$����h��3V�љEFe�9�fadٕ�E�Q�a��D�2"j�E�e�Ed��de�����f:�k"�d�3�,���rb,�0�p�#2d�ʇ$�S�EQFA��&h�l�Ȉ"�,���2�)�&�a��'(rs0�J2X�a�dZ��VXMUV�FVa�9QfdSFY%a�c�YAc������ŭk�@�~�R��/�$���T������3OqS�����ỽ�j<A�@��C�ŕ����N0X{D&\EAۜ�~�S~e�����>I�����se��D��f�B�j�b���S<gIcͩy��T/��1r�T/�C�ǁg���:��E��YH��I�u_jT���E��k��g�A�m̘!A�DO�kR�{����q���6�dv',��e��D���T�"�ꠁ�,���<�X����g�(�f��o���;IA��:�F�bJ^V˰�w�o�
b��P�gXeO6Eznc~�`��j������.��,��&cD���� /�U���ٳ]6�=ŒiǾ���W��w��-+������3��{�Ι`k�
>q�"Z�$��W��^��7�+&͜z�nf��?o֚�>��,ʦ]�\B�03����0���r�Y�����T��A:�6��V�� �����i�/%�<�wp5�@�۰��Nf���*�4�0�͍���d)�Y�57�{N��o>����XdI�+F;&��H��I�^]K~�tUn��N�/��4�
�^���A��x�y](�F�\��^�2�L���aaPL��^�?#=��]�5eW��=��,��!������n��+�SN�i��3�i{;�����tP�X�N��w���GV�E�����n��v����gl�t�bs�ڛI�wˎR�3l��l&K{8.mv��u��=E�0�v��3;� ��-�q��k}���b�����s�N�{L�f���P�WKP��A�#ir�_�Ȳ������s�9��n�Y�����P�v�&_��4���/>5���T��})n_��J��.�&ΖM`��WN�颱*�-��0���y�/�f�bWE�9L���ZOQ��]s�ϸ�mk�,Ͻf��t� �p ��:��}[2j�u�_A�+ޝ����=�w�������Xy����ف☡��<҉z���
�+ڬq���K�Z+	>�Ve��t��nGَ�9޳�W�J���S}<(;-�"�MB�E�=c�a�4��z��u��=ْ9J���w�攺��Wl�4tr���夆���U�5���]N��<�8��<����Vj�D�V|=����
��p.�L#'Ψ�o������ޚ�]�aA�i	�̞�L����\��܆���`��Z:Y;���A<7ժ�o��{�j� �}f��kc^�\�sҮ.�]�g��K�,/9l�Ӏ�{kjK���D��V�*$,������$P��h�P"�*m��@�sooi�3:��c7I���Cx�C\��OF�$e�Y�7��Y�!J��.J������S:h��B�+�<��p�ɖ_&���]��AWw����s.��+��&e��ڕ��
�P������̯v�-G�N��l�"Κ74*g�z�;�{s!�޻0ei6�U�F�'���6������^D�E�����o�]���"]T������\0fĐYNC�����9�b�P�v�]���(z9}�����}=K���TH��<F)��y�F���f���/E3�����-�fp�a���}�2u���G��U�c���:��R��崁hrC�����
e����r��.�ҳ^xm��e�2�����o�M��en6[�|b�����]*E�6�[�%~tb��L<\ڇu�����7�3�-��Vd�n�����y�����3���t{�|��4��t��Z��*�7�ۇ[+�/8VO/&y`��0Hl2.Y���ѭ�E��⸸�ʏ9͇GUl5�y..�!��wއm�����=���=l�0��h��RO%���yB�����U�\�ޱ.�ݵ��wӊU�η�8ԋOL�9�'�ȠG`����K��ZFa�4�|{<��I���8�tQ.��u���[ј��Ԟ�t_K5�N�ز�F���WaaP�i�y�H�J=&� (�ʜ�m����*ꜧs�t+����q���3���JC&n�{�7����b��2Jhg0���M�[8�җ'y�N흰4NK��]I��zK��IC�+��S��92���z�x�� �����֏{Y$@+԰��������[j�:���8j��3¡�f#�U��y�[9����3|i6��L�]TL�`�/��Y.x��u�-w���b]:���[�g��Z�(�uP�%�A�Hß]e��u����u2��Yc{|�fӢ��t}1����O{Ev8V5�tC�^�g���/3ʥϓ21�����={眴�m_#P�/�s	�:��a̷�x9[�;�b`�Z=K<�t5�(����L��;��iMѽ�H3�Zg�n:��<��}�-�V2u�C1w䦎b/g�r�c��y+��V]G^�yM�	Zk8�}�l��b��\OVz;�o�����f���~�糲�X�ч,�0t5g�
���UBM\*�P`�ٴyE��+�.]ױ���y�s�}��=�|����[�0�,�ʤ�>$���z� u5�	����,�|�{�\2۶*����s���r��aF�G�	��\�= z�.D@�W�%�u��X�bޣ�fYڶ�]͏0��N�����w7�{ǭr��;����pR�ʹ�X�_��C7^P�K'ϪN���f<��nZk�K����uG��s��n���8s�;�cܳ�|�X�U��7��j����e��>y0��R�W�^��h���L��]�~߼�Y_{*5�'�(��
�񠖥���M��ڭ�]<���K�<���\S�~QO\#�,Py��X|�x焠�KH�uH���fcw��4��� l=�J�]G�����j�u�C�p���<&K�d�f�Њ?�7��{<�����0{ @*� Ǵ�:+ب7���3 �0k�R��8P�Uj�<�����\�wk����yl���P��H��I�u_jTGP�E��k��r�~ջ��!hP:���[��u�2�ǎ��р9br���i P�|6�*��4*������<��۹�Dj�\�g���+��a�.�9�H�o�)y_�.��;֋7�L[��i�5�q�{��,>���Xb�__5�`���\�U��h�r�&�J'��	�;ּ�fxF��e��uK}�:Աr��O�nxөx�q���!������plyǈ��bz�t��|L�)�g�� P�f׋s�O0��[��hѹ�
tM�޲�1����.ejȕ����KG��ZF��I�Utҵ�랍�E��oj�nFN�T�Ws��E9|�_N�Vgmɛӂ�{z]ri�Q0գ�:����$[�{��S�r�Fr��U��:���s��Z�r����S�VX��n��2R^u�SrJ�u�l.���
�u�eKR���Tb��K�1�y�^��^(Ӿ~���^��;�'Q-��g�w�%C�@ty�|�Ë�2�(a�lצ�V܏͵�<�g���_Z��lU�Uf�L�=�x�/����-&6��|/1��J�Zrv�ww�[L��X�\������Yj/���� �X,b�'5Ɍ����M���F�]���Y�p��X�u�:f���P���<��g�x�>�Ho��b(�{�\����p�+:���/�����G�����ySE�s	�����՚�6��Z�`K���"9��vW<if�,��ل�Os�g���GN�j�U{v;������G��4OD� �qv��k��-:�OV�ɍg�;c������3g��Q�.��`�X�i�wH�J%uLƐ,��T2������z������ӝ��o|o���ρ�+9zz�!g&TłxPv��5�:E�b�B�.����=��1�ClG2׽�]�<�u�X5t�gz���HLe�yrP/ól��6�}ʘ~���8�;��@�A��-zY���<kGS���c��� �'rL\hu�5������Ǜ�(>����E�^��]ϥ�H�0����
Ώ�,�O�f����Zb�k>���WlZ�pL�E�����ZHV�\�1ٞ�{�J������jv;�M��;�^\w��W���>�
������P÷��"�y�%�y��k�9P.�d�z���t�-����,y���h�L�ޖ)s܍Y�"���z���e�	����������:��,!�֑y�k%S\/���/�8M�{j ~}��
�Hv��}�,�/f�o%f�(Xc����d��:���xe��Լ��ٶ�P'�O\������.���eת���f�����`On��{�5Mc�\h|V��r��Wx�H_m���չ�������xޣ=�4z��t�do�FPcӼz}��7?0���	u�������bO���i]!����՛r����,ܶfS��|#���wV��p��{E�Q�(b���s+z��c�9ޕ}X��B��A�h���Lm�bu9C�9c�&���P���ʣ�4��[�U�<ݟ+�t�5KiM�q�1C�.j%yъ,��	��s��n��}{�j�2�J7]�E�ڳस���Ӗs�FR��8rf�P�����]��j��@��jݱ����Y�GZ�f�K�c��<�[A\ʏ,�9�뾙Zñe�B
 y���v eu᭥jG�l�m�����%,m�w�~|�����>4=߮���V�a<E����$�zSHV���C��rv-ٕ��>�f��(����a� �l2%7�ݭV�E�+���ю��=[�ν��x�FN�:��|!�?��%�⬪������/���h��@mu2�Ù3�wfN�T��[7>;��K�iς�xw�ߏ�Xx�zfq�O[Ń〇N�>�HG��yN|�񈞤E��ǎVq�ηJ�顝%�~�Vg�x5S�92��x��Û^�Β��5�D�I](Uҍu��;UH��)5��`�⸃����$�y�g���5�_�^,Eǎ�yva��i,��t��uZ�h�sG�?9�Xw�����GT�>}�}^"��f@pGE�Q>;�˸s�h���)�����˼�9�	���1�~��g,o�ԫ=��C��$N�	%��X֥�Q�`n]Ã��^S�9�jt3�U^�f��b��Fs	k�f_�ߗͫ����k�J�P��oJ��[�)rʛ���A��Of,��Om4�^�}�u稗5�"�<nn�E��%�ffW2��\;囙�糶F�`i%��7�7�{E��y�o�(��c����Z��)��	�}Y\ؚ}3^����ީ�4B�
��f$(�f���\�.�)����r��JLήV�*Yz�7��Y㶤[�V`}��`N+:s�<G��n�}i��VEӓkSW��<������V{>��Y�,j�2�"�U0|9�ܶf
w1i'����;1չ���"y�V�V��^ �Bc�%��%ᄹ�T��Ү����)��T�����;�'+o��Y�'�O��]�df՛��iZii��UW��W¡&�mY��j�ݻS��Ӕ^��}�f���&�]���mW4�aTM��KSZ8��Y���?o�N��z�A]}��	�҉�=;�無�a�'�Y0��TF�	rL��1Փ�%����������K'ԩ���C�S�5x)�{�,��<��,>~�X���s/��%�8��{{tv'���@��X0$��C�WRg~��j3*8�x�����>����Y���vK�wɵ���Y0��OD�;�_ZY��>�{T�&fU�s�i)�3�of���n-s�(=�������ʳ�,�s�&���GR���س���Ma�����,���`��&����e,��N���T0Ө�}W�{��b2�*�5����ֺLM�N���`	��%會V<5�8�|�JZ5slI:�
����i�V�]�(�טv57q�ԥԹG�=E��Wv⻆^�9����j��L��z��};N��+r`��ǎ|�Z�5t�e��o�d�襉p�yte���ӳ�Aǽ��l�i�9�.������탁�$h7�����������O*:º�	1�Ϥ}�!�qz�j^iu�c��QS\�U���a�L���yV!��ڻ���\z��I&V1o�-C�h��nǷ�q�P����S���k�
;�j�G03�s���S���%�x�m+?Ek]��u�ּV�
)��\�rԙ�~�ޠ�%��{�w4'�����=Q����:��ڨ����ǀ��ES:��of@v�;����l�r��G�2i��=|�v��v=tlU���-tJǡ�.X��n;��6}Z���@��p��g��d�t��r�O-�8�Ɍ�Yj+ �5�7��.��Z��'9N�b4�§�\\�G>�"^�.m�9>�q|W�A2����ϫ}5֐ڋ6�y����x�`#�K��	�v�ㅖ��1P���&\��0����/ƣU������z�n� \(MݻLf�c��o#jŵ:]�[5:�;z�rBG�������уז�
��qUy�Α;f�WEJ|ힽ�R���=F�Ի�b�.�=g&ڮX32��w�۩Gg:�ڝMWu�8�o��F٢AɹO:�R�V�]�k�ǦJNVp����p`�2U�ܤ7��]��*f��p�2t����+o�̚���@7���&��EL�k7�h��NU�6�� v��xd�6%���;�桸.��)����9aR+2�u��X��F+ uʐ\'�6�l��pml;��qd&s�"J9��_as���4�G}�]���.Y�����B�A��N�z��u 1�{����@����@ӮL�h�Z��:����镽@媛�#2�˂�IS��\{8}f�Z��8�ql\r[�ޤ��Pء��������ٷ:�u��ɩ��8�+6c�[�Ņ�������|�83��ٓ�&p��ͺV���[�9AB��Gy[��M$���L� �����:3Y)[������[��t��v#��WG��c7��q�
�ɢ� u�ZuP�v�@�uL�A���h5������|��S&*JI%_�I��?p�+*ܴ��F��7ׂmU�����W���&�B��2��v��vq�c��ʢ=ݒke=ڬ*�-�>��B;�)Ӭ�gX҅k�vJ��2z
ѓ�գ4w\���k�'S5^��!G��r�';�t��]�[�%}u\�O]M�sWr�<J�����̾J�g%�m�z�(�;�y��8��-��ЬV�C�یA�;�.�s*h��B<��+8;�5}VU!&V�7�Ȱ
���o�=�W[k��k��&�Ժ뤧Ss���Z��0��oU#�A�.�n�aТv��9������E'[S+�b叼�[=�z��<��U>Z�A�jv���|9�K�["���͵��y�sX���	�z�7��ÑEu�y��K�[J�=99A����3%Θ�eL�܄H�B���:�p�1v��wb��J��s�>)�w�RȘ�O� �P}���yc�@*ҭ=�#��ME���}Y��T�nMdzXo����sm�"`�V^0�]m�f���;�ja��I}Vu�E��tI��t`ŒS����RQԺ���/A�
TT;�A��ϳfu�d����p��&T�pрshJ���+�i�J�ܿ�^�+Ѡj��PާA��[�ݷ܃�N3������5L�݄�^�v����9�\�G���hi��(:��'�v��)^��s�7�W_wv�8�H��F���o��`��
Q�P�t�2�@��
�m�S�q�O")���6*|�\�<x�r����!�1��v`R)YBhZ�W`�7O�wP��b]�K�u$]c)��v{���xh���+}{5D�P��uJ6k�Y ����övn�g��(3i��a�b�Գ	;�]�#W@�B�ē�L5�DdeA��3��f.���X�a��adU1���1�UR��Z25����f���4N�Ȝ""��hh�VEQTQ�Ȩ��s(���H��3*h�,I�,�0�$¡�3)),30��j�'"�Ȫ)�����%0�1�!+,�,�
,��j,�1��j�
,̪��#"�2�%�*�2L��0ĉ����J�()(�̌�r(����L�* ȳ��1"�� ¡�2
r ȧ' �2����b�h��	#10��3	
��r"�ʊJ2¢a�C'
'+0� #*1+,����(����1&�� ɣ	��*Ȇ��2i
�#��hrH�(b������1Ɉ�(��0�*��Ɍ̊b�0��̳'$l�%,2��*�����̬!���"��2h�*h�rrȪ)�2�$�""�����$2i2rL����(+*�i#2L� ���L������¨�*J��*)2r�*ʌ�
�p����0Q���0��=%ӧ�)J�oH}|���ǖ�X��O5.�s�S[F�J��v������s���70_IwF��]�t�׷s���l=t���h�Ơ6\C����r�v\��3ݳ	���klE�g;����߼��/�����.]#�QD�:Q+�$���ԃ��W�u枧R�j5K�w�<}����~h@����qB.�L�ر��.�>�Gē��qQ�I�\rT�lv�6������5=K_�q�j
��xzf��*b�<(;��hs�ZWN�wY�=��/L�w{ޙJ�{A�a���س�ڍ`���Wl�	k�ɕ��������}�K�֊�x��D_`!��g��u��g�k����F`S/Um�OQ�:s}8�>�mo���������`����?+��m໑<�ȸt���+{��9�	����EG]�ozne{��J|���Es��]�<�,x:��ߊ^+���"��{j��d B�L�O�{���[�[A��6x�N�N��p�8F�Ϧ��j�e3�۸aT�F'��}%�>�����r�g:�5�C���ƖzW��^:osw�Zǂ�����w��] s{l�R��zq��TW(J��]����ֳ�z�ߪjk�&��W�n�/t�
�b�18�3�#�)���mlƨd�[�����2���������,w��0b��s6�=hЂ<�G:F�2%0_@�ka��Q�f�;(�;)b�X����u�iw<-C��]����P�r�U��R{��`թ\K%�N�{*�ffMj�}��*j����V`8<���n[3)�ñ�~C=3��Q��\���_���m�MX��Hџn��H�!��9X���.��L��m�eӹ�|���ޮ���P�u�]�����SfT/��٘+-6��3VڙJ�`S:�5��F(�,�]I�~{Z.�3<���7�m��5t�^��}8��K�x�Ն��I��Ȓ\f�u�Sk&�X]Д�1�?L�s��ܜ��3��-\�옼a�q���f�����u"�<\Z(&f�L)m\���*��]zs:�̶&R"�8�y�xK��92���!�P�U lj�0�����^���>Y1��dPw�>����4�
e����K1�:zzfqɔ�p8q���X�*�&{�qa�`� �Ĭ}K���3��ιJ��M%��^�U��<D�~��/�˲Q��5��<߷�붟U�YIz�b���k2���w�j�(�p�خ�{����>��鞛��A]nG����B2�t޽�n7�����u�Xp����Q6�Ϩwq�7��(X:��`p�b�2�&Q���oLԶi-�˓.��F�vWn �̢d}�^3x����u�(�Y{��km���wU�ϛ��٪��9n�GDP�nFǄ��8V���ia�f;5���C��9����`����Twlr�\1�'M�2�����΢F�9}.2y�P'�'H
�v���C�3�*�󂂟Ia�a�Ƶ/t���.�� �AvP���Z�/g�ev,�Oy�=+�G�n^UiZ����)����w�}�v6�o�����v�8Skܤ!�Z�r9��ύ�6g#xd�k��~6x���u�ݗ���<G>���`.��S:Zy��(�;��7=T�D0L���I_*��aq�
T���Hؠۦg
w1i�D�~�V�9���{[3O�s��e���X���;И�Ic>�*�R��P������-E}���I��v�vy��e�̍� �vc>��B5��:�VP^qzRX���O�r��*�>}�P	Sn��f]�a4b�j|\����͍hSA��@ꤼ��uY}n�(�sq�t�w�^����yR�H��(O,�zQ2����s�P���]� �hqDi#*_�|�:^�Ջ����6۩�̽�/��ö�.�hCE�&�j���M��m�ܺ�L�J�h���n��em?NĹ�9��V^������{�j�����D����ᝂ<�Uʁ�P��7���|�VE���#�n�I�����գ]s��r�b����},�@ʿP�81����g9sW���G���y��Xx?G�9�(;Y�AfϚ����wm��G���"�d@i&��9��}i��O.
z�ײ�i'?{
W�|�oW�x��.ݞs:>}��Z�r�z�ɔL:�D�:D���!�U��{T�0kuGWpj���}7���7�hd��t������C�a�k�&��T��VG[Ϩ�/��^�o�B��g�X�{���A��>�����x�r���')�%���P�|4®��p�dWpX�K ��U�����i�87��V�0�]�q�$h6�����y�z�L����rWrG�{�R4 �fz�kךp��t�)�zU�k�J���a�L�`t˴{ա�-Bd�d�������hB���hq���f��
)�o	L�#�����]�Q��#B��y�Nv�����;1F�����QZ�~U��'3�x���V�ɮ�L�#�3�� ���==w��S#���>~w��gw�<oN��8}>Kp��\0�<�ӶOP>@�r�w���u��RW>��n�]��x���:�o{��~��˲2��3�Fe��@�3�[�_�R���g�kN��p�]p�[%����]�RΝ��0Ț��v 'f]�B����CP��2�q��x��74�wݽIWeY��1`�<��խ��ү=��;�����z���n��v= �.͖�|��C)֔��r���>�rZ�&_
|�z_I��L�����oT!��O<�n
�QX#���I����5�L~wn��m,����p>H瘩�K�Zs�@�~�/��kY2����o��d���};�6[��(3���
T5���ZZ<�C7�0�bzƘp���[�ηB�\��N>F-r�p��Wn���y�o丆I׮]��\�j����L;-'Y�3}�v���S����p�es�xHi��L�xؖh�iDA�	i}B`�ܞ<Ŏx˓g�V�0ob.{����wǠ�+|�B������j��.��҉$�kh&D΁w�?!�^CW/y��ң#+�_5�՞�[ཧU�-��^���Yɕ1L=�y�Z[������t���n�_-���.ٞ��3��>-��}S.���J�-B4L$�ʨż�w�-��=�k�Mz��d�>q�w�����z)W���S/Um��O��9z�#�|��=��Tp ��7(,'�������J���{��O|�P�����m!(e�+�cS����XS�;k��re�+�k�	�Og4n�Cg��#xv=��Nr���Ȥ}\($8y{����u���_6FӜ;6K޹)<�l�'�����I����S̺��S7y^�!�S��T�h��g��Ι�oL��j�i��(ٞ��ӣ�ꗟ4p7EMK'01�XC��!�V!�Y)���������Eu�Į�o����r�;�������9��:������8p�.���`U�z�>9]�s|_9
�������L��X����zW��/���^���c�\h|V�>�hu��Y����iO��R;/Hw�Z�w��/L�%����(g���\^��Ou�k���
��I��?m���	t��Ykx�M��P�Vpw��Eސo�v������^���Zɻ�;r�`�~��+֏���W�>�����V(0B�\>�
e����N�(^V{���U	,��!��S�}j��V���G��5�U��(q�����W�F(����kaF%�~��]{u��#7k��[�IƇ�]�ǅa�6��F�\dXUq��9�H��7}o�s|�b��ʸ�����k��<�&!5lN6%�n�j���b��⿾rj�`6�j=�v�+�W�m�Qϖ�xn4 4�F�{$k���Ϯ�J�S�
۵�+��m=������.�OW4�Z<��t	r�P�'&C�&b�M���mA��#�p��y�`���\�f4Z�i�KUs<n����ơ�]��3/�>y�o�,-=麜��6�S7;��Px�wNz�kL���r�yf.�jD�H�ʾ�K���z���{=�P1:�3�˱�n���p�9��}��Q�<}=38秭��蓎�����5����!k5��&�e
g��R��%�CIc_���eKZUS�ݳ������ZΞ��G�����v[??Y,�$��qWI�חa��r�(p&{Ʋ��Z&�����=�P�.��IY����=�"8�������c���������G�{�3Ow�����*W&c>r�\0Ih鹗pJ�Fϴ�LX��ﾣ��ڈ���s��F��t�����X�	W��/:�.�[A��p��'��Du�b/��I��D���{�u���x�S���x�m[E����z����$Xs-�]�U׸�V/�F2.���.Ls�^���7H��hB��1�x��ǫ�"qYӟyǈ��ʸ�ϓ���t���r�o�QC�췛~9�����l2/�SÐؠ��l��y��?x4e}�����X(�ۓ{ϰva"�X)j-���%���r�:n̆֝K䰌���}��㨦�r71E����6��m<�H���Y�8�^Q.�'3UwWi0�8���1��{8��D���S:�en�]z�Pk�?oKC�«e�U�#j	��wwb�V�y���릫}�Е�
ëИ��Xϧԗ�����J��WU�g��V�km5�u�'@�}Y�]9���oW�j~��]Y�o��Y��X����X�|n��_��*&_
�N4OB��NB)�o͍hSA��@ꤼ����f��k)�;�f̘�}�}G\\��3;�#�	�҉�=;�羔9�8'�Y0��y�S[Y�w��+5�l�u+|���)WI�gE9sW�S����&�y��X|��*�h�X�sl
���C�̉+9A�H�U FC��
9�_Zg���^S���x��>��<ˇc��&f������)��D��D��H�Dq}hPq^o+=L��w����]ۯ����1~;W�lj��g�J���=��;0�=i$��_3�s��	4�q�}�-��9mLo�W\�5�>��"�8�Z1��	�P��IP�Hu��d���F���f����a!K�U3@�^�����ޗI3/�]�{�
��#g�UЃ�m���b��{O[�Z�g��E��1٢�.=��j���w�oOr��ZOj�t��_�9�"��`�m��C��`E �W�$_(��e�5.XEbB�{���WLى�%N2:���qi>	ʠ�7]��>	כ(�����\��JȻ� oƂCk;=i����g�L�ǹL[Ҩ��0�Y��
�G��Z�n>�m9�m��S9��E�!3�o��C7G�"�������'��(�Jz�uί)�훮J9{����na3�s�Z���u�xdK��U��ZS&����#�xq]ʺ�3��t�Y箇b��M�������r��N�v�D��p�_�<�;�ܞ�|��ۯ�Vc�^h0nT!�۰�ϩ����T-+�ܭ���|����t�V+�gxV�Lԡ�4o������KU��&}pSh��t��r�O�P�y1�v7+-Dgd4���̛rWM7��V����څZ`��H瘩Ͻ.\�������j�{�6(��O�N��빧�Y����!a3C��ԝҡ����e��3�6a2�i��݉�)�M�������p�����ם���h�:T�q�H�j��v;+�4�j�����L�ìٺ��c���nsd��{lY�+{��L��e��ĳD�:Qq��8���uj�ޛޭ)5��ͫݑ\󩴌3]�|+�����!�q�}H�{����3��]Ǖ��
���U�#���,]BmK=X}������C����>b�R;��~o}�uuP���~,��$�2�nۋ2��Ih��������N��}�\�Zu:��2B<;Ŀ1]��z\7�^���ΰ�?��AV�>%&cNυ!�*��/��T�>^�A�_��O�.k�^_�ܬ��ꘅ��eByVWot�*��`��:��V�]�ۏ�p�>\�y��k��tG�N�v,-��T˅�+�v!)h=2�[s������K��c*fZHP�j%qq�˸z���A�k����F`S/!O� ����1N[�n���}��K�<|x�H�|B_�+����U"�o pK�O�X4�]xe��ql���>�t�fV`6#�,,����E����;i��c5[�i��9׵E/���2��c
�����y�m@�V�N[��:�Y>;���awՇ��}�OY�LC�yU�{vζ
�^�3�c/@�_b���q5�cpy�igޕ踟,fL~쵈�XO4[ͺ�8�-읩uz��е�Qh���D�ˏ�G�/L�%��y�e���|�%o+Yܻ�\�͊���t��Zާ�c�����]�G�]Ȭg
����Ķ阜�>�Ga� ���I�����t���4rlV�/��o���V�Ps\QG6�c����l��L�8ܣ�@/��.�sW�.���R�{e�3�|o�_VQTF���~�T��>L!��k�7SZ����ӳ	�E���tՙ�j�t-�v���Xm��h�!v�絛�5[Ym
���W��2h2���hX��E�DZ�~��C�k#��`b�H�z�␻͋�5�7n8F��L���cC=��is}O1�c����X*c��cF�qo�=��֚���̨���1ӢpV<t��m���|��� ytҰE��{o��̀����wi�\����v��}x�u�VRn�`�d���֎�]��븻h^}�f�ب�ܮ0:WW 䭵cW�k��U�׸/%��I�������1-�Q��l��9ef1�j�Bཨz�f�(pgj2�4��b��-��^��W4PÈ�c�*[}\�ښ���X���l����,E5c�XR�,/���7M2�$Ty��ZW��^g(E�C>_2@y�f&�*����y�(��d���5t��x W[�U&�-��Z���vZ�9��9N��;7o2,��g��s����3�Z}JgX�������xGz�S���º��Fɷ�7�3s8�6yAj�S�ɋ��wU̬�n�b�1>tuu�Bx2[c+�T:m-8�,*�)l+V�t$���U��ڳY��Y�o�֣!�KF\��P���R������.�&.�� �T����S,����'�a��{;��)Eh�؄�/)�oz��)-rbK�҅A'�0��.��O����7};�RCI��an'u�?�iQޙ��Z�X����}�,*�^j{P��(U���5ñ����鴵�?Z����*&y`S�E� �=u{��W��|�^,��{��	Rc2��[15�"����Vތݎ
�-�6��]���Zy2�S���m���[�m%|��3��rd�7S�o�mT��\�����xZ5*vu:.�)������ν؞Q�P��d��|�/r
b�Z��8�t��n��7E�_-
�~��dFj�fr�Gd�7�A���ya<ڦ�$�uy��<��X���yɝw$�o*�-l��u�HG��	|����GNV��8}v�Zyz1M�yکo�VD��3����ۤ{:���_�S�ub���J��ƍ�;c%�W�fJ����ږ�T���]�1jV�ѥ�k`5: gȵ���t�m��.ζ��7W�Vpl�2�"b�#����W$dۂ�ܥϩv<cN�:��e1o+�`R����U+.��w�C4!|��B�0�Fa�R�R��\m(�Y��+A�͘\�7�D*��.͜Ȼ���{+�:LZoj�pmC3b��r�9�u�
]�ziޕ��TI����j�GL���]���d2K��P ��$�)lrb�%�0�J����30��K1����+'&��3j�k%���2221�2L�3	�2*(�3�,��32���**��*�2"�Ȃ���31
&31j���b�(��#0��L�rL��j�`�0L�0*F�h"*�L��"f��'#3 �, ����*k'	����2"(p�3,��&%���33&s���J*�����"�[0��&�
B�� ����J
��,��Ȋ��*��2Ɍ̌��*i(�(r2���2H������!�J22�(���ʲ3033## �333�b)�2�̲2���1���"�2�32����(�2�(�"�2L��*l�
�#!��\2�*

�"��,��2�20��K3����)���h�3��2Ɋ,�32KD�0ʨ����$���*��,�31"("�	�#%��q���Ƞ�h��b$������31�����ć�}p�H\�Q�������R�J��rIw�}rJ�?u��{.
|�u�3�5W&N�&��\JD�/a����yӹ��3:��\3�["î��,�����V(0Eh���S-g�a�&������}k\�GB�=2��f�nގ-����Ic>����]YShN+[������z��l<�l:����C�N4=��<+q:�G�q�gª���`����g>�9���Dd��Vq���e��\��<�O���
������Du8F�E+�O*Uu9y7\��n�5�PL�λ3)�~C>O-ͭ2.7=�<resY�CԤD�V�5��`׺����ߐ3%�l'P�)�y��L��L���:�iϚ�A������@8�8}�r��4����P�C��F��H�]�)�ΩJ��M�,k��� �t�澴�w7\����Y��^��/+���� Q�GAt�x��v��^�~��#�*A	1S�0��N�:�[��=Ց���ppU�(C��˳|�i�جRge�y�1! 9�*��.�z�=����v��z`��ʄT�lQk�	-ѿ	�Z6}�
c�ۙ,�>���x7ˮ�M�x{	ë֘��T��a?h�{��Y�%:s�gj��������6wP�ջKO�4�LV-����`��i�1�p�+h�R�RrVm���.��ܙ��2d|���s�d�ێU���R>^�[ݧu$�e��'�!nϏ�^��W�)���9��z��X`ە�j^��V7.�z��vu��)��_Bor�8���pa!vP�	�}�e����Ύ�^4y�,���Hr���,�z�Mh:��IؽQ���^چ��Oe�u�ڗ�o
��{�5׆���Ο�'���e'{7�cE�</ѭ�®�wP�-�m��E�Pչa�W�탟r���Wr�)���<���>��o��=X=9�V]?;=��Bc�%��%ᄹ�ϵ�*�Z��=]@�+)��̶9g��q_��d>]-��C��,2=b��7�m+O*��X�M���ng��H^׳�a�/���+�7�D�V:1X�r9O�x͍k>��P:�\SF+��ٷ�7�$�J��S�H��͎�S�9��BygޔL�=;��k�R]F��̶�]���?msYA�Dq��JN�*��];L�*yr��G��`*�o4��z���6�ٽѽ�v�f�Ԡ�H��x�	<��
�/�2����z����^��'{sUǏ%��<a�޴�}o,���;W�����K)Z]��t�%;B��W�o��;�@(�o}OA���2���̅��ہ.��&{��m�o���U�x+� ����+��r��Vb��luI�X���h2^��u�w�˯q��J�X����59W]z�8�����}�y2��YD��H���
+��a���bT����ϴ�ݖ�ɶ�}�Ɵ/����EB��J���\6{��P��#� �g�t��A68U���p������>�i�Π�E�TɁ�+��Q��>r��¡��RK=�� ����u��Uä->V�RipC�_��e�;ҩ&ag���y�G��J^]������۵�<�r�����Ix����ۮ�qK����3��4�;��p�*��v)��.8���+���,�[\sk��hB��Ƈ��i5��ZVV�Z�Ӌ�7fu����'�����Q�_zC�L���[�^�o]%xd��_���R��x���S���	'�0���8+�AY�d�yo\����\�~�I`cƫ20Ng[ �QR��[���b��Zgٯ3��ܮ" m�qe9�6(ZLdwrяo�yx���x������Y��Ľ�2�XL�yp.��(�N#�w�s�fe9x'���B�+���ˣ{'���y�_��Թi��w�T�d+�B���9� ��N�Gr]���a�n]��4^S{\�b��X�*��K�+a��Wps+F�A\�޼�ϝ�Y��v��j0��-������]�g�}�6���|�B��NCG��A�C5U��b���S�b�K���bqu�"�3H^����o}OY��}�Lȣ:h`5�
�y��=�K��T3}�	��ebw{��ܧ�<�o���e�������k&R=r�'J��tW2Eo��l��8�V��`W<l%덺i�y��=�%����L��S�3��3�f��t�6
���]vL��DW���t�_�|��S�v�+�=[��!Os�b��B2���[��l;�4��{V��Ϡ�*�z'�Lk���)q-��2���p�^��ㅹY�ӌ�Ys���i��3��R�Er�������u�p���"�gZ;ڍ)u��;�(K\
�+�:*��J������B�" ���,������A�k��TcS-ë'G��]]e�,õv�'�j���ב3�T�p&aەDB�'�
�$_-�s���[�a�h=;;&#:C�d�4)O��b��৩t�}�Y�͎Gz��ݺgڰe3���T���Dג�����.* Am�W�<GP=���2�;l[��]�"R�/� ���.��0q���1,���}6cEw���oυ�1�7;X�o���񓕋�7}�X�ޏ����om���ɉ��/��Zi��eov���}M8f�'�V9G5FEz��m@>�¿9��:����6�E��VZ��A��|3��9,C�w����e�����{s8���P:W�
��1����x@��z��\��"�Vwj\�鹳��ۥ�Ƿ�p�Ŧ�>��",v^��]�����P�G1�4��<���}�,���L�C��x�X�����{8U���crٙNfN��ߛ>]�[�>�,W�>�t�G�}qV-�ޚ�����H0F
�.��L�\�H��^�=��aL�y����L�A��v6ݽ)FF�����K��+�.�!jQ!�3� ��@�Q��>Z���a��T8��N4=�3⬮'Rh��Eo�e��M�{��D{�=�p]Qt�A��yv�1X�}��0�Y8�dt�Co�v�|����x����u���|s-�B|W�˼we�a�	幵�ȸ��<��	�潋���'��m��/��Oow���#��h�W%���Z	�}N��L��6�sU���w�3�!���"��'���ZN=�Fmv,�M�H���W>z�#�y@	�z}�e�{o���������?fY{8
qw��ă��-��z����kwIA�9�A��W6&��z��7;�f�y��q�N�����4��C���st���N�*�݊f����k͜��s��A� �5��X��vB��ιJ��M%�s��~~�O=�-=�s�g'�S���E|�2�ܞ�Y���B�].*�']P|����D�����ז<��6s�W��j�z`�`9Y~�����
��!��f��¶H��5���&^��ORW�0�<�V��W�)(�EIv���+�d`~��N�l���W�Pس�x�3ϝo�>�H��fn�7���5���+బIa�ⶼ���ʸ���ރF-���|��w$���~����qa���T�I�	�~��+o\�/U`�咷��$=�������{=}�W������1M�?5�	�,��=�/~#Z�x���u�ò��kF+3�R�nl�����=�v���7W��=+ob3C��/��aG\)�%��eC�7T���/y��¯3�|k;|C���=��Z��XV�Lt�,g�/I��T.��������>�4�G�YL��s2ҟ����O��#��7��Y���>��PIL�����e�B��I���]����QK�,��;y~R�s��A:F%�d�s��W��aySs�����㞲������s&���rv^�ԧT�P.Y�*+膿/�)����}�������ِFB�L����cy<�8��� �Y�1$����_hP�|�����{K�j�|���9�����օ4FtQ�}�:^y�l(�K�g��g�
U���.��w"G6
�>��e���g<%k������f�o1�z�����C�#N%`�[�J�����g)˚��G�U�~Ź�x�)�y�%I�Y��u�~jvx羔�)uH��	<Ԕ(s����)��Wb�6�u-SӤ��;�sܨx�'?{����z���zɆ��D��h�/�
,�p^t:zgT�݁��mhx��.�����K� ��K[|'�8'�Cs#_��^�'�άU~�����|l����',���j�Pg�ʙ0?Ev<p(���	���K��=�X�7�������o��j�i,�WT����v�Ãz]%5�>�V{�wN�k�P<��~��7 �׮�l�ZJ�R��|�f��]�7O��f��_ݾ�!Y����}��>�*�M�X��o�BM��*�5�+�G�V�i3T��V���L��;�d��;���1=B�x�>>�3ۦw`Ld�QN�rDI-oJź"p�)9���o���:�RaBb��.�wP}|�fF9���©ήh0Eٓ�o
�SI�B�Y᪛����'p�n����b�W��F있���U)˥��9J�Ko�G����"�E=��8��.�H߽~�w��KK4�K��W��5"�`S3-�����������LL{���/�[K==l����\�~��<s#8�3OG�M�3��{t�Pt�N�`�ܮ"۰�ϩ����K#�wW{|{�/�z��Hfy����æa��Ip�bՀ��
�"9�|a'i3;�ua���^�8��nӹh��7��dcꝊ����]b�]/Zx*_���|)Ď}�R%����`�X
��y�u�;�m3�W�;L���Mlԝҡ�.�<p����_����[��#��ħ+��S<`Oo�{�ƣR�=��6�������ܻ�ͅٽWS�ۓ�Gp>���j�T������v�`μ�td`u� �� pp܁x�f�r��9Im�!��$GW�7:/|�y��yNB^��zׅG��YϺ����B������7A��Υ_��]*J}TϢ�(."���b\�6*\:ׄ����g)�h����x������2C��>|�T ߗ	�sq`3*�kt�U� }�'�����wt@��*��X_]J��f��������kT�3���
��S���c��o8��T�ꝶ\;pq�GU4��}��p�sB����D��X�i�I��Rhq�z�8����q̵Ӄ�t��:*�q/T�]�p��u�]��h�Y�mF��\/�]���hMy��ls{k�������X���I!��K��uP���r��q9�~�yb�F�8�֏��tK��U�N�>G0�ʢ!��З»��n�D��g�oa����M�zw0���=�������+,pSԦ���8J�!�u�z�Jk���~U<a�s-wg�Ԏ�����OgF���K>���-��,,��:a:l͸s�as����Xͺz�׺W1s�ٸp��+^��QL�_�[�Z��[O�[Mw����^�ܛ�������[}�U%������W����3m]i��zfIvF�����h��y�w�ݭ��܄0��x�pq��+AT]K��L�+��p�,Z\Kn��=f�T�nf��U��W\����{A�����'\=�^�|l��,����WA�+D��4�x�w�-���7O�z�.�����<pM���_����G��5ʭ�C��*�-���xÁ�
@�\ٕ����iN��tۦo:jҬ��U�t�/���⹹̐���7[[|���N��|hm��Z@�t*kl�켔��>�in�"+�{�f����nS��d)1@��TB9�����,�d��L��u�پ�½6�]E���r��d)~���x��ÝP�+y'왌��Xk���х�au���n./�(6��<����Lթ�Ui�.��b��(3qO.�e�	��1y�bq�ȔPܣv�f�Wx	�����X��j�'H���5��f^;��S���wNz�ȸ����=���^��=�C:S�Ѽb���wsq>9�D��:bL���P�e����v�Ӈ��.�o�%�x���n���y#��w�3�zz�,�Z�D��\��E��Ր�}!,V�F��KW�O�;X��ឝY�=�U1q��E|�	����ȢH�t���]uA��<��nБW�K���k/��M��5�I���Y~����pU�(C��˳ �h^U��#|zV�Y���������Ar����X_�޵`ޘ)+r�%�C�Z�KGM̻�׮���û�g���]y�ٿU�*���~���]��kiB���W�
����cZ�w����o�Zț��)Iu��N��\G	����wt�����<3o\�/U`�������)�l��ǳ��gV�{X� �c�g;zV�fB����L�8�*������䆐�����;u"���k��tʦ.��JڥRJĕ��3r.�CS�X�!�a�w���,��p�︖2�\;j�66�G�*Bu�0�U���9�lQq����grg�}�k�6F�d�:�8��ŝA޻���qj �`�4��6�6�ז@w��ԶR�Tv�^dg�f�i���S%�����;�/-R�fW3du7�ڎr����ې��J�УgR��Uׇw���(W1�|Q��Ag����):����^f\l�~�	���E��4'C��e�_�,�N�r�*�nn����z�1dz���K���]ĺ��݇�
�tWk�Q<Z�֐(��r��u̙�����Ju�	�S
-��*P0LY*5ͱ;�1�u��Kw"���#��I{:5Q$D.p��bM�X��o[��չ�sN�@i\8IP��j����yW�6��][�0�b^�Yֳ[7;�R�";�����E���M+78SQP�K�����C��b�5��$W�U���62�M1��P)s�V8�1�)��T�i=�j��>�Ti��t H�����ۇ��q{V�c�7�≠;�-��0�]��4g@�V;��}nڢw\=��:]8,���aSʗnѮ\g�M;]}�fm$�m��1�6��\�ܟN�:�i�^ڎc�nhR�G["�Tj�J!��p�<u%�%ǲ�4E��ۘ�u��u��n�ą��e.�ri�wf�#�nT"�-�"���
Q�f;x�ǎ=��/7BJS��^U���L]#X*���ٻ����U��Y͜E�����}���_�`yZ�l�Y�Me�Yq'33+t��q@��wQ��>ӝ�ﻤ߻`�w�t���vEn�M��b5��]䮏'U�ő�s���n�u��Qm��6�|�*N�SZ�n�+Y���֑��3�������b륬1\�n��[����Ss*f�6`�\2�v�
��W]���Ր6�Ό,���F�9�g�n��Oo9�n�yk�`�li�����jם-
7�����̪d�¾&X��*�ߝsŀ`)�ݗF�F��%!eX���lR� N;�a����'�<��ޮ��c�/��8�w�oJZ��3^�!���u}�9��x����d��{{�db�/����L�Rz�x����9-�S�>;�����5n�(.v̠n���g�0"��|*WK]��� \�~,�wZ���Ncm�4�vh�D4ڒ�{�9f
�P�'3;,���F�MH�l�0���
���:�7y�ӫ"w��J�K��]���V��
���gK�G|�DbV�����Xj�u�f��-͑�My
�R���WSx*�$��k��.֊d��D}���gx�H��W�x�ϵ�"�0�q����ԕ"���zV:C��ۻ{�z}���ֵ,E&fU�9.A�TUTaAf)T�e5,EDQ6FUPQ��TVFESAAXa�@Y�LIEQHEA5L�I�fT��D�`�KATUQ$�ET�9d��e�9�NTAP�YQ4D��QE�œTSAE!��14RU0T���D�5HX�d�LS1FK�LY�ECT�A���E%MDTUP�HMAAU9�%dٕM�مf!�TQ1U2�MDC��$�U�Q1�ITR՘��0QLA$DA%Fc���44�STETQA$S�N�Q��a�9���Y@FfԵL�UTf.TLU��PPREA0PS6`e@E�fSFFD�SBQEE$Va�a�3U%!��d�@URD�U35��UfCTUE�dL��%!C��C�a���T�E%4519��!�Y9fQQI4�QU5�QAT�S��PIT�NK�D�`SEVf3E	G���E ��Uvxu%U�l���z�AP�zd����2����q�L��Cb�5u�B���.7���&j��g��.�:��p���ꦎ��_{��j��^-hBx*��#�8���<vԋ�o����à��mקI��W8�Ppm�*{�����
���J�؆	Y�1�ߋ��Xb��Ɲ��o�z�#���lUh3�����l��Z��\OVGp��Xp�5�`{�Yim)������+��7�w{���B��:�Q&C���3!�]-��}�nS��9y,H��X�ed�q{R*z�w
3�h~3䗇/ ��f�;��|�W�&-���֪�W��s|n�wr�ǝ �P:��)�+��Eqz.]��H��
��.zw�Ï����џey¤��a]ZĿ}%��x�Tі4��rLKb�J��N�;N\��=p����Y�壗��g�����L�W~�k���D:��H�@��`�\��9��/�3�F��`뛳��s�O�@�����i'?{�S0'���=d�L4Mt�4G���z���wӝҮ��)A����S=�),y�W�tP�Y%L]~{!ÂxT6&Gk+Wʳ��K�q�V��}�g��r�tfm�j�v�JɌ�Ȏ�T7�����1�ߚ��p_E��(P��A���C�:��?�vP��R�<s��睱rB���>X�2J����d�|,�ܼ�1�Dǜ3Cm��uqc���;�����R � �����|\��Y�3�?�d��>��x�r���'#]�ͷ���Ufo�z�Nk�3��IW��3�E�RL�RȤ�;MaޕIpCȮ�+m�crQ�*vc�����Rx��3�y[˱�;֒f�৕ԭ��u�S�]���>�f��eH����;�݋'o�V�P,=1��;�J%o���-WX���m&ii�)�zHK�N}��l�����\U�
7�#��ORΖH��~�a����ڳ*��W�^u*�¤�-wZ��]�0nWb��nX؄�x��1��g�j<m\���<&N0�>y~=�Z� ]>���,�����L�>̀�r��0m�qe9�7ҡidu��=�=8�f].h��r��Y՜),�=�V6�Հ��_
�����Nm�3>�/�.[���ъ�Z�}ݽ4q�(B<W���: ��Mz��L/����N$py��,����R�$�o>�m^M���#5�g�*��\��4�:��J�̻��&Z^�f;�i���\��v:�Z����i��u�Ü��l쉳�e,�#��qv���+x��5` ��:,5��m��J��u{`�\/7��.4���#l��J����<��K*n�Ba�M=l����Wܻ�OC��O�oޔmG;  N��17'g���������h�	{]���Q��e#���G����җ]�u8N֦V��g\�6���=,����z�(5afn�&=���[ޯ|��Dh�0�U���Ǖ,y�ߎ�G��'?^��q�q���sǫ�:�OV��;�]��B2��;�L�h��^�B���'qz`�o7�bR���A2*���Ys�ةp�^��Cr�W=S�O'�+�^�ݷ��N���?
�-C�"�MB�n���XE�u��amF�����j��QD�b�m�~m�W��ðm�ϦT"XBx<���}y %�^�)�
돰qĳ���;�s-�wtp�v��%����v��DCo	�8.��>[y�
��ؗ��^�I��c�c	u�sưk܍YȬ�m�ORΖN�
�o����,w�c����a���,)u�<�3g����t�ޖ9,�\��`�e�.�O��nm��W�����ջ7�<��uҽ#l��d����e2}~uQl*�ipP�sY�^����U�׬j>��;��b��XeY��O�����TYz��o��w��ˣ�w��s{Ak����@ž�#�tn]ҳKVf�<y�aغU���j׿X��-ڑX��CJu�c��B.�w��|j��iu�D~m�%���w��"=xw�>ݗ���g6�;�3r�T�k�Mc�\G��t�X������'�q������z	.��m/;��W2�#�m�__���1򸽫���Zu*����]�G�ԋ�8U����lT6{�(��\��5�-{m}���(��o�c>���Z����Ŕ��-^!��z<�����#�8�+=�+��+�[A��S��',x�޿��/�e��֚�%��S��9ޛ���-o�Ɔ�!�6�^h�za0�:����hxN4=���g��Ѷ¿x���/mξ���'B���Zʪ���TG.���S�}��W��옼<�gӍ�~;���:G�z��wT��$X��.,������<C@�环����d�Rr�d����ǯ/˱C�ڸ���h��@mu2�L�M(��#N'��O]���Uڝis��5ݹ�遲�m�>�2���8t�B�j%b�5�B���)@ifcv�9�}w��������{��>������b��"�G>.��%�A�(�#����m�����f�v�<�.O�mge�^n�k�dd�g�ۦ/9޹���	 V��P�����B��q�,<=�2���Z�s��K���lM|�bUbeo:���p�gn�7��mu7��yM̽�Mh�V�뫓}mj�o�#4�.�!�|��w0SԷG|���q�`��>������+"�]�^pU����˳�qd�Q�^����t�`6�p��P�ޫ/F���7�
JÕ�.�.#�Dt���{�1HI1L�ǹ�uc�Y��o�@T
�pb=��u.�X��Uk>�.��pXV$��k�{����)U{�O>d�A�sǾgw��<�]�+j�*�)1�9o�xem�E�B'Qz�zu�S���oi��+�"�ޑ<��^?5�	�&	�=�/H�W�mH�e�.)�^+$���{_���w�w�۲��E�����nE[���-/E{Rơ���i��?(����O�Eރ���f`�s�՞��R��V�VZ���ĎCz�c�۸��z�Jઅ�y�Bﳨ�
d8�S���.��xơ����{prP�j�~�y��d�΃��0l�i�«M�ʪ��\�o���gQ-��]�&-�������y�*�n�?z�Y�����X�*@�w��LtEh�����D������D�I��沌�:Q��������\����c4񚝎�t�v����Rڇ(�'���.��Z���-��"���8[��G�S]�����n�O���i���M��JW�T
�]\��:wcA��'R�`������[{
�q����WSt�d��m?&s솔{QYHmM�J�p%�0l%�L��Ϯ��S�<����
[��q�ӧ�r�ݲ�)�~��k���y���be#��@�<C�jxP��\�A��`��IgL��<��{)3>�/����cH��f��<���	=l0@�$���_������?WV�YW>B���NV�=��0k�y��T/V	*b���C�`P�옺��mm��s_;��F��%>�du+��v�lY��k��gPg��S&Põ����Ǎ���t��E.�˄����n��Uo":��yh��.�ߏ���Xsz]%5,�Ř����35F�{3�"��I�t��ݖ�����x:���/�^Z/��k�}Ct�Ռ�{;�����΢���&�q�n
d����j�쥈>�[�0\����ȆQ}�P����OU�.ki��-ü%��po�8�3԰t�Ez�b�^��j��z�?_CR��F�nz���ל��0C�+�A��E��)�����v�:x�-0��2s�Τ�lP����$��$-o �m��QT�Kva�ї=�;m��)V6���Ȭ��U�=1m �rf���Y�B�yQED�
�Yz�H@K"q���*R(2�3���,�ܳW��/�S\�Dqc�K�o��9]Jo$�ɹGu��ُ��Hޤ��O�ф���ӶOP���Ez���8�
s0lP��Gp�*�z�,�op����*Hs'�5�k�]+�A�s�Y�JҬc�j�T���w�pm�19W^�d���M��r>����q0�	�y�=e���SH��R��L��H��b�K�K�V�Y��w5�3=�w�"�v�����k&T=���Zh3ԝ�T6U@x����)^��������<�����k�e��a/k�wύF�L�z��h���!�ۭ���ol�v�o=�Iw�Ht���;Y�3vY0��x,����8S<��h�f����'�"��?^_�5]��zQ0X+N���w]1��u枮3Ps��ؽ=P���j�g��3 3W7'��kӃ�϶��(��PưPL���2˞��\:ץ���nVr�e��X�)�n7�����,���X'��<�-.�uP���"�:�ذ�j�\�W��9.�_��Ӂ&sP�L2���Cϣ$��8-%�Z<���k��zk�CEh&��Z��~OE����t>�뫮ۭ�y�HS <�Q �s�L�2� 䛗��������s�Bx�T�H�uѱ:)�Ϋ�rg07Do�g9�n�]��*;ʻo-�/�M���-͢�v����Z���h��u�����W���P{e�fZ�«�,8)�8��bDC���WyX��m�Vأ��wL���Q̀h�|R�x:��FoK����+,pSԺQ>4Q�Y�7�|}τ;�Y���h����9��)q^vq~s�Pެ���cXY������G��=�޶��v^)��S�����L9qp���y���(E�v�,ny�iu	���wTk����t+����^�������k�e�<-6��e���+����u���������XF�6�(`�s+�ں{��gڵ+�>��]���w"�2�o��iݯv�Zr`Rs�u�;h���;��=C���L���h���~1f��Zv�yz3��s�5�[�%p��py���f'SS0'.�{5A�Nގ-����w������י��M��4Ԙ�R�*<'%�Qw��:����C�q��Ϧc�i��ɝ�o��~��ҿ|&/j��UW��뮶�ϋ9ձ�ϲb�π�My㑤2�c>���˷[�ju�wK���Ky��[������xR�;T5{�&{i��]��
eg>ɢC��]g�'��U��hqo&t}��(c����!� �=Y�@��)�T��R��������Rnv�������Eq�{���w����'Y���kU�H�eqq`���������1<�6�"��͍��b��g�\v��>9�\�b�j�$IT���@t.�^P�e�4��F��{��w��uÖ�������yg �6�k���M̮���@��Q+���K����6Z��v��Iy�#���.�%6���U1q�E|�L�ve΃d���\W�ؕ�#�n���v�3	���8:�cT�FӇ`��ޯ8*��!ۙva���#{�?(�<����]��DYj
\g]e�C~Y�������I[���1���-p̐%�P}\|eN�ߏ���H� �]蕶��i����o���y,vV��|sz]%z�s�����fnK�g�q+{�jP�_'��CK���N�l�j�ӣʥ���Yᛩ�UD�y�M�x�+}=�9*Y����6�'n�a�LJ�mq��K 6�e;ڼ��|5��<��:z��ֆ�5�7ԡ�~#�6ݟ�{�����l/v;��(rݖ�1��J�e=��D�ݦn %�un��L����7��j�DR:W�*Ñފ��ĦS�Yu�d��DbN�\�i�d��`c�Ba�{���ܣ�%�1��ͬ�]���#�Pm�Q��r�uȍ�&H���L��ƞG�;�W 9 ���1J��Z�ӳQe)�|�y��w{���X�(}p]�8�ܶfS��O�.'�=�6�aâxׅe:��+Y#�~�ڷ��c`~KY�
�:�0������-E�
d8��s2|�[���_���=uΫ�;��b��*ͳc�+]��M��UWR��	7�D�V:1_�)�A��11~��y�5��E����Ц�ڠuR^K�Y]V^}J���v^S�86
˥z��n{���S�w.rW���{�^��C��8��,��Qi.I�`%�L�]|w;GZ����.�}�:���Y_�tO<��,>��<�ȃ�-#���"��'����z��Fq�s��t�ތ��v��Q��৮{*Ƒrs���	~~�/�[�'���� V�����\��z�z�"@�\/��J�K��ץZ�ڧ�L���� �"�z��*b���C�}����{����W�mkYH�5҉X�du+!���q~�]���g�b�L���s�X�ˡ~�y�zI���:>LN���Cs)%C�"��\Eo�L�;k�O���ޗI�>/27^��U��c/.Z`إH��O�Ӂ�N�gmu֦RZ��]���N<�k)�̆�,9�<���%�(��,�[���N;&��j�9�|���eAKwv\�.��� &���o`LoϗwD6���k��W��}�:��X�%��+��&�뿅�8�i��]	Bb�)R�x!��Qn�^7��3�w��,�����g3�����/F��}�a���DQ�6���; �X��b)EƏ�y(j�˾���7Z%Rm.!��β���|�ޖW/���!K�rb���B���H��q����8��/�Tg�j'2ph�Ҍst*�q��+ݣSGM��&�N��!*Jk�fŤ�U�d�+zYf��M)�jZgn�Y4��h��k��M*	M��o}wsWV�p�U#vp���+���:�.2���8�n��-�]�b�gQu�Wu��:V�*Jn]Zdr���0�z\Ձ0�5��=�gZ(�ȏ6Q��L-+#w.P�j�{;*c�\Ҧ������v�}*�A[l�T�-�=�hɴ����&[�i�z��+z�}���V�ҞiQw,▯VP�.��U�Ј��N^y�ot�ˈ�>�[����Ã���W1=j��WQ̳,�1qu���w�+eY�eԽ+e��J]�w@��@�����ynr[�:N��ӊ��K�BS�B�[pJD;�{�sm�d��#�A��q���=�+�+ hJ�wD�����%a�쮗`��9Lab��x��f�Xf��a>�V\tYv��6t`7TkoPP=FvGY�q怑f~$�g&��[^�o��Px�EQ�94=wc�/B���n!�C���n#��tΧ Ԕ׏0 T��)����a��d����κ�-� *���ڊ����׽���F���n9e���e���2�� ������11=���8#%d���7j�swp��vb��]�pћ/n�1�>g��	���p��xq.;���v���q�����&�«SǓ+W8+%��=��A�r����ƒh��N�t�(�u7jV���� ���ܭ|�Jz��cwV����m��sf� H�l��:�Ya�9��Zhރj�2�Ԋmmvs[���=�ɐ��'J���W�Fٵ(K����a�[r��p0�tR�F���޾����$��I3
���]�f�6�s[������nN[���"z�>�,��N�%wS��⹓�m�`�']X;'!�_^�ǂ��:T[��6/tmbo���@� _D���Eִ�ܬL^�����4�l��D�v����7���ѫ�{���e�y�o�Q�ۋn
"d���v6h�e�k���<��WX�Л�h ��[��x����+w�R���뤫{����*k��<���|gY�����������P���:<��s�}�߼��;��S�=*���(��*�+3"�������&�
2�%���"���
L�)��� �����������&���B�2�a� H��r�����̘��������(,̚���l�r)(�f"*�����)J&'#%�,+0r��L�h�2̘�k3,%�&��,�R�#*��������*��,�`&����0������b(
��)��R"��� �Ģ������ �����
$�ɉ,�
Z���������"��J�*����(�`�3(��������3(h����j�(��������
I�J*H��h�����#��*���������(�h)b�����������b��(���*�����������*���0()����3)(f�����)f�2��(�*����ih�)()h(���B"��������
N��믵����:�\���FM�]�'Y��/8� \u���v�]rC6"�]Z�l��YW�{�G�i1����������J�L���o�Q����8#�F��8��˰�'���=���y7\.���/�C�&׹�zH^7˼���VL&�&cD�$�J'�U���^A��+|�\��C�
S[���=���sWRY��}5��^�r��qqV5�q�8f'�Oe�5�k�j+Z�0�v�W)��#o|��ռ�pVb��:)�]k�k�1�C�w�@t��r�X==l�h��(��߫F�//lk|���~Ss&��TΥc%C`c����qg�vYNf�H|g�u�d,������;�=F=�t�Cs�1_�9��o���GG��t̞�}�x3��rۓn��6�`������g��WJ/�SV)z��*_���|)č���r��~��Y��d9��g��m2"s�O�=�tFkZ�2���� t��ܓ�T6B�b.�b��y�t}ݴ����~b���ɎzƘp'�ܟ912���]����P%�����L�:{6�K"�#���b`�x��XY��a0����1+�fڿ��p���#E�<���:���d��y,���j�Rغ�:�bhe���Jz�]��%WH_�>\�z4��h���+Yx����CU��_c��|C�
��W�C	�G�9�w�1[��X�8��ν�Mu����gyq?]�Yx_k|�c��48�6���E�N��u�͚&gR�6V�l �au �
�W�N��ռ�!=�����H��Y$��'�7����}c9@;ơt�9ҔJꙍg�"���a�eͧ���y~;�Z}@��'����8������Em�G�?*�����
��K�r��>o�]�9��^�����L������x�n\=���J�-B4L%�����%t댺�x%�՛�t铙�q��b��S�>��=�TcS/"�h���O����l	TD��b�R��g��Z���Ԍ�w9'�9bS0�۾���^P�S���sưh{��9��৩gK'l+4YK�/b{�&P�<����^�S��^��-0i�җ��N�"��ڀ>�e��uY�^�'%��z��]����`#�c�
��T�Ex^W�����[�Z���u��[M\��
�v9�b~국��Sx� ��z��Yv��󴮗+��K��Gaۥ��9�&�w�u�@���Te=�����{��`�+�."�&G�[��]N�)��N��e�,6��-e,;W���A��٩{`̢+���2�v0�w4�镴 �"��VJg�<��M�x�X��1���<�A˅w)�:�{�c<u�lդ�	ڤ�Ρ̵1���U��m'
X��/5g��x��e_vsؙi�!V�����x�18���J�[n�ԇ�p�޿����a���>��'\=����oM\H�!��l�c�d�s���.�{� ���������P��l3/�w9C����7�-ϵl�5�Eˡ;Q�v��y�����Tn
��0R��b�Z�V��Ͻ0�l��'/��h{�ۭk���~��/u����0Vf��҈��ŵU�e�˩��r)�b1?��d�H�sûIe�=�#�l+�X������b����k�,�.$3@�vZt!�3����i�oF�"E�����G_�8Q�}=|ױx]�I��_j�6S-�єҊ>}�ٵ����܏�s{l�'n����8�k�d��o�z�, �!�t!f�W�.k�s�e��G�z':e*�O�o�3�zK���ƿ}+3Ǽ����V��L�w>��Y��`����#!�ܞ�����W	�\a�w+�x}��Y�&
6��8j��|�<"��1��L:y����o��}�1��C½G�<�x�?��X_��E�7�
I��L�	���̾ԗ��e"���#�V���G����h�ΰj����.'��
��ث_��@�V�~�٩��kG��*��.���C7�pn-������gK�=��j�.���-�{i{+&�$�s����Ԕ+K����i�R���E�2��ξˊ��=^�d`uѿ	U֍�J�@�#�?R�%�ϵ�oK����=������nv����t<�bb:Ƶ/}ҏ+ܻ��X���}�Zt3�*�5���&dv=C��yNo8{����>�]�J�;��n�aT�8�M��!<�5綥�Pr�d�P�z�}a�w06?54��U����xm�5K��Y���U��p�P�-����lN��޷��Sg��YJ��,5yc���w�x�P`��N����*��²꟝��.��}��Bz��z��,�gc�VhLtK��\0��5>7�E��
d8��s2 �[�,c�a�&OsNo��0�rx�z�mf���h��I`|bKG�S�=���p3��'_^���G�;Ϛ��O�df�8���:J�M���1���?69:�"��B���f�Mv�c��Ou�=;��k	ƻ�}0��ӉrLKb�J��|,��Wt1��g1���
��w��C�}t���UqZ�6�y�zPv�L�u� F!���@`��X�}���M�8�}��SA�(mu?�q��\ݥ�o���@+o*5)�������z��\a�l@�+rn+#���R����57�[� Ob�0�5x��ص]u;�1�|s�-�q֌,<3��k�魐�80���5':rɍ�������Ln��|�̨|ؕcH�9��}=.yd�f���&��\���=����&�"L38�$^��a�3�Q�R`��*��?�^���d�{6Q"~=$����Y}~��ײB�G�t�
�]
��3Gg#����D����L=��I��Ugs^`�mh���>�����ґ~YR����F��S@��XE�U��V5̓e�����Pyi��Ev�q<�(�ۙ\�- u��7=��_n�[�o��]M=/Ӫ�1���� ���]=��f4N��I��<�;ּ�ϸSCû�B�y���'����Q���!����P����p|�x��Y�����z#0�ْjg���ص�֚��ي~��\~Z|+j�d�Z�k�1�cb�M��-��zz��Y�ݏ��H���������!��R���ՙU�y*�2��� ��aŔ�M?Z64-ū�zud��,�����cѢ
��͖��g,�`/��/x�|�x F�'Z��%/�4���dLB� ;h��u�P��ʰƺ},tV�R52{���̽L7[Ou�5ů�Aa1�����`
�{�Fy:�{������/m���igr i�y%�v����i8d�x��[o��*q��;����[�q��-�8,L����m��|c\]�}�i�W��axWxs/�dQ�B�R�Ѷ})y�.���x�޾Q�����s�����W4�*\��=�v3ZԵw²�!-4
�z�������&�c��w�,mfAv�f���J��C7e��4ß'���j�cf�j-]�����z�9ӎc7@��q$v�ꡳ��,Յ��0�lOs�g&V���8i���Xwj����'3}�N�g_�g(�`�J#eqf�qvR����'^i��S�����Y�q���E푪_v��X����v`x�x�6��҉$�kh&E^��&\�~��íg�Ś>فj�nn���2V���0�u��'�be�kD���k�t�J��.�]��=�yq�j�7�^q�J����Cܽ�S˅�+�w҄����*b`��Hf�\�k��S�w�Y�ể�ހ�ւqK5���z/oU�x"�h���O����bDA�^��t�n0�GF��^�gUʳ�
[��]�B���g�渋cz`�or5g"���৩gK'i;��t>�K(���A�X7�vl�0�%��j���t] !��&Qz�S�t$�TŎ�Q�9��%;��{0Зj�����
Qq]3
CNwwS)QoN�=���,ꜱ���	;*�c9N��u��D�uY�Y(�滘kfs��]dd����F���\�8@��վCma�s֘(�^��W����S��`O�z����1���{�qJT�Q���ٕ�ӥ��ǫ&>�1ת�>}W	x߇���G�烺.o�N�^ˬ�P�g>��C���K�z.K�x鱹��m�G�m?�+��kā�v{:pb��oOj;u��IvF��wC==�&'��`��|	u�C���RK�����utt�f���S8U�<��K7-��S��}�v�����ѓ��z��zUE3���wn�gT�ʝ�V�/R)C���B����)����N�({��ub{5�ۯ���o�^�#<����^�e�G�(kK�U��*E�PP�\�J������T9�r����.������v�s�q����̅����[I��W������+g"���1y]H��*��	y;}���S���^�!�\�l2.Y���֫�u"�<\Z(&e�we�;��nӡ�)H��ۭ9�"���+=W�%��S����pD*�j�D�_K�����˩��P�dVL�>soʁ��[��λ��m�<������unN=R����Lmc�.TgQiG}��w&AwBǼk�mg����bh}ͦq7���ӥ�`t꽹����s.�M���Q�6h��9n�r��w�d��kYb%��E��-���9\t�4��g���﫦iϚ�a�r]�z�,��!�.��X�c1��x�r��D�>���,d�J�顟t�5�w��5S"�G�\;��K2�g}����k��w�u�nvx���{�h�Z=�|�v�WܮE픚�&
6��8j���Q�~�N��9�\���Z������R>�����R�.��]f��%Vo�RW������v�Uԏ���y�V�k|wQk�-2�x�)�D�4Y��K��{۞/@�jo6��|�������~����Q�
��q[^KzP��7�:ѳ���/?�*�>Lp�X}�݇J�t��8g��g.k��U����i�����w	"��zW��[�{�M�X�.��Yq�~��&�I����n����+��O��~������n�q�8==cu{�i�κ>=�L�9Q��[r��jw�>Y�t� �%�2-u��!|.�8��r٘)�ŧ������맾7I�]6��wI��?T�ڿ|�V/����X�D�0�SԩU=�]A�A��S!�`S�����F|������gӨ�3�u]�s�[��jL0QaFŲ7@q�N���KF�ÜmuT�Ztw,t���(k4��	��g_ړ��n�+�-�N���a�I��v���u�@\p��BG7�%��+�jٯ��Y�:sw9��W���:�VP^qx��RKG����| ���|��4�k}�1�`��yѵ>�܃ϋ��tf��
�4�{�l�x�Z���ҩ���37I���~��e{_I�g]�F�;��'�c8ġ�a�Wj�P҈�$�ux����������-�$`�|��v�Ϫ;����=�ɧ����w����H����#����3+�$]Y�=�B ��B�vWR�@��j���}o��i�o�9#k�/o�+�z�-gO��/c�^�L>|��'L�4Ms�I���Pq^o+���=R`��W�A�*�����h��y2c������W#�o'�Cba�k�&��T��Vgk�س��I��8�Cgj\sjT�GW;<�y��5v<r:6�`r��xT72�U��H�)K�E&�1����ѻz�}��(�nsF����o;������]�q�$h6�+.��޴�7�O+��q������r�HV�^˞�[����Lz����*jv�ޗE_���j�LƉ�2M��E��'^،5��V�X���+�a���ͻvx��;&'-"{�ƶ_L�e�S�����m��j�<#E���L���0T�:�pG
�e]��n�20�o}�!'C��%-�gJÝH�W7�ݛ�QdA�o9-������m��nM����4(�9��Z�>ceZWv���Z��yݣ��Z>�V����B��c"��n)��\V�����<G��������z�U�yS�<�O9��];�SV��/�11�zϋ��[�L����v&<卋P6<崸̤v�V��VW�c��w����O���>'p��.K����v���E��ͻ.1�ur�&�l۞�V�G���%3�2;��[�iӄa���t��b�u�^;&��n���rff*�f��>��zt�����/�.[�胇��K�Yg��+E.$Z>������Z|h�qo�����@��SR>a8��.m�����t�kY=b��!/Ц߯R��xvG��K�o�J�C�]�,���J����L���i�������	��HY�M}�����9���5�o与���\���Zl�=�f�;e�nQ9ڈ�0�=Μ���;���GL�Y�k6Wm8��u��'^i���r�	�q�u�� T�l8��l�k>���z&ؖ��H��4��(."���\y�w��|>��Q� ����QpD�@* ��Q��
��W��* �� TA_� ����D�
�+�* �`
�+� TA_��
��W������D��TA_ TA_�����)�� QD�wK��9,����������0Y��*�
��QB�A@�,�j�
)R�%u� �����r��QR�A!"� U!U�� .�F)Bfp�k.�R�g!n�3*���m�G P����i;j��`R@`JT`(  
    t ��[6S�[
2(�6k!!Kgn�JE������c45�6ʈ)Nt��2�*�+1��M�ZUR��m� V�M���¨�lY�d�[Sm�K6��h���h�U�ml��kd�e3j�!M4� �mjL�P��j�F��i���.�ra�$�jM��V�m�-,���
㕬�����T�����    SƌIRR@ h4`	�� O�)H�@`��h���0sFLL LFi�#ɀFO��U4hM1M2d`	�i��101��&%=$��0�i1L�&L�L�d���_��?O������5��/��UUP��YVUQEUP���X*���(��A@�_�UU@]U3����?��5��T��PU@$C��SUEUUĪ�!t5T�\h�����w���?������??�aAUT��^eO�}��~lO�o�Y����"�>�~�ݿi�����q[K+��mPvجO�z��gVcկ�YN�망n�sv0��M��V k*�,5����d���4���IdSU�P�fP�ژ ��xRSN@1STs�&Vʂa��r�w��7i�"�+��X�橚m�����y0[�܏Nb���s6���d˱,ǟL�J�۽A�Dv�CZ���	��\cM�M�E^e�yf�+ ���36�|΋T^���B�"�x���ΌEn�j郅��o.�d<�.��җJ`VV�J���M[�o��%���7�����E0آ�G�2�^�-�da#bLVvwJ�n���Qo�ussH��[/q��N�Q�l,m�]���6�D�������D`��`1�f�m�\9����a�+��<us�-[����vҔТ7�� :�Lٳ�3/%^�y�Z4RCRȫ�Kj���v�7>d���Y{��Õ�2	Vf�Zw	lCna�9����5j�B���� T��v�Ф�W���:����tn���0��b�n�X%m&��%{�\V\��0zm�����,�x�=0�JB����(L���+�\�KN-m�xUa�*Fk@H����,��l�hJr��-Ю!�����M�0�����J�f,�1�30F��[xnVV�P[��6U�1��̤��P������M4����4]l�ڨN�EMn�%�X{C�:��*�#.�0s3Ł�	���kݤ���n��ӂ��U�ӭ�Y:Hp9����k1���0�ŝ�w���vo�t�Q���e��f�\�x�]+}k��-ae��e���iX�\��[x� �oX�d��t���2�nn��
|�*wB�وЬ�ܘ�HG@3^�ڰe���j�2ļY��ˠ���:�5.ݧ�@-����5��6�Ӯ�+���tR�khǌe�@Ԗ�aR,TT�Z���[�-��I����*��Yf�z��On�|�כ2�VL�da��m=?q!p�����m�����w���^i�REN�r�mX�f��9�D�`6���Jc��ӗm䧯"�nR$h�П`Ə�(���-��xr��v��M��|��+�#I]�SiV��V�`ٚh�چ�iwdXh],6Xc\�k,��b4񈀥����.���!}O�+��x���RUa���m�D� �Ŋ��e�%�{yXYPc@�[mfA$��[1m�0�X� �Ȳ̳��zV��,�ܳ)m�Q�NiØ
5�Mk��f�4ڸv]��ge�%���ʧ�)]I�h�B�����(n�;��yy����Vn�%��n��ԉXnKт�!$"t>�a�/>�Uh�f�fԫoL	#M��r��z�,��ox�X֨�d�6]m$(EL��q�/A��N��r7���ZF�U��=�z���Yki�� �J�����yh���4u2w�nl��^��ʽ�ڱ�ke�����+�@$Q7γ��/���WjѰ�^�˷4錫�J�	
��QW,[͢y�e�Ǐ�mf�-���®�㩸#�O^C{X>�0�"�YI�
��AGv��&aw�ę�x��˫�ven٧��Gs(�`ed���k5Q^��/u��ʴ�^��GAV뻧z͚�r�����y�Z�ԕ�U�" vޡ�m���a�ՙ���:hj"�t�oU$3R���dѳ
�6,���Th+cq����f�8���+��ޅ���BY��r��9�Q��*�~���q���Y۲[����7cU]B��]nDYl
���ndv��k��۩y���{u{.�!U��E v�I�ϲ��(�݂�:�p�c���7��RX�M5ϳ�_5���=w��]g:�$]�,Ӧt�Ǥ�y�\,_Q1���WV�ҫ{�Q��f�m�������t��S+F�u4�{7�8vUve�,�CJ( �|��g:!}zq2S�O��l��5�ޥb��Ҡ����2 �q�j]E`�O�����f�9��_���M}��h��+��)?�u�H|���ϼ���������z�{��Y����� vd '�c�Gj0f�q�{lK��e��U��68`)��U���0N]��܏��@~�&i�0N�6� I	�tW;�W��Le�+��O����,*��u/j���gq�y���+a<��v���A��=
�2F,�6�^�]��M���ZN��On�)O#��j��l�p?mnr�}#��0�����]lً�/�{��[�u��M^X��ּ�y�\ b���㒦n���O����Ty�QƤ�wVV�I�YB��-]C�ۈ���̼뿗p���1`[@h�,y݆�ٸ[o	E�t��8b��ℝ�S:;{��Ò�S�V�]Z��X"6�cf�Y"A�kt=ħ;@cghp��'���^мq���w���TՇ��.�kj�\Or�޺���ę�n+���>Gpb��] [�K���F�m/;F��&�2�YM�u[�j�{���e���7�P�Y7�V���-WWum6�Ɯ���C���_af`vv0��e�N�i�����z�@o`P$�AM0f�ekCw\���r��qM�*��Y��s:�Z�GWiO�*��J��j���6�]�bG�Pñ�|E�Y�l�s���-�/�jmȍ���p],&Ma]+�lc�2��^�k7%g�[`o��}˕!���W	���6�wt�8��dS�J�<��g8�^s�r�Q�vq��q.��a맻7�K�wR�k"ݣc��j�����3y��)�o=Hu�T9W�˸T��.�N��O2��Oc�.�4��ʺ�v���1��oF�Q��G�\��0=W���Ni���k�n�j���0��'vF��rxk$�巋�����Pޅ�;չ���r����6y-����Ϻ�+�l	�DU�:�[Ն�[��}:\���w]�Ǻtmu��Ӽ��c���u^��-��\��l���(Q�����6�2Ռs0-�Jׂ�63���WsU�i�O0	��N��)�{�ά��̵�,��1Qy|�J��ɔ2,ͨK����-N^)qf�v��uJt�-�hq�<	lo�H��ռ��ƍ��$d����yS���w5�E孷���6�/
�6�)�aQZ��>5���n:.�S�=�	5P9�6��Z�6J��uc�7W`\�c5K��_:ia��֛'�	�bܑ�n�Q����ĭ�r�r���@i����&��%�����إ2�E�Z.,B��F�ZWc]���)�i�f�x	�wJe3ט�a�q���7ݤ�١bKǬ��$�>�oz=��Lԭ|�˛M�Y\\�^v�و�{[���9���k�~�wI0��l3�,	��.���{���p�����n���]"��k	r?M���M�ھ�Ine';��w�3Vx����{��vuj���b-U�	�^p��gw�C��G��V�k�T�b�	V�5%Bk����-�"���g2_���,���\�ƨ�pmE�VR�}*�iK����wg�s��q}Z�9�<��H�qC�7���ٙ�B1���k����kFywd^�r�i��['��5������Yiˎ�l�$A�o"�-�m���4��M6�m��m��m��m��m��m��m��m��nI$R@cܔJ�ڙk*Dv��;���WlR���=�x� G3Uja1e��ҧR)E��ކ���#��X��*=q�ڛ�LC4�)u�h��y�<PXh]��S����8cY�S糭=�Fd��$)6�:�nF���it#՚����\�q�.����� j���=OOU��K�w�%�q^�a����G�ç^MoVwj	`�*&	�/E#q�£�g)Hoq��ǬNՀ�]�*���l��oKE#v�8R�\�t�[�ݥ%�]����ǋgm�`B���;��N9�4\:�Ʀ\���1����3�n,rƅ��p����0�+sה.<�G���#�}�}��ݹ]VruU�y7|z��enĦ��lA0<���'W��OgC������1�������b>�����'q|��r¨?eW�:]UUP�6~�o�l�k߰�s��5��s��0v�e�n�}I=��c��t�t+��T(��0
�̠h�C���@�N�KZ�إ&�ţo}L�ʄu���c�zT�l�]��UZ�խ�<��C酠f�4{jV�]����<,�2�n�"�303.[�ݒ�����AVc����oF����kY�7���X �BB�cK�u-q�fՓ����L��.u{)SW`g;θFi��W}<Lz��h��6�F&��o�l�������e#s����mV"���I Ա���r��yΈMh&7��.Nӷ���a��0���� �|z)L��F�3�)�Z�u�K�,����/9���N����GZ6N����.�#:�o���K�ܽΓ�Q�+ݕ�S�����#�"�]�Z�F�R�m��٩4�wwwj7ϖ�h�Z�#[��:��+y^Ӻj_n�ܨ���f�WM(��=��j2��̺Pb���f�����R�E(gs܆����ף�Ӷ��:��v�A�����G!����u x�0Lh��0����̿�4q�t�g(��)42��]Y1�IW�����u��^гgr*u�x'�xQ�r��]b�:�V�j��(��t�	��>�.�ȝ��;[��C�E�Ԝoܕz�+�M�X*�:��4V>R��ѵ�*sf��R�	�䐮D<���̕��\��$eg-�n�� .�����(��o"0 �\����{�fr6�wx>(��Sf+i,K]��aV���j�Y�]`�s�uZ�]�؁��[���=ڸ	!M�rI|H��a�o�[��#�ݽ���d��U��m�h���9�].�0̴)��tt
��kz��e�#	���uud�n��J� �r���MN�y�%ij!`�Γ�9�3.Wp��k�
�5�|�f1��gMJ:8i��#�7��{Q�j�a���.J��S��h��㹡vC��M�Ն�����{Zr��ba⼬���r�j�CP����]K���u�0��S/7r_
j��fD[�]O���W��wZ�O��l��(O�z�A���Z�c\��:�t/��Hˑ�yF���:�L�FkF
=��s�Qވ2�u�ɖ����g�e������!-3*�.����G��k�X͡i`[�8�'n<���Da�9�[,Ca]���ن�P_{��B��.D-8+��5;���ƕ�B;���kT�w�tN�u�F
��oR���D���R�tK�J�uL�
�n�nIQ�$_)�fG(����+�[M�#uW5��� 	j�jn���K�,�8 �Vsu�nJ�7���2�6ޖ��)��w	
�{�R�%��4i�ܬ{�����6�}�CKݓ���;UAP-e\�t�bأɆ)��jF��S��y*��7������~����=�� B1�h�8a��tآ(�C�����cڜ>�/"�L�:GL)EZ�a74���D�-����@}�c�,�E<q`�mV��Mh��wB�:�vV�l���9V���.��dk�ҙ\��ܺ��}æi�	-�[�Q������_�y]�f���9�7�脯�ϯ��
����9P������i���-�~��K&���e�KU�r��u��M��d�'gWu!�N�U�*'/�=����0� �лD�'���.e�L�]R����E@-����e�f
V�V/�D����@�����ÆC��RF����
M�FRWIh�E#ݳ�=ݮ�|4#A��t�0`G�i�uݕ\Z�褢È068`я�[|����M+ӑ����6�w�܋�;TNdX�(o�TnL�]J��r��H�V9;�'z�Z�u�(���Ҟ�7�
l�ݲuMyQ��^I�\�$T��0浝���T�oh1�[F�5��2��7���>�v���W-w�k�؋�y�Y��R:k�����x��v~��k+�'��c�ƃ�k�+�RY0VWb\3��S� �44V�,��Bu�޼�l�y�2�ʵ��W�PU@ �R�}(������ʡ.���>�/�w�8�YL�=\��[ъ,꾆��.�4vqp�P=]9�7��gc{�n�m��5���)�]�֍��b)��!үz�SlQF��$9��b�E���A��6�^�|���+�t�5���rt�8�OO�(�=Iq���v�!�G��GzS΍Dp����$�7�[��W*�vs[�Qm�H���5ei�r�H�u��<���k�²AE���˵%��Լ2�r�E11ui�U$[���2 ��ܦ �H���l��M8�4�m��0]�^��2�ᨩ[30�K��1I�dhnR�1c�ZF�%V�pʉ1wR�#lH�0��--���j� ��Ѝ�r��$Z�Ux!�IKXH�r��j�[wl��
��0�Z%Š�!��ݗ�R�b�p�b0����n7�����܅�4�d��T�W7S�?��?ߊ�x@�<�o���P����N1%��H����ܵ>�G~y~e�;Oa�U9ሟe�1'�綧`{U!��:'�q��!�\_�"em̻�iu��6�-�φ���(ؘ�νfƸfw�CË{y��pE^Ae��0�v�#/�{��ȸ�ag��2�������}1g�z#&��k[L������z�[��6�����`YGjF�׻�W}�kM��6�ȣ�4��
/�Ӷ��ۅh�̯9<w��,n,U���^-���*{��Q�q譼��E�y�d�pֈb���Z��VWdc��o��y������;^�M\ٌI^�WI��\-9��:>����fRk!rK�ljQ�+;;G{_��n(KQ#w�c�X����6���>�7�o�/TCS�t�ַy^9E�$ͅBE��&�=�V�u�x�dT��yx����l�h9�\���v݆)��~��}���W�+�^�Ag�
�y�g��*й��?3�2��m.�8LD��tt��dV��c2	빅�;��7�y����ա/̓�Nۣ�B���Mz͍�ng�7&���7���g���P�LW�h�+|��;��J������[��৤v̊�drh:S=|�omqrz+m�����s��3�sb�'B�Z!�(�� �x$KMH��:���ړ"��ɛ`]�V���_Ηo�2�fӯ;v��&�<��ps�>Mkw��S���������h׬ӧs2��e�k�����ϱYiK@���93�m�\l�f1����mQ#N%hC�*����?�j?}��wH/1z���ay��j��+�1�r{\��=�\p��U�CIiYNo��5L������3�4Պ�S�1���QCtq���{�7[e��ӛ��rP\T��H$��L�����>����0V�p�Bsn99}4xk���ζ�jɻ'ahw{�5��9���i�gSL�FS�b�9z�}�ou��f�-y�N%ZM�w�o\�3��<e�fT1	�o�i���)�_w���O&�S)��\Ĭ����5���<S��f��>�f�q|kW�U��o�ܩQ6�ƭ5��}=w���P�%e��4�-��c3+;���q�i�jy�q>��֊�AjM�$n�צ��l�#8�a�;4��a�N�C)����7FǏ�8���Ӊ���g]�s��WZô�%kp��kЍi���{��hClI���/�>�zk<j�z�����F�����'\&��W'���{�o���[Yp�`�
��J�,�nh���a���٪�(�y�#�n��Q-^�hÄ�|���:;�����y2��LAf�F���=ȬR`���\*��d6����qbW�!����3��r���N["�Enj4pwH���H�M�����7;�ԗ��|��[RRϝ����Ġ������1��W�]�=�CN��ƹ��cG9�	�^������W�1�|������
L���?pc��=���U��L_/�6���Oڪ���xϵ�l�u�S%nf��<�r����x���q�R��a�n]'xy��Z=��NB&X��'�y2�����.�O72��	%q:��|ƨ�8�b��U����N���%��oR��E��U�Ώ�5���D�'hf���, ޷�7'>���5�ѕ	��2~�����`��ć���EI���k3�[p�B5���N��ʿ[,��8;��m8�j&S͵�������9�r��S����{��0�z���z^kI���y8zN�M�M�k�-��s퇒!9N������a�i3����@�I��>p�s+��q��5��k�� �p�96�Fm�����]u�e(#N!�R|� :r�ܼ��䂞�b�^{w��9y�eo+��^I��ڛ2�kq�$W$��.�y�
_�����DM��º��>5Uˍq�zKM�Ue3��8�r��Sm�1o����N�ev�ס�8�o�e��{N8h��p���Ա\>X����ҬW��>A���|O��s3��o�����nV��a��P���y:ܭi��?p��0�L|G��ͽ{�g/Sw*bT�4�hc��ZM[�o����r�+���^įv[�N>�l�~꯿z~������1$"�,��R���9�����3sav����Nk�B�x�A����a/kG[̉��B�$a��� ��ୱ�{X�5Y.kvc�5Ի�[�Ҙ��9!�]g����a�ս�|���#�~=�m\��v�:�G���[M��J3fwAw����
�Ԅ$�{WI���m�6�hI�������X���
d����۵�s�wR���E����^�/l^�X���>���<��������{�+@�����8�;^PT.����U"C{u�Y,��ȦCb�d��=��!gqj�TC;���؄�{��g
���,�j�г��T��Ci��f"���ɮ�2oU��I%f*��^Wk����A2��y���/,�|�g%F˝z��]ɧQ�F���X��)m��g����o0-pMT�Ө
�0Y��Bc�݀ʈN[�����]�]����Ą�.6����ж�F.6����"�a0�d$!��`�\���13r�0�[a$c��\Y"AiK�.챸0��A��$BU�q%�p఑���d��ݴ�	d�-F2E�%�	$�[v�"�\��.�Pj$%���In�����蘕b2-f��K�Q�]�D[��m�촨��˪�ܿ����k���X9�� Ĕ��_f3�w�������|�5�f.7��>��@Ƴ�;�y;í_a�0ф�gR��~���i���ܬ�|�}�D����nc��^kN��[��[J�'ɞgإ0�ì�7�Y�%�Z3�c��;�����>N�V�v{P1��o81{��4�Li�����>N;�,î��;�dj�į5�����7���{s�Tk��cV��]_��)��J���a%�����<���&WF�S��Ɣ<�>g����)��om<��M�қk]&K�m���>6���a2��w(�i.��o]�}��B>Ff�ڍm��
�n{��=��w�m��8r4��9�3/��y5lN!ƴ�C�c��gӽޝb�z��ZxѤ�8�nS�ײ��ٽ��˖���He�r�gLnb�T4�p�����>���3smhi����&�g7+�qۧ��c�������/��8�a�K|��^N�ȩp���>�ʈ�V+��w�y�W����V�p�:�����)��z=}�ҭ��v������Q�1�Ld���uY}�!��5�_5�;yp场�ku��	>��X(Ո ��D����y�sxh��M�u�ZkL�����{���]u��z��0�5֯��ٚ�מ8v��^H��.�3�y��ֲ�0�x�����+�/mu3�Xi6�h�o��rko���+��5	�Y�nV�љ^t���:�i���e<���m�o�1������=@f���s-��k�W���1�������RcA���f�_��>�}ޛj��B9t����|�N&[5��c;��u�8n���\5���y�m����O=z�Z���!{���>���˾��䭼@�Q�F9��Dx�]�~gVa�U��<3	�^���Ŋb��놞���C��=��U��C�i�nNJ�^��9�w��KN&�hoP�����y��!ֲ�@�Y4Ŋ��Q��H�e�}��+?TG���TCxф!��uץ㱙]���
C��U�Ҹ���?��!�.���Q�r�_w�s��~�
O{�>ϐ&����˦��k2�wZ�g5ֻ!�������M̴�V1)ެ���j<�%ʜ����o�:�k]�9�g�u�V�D0�N5�J祸~��Qa?1HR�W�*��f�I��l9�or��B�-fT׻;���z�ܽ�]��M��ҍw���{��֜���gZ�U��c[�q�׆���޹|�fR���wE�{���9-2�ޥ����٫+�����R���������['u�n��YǸ�O��񰴡;���K��f������QU��~ƪ1'�_;u�Nw\�L/2����o���^�άV��y8��n��oSmTkͧP��_d<�ሦSubU���o��=��Oژ�L&U��E��f1�׳��z�s������b�kӼ�7[�	���I+�P�`xN�{|��O2�--���\N�|��4ss�sүs��a�C	=��{�4֓�S��v��&!9�f؛�����ؽ��ܽ���л� ���uYوxþ�t{b{�Ax�8������j��)�>5��g'Ƹ�jV��汋���@���
�b�~<_xA����1AĞ�w����Ʋ�57�ɛƼ{!�i�U�/�#��rg��!�I�\�4I%(u7�k��$v�����R��PC�O<�Ls;ޥ��;�q�2Bйvs>g:�Z�B5��9:ѷ�i��5���{�k��Lk�ssn(a�r�7~4n�
��t�|ӹ^H���s��<N���]�����#a��:+��f��$�֔�泑s.9_ʪ���9�}�z�&&P�ilLfoo5�j��S�g�i)4є끭9����MrԬ���a�jVP�r��oݼ]�u�1)O5�b�i��y��۾8�u�k���Q$�|�������X�c�v��-������5�kZλ��vm�̔a"S���s^�~�8n���^�n����w��Y��èi�׹��h�%�!7��{�g�oSO\�L&�!~�x���'���5���B�ݞ�Z��}�~�Bd9�N��D`�ۖx��p	��U%�#��ﾡ�}�׳��&�9+N�Ƹ�������s�xj4�X��{з���=ٹ{���(�UoS��ɷ������d�Y�8jQ��n|������^/w�n���Z��;�Ft:������mv��&��ɖ��&�=�gY�5�yM�t���i�=C���{=�˻���e��ha'�;+���^���c;�뷯�Xk	2����������5~�P��k	���G���]��s��q��h�|H�y�9d�ȑ��F�����\��}�US�{د>~N�&=˫��Zm�g8�㽕�[\v�k[��K�=�G��>�q��{��/5����a5�|�~c��y�hץNM��}g5��r�{Tu��ƝJ�e[��9�w��:m�!��UmW�g�ޯ��9vx�S�ڨ�[O7���L�4�\>�E'�1*n3�VbT��߹���sR���y/ʸO4[�a/��0Mj�[����0յ;"�W��7��������v!Xs��;G�eo�����B���r�(T�1�YJ��@ފ(tې5��VT�v�������Bf���Y�ǔ��6m�V�6��&��m�$��[�Y:�%�6�^[_-n�l�`�ե�RZ�:���J��Iv8�땦9W.�m�Xs�d�Z(vpr��73�Q��*
�{���U�Ԯ�ތ�'b�6�<H2��8䳒�fE�&�˻����ia5udP��ƺ���I�kQ���#��:���ֱ=œ0����y�.�6-i�b��Sַ��
��n-�5K��]`ٔ,,�Į�k|wt
�ew��H@�׃��F����r�0k[д��ի|�Γ8�oLʾ5�\���̉x��[���˹�G�#HcS�FI�RBiG(d�[�5�ptG��6,!n�z	RA������L��ce�/�^��Q�L�[$�HB�b�ƒT����d��.�i�RJ��Yd�I�X�I%I"BAV	�E.Q̍�1%4�"�ԅF�	W!����U
ZH2���V��%+$�UET�o�^�/�b�rb&wa�K�miF?��_WԹ�ģ�R�0��q�5SHLo����?V�2�����i�r^�fSz��_.�ӍLb�������Me2璯��2ֱ4�7�����J�j�Q(Z6��҅(SۀZ�y�vQ��j�5�J���A��D�v������/�"�)B�)B�h�B�)B���m�"P�h#Gƈ��m�(|kmZP�/�!���)�ˮ�ma��B�ƈ�)B�(
)B�)B�)B��ZP�mW��Z�U����J�NMd飭(_4mJ�4D�J�J��D����4D�(R�we
P�����)W��>k1��A��D�h8ǍJ>r��GZ"P�
P�(�
e%
J�B�imZP���@QO�����ݜ�B���-:�2��M�A.D�z���0�P�y�)B�-h�Z�(D����-#A�\��y�Mw�;�3�d�=4�j�4z�rLBB^�η����f������{���(Z0�2���Q(Z��P�TJ1!B��U;�[F�#F.QiB�~��(�
P�
P�Fn�'u��6�J�@�D�j���B�-R�Ѧ��w�Ҽ�JR�Z8�3�QiB�^eZP�m���J���ݓz��E(R�(�
�h�.)B�i�[H�P�䴡J�WĶ�4D4jiB�-(
-��/{�y�%
P���-h�B�)B�������Q6���-��D�JvUZ)B֎ʫJ���=��%G��|�J�nJE%F��F�D�h�Dh�DJ4��EJ�B�-y��B�m����5U��J�Ei�(\�(P�ָ�J�iR���Q(R��ZZ2��5�!�j�&w���{�@Qh�DJ�h��-(Z8�R҅(~B������)]CW
�-�w
�h6��J�~I���y�P�b�4y�&"P�
�UmD�J9!B�)ְ�iB��%
�<����(��k��^�w���q�m��D�@�GmTE([�)B�-h�B�Y�iB�����y�4c�҅���J�F�"Q���|��6����:�<����Q(Z0��(Z�UR�(ZġJHa����C�Q�����g����̿�r���k�6@R�	j2�3;��Íf��o���@f�ߕ�(Z�'�҅(S뒋ih�Dh�DJ�(R��M�P�
P�FnQiB�)B�)B�-_w��3T�)_HF�h���(Z�9h"P��6�)B�čC�iB�)B�-�%
P�
P���w�(�3(�PZUm��Ui+mi*��q��Ҩ[J��yz��)B�p��h������-�-��Ĩ�:�%F��J�5�-(Z0��%
P�
P��|���*%
P�A�4a�%�&\�mm�'_��&����Nbhd#>J�^�-ۮ�>̿^0m�%q#\ki���k7�Ƿ�Z�C�c���u�[9��M�MB��p�8�s)�������s\�-�L�u�W!��v�����[/76@��iD��īWQi�u���X�v��!>��11�P}o���}T���y������%J�>1��^�z�d���vL���L$�6ײ�]뽟o�1�ER���!_i�齼�{5�op1�Yf�a2�ģg�}�^�+|�12�Sr��ݕ�M���N5�9��Zk�u���<��:���jcm[U�B�r��ֱ�M{ְzk|�y�ife��]z�ĭr7�k1�{��kmT��W�]r��1�>M��l������>��`��iT��~�:��t�=S�v���c�4�ʠ18�)�>��;�s���EU1�M�<N8M�kY���X�^q��{�ه�q0�LnkɁ$?!<+0���LV��>����LS�ܽ~�=+"oj�w�����%2�o�B�+�~�x�f��x}��#dtY凩�2�������{�^�~լWiC���#��X�%?(dmL���u=�������|��VkJua�bb��gY���!�:�ߣ�#�t3�}��v�|�"��������yi&<ש`wA����O���hL{���:Һ�����2��X�qs	����u;�������l���J��03��zl�DI�l��ô�����Z�����}~*�̂9���/
��se�ֽ��}�<�~���5�.g\�Êm*�QS»oƵ �Ս:�t�R���Ȃ�_�lk�>pl%D��WZ3��m o�t��u�)�['�l[Z�\�'/�G���.к2������c�����t��o��B=6��0�9Ξ�C�x���=ԬGs:D�%���1��UU��=��������w?QzF7�6F��y�;b1z~�}�	�잢LC�;3=�c#oC�ǚF�L-��0�����c�]4g��i՗D	�����&�^ )�ػn�)����+Ġu���/�<C�/G�ux/ʕ�[����Zx-�Rj�봩�Z夜���hF2�}����<��=Q㛰��͍�u_f�>�Cyn�YZ?:W�RϴL�\�DT�}Q�����}]��kƼ����od�}��:?O���n�ެ����y������e�=����n�k(=��\l\��l�����ʼ"dy1܅%�'�j�Ӗ�Z���,�n�7��a'I��a<m?DDG���m�-��Z[�����}��{uOl���&�դ/;2���&���^���(�kfÂ��d�J�{�QFFig{���}����)�W�y>�E-�[��&^�e�;i�t�(w\'����
�ܞ���?7R�F⮳r�p;��͡�X��޻82�Rۂ.��Z�U(��F�I�����$yN3PU�K�n5J�lm<aTA"v�v�4�E	���ǂ�4��H�M��f�����E��k���ݶs����gբ!��X��k�P*�Q��qӴdg��7��������c��s����Qо�3H	`�P�yVl!kX�sK��/��&��/�\��Eg2�m�y��È��#��#�OV�<�y��HS9��q�*�X�푋�4�jvqt��d�D(/�����6P�^N�Ev�H=��M�Ɔ�tS]bu��r��W��'f>�"�]�ӬѦУ"Ժ�Q����+#�x\�Mo0�r�|�z2��ܭ9%�;�V0S)dX����Y��Z@h��(���)y�$Ѐ9�T�+>�L�D�b�e���>�"�1��_�j��PY$j��ҵr4�(�MB�J.DH�DA��RҖ�Ti�Q�X���������"�%�U�$c��"�\ ���6�"�մ���"��4�8e(���K��K���"!���E*�"�(�\��7�ǝ�n���̗��Ԛ�O����������E�
*�(X�!��ٽv��G^��î����^Ղ�%�S�X�/�w�.	˄�ɩ�$$f�_»�Ԇu�+��/�u���P��4	�Q\-��.3:ƽ��,ax/��7{�~�O�O,~`~����a��)�ȑ�VJ��o-�:�6��-4�0�s��e�}�����V�����J�����X8�m������RWw��j.b�O ��}%��L����y^s���u@�q�V̎+��2]Z��|�������q��sBVSzN׎gc�:Z�8�0nE��U���ժ�˾��4DLm:��GW^����&�l����I6����*��xn𥳐�Z:�{����?9'��o������ġr���'*�n�{'.���7��SǺ�U��[���8<�c��E��ObqJa{�ee8���*-�}�g�ب���򾥰�5�-��ˊ<5<��%L��,4&�ZYzė�0�9_M�Q+{WX(����d2��Q:tm�(�_�菣�o��z�
���d����5
7�]oޙ'a�[��{�{^6h����ᓙJ��Vl5u�Pަr�Z�2��,��)�N=�d:�0��Jl�{Y�����Y�I�k��YN��X��2�i���7Z���ݽ�����2�PW�-*��Uݔ�=Ε$M_Ddo&�x���}���{�����^W�w��@w�KG�g3c^��JK<�&i]D�^E�s��]́���uk��>#R��K�:Z�ǽ��aC�^�ۈVN��k9�˷���l��(.����A����
�;���n;�LL�6y_4zФ߆N�j�%Ϊ��Ü�hA�[�V��	��">�<��o=��r�σ�<p�,�����iq���62�����͸�v���P-�ghŃ���U����~��3^�rQ�g�}�d/%^�6�ٹ���j4k�M�,���"evW�o�߳��||�)�ܽ-�� >���;��3��WE\��C��8/���
�/����UU}���z�L���B9��nӥ7\&Vzt�����k�ި=a��9�B����^����D	��l�V��Vvh�!)@���չ��O{�����4�Ȳ�"ׇ���f��a��������'�<��0��D�]�@P�Z�Y\M�)�׷��ӑ�(��;T,NX6˒~����޿{��?���-{�r�|ǙpS�޿��V���%=�x��exÚa��ݕ�r�bǼ��4��ܽh�zϲ�^�-�j��4����o6�A�v��'+H�L������TZ9�=��w5��}��粠D�GNfa��V��_n����V��u��
n	�F]f��?}|��f��F�0�Z<���f��=�3�����ެfr�Ԁ�T?`x3�R{5���W 3��i-����N�'�\!K�����
�Oa l>y+�_qB��J2(]O�3=֜��:^�Q��5v�g��kj��V��Ǚ�&L�q�]!4�BSi��F�}�tߥ�ʍ�[y�����罒Ǖ�"�����~�8����ҟ�r�6�8��!�F��$��Z���Ȧ�z'����w���M�o��|wzZ�|l����9�˚)�l��5��ӧ�����]R�q�nuh��^������+D$���ۛ\��x�����+5�nZFu_b�g�C��:�
�\����5y�H8�ʶѺ��X"n�ܱr&�"�%<�o��%�nQvr=�ѵw
`�HU��,H���v��X����i��o;+o��5n�Xw[O5Gnc�Y
f�ͤ�n�s�I�� �T�n�.W�qK�=����ű���[M=B��ʴ�H�W��6��T��ݔ���ɷ(�7�P	��l�Z�����:��rQ�8��$��>����P^l�0ε&��v࠘�(�_H�c��9��M�8��Ջ�ssn��� ����;��ˬ��ٜ1ά�f8�[f<ɕ����j��ۮ�xvT%���s7��\Qͺ J;%w��*n��O��XT�(���8��#��+��Cz&�H���g8���u;��t�g}����V�A#H��E�\�du!p��d��#DDQ��
�$�E�F��E��E!!Km��H��Y$����&�
7LE�0�#%HBIi`�F��͗q�fKd����L��F��)�*$dd�L�@�C_Bq��\�KY�9��U}�g�s��e�߫to�V�M��)�nn{v*��	w�wC�
��,��3ayoS����GJ��W-n�w/�$�n�fw�艘�F5�����;CI���s���������Dv�=�<֮s��.;�ѭ7W?˷.w��UĿ���Ǥ�{��nr���'͊A_���c�\=�n@,����}��&����(s�Q��c��������^ô����=���A���FG�).�V�l���f�w�y�#�n�4p���~������3�Vb��Q]��k�4&��:^��g�>��+�D�I����w�[�k1�����.�
Ψ��sit �֞_������e��U.7��He<og7����\����@�z�,윢;a[_�U�Ֆg3�/Um�$C�5����.��pv���*���ߦ1���dǣ=/��}��SY������z\aGjNR�lܬ��y����p�㌭�5Q�������|3��tM�#Ϝ�+��=�W�õܗ
��jg��e&�$��1o�_tw��v$��˶,{T�ɺ���5�@�[B1ԉ�}*�'��Ĺ�*��d$��^�s��o�ʣæ�7^dFy�����Xg��`�^�w�ߖ���*筇!�����;V/��kN���{5�ź(j������^�G�]��1։�	��>�b�]֭Ͱ�׼܊/J��se�ֽ�>��LE_�Oy�������{���թ��Y=����������y�9r[y�pr�1�\�l-���_{�^�~> �r,y����o����Yb%A�A�Q���W�jf�����c�#R���]J?:��
|�5�������F�0ދ<��\��E!�/�i7%�'< ۅ����j���zv0@9��±;^:$��[�n��C��3��!L�ö�7��<����k�i{�a�]})����jdrp�,�"�{)�}��O7�%��&��.7`1����vh�.�b�۔����U�x�`Px��t(�rs�&��x��}��>�J�;!���JK=�?8���{��"�EW;����W�\���UU�K�,�`׎w����`�����:�]��b�S:5�Z��Yv�5�]Sɾ-m�L3�3Ӆn�G���4jÓ&	����ϸ����/1(�������be��I~�n��'���v
�@�-���ڙ����ʙ�5��1��z�~�_s�3�ݾ������3���l��[��ce���z�C�Z3ݏ��\'��{��B��g��	���4�R��p����K�W��i����F8��9������)C�>"~��i�X���Qx�5�%��oP�ή��-�Z�in 5�#R_EL��O���k�lݡk=g"��y9�d2<G^�<Q;#}��^�����)��B��]õ���㬺gm���m�
���ت��uܬ�+��[�[X��x�^��vmbʩ۽'Ge��x��7[��V��}�}���qT^�}�4ڨN��� KwV�C9"�[w���r[t��OL���<l�ϣ��Q>��w{�3��\'�Y"�e{�)^�T��-��Ǝ���u�xi����kzK��uΛ�x��]6�<c�l�.�:��9�;z!�^����C
Ź�� �=�c]�k0olǭg�y�������)���O�sS�-�춫�ĩ���{Y)r����㆐���nvkK�-iQH�L^�$�ۗyT�{r�!�P�A,���⌶��h�J��`�ޣĥ���7�xKX~�F�Æ3{;�P-����჻����|�s�ħVT�g��9d�l�NO�d��c:HHf�C2�ƻ+	����\#�Q�U�u���͡x�=�th�3�Ir^��Ya= x@�u��|��ń=���0�51��i�6K�sT�Q-vmo[[3��6���9���2d��]�T@�Fe�%�1M���8�H�e��;s���tZ���Wp֞���N���5�EF��j�[�Z�ʆ��c{Ď��9ۏ�;E,{Yq�p������&�q����6�E���܁;����R�K�D�f����g,]�-�.�
{��+}�޸ww��ˎk���4`�BRG0'f�DK�d%H���	d�����)	!"��F8��4��*�,��D�!�b�T�"�
�`�-�V�$�UU&eZ�-I%-1d�TcUEUO�1�?Vv��S��N�N�v�p[M$��D*���O��4'�MoY�֬ �0vB�r	�mp�z�：J���u0�!�V�o��<%"�^Z�P�ͯi�~f^{��Kͯ5����Y�5Z���t��>���c/��J�i�=Mi���H�}<�.�yt-�jtk����#���ڰ��J�e���nt0�����|2����RR���g;���R*=��ݷu��%)G�CӓsmΥ���Qy�ρ������ax�7�<��xCN���
d���gxR��o&��"�'���K�o��S��I��^:��Я.m[Gլ*y[�(/T}��ڎ����ͳd�7�)���`��~��{����C�1_	���V�}@4���5���y���ʵx�z=<�W����de`yy�s.�*~����q�Ή�>�gId�!�o��~�"���~������y�M�l0�b��bsM���j?RfE*/����	��X]���̩����Z�PRR駰'V܄=�n3�9H��>�ϧ����R���^�N���6v���=^�f���G��u�y4g�U�'|�O�9^C\�(�{<gC�����˴��vԊni~mo2^����rT_?-���ru��\�u�S�ʭ����X�g�D!�(C��j��E�}\),`���b���^NE��Z����E��}�|*�l���#2;S~J��~�+ص�ӻ�En�S����3V�;��:��]�Y��~��/��ݜ:}����]��d\J���� U/a�����f_����Z�P��y�l�l�w���'��U�c���mWl�r�]*n�z��rF^�2Վݵ�bt4�����M�DK����U����Ecu�0�Ϲ�����[?'�a�"�w�XZS��P/p���F���l<�"ćV[��{���)AɊ���>;��� m !�0��`U��X��R`�BG��5��Ѧqfo�K���r3��n�ƺV���]v�&�6K,�I�X��#l��wZ�r�˭�Z/��uw�?TԺ룻�ܗ���B��k��{֎�����v>{j`�%�Y�7��vټ^=-�@��_�U�Ag}�}6�gO��w��C׮.�da���
�� 뱝k�Wf�E�����c��.�'(C��������a`�W�h���ڣb.=2�\֨�l���M+Z��B��w����o��|2����&-�d�ޅܸV�N�Z�`]�8��R����������'��.8�����&�m��ݺב�*�LE�������y��u��SΡ�潺�@�zJ7QG�#�q�pۺ����x�H�6�Pu���L�t���\��Y����}Y�=��c��r���ߞ�s6S>��C�~����N�8�I��������ǁ��ˑ]�{����9�nm���vd���t.���P�9���V�R�G�1����k�����e���_��}i��^�����d
g\��J��y��tU�
Ho��ԨI}���������yc=p�2Ӿ<��VToT�yɽ�ݩ��ґ��qI}u-��vP�n�;�� Ls�XšLj��ׂ��ŰAx�/;#���5|�	WJ���+����\��N�O6�k^���z-�z��m
WN��B��7�J%J��ky\�]&�s��!���y��s$u�#��,gFU7���m�Y�1�T��y#*�GY�^�oDt����"LK��:U�O {�o��`�����q��@�4{�Faz�x��ҧo�ttF�^\X�����{�n,Y�e�̢�]�McdW�pL��z*�U2�k��P��tE�L�ՙ��4�3,�Ә��CR7�P��;��=�3���*����@����9t�Rib���Lз�^ƭl���W1E�iĞ�}Q�>��S֮��U2E�	]'M�tV��ō��K ��"Z����H��ױX����`�v�e�0e�ʵ�.�/-ֶ�eBl垃�M\ɘ���E��w��oL;S�ez܊2�o�����=7���ns�^�,���y]�f�Uh��"m�-�$���RIK�7P�Kj�F�I"e�K#*$V�R2J�Q#HA�Tj��7!B4Y%2TEJ�DE&X��-)H����P�U��@F�&��;��:����o�����""%ww��:>;�r��8�k���&�+k#U*��v����}D�[~x�>�n�g��T�__����x���}��r�}p�$������쌋h���F����R�,�\�Ӓ*��|�~)^��[K�����T ��Xo� r����Ae�0U}J^�͙I���/%�E\��A�R�e��g�bd�)o�u�bB���5�}�uvk~����K+Խ�\�d��9r�3�b�\Wڼ9='sSޓ�1�fQ;�-\��5�}���1�?��m�ػd:���P��F�|�㿷��O2�����o���:/6�l��Uґ�$�����M�^(!������{ެ@nnO�=��"f'̀��qb���==�k=}SQ}��"�GN��2�KY^y�$I����t\��U�W[�塦�u�舊��?b~�I�^�yw�A�<�A��ػӚ��vu��G��Jc��*��K��_"�5�}ZY��jwH��^���4RƸ��Y�e6Z����>~�n��};-���5�Czo��bOڇv�#��w��٬������|��y7ֻ����{�e�ޚ
���/P���q�����~�u��Z��ܺRGK���#9ӵ�f�����7�v;��')�ǵm��OB=�̜���tB�Zu-�b�W��׍wt�X��5���oV��p�E熔=�]vL�a��+{��d?Z�D'
�ȱ��=�i.*����?^M�>^�`����4?�,��ܳ�4Q �=^è�|=����C��HO��ֲ����.����-�Y�L�6���I��yT��������|3%��]9?_yge���z���e߬���w�	U�k ¹��<�.�Sա.:R�|���V�]OJ�٩�����6�g�n�" Neu�X��{K�\f>�7�e{	=��5�&�w;��M=����b��[��ޖ�ue=c�Vn
��v�%q��u0cY!X(IL��i�m�j��d���0��7���z����j�ǝ����c���]���=��+԰�1�D�r]���')���[{��z<��j֮�4+�qg�k�x8��]�N{X"A��<��B�Q��=j�����T1��/z����ןOq��Nf�̐ʽn��T��{V��-���l[6�a��B{��}��������?N0.�L���Lg������3��5�,��R���s]ye�^���;VA	ĸ����׻۲�t'�[����l�_�+P��L����V��[�@���R��y������N�}�i$��"�t|�ӇcF�>��$�+�g#,����s�C�Y'D�6��E��M?DD+��F���MϽP*��Pv/pCݹ��<��E��崳��_��G]�e3:�3\H��{3j�V������Hy�~�:0{3-s���d2�_<H�_� _pU��{~O�j��k�0b]+�|�����Nw�Wmm+�^�~���T5�S��腾���g���CNA�'-깃��O�US�{�~���ǋ�`�Gw')BJ{��y����2�_�TLn�s��3},R�_"}��׽Zڷa�Z.��OO/-�t}�S���y���c�����m8nF�fX���� �Q٢���v�)�D�������]��q���'U�Y��S����+����k�RJd�.����\kk�e��5�:�bD;�cs�"�P�t{-'MP��x����s�bV%�R��]��}JP�|s�Q�Ճr���gCi�%G܏Z���:b�w�2p��e��#n�� 5	�C��0m�6[��yzZ\On�;���^C@N�0@����p�(���AJn�p#`�S$�ڐr��o���A�r]_ �o�Z�+"��,m`
�梾Au�N�ٻ�7@.��C��e�4�	�Q�S�OW��h�0�9Tp�c�z�'wj�>J���٩ۈ�Q�����
団�fm%��.��^v��\�,֗؍�˳Y2*�ț��4iyS,RA6�G��;��b��S�(4��.ƶ��NS�tSL�]��o��2���Ҝ�E6�bܫdnQ��ё#���An�Hբ+v�	w,m�Ʈ�-��
�G�/ea.7u,�UE�YQK�䐶��K�kr�\jBۗM�V�TV�F�.A���o
a�b]�l�E��cJ�j�$�P��DI\ ���B䨖�H)$nJ�����8���������4ҫB�@i�J�Q�fD��IXm�m��D���X�.��mIZ�n�X��!�]�E��m�� �@-	�/dC����.������}}�{��Ӓ+�rT�XΉ��m���&�lK'�!�f��SXO���k�Հ��ݧ�x��8�j��u���>Q�$ �ϗg�;�����?�)�c(/k������������V������Ή@���q�\W�&(�Ƽ�
w�nyDՉR=Y��1�9���n����w��\��>�꯳�OO�U�s{�	k1�FM�b1��4}֨0�*��}w^����^f�i����Q����q%�u�0g�3����K�,���s /F�EbUK����9����ޔz�VE��򜍞��u�,� ��(iRA�w;(?`oM�YN���e�n
�LteU�w����[r�Z�t�m�<ZU�0s�e�>�><;�)�ս����{����MuP}�7�c��=S� 4�������g}�����n�L󋏺��G�<at�.5:���R��[�ͧ�n���Ӻ���k����ԛ��9��G}u�ߠ�1�R2�Լ�����lT�����������x؜k,�l��9�θ�ZI���!Wwzcg��me�T�mоy!���l־y�;�{g�Hv���ݟ�ܝ��� :�����q��EZ|6nV�]�/Y���Z:J����B�V���#[���MB��������Hʽ��L�.��1�_��p�����C{���g��83��@�,c��IRR�����ޣX|�w��U��#������j5�l{(A�o{F��.��;~���7�71M<Vn��h�7�w �^��z:N77ފ��2��=U��:�wz�tB�1Qכӳ�ԉ*k��#�}��
��S��x9�dߗ�I��a�vc����";*F��א��&����}��L�	�k`//��<9E�޾�����W����``�����sb�+�Ł@����.`���w���w���5��<Y:��qW���E�&f+9o�lр�.���Y�[zMx��}]��n$k)*�7=�X�K����jߘWikô�!ayi*��t�[#�M�mH^k8g#�[��_�͖z��ጒϷ��s26y@g�᣻8#��9����J:n��������V��WT��,��3��<�T���͵\�Cp�����X;a����M�R�}~�jk�z�M�I�qp�^SC��+W�V9��f�^��3�b�| n�#}ªK�F8�9�vT=SG�m����oǼ�Up��������Wu�G�ߋ ج�>5������r��	�#*���#7�Q},��P����2;F�oo���=�d0�9c5���QԲ7�k<�f��/*�X�G���h��)
)���)��y���v�[{gn^[�3	�G�9A�PZ6�R�\�W��|����u���{嵵�M* ��w���W�ʗz��,1�V�zV�.�hCƣ��Ơ�앃G�c��;����E�}�&z!������[囙%\����yM�J������W����0��p����V�R4��������W�M�]�ܟ����W0%qk����L#�}�֮bx��4�T��Ϳ�C%�W	 x��{{�z����{2�U�ٖ���ؑ��5�ޔ �ܰB5�x��"�D~�]P�z�n�d�7H~O��N�m��)��k�a��b����*w��-�⯭�dt������^�� �Cn�r^Ԑ�wv֫m��Ó��c��Q*�l5x,Gmm�YY��*Ԉ��#s4�PiY��[�z��m���X�r�
P����K�x��ܕs#��C��l��E��v�c��_6p�;���mck�����Lv[���ו�L#�/M�+*iK���;�>>I=��}�l��Ŏ����B\�0���r��KF��(7��c��N�C�ݾ�\��1�!h�Q�r�G)��VƐ��{��˗{��fF��uĭ�gEktYh�z#������jF��E��G`Uihf�1dr�!1�8���t�����[r�6�+6�8��Ok;~\��[�j���������&�YX	���mh[R,.��ч��h�i��2�Nkm��éL0��"�=dH��=�f��Ŏ�B)���nk�9��4�E�&f����m�m �DF$���V�HJFڎdU.T�E�UH̤ZU�S�[rUH�"��)���DQQ���Z���"2�n��!��-* �j�4���Qd��%"F�X�cB*\���V��z����=�{n;�k��(rHo"F��T��ih��I�s*��]q뱋���;��:�kz�ټ�y�[|q��;Ҡd��tᳯH�[�V;n�{R��mJ��s��2;yvE`'��b[Z����ޛ�Y;�;�u��'�򎋊yw�B�Y����w�:�|�^>�]�f�+�M�q����K�)3�ԝl8!mM7E�ޮ�/��r�Tݧ[<�����Bk���n��y����U+8���.��Ik�)�J�u��1r-&�C.%R���f��$�p���{�x1�n0G4�V`��]�a�0��وuy���^ռ���Uc$���Vs��a��F���=ɞqIc�\=�nlS[-�51��žI��VI�u��K�5�� �������
D�ky��o
/Q+4�.bԅkm['�!�"�ђߏ9��v��w�}��e�ͅ���ؑ x�;�fx�y��WS${ɩ ��[o���v��k0�r�pޅf�b�W�ʡ0��)����Ɍ���g<�r�y��XN[�f)}���[��~H����ֺ,'�ޝ�������ckuo�=hJ�xWgnߵ@�+�O|A�96ߑ,���9�
����7K�JøL��?]�jv|ȎN
�mdJ��̶ː'�fQ!{���6]f\�Q�������lE��I/cť�:����uU�����++��k�c�H�كcs�ZK�^z��y+�^����=Ȫ[�aG�6��Ǵ�N�e^�<�[���u���b�v�Fޡ��'�m�2�^�(��Oy_�nX��V*և�8�wv��c���W&B���P�\�]޼ɐ{y�x�׶��e���N�N�hOd�-t�HM}�����u�{f�R�������P���#��9�sє��Tq�e<y�w~kH tΘm� ��)`��#iӡ߹F,�xr�Mw���R���lu���9��uQ��u�o:�
~O�n`�DGdBR��m�O5p�$r��u��a�c�-4�N�H��Yr1����qÒOW���[dƟ�M��=��}lMz,ǆn��w�ӵm{J���S}�^�����Bq��q�u�z��u�v쬯<�RcNf�~zv/N/O�w�sl��m������+���Ka�����vپ��1r,?��ٲ!���iW#�Z墤���Q5I=^�_5�E��@�R4�����+!x�1�����cK�$	��P�T>���7=�>�+]��Y��S��Lv�Ή�6ea�Oa÷�����B}YFi,��oiv�y{W@t����^)	��{q�d�]�o�`��4��a4b���n�e�	�cw���հ����a6Zf�Vp��D���/��]WS>�ك�k�X�=�+g��Ww;��"����Ow���RLW���Ё��3A{�����+7[�װۙ�����[���������
��Sتu�ˏ�R�5�7�׮x�vp���:��Pb�ڎ���Eѡ�dv���-��a>�J֟�E���܇��Zr�|�"���44�\!F
�v9���oy����ݭ�p�Sħ"Gm0G/n����NM�8���"���
U�J�R����F�~���Ǜ�����3��?3�[~[�/�챗�
=�i��>W��x����/[���?μ��J�^\�K�T'.3d)��Q�:�U���y��$vG�T��T+�˙N�ѶT�iM��ŪF�ws&T^]f��kʴ�G���i��u��2�_kS�;Y�#Iw�p!�6���ZA�1��ݬ�����t|0't��\ze+u��4���U��DLY�6�*<�A<���-��wS^�O�ٲ��ݢr ǽ"�bFQ�E�A|"��J��R�[�e'C���6;.��hRw	oSUA}��E�#��!������o�M�u*���d����]�0�s�l:�Ŗ�-��Q��̨����h�G7s���:�R�$� ����\ۉl�3x�H�^9�Q�gQq�ы��9L,�c�[udI$)��;!�"�<ƥ�C]ʂ�{��{*p-RrǑ47�ΘW�ꥻ�Õ�]UZ4y�(
�B4�����]���Ĕ��-Z(��Ц�2��JUR�!wv8�Uģ-e0�"V��[#DG0��!QQR�]%�h���k0�"�b�)�˄dd���KV�&sw�H�+i�uff������-���a��x�e�l~O�e�y흪-�a��D�u;�򻣉7��>��cR~���d�}�2���.j�~��sn�R�R���sG|�ܼ�WE
�M��~?f��ǖ�FLٛ����1��g�iѺ��#�ݎ��hy��
R;�'�wvQ�+H\��n�6Yٮo-E�SnR�i��f[{����^f�E͉��-]�|ќ9no��z%JǮp��G�^�x;~>�Fg�{g��E�⥧��?g_b�w����N�ؗ�r�tg> uo��� �,��C����e�hڎܛ7�p	�wI�@wq.z����ݬ�L�]�X��Ct�Ƒı�nv'�J��ji�"����[���9�t�{>W����F�ax1#�P���/9dl�rF�������=Ɲv
��/y4H}3�Of��q��=��Wrc��,rݾ��/�O
���� Ԫj�iX�m�y��w�i�<F}�t����ÊVOK��o��αz%b��ͽ���_P:1�1ArD��A���]$�Y�� z�G�����د�#yʦ��d��G��jƵ���>���ƛ�����s՝��[���r��K�n�sa��٫�+.�U��_���U��\�/j#��1e)m�<�q����������-b��^Qb�M��C�k#@�Q���vؐ��n8^s96��c���3Ǻ�(>8��p:M�1��\�����=g`�Ostn�odorGK���qY'��`Hgd}�����[��}���̘���������{��9�ٓ��b�B��t�m�2�,�u�.�u�'1\�S��r�^֊�E�<O�^\�S��D��o��Iy��'`����cRԐ���N�Ô2�g�)s�T ��Q���r���R9D4�Y�ɜ{�^G=~�1��Li�ټg��C���sw֢�U`����#aK�t���H���\�J��}���<=�F[4G���K�H���j����NPpQ�wrS{Н���rQt՝��Ԓ����l����7hO�7�-d�A�;����,�7؞���5�ep�����k7ߥ��:?T��;.��҃�alB��-/w�p8��<.G���3nAܸOdkOz��<����ݣ�Y��pU�dd�[���$AF��oQkv���t|�6�-ɉnk��Fwo88�J5)+=U�{���i~W�|0Ek���~�\��
1i�_v����\}ġ���z%=��Ii:׃�q���{�u��_N�k�'mE�X C�4���~�=�o�Ӣ�J�ժ�wW�B��X�qk����m�d����M�ە�Ln�b�]L� 2Gj\�Q�z�P��wzgd��hr8Ԝ�ڻNe'�;�����z9�X�9��p��e���]������1��7��aR>�	��X�0%�۲��S���v�(�������u=������dg��{�~�e_�� ��*�IO�`�U��('�y��~|��c�0�w�{-����m:+�qNe�.)%M��	,�<~�ei��3o}t�裱��㾿���^�;������ �+x��#=��n��&-���ҧ@�㽖������ig�2�⌦�z���ܚ�}jzy<���y�������'�b�*��ʠ*����������j�t(*���	�H��&� ]�#�����?�`�/�!�c�.5��
��";�HJ=B���C�%U`0��꯵*�����(_�ʮ�o���w_f����x^�t?�Y�3��g�@���o�9���|�Y��]�BS����kyٍ��
��?�U���]���J���?J
*��� j�U@ƏشR�*������������3U�5V'�=z��������C����!� �������a��@����@�+���hh�������Sʯ�V���	?m�}߁_���w>�~��Y��!���@����^�~9�'ۓ��n�5@UU�R�裡s
�W.�Y3�<�K��y6��_^�`�~𠪪�V������}���iU�r���z-|*�����|�:}��b���������(�����K�e>�0jUP����_u>�������d2\����+�@ h��_���Oҿ������?@��>}�U_����g��q�������i������|�
�!��?�UH�@UUU`�a��UP�����??ڕ��%W�`c��'���N�W�d����,(���5Z>�F�|Պw�+�wEUUU �U�U�b���:t��cRUA�SUuZ�?���J?���%�a���(*���a���� ��~5@UU������!O�_����G����WϿ���?
?��Q�UYE~�����J��_�~���������AG��u����������*���O������Ģ�_�Q�ꀪ���F?�;,����G~߇��}Ux���~��g�2U6'���"U����T�Q�~��C���:���g��?��5\�}�~���j����>���w������������}�������zg�����!���Q��ؔ4UU��J���?����'��M���젢��ʫ�?2�ѣA����h3��J�	Y����+�E*����q ;ꣿi���w$S�	 �S�