BZh91AY&SY�͐�L_�@q���"� ����bH[�           x� �PQA@	��5�M  Q�ֵU�@  h ���(
 (��4  � 
 �w�H�-��V�Vƨڔ1ZUV��dR� A65��SJ$&��D��̙�5�Z��շ�R�0����Z���;��hkpuE.�A�n� t��  ���j�H[iV�i�F���Ph+V�S � v�)@  }%)@  ��c1������Y��WX�
ڪ"��+��e���pZ�����JЩ�(( hU&�hh��|�J �/�Wݾ� �=��wV����^���s�^�ltz�w�QN�{�>��h�Z��8k����[����-ރA��t<��������==
�����{����wB�E��H�ITo��R �/���\��[�@�{R��W���U���J��wcn���A�����W��oc�������{�wc�)�;���uwn4۳<��mJ4<s{��=��^���R@ilХ��R�ޡPz������k��o;�A������/8;��uN���{���kN�}�ϕ�ݪ
�I�{�4:/c�=�����u������ww-�:���hY �@6��R��n�}�E)GE�{��G@�;����+JN��t�j��秦WM�=�����Ũ+Yku���PkCN��4���A�k���Y�[���� �!���44�
��� w�S]:�!�h�T+B놷uvPVn����
{�����(v���u�.��l�譶��n�����@��8���.�;�@�+i���G@�Ҡ���R� q��
�����t����g�$�/p�$�湣C�s�h�$�{ޔ=��.�a���Ĩ%Wxۃ@�8�hQA���-�l>|��� w���@7�rM�m]}�:�,�{Ɣ/a�]\��8�`
�3����*r���Um+4:ְ��sJ�.9�l[P ���(��)%  c�z��UJ;��uJ��<(��<���U��^��R�U����c���aP���F�J�YN����j�B�d�@( ��Se��_>�R��>�&\�oQ�U-�zw���V2��T<s��@�K.�U �6�)U������J]����w9U+mx�T
�   : )@ � ʔ�2b` �F�& ���*R�&A� ɦ�#A��d�SM���    jx@����O(� 4Ѧ���JH5* @    I5�$�&�F)�Sj6�f��&�?/��'�ʠ��2��H�T���͚����ݸx$�f�y��7·���n�w�̫�}�
�����T� 
�s�H
 *�A`��3�����?�?� *���I$���U ~���1@E�����x~Lt��X��m�lb�L�%1m�l`���m�`����`Ķ��m�lK`��6Ķ�m�l)��m��-�m�l`���`�LKb[ؖ��-�Jm��&�6Ķ�-�lbS`�L`��6�-�li��m�bi�l`� �-��m�l[`��6�-��6�)�[ضĶ�cm�-�l`��6Ķ%���-���-�l`��S`�L`[���%�m�cl`�ؖ��%�m�lKalcؖ���m�lb[ؖ�b[�:b[�6���-�l4��4Ķ%�-�l`鶒���`F�m�lK`���4��L`���-�la�%�)�lb�ض��%��`��6�-�lb[�i-��%�-�lb[ؖ��-�L[b[ؖ��%�-�������%�m�lb[��1-�lb[�6Ķ�m�al[b���m�lb[Ķ��Kb��Ŷ:clZ`���m�[�S�%�4����%�-�m4Ķ����%�-�l`[ؖč���%�-�lb[����-�l�%�-���-�lb[ؖĶ�1-�lb[ضĶ-�l`Ķ�-�l`���0��m�lK`[ؖĶ%�-�`[�Ķ�m�lb[ؖ���%�-�l[`�)��0B��[b�*��F؈�b�lTm��LA�4� � ��U-�lTm���E�&�*�Z`lPm�lPm�-�Q� ��SL؈�Fب� [b�lm�lQ`�l؂F 6�F� �`�l@m�-�A�
6�2ؠ� � ��@�*6�F��b�l@m�� �`#lm�-�Q� 6�F��M1m��1�*6�Fب�blm��T�1���A�
�U�
6�F؊�b�l��(���� blm���*��� 酱� 6�F��b�lTm����(6�F�	LD-���D4�F�*[` [[b [Zb6� �
������ �� �(�X��*�Kb�lT`�[[`+lDm�����U�
����-��lPt�KbSB�
��V�
� �(��
`	lQm�.���B�
�@�*��1E�(��ت�`([ ب�m�1�-��"��@��� ���@� [Ŷ%�`��6���-�`�-�lضĶ�t�CL`� ��m�l`i��i�lb[ �-�m�L�)lLB��m�l�b[ؖ�Ķ�m�lK`[#ؖ���-�lKb[���i��i�l`[ؖ���-�lc`��6Ķ%�-�l`�٦6���m�l`[ؖĶ�1-�lb� �%�-�lm�b[ؖĶ%�-�lKb[���	l0m�l`�����-�-�lK`�ض�Ķ�-�l`�ضĶ1��-�l`�ؖĶ�#-�lK`[ض�-�l[`��[غ`��6Ŷ�l�ضĶ-�m�l`��G���F���\�G��5^�����t]Hp庣�V7AQU��n��ﶪD� Ȗ杂��w-�[aj�����
(4]��lkeki�W.��Y�T���X'��*����j7ꗌ1��*�{4�e-'H�\�F]�T򒔎R���Ud�B�T������-UɻQ�M�{Cp�����W�rwp�f5*Pږ3-�A�2�^�vӖ���ŗ����D/l[��f���0\�LX�W���+�Ǵ`RԹ�oFK�F!��iDjw�=���fLQ�S4k6� �)�TlV�0v��Y�#���e;Y4���ݓ(�p�#F�����(G��CɡSN�Y�2��d)�4��T:I#t�R5`۽d��V�0j�`3L�a�oo���̪ ae]�f5\��H2��e���n�HCYJ����yX7#.5t��FҚ)���"���uY��+�B�Z�2��� ݬ��̐Jv�b\q��̺�9�{ʄ��f��N�ꆖ�̠^�b�i��%�wZieU�4]�]I�1�xv D�n�b٪��CT�V:5�P�m�WZY�J�f+(�yChn
'n�G��dc��T�W1LM��f� Rt����,���M���������Ȫ���aT0�(*,i� ��Q�Cc�uU+&�5�e<�5��woFHn��{j-�Km#�H��R��\�w�ʈJ�Vl��U(����OrYǹ���۩���U��l�8��aڽb�n��1#�롕�ʻ�.�C�b��)�u��nz��L����[ɗ{��77�^��M��aR�x���6�M�Y�]�A�&s-�rX�4V�i@�VD��fe�fLy1�yCGo�f�9�-�岽�%�2��`�fZ���{�Y�*��,��pf��{���*����q՗=�^n�%��։�W���wJ�5�%�I���.�e���AV�]����t�TB�ZR�,d�L�(H�����#�����Y��s2kY��lS�6��فPۤ �CoF=EeA7"�S���"����Ψ��i`��`���@�ۖ�^��,�iE���.h��gm6��ʷ�U�͙p�!Sf�0ND�YE2�6��a5f+)\��M��-H�B������Ia�:+q%nb��ɽL4`I]��$�yKN%il��h�^27�3S��4F�ö�:L��SD^-���rf�d�kUe��b͑�)���zF��k[s4R�U�L��b�"��PZ�{���2���Cr�	YU/`;h�k���S�,#�ܽ��J�e^f�`��GCͲ<��ScT�zueז��{��q׍�/H{Z)f��Э)�zu��Yy-�亴�2U���W��B�`�b9R�*��DI�9B�#��7f漨����0�F�l��P��U�\�
�+��i���JEӫ;I���؅���] *M�`"Zf-ݡ(��X�+�#�3Lt/QkpP9Fߡɶ��Q]93w�Uv�ܨ�l��&Դ!�U�/\ED�mPa�Y׷���};e��B&���Z��
[jW�t��A��]N�^+3ʞ;
"A�o6,5V/
L`f��2.L+51j�܆����Ȃ���-R;E��-��m�w���wmT�Iܧ�vD�a[���p�m:���D�ee��j	�a�W��M�F�ݭ2�L�Ci;�:��Ui5b&��,!KƓ��A�1��e��R��	װV�nUM�qjR�Z5�E5��`�#�TUEx��0�e�CR�4�����GUDd��RJ��hṛ[��(�%(4�x���I�h���2���a�䠎��X{�&��2��U���m�
i�5�t���ن�^��#�ʕ��VF���u��͡��n�cR�8`M�NIUkn�l<2J²��׺M���f�DH�����F��`uwy���mh#4I���Ɏab��8�PVK�K�Za�	�L0�
�^k9�!�nֺx�B#KF*����줅Y��&�-j�"d�Ȧ��X%�5[�K��%�7lJ0�
��������L3�^�zb���7h�^��i��-/�r[��6���p��ZX�%c*��t#/V���T�D���N�nV�s�ܷ�b��{T��j�VYc.9�V�f��7x���\�5�U��
�7I�c��F�cf�K^���J��ZT��RL�n�U	;&�VXd��,*v`R�Q.FX�<8)�U��g(��z�ݫ2����A8v�KX$�㻖%�Yi��4����Tb���k�^]�����eN(�j����A���rU�ܨqm�.nV�%թ�^�E��F�X;a��%<�OjyB�l�T��[J*Y[� qi��×*��v!*�PUdf��V^��d��/3pj����<"PP��PիT�e�W�%�!�J�튼.��t���ni[��vM$�v���U�P�
�j,\F"�l�Z�,k>�Vl�gMe���)�QͶ����^�&�C�t�s5�5*�a�Om�&�$�(���&0᛻�\�q�+֍�4^?!o&�{��l4�Q��H�۽Y���&B���YOB�~9������߷^M���Q.h�n�&}5�ٌ+8�y7��8}b���bݔn��"�oN5�U�^�˘��4�a(�&"^�v��8f�3�xM���kbOST�K�v��4�UW�������9��&n��L�q�,�H�,.�P����7Vl�ͬ���R,!��Bqh�H"��Vn�vi6Un�z22!a]�:��KQ	��nk����ҥ=�*�wF���0JT�ɉZF�֚�V]yjmU�`�2m�ST�P��1Y�&�꒴l�Y"��=�ٺ��R޴DNR{7q��F^��:��D��t�9��U�Y�Z��+�5�wY�Sy�.�j�v�cITf��*�۴O�N��f`,��Ywꫴóm��ʸ�)cIT�q��gA'*U��J��լ��]j��/��J̷�Yv���[��d��35][�9�&%�q�Ea@�.�Z��K�K��HR���)����-8��-v		fF��j�][����P�Z���ݴ�͚$ڑ70�,PQ�����8���Y���5��q�@���t��@�.��b��q�ҬScG\���I֛��y�Y�A�9�5ێ�l��$a�$��ʵ"l��7kr�L�h��Ŕ2�Oʑ��F�P����/u�"^zj��p�Kn���6��[�E�����jR��x��"�p�wPe�l-^��&�5��-�����v�kX�&�ctfP��NnS��T$���Ew{�-�;ib���*��R[�Xѫ�*����e�"��.�Z�-�k%�ڔn��o{x��=�W.�T�n���*l��䪕�茰s6bʎ��61�$��m+��Ċ�����J�ݽ�[���N�
�(�����e��n���,��7���!˞�B
�t֍�Q{Yx^nV�j�7v2��p[&-�
nD]S�p�\pf*
����W��vm���X���&�8S�kEѭ͸����F�ĩ�hf��Xٳxr�"a�)�.ɦr�bY��i�Lr�%Z��ei����mGkN�t
6���.J��2���IL��	�r��(���%y����+3wn�$��`F�+�jyUW�u1�/e�m�L��9�F����¬��ut�ʅ�yD��V5��Lͅ夵�Tj�mc���hk�&��O0`�yB�EU5ٺ{t��v���`э�I��:��Uʖ&��5VH��)��V]�����]`F��nU�r�I�Р��L��v'h5D�RB�˺�iC�)��1��wt���[z�Kr��n�/�ˎx�~��hÄ(�c��Hmth�֑n�;0�^\���R��Q#E��h�EU�(�C��4e��i�i묥{s
�Re�A5��\
D�+m;�ѬRM������+v�T�^�H0\��xF4NL�r�jQW~�eX�m�X+&�JءiJ�1l�4�W�RK2��m��8H2i�d9��R��X���U�1��壂1�,@��=Vf�&�f٘�E�.�'{y�ɲ�Vͺ:�cܽ	��&v���JN����Ha�2�1+,���ڮ����-͌��]Xd8Vk��(h�3#�RU�D�7.ߡӲ�]kcf�ȶ�m��en��t����%���$%1z�V���bJF����f���bv�[��9v��v��L�L�
d��u�U(�u�U0mXo\T��V[r;)�����mYyکWk�2��s}���֊�l@��-E�W�!�ŗQnn]RSk4Ҽ��Z�\u�R�8�[CG���X$��7&��0X�p�KhcYX�M�t�6��K�c\05�*']�VU@�m�5j�U;6��P �qL&nʻ�(J����+J6�LFC1-�aUP��>�J��d��+͢�m�B۠݊D5�Ar��ʌ�2�.��Ģf1�H��n
��,�R�=ӏ��ZN'p;�H:&�m�@��=��.ueÖ�n+�0mn�fh�X�)"ԯh�,cp�#���f
4^���xw3onж����u	�~��n�rXc2UCIJ���Qjظ�x���d^\Eз�-߈�4���=�j���$/^��嗔2˼���;��R����_4��4��B�٪�������h�U�u�D:����9~���P�V)��u�
�FZx�I!w*��Yt�^�Q�v�! �!@�6��ݒ�:YW�,R�9��*�2���.���53��ȈT���<sI�6r�#!�p.����SZVe��T٩�X96��TJ�h�RU�)����2�ߞ���Y�m�F�DL�մ�cB1t�[�����v7^mc��)h8�ͻN�;#�j����eULV�X����ΗR�ܛI;T��M�d�ӗ%�q��Ll��v��w�S.hF�f`��;(�n�V�����D���Ws�U&c$ᬧ-�HҼy�=^Ÿń��*�K$D�a!e��)y\�9�LJ�ke�+E��V�؄V�y�94۴3u����-�K��v�
��ȵ��H%��z�Y4��ꥄr���ŹN���r;�ܫ �Ph�#K"��)u��������ځ�f1�ʺ�f^4����ͫ7Gh���,x�n��b����H�ux��\svc���/
l�mğf^�QvM�H�*�ٔ��k�)թD��w�¥�Dh9��$i���׸�;Uu@�͚�]�<����-*�~e`D�"�sJ�y�o�[�u��#1�s!�w���,�a�T��h��
B[ܒd�V
ћ���
���!�(�
�R��Q�'����YSH��^��cS���Q"��Q�6�&$7pm����F�*n�f�J��rS��\fěx*�X2����]�ڲ�朷̐]-�A��/+}!p�T�dx���[^��X�������V�ja�n���)��f��t��J�iD+hnފ.�[El�r��U���i�
r-ӕe̐���{P�m�4�J�0.̛���5��A9���&����լ�	�
���F]X��i��H���s֭���q��q��&ꎉu�w��du�╎�.�O*���ە\���l^e����*�)���iB�E�Mՙ�����kv���e�ciY�N�� 0�xi���,���XN���d�����^`�
"/~Ad���lT(��9k�*`���ł�L��9e8��7RК�z�[�1�L�8N�i��v��,���A�R�Y��Ӫ[�-yݤ�'�1悤�
�ժ
J��(������fdj��nݢ�+i�=��Oo6�!U1ɢ�m-�X�����3AE�M<� N\�ă@�2�����UL8I)���IoV(#�+4Jڲ*����Z�j�U<݁m�\";{r�˼��˴��PIܤ��$5S4nԕ���N�H�LL�jѶCص�,�80�&�B�����E'B96'(��ʫP5G*�fՌ1)�FK��kou䪽�ع벤j��i��ïg����قK�Ꚇ�{m�j=Ke�\��}�V� ���J�b�S�O/��U�H�92�&������tyn��A��ty8�-4iW$ֵ֥֫�W�Z��&��y]*�mm#u�M%Y;���-@�r^k��ݜ�ْ�5,F3�2POe]UDf�T�t�*�m�Ir/��;19Q̥x�S�R��Aʷ.��]J�<����vk)w+���Kkf�d՘�*�1g)�b�:RҊ�v(�rԮ�`>ޫܽp����-���5�&��dOU�����e��uKR%���\J���>�=/vc�	�bT�����-.\�r��%K�i:ĒS��$�dU��^)i��Z���R�&�s�Z��"�bU����*ı58�y�YgVĹU-�-lGIǖ�2�7`����$��:J+י���)o�|�&���Q\�I'�\O�N��ԱmB���"�w.H���5 \���7���Έ����]����X�)iikD�Hڸ���]�b�T��4�}}��5�"D�4�7J�(�M}
[PjȻON�\�F�9{���U��U�J+�&�Pv�p�J�wUnDLDu����S��UJ�+J�R����q*Ӆ�$�l&R�.B�^+�qUm��kuU�@�U]���\R��g#��M=�3:n�IZ�*��Z�*�]��A�[JD�l��@�'%�Νu��(��co_��+I;9vumP7��R�S��L]��W�$�RR)�NeL̭�Ÿ���J��I�M4�R�+��z�#JFe��v'�Z��2�-YK�R]�Y�bQG��])8k1NU�j8���Ra��y�kw��6�V�ڢ��֖*iE�tywp�p�=Q�c*�X6��;���:�҈���%m.[J�;Z���@y��[�2�ib|���j8�mh���j��GnK��E���-v^���U��J��@�]J$s��5n,�"Z�u�5w�a�{G5f�.껱lUQ8�/����lږ'5�j��KR��M,{YR����O���v��u�˥�X3U�u$��j�<\1b9�
z���ZN*���:�-4�K��5NJ�i+���b\��j�`8����[��ߞ�\�>-�� ?��J^��`ߏ�����~���m��m�ۈ�oS����ek�*�l��x�3Z��M���Y�i��1�u�6�q��\�)��������Kj+�o:�l�.S.!��[[���+p���n�p�Ҏ�T}s���sHw�-݆�[�-͋�-��j�\K	��v��b�+:�K���[�Y��,��z-��ݧ��N���5e9�"��Z���Sq��YK��e����F�n��$M9�m�ul����^_r��	�SQK�wJ.�J(8��ӳn��IB*
@�ٛ�Y�h*���E� ��jB��:�Z�[�`�թ�U�f�32W����˛����X�t�"�
�uqx��<����������C����0C��m�ҋ�T�;�X�#z�	Za��"r�����惃Uv0j�Q�%���I�8��1"^���W?\eZ�m��]8���#��U�j�[��{�����ϥraӜ��-�ĵ���G�r���	*�3/�+���iϛƨhvYD<�͊S�SJN�N�3�*��W��=(�ȶU΍ɋ�I�Ȳ��Eji�μ��ګݮ&X����^���������+	���h��R�\;�y
cg$0ͼzI�34����\wU��rc��������*�^є[M�:�ۼ�^��(�F�EN�A6pkN�2������\�Y�h�2�e���0z�6��T�NN����TS��#=�kD@m{�j�n5x�E$��n���Jo�.�^�c2���y]9c���qwd�A�$�6aɻ�r����L,�dU��Biٺ������E]1ؗ�va�E]�c��X����g]Qxr�����Z�R�&�nrw�q�˝݈�j�kx&�e�N�q�b��љj�ʧd�B��vgU<ۼm@A�tG�~��9Y%���	����pғ@a&��e%W5��g-�ڃ��l�U�l��&lI�EU���ҽa[ю��%'�;�%����H��D\mI�09�p�_�RRÙ�Pm����R������mg�ftε-x�6E�t^oTu��V	���BgV�p[ͦ]\�U5��F���ܳ!H8�蕘��{���U^�G�����䷺6�sZ>�����v%"�]a����Q����n��^d���Y|������K�#,����v�\p�(]9Y�gQ�)��9]'V���^b5�cުZ0P3b��WL���ž�훍䖺�)^wX}՘i���Sc^0/�\4b<5�֬V�9�Co1%��fŕ�o��v�9����z,�W:�w��~���է�%_bU�J�:������^ǅ��'�M��8(��)�Qu:�rᴣ".&��X[=��6�%�3�1c�c,�b�U,`�zޚ�C�TN<B�E�[���W����h7,j��g�|�W�wXXT��v�/��X�o-��cpt�B� �W�X�p�ᬧ��r�)^#�{���=���f�`ћ��v�L�
��[��[\���e�8w��5v���l���zV�j���@���7�[�����N��
"A��w�nb3�M9E��Ӿu�ٷBQ5rv��\6��QUUR`�f�����%�.b�C�=O��E�F���1�w[�t��4n*Gd��vY�-^���%�[�ڥ�]�cA� �9�h�u��s#]`��B�vK�b#��T[rմʊ�:�K�&�ܳ��T�pڂ�����N�I,�rKA�9�����,2Bm9�vUі��yyZκ���j{y��j�=�a�ˣ���;;iۭ�,MӰh��OE��J�]�vˬZ�!��MY��X����p��7	�j�YYX��k'q��g�v�����U��^��	龪�UoNM�8�"&�6��{h5tPN��T,`[+��i.����%i�6!ࣥE£�L�u�e0䤜��Ó��z+ɷ����U����M�`��V�+��Ea(p�#=�⫩��w��{6�h=��ܬ�4�u�\���E��kaˣ��8����3�6�F�}-mJ±<��.U�����FEЦ��hF/�����p4��ɽ�N�]ջ�CZ��m��5�ĕgm��am;�:�'�	ɠ�0z��,�KPd�}v�e��8X޺��N#5�2����bYyM0f��D�{N��Th�C�Tw�6�#Yr��tk5˩����Q��zm���zU��gldE��S��6F��p��mOƔΚ��ԫ!旻QёN��-:.fU�S]���F
�����q�l��=}',&��=�Z���G���ˮ5�eU�����Hw4�F�B���l`�E�Z�A��Rz��S�R�u5���[(�!9��n�Qm�nR|��0�х��Օ��g�Yf��Sي�Z�b5tq�QYF�J�:�zN}v���a[��5�|Ԏ�.����Ӕ���9��lv���c��dN�øyJ���t¶r�X�e���|ge�|�W{V3]Y�J�H�ڼ�ۖ�YaD�B�j�b��cŴ�z�j��ZbV]K���,�S��J*:j�M��^b��P�����h��37M����`L�n��U��̥u���U�7�R�[@�fQ]��z�����T�ۤ��,�4��ĥ�񉧒�wbוR��y��ۋ�ѽ�(G
�c�%�wb�����Q�U�wB�i����*�EN�t��lc#Y�F銗SR���q�j	���{�s�	���	����J�]�h�EͦkA�A�ep�/`tx�T����뤉����ئҾ͑U�:Kzx����#��/p��:�iGV����*���;��goV�\f�ƹ��ܺ��h�o��EN��x���a�*��M�u�mI��fd���nZ��u�Z��B�v�;�ph���eJ�*��{Ƨn$��A�ݣ7`x+���R��CUʆ���a`���\����#T���U�����R��Y*�f�t{��&�aŗ	s30��{x�+:v������q�$;7���Ԧo<ĉ����zpΙY�ƍj6k	o�l��O�(R��XK��=������^��Yj��6���ir*����k��o �[H����K]�݄'aZ�z���C��9V��7��z^{����e�j^ծ����H�7Dd��F,��j-E��EW��f��3/�o4�V_;�I�
�����9�}���嗙�U]�Z��U�-�,hz�����ia��rVҤ��*���kFx�.�A�w�jݞ(�Y�����S��n�����L�W}��	Sʤ��fD7oP/�srB�&۲7&w'j���-
J�Κ٧+��,���+lO���'a�X֕z���z����P�}���$���f�3�m@��o6j�KĐ�]ĩ�����x2ї��f�O���WW�|wq��Wb�{�A���S�B{�{�{7P�2܅Jh��Vص�2I�WJ_:ڽ���N�/D\����q�%FT��B��r�Z��K�r�vM��i��L�t��U�Y�\�z��o�*����η�Uo4����T!Y)��kmUv�f��9u�^��Xkծ�S�7��՜�1�a�[}Ed��������h�_W�6D/��m6i���b<o�ڈ����{cj]��u�#�HVrOx��׳7��K�ҹU�Ý�+U�{���r�rk����ۭ�*yT��OD�Z3Y���=�o8-�jW��0���^^1Kq�b\mʲ�=������n*���C"��U��i��K�9�[�N�vԬ���\����mV�
�[�6:r�%�	���������&�4Oح�����z%
��1��*ܮ��������6�a�V38������z�j;n�#^�E�r��觮�,�&o&�X��73i�*�����RI�ʚ&�[R��᥍�e����-#���B>+��_o�B�j�v�'pc��4�ܷ�idǡ��r��W�P��S�gr���ӗ�q)˸���uwW��n�X:J�6�ޤPv֬�̋�����p+�H"�_���e%�]Z�b��E��>�To3%@ft~�2�Y�1\u�(��"��F/Bʛmɷ]3�_�aM��1���/�ԪYmҕa�׍��z�m��\nkݳ6Դ�#͸�pK{�[�qV�gQ{a\�V�鏶�r�,:':S~��T�'7�׻�P���|��h;{v�V]����
��cL��c��7]�3	�+2�ܑgc���;1�Ϭd#�����ꂻF��D1n���蹎̩�T��m�+���Z2�c��<�*���5Y������؀b~�p���n��5�\��q�9]
��Ժ�X�=��nt�:|ɸ�)w�Zzu���[�0�g:�_��L�6�t���f*�ݐ��;G��]> �";+.�@�Rn���Xڧ\:�2(��Vl�eGD��^e�B��j����J���".��/�zb!�6Jl�q�l:À��܌�R�J+a�f�e@-L��f���K�URܼ�a�ۻɺ�#e�Wٶ�w��(���a�XG{����|�6���Ⱥ��d��݈��2�=�pt�KV�=U����M��De��x۶!o��CT��W�,*ɴ`I*t�40\ܬ�٩%͕`=�����m�Ȼ��E*f�a�Z�-�v�!�VVa��k��2^�q������́K)J(je�=�G5�s34L�p2�Y��V�3� �j����g/�)�7&6�e����7�_el���ԃ��vڃ�A)fp���sw���\)�V���u%^r�y}��`��uV^#�X�싷�ؔ[�Њ[��Ld��}V1%��+Rw��%U�idF�F�sH�T(#��ƹ����P��.��Ơ��W`�و���U����x٩�I\��)��B�:�/H�"��T(I��ۥ���ѫ3*2m�S�\��T�h��cL��
0M7�����`�DV�s��Uڧ6d9�Րd�[�QN�I��E�.�mZv)ꁼ��:eJ�Oy�[�z/����u]tS��� {D��8n���$d��T9�8�UѬn���㺣��[J�e�D6PHN���+c#];U
��pD�G7�jT�4�X���%���*�L=�M�x�ދ/�v�8����;,��)���&su�^�f2�:�ƛxs+�mmL˷��jdZ{hEq7��yʥ�� �˞�����Y&�C�y낥K��e`��W9qf��J����/>�FԳ�\�Ūm��^����[������l��vpj�(���&��l-�3)����WN��mm7���D�s�ނ��%zE�7[��\f�m��Ubj{�ه"��]{N-�NZ�=q���S�c�"�T�T�Qu�<}�E��R�u����Qט2�8���\ѾuX-�0g!���^
\#����-���f�+͈�52c���Zӛ[���Ee����y�T�󪣾ra��N���1�L㋉lk��c�['�cy>X雇7��tJ�(��7��2�K��5+�՛^zp������tܰmhvU�����Ⱦ{�M��D�.�Y��1j�H��+MH�t���^��2�M��e�6��VyI�4��L���Ss�F͘S�r��Y[�C��i��s.U��a%�����AԚ:�1�s��c]���͢�b���[v)X�MZ�.v�����ld���^T#6��4
Yw3�tZk
ɀފ[;����멛Z�<h�-�����ڽR����R�ѺA,{QWy�\�ۺr:��v�^�7p�xw���k+c �l�8�L#��aeaŌS��su�oF�a�J�L�'N�[����[��J�	h�OZ�V��.ј�!��T��ӫnJg�/a����Nf볆_&��d��s�p��qG,��;�WVf�ܱdv�y��ԣ�0�KR���Q�O!OA0kwP�"�b��q"�OVi�vQ왷:�_>����Z���0��f5�x�U�}u�\3�w��2�aM17$�{�\:T�aJ�R���$�x�ڛ�p�˂���s���]�˸#%�͌j�;
,Szb�-GS.�
n��cx]�sb�t���:u�9�!�i�BY̷l��(:��/M-�[0�W7X��o�s'Y��)t����޾�;N�ovJ�̾���ק-#�a����ݫsRS�rH�!��&��iC���D��B:7z��G)���
"��t.�Q\ߜ� :
��b[o-u��������k��[�r%���@�.�Mj �]�79C�Pd��7�{*�Iy���Ըd�ʸ��C�C">I��XF�`f��#�#	�xa��c� �؝;@9�4��q+)��	9C�t�����dN{H��NF�����0$�|� q����-3R�@=Ro5_���{^��7I��,�g��\��R�)y�������k�f���Ad.�qڤ���zO��-�&� ��� Ņ��v�W��E���ׄq {��yr���_��l�.,� ��WQ�<�,�q��x7}�u�5����'&���G���.W���vT���������"�>���}����Գ�D��?��>����o������������|n!S
;6^�Y9Qëp�ý�+�:H�j<)خ�s�u�C%2d��T�MT�v�p5\���a�)"��m��6'q��O+��#%��J\/��z��U��i�U���d�⻺��ೖj�X����]%F�xv�rɮ+.�G2JC\M\�*��a�B��[r��}��*�m�ʵ0�R.	�A%�2��c^f�U�w�"����|�-^$f.an��(^�rSuѰtC��O+t�}{���0�f2gn/r<���F�C4�d=*i7��1�Z6.=V±L�{bʾ�K��lb�1���d��Kr֐uc�{/&�`�����wF���0ʅܤ�|��%י��n�1���q��<g����Z���ߠ�Ԏ��z�ū�,�n���Sz���"+XGjŕ2�)�l�O�z��-��ָ�i�r��r�D�2�漩���2�
C/*�M���R*�����\k�^.t�fiKQx!QZ�`{wU��qK��U�#�ui�]9Z�u��[Nٌ7���ر�Kk_��}�t�A���A_Wʔ�q@;���{JQ�#��5)�k.�	��7li�gtNuY�L��#��j�9����#�F���dXkJW7��Y��Y8m��f�^>~��W����8ێ8�q�}pq�q�q�qێ4��q�q�|q�m�qӎ8�>��:q�q��q�q������O�8�>��8�8��q�8�8�N<pq�v㏮8�q�q�q��i�q�v�q�q�x��8�8�As&��y���.�sJ�ORՙaC�dͼ�[RM"�V�7R-�eC���Yx���u��q_7Ao>��P��+{��n�F��vz��來�qVR�w�3�Уj���e��E\�X�+;j��Ev��;A�,^c�i��k��:5N��ՏP��yԯ+EޮZ6�^v�׹�)��v�KQ�v�n櫔��N�2�pf�X8���,�����k�H\��ÀǨ͗v���,�Wc�6'���2�w^���Z�WrZ{�.^��&zh�n�&K�WjWX��d�%�k�C�8pٽ�3��U�qW��[�������r.�6O_�x�Al�	�v�+�SФⶭ	���W��mX�S1��Q�+FD�ڨȼ��FP�t�ق�?�1�3j�yUj�1�7kE�B4�jf%�:��Fvg.Ɩ��Y`�Xvo2Tc�/+9�J�"b�Y����F�9�����v�����uj5(osk�����ݙ��^�����!��p�N��S�vʮ}c�A�j4�7ckq�:5��imY:V�h��e�I;��h���Fc�M���S��ۢo��n�{�s.�kSf˒5-�]��ʫ9ܘ-r50vYc�<�T�#�WD�nu��މp��]䕋B�~-��wBa�Mݻ��٪�M;t8㏮�8�i�q�q�q�q�q���q�q�88�8�;qƜq�q��q��q�q��q�q�|q��������q��q�m�q��q�q�q���8�8�q�q�\q�m��q��q�q�q�q��i�>?����f�3�m	q8�Pa����E����gg����YH9�<���dX��xcDT�;���&�z��ٓ@���l+E�n�Cz�Or���;�ؚ(8f�6���z��Z7�*-�کqeۭ\V�	u���o7��մkys��H�n��b� ���"��kg�2�UYSwa��t�w�^�mp��\;��,{��qȶT�1��9q9ե�ӄ��EWGu�J��X�+a��ܬ9$՝w!y��.Ɋ5�l�췆�N�`x�J�A��ɭ"�]���Е��T%RUWo,�������plU��N�\g1{F麷Op���h�{�ɫ�\�3�:qeiR'�ʴvK)W���י)64e�:�#�53v���W�A�ƒA,{W�r������)73�+���R���e�ϭZ�1��%�3�	��i�U�B�b:6�/s:�n��3������*h�;�@ŜbB�*�����(��n<
�S
�:�S�u[��mgC}/��4.e�v��ءRUMYf��4ch⺕*�WxSUZ�s��^��������*^�H�˧ ����`�ï����F��t�)6��6�c�
b@�U
��nq�����R�F��/N��w�+y[UD�]%��X�@@��Pˣ�1K��s���T�y��I���c�o8�<pq�q�\q�N8�6�8��8�q�}q�8�8�<pq�q�v�8�8�8��8�8㏯������8��q�q�\q�N8�8��8��qӎ8�>�8�8�;qƜq�q���N8�8��8ێ8㞞�w����8gUnmI҅�ʆ5K*�3J�1��v
oj��h�Û�Հ�ҍ����bM��sֽU]5�xm�������1��t�Xk=*��^�n\�u��ˎ� �"��k���0`OѶf�0��]�1����u��oX�8�Y�n��o
�O/{)u�ɔ��cI�D�&)��0�������5�+���3/8تX����u�:-�p7�[,1x�[
��ljʡW�9����-�
�X���(�tn��z��+/�uD!vf�ꪎ�0���)��N�V��[�߽�s^@�TB�ƶ�ø�%(&���&d��UJ�	��q����{��R�{N�!;q�lvn��dVX{i��ݱ|o��qؽ�_\
�8��ٵb���73�eZM�K-Z�%�z}�I���!��jͪK�m�5:tX)�1�i�����v]U��d�n�(-}[%�ަæ��|0�u��d��r�����*��`�ؓ����+�»��Hj(�%sD����K���M�����-jW����2k�$�zOf�SN�-��/K9y+ M�V�R2"Qtڍ�\1%O6�RYe9��ԉX%.0��swBK8�D�V\[�Q�u�Td���{1�e9��-���rF�z��f*��*J�ͺM^��fhܡ�|���m�ӎ�8㏮8�q��t�1�q�}q�8�8��8�n8㎜q�q���8�8���q�q�q�q����>�����<pq�q�q�q�q�8�q�q�q��i�q�v��8�8�8�8�<q�8�8��9z�����k���$m:ȸJM�'!��YX�v���X^]�a<Q��;��x�F���#¨�M�Sr'%lhvh��/zu���5ί�Z������{za\�<���L*����YR�|�NRY[�t�vo�r�^����ŗ:s�,n��^��EʆqĨ���Z� �m$]��QͽC�j,ȫ�E�h!VF��p��iЬ
66{�*�h��p�Z�>�ZlH�?x̥:m�랼�
���2X�J�}�ɦѻ�H՜s��%�(�X���,A.�E�*����i��S�+s�NqT�p��
���-:nu�C3e�������׏�u��94��� R����{V���y4Լ���v:����Ə:i�!���4(�ڡӋ��o-PJ����K�,�2�7J�����H1N��X}s+�����`�y#�64��Y�Z|�`�^i|R]���A<�1KѻM�H�=C� ��'��sU�H�i�yP��w�kd9�V�h׭��4��)��l������ R��ͨ3·heCV��U��Z�ñyJ��j��κS,6!%��9`�؈�T�`���u�b�Y����'+���Ӄr���F)���b�,�)u!"���j�I�XB���a�hfPS�{ne��VKx�Ah^��,�J�q�P�w)U`Ő�[�S<=�K;w2-$f����Ρ�I¯���x�4���I1[�n��9�Pc���[�m�R�d�2�n�� @>�^�b��*�R5H��{vT-ʺ���P�}ʥ:��	�j�6b��7}/��O���T��Kg���aƃ�{؂�j�$Ҹ۱���\��Yb�9Q�g�e���:5R�K˳��g2�la!�*�1.(m[�h.�^�z�Uw1���-�+��,X�7���L��X��Tn�풧-d�/a�/2��ɜfCD@V��A��̋��[�4%U�O:�����  �z%��B�Yk��T�ńØe��*���wwqI\(�əU�g�(m#���D�n<���4��-��՚�n;�HV;��!i�����y��٥$Ṫ���.].<���DGM�J*~�>��>H�`a��DB�:�R
]"u���bo.W�]��#�!q�b��,�9P~9��b� f	�^J���z(J�V���t�ZY�؍T*����o��F��c�$R��Ni�@��j������r�mVi9�oq�A��N��$�4����n��&�s�}���әᩴ;f�Fؽ�8`����^��	Mw��Ѓ�s2sk����5��އ�E�fvw+ĝվ�ϫVl=iR;p�ڇ��j��}b�.��j̩�ި��Yk��U����M�z+)��,�b+��w*��]�kN�	��h�&�tM�z���MS��a��C<@��T��h��)���rU�#j4܍J�Y{�ق��U���,W4[�~"��pRKG�fГJ�U���U�9�'n�n���s���b[ ����թ2�P&(FT1�܍	1�MӖsC7x�A]�-Zs^�H�ǃV_R����i@�SN<��<oɒ���r#�c�񗓉�;�-uw�8n�3.$PHŹ)oU��2�g�.���X���v�Vν����5y9!���m����v,�GN��x
���+����u�)�P�H�ܞ0��щ$�C��V�MN����
H�T�W��^�����qAT�xi�U���A�Vj����ޖ�.n��L�[ɝ���E78�͒��A�dM�al�Pտ"jf��ۑ�8�ۂ�M�Y�Tl7J+���ej��e�"2Voi�R[8�W��iʯ�.f�g^Ε�Z�h���Ϫ�֭܈�rQc�M"�|�k0,J^�'����z+��*WcJWe�WM�Z����a���(vv{9hAb��!'1��u^[DH�w���
Ys�yv���/7vj�('hC�§z�Y�)FH��I�8ޭ�
����nޓ���7��/A����ٌ�����\*��Q&^6%ܮ2Ve�u��S���,w���o�ʲ�f�<o���FT���`l<��$=Z+�8J T��#�E����ﮔ��*bcY�ђ�m���oC���8*A�%-�d",���n���.���@@�WwQ5��d�C���8��nڪcruf�b�L[r�'SZY�z�sh;<慎.���W�9�FJ����Ž�#*��zOIR�է�]ثkv񍱂˧R���ö���{�eL!�(gT�2)vW*�+=i���ɯ�L&�i��7�s�?m,PUK1������h�K7N#��]U�<��)��f����4 ��5�^�x�B�B�����:��I��k��Vm�/D��Er�S3�^s�ՠ���YM��z����e-yԋ{E�q���;ܰ��[���e;��6������:ײ�o<eM�F8�rlr�Y�XP�P�
�vQ��?op�%0��qλ(h[g.q6��i)ѹH7���n��P�v5�-o�[�4\���{f��*+�qj�9Y2+��s/$�L����+��l4t�0Zp3H��!��,�S1VCW����-��*@�s"�j�܅d���f��뷕{3���=]�$�i�T��uXLE�]�I�l-GI�T�8��Y�d*�Z�!9lL��Ճ��8��H1N�`���AG�n������J��-���ZNoR�6�ސ�
V���T��/]��n-���9�ȋ�������COA��*����e�Ruؐ^�,��fg`�dx�2vT��6G)t ��޷�`��w��X�-���%���Eϕ�;U&n/��b�QE>���p�g^����(e��汎:�o2�p,R�Hѱ�,�q����osgnHuϝ�`�M���g[��UN�pA0U����T4�[k;Y밳��j]�sc��[{����z�c̻�4���8�8E��Dv��b�.�Iwy�"7wh�����t�uI�mLk�Uj�o�������ܽLV\{�z=�D<s�9a��Z�+S8�|��3_K��2a�f��m��zi%��,%S�����!U��D���v�U˔(�奔�Noe�G��.:ۓ�j�aw�Fz��#9WƂ쓞�;��[�%+Y@��v_eoK�t{��4��M�c�$-�.�gvf�
��Y[[�0/"�6�c���b��U�bt�"R��M��;J"�2�{��m���wgi'��Qݕ�l���n��b�9�(��ͪ�����Эx����JUX�-QN�-/:^C��
H�2�M^�J8��ռ�:�]�V��-�hnܺ6���شEz�Z1����-�cF�]7G5�L'S��ɺ���w	�s�h3��Q��ۏv�=�Zcl�-H�
͔6��]
Չͼ��qdZ�e�s�Q;��������{U+��N�%Q[x�H۽�EI�B�KJ����	վ�{v��nVke
Rq<n�[�59�1,��fdd�n�;6�h�}�8ˑ��W�����1Q��w��m�ιPT���m��X������rȾ���n�Z۶�+�5N	��(�8b�8�(�+r�����d�.�֨%9%Zy8Τ i��\�P�̵֯�f��'�]�<�s�*��S�ɜhnB��湙
�
�+U����Yu�O�u�3pQ�K�Ο(����ћ]zj��Flrw��V���8�v��S�d{/��k�Q:
(��Ge���LSJj�$vkPe'�^��x�ѥ�Y��m���8]��;���{i0yw>��,�i�EZ�;���9�K۸��57o.[�{t
S5X�a7�a�j���eǊV�ޜ�lf�e��ư�؎l��
rKC6��̣<���%m_ge*-NK�=h\Vc��6�t8
h�lE��F���@�a�)�B�;ǩD5��t�K�R�4޻�����W�=+ Ωٸx�5w*��{t�Xp)�uz�/_����Q C��������������������Q��TFA(G�@ā
�I������a�BI$'�Ŷ�s��E�DP)���%�����tb��h�	#AA-4�^%2����	�4#d'����l�U�'^+ėU@�A?PT���F�B��&H"�½�B�x��uL���0F����I��шܑ4A%
B����V�2�*���2@�f2L((ˎ"5(�ّ��j����0�(Fy��!F�@�҂���?@�*OD��7�y}>{�3��2d����a��<R+N#yl�B����F	��D
�7L��$�����iҪ�Y��E]X��]�Z�*N^�-ݻ�	�������br��Βc���2�ٕ҄�^�6�}[�r��t�9f�mEl�.V�)���^��3�p��!�]��c{��e�Kh>�͛���9N٧}oZ�<�QIw��{�ʸqhJ�����۷T�!�}��~6�45�J�J[O(n,��p�R��P�*cf�����I˹�+mu�]��s�V�p��S�V���)nJw.�̶Ǎ6�Ye���!1ǵL�F�á����U!ef���ի*L6�&,[wu,CuT9Lm�,R�"���HW�B�4.*q�ۘȄ���A��7G�α��Qk
"z�D�{��M�b��;h��M�%Iv��C&��V�d�:�9���mV`�VÁh>r<��������8����U�+r�2�8��7zm�Pr���K*��{�e�ҳ�Z9=����Էn�[�����9쩗�c;�hv�'Q
UZ1�[Z���I
����Ut�K�+�����`��Y.j����ԃ7;i��L����iԂ�`U؆g��.N���E��U����(a�@�M�mCE�b�EA+�0]��F�D�N�%�|� �14��D	�#[A�Qj�m�d�8De!"I#$0�
dp�?T(�	�M �A�h���l�Ȟ��H�ӑ�ʪd
Ya2^i
,(�M4Y�e�H9
���q�<dd/����@�d���q%�4RdOH#!��-�
-Bl�8�-9J4�&$J����2�i�[�H�rˉ��d*0ъ�iHd*B!�e DA��e$I/2Z��ˎ&�E�	��qO0�b2҈$����$(�T�M4Y��	�#�&�M�#Q�a�ňO�,����$,�̄���QQ�$�9
f�,���DFR$��D��9�(�"m�m�,&LMBH�D��8M0W�b&��2���D�E�4	*�mCE�P��Ȟ,���!�KG���f$��@abAP�O&CI�A��@��a;��=� �kwId�!��R0��-ˎ��yE�)(-2�aIJ�	Ӧ�q��nݻv���<1!$�!2THBh��ؽ�#�ͦ�DJٲ���/x�Ru�j��i�N8㏮;v�۷o�q0�Cs[��מ9�Z�=;�s���>.ȹ*��8������8��ݻv����9$�TJ������#kZݎ*N�IS����z�/��,9N<��i�o^�z�nݻv��Ǯu��V��5�ml�箼ֆ��D����2Z�ge�YY�u%��!w�|��	_7�y�z��Ӯ�����;���S;�����niQduq_5�ۥ�󼎻���ݽ�kY�۪��֭�u s6؋�ȴ�ew[O[E��b�7|ov�w���r��匵mh���P)1;��ݷ-�gm���*d��p�Yŋ���ۙ��̵�����e�1e��Ս�enݝ�%�ߧ������z:���ndk[����Y۶�e�����ߵ}-��wy[n�N-���vV\]��)�b�ugd��Im`����Y%�E$Dٴ���@�I�f�\���/��y�	F�q�\%H�&Jh�a-
���rE*/!-"��X���\��D�s�fhS���*�<�E�)]��ֶaK]�����,^N�8i����/����kq芉恄�T�[>2܌D��$��")���a�
��@��,�L�R�,�I
���E�B��V�'��)�."��M��>]�= �l���X�ҕ��*��JUPp�"��4�d���H�TY�H)���E���Ao/�;Ǡ$�Aә5/��կ&�Me�Ic2�K��|&n�f��Xx_wc�íV�{;X�X��x�N�:�Rۥ՗��`Q5!��Uq�����S�'�6�̗��7<9k�<;H�
/9��J���v�|����_*��$!�L�A3�:��,���*C۞4%Tu�Չ��U�.�*.��:�'�m�&�v�����.���q�!������JIb:Jӱm��y�6y�]R�F|~W��&�X�*s�=��Q�Q4���́�\��X�Tă���8U�٫`��N� D���3�3�3�I*�y�k�۪P�T�"��������t̵��)=�	@ܥN7������N�G*��|�uN�f�[��]<��"	����)[y�������^�O{2ܰ���̻����Y��G���"�Ft��nM��Aޕ�k�2�%d�T�ι-�ÔSML�9d�Gݛ/t�ل��w;�q�Ų�o��˶M��d˔���0��6��#����J}�^	�WHV���K��*P3_+�22��bzC��HŃ��Я�X�|v	�M�sa��U_I -�G2�=y]�a�3Bd5�<��O�GM��6J����Wne�Gm��]\� ^_V�Bx��%5��Y;1�/�T��Mqgyv"�����a鎪�}����v����來��p��8S�w5}L�:0���!who4rY��_lS5=�,��zɦ�t歙���Y��N~/�!(ݑ�W[�ѢV��N��\�u��\5;�n�r͵��yC����&U��j!��4ٴ���QG�hj�[��>�7�rx��(�����͝hLr�沩�h2w��TQW��9�)�>Q򶭍�:N_MӎSu�Lbe�4-|�e���ۼ���/bI��
��9y2�<&�Z�M�̘7�y�Jf`�/�S�J튑�a%��ٶ�{�Z�l�N�W&���,�#�6��:p�m.�ȏ���"�e5��D�z�9�{�k�
_\���C��g	#|���Ӽk�p�����<�5�OU�t�]+��h�U�~R��r" *����,�M�ȋs�%_L�)Q�=w����9���:�{9��R�u&��(�Ȏ18�^���<��r����ԆowI�%�|�0�sy6��O|��M���ӈ9^��&�]�� {o���V*.i^���s���8Gs��U��؃_�5�!����k�N�VWa6��A�'����}o؜oץ7����A��B���KuO18|Tk��to�g���6F<eK!��'E,��+�զh�V��NW%��&R:����x�+�w�H�>�52b����n���|�}g6�NB[��*[��Cf}�HRT��*jz�ݱo�#�V��n�Y����o�%:̣��F�C��+з(%]"';4�(O>bʃ�{5��m�h�{���'y�DS��տQ��ۤvB�h�i��qY�ۚ��CE��I����0����q�m̪�&_��%"�{��s���ßQ���N'ئ`�v��{gN�MCM��;�kX���W2jj��s�z+@�$���-�^�nh��k{,׷}��*X<9JD���F��F*�b#VV���C��|�������:��g6¼����uF�_X�#��>���1Qb��s��'.�n׵��$��p��F=9w<�=�2�NS�Gx�xq��0�����O�+v�60lu���Y�_h��u�Hn Ѯ}e	ш��?6�9ϷQ�F؉=7xj�$؍r\z���[�y)a���9��r�Ω��X�o:_^��ܷ�;�]ۭ��&݁o�j�{�v�霝(r�ċ��ߺ�3ܞ}UW�8�1\�-����������ԝྃ]����@�#M} �Q�H��M�3N��|P6��rՉI��nu������z�[����L���J�_N��Bzb|z��-��>W݈�SA:�	��ç��]�v5�\�r�ԞV�Tn�sջ��f`������s���Sw�R�w�v�2[Q��3�J��/2Ru%�:z�hU�ԕ�s)m�Cn�#��e�.�xq-N�k5V����77�V��C��vVatv_3-%LO�
Oj�wF)�J�IE<�6�Ρy�*�gN�eL�� ��=���?	҂��g�E�=:�6�}:�i5A��׼G1�Vp���P$��&a鎣5ہ�J�`��fO�������N:���ñ�~������$.�)�g��5N�<��}z��	aU�}��gl���>��1hg�w	� ôxB����z�]�����2@����42׻�
뽫�Aڕ5WF�(�j̨��vxr�\�f�Wp�F��/��޾δm��*�x]�u\��<&xsp>A���|�'W���X���=j��X�s'�ܣ�{~ت�㔊���ݯxJ�q���,ND_SR�%���P�1�f*&d:[�ӯ��8�3'�}!e}=�C�9v�.�:eaT�ꢊ�Yi'\���{�&��E`:6gGf�v˂��#�A�Z�`7^W���'�4R��hU���I�d7��wg������0r�JSz��T��xYG�w�¦�J��U���4mBeܳF����Z��P��B`�%T��#�-f`�g��:��]n����`|*;���r.��(���Ϗĭ�>�)�]L�q>rb��MĮ�"7�� �/���4�'7���,g6;����X�<�In�Q�}���3�t�����ו]V���sw[ʛ6`��n&�z�_v[�]"���x&���-f<y=��o����Z�vK��9Ga�|3U#���L�L����V�zy/�B��u�o�N�yɻ�µJ����;�=��8����ě��T�3;�8�C����4O�ؿ���5�er�����1<,қ�d�$��)ֆLZΫ�y�yn�it������+�B���ˍȾ�ᴣ�B�C��/+���s��wu��_+2�5�T��Vt�fs3��ˢ��A%͋�S�S#����8�2�r�#��0Vb&�Vh�	Jg&����̐�r1���ki8(�7j-�W�r暒���s��!���N�qPD��j�*5�\w��]�37@�Ȫ+.�)܆�MJg%��6-�Le�mMP�j�U'��mՊ�}�nї٫8L��SV�i;Q����2}��2�������J��w�z{e>]e��(v���\=��;x/��9{ ���|�_,��OP$m�H{���sFjqk̺)��\��[���as )�����a���}SK�O,�C�"8t�f�^�C�㮪��:�}�b�+����۷�#�5��c���;z��+�Jx�)��3��(i�Hmd�=�t�y˶G�V��ww�l��jv����ӽ�﷠�����8s�&�:60����K{c��M�E�s���V�o����n�����~_o`s�~�ޚ͕3j�r74�g ����5��=5F}5 ̉ё#�}L-����%Cr*���ϔ\��ꪨL�WΓ�G�5P��ÖPV!R��,5�Y�K"�R-vp.��F�c���`� 18[�����f���5[So��nk�}A��ɩ��+��î'su-�H�&�����ʫ�w��O���f�p�Md�-�ش�͛�-�M8N.�Z�I�*yX�8m}�:�Y����#9.�(�Ʀ���Kz� ���ܼ�Z����3kpZ�q�e=�s{;,1'�q��&�R,vU;���}�ivً\�k-Vb��8-1�f�o�S��y���ʍ�]i][RQA�|�MDEvv�dJ�V��AK�*����a\�Z������GA��M�������q8�>�����ʻ�isny؟'r��|Ӷ�w�@�{�첆�5���Xk=7�s�k8�^�N�|Î������97��{)D�3�b�����gs�=è-0T���M�Z+���C^	�ę1ƫ�ur��P�~��㹊{���&I=C'��c��7T���)}�
�k�]���*�:P������5�B�ύDpn=c��'FHQ�W�B���f����Nv��a�Xw8˯��6�p����+�U�����n���1�{��s�J��RU�EVLN��gA�r��)�\/�كlM�2��;�W�+b�v=8KC.G�GP�|I�Yx�"�b\*��T��ueOf�V�;�C�+5��7r��&��1:\�)���KҘ�޹�2� ��(5�ٜGj�J�7�zcn]u��^�ˣ��#��nMT�U"�lB-�^D�/�v���Ü��|��#���1��9�*6��Y�C�Yڱ8c���-���b|�'y|ho� t��8w�4���D88X��6����D�@���ۣu�);M_��_3�:�v�vU´�y�����K� ���V�rP��'[a5����1ӂNd�zOn�~ Ϡԃ�p4��#d�X�� oS�>W�W��#��Ϋ�j'�W=�f1o�n�JEr��+���#5�lw�k���n��qb;��0�=����C��CT��W��	��`���Գ1�Z2������ո{��������
�h�
�5N}�Eܻ@7�vFm�K� ��+���Q54�#���k��P��5�i�|�8����C��c6��=bG��[��]�=��U�׼:�����;.K���,��=jbظz��D��)�4�inr�)��e��S�'Wfo�P�q��#mÓ��)�7Bw+Ү�G2'z��k(�����*Q���P�k ���b�,Y��v����rH�UUU�.�R��}��I��{���O�T�ģ<ƃ�@�b]��}���*{�vl3Y|���Z��9�HE�tq�F$,��+:���c�c�'p�]-5�n���W���\z�i��j���������Ƅ���<ŕ�*��4���r�<$�q�}�u��
m��	&�bǍp�����5��729З�y��k��Z�M��>n��
�g�3rjҴ�L��!I���\C���"߹Vd��K6��+Ϟ����^�S�w˧rYඝ0�T]���J�q��~w�AW�V��������m+����)o9�FkZ�������ІN�N���� ��Qwz�v]§̎�ቢ���g+�b(�p#�̑	u�L��ki�3��_y��8��T�X���+~$R�?`x�g��#�xx��	Ȏ���{}S�K&���C>����a��,�#wZ����8-͘&b�4��՜&����w^F��z�s�U�2�R���5$�&�+1�}�z.�{*j0�椹aA��NP��*5��5�R����u�ÞuoV��]��l�p�N����n�c�̪�&�Ú7��o�����Xmb�fLr�EӼ��X��'w;���;�U��V-�vav��z�3��TN9!��!d��s-��te��l�#-8��7�R�k��s�;3ر]Nv��pv��;�UW(�ug��H�^�7E&!=�S{it�4�m�!.�X͋�:�c�:T3n#.�ٷ״�fX�R[�H���r
���K��UI%�_$�l��	٥K�r���,!:��#+J��*uS݌ƕ<�1J�ۢ��^�{�g;��Q�*��ڛ�����vЪ���nCZ[�4�m���(c�H�%�b�L��S�6�:��R���a�������t�܁�-Q�m�*�AƏ&��r��sf.�꺷&�����uΠ�5�z�� �B���ް־h�pU�p��VmcFtO�̮�S%�Oi�vQ�ÆYq����
@�
��y������y�7�.mB�׊�u?�VѦ�
42���v\����l���L,+w��zs��CT󝭱ַ]�9�݋�u�V�sD��sx#V��e+%�Xw��RձK��oQKv�03lt��b�������8�L���D���#G.�#��C
׭
"Q�تfY��T�Y�9[(���6�^N�a2��	ж��kp�/����Δ��8�kK�޼��_l]�:�3�tt�[�x�ݎ�0v��f���b%�����5��2�c��Tr�����&''U\g������I	�b�b�N����dE�u�2a�T����|��+���ɶL�#ӡ>����v�����X7]�)=J��ʽ6x�����Kc�dɷB�P�$��9��w;m@���Q�Y�*��샰vm՝X&eS�W�˶��A���F�	���zUI�Sݦ'Y��|�����$�Y�8b�"�,�1�͗},c���]�L���JXU��1/��Ɇ�q�3P�6�ʫ�s3cX�e���C�Vr��x#&�¡R2P�Z�6솢Z�#e����iq�A\��l,�V>�}���-�E �Q�>����R��u��t�o�u�X8�1�ͮ/8c�P^EQ�|T��*L��kn�o�CTb#i�c�[��út�G[n܎�nG�u�G�k$̀�PZ3&^��}���4kVnhf�#2i8���ڱ�8��Y��/Zb�hHν���
J���o���fS������7F���/��$}�I\�D�e�q�߸Ԅ	HSM>>�v��nݻq�Ǐ�{��@�I!H��$#HRNEE8uI�������^�z�۷nݻq�ǯ�}�ڄ�:B�: �us�);�q8�
BI$)�=z��;v�۷nݸ���}�����9J�w5�W�i~��㩣�H9#���>�}z���;v�۷n޽pW\q�WDG)�[�:�H��NR�s���.8
 �(�8����9��nӢ�J�+;��(���q�H��X\�@��I}m�'S����X��\�_K����ˢ�;���躎�*(s���$A �	 �x|"� ��
�TUow(�7+�r�#	a�0*h�X��v9'Vk�2���F./8�X�"�	j��z�t��� ��|||`{+�h${�����ߞ��xd�.<릘C~n�� ����-���i���D��;�h��R/��o��pa����{������a�����M̀|DF�G���&�,��]��/&�[��+.�����҈G�҈���3?qi��c��>��=�ұ~�7�TdD>���wв��Ԑ4��g6��P
����} 3>b;����K��n�U�"��H����o��/}�'\����o+���/���w��ߐ���@h�V�ʭP��\���\�α���js���0f� �Emi�'nH�L�Dhok
މd��SL�*4)�I�����৷p"A�i��q���LN=3��U���������Q��!Ds�_DIxL�8�=�+�Z��lz}n+�2P�Ќ�����gf�����o!�}��a�7H����}7���z~���1��Z�msxsW�E�Ȼ���R=�[Ӊ{�M�_k��;4K�{�{WE�x??�c�������+D@���Y�={��35:~[�R�kH����o�zcVq"�Ҽ=��h�%���G �8}:@��`9�?d*�j�#���>�}T}�w�p�+�����]U�����6�$l����0�9�Nl7*pܶe̸
���#�Wk��U��L�SNH��H�D_h7T�j�&�t�N�''Rp�J��Ȩ����VѼ�c-�:�U�,d�s��'�Us)�^{Z��s��>1�c�y�k7�^��^ "�a����|��g^�c�l���B�#���H!���#�g2&:BL�����y��� p&�C�5o(}¾~��h
!Z �8 0�T詇 t7]S�������>�4[wԧº���@7F������3�[iM"�gwY?!�llB�}��������c��� 7�`9���C�w�B]��i�`���q��=�L8���2������v�vy�-S
.�J:� }N�ܯ�f��c�f���[��n��O��4]q!����l�Gy����M{z`Ǎ�[nA~�w�P�7���^ }����}�����|�������AvO����f�ؤ^��Sb�BB��7~���m�>nE݃@��|7ja��5�����V�N�����·g��Ķ= �M{\{���ޫ��1����1�:���C������y���ٶ��ΞG )'c���/ߔ�<>�doܕ���Z�W˥�/x|� `����O�ڜ�������4WV�׌u��@eE��lgA@��[�
,?z�0�cj�({�E���ߏ�Y���;��ԟ?,�[���9w��1���X��*�>�r�kv\���I��|*(�@֨<&�P*�*��E�Q%�É\�[x�5Xټ�h��Rw5!�! VvvQ���J����?��D �KB�b�m��A,oR5.f�+���j��Z����S(���8�q7F�yH��f�K�򉗹��e�[!�1��;�*�v��$���x������0'\��^Sc#jŗl���ۯ�����������9�~ \_�,�`�)�8@�t�Ͻ���Q�^
��N-�?Q�Z����A�^ e>0�zh/�5�C�m�g�¥�e7�E�͕I�{D7���*vN���m�н\B v��tb4)�+�
w�xa!{v`y�N�x5_�Tc��Z�g�oD_Ej�o�Tn�� z��wLm�n�7'\���,F��5{��H �8~�hp����4���7F���qmOSE��:C�z�Y��fv�J*��<��f�҂Ƶ|��&�qf�_]�ì0t�gk�ƕ���ŀmwH҇���0^�^����|;p��|U� s�R���Mm���� A�-)�ЂQ��x����������%�DdH��L��R,�������\�¸��r�����a+nu�03�[j���r8Gy =����`� y������������M7�P�z@�{�B�'υԒm�j�3k\�^3U����[H/A���E��<(Ak�<>c�8r��=�"�P	�_Iat&V��ӕ*��uM!�_5�������/��<�Ou�uA���F���Y������ת�db���{����-�7B䭜�->ظw^޼�{F�r�L�l:��]�ܸ:,m��!텒�mE�F�l�����&`���W��,v����ʰ���������}�X&�/����[���&}��}/F�xek�{��꒘���|�s>jT�{��f{f.��W���z�?�F��H:ĳ�� Q� ��t�>A�8h��
Ll�k������� �e��Rzj����I���r��J��B���Nq@6aL<� E��Ů�s��7���+�vg��^.�\0�!�+¥:_C��*������A�:�� q��[�l5;<��Z�-�Y���\�l?.�g�Dx[X�Mp�� ��U�<��%5��!0
��P����ʌ�O����� �N�>Ǿ.�	Đ((e�B{`,�1 ��5�Q��D�<ԙ4y���O1�6������۱����PW�������R�����m)�}�	<y��e��L���31㐽�s����hz������C�%����	c�M�A�+�S����Z�ă���kaL�c��6���O}�cCy��n�ɵ=~�y�:a���]7��Q�j|�5��r=�G^�7��<�Q��{�)��?HP��`	U}I�H�2C�����PcZ���W��`*1[㎇����0�i� ���b`鹤��;:ubc��5�fǑqv�0�j5�1IP�},�ܘ�ml��L�q���NF$���7ʭl=F�9.����:ő��ebޙV)5I"3Z��ʦ�5�ts��7�'�)ׇ�bU<Ҵ�b�XW�6�u�	S�1�o/a�S�F�6D�;�9C��y���n`�D��0.�����{�7k!ۚv�ݝ��r�Rw���}��� �
�c�T
ڐ	�;�8�����
lV&D��Gus
�R�ᐓ!��XC-ڴ:۩�f���:��m62����5�
9�?̑=;�n?O�TN��=HCϷ�ը��wz��@�O��kޏA��Pi
�� ��y>�����O�ǀ����:��1�"&�9^�}w�L|7�i �g�$���ހ1���5�'�mz�{#��c��=��77��~�Tk.۷KZC��w�#�Y]p�@w�t�Ӏ���CP��^�"<�MC ��q�؊��Bx*�;e��e�9퀼=�l�"����B.c��*��s�К��J򸊯��^= t8R��1��7n��$�Ο-_~�����{T�3T;��/����Ӗ�7��X	`-% ��dދ�!��	G�n<�X��|T��`�s�/a�c�^
!�L@tP�>��������~�R�TUa���l�s��3��1,�,i��YE�'�Y]H���g�Y��~p1��W�BY"��x��79�ҁe!�c]^��[����\G&�	��pN(i�d�% K"�Ъ	k0j:���{}�����-z�V}K�A�bU��C�\یO�ĺfk�h_G�^C���k�u��{n�R������j;#j]z��p땏?,!�KD\�ss�n��u����6��X�*qlQN��"�F��26�]�����)�^�N�u��\�������ҵ#MSL�F4��A�O?����2���X;K��z@L&�
t�������0-�f"�n��&����;"��ʭ���/����A���7��i����@O�9��H�]�'�ԩs�tż���Q���s��gZY�f���Ө��@y��3��A�<�6 �>/PK��=���?��3��9�P��-?#b�b۶)^��j�@9���4�@��xOtw�=���Zjx9�]I���4�����Rv)�>n�����������xctLw= �x?��jV@D~�6�� #_�}R	�����Y1�tL����on|����o	gO��#Ъdel[�Ư8z!�ֿ�-�h�H@��γ�G �(�����d���I��:W��zqZ�v|��v>��ڶߟ���Gf����p�{Q!%O�V};$p`��� �SP��f�p+��ύ��d��Rq��,D��}� ���z���;6K[�rk�:'�>;�J�p�eM
r����	�J�Cc���^7�K�0��*� �r�9����o6�:��c���"��t�_g�xD�q�`�������p�z��c�9Sr�)���i|�V���(ӹ�"�n�D����x�y?t�U.����ri���7�.��x�-�Ț�&��Elgf�[\ҙ�|ot�߈fձ��(��@�rl<�ʈ�_��M��Ǹ^�e��j��q��Y�r�~�9'�Ԫ�=�#����*$�hB�iZ� ���=�;��^GyE`�ӥ{CN�E���M��&�P�1�=8��T����*���9�c��H�|ko&��6�v1������y��*<���f�A�X��D��Γ�q���/x�-�n`Y / ��7�L��1�9iwq�S��n���Oeԯ�cP����mL\^+�-��$��v�	�Y� �]\�\��g�b��lx3I����q�o\:�%�2��	y����)q �_���~������"82��� &+�\���)���E���P���3�-P8½��u�l��!�� (S�u鄞�Å�&Ɯ�Ls��N��*�[l��;��0gWW�;���g�)ƻ���@�[AQ|oG�=��p�} g���i@�{>/+���`�d��Mv�b�Do ��HkȦ�jxЯ>�s�^w�xa9���|k�M��>1��b��������ވ��:����S"�9���.h�d
�;����F� 8ܶZ���U�3�(G0yn^ΐ����S{��ܢ�9`	�i��%8�#rݘ
m
�ݕ��JNU��g����z#�[�З�~�3��/�����|���k���Ҡ4���ΐ8ľ����|l;�ߏ
Z�N�xEATݘ���Čܫ8h�Z�Z�yU�n�vy���w�WQDo:�wT5�n!�au�:��"�k:ܗ}B���p��vR�AE��ڨ귋%#����vPy��NV����L�V^�BO�c ��J4҉M4 �4� T�TI��y\���� �@��>8Y����`��E*�r�
zV����G0��]a*+{��̀��F0kۺ�.�� @�1����b|�;2�<�מ}��`���Bu�+]\^�P�\�pn�Rۛ�V��z<HOA���(��q^2�O�LL��H���/d�,���+wh���@{s�[�{:%={�"j��0����B��`��/����3�@/I���[`U�U}����t������	�Q Mt;�oO��� l���^)��p�h(�._�^O9�Mى� <C<8^��=P�"�����}�E��}
~�͏�{&|�pi� ���Hh\b� {�	�߽�i��~�x@�%bg�vz�j��m��(19s��<h��n�6�̫ӊ���{���{�*=���3:-��X0�}#���l���o�68Jk�3��=`�fW���g'��c˩q���{C�]�p^sEy祙	 ����X����!�R�e�g�霻��؟�P9� �fD���	��J�o�V�g������FCϨ8u���'wA�y�$�I�^���u�Mҗp��m,N���Z����ѧ�A\�j�s).y5�G0a�tR컫'0�u�d���J��=$l#	�*'+�yT`o����Йtw�4�Fm4�����9:�H�^`Z�dьC��%��an���������@)M4��MTD4�X��Y�VAIdAd	FE ����0�$�9�6H���gцgS��,Sޣ���I�>�s�{���� ��zu���ޑz��=m,1�:r1H龔�8��'�&��E��W�u�:�X1����7:�g���XY�J�Ѥ�����2���09�}}"M��	�pge����T5�K�4��e�����p�6P�,��@�|Di�#�>�S�(w��V3]F���1Fus:�ƶ͜=�5�N�" 4D�wCnb��~�50��=#�#�����i����Y��'�������3r��I�@{��ˠv9=��  @U22�Ű�������;k��vl�~��'��Fjf�v]�����nP�e�/��q���z�r�Q�9�@�$k%y��_�[w�g$�Y�g"aˬ��%�I@z�کץ�_$\m�Oܶ�?C���oW�Bg����x�DK�˟�����ϭni���X[	8��!�9���*0��@��dIc2{��>$uwr��<W���4�M��R�*�����a��zC"Y�w�h\sL9d�m��O�
��C6�E�7 �����e�/�c�nd�z��g#�U+a@��M�v�ڧ������\ӇBO�ڙ�O��j)	��D��E�����q�YS
c}'TS�sp�5�T4��Yv�k#mZ�SZ^�-bT'Cr���Xo2���'n�uK����"��a/���M!Q	$VAX�HB5ڳ���n�ue�]]G
,�2(�"2,�$�(�qu�]�wGQDwu�~�n�(J�����zq޵��F<�ňM-$(������Ǘ��{h��T6�=]��y�;���5$B�f�C�6%��VW�:
I��]���<��A��®a�>��B�����F[6G�����Sq��@�~���	�o����ϡ�mY��Xp����������4F�Ư
��b�o�^mߡ�w��`WO�ށ�����q��<�?��+�B���_N�1>�&e��pt��w�Y�<�<D��~q�Lk
�������Ľ�b$�*��4���mȧ;�ԥ�]к$�=�����ϕ�c�D����k"�y�H\\[RO�!1V9�Q�!7l�-��7�_���D�z��_�綩c�~�d>�G�������zlbk* 5.=S˛�be�,�Y��9���s�N�B��y�ʮn�觟��(֑G8�xe�Bz%�fGG"v��������^9�%\w<H�!7w�,�w8X�0�;�Ƕv@�`�	�M�u0��!L8\ԯd�i���cY�/�O�Sc��գ��qK:x�])怪delX�$%�+��M*�7>{��_=�ʣ֦��MԊ�cB��mgm�s���pj�f3B�tELS�-҅\"l��:g�J�+����ۚ���l;K��z�u�/^ WS�	��ܰhq�s`�ka��z�uL����.qCR�Ѝ�n�έ{]���Z�(��R�`4�/X�T���[����Ԏ�Nm����wv
�I�A�nGb���G�W�����uwWf�#������x:C���v���Z�����'A���ś���ut;�m������b��P�{��̮X��b#�co,[��9D uY�s�;��f�]gh�ƕ@����^��kZ�a��b�V���Z�������IG*��F�n����N<n��Ɖ�W8v�j�g(K��*�ӭq��M�nո�-X�޷0��/�jE/�Z�2UR[��ros��'�
��O�l�YV��S�I`<d����l��$��Y]��e�ɠ�n5��Py9!K��vcC\&ݡu.ꃫW4�zв��R-�v�*GU����י�q�I�bVQ0���:���oX���l�|���Z�h��i��,��fe��؎��FU��h٩/{:f��ᓐ��]��3Z���8Mw�6a�{���\EMgcF;]u�"j�;7aܻto��_*����<�-�+4i�(\��9�T�h�rlь�~���7z���f�B�Rpm_Qf&9uH/Vc�Ew�-�"!ԉq�E�N��7�a��͑�ݼB�C��<	Q�u�y����=��l��8UQB��@��HB�QJ�q�%&F�L�����b�ë�[�2\p[Q<Ӱ���;!ޱѷ=�,V���Bd1@�]�uQ���ł���}<�Uƅ'�h���1���Cgj7��¶���]�rβ�ڏ�����+�98�i{m����pʢ�Z5�*;FUe�vUw1�`�䥒��lߘ���\*'M2�VE���$����ky�5^��m;��z�]���^N����Tl��7͖vҚ��G'���U��˙-�[k$���/�K_9����ܽ���&�I�8�ial���n�kN�@��&�#eK�r��++�[��d �n.3S������8�
�׷1���$7�]�Of�kk>�{5N�F�ު�z�]�p&o�����G5���$�7��,5)	�p�zZ����P���Rؽ�i�썐J˴N5͵W1��8�v^kDTZ��B�;-��dCۆ���;pϱ%['z�QT��$ڻ�2��
B��F�2^�>��f�WKI�EdL�S8Uf5@��R���F���Y��SC�W�m*�o�6�,��N�J"���J����J^
�udk��l��Vk�ͼ��T����@�r�<a]���
w��'c�OZ��.�v^���殢����x5�ٍFQ�{n�Un�N�W�/f���t�}'_��w�~U>���DwE��W�j8#���"����:���㷯^�x�۷n��}���rwG�q$9�$\�pq}�/�:"�����qǯ^���Ǐ�v��Ȑ$"��]e��]~�����@���Ɲ8�8��Ǐ<x��~����9"�O�W�RAT*!ʨ��RXƛq��v��Ǐ<x��,�� ��!}+.���:�#�+���.�#���.}�GE㝥GrDA���GD��I�q\�q�qE9��JΉ�lqrT��t\q�t��k�Q~5�:r((�Z��I�s�QQ�A'��ϓ����n���`����-���"F\n�,��R8I��%Q�I��g�<��DW�\7��g�ǫ�L��͕ƽ�'�hL���ZE�W����'��ئ�����D�aQC2�"B�"C��T!�G<�M�.6�RBi8����!��H�� �\(�H)� `�[�����Te9	E�d�fT�D1�I��)���@%FA#�* H�ƚV��F�� F�U
E�� �H� ���"�ɧ3}�<�ϙ�w_�^	���;��"l̠�(�2��U[���O�d��;S�z��O�(Y�k�zy�s�rz==�3� ף]�;B��b	�xg�(A��,<�BhtɨC�az��'���$^�'lzi�"�A�*�z�8�k�3j�ѻz�?G8>�;&B�� ��!�-0��.$rCcś��^q5��4�P����[B���?x70FX��uȘ�A�b]iR���zkNq���3�=$C0��Z��=oۮ:���e����[G���ړ�6f��$u�
�'kc�8��r���I�$?v�ky{��2�S���&��IQ��>�M���-�<�����v�i3Q�c�
��C�z`��ME6��I�ݰ�zYX׊��r�N3�1P�X���*��4��'OA��0��a
�q0��6[�@ȍm���X�X�RRq�\�~x���k%�n|[�=q���,����~�������?�S��G�p�M�~Ȅ������0�����΃�wO����`8�D^\�;�d/�-~�JO�B�R* ֜:�d4��������������ᬥ��,�d*p��>4����w9�X�5A54��Dkz�'Z��P���Y]�iNKj"�E�u�8Tz��ǔ���5G�[ϔJKra��ؽ6�aF��i�^�*R[�W������K�$��D��Ѐ�M(�4ЀTVEcM�EYBE�����Ҋ/������x�s/H����
�\��v��Fd�vI�&�2�!��"!KSt�e��!rڀ���CZ���8�2.�Þi��m��s�~{���| ��j�����3���Z*dB���[O�Ǒ*��,*�<7Y�["�9c���/'�q����GS�J�r�!Y���!~kmB�ܞ��ԙ"�x�y���+���j�M�V�Mm�0u�!^ڗj��bטT�>�R=���s��#YW�)u����O�c�AǶ���&� iyY��yժ!j䶵;��8?���i�;2��`��)���q�%�D��i�{���\]y�5P�V�-%�3�!����dD��<�o���>�	���tl�p�<��n]&��)��a۵�q�l, D���_"�������E�i�Ro�(������5_9$|�e܎��oH�hwmI��%�ȕu�<�VD�9@��sV�\����V�o�'.z$�Y�?T7��s�j�	z*�!A^i�a:�@�E�O)�����@��ۢ������ynIY��UG�2����ґ�6�c-:�Ot���ni�#:#V������]�Q�6�DɁ��U�[7Յ��v�RWQIZY�d�7Jv�/֟�`~Yx�1�{�M�38��ܞ��k������v%٪�"���EH�4�4�)�#M�X�@�QT����$A	RD$DY(���9�p�����}��x��, Ps��+�bX?mH��.R-�rcG2�(VD	h���[��t�2'��6��ʔ��XqM����A>2U��� �x
w�p�OB�7��c��M
s��81�l�F
�F��n�	z-
����~������/t�����R��@�3���Փ)�jRU�F�����3:zkw�Hql��iyŅm�y�F��̼ފ�HAu��7��͙����sI�X	U�V��aN��wn�W����������q�B#sL>��t|�K�r�/e���g���.���������At�R5':{i�f�\z=Q�u���M�/dI��N�E񞇩%����t�w������� ��r�,���N���k�h�?��scO���q���3Úo��w�Q��p+睶i�9X{��vO;�e��y^	=,�>�-N�6�<#Xt�G�2��xl[2%��g�f������|�^V��nt��E����yN0mL��+b�l�������N�FS{-�B����Z�0�&蚄�P,+ݕ�;}���*
�u����ðQO�����	�9��4V���N��fWT/^�D�\&N��F�!L-�nP8�2��f���U�5�m�V�<��*Q��y`�8�U֦o3����>�S��hB����F���"�hF��F�E*"�
$"H�H��<�y���i�5�Z���6��S��m0�%�-�Li����5�W�s`����Tٙv�=�	�m��1��}s
NȈ�o��������� m�.+��LZ��vS	W}���O�Y��E����$E��k�*�	8��ؗ�]^��/��Cn��c�I5w�x�p�ڳm>��8�c���7Mmp�>����ߗ{��+9�竣Bhf�0��MI�gUN���{hX�3'愼wʀ�-3��aqg���!��9ԏN���]�v��aQ߭���s^ݴ�d�
� ��	��-���6^��1�m!����?x��f����Ѧf�WK9��+fl�:|�I�����oD���u��|�7^�;3�[T�K�.U�nӮl*g�Z�Hky��H�M�~�� ��1,��%4�������c�O�U!����S�|s��Q�?b_��?G�=�rB>!���
�X��Y�%�LD�V
>�l�
4��D�n�r��}M}�B����<�i
��;peb�Ӭ�p���)9wM�o���J�FK�*�#5�1���-�����Y���ȵP�G��Uc�u��6��T�X��mQBSi��ɪ�u|�G��u�O��/u�a[�$�ڭ&��k�g^��<�����.�ڴ�:�L\i� ͵;�ڪV���&��9��\�@��4�4�H�4�
SM(5AB��IQ�d@�D$ ��9��ϙxc�fvp�B5��JiB��b�䊋����Q`Z�1e�>G�V��R
=Ȅ�@Lpm���K���V��+��㪧�cy���vE�n�%���_��:ٮ�|<�J�9L��]J�\mF�Ov�n��F;^�	�=%�3�/����B� l���v|n=�%�{�'%�v�0���zdJ|�0%�cv�]��)�,���b��TG�^�z��3^��9=I��mި/�6��0��N���΄*0�>��^٭#���vג��%����!���O|�ߚ+;�׭6��)�1{0#�H��,T��N:a�k�r2oe'a�M0�-���c�����9�J�[�~mj�Y��_\�5����&&~q��E1��7��v������F+ě�Mp�Y�Z�ŗ�v}��{��V��%���o������s8o�!D��~�\��u�34�?{�6D��y80���Fa�>��(���
�H�;���L��`�{�x��JC����-X�j�Sq�]鶐r��l�ɬZ�!�0E��.qL��sӻ.��=U:3�����$��ظ���Bׁ�8�T������\"�)��R\Q���ا=*oKi]j�N#7*%�_3wJ>�����/���,O���{�h)T��bл��2ƠM��[�I��j�s��8B�ԟo�\m�����wL�K���޷��9�{� "	 ���F�hP���j"H$�F�P
����"�{^�dB��a�|4=�v(C�=0��	\Sw:�(�=P�zd/52�\k=o���{��(�x�c��d�l4��܀O�w6���J�p��pӋ2y��oc:
A'*�1
:wou�;��&O�G�y4�Nڂ�����0��T2^S�y�S�|l�D&�|�������Qף�Y~�����)��d�*���5�ug�9���4L|
�8tJ�&ߎ���J�9��~��z`s%|�(�x��X~� ;5��܁�硙C�~ʕ7�sDl�aF��j<��qr)m;H�)��M|b�X<؏����W"A�iQN�y&���)���kDs�K3CD��^
iOA�<�V�OU�&�5�t�xk5�%�F���'�z�#�8u�E��5{i�ˠ����聭��/)�	3��/�3��f V�a؜%�MN?�V�okʾ��ϕ�/;
�?\(�8E��D��(T)�k*0%�'���ҵ�����W���7�a`�]�Y�>�H���k���
4�I��Y����T�=|�`�� ���B�F'%M����wF�x2��!��/Lۚ�1f��N�1e�#�,�+fޚH�6>U2�X�Y�Gu�5|�(޺�f��]g��\��Iԏ^cz��2uof���ۡo)�w:մMDl��5�7lجvS�/���Mk�x�4EFEX�@�Q@�4(#M+PQY A����7���缕o� ��:���}��)�OXv"$!�7Y����ҫ|�a�ĸ�#�3F��]��{���g��Iza۵�q�t<1��l��lz&B�FW]L�R���l���}�����¸d/	R��萪��ʀ��|����و�jt�<��J�w,��j4e�/�`�`n�B��ry¨NA�2��=_tIw��諐�My�*ތnjr�76�>���j��ʠ�#�yw�+�)~ҧ�#��25b8���r�œ* 8���hfb�ݕ��l�	^����z�\S<!��6�#�S�-�-a^A��w�#xL��O�M�f�����b�)�e���,\3J$���?�_��E��U3W���+�+��h� �,����Jua)LR��]z6@�|׶t���bC�g���؃'�����d��{Sc͘&��3fQs��%�{�ģ)�>�s�ܪ��{^�Yntj<W\4|$7��*"!0-" ~�zB��.�wИd*�]`����3Vv����uWJ�^:�?:ݗ�MWb��r;6�C�Q�GXV]�7�$��f0�a��zAY����>J�Wk<��;�uT���@'��5>��n�놪�uN�{r�@��S[6���v��t�ij�:K��Ŷ�r�m��*�{]�ܭ?�<�"�"��iZ�)h��F�QZi����� xx0a�o�Ԓ�*:�c�|�����Ht>���g��{�)�=25��S��K�;~��*�|�~����`�m;�,!�����M�0���z�H�Lar�p�ӛAM|�\��ٗXlrrpJ
&!qɏ�p/���ܿ/�I?n0���s�g�~��3���gf�3ͨ�ӨL�!m�2�j0����ߩ@�S#+c1���P#�G� @�1���Pp�N%�t�i�������WJ8��A�ڮ�{��ލ=u#�'�ǟ��s�R�]�+�wg��BG�~��}T�p	�:EwC��6(=��}A�W }�*�������7Mt�Q8?C��I����[�	�>���,�����A$ȓ�рw	V��\Ì�e��[D�m҆B�N�Wz`ީ��@�����^>�e�^�����W]BR��m,�П2S���|�@c����/?zb�;�*�̥
v�B�x�ͧ9�G>r;a���,��7)�X�Nf��t�Jq�j�Gh>lR}�f>���'�B,�?tR��uB�Jr%���su�f��ADh�ĝ���ɠ����'W�F��P��s5<b����A�Y6bi\)VD*���b�<n�A�#s#���k)�������Ԍ��Ȇ*�4�򐻪�nKĖ�«hn]��=�xu��l5�Y#{=a:���M��T���~�E
i�F�	hP�(F�j#"H�"�Ȫ���D܂�X��f�s���恓L��2i��F&���v]ئ��;�2�o� �h\��BS]�2�&�Q^],w�XwŎ�w	�q=	�1���fF��⒆=hW�x��
��	K_*_[nw�\ixd�y%4�£B�(�|f���fo��hc�1&|���
G�zF+����o6��:��o'%�q4,f���hj��|U�k��w])md �皽ʍK϶�eh�yX�R�ϯ)@eS���T���$����m욎�Z(�N���-��~�J��Ù���}{aH(�"m	��m��$��s�ɨ��Y���z2v�;.���z��Y?,e#�||���W ��	u��24P�(���+�����$�-ne�	ؖ����Uj@\�Vd&0���2�q��1흄yd��C+�k�\.��K��F�(���['ѻ\���I�,�uq{˴�>5C�q�'"!+����x�g�iDDr�<��@b\!�:OR��"̊U�<�i�5��=���S+0t �S���3{��y�rء���8g�,Za�|�����#f�Rq��a;/F跾��S0��?� ���K����1��[2� V=d疤
��z�wzP\�bWS(�ٵ��u5rL�	h���i�����P��ɴJ�Be����(�ö��LC'9v��m<S�����~�3	�����w\\h�9����{�}���F4�-EcL( H�B+QB@ >   
K��3��~��?��Կ���P�'��E���M����	����+`@�sֻn1���k��{����}打�8Ej��+���q�3Ô��8����َ�����y�y;>� c��T&�e'��x ��c����Zz�x5���)tʊiS���7	��@c��M�;{_\����⽹<^Ĥ�kYFCH��e@��p�^b�y"�z�n�k�s���@�aֻ����G�A�)�:>Q����%c�Ī�g�4͝�Qx������x�5M_��,|9�����F��{�e�
��`<��<�{\{�2;�12�<�%p�MIn�k���/�E�VWT\<���ƒ�����S�.���+��Z�Z��b��<�C�[�
>�35�x�L̗�&�H܋hU�oG�=�'I���t4^�Aͽ�_�Ch�/��|��?1�x��y^�\h6�����Я�[�}k�E=���Y�~�2����9��Y1��S"�z����|d�5y\j���ڨ!�N{2����F�T��j���gɭ�s;��K$))��J�Y���j�:=W��M���k&�qr�"��܅.�ռ�q
���9��H�7I2^�,R$\B&N�ӂdjl+{�z���,���ʭ&���[UE^�q=qRa���������)iCSaoq��8��a�ɰ���X�B���,ʴ���y�T�Y�]����`L�R��T<�F3��uH�Xu�[�]n r��E�ʭ�Ĳt���N��Z=O�Z0�����A���rRp�O`"�i��}[���p�aUJ.k�&���И�*�Y�T����tࡴMӉ�:���U*o*��(&��O��::���p�+p=��K�*�oVD��Y1����dq�P��D5�E­q]���;�հ회*Pj�*��Ц�Wd7���σ�XM�K�L�S_8d���}����˺�	��}zSe܁��ʅ�͉C�����۝��ܭK4oqU�U��ds��+*s���6-�E�S��f2��U�݈I���a{�/)�:׶k�x�e<��t�}��Z�s�l�n��ڍ�9�h��	N����+i��q{
��xf-;;ZF���v�%i��h-�G%z5^��Yk����V��U���p�*�P8�{�`�VVf���������9v�S���i+kr�X�P������^:��E���.�"f�Ȇ���IRXda���5^+�����%�����N���r&C�V迡A+pe2E���v�=ItK7Fz���Ib)}d٥�+�U|�n������@�4t���k�+vhs�]�2�mʭ1&0`�R���K�o�E����GW{�.Z�-���Z�n��ѷJs�ؖNF]���ַ��ڌ���A�9��ȷx]M��׶�)2�$����cW5�5�}K�`�Z�,��ݨ�FܕKڴP��3��me��T�i�Q�r�夺1W|2�0i�_I��s�xm,�/zF���;SТǏy(�����Mݓ�����׋5�QPҷ����Cp���dγ����RK��ʡ��(�F,9�lR�13���aٵ)�Y�VJ�2،6A�t���环����ZѾڒ����R�N6[�{;Q�0?D������#��]b�^c��4��D�K��8Y���4��ՅU���S��)�W���UPO �q��"r[���J�ū'meJU����ZV�l�(�aK+3"H�C ��L5�o&�ґ�sf�z��.�k���;/����\�v͌��5�u�r�:X�טCF�el7O�T�:f����7����*J+xoKU�B-S9��O�P�6w4,)$D��x�*p��3��#���B �%Mjք�r�������b�M�v݈��{�:"%�y����|>$|��ֵ�wQ-���Ê(�1�o8��n<x��Ǐ����u�~�e��W�e<Ԕu�!!�Z���4��8��׏<x����$�	BFBA�&��H#�,�R@�e4�8��o^<x��Ǐ^���@�5EBH�%��tu��u�4�4�8�ǎ޼x��Ǐ\1�$R��ϽvPG	W�g!!ϝk��#����8��N���/Ʒ�S��qG\u��Gt��uQqĜqݶ㈦�}kTt{Zμ�Έ룺��Q�y��q���w�$x�H�H�'��FɣI��oT���û�f�[]w�d���Np�t�Z+6a��\۸��.��0�%3My\��h{�ɳ5���,��i�$i��e"���*(�"��x3x3\�mԣ�X�p�032���)����'z���P#��0���]���.��8�]�bv���'q�d���ÅJ]�eͳ9��7��u�nL���E���c9�Nq�3���Q���m��?Z�~^Pr����}b"C¡�'M��5���?O�nU7pyW�t�to5�j˯�Om`*�a?��4�g�����$~q����=UR̰SK�h�&�rWq�s¼��2��l�k����C�A���|�����_;8cBk�&��u9�8��ן\y��I;�A���w�"���B���!���9�*{�Cs��l�����o3��2��5�f�(0v�BK��Y���$@NQ�r7wӱ�8�چ���}܇������p�T���Ү4`�_	g�D8��T'����y9�5y�r������s �q7��0��ͤ�]����)~�x��N�$O�O���r[�4^>�zEW�W)�8�I��y|�~ޢ���wlw�}|�N|U�0C�ئx@�����~|Ol�H��S롏9HJ�.�K�_EE�LMd*��K�Y�D8�J��z�L�p�׆UX���#x���_)���;�ku����i�m��M�	oF.70o%^�y�9��s]��X��M
fY��B���	�G�{d5ӵ,��\e;5���A�Cv[�n3�o�k��q?f��"ƚ� ��* F�
����=�	����Y?t�r�����;���	�,T)=���a�z����p��׀�zϡ0�؊�ؙg똪5��u<���P���[�24Jm��#��`�AR1R�2���^��ə[�m�x�ŋ��`�U���C����s��$Y�G�fQs��b���ƁF�
7.��nʻi�UY��F$�Z�t9��M�3�@���A�
o��C���=��U(��ybeںfr��u����nJz���S�mv`�/���*�p����Ǡ��}|�?4��S8���d��籟;S
��1尙P\�]��'�4����-�64��Qb��}�N���v���U�o���#o�]�F�F��J�s�q;/N���,:=í~)�����t�{�Gmڲ CZ���+yJװT7�����G�g���ded�p�>(a�>���g�7��%�8ж�C�>�óe���O��a�Ϣ�ޯU�ޝ5���[:ϐ��̪%b�;PfB�@|�a	>~mO�0�T���0N+�(t�P[�O> �k��m=R�����<"WO�"	�YwNU�S�Q��9���OT΅D�3xl+1BC�N):Qq�n){�Fu��o~A=�{N�dIi����ț����y{r*�=��Zs���SV�V��*o���3rEn\^�8��+`��0����� }�D��B��@��@�X�AQ@�A$@/�<�|���V�7��b�pb�V�)ÜJ.�2L��N�\xs%$ok+���}�m�$����4X��c��|PO�z,?�d����ջ�`��M,A������!��/��IӁG�ɕީ�sF'�$C@B�d��z���d��s��C�Xsէ��/i�hȵ=���U#�M>��q&�(��O�X�/��PU�[4'�n١�/]��3�j�C�k�G�j�]��$��&�Q�C6m����OH��D�q���V6�:_�Y3%�p�nA�`��O�
Q�׶f��u��	Mw�Pb֞������͚��)C���N��~�L�e3#kDKw���쐨b�iAqCLK$���ej����{�FB��czg7h�֯{ε񜼁o��$xN.�U�E��&�1�D&%�tD�O�60�,���=1�S����(]�0��V~��>�^ۗީ����" [H��n���^�;��i��A���t�{��s�"���KzYtAd��EW0�LYz|�O�b-� ���$Rn"�Nx��]�g��w�h��R�|їi��̥ۋ���HO#qsH�+�V�wH��B����c]�3������r�N��S�^�|8�t�u<����wi_0��V4��sp��:h��W1k�,��z�f��
Y�ȉ�Uce@j��<�C�v㐩/���j�q^щL��sAk\�n�$1�d��Vj��o�a{�0�y^�B~�� �������*$i���������� �s����C�+z��K6ׯU
�}'�7�d&�~	�L��"7ӭ�����>�3&�en���`�b�8�/B�M	�:�0%��^��|�c:RqAgO��>�S#&-oCh�{J��L�6��$s��� AT?y�D�����~P�0�>��_u@\F�ӥ�=�/{+s���c>LXO�}'����2R� ȱ�����*:gX��t���U��<s-}��&���k�Ə�ƹ��c�ɫV3͍(�>(�`��	�ֺ��~?�0��![[Ms򕻳O'�n}�2����'N�A�J�B�lƭ�Q ��ܯ?Q�i�<Bn7{�)c��g��ݭ���W�<�=#+6Qz�S���3)��Nt��v+�R���2��l+C|1Z��[jx���7K��#�J���Q�4�G��e���É}|J�����l��jy��zaQpÙк|k��z�X��f��,U=��;�� �\�+����/=E��`���aϐ�������Y�s's�.c�J}vJ&�u\����[�[��2�"[�e<�j�U��n鬔�]H��лsBEV�dI��l`K̸L�6���h����n�Uw<[�l�T�a�9m�$Y�ɛn�K͍iM����n�lJ;�ԙD�D���%4�-4ҥ4ҡS�f�37��-(+S�5��ܽ�=�<������I���8�}=A�T��0�c��ට"�<�&����n��ϼ�"��]tD�W��
q[������Ƌ�Hkl:N;yd�)�V���wf Ҁ�lk`i�#6M89�J��Qzm{�B2V��"n�Y��_׎�]�Ը^�Q�ǔc#|�¤������1���i����8�2.����4�o��?D4;����۶üDk��p�9y�@r�+*oc
��<�CP�r�ޥ1�rk�Gsm�uQ�]��p����}�~kTHs+�.����*�b�S�:�����,)��=捭��n�!k\����,ὅ9 ����Dat|vs�0�>:���j�/�^]�D����謠o2��IװT��G0�-�֡�it��c�^����������C�Μ�f�
��~��-�a�h��۟wH�^�CM�k�Ch:pȺ؋Dkt�/&ۗS�[�<Ek�޳�p�޻6����������_���ᎸȞ�Aͭ�7;[�u4��eF�U7K�eԿ6��b�����k�E��}.E�W�J���Q�i����I�ӵ�\�Ȉ}��뺘GL�S������&�/��m�ڶ.klN�Ѣ��Uvg;�������ٚu�/�����{��8e���n���R?f�)���t�����n�W\TU�uD=V��n�w�*�C��!皘F0�����~TH�����o�;�绶����L�31��Q�#�'�W�P��Lw��'~B7\=��(�W�lzj���E�nBO�0l7<Dg%�ہ�g�r"������YIl\y�kuB��>!��� wr�W��Ϋ��U�
��"AIefJnv�n���X _(u�N�z�ȗ5���2���c���h>DLej�����5۲Шj��]>q��"S^�	��,pm6;��7�����o>��v�[>Ч�U֙���w��\�ֲd��O�4iO5{z%:�%~������N�ˌ�s7�1%~���)���և��uϕ����f}����,Sި�5�&q�N;\��ۚèMu��p�Q��zD@�r�����t7�]���E�S���㋤u)h�V�C��8�&gY�������٘]���"5��m��Cy��Jw�oJQo4:�n��GVn�u�ȾwL�PX���\{ߐ�����=�?�����LOG�Y_}�;,��\�fe�X�,X���]nMd<�����hvqWUDC��]��X��Iۉ2��!�-��Ze��M1��l�&�>�HP�$�c�[�h�y�OQ����Ak�b�̵�1��U�⪷�gb���gT�Bb-R�S�8!ٻX���{��D����a ���04�5�4A�HTG�3{�n���ZC@�ȉ��Z�ٱ�,���Y�e��6�f��¬�y;�W�.�Hч����<��1װ2iAƾT��a~I��#��uN���B9�I���r�1,��$	�"7k�o(X�?sԺ��'��F���}�:��`��iM�m�u=YNo���d���̟Z�;6o4��P�T6�n�O��3���9��K/`@}��nW��Z�P�	Z>a;�A�{�5�~*�?�ALlVO����m$E7e�w[d�6�	�"�3�����B0|W��y��8RDd'��`������X���aet���lth��,̓����-wW��f
�j�E���d&]��a���[��~xi�����/��B�����������	���C����U�R�3)۳�v!8$���)��n�{�C�m�jBcяM-B�����`͂R��	���|ؤ��l�GH�z
7V	�k�\/���#�5�!l�>��q鑑l�\��x�Mw�Pd�j�4^����b���kf�zjK������+����ҏ�PH�$\؉as9�
���q��%�{	)�N8$�dj�3ռ*DlFoM�>�8��]�\��V���P����k���3	t�͚�hoˑ��W[/nE�y�+W�7��pI8vŴ�Px��ԭ|�;g��z���8�2mC����b�w�[�� ����Q�H4�@�M@�O���s>'|]�Ho�
}q�|���"�����HL���	�c�Pq�D&%�6���y��'G\�����-Nhpm�<���e^P����"GdY�°c��j�R&�)��]�gl��5q����F�U��AD&*ۤQ����9������}z��"�؂�C؅^s�R}gw��{FwD+0���ӏWG�P��	���~E<�i����w҈ތ.��wF�C�?�j�^�KF"�G80��Ϟ��^�T*���x�2z	Gs�e��û��zҼ���]ɂN�vv
��"���zdN���-���E��[zӄ�������A�-�y����E�SPv�	N̏|�p�H}�vd�	}l�V�<�_�Ѭ�͕ft�Rז�|Qٜ-9p�U��0����� �!�$�#������vO�����q�i��Vi�^J_^�R3�oi����7���F���`�`�glv`�S�+~��;U�jZuD�j%�Ơ���6<z՚�����;H���}jg��ȗx8������pt�y5~�8Δ2oB�^,�I5�R�3o]��xLͮX�!v/���B�>���* "��I�;E�V��,���	+K���4�a(���aY�3+V�}2QO���(4f�;Uݺ�D�Q)�S�T��-��V��j�A/��  ?�R�4д�@��@$B(Df���X���ͬ���LYp���dy�][�K��G��ƴ��y����"9��9����E��N��P�^j�,#�qm����O-�ϥ;���2M�J2V�ڃ����9��7�e,nC���@9RN�������]۲.F>�k�'��t����p�6�����Ԭ�	-��`�u��B*T��$t6g3�|�%�=�i��F�̕YYא���)�UBg�B�=�)B����-!�����"�1�#����Iו���`{��V�g:��y���Dk.{�[�XUAPS%8���a;�m���m��x�Ω5�j�wk�U.:r*��֠@��V�s�d��I} �^W�~~�/N�o��
:Vi��h㳨/h�->�ÿ��|��4��}t�"�����]�-�&�{�#lC�Ö�r5䯞n�;4�:�	�4t0�C�.z]7Y���t�{��y�Y��]e���s�	c͐�o� ܋��f~�D��q�Q!��/��H?�|�c����x���o�n{��j��h����	O6ӷ{�"�&!\t��{5��d��B�6�$ yEH�={��"��}��f�<z�j"���>���`OMj�XQ�`�Q���$us7�Ӿ�=��Zru���P�$�0�gTL�e(��h�̿y��'���4��
B4Ѓ� _R�.���V��nl�)�)V�Mm�ռ�'�~=�Z�ha�t�TՍ���xK��1�ϓz�r�@k�A/m~U�V��P�~�t_��{��'�S�Q�0�@~�"���bNU�X�ޥT���@�L9�3x�9���W���	�hsH= ��ހ,4C3�����u��;�3�}(�z��m�i0q��K7'�vl�\��PD��O`�v<�
��_h�S?"O�+�d���J�]��a_#������|N�텈��F��fgb�����p��~Y	>4�Ͳ����Pʐ�mg��7���8(�5/|'%H��]}���)�2���F�	Qmi��e]�'�3��b$;��Ckd`>-��~<:;jP����/ߐ�;~��5[�Q�۔�_��l��
<(���?�[�����
��T�dQ��h�!�5'����Q-��§�G>6�j>�BU�L�ʂ�B��U�A��O���'Qf������}�Xv�{#�hL+��%;��3�`�
pӫN�)LPRU
����@ ��{�xʕ���P��:k�`���)Ȉ�	H�Aw��D�os
�wd�2Ûg{�^�5�Y	����f���%w����E����j��[�cq�Q8���Ի�ڣ[\��@�9�V�YCĹ���E���
�m�������
q��Vl��HЁ�����k$�`ʪ�Ɲ3y660���"]N�26·\-���6�ADBsH9C7ط���{[S���UM����nE�#�X"���d���Op��15�rf��w/v�3&B����V˗ei�ۭ̌j���5[X*�s��u۬M��+�	�q���0��\�y>�%�\��ӝ��<��Zl�\�k�� ��Kq�KgU'�jS���sݮ	z���U����i�C���S��L����:XM-��,2�.n[l���6��t�F��H�Gp]�y���#�Mԭh�+'�,8��c�KS}���4x'V��7*��F:M���;��#@֩*��ۢVn��m�&]��N�:e>����P�SJ�)�:�mȔ����^.AnIN�$�l�ح���N��3�-���D�|�'J5��
0�v�'՜��SBz�1^�w��i%H��h�������J̘ڽ�za�0+aUŻ&�z�nT7�N��˻)ee+�v���f"��c�C���N�M�Y��7
���;��T�r���J�������}�q��=W����Z:�[�;�q*��²߰��������.lZ�զ�EA�_[wc��M��P�C���_�]��ep�����CY��έ���{V`��
�Y����<��&3�G	7�#����]9N��Q.������Sb�w���;��SS9�Y]����lL�е�f���M͈&t��� G�h7۳rv"�WZZ��y]��d�z�/&�m�����ﶺ<W7B�{���/�����W��o���̻^
[';�%\�U��tbJ?Ug����Ę��JƬɈ��X������ԑS��ى��q�=�G�D��EG�%�b�Y�al�ht:L�S����5�(':�
'zԁ6�ݸ���c�[������5؜�1�EN�j��?X9��Γ�<���A��b�06�q*V�BB���Ů^:�T�zrs�]L��ٯ���ۦst;��Z�o]��#e@���UM��i��s`]�!����B�9ͻ��C�)�y�$Xc��x�G�"��>.��T�0P�W�V]*�����6��M��b��$�[�/)g<p��lo��ܝtH����/&a�s��w�[fAx�L�z�71�e朵7��W"#x#b�n![�^]&pKr*�ʺ�X×nH_r�����A�el�R�p�
�j7�S��t+RL��ko|��W
��:t��bp���$���$u�q�RA��GIG-��>��x�ǎߧ�<x���o����A�\]Ą�I H�i�iӎ8��x��Ǐ�	�� �TKZn�?��;)(?^����*�FI$�ӏ�;q��o^<x��Ǯ���¥A���5�I�H�I�i�4�8��x��Ǐ���"ݨ����>���yr~%ݕ��gDwVeɜwwwe�f�h6��Λ����9��g�VV��++.mgk�����+�[�3#�f�(�r�l�mӕ����Y.�Dv������
�Σ,�#��:�|�y^W�y��l�80�.=�<lcm�L�2�y1l��A�)9>j$S��}I��*್��q�ENuK�=�Xvo���֪���@�����뾸,�ם��W�j��z7}ֵ��܃YA��H	$�J�(�08	�8�ĜPă�5!q6�L2�5�S$D�+�9L��%(��D�@���h�QZ��.QwV袦��u��H�G�z=� �G��iwڋb~<�ܷ��ΘLc1��l,�	n)�5����s�I�k�Y�m^��'�S򜲄c��_@"�z�fQs���8��pl�ֲJo��؋�#����d��5�# H�Q	��e�7J�
E�{����t��E�+�Q�;>��!��� ��<�O��1�a�_��k�mxw����C���Bc�6�G�T��N5�=��Sda;ӓ���.Ξ��q�O�`%��.�Ʉ1;e�P����P�1J(2g��X�]~��a�n�W�)�4�oq�w�*� ��YG%Y��{l���[����B9��;$l�N]����@���_���/>�����������(�del[�t��k�"*#Uf�aP082W���"<��7�:���XHC��1��������f<"Hq�g7ln�!\����A���gA@r����]�䋀�q��E�s�}�&�"b�ǅ0ɫ�X��X�r���<=�%��($pji1�����`Ћ�*p��.2��LEf0u�����wTH�<�{:1=|  ����o�P�Y��hA�ӡ���t�<���Ai���?)��(��7�cY���V��ߠ3�����E��D�#(�eO�֜;���#Ut� R��'ÞYZJR�7�s�ҁ�}SE��q�ӺS��*�܈d�9.;�6Z�
�;\�E%��ݭ�nJ��1�@�/|����p�ٴ��v�Z��}^Me
~��"���p^��g�rb�g3�}c��
+�$��_��߸�p��b}�1����	zh�>MB� �T���
;A�b�O���9��3Q|���ŎM�AG����8��ߔv�2b�%W^�A�%6_A�U���ӌ.g��1�"���e�NJ[`F5^���3i�<0�py�.��!W�O7;��g�D�N����L��Ţ*�sZ�ҡTu�5s�9y��x	ุt�̄Pgg���1�t�w��[+��M�f�R�n�!���[���R�kk�����`@0-�JD��e^�D\�3ܖKp;�`�,a�:�'ܩRO��������W�<�;�i]����ѐ�^AG��-���Q=�v�T�,!0�d��(W=�v�7��2�8ŧ<�5⁇�f��s�蕮�77l��������s�gn��>3M�3�����Ix�jF������3�^�d�"b_�{;u��1w����3��a���s�0师��&�ȍ���N������f+î�ȃ�v���
��Q)ܘ�̬��[�{K�2\��i��`	E�G#U�����L�r��5*�SU���F!Z�oX��c'e������n��߭h��I�\9�;4;��՗N^�/sUa^nr/fX*?�`G�g�f����w�u�%u�o����0bpl����z���0%gE��,�
�'3z�z_�����4�����=��O�M,6vk � �_�qMa�^��>vz��T�T���Y�����q�����3��o-4:9F��"�"LO��N&��2ߴט��>�S7����9)s�.��ć��C6'�;���[����P�et�"S^n9*�.���[��v�H�?Q��P�
k�V��׏���]u	݂]'6$c�[��sN�����]O'ڮ��Z�W<J>ϣ`L����<�X��L��hW��~X	\��r�c:ˊ�K�c�nHeJ_��^�S�~�
a���ڄXv��W,�t�ۅs>T��oYGAT�7uyj>�oj��:�:�1� �>HlD�v�MM�⺱�<�6�6Lڍ]9������LF��|.��2Z� ���2�Ք(Q���\ø�ﴑ_tL�I���v;����7�.���{sJ�

��liȎe�~� �)O2o8S8�tȯe�3�V}���_A��޹������v�$���l#t��֦�ɘ�H�X��
r��vs��xTm�P�>]Ua���!L4�Eg½J��ĩ����h��q�z��황nЭ�(�D�`�:���;8�V�	���O[fD�.���Q�1wX5�|||�o7����h��u�^�N�c��4���4��<�X�]�
�Ǜ!U�/Q���
U��[>��Uk�F}bD�!F3��s͸�S�ާi�<���E�3�Ӂ5vL=��ه��T^��@�'X�����1^j���`��������){]�'l6�Q���R�$A��[��AGL˨�;���|va�d��g?K�uRdt���:�Qe��-qqKw���k���_,"��3��
# �� a��()�m{}��^��¹�X��4�a�9n�8��е�O���*�j�Rܝj�ѐ�]���i��
P[2��ʃNL6��ҘI�����A�('rT��2�{��@��=r������y��c�|���vƩ�;P��?�0��no�ܞ�bgg�^΁������e��=!�g�U�]�Qsx	/ь��2�ƾ�;�`zw�"��k�.T������Z���2�[�'�׉>#3���״N���S����`��>����R��JqE�se ѩ�W��}m�F�T?AX�t�!��J���z2(1#�>�-�"R�m��!i��� C�fl;3+����RDp�ZqKW�R1�jƗo^:�IUH�v6���B3i�}��7g,ܪ.�y������1�~�|��o&�.���߾��X�����2:���+pv��E0eMs��m���JI�?dY�W�����'���ץ�6�5���y���ǬG0�ǒ��H�|�/��Oә����O��r(���G�e��=>�6���;�Fy�Sxg� ><0��f�U�?v�p�YC���[�y��$;7�\�-r4�L�+�c�����zbt�5?IH���Pq�hJ9��Kۈ��Ϩ4R�`$dw��-��>g���5)*�� ����Y�e.�����3 �|������1P�=Fs]>��`X~j���t��r��㣫�'M��ף+l?!��	yB�IgK]r���W��ɋ�<g�!���]!]Aw�h�e�/�]�w�͵:���3��D��btj���L�ވe��X�B����/}���^o&!��{vq�!h�C����',N�.�Rqw��"QA�T	�(Rg؎h��sB���<'����76rR(������t ���<��I_��~ ���ǻ��[��� 6�B�݃������\ߦ%�*e�Yn�0��^T��r�5O����v�uvd��A��'�,���L�]k{܊Y�����7:���9�L}�f�1d����m��e�ێ��ɝ���J�$>�]����iɕ�gdU��ip�Z����詛��m�i^n�i׺�uw�%��*l�=�����:~1��=��7��K�}�!9����#�=2NG��N8[��q��Gg:-�N;B��e���Y���y�5�����>�G���+�9����Q$��Y�>��f����������8�E]�D�/s/ib�g����:�;F<g�'�a#��yf�S6�=/��3u5=+Kyl�Or�ݕm-,��BNN4 �Px��9���S�דF'�"L���<��bVh���2��2ݗ��2�^�ҿd���_!J����@�!�[0(;���Q&��,�U����Ęhڻ�O�OX�p�	�/�}���OMR�ñzPg����/N��Α��[��C����N�88{�D��EG����3�8\D�{q��H2k[\�1���,����ɮoo�`o�p�ͫs��~�`\؉as�y�,��F㷶 �⢟�9f���9ڒ~/�bY)22��ơ����SۼzA��ˋ�L04T��8�������ם�}�;J�X�4|�#�Aר}�f�y� ���	M��i0����u]�*i������/<�˼!��KIҽ�ST�މRf4��Uvш��9�&Ë������9ڢ�E�Q4>�ş{
���|�Ѣ�����q�څ�r�K��q��n�w�c�	^��"�.��V�})��pak�չ�o~��������39�n)�}�!��a�-OL@q�J�r����r����iWt��#}>��ز*�Ouy3q���[�Q��y�?7T��О+T�������P��-98�G6j���U�홥�˫�V��Xh/��]3C�-�i�m�!��~j��\�b̄�'�}�|���֐Í�K8@cü{���� ^";b��J|VG�M19�K͟���W<N���n�mu��`;�B:�5� ��r����l%�ZC��o(G���ץ��N4�T����芧z�6���L+�H��nt�C�^K�< �<mǲ�Â��>;^�Qd�Y��҈1�0�Vo3�8�V��jJq�Ǧ�Wc��}\g˩|k�a ����l�gO�jE]�+�p�x��mUt���f=6��wI:w�x�`�j$)ؗ����ɧ����T�<�$�8}8jj{�L"�9��@Mj�3���HI@�c��3���� 9V^�F�����^m�<��.�H� H�+X5>6���zf���.+ױ~���B��v�̣/���y�ڑ+J�=v���^{�#���N�^滟n�v��5[��Ehc�ac{}۸ju�+hx�^ ���ǵ�mj��e0�n.i�bٽ�F��R�;�M�e���5<��έ*	��n�J�X��Ĭ���E���������*���gS�0~���y�(�sW��%c�(b��#v����~V�V`w��hH�
�|�OK���}dv�(�P%����x鎷.b��ƽ���
Cb'�A�����]���$�6��·�����]� �Up��\��B���aEv:�����c�}����r�N�m�[=LE������ݲ �P ��N�|�=2S��FM��hȳ��Y�p�M�n�:��Dz9��8�����n|���Wi�3�.��Ȣ�W��假�U�P�땔�~���l~�'���_~[Q����Jޤ`�����1L��2����]V��jչ���v�˶�� �8�g� 5诣A�az]1�}�QWԘTS��ݼ��q�r���.ǝ�nJ{��.5$'x���|��7̛v��M���T���7�+�Q��g"�Q$�t	����S����E�z�N?M�֑���5(P����=�$�$C6��r'"��T�*b�l��R�a̜qǡc�PK�XU�V��`r~6.�B9�[��5sx)�6b��̸d�"�{]Us����G�7��<B�3+���y�e�vk��d�{N�^�J�J<��>Ąhm��y�j3��;���'\/k;)\��V���A��Ob��)�^U}z+3�Ǚdj�`]ǂ�K!�B��>>>>>>��Wm!��NΜk܍�r�L����B%21<�9TA��.9�@t^aٍߨ](�@t�3��Ǧ���Ǆ�49��ڡӃ�5U������l��_��>!��Z댟��W�^�Cd�E�^$�v�u�7������ہ�>AB%�����yw �oV��?9��dP�E�}c/Ԁ!�t[�EwR���9�����$�|����4���^)ẽ���!��}p��Bp��f�p�ԏ���譧����C��ft�5�q��&�f2��� ����qb��.�7������"�}�2�)��H��v�I�����yL�S�S�L(�Ɵʶ�0�%�u�5�
k�����{d����;�7�,�A2��Z֝Q����ȑ8����wsʡަ=�y)�L)Q1_ֱhik�C@F)W�k�w��uE	�oD�V���	�y
֬�ݘuf���{x�wy^�<�D�r�)��$8��]ʗ�C$���Y�Ft��Y��hݥETOfp���a��лb�P(�aJt�p�m��� ��\����x"'�3P�`�`#"
aM�l�b��C�ѭ�*��9�6��݀�J:�G�۲��gv��Vt�fj;.g�M��F���}T[��a&���{���5�J"U���,��+C�3	����M,H��u���Н�a6K���U��Xx.�)0�l�^t=���Y�����"}��������oo'3��7;������
� �Y��N�81�:}L��%��$��?/F5q.>��͏�q�����8ff��]"v���|���ÌZ~kJ�%ߚ�q0���|����~s���<*u�6�|	�.s�����e'��3��+(�[�G�i����v8�0��X�%C��d`$�;�
���3�ɡoL���;L��Xt�
=cc��X"Y>��8�P�쨂b��8g�a���f�V��:��1FͰT�a�ؒG��ꓑ�0Jq@-�yN}Ch�q<�ux�Y;�N������>��1��'*:k���|��iϕ���[����T�#s�}�=׿��n �?,�����5�f�"􈣥k���ψ���|�s����>0o跚��������d�����4�u�'�CO�?R0|�Z���]C��Bx{��I�P���;�����f��=���/N\���rsj��������R!粯��M��rUX�����ǚ��b}��(Z?0·|���/��,����Gc�4����	�[!� i���GkA��_u���C�:����Z#%��^m�D:1qH�f8e�Vp�3W��5��2��V�̼ye�(�m�s�=��a*�N�a��-+LK�_5n�Y
��HY�nz7z���b�w&��#�̳�~�98�
�[���z��m�ڔe�#���x��hVd�p0҆��g���:�U6���xwo���۩�ʦځ*Z�l�Q��v��+U��3��5�2&��;���$(�R���u+N9�{^$E;
+�*�VG0�C5^�3x�Q�%ےV�Ba�∪�V��?4
bڧG6ak��q;ZuQ��SoT����C��zf
*3��ΡBd1J��jnKyWr�l��Te�M��M���L�̮G,�ӴB�S�h�l>]�ӣ�ıJc)�]sV�t���oJ����ӭ���hr��%�[w2�#f����^�3d+[����^W�9[V2߶0ۍS%\�cN���&���%5������c�u.;
�wo9��wCtd�ݕ��ˡ��:s�.b�7�W;;?7O50�	$���b�!�"g/�Ku8s�zSe�R֎4�t6�^=�eh�J�]�`cv�m�uWd��t�t�I��VFoc���fT�ȝ�ڑ���a0#yx�XЮ�Tuڦ�gQ0藸[W��w�za��D��b޴s\�lK�o6K��=��tTY��.[Qw��˪���n����	�ؒ�6j�G��C I"����d!�g6Ni��������Cd��b�&B��c;Uy�9 ��7�B[T��B�q�˹��P�';����.��ۣ� �hDlP�j������E!uK*%��gz��u��×�4"I�-�V�.T��Q��h c"���*ofⴶ�9x��W��ݪ^��Ǣb��!��b�����V��gcy�T7��d� ����麔;�;\���W����c�Z\��
ǡ��j����Vz
�v��&�6��j��ðu-����Z1�y\6'ZvWl���w0��|�OC�Y�;36�6�����uH�%ݨ��Gp�+^���ܻv�t�(�Y�[��w��FՊ7��3E�b���BEu�ͳ�,Ȉc�u=�U��b����UL❅��!2�>B�U�H%K�yl;�	�aQ�әL"^h_P�Z&��	zef�Ź/&������aE���
(�z
��rj��z�YWw�s��1[��V�_�ŶB��z����p�nt�]�-�,pTu#�v*�6���|����#��Myh�;��9تK�g�U�y#�EX��2U��Y���wR�)݌���\��3�گ�5B�
F�]ա�͵�˽{�֡��9z(p���R�����]�Y�l��Q�O�Tz����S��/Jj��nU���OE��ݛٌ"we'�xL�'�6ҔD�o^e:�����(V0M~��Y$x�=đ}m����e����4Ӷ���ǎ�x��Ǐ\.�_jo���qgFq�e�Qh�����.β���Q���O\}q�<v��Ǐ=s���۬�⎊���2(����sb��{v\ҒB�SM4ێ8�;z��Ǐ������u�T%Fv6Ȯ.�ՑGM۷n���~�qǏ�x��Ǐ^d����J�BK�$�)+r�ts淳mn�g}:𣾶�Z�w�g���<�����;[QV]g����2��Q�e�Y�o.n�-�#-m_�W�fU��wdDwGtڍ�h�e���_��\O:,��w���v\Ϟ��쎊��;N�;�:���:mٝYGu���ge�[wy6�ˣ�;,;���3�YGu��)�0�!ۜF]��GTF�:�5�Ԃ���J�a�Ni���������Ǵ;%n�$����أ�`x�������Y���`�$;*3�f�D���ŴX|/#�q�����"S^�A���+5����Loen�)�[n��^�O��u^���^pL��14C�"琛 :j�
��J����b�������b�7K�S4�Q�6���ܬ�ʍ���~~O�b��F�9ʇ�(��kuC�m��tYy��z9��\�1E���H!G/����{af�ۺ� ⾠\[\u��;H��e����ebe����N�}�@*I˺b�t�4Up9���t�'K�h�Zj�̚�9����H�ѯ���^��w�ζC���0�^~d_G��'�ng��[\����k��ܚ:nV2f�>�;�� _�W��qBSО�m�R��\�Fc�~�{=׼�����z����}P�>���Eٞc~$�����6���cݧ��>����w�:��"b<�G��o���?�1�����D>H|�%�xmk쑑�#QJ+s��.de!���:è2�5E�a�fJa���}��DA�� �Ё_��y�V*��~mۻ����R�M�3
�k�{��շ����]�\����T:֡8�`�p[k^ʍ��S�8$��-]˨+f�J�1e�`i�~jx�]�Ћ���#3��<��\ތ}r`�v\��ZU��k�uխ^p�⸓�||||||��.�%HgzU�S�%۟$P�V��9�P�=`���&̍����j8���>:9ឦvd𛄦j�Nlj�3��p����`k#Y'���0��^7�K׉�nia�;��\|u����QY�(m)�e��o���I�A�0[�y����$(��G�U�P�ݏL��JB�\Zxs�|/���\{g�T�of��́8�/��-�-�x��<��kS����nDm���^4ux�!G�;~��ŏ ��ɦ\��	����`���?{=1�����想�w*�¢6^��NW�������Ёs����Yx/���0t��z��02}b',�VD_S���H�
ᡰ���T�(��U ��s�1X��һʫ�SQۜw��"Օ:�A�l���G���}���:�^E�B=P�|2!7s�'RQ�R���w94��6Ț/Y�9ҷK�o�j���H{h	���C)�[�_?���T��<�X�E�!��K�}�F�8d.ۏ��:�^J�2 �;����˟�1�J�,���*ߧӽ��h≗:��ϏՑ1�H n���_�L�f*Lc/k=�/&l�P�!2��ʹ�r��#��5Ğ�܎b�d]���w����=-C�jiY�z��gU��{&t[�o�Zi�(1n�T8�F'[W������o�������}�q��Jn]�m"��ZE�C��d�^���6.�|N��+��~���s��k�w����d�s亇�"{x${���-�;�8�9;k�N\n�2�r���ޘa%��!��.�b]�Bmw	�a|P�f���i�BǊ��;F羷5"ׯg��[����k�G��jUְ����rf�� p�u�7�xں>�E?!�`��#XÌn�Sliq���׊�^���N�嶡�L��ܓ�6�o�e�>8U�}ڞ������+�W��c���*y�i���z �r\��{�h�=�r�LD��mU��v&by���^���	��
D~����?�i���$��ߕ
E+z�E���x��uJ��ե��`�N�^��{0D���]s˼ `G�>A��������2Y���R(--[Y��ƣ1sEd.��-^�����-�s�<6�w�xJ���\��u�ͧ�.�uE������.��'�ִ����w�<�V��E�-$h���[��S��� k�M�Fƨ�U�.�!��=�"I�b���,d�-?�c �5�d��N\9��Xy�ȱq��gW����b��7�J��w�k[�I��ۜ:����Z����=��,�R�tt$�L���[lZ��l��*��s���"�՟\岪]lc�Rlᕑ����4�V^Y���̢�ڷ��TεXL������6s/���X�1��<��wY�w��δ@Ɓ�F��S �J�c�#@�������da��R�RԞvо�-�F�=�Ë�#OR�~�=[�/Y�k@m��{�Tx��Q� >7��i����؇X�TeCj����j�"d3¿�qC��v�^.��e���$�B�����1����&̟0��上���C�վ���;n�^�玧t���6��F�
��|�y]����������`h&H��g�i��f�R�u!�wN;ϵEL/�J.��X���8�S�}�Ϥ@m
�U�ǾƁ��w��7!K�L�"ύ
60�yD
V�WK�'�N[9AiѪK�5'���l��U���\-ټ�k��{?�1��ɗ\�1�c^�"��Uz�k������9�UP�0U�� �Lpî�Ԣ�&�6��������jّ-�#v��o)Z�T�.���J~��5[y��V��T�A��hd��>�A]򁣫�D��m
�G����8!�k��Yc[ǵ����f�������Ǉ@fq��x� "�&0�B�A�.��t�ҤfYP��m�m^�b�xC�T�mWv���CR�}S�qr+"��6�����2�}�-_����㾽3��0�ⷿ�����t���{LE��&�Zh�^,f��њ��"�5���1U�6h�f���i�p�x//b5�9�O���� ���n���%V��	h��s�f�����@۠�}M
�q�ELP3S<!�ψ�Α�P�4�v[�]�pO�|���ި�\�kcԈ�&{�����PzP���VT�5�nF2�$�]�G���A܂88�#(����J+�]z<��*�x�����S~3s,����1�fS�&_��.���ʮxeo%1���_�a�w�}~���΅�;��A��eIN0M1��g����]��s��<�*�P���_<���lҺ��kAopl�Eǧ��ؘ��"S[���Ї��
�z�E��!<�S����v�qn��A�0>D��C��!�����V�e�^�b#��rڍ�L�#F���I�%4�£B��:��=���M=�Ǩ��d�f�^&���
�LTP�{2�|��(x�E�$�"�S(�l�E��ZD�T���O�ҋ:K_J@�{�#��-�V9�R��ߚ��0>��
�/���I˺nI�Er��,F����dkQQW[�}x|�dO`�#�k�f�Ay�Q0�-��z���{%cP,@6���@��c���Q��*e�[6�1Hە-�Z«�c�m%{c=[Wt���/^�݈��L�i��SV�qG��Ɉ���W��}u��j֧�©M���0�v	sgub�ڔS��FbtV�maU���&�A���E������1�c�}�7��9�n�N���`�(��ag����<��YkО�m��B��s�hp0��2 C!*��#��0��\	����.����^��cCخys.��z|D�r�Q�wr�vϺsoے�Z���ѐ�1��r<<]�����?W�Y�雈H48F��Ø%�E��S�.��k��2��	n6����������6t���ד��U��-Ǭ,0�*���X�ߺ��n�J7t-kgkl.�%�_'�dd��I�_���
��;+�k��_��a{y[V�@�D���bw.�� M,t&���z�����Y�r�z.��'��y�e�S��8ǚ���<D��K3Å��ִ�����B8-p q���5F�/��u�'�]��P��'�_p�fL5wo��6�;��o�NVG�ا�eb�D��ۉ i<?�V%�JP��@kX�枕;�⎽y��M��'C9FC^D���-�<�zw�`���<��.&)�!x����5�l�s�M|�^�v�E�bVS1�;w!Z�1�� ��}>*��R&99D��G�n[Ϸ
&�kAf��
h���mż���㼇���gpo�X�S���;j���Fۈ�Y}'*�I@��7�)ȡ��ƌ�u�ⱼ3�.�((��o:f�nfޚ�i�'&gz�ۅ;�g	\.m��-�~��������]�c��U�֎���'\$��t�L؝�`x����yW���bn�~�p���=�{^�>����Q豝���&9-!�e�/T��fTa����h�c3�r���
�Lj�`-��65;��~�N��A(��R���m66٢�o�B��{a����1�P3�����������W`L���%|�=�$q�'�P��ӪZ���$1��2���]u �Wi�=�����~�?�g���*O�ڃ�����/
Z���ù�ˏ-�Cv)�:��q �b��r��r����K5��;�|�g��E��%�,m,����H�����I熠,ܢ��5�ơ���qr]��`�f�2��ݣH�HSW:�����y8�Uo�Zz�U�g���&"� �w��66Ҷo�ͭ�:�!�c�鳯�"�O�ȥ^~�8�5q�V�9/LJ�,(V�N��a�v��fndh��t= ��`�#�Ά�4�|O�fWQ��ɯR��L�Dxr����:��A��"2�[��m���Ǟ�:�!��#�o4IX@x��6&�|��3���k���
�'l�DH˜�6��K\�E%�*v�WUme_P����UY�@������E_p�WF���N���Зv^<���&�W���i�j��^�dT���/5AeN���۵�)�K�jHbm�!I�	���2����f-��U����S�y�.�d�i��1�`N_���g|�9��|pl;-z��%�K��h/B�b!�Ca|������l�&e���ò���C�F|��sW���V|���p{ڻZ��$htt����	^�>bA�;���Q��-����D��q1q%@��,���\����M]1p��ئtWz�E�4�UO<԰�p<��"�����/�
�KP�2-�r81�����2u��+m� �`����M/L"�r�~
)���5�l?�s��KFO�7���O�&zX�R{�[�����a�k��sH/Z�ǡoV�oV������& *|�Ux�60�!�"|��m��Ga�����`��/i�`�mRV2�sՔ��l���{w�����P� �/� ��k�9NS�N��^f���ݻ*YsWOcTS(�aO�\����5��0.}�cw6�CTˮFl�ͧ��Ҡ�7dl��W���0�0���x��.��NY�6>�p)���xV�s�S`Tpb�|��&6�@����'q|c����ߥ��ZPX׵Iw栜K1�w��~�8����Ug[��٠g�"L�����/r	��!v[Gt\lV���ɭgo"�b�d;XW��p�bk�# ���S�+v�ةr�`j�ն�0Z/���]{�\��Bz�Y����1V�e���㴏Vn�}��������&\��������:����F_�b�>W/�\F���{�dTa���Y�%#���<5v��牙̲�צB�{��9���tW�LZ��垪N�7h��o#�\���Yp�}�(q��}jv��a�K.�J�؃�`��C�~�.�g�Fu~�Q�AYY�=�M�hz�u�0�9Ë�}I��d��k�~m �I�Q{�y�7��D"�!���H,�v�54�S?����΢����!Vz���#�:�!萱;���\8��T�53@p��{�S�#�������t+�D��xlm]�"���4��%�� �$�4��o�w�WS��䍰�iJ�/�u[:�Br������޶�~��]t���,�����Zf�l��J��3Ϯ��s�y��ֆz����q�qiՉ�Ay�p;�'ɨWd�+vt;gz���r^ڼ̬���\�u`���{
��|�|���b�� �LC�J_����L}0LSY^��.�<�z��j��tַ}4^���0���V�o�[� �]X�an��<򳖧�ھ��AQ�,��!S8h�o����ЫS-t�c��K?_�R����{���;�~��b��de��d���X�|˴��vچ��ݨ�.-&��L�0��KA�u��NQ���iy"nY�&�Q$C��G��}G�����W+�hu�i͗ü�`7���SL���O�\Ycb�}����C�u:�t3_+�Y=�z;eB�qq��`��MBו�/c�$�aR-��4����,�2�����+����a2	��w�2�l$W���"�hL@eO�:�9�w���O�!1V�Q�Use��.)���(Eu��K��E��c��Bm��ۂ�Ay�K���"�8ŧ�n��u��Y�!�d�U9��5cY
d&�|��̯Ǧ�O��?O�-��Y؎qp�C-z��M7g)��7�!�l�TXn����׾FÏT����
��x��?fy���E<���8� Ӯ�V��!�Kwb/;{�ʩ�x�w@�-��|��I�����Yϱl��m��7EhQ�����\��	�� r���ߖ��y�>��
���-V�G@��n{y�h�ʘW]ח=О�hQ�KM@��W"�-�/�F����>2d��n=ONfD�sM��D{f=��Mx!�|Gɯ|�]\F���I%���~EK&zv5�-��ѫ�%�5{�2*��V�ӗ���O\R��{�U���R���vne1ܞz���h�Ε �d��;o9mK=�����&�M�lqqz�K��7!=��F訖M�Hnf�RD�Ʋ�&�B�{7l��J���2���d��=��X��i��=ەn�����w��q�G�r���x��<YidX�3�G\�y^y*�1f6��/w���זzrV��}��v�O]a���]�d��ya�����.�j���9�������F�f'1�n�Ipg܆\�0ꊍ�ɷ�UTKs�O+����$���[�����Pr��a`�-F�]T��j��nn���F�èf�qjuZa�t�k54��bD���Ӛx7j-Wx�em��b��KNnY�b�Bs	��WC���V�%1�aS9A�xU��x%�X'V��˿Y��S�X�R��QyP�����_(%C�r2_kUQG�,YW�'RF�h�UŖ�W.JL��1k=γA�5ʬ-�E�������z���E���θ����C([pv�����v(�#L���Wȭ�����+��}�;��
�B�|͈���l�fe�i��K̼�	��.ŝ|u-���2�Fs��ν{$����b���_w�򺫞�]�{cCy�7�Sse�7Urn�U�;�04����0H�N�`��1�
f:����˼��z=�2�Q�.�*���6U�Bٰ���c�Q
�F1�]ʹ9���Z�@�k���>n��X�+Y�7��or�x霴v��8I.	��>G;U��[t��}��^3��xmuNT�#�Uh�9Q���k׊����7�=@�^�\�e-�C�Y�M�ywO�,Q�Us�Ŭ3�1�r�s��FQqs1�{�T���Z��F�3�A.�s80A�FV�=gX��' ��{u���\'m2�	�+.�甖��^RwYT��7R:(����X�P��e:i�[���m�U}{m��Y[�V��֓M՗
.���D%( �ʻj���-�Cy.�1p��vn����g�gG�8�Yv���v�zN`�p����:���Nd�GEu��$�/MU�r[�6e[�5�q��AC��.�P𻌌5�;��ʍ��u�M�����E��Gk��e�#�ս;u�u��_b��U_�ͪ�7��;�9�����èg����CA�3��vL�a��83�Aײ��{}K�w�«Y�Ly�37@���g����\�[�ET[��Si�5�s �3[v�a8u*�cd�!<(���"��Z�
���2N�����m�]e̕lOf�f�]���+(��1��Et\"��U-΋��U�w���u_WAϔ��*�>]����yz��I9ۛ�Jta�U��.NRwxVe�iܕ�wgYq�E��Z2���m�Y�4��q��nߧ�<z���Gm����㲳��8�#��mm����N����qǏ;z��Ǐ\rv�(��T8��8��������uT%P%��z��8�Ǐ�x��Ǯ�d%D��!!Q$�K�;,���m�m����D�JJi���q�x�㷯<x����TI��� K(�:�+.�ggQ[����¾V���R���[c���h���6���"]�qqݝ�^^Q]�Tێ⳷u6��%�'tX�4�u�q��b�(ꣷfMÎk]�tE'q�k��Yq�Y�Mk�u�GC��H���f�ݩ���mimi:�����b��-�{�	8��J٬mg%����&�s8�m�eZ�ݕ���G����\�[��o{o�O6�*&�s�$Y$	�!L�4�l��IH�a�M\_w�.>��e�4�:\뙺+Y��WtݯZJ����1J彷N�fɼ���W�룻Gss���9.$��˄���~1B)��$��A�L&��m�F!h�$ �4���.yF�)��	R!$�$�QCl��i$�
�R([rBSA����������
�n�R��D��o���[�`��HG��1S���h���&���C7zvE_�������|�vIz�Mk��t����f��u��8� ��k-WE����|�e����P0��N���T�f���֞�鸫J�2��>+D
�S�V�zY�Y��	A�Z��謆����8oCuMJ� '�g�N%t7 @�&���z�TK�,���r��@�6��<��6	�i�+�ۭ�g��}���^���-��Q�"���Cf9��sG�A�J�c��9�Ғ����Y�닸��4��m�Q���}���A1��q�\�� V��yЫ�tm�1���O5��¼�x|������S���l?�aNd��Ɲ�B�|=�F�옫����g}f��Y�s��|�[=^a�����_��,o^�f��Sx�}>��NP��	���ȣH�+�Aޟ_�%�!mU�Ѷ�ǲ�'b|�ʴ��Td��Ũ!7��s0�H[�����[}�+캖������-����E'�1B/dY�)�EjM��M��o����Kn�s<3�t���V���.-�bGXa�x�{�7�F�S�~�5|�:n�z�1�c���rw�_xo>u��#y�"��[˕Z�1J�d.�tĴ񙘒�4�Uʮ��L$v���1؟�f��q�:���Vv�l^*Ƭ�{�w����TX&	�����\�@<>1Ìy�&�1���7�u1�-���]g]�y�Ճu�VO]��c0�灒H?m�{���{�I3�b5:��v������@��I��'a� \if���xLُ�5ϗ�f�9ލ�	
�|�s�IIs�hh/�/��07z�R���ݲ�^�׬�m�a+��Y蝽�G8͸�V�ud�ɕ̛��N��e��Z��ɨ~�>���9~�> �;�[v�����8t�[}�f�����t2��S�f	�_��Jm���pWch���5I\��������n1)��>�ם?�%2ω�O��Ht�l���� �Ω[�2�a�iEf)�X\ї��Uq�+K.XD:Rbm3�NX�U�9�8oV5V)EL3�K�-ڞU
O{![ec�7Z���А�;#n�3�Y�px�����B�ؤ���ŚsVӝrf]Ͷp�D键�&)�r�"Ƃ+߇�������7]�\ܸ�l�f�hτ��h�'��*t;���Q4��p���r����y^㶃�`�iF�ls��ا��\k���N��T���F�l�޵�ƳҀ�dnt
�ћ<�)E!�&}kw�xɬ-@K�ý�k�_�֍�
��W���?F>R��I.�/(�-N����q�j����/am������Dv�����|��63���_kA�I��[�0��j��,�2o���?3�o2�w�<����� V�+��s�(�i��;Ԗ>E<���[g<�@���� �۸��h��;��/�;�b/o(��<ހ�{�c>α��̀G5��Ț��qB�CK���d�}_�F�4��~��M؂���&[�����}ӂ}����Ĝ5��>U�ⶌH�FI�q�$�SlavNע�v,�{����
�R������{���8���C[�aLa��rGsJZTX(������ ����Ěu����oP�V^�Wx����E�]� b6�.2�J���f3�5J�9#`M�u�X��Ԣ�1��cƹ{���0���Z��A+eWO2�K��v�jLU�yl����m�ơ=�:��>��ǗW얰��mT���UbK�"w����oa�e�]�����ݡ���'����қju�g�� ��%a�[� ]ϰĲ��������f��*�A~9=�Ռ�͏ iLt�;�����aW��C*(@oײ�[E��06Z�2Ɵ��n]������V�{�<�G�%�P<c�Uܪ��qGt� Ύ}o����ό]�~D��E8*�&|C5K�K@����4f����Ĉ+����	�%0*tz��jw��~#�\�ͳ�M�,x��俷v��9��Ez��6c߆�8���Dp�>>���b�w:�Z�g�B���ΘzV w8̹�F�����m����U�S�QF���uCW={�fw=�F9.�Ռf�3�2Ӂ�T���������Y���K26wh�N�L�7}q��d�W�fK1w�[��z2�iN$,YX���IHQ��lX�k9@,�0,�O���h��\e�$�!Ц��e� ��Ŕ�k��o�d8Mt<�+����c΃�}k-
o����7���G��
����>a����A<��G�UZ:�}Y)6������[�����
doMIQ�S��|��7#m�!�_[�#���ל�cf�nװʗ'tV�7��Z�3�B<��L�����\�o���	�wu#ǫR���m�8�3��aU>xS����0Ǔ��݈>/���4 ��\�F���H�x+"�_3]�qG�nu��h�Ě	'��_�
`���~Ǉ�т���SE#�����2Y�t�G��fl�L�{�����i�ȍ����Qk�n���'�u��s��!�jvV^��A%<8�Ur�U���".�h�|�!R|�V+�I��-���o�Z�l�h��c�x�����MO^d�--�W��h�ܱ`z|��:>�uw�H��mln�^k�6���Ò8I;�u�u\TK�����j��s���n��n'����ާKe�]d�V�m�U\��V����8��h|�07��ѷUU���L:�����T���t"�7�^�_<�]t�kܐE�B��̽��uv�m�ӹ�kd�-W9�v^�છި�i��oR�hP�՚�'�6�L]dS��1j	�� ������n����=.�I ��sؔZ����ّ"ܥs�_O����\���C�7Q�/���~�>�\�4+�����{��&G��(`��y�u�A��U��E�C;�t	欂�B�#]\۠����_^z�.�:��v�y���۠� �1���Ǫ�gեU��4i�[�c��;p�>N({���%4+W91TX^�t�ׄG'=u�j��\�ֻ�Y��,|k�^X�k�A1���7� )���vo�a�>rV��O��7�K��2x�+��}�w��΀�{��pn�J^`���<�?0Ł�za=�}z�}&j�F���6�N��Q�}���T�_`����q'^�B;��3�/5X�f���o�0�e�T5*x�{���g���C8\��ؑI�/�zw���PƺJ(�`=�*vRN�/���ޚ�1EK�5Ǉ�j�zo1��Y�k�d���R���m×=��v���m��tIU�l��ۼ�,s�u�e����4���W�겧Z��C��W8=��K8��bV���j����Rq}Eunm�P�9�u��Nd�`|c�0+7���v�@����XdDԪ�ȼ56��#m��΋:�2a���45��>ډ�fLAP.Ms0������{��ڙ�yS�"2�M�1�u�4��.i�b3�q*GuK���`��{0!�%n�Uӝ�6�`�m �ȩ�/*�c���g�^�aaZ�������Z�twVց�mc��z$�R0��m��m2@�g�վ�%13�d<^Q����yJ�y�*���8��Ub��W��G|���xU����%{�%+E��Ћ��d��.�}�9��J*<3V�5� 1>��؝��F�G���;�=Y���2=X�+���R�i�����1���hs��g`�Ｇ|��nT��p��Lwl���6�:P�G�����ܷ�us�W��������9�?oF��o�����������0x��e�b����wB5�b9����^�(�,(O&dm✽ES�����әE�:x����T����w��vͳf��ӔA[i��ެ��\3P��w�y�[���Uw�����e���;����'��>>>>> 9'�b����=A$�hJ�A���o��C#��}f����
��:��!8c�I�w���#p�nJr=�~|����:8���=?��]��
�|�&D�5B�b���=_a��Cv�XBj�B�H>w�MWm�ޚ1��'V�1�* �����zJ�,^���3^�f|H'�x4�g3x��9-�qū�Kơ�΃�"�9)lO�(�boO_�q��۷5����������Q�]���Ȳ��ү}�d�
'z��)P_O+�}���s[����J�Q��ʩe��g�n�6�ٕ
��i�Yw9K9��\�N5��˽!���'��sٳ�NdPd:��'��dϻ:Rпo�v�8�s�.��JR��;W#U�f]�;�6uwo���Ѥ���>�@c���k��G!:=�����EW��F��);�G�㸗�|�]�]�m5U}wW
�.�M�;�'p�<���q��K#T��tU�Μ���nT,Pb���h%���Ω���43.4��פ�j9����֌V��\#R���u��;�w�^���k&M��3��{�0��~����&g{٩�h�ON�FS�xhM�ҚF�U(Ȼ�Tb���/BQs ܇*���S{�zJVt8Lj{#���bn�n��1{�E�J��z�|{m�A\>x��lS�5��pb��g�XUCZ�ޔ����ֻ���V��`��������\�QQq�vP�ʋ�������Z<�G�K���t����UϦ���vw����'��a'Gc��)`W��BJ�S�5z�N��4^��M 
`���3��d��0�i�q�2�t��[�e{��oT;+'�yF֣��:�4_�x��f����X����.��QN�`��0NX��e,�}�^��X�@�L����1>ǂ�w��X󇍌�����P�^Ir/�H:�	�^˃�C��r��^{��s6��fK��f���3���o�c�^�o)����j�U�u#E���+��9J*�;���^੧5��ʺ��Av�uM^o���^L�m���u<�ͦ�*<��d}�XO�+hUmQZ�/�~���<U{޲#a������˒f�>�3��$c�s�S
����$�ZZӈ�Ùy8�is&�]�pu�ZQ)V�J��E`0�������ջ;}�m1a�q*)L�:��OW��
�����\+��C6��Ϩ�vó}�ځ�l]�T��J}t��Z���E_�4�ԕ�l�Wv�3vwd�l��nF�jg�p,B�LD/J�7�����W�K+�*z�>ؗ*Ļ�O7�����W=MD�3����s*����
f���)���ъ����yZu��fG�����g�8�O� �Sّ#=�Y",(����2��M)m��ݙz�^;"@(s�+���vCU9�����UKҽ��M��l���i�R֊�J�=�W5��ͺvz�b�^ t{R�,�=�w��ˤ�g?OP�WWǟ������u*�l�yRo=��E�wl�w��Y`b<�w�D$�Wi��ɽKtt��9��t_:d��=x1jj���L��ao�	t��VgҲ[�|�k�	[Y�^9�b�7S����GU;�4x�sL�zNa���Ƥk
���j�t�3C�"8��e �6�r�VT���[R�S3Q�:Q��+��>t$��w��ص^җ:&��Qxn�}�p�W`�­�H��l���!�T�M�{�(Fҫ�
w��Jܳ�u,ۺZp�ʡu�]����.,ƣA�7�f�w��q��F��C��omc���W�ԧv�1j�"+f��e1A�	��\%��@��ג�Uikm��fd�ʒ�kʠ�a�KZA��1i��T��{�8� �)���T�n�ZĂ����f;(T�R�ݖz�of�JL9��[��&�:���,��*8�}Ճ`���uT�cx�q*�v�h^�e+B��j���#�՜���z$��C�ob���UWJ�(IĨ'e��5�����nӷڝG����3�N�;B+�+��|�(����6,�r�ܔƽ�'&t=%2�uJ�JJ�L�h#}�h��J빂�a����v�s��AL�)�����\:�c,nٓ�u���\u�*m�ʼ��7Wf<��1
9�^Z5��5��2�tt���y����h������
8-Ay(���X6J����6N7cR�9X�̹�%]�d�b�F�ZXr��-%�h��W>��<L�+�uŗ����5w�,����s�b	�,l��f仸����m�
��I#&'�"���U�$	����}��ݝ����Cٰ�N�׫2��~�����|A�[y�h�kn�`�E;ju�4��A�n�gf�����|�pܴ�][/��R�1a�3T���+��yvq5-hR���gGݎ�dAYS��o�qr���%�A�X�W}u!�-ִ}��ųs�S"�B���S���ŤV.:e �l|�sD7(B�3�KK���Tl�v�^]ƑƄ��Q=��뚅�����Uq.���cq�n�X�j����`f���>����#(���Q=���<v�y�
�z��q�He��E�Qz\�Λn�va��2���V�ݻ�Me�c�r��3�����ؠ�ɽB�,���U�ÝѸ�X�ܹJ���dd�ڪ��l�8i,6f�l���-���/kl��IԳiV���v��F��$��l�A�l�+F��n5.�tœ9>T��R�Ӿ�9�iVU�a��y�h���d4�"�e��7V��{c*oIW��y�dx:�1�qٶ8��LOI°n�UM�W�v�Y�d�9 ��N����7Z��rU��G$��*ۦZBʄ����5�����7a�O�Sw��Ν�Ҙ�xN8M��/Fg\a������͇�iޝy[����dC;��U����&n��x	��SU4"��%m`�R�8�q(��ݥ2�l��r5���(㭵$t-��mu�QJ�Q��i�n;x�Ǐ���Ǐ^��a	�	%QjB�F��rVY�ٶKkq�$Zd�F�J�dcO]=q��<x��Ǐ={�;
�P�T �J��Kk C��v�ݥɶ���VYe��dvڤ�	D�T�4�׭��<x�㷯<z��2H��(��j�	!TT��Y:찠�;^�s�Y(P�tnt��Z
$@��i��޸�<x��Ǐ�����d�$!���~7W���w�q�$@C5'��(�"O��ݙ͹�v�����|��$�희k1�j[Z�$���8I/{�v����Y�*<ױi6��:�՗Y�[j�mm�N
H��6�{I�j�0�Jm�eiS�I��km�ۥ�%�����q2Ԏr��ݮ$��f�Zt�s�I����I#4Y؉��K-��E;8��r:$���,�-�����4c�{6%Gfd<�v�0�ۤV���R_�OSZ5��g�ĝ"s5	H='ll&n&�6�q�s��3�����������+��� �n�TD_I�Ʋ<��A��o�h�r������!¸���s̯�D�$�^-rb��,��gq���gn�'�}�:�C��=Gs�b��M�d����'��Ԥ������g�ƽ��wu	���ѿyEO����I���n��GE;<�}�^rѵt���%�y����C(9�_:%	�.���~;]+�_���>yJ�q,�֩��Uu͸�] H�1���@���r��qpu!�w!��ޜ�x���U�G��Kߢ;S�j7�|m{Q�#��7\鼰�š�f��UC���>�	o�A�;�dYk�p�������m�4^�ڊ�Z�*��{$�\T��l���r��E%M0��n4�G�p����qG�����%A*�䠩���n�4�8��r�}��K=����_�`���J�vQ69�[�胼��t�ӥ=F{fjZ�����;ga��e��]�TP]Bgy	�P�ag��.�ma����^�mB��OqNF#�EM���)�q%��2�����9F,Z*�iJ�P��(F�T�'�3,�^��R�V���ӧ̫ȅ�\��J�����0`�60k�ta {߼�o7��z��a�v��րW@��y`�-zJ��I�U���^��ĪŤE������£�n�jMO�9�pY>�U�={��&�8��z��-I	�[	�z�V3xO$p\Ę������O�u����p�b�G^ޣ2R�u�����JJ>�㫦�u|�u���b})��H�v*��Ș�h}�����]��6�.Eo�+��<�35)��f�ؽm��`G?��'��޽��V{k��e!��C:�W+���{q����}��ЄK�=B��_xɽ��n�+`EG"\��Amy|\�}ؾ�<��������'PD�C�y;�g��^6��`�jg6_}ip��l\Ǩ�y�T�L�=1\�ۓ��5vn��'v��BY�FC�{S0�Y��қ��6~�����|�J����}���2�[��t�|�鸥�tSy��3�1'j�R����]~��Q�B�5,��;�Xa�YG'�Jw����7j	���PU��Yn��HR̅a:4c���4�E���E�s�ʁ�%��Yg"`��z�P	��'V��,3tF�fL��V�x_�qV��gSY���90Ѻ��p�����uw%i��1�bwgr�L��+�ٽ�۷�s��FD8���͆��f|�����n������R��C �J�Q֑�JE�-��
����&%��A�Y�7��X��T�q&��턏5�/��O��*/N��XV�L���满�p��> �́ؠUϢㆁս':������A��=��H����hc�2|Q"��1�!�G#����ʼJ��Z��qd�| O$ߪO=fE}�<%�-�V�4;a*�G�5M�4oJITU4�5�D�oL�oF+4^�M��5ƻ�f[1��p<B�#i�e<�Bs}�ܰ���ޱ�]�^�K���l������U�;��68C\$�4�	�\�j��Uɸw�c�a���W��y.�仵O��<�^zz��Q�z���=�ͯO�ځ��³�*�MH}ު�I^�L�NN�O�tF[;�ܚ�[^^T@��y�q}�eH}�!v��j��n��h��3�h�E_�sg"�o�@#"�mNTk����K��'6�P��,�u�'L�S��}��].F�ǽ���Y���u�UݞS�{��_)�j-�j��.���5��3u���1���W��w8��.a/��c�k���77ߛ�48�LC�#޿H[uw�Զ��N���Iyv��Q�|;��/Q��:��|h1���4k>�꺄qK1Bt��5�:�q{st��<�w�]^LU �oV���a�;Ѕ���[��C�,����&U�;l�.�����}��5��ԗ{^;�b�t[�3���Wv�U����(��j o�����dUm��/o�
UB� g��r�U��ڙ�y���yLU�n2;��H��Z�*��O��r��#��yEi��E�bu��^��h�Ǘ���qOsi�����$F{>u^���� ����}�Z���RV���'����.�wй�.��R/�?l�)9 BP(�����Sw�[���9��}k�׵����T�I�;��ә��%nBX�PK�ݼ�ퟻ�d;�����{l[,����6�s�X� �9���yl��&G�r�D��۾����Uk�Wg�8η����X�ƅj��v����;ݛE�&*� �)Z�Wgv�jP1��ɧu�"֩���n�V�e���ݪѺP���Q���C�M�z����e��R�S'2O�-�p��^���> J�w���q��.WӴ�L��o��\H�F}��tå��[�����c�4��W_��>�ܓq�˙�_y�H�]�y�k@�h�֪Y��cMǭ�ZG��]���L�>�b��� �>��c#HhqU�q@컻Є٭�Z{�i�a�6�a��.���j����?q���Ǳ��$�s�*��NE������fҝյ���Ѿm�o0Şx�*�uo���\��l���廇����,N� �c�3>��(��NY3Gu���s��ް�b��E��}`>���s"��s�^�N�/�P���1�}B���X��瀃��K|��y�����cl�:�gr�7�b�B&ډ�w0�S�7���*��y>�ƽן4Ŗ���D�{x4�ڤʣʲ�ż�ul�	@�awDn�5ꀵ�/K�[�
�ؖ�|�)&>������7ʚx��ۻ"�'u1^��l�Mu�G4cM5yK��;/��.wC �x�G��f�ɩP�D]���Ĉ;2��t�oJ�&7]�m�ø�]!VƯ�l�q��t��x����]9�il�}������>>>>>>��Q�\o���!~"z��1cN{_ו��p�S�����i;�<��Ԣ�c�;'���k�y���	F�;��6_��:�m�e�P���Th,k+N��=l!�+
�n�9�UR�%U>�ϧY�	�w�7�x.z�-�\���}�*��,�0t�炱Gh��6�Z�(��x�ܒbM��H|Y"4-��*�ݽ:�����YO&��&gg�|�X��|sь۶�P�j�^���[�n��&5l�����1�~�5\�jc�D��Usb*��I[źB3 �h����k1U^�5��@�*�<�
����/c��-��?�T�n��8��3����O�y���<�&��_.3��;{�8}p�V�Y�SBS��Zoȥ��G
ˋkh���>�{$�>B=����;3�.����ۊ�|k,q��h�j��Ww�9L?�h���'���V!�c�k5̼��2OH8�v�K±=�G���N��{�rL{�xr�]�}�]x��UO�Q�Q'��y$�Axl��i�`�=!˔6�q;�jE;[�ejV΢�VU�R��C���L��kL��zZ�:��o&k��e��>>>>>>��ץQ,�J�f�A�����6��ꙁ�*ܥiU����d�����~a�+�-q�X��wL�ᷞ��ݵs��:cfi��akԽv���9���³B-)�ߙ���'ͻ��~;%���Kq�|���>5�b~��۹1�#�ٍ����V�;?����
�hRt�Yn}����W���nk���
�O�ȐC���V%D�n�����L�BN,ꝴ��D����z�n�@�g�l;c���6�bT�c�c��O��.���~�֔����}�qQ�ˉs�n�NK;,�m�w��5��`ǲpJ��b��U����t����OM��MFbɶf�������zm��U��Sb�Y����k�!sP�j���pa���Y�wo<G�l���o��R:��E��~}{�@� 5��͟^�'�����"�� ewd/}��W_Q6e�6�WNBَ@1	���菢�-<���p�5�l*��ƴ���Kz�[+N5��1
f�]���y2:"-�ÂSu+�(��R�k����U}�O�=�ݳ���i��^��
�sn�BB\UaL3���	̺3{G�+�ݝ���w߀>>>>>>{���Ĉ����o��\W��5�����S��kqi�3�8�Vg��S��q�H�}7���dWy���v�`LI��v���>-�+A=R���U��2yW�X��aNG���-��o�ޠ=S�1'-NT%|�5f1|�p2����؍�[қt��[�g�	�Zy�!|r��h�5�}F�He~�k����#B�L�jY8�UCd4�[���N�^�(��|�wu��@T�o�4ns���@8�uF��[c�25�o���dS���31�G|�OhH?X}�[������| �z�^����*V�/F�M *��<��|��=�,�E������L�����ô5���齭�~�v��)QU{��K���\D^�m���/q ˷��?+��Cc~��/gy��\�@�#�P�z1�/�A6C�G�q���PU����]9TK�\6o�(FK��P^y��R��#5�b����79+E�nL�BU���YY�n;�/$�.5[*h�������8#�,�b̤�]��]�q�ӹ�+b0��M�8�MSΊ���b�w�[�D�~����y��'��糱�*�\�TK�17t�ÿG�#7����Ś�:�ܗ�Ԑ{�L���� ~ޜ����>l��x�\���&����aR$>��[���݈#!f���T�%F8�=�ܧX;2�r���j���s~�.��10i���d��+א��pz)_<�+�zC��S�v���OR�*�v��4��$Y*���
��+g�F�\pc��\�"K��Sw�O�q6�[Y��S� /�<�)7���j���F���vgTF_7Q�=�+���f��T��.A�:2�5m�j�o\�O}c/����m����a!wn�+j|٣��s�c��W �|P��w�3�޿Y}�}B�ٍs�X�&"�DԽ ����3�~[���_@A��N��|�za�4���ǂa�&����/�M�ȟV�{'H:L�c�o��y��؉[��s��4�.S�X�ĭa����dM�1tY��O��7�q�&��ݼ�n4ۭ��쾫$�dq��yj�Qл��ˠk�v!��vn������6�g�t��I��gz��HUac�������x�tz�ɫ����������Kn�9�fZ'
�xg@)��&������1��_�_W�M�FDRsp�e�Te�� ����ﮭ�`�����x3�Q0C]��j��Tٽ�|9�gue�c�j٘dzD[K�&D(�e�c1>�W��n�ow��g���ڛ`�j>�s�.�W&W�����C�0JLnҸuds�,X7Y�z����zh��n�/i�I�3�����w&��5!�	[�r�ݑ.��� �t�#-�Q��:Nr*���]��R�L߀|=���a������r�����lH����0���KI)PRUP�s�P�F�SNōQG:7��c`[�ں^��[����D�炨b��<mA8���&֥R��i�:{���.Km9��:[Ö\h0j�pZl�W�T�Mͫ;�3)�,p��q��U��:���$�����jپ�5ɐ�	������㞊��X\1m�<�6�ӚJ4��f��μf�o2 �rj�(��m���3��ZC�'Ax�$��+ =�����p�������\�r^�T�V�'q����8��đ$��
��#*�l���բ}��Z�����������c�v���$a��֕J�1L�L�cP�PZ����nU8�XoQA[}h<KzF���D�*eMTT��s+i���[a\�݌��L�K�ͤ�*�0L�(�2�MKcLb�A�͗Ug5zK"�\a)cpc�9�a�v�Z*�SY]�b�tR��ָ�Vc	fwYK��X��s�u#��������3x��uӋ�L��רDn�oI���.�y�
�W���aJ��f�;Sb�07p�x(�aGU���7�Z�ƣ��}����lݑKu����Uz��rR�YvT�',"�X�VD�BYv�2��[J��14����WKڷ���#I���7iIƫ9L}uu@��/L��Z���($t���Uk�̨��ar�u�_f��%Q�ک�:�vk�y��1�p0�WY�ފiX<ԍu��;U�qhf*�{B�nuQxhUYxp�U=��U.��x�
{�:���U�J�>䝲���it��r�Q[~w�רfں�9�ʺʾ�k;��n�9w�M�׫�`�ϕph=��H�S{��sצ��9��5B�zۏV�r.£��Z6�mX��M[Tsr���;���|��8��1k:���şiG(����M��'�����2^p����UL%�98tP�iԆ0��j!��񼛤�3f����+�($���Z(��ӵ[������e�Aش�ozi�%W潗�-�{.���;���ZÚ���d<oP�װ�K�ٳ�<�����LTVh�+Q}���\�ŷ��b��U�Է��R�eT�L�{��8��)M3DxmC�}R�7{#�g'K;!�^řX�N��6��-��p�ӹ�]Ժ����B�f���v�JC�޶�e��+y\8d��|Gm�I�V�Y�>�y�j��ȍ�� *��I�@�b�Ě��!���h�]`�u���7BE��w�v�2�E���12[3�,W�n�lH�7ϣg	�%'��L�P�U�+�;[�h�&�:c7o����]ۛ�!˷]�C���p��Gml���\�k�V3�gN�b����u�K�M�(�ʥy;�5��H���K���$u ��wYt��x�yD[���J���aF����)긫�Y��
#c�uo,��w{V�ruO��%���c5uټnŌ�F*?�Y����X��D�IT�y3��۷v�U-�Ź\��b�-P�m����R�p�}��y.�.Kyu�6�b�ٲ��$���m�2�'ԓ7Cקzh�c����!cD�[��ޥf�S-v�t�C��U��	�m¥����������{ �,ܣ�̂�6����:qH���i,ͭ�~7������,.v���v����v����N�B��HIͲ!����m��lS�6�ffp����e������l��,�YZq��׭�8�nݾ�v�ǯ;�����ڗ֭��r�
�m�gv�d���9Ӷ��)��*�����#O^�|q۷nݻz��׮dgJ��@�J�UT�J�$"��[i(A͛����6��nL���9$rm۝O^�|q�nݻv�۷�\� vT	$�N����m��f\��vړjl���g��n�e���p�����m�dm�k[sA�iu����w{F����͚6��\Fۏ׵���t�c-�Fͻ����m�m� n��wt!ֈ�XV��j._��A���'nD�Ȏ�9����;�qX8JE�Vج!&e�.P�)��vL�Q �-����P�vw�Gg1���wQ:��쳱�h�H�BQE���Ϛ�w�ޱ�=��aR	�,/8SM��`�	F0�(�
8���*Z����5SE�5�
��ɷ���u��Sbت�.L��tj��mE��mSS"��J��Eu��z��(`QK����Ì�؍��9!P��I"�$0I��T1Di�Ҍ�#llD!E��R@�$�H�Ɗ��LnHa��E�(22�����`�$�w�������T.5״�ʩ����VV�Y�c1�X�]ӗ����7�euOq����r���Ϛ���{Ѽl�n��ל_5�H,��mŭ/�Ku�!Z�
g��z�
6H�\V�c�F�<���mw�xo%��50�I�>͠oz��x�P�WNoz9�2�,�p��]V6H��G[��-���;��2/��-FMT�yO(���C��i����ŷ��r +��b�A�OB�s2�z�<��Ui�Ig������hGt{0�^ҡ[���ú����%X����-<1���E�FE>������oqE�}R_z��z��nwS�95q7�#Da�s�ʋاf�4:����N�<���)��9��i�t�ީ��>�!I6�u�fқ�!W�[�����ͺMV�����
X3�%�i"�N�K ���^{_�i�^�̃>zγ;�u��N,�yR����4t��A�
��$�t?��|�=��iO�ar�J09g.��=ٓry�Ϧ#;�7TÚꔾһ�з-�Щsl�XĦk��y7n�^�S���x:̤���_u�y�hW�x������sw�Ű�c�����
�и⚿[��u�ǽ�z��Uӧ��R��)�ۺ�F�}�ߦ��@�$��B5�,m��'^�7t�Z�!QԹ�K]����w��3�[���n�S���SF�E�VN����l@6�O\�k����zG���fu��7��"�gv�Du��8d\�֭\�x����-kgd,���S+΋f�O﷣P5�� �ꘌ��tl֩�Z�&���j��3�v�I�� ]�g�ulU��x�U�}�0u^��7�{�;ߠ���pi*B���V&��Jm_VD��S��k@�����ּ�A<7��ۏQ�/�v�v�+�y{��V�������3�{�l��rFx�<~������}s���$$�\Eˤ�ږ��U�����,d��L�ƾUq$zb}��"ʐl��U����m�����1��,�X7����َք�p������Sh^*�f�"d�B���
Y%�g��+3���Cp��]��]�X,�w�=YKi���]^����w]n������9��D+�'���sU�=�S�c����}�0��Q#ִ���{:���l.���SŐ����:�ݧ�x����@��?mw�7���|������N7��<r�T[��U��!M��7���wAD�`*�E\Ȫp����A%�AA1�P"�!�!��]�ևӓ{6��k�^,'�T	̷���rG����to.n�1y��gSu�A��p�МX�z��]akA\X�>w�@?���^����m/�۳E��d/�&uW�E��4�x@3���B�O������IԚ.�}`6�l�{�����c�P{��N�vdzE��[b2��./,��Z%{)ס	�H�@�{�K�t8L�����WS�����F�o\>���ћ���fDB���gL7>�����h��U���\o_<�����.*��Q�6}i��N���:�'��|�P��Ϟ�"w��eDČ��_{�:��[*c\;�."�	�=�^:�FC��D����2�'@�tU���!$�Haez�'��o���8��q���ER���q�Eh��-���V�u����٭�Q�jw!�eQJ`�qU�������>>> ov��3�� �\�<���xu�g�6��r�g�MΚ�`�,��h������Ksgܦ��J����m�o`�`�⦄_����b��-� apug�����y���ߖ�k����|�"���پxXN��/m*5�z��~������zCv��J�UTrf�{�ֳ����1���k��U~k�XI��H�>6��yᲃ�f�����n7Z�/
�<�������WO3�G"D�"�k��.W��'�aM<$����g�=!0�����"+���K�@�Gk�-�i��l�GxY��7�[ois���g��!(��ɯC�ՂzN\:�T�J��r�vO�%#�ͽ��S��J:���!�cw@�.p�Unn6�*Q�l�����*���BҔ���؝ �GRgυ�jWh�|6�D�ܤ�<z-A�nw5�)NT��Vs���oj��ZY���V�k���4g����9��;�jD����l3��'1�湧�%�"�*&ru�F�V%6qF*��о�<���ճ}I�ʲ�{ǰ��.��l�ߘI�'����1�U��g[�d��ۜ�P���35X�L��d�E�ˡm�L���Ra66�O����ք
Y�#�:$�T�T�l�gv����ho
Z��wYq��X���"s��'��^�=�.Zb��������k����:��yr�-c6{|���"O���9��gVGO|Tc�M�ܫ�m���!�eշ�z�0w [�r����m���2U��͞p����*��x԰��_����/q�cqÕ��^���\w��O�T^��;���mƕ�Q�$+���k)�S�^��A?]R�5����o%Ո����b�e-��J�sVMN��U��x�����7��٨Z�n���G�p>j�>R��/�4���{���q2	��_�g�p)0�F7�!��1���P�~O[�ˑEB���=A�� #��X�6^�I��\��Q�r4odΨ�������˂�;�Ef溕/9��9u*��'7H�::�O1"F���+�	�3j�����]���y��NƆR��{A_����s�\�VE���Bs�OM0�D����ٜ��M�*F6�y��o7���]�\i5�a�RE�v	S�OӐϡ�+������U.���ZӘ�ӵ�����xQ���n74nr����F��X��Oy\ T�w&�������E�_�J�7G���������(�����CQ�h�kD�70�ܫE��Al���v��\B�(.W�mW�'�<`��q.����9���^��^����"@X����oP�i%]d�1S�7|f[�]u�^�N�|�ɘ�oР����u����6;&��U��9��9-��l�ę�c@���~�t�K�Y�J���ڽƋᛗj�[GH�X���νƩ+.x�m��:��f,������^D�{�s�~�g�B�[m���bO�g��ҷ�	f��>��W�.�ͨ�V�-p!�\�U5b�t��n��{��m�K���.������,NB�ig=����ؘ��݂ì��w���8���nځ7S)d����{P��6�ʺ8 ,���x�Z75:�|f#7�dT����M��aB�.%�&���EY���'�������y-�Q;��g��73��N�x�c�1�������މ�vk�L��� �t\dDgyT��n���S�w��>���c:���88M��B�����ћ ���Gf2��ib���G;x�I���M[����+ˍK�4���c��0}ʇ����:F3YH��gʢ�;��3�;���_���u|�$��h2�Fz%��W�0��r�-z"j����L)[=ʽ	����Q����)�xP�ɢ-j�����"��d<�7�O���h}&RB<{�}<���a|��*"����l��$Z��h�U��+Gp^�2��*��e��\w�Lېd��U�M���B�{��,��˽q�����Ȳ��1����X���*��>�⢢\��dX��u�U�1�Sa���u�^����&M�0`Ǩђ��ӷ�:i�i�����æ��x��S,P���۫�v�|��0�{z\���G1���ZؤΛŘ��pk/sKU�w&�l�N��/.���wTq�޳��^<�l;���RC��q�6X})J��
į6���]�bC;q��e�֩�9
�,)����w�i����>>>>>>�6��݅�ӿe���E�+�s�y+I)

�nhv˫}����p����j�Kñ���t�g�5j�y	u�rR�sɒ����E����)�!���6�f�ϭ������X~��	�[�^����G] C�6�X(|�*��l~��n5ӳ�l4����|����U��h�&)��>I�*�ؖ�xw'9���Ĵ*�0#�ey:��	J�ԫ����ۋ"D�U�\�yΧ|K~��}Y�?(�j�q �|�y��}<`Y��J�Gt�D�~^�rQ��Vq�Ut����6|�Ǝkj(���u�*^�n9�@�<$�g���7�{~ �f�������u1����ϵׂ	��dE���P2��)�g��w����v6�Q�+�N�DZ���%�j8d3�7h�}������w�Y�����Eg��A�0��E�
W+w"��*�Ss��<T�c%�kN��Z��A=}k��B�|��6�����2�7i�aP��zv�n���
�PFZr�7��WMĵ��9Uf�-�\�`7��Mj�8ғW��|@>>>#���u,u�+d����m�L���A�Qz���mf'1��
W�	핑��q��C֫%�ؐ1 !f�x����r"��n{+}��Emr*i�a��Z���JDX��p����|+fp��K���j1�8���^,�^d�Ǭ��*j%���!t�*�ȝ/6b�98�z������6޽ �)M&�g�l�S��^��v�+�otg2���x��z)�)
#E,�#�gBT	)R�����	��5�ݢ#���]6�3�[��N'xD�-�O3��Ϯ���S��s�asqG�on��	Y�����?�M�:���=\_γ�C4� ʸ<�o
�;�W��s}{��>y�E��S���#V���vC�C��R��!ꏨ��cjO����7g�;�\�y�"ѕ<UM���B�W�>���w������3��v��Gؠ���W�,i�,�𧯝��+��[�����ʊW+�rf%Ysd(�z���t�5T%�IZu��;Z��-�ևI)���{e���nwB��d�0��q廤-�i�o�6𹫊���9�t�b��v��B5:S�b���^�X&e
:��tNp|�ϔ!Ἴ�o7��{�^`<����
Lu��qTB��έ䷽a$�b�u��ҧ1�骮��$�]v�O�~��!�66"�s)yS��{w�ڴ����[�*�}�䳲���cOU�g2�j�dm�\�0+�G�O�!&�Y �
-qX�j���3F���:losK��j�+��c�W���Xh����³^�I�������SO'��ʅڔ�A�I-�"�dS쌆p��]�sZe��|F�v�QJU^���^i3��=ϓWg^_������o��
<J���[�����0f3��)KR���w�AN's=���eĲ�X*�R#pͶ.Y��\X�w2:ɫ��+҂�����i拝�汭��x^�mo�=�~�Hb͛�}�A�&`�F��>���l찝�F0�o��Ӻ���a����|7�+
{ƻ֎m~�l��y܊�@4��MZ����Y!�/�o7즣�1ڻ�v5S��5���$��
�V2��+�����9gM����f��[�[J������<��\q�V���VXB�c�br7��v��X�i��Ӄ����$A�Ec�nL��[{�j5ݸ�I�a���۪�T8VF.Gz�aG\T��3o�}R�Gr���S;x<u���e���lRB��,8I�b����w.�f��Q��-]�2܅hX��5��҉6�M=VK�A�]7��Ӿ{����+��v�s�w�'�;j�;Gq��:����c11��.6�]L���ٹ��#5�d�3��䌑��p<�w���}䮻vw��|�(�
Q!uOV�wj�n�Z���4�����0޺��[c�n���[c ��l=�m�1��Ϋ�%_IU���5Tշ�=̱�12μ�3�^��V�h!
���w[&nKո�����r��]�U-�uRmc[Y$;������11���؋/|�����du1KeDzu�a�q�G��m���۞�RA�cɏv͕��)I󜻯f6����tp{���Vu�3��B�+9���e�T�]���Lޒ��K�4�'D-N�Nu�x���
��*��ZB'.���V��=�����v[ǂ�|�S`l�kC�P96Ԇ�Xj�X��WpgK�κ$����1�f�0_Gu��+��Z�{i����#R�������S�q+Sz]!7�tL�B0�7b6p�o
D�֧�MQ4rn3oLX�3]ȵ�1:�Xk�9�wMF������Â�-)��J~��Gm������9�!�Xp%j���9<�"��Z�7���؁V��Ҋ5@�z�u��8l���X�)Ż�Y��D��7*�qkv�mVX.'�N�.��ww��P����+d}��N���E��7k��Pk��<[ەJ���7��S�屾k���"�-b�v;�sr�p���JYou�Ðc-�NA]�ZoSS]e9ە�3As���m�}�Ĝ�\��UZ�c�7o{2�xũ�w\�^h�ɰ��v�J�V6m�2�:�HF�8v����16N-H@��b��1*R�]��]
���s�[s`����b�U�mc��0a��R�˃���h�l^b�;6e�7f�Xf��R�a��3;v^�ĭ���P�λ�QJ�]Ubd�2[�[G�1�9��Q.��ƯR)e�8�=��^>&���[ę�l�3x�0�75%�:�ʹ(InD����;�R�����Rv�ա.Շ�U׫x�Ji���T]����WF��]���<����{36���fJ�rKd�ԙ�lg_f@�D��/�����C��ۻ���>���T����\[��z୼���m�7 ]l�jJ�HL��t)dT������J�x+,O��9&d��#��{�@NND�E8�G��D��4ӷn>>��۷n�_�߾����I�9�N�"���� 6�̷��D�d		@�P�i�ׯ�\v�۷o�]�z��H5
$����*W�Iq��bs��#���dttkb�)۾�ﾻǮ;v�۷׮޽p0��R��ŨQ>]�^�Rݫ�9Ns��^'9 ��D��4��ׯ�ݻv�۷��z��%SK���K��qD@'S�]���k���+m�vZD���{�|�ޜ�LE'bt6�q�m�!8M��>;s��� ��S���Y�kq˒�.q�s���َ|�XI�`��������.S�դڶ�wH�D��V�t��j�I�.��mօAe��~����襷iiP�kD��(��;���^n��H>'��H�}���Q���^��p�Ym*�[{w��4�d[�	����6�Y�Ȧ�B��Uf�
�to<�5ݰ��6N{���r��6{��C36�����g$�<�QUA���Ս. �Ka���@�W��Ѩ�n8�œj��~ޔ�����zx��h�lǍ�w��e����7�I��b>y�4tT� ���*��Pir��mO��^�R-\il��[q�ym_��Y��c��^}�"8��kV���PK����][t�.���:�C<dd�.����3����yl����V%'���g���{�IrO��9�"q�).���g�a�b|��oK�����a�O�.�j�n��l.�Xr�����F�p>o3�P���Ţ/�/��@�k���c�7��Ի9���\
;�<B�
c��=�,'����C�4�m����]��(�YL������ǖ��nOP�7���� m�[�Ӫ?qQ5~�磻v��
4#c�_��h�cՁ]�L��c���+p���. z���WS�\�<��y�N��V�.�a�]���ӛ�WgT"�Q\����7+{�]�#,`���R���GZ[h��F�/6KB5X����
��W��j�n�I�Ggq�����j@���
��wR���c1{�3���W+�7������c�&zA .����%5IG� �m����R�2l��h齺�#�}������h�(}��P����]?GRa�����ꗷ�q���^;aY������uH� �lA>�h^3F���6)��۪���i/q}{�{��+2h�TwM�y4lxS�èEz8V����/.I%�{h5<ڊ�^�~���g}���pI)8��m��麦��Q�N��qn�Ł��vTpQ[�+�#Зg��]c�L��}�SrK�.�:'�6/�J��"�������[A�w�TB�李Di����^lH�5-��!�>�Ύ�+���DdH�s|�"�J}^��Q@��E4i�IxE�-�P��J�[Yv_��r�?�2'�s@y2Wz�x���W�l����i��UV�*���n�W���|�8^HpA��W�����_8:��� �h��f&����5J�>��M].�?�~��V��ԁ���	x
��_^[���MY�g�"��Ғ�����(%�M/|}�r�S��}�g1(r�2�֘�y���5v�xp�|Ok�0ef�TQP�-�������3y^�T#�#�07�9�o�1��+��g5WԻ�oB�Za���v�n��b,bRMљVa��t�UK�L�~�7�Y�/�diՔ8�Re=�K�������7;~/3e�s������l�3T����u1�u]��d���$u��Z-�)�7gakGd{��9���E��J
p' oA�Ď��m8�An�n]�-#�n�?xױ�p\-c��B*ѡ��8�f�g�wm���^�}�Y	D��=����6E��ܻ�y�5� �{��ޱ7�F�c=`�uK���q��5mwlhiz/Vu�}{VC?��aE��7�^��SZ�F�v52a�bo��cb���%i�� \әٿ?c�&cH#'��u�5�M��u �G,�V�ʽiJ���N���|��ZZ��u�����.b2& ����aoX�-�Nko]��t�B�^>d�߮'��a~���Q�xn^D���}㮩W!5�tq-����S����D˽���층�޾�~�,Q�rU�W��o������g}�>���J���*r����z��ԒV�U.�}C$U���OU�ϴ�S��{����0�9�7vĭ�/$��:��	�:ˍ��[�����O�������4��z�@> �W��c'�U|��o�>}앎�r}j@���")�^~_O`'�_��/�QO�����4��sɛ[��]0��A.)�/
���L�1�Cp�
:��N����kI&F��(���Ϛ��_�q"=f��A[@���@ �d���%cR5\Ry�,�wd]&�K���A4�#{���sܐq���1;���἖�H��K�a�i��k��h�:�-�}�H�w��:|G[02��jڑ�|��m����m$
�b0���K��]a�3��s:ÞǑ\
-}F�,*z��lEt,~�ׇQ=��g��v��C�#�0#�YgInc�� �ì��2���Ԥby�pI��}��e��������m��*Mk�׾�N]Yǐ.]�g���n�s�Ex�<Uѝ�}߹�����M}�
�`]�%��1��9�f��ui$2�0�lE��:ثO��ma�a0�,fi@�j�2q��qڛc��5]s���م���D����zlx�u��y&��⪫�i��n�c��yk�8W�n*[ά�4vj鴗��������1�h�=��Z�)T�X��h5Vk��R�!���{Z_����Mj��uc������2���D轭`	�t��#x�HWCJ
�c�U�m{��=��������/�����J>A ��#�`�ye)(6�hƎ���=��1nF��zU
V�mu^���Ux� �����L�����wTɞ��Y��o�G;ĸw��2F�o?����I+��ځ�N�mx�9,�IC���O����Ȩ[z�7�%c�q��W�v�Vٻy�e��~��֍���'U��Ǫ�'��r+�.I�}k[2*A�y�h9�n�nw=76�&��2���D?��kP5�^k�17u=���D��<F��BuB�[�%lmU�|���Uj�2eΚ����d��C�a��V��iJ�U9;L�q�`Flx��pR���(a]�ڬ�Rv$���H�~5�{a,J�[P����V�mc#��]���IN�B�*ӗ��])�t�
�3FΩ�_��7�\rD�������"��f�d�]{��*��W�u�vc��[�u���sW\�@�}��y��o7��ow$�>7���w�#��>|�u"*�-_B������|���6���ۙ�A�ۉW��wSP8ݓǎ��Hc�j1q=��n�sj0�zƅ8g�څ�м^g�,ڱνa8^��D�E�N(��ꝿv�iE�su�x�f
e��<�5|�u�#R��ݣك#�d��ip([k2{�J�o~5����B���県�W�j���ݮ��S�[�9q��A�Y��M��&uS���`��$�Q�G�{q*�=�_�K�e��ē��&G7�}��<�&��ڪ'��C~�l���R���k�7o��q��bNm���tVr2�ɯ�Tv�}�OL*�R>]]�������T���	Wm����^Ij�f<i���=K��2/x����[�I����^��7�pl�WO����"+�k�OٮJZ�C��б�*�x�cf�WU����:�[�Om�[��i�DP��*��}puU�Uk8#�MNJ��*�뻻8hUՎ�ݏ<@� ��5���Bܺ^[��I��:dNmՖָ�ޠ�Kf�����U�})G�j���ne�*���Mo<�1��1�`���{�/���sf�r��̒�Im`�٥G�x���۪��+T ��s��2�W -���>�	���{�X�E[��h1����+���í.���X<�+f^>c�}+{�%���Y=
��3���vw<�h݇�'�����
�ϫf��n�4�G\�"�;f,�a�"�xV��miy-�V���pLx�8V�ʏnk0"]W���ӂ�a���>�"�-�>�>}ޑ��P��J�,�������#�{4x��CG����f[^�^A�g9���-#�u-�s�GleP��8�����`,��$<2=�<Sxgl)�����#�aY�5_vg�?u��vAO�Y��Ћ���;R�L131U�&�o7n� ����Vi�D���y'�-��.p��w���L8��zp�}w̃�u�u)�?��Ej�q����<����(v��D��J�5\g)�ߡ�7��K.U�ϵ��N&��C�iwyS�M��|��Y��Y�򌙵Ĭ�n��f����8�(9M���`��׋�n��^�%������uV8Ԓ	��B�[N��8WY{\��c�1����vo�_�{�wX�ҋ��}�v�{Ϳr��Y��u�h���6����U�wF���|è�H�2�
��DZ� �C�}fS���3�&d�]i�]�����5 ��<�J����Б�7�oO�Y��-V�J��:�:ڣ�L�8���d��=�gu����ܜ-96�~G9M.���<O��냔�:�����/�gϠ��uu���-o�7<æ25R~]ϼ������\ZY����i��s�!Xwpi�/;�33�4£6�O4V�y��-V�Fy¿��Q�W��F�"3W�Rw��A�Cy߷�i�N���+�Iݐmd�(�ժN��YD3m�3��&Lw��*�P�[O���w7�{��=�����"�����Yf�>Ͷp��'J�ĺS��x����;;23/+#,�OsRzႩ
5:܌VVD��p	p��H�W�!��ݶL���p����b���ݚ˥kp��v����Y���G�E�x��5��z�NWj�X6���$�6��н��i�h��n��T��b�U��-4�y�&n	.r�˹̶�n����]z5}��\�EO=��6���ϕ4TJ��;��C�%��
F㳛���J.;���V��}���{�}ǣǤ�^�gC�0+���[�x��)��ݺ�#�ȱo��S�L�;}ō���M��Ϣ�oa��ˬ|��P�!�֊G=l/-���c�¾�rX`�/)#���ڽ�';zȭ3A�����c]H�T���	���g/��m QJOL������O	��r�79M���A=a�B��v�+J��z#mMVMb^������rk|�=��[���a� �wE�tS��l:�����=���j���JeFI;y>�oDӻ
cSF�>���6I�=-W���Bwc�ּ\Q�QTEmi�ܟX-[��A�=������u����V�oBJ��m��:��z�x0OĄ>̆���nt�/b�8tEhڜ�a�i2WjPN꫃_f��U|��}�;.�,'S�^􋧫�Y������4WNqVv��en�3*����@��v�۬T����!��/$a�Y������;s{S�]��Z��p�Z�2�a��!�Ww{:f���ȫ����pا3����P�+��PtV��l�&;u(2���K��aoђ��y���\��׏�fY�+��ڗE��+�5#��q_�\ś-��{a�yt��>���R��h������U�,�'�u<䛾ԝ�{dl���3ip�o;<����یB�=������4<p́�ָ�в�F���f%�o������(�Y�e�+�Hm7l�3��^���7���nT�ޔ��ً�*���W���!�'$����I�5���oN ټmS�"���F0��ѻ^�Z/�Hb���(�'����.)$����^MnU��Y�� ��ݑ����.���(Ǟ����>���p;��]�,n� ���5}��'��:���R�WN�y�������_�U#��@Z�PPG���� � (�#���h�@`yj�R�A��*�N9uӎ�]ҹ�s�.U�1	�@b�FA�V�
D"��dF(.NNs�\㓎wu�.Nr$A�� 1	��d�wJ�98��]N���K��wU9�N9ur��u��S�W98�WN8�wt�����s�wJ㋓�W9�]s�Ur�]t��Ww+�\���N\㎂�dB"� �a(EK�wu:�s��K�9WJ�$B �d�@b#�$(��@`@b��$"��$*D F
�@b!�$�� 	T�)�$�
@`)�$��@
@b��� ���`	�$(�
@`��Z�0#���4@�b(�`�"�`��#��������(�^��ب" @n�@("��������"t�B �� 
� �� 
� ��hB���������(� �T�H ������*����  ���"�@`��� ��(@`)�*d�U#P�D$b��� �d�@`	��dB �
@b	�h@� �D$`)��*�@`A�$BF�H��FA���dB*���b),�@`)�"��D �(��y���Q���ª�F"$����bϿ��~���c?�������V������ ~����@H��Z?���Z�����������@_��A����?�QTE�Q a �O�?�| � R�O�/�O���~�?�� ��?��?`��s�_������A9`W�����(��`���	A �D �"�$D"�R @B$"0�A �R
DB$T""@R��B(��A#H(@BH"@H$"���"�B �Q �@R0D��S��:�U:�J�:�] I	HT$Q$ EAP�I	 HYD$� �TA@d$�躢����!I IIDA$#E$$Q����*�J�\��*�!H$D#H���D�~a	C�O�G���

Ƞ"� �H (�}��k��_���� |�����~�@Zփ���/���8_�>%��4a����B��Y�>��
���Oˮ��� @~�W�!��x�>��@Q�����  �� ��(?�������r��_<O��#����
��z������� ���@7�o��o�~{�}����?���Ɓ@_���%W����6���?�y����	A��e�?/�����M�(�
�'�$��Ґ?�X��h?����?�ߋ��D_�|`P}�,QTE����=�x���!�'��(+$�k#O�@���0
 ��d��HG>{��]�HJ�����m��Tr��J�5(���+f�SUT�JP)+���$ �)iQ��ö-]u�P�Cm:��M��c�f�v�v�7eʒַNm5��gN⛋p��ugk��k]�fӛ����鵶�m֗;�w��W��nwR�t])�;����6-��Z�n�u����]j�:����ݧv;U����˳5ηh��tn���*V����k���*m��uۊ��.��ws��k��V9�sk[vW3]��l�-8��:�7wh��\뻭�ݷo�  M��=v�[jYN�)ʚ�m�Kz��H�ݩZ�m֦���ZC�R��M�g]kt&��7�ݽmi�J��ux��i��[G��R���I����f���u*w��f�[�Q˷n�skk�����g|   �X�(H�"}�
}{��T��+Lm�$,u}��W���T(P�9��y��۵�X�Y�U��k�S��K*ڭ�r��H��mZǷ{�p��4��N��jR�MW��u[��Uh�v]k�nw{��{Z�vۭS�×  ��t�����o�vm�J�[:����sVU�]�׶���mM[���4�(�{���ͬ����o9�픫m��+ݶӭ�ѫo�z�6kU���]��U!ֻ�y���͝�;�ݫR۷n�v��ξ  ����5UU��Ukg���N��o�^���ѫ�Xtڊ��À�{���vB���k�������W�`m��wS����u��ݲ�g;v�6%�T�v�u��  ���Uɭ�m���
y��U�z�gOi�����v��{ݵ{�[j=;]]Q�1�n�B�{�yh�UuF����p:�xk������{�t;��.�Mλ��v���o� i���
���׽P�tl��{�����۲ٴS[�vj�5uzު{�׽��S�p��u�J=��gz��:QZ�@4��;��m�n�ܹs.�ڜ�[]ښo�  �_  ([|� (N��{�h ��� �8� )Aev� =s��F�����=�`  =��ƨ({�w6�kwW[uv�-fi�4n�ho�  g�� >|w@ ڹ��� �:�

huk�;�
 .s8ZP���p u��`����� .�p+v9^�*^˹�k;�6�u�k�]ٮ]�5]�  ��@ �}x  ���  6�P q���  =�m�A���x N�OU�S� k�V���  ����]��n2Z��n�����   w��Jh����zP��{�  �o^  �\]�P)�x��  �q� :���]@;t�P ���t �"��M��J�� E=�	)*��h�A�{)�j���1# #S�A)*P&�F*J�� �$�JE1�T�  3S��1�������9��I7?[쇼:{y����/`�Pދ�`�$�B������}�;�Vֵ���UU���kZ��Vֵ���[Z�٭UU�����_}�x�?�F����!Q��ŕ�nK��X��t����� 2�����Y�L:U���H[D�OQqIn;�VHVBs��4E����G4Xd^��HaKm��ZQTŀ+F��Ă������b��Nꩰ��iݷX	�+0ּ���*�j�1����8ޛ�5k`5�#�Q[��Ʋ���6�� r�����Җd7B9n��y�p�"�<�2JX�ŲT�mX7Ke)����)3�Z�I���Jט��{!On��[�H�u=Fڲ�S`k��ɼ�0�KVUܦ�����ثx�:��]e�pj.Q؀Iށ��pк0Od�$0&�ǃ~�#<�b�t�"�����ۚ��q��nRFě�+[A^[�����&'eǴ��%;�j�B�Xtο��U���Ǥ���$���*�L0Z�t4kCk�,S���v�I1,�!'�Zv�q�(�P:$4��j�-0���Ard٪З�fӖ�AĞ���Ź`ZV D� ���'a�2�Z{%
­=ж,�uiVD��Lb���<9Nl%��f��*�$v��V| +
�`[á=3�y�AB������ô�4�IZ,���Pc�ƫr(��C]mYWXv(�Yy]*l"H 	^�TeDX&fg�3+f^�N��2jA!�X�)b6�i�R��@�n���p3pҟ;�׊��嵆n컬1�Q�Uw�LR�� 5k�h6,X�@:��wP-���pG���V�C2a80A�؎=��B� ��6�)֫_�ʺ��t.Ӧo^a*=��1�P��(Ӕ��]&�m+����6���Y2�K�,֝YAe��,�#/������=���T�'Z�0	�j�sN�L̔��f��Cv���zU�0J�VSͥt���Y�e�eB�f�{ug,,y6K�6m�G5$@�S,톫5aVE�u���yJ�NX����U�ȣ��Q�"|���[�n�@����}2�ZCLMz�E�ֱJy��q2��Yr�ڈJ����+-e�括�`��NB|B0�nk�Y��Z�i�I�@�fh*�u��1Gi��-(m+�����Ru��X��+
��©��l�h��w#q�Ȝz	�E�3��o܄���e|�N�c�6𛷵���b�Gk>�d�n;f��"m}���b��h�����M�z�����tj�H��Kb����X�f��V8�9D��yu���B���_4W#�M0�Л�z�6�AaXaP(�v��2��Z��M-�z�P9F=H�Z���#
�9R5���tI$*�".9�E�Ǐkbi�wX�:�U�^]��>ZR���Y^CGw6��I�Gm�7Wי@^M�#���ф�%�lmc�vѷ��z�Qv�+2�MMT�m�y���,��[��p*�&<�T�ɔ�;�FθDU�40C��4��0����:��d��� /e;#A@V��⺰�+�mU���7��Hbö ����k3+�0X��ʺ�� ����x���L��w׵Z��
��uwn�yG�V]�Mb#���nT`6
:���B�����)͹���{�!�/d��`���GH�0[I�����A�ӦM(�wT������n֙��A�x�՗S,�y@Z&M��P�0��u�L\N��.����M;z���f�y�*�;p�fnR0�B�Z�~ͷ��Q�tv�x\�6���`���5y�< i\�yk�ل��	���[�rb-+���*�\�@SB��x��ucY��n�8�S�\�h��`q���4e��9�lM����y��;ܜ��:#�9�"gd��O%� �$�4lO��`:|=3�bȈ S��nshјҙ���&�v��ͤ/ij���(S���ѩ&h����Me=��^�õ��������F���S�Xk6�"�Sl[r�p'HD�OJ�;��Á�/6�*�7zF]�J����TI'7f���S�YMRӹ����d�6���hJ���!�V��2�&��rMx�M������l�.Z���r����-T�*�g �w�ȼ׹x���hf�G[s	;۠����bfk�p<ӭ+*�M����,U�f�e;���o4ս��H�Uv��S��%��)Vx7^÷���qP1�V��6�A��h��m5Oq;�){X��Lt�-Lb+���JbDc�|i�l���\��a�#-�f�֚Ԓ�X^�z�Ǧ�h�L ���򦶯i`]�Bۄ��l7b���p5�j��e,��{A^ݩ�,״���j�,eV��. �j�ܺ4Pv�#r�4�RMsY�́����&NTB����i!XmU�^��cF�&�-�Cؾ�ԫ
���b��gs�j��K2a��i�5E+M޸�$sM��r�X��	��Բ�کX�Gd�Ź�嬭�Led,ֺ��.��j+����Z���]������La�Nf儱S��]-P�dnU�ރ��nԣ1�W��(�\n�!Y��{g-2�7�f�N��XV���~2⚰j���#�r^a�mȯ����k5σ�bhR���Ye� �Y:r�*��qXW�v��Z�f�V�Z�� �w3sf=�Ԇ[ GRV�)7x6\)�����̝0�lLǷI	���"u����N�h\ݻW�Y���b��4�X��b�ܙ�k�]d9���!"�X8�SW�$��*�[ܡ�V-�[Q&���kT-	C�^+�`���P�F��Jd -�J��3twF�˛�$b���hl�OU��ɑ�`%F֖��6�,�e�1� FÂ2F^�U�cIb+1Z�ݵnQ�3>@���ء�+MW��
�'Y�]�� B�3.P��m=Y��ڷ��C�&H40PH���[��Aڔ&j�1��v�1���!Ͳ 3kU�w�yIcQ��iMc5ˤ���� ���처T��k��b�۶owaiL\��T3�ĕ�%V�v�w]+����ncג�7�hOR�������]D�OX�)�
����4uD��9+0n��$�tR��nʱ�H�)q�F��R���Tf%<R
�+/Dj����fm�х�ʭk�$.�A
�>M��3�N�"�h�+%�cB"TI��.��rL�	n�c֛C�Ѻ�T�4ñ��2ғU�� �Ҟ��0Z��شK���rhǧ��iS������8٘�0Ei�U�R�c�#W��;���Sǲ��w�i]lX��UݨͭH f������/4��e"w ��-;Z��8ٛKYch��ޣb�e��DJ��E����8�8����{R�\��qn���E��Y�;��[�i����]�7�魺[J�ța�&�Uڛyy�)�H�%�'Fk~�H�y$͌e��H�)�����T�;�YR��w`�
{��o����L
�d��a��8�d�t0�6�b��qD<v���N�FE���#�	��];��$�MX�Wh�YLe
�3`f<�0�r����j�m&vbY��m �����{e�U�E�F-r�؄��9�mR�$��)sw+i�����	�ܱ�3xY��rB����Q�ȝf\ɥTV3_�qǚ��2�L�(З�ȫ�L�H����f�1�I'� ��q��9�L�����W ��[bK���ť>!q�DA�OEW���a"g�0	R��j��5B��8���{�6����n���n!��y�O�6r�D�L;�S�-k�eԼF�g�1�`��@.�	"q��e[L/�1�^0��+ ӊk�ް��L�6e�6����ҪR�C�lCe�܉���"emetSݬ�Zhb4D �Fݗ�v�὏�ؔ�B�����d(�aG3 ���w�n�N��������`�,��8��F��-ѽ�`���!W2�8�xs&���WڕoS:�t2�˴�db��r���H7�&PHe:��OT�CQ���Zͱ��Z+#���l)���(��1�*�#U�D+7vJT�R�/cl��7C��`S�n�#�dʗ�G[ܤc��{�\�J�f�SF5�(�&Si��t���Ǩ݋M�*��NY{��%�MM�����CNՆ�Tm�ۢo�ݖ�"{�3��$ �n�ް�8e�v�4���1�6`W��@������V!�w$k`up
eEN�`W{��ܩ��s��e�{Knz�ݨ�jY��x���f��0���8�j��	V¬V�ԑ�h�m��Cߔ[�m�����t��ͣ&/�K-VC�����rDӚ���G/4�ے�5�m�]�0C6W{bd	�re�n�ŕy�R�H��\z��O�$�ۀ^�b,��2����A��na��A����c+r��!��Z�;�+l��ot�b�0��sT�ǆX��Ahv"�B:Bɒ�€ܩg��ǈ�M!Ǵ����H�%��S�R{�� 6�eJb�6��2������P�
�-<*M�2d��V�8�^C�֦bof��Q��܍Ġ3.JE�'mMˠ����J�5�?��
�Ńct�H,m�5��2�*��f1RYlE�H��^6�T�F-{$�h܏Y��kǡ�v�w�v����vh��x���E�Xo�;u� �͗�+�v�՗����"��ld4J�5���*�ݽ��{��D/"�#�"5k�w��:c㔞����/C���d���&AV���A8��KMHQ{�#���=��xC˽�"�{�6m�p�l�ȺWA�1�nGr�2��ө���Q�R���*ms7�@.Ц�lf��n�L$=2�o��-+!ummӺYM��#Gn]��h��&`̕p� g/��,RXac�R�fRe?��{4&k{I:�"&ue�{�31+��<u��a���ҫ$�艻�/p�n�����R,M&�前�Y
��T��)q�m��Q��b�Mò�k��2άJc�3�t��H���.��A�u��B��h#��ڳ Y�D=��B�L
�A`�ܦ���ڹH�k����M��AY�"kB�f����S	���-�#-�q�,T��V�jV:U-n��2ؐ�v3[m�X�~%&��Jań^�H�X�w��ն���V-���-����T���F
�;(�g/��F21�th���U ��l�)i�RR��m��hu���.^ԧ%��%w��$���u�o���ţ�y�ŚY#��wrװ��D��.�~i ]�H����=�Ā��-i��6{�WC6��;B�)^�%ZR;�44[O����72Bn��q�̧���N^V��ٽ�ow"j��HGFJ��c.�C���u��YS�,X�:n(��EB�-�V݂���g��S��dc ���,c�>i�lح�bc�hffekxBuj"Y��7FXZU�R�*k0;N$R��VV�ٚ6�m����t�j�Xëw����4VK�h$m�Ѐ��I�a]�d�����XvtT�Tݬ�$���f��2�D�3'$�g#���B ��S"Ɍ;�\���O\�<1;/2G^��	�����*�@&��l�7Rt�X��mӺQ&�ͣ�V:�p��-�"���[��8X���,�xB't�!}�r�;=��A+�sQ�H&��l� ,�.L��N
��A�IzaV�FS(1�/l
m+�b��T������-�yWJY�R4��ݽ�ES�J=�Zu��\rH�U��X�P�����!��L�֕Z��i�1Vt=��� JU{PB��K^��e ����,L#���s��;��ڻ"ٰ0�+��F/E=�l�D�M�w̭n��l{���A�b�r�e'%��u�6V*��Ux赹�7c7��nS"���m%�66�胩A%��v��	��Mf�8f,m_��ZA��Ghp�Y�Ʃ̇�Ṅ��2xf�e �h��me��K�c��nVnK�Vf�����e���ɦ�EF
�Z-U�CE�iJ����yn��H��Kh!f5X�bSf�Z\�׉��N��""���\Soq�o+�<�RӋ�">P����]�/RJL*��e�Ŵ�]��^�ajN��
�,��ޣ�sAv�e��Um�J�+n��5�`�w��v���MES9c1��ڒ��X(� ����sl�0��-S���-g�w&��&o���۳MǸY�֫��rAi� ��I@앖"�h/����ʲv�4+-0�^�A���l:z)�� �^�*è��(X�j�38�;�c݌i���(<�p��k��oQ�T�l���q�\t�]4�)��h�X�3R�4Yv�v�,ml��;V4
{���N6se�Ad�7v��4��.�㛘�2�;�y��M Q6īҦ�)�'cnu���د$�WB+�5�m��k1�A֟��w�n:ԙh;-b8",����`�6�w��k͊,�K�����)��Mܡ�E�B=��9�c��o-���Y�@/�Đ�[2݋�C^GFd�o�m0�a;	�O�c"�b��ym��)[��KK����{m��e�U��ѣZs�n��{��*J��]��A�{�@y��;T��LQ[;���(�5w��do(�����<r'Yf��׊�cC.���)��RJLvl���Dh�K�me=h`j��h��.���Q�v�V��P4.nF�M����chK&:V�,�u���#BԆ�+�!VF�P���Zò%��WƱb�.���9���hS��/xy둼/�/F1W/�D�ոv�G���*b� �E�M�҅`��ڡ�[�ȵ��n�o6Q�t�?[I5�'9�c�1� UF�j�ǻt-ԫҶ�?�m���nS�������\�='۷i3��G7�K%U؈��YvK��=+���ݽ�Of���5x��L+nb���`+��c��L奅�ŰN�����O��)���Sy���:M�`�/y��̮����� 8�k���`�L����%�q�D
X\���}IC��ǩ� G�gs�#���ގ [�r�;hV{��뇑��qy�#�+iJ^����G1�v�Ɩ�C�z:Ï�t����2�^"��3�=�[�}HVW�U;/���ܹ/�.�\w�j�ԩ��΀��95��,�G8��=�����.�L�s�h��ۼ�U�u��V�8��j=|.�Jh�/x��&J��y�����7{pX�j�Y���ӻN1L-"�+��9�|U�i6�DÏ��������,�M=��g�v��>�C5�bw��$�,)z��L�L��`1����� l>�o���'1D�z��779�=�#�q_GS�s��)c�˛]�[���x�3���E(����+h��X��hdo'(�d�_o.'�ҽ7ݘzV�� �%fuVU��?��0]gY��B�S9C۱p9��a�`��}���c�Aū>�ɘl�Y�����묶��;r���S�6�5P�,L�T�`�w/_��s�][�n�T֕�!֒7!~�
��`�bs��w\O5��44����e��k�:�,F�Q0�s�����fi��Eo�N�ָrl�K�C^���<�N��w\U��C3l	��'���|2�<��0p'n%;TI��Mދd2����ч���;�B��W�c7:_��l�^�[�@�����X/�`N��R�s���i�\��w�����25�d�t��b�>lh�-+��_N��ŮG�O�B�j���i�$��x�_mі�P�7k��̆���dC�Y�I���΍��	���D�:�F�^�`6��^9�vk���Kgt]������3wB�u��g���&g+M�=+4��NqͲ�v�k��;c;
J��W�����X8��R��0w*�	ԡ�/Fc7�(ĕ����h$P/W�R�������+x.D>j��t;6u�ٜ�����+�)�p��$��W�T�M��~ �(G��������M�j������F��3/�(�j�ʛ�ڢ�����+W;��鋢��<Y�䕲�f��5��įl�mlu��+���#��m�v[���r�t��c����M:��ɂb��V
��ą:q��M���T+*�_0wMͬ��g�������[]n_� $�L�$�i��F�Z�B�ХB]����c^v�,$Pm�`M�Kvh�g��iX���;h����ܡL�sZbd��+\hx��o*i���#b�;���R#���Ҍ��0)�u(nU�/m��
:���$:��tq�zZ��h'�-��Z��]޽wfpI���t�ŗ��#oV^$nm���cc�l��H��@^>hSF� ��zl3V}Ɗ����+F�N�ˮ2�O�%5����+���䃷1!{X�L�NC6���zA�r���PVu����ń�����/m{��	Z�AH\w=޻C\I��x5��:��+�j�Y�:]�6�WI�Wy:��%b���jOW��ҳ���e4��N���2Hhv6v����S8N'm�6r;u�([��1��uo-*�B��8� ̕�G�@�[ON iAB�So���:�I�b;�yΫM��8���� &���s���jk��Ib�m��rk�JX����Rګ2�on�M��J@������R�0Z���b&���ܚj�l�]��+U3�[豑�(|����Ҙ"�;Z>s&K$w#,fV�ۀ��e���sDJc���jJ	�3��B�gaƴ@1�WR͖MSȣ(\O�$��nw���=�^���6�K��o�G��i����̙H���`|yV�4���,��ZxNy�JfL)��gq���P_9�m=��؊�9,r���B�O/:g��:X���ܐ���ư�lF�Ҋ���2ި��LC�3����j�p�V���[N���a�Y�YW��ݱ�FP�C�����s3z�-IY97U�j�B]�w;��h3m5�U��,�s	~�9�vٳV�iwF��a	�[	��N���fZ;�JcU��"�Q��g:7&[���9/T�}��a�2���2q�0��J��ԡ�c�(B��j}&���g��$X��ƙ�D�gKj��}r���/7P�p:23FL��_Lb�p֬����c�.�SVkK�{�[c��搤H�qu@�����h��M@�2Ͳ9�푻�b�m��8H"^�\�=�!(ɝs3�����@zΆ'`@�����f�;�
�o,g:��5m��)��r�K�����Ǻ4i��Vk1�Yn؍����Z \�L�ְj�ck ��]��v$/Ƭ��f�d����OY��V$�vv	E���K�=([��1��F��)��Úb�Q!��&���9�2y����O0��Gjpٻ���v2^ʁ���9�֘RwU�ww*`� �+��,q��R�xfRggNVU��f.���ƪ9$��OC�9�&�Ԕ7/�"�%��&s�x�ƳJ���fe��yOq)��Sa��0����X�(t8�J8g\ i�r-���)��n��>ň�M�;~��6������6R�<�Mr܍���d1��p!u��#�qڭظ�R�9ϳ��f�m;`�K�-ɨr��,֮譄�!��r�T��WV�gPl�Pʨ�.aD^мX��i��9�Ӳݍm�\�ܨ |E��l����t�5K�E��{ېZ!���ҜxK�/jո]��J��"�s�����Q�2�NЛ{`Vq�':�;���\�3j����չ��( �R�f���(o��/��3Nn.p�K}��%4�d�^zud܆2��Q�j�R� �������0�.��S��\��ob:�i���A*�[
,��9�.����E��64,ķ
��U�:���f���\�Y�|]GCI�!�9�3���{/��[��[x��7�:���rD�Ք2����[���6���̰F�>}��-��1h�匃�r��],���do+|��r� �D嗀�Q�ڵ|K�����ҥ--_`g�1�����<��b0=|V�����೭T�TI�=��̥<}�"�Ķ�e�n�y��nɌ��y7v�<��h[�ʮ�,kV���J��ml�&��]-򎝮�>�r�%#�m�j��YZp�4��j�K�r��:�Z�%]�$y8k���M��V�0�����v��B����b�.�˽u��ϩlu�1���O����
g�!�$���ۡCb�Ut������`��k7��m�(#�m!i�o��qPnE����z��7s*[�]�h�m�V�Ť�÷�0(�
Jju4�ڡ%7����S���:�F/�գ%ޅ�1��!b�ݹ��FE�-y|����EaGT6���"���3N����c.��;��i�t����i��q_���l���o1���K�[�v:�o��`�^�)�RP:�����!|�`�Q�8ĵ}��-���M��p�7v��p]*�%.tA���gm�Ʈ0���ӡ�wYt�p\ �:X����,]�U2�,��j��,!4�,z����#�fVj����[��J_p��j��2���>�e�Ke��k�|���L�w�q����h���mv��5)�]}Xfek`��7Y'k�����f��+N
��50����⢓�R���f��z�E�_��ݒf�9�����^�yǚ�b���QY{���!�͙�0{��ͨ�Mpyڅ%d���CIU��Gû��#עvZ��K
X��m�V��t��\7��%C������n�&x���bb�8��u v%��`�9{o8V��M&SR^�oc���G��Y�:;[����2�27;+�**�Jȵ���L��)��j�o��g��q&9L�)��ňZ�Q����J�n��� 鏜䟫���$���+(�{�7��+2��<r���K/HE��yw����MʖOڐ9�J�7X��[n���I�����,�0o.�R� 7cK�A�4��ܡM�Ux��v]1A��p�>.bit̧u�b�$�������u,�j�+v�X�-��3���K����W���*v�����R�ŷĕ������v:9���YY�(�kR}�	P��u|E�%�˖���m�G_��
�Y#���.v�=�H�;�������!�|.���v;%�>H>��hvq�;��ep�{��cX��y��r�:�G�N`�X��Ս���4�㻤�hZs3�:�M��f�n�,;d��6�����.��4p�X̬���Ѧ��6���̈́k�=��O$"��^�p�. O.����]��7G�Uґ= :b�us*Ȇ��-��hb�S�aw3)i���@���=Z��� ����#o�S��ɇ+z:�w
��9��.�l���+�-��H�fI*l�6��ma��Vޚm����WOOx�;��4q���˽n�U���X�ͧ����j��q{�s���U`ؓ��u��
 f��$PW��s��T.��)�xU��Cr�ݜ��M\^��;�_gO[�X����b��[���J���b.��Ne��4�i�r�S��	ڊ���1���nf琵����Գ�5��qվ��^��F�qkЮ����z��:�(4DRӆG���s�ܭ�O/���Z�883��+2]�$�P8&���Wg~�%�������àeu��G2��yگ��x���n�fv� �8���{��S�|oXj��7�]�m<��/�v���:��K�\��	{�^��3z>�4�;[��
���-N����"W�1&b���p�����X��ht��F��:��(��Y�a4��I��`�|�Ff�\�bT���uY��b��6Ո�ec�Pajehs�֑���j���W1:(._]%�:�$�7\�:��b�_ oxP�,���E��B��@����b�A�'+6��]��f������q��h�^�X|Wo��B��F�Q�.��n����V��ҋ��v���/:�[�ޘ8B��g4�ˌ7��l�el�W��-��nS��*�Z�	f_K;�����tNB�Xc{�3�N7�f�*�+�&\�;8�[ԕ��t��k	����6����8�E�w>�ңO���$�i��y�f�3W�5�W@�5�o��m�/b��q�Ǖ��5�`X�˃�lZ�xX��s����nQ�#��e�U?1������c-���œ�<��n�.����a�B櫭]��i���[ǅuJ6}�+��xƵLn@�<V}贉ף�V]n |Fe�t�����_`�bk�X�&ّR�b�Yd��$W���$ʻΓ')�hW�^�傲�*�=Axs��䯶v���Ű��p��g&d��:�ə���� �m:p(�֞��E�S�J����w�L�1Ӳ�q�&rv����u��6m�a��=(^�k b�O��|Ms��z0�ždKzy�)&Q�-l�uQp��G]�cd�"�یt ��a��J�	�S7��e4�mƔ�2.{�ԙ�%�[�Lz7{|��c�(�m
V�$m�~�{�A���C!ѻ.�%��U���3)*'g���nC���鮀�44�(�#u��v����������|tR��tU��Ȏ���6K�vV_�#�r.���_��k�ͱ]X1>Ku�Ed�Ⱦm@�i�ۤ����8$��+���C8yY�t���W�ѯ����έ.�}�2�[,+'L����j�i5cL�VU�@�U���sT0�0�oP������/U9�����v7�4�L�`���o0�Κr��lb��j�_R�,N���z�8B�^�<w�]�%!�#7�@`c�^��Թט[���ǤEJ[���4"�:2�r4R�k�[#�>֡ضq�{���e��N�f+��X�c��\���o��GHl#Gk��2����%r�`t�܌�[J�wU�Ee�kGH�5r����i'���"P����]�+�f��w�Y�,�W;-��t��ԨQ(�>���gE�	���l����`��,�:-�w�hY4B{;�JꊃqW�}Ba�(��GR3{�a�/�����g:�dbJvs��3���.����5�Q�3�@���a��%.���Wۚ�l�v#]��{�鵦l5����r�v�ӝ�(L�Ⱥ8��_^�n�a�(.Y|1�`*��=������ۻΫ�����ψqz�fE�7����M|��[WȚv'+٨����;tS� >�����}ȣ1�<)Y�g����W.��b3��hBD5
S���n7�#F���ickw� l�g���Ő9d�篳 �WH��U���W�s#v�QA9�aVlЈ�ӏad25r��1	\7C�����=��!�A(^�������Crj�=��8T�^�sN�tq�C�u��oȑ�����j��۩���	ک��=�n)ݽa�p?�������o�yy�s-�\^IKk�Ւ��J��3,���C\����\��԰�p�a�ɝg�1TP]SA}�u^�Z����n�b��e�m���e�JI�-�j�N�#{��J��K{�j���sr`�:�O�:D�
�=�t�؂� ��e�T�3����ֆ:}�$��ѣWo�3RAyIMC��%�h������(�P�Ļ粔R��I�̩:K"��7������X����Y�ޮ����   ����������¾E~\��l�$�2V��Fc**9�+,��嵻N�\�pM�2,t�����K'�mf �M��-����l�bɎZX!��L�,yW	IaΫ��[Z�6��Ac��vʖ/�h#]r"�Z���ژ�^ݝ��QDU��v���S�S�s,��l�l�C9{����$XJ�X.z�Ee��d�[�]u�e����εB�o��W�m�l:J_EvRγ�|T����jh8��K�f*���r��"_f�,(�m9��{K$F��Z��D�̬]��������n�J�t��6�Oq;�տ�@+j������W]��L�}V�ˑG��X��^h!�X��R��zm�� ��c/]5��.�KF�w����I�n��Z���b3�9(:۝ieXхꞝ���zf%<��ټ��v;j�ꨈ֗�CE�����}27ٽ�[�*�e[z'af�pt)�2�LŜ��R(��1�;��XO�$oR��s	��,�
�|,�-.��`�٣�vl��s�i~�Zڇ��N~� ����᝸���h,�����S�4E{��"��ZY���^^[~M���㱪�tǾ�.+k\�T;�=�VC9m��<(�F�yg>&ܘ�[z5 ��XǏL�Y�0�Îຐ9�W�E3���f�ŉ��v	O��m�����*���D� ��Z��R�{�\�n��E�.��ܥ��j�5ibX������]�h�80Yc���&xR��n��� m���2��e�spm�I𼥿!+n��c^��VLO��d��KŖ�h���O�yr��g�7��}'Z����i]b�C�t���8�q4"R�y�{��S)��C��f˩ˀ��v�7ղQ%��"=����	�&��-Q4���kWd7��33pJA�=Ɛ�Ѻ<�F}��c\�O�M������҆t7&v��vs{�_��H��z�E<J�&��όnybWe_l��!p{$[�+c	�n��+FCp_����;��%�Z��d�%zw����WOs��Y�9�}9��b�i�1[�uAXr�jiVe�H��n�瘾�oX��]�u7AD��G[nx4��R��NH��*�K��r�!���r^e�DsO����H��B�͙�����Aλ��c�I`��T[g���frzf��]�V�|&t;<�e��[`n�mJ�ZL�T�����&�sz�-ÒRW�ٶ�}�EŘ���h�Όn�駌�q���Ȭ|�Y��6vRg��E���6�0��2���uÎ7���%K% �eVE��Rb� 	R0�0���΁�}��'��k�j���Z���xƗ�+��8\y���/�$sჵ�r�w9�V4�f�Aj1KrZ6�9���=�I#�#���u?l[`����(V�����Q̻���5��H	��?^�;iڇ�R�gͻ�U�[;�5����Ǹ$��&��n�U�.��S������Z��`��7��qGϤ9����B�Oi�zv�a���/	����ms�_T:����(�KGtQYPο;v��� ��7s/���{�7c�b�z�����1=Bz����Snh��+Z�ww����r;7lm�WE��R�sy��hv�!�i�\fW�}x�Y�IN ���Zh���y�{j:�bR�Q!:�e���fV�=M�� �U�U,���
<��B����w��M �qlΡYx�e�k�û�S���wl��g��OS�	�hq{)�(k'X�夘+IӅӠ��=g$���.�C�1�8�rNګ_K�v���+b{G,��׭�5ֻ׋e��̍h2�<�:x}�Í��KI8v�J�	%i�f�JE�ʒ!�<�ڢ�0&vP\_m\B��.�Y+��Ր�>���&p���\2��*���h�ub�Bo3�Me�P^�]����t�wթ��o�������	���$���n^�4����xckc�3=J׉����{M��K28'u�33�m�i���Y7q�g���v��11G�A�u�!/�Y���N-d���dʸ_:����7Ӛ8�r�48h�1�D����uk�*挻ǫ�!)eN(�J��6ѕ���M�b�,���ǻ���,�� ���մ�8�n�3Z�J۰�p�'2��TW��@�����B���f�ȏJn�e��`���l�lJ^Q�Fy��V>8ŷ�����x�m���7�G�k-���`�TQKF���R��f�^U`�i�v�����ȾKs�=��"t\ʪ��Xk��B�5�=�y�%��;�bt����SY��n 1���ޣ��q�d�"���y`����OٓAM��%��c�w��ƦMޞ�2B�n!�WG+˷��]��9g�Tch�D�����u,v5c'uf�����e�«D��l��35����)W��Lᛁ�I
�����w����QG��'��U�)V3����|��@>n�g��\��_��b��b�I����]��*�2���͋���k6mo!�S��q)
Dl�`S��:k��Mv]�g��"Ֆ�y7�=�צ��-�����:�1�q��I��+��RV.;L�'Wѕoy'�3�E/��2�g���"�ފM&_bS��Ea۝�H���rbAY�[d֞9� �sCnQ}q�[@i/7�5Sc�;�6-�J�Q<��[���h}	 ˜ü`���t��4�:�\a�e��.�A��;���ޚ�yQ�\����V�v�_G�{u
�1�@˿���x)P�ٰ�:�FP���6���3ݹ�����SO^	���Y��Kpa�&���r�3Υ˶j+��ૈv�ץ�-��h�Ѵi*��n"�w|o ��#�`�K�X�$�̾ek<;�F�i����5y!Wce7~c;���a2���\�y�!���yF��ab�:�:4�[�vz���qxoiZ�\�<,���\��� ��vvW;��Z���.��V�r%;F�*�
��·�Ա6ɝ�ո~y@VTw����Ŭ�ǜ��I�ђ���8_	��K<�53x�D�+M�(� K���ǗC�p��H8��6��ƞ�(hf�y��F�0�^��>�Gv�C��_Ef�ú��0A85����[!�)���ﯰj�m97�����貙y%f�S�Ϯ�n�*� �#�w���<��t�޸��Nc��Rm�Y��ORB(nl�>�������޿A���h{t�ոFf�M�nl�V��)	�\9��`�e�K�V�rnu�J��VM��3�-��ֈ��W�0��ѩV�O�`JK����+�V���.R��Z��263^��5o��olʖ�e�5X5���]�y��I����'�jU0�4�g\�>q���o�Rt�ք��+J��v�b��.Yt���Ǥ�#�v��3��:�ͳ�V�\��\5b���5�*���t�%; ��Z�]�d�]�;�1��A�8پ{OĦ0f��I�=2LܧR��Em�´���ę�V�Ĕ	efn��3|>=�k�z#�(m#4ڻ��-�oo�mv]p,@X���
;靮�SX.�a�g�7��Ƭ�s������+.U�b�Մ��� \�$nX�*J呍�l�IZ��Qn�A�7�-�d�*��h���N$�Խc����|�Ƙe�=o��|�`�P�_+JZF��!+*Z���/F�Ow;^Ca;�ckL�$Qtޥq2r��2��{B՞��{Z�Wb�m҆�K�]q��h`��;y�a�͵7&��[�j%��v�3ܘɦ�W���ƅC�]��gL�{7l���z��ǒ�����e�S?U,��1U�F���Zʺ*жb~��;�2#5���}OF:ȥ���%md{���},����jΖ����Ip#6`�.�,� 4��ɲM�`��;��jPy��4�f�[7֚�K���)�3V�D��m��o���ЈnRзs�~�N]��f��yi��yǘ�
�\��P�6�>��'#2��.>�ĥՕ�ld�qNÆ�M�t��1�8�E�eMN�t�� ���AP^;�ʊXV	��j�0nj�XY��#I�ݫR1��z��f�n��cE��x;��<(%z]��w0��r��7��u��Ϡtp���/��[s�5�4F�V��`&�:�h�9��`y�ք1�v�3��m�coS��pS��d�K륥m�ڛi��x��ZZ�]WN�q�Y���y�JNJެ�(`��[fU֫�����&ځbe��������K�RU�#n��_c�Tn��i��C��7��b��;2�X��D��4"4)˨=<8B��e6��)�˨z��c`�ܾ����7r][��L4U᦮+�=�V!��{����Np��|�,��t �[��ޙ�;�ԣ˷EY*���%\��6���=f�Jjm!�f67�9�*�G`[�q��5��t������f�J�Ξ�-k��9tx�Z�Ծ�o\K������(M5�e��L@���S�5�q���9�ϫE�Z����XC����lf�Vf]A��h5zihȃy�nqe��V��d��W�4��sZc�s%4i;eVf�����hi��#`�7�I�ed��X���/j��8�u{�8�Ò���Ζ� ��f�<��:n�	���2әp�)C�w�ލ7Sv�K/��ˁq�+˳n�:A�H�r�tT��CMR�'�!z���ټ���wk��������%&��,�=l�בB��ޭ�A3@%�U����0��I���-du��.�&�Vb�)����|]�Qnڳg��t��&��-��K{m����Z�5���|�.���#�3��#k��G^�V���خ�Y*����G���[�@S�[��p�d HC��3���+��o�jpP�<*93Y�Ӧ˷�B�ޥ��]�Pi�P�|8�TG�q���d0�2�Y��O�YԊЪV�� �('L(�3ԫe�J�+A�70����A��S:��{�e�B\��!���78��z�gkG:�KN[W;��;/�Vڂ�>�%�E�;v[�T;��9��0]��]e��dZ�U@�R��1{i3N��95��dDսs��4j�E1�޼��"m� r�;�4p��L�5�տ��v�LY<T,>�1nygm@���5.#�Ũ�K�e�$��귝Qݮ��ə��KE�����]�J��U���|�p�e���d>׉�|.�Õ����c�]J;E��� �0��|�L;fjH��чo�]��3sr���W5��W(P]������	r�\����+3m��R����];	3etl*@�U�!o��1Z��);��[�ؕ���-��GL����E�,�a��s�z�T�aT�!Y��Vl�z=��1����Չ�;W�2���?Y�q{��+0u��/
��3���wy���X��	���1c�Vh�b��f]���1 6Y�c��E`k�n�2�3
���}�6`)l�w/g�TF�c���K�.���N�'U��f����^o��mU�0R��y<A�\߳7c����P����u�S�T�:�U�`�y�	E��s@�.�U�͞c�78t�p��vQ�P�p�hr��^��lZ<G����A��D3=��FoHuȬ.���#5��OL�(�K��lt��p��-�Dn�i���+� ����*��4�`N青�shЭw�������=N��ґs4��"1��L��r�*&�m�3;#F�r`}� |���p�M�C���ӶGKr������R,0�1������;NDEδ�:;mZ��8����u�WV˷�]��D)JPK-N �7q��8㊹�������bQ��d@�9ذ �P�ũ�i$��w#�xd�&y7$����!Qy棌@���WE跺lm���.(+�
��+�$,���[�qA�˭�"��L�n��j��-���;\M�5|�|i��+:���JMb��c�R��ܖ�5փ�Ē4"�����!ن��]IZ�T��7}����A@ֲ�9�rB�����L(^�WU�0�J� �X\fN�Wd��|�ĥZL{}��I��9��b�^�{AZ�A[�BY��K/��s�}*rΩu.�R�fOVT�;2��
�Ěz�wr���S4i,w�u^���1�6�)�������'���Z�o�=Y{��"�F�۫��J��sY���q�x�N�6.�Ǯ�_d��U�RǍ�j�![��k�0&s��+GzM�nq:��.��w�2�eq�겴&��m��Q˳`�Y`m�يʱ�_|�ڵ�
䶃͑ߑǷY�]��Gl�,�˒Y;2��r�eS4�'�9p����=:�nW����Y)U�|��ț̷���R����־�ט�����].�t�J���u�ž�=�*�����t]�����s��R�ebj��yI�Z��jS���ţq�S�_�Dd7+>�kMk��R�j9ù�i�ƻE�e2����=��V&�����2�9�=�k�V;���>�xf�JAF޽4A���4��N	:]ŃY��U�0�)����tT�_*7��N:L�����״��q{ٷFy��t�VY-ս-����r)7t�[��.�Cɢ�4��^�j��|j:qc{])��A*ж�٥��xd��NB�c����)5SV],�Y��ܙϛ�I�u�h
]����7��7k#�HF%b�7�O
�o3�V���Q)V2c��IACUwS�6rqV*� y-��r$+�c�1W�À�J��/j������j��r�.�t�`��LBtcy	�C۬�m�'�ow�,ξ7�jz���z-�}G�����������9��l�;79� 34ձ�T�Z�9(�t[\d�B0*: d��,������𜴰�;3G6㼑N�l��G��bR�Tc��n�G|'V)���E�|nr�D��%M'n�w:eXz�-yͫR���ڷR�cz��m���|s-��d��C/��o�uki����G���6�F�HxKD�B�f^�|{��/)�Sj�us'��̤N�䟛�D�76η��N��u>I�!N��EU��r���ϖU.���%�1�"v����w�#���S�cff��r��El`��w�!v����嗙N�V>�!_6��;��1�qn֔X��
�,tK!9�8�)�]L}���cH�ٴ����
�ؔ|}0d&��K�����)���v�ю\�9�*Rp4v��=����SJ�ɶ����2y�W{:�	�V�X����	��.�EL�<�rV�!�ur,�| ���<��3�y4ۦ~ؖ���)ɝ��T�ִ�WL��)O��5v�|��(E����g�s)U�YC�!C�9m"J�����Z�	3y��F&6ڤ�Vf��N�7>��ͧ��y��ID!n��b3�T{.����n|fV�A�SZJ�6j�Պ�FZ(��|��ކQ�«�}n3(N.�y�q�������h�݂r��W���J�zy�*�S���j������������!b�BMΨ)���f&��C�II0�fP��Βb$븮�)��nQ�v�SJl��݌]+����	S���Ic�$�"�1\�"���n͐h�D���E�]�A6� P�1�h�)����e��0���BD�BS �T�+���A2�
"$��-���nR���!d)C.��;�S#iLI�Ɉ�4�.�q4�,��D�2R�&I�.rD��G7f,0f�wW0�"1�����H�,���,M	�46PI�;�2��@U@
����y���ܰT�{C��:D��'�rO�V����3-�;�Yθ��mI.�%7��:S�H���o5m�̜s���y�-8r%�¿�TO��fn�P˪x��.E�m�1��P��G��5[�~.{���:�v@SC�Ř���W�?=#ƃϢ��4���j����~Kr�`qN����z����2� +��b�y�J
�F.(Z������k��>8�����8��3�x�����=��G��etWz�	}����H.�Y�	�tk�UV�u98������b��?9s���%z�n뿍w{g��~��=�
�
f}ƀ���U�^ 7�p��B�s}�%)�
�p:��>x���	����޸.���7_{N���2��O��w���vc)s����}�����it� ��Ƙ*0��Jnj����gkR{�2R�~����l���?my�9qQ� ���,�4k�X���}7��^�07�ĵ
q�ZmUN��g�k��
��w	>����>�|�!���I`��uȑ�cQ�Y���j͉t��{�"�Y������!��@��=_6���yX�r �D��A�����0_1B/-��n�,ɻe��q�γ���hm�����YQvRϳ7E҇�m�fڱ���N�[��^m3VF��41��\�9q��x®��w}\F�"Z�"�6�v|�<U���8{����
՗i�M5b��=�R�����G6na��c2��BE�_��|Ԗ!�Y/����ץ[[��]΋�7~ lL,����J{�����`� '㓍Md�L^��q)m�*s�6��n������;=̊��ǻ��<��O�劂.<�H]_��͸!MR	�V��xa"�W� �����X�~��1���~�r�pu�����0��z̦{Ne���]v�"�u�*QlnS��Β��8F�4l� �S%<�h"�K8�T{��״�8:����N/2(��N�Ӟl�X�7��먑PܦL�M�����ګvr�xP��;"X!ͺ����{�u!�[z�}�~5�yp�'wF/���n\�u#=���.��wֲ��x��͙��sނLw�M6�~5��ϭ1�앵�����+�3^�`�&uVMo�8�׆L��)o\���;�K������5��za��)+�u\i�|
R���ȃ� 
�pd��r�~��/K@?�]��U\���EV���Xt��������g�$��,s=[~�n�'h��uB�4G��b��"�l��T�sR啽�7��G�����ɥ�>sM�w5���ṠSu���wz�{��3�,mn�"�ƈ�)�G���E���Z�@�Y�[�0g��7s�5ܵ˅�a{ԟU��a(�.خt�TɡԲ�>��"E���Q� ��XyRo�X5���o�u\r����յ�\z���F"X�Q���\�^OzW�_��:.Z:i��:	`�����v�f���V��']~���A��a�au��YT[-�QM_�e��<)x��A�Exo��d�-�q�|�0�����qU/\�2!lx�c�����*q��+�g�q��\-G�ZO����μ<�c$�U Ta��*�$��贳�E�*X�pЖ�\?IG�X�p�������Uz���d[���F�Ѯ`�z�R�)'����Ƌ*�����>�wVh���%8��E���6��q ��ܨ1��u��t�߹N�Y띗�r���v����XR:M��_�}X��n�mú�P�$�kG�B@����N��>�����+�j�s�������.d¯��h�5��'�Jq=��;�by�H:Ԉ��V�V���f�&�wm0��]����k7jB�S���|�vYϜ�G��Ut�Őo�����[�f��˅̣(�\qw\�Ǟ����ڤ�Q}}�iaT���&�`�Tn��n�^\D|cF���Sf�u�F�Px0�H�)�KsyŔgS�E+Q Q*��w�w���BCҜT*`�V�1
�q�}��1�{v�t�>�}[;�H��+}�:�]>�U�	e�vy
��k���I]а�
f�nX�3��d ̛ę�2݆����\"�����z�v|Y��n��^�X�Xb8���m�]�k/~.ߋɎW���4 �׾�LS��[B�g�'_��(�:���2��a՝�ws'���?y�ѫq��9E��B�S���s�������6i���V:S�𡿉���&����Ʌ�ڮ�[]�1�w���=���|��	f�N�lܤ�[�y}�W늸jE{SN{b��+d5>S����3�)�eI��n��/�9�?1[��.x=>���L��-#<
âElЊ�!�d=߼U��S,D������*J
�#K}�h&f��=�7��I���k��+���|V�旴ϟ +��c�`���kD��vb�=�I�&���Y��C~�.^V��gЎ�u���\�]�|���,����o��8ݦH�k�˼gM���OW{E�8�m�d�Ն#�U���R:������2����ػ�og��SWAB�S�ˤ��-)��%���3.5�j���]��K�w.��uΗ�Lo���ƹgg� ��6�o���g
�K,�y�&Q�f�b�t��@Ƌ�(�x�gT#E�o����=�9鹭RzUY�;d��s���=�Zrcz������՛)+�W�ҽ�Xxm9��{$V9�B.Uz9ǫ����F�i��w8M��īC�{^Q�>�eA��G�����Kvـ+�aߛ����㨟:�e���k���o��ԍ}~}X��9�P��&��V�!�7���N�C!�VY�b&��E9�qN���+�
_w�l�ݐfk0�3}AG�8<��'2Pu�r���?T6�Ix̰5��Os�Y^�>��<���8�6����҉�2��N�k�c5�iպ�J�����tT�����ϱ'�|�m�!�������0']C���騀�ߏ�5�ts�X�n�ʸh]O���\�9�I�\�lv�]>}�ǩ��w�����͋�g�Ĥ��h���Z����K�I����%'���[w�%�h��s+�Q�ޭ�
��}yʞ�^w���O�`R��Q��O�L{�	XN�4�Y�o#%1��!UU����YT���:{b�H�8t2�w�7�x��Z�e_�@��f�&��X#c
�V�=��O d��#��}�5A�q�������Gfĭ
Ǡ1k���u��j.����fD�A�C�����yN����'>|S�7~�Kƍ��[����6�}h�/��þ�R��� |�M�P�.����P`Vs*3�@�{)S��mf��kX<�r��֪.Au��Q�����\��r.��R�G��l��|o(u6�� �@{�`��I��]!s�c��V��E���6��V{}jڪ����r�n0�1��_1�V�UП�}^@�֠r�8�C�[؛���ۿx}��pً����^��Vы�:	;R�C��Hh�V+�d~{�u���7X���0e�7o�#\�_�xB�ڸb��q�QԤ� �r@�W���s��ւ��gۀ�ml��S0��J�!"ŏk�D���'G�I�1ǲ�����z�����r�,R�,P5`Tuw�:+&��BR���<�e����?�2�J�\Y�-���^�����Tp�"�s����s�5c�(*�U��Tjj�Ϝ�k1���^8zf�{�u-�\���xU�"��Ti���#
��z�g��X_xM«����==3�F�'�(��%���y�5����zO>���T�Ev�q|��?���9�:�iЫ����M�=%�f����EBR�2Sr��l�@L5V���>���T}a{��X=���Vb��� vqt��mR^/;R�U��>�~A�kʐ�5�,+YX�;e��LV\(�B15��t��9�k]}P�9�C��ytf����}��};p�9�i
yt��:N��t�JM��4�dN`�N��&di�ȷ'-a�����8Q�U��tQ�����{=V�}ɾc>L��1��x����TY��Lhu7	g�}�VM8J�~۫�� �Sʸ��Jxe�\Wy�>�'���D-���`:C�$)ɇ��0���b��P�����N���>���Q�s<�+���O����z���EWYc�����t� 7���������!b(��r�];��G��=�G����ע�p@+@q
�:���U�tb�z��oB{�5��5M矜�)�,�?-u���U��)��[wcS�tl^I� !Wg�c�뱊�T��~�a���9J�aҐ�a���]@���U�ge�}��\'(D�:H:�U�w��Bfh�38o�:��*�L�12^��dF�L}q�!����WB�G���<O�C���;�+��I�=UgI8C��֕pt�Ѿ��u�B�K�	�J>��wP��ډ��\>�J�^,�+�s¾��e:��w0�˸Ɨ�{Α�u���~�6�-A�z-�F)�;i��#�J�ٗ��`����ܸ��-��"�^��t�I\�=`q�a3Ҳ�35+CQz���֢t�6��%�5�Y�-cΊʷF���KH�WC��'��թ>�T���=�2e�W
�z��-OYNL|F��i���`��Js2�Ј !#��J�W�ҙ��0��=����5����[��_2�j8�pBG>s��m�r6���I�*D�z��P�(���S�G��:�
T�g-�+���20��X~��U��8\ƈa�H���x
N���� �R#��k-��Tf_v`��M�o�C/*Ѓ�p��v}�{��塣O䓲�C���j2�d%a�/���M�y�S�{��߬2+~�=�g��{B�5��$��hL�3M� 8>����<םV�����-o��q���2vP�����?:^Wf|�
�O���G^��ۣ(m��xL�jvT��o[;#W��1��LS�}VЧ�yu��m�t�[�2�]UHO8*�wV�e
�Z�kleZ�����m��9�'�ݹ�>ʉp��8b�v����_Օ^#O�;Oy���c=�c��Xz�*�앷Z��-�+�o�|��	f�Z�8p�/dL��܍�t�7"�b������:."���~,	�U���u��ȉN�+�Sb3��i�g��>���~o@��+ٶ������1|���/�V*đ��!1^���!�z�b��6���0���EsN'�Z��r�՛��K�]#���Y��u���]���n�im�J��&��Ö��\���͸s�}%��c�Pꔒ�^�t�X)��fyx�{�*�U�&Jo��ڟ`�)ߨ�#��ZxJ~LS\��P��x��+�X��-�ȧZ�!�}�7ᙞ����fd^7Z�����2�� B�2�����z&��S��=x��57G���+�|J�РX(��Nu_{Mt�Wq����7P���+D`�.�ۧBk4�hl���,�7
�Z3��>������#�*Gʇ�"*],m���޷VƸ�j�n�w��%����0�ӟ=�#���deú�V>WP{) 2��e%�i3����+�s*��!�T�����=��
Tc�]�X)���r���ŉ\�\~G�32 U��	�E�z�D�u�J���X��l��W��P�;��N�@6����m�ѓgmV��F����-y6#x��)�Gv����(vWV�y��C��-s�nt�����2��=KI�O���*ʾ�`*�������iD�L���Kk�dC70�z3�-�q��\��7�~;7^TP��C�NX/ )�����V�ב�@��#�����>dk�N9Dƚ��4�s��Ϟ[���׆�3Y��ݼ�O Y��7:���b�f�t3��V�OSWZF���/��>�<�G�x��Z�Uݡ=��yٜ�9^{S"��.cm{B>�?^���cރ��m��87z����9�'`�u��6��i
��$Ť+'Y�ޅ�/Qc�A��lF\-wzs��M� �S�b�y�J +F|b�Z����#N���M#�T$.�6׷=�0~c�ӿ/�����V���TįL����ɼ�m��mQ��:S�-y$.f$S�\�l����Y7-xs�uÒV>��=������>�2<�-�ވ磞ԧ�Ei����U`��x[�ٔ�x��Uh#e�]G���~�ܽb,�zgn����h�T�G���=0�'X���g�Z]>@{eV�X������'���d���k7{%��{e�k�t?o�3������ώ
��u*��N��AW��ed�>���U�/�>`:�����1q-S��z-j����t� �{]t�{޼'��}糞mo��3��9:1�K3Q�����!����|ڸb��^|=>�D�6�7oMm��p��C��Zw�O�U�gϕ|j
E����>��������b��|��s������.+>��k+@@׀��jt8VT�<�mP��;�0����}r{�B��[��Ιv�pl�w��s7�!�"ĮWՓ�P�v�mI�AЗN3����V�L���Ռ�Sk�L�BeJm3I�FDK���R���_��a����z���X�4�����B+T��i�F`L%e|�x���l�v��Fє;v�[�[�
l[f��n���9�PXj�����Р��3�`�Ŗef{��R��[�g���dz����YL����]�*B�l�����3N(Ov��槽�{�Ǌr�4s4��كɛ��+�'�GW޼n�x�C����#4�ֹa��Ov�=��x�~��k�c,��`��]�N�ىt�q�	S��Ҹ�n�L=��@tml���!Uv��Ś
��;�&+q�Ok�9��o�rδ���P�w&<ҭ�ňPk V�9���)�ɫ;�s|�8a���%ꯥ��-�e�c!_h�z��dN�D��/x1#���^70�Y�Vl'tCx��l��՗s�7!w�6Q�u�F��)V2����.Y���`*��5w٨�8j빕N�M�����~8@�U�}m\����䵹�h��)-�3z�f�E��6�*y��F��d�w�N�uP� (<�X%e�9G�*�є"ҡ�@�\�R��v���jY�n]��ʊ���Ɂm��F
u���
<pקW��n0 7)��C(=7��u���	r���[&pt�""k�M���[��yz[���--�S=z�X[qot=��������K�fJ��U���Fr\����r��
o��ͅ���	"�-�gm�o��[�xM�̢��w0n��kӁݩa{�Ρ�j��*���۹*�3�Ǒ��$��q��CR��;9g-�ڻ�o՗%�e*��J׸Yx�-AE�bf�l���+�\Cѐ���\���-{g%�i���O/L(�gbz�.��VY��jɓt�]��&J��>Z����Kr�G-c��8�����,���W��֚�zТj!**�xO�m}Z��l���7c�	�PJ�!��Y��D�Q�8qug	"��㝇ѕ�K���e���I��E��nhK���R��`�ېf�)���!�p#1G��\n����v�+k���yk�'�����vUD�+#8u��Cv�f��c���}���E��8��o%�\��>��\r����9Q�֧)�Ȋ$��Q���	z��<��Τ��2��Ӳ�Lv#
������4�tȂ+�!�/�;�U��ʹ8/#	�X�$bɅ�C
h��7םcq�ϛ%z�d��	C�N	�h�gX��nc[����i�$b�����	�gj���2Q�x�-�u�r����t9�M�±v����D�Z���o*O�����r���:��,wH�;nQms����t��E�]'j������y�z��xK�Cb��m�[ǆ\
�N�O�e��D�E���e ���H�TQ!D�L���J$HJHF�F(�+���22b%,ɢbRb�6k�� �
�SL���I@�(L�1.u��QM"�dJ(�)�5�2$Rh��dR�L�(�B(Id�&�i��� �))�#K$��0&����a�($�	��l�B)	.�#$�2)!�"d�H�1BR�1� lX��P��L��ba�ILċ���a@���'wcf�#�$�`ň�J�X HB��w],"�0&h�"Œ�P0�&��~^�{������Hwe�GlA��5ee�L��yޙ�6�+Z(K���wx�X�(ސ�U�0���M�Gev�� s��9{�k���`�f}��<�|}�=����׈��x��ί;�77��{��J�so��ξ|�����[�~6�o��Z|��������or����~��1��DVJ����s�<oU^�l����1��"@�|�~>�G�x��|��ݯm�ۻ��]_���Z7��v��۟*�\*�-��������v�׍�y���^���׋�����k�#�&�} ������,����9Կ�}׊�Z{���ז?W��6���W��m�v����J�7���s�uE���������ε������������;xۆ�?���u�ס�׭�|_��#�|l�F9;���L��֎���,��7�[�~+����j�U��7����Z�{Z{����{[ҹ��Ϟz�����M���|����5���������r�����0�ڹnoU����[����ȡ�N�� ����"�S���2�;^����#ﺋX~����@Ϫm��^��W{����7ſ^5�����^֍���Ͼ��_���Z?ߟ}z؊��W����o_{csx�_����U�so�b�����" �"+<.�sT�q���җie�D �ƌG}�#�c���w^��mʿW����ߏ�/w��������W����������^�]��\�w�~�{�����Z7�Ͼm�nx�k� �@��|co�½Q�%�����oF���,H�����#�/��[���^/�w_���o��x�k�^->u��ץ�����������m�v�W��_7�����צ��D��1�����`�9�{/7P�W�D�b>���Ds�X�� ��F�y�Z>� ����/�V
�U|p����ߪ�W��yzZ7�~7�{ξ�����^��+�ߊ�������R"B�DQ"�>�>�#�C>z3��d'{��uNVd�jE�X��"!"#����ڹn��1_V�����z�����ү����������͹�Ͻ����m�~�μ[�x�����j���x��:�߫�ѿ����5�W�^������P�>�]x�z�JG`"<"�D���ڼ������Ͼ��\�����[�}�U��_<������|�����������6���ϋ��m��6����_������{��o���]��y}�V)EOq���#b
���|?nX�����6s�7�IՋn�8R]�힊J�<r�{����;�Ya�kƃ�R����]2��k���r�wS@��3v�=d,�Q*��&���{�7��;A hY���{N;�/���6�,�8�K'���((j�غd������k����}z��?W���������>�~�������T�~������׋��׏�{W��}k���{��|_墿�������_���Ͼz������菵e���wVr�5���A|F�.m���˻x���^u�o�ַ�^��#�G�jb"��|����1x�������_Ϳ�����������޿~t[�T�t��P����>�">� a����W+��[��x��{�ޕ~�k���y}6�W����Kz|j��thDP�B>(���cuh��""�f~���}���c��Eq��>�bѝ���6��N[iBI*=�H�	���s�Z��oǏw��+��W�h�_�y_��^���o�u_��z�w���ln^�{U˕����7ϝ���՚B>�>���q[�p��@��{�1������R���ߒ���|�1��}+��^�������z�����߫ϗ��V�-���ﾼ׵�:�7������m��zU��:�wmϋ��W��Ά�E��1����1>��}c�!F3��,�}��?V{} }",}!����W�>}�oo�|W��7�^o_�\��1���c��2c;���`��G�F}���,��E|�J�b����}DN5�1#���I�����3��:�TT��{�b7Xz<�H�(}}�dG�#�$D}[�8���_�⿿<��^/��^��z������W���=-��[���������^/��zU���_���7���>�
�����꠯�c�>
����ߡ����Y���#�Έ�'����""/�����۞�������o���x����o��ޫ߮���o�y�zoKţ���/�}_�o��~}��*"�W����b>����G8^�\�s��Y�l�mz|�nz[�\�}�>y���߾�o�o�ޗ��+�ݼ������������ߍ��k��}m�x����h����oQ��#�>�F|ۯ��f>�>�蘭�b�P��͗�����8=����̞���m��s��|��KF��=���4������<����/Mx��=���5�w�/տ�E��_V��k�^5�����W,}_����j�.o�������P�� ��\u��}yj^fԞE��5&I���5-!*D��8��Q�1�h2o�?���f0��u�@d�Y4,'�q��%��i���=�txv!���� kz�F[�͢5����V��� +z��Ԧ�,���j�VR�ϙ�)�_�|�U��Z6��-���p��y�XM8�u���P꫺����W�;<�������/�z~�?����^��n����~u�Mp׿߾W��x�W�^��?�k�꿛����~�kF��^�~7������{����o���K@
L���}���\}F>�";����`��G��U_D�cG�H��o���[�������V��j��z��������o�ܷ���/��m鹿�_�|����vߍ�ݫ�����o:�W�ε���n �دo�����%P�=������"Z���x���k��^/���Us�h��������to�>��_!UDQ�|��s~��_���-�{Z�~|�z��}W�������x7�n�W�*�^������n;��+�U�B��O}����s������E�[߮��6����\�k0��Q?|�B##L}#�|I��;� �AW��|���ޯ�����m��o��^/������-�~��{{_�/����na�/�b���"_��]��ߍ�禿U�}����c�|^���J��o�^���]�[x�������޽�5]���}��}�阊X��#�|��_��ѹ�=ߟ=z��޼k�\7翾[��#�H�C�}G��P�r*��3}��;�\ߪ�/��y��W��h��~y�_��oM/��ݯ�\����i���;�ͽ*���׾�5�}6�����r�|�ߟ<���\��w���m�,}�����˽�O�=����t��~M��7�}������m��/|�E���ǟ;_�z��\����s^7��o;x��x�k��{�-�^w_W�Z|�{�׍�>-��{���}���3��Y�J�}��ܟWv��Έ��堾�����޷�x�����z�oֿ�|���r������_ͽ*����}��^Ƣ�>��+�������ޛ�wv�ϋ��z�o���^�����@ G���j�^�����պ=M���t\�}���G�D{T}�0G�oK����Z�����W��痡��ύ"'ܪ>��D|�����"���x~c�DC������4H��\W�����)^�lr��k	�Q�5���#B!���^"[��^+�s��N\;�ŋ��@��B��g�\Q��j�H;}Y��]���X�r˘�W�1�"�c6��KGˌ��J�[{p��A�;���]ͼ=��9�D.���[�[߷H�>>��g�J���)
j
㪄	���$�F.��mu��
�qwz�׊N��Y�z�H�U��G��v}Z�-����ـ@��:�4.��`��w���"ڲ�-x���>�5�)=3==X�/�֧�9�4����G�P@Q�N"��4��w�뮞ςh��z���8�Ƚ7ܠ��sFtyDF0�1�)�toL�􍩌���#H����u�uq_H8�ϔ�����:�7t0E|ܰ<^@SC�\Y�?k�rT����ح�x��"�{ꁿǚ��+�����q��a�n��9^`yg���B]g�Ĥ��hF.��VUf?Lؙ����@�>�f�}�>@0j��iߕ9��(��V�����T�!�4�� BgylŮ�7w!:�@�>ֲ�b��x|�=�~Y�yH�*�J��>���k9���:�n\���IJ`��z�'��F�(�f��� fW�cD�Zx:q;3������o=g��޺�Y���p%��Ң�ީ�<^�V�>���Cd�J+��ZςҸ�� �2�
:Ɂ��{ݣ��/������W)��5�o���=�տsߧ�3�� �~��,L�]z�y��f���N��R�܇�I7��e�	K�n�J�ț�����1.���-@ŮT�-^W����|���]��Equ��5��T��b�+7���&v�M}�k���i9z��,;��`�\θ޸�����S]����ڭ�)�z����}�G֓�@�X�"*a��F�@Ta�w�6b����++F�U�b��$�Df;��jy�z���r�:�^�>�s-�����%�Nߎ�x\C��5�4;��[�y��Y�z���E8�>*fH!�M#'�Ә��3��U�v��<�{��v!���T��c���'���wT��O�m�2���V�B� ���jw@�7�wl��Z3�siyԑy"��ӧK���ކ��W����{(�P���@�<$�@�^�ۂ��=��)K�4�q��2V��s�ٌf<0���x�X�*��Ti���-���٠�Z:���}([����z$��z����3P�&�u�����`�F��~��j�]�a��چ��xl���YZ#���F��'��IJd�M�j�[?PM;/&���2"4_)ݣ{=�*N�@�,��ħX*�W�G���g�;�1q�~D�r��3�m�ws�l�'jJq�W<���:��~P�Y�*���Y��+�Xx[��&k��gy B��,j7��;\z�^J��Kܫ�l��+�����5|yR<�L\i�6��܎�,���Z���`<���z�/{޺5�H����	�Q�E�Vy�$��S8�K"�;���,�S�q���э>ji.�d�W�^t=�mH�Cz�&ir���K�� ���}T_+<}�=м�v5�J�����[�	����n�t�����`��o���������M��^�P��퓱}=�t +�~��Gm/�c�2��φ�k��{�����L���b�&, ��������;��ў{,�-z(��a�I��e��tw0���K+����^�z�m��ǵֲ3�U����c=7p�F5^��*Z:hg��u�N�7�
D���+��U�>@huiW�Ϫ�:��><̯9l��j��(f�1��7ٛN�/z�b�>���Ψ��Ep����m{y>2!lx�c������|�H7�5n��N*>��3��|*��� ;hc���xF�p$�o��u�B.^<���ll(�ӳ�v�z��"�]�2:�6��ҽcq�3��o**��=�G˸Ϛϕμz�"���&��t�J�;j_��z}��i~0E�!	_'U.m B!Y�O[��A����_ V��da��ƳX�o�)�D3b)�Vq�n�l�G'\���G�
�6�玔���7�U�8���%b痕�5���li��@�^����2	��w^x@��vL]xP;-<�Z��>�4��o�/+���f��f=���Ep�9�2�ht����/M�L�bk�w�6tc/���8i��[�ɍ񹔸��$��т�Qy���D}��cN]�6p�6"���3Zk��Q�m���ha�H��׀Nm�I�Ejb�R���;>�C�#2�1t�W�p�4���.�u���1P�vYϜ�G��������ׁzwZ���TL?�P�F��F�S?lf�b�3���\�5���{��������Ư3s�=������� �q_XuY�A���Q�T"��TY��������_��C1(�2�*+Z���N���V"���b��M�4"�\eH��Dڰo��q�V�����Y���I\�\�a���6��x%�e��`�{lC���וc��D�� 0���\&epI��'���LO;o
�l�a�5�W]kOx�h�gy/�>�y�>�`s�zWz����ӭ̡7�-�1}�b8%�;��:>͗Z��6vM��ȻH=5�S��t�7 ��^p�Ѻ�σ�p�ϩ�1O��q�n��� �xz��q��[��_f�蚕�����wZB�ӯ{�-,P��Ҋ��U4���H�L�7��_9ܻ)��U�f����3��X�4 ����A-�Q������?`��vŵ�=�J�;��mMB�,�kx�teK�T�zZ�W��`G;qH]��O��MG����.�2��ݙ+�г޼�'������RB
��c_`�;���V2�着�����a~m���ѬL!�釲��eehYUc�@j de{�*i �n�v
#��1>��s���&(z���>=����<k%{�٫�w��>����� �K������I�+|ԹK|C7U������뉹�7�/�H�U�dc��V�τ��`�u��+֖�7�<<h�)��@��a3�./�>e�l���'1�_<u��g�E%/2�y��߹[���m�3��Z�2��&.���`��|~U��amYg�~����t�����v�^��ƴ����Z�҂��E��i;\={����kf�q�ռ�c�/N�ʟ�~�K�e��(���>ϔ�:7d��mLdD��Q��0�L��^����i	^�����1�����iUѿ��`��߂��.,���P�福�õi�`8�U�P�D3��1V��)^R�k��W�Ǔ���ȵ�C�7pX4'^[���Nrm���y�����y+�0�x#�~�9��(��V�O۾��OiR�U�G�c��. z{wי®�P���)�(gZ><N%�Q�i�J�H��ıa��j�m�^�E���܀��y5c[�>em��}���-3���/�g2��wwP^���5�\|:�3')��b��TI���^����*HUM�C�b���U}�y�Sީz�wD���r	��la��*q��+&�Z��=�\/�m��Ww���-�n����o�}q����|�E���(�0QVeW��U��i�n'f>^:��(�W���6�f)Ǟ��{N~:מJY����{i����8T��e���
�@vJ+��|�O��0(�<��	]�6r��@�� �t���,G��/��?gdCo�I:Z=�����0u���7Q��)ث,F��qL��K�0|��n��1��z.��5�I��)�䀚��mo o@��.*d1X�l!(�bv�u���#F8���e����t's}�����,��D �r�X=ܪ4�|Wr���Ňy�G�ԟ�iN�}TǞݥ=YW��9X���k����+@_\ G�S�²���@�k���>���&ojΆ�&7�f��zR�>���yQ�|D����=��L/;��X���k�T�|=0D���C�k1��xa5��<��<(!�����/�F��=e%��Wڵ�,U��§@L4Ir�E�p�CSu-�w�9��^�6��v������Z��٫˞r%6l<���;@�"�ܽ�%�=Y������M��,V��y���Fm��*0j��R���	iJu��K�	�c���N*��">��<���
+�0�����f��%�n��׃!Bv}`�n�n}w]됕nn�,�t��?����}���8��B i?����S&N���5�^�g��wg�<0�ħ�Ӽ���a��/�)�0@�yn�[�FJ���\$�U_c��5�k�; ����wk����0����0�p&0*0�ਥ8�_�(f�r�3��O�C��N�$�IME�rmؿW{*Xfq�`�&u=��Y�ڰ����{K����V�xp�Bb�]���=I���V�̸�3:|�t��k�t�g����K�^�&��v����Ec��r�:�T}�b3�����w`���_sn��^ڮ��z*o���x�O��7h��g!4���/��x�(sz��>��x�T�W������'�
�|��Z��4;5��^�Z%�����ܠ�rg�w�/��� � âpw�i{UJ|��d�aL:�eQ�n[+>����M]Ed�����f�@�(��ł���u�\5��pik�)���u91]0��}/�����Q˲<���g�#y�t	�n���[���m���TD���9�[7zH��]���Juw���5	�wuw3��Q�7�u���tb�&#ݙ/��/6«�ŷ�"�Wa���~0��>J_��w:~9��{���qc��y^����	������1Qp�h>:�9��Ρ]	��Yv��P�Z�4SxR��xe.����.��Ld�	؛R�����oԩ��g1U�ǱOj;up����r`��*t�JI�W�7^4�Z�����G��Dͬ��{z�N`=��i�<t֊�D���BX�ik�̧�0����1zc�*;��%�,r�}6�~�u��C����^���feK$��Զ�:t՛�qn����u���d�0�p�;�F�N���v��H�����}k;7�-������ܗ؂�y��)s��1s�
|�Ռe����vO
V�-;b��j�<�$@V�Fb��:�*ٰD�M�Qp�6�[7���b4�PWW	�*�TO�m�>{�=�]��:���'�7���K��i�-MQ��p�Z�+�>��V*�DႮ��[)�[�=�)C�n��ё� v��^Ȟ����m�VMk�1nQr>�s����̗��U�qxUJ�	����ǽ`�xn�T�K��w�xa���"x6X�v�zQ�/'�^���j��}Y0O/zk!M���w���ϙxM�4_!��n�o����Q�v$]7K3'X�ƾ��c[��^����:����d����, �a�2#��)MJl�f����)w)����4Z��龜*O.�b%��A>>��������.�F.�Mi�N��L{I�R![�:���w��Rܫ��C�W>�k
�níeL4r��U�m���F��M��V��#a2��]	7�.��4�x�󆴱rg���"�I-c�R�\3W�h������y�KG�*wf�w�[eu��uz�NXB�Li�3]�w�_}�;gu�I�Y5X�����<Π�k���S�%(j@�h�0P�ԴΗ,�7dܮ�6=��̙��`�l�5��\`5g��5����������N�	��s;�|��1�PmZ�v�Rk�+7(q��]֚�jFڗ{X>�4������lg۽%ɹ�
�3��G�'.�8 �}6�	��Yr}h7,
*��n h	#}Ԡ[� �;����9n�F����2T��Oٺ���b}�"�Үr�� v������s��xh@Ub`R�JT�+g��`�N/���=ۣ�f)bҔ���JY���R�t�REe���l\�Bڡ��Q���:��ᚵ�Ik����K�<��ieF�����)G���S�P��s�H펶x�X�_<n��6 �3%������y��j�*���m�.v�b!��F�#!��5��z库�9{*n��7�I�b�],��'z���<^Yf�z3�+��c����`��|s�4�a4���	%�3(�̦���t�iSI�wq@i"�s,�����9����$��J1�c$N��`+��()4��k�q$H�fM,&#�0+�%	JHld�&#Bh�6@wt4�
.[���І���"�"���̨�&$�H&dԖ1gw8���ф���RB�)"3��jL�1	(JPQwr�1C���M���l�QG+�3�\уd@�,Kd�(�a�Ww%,b�2d1f����&��%� |�TEV�
��-�K��o���5]Ι��`�W=�E��>�*��g��y�^B�>ﴣ�s˪���k�R\ýIs#�}U�W�=�s����PF|���«��p=��GI*��	��)�\$�o�t��5�zmY�]��y���Ԁ���q�Q-���(�ౠᨄ��8ܙG`}�ǠO�R�*��J*3�OV���=[��~�_c��%;�U���7D{M�L��I�K�D ����h�IO���J{�{W�����t��N�-���t���$|b����G'\��t����%Y��cI[. � �ZX��$�3>鯰��U����As!�M"V�^&�g�&�-�w;=�˳�����m��#vP��yW���N�x��ևO�h�0�tYQ��e�s_��J��"|�F���^g��4��.�V%.^��2s]��,�Ymӽ��ܽG��f���8�i9`p�����*k�2v��)A���$2���{7�CҜ.�E�\��U�Ah�56BN�F'!�PX����LS��[B�yu����]�� ���K����}�^�b�C�*]+�B#�^�6ƒt1F:�'r?v���*$b� َ����sf�Z��b��u���\����/�xG�uq�]u����'��o>'AXK�t���?l��Y��/V�
�ËY�Z��s�-�_S�7��`,��Y\���1���M��l��}��t��i��dɂ�P8�8f��+"�������UӶ��{�^��-܆�x.eV�N�93�#Y8Tx�~�]���#�g��d�y�צGUw��-'	Sšk;��`A�ko��na��Qg|P�G�.����TO�؀�{Y�t�<��&��t����_��i�����\#a�P��qͲ��/��Wn�+N��"#����R�7Ғ���Gr"�hk&Fi��׮t�5|~�(�|#K�gϐڍ-7������+���G�l�x2��2�0�)�����uI�+�?i��h>8<�4�U9�8������g�eq�G������C1����o�HnK���zrJ�� 7�����T����;�!xxy�(�i,���Cpީ��{$G�߈�~��Ü���}����WkX�d�	����k�k:"�/��׃Ȗ� W�ð�Ǆ*�[����tä���<����O�$�bW�kǨ[�L@:�4%b�!�;����11�~�����x����m�C�]�w?���O���3R#�P@QӃȺg��uV�z}U�#NC�U{v.�RR|¢��
��&!��Y~5��5eSι�	m@Z�N����ŝs��`�i^�]�����rѝ�Q�^#Ƿaz������e,�:�X �����$u�d�*3ۓ�-��n��nk�NM`r@��s#�<Mt�{�hq�چ�۴?���>�����:����R(~��O�ۭ%�3,rX�t�Ԧ�ѽ2K����Z
͵�@x����}�����i��8�Z	*�7�CSr��yM\Aqfƺ�%\�����V|�TA�y���i��*�G�E@�ee�7L�t�U�09C@}�	|����7f����Sէn]�v ���F�\ؽ������kN����Wz�x'��^p������~���~p�Z�p��#�]�`տ�p�-X�����r�nU�\��p��W���^�ny����.O9=]���o�ٮ�,ؕƀ��\>��	�E)`�P�����[�nV/Af-H�S@�;�pK��;�Cu���k�h�5��l��E}�����ǳ]�4{=��ך7`e�i�"� O�Rm<�y�V�-^{�|�����-$�#���wu�E��A{[߽��z��V*�F�@W�~C[u�Q-S�J�躩1`��\����]�`�O���l�h�ݨwS#DTD�5���8�<;�<lJ+E�k�ϋw��6T�0�f�����蓟{h|aAbX��nnR�7v�T�J���"���TL3z�����|�<idb��6��r�Ş�3Et~WZcf��&�vVr?M���D+ݬ��i����1<��B!��ڵL�O����vtJ�������~����:�X�-9�CV�=Ȃ �ՠ�ZS3��%_�
E�ם�a{�n��[�y��I-�㦚�>��P�8���� ��+@@� [�N�
ʛ�
's�δ.�r�[��z����(y���x�'�T��N`�P���	�b
TJ���zu�@	�g���#�o����j��9Z�1,�|ۯ ���z��f������5�X���o2�4�v�k%%T]������{�P�5T9-��Zf�"��&�`ڪ�S.r�G�V�o�x�7=��vQ��s��M=>�q�}���zbB��2d��4z�W�S|����mOD8���,�8��b�L`�/-���w��-v�ww�f-��R�#���jk��g �Ԍ{�0�������X�5�6�~50��2(!�0�P�ʛQ�П��[YW5� �f8�D�Q�=u�Y����mXHWܯA�_Z����~�E�Ѧ�c&�Xo�Pų(���ϙ����}U�(���v+�_=���F�kG^�`�%x��Y���7Jn���ɜz�p�/<ݿt�qSZ��-Q�o
���(��KJ,'l�`Nc�.���WR'g��}��:3t�#u���nQ���-�ߤ�kq��]�C��W)x��4��3�%����k`Fw��DG�ͯ=��[����%i;q0��m�������o'�7_�A��E��V�v��B���o��t�6A�Y�z��V�Y�Q<@Y�{�-s��C�5y=�\'20)j�c�y�����EkgC��Q>�KF��T|������e�t�|y����*��-8-�)���&�>y~�b��%�}�\)xǨ�����
���D�׷��NLWL>~��bg_�œݯc�t���e[��m|�B��Z*\� ���>��\/䖍���ܨJ�[0���>v��#+P��T��Ḗ�?�icA�P����}R��>�Sc�&
T �)�5NPnwVx,�������Α�u��U�����Q�eC�MBuR�� =F�RʓV���R�"���8�UP(d��Ya�[��NR!��[����C6�����!��K[��v�ǉA�I��� A�k:"�J�c =;�
�m�s��4C�D�)1b�ڞ���g��Ո$���bW6����x!f�Y���;����K�]k���؍YH8k8�X�Fݘ�f*@���s�'' �AF��}~�uu:>������0q:Ӧ���7`��3�a]\�K�;p\�{�y5l�1,�(���{�,ѿ˦Π	���h\�:�hW�#C�=쮰:��g�?�����{�ёt^�v��rUY�����y� =��3*�/��95���\�e�\-���i��ߴ{۴�g�ǫ~��wt!��e ����Gj�y���WCW��� S=r���kstn.���y�X��3y�S��1⇂�e{Ɋu��hS�����6�y;�&�U0*3e�'���T���]�[5��ҽC�o�z���4�^:�'r?v煾ʉ:�:�v�##�ߜ�������a�Q�c��Ôϸ�2��G�u�Z�� Z>�W���wbG��W6��_n�cNN�b���N��c��&#b�!�R������Y�U=x*�N��n��KQ�4"�ƫ�53��*�A[������ɊuIHGn0��Ӳ�V9���~�6�Ő�^�E�r�ܧZɑ�b�^��B ��=��^�Ϙ��k�u����O�y������0��
��2���{��礫�
���GI;F~���y�lm[~7?2����x�С��7�y
g�E�s:�g��ƭ����s3�0��Z�U����9�*�y[n���7p�?@��nQ�������W�2T���ǲu�Q
2���an��jq�f�q��M"�tw$��\`p�`5PQ#xb�X'}�u%�9xv���x��xQ�fȘ�=��s#sN��B���A�>7�m������ꪯ,��>��0 �!���l|���l�=�u;�R�p�3T�ND=�#�ݑ��JL��~ݻ~�=�5�X�[Di�H_�A�1�苏�/��׃-�f �;�)t�����X�[����|�uת�ݵ��g��k�P�(1P;�LO�*��;��(㊆d�^�̗��̠���VY�E�jw�3N��M:7�$.�8<��{$��ã�k�����=��j����܆/����ۭ%�2�ןQ�',}�)�tn4�/M�ۨ�Ko}���-'~�����e
�U½W�v�Jj��pܰ<\##<\Y�1����#o��}�����d2�z�<�v�T�+�S���0*}���]�:������׾��=mf���G�ؙ�p| �ţ`���/;*��'�;������iw�g�m��>�c��<B�^n�t��B��H.��@��^t-X�T����\����eU�m���=Ck8�ՙEmg���s�V���zl�ٖ}��v�b��3�р3* �!"��'eq� �-�ي0�3���n�Y�7^��r�W_�����/	�,����Y��.߫#oĪSl��*d{���f��Fu���q��f���r��{�"0�N�e� �@�V�`ޡ�
��}�os��Y��*�+8g8e�QZbЁ�m��Jva�V���^�z�#\��<�y��V<w���T���K�|"�����s��x*!��3�wn��5�:�yN=��[����ш]��4�Q��=�SsK�t�m�K�<׫�^�v�9 x,O�.�j�w{|gOxA&N񜯪$Ǒ�@�mL���.�����l��T��^���l;�G���H�]�;���]�i��%�/���JiC��!(�F'o�Y�,xB��N�;<}��\*/RۙN�BR
󇻰�8��T��F�o����,�Z���5z�ƙ���r���VL�C^N������c�R��3�H0��^�{�P�"&����Z�
���o=��O�[�A��/��I�{=)a��}_'0Y�����J��[��۩�~�����oǇ��0�c�!��SV�G�r���f<0���m�R�2$!Q��]οy�/*���؜�6F��q�gރ���W���%�:P�x;k�+���>��&_�}��y	q&���"�8����5�8��{��[Q"�JS&M���5�1	Ml��������!y���"L_�]\\���?�0�Z4�ӝ�+�����Ǥ�ޤ�Ǚ�r���.:���El�$��c�\�@�@:7��r�S1uc̫J���j� w��Pp��U���}��r��>9ӯ69��ɒnv*���l�zT~���"""^�/ZZ\N��'�W��ժ����~���v��j=��!'wF ���Bk|-�.�_��e�.����%o�*��a�i�	������}�����)��ZS`rb�>���H����܌�t� q��µ箰� ��?m|a�&�eA�^��h�93ok��e��_��C�<�ݾ��=�t ^Y�{N힘�l��B����w�PR�b�V�
�Jd��� ^��=�����o1�J�{-x��NLO�5�gI�-l"KL�U����j���g�k'�
���U��u�;�,�f޿&d���4��VΏT�t�	`�M/j��/Vez�C��hNô�B�N!��^<l+���i�J��iL���l�u�W��P��药o'�
�V�c=�*Cשd0s��n9s��g�^ʾކ�LB����R�wr���8o�3��77u�O���+Ώ��מ�����3�|ϥ���x�C����A�����_%�mC뿈���x����Ǔ%7V�1wvZK#�ˌY[LQ#��p���K����c�����B��`)�s0�&��كt�9/�]�U��6v�*��5���ٰ�6w��I��4EZ��N`mhǕp�:m�t�Vv�S'2�V~�U{�UK�g?��?hn�z��D�a���[���o͌��o�:�5���s��"�RUbU�C����"�����^�����SI��I�`�����^7�ñ��>��(�y�f�Ʈ��q���o�(�;jt��z_�έ^=��,ŏ]����#�1��ҙsQ�-�M�^r:_.�U)fˬ.�l6/�<hA�1�{^�عR�O�;�\y�9�\N�s�몶r�4�w�Oz������d�zi<���z�U5i�5��o#�.&5�;Q��Zy��!LK~q�F|�t�qa���$sy}N{a��z�7���Ͻ�g��긬��{�&�7�t�W�Gj����g+[J{�Ơ���S�^�j��4�ڄD)�`~̿��ClAfC�$��B�(���U}F?gO�-�{Ϡ�E���>�qy{�e��q���o�2����9���F(7�A���"ĤdU�k�I�[�u���O81��t����& D��
�y[�vԑ^췥l�A�B��g7N���t�i�� ���Q�9O�'T��KR�|�D.�)��v��nK�n�B� @��RtV�[�R�������[��g@1u����5�!���R�Y�׃e��{�]�N���V����|�r�5yt��,����̯v���9���a��yc��������˺�N,�ȗM�K��`��jټ�����q�1���F�Oz.�]�1����3U�G�
��cE�9�7�j�&�ogd��[�}&���_B������IW;�Ⱥ7�@R����
\�ZR3�\n���:�0V��K%�M��S�G)��g�b���Ѣ�p#�즫)�����KN�����%DZNʊ�#�3E�"չR��U�iJz�I�rs����s��w��܉�����9�t9>Km���s=۰�
XWf\e�ʾa�2�w2�]8
���;�(�Pv����|YuиzA��
��w��e�uJ��m3v,��&ra	�#u��
u�;c�h�%��l��R0�j���Z�Mvz�Ұ�<؃��������J��e�AZzM�h!�-�/nY�y/
zsyMP\@�Y�]�o}�/!�o��E�x�(R1��ku	��+#���łU�Ƴk��30"�7R��}�L]��>O{�t��	T7�əu�y��)���6��nu:U��{���igD���9ާ	ycG�+Ct�����ĺ�q!��iFX�b��qg\�r�UxW��d\�NY�n��4".�s�,($'ZN�-DI;2��vl��|n�vr�^z��l.��?t{��ag�|���^ݬW�:o�`'jܾ����~��\�M� nn�r�\����V`��'����ߎw��\�%���Isދ9HA`��W�c���ZƛB���c���2�KkwKh&4N�wg����c�O��Ǹ�tـV�%'�X��%�8,Fz.!��/yG�#0�;b�J�Y���ŨL�T��v��񘀲�->kr��r���6����z7����T�0/7u�?d�Գc��zˊo���:�y�R)�Pg1����7���k��[Tɴ�Bs��Ż�L׮�k�p�m��Ad�	j�c�|u��ǯ��Db���|tF��1���˺��(Ş�<��0���ĭ�e�q�]�a�/yL<+�L쎙:��,�V���2�N=��ɠ���E�W�w��cSg%\�N� �R�؎�8����%�wC3��m�N����"�#!}d�r��f�rT��ً4�������/�$��L3-�"7��j��W>c�Y���2�V���Al���D� ��[w��,����䮇
jm=��V���?b�g;w�r�HFWv_zY]�U��^g4���}4�e�|>���2X�n�H�ػ���������D(#IS0iKI""�I�
#h�1N�L��� �i9�I�;��i�D�I����c	�DE#&Y��Y%9�щ��a�CA�ۑ��nt�F�ܹݹc	�B�"�� �;SID�E3	�.k�����F���M%(,!(�A�@ h�u\BH2�S"4IR(C3)���r�4E0�!,�%�œI!�-�J��!LQBdC�Ʉ�$����D��
 }�
 }�%�Q��3{V�On���|�(<2=�����qf��pڊbñ֞�M�����R`�ӥ9�q��Grǝm��UU}U_>(���g�R-����x��)){�C����*���M�T-�t&\������!���fc�\M����m��ר޷�|�@������LnԈf��������1����j��c�R�ǋwxᬷ�����f������l�:�oЕ'�c���fTI���V�DV�n<�\C�^���p^6�E��j�*g�cI�s|� 7Ծ�>�_���$8�|d�hH�\��|�9yL��-�f+��(�b�6�©}�Lx�J${^���/_����&*�c�)��Ml��õ���|�s.qL�Q�-��W<�~���o��
Y5a��<�o�v�c����w͡P��S�s_)�5�-����٣�#�)������][�����x��BZ�z1�#�0��P���h�@������r��g���]�l's^{ɯ�d�g�+ITխ`�6���������z����gf�u���1)�7>dm-N���� #�G�S#�J��eٯD��s:�B�V�3��'a^*�'r��v4� 7��{�n�`��eŊeK�[��]J��7�:�	���Ys�;�/�D7�$���Z�����ܹf��ˮv�Q~���ﾩ���~i����?���!.���j�,SO��bp�[P=R���6��n����-j_z�ݪ�U̳鶗"�9Z�=���Ng�]euZS�o��z���s�O��+�a:�Wp3+��~��ߊ�y�w0sI`�2������5�3/�������=K�b�d�s���É�,{��&��<w<��
i���V��S�܈m9<��X��7�5��B#2ۮx�'�ŷT����'*%��£k�*'ړs-�(���n5���D�7�=j��޹�xX��w0��/J�^��-\x��P��m��Ob�V^��~y�/�9y���l�AUIݨ�z���X�ˏ8k6u�ĩ��:����l�-���+���s��ǻ�#�����zڭ��u7$����o�G�KS~>�����2<���T;����U��:�3�;�^-�m�J+mL�PtB
�����_j~j9��E�Ġ��.ct|xj�����\Q1)v��'ܗ�V9���V����$1�a�,^A9,9����Tp(�T��#;ݪe����R˰�Z$R�[�u�V=���_*���%��ӵ2hw�DDC~v�U�Z�+���PSݿ���ϓ��|�T��9-|נG��aA�W����P��O���3�;�����2�o!ÛsP�J�OYs��΃�ĵ�W�fy�^����{��ծi���l=G"�0����+V=��,ah��i��cT}�M{m;�W�<��ښI0b|v�VVL�׼�%WY�9V}=[Y]����ګg(tH�yb�ݘ��Iy�V<R��(�rg��Ҡ5=귵=�~~�X�W2�=��k<���f���U~Œ�ˏ1��ջ��m���5n���s��y7q�&��������Ym�c��;�z�H^Ǚ��KZ�e#�Ʀg;���?g�^E���j+J��j���Yu��������5�����W�57��θ�/�r��y���u4��;�TS�d,����[㝋s��WT�C�>s��Gw7_L���4�b <�H�j�� ��\���7�݂x���]|������q��!-A�u<��@~٪���u��]�8�u{Q�tGZ�����h�m��s��r>���g%��[���ȏ�ӎv�+�am�g_*�M�Z��:�I�qo��着���.����O��3U�E�N�f������W3cϐ�5x��3�g�)OV��r�Kn^�
�ɯK��6K�V�	73Ӛ�>�wӖ���s�r��~d�����8k-�/T6���Q�R��)>���nS7T��s��Exʓ�\�h3
����\���y��+G Ԉ�}�7�!����B�>���YKv·�l^l[c*R��[�s�P��M�f���H�Uw��Onz��za���)�^I3�\ڙ�-F�N=���[]c�{�sJd�#��#�������ӏ��/pL]p�ݓ�?N����M�;�r'���)�5�-�M�W���9�&���oM?x�*�i���m�m0�̸�B����]������+ٗ��Ɯ��"���73�[k=����^��͋N���y�|�G�\Lk�v�R�N����n����}w�&���	�k�����{���C�*k���cZ��צ�]@VM���Րv�ɞO8'���z�̧�>�o\�h�ti������IzR���Ѵ̵,��+�ro����ER�Y��f����T���j>=mH�|X*���U_}�g�毻�0���c^o��oJs�z�7����9�#	�/��D(5��+��zi��U[�I7�-�+Z�����.�S�R�xM�������k7�i��C��ˈneL�K�!?Y_.�wύL���{<���}�l˼�Խ:��y�=]�L���������C��En�W��_U��&��'��r�54E�JJm�}.���7�Ʊjc3h�_�ז�e�`�@T0'=q�U��Q�#-\Fz�s��ۗ�o�9��;��l��E
xP"��i=��N��U8�9�ƿb��<[��c�~/{<z���<�ajxfB�0���W�����d'�%�R&/u����\?����L�c�"��BWuu=�M2'�����07D�iT�N��_�5[^;�i������Z�jKd���eF�5a���Ӳ�1}Ֆ��fy��{ۥ����e[����T���H�zNݙs��;f�ilɝv�,q��t[�^��%M\�}�lt{���ygd��$�붃THGŅEo��}��[��Ƹ���;�xt�	��T!���=�1�'%��שֻ�v��>���?���>����jܷ�zR�my���n��D)����oޡ��_J�Ƴ����OT���{��ƿ.���$Ұއp͡P��T9�(�9�-��3f�d�Y~U�Ua[2��&����.�-sM��иI�
m˜3SC�k'Y�=�%��]L{&�SɬY�v�ٕ��`�Cn=��{2������s�"�{���VH�U����.Jf��
�W�sڕՒ��o~9Zӑ�Y�y�Ʃ�\	R���л�K�n�X�W�UqΠ��#XwU�Ny�tuk�Nz���^��i�4�V��L�K��l��Ncx�b�q/rayp]������ޯ���*~�ix�F�ZW�j�:v�ջ��RC����.Z
���Z*6^�����7��y��y������T�w?{�Xܵ갞�<U*��\nխK�m��/s�b���$#��Hѵ�O]ַ̫+��Ma�	���*b�lۋ,�=���B��j+�e��c�[������^��i����{ڑ�9V��{o��H-��R-e���#��С������T�a޷)p�H�W�J' �d֟Kw���wC���磌ꪞ����/�ҙ�DV���W^�J�U�Z�����j�{���F��ku�u������Cro���q�˹�A��ưI������ᴓxǒ�;x��W��1;״2=X�X�Ri�������hz(n��"7_�f���=��L�o4�d���x����f�[є�7c�Z�W����R�e����o�׻C>#�y���e�;�?U��k����ʇT����|�1�r7Z���(r�h�w�S�F<�UD�<Ұ�1{�SI��le��o�_C�r�X�����ڸzhB}K-?*�<uYv����hB��#zf�zr�v=YM=� Ì�b�L���=��5G�����w�y��]��K�sw(eNcyib��4�ƿG��Yq����^�S�C�C�q��5(v|��+{��S�V�>������U��U?R�~��Uk��ip�9�yBf�L��z�>]�(��EL(��T5oU��m��Qma�P�KȘ~y��-d`�}rs��Ⱥu��������,Z�,ɥ���)�їs�-�Dۺ�p/+Z���L�22>�PjV��T#M;G/*�wћyx"�ֲV	���\f���rb�K-c�>���ל-��c}���.k}�y}��5�_�Ϫ5�Mߜ�ov�Vj��o6e�4���󈗃*#����ٕ�p��y�;c�T'y9����fy*��t�� �*�{M�TKCk��]�=F�y�U�'+��x��0A�<1=�H�\zx���io��,8<���1F�׮�r��"����٭�0����&g>^�V��~j���Q��=+��c����a�O�/e7�-�M��z�+�&�.�����;�N�E*�w2����/W���Ί��x7[ᬷ��y�����Z�|׎��W��sm�Q�H�ӓ��);����3��f����y@����2:���Yi�x���������?�2|٢�����W�i�����7;v���$_���9cs�f�>���_ue[�L�{H���~I/WU��5Wv#%�²M�L�{qR��s㢼�����F���kT�+�Q㙢����w��j}�75�hZ*�\��<���<�l�m�Q䥡��:6S��ASl��J�rwL��.��Rl�S�} k-`�7,�6ClΉ�&�#��bv�����T}��	;ֵn����C�gյNiL�_F��ںu=0�����~�c���~k�u��C�����A1q�ۚS.]i���&�m!�i�md�w���2\<g�lϒL;�eǝ��)�ƺs�^�6>8�{�C��wL��x�k�R�~��X�%SV�"ی{�G�\Lk�t��_��e�8խ@��X�۩�ax��Y�:x��w��O��>�2 ^�+���]����(	���=7�K�X|�9Zڥ=�#��L�>�S��@���ӷM�|P�7��k߷�ߪ�߇�Ir�8�쟭m.�G|��VdG�V�K��s���y����=w�N�s���V3\�-r�����R���B�����qe�����"n�߅B��/�{��<�m���m9���:�6��K���_	0?c��v�2����ԛ�m�}/^ڜچ՝�=O�힞�20:M^e��NOc��̾�߅��|��{ދ�zQ��F`����r<<�J�vl'�A*�c�3;hj�nfO_/�n��y̻�xN��"�j��FU�W��ӋT6E)}���we������M�����<�n�8TX��H�����^��9g�l�=���N����R�����F8k.���Z{pVj�A��
.&����^�k=$���z�K�%긊�2{���]�y�;���s��P9q���8��
�X����>�7D4�N�RX4wE[�BV]�� ݞ��^Rd}��Ɍ��-̭PK�Rc����׳�9>�7m���V����N
z�ז'�z�o�yq'�~�_P�47عg�����5�!�NW���#}S�T|Ƕw����ݳhT6����B�s_ifs|=������B�����x��O^mgyf�����Z桷��C.<���;`dxNz�����	ny�3���3n�z��5���W��%3���Pۏ=��WS`9���H#��X�ԽF��ǳ�׾���"[U���K����Ol�^k��oaK���J�.��o<�Ty���������Ҟ��h�(�p�r:��}y4�+;��/�WYZs�k��DbF����^3Ό��먼����B�g5j-�f�x,8v�����J���V֦�J3a��gt�v�أT��4e5�*;���;i%o:if)�&��ˋ��ޖ��S�V�fs��Y3gp�EQ��x�;�L"������t-��+�˺���0���"IsR�:�.h�����jnWK]���;�Te*h�=+�U���o�u�Qt�q�t����z��]���2u�Յ�z�%�V�,�ݤ�';���+����.�K&��+`7��(%@q*w��=]�t9]�a�x�,�%�g�ߞOE�z���
[�xj�X�)[t����܎Òb�"�=!� �N��"��}Pw\m�tE��n'Y#�(�D �uXl��B���#�1g�֮�T���56�t��Y�d6k�
(iyq���v�v��f�(��-[��r��Y��Ͳ�].�S]��L8)���r�a���^f�]t̂�ё?�_26\b��K���ج3�ը��`�e��³�#D۔�bܭu}˰��vʉ����p�|o2�s��V@�o3��+S�6�"l�c�@7J�Tr��%P�nuǖ���8M˃\,k�y��Zb������C뚨-A�y�z�kږ��L�6�ܖgD��{��m�.�Q��z��(r��BY��W)�ZƮ���W�vK��iǞ�j�q��(vג�5�'��G�z�K*�#���x�"�1��E�\E�B˗Ջ�y�S���J�Ka�3�����i=�G��Dֻ�5\���C�1�bv���9�h���}	�	8�=��㰜���t�[]em�G��P�b�U^�c��Ԟ���^�S}�=�y�(-�Au ����Gn�"�)B�d{��5�������c^%+R�O�mSM�kq����k���ȗ��W�u�B6D����Xj�/q�/��D��Q��Ⱥu	�]+�c�(��e��U�vzz�����ٳ%���,&�ɡX��^�k��c�G�q���ά���̎
�O�Ga5,ʉ�Ŋ�M!ƚh�mV	}����������C�#�L��6�O�����3o�Z2�0��R�ii��g��x�Q����JJ$-51�T����;��1d��YZ.������Ե��k�+�V�"����ս�z�03C�k1Y�f����?kݣ�%Qu���q�:ǻ���9UVރ1�j(���{�XW@K��M��h�NcK�6�L_u����YX�����k�\Q�ܵ���`$�i�o	������E���+6�`��u�����p�r���	���a���S�i��Y�%E�A��
�i^�&f�����D�.]�Pj��p��7n��Υ�6kQ�B�.V�dO3�t�*��v��遴Ǐ6�\��1�ݽ�ɍ�V�mU���X�����F�2}�P��|  |HE&ř�,���$�g�F��@��ѻ�chir�m;��b"#D�h5����T\�J��1�.%�X#	i�� E�r(L$d����Tdۗ4F�F�X,i"�$"BQ����qS*1�آ9�wv�r�De(.c���H�D)�����8E�r"��1�%��sF˅wU�I1�w4`Ѡ�s��n�0lQ7I,!!�,��	$I��͍˥��뤗:�؈�33679"��'u�.u1��СP�S�I�,cA;��Qa H$D����]w��0�,��0�@P�Q}DQ U��طܧ,�s��K��j�王Fz�uu��7������}P�=	�ǎuq���G��1�b�:{�S��L?� �:��.�y�>է}�1��x��}	�ʿ8�^��_M�E%�J��^�޿x9�Tt��OP��p��;=ޞ??g�~f/��r���ł�%3�n�g���?boاJcm����[/\\B���n޿mc^�Aг��G���T�=�{��wz|	�>U�j%Cڌ.7��jM�SoK��8�NM�W�����C�z{����eܒ�A������R׃�E�Z�2^�%_?��6�d��9ʚ���gѽ�Ϣk&�wo(*��8>��ͣ2]W|�J:�Ɩi�H�n�����a��ecw��Q@S}蘀�~Fiz���ٮ�����J�V�!�=�/q�>�KR�ތ����}�~>�ʻRh����	���V���}f/�m�qBF��o�uG�
x�S�SP��s�Ŭ��'1n M
M4���~葹���+SI@w�ػm��liD[q�o҈ô��)�g���T�d3�d9<<s�U����P�����Ń�}��+��X,��*���Y�i�r�5��a{ 䴠%��3n����l)�$;��x���/.H�#@=�c�!��:\�q�YOV�ƥsh��WS�6;�zג�f��P;=�'ȅ����of�{2�'{�y��7��f�E��=5���m�=t���	�����Jy:�#��c��׶ӫ�W�<��ᐿe�Ţ|��92�v{��>���S�q���:^�㲃���WǶ���@�g+�6�^P�O�u�gdz\<��Z�k�Nm�O��[Oԩ��*��j�.���$Q�M�����X}Y'�|�>.g��w��O��>�=�x�&����>�"��H�{�����.��9Z�]�G_������O��/4���[U��˨�m�=��=IZ[T�.XqnO\�]@�Op�(w�C�&�pў�<����e��|��^+����8�Xs~�bڬ���]S�Ag2���i�O��d�H�^���缙��|��$�rh�V�Y��hu��N�7����g32�~�L56�z^�_w��˹�=*�f�u9�v3�Ԍ�����v�_X�ie�GD��:̸�Ћ˺%c0��&͙�|�r�Ťh'���2mR�2�����λ�R]�ۊ�q�V������M�\��] ӏ7�^DO�o�ۻ���jv[���g�����ꇬ�W�0O�| Y��F����j���t����5i�s���P�8�m�w��gkai^̬1E�1�;�ݸ��!j������p�'�U^P.�{�<}�	̽ U����ޛ�ՓO�}������CH��>l�Kv�+{�z���1���8�WM�tz��uf�`��
C�%eZ�<ۋ*��.}$���Iƕ>��*`��q1���`�ި�����S��2V����{%y߃܋E#���{ۺi�ld�Z��7��C6��g"a9���zGk���%2�!}j�^�~�nR�`�z[�?cҪښ�$ö\y�iWz�d��o�z_��-0�Zf��x�|�<}�U���<�œ��J�ӄ[Q��ߗվW��T7&3�Bf$bώޱ���[V�߳�nr�4�e#����iw��h�x>��z���	�p�����=/^�U��CpN���Jz������:�,PWm�r�:�-]��=�{0u���j��H�,��a����ͷ�Iih>s��Q|;8zdi7u[s+��z>d���iNk]�0��b�[{`w�+Z���I�.�F�<�����V��W�(���1��G�A���q]�%��Δ�&�����W����H{�2TVrs�o�~�}nqt�A�������֮���č��س��YE��2��6ob��W>���E\�z�&�>�.z���r����`we�;:���K���|;��_g�g�s~^�֛�hq�xI���^�'�q��m{-���鴌����z�s��ۉz����6�ꜳU���sYy�n�@/�n/��:G��uo_�#Ż�p�\?7���{֤-��v�
���:vq��J��η@�G(�;y��U���Q��ǜ5���<~urK�g�r��E����N��\!��0*m�[H�O�Ia{uw�j.�'�˽c$���6��Ϟ���/�꒸�_j�1�][nzd��JxfR���;�^q\���&�:���'�
x�S�s_)���}�.��a䆘��+�y���;S0�+p7o|V��	x'���S�sP�|��kt�����V(Ros���=e,�e;#SY�}\�<؇u���xg����!�8�vW/XQ���b�˵�0�˗m�^"l�ƃ���>}*e�l��&y�R���3�r���r��.ts��X#9�Az4�tLz󴘈Ѩ!�jN\C�8�Y�W�u~��W�j19�Ҫ!-s_6�;eǝ����ڋ���ћ�����Ŀ,+7��c�Z�޴��Ӳ�����t5K��^$7��,�ȟ8
r�5�ĪmX�M�}�Y߳��qT��]��K��X��m-w�zV����5�[P=P��Y��W2�M��~�%���}���p��Y�fvj���:�[��mr�y�%K�zQ�Y��I�{�&�nRe��_,H���*���S3�������<�~�{N��0�="����,�k��Ng�nV���6��|gKٞ��\�����Hb5�Yn��n��.�Ibc'��9��*��\maQ?{Rne��S�4�L�U�~������^��K���]��tϬyTI{Q*5R-Tap��c��4��ޢ�/5j��W����US�Y��ܠ�_�mV	 ��H�us���(���B¸t�����yQi�	V��o^|b�wF�	�7�<�˳�$se,�AI9��[��걛�3�.�F�Q���~�P�=���t�s���ڶ)�pn􆱰���_f��m��ݲUYU�.�Z��v�7+��^�ЛO��ju�!�{�8���D;���<��ᬷ�_6������Z���,��g��į6���;..Z����������kע��[ѕ	�w�]B�{n��ѭ~>���7~��;���U��n��z�B[�[�d'�
x�S�R'dמk�7 b�H�溻yo'
k�)�G��\L�X^��^�M+�;�l]�2N
��^��0�f���wѶ=1ѓnk�2V�ۂ�����%��)�y���@�Iz&Oc��������I`��^�6r%;b�M���;_����}9�:�p?S��&�mef���g��ѷ]M|�`�����[;b�Ǩ-��^�Ey lȚ��ŕ�����N:�{��ӄ[P1�k���W2�sY��J���`y�7=�@��Xb�Ƽ�H��Ng��W�Q��f��s�'��u~n슆f�W��D����lfz�鷵/W؜�ז��zz�<�)B�쪯d��9U�2�u�V��^my��A��3�pR�7����uf],�u��"'6Y{J�.wEԫn���O&���I��r�aV��Ľ���s�Ijw��Bf�ڵe�f@�uB��/S��C��i�S�N�-� �ȝ���ƑFs�������C�|�k-��T����ٓ�Vڷj���===\x����N�j�X��(qϬ9��ſgW���Ŕ�Q�ӱ�ߒDb�������q)�򯱯NϜ��9�힩ʓ�����u��o�"��і�0���A��m�/_��ڈO�x컙��2��	R�:OQ柞x��z���2��ԥ/�q�X�l6��
S�[C�>N�?J(�7k_xM��˼��1�IN����>����_��?��o%`�a�%J�ׯ
.��qp����>�(�Ҩ���͐����[�f	R��-�'�'��!Kգ6e�'%��T���zc�xc}�OGB^�v
oɡ�����&���`����r�+�/!�郟�I3[�����r�ս��wyl%��6���r&�(�9�-����	�f�J�w�*zn�A�2���+w���@ux�{�ٹ�$��vY���_Ik��R��o�u�)�����X-��;��޾Ù�VA���33�c�e�t��#z��c"�g�#_�>��Z�C܂RYx����(��C�"� IЬ�M��*쭩q7�5���U�[SI&��=8�.�JU��V���F��_f����w0}�˔�j1d�v���N���?W��=o2���N����B��lM������Ks��|�<i�l]��ǂ)�y�&�v�i,��j�Rq����5|'���t�����}qgT���z��"P|�y/'�YO�j5\c�v��_>�9k�fT�����0������x��&�R��Ψ�)�6o-cQ�+%9�_��u�,��׳���W��d��pb�h��^�	���=q�k���V7wZ�^UD-�m�ރR1�9����p��*&/Rnr"�{q/\�g��n\���5W�y��K����.�{���*5Z+TG�wc�����K�O����ѥ:�ۛ|T�U�=�.�`�z�K$�WJD�{���W���QT1k��U��i�$�Y/����-�WV�'vQ�olYчa�])�Ӝ�:F�T�0bN�}1A�Q��݄hU�b�k�\�X3Us�'-̃^�zi�3*0n�^]��#ɞ`nѹ��O��c���F�`
G�#ՙ��f-J|8^.�*���jC:m�{'_���^���©}�O���?�I��z[����zv�7�S�O8[�3�G��-��꒰����x�Jй���/ْ����VQ�Lf�O��i\j.��+5�|8�O�f`��;���+�:��:��٫�3Y��G=�({UM�ε4�7��3h6�<�ܜ�ث��*rmv?9qg��6����o��f���JA�k��m�w��Z��	v&`�j}��Q^���MOH�R�e�T�֯�{��6�Hr�����s�f����<2����
r��.']�W�=n�����V9�Y짣�~:�˧)ö����pӭ�n���z�nr��0ל�^����$y?3f�w?5)v��ޫ^�{)0���w�yxx8���Ӝ_�ҿH��5��4��a��=���7<�.�G|��39ٮ�O?'��^+��k���k<�h諈��{�Ef��ǑDǍ��鏹j��/{��(�_0mۣa̧p���{���5�hwo_��*�a��A�B6Y���M%i�@(��Zq�WY����lP=="�Q&)��<p��-�p�W���{����Mj�V�� �
��f�d�6���h������n7��W�{������O�qh�uǞ�]Ս�����K���P��0��
3ړseU f��i�	m���N%�[�qCU�E��B<����>�N�,�h�J��&���w�DZ����+�^���y��8���.�Pt/ӷ�, ���u���c���ץ��m���X�ki������Z��%��[*[Z62����o�"JN����I��X��=�oF'-�Ypm�Mٌ�[�%U�>�A�03"F���~5-ۀ������H����:m��|x�O�Kln}�/�y�+.w�}qekBs�6��̙���zn�'�u��-v��J}�Z�'\��v�XG{S��w*�zo�0Dǆ*m��[*[Z�b�z�D�v�|����Bځ꒼��K��˻�@]������7(EF�H����3 Y�{x!��/HB��d%j�}�H���{:�8^ꝃ^qYG,���q֭�J�nK��a)F�b�]]�{�q��-18n3��Fo��� �����\V쑩Y[΅��`�Ղ�dg6�k�����Z�1��6��#x��˺�̸v 4��3jy�ǯ��47�d���s�pA�!�H����S�����f`��&F�|/Dѽ8p�.|��i��u�Fh����dJ�����V�r�cj2`H���NV%>�|$eX��͓�v�6��@��.e��y!�{l=vҁ��F٬:��vx�v�-�݁Q\��"'b��[Vz��;tA��ǔ��u�+�+"�̦u�'���]��wL[�&�:y�7�ot�/j�7ܺw|\Y6��4���(/���;�PV���ڽ�������Nl�0{uf�n�;P���R���v�Oi�6�$�V�4ĵS"�*�賙��{ka^3��Q����V�<�C����8åŜk��)ۑ��\'q\���G����O]��c#/�U�Sb���_�y���R5��1Ty��ąړ��7����q�m��i�u����:�)��F4b�Ҽ8(7��sq��X���r��y�=��w2#�d�����!��)��ג N8���I
�C����o���0ѷ%���#Ea��ʲ�d��u�ݷn��S�¥�3ܘ�'��mC9n$��������f+_,��ٖ��{x������4�>��sjN��b#0����M��gkM#�6_,G*[���d�����Ԯ�A &-BN6w��;Qla��زl,{�`�=�.ƶ��{1oW�v���Q������\4�\`�n��s�ޱ5Ֆ�\���<��z�:�������#pi��TuMc5���̫��+�,�btg&����ZU�(ٱ�'[�Up�y�{%���4��;U�[���C3i�f!�1lq�v
��uln��X7P�tYw�C���sU<��>�q�IVi��U��4�Jj:�mҬ�uu
0K�F�J��w�H��m���iX.'}��yneeT��7��R�l��nq\�����6m���2a�2o:6��"s�L�]��Ϻz#��[&p;��U��68�.�7��x�t�4��\���{.�|̋:εLq��t۽�3m��hpL���b�����V��&`���;�@ V6�����;M��@+"��}j���+Dn����-9�~��[X�C���oH�T�8h���IۻW&�އ�^i���I�_-���{3.,N�|
w��E�h�꒥h=r�8�J �]<�.�����XvĽ���J8d�yZuC�x�<�ʎ��wb��iӂrږq#�hvq ��e:�����Z��n�p�cbъ|2�y�8Pv�n�u0�u�P��r�� N��6��7�8�A�@;�Ssn�wj�ɓF4H]�2k��4n��1��Ҍ������
��H�$S�vw0h�#�w[����:%AI��\�`�h��.\�1�������H�F`[�u$�7ˤ$�ۜ��QJ�D����#QsN�i(�ʮX(,��D�$kuب�+�wjNm˜��[�k��1�Q�u;��F�c��E	�rƈK����]֋r�݀\�T[��D�d��]�eݠ�F �9I�n]*(���5�t-˛�u�D333>8� �g����cf͡mYw��,y�̕�ݭ;"Aw�n�A֙V#ና���,��װ� T��t�8k����ܩ�d����9f��ž�p�`�&����r'�.&�v�=>�����G�F�����vs�xVn���ӄi�ծr��2'�8�ܘ��������y(���g��nyy����K��'�[�}mϝ�eޱ�O�i����d��Z��Z^����֮�#�k̊��|q��J��ΤvsIN-������X�V�����8��ƺ������g.W��+l�:C��yܨ������y8g��^+�V��9Ua���gW��y�C{w�L<�S�K�Y�WO������r߾P��c�m�/�aF\�[a�����1�i�J�m!���CՔg[Sp�{K׷f�k��@ТB���5��c�A>��ĝu���t�+�Ż�Z~���W��ة����ZͳI'~�v��y�z~>��Z�$�Rw]�Ia����{�y�1v[N�UWS�j��zB�3Հ��]���[�mʱY�ÍG��^d��[u��}�����:WF;�gJ=���חS,9lv^�C/�ʋJǃ��5_�s4,��RiZ����m!luv�0����Sb�9�%�Zή�_�J6g�הz����C�A(��4�蒲��6j
�_j�k+���I~��{'Y^>��uJk�亅���1�J*�ٸ�X�V�"r��?cލ��ۜ��^]D6ϪS��L�[!m@��k=Ś+-7
=v�８�1k�j֐oCb�[�Jv��4������a[T!e\4���Y�2�f�%<��n~�ҩ-���Lx���~<g�ޣCp�ۓ�2��z�.]�x�seŗ��z�f\Ky8���P�����b��e��0��7)��q蛛Q�;l:�^�G���[Y�̾H��=��zbYR�X�H�=��j���\'Z}q����u������wΔ��]b�^���Nõ�Cx�[�*����!����;q��}NoˠfQ�şM�E��P;�����x�ۓX1�pb��t�p�q�bes����+J�g^{Fy��������W��WXǀ�Z1�߶�Z=��&]��rQ��%NB�
j&�]%Ǝe![]�����^�\�,�g��;hS�� z��p�k�u�=��n�mpb[�ݛ�!'j�j�$���!u��3չ{�
�dP'��=���K�ch�_:�)�&��,�Y��ߗ�^����SoK��D7�kӹ2���9�c.����n {�2*y��ֺ�]�{qTM�M̶������O�M�!5���~�T�/{��6K�UD�����X�/�c5���j�wY�{TMo�C�d���ծ�wo���Â"�R��*V��QUu�kq6����k���j�����K�S�F�,Έ�D��d��!�ny�ۜu�AOr�V5�E��c�^������֠=�B��E=����U^��Tl��p[Jÿ/'�5�9P��ЦJ�F9�&�j��U��/��Q��SR�������V���oC���y��W?H��{�ۜy���,ŝw�����Y�f��s�jz���f�5Qٚ��4�*�Q;�W��N��zG��j�e���Zw�y����Q{FTr��zM��8��� 4Kk3�[j�I}�}����C���]��nK=O��tG�;h�[v��Vj����&��E!nVMW�fN0��GOuԐ=���rGv�+.�
w���e�=��˒ƚ��y��F�3l5���|��n峠��MC�3 <�Kr�q�0�g����6�ާ���-�~�J��ˠ~�����'�������[�t�3��W5n�����ځ��k�!��q՞��}a��� �벴��	�a�zZ�;����ީ����9NjVG�����cR�ѥZ���H�����Oc�m�u~�Q�:V��;���~�8��&qbwRn��fh�=:jS�@�O%imr�8�Vw�j�gK��ժ_��@��G�5��~Ԕ������Q�ص1���@��k�]^�gն:����1�g��8����\�������קn+@����|�{��Q�ݦ�j���ܬ��Ş&r��-w��{���^�m�נj��j�����Ķ�y:om���$6��[���qJY�M���Yp�����V��aU��3~idsL�ֽDJ�^;Ϫӛ�`��{�߇w���nCћoE�:n�U��"��`��@���s���u����/�Ih��wH�P�>�"���X����"��-�xT}�m�PV��l��}�SL�퀖�	��X�jv�u��ϕ;���_ޞ�.��HV�g �����!���-�a�}��o���]&N���_��Wެ�s�_<�<Ǝ���j��ݕ���y��x,���(��e�VMk���}�	|��@^��^�����ux��ޱ�����z�v�����<�W${H��Y]�Qv]χ{qc �0�Z���l�Q�2᧳P������?'lW�m�ij�/9�g�1&�� Er�vy%m���]�λ��wz��7w�LG�\L5l�K���ndO��X�?f��d�T��a�|8�5��5rS7�u��֜#Pہ��\�y�C���>�מc�������-������_,GO�3���������3"�y�-��ݴ��mhÒ�;ɴ�_�Z����Ԭ���>�r����R�Owoy�ޯE�gj���\���+��-���.�8��uW����U�6ڏֳ��My�t�P��E�'�K�c?r��qϬ9��g�6���ar�Wu����Y+Wkl�<�Vs۬+��D=5N��V�3��&8��갯i�5>FچfI��A.����H�>�k�<C��,=sVWZ�CO�"G5������6ʮ��ݞ�ެwl�E�����m��m�ڝ��i�ٰ޾B	3�vP[7��o��.'ڵŔ��S�\C~X�N��cu��~�n�*nzgZ����d\��{_�Wm�Q7�5-�����ͨMz^��P�i�s��\�jo�u� O|dT���t�j�RߣŻ�p�[�^���;�vwcA�Z��š�Q3�aU�9>��)TI�wIa��ˍpצ4fMV��]�{^�J��m#������*�ڧ��0;�|=���t��'�܃A��rÙ=�}���nU��t��2_K�PL�~O!W%g��L^�`�%�ڤK�A8���;ko�V��,�}��m�9�9
d��e����.f�s�����:���¼��{���Z��oC��mp�Bt�!L��*T�O�P�m���P'#�k�]I��ԭɨ��7J�KjjL;�eǝ��soT#j��a)�}�7��Qgs������Jy5�3]��eZp���7OA��^�6����(KwK�_��&����0���L�c�3i�$����x2�PZ��\����rn�����7f�!�p��~�"U�/�Ҭ�ޓ��.��.&5G(B�*Wy��
����c����2&�=g�b�=԰J4��d��iL�}��,U��?�����}{�k�G���^M��GOT�`ѻ)�j�g�Q���GV�{���pM�Z�W������艷��bQ��y/�Q:��nW�x#��wZ�̯\$�]�v��P����~��#1g����h�W��c��q�eF(?]o���4��m�z�y���'���7�F�o5���~�m��TM�T��������)�������o��#䣝�1������s�;��q.v�B��¢b�&�>��{nj�S�b����Ck�|��')Ü�4�짠j�ځ�t�����w˺a��Q�(���/2ko�4��%�Z��{����hNr���;����X$8>s��g����=��^�Ȭ�n�����^���e�v=�R�T���/(̐�Z� ����NN��'��)n^�kq��U�2��%a�u�T5������ڱ����]�yY�&�vF6VW+{G
�0�oI�fpy_��7�Ēuv}�4r�xr�$f��MH��וlC|�{z��Xݒ���z�LzN�Eg^�4�9�H���w��/,��.�<�18a�+nMd��l܇]�r�\��F��8-�^^����%�F
���|����m+���	���7�T����n��B�;��K3O�k�l���k���~f��V����3���V.�YrA�w�FW�}P��#{B�٨�Ё���ԯd�'?Fn�_%�`�;zS��J�,{Ig�����<ظ����}��/Ҟ�`�T�7Y�_u]�3*Ɓ3[>8�>V6��T��ްk��y�9Q��Vʸ�Ohz�DN�H�b����-]��v2^`�zz;�qջ�uV�p�Ouu�+u��-�����;S"��ռB'7п{�~�xk>��+Z���<c�/n#�w坸�3	��6�k��l��V���D��9A1�����K�-�P�����w��?g��ʽ隣�x��f�zE��v�,�>�U_N!޷Q�Z+e�4*6/����8R�ꭽ�ߪs�ܲM7�����o���Z�R�#��A}�w�Ef��t	MLL�XڑL�� eJ�L�׷	�ҕ0e��������&�5��g�
pnЫ�vw[�/yݮ�X�s�澹��*(J��7�ҥ ҧm��wb��4���k�j�X��2��w�ܭ��<[��@��f���@��fs���W�v�9M����놼�>ƽ;:���|�$�^b=��(�S�ic�ƽ-��.&-B�m��-=�+6��Ү�������w�M�;xqת��ʙz�)J5�ˏ8k/��M�낱�������or��Lz��;U� K5 fi��w]�XBN��5�E�����]���jFvt��������B��<^��"����t+{�Eja�-�&�V��Pm��mS�NK���L�	|��|���},���k�tr�K��n}_~�snj�U����J�dƵA�.���j��y�(^���G[z�7��H-;b�ۚ��Q���Ǐ�>�u�L��[>��Fs싰�}ܘ�FpĘ)�ƅ8��v�t�U0>E��k}�W��/UY8H���5r�SO�ۛE8E�=�r��b�Y;�}w������	1֖�c#g;:�K6r���L�2Cyq��v�� �vC�r����P�-C��X�n�`y[¦'��{X��V	a����EP��	b���b��x����!��2).Pp����am"s��nMN�:�ܠG��.��^�깕V��K�9-�9y�|����zޯso�w�Fl�Yf{�tO5��Nǵ�+	���e�M�K��u��.��]�hHT�w�	�%�d��D����Ã<���V(l�������z����z����J����~D�8v��Ψ�)����NO)>^+%9a��_�\��VQ;���>��`u���1��==W�ٿJy���Ʋwb�n�>z.|�E�:y�y�dd�3N����^��^��{��?g���^�:v��|~������RS�ߪ$��U~��+��iw��ȷtz;��D�>ϣ��{��F�Ԉ�x/�y�qt
�D����Oe]A���C�2ٺ�Aq��v[��'��A��&�������ܮ����)����>���-�s�t	��@�-�Q��d�ǲ��C�t�T�^z���=����ӜV�wI���3z�٫}T'��!Ha����EP���e�l?1��T,����~��fS���˔8�N�a��əpB��9|U0����/b=*^�!�0a-�0�3L1F,o��</2<�1؅+��J��uf���;)�1�i��Fj�ȳ%�5)�-اQyX�[5`	�Mm�N4y1��'��U��);��-R�\:��9�v�b���������uM.9�<��|�Eb��"�B����3���4�3�s�'��̮-�a�^�(��g8�b�\�L@��-ԓ,�}���R@=Ȱ
E�����;�O�e�F�����3ƌw����ݹ�S��%��7��;�����5�={������v���aV__K,�K �7���&�Hi�tz��qԤ�3%6xi]�t��y6�6�M�n�댷��#x�,q��T���R6$H�ħ�q=�"/FhgݗOq$��|a`mK�v5��ӊ�c�+	
��������󖣭8:^[%��$4���9�sq�{'�uY;S��4ͤ,<'K���=� �5�t��KG��6�G)v4���l�7b��a�-�]{�U��C�w��+Z�ۃ��;/�]gه��TK.�b�m���)<�;����)���Wn���ؖ�Q CZs�±�╁I'�p��N����j�v�A�M�����u6;��Md��(�F�jd�ot,�3pŝҮ�e��Yӕ�l�kF%F��t[�� 0<SzD{;k�g�k����E�!�R�Ǒ�����#�C��0ڑ	��jD%�x�v�A��_>�D�єp�K�j�m���$g��W���cn�9����N��
+��a� 
*Oz��z�T�(hTѯ�|f\��(��;!�H��ng�#c���wއ��LU]^����{�A<G�̰o����4P�ԇ��h����	���m[�N$Z��Z�쮦�i�V75�Uo)f
�q˸�E0K�ǩ��	�T�opC^�5�˨
�qûx٢:���5蕁��v��]l#Z�:��P�ہ�͌�~xOkZ�	nY �Z|�)a�Q(v7�d˶6$�v&�Cw����b{@���A�G�yA�wu8�	<��t�m�4��s�ss¡)�Ҹ�Z���'vu�@1�B���h9���\��s��b�8F�3rv�9f[�O�ȴ\X�
�g��Rˆ�#���h��jE��'>{NO�E�Wd�1tS���A#�Ƭ���M�
j�>�V���:��1%��w�a;kj�Z-d�&��I`�L�w
�>���C։�Ǳ(rlW@GT��I�Z�j�7�z��+�E�X��e�'�"�Xkk9�\s��z����a����&qfg�=�:�ΕeJ7�v���T�r[2�<�Z�zH�$��6u]�Y*�h����
���gB��E��7z�M][�b�� ހ�XuRR�RɾH��fV�ͫ��O�>�33ᙙ�Ro�㻤p��st��r7wI]��Ksr"8�\��9E+�.��]���DW6�G:㫗K�;���ݨ�ME�v7w[�.W-�s�s��*���nU��iw\�$b���w]��h�7"f�sEsnn��mwu̚�.nv�뮹��9��n�M:�Qݺ�9\�vܮlm�.]-��u��ss�r�1�vӮ�Qͷ*f0�ܝu�tnAӻ�+�#���p�ιW#'�.�:W6��\��r��:v*�]wI�b�guF�-���b�*�N��˗9�ѺS���gv吣�sn��'v�(��F��:u�7:�u��;�7!�wtnk���K�rˮ�Y�&����ܳ���#�]ر8q,9k2J��tVN��������x�؝z�уk�ԟ�w�ʲV'�V�ӱ�
M[���uj�iGS�y
0b^�^�gְ�mJ��;gG/���c��6_�3�&���v���зURͪ��Gp2T����ާb���M���}���mHz��gO+<s�|�y��@��g\V޳�=u���>J�|���g�Q�d�W�/k���Z���X��W!��U��\Og�g�޷9$Ō1�{�T�5����;�2�T.�Tm�1����E��\G���ep�m���ݵ����ѭmybݵ垔���^������ˁK�ʰl=7Ӂ�u{��ӑ_��//����=Bn�cX����ލ���h�}����T�>�p���oz@(������VW9�}���W4��Uk(;�|{�_�^�,U5�c!��\s�U�V~�{�qߧ8׎D?����	�{�`����Iz��;�S�t_����X�ې�|��������*�![����7�]�������4��~�~�$߸�vP�#�����@��`LF'hj�v@�u�ҽ]X=���J�����y�-%���n��Y�R�1�k�;P�rW�T8,�tF'O�k�Q��7�W��8�$�_2GR��L�s��+#��:2���.�hg/�T;�|rHH\NQ��Z�+�!�N9��r+�ђTL<��q�HC��\�%���
�u�4�$����͡��Q�W�/hY���X*D���eI:6R�,��8�)]Ѵ?+��o����g��?w=�
�$��Z5�P��7�3y�0،��ڣr%�����i����${��/���r���K���NI{P$���'�ʡ�T�s����2��7y�U�x�׳\f��w_x���8�9�Y��~Pz�ǲτ�n	��1�M�����)Y��`V�c��Z�ȶ��n[�<3�����G)>;q����v�<�z���痔]����y�*�p�@���=��X�]Z8)�v�A��w}�� ���c�fOן���<ֹ%-Fo#��VI���D@j.
u�d==�&�[��O���{�ո�w����fL{c��ū�����]ՠ_α�S����2KF�f��7E��_�����l���b]`�ݥ���^�<���dq� o18�e�6곪b���#M�{^u/����Y��p�7V���_�#��Ǖ�n���ɿ�����ꇷ�Y�u����
4��΁���.�Hw�Q���s�!_��:� i+ˇ��]���]&��;q�C��0�oH%A�7���*zj�B�=��^a�c�/z{������o��@8�BΑwzu���{�=Z;�Y��#YX0��O�>X5Ӭ�wC޾��i�`�voAX���Jz�t��Ԅ�mY�}Z=S��xV$^a�_A[�p�G{!�˶�涤�U�[���\�}+���ω��P�eU�=��dg�1ߕ�~O�]V~����JX��=]��(�_��g���X	o�W���!_����ӟ��0�_m�����9�r�>��������ۍz��nO&������>'����wYU�t_�,i�����_�N�B�&�N�ߛ��2���R"m�~�[Ee���vr�B������r&/uL�3io��_o���z��k�3�辸�*yTg�9�1�s�<�N�%�Ψ%��b7=g��Y��/��^gg����}JG�o�9�/4�@�}g���{����� ��{+M3H�Wv�m[��u\�պ7��k�y���q*�\UO'9nh9����(c��}��s���.��;�4G����Y�s�K$���(��g@��"˖��L��"-��q-��g?W2�ʏ��':���ي�:�w��z3�4{�u�����f�:�1�&t Ҹ�����Q.[X�޳�`�h\��u�{>Vp��\��i7�}wlU��鸆@树�`�P#K���+�>_��π���t�k���?�r@����og��SZ�W���b��;�ڶ�5�����ykY���aظ��3�z����6�ZW`��c��XxP����fܰY��{��������Ԛ{�p7��=.��:���/o=�w�Kw�$�WG>��}�9���:v��w^�uVq��URX�RZ�$���B����9�}/6�W�_fZt>��q�{���o��<r:g8�ϙ�O�8�����I~F�Q��Ni�{}���������V�x�ǥ��zd=��wF}FJ���7���F� 9���޸�;˽.�V��۫~��ts��v؝������j�,z���1�u��}A�����i�>�k-״o��5{�^���I�8�&wFN���>�q]^��{۴ǅ{/-��Uț������q�D���ẽj�p�=��̏j��P�ޠO����|}�u����|n<_q�Ӎ���ӏ7jk^�˾��g|OGup\sz����v���+�|��=2��ǧ��eW��7�n&ĝ�^���x�I��6y��8�\<�SK�/�Y^��ƬZ�^��U灆���\O7�
C_�ȧ��uO��WH�7��*�w�WZ�"__q^��.=��z�_���5b�X�nݛ�5�}N��7�I�t��
<3��n"��U��^��lVGuw�]Hrۘ��yY9�>�2.����C�@��C��3n3����ڼ��3�[9�]	]lRXF��ik���FW�,�>1�\}2��N8m�����+���}�!�W��k-�7��u�'0�Z�Eu�wm�[��j�kvڇ'u$��LT���n�!��D��\�q=��~�+�m郴@>�2������O���a�����g�(}�U<�(<�7��r�Y���:�N�Zr"_��}R��(���l�a�Q�����7����{Y!��^=��奢�wm��w�H����F����9������l��c��6<���Мn�c����z�n_ZG���;���wQ�uճW������jm���U��>���Pex�\�ݞ�
�_b����lÎ��l�:g|OwTO����URϦ�lV��!�cWj�`]��� ��B�w�� 
�m�w�j�1�<���q��q��	v�c�����ּ��7��ԎG���=s�?��-zj�,w��oͫ��n���ל�s�Ӕ��T��bT�]r�C7�F]Y�v�#`�?A�M�������5�]���t��u��^I����{zǶny�ﻝ ��p<�9��躁�Նe@����p9��DQ~=��[2�E���7VϮԅ��g�/.<�Ui^}@t�κbw#��j�3^ޠ
5���z|�r���~��{9�{�x�k��k�r��f��D1������HQ������;���{z�������Z[���b��N�l�(�y�y�@��J��%�23���!�B���*��]={9�3��I���*ݢr�h��o�]��a	k+-�[͘67WG[�S::gu���=)���{q�
��Lg��E.>��?~���������}>�P�D��e�]��̺|6M��ղ����܆1U'�2"_^���5�W�޵��X���]�կ��)O����a�١�ОE��>>����=L	�N�!O.��u�һ+6=�9oj�4�􎡖z5�1q�{t�Y�R�0���>��F��_�P�����3�tc�Pn�����ձ��rk���k+���6;�܅�r�(��ό�� �2�:����V�=���kNߝ��������s�t�/���r"���K���l�KeJٝ~���
�!y��ܷޟ����~��^�r���7��szG���|��+���8��,� '��UU���?N�!��g�*t�wTĒ��~���n%�C��[Gܤ������wlË�ür�>�c�,6�ǡA�|d��_(�SP��ף�}=��Ϗf���n��o�   5�E��x��zƸ�9T�+��Գh�������7E��`�j�nHb�>v���ܸ��[{5��]y���VZ����Fh$V������`G� �q�7$��v`E�}�I���<����,���>�R�r�[���f��)sS�f�&����A,Y�G�r�甩ȲY��n��[��y���3�}WQ#�jl��ކ�~�=��+�����VvE9��|��Ѹ$i�/k��zr���u<"�v�Mx����������]�.�G���8� 7�������gT�<��͊�{^�^����ۯ�cG������$��5$���g��I��7�̌��#���s�nx%P�mXF/�k�����ɴpuo��_��~5����ϒ�c#Ϣ�M�Kn;���7�x͟f���D��U�s��*һ�Mw�e~T�[ts�
���@-Y/���޿��?�F}��NG�k���'_W.����f�m����)�UY���xO�a�Օ�o�s�}q� ���aL��'�Ȇ�:x���G�u�
��fz��ˎb�دW�:'&�QU�Y���N����< 8��i��6qᫍ��h�U�w�N�#:���=�:7{աǹ��Ys��뉗���B���MM�M�[���%ީ=�=g���Ǩ
��qꮨ�;=�����"�}jI*�e��m�"pI÷O=y�+:�h����L\Et��~s\^i�X��G#�{��u��#oei�w.7˶��X�Z��t���t(V�?�Vh8�7�۫*�� ��:��A���8�;�(.i�:n녛I[�N{��ޭ���C's���J7�� [X�7�Wֱ��_0�B�w(��ju�xP\�Ofwn�lͮ��{o�7z�5	N�z{���A��E@�	=(z*��9nh9����(gDv�go��v��6��^��x�8��1��G��I�:�)(��d�l[y�"����3����S��:��
���g���Tx�Z���N��ᾩ�pȀ�A����
�����N.ډ�����=g���:�K����wϫF�������}3=;�9�A#L�[�e�����9ǻ�k��Ѫ�A��<�P�!���t�i�>���7�נt��C��,Z�-M�ξ	�|�&�o_��sY)u
�xpg@=Ʊi���u��<r:g8�ϙ�Q�8�:��5"�;��b(���u�*�R�/�[��{?�ޟ�:���{z�;�����Y�p�z�3Q��R4�V����*��H��+ \�R�-�M~�/�����39�<2��Hž��F%>0��gJ�q�^W�� ֫�g������FQ�W��kҟ�c>�ۛLxW���݉��O�e�o�o��[O�ys���uXs��d{av{(foP'�D{�b����O��&�Y�����e���%(UB��U��!,m���_�0�{�Mɫ@��Q�N>X��au��ͱZۣ;�'����#�g4;"�bVd���P.�ԧhDc�>�D��W�|N�!��	+��Z�]8�7̰tǴ�Gqd_3��D*��%`��Ӻ�=��՞����Ϊ���u�qϷ��J�v���Q�B����eᨃ������'ލ��OwB��U�-����M\vD:�\@ȗլ�Gw�5d*����=�	Ñ{�!{�Y�#s;_���3�>'d�z)�J|8�.�Tj�\`��u�]����1뎬��:��s������i賄�pg�@:Xʙ�n)�e\x�Y����1��wOqٌk}��8s�f��co��{L\.{u�,�J�1�ѕLI)}U<ȷty���m�2���Իi[��gܺ�[p���9��R o�Y�Q%���0yT;�-���P\j�����	���׾�K�N�x{�G9܎�!��*���|; l�K�r Nj$��������{c�^�et��(��޸��n�!��Wt���#6:�٧�"x�C�m�?N�Q���9܂^X��@���b��{MDb���_[f3�6�>���7�q;q�wƄ����ia����V��x}��*�5A`.SBY���mH{	���t��:g̖f��T�֕řs3�9�Q4D0���p��6��͸�ҡ���g#{Ga���+�ڿ��3��\)���w�Ί��JKX�vс�s�F=�o�=CM=� Z�N�:8@w�o՘O����]���G!���(���/`G�x�W3��!+��c{)e���׿?���EG-�;f+�{]F�(��;|��b�m]н��cV�-��u���g�/���7��7�F\
]��n�y�Q�������1װ� %xV�lO~H�X����Ϫ��wPn;�����sC�U��;)u=�Y��O��(����a{�ou.g�O0v������5�ˎ���������T�>�롶���oz@(�<6���Vpܰ����u�Օ��{����f���!T�i���)q�uW	Y�~���9Ƽ_�C�T��>��׮B�^7�����CҚ�pG�x�����+�~UI��׬�wMqԬæ�7�N��W�=���i�(��ʦP�s?|fA�X�d׍�9���`O؝�B�]p!-�]r�����������4��9�Ճ�r!=�.=�n�ȋ8J@ó�v��L�� 5~5C�R߷G��)W��]���F&C��׾����z���~�;��BW(��IhѕP�(�#ہ��^�z���b�p/}j�v�����8�v�wl���pY/փφϤ��(UL�
>� ���=�iq`{[
��A՝:Z��BWk�82K�D�A��2%��s#,��:���2q����#ʞ��6�F�b�_��\[a��`�e�g�Y}�O/���Z.Q0����ft������&�Z�Z+x��� �Ȯ|i�W��D�	�)�6�J�[�Ѯ5�X�07��-C{.;�n����o/�a����O{3(4�b/��z�%:[ ��n��;�hpS:1�@�J��B}���TJhm���2�rh"�5>=#W��˰sL[ϖ@|��>jQW�b��d[�־ȞL'�l���R����}����.�JZ8���Rg,4�Ȕ�v����^��i�;�kK$`�x~��ias0]yh;�ѰQ�*aw饟x�
KG��t髬�ۑqT9]cj�i9�㨨;\嵤�|Og$ޯ�D�@ �W�ґQ��2�R!I��|�5��w<4&m�1�_�Sj>�a��*9���NW��t6J+��]
rp�:���c�:��I��ZiX�]�����W$������\��;|��l"����Bv�U������!����VnC����ϵ$��.�ͻH��}��32WE)E���c��k�읡[�=T�`��y�\�(V�ؠ���;).�F�h�No8]&{�8��^=�{��i�3 �烈w5:�e�Va��S��T�Ɲ]ѕG�^����FM�e��*�z�T�|�������W@���x���a]�}Iu"�@n�3�I�
Cx�w� {��L�%/�v[~�
�H��)�{���K���z�+�*9��D,�G�f��߸�I6�q��#�i���+����Cͨ]ƛ�^�'r�HsZ�K�Љ�bH�1�1��->\Z�*�CA13=s&�Ŏ5�[/.�7�2�굍͒��u:���\}p��{4k��Ƿ|�te�9�Ҷ���C�nnm�8һX�����-�/�z/ �W���m�'v��wx1��Dt�G�L�<�xfpr{��ŧ�vҫ�+vR�O�(׾�l�7b�	����ll*�ٌY�����v�Nҩ!�8d�9O(�L*e|��Io�Y&�[P1�Y���|*�i�Ti5�,P�ӖV�g�:6�=ڼ����>�P�1�O*�c��r�*�����xr��)b��t�ɉ_��ݫ9fqJ_�7^s���s�)�42��RsT��ᶮ����D9�wg��xT��īw�!��K�[3��1�Mw�q��2��,�/��Z���k4֧N���<=ٹ1+/������7�2o_m"IE)��
�m:ua �j/2�sB�Kv���^��uHG��f����a]��GoY�4�+�[�sh��"��	7���B�\�/՞��z�u�vz�w7K�nlax[�:��2�N�h��e���gh�$3Ye|ϴC|Ĭ�rvzӞ/v m��j�wx�c�j�Mu�Y*�L:*���4��ع�����!��h������W""�q�N�G:�w;\����w\wN�\���\���FFRs��S��#�u�t��M�wu��p�J:v�ỹ�N��].n�������(�)ݹd�&:I�ۻ����9��W9�We���华��\��;�����iˮwu����\�u۫�\��-.r;�F�E\���s\�ܑ��b��̖���Iȹ�nA�N�n�(��tS�؋�H-����wt��l�qD���r#q�1�������]�Th��m�N��؂��+�th��sh�K��#r#��Lnp��\�sr�B�s�2�]�np-ȹGw�ùwQN�r�����'wk���f�{9c~��G�>�V�GXU�-�����p<Ե�\?r����*[���;�tnB�����U�����z�:PR��tp����ڂ.S?���3~n��x�/��v�go����q�ӂY���VГ��>��X��G^^�*�́0=>�o�.*e>��n�&�[�<Χ��r���Prc�D����WN��ٞ�qv:p���ϏG�������k 6��ף�D�;cf��CF���{���KV��d�C�q>6��✙�|���	@];FC�ؾbې���3R��t���O��j��+���2{8�M��ՠ\ugdS����2KF�$i������*�s=|..�Un��{P�G��ơ�*�*;��=�k���x
}��۪Ω�I�;f��aIY�y]mRB�ek�]R������>Օ~m�Ѹ��&M�u���\oP�+�u���.q=A���yo�|j��Z�>�l{�N��w���LUǥ�ו��ϡ.�F<�'��Η �uH�pT��/t{;dzk/Wyh�<$�=�	q����S�>N|O�҇W����呑��O/y}��w�j[~��3|��i�}��Û�	̅Wk�/�w���/ #����`����Ty<TV]�yk�劎��*�����.��wc���55s�3��Шk��U�&�Se�*���0#3��h"�2��v��;6�%IhE6�h5�=jƞ�Ii]�*�ի����I*�1�:�dPɑ���*,�I wn�}��)z.�]I9��ڧ�F�x%g���_��
�Yts�Jv�=��3c��5������/ ��d9�L����>�� �v��[EQ�P�]��;P��5���ꐼ�6p6��-�}Շ��*3~=W�P��=N�㸬�W܈����u�PϭI%SbN��2}`���l{��R:d��3�늙�1qNBs�g������.�wOqY\�9d^E��"�s.=5����ub�I�^=�� �3�O��,]J�/���-�7����z:X��Y�yʩʭ����9�x�є7�o�=^������$�t��z[2J���	��}{/qT�n5�����es�>*� |m���d@�T�D��l	-�vWPa����c�bb��_=����G�tI֭��\��;�F�q�q�v�[��d�j	d�P7��䐢�d������o
抮�0��v��O������};^㻯@��^��T�-T���ц�/w$�V,��ׅI\pdʌZj�j���Ȟ/�s��k�T>��-~��lW����pS �!�`Z�S��Oxz������g�_t��'[hHo-߁�T���δ�UM�(H�=��>һL��j~w��j׽�Ҕ��3&<�]�{J��3a���ن�J��#�u&�j'OS��Q�cU�ؼ�t�|�=}`��V����dVs���#v6hd��4.+�x��_���C�m]ыm��/�@�nڹN����g����#�c���C�Eg����`���,�Q�=Q�w�����_?=!���E��-/?=���J�)� }�~�(k�H՗��`�{��ڼHW�G�Ho�_�nm1�;��C���ǻ����	����C��SG=�C��M>��顷��C3z�>�pr#ޘ{Y\����Z��x��ѳv���|t&z=���|����n�.*~��y���'g�~Z�5�c��5�� ���W�]����gg:�M���Q|J7..U�gx�S�g{���к��t�%���w�M��^O�5�Z���C ��gC����t�r��`*�p+�]k��}}�O]Fx"SR��Ц�{u?b�Z0�ю�v��9g	J�2�P3����F��!�x�Y.�
��[c�Ԁy�H�+²��̈́�م�7���,.��\>{u�"�$�c�KS)����E��ùX�	e<�R�ߧ7��n��'��v�o��c����C}RͲ�.���Ts�FW�FS���z����ԬH�h������@��M�=)�R�2X�
NS.�qItk4�c-��*�B�֫1�7O��ه�Ȇ�7���TǅG;B+��,�r����q�rr���#��۝t�Ìjĝ�"� s��r�Ӣnv�j�]K}I#�]����r�I6/q+��.�Y���5����_x�ˤs�Ȏ�!��)����8��)�蓠ʵt���=Y�w׾]eo@�r��<V��O�rݤC7�x��>;q��G�:�٫��P�=�}�I?MY��Z�����G�.Fm@�.�*Ӹ��<��ٌ�ٶ��L���w\N�v�\_{�9BZQl�_t�����D�c}�\	d�Жw�l@<}�nC���c:yY�4e{�J�O�����vb�����d��j=�]���S]F��X�������k��W!�<����_k�.Zv.WP�}���3�oc7�]@�]��%�?@�=4k>e!�}�"c;��v�gyU߷����=�{�z3���c���u�{"��ތ���ʁA���Ӂ�uXt�O_�h����g����w��^\<�W]��}@t��κbw;���.�雸�� �kr䯷}��q�r�J/�g|2t;����~'���q�e���U5�c"��>�uW	Y��׾!��b*��V/{K��[g������8�%����yG���>�K/���U'���;�zq��W�[��[��5���j���9h<O��1VV�{�
��F-& ����2�Mx��1Y���X����``��Ǚ5��l����w9@WuhSV���Ev�Ƃ]��!NES:*m�]`��O��ݙ�R�8�.��2��r�c�8�r>�=��t�O���T�&v������Y�Vk�c�ǩ���M��t�1Y�߽�����K#/��=I9^���ӝ�H_���9g	J���_ڇq]T��W����+��syu�ǭ{�w���8�Q���MWO��u�����sې��J;%�
�{E�j����f\%�gԧz����G�W�����{�q~ϻn;��s�"_���Iw�	*G{��.�*��\���A�W�2I��tT�L�2��Ϸ�qzs�K;}�p�W���uo�3@�&��I������?e������nbIO�ŷ^rݡ��u==���HT�� vb����G��]��;�,�C�u�6Al�Ger�����ף��tå��#Vt��C��v�v|��ް���I��\O��u�\S�2��@�N�Ȋ/O{ L5Ghi� ���Z�yU?o���P��2u"{�������:o�)��T�FIh�4���^�f�o�Z曍�{�9i���r3�6���t�y� o18�}��۪Ω��L�S���6���h��Q����K�'D�-��:�Gg/W�����)X���lD�Om�c���#��+�+2���n�n��N��3V�]:�**�
��R�dAS.�V�����jU�Ol	2�-외���C�3e��F�Y쀪��H�����������5��\6�U�W&�����ꇮ7�a:�@��ֽ޺�k����E�G��'p����W�~>UuЗ]���]&�:\��B���𜼙���Z$���<f;�J�1�=>~������_��UXcګ�E�R�5ۑ���N]y-���˔����eg��i��g�����	���ݟPY��*���W�yX� S.i\���ꔽcr�GGU+�{�������S������k��l���C�mx��u�[���/�s��^C�}�'��ږ ���ȿ�:\F:���d�Իm�:�+.p�l�y��4?q+��sFse.��Of��@�|���
��q�����er���s�c���P&�=5p'I�}ԧ�l׼/�>&��C�*g���9	�ǜ����}���tr;����Q�G����:���0_�sں|����K�u9y��O��X��H]T�s�[�o�>����f��i����]gK�y�%�p�f��p�>.��; o�Y��D�Ft	/��ْP]M�	��4T��ʕoƍ�֌R݂�~*X�<�=�0��=�W������n���J����gg:}�U����u�����YBY]�8��':�Р�Y�aH�|bj��w^�89N�+l۴�����C�Bv �~P�d+V���FC��c����}-
��n��w�^�I"=��5�w��q�H}}q�}S���1�$�@+��m]�j\�<���X:��+��|����uh�n#��#o�튷�S�l�9�OH�̔ꕑ�^�Z�}��"��]A���]�}m����=��;^�����5�uU%�=�<��t��x)����7�R �=�®*^�g��5�MC�M_Q��O"x�7��k�{5��W����p����Z���H��s�y̐���=;ƅ�J����oT�pڻ��o���!�E�&�s��o���+y��E.���z�߅�r��b���`�~_����3���J��~�~�yB���ޯ7�E����9�}<�]�^7���^�Ȍl�z�㿵�kG��2(�r� s��[WW�*��y��a�]1��M��f�Ý��#����P�ޠO� ��z��qίdT�HMv)V�mYΟuQ�ȟ��}���L��)Og���J�z�lC�Q�)�>>��(Q"�=�.��or�s=XzN�u�^7Gx�|:�r���bS�ez;�q�"^�Q��r'y"�0{ �1w�W@�Xv3�g^g8��\m���^Um!ag����L���}q��'�0b�	��VQ�h�����F��]4��$<�K�u���A��EU��G�-,7Hd�a���v.�84\Pu�-�j��'��N�]ǌ���
�C����8�9�<2�·qR��]9����#��
�]k�������]����y�jH�D�e�״�{��#�E�%+�2�@:X�yd3���
��.L/w��9j�=��3u����Y]HrȂ���s�Og���U������]�6��ˮZ�b*Ns��;����"����=׃";D�>ϻh���lv��~�nL���$�c`_ǕC�sj�0'Ƿ�����*u՞��P��}뉸�n��"H�;�$?�U#���v|6}%�9 ')�ޞW�g)���>��^y����P=>f⌳�r/����ݤC7�x���O��FwY��t�j��A����iC|m_lm�)�B|z!��@��.��:�P�N�-�"_[f2 �m�x�#�~�M�X�Ε���;���3����?smZ��|C|P��g���q�ٽ����wՍ�~����[��Ko�w�=����&2��u�_Φ����Hj�혩{]F��;���1>0��:�~+��`���t.;�q=����x�u!v_Q@���������VJ��yhs�@�i�d�mhR�L�^�����_�s�������%1�	\M��*����Tl���6�\e���6X����c)�Ot6��@/� ���8�$��� �j�Z�2��b���|����Y��\��Xn
��ݼ����]���'M�զ���ۧ��3y���m�ѿ�� �������^�e�]6fW�������
m�.^������>�������9��ײ���ں��>�:NuK�롶���n5���Y�/�U<D�Zھ ��&z���;�V��~���a�~�yv�v��o���uW	OGs+�f���;7�i�������'?D�C����}J�K~���cRy`�76��V]��sn����y��:���^1ӿ3�}�0��,N��9�����Ccswru��I�-u���D�wt�WViϻ���sۤs�8JVf�;PM�wF���w��[��z�����t���>�_WY]hpY/օ����,��D�j$�Y����}�>��V��^��t_Q�x�Q����T�����r#�#��v�w)Ȋ�\K�����,�p��j��E>��U~G���I�}3`Hݨ�%�Ǣ��3L�3���szG�;d��w��מ\�sh���l8�9�g�Y�p@]Ft	
P471qS)��^Kv��'�	�w&5$�g��A�뺹�����z�y�p���㒀�ɔ�q��7�s;��yQ\ۖ��9K�o8zE+r�׮��\��kc=8�c��9X���\k,β�.1PYف����f�������E�}]S�X�)I�;�׸��rT�28�]�j����񇃽S��p@N�� �@����5���.�P�!�fϙ��+Һơ�\�AY������n#���}w�n����D���J��7E��+L��
;���^�;����(���k�vHA�t�=ԉ��8=�>c�;"��U]Sh�-$idc�ɥ[���U5���=s�����G\Cj��wJ�K y�5�*!�_p곪b��\�y_dݛ���Ҭ�_�y��f�o�G>�����>m�Ѽr��=� {�uCΡ�w��{]�V��,I�X=*s�r�����+ڣ�?��ϐ4����~%�����?�ڼ������̫={������2w�0�eo�'��{�c��a���	�:�O�%_��qO�h������::���\�'9��+>�\V�}��üA9�f9P�xú��7������3=.��ҽɧ�8�� ����T�A�n�t����9���^�ܴ�� �������LG���寴£�f�g|H�G����VE���qg����� �v���D���%�UWv���B���te~oj,�zg*;���9���~n�[ĩe��@��L��l�R��Tz3TZ�h����̧�����rrĮ{��Sk%Ʒ��U�Z�1da�˃4,*Lo-���d��ǦWG[nԘ�)��^nr�CVg���9b*���T�Q�٠(�>1ޚ֫�&kV�Z�d���!���&4�$������f�{GB]���qB+̙�Z����ЋGH��[���=P<Fk��ˇ����_W=����
�4�7YZ&lN9<%�}��	�񻹺�{F(����g�r��
D�%E����R�5e�0��r��r��+��x(�];5��ԃ��nƉ�i�)N:{���֫�ArV�� �S�L.�٢Q�	���ӛc�<���oKEQ��Ӫ�w�"5P�΃�o��cxu=�S78�MGcmYs�����
�V��f�r�:?@�:��ާ�����)AXs^�ݔA\�ڧ�]��GB�Ow7EcA��b�IΫ�L�r�&uFp���q͹r��rStɛ�B��Q�om�-5��@�okT�t�i�8��ݹ�&u�̕w����V����/Gڝe�v����9�_�����-[C:b(�ҩw;
�#'k3��:�c8�F0e���&kt��"[qnd�k%�L��A��0�F��MS�c��
���=�q*wk�	���]����3d!k�m�oz�S���PJW���΅���E��%���2h��LB���b<OF��+��eh��v��3��sY0��yp��TA��y����z��p�:�6et��t\�<v�9˖�q&��y��L.wvyV�!��.�#8[�n��e!N��2�]qe��	Gqi��V;�oA[ t�q]aC6)�m0�u:7�ZZ�0t�Z�����Xpͽ������S�͜�򩱗��s�EhS
 Թ�>����Iz��̨�w"�9ͻ����$+��n�m�2KoT�9Z�}[�l5�c5�X� oT� �%����4�kE�,�7���**u�(�8o^*�SQ�ó���l��oB�WY�M(fY��E��_�S�{�bI������[j��9�N�B��bW�ܽ6�"��o}�$��w�]%��8M{�56R*�w9<�FR�ۮ􇵽{��蚲�J,�Y��J�٢�9���]�g$L�3��ӚsA��<���7��B��:mF�$�]�C����4N��:�e��
`⻒�O@x ۖmq㍹���d�w����Y���gH]u�YOܭ�S�֘m��i'���L֗UӭP�}soU,��}C1xi�Y��;��7`zz���!>��iΗ��Kr��q`��^dl�,P��AKW0c�$�)X����,cFt��-7\)�x6����fvm� �E+�!w��5ΎC���╌��E�ٽ=��ԣ@��:�<N���]���`���Y����D�uwC�����������AK����R8s�������u��F#.��Mwv����ۛp��mp	�lb8	��r�.]�F��Ή\��sN�6;��r��WI���v$�����9]�1�\�r���ڻ���W#��c\��廛����i�B�nnp6��9�s��#uݨ븫�;�r�4��uڂ�]��QG.cp�N�;����sFJ�ut��G湲]wlr���\-λ��rs�,���"��$�N� �����K�����\�5�ę�76�5�r����R�
lI��;�1��ܹ�nX��nH�Ү;���\���8��4�����nnl��˗]ۢcs��e�fb��X�7������������Q�;$������Z9Y�Q�(��Z�~�W�Zu+w�eLB�_hK3�f�}�S�s>Y%��Ӯ�xN+�I4���+l��|g�����?�s���Djt��z/�;�ϫ�Ƿ>���«[�L�~٭~=���će��������c�S����s\^i�_c�<]�◒ű�Sإ���g6��F�ޅ|z�����\s�RAU�A�X��HL�Nv-�7}�<�C:c�.	�>�v�ޭ���X�|��;p��v�9�9�K6�$�3�O��H���ٺ�At��뺈�&�zn}+70��f���bGJ��}��W��q�H�����O�D��l	-�w�|�q��+֬�8v�ƳX�n&���!�^W#���Ѥ��d{z�ث��S�p���PnNHx����GV
,#�n�N�u;N��P�>��GL���Ӏ�w^��7Ɯ��d���S�{j�b��%�I>��@ـ����z|=��X��;���}<��3�O3q"�0D��͐�<���ҏHrb��C��G��#���.w���^5z_�G��C����Iy��*��V������K4�fOD.�����z+z�*eu��9A�1�ׯ�>�=�W�c�)V�#������|���S����QC1:���y\��I����/-�.7]�hJ��r�	�ۮ�����ot�-�G!��gG��ji+���=vA��g#��W''XX/�Cv����g�V��;pJ�U� �z��u�������Z����}�2���]и��g��ˮ'�ޏT
��2U��{	��;������zfz��}\�o��,r���ʺCڪ�9��P�7�V����졙��}@��I���yT꩙���Ғ}]�+Y��'�Ǹ�{/m�UT������L�^��}��>X;��r�.�o�Or��^����xF��VUx��J5���\�;!���}>gTwz�Ui�tJ��g����5��ѧ�]9��'��<2�L�WS�|/�r9M��x��Z��}7J{ۆ4�Q���J��v���q�ϓ�f/������pe��t�qS<��9���{�ڲ���M�7���F.� �Ewϫ���C�9�0����Ȳ�(�s�*������� 9��tc1��_���}E����{t?����dv��}������iȗ�A���:�$�3y�����a�l�]x��d�9}�Q���X|s�o�q-�x�ˤs��������ti�-FQ�>׆{���).�yxxU=l	�@���(�9��q-�G����~����ߴZ/�W��7~6	i!y�Nf�8fջ���C}"��R�<7\te�v%�Ѧ:ә:䎖f�p�{�u!���%v�G_�A��Hܯ.^��X��#�gAx�"�wWOhӤ�9L��gh�ˏ�1t1U���}�CV���5>���wy���K;�i���t�ّ>=�(!��6�5��H��ŵ�侶�dͶ����'�;U�n�t���,���q;j���s3,�T����6`�h\E9�>��n-���9��v{���bع��)���>d��Q���*�Mu�2CPv���TQk�^^ɪ'��6�ՙy��=#�WG{�F���\6�������x
��e���}F�FI�l��l��ݪp!ۮ�Z:�Eo^�	��Tw�y?_��WF������<y4=qї�V��k6���]��K�M���Ǿ98:�+k�7G�^�ǲ����+�>�:M��t��uH�F�g�d�r�*��Uv���fWoP���pv����R�O���ײ���Ъk��|�E.+��;5I�d��K7��^�}�����5�� ���O������qJ���&2�rUnJz�������Z������gMq��޵���֖0��|fW�y/�ɯdX�1�ê���,Y>�������A��.��W����wm!q�{t�Y�R�0���v��t�8���y�T/H#H{�����m�gR��G�J5��}W�����۳k�j�f�e�t�����,]>�K�f"�S@��2�'�����ԭ�`�DwJ��z�{�D�ش��\�� *h�@`Ճ2fcQc�faZ����M��.
bY�:�uu�\�]�)�V�_�ƨpY=@W؝>����=Zޗ�B���Y��$�W�)��(!�����<t��\Q�����7�T�ϴ�vq^w�ٖ���~������/�-~dG�r�`_���1��ÕG]L�1'�3�晛�7}�F�/Nv�gsMw������y��(k�����/τ�p@N�΁0�j nb���O�-���[�<;�W�������zwΎu��>���>�>��f@�T��2�l�ger��X���Ou�β���)g���lX����ٶ���n�}��늷SR�Z$t��қ4a\�|�Ǯ�Zu��a�Fv�	�t�"{#��2{�|�gdUê��@��W��6;
:��~��,a�^�tWUǪ5�C�m_Q����=�Ƹ���x
��|� Fɩs�ض�z��V_�Ltd�푦�DOmxU��Q��^�������r��7�wP��h�x+�eI9�ݣ�"{±Ȳ;��9s�b�:P�c���	��?����/:\�]wu�0���,�8�N�싌���⼝��A�^�w:y*ܦ�`�m�:�j��SNc[�s��Z�I�l�xW=2Q�Z{�7`�3F�9"�����̧8.< t������g��8Egh+�1ه�S�߉���W="�Lr���ƪWL�)s�=7�Rm�];vI�}*�]t=q�C�l�JѓX�x;����ω��P��ո|jw;glj����t}ʚ��wP]9��k���]>��N���,��+�>�HW����j��s��~��>�q�v��`>�\ ��5Uu�9�u˧7��j�o*�vz�{>s�}���<5|Ƹ��t���)�tl�Ξ������VE�*�\FC��O��Ԃϗm�~�[E{#�]~o�4l��L���;y^��M�w�9����;��d8�Ǐ@^@��x�u��qY����w5?
�N���y���ǂ����DZ�J��aP���yL_��'7�5��i�Q��Gs��~[SR�w}�J��{�ܵQ��בzW�2�IT�$E�*P�T�s�nh9�F�22{����Ҽ�#��!ܣ��dGmv��v�|]{�v�K7�K�3�@H�g���ӝ�%�qNs=P��Y������{��lG?W2�Ië:�>6������{c`]���e���N�ҳ�����Ղai����n%��s���|<OG{�F��wlS��uބ�7��q��1��9�x�v��,��%a�2l���t#5]2���t���K��Z��q��5��s�+ܮoHly��b�k)�.�Ja�o����^�恵���Cy|U�˥{��^�o_b�Щ�=��)ח�6����=R��� ��/K��0��b�P�>��GL���Ӏ�Gw^�j�R����8�z�J5�ꪓ��Ijl�6Gu!W/O��>;�-5�W�nO"x�Q�Uz�C��>�m�v�-���K�f�.�d�u��Q$5�j�}.w�	���}�Rc���W�2��gg��{N��tc���2o�}={"��V� .��*(�j�;�*%�_�E9��˯Q�����I_�]��;Etw��xg�u�����wO uu��ތ�{,�V.a�x�^V���]\�P��P�~�ά=��n�7�y|3UW#�}C��M>���m��~Mm�?m��^���d�(�ɳU���P)G`�=�ͨS����||�^����9�u�q���ݹ��{h����9��]��9�Ew�����gp�>��^6�ap';�ϝM. ��v��%�q����߱5��OVO��|f~W�h��f�/�tk�8'��r��ŀ�#����j^J+��?:�y}�`w��i�﫲���^f��H�%+�,e|�b���FY�/A����Q�>�3��ɗUw�.Q��%�^�w��oD=�c��9b�&}73r{�f�%s'�L�r6�I��eu���-������VE#����Cf�Ʈ4����z�6���+�y��W��ZVc�M,J��R_^��k�=�=pF>lVwWqYԇ,�.��_��nx�I@�"
�=?_�8�n���:�DUJ�u#�Q���g��'��{����i�~�@�T��$�\[���zi>q�A�P:����詖4�`�蔯��.��w�H~*;ʤz�}wúw�Qy]�����5�2o�@d��>���l��e�"�z�o�n�8\����|v0LwI��nd%��T��i�]���BY�"�&@��7P(}(VD��b����l���{]T�d��o���O��;��|�}�nu�����p�Y�RCP@��Ж}� 1���ؤ�����i{|=="�u���g�}�>d�ϳ�)ɞ��2CWhD��k���{�Ay��J3��y��Oك���8{��b�wB�u��}�x���� �.�b쾣h�<��g���Q@t\�F���n+A/��g�~C�C�Y_pU�޾��8�@r��OC23�ї���ɯ���b��N]U%��񙾈�`�x�������?@�1�kʧ~'�G�P&�:��,<蝫ɨf�0l�����&��Q�B�e��dҤu�w�ؾ�=�L*���z��<���y[b�x�Q�NGt��ڗ�j���LՒrs"��^uF)%�?�����Y`�xX�U���ג���q��7_	�m�D�A�*�>kwVbή�ҽ�흡�����%%w���kç�1;��V��~�s��w�ц���7�j�އ�ۙ��B�,�Q�����	Y�XW��?�߿�8�|����Ń��81��O�X6/�o�=��WV��̷;�����g#�k��F����g���>'޲���/�|#��fs����M�~d��&�|뀟���E�����wN�M�����B��n�ȳ��;=5B'Eb:�Z_�=�������P��.�M�	��r.��N�t�t��WZD�Z�sې��{�N��g�����sk��g�a'Ǥ�vc�(�#t\��y�0�4�X�C+�m�r���\ݼ���/���{�=���)	+~��$5P�*e������E��f��w�9�#��o��g�,n�{�9j��l�f�9���]{�`��o����j nbIO�m��8�랷,��M�o[7�"=|�����'�o;��:�ه�<v�[ +��h�0'�����n�ݶwV"��ζ�|팃ٶ���n�w��|o����Գ" 5_	FDB�>�Vd�Vk�5����J�u����Yx���I7@��-"�Z�9�6�����d��*F��1�t'���vU�X�$N��7�.wڡܫ`�Zyn��!Q�h����Ff"�Vv����C�`��6���d�3�Ү����r�u�9�bY�`�Tg�_�`L~���C!��R=H��3������ugdU���O�F����2j�<�
��%� ���]F豓QP��4�C������@�}Ƹ���x��{\ϢW�m_��|��ѱ�X���r���e�o�?2��ϸ�������BUL�9\L�2	s.�]��/m��� +_ê��P�)���� ��V6pt����\*��K�+ˆ�@)e	X���Uy��CV��;0��Rz#:\��t=q����UD�jǫ���=��qN|O�X�e�7�-)���ywUa����������\e{�'���U�� {��(7�Qr��Ǵ�_fg�'�gO���t�}�.���UN�緧�d==���o��C���������3g��k𹞊��raT�V�����W 'W��!:���;�H,��htDL<p3��p�Vg�%�s�T@h����]>|�#�<*ʁ�;@W��g"\�gn-���Ƞq�W�ѯ}�i������Ƨ�tw�B*�XPN��S<�.��k��.�,��j�����E�^T�Eҷbw_�;��¼�����J��D��Ή��ő�8�_JF���N��x�����z���N�8"�����	��gi5��K&АL����R\UJ�QlԹk�f��f	�}�Ԥ2���:����`|��L��RtV��ah��~�xr���M�\wƙv����l�"��R���NL�Q�n�z�{O�y��������{���dv�gn;��n^���GI*�� �1�E��L���{.zw�̓�}o��Eķ�����ʼ�@��>��쁾�����M̪���w��?= ��: �|̈�D^����mb�r;��i���R6�:�ح����f~��*�ܵ��\�̀�G��w�x�z���X�����t�il�:v�:�Q��1���g�_����6�t:����
��SpH#�D�EJ���_Ŧ��ɫᦪ�a(���Գ׾�u%��H�z�i=�Ƽ�1�9]F��\����4.��+�.xf�Vצ�}խzV�#;�]ы����>�����G�P�B쮣h�*��혩{��/kދ���m��׹l�`�n�f.ӫrN���f�x�]q^7������sP�/���KΞ������!����G�=�����������sϨq����g;����\���)�)�F����=��<;t$�v��d�h��8��aʾ7��h�;�tMd�����۬D��[���͝"�H��ax����g���]��9��E�p��r�s\Ц���UZ���t��	zC9�!�z(�#��ŗ%c٢ҘL�d�6Dj#�%������ٮy�wr���Z�n�n��(�U�9�]����`'u4��~�����K�]^�p��w��?d~����c���ޱ�E,�h�F�"���p��u���t�*�\�hct�v%87��5b���ؚ�X�\�3J�̩YȘa<�]hz|���8������sf<��*ܫ��ٳ4LE�̮�k�0[\Օ���Q嗴$�v9�dY�m�w�w_�)��y��.��	xW�P�i���s�(�WlD����4m���3�yݒ(,	!t��!\)�	Yr�պ��F��wT������A�
g9����a㫌/jk���k�U7��W�ug�5xttxX��C�}�'���j��r��a��vYB`Y aݟ[vz}f�^L/�:dJ�ܣ5ܾ��2��<�;i�5y��be�W�����ň�H��N��.Gd�Z�q�I�vG��HT@�����jk���Y�c��ua���m��p�o�\}.{ۀ�D�o5w���WYD��t�Xk�~v�Qεh*Ί)��/Ut۟8�>��/MX*�D��s��|�^&��;��/R]L����������"L������V�t�뷘"�v*��UewG[G j���W+	��ㄭ��;D�9�U�o&�vG@l���\�}ZV�)��VZ�t��s�4�\t
�5ݻ-k3���sgw$]�HJ§y��tr�.tĊ���r
���u�Q�Ȁf�
�+i5��q{����m^�ם�@l�E=~�>Z㝝+Us9fE�������|)6p�ȃ����n^��w��%��o�ҧDg��H���4U� ����I��r�w3R�;,��i!�
+k�e�Ƽ�Lձbl��3M�2����d����)nR����\;]�|���4p�q&�̈I�M4���1��"?O˅^����C)�Ф������C�x�ݿiAs���BF���U�,�Nҡ�Ďm�'��@׽>cidG/���wi�a!��͹ϚI��%��30w]�S%�úf0��ơ�u>�'k:M���"��V9ۺ�UIa�3e�G���Yh����D�1N-��]�NN�i��`�͸�h/3�CO{:�TD0{o�ǹ��gd�.�{6�i�=Y����a��k)� �{{}� ���W�+yNnV`���8dSy�=I1O�Ј������ҫ��\�\u��!�{&�V8�h*�+��z����'*�^]��VX����bY�N˪+����,�T��,y�"^c�K䳧gM�g�
9ݗ����������M�t�&��Ѐ��N�]q�$Q˚鹫��f�J�E�Q��s�08��W
���a��9;��jLMΝخl��ر��Er��\�4]�E��n����܄�˦��F��s	���㺊�$��۳r�wWPW&��b����cFH��A&����*LL�JDF�$dfc��7';Gu�`���3�n����%$hw\;�D����.BEΒb�Id�23��G8wF� i1&�J($��θܣ��v%M;�ĢK��C���4�wD���"�� �0 �@$@Xć9Αs�+��؄dW.���r0̆I2#1�
L �	����F%�t���z����W����h��9���bp�s�Z�f�}���R�.�Ń�`�ˬC{�=o�����jT}��v�:v��	���sl�y\�&�a\}������9�s�q�uW	[�l�6�K�E����~�Ha=�;���`aʂ��|EeV����M�m��SI�<}cw^]zh�W`�UZ�����G���x~�~�p�O��?���r��̫�:EOQ�r9M����|�Ӭ���h�]b�FOu�=u����*�ψ@HhgZ�Q��������z�t�&���o�+���f�?���B{���*zP�_^F/��ȑ�������.������&c�f����Y�S?�~��ty������'��{��S�_��}Rϸuty��Ք{G��R�zI=�1P'��Tu�Q������sq+�9�s���!鿻ʣ�2wE�S����(���di�+��MI�!:R7Ft�9����ܷh_��qZd�<�*��;��뽽�˼iF��OkV�Ю����	�nE�� l70/�w���x���x�#�f�iɌ�㷷�e��=<ف�������Gw\N�]��Y�@j��ʾ�3o<'�V]�����͐��X���gI�[�;����^࣋h��6��5�Yz�Ѡ\����F9C��U��Fsor��9ZKY�v	ތ:>���B�Ch��ע�=�����͑�TpԵ���8r�xl���^�瘉���g^�t�gb��iEr����j�{a{��wg\�7�����Vx�tϙ7�uG�S�늷S]F�S$5p'�3#�\쓖q�*w��B��޺2/2k��ë�%r"��t/��q=�g��b� �ϲ�R쾢2��Cv!�K�0�"Ng��zԫ*�0"�(%��}�qڮ5��?�~۫�q�x9��Od4=*���14�VnϺօf����*���l�p;�)׼n(����b��y���ϼ���=�2�=�Ƚ�+�ּ�J�=�k�;����bRo��6�]V:S���װ�2<W�e�:�mAN�w\��5,f{��W��f9s�L�{��J���o�q_�99����C�3�����8_��m�2]W��㛌���\1��N�7��W��\uz7�x����A�&�w�P�6ߤ�2g=����}�G���<�;@�U˲K�gs��{Nwm!q�{t�&j���S]�����!��b4�œ�ψo�G��NW9�r��u�=�s��w��LɈ��R������H޹D�k�<�A��Q&{M�QP5�*�>���C+�;�;��G���Fa�ݨ1�6^eg<@��Tb�!u���4���Q`	7j�r�d�A�O���DQU�����5�C��a*ب�p_��xZW�Hk�LI�=nv�q>��3F��x`��s���ӯ���1^�l��/����X}Ya���/�'�J�k�P�!}=��og�zܠID���P�Q����r"��3~]}㷹΃v�;��{C8i�ˤ���WrW��@��m�@�
P5 �sS+�{�Fl��GՕ��-vg��'������#��m}�O��gT�}v�<�ީ�|���1� �@^�C4�.����j��>�et�f���^���j����պM����ꩉ��R͢ 5(n]�uSx*��^
<��7uN�k Lv�ې�|�O�}��d�wuh7���W!,GJ���s��l���I���G�:�7����Ʊi�v����ҁ�ƣ���;�S�y��W��d� w�_q�L"N�M
���b��9Gþިm��"�O��W�������|�4��d��7���}�BȮu��ND�
��
���p\R��W���U���2%��fw�zspek���،�r{��}��C��<cx�W���W�����J2��z.�_��[ٷ�;�}�t��ʫ{Ur�ȏ>��󦙝�7��Xr#zA>�9[;S�K8m�ǜ���_�R7x.��k�ү{�2O/�-lֽ�F7�6W]�Xh�i�(>��T�
W#1
O� ��ۻ���}h��j�y'fa�twv�����]\��dԺ��;��t��N��L��� �s���Yf�lW�C9���$��墾����ج-F����c!U;�r!��Ӽdv����p�=t=��]W�4jo���f˹�`�L�0����_M�a��̝�� .USԸ��U�Z�Dwz�Y�Õ��X��TQ�^��]����I�;�]>���	C�=��Y�uP!��>����
�Ը�kU雿E�\�|�%~����﫺�ې���u�PϬ�UL��L�w�L�r�g�~9�i����6�ک�پIk�wy�eQ���VEuGm�U�o�Ҵ�9jH*�3?ȱqR����|b�GZ��g+:���O^��w_��c��E���w�]xC��F�$��΁}�q��c�����ã)��a��&�i��a�[y� �Ճ~�s��v�e^u |m���d�H��>�ݣ�K��^����W��0}���|n�?���!��r;�����$1�F,A�F������@�_6�P #�2R�=)��0�����ԑdߊF{�)�&�auW����Y<��}�p���s3%�|�KSpHtM�R�x{>�Ŧa��2�s���ׯ �1�w�.�V�D�{}3�-�ܱsS���R:N�\t��g9�|1)!���S���~C]]��8>Y홽LA	�:��o��ǐ.�O�],׹FM�Kxp������f�2�p��"��%.���H�p%��Z�-��c���O�d���^��g��9]F��\@ڰY�4=��4��G��O��U=�K��y~ll��=�ꑷ������E������z)� R쮣p�r�;f*@��O�Og�*���:���Ld�j�b]wB�1�3�xl.��ޏT
]�d���DBHU��^�z�_G���]~5���?!��e�4�{i?����P�7�V����Cg/},���MmW�h��}�K�D{���¾��7�ƽ���D*��9��v������o��^Y��D�Dk���^��ST|^����eV����_ap&/{n�gr��s
���;����wۤ��Z�C���ڿ����;� ���������9��wX��bl��ʩ\�׼����:�5ԙ�_Sg{����u��^���'w~+��V�������j��z)?�1=�|��Xz��.�f�/���B[���u!��#�nE�$�m��|+ї�ٯ�;2z'O|g��I\}G�w�ty���gh�g��{q�lv����A�eW��hAV�A������L-�1�r�dY�m껭�6�\'T�i���ܒ�3�����;%2�Q��u�Mn@N�x�&�[2�.]��wZ�ͨq����{v�g�v��8.Y���[m+G�v��(�{��O3�Fs���/�Tl*ܓ��e=݈���?! q��C��)��aq�sq+�8�G9܎�!���]�y�أ�5�c��]g�z܀���L0'�ґ�3�q��Q;-�D>��������c�)�:9Ӧ�L�>���G����}>�����6`7P(�n^;���Qj����f$�ַ=-��}i��=�ldwO�M����w|h[��f���Hv���9��o������xw�K��T�ѩ�3�Vx�}�>d�wTz}��*���Q�2C]��|4��R;4�%	س�b�����^,=�W")-�pۮ'�8����ǀ��p)��UJ����Ff���j�h�+��F�%���n����.Oqʼ�~5������8�=���o��t<��LO{��Fb���n���
�ї�VIW ��6}8�������ᨌW�5u�5Y�Y�os��4�ymj�,��d�}(N�g�ޡ雽� �0�����+���*_���\{i�U�wlq�7����pd�'�w�q:�9�'z;���ߦ����A���>o��[
T?��G��5�����g��99wb�'��>]�.����Q��^,?�X���ґ�g���f4�� ��v�컬�>��x�fefz2WS�>���s��+V:&����h֓Q�X�eh��i��v��)V\ Ƿ֤��:i�ꌌP��Y��ۣ�l��&���e��!�*����9�t�S��)~+u�^^G��3��?P6�7�88��{�ttW���s���p�'hj�v@�u��{��5��H_��Hˠ�;"K��=T����xq&�3���C��o�r+����]Q���·���~2��br;����?|����=BI��n�����Q�-���;�<��p>s<�H�W<ٚ��X�=皷��
�p�y��W:A���U�^}r�%W�:r�rJS�WRg"��3bGDH��WF��|���Or����v�go��v�u�=�6|%��jH.�΁�n��/��j���뜾�=���g{3��{��7/�����z\r���r�>}U�9}}S��=3�o((��E�^����mlT�����n^��@(m}�މ�H"��ϫt��TN����[���ٔ�OZ�d���X���A�����^)��{X�$1B|����=�Ώ���#"��4Q��~˻5u����Ig���UN���Ѹ$i�=Ԩ�zs=a�Ŧa�&���wR��mߦy��OG�-�Y�G
�����YqxG$�F�w',U��)jA˨z�4u���oA:�����p���n����l�1Q���z���}&�Av������LB�w�NKY������]��ɭ���|�R�uv9���wɮ������/��3^u�Ϋ:�-L���͂�xW���^�Ly�s���?]MO%g�����y9�s���u�&��P�x�FG:�ҧ�cgD�^>O���P1���v��z�M��vC�=޼��5�tb�E97�����ޡ���@���x=���,р���e0�\���+��c8;�R��l���]��j�Y}#�\gM���������O�X��*~��5˱t�Y��7�y�'4¸��FY�9����cS�!��ӑ�4:T�k�j/�z�p��;�/3]{�PXp��c�x���Ux�\J��0�.W�U.#Wjwܱ�ц'���oJ��IO�u�F~]��_�עx �Y�B�����A��_��@U����N��q����i�Y}�GOT&w+��۟wn1q�u�Pȼ����X�:�L�r����ʮ2:�i��Az�x��a�q�Q���tr;����Qڋ�#o��9�� �x,Qa֜��F��\�1���k�L��=����4������c��Yۈ�w��u�a���;�K�� ��w<=�E^'�&pfڱg�F���T���ƗC��ƣ:�mε:��?b��@�o�Xŉ3�����ɠb�(q&������b�mC�3�V��gmz��o/Ȯ�I�g�E�J�޳��R:��xu���^٬�)].��l唓�K0P���cY�Z|.�u��XO>���Ao��1<���g�3��>���Ͻ��{*�o�Kk{pOM�}�c`L�A�l�T�?��뉸��!�^�5U����U֮ٯ����VS�����WG��­uT��d ��4��@�|Ud	���n�<�%��v|�_��z�O_z��ا��=(�:}8>둷u|j�uU%��T����6`.�*K�� v�J.јڞ�g�C;����Q�=�ϭ3���<s�q��8׀}7Ƈ�UuS$54;Ɓ��ͫ�����0k�4�3��U!�ͫ�1m���":g�od3Q��0�����r�jI��F��+�.X|{t�V�}[=�W���.�ۻ�c�f����7���ޏT��j2�˃/��k&}4������s�'�a\WW�n�����c½���}���ϼ��Κ},Ҳ+ ���ݺ���oE�\�=r.۠J�p4G�0�++�o�/���.;콶2!UWiS�tL�ߘ�s�/([�&��>�Bw<�<-�W��i�G���ʭ7W�~.���]s����P׾;'��n�T*�V5I�#n+#��������llK��~{���t�����^q�h�����7S��AP��	Y66��	�1c!�����%�2���
��3u���r���V����i:�����$��Sre�:"{�Y����׸��Nz�F?I��Ix[�O��p,
u5����U�i��f��z���b1��7�k����W���۟Gu�1~�H�% X��z�ٮ�y=�v��3���qW3A�������﫸�����ב���(�몗���ET��Ԫ���'��Y��p���FY=���0�4�^��O3��WY]lv����NV�r���C�Q=C�ީeI[c`L��`��3���F%}�x�s����]Wv�V�^5�$��!QﹺCK���Ϥ�r NjN�0�5���FQ|r-�\K��'b;����O�=�y)�姣���Gܤ��wQ�uղ�O��"�nu��*����뙹���f�VY������1��m��>�*#����]�%W�k�u=� 5�3+G��[�{�{��3~�SC�'�}� ��mHi� �t�ǉ�N�u������*���
�"�؟#o�7�VG ��	_�N�������ې�����n���`{~U��Z������km���Zֶ���jڷ��[mW�kZ���6ֵ���j�ֶ���k[o��Zֶ��U��m���Zֶߵmk[o�յ�m�m�k[n�Zֶ���m��Vֵ��������*�ֶ���kZ��[Z���{kZ���mkZ��b��L���9�<�� � ���{ϻ ���ç{��T�ժd�1��--c)��R�Jd ���m�Mkii2m�M����VV�l�U���e��fͪ�,� �{W[�Ͳ��6����D[6�m&ֵ��ۭ���j�Vժ���j�Y��[j�5V���=٭γ�f�G�9�5��ʬ��55��6�UZе�Z���m����c6�H���5��Z-cZ�6VQ�l��Zf����]��Y�  �q�J���p���8A@'Ct�@w���o^��@�5��*W{���;����1�J)���kl��is��ֶ�;� .@z��ۺ d�] ��}��Q@QK{k�Q@�QJ=ޜz(
�=�)E�E�8iE(�
=��R�}��ҫ�}ei�m��m��&喵.� ���g>�� RoY��� ��	�q^��� ������k�P��n���Y�̋��&ն��w|_Z�Vi�l�;n��������Q��W[Y�;����]/c����������n���ƯGt��5�뺭�u.��i�<w���ݭ{���R�Nnv1wu����>���e���w�n�A���^�]uٵ��w\���N��7n�Y���6��F��x�Y۪V��GQ���N���[u�ޞ�I�ݫ�;���+Y���R�ݷ��5}UJ���\��U�wu���^��ҽV����ww.�vz��R�֫u]�m{��U�����a�K�k��R����z�s��y��M�mݽǫV�u�mh,�4�wh�&fW| ���f���w�ܥ#�y�{ý�ky׸�^�-Z��z���{S[.{�*��W����9���<�E+^�[�w{�ksUU��{���^զ�cU�����Ӿ  {�ꛜ����^��n�{]��m���&��V]�m���۱���=�뮸�����{Mƫ{�{î�]E�c:��{�=����ֺ���Jm��i�r�X����  Z�^��-��kֲ�뮳��.�m�Q�{{zٳ�U���Yj�v� ���[�ˁ�-���-{\�#����[9�8F�w� ����',���|�� jݷzP�u��pw�ѽ�^h퀠6{{ν�ʰPz�����b�_      O@b�� b`   �)�IRUM0�C4�h O��J�&��@4ɡ��i�@�~�UJƀ   & S�	���#       ) �#Bi�!��$�S�����~Wߗ_��������7�f�9&�$�]�M���!INο�*"����^�"����hp@�؂
����G��0�@�("���������������z��`�B�A"����2a�'�*���D�H	HJ�(P�����Y�y���~��?����T��/�uִ��~�8?��:gzO��l��S�Hkq���~?.^c�;�u��k����o.�$rkð�a��5�ˤ�c�����*[Ie�����{lT4Zb"d�T���&��۰�j|��)���e�*�8Mc
�]7Z&�c畺��.�:�ӱV��ot:H�Ƣ�kC
6��#�Z��[�ݩh���KnD��ڸ�wf��2;�d%N����<��<�\���E�m���BS���R�;�Ak���IS�f��p�V�4�s"o@:�ګCn�&�%4f@.c�z��UAmX�5�\�QB3-�a�iHR�r���^\����q ��=������jZ�cݭ�[P+ݷ��.(�YM�[�+��t2��.���3�#t�U贕mAsX��'�^4��IaB+ѷ70�aw�Px4��״.�L5U��x�.�0K	]8p�զ3U���>	��]�t�7��ƀ�&K#��b:���؆[�FB�;�E�
oZ8�A,���n����à��k2*HՔ��,b(eak��Y��Иr^�V춍$�̹���!V�IU���4�L�.�Y݋�L`��%Z:���̔�Hxt*] 0��3r���Z�����&�Zb�F�)ؗ�]J�gk*�*��m�8�SFJ��MӦoSe<�Ô���i�2!m�V��/"իsn�+�.d�oB��p�+q�N[Cp�5e�[6�*��T�C�[�ᱏ%�(S�b.����v�6$��!�ѹ�/�_a(nfD�R� �-=q��4�V��k�"�m�V�kW���Z� [�����Zil�S3Kx��N�nbP˫5�%�ۈ���q�
8n��l�5����é���.)�P�f��e��Iq�{�MCǘ��DK�ũq��;)��خ��Z;1@�=E�R ǎ�U�É����D�V��t�d�A��7i��!.ܷ��N�%���t(�o`�'9�Zd:Wr�
ʧ6(qâ�7q4�j�ɺ�+�����
��RKaU3i��!��p-qc�&�АM�BbBzE9w*�NG�F�6H�q��l���N�˨�[P���;��ZH�[���U�.�z��fl.�i���*/q]�U,�Do������*U�m�4��ĝ1q�چ�༕�ECu�IGÚ(肥�%�M�,u&�F˛�/�t�F�8-���JY �p˧n�=�D�7���t�6n�54k$�%�dO)%4ʲHN�NKWM�JU�����K�2�|H-2/r��}j�N���b�3S$�kFb�����SQ�VS�*�hi뛉] X;���:r�bA�tWƞJ4�p*���+^e*Mn�zBBՌo{��-�69�m��n*$B�Vӛ�R������!7����2��V�����Ei��t���mv+p����	n8�ܸ�K*�E�B),�NE�$��cw��i�Փ�1�7D6�x%���Yp21�wcA�j��؅JZ�$,�tr8���9�����&��e�̺����:���5e۫ �/2�5I2)6�S�V��nL҄��R�)TXNT�S]�B�V�Y�1�Ă��%f5v�4u�(�Z�Re�����fX���KìF�h���%��m�SIPZ.5�s	.�M�V(��~�d�A�Td��4c_Ć���T�B+n�Հ+p͵c	�%5��R���]�<�}�J901��E��Al�1P�:s$�J$f�u���YV�*��i�m��]���! ��v�\���t�Gi[ǋ1vk��
�[�a4M��.J�� 9W*ͥ[�h��5�pR�@Yp�n�gH�{���:�X�b�����.^]�(�X�gd�!�(�ݦ4k�M 0�!�Ġ+K��԰�1�C� �\9����m�\�%C^�۫{�V�&U�0�ä+�:Rd�Rb`�Oe���f *�-�4�j�<�LZ����S�y�6G����4�&sQ��*@lỦ�����b�/()cA��ƫ&���� 	ht�&�壳)Z�|��:@hɔejҰ:�Z5�iA Bi��жه�ݖ�}���؋Zw񗻔ޥC`�S(�0�ǖ2[+jE��f��hʏb�,˧Wӓ%4S�T5�op�ve����r�4�W��`j�i��s3^n��2�[��MA/������j2+> �P�陙lM�3Y��F�4Y�T�D�[f(�v��Вf���Kt2����J[�S�֕�E����+4�������"k���x���2ɴr�H���+e5�n�z��M*Q�J�6� ���B� �%��Y��,���wF	n#f=�ţo�������X���Xv<�e�3+(Bĕd�׶�P`ɈViʽڭ�N�l�hJv�l�T�����#q��n�E�X�{�V�|�iմ�ee �hN�d��r�Õ�$!�R�R��&nDԎS"�o�$*I�@VnѥD\�����B�Q��� ��M��E���O��m���u��C��^�Bږ�ˏe6�LF��2��f<�V4�������h漹[�W6�����u����f�íhk����0�8�%(�!h%W���B��7OR+C;uQ@ӑ�p�l�g��У����wwN�z�Z00U�/�ZfJ���9{{{���q�weQu�B+Y��pnd�I!��,�A�i�/6�V�k��y�]�S �Zȷ58�%GjJ���ke�aLX�+o6��;T�ѹ�$��M�R��W42�.��ŬMȾU���'�G[y1a�ȝ��(�u	��u*�A����IN��t[���m̫�4@�ۧ�N�!Eml�zN�gL��5tj�5�Q�؛�Ӊ�5�"�9Knf�ini׊Mҭ�)+�V��e�x�F��jH��q��NK��`�icx���-��+"��8�Ǆe����4�M3��7���zػB�[@�gD�VM��v%�Pa��}t�Z���H���6��4�Y�Ra��[Lz��k/K�su"���ܬ�����b���� B��С��	�����\�pL7�w�Z��K�V
)�fث@�;S�/B�3+Qס�V*0�
i*��o%����Q�Ԟ��U��
��V� e`��"�hW�-��>�I^�.bO)+�B66��0&�\4a��0��72�ڼ�tH z%$�u�@6��#LH���eM+Z��)�İ�Y�)�(f*��Q���^V'0�&��6�E�9Fф[���M����ʉf��`ա�B����Ñ�%��#\8J9��C)��iJ�\�Z2H��2��#KWEF��Ê��1�'"�V�j�ad�c*]�Qn���x7eA&؛����������d�a�,Sp���^]���DfX7a���Sj�ӗH+v�i;f�a���������R\���H[7�h8n`q%�k0�K	�*  61�ǭ�%!L#{��������&�L	M�r�l���+�㧺Au�"H�Th�Ƨ�A[b4�a�Bx.-��E] ]	h
e)>{�)F`7�v��嬫.k�%͛�S��E�f�T�eT.��i��k@�����o�G-[i�⢲df�!����eL��`Ԧk������R��l�'Kn�@m;��S��kł72
/K�����%+{aK�y[���x-`����E�����Fķ�ʤȻ�,!��P�J[tm�©��`�-%�-��������C�P�Pn�v�/�b�� �)���yF�
����Yh��t�˔Ww��U���쳤�ژj;����֩Vr�E4l%��o`R!��Ȯݓ&�ړ(e�t-)Q.<�:Qe��xf�EF�1�N���%
5xnVֶs"A�"��`n�����ֱh'[��V2�=��3	�SL��ih�th嚉i˕(�qhE�+�74el�&���(�{K3��X�߱<	ih-[{�����f�ͬ���R�P+�w#R,�%��5%��[���R0��bN���m�o>qnBh|TRsN�f�^`��Bn�ig1eLJ�j0
��e=�$ٺ�'57A8�1Z�'���`a+��Wb�I��X��	pk96v8�������tnat�
�Ϫ=��)5��
�	�)f"w#�l�&B��L	á���2��J�7]B�+p�[��۲kbz�7%�*���tE,�eFH�P�9kSK.HL��?��[�n��d�u����2���[��Xk4<�nc�1��ʷ{)�*fWZ�c��Yj�d��-�h��e�$�۽ H����.�+U��@�(f���*���.�ll�tĭ�w�Q�@�^���Ẻn���'.�Z֑����Rl:��;f�V�	aѻ�
`/�&��0�i��e�[��7k1��j���4#��n��KI$��JV�X��9v*3B�Ō嚗"��7��|�w��h�T�)q:5{.��ȉ*7&,��3]#N,�i��M�okM����ՠIu��ؘs���51JԒU�X����<ɭջv��-�J3�Yy���H$�{����H��V)ۙJ��-9�I�A��-�wr�l��+X��!y�.<�sE��)��JUռ�hZ� �ѭ���V��Q�2��7m�Ud���id�D��(����[�^n�9,w�Z��'"��ܽ��T�M�i<�ِ�m��5e��0%�m�6,&�cg&����;���u �����Y4 �/^���E<KeJH�f�F�*�oe�q��;�[�B0P)��W�=�������=���K6�9)]҇.�dMG��f|��_�z��2�^����g-�CXæ$�eX��uh�w��hAu�� �)�dEn'�$�|$b�*9��	I�SN�M@i��ӊ^�4hն�cm�$��ø�h �%�W�Z�B�2s0*"�.�������+o",�x�6��hZ��Z��d��q\nH�D,��i���4H�w�5G��5��0�Ь�`�Adz��m�5� �Kwf#V��4��� kЫ3#٥m�1���0Zj�M�iIQ�gH�Nʚ���/S�N���S��ӫ��[)��.��ɂ(2�B+(�Kv\7�l7hֺV��gu댫sҍ��`�W��T͡�����`iyh�n��u�;�{����p���k/�ڕ;^͘��.Xp�*+nR�ct���w����c�ƨU'��cn�m��#5��tH!;ChJ8d�]�՛�%�R)s�:�::O�DM������O���~����8v�Ο��~������1?W���?<8�������
I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I/夒I&�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I,�&C��Q���;9s���O��5h�3�.`|!��v��&���_S��	evn"A6����Bs(��}a]��n��I��ʜ�|��݇gJ
��.0�Aۮ��H,�v="����@���q]	eN��f)��d.����yu��1a陨�)�uzv�g�Y�"(q2�%s��:E�����V�b�w*-Nu��*qwݠԒ�S�yҳ��L���g}�cK�Q��Dl^V��Sx��lW�#�iխ߮�ؙK}59�j$���p'�if�1u�g
�:�b�M��a,���h5ۅb�j�����Q�Y1�����t�"ʶ�C픒﭂��1�����Y�d}�zVj�ž�[q�b�,:v��?TJ��k��CQ�q,��]���;QGI���|Ɠ̚W�
Z�[�꼥f�BH�X�N��s*�oI�q����м��@s��ub
7�#Q�B%؅b�EE�U-�A�dh;)wlk��;z��M*[�ggq�����_KR�]i�fR��\�0�7�c�H��vn��S��.��n�o.��M�noX�IX��;��]�]W'B�Ǉgfۤ�v�i��Lȸ�:0^;����J�*�`i���0�̞z̸0��$X����t=Wp\�qq���+b���it������\V*
�m۝��V;>;��.�j��i��ov\O:Gv��jR4���Ք?2g���ޢ�np�J����:�bS	� �,��;�P���;�a���[���/{�4eLY���5t�#�a,8��D]a2(vmD���|5NX�Y6�4��|2������cT]p(8͒{��g�@<t������M��K$�ۈ��ks�K5��])̫|C�.`Ž��U�9��*o����mffJK�<��Fj%�j���T�ݓ�Or�Ca2�s��k.��nԳ��wK,�3-�O6�qosh���c���/��k[���E�alT�Ł���t�p�����.}�.�x-*��[ڻ���\Ӎ]\������cfF��Q���nJ�ͼ��ћv/b�\M]p�}���^�wm�<��zG����j���@���A���SU��r���jZ���%S�d|��Y���_�pu%���� n�=[��%��/��ǥ�ʸ��
���c�}!�:��{]EI"�٭G�t�z�R���=/P��Vm�F��E��9g+,��� ��K7��&��٭�w�-x����A&�""8������mn�� ��錩�81������;�P�;@0Ǜ�,)M����Ar����`��
�N�
:�ղ�)�+:��Ƒ��1�`W1*�a��؛v�b�D�+�$j��O:������j�;;���:����%��ʕ��u�[U돝��qg<�`�z8[ح��nv9Y Gf�M8��mt2�K�й��9-�9^Tն�P���x&^u��ﯜ�G4u\s��i�5˦-ݾ��mm;'���Xu:�Q�5�I0�bҧU���X��*F-�!��D������q�{%���:�9��K�vp*���vT ��szm�u��ͭ�gX/]� ����u|��Wʋ�Z8�*��ڷ95ӨO`��E5���5�oX��P/�Y�U�;��OAx�ν��E�V�� �]�%䁮���s뗴Ȳ�+�'|��e�lݩ��1Puv��/;x�c�;K�:��r��G������1	+�v}o9W]�W�C�A�ɎWgV�z.�8�[HH:��[E�c*}�d��ovHl�[���u1�2��{Mx�H�w}�/�^}� ��a_lXY+�^���9	��,qH���^�ml�Yx��+A̝�o[�t��V.ڜ�}t�)��_l��F�Z��6�k��V.c��O��
�.77鮁����q��_O ��=�u��\���ɱ�v���̱K�Aol�9S�2{��+2��]��Ϯ�$c�t�P�el�er`U�o�f;��%\�Hx�דy<9��+�)�S�,P�yt���#���MWP=��c+h`]S�*[�(��颪'.�7X��\uG˷2l��3�ul]�Y�!=ڂ�Ǘiiv�j;��n����[CH�r�M��6��-sT��#�:�eGv�r�����:��3��R�,q)s%�R����2o���<�����#;�e��Q���P�Hk�g!fpi��f���3i݇S��.=�E�\]�A$��و	��G;%���Sm]]
��xe��To��sg�\yr�T]uc�F�je��[� 1EeI��!�O����R��'+�,;��_���gN�g[�a6o�k�"	��$Wk��IwVlg8p��J� ,�*N�n��/j-����ﰩ�jOw&j;�0�,�y�:v����#Y��Rs�,U�!��-�H��6�R��t.J���0yHT��b�x]2��j�྽YO�$��5�*[e�.*�F��%r�y�
B`��[/�u�+�჊>��1z7η�qT,�.�۶�;T&f�Ϯ�^3SxP=͆rur���dR!��r��<8���n���0{�P�����rf&z�I��˫�nu��C��K�X:��V��\[N����mݮD-�P0{_T��M�������y�;ʹ��kH�p��W9��qo�7��	|�6���\�)]�9>|2�E��	�uYAXy�6�h<�n�d�]�)ut�so�鱵���ږ�6�e7i�{ԢA�y�.�M#��p���(�hM{B��ɤb�-�؇ݻM����s@��S�h��qwW/�)F����F�8d��o��$tb˩,�wΚٵ�.�m�e����-�r�QN #c]i s��Й1�ʣԐ���؍�e7�J��=�#[�wy��תE8<����ô�lk�SK���ygr�����@Oq���y�c�AT�)h��r.T7���ɅS,s���	�zHR9x��9���Z���))>��z2N��
��*:���ʽyi�&E)v��͌A�����Y-�+Mj�s�:u6+-�h�j���=��u�F �l� �C�}+8��u�Z$�\�ywTV�hާ+�P��{0SF�<�����������աE�q"��^ÀjW�;�ٮ�B�4�ϋ�3��6j�O�n�]���E
��]�w7H����.Y �����gK��:��z���wxx�\Kx�;9�D�Zt�; �iZ��@��tlz�u�����C��u�B��c{\��vw3��z���G6�u`��YQfVp.��d�v�b�o,�����r,͛W��{���� p(�Z���I+�
'iU��bԞr�"|L�bqF�w'V���ӑI'I�mWm}:��ɘ{wge�ptcj�#<��A�����n�n�����\�uJ�N�#k$r����.g��
a6q��GC@e�p���*WY^U����	v�rf��賅:wwv4�2���gĎbI����j�.,ã�ܹ��Z=�i��vF��K��}$sw릋=��$��VG�ϡ:�x�nu�U�9�|�a���t=x�u���;��GM7��T��R�;Ndp��vv�<+	�p�M��)�j�1l�%=��U��=��G��a��&���deJ��]k]�L�]rƤ��.�V"�^�],Uթ��=f����&�D�pBG]]�S��N͕0@.����H���wT���V!�/����MV9d4��ضӅ�h�����ս5����ٹR���r��EI�,��-�be�c��ic��/{���������^��kgv�Y\n�+;���		J틍�F�>ц�e��`ڇ{�ȹШ8����g�k��kQM�TB�ӗb�Cy�/p�����&��3FvƐ0�\^��kazͨ-�r���v���N']y��:��J!	J�f]o*��v�A�K��#�0��'��ՔhP��`Of'[%,��R��0�2�f `��]�˹P�7��2�=|/w��w\�@��Q{���;XQ�ZF�c;eY��#�ld�zmD��Jc=hz.s����}ݝP<�SKO v u]k�rWm�q���yp�<�f1��z�Z��Lߍn�5�I1�,�Ե�RJY%`��ج�U<)\֚����
�{foPt����Z=�G@������xhՓ9+M:=�
zM����=�k 꾁'֣n$��-J�kM���ir���]DU��V��oT�5ku=ʒ��8��sTK���:3����¥=
�5�Ch���WZ�d���+7��hP7�Wq�4��w��d�`F=�C��5+�6h[NJ� Ҳ�\&�u8u��Z��]���ߍ�>n�*av-��p#FG.�CX�;;������R�T��3�)�r{��m����^�]�uv�"����ll�e�|*�6ԓ���cl����hM�=�)!*��H�]����/kSE�M�q՜ӣRnp
vU��	��c;`�U8�qc�!y�y��v�VŴ��]���:�A����A*ע�,��Y���т�k�9Ƚ��v�K�+s�僺+�;�J�[�7NtJn�zb��A��5�^�u�ʶ�Ad�=`3:�^��/c��_�MJ�z��yu�tl�}q��S+$�,�!���%�t���	����mEQBE�,���V��HH�1��j.�Y���v���#������m����ŏY��p]��cK�3�}��ܣ׵c�iT����M��.���ʝ%�Ұ붺��/��� ��A��ГB|�M��q�����`�w+1E��X�E�����F�W�����T�k��J��0��4�;fG|��pj�wiF�r��x �,8X}�YW�P��yY�ǝ���S�d�9s@L�2=�6%���͘G})X�dtԻu+\��{�E�����7q����Z��t��:��x�q�Yu��-v�3B
��L�������J"=����4T�N��f��4m��X�A�{��j7ڸ�&�Fg#]��F�,.�G�G}C7WR�$b��2w):�=�YӚx���h�Zc�BZ�Ojv����#�b�N���'R�C���n�:�g=o{O[�]��[���y�����m�w)�ؒ]o^�<�>0�⑬����[��(�q�ͫ�0k��vD�qۚ:���h��FL���T�ܦ�H괉]1��J�=(��C�JD���QJ�QI$RK��"9ZJ�()e�w�v�d5�hx�����,�vNM�7r������,ZQJ����I$�I$�y$�[��I$�I$�I$�I$�I$�I$���W���>(��~}�_���z#�Pm#�u�"��׺�'�쌜?�P�?�>���<����3�Zb����cU�h�b��ז�阉cvZ����d5���˻�1�.YRl�\��݅��oz���p��+e��o>���I�ۭ�%��eN0�5�!P-�̳�ԾI���ovm
��&A8A�Ct04�|a˦ ����n��oZ��A�B��SY�k0�&��7b��c�kM���
6�Q`4n��}m96�8ę�hVq���Ss�f�0�ػ��]�\��Ns�;��y�z�U�99�Y %��n���<-A�f�0oh��Ee?�Rn�R�m�ө�j�Xr�T�/�{��-�Z�	��%_��Y�(u�y�5Ç\.��Wz���r�PŮY�0��6����  ��}K�I�Vn�M�JA���ړ��u!/v�^T�{�����?U�p��9��HV5�yY �>s�=ƥn�KCmZ2�˥bnv��Z�m��0�ϛlݝl�=�o0�0;�	t1�K�$:'��CI�r]ي�cj:[r�M�t�r�����y=Y��mc܁B/�`���{mr�掱žy\Y�[�Ģ����)E<YX���݊�RgvQx��M�w���Ul�e�ų[$���ya2`�^D���yn:玭n|Β�vtö����qiȇ	��f�����-rҷ��-�����^l�i�7Vh.f�ة�AQ%b��Xmv���e_F8��Y�P�K:1Q��{v���&�m�M�K0��IK+V�V���V���*=��g%@��yү�n>�֑��a��.�S:�1"��{9�U�Њ9[�"�*u�|�,/�T}w[�t�������4 ��*�,�$RUf�� A���)a$ -�����6���Xd�`!ڝ�u���vjcU)�fm��1U�'�,Cb�z�����3{B�V*}�-`1ni�Y�;M�$mZw����R�gD:���v�j2r69�#�@�����;ĩn=V�5g1)�I���<���N�fvT�5-ub]��ܻ.�|0>��jy:�r�v�o�5X�?�0�f�e�e�/R��?��k��U7�t{�D۷�Zcu]{��V���	��4�YQXrcB��Z��ҭ�"�Non��H�V�Ә�?�U���s���Vz�:T֤�A�WNM�h�?vȭ�	�A7-��T��X�Ef���wA�q�b����lGU��(˂��kH�̵2=@�+$���:�&�6���<�R.�t�k������Շrѭ�ҩ�S���X��WxC�v"r#AB1S�0xHM)��ӟ7"�.�pIہ�$�Smئv�w]�Gu]e�v���N�R���U��E	�A�(��A1$���RJ��|ܗ�n��uq��G�;N(�Ӝ;Ydu�0#,0﨧}���Xqn�SbY��zp�ݵ\�ݩ��]E���͊�D���Ôn�]�v�W1-�K��K�Ĵ��/_k����3Y���Z�A��*
��k�a�vnL�Z��Կ�����4m>6
�u"wo�Q��#s���*kҔnQ&��6����W����K �e��,M�d��)�be%uٶn����]S�q/`��_�Qq4�n��9�f��u%����g띯^]��d����4�]X��1/p���A��[����]�ɗA�u��, �@	��w�V`��We���\T'P(�DWmv1�I�09j��V��m�`��f�i[˓����JѮ� ��%*7kn���l�z]���z�h�J�V�.|�G���[j�EAwyN<"�C��w)
��H:+R�6𛿶�s=��^��=�}E1ͥ�2�P������qhޖ�#�U�"����묅�|i'�z�S�.����>g:#Ӻ��
� ]�%�^+�֗SSh�P�c� 'U�z#�.�J&-�{�ΥO0X�N�J�'U��v�.�
 �\�f�%�U ��U�r\F���p�M<[8��4�^#t��7�����,��ofE6$�K(ɛet��l�Y�1["�[�\�:�ݦ�/�zb�kZ���YM�6�r��g�7�	'ys,�/K��4vn�iǺ2��R��0����"��>O�`�YSr�;LU ���c����c��Wт��6�0cf���I�N��\�tk��wŴ�5�K��N��[0�p])}:���K"�&v��h����		6��i�#HU�[G9Ky�����+�+R,��9�2��b��Y!�Գ��ȋ�bLuqfÐd�`t�9��g:(�a�{���]J�.uסe�{� t[K\yL�-�͠v�pW3t�m�����`H�f��=��t:!����s�|�#�s�����tIĈ`u�h��`r�	�Mq�o�a���/�f�L����{����O��
���R�bvԼ�ٳNP��������3 'o-�9[�uY�#ƅ@Co6E�N�K-/�K�Q�Ѝ���w��GC�����<��%����#�Y"Ce�4�v$��=�[`c&�d)����cQ��]Gs3H�Dv�uܹr��ڒ����ܩՓd����J�*���e����\�����vwv-��v������t��F/�d��^K�m�g�)[�A��R�Əj��'kR�2�e�<镗KD�U��-̌�)a42[�PH���o�S�]�23��zٴ��I���q��Ϙ�L�9A��\\o�:VṚ�5�q<�:��dy���Mۤ6�r�)��j����)"�2r���\��ɣ7.͇Hd}�H�Z�=�v�ج:#t-Î�km,}�t�Y\��w4ݘ��nmC��F�WR��h��p��-�x�`�@!��{Z�;�*[9�XS2�2Ը!���E�z-�������8a�6��!�LYc�}�e)t,��k�e`�52����bt�ʇ��#Bn��/�:�-�ދ��Qj��.���Nm7ۚ��潾z 5 ���˃
!t�Ɍ�Bu����/oѴx��zε�3X2��:z��{����ȫ>�}gb�R'�W+kb�f�Vg|x�'��Ck¢��4��,]�A��b�t�ܡW���õt�6ᶋ)CK:]���k��nV�=]��3�#�sRVV:��F�}�S%q�\]h�m�Pʷ6��A��\4�cFl��[��I��h����}��I7p�㯧V�۰�t[���\]�(f�6�+���8��[�%iy��Vz�+���܏'^�Qd�j�ʯ.�� t�튑P���J�aF�nck���ނ2Ѯ�P��=ɳ�y�q	bcۜ,q��Q8c��Af$�Qm���3�2l{�u�V�_R+��%IN�<'����w[vT�$������R����"�7�*Щ&����]]3��[A9.�\���byFVV�-�eu����Zt�o_q�|��7����Eu]=����̥Ӂ˶ی�Ulm[��[��̧�T�U�f���ST2�P�L��+��"�oR��A����s.�OO��t�VJyۄ���1ЌH�h��Onhf�.kQ�Y�n���]Z�,���0��Xy*��+�(�2\�0忲���Λ�� =Z��J8�j\��nœ����*3�`&�n���҇Li�݂oa��T*�[�\���;5��� \Ǵ���������@���p�Z����R^��5|�YY�&�r�7 ���fS��m>�9{�[�S.olVs��iY�8	�C���V�u�5�Б@��V����Q�U�o�k]Ƭ�8z�d��M��wY�᭱�(T�1������V�����m��i�a�ޫ޳������%L���#��l^M��L!��ˣf�
{
dv-MU��N�S�@����&�FQ��qn�T��ސ�sGoZWZ4��];3F�ѐ����֭F�j��*j���)ɔ�ל��ZF�V��	F�'�R�*�}�c���+�'��%$��Q�!�V5���6CTt�G2��71`������;<�:�
N^$昁�7-��,&�5u���E��]G����̀�C��+�W�	��<�emplP�GX	ކGnt�]�34�,5,����4ܧN��������.R��J!4
̗f[yF_E�̳wu�3[�m; m� �X����T�2��_)�K�h]e��T
�����z�fQ@Y��arYK�F��{�q5�ί�;����q��f����7k7*��Pr��
� a�����ĵ��@��������F]�f�*2^�����[�un�M��H��$��c&�:T�m��K�Sdm*w��X`� �a�Q��J��=��u�6�;¥�M)����&�=2X�S�m7��#�Յ�갥:�+�P1�H]��VҾұ�}��o%��=gAdAʤ���1�!en'�[#�}"���Ƣ���r���X��9լ���ЈF@�Mu�T��s�v�J�
�b��)t�=�w۴ RG9�m(A m�G&�e�w>�����i���ܝf����X4.Uk�j������orO��t�L�[b>|/93.e�M���,��q+s��~Ρ0Kzh���=;Oc�1��HEh��Ve[UD"�l�&�U�H��bݝ��[IT��1��}a�ɣ�^���{3�\���l�V:��$$&���Z�d�P]>�,�1�LK��rŘD�	��U�]�B���y�̩�JoȒ�O���a
��8E�������ؐ�m�1��酾��濈q���U�f���5���؇'��^�[�ˬ�:,ٺt%0K8�)��"\�ם�9a�nn|�P¦fUQ����R�J�T'뻹���_N��[�h�t{��y�Ծ˽�+ha�].Ww#Fԗ1�+�p����n &������k���,-��Sػ�|x�ԲY���)���Ӣ��)b��v��"2_�
Ir�z>6���ENo��7�dPv&뻴�j�yWE����k�o
&��$���{�I6BjKd����B�N��S������iPz�9n��c�u���kѧӣ�2їj�RSo9��l�WcM�7����g�[oeb��{`r����5���X��G����F��ٖ���Y"8��28t��Δ���;�X�&�ډ#����7�8��ǅ��g0P|Ē�$�D������g+m����8�!5�N��M����fC\�����ʬx�mm5P�o�����]^H�r���u"*u���Ĕnʌ�����pi26�znu.�^���^��i�Zf�gz�6���fN�s0J���wT�b�o���ȹ�}�s���)�b����?C�Q��hp��c���=�}�$�I$�I$�I$�I$�I$�I$�I$�����
�u%���;n�S,��������xgU�������q��v�ˏu��J�$ULb�צ�- ��T	�֪�U�H�DO��1��&J��v��T�K��S�
�:�'"(֚�f1�z�
V�;���9k[2���F��> vS����V���^���h��v�����.6}·a�+)�W*�.u���)�.)#K6�A����١�`���̏��z����ղ�$@U��K�+)2���3��nّ������,�zEsv�䦝�G�p�\a(��5��EswpK-�Ղ���9��[M�����ZG%=��+XSx��K[ƚn���K�"v3D��T�
�t��Q7�ۣʱk�����Ҏm����Qh�Yˣ͵�c7���՛B/	�P�t4��{�o1���g�Tő�F��a��[����t ܊V����M�1�Β�ɪۼ�]�L���̨��:�@+܅�,�Ƕ(�lp��v廰q�����H;�n\^%�����AD�R:�H��+��'д�%PR���MW��JQ'1��4�!ERU!MJUA�d�-!P�P��d faE15I@D1�IE4P�Q}c@QM$>ɇ8��sb�fMT:�
�,�D�����	�����*��((�0u(d%RDR��L]�a�\���h�8�R�k5V�(��*���&���b�����fPd��X�5JUP�q��55KE,@�P��U-UHSE-�ɠ���$2K�W������bD�=Ƶ�d�d�D+AT!AAI�2�(�2����5&B�)�%4��$Gr�P-J���@`CIY�AJ|�?�]��pwM���u�K{��}�O��� '5�M�z������e�|�=��4�n���K�$گ���1�P���W���<��=������ep�H�k�ܮ�b�E��"G��!��mݗ:�4
��N�>E���lY;������hn'��^Q*����\�P��vJ�qK�j�nB#lv����x���+�����G�kiku�cF8�������;�[������ f����>�h3{�F��1i��輜|i��L��}PW9,�Ǌ��Wp�;̑>�"�^62�}�Fţ���ڞNgEVSl�go���b��!U�������LZ��d,��������A�;TT�������9��S�Y��O��ݽ~�'���vΫIO���,�`?N���Uƍ�{i���� .��ţA�8�%W��5c�ρM���.�R��n=q�_��g�e��V]Xf��M���M��=�<�[�PkD5Ϻ�+�b��
�f��%S��T�angRiz�5�^�lx�����S_#g$!����u�&/��%b��*uijqOw����P��W&0�c�㧭�<�gq�H,����b�+5U@%�4�1��Z�����=��b��rK{��z��t�Db2��K6��aZy:��ס�j������Ҍ^򸧼QoF�[s�w��7g*�8� �ۓ�ooձGT{��d����ۮ���-�Џh��;�_2�v��+�u�V��	���t�*�Ss]M���]m�y͜��/�J�c��ax�_@Jlml�s������6���\;�q�ގ�z�mC��=�.��!)U\~͆���ס���rC0obWm��U}�}�âҞʙ�\'e�� 5�
��O.��Ǟ0p#{#=uϔOmT����ĤPF�pQy&�����Q��i� �W���W;�ވ��c���;2*�����������CFtk�,uA��k{��^�.�t�g9X��lr}[�k�\Y��鯭4+/�����5�������X�jE�c���y�^N^6g.��藺�4n18q�S���&�vۋ��+i�{�I�����������K���4�e��E�uw����`���Ԑu7�\Z�K3+'�S���WL�.��S� ]Zȷ2��;���I��S�l�E-ۅ5u@�g+�6+fu���;�X���+�O:=8�=�K�.�Ϡ.c�D�	ᴜ���e
���+%����k�ӌ���߇�,ԯV�^����ګT�]D�!p�)�{R��^�C��ו��m��me]�Du@:�s�<]��3S��R��Ҳ��{�G��n!����s����9V?,�%��&z�l��v����ۉzx-ù�8�=����2�eq���%9ʸ�OȾ뎁�.ӕೝ�i���n`�'n^iE�����JWBi��ֶ
�ڹwfV[�!v�)"�]ΝFr�'Foqv��k�__���7�S���� �w��-a��6q�r��;���+�)MAW#P�esk�������*�;n�;�t��3&��D��Wi����C�<`�ct�����ڞN2���J&�L%p����7��l�򻳛�V�1�[�M����}�O�(�i�v&̻ۅӷ��y�,Ѹ:ZΥ]�/�ͼV�o�nw�@�u�0��K1x�W	�9�+z�5{�Q��Z�����0��=hɌ��P��;��ZoZ��oOdvt��>a��-��Wٸ��|^�"�0����V\s[q�����mn��͌�3w;e$�wYOA�0�����˄���쥭��[DL�j�������ګ��v,3w�4z��A����.l�D�EV��&���P��,8�':��3��µ��L�y`�����!O��j:��:�*�9u׶�#�S�P�ݥG��;\��j؞�!rY�-�������E�_"�-:�{=bV#n�o���N%gB�2�)ѿJ"����jަ����ܽ�g0����
���.͆:�-w�̝��r�"�y�r�wS�m6��1�uOa%��^��C���ued����tu*��I("�xs�)��ܪ�eH�9體�1=���Cr{��1�􎷻�o;"WCy�S�\�el��Y!�z[�BuL��0���Oc^Д�.�};yKj�Wݨ�r�Û!T�-����^��y}|�5gz��VGx�w�fu�߆ʔ�P��=۩|�J6�]��{)��F+��]Ɨn�k�wc[A��ˢ�q������giz��` ���������+��\�)2�C"X���U#�����\�7úX����Q
Z��N��bA�r�����¯h;{��p0��_v$NEԩ:��(^�۩��ܤ�댽���[9�{w8{�̩��G���/�>Ϋ81��	�<��c�"���Oc�m��n�ט�>�+�k�O���oe�)�2��;�wi��F��}R��Q�z��rxo7MN[ޠN]�ԭ��[Xf�t�湨���<h�s{�'I8���r9��mmĲA��m���[Ln���&�n�N�W��v��ᓷ�Ӎ���_���9 �t�z��:qenm��gp�X���R�w���\r���a���M#s�I��N�+�'S�H����rʓ�tfZF��*D��<5J��1�Y�r�B=ڝA�W[�n7��«'���8g{��>��'�{���{q<���wRn9\�f��˩V��F�w�5��Zr�v�M���=)롤��mT<�5��l��RR@�=��Wps;��v�*<[GLpu�!���z�hڝ ���4��t�]�m��k��!�wr��מ>��
��I�k��b�@6<��l�jz!�8,iҠ�K�;����f����>6D�+��V���x�e�S䥻���O�hOV�j.�����ʕ�S(�q�mvx�km_9�:� &��T�嗓o��/ܺ;w+{N��r��/��K,ӝ�*C���~U��o4�U"��Wk��+���0<{^Z깈�+�X�m��l��E�]�d�Sz�k/'�Eྼ���L�3����}.3�$�\�v����m���tm��/SyG��&T"۴̖J˂�}�m�ȇٜ�cp��tV�eV(n����6�z���$/K���������,V�2�^T�o�gk`7~���
H�f�H�^�u��^.뺊i��F��8�����/�V�k��20�{3�3��]�K��;�vvt�AL`i�#��}�WW�k��̎���m���g�m�Fy,$��o%�NVOBv���bT^�+��.N2i<h��}���S�F�ň��/X%�\IᅼĔ_*�{��qudFu
�MZ\z��^�Ak���Qf�>�<�Q{ɨ�ko/n�0��ۄ�� �m�s��d-��դ��^A��HM�w��}['5˟4�w�Y1E�+��»�m�wq96��&�@���P��J��J⸥5\��!¢W:�u�d��]�����,bg$J�5I)�Z�Ǯr&f�/z����=��x��	�:a.�CZ͎C���-+6K�;8�W�]E߹�u}G4>귇#�!�t���,F��M�Ӿ����l�xb��Q�+�X���0{�0���7>�t��;l�qp���Os�F�vE��:u�J_E�r���X��*����;��c<��vf�ó�8G���CK��J��Kc'LJM�C�R�
���vcBH�嫑��.6��|�lb{���ה{4U�{%�x��n$������X�(�i�sC�7����z{#���Z)n��˺�t��;z��������y�Yq�n"��}�f+��ۤ��)!��[l�N 8��>�j.#8�~��\����m�"WuZ�vK4�n�,�0��I��E��K(��h��]���+dQ�\\D�qÞpE]:!��^��1�n$��i��JW���j�a���g�Y�r�	�jQY{��B��ʳN�,��ud:�y}�Hl��F{��guF$�Z琕�Juz�y�W�N%�0Lp�Q��oufl���㉎ul:�������V������Z��¹KT&k��D�4��.�u�*e�6��sMB��ܳ�+���X��"�{"Z���l��;i>�RŴ��';��t{��j]�ʻFgs&�ȷwk}O-8�	��w;�83zw��{�x�=�c�ݍN�^ЕJ%w(rOE�X�R�Zƛq���e��S�Xou�	Ř���륡cѥJ5C���Cym���׻E�n]��Ryf�x:s�_`��q��m�hkwT^N>��KZ�qR�?G~y'��+�A�t�q�(Qx�/zgU��f̜�F��x�ujQl�J����bn�!J�ҷ������ɘU�pzI�k$�0�j�/���.o9��Sؗ�e�x��)���)�m�_gM^m���sQi�ˌ��h�=#"^Fa+PW���)��9��um���/�����}7�P��Ņ'hM��̠\v�Eb��6��~/T�%�&�?�D1=�����~\���Y��3%�OM#!uɺ�6�;�ǮMILO�sj�f5���gaҩ*
��l�=�����)wPհ�^_q�@��t ee%���@E�Ԋ�h:����T��������(�������:���n
u��09�V86�kX��J��4��+��c;����Н�;�K����P�����$[*c]e����cJ��,�xŪq��C���oGǷ.��!����)�sML�S����.f+әؙ@'ս�`��x:���u��KM����s:�G.99���s�ap-�)ӝF�Q�6ʼB��M�K����#܌��L\�O{b�C���v�97y�xr*�K�V�.�1�3*���]�.�����j\�R��Z���4\��Xf��=�$8j�����I�Wږ�8���:%�,�PA+(�r'�V>���-7��ŋ�K����h,�<P7������[i=�=Y�gXl[$��*�'�c�"��uˢ��[�Xœ+�A���˰�dj��)9�̮��&ޞ��|�/�q�#�T��e��Pn5Wm�e�G�ΰ�{Cu����U�(���	t��m����8s9�Aʃ�k��i�!�ދ�o.��b�_�>����'���$�I$�I$�I$�I$�I$�I$�I$��͍��)m��[Z�*�k�m�9�ei�p��gNp���A2���u���7�{��U�u�Sub|j)��(�帴Ӻ���!����rs�*��Iu^���oR&���l:�:*����0�W۴p��tW/Mn��-��[Q�f�hyH�F�k�=�l:���?p�V���N�w�
i�y��o���l�w;���5�4hj��
�nʽ:�UV�؅	��� &j&��r�����.
��-깧v1�k,7ӛ�ϋ�U�4�\ߋ�Y�}Gj�'�ۼ<c�b�4]h��T *�6ow�1�\i݅��ͧ�oyɃ���,YՒ?��l�σĶtV�4ig�ܼ�a-�x�-Im{�0L�xz��t��D��w\	$�\Y	T��_a瓦�,��в��e�/�hT'Pǥ��'r�7��U��-�� ��fs�'����]�9k!Yr�]�;�5v��`܇�r���iX���_WU�c,�'KM0�m��o-Ϸ�Үcd���쥻JA�Է"�Q%$���$��{�3��������((��%(���"*$J��V���"JB����<�Զ�)Z�%�ZF���h���Z@�(��(j�eLYK�� d4-SEQ��%�dd%&M"Rљ�R�.@Dд�4�IJ44�d�4�L-"۰�r���JI����&����D���bF�:��*��-#HP�%-%!u�d�!�E	BPCP���i
)
�)B�@3#�2b!G���|�:prԃ�eAY�u9P�p���w�����������*��f���-�f�k�e�9ې�(
���D�Z?"
Os�U[�;�Cב�
t�F�x�,�m�ټ�t�)n��U���g�Q�^�����w�nv������zy��؄[%�~������'��j�X�[9J{��sK�p�'�pؗ��a���ny��\�^�w�p5�[�����ܛ���4P .5+y���������B�Ӓ�=����7�Z��jrG!�:�]^��=����=�|_:a��ÙUF�J�n�r���]�dpR� }Ǖ����7k�����T.���/g��}��G4'�G���B�������`�"u&6\�`�*>:-ߺU���K}MIز�E�x.Ŕ�d�I�Y�W���70����~�a��z�֜���wJ����k�vaʹ��˩���k/R��s�њ߳���ݜi���b�Y��RI^jB���7\��L띁m����yڻ��i��'u��s���e���?o#�]���ؿ�L�Q�z�^��.p`�Woo��Z�]K�{��sk��[�dD�8۬��U��!}%����}U�,��}���e-�58�s��}Ἱ��F��F�����i���q=�|��l�R�p�&:21��|Jϓ�k���U|+��/Q\J���%��Q�Btk��*��qc>���}��p<60���J����b��ueiة;��so��>���mg��:�o�1ʬ��`��N��Ujjqow_D�߽]�x��~,}Kny����`�!m���Ge���,���J������iZ��'W1�*W�˫�[f��sR_�舛	�џ��⒫��Y"��b��͋p"�oU�SVd���;"�S77�H�"�0߭�7�]q�*���+�Xýx�����v���~=(�p�02�8�J��q�M��z�>mJ��O�Dƻ�E��P}۹�;9��/�S�����6���xv�+�Fi�Cj1Z�K�J�Wh㢷{�f(P�z{�c��2��:e�츫�@o죦���ue�e��CF6���^F��{)ΪX+���I�Cڐ�"�\jE�%<�9���T>ɨ/'Ρ�V����=�k����~��W�m�L8/�����ہ��������j�fv�h�[�㖶��rB��z�o7���]�m[��y���T��m'��iUV\s[x�}�o���꩓)"Hם�JY�3Kf6浨����uR�O/U�g]ӶaNN�}e�X�=��B��T��D�b�����#��*c�G��=��?b��Z�����P鏡�=H����C���K�ӛ�@�����M�ԅ}+�Ƥ�jW�a�O��rC�M������R]�e~~=^΀���}M,9غf���+��r�KlH��o.���������"������Y��KR`=�[�W�s��Z���!z��m��,�`֑
\H�>k�6��˕x���N�r#��#���y-�p�z��"#DA�G���7��<��Wr�������>�Q�2S�;��;�qα_&��"���>,��V���?}����C�إR�/�0o��q�Wr>��n���:�zG��^{ކ�>�ZSP<����{���0!�]��6̜s{�������F|� ���"���_��(>��y��$>��>���	Ʊ|���q��<C�J�D8goޡG�������~EqW���!���_c	��vs��%~�q<��N;�����k�G����1|�!x5����~���j�� w�6���4{�"#�_�B$G�=ϡ�}���X�r�j�G�㎰>�G�89��9w)�x�+�8{�7�F@��u�������������ͥr�N���K˯y�rs���u��9/����.�/x�O#\�qu#�A�rܧ7ҹ'z�9ݼ�vl�o������J�5)ԇ]�(7.৓�&Cܼ�\��N��\.��{����C!�_!��;�b<��>y18G�*�%�����T�~���hd})���W' ��}���=�pR'�ПC��9��!�^�dx��w���]��f'��{�e�7�yu&t�����-l}��S}����|��5���A���r;�e�2�w��w� �xܾ�<���z��ԏ��={��3���Ǫ������z A����`����O>���/pq)��X/Pn��g��_� }��=C��|f<��Dp�����hS�zݓv�0�xE�[�1�Y��5d����-f�n�� Wb��ۭ�����h:aÁk0�,T�XSQRiU�M�n�j
5�]�H�Ywrbg2\ڎ����'�TG��{s�f���r+����ꤎ�-�x�����jG��{�C���ҽ�Op����Oe�x�A�~����`�w��z|�r����{�6m�Ϝ��\�=����}����"=����p/��և�R��=Gr9���NG��uǚ����`?G��1"<ǣ��B������U��/9ߜ��m�ǒ>ɽ��]����}.��^�ޗpCݯy�rC�=���y�:�$83;���ҽy��}���t�(�f<����G��!����l���}���}�wr?yb���}w�.�xϸ��(;�����>��
=���}{�Y�����:�|��7m8�:���~������.���S�~���ܡߘ�w�<��i�ݹ|�%+�{����r�-)��S�Y:�^J�vW�M�ވ�ǽb>��ԏp�9x��8�������XK���O��O^s��_������'�h_cr�o�&J�7>Ǿ�}����׾�9�bjc�/�Rq�/p�x4`�C�����G��>�w2����/�w	������uG���#��U��F��s�7�>�x���{ޔ>�����M@�;�%�2^�`��>�:0q��O,��xq;�wr�������:5�}#׽��y���898���ga��GG�DG���k��8�f��s+�=��.�{���}���X��/�a���9�v^���A�=����bc�>9*��§����M��_H��s�!�O��1O`�_�Ƃ����\.�!x�>�%�B��|�|a����?���y{�F�u�?��rև7�����I��@G�s+1rd���(�9�sҿR��ݖ�=��q?_�O�{��汐�-�NuAW���ڹ0�V�2�X�\��bK���gAl���M�@�(ԝ{���*-�{�<�ߞ���9q��q=�-�q� Q�:�r�uc�Oa8;�IA��AO?}������.���]p��H�{�c�{�h���;=�a���o�R�/q�>�};9Ǜ�_ �C��S��7+��i�+9��O�;���~��ϾЙp������}��������sm�����ޡ�=�>�}�#���X�����0�8�r?Iט�3ħ7�<��u������#���I�w&����8�q�㯻׿g�	CԻ��yʺ�Ϻ���W��Zn�(7!�<ێ��>��q�qď��y�jS�t/0}'�pR=A���}򋪙�5�$�1�!=�{1<w/���!Խ˰߽�ʼK�}h{��s�-Wrfu��Odx��P��n^�ܿAw��w�3|�y�w���ڇ�o�;�!y���%�2S�~�컗w���!Խ������|�{�����|���^�#�SϞ>?K]ۙ���֥Ȉ�������#'}�>ø8=����7/�2=������C������.����C��ig�NgR�}3��]��>o��<�μ�y繷� ������;��~��d�_�'�a�{��b�I�}.�w�!�z����K�a�돺�<ǽ
�ܻ�-�ן|���y�Dh��`���u!GоA���pR>\��FHw��n_��S�~��q�x��s�C��/?yi���=���^���o�������m��o��Jg!<���K���C����_,��|���e�]����)��I�8x#�b<�<C#�g�5�� ���t*�iJ���!Ηz�ۻe�s�w��k�WLM�s^�w�O�hs�y.��7e���)''�%ן�w|��M/X�����f�������ib�nI��A�v���j���ҥM��%~Ǣ#ЄD{�)Nj���>���w�o�H�w/=���|���Nq�	�<�}r�9ъ���8�����0=��G�"*4lr=�<����Rz"���|���]é��w��̾���;��Қ������!@{'�������{���S>���*�Sm�'g�~��>�K��&��w7�s�C����wnp�b�H�}� j^��A�/�r��\.��x}ϡ�}�� ��!�;�G,��W�Z8���p����x��+����˹N;�r���2T���!�x=��O'h`�^O�瀥~�C��������[ַq����wǛ����vkr�.�#��G�|����8�p���X}#��8� ܯdd��׺J�>��#�Dp����^TW�쿋��+�f��<�óz������s���;����=��up�A�X��y����9=�>����J{	��|�{s�/x�>u�u�oy�Y���^aٿ��Iܼ{�2�������]�ۨ`�C��s�)��8��=��t"�G�2X�D�g�N���Q�ʋ�~u��#g�w/pP�w�=C�~���hL��x7�\ j^����Ww^���y!���H{Wq���è��#��Ԡ�ؿ�,9��e�ވ��#І���l���c�;���ߴ���d�}�ܾK���ex�����/��4<]HR}#��>럋��2��|w���by#��c�C����˓��=����W�����rS��˻�w��p���ǲ>Hu�Z<E��U��<�[Y�/z��U���XptY���}c���5��I��U��0jx�)1����f����#�ݎ�ת���[�\��Dl��u��V�P�m5������bzD��z-��_oq��>y���*#�"#J}�7]���y���?#07��w	���Aħ����K�9��O��>�J�=y����G����K��{9ހ<���9��+o}�Z��~�`�BɏB#�">�S�������n�����(z��e�dw#웓��>�>��3{�l�<�,�� ��r)W�ߒ�R��r�9ޗ�a���
}'��<A︧Sć����~#��O��u�'��rC�q<��}��z�=�c�<,7���G~�\폡�=�1���=��{�@}W���_�~��:�M���d��pw!_J��C�����^��1C�=eA�Vw��|��{mO���{���8�n�}����$}�2W�w��4/sǻ�}��pd��P�AԻ���O�������_ˎ��(B���*}{�l��&`{/����`�:���]F������>��� {δ��w����=+�p��e��Tl��_k`w��tb�ɹ���y.��=����$��7��wyd�F�~�Ϲ�=�0���~�5�ёUs6㾻�<K��� D{�s�P�9�`�ܻ�tb?K���+�q�'��)���y���X��>��u�/��/Z�y������^w���`�0�|h9��>�K��^�ϡ�}���X�r�j�G�㎰7d��s�˹N���]����^��/5�����:��DG�DG�
} DPS����>�>�HI����uǙ�9/�b���_%�����s��}���Ö�7���Ϗs��z3�z��ʆG�\���F�/��ڹ�lh1.I����;���F_�ٺ[���2:���D-S��	�))�h���au|��1a9��'o=u�<��~=���u���� �̨�@*Ҡ{��]yϝ���}+��~^`J�5)�i(7/�S���!�^�ew'_k�P�t���q�����P>�n<�}t}Ʒ�o�vx^o�}��;�6qo�C�ܧ7ҹ9[��W#��_��<�	�;���hL��w�tq#ľ�.��w�Ɉ���A1v$���ي5�s�A�{���8��p;��q��9�y�pp����Gq�F@���������_TDA���l���DF��y�.�{�7]��q��/${�����Cfb}+��p:�gP>�ԽA�O/:�z��8�;�:�#�~�����=C�w��0�_�NM��{�����=�����"羴=ڑ�=������{���=�ԙ)���7/�W=�>J��l7����k�tR�%���>�{����3+�^0v��~�(_CN/y�L3�������Vri��7۔wl��yU54z���Tm%���X���ϸ���hy�p�dQ��V�3�o��	�Zޗ;X�E�cc[��[ڎ;�CǮ9y;z���Z�xl,8$.9�
�s%�S��]�ԯyu=���Ũ�aF
�g�x�W��� "�&��-y&Pu���]��J9OP�ղh획F�����~1�~6*T�ȑ}r�+�t!��sD�)�uH���9"��zjM���q1ׄ�򰸯�G���@J�F��B�ZAi�Z�J �
������
B�������� �y��p�Ѯ�8�I	ـ�^�Gyzf]�Ļ��>��8�V��5�<ƀw�9�����#���,�ߕ.t�9.��|VMA@������[�%b�9����++�J��]�_�Uµ9"��ux.umכre�Cm��8�vB�Ő�J��ꞩ�u���Dp/6�[y'L��s��ҝ̻����"ҭPP���v���/q�AMZ��M�
TK9����uի�"}�(Et�ao��z�_M�lieї���sEc��R��<����s�S.��V���T�:^O^;�]�E�7k���j5x[7H"��r�]�"�oM��ov��|�V��_�)ݘG�T��q�P�~�h��Q�W�Հ��o:�Ԝ�9Ի2s8&ϯ�Q���v'I���1��iw��7�q�Q2�}�J��m��E��iMY�4�_}�g#yӏ\�TtG-��}�<{��u��&�؜eC�ž�E��M�pgǅ!>X���a_$����?
Z:@�z��;"�-�
��:���Q�W�n�vG/5�↨N���xGe�������`Z�;Q�R��s8���ծ���A���e����@��M�U��k�vE���hv�&ҌWmg==������Lc�����'�n-�[{&�^9B��Q=ڰ%�,�В9/�e����qҬ�6����R��<e���:ge��l}�9-\iC������8��2c��Yt�Eq��b�Yr��8�`�����Z�]%,ێ8�0��:}k�ծ��p�TGZ��� ]�G4#N�P|�֯��۾�l�5dcpb��;��0H��\����ղ�;�ˣ��^��PU6���Lt�P+Xf�b3_l���k|7 N�\=:'���k��'���OoS�Pxu��7=}oP��\���i�oj�o��9ѱ�f�B#��6�s�g~����E|��$�I$�I$�I$�I$�I$�I$�I$���݀�[f����F��G԰V�vS��v�8�22�f��n@w���sa��B�Ѓ�+'{N�u�-t�9;�YMw�gQ�j̮�PJ�'G�Ⱓ�)��ڝ�4�}F���r��h{}��]�[n2���u^Gp1U�8��H��4��"�0$c�,�'z �q5v��5�B��K_c5d^@r�]�z�J��X]ta,�Cd�ɘ7X�8����̈́M��(��˻�U`��;�	"[���@c�؋[t�6�qp�0mb���p��I�a�NRF[PTx��n�T�;y�PT�P����ǘ���#���Uf+��k{ �����՘L��:YX��fV4����{S� �.�ڋ8j�'4C�q��I%�[�1-L��
�p����m^���F����N`lib������>��9��$�G�%��+z���V8��E�o��k�^L���i�
������U
2��Yu�'rڙ��n�l��g�F���B�[��p���u>��Z|�����7[u�%$���$��~y�Z<��=�{����y��Z�(��)Q�ʄ�i�8��uT4�.G�↧%�

]�d�IM1(Qk����AK�M �%-T-)T�&�š"
��&0�ER�s�<Ò�BД�wd�Q@�S0�=NK1JdI@�4-PU%PP��ILT�ݐD�PP�U RP�QCE^G���z><J�� �-\mW��eP�Iq�yK<ƾ����%$�2�r< 6bɅ�ز)`��ڽ���=����ݹ'p�o����L_��PUTo�>������짻n.�5�D2q����m�l(Di~�n�
B��+����=-��X�P��q�Ŭ�����u2)q�X�ebT^�+�]VК��;Y��(�-TBx�����O
��R���9Y�FL�s�:����q6P.��9m^�D;<���OR�����ҟ����2��'7���-���3�/��P<D3�tK�|	(H-���]��Q��p�VVLQ@���]��.;I�:�y�
�+�0gL����c1���]C�[�Q�XE0�%�ې���Ry��>�;�ckz�|'%y}!p���Y�u�CM�i�]C�)Q������v_��V��0��3�����Y��].��zTa���د���p��K9S����3[�/4� �X���	Op�͸��7�Y�v��F�F�_j��K�
w@!-��1I�ȹ�E��v��#�3u����VJ��Dz=�@� J,#��s�hk�u/�+�4m�;[<*�P�>3��ׁM�sk�{�{�s��CW�d׋�Ǟ1���x¥V���ũ�govQ��T�Lr`�lt'�l���U��\@"6o1bgt�VW8���F�0�u���Zor޸���"���e*˙ծ <r������*���s[���n2*�6hGQ�ѩ�
Y�ݝ;y�Aĵ1�E�8�q������7;�%qa�5�.-�ҳQPr�.w�b�|H����q��\b[��E�]iZri(���	�=�Vӣ�E�ב�(2�qor(_���q����7��q�ٸ��T���;;�-�t{����N弄]�>��/[)��p�d�5y{wRҾ�r�glg���\�h}��qb&.�,ۢ�ȧL�.��b��S �]����4�4_����"귆�V}�ާ��N�q8+1�šM��Z�NfAF�:)0�
��v�]��˘�u�;�r��W��DDOu�km��1�;���v^�<��vJg{by�[]ծ�yYs�O2��q��3�lʇ�{J��.�� �� �����T����U�4�|u��{ޠ��$�w^�K��*t���J��H�r��\��p�2�u�Ꞥ��h � ��FJ�k���P�g�����j�=Jh���)�K	o��l<�ʔ��9�U���Мq�.�lŏ�˾뽮�c����9o"�ֳ~9U�Q�N�(�l�ou��;�7��X��ћ^	jȬ�q�]q����r@Xf/ԣ�=6����_�8�Mm�V})����x�^�y�*[N.�P�j�{�r�=5l��k{����騼ڀp5�o�F_���O��l:���p�H�!Q������~�mO�M45�b ��
�,�vo�~IKu��9�ڵ`����0��{�v0�.jA�Nj�"ڋ�tm�q�*�w^G�s7/�t�K��=���=�{-l"�����*7�Om4Է�'0�#/'��`�rbާ�)զ�1O"�8�x�8���+�G�s�@T�h����t�OZڵS�J�-����J���>:��H�[����;���l`k�tn%��^jF/y]=�)�l��;�|V�6PN��5��]'�S��Ƨ����S4���:�s5հS[s�� x�s���z!����T9Yf��cN\$뺔�@�0VM�\j�s���L]����;�y�^G���o���W
�NH��9���}Km�b՝h�;S��^��;!�e	:a(Kwo��3��T=<��̐\8�=�%��,����0-*�PP�o����fQ	uC3D���_(����cn�ޛ9�0۔��ozmn=�E���i��T����;���b���݆�����,��ۺ��L����pܝ�,.���p�%|O\��o�z"=�X����b�}�����1�e��R�몋X+H�vb�KB��KoP��^t���+!m�Jb����!Vˬ�kL��q�ѕ��*-�i��;�{�*�f��ZIޛB)�GEҪ�s���OZ~�*.5�:��?�Oy����b>��Q��;k\1[�7JN؜*޶/J��Z�(���l�˛���N���,Ȧ����湻�,�\S���[�W|�5X�Nd���ibt��!tfB�*:�W�T����}0�V�XGQ��8O�V̪�]q'�F�.�H�vus�/Y�^Kz�޸��ۯ:��#�ٮ��<G5�7{J��gX\�g3[����y7�8{��~�p��z܌�4��L����TbX'��#�Ija�mT)�t���h�Ȧ��BŦ��'�6o�a�Z��2��⻺Z�F5^٭�;p��B��k3�J���\cn��k�H]d���yz�d�F�,�=�� ���%��.�<:�-�׷]GkwF���miY09�ݍ����k�j��]��xr��ktU{�+��D�;7L�W���m#����pUJ՚m��&��
�_�^�}4gN�#*&�Ss8�
�F�瓥�Uo:����>�Χ4�7(P����C�dd���sג^ݴy��}� N�zU!?f��1��;Lt49��w6Ɍ����}=�Ї�iw7��q�r��0�7Ɋ�����3��p(��b+J��}:��L����F�7��)b9���@����]I7K.��2�0���ϫk��zQSy�m�x��ç�����엽%��-�-��j.3�_H�
����l�[r�5��.0���H���,��=��Vm�odI�v�.moK%)���"&��c��}�<��
�/5�v�B�z�n��J}Y`��V�up]M��l�N��1�+2��W����J�ov5L����W-�l��DW\���R�LmB0�Ղi[��1ˇ$�VQ���&�v���s�(9�4;�n>E	Z�1X�^Q�Į���f�QOl�L���V�κ�D3zy��4�=oWz㣀j'kP�{��������#��;��VU_<��d�w�'������u}�VX<�`�q긃�1F8� �a(��N��+�*��4��S��:,moK��;5l���P"�w�N�0j��k��F�ˣ��S�3X��,�*�ZB�dr�s����U�|�(0��>yh
��^�`Lc�d��	BC5���S��������H՛�F�^�N�j�0;��ģ�bW�g��[��NlY��X��}@�`5��93�9�C�l��0 l�Zscr����d⣳�n�4 ދ���趶���
5B1m垵�#+{Tb���'|���x�t�r;�]5�n���M���:.u�5�k�ޏ{��'w4$�^d�Q�@f�)O�Y79v���(TAx؛ͽ�j��nΫ���l7��$�O]����^��aj�����p�ovy�NT��[,r
{}�'#J�]L��3�"��/Ī�S�Y���Κ�͠pT5ju�>aӬ:N�3Yx<�^�G��M5���r���2�z�J���7��{�3���iB�.1����\�mׂ�3�e[Zc�\Mr���}r�.r�"/�ũT[�;�C�G(M�{E�T�|v�o�����L�TC;��ԍ�+��(�[���L>C�[M�0���P^��;ؾ�V����t��wc*ؓ۩�n��]�N��'����m"�Dsa �#ŧ]��-Hۛ�QcsǖӜ���J<�hi��Y��7>O-��V���`�B
�o���p�m��N���n�r�mΥܠ��R�������O�ڊ�A�To���s�B�͢�l�ٿG���'qK��x�\�u�J諹6��ҁq����8��Kr�vjD�oP�31�a�	Z{���#�3Y�33��e<D's�����x�d;W�Mi�����3F�
�y�M#�J!�r�n$����r��+��lB��y�ѹ���c�~/g�}�nR���b-`v�t��A:W3H �n�hw���}:^Θ�л���0���F[���1�)�9\Ҍ�������gz�ۛ*�fנcD�*� �
#4�"�~ۧq��.5O:��EY-�,����M$�P�ݔ�7�:l�+�AU��VO)����u�Quۛ���9s8�ǅS4D8yx��_D/9ȕ���c�5������^��hP��9�Y?�Tv�/$Bx��he�S`���6��KRN7�����nuG�ʱY|���8�9v�3e����>�Aj�8��G����NAovRNU(�K�va]�vI_z=�����K�6��z�b�E`� �����Ư\J��30ｚja�`���8�R� ���h"%��B��/�L#�$G�C�ג˶�^��8[�/��pm�.0��7��D<�`��6�ı��11�e� kyoX ���!.c螯�rd�[<���m����;'
Ůˠ\ɞ�W��eV�Z��ā�%qb�l���;��˕r�y�X�%��:�7]\�;�򭃺��Q��,7ж	�O�a=qDk�ʹ��4O{֋��0N��V�D
P�Y�M!C�^�N=2�UC�1��t�Wϑ�i5ջ8�M���{���U�>m��|��R�g�.�.�b�s����p����].�a�PJVB>5��c���٣$�	�gq�hz�A7Ui���̾�yw�r�W��s	���5���R8f4��<�1�3���(d�М��8=HڏJ�fnvWTw$ט�������y�.�֋�'�X��a�A������5uE;oW�2���9�����.ڻ-�\�fR���v��.o������oTL��y�'t�L��*S��I�P�����5<֭w�1�|z�ʗ�ʆ�t�^��vN� ��1iq�O�J�8iش�Z�i��r����{F�@�wl��Y�����uV���C�C��Xzj���i3�VL;3:2�)x��D��b�B���}̮L^K�oq���_,�#~A<������-`��VVEL��)(̕��
��S86I�N�r���Y̓�E��'p�_fV�C�6�*���NZdsLR�j��ps���bz�\�ݡB�mA��'��'��1B�JK5�[�%|j
�,g��vsOϟt9ٴ�R�ʇ&���m�w<IXwб*fsh��x�a[�)0���\tj{�ޠ��c%X`L�"3�����oWK�}͵6����[�&�C���l�;�71)��+�h�Oe_)ԣ}�7��Mۛم��,���d��w��#)Ld����}��A^`�h�Z+Q+v�Mم�u���i$�I$�I$�I$�I$�I$�I$�I$�Y���*k\�Ʀ]Y���ܾI2�/�)Y���˙��>��ɋ��e��]+�;�	 �J��s�]N�xL#��{ښ!}�mi���J����1�]l3�ͦ�����Nr�:z,yX�"�^�of�\�R�b�̅��=a��R��� �{m)}���L�4%��V���d�q���q�����Dɇ�W\],���YIj��m�)3�K��Խ;9^V��p� -.�+y�4����O,�j
V���۩\�ڤW<�_X2%զ�jlm�R*b+]�C�æސ�s@�v�#�,Rx�=���48����gq�����ղ�TY �us[�g�eI�F#��g9p�нit�W�c�0��:��"udk�R��yF�i��[�K�쭁�}�lJ:�G71�G2%�ör�әm�meG����bG�uKP���'��.r�/Aa4��7�#X�&�uuu�nS�/�{��b�/�Yx�G\��d�Jl̃�����ONgn��[�zn���q$�qIV�N?���1��� @� ��^�0���a1�s�AP�Y�HR4�N��N$32��[1�!� ��2���#���@�1i(����L��$,ĳ ��� 2^�Z�!��.�)nq8��996aB�EB)B��+����!B� ��2������,��% �4�49�K�{�S�"suC�g]���v�M̅V�r�N�m��|Ň���}�<�$�\d�j�����=�z"���f腆��H u�yK��XC�0��8�o<�%�,>576���.��Ҹ��J����r9����>.���ᇴc��#�Ґ��N�I�k�<�u�rsP-�]L�8��E��p�G
e;Ю+=��=���N�n�֪���a��oL8g�f��o�I�2�<>��P\�!�(�v�f��P{�
�,�CP]:4n�Ftڞ]Qþs/�҅NyJ��i�`ܼy��I�G��(H��(˜���ͱ���W��<A	yL2	�8Y�q>�ID��s|db�"���|+�l��f�����RȘ�q1���6�Ǽ������=�6'������%[f�-��~��,mӞ���r�������;g%��/�>2��2֑GeQ���U �w������P��k\b�۩hu�<;�!�^I���Z{��J���}^��:uuN%���݈��C��K����3��l��䣖�N���#����Wl�qbh�u��_V:Ի�9�dș�ʅ9%��XR��4XX��)b��R7}�DT�h.��-<~��{Щ\R�,�t6#������l�Ky��&�l/��\fU��/��I�4C��#o¨�BF����4F���Ӓ��}��;<ѧ^��\|*eu��qG@da$�0�5�����)2��c�S1h�I�
7�$�OgV=CDg�Z��o[/�>$��E�P��g!����٢r��Mgsa$��ёaX�����׈qǎ67ls�W��3o�2��^����L�T�=4;slU��X���g�(����΋������x�T���|7i{:ȸǷ�9�ľ[�Κ�|�j��Q�~�����{�k���zR�n�G��s����\�c�g1xt��csU
�ʂ\q ���]�J�L�h6t���9�TF��K
�!�tw4g���C�Z�cm�-r�u��A�L�̡�f��HHN�:ك~�6�QƩaNQ�J��-��#U���3/��C���+��xu4�hڙ6�T+$���I�e\^Mq��g2�)���B1�[�ٯ�K�f�h_VG3m���+}ȶ��y=h�Yi�rı�����DA/O3�]�L�͋ޫ�����$<�]����~�O�[�Q&7(���Y6��O�����$�d�k�X}��g�^\.��
p��O$$V�x���.C����3�`���#�]Ѝ�b:DΏ55������q��'�����������ޤ;�i�>a-ˡ|�@ �"&��:�B�K�#����0��	����.�|h��W�i7�L��fv�E s�m7���/�8:�(1K�=��m�&en��9b������[�E�Z҂F���s�P���j�^b����\o��	�v�Fk�Es�8f1�ۮ��h�C�x8���|C��Z�f�.�����6�MB8`��@��Q [U#n��/[�'����=�UB(�7�T��Cܢ�U���������}�c 2ԉld����Ŕ8j7�A.;�8E|h�#��Ө_0�{:�Z�)(	�J#���׆�����|��VT��*M}��������AFw]+U�O`�}���>dn�j��"Lu�9ÏVT]�+0K�,�;ѼRu��~}_U|��q<���Z8H?eF9��`�.f�Sza��Bk�g+=�g<՟��T�{.w�j/�Z]eW|G�=*��\�zɶ��.�1΍K��;-n�wA%�G�M(�W������a'��5�-�SK����7[g���%d��>���h�cD�N�Wq7��A2��3��6��Lrިmֹ�0�K���/�٠B)s��>>�q.0�O|y�ڔ{>��1N~	��TU�]�����C�;"�x�	B:�H�-ʸ�'�������҂�փe��1�6P�: ��.�������wuK�o��5+F�MfQ1�ES���ldEϝ'q�%	`��S̜��Y�=7ye�r'�ܣ
��,JC�!�GL��K��.��-ѕN�ט�M�+�m[�n[��<�8�����@���'�p�DEex�2Py(v�+P�7=���D4��[�����v)�r�#:�o���Kg!����<��8̹�v;.L�8uࣅ�C�>Zt������u0�x/�+�Ss��X���[�O$l��+�z=��=	=���?-κt귭�i�Ik��;�o�p��Y��_"=8d�5r|:����>��S!���>�͑ƹ�4+�z�4z]� �^��0J�������w0�~(�g�@����h�*,Üڴ&��b5�'��a����=��>/�G�R�|�/c	�Vx�s�n4Y�t������}9K��b���
A��_��6F	��WK��2'O	;U��'WU:�cG�R�uG��D��ê��X;Ċp�E�3�p�o�q����
g�Rر�~j�j�����"�.1M���g�d�U���xk���ͮ��!��=���j���T���By+�X�l���&�:��(�(j�+T���=5�]�\�{r����qb�s�Tu7�J�����l���OV��V@�f�)�����<A�{l2� �ʥ�iخ��`�*/��mۂ�+HZu�3�St��{ACLr��0���!��u|��u&��:���o�Bc�.�w,B���ķp�n� ��s����n�LQ��5���Y�W��؝���1ݞ?�^|e�du74�"�V�U\�q��y\��w��÷���t;�6�$e3�w��Mm��yo���N]l�^�/mj��Rt�]�E�'f�Pt?eS>1/�O_ʗ?��;Z*��ȗR3���OE��
�ۮ��zji�:�yF�\��a���a��Q(|/_�}haQz�I^�����4����GEu�U�!d�u�YA�VeFb�����w�9���F梯s�����o��b���U��c�*F��M��Y�=�r�zQùNR�P���:IdB�5�f(,Gr8Xyt�}��Ր�J�2��E��ֱ�2�(z��(_4��
���eu�����k,�e���p���z��<~MҮ
�+�8�Bqny��c;3B�+`�?>��+yx���c��(o�<�G�������
nz�LTHz�������f�n�i�����<��7����SF�dj�bm��a��&oe�ԏ.n&�y�l��3����=�r�v�oJ��䊍2�C�'Sw�!�����v����<x��G�ɲ	jRЍƂUH��e'\A|����p�3��F<�����u��\ݾ��f�1��\՜��s�������Ƿ�\d�J���i��c"ޖ
�Ц\7Q}0�Xa��T�q�#9�醥�N���nĮ��Iw���$?}���W�8_ծhZ{����^ڞ]�C�����\�ut�����Ԩ�s�K��T������v+�Ǯz��p�p��v���j�j�i�*˥	$�&Z�V�NR�a�ƆG�Y���o���t����ZS�pT�so�C�{�+�:J4i����(is���,����=L.�<si�4��ydfyW�[uC9Ԁ(AN����eT�����+]!�LM1C��z�m�v�	\l����0E�I��Y�zDj�>�X�K�Zg���)x?�C۪��zYP˫���N�]�F_=9�F2��������vuS��+Ƿ���yEa�]F�9��=#�3�6�m�u9V�S�Iύ��nhuv҂=�w8��w���p��z�_SN�V�{���Z�G2;�β�fઐE��Hiq�*8v����F'��P-�9(i�+���������"�58;���q��:�^Z%�.�
c�� �>�����ܞ�y��C48I�H�tʱ{=O�ZQi��E�.�0r��ƽ�{uMr�6V�(�l�@�R%��=��a����5��<�X2�p�ve�Md$!���4�*1M��=�%B�*�>4&�he�3����-�L�w=u��~,x/�fp�bd���fJfɦI�.�Ox��n��:z�p`��=�B�**.�� ����.ñ���x;iE�#V����K�:X��5aQi~R!z��Ťt���L�E�+�t讨�i�!��ku�"�����F�^���f�\:u]��_1ԇt��:�Y]dg��V�����h/�A(GRDqK�QɎ���VV�y���.���Þ�$j�PzW�E*�2fg�y�/y�<AkQ�舞�x���eJ�v��ID�IdK_M�|e_$��էq� �}ձ�F��N�[�� b�����h�i9���W��˘���z��U��8���Oc��f�!<�; �]�	̃{��6��ۚ��Tx�E��ZG�W�[�6v9S�m���4�:�,
)V�NL�U����PKN�l.!֖:�C����֙C}.y�E���^ڲh��>J�u���,/r�'2�z���xm�T+XLC��'�5?R��;����[�o�4P��jHqf��������f2pZK\�y��,P�+�KE����,�z!������׬q�sdpu��t��e�H�>w�|<5���mR�rt��_a�|�s	1*X,���w$r*,�ԕ!�k;�2���l����7獝=Uզ}�)\@��a02T�E��Y#�9T0B�ꜝ<Ԧ��&<vͭ�?}H<�v}�)q��r�ķ��#۲Թ�8�,�n��Q���d�.b#Y�vG�dZ�&C��8���B�DZ�	ܱP�1���'<z���y��@�����2
�������~L��Y�K�u��)���JL"��o����R�I���wa���q��pJ�50�9n�|�ǰͺٺ1k��.f�ψ��;��WT����������+�n��-������j�V����c��<�Sd0<�Mn��㳺�n���f�5��Py��������"���F�|�i��_f���q5Y6H3�B2��,ԶK�v�;o��
��U�&�b��gn��IȰ'�C<����j��0���|jx׳�!<A�=�2�R��7�M��9i]�#�>4ze�dm7�Uګ[���W��V&�
�+�s��eL�szM�u��BD���O�ty��c�*�5�z畡�5z��G@���~�^~0�80�*����4��.3��;��#Ī9=Lx���T,\��=E��u˷��Dk��("]����e9�0�{��Ts�9�X<BS�,'�� ��ߞ���g��D��R6��Q&C�k��&7'�1����
����G���n�:��>�@��2OO]��~�g��d���xh�/��TB���o������P�"iV);Ǩv��!T��۷i���(C��K(���Q�.�,�fR�97�q��3����b�Y`<{|�2��֓�k6�����'۲
4yHo���"D������)����=ZWu-�t��ਸ˶���/7hm��m�(�S$8���ժx�	�g
��mh�����Nga�K�)'ڹv�;:�������x�awow�0�]O�&*��[�1�:�`ɗ�]�DD���z�\�S���y��ݥ�kb�9��;X�V�)a�sTN�Q����X�d|ݻ8�ȷYU.&vP�����pܔ��f|
OB����,ü�0��*�%V�8��� ӓV���%D���C7�}@����Ƹآ�ֺ�q\kNP#���vu1��.��zuWi����jԽ���5�.�Ig\�v7��]��/j��gZܤ��L�j�
`�`ջ�դ�;��:8�^��ջ2Q��"�+77yͿ�8�]vV��������c[&^�X�a��dbB =k���i��t�tӁu���2`��_�ڴ�i$�I$�I$�I$�I$�I$�I$�K���PE�
��R��uݐ����`�@�N�_�=ٮ(\6����rh�vG>���<��ݜn�Y�-
v�.�W��G�W8�HΡ��_	���3i�cg�@�[�7��<7�㺝YÀ8��kr �R����T{Cҫ�e�l�U^Bn�bV��J�'\�#g|Lz/��ɥܱ��萦�6�eu�9Ӂ�DX����s��̲��e�U�=3g4�5x�Rl�/(���+0⿢;�T�H�;ўJ�Ju���w�۸عuR�n_t�o;p�or���W��h;�gK�$moh�̊KҌ2�k͋N����!'��oq��nl��m�X���f�Ȱ)����:��j��xy�l@gK����u����+snm;]{HQ]��p���p�Ծ�ڔ<q�MZ0�{��N5��wYK9��kv���6v�B;޳5�սrg��%�)Ź2A��;]rgO,�u��F\<�>D�mG�};b%��S9&���@�݋e#{��V�Gwm�V.3U��eg���A��3�ĳ��怣I.)$��)_��Ԇ�3�$���C'!�O � w�Ek� =��y.@q�}:�Q���Ɠ#&�"\�# 2���)�Z�P}*e�Z
�(\����(k%��J(rr$rrJ\&�p���� �u�9>YQJj2r�ȥ22;��^d��1�2�2Z$��B��_���A�i�ܧ�7�x%$��,��s��Np�5k���]&4��J�{����\{5e�Xyj�"=GZ�T��:�����M����(�da%���׹���)y���&�yR��흮�h���=�
B|8c1���o]2����AbV_�;������������p�wF�>0}����WJSd���(�������!HO+$���qY�驹�*�)b��,�1}h��`͸�����wÌ�h;n�E��E�=�}:�p9��vt�2��:�F<�K#��+�ݾ+H��_/�E�Ǩk���P�����b��c�EP�ieⵍ���8i*~�P�^Jgܧxݑ�^�3,T��� ��v�r�]R7'E 8,8�~ f�;�C¦�q��7�ґvN�?V����G(�("�Q�4Ĩ��tij��~����q"q�g>���I'Y����1�Q�$�ШW.務ED�W�/b��Yu����~;�(5���^�s�����%�YO�YB�ا���gu>	�-+��%3{=��������H��8�!݉p��K8�_q\�Ó��]��VPv�w
��˫x�d,�����6�7S����I7�_}/�n���_�GS
�6�!���!��B�{�>�AQ(xѧ6��z���>O�5�C�Od9`��=^;ֆY�7z�_x*���" �)sv������x������B�S��8sq8C�!_a�<���|[�S��q+�;��s)!��$��B!����/,u�L�[N�تb㦃rOMvv�����LvB���_6�2��,�-�.�e5���t�fuc�&]�ê_t����	#���	.�L��P�=k�=�.��g���p� �zR��u�y"� Ǉƽ��M�P2�^�S�&�W�>9��ݗ<w;g��Li�m4T�J,�@�R%ce/���^�z����Υ��2���^����P�+�PަzШ��l��nf��},h�~f�P�u&��s8wHꕳ�3�t�ȼxପ��G
�8�J�v��U��S�����0��th��q�:]���ʌtΡ����+V�oE�T�|}D1��f7"o&�Wu	�gvCH��(�K4Sݭ��Wȉ:�h�L]HƐ��훱���(��Έ�em[��ȱq���{��Q����x�h�N��ٓyZ8\J��Qp���Xts���N~V4W=��z½�~se��uém��PQJ�PZ�K�D/9Ȓ>�<��S`�n���8�w�T�T3/U'0��ٜAҨ�!��F�y�k�r����e���~*�{(2�4!pWY���x'1����i(GI��U��U��7��(�6:9Q,���C�}��e
!�; ��P/0��$�;_q��O��B�yQ�jϭ��c>E�agb���q�)���⋅��<G��$&4M&����B�tj{&�⿔����:�'Ք��{�$������	�)��J��OXn���y5	��dYf�ߡ�
�w���]��)����N��D�Tഖ�hwT�����t��m�(���{� �oZ;Hiƙ
�|z��>��TG��7Rz]�;O���4p"2�E!7Y3�����9;e$���*9������+P�v�'M����$�u�.L!"�_4&8�:QT�)(�x�{/j	�|��|f]�Z�s$kV. ��]�_5�_H1%'L�\4~c��uƯ���!�T�]Ǹ�3ɋ�"�zo1\W�s7�X戧z�gL���e+�����3U�1N�p�z�jwܯ^*�P�sH��vcd+�6k�\o�XD��8��=�u����^]f[:O��A�6f��J5Y�qC��+��e����^ي0���v�pG�P��b�g� ���{����p�*��OhN=�K(W(��R�YR��W	ݍ3&;��v:���eAu���1�yP�%:�"�\>�,�"�;03z�Sԃ>T��`�;���i�{��'�J̽ĭ�r�k�1\�I���W��6��N��|+��	�vZ�/$"'�c'�F곌X����G�X������;S�$���C����E��W�Z�E��l���.h���+i�͞�͍�-��~�� ��<��4��E��ebV�,���b��$�J�l9�W2����G� �=�ER:���ߢJ�X���4�aۛ���j�i�D�ؾH��j�;�8�^�j��yjh�Sx�5m�n�Wj���å/�Ф-����b�Oۮ5p!�vU3^Q/K^��P}���",~����g�6u�7��\��Ų���ޟmw�	]u�@;0�6�@��D��]\����/�GչPf���ሞ��+�`�x: a�ص��HEQ��b�X1�x��y^��U����K�"�F(FP�48&z������p_U52iF��z�ɞ1��p�V��5�m�8�򺜨��4Ί�AJ�� ����Տ�1�F�]1�[hs�XC�3��o[/Ư�ȓ�����Z��Un�{΄�ݣ��ڰ�S��*e�6U�ᬟ��v�8`�l_�y!u`��-��6X,�z��Nv<]pΜ�ŷ;,(��������G�s7}�jJ͔}K�`����ȸǷ�S�"��ޛ���j�N��q�i�v��ƨ�TD?]S�*;k��4�tg��/�#v-^��O����1OR?#����Ӄ����{v�y��ǝ��>w*�ӯ�����J�t,:�܌�5Xw$�*N�t쾵;E>�&	�T�y�7%�	������o��J;w+��'z�^m�_�&�#SN��u�W���ᄿyRz��;<<Z�q����:}0԰�m�i�7��J�i�K�]ufsG([�F�K�Tp�Z�&�i�*�(F��ʄ�E�｢><��ܲ(C��A,J��D��c�qL�S$�d�ܢ�MR@��D���ޱ@��1[��G�qc�JP�D�a)��*k�Ⱥw( ei�i���/
�ţ�^88]?M���[���K�~��t
�Ά|}�Z�㔫wy�f7f�r�z%�:���C"�0�呙
��۪T�Ui.�F;`�|]v$I�iqxP�~��<��М!�B�Zr�����T��0����)���դ�Z�P�k�9�pУ�-3��hJ���a�8�fW;�>���5�ǵ@��C6�lh���>������1�����o�gH������y� 3��*�N�҆�.�N=>u�\)U�g��y��u�T.���B]У7��;�M,��|1ǄW.o1���Zy���E-@P��2=�h��H;��ʋ����#+k&JW��&��%�1ҹ|�X]�GRβ9,�\qJ�ŷʌb]��{۷�{�F0{z�MC�<��*���\l�[0�E-��Ho,�������@������|t�Lc�3����Kc$vK�_Odr�a��/3�$���N&H��C�Uq�L�[�����u�z&4pY�^��U�\���;Wt(3��;�C"Y���S��_���p�J�������=w��9�^�����F�>ʹ�S�6�x��F&p�)}���z��f`�};��+�~?o檕�
����"p�x/�ќڕ��kf\�W\#)�Af�s�C���� �Tp���뷼r�W.Թ�t�o�i��a��t�F")�������XS:�>�*|���Cm�y,��f�T0ި}��e
!���9:�3m�]�mT���c>4i�Mo�����/��'~g�J��i�M�l����_�7w��h���������P����^VV�,S�V'��Ƥ}}9ۭ�X��v����pJ�uu��C[1���ugXGu��gO_.ӹH��_DG���\���q�)	 �����  T��%
OB�f��Q�ϑ����)
�Okz��C;p;�r�x�X+*'�P.����u�^�P�'��ؕ�H��V�{7�ĽDT�U�g��\)�t����M9�i.�-v߆��Ì_�ۥW�.�e3�@�z���
!އǴ��ͱ\/���2͡i���f�����VT���V��_Ta-|Q�Η�r�H�TY��m��k7dwv��}n4=xu*YJ�� �c����3ٹRwX�<�ͤjQ�L�h�,��fר�w<�Jc^R�x�� aj�&��3�0_g��u�PMy�%����G�{<@v�+>t�fƲ���V�93�C��"�q�}5�/��P��b�G�Vfk��~r�l�!7�;^&2�[e^��)`��INGJӻfLv#i��u�ܬ٥��"�:�&t���>yc�M�}|&D-�e0RVͭ&��Y*CX:�U���n�ܼ�:�i�D�� ���՛�M� �q1,�zWHd�Y��uAY	���ړ�1.X�~���c����.����o�v��/�_WD��J���Ea�zPR��p������}+����s���p>㙀��״�!�c��xĝ/jՏL;�jr�|+�ɫ~�כD��( �m��U'L>&.1�G���C����R��h�06�}PW�.Xb�l��LH�\}:g��Q���(.{1����s�'xo�����.���WE��m�<�^��<��*��}m�+5�}٭�!9�y&e3g����d,r�m���tthR�h�R;�E�P�0oY)�S�Q�"���^�ɤ:h����:��Y��p]�خ��ܝպ���pUyd(8�����"�^=�
�	��A;��䕛���l܈"8BtgZvj/��X�/+�����K�ͼ�Mm+Op	��ۆ	yb��Cj��89�3,k$Qg��%�`�����ר��m��.�E����M���F����ݦ�F\pD�]�/B�) +��/p����_yzP �{5Wj����c"_+��:+�������N�e]ꩴ�����S[ՂJ�Va��oT����=
`a�E�!@�%�R�K�˱`r��K���W�&ږ��ب�{�L�x��! �Y�|S|~ceԅ`������ը0/$)��o�{[��o��O"�z�p8١�M����,�r/�1�֎�=��C���A�=9�ɷg9�=�mB��E�1�Q�>��v�E�vp�^?���]�r�y�;i��U1x|N�'¯��j.1P{���yŏb�ˮ�yh���Qa�P|��8���.��nI		͖c#����ڶҦLlk|�W��B�4�K�C,/>-\�NdS��Ov鞾g�<%�9G��_I����\�y9����j�'������|+Ԟ�\Ƚ�|����Y�x���~<hl�ؾCb���r�l@b:�qW'��kC��!N���,��˥�����Ǹ�Z��db�1���.�_W?E{A�3Pcd64�]lMq�^~��@���S	�%F��9]+��l�bT�N�T��۝�ܼZ�k���'�[(I���f���ࣄwd�8<�T�����F���k�^���p\q"��Je ��7d0;ue���8Nd�\`ӥ
�9�߅N�������*x�q`c�W�J�1b�ڮ�B��V3�ά���k��Qmc�3А��Ԥ�@f��۾9�l�m�3�:��a�6�ej�SS\�Ạ�.�i='Rsbu�w��]��("#Y���{r$4���B1�A�gFئWW;
�`	.�y`�!��&����M�s/��n|�z�V���{�3V��{e�Q�m�\o�Y� t�7\�H%:WK�̬K��~�C�����	����q�ϙ�]�����3�������b����ߓ��99V�[f��-at��uK� t�/�8#e�u��I1ٗ(����t!�ޭ��+j�5p��v�=k�ʇ0mб鯚[���֮fP"���R���F�nmL�c1fP�&]7 ʅ>i3Z�&%�ʵ��X���*!Z8�
�;��l1�#���ׂ���J��]Q??2�I4�I$�I$�I$�I$�I$�I$�I$�If��3j���N�x<�Q�����ϴ^����M�����nQ�ss��q�����w�5��Rw74̩N�scs7p�ֶ������j �Vw�9wZ"�;[���k���+ߜ�]��ݤ�Oe3&�J���G�F�åMc�H��k��ԇ�^к�'s���]!d��:2�8��At�0�G�;�������yz����~�VQ3l���-,-���j��Kfj�2������8Z.�z��/�\�e���KR.I�qp���
]�G��bx��<YK2Fk�;3$�}��()�f����g��oKT��F�]�RR����OAʋ���k$�4B� �N�eNѻ�6T�G����Hxkyī�����&s�Y��c�Χ�J�������gPެQ]��5�E�N,�A�XTՆ���niē�]|^�J��\W��w�����6Zy�6��)�'&4e7�iU�E�&VP��P������]�_Z���@�:Q t���PK�	f	�K�\*zf�!+�F�'Rގ7�(IW$�%"R� y���=.&Ǽ j���JQBa#1��cq�25	�T��
�Pf��e�����H��)�$�'$(i
ru�5d�eE�dOѣQ�K�I�d1FaS��MXX�FfY`eqΎ	����ɤȫ2�&�}�ueS�dSf4dW:�_c��0�̬,�
�,����L�����2l�̌̃#&rr#,�,�����',����*����"���y��׹�x�T�.�qo�
�i�{$]�A������mu���A����O����Lr�Qk�����sG6�����T��ü(ׅ�j=y�v���
b�F^W�ғ{ۓ�\i��ń��fvf+�RԨ7�i�8��a�V�b�=#�b�0x廕M9�r��Mh�'9O"���t�ؑ���\}�a�)Ōfot���-����
x`��5�`i5������B�-�O�����sg��v�P��i_)���(̉p��Sq��;�7æU�=O�ZGYs8b�̬Ǔ���J�C������A���E�WJs8]��DJe�w�8�uv�B����ny���7���l\BƜ�YL5�L<஖O̥$H���]F�ۭA�tMN84K�uu�m37Uga	��[�j֖Bed�[<b���=B|�`X,�g�o�
��Ӯ,̘��m��ݚ��=�SK�ؿ(%��uB��E�4к��r�͕���dM���c=w��;�\ʖUh���uV3�XZ�(i.�[�� E�D����Y}��ޤ�\颵oS�w��oS���v�Vu���[Qs8�S��3��9b����ѥ}�����9��g>��u��u*�c�4��u!1�<�c�p�>�+�>��]�![=^�����?-J�Ǭc�9F�8�!p���u	͈cNj=3ѱ�x�M��ЃU�)"!Q��{^J�(f^R^:b�LoM��P�9�%V�k��{���h��#ǳൠ֭-�;��^����Fcrn���3�Һ����R�m��aF��G�'��Ѭ�VMc��2�Z�y�gC�ۮ��������B_O[��N��x� �Q� !�1�����wgXH �H����E���T���54&#���S3r�>å�ap�L!b3f�#���2��X�8����v�D�l#9�zf��Ԡkqu]P��>86}1f�f����i�Js�T��QkII�u{gz���m9���w��(]������	{�,����{��ۖD1'�Ee��	o�'J��i�x�D� H�0�eÆ�wt����dP�Amh�x���ȱ=$���ʾ/tc�y�+��3���ʝ%�׆��%K�SwKݩ�S+�k�o�y��><�w���D:9����s�#�4�CBɌ��O�㵏)J��h���K�=���k�k���Q,�x���ѱ���@U�1+�X�U���;w�����Vz���/������f���G������L����O��E��� ��C����B����B*Ѵ����t�z��] ��U����\��0*&��j�6Hs{d3(!��`L�	E�`����9V��4u:U7y�b�ue"G���:^ժ�����;��M�Hd�l�cq�ȯ~/��a���< typ���������"�$�eۋ���ְ���&\.X��J��Q D��h����c�*�P���vլl�d�8��1Y�.�:�;;*��<�^��-31=�9�Ѻpu�����#ʤ;6�w;���P�Գ�EwEF�eN���x�%_0Lhn���ʞ������u��se�E%iΛ�K�YiثB��eޒ���5����3_�D5d�RA��ut��V�Z��8[�oE�ɗʙ��lڴ*�[�u��~)�f��%l�zV�J7�/��2��\��W���S�C~P���~+��KX�B���YF� ��n3
�k����C�K��׊���U	�Y�H�?h�Z�]���c���Uf6g���>M֏E���h� �k�_[˩x�.�6`9�1^	���b`�(+!)(I(xѕNVٞ�H����ʻ�-\C����j��5[�{��u���1�^G%ܖ).�w+*Խd�k��yr5��q��>#��=ʱy8�+<�����l^<&�ث쥈PЯ����ژ\=C3jP���䊁R��sasw
u#��1��h���b.l�
꣐t���/H�y�2y�)�4+|z��Ϭ�^0d��[˷y<�Rv���|�cz(%ªÇ�OO
8khxps>�/�ߜf�Uӏ����XKL�|���C�-���Q6�;4h%��>,^�
cGp%e_�-���a���ݻ�]K�|@�bZ4U�vX�q\eP酜Kp�>���}��l���V�JN���k���t�=�n�����kU+�t�+�it6���%в��"��e<~��^���#�Sp����i�KP��i'f�8���]Cp�.�\6xFo^�X�ّ�a�B��"�eL�	�u|��h$Nf.�����{��4���¤�[�7,g������A�����#�so�GZ�ȍ��o7c��Zw����%� �L��!AG֬J�u1�;ֆE�:"���Ⱦ��t��N�K��p�.�tȍ��8��b�Lmc�����|G����e���B���L3�o��!����7�i�G:����3#���K�L�L�����ύ�5���bD�;��J�Ǝ�Q�.B2aW�}c�3;����x�o���DH�wU����g,���m%<�\.�	ا�u&%{6��Ŧ�z�B�>и�w4r�eX�6z�!:�+�!0W�.,�j�u:1��^�\UJ��
ǥ��P�-tJsD?���d��b��.�:�h�<�B����j/�P���Ý;�p��%�:�Iu�R���:����Sl��2f�W2��Se鷮�.�-���N2�f캚��t���V�Li�� ���_D���}J�H��܌�W(�|��\oS=Bظ��B���	j��.�yN������X�H��V��iV1��i�ބX*;��GX6��3JP[-��1΍�'�MV�⢢�ک�m���y@��CA�B�˫�r�P�R�mN�q���Ţ�h{�R�	y��g�$��Q��r3_D�ψ�C�y��,�{�D9�g��`��f���.�4]���GU��
��.%�ŢƎ���
j����缆�t���_f�%:�8���i�DB�r�m��%C�2���3�b륦�Λ�&���&�M���t+�Hx�-h�J�[�6x1[X�y�U-�wk�5^s�Q�ǭX�X{�L����KN�0���;򦓩��+O^��6jG�,��-�I����z�<I԰>~;a�1+<{dPz˄�Q�kV�r�(S�\csob,ԳiPnC��X$�W���#.}����cm�(�w�lT+T�<���ue�-ؖ3�k�\���f�W/Gp����"�j�ʴړ�u��Rv��P�ʈb���=SPB�Q�j-5R����4慤�L��-ٕ'��N6���:`"�1|�"�S!Ƙ�A�C�]������e���T�)W�P��u����������"�$Q�))î[�N)�n{^�+��D�a�H��#mDj8��w���B��7�C�h�v�n,�Uh���:�#)�h��"Rf�'���ǔ�%��)}��ʹ�]�>DA�c�z�lyK",O_���4z�h�DZᗇ��#����H�M�4s�xz/�˸�]b��Y��Po�O�����1՗���jȫ�[�ns��p���0�R�Oi�*�؟lp�bp^��>���^}��!O%p8t�v�vi.��i�a*�gE���R�V�T�<�j����W�s48�Z2�/g��b�N�vVb�V#"�6�:�����E)�{�޲�KD�u�/��^�y�}�z�p{nA;خ��g��f�AԪ���]wٍKj��u�;��Ɲ�.K:���Jѫ�;�w$k�-gq,����z�ąΒJ�!B]�L*aV�����K��ay�Ǘ\�ƾ��S�*���kxx��iu�M���9�q�w�UX�cv
�  :�F�n�p���B��mT�n�<0�&9���ycn��b���@��f��K��^3��Q�H*cpc4A��#ʢ;6�w;��v:��ֆ��적/s�Q��H�/���yu��b�J�ޏ����a�|hTEu��Ϋ��vJ�iZpO�#���,n�Y�S�8o���<+�6=]Y=��>�J�p�"n�{�C��%�ҝ�He����Q��YBYU�wv��cxhg���J4�^��<�Pb�`�-�����)s�49��/�¡K��^4� ����W�ה�T3��j^�t�_;������E��A��㲬^N~�bj:��Aym�7�Fy���5�������w󭿵a���sK�"_Y鳜�x�+����9Y}l.O�:5V�3:�v� ��__�ؤ���~�)�I"9�{7Cn4�z�P�[י��=k�.�[�w��&澷���v�ѤW,�鵛'>�#]��ٸ:��^��c�2F��Xu
u!cۆ�<;o(���I[s�u<��ʄ�g9�2y�.<E�1��R�~������Q�W�{�	E��U����g!d��_�(h��r���)��Su���$��4�ڇ^�at;O;��}����LX�&�t��b0�*��[����O�H��F���_�/����z� 6!}E�0�S1��mzm�x�.s葡��4-q힡�F瘭��τ�8�P�H���� ;`����b�)|_�^t�3�ÏM���Ǫߏ��c�بO4|��i���z�OT���Ĭ��O�.r��b����7Jq9�@S��f�;��'�	��3�t9̈�sHB�6�������_��o�h�u�q̿l�)C��5HM���p��+RK����P�t�c�\�5�p���kq�����uP.�n�qX��l����)du��TER+̬H�"/*�5�h�t:�ۉ{��i)�z�6^��>�.j�v��yF�y�8+�w�i;k9�AjwΨnI'�W;8s��s�;MH��T�	I�Nr)�\Zx�/|��ꏖ�D���<��U܃�W�.�ߗ�11�ء����H�2KCݙ��6욕R��_hU�K��w�'��˳���H.�P6�hu6�
��D�5t��@�����r�ڈl��$t�eW��4����ZQ�.�U�����T�w95�"It���,x��&\���J�cS=Bظ�6�2��P���ʸRf[ݾ!�L��Ό��V�x���m�l�0[�4������!Q��u�`�fz-S�kݗ���$5	�5�P���>����Z����:�!�C*j7�-� ��<��f�\B����[�>&=�1�&g��Or�^�d|kD/T�O>!��
�=��'O�k�`�Z��:���ٵ��=%ݟY��O!�uP��|�ꇴc��ʰpu��:��S��J{��Nz�m$nL�.��x��5�$CAE�V�]��+�>�̇�ƛ��j}�݉�4��<�&�i�3z{M�P�j�2܌I�j�Y�x����vaS��p��8�ed���H�\uᇃ]|��u3Yu^]ɫ�T�F�`���g�e:�z�:��I�kV�������Y;��E�ڒ켇1}AlZۓ�V�R�:<:>j�L�X��^�*uД��1]n,ޭ�qX3K2��B�SZ�H7����hcb��l��߮�C��07I뮜�3v�:�nc��΄RU��ygbAD3\���O �mr�׫�S�ڍ�����[*��mX�ٛ�)��ܸ��ݗ��R=��Zp,1Nj�jBT5;�7J��V�p<MX��ʹ��q*W�X�'em�o���V�O�o��G�zG�Ý֋�p�љ8e'H��Ɔ)o*�X��$�C_Q�+W�}�r����/9����Y�V;Ņ>��<��nf���/4��Ԏ,aw;���$�zƩa���dz��ԑ������ݍ�߄����D��X>�0m�>d�
܊m�J�	D|���ˋ�]c���b��QU��)$�I$�I$�I$�I$�I$�I$�$�'v�����#�<�P��r��P��YA�w�('r�{0�F��	z��P^g[8�>������ޥQb@I���Kھ\y�`�>��n�<4HS�3R
�j��j���:O�]le�ħ(�P���;��">������W�:��4|+�Z���w�w�
F�$�;�N���)��t����Ϫ��Mt��0��92�w��RS�ܭ̻��BM6W/��E	u�M�N��0��w��)�VKJ�f�4����#�}��v��/^y^]n�������s�����ޱE�Q���#\7G'W��G�T�C�z@�݇I���=�b6G�.͓�iH��U���J¾�S#��Ȣ���/���xi^�P�dX"[����k��e�w���D�m�կr��;u|t�3���5Hmƺ�Ӹ�w�_3�V�h��j�.�%�e�]WY�dM%��P�O��;vE1�udc
�<B�����~����F�@�e��[Sz�����.�N�W�o>���s3]
�=����l�BH��$�)�P��O��sfE4feTPdf`���9Kde�I�YI��KF�іYef�Pf�fX�4u�d�S�T�Y�cUj֛2����%�*�dUkZ�j�B*�0�+XaT�-�rOp�fqck(%���2�h���2�Y�UF�dUUDq$QV��,ՌWq��b�� �,Ĉ|��5�TLFq�4Fw�Յ5Yd�Q�a�0+X�іF13U�j��(��ac��dֳ,� ��\��0�;F_q�̾�5�Q�܏s�O�7�TŹ8.=Ϻ>Yf�Y�Wȓ�٤�j����u;i�o���X#���C�^d�����-p�=s��O�3�M:
�^���:=�	Ŏ������}�F��D�ΣC�2�y7���ۂ�M��Hn���2.|K���oKq�T�aF��+i��q2�1ZG�%ES�����g�B;>����P�����N�����l���q����� �E@EMx`c���5�yWC��Ӯ�9��4�b�u��15̫$j�������gcC��8�L��h|zƱ���R���漼�$����Gh��9Ib�lq�u���/�PJ�q�Q��[8���+�˃z� �����֨�$��G��42���eԡ��+��D#��������|{����4���	֎-��Z}��t8LV�^ʝA7x��jByZ�h�7C�%�\Q)�C�z�TplDu�j���U�	��[��U��Ŷ*5!5�Z'gAt�m^,��hV������;�[�/��xo���g�*x�+�)Ē��;)9���Z����ce^M���ޮ'V���v����8�鯯?>�-ܒw�H?�E&�J��G��>��s���U�3X�X�3�y9��rH���l�1�4�[I�t������F��1�$.N��7��R����&r�g<���D"��\2Lm�� ��Q��S`��sw��_��q';��VA��s�	�P�nnf8E|������U��9����G)3�u0�HmR�{9;B�!D�H���T�˯�DO`���3��]���!�:;TޡCc�����fo]�'��9[^<"u^�V��⯏��C������������m�^&P>�a��{nN#�O��*X<�h��
c-�p��g�w5����'(��;�y�)��YA �&�b����ߔ9Յq��8�rzw6���	�U<-ӼB�����&F�S��3���,�N_(xT��%t�PV����c� $C�����d���,	2��J�\Q�`a����ˤ˲n��[�:�ݮwxsM����5���K9'M���L�zJN�>Gz5L��Ǔ�Q����_W)���r�k���5уG>wu��ad:* 8O5���=�c�:�x�9�H��kvL�w,��K�s1A#}�N��S3Q!�<|r�oL�7XN>^r�X����^��U�*��������䯹7^�n��X,��C��2��DI��.*���,=�"zP�wM��c�_zf�f	��y��,G��똶uU޽C��(?�B�"��X��}n�n��N�\cۆ3-���5�{�S._�/���̅�_!��5�u
d���X��F��ǳ���ݞ����0M�Ef>x �z8#�T�9�ta/Ɗ���^^)Uu�=��C��ݻ�&��x3(:tǲN^@˜ лΐ�׻��̧x��g5U�!�g�Bsڡ`�!���������,��1��Ĩ�&rwo
j��.{syeQ�m	jD���J
��w�,�ε��q/%�%n�r���5�����H�:)8�W���i��w%��E�՘����6�,U��Z0��Wm����W����SkdD,�V�N�M�5�m��k�8��.�to8��u��oZ��j�����Wӧ3Am��8}7��L=�w$g�Q�T�fF�
�+��0��ɥ��'Q� ��Wi����X�	6e���.�HR�-X\��(~�竃�'b���n�{���qz1�lf��t�z4Ci���6x��~��L�;rg��i�P��a��m�bu���4��GI'�h�\"��:®����uwx�+C�CB�O�1��(���N�M*:LZC�J�zA�>���|�k���x�W�	U4�[Bn�/�ۮ��Z&���k�����z�Շ�p�.�8D5������%239ލ�О.��J��	'��8>�_5��긇�!��T� N�+�Ij7��.�+�P���ۓ�,�S]��t�����+�Ҟ���*1��孡�i	tS]��P!b�Pdʆl�������j5��q{�B��Ү�Ǹ�����Je$�,;A
�ѷ�R����]��B�E�u�l9���TuW5R>fM7·_r�����E��5XC,BC
�ò�b�P�D��w�&�gb�y�.O�a��Zz�d�p]��љ�Z�c��&!}*�ڇRu�哽Zn,8hb����:�;C�n�6��׽��)�@��\��!�Uq~�Kg=
`�}6�瞱��CK�V�J�I����L'���ה�/WD��|F��Ϧ1c���\���6,���,Uw~8&� 4=�U�%Z����W1������r-�+���V��C�QN �q�_��Ե����V>35f�Ǖ�=����j
�>�&l�P����]�o�Dk�| tMA��4<c9g�o>��弶���J�~2�^���>TU�d�B���и�S�q2As0�]t�r
I���!��$6��kOo�v(z�3�����3d�̹��ֶ�[�}�l�9����눊��أ4a�Xv�WtO,s9���2�HI��*>2�W���dY|Ĥ!�S#4.<���>�K�Ө�c��E�1ֈk3RX��� �k���d6�o��ˡ,���I����;"��|���:��vl������ᣩD�j��+k�z6��ô�����|�<ǹ�!���	U�>T��� ���lCN�?z����"�G�0[0�d�<�}�ǎ� ~�rG<#�F������m�P������0���ǵ��J����9�ݮ��!�u#g�L�Zx�{[s,����㛌����)4E�<��P��(�|"3�꣛��Z��y��y2l:y���q{V.6t skBs��u$&.1;}:�q����;=�9��/;y�Sk�E����3�Bc�X���7�kEv���m,��y[�v�V�{�Sa�iL����\1h��(k��є�:sn%��7��,�
テ��[�v��[�����Ʊ!���<bT}�VJXz�y����M�
py����W���"�}o��b"gǗ#��_:��9/í���Ag	p �����b�.���1�WK'n� �T�5�[X�`6�&wnz�=݄	t�cC�]j[&@��ζ��N��H�Ny����6q�����(��|�]�k�(��g9�Vu��L9ڝSf�A�����ah:U��|�i��t�ݿ�"v��3��o��F[b��ُ ?j�jS#�A�8�WW�2��<Z�R]���x����g�����nf��ظ�<�^�V_d��A�@����i��G?>��!��6�/_�1��q�󆇣��i�c�K��<��ݽJ>1�ö�Va�-|��ZU5�΅P�*�X�j�u��NGUsoP��©�parwu��児�
��y��k�S�L����*��_�\� u<�1.>��ICƌ�p����Hg�eg��D��joG�s����5��b�a�Cab��#�wPX#��+�^XZ��`�MA����Zaٱ��0��hl����ǅ��Ww>�3���X}���A�_����\X"��X���=#�D!|�`��d�L�Xz�Gq�o��'#\�1�-?TZ'����
��codm�i��
���f/�l�|y��r���꺇F���וӛ4�N��Q���D�މ&F��h�!����c�(�옘�0`dB��K�	d��p��e��)�v��H�Ğ-c͏�Rձ��Go��_ME��N�J��h4�_�\fJ�>����^����5K��������Q��@�u������L��Qufv�n��V�'C ���6�Q�5J� )� ٚ�2��qхgc'J�9�A�[�9-̌S,���w�:�|�|�By�.������s=�e:�����KqDT9�RD��S��������|r��XV�6��bM�7%L��{3���2�c6ߚ��-X\��(@�:�7��GQ�4�s��DZ�0��и�DU@�^����������3ؤhI\�D1��듐r��<�ɘ%Q�Z\+C�EDgU����w�SW�x|w#����L��:+X�~O.�n�k��u��4����	7�(0���b���l<�H�Mhj��	{U�"t�ÀB��]�c>{7�N���˝C7��d��'P�i��`�M�4�{��N����~��ANei�I_vǫ�:�8䚈�F��;o�ټ�N�-Zx�])B��E|Mf�m�e�L�3ӡ}T�U2��^��j�m.=�͍�^��{��n	2�_ޞ��wִ5��w¬V��vn�
�A޸�{���5@s�/=&���^�w4G�K��l�:xC�d���J�*z�h#��\{]<ԽP��>:C�z��p�P��{T:�Ds�/&��ȿ?%��}3�}�Ճ�-�,IT.�\u'Z��^�� �O���[��[-�w5���+�����!c�F�AUqqΖ�)����:��_g�\��i,�J�x�QF�^s����%~|C�a\u'�	��K8�m���͝�͕*�vg�����1��2�įT=����Іi�7ӓp�;tä�HOa�
1�#�!����ԑ[�C����`����p��;-�c��b����P�8})���Gh�|h$<z�ZЅn���L����C lf�9	UU��%f��|i����VtJ�-@�
�Y��4�u��ى��Ej�V�Q�c�˧�=ÑL�e=����v��,�_���3:vlo3���\}�܅~R�n'�����L�O8n�u��8{waq(���<j��8ן	�7#�v �����OC׎��7҇�kd���Y[p�ۨ��c\ܞi7}�q'�zڠ:� ����D<���(�?�Z+
E��~]��ܺ��i$=�y!���9k��hW�L�q����j��{���n����0��Tud��֕xu;���ƪ�Q=�d�{�xj���q�"l���V;�>��ц�6�����42��/u(D�O=��w��<�r��	s�O:�5�q�u#fKl�Ze�d�;X��|UY��̒`�WP���0Z�$^k�lyK".z�tln4y���P�_����X�-bP�3�Ν�fw��ly��=�	��vў;-_m�]Z��k�����Z���3�1H������c�o������g���?��b��T�47eV�a)xզ�!�郆�cT6�&���Ps����Η�X�Z_;�����r�S|v�{#uuzz���gt��j���L=�$��˕Y�p��2ۗ\w�9�s���y��\��z��k5����_+C��J�NL�:/j�c}�`�u���w]�|i4���X1C|�����fʫ���s�ںܭ����h�����=IZܑ�2�����	�J5�\��vs89Ԩ�7A���4�����jr]����2�
ϠF�bw��ϙ�cu�Ӯ���)_M{����V��n�.�E�|����;�9���%�;�I�
��a�]E�+fqku����@{*N9+z��������µo��?h;��+|��l�����lAj� T��lbS��YA��q�ʧWW>�V{m��o���a��d3ck��@Rʾ4��x�s;'�X��̽?
�M�J喏%Ԩ�t��;�i�e�,�D r��J�G���4S��]����6���\����F:b��L1��S±� 5:7�*�ՠ{��tڳ���$�9ԝ���r��#�1�Z҆�ط�Ҫ��$�I$�I$�I$�I$�I$�I$�I$�I,��'@SK�&��*p�Ff.SP'��ݶ&<EiM�h�a�+���8�}үe�|�m���aYa]ɠl;2Z]��̊���9���Ļz�J��8Br�)��g]�!�Gg�Э�aooû�^�C�BJ$�D��v�����k��t�9fYl�yvXS!\�kC[&�E�'κ�x1�B8�:��٧(������㜾ُ����T�.NV�B�	)�׫B-w�f�o6��f��K����s����sa8a��lٍ^�H����Ŭ�m`�_����z��tc#�wqz�V�F���}y�.��9]��u�A_sދx�ڷ��͡Fgo[#]����_Q�Xt�Pw"'�%���^݊��������.���
�mp�3rլ�^��j|x��V�.�V�Ӈ�1=*��U	�Z;]��N2�x���X���7%3�zJē�+��f�����^���.�l�%���=��LK�p�n-J]�K��Y$�$#*�(��P�3��b��kG��m���}�}��w�e4Mؙgq�AAQ�#&##Z�f9�DED�c�����8L1UT56T�ISa�Rwd�UU�,���1��P�4F`ђAU=fQ��`�ř���Y�ё�PĦ��A�bPAI\ڌ�b��2���QES5	��M��H��=�2Ց��Rj2JJJ�(�)�0�YE4D��C̨ �B�e���Y�eT9eAT�k�(��Pe4CA@SDQPUP�E)IMQ:�Ց�U=ˍ�ʦ�0�*��&��"�Z*�*��"�1��b1	uo}ӣg�����R�b��2e�ⷓ�2�P<�Ż1��^H%F��˫
J����MCɵګ������73U
��G�6�G����+�f�	�!�|�8�Af,>F�X*T;��xw/�5�!�Ӄ��%�EA�T[D����%ֆL\C�^��'�Eļ�2z�pC�R�7'wnSL�n�I�����;�r�|S>�R�K�oC$�L�kV��^I=��9�R8<�!��U��S徊��k�=��b�(9��%��g�]��os��f}�R�i/L=2��=B�"��O�E���~9�]A�b��8�;͎�k�ٹA�a�b�vS�q�~p׼�x���4AjW7.���o��Af��c��g��t�����T����f���Z�N{���Ce��/�h�M�6Q��q<'�B�(�+-ol+�;�-�U�uq�'��K��s1A#Dmê�2k$P���Z�ʘ���T�X~�n�-qX�;rv����9���D��a�Kɫk�y���gP���6%���)��#�tZgz;@��,Vh�s�]D��S���k�Gb����S��e.�I}i���L��w�Ln^�X�1�\i'��43��J�����2»�j�E:��;%H�U��&��=I��՞�=+ˏ��˩
��{!5$�}ݙ;6ý�[��~T=\~��͚yX�q���|o"�F-�#��m�Uh���}��P��Uq3��hE]R�*��kԮ7:T���ոt6`����Igbm{�׬�hL�����Sy�u�^�w�=�n���:��轭���+�q�R��,�xt������U��Vzzj�1	���9HE�$������o��9N�bCM j�]��Jϊ0.ze��6��H�!�����#s�P�.z?t!=2%�ȶI��>]kƒ'Jb����Y��^Z'
���[X8z�|.�0�8�c�z����ֻ2!�� X}QQ�n��>�8��Z@zK5��IMw7x��HtN��s��3v�9�o"�*��/��^�����%��2��R�.w�!��39k74⢪�#V.���N���u��5�;�|����G��6����E���9�]�Gjs����u��,+���U�+�r�_:�G��b��A�WM�5��٬���������8���ѷB�L�69bB�UI��B	?V�Ld�	��B4^pbR�b�z4G��f��,\_�˩��ָ��m�U�d ��uL1Hu��"<PਚJX(d����xj�ݙ�;n�Ȳ�B���>~��Re����>D4Z�眞A�t�b��8vF��$֎W�*��nМ�"}�|)3Zx�k���g:��C[}���(Ϸ2�jrS�"�0�����F��%�rc���\C�`��o��kQg�����r�_��P�P��5��,�ҫPqY5<KIu�X���]y����`˪p�[dlU�:��哽�mx��R4��=g�Ӳ�Vx-Rz7\"��W�a<p����Zz��^��X�[����A=,%�<��5x��K(SKq�3dǜ�Z�ÀThR�nV���G_3R�j�J����nX9ʝ����(�i��ۺ��x
y#&&T��`N�2zc7��e�H��ˎJ��zu4�oQ���t��;b��u� @���T��q��Ϣ��=��-�]u��k�~�����'�3�O���PT<�3�U���g�O[}B���j��c��*�L�˗�K��ǌ^���5�C��8����u$G�wq�k�[���.8z��!�Ԃ#��!�T7��ԏ��c�G�Ç��
�C��1��9��%�}��NL񕳱�y>��u,�oK���u9~�]�O^o.[a�'ʼ�OZdԼY��q�R\��*����b��{�缘����C@�,X<�K���:Z�2��!���Az�@�I�7��� L1{Hg��J�kǝUq�(x�ׯ���2/+�-c�ۜO�����t\�����Q�.���ۯV��:��O�ϒ{Y�y�;Ǯ��e�K⏋�r�H�TY��6����he�fO+�uV��[|��:Z{ci�5Y����n��J���.r�a�Gkb��3b�$�xݼD��1���^\Qn.u>��{����Bf,p�������,���җjP�����f�jN���*����^"��!���' �%@t�1N�l��L�HQ����z17fH�7�=ݶ��딃�c�[B������-��B0����(1}绷�����1+X��,0n<��QwN�������)Yfz	��ؙ���W��u��8S-hU�0=��G���e����:�o�B��Ls�>53{�*�f�N�B�*� ��\��񱻑o8n�Μ��=5��p�FL�bݰ{mv��~U�73"��Tuw1��z����Wqs"�pwI��A���2
�	��vD)yhH��=.Ei�nN��#ꦾ��>`��I3��8��8�TEyh��+0�w[Rn̤|㧍���@e#���G���_-���w�6��F,;[��.������z����2�^��&P>����)����(5�>@Me7�m���5�����ެ��\E������+�I�p{�P�$Q,X������3���א;ǳ�ٺb0�������۩g�׈�t��}���i8D论]zI�VI�%|�
�&��Q�]KC��적�bH��0�0)Đ�Φ/�{:ֺv*�u���,]4xh@��Җ��~[��7T���Ӻ�E�Y7zS�9f��L+�-�{A��KG��ɺ��!�8T��ouGE34�I>f��k �oqĸ߹����>2����0ήx�m.����EӇ�7�U�X�W�^��}�CAȴ�[�ח:��@�N�	%vL!bnQ�89u�̨Bb�:}I��g����������;`�,�Ӄ��]']�k:�/�|�U��̝����IpW�r�����C��E�=�c!:��ώ�#���b����|������M��^s^Dm���\Gj�#�.^f����}�¯_<]{��*�YL�%��}R`�6xf{�=]3�V�yi�A����
�g�q��J��[ug5iz9{dmx�f�Xa������l�5�{Gń���ۻ�<_�u�C�X�_���h}Xv�u�*Ct���I�ԩ�k��;�񟛣y#N:TT@�������\��)W�47Y��s���[�w}��I����\����#f������@�*�1HN;0n8ۇ��g8�4�q�t���d�X�aG��*Pڷ�#��<{�z���:{����oNś�-���KP�N	L]m1�ܥ��zs�"���_�GMA]ӌ�c�!�qK#!L/�Gr쿫��$ٖ��u�B��-v��wB��_aOP� ��=Kz�ȹa�vF)��g�"0��B���mr��)�d]�eo���'��C\1���Lgދ8o&�	�yc�ˑy+~}�H���ƅX��쏃C���3u��u&�	p��N�2��$h�<�����0�
qc�����(��d��Vd��=k{؞糄�=�mץi���Qa�q)U�6�
��	����b�Z�d����!�����F�x���SZo,Uq���UH�3	ݵ|�:��&m�Q��Ҟ�$�Z��s,Z�(!{se	��5,��qV��/��m�b�[��9ԀY�|��R4V__q�@�}�inغ�;�gjH�Z�ͽ����[���d�Β�>��>�^w-̦�DTC측=�r�̍w�Lx�Җ.�xl\�^{ٛǵevv[/k�V�T3���Z#���(TGl������,_��+*�E�h�4�B�qԫTE׹���g��~vwK�s�����j<*�0�=;�"Ϗx�ryKSK��G��U�1�OA�o�/�z�l�E5T�F��^r!y��V=HEDP�i�Z����P��T�����c�l��y�*,ә�4���8��yϨ�b�'�p���\)���	�C��đ�ܪ_<�^؇�S���m�ycoUj.	�ˮG��T��Pѳl�a�S��+F�+���I��)�����u�\�B����D�꣓q��6�s�ҥ���VP��!��V��2��X����t}}�0J������ccC�V"��`�.�æJ�~:]��|�l%Tz��n��.l:*��m���%wI�ΥZ1�]�ǻ�Ş�MF��e�H��;��-dWs�V��L]gtO+�����i��*;�3�@��Q:�q���Z�O��_�#C���{�u��0{{{�G���T���i�д��0y6�L>%Y���	�f��n?nM�!��C˗�4�uJ9e����u��>
Ϥ|#s�9ɋ`����u�0HC\JR���ᤑ]�V�Z/2߃C������WP���}|�,ladp�P�ꑁ���b�+$�t����Lo6r���+N\l�%�m����\���.e���#;�vՒ�Wuv=�8U&G�B����0p�QA�^_5��i�aW��Ϻ#7��z�ZϪu�w��W�j#���G
e;�`��E��B�z��D��X�`�n���f��1�S��X͞���!�t� ����Y.�[Q�

\+�n0�s5=~���f>�����8MABVc-¼s�J�~G4�b�{L&/0�Y�0)]u9FVҩWC�v貙�D�np0�2q�K����#,ҕ�;}���{�ԽK�U�sD;X�1��Q+;E����N�� ��m�}#��KR�Ɯ�k�~7���ݞY_�É����W/����|+���������=*���d�1ݞ1y�O�t�DC���L�|g��.��4�߳�2��Ϳ'��w��>1"p9�e��y��*1Q{Z<k6����P�:�V3������bH]C���8���tv�������A��\(<�r��G�>:�w��2�h�.�F�,�	H�8h�K�2�t�;�*P�R�v��i�H.<<����S+��w��_���(="]Et��y���\�*�7k��zhD�=�:��犑��8m����\�,G��n��:�����s���F�����J4eS�xz�Dt5����wL��(����*���V���@��O%��0�bݾ�v����	�dp�7+��>M������5b�c��=�w�ү(lP�Z����GhL�c;�*ةI=C�(�z���-W���Ʋ����$n�ll����l㹨 ya��r��f��`5������B�Ɲ�_6�k�h�q�)f��Y}ZT�x�K']_r�i���AH���v��i���}��ΜX�/��w��l���7@��yt煩*�北*��p�-�Ks+�::��kK�g�q���I�� J����_���w^�<�,��㮦I���Z;�.��5�]����s��L-�{��[���9+��)��	8΢�.i�Z�@UׯtIK����D�MM�n���m9�n���3q]�E<�sy+z��WWt,�k��r��L�;�ĭ�{���&1&hPR �S��j
��e��Y�{�S�A6�K9ڎE%�:^l0љ��%^�]�/���6l�R�Ȗeo2x������
�N�8#��Hq���u.n���Ã���R���\f����	[I7,,�`�����2��T��٢�&P��[j�u*�>�=]4D��K��5<[�W#09y��U����*�
�Q�ϐ�R���'�#R���2���l$�o��w�(��vS]�"$1��,k.Z�:믡��=[p����RI$�I$�I$�I$�I$�I$�I$�I$��ޘ$���:y���]�QK�(pJۣհK�х�Qw
�U��4t�)��i�-삮�$]�Щ�<��C2Bz��,���JB��;N�{$	J��(ݚg\N�^{��m�e�lƦ殗t;���Y|�&o�z�؜���S��MZ�"��jq��QB:Q�q�
�Ы���{x�+�r�k2k㸟]�#2R�*rgl�bmu�)5�C����@���N��^�lU�n�mk���V����vbBH,[k���spoJ5�OM��V�U�]��}��{QkH�D�.1iI��֡��h������i�Ir�}.å���>y��ϱlԟ���B����eg�h��fb�U��v��u�y;�c+T��`��d���%+~�xa�#đ�[+]����s-f���⌂��Wfue�bo[�8��#Nܷֹ�ނ�%�z�b��gS�HE�+��L����;�	m��L
������N=�+�W|i9�`�:����!�d���J�8XS�EqIR�"f �@KSEDQQPPS150�RV�(� /pʀ����()����ʋXQDQDMEPU�ED�$BRATUTA�T��DLE4�5AVf1k0� ������i*!�i���l�%�<�j�����XRT\I��RSMEI@PU0S�M%��&REDLIE44LSL���D4EIUM%M,�IU4�$UIE�(��$("k�\��""j��("�����Jh�f&��"B�ZH��.r����`h"i��bX�"�bJ��
J��
F`��i)�f
���i
F�*��`��())3������ӳ�j��nd�z�GQ賂$j]+4Lf%�5����]ep:&fmH)"ټ%%2��+�i��=���e��V�K��=o�X�R�立[Zh��x�(D���:�)C
A=Q���r/�1�N�vs���EP�W3�������2��������v���0��:�^Qs6.���^{������8�����p�]��d�yVK���1P{���
��!ڸ�*�mՑY���X�ے���]�\�	a�.��*֞�#q���|��_-�C���{�_
��X��,::����~�Nd^��/%e�C}����jj&B;q�'��܇r��$�6���ck��-6�Ӝ�|ulY�>�mKZN0tq�6��d)�����u�̈b: ����1|뷘�#����)3�,�.'����ǎ�!A���3y���t} i�4+O����v C>�}]�tO�𬆸*�c;{n�~�|.��5&u{�{�6�G��S��`%�v����.m��W{[�nPH�J�&hh�P�[������np��B��;K5H4@�w4��㓡�r�{�iM�Lǟ���MG�^o[Y˷`��j��x�n�ܩ��UX�Ql\T\��ædz��8k�&en���cn3�9���I��F�YU ��DE]Rti	y~*�6�D�x�K=�������E���:�~㙑��멘�rn�x��R�\l
��S2& 9{ݱC��xp�١�+���-�ٍ�B9*��܈��"�0@<�c5ܾ�܋15�YzQ��`2�D�u"��b{N�*�F�ω�/j�C��ʺ��m?L�>xg�;hW,0�Q+�ʆb����yh���|N��wy��ޖr����YT+谍-�.J�vJ�@�z�#����M��=���Yb�SfPǋ�s«O��at����{L��ǏD�-����Ga�o[js�,(��R�����^R!��%cψuʦ�$l���������T�eC��o��鏂�y��E`�'Ҫ;�6,әc�h�Qp�����p�]I�H�VvCIXv;����cc��B�2xW��Zum;�^ؽ��r�8�ccu�l9���������G��]�t�>&uxM��]��ap]Ֆ�vFnp��\1.�Z��H�~����K�:���4øux��zhw���:1�#�!����u)���B[]�ֱ&�WZ�����m��9c��7���\��F�R7iL�)���y=k�Tx�,��@��^�w��|̾�ܫz�{�V����-ʊIʲ���֢t�H!��=-2j^+GG��]4w���sH�=Ʈ��zK��{���=l�N��|�v�|eST+X ������n�h�m�9��Oڹ�t��L�Nm�M?����k�6�� � ⬾�O�3.���+��Y�Q����i�}_q��b�Z�T��yp�3�B_�F3x��mK���a&�C(���{��訳���+_kų5F�2�h��YTR�X�\����*_jb�֎�)�H[�ͩ��U]��2u��<�R璆�ה��"����|��"�H�+7h��ӿE0��.��Bn���ƣ�ڼT���`F�KY��8kсMv��rw�۝Q鱻[�q��9Ŝ�=O�&�w�,7���+aA�.����3lb۷��&3�K������nLX����ڐDEd亇u�qX�`�(;���כ�����/���T�Ϻ?j�j��o�?)�N�X#��{ǖ�5�v�Ѽ�!(�v4�!ͧ�تb}���j�V�ʗ0XC�pV���ߞI��n��T2��\x�B��P�f��wWŢ���t�&��=;��B����)���Rg=�Q}hdL_�
�v'�Eļ�;(���#�O%��!�bG��]5���Ab�6˫;���:z��
�}��%V�u�>�.g0�H�0T9���r���4��ُڞnA�{dbƊ}PD�C��s~\(>ʦhyD�	>3 a閴����K�0��5L\co�!����QW"9f�WN�F�JM�0�T���<3�C�cHo���]���w�`��}a8X^@�Qh㩎�����-����m�4�!�+�̺�%\�C)�����/1iT����h���9ح�u�tb��4�6t:��̛�Y��5�>��{,��>����PE3�mK\&d�5+����1�_� ŪOG�jY��+�0���T<*_�-t8J��U�r/��t���8�C�;�1�u�;\�b'��K��s1Am�pv#wWϱ��Y�:۠�Pdq���YC��P�i'�-�w��|�ݐ�-������{��}ѺułϝjB<���p4�����e�{c�y_�D8��w����5�����qZ熼�I�WLb�ΐ��!�#*H�КO����N�c���C�hԶP�h���}���p�Us1����.	���|
�K��)�چ�V/Ya�.1+b6�`��օ�7LP4�V��Q��'��ճR�3��������`��1���-
ܮޑ�WYgISb���oΘ�,E�����/h���� �A�^�l��Tlh��l��+��Z�Iv��y�mԱ��O�uc�z9uaFU�J�#w,�I���[Cf��	������Ǟ�;��z���7�	o��z6���
��ȮW�a�{j^�zi���]��Ye!]2�#vg��EV�K�_(6���.�q'B�Y5	�!⹓R�%�9��醮�����,�>j���W5�Z��:7�LiF4	���|y	�9��>�*����
kns�鬎[Y�v�=�hʥ\��9� �ׯl;ۉ3�wI�7U⋁�nt�%�c6��C�D�;����&�eaz��Xwr�|a=n�:����Lr����r*#����lR��5��d9�,�V7J13���L��sJ4�8UR^S�::���]�+b*�	�YV!LNeT���Daw\�mtu�O^_��):�[�U��sI���A	�}}��������W��gf#Y�����ԥ*��N%��n�q�Ŋ+���Π��鬋ͯ":�+�U�^����8JȬS�O���o�^in�;ol��͌��ׯn!��{/�{=28 ������F)ԇ<��knS�z��펕��\������ѭ��Jkv�/�ssBM��Ϣ^��Q�b��3[���EYoh�V��q��K8�s~����T��z{���[��%8���%�ao8g��{������yPb��ַ�X6M!I�V'b�L$�h���)��KQF�.w����ԡ�n�;q�e���
N�/U�F�hyؙ����=S)�Qu�}��Rmɧrب��	�j�޸(:z4��eVӋ���\����Ju�P��y��Y���L�\�F��ܗ���ښ��ځ���lu��zX��g�X�X�YR���6P��6��6���<P[�����y����p�T�ތ{e"��K�b�4'l;y���0*3��ߵyS���KP(P^��Hy���-!�Ǆ�r�����,/�@Џ�4ӍVlb�(�JA�᎗8����vۮ�h���f�V�ݡݩ 8�[�E�v�,�H�X�s�AV���>�
j��B�z�)G7�?=5�j�8J��
��]u'][ь�v`^�&ث����ŬL$���[�9.oN<k�e��+/����~����,�E�%�1m��|��[��w��6�ܸk'逍�z�u�Q�kJ�b���T�P����z���Ǘ�V��)�4���֦g��e�^0e_i������͗p`ς�Q�j{y������ܬ�.�)ap�e�5h���m�{�:j�j�^7 vu�Nؗ���Fs�w�˄�Y�nQ�EH��h���+{�r�N�LSb��юy����������T����(N��1�w�r�.
1��a5���8�4=�+xv�--�lZ��� �n�X�*���u��{�"���H�B�x�$#�r�wo$Gs�ku{���ƙ:�w\q8&�C�ͷ�VimA*J�� Qޅt��gwi�;��O�9�N�Z�E_Ń^��X����;n��8���?�vq��&T}��e�B���$��m1���-G^��Ok�q:{R�\Œ�T�ڝf���qUrj:4����a�dh	9�zp"zO)���O�l�s��읦�� �Q�^�ע���M��|����s�
�WqJiN[�)+9,^��yLd{�%l��X�˾U��1NI�	@}WS�vY�G+8�w
�Z.G3���Ŗ��c,FFFF�a�[Q�[Ci���m��1(��M5Q�F!-�3��^��l�з�9ZC9GV�鳃:+ ��oC·�R�����a��U�V���*}~���9�u+S�#I�r����C�]�h��ݐ�.q��v2��r�;޾��BVx�1�gm��^����7�%����2F�b�\�ɕӡez���}����=)�=J�u8x&]oO,�Pr��9-��ﵕɩ�ߗMe+z�\j�uz��[�[���LN�^'x�^\g�.g��5��mΣoSUU�aE=�ޖ\�����Sݿt\��=�svR��\��λ����H,��X�=��X���2;�VX����F�e�Gv��,�p�\��M'�8t<FeT��QhSs�Ek$��#������ �[��(�:��]=m�1L�Ѽi�tJ�w7Cg]�yT^���(>[r�-��3��J����s	׬�W�lu�/}���W�WR���E�2�cv�7��Ɋ(�]V¾��!���3VpZg�7�r[q�>7�7U��8��.��6��b��
}��
>UU������5����h>U�|9��1g ��Α��^�"�Kg�O��w
ӝ�H�S�̈饚7�������kE�K�_R�F��_�/d7�l�8;2���H�ȭZl+ޥw\$�'sWx��H�rf�i��I{�g$xn^�����,U�Y*��uj^=x֞պْm:&���:�M�Oh���b.c���R"�b�b8$}����s*-:F�d�L�1��V�Ή�z�"%$���q��M�$���(���k��ۛ����8�q�s�2�vj�C�/��I 5��h�Z4'\Ω�L�ũЬ��w��ٕ.�N}e�$GRE�~dy�>H��/3���)̼��f��n���a#�R�j�V��<]������wǌz([���H���vҹ�x���+`!PLb��S7h��c���yaP�s{1��C�̮m=W����C����<��hA�Nn�:���ǵ4(o��b�efRi�`o*�1<6^�bT5�U��9Z�h��J�۝,k{(lR.�,1rn6��
Zg�'3'<ͻ0��I��R�n)��ɦz���w��][�7�v��corM�iɴkF��ќ^鸚aR��5����I$�I$�I$�I$�I$�I$�I$�K6;��0�ѾЮ/q%;�u�q*�F_3+z�<��Y��]ol̽��{8���v��9;
��L���x)�ys�Н2T<[m���5٭�M�)���S:�7�HozF�k�	-�����3�,�z�nV��]-M�++PJۛ�-t,�;�T-����۵�P����CqՉW�3�ܝ�)�%ky������4sԡ�`R�f3�L�z�b�n�b���9�*'PuZ}�.ٜܲX{>��.��N�8*�<=ư*�r��o8]������9ͺ�����뗸H�R^�N�yr˛��V��w��A�&�f�y��0ht�K8�a�-��Y�m��2��k�z��������{[�B�?�,f����ٚy���E���jxs�Pd(�O��7*`u
��/�ds-۷�i�}����ɻ��л�˼��+u	"(�E}����#�Z5WM�n9ϗcoc����yi��-h��}C����>h��y�&����X�1����,�}'-��|;/��={;(ٮ
AEr\RG�\W�g��H�����*(
B�(��HbV�)��i���a��h������CQIO�eIM�PPO�TE�Q4SABUMJ�+T�QAZ�	
�S�J&�(�J(
PU������$ �J�\������(bi&h�:��Y4P�C��2��!�(ihi�r
iY�����JV�C���PSTT��Q�q:�h��$���*����;�ɠ���"Z{��*�L����j�JJZ�JaP�@RD�@�-��;���� �땱pѝ�I�v��sT�z��H���s0��:��2�oT�n[6:�%�uj��
aef�트����/��,���`-����sˑD�H�T��ư_p�d���I!��[�S�����^Z|,�ޞ��y̩�vح���v��hu>ɨ/'�yg�����ٸ���	�n;(�Fcn3�ca<�}zV�wjSK�g=*��S��tVd@Z��j�oL��u�^��p��5 s����v��-���˾�b�V�_��zT��VK�h���2��}��U����O�Z�M���ng��|eZ�PR����2�o���KjPr�s�u���&�#+�]�k���aT_+(���IK��b��k�KjӁ��*W�dTc9xM[�p_\y��rW�'�����"�;���)O�ӧ\\Z�Z�9�;)������'��\X��<�Y{Z.���;�vp�Ykfv��)���K�^��Ht�*oC��r2���gq.ز�t�{nʜ��:��k:4T�K�q�u�n��� ��]�:��7�g!}��N���C����+Z;rA���^
��}���YU|��#��)�D9��$�U<{�����q�온1��*��W�3�<�>~La;�ܘ��6	*rG�Qs��S�8Ae3w�l�齴��L幡����]{^ЕJ%W���J��H�r�0{$�ͳٸ�7�jS�]f�b
���Bּ��(wbK��f]�1[�WVY�ޑ�����^[��V0*�į�FsL\����N�[n�6Y��<��j�Ն:`3y+kY���Wj�)H$�Pz��-�$��0�}}FŢc6��u�I[���&N_��z������7��/N���h-UG ���B;M�i0�� ����)��}1J�e�@��I�c+����B��7K�#t��TR�J���TY=�2�,��+dG�ҫ.@)�_�˗:ʊi�`w.�u������\�O��-�;Z�?n�̩��U������W�:o6:�����y��m֧���r�4n9��M5��nQ�Y���
^������.���z�1� q�Ӿ����s�ˢ�K�G���`��"�5U]�5h�-gjV�"`��[������� �v��+��2�쳈��O�	k�:/yCu�]����[��*O1�^�q��1u�碲�cJ��<��Ƴq���qE�][�ۜ�8� {�o�Ld�Z-Is��������u+���M����X#�cs�������ɩ_�PZ����>�9�����e������՜�B�o`��Zv/�]y��j����q��ǒ߮�HflG�$h�WP���E�taT����i���=��խ�Cvwyq��y�c����:3N�K#�Ե�z�`��&���Msobc�Mm�	Y�[�\JJvv{x��3��h)�ۏ���n�Fh�h]�;2�����_Ir�o��o97(C�ʈ���7u���0r��[M<�Nl�饬�� �����l������;���z���R��X�Sy㮶���Eگ���,TZ��=��;{+�t�Ű��}��#���|���Qz��^�*�o���t�#a�e[��i�̶����Ez4N��0cJ�*�Z��.�Iv��s;��Sy���t�KQusp�fk��)�-���Tj^�����������V�tf|;�Qe�j&�n/n��U$�c�8-���}�yM����:��Or'�xq����%s��F�5*�U����������"�|�v���9ՙ�$�s�ͱbԣw֭�v�]�r����0;ȁ\\�y<Ķ���}L�R�d�b�w6���3˹.ul��N���5|��N�b��r��_w~FU��.�W�Lk�5P\wڝE�+�n��(2E�q�u��t�����c�ߢ`��z��uh/q�F�����������q�&(�ED�7+��U�kS��ޢ�ur�� ޱ��=;��C)��0�Z����(ne_�+|�g�`켅_	���{�}��"���?��t�9�l\�=U���Ȭp��a�9GL$��	��f�=�H�;����Rwm^eT[��&1(�i�����ʦ��A��W��vf�s��zj߬���[q1Ɋ+��뭉>�fUMf6�6��U�F/(=|g'w�;�Fv��[�#vj19�Z�D7��
�o�gL��Yb���&I�әdw��x��lR�]�龎��;�<�Q����-4���6:71X�W�W�%�G��������c�����C0��S���Z�����(�����uA}�*f٦�����D�Rˊ9�ݧ+T�g�?{���[����5�k:v�j5�R�t4��E��C�Hie��_*o&��E�h�ޑ�7V�w�7ŧ�i*�q��|����ri\�w�8L��rs���Յ�T���g/	�����p�9�ێ���{b����v�_�_X���崙�!�!�f�ݡ��ɻ���������;��VT�F��^�AtUk�쎁!����P�'�I��gvv,ʑw<4�0h��N��]�]�^{ z��\�`���pn���'�3KJ��;��i��$<�\���n=@ձ���k���R�j�܇}C��Ws����!`:��O��\c����+�����TBE^��)���+��$e���ڂ������X]d.�Rs�s��h伲wj�۠�H��7�]P��حms��Z�,������D�|뤬��a��ݽl��މ�a����2�]�O�r]�6^�f.��v�ր�"b1(Æƕ=���"�r�dmA9uq�u᎐��R�g|r��N��f?ůU�[�k4V�hd����F/t'Z�+(��g(�p�kE88���46�7�	�/F��1gBЪ��B�n�֌�]�+P8��+��O�u�;�Vro�����Y/j8��F�~i��J/��8ѿs{i��)��lV㬫�e���T��Z2�c{�������9�:o�ѪF��:n�B��/dQ�Ѡ�\�`�i��DV�"5.�xQ+�d������� �O١⸙�t�ܳ�n�7t�+�e�Nj.���޲����ʩ�)�SI>�l�k3Ս�ۯo7�t�A�\u��b�rv���B)}��5ܓQ.�l�\�tt.��xr�ft�7�/	���y�GMoB��yO7��!�4E���}՘%r{���H�8�n򏍺���y	�9\�S��WE�w�e:�ܚ�8[Pi͖F������<u���1�L�K���H���y�|j�J�Sf[��7nZC�D�:�}�epʌ/^Q�z�G�r�;�w�slOG/����!rqA��zq���x�c@6����N����"��cuM)���]�%׮�\f8w�����Vq( 6�V�h$3|�]����G7"��;�ow�qj,s�.:��F�K��q��:K��1{���Oi��6�#%Yt�eg�M]�n2�������ޡ7���ݸ+�V�d������y����'
Οs���E���9V���n��>+��+F=N�!h�+˼�S�;��n{�.o8VR��}&��$�/7ob���D��T�[���tE��E�}�5�ܕ���AOzh��G9�nfk���۲	�}��Ї+#���P�X�����rfWM��Vh��\��R�ǝ]�I%|�U��KX[�3����=+1EMO���sxR1��fԷr:�"ܰ��}m=�|��l�R�p�3!s�R�����7՛���X�Jq�����+��������]yy��Rlt������v>S��NؽN�gZ�<K(�������s	׬��~�f�Q{����^�9�tf��KMq���w���VB��ջ_kn�mT�X��/yl6�9kWG������a_�OxՐP��xT����1�b�4���:��oY
p��G�����tO���?3ʘ@��֝���W)�[
vGGV�s8
��@(�G��������{�;�;�t�0r�s�Uj���ǟ?S}V%��]ξ�]��Z���d��xrs!5�qн����}Yw���%���M3��8�0
�q�m���/�>��u#N��X�NW��U�t@�����<�w9��.�^���;�B��r�������lq�EDs��CC���o8�C�yy�)��N,�Ρ��ە�m�|�ެ����Bg{;D���7�ɻ��,�E[�P��U{q�;�MN�`n�D�@�8zE[or޿7����߰ς�Q�kk�]�bJ`�#)9%��ޣ�x�����}7����t�T��{9º�h���>�j4�������-�E�Yw�f�;�&��c�R�ldE�"���yhyɥ2.1�s�T��	�]��t�lQn|�Mͬ�S;fxC#*@GRױ���2®vl!е�O*��7,��^i��vzv����׌a���U���
�i���:��0+�^������G� >���*?^eMU���"��:��?⊂���	��*
���"z�ph�N�����]g��8?��G���*(@��G��*(��@��Z��5�f�9���I�u��~;���	���p?�ӗ��)����q�`�
���"���}�E�������?�&��A��6�Di�y9��������N��'���}�~=>��LѠ���w�o��(��}���~G�����X^�?`���`��Q�d?Z%&.�ܟ������`~����z��NL?���y��i?i���^C��������?�O����~���1�Ma���NO�?�8!;t��!�'"^��F��3�|p����J����G��~d�������#�W�!��&"��1��91���u�9�_��DG �(�o�}��yt`r��3A������g~gH~[����h�(��K��:���?���A���9L�M��ߏ��~��)?S�)�����������!�O� a�?�?�W����� ���Y���?��������?����?�GG��c�_���0;�/�g����u�?xK\�漃����<���~�/_�?w������ �(����y����?�?��r>!�h��p����0��8��TP#A�H�(�C�C��H�.O�@��?Q�8����p/��#Ô�S�9 �`�~ZE@z��:�) ��4�N���k� T^L^G�!O�~��y�����Iֲ�p�b?t&���BC�'�`s��㠯���yЪ
�������b��O�
������/�
����� C������}���?�?����~����)��?R�0o��h�3�A����~�2�����~�8����'�����`*
���|���0��L�����Ŀ���C�������!��z�l?���>�'���t~Bg������N���<b��p?���/� �?�������*|A������/�i;O��9�����t
������X='�;��-���$��������0F�?d�A�0�����Ñ8@���S��?L "�����t�04��B{���o��3�}���~`"*'�$T�����H{���~���[��|d9�_ۤ?�Z��OД�'�H���O�����{�rE8P�0���