BZh91AY&SY��#ps�ߔpyg����߰����  `�T  >�   4/5-h�   k}��|�               � ��
ǁ���2 �    ��{맣_F���o�η7;>�������[��o��#ŏ}���N�����z�ϻ=Z���[���]U���)���=Ƴ�s:κ�l|��˻�   �����m힛�㷞���^�G��n�Ub^�s׹{�Ӽ{�����e�7�o������ލ{cӮ]���\�x��s���n�s��׻t�4;t��  ����my��9����v��v�[�ڽ����u�{�Q�H�}Ͻ��>��믽�[�6�m�;�l�ݛ�;��w�  =�/�9�;W7��yǯp<�s�u�{��Sn��=v�����B=��{>��m��ٺ��y���������=w�z�0� >  �@k�7��]4۽�=�{�k����Q���p���]�� �g�͟w.�;׽���{t�{���/��{7c�>S쪂(�UJ(�U
 P        ` ��  *��h~�T�FA�&C#����J�F�#	�i�#i� M��A
�!�&a1h0LLLA&�)U ѣ&�4 M LF�D�!�514MS�J~Se='�~��~���G�٪~� �L�J�P10	�L���4�L�����Td��X�%��ī�ܥ�C�Ok����Oz ��%��|r� ��� A��%[������-��͍B\xXu$��@G
��1j襡�����t�p����N�*(-� ��P ���u��z�o�=>�_�/u���_2h�˂sBw��'4[�sŬ�>=\&��[T��ě"si:��N�
xMl�������|Q��s���$�^�NH�'�#��O}çJN�Oi#�,��s��_A��9�;�އR��h�in����.�)��yӇy�y5�rt�$����N�)���(��]l�������7�f�0Tz��k�����#8K(�nO���Chq����Y6V���4ɦMi"y9R<�~�蔞�d����N����<����O$�'��C�'Rd��G�S�$x~�d�	�=�|�a<t�#�ï�Mu�'~N	:'�׎��?x|{�!d�F��丑�bt{�P��8y�>�͒���H��%9��>JD��&����y'�-�>G�"Mp����O	'I�$�DJDGŔj$D�X��
�%�'���"%h��B���Ŕ����O��M�DK8���,�Rp��A�e�D�\H�]I�E}�D�">,��H"'t�:=�(~K�elD�YC��~I�z$�C�O	�DD�6A��6�6�/�8;!ϴ�>�<�t��l�'4D���G�%��G�K�N���V�.~_�xm���1Vnx�1��Iv'�cg���$N8�9�<"�ԃ���MY���#����K8�+�����'hG��㦪tjtM��Ԃq�)��wǓ�%Ή�	���z�9�f�}�{��b5�&��f��5���q�'4"�>'HW���=��N>�mT٪�Djʛ�e��N&��u;F�h��i��<>�+���4?Q¤��.�>�^����t��G���F��yu�Ӈ�/�~�D��,צ�Ԫ3�ӇxlvԻ�|jY��9ƧI��|��9%�KTp{�TMvCGH�HԹr�.\���t�8pw�,���kQ�""ĳ_2ϐG�Q8m��ʈ�"x�O������"�%���UDG�Q�8:jt���"�p��#�TDޘ�4��">$N?#*�"Y�JZ�"v��ڈ� ����Dw�¸��I��d��	Cŕ���U��ؔ'8Բ���N�P�r�#��Dޚ�A��GZ����B3�9���y>DeT�c�����;�֧ȏ5Q{Q<mjP��R�>�':�B2�":�DM�D>Dݍ�DG��G�z�'6Բ'����DѠ�R#q��+Q;�iw5btOnx�KO��}ϡ��W�7�s�{(�Ẃߎ��Q����'�O���І�F���>�\{SǵҸp��HA�8#]���#MOԱ.ښ'�Ϡ��w.Q��Ӽyg28:�ͪ?X2|��>A��g�
g����<���n�?p�rx��D�GsBu9��͔�9��n'�R'�-�N��>�E�D�T�����Q�E}X�uL����Eö���;�w��{y4H�!ƾ��XϬg݌�}�f}��k2#:}c>��mf����|ϻ�|���<nN�%�[��r<��9Q�*/�}�~5?�(�
�������D�|���Ժ��H�uS��f��ܒ�V�7�))9�J��rO�V����|��jsh)P���aaj�Vwr���ǽ�<���57��w��Ӕ?s����2��>�X��B��t�s�;S�nD��:�e�Qڞ����'�l����t����=A}L_mg�*��_i�7>ckC�Y�̺yN�������zX�_P_`/�{9�.���59Q9R�NT�K9'#Pҟ��	����F�XϬc_ZϺ}���f��g�~K:���Q=�I���_�ʉ>��ȝDt�C�����D�:l�¸i8Q(N$�Rh���弲�����'ݓ�:]��C�tE�W�Y=���Q�%""r��c����yBV�)8v��ג�ïJ����4:��d���� �"<����htz���֥|��Q����9+�~D�5)�؉��W�ݩ[N�"qܤEܮ+q/q4�R%���G}�D{�VAYD~��DG�(}���5)N�"q�".�x��%}ݏϥlM{R�M���6�������w)C؉�2�h��KvW��*��,u<�RhM}|ԤM�s�<?l؞�N	|� �"Q�M���D��I�ze}@�"P�"p�8Q��9ɲ��|�'i��}ϮIe2Dw ��Rt�~G�T�ҽ��D�'Mjt�,w�Tk�y�_����j�x��N&�����k������^��eh�t8H\�(� ����D�U�}�u9�fǑ"{������+Ǹk��=5�4K�n#��=��9%�D�Ǖ^<����M�"h|H��H�IӬ��Kd�\���rw�M5֪��WI�A�jD~���tOn#�u�܏�+��jt��㽻ޞ�o/x�ٷP�3�&��n' ��\��_Wa9TV��5��n}�ϼ?C���{�owy[~b�b�mtg�\��fyQ,�Z�j�jF��S�c��g)�^�;&�����>��/��U*K�%j=�yg��\g=O��h�[�oW�}��xt{�U�eꪤ�Hj&��e�����oŲ��_I-��)��S�p��u;TNCC��7
�V��$�u<���]�l\�tuɇ}��yƸ�����W��Q�cA���?=xVS�/}�wv�K%�XI;L@�5Kz%�N��j��ưu�E���x*
���mG�-̃k?���տ{�^�����4���72,&��GI��4^��>���a,l�.���3{C��ϧp�����K�� �w~>��g�_��Ǹ�����i�w-��ǷO5���Z+t��v����|��۹�/����w��cϯ9|ܽߺ��n��� ��7��w�:a!�{;���Y��nY�ܠ[K>�!鄡� �N>�쟧{�K��(��܁��s���d.��]둣��_f`�%���v��0p��3)�ڲ�v퐳v\�f�f�`Py=׷"'G�vC4.����]tݙ��L�5G����~]~������'��v�}�5�=!+S�]�}��cΖ���ɯ흹/�.@9��~�g���M�郇r~<��ڟI?d�u۲��1~�"�ܥۙ��?C�w�y7��=�����g���c^����M�Xw����;�f~�w�;$��ٙ�ob~.g������	�W}r���^�=���ՙ�7�f�@c�sۇ��C�eϫY�����:S�{Ǎ݄�e���׋:��;�<1����>�&���YS{-�M��Jx���Zd���f��;�?=����':��&�Ε�3O�N��ɏ.��s��5w��9yv��>;�3ޙ���\�2��.i��G߻����>"fn~���(d����So�w��2�$e��&��&L`�3i����� `F��kM���A���ն�%Q���՗������x<�M��3Z�w;�Š�]�>� n�����\&(�p+��`��k�:Y%:;G'3����tדZs�ŕ�R����v�ВQJh��'���g����M(�@�i�cO~��Z�w��k�����v>E���缱|}v3�5{�S�����1�ǔ��l���D����p��7������j�*�x���V[�n۹Q}����]�dCD~[��9�����}�֖x�����7�m,�� ��H��7"��:,^��G�	�{x��Z�*���C�Q�3H�:���1���_O��zo�s�VX�	���]�8L�sūc�����w��� ��0TK��k��~��K�'���%�FC�3�l����d>=%����:W�1~i�Ɠ��ʥ:����P��5���I�5I|i������̷3=;�5���ݾЛ*#p����wJ�o��5ߣڙ!&[�|�<�;��:��j����Q����
��X;��^���ܿ����~n�m��ok�>_\=Z����g�O�ej��>L�/�C��ѡ�������H`�U���ب}��2CtwS��fV�æw���3������O������OQ��%�a3�K=}ޘiHA����ְ���k��߳0�_�˯G���e�������2{��s�|�K���/q'������p/s3�!�/{��7�3ٞ�o��?y�-y��Wv[a쁤1�[�`���33'w������w�
���o�5~�;��}��^ioM��/��~�}>��:�{O�y茕;������|o��̉��@J�d��1���e;�ڳ���^Ğ=�[�]��0���x��_o�{����+�CN���w����rz����wrG��V&���g֙����ut���n���30ݣ;����ѵ؍[�����]ki�&�}2g|c��{m�ɾ0ѭ=s8��=����a�h�K6t��&z%5�����=�G^�X�ǌ�)D��OOOo��k�����)N�_&��{}��Ҝ�1͐c�l�A�>y!У�d�>�w'w�nO����#���fM��w}>���I�
�w:io|ӵ5��l�a�>�����T�_6�o��~��n���oG=���,�~�[�m�s�-���S+��w*�G��^��4$��9���4y���Ǒ�$wۀ,6m�w��0������7���^�g®���v�]�g���<P�4��it�ŧ����2��|x�wJ%c@��&4Y�������o?j$cG��8u�ێ�	,�n�Ok{6ru���޺n,�)���2�J~��=Ϣ�pFo}-ż���r�ً��d�����%����"eRs9쇣:}3��ݘxdO�џ��e�jb���Q�������r�V@�do�e>�*M���U��ؘj�w0��7`ϻ�w����]o��4ˏ7��.tf�q��ت�ޖ��k��� �w�v�nޠ�6��4ó�؞9�ל�{���w>�^s�|����?�;ɳd3�Nt���?ﷶ{��(��%{3>�X~��՝?O:?I�i�����瘛A<������N���y��O��=ہ���~�}0>�r�Y�O˩{�v_��߶*��M��8\�&�	���<��E���W{��g�Q)�W�1�����ɻ����ˋwu:�At�>�UC����}�w�2ϋ^g��>���g^o�0�o��v/4^/�gx/��ݛ�s+��w��.�M������M���d���ދ�D��wDg��t��a���&+��4}8��zwg��v;$�D��e�u~����_զH���䟾�{�H�'���U:f}��ڟ����ʨd��K�|y�b��G�?�o��7�}n�1�%{�/U��0�n�<][~�Oo|Q���Igs���r/��>��U��5L���;/vv�	�?z��L	���7����i�>��߽���>�<�>��Ф�r})�:wr\ٽ�S:����0��t��nO��=ո8�	� �S5fjȔ��
�7����������{K��Ǿ�i=�k��������Ǐ���t='�uC��=�oA%���aܞE.v�����K�y�j^;Q�J���V��R�m��@�r�s���(�1(�R�]��)cq�m"`>6*�ĬT$B�(�R���ę\���Z���1�'j����O#jx([8ӜhExV�|����vi���(�M��j#�/%L)]%��9T�}8�n(A�[\9 N	�6��C�)��M4:�CuFԢ�C)2BrDҤ��Ukn�"r�"-F7[+n)K	$U�����P�pq�s?���K$@�)F��ڐq��"�,�+�b�6��5V7������9kT�+���"��&��$�KXVWlV���H��)����LM�A19�F��ն+f`H�c���Yh�/\Ǻ�u��\���V
�tM�e��ªp���%$�q�Y&*��v��r+9#�
�H��de(8 ���&)T�.<�f)`�f(��/�4f-����,ŏ�K,d�
����\�u!�U+�c�������n*u
�
Զ5cm�!)��X�(��#�����V�;��'������V{�����lc��q�3���.`c/2&7W�$M;W�Ǖ��|�X�����+��X�Dz�QZD�SR�1We�9U,����U�bbm�Nqb�eR�Mdm(��4��x,��
4��Y�Er�ִ �EdmID:&Gx�2�c&Q�\���n@4[�lS�	��+S��K	�Ў�2SlM�K �T�BK%�ư���qK��˸�L��DrÔQ(��i3nK)�圜�lM��v�I�S�"byy+��,�`V5ȥ��O뙒�V�5hȪV����cMk�T(D5P'������do֮��j�ؿC�qց����y$Xw5~�`u�;*<L��ŋ!86;J�JR��켢�9�r���M��z=�(����SI�AYm�������o0�l�Z2Ď
���J�kq�*�R5�,˗���W-WpZ���n���m��x��=��(��;�Bo��Q���y��|���y�r�����?��=��==��y�O�O����o���UUU��努�V�U��U_"������UU򴪯U�Uz���ZU[Uڴ�U����V�t�{Ң���J��U^+�U�]����U^+�U��_}�BX,�"�AaYJHC�$FB(D�Y ��)I��
R�-�,��`�$ffg������U^*�Ux��U⫵V�k�x�X���iU^��UmUmWj�j�V�U�*��iUګkUV-�w��⮕W���]*��b���*��iU���fffvGu%�"���z�
H�",�P�H(�E�[	-"ԕah[TZ'��Q>[�u�W��j�U[Uڪ�WJ��]*���Uګj�j�j��WJ�����ҫ�V�*��U�UҪ�]�~�t����UUEUUEUUEUUEUUV�tX|��a$*"�`B,)
d����
E<2L������Ҫ��*��b��������V�Uz���եUUEUUEUW�V*�]y]*�UU�V�v�V����UUTUUU]*�t��V�UꮕW��{�p	>$>��B�5�-D*+QZ��!�"H� �
���!@�Z��-AJ�� �V�P
�� Ȝޑ�K�J��n��TU����������S���<�3��d��d�4z����NN���:'�DO8%�DJ6""'��H%��'؞8"X�؛4&� �DK<'
DJ�<"Ȟ,M�blM�BP�p����6!� ��h��bp��	��B""pDO$�"%�b'DO���f�CB	dA:p�&�ѡ�z��~κ��Һgv6�x���%r�#j������#0�uH�&7U�ddaU+U����'`��-�Q.c"�
��6�:��Bژ�j�ƣT��+Uʭu�*[P���"���[3*��:�b��O#1���[���W/�r�d-�B)+��v�Q���!jdt�����uP-LV+k��h:!���!d_�r�Ԉ�V\G"q�1+NZW�Evړ�6'J㥑��`�b��;F�9o��і8DЅ	�JAB�cv�%+���]s��>:��%���dM�*ۮ�
��ҽjE�(&��1��������LL!���H�r�'eq�J��&&�QC��,�R�j�'ibe��^E"�BR��+V:�଑�b�Ԏ7���'Z��n5%Q�$nA��-�$r�˒'�j��OVf�der�q��,���cqX�h�h�n!ƣKh�w,3�c&
��a-m���KD�.	�
*��-t ���Ix�
�p�Q������QJ5QZ���;e��v6V;r�Y�Yh��QRʙ*R�W[�T5R��2UJ+$��!#,�������l(9Uv&�"����)b��Z�v���R�X81�$��-�q���BT������a���^G`�le'��U��8�Hӟb��bq�M��7L�H�5R7#P|��Z�"��ѥH�a]��MGb�F4��؈�m�9Y֝`��Z������P�!�,����UW�!Y�v�9#v��9�mZӱQ��5(@�N���3�^]���}���3333<�U��ݮ}�|�3333�^]����}�3333<�U��ݮ}����z��ǎ8�lm�Xٳ�8l��{�{��Yd$��Z�cx�3,�����[�fG�n�5�Yjy!9%�������Q��q+��+`����YU���A�;SdQ��c��&�.��y���E�ۢ��+*��� 5B��*iN1F7NCPq0q���\M	�:�� �Bx ��~�2�fe�7�:t�v+�c�(��w��`1F?u��a�rʚ.1B�FЉ�WG1rf���2�&S��Ҫ%�4x��'NC�Ī�D6w� M�K�y^�y�]����U��d��6��ьY���v�+UF�)e�aDڸ9��-�������clz�Ͷ�^:kq��F�s�U�%��,�0'a�d��,��ٜ�q�rg�a�n;gMB�p�~�j���ɝQ;�����kˎ�[vY	Z����\.�ɨ`c9թc7�2A�F�d����,�bX�:xO	�:'�Ǆ٢�a�	X��,��b��37.XX��ܱϴf�fr���=1��=5���[��[L]��"�r�3*Z*fb�p��f�D]X��\�E�WhÛ�Zx�Q,��L�*�Yi�
F�]�ef�����;�m����#�5c�?<qǍ��lm�Xٶ���M��phl���Vf\��3"YC7�<!����1�3�[12��ۼ�f9s!tesV��=��[�Ȫ�*��9:�d�!V�`�jzꪵ1���uAR�]��"��f*��!�6N��T����j.0�^�Hn
1&�?:w�cqǍ��lm�Xٶ���<��Z�^K%��D�[��8��~3i$L�x
5GJ�n��H"���Ƴ$��A�@���GB6ȫ,eG+!5G����s���V+��R�g��W��"Y^<��=3w���r�!/�UAw��_u|�}8��X�#1�y�F�.�ӻW�QA�L��(�����a��F%��sLP���V�x���֎U�yBY�s"�9����!P��ZD_�\1:�A�J� �� )�lz���--����t��m��lclm�Xٶ���L<#��V�tr�ܶ�rqUS�� ��+:��v�t�n�4l�:L������h�4n��ˁVVZE�\$0UG'x�1N?����`�寒�[>�p��j&��ի�,72\����U$aG�\ىe�਌^���	Z�/�>J8ag<xO	�6t�p��4Y��qKl���UN�GQ0T@/|n�-ⱋ0h���)�]�T0zr{��]�N���Q�%�_w1��q���9e�91n���l�鹳�C��-�j�L&�X�6�UZ���0��j���G���{]М��G;�	��n>q�|�c�6m�z��<��aR�����⪥��˜����^{�s��k��+���eʲl��yW����ʏM͕.�HѬ
fQӆ9X&��h|�:p��7GhW �:Ys�(Ka������������n={[n��8�Ǎ����_/%��.�Q}k�U	�V(��1�ZҶ�+',�-.G%���r���� N�]��X����lQ�c�(�|����j�G�ET�Ȭ�F` &�r��Xsݗ��+��R��摕6�1w��ܑ����Z�x��F��X5�����M���bL�j�tIJ)O)��,���a0����L�n�..�.�3r�I�c�}z�%�;�g�6��MfX��-:����7G�x���6����::C��7�7<����I����e�D\9�ޕU2`�F˂ X����F`��h��X�c4jM������S����fSÞ�V|���gC��kR�K(j�}m�mcm+TbV������fh�D�V)�s��d�5����f���45����OX���k���N	�֧c�6|���[Wӌi�q�_�Q�p��a
Hx�0�TL&��
�a0�&*��0����(��VG��~]���O�|'�g��/���CÁ��,|��'�k��|?+��~:W�C�|8aZ&	�
�ea���2��G�d|j�Z0���-�*�����¼�#�W�DO
4>4UyS�xg�hr>:T��p>�EO	�����.P�;O
�ex|8eO0�dL+�T�HaXL4VS
�a<eI�I��+�=Rp¸B�k���xSԨ�|(�|�剡2%�xp'�0x��=��aX���3l�qDE~��3�Ʋ�i���ϮD���2��oz�#|}�>�ެמ/���}ru����;�y��}�ޯgN�4�w�D���ze����oz���k�π�^sګ��c<��~��=�{�{ʭ�{ڵ�|fefg3̙ٞ�������}������2�2�{�c���Y������fr���c��YӇN�:p�<'��������K8a�T�iҪ��j��4D��"�SF����		.���I꼏�h�Q�MɫפȻ�)D5�)^�K'I�6djH��CԛJ�WW�朷n�\�iwv�nl��f���5G��\�F��tCM�
`'	��Q���E0�
*Ii�2S!�00K(��bI��c�0�X��l�e�E	����$y((M�FO����R��G�3!*$�����\`g�Rj$������=q��񏞶����q�!��eT��ժ�����ұ�P�v�U]t�kR>Xb��Q�����(d;I���_�Ũ����iR�u�rd�0@�2|���a�2L��ȐI6ʁ�O�Tx�6�2bvb��#
M��]H�P�ĩ%�Y��^��w?)��Q[5F��K�8"�$����r�͊H�N�/R��f&P��2!��^Xy$�,��ijY&"f!�*�@apIHB�,�G�fbTȃ�'�<t�|�c�6q�V�=v�i�k��bj�tR��3�YX�di��\�n<�F�ka���Bų-��ys�Ql�kM��H5�^�Y����)lt��\�:�(��@��uK) �N'+��V���b�`�D䪉�4:(����*����L����!���C�������M3��*�DMT�zW.���}r�q����n� ^����ւX0�&�=
�XND�]��f�	�@aB�%I80��q�ÅL�gJ��>���JbFZE��A(NF ě±a��`����	���}'�ڊ��3tC�4���p�Tk �HͫF�X�6T6�dd
A�ټ⩫.1J�ō�`���ɟB��p�(J<4b>e�k��>�Wvٖ�#x�KtU�,2H�e'#Md���T�m��X�˭�hBȓ� j\.Y|J5�/�j��%]"[b&	�T��x�&���4~��xN���Q�GM�7[�։W�UU�e�VB�ԣ�(>��2$.	luQ~��2��(d4�FBD0 a�R�'D4fR'I�"���iC��I�<���@I�0���U�na���+!�"Aa��B���zܖ����L�-#��guV�Z�$��!�"�a�.��	e a �Q���U�h*h��b\��4��V�R7�D��%��)� ��Dj�+�$ܱ�m���m��c���t��8a�����)�*�axy<UUQ*��ΥQu5Z�2&R_����*$؆A#|!�V��	����5�8!*@�2�rD/�U(�q�Aq��5��A�
C\P��H�UC�@��O�c%\b��N�H���a�4ԮG�K$�P�NTt�7�;���j�w*F+Jj	��RM�TJ��4�Rla���LHo��c	�FN��
�TSE�`��T�A��"-�rU]2�y�"\���7i�����:��������c���ǧNpك�`DE*���[���Y����UU��ՊV��ag�d?B�#c���$a��V�2Ĥ�D.����xI)�CɅ�m��tS�}����A����j�ld��d��l!��hts��UK/	�t4`C��"M��O�3yd2]:`b�Eu����Qh���a���v!�`�C���R��cG�l�+�U�N���
p��<2x�I����HP����;mc]F���9+��J�Jg��J!`��	S�M��<|�Ϟ>c���z�Ͷ�M�v���O����W�al�TH���dX��0�����T|ll�Ibq�;�7�Kn�8��S��ƫO0l ����E�|��K�7p�qn�I������UUQ.g����0�k[�#�nW\�b��e�l��:.��њK����0ٹ@a�g�F�+9Lŕ!�)Kv"[�*�*Rӫ�b �!v���*�� r�v�se�+fς����ɂ��i⡮JlW�-|��D� ab�H�. R�"����t���HD>WN��Pܫg�Q��Ǒ�X����$�"r��ܖ��-ʆG&��!�`����!MQ�eB��b��F�lԣ>��W�Iڿ1�z��ͱ�z�Ͷ��NJ��s�eS"5kCn�O������IH�]e4p�\y-2@tī�M����5ır��Iq+Ma�ũ��3c*Ҫ�B��P؀�7nHϲ�E�3�!6!�H#.n6�����ĵ�-���bČ[��}j2Zn��c�}MQIN�!���QI���	vcq��tEㄠI�B�, A����R�4���^��6���=c�ͱ�z�Ν!�ӆ�y��	�9zUV) �t`��Q�F7K�`h�Ds[v� X�hd�&Li�!�$22K�Cw�IM\�����f���YFk�t�I%3NfKjBl/�˱d�wy�"ȍ`y*��O�T9,k���KS�ޫ�U|P��{���pj��C�?B�N$��`#>�R4��0�X��7.F=ȆMX�0��K�Ka�c��b�fߚ��]��pBm�@��qj�����O���׭�q�Ǭl��6xق�Za{ъ5�7U)���"]��UT�@>K64D��b�UE��ə ��!�����8�>�U4t�V'�wt����կ�!�%�K�a,�
=��d��n��6060�� b2P��O|"�Rv	�%%2h@`�#��K�*OFB�DC�ʒ!B�`�S!<'�j2"����M^B\B36!�!�IcJ˜#HxM��4�,�;M,�T���O�G�+�&�(������cm?��qu6���_�M���mƜcN1�	F�0�0�M�0�"aH��*�(��a0ц��p�&	�I�J(|>	g��sM	�ex�J�Ύ�<:_��FD��p>&�Q0�°�Xl�XL!�t°a¨�+	�
�a°�L"~E~�>�D�������0��F��l|])����娏�\'���O�0_�|����'���>�G�84'�6QFG�045>J<L5S
�*aXx�0�D��(�$0�&3Ra0�0�&I�I��ҍ(��	����OE|*�����j�ƪ�WJ��\\%z`�����ݤ���$�&��ї�Y��ߞ4m]$0ǋ��O*�ce�v=�5�dǧb3ͫ�UP(�#�Dw^�}�[�ފ��'���ʮ<>���l �y��ؾ��L��l�`���rL�5Sh���݊m���F�	v<�[�6]�����=H�{ *r�	��x1�Г+�h���a�&V��s�ُ,��t׼"��sX#,+J8O���0�M&5[�e�d���Kbב����Ӿ�_o{��1�����g�ֳ����r����=3��1��;�c����[�Eެ�hw��}���z�;���ٽ���	�\�I��,����dX)�������d��L&wnz�z���x�b�����g|��C��t��ιG�ٝ�Y���^��3J���R�ƛ�ž1k�N�X͟���VU�V�ُs��^�w��-b���%򙻛�po�u�t�־'��ػ?9�3�nG����8g6>�����WB����WEx��*ت��,���9�`�O#�pv&�r'jpR�ծ�c����6�吅b���9[��"�;Q�F�cad�YUc圐�&�eyaǘ�d|���X��u:����:A: 䮍D�h�;"����v���.,����x�"	D�G7E��o5�ߖ~\V���/{�������⴮s�w���33Y���V��r��3�ffk333��\�9w����G:t�8یc�6m�z��o�+�s�^�y��P���2Z�U�@V8�+	]�e��v�)����8aXG��ڱ��89[�\T���4�A��NX�4㔱G]$d��2�c��o1N��50�uB@�U8D�AQ�Bq����N��Ycr&(�j)�6�Nި�u�\Pʜ�����6�m�Б)r��#�O^��d����4�믫�`+vg-ykY�{ztO2y�t2�h��i�,٢T*��Dq���MC�ͪ+�!�25?7mQ�<��H��)��ı���� �(�v������p�a��!D�f�8�e������f�+����{��	G�	����!��͈lI��%s��@�ϊ��`@�]��.lBP��z7�|�T^��Uhĳ 8�]a����C���Y[%?P��&J��)Rc�|����j�p�<sQ��t��o����8�=cf�!�ӆ�x����8����� pa�����,I�}A�Fꉓ0C0�5 O�Y�>.PO'%�Q@t����)-��u�%��Iaԃ�g�X�ObCSeC{�B�@�B���P=�D�TH{F�J����� ?�r�e��mn��V�����q,�!���l%�pE/M�),�,@���O�})�u;:�F�Gn�4�����|��Z��q��.;q���1���1�Xٶ��]��ݚ�z�ԫ�m���������� òBR4lJK������#�ԚH�t5�@�p�'R�^T�W�!ɀ�g�����P̕P{P�9оh�Q�󢕥lw�%YO;��]b�F���,a�V����b
eN�ɘ}C��F�LA5Y!d�&�%ӄ��� ]�F4������}9G�ycC
5V!!"Ĩ|bh�b���T17��pC��a��C�*N1.���e�c�<|��>c�1�6ڽq����JT�d�c疪��ڕ�Qf�:n��3Ϗ���{cD�ڙ�b$��Qܬ,:y[r�\'ɘŸ\�e����ʟ-��I '�/��J�NOC$<o�q����FΔ�{n���=�
N82\�S�����H�,��Z%Bɛ��,^�Θ20D:!�U�CZ�L��֪zd̐��0�xF7�����R�F4��h��Q��͉�����w*�k<c�1��|��>c�6t�p��<l���L�w9�H��-�����aU�DW�U�	+#��Ӑa�l��1NG Z(ǝBΊ�R7�vn�$'��ƣ�G!UUTObN1�Md'$BmL�]$X,d��6����n-�F��ۘ�py���Z��1�M1R��ɢ0��7u�����˯�n!5���P�*��T��Q+E��.��|,����f�K&�a�����J��ה�i6����OC�
0���3�L3ӅB��w1g��JKɐ�z֗B��٣&a7�cP�̆��4H� $�R��zk�.�8p��ϻ����.�ۊ�q�ZBbN��j����H_	uYSQ��b��ģ0�
*��~��;t���8��1�z�c�Hp�醨5�UT�V�ϻFT;BQ����ݶ�f���%af��}.��0!Í�4ft���2�%Uffe�W��g��F3�1R� ���;Jh���$�	(�1�gʎ�CGJ��eA�sR��]�cX���:��%�K��!��B�y�-���o/�.3��~��ėu�e�ٙ�)�H�]�5�&��,֗1*
�2���,�cOc�ۚ�X���|���1�z�Ӥ8l�Ѳr�P������CS���EC���\߸80��E���J��S<rr�G�T�5��ʸ㩲�D!�0ȘԐ��5��e����j�	�����\�n�6��}��-�F�A�p��6\蓦
H!��eUUӚ��{��I���r�NL�$1�[��sKw[DLt�Ёd1yuE	Mfnl���\2 ��d��X��ӂ4�=k�=%z�>|�X��q�g�	�E�:���*(��d���Jj�-�����W*r�h�ON�v@�9=�ndȈ8����MYˉs�ޙnk�\���,��2�В���P�B��2���3P����z���E���>�M�A6�;jwLP�j�E�L��Pܪ��L�.���8n��ƴ����tx��֜v��c=z���.���yy�TUyM��l�P�&V�Q�AV�*�7:,��ƴf��.�.�!%T��r�b"�71��k�nǜ�|a�P�&dRU����c����]���ꪪ�7���njYc��%n�4eQ��I�j�6�n��~{������fb�Wy��n�����Ss�x4�MnNW��L���Y�!�+9��U'�K!�SG�d�!�A�]�0J�ҋz0 �}�a���a���N�gSS��Oɨ����L��xfqǹ�&����.��dqIA��4�rG	�b}�IÆ.S�����%�c��[c��m�ǭ�|�q덛mN,}j]ԁ	W"�ԍ݈�gK�z�����}U=Z0=���<��cv��l�y_O=<,>���4���f���:o��/
����C���vm~�.'bP^x���'a�A�m��cFf��R��<�R4��d��	�d�b�f�Kn�h���ΐ��*�yP�{\(�ꮪfn.>2t3�Y��GFOys\���d�{'~�������Gɓ����t�_�|����6�"C��(�+��&��&B�°��k��6aP�L0�V��a0�3��L!��a6V	d�C��"a[��NɅYE�ĲY7RC	++F��a0�"L,�&��h°�p�XL"L!�a��Ԝ�
�a�2OD�zK�F������B����G�W�(υ��E=K<4>�6&G�<:	�<p��E�#��i|Rx�����_I�a0�XL�Y�&VSFL*��
�52�I��(Β�W	���_x*��x�W-�´�W�q�Gn4��wgd�.�^��w4��_���Ǉ���w���T�ם��vd_z��{}.�v�OHǟ}�k�ٿl�.��2�xI�6�u��_۬;�8�-��339{��Q�߹?=�g��?�Ū�o9˼��ffo33-WKy�]�gs33y��j�[�r�331v�ڮ���͜:p�ӧN�0��<a���6Y��M��UU j��slY$��T:2�٪�զ�y�r�A��Y�G��ݭ��+(���Tr��5�s�r�u'�a��6WC
��\5���*����ӓ��N�s*�:���X�SGL�P���@��٣����1Ѣ��Mçeh�|vc��t����y|J�22x��lv��6���8�q�m�8l��$e]��UUH�՝�P�@�+P�uk3��6X7]�i^�ȹ����n"�1�8^۵q��72p�G�#,�r{�0n%M�(-��m67�tÔ��6Qp�N�p�����ْ��P��׾�yh�辜>�_ߍMM��Ӈ'�t��ӹ���n�ov���G�%����=q���\q�8�n0t�,���>�"��5�Xe\'
19�2�lF<ʕ�#232'}����n�1�Lhy�j�s��j�V��[��l�̂��1R��dl1�T�XЛ̊�Tn[�*�%n"�SQ�$RBHGYnL�Yb�.��9=UUR,��T�}4��9�٘���6,��I�ɽ�����uPB_���������6zz���Ha��h�tz�Q>��"�PU<�(�u���/�N��rBBL�d0��i��}���d6�KE����:x��,�.V�L5t	Y�n�z�Ӂ�u,���/ȴ������^�d$b�˲"Ò�dv$���Cz3�FD�^�F�3Q0���=c=c�6�8ی1�ٲɻ�	!(��UUT���48r�F����o'a�F���~0j�N}FU*gP�'�g⟆��R��&憋C*0�s����oa��?~]��Ɗ�- �m���k�&��	��Y���/��uB��8:B��&	A�O�>)S'��3ݺ�n1������8�m��8h���i �X�j�)
oa���D��UT��r��J�E�Z�U\Ҫ��6C�.��h��X<Y��UW�>�J���'��@�Ψ�q5�uI�[U�I���,GNZh�=9.@ظ3DK��O��ՙ�h0Q�p�Ɣ\�P�_z�N�N5�t����q��Sl�r�J��d�!�����vrv➶�O=z���|��q�1[8Y�('2Y%��UUHܜL8HQw���i��)�\�)�95E������,dcm[ɓ�s��anr���,MYg�����'� ˌ�2fjYe�ޘʃ��ü8e�d5��HJ�9���aM5tzn�8x���(OYGƮ��4`�<�&����O��S{6�<q��m��8��8�q���/.���#�QA�����S:Ғ�cN[K*r�f3
MtY��i�Q�),Q�" ��i
����^B���r�0�3����U[|hWV���i�nn��[�i��r��3���V.��p/�jHO��+IE�#~T��VZ��G�AB��p��vn���ҩ�Z�z%	�����Y�1J�16{pѨ�*d��D+E���F����4x�T؉�0�#��:Y���!�=���0�3�T@emD�ӕ�Z���v�]+���g����1�8���[|�q�q�1[z��&@HZT�as��UU��Ȝ��܍�=zU{<mޣq����WJ���gƏC2h6wK4Q����$��L�6�M�4M���� }Ulhn�!���bP��mY���qy)��׸^E�������XV1ı��v�X��m7ϺzyCC�L�)��rr�f|�0%��.B��Si�$.��V�����m��=m��1�c����1��^�����!t��͐��>4�m�3����zb��,DD����ᒽ��Fl:s�6�S�::K�ݍFT(0�j�I�&�шh��Be��,�B���Y�DM�blɒ�>�aBY�SQif�h�~W��*��4Cu_yF��9�tY�r|ŞL�#Y�7	fGO�ׯ��������8�lۂl�g�E����'�����Vn�����<�UU��%%��]��ފNiGL�K��|�HՎ��&��]  ��U==����6�78����S�G��E�1�Ð��3$<\,��Y�h64{FC�ѣ����ؐ���f>�FT;<��̛.�hѸz�Ĭ�(������[|�j�x�+��q����q�0��J�$0��x�0�0��J�:M�a�a5��&��a�l�T:
>�x|8�#��'���$�$8aGI�;&Y�Nɲa����5�مa0�a^0�"L,�&*J�a2�0�아���aF(��0�0�!�
�	g��=%�����x#��P���<�(���<_���/��v���kK�ʹ��`��fJ����_����?����)�=o��>=k�L+�2�V	GM��0��4C	�OEO
3��|(���-���yrTǆ�	���{yﳟ#��&�5꘤SI�w*�Z�B���m6R8�U�nA�S
۽�1t�fv��F(&�t�H(E2\��eC�d�U/ۋ�������{.9*���~�����}nu�{�0�\k6w��)����=���>�nu�o�S���8Ly�Cl;�j���a�1t�=����<ʞ8\Ke2�t��źFɟk��F�ߧ(Ta�L��?��z��UW�w��5��v�]�Ν>�S~���_o����ߛ��4��ӹ��}�؉�YN��;�����ts�I���}�-����s�jɞ��D�~~�c�����GZ���]M;�{�ڶ��%��]�٘��V-^���f��O��gy�>���w����ϼ�{Q������D8rǇ���©W~�a<{�<�ii�#�:���w黯����s���7�������h8�?��c��ؾFW��O�c*��Q�\�Gdw��(�R�6�r^	��YT%��eRS��l�r��P 7�#G6�\V$��$M�^r��(ܭ�:�w�>��Q$N�6�I
����5��Ȋ�w#�N�b$��L�����O���SL#�Y	cc���pjy^6�T�5-h��sS_�2�o/ͪ�n�.]�g333/33j�ۼ�/333�v���r�0��[Uګ��󗙽�,��t�1|�������E��8AQb�;DExYsW�Q�<P��RR��FH�vL!NDd�UYc���R���l�Z&[J�T�QJ�q�Q5$�v�J�D벼�+�K �R�K8���Pr;![R2�5`�XX�J@�;ka9(�Dm��(�7E-N&��-8r�A�����Q�6^u���m�mZ�Y}``�r�re�Ֆ�F�U�pb��GOǔL��Cv9�;>�e��S@UZ5Gr��|gB�����U����Ϣ��5�OC�J:�Pf!Ó&S���o�a�!���\8Ub�,D�A�p��V.�#�h��.�P��?lvH5��+�֖0�h�"�E@B��Rz�*DV�������zn�skD.��`VK�6l�����1�8�q��m�z��]�Y�MC5&e�s5�_<UUi!*��ML(� ��9v�wH�����;�TOCSS&��^e��䁠4l�hN��!��d��zT�T=K�c,StP�%*��'Fj�K>=����=���\ K[����T�[j�WMh��jꪏ��0e�CFa�*�������"\4zY�2&ni^φT3>:���gǏ=m����q�6ٶ���Mk�Ԅ�]�,�!
$�{ꪫI�G��0PѓB#�T���&�)�i�ardF
a��B����&��ɣw똤H�QS%���k$�d���9�I��P8	�}�_�B��P��a[,�=�39,ɳ$��RlLMOW�M�����DX\<c��`����
,�=���#��~m�^���8㍶�t�,�z��o<UUi!�=�+U�,�b�r��ad!�Н��KZ�!w��H� �uJ�%�UQjp,A����{����V��hț�7�ɫ�̞�|4���,NHʝ����4�b3P�g$�>F�FO[���m���^���ɧM��W��+cb\R�,��N;~i�nr1_�+�����Q��O�6+��xǭ���8�m�m�]Z��0�b��S_X��|Ǒ2dq<E �Y^H,hl���jÚ��T�5E�X�6)��R�+X�+Pݮ r�Z5b�e��ڌ,QKi �n���uU_Q�ݞ�٢l絞�u�t]��o~�H�l����|���G�ÿU����m��Wy�֗�zC��rO+���e��.�<��F'������Q�9�[E0db"'Ά�\<v�t�� Q�31�br<iK22bf`��ˇi���&�%C�X��kE�����N[%R��I��Gg܆��2t��V	�uOj��꺱Ծ�6|��z��q�X�㧏8p�p��4Yj�F-.Z-|UUi!�h����p�����.�[t@𕳓}���QB��J>���wV7�N�ˇ��s���}���¡���ӐѰ�1�Mx�_��B�L�e$̲V�dbl�bh8p�BW�A��()��
>5�6t�*�ɺ0�7�Z�AyX`a�8h�t�O|��|�q��6ڽx����2�⪫I+E�<�Q�9U� ��1�#���{��UWs��zp�x^Bے�4�2ܠY}��6�m��Vb�x�lż_��M¥��{9<'��Q�.0%]��[(����)Ã'M4�Z(Oqz����}�;B��4d�����.��	�ɳ&̖M(�ɮ����x�f�W�%�^�5�9	RK.����C�>'<����nDG�e�B���Bk�}BZ9�h֭������$���F���z�	�.��0�b�6iSF�g�����u�4X���K����Yf��fN�6O1������f1��X�lCp��D�9e��b3��~W���d{�񎝾q�Ǎ������ᣧC�Hp�g3<y��ck3t�?�f,mJ��m�+j��"�8M�*�-�W�me�9�F�Gh�%en(�c��J�5%��Ͷ�o�
K��.9=�|iom�3�8������s�*�w��N��:�`����c]CbTكʊ��С%sf��g�������d��'����"ӨT�n\����r0��}0}IeA���bWNj`əp�X`74DH�,�">��1TЏ������-��E]�� u̴n^e�r�7G��N��jă���N�3��ɏ��������>q�lc�8�x�j�O^:u�T�sGz���d&���Y{UUi!|*D�]��S�c��gs�ۏ����2p��珖d2'��(�h�1��NH��1=��j͛2%�T�Ta�Q�_�=�+%��G��2Z!\y(c0�;�F't;y�|pM��Xd�/8�!�	�ˎL!�#�oZiD��8C��g�r�[��Il�R;�q���篞��6���a�<'����bx��B	�B"q"'M&��B&��<'�:pM�e�4&�"A6""tD�H"&�D���<"t�6lHhM2P�%	Dd�"B!��ЖX�æ��X�_�v�a����q�q�ƌ��8"xDD�͔ � �"	E2&͉�?�K���3�[��!̨i��\�l��[i,Z%�#{��I$O�h����g�ɝ}�g;�����/;�l�3*����]�mO���O��=>9��j�vj�w<G��z�tr�n�U��wn����?��7�ZG��ȩ��6<��-�6fHb~sՎ�>��Y�o�zi������t����fff/ҫ��󗙙���WJ�wwy�����x��V���8lٳ�0�0L0O<t�D������UZH{M���i����j���/�~t��_�˶�l�vj�	�;�w�W��rf���S�E'��"�]��,_l��Gd-�,�v=O�����2`�c�i1u�`.CA�a0]!�0��Ĩ`�����!�fhFO�a�GY4#!�c���:G��O�<|�1���m�m=xM�[���[������Q�Cp�L�%�ea�L�J��%	�n]�,����DxF���g��&*�n,�>�>������m2�_+�}�Ht����zP�[�QF�	��.sB���.p�`x2d�4Qb+�K90�&ݐ�4C�"eV�C(��ɥ�Z�rdK����hD��5U���m��ù��X"'
w��������0L0Ox�t�'��#M�
Y�Ҧ�	���j]3eCW��7�
���ۍd���Ԗ�%b��"�:$m��#�����i���'�t/+v�m����y	��|�N�~Su㵽[�صm������Lݛ��X���wx��'��xa����Q>^��2�ܣ�Oㆄ���õ�:t�����f}�L�1o-��%��O	�j{5��&�C�=�R���!t�)��[`�!~Xf���O�����L�Ϧ�q���"w����g$	pȇ1�+�"hiLp����'��/��X��5��iQ���>c�O�6��c�q�6��j�G�;�yd�Vʘ��*����	�K���h��<<|x�&I���U�c0�F�4X�L�����	��lD�������2"2¦!�Mm�\'�lD��Ι6d���檞U�e��L�ڬ���r��]4l�7�,/i>���*��J�J۔k!~�L)���6�8v�����;q㏘ێ8�ݶڶ�֯��(����}oG�,��Z[6e��V}UUi!�@�m�W>�k��xNϡ�`�P��\���P���L	���C$*���[��Y�N�v�+�m8F�-�E�ʇa4���&Y�>6P{&:P���Le�Y\
�N#��L�B�}U���f��Y�2��~�5S���pJ!�g&]N?<jm~q��x��cn8�0����C��(�<�UUZD�;�Z�.�Z}MW&�O0�qw��,^�7�F��̒Y	I�MDZ�&Ծ���J�$�}Σ�;8d�0&2�1?`�6Y�\,ȉ�8bh�dO�C�
����=<B��]V�'L���D�u����'�*\�͜hș��5�J��*`Oz0�Iҳ�<t��n<q�c�1�M�������e�j����Ƞ7�D��YK]DC���f6�4S�ck&ř1��2h�[S@4K$�"��ԯ���:;P�y<�m��еmѭ%���=�w�wsnj�fnw0�ͳ�S]�F�ky&�C�G��Zi��!�B�쫲�x^�0'����FC�p�*�M�lG���F��aG��.}�:���b!C��b\��_��?#S�gO�y]+�i����%�4CD!�;�թ.&�p�⩵��.�MT�=��p�fa����0}�C{9=�ѓ��:h��6�cn�m[i�ǧVNY�r��K�ꪫIЖYڔY:߼��xѪ(I�MO���K2%��&E	��χG��1>�L�h�.�l�}�.���6C�HJ7F�Я��_�?��1�*����kj���d�asҒZ*����6'��d*fd���O��
Ɠ0���G�؝�%�O#�-�~����q�n>x��>|xt�����gN��7L<��p����Оt��3U��s�lH䀚��YR�+��8/g8(�,O����~]J��k��; �-t,NJ<n��&�u��Μ�8	r#D>/�Q�,���}��	�n��Qd�q��s�����J��9�5>7*�b0����>�[���2t��m���>clq�6�ն��dڛĿ~��nd��D�u�N8�9֦�UUhM�r1�����:j���9���_�8	�s�����X)\2��l�.�9�z���Hr�}�;0bh4cq`ଆ&rq(,�x3���Tѯ���ǎ݆ϵ��X�����:0�è͆Y��u�ŕw���F������������"z��AE�����G���۷>c�ޱ�tN���tN���D�e�DM��"P��B�D�ı:""x�bhM�lК ��6""tD�H"&�D���<��,M���&�(J��2|�Q�N�blK,D��:]ĳfl��a�0D�(C0�a�0�:?p�%�(AADJ(Dؚ�eI�ֻU�kaz�vni��&����gPR��j�ڋZ/�n@�G_��H�rF�X��hu���uK�,����A󬕖�77lO�Ή��	���,���;�ՙ��<T����0���U�(F� 3��N��:�m���1:��X�v��⸘��eW(�����)[X��y܃�7׳mT�g�����_�_��������fͥ�T�s&��_woÒav�ʡ�|ßW�7q���L0r�V���j��>y��>����2nU�`�+��T(߭��Yn+�zjf9�/��v-�VYj�dV>�km��6K(Ьj�+u��V�Gkm&�����r�ɊW\
����"i�§$�9*���-
U+s�N/�^2[���U%;p��q1:��4:�-��@��m���������T���(�i��<��&�R�T@X^�x��u*�Z����+kz���Ӯ���U[���s3333�J�wwy�����^�*����fffff=ZU[�����gNY�`�<:YӤ:'����I�]�2���I�lQ2V�c�V�)GTQ�1��P~��U�m�`�@�-�Y!�s`Gl՚*�eZԃuYP�nJ��!4uf<�G\&ZN
׹p��XG�rL���VԔ��br*�
��M*ȣ��dO��g315+X�'�աiD�c{��m����w�t��������{�&N���{�e���m��{u�F���AM���v�8=�xr���~,T��u�\O�D�R�5�S^&ˆ���=�*���!�]*�Ӂ���zL�����*���!w2sWt]ݵ=�����S>����s��R�����+r��F�^)!�o�S\:y�CRF������z����z���8lp�E���;UUhL���Y���`Y�Q�N���<ٕUF�Ek�'�d����U��sP�ϲr�f&aP�`���hy�E���ʪ�R(�f�p�ܯ-�Z�Ikk�*�,.�j�6kߡ���M�_�m�zd2}��gM������"��=8d��O4qǮ1�8��m�m��L�V���e�J�������'�{�$�d��mճ�w?SǊ�<O��������+BD��l~#�p8er��g*�_�_-KT�>��6��m̘���lxs��]$fD�q�Z�|�NM�,��K,����1�k&�Z5`���]�0k�o���d.P��?]E*3�*EoJ���Y��>u���s��8�o�6���1����Å�:C�pٞKc1]���&�kg;(��Ѣ�;D����(�ޯ�#�(넣PI��M�7ST�2/��r�3,���͘�?qyo���bÇ�yT]`vML��'���8Rz�;(2V�;����%�|�N�6tXd�OB�TUGAs"�(7|�)�!c�RC�.�J�`̀��T�f��
S&�4l㏜q�m�8Ǯ�m[i�Ǔ��O�O����ebqU��2�Er��"(�6Yj�ܘ�k�[Zkm�����SI1���Ř*������H[3
 �Ƃ:�j+��)(J7���m�����{<�-�ǘ��2+-�b3���O%j�X�,y��۽�˼*Q�ޒe|{V}H&��Pp�h@٠�(�^�͂4'�'���d�"6�"�}�3���5�S�����>�9��5�QU�V�T�W4}�N�̘3�Y��A�1�� �rg//��+m�<��]OΖ<��=m��8Ǯ1�8��m�m�����o][VT%�\��ͪ��'�W(�RY�L��ݥ�ST[z�EW�!�.���G����O����SA�1�Y���aGa����Ѣ�m�R���
���P��d�60K�9fOH�V�g�G/��h��@�1p毗f!�M�O��%�77�Ag�JW�)Ab��6`�v���l�ك'ͽcc1�M������Kj���ꪫB!*��!��T!�h��AFC' M��ډU\ک�{����rLb��h4}�x�0�-nX'cLLl$u�yb����B�Z>:xl6klR��j�6|���ld~�u6����)��j|>�N�j���|AZ���p�!���Tc_-[�Ϙ�ǌ|Ǯ1�1�������vRw�i�sM��Q�k�ꪫBp�U�MѺ72�U4�H^�{'���[��� l��ڽ��?My5����q�&��\�s ��C;&`�>��l��i�p8L�[��N�g]Cr�%j'�ɿ+����f��|c릵;?;�Ξ<��'��c��z������[m[i����Ny���o�4�&:���qd�������}��+�D��K&���W0D�9-t��+d��ٝ���*��'8��X�U�f:�"N0��u[�\���9$�f]�Z��*��<���� ��&��E��f55�,��C	��9.V�����ѓ
5����@�t�J	+�=�mK���(? �Z=��LާLό�
(�/��*4rѪ.B�p�9a�0���Q�F���M��I�%���b�wۻ���]:JK%��B�͌1��N���ߝ9m���6�ǯ�����d:'��;�4�2`_t��s�UUhM��_Uzl6{��#�Yvj�_\�Cu:}4u���1���&�G�0�<O�ɰ�s,.\+���G�
t�C�BӉں�ܘ>��ܠ���J�(��Fۥ�SE&��Rl5d�𻦦M(h1Ma�C�!�ɯ�z�}a�S��͸�xٷO=?D��xO	�<'�DO��"A6""tD�A(M�"	��pM��6&�	��$b"'DN�D�"lDN�̜�؛4�F�鎘Ҳe���L0���<Yb'N��X�l�F$6a���"A6"'��0�f�Y��AA(�4Ț�����I͏}�s��[_d��?�1��}��%�I�`�I��'���_T��Ž��U��lNI���7�9{߳}U�u�Ŗ̺=Q��8��+k}�Y���~T�+���+�ϡ;�}�۽>���u���?�or�wݿ-���ٲޫ\����������}������Ӧ�K�l�g�Sɻ��ŭ���rHl{v7������Rw�IL�������~�9�*����fffff/���wwy������b���ݹ��������wwv�O�YӇ0æ	��!Ӥ:'�Q�ڪ�GhZ�r����$����boK;b㦒h��'3���s�}w�\]ݘ����k�Ù��3�Aɰ��J�l>�2nvns!�S���}�&���i^�V�Z�<:�G'Ӹ�����|���mӧ��Âp������V7���}UUh��<�hIgƎ�̄�K�z���mQ�ڤ�bR�"P,/8-b�Ės��Wd���Q1LB�$8Q�t��>�5��\����Av틸a�����FCf������g�;O�*��kO>�<��cq�Ϟ�clco��m�m{o�{:����bn���ւb�k�E��+�W,Q��SW0d̓�j��EcJpJ����*�jJ>E�Zܪ�mp���D��嬗��m��N6��Ι��X���O
��	�"�\�������S���^�H]X���ˋ�e��߫%]��N�5�~.&c:i'�����NfR򪒩����C�7:,��2���B�i4�d��/~ir%50��+j����wn.�蘞�䇏C3���M�X��uj�����Ͷ��cq�:C��6{��On��/�������,��8fl<Sd���3Ax��=�R#XK�����ss��������u��ќi�d8CD�ޚ��0�$i���n~Ib�T����\��C�|\.��U��rn�F!@�ag�������F+Gş=|���m�mǪ�j�^��:��0�h�S&iڪ�CG��F,�;�L�����=Q�5%͚��Q��g�%��VyA������{�mn�r�`�JH��(dÅv��u�&Z�c.6:�KQ��O���s����Rh�36W�8��x�7����yp��l�
i9M��r5<\M�6�t�|��O\x��ϛz�����z�����;2��%⪫F�f }�sa���|O�����K�??ﭐ��Pd#�����{�g��ڊl�d�d�qi���I�!��K��su�I�6rX��r1��F�u�O-��8�(�a�x4���>&���ӷ�6���m�m��m�m�CT�&�?/V����A8Y��	�ÑǑ9��q�(e;tJ�5��k�fL�p�V���lj>d+R��J�3�G-�0��ʕ�m��`K�UUZ7G{�}����31����4ޭZ]���sy�/75�i{���r���Ukj�9�A�����Υ1.Q��8`.x�I�7L ӡ�M�w���r��͜溾��97'�J9l^��v�؉ ����h�Ѫ<����H��Ț�Ƭv1������ާU��K_���;�h79���ӌ|������z�����3��2R�#�UV�����0�#)�$����L�s���na2�/�a�s�6f\�d���:�j�Ֆ�h�3�I�R��sM��we�*�ᑉ���<����%-�E��*�XR��C�sa��UQ��)��&�ĢW�j��4��E�_}">:l����1�1��m�m{o�m�4u��:��犪���!4'՜��ف�bp+��̘7*h1~]�4�;�����������̾OU����
VST�P��}n�[W�3��`�Pp�	��%�sIv�#��ed08�~6f�PQp�,77>Э�0�G������珛z�cq�:C���dIV����B������%�Wk����n�+⏨��B���5���˖��m�b0��m��[Z����(�g}��2 ��p�ha�这2W��~K(8���J�7�*��l3��=�Έ���_]�.l���]�]�nߝc#o�ޟ�돞8���tM	�'���xDD��:YB"P��:P�P�"hDK�DM���l�6&� �DnDDHxN �O�'���؛4"l١6%�d���A�6t��N��,�blH&af"xN �D؈��<"&t�,�Q����� ��&��e�Zw�4Ml��j�f
�K��0�O$b������vX�a�!uX�8�ȋ��&D�V��F\#����#����޽�Ε�o�5:�,B�b�:��Č����TT�Y�r��*!�,--��m3����!�-w�8~9�E��|���1m���ſ��wo轞q�&?!-��^joԴ��"���,�����xS��{�v��Vv�(��jozL�)��؉f
��}�d#E�H>���3{��z�*�i��{.VÀc�K@:�=���85x"����E���:v���k&
UD��9�	�bjz�$�c$͏�1�Nn)V\LL�J;X���N�_+j>0�nH尨���G�\�n��QR:�dV���%ER��2��]���j�u@r�B��U[c'
��(�r+�����.#����]]�D�L�< �	���X�C��3(�tj������u����e�2F�Cj&[a[Q�8*{�ݙ3�����ݿ�ffffb����ݹ��������wwk������*�����8t�ӧ0�xD�Hx��T_��D� G�*�5Zc0_�Ǎ��r5+�����)U�V@u��u��(�:�-j(ێF�v9w.NH)�Fa��c��R
��-̛Sřx�VFKƎI��R:)%Q�)^�6f�V�L!�u������j�I��⪫G7n�'3]sk�.o��5�7We\�r�2-n�YȰ�ZwR�&,��˥���P�ӱ�p��4Q`��{?N1�6���ߚ�~/��v��ӵ+J�5�*5������yθ��#��ԥ���pQF�g��'���S`s7Q��7��r|���[x�ǯ����ۤ:p��d���Z�%�]D��Ua놥�
5���l�nTcFF����[����4pt��os��u^�11����tC0�g��sأvX���g$MR6�V����؏�Z,i�J-(�h6bs�{���0K.r
�<E���>��G�6ǌc��m�m��m�m맳8�y��w�U�ngb75�ycE��9'g��(��rf&�J�6	����Ó�bvfPz��-n��*���݊V|xΕ��6	�ƼbtOu���6gS��,纬4f!Pf�g!���d,�K��	�!c)��y\?%x���ͼq�\clco6�8l�UIxUX}�Μ�C�!8ꗝbX#P�QV���dd-Ozj]ڶ�wht���6Ot��̖L���������@�1�P��A��0r��p0:w�+�S��Z�4	.5gN�}(L��Ū3&��)�z�HcQc����1��1�m�m��W�TO�_�>l@*�E����蜹�c�k&H�����r��ة&�DA�J����;T�ٖ��Mbu�)�ڍ��⩡0'$B8��ܝ� ��+� 8�[�]��{�ܑN�;�N�̽ћ�����oTk�v̜n+�,��h��к0�Cd��2h.QާN�T�����Q�^�G<�#�g!�2�6`������`���{EK�E,���2e�a����,cw��>,�$���f�<<�,*}��k`|�2p�̜6h���������t�����7]X��¡R������5'Nuh:jT��?9�����'����7��mWo'��ѣ����m�݃��8(;bV���q{����NΛ�D�������(=35'r4�09�,�͘k`�x}������Gϟ��c�1��6�6��շT�����q���*$���8�ձ>�l�.��˙�5O�L�b"���h���j��f!��>2�xԪ���FH���HR�X+�p�)L�tX��s��⥘��'�'ȳ�"�>�o`Ȉ�f3U���@jk&�&���7��w''"��w�t����q��1�1��	�e�ѱ��J�RR&�V��\՚3����)s��K^�2�D�FV��YUkC�V�ե��Q��Fl;�)K��V%���rNCfL�\���gjn����:�i�Y6���J�4�,oo<44�6n|j7ɠ̛OR���)�8ƪꃐ�786T�,�)�q�f,N�Y�������yuN56���*�l��B�%.Gn:8�����CY���w�&��u��J�Z2W̔�7�ʶ�m�C����:���I'%��c��2֔a\j� 8��9�9[Um���l��k ˳.���9[�Zr�F�QTk�@��"��!�wx�ٳA���l἟l=�MC�(fLCP��Wȼ�Oy�A�����aQ�� �FQ��x�YFk0a��A{0v�M%t�_�fK'!ءu9�'�[UCT5]��D�9'@�2�������M�q�<q�\clco6ڶl�>S�R���m�,Km�+�Z����-UN��n3yZ%_�in�ԅ�p6j�]��p���(ٶ,��x�:b>��z���%`�5@k˼��w�t��]��AX�7Z�\QZ`B����x���<5��+�뇫�v��gŘ6x>�̝4d��f��]]����xO	�<'�DO��"%��t��(D؈�'����:'�f�٦MA��""xN!b#R&��D}"xN�bX�f�M�%�D�>C��BA/RpA��Ĳ4&�x�<C0��0�<'
DJ�N��<'Kĳ���F�f����sF��J�數��tڀ�4S��U�!۫�_�r��_��<s�36���{����y�Ν�����nfz��<�w��ʁ6'������_��MY}�甛u�������l��Q׊z-�}n����^�/�Osء��ǆws1����ۻ�5��������Ս��Fn�vRO����Y���߾}y��׏>�_w�W����&I��}[[~ۙ�}���/k�{���۽�Vw���o�{��U[���s33331V���\�����EU���\2fffff"���ݮ�p�ÇN��<p���6YxUX00t�ј�eA��j`��7t��enhČ4�p�cB��$ːm'��Yv	̴��5A�\*�gM�d�BQ�,̠��&����d5*4c+�J�W�aڅ�G���̏�T�ǋ<��o�c6���m�m��V޺=���������4��EمU]��?��I���u��?+;l�i��Q?�R��L��).)�˳����`��`�.��!u�~M�t�=��>�Y=~�k��gL�|��`U7�t�(��:"�r)�ew�:k�^L��]�;pjg��,���}�mr>c��8��=|���͟N�����!�S�H̹p��.�ep`�e#�U򺰸Ia�Fe/&:�N���rȳX�S9'+ǈV�v��4&��S����X��P,] !��~���ۥ׽�]���V9���nE�����U�����`���;>b|0�6e�,x2M�06Y*$���fN����MB�x������7`2�xdt�y��'�QO��v��ic����F�y��:]�s#YI3%R��� QƫP#���P����WC-�����6�lx�o\a��æ�C�Ht�u�J�U`�%&t���S�C��M��`�u�J��md�"�#=QVcFa���U�t�`՚�!A�n�(�Ik=�C�[ }_U��,��ͷcU�7#�K*.�MQ+��hʯ��.�S�չ��خa�ȼL�Y��/�4��*{��y4��=|�m�m�m�yy˪,���I��WD�U�����u���gr|���B�>�������x��a���h[�B���9�ƥ��3�"�Dj�4�7h[�Z^ɷ���C̖p�ꪪ7:f�{,�Q;�-0���#����n6�1���4|8'�Q<�0�Z��)m�ޕVs��evhI1�E�;��P�/�s�|��(��W�_.[��R5/Y.[��&�m�S�����p��S�R���%Ԫ���A�ɓib��F�+FÉ|�4�/C�(hЦa��,�Ǟ]���k%�'�'C��ѩ��l���a��2x&f�.�*�7��p�4Q��Ǎ�	�:Ɂ�:p��GZ�v��Q�t�࣑��Q����s�1�0e�l�m�o�2Ʀ@n����vX��Xڭ�)jB�㨊:W �h�UY+T⭷���|��
�\�[n7d���0��ԓ6����j^�`��^k�[��z6]���CGU�fa\�{�b�>��T*|fK:sȪ�J*��2'M�OL���jt���)�6q^BE8v�j�P�Vr����I�&��F�9My��I�F��u����JT�����#ff�K*��̟��N>c��Ǯ1�=c�oU��Kz���[.Ց�K��]��*��L�sɣ�Ԫi|M���j�a�9�|�77�>�JJ����xi�Jipɲ���;S�8��e��mdv���8䪺�'�"H�SS���A�U%jjM2hc5#3���Ӵ]d�H+.�|a��N<tD��Ht��;1��Wԭ0P�Ubp��sй���2��a�
�*eQ��b�N�8!�&BB�>3~əI�7f�%Q+YK(�i��o9��ub����"�-C��Cl�ɰ�`jp�Q�ףI�B}v5k�l�S]�!��X��A�!�a��Ǝ�4h����tL!ӆ�r��*}h*�[.��UVg����J2y~���_�G5~��~q��
��&F������4h�p� �������.l4w��3��tL�U{;�e�I��/:!�y7EG�g2aɫ����pem����':�#!þ��_G�C矺~����ڪ
��I h��}/�|P�����($����b�悂�"
7��&�LOӫ�)��Y��Y	jIjE�
n����""0HĂ#��q
�#`�`�DbF�b*�,��YKT�R�,F#�H� �D`�
K)eUX���IR�V(bFDDbDF�Dd�E�b�U*�*RX��T�VR�%�Ub�R�,���J��VUU�K)b�UU�YIb�����)J��e,R�X����X��DD��0DF"#�A��#���Db0F"$*�*��KJ�QUeR�D`�#�A�EB�"#���D#�"DF$#"0DF"#�J�T�Ub�������R�YK)eEU�UX��D� �b"1F�b�V,�U�UeU,�� �������UU��X��U�"A�"2"#"2""���b�K%UX���%UE� �b""0DFD�����U�J�T��*�eUX��Ud���X�#DdFȈ�dDDK%R��Ub�V)��V*�d��J��T��U��T�UUe,���T�bFDA Ȉ�b�J�QUb�����X�U����)b���J�UQUR��R��UYUH�#"#DF��UT��*�,UR�YR�5CJYUV*��R�ʪ�J�UeUUE�J��#D�#�DF�Db"(��F��R�����V*�ʪ�DH1 ��DA�Db���VURʊ�J��T�bA����Db"1
@*"#b ���F��Db"1�A��D���D�"DDeR���*��EU�JX�""A�"1"#DDF�� �#b	1���$���TST��(��Y"�$QbJ,�E�(�YғH��QIY$QRE!EIX�HQBu��N�E�G��	4*D��J*D��J)
  .�6�,�I4B��QQ(�
,B��$QH��P~��'P(�Qd(�(�ED��QP��E�ƪM!E"�"Q`��X�T�*EJ,ғQY%H�Ģ�E"��E"��4�ԅB�"�
,�,�%
,��B�X�T�T(�(�E�Qd(�P�(�EB�
,���"�"���֚(UQd�%��YJ��U,P��)b����X�Y�Km�,��K)T��K)K�K�U,��%)b�ҩh�,R�i,����X�R�b�K%*�)JK�Y)T�Y)b�K%)IJXR�J��X�)b������U,��U,R�T����R�d���d��U,��%�,R�b Ȃ �C�b�`�)b�K%*�)JX�JX�)b����K%*�RY)d�����U,��Y)JK�,R������JU,����JR�J����,R��JU,��R��JR�K%)Ib����K%,��,R��RY)T�R��K%,��R�d��,R�,R�JR�J���JJ�����R�)T��)e�T4��X��b�)T�J��R�)K�YK%(YIb�R�e*�RR��YJ���,R�%�T���ER�U,R�-*�R�eK)T�B�b�KY)JX�RX�(�JR�)K�J���K�YJR�*�R�,R���,��T�,��ZURU,�Qe����K(�YJ���,��,RX��R�)JU,�)b�IeR�YJ���YB�e*���YJP�E�)K)T��RX��b����,�RYJ����K)TYJ�e*�)TX�5Z���QhYIb�R����T���)),RX�QIb�X��X��%�,P�X��Ib�b�Qe(X�X��%�,R,R��Ib����:�U,QJX��H�Ib��),RU,��"�YK),��E�,���eQT��e%R�K(�),���Ib�Z�),Qe*��YIe)V:�����(�E���Ib�(�E��(YE�,����J��*R��E��)Uj��YIb����w4�,T�UUJ�YK�UR�,�e%�X�e,RYR�*R�,�E����֍���w1p��4B��?��Ɉ ��(�
F���bƻ�z?ֿ3�k�__����P�b��C���uψW���/ܝk�7c��߮�!��ǻҘ��Q�_�ߋ�s�mn�<���s��_�������y�w��Tw ���������������DO�`�~@@)BP?���w��.~���C�B�B%
n��~c��_���;��!���@x�S����$�a+�Җ<ҏ�� ݟ�ߔK�XY��M!�}�))>���x+M^��\9y�����0�s��a/�`���}����%$DTB��XQK*���*YtF��Y���8��LE�T| ��A��D�������M��5��\w�c��N���� �TR�i�U$E�X$����KJ���ҩ ��
)-�g�>�"i��w�zb>�z0}�p<�@,y����S�R?G��{��>^k ���z��%��?:�3�އ�C>��{����r�Y�+�_do���>M����/��]�@?j��q���>�G�'�����>�r��ֲ߲��Q�y'�~P�w�h ��p�a�TU�=/܁�ϧ?[�(-`=Wto�-�p��m��]S�b�Å�!��>�����H6O�'��S�r�<V�RQ�J|�|��uz>F6#h7,���K��8����r��I�{~/��,�e}yTU���� �ϙ<? >{ C�wl���,z�rY"�|獪z��O[Hx����g�� ���G���G˰�-�EEP�}���������_r�� ����G����q��;��w��/��g��GI �!CߏO�� A�A���sj�@=������;�d;q�,.S=�v��nz�**��?a<�vH]*�O5�=��?�P��j�?/�A�xM��	=D
�K�aF��t�\���/�"� �ي������+�_f	��iDN���st����^s4�'��0�����Y�*�,��rk������"�(H�� 