BZh91AY&SYl����_�@q���"� ����b@^�    {���%5�mUCZ$�a-�Y4֭a�SLDI��l�EI�
֫Im�B-�jє�jѤ�KaZ*P��[d(��ZF��&�ElЖmaIf�e����[R�6f�UkdԲ�E��jچ�6���,f��լ�E�U�[flՍ��km�6�	X�B��V���H��VSV�6��Z�l��R�mKj���mX��6iCQSBlZڶ�l�����PU��%[-+M�mf�m33Zʶ��S-����F���3rwem����fX8  wfz�$�v:V��q�
(����JAU�-]5UM��T*ٳu��5 ��zv�ڴtI�n۲���ҌH��8�	��E�M���Sm��  7v�Ӡ�@0-$d{��@yR����ۀz��Pm*n��"���d�� ����ҩ Qw)�PJEw�p�={���-�*)���l+"�p �}򾭃�=�j�R�H{�ڸ:z R��^=���枸z�lIT������{���R���W��>R�mAKξ�|��C�n��>� @|�&�Ze[j�i�4��| ���J��^>��=ZR���{��z9(w|���+�Jzi[�'�O�P�}p:Ҩ������(�>�Ͻ(R�}\uZ e/��A�U(�=��M�+mmL�m�m�[hJ�  wu�BT�[�s@h��y�U{i�l���U)6�ў���=exw�z�Ezg��z�ԥ*��� ҩw��AU������]�Ǿl�բZjm�j��m�l�p ��˳@�l����z���Z��AT$�O��()oR�]%J�=ǥ�;�G��qѧ�H+��w�(Q�����T�F�n�$m��z�ՙZ��2��ҬĳjZ�p  6��������A{hHW�{ޡM5��P���^wSsЪP�=���J�{��n��ק]�2�H�����\ *�w���@_w+�3j�YYY�jٲZ��  �} ������^ۀ ��x(
n�� �W ���Uv��(wy8@@�� ���m��
e��SFl��U��f�  ���A��=�����uT=�*�(��w�u�{n��\ ��ࡠ9�\F�9��Ω�ejd�i�����Ti�  �� o��=����^��� m���� U-�8 ��
s�� z7��
�9�:�{�       j`�*�� �C@i�Od1JRU�a0�h�����)��	JR�� �` LL�FD��R �� �4 ѐ��h���� &    JH'��O�єi�F���mCM;�??������k�T����?��1�ȯf+��s���;��e�l������;�   {��� <�*� *}Q_�����  *�A���3��̿�����%�  *���UW8� *���%O�_�y����|��`N2��aO��?����?������'l!�;a�C��v��l	� v���l	�;e�3�v����l!�vȝ��l0��(v��vȝ��l	�
ze�C�D�;aN��	�;aN���;`�@���v�����L!� v��'l�(v����{e�C� ��;e{e{e{`�^�C��"�T�ʪ{eE=��>���� �eP{d{`P{`{` }0�=�=����N� �T��Q��U�U���Ae {d@{e {` {` {dD{a{eQ{e=������ʂ�Q��U��� �ʩ��� ��� �*�E��@;d8���"�Ȃ��(��*�ʠ� =����N�US�S�U^�C�P�;e��@�;a�	��;e��D�{aN�C��>�3v��'l�� ���l)���;`N0'l��v����l�� vϦW�P�;a������������^�s�����l�Vw4)6�m]�cn�;�uK.^�ouพ�@�8���Af�a��
�\�0�D����sC�W�lv��3�\B���WYD��Z[��a=ؒ�M]��PI�Oe��Flc�(	L�YpI�25b���浚�����"�OF���F����ʍ^�sV��eLɯ�ۈ��v[`��Z��í���^m3b���!nG96�#K�T�X-���ݤ�3Vڛw
�4��P�m2��,K�8�9�������)61���w7VǮ�,�"p:N��f�)-�Q\�op�jݕ���(��P̼��໧�`[V���vw���b{j�{ ��F��q�����"�o)�ˎ����
�J�|��ôC��Lq��������j�9��H�%2[��T��c�Y��D�1 ���S�����4�olM��iXku��:C1'uu!�[�GW���Y��jn*�����̦4�'�kML�#pU��Jl��(]f*AZue>��&Qf�
�`[�[G/���Mщ��<�ɑ�n���U�4��L�*X�e,�76�՜y ��^j��zb��[6T�	\�#1a<�`&+BՖ����1(��ӶH�Mց�qd��s3UX��+N:9��)n+�z��n��B[��� ��Id5��:�"���xq����F�-o1*�ä��%:D1S0�[�v���f*fx��M�c~�ں7Q̫u/rU)z�Yա�2�[��*��rA"�p\N4�wL�K�h��Zʱ��z��X)T�ʺ$߱���`��G�C{P,[�O#(
F�M��	�Y�I�D]�wNf�$V�A^��J��'kN�,!l[U�2�^��.�)�����	�Ҙt�ʪ�荼lЕ^��h(��^�r��^A�g58���dQϡrT6�������`U���n�v�)��RsA��QۼX*��q۸u�zk�F����$E?�X��J3@B`�f1�!Lr��yH!F��Y��O].�Y��{��B��Ӫʕ�go,
��"��Y� R���1�x����3q-��1JX���i�+V����Y6ƀ��Y55�ճve5�+�O*��u�[��/3u�lQ���B��:�F��q��x.���ł��#SU����U��k%�Rӷ��a��'P��6T��@�vm3z5��f�梫"M@�"!��*���ӱQ�1n�ot�C!ٴp�dk�2���S<��0<9%���CYW#��Yb���$Rdu�Q �J'�͛n�eK/E2�hP	�LM�r�-I�(]H��ga'���S��2�Vl7i�Y7m�.X�����,�Ë��B���[e�[e���kH���h�̙�D#{01O۫L����5D�И�T�zu��I&n��ײ��pӧ��u�{3��]9���8݃Z�֑�V��Ïv��̘@�|ָk͑� ۬� �Ѹ�$���sxA��o.�Rd���+�4Xbޱ�����漵eK���հ�e�5[�Ѣ�A��M��6o�4#m���mm��p����u�
�	Nl�XR�n��w������V�V ��m�u�I�Q��Ѧ�ycj�H��ͬD���n1����ƪb��l���1�+���c41!� �H�(ډ��^A)`C�A��mݦ�5X6�,�[pU�v��V$0��͛HdBӹw[���8����Fƶ>� �;X�,��1UE�1uqҬ��5�Y�Ơ�vn6����4&k�]]hI��e��ZE�L�W�;��m��VͧZ�ӱs*�e�n[9�F��St,�9��As0랽q�@�v(G`RŘ�d{HM����e'>���������^�M�ul���[���Wm�����֞Kɥ�(�Tw~t��1@�6+0�O���u�kS�kn񍧭�M^ӎ^`X۫A6�ҍ�u0鼽%b�����N0��c̛���f���,�"˒�K5U�6��w���˙X�%�F�hs���*9��km!@��i��Ev�N��4H�uZ��`�t73��rJق-���c*���u.d���2�)��D�FxU�p�oq+tF�����H*S+&�%�p�y��P�]M�yy)�+n8q��ʼ�5k��J�r�M��3!�.�.����,C�A��a�й�ki��Wco+]��M��M�{xQrD���A�b.�Ԭ:��S*;u��a{[����F\��Ͳ����4֤���:�b;���`��#�qkU7 {�+m��.T1ӡf�aDֹ[�:[H;�/c̫ٗ@-���əL9)c�Q��@�!�U�Jv:2*ܷz��&aY���� ��!3�t�v�Jt֋����-ג�965����mW$��n]f:���2�\�E'�oYw�Ħ2d;�9�"++����v�. Br��j�F5��ӹ�BD�Js�C�^<�q�Ò����8D�����J6�A!F�س%1i�4/i����ۧY��A;��u�j��Si��EcJ�{k{��ĳf;6,��P"㱷Gm�L2�c+(Cj���/dObt�	r���J������(<	e4P����O*�a�v�]�l�YYc]<�M�h��D��xC7)�^bp�f�.��]ij曍k"��T�E-U�C*���hځ@	jb�a�转�cU�M O���`�W^6z�qv1'�� �I8Rôn`���+ִ���2e+[��a_h`Qq�)ک����	L�0l���[�AmnZ�lV�7�oe�w���
ƅ�H�v�h���eɭ'n�-�U%����Y�2�����CY�4�	��n�����ia��$�S7RKń0�it�; m<uf\�m_*�qx�m�2��UN���;�m�Y�v�e�Lz�jZ/��E9�32�;y��v��a2�~��\�.�'�(�,�O́Ӵ��ǉS�m�82m������-��T5�u�@�׎����Z�i�,u�<�1�J��T9���!�3hɀk'�$!\�5��^Zf[�G���fhǻ+�@��f�DN�s4=�v��Z8�x
Cc7�rh�0KB�8�7�P���ۭA�X)S/Y�-�rV�[[@V�2���ǔ�8ի��!�7kD�Q,�2d��w�=:Sf]���P�ܓd&����3��ᮊ�����Q������T*`����yf�P���KB͛�'�Lg��������م]��V��r�S��{���%5��cj���j�Jh�Ɠ�V�n���z]^`��2q�>D��+0Q�il��i��
���j#+.�Q��7�=��$�״�%�s�i]s4`hƲ�+&��a�Pm�b��wv�[�ՒC�����l�mc)ݶr��~)�c�!y�8j�7&*	����kc]�gu���Z��ot�B��`��k�XG`�c�,guPiP�l�%m`Vk�ͅ ֭��lF�!;�@�,��R����Ճ��[6����&M�$��nk�.�:�u��3p��F��l	��z�oEX�_,8�k�n�2S*��Pڷ�[����ׯO ӼH<*�.O)�K�3h�:e�
z�9BU�ׄ���B%wR�j�'�su%, )���I1����j���wY��6�ɩ]��fQu��15�gB�H��K����a;�ӈ���cZM�9���4�#쉟'��z Ֆ²ކ�6+YW��F�b���m�'Hki�����g	�$h�m��f�C6�ݛx��܌c����\34a�E�֭WZ��mՑ�Y�&�3�oR�m�i�ncoq͆�*)S*�Z);:�[�G2�yf1	�S7.�
V�L��nh�Z��Fʥ��K˨�����ʖ�J�J�b�g4ҡ;v�:L��8�2�Q����.Kb�ѫˢ��!�T�h[�i�3V
[���{L�D��6k�a*Lך����f��0����vi�l���A��Ǹll�²�j鴞GN�lhD�[�c�ɺ�
�phK�71n�6��\�e���Y�w@k���S�D����)hz�����V�NU��!"�mco+��ˣ��ʹ6,�`�w(amD�
Q�E:u6��w�0��F��P�AV[�/HG4���.� ��)�����m��We�Y�tc��̢
�Or��	�y�k67q�ʢ.���Y�Lޖ���Cj;	�I݅����ݠmE��!ט�&�n^ї-��z�-t�1���Wi�kj�:"�%j�M��T�w�8wk`'.�ܱ�X��օ����%��e�K��Bj�&!�u����՚>�+Y;�{�a�`ATڽ{m�e&���p�/rK����i��j��o6��ZRES��;�"�SB
�ʷ�<�V`���9V�u�bv���D�KU)JX�z
˴PDʔvZ��J\ui��e���g���{����]aܧ5����h�a��E��&,%X� �]L�"u�Ӳ��0�1��e��H0�˭���[͋4d�N��ٙ�F��PzJ�ڱf�K4ީ����qD:��cu��6���vG��nʔ�`�e�+/��L����zE!v�O=�krT�'RKW�"(5Sjѡ���@B-�)1R0�;��l�w`ݫM�ϰ�wmr�K���hC��$��U�kU��Wn�*(f=ֈ�nl�Z�^v]*��*h{D5���;4���[�Q�CM>�pLp����.�d����R$l84���O@V�O`�t96�&��)���h�T�U�����v�����V�!%"|��W�]�o2oq���j��W���݆�>ݣkS�֪�1�[{w! fB�A��@�x@x�)J����t�`3�f՘���;��5���i�5��u��Be3{��4�E �:�=���35���壣)������$R�1"kqdT���]�����C�K�v�[z�7�F�PiƱx�� �Kǵ+j����i�t.d��b�kD�����I�`�K!�C��c*�j���vd�ڄ���`$fu�XoX%���D�os	�Ɨv`)��K��X�ެhnn��to2�׎��6SDdu �ͼ1ͭ�¬�4" ��Jh�tR�ۏ( F���O)*w)��7�b/B���%V5f����`��b����i���Y$ۭ���o�Z8��n1��v��7vC#W���F�e5[��������h��L�v��[�e�w��Yt�ɡRf���!�B��O�ޅ�Ӡv�5���[�E�t4,'�k�+[����锈׭���Iu=M�&�(cvT�����@]�{�׳�� ��2]��gv��4Kf�85�bF�8i*�59�۹y��Wb\���M�]�	����LŚ�J떳���l����t��
O
m�l�TQ7+*L�1�a�5�SLi1qY+*�T+1��e���k���Z�̥�i�Z��6��h&���y��ڕ�2�PViD�K��X��5Sp�W�݂.dNSs3ą�[cAX��G0�m"+Umi�,ڎ;�/�j(lZ��%a�r��Z���C%õ���i�;�k%ђ�j�.%��C�
�1�ʵI��l���U��!N�[N��n��NG�f�B{0b��۩xQě���ф0��X���h�N(��l�R^�f�N�e��qn:������̏bnY��f����.�zo^Z�e���sENnָ�R+�KQZwV̭i�����Ⱥl�B/�3	nYi�sÑ�`���k͇4��4�=�
9l�Y.M���Qٲ%�w��{t�lc1��ۼ�m'S1�Hf�q�&�������I��ly[�(f�� h�i�q���6�v+\��J�h��;�5ZL:�����:jn����]�2�=2���e�#tŋ%�O�0���s%���'��ϯq2���S�q�¬�r^�YKP�3�	[��֘wsY;PL�b�eb�I�u��OV� �!CD�@��]ӆF���XN�`r�˽/e��];i���D�k�Y�ؙi"	X�Rw`����YCuA��JX���֜��I.*Ŗ$3 j��o^�ϝ��?M�Q����,�M���z+sY��,�H���I�̙�@�l�8� C�{�	�#�гs�L�Ψ
�W����� ZT�͛Y��=ח�b�2]�o�ef �f]m�tq�S�	�p�����r��f:�\{u�Vf��RO�\Sw*GQ&�Y�{ZE
N�m��9-�M;w��,,r�b�m��l���i���3!�ʼE�d��a�8�n�'���;H�V����,h�QjF
ǫ)[�f�Ѧ�9*T@Mպ���^3D���F<�0���N�~[xv���dM����a���ʁ��Ď��GX�b"4h-��Cfn=��qԼyn��
h���z�m���oR{m�C
����l	�7�R�w�ŪHH�5ф�`z��.����������VA��mUCN�ѥL��e���v_6ѺX������z;N[H=4˛��Ջi�BZ-n�%։)����&��3^n��,�u��q��+M�3Cٹ�����]0Vy��d�`էtT��fX.�積�r�
�V�y�i��/6�<�kh�ۻ�Q&c���c�&G�IYv���s���熚;�4 �t~\]G2��Ъ����|��!P�f�d��Y2�mݜ=#��D`U�Z���E��A0^�������a��W0%�;���W�:	-У@��S5��52��pIɡ�K1N�xdC�z�6�Xy���<�$��*p
�G,��Vu�f�����"G�'.�XX��[yM���g6���B��F��q��$�A�8v��j7�,�� &#Q��ө=�7F.���0�]��>��b̄{f��D�u�h�2U��+>�b@ɔ�)5�Y5u� �1,�*���ߝ����?{��}����������<����~���7~q¢e�P����}��:�}��2�ک�Ռ9�$� �p���y �'�j:�,��u;�v&�0���]�l ���i/��ob!�
c�.���N���K�a�iu��wQW0}���u��Q��g �lm�u��2����R�m,�f�{��W[�h��\6Yyǌ��>��30��]�ox\��o��x�����@V�ޔ].��L�O��i�z����鶪M��{�ʧ[��"���<B�� ^}�r��!�`x��w���zk��	V��ۤ&��NI�p��gۻ��ĵ{�hl)%pӊ�</F��Z`�; I��h�.��L%Р�U�;t�8U������="��2�V���i?�!A�qh.f��+t�e�Z�Lr7�Ԕ0o_l�T�v� ���+z�{�5�ݺ���\D�5V:]t<�������[{/N�\��q.���Q��u!�n�����z�*��uw�j���FJ{���\���kpl��K=)�@�PśصXE�f�b�Y��b��[6�<�p�ۄ���jKB�g(��4x���P����T����zС�zS0��d]�]Kr��;w���{)ƽs���ʠ�6+w��p��k#��iAeNS5��q�]��ϺLZ�t�$�,(�M�[IoS�2V:0�����!�]������p5Vѕ�پ���Os��6��H}ǡh��(0n�f�Hv ��v&�s�{t(���E����m���fc��nkUgP|[�aʓ����M9j��*�Ynf�p������}����ܡ+Wn헸��)�.��F5-�ha��ꥄ�m�
��tMXB$�X�u.)a����]����v���-�tvU���1S�6jX���t��@��+t\��"זDS��[ٗ�T�GU�=+���E��G��m�L���7:3gV��l���{og;��z>R�&!�4��cb�t{Yp�T�A��cU���W]���9���6��J�����Ӈvd���䢃x�m4���va�Jf+ڷO$á�p�ɮ�����
�	w�N��r-�w0� �u՘Yss�֝iǵ�+��%d����7�\�O.s��:!`�� ��Nܫ��h6��ն̸0����27�pwW��i�LgN���ĩu�$�\(�k��n	��s(2�>V�[E��8��(fu���V�'�ͽa�z��g��Qs���7�ln_Z�˷@n��&��o�V�CF��Iͭ���������cT��գl�xT�`[��4��3��7����5hH5ßt	u��)�Nu�kd�����9_��;*�D��n��_�%�z�I��"凰50j36����z�^b�ܭ�:^ھ�C���:�
E�i㊻�/���##�!�*'P��b�%9�d�G��̽��d�u�Sx�sz.�V�:v��S��m�
�}Qķ~���K�q�x?x}�+f��6��kǔ�Z�.��&&��K �5��|_��óS���G�n jR�1I��r�ǃ���][�ZC��)Na��r�������!�ڋ}%�(�ێ E�3p��*-���
���"���;g�M}�7n�JX�PYݢs`���X�H�N;�X|��X�mvb�)d�ܤR:�|��%iލĻ�����YH���� �|�u���}!�6u�� ���`Ǻ����HI�Fsy=+'5Wy����F^R.)�!�|�q�z���������C7h�Yƥ,_
�&�������W���A�+F�P�$����t����O
� [9F�ʏ�t��x�L���I_m�]3O<��Ss��-7�Y�.T1�hoV�X{�{�1�Ǵ����T��f��$�ү % ��K�j�R���RӼ�Д�y��ϭs��� �h����υ�0*-����F��=A'M�Ӯzd� �];8�+����a��\)�c��"��m������V�qa�8�� �T^�-�l��l����:+J=�,��
� L���l���f8v�5������g�����4��|)�K
�\��ăFG��Vt������ڟ]��oz�,V'� �b�y�skz�vԇ*���^b�����çA]l�gW_&)�T'W:���ѐ�' ���rK�6�.=���o앖�^f5 �NՊ��#��q�j��&�W�Y�#EMƝ�ΥO^ձ���rS
8��>R�a��e3�i���f��NsU%�[�dƵ�I�j�9��B�x��Q��af:�.v_��V��D$dg���ժ�������;[�vQ�ՙLTg##�9�YX��\��I�r�������wgI�&�-��C
%�J�i��F�7��΋�^����Y�fn�V�S�m/^�u�]E#�1�t6*oF����h^';ZJ=k�oi�B����,+��z:#j7F�"n�#R\u&�(;����w%��+��˼�$q����T�@�F)Lu�D�VGG�]�(�Wo�q��.���w:fKj�hu����v��>͔��`�չ�\7����P֯�]��Ӎe���/�������%�L�SK�Щ|t��:(=�f�c���FJ�7(�N�;�tPBt氬��1s�H�w���`���zXA<۳�c��n���\M�i��F�aOa����F-ټ�5��Ff��9�����Z<�����L�l�N�GFL�a�n���4,�޾3�H��^�P�N�z�p��Xnh(f��WN��+�ƛyQ]`���mҮ.�os������m5�"֞w;�%�zB������ ��U�vI��0[��u֖�u|[&�����=	��H�Y�M��afV�gE�Ū��Qk,%v��kIM��/8u`Ȝ�\ s���6+�ҭ_Ff��n�t���K1Y��a��p�Z��Ve�D��6�ы����ʝs�^��|���Ra�]}��ٝo.57z �.�`;�5�g��s��2�z��n�WJ�zVu��5&�]t����*Xڊs2T�IxP@3W�Ղu���C���� /z\�P��9�;(����)�L�˵O��7��l8��북��N�L�q�/y��.�d3���*��C�Zq�!����%G27��xh�Y�M�A��og*� �<��y��؍=:U���7�Ԕ���N8p�V����
����q�\?U�tMq�sL�z�FmH�0���6q�.��|�\#�u�H�oL�Hov��uMP��ҳ�6)�sS¡�cB]4=μD�]:y8����wU�]�#:^w<1�,���7�7Jt39n�#��rF,!"=|�6-M�K�P�VQ0m2�9J�_nX�F�cS�O���rfy>� ��c����t��%u�kȇ�]��I�B=�}/�H�S�k�;��ݹ�̧���nd�۔Q��wJ����wbVE	���Vn�j+EIX���8�&$	$�=�S5q�Or�W�Y�n
͕�"��6ޚ9�wHc�--���v���z���z�:a�H���P�):&��ʉ<�{D����[��Y�S���3���l�������'��NI�y��Iٌ�3��0�D� �Ȫ�%����.�+{�)��2_����o/P�oNE[l��f�9�&��jb"�S9�N]��jA��a@pr�����7CL���}�S��Q�m���JMZJ� �Eja��@f�]�r������	R�Hx������{eR�cwg� s0�4��]W��A�ƋyJ=���[��)�`�/4&�C.m��d2����杙��y<���
��8�S�����[s���L"��!���ڻ��q4�*��ӓκ��:G��6Pv��'��6���dI�7�3���=Z�s��X5=�ZAR������@9ݥ���bm她�qm�Ͷ��˭t�}�y���N���mӮӕ��=���N��Y��X��N��@v���8�|����+]GӅus�o-W&G4���j����P�γZmm��4�oXr�!/���y�9j4�K�C�ۊ7Y�u��N���	���������|�=����!�N �N�׀(l4&�P<ܾ�Co]�b�R��1�.*:U�iK=�Ŝ�V�@��F�ޤ8���\z�n1�]����f�+#e�"��R�e"�L�\t+�S	V�y#�#6���iv�qa�z�K�@�z��;Jo8�V��sa�9d���\��Н,{W�rG��X�R��T碲����٘�aS���]�ܾ ��_:�&9�R쭚��w�FGzBҌg��j��ݏ5� ���H ��Y�r򤗇�$Nt;M��:G9���#�-������T�v�<�΁θ��[v�F�>GE�]n:*���v�AsB����vV����\�U���MְwG�`5*�nx�7�y�/e-�=�X�[h��Q'7(�{���(lPq�6�\��S����n��<ʘ%2�'Q�m`����'�2]�U��IJd��9�ֈ/��j�wM���bU�싪)�)KW+�����	;��@YO���J�������x��}�0���]Ҭv�o�������8@���%����,���&��U4�sȔAVS�z��
�tqT/�
-���Rൽy-�L��\q� M�wu����H�ٔ�n����S^k�9oLR��c:ͦ���-^�l��BT���[���֥2 ��}�v��5v��ed'Z�l&����%k��a�i�Wb�ʔ�k���s˩۲����{�G�0G �U��O&,H��]�N\��[�i���KI>����wI�s취��|�"U�`֮y),Ž�F�A�Ge��E�D�r�w��y�8�ubScj�N݊n�S:�t4v8�9n���J����Ыc��I�ˌ���Fὠy��}�~���C����1�N^Y��n�/T�!.�oUP�WK�֞�O�Ai5t�'et5*H�u`�ĪDQ�]�A�kpqÑ�ܔ� V���ܳw��E&�
)r\���L��3m�N;Cv�'I�����*�-�;��3t12��s�3ld�rm�2���íM#E�3��q�++��	�r[F��t��5R�q�u%k&"�����D8�s�����l=��p���	."��Ü��UU�vJޅ�<%=�Cr�v6LOeEˎҥtn��� �	��Y��@T�U$���Ӷ�t�-���*��\�șݚV�� v�h�� y��C���zOay�݈�]M�kB����Ѿj����QQ=^[2��X1vKi)�v6��2�cx�;7X�<���颕eQ
�2�gHåU����]E\s�V�W�a�����U9��(�k�����ʂ���Q�γC9�jl�x�t �;��d��S�KL�+N&5Die��B��v��,Ty���{��-�a���J�*�h꒎$����V􋸀ٷ{�$ѩ�Y��r�M'���Μf,+Z�-��j�N�L�u&ꢪ]�*�3{�˻>0κ���5( ]�瞮Sd�5���>�1�Z�l)�{����p7�!�6�i���q��:�
,]���;�׉N1�I��wӨ��d=�n��>�:�wgK9]3��;[�;�	��Up�-��ƛ�m�8�F����&�fS�bn�,�ªٴm�b7���ȸt��6>�2�i�NQk��t,R�k����D�e�w�f�Jd�����R�[u"�"N���\��O:ˠ��+�8���g(k.��8^�p�,������Z����y�|���Hs�.��uU��M&$��*N�sU��`�y#t�h"��V�22����l[װ������Sj`�N�G¹9[�V��#)k"�i*.e�2��s���ۆ�ؔ^}S4� ��N���Ŧ��E��ͺ��6oFYېb*��`�͏5h]s[���[��F�\*h�g��c�r;�FN��z`�����7��yet5��.��r��t���M4ӟN��l2��F8Ģշ�Wy�y-��CSo��͕3��<s�ue`�}>.�b���$�S���Z�����D��~�����f�zD))�m���d���<�u�!O�Wa׸��S���^���J��	�һ<�$�t
�6�G����X��nsU2h�`�*i�5���'o�3yg�S+��X�t˹R���0kk�i��6��a`��Z/#յd��f��Άbi�7tiYl{�M�����˽�9W.�{BN7Ƿ�J��8P�U8M�Y��wh�!�zN�{+;��8n�e�7��՞��D尶����.T�m�n�_!�_l����|��З�����:7{mż}�v��ޱ��Q�H�Z��z�I�%2w+����".f�n�����m��3)��"�[sc�ֶ�S]��Ж�8�o�Sy"YC�8X�B=�y2�9x��4�����K����(Y��vj� a�x�.y��YBB�}�rĖ��v�k�<�亶#%���J��|�X��(�GRq`"Mʺ��MSjё24۪"�	�f��3��)	Iw87nV�8wrjU4���������ֳ����5���ř
����&
K:�5�j��"��Y�����{�L��e�n���B�6*��x����*��������#�/%ڍ�m�L	n�]
vx��V�k��fk�D�O;���Ty^K�.�Ft��W8��4{�����9LeiW"�S.e�L=�v3;��ܝ�ݒ��2>ٶ�`L��+u)����9$�H�I$�I3g)$�c�H��'0�ʙ��U�V���J��Vt|�װU>5\=����kET��*�Zױl�Mv�� �U��&��''�u�9��))<G�z��Uh���lUk5�)���Xm!�.%���Xk�<�lנ�+,�|f9�x���sz�������QQ~�S��B���q};���w��P@��/�;����}>��}Ŷ�^/���5{��2�#`��yP;����	@��g��������E��k��x��Hr�t�*,�v��<e̥�[��%:]F*����:�f����lh��U�fڄT��������O8�UjT{nX��SE�𮵉o�!hs�|v���I���i�sj�b"\h��QYg��jU��i�w&>Y�.C5꘢f_K���9�:oM6�5�n�3�yJ3#6/\���Fv%��e�{z����qNm�����à&�a��D��S�
)`���쳦��O�.�T)��\:���&ImbR�;�}5IҐo����yk��|��W��ݜW2e��A�hn<�V�۶;n�	��*��Q|��2�Wlt���h�J�Aոs0�P��"�]e��Jl�F�Cr,�S�VU���-L�C �6��p<���HLJ�d+�Z�������.A�����$Еf 5r@��Yp��h�D��a�ނ��z5�j�PA�]�2El���t�oxo&��^R�[Cdxn^��G\����^3بƶ�Q�ڃ0R3*��v�C ��:Ű�ۃ���j:��hW�OW!xN
��1������V�BÝ)�<Zԯsj����4e�x�$�g/�8:�7�(b̙:1��R�,�	� �\c�Q���f�Vwfl�̘R��P	ۈuݭ`b�˨-VQX��<�Shr�{˟0C��¯dѼ�ɤf��a5f�"lp�ƨ�kv�x�ȘH����1p;#j��H����*V\��*-d�fX�,����6v�q͒F�^+L��p�0wyb�tX��I�:�A�s3:B��ʛ kP/�тr��!��2�4GR*v�O�}�q�;��ʗ��G���#7SA��]��&����u�{�+,��Ipp�U�ύ �t�䭘�x���K(82�i�i� �*\��
dY�C�E$��nk��"^dfե\W�{�>.*�]�:�[��:�����u���)���)�����Z��+5M.X�����BX�qoDm�y����*��@l�O.�m�7�58�D�O��n����f����
�.|l���kV+����aDYg����+g
4���J�6�U�9�M�@I.�����{�|�Ӧ�[Φ��)Y���;��{Ev:�[�ɽ
��װe��:��p�k����5�e>:Ht�=���ڴ��Bm�j=���L�51�B�2����[S�ڼ�۠�.�̃�Òd7C�ڽ�Zn.�;]��3\�Qų�I��ӽ���6cF����R��飘G��f�yPo�,�J]�֣����W��!)K%�(�%PN��cf�K5�¾����m�Q�׻w��[�iT���k��r]f���ơYB4�J�8�iY%��۩�WSMYX�H���V�7i��W�v�=Ճ�Kvږ"uЇ�T�\ �.���6��*�[�C�Seb���Y[Rݛ%��91z���@�2�va�޵�Ѳ��^�j�"�����:�ڎ��8��B��v"�L��ݫ$��] ���z���Gr]dB����﹆қ4��a���-�a$Fi-6�6�4�8Q��D���#yc*��Mj)�HmGt��0�Y�3,M���E���dsu�I�=훢"�>�5��닲�靑R&�"���;-R���h��VG�u,O?Lu���2��n�*�Ӎ����L�LS`�f�d����=
���r���hu\�`�M9� %9|U��������� R�.�v��$�5�]�`]�^����η"��N�K�[��p_YC."��o�ae�E[�g�����4�����ڼ��(���S_(�Ljn���^�(4Ck��JB�{5*�w}�k4˄�6h1׺���5������fK�Sl�f潠��JWn�N�U�U�:*8 �:u�|�o3@9�Ӵ�N��������.�%Y��3xe������:�`MLķW��[լ���W�c�i�F_l���"�A<g��UԱ�;9Ң!ƥ������̶�*	��"t�oY.�e$��yw�PCz��zHX�I@��[e��y��T3�O�U�әB�f't)���yepC�ʥ�c�8]����x���p���j�U�s�<3iK5�]>��6��E8Q�i���b�Y5Muw�S/cT�-���OWWq�,�W]�6æ��r���8�v�oL�g�TYig׳��o@��]�J3��V�3�e���bo��"y��U�S��8;����*��ٔ;���^�I�L��R�5i"��C� M�(ѭb���Q��jBs8Ĩ�<.̩|,���%M�.w�:�|h��U����%P�Tt���w[��Ƿ"Sln���6v�Hf��o�G��/)��i!P�{.����}�:�4��OV�<t�6�i�8V��"Ň'i��7Q������̿�޳tݚ-m�O<	�ՙ�Z�*��{�N�+_\׼x�k��We:�U��n:ޅ�H�㕒�#v��1�iz�{�_F���uH'ʂ�.9������Qop�]�	����(��8�,�j�������qe1
�Cu�[��L)��r�w ��o)�Z�F%��Y�'�c�b�Q�@4�s}��QI^^)}g��`�X����JԬjz��H�ҹo^��u�u�=�
�-gJ[�.�`=�5��
A����v��,�E�ͤ��+��;wT��4�j��қ�Iw����o���҂p��]��а9�:��L���s[�*s����hFK�$M.��(��%ك\�<w�Z��k��y=�%��5��6��ýMԦ	i�K^�w/�2t��u.a�A�rYu����̨���xq��* k��U�j�[e�=�M3D:�(�QOZ�mQ>b�Н������;�2��`��*��s:Df;u����MN8�]��nIi�3j㹡�]�63���p���q7��p�i��Sn�%���E;��WX�[:P6��z�������G�lR���-�p�Y�e�D�QŠ�
�#�cuyG[
ҩ-FY��\�1(��]��Bj� ��.ZO��J�ٶ��S�W�P���%��(♎ڨ�7�{X���tb8�j}��d"�/��u�ft�YօН�k�)�]�Q�必k����S����Q�꺴b4�<�t�<d(pLwo*��Z[��J ���@G�bQ�df�<���N���N'sK:K��Ĥ���f\���`Y��n�|
ڗ[cf(�Yz�n�P�o
��Li�����uL�w�a͗V[��q�y��I�ܶ�P8;�
�s�Sژ,],˩�D�k��JsS�����<�}�E��{B=�\��t���hѼݼ���|��s��f#��ݮq�d��S k�k�k�m�TW�t���gj7�Ǚj�5�e��]	�0�����u�u|��̻o�f��u�]M��z$Y]��;=�㳹C@fKt�Z�NN[�
}�4��KXg鹱u��z ��P�E�-�ZGG|�f���4�Rvܮ =�om�A�������I�w\�uMl4���V�V=�&m��HjU�DM����n�>��5�����
��]�ŋ���G3r��(��J�MY��
�)��=
�ʴj�;�)z���jˁ�۬Nd�ݔ�O$;�;A����a�!��Z�i�l�n�����J�M�f[M��)ݾ鄍=-+3�״+UQ�V!I�8��ȡRY��].^�Ǡܡ2sx����ov�յu$|��gZ��Jv����L^ް���ŗ��w �V�8\�cj�Ӭ#{�lJ�[ Y�O֥�\Vb%��:�ri�9�U��=�� ��	U�7����v��dt�3C-��z����6�����҃j�˄U�΍.]��fa�91a�3	�t����F��,7�z/'n ��F�dݺ��z��HVC,�ù6�P����@Zx{J)�[P������lsd�9�X���e���I�!��ʟn�ԁ��N�5�o�o�صV��\v��Yshuwp5��=id����̬�!o�P�No���_���hv����JCo���h�ns�Ζ�����׮��t��Ԑ��_w����ب^#V�����Di.���U���ePF��,]aK����_l�T����cL6+/��α
<R $0�.t�!��U�h;��y8������
�E/��[.;rY��=>���#pJ���ݜ�7��(��m�;Z܂�r1�����{�%]Vfu�m��hX{�n�*�6˂��%f�`�:'f�`x�7/��6>�� ��B�۫�K���T�r����əuzP��ާ)���hwHb�1�X���{�^�Z 8R�J����5�e�r���4\�.g���W��^�P�&�9�/!ק����tʍ�(��Ӗ8�_R�ku�_�V��g0�{FS"MV����N�b��^�1��r�� ˰�\2��s����6�虘��;�bX��+����\bGl�鵂��9��Y]Av���)���	n'��Iًt�J��ގm�Q)B��w*����<�pJd���  �t����y�F���90sL��y��4T���L�"�5�w�ا��v_�p�ɕ���ܔ��Bw��|&,�}�M��ꝰ`͒�;�N۸��<Yy9l���ﭻH������0jD:d�1��H��φ�y�jv���w���m�6���)Vm	�k��E���j>��qM�����ַ��'l,N��%�*Us�X�7�]�8�)+�F�*PW���o	�n�Ý���nc��o1
�Rd �[���{
��+�Zç���x�PԺ�Z��N�Y������ŇgHz�x�.��vf��n��k�u�`I ���U��x+�J.ԃHnt�QU:wT��P��om��6;��L�J�7C{�dv�\�C�[V�b����lnuFKr�j�:��\ҕ�&#xH�3`+K coFk�KE8�=4i�Vwk�����~�f�v
�Lw@+4s�&�֥K�a�.w�)��vҞz`�����H��-F��֘�ck@�s0��0��v;�Y0H�.7!݉��g}��L�F�X�W�.�;�B�k�2���c�3bt�M��Qm���v5�=㕅;=��A�t(^�\���D%�)�K|iV��ӵ�+��yj��d%Z��gD�8;ѓU<<+����rŒ��*lAQ�̒Q=`g�u���5k�մ�>o*�)��T-+?nP��)	ܚ���:]�Pdl)��2����N�u7�����/m]ӋH�i�W�t'NI���������M�}|1��f�NĠ�p�ɏ^�^�d�|�/k�NW-,���l�U3�a�p�Ip�8gS��np8 ���R�f�X�}akgV�݅րo��N��;��:���2��5��]J:�,��V�'y%�ӌ�L�Ǌ"��y�h����/I`���0+�Ǐm-�hu=Y�y[�V��'3�2�b@��n��)P{���̜�i���N��bvMq����z��hǻ��Y:��	��r]��B��vm#6���\�cij��iȺ^�o-�m��ʯp$�e�/.����2�:3n�Ss��v�ó��f�G����B��7U�x��ko8b�W-�+oV��0��/.��}��0�f�Ѳ��nP��汚�xv��	S*7��c��e\��P�d�:��+0�4�^�mv��0���X�!�G@��XM��r�Ph�-����t�����-< �:6r�ؙ�>��ݮ�9�5Vq�-���b��O���n��ݍ��(��TFL}��S���"�u��y��خ�!t��7	DS�)��t�,����Z鄦@�K�t^�z\���Y�z)%[x:���L����L!Bn��,r��]�L%A�]�[��Δ���Sڲ��3�=f-�[b���w���ޝ�Z���=�6�Mx��'5���T���T�2	�,�O7���ؒ��ٗcPo� p0b��u�i�X���� 4�ows�$�)vSʹ�l7�0��9T7����M��
�BEݻy����i�=؄<����3�FN<��Z��k�b��h<Yy�3�Jfs�F-�ʻ0rCs]s�#H�ƫ���Μ{"���+K�WݩP�eC��L���:MU����F1�*a�����n�YX&Y�.����]�S�>xsU��L �ͭ���p���ɮ����9�q�भ�y�w�@�XԺJ����c>���j���]&�Z���p\.MQ!b=���mluzUtv�Zא+���5�.�7}Q�^lwf��J����W�+��|jJ�Ua���F���������q4 �0v^�Cx�:m�o�l�Y6�����1k��	�[Γ��X���"��n2ƺàEl=�V)�i-��
�fA��H1טV3����w�ۚ�xͱ/r	Xކޛ�:۫LKn=�����m��M�ա%�;Q�\�9W���!ybrR�Lf��Ԛ{zݺ�t��}���5%�B�'mAWM����B:�3�X����;ٗ/a�E�7�tڑ�me�C3�OP��̘2�,�\r��A���٢y��c}���k���&<���.g}���t�Pdpts��a�je����o���آ���N]��"'3�bydQ���}̮�D��tZ����5���%3,�b�+oj��}t�Q��mͤ�Po�N�t��&���q*zk��{�W�.R�'.�+̲�B#*�����;��$��g�RTWS�zVSЈ���-��	7�ܬ@�}F��huY�̻�A����l1P�Xe,�˂�����f勡�-�ݙo�t��B��KH��Ҷ��@X�+P���5U�[r�`�q��QJL�٘�?��k���Q_�F�_����?ҿd���_��_��_���}>�O���?�?����5��v�=�^j�Zۜ�4�T��P��2L���9dR�a��Mh�J����	�U!H���o������A�-��q�y4�Gr̾kvA;�ιX��
Ue'Eɓ�����G{����]���m�[C5T��(h��Y��>�^ɔ�,����Sh���g��٢D��A<+8m����)�p2b��x���o��5[��%��^�Nv�}�>ə��2�-��6���M���tm�*�+mm̫9�s3r�ڪ�ԓslnY��w/WR|6wG�,b���W��;�$�b3R5�<{��T���f����C�@)��B����@B�&�� �W&��L��\e�w5/0f�u�U����W��`3Mr:B�e��K���vںs�qm��pv���h�v�s�=�]g	:�t��¶�pf!��U��֎u8X
��w!.�m8����7��yn�P9"�����u�i�m��p��[8���5X��Z�X�N���C6��{��c���܅�r`L�rc�Z�%�9Z�"^mJԊ�O�)��fGu�\y�7���خ����X��1mJ3����xeX�@��`5�1�+��Z�3�6�θ�L��lG2Z�����/�ʾ���Vޞ�)�t.�o�J�B�7ف�g^N��`ʮ��CҘ�vﻃ�����{�Y1�j�3��6��Ρ��͔��Orv��w7s:��{�srf�:+(*D2Am���4ZC~Ee%EQ)*��Oʨ$l#�I��T (�D�@��� �U
&�a6@H"��XT]hMQ��`��	 �I��e:��:�u\��]o4EQE\ڢ*��"(�����"f���*�j"�� ���(�(���)*�����: ���H���")��"*h��h��ՌQ%5QT�SmMT5MEMUTPSQSI2j�$�

�f�
����"����PĒ�QU%TDPSA%ER�5D�GY5F��&�#s���u��TAQQ%��TTTQ3F�A�b
�`(����j"(���5x�x�\IE4�$�i�m�DTAMQD�EEUS՘���*�������EMW�4�*O�*(
i�H�
�(�&*+IF���*����)��H�B�)�o�T%STUxآ"*h������Յ5hUՀKH+7��cͩw����P���n!�\ϒ�:���K���P�6���Nwz{rܔD� ��Dvn�΄�q�K���@]-D#t�HID JT��
�z):���;^����Sc�c�Rv��H��ZpLYb��~Ït���^=���w�D�i�3Y�r��Ll�r�&̗=s�Y]�3%�Ҙ�;�%�K�/=.���?����(��;_���\x�sƳ�hzj̒f�[}�.z����4��{��%{J��c���բ�A����:w��)���E)�o^U�$*V߼�t����z�=D��]�xZ�9!F)=��c��2ey@�ɕt��W��u��>
��"fz����̥�r���,���ai�'^}F��wp<_�!�cg���y�`�Qy1yOs'�w�g��tΓ��A*��ù��ݮe�WKw]����NcU�K���C׸��vO�'链roN��{�hI� Ԍ�"[���n���``��e����|�Y�HhR���Z�O<���Vߞv��B=�[�����+�S�~PuJ�僺��Q#c�C3}@w��]�_�Ы9`gjf�*�c�S[+��+6����j@���@��L��LJA��qR��vw��=~��M#�N�YmY3M]5J�ʋ'Wɚ��!ShMd��:j�=d�wy�j�TՊlk}��vmY�����ӑ*���'i���wS�UΔ�Y�^�@�ɥH־��$`��f��b(�^�?n�!�w�ꐚ�WH��;�K� ��X6��X��$�3(��;��o��.����S|s�=�����qVmR}�Ǫ��J���7J�_w���wɏɳ\�Q�}{����vk{}��4���I�#�I}���:�����u�٭��$m{��n���i�hH�l�m&��=��cY�$w6��mC���i�&�2b���<7�=�G��/8'�k�����{���~��r:�X�r ���|�v[H-�e�_�����m���;$�7�G�۴G[c��`Ү��������j#��7���lR?h-:���/����������]L{Ջ������Z�u�������I��'��y�;d��y�k���S���R�C�x�C�;���VSX�,���Y���5��m��
����+�a���m
���C
oL�kKx#2�dN��]f>=o'�'WswEිT��.ֺQ�Γ,e)�ӛ}Ξk�bSY���w��ܡ��%�j�fK���0 pR�gىU��f����aTO�&�rF�x��ɡ|h�^@~�?z�p<�����ݘ����	�>���^V��F=��ǵ���ܧ�3�C�<��h�M��FQ�=>���<.���z��ohU��^?m�*��G�Ln@�h�5-u=�t���ѕ��s��#>�L}�r�zk�i���I�謯K��]-�7�_���3�<ҍ}�`s�Q�������;�P]f��&Eu�ʼ�3����Gy�����Ⱦ'��&��|fW�w�mX��iS���Ef=�ʧ��*/P3�E�*��zs8�Jr�q�Y��c#L^wt��K�`�S�L�c���"I���ך�u�';�H&���r��Y����@��_�N������p��D��U�i8H�"��Y�evv�гO��i��3�<��6��r���=��:��	�=ܚ6M{&,�9"��<{��n[����#����XO+`)��4��j�Eb�t�1�G]���U�v��y<i���h�H^�뭃�D�B�d����:�ڨb��U��]X�㧟!{��k�����k����ei��K�ijd�5Z6�WS\ĺiEB��ԨI�M����:��3�{j>���3��{Nѝ���̉��������zF�(��@����ؗ3Mp:kڗuzm�����9u:�\��t�\�bx��Q&��gC�@ۧ1Zw(Ց�����F� dp3��� ��?'���秷�2g�$%bT�G;[\!=�8��omL�x,�NA��:E��-�LP�G�O;Z^��t1��x�i+�$"�[�n�J�"SyT^z	�/�{7�S����κ/1y)e�ة�n�vzL�@�]
}}���י�y�3'��k��7�>q��]��}ۯޙ�o�k<��)cۡK�I��OqYI&�*��v�7�t��o�ɽ�_NVO	�>����ʹ���+�ԅ>��w���x�ǜ��;$n�'�����E�;�b��k�ުv��U���o^����T[8ڨ��s.�Ç]��HXC�x�����
���.�J�t#� .?��z��.���.�T�*���4F�@WVL���67B/Y5i�mj6<-����fuuü������,��	/F��6����;��͎�kҒ�)@@�[�@���z��UA.zU�{i�f.���2���R�^��ܪ�m�z��9\U��ۅ�Ut�}��[ޝM���.�m畅)_�ݎQ���Tk�:2K�Y�ǀL�WTհ��������Ȥr/��\�8�|Ҕ=���6��y�Uɑ�Nge�X�	��>M�̜Rc|��~��d�7���qz���G�}�6�eߓ]1�M*���dk�l�+g�d��S��(חo�w��%yz{��w����[��Z=)�8ݮВ�W75���с�[�'�m�nH���ۯ��W�`>��Oy5�<Q�;�{�	P��
x����p�,?u��z��4��K�{/�{4��k�-~�'��귎I&@m���s#1�����N�o�| Ý~��)Ŋ�Ǳ���b��+�1�7��Y��힖�%�[h;�0p�3L:�h�5E6U���a��7Ks72�䲽�^���Wb�����5�*��ō��ԆS�XTUX���[ лD��R�e�F�d��/�Ӗ'So2�+���C#�x��7�v�������X�m`�V�7-��ԝ�Lo�_{�G|�{��Ͻ�ߟ�zI^p<��n�Eh��^�[��w�JȢ������}AW�g��Ft�79�3��p�y��kʛt���m���įO������ð���α�k�M�ӧ({�nmg��s���*)Hsݮ�~��h���F���pF�Ka��ǹ�f��uy��z9�r�y]�)#�zlC=�qYM�I�s���Z�N�WM�����Gw�,�1�=���#��Nn��S��Hb���ڸY�T�U����K��Y�Ps�j��b���%�^Z�<H��`y�v
Ƈ��Uc��B�Oo�~$v��7P:h�����uכ�//�H��I�0���9~��^�;P���h:�g�7|��D�y�q`��Q�ާ���wL���y�Ѡ�'Hy���}�����C{գGt��b��d�n�9@��c�QɆ��FX�ا��
C����/i�&�o�E-*0���۝;��w��.�Ou)�q��ЩǼ)To���|��5jK�K�y�t�C3v�0q��v����M3�k7Y5Y�uŲ��7FA�*k�K���o%�6�.{��4^���֭�E����R���]M9�k>�m�[���#w�֫P��q=Iz��Ϝ��2����G���䗬y}lU�}��/��b�=��t�M]��������a�W��O�&�>ދ�65������ۣP{k��n��@��dYe�vI6��1���R�ʏ�U��=}��خ�?W���u��A22xl�^ܚŢk��Q�?w�y��|;0f{����~d�;7\�]FG����{���5{���K�T�n��l{�_�����_�3t>}b�&n�"��Qx��fL��n�\���{�ki�)���褋=JI�k�>���[�ۤj�ҙ�NK�SU~����v�;�k�����U\^�q�5�]Lս���v*W�;�b���O=��{�y�4"�쁹ͳ|OQ~�\[�����C�V#�h-~�3V3U�3ps�.�Y��R�V��s)�t{�iں+�����~7�s�LU��I�XL`�������E[#M+u�a0��4�����ʃ�ek씖.�nc����Rn�[3Sa��D0�ī[��1��5{ؒa�nٛh�-�O�+/ʣ4�m�����c�+*��\vb������I�y9<W9�lU* p���&�y]`f�����>b\Y�6vP���]0	�6�k��bdp�bgn���\�����{0����W����~J���푰G�ct}˕d�^W.3�0�8��`����x�^���U��p��R,n����پ3=�וvvh��x�^v�s��l6���������@� ���N.L��Nj۲w��|6�@U>�s�?!*aՕ�����rM�=^$Ѡd�m����H��Ȓx��y
5��'��+��R�,�f߽�;��Zo��~8%`�5Xdұ{���*9����`�\%J�����T}���^��=�����%��e�0�)٩Z�}*,t��֏W���#73��.c4": ��Ϩj�o�����u[��a䥔/*�&K��8�f�K�չD-�t���;ZJ����X�����MuY��N���ٱ��;Q��	�F��C��^1�3L��gf� �4�^=��]ڝ��xH�t���br��uLBJ����.�x��E#`Lu��P	���y��f���>�D|]l
��W�Q����u涐���if�ָ��Th�]V����$�{�ǆ[M����)����l��v6'�)�BS�Mz�?v����=����/��n�=3ϩ�ڹ�ea\|p.y]JAG7���e0���H쑹�"����f���}!nI��W�>��'��6�?vն.H,���lI�������w�`�����ȡw$���o�"��~��c�G��*�J�?��n�quu(ɑ����v�wh���$G��h�_���=Y\�z�*2{͑X�k��G7w�����`��.�(=�=S���IF���L��<���B�K�S\Ɠ9�0�_mV�{�=ꉹ뇣���a�Ga=��V*%�z��eI���-Bu�7w�u�jQ���{,�1�5��x�6dנ�Sy�ēOu㑔Gdy�,m����;�d�5*��n�T�zGc��+j�n�(<8��f�����k�=z�c��7<X\�P�G4���C�0�T'A4�uN������S��p�֕@�vBE@�{f��<wBE��Q,#gs���o�[��.8�Y�p�T�������m���p��4�<`�N�cû�/���G�5�U���33!�U��HyǗ_
�ծ8M4�EUI�y�N6���/�Hm��a�zA$�ml�S��UuA�l[���X�B��=omI7�p͞�\GYj0N��Ƽ�<����z{�qg",ď��4����'�&&�ײx�Ɜ��5�^E;C�t���Ի�Ƒ�Z���8�O��Yꫯq��Y��Ft��;u�A�����y��^y�t�L͇�}�xf�&t�*�ׄS��k�a��h$�4���uT�]���Y8d������}����;^�P[�mf���=�9�=�gԽiy�ǽ4)�}�{+�/>��dڹ+*�K����m~v�n��nx2�Q��{.'�+���7G	�m����w��t3�_E����{�W��������=��g���x�#��[Z����K�V����UC{�8��[
�A �u��=����8l�.��k�I��1d�jVr�@Y/�ܬ�bn�h�2ųt�u�Wz %ٓ�kAN��5��x��WVs��v���5�k��s�u��5�4�X�<��d��I15Ĝ��P��� �i�g�mL�c�jSc1��)9���9�\
�����/�!-�J�>��ky[�d4(�*�졻h)�s�����#H)�A�[)Yd�vH�R ���b�XѰ#ݜ���R#Z'�b�9X��A���ǻ�����k;����0V�m��]u��R�+_-R�ͫ�:Y�yպ �oEs.��*o����+���Yx�厦Ԝ	�Ud-M[�y]5.���ҙL$��c;'�3{]����.E)�b��w9GEzV&U�Zn�i��@8���i>О>A#wh�	����B��u�)�ZA��a[9̣Z;2'#�����9:rEη)u�gX i��zҙŜ`9��n�|um{9c.�av��P�!��Sr�RܵY���P���El�9�Or��=�z�\��q��=]�b��c~/�����]1�4[���EY������a޾c]rA/3L��X筁KD�<� �*<Qvh�hJ8�!v{�΢�HѮ��{�Zv�V��Ӳ��˨Q��������\<]�+!<�ƌB���+*o�H��a9Ӏ��qR��+mR,�#|��	}Q�1�-��K��^vq�Zٝ�-��/�U�OI��f�L�U���_�)ĩ�����X�%m)�~Oea���C�d�1�s=l����u�Z�G�']��c��c]�o��C/�.��C�X�i8�Cf�����l�b��=��oM��τg�y;��������g	��H��KE���Kv�`�Z�U�e	�u�S��au�J�t/�5�Qk
��Zy�����U��;m,�p,pEN��𭼜
 �����1�l��wÁ�A��1�~Y�
].xŅ�����ú�]o/D|��]���A��{�ᒰ@��P3һ]��ͼ;]f�M�]��G�(�}��XS.�女,⌲y�h���z"�.r�0N�u����`��W�'P�bS��	J��1r{8�*j;�V�؋*�c<��2���qg\��z���g,��X���-Y\��՞�N.��m�[�7Æ�S��!�,XAbX`Ǎ�^�Xi��u�g�t\�c;1�9�fg��Z$0����_5��@�@����U��h3�Z��FM�MR�X�a�p�89o�"��j5e	l<�\�n��ҥiH*ݙ�����'\�����l��^�1��� ���G/+�W�vp=i2;0�w]Mf�����k
*FM�����c�g�@8��6C;���6.�V[��V2�M��fӉ�r��Ί9��7Ri5�˺V�p��׍����[���b)�f
�*�i=�Du8����H���j9wÜQQU�*���z�
�5DAQULTZu0[8���5�b�cMQ4QT��
h(����wj����T�6妚9:�y���C��5�ɤ�����RRRI��4�SUAO"���j��mQ%DM/-4U\Ƃ����d��+�Ӷ�E��MEm��:"`�[b�yP�iڜkj�馜Z���j����cy��mW��ͪ������Q��[���mcE��F�͹j)l[r0r�u��TPr�D���<�pɭQ�9k�sm�:Ѩ�˫d�b.cF��	w3ˑ����bMiH�#$c`�i����@QA��颩��jM��4�"�MA���Ar)��{�4�UH{�����6���)��b�VQq�G��&���Xj��u��Z�ml�;��f���e*��ݽ�ET$2kz42�AO2���*�_�����w�룫zF��'c���o��
]�
ޠ�h���R291k�Ȋ��蒏�3#��)K�uV�祡�:O��z��ǵ�z��͛&Y�k����P�?Cx��U��ն����.��zY�vry�<��֖�&���8*��o{m�rT��aM�1�`'���9Z�껗Q[ӻۈ:Jq=z��]"��`qmÒ�"��V0J��z[�;����5S����MZ������pj=�sM^�ψ��f��0-U��^�$�p�#,D����!��u�.ѣw{z�9˓��� ��^'�Q�er�#ie�>j��Ҵ��ܣQ>?uܨ�P:T���W���#{�aHЅ�֚Q�'��%9�.�LRR������͏P�@���%wDN�J���L��
�m�W���C+ږ`�B��J�v/)�ց%�[Ø��p,�Pa�����b�ں\0��9A�S��y�9m����C:q���
�`,�n��r�O֓�%��vd)m�����OT��޷C�mz���4 �~��x+st9��E��KƵ��"�~�_�V�(����P�ׇ���t���ۧ��b'ו��f�'E�eAgh=JnZ������pUmU�_�U��gR��. AV�L�7�i�Z�7v��qh����.L�a4�A��.���;|�a)3>@7��˼y���հ������^�ņR�_i�+��� �r�A�ؔ� ���@���?��\�+dS ޮ���uFb�Wé��4��<��GSɨ����l����  ��C��mi����r�k.9��lCR[��}at�LcY7��ܺ}[f���������Cs;z����L���!��?�� �X�0����A���I86��0E4��,'᎘�
ɽ���vs*ٹ�Y=��j�t�k;E�	�&9������6�ÝBhq�.��]�q~w�~����9���M��K����u�~�V_�� ��sH0����m�8=���]c/!�'��k��4�.h������e�b2}��J3���/j�5O�]�)� �`L�#C�z-�p,	��Wf�� ��4�Mt�����5�{ںÅ�475$}��1�����T2��{=+B���-<��=0M��3��19����#n���]QXզN5��׭@�4��z1���/P��� �czuv�a����oSJ��OH[��p���.�d��ڒ\��ُ�#�Z�B��&�~ѷ>������^6��+ˁ��)"]��~5�	�ڢH��|��y���K�FϮdފ�L�S��Qྣ,���J����Qb�f7Dh�}ީW��ER��%�o_ob����9�<P�wܭ��mu����M7D컉{ڱە3��M�����sm䴛��32�[�Mh���ʹe�_���p�_J`9��$�ħ6-'
�,UW�P1���vɩ��j�����S۶i��\[B��a�>3�Aƍ�!�_K1"�˴�z�&X�b�M�락S}�v�ގ��p�\���˞ ��@ߠ�����tW�D��kH�!9�I��ʬ�vo�:u]�zM���Wvq؇���D��ٳ��J�ƤenM5A&@@5? ��;��[U���Z~�|2�׶�	��p=���v�
�Z��V�@E�z4���A(H�伈>9��ş�nm�9������9�[��n�Bz ��$���<fo]���­t�)�U�%=�}4ՠ�� GQu����%����cfBv�1b�Bn�'�snr�K��X�t,~ �%���P���#���Fd�)y� �U���rǵ�(�#�W�'�K8lNw�R�oi�,9�
T��{a�q��s��S�j�����ydj�V
���0���R��N��J<�X�n��E�6��n�Es�AۮZ4�c}��f� g��fQ�
��8V��< `L���C�|`�P2/���Ό���w?����Z}#�ԯm��ҳ���i[�TŌ�J��5�S`Ҭ>��4�k(f���(\k�]x8YP@�m�lk�fpe�V�N��TO:� �ݼN�R�,��hJ60�z��+#��bo)iq�������y����b��P�Yf�f��hwH���P��F]��-��6��\3x	�"˷�e��[c��U0d��W�gM\>,�Bj-=�����t��p9'*�&�j&���.���p�v�r��Y�V�ƙ��Ȝ;5�\�`�>s���/�Q�m�*���_��A�,�m*<��zq� �!���,�m����;�ǡ�(�v� ���0L�q�+g+��KsP�"Sm�!2�iP���\<�r�B��l��G���~�����h�v� b�S�!�R��x����nj~BS&�O��R��4��ܢb���C=�B�= {ʄ��S���)w�:A�Lоou̕��Z$<Ի�M;\�s�yz��k�Q,���n�b��Ã�_?�]D'�k�H.͗�.p*�_T���X���Me>����eA��5{Z��\Fv���O2���q�����6�L|�1��ͥ���DU#�L��0Bm��	�a��xi;��eWC�zN�ѧy��e����uNR<%��e�[}(9L#�`�&֑#X�ħ[&q�l&�W=���s7�T;���Ճp�����	�z�<ܛ�.�ݸ���'3u����V�;ْ���弧�������M�ntk��(�l�uٱ'����l���ਫ^�ݬ���������4<��ۚ()�7�̘뚲����Z�cU���\�f������-�1ݦ{>������X^x���"%���PL��C��؝NM��M�b�a\�V��V���;�Kdv���t��N���r�q＄:r(�����&��d"�W��͞?k�X5����9��\Of��>X�>�z&g��d����`����% ��Q�;P����P���mц�Ĕ��#���ს<����+�E��Ǥ��-������ų�b v2:%�-�k�m�Ԉ�d���<k�es�{�D�4�mcޖ�a ��S@Byv-��ױ��Ű�g[D�C�z�23�5K��G4��&L�l��=[���76l�f��é,��r��r��s��F8�Y���:y��Z�H?�J\�_�<�e���^|n����rT��aM赧Z�����k���L,��PT=��^2~���RQ��B�XH��ǧ�U�����%��Z6��ṣv�f�h���=���=������/��ҍTm.��"H�T��~`SFv�M���[�]���=�D��栜h�(=ɍ�=s�@q��՟5er�Jґ�x������U�]3�aC)Dʟ�=�/C��r�de�B�s���u�ݭ%Z�Z�;��8���j�x��5�o�����=�<�̝�&�&vؚ�+�)E���t�m�-۔�s�!ymtQ��QQ;rLf�i��y;X�`�$5:`|'=�C2��b������3z��S�2N;5|��ވ�#o���DJt���r�<%��%����y�>E���y�X�+b.p������|�t3[H�e��ڒVf
A�P�Gu*I���)9Y�"�-�Ø�Z��U���}�k�����ʈ�}���x�L0^yϯ�z�'zQ����>U�����L_�-��:VWc��z�u!��n�x �i�H=!�C�|�G3�s�
zi�����7^r�koTO]�h�r�4(������쑭��8��>H1�,(�2����G��t��M��i1&�m0�|9x�d��CX�d���=%9k��yoZ��l�����XL���쁝��)9��.�l>m�Y���f��z�:��hZ�R�u1�e�ˣӆg����a���O�C��хE����"'�y��gZ!2`$C��z��/���A��I�Lb=.M���W��a�d�fI�ʫx��ϛ�gs:�C�A^�5á�������5����>ÝBk��v�ŀ]�%���Q=�2Z�g���k�Ap�OI��@���A�ȉ���%ώZ�q�]l�ǯߧ���60݃��}JB��*w��nz[kF@��"L��n`��/����g�2
y���!yZ�u�ӀV�ٕ���c�^'������a>���#=S�9\�1����|�ƹ����Z%}��2��!�t���톶�k^v�{�GV!���������eY���wA�p;��.�}�m�5���2-x�*M������3�<D8�^��ϫ��-)�pƵAeH�v��i��}!�9~������#:�C6q��-�?4�Ճ'$�]�G�n�0��u:�ؾ�\���5�d�n*�y�O��;'��%�%լ�c��*.׮0�P`b×�֠���lK��hp��BbS���F��gLir�,}�'KT�Gҩ0��-���P�6��"���ٗ����١e? ���?7�B�k�;`��n��M�C�$�^���E�K��y�5�+wCn�.����Iȶ�C��|k��2��f!��;oJ�Ž�j72{"�����-&�p�i�O�/�o���5l^��/Z�0y�x�дrt'�^�ɼ�8S/=U5Ի:�5�qK�z�˫�^)�ٳڻJ��Ԍ��4�$�h�f�!��EJ�]�=F�ŀ�����7�MGkG�;�'.����̮xj���^J�ģ�$'�vh���[����5W��mp<҄@�X�=�_��7�q�߸�,*�O2�Ց�9]������VfǧEa������/��д�L���Eb���c�u>
����in�T�+P�9�]�"���x��±�y5�-����n\�2�w<ֱ<Za�K�)N�j+�VK�ȝ h�g\hv�9�\�F7V��mϞVG�`>��ib���C|<<<<��]�x���1�?0~lg�(����4-Xu+rn����A/mbT"�|J�(�^+6��q۶.�*d9�%�p\#�PC0 /r�ROe ��l)H%�Mc�1۷�7%tMb�x��c��g��Z��KsP�0�j��J��((���O���ܒ�ޏj�t:�Tٵ�FD��a\���˱ǠL�;�Q�8V� BU�`L��j�
yx�l)�67UA�k�q\���yRĮT� ^E��@�C�Pm�#.��\���� ���~���#7S���MNMA�o�{^����r�5�g1v/`�xe㐂z�+$ ��6�q����zx�n �9V�B����mL4h|`�\��d�}��j62�[�ܤ.{aT̡Fң���5
�s
�9sk�z�:{>�z�*Pئx�Ali&L8�v��2W�R���D��FBd�y�O��:D�)_�ŋs=|*�Ng�]�9����kgk���H|����_W�i��S�<yFA�ն��v7�{�cj��N�_���5zT-�.���¨o[�	��&c�/Y�9?{U�F���ӊb׃���lL��ڪ�\�K�������}�,=Q�4n@�v�U�VHhk
%�l���7j-��~�7��+��G.�p\�M����7ˏQ�N=*`�g�κ�Kn�Ι]��:� f�	 ���v�'���Ck3�������}�<�IS�sv89v��L��Ĳ.�裵ݵ�Rqmu�ذ��O�ا�y-Aɺ���zes.�`�V"M��T��0v���eI���E�r��8s.yN��|Mh�~����!	�	��7B��'qUeWC׭���6	�{:L?0�����CNc,�]�=�c�SP$0�l[Z}F�lħPb�>�-��
�0�j;���mq$����������<&�Z��V�x�4C#~k�.��	ɣ�r�M��M���Ln=Y|���Y�܍9��UK�����s�Ő�� ���������B9����r�������딶�ms�1	�^�#>�rb9��3b�;���p0�E���,����%6�v��:�|�Br9���>��_��zt*L�݊�p*7�b֡ 5L�=j�%��yz�}�p�0eLy�ĩ�x׽t��A��5��a �S@B}�ӱm���}h�����|fkvu�^A�}W� h�ii# ��{d������ޡ͛�Y�� %�o/+4\���k��m���]P�S��W.Q�b,*S��bd*LʈщGZw˻�����K�tĤ-���Ó�`*y��E��׍�ː!o
�y�a�&KͩKvդ)#�39��^�󀃺���ZB��C�ܒ*�c�z�n��W��iK������+�$2�������x�n��2�%ow��3e��xi���ǬGO��HP�c#)��jO�Q|�mG�3s{��i�LMm�zV{^�v�9�l1��}�r��V��9_Dx�.�".>��U�U��UD�l4��5�f�pܽ�0Ak&b�Z3IԘ�E�ս[�{lw� �d��`��0\���`�3kU����Y�;!
�a�jЂq��~�Fi�#)��7�9�<�۸��ݨ�C�N.���,Y8����:��3��� ��y�%:O�bS�]"��J�[?\s ��ZRA���;��mj������زҏ@N�mPT�m
�q\��,�H̕'��$�^S��<�O��i힚?�=�ONs�JT��Կɕ�~*�� ��9�k͵<�:q��c�.�,�noC��X���1�*�A�g,��^琋���:�M0� ��>0#��gb9��tK"�$�z���ۘ�Ob��jY��_���#��z�Lr�Aꄍ�7��$HP70>b_!�ߎ�wL�)N�=�MAs��u��sX����Г��ɷ�
���U,�^طvm��Cs�ooO����?/�����}��o�����=�����~AT�&*E��q=�Ff�xi[[�|-n���l4�]ت:"6;��M%�:-�c,�ݻ�PNi�4E݄�e`@]�[����#/#��v����݄h]��f\o�L�j�]��{BJ��g�VS��������]��a7"�>&��ǯ�L�o�5@	�W�
;��4��ɂ��J��!7����Pc/�+�9��q=�/u_�
��8��TH�ZZ���횿������ە����S
�DAV��d����&,ue_B+tXE&����^
¶�T�Z�x(H�[3����[���1��:va�r�oR֩�h`cm�
��
yZ���nSCw��)�f.cS�Ӕ���y�뭁`T*+E�=o�U��]'P�m)�^�2*�ͺC>x�Ь�v�U��ň/��U�Դ����tS-dU�%�w/���l�L;��u*Ĥ�����I�TWYN���AnR��i;����Q�;�M�r���5�Ӭ�'^�w5f���ڵ2Â��-����:�]X�ܘT��C��M⫽���j[��Ϊ�7�~��F{��R���͆s5O4:����S�o�mhk ����or���\���t��)���v1���^�Aru�g-o0ؐ�F�ݶ25�cY��Gw.(�oqW'� 4��my9��;�W)�p'�VP9�2l޻�T0*d�|�v�'�x�%���{����gW?/wzׁ�X.����Ս��^��mr�`�ܸ����l���Nr����0�Z�\�=OUF�)��_:�C|�f���t9�Eb�f�ۧ`*�����4�=��s���>�թn���I��=h�}���"Ғ�����N�mjm�أ����|�_AY4nA�H˹2�}�p��fd��t���h�E��r���C��lB�oI��c����6ބ���+
�{dG(	��2wW4G*�65N��j�b�/Y�j֊�a3�T�����[�Y�R��wy.�j1vbGE�.�Iw��L�Rʓw�73�'�f��Q���Ar�s6NP2,���Er�s�s蓁����[9�f������:q��M�NW4d���Ygq\[-�zx�WV�IQX��j������c�ɬ��kS���J�v����{,��]�eL���8�
�Å�i�6���F�.T�sb��Ч�dާPC*���H�}}�U��%<�|\tJ�RZ��X�F�*_8#̹�FHN�1|E>�6���Y��'#%Į`gVʚ7�# ����eI"̡&L1;��N�<���9g�b�N�&e�\9����9��a7B���^K�g�MX��`p��:�L"�y(K!�k�똇7WbM��d��K� �M���{��'Vo�Pu"��v�֝T�	(��������xwAv�qU�ʰ�Ȓ�;��;�
d9!�I��'*���Ϣ�:�zh/��gm����M�E�4��NPR[�q	ZA�J�����㬔�Yv�Q�5�/c�t\��JJ�PREC����Jh
��JR�4��4IC�<إz�HS[o2�
Zh���9#x܂�"SġZ�t4�	�ORbZ�j�6CS
i4&�E��rV&�9�N��S��(b(
��A�4�j����"�tŭQF�4KJsc���P<��4[!���PQ͍.��J���/#�4<�E,����m`��]�U�����z�:�N��"�C�a����3�$��,rӓ��^nL)]�X7{ �5��������E���Ӯ���`��e�ʿv��9�aR$V�TB$(�6�0|�4�K���UW��3`ɗ��A���4D B�XA���k���A��/�ԦA�k,{�.�V�y�����=B�z�r�/Q�8
G��h��L��B0��Ϛ�Ӑ�e �h'C�]�m��f�+)���Qn=�W\eE�k�lܝ��M���*+�/�
������X���M"&9���_u�Ý"w�f��b����nnV��u�6<T��y������/�56�h�)@���`�fDLw.�=9/��w�̒k�e���ѫ�Y��I��Os��̅��.�.Ԍ� ��˴��Zp9�=q'jE;�e���T2����Мz�R�竇v�/D�kWl%hBZ�VO���g͋e�2E��qd���|:_0��~WtI��w3�ui邹����j+����]�W�Uc��߹�/�.Á��D}�݂re�e'�m��������1�\:�^�k�1IխT)X�I�4�N����`g�]�F�I���2��\:��F4L�-����L$�B�Y�O�%75��ܬ-��ί�젒�t�M�1;̽6g9��S�]V�|:���o@�DcH�H8��!��3����T�{���{�#q�5�n�{�+��*=��L�B$n�'����/�s{�����*�L�u&63�e���䋁:������1]W��R�tck7Rn�	)
��̔�D��4�ؘ]���f]�U�ӛ[ΦTf^�w|�˳��2:h�;[M��������<��0{8�gso�-�\sq���(�$Mb��|��� B�g|!H��	r4j~�炩Ur.�Uģ����E�G;M��<��H�̎Ƥe�4�$�jPV`pC�fO�fI솣�6�}����Z���U��7^la�¬���Z�E��T�4��G�Oܥ"a����/#q)���������D@�<��άI�K���U�9��U�$'����ef�4���͑���
����.,��;B\�r��еn�c�Mб��%�D�jYQS�����Y�
0�v�p�rĦ��ù�`0��f�69�@|Njv]��mՅ*�n�#MCgM-nި��q��p�9IT�5k��U��X1��%(lG(���NK�N��iͪ����]�r����VnV��F��v��ٕ(��v�p,�S�R�E�P�[�����o.����Qό-zs)7,&��Ȳh�C�Pi��I�ʇD����N�
���Fb�0�tr����AO�j/�Ƿ`�׷a ��,�	諐�F�y��`�o���5^��O��(�vU�	�ɝ�:�hum�զ)����p�6�Ҿ$w���n�/)ōU��tw�.rJ�]�$싘�	��G7���e&�gi��B����	��vlD?�Q����� M0�39��MV��1�8�Y5p�%��;C=v��׵��������97�s��"a���g��%�������	�Ʈ�2�[r����PY�(�����~��ӗZ��wyp�)�똨~��g�DƟ`�-0�9�B��J�کnnr!6z�\n/Q�4����Z���Vs��_��d�=�0�����!W��lXG�pw¶}���'#)DaÙ(��m�˩=�����A<Js~�)�j�U���ʾŞQʭy(�${���r7Ë �;2^�pd(:uoO�ޓ�N�<^%�t9�y#I��p�Q	���̽��Z*7��o5;n�F���B#�-z=$2�"D�2��Y�N�XF�X9��#N�^1�姡b�2�wyWت�n���C/PP͌�����n��I�UYU��-E����a��yM��k*.�td�������`>��q����@���[ۄ��qTaԫd�����ɽa_j�{�]Asז@��j�<��p�F�.>���@8ȓ� ���-6o��iqB_��g5�vo,`�eOk��S�Q̮a�s���GH`Xh)�D=H�\s��[����xg�S�B�t����qG�G~w���OV�Ll�0o[|�"t�W��]�m?ocfBd�}p>��lfPV�R�c[x�ꕗ��C�$SF�*�z^��`YYX�M��
/Ch�_nT�8S�qV��#x�����mYxb��<���{�����wwAs0�];A��'JSGS�>�z�3<Ǯ�����Lg��is�3�_kU�n����M����V�.N�̐NM��N���t*e�vW����lZ���ggqZUwj��ы�A��`t�H�Se�^��<h9͜`����A��4'��fq9��7{IF�#���[��K�z�*���C�CPC ��{d���^=���i�i�kݒXr�6�1e�!���ͭ����BB���\�>7�.�
���0���/��ŖLLz9�^��>Y�ԃ�9p��Ddm�u���~@uO9�����Y!��6s���V�="��C�h�"���*2n���j�]�Z:�7aSv^|�y	M���xоٮW�Vψ��/ʭU��Bג8(�c0,�Ȩ�3voH����Z! ���EF��'9D�Oe�W�F�]�����t�lu���8�1e�o�\�@�P�>�du�F[�j�D������H�4T�ی�x��Ks��Z�n����b��z�U������a�`��$wR����NU�=�#'��@g�L[x5������5S�匡 ^�\z:b�hЁ��$8Hޛj�^��W��3[�����u��\<`Jeu�fv��:�l����Lg1`7n�J-�D�v\�Y�K:1B��׀�ޛP�aD��;3:v�K/&�D�?���W��L�<���ek��WR�W[f����k g�E�c�e��Ϛ�-�<y���&86p�t�Q|*��Օ���w�ۚ�u�/�� �A/^\^GR� �/������k�]�ϯ���Bq]��W������Z�`b�^(,��eooѺ�rĆ�D�ux��A�A�ڛ7D����{+���V2n~�q!��%H�4dյߏJNs������}5R͔�v���m���J�M���7�Oa@��80��?B>[��Ak+Ϩ_X]<GW�Ʋǿr��m�j+��J���0ñ���N[f3�K�lUƇL��4�&v���;�{L���I86��0V7��sC�G����ae�ko��4�-�}��r�妹XHCPT`�Q��*c���wPny���4������Ɋ�_Vgr2������p���1e��/ BV8!�T.��K���x��%"���ӝ���3M�<�S ���2-x�*M��$RQ�����"�O?E��z%�'���ʮs^�MG���b��l$W�BZ��!�#:�Y��� Y\��K~?C|wC���mC�v$�����u{P]�s.�y�>{n"�_:�'h�?
�O}yz�&���l�z��-Lw��QYffȷbn�\a��X�g�ܻ�u�U��|1�ݤkL͔�r��s�XѰ8�/�����.ǩ����B���?v.�en�mo%j�ܙk��~������}y�׿���_>Ϗ���Dg<��=0W5�	�y��7����]�d	cIuk=�|c\�K5$�&sD��z��й�C�p;^@��mh��S]�gX�d���2�E�:+U
MٍҊkq6Ue���9�܋k��n��r�q��"y9�k��Iڅ��}ٞ���&!2O��BUe҉��yE�)T�N(�ٶ�Шt�z$�!�6�Y},�4���lHd+�R���J���rvB�ukvPa�EH��/���0ю-#a�OŏV��t���gs��[!@� Kɧk3	<�)�Ev�}�H��MPI�Ԅ���y^ɺ�Q՛-Ey�v��zz):�I�p�a<,�熯Z�E�ʒƀGjHO���7d�mJfJ��읾����-7$.-!��󨦺��^���!w�E�Z��3b�k�W�B�0�M�i�.�{ )<ՠ� ��a��/H�jzG6��4-2�n8-���f+a�P=M/k1��K����С�ĳCU���Ub>%}����Y���rQ징�1�ȍu����5����&�6�p�f��0�wKu�0З@~����w�W�`a~rq��� ���%��3/�+V	nk���f�쑜b�=��t[�2�K�I҆�F�(�.�O�����w}��6�󡜩�ޱ��׋ߏW�u�} DO�����{���R%qt.%f�!C�M���ӄ�39��Wڬ��Ȕ���U��!De��g]<���
ڴV�#�;A~^͖d�$��bu{(�ṇ�hQZ��)GO�i�&$BT.�g��Ї��G\�.��fyC��HzJ>岌�Y�&�C�}��+�3�
3s_MI�p���q��$�K�=6�<�7a ��,�	諐�F��|`5��0��Ѵ�qf;��e����
)�0BaÔ�D]���Ʈɘkl�ʂ����,n�OȻQ��2��'�۲�^d� ��dp�T�.������� C��i;8�l�74�(�c���a��npX��9�zҡI��Q�`���V��+(��f�!:�L�i��7��'hen��S�ݶ�C.*KP~�I�x�J|*�B*��e��ކ���z��y?R��m�eVe��/�N���z�|k�7�Ru��YY��44�P~��tˈO��~�aa=!Qmv<��^�a�$D&	=	�A� B�4����Rt��]/s�1�b4����l0����_ �*�Y�6f��{��2d(V�ɝ�~�ѣ���w{'�N��ID�n�^�c�o��sk,��dǷ2��֏\���6k�Y�
m��ih�b`�l\��2��AR��ّ����yF#����ԇm0�$�$9]v�7|�T���Ql�(��U�}�$
ZP��|<&��7����Uo-�wop��A�li� �t�Lt9B���*��QQ�L�U��Be+�k���b���pʜ����((�O�G� !qX^LItd�0-�܊�kcu�!�u����[P��-p܍���u�y
k�A<A
!��5�bu94s����;���k"��ˑ}��X�t�8�\�J	WJ��?uԓ�Y	�a�P4CՑϘ�nY[ZӶ�z�������vE�^����1�����dz-�fy�\3��P#��@f:�y����0sH�y�C���Gj�S�ج	�\�dc�_e���lc�C���;	y>a�}lY�սqJm����������-��A@��w��R�ht�|.$�6^5�]#�4��0R����M�+���f�Ġuafz���N�/'�o�=3r���,���҆B�=K�$�^��h�C�sqSw���Aǋۋ#++n�Y��v�a9�#B�w"�o�56����X�d����G�Զ&>���|%�328�7[�ܵ��U3u��R�����z�����o
�E;�,���U�~*=�㊠�ȫ��cNHf�)��N?��|;�äQ%�L�W�ؤ9�ʷWS�������[���[�u��-���ϣ�Gj)����tiF���w��+�Dw��ޡؓh��#Ӌ����nj(��r4�g�v!c7�P��;_Ϫ��$@�R P)T��(L�w�1i�zz���UZ�+��W�w)����ɪњOaQ�a^�0��\+�Ä�����y�ߚ�^
Aʺ~���k�KhL��ϯ�B#sS� �W(�I�1,��I��F��_C�HSa�d*����y��E�g�A=����2@Q%ٲ��	����<���'��%9��)�����fv�,�r��둻��̲.�;$�>E����3cH���hmOU�Y�����t�I�F\3Q���%������z�9�WP;\Ú���������RG��C&ݘ���Μj.�K�`>B�Ȍ;p�%<�N�R�m���Z~X�A/AqyAt�=���`k�tY�Zp|J���r�F�%��v~ZK�TKj�խv1J/�5����r�Aꄍ|���@qYb�|�I��W���<ځ�u:��hRurdS2j���O�}����ū�B��l��wfԭ�m��{��27oWɃ��P~Ǒ��zP��Yƅ�u)�S�X��S>��Ӳئ�G�/j���C7��<�-�� �J �tȄ~��Q��BX��H�I86��0Q���e�.�{�6�Y��V����ma��Be�{��^�쨺���uAx�X0�՜A��y��o��y2��I���Y�;X6
�x�S�f�RC_�f̨]j��@jٔݣ7�҆�u�gR���y��;3 m�
u�8o<�@��I�X�}u��7ǿ��}`Z��A)P�
E�V�B��}u�||�o7�l����E3M1妾�a!5@���0(-10�͉��_u�4��m۲�w�'g�S,��.Dev�J��k��GKՉ�z���Y"W��A��\311ܻ�(�}�xZ�'9�Kr-ưҖ��y)�z��3I�<�S�z��5���6�hl�wq�ͩ�����y�/�k�&E�	��Q���^[	BX��.�g f�2��-�:T�M**!Ϣ�t����.�"�!�|Ǧ
沂[/6���!?5�vOAd	b�N3�p^���P�%wf��;z�^���sW���%�P��N�jɅ���2��b����-znLYX����{f����ע�v��u�D|���t�z�,�A�v��n;%73��//*��Ua���n�-����:�e*��N+�f�O�"�t�z$��q#fd���ͪO�<�������d�K��F� \&)y�E�$`�0 �f�xaz2�h����_�oL���+F9S�OC	cVU;M���Q69N2.���+y�m��~g������>�_������{}��o�����յ����c,t�m��6+�%��pP�)b��z���-$,�T��{��M��J����Ƌ��"{Ё�����Pf'��0��4��rb�S:��B`��M���Ԑiκ�-�9�e��F�A�R��g��ݬ���?k����	AU��-�d�5T��������h����e�����5�To),;�]�w)�]t.��\���Bsf)2�>��Sg+��R���|cv��3Om�]j����f�˙��O���VF�پ2��	1;d��g$�A����7
��ff%����_D�|�]n�t\��M�WY�d��%M �������V)Td��/[�i[G{�k	�E��ب�*
PN�Jݳ0�Ű�t�t�脚�meԶ�N�y��6�mҵ��K�3um�.������g
7(<�=�e���N"-k{��ʳ�A2�d;35D�׷�PbWj��/c4��A�XȮ���u:v��.�tj}��t��'8Р)�W��g�#7HF�]r���nw���ʂ�=��ҮOC�3ipQܳC���	�W%�s2�_T�yj���{H�㓡]�S+h�v�ИX��0B��pb}� �u�E霹����K���O.\$X��bޭ,���B~FƸx�5WKz'-��w)�z��GW��K���0wkP-�Ի�I�Fn5�8��knB�G�LKj��d�ǵ�gpz�����wH���sZW�t.���Z3�\m-�|:-Ե��5��)\��;� �p`���t���ytjo��x���Z�l�;SdYS/���u+5�x�bl<�6,S쭓5�1\e��5��@\ƸI�ٍ������`*JR+V��b�i���蒸+:�.N
u|5�*<Yy��7W\�Rb�2�6��yrݐv��hӼT�N3�q,f���jFXy]9n|���;�컬O�fnҮ��d���m����f�K�[��#��a&1K�n�Z;I�15 cv��љv�',�H�k@�:n��w�*j,�r�g(q�V����2�ƻK۴vҁ�2
&m�K�]�H��s��L���XT�7��;Nd�f���7�,kÀ�p8��E\s��Y�im}������yA�P��Gb����v�N�A)֝����
U`�+�73�ek��0v�pGL��%���z�*��X��k{�� �{UN1�9[�%V��xx�2�lS��u�fr�e�Z)���E����f���`vVSŏoP�!��83��+8ӃMT�2�vu�j�bsqVn�*���	�F^��`��SӔr�{�����]OWd�:���(S2K�7X��c�6��Iρ�x�'r���Yʃx�)�L���E��^,w��1�T���M��#��uYa��T7[Y���/D��Ƿ�Ƭ'�����ǚ����"w����7��X�S�n��z����j4k@h(:���)J���s��B�h4�h���97���
Zc�V�g�:9�i1��l:[m:�Zh(��.��s��4�h

"GHh4&�h��j�4RR�&�M<�C�������Tѷ7�PA&���X�m�"RSV�((�-��QE!l�
(�]F���!Zt�!T�k�G�<�H
�)5Hm�)u�5��%[b��/!(s.�4�Ɉiкti@�J4�j��QC��:X��N�un����>7�����S�������d�il�Z���S�0d	_o<���{�[Gt�݇��y�����۱uP����{���y()D"`�B 
��\dq�_3�\߽��ב�$��%Ή7B��¨2��Z�E��T�4�*�nmv\˻���o��c�$O}5�	p���-�qzQ\�Ĝ�e�q[�*�
���fљ�d��:�bcwMwgx��t�U���@����ళ>��1�	��Yƅ��X��`����MQ��ꞌ��m֨%�T���Z�%�6	�����{��B=��v5vҋf��W��3љ�=�G ˦��f�&a���/@��d���iR�e�"��NFe�woC���'%ؗV;����,8�me���3.�7[�m��<U)�)7�߬И����Q�YJ���'tF�!�>���mX;��^=���Pi��I��}��:q�jT�ɿȧh����zP��P#�^����Y5�f�#���#�(5�0��E����=�ꋅY�,��������^dr��Þyg�XG�:N$E�֫�j<iߪ���>���r�(]�S���.m������n�
��G�=oN0�\�C�ئxB})������.�d@_����	��]���t��3آՅh1�X��!�#����{f�;c���È�y~{3@pe�z�����	Z��w�'��YT�eMU�©ou��(v��L�����i�ƓV�/�����c�w��=2d[0�W��Q���t"U�1��"��yu1��T��/�+����
Z))@f�f :��:'r-���%S네&UiP�������ƚxk���1l�A�����2�������W/}\�Q.� ��g����X/��c��kس�9U�$�j�G�����d����9���o��zw�Ru�/Ⱥ���#)�?E�ֹ=��}��������j-�|h3d� �\�'��4=�H�@Y��"�Rt��5(���Ƕ��m�T�T+m7W=�dorv�X�� P�*�ޯ 0Z�_�>w_��a�l�*�,��xQ�1����<n��Լ{q��;	��%������G�:mi����3E���KTj{F��@����ڋ��@��R��~�5��Tz�Z�#�#|F�Ѓ�s�p9�S�>�v��6�b�Z��	��r�Z�PK�z��(�W0͹�!9r+��]�]?SQ��	�X'˱�;s�{wd����6�ʔĲ���ϧ��m�Y���k|�a�TRD��"���!����|���^����7d3l��E끏IŜu�&+�xz~��Ջ7>��Jh�,���81�����2fdx6�?]t9Jx��f���^t�2B�RZ7c6�s�˳�(����:�xK���4�V�c�%��<z��7Y�ʽ�e�yp&����ۻ��56V6A�c��05�R���|y�kߟQ�σ�ν���}%"�R�$"���h)������x*&,�8�Z�[�=s�ʾ�	Gk��h\D0��H�ٽQ��$x�s9���
��\��]}��-�T*]ݏ'~��ѽ�:��2t���CDi���O�+=��*��3o5m&�ۛ����{��i3J�Xu%���I4]Ls�qp��KzR���_����e9��ٹj�Jv�rr�]��q�38ˎ�f�;(2���RKˬ=���z�o
�H�x���b��}m �ұe�+�y�\zH�*�`����H$�B��є5��d=u�C�~Cx�{�umޖ$T���r���� ���2
"�dQ���?B	�'�I��(J4�빺m������+%�o�x��+�Ҵ��$lr�D�Цx��lH�n5��r�\���Ǿ����"��^�g^<��k{w#��E{����2P]>�!C64��,�Cjx2�a�#�o��z�R��B��VcL/<x��61<��(�X�$R��XcP��?�s��[A�yȄ�[S����S�D)F��۝M_qh���-e��.�君��='�|�A/Aqy�%�a��ь�
8J�����x?QL<Y��	xԠ3L��_��g%r���5;d䫼96�.U�㛛����;<D�)Y�̡�\ܩY0�����V��='"�2�����S�j��Mj�a�بm���RWW(A-�99�	^N���ʁ��e�ݧ�J��3��C��UP
5@���H��R ��&eԎ�Ǖ�\}�=��n��Xn�6�TWzF�[�ڮ^H9��(���g��U�=r�)��5�A��|u�0��Mzz�s�dS�V�cL���� ,�*�f�܍�u��)ӗ�/k4���H�w�dJL��D��|��?>��4-[�L:�Ʋ�����v��YC��k�)����
�}�h�0]X�Жҏ�^��A����RSh=SIpF�j}��7�<]Y������XR�������&<�֫	AP0C(���X��]Z�<5�Ut�YK60+�sy/ݝ"��j�.ŧÌ4��U����C$JQ�1���w�U�QIS����:��kof�������;:�npoO�ef��='��%6�5r2E�	��L�f�2W���mva��z�g�r��aqm���W>��lN2�H8吃�VIA#:ϛ�o"cpP+bf�u��k=���2��ʒ��z�!'v�y`s�5�ͨ�m�!>� vO^YX�X�~4º���	����-e���^��N�(p�aF��	�h�9�M^Ʌ��t�����W*yک�1�X�#{"�*�Q��n����e�CQ%av�o22�#��Avt�L��r�T�����e��yJ��)��~۬���WX�mY�5���u��3��FD�h����7Z�`��U�S�����1j�۸���l����M�UJ/5Y�d��1����W�ՅIMR�4--!LIA@R4�4�O�^�=|���ͯ���dO|%RaMAnN5��uB��� ����]4�N���f�z�����Rc��kb���A�9����%:�Q�jªK}2fm��E�*���	F4änx�X���5?N�6u=�;��:��-�b@�e�F�*L�0a�E�$M�Gؼ4��e:F��uߡ��[���5:��C(}	����ʼ,�v�0��(�\�Ʊ�x��s��E��������uw�寬�����b�Lާ��Ӭ���J�W0�es�P�r�͕%�5ZZ�h�&��<�{֡�3��f%k�Ǿ,��^���S]s��{`-��.��,B�^��af�����y�q�z�qnB���A���3 �cS�9��k��b`�T�F�n5��63Zޖj8�=�a(%�T�u�-A���y���=�9�w��ulc��v�v���>d��L��=5�K��=���}��HīU��vD�����m�	��(=,��+s�r��^�r�'6;���a�,(gE��/T1�J!�hzdG@�t���b���#1a���ro{�䅩��튖���Pج�L���^��@�nx1�g�sr�٦,
-��Ɂ'8�f����RC�o�b��i~W������狱뭘��C��J�x#a�\:wk7F������r���^�7��n^n�̦u��Y9�[	_F��ڙU>��44�LL�RQSx����.�X���8'�)����2;��f/"�y�zA!�(4�2��Ō�&��Sox����
[����2��&P�.&3%'�&���6>���C|a���feZt�fm�S����BF�O���-^鋇U�`, Xt��嵁�]�ݿ��������=�>��uqυ�7 �(Q�ZVy�ׅ��	���5�L������K]��]�/��9u�ww�����*����s ���h�L����vNk�ǫxi��v���i�����2�Uf�ۮ��:e��	���{^!���5?!)���)Օ%�j��w흭׻}Ǆ棚���ַ���
��_q�����B���*� <0קze'XĲN�7_��ߒ4�V��)���c�u�|7�v6/�m\�j�5pņ ��O��9�	q��h�*̧}b���E�C�i�2��Uc��y��.��G;a��I�Tc�C64�8Bn逘�r����')����5��7]�#$��#�ŝ�s`Be����K�:�����&��#[��������s�@'Z��M����*���(����#ߘ�ؙV��.��Ru*�	K�%��DXz�b��jټƚ��a�{�P!�w����s�F���Q��tV_7��6����]!��ƚ���1�j��8L�9��p>Æ�n������>  �a�bF����珞��u���x���;����7>�%F�Gs��t;����@��x�G��`e�G��9��1�Q��z�f����2%��&�[+�c
��_tn�������RNPqd'!�|P*���=CB}�h�]����sܦs���v�z��c~��1X���3�Ǣo�\��b�f1�����>c�0޷���n�\��@fhP�ϡ�_
��\�fH'&���5}=0���艚��D�U�SQxemcM�}��TY��!��R�t��	��V'#ػ������
^4gS��Ɯ����]Yz��\3L����X-}#"*�D��O��R����=	1x�cb�s_8i:�hӝ�[!�����$���YA
徭����U�mA�U�#L����Ǟ/y4dտM��H�Ӑ��&y�޲"�uL�geK"�Б�^͜OC��P��j;\vb+�,T��xC6��u�(*�`M�EzGq�Q�1�f�Ϭ+5L(�^<Vj�u&&�&�����]'�x�$`�`r�BA���S4�p�(=��l����a�	c�w蟢��R�:o�m�C��nRWe5�Ut�0۽[{{W����L�}����x�uł���O&m����=�8�92�^��mF���袩}p�ɝ�e�p!CGA�����ؽ��!
�:4#���cX�3/Yjn�Gj]�W����j���*(&�z�翟�|�<m���C��Y\���#P��N�}@�qBؑ�E�֫�<��νhTu#��ۼ9�a�Y<���"��%HA)v_GG���ʼ@��߬z�~xe�*T�5��Qm��{�]Z�ݤÄn���E'+9�R���j=^��}�l!#��M��S��c��^���#+�'���e�A�M��9E��'�J�z�:�4D�p�b�ۖ��[U�8���h����K�����d��i��k^F}�7K���׋�����1җ��2j���h�;���!kR!��z�s�^E1�dյޙI�x��yU��n���E�$߭&;�O�4��n��z3��G����k��=ϵ�hZe	���������~�pr���5�0��M/TVg��~t!!�}�2�.:Q�e�v>�i��&�xƉbi�c���"�{5qHSL("�;h�[��m/a�@j
��GÖ�&;�v�'z�*|5XO�ÝbW��2y[�B(q�.��]���i��W��Q��%.gЗ��G�;݄.�sx�� g�,�#��Ī��d�Y���
H���gc���˹C3��H���1O�:�i�=Q��+��w\ͩ;�&@��wnܻ��<>x)�^b��d]5�H�w6V�����0����4ib0��0+Ry�H�*3o߀30f�0��u�G(:᫛�D�N��ןm�v=�זi�k���v����a�m�?4S�\�����aB�c���!�A�e�Q���Ea���
!-Ed����;��*rQU��ݮ��'x\+�����c�z~���0��DP��߆TV5yt����A:]FUFuQ��ˊv��ʢ>�����#�b�a�&���uB����P.��q�&'��F�mɅ��ta�\V�y1��ۈ����:���B��T�S-���z�]q����Y���	;q�c
ɇ3��ꕙ�-[�i��L�L��$�����F��
�'q�l$vE�*�� ��ޒ�%V�]��/�N{f81�_K1|a�=�J�,^b��E�)'�/ E������6{;E��T��Du������!�N�OH@�{	eBʧijRy�Sl��EM4�{�� Ы"\,O]����۶Ew�⼻��a�"کqZ���Уxi0�0��W(�����>~�*�h��]'8<ʏ|������),.~!qs�@��S����}B��[;�/��o����ӱ �ݻ�P�x����.K���$�omn2���6WD����(otX��;aw\�
&ք��'�2��:ҭ��� ���x3R����C�h��Q5S�޵J� d:Qn`���%����"�P�����ѻ{���� &��,�ЧVor��%�ʝa���P������H!��Z��yF�_�&T�gy�L���u\���[#mƠǥk�*	{k��-�]���eCWBQ�b�ަe���ܣEgB��J������M���,n##�e�Z�L3N0��@��3��2%ޫ�T� ��^z��D>,x�o���v)���Y�p�^��nǠL˴��cU��Br-dW1}��w�!���R��Lp_G��U��P����nI���zA!�%�z��h���d�.�N�$"�v�f�����F��ˌ��I�j/�5�2	v�xj)U���WVrf��\%�I�4�e�j�L\?PqEx-"��܂����54�v�Q���]�w�{u�r-�������fP����,��T-�ɲ�p�8pBҷGk�I�����_g_:]��Y+j���?!)�����
��B�ڣ�.�ϱW�Z�"��|�cs36h)䇖o1g��ma���(O���4��<�W���Yx��,EP����4{=>�_����������o�������N09&z|�go�e��T��uL�7t�h�3���KR��Y����::\�阏<'h[\��[b��wQ�f�2�j��$u6��'.���y�.�s��vU;
�|��mu��/�u۴���|����8g4�[��)U��P�J2�,r�����o`���[�:c�z�&ӫO_l���1guSYY*�]��D}�S�M��X�F7������>��K�jm6���K�A"���{��vc߂T��������#׌G}� ��#T��l�qB�ٺ�3_t/)����!ɥ�ŧU�o�C���;p�p;j�Cu.2s�x�����r��0u�d�Cur��M�]}�hc�rz]����Υm	���Ag-�rTԶS�X�>rrAut����b�vQi�W,�p΍��	kG�\�F�.��'�Q�d�ז�u'3z^���n�H-6�3y�O:%{ǥ��w��|��K����74��2�]���Q�f]�j!#=J-�+C13��?bp�ۼ[��4��NJl�yH\�Y�����3&�a֣N����E�9zgLF{ٱS���S�;�/�u��<w.��Zͺ5ݰ�)�9$�z��vnuѥ:<ېBԢ��q��9;/-�P��xj�"ۧB�8n�۝���壊�(���<悴�N"t�DF{��k�9&>g�1:�h��.=ɿ��{aB�8=����J��b�����ä��p  ��6�L��o˻v�7�\���3*�y�1Bm�{��N�-"��*V=�҇���ǹ�}�;�����*!�-������H�ɕr�૾�
�!氮�z�[��j�|�SN?���ֻ�ë��.���4�q�7�Uɖ�{�S<�n���0��Whk��%��������z�CJ�����Y|蒹 �XM��q����Ř$�7���gVIy�ЅqoK��6Cp��͗�����0�oG'��9��U��CL�qj{[7@�n�%����)X�whfn7����ui�zH�T��6��k�����j�ԕ=�ie��۽J�N��r������ؼN���롚8�450K��s���Z]��KC�/�vݻ�h���R�<���w���%f��`[��ԡM��	���n:��P�eu�m�]�e
Tvf��ٳB�j�ܹj��v��|cF4��`�"V"�9�`̴խ@�����/x�N��.��.sV�*��/rwZ!.�Cܡ��K
���i�x���r�m�u���f�I&�M�.�V1q!!�*�F�7���>ՙ���l��Ű��x*�mgmy�H%%²�m��}s�#Xy��y�*�O�����i=���8�hWL��t�3��_cR<}tIb�e��j�5+AYv�O툝�c�q2�P���"�e&��p�K��V��WM#mtYz��ӳ���#T�����ڜ#�8�6W^L�tÍƛ]���_���ޭG=�{�|Q4%--.���T�S�4���٤�����l%��#E	�E#BR��Ć�cCE)BQK@r9
rR��)6�h�4�(� k�<�6�����-��&�"�+T��(�9''KEh�4��:4�i�6�R�.�4�]����:(F��M	C�
9�:4��C�ZK�N�.ً&���`�IF�SKM%&��WQ�(��/R��)�ѶB- ��!\6l�UQ�@�iNH袐���r[�Z9ptD��' �ki�˪R�LF�@kh�kE]+I��)�)h
Zu��Tѡ+?G㞣ߩ UB�"7�?`W-���S�C����'1�xLU�cK�1���b���Ð�R.��y�[nJ^4����;�'G��]t��4טt���4I�Je���y��s�{�>f������
�5�������3G*� h~3�ޙI�g�I��W�2���C)�����O��٪X ����fT��}h�l���sО�װ���i;�b�q+����M\�_��O�/��aRs��iCa��I�
�D�؆#���	��ȓ�0"��	��u�SA�E�r�k��Y>�N[�,WA����K���g�#��M�B8F�S-nc�^`�U��Tٗͯ/�˩ʜ�`Z����*�*�mmX�گ���T��5�$��M��b��7�T[c;�Ag+�sG��Rkeb�aO��R�I�=S�R�iWRN5D&��#�q#h^pͼ�A�8l�v<ñrӓۏ^��6 �LB~��F}8��s6f�5ީ䎩j���d��ڠQ���W��P�Ԍb��Ĺndl�/��c��e�4�Ɇ^�Ƀ�D�P�p�=]����ZŲ�C��bR�ZDڄ��z�	��.�|��ݺ�rկF�tjh�[���2
�4=Z�iՂ�ӑ	עJ���<=:j����>����]׍*vJ�@�m~X1^n�j��_rpO0��>���s+ʻj�ٔK�!R��i!��R-#vI��秩��{�B��8v�m��k�2�Q��^
�m�w+tɌv��vs��U��p�5b�W��J� #.��*;��������%C�Fnf��,;��PB�Iw7�i�m���)/q"ag�ޗ�
�&�����r�s(�T�&=��g�䩛��R���#��l�z�o�Ǯn��ܺ�bv�wtq����"�҅U��6���D&��2�&�Fi=�Q�`�Z��EJ�wN���t]o{sqM���x/^��x��de
,.}	+�Ab�j~����;D��CW+�OyL��^��E�z�Kp�uK�(�����/�Ivl��|$>����˩Vޜ���S�8k�n���Μė+�KIRkk�<��\:�ty���	K6���d�E9����G7�3s��=&Iv��W��R[%�1׾s����lA���,i�Ot�osLM������Q{�.��M���Qi�by�{yH��]4�O@~�jd���4�������(֑�q"6%����k�n��kX�2����#ʭ�mWܼ�i���F*t�P��4�O�]��q���<���@�`�D;|�c�O:�I�Lk�M[]�2���`��y���u�΄�ޔ"�ޫP��֛�S�xU�rWk=�f�Y��iVE
��Ӷ����M[Tm���XFe�3`���
�n�c����5������|m�5j��C)�7��cy5\1X3p��bţ�a�E�sx�)ea.Sm�V�hli|.��{$~	�}��q��+�w���Y��Ͳ���d���_!�j�.YC�h_X��o�6W)ozj�q7�=<��������¨�b�a��Br9 �
J��L�X}��!r�jN��S�R����/�dl��u��h�|�h�z`<���}��-:h$ExS�,YU���y_�6w�v���ݭ�p�6��$*��7<���#�Iv��]�O�B@�z�56�k$JX<ڏ+-��S�����S�\������~e�����s�z}��3I�<��M߯Ѓg#.ӯ�i�6�#��3R��d	'S��`�5�~�P�A񅇸�E�M\���b��l$Q�A�P+$�y��;�5LL�+|�g����6Β�c^��_�]����0BO"1�D܍�J�<֎Xe_��p��̕��Ǘ8eOҰ~��e����� �`�=���~�`�]H�.2�'��t�&��W-;+�]��Ύ���۠&#C-{�*):u�xR�%��]���8��:��x��:	�;c����N NL�ۘ��h��b����L��xN{��U$��b�u�4.8�o7��P͚�s&Ƶ�lm-�����^_uq!����U*L�J{�ԦN`�8�D�YA�6x����f>"!7�:h�j͔��7*��5,�ݲN�:�h�Gz��o�JV�&�.�.���P*�@;��pX�0���W�f$�pR�V;�6���*����3�
o��feB�Y�i�˴�R���LU��EH��3���s0���Em�CO�����v!?`��Az`K+/�0�f�D��q�u��cp���Q�J�]���n�_s���M5A.)��v$t���=�B��«�es�N��ZkN=g �MgZ�)�s�k�*�P�0�ȃ�B����ꯝE5ѷ"�%�Rj���*}��GY�ڎj8�¨��؜-*u��+���j�Q�Pа�!_ؙ���˂�jL%8^8�Y�B��Bպ����{�F��;(Nj�N@pq�<�ՙkm-����Ö2��>ԙv[]��sW��@�.�ײa�{XX�[��/V�i�Z�Z�~>���ck3��#:!0gso�9 ;$��t�t��,��%ڇv�rb�&�j�[���]��n]�'z�Y^RԥÐ�ڲ��*<{Xn��z�k��������;�k��R��$2Qc}��C�U��(E�����^=�k�H�?��XC�3wtm�굛��-a����-�2�T��
��6U�Dr7�
���I����T�k}�
Q�]��<��V���;��cevt��XBn�{�N��b���Յo*zm7��m��m���\�P��[[��h�ۦ$����\����L���Êi�4�[���������%r>�R�4�����:b�sRW��(�E�֭�;-�k��UQ�ݧ��mg�������ƭ*B�vd��IЕp��8�nb��ؖt6��`���6TY�����\�C�.Һq�XU-�O�Jm�#!2�F�'��vsf�cռ4���<ZrΈ�i�
�g�2d���
}^!�sh~BS+/�X*K�!B���·��L�\�e�������([0��{��AX��D1�s�|��m���t�Tf3h�����ǍW��j��,+��qa��׆��zA�lwL>	�!�a%P�I���+y��y�l3�V_�!�R��(����=Ca��I�*1��li�uuHLs�kMVISWz�[9�y�r{(�(�'qV��?Z�O�S�$.���4���:�)y����h�����W�#�фs7�7��hE�xI��˓6����z�w���c��k��85R
>�{�����X�=�F,b��A�������f�U�Rkea)��>�UҞL�]I9/�څƬQʋ^���7��j����61�ֳ����i����s�%��{�*�^��]XV��<v)�-�S�J�l�l�,6�i5ܜy0�ӻ�+��em=A��9eKCb����&afI�x�W5d�$q�{��mo\�Ym�Z/��������l榒�p��z�0gѰ�]ٵ�^L3n=�Gz��1��:�-��X��)�ˋ3cu�!�ln�R��K�jl#�LO�q{U�B��2A9?[����f
fB�EFV��ު��p|h=yQi����tӱ츔�pZD`^�&%M��N�k�L&z���O=��:m��ݝ�A�{�ki�Cף���Eq4�[�?�b*�Ȗx--(d�	�1��az۽F��c�=�@oP�3p�4�zt�C��8>�H,�M���%xc6Ov��kf���ЋS/29�'���;�t=\�q�J��� Ȭ�`Y#�}�8��Kn��;<Z��I����K�T	K�Y��H�����ݒ��7�Sm�A�P�f��ZY�fds��V|w#r~�_�x�7��>� ~�^4�aw	�`��[���v�Q��C�@����渖6��%�IjQ��C���ȧ�x�J�.͔a0T/D�#�sJ���i���'���cњ�:�Nm�@�I����<��\:��@.�m^���������O�k�aȥ����T�׳ە���g5�j��'�­;�[����L+Xsm��~����i̼SlIC�70{k�A�kϨU)�!�P�W�yu�^����pꦥ+�� 5���Wf�����3N�3�Fi�x!�-Il5�����.�Ov*��0��y����ݜ:2ȟ�1�,�`d�a����$�^Tz
C�E���,9�=�����ly�י3�lğ���{�����]RC,趔��*]��&�z�����w�K� ������/�����T��Ύ�h(0�a^O�`C��=Ǟ�=sM��q��.xV�kzGs�0Я�.l�[n�K��g4��BF׊#��:|���ٓ�<��L�c^2j��L��?����/�Z1(>��0���L�D��V�"8'���xK��W�{B�^�8L�����Mo]��	E�6�;\�N�ڊf�g��~t!.+k���ŝ���U4�� �U�4wd(���Ξ����[R�z '��8���,��ǖ��a!�*0C1	�{v��)y2���wY�[�vx�<9/�I�����A��Ρ�h�W�˱i��$�,�jmF��wP�	U�P�ҋm�s\1.���t�"a'W����s����2�8�<�A)�A�F]��'��tCȻ�R���r�o���E��z�Ȥ�x89�u���8�_=5���Ί�Z���ϏӺ��e!���E�vD��Y��jpM���kB/���vΣ�,�ǨLk��_bקoe%xP6j����fJ�o=n
� ~y�x��Yve���2;w`�����u�V�^�3OK�"�op��1�z��`�����{����dқ]������l��S��ٲ�6�F3��8Ƈ�Y\��J���ܽ�/yQ�M�����C�l��C�Re]�ca����l1�����XV�j�ʨ[�\P��k���"��E��J~��4�LNb&b��Qz�k�1IխT)\�L)�vN1�����3��	����A��ŏ2��Y��LԚa'j��>���~k��&��ħ6
^V2/ʩ'b6m��E�"n_^cQYV�B;s�;�'o!��[;"l?\/���ö�J�,c1C�I}	@�v�I��L	��������f�x`� @@�Ƙt�OH ��l�v�5)<�)�E�Q�FSoM҉;=�:0����e<�j�e5!f�;�Cw=OE'7&�Q�4�V�:jl�£%OwkF�n�%��ry�,H�z�'�vmļ� �\�.D@���ĵ�kGQ�$E���KSF�}����+]�J����ua��,5�V��26���-��i��C�T��ݭ����n��[�¨Z�R��Xeҵ�%�J�a+hN�h$�W��8<����d��sx�#.��rȜVmhLV�.��m���c�{(��v9�fa���/Ɖ���%�����1�1�{��e���ɮ��{'7�]��v�t۝;b�ۦ�j��"�:��N�WǗi`�u`�>/�q��f������UW�Y|4�K6Ep��������7����'e��l���@��k\�f�&b|���/���d�/�,V��۾�[�>*�)F����@Qi؟J;˭�$�{}ZE=��k粋�Y!�X�L+�>���f7���1v�V��b���d�H�/q��Ƕ��D_��)��(�� ����H��{�t��q��0��T:&���fq���B,��Fd��&���,�g� өj�x	����]��<50�z�������7o�C�.P�ʏ��}�?~ɼk�'�~
+�"t�:Q�G&a��.R=���*2��h,qdT)��RU=c�v{Q�X�#/n�<�2�1�>�]�-�boj���?)�ѐ�U�B�ڣ�.�zs^�5�Ϊ��"h1Qi�]gOr|xd���ҜI�0���>�S�ܼ!2,�T�	��^�<+��7����緷�Yk���T�%Bc�p^�f�z���D���L�����m��x>�ھ8��f�t�b���t��8��w1ʾ�ց �6H�L={Et�ӄ@��tf��oc�נ/EP�0R�}K����8�Օ.]��n�}ȹN��[X��p/�=�%��d�͘��p9�N�D��i��-*�) }L����tа����E��I������}��嫣Ȇ������P��8�)��pf��F�g���`�/G9�Es��Qu��Ǳv�����A�_���Կ�|g6��K�	i��1
b�e
Xd���*����L�ѧhs���r��Ae�D|�Y{r��r�;'
�؇�'˚S�h���h�6��'(]�*�=,��5j�w=�9���gN��N��gz:Hp�X\����κ��m;��-l�)��]+^���O)����z^Y(��~DN�MaS�"�<Y	��Appp���������6yoO�U��Z8��z��Twb,Ԏ��̇�c!�R�K�g;�Ơ�v��8����.O28��c�Y��oo�L�v�p������z%�%��tE�jb���w���h|.&%M�~�1�R������c��l�_%A���X��G�D�&����H؊��� | ��-8qSmqI���ѣN��1.�������Nnf���u��ϧR
o�|�56��&�1����"Կ�i�,:
���U��ϊ+D�����[g�%L�`��d[ڑ����=�/Oo���}��o����}�ߗ���|��߃��E�e��W�d�K9�����`���l���M'w�j�s�G�7�V���C�u���*��ē<P�p��a�ZR텮Kzk�x�f3{�GM�Y@�U��f�5,�U��$SY�*��H���Ub�솬�æ�2��\_E�u��㽯������+�i�5)�:u;��ڻ|)J�"�K��Z�g�@�}2c9�H�:����:%Mт*��\6�0���Hqt�K�;u��x��68Vک�Y���&�K�k"����M�����'q�ݛ4S �L�p�+"�{��aٍt��$h�J Wnf�ʾv���%Y(�՗AБ� *��Y����ۜhsq�����vdv��q�ia�qfG7Xέ"-��B�-Ŋ
�:��n7|���i���;k�fl٧����+0���k�ÙA�w2G���z�s�vv�dEK�/"K,c��i��!L�)�u�f�%����Oe��83����߳�	˷��T����7 ����Y�K�s��p��Nd�Mt��Osw�*��W���ZGm�}��uZ#�)��T���e�B�@rc����s�S�D��`�@���Sw#��d�ݮ[۝��g��\����Z�t�������3�+�ւ�%��q-[�u����1��t�8�H��Ke�h�e�"�g{�j�-�^�)ס�&:�Y��d���)�H��� ;��jd�jV7)�\2]
�j��7W�-��z��9����]���� ���5.��u۝���	<���v{q���Dwd��09��ˮھ;� +ҋt.�*�X��7ϰ�p�u2A|[#j�)`Ž���P��T���Ď^�*��WaL��:W���
���,eL��ˮ{��K{����9��M�)��=�4I�,���;���91�L��QV��^�k8w.;:��.[���Y�i}�*�tP�@�M���3q�	r�d�Ĵ�;�=.��b�5D���R���T���5�k�©R�N[PV���vZ�hk�X��we.�o������n��3�9�O��w���r�q�rF��J��r��$�5B����8�y*��޼��m�M�&�������#�$ua���d��i�u�2���v\F͞�kk��)=L>�T���TisMT�{�˷A�T�L�ngr�nU��ḩ��"S���N�=e���m���Y@o���+Lk8*+xrM���Э8��
b�*��6v^k�����o����;��W]s�O�[��<@>'^7c_\�Rx}��+5==a�j[�s,%C��e`���r����n/z$�+�������6�f�<����7�Rd�np=���ZC�(ǷX*X��7h�La��#s6�Տoy��+�V[���{i�4�heNC�p[��Ji�O��X��|v���;�"��A�o�PL��"ϙ�uL��ԍ��{�F��i2*���P�Dz�
�9A�mf��r�-��	�t��MP�4�4P[$I@V��֔��m��4��4�CC�H�4rMR:�!B�-m��A�E���"�֓ZF���	KF�T���i4ևi(M4���ES@u.���'Hh6�Ԏb��P��MQUL�襠�JJ�P�M�*�IȠ�
5��#AF��(��T����ih
 �
@�M�
C�A��'�uJ���h�����i
���W��:��$v���

�����I�
J �����{����^����*������Ht��邊���^H8���w��_N�҃������P=�]`g_�6F�	x���U�w�.�/=ӫ�-U����x!f,-� Eǧ�U��y��%6�2�&˦\'�V��TO1���$�`��۸��N��
n=�fiG/Z�Q���$\�й�S���_�,��֝�h����FE9��q�������,P�i5�F�5���Ξ@��x􌁒Ivl��L�]\�J�ⵕ�ќy��G��\�j�MlO-��E1�
T���s�O�p�G��3[*S�T�W6�N���,:�1]RC*�,�HY*wJ����'+=�"�-�Ú�F��}imf:Ňc�3ݧ(7p\��t!2��!�:-����[����-?,	����Ud1
�*2��j|��8Å\�F�Wʥph,P{>ȗq&����w��};�eB��Q�K
�%/ѭ�������y!��R1�D�!6�B<�Ժ�X�(���7��_������X�v{�yzd4�6�~�+�%T�>��H���:"t'�~�qv��Dd}+�&4�����:M�O~�2]M�x�X�=˧��h�j��z�;t���8���"�7�F�z�G'�����)\Xt�B9Ւ���d�>SP�9V��S�Bic�tn��Ȏ�=nJ�J�)\�*�;u��P�.�
3��}��W(*C�}N�r6�Z�X�uҀ�*�˼��D��{8K�{�����<����DVR�Q�ݢ��PL���TޣϗzNs����Mç4!��߃�٤��h����8wSZt�HXj
�ۧ&��D6S���P�*ge�9��&>��5����'s�E3Eڽ�]�O��8�tF�Zʷ�Z2v�Fn2�o)��uФ�`B��yw�����O���/,�4�����dk1���8Z�Yf���]���sV���l�w����B1���E��W>��y�X�ou�ęڊ8�4�����n02$γ�l�/!Er�j��,lO�w)��������>�D�S��r�j ��I���������ʻ�$�w:µ;VnUB����~U.R��ra�!��W������ɂ�v^Fu�VL.~wA�>�b��Z�R�*�
jrq��.[�=�y,GG�mtz�k������`�1�����Y���-�A�$��%9(ȤB�I�ߣf�L���c��j�̕��cF �[�$!��r��ق_C1��]�oR���LU�H�����7]=�蹊G�o8v��hC�4%�PFyѢ<dZ���Ѫ��YU�N�,Ԥ�>M\�j�9y���_�s�YPe�w����2�!�pp�j����ݞ�pį-޾)���N�t��"��߰�8M��߼U�t�G��ڙ���R
Ԥ���[�fc�6�Y9o9���H���L���Xt9M��%7�^�㲿�U~qi��Ό�,��	��HI���y�pee}�4��MO�f;:k��l
s؃��Fڬfz9o�����X:��Pi�kS�ӧ{r`��	����6�M�qz����c��B�\�9�,��n+GE���c$R�`��>�|�A��������l����=��Y	���M���Z��V8�eҵ����Q�%m	֮{�t��)媗EF�0���X �!fHط�Ϝ?s�N�T3�v�a�@J��]�K�E�MKs=up�F�n�+����ܴ#�k�)��}à(�D��z�]�7,�#Qa\bK���4$;QB��Kvmvi��V�����9�Q�r,�U�)O萄@��ay�>�c#�,�qP�F�L!�ʧq���wj<W�H�A)��&a�l�oh�̀�����\>d$�{����$Ii۳v�*s��'��<5ǌߣ�)/�CO��8S��.=k�9���I^H�\TX�k/����;����{Q�F��R��)���A�yfP�a*<���ӌ&�*���>�E����Xz�n?pԠ��E��cu���u��cHr��چ�k������$�_#v�����"���1q���`�tݵ"�㜃*	�ή�W4�x��9��u�{cCכN=�+D��o(�rV�vM�S���6qk���w�$���n>��㺝�����C�N�峌���s����i�<�Be@Z4)=�����eb��돈e<�{�z+s=�k��V�Ѳ�~@Ŵ��P|����_W�i�y���ˁx���Ftݢ���G���al�y"�=>�<�U�% �<{������7�>�5�]=۷j��^.2汎�uk�G��c�]ctS�J�
�|ᮢ���H0͓��s�����f:�z���$�7x�f�hB�\�u�QI�Ԣ��Θm&:��0m{p��t�kw��%�µ��15����ʆ�F���������Z�O�Sy�����&k��<���q�5�9G�FgnԼ��d���\D�vk�\�&��'(]�Ta�d��Jb\�@�0���7s��N\Uki�m���Bn���H`c����6%�l��V�V0�е�(%��f&��6���F�����)]ܬ��'uQ9� �À�p��D#��>z��3l�8��WRb�\�$v�$�Y�|�ܡ�b�F}6�Dsh=��K�gm܀������ڦ�����ɀ~�5,���=˗���3��f}����U�MfVШu���P1K�r��~}���o�v��L�m3�8ӂ���uzG\%�cz�j�CF=ǽ
:,�M"���Mr�%�4D՜jt��4=���t1��C36z��{��Zv����o�������!uZ~�1�!��;(�:"ص{�C��z9a����y{P��1���wo;��u������3�X�OA!��Z8�v��,�z�G��W��ߪy���v��j��ihS����t&v�)�L^=�ޡ�9�i�i�t��r8c�Ԃ���|�*Q�T���R�#����*yg��-(M"22�ؚ�O=�E�.J�����E�-{�t*Ϫ�r[7ѫUc�Ǟ���*Uj|�RQ��b��S�\},WUx��?{��M�E5=���Rl�V53�a���f����ݟ_k�yU���Z�P8tH��an���2�A�F��""�ե������L��9��E�f�\�I��7�5er�V�}#`zz'Q>�^K��W+%�I��Ap���I��xN�����E1)Jjn�<��ȸu��֬����\�fr�'h����3K(*Y���A�a�`��%C��I>9�NVy�-�Ú�FN����rk5���k�W�E0���?M����YӍE��T�M[M��Ԣ���'�K��7K�-�ت�R�t���9�G�4e�lSϝ3�]�������׀*(u�L1��k�ۮj`�� �n PU�i�.�J�iJ�Ocbz	�v�*�G0��z��z�ݖi�/&>����R��.��^�X��Q^U�}�Ws؞3�H��S���w6��7��n��ݳL'��a�y>��r@|�e�Q-�3�k]�^,�bێ}lc������"_z�p��9�> �bR1�D}� 9.�vOƧ�W:�&E1T�����Ւ���m]��<��a�\�#�M)�S,�Y�9# ��Й��"7�}�Z�me�_Xuު��*0�A�n�t��{pеaԦ@�k,{�.�W[z�_pW��:�;w;��~h��cy�/���Z�opI>�C�:�]���A��I��23L+�Zeb���rŨ0zM��=OO]L��Ϙ�D����8�s�5�f��U�Nf�{�.^U@�fx�o� 
d�{3?sQ�t����.�J��C@�q�10S���s�oO�^Y�i��y�)]�mp���.�\b���Rkk5Q�xfd�gƚf)F��Ixj_p�
��e[�����z/�>���c/�q_{_�Mwoj�:�O-bVI@$gY��>=@O�Y\�5I@����R!{ʈ�}Q*���wz�Ǣ-GcgKj�-'����V50�~k��A���&5亵��c��*.3�q�6y3����[LҮ�����܂�.�A1�0�Т��g��6P�N���J�쮎�)��:�7N>�IA�ή���,��lknPt1�}�üֻy�L���m0F�ZK��M�3]��<������-��B��-�z�Pܦk�^-��V�뜞z��H�m���.��v]ɷ&?>ze�Юa:���(R�KjܜjꋇWl��'&!�flbt�z+y�rvt:���<������OV[�����I��L�0
4-Z�I��QV8�Y���l�^u>��R��8Я�[��#��0t��},�4��.�ҥ2�n4�z;(^n����柫�4�T��\��w F ��P�!9�2O��2���/����1��1i0�si򆙶%��̎Ƥeɦ�e5������b�sׄ�Rr��ISW�wC�=��r�sGvdv�{$�j{R����/6T�4ڂ'�$L�^D�ƌ�B���������C����/%ʓ�,ۙ8���Ui/���uՄH�t��AG؁��b��a�qO~�K#}���작͹�E.�c��˥kߊ�^�Ĩ����\�q�R;���K͢'���f ����zvW��k:�j�Ԩ�.�װ�i�"�b�E�j�1�&���\�����V��,���Pg86D�Ơ�`�"��N��J=ˡ�%�ܢ����ɞ҄k&�U0�|��`n* 3����ףHq�Ŗ��*Zo�e�f�y ��s��J�er�z�b��i!�Ib�-��FRY]F�G/�,��YJi�OH|�#N���Fy�8gۀ��Y����s��PWl�S����S�A]�5(�k ��
�C��ak��]����0��k;�v�4˶��3.�C����8�(6���"��#.q�\Lf������*��Ef����tb5����� �C$�hzlǊxb@�����Yv�w��7��v,��WgNd>,�Bj-=�k�U�!��G=y,��#>m �	�t�f29�2�qP��}�۳�I��E�!�=�Ix���ܪ�Ơ���A��B����7�t��Q�#r�s(m�ںS��.��S<[F	��#�]���Kfa��?)�	�.�%�fi����kwv_wvp���*ʭA�VQ�dr�z�>		��x��Q͡�	Lż�ס�V�oP�CO<��p�x^Ҙ�EP�Ȼ`�g��y(������5��� Y���2lK<mQi4��o/*3=���%�u���l�ҕ&��)���k@.�z"�Nv����Z�},�1A`�&��w�Y�N�XF�Y�Ƽ��u��i��8��Y=
`-�үr��*�{K4���huHL��r�y���'qUeWC�b�N[�,h.��Iĸy�z;��&X��ܚe9����:�2K���+i1��ifm\To9,s3bc�u�':�|]��ty��L�g*'{���S71Q���K�V-��&���{��Ht|��\����e
���ܙ�v�Ln��8��*�څ��g,�EG|Xff�f
V>��V�U�u��9��z��6���T'f��1Ln�.��0�-Gs����s�F��R��U�S��X^��.�Ä�`����k�zvi�\��V�V0�]+��$[�׻dvg�u]��u�
<�Р}�ʊ��]�~Dk�v�L3n=ޛe��0v'p���,��"�7�5 �>XF}8��fy��,ƾذQ�` �c`,�#�W�h��7T�q��s��i�f�fSfx�[�҃�݊�~ZF	��߄#�BT8-"6��6�1�Yyj�nM�x�D��W�1���q��۬a �C��G(��_bS	��������K���sK�׈�im	�`��I���x�w�knnf�vu�%��qR�Äg��6��=���oo��:�>?�p��,�K��0�Dde9��G>^��P\�3u���
��ҁj�X�uA�/=۪�[n�Hu�>�CʭGPE%�0,.�".>�(uV0J���#m�̃�ʵ��MwOpX����U��O~�gXP=�Bޭ�[� �f�q ����J��9AE	a����i�Ң\�]��z�b�N��p��n�`2S�J�<Su���R��D��8�����Wa�ፊ7Қ{�a�u���-�WsMuʽ��1}�1�|�V�2�N,d�m��1Y޾�;�O)	*;1���bo7G>yB�ޭ����ڃ��u�~���{U�l���4�3�ƃVW)�)����N-��c��Ι�G��i�`h^�H�����yN��9%9��)��'�>��g<�?�14��KO!��y���y��!f�RC*�,���Ď�T���'+<�T�a͒��X���Ӱ%f��Q]�*��|�>O�E�@��Bkz5�7hΛj/xT�[&���Qi��M��e2�/�f/q�Y��я286�6ڡ:�Hւ��#d��i�s��,��O\�u�*־ʥB*��˝�7]�F�wr<�An�����c��f�5�Ǌ"8d$&��<�Ժ�'������uZ��g'E��{Ҫ��j����FM�ʏ)�f��ͳ�����p����͒ �)����;q��΄�:�O��BՇR�u��tzw����w(�|��G_܅�%~)�
�>�fe����1x��أ��u�2��D��gh�@�[8�@��(�Ys�*{�=v�Ͱ��PT|<!3�x��؝������ �u����|wֻ�������}?/����}��}��~�ޕ#�� �sU�hZ4���N�.�WW�2��YH'��R�H���m���%��-� U�;�7
F�с����!�n�k��6vy]�X@G�·F�������bDtNaYw%��/}��.:烀�]rl�����i�n�b�F!�4㻉-6�ܧ��R�3�h��M��e c��ڛ�V��l��P�5۩D�;̮�(
���k-����B��3Oe�u�4���B���A��W]�.��Ԓ��G���'R��w��ͬ\/u���ǭ��`��)�]lx��R�x�r��,{�WQ@;4���Q[�k�0����p	����5ʂ�9�7)Q&.����bG�nX5�5�C����gm���:�[�7+quZ:i�7�݈GRT*4�ʳ�䉛��Ho7QucZk.XW�4(�w���;=1���Z�7}����$�o+��a��� yj-��M"��kS����l��]��ق�!r�]�3ez̵#r��l	!j��Ժ��R&�7fhSK�oG��#��t�hh��fu���9Q�"�d��%�=��S>4au����v���� D��ϙ8�7���wn!v�2�Z��؋�a�X>Y�Xn/nQ�n��(� �o+�[;��R�V���7�7���������ڀU�y�3lh�b�����j�J�����kJ����s���,��f�> ���#5�����K��-�z=Cp�1k���Ƨ���EN�63�
v	V�{� �\m�,42A�u��"�XdIQ�H�m�����ۆ���z�����K$�ɯ��"��8��NAtw5e�eT�H��t�5neֆ�sŨ*�d�rnaV�W�g]�ӂ�V
�y=�.N���7� 	Չ�2V��׮�� �t5�q�����u���X�!y3cK����뜬���M���Zi��6���XR[0Z��OnPz�9sM]��#̬�R;;�N��c�L��'�`{�]:�n����=�5��ëw$��ɝkh��l�V���f�6�1q��M�E�٘ve����K�&��]rn]����A��]^n'�*O�������Yy*�|�~i+T�t�J�e��i;תm;�t�ol`�.渍�݄������b ���Y#������2�^�h�5'8w^u�7�wC@(�,m\�q�s0N�\��ٽ$HJ��ǈL�{��J?��_�%�ܥ��!�#�EWR�#��8�r��q}/s;���*!ٹ�v�9���=Y%'I��gSZ \i΁Ҍ���jt@��͸�V�]�"�P�S�>�2��nm$GJ��z�:�L���b̦^�[�v@3c��r�M��,z��qx�j��X*�� ���a�^�@���]e�:����>`�cu�'�����p7��YR���5�K8�w1l��} 7��,A�35t�H��^��Z���z�U���u�D�m�s7p����r�|{�Ǯ��]u�:��O�t�g`�%�)�d�B���i�Jf)�*��
�tPi
�t�X���@h*��3BS�4�-�UҔĳPևF�%!K@R�76������N%4�������TMDE Pr4�U��
th(i����b���j&*]�("
N�9v��M,Z$��Ɗ
i(*�ꂛm[j$������ *���)i����@h
*���F�����d�A<�D76�"��IKMU%V�ADKT��uM,�DDCClb��"4��H��bZAZj"Z�T1 P�S�֫��CAQQ3�|ow� l� �nGL%��޻�ζ~�O��{��#*ɦ@֫Y�TEB���ɚ�k�����#O[�ʹ��R��0�"�y	S��%$�H�IF�H��+�9���x{�^��C��E��mGW�"R��8-3q0���N6ۜޟE�f�E�)�n�E@Z���{#��Y���C�{�DmC�r���m�IG�����x�j�j��7_`����2k���˷�V2�����&*� ��g��8ɽ�)�?k�<H���[J�ɷ�QTo�+)���J�{`�rA7����O��vPOk`K.@t�>��|jʋ�5p�e髄�͢�o��FҮ`̅�x��ħi]:ɫ�0���A���.&��.���R��KonN5D'מh�ܪq�Os��G����
�KG��/�����"�:�N��Й'b���4-��si��j���9�_��t��6�NE�.�o@A���6`�U},�4�v��T�@I��Z"�҇7;�kN&��C�4��.͔���n@���"�����Yb �%ےJ��-��%���l����m�E8�=����������C)�Ax�<à�ΥwNv�TճH�\�"�N��rg.�����\���j��IcH�N��D��؎�G�*υ��:p��R��l��L�ǀ8;T��R9�`v(��)K�A����k}�RSG�z��x��#:���U��4I��4FÛ����W������6�JJ�2VVk���\�@��&��K&\̬35�/�>��S6�2׀×H��a䫩Y���3w�Ug�rO�Fw�~��Yc׺���r��d�@�⨑@_9gf��WAa���ݖ��#a�W>��1������,�OH��ƅ���k����k�*	{k�9�����ec2�~�iaP2��|L��y��lsL��e�mf�XsJA,�k]CqM�n�S�y��g�U��b��z�᡺F��U��[#dJLj(��-���2?~?���E����aR�%�#&No+a\���d	�nנze�N���ej��R�d�R)��3#Z��7j3j���,Ji�E�Y'���;�2� ��e^�xcC`3?�܅OPɁWJ���Vy���
0�OsQx���؏k�� ���; �t����Eǭqp�T8��r�~�J�Ω�W1D<�"{P��Z�V�R��ܤ.s��"�(Q)��ӻi��6w��>v�ϥ�¦*WE3��Ali�	��#��l�%�0����m	�e%���,�lr����Zn���B��α�3j�+(ƌ�3�!:�`ws�;�/7����<FC\҉���+6��$$��~��8�0,"�1��.��11|^����k��Y�#�f�i���tv�.<����&s�]xx]��We?�q��=	�|*�Tf� �u�ǉ��1�훒-ө>�'j�RV��ɥ�z�+$ã�X����챼��;{��m��N�_���5EP�R�ku�1U�%Bc�Y�p���M<;�Tx�1��%��j����{�«��)�1�d�ctSIRaA׌�qa�&1�k>��0̈́OIjPno�7<�,0�k�b��$ŚN�f):aa�]s<�妢S��i��χe���ֹ��Z����e��64��t�,ta�la��*���z����,V�C�3��k����s����#�z���4�YUt~_�ޝ��'f������a9B��0�Z��3�X��.�b6eepy��z��~Bme���T�� ���<!��"s[B\�vߧ����*��a�	��ƕ}،��)'�xH7��e��ݵ�C�BdʰPa�P4C�0�.>�Nyu׭�Z�w �^kK���W�������O����w%���������`>�E���'�d��m�#*Ν���:��N�۲�}}$�Xc�C�gd���lZ��#��R5`�}�ӝ��V�.Dw�s��J�׹��t��r}�X�}�	Ŝ�z����o���FGZ�}�@������ZH���d1�8�ᦈŲ���ޣ���;��n�<�+��ڞ��s�W������GZ��uZ�G#6p�;Y�{GmVX#��u
ʝj�4�!�s����}E���!Y��C����v������0>�J���N�ݚ���G�}�0��r?�!�6?�F4��2O�=�OBz/��C�}�����d�A,��uc�f���"C_�zJ�o;�öm��6��)*�fN�\2�,������j�?w����6��baVj�Suڸ4����	;A�f�'�1��@�{���<�r���d��Z��	wm����
�!��s�����^@�	M�R�&�h�'�J3�=��[�z��A@�"X]��y��VQ=}�r����9�E�N�~��O���,P���ie�,�\��T�ۋ#73������w{P�6$�1��`���<���'�1)��t�cE*Mmq�<��. �F6�'�n���F�Ő���@N�mB
�m�6���'%C�ԩ'�1I��%�+��?>���ު���Kdќ����찋a�9�a�6ཞj/�C������?"G	��C�<�bS�G7f�:\^GW�M0�@~�l�Q��G8�U��e��;��u�è}��5��������V�kz*;��㿇O�K�.X���Wxw��{����D�İU��1��y�a�U��kdq�[�/:C]r�9k8)'��1yw�;'��F3lW��5�vc��O�����/_�J��o�__�ދ�����<��ч�C �X�#���׽%*p�NW0�'����Fb�F��n���8�l�j)U�8]w:h���9V�e���r��ƺUc]�L���o7J|�!�,l=�3l�0g!���u��e$����9�9�D��P���}B�����e�~�}]f�����%����T���y���L�𣺘2A����Ƒ͜�V˗����{$��#4¸��&+����7y�N�\�f�y�Ղ���}�
��ZT.��9#u��79���'��}��z#D"BȾ�j�o9=�$$f�T�ڎ��%.#8.9��0����s�z|ҍ�4�c��l������h�v&iK'{�a)ư�9v�^7ʃSj6�H��xl	��!\Y�U���^u0�/t��7�;������j�zY㐃&��HjHγ�͜e^��t���B���s��^�)-�&���ui�D܂r^m�.��t��U�?߹�>=�D}����U����q����!��(}�$��bS�uzu�n�+z�k��'V�P�
S�"��`�,���h܉�ܓl�.���\c<H�ހ�K5�i���^�7	�����	�{bS����aِ�(jѹ[���Z��{&%�8>���e�T?���D��]ﲚ:2G/;)�B�v��	��k�cF�����`�B=����E���i���s2S���:�Y�b
˛9�MJt�u�*�^|h<�2"���F-�uf�IYJ�dxo29��/כHU�z\fFM��zhX:q� ��vH8ݘ!��f!��˶�eD�/�r��~gso�nM�a�E(���/^�����<B1���@OH �����ΫNr�=�[qS��U)<�=��T{����T�)�AY�v������_]'���:b^V�u����u�Iц�
�Y��V�Qy�T�4���%����/*�x}�EriMh�z�K�6H�Ǟ���W'(Y��N8�U�9��J�����l��{�s��0Ry��l5�9��`�P`飞t���m��Bպ��:�-�R��pK�2�l���"?5��NkVt��V�7�ׄ�*�'.1��̈ܶ��[�%�7�P;�Uˍu�޾�Tcy�kZ<�uIk�_k��T�n���F�P0GR�N=�.�3��aغ&,�,��;=���]�Xqx.�8˷c�3(���+T��8���@�Fr�wMˬ�����Qό]�nY�L�=yC�x�Cג��O#.��,�m�{ ��ϗˡ��P��X=ށ��t�ֿA�����հ:�֕�;���;�p��
t;f��`����n��?p��mN��+��w�|�v�n�2G�U�fYr�TNv�t�P�}�{Fr�m��+��˙S��0�)���c�֗$�.�k.��ll��J4rp��S�����[X͊i��yj�9Ҹo#^i��t���b������|�����%�h��,:N$Eǭ���F5u�T�5.R=��P2�������PqQ��gw�k�4(S�-�MV
�}K��ײ��?#K�u�^ߥkv8>�/�_�w9Oخ�ϬcQ��ж.��sR��s٣�.�Nk�=[�H��v�1m!8��S!"��Ch�NvZ���S[%�\��؀ܡ�|�%��ħVT�	�T.�#'1����	���0������dn�:�ӗf3a\i��.�3���JN�xd�ktSIRaO�m

�c�b�G��]��>Ete�ط3���#�z�C_z����<����@��܋6��ALd�z�n97p{�C���׈j�Ho��xy��F���.�0�f-?1NXᵏM��*w�-�_횃�t>��KwD�O~��<���֘��]l���a9^~�öSYUO��sYS�%`�&�T��pwC�����5R
-�s�����j��-l���
-��<�a���9��F���+�<�$ww:�=)]l7��Liu9�:����hD&E�9#���Mܤ_�^O%_�q���s�a�Ѯrq�WWP��雝�tH�t�1v�P�I�B�E����.ήC��o�O|h)����7��IJX]3%	r�R��jγ�X
�$S��[Wn��ì����I/��)Ai>��m�Y	��!a���D=S�#����|v�������ˮmL�]n�W�J����@�>�z&{��GrY����A����U^W�v���V�3��"W,\!M.�	�\���s������OJ�v+�����v!��=���DTzr|�6�2�9p/ڱ�X@��=��M)��9�	@��Úz��4���ň��Zv��9LNθ���b�s�BB���a��Y�6���7���"$m��1K#..��HY�����g'���J����0~�yc��J�ɡ��{����\���;t��z��6�+��d�Ԏ��0�W���+�qc�ܱ���UP���\g�Y�؞ճ
A�����I��Q���=�[�?W�vO�%�u���9�Y�1+a�چ\���X�+(�*�q�|����,�<�D4�Sb�̴��R�pǧ���Tk�%@g�0vuf��k�c�t�a�Tk%�!��or�g���σo������P1�L�w�2�xi���{{B���?,3yY����~�k��d:�ʬ7s�fkͨ�{oeh6-�ƧL�EhE����6���ŝK�+�Өg΃`��)���+kB�oKOR���Yzc��ʲ@�nj���'�.���"���S�m��$��W�Ym>n�m��9u�ww���]^=�Cf>�m�B�˲�8lxV��ɢ�٪��ͽF�؇û��Cw+Oܷ�w�eO�7@agе܍鍕Ʉ�z���!8���$̎ڞ#��W��#j���+��L0p;ްú[�n��9��]S�*�����$��ɦ�����ݞ���T����X5jg�}{�a���ݡ���;����n��)�Z�����5�GI���Cu3Q��vYNhk�X���]n��}�[dz�<B����\�W��S��/g���'w���4@�g���`F xV_�Gp�7�fi}�q���C}�R���ה���h:(��"��dd3�b4_@xH�u�i�A&�Ә����*�~o�[��;������Z��s#e�B�y��n]Y�f�F����D[ՂR
���>�1�
��4<��v��N�6C��i
���y��n]��jN�![ �����EK m�E:�w���F�"ɲ��З:�G3;���xJ�z惓)��Oc@���.�L̝�G��畛9'7�[ߎ/��yHg���3q��J�%.ƛ�R-[���d�;q�KV5nUOl�n���E�w*�l���\B��	���i=w5'_�6zyZ�w��g�����~�WIG�R\�7u�V���G�z���gMV���MOt����~���j�2A�u"���\���֎�s�JK�g'M�����݉�������T)H�RfD�2�/`�����/�����:�3���s�Ѽ�g�sm�E[s�%���6�.�!��y�LS>F����E��x4/K�_
oH��5d�Q����K�󮐷�g�g���aPvpK_^�m�ƈ���Ҽ��t�BOU�@UY\������ǱԨg�E�ەtӶ�������n,:��ǝU�<�A�4���ʅ�<O��U�֯P�H�^�xk�(��6�:�����4���4�:W�j�������}>_O����}���������N{����w֯gf�t���$;�M �#�U;�_�93��"�䆇��&�1J\5�S�Z�:;jV\��)-:��0�JS�4�Q�X�m�c�r��oV����w�n��]���M��Yd`���ĦT7׉�d����z�1#JG�i�� V��o�G�Hd޽���p�c3���{�V��.ֹ̥oR-I���>�[&�Y@�wu>d���|fj����%�n��Ո˺�Q$ayy¸��u���u5�Baz/�RUw	���t�U1&�����6�CIR����ֱ��Q�o���Ϻ���V 	����/��Wu������N���ʱ#�fwp�6�{���T.��T�ظ����JwǳA<z\��"�b㨀��:-�rKp�S���ٞ}�����u(�!�@�=�q�ٗ0LwE�{��*�k��Do-L$nR�+5;��|���Kn��8�"�u�Gէ��!vt��`P�澊���;Ư��B�p���t4������6z��&��qv�P�꒗ )�ՔQ�\"E�7�%�x
�+m>�����]��k�sFPBL�\�G��`��r�zR���]\]p��G]w4����P�Y��ɮ��%�Ri꓇W#��UwX{1.�[*�x;o�M��qn�8-���֦�Oi�B�'E��z1����겞�4�X��4�����M=�*�jg6��T5��4�[������PO%A�Aq���i�G�T��*�(���г����k���e-��gK�2>�y��rS�Cc�S�f9K�Ҹ������\3 wvڦ�_h��,���3�L��lwu�-�F�Dt�CQ,A��6������aomBN��?_>W��N�#�S�],:2��;=�>6<lB|�Z�^�V`qt�Oa�Z�t��N����2�8�Ū�X%�Z���s+6
�j�0�F
�FiSV�p-G�v�M�:Q^V=�y@w��"S��Z&�c9f�B�{v+x��`��)�"2Qg\:��l���N)�kf�4J�8Y��m*8C�E�Ā9;=}V�"wݘz�ͨ�!L8����u��t(+ץ;�R��A1�Vi�}�f��F�8����#9���k��3aU����;r��O��4�ߺE�W�K6��B�\�-�]3�oP|��xQ�݅�d*PrI�7/����ޫ:
Gzl1��C��+�f&�bՍ�>�Z�)a��̀j�g\k<4f������u9*��M�>�ңW2����a��4�ld�k��c�@��6�4�̭V���6�����\���˸^��W8�Sz>��hPTm�r���������6�l˧4����%L��mna�Y:嬮���D�V]��Ì�i��~r�Vf�n�f�Y��:aG	B�)���t��*e�����!Y���3�wvM��*1p�I�_� xh{�M%�QT�E%1	��D��P�LD�)HS��j��j��QP^�L�g�NQPD�͂��j��ӪZ(���8�*��Zb�L,ABiSت
"
Ӣ$hj���$)j�"��4QT֝)LMAMP��F�Vڊ**Y�:H�bhb��"j
���b�9Մ�Qm%RQHRU%4�Q@P��qRU%TEAJrt�QQ:44�mF�)MAP��Z�)�B�h4:�Z)i�\��&�*��9��������j��&�a���*hz1�4,sb*���)����a� ���)��Ħ��7-A�̅RQTSUr�T��Q��UMl��%�(�Jh���AUDQ3]mEDLUE�	5@S$UOkY��t��Jڃw6I���:If�a�2��j�l�������Pf�݄�[���̹��.��1���ѽ��0WlRe���(���=���4���G3�!�q����E��\(jX�N[����E̼�R1şi}Ͻ��������x�省�<u�/��6`��C�����7�x��-�>&�Oi�=�t"�G�m9����?p�/U7���tydD�$HI!#�c�W<������	��#Me�N���{�hD��^nǯ/ȉ��:|����@����S�ú��D w��6^_���U5�����v��.�I*���m�6g����.�þ�m��|�SsN�e݂
����n%�1�51�MGF�ח7]�40�m��}ط��*�Rn��o.%��U��mdx�!����+LYw����5�H���q	Pn�k�y2aL��ʭ�u�U��8q��s�י<%�2����L��-:Efy�M�)Ғ�D6�J�?_Hk�@g��ݕ�ߑ87ܐ;�G�[���c�m���Y�a�b�^��]���M�ui���&M[�0=�X�C�-)4St�]�V8A��)X�5ղ�.�c�r�'e�ǭ�39>*��ڐ�<Lm���L"�d�����ǩ�����p��Q���ͼ5xS��� N�O>�+(���y"ȅE6z�IV�"�sɐ��7Z�iX�j㶯�n���̚�0�@�d���p�zN�M2(�zR�d+P����b�vO�P����$������a}��7�ѲU�'	���F�k_�@��W�rI���7�k~���n��?�ކ�p����ڃ'�D�缫���}��oԻ������X����ɿ�����C�"������Nۼ��f)�y^���p����֕�	���	��c�R��j1,��\`�s54Y�E��	g7��df&��{��I8�d�c��E��&A����Y�{���A��6��xVj6�-���#����ֹ�(�3=v�n�:)��u��vB͇�J�u����Dt_.-r�T��ݘ�,�w^��(i��vz�R6)����A,����ӝ��Dk��wl�ӷn����dU�Xcj�&��Bv��ve3��uv�jQ���B��E$"�B�e���&m��[��
����K�f؇�R���X1o����IC��djX]b35g�n�YG�D�}7�Qd�"����`�OEw�WWgmC����)�/��#@�v�@nM�;䎴��R�:�l��t�un�0�/:��k�n�e����K�ʲcg���PT���|{2E�9��ـ�VK��Tc&Nng��Z����P�p�jh�(׊2�B�T.*��j���H���G�?/,ht����U�#o�N�$G9�U1Z�LťeGV�UWfs�ݾ��k��s#T-��<��+
m�%)h�]��ױ-�x�{+r�p�WP:o�Y�6c��NBٍ��������x�̢k���������F�+	�����GǛ��,�`����7A73I��]B�i�85�x���g�����f<Wr���a����oa�옅����U��}�`�ncd��$��>җP��QBJ�*����gSö�X�
���Ѧ{������zek���}YC�uu��_�離�(W*�H��?���=���rg�v�,�SBk��WMN�n�8^�\|v�n��d{��WRS��ϵ���}<h�������.hX5�ೆJ.3�y*��3�1;���Ԧe
�vj캝t�u����I({,27�}���Q�	��@Y��9bt�������~d:�s�_m����l���*:������h��Թ�/���M�l��A�t3��p0#���ףsR��܍��`z���u�ٯ�&���/�����<y��7�Ng!� b�0ΐR�vQBJ��K�Sɫ$�	��w���T���=�	]	O4
Yk���]���S��Yl^'j)��ݱѯσi5tlnƅ��RU���ICv���ۡL�9��V^	]��|�ǌ�s����}C�ʨ�&����Z�vM�:�k��t(h���gg5d���Tľ�I��9 `����q�J��,�e�ʾ�wbn+�ky���|R��Q��3A����!A��#իyM���#E��8ف��sQ�-������j��)��{2��>oBBvM�9̝6(m����u>u�!ԉ~'[�E_���N��;!��ϳ# �"mN-hs5p�q�3zG^wh�ٝ��;�6�g��k}�F�CT"����G!�[fN��,�.��b��u\��-Sr��V'^����T��>�Ua�Z&;R��.��*{�[���t��k"f��X鏮G)�31�._<��E���f�~�ߙ��h�Z�q�\��읞�T�������v;m�G?"�X�%��&}f���*�+�iR)wp��t���so��%��9c�u�1-pv��oPٔ��=S�˕Z�0��I��3R6N��q��센ґ���?��oHa��#1�Vr�Ε��׻!�v9ˌx}�f�5U�]��|w���W.��:��o�G3���|�2�fWsx����j���[ze�gm��i�NR����.�����Fi��
��K�ξT��g{y�����ѷ���${�u��;t�<�aK͜��ۛ�}�֪;���:��B2�+â��I�D�$��@8*�����Ix�<�_7�p�l�я���B���f�7cׄ���vB6C��km���{�.j���=\�S��?�w����עc��.V���=�9�OV;���5�9�l��]��1=ҭ��:ͭ��f�����{2��Q�i�8hÓ�b�.[����f��gf�@u�]�[6�T���W�0ŋ��Q�Y�S����̩X'i�.
�e:��s���j��o\�7[܇=}��gkn��K�U9�ܻ�vh�<���נ�s𥸓]NtJ�n�������q���p����Rl���ә��pJɍξ�����3s7α��y�O$;kr
WB4J�%4���|;��[S���`gY��'��.�y:8����D[��Ipc����$�O���e��2�mŮm�e�q�ܖ�w��D*)�������R��.XtN���b���9�{X��dwv�l{!�l ���d��]C;$�M�����K���6[����!�M�־�bC��\_�����_@�~��X����h�#%�QJٳ��f��y���|N��0}ƏG�����0t1
ފ�k��gZ�����R��w�TT�0"�e'����ﴚGAO`�J/1x&3p�f���;�/:���Hn��*(��v���>�j�3�hO��>���q�r��������� ��}*�f�ܞ��p�$��W�-����N�
D~
,�ZXU��^b�޺G5 {��N
�����Xݔ���6w�˭��ޒZ��h�͍��W@т�x�.�ѤQFk�ʁ7��Q�z��ݫ"蜧�V�s�P��d�ּ�}���8�O��k�izM'�v���Z+��{Zi���'��f��9��#MP�<{�h�Ψ�Z(f��_Y��H�.����P�S=����f����f	W�NqڼC;+�?$�).3mf�ˊlTn�M��=�bqrW��Z=WJv)����A	�cTJ�������̪ ��f�p��f3z�vn�:x�5䎴�6��2��P6b[^o]�X�+�]����ң��(d�� �B()��=j��K;4xx_]{�?~Va�rA��\�Q�zW ABj�p�CjW�<�,W���L�k'��p̊�E����y�V?�[���@.�
�Њ�/G���d����<���ym���7�d�I~����+î�N� t�#����@�-})8��u�>;�!���מ�yu�d6cƻ0��󐱧Ѽ8����FN������>L���@`w_5�p�nqGO��"��S�/3J�g�����5�f�!�]��j�*P��[[F2���l.W�p�(VW�E����2���r,���F��)�1FR��A<]��j,C+�����F���{��ì����2���x��J�w7Cp�yt���j���~�1Q19gL�͌J2J�S�|fk�l?��b�
����@e�?+�{9�����_�_;Н�:k�Q�9T4�4�LAJ`[�>[y�N�N+;^����}�/y��P���6y�F}�>�4�������Wf97�xq�����k����=v�A��>�0!t�F�Yl�ò,��s�N<��c�Q���M� %'l��c�!�u�sFU�_$���!1<m)ǽ������њܴ�c�M���C:0_/y�� +]q5xoe��fׯ^_����b�m����H�UI9ʅ=Yo�$��#����񨚺����ԁ� ��Yp�U��i�7��g��Õ�w 9�)g��A*z��7�&�6�-�s�6�ߣ�0����ג9;��6��V4�҇K�8n������f�ӕ�V�0g��_�:���؟��n{»ǕӔӚ,w��5���h�v�nF��'ά��l"j����.wfRػu��[�&k\��D�J���"��I��>d�Kwj�c{�0�wN�v1�
�}�13��`ua܍��{e�+�vީ��g̶�x��͛��}�(�藉j�\�HEof�O9;���u��������L� ���5Ov�)� K�P[h^gP���Z��L=�Gtp�Wt{6	6ܑV��N�Ί�7�����S��Qϱ�R��a�x9"7��|�P����U�W���}�u�k��k0kK7]�m]�����D@>��&��W%5�]R�h%��yn(V�ؙ>&�3�%�_�s�?0�5� �?��}[�̕^�fE�����Cѣ�ª0�oQםPgJ�u�������½�\�6�W�9��Lde�ϳY����	kz;���YǶ���W+�.��A��7ͣ��ޏ8��m�����B�kZ��.f;�����J��"E`]3��v�N6�O��O��%�?%�������Quᵵ�� ��r*K��Q��a�^�x��y�l�t_<�i�C�2�r�tPk!K��ph�)�d�U�w��5����4���}�`|��
�˵�4~�
��v��Y��� �7�XJ4D�%vx����&՘3+O��#�u�1��Fi�)�;��P2h'���GGt]�6	��iTe�6;�E嘓ĉI!#�i��!UÃn��{�{���=GUnO0�2��F�r@B�=%1�uכ�xH��Yݬ�:��T�����w����;�^����{���:E�}ﶿ =�Q��i�w�c"Tv[����_,�:9+�)v4�^Z��s l��
z���pVؑ�m�Y>�K�n���sv'�!ϻH8y$mT��P=yQ/w�VΩ����O��YM�0õ��Wu�'�.�B�aY�Oa��)]���P��ʫ�emS��ƍ�YV�5|�A�l
P�F�<��2����"�;A$�\�F%�ݹ�i-�9��6+�n�y����)�[�!@��3�����Ҹ=��5-4���̝��#36Gm�M�S�p=�fF����4SyO�����?������}>�o������ǎ��en���>���b�ec��jo@�*��*���k�a-�&*��욉a�\��r�Ρ�)�w"zŊ�Ք�
S�,���8��t�^�xi���|c�v����=&]�w�eg�8����{J�;�� u��o%�1z�:)	]���ԁ�Xq�٭�A���i�cu��4UnA�`Jr*vwZ��w�goU�2Z�����a����n�?H't�S�頳�3K
���T���+v�f��v,'�=�T�,�[qY�����HZ��Ĳ����Z
���]��o'\71KU5��Y�kq���p�Vt��q�,��h5ɇ����$�)�Z):�>�#�^����H~ũ�BP7� Iq�9�jXtR�i��$y���^��(�V׶f�gR�LS'8���L�>"��L_Y5_�����vz��
b�g&.��4[�α��q�y�
d;M���d)V��u��*X�Y���ozT�z� <M��o[��}j�q��D�j��vA�{'dv��t*[���}�Ɗ�\K����K�k�5ܾ��˻NgB�R��^Lzel
���>�V9�K)�Ц:���.��5���(R�a�S�Sw������������\�w�B.�I�A�,E�WN�*E7ua�s��%�6u`jt���'��n��P����\��tGC.RR��CJ�W�-�:��,B�&�|)��7��w.�*��t�p��P�@z6��TSHEvjF�qȂ���v�V�d�g�ot���u(]f��g��ƓΆr�3[SNt�.;J�K��0U��Ђ)�zf�r2̭�{�r7�0'�ٻ�1�[�S켿�&��3S\�n�39��"̝��qS�㓶����9��
�wq3�n^<�%� ����<auuY�Cy`v�q�#�$���E��L���܄	+)eCD�;+���!��z�]�ø��F6
a�׼�A�-�t��Sm���\MS�t�*�!���u�Z.�9[���^5�/�Z絜�����!ǈ`;������CB�K�$ɼ]>q����F�%n�t�1�h̥�;%�N2<n������>��{�nu�}�vM�
}��f%ֳ�Hcf��ۭ�)7�Z��J����ʌ�����.�fH�8Wk4%�FJ83�\�f��Z�.!�w]"o���}�ۑ����7����fr��}A�6`|�r��NDM�,�(��굄s�T�30��Xpk7��H��A7h�Dܽ9�����.[�(����p%Fe����^�в�'��u���N�Jzxf�F��u'eh�[�"Y@� ��4�N�p�*���S.�( ��䓥���l�ɛ����s���9�j��eV�9�#$5��u�]�Q��hb�3�N����������������e��̗��f��O�J��{�ξ�wLSMQBQ���h�6q�I@���A\�J��(����Z�(���d����"�f��7�DRE:�1\ɤ��lW#ESTP�T�DP��TPW1u�QE1V�QPSAQ0EDsh(���ۮh����cS1J�U4N��%Q3IQ��:ک���\��Rx�AGP�b`�T<�Q����M%Q$Q1WXɡ0EUMU�Պ�����M��*墘"y�ђ����)��H�f	��*���wQ��������(*i���j��%E^7�f�*"�f
�����gŀ����EEQ��D3SK؊�F&����EQ-ESEu�CU[j��N�b������K��GQ�N�ET��(:٪������?D�"\¥Q�wSS�F�
f��%�U�\�����t��^���-���������c{��ԍ1]���&�EX%��YE�:T)��E'M�6���v�X�t�����?}[��&B��!x:�ap�~g�)��>��¦��T�ұ~���dv�(��)�:$�>6�|i���p�����vyQVr�%Vn�o�Xn�2N��Ύ�@�y.���B���e'��q��NR�����3G�tE�o-�����9u���6�|�r�&8�f,qy9�2)
FQ����.k���+�	�hJ홌e����|�s�C�v[��j�����֧U����Z,�T�����³Q��kn���ON��WM�i4l�/�=+f�!wY^�K�#��W~cU��w������5�\�٭��^�X8�t�p��Z��!<�@t���C`��A�Z6i�(�j��9����k�Rh^��)rBA�ƑK��)+�Q�+-�'2)�oT����P��{�4�&�c{�Y�EI�֨�>��Kj)=o���J�����Vc�s��+��!����ʷ���@y�ypcw�V�����P�����Jʛ@�`��-괁[�e[��(>q��K7�]�-�1��(a�)��wC�K&�\d��#z};�q�L���'j���|�v,uX���ɮ���l{�Hڠ��]�nκ^d�����^i����ݽ�DV��+u"��� ���A֬��5��']"��;5��0�-��}���P)*��Q�u#K�t�dpR����q]��D>_�v^�cb��dƟy��^מ�yq�;��x��t��[�=8��d���մ� �u��7Kg��+��f�`�>�n�Zu�q�m�U����}�C�*Dt�Q��|f�k﨤b�]˱�
<p�e1�q�S�5۹�,��A��Ly<��Vt�4cr��R�[�(IWtͫ�ң�qD�e?�,w�BL3�Ϡ|7�#1�����9+�'՜�"ŗ�$<��n�>*��+'6Gm����a�At��F�Yl�ûyl���e��}���E��oR�&*��-�$�H;f@�c��G6!�W_���v�v%�Uh��'\;W��z��zȼ�@~�R�L��H�ҧb�������CyL��ѧ�s�赵�.�!�4�-V�N�M� �
�%��b��S#b*�V�6$38�����|��ʕ�Ձ��fc�Rn����+N�r��ˎ�Π�;YG�_H�'���<�tQ���C _t>i�}�0�+r�GJ�7O�8��Y��꼲#�D�F�k��q��ͿՆY����Ux��9�Y^�F"�P��TM]P��u N �dI]Z��v�љ~���kin�J���g�[�ae�=T�D��ɋ��-��	ӷ2v�Ÿ�o���1ި���W����ӽp*%��?�
�9��@Yh�;H�M"Y��p����Ci���|A��̗<�N�H駚jР�t��Xi{�{!��,ޖ��x��r)[H��n��˥���@;��d�M-5��nTG]��%�Ev��B�Ҽ�8e��0H�A��F�s�cD˘�ݍ�����˞�dE��s��#�9&G�H�R�YM�)W�J�z�����{w�U���C���>aN�\hG'΁��pY����UVW=)E��7e١/GK\D�2�=�� �OF��y�	�1R�x+7��9z�>�ꖞ���hk5h�/��mm��L"�k��&9���E׹���x^Q+1#Y���������w�)��e��3zsA�n�hd����S�Ҽ7�3����ۉV3O,eH"��[�q���)�o�m!��n�r�n���V�{fJ�i96z��DE�J����=�#�{���LT��]l����n0r7�0�
�|�2�֟��yGI���E��O���ɾӄ�u)��]Cz[�6�goM�b�^`�L�^�qy<�M�<�0��٬�haH�.��E�ѽ��xwd�B�CgTr����Y��
b0򘕗@F1R3;ͳ|�W#�ua0b��e��N�e����������u��_K³Q�����tz��I�D���]�NMD4=}�Pz��۬O
���"�^@B�RV.}�//�ۻ�
�J\��ݚ������w��>�NU�Oל��7삅�q����v��re���X;ws�����*���yjE�9�l��N]��^K�
�S���?_:��J���+�IU�*��r��й�2*�~���~'=V=S`�2�F�/�Q�N�����s��k^���d�����u�c��]���q�ϖ�l�����z�$�o8s��]Smú���0��R�6;����%d#�0^V�ɚ6!�:�Q��S�2���x����ݤ����Sb^e&���E��w���E"}غ[�K�y'IK]U>rYL���٣33��[W��t������[�z)�#^[=w��;:�S��둻�>�KϹ���S8�]�.�gx)B�E6t��2xW�E�y��J�n]�y�mtv�m�M�R�`�GM�u҆�W;�����ʃ���g��V�S�]��J���9��a}��~�C��{w��t�hsӭm�z��ʡ�W��tϭv�l���USi�Lq��^o�pd��W1ғ�~�O%�Q5)�L�e'�j���Gz	��M�u��r���{�X�-�n��N��q��a�������r{\>0��A�13�΂0�fDc,�-�|�Pc�xgv*luy������Юs���~��ڞ���5���Gt{5�#.%b���٭�:�SƬ/����u���I�̷e����4^m��,�._1yӷ�r�6�����>\w��
���:��D���k»se����@I��LT�ۧ��s�dT8�����c��2��r��=}��૽'�o�gv���Cc$�k	�E��7<V�:Ͻ���f*�c�~��A��_3��k����́*/c*8j�y��y�舟gr�K�ȴ
�R6)�䳁c��lt�~-m�'�����O��u�&�{+��
�B��m�GZFm��e�q�S5�����2���om1�����r�V%���BĊ
E(2OZ���<ҋ��]_n𽅹�EM?P�:�P�s�ڧ�g]�r�j�>p�Tk�~�7Gl����nH��??U�)ȩ�hEW�G�\+.���GO������m����RWL�=�N��.� dpY*�S��w��;�i�s�"��e0��ܸ���O.�'����� �Ü�s5�ꚵ�2�t�sL͋�"����\[�%<�iA>��|��R;���z�f�����4���ѳ�^���3\���F+�w.�����QsP�"���֩?
�֩����9X����N�+P�YY+����1-�q_ll;q�ᝣò����8N�����b*rXT�B���Bn88&AS>}H�oF�9�)	����mkO�Oan�`4���x��Z�jvk�u�Wr.6�Mo��Ǹ�.���ߘ}���О�Tgh�79�)���v6V�S38����̃����Hԅ#��8�3P��	��ze[��7{C����OT������#�yR��;cg�7w��B�~�h����㿅�U�oqw{uD��xr�#}����X��d
1�v�Hc}��F��\	��;`���]�z3Z%^�t��1�w����c�O_���6�6�QS6r��K�9��m�K0���ĉ�Di��-e'|蒖O[�؈ؼm��oc�R��h�M]P�;+R� �Q�CL̮��0'zr�=���U��ª8;�3�����g�_����x��2b�.Kn�L�9�Q�U�����C��k�k�xs�?�Wa�y߄,�a-�*U�뫇��uM;���ح�-�RR�ɯA�Gn�i�Р�>�Fp��g����X�6*]�RT��ӏ�r���o�\��6�y�h�� ��T��С�,b�=���=�Q*���uÍp�_,�f�ͧK�A�'���K~��7Ê9a����u0�����'B��f��l��Q�<���:��vFn��\ӕk;8e5�}���%~�����mI ].�EHI�{�;��GfMF#�_���Q۳�}n|�B�$)���l"o��a�JD�kgC��n���nm_6��ps�	yc�d:=1�t��ʯYM��At�7���YZ��9�"�S{Q���I�|�<��*���X8.��dY���J���f,��>�̞Ǜ��՝sgt���S�ۍ�p�d>���ْ��=2-�8�q�mf��m����<�Z�1R�e]l�������ȡ^��r,�
hu4Z�g~;�Ok(��mPt��#{VW�ޥbWB�#��}:9��)�ѝ�����7�_��-�n�XR��#L�&ݐ����8h�c.�V�����{UWm���^d�3�6�׶#����q�#�Ż$���?�u���k��a�ҷ� 3�Lh�`<*5x������1 �"<���7%@��
h��/0[�%]kw�|�U�⥗� z��)�,���6s�ǙXS�.t��7xDR���s�����W=�Q��4�_
�ۊ.h����3d9N��;gY��ol5��X�غ��9n�lSS,����PT��p�+��f^�����њaՊ@W��,-��k˛�Ba�)������)Y��M�{ƛK{��,��6D�<��<��3��J�K�;Ox%Z��͸��6Ǳ�7^��.���ve.Ƒyjni̍�B�V�5T:�?h��t���X;�����d�ڂ�#G����u���V��\z��Z�	n�9LnAB���D�.���Ѝǒ�	'���)>	���Vѳ۷6}T�=4��
��!�愦���z@�-*k)n-ӧ!�sq~���sb��G�u�������
�Sɢv&�$jC��O9���ܑ�%X�>Y�#��|Ŷ<S���̍]�Y��9M�j����=͓s�.|�Y��sW힓<���`��]>SțY�.W2�i���3�z�����^���������Hc������0�+��S�5C�z&���܌1���K|<�z�����O��x��-�`cڥC�E�;��iD=G-���l�',�����;�SO�.t���T����s4[�uf��5j�5w�%�A�]�����QfU�R�5�Fy�d ��M���*11��;�4{�}� �I=(J�����N�Ʈ�t���4%�1���i���9�}�S}�Ij�O��]`8�gdnOg?�S��݆�iS���.�y�nNL��x�v�q��w?����S`���#���,�-�/�躑��&7m��=���7�q�E��Pg���˰��Dn$��.�_�۶�ɸt⸤����S��O��U�c�C ��A������:1���������Qv��O�5��CI�J���}WJv)̌�&��L�EZJ����_V�n�8c������1rCGZƑБ֑�jp^�6���ea��@2�0+�a�����d��qQAw�(6�N��:7(G=���k�w��jEnϮi�
A��u�x.Ղ�l�k�USd�4��Y7̸f�{�g��a˹�ԁV� �NEH�����O������{=��g���{����	T:X|�\��#�_V1x-�HuY�Ve3�r��B֥}7dڱ��<T"HZpn=��D��T��X��[�jM��4��`���n\�C��*I���3%���w���H;Y��mg���{a��ńr�Y��#n;�ze���]��կ�:l�i�19w]�V�pe��}�|�%F�yM��۲���E�CK<�@��8�t�=�t�Ȧ�
��p�$��wD������9:�����:ְW3��N���;f��[��"�Y��Z�Or��<�ˏ[ڀ=�n�.���R��y�|�	!Of���v�n�ޚ4�$��,fh\�%.��Wx�ٖ�Ʋr����W})+y�׋�t������o�j�:n�kָq��C���qt�OB��2=�Z��:����obȀ�(���OdW�2����}y\L�
u�8�"G���~[���̾��ݥ�`l����s��4KV*L��O�D��;:��s�Ty�zt�C7n]�C�[�]�ѷtD�3ٽ2����>/i����&�+��YJ����v��gl�9-1̗\�U����v�6�]ʜݳ���c�d;v�Z�����{��(��}kW!�_Io���P$w�QDRZ�B�\�/E��FħH�[��t�sc� �a�X+׵���x`�n��ܑ \��pTݥv���d�pqE�����iJvkSLzXՙ�g�˷n��:��)cS�*"�z.1q�&���h�m��N��2h���0����v��lR(/w,ZZ
�?D8}ޭ�{ͼD������{������-�ǖn�!b�]�T�v���)����A�L�qv�0k����J�R�*�䜚��ʼlṱ��l�5l�
�w=��+���"Җ���]�[X�;�6]����Dz���O1��Y�:^I��A�h�-UĮ
M� &f�ӌ�i�&�,
�k\lݪ�I��ؙ�G�Sǎ�S��u��9ut��UA�&q�f�P�缂�G���n�y��̥�y$��#A�i���n���jowr����N[y	���B��jƗl��O�^'3^�L�\yٷ7]���̘��y�����ӡ�6�̮�i��m"�tP[�#�a*�`f��r�Y#g t�����b��PkBmX����MíM��&��L�C��e��Ε�v�	���vu�]3-�6�[��� �oE��25���h���fǧ��L�M\}�9h�������$�t���r���ӎ�&d��wT䮆�:�H�C}ާW�<�f����M��k�o)D�]F��8o�ٲw+�\�z�P�1�:��g��F�a���UN���jf�xh���՗\�R��n�I��Q���PtF>=#�F��+A���w����1b2�7�^WN�x�w��j�B�7q��Y��Y/�'��m��v��$�82\7�jn.}�T��0P1UZh����jj��&���gED��3TF�4[h���SF���i�!��
(�5Q1ぢ�*`t�#�L�Cm�(�����\5\TQG �ܳ4QM5D�1SUES4EUECAC5EDMIUE4QA5EDD�L���tT��S�����$�*
)�����**���b��)�EUDE�������Zth��l�E0L-PSSUUEUU՚��CMUr�X��]EG1��*
���b����("���"�"`�H�����E�r�\�DF�bH��ME��K1TA��4rqUAM��EEu"�֨(�cLU3Nƪ���W6`�lL�T��z�A&ي����l�)L��UATUUEE5TL����{�>w?��~|�{ny-�������.�Zڧڨ����g�x�=v�"6��u���C�"��*�(%�G2+FD�=�v)�������+<��y�t�M�\K�v�%���UU-k��_���>J��4q�J�ܸ�מ'�q�#1�RYN��F��>��J�6���B���i)�ʗ+O��_$vJ���#�kN���~�mA������F��Ɏ�/��rע��wǁ���r��#��.\���N'�3����=�R�w�h:����`�PROf�}� df���F�r�E�:�@��`�<�#6���wd��K�����2�pg5�vo)r�G���{�����Ӿo���G�Dn�DT\�w��1иk��|g���z�Ԫ[���;fz���g�͚�Þ�=�i��r7�qg&�RD���r���>�n3�y��E�b�3�_��\�m���9ú\V1����VM���DH<H���n������췲j�������râTj����"�5�eM��2ԁ84���O��o�9�b�����-f�!�f��C��;;x�2���Z.�\�E��z���0��[R��7i'�x�N��$�qd�U�R/^�5_R�h�k��}dE���*lfv�)ӗO+�|�k�{�j&��0셩@�����[j%�.�OƧ�fA����9ֺ\�,j�P�U.���~�K#x��0�Fv�Gu�n�|�=��̓A.֓��p���Ön�7'5j��f�;��Շu���:+ȣ&̚yPw2GM<�P@�$_p���c-�̥��4�:* ��#o�CjIt���9�U�S�n��a琻����3W��.l���H�G��fߥ��"���d$N(�r�.������5%������h# :]"4��_T,��>��˥l��{��X�-G#��N�?6�ϼ�e]!u(��]1�ȳS�/���b�-��K ��]���g�w��gp��瀘
R� �l��@�{b
��8�e�mz9/��ai�2Gmq�껏*��b���
�du0}�l{�0��x�eS,�zk��Z�?P��E6�[y(�;T�]�P$�c��$mE|��-��VZ9�Վ3^7Xo�1�X�9�Ƶ0�H&ob֩��z.��^�M2�E|s�Ӎ�}9������>Y�o���f,B��/%G����G#o���u�t���=�S=h*i4r&;v���vs3y�6�{.�僚:wn<D��Qi�+�+�Z��Ou&�\��Sn�]Y}<�"�WGBd��ܚ��V.8R$2����= j?/p�A�{o;eOb�����xȐ��Y���/�1����j�\d�K�7�ҢD�3��Y8۷bsF���t3��E��£Q�������"������bk/{`^���bq���@B���@ں��d����
Ὕ�E���M�i��yjGE<{a��t ��Q��jz���rk�c���J]~:��w�]�>��"���j9�O���½�(��l��[��L@�!e�*ѿR����krr�^�hw�ݫ��S�{�/+g�q�r�$ Wa;Ag�B5ǀHE8�~�~'�J~�õ�v/R9!�}Bwd��Ͱ +����_��+x�������7���
�����e�y$a�f��s�T29� ��}��D�.Á_e�
��L�$3�k�8p6GIc�M����W,h���f�nY9���s�rM�)�w�'e=ktv��=�\�oV[�p!x�V�տ�9�p �J�����fWH�0��+����6��&�t�?!��.���tގQظT�97�y�o7�d�5磝�iT��y3坳�}!�ly�8An1���=��Nb�$l����ʜ�5d����Q�e!q~��z�|��a}����j��Lf��gD=Wl�a�	}��3�UqE�y^tH�&�H4�<�x��1�5���:[���Q�T�6t�BΎ�@�\Q��iW���D��3]Eu���اv����;=0jR:Gdޚ4�����~�����-�1��s�dl���{�6��m��B-�n1�n�]�Ź�Y��å������}��y�l�@�Epn<;aG^�٘�DH�#���|�_.b
�e��4�8�Ӎ݂��Rk�����}
i�&����F��tn��W��Wgm]3��y,By��Oڬ��u0K�վ�{r�0c�*;�I-�©�t_��&ʽ�o�	��,r���}��0�����*e-h��1�1�ب��Wo�28i�ш�0��Ɩ����w;�Bbk���匓��b�/���p'�s40\��B���W��7�Cݑ�X35��ݍ�vcT�nۚn��S�z�������M�W��4�;�z��GY�DTQe�R�1��V�t�q,₸8���S�vLl���E�w���v9�����݉�˵�v�sN�PAT��煮��M�;��ku�#�۴A9ۜ-f�j))�F��V�j�� �NEL:�Jw�d�q����nq��k{lp�� �^n���U)*n�t�}��.��6�%5*�i~��FF��Z�_ބ���q�|�q%�PlǙ�g�P,�D#m���i8&A+�t�A�M��%5�T�Z}�k�S�z��X:j�ԟ��ӯ�ps�;��V�0�á�1���c��L�-z)k��=��������K��]�ƥ&j���2#gU�F��Mlܦ�UD<�H۹y=xЧNovV��G#0-{i������?
��	}>�aè�#���$�ύ:^�4e�o��lʖ�'wXq�w�N颬���a�ƍ��4{l%����"�U�өy�/^�|���~��]=XR�������`X6�&^�BGz�D�ƕ��ev�,f�.��^G����7+�]�GS#���%M� n�֍DՆ�\��:Ms�A���������7:�G�{�7�]o��4+�s�[���U��Hv�l��Þ�Up;x�d�'l�<��W>J��0�wi}�-�X�`.�c�)f����4�	��@'��1���Sۏז�D�>��U �X��ctǳl�<HԈ.��v�I�yf�#78e��zۭ�ՠ�ߧ��!F��5uC0�H�oX����:�u���DVU����\I��V�zY�,���:���͓�rU;�m�E����q�{=��|mI��Z|z�\ϰ���<,A��!�_�ͪY�o�8�Ud��tR(�6dЃʨ�fWU��D)>�~s�y1}�V�Q�Ei�v[JJ�xJ�QR�Pv�m7Y��S��O�}���e>Q�TO���:HW��5�:ܑV�'=��T͐�b��["�<��j�˔�����ќ�c͑3���$�)V�a�'����Q������;:��u��3��9	���)�7�!�7q��(�Y��<�����iEij�a%�Iq��� ��N�J�v��O.�0E�]�e'i)�r:�|���
�ؖ�id�J|�����������j�R��e9]1�t��ʫ)��e$6�$75�l�C�*� �$�v�Vu�K���_0��cp]qȜ��
�/��Lsa8�3��`�7�/Z<��4����P������`��oP��@���fSm����7g�]�=u[ǕZ�1BV쫭��7?��q��, ܄�1[�C�h�_K�%g*T+��VQ+��\�]o��D���~�Ј�#�	�Hۇ��܁Y���#L�n�GH���sJ��O��b�?.�w�?S��� ��#}B1����j���&��-�λ���quˢo���O�� �=~�p!s��\x�)7x��h��fy������M;Kw�:�%!<�G�
և���9�B��������&�gs\�FT�����@f�>�;!"}��x���������2��_���ܙ���z2x��~��1�]M⽧�O?Y��0�²�7�|(OSggsȰ������f�nc�OP����U]K�\x<Nv�Xw{�������D3�22Ts��ܧ1���p\��2�����Yڳ-�<�*Wj�{�fɁR~�g�&:��Δ���vg�.Ƒyj}sNV4�qC6��g��2Tm�v�1ᯠ�P��K�bi(I䕌[*���[c�ђ2���F��Ȣ)z�"j���,��!! Wa��7 �ڡ.�I����O��a�^ҵ�M�V6�Ǆ�<�H�����[�;�xku)�Y�7v�t���	'|���t�@�q �dWd�	�u^�v���ط��l��D�~0J�i�F-���m�-�S�`�5�C5D��f2�g��D�W�6�2V*Òl��+^t��`�gˋ��/[e����JƵ�3t��0X�|�U����7<W:W�wt\�t��K:�u3�k����$��r]v9����OGQ��8(��~��Yl��#�9�kȬ��� t�2i>�Ϸ� �8��Xi���vυ�A�������;�wW�kV0�)81h��wjǭ�C_қ`s�`b�X��h���ln���⷗LwQ�t���=����Ԥ.������̣�rA������
53e^:`��+`G��D�;c�J4���e��]G4T[�NS=6/X�i�hR)��/�ؿ~�y�H���9���3��Yz��\�^��_w֎Dw1��/�r��x�l�'E�A�]��wG�"�{m]�y���n��gv�f�k5������#�:�;��2��~�em�O�Z}�C�:P�EP���y�tm����y�X��ȵ\�Vt��0rH��C�f����C��ܰ����E㣲�2W$:�C�q�O3eC�̴>ƫ�0�����l�۷@,�ńZ��ī&6F�Cy1~]�5T�Y\�w���$���j���e][�����A�v���o,Ed-�в�wL��H�z�׊R��.�S��g �r,�l=󚛩̗��v�R���85�#��*{�2��@�R4���stdC*�:�S}YQ����Dtp2+B3|Z=�)!ˎ4i���P���D&��ɂ	+Jiz}ʴY=���\��x�Z��h� jm��*��c֡�����ݮw2n!���!Ǫ����X�wSE��ٜ�@V�9W_pV�,��>}rj�*}n+����C-;��^-E�,ͮ�*��[.�Y�u��y�;�:S�a�؍��/��&�u�*�r���}�����Wmnkɚ�m�};���t0�-�#z@�������N�o�i��3 HS���k�'�%��9M��]!v<`�m��C6�q���B8��B��:4Z��n�[m]�ק�ǤQ�1)�s��a��� ��y�0�8wK)���ȍ2ݚ����Ĩ�s-[ș1�>'pl������C�YRͯf�)6�=�Y�8i��C������g�Q�c���^�v�u3����1�Ry��idxM�_uh5����J]ø���#5�����
 �P��2e^oK\�u��T׮�Q����a3�Z<ߏ.�Oz����zٮ���Kۄ�f���#_WE���Z����ä�س�
�ۣ��������&�S���֪č��UN���K�?��ľ~  ]�DT_����E��J~��p�X<ϓ�� �e�f &�V`Y�f�edeY�f &�F`dY�f!�f &�e�	�f�eXdY�fE�V`Y�fE�FdY�a�f�V``Y�fQ�VeY�a�	�f�V`eY�fE��� �#��3̃0�3"̃0�0�3 ̃2,�3 ̃2�3 � ̋2�3̃0�3"�4�3̃2�3 �+2�����q�U�UY� fUVe 	� &P �d	�@'�y� @�DdD	�@&E@�e	�& �@��<  �UY� &UVdP�(��@d 	��U̪�� � d 	�U�UY� &UVeUf �UY�U���
�0 ʪ̀2��( L 0̋2��0,ʳ"� L2��ȳ(���x�0�0,��̋2���*�:p,����02�³� ;�|����}���&DE�?��ݿ��>}_������������w��������ϯ���~�����?��~O��ʪ���~�����O� �"�>UU��������?�����������!�UU��������Ā�!���)�?s������M�~���b� DaT)@P  �U� %Uf  � ��  aU`	   �!Ua` 	F �!Ud@�  �U� 
U�@�U��H\� � ���������@�E(@(@( o����o�����4?����?C��}� �݃���������=��bW��?�?0?����:?�  *���?N�~�� 
�z��+�(}��PUW}�y��p  ����0�K��#�}�G ����O�xx�����  ����O���  
��=%��������>�ׯa���$�����  
�`L���UUE~�>�C���t���{�����@�{O�����{�`|��a'��� W�y�d���� ~����8��{~S����"���|0`�>zQPEכ������?��C�O�����)����hcv��8(���1���
��TP���R�"%D�UR� �T�)EA"�UUT���*�*Q$E*�"�")TPU
�TQT���!%� �R���%E�*�����T��("�HID"�H.��IUR%(BR��RU�V�	D]�uP�� ���zeB��BI*!R�TT�JJ�����(SZ��Ҩ���R����
�����R�(�PS��JU"T�� m"������8n��W[kn�������T�M*�[e�٬iF�3�lƭ)�5uR��ꚻ�p�i*����꺣l4�"��ݻk�i��%U%J�)@�I) �СB�
7z���:<uw
�P��C��tn ��hP���`{�:��Ӷ����2�n[��(:���2P�ڬSC�]���]��V䔤�� ��$%� c�^��������Jշ]6��wS��Cv�f5��rwdHhv�p��Ѷv���������;5��)�v�Glw]�k�u����K�mXJR��*�*%T� 	� ���]ݵ5.�ґ��AmT���N�w`n��nͳ��T魕;u:V��Ƈv	Wkf�h+V�
ژ��A%�*��5H�T�;� ��V����P7�Wl40�[j#V ѵ��
�ъ�T��m�M�V��6$!��B����R�  �
:У6�(-�Ƀ44��G���ҥ��ֆ@e�0��I�a��@U���PQ4�H*ET��A�"�� t�QE�M6��(hV2�3lC1a�Y�� V� Q"�� zkN�aЪn @�QR�QU*B	R�Ux  �� ;�� �L�l`�  5�� �J�� ��  U�@ t�:���@ŀ]rm(
ER ��  ,y�= )�X@�3�� RΫ��( 7kLt4�uC���0  C �@��k`�I` 4�T�J�%R�R�$�U� =�@an�4hu`  wh ]�P�0:�Ϊ��C��@Bn�P ��� ˄��S�)J�A� �{FRUFC@ё��SɓS�   �~%*��� M� �E  
DLj�M  �T����Q���dh�+Յrg���6��D��b���U����伽�F\Ν�<
�+∊��ڂ���r
�+�TYDEQO=���u���e�?��Ǜk�)A��+U�r�V��O/(c[{7*;#I[%4FU$ �����IC�a�RO�X�J�X8)��S3oFYytb@`�7/��Q�:(U�lm֨��[!V�*\@�ɧs7rCCjcȃ��y-�(�
��`���~�TaG0@��(�LO.��km��ૉ)�m-ѣ,�[mŭX�2�3�*]�,���$�x�	��`6��Q���֬VP��Pf�64�7�*�h�U�G�P=��T�\d��z�xs	����L���.�4��f�x9���v�u�f�ëj�/��a�,��־h��j��s7��%)�:���׈��m��wZ,V<
���[7[����J0뱥�Xu��.���Z-lMM�[b�;�.GU�L�b�)4�6�\:�+��oM���T�8l|1�c^5�A���&D�M&n�ka��Xф������� ̩[[N��je�)�+�CN��Vb���j��jVe)���f����v�6���Ϛ�Nm��r�VS`�B��2օ�nF�VT�V#"�=�t�S�,��[woB�V���L��m��dH|:���E��Rhض���)�Dyb�	��0BN��"��D�
�7P���[�e(��sA�R�1U�*����D����7g��f���h��4�� ��&*�qY�r=ѢS���fAV��˼�R0�{�f�2�;aksM )�źʼz36���Fҭ՚�LC)f^^��'�����q��i,�wh��e��6��TMmA!�=L*��p��z��
n����l����Ѕ��X 8��e�"`KtV��4�)�Z6����@�.�oiݛ��w3#yVCAU�뺴�2�%�a��,ͫ
(LUd��{aa�)k66"�E�Zѵ�Y4I��6=��l�]�(9��a��f
0����"p�_<�i��h�am��q
͒�h��[���[�����U�ڻ��k\�E-C�6ġ-��\����e�%K��N6�U��^��4�kn�4κ��aȁLV8��ڧ�Ɇ%k�y��o�mG��v2�ݖ��,j2�XF��Yb��L��)��K�ۚ�JN��lOr�,j�0*WM@Y�C*�Ez�\J�t^��Q�an��f�[�kR�5�Bt�K%��lS��&m趡7-��UK�q"&�����ú؝�
�4�N\��b��O��������@4���-��Kp�����世�@�ō�n�1V�x�̘� [��^�������35^���u�&���ѬG���&!Z�4p`E[H�ۗe-0�Զ���'/[��n�-� �]����m��*���٦���+/�-�L�c�HS�'[�mH�>KR$޺ݑ�}��S%����b�dn���Q�\�Sb:m)�J��<!l��	����ǿ�R�	N��x�Ѷ֜"�VSglب���k^\��"b��v:��x��n�,3U�4qEu�Q/hR��C4$DXh35J�KE�&?������(����ٓE��(�z�L9m8@�*�k�?�l2�S��4މ��U��[miPҧ�^�@���x(�p̎<�6Kz��C8f;��:����S'%ۅm'w&e�`��m��,�6�&�,� �m�_���9���B�ߍ���!0w&���+�H��T�jx�J���,ƥ�3�i�$�ťQ&y+&	w{tX�!�1�E�x�ޡA���j��v�o���1��h��Ha0z%GT��b�5uf�����8c:#��+��݃iP�Ĥ�cD�͆[�I���吋�JV鱂�'Y�|6��:T+eX{��Tz!s/3+l����=N]+Y��N�JR��ť
9J�<�w0�G�5eI�˲����*l�u�2[f��B�چ� �ۻT&��ݦ�m�vh��TǏS��&�F��C��?I���Wl���\J�̺����x�̚�����h
��60M���"�n��p�8m|���kĒ՘m�g=Wb��T��!cDJv��[�Ἱn䕑}�[�V��ܽ��S�f)u�"!�,�Aؕ��usC��ib�X2�/�	��o-����wGn�y�6&ySr����/RVX�v�d�k$�L���͏)Br�Я`�R�l��m�+����Qˡ�CQ�3t,H���4��ݴ�a�H����-1��05'���l� ��Ÿ���V�e��h�H��e�MVO��jQ��٦L4�O�ܓ[u��	JIW7B����-Oh޻�W�����ٛL\Ö+E�z����r}��dFi�T��b`n��ɔ�ށ.�z	�Vn�[)2�hѳHeY��C#���4��8�@ݺ��v�4�w��Zz�6��6�ۥd1����N�L�#.�@ �#����J�շ/R8^��Ǐr?���&-56'q��z�4r�q���d����A3�F�7/]gK*��])��qĕ�SSɰj*]�$]?��������`�k�j˶؎��U1�J�Q�SM �e8�m�H�i5�V8&5r��=P޽EYo.���y7v��E^�i�q��&�̲��^�)#N\+&�$�Z9��R�޺T��c��Az1 f�Owi��12�s&[La�Sf.L�[�Ӽ�V�YcbY�U��qѤ4겅���on��+�JT�#I�'��B��`m�۴h'f�!�I�X�*�PM���tB�HeD�J�]�Y���
ғBpS���/,C�R
�8�&T���A]ml'h$�[4�KtԷd���������,R"k���3NYlZ��ۛy���2v��h�o\��M"���[Co�a�K�s5�o�ܼ@B�Y��hS5��ۇm�QT셌����^e:��[��7E��T'B�԰�m|��ŉ�Z�7W2���b�.�|����n�ZB�槰̦^
L`���#5H�oV�Ȟ�?��YLŰ�T	"!��&��,n��x�,�9e3�t��ne�n΃,�L鋳[�.�;�l��3��ֈ2��DOSf1�
�t��fa�*�d�C�X`t�Ʉ*�1��4�Jf��(n��]!cr�n�*E,��� �*b�"���U��O@
*�9���W�F�P�7fG�sv�ڽ��鹯(Ǖe�
Q���zK�m�ue�[fR/.;�S���RU:.nK*��o^<7���b*.�\����l���jtFj�j.�ս+۽�f��*��@EJ��-�����-�-�u4G�	�z5����v�淲���e�M<�����ux����Q�1̈��v�ja+�/�����o~�*�nn�i�ur,Usm�(S3tZ�If�/%
a�ԕ�m\����:PV*�)��4PD��צ��ˤHR^���P�ٻ�I(֪��.���S^��FQ�/�)���c��hЭ��f�wn��ib1���i,њ��[6���Lp��6[Y+�r������riU��L��նũHLUz�^Ȝ�;��%T`��8�ֱ՚�mֈ��c���r�n	�����\�.�=o���݊1�{d�M�d�y��p'V��nL����$p�7+]J����@>[�;���Q�x��rբ�"Ti�������;R
 �RjKŊիu�(e�Z+J#SsiI�#/��V��{�ݎ�Q
)b�,�cU�4-�5�ɺl60��̢h��&J�xV捲��3(�`h*�N� ��(�Sr'��eK{�Y�N��V�DE:��A��mk�E��L�2�X�P#�Y�*wG�N�]jƜ��ay1t�J���)J�LQ��cӗXU;y���:����X�q���^ݳG&�ٖp�5��*�֥wc29����nMޥN�{ABh[om�m�e�d������܇a2�!	�!�6�6��7�����"�������k*���vE��V� �F�X��C5 ��M;V^ͻ�A���V �(�Ğ��6���wCH��b\���2[�x����d�J1t+Y�Ĭ�WDk����.�#$�ecE"�wu�:�YX��u��$��g����f�ԙ=p���H͕v�&*̿�hb�K4BM�2�f�oi�"@C��Q� JZhk��cKn�;�%�Rb��Ù�Җ|"�!�h%C>�����h��M�X�q�D�	6-��d�%�*�c�t�ڹn,�اV��o%X�%c)�يl���nJ���p���E���wP��7[3E�.��Sw��QO�ܗ�b�{AHɫ�n�kq^M.�hբ���<B���4ō�$f��&��6�蚰^J�8�8�l۶�b�Q ��,]f[tQ�2�K�O^(XDiY6w/j�x!A-N�5��8#��|�n'A-qj����O�#0�mVQ��ޕ�����@а�)jFbԒ:��0�Jn��V\F�Z���Yx25� �-����ՇE�ר�	+��9d���3wNU�G��������/Z���b���z݊9W�Yj��N���*�7�29w��i�t��6�ZU[�h��Ʈ�mC�ހkm��Ǧ����)��T�hQ������Ϸ#W�^0-�$�5��t*S���)�(V��r�� �*5o��y�'����y[�^Ы-�&�<�]a�S676A�k12���Yq"���R:��;[�} ("�"^�f=	ލeT��\�E؅nP@V�Y��b<,��3ZG��e\wB�sm�ۄb�L"9P1fT�J���{�d�FeѤ�VX�g�/��tm�۴u]���Y�e\�[ki5%=�Ǐs2�F�-����j�⫹�E�)�	�d�$��ksՇ��f���!w��򙙬��#9jV�\��.aɢ�πLQp^�Mj�w�8%Xp2P���M`���3mUr���qj�'^n��$n,2�^�Al+ui�`kF�ck�ֱ1�V=5�X(gwu��ɶr퓚�ZJ���Y�dn=�W�����P���:AMa��=��[���Nl"]��+t`�Z���cn�D�FC(eow.��]�C��K�͐�jlh���A:#�Mސ��3�51�R�;�ZcN�O�4n�s��١��kD�k�`�E�֨�5Mww%����̋j�9J��6 �ci;'Tj*יB������t]nC�P2i��"��R�Z�}��a��N�A��{���_X0�E� օMhd�,��rA�¬�hi��W�I�ՊQ�,6��jܭ�0I����J�:@���lbD�ޤɡ%�X���r�u5t�6m��7�͒�*�3�������M�J�m�oe��S+6R��mQy5����An�m�b�� `�����[���=���F�YvF�z�(�F� 4fk�.:
�u�r��N,6�¯p�h�
��n<�
���"�I��h7���,4X�iiPhǡ;�q\4�e�c`$4�iQ`Y@͆��jy7"&�-5pYl��	�6���H��3"��[@���I���Ū/�i��r��5��Ɓ3*�wR�TY���*᧦���b�8I���E�EC3%�UhK�w��
�����0Jl�Ov�����w��،P��Z�"j���vC%�a��_:"m��M�Oqe�Q�c	Õ%az�)�@SE�X~�M��\R�qm�řŁdqҢ.�]KW����2(�c��k[ t���)c �[ɺVlvCj���cR*�B�;�Y�Yh�X�'+u��A���7.ZQ�g���cX�ߦ�B�n��e1#f�]�ED	��r'oFem��Ռ��EkY��i����7K+�.so.<N�ƍ&t�6��"�v��A���/Rmᥘ�Sc6�Ы�W��V��J�%<a��(�9G~CBf�DUiƳ%Y�e`fR7)���D;�i|a�Cwd\.GM⫊�V�=D�X�T�!��n
\���A���,��-�� 6p$2��J&�b���\ ���5XB(e��ܕ5�x�C��7�����vS-È�[d��Q�:��u�yiHx7sv4T��le�1>��%��0j ����i��m�W���/�ݩ3R1���Ct�;�7���N�;��� �&4U�����(�HԒ��H�EP��~#��[����Ǭ�hLչi3��[�(S�kؙ��{)A�R��,�5�jk��Y�Y���P�R��WL�����k(P]�%��	� ��5c�@2Hm�	ޥVo ���X��6:j��E�P��3��yb� m��ʚf�Q��M:�;0U�z����Xs(FT[۫�@Vۙ��H�e���LV�ֻ*�i`kq<�T������KH�3W�n��n*�����;d	�"l�7��Ur"�^]���dh�.�N[e$1F�͊�ԡ[5\Q$n壵�$��� �U�0>݉���*��e-4�^!�cJ��aZ�x��x��8���0�:�W[(��� �ݗY�%��)�I��dlςb�6Yq�M��	����z�R���Ѩ3 bt
���:pU��A�◩##�wPY�V�RTΙ��f�MހQ�{mPA�M�㴞�b��j�2셓4��b%5��m
Ϝu��lK�V���B6YRk��Ż1){�^��&ļZ�d�(����U�!IG�4A���(J�ݜ����*IJ=V�-�H�nB�T���#�H�i�Ȟ�4S�1R�z#n��.�d��� Ӓ̼ur�Hm)6��e;�%����n�E��ԻˀŰj�Q�;�fFҴ]��Z�O_�n-膥d��,�<ږ�'�f�y�
Y=�$m�]⻃^]��iR��zw.�݅��h�v�zr���+y�h(4�t����HR��`����pQ��e�S�eI�{���}�=�i�rn�5u�bY�\�y�.O�7��)�=���z4��M��8��)"8��x�xf��}3W	tc��M��o0�i�ܾ��X=(f��-S�JkT��W��ꏺ�����Np�RѠ]u|&���*4�,�p0�W1`
\T7���՚"�%&�g4��Z�LU�7�Y	]&�v���N�����V�-v�C����k�j;X�}w5�<�;�>�39�*���\ҵ��8<��d޾��tʙ]��hI��2�:&�*��'5���zu�a�B�E;�8Hv��Y=u�2Xۨ������v�>!�8�&��_78g�]�B�P�#�@:�nӻ4���q1�\.�K�,��������Xx��Crӽ��5��n�ֶ�L\l!����D�WJ�P��]�3]uZ��w�1D��qg' �9	=+Fc�J�s��R���=��tv\�jnJI^Ko]]Z�;뽦�U��o�2��S�����,�*�˓����QVzq��P\ćS��Yb37Pt��I�n@1i���*S� U���3;���8u��q����}y�i��t�z�J��b���a�*%�V�r�eR�s�!c\�x��,��W��4�u��k̭��L��.�˗S,;�#c3;��
�U��Ǌ� �-��Ի��i3'XΙuΤ<p:d��A����U�����O���u�y09|����j�ピÓ`����ew�Đ��s������;�
�z��`��,`�w�js��D̰��Dr9y�m�ĝ�	���� �V�Z:��Z�̗����j��b���=V��S�:5Vӻ�,L�T͚̮z�O�:I潓g2^,��OY�Ҁٛ����s�=2�z�\����Ï��;��n�J�b2$/���jA��Y��B�J(��32�5���3X��oCȄ�����Y�u�©A˲�瘕lq�/ox&c�ݾ�{Zza�ɨ$���L`�0�I�L;sk/��ޢL���=\�U�ԑm���굪�]�*�.u(�w϶D�fEKh��RT~Cn��|S�
��MދV��+*�I�Ȩ?��D��]z��WN��/H��<��VtC,��U�9F�cϞ�T��6�'��}�M�:6a�(�kO�4Aa:M�C�*���q�=�*㡵,��bygXx���k�ې�З`Rf{�'��ЦM�t�j��R���@�][
�o� X҃[Pbb���	d�K�jm���ch�;xqf7��F�f]V MXb����e�:5-���"\��x�rt���I��	nվ;el��µB˔�k{tr��Ä́ѽ�`e���gt�J�dΏ''ñn��rY�(B��ǙX���m'��_�o�^8���%iE��N�R >Dai��܇�WU���"��,�m�`�+D�h}���LHt��-�y6�gYtM���R)[]R��ӣunN���;n�p��\�>�';��P˰�K�ʅ��A��l|E_lOR�x1�AIf�����;#E�̾<Vk0�:d�v:�G�7N���<x��&V��/�P�n�G`.����T�턓D*��zv���oP8m|�b;�a������f��&�h�m�W���q�7']��ո1mbg�֭�L�C���#޺�{��vn�ޤ	�n�'b� ��^x�h�Vd�qϚu4h�ʋ5C����I򑾶��óq��Ӥ�|��X����X��X�t_Gw�D��kqٻ{��S�%��B�����Ybٗ����p�B]H�qs�ϰ�[�[+���r��l���mޡ�Ѭ���!��oj��=��[�`���=(�V�O^�(U!�M�4�[E֢*Ke���s�����B�u�Sh� �l򾍥�݃J��}H�����oV|(�C�	�GP��no��ق��'��Z]D��Zw�����iZYw�啣���t�k�����>v\�N���R�=Է��}�Y V;�n�U,�v�΢���ס��0.�k�3�Rkb�M�/�f��$�D��9�1վ<�6���]��:�ut��ᆅ�`3��C{V��s�����wk�۽��3S�����I{�,*�򶦘i[/+M�ܩ	eZzC�i*UwO:j�(m�f��ld��K����*,�}�s4ưW*���r��Ҡ!b2 �InH����%@̺��p��e��r�a�2��r�oj��N���,ͨӦ���kv$N�.�$�k�jqÉRZ�o;0�'�C�$��]A��e
VU
s�@��p����[�]�g�6Nw�X_

V�nv'o��u��e=��vO;ȓ�v��y�w&�T �Ԗҝ��J\��汷��e-u�܍���qv��/�[sZH^!�L�Kf2J���K�]`-��;l�/���P��E�.Vp%�֫n<r����W�Ch
T��sN� $��n
e�טv���-�QJ�\/�{6���My�3�[��yu��X!C�i���]�8�2�i�]����]�v�8�_s4p�脬R�fS���BM6��Y�6��QCR�SP�R�0gA�w\q͇(���/L�!���:����ǚc�9Q�w(���f�EZ4*�&�ށե�/��z����쩀̣pMf�r[�����]}f�MA�ޮ��jW'W`�)Z���[���5���t�_cf[�[N�;"���,��B� ��pi�)p���}�_Z�e$�����'����ѷw]t��[FT��i,���vnu_X�'@�֙n�:;Wu�/V�M>�}�vIV��D�rw_1%�
�^�ԏ0ݥ®Z�G)2Ľ�+����Z�es�0���\b�J�v�V�a�U��O{���F�K��e�P������n�J	�,�CH���j��v�0�� �g�Z@�*��1�XȲ�`�B��#q�r;>3�RY�wT�J���a�E�����m!�5^,�t��vT[�Q�-�?/�i�J�J���\���MP\B8a�uj��w��y�v�6+Yܻ�)H�V؁�}ûo�r���F�̪��;!�wx�<���%`�5w:�gszPnm�Eo[cLt��btהӦ::{ED�#�]�u� G7W�k��d�42椴,�$t��5:��jU�]��������)M�Y}�i���"%u��� [PR�����m�/K
��9�PYJ�Z#�3vA�����i�*^n�R�f�9���K��5h2���4�u����Q�uk��$UL��#���*X���ȃ(E�Z��]` ,9�.N��cDsk�;܏6����t[�]wK���ʂ�s-^�3�ң8��L'���+��cᒜ�'S�r��j�J.w��*c)v_a�
�Kl�FQf��u�i�RI���76���-���*V��n΋���2�s�n�gjW�QU��#;�V��C%�����˭�I���4�xt²^R���'�u��� =����z��֜K�v��:�^��RM�Xˮ�l=�.�Էu�v3&WCEN���M����MM���F�e��2I++*U�/l>�+��0z�4��Z��,X
�w% mY����C�P�CuD �X�VDܽW�w+vmp+g7N��g�sv�&�_�`��V=�9�����zB���j�:���OfY��V�ﴘ�>c�������A����`k �VQRK)mǣ7bE���3����(h�2�dS�ne�xM�9��Xl�LnT�q�:A�Ofy;#뮎��F�������t��ޖ�n���S˽Nٲ��oP��N�`Gmsb넲l�G��t+��/�I"��$d���\2^f��e;�qe$�gZi0[�Y3�S��z�Z�B�}�l�hoLK��O��]$�n�b�@�h���Aim\5�a5N`2�vܖ	Gg��u�c����7�-y��u>M��Z�@C,^ͽ��
wZh�wu[{�"���T9j�]�V�8�ʉV��J�5�Ț��X���YY}�__[��V���R�8� �Z%��i�vh��W$oJ��"-�u��(:�k�͇[�&����*��*rѢ�u��dzP5&R�X9��!�����<�R��>���İ������wgC%M稻���dû��v��t]�*�I�Z�4
��r;��/��ɒ����d�ފ�����M�'t�X���U�A�w�0GQW��ꋁ���S��Wf4�+�Aշ���Wa�4���ǖ(Vv�}QJ���������bM�7�d�z�.HƧis�w��p�le�r�����e#g:�9�Ϲ7��2�4���žf!�����ܨd���)[1�;9&����U�j�e�Uф�T`J�0�nKD�Y������v���__U��݊.�,�s�ʙO\j�\,�L���%toGdRvܨe�"����n�������y�m���:��|${��m�=��PѡQ���%7մ���V�>��YeL���&���}���͌K�Klnk����up�_�K�U�v�F�Xk�ɼ���`R��n�����r��XGp����ճ�'7c95�5�M�#cr��&o�0S[ڝ�ԝ�g/�+��%\qd�mɦ@��LR�v�*��Wow/�B���S�+����鈄�tr�l�]7E�:᝔�N}�V�5�N�\bM���(�*Z[��U���'k��DXac�yWe.]�ON&�Լ���=��k��Ύ����"r����A3�3ks�Ǝ�Z]YSf������4r7�M���Ò{�a��\}�6��Vi�C�˫�(,��m�{�x�"�-Mۙ:���f�H�Y;9��2�r/��ai����b��BX��v��7�0 ��;N��F	g�I�\Ш���]\V�4n�w:�8�ַG�O���b��vJ�kQ͑�����̃Х[�|Uhe���ٛc�J��������:AF_D)v i���3c
�A���pڙ	9�>@i%�r�B�nH�9�t���7��z�<�O���6�9���d�N\�R��H̜�����������=��v��mրJ�YF�M��n��s�ܓB�=�5�ӵj�)޽��Y�(PL�uو�J��_�������}��5�Ѩz���z2�t�`;L�Ѱ����8k����z������� N�_k���N=2�e�܂���q|�3�_02�S����{KkDX���;�~f�ТF�N��_3ڮ"p-�&�;�ڡ�lmf���h�.�sѝ�k{EA���XM��Gn�R�Y�b��uR޵ NI��>��;2�EC�V��u��\��.�[�]uvx`��)ި��1)U�t�oKM��v��-�B[Ѣ̼�۪��0�Mx�W[��7еvIz���|���ͻ�7��0oQ�r��)S�Qۄ��^ʕ"���v�;C�Z2][��9+';L���)����t k�㓝�}p[�7��k7���kcn�����U�ʗ}c���/)��7Da�/��󫕰7��δ�u���I�&����w�:h��s�2�ܗ���[�|��0vP��>��ڟS�O��-�n�M���ҕ^� �?9C�%K�-�A&�rq��[��[�Yۅ��k`|�L��Y�vS:����4�9��)z6W�isMݥnR*�DjNO�Ӽ�����n�ǻ��>>;�I���q�Qh~FvWi&��;��XE�Fv�ūy�&>wZ�bv�C\1X+�;^����pU2�-b�\��Ʒ/}ZwV_j7#�hi`F�Y|st��z�.Z�\t�{�M�0/y\���"��:]��r���{o�MD���qv	�L�0s��g@m[��n���;���k{��3\Uu�>$�Q`YԴ��Ge��3�����d=�2��3F�k\����;��`a�}(n�!��8T����C�7v6��&R͹��ݎ⁸�m�4�e��6�C�uh�k3䝨��'�S���6��ױ��J��+�[[°�}9)��y&�Ruh�P�Z4�1;.A��s�S]չ�������+�/�����`���2:}i�]&�ӄ��J�����	�ѳ�	}�3�e�@�]8i2��h[��;X�Ivs����C[6 ��>b���:��u7]�,��H�ړ{F�fй�R��B讀�=`��`�{s� �V��_vicf�����]-��e�_w��i�R���n٧���y����W�T��i�MefRn���y����Ȃ�,A�j�쾼D����Z�qf_v� 	����[��u>�[���9l1P�t��V+.�^�o�S*,MKG
<W��h��%j�l��f�)ffxn��uϲ�%�u���I30���'r�ݥ���bTx�u����$��]�trCfB�hCj���u+��_i(�t�ܻP�\��hkX���Y�{Yu��Յ�*�LSB"Gdf�fF�w��ko��f�;OcP�}͋����W|]���.J��χJ�s�f���������͍���X��ġ ӣʤ,5ڞek��sh&��g�+-��(�(���DF�|�_]j�/.���p"�E���+v#��1���+(p�-��V~�W0,�v�gGC����.`G�;/(]w6;���]�cy��ˮ����"h��I0�\R��e���u>��f�}�^v�S��cR��6�h�#�R(6'__��=�zD��i�]�nP�_C���=6�T�����I�q�B�ܨ7r�wj�A\;@�-%�SՒ����ݨ���{w�˴`yY�pI�x����F�-��껥�D�����3n�3�t;U���۲�u(�`�R��\�u��_O"�%����~��k]u��}�����)��T_ݞ���W&b�eGg����������u�s{���b��_:8�P��j�=���V���4��;��RWR����ҽ!ˎ4QW\��ٍ�Y�]��%�csF ���f�{����җ]5���Z$B�תa���U���z��i��m2���N��^��B��em�DSw
|7/LW�6>y�}�-`�f^T�t��Rf��
4�Wa��̂�':�uj�-��>�)�t��
O~�3k� ��io����*�m	����)�o�/U�t�" ޷V����yæ��I�6o>ܵ�Z����0��pE}�
U�s]J�����:�G���c�Ƿ�V2���Ẇ)�il;����2��1`Y��ӗ[�D��T;hA[�0���o�gG�ӻ�� bU�5���kz�#×�뀚���Ŧ�K�~2��i]|��9զ�*�yx��������4�3Mf�����L����Mr�;wtr%N�k_P�T�&��5\P�t��]���;����κ2�"�e��
8�	{���.�p�*�_a{`<W]�pY}��K[��a�d�EcP�k�-��]���ّ96��}�t]��p�Z�U�P��Q&��	Փ169���1�,�;s�yη�w4��_��r���:����:�!G�$�ZʄX���3��7���r�b��5�z4�Ƌ��.��(o��IӼ|��xf�4����7����+*�ޒ�OK���B|���[{���0굌����R�D���5�ifd3�a��u��:���{4H}�f�,.o��|�V����N��mTs�Ga��EAY}k��(���px���%�/YVcWuB�.��-6���T�^���d߲��i쌓�jG��4�C���ep�K�Q�%i�<7��C��6t��I��{�y���t��Gjr�omh�#�S�֨�\_.�9h�h�6�������Վ��0+Nn�z�y||C�WV���MDֈ�K�Y���.�J�������u�+�g/��4s̡¥��y ��ỵ3ƌ%��cN��z�RI��ۧU$pNp���,��yu����W��7�jŅR�������[���
����:ء�V̟զㄆ�0�.�=���nUHE&���k���2��wK���i�"��筒����
fWdmS|Q�iwt���+,pN/����D��QcPS!�о��M�렔�ٱ���vxy�+�:7R���25�Sh��1�ǔ����������˄���|�|h
e
�(6��Ѯ��h���������)�Y[eSON�hW.��eby��n��,�.��Z���q Ȗ�%pL���2�[� �(��\��w΂�Z4+e��T��j�c]e�\�7�q��e�Ef���,�@ve�E����Gj�K�y֋�ۡu
\����*0��1'���z�Q8+��Itʆ��*�>*Q����kp����y��8��6��"�;0f^��}��M���fN/���y� �Uq��+�]=
�׹i�rދ�Z@�H�/���Ք�G�I\顛�jb ��[�o]�b��.����fd���M�í�Ա<��=����v�r�ށp2�/1� ;C�`��g/{���],�����=t�!�P�"L7���)�7)���Zrȫ�Q[����:{6�� �%��ڜZJ�<�����µ��=�.�� �l�A�Fe��*��Wɔ�f�+N+��)F] l�2��Ooz�Y���.�sv�\�*�����nV��)��"q*yМ�)���)�/M�he"/�-��(P-,��P�1I)v++2���6�����.��n�P��W�"z��r�=�M�v�Z�����@"�}k��'����w�F�.���ϕ�t `�g���GkTn�9��J��׷�\���$[ћc��1.���l��Ǆ��r`WaR���6�&�[�H� �n�`�0}b��d��n�"��/x���X6�)-7�V��T����MKVZ��p��m��-u�g=�j�`�=ݗE]",pS��t��Q;��4���C�T�_�8�
�L�'�N��+y\�,���;JA����3[���RI��)����.�kw���I�U�]r��M�s)a��v��1�gze�Z �b3[Y�;��G�)���ubS#ٽwj��]wj]l�Ru��P[\n&OY�9L�n!�#îk��(�������k�{�qf�s5ۂB�L!^�,�D.Pb�o�3�$���'2��@��[��z�ʱ�7Z����Gx�ħ�v9o ��z]�u�̽�MjϞ�vN�#Ug!���(,燰�g8����Wk���3E"�\���\+7v�����Ozs���Q���UX�G�go5)0��Sr�([}��c��T�pQfm����0��!��3S�T���"�@�Uۙ�v>С72.���4�"��g����k�d�NFͺ��A�|�B�4������kW�o�p��Jt}�'NG7o/�G��΅m.��oi��Z�k1��(�л�6�t��W�^޲{q�MtsowN��u���ź�&��I�-�/��;��nu8��u�p *�3`s�-ξXZww�
u&��m���.�G���-��>�a*�H*�U��*ͩ�.�`���E���(ֲ5�N�����Z����s���HPP0��Q�o�d�/�V�������UV^��_V�9�Ȫ��8�=����{�Xmȋy%����orŒ��w�@ x�gXQ�Z���kO����a�{����Rv���[��5|v��w�*֓�R�AL�Ю�!���u�6*�kK1bC�Q�C-�B����ե9!�>���3��[����5�&D�tq��7R�\;V8ev>9�O�fM���JX^��pB�,ܬ�.0�ң�7K�ˮ-��.=WҲJ��QC�6�r=[�S:iU��n��2�p�3��N�9���X��-u�W�7O:�,%��s�>*v0�=����m����u.���5�^t�<6^k僮i��K�����ri�Y�ٻ��[6�;G*"������)n���)�Of�c�n4�ٻۆ��+\����b�aV�U�&�jg}�T�ꛝW��5��� �yb�;��p���k�-y�b,���Y�2%+[]���qi�O	He��r*�˾�ش�`A�U�[����!���g�=�t�ue7�+vC�F#��{��݄ܳ�gKx��/y���*�7��SY�4צּ��-�� 팹����;M�{2T�Rk
f@�� ���i��L vQ}�f�V��߆4jj�M��/w/)�U<�"�l��d�m�QY&ha����et�^���R�Q�}x���Ǜ�SQ����#7VӘ[]ǃᵍV�4U��o@�vos�e2tį��P���R�N9B�n�6��Jwvj˅W]��	��ǵ�s9�ާ(����]�(ct�P������d��~y��y��.�L�)Z���NV�̽����G�Οn\�inE�iܩ�R� �M㱂����JbP�Bk1i��,$#�yyXo&��ޥ*Y�-��AT������#�i�2� �k�]�V�F�t.�v�+��kXx�c�4YY7K�hrX�����$[Y6�:i_W6�H��ZҨ��C�`wIL��殗��A����w��-� XxZқ�Sz��� H�`8��Ą����}��}d!��sz�ƴ�RW��:K��v��Z�[[YC.���t[\�6� ��yom�<u��8���V=�
�z��>�XȶuU��^v�v��#���������6}%+ŎZ+�^�&�
�J:LB��/Ix��}1h$h]j��z5W9��10��ꠧ[ш��d�CA5��]j.�c����a�ǲX�&x�g��Zs[n]h�Tѝ������-J%�4ml4�֫	�>�5uΨ�zR�f�C^�.[w�����WPbJaĔ�J��#4�ì;����Vǆ�E|r��w̢�"Ѣ������] ��gA\�I���X����]�it�w�r�����Q����������Ri�H�L3����e����2n�,�#���S�l=�����)���ئ>����+ˈ�# �v�S�s�	�S|QWur('�f�޾���k��4mc�{�R�x�*���kM.�t[���Eu����i[�B�Zn�r�W����!�gu]gv�J|���D����A��&�.�v�ƴ�dM��iм�򚘫�ݑ__�i�u��%E�[n��1õ����YW�~F.[�H\b+�뭲�ǲ�f��蒹:�h��n���n����Ձb����)�_a(8�G�B�����VФ���ԁ���'��'0�yZVrڡ��K���>�rk9g5:��ƻ���k�iN����W�;��i���������9<���hO9-X�f�\�j�˶�����^���6��sQ ��GJ9wv9��ϰ��Xf�������\���Wݠ!6�	�W3b��zОڔ��;
��)�Z�r��u��o�N��X���ċ�ڟ�8�X�d�c�UE]�K�͋q�a�r��͇q!-vt�ծ�{-ј�$Xs.B����A�:K���)�`��Pƪ�8z�72��-�E���vv�����ń�����Ӑ�l��0�u�BJ�t[�E)����cLh���$x�v��᷐L�n�uI1Ef��Y`X70ht���ڄE`Ȯ��B1x�d����2�8��"9��Az����xnkqخ�f�;N���3���1϶�R��A7BaY�:j����kE᨟Z�=6L{z�xb��b�ݙ2�"c�i�1�8B��`��/f_&������v3�7ݒٝVQ�)J�u�(��*��vV��)�-���M�� ty4Bh�u�n��h���h����U�N�ٴ�p��Zu���w{���R.̡��Yy�S�+��P����dO�gr531��G����qM�_^���*�2�oF����jh�W��e��I�w%�"
����l�M��0�d/iԊ�QwZ���/*�^�����X��V��ܭɮ�V�4N3�����C��mk^���U����I�"_Vok�I�Yp�;�}��&:=�r�O>��V�������x����iX��̝H���α�צ�_o�����rb�-�n�-��j���e$�$�������.��bX�[-L�0-���#TT`���x �����ӗ�k��b@(X��O�����J����Y����y<����,�Movs�kj݁L���%;��R��kǩ^��)q�n!h�*rSj�D�vٺ8QXU�>j�8�e�;�fӿ�Ռh$�o�<�Y�[o/z08�q�YZB�h�L�[��받���ip�A�2�%��IIf�|���stζ���,��<�̅a'�3�,\λN����br�˻u3wjb�S�Ɂ9J����i�û�f�S')֦��z8�'5�P�l��cU��7��Z0������<��c-������UE��ާmRV�{(
�]�mq��.!r��Ԣ�1�mX�;������%]eup��ݭĬXb�Q�;Qj�h��w�9�Nn��8e8����_�6�yv]��u�:�j�m��#���)�gI�Eǯ���eV��2@��9��tE��躣;�)� ZǕɮ3�	$�̇����vr�⒙Z�*�7w���<Gc�-�9Z�d�ۭs���XZ������6����ԩ�b�����m�6�l�a���u��M̶pi�J؇�z��1T�ϱ־���C��5�5��%	�E[.QNc�jL�/���
uo�J^�ʺ,�hH���*�ΚM�\I�J!I/�EG�ڳZ�ZZ#�Jf����QE��84c�Ƴ&��󒣙�7��	��#)p��R�y 3����S�P���vw��*0
ͺmD���D	.t㯥ueh�2�c�� 3�WԎ<)T���`�Qo��]�s-VmůF���rubC�]�2+'F�WP���[�J�;��Mu՛p��vy^��u�٪�C�H�a��U���	"�P�*R��m־��&��g{,_[�N&����>}�/6Z��5��Eeϗr+-�z}�.����wz�ͻ�6h�R�֜8���]c5���0<z�l1m��x�w�}V��o�#�� �ҕch�/���d_Ko�E�=�r?�S[[]��KĖ���L�ERf���g��Ժ�4��[{��\rG�Bq�J}�+xsv��WQ��Z�|��B�@Q`|+)F��I��
 �{Ӳ�����,P�z+)�[�X���W5�KGh��	꺔�k%
Cj�D|��&���U�,:�ץ\k���ZMa�뛪nJO����'s�u��#u�,�ҘZ���Nf���!��-�X�VܘE�Wqڬ;���i Z����#���ΡSe��{ŗ����`��k�,��nB"}�l��R�A�қ��+�	t�EL\�iZ0V��w&;�(*��5���9A���P�頩.2�Rġ	�0%ÞkK��uk���Fn��#�:"c�zF33���0���p�[��!�=F1f2\�n�Y����������I��d�:w1ݍt�3mNM<�O_άq��z4��a;1�çq�Xڅ�OcRs��/k�Yt�B��KX��!��I�7n��^�옝�}�YWu��v����	X�Gyض�y��6"���͍j�G9�ð��LVL?7�8�\�Y��~�)Zuąd[��/^��ǹC��3#h��6s�JS�3���*_J�C��}׼z�����Ը깘�<��伽�O���)�g\˽D�mF�XD�x�
`N�вJ�ގ�#_�v�ml����M���)VL���P0�km���LJ���@�y��!Ye`&�֤5�H�25]��8�^\�t�V%Z�-J�]W��P�'u�cz#���iaV1aU�ҕ��,}���X�-z�/Ic����{����v�wV\�o�v^Nht�}��:��2�tڎ�{��띐rk����,|�j�b���x���إ�#�wՀ��W )��n�l'+b�d�­<��i��١ĩJ��p��u/�6�d.���,�X8N�Uʹn�=��V54��)��вkj����+�z����Ov������6���y���/W&��ʲ�a�yf������2��]�z��sw%F�5_�2���C/�|ԋUn9��e*����9��Ȝ�|E�F:�)�h[���RC���μ�\E�J�Ň��*���'Gr�uoX����ʸ�4J��gn��8{w���`g����;2p�%<���[ӂ#]k]�7�\��o/������5Pƞ��|(;�ES;5���4wo�Qr��v�P�S���s�p�YT�l�*ouu��1���GȚW<ʧ�{x�X���`�t>��u,�x�ıѕ��,�Lx/k!KZ�9�ékR��cI@�'�>�jΞzo2n����	�u�X��׮��k�����vmj��"B�8e��AM@P�`P@S@�Y���u9!JDVBaQKQ- RT�E�Qf8B�%$Nf �CBST��QT�Bd%-�U
R�!KJ�5e��94(P9�%C@�	������)��&5KB��CEERCFJ�PP�%#EBR4�Pd@L%(5J�D��!CN�r)�(J SB�P����4��B�Ѕ�˲�Ŋ��Cgz�j�Jùx�W|�nȔ<_��Y���#G>��wbwN�z�a��p�k嗏t���ӻfI�M�N�����\hF�ͳ\-:�+En�u�ݭ'8YS��3f����){��L9]i�����v�݄BƯ+��Yi��V�.�w�rO;5�w��`r~�^�|�����@:s�l���]��/&pC�QC6���������N���c)�Of��众ȥ}uE�v�����u��9K����5���jٮT-X��:��͠�%���ٽRtz�@(��h��a˥p�d:�G���Y�1�ΝF����_�m.�v�%Q,�t�vn Ӡ8\	�W��Ȥ��/�T��W�6v}�w=c���"Ԭ7 �^��XX�s�E}'y�����'0;�O�_�[$R�M�o�)�Z�6�
�O<���S�66��cζ��e�!'3HFU}[SM}ʡF�xw�Z��dۨ��4屝��"i�pً�J�ܹѐ��O�5���.�[Y1.j�ˣ��k�/>�Eg"����V�mIe�ϴ����8�EX6��JF��T���;���* �hF����6���g=�����p�A�F�E�E䖳'��X��Ϡπ難6KB�Y/�譽@���l�qU*>,�[�O�i�ά]u/�������}�3�KnVgP�ׯa���WD#hA��-��@�f�� Z�N<FMq��uY�S��,h����:ԝ9*����k-NO�ٓɜ����1��6㻀��x�"��0���N��N�hϝ5_�����q7��7Y������֒�&g�Ux=�{���9�9�1��D#Q�u@6j�e�&xR�	~}^�@*ѧG������մ��p�7�ґn3��q�J�}�"����f�+�u��"	c+��nk��]!�
Bt��0	�T��GJ& �����6�'Ȇ�.	����D��wn��y۝��e��PC�̚<۠9�{v'�jUj�:�\)�< ����n��� HK]�'��m�q�]]B���v?�����+�nI�c�+͎��p��rI�y�n��9���kp�qj����A�A��*}���0��|uہ�[�j�횑��u�{<���d��?�تJ�Ydx5����fh�ù�|e���3���=�%7��
�@rz�Nlq�9��(�Y/8��+�_�>U�c %2{bH@	�\�F|�a�f`ʭ�<|�V{/�ا���n�X�cg�B�^q�a����j}s�K��5��E�}�wc�w4U)�e⮛e��G��c;���:h�l6�V|*ܴ��P�GuGot�(i\���wq7Ż�b7�����7j��X�[ww𶻪s���>6��*:��9\�P����,���l�>>K��������W��Kü'Y{`�<�6����;3��+�6K͖��y0��1�p�h�Z6.r$�=(%��<o�T���h�3'���opГ�~ץS��e�岲)��DV���RAڃ(
�p���Z�F�>�#�6ݖ7'��{8�*Y�S}��\k�Hc0��5p�>3l�_@�:��;t*�;x�fs�]�I�l	52,��F��D��󄋉r��ь�}'�8;e�щhr��[T����<h}��R�&��6�6Ǳ�m�J�O�+y�;��E^�R���IҢ��l�xU��m15�*k���)V�zeq{�Do�'�7j�
�R�u��[�Q}֋*tG#��`)��:؃*d���Ԥe@㢞��pb����9���Ү��NZX+�od���c.n����O�A�ƆR�����;u{�z��”G+<�!�BF�;=�zn#S�y����A+�ҾZ�,�-�-�v�v�g-2Y���29�(�p]�+wf�W/(��Xy�@c���	�n��>:N��P�T6U�#2)��Gv�`��NL��s2;��Ū����h��΀9���3:Q�mc�R���q�o6󑡨�OL�}a��벫1vI0�1+�l5ӣ������N��Չo_��5���d���{�!)���O3c�1R\������ƻa�)�K^X�ݐ	�k+����۞č�\����Yb�*�"�:�a������st[� ��f$Lg]H�g���f*�v��#V*�]�+2��`��q�+��Kzû��F��7_4m�����^��Lu���ٓ������Qk�#�^�7�ͧ��P�O��+�LCo�ϥ�e�)O��_tޗ�CVo��r��l%���y�+c�����їk��P�#K��br�㘥�R��Ur�+KBL��c35��1��ͭ��]3#`6EFӠ�φ���\�,����L�|�=�<�خ�/%�P��k:��j����C@W#��U��xޯ+���B��`Q�&ǲB�9�SU!w11u[��w^����>is�@�<���s��ܙO�����n�Pʓ���m�Y�Rr�}KD]	1��臦��T��U�0Y:��@jt� �*�0w���p<�Ͷ;�[d��h΂�N�}w�DR�C8%�f:
n�us�e���de���}�F�IP)(�H��PcD�c�.e*g7S6�e����dz�񥇛T6�a/��o�����D� ���W"�h��R�h�ݬ�{I�Fm�8p���b��.&���=+=��A~0�a�N@���쌿��3Jd�Az����_K����d��u�7m�X/�����΍�T��NiH�s"��r�ߊ�#ܡk�QE�����X�I$��Е�g|����������� S%pu�"�'6��:'n���;7��g�	V�,Ӥpj.�]�'�Poz�A��~��*d�X�c4�h�-���]S� ��A1�v�
ʂ�w�l�W�p�R��jk�Wn2�)�ʇ=����P&j7�n%�A椱�2� ���Q�v�΃�'
W�8EW��о��H�mD��E8i���΀t�" m���<���9f��C��f�¹���h���s��vie�Hi���J���I���>��6�fS��U���$�f���I.�kWV}<3��wV��OSZ�΂��n�i[�d0\��!GΧ�N�wdGVp�^[�bq��'5�3QW�6����vg����w�N�/�,p
��o�I;�[�L��0�.w�^�����	f����b�As���ꍊ�9��*��{�������ᵓJ��\�8f�o��
�]��o�_"�	�Z��]{��̵hN�7M ��3�X�*���h+��.�'�)�IV��d�鯇�,ڗ��j�uR�(�Ve�9�J׼�`���ݥ}'s�^��	g�]���H�Y)��wvnM��b���#���:��W�o���r4.E�N�����W�c���I]{�V!w˦�+�g��u�we��/�f�b��x6|&��xq��W�W]=o�x�m5(�_Z�ʛ���Qg�,��g�{���Y�k�앭(#M�ı�b 1?�ݍ����=��h�.J�����s�n�5X�㖻H��I���*��ID�v��y��M��ӝ�b��$?���@��Nt:#�9�W���(n|�w��.�R�N<�ܣ����
O� "�D��1q<��\��Lb�\��I�C>r�4���m�E%��m��Զ⅒�ڭ�OJx����#ŸΟn:	�}�"�W��
��{��8�ج�[�+7%�'Lİ���1
�I���L@�>���G��a�v�}�{��$:vn��_jgVmm�����mT��&�j@ή�Ǿ�P��Uq����N���LI����{�D/]5|�<����iN��&z��b���
�u�3܋��<f�$�M8�Y����:sD,��բb]K5�]��U ��b������w`��	K�L�k�N�F�]/�k����%Ĳ�gYi��7C3zFa�4�Ջ�����C����U���N��}?95僷�پ/L�� t��}��[Nv5g��N�1�����I�҃Q�B�	S쌍N�
��	�M��.��b�b�nK^�.͇{x9q�w)�MT.�C��<��gR t^��-g��뙍I���2W-��Q��S]"��?;wR/�'0Vx�:QU�R��H� *���C:�s�9�oTl��M�2�fz5EY.:~�پj�V��و�3��\�K����ϫg�gY�h��[05g^�B���<�I{ڤ&OM5)��/���7nG	�����H	�n����]�.R�5�9��4���8��+�aý�&*;]|�\�y�]�����)��F�݌��LZ��&�W{Ȅ�w���;�;�R�Ҙ�kS�>|�i�u5P���?U��T\���w�/x���'A�.|�E�鄍���w�p�Yvm�<��)W���˟g��M\u�N���z��4�
o.�C�fJt�#�V���-}Q]��|`NA��_ENRď�Z�F�:��;�o;��6>m��fA�jj-�u����Ω�Pg:%�cԋ��^]vkʻ�
}m�ږn�	��D�t�P�Y�u��}j�we�7�N�t0�=ֆ�k�4;_s78����
��ok����������:��]��<��D�s�Lw���n��q���!(��8�����v;��A��҂8���y��ߣ��}�+�Y;��\�����&�@f��2J�f�#d���T�BoU�e�V�t^�w�qП��f�4�1����U��'��'�9��>IƆE*�wc��/����V�r��1�E}e��/M�u!��d��4�Ѹ��#\%N��D�cX)ͻ�[]^Y����oM'�C���}5��ī|���b��O�����\"�s5�r�'*�JY;��Vy�����>�{m�]j�u�U�G0��.sQB�����ULA���ݡ��\ް}m`eOW:���DJ�F�;<M���|e�])���X�&��)q٣+'���W�CԸOwdv����捵u���.�X8b����+K��Z�u���~0��绎A0r�t�s�WW�cxআ�.}���jacn�E+�� :��՛�^RM];l���E��Nҳ�u� ��b+��,r��<#6��Y�0P8\@��ѷk)�xwW��׹f�����%p��%�A��f�T�sm�T;�t/���{[��x�6����?o6)�һ�cثOQX�h��S����Z6lĞ]Y��*�D���/\W7�5�2�j�yP�{��,:�`�����Y�Y˩�^�{���p���\pH�28Fʐ�ᮬ,��+��')��w\WG �EC�]w�)�;�U�����L��#�á�5�E�c��i�ʥ+��u�F��CH�ׂgl�}��g�ݟm���%4��%�����U��K��Y��� 5vp)k����y�t�fB������E�s2�f}��h���騒��
a������u<�Qum�b̌gdtξc�'��c�ʘc��Brm}ݑ��Fk�2��:��.�W�Q.��wp:'�^�-#����xB|{�]\;>T� ^���s�e{�>���K�%�[���{�ݔ��)�a�����^V�f��C�������]l!��e�[%Xu�Q�1Z�t�n�u��b[�'j�7p'��D�M�\b{e�+!�:O��S%��S���kw��Ӆ|��a�s�=,λ��{�&��:�B�պs�ن6�j���-��s�Г�%mV��ѽ�/�Ȁ�|ܰ4�j��t�gX�	�m��[��r��i��/s����e�Z|��,�����qBO<6�Ǖ�����]�S�BQ���닻�)l���w�{,�i��Rw��☆�R��Nﴼ���q��s��R��y���,,���[b��-c馵�j�](S\�t�����wɍ�������B�B5�ۻ�����~ڄ��pw3b�nP끓��-���Z�r��\�M�NF׼u� T�w�P����!J��6�l�}���=��$�4b�WxS��	5������஧(�P'K'/��`Tn5��}.����q���I�
�(͑ԶN{��� qTv��Z>��T�va|���� ���(]$��p�=e�|-��$���+}OZ��'ѧ˥��ʮ������,�Al���E�d�u���� ��2R��$�Ec��*WN���w8�S�W7>�*܍�q'�wŕ��W���^��/{f�㜔�z���1�/�f�cN�DƄ	8�e1~�\1�dT��{]~C�#�)_�f�&hN�OO}�2�某���\!d�=��{D�����׻�P\�3p:Z?_�j�����_C�8`���-�E���0�%��*���>�H��qn���B�ME�`�0/h<��z�Nx`�M_�����>�����³x
Y
�����5��(�{��Y8 ���V�	���;UЉ���tk6�܈��n�+�|˂���V�¬�h iѡ�t2n�=�M֮���]�q��D��=$w��1殝z���D`�`W �t1�WX3;�^N� �RS�z��S���}�n�m�|���Cw�6B:����g+3e�a@C���7o�+2��	A�ˆu�R%��vw*�:�˺p�oL	�F�5��s8��=�ww*WD�O-�;�X�<��i��˫����]x٭�<���X���ј��u6EX�J*teG���I���es۟h��d�mZ�w8�W��m��rj�˄��$*�z�Y������c�J�+�����k>r�Vpt��z��uѸ��ĭ�r�j��Y��̈́]Իt"&�Ga[� ����T��%ȫ�ԅ45��<:'k�&)��,�6c��/&�f2��Yy�I�{w���7��w�vA�k���-��Hf��Wc!��#M����OoUG}�'�=;Třj�_8�J���#����\7&Ѓ)>��WK���#���s�[��ג�gy�h�77j`3Dn؀/�-��\��Pw]v��Ǖ0-����R��p�d[U����D�!�]��h�+$�|WP���V��2�!Y|��:g+ ?M[K5������O��nST�^��s_�4XAS��L�.CdW�ئ*��>���U���ĸ�u����"S�*����.�m��-�b����i���F(��]��B�Gt�u1τM�-�eN/@�zw��R���;��s[�@�ڻ�������6��˫�{j���y��e����=�]}���t��+���jXje�F�1W�A��P�A�J۫ZY�����W��u����x3It�̱"�4���7��L�Xb�V�Tf�t[�v�bS�=a(�1)ɋ:s�?y���ʖ=�sr�C�͗]sQ�e�E�qow<Y�(�����c�yF_ �SZ�7W6�#u�P���2��}e�#{���3� �s![R�}�g+6r��l.��wq��lv�g�wQX�m88V%'Y�s�Ծq�wƅ>���7e=r4�b}ʎ��T/���Z���2]W:�f�};�9]��X6=�&����Pl1Ǯ����rF��)sz��No���P��eɝ�)1y\wl(d�Z�*ήbHka�(��}O{wcc�J��8�K��+ض�ӽ*,r��o��[�����X�0�W1U��w3�W_+�Z�o9���[dr�kfm��9�1�����ԍӋ�Զ�Vf+g�[�����z�w$��h�]w{^�e<��c\pX�U�q?wbn�� R��8/��06���l^�q�������}�V��8ʵ\�3{9�; ���.V��N*޷�Un��"�{3f�Prf0�S� ە��F�׸3_�nu%�㬫���W7N��h�v��k�'r��u!�P| B��HQT>I��CJPQIMQBLA@RRd&HQH49!��H�ACM%%&A�Ҵb4eT	@d�6`ЍAHSHdVE.H	�9SB�	J��Rda#AFYKH�B9 �*R�I�4�Ԛ���)B�)�0�23 �&%
��4JU-9!��%.TeBӕ )�� ���9&B d�
eI�&@�.NB.C�&H����R� fb�'����R�3_W��2�'��%��Aƞze��=ڄ���B�u>΃+:m#[!YQ�cz^t|����Wi�V.���^^S7Tfq��_�s/&o;yc'��<��BU�QA���g��'��t��%�j��=�/^������;��\�����u	y���}�{�%�##������\�[׹��z5��K��Y�K�w��b!�}"$y̴?���u��؛���c�:�BS���%�Z�}��0�HP����%ְL����$�9Q�{�����MG�u?��]�U<�/~��uמ���Lh��]ʝ�Z�V߾�"(G�,�z#�u��cr�^��r:�e�c�y��yNK�fW�C�?}����;�S�:��}jԔ��u.C�r59ɪ�����7p�X��yw��z�o.�{��{��G�"8}""�E����Cs�Χ�y;��%Rw�>�u����k~��F����9��u&I����sI��=����:��u�S�K�Ծ��������0�����y߻RHC}�wNuחB�X���}C�z�߸��U!t~�c����α�1r~���?}֞�J}��~�����BW�{�������]����v��%�5!߹�瘺��5��Y}��7Ժ)z��ƹz",}���&8Dn���vf��.@r:4a�Z���{��n�]F��i7�e�{�}l��L�K���u���?BS�Ϲ��0}�4�?���׸o>��}��˛_B��S�/�7����7�[yK(��jϰu?F��y��A�J��o3W�?A�K�;:�p�#�uI�h>�����a��=��9.uߜ�
A�������?A��u�y��c��*g�w.l��J���""0`����4nz�!�<�y�ܚ�
|�Gq��;���s�5:��<�֍�S��VG'�7	T�����k_`�F�a�޵�FI�du�5�g6���\n�箫�#�G�"2{އu�^F���7���g���}�ߥ���;=��w>K�u�y�b�uR�a�~�Z��g���!��֧�Xn|��)�}�GRuu�1��$teɳ9azx��W��� ��  ����oHo�'۷Z�c���5/G�i���]s��9�]�U�>÷\�{�/0�y�}�%��7˻S�\��5j]F�?kP�\�^^���7�-Bq<j��nQ���8�Cj*�)�]�+^�$��.�W�*%��p����ʄN�ks�2[�#���r�*�5�dȘT���+.B8�#xǆ�+���K�2��H"R�])���b�����Q8Z>ml�v��C�`�$Z��{�V�� Mw�9%���}��=ǒ�_~��=1��G�������n7	]�w��z�ښz>�^�(~��é乬C�oT�rMG!��~����Q�~�9p�On����Hm�5�CZ�e�H=�y�>��a��[QtG�Uw����C{�z�-Ǹ��K�}�κҺ�����7#������ ���&G��s��	A쿣g�h�W�<���:�:���ܹ��>�����=�����pd=��yy��5�����ђd�sZ=�����������ԝ��k�:������sg��\��g{涼�����{�?�똿N���g9�os������>7�K/;z�zY|���y�֮���~��)����rj�C�`PPr=��	}�dtk>����u�3�y���{�ϴ�	O��O�>��d���H����'��}Y��7~y��מq{��\�����u��S�}�C�{.�_��5A�q�1:���2w?A�b��7�d乘?Z���9.BPkX}�S乬�O��$G�}��O$Jݗ�mn[�E>GRj8~�͆A�%�sC��>�R�k�w�C\�K���7=˚�Ϲ�K�>A���s}���a�ܺ���j��K���Oz�RS���c�}<=Kw�B�s��B�!;�$8{ַ��5�����9:��5��Q�J|��~�os��Hv}�n`�yGo7�7� �j�~ϴ�@y&GG��:��v���گ�,_�K�����0��lL��T��������A�1�:�����D��N�ˬ�����}��.��|�~}͇[�2yi������j��I��M]A�=9��(��9w�i�a�#�Y`������#y&��0G�(}�ƣ����b��N�3����:�u�pj���=�������'Ѹ俭OQ��P�^K�������2��iz���d��������=~<���M�}�qy�^�{D�z�z!�}�&>������.BWq>����\�G�;�F��{'Fg��%?G�v��y�j����w~����{�o��������r2|�;��m�]C�2L~AXқ�;��c��v'*^��2�_b��d�b�1!��8�zx�K�rĸ&.�t�s��҈�5�����n1Z�l�Ȧh��B��:�����Iږ��d�b��������r�^��>&
�ṋl�쾧�������'-�Uj��9�zH� ��4�:������~�Z)�\��嫣���ːl�Gqԛ�*N�`j�Q�?Iљ��L�`��;a�GP��w�?������㪓�p�g�>n�wt�G�g���1����{��^�9'�z��#���n����%\��5�>��P����N��.C�r4K���N��p�k��֐�?Ov�����L��Ώ>�_|m?i����n7�1��C�"G���h��5&���~ךu-�߶{p�1�OS��ur]F���=}���xsA��U�g����5E�:�U?����F�R��?���;���\�o�˟|k��;�.��n7R>�[�]^K�k�/ƺ��z�_��pg�:�K�����u��K�׿kp��O%�a��h���5����2���w�=G�=�P��w�3z�5lg�[�ݿ���3��2N�� ����k��tkp�����5�|�P�]���9�!OO�i��%���?����r��ܔ��{��&G#�9&T��4;���jg|������t3���i����`����\��f��#P�t}���z�� ԝ��j��2-���/�y�ѻ�z��2{z�GRuۇ���gz�BU�/[����	}��uͯ#��\��酙�C�}%K���O��2���7�z���uA�b���wR<�-Z�pk�'��1;�&��Խ��MF������%R�E�`�%�'}y��~��W��>����S�b��
�E[g������^����@ G\�k׸?��?�y��a�uS���@j2>��Wo<��C�2�{�:��B��]K�׸�^��%����n:���\��[�y.T=������]����V3�_�`��?u�Bd�ɨ���l~��)�w��i�����T�������y��ב��9��Q��{����u�����fHV�q(5/�����G��+&�����.���z����97���))�zs�nc�Ԝ�*�}�C�=�A���v={�d���9#P�X����~�Q���7R~�$���7	k���GW'�BZ��{����_�f�jʱ�7�x)�֭�\�Er��AB�NYy&�>Z�|���_e�O4�$�v���R)麽u��.�ծ�P���-\7�����.����i��9(��ۂs軯�;��N�;*p�B�����u7�}!g�T�JdX������7nt��o3�����0G�(}�O�"(	W�����u@oxk����r߸�F�y9?�~ևp��/n���T���s�w�<�>�2?k��?]ɩ�jO�kI�ܜ�I��5z{�xk�y�?_u��y߾u��J���sA���-���.疡����p���N����BWF���s�;�S�wޗa캩����>��K�=�}Υ�y]�5�ר�HP{���s�<�w�����>�7�_�DG}"%��s�����_._��T%=˙��r�өr���MC��5>Aј�x&O���9q�Jo���y�jO�y��O%ᱼ��ॗ�p����󳐎����u�9u�u��|���d�2����I�oy�xg�l59.s2��C�22_ֹ�����:���(9ujJJrgP�5��=35R?G������x&O������#R���;�������V�MWHם�L�߾��}#�xDO��퉺��2z�������ￖø��]@~��Τ�29u-߳�'pj�1�����=������g�w��������F��˸~�=��o�� /]�O�{�5��S�}�� ��{x{u�g��;�o!�Ԛ�cQ���9����A�%R�������B_}͉��r^��ϴ��p���{<����j���Gr�{�V����K�Sվ��;�<{����$}�>�a�<��`���?��|���ߥ�5Ru��{�K���=�W���G.3�WF|�q�N�wz�׫�L^ۑ|��ldQG1�PU�V+�n�^��DJ����_3#>����V2�f�_�9S�;�����ؚ�stG���u����'0;�O�>�ga�Q��{K������:[s��\�b��o�*.$�u�;��:ƫȀ8]�rQs=��;(��M�4�dC}�����\�ۥԖ⮙��ʛb�B^=��2Ћ�����Tֵu�_k�-Q�Nɛ�(K쵫:�|ֺ�N��U�/vo+������`uf���m��,����Kt�|��U�nB��^���|rz39OM��u����r��>��1�&a�Jjpl
&4p$㉔ bz*�j%3z��AJ�܎u�\c�B���@lК�j��9�e��?!�o��&�W�`�z���wa�j�j�.�ov���&��/LƖ�ݓ6ˇn���,p�r�ijN��8��ʠn\m*-pm���Q$�p���P]2ai"���S��:"��놇-W�<�Cd@���}YN���Bz�Ւ��tς��
tݡa4�o��6*���1��u�'9D�2�����iE��:z�1l�M&�@�n�jc��#I+iѸ딏TIٶd��z���ng}A��Q�	�95�n���0�p���"�j�~@��gW��qe�=�*)O1�)(C��3A��n7�������P�y�F�t<�=��,����)��M���]�ws���f�>�C��+�=��
�U��Ϲ;�cO�ME�`�{f�d�v����]ʢ�x;D�n��1
�m�����Vk<2(0�*}����΃�eL�w`£.�����m���;Wr�j���Z��T��\�K�j������;�j{:)��ZJp܅D��[�Z�Ӣ،lم;�xE�a�����#�n�a�h-b�e���* ��A���0w\� c\���mIx�"������Fv�C?F���tKCEE���&3��	
�[��4�aP���g�xKѻ �I����L�t�z:)�{��{�m����(��Y38���{�ڢ���'v��gYъguMϡ�v� m�y#!\�d�9���5\*Vła���L�>�,�u�S�}�5�wZ����WQ;���{2¿��Y5	Je����V_�s6/f�ี$�Ub)h2�t�|^��=���vF���EmR���"Lj�_+�9���i�edSw���9��p���mU���-�}�E>z�<����>��{���\o�S�L}�>��s3 �{�s:��yO���L�j���OI�P �9�8�G�[u�)��"��"pL+g�R�5���J��f�p��;'61Dll-��搛˱��Y�ذ�̬Ȁ���h�4\�1�]|�;�lS�[p���|wS�8�f �uHM|�J�� b`1�Jtme1��0�^Ua嫷�\q��9�$��/xOړ��As�9�`6���؃0�I\D��N�C���fZ�^$���ۻ��mWb����w�f:����/9����Aw^G��hmt��yQ��u�Gz�C`�*�@��\m-�!�RV�aܶ�m���v�[\�9
ҳ�x�pˮ�ʘ��B;l�T�`wi��^���T��W\���7ɺKe�Xݎ2����lr�tn���Ù�K�� �$�lǌ
�4-�n�W��Y�J�A��X�B�S5v�懃�2cc�vh�s����;�~z�idjs��8���#ˎ�������*cK{|Ʊ]jWB~�5;��r����V5'<��L���� K�+<���^']U�>0�וٕ�p�m��	���ެsqyMp���R8u\"�����Cs!��a�B�B�1-�Iwn+)�n�d�jSk�7}ӎ�,򞕷yqa��[H92�����5u�8)_:l�$T�d�����b7���)ԵՔ��я��6jZ%&#~�}p�U&Y8(Z;Bj���?:1����[�d �N��̞\�8S�e�~۝��� Ӡ���`;�MC\��`�S��eOͱ9f��NJC�ロV�q�����+�҅�E}��"�\�Hk����������Mf���NݣvJ�{l�pQ�ʇ�|�L���%�������݋�A]��f<����QUz��N\+i���SF5�:�h��ÁtVs�3 ���>%2��S�L2�n�h��� <�N
i�p� �UT!���
@��*�p����7�p:n����J9z7��K���٣#T�F�u�b��܋Y,�*�uML��/$�����]�s��hZ��W�d�O��&�l/Oy���5���H�y�!e��ZŦժ����9g����W��m�^C��[�L�� �B�c��P�d�Qw�:6eD�Z�H��=kj��ϩ5q7,w���;N' F�[vF\9�f�S �{B���Ύ_��(g�d%|���xFD#ƣWR� ^��u1q�=��Q�d�4�r��nd�7��ƒ.O>��a��e�e��j��֤wl�j WI�}��2{3k$'����?Bx�иL3�
<���#�r���u �*!�oHb��oV�P�:��j����%C,j}`JuGK���:�BO�e(�\�kej�M��8)�nR�1�=��6���d*!�`iy�[V,;?	�����MAɱض�o����]/JlҌWV\C�h�w�ƍʘZ��㐹����?jwL^�ZW(ׅh�P�"r��՛^ɣr�����}7\3�W���3�J�ó�k+~j�%\F�i��}�PDl�Е�������iN�ݬ���a�t���B@r����qZ ۯw���W��X�O;y(/d���V�v!'�o�\�����ñ�j�B��Q��Z������U�o.�.n������b\xn�9v�h�][��)�U_UU|I<�o:��d�e�#����]NQ��ON\v�q���WFC��y�LNb�`��n�'s���mV3�*t�����*�k�T�����)I��9��LT��`S_T���f]yma�C����}�������s�I� �'��y����囧�|��H�����1�����#�4.EĜ.��Es��Sp4H��w���0��i�a�����U��Ξ���/�f.*cr"n�u�d��@ �X6��=oB��ׯi���^
�XlК�5�|y��������8�E�O!(@�P3m.�������8O�O!�#1�#�Bڬeӟ��4Xq�]�w���$�^�Z38�s������[hsH�3fB6m�O�|��
tEB�\4c���.��$�Nrh}x�)]�Ӻ��[9oF`V�"�g���i��Pt���u�oP���&\�����ۋ�����(8Oz��.�*W
��7�-�zzSǄp���-�;�[Ǔs�en�Bi���N-`2*bk�J��7hn�e�粩m@G#r�VD�M�`.^��Ѐ��yl^�χ�+̇t��{�*�e�T��R�����] ����b9���]���k��7�;�y	�@�Ve;��M9,�[-�R��������W�UT���<T�{.oNW��!O���J��M��3L����&x�~�&f���T���Vk��\��⺴U�����z_�O���P�y�F�@s���\ADD��XO��;����0�wNg�����"���_e=�+���^\,���F3���V僽�]s�ﵱkf�����2�wc�:&lt�]nK:���Y��s�jU��鉈<%w?m���z]�v��~F�79+i�5=[���p1�D�4.�!�Θ�ʇ]d�1EC�vu΄���/S�������|U���ԯrc0�e���hI������|l�0��TJ�t��n��ŶJrF�&����a�Ck'y��r�pR�G�G3�Y�q���#6�(Tf̘�z�f`���v��w��8#5�/�_�p|c3~u&�nN �|+�ڍa������vt�w�keyE�k�\u�ak��c�
0VZr�Y����6g��yj�n� ��X�1����2�@�WK��u�mq\igzx}>��>覆�@�O}�"�^���m��&�(#W/ky>��t)��2��+0�(�F�*�+�Nc�%G�'_f�)|Ec.��K0e�w�v`{dP��4
�Yt8`=�:�Wh��Nԑ�v�3w$�h�Ԓ�\�S;(��e�#��m��K"��_,�&� ���g��`t��@�BU�n��No<wK+�G�{��L6ېu@�3����u%�����]Qؕ{㓤�!HGlb�b3�y���6!�I�TXm��N�t�mhʖ���Q���)��];���⍚�c�ЫXz!�b9��.$A+8�����S.�4ls�6��̬��o��Jj��ɳ�\�+1}�eK���2n֖&�m1w(l��#��ݿBw�Y,��h^a��2�2��%�I��D5P��"�����m���wƘ�Y-����q7P������0YΡ"X�:�@O+�I׊�Y�͎�K(�-�hUÕ���!�'Z+@wlK���+Q�Q�y�3����wР㮣�ۆVj<X�l��6`<�L��`䌫YC`F��gQ�ʋn�w
�Á�0�T/�\��t�L\�����v��Xm�z���b����K1�ZQ�Q��]��Z�[N��;h��:N���7%.Sl�=jr�m��cS�yg7�5¶���ׂ�VW|��͗WH�gY�ج>���i�]و�؀c�{�<�+P[�����[+%LFC�;�<=�����˒屍g�W�M�|����΋�W������l��.��'r�{m�,ۢ'O��Σ�s:�F>Y�-���\}�VX�om�n�S]$%ec��-�7�Х�A����^����R��Ŵc��_�7&���F�G��.ݚv��z�mA�MZ��Q��Ոz�_:�Twr���l��%3Yͨ���n�i��ճ؊��bup�&Cuɻ7؆B�`�E����-�\(X��Y�L*���؛V�h[�6��"�5�S���ܘ9���EWa"��o��v�nujA���t��d��"�ǳc���X)w�����&��T�q�c8��w*B�;i�H^K��s�hf����}���]hq����º���KL��TP��;wڕ�U|��:X��si>�-�K�w^l�]�ď��6��M��^힡��z��3����9[Ϣ���5wr��/��IM��p�gfk.�t��;��������`��ku�e	̻\�G{��:6�ιQ�T�c���>�6�|Ծ�T�vP�WX-��}�������zq��9��DdT��v�N��Ťgu�����V�,��	�|%�3�4LԻ������ML���M��g(���Yz�h�H\Y����5o��t6��N�J׭eJ�O�oi��
�r(�1J�3�A{�:;��^�or��b�ۛ��s@�Wv��Wb��1���%����[a����C�}�ڒۨh��5���N3��^�WB����͘w��!�B�.��7�wy���3��v�ȕ܆B#@C�����FBT�J�P�H4#�4�J�d&E*VBJ�H��	��)CB�f)H���&JAX�&�%J2L���2J�
C%iR�
�hP��J��JJrV�2C$
R�!30��J� L�� 
D�rV�1�+!)30L� 2&��hG&��P����Ɓ���"��2�F�$J+$4u����f�5������oX嗒{��T1m�e��q�it�T�6��s{.ܦ�������6"y5M̳��C��G�������<�aGrvL���[���OCC,gÀ�P �9�g�6��%�7�$R~ �E.n���UР�[�ч���,sF���isHM���g7b�P,�kw��>Q�������輺I�A�f�QN��}�>:���m��:�&�L�< �@c��αk��y?wEp��a$wA@��V�Ʊq��t���D6p���7z����L���5u�,1��j7K''��K�& !#�+�_��S:8������s!�s6�yV����Y)��:g�=�yC�haTT�v:�a�e��a���C�/�H��{�F�1o��;v�<�'�5�����e�t)�s��Bj\1�(O�
��)S�Za�]w�>j��ꋕʧ���}=��:9[!�� �i�`_s�k�v*߃r�=��O�TO�K�.�-�<̨|��U�ū傇	��)�!�t<W]y����Чg���3wC�ս���oI����8l����S*7o���=S6�|Ѷ��w�֍����?1G�j/
��#7Vf2�Q�'p	��!.p;�����' xL�s2�Yk�o�RXd�&�C�JP7�k�4��S�� �k�n��Db5��Mt.+|�>�0���_�ޮ�u�%��|誸� .3;)�1�M��T˨}j�m�FW�{�{�{;a�����(����QQI�R�t�q��*S,��\q�j�뎛�v-�x��409�2�]k��$Տ}����%�o�3�;*��*C�Qe��4�1�y�E:l���Z�qu]Z�֨N���i�fe��^�W�XxFP�X��=�5Յ�5��i��2���n�eP��sк��{"j�>r��u���1K��e���QZ�,KW��$?u��ߌ�x�S����Nqfq��!�W�#\L!��6�-��X9m����߇��Z�6�^q+{I�os�:1@�b9�~��F��Oq��^s�
�u��d���k����>� ��Q�U�ͷ��~!M�2���`�kj���M\M�2�q�*a�ӟ/e�=>��{7�%����2�e?rM�E�q�;DLKu�)�!�=�1���Op�Y�W�uL��]M¶���k�W\���|����uZd"JS�A��P�"b$��<��	Þm|�[S����R��d4_r�&�k*�P\�]���>��Y�ϔ(rۜ�����|=u�gz{B�jۃ����]�B��a�bz�G3��;0>����mV
0�n�ec�1�T�gmt�W��a�&'VW9�5��v%�K��@݆)ʔ&Y�0
�n��H�����4p-�Qm��5V7]y{Ӳ�d��[�
ͮ���d=f5����Q��Y�?��%�%�[��������q�?T&���9`k�_[3�B>�m���
�E1K��Z��Ͱ���*��\!�����c��健�[V/���&#��� }�O��zY�e��O�=qa����@�U�z�5��b����	��|�1����is^�`��t�Civ1�ӻz���F6)=��֬��1^>�Y��Ť�YMUD�e�^�8�P������ �-�%���;S�l��	po;i���
]+�!�vz�"�K�c����(��7�hn���1X�! Ud�>|PϪ�٥@1{c��`٤q*���
�]�����\:��*��WE��嵆C���_@���|)�b��'w�M�^�ɬWi{�;�]B�M�;�#�K�nD�}�S#2.Q'N�������|'��s�Sܧ�~�a3Q�]r�?0�Bf�LnMֈj��q.��R
�uչW��D\������I�h]G_��L�
�44&��j�d3�F�eE����$]�H�"3.�󮣤3D�U�����p��m-(��ූ��e�"i����+��A%�8�����^]LV~L�����ᮤ�T!xm�堓`�Z�ٖ��s;�,#xj���X�v7�	Iԡ}}�%�;iwe1�������y{x��f������W�UUU��:����}����|�����΍���j��N~�X�a�-v�9���6�������=�'4�3�S�b@�(�t;��艉0��Pvy���)�����w7U��Y�־ac���wy�(�Y���D�c3nי��Ό�}��֤Su.����Cs��Ϸ0�S�p���S�Æc&�7Z�wP`�Sj�����h�s�5i�����|/2���;N����TjSOBn��2� �}��)֮'�gcű���sG�ݣ}�gḠ~,off��q���p��"�d�&���y�ت��ll�5BI[�;�\Q'�#��JQOa�>�[lVDN������1�>���12�I�"��;�Y[G6��(�E�< �0��L`Bj���͔��B��]6y:�W��:���=�|v�C�i��!�|z�*�
�4M�s����P�T:����f��rH��˙�۲ ���8��'Y�������z�0Ъal����<���ٖ"vVő�(gu��`|j'����N��y�d�6���E�u�:�^�U��Q{ګ�+5�bA���?�r��6���f�Ʃ���Y/�nN������#4;Q�h+y�K���5�^�Gfcũ��o9
�e8�Ljį.'a]�����y/yNv��Er�ŭ��Y$ ���1\�d�"�N��W����V�6x�8oޞ83��	����(�����q��8���36*���v��&�Je��<�����f�������٭�ۼ�V�铂��a�,*�3�]mS���"Lj�_+���7��7��oj/C�v�t���f_PK~�U�Vt��A�Ep
��cؼo�k��Jb��鏅N@�L�B�&��X��=Bр�8M\>��E�?qd��(�dgǦ7-��{��նlfj�C
��Ykz�	\��q�)���8v���e4���e!ֳ�v,�lxYU�r�{���j���}qW��q�໧�u:���9�2�RJd�� c*oq�����[S#�z������"3�Db�_T$�"���yX�n���{ХO���Ea��-�x�a4w�|�A3	6q��d>�mx����&6�.�&Ә�[��K:/o�3]�%���Y�wVh�t̊�`i�3]v.U��6�g٫���4=��k�_;��`�<Ǿڎ���(i��ފ
�!A��v
�4�aX�-�;�lv��o[�k-��d�:����b�ܸڻԆں��;��)��\�Ku�[����Go�c©��k]=gp덣����}��Z���fv��d�aTյ����Z+���&��x �n:Wқ�L+~��0��MO�:DnLX̥OMg�0��O��1�e9�����w"�`9���`Q�p}Z�V��[��=i�ꈘ~���訢i����]=�"�*C�YbҪb19���@p�Ag�B�q2��A	촱�s���9��aL�qJ�&0E�Δ������z�m���p��N��ѿGz`�vz�.(��x�G.�֠t��*FҚ�]�84�n�NvB�_8��'��O�Y���^�*H=l��������Q�N��c(L����:0Ҡ���`;�P�TG)�X,��Ī�Ԭ�]Pgp�h?nK���+�}�f�\#a�C>c�X�8;e��2�̸7���w������<!�')�Ϝz=�T�]�.,Py���U��xޯ`&?s��SH)�9�~K��ﱲn����Q�&ˌt��;�鹩��.O�(���*�����k�[��t�	�:c�df����g���E,�n�\�O��hd����sS�� �cթ׵�劃b����xʻ���+A�7���o��g�f$"�D�����s�	��)���.���|�4̳�^���	U��刑��)S����3j��9�ں�z� {�b�9������V=�Ƴ�g�h)5
�= .����>����ƕf;}��y>�6i�cBE\Bڱ�r�WKǊ�c��rm[vFQ(Cn	�3������ ��#�I)�h�L�E��]\;;l��R0n_T9�/���]od��C.J{�+�ö����j�i��}4.�T1��2�g��l��4i�UOܮIE�PA�N�02T9�)U�q8�U����<�ȻM/r王zPn�ٵ�7�3��m����J%8�偮'��"'�(��BӐ^WۙN,>y�� �!&���8���qNa�چ#�<�3��\��T7,/ -���O^��+�.�[��鿎�&��lrA��e;ְ�q��0/�:ӝ>�O.��K|og��彁D��,ȓ��x��eP���(�.}����9��iC��;+�Ww�xL�o�E�)J˫M���{���P���U��l�
NI� ON_m +q��;닩*��va��s��;�Wn.w�܋�zi�_��3�v�*�/�W��n'd.@x
н���Ғ�tU֞w-k�Κ�h� �υoWp�Jg=�Y<���B�ν;S���\��N7Vm-��u�Ep��IR��9,�˕q��ݕ�n�+�wU�O�Ks��ۍw�Q]�C;��&ڕ�����Ɗ+�J�{e��hJ��Px*=����QV;��}�om�#>���.!�6{�ۦ�Ί�ʝ7Q-�'D-����)2�ǊVOBǎ3�/�{@og�]���d�Y)�퇔�+�\��r���Q'P�/�`k2�=ysځ����ڬE�CC��Į�gÝ=9~ae�;��[�LnM֎�7�o�@MK��<e��Lp�I�xT)�a��W0Y��6hMkV��9�9~CP�Bt�߶-F�����@	G`P<_A�����fll�~��mV3����NX�/u���*N���֫��8�\�ip��=d��T9�!P�x����B�F�	��r̡�s�o9�0��OD_�[w�و`p���a����э�6%���,���ɡ*��	����C����NzT�~���3�.�1l�MBn�N�t�f:��}���T*ۇx�m�{i���Z�H�bW���Ԧ���p>��_� �`r\�z������x��]�ܮ�����0�D"����)�Hmgh�ѽ+��}_ɪ�d�MH�\�GdC�n����M'��:3]�O�ٜ�;�]���s@U���O7��U�s��|��kw�v����^�b��HG3�1�w�`]q�>�8�7w
��-6Y��ǚQ��ֺv�j�T"b�Oe�-͜���hk���^K����j�����ǉo�
@u������N�������d�wGay��r��xS�T䉬�cD�%h�Y�`��v�,��c�Wq՜��)_]x�o{P��uu{�U�u�n�S|�M!A���S��C���eX�Y�D���C��U\]F8�޼�ӹ�n�!�B�N� T^��-gW�{�Sܘ�7Yk�Sѡ%j�s��JF��+g�fC������3���}`M��2��d�"�N�U�.:�E}��~2�iK%`��M.��ՁN�8�ea�vu��7�1ٖ�,2k��_m����^$E\��+(t^��\`u9DlJ��4������~J�l�����ƺ`�C��1o�qˉY��5/���:e4�ћ>���da
9�-�W ��cؼon��>|���nw�U��R|�}����q�>�9p��ʇ��g�#�I���`�2,���-������T[���㧥bĎ�,>yM�}'�Ŏ*U
�Z<]�ڨ��n��l)�3��\x��Y1�Q�T��4�,:'�e��)��O�z�.��uwbSN�,�n>�S�����e�6�5��Ax�;����T�4�[�u�x�K�-"��R�uU�X�	��>Ƴ�p7�t�����7�������mz��Wm��IJU�2�v����y)Y��r�ӷH����2��W�)k�-�p|wS�M�ق2�RP�J��t���m�W׎Z]� �����Z���nđƾ�ƾ��$C8!����n!7zL�
�Ⱦ���I��Ϭ��;�Y(��% L�o��p���Lޞ&5��%3!
UHֹ�u�Cw:Z�nvjX��6���Ӕ��40��o��a��^8xn���ާR�
鼼;�۸s��t�r2$�e�I�v&�Sg@�Xhd5?��f*%uF�/5w϶o�ɼz����D��C��܄g��5��}P�E�Bju������Ef���=`I�\t�W�z�EN�e#�a*�!k��r��X:i��?k��7����mh��kE�᫄�e�WT;��H���3�e}�}l`!ꙶ���Gk�E�s�l)ʒ=���u~~��B��� �#�=6�;�h��+���%Re�����bΙʔf�ܥQۯ��=q�Sg���ԃ�)�:N��Ҡ���`=A��BYr6wLÉۼ������针��I��gs�=UAru�Y��65͔���h�KzNl��-��`c���r��я����ӆiƞr��g�WEN�&�G��(ṱ�]vjP	�$#�
p6u%4�u�����v��N:�|���[�Cv�G�tN��;n�v�O�N��;�e>����q�L%��N=���Q�h�8�x]�	���WR}ъ���G�3!��;czq�T\�E�]kh��о�q�ə(Z�]ט�;b<�� ]��lF�\��͡�$��y�����ΑLoNe]�Iu��>3[���)��K8L���7:��b�W!([��z�y�&]���C�wuajWͩ���2��3,)�.�bt 8�R��޽�:g8���H�ҴT�,���&d�t���v��Vz�V-�I�,E��n%�U���M�����
^�Vkm��_D�>:j� Nk@���r�D���#���	�h������B�+��.W<*�u����i�����#�80���v��N���Y�w.�o:�JS�.��yƤ�oZk.��/977tK�R�=a�\u{�(���O��#����T��;m� ;��}�%�b]/�v��k�S�2���Ү��7�b������O�w�ly�����Z�out��
��-☥	=�j宲�f�I`�R.� �E�gX��QX�k����{���e֭��k��CR��-,@C}��M�Z���ʚ�5���/2<���X_,<��;����L5`��"��'��;3d=٩%c��k���P�Q�׍k���<���/��\P���v�]�k��~�y|���-�(�{	�ب�S���
(i�/(Jfwho'" w���Z];�)i[ص��#4k�,�za�@�q�܄^;��b�:G�] E�O:�u�B�|��4��޵d2�2���׫�3~��>�~����]�Њ��+���4�#�W*�`���E;�n2��Z�����x\ﱩ�eG�v�k?��qq��G����[�Zd�`��+WP_Z�K���e!N��b���3i�Ÿ $f��:��h�{�EHxCQf�9nT%�%�o�T2�w��	�����&��hk���:5��U�vBMs�(�ӝS2���v7��xZ=қL��wǶ�r�+y'�Jy�^��w۲���w���C�hU즟��b�� ���x����ai���Dx�o=[a�k#9��w,����Ye"
޷�{)���[�!�;�
�{f�Pf���S���$�T@j�V��:�w�r����$c�����l���&�u��u�v�VK9����._=�$��?h��ܩ8��=�%J�q�Mޙ�^P��r �-N���N%Vq*��8�]b�J��{}\�=]�Ci�9{y}V�
#�M�[���Z���ך����$K����.Hd�A��(dHeA��%J@��R�Y
QC��ud.H�.B�Ҕ�H��IBD9!��M(ґ	�J�)P,CH+M!BP�Y-.Jf`�4�H@R����A�IBdR�%LH�MST5@�-��9.�5@SM4�%J(��CL��(h���J�$�����K@�@��-A��d&I��#CUH��PRVC�Y�d)ߖ��]߻I�:T�F�d�כ��}�	�����NV�ňo�a�+�>Ý� ��u�<���3{o[���.�����%���y߁� ��پ�0K��v�)^�f�W
���G@�<#(xS��q힧3��U%���'2�8�p���x1	�g��p}�o�T.ʔh@���A�� �i��#��l<u&.6�(�IVK�c��؅�[��a�t�K�}�JO/m��\�0�5�*�}6����͐�|J�b���énL��}Y��<�f1���{�#T����5y�.�yk9y�I���)l��=�&�${�F�.�#e�ƃ����U�f[��]{Dr3�x�D>�8�J�&%*�T���_��ò!S��Ti �\�[��KӞ�!��(�{��F���\��S�-}�b ���/���e�1oQʠ�,�pc|�].��4��!�Ֆ`
d����T��J'hL����"��7���J3̻��=���W�%��VC�Q��䩒��偯 W��PDO�Q;@�ZC)D����<�m�.Uܨ+�p�َY�GB��Bj�M�1�l�0��j���߮��Β���}��>�]�}2S	�mE)�ud.���J���w�GW�>rP:
�D�AQΒ���~�V����Z1cց��ݜ�;��+y�$ݞ7����N��Լ�����+_&̶��f�I��}J�V�#�o�����%s�{�:�57�ϑO-��tZ�~ô�����KRw|r:ӝ>���)Mp�t�]��˿o�c!H=^>��Q���65?���Y1�^�*�����Qj�p�\��ZXJ���92�8N�%\lU���$�4BB��E6�=A�gÃ/��=���+op	�2Zm�f���%S�b1��=�Վ���1��t�# ]�\>���vnT��纠�5��}���O��c@����22)'�uM�����3��:���ϡ�}��ǭ�4�ݢ&%��w���K�p��\.�gPdqwc�-���LB���9b߲�3�j��՞�l�+>��"��NN���\:�!���#ջ2���ON}��c�LÞ�1˻U2���/�{!~xF�8�J��W�ipT)�a��s����SӬ�V�rﲻ���;ø��8����%ޫ� \{��{DO ����R�.��bQ��ۯ�v%q�;�c��F����B����#�ԝ=d��S�B@�(�t7]Q�!#]��qo�`{�_�լ���5Ѫ7�C�8o�׷��ԭ����t
�t�����D:�j��'�Q z�:�p.B���{����Y������]��vB}� ��V��'���P���Z�!
�+���_u�K���z^���Գ5�Қ���m,諅�*������M�,�.��D_d���5Xy���u�M�w��g�F< K>�©��+����XjJ�H��{sv�5�u�)&�-�&.������Iѣ�[W+zO��h��?^�����K���2�u떏VBW���j6ҨrSs���0��%7� m�3�cճr�ɩ2�J'�r4z~����U������{_?�UW�'�4hJ���a��6�g|���;_�]��bt�WF�
t< �����������s�ly���R��pq	)��I�P8��<��� �0���F<�����V�LU�B<.��I�ǂ��4\7O�3�N�Y��=_eX�S�qLp��{>���%�jS�F⻚�<]8�œcˌ�`
�U Y�e9�a����9��ۺ�w҉�	\���E�{;�n����N�W�<���3��Ȓo�<��Ja�l��y��s��(�ЦY��0z8�[�2bC&�'����VΑ��U{����TK,���)��n�c�"+^�0'W!D��+�M-#�U.�S8���L>�v�N����c�'],6���y�e��K[*�q�[0�E���l[�����p�W.5�.��Jyu�b���K�
�ڀ��4p�z����ڵ���Viu�ݷ�촇f~����FK~��hGN�U�X�Fĩ�I�4t	`��%S��4������?n��|�L����y�t�<�s�IGt��
lZpQҸ�r��\Ǳx�q���|o�D�bt��&j��.s+,z��P��HfC��|��}�m�� P��G��dٜ�̒�nV����6��V*�sZ�}�޽JF���MN�E��A�Q��H��-
��[��Μ�,��c�m5U�����������F�U�㺝p�m��N�	�x�=��F,��kS[�&� L1��S��+�ݒ#8�.���t�������ex��]���r�{�� �g�I�J!��A3	��e��[]�x�0��������ަc�|���.�V�
�����>O�A��}dSG��gh���b���6��Z̠F��<)Q9r��ZҼ�l�5&*N�'�Ε���ǭ�FhXhd5��c���鴮��XwG�v
�����!��ƌo��B����_Ȱ�|ܰ	�l}��hX�N՚�T�3�>��3�w+P������w�u�2�v!3>�3x>-ST��Ew�e�t�O��;��.z҃W/OX��p��8�>�T��v�$�������)���yK�ά��c.�ɖ�yz�}x�XU0:�oV3Woa�y<���頺6i;�5*��D}���}��Bx����7�,C��cE��ťT�Z�A�X�,4�HY�Ц��k<��9�7������C{^:��������>�X2��g��7]D��wM������U�J�sC0���f t}Ӂ\VUi��Ox�X%js�WR}��v�,bڛJ���b�����8o���3��9).�	}��?C��cܬ���,���lʪ��ON;���ݖ�>�M�Ϛ�W���ziـ�b�W��\#a�)�D֠e%7b�%��[����g!l��5��R�鈴�3�������m��C@V*��x��6�����v���ډt�w�������c�Q)]�Y���F�5�u����O��R��&��we�,���k�Z4����G3Q[M����Y���?T9T����3q��zoQ~Av��7��8�:�壴���ƮI�� �jK`)�"�*�mX�9I���2�q���<z2�M�M�fv��S@R��ބ\�'�$�[DiּșJ�6S(F#Ʊup�YbZqח4���۵J�jq�� �n�av�(�F�E E��ue�2�綖f�l��e��'+^�E�U�)�}&��OȾ6�Eg#ein� ��{
�r��J�r}'��� �f�v+2�z�����L�f��*q��pɥQ��Y����*�'����{qt�'�lK�~
�4��S([��]ô-w7]����H�1)�:��6�/=�\�W�۹���S��k��j�.�W�u�.\�:���[�l�]�ӿ6]j�Om�B��u���A�TC
�?TrT�y�5��@g����7zT� /�N��@���x%��gMl-y]oM-�B*<�3��\��Sr���ڱ=���ݕ��Uj��5�t~N��c���Xo�o��Y΃�N�v�ۮu����\�Nq��5�6�*��"�;J#�����W(ׅh_�mY��M����'�gxP��f:��~��L�竑]�½^��ß���4�1�W
�$�f����?���g�����pSp��їUz��ѵ�Ro^Cʨb:�G�!:�ݝY�+T�F ̨3|��|�v�� �Ltv��c�b�E�kh7�������H�G~lv�n�5�����8�{�ݮ��g$V��f�'�	�����n�K8������nu[�#�%�;>���IwV�^~t�X$�Y���ռ�£.=NjgX(QU7�+ �
\��6��nw��:@^�u�b��U�-8��X��#\��!k����'�^�>Y� �����=m`���:�D9�G�C��V�u;��v{�v�ӗ����ըAT���{˰��i��$�_Ih�U�mL944 Q�Į�gÝ=:>aZ�p�������{ ��,Mj�u��8�c=@�ii�IƗ �{]rԑ�:!\�f�f�ֵo�{=�S�UEm�;yj+���LRk�!�-��M"��t_�fll�~���c$�ӹW��C/1�ǝԾ��0s�K��r̕O�ꄹֲ�hsH�3fB:|�jρȷ��F����,�z���~z놌��W�e��n���n�����F~�K2�ω�Q6��K���RC�דJ�=�GU|���$Ҹ���1���t�M�5r����N�[N�Q� ��ڦ��l�'��4��D&�;�\c2`㒚�Rʝ�^�t�k��W��U����Gg�s��>��{�*�{)�ݽ��4���ԌB�	k�5�uZ�Y��ۑ%���>zg�z�s��a� ���$���N�޸sm�ߛʭxm�xj�л�����T��2���'���ӷ�EyN��e�sm�3+7s��9�'Tȉ�����dY�rS��gx%̀���g�۱�@}�p̋��w�#ܻDEZSz�Up�̎֍�1� .�SK�ұ3��+�Z �ޡ�Px���ջ�@s7p=��	\s�em������ɵ[�nҗ��kZ�oF\�;7�]����t�(�3g�eWG8S=/�[�%�ˌ��c�je�8�4��n��[�zUlh����b�Z�����\�K�nr
c�
�����JM��ko�����f6���S�
�;�w�rX�
�ި��S[J��talW$��t��}�vD�T�oEv"��Qd�DSf9Q��F҂��Y1��־%�MN����WTbe��|Zy��c��U 4(���S�Ŧ�K�2#r����[x�b2�wh��{o�YoB�M=�4�
1������cd�W]�o;��*R�/w\B�.�%�5���O�mD_�[�]�1�ko&������%ٽW��Z�w�nA�b�Q��̈Gz���-�\o�!=��1�ٙ+�=;�v�=���-.�o�x%-5s̄s�q̈́�W�y�������!�5���H���LWZ���c������zzoaS�%�Coq��̮\r���F�Ϋuy���}�i�n���f#[�G�=k�R]��ٵ����jل���r�̀���Y��$���~R�6KK�j�`u^FZ�.���5ͩ���4���4=mdS�g�B��JU@O��'�n���|wy�/�����F���5|���.!� ���Y
Q3�l�·\�Z��G�aL�ݹ���ϱN�p�����o����Pۍw��9�kk��J22Ar�WN����N��J엚��U��N�,p�p7�λ#��]��j�lky��kO�ݡ��?Fg/4���I�/n�r���w':�Tr{e��A��ڵ��^��N��R��K�[���'�E�޵EMT�]��Yۺ�_S�d���k�b� ����F�g�{ï�*&/�<�ΧG^Y�+�_!ũs�'s~��H[�>!mOZ[����	P��[�ν9���X1.��8�8g��ͅ����Wf��:b��J�
��ENP鷧�*��}�b������]+�b�X�M��u�l��m����M��� yV%玚3��ݙyѰ��G>��=J�6�z��S�B~T�-+m��B�(w5.�E�F��.�-�h*�d�lw�]F�I%���[t�H�u)N����Ce��2���Φ���Z��v�p}����27��8w\�y{���&�ܡ�i�4lN Z��\��Ws�;��;�'e�WXu)R��syx��:Ol��h��UX�<N���.GEʢvRJ�������[�K��<`tK1n��>,��+X�����I�ԗ|���"S�P��8���?�v�����gTm�jQx��QQ�D)���0ѣSY�#�{1�:^�q�Z�3���j�{���+5,�0Rlc�/\Gk����Uǥ��d��Gӳr��_8����"�=��5p��aXy����)p7!���ν��{mNޚ��훎�����5��}�W���6�9;UN'ڹ!�6�@ۘ;��)��f���<v��K9�mƺA����w�8�sݔLӯ�ȼ�s,�ڴf�y-����s�9�����|q�'���V�o9Z<Vf����[�O_�V�{��l�v�������q�}��liA������Z�H�$J���-m��(�� з4u�i�y�8��C험h^m
iI� aI��{n�g��͛ԶG�Ԭ��4��9�KŪ���L�)f�O{#���zz3��_#�.��~� ���&n�������:rH��\2���rV�>�ٶ��1�G����ow�WڱW.Vh��V\�h�(٩Z�����j�K+*�f3�Pg%*��7��w&(�����Pf�]�Bn�ײ��u������:�4u�Q3֣\cߡ�KYd�i5J�kZ03Goh���u�H�
L��X++)k.�����'O�a��dѮ�؝<Ӯ�=wo��t:��w��쭉�׮�3of-�io@��\��� �e������Z����ӆ3R�^��4�h����יW3%�8�V!Օ�b�6Z��ڛ����hS�Yݭ
�Ra�f��2�iP�X[y|�]p],ܞ���m>κ�r�"*�"�nQm-|7��d�Uܾھ�,�4��<����y�ص`E���#��M�# ��g����A�m��J������ms���"�J�6�؆�Wz1��>�X��N]������:s�";�Bn�U�S�v6��0�XQ�o"b9:�N�h,�O�f)�	3�B��O2�j�
2�<+3eJ�h�&�L��`���-Rz���,a$E�����t�*ya����g
��y-T�J�XH�y�e2g ���W���v��=���3�6S9d����^es��T)��tuIF�ΈT��Q)G����F{��P�ڽ#o���5��ؾ��(M��0�f�n������M�uNR��O�5��ؒ�}x���+����w�vo��/4��Q��n��Q)v�J�"��U��}���u1��
�s���5��
è	�}����㋆�8l�}au�{���O�S��А�Q�y�\y��.VY{��-ή��+uR�]E}�����Ԛ�}ٻ-��-�{���;űP�S�ǫ�j���b�6������諲�2�7�wU�E/F����+�Wbyq�x��˦�r�^p�U�[�u3����MK����!+jV����(�j���څ�ІGҺ'��qG�Rq���c�S<�ށMr���nGN��yJ��ٷ4�*�9׎Ky����1���*�ũ��+�����
��%��{T�(��*����_.+��y|�0Z{E��եB�G���;��wn�%ˠ�< 4R>\1^j����.�:�E�W��C;���Бf�o���H�|i��Q�6��Wi{I	n�sz��`h�k�`�R�<K*���YD��Ve䰭�mj\�'H���:Ϋ̻��t"[�̜'ew]HdYKZ���JW3��ݮY��� 3[�'D����U�ZЬ���V��oiBk{�V��n��HJ�r�F-��3�f��E:s6���*_d��P�,il,����_=ḻ���IQ��P��@VY!IIIBQAIM	���4�Ҕ�d4R4��:�)
��)()J)��"�r�!���
"hirM@j�*u��Hd�RP�C�d�@D-H�D�AAIA@�&��V-%*P���P��%D4�5DT)KC�L��rr�������P�E-(Ƴ$(h�(i���F��*�Y�CK@P�)H�1��E+�dPfRa�IED���RS�&ERU1T%FDUMQT�����������=Ou�8�J+
lS	[�!��|]*H�k{�p�Z��h�c4u�.�nJEn2,�"�_T��O���[\��zup��g�R���-Jx��ɾ��K��Jg4�RT��l�{ַv��^�|���C�}p�n�m�9�G!�_s{u��3�<h�R��E��Ƿ���V|gOY�޳^�z��ktY
V'3�qT�@T��^ɗ��g-�Tr*��uM}��+��^�DZM�So�_>K:�g�2E;�4y��euW�[��mK��PF%J5���P�I�:��<�MY�Pvh�v3{�����+���e'�+��%�8'��{jq���\5��S݆����|�J�(t�Ϧ
�����-�|����yM-��\º���kzj!��Z�d>���2��Q��ﻤ�2�Cu�y�����G��f|u-}���9�q��V��r̢�i�-u����o+����G֬�zr�v���&���;f�M�
+3�j��Tt�5u�_�+����}CWU�gpU
���Q\.豮���Y�m��j�I�,b�Ư#�x�ZW97���� ����oE7x%0�1ʖQ8z3W���Q�<f�����6P�⯮r��26)�x�.ɝy��zvz.��tv";��NUC:v��[����zWd���֎��{�M�{/Uu�\��[4ݪU�ȗ(����:�s�ͣ���y����z�����zӐ���ؚ��k����vD���{/>�Z�MP����G�1�oT���ۮ������o*���:~��f+��"+��ɣ\�._��u��g��^ܚ��R��8ֵ�ތ��F�1�:�>H�d�0��T�/w�H&���m�	���V�O��<�*�Ow�l��qp��R�`�������{�O�{yҊ��aQ1|����.��J�aFP�:��ܭǭT��n~���������w�6�Nʆ�K�X[��2�8�ܫuFw�3��Ro�vmþ��l�7 �U};,��J
����d�T7��ҥ^q����yp�}q-=�{=�z��P|�=0T���IeuWtLut���c�z�����1�Г[a��|�Mm��wp�K3�M��sc=�6&)y�u�@�*M���׎�/M�:���Z�	!_޺\:����]5�~��|2��:��)i�y��RӰ�*� uº��*���b�I@�l�p_��R^�}�q<�߾wgk��F����>e�=k��ۃMW�(t���,S�e]_+H��t�j
�45s��]D���O9�Z���u=��ܻ��sX��2m���z�]��	�<�b;������S���-L�>�*�ѭ��5'��|���=�R	h�\�}�Tb�	4�h�-����6�rW'�Q�m0�CO"�t��!uD	J�h%>��]��S�v2h���-���U�q�x�ɾٶ+��(�[�;�6*=�M�齺��ж��ܞ�d����ke�'�j9�&�q�¸��27�]	�ɚ��ϋ=�f��]"�o��}�y�WM.NKX��no<��xE�ͫGx��y�}q�#x�>Tm�]�y�/^���w&��/��r��{gN�a�;4�
�LuTM8yf�d�-:�f*�}`��N�+�E�"%S
�0̀������X�
�h7�ͥb��\q��={���	v��-7wo`�6Qb�jٶq9��o���Wu��.ع��oj5q	I�B��[��t���Y��kr%u���L��5���z�z:�.W�݉	]rP�=�_t��L�w^�G+�ד�F�;�0:��U��^O��u��uc�����r�r/5��[����:���k���ٷg+�̪����g�"���t��5����F��q��e9\���u���Y�3�r��Y�ꂬ>��j��87���n�渉��Q����t��-���������=����Gm�; ��|]9|��{z�^�"i�/�jT��bR�c��pը�i���k���o�_?:����9����h%A�Ғ�tYoN�S��o)�cV,�ͷW3α�B6��C*!JT(w|� ��b�jJ��qO�
���n��S�$�+o���;\�cZؼ�ţ��!O}�0X0R�P55��ec�L�������yW��n�\)i\��@y��M�e�D.��@�*3p�H��&�Ջ:�XR���[��[�����桾C6�\x��r��\�>g�X��a��L��^�,����{������>�m��W���Σ�U��]�dJ�i*�thaX$�.��A�WSn��YưT�uQ�-f��c�	��l��*�̨짘:s�:��2���|`��α�<��Ap���������LqW[�a.����7���B}F�&�.1��x+�����2aN��wT�i]�!� ���J�ˈ��y�W;|��_,p���ڒ�uj��fcy͌���*eG�-��^{�Y�Kb��Z����s����ߩ��Y��
�E��yyI]<�1�ڄ򫝛�;~����m�}Դc����3UiЪWd�-o�^%�V�퇰�IԺ.�"Ԫ�u��������Ɗ���4㖧�	�q�+>*y�����kg�^Q�gZJ����~C�0:��&�UD���q79P%�u�Q|���͋�M���ۈW�����;�ot�+��kt�u�]|]���i���J�.��lU���E6��7f���;D�
���;����9�������s���s�\�_���Eu�Uh��T�q3J#�}q-=���T
��*�*��I�������l4��^���ۤ��{�U�-p��Ѓ8��վ�'[�]�ȋة^�qӟT0��տ1,V>��Q�t�\m�ꈌe����h\r�4�Y�NR�C���<9��&��媹�=�����q/v��Yo��"?sn�l�?��W��o^*�Ę�v��m�m놷,�|�JZ(t�|�/���.+T�2[�9�����p�g)}=��Vֽ���Q!w}�A��&�K2��-5;��He_���,��k�rҶs^������Ӗv��f��$�5��^=�����'�����U���$ҿ�|Ž�;pF����[D~�_{�����Ş�|�E�Z溗l������ڄ��ȴ�*j�SѮ��%16���a�L)D�r0
t:�>+rj.����٩g\-ћۉJMLi��c�YJ��t�9��MƸU9�C�U�{W�ۑ,;^wqyqgt98�7��T��[Z�����_�\9�n�yU��7Q�t�]m�4���,T�<�:j*�%�nV�ѹ���6�����Z��C�.g�vn�tj�J���{L�t��^8<�1���+_��+>�S/O_w�[�/}G�,�de#�ƴ���1s�0��Q��\\�"��Gu3trm3��ˣ�x�0�mЦܥu��8��Y�I �Ve
ߓT:�"u7��*��&���×L��)���vS9M��t(qO0��n����!�'mӷp���B2����[e�A�"�L<y"�������Xqm�z�AE��J����s.L���A��J�o��͛1UL��χ�s��~i����4�R�!gCh:{�;��T��Í���~}��c,���o(OeX}���^!+A|�ձ��V�l�[��E���`��C��Zi�i���=��У5��]D��f5�[��vV�|�|�i��4��޾Zz�&��ƚ�:d�]��O"��4�6��:���=��q��]KzjO.9�\�^t[�/쌀՘m�ݬ�[�}��[�C_˃�,���fB;���t*{��ԌΞ9|5�֚g7S�QF�x�2�"��%0?�U[���a����H<������/�F���*!7�N�@.�)T�L�^�6���x�=�'Z��M.��Zu�g�7��L>��&�g�ـy�î� �os�Ԁz���I�K
�F�~��].�k'Ej6�6k[D�m�7Z�-��^�.w�Y��>���(D�1�FpV���ZT�i��;%n��e�<�X�t�o����)��r�`�+��:��c�p���%׽#KP����I�����+l�wW\8��ٽ絩�_'�y�'������Dr���خ��7�����-a��X�e��\�o5j饼�X��ns�Pp��gފ�yǦ�S,��S�%������U/2����x�7*��R�ָr��G*ݹ�1�]#:)��>��w�s)B.���_*���&�P��/9:����5��,�٘�V�ˬ��uqp��p��fw���3(����TM�P�������U1����i]�x�e6�j]��>З�֕����6��%��'�:��K���1¡����6.%����Еo_�6�ɍ�a���Mb�ײnS��F��%c]+�إ��M�Q�����y�ˋQ�&3�'�i:�S����w�})R�n�1�Yq��X/`	�7SUB�{�53ɛ͡C�9�T�TmJK�u-�=哩s�m#i�mм����s~׮�B�c��'��t��K�-��n���c�#m�ى}�+#`8�޸V�x��Mvn. �5y.�x� (��5e�b�M�]�q�ifh7uu9Kc7�޸_51����\�ez���v���a�p���D�=����+Q����{�x���͉��hc���ڈ��*�:�}%A�LF���[t0�CF�������%x�Ά�m[c*!�(�wtAKGnwdOR+���Ǐq(X.��׏��KJ�H<�I���D.�)-y
�B�P��Hpz�iR�6��ڄ���vͰ�<�R�^���[5[I�93g6Cke�#���p{T�].ٸ�N� �>�_G$ÿ�q�e�]QS[Wv�AR���\.ɨn膆���«�
�ˌ�{2���o�ҫ�̊A*Ĺ*��Ωug�Ϭ�f{�Ο�������Q�GcǙ_e-}�����-�*�QS�r�Ė�S��]p�Õx�mByU���k0-u@�U6��<��X���]ʫ6�SJ]�ڰ�&������N5��v��ѥ���E3�f�yo�4j�m��a8S=nzv�����O�=�^��k���Y��!7Y��{��~�X����5�t&�]j�O�5�&�3xH�9ND�Or��"�YëZx�w�����IҼ�L�]v.ܚްcj��>�;��ߗ1	fl�f�ù��o�N0R!�Y�����2���k���b���	bvk�u���k;}ՏK���nK�-OPG/�mD��	p��b��̕���Of,7�ћf�0�S�=(�ڷ�Bڭ�ɿr��3���+�=VRܖd�3e��^=�펧a�oW�9�z�d-��۹��Ƽ�,�}˄�����N���o7Y�WUK!+q�>�i��oz�P��9�|�\D���˨Y;�mc7�Ův*ѓ�%Ƥ���[q����m���q�>
*ެ�|(r*�Hou��v����9[Z�^;le|�*�A�k�B)g����|*�s�s���6�_mÖ��9�[��[csb����Gb�ՙ�)/�s�/�Ɗ<�kis܄uR�P�J�7��1zb��i�yM��i�Yua�[YȄY�*�h0V���]�ܚ�Z;��a|�Z��f��f�_�Z
��\"��1@)�|:��&��ˈ�xܲ:$�[�,�l�].bq]^�Z4�ȫ���t2:���i{&5[hlW(V�����Jgms��
�3��;WC@;K�4.�䏒]w-�]
U'ʾ������޹�+��-��hfO��8�RI1we��םY����tL]ƥ�|�n2� ��nj��g]ۣ���rT�7���n�8V:�]}g^��!�˱,Z�7�)zz��R��$cW�2)v�upd`pZ#x��M�\0P���{έ�X���fmT�o;yxUs�SV
	���3�-,��[qu[m��ŧ��TX�ޭ�ސ4q�8�nA��7TNRz�*�j�gWq�J+���VUܘ��_Q�k�կ7�,�P���;iW���C'��.�О�8;Y�����r�R��>{�?�O:���{_';��E<h��������u��wZsbD�,l{Y�6��wn���к��P���j�H�r���L�:�גb�ۤ������)������lA�]3�Iv@��5k`����L֐�I:U��q���F��Pbk��gwe�%�=�@(G�3/R���,�ʎ�Ӿ����{y���,�Qш!����;�}˸���/G_w�������|m��Z���iLuY�H]Ͼ�n\��
���0kӳuڮ:Z{�ڏb���K�R�8��y�5�5|�������X�Ϋ�\+N���� 6h��s={�S$�a�]�n�S4i4�egív�w�`8��u�o�U*f��U�Wd��p}r�ˠ���޾�X���h���Or:K�����.aw����x�=Ov���Ǚ�ceԛt�|9��VԆD�!L�L�|�wm����匰tg7�����-�ʈNAN¬�˅���f1ն3����}r�N�*�{+i�\�z���nb�����)tα�ު5r�ߢ2Ɩ�֕%��v^C�\��J��4���)�9�(u�&�+�:�_i���[�}m���%�Z����f���k��x�1Wo�'ܖ|���v[�c�[��)��}L<�KD��
�v L��	�b�ٮ�4c�̭��� �kp�ut�X��j�~]t4�Sq>L���/3����!j�%h�vs����\����I [�ò���Ϯf�HfU������F���%p��x�0��(�jQ]�Y����v�� H�q]��:�cx�yz~޼�1dD�����ۨ�N��*S�^���]V��V�V<�(ŧx����ƄXa�(��4+k ��/���=��i�D�����޴4tDԡ:A����i��- ^E���+k#ɳ
wQ�ef�ruE5Y��b�ӹ��4�3Z�ӛ��z�4������G�Q�x�ΥȽq��J�������a�Q2`=}���1ve���wk2<8[�0LX����)�����4�r�
!׵�qϘ�� �%e�ok��X�6��� �n��pg\���9:�\���I�*V���/r�=⪨P������hj"����2H������(""�!���)���&��)� ������*����
�((����("��������*��3!�*�
30
� �((����h�Z(*��h���$�*��f(ij��*������($�))B"`�����*�	�2������
�&�J����)b��*������j�Jh)���j���*
����#
JF��d�d��
J����&���Yi(J
)����H$���*&��jHb��*&�i(����b*��
R�;���Wh�g��~��Z�Y�&�fU�a�/tVH��6��f�ђ�p�s3V-�R{���o�I_q�e���+9#��k��z����g15�n5��Lƺ"c�ف}��v�k�]�R���u��4�S]7���U�Ns��sQm�چ�٬�;�G>�0j�#��� !S]��Kf��4�{i�>?wg��8ֳ�t:��&��U^�ে���S&[љPR���"m�|%`��Q5��x�'�k��X��U��f��e-P6RJ�����.}�.�9T=��En���TM�ᘜ*�.�S�+��fy6g�*��VB٩�p�/B[��8�Xsi�*6�5���Fၚ�*/,j�%oi�l��4��6��vm�齳�H��bշyh����i�B��ˋ��NA���F�:��O�%��og��Ju���*ӿ,՘��� �^���y��Q)Q�\��k���x�,pi�ع���'�QURo�ܽ�1��6`�υ���EԷ��-<�mk�x3��uI��R�wJ�7^�G8�eLڬ�ղ^\�g6g�ܶ�8��1����砖�ؾ�����X3�S3A��ŝ����l�X�1n)��{2U%x�aJ�X��̴����TһF^TW10�Z��i�x�rV��Kss78�������"RG��yX�&��<�_{�&�
1�>����P�k2Ψ���o�ba8}7q�*b���+�鍙�m��(�!Lw�LZ,j��y����F�rG8���;��4��Vky��ƺfQ�JUA��N���u���ѹ�nZ���/@��t�߻ޗ��6ÿ�ȘR��!�>���]
�V�N�:�ک�^��].پ纙|�Q�I�m�8U
5� 2Z�f�ۧ5˗$�gmc�/>�Og5g|��_'F�c�5�O�A�܃W�ӽ�i��"~�s*�:J<�[Sy�'<�����@�ԯ}�Z�ڇ��$�]�㮉g���]Mqv�m�D	X3�3"�F)�u��VwAnuA�vEsǜ����~*{�����x��ΔW��c��qݰ�w�1��S�;����C�]6���fݜ�.ª�q9q����/��,B�DE[�a�Ed �8l��u�gR9�bu�I����n��^��:��j��-��v@��c6Кr|��9����ǹ�zs�.��T��T��	W}�hX��LN��/!;5���k��cAF���m܏yxs/������W���׫�{��t�����lL����gv�y��u��e!�i���V����҄��W��B��\&�9�k��ʲ���׮�
�_��O@�G�@�<kS�c���m�}ᬻ���������wX����/�-��
?s�
�-���WE���L����]s}�;_]�>�oo=��|2��P(t���*�&*���\������ܳ�0q��{�k����۟Cc6��Q@+ﻦr�P2�>�1�gXif�̈G:�w"�_��@y��c)�(��<c"V ��j�;S���q@��u>{��OxmD%�[/�b�]��ج���8����Jv����t6��9�].پ�� ��;�0��#��}�|7�h��WTn���.9�����[�q��f�3V�.xӫ�-]�!̅��͒Q�]��G��6�*�X��f�=�Q}��Hu��!rF��z�r3�Q��^MJ��<_:`�����v����C�	{s�S�J�34F�ޠDܬn��eNhK���@@W�ͬ�]e���_T�JV�=��NW`�����o��~�8�����y���Y䶩o?G8����#]�,�J�V�䯪[U|۝�Z��}�WӖ���O�Q�������n$*-��`wo�v�W�;g�絭�4;<�w���zh������J�.F�bũ���!M�$��	���}�����:P���j�5���/6��$Y�]A.����M���z�>Us�%C���YJ�Ö��vط5����u��w]{���*9K���휔o�\����SQJ��=a!�N�o�i�Cv�zg������Ro�%��[��r��0y�<�K���|}=�˥b��=��OC�T=W���k.1����7�B�O 6J��p�O}ηz*�Nv�k
'�v8wG�S�_kOo��m���E�[pi(���>�L�Quە�9Ԯз\	��OӸc;S[X��鯋}������le9K�t��)��t<s��,wV���[������\����U�A�����$�ɡ8{��J�7{u��r܃����w�o��s �K\߹�{�3����h����`=���ޥggF�N���Q��ԓ�n旴�ZVP��(<�\����m��+�}���S��_}gR��9i\C9�r���9Gb{8�ڜ�o�F78gH������{5K��:�o��G�hU�&$b]�Ki��T�oECOb��3�"�@K����.��O���̘M�{�]Ϋ4���pˌvDL�!�
q�enL�-���}ϻrnwOOl��p��������bi7��tG!�/�	����e\ֹky�6�[KԶ��o���յ��ru���jہ��UF�7p�,c�e�%'Ws�#]��s�mM�K��{2�����S��*��%/�18ֳ�t:E�`��&�=�x�d��/�n�;�e�]�X|�r������ٞ\"�;>~�=�����|�l�h�wN9V����[�u����>�N%W���:�D��A��񚛯(�o�	�z�g�rr�xYu�U�޸�tL@z�0ܿ���gl[AED$���h�;�|������uӫN=VT/�Gj��*�#G��N3�e\-�֘I�1��V0z̸�\��y+�Nt��-����k�E'd#��/i���v��;x.bV���SM��	�2>��n��)��56���wLn6v:�b��or"�}p�]v�휯��y�ѽ%��3�;�ƚ��f��x��Seo���m�������떞�����Z��N��Eu_qy�{���thOcX���:����ou�V��{A4��S5�$J0ގu�;�Z�(d��}�2 gw_:.�[�PZy|��]��Ot��G7/�x.��"��
{��T	h�毾G9w�E�W�g�ӳ�1��u�ѮJ�{�mWdW��G{nNG�S�=Ȧ9y�|��̫�kt�M%淐`��y��B�)`у�Q�쪂67u�洡5/��[��<|sa�f�7��6ø��'�(rtPF\��A<q�[<��s\�)tܮ���[����G$��͸�p�f���R�k7�N�WD4�ŭ�Am�FR{7���uZ����P�Ù{;j1|�6�������%&Wfrx��&h�۶Ō�e����Nb�����;�c:��;)��8)ڭ7|�rLnj����du��['tf"�'@_�fa�h;Ff���ώb�c�*����IΝZ�*�*�[�Wi3fu]��	�Kh��S�x��Ʌ�η�s����?\�Ή��<�����ִ�W���b��~'�m��{�����tq��ٺ�2E󨁘���%`����^�q�[
n�e�R��i�V\��Z�9^����1�E��=���mn�c�٬%�[�Z�	�qL_.al(�X���q�?[���ڦ�	_f� %�(5,��V�ؗ	\ap�cb�&��Onvm¾)�yY�z��`��Z��Iɱ��s �ڗ5�҄��W��P�7�	��,9����%�B��o��qF���v��o�`�@w�5����-װ6�c:3HS;S��w�k�P�����?����i���P���%A��VԤ��WE�f�ێ�*&Ȣ�:^Zޤ[���m���[ሥ�(w|�(߂LnЗpb�vr��AH��i�uķƾr��[���mE�1�r�����l�e�8=d�"����k"U^Q�r��}._[����#/�u��oh��]��X�{���}1t��a2���AMv	Xt�� ��t,�睘�nG�\��Zs.��@v�r]1`��Npl�}܋��Na8O[����Q���x�Z��a;+�i��/�P�.��<�uF.��ޤ��	�{Y�
�o@��p�vCn6�m��㧶�S��\��hƗ52�6-��-p�
CW�3r������ٰ�٘E���@�\������B}Fv���J;W�:jau=���bd.�y	��o�
����"�y���nb5�\R!/�O��s��YYK�Kx��n1�YU�Ș�c�Z�}R�4Z����^����>�[o���ܫV����r����Q���j�p��Gs~���ۋG���٤��d������^�����"�x���綦�=��@n㐻��z7����nr��qڢk;�������nՊ�;�V�ӳ�r�u/7=���R����#�j�җS3��Ξ��$1ɲ!Q��Sr�㲧���!>���Y:�/�}cUm:��P��Ҏd pvE�"��cT�Ljv�M���gN�nWG��\���D9`���<yow�]L��{��gR;\���l���{��e����|y����X���*�8őa���r��Ҥ��ue^l�tj����\�
lZ�*﫹\'�j7�+���v��[z�_>����v�ʊ@l�p9_Ӳɭ4r;�y���)rZ��Z�0)fN�r��5��>���ٽ�:c�0TNzܯ3g�Z���;x9�ŎEU�G�%�5�=�p��ю���G�l�B��滜����V3_s�c[V��ܷƾ-�r��>�[c5vL�&��žV���b�9S�Cf˦���fS������O�(�ޞB�yD��~�d�4)!�J2�S�|�h�<�j6�=C�g�}1si����.�Ԙ�a[6�|�د�3(�����Z��]�M��#i�;N��]��#���݇'�j|�.1��0�<����C��<L��zj���RP�T���ٸ�{Z��Ԟ�s��}N�"�9l�f*���e��H�ݽ�ç���o�c�O��uZ���V�r���͕4X��j�V�b�sC��s�3�W��\+����{R�z���`���oq���+ju��ڕN;��T�ُ��1�4[����z}tF%��Y���M�8�ҝ>̇����P�\��Nk�7ܱgX{M�+W�'p���\9-I��z2\[+6S��F{���2mZ]��Kf�<���J_\bq�<˩���{�9����z�Z#��}{w���w�ﮩOc�e������p�
� \N�KA���������v�og�vo��Ȃ�C�Ss�%1�:m�Y�َw���Wv�m�r�9�9ܜ���-��ߨq�|�H�[�<�z2��cz�K�����7����=���2���]��K���l�*�em澓�:��9*
k]+������O�O8��u���;�Tt���%��vt >U;<_U�JTj7���k.���R�:!�\]VwQ�3�������L�p��wu�΋�oM�d���j^�y��i�'qb����Z{G��_

c�}0T���j��;�<��S�#p_vۧ�؋��u�o����Q�B������t]ૠ/]���WV�1|����u�rWEqU���{���BY���^d�%�j�TD�rA��"
� ܣ�;��E�޵�����y�r:���{�T�|�r���2�8oh�7�k.��š�:ip�h���	����]�9�u��eM��m�52���qipu��e��u�r��q�{�m��i�vh� ��N��7n,c����x���2�ⲥ�Y�Ѐ�.�(�nY2���k*� ���c��������n�=M�ڃ.¦u���G�.�&)Go������œ" �[Zv��:��v
\�w�C�����l�*ek�gY��!�,ԟ���2T�eZ$_m���|m.�6\nN.�\��c������C���Ug#�`���:l�t+�(X�Eev$�]E�H�n��o/�D�z�F��{���W[��s�o Fsa�Ң)N�9V[�@]_X��ȰX��i�;���ܭ��B��Rײ�&h	W�+T�{R���+�7A���u��e�]�E�`뮅��֎���WN�����{�8K�9��.oN�[dNξ��F�Ev�颀U6]������s5'ȅ�=v�Z�Zyw��V3�Iu ���k�-�C��i�O1��k �F��Xj�0R��|�b=�V]��D5������)�9fX:��z�dLT#�)��Gz�pZ��Z��1;�C���!1�6�YZ�M������goZJ�S���;�3%ɷ�w*F#cl�ȨQͮ��G;4݁�U�.tٔ�1�]�	��0�$�M��:�ܼ��XJ}3��N!�woA�w�D�5���77�-�?K�@��|������c���Ŵ7R=0���D�p�[���8�)8�ʙ�6�Rz>Z�q^"
�Z2�v��]��PA�b�i��H���n��N�}�K<v��Ϳ��T��f>�]|���G=�:��]	�Z\��
׽��� ��ܰ�;�Ns��8���
��č�"�n��x�3��G&Au��<��c���C��C*���m�`�T���oW?�!A��
&���\յ{��6x�豕*�#�>�y�ћ��$>b��q��x��h+l�B����>A����᮳�;7GM���yuP��ET*ܠ&u1[����oCB�Ϯ���̖�FX���>�rf�;�l�d������m�N ѫ�Y�&�;��-����I��x�d�ZR��Δ��<Kā53F��ӱԗi5j�
ʀ�S8�{;��6;o#��{�WW+t`��,6���µv�=B�Vnд�o����8Yi֊r�ծ��j����C|�+��B2�b�AwCovm�C�V�(0�����бWc���]8`�4J�������[��a��#�sCJ��gw<�,SN�\������g>6bÁ��VD�y���	���7\#,��wV޼��ْ�S�F���Yn���R�SLS%QMD�Q	KT4Q3TDMDLTQT��U�D5MPT��%�1EIT�4�PDf`DSUQSLE%4���PQ$�SAP��0ETD@��4P�T��RP�PETP�4�P�E	QP�DS1�TQUM$T�D�T4ET4QPL�EEE-UPSIT1DD�PETUU%AUADM1E3!CSASITAS�Y8�QID�HC4��RUU!M$L�U@LD��E)%ERRLU451U	QTU4{��_���,��B�Ny�j��}G��[���{}��XӒv�ʹ��%��5�ñ$��tw{�'����ƒj�l��-��
����<��]m��G:�1��I���wa��)�2�]P%,u�g����Z|/�F;h����f��ݻ�[��5�e7��f�=].\���\�*�}Qf�/N�
�rwzj.�l�w-�����rLMCn5��F*��uz�d�Q��U5�?{���]�tH��<?R|�f���X �0#5���[Q2�V����V�#]���{��6��L��>sπ�J_70�M��'q%T��=�\9�q���]��V���%��>���'�F�o/eE�9�wa4گ�k��T��u��9Q����u�f^��}�WC
���)��Y)GL�9�ځ/�_�_>ah7X��]��(��2�)��[}�jI|����W���Vؗ\ap�6+�l\���vl۴-*���^tV�W�辳�������sQJ�����|�7���L/�۷W�`�R�_L��Q�mY���n�7�O]x�ѭ',��x���N��n)t��n�����m��w��j,�B�A��g�nI�x\���)q����r�(
{hV����0k���,��'vi�)IIo`�h�1k2T�=Bj�v��ןFD�X�)�ʣjzjv����N>���mk2�*��=������Έ7�:�0Wϕ�Ԥ��3a���9�O"�B��m�f��-�یp���R�D
1�>�iA[E��ؚ���ZE��kk:�S�P��XX�[�m��r�J	�RGV���˕�^�ߪ��E|5��_wػ��5,��&�l�,�F����kis
�D>)��Ϧ��\�m�Թ�e�v8V��Y�����x���z�yqZx�wΆEG���ۊo'P�Guwٹ �a�ح�·>B�KZ�W�.1�Y	���Y���[�q�<�~����tF�A�<'6��S�C��,p�mƸW:�cP��2��^��v��*� /�j�j��Ϸ��nU��οW/O1{�^t1�pߟyn�*"��1��m��Y���l����#�
q˅�!X�'6m�{�GC���Svֹ-yp���,9J,��ӒY]H��[��S����Ɛ���Q��;5��]�d�8���r+V�7a�[��:t�1�oknay��L�+��鲺wt܁j����Xbڛ�m>�}�\�
��	8ֱ���ɧ��RCFՇ��y�}h�ھ�i�$��wΔV�O1��:�󲧛m틎1bha�co %X�ݛIN���?Z���e|U�|������Q?_.ee�UڕUe��-�ɏk��-��nٛ���g���?5��(1am>�����nK����o�܊m����o{h�3`�傝TSP�F�EE������t����=f4�D�����H�@lּ�e�^N[V�H�O��$����}������^�i8[V�m�KO`uq9����<�msj�-�����C�j���;�o�|[촱���8h����,|�Lt�B�5ض�'R���wI�	-7��:�������u�k�\Te���`2���޿���͇,�!O|���~<�vW<�9���ݳ��+&V7��@����x�����%P<�Bũ�q=�y
���]��N`v��"SfYʐeLR�fne�Κ���*v�k��H��1V�m��&����5���ɦ�^���_s7�t�l�O&\k����F��Q���05
�Պ�u������1����L�,�@)T
�8��o$f����jyN�e�K�IV�v�.sI��q��ȟ��g����o�7g�K���o���s!n˺}�{�j5=w	�4����7�)��DM��_Y�����4�.\f㏃�{/>�z�5g.�W�m��m��lC�x"���g�hf��Dι�U��ip�+����֟����{w�k��g|&3<�1nR'��k��̹��g|�|�Oc���ʭ��4�.ӯ]�%ni�ԣ����X��Ow�t�Ϗ�;:��r�ӷ)�z����;�����=����wY�1��s��yE�����J��~ₗ����m�K�=�'U���K�X[�7�M�sך���V�\M��C���SړT�\�n'e�PU-t��*�4�C��9�ۦ�ԐoeGd���,����Vv����_W
[�r�W1%��kXW[�ؗV�A�i��VD��˲t9�|���@ظN�d�&�����Xqf|�,�X�����	2��}�.q.�Gv���e�=:�Dk�5��|:$6i�Mm�O-�i)��h��Nf������|��/z쪔��.ou�W�Õ���f����H_r[pi*�C��0T�Fwu��[Ӗ��8��S�j�5�uN�]��f�E��Q!o���}���q��E֍�j>ܙ�L�w�D���ې�訋lc(�!O��S���uS�\�QwsYQ*8�uvb9Ջ���A淟�w�D.�or�T���\����j�_c�����_O>�����j�k��pͰ�\.&�͓�(�;Д�[�ˆ�-����k��7�k�L��>�Q�1<�_}[�MtZ���vsީ��U��cb�;��Y�XW.��z���d���d��͉��nn�z��q���|ہ�򪟐�땼��7<���~��e���p�I��A��̤��}r����Oyk�)���X�sG��o��ۨWi�*O/wA�SE�h��[=�PP5 �B����5�ǝ�XtO�L�f�\4��)`��Dx�mQ��K��i���}�w��s�(M��>,G�帳6�Zm�^�����ss�{���A����vEʱ;:�3+n�\q����mh44lx��7A�f���ռ��)b�gyǳƇg��ˡ���[���{�ڔH4y�߼3Ц��wx�%�6[���nr�N�_v8��|���:���{�Y�	�����:w�)W)a'`�_�uN�^��\�`��FC\�����S��M�n�VQ�����\��Nj6�%�w�[j%�Ӹ�V���7
R���3N9���=�[1�d�2�9�w�#j\��r퉅W�:��&�.F�g�Y���Yx��i�ޡC���`=�z>q/tP��71��?(�V,;��>�I��p����RU�O|���R�=ֱK�&�U0�`���]�v�"�^�Z�63j�P�3.k78Gjإ�1Ry���v`�1=5���os�j/��8o0XlŐ}k�E�N�o�ؿ}�e}�j�r	�_m.z��2��B#U�IF��r�k]�T;[7�旉h�v-D�VV^R����Ͷ���m �y�U�)��K���Z�z�X�f�~���x�6���w=���p�d���c_#[u�s��έ�]�^Sa_Ue�R��؝�UAX��m�	\u�XnM=Hc�s�虄���u��o�m���'~�Q�(�@<�n�5Իf���.SCX�o0-���:�����ٳQ�0��\c�q�@���sn�#z������ދ�;��K�Kj5Z���k�9m�>�,��]�?ti�]��ۋg�_7%mL���+)j��YQ��$�yk�5n2y]T. �J^�Ӹf�����m�[�O����Դm�Q�N�������kQ�N`Œ����6o;Y�)��5Q�0'�0S̈�e�ڢk0�c"�FN��u�w���(��	�Hoh}{��s�AUy�lʒer7S!�x�&f�)N����q:���G>ݿ���{g*"�r@��s+yl�?�[�NK�˵�;&2�����Dor[����5��WeRf ��ݨĵx� ��!=�l��mdu~߳�(���j�OWΓ�5�C��Էo1>�Ux�Êd�M7Y���v�^n��MJj�,V��(7|�&�s�t�Ig�ih��I;�Ԩ�8���T�"lz��޹�Tj*Y��|/oL�O��[ѳ�T�]�DN�Ds���-p��=ܗb���4�r�8ӵ��4u�*S��������M�,�[�K5[ӧ��UR�����[�i�fP��2b�ݛ R��WGr�W-�wIp~���RWi�oHiޥ�t��oI�fk6�7Y����v��J�s>zew;6�W9�d�Y��iǹ��]M^�֚8��}����#�~���\�Wꖏ��ɭD��L�u��ة!�\�j�g��I�G����>7>�ՠ{�M��}d�e"4���[f�!��lxnw�Z�`�D+�g�%/��|�G&��W���O���� �@�4�d �O�i3pt��8�=�s7ގ|,ϣ�:lTK�ƆR���9S�s�G��]ɋ���4o����|D�kQ����D�Ŝ�u�����p��pb�v[?P�ϕ�S���W����j�	���G�{gΌ{����DycG=`��4X���Tq�*�\ǡ��lW���w�/�>��c(������#Ӿ�<����3��t<^F��>��[�C�M��L-��P�TT}���a��azg=Y.2�az�bM�]cI��ͩ�ш��}�Ww)�R�Ub�E��'2���[�z�������r��A�:�4[��Ԑ�رi�op�h�si>{;')˹ǜ$'�7i�߁�R��^���|̩i޵v�z��&hg�r.���F�f�o�NS�_������G���靇��9wQ�S�{Ӓr�R�ӷ2��A�Åfb���6�N(��"M�(�*�5qeJe��Nq���,�YƢ0�8*9���4=�;5#k]�'��>[gގ��J�����3�Ɵ_�����O��u;��u��ֆ������"��xf^J���O���z�σ�g��^�q��2��A�����z=^�?S�U���Ͻ�ݵ��js�Y���{�<P���K��2<:�o���2#_Ӌ2�]�yb-�z��,�`z��/c=Z'_D����{���
yu��	�Q�P& �T)��q>"�Z������ꇎb�Ykz��}>�ZW������|s�H·Tÿ��f>� �MI@O�*�>���*r�ޛ��GX�g�y��Q������֑��<W��tu�dmǦ��s �JG֬v���@��%yL��K��o��#���IW�'��Op���{�H���}޸ۏM�����'{H
�pϢ��ny�o��1�ਂ=�E�r�g�c��R7��_�?yQ�~��ڜ��A�ث��U�/�ݍgqSgc�C��f�U=�\�.6l���)6it���R�5�.!�V�|�J���{���jp��\�[/�=j�]a�ɞI��t`:��y�����/tC6��zs�J��7�Ē�:펷�Q̨�{0�sj�d����&�={��	PuӤ?���W�{P����܋�Z~��	U/�<�25�R���p���{!���Bx��n7vo<,���5<� z� �����z����+�}[�6�x�f�Ƃ�<՚�}�{o�n%�nǗ�]�o�U���8�d���mH5
|J�p>#L-�Va=����]9�������Ozx�>��}��o./�^G!��S��eD��.�
&�%�PrP���r M�%KۯWdӄ���R�*:��N�]/��:�ǲ\״�Cs�����O\�j�3��	����T���=�9�=���gGmNQ�q�x���ы�#�>�K��w�Z����;�������&��o�n��c�~ʝ(x�̓1r��W~��t�}���W������e��g��̛�B�������Ӷ�9���0���z��k��7n�n;�BB�+�lc5S�enr7��2��G�Kgs����Ͻv��dM��22"�$�+Ơ�T+���KohTL�I��/��E��Ϣ=�w '^ӑ�/r7��qμ;&낸�U��L��k���p�=�ZI�a���G��]�6ɮ�Oiu�4�5�غ]��:grP�DNuu��l9̈́��B�R�_�z7���:M�zX ˦�X�^=��^v��kPx���R�7�2X���1J��U>(��b�k�Y���B�k��Zz�bƦ#�S�Ӎ)wY�a�}��o
��ʶ�j��uoB=]E3*+p�a&��dm�<gk&����L���m�|
Ċ>�B����Pl
uK�Ļ���3)�|�Z�� ~êud�rvd�'jf\:v�sI��r��ј��&��K(�벡:;{v8�aeW-��i������:�7h�R���Ld谥d��MAh癇>Ptv������J䄩R��_p����<����Stm}�@zz�L`���k���˸��x�LuX8��C���	ǆ-��3�
����;f1`s�В��ަ����i��X�)�#��f��#@��`�7v�f��v� [In��g^�0���*���"�Oo���Z�X[�Z�
]�f��ͮ�K�#Pk����w[.Ju6f��+s/�}�՜l�W�<�%�gZ�t���f��PD����[��Ýj�r�*�/�h���Y��C:����/����,���&E��}��CVn��(L��sCgK"��;��{;�g�r�u��nX�wi����L�1չ����ah�2���]KA��'*���Z�e�,����[K�Å+�P�KD"�V�>��-����IGջd���,s������������mro��y���|�MMtq�4ve�{���O�曰@��0u��R��*�
ÂEN���Yl9+9p�j\�.�:�<���q�X��J��9`�%�7,�g:�rYB�A(lʴ��l�N!�PS��ܨM�	�Ռ��6&�g��9�6�Z�w)J�X�ơB��:��-}��.�N�ลn��b}[4sM2h�F_<�:�aD&��zFɝA驥��nD�Ss�X�ٍ��U#.}��8�p�Z�	��7�B,3�������	l7�3{/�wR�["�~_��I�w}�Ɠ�*��z�If@�\oxU��r��n�y��	��9��U�'zN[�;y�{o[5:��%D���q'`r�)$�Ok�����yt�Զvh���XDZ.V��k�O,y Q��{d����u� ���8��;6�<4*GR�s�QƵ����C)hq�@m�t�Em�z^C��=�j1�?[�ko���tQ��Е��6��E�"w�˼��+�;(�.�a�)]b�ki)K�3w9�/f]$fR�*%)u`Ҍ��iR]��9���O�fV��F���ˢ�\])m�%NWP^�HVed|&f,7;O<�S��4����o,��8����r��7JP�v˵b�����J]�p��֒�ӱTS��X*�X���Ҹ�XM�LR�ҥ���lHu�Y[ݑ������}�}�;���&"���hh((
��������h�d����&(����"�
�"���������j"�*�)��� "��`�����������*�����(��3D�ID�aA�DDERD�Q,QL�RT�U1!UQ�R�EL�T��QUT�UAUSU52L�EID��UD�PQST1ET�QEEULUAQQTD�D�UD�USSIAL�DA�DM3T��D�QAD�TULAD�TTSR��U-AE�UQAD��ATALLTL�PDL�3S5TEE@DEC$�EUPD�55Q޼���x�o�c��9oJ<JW�����ڐ�Zfg�t)ܾn�"s���w6&�8M�۬U�AI�ʙleCɤk7�o�T����6�J�˩�z��sw�>d��.#}!��*��6˰lf��nR��8���vwk����6�:@�l��B�g)����zЋ�=��>�8v�ꃙq�t�İ\�M��m�A�cї%��H�-��g���|����C��:a�o[2�����>�qũ��>��_}(�W�О8s�Z.�L�	���u��h���t��������/VO�Q}>c�*�K���_� ��J�2�z���nLL��7�h�Glj&����^���B��|**��E�>�Ƽ �dZC� �t�tW��K8�W9Z�*6�K���/XRZ9G��>���������=�F����Ȁ��\q�L��L3=}���OFng��Ç}#���Խ:/mu�f��7����C~�F1���F��k�N��� \��x����4}3��a��8���E·\OoKv�ǅ�u����C�/Ӌλn�����}K�zD�z�Dƻ��zY;��N�N銛�i�4����`�W��ޛ�|��߇^W���Nm�ﻫ�����TK�^�N;�eFM�����z`ƭQ��U�v�N����m����@7�(V�c7�<�RT<��2�*�z��MX���"@��x������">��b�%��~;H\Uϥ��m[����4u	칑�[*6�-q����YY�c���ƅ_T;Bӂ�P먄}��}d���yX���@�Us긙�O�P볽 ��r��9����yWǕ³�$��r��]�3�
�-M����z��E<X��yQtv��L¬.�7�S/��q��^W~��ܝnI<罵�ο櫔��������g�	T6��W�<����V'V}���~�>/?O�W��{W�o�˨�g��ˣ����K2�����I�`H>E���~
nhN�����;��b���f�n�q0M���y
��'�3~0�\�P�L�$�2,���>}u������������{�
��o�83Շ��+=0,�ΕB�%�"�|g�n���x�PF���J�c��Pho�o����u[��x��?RM�Do�`�*k�)�� �O�=o]�u'���s����r7��
���m��>�����x��_~���̓���������b�"|G�}�­�$xd%>��#Q�	��~�"|s�>�����䐟�^�?��P��st�w�n�q}�h�9f��ǆ���^�7K0ډ��ˊ��*�wm�N&���Е���M��,Ü��X�^��=����3:�^o�k�[���u2�"�b���KU�Ǐ ySo��Dm�!cz�ko�^��M��Kz��ٜ��v/��'�.}���	�/NF.W:gO�?}C2��������k��:�0���LZ���7����W�`"eglk�����{�k`�}��p8|��MN�%3�B�>U`��^�ަ9��r~���vR���C�Y�si�,��UO�� yz�P��mH�>%T�}bwL+��[��W:=ٽlxo�p	a�Ǧvj�����73�q9�o���~ɡK�R2�Y;@��9�r}ǏP:�@�mNڽY�W��{,�}҅E��c��o�v����n��߻Ӓr�KN��2��@��<����S=-��~����Z��鿱.�}��g�8��;KŽҷi-����o���!F�ԫ+<�:^8_�e���uԬ�O�y�����7	������ǲ���z��3�B���.���3z�o*�i�}�*tݐQ�P3ŋ�����t}���xoG��]�oFz�2�˽���>�+��n|<X�.������_3}��"��O�>Y���o,D�FZ^.��||q�9x��[U��[8�H{�~�=�>��T*O��<(ʢ�e"���ާ��0͖�g���S�S�8�K�R�Xu�Զ�Di\�EӖ{O�X�<i�A.V�6��Eb���?*��
��'y�u:�(�U�z�����c�:/����]��1*� �z#�͝y�n���%����zc��:�,���LޞVTuj��կD�ͨ�D���8�>g��CҾ�*#m�0�Q7��=�������Q��H���>ed>��o_�����ZG>.s�q~85Dg�dmǦ��H,��\��ԉ������\�c�Ϡܐq΃�g̱���:���~��a���t�wI~�F4{��E��;Z}�yِ�/gƦ�Q'�dO)��e�\o����W��T|O�|=�bzk�����X��Nxz�`W���'��3�wT��Q�=�v#��w��#�zB���y��n�*­��s7^��w������q�S�܃_)d�@0��T�ľ�ӛr�z����v#'��U`��nR��H������U�{���SO���w�dS�UD��� S�����u;�	i�/U�z�Ȥw��7�yp�]������{��y�.��#�ˈ��(����[^�J;;����g�9C�YHmº|O��\gZ��D��i���]��<��U���vZ�?~]S�Ը#/c��z��3㳤���l�w9GE��^'r!u0+s�#�%��x�ֲ��T�*�R�h�TNA"���q�cJ�ٸ�x�p(o*��Q�e��]b&�����F�h�g&�v�K�Г�jY��.���em���B����A��e �7ۯ#B�'�Jy��$�St�ܻ <`�p�74��wH\,��=�Bp��wr0���ᝡ�[���kr��V�$��"�Ы|b�T�E��;��XQKj��A�@y�i�O}k�G��X����@�C�u�N��R�"�Jfu>4*ʇ�R����Q�.�d�3�� �z��TI�zD��}2�x��)�ҽ���<�]���7\*eHۗ�0�'7��]�+w��+�טN|عa����<n5z��{N���7��}N|5}7\�d�R�'�Á��*��//ʆ�9���)Tu�]SS�.����z�M�w�9��R|_�Hg�<�d�^�3'��g��p)Vz���x� ;A�<=)����c>}u�9�{Ԅ�z�hh�O�m��N�����V/���٦�=��7��G���!{Pͻ@Μ��Q���t9Ю5���z�����͹"���3#.;��3g������~�<o�W�&���B 7_	�b~���7r��hu�i�/0{p����ݼ�].�c�����>�"}�3���C����_�&���eX2#�/��Gs;�[�kݽ���u������7��G[j�F���HxO��hꜙ�R��Pf_�넷g�EE_�ö���f9���|��K�>SP�a���e-�hyMdK��Yk�t�'bs�9��H��!yg��_��m5�E�q�<��珻����ە:�$]Y��H�R�2k�仔�����A�n\�ƍr�3�'KG�4^����l��t����=}q����O������~wrn��4n=�P�n���L����U=�Ӕ�s��cO��>����9��Zt^ߺ�+#z��w���0��>����{~���1퉡�_�|��]�����B,�_�j�ևu>Ӣպ�{7��\v������ m����^�I�n�{9+k�-_��v(�ߪ�n
�C�������	����Dʍ�ҷ�����O{AR��?Wx�9��{���Y��'3L��Gʡ�eV����{��.�ڼ�uMj����d�W 1yz�/�ܯzNG��_N/:Agв�W�Ӓv�'�	vL�=��b[[ռ=�����z7�m��7�P<�GL�=�М�v�_�=��������9'C�$�=N�Ʃ�B�ܫU���D��|&XW�Nf."��.o_�����+�G���~�x��[��
���Yw�{f����O8���<nԐz��'�|�]J��eK7�7V&�9��8gz=Lm_=�P*n�ƻ2�c�(3&���}��a��䢇�(��@�۔��'�^�p�EV��z���*n������U;��{\����Xe��A�-W�>���s_.��`�v�.ח��s	v Tjr��W\�/.���n�:���)�n��UY��_R֭�Z�W�q�.qUκ)ico:B	�7Ln�m�0Jˉ�3P�NV�m�v"��cѯk̮�<�ԁ�n�C���f�D@���n��=+��si�8��3=~랗w~����r���ז!��uC�!��g�Do�X�Ir� 74}$(������VFx>�Xih>�3̭bcQ{�c[~����>�zv�~�����f�s$�v���/�^����z'�ˏ�*H��n���u�xr���5i�����'��߉��@��2&�Y{��7�qM����d{�Y�31�_�V
�s�4.#-��Yʟ����w&/��>q�eY��5���g_.�sw�z�k��2M|�'�>�>�-m��s�4���j����xa����{����}�P�Mǽ> ��ࡽ��|J�0��>�¡\�>V�`�r+���������(5WZ=��U�u�G��������\ȼ,�P�7fŌ����e���#}^�N��A��'N}�+��_�C��o�w���9���N�����|X8s)�s�mFW���%ޮ�����eV��S�%ٟ@�^Wɕ�ɸw>g���Jo���Ur�?�/�� �����<��cd�h�ST�m������ԃJ���sY���^\;���֧:v̚
4�P�[R����쩏��)h�rEu$yjW	pU�5��������dmM4�ݔs����	`2�rY1T0֭(ڕ���"Ve֥]�7hwq���X?v#�'�xe	�z]\�)lπw���m:~>+���gqr�ݟ
�e�uπ��c�y�w��P�?�	`�>�����2�z�<��#�`F�*Þ�z+o���H�P�|�^�Y�C݆o�T.ʔn���?�2����S�ȅ�Q/�Gw����R��8Gc�jqnq�^�{���A�8��G�߭�qɹࢉG!ITf	>UY��h{=��7y���w��?]ģS�\Mϝ�J�s��u�甑�e���T��4�� ���ѵ�+�7���,�8�|�hg^�\�֑��<W�~���=�#o�L�\+!����Mi��;ž ��l�OI>�p6:_����7� �z�1�����>�~��`�����{g?VM���<���O�3Wh�9�<���E�X��m����l�w�4a(v��i�wc&�Y�6���V���=-~@��L�B;�n�[4��=C3(������X��)_�`�w�܋~u�}�=>}����b5�2݄��~Ȼ4����X�J��mf��빘��;m���]�F�����P?l�D]�J
W�5&��xk��n��]��&���>�{��B���͍� 4�)��c��_+�:��WE�	gf�1�r��2>G��o����p ��-Y�w����T{���nV�k�#������C��t�B����߆{ή����z�`�8&���u��=BǴ���z��^+��?�uO�q��{�G�����4���/� z����Q=?nX�}�9u�w�G�&c��q
*����r��ǥ�cgG�+)�����x���:�ǋ3�1�߫�^Ǖ�J���b$͓}k}=2�~�?�G�����g��|6t;��:,ү��|���W�t��L�ZJ�L��ۆ����V��$����%�+�"�U��ٰ��ݸ3*�.)m_�N��ϴ׀6�G �L��s9��B�Us��#������?���'�geN�����^!�^?C����ޟ��4�l��>������>��d=/ޝ��{�hxv}7\+��R6��xԕ��}���v�=����p���S���wp�z��7�<^�o���ׇd�pW�6J���0o�V<�������V��&��<;��3�>
>yu>7^�X�n��G���|C:����tߤ��ɡ3�-1Wܹ�9�����3�$)^3����|r��Bn=^�4b}�h�f�{hz�[ꬩ/�p�3��c}������ӌ �*<�L�0����7V�m�퉻n�9j�V�������y��R��;����(���I_#����,�v�����W7Ǎ����,6���DW"h����l
]���t7���o���ײh�h�u��{�������( %P}DLIo�����9�t+�~�8yC삣ޝs^�Uv������W_���o���&�3޸<o�ꉨ�d�H��@�&&%z����-v��Þ>Y��
]�����0z�2�H�x'����_޿\K'�+`�=$v�k�����=_����Q�Į��1Q�ڿQ�{ԁ����AցN�ɚ�,�{�^��c����kM������Q-V����3�q)|o������M��^&��ޠ;��Q�t�(�#ۂ}y��gW���O�s=4rX�pz�V�����ާǝ]C��v�c�Ez��0�VS�5��%�G*���~^��"���>%T�h�o]��~a���D����%_낏㺝@���t�ub��q�^��F�O���M����C�6p]��~Eغ�T}����b��h��vX5����H�h���=���ȟW�Y����άw��ʑ��s7�0��)�o����&�{6���V8��ύNi.6X�^��W�'=u�s��H,Y\+���;w,������<�<��)ҏjU�ݪ�C�*��{+^ʹz��%�Y��*2�7B�'�����]s��ot`7g��1{I�J�i�Tˠ���y���c�7Div�J/�������6MY��\��;n ��H���&��.�xU,	;�.�5��P{y��TiٴuS��S��H�\�J��E-�w�l:�`�!c1ޝb�����hf�D:y&�v��|����o�ކڣ|ӡh�o*R��ʡ�{�:Lmk�Ջ�b"k���y�5��X�{&��<٤�U�R�Mi�����q�����]�7�bU&%�Du�7z3��>�fJt��lt���=��V�7�+s!���zw_^����EB�/-��?*�{���_<H�bkUuy٫�)@|9���c��V=��,o���G*d&եc� 
�F�s�LgDv��Jʑ��աe*W���lAn�����F�7,�2��q�חz��:�,w 9HԻ){ԛ<�Vv�UO�%�{-��wU�v��0Hҵ����Z�s�BY{�6r�M%͋�:o+��m��oP���T��d��7�7�p30_N�VE�t����� ��;��N���W<���h��7X�1V�!k ̭۬V��r��j������3�>�.����ڋ�di���e�øق�*���B�]�`{\8cx/H�n�q6_XW�Cv7�Fƍ2��,���|�F,Nk������ʅ>�,m�/]�x{��\�*eP����85�^fetN豬�T%]:����Wfh��et��7.�C���ZiN˵��)&���љ�6�0�Wf�l���$GT<�ſ*K�ʏn�o�̗�w�;��B5(���;����"�U�^��uB
�,�Ǣ��v��rJ*���Wc�E.�;��m�,JT;o�ŷ�ģ��a
-,@�m���÷�)����:�^!�����q�F�Q�Kn�^�⭮��ɂv3�r+z�[�c�,%q��K�o�X`K���������4��W��6�dRS�^mCZ�Д���;(�K��&�M��kj�fL�B���dnuu.���cr�X�����9ֻҎs1p��9�qq����q�/���|/�/x���]Ų�;��3�N�3tv��w�� ��w'5�Lq]`#k����}�e���*�tR(���s F9�m��������N��}K��١�4�wm�`�D�	u|����^���Z�7o��˼�|�Ç��q���3F����X��[�S�ҫ&���&�:��	J�{X�a&�$����7���qF���GX�a��]��m�E�5�P�����a�j��뭮�ҶD��T��q-��Akԓ8�>� ��\�u��9���}��c����ޛ��Ԯm�8�򣯛�cX͘����	h�U�_wq\����q����M��,�s�x�p�f������m�;�Q�t��u�"MƵ�~w��{�~��i��h�("*�&��Z(����&d*�*(���i��h��&�b�
�������"$&����*�����bf&i������*""j�
&�)�&)i��A5MTEE��TTUMQUTđ�a�0DKI0S�PSED�$DDDPUDTPE2�SCRSLITQ5�M%ESIA4I�PUL�4�R�MQTT�E%DUQAEAQPQ4�MRSDEUUPD�UUEPDU4ĥ�TD1EHMLIIe�RQ��W�|@PL'��=|Q΃l������ֹ�N#�]pZ�	���Á 8�����x��b��jJs�+;]�O���M96�%�s�?�G�U��]Ѹ�@l�>i�x�������q��Ey\od{m�^��zka{s
�מH��SQ'�/�΂Z=)�����0\�k�Xy�W��m�"��)t_�4��q�Y�2=r{�=J$˄�oO�(��H<��,]u+�w2�}�X�����*b���}=��u0�x#�������;�v�w�(��J����pz[s���}G/�I��Z���Q�.�����H/z�y{k̭򣧮3ԁd���t��8�hɾ�C�gGt`]�A�{����}���q��z�Q�w��\z����y�~�8��z����LM9��s.;,��B%�<��v��)�蕕��Z>�&7�|�G7�l���>�߽;Z����.=7�=��:���5p��q�27+�g*��ޟ��"FJ�!J���y~7�F��U�*!�|���L��>T7�j��Ǻ7%�^�=鮙�^>= ��ς��h^[�Ʋ9S�q��#��mc���NL��țK'V�
/��w>&ϩ�a����MN���ϥ��N}�����R܊B��{�����],�>�z���GFfpޚ����uw8��I�`Tn����I�m2������\�����NA�t��_2��j��{s%����Z*������&�ѷ�m�ɤ���;��ho[c�$�\yEW�*)�l#r��!j�W<��ڧ�S�=�����=SG�> ��/f��ڐk�Ī0��>���pc��z��N����Å�^_�s>Ҿ�~��/=ׂx�{&�G{*F^�'j �m#k�yT� �y�z"�w5>�t�к_��u���uU��οT/9�΍��Qޜ����\�+��oSk�Jw�`�^�gp�s��+*��A���ߓB���}I�;�௥댥�w	yɽ�fn����n�;���aܙ�|��ۉ�2��u��<0ӡ�9�>�}���n���M,{�zЍ���i1QW��sHn��^��U��geN���|�b�,w��^���2��Xd���V�^���}W^�G�Ln{��Vz�,�3|T{r���I�d��~j�����M��\:�|w=S�`y��7����'�Ѿ��q��#�p�l{�M�p.J5�,���3���m��k}t�C�#��9=ǽ��'���뉸�;���<�_��|n3ʈ�2���Z<EfI��o�=w��9���Wxy>�6��\�:S/U�F_�D��z�8\��?H���Qڽ7:�~v�l����a0J	�h/dq�"�֧>�n�{Ӷ��W�Ϧ�l�k]mw�
�ďx/�b�hF9�}2�$�^E�qbiG7�����=em�n9}fan�m}T�嫺v�!;�\�wD�:�qgZXx��Y�q�ʲ��Et����,˜�Cd�tgV_s|f����<UD����끎/ŌQΣq�R	ϩ�ٴ�ݟn���S{�ڮ�ߪ��F{�o�^2*�jl��q�FI^SB�:^=�χ���N�٦_��p;�+%�6�V��:��s�9�^@�F��N�iK'�L���/��o�k��_��Z[���7�����lof{����!~�&�����o���*!��AE���ģ����]�!��'���(r�V6���s�z�z��n�߆G����=�����i���w�d�>%t�q�뇇T�����Y�GO�N�AS��N�M����w��7�yp���8����{��z��r��nj������ѵkF���>ڙ�9@�:=�Y^j��<r7���u��g�潦��T(��[5��-��eĿ�l�~3g�?���L�~��·u9G@�?�ͅ����,�+s �l�4��]!n��p?t���%�)d^
}P�Jӂ�P몠O�b�m_.@��~�T��^�ctK��H~�����o��s�S�Y���|h��{&N�G]C뵷�S�Auk�׽X뻻�7��-	���D�j>�;5=���}ʣ�����Hk�P��j닣����\���������tЧ}ݭYw��/t�Y9U�0�rԖ��W���p{K���r���cD�ޥ~�<����;-V�ݧG�F���p�H�Ab��n/ʏ����8��C���Y��~���+��>��Zѕ�m�x������.���dS��r�>���>,���n^2	Q����eu�{NF�G���C�K���ò&�߼-����=��6�ϗx��r�%��,	U㮩��חS�q^�X�n��}�'��Ϸ����>�e���Gp?t}	�ߊ���YP ��2�����1Ų��������Rq����yg���׍�N��o��d*������d���E��#������*>�'�-��pzW��3�d��>O�g����޾w���0{���Φ5G�]��{�����D�3%� o`O�]F�p�uV-/�9�{����q���9\{���;c=>�O�����.=~��s>�W�!�Ύ���9׷���%��m*7
�#Չ\{���b����������� ;�� s.L��t�����p��-�/"tz�i�Ӏ�N�،�~=G�zW?uǳ��w&���4o�{�z.�邛�w�^J��2s!sy�*L��{&MB��S_�:ǧ���F����z\s��x��ъ�ce����١1�&��3ôue�\C�)M.�.�j�\�ŵڍ �.�'�`\q1_ڶS�S.^����@�w��)�Zq����{��0�\	���� ��.��ۡa+k�Wie=܀^�9	(,�Xw�j���d�����)�5-n:�,�B�,��a^7ӨrI+�N�z�V�+�����\/^پ>�8o��T2a�����������ǽ|�׽���p^�e��
Ɛ�1���%����;��<�ĭ�1{*h��໔�[�.��a�����o����z���Uz�^�� *���3�U��ga������;'�z�E�N홇��r�R�A̿Nz�RC�{Ѿ�u\nO�+׀��H�r��9��Ӑ��\�^��Ρ���ׁ׻��\���'C���Pg�}j��uϠy�'������e���y�q��m0X��&okd_z�W��s�t\Z�O���L�s�>����B\޿U��GW��m��2��������O9��P|��V�a��H�F�H=�`H>E���s㐳*Y���Ę�\S9^�{�����)ر���|�I}�q���t�����SK�B��5����~HO��{�S���Z�$�V�M�]Zq9��������^elyQ�'ʾ�b�]�4��{FM��sK��N���Lχ�v(賰�	#�H���1�}��+����!���#���IQ����&��r�`��t({���`*K.t�|������+R��|�Bp��,kiz#n����/���to��>6�u.nL�I�`�yK2�빗@�;����?�����Kb�|�>��![c��f�/5����N�v050�RNH*}���t����/�����R��`��A�"g]p7gȽߙ��n!Q��~��DN����N�޽��>u��7��)r����>vg��W�S�=$L�Rj�õ~7�F��������'�x8�ݍ��y���,O����h2�ddB,�a{>��D��n��/J��������]��˸£���<�0/���I���M�.u8}���Bju�>g��	�nm�\�}�Mɇ���W�'��yx$��B��xϽ�]�{��^�����,\w��������;�z���3.G@��O~�?ק�����)o+��W_�7U�:�#�S�KL���7�HK�^''��M~�Xn�ݯ\��Av*�Ja���h�ƥ�:s���o:��dC��o�wި^s�S�u��qr�p�N�r3G�Ƿʫ�&�X:v�ea���M��J7�.F/;�d�~>'=s��VxEB����72�W��^�^U�5��֖	ߑÒ��A-������-'�5}~}�r����e�tЍ�f��*�=-Tf���Q����vY>WX�x�=3�;�[�˵G�2��AT``���=~*&��uuᗮ�-���[C.s]״��0S㏖�wgS�A�����������NTU��n��(��򼾝�>4N�����ʕ���o�w"y
=p�'��pbe�3x��@��X� ��[Eb�����v�"NvoT��>������O�/z���]!�f��.ʔo�,��f�*X��F���z��x��
'����ٕ�K�b#�^���O��t��|�l{�D��QD���J���r��i�k�٭��p\����ڨ��h��TO����^�н#�{>�u��ўTF�Ω�}��f`�imy]�;Ğ�Ht�I@O����:[/>}V5�~W}�H�oǴ��i�'�&�ｱ�U[˫Y	�F|�Af�PB*��DLKu������3���� �z�1�3�}NVƫ�����1�^3��t����o�^2*�jl��q�FI^SB�:^<�������ѝ%�oc��nE����>�㞙���6}�DҖOT	�^�=�+���4���>�)����Y����d�;&��0�Τx'�w"�M׉�|=>}��`��܂�'������U>�U��sd�_[H\���zyWiȭ�#ןo\{��^�������{޿��Ջ�eH/(_�D�~Cf�\^�崹{	p8g|vp;�V齹�#����ˇ�߮�ϟz��9�vTO'����K��X�.rs�R@tļ������F�h��࠺9�@� ��=kq�������}n�q|� [/^Ny�%���V�rwv��WU�\����vl(.�C��C}بhօkx���C�:"�ͫH�;IBevX�2��Y�0K���n���߇嘸z�2|��r|3U��x���εq�5�0����XW��M�T�f�wq*�Vi�g�3��G�gn"g��|6t;����J�����`EwI����ݕ*q���]3���^�x�]k+=�ݝ[�3�3�aN��a�"��-�����U����=�^�������B�Z�-�����R����xTgeN��.��<=}�>����幺���l�/�3��5�P|=T!��>��=��Oo��<�T�����P�*F�w�x��d^����_b�p|���[>�x�&1��'��2��>�i��H�{���9��ׇp���]r��鼌�s�.Um�6N�C�	<K<�u�7>��|n��7���}�'����k����8{gy�	5��w��_@6
4���^3å��C��zP�����zc�K����S��an�\|��,�^���\��8]>is�Z�m�>��o���Ҽ�u8�L���Wb<����YJ]���zu��ϝ0Ϸ��߽��&�=����z�X%�D�O��\ǻbּ�����4��,� V9����u�gAU�a`u�I�v�ml�y�]J��B���<��Sb+������%��k�I�������P�u��n�=��@��fԣ����U0�B�g�VpN�l�23Eqƞ.wܡ�D��b��nJJ�G��=�%1Cû?���r~6>���XF��o������>���n�\��q5g�+}��z��W�|�z�O{qH�Kt�����f����?1Q�ڿQ���Hg�x����ؕ
�Rz�VԦ��&|����*pT���+�h�r�ǟ��Ϧ|}ex�9�)��.��ʭ����	G��{��ɨS�����X��wR���}~����{���~�/��98@nd?�sy��7�9��w���<=�l���F·�>Ӣպ�y��u{�]LuTyB�'nwgϋW��^���p����##_�w��yU�W��
�3gC�az��qx�9	v��G/b>5���F�����_:�^�:�K��X�9�<3�2/!K'u�&���T�`ٿ^�� �x����eV�'�J�L��\��{�s�Q��� ������<6U�3)�L�&���ۿ��T@`�xC���N���E�<00�9d�G���~ޯX���ϳ	�J.����N�1�#�|+:rN����z�Pu���1u���_�����9���:�T�s�G&�r���`�����9�v�P ,��#zG78��{O����wV06���篔��Kq�]��K�WT}�׷� \�bV��*v1�+�l�W(�b��q#G�)��NT��Z]��p̩9�M�]�T@��κ�}�ˤ�-9�����x��xѫ>�����:�j�7Ƒ�2�Ź �,�"������R�R��"b�T��1�K�>�=�8gz=Lo�K:��ǻߌ;%�P,�/L��x+����g�{�.�k'��Q*����"�|�z2����*:{=(<��;%��D!� �yw��7:,ߒ���F���:�E��E)��!�zr��o�ԇy�Q�%G�}����zqj.�8�s���q %!/�~���G��Ƣ�|�G[~��N�����փ��k�^�p�F�wϲ��~��zf��)���f�=$�P�WM�#/����rj�G��o�Ͳ��9{p�C'�Nϡ�����)�9��,�a{>
�TD��H�z��c�7Cw7�X���9G|���/�������h���7���3���(2v,��}�*Z�К�i{*�edR������y�C������\=�T߽> ��f�w����*�d��[���g6��/|Uz���*�=G�}˕�p�μ�n��u�G������B��R3b!yJ����+��'�U��#���Ř?|�d�O{��2�Ǧw:u���S��|�S�i",�z*	������_�F.�ڲK&c�4\�L��:�;f�Բpz��D\�u�yM��j�e�[��E���D2�c{&{4�s��ƶ�A���t ɩmn��=3Y2�����a��e'�[���w,��˾�ѐv�y���u�9��kĮ��| �M����v/7������¦;_���N)��q�=�b�r�gc������!�H]Љҫ{�N�=Ҿ�{wH�s��Ո ]�]S�wC���NuI�����q��V�	�o��A��Z�+4���g�U�j��9&���n���ٺ?��e-[���/]u���b߄��5ph��*@n�x��[ԍX��/�l��L��/e7�w8�htr�ri;�|�%Gd��J����y�5u0V��w�b!b�fຐ]]�w1��tF�X�8�4,�ݬ�2::�q,��)��o����!�ѫ�yI�9co�#�Z+M���M3�
u`C��Sᒴp*��+�r���I�ں�B歜�
B�犷�G�a緵����l�n��u�]y����.�p��e0�g
P����t����9$_���,�[K�U���0�,�I�|�9�K��73϶+�ʥqw���&�,c����AYոU���u�4q��'i;�Ӌu>�gm�tF�)7�%�Te��\�Om�j�\�p�9us+s1k8Q�E��=��w��753�-6/�{�:�S��O�]�w�4��M6�֍��Ŝ������okk�t\�5�v�`�i�#���j���]�\=פ<#���&{B��v�܉��yy�������:���a7�YW�	5�y\���X"̺
��:�K�Q/��鮎�h��E�i}�S�37�ࢻי�-5ى�vO!��kVr�
"�uE��<�s�[
n]C݃��ku�.�ٴ:�t�3��ih�]���m6Lz�9�� �_s�e�\�%�R�ֹ��emuB����MT�iHF�gu�Ԏ�Da�\-��
�pk�]�|�!L�co��N��s���ը�v���@�W�n��m�y_vwa\�Q9W;�fsU�G��8�x��q %�,��Zq>�Y�:��
����^v^�t�.�4X�b���qQ4�vo*t\.+8�������܃4wR�Wr_�=m�z�,B�7P�Ԕ�I��VQ�<�eh-_�f���V�vk^qZM���N�[r�鷔��2B���5��GP}I�.���W������KaCw�l�c�V[��j�f���bɥ�nS��
�G{�o>�,��=v*�0;�Ht�����u�k�����N�ܱ��U�Q�Q-��I٩Yt�L,��cW�9W?�ݘ�"��*����3GB�0���o+�E]$^_%��i�[�����E:���v�=�G�������kw8��k G�d�}K�e���͡��(�b"��*�*��h �"J��J���)����*��(*�����(���*�j*�Z�������� � ���A������̡�"j"B�h&
bi(&Z��J`���������rp���)��*����� h(ZB&���Z�j���d��!����(hJJ���$��(h����
�����j���!ij��)����P�b��Z���j"��b�����!'��NEIEJ����y�w|k�?k5���|����r��	���)�w��E�y�Lޛ7���;��@s��֓Rö�zEh�|���:GukmXQ�'w�SSf��p��EF�>!��ʽ~��Yj�2%�{\����9wQ<.��eW=�����T�z��g$��<p7YU�I^%��p+�^WȗO�����j3޴z'3=�27Д_����\$����}�:�Û2�T	�
���Yᆝ9͙�q辤cA��f�'��ϰ}�^��9^�x�SW��Q����qe��fX������^�ޟ\.5�����Z�,Y�@�U����G��r=�~+>��Y��1U�mq��:ʯ~:�$뷠H�w��Y1�U6���^�	ɞ��<ʉ��t!�#�^��D���I_�����D�vǎ+�o��n��w���3`�T+��x�}w�q^�\M�>w�+�yοu��FyQ�`FU	-�tv�_r�ld
'=� 55'�L�������cQȊ~Wq>��C7�ϛ>��J���Ɨ�ŭ!Q^k��Y~��s ��V����n��t�7Y�F��A�eC�c}~����-Z֋�c1肷֙9��?z�����ED9��٩����A�hJr�w+���1����&��o\n]��/�5S��<�>�,,|Vֵ.i��W����s��^���$8d2��Cx�T��nX�Gx[���J���:�d��׬f��m�8B�n���8AM��!�6D�##��O2��9�P�۽�;9Nncb��\��y_��T|r����uy��i���<-~�3�ߑ�/�Z��wY�p���__[P�����.�JX��vG��ɺ�>�����0
����{��s�=T��2�=M=,6}Bt��TT�V�)��ڇ��^���y��{�Խ��}��X��|c�ә��t��(Զ������i��+պon_#��_��x߮�}�ԦK[����o��պWV�d�%�ˡ�+&r�|
4rXV6t;������ T�{�*5����B���G���؎.:��|�Y^���%_��f��38o�|vt��6t;��:,ү�����W�S7<g�Y�H��rx�������޺�V{�̤�/
��{'�N�C��g�Nf���,�4�
���/�b�dNH��4�����#"���T�QN��/�;*t�d�]�ˊY�[�7ޗ�uY�NT��_]Ѹ�� �Uj4��E��_�=����Ͻv���CN�2�Ȯ�����w�%�}#=sĖj$���*��\ר����f���x;��9����>�\?)]^�E+|
�1K�X��n�����F�'6#��t�KE�U΃�E�*�6�g����:	�=��MÛ�۫�����wwÍmN��p���ա�{tͧ��j��Օ��b[q:�{,���Ew�l̽�Z;99Y�_\c3�e(����M֎�l�JX$�D�<�G]Ss�.���ޫ|����yLkQ=�{b��z(xɮ>��=y�p� Ͳ��lk�*2��W��@�l��>��>��'�dܑ%���Y�^b|�m�޶�ǔ�=y�\��S0��f�P@HzH��-��9�?gBۏR�4����
��K��ӡ^�և�W���o[��wF{�����D�2Y@�+�nQ�2#�n:�|+��I1�Y[F��Gݡ�s���ߝ0���D����=�����_�'q�+�A��^J���Vә�!������r��ϒ�~7LTu���}�J�Ƽ �Wp������sc9�/ ���Lץ�¢�fʜ/�EeJ��=�_���D?;�4��6���/l-��b�h�9��σ۱|}�&��*jKcӁ�Zpo�o�²#z��xA���|����p�k������1���^�y��=~����3����_�j�mhw>ӣ;�I���g��N_���|�^���s�Z�C�/~��6�P�^ʚ&����~���1?G�l�{:��L��gaԯ���[�'DyI����C3�M}�i:���I��!y����i`���h�C����3ʶ���*�����yP[�<Z����=y�TA�t֥Т���{F�ev��/���U�{�]k���2: ��S���(��#�7:�?o
�ս�Ck��ڭ�/|��:�^�;Լ_���=�<+=�#�	�)5[.7���\y��f7|[�W�Zo�R�J�,���H�w/ޓ���ӋΐJ����ݼ� �g-�{γ�=�9'n.|Jq2�ў�]^���r�y���|����m�~>�	o�\;�Y���j�N��?TA��ql��b���$�ĸ~a-����T�g�^R������ǔz�wf��e�׬o���;���}=+�<��(}&y�2�g��X���s�8/���?w�9˅��կMWmX��N�8dw����{��������t���!i�~fz�9�.�`��6Q�kǔ���IND>���׽�$\���b�י^Rp��x.:�K5���C��NfUp����� Vx�X�:뉸�ҙ{��j7��(���^��#��Hq7���7���h�3õt^���O�d�i�����Dķ\�h�u��E���#���>�0��ӳB��lޮ}�\�U˰m��=��2KF�Kf�I�P��t��ڌ���5�O��xFo���'�-�S�+�λ�5٤B���Pё�x�S̽��'Z��C0f�v;�(�J��A�z�?��OUͯ(�Y��V�u�Nz�^cy�ܞ���9Yb���9�{��3yBn^֎)%N2�dc傗m7��ܡ}�;���
.��6��k�fNG3Q�s������J>�L��9�5�9��= �^�
�{Ɔ���q�I���w��D��ù����Ϛꐮ�����4}����u��d�;�&X�a���� Z��moy�$�(��9Zk���\5w����w!�z��,�^�/�� �t����(���*>����[�a<��L���R�[�Q|}��W���:��1��q���2��u��>�#y�j�k��5p�ysܪg�+�x���p6F�Ǻ������;��~7֯�"%�{\Ͻ1�S����s1��Uv|r��t�����w�$���t���?���t�*#	D>�U��h�o�+�韄U���S9r6κ��ò;���^��ߺV�-����w���9e�4�຺�g�A�C�S�c����Wn���\��s� /G���/R��9^�x�E5q������qe��fX�x���_{��G����ҳ�����di�@�U���!|�z�7>�z���]!�o�T.ʔn,�����/��}�T]�r,�|�iQ�]>��eD�[������>gs�D>����M��wh1@��k������˙�^�	��z��q��e����[/_d��\�7��l-k�o���G�U ���X`<%d#��,J�f��w�*Ίu̦�Cy�"�.n���<Ꮰ=�e�mҖ�z���=sOgu��\rhS`+#��;v���ʶOw��7k`��S9���J2;���&S�O��뉹�iϗ�y�g��|zE�ڗKlQ
�o��z����T°l�J@S_I`Cs�c�e��U�G)�\I��"�]��'
}Ӎ���7�Gx�ޑ��#=�#o�M3,�Y�"�}DO��p7����΢��F|�lK�֕��63����^>���*���_{菇hK��הC�v:����)��-m������u�^^�(ά�v��A{|�Gy��a�}�g�=3�%Ǧ2�1)K'��3���ve+��Geה���u*9E-������~Wr-7^'���3�;����V�66���l�_�׬��߼�U�����$��2�v����m{o�>��]{��~��>�1{�bd�0�\g_��(���G�*A�,�_��l-�V齹||���_�����]�;���1�W�Y�VN_z,���*�}�yQ=q�nXC�3||e�p6t;���ۅt��9���s��:,��.P�z7�.ii���w�߼��U���4��g�����χ��l�rrN�!E��yh>{��p����H]:��/��
�S��O)�v�����yp5�z���w
]�U�k��AM��^����W)��ݝ�Z]�ܠ버�I�:��Ue�
��[�����i�"�t�`)�\%+t��B�pn��Ѱ�Z{9�vN����Y�{<ů�/����l�ȼz��{'N�^v#q�=�l:gӍwv�ץ�5�OH]k�R�k�FS~��z����Hw��K�Qn1�=ῳ�{��NG0�Ɖ���c��u}j��[����Dy�z{c�^y�CÐ�����m���ȭ�:�h��*F�D�;��x�A�P�:�F�X,�uP��W��o�x�B=+ԽTiGw_9����Jjtw��T����,	U�e��_<�����Ę�߁j�I�맙�7����ޓ��;���T-pf�w �(��@�,)^3[,c�������w�L�h�஭yi�EwR��!��>��w�):z�޸;~�f�.K4�����UW�-Nj<c��ypI�RG�ϼ�a����z����c}��'ў���~�TM3%�r��T��ޘQ���o��T���٠�>E�9�oz����3�O����n�\�[0.} v��9�2��R�N%��;�G�G2_W�ڹh�d%p�n<��������z�>kF���ۚ͸�	�V��f;,IZ�Sjc�`�(]:��h��t�R�W��ؠ���#�F�|d޴6v^�NVJ�+`�(v{�:eH[��T|����M�Cjrk���^���rc�Q
=�Z�����]L�7O��Z)�$� [�th�5V�NAwy��N{� 7P��_��+��Ѧe��8*_V��˥��y�G?uǮ�}i�ō7j��_W����Ϸ���|�۱|}�&��*h��=8�JӢ��}~�Ǳ9�`�z\�L���%������g���ь}�Q�����znI������B���]
�����K�8�;8=���{zP�ۼϺ�k���)�<��P���q����,ї�5��>NnV��1�yE`���ϼFűz�����9�V3)���ϼ��q����!��	B�"q�.��)'�7�Y;�f�>U������VF�`Mz�(w/ޓ���}2l�c�Syp���Okɥ߽ʎ���,�
���;w,���xk�=P���tz���t����N/\���;2���e�7����y�qݞ�B��$踋rIꈙC�O=3��B\�J�^n��{�.����>����~�>>ӏ����w����C��;nH=QX�c^l����_Fo��vRa���NG�*x�R�X�~���7>�Qg���{��4��i�4�����>xUH��U�����r�uJ�r֋�>_k���Y~�>��k�p��󬘇�\��u����<ѕ��u ��,��k���5Դ&Y�M��!�c"H�����JW}��/���(-O��2k��R�Rs��u�}c�K��M��p�ulν�7 �WM���m���`~v�'�uyzq��O�޾:|�z2!{k̭�*:z�ԁ�p��9�r��ď�ףfz����h�@���_���Ҽ^�u���+���yb7>GTC�!��h�9`R�N�tnu�V�լ�����S%� 9��"b[���G۬�r7����M�׻F�P�ڟzv�"o|��K*�=4q�D���y���s$�nKf���_�
ϡ]4xv���x���A��R'#��1�enr�s�Ϣ�}j��O�>9��s��>�
�4�d �H&��s�4%�� ����'�"�{d��ס�|o�������^~�G�>��PFWO��(2{FL>�#uʟeއ��Ș�q���\��Q����ѷ�\kzX�]�c!?]ȿ����o�����^�/�� ��&�B.cj��{Z7ۋܽd���p'tú�n�W>����8gU׃s>��~��/=ׂx�E��b�M�k��%TW�z=�R2Ԣv����C��+ȉ/IÈ�֯�"%�{\���<���b�����ʛ>�˟'u�qmy�ӕ)c�ŗ>:�G�m����߃J�~M�I��Z��إ��5�G���yZ&&�YX4!�vŽU0*f40N�!�F�o�Χ���'m��)�w0�$j�x9���!�l���4S���78�-�d!��̸��C���N�s���C{)x�
W1��� tK�Zf	`Yt�fVtuf���F�>��3�Σ�*�5��3�x�8K�g���Q���;Ӓf(�-x^���i�t�%>�>�h�x�X>��{ǲ)���Z�TFvT鸲����ռjĚ������N�=[U�U)-�Xx7��E����܏z���]!�o�W˲�O˅>�a͘��&����� ��:�!!��i���祵Q�)��!z�do�|�纈|�L{Lӱ5�ޝ����R�#�������D�_�O�C��a\-w�u�u�ܷ~ӟ/H���Q�"+�^��<<D��S#<�v�� yNĖ�n�����U�G)�\N��(i��h�U�/ַ�ϊ��|w��z�޲6�4̲Ag"����Anx�/ō_xܝ�i6w�{�Z��o�����u�l��u6G�a>�~��ۏUx�d��I���"r����p=1P�������ZW��Е��������W��|}�g�#�9�^}�˘�R�LDL.ք��<��U�����=f
S�v#.Z餦|��-:�[��w�gݷ���t{���H*�� �"��"�ꂠ��
�+� �"��A �P��/���"��
�+��*�� �"�삠��TW�*� �"��*��APE�W� �"��A�T_�APE �"��b��L��/��T>ɿ � ���{ϻ �����>�J�Q@ P � � (����$[0
$BUEJ�J$��Q&ڶ�p�P�Q%R"�)%$RR�*��&F*w v6ժ��(Z�[F�2՚��f���˸Ԩ�n 6鍱��Q���  �  wgn�i��F%)V���T�Z��lCJ��ZY�[lĠE�N�+k&�Z�M���X[6]����M��E$7R�9��ɒ�훷6s�\�1n�''m�;��j�qv���]�
T�Cpr��M��U��S���v6��f�e��n�ӝ��8;-�I;wiu��(�����m�ml�[[Q���(Y0i���Q)V����V�3JYkIV��L5�j�5�ҥI��Z�Q�EkU��mh������%������-	B6жʕm���Ta$�[�     L*RR�� ё�d�M41�"�0IIT�      4�ɓF�� �0F`"������       �&MLL`��I��R�2i�<�1MF#�h�CdM�'��>Ͼ�W��?Vs���Ü<���B��a����!��%@�  ��I!XC��4�B�IfO���?���Q���?��aE	�
:�BB���!�a $!$>�ۯ��g `������������C����,*^���iQ��K�������_������E�/���_��߷���8��̣��S�FV\�h/�%��5*��AfK��f�3 �����ޠf"rR���J��;qj�r���'���<v����/C���W1�|y�����q��d�J�zN � �V���8ݩ�h^GAS۸��X���J�[L֔ձ����#t�mP˔�5����YHeU�2���(�jՍ��@��o%�[��b�e�@�,�� 9`	���LRَ�yG��юL����^e�r��3�.��r��,�IQ��*�>6��tg�c� 9���f������A�f]�(�rt�J��R�YgF�X�y%���s��[H�o=$m��7�/F;�G3��U�fMT4dq7���-iƚ!��G�+.�L��4P�zl���w2�Q����V,쵲�Ae�ݐ�2+wv����m�6��'����)
M^�q��Mj�Dg/$������6��Vst��XP����o5͙��jn��W��3v�i0i��+ٛ)�pC+%� RXi�(���X)J�1o��˲j����J��K-��k+YN�ܫv�^�5�jL$�Ytތ���	�Y���]L�ޖ�H�b%UҤ��jNeX�e���c,̵���X*��2�w�B e��%d&r�u�Ӵ�V��VQ��T�`;�4!�*���2]�p�Ak��:�a��CA6�8���fj�`�e�v��&���Y^���7�`׉��ڛ7U�Gu����k�.J�t�n<��홆-k7�d��T[u��j1�Ǘ�Apm�m-D�bl��{����7l(�Si�Z��++�[yM�KE�"���$��U�-I-): AF� ي�]�X&nchZ�6't�0 3f�4���a�D8��׵��CB��2%&�1]�q��Z�	�,�u�3s���rK��Pfڛ��1^ٔ��(��i��^��Ƞ�V��2]�QA���_���M��iX[:8�NЬ�c��Eﮉ<ݠNfk1�yn$U����.���.�Ǚy(
ƪd�vj���R��]6���F���l^i�z�in���K+4��f`���q�~[z�K�*� �K+�e�*�Q���*���E���^nn�.
����h���2�`�n��2�ɥQ��E���sU�Ưbu-)xP��I��.M��j���X�xMf�e��LHc�*�o$����@Zi������@�H��ϲ���Œ��f��X�-�R�^&�1bhV,M��n0���kf��A� �9�5r��++d�1<����0�ZK��/u%G]3oy����썄�0����k�;�H�p��{��Ea��lm�d�;�Rˠ�5[h%Y,�(hw{�V���i�Vn&f�e��ܛ�r�&J ]�X��qV���*�gw@� ��u�glu[7����0`j,>!ȬbmF�n���<�e]#@�}���y"U�(1�b�ւ�"�י��h�mi�+�Ҽ����ڼce1S(X��-^`��7���֑/j^)��4���3�oa��36V%�#�r�+ϵ�f�StU��T�)Y;w��Ő��b�YP%���e*���C9��R�ƅc�Z���J��.b�T���"�@ �z�8a8L�h��@�N�=�w�q:FJU������%XD;lZp\��t�!n��ٲ�ʖ^�j�e���dʅ_�td.�1�+ܻ���6���vq�UiӶ�21]eWw�S=WW�wt���!a*�V�4q��Y����.��V]���M��Efi;�22V(�[t6MO2U�k 4sj0�[���pb8eD��	d�x�Z�uz�q�t���d�20�.^X�[In�9{b�ʺM�_ƌLI�8�� j�c0d+)m���Ѻ��KwD4�
�9���6R��ݬM�t7* �Mõi��ڎ����.�0����Qr��`��l��Ke�]�F�S4��� ���դ�$���Q�kn9�� ��/�,
u�/ab���XԒ�;s*�O//���R�-��2�e�z�۽�saњ�waOmYhj��$k�0��$Z��Il.��T�����u�]pc�����#VްA *��3�������e
�+;m^�)��%�X�v��,E�\���J.��ee��=�D���.���h;��:)=�IX�U����]�7礞�6݉[�"52�5���(�L�
�Y�\ɗ,+��!cAi"��ތ�6�ӎf��^�!4��"j�{�m��<St1e�+�_X8[�:��K�i�V�����gu��h��nɱ2�hSp4�*LQ	F�[z)�`���h�gb4��G0kMn�/0*53"wv�j�lT�7Nݜ��Pr�\y�t�y�8D���!�і�-�B�Ճ�z����ba��v��L�JӘ\e�f����C����Ħ~�̡1��\�pH˟�C�����uP�)�}���֍
?�A��� �A$�&TZ�ʖ��̓�容�r�M�:m[��P3-[�H��k�|��@AN��v�����SC���{ ��//��mnγ���:"��k��k�L�[�%����0oD�.]vc��h�U�)q�,����e�ǺH�"ݻ�,��!��ڢ�w�O���Bok�w+��bOMͽ�.WkW�a���V��[�휊�\�۽}',fJ�F^;�{��Nd{8v"(��Һ��-wV�Ƀ,���p�}O � �1+��krb��u]������;��`$��dqc�r��n*���&�j7b��'ǻP�H|ي�k����Y�5Z}���5]u��!�w"����}w|�TN��o(�Si`U}�ؗmS0��tB�0�,��,@���K+��NۥL��\�����yG9�uh�����`��1���e���wm��A]1?���:o0�Yڡ�	��ن��;P)P߬���$u������4��X��.Ѻ���`}��m�keMU�;ju�q�E+}�ܥ���V���6�4\4��	L-�X1����,�y�:�̺k��r�4���I��E!�Y]�(����5�Gv�˼�$����]�B���+�z w�z�8��1sm�D��ۧ�ʕ�$�а������5܅Gd�7��õ&�f���*%�B��nb�h�X�5t�xh��B��@���QV/�sx��:sՊ�ꘋ���a���͍o��`�i��u 7J${�Lhxn��މ�ԣ*W9BPW�r��6��;uA|*t]�nԼ�¨u\��Xo����1k�S��V��	��uZ�������p�SCY�t�L�̧��\��-3[ءAh��5�(���Pq5 � ��"w�U���"Q��Y��>���B�˹�r˩�����&꽒�7�PZ��/F%�*P[���e��Ӻ�y!��}�������e
�(]�9e�A�ъ�N�L��vĀJ�вo���-ht����N������m+����yH�/-ѹ�(���w���W�:�V��6ԩpßt��dga�v�X��5�둳+r���ػ .��*3{]�떴t�k+$Jv�������.�_a�q���gw
�4;�ECf���9�*���q������9C��º�`#iR��Q����Fn��Φvn��f��mu�GA�X���=�U/��.��_>����5/�BZ�{]�`|.�9�)�B�>�����[���.�]:�\���%ΧV���(��f�͙i[B�pO)g5g�y]�$�AV�o"��I�:CYƉ P�C(�y/�un���r殮
U6���Y�dT�����ʊ�s/�a�w�&�-as�V�7�w@�`�� �Na��N�9#F���?w1%�,.B;��m�t��*�\��Ɖ4��K����I�Gmn�"f)ٖu��*���@�'2���2�'3���H27�^s��w��lt�.��3"�ԥ��o�Ω{�g�V$�K��ի���f&�U	*^8b/4 {�=ДNSe����i>v��b���dM1`����&@�v��wM.��Pw�{�^w^�k��h�N��l����r�_�NŸO]b���GE�kS(��}��:���ۂ_E�\+�EDb�b�M!,�}6\ҹwWV�w�tn�$e�e�.�8b�A[)��B�h��s��C]���v(fr�C��#^��� v�xm��q�6_8� ��ԛ|�d��C�]�r��2jĒ�g4�Xܑ=c��四�*ɣ[*fJ��u�90�&�P�L^.Z�S�u6��SgZ�Ԥ�3�z5�/-�˫��p�3�Ku��GjY��\��z���v��x@��|�0�)�x�s:�`��m.xX�t9�4NT6��f:��%�y�)'&�-�c�n�3be���~7[K_���}ZR�n+a����m�7-
za��;d\���`�n��]pN���X�[�dz�Ks�s1��M�+���N��e6��}�f:y$7�Ց6�I��|&G�(�sOkΩ�bb�/I�8��2���@��/S����h>��*E0��&Z����|�q�*8�KB�{oE����MY-i����*�a�A|]���<�j��1]ù��D2U���׹:ڻ���弨�Ub�R�Ȥ��X�w]Z<��|y��C'I8�d3y%����.��$�o�I$�I$�IVn-ٳ�:��-�]���;!�0�j�M^�sjp-KQ�&��L�(�%�v��yc�Z��"FL�9= ��I�6N����������MZW!��
�ܹ�Hp$�H5kw�^�Q�}��yǜ۲N�.�%Ac�4���"I$�I$�I$�I$�I$�I$�E$�I�I$�I$�I$�I$�Iw��^�����o�~�O��}���������B��L���HI!��d����~��?yH�!���3��>Ͻ�h��?n)�Ѣ�����ח�K�#����L]���bY�dR���F��qWq4�j�F�$|3�JXFg\�M�Q;�jff�p����d)�c�r��a�Iξ/�M2���v�Yȋ�&.���`}gh�l�\�i��;GJ���\�ϟms:�He�8��I����� A7����A6%�)@�U�iK�y��
�-�q.��B4�؆����Q��7g��z�>y=��Ѭ�b;�Ef]��,���ܳK��Է.�}%Y�N��V�0�(Y�wu��6ӥ���:B1}wB�xJ��|]'5��cv)h��es,���K�
��rT�%k5��s�{$Σup�aYľ�[�� B��鮥�y��R�v)�CzἘ*��ྖ����F}����r�:.��r��f�:�\`xf��TCE��l@ZE�_\�osQ4==ҳc�.�l2g��i\�5��@Vk�`����������Q]�/���,���	�,wsp�9icl��aA.	�)>6��&�"��E`����E�<��vt�J��KNwQ��`��ʋ[wWb����m�O�q[�
;+�)Ɗ�ُ�U��� X{��V���Rl_3Z�7Cw"����Y��:�i��̰�MȹV�(ZW���ϵ�j�nAy�Z�'�^g6V�\�)�5",�2�w���jeՕ�N-�e�۲.�����S�C6.7w���\)�٭Z�f������N�)m����t�j:�h�Ȟ_ZD<�0K��٩�����u>��v�V;/���-����K�1v=Ɵ;ή��pClR�7�1p90���
f�����!	�'R��q�7E!��˱Γ�	bb���W�/���c�����:$Ywv�n��A �x���C)>���}g��P��9��d�l���l=Y7�[܊��Ge�[5��遶H��	v�h#"�`ٻ��N��tl��1^RXt�����m"��j�J�YB�M1x�e�E��;�Di��;d�U��Qͨe��#��Ì�ΡR��sjuca�|1Gw�t0[���ٛ�j�k��2��)�nsT=w�Hm��}djwX��N�r��� 'x쐈2���Wa=��f�]Z��oA�:�JtVl!�VQ7wS�
]���v^� ��K��d�����Y����v�RL$_U%��<��j�@2��2���]�}"���FѨM �B����^������Z�*η�P��N�xMɵd:��%���/�B�*P�Kހ�ҺR�A�;��m�6�.����碚��к������zd_+�U�˥ ���ݻ��;��s~�6��y���f���<�F
NJ��X��F,�%����he�6U�.���C��1ԣ�0�L{��ª�u�][)`��R��M��Va�We����e�.���]���@wcPuÀ���J0�s�'b,��w������W}��np����]�T"�λ(ж)Ȏ2��-�цip-`���^R@I�z�搔n<X`�5,��+jq�*��WhǸ�Vh���슅�ҽ�Dh;Eԫ�:uv
*PDNƪKu�ڧ+qHm�4�4�#��3�-��}�t�t^$<���ڼ�U�`��q��h��亜��K�wJ��j�ŏ�n���J��P�Y]�ԝ1q�-�j�$B��HeqȖo-�;���c�(�F�����"��k�I']mN5r�]���wY���S5�]Y�4�q�҉"D�=y�G�9 �˽tV�/��|�o�k[� U�s����neG��72����m���ɹP�ҥѮʃ�ߌ5+6+��B�I�7�Xv��srv־�]3���P�+��Z�(��:lP{�l0����\)'ö�����6��1/*|.�D�R�Ӣȧ"��x`��&��9�*p� NZ`7�]ދ�����TK���u"(�2�*	6�k�F�ݢ0�����Q��RXw����/~�DB�u�R�yX���7�� k42�~A�5�շ9.�p��ھ?zh OGjƛ�WJ,�����dHxI�����ʽVUi��s�D�����	)s�0�[ՎN��y������d�P�ASʌ���ю�-�ٙ0�$���#���W�[������RD��t�B���Ԓ�j+�g_9Q�$ז��� )]���;�d�j��o;u�:�2�&�[�����[=͈�3X�P�\�w�U���,���`KpY��#]���n(6e��� :Usn�o^��i+�Zn䦴�r��&������	Sy��H1c�լ��ا^��8r�ۨ�D�ffih��[x�$�W�Ʒ�p9ԯ�����:G��m�s��W��M�=��!��]�Z;q�Mm� $t�z9����Pt�>���p�b�C���)���Ϋ���֩����Z��!a� b���h�:x�P���_4k�ߧA�G��-;Ժ�����{r�Y��B17#��{sc��x����x{�|V�o�Ɏ����u�ѽ��h��M�
�֙6{.�*\�֞���"�ۨ�7s�Fo^k��l"����tݷ�m��v��H]�-���}�!|Ќ��bG���-�QR���^��ˊp�wEC�x
RY�65&�9mq��Q��VQ��r1�ݰ���O�6�*�$j��钷�!����	��E$�	$�|��}����y��e<��@PE`�aC:Тl����Q��%1`�Qb(�訲b�b��i�A"a��,4�(�˩"��hX
(�M#��1T�n�.��Ri�L��CL�(*"�-�ڪ��E:B�vL1��a��b�Kal�%��AT���M�*�RKQ��j���a�?vO;�$�]�W��_B�a.ͳp������dwv��)������E
�7a��+]11ңH���eo�m�FOlr�z��{NSw������@��x�x�T4�P��<.�K\�����μ��Gx�D�@�9r"&�"�;����{�u�<e�]U��PQ'�ꓯ�Ej������:����7����P���ܻ�B}$5fH���5H�t����J��՛��+����>CM�P��
/5����"��fi�Fc*֚~�+O�%�lp��-0f�]�|0p�d@�b�;���v&��,Q����oBb
������x�]
�g�V5�U��zc�4��`�C]����ܾ��l4+�a��.�vwϧc�X�m��}2{���%��+�6��u��AQ���7O;��[F�oTu1n��:.-��+�u�cNǧ�di�<�)��ˎb�D��*ښ ��4��>�_�=0
���F̘Y��[��.4=�c��ܭB�����q�������k7	��eC�TW��gT�������C���.ש=�i��|�yW��L���Ȳ������7�*����_�d�ׇ��N�$�49v)�[�q�l�ͭ.��gF��;�j^V���	2�+1{s>v��*˙WK�q!ݯ=�drB�iKy�%�Ey*��s���D�"��%�n�}f;�Ĉ�*J�4q�ee(��W[��o81�Ͱh��ֲ��9g��W��|�=7�����h��k����+o�����
E�qz2^Y{�i�{��j�"6��[ ޥ�M�2�@��́h�E=���D���A������\��8Ű�tT/�<�gcR�ay�73e7i��y\�}PjzTZT@�k��5	�u�J�@�X:`�}����"='���|�s:�]f�-�X�h���f�	�;�c5r����]�j6��=˛|A���c�Ϡ��k=�m�!�<P�:�GPLF�A�ث<�ݦ3��vy�Ϝ(��A���4��zm^�K�53�/ޘ�9�c)^�E���fH�s�m>&F_x�;el@e?_-����ڧPt�ȍ绥�x0g�R��V���t��(�*�����[�u�;�t�O��Z��]��d�7��,�uۨ�+ܝ�<|�AY�����>k��2k��U�J��{�t;b�W�,Wn���ݵ��t�ǍU�{���.＄GgW���^���GOW���&�1ʍ���se�M���Nt��lk�}bL��`t�[�5�j'K��	[S��l�h�]���! c�F�Xx-��񡣢؄"��ᴑ������˶��#	܁�"s��<�Ѧb�&nR�e�̯5��$�<���QV�N���Z�FMf�|6���9�mx��I'���Dc�λ�q����8yDaw�c�۝7�!��d틦Ŕ6�ì��
Y���]��S5�i�J��RkǪޞ1���gc�n�FM�b��h8��:��X�R�O/�޹%�u����X�<�ݘ��}��= Ќ���Z8���M;�����ƕb��Ѹ��ZL�#;��_��t�r�l�2�^ފ\�7����^��u�.�3����'^�����A��Ӻi}4+�qs��(�v�	�Ւ����Y�ӏ��]6��';[4 �N�+կI`��|ױJ�z/*`~R{�=�QB��SC#�nQ΀zFPX]�wV���Y�F��f��RhK�a��VZ>�H<��vf
9�珷��[�����Mg!�s��z��7@(���,d���L���[J��.^�9�rv���Az�JGk9;���l�Y�.t�ψ\\{ºA�A\7c3#�G���k��߽u�5]���:��3P�Q�ɜ�-��՗��IJ�3���u40��WQ��4i �*b0�_,�Z�Nac�Ò�O��<��u�SwF��ټXJC��9��(�V.�7��6�
?�wYt�]v�.��/�r��3VŸaU�CU,4,l�j{S�ft�`���-Z�J�鮮4;O#	��,�e갬�pf^���}���q�X亦��Owd�H0w�m�YJ��T�O����0f��h�]im���j�T_*�V�J�k���3j����n�N�8 o�zy5)W+���=Zjز6��g%m�N�3��bSQ�E]۵s)��M�|qx<���`�cu��\"v�+��wf���'镑*���������C������S���>�D�쬪����$eM!�(�^�4�DS��![$�1��}���Xfe�q�C���e���U1�\�g�r���pY�z3hn�Z��6WX�^H��L%L���YC�����u�,����(�f�#
���}�������,Κ�L�M�6c�r/��o,���V19O��Ա�Cu���d��M�'c��j˝˦�����vQLV��ԯf�`!	�ls�w���$GJv�@���I$BI%N>�WxҺ",�4�ZQ�������R�*���f��Xa���V5KJ��.AE�2�e��&1WT,QU)��h�!B�3WB��I��b�IG��Ѫ��YE�5E�nUQLU�il\Q@�-�U�)�P���`�e1b̵QTQF,�INwK��,��J�b��2-�����������]����1� a"�*ꮡ1Ta�L1��@�2ͦBj������kj�}��<���abPGK�V
�՛:�P�;���z!��o�T]�~W�3H��2����w�T ½�h^�-92j�Ϻ�Ε��N3W,Ԛ��g_ٗ�.���#+���7���v\�}Ր����܇��ב����{���E�/�Ӌi���Y��8.�Nǟ��mH��{�Ie�R��9�5�Q��p���$�Z|7���@�6%�˄�л��S?C�� ���H]!�`��Rb�ų��m��_UG��X���B����=���'���E7Ѹjt�pd߇M�=���S��5�kR�0�]W9�	�y��x{�<7���]ˢ��ek����
�] ^�`P��e[�^q�<��- Mv}1�yS2�c'{�i�He,�G�����W�w� ����P��.��m��Rd�j��9w�@�ru{�XL�86�T�է�$w:T?=$���?4���b�����2ĄלGU'�1f�T��Qĉ�z{|:AI���\��Fn�6D�_��g��$̑�g!<�Yg0��wC��n�U�eX���Dd�
Qm�r^�#��C	\�3� ���.��r��������CiU�z`�R��ӓY�MtT�y㾠q���5"���.��rQ����@1E�7���"�@��Ē?����4O��0���&m��w�5��Y����_g��==^"���ISF�R�\����
�.��vh��Fq��Zp4 �h��w#���+��PɖM�,a!�2v��q�wܐ�!�5���{�!���u����'
N������2���9�B�y [�HL$���`O�!�
"Ԑ�I6|׷X���;$6�i�C��m `�Hm	������He6�P�`u��@����R>��}3-�3�� �:��v�Y��ju�.�T�@F��W�m������u�g?B��!l$0ϢCJ����T�C��@�B͙����6W�y��p4ɦu��@)$�	`E��Y4��!�&Rq��ϛ�Y���:HZi�4�HC��H#&	��u(@�$���@�w��zǵ��`)���`a�Hx�I
���a�a'Ą�Kǜs���!�<�X��!�@��� i��\����	� ��s�^�ϟ>|��-�l!�樐�8�d<��0�
d��i$�hM$_5�߸��|��I�C<$�`RI��N2B�� y$d��\I����~�����M':2A;D4�I&�*�O�CL�Hy$5�!�淼�����l�	H�ku	2�XC�$�i"�5u$={�j�|Ƶ���L��uD�n�0�@��N�C��!�HS�I'6�����}��1��1�_��Kwg�w���!��Z�̱�U�_��$��	��:�*�F���zv����� �_s�!�AB}����T�d�ʖ�:��!�k��Hm'I����s܋$2�hO2@���3S��C*�K9@`(C��/��/?5�C		0�RHx�@�q��@��l ��GP�X`,,9�U__g|�I�2O2LW�0�I�T��I-0�$5���ƾr�g�-{4a�$��O0��)$�X��	l) Y���!��뚿��u�x�HB���!�L�-!0I:�L'��$>{�:?=y�y
Hm,�P��<��R@�h�Y��X���g�7��x�����Y䐧�a |d:�Yi�o�$2�8�|a& f������t�a)�J`O!�a$�|HI�Ba q3�C,��I�N�wn�^�9$6�����&��]�!�8�8�q	l���>Q!���뗧"�
�{�K�hB�pX�\U���͹Ƈ*��H4�.ZӪ��]�w�o;�BBNw�Ϲ��L d�!��!l�Hi%�|՝��}7޻u��������=�1*�R�O��Y�"f���*bZ*�l��W,�2��E�s��1Ӡz��/κy���mk'�B��Ye=����aL���g�8��r���Ju£%��t@4ob�=Y~��9����)팲Q����v���&/�C�cXjl�{�;����9�<O�~C`��|qF�:F�v���D
p��?z�+J��'t:I��T�k/L��8/6w{����g�B�t@��E	$�X_��{�Hޥ�6)Z���G���ߊDaB���d�f�c�J�b�GeC��jq_1���r�`�q�d��d�h�%�>ȃ�o^,d��E!3V�5..�b��ĎW��}�Q�7�+=J�7ٙ��o�\���&�ȉqMQRJ������)vo�����VP����PA�����Y��r�>k6(z��2{�;3����C�d�B-[~�n�<�A�[�SMs���Xs\�6E�?l4~��p�^�YƼ���mW�f6��GG��yqzmI�{ˬ�����������ç+�o���-��쬟z�{�iۤ�r������S�fe���'R�@�w������������?m<���39�zA��I4��y{��=_ߜ3߯�(U�F��~�a1E�3��7{K�{�,�w��X�F����!mS1u;˴鹣*¨�Ƃc��A�V,��WA�z��c�N+���q�Y��u�Ե�}�Г��i�	��C~_��dJ�7p�OD|s�Y�m��.7%_+yLzoM�*�����=$���rR�.>\�6E�MhR7����O���l�>׶�cݨ�W@������l�9��qV���V��8藅�[N�lB��;M����iGZ�%��7*��!���]�jK����՚%�Xzv��L*ٚD��0
�U!A�եh
.c�+����NX'' �V����v��o`2;Y��$����5<���ت�ӗ��dߎ�J�,Wo�Bk/��:_��?_�V̈́k�;��w_-�(^X��s���[gS�#$�d��V�
�P F&�O7�R�ّS�\��gN�
;^t$dD"V��ثw}כ)G�E�S�o$��Ma��˞ɡvukY}�0��2-����������j�yC������ǎՙ�����#�QZ�E�e:�3�qJ�9�n��w��aE2.�S.�Gp���wx��m���'4r�w��"Ea˹�($JĹ�$$�U����,{��'��c�I�Q-�$�u	m8m-��(�
��a>3�-U�,PPU���a��P�PYi��L0�@�(d�C�6��=s���C��oH���-5&x�Ԓ7]s1ZDc��G��G߭{z+F�~���S�)-q�����Q<!�"���4�8�*C׸)��� Q�X'+Þ�z�J��!:)�]I��eEG������R}�m=������G�&-�0fx��U��{%�οS��j$�6���h�<9�Ӂ-༁C�a~�Z���)(`�D�l���Z��*�t�O�Q�3���mr��٭�C��f�C�������x����?�53�{�p�?��~6���L&7{���ۤ��*�ޟg^���Ȱ��tG��CN�"C:�yV��f����f���{g<aU¹ud��ϸ3P�=��~����`�*4b��۴���ќ��"�jA�1��
룒/q���QS���d�:�|�+�'1mʱY����u��('�[+�G'h��������m����Wʈ�|�9x(1�M6����6��e�|r΢E�H!1��v�S�df��>՝F����Fu�J�5o�yL5���=�B@�7=��1΢�^���(�al���,2������k�n.%c��vN����'lߤ#����kpud_��q�8��v�ҕ�gwc��Ap�;�:�=�{�eoq��N�c�����1�C�)�Q(H��:|7���j�}Go�ӊ"dcj�y�\���Y��)�,u��&�Ga�%���,��m^dO`o��.|2�wd,���,=��q_��w�A����^�H�OGa�I�)"�a�<a����Y��M�{d���GYCp�hÐ�v�*�wNqj��X��N.�Rk�f��v����K3Yq��E�T�W��f�^>{��ƭꌐ���4���&i�iW�6?����>Ô����Uzc�/gE�{�����Tw��y+��I��
�x�җ#xU�ˊx.��Z1�Oߓ����}r���i�D���ҴK�.�GA�ص�t4т���n;�Ow4��V�D�\V�;HĠ�O�鐒괣vE�B����Ͻ��G�y-�d�+����9�o�I3�յGnf	�8�+�Ml���Zv,]Q,@V�׃ü����n@�{V�Cq]{~���݁v�³2�Is���8��gB�Z=obW��׸WG��~�2�p���~�ű+:�񞹫q�6��ς�ڂ��y��c����Ϻ�(ݶ:��^Y�˅��+�L��'R,�!�S��4����UW����ڂ6��=�(�;?@�^�q�xH���-%�w�^/J� �����&s*��Ӈ�~�xҾ��3���^D*��쨭D л^�m���Y�v�w���/[.�u���� ׼�}N���޽|Wx��53L���y3����\]�5�Y`��ɳ�_[���}�n�)Ni��<1/vӭ�|�~���/3��H빭]��	�_]��G���C5�ϫ�q�5TB13�s�<��gP�,9���J˗N��勭I��3�|��h�H�����|��借!�\�X[+Pd������y�B�����1�l�w��=���AǙ���T�(yw!��d�w{����9�s��Y�{�f^�s�f�3G"Ԩ����mE6qm��r_ix��y*I�/�U�W����H�~����٥��!Y�kx,m1�v˰/�o��x�Ht�e� �p��N�:ݾ����]�Y�nzLu:5Դ�����$���j��4O;c�7��ZMLi�yܽ�N�p�����ݜS��KXk�G�E��ᒡF]Qѥ0XߎU�˴�iDZ9C�ܥ6�6v����c��=�dN�ISxm����Agu����c�1�.�O�pm�n�Ϳx]���İ�x�P3K�~ʟ�;���X�m��1J�.�K���)�K����%��Ĉ�{�)�bu�!�R��y�L���3�����S���E?z�Ru����� r+se:��R���~�7'��;���(��0������S�樭J��@6�������mZb�o����0�룕^63d&d"�:Mfee�+�+�k�w0��S�pM_��Y'.���b�[ݶ���;@��E�����\�W�1j*/^���,�a�0��zn�'2�d�c���ڸ	����f9ҥЮhj��v�+�5f���ê�&d�Gk��|�00�Yc�uL��]3��	4Pr���Z1:n��O�¦������8ay�	�uj�&2���T�ik&��=M�����z�^���?�:I��0uvkzoY���R�ٱ��u���^a�[]\�V2G-骺��q�/�v{Svm��$F���K�^����{��.�1N{S�.�ۮt�����$�����Ԕ���T����.>�٘��$U�yoTԻM��q�θ�
y�̉�ghl�θ��Y���V�����w[������u�	�'k��
ˎ�>2H9�͗��-�о6�-����|n�����sU�]��/�C�hޓa��y�����������u����9("i��a- a2�["�L�,���_��i2�i�AA`�,�Ȫ*�tXhFZJa�,d-"�E
��i�4��ED�m�h@�[$�HS Z�c�7�O���*�;��+BX0̐�-����{���������Ԇ��ͻע��݈���C�\#y쪶L��5�<��"� �L\L��v���݌��.���� ��g�ρ"x�|l���=\0t�����y�A<<�8���9��yzaq�� yv_m12AH����Ws��>��o���]�˪y�0�@Ⅾ�Ժ�s:��z�1�0_o�Tt&,���F���G�7�>��J~2*}5'�ũq�~�#�F��̓��*T ���d8ފAK�����F����F��x2o	�{y��6�E꫑o݃�N�����Y�sR�N!��;����ƣOPB`H�����<^�OS���)�Xhl��NP�YB�{����8Z�{�sx<c���!�GAJ',�uZ��q�+� ��ٿD{ȍ���$.v+�1��	X���M�����q�Ѝ��۞�{31yض��7��sOR$Z~��W�o���q�a!M��5�ړ��qW&1�C���K���Kѱ��B�uL�]�X�٘�n[
�*�㹀+� )w['�Ѧ��uﲳ��`���B����l�B��փa��Ԩ,.|_d�y.uc�֜�(�n�8�m�����B�l~@����K�?eJ�"~�v��N�&��R�������x�?Uə�S��k�/�tl��-�ܨ������~�1��3nKW�Xe�7��ݛ����U=��[3��Y�W�Y�;��ʬ��o��{��Ú�Tk-���K�]NMUF��%hlK��Ծ���^���p��8#;�t�t,���=V�9�*3�oM�O�+vŬ�3��B E㴁д��S�Gu��.u7XlXp�G
����M��*-��."�ۺ�G^0��_b}�aΈ،1&�E멇>�R�N�t���{��3q3k9KZ�<d榆�Գi�����"<�ԍ�eT�Kh���+�wq����M��ϸv�[r�):�c�w��c�R?Wսс߀t_�J�@#v�n���+�=�hW���c%������=o9g��g��;�&�=��b�U]����c�bͲ4�,��zp�\�*�P��^$&o�����}F1mJ�7T3��b��gH�:�Wns��o��Rӗ3f����=g���3$A�F�kUvS}�4z����J�x���l43�;�_�<�-~���>'L�ւ���9a;�+��|���Eu^42'i��m��XŜ��j��=�x��~�J~d[û�*��J՛��WZ4�Z��r�\:䳶���F뮝��n����D�#���3N�r����T�ȓ��"nzjc���GH��9P�4P��P䪩�&�%ְ�}��:ywD��eEr��N2\���������غJ�"�tr�`���G�;�\f�5�i���w�mxf�K@��ވHf��0��>��wPʦ�8�i��r�NZ���O8|��ڢ�㤴�z���޵��=t��tM�^�a-�Mg<泍v��P�c�q�䨱3�p�غ����+՗:��Df��Yf|gMD4I�a�O��ʋ��>m���B]e��"��r'�e�����(<u�<�7���{�����ge�ن����b�~N;[��}�k{�[�Q�۔-ɉ���5�5Q�[FP�6��_TUП)]���]K�T�ި{z��y�ҕ�lV(6"�z�=�
�Z:�iޢ�v2�n%��=�>��������-��nX��.���f�o%�$��œtU#�2�-<��u5��^�yｬ�u>33�j*au]W��d�&�����O��)�Q��;�ZfbeS�������J��+|N|�}�.��Qr[V̏�n�j���
0�9i���Z�+��)�y�`8�:M�J�n�:��sٛpњ:�ƹb��Î�Nُ{�e�M�J���g�8�C�4ӂ�

=�A����^��GM�Ø��Rf��S��ҫW��YV�Z�{�
��-Ck,k����Ѽ�T�Um]�����z
9�������O�'�Gn'�_LwQ�}63]sB0e܉�rz6|"T�TL���\X*�l���^|�NC��q_Y�x�=�Ѫ���t.x+���pW���y���ߵ�q��4���Jp�1u�<�\��o�еu/o�|M�*�Ъ��)�w
@���!-�]��ז�AHѓ30�t�@�ν��5���l�ϭTרӜ_����S<h��q�I�I�`N�w4R���=P�@�uT��O���Un����j2����u��y�|�b�A6ME�N��*�c�/���BJ\��d}&%��#jKKl����d��Tek�H��E�e*^�4�=6VY��U���z�������c�{�Yx����Uo�b��4�1#����$���>���[D��hkۺ��.�SNde��t�֝xF�#���N��f�(G	u������*��hC��*S*�^�4���ռy��f�e�x�L�vyd�n�bYz��o�wKuE��y�u�+C;]�6lN��-v�h�˘J���u��钋���k��@�<��rM��:me�l(�U��l���z���X����s�Wx�J+a������i�tEI���3_*�T���fR�4��:�8A��(��m��)�r�|�|�����Di��Bk��w[�#�N�Һ���m[�泾Ԓ��^@;g��-��jf�r��r��dw8�b���I����+XҘ�!D�����m�s��*�7v�e�:��K4�R�c�b�AZ\�IIN����S1��L� �
�M2a��$�a�hGii04�
JE�!Hi0�m��U�L)�V��"��e-d/5%���p��C	�WJ@bL�	2�=��\2�L�=�d�>��^��G��V��7�k܃u�N��G��,�]�^�ӏ;܂q��!ײD�3��˘B�\�Lt��*yy߹���Q���R������Ӫ��y�n�r�|>|Ͱ�J�L^�{���
Q��kܪdϠ~����,�*�STu7��{t[�Q���hw�^t�X��=C�j����j��1Y�������s5�޶�v����;�oY��ǘ��˽S�o�-6��Q�^{�Y۪����t?�<N�`����j�����Yt�ٻ��+������:���p��j%�;wc'���w vUW`�Z�Kko��Һ7w�d�ӳ\�}�{�+�j.}����t$ਛ���Z߳�{e	�{�x��n��9*�`I�5��� ߶e�DL�註��[0f�!U�Xfsx�t���T	����ٙ�*T�����J��xu��񖄿�G��.��^]T�	{�����J���Ϟ'D�5�\'�5�gim]yBި��ڲ�gTZc��c}�!��^�h٤)hU?
5�W]c�kd�u�,&z�Q|��Şz��4�����V�άc���U�����b��9�����~���m.��u��r��גqm/�ݼgş|i2Ӈ�]Wcvy�ѽ4]|q^�g��XZ!M�f��v��ykǣ�t�`����B��������㾤þ�*A.��^���+����r;/i^��6y�n�|�/�n���3�Ǵ�[޺�_jf���t��r�<��{7���WxPA_����U�.��]
�.Q �*:�|{&2\�uL��2nu�c4t,냆�b�xL	�n�\���u���o�ި�8�6���6%��:��uk=<z�1�*Ν�v'���C����5+�H*��Hh��D�x��ykz�>���O�ם'���>&�oQ��J��\s�5ڇ_��W[��]��Y��t�ۏ	>(��w�]P����ٗ[f��o�x�{}? ��u��+�%
����:�4v���{��IN��S�D��FU�S����	}PT��A�k����&+��ΰ=��2z^WK�~�Ju�A�Y���zf�迨���Y��r���Y�_�����{ޞ�i�v�MUhf�Yz�3G���\�g]����2���S��3�U]R�'�K>�����/�Ni�zg�-�ٔ��zђt��k[�.mhM s�_�зS�u�鉟vW�����*x��Mfk\�o�te�c�1�ݶ�S	n>�4[��UU����MѴ��x�v�w[M�)^O_y�q��k�g�7o���m�(3��7�Z��ٔ�7ez�7�+�Q�y\����:՝x�u2�ڣ��X��0H�x�[F�'%L5&�&צa�%֑-:C�������h�R廗��Ԯ���-��3��C�P�3M�\�r�\2��{ߩ��fJ��t���.\�+��g;�,�{}�Z���Iz��P�9vU=����2�c����nPE_q��U8�^އþ˭���Yf�m����쿙�C\���nS)6��|t���Cn��%�y�wZJe0���a�v�J���g��2]��!Y��Vj�*�ϧ���OS��5�����j���`�Һ������~k�Y��i_�M�ɕ"L�
��x�C��TL\��uO:Ov�<�Rq��y�7�V2��ʧF��[�p��׶�� �o����}�;1�*D�6fc)�J����������y�5��Lj���I���h�&ܛ��"��U(����]�޺<�m�Or5�r4\��S}�lX��;������GW_YY��q����Z8ͦ���o�ԴኽV�P��G]�6�xj�='�'��K۪�r݋7G«1���]`�#c+o�eҴI�6���ы+�����[���;tR/Y��<E󬛳�S~�w߻����2�fZB��r����y�mw>�ޙ[~-Tq�l��ڳb�Sövz�>&+;n볌�����D�T�瘼�}ް�O4��ٔM�L��eL��X��P�g&��
�4`˥u// ��t�ҳەt�弖��1]f�����gk���\��G�[&j�fg[r�iټ�_��=���g�6�'+Lӊ��,M�S���PCz?&�Ȗ����l��m)��3s�S��d��5��(̥�˧+�2w�9=)f�i�+�3=0{�L2EA5�A
��B<���{f
wW�UW����=P.�b�	��F:�s����Q.��l�q�׽�ִq�0������ �7�h���A�j�a�VtW�lU���6��Eb��<�q���F^��ԧ��+Wta5�`y��g������W����(ׄLt���ˑ�f���+3��|0UL�4ue<U['��n�7x�+nd��et�vq��r����Q��P������V��+_/��Ȝ���{��x�yej��8�%�c����NSg���yqZ��yg-�L�Ob��Cbm-˃�S�6�p�]Ao�t�|n���32�eC�(p�S��7Q���.s�*�ݵ�1��QT`����:T��Q\�<�a�����u�{ɧ���KWJ�����_�}{u�L	�f��|DLT�e*���}��y��6��汎s������Zm3m�^T�^�a<����K�{+��.��K�h��H_�:�����w�Z8)�6��T��s
�ц��[x��b�t`d�)��y�.-:�7]K=OʱѶZe*�Ɇ�\�7����uɪ�y�t���p�cU�W5A��\1ؽ�^�������ϕ��^(S�x2�j��AF���8{��[�����a��,�kI�ўW^�ִ�|߱���0ۇ��6]y�Q�÷z��s<�&/e�1E"�4���]+U��~o��t�⯭��f�X���}�.�>ᷧ;f޼�l�ctt�Xa�wY_V=�s�b�*��3Q2d�r�:#�\#�I߅��ſ�X_��pd���֚����xqE(�����΃O)b���ڒ۩ͅb�(��P���-W<��"�e��ax���4���W�0�A쇩��[Y����Q����1Z�f�{2Žї���o9�e
θ�(��ذ�������"�ɍ�'�rK�6�V;���qUt��RW��*�XU�,��8V���w�S
nl���4F�+B����oRwW���^��.�S㔶�h����д��H$�.��h�����^6MC�h΄���>y޿6U�tk۹�@"	�3sl�R��u��Տb�Y�O'�4�_W4�m��
v��3�V�(o�:鼠�1��Ď�p���&X�Z����2(y<��VB�[i)ܳsrK")b�k�*�ݝ8=w��3I�m�����]����v�w֙����3d��ܬ�zC6�O�D��ӫY�c��D"��jQ�Ѳ�R�ﻊ
��9G{�k"�&���'F���X�'
��%$�%$���a�)�����iV�J�H�ƈ,��!b,X�H,U�e*����e'ƕQ�%1ZJ�UETqE2f��Qp�`a�R�UuC��Q@�R�"�*�X��Uj�[B���,U��(̡�[M4��b(����fj�a������k?3W�#<���M��Z;;=?��N�w�{���t�z��7�5���5u��cà�/�3z�\������Сt�w[ujEDaS<W����²��U��̪8���ڮ��8|��jy�����Ӭ.��a���.�ڻ��w׷.<N����3f9��N�Mv���^�ۻ��X�LuR���ڱn����j,�P� �2`�T����M��]Sψ�v^P��N��2�m�eԿ���r��Ŧ����w�������F���7򺬱3n�u���󋱛m:G�W�q�i�^����vU���I9�6���k���%e�݌
�P�;��DDD5x�wt�ݑ����h���
͋M��fV`���v��;��sTQu�e-��ڮ���m�u��|i薯n����W�L7�Yם��SlҦk�q�(�y����׀�\�5��zrc���F�VUy�w��^��]z��)�ݔ9J�y�7�[²�;��PBS
|@�nׄ�E�4����CuG���k��5�9u8!�ݕ�x<�^ۨ��I�Ψ�o"ň��7�~��U�ozN�{�a�u�n��է�C�q1����7�^�6e�{�\��s�Uޖ���w�k��nRz��G��\��"�weq<i~���}(]m��e�q2���<�KeT���}vtƮگ)�>��|j&���GaZ�9���n:\L^�^>�{�J��1Ѵ&/��w�N߫��!�4�{�߽v���q���e:��jq�A��Pa�����T�S�VN�km�&�s=ν��*q+Ֆu�u#6��U��|��얙�J���w��gwu]�X$�f���FV�N�SY��/8��s���ܦ]9T��QZ�=�r�R�A���ns�_8q�羫u�F�X垼�j��Ƈ�w�x��M��2�V�p�|�UQ9��:���Q���6'�&]�i6�7���{:��НlN���ZY���l��uޱ����g[-�6�7�����Y]���MC"竼z�����>w����;�/���1�<�����4�|�4��&�\W�fb毸T�ܽ��|���)��]7�+�Ξpb�]u�(_��M���[�C��򫕌w�:��+�uA�U�{E��x��M{5�oY��E9iⴍQ�OP��)�����^�L���P��ٹ�;7t�&:$R"/��&�36�hY��=qG˯Y�[J�G�f.�aG��j�ыT�4����)߽ѽ�uS��U��HP��K����5b���V�I�nΠ��-0ᶙ�V{��s�m�B�`�z��;Y��yB��囻��v���P��u��|�No�8�������}֧�p�	牫�Jt�L���k���^j�ɧI���Y(���Yh���ˮe��~���u.�b�ۖ�!�X���5���N]��=ʜv�ѳ�8)�S)��k�qto�w~8hp����h�T�U�����E�u/�z_��Wf�4|6���U;�԰uy�A�'0+9Ô5a�szX�[�u�i�݂^�r�)m.�8M�������??�Wx�_��t+���R�*�\:e{[ۜ�N4z�fY�Â�T��͸�5��{�9��V�wED\��Ƚq�C{��ܺ�WY�S���_Լ>����w��L��ѷw��yB���Vo*�p�Vy/��ڨ֬����4z�R�3�Z�}�$�e��cx/շө�����{��8v�r�fUQ�;�	COJ�\ˑ��ׄƊ鹎���OD$����^����^_�=��to�.�묽խ�K�f��l)q�EE.����O�n6�w��XL���:��c�	 �~��a�Lj��7v��ɺ��Ϗ��|ӧ���z����y۽
��C:p�K�����"|g�Ltķ~�c��}�k:�pyRU�u�]�O�݋�q�׍b�����u8��i�he���.��lcZ��
x+l设����;��P�hG��ӼB�0u]l������O��Q3k,]k[�)�M�7T=]�a:n���~�ZE��̻m��v�%�
��7۴8}dR������P6+,�;��xzZ+��#v���M̢]�X�qm#黕bu��Լԝ��&Njh
�������B�{�AGu�1�Ez���ͨS]�0F�F�s�E�d�5C�~?U��n��_��M�L�R�ꕘ*���o-�]���׽+��n`��+�w�L]M1��۶�S)U���3��Z�����f(�oe�v�kwM�+���8c�X�h3]�r��9�:������s����wT�B{58��N�1�g�G�vY�{\N�����}�.���_;�5(��w@�Kٝt��|��X4�|9r�h�����*��[��ZZ����$�5ۿ�8�^ٺ�����Ŷfl�%xAJ�'Wk�y����~�s>ᤘ�������L�v�ڔp� L���7�7T�+�I�t�4�i�0��s�c�}��N���P��
�%
Vi�uOE-�e5��_�/o�`v.��y}�2x{��Ϭ�-�.��L��w�;�y�w6a��J�;z��5�,DAY�t7�~ٖ}���n�+�u˘�>Z)}u�-ۛ׳���7^��a�h���p�,S�w���{�/9Q�i4�4&�&��u)�7������]M�f4U�c�B�T�j~��G���^c�"��!��"�TE�ܒ�	Gkq\/��uh���
]��y+ZL}P>�:���G;XN&�&;�>[���3X�*j��ݼ�S>��_�=��21���:UWF�ѿ���J���%�ԫ�=�A-���5aQ�V(���PwT-���\l���^���m|xW]]��۱f��kL��ϲ^H�WY~����tm�h�����團m/�y+������Zb������KS{R6�g&	��Qj#��ю������1���a6�u1s��ۣɱ�r*���npWkp�e���e��F�D&o�j19�$�)j�6���;ՁP�ص��L��Y"�⠬"���[Yb���vV;�{)����T&�Ok�_gZ�
�ʲP���Ӵ���D[ �OV*�� �`L�o��{R��`�a�\*m�����v��*�E�[�%�5���	���ŭ>yR4�c�ڋwX{�]�R,��+���H�y�.Z�� �-��~�����:C��+����Rֈ*]��`��>Rd�,�G�t<����ǣ�o4��H<ss��p��XN�e	���c�!��EYY��<��RԷ����$i��ܫ
�R�k޾x�$��Q��jwPP�е�8�n����L)%�4�9�ӯb�D�r�c�-�����h�j�l7E�{���E��3��P�É�ߐ���f̧΍f�dyY�Y4�_I��R��9v���ڤ��o:��R��x�e�m�.U���$v�����-tr;�Eks&�zZu�I�V������l�$�zI%� � �wt ���b�b0R%T�4��bRS5R�@bDb�b�Ԧ���Gm��EF�U����QTZ)Cj�Q�*-�nġ���*R�i�c("�QB��*�@�T\Rң*�P�S��
�i���EF��RUS�
U���Zh-�U��EhX��"�b8hD��)U%(*�*(�a�[��EKj�����K��qs�Z��hVxt�7Z"���z5,�P&*f}0���3��#+i(��������pM���s�G��IU�@�z��5��<��1�����]>�Ȫ�:��2��Q�S>��3�H�5n��ҿY�����~F�QR��9��Bn����4|�!�(<�_w��߮�H]ɤ,�T@�QS}ڷ� �0�S�q�jQ��<�u�|$*���9&6��ܮ�sC�>}�`�Ӽ�1a�ޱA�kx�C�g�6`�ed�&.1iD˘�<����b{���׺;y�\!�������q���tF���D����'��X��I�j�YG���mM��}|z��迊=߹^{*����}����c����CqXyf�aY�F��Y#P�#6<�_��/�4n�]���G�U�DKFu�i�9{*E�T}�:���o�y#pl7O�=̍֔蛈"�ٛ��	�x���G[�GV2w��9���0��on�[|�$��U鿇���!l�qf�S
�������q�ԖlQ��^(oKD�%���x�~0�{ҡe<����΀�}5`����m�!���D��d��4/������w�1�4�ж�ɬ�Ota�������b���1��3���XO^�����'K|ƾl�w#���]����4�Jepy�2��o�^���+0�V����-��ɩ����ތy�bF[�D����VCO8N�v�c`P�3d�V��u��1�=�x�M���RGBe�؟#Z��'A���䎽k�Y�o �փU��\���Zrc-K��1�-teUU��<9�@Q;�z�U�:����|n���J׌�#ԫ��C�ky�V�]����I�����4m̽�;�al��S��-�UOÒ���zyz��:�yV+.���2O��Z{xuz���â�9�-�6�2u�}
�^�gn�y���8&��}	�a�g�)ً��;%	����:��OiZ8n�)+3zp�&���WM�j�%X�*@;�*�f���7rt�,\�Xfv%��Z�P��+bkM�}���c� /I�2�����^��m���m�WN�+tO�۝�]u��`���Q,�m�}� �ܶC�໇�p1�h����룗�
1N𭢜���Mխ��M]դTi�f,�F�p`�l��yx^ZZ $��)񲪪��SW�����úB�:��qhw�EK���T76�����o�����=I��F��@��Z���bGM�:��<�^O��&��[��<_έ1�91�bc�{ED��l�����v,�Ɓ#�>�9��g�B{Jd��</�~Ԝ�ָ�{�Q�h\H�*�CQ��*�Y�����X��25N�蘩�˰�K�u�9�ۍ�;MeyvN7��G��tp�Gbw�Iu�H�&f��zP���ց3��N�Q���D^e�i�'N��'�	��v7D�j�������٥T���!�2S��ݷ���`}��z�E��X��V�3�or��A)I$�I'Ӹt`~���_���?�{W�q6"R��U��1�js�����Qn���xaѨ5��3�T��~�ʽ<�E�O����ju��/{����ʖ]1�O�o��������%��FD�3ϔ�dM�WHP�O2$=�N��CGx� N��}�W:`�q<j6�o<+qE`t:��C=vv�ǞJ��5�����t�&���52��I@%\eߢ��ѳLG}�v>�-�
b��n�Vn��;]\�aVcQ	�83�r(�Խ;{�3��˯!���TS2�J�Š�鉆o}�4�Ł/z�oţKOC#������і!���?FG(���u3�fV�^t��z=k>EZK[�-��b���t��^=�k�g��̅P���rh��8���G�uҎ���wt!~�����HD� /v��Z]�n��;���Y�7G%C���2�f�(#r�0w��X���]�N�[���f��%s�p�,�x�ߩW��ʲ�4|���&���k[s�q�[�B�Z艟vJq0G�|Hl�����]73!9�}������+:�^����߅�kܫƳ]�����v��^۵�9uK�I��y
�mJ��X,�/1.�����0�j�����Qӻ*�o+���AY	n�@ǐM���uw��y۷���D��i�Xj�Y�ӮU��V:G(gQ�#���*:�mj� ��zv�s	�ծ[у�!�.�c�(���Cs�ʭ%;D���#�u.%�y�Z3zIM�+@�K�x�\�8�9N旵���-÷wXUcvuI'9��nb+��ڴpK�����v
�&t
�=�.�b���Y����+#�;NNF9zV��&.��۩�%�mR�|�M�w�O�j������QoD���+��R�B��$����3*��ΡۨwM<�bvn�*��q)[Z9��$$���|�TU����U��XL�7��'GTÄp�s��D�t��@��Pޘt��n��yO4If�5yw��e���}M%R��i��7Ӳ���8�����vîھ��&�d�Z:�{
�3�v�(�WZ�\/� ���έEj%E$�	$�P%zEL�&=5EG�Pb�(�R�b���*R"(�ULDc"���6���F`�#��EF�-�+)�(ėwm4*j�ꑈ��eQ�)F1Z����-P�����"�7Ea�QET�-(lh��U��c1T�-(��]4 ��QQ�R�U
"�"Ȣ�悮���yu+�@tHd�xZw�2���ڵ�g]�w�Axu���F����&�O$��m�m�|r��N�O;�;�������'R�=�-��mUԱ���$�8����ɛ��d�ז��Y�op�ķ�t��<l|���� z̵�3B��7F[&���W��*tN5�+,Y�6EOL�c�)��o7��9��B�2��S\*hK;�lņJ܎�����w.q�x�pb+ƹ����KLO��Ǜ���ƾkD���#���V����핖�����׏sr
�b�='�Je1��	�dC�/�s�e+1ẅ́"�ܳ'�n�)�9���W��%�������
���V�	�~���[e�^�B�`j��F�oR�\�sL�'W���!|O{�H��0�fS�n�F��nqe�^�q���KO��eX��\�Xm�,a�ٯ��N���+i ���y��'�������ݛ�	�w�:ӏ--����+�ďO �Iw�hV�z����3]0.j�7 �꺛�lQW���m����?R2�-E���B����V�2WLԲ��e	�N�`y;=���ٛ��	=�C��],��_r>��r/`��w�Avjv㼾�*�U�����޺&C8F��h�a��ɚ����S�"W(O������Zg*2,X���^��r��XX���l����C�@���0.���:�0�e�N�O�_�HY���U#���Η֞�J�,��r;^��- \�����-�f�P��&��R�e�>=8�t���4��WB�žR�/w��k-�ʉ���#*��l�33Ş]�/�[�@�{���������r>��j)ST��4a�H�������Yx���B@�@"���8�o�葟��L��T���I�9A�_q�/��ͷ"�"��&K���ǹώ8`N����9�VS޼��MqH�݌'p�]�����Y��NOd�u��E
Z�fh���l�����ch���1T��D�`\R�_{/.�[�&Q�n�ʷqiK�S*)"�jY�\�t��`���%�$�_�N'�A�H�E�ۍ��~�Խ ^���Q�ʼxCBW#v�f�uL�`��]5"	�n��ON�2��7GW6oh�S켳($���G���ͣp��̛����ig	qm��7S��]����<���,�=�8�|$��ֶs:��ۏU^�⒮c�9 ]ulRWv�O4��ĮQ�c�w�S�<�~Y�[��x�B�%�q(F�=x��_S���*!j||+��i�t�M�=����q�,[��=�xG�[L�I-��F��Ʋ��*�A=ݑЍt�UKbpl"Ü�0K�(alu-6z)6�9/�������0T��Ң/�6�0�W+�ސ� ;=�]ύ�+X&���n�9�h��3q�v�6[��Ip���w�&���Ŋ�OM��f��;(q~��I��46�<��v���e)�y�Y�:nv�;����G�g�!�$M������c��=�;ni0�����Z���/�3�6Oy�:q��vy��d6�����xz$t�p2��[��}�X<�Wz1��V:��|�V,�t��8m2x��}�W����SX����� \�uh&}�a�5�����fw>�>���;>Hf���س��î]��'��S��DQ��yZ�\:�ej����&3O>Q�����ލ�>J��&F�Ҭ��Ruc�}��j���s���J1��-h�o��7��@�x�-k���T���[�Y3qڳ�a%Cd��N� �S�ǥK[}!��
�N����M��2TeJ,xc4cE��P���s�t���܋;�*Lp;������'��δs@����^x��h�ST�t�"��͉݃v�ݛ��:��d쵥{���PQ��&ޛ��0�z�_a�'0;L^
��<#��X�hu���e��,�]�IX D��;���Ok�h�nr �v,t��MW ӍU4�zf������,�ju����v8J� ��V�c�2Р�eXc)�f]��V�d,9wBKC/32S��S��,\��:��7J�H�~�q9}oh}�:d^U��Wgk$���Ow'D!�l�A	t��;cNb?t�z�f"���,v2M�ơ���pdP+���&��̒���/�:�!�7�I�*Y�c���fc�b�ѳJ���'�]YS�������WӺ���lE�Z元��B&��Vcţh�=��aw��ӣn�����oo+���6m���n���d<��R�N9(��n��Gd���!�S�1)t���g<e��ͨ��F�T]�¬��+�y֪Q*��+��;:�Z����rh��iɮ�	J��Į�x�N.9�]����h�{o���%��WNg��&�e�fP���ޢ�ac�Lv��ꊹ�Ik�[:���\�M��O.�y�GB�,�a�l�kG(7�/B�/��db��#��V�Gf6�Y��4�H���4�K�xY	��Z�mr�Tr����q��1go@����E��I$I)�����X�Q�
���JJQ�*�iU��1AH��D�D�H����a)TQ-"���U`��j�b*�0T]4��TEX�,5TDE�F0DDX�1Te�VԦ"����YtVR���"��)��#U�P{�k.�^8s׾o��{�sV�b�?^���e4�t'�w����a�2u:�tY:�y�+$�vӜ+\��3;O�5_����nxuzd4
Vx�������h��5� ׏������iۺ�j<����K� �v=���������{���}�Q��]�K���$����=�3�j���p�@���k�к�B�NXsI_/
YN[�"��Ok��͉�vk��iF�tWh	��l�Ҫ���X�V���$.�}���퀾�x�Nr^�̗F�B4�VmѰun�N�1���YD4�>��N�5\�'�ت�Jf́�7<!�M��R/;bn�����u�X�����̬}�f�^,zo��4��媍�fP[��}$~���&>���R���yY�%,������{&/_������c���c1Նk:�˒��<�;�;�OÒp����k9�?i��X�H��=A�y�ju������%�,�5j��y�:�H3�Z�[GgAa.����sQ�v��N��c���:�c���Z��Wh��5�>Ee_��+E��ȴ�m��W��L�S��7C�#���[G۾�x�����VX�y��z�uZh|���ە�|�kn��O~�JC[��7[�]�g��v��ty��,��'��]�Ͻ��9_���6�:�p7�Z�8 ���`j���<A���7]K�Y���"����8�Z2��ެd/76J�#���I6)���l��Oa�g4��+��reI�JNw%�K�|9W^IN����:�8{04�^
�^�׭�朶��x�/n߮�� P#�Q�=�|�p�'94�%�Y6AB�K/���4ڝْ����l�9�@����jU����|ִ�u��t\L9O"�}i��_m�sy�2�N$ȗ��Q�h�,^���LW	��iN���7^s5�#�}�Q�_`w.��NCy˸���n�
��K�h&��)3�}���`C&��Vn�|��'�����,�0��~�ӳ܉���b�+rϴ�EM	�T�M1ΑrI��N�4
}���z���ai���Y���D�Cl�@�xK8ޖx���M�b�Ī3��R��%��Z�<�KVSA!N����%F��Z�23�{u�0��*9�7�i����v�/*Rb�gj+`���������nbƳ/�k�|xf�FP{&e?C�|s"�����H-��b4Ԋ��ME� ��=V���r����{��3���Zf�8���x�M�0�tI�:��f��q���c��5�GN�g��K�^,p�ܖ0:
����jӫL>��]&�����<��5<o��z=W��k��/A�9EW�f��0V^Kse#���4�Wl��#���y_c�@k��W��[���Zn��ӥ��t����a\���[�����s��8=)��ܗu23��z6f��wrd=`�f09U�y�4.��*�s��咃,�c+OE+��Za�RD���k4)�I}*��}:t9��c�"^Lޘ��Et���05��U3�Z��չ�at2\�׊�g;�E^o�=6���Ы[\o�<AYAMFO'[ef�,;������aN���34���"�W�P螄�&8ŭ�Q�����V���d��ޢ�s6೭��K�-:r��Xۑ��S�����ˇ;t�@whY��r����:�M�~Os%���+����F�w�@�tA9�K4���X�1��P �
 le	�b�6�M�>�#�X�L/oo5Gj�;�ۤ�%C%kT�`6��.��Tjޏ��V��J�Сt/l���Y���y�h�n��)�<��`���<x��2Xa�\�v$3ն�f�:M��^v�u3 ��*o/�ƻy�r����ߠ�ʛ��C��[Ct/�u�)�R��0�8�z�V��&H��3��
�)W�4]߻�<}���-ipwf�"|�#5@T��
��R�a�7�ʭ�X�'��DI�X�ƜE�s1\��*{�'H��z0Tv�3�C�e1�6�ia�����=�?P������d�j�Ň�~�f]��F�������S�ɕ��mh+PCiA��B�u���.�,�r���,���Mǖ�X�8��=�z5yP�p,yug�`F�CS�i^�]��+nE��ǝ��\������y��r���DЭT�i���D�W��S�)tH�z�I��ݶw��'J���.nK��pҜ���Y���fۨ�Õ#�h�@AYET��r�=�\f^�۴c׭��9;N[��!��L�X6���u���f�yKt�wٝ՛b�S
�bd�y׹-���5�7����kyg�%�2N*N��XH1n�f�g4��'U���խ<ʸ �o]ԣ�'���s;��gGu�u�1���!*s\���3@�KT�fEW�&1!��(�j»�r�+��B8t)���_�V�ʛ�/���q�T!�����u㑲�.ȩ�Hp>�ʽW�^t�.ԑ�d�ǝ:�aҏ!�.,�R`��4@�鴩�ݜ[����(nN��:l�&N�I�'{���ŋ#tj�5B�.�dUU��*
DH(���R�1U-)TW-(�W5)TA�Q��UCR\�H�2�G5@�Ҋ�REr�m *��j��cL:e�H�~���IJ�F&��IH(a)U�+PUAn�Q5AI��EPV�e���O�����9�܇b
��]6,�Y\m��*��&����=�W�lW�Ã��KAJ>����})R�&��ݹ����!��Ȼlrt��Ց��y�c+*��Z�D��]��V����j^�,�:�=zƶ7E��kng[V:�y:g�z:^ɏ�a�l�ךr�p��[�A���î�X��ȫ���MU���)�p)u�+9�Ph��x/)c���޸�'�9lӢ��gl�ۋ݉��iFf|v�0�'T�����qW�-�9�ةײC��-o�{l;w�t�w�lLq�����r�ǹ�C�$l*xt�n���vyQL@�a�gK�״�0���O՝#�g�f/�Fa�ke*e��Æd�ڌu��RV��{	>�e�*��u��r�̹�pۚ�{��O�Y���:��֝Y�Gp�SVzl���$@�sw�92h�֗�0�~����{v�5�dGk�Y�܋[��S����%?2���gs��5�> F`T����ږ{��=��l��g��<4����owV;]CFx
�F��rɊ=���T�:�(SW���ʏWD����کI!{G8:{;{Eex+�8��y��d��"��Բ�v<�84�.·x�z�z���*�l������Mè�Y���I=�*u�1Qb�x��/�P/L��k�����H�O�e���2�O.�\�/,ܬ�X�~N����)Yj�"�_�+7���Tu�ǃ�<4Ha�A�4}G� 3�k��[qou]�	��#n
b���40Ƕr�*�SB�#Ew��Rݾ&v��ݱ���}x����I;+w���;y��Ԩ�NK�&;8աӋ�*�{:�q���p��ٚ���I���E.��F����Pf97�ZYQ��U�Ԛ���a�:NN���k�톔L'�x���	~.�*<�)6��K��������Nnxs�]��]Ť�.���+(.�����Ө���TK��<�ٵ���5�e'"�o�=0Z��n��#�o�yln�=�{�#��P��)�I�6XE��;<�U�O�0����񓵝:���!F|�n�xQb����3��TNV�u���mq�)���f� �������<�M(7W�E�����}ϸ:�=��"|i�O_�Ԥwv2J��y���4�NG�m��xY����I��V�N���y�U���6�6]x���V*�`�\+�
*�]o:��]��u��x㳹�t�b�#�u�j:�Q���C�yE-����HD�\�ˁ���R�u�n�,Tw��+:�B�ׇ[��Gý�LjV�e{8�O��&滎5���"��)����|Y�|X�<�=ɏ�M�.A������{��\���t֕�����t;@,.��?w0�]J�l����%]{���>l�Gel�k.fa�ܺ�Fo���;������6�fRq�` �:�).�-�{��\���ҽ�S�ͺK-{�,m�"s0S��B�-QQ�Y"�OlC�=���$�����D�£t�(�*�d��m!;l�ŗ��VcNp���q����vl�C�x�)�\���]Q���Cغ.o�Ҕ.˅q���S�K��+2�#���~:�N����z����_�7'���薒�F�"�@��І!�;��U�bb-��w��h�Tp�iX
r@��h��*C�tn�������.������rՐ8���L���̌������C��cs�ES8�ƶ:���\7����V<�X�@�7'o��r���Z>�7��x��Q��WN�l��Z{.	L�@�H���B�krxhv��އ*�����g�M��^d��/�ks.�L2W+o5D�5��vUj8\�6�.����p[�T,��X#��P���='�hdx�ku�d�K+yP��Tb�Vw�,��9m��
ث5p@x*'���������9��'cݎ��نG�_�z�.��ȵ;�ܻ8�5�6�:�(��-�wW���a�kZ�g�>���?W�>�)�UE"��B@�!m��C��N�@�!�1D���3A�!F����}@�ê����ΌxO	Ԩ20���
1RI	#?��1yټ�E�ꂠ}$M�+�D7�H�jS��P�*J�P�~�А!"�]�:���_wu�k���>��|��(D��2d?N.~��^
!������._��MN�Zܛ�a@6X|�2��~�B���=���/�~2v��$I6��!C���a$!��%�������A�C�����O�C�������\?����>�����C���ο����$D@����$�O�����ܰ�k���2A��(�i!_��!U�ԑ������� ������4	�w�I��	�p��=g�V�m�D�H�1��?I�r�@�R��Уl
����^l��������?l$BY4B*�G�h?(hL���c��?y�­���T�2`s�}d3��@?��O��� ?�����������2�!C?�*Fx�pI����������?��
?ڟ`k���!A���~��o�����`~1rO�L���~��8���/�$�激~��?�6~��	���2 ���o�"���p�d8"��p~!C*�1�$�� �Xd$B��'������'��Z!�:2P}0I��	�0���� ��4}nB��@~�D$�,E!��	���	!T2T�&�I��!�2?�Oa��i% ���	�H\�Z�?t����f��L������$B��}��~��!�d>�!8�����I"l����S��B�>����C���>��a>����'���#�"?i���_��~l?�?�	��C��}!�c���($By�Ϸ?��_�/�!TQ ���Hr�	�I�����Y�p��?��>���^'�C�>�%�R����7�8!�.	����XK��������>�h6~r��>���9p�:x>�?\~���$B�~?IC��?��ֿda�?v����B}�{
�o��}�2C
�L���?B B��2O�.@,���{�'����;�����!C������lh��j��D�g1�Q'#;��p?m�MH}`�B�	�E���B|�f����H�
|�`