BZh91AY&SY���6߀py����߰����aO�    uB�    @  ^�M  Pn>�����woM��Z׏lֵZh�2�a4�wL#���-U���  ��ö}  � ����f� �             �   ��� t (4���3����:�������^��O{�C��j��L���{��读�����v�ځ{��>�}�[=ۚ���s��Vǭ>��z
9��jޖ�{��Zn������՗��kG���C�` � ������t��^���ݝ��7lGr򧇡l͖ǡ��h)��yyv7��<=v��ׁOW@ �/J�w���
{��h�s�-�G/;:4��r:�vE�=�́��˳�gn��l/>���( ��k�{f���v��H�7fn�+����l�:�-�%wj�����Z������z��$��jz{�nݗM�W;u�����x:�gI9�!6�^ �b��G`   ���'�\r�Y.��N���ǝ'�����vݳ`7:������ ��oy{���=z��k��wn��u�tk݇\n�e�붺�W�m
�6   @�v�cn�����=/{�y�7]�i��wPf�\�f�pP�K���]*˼���j[M��e�=�W��n�l�ܶkݻ۷�@�     �@           �              	T��UJJPz�H�� �4   ��BIR��`&  ��L �ڈ��R�� 	�L  5I��4` L�   4�� �B #B`B�Q���x@UOP�J�!�L��` #0���~��/� \l+�C��	�����pd��* t̞!C?��� J�����/�V *��0�U����������G����I��P�"�����H.�@����*	RI?��DT �T�
vђ
*�&�ˠAw���G�3����N3�JO�7'�V�^'�b��5?Q��Z���ݐ�ܢ���N}��N�L�jjtΕ�w�;�{O&p�r���O't���]��9�<�LL�d�E�
Jh�'��+"T�'�NԜ#d�"%��3���%�����俒��g�u(�h�w&Y��~��d�gϤ����?#"{ŞD��f��8D�%y�Bh���^K����Ӥ:���],zO�{ʭ:VĢ?DѨ���""{�N	��%p�ؐD���L��1��F�W����cq̑�'?��'VW�1�'<x{�_#�
-�&�DGޕ�?"_�R#���+�2�pKy)�%"/%x��#��;��,��͕�	�t�?DN7)ȍ������H��WDL~��nV����r"V\�	�ґ8���e��@�nJD����_���_?,��[�D�r�5�,o���ԤKy)��nV��������C��^:q��N,����E|�R%�)����~�w��'���eY>�ݒt�Ii��	�e&ݕC�;R��[���������J��|��x{��1���:���858\���~���{:ʭ8_�Ht�C�A�ʯ��WJ%�_Po��X�rR,���x�DGvV��y5&�Q��sD�<��������}U�k�^�=�T#��:`�U&�4� ����O"7<vL)�f	xʬj��� �/�G*�4ˈ����͐vC�h��LɚOh����;SL�}��;�ώ���'æC�!�~�~�w�R���rVt�d�=���Y^����*�ظN�{�����~�w���p�<#���ʮ��}+�J����,�[*�j]I�|�ٝ�����&N��.N�)��e,��egfW%T���'�8�Ry��l�1j�Ι�ܓ�URN��{�_v���o��f�Ȧ�I����z���9>�12�����%�W��t�ɉ������'K���uI��ɇK�N�'�LxIY�I�:��#��I�(����I&q&麓�>%��&��|Q����~���v�y:&�&�!7�3�I���F�7�Ͻ�K�|��D�:���12�OY�8U\�e<�N|�O&9&���T��%��aH&2LHc$��2T=Bz�=g|��;���m�a4�����>���>FzO�l�V��C�!�b��8Qd���X�i2���C�G�i1%���D~�DԆ����?Q�O'�2P��D�"o�"iN����-9�	&���|��a�s�jxN�'�æX�T,�	BG�&��0p����i�t����H��H�x|A;�+4�����~D�H��DM����>JD�$KBLIMI���'��DI~"'QD�	�*�"R"[��Qq"'��O?xN����(v4��L�ǐ���DN�	Z�L)��	��NRDOy"$Ԟ4O:O,Ǥ���eZL��|q�ae}h�<�":x���M-"`�B^�'�âbx��&ԟY�'KBh�9�	�I���"xL�Dw	��}oI~�y��t�}��<�<�0��I��'�w�!H��D��Y4IC�N��:r��MjJ(J'��	�Oq'�߰|Qo�OԚQ�0M�&���ɤ��Gr�{bx��x�rx�G"e����x�ق{Dʉ�p�C(�C؏��a�0K�ƧO��;<q�Mԣ�o�/����&�?p��N'��P��%H>!�g�:#Q7g��s�#U8]]Dk�N}ü:�LK�K�����ԯ"8���~�%��x�<#��O�W�:���,ߨ¤���������^QT�*J�<�=��Y1y��g��+�֧��jt���S��#����]+�?{*#�_d,�%5;;8�e���ҸWcuQ2�zO�DG"t�ϨO�D|H��:[>�_d����U���TDY�Kg�FUDNX��",��S䡕Q�j"2'�ژA��n�|�+���D�'���%'�E$��eTD���DN-Jѩ�ϓ�,���L��O���H�}⬑�"&��t�����"�DӋR���� ��v�R�gjxF��'-�D>Dn�P��R�cSD�� �|�ʩ�G����">doja�����"�DӋR���� ������P��DM����jQO�;���N��ͨ��5:A����,�p�r�>���ډ�jx��(�R���S���5���N���*�{8w���TGg��$�
=D�C*�98g¤Y�:i�t�x�5u ��xw**V������Zh����)"#�d�`��T����:��d �$᧥�Wǎ���t��<t�G�ÇOQ'���}�b�:�];ŝ�X֋�4�I'G����Gfiږ2i��0~��ͨ�DL��a�ғ�9ڔs�	Y������62]M2�ʇ�rWNr&�5�T�E��qf�SD�|����î3�[;�gylyl~�;�7l��c3��v������>�[��G��ԾƻQ����Su����s'��7t�Gި�j/�V��l������G��Ԯ�]G{Qɞje5=MOT�m57Z�ʋ1�ܩS�*v�D�':����0����x&o�N����&=Rӵ9�ۉ��fD����g�YU_{�'�G����6w�'ܹ��S�]�`�}��G'�'�VD�̓�iʉ�9���ܩ䲭�����ʙ2����2o>�̭�ƜZ4�H���}܍C֪�ri�56��R�ҫ��*{�/v���l��g��ԫ����T�|�=���;��M����&���fV㾲}�5�i'	����
����*=��#\�� ��ڝ=��I�%���!�%iὕ��2�X�D�$G��,����"uex��tn�|�Ģߢh�D}�_#�%��Z�DL�C�T�	o%"a�e'�W"$rR'q���?"9��CD��D~������J~��ԤKy)��nV�������yr�'JD��O}�x���{+�[��=��,��F�W��+���:ܤMy+K�}�5)�JD��D[��N�=�_?;)0��]��"qe'�[+���KrR'�����4漏O���ʲ}�$�L�D��uڬ�eQ�h�)vV����au0��8<�9�>����'�ƫ�ǎ�����F��Gg�9�7ݕd���!�C�чk�.�ev�խU�i��0{8'��4u����Zwe���K��OH<���Gb?a�:5:&rc��=�J���K$L�X'Gd�u�~��A�Ӳ{�N�=�4�eW��0�A1 �M���n,�}�2��vC�#�}3&웑YK2�r��
���>9�v	�&A9���B��n1��{��u�V{�W����*��T�Qr�ʧ�^:�;+����Ӆ�ʯ\�nU=��ҫ�'���+ײ�d�9M�����ϙ;��rK���C�;e�]�D�N}T"{�h�L3�'n	߽��ù�OGa���H��~&o�����h����?��8O�T?���M�V�P/����aĥ�o�S!P&������d�,e3rMNMML�.�YՅ[���UM5q?�����-_$���|?q�5�E����)��5a��Mu|O��|��(���j�U^Y����˫���z�x���rx�������Ԗ��o��MjԔ_-]Yt�pJ.*��qDב��VB�xD�_(���>�����^}^Q5���&��%Ē\]O�Q5U�}>>�l�V����k3WSMuuq%UZ��E�M7��QEWWQ�UES^]Mq%�*���uj�S����l�G����̹r�%IE��}<����w��ά�����:�������x�\�[�ܺ�W����}��m��]�l��s�NJ���5$ĝ���3|Ԛ�^�wwWU|�
�u|���ڼ�/�Ww�2�MG�q$��1x�����73r�e��$��ܯ�4ndc9;.I����[�_��'s�s#c�{��k%M�j2�FU���-[�噫���_/-+ի=���'���'�ɳ��d���=۶UmՍfw�Τ�]Z��K����W���|��/�D�Z��/�g��,�q�\QE��*����������8��.,�T9537*\�����w��r?�3s�����%V�7�y'�NL�ܫ��j��ݝ�ʿ.��:�Uyq%������x�\�]^�U�[|�U꯷��S_,�7��$��5���T��ͷ:����'�r|�K"̋WU_(�EW��<���I&�z=�ޞ�j��,�d�;���#9.|Ͼ����/��܌�ª�23���g�L����l��V�62�=wu�ϳ�RU%�ĔUsF�<*�%�έZ���z����ur��\�V�g*�^...�WvcF.8��������{F�&L�rٳd�= ��z}S�;��d����Tj�KUIuE�������y��\�^/v�m_/w��Uʺ�[�]M5��//�Z��3ɩ�߷�.}Ƿ���|�$ْ�2rz��쭿FI��rEՑ`�[=<���^UyycF?��$��N�!��z2/c��Q���D��e8����\}�fJnb=�P�R����z>���ܔ���Rv<�I�FC%-�}[�;�����U���j̚SK���9�Yh�G^��6�2�p��Q]��L���u+�������V:�hrj̘�F�O"�͟X}��Uochѿ���>���T�jf;�����'�V6J	.#�����3�����G�$dYVU�f/q59E�5�+�}������fz��=�%z$evUo�4nŕ]�)1ř+L.���J�
̸�W����!�^�,3cލd��J75��r����J��#>E�D��U0YZSU1Q&�|''eÒ��+h��}c�^`�19����e����{1ՙ��g8<�Mg�2����VDTYVeѦ1#��6�"xsJIG��y��T�Өf(��qѢ|<F��z4\�*���D>S�5Y����FE�yd�sΊ����q���\u�Y)$w���FE���+
���y�Yq��&� ��SM@�u�C9��yv���G�sCd啘n�c�+��sGQ��o�{�G{+��sCاY)֊�dQz�(pd���:�%2�+���ԭ���ddnv�����}͙�NGs�[�V��*��jr���G#����#�#�2M^#�|+Sq�̸�r>�Wұ7�y�J�W5NǓ�VqU�^Co�yd�D����>�}\Y����F�wޘ�ĕ�?�Ď��X�z:��eÄ�J�7�9N�NG�VW*���ˮ�uo��{��{���Z�y�ؓYի%�/{��������ί~R����)埔ė�*���7�������5$s.;�3ɢ�7MǓ~+o}E����J�Gq̸�f9����r�V�c�r	��'������=�L�~͹�G�Q5uL��CN�a�Y�-/���o�"�=^�jY�ucIf����ׇ�F�Ԗj�TX�YV��ɟ*���ի<�,�3��'�Vt��w��ތjv55LǓ�*���]�1�+��}��Դm�g�-Y�՚��TX�߇���Τ��z6�ϗtz��%���iU�����.��5q*6�X�Y����8���ş,�q$�}s�ժ����s^*��ۜ�Z��j-xs��VywG�,ԖT�U�:���=IdG�y�mdF��E�J�ʬK�NUj�j�˫}��r���u��}��jS>�<�}��\�L�jS'ͳ5f��`ugYYYtm^��v��s5M�>+��iG3����s[��{s�j�j���O������n[ݹ옶���LCDs�[+��e�Q�w�\)�1ڨ��j;���O�X+VqgVq��y��Y`����d�K>Y:6��n�u`5���\�:�Vug`�������YŝY5�����Y�E�",�u�c՜Y��Պ�Cc��x�ϩ+U�阎�#���:����j&��G0�S�c4�5��L���X�dfzV�x��MG�u�u���x:���,��y&J�����:f�(�0�+1�K��!Q�Q��*ʱQ�����Y�k8�VU�g�����Q�=G$�U�Ñ�TdqG��b;�P���Օ��9������d+q�99z�1��q�,d����:f�>�0>�?J���*�q��E\�4N��G���Fw�|?,�l����*,y<4����Nl�GP�.8�H�B���Q�
�J��G��Ȏ��oH���r��6��,
���t{1.���ϸ<՚���f�?�Nc��,�#�R��5b�ş���qj���bg	qfT\�1�7�}l�G�+�:NGq���3�hʛFhu+u���ɐ4Np��9E\y���[�7��6�`�[���0�J�sP]z2Ʒ*D7³�R;�]��Z�cP,�\�kCr�+�ذ�#ޗ�Y��]��G���5EH�9�y��Y�q���=�#�v27�`���9Ҳ��{+�ݕ�+�q�y�qƣ��s�G0�*:��µL�c��;�㈕r�棈�k�+Xy��en�;���;�c����#Q�s��!���r��nW4:G��WҔ���L���j7C���y�e�ʩQ���=ٮa��s�<�Ϯ�F��eJ�Z���>�V%��'�>��UVu��W�W^^]]Y�k��W�Uj����V�g��\��^�W��-�ϗ*�y��57+�T=�1���+���������~~_}��!�ͧ�������b�X/}��g|�,���5�����f��^�ϋ�nY]�םeO3j��ns-���d��;�תr�6�.�H{;�gs{��W�#���_(���%c�.���y�z��}�Ԙ���{M�9�94��y��ۧ�����{�+i�7�.w[c��,��U}󝂢���_>s���O/(�N{���g�M��r=�|�^q��=��x��W7y��7z�|Z8vq�zu�����Ƹs;���f�W���}Ӌ��b����<�Qɩ&{�Sj��V�t�G��vogd�'�ގ�.���5ȓڷqm_n�~����Ⱦ��97�V/3ȴ��ZY�8�W�ܑ���~���9�M�l����s��{��=�ז��.k��mw;��7���d^���!�����WNs����q_{�^e�;����|p�Nou��~\����9ޮwD������5]���G"}]9�uÏ�[��w�{�����}�7�IOn�}:�]�Nxm�{�w�9��V�œ��>�s�Jk/{o%�'�ԩ�j����N�]�s����{_c���|���|�u:��~뼞���]��s�}�}�6s�>����oQQ�8���|q���������d9_����	/�/h���M~�� �����5��j3����;�.����jʂf�8��Xs�X露�k@TP����
�������� �A�5r	"��(|@��=B�9��w�D�i@̸H�"�\�r*T_@�(�n�J�e��"&`̤�S1.
HLT�!pK��#QNʋ�!P\_/$�����R�E�oxB�"�ʪ�Ȥ�� rQ��hԨf)� �A��ꔺ��;�MQ�*%]�6Bx����� k�&�ȉ���D4<���@Π�����7��5 ud���H����h�"h5vl,�xqdXqa���2HT���.QO�nJ��\��"]�f���[���t@ۨ*K�!�UYP'fae�!�VdC�%��,���V@�h�@£UFbvUfvK�k3$�S*0���͌H3x�:���v�=>��g8���f�v������Dnj<� ���<�'yj����Z���^ =�q�v��M��wF�M�w���Hg�/7\�����حL���ϓ�n.��78zW+����A�WK@�i�@�#A(�L�
�&"�"b NR��>�d����"��M�̐�^n�@�C��
]�Բb��p�+D�D�,��1�W������JP;	s��{��rA�1i�Q5�Fj���3�\K"��b5J�+P�9D7s�Z�b�$�$s�y7��N�Y��;1���?��u��QAA|���x(?��p}�_�ݟ����?A����������a"���HBT��?����������4���U]b����Uz�UU�UW�ڭ���^*�U�U򴪮"���UU�UUu�j�\z�UWQUW�^*�Ux��U��U^��ZUW*��*�\�ڭ�ڪ���UUu��������U\\�|IO�YW�rQ��qV���|��e1h
�Y�VS:�8�&�NY�lQ�k�9b��Yՙ\�&�[kMX)Ճ�n���U`������TUUU�������j��[U_,UQV*�Ux����U�^*�U�U򭪯��UqU�j�努Ө���mU_+j��[V�\]�W��UmU|�UUb��s��U\ZUUTUUTUUTUU_�d�������KlQ&��+m=[g&�5@�ճqck!X��D̦���M����Qdw�X�w��}�k�UqV�Wʶ��UW�ڪ�VեUqUqiUU�y[UťU|���Ux��U��W�UV*�Ux�j�努�UUU�OV�UȪ��J��^+J��*���Ҫ��UU�[U_,UUՊ��@��H"F2 �${�.f��Vx���څ
lH���©Y�O�I>���s9����U�U򶪯��UUEUWX��U��U]EUUEUUEUWX���Yj��Ҫ�VեUqUqiU_+j���X���UV*�Uz���mUqiU�Պ���UUU��U�mU|��UϏ���I>��>Jl������r�q��c����3���"�H������ �������5`�� ܶՌ�倠B�nsuJ\Z��ԨH� H�H�#qC�~c�~_�b��#��_����ƿ��)�A�Q���~��8�t��C���"X��'H ��"'DL4D�0�8P�!B �"Q,K,D��"t艂`�a�h�`��h�P�&����xN�DJ8""&�����K�%	�P��<'��,��'ȐDD���B�B"tD�h��'D���P�%�A<2DK�pH'��p�4�M4O��DJ�&�"h�tN�(O2�<m�"�f��f߱�_3���:���T���brA��	H�j,lj4�IV�,n�j�v�-�n�n;T$��4X�ZϩEEfO���b�yaũ4���
8��&WZv1�b����"�"�i$��[���p�,X��rR��t�Q��(�	Ċ6QK����"QLv�8Z��c(��YY`��	1%��cT�*E�%R��r!JG%���Ujf5
���F�i:6"2��LB�[U��v8�aQY ��VA�����#($:�B-TCti1������:�pvA�$��%V�ۉ��%v��QR�H�
JT���W��N��i�$꘥�72�8���%��TmYdX���kɪ�Ѭ�Gl�F"A�̩�ɎKU��Q5�K]����"��m<�
����\L�QKKb(��jQ�K�O��X�z�cVT��GS���vX�)��qTXӰtJ���e�4�-���H�uE�	[l����S��4�Rk��c��"��ǒ	H�	�d ���Q.�e�Zy�7i�=/��׵��)h�L�����*�LE�*Q�R�h��D��$m�Arƨ�U���!�8�����d��O-HX�Hq�;��j�-ɈlD�Xĕő��
�������f�N���I���7�1!�-v�,ClU,W-&:��B*%���X�ۨ�j;V���5Eb�-��أQec��"U��(�i~e�j�ڄ��q��F��x���؋��k�o+#C��K9����V:������(₅�P����,���c�m�b�cJH:I!-e-����BB������P��% �1L��tlX�H��d�eDB��q%���/%�M)
�	�R��we��TP���D�KJ���T	+^(X���"\N��N��㐷�z!�M��R���:Ek�B�x�&R�mD뢗V��L�����Y���ǎ7-��V"�Dd�u,p��FŖ�x�Dw��Tj�\j�Ғ�y~�U�,�	Q8'J��Y���Y.(�F�J�"%Ȅ*&Q��R&�ƭ!mx��u�
QR4$�I ��U���N�T����RS-���.7H�
����%HE$�+����Ȑ\C"쁢�E��G1��m��)$�af%*�%%V��E��,k$��<� �tTC�����tYD�ѡcrJ����ib*
����U���A*P�o���)s.J@QԬ���H�KD��H8쟮�F��
c9
쮊��--(�eI�$��E��6�E�c�a(� �1
 �~�T֡�$+J,�IĮQ�
R�Y��pdF���%.Q+v���),��V�q�Y��F\N$B�e����%Vc����$CW*ō�!RԥD�P������"���$T!!����.G���]�ȫyP�[��.)V�x6���!��GQ<���+ ������!*D�t��\�@�+�Ҳ"!!�$r2Rb"B�� �E�J1
�FdxR��U���CH��iZڶ��1�$ć
�T��
N:n����X�J5
����t�����GA�!\�%$(2��D��	��pn�:�lL�QEEid�x��"VH��P�fF6$�,JR����!1����q��r#.**!���Ui ��(&(ةV"�+�*;,#�7�L����U�+���6�kd��iˑ[��QJۅq0�%�������i�r.q:"U+�'Q%+(%Ui�(��eUID1���	�D�y����x��%Z�;#"�6�%�eq�'�����IHG�N�d)bV�H�m��̑Gk�6�M51T9���ƚjZ蔌R��+,j��r�Q[T�բJ�F*2*�F�q�\r��¥��)
WI2�1�Q�XV+cn�(�i�"�1�D�S,�:���*��֭%���ҟը ��G���#C؅\���
��bi�#I�$�j���J�U�ą+\�-Q��T[h�I���Ƃ�"j���J�*�$�����҉QAK]C�&�IѨ��R�T"R��ccR+VB��A�i1�޶���ĚRLC���L�Z�J�`�YQ��`�QWn1��H�v��e^Lr$��DN�X�I��[Upeuc��r�Ԝ��J!6�y��R��"V��UJ��$r����VT7hșH�+JGJX�P���1Il,��[]��N��F8&�Vأ��Vۺl��G���+�"T��9S�1���W%�Im!F+��e�)!*JԪ�֪�QV)D��cr�UFF$�n�Un(�
+m+���RG��k-I)KQ�R�,��$&%+M�*�$b�G[i��G��X�J�:�!":K-�"T��cX�J�y[��%&8����V��M�W\uՔ��btMڒdtR	��M:�B�9[v��Z��)Z����)j���$�lR6ۨ��3�s�CTIH��܎�ڷ=m�2Cv��bBV�Ze�&��N�2֕J�T�M��VK]�K\�m[mO�c��+5G��"#��R(����u$H;�+�	a	\K�Z)�i2����)b�TY1$մ�7J"�!	J�X�%m�)E%UT��RI��
%j��Um��I�Z��p�M�#�(�QAX�i�$�1Z�D� �dJbV:���+H�J�,n�X�"�2є��v���Z�FۑEd�T�Iܲ9-�Fy�ږ�ҍ411Kch�	)l�IJ2�Ș��EJ� �JMUU���"�VUE(�m�8B
�U]�	��bU�$뵦�Ig��:>6��9�����UU�Uy�s��>��U��Uu^s�������iUb�U]EW��8�����V�W�,UU�Uy�s�����}�~)H�0�ʔ�o<�2��0���8C����Ib^�mR5Er��"�LV4G��+�YP��[��A\b���䒼.ETp��bn�$hM!
�J���T��5.!5X�k����Tc���y���4��'q��b��U%bu;d�R'��jCI�LyPյ�����YFK+Ea Ć�% ���!V+�"1�	11�ȕJ�u�jD����ҔX��:�V����5DF�@J"+�E�e2�� Վ�&c�G"b^)E���q�46��*Jc�p��
%m*b�N$��L�KAȲ)�cl��2 �y��),w"VD�KcN���w�i
K>1��5{H6D5j�TJ���8ꊦ�V&Д�)jj(TT�*r*�(�dmBH["�Qj[\�q�6�uэ6��%�++*�2�
�Yl��q��H�:%bj�$��V�1�W,�"��\+�;l����+UM��mi:�c%���m6�B�G��C&EA� ����4�q�ɓȚr��*ʫą8�mn�E+��椒P�:��k�)o����'ox�~���8n��ƛ�ލ��s�<��9xz	�;����è����[�iwDL]9�^�I��Ȓ:�ĕ{�o6U[�#rh��d�W��}��8w���S�8j��Jm�J�G�#�!xr~Z4�}L��aP��zh��'�ʢ���p'g��eԱ[�����u�܄$,�o����W����9�#�c�9a�������!GfI!���!�<Z'JB�ks!E��,��]j�+I�OvsH�>�:�5�>��{$��p�!��66ܙ�����x�abpO��DӢ`Ϗӄ��y�R�2��$�6�0�Ti�᳀[�V��YC��4n��5+a�6t-�ߤѳ|&�t��;���pe��2��L9�2�V{4g�qQ�d�O^=}�&�޷�5��N����vܜi�M��l0L=s�Kr�kI��L�n��2�6��:�6�<��l5k[7����eMa��_0ԒI�z�22�Ԇ��9�c�KE��bX$.f$~Ha�k&�x9ll�`X��,�w�Jd9[!&<v�BE�d�f��zNg������Z3ZDd���4>2
{����7�[z3L��d�&C1$�X̸�c�BY׺�їQ�g��h�*I��ăJE�˛�gN���O�p��"��4���,���"h�'� �i�,��U$ܾSo3W�^I$�2���e�J�&���y$ 0��"Nv���bn��k�S5�S��Cc.NTv��I6X�ՂB3�SL�#��q�"�<���3�L9����D����
[}��ޠo#��X�<P��7s�T��6A���^L��c$3&Im�]e��q�]So<�:�n#κ�6í.ַ&XZ�뱳8p�-8R��2�p�*\����Kx����V)ĒI%9�"}�g����_=�'(�p���ח�=0{�M��/�|���&Am��^�����{r��t�����{�Zs��ո=�+�㞇Q�Haya}��	X{�����p־��Eܝ�M��35ל�0�Z޹�U3�\�;�{��ͨ��&M�L<Tw���Ew�-���xr��}���I+���]��u,��E����N�;���V+c�"F&ޖ"e��9q�6{!�:m4��z8A��:|ч�gQ=Ƀ���3u	>�0�Gm�A<�!��87���%x1��D)�!����nސck�)��Gx@�I4�te�TB�-D��^wd�ș4ё�鞻����t�ag�?0�'�D�4O#�Ǆt�o��O"6�A���7>I$���c��gp�	�FIe����:��;;��m
�~z�k�y��b<6�V��̒")�U�2}8P?�8,����=��kn�!�I~�8'�%/9s����ĩ�9�%��4�ӢT�B�}��/�p���ٟd:0�RPu�'EJd3��t��΄0�O%���"h�|p菏ӄ��KI�Ɏ��Tbw� �K4;ąey9*T((hR�ޟ��(8g�IP�BBD����EtT6�� 6��Q�6��d)�9�=��R�{��윥��y9�����Ӯ���9�R��;!'Lty�=R���^�o1�1��!!��m�!�E��e���SS-��KCn��`�f0OǄD�4OA4�x��珹[K4�*��Ӌ�S���ʕ�LrI$�2���@���O*����E��?B��H��;���[��mٿ�6ǉ�%�Z�����7X�a�:n[�E�]od�480�p8W	��D����[&Y	�*@�=r94;:I~��ʻ6d}��2�AOL4l��K84�FCc{lI1�ml�]���.��o<MD�4�x�9��v�����ih��v���|Cbh�ۘ.��m�'ŉ���X�j��I$�=�'_z}�N�|���7�Z�w뺾ӳ�xʾ��K��6���w�{��ǺC���ě�>=�,��vK2>������2�s��{���x��oa:Bty��q�_��U�j���{���B��M���ju>#���C���w�{��Ҏ���o!�q�ߊô�o��ڴ�E)ln���a��z<���!�DÖo̒L��e��BI��}��89�}n]�vI�!�3�gx_�H@�s{���p�����8U/4�7�S�=�둶���S����tA�e�n��x��\L�~���f���w�9�cg��Ox#z��3�/E�מ0�w=����&��!�<t�,N"xDMD�4�x��L�Q���AJ�I"��np;�������B|c;�	~��{�*R��n��f3/ӷ�n�*A˓��d0;�UJ�)�ҺL�$&c��d�.���`��)��grtK��]*ٶ��7�4uƦ�?gӉ,���zcŋ�R�#�ph�l�G�v��sΥ�TZ�LkX�	:u��H�Z��u��M#IH�iW�(�QW��0�%"�y���lbR�K�Sү)vԽ'Uy�JJyu;y6����bJ^*��IyR�G��B}#��B��t���N�~!��S�%��]��<�#ϗyG��˩�ݤ���ԞJyu'��_�^��/��qM1t����/M������S��:�Ra2�)zFR��RmzJE2����җ�'$��&Su|���J]zOfK�K�S��u))K��JJR�R����U�ʗ��uK�)4�	����g�Ic�Y<X�<[���K��ړ�'�-�-��KRe�E%�M�Z)-���Ǥ�8q�8_O
N��<^)u%0�*�ڗ��%'���]N�FԾѤĔ�U墒%I"6��)�]IRZ6�#�0�`K�=��?e�s�~�x�7���'~����Ϛjܾ��w~���޵
�ɩ}���[�^��Xx�95dQߓޣg*od����/_���yL��w��W,�s�ۛ^�y�1pz��}}��v�跞������<t򏼗���"2$GW����P�tZ^��yv�N\��N="�5��u��V������OL�����p���������~wo�����zJ�{�E�驝�F7�k6ۖ��Ny���!ý�j}?�d_�p�	:�߻��E��{����������Uqn���}�������W*��U^����cǪ�Z��{�����UUꪪ��=�{�=B����{��oު�UUUr�[������i4�K4����4M�"CK0���,�Fr���`�b2�?�i����-��at��1m�Y�0����ч[��H0�4��(�*S}�cp1,������%���̉�Ia����c�� t`��E:��L
2��L3��xx��L�'�SV��u�oX�p�M/O���a<�7�K���L �
9Yr8E�Z;,�,aŮ6A/aC�e��::�Mj���`yV8��gTG5r��0�ō��A�F>:Y�`Z���l��H�}H��R����6�7hy"يK[$��],����ke�Ѧ�u��R�6�:㭼�)��C4���X�-�/j��S_ ����}�m����WU�UB���i�B��a�l��TY��~�a�~?���1?��%r�J�N��w���ZX�Z�,*��4�����8�73$����D�]n\`���Gݽ�ioC�p���+!�:`i(�u�k�8�B�1C�����W@H\n��#rJ@�A�`S;��Ui�����	�˶��4�0"Q�W�
�`v@��6��(�vy�Ŵ1x�iLN�"X�^�գ�8�ֆ�F�a�2'��D�0�!��(�� Ow�b!Г�HA1bg���,geN4�ؐ]\ob�"���EEEA w9����}��W K8o^���������W7�d^�ϝ��ÚY;�=��>.���ӟo�ᷧˇJA���(�v4}�(����3�$y��RTL����c��g��o�;��$9��s����*���-�W����61�����z��ޥM��C�}�|�~�ϔ�su:r��kr�djJ��<�
O��G�	�:bP�tb�& �d���ԄÅz?4�kH&��6Kv,�q#f�,mZ-M�{�>��DJ���{��3sH�adB���<h��|P:����h"�狼L�P��!(����� gUR�:��"��
��>h�����t��tϟ���B�&�P��D.f	a�,�Iu�F�bZ���y/c(�'vJ lb8Q��HA1�!���<�tl���h��~?��D�4L0Hi�J4Á\�U��9k��*i����`Ȩ}�J�h:;�!B�4B!�0K>����I� g37��dE��P�[�f֋g���F���H��k�:��S;���L���I����Cĵ�!-.e�P�|40�b�A(��&��+H!�F�&�Mέ-��eh�d����!Ν0�[¬����	��ñٽ��5&��х�=pT�ʇ⠜���z
����f��>�P� t`��|�ۨ���|�zӓ[	�@�����3G�AA��h,ݛ��	����0ha�)�(��!%[+r�Ţ�d��R�g�x�h��m�)�>m�u�q��8xN;ݬ\�h�1�ѐԭ�hH���������^L��Ԓ��o�}��|'|�h��֋\��EE��Kf%��3�
����	Ԃ �A2�*�]rl�[�����ݛ떃�[��A!���T.#%06�K"�E�E�h9�11�f#gx���8g��ԥ�X�Ê*�T�6S�AOH�$0s��=��Tr�P�P������֋b���q��Z{#�m�K�������`��v�l^��xF���W�RKd3p���9�`ҽ`n��"D��l�y��f&4ݎT\��QVx`h"��t��,O���?��"h����먧\]�H�%����<�K�I�.Q#R�d����QQP�#�o��B�;�����J��M |A4�pB�ҰrН�{!
�R��%</P�aQ	�/��'4��Ҕ���Y��a��
`h*+!��Cp
 $KhH������&m{D��c�a�Y�!������IaLL$�Za��	щ~%
h Ra����(���4��ʳ�3;�5��*���7F0�A6D���.�F	�H���ٞ��T_��BjK �l��DY�-r��lA���O0����ͼ�μ��8�:�)�	������˗�w�h���VD�ñ'�Q<�'s���q���6��8��G��_�j��G&����%��p��9%�o9��u~<�w�?x�_)f��xã��o\��Ǿ���;��p�"�����g�sg4�Ɠϑt���e�C��v<�W:�'wl�Mz�����sw���I�;���=<Lrս�L��2{��'��z!+����&�d6����|�&țz n�P	���c9(-"�gD�5R��0h�a��2�,>�,���r� ���ϒIkn.Ɍ����,�bA��a�a͊��6��БV��j�o���ϥ)b����	�ٿ �1�B��$�M��d"}��$![)��4i.ʍi�C���66�!Ty!��0�$6�C�B��M0�>da��u����u��~�Ht��<t��)Ͼ�l�f�$���6U˼E���r\�̜(�=�]eCD4R��44%J ?8`Q��y�|I0�[�2]�q�a��>m�h��`��H~4��s޻�+�^���.[2voDO�TTTj��8z46�	��y�����]]��W�ه�FB`X������X��!y�4&݆rFA�M·1�!�1��N� ���gG-�a���p3. �p�n	;�y�C5 �u�#���ZFP����@��ǅl?_�:�Y�m��&�fi�޴cK(��:����0P,,�K�q�2��В���O�,�z����2B��y��Ƃ�b�A�u�l�vT0�� �nǃ�\N��ĳ�?�����"&$8p��!��Z}�$.����W2�%�.55�&"����<�۹��-�퓹�����Tdː6�+'��?8�:�G�OÊrbpG'�_tx}�/��m.Nɑ˃�`B��N0%7�9�\K"��,�d
Qd1�({}�UĽM�8=|���!����Ɔp}���У^
r]-=67l�C�& �۵�d\��s���--{f�u=~hl�PP��Q����>���}_V�_(�e@�k�H���C��l:�ht��&�
ltoıeb-OZ�5kE�[FG��K4�?��"h��`��Ha�賧�A���qW�4�W����i��¡E�����>F��������@����Ya��@����p���DPsH��~r���x�s��D	�σ�2�≔ٛ˱��B96ۦߏ���e����T4hz8rG�ކ���t�Jt�I(v�9$$4��mBs��H�ȑ�kuf�V�u��d˟������X�F�
�um�R@����wci�Ceō!�\���,���Z-� �p�8���r��&\O͢ڳ��n��[����/��?��O�J�'�W���l���<'���ǧ�������\����X��:Ȥ�RS˩��R�F����Dw��U�R�-�K�'i�q�&QL�l����R4�ԍ�\��y��R�i�>]�|��<��ԧ�Ry)<�����u8�R�)))�1IM�IIH��<|)<D���������?���'�[�W�'�.�2ژ])9%/�)}I�L�S)k�$R�Ja�3III�/Jy�F^�D�/I�/IM�J^�Ȥҗ�씿�IƗ̒����_	H�R�0�RK��K���ړ�'J[����R)�R])JM�In)uԻ��:Ng��x'O����L+�RmK�Sג��IO.�mK�-��RD�*�J���%����/I��E��KF/1�s�_���c4ظs����{���y��ͺ�N�Aە����}��WY��vOoi�W;[���rBb�P�[q�Xv�����RO<=G~�	!Hee�g~�9�6��tx×�BfY�\#5����4'T�}��=��4�w���M2�z��W(P�_�g9.|.�S�RS�lr����|O�����d� �<r��.m��
��G'+�0���u�/�2aw�^����x���}��}��N�NM�jYkի_���O���94�l��_���?.�k7����w��~yWӴU9���;��ZM6Ԧ�"W_�����1��������{��v��ڬ��[^�1ϻ��~���UUUr�U�b��}�����ߺ�j��~���߿]��O�ww����UmU}������w��ۻ���������Y���ݻ�� І�CM,��4Ҕڞyמy�G]G�25�&��G>-�Z���*��%��H�y�hN���e��ˌtI��e,Vd�T�mKZU7Q�ڎ�����m6Z����K"jv��9D��أ�u!�B"WDt�d�;��X(���+QV��E6;�b�i�r�c�oTEQF���TȆ���$)����I�-(�H:ݵD$��po
�q�HQ�F��R�GJ���ДC,BP�X(�U"!�Ђ(�����dȝTMB�����d�1h��]��4�.[B:B
�E%!JL���
[�En�d� K.RF$<� ��I*))m�bn"�Q!�[YD9F�er��2��D�G
�K�L�i2h��V�&յGcQ)bpdP��袷+EbLe���P��pc�B�K,�L�!Z��
�Q��G��lPN�%
!W�2$T�U��.GYbU�V�r9aR�j&�Q�ꭦ�j"��r�L�F�ԩDQ["��K(ǚ�IJܩ�9HT�b�(�mQM1ܱ��
�-��6�PyRi�rX:(�RV���$c����n���$q�u��}�1��=zM�]�w�����{�����Þ���<��J�
-\�'����#~�k���m��ގ�⯹�n�x^Y�1����h�`�N=B9���a������|��y��}')V��ʜ�Y�/�w����^�Cן9��ϥ�����s��O�����[�s���|��c��-��7����?�b<M���B� �V%�$�#�S(���;�c�+�n���B�p;S�Q[CaV�cd&�T93eZ�`rϫ\>3�Q���ku[�}n��F\B
D�-b-�^�nZ����̠c�8�L)��!D�(8�ģ�%��d$���4�|�L.�`�x�y�4�
��pb6�\��}!sowv�#�FsH�8[Ͻ�!�~�g���ܦA���4ń�߶�*��������~,��G�Ǐ�&���	4�� �UW>��^����c�@`x���Fe��mB��e�V��
0诣!fC��c���d� �r�����R�JJ�L��$hhy��a�
*��H�7ic��΃N����̐�!��
(a�(A1�#7F
�3��Žm���CD0�V�!<�޶�&�Ӑ�ޛ7�GP�c�8B\�v����I��̘���ӄ���Pl4<$��4
(sF�x	������� eH�!$$���1t0ᄠ&�\
4�۰��\�Ppih��S�f��kF���:��y�ϛS�"&	�����';>>�Ev�r���neʩ��ky�1�4@v~o�[䶨��80_�2���1���$!�!���ȁL}A���'�ZA�	�Td d Pǭ��};���Y
8��z����Hl��aM�I	)��AЦ�=z��03��،�o����ͩS���Ů��7���x��с�wid��.�&�1*98��v����(��-�����-ݜE�cF���h6�n�|47c��)��M8F(`W���A�¡���j��V�������)n�{V���?h�2e�cn\HI�^��I.�1�2�ܐ���M���AJ��YqrYk��/�u�J|ڞyמyǝ:�<pzʄ�߳3��xG~��c�@%x��@��T%i+^��a3�+&G#|2;!(:@���m̎�U���N�lh8@��Cg�������$�ŐSV�Qb�[ʯDb>3���"�s㘄��W[%���έ��F�X��$MY�f�"�ZC$[P	0j�,85�L���+D �  �Wk�d�#
����C(w�_�Z"^��lZ,�4Ƣ� cd���$��I���Mh��QDd$�����!3&���&rљo�D�shq�[�]m����#�����瑆�e�|ҟ6�<��<�ΝumL-7�?υ�=d�2�]KX:�!�$,me�Zcm��w5�Z��#�Y˟F1�c {~�}ӿE�޳����޽{����W���Q� ��������^e��G�2|��9cÏ{�=�;��K��EozwpN��+Oo����vßp�w��}}Wx�ݏgY���ׯ��aG���z_��������9ˤ�����߻����6�O-Q��e\�ee����"�S�$C��bj�����`aˠtA+�D$�q���$S��d�c��zƀ���Px�!���	r�y�:�!	,�ś���sH9�K�y|YF�[#����h����*������p&a��֤�2�ق���ta�9�Ue0�` 8�G]v�z5	���	< wwa#��q+:��-{@�-	~��}��Sm퍤�}4黴z�Y��z�^��w���N�!�X|?�5I��K�b�2m�����C�%I#$��e-mqe�\eO4��jSμ��<��Q���n������6I��3���;�)9��8v��i��h�������3������C�p��%�{�I$��0���{��0(����rv�R��L�{3�ނIu��Z#rK�>qs)k;n�[̗8�������$��FC�=`ܜ��%pa�
��([t��$�c�t��C��l����,3��YE���H�t,���W����N?4���d�jx(8�W�)H���U�њ$�@�����C��oBf�����Pa�����FX�cSE��d|ˬ�ʟ4�ͩO:��8�]#�EQ��
�i4�뎛�.��i�	 �60a!! ��S_��T%U�yz��)��ѧ�H�f�4��dL�N�CC����M�!A'��$<��Ɍ��L�,�t1�%�����Q޼Z��9���ǝ,$�4�}�.ɛ��0o�!����@tu����`d����%��s���NI�L���MUIM��$kO�'S'����DE��у�h�ĤrA57E�%��?_��̸����j�k�����$n�20 C����ǃt}�q���06E-��C��7�38y�-�9j7�:�4�̩�^i���~DD�44�]�oj˪�.�7d0�G,\2V@�u�j1�c/����]�[�fȶ�|���\�� �^Њ���sV�Hp<$�%t�|b�`�?"4n�7-�\�j6̂����g��!{f�A��Y�z�:���&G0 @�	췍��8��c쒇�8�q��#�r�'*�����{��N['����e	��U�(I�e}
4J��)��d�r@�۪#7����`F!�i��)0o��)��!�/�4䍻i`�	lK:�<�l�e�4�ͩO:��`�i=��J�0�_����7�!���-�X�*��M4�M0>5�����onY0��W��r��'�JqNu�s۲X�o���g���٢�g%
z������{:2y�M��B�����5���ϓ����Ԭ�֛g���(˜�}&kQ]��{��J����qHm\���?�(�˫!	%B۫���h��N�)pocfN�:����1�N�KL
��4@����"�26�;���:�4@�B��k�/��}�vݶql♖0ilB�8�uwR�Kp�CwAQ����^].���c�Ş;afF��a�/}�q���2,��nX��J0t�����IV[�
!�&Gt\���RK �_Pd�LnUNRW+DA s�'�ŝ��f����щ�IkQ����x�Ф�W$d���(�5ߤ�����)��y��� #"a�K�h��2m�u��u��4�Ǐ��4DLCM!�IR˼�q���EDx�,I�����!-T��1�c	�Қ��9e|A*��	���q��a�Ld@ŀ��y0>X���" o�YUD)�Sm�(�D-�)��F�C-GE��O��Pp�T4}��a�c>̔�0��A�N��ro�Z��d8T/��` d����	3B����[�(��`���
x?��2
��7���[����G:`0BvJ��E Pb6�Uj�8P	���!��!6� �ܔ6D,��DD���ă�V���i�X�@�,L�p1��wZ"�k%����e.���eѬ<5��h�&�#'��^R�)zJuzJz�SK�פ�^�y�1II�/IO^U��Rq)��Ի���e0�i%Ih�T�%�"(�m{�""�H�R[i�S+�*]H�R���I�Rq�<�FS�jyu<��^�Ȥ�y�z|]O��)�ë�4�tO������^����Ȯ%�R]K�(�eu%&���N���'����R��RrJm��K�II�e:��])*�_�]�4�%%%<�8�����E�%&�%6�))<����~�'�I���R|��|�>_	�a0����>^�>H�"%$G��N)>�U���;O���8�6JB�]It�w�w��uzJz�b�I�*�
b��M�zJz�T��IO.�%�R�FS�IK�v]�-ީ�;R�Iڪ�K�HPY����?�����{<�4���I�5��}'&|CyٿM��<�?u���,��(w���v8�Ѳ�|��M>�3���u��ͩܫ3���׽'�]Oêv�>�sb���i�����_��~9���a:=��4�|���ǻk��.�!=b���<�L�z_��
�,�9���8K�H}g ����&�~�������5&�ս��[s��v�g����w�=l��m<+�L���QC��]�����w�G{��H�������l����׫���[U_,_߻�_�������߸�j����9���������Ux��b���s�M�������W��V+���?s���Hi�Npӭ)M�O:��8�]G��V��1��/�ة�a"�,a�\U^Y��d�t�:��o��ޮN�0�0h>v!Ԁi�6y������)���y7��� �h�x��,*+ `�oYn �F��Gc���P����(: ���q�ZV;���,$��F����Sφ����`h�l�!���ru�c��`�T,)�⚍"Fr�A��gJ�ƀ81l��!���!c��ID>�͔<��� ���C��[j�V��CC/� kp�,��C����ǁ�m�|�g�4$K(c�BψxɓYy�o�ڔ�<�:u�rۖ�*EJ�.��W=����А�A����Cy86b��������v��B�	;FPǴ��T0X��<�T!O�4�mD><t��!?r�x�d8固qp��׍?�{�?�F�����w�sA�RƊ	��Ѩ��Q�K�4P�i�����6�CT�D��,��g�d�n��i/�ݏ.d/Ŋ""�����V5E�V�SGË@�#!Id��M�\ɘ:i�;�:1���,uL�)���+1�ƃ!�CC���t��mm���w����V!em�]e�ͼ��)N���<��H�'���Ѽ¸���Y�G�J�Y���z%�KcsQQZ�����b�/���6�7�_G�i��s��wzM��(���s�OY��M�̝8٤7̮��g�;��$<�����H_9��v�߇��E7E���y�����N�������W'g�S�M�Z��oy��]۞���	���ͼ���3��8�z�WOG�}+��_��M��\��G���Kc%2]]Z#���(8WS�!��h���8lcq��ςB�N������J�@�Bݑ�2P��i<&�ޗA�c�H=��2�`��B�	Y����r�I�yuj�ٖ�4�;�CC��58USfD>�cY.��G.H#Y�!t�KU��dv�~x�m��3/L��4��f_��rSQ�"U5�
j��3������.d2�I&{�i��m5���4l�K��.]�Y��Wav�aL4�����)N��yӮ��%��Kሐ�\�JeR-�i�!����\�
 h�~�ˑ�;�Ό�`x6Z�����l,���M��������{��(pv90߼|:!f>��6;6&��h�]%q�CM	�ɒK�u+G�4<t0�	kI��K4���W*骄0���>��ug�ډ��"��,�ɡ�6��� �0"�0v:�웍Uhv��_{�И!> �+Ԓ�%IL!h�6o���r48(�Fp��N���R�S�8�]G�����Yn�3�.��{ZEEEhHo>HH�V֏�q�M��z��@�P��@lv�!�hj��lrX�kٖ&�m�~c�����QpᑎL��!������.P}����=�^.�i7�&�s�ɷ�����~3�x��Η�&�1>���g�8|c:g�4�hlpPd���ӓ��80p�}MfT	*D��C�!�4۹'M�	[	!�cCC�q��Ijh^�kh�4����Za��ip������ã�c��N����
(�u8Ì)�[|��)O)�yӮ���Of���(��*���i�!xM��QQZ�5%o�F̎hr�-Πj�c{Č�xd���O��[�s�n����Q���w�WM�{4F��4�����h�M��%��|��:e�Bt�nYc�0���p�J
 tx;ӭ�����T���}��!k���:Y4�Iu�n���>lo����kK�$�btlr6�����URJ��c��֣*��Ǧ�~�d1�c�����Lr-sn0���|��mO�R���:u�q�f�0����v��= �*V�5;�-4g��q�!�Y~��w=����kv^���\_C������q}��ҝ�g�ԃ��]�I;=��~x��m��{�U�z��b_ՂV��+r�_	�	/ؙK�RO����r���%�V�Me{[����8wSK���׽T���;�UԽ3�?^s��7�Ν/J��*�4ݻ��2VK<<S�s��0~4a��;0Y��$j����I#)��L	D8B�Fߘ֝�����n�I�a����68N�((�,�pm��ti�0>~,$����:��X9�1�8hv����w��$XA����Xq�ca�,!�b>�����t��	 ƍ<a�V,���������˺Ź��>Ĕ���>N|dd�2C�F����e�>x{�����49f��.���.0��R�R���:u�q��nċ�����cYY	�2�m��=8���А�Թ:4��~,,�����I��x�T,r�����|���������,��x�]�bG�g&>Z�wRL�XBo]�r�(vdx��ي�6=�]����UƍӃ �Zl��𴬆�����-���X��>t�6j:�ئu�S�����\�^b�����vh�çN`��٬4�AD$J<Z�e��϶: Bn��Ԕa��V�����d�H��Y~yM���qJS�S�<��Q�r��gk��3�bI�i�y�f�QQZ�ӧ�Z����<7�!		�-y��� h�aD,PԢ��Q$��~����0!�R�Z,��-�5V@L!17	B��!g��i�M�V���>�|χ�:C���(����46V�8t���Uf�cZxƺDKf��I�}��塔|�L�#��
$~��ຎ��o;���@$`�ƞF��E$�G��P�0�֏2}%�0@�u$�rp������^F�q��S�|�8�)�)N8q�m�z�Ʊ]�^��7�!u*���h�{�EEEhH��]J섓�k�65°M��х`B?�H���=��Be��p�$6VW�7A�����H��
[履����ER�[dB��<�|��⣂I!�#$)�K��L|;����w.@�]�ٳf췍��>;�3UK��T]qh���f���h�6�g��T���Ô�m$�zPB:�sU��=������v����Y?��~�<CG��0�!�>$R�Jb�/LRRS�ү:�T�JJ]|��פ��Ĕ�R�U�W�rK�J/�i0�E�EZH��j"�%$q{R)&fL��4��Iu#IH��)��G��.��]<�y{uK���<�O)~���yK��������mz%8�#��Sk�R���m)").������JE&R��N�H�yK�R�#�R��jcrJM�S��o����������Cg��~����DO�<>!��������<N���]��Rm���JFR�R/���S�H�R"�DRD�DRIڗi)>�.��t�O���?�~'	�_��~"O�ǅ�']_�^N�T�JJ]X��4�%%8�II�.�^E:�$�ܔ�Ѥ�Q�EZH��j"�%$E"�'Ȉ�e�n���O����>�u����X��{7���;�﹫���.�Ϲw�)����p��lԲ��&��\�iD}|u��zs>��z#O�����=�G![���S�^#��a}L3�4}��,��N�&/,�o�^����w�d#M=�� ��t�Kb>��N�q�Ru�������m��٦�Z9�E��r���O(���
ə2�����Sb���6zT.N�0�߽�����I�����˟����.ܪw���{�ܽ95�������}=�_6��(�K����%AAR�5-�e��'N�T��w*�(��]�_~�����Uz�/?�������~�W��U����n�����Ux��Z^s�9��������j�^�K�~�?_Ɔ�CNpӆ�ҜS�R�R��Fݴ���1�8��#�IhTE�e�d-+�@P�0b�!R��혇D�˖�;�����!ƣ����h�$*�8�\���2���$I�ؓ,�b)Y(�r"bd�A!�V:�
��c��et�lUʠT����ebI2�Gc*qK���Ia-)cx���*V�۶�#�9Y+f,�6V+�d-�U.ۍ{Ӎ�����%��XԔI$IQ)
4�,h%��*�Z4B�$�HJ�Ɏ����X�ꨣE"U"e�؈U�Bp��Uc��e!q8�(�rAԁ!Im��9
�	ڙ^bn�C B�Z#(�Lh���DD����FE0�C%����M��D"YV6��)	-QR1���r�J�ҎK)`�n4�B�ē��BX�KbCm�R%Z��`�Cn�U�$����m�7k��*�Lm�2�#�\�D�܈U��RB4�cj�;E�J�V[Sr[J�1Y�;-�+��]r��MʚҕV��D44Be��T6���&��h�C�șq(�"���W�'P�"�)S�Z�e��KD̗nc��̌���TTV�����>���%\��5��{�m�>�/��׾6���9f���w=�:+���V��������5��8�h�x|����[Q��ǥߞ��<o�9�������d-�+^���q��D������9�)K�M9|Ӂ��c�s�=��uZ����r-�ª�T8~�%܈�?�Y�w$>�o��;;E��W�5_B�}3L�!CD?���&S:S�#L��%�23RG0�z�6�á��[>;�A�U��f����O����%�!l2:�à�&��*���!@Zz��2pc�&�Cp|�����\eo�����|��8��3�kU,oǯ����m;��ƔV������K�vp����:�K���s��f\������J�CfCAE��.2�/:��┧��8���ߍ����T$���iL��hӲ>�QQZ)+U����ԝC��&F�|S�&HhN�P���$D#�S��p�j��&� l��cf9��c��a��À�y��:ی�+\�G��[зR��}8����ξ��:<���K���/�5y��km���d3���x4(��e����>���
=@�&�lz0z94�CY9�M�tlg� �-�H�K��e�[e�Z|�R��8�6��w�^��_F����l���QQQZ���Ɔ�3:�D:��AΙ���?��7�ɱ�'�:izC$1F0r@��<2h��r����v;l����D'jq2�l!���I%��'���g�t��B��!E!@��$���o˓0ٗ/���PY�`���R������*��2CTHH[�(c�O3�X���H��c4��D@o+q�\[n��KcrgY2e�y��|�δ�R��8�6���#���:��f��daQr0����***�C� `���d�2CT'
�Z�l����Y���E�"M�P�������tC�o8�m��߈̡c�l#&C��'v�k�G��.�u��Ӷm�\v������S���HvIxc)�3���
$���v�CSF�un����O��۱�{{mټI���a�yk�m3jeL�d�Mme�\e�Zy��)JyJS�qj����h�A-�
6V�
4m8=����j��EEEhH;>�����������]�s����ݿ|.sN=���+��W�2d��^�C�C9U]�]��:Uڼ3���y�ɥ��蜚w��l\��'9�y5b݉�=]S���G����mͫ�h��Uc��������]�b�D�!A3w�.l�'/��t���/G寉4!рg��d20�O�O�e�E����0XB�-�0�!�ĒN��}�����뚩G8F2O�Ͷ�� l�`ےPQ8}'\�y�k�:]U�����-eV��l�F��K	���g�,��ˬ��������:�����T�Th��4C�(���H�D��C����UƟ^�8y�e�Y|�ϚS��R���Ǎ��!�<�¬�D*�[�q�ƨ�t�x���А���Oh��-Ș!y1�U|d ���ύ�u�B��06?�F͵F�Jӽ"Y-}-���ϡ��眷�[gG����R}�8�[�d����:e·����gR�H"���KH$�m�������"O�ǆg�2倅���_�����D�������-M2/sh߱��[em8��٣-���e�]y��>qJS�R�p�����]���8�&$R[I�{�EEEhHs^'FK����FU}<�ە\�HI�C���$�8����C�����B}��p��=�{|�^C����G���:8�d{�ǌ�CD(�x�-�����W;�v�9t�\�%e�����$�!nK���8|�	��Ds8̃�4��OZV��qn�u���m�����'�$*2�nL���'�$4��՘}�8�[К ��i��a�$e�S/�o����<�<��9�G��V�n��q���6�����:|��Ǥ<;f>�׶!���b�m:}���Zi�V���.�C��,
!�8|'Γ�nJHZ{�D"����49��5�����6>v�2%�b���v�����C?w��V�p����f�v%l,��R5��)��+U��p484�I�.+{ �vm�lbH���W���4C��4l˯�8ڜR���q_-�</�@x)��d�8tgT(Ⱦl��l�̓�_��QQZf���Y����wg�ݜ�W�ϴ�h����w��{�x�����>�S�HIf��L�:\�y��ƫe�.�Ž4y�iH(�p��}��z��WW�����v�	�~;�{��5ik���4��s�g-��wd�����c^o�t|������󟒿��_����N�w��������|��"T�[R��9�����ܯ�7��l�=$F�4�����a�<����f�6|P�r92!�1E�����YAD;��x�|ۜ)Å�����o&��s(t��h��]�Q�6>�\�����ތ:z%��!{>�'�(�a\��?s	�8d�G�3"m�.Q$�m��u6�ƭ�
�ˣ�������ŐFBK������x��4�_<�8┧���q�qw�u4TBc3�Ku�ĳI�$.k9��QQZ���t�P!}�d띚`BL��{�g�l��k%�{ۿb���Ø���Bxp9��������8���a��;� �p����s&�C�4�FF���t�Q����ҭ+�u"�7^-$wuɺ$����=FO�~y���	�#	�`�aw��W��BX��x���W��[����qHD���ɓ��>x���8Xx��%�Y������ �"%���"ab�DN	�&&���'��Ӆ	 � ����X�:"xO	�`���h�&��h�&��&�x�A4N"y"& �E�Ă"`��i��D��<'NYH`��CD�'舘&&��:h�(�bX��.����^<R�)m��S%)v�<��뭺�u�)�����C���<"h���x�D�e � �������s����S?C����:I�޷Zܡ�)o�Ֆ}y�>�4O︵p����'vr{�����Ne��o��i+++�(���q�s/��w'�$�g{S�����w��躗9&�}.�\�s��;���/vl}��r	/���hs95Ni��a6�٬���������y�K3������w��G�vo~�����j��{u��%Y���H{.��K[7}���y�h�\j�k�N��佭)���տN�p�ܪ������X�ן���o�?�Z��W����׻����߭Uz��[y�~�������ߩUz��[y�~�������ߩUz��[y�~��>�HiF�Y�NuN)��<�<�#���;��^먨�	~�����x?<Kn�Ad)�L���'��HX�s�����X���eSis��=�(�d_juA�ḡm��Wt]ݕx6�О��h��m����`�2�;�a�T������9(t8C��á��р�ѭSTM�4C!]9.K�+��	�����20!92�q�m2��o0Ӭ�O8�R���8�Fp�_�Ԫ̋"T���#5;$F���QQZ7[�ԹMM]I.����>ߏQ�����>�� !g��~?����ڻv-�⦌�k���ͳ�r:����g��	��v�tx}�XY������:hHC��0]L�G�f>w��~fo������8!��F��ZW*���i��O�]ù�X&x�2Bӻ��#�$�!Gãc���|��C%0(�JtQ&ýq3ԉ��n-�x��8��0��T��>q�)O)O8�������'ǈD���A�)u����+vɲk��TTV��>����}������	r�ݢl������B�WWy����=>���l}=��bF߈�n�����^�(��l�,�ۜ��;.�����{�;F���MZ�="C�.&���[6ϔ[�E�:��_'�ޅߚk���Q}߮��-�7m���z�o{Æ��կ�7���qR�P��S<g!�u��X���%Ǥ0��|;��;:���z�!��({�g��rv��*�"7cy�j%׈�I%�[�y�[�G���w���CY�?d2P�h��Ӳ��j��(vx� F�������K+��~������{��;�\!����ӣ���ۭo�Г�~{�P�f&c�ƙrLη������:�.��S*y�8┧���t莌��_y�DO��VH��M�*L���**+BY[+*�5��"Ku{b2A-���;f�r�#�E�*��4�ٶ�L,��5KbK��aZ)�]J�]~����a����jO���B"��RSf�D�n����ャ�gп>�S]�;�G��:>B��vox	e�Us��cu��c?|�~(�z�g�M\�2<�C6���<h��A�}��|��.2:+U�_�dVv���/8i�qv^a�̼�S�)��O:|||C�6]3�6�]J�/����&FN��/�>,��F\�}�I]���2�À��$�lc��
�)��n/~�2_�)��j�C��������]ʛ������RNI͔�[����g��{��t��G��s�<�0|����Ϻw��� �=�B�ǜ>�h"���>jB!���NX;83G׫�Xd0dyZ�k\�[������Sl�yN>m�)O)O8���f���BO@e2_gȨ��	��W�Hi�c�����Ȧ��OP@�<����y��8	O�Q�q���uR��a�O�>Ě��E�ݺ��2+!<N��[�CƊ�<+*��H�C>���U���hh��(�$�QWN�5��|��A��ٽ�����62<�Ӡ�0z�i�8"���8Í��Ϝ|ۊR�R�:tGFp�����h=���o�E�zB��ûa�\�y[_��w����	ϳ[�����ٯe�gѩ��|8I��>��wގgŦ��r��{͐��m<�v���.}M���u�w�����x�=�J+��o&�k���*�Ym��b�'�]���՝[��gv<����Y��˻�W��[K����Òq�K8��Z�.bZ�L�PPcw9>w�����(zNhӠ���;9ET*�zxi����8�l+�'�C�ǜ���}�Uwe�\��t1����Ѭʯ`)y�8v��M���|4��і'ü\��Peh!��6(����MC/Y�IY��z�pur�T��z�6�v��u$^/0��\)�ew�a��|��>m�)O)O8����-�>N���I=��;\�lkgշ���h��B"KO>&2��UU}w��_����9�>��J�-����3��)�8~�Тň�|�����Gc�
->m���[�'�8UH�m��t4|C��B��?���f��g	�R�\1+�X�R8ۮs�݈ϳ�$!x��RB����	S2l6j��p14_	�UYs����aM��l�C�̎�G���v�Z�[�L��.ʘ|�.)N>m�)O)O8��헴���,]��NoH���	������5F��v��p�d��,(�@��q��s�0����Z�m��Z��2�[���s��M-�_t�_3�ev��at�+8�d�`��у�	���aOA1�i�y�4a���^�8�y����0��{�O;x��Hr�w20�N��:�٧mm�I�!��9Y�����Z.���L8�*S�ۊR�R�q���cʆ%Ў��ڑV���EEEhG����x������C�=���W�$$:Y8�x��>��b�6Qs��7p?}�x���+�ĒI$4�x}�����(����N�V�r�R��8谢3�qa�Oƃ�73zs�����6�E7n۠t΂I�ۓ�!t�a\q�A�o$�N�2dca�!��χ��M�C��Tf�|C����~?�S��4,DDM
D�"pDO�""a���,��� � �4K,�8%���'��&	�0L4L�4DD�å�D�pA<"ab�D�����h��tD��&���NA&�0D��,D�"pO	��4O	��8X�%	E	dd�ǎ��-w�]H�2R�l�8qƜm�<��.��)u)L�J<~?""`�����AA?,�s����|x��~�p�32e�������>���#�C���g����>��a���9��ah!19������!G��AOO��o7�&�NW�ew��Wo���m��=��M���9	Jrde��<M|^�����C���9�V��4�oM�τ�B�Q���'Mg�����3M�W:ׄ}���g��s����w���ǿ_�c�٩�}>^��r��Q����k�U}�R��{��~���Ӭ�6wMyi�ﻍeH��[䑺B�5���իVM�H��L��s��϶{�߯��n[��9�Ҫ�W����s�n�����Ԫ���[y�~�������ߩU_+j��ߦ������U���?T�������ۮ��8����|x�����H��diEK$e���+wP��L���
�v�G�d�T��DU�����&"����1��&Ic�EP��5Ċ:)��+ő5%*�R��j��bĝ�pTy"ı��cɓ,d�Y$VP��L��S&!��"M2�B)[�P�[��
�l����őC:e�Te(ؖ&�
�ZRT�C 얍B��2�Em4��I)�����B�I�[���V	��&Q�R�(����X� �dD�J[-T����)+���R\�-i1�,b��ؠ�."QX���Q�F�W^<t�d��R�H�L�V!ԅH��4R�1e�""*"��R���n���4�#-&Ue�bE�J��Q�2e����ȪM�)*�D���I��5S+r7J+��6(� �I:�&;lI�X�*X� �-I�$�#M)��(%D�d����ӵH�bU�
�i���:����X���V�2AY��X�r�A��lV�����S%%i���c�P�!Z)b�Y1�--R�T���-��m[��1��u�3&%���TTV�]�g���7�&MO?�>��d�W����Y;��t�t����t�9��(�G-����m�\��T�^H��}�/�{�8s�7v�s���V��U��-��3KaDV?g����V��:/�N_#��F�p��:GV����~>4���&�����cZy�8�p��``P�#HY�2:��>�+�&��0a���C٫�;s�ۣ�D�מ鷃Nx�ofs�݁�́oa�>hvw��2��l�t�������y����������zw�s���d��[�e΁���Ι�嵅�����^���]0ن��i��m���>Wd��󎸎gl��C_A��a:�qr�6n�M��Sz�Z�/�|���П-vm��[Y"��$�ٵ7�>��`�2qP��T*0�P�q�Ȓ�J26!ǁ0z<��N���$ٟ�0/�%W�Lx0p�`�Y1k	�#�&/����g hGH�5٫��s�Y�e
����ϋ�̒l:0�H}t��Iг+���$���������n�UZ�R6��0���y��S�S�:�8�nig'$�T\�Ȩ��	��DjD���˴>A�O��T�5�<��܆�=y�&/�C�q���~��d��	�����?�n�L���{u��1�ok�~M���?�Wp��T��ê��6HS:4��Z������K���Ӕ�Op]o�h�t�|�ɮ�����y���e���l���Ѧѵ�S0�S���jS�S�:�8�loWg+�Z���ƇF��]H��qcz������.�I$ �h�9�Hh4l�0g����Ԓ)��K��e/�D#�2B�N�t�~��}K��x$_��� �I�$�.�֤�Q%�'�^eY�E�.첺S]�y�:�Q�>��{�>8�7:,az��4�$���p�b)�0�D�tvc5	�TM�]�����)p?�����b:3�0�
q�8�N��<�<�#��>뱔��o����n�j��l�sf��Y��v��^�EEEhL�?}�]�[7�.��\3�=�\{1�`s�N���%V��G�m���oj�.�����Un��o�|��{�X׼floԄ�Ӝl�&�k����������ovp�W�}�6��5ۉ$��7��^�G7ɞ�/�k�� Ϲ��cyx1��r�Rk�K���HwOP���`��^���tm�
� ǁ
ym�h(��艺�B�Z>���v�R;��-��0y	O3aBO�ـ�#��m4h4y/u�sGM$��G��< SҾ�I
�p C��]���W��ђa�{ۻpv;�_��e}Ҷes�vK+�[�ٕх�q��|��q�S�t����M�Gn�fƙ�(�|�M�K	_,�CF$��ތm������ha�b�!K�ͼΟ���c�������.�%X�]�?j���R���F��gq$��Ñ�m:����l�d�ѭ>�HBۀӷ�=p;��9���������Yf@�u&)c�Q4�."H�?���g�r�'k����������,�ܻ�z6_0a�N��<<�l���Ճ��'�٦���|�l:�^qJuM��)�u]�vr$*БǱ�3z�"���&�!;G���W߿7r��r���� d�Rǯ_�񯉥z�7KE�G�ms��ޅ�}�B0I?꿣o��8v]������Sc�R����p��P���E3Gn�/�{�x��e{F�L�e�mX-h�l4g�HEa����eXHi9���0=�r�<֍ܻ󡷥��<�.�Xm�:��TڞR�q�Q��k/-!/y	�a��b��oh���	�a_�~ӝ�j�%�7O9����q�m����T@��+�N���ס�����He���JB2)#󂇁��\�)�t����aoxs��n]՜;(�>�0):��2��x��Yh�B��fB�*q�܄��珃�\� ט@��(��ì8�|�TڞR�q��:3��㧴�O1T�ď
4ZM�1��+��B:.�9�9%*o˹��zZ**+Bj�s�n����W	����g<G}!��b�=�w8�:��SDt�����N�5v��M}e�������ORȎ
��|r����O��4}>7]w>�7Ǫ�d�cM������Qs�P�{^��9ǥ�/p�����g��O�7iϛ�ϖ�v�:]&�f�sI{��a���c��I���M?h)�:C�4SL.<��ߞw�G;#U���|p�I*��0�}'��S��A���q-��D�V�m[�Z���A0>�23���)L�=E���1��D��U��1��١��Tx)�~��H���I�M�zs�����[k2\�b�P/��{�H}�m�jxµ�L!�>?t��N�|�T�R�q�Q��fcF1{ˬ��*�}���TTV��Ma��+������'�&�I��z��{A���'�J*��tw����m�
,}AF�0��pY�$y�!��#�[��lk��L*|:�A�vh<S���!�Q
"IUF;􌔸.�8n��X�8+i�5��֏���5Z�n��D���|Xh�h��(�Y�:p�a�/۠��w�B�06pv��խ������N)��e��q�"'DD�0�H"'D���"&�tNP �A�QBȖ%��<'�0LD���4N��h�""i�a҄H"'N�bX���&	BX����xDM�pN	�8x��"C�'DGdL(A�'D�<"h�'���:!�ĳ�	BYe �!����yK�M���Î4���0�H"'D���O�R�iM)���Ǐ<x��!���|��y��#[���oe5��>����s4��Λy̏S�3�3��w��|�������ϧ7�jC��l��b�g/�:��>}�s)?w}a=Ϙ��~j����g?-~�"_/�Ҝ��՝�u9ͫN�{�V�r�G��A/O�ww�:�u�t_W�7d��;����t��O�<��kg����w��7���2t�J}N�u�o�!Nμ����ZoU����{�����EU|����9�ߡ�����EU|����9�ߡ�����EU\ZUy�s��wwww��UUťW��8�>�H��N��.��R�R�yJy�\!����vW�".�������i�vd��Q��;�D�C�d#>�i<����l;���k�J�h�r	�:6��5BA]���jԾ�3�3�O���80�:i�m��.��<6d D�p�'�}�ͻ��$�!>���5�v�����a|i#���ol�awQ��O�m���)�)ǔ��<xG��n�/JE�8�G� �i8�ދ�D��q���W~&~�`q̄�1���O i�Ɗ�����ʱ�FƷ`��T��G�d�$%u�`��z����%�ف�t�_�*���&�I�Tj�݃c��t|=�>�[��URU7,�U˪�%]|l��c���u�;$6���*��7�] e�vw�Y@���dX����C�����a�_<�|�T�R�q��<p���q�J e�"$R�,6k!72�tH�5�i�[�?G�~�ʵq/ݷ�\�gZ�t���b>��ｿi��v�����\�f߮^p�)�}�!�z}
�w~����p�yi~�
���s�'
������
m�{����~�j�މ�ov��U7u���zw;}t����>�̏��9������q�Z�����j�Og�}%�x9��A�ѧr��� �ߎ>iIҍ�o�&V�Օ���G-$�Ä>g�;��Jԟ��.���BK�(~Ϗ�%�I'��U���t`co�����:��d�D�lL������Um�|F�+�Pb���
KXt�KC;������C&�F��u�2��S�S�S�)O8���N7��3i3|�vc)"���Dر�.�?1�6ʪL�Xo��>!&�ѧHlw׍����a*��*A����L��
���������K��P��r�<2^_�h�ރ&M�R�_��Q��������n��xŞ���[��`�_D�Rݻl$��m:�e㹢H���ƍ�̏���~^S��х��a�_>y��T��<x��Ä8;%Dn�b���9���Z�!p��MY��W�����m��* ɽd69f��˂�+�i�b|=�8{�:(���ݭ�ޕI����E.C�=��t�A3&�&���2Ӏp3
�C2�o���p>�ޗ��������G�@���ҡ$�ן�z6>�G)�QD,�e�0S�<��:�6�󎺎���l���:�X]�cQ���**+F�'�
4L>~�e5���X�)���އsHľ���;TF��E�ڤ���o9Ě�Q�_�'j��	A����,פ���F�9���9������jJ*>:����'~2|����7KR�m�O[h�
_���u��6Wá룮��}�ޏ�J˧���8y�D��}��G��Տa_��e��<��:�6�������<>w�vƂp���M^3�":ub� �4�4�zI�^KYgu�TTV�����ӧ~��%u�r���W����ߺt�4=�����߲T"b{�=�#&yӧo
�K�w��t�y���w�|F'�$�;�N�&�x~����'RvE$������9mHSbY�vB5no��<��W2�{F�*C��'xo��k��^Q|zw��}DIDV�͙]�ٽԔG���lkrM���m�Xv;��$�6+l;G*���&O�tEd6���>s�7�n�'[tt2���%���	u��ޫ�(�/��G�}���7Ghpt۱�ɴ����T]k�v]��6]۟��������r}
��<v\C%p�,�gT�ϔ���S�:�:��ՋȄ�$�jy�TTV�U����>���t��롰�NQD�V��F=2�����%OCC���~zs���l�/�M7�|o��*Xr�z��a�
)*&�;0�zVn1�A5�^����8��i���)��tJ2m�n܎���סos�	���ڼ���J��������h���2��m!v���aL��y�R�mJy�]GW�m��Y�pJ4����n��r�6sԖ1׏d}�ߔTTV���.����J�l�8u����n.ކ�j�ꉐ�Y.S�^�^��8������	W��~�^�qn���� ~2}�T$�2���G��~Ɂ� `4:e6�;Gzҁ��B�l��%Q_��x�݇�%`ĭ����g��,Kx%���-�����l�n�)ti~&�u�So)N�O6�<㮣��1���cEؔ�m��TTV���&�+.�96;�N܌���������c<x��Β�d��ܬ.č�f��j,Q,ڷ�����C=��2::����נ����#����OV��t3�E$���JZXW��|��So�}*]�]Wa�K]�d�""+D��[�Kb۷/%x6�7���Ñ��,�E:_������tN��4�"'DDM�"A8""`�""x���'� �A��%�"pK(D艂xL4�4M0D�P�&	�"&�&(DJ8""o�L(A<A�D鐈�X��'����p��p���dDD�<P�$� �4M�tN	�pK,�(J,�A0�	Jh�8�eN�q��mJu��x�DN��&���:~??-u.�(��<xꈋ���9�+O��g�4s����o_���[�l7�|P��i�ӗ�����
=�R����9�^�)�fWy��/L�����s��]�}��{��V�&ϰ�Ok3����R�/-�%����z�Ҝ��vl�g��Db���>�+m��L���<S6�m9�a�z�)^�|p���_�Ӳw�u���W�͇'v����熆o�n�}l99�gth���9�$�'q^��t�'��,�ߎ���D��~�N-5�s�u�����������co�]Wa����N��ܼɐ��c[�UW���mw�0�C;^�i�.��uWΕ���sz�֟������j�
�a2w��[�T�[�i��YH���ެC�\�*}~��v�op�r��`�s����?����J�9�q�������Ȫ��J�9�q�n������������������"���Uy�s���Hi��Y�4��R�R�mJy�]G[a��m�}.=R�ۄq�Pu�-VDУUD(�BJ��^B	9�$���:��Qb	��T�+�h��6��KbU2��;2��F�tC ��C�&1�!:'	(�+Ir!֝mR1�Em��Gjc���)
��eV���7GR���CH�VĄ냱1�$�R�J$�JIBc����T�x�ʄEb��p��	E�E�THJ�r�2�E�'(�n�A�q!�ҫJ�-�Y���K�Rc�V,���e�E$'-*ɅX�R�HN�
��%(�"YAH�I�$�6"�ʢRV�1#E�̵���JWRvɊ��1ђ�5&2GFZ"�1���
A�El���X!���x�Hr�	�%T�jX�m�Ę�*���ݕ��"Y.&��$�W-�4!��6�xAƕ�����)[n[�t��cO��QV�]�VR�V�HEi�jGT���۰�V�QGX�Q% Җ����V���TvD�R�1WhB�GS��H"��V�*��,�v���!�G���1�+��PW%ob�*ؔR�(�ܴNK#V��r&����̙�%ۋ/��w��**6��Q-���;��p�/���+!���[û�g??�����������JsǴIw�=���G���������d��Z�;_����f�R�$'�6��vz�=�+�s�9�m���︔�W_�-�^A�{Òݘ��|�`yZp�c�����$�|κt��$+�y����)ك�X01�8��'?��黖~&�E�o	�.�t�s���k})a��/��@�>�#�-rZ�������lhʹ�-��x�;-�64�+!��L��CϨ?IW؏��[J2*�3t�q%H�����B�'��A�߯'\�n�"�0�4�0�/�y��)�)�ԧ�u�u��H�/.��Ia<U�a\Nc����BBXG��!%�Υ�pA�7�'ω$��>����Xy/���&�@���>+l���c���[p0G�z�%U�.L�<8_@�|��vG�	*���9yo8/93���M�$�������1�F����c�L���6E���֫y�6�ʵ���2ݾ�6�A��e�a�0�.:��)N�O4�<㮣��ӾH�c��+�1
��
�V;����Ͻ���[+es�B�'�t����L�p������p�Rx����?��x?�:xY%v�]s4�+�MF�*��5�h�v$�B@�m^W���Z��U��crUid4�7�S!�x	���p��ac�I	 �ti�#�9p#!;OK�h�p�oam�Xq��<��)�)�6�|t��:Ag�W:�����8�j�zޮ����v��BBBX<��IJ�T���i˖�4:���A��dVQZ������l��ǹ�WY�R@������7CU&�����>�G�EC�0gG�0ZoA�tJ���W��õ�YpDj)�����=G0���� ����р��)�nG�M���r�4P��c�B�q�a�T�;R�R�Sjy�]G\a�kR�]�a�e��|����H-Z?�IttG3a]���!!,?j8�s�ԇ][q_��N~��d4|�wO���e�ݜ�7��x.��&zt��{bW��҃�vB��s8��xy�w ����s�Ǐ\G:B��I>~�!���-�ߑ����{�yYRS���uk����۵������=<���*W{���f��B2�.d�	X���||2
�rato#��f<�N�=�[�Z����h���N=�����XUUշ.�u��������G�|=�Y��;
J�9ԭ�"A ��j��$�1�2P�~#�~�J'˽�n���p�����MM)�O���U�s� �>�^�0�:� �ʪ�u����G��)�:�o��T��ڞq��<t��qi��V��6�pX���YDm��k_4$$%�L�gr�ُ\���J*�����2��6쟊�B�?qlle6ݣ'
��w7_����&�XӁ�����BBI�c�Q.mk�:�#�:>{kt��%���������Z�O�oɬ���.i�}��WtK��;;
)��)�$O�BB;q�����ӧ�C{�L�1�,�m!L�z#9���P��L2�L)�<�jR�R�Sjy�]�'ߡ�+��Oj D]@��G��i����>Y�A�q~�p6ry��Ӿ���80�d�ì:g�Qf�wC�q����x�$���ۼ������9��_��~
t�|`���>���ua��EJ�t`)��'(�U��پ̜�
��2qU���%Hr��B�������h9o[�=�������p�(ҘS
eO�6�)�)�6��u�u��q�vRɀ�mU��HHKc<~Җh�!$�!n-� �K������s�"b��Q�2�֝2�5c�z;33r]<�CvKM��JC#a�࿈B=��3�<:t�2�(��VXt2%���E���`� �N>�d6O�:p����t;�	��e�j��m!����m��|�|�:�<��󎺎���Iixy-�1������"�Z>Aʠ5-P���G8�W��		>*�̮r��<�˿�6��g�0�C���z�xھ�h��I�{��{��v��9���O�꬞o��|��^g�7�U�9v�^_W^�̑��z_'����f�׉*3�	�Oou���/�w���f�ffw�Ok��v�T�-�� �gN$��0��~:�[Gc���i�n���r������,B�>Ο�׺�壤�!fk������8I:-4�uɼ�ے�N?)m�'�z<�������C�NG��$C&g�|r8y,4�`hr��	:�n�u�a�]R�R���S�:�:��I,�״���$Ig��_y��ZB"I�1��y�{�3aA������Qԓ�tf~<�����t|��KFo��a�a� �����ƃ�p�~���������hk0f|���Bg�'�������i�W&+f9�:<9z0va��HeۤtK���n�ˇfGc���)'���y���Cvu��q�]e��m��GTG�'DDM�"%��M4L:'D�e	� �`�
Ĳ��X�'DL0��4MD�MD�L�"%���a�,DN�M�O	�8'�{%�O�D��D舉�x�F�D{"쉢`��pN�D�����AC>Ays�2��ͼ�)�]u�uJt�(A(DN��"h��a�i�S
0��(��q]䀎X�6r�ʫv��f�g�ܽ�̕�k�n�Z0s�y�_M�����iP��k}�θ<��bw{ѕ��r��ܻ�֮9C��N���co�9o6����}��}y��H���_���j���}��{���_�̉���Xog^��ɝ��f��Hݗ����������|��̜N꺜��P�쟛<��\��~)�e���\~�g��;����;�5��\9x���9���EUWX����7www��ª��Uy�s�훻�����UU�*��9��www~�*��*��9����CM0���mO)�)�4��u�u�e��ĉ'$$$$�+�=e��P�Q/#�P��6��&�*����d!�kHl:`�w�;�N>|p��l��Ř����^�����1�Х����v��D�;���j���%5�rHw���W�����F0���GFΓ�S���``�Ks��n݆�F�a�������S�:�:��IS��"B���I$7��$M�z;8�!���4+d�����;\�UQ�曗.�̝�M�z��rm�J��g&d�)Ӯ�:8=k�t�	�@��iW�_�#bܛ҆o�a%�Q��3��n��F7*|#cdԓ�,:�d���[&Fa�e�T����S�:�:��"���'�a���1����Q�����u�4͚��-�&{RI$\=�v�8�ޮ=���U���o�8f.����폻.ޣ������=U�x̿{�}zi��P��Ӧ���{����za���t��F#�k�J�*���#�R��o���	�k������2��n�u�'J�rv���q��O2�}��ݛ���#!Ìہ�c[�pr8�(<�"O>�?y����Ð��)��HC����	��y?�:I��p_��ݥgg͟di��!��è�{6܎O�r�&Y7r���s���H�����&C��Hx�r#�?��7.�j��p��:�ͱ�r�㰉Ǒ�C$8|>]���]������<E�M0�2��6����S�:�:�ȳ1R�-y���K�K��w�C5�����D�If,6:��8th:q�@��8:?m� ���|�o�G?[Ed�N3�)���'�Yy�kn�l�5c0^�H���8l�^���!�D2T��ٱz�m{3k{*�n�ǚl�6��V��b�b9>�K�.�6l��ၲ! �3>�v�6=T��ݕKti�a�a�_:�jyǔ��q�Q�{ߎY�M�Sr��q9�[��$�G3���)a+|l1�$��(�$!&O.b�:&��-�bI:�E���n�m2f�6�d0�S����H�doC�ebUpZ���{�`�����]��dR�w�w���Q(����x92O8���4��L�<8]�G��pz��n�<=��u�Όg�~'��,]pR:�
_�����x�I!9���m�lպ�GF�a�eO)�<��S�aO8��1kb�9{�R���ؒI!�HD���(�m0?`���f��tY$�?B�����sVp���G�`z8��M�*hx94�`�g x~�i��fLL�\�RI��6o^0�G�sN}�j�E��m������|GC��#��h{���y�g�ve�����6=â�G��'YA�T1veS��ׇ��
8��QD4���.)M�yǞS�]ړ�#�x[�K̢:S����4���ưwM�'ȧ�$�H��sC��C�W��7��|��s�8u�B�?/ü�8p,�n�I
�[�>}��YBap�õd�=Gfe��na��{E������xan�t��oy�d�v{���|�i��.k{��]y���ݪ���چo��xo{�S1�Yb�w�_?�&���z�K�����Fb��:6L��;�<h�p�86p�hz>�P;��k����J$�i���ن��t��������H�4ti��d�ÓfZz�c2H`s�O��9J�ߟN�E���n�����2��-u
�~+g�T9�����"^]վ����0�?6�̼��m�yǞS�]�:�8���vK�+L�k���J��E��I$������
6���,`�F~3�?3��Ţ�$(�V�Il���<69���pd��d$��l8h�$���8K'�b@��]�	��_{��]8U�l��a���f�6�B�쓎	��>f�4ԃ��UQ�ݻ>Ŝz6�����<p��)��,O>
3C�T�N60CgS�|�;yǞS�]�:�8�
x�â�7`��DT��E�ў���2�H���4�Y��I$�ƃp��<���<NΑ�S:8:'���w#�q�L���.5�O�u�t��BT�h��n2�n�=R�q���4�|d�!bR�����CC��M�J��sG���plz�̆�m:�8T�>ā'ŉ�_���HO��CEh�~�CƊ|�
,�M�h�f�4~��4�i�0�dj�O���ީpH��H�f�Ha�r�ӟ������s�z�8|QfHQg�]��̳���#-�h�Ok
����ͮ���[޴��ۦ�Kq�AC�:�S��c����=���q�pi�Ĺ�;:~�g� �ũǎέź�I~��)m�Ͱx~����~�o�߼��������*�66������������O����윦�" ���.��C3��ť0��o!�*� +�,�>t7���(��5��ȴZDŢ��kE�"���DM55�"-5���Z"kKM�-4E��LZ"kY�Cp���P�X�Z�!Ů]m�DD�14�DI�4�����M"M9�DI,A�h��KI6�L�ZZD��
ZMZI4��--"ZMKI��I4��M$��KI&�I��I6��id�$ւ�&����$�Y$�[KK$�I$��$�K$�M,�M�9��i%�K$�$�ZI$$�I$�Km���HI&�&�md�I�I��I�M�$�K$�I$I&�-$�&�Ii	$$��M$��$$��Il�M6�	$$�H��HM�M"-�I�HI6��Y$��HK&�HI�$��BD�&�iii$��m		$$�BBD�mi2BI		$$M��!!$�i%��kH��K$�I&��t�qd�[$��MAi�-$��,�K%��Ad�Y-��D�kKD�iiKC���$��I�id�i$�ȚY&�I��!&�&�I��B&�ZkE�MI�Ii4Z(��i�ZIii$�k$��4Y&����D�KKD���kDI--$�M��m"YD��--,�D�M��KDI&�M�H���"�ZZRM4e��BѓF�eKFM5����&�i48��m25�ѭ�h�5�F��CF��9�F�ѣF��XF��cF�@`$
�*�� 0RlF��6�fF�#M�k5��zxu��K%�i�Sg�CF��fF�h�4kf�fѭ�5�#8�F�#XѦh�#M���[��f@���E(�@`�(A��5��F�#@��ѡ�L�Ѳ5��6��24�#L#M�6�4h4kfF��[�шш�m6���44hѬ�h���di�i��6FѴh#X#CF��4�F��5�ѣ����F��6F�#[�؍f#Y�ki�����0��жИ�2�[f�2̆�B�Ba	�cB͐�4,�	�	�[:�E"3B�4-�BcBm����B�B&�l��4̚Ѧ��kf�5�h�kf�,F&���i�&��&���bl��٦��̚l�ؚ̚٦��Y�e�5�4���km4i�i��XM16XM6��&��bkl��i��M�4dѓM����&��f�f�bl�ɦi��XMm�XMfMi��i��3��i��I���4�I�Md�i���M&�Bi=q�R��i4�D�M��&��M4Mi��i��I��$�&��4�Mi�4�d�I��I�КMi�l�i�M4M4�i4&�M&�Mi��ɤ�M&��i�Ți��hM&��hM&�M&��hM	��M	�6I�4�I�4�I�6D�M&�M4M4�4�E�L��4�4�D�MBi���l��o�hM&��4�D�M�4&�Bi4�"ȴZ2"�4H�&�D�FB,D"E�DКѭ�D��-D�"�hDY4YD�4H�Z&��B�h��-��$Z-&�������-��,���M"�dBE�4H�e�4H�kB��-��D�CH�(H�HkD�D�E�bDіD�dM"hY#$Z��E�!�Z-�!hkDE��4�dZ�#�Q��E��$&�!��DBE�h��E�"�hh�#M�
5�FZ1FZ��4Ѧ��-h�Bh�h�F�$M�릞8��&�4&���4Ѧ�4mh�F�6�4Ѧ�DѴ�hMhi�M"h�F�F�4���MhMZ5�Z6�kF��P��Ѧ�hֆ��h�B#Z�E�h�քM�-4D�ih"-�5�"kMAh�-�M�kDMhȚ�A�� z?ע�������ց�4Н����?���F
(�
��&`���75���_�5������=~�������?��w_�����:���X �����<��?�kY?������G����������?"���?k��͛�O��Q���kI�o��^���T~ �����������_����b`(
?�H�_�@��!(��������~��,2��Q_���Q��!��~������_������B����������H?� T2��͉c�3@?��m���0�alܜ���q))?��>"-4�~�k�t��OL?Q	5����b9�!��������X�� ��5��h
�(%���(��� �RQE`@A?�HEE#A�QSm�������`��W`5�o�?�݅a? *L���O�t?������f͛�9	f�lZ��j6f(DT	 �A�����D� T?o�b��l��M��@�#���@ �q��pB}�����Ҹ�?������'� 	�_�����u� )?s@r�`~w�@�}o��q�:����d��������}��?�?��o�2�'�p�ަ�D���䇿3����ʿ'�����l�?@������A�ί�~Ց�g�W�?zw�ޟ����(�� a���������PW�O�5�V'��h��p:C�����0�<�n��;�X����(����~�!� 0���G�R�� 
���i��?PئQȔ08m(����Jh���b��P�y�?����`�_��._�4'�uO����������'�|?_�Ҁ��/�S����t���\�U�@�����������?W���c���K� �����]O�?ʟ���#�?��xg����*~��#�����Bxp�(
����?�p( ��_�/��!!"���2�j��P���Օ��+SSS+V�Z�(�Z�V�Z�e++jՔSVQX�������Z�f��jQEj�[+R��jeaZ�ڍYEl�V������mE6���V+��b�AAAAJeb�X��V+j+��lV+�Պ�b�X�V+�Պ�b�X�V+��b�X�V++��b�X�Vڕ�F����(Օ��)Z��J�VQYE2�)B�)M[QYYEmYEmJ�)�S+je��mEe�VԬ��(�R���)B�+)YY[R���emJ�J�J��5m�)YYYYYMJ��ڲ����MJ����Ԭ���eeee�+++++++��B�Օ�[VSVVVV��YZ��b���mYZ��ej�j�յj�L�ըV(P����[V���YB�P�L�L�V�YB��J�mYYM[VP��
�������+VVV����YYEjՕ�++VVVV��YYZ��ej�Օ�j�+VՔVQYEjյjڵmZ��YYEeemY[Q[V��Vիjիjյe�j�+(���jڵee2�2��YX�J��j�VV+Vի��
eemL�P�V)�b��b�X���AL�Vح��b�L��MYX�V)�(V�V+j̬+eb�@�X�VڱX����m���b���j�e2�V��Q�Ej++����e�յ5l��V(VV�����5eJ�YYMMYY�e5eel�YY�VVje����Z�jի+V���)�P��e��(��Z�ՔQM�R�(���eb��SQF���j(��թ���ڶ)�)�
ڵVSQ��+j
�X��V+b��P��Eb�X��Պ�b��X����b�X�V+��b�
�b�X�V+���b�X�V��b�X�V+��m��E���MZ��VQ�VթMB�)�(���jjjյjڊ5���jjj�+(�QB��E2�mEVVՕ���jVSV����5j(�Jڅ�(SP�MB����թ�P�5
(R���
�++++++++jj��ڲ���j��յeejV�Vթ[VVVP�YB�+(VVV����YYYER�E5552��A[Q���MMB�b�[b�Z�B�MYF��+jee2�je2��SV�)��+S)�����5b��(+S�b�AX�X��V(((+b�X�R�AX�V+�S(+��b�X�V+j�b�X�V+��b�X�V+���b�X�V+��jQ�j5eej��J�E2������mJ�J��S(����������)�S)E2�mY����[R���+jR�J�Z�)Z���ڕ���)��J�J��m�(R���������YY[VVVP�����YYJ���ڕ�����Օ���SV��5jڔ��)�VVԡJjSSSS����p��:_�'� *� �g�?����N?�?@���Y����.�E�PeQD'�g���&c�+c����H?��E�����o��*�0�>���g�\7�p��~�ʀ���)���_��i����������-���~V?�WA�O��=z��?��H�$k�9�!ZA�|~?�pv�������"�G��#���bY�8A���~/��@Q�����Wp��t�v�6�~����2?����N?y�J��*~�w��w$S�	nX��