BZh91AY&SY�uL�߀@q���"� ����b<~}@   >�R�D��i�E+Z(���*�kDZh�j@��P(�ME5JЊCf��Z2*��FK`d����IZ�&H����ImT�[-���@4�ej�H�f1�0�12�*�4JًKe�H�JѶmVk-5�͛jٛ6�#fV����CU�lօR�=��lRUZZ�6�H3,��j+-�L�&�lͬ�5�mi�ZՖ5�H٭*͓3Ym)V�Z�Z�����5,�Q��2���	lY�������x  qG|MCV�X]f�fNN���v��R)YR���L��P��F�V�:�M�U�r7e5X���s �=ƶ��L�6ղU3I�-i\  ך @q�9M���*�@t��:�R��*�:�  Q�  �.� @*û� �S��)(��h[,֬�-%��n   N� �,��t6��k� P�q�(PgU�Ҁhm�� �À(�y� =�=�j  	�� �ך��jF�k5�Z��Z�B[� [� ��� @��^x�  ^��<=.ƀ=����@z�{�  wQ���l�v=� �;� +��v�
�֬�6�����C+6���  ��  x� c�Q�PWM�؀���pG@;��� )����`t �q���S]�`  {t�ec,٬��)�m��Y�� 6�� �p2�:uW8  �p��w#   �� 
 ��p  ']W 4��:��u�\� ��RA�6ֵT4*��o ;�<���s.� -F ���q�4 ��M9w  (����7] ��N)ւ��8( !��k%�-��֚�d�l�-< w��L g��
nÀ�� (���� 	�`�R� �uS���2����Z�i��hض�  ������ �� uܪeօҘ ��� ݜF�:`����Ph�����t/k��i�$Xڠ*�  c�OE��[�WUU
�[N�@ ;�N  v ( l���;  7v��ES����    J@�Q!��2�*��`   E=�LR�� � F�����Ԥ��4h2h i� �?��� �`  !���&���&M4ɡ�4$�J�iꒁ4ښ2�  �h�ٿ~ّ.2�p�q��:c �7�elgk�K�q���x��c�
�)���lv  
�j�V�*��m��j���-�;�.�m��0�����<�.�⪪��|e �ժ��o2�)��zڭkm��_������e�����k�2��|���j�ٵ{ͫ�f��oݚיj�+^ek̵y��2��6�2��Z���m^f��Z�ͫ�ڼʷ��y��̭y����ּ�k̭y�W�Z�+^e��ڼ�יj�&V�̶ͫ��k�ڼ�יZ�-���{�y�^e��j��W���-^ek̵y�W��y����י�zͯyW�j�5^���ڼ�W�U�Z�ͯy��[[_��m~f�����ߙ�V�����*��2����ռͭ��VיV��m�o3mm|f���-j�f�[̵my��o2ڭ�mV��ky���f���mZ�eV��kU��mk��k^fֵ�j���j���י���f��̭m�ͫm�U���Z��*���շ��j��my�ַ�Z��j�y��י��y����Z���m��Z֙k^e���6�����y�V���V�+j�eV���֯3[�+[^f�Z쵭y�[k̵��ͭk̭my�[^e��2��m�-y��3U�*�ͫ��^f��Z��W��y����f��V��k�-^ek�ڼͫ�ڼ�k̭��y�W�Z�+^ek�+^e��ڼ�k�ڼ��9�3U�Uy�W���-_Y��6�2��V��k̷�[�<�?~y|>�
^y��(~��;�EQ6m#wc�EX}�׼���{�g3��F�fs4]�27�1ܝc5��pv�ȦT��׺\��[���"
�Ǒ�;AS8�\�[k�"��h��n�����wj5�����G�!�	Ge�K����9:�[ŧ��_���������N��
�D�n%P#�kj5���z�8�A�
��G��o�q>Cf���1���hΰ��R�d)����z��nȜ�)�͋*�7	�~XGu�LL�r˴����)���B�]�zr��Xb�`��s4uXn��"Y.>�i���ι���sMoƾ��wM�Q�		�fbݻ�#&�X������1T��F��u���E܇tS�&�����ҫ	�4��7z�lhBi�$oWy.�o���lR!X�A���[�";R�\��ܻ�W0��'��'�V�I�q�8�e;���w'���z T �\��]:,f�c���ŋҭ��q΃�j������;�IZ���=L������izޫ���vR�"�	��ٲ�%�S����\��W�rA��u����0�D���ҍ��+K��ާ���쁍�ޏ�;*��ɓ�10X0-�7�3�f�E͊��6���Bc.f�����c�����qo`�:�%��ٳ�!����bp�"W��,՗7��^^��>�&����X(��Y}yA��k{�~�zpS��dYv8�-�n1#1�$��v�V�[�
�E��ãu��L[����ӍO*�F�����,â��O���
����3F)j���8K����di#w�LK�qc����bO!�s �d*V��u���g%6�v�8N$+��;ȧМ0+��L+�$L͸��4�,�\�w'�QC�VKV��I���F(����;*8j�T�&O�cG0`iV�Ɔm�R��mm�lf�r?��ڟ*Wp`N�w��o�F����� |�ŭD�X�;��U��iy�����1���s�DG`�P�s*���
gq�x���7N׎s\]�F�u�����|����ݣ�	�V�{�Ӹ�wC�uP�1d����qν֬�P�s�T�6�����P�i�k4M��H��g٪�$�V4`w:�f��b�F�я���f�u��ާZ`sǩ�/��:Tg0��p�[�4bS7Y�ڣKl�j�rkh�>�ES'Lu���ղD=4���;7,���5��<�ٍ:��l�뱈�|�p�l�k��k혀%l9��֙.�%�Kŋ	�X� ��-����#k+N�&�����@�
�:1�ے��b�mf�-^��)�4^bJR-��x�ܕoT���z�F\���w�yBN�A�ۯ�u悹�0�_ئ���G��M[���2 ���aBa�F�����͠�J�#q�r��&'0�=.�vQtu����.����:T3]�ӎ�&��7��
f��{�հ�au���Y�Ȼ����Ⱦ¯\�5�JJu��L�MZb˜D�P�VJ�Jq�@r��t�D܇�<{$|���,8:�`�&%��E�8.�z�}�6�M,�i�Ӕ��UR�Ǻ��X��(��gq��#L�43����.vW{*��-��Г2@�aym�g{�gy�qA3�6�7g=b�T*)f��­�ܠ��#4�72F@�
�vŽV�]���$|���E�ѻ5-�[7i�n�"-�(�N�x��ˬ�1ߩj췲 vfh"�8e�;x����.��,BZYX���4]���%6�n�lۖ�B���$�':Rֶ�]��q�ˇ���-�L�۔X�7^ֈ)�і�Z#R�D��"䇯f�Ԯ/f�ܛИ����yˉ"�4�6�@<�������Ŧ�����zGf��a�A��H!�XOQ7�o���KI\,svF��S9T�m#��t]�T�֖&�9aU7b͛h��*���[y�F;�E�rN���Ig^kP}�K���ӒƄ��B�Sh�oK�ww����q�\wU���v��㾪ib�2�6�Ԫ��l��Um��k�ի��o䒨	8�q�Q;f�0%Y6��lUn���Xkf�O.\� �t��@j��H�r���듅q��8�>�������F�"d��9"�d���4��/o3��w���R�Xa4��$U���oaX�����U�{�n�.pЍnņ��x)�bc��n����-�~A��BWjyM���g�C���6�T�[���s��-�o$���WJ�����YY�ss�0�-%�ĕ�3�ث���aL��,���N�O:lSI�*��V�b��0ECD+C,��Y�M��
|�V�Z��kv�]������KG� �K���0	v�H������L��I��9��+at:�2�c�V��C�/p�a계�K&5�����biO���0u�l���7zrϙ�/UJL.�4#�tb_q���ɛ�jiT�㳩���N���,Kx��o�ʹ�g3)+m��FM�`�J�YHs}W�����b�eM��G���BE��O$s�>Zuy%l۲9/����e0�d:�'a�V�k���n p8��ͩn�D� ۨ[̼�f�k6\�c:��6q� �9�˂t�{&�Rޏ}:d�lˍ �S�]� �&u$�h���]���(ܝ^�u�\Я*U���� ��u�E��9��R���2��؀C'}v���f:}:*�>U�2�q��[Z�sDգ �V���B���tb$�C�.^�-�mQ��!�bo�Y�X�s�G;J���K�*� :��?�U0-��j��n8��M�d��Rq6��٫�K�E�7��Ȃ��H��;��:�F��K��+�b�U��Ü��s^1�ծ�������K%u�z�����@��T�!��>,��a+^�Ҳe�▴_�e�qi�O56ݽ�\|v�V	�jO �vs��7V���3*S����tJ��XcM5B�挴�h�2���f>�\��Ar"H��ԝa�MR�r�+����["�k^ȏ������"�I�R��p#���0��]A�y�y��8HfjP6��4�]��+ܭ��(�W���J�Y�cwx �~n6�4����3&�CgJ����5��,]�.f���m��
>[0: �]
�[�KG�=�:�sN0.n�R-5���J&*i�I��V"��]��Ԕy���1Wy�2�ڨ��M��X+��˻�`�<Bs6r\��-7r�K����+.D��ja�U��$.ُ�+ɹ�gI4[�n۫��h#/I1�ڶ�ϋ{��h��Y=˞Cܧ'�=\��s���� �Eur��;���4�U�2v�׆��Hww��ќ��κ9��6�P\|�;Z�<�'H6�;�
�Т��Kx������!*Jv���㣗3[���,��7��&��mP���s���wI�t3Va����V��y���L�l�xa�F���Dfn4����.�^��nK	zu���\vj�@ �Ж��x�&�M,#�le�iL[h1��)�c�YQw\�,R8�-j�aZh��XǗ�wbb�A����i�1�i37A���d��X�/{f)�5�u�5��e�R��닧Ma��I���,Ƅ�Mۀ!y����o8��Ǣ.���c���r�c��n1�;���=�qh
�`��R��=9��W���"�ۃ��A�Mh��n��twx5]��e�֯H*l-8�oqѶn)����l+&���#&;��k8�b�D-����Tex��=�'�.�aj\�`�����{�U�d[n>gp����]$��� kӌ�5�֥^kq0�;X�T����f�"�|f��R����װ�;�y��'�;��%��)z\n�d�^<���O���o^��8��p܀�������ٺ	b+���>�֮��a���U"���k1X�_L�������'e=К{B�5�@qͪ�T��v�Λܣ�Sd��`�rD62��0d�`���%��csr7'IHՓp����ӗop�54���{d%��ӗTz�;������c�X+	C^ X�]���ٜˉq��׹��C��\�\�r�,'���ND���s#�ʹ�n�&<�dl^3�ʹO���)
����(*u�$*=��M�"]7�c/����v]*;��/K�@� ��h�X�dڪ̘K�L�яq�`��5�o*� �(F�k��̲��0�o6�;�^�Ճ�p�O֨޽8�d��d`����r�MS�5g�-�2����C�]�r��b݃}��oj��K��t���\9���ε�������6c��v̪�n��,�s(۳�����
�zk��������H�LuM����=���~��o��e�2���m���b�Q0�F���V�+�s&![��%Ch��X�`:�e�t�m�!�������h��������>'�h!�ehҾD5�����L��ޑ����3e�/2��7E6�c�d0��c�����l��_kI�I=��t�MA�ʻoh?1H]�r}�6o�d7��v�{7W�L�pnK��&Q���q�}50�4+�»xJ��*u�;�m't���+z�
���k���wlgb�F�}�F�MG���{��foFC�ЍD�����|�u��/ͅ��ԣ�s@�V��6[�N�����af��E]�������9P
�T���-xe�j����*j3st`��i-�hG=X��)P���i�k�_}&P��%�@Vb"��Ꮹv�	���pڡ�#"��rvQ�+�f��V����F;�bO���K-3`�X؄Ķ��U�+��ɨ��BVN]�S��� �u��m��7oH��Tp�X7%e��U�\����*�F�{zh����ӎ���.^�I�<  .��o��J��oi۠.�Ђ��+vD6���t�i��*��ab����R:��(:�5Ww�ƒ����i��G�0��i���"9`��}�Qx�yRd�>ۏ`XƏ��Ĝz���ǧ�W�t;���89���:�e[���E���	��O���`�@��_hKPݡ�-9zĊC	���.�UP֋���!(`��|��Ǘ`��^��;^�f�C�z��ΉV4�nR��������]�B�9���F�r-9ir���
��,�2!�c�ɺ���A�h0jPV_q;�o=0�_jؖ�v�Iv��˖n�m�xIkz�a��^f�S#+����:!ۺ�
���ź�J;Hȩ3A]�����*Rѹy��ێ+��'ʗ)�Y�,�5�����w��VNAǻ8ol���C^��	�Kɳܲ��[w��s|��:�%ƴ5��pլ��i,}yxx��M�=�٨�s&"Y��g)^�vI��9�]	쨭A<<�|3�5f��vcz���X�;��m�IQo��j���0�;�N۪'��십��[.񛔮9�,Չ�r2,��91������6�;,ԙ�mLIN�e�0�;Z��Í=�*�i���z�;bQv���M�oF�UF,�貭�n��W"y�qT�,�݅��ZA�0:=jd$��e�f���ݛ{��ǪQ��x��z�z]룶#���ICծ���K��N�x���pat�f���r|3z�b�^N�^�/c�[:�cjdE�^�	���Q�c�Ƶ^$�Okkz��m�ƩC���W�������!ҁQ�u��K�-ga�R�]��M_ҭR�D&�Y*u��Y�{w� �m�l���w6�⮪�:@p����א����CmM8��kyF�0h��z�K�9���憌v�oCA�Z�qW��\�w��!�x��&4?ws.�� �n��s��;�K���]W��Rv��ْ��.͚�|l��J���jaPVPTV��8��ڊ���{~%��8r���ז<%就R�+�W�:�&����:[{��U�茥B슳��so雡�a�����$�z�9�w�Ǫ�YNw&w|~�t6�g-[��m�x�%�he�!|M¾Q�&���ޝ]Ԏ����+��Y]���GGC4�9���8�^�#m�-�s�00�d�)/&(�E�@t%�$+y��o�2M[�����fQ �5�٨�y*v�囕���*�ޞ�]ɳ8C��Npm�s/I�I�E�R��h ��,�Z�ɢ�X۸��z��}4=4x��@@7�J[ӦS�N�ݽq1�C��ϤÆ�HL�w���4N{��\����3�I�vp�N��v�(����;+0⢰�� �Pe��A�X����0�A,�d޸�`�޲:gu�\��2��l�w'HP�X�/_�7� =�%e��$�A+ѱ,��Yw)�*��n0�h`��}F��u3����]}nվ�WO�&��$!�8��vf;��dʍ@�Mg���=xV������<I�-�-	�
��Qע�S����ܦ����' X`O��d"�4��ڳkM�:�`c����[���Y�ץu����3�~� �v��swsċI�ȶ�J�jv��.I�MT�SR�A/,^�����H�{?��"/�!�Ô�S �oT��y�H�to��t��V�2�l]uj����`{��"0M�  � �o8����:�m�e��x��������{����x��Sy��_I�'`8=�=�b�x�d(�c (kTGfh2%�X����h�k;{t���h/�Ip�Wm�{�}��ߌ�qo��A�� S_�!ϷgF鿋��U��\�`�2����Ju���H��ι�m�;4i��j��"�{����Ȧ�eN�C��w��9N��bf�ܩqeH��fG��M6��[�yc�Ҍ!]�C�jX\��정���3��Fa�q��g�	�fd�T�}<α�<������v>@+��|,Y\��*,wX8U�9wƅqgr<q7��I>�ß��k���1�jV��jS��vG�*gFt�v�I�9��Sk�+���jΏ�!Y%ނ�'cUt#Q��M�r�k����_P\����f�謇S{u��Ľ�h�mo5󝧶�A;�c-�7y��{u]���A���>ʸ3g&���Y2 �ۧ"�4�!�\pt�P[�^�6�ީיU)'����岕������K��{k[�oH1�����'1����;�3A�|v��#oa�zL�34P�(��n��ZrQ�i���Pj����[�j�wV0��h������a#b̘�$oNi�T�,ЩIr�p[w>��Dz��A=��Ki�b����瀞͋=�
�_�H�<�[���gχ����u����5<�CJ"��`���)��4;f����ϳ��Tf�j<�n��VM[��H�����Շ̯]e�Q�+V#���`�	�QV=��f�2s�v�d�r���]k%]���\Ÿ��7���sZ�R"x����]���s��Y�����=|{�.�'N�� `�o�cy}5���:�����bT�'�7�89y�ǑbVՈ'i9#�iYWd.��kggR\��b�9���8:�h��i�8�gĆ��Zz��+-�,@c�c!���Go3�u�r)�gx�g��ﱇ<���Y9�>\���	K�ft�2S��&�\�>�B�6_v:�+u�&��Xp�HAj_e�d�����ebr	M0��s4P{� ��_�P}�Ք!W��� �8�n>�@�q<�b��z[��Wf��)S=�A��Af��@(2�헽:'u�r��]��Ѽ��Yq�����ž���Kˠ��3.�ӓk�M�8��C,SLo?�*}gO�h�̭�/���y��/���"sD�y�e����{t�JqC����{����=�`\������S�����|����B��Ӑ�ˁ������}��ps��#۷QX;846�ɞX�ti1����Y�N���J�|1�ZC�����;zS*�K���ԅ�擵��b�/Dǽv����vI����WG�ҘM]'m���'G�)�8E��/�j���vxG�S1���k��<�*R'rnj�N�}0ἵĶ���q��̮q7eg���\�v�~9><բG\G���OYwN5Lf�$�-�K	콬FZ������]ֶ�¸����wd���V���M@��|���{IS1i�R:gJ]y�m�O۩��NN��t\)f�kf;��|xee��f+�krL�\����\�xl�E�[��׍����5��}�c��:{C�lR�	|��Ayxt�;:M镓���c�ǚ� �o:"4�g��t�r� �J��+q=;N�����[)zm{F�!̗�M&C�:�.�6oz�rO�^�i6__�І�LG��%������d��C{@u�fRǼ2���q�Hf�9��s�<���zce�e�&����<�oheY��/�KFK�4I=m�nO._.���$�
��R�qL�{��$�rq�#���)Q�'�a��t� u�V�^@Ĩ_P1wi����p�T^����B&>ٚ �4�{)�bH������ڵ�s����`�ul7l��˽�*T��򷷤ee7���1J}�0�ڕ�;pi���R�؝�Ge�|b{]cCX�Gi�>�["�c��W�Xx�^ z��79���:۾�[,�ټ���n��Zs%CFv+/��.�Q,�k8���dVe����4k#�����m���`ke�v�5L�(��T��_X��q�E�)h����ܷ�c�B��kRc���P��=�w�.�,�	�t�sc3wCS1ڗ.�^=�nuB���f$c�G7owD���;��7L2h�}"�n�N֖��*���v���:���SE��8(�[�^�F��}c�ޚ6z�oS��;:����d������Loq,׸��au�^f���/߃�;��9����y8��I۰��I%%x}X�ɹ5��&����Q���1����;r���^�ѫ#��,-y��uv�7Ogqc�S�ړ�ף��p)%Q�Ӗ&r
�^�j�V�Ke�����=tt��t��^z"Bb�:��NݾN�uKk���Vp�O}�QV�q��\y;�L��=�����$τyC�*�vTɇ�� �:u2;r�=":�;~��:�5�"D��P�x�䛓Hʲ���*-��×�����*����gZ*hʙ+L&-2B.�/u�f`�kÊQ̳y�w�����V��U�̆�l��������:�_k�'CS.��fE3f����)Ȑ�d�8���ó��9�vZ�O21�zjt���V�;q�@���!��L��Y-'�*�op�Φ��P��R\�]x|>݃H�A������[ �q��x��=�� ��o�ήC��#�t���Rb�c�e�-�=�
H�%�K�uqØS��Ru�����{j ���z��5��:�"�[\*sŁ�sK��!b��,4�$,Z+As�e�m�jMܛ}�T
���\p��w�FB� r9�F�����rV�R�=�:l��&�wӺ��houd�!fR�C�m;�5��yLt���v�J�}�y�s�k+��e�����r�{{=� �^�7P� >���G�r�`�1��Ү��j�Ds�uU�P]���"����o�Ú�������N��;ܻ(���Y�<��3==�F私D�{�%+��z�#�)%l�L}�������5�
ҏ�H'!тPőվ��f��}<h��{�>�����8T8�։��{�C
��gC,�w�gR6��o�;2g�C"��2�y�Ú��E;�n�\�V�7�{K̮����Cm����A\Z5�;�mU9ѕ]�h�������Ds��7���An��.�mK�OjLY���-�-)�fN��l�v+N� ��z
��tY50��m	x�5�4}�s{2���%];3h�T��7MEM5B�g�K�"6�úi�[!ɼ��|�z7#,�Y���y��ս�eb]�ϡJGԲ:D�a�!}����F]`1��;��n-��|�PӮ\�]v�̺=�c�� ��x_I�HۛpZ�G83�:�m��������䕰"� ��j�dʲ�����[8Q^��Z���
�a\4�ܨ�2��$_�.fwa��e'�z�V�
E��2���uֳ���,wS�عK71��tf�	�%�1������NB��7�&��E�L�����G��@ެ�I^��:Oj�_�ǧ	��/.�~�:���f�rN�c��u�q u
�yj�H����4l�)�ͪ=O86g�l�I���vЇ����y]��,1n�7Q�z��b�cOv\���V:�[ �[8��WAmc$�K��.���*���i�����I���/JE�� {�1#)]���5>��0v�[;|x���u�	b���G⯔��ڍi��e��f��Om�)\[��z#7����j?{ϗ�Gs�
�X �+��p��`Ԡ�Pֈjá�qn��$�wqPN��_�<�CJ�sX:�ni*6�C.0��PA�y�vZ��Ly�
!�A+��W�|��ǘ[D#�U��銎z�A���k:FJ�B�A�����;��T�V"�ZI\G*��T2�d�������*�'�&,�����);=a$/a4�V�$�,�2��,*�_l��b0��"��omCg_�xwVcn¹����H�#�p2��]{P꾰��k��=���*���f㼅̎�Y�*�&�J�z�ʛ�O�-���u�s!������")�.0�e��{ʇ8
N���-�����CP�EG7v���z^Z�қ���DV<Xe��hW<KJ�bʶI����=�L�vz{���ΰ��Y�N�,���b!&S�j���vge'�����'��7��v�������ōW�t��I�U�FZ�xr|�!�ɆO���1ww��pڴ�Sz�	&W���k����Y�3��ExW�ۤ�lgT����hS�T��������r�����3f�n3�.,���Ϩ��O8%���w4B7�2�{I�s*��������߼�ӣ���j��
�9:�@:/&�C��by��5��y��}Ѧ�(�\���D�7c����&nœx���j��׫Z�c�����ńf���Y!�&��r�כB��L]�ښC��'�YQ-"�
���.�`����b��Y�8J�N���m���W6�Ji)�7�ߥEv���e�۳d�[X�7v��Q_쏫M㻕�dh�ڝ�ܦ�ZW|VȘk׃d^��M�J=�C�Bm��7���]�W/���X�.'2iU4n7����B�=���w:��
�ۗ�_O7�@��t
Dn����uL�K�i�M.�ܾ/�%^L��}�8�Х�iv�̨�����N��8>�o�{�[�qq`��T��[�+R�Y��nO���Y������t{�D�����x�#�f��[�2"���=�=�ԓh}p��$�V�uF�
� �K)g�;R�)�������z0���!��ns�e�c\��������!{sGAbX��L<�Z�H%2�>�-Q�uڧ�3gCY�5��������݋�K�b	>��U��]&�9��Ɛ^�� /�h+���ɇ`�h�������ȼ��kPeX��2��fu�K{d�@Lv�]<��x�����uCv������3�\�e�0�=zT^ځk
\�C�]��w�P���P;���B#�V,�G��Y�ds�mnѸX��D�l�V��DW�.R.5�'~;L�t�;�o���'	�i���~��C'��}|'B�ˬ���n��e�L>�)��#*�f��)f�W2����ɜ��[}w���wԮ6aSs��R��z���ڒ0%s�ΪMLp�æU}������9�в����rΚ,V��Re�Y��������:�.�G>����q��Z�kCW�0��dp���oS�%��5R�+)��Qk�6�Hx�rC���~���ы���`PǕ�9��r�M�����z�:�4�*�Z.]m�%�N�;�#0���O��~(X�]�S�WL�?pփ�>c������c�S��t1}5�����Y<�=t�F�i1q�x*sg�m���w�2}�*�}�nP�^��,��=���Z�
i�ɾ{�B�_�㺻;��n2���p��"����d�N=��= ~fO��.�Wa�ͽ�m:�[\t��C�d���u�X���γQ�V<�8.�v�eͅD�3��6��F�u�@�fk՛Ke��Z���A����_���mDkq?g��.o�e*}F�X_����\�ySkH{�L&3e�/]�}0���j*=�x́�?
���b�����:��>�w]��Y�T��IWw��edU��]kw5�����fN}�j�m�̕d,-��8�ͦ����k��ux�(��v��q�`�Ʋ�e�F�"���g8ի�tu\:,Ð�i�R����;��%L��$���*&�t��΁T�u��M�0z���\��&ޑ��G�3���@��/g���=|7J�a��� 6���/^΅�Fr#t9�"yrΫu�3K��l�8���'��BF�)�)�Afq���C��d=��9{����k����W�y���T�k`wrl�)I{�)��t�XF�	�7a�j�r�m�J
���Mҍ�N�+��K��;涤���ӷ�\�b�h�ۦ�W/�h��@�٫)�#]Lq���t�=�n��H�R�S c��'�{�6��뙔1r�K4d����U��iMˍ�]�fKN�zo�YA�)����v���v��"͹!˾��Mԑv޼�57�E+ΎT�+_q�����A���vΑu��];��Wz �d0L���Z�:��}{|�,JK{j����t@��r�\���(n[ա�o�o*U�Q;<т�E�ʞ��+q�݇��Ƕ?�;=#��xql�av���d�5���1>�tJ>*���.V���C^v�A[�qI�]ۓ�R���^s��a�ǹ}��#�D���+ѯ*�WWYKw��Ȉۈ��x^mj]�!�H���V�M�cz�K\�R�l��0LG9s���4�F�Iھ�q�2h���Mb�Eҗs4'�4���Ӻ�*p�AԔ-P�9Z-.�[����+8���!WY���V;��m��I֐��dR�m̏+V\��q
�s�d�9�.�����+g�{��!uYe�L%�����VjN?�'{�Ԛ�.Tmau�q9L����(os՗D"���M�VX�B"���S���mSo)%2�p�kZ��c���C(�U�>x��͙�J�Æ�gU
�欚��G�q*���c�F$����;��(���òJM/��@,��=F�H�d^Ft��Cډ����S��h	�v�:��:�rR��u@���-����)	 .lӭ� �	Q���ob��M�� �W�fRӑ(M�<��w�-s&��L��4���nr���գ�\���*v]���5n��V.Mw��rxҡ��nMi�y���2�s!�&_�p
f8s����|���(�NQ���GدJ�^�{��[�|v������k�	�z���bH��-H0��Ȅ"4�x�5cn?
9��T��B0T������*/�X_�^��� a� %����E8�8ľ��=*���C����A��QOwXf*"��#����妲�Ov���&S�xmYTf�lۭʂ�%\�6�j�v�d:�����z77e��N�8���u'���9��ҦS_>^��:�r��W�RZ�Ԧ�둘񍖇s�NG0�wtQ˼�Ǵ��2�eN�n��34lh{|��ѯ�6��"f�b�@ݣ� �����v��X�j��s�|�^��jKT4�:���imԵ�֖�7����+�W�%�|��=�Ɨ�4G��ڹ��z��j���@��X<b� ��ypQ#��L�i�q�_Jv�le,��v���掓l<��P�+>
(�R�K�����#wGH���2SiM��L��0gx/{`˚�^އ��N.�R1mh�`h�λ|:��<��n.�u�ȫ�D�F(�pm[yg6�q�,R��wywj��@Q9�f�w�/����걯1�I�vs�([	Yu�ЧIvK����GC���J��'���N:�`��W8����׹|��
wgw���"�D���F�B[���6�*�H��R|�Z\�Ff�fwrI�������c9(�/B�X�Ȏ��a����Q�`�(<[$?�Cl�����-9�W����X���u�>=E��W��ڏf��f�ҦQ0�q(�����6-�ظ�&���J���/�͍�>������>��'��y�	�֯ku-[�+��;�d?�N7�/�*�r1�}xҢ�
������D=S���P�;��V��ر�z��a�]�w�ϫ"p�.���s�{�7ڪ[Py��X6��b�vƹ5�����j�o� o���s�t{LU�˞6���Z�BG�.�mJ7V_�ȥ�̻X� N+���)�3�4E�i	vB\k��̊�C�g�u�g���5d�Z57>��=���{T�����皉�D������]�j��2W�*F3%M��kw�7�>�%��5�꒲(/��%xP^�ctiԓ���|���	%v������צ¼z�T���Ἇ3\cx�)������}ڇGI]ӄ����޻�ZK�W��.O�&���e%%*����Rk�������W����XoL/��-��{��n��nM�V�Z�����*��@y�XZх�X]'Tzc��qsS{u*�n�������g\�T;��C�����s������kUq�K&TL|�4�cg��-*��2��a|�,G;Q����;c��D��(�P:��=��k��Sk^��U1S��	RnfŌF�#��L�)xo�kC/b���P�d�ޒ���V���2"�����1����+��7!^���04�c�sL�^��Q���?I!�˦{Q������m(/`��wӱdU�z^��Q+P��,��o���@�l�:�W4��ô�u)���/E�o���ɽ"�h�N3�ᮻ��t搦q#�#�E܈:�v� ���~�q�)�{�.ų{Ɖ�����s��7R��5I�&
Ώ��y�@h�V�*F�����+�����yxc��KZ#GZ2��s{�-�n��ďg�b��k���#�Q��;��J�������\:]�s��/�6�˥s>��j̷:.�����YIt9%�s�u�g�YPNu*rM����ukSӏ��cs����n=�C�Բy!h��q�+�q���LR֯tv����ˈ�btC�*���[��W����mvA��9���&��#8p��e�ud�ð�TR�?<�T1��9;7���X�������5
�w�'n=���lnd�deO:Z��#6S��
�U� ��I��E�7�HҪ�rգ&QX�K��9V�խ(p�{�ڳ���:1�y����Ӈ�V0��B	y��NCl��Tn�x���݇)&�w�o/�n��Q���:`���B9���\�sD�-�����N���*n�9vi�6X3	:����(��|n�m)M��5j42�e�Z-�+��F�S��#�9����C m�]	��~��f����\,��û�8��1�-�B˙4ɗ�s�
e�KR�\��Ŧ�9pM��\sZI��ck�VF�O9ތ��`�:�=�1V`��*�+,��{x�� p��,`꿂�v�����e&%�^n�z�k31���e<���ȼ�ѡ抜*;��W�����w�(=�E���s�6;tW�P�Pt�g�uR��Y.o;���RiF�2+�5ϒW;�ީ[@.���ȍ^����y��B�\'F�b��ѻ����'�P7'y��[[>�lsًN�A�*��@����o�|�v�#���;�n�[�ԹLT� MY��(�u�}�݇oR�֤6]AgM��X��������:�);�1<�ݴr�Snf1ȁ}x�0K���us0B�.ع��ܼ����r{�\�_� '�%���m's���w
N�G�V��Bm3xp���QޘYK����a��ۇ�{��T��,Ae�^���Æ۫�F���NM�_�.��,�����Hk�5��a[���^0P�O0�L_dz�GQJ��R�U�<�JA��}��|�7��c�o��A�Z��b��qZL��]|ٝcɩ?�"�q���/5k�>Ν�����>�D�]�TAs�;<���Ĥ�ݓ�&�	����\�^L����Fo7 �]�Ø����:�ZWw���ui%���rq��Y��*rxy�� ^���*p�:y.��X�[��.�c:�볩I��gr��b|�-K�yj��G�^*�	�su���j��wgG6��CV�e}�ULk	�s�G<]mdfs��h<L�uP�C�t>�ӂ�����kz}����{YJu;0��+;�s���5tB#�s��{/�kQ� b��P���yېƩWd�Y\�aU�W\T�f�I��ﺰ���[�/�̀�"�p��b*U�yx3���5�h��ia�x�,�oc���^�a	V")�~���5�5gFkbif�`�/T�\�'�y"�.v�{�+�^����O&���2�]Η�S�(ʝ�gf���s`���ҝ&e��Ϊ�&_s��)��q�B���g�����pQy�EM��Ķ�w��b	�e�f����^NH�������l�Ggz��r%�4����T��`�Ԛ	{޽����2+��"�Z��1�y���C��1�h�v��>TVe��N�$%e�75����>�A��١���R�8�Ƅ��
|K{�����Y��9��(���YϮj5��7�ї}�V~s~;d(JN�Z=4tא��tݜ���;��SC<sPQ�7r__g�R�N����� Cj�{�l�Oc1�RsY��F��E��mW,r�%��qZE���(�u����3����^Ιq3zyzKJ95��7|������)��+Y�m�oiQ{��X��K��*�M�ft+����3�BxjdV������6i6�F�ڔnP���qʰi�2�c{��K&��K���=�*�����0��{��=�ْ����<}�P#uٕ+P�d�gd�շh'�%�z�vq+.6�MԒ��DW�q�O�5[�T�,�����TSB��*�OR��v�����r|�R)t�jԻ�յ2ڛ���J4�SZG=8�J�K���i=+�A)�R���EbJ<�D�C	
Δ5]Ն�ffo^�y,��P��뾸��������!�u�&^>�~�h�v��ⶽ���k��m�޴���M���MH4���M��Q�����ݼi��OTu��6�w�V�v`�cl���i�wz��h���2>��]�%�A����C���2ok���l��XW}�x8Tp�}3��AҖ�BΜ<GB�IzW{�7�����sLh��Q�ڲ&��<���\���d���>�xz6�U��S�ou�#U.s��gzj�ѽz��w5k|eo8j��zMv�_b��"��u��x��M�n��;�`��}��Ḉ��OX�_�%4���*�L��^^�O��-�*n��8:k�k�ƙ̀�1iǣ���fD��W��Iv*�+V��<�?xٜ*{*�u�{T�~+�g\t;+m�6�Yn�ks��6��e����-K���f��NUs��2;�O ���9=��&�^ѩ��M㡡ZA��c�h�5�s�����m�D�Z���d��i��?Tk�[�{Rm� �0;��w���ͬ�@۽�wu��r�\�{��S��Oyj��%��6�k�'��+�n�}��E���ќ�����AZ�i���	�o2�o�j|&U�a�ͼCq��-�W����ϗJ�6}�����*�2vݑ
:����{�A~�m��l����gv�z/#k[2 Tn�G Ժ�gVLa������Gz9��L������r5BS�ir9�Q�7��C��lM�`����'�����۪xz1&�z�3r��p�K��u*�jۻ(b�j�LK�RU7U�������f���?M�z�D�=�p�sx��|Z@�8f���r���%�{'�p;�s�Y)p���t��Q����9��BZ���ٱ8=�F�
-��ۍ�پ��u��u�ӈظ��X����|e�3e�o{t����w�pX	��Hnó�f���rNi��!w�5^s}8>Q㱷W��Mh�H̻�@��ju�\�_�?�����˶t	v�bq	i��*u3kfK�d8*�˧_yI����Cǽ�`V!�u�N5��yzU�{F�`c���sq���p/ӽ�i9�*����V1�{(ͳ��
}��J{7�Z�-��vJlnX���ϸt��w�`X�؂ə��5�7�u�3�WfpB�a�NC}I�畑��wj�T�\Tɤ���R�]�Ɲ��CMj�\̔�sB�>�o�R��,(�5��h\(��H޹6#�7�q*�ͼΖ�T�����2Z�B�4�n�e�v��;JD�\v��SI�q`�o,!ڢ�r�G�`!���KԂ������.kf��B�V���xP�
z�[M椞t�_t���;8ms�a�������}�ǧd#���0Ex*/�� ��j�;Drm�t������6�Q�XE8{-Vc!�֮��c�V��X����ͳXnK%˼Ә�B��[vy�nKK%�i����	��m�����4Sه��vA86ޤ�خ�r 2�܎����l[2���6%Y�̀��m���U�O(0���A�d#u��N�G.d7x�	S����:���ܗ��,v/�K���VH�}��[��r&
5�])y��g+��+P�3~�B��1�t�佘ow-���p�ד�3�+8/V�!DL �+yl�6�C�N��;�}c���.Cٮ(m��b�޾�,L)�;�g�}}N�b����Z�p:�ۑGx*�.ge��-�ŕ�q��9�-�j9AH�ʉ��xu223��/S8�ḳ�Y�8L�6A[
Q��gUn�ۨ>}p�,I"�Y�J�c�L!����xT�c��km�3v�a�n���ϔ	*�)l�L�<!�����;Bl#�q���=�y��g)��t��kI�6��
S��\��ֹ!s�R���ozbx�^)V1xr%��\�D���Q��=T�u����ڱ,�s�t[�=�(�|�H�L;��s:��R$�5]�2�5�qr�RR�����IY��V�F�0��ՕK�����\����a��#�]p�&IQ5*��L��m����tFm��DfC� ����1qԔ{9�m�\X�r�1�э��%�9֌�[@	D�����g��i�����aǏ��]ko\��
̄�]��t�(>w���G����$�;":�"QBS�z����t��%Mǽ��-1R��n�R��zt�c^�8���v¹�����)�V�ڄ�hEJ�ǘ��[y�;����AI3ܪD���ꈒ,u���'��ƈ�l0r�������p���9ʊ�i.��[×µ��uv#.�x�S��PgI��7e�ai=oib����j��̎��ݰZ�ʑw>�H)<�@=�ab�ڹ�Q7���3�E��²���P3f��w-/����|�&��C�t�V��čǘ��8�+d|���B�bGn�2}zJ���V��:������!�Hس���z�c��RJ�w ^`�Fj�2:i��DU��و��WK��SdOq
�X���y�1���Dt�a� �l�٫���;��t�ƕ<73�f+7v?�p.�kz�Ū�6\z]m��(Á��ˤ_(\�;urOBW-�s���10�v��Uc�C����7�`�%���JP�gG��铧�@t��8rs,H.��^��X��G�o��<2e��*���E����6��9��)��=[�୘��@{q�30m�1���[1Aȼ�:w�Y���=�
⧻tn��H8&�@��<�� ��ݭ���i��Nީ��F�x8�%#�\�R齂*y� ��)��^k{KK�GegN�$lWK��\zNe`g(�k'^:���+n�:G�p�SkvLܩVO2e�����ʙ�Rv���N	�țv�r����U�I�|�����s�6��wZ�ׁ��s���h6(��sv��g�x6P��C�!�:���͓����\:4{2�8ޚ��l�=2��w0�c�}љ�'S�_s�=�v��|uM�N-ùǜ�Y/�~�L:"�P�
�T��,��q;��Ǻ��6"V��w�� =U����q��G c�4��m]>r��C��37�Cy�1�M�ק/4Rc]¼+� ��� �3�%q�JMΡ�fǽ���-��Oks'6_`4��^e�6oCQ�h�E�xp�j�F�T�w��<��\��.1��K�������tL�5�V���[Z�_
�`[~��UTWsv�S�ç��v����y<]^/&͛6lٳwQ��@������I��[4�$���P�B��1�hЃ e�.&�j8��1�TNMƌB�_k0����u�|M%M��{�늗�w�kGj�|�t��q�����f��9{�����[��`-/���:����s%�փ�vVf�G�T��E]vh.ފ��d���n�
�\��mX��@�]�'6cL<�&5����f�"9�������V>ڽ���5�n]�2�;ݣ\|z�93�9l$�.̻�A� �ܛ�-�1�Y�%6���K9��.	K��^ej����Z�ז�R�k���^�S�L��WǻH��o���!/*׵}{�#ZӍ4N��ဏ�]�GӼ�w���<���FǾ���
�1�����������Qfcln"VnK�>�R�_T�ژT�5���6�/D_s����r�#�f�*�����`4o���7N��Jҝ�[��^�]f��X�H񚻼�<�Ah�Zk*�зC���U�߂��jh�w���q�^���>2��g?Pǋ���|��>M��M��똆�M2�<w��#X�w�bc�c�Ɍ�Ń��+;�[mi�����-�4���]���:�;R��W��bV�]���Yݱ@�N�ém�Ǿ�li������;1[���g�}�I�[��\6	��r#$��f������zw{H��������̀���r� r��Ro#��SW�t��Rt��pѣ��$��c���2�V�xiV��j3%��
���l������4a�$��
Y("�+����A��-|I��A�������F�)!���4�bFKJ+�*���2B�Q��-��2\?��/_;�@cAF��&,hS�JJLY"P$�D��n�JaL�$'9��MBL�b0�F���I&D��h2Q�Di�H�J2�)
�� �"��TB�D��`���0�&"Li�I��]a�4(��b0"E�)&&2�JH���I34@���4��`X��(
&�Q	���1�aP�J%��f��`a46&H�!�	�e d
SBJ� �A�
E$K2����	���B��DQ�>6��q\4��H��u�O7yOQ��I�qc�N�N�>ӔHɒ�lA�&^Eh�]�����N���i��wΏ��s#�T�v0`�W[t,`~),�p?}��g��:�%p�O2��-ô�[�*N�k�#���扵Kl}o3`]�"�$��N�<��.�����4��{�y��h�������~�׼jD�/}9p�}��O�E��[� ��9�c�$�	�����lqq��y�A"�b0�ۙ�wa �y�"��0m��F��7���Q����z�7y�ۺ�?>���n����/Ax~_1��^����I|'��g�ey�Y��c���ޥ��<ڇ��d�|�ͯ&���"xx]|�{f�����5>�*P��^�'6�͑3S�y��{.�V�����[���	�yz�h܌-��v���A�7�;���^�7A��ElU�sVϔD�y����{�(0$ϣ'ޣ^rnOi���Q^��u@Sܑ���s�Q�h����?V�r�9���˺�6�?�__�{f+�0"K��f��O��X��K�6m�������ʽ����.��y�������a~~%��	���:ݫ���/�ƻ�T����&��t�G;#�4���Gm��:��چ�(����E�t��1�LU�~���GnE�d:�����w:j-i���Rf��Oj��*�u,*���wدϕ��~�H}z��;���ܑ�׫���3"����<�χA����\����h:|��ě���"�5�*�q"A ���~�41D�eo��p�$��=Luf^Ol�"z����&�t�ڢ�����W������׳[�ӳ�z��m�L������٬��4���A�w�Ǳ��>S�*���\}�;�%����T��§��k�1 f�9G�2lɶ��P��r���	n��G2�ji̊kw�n�6��np�pti��&��0~x����Wv��/׽:�~�U,��h��(:��|;p{�]J>�*�1(Zג���u�Gm�?A���{d�������xӱR�<���:�5��NƘ'Zv�q�l���$�����=gw@��l*}oO(�`Y� �۰{������;�B�o�S7�QVs�\k�`�����z��5��G��#}ؼ��e�#b�	�I������R��Ǌ��T}�V�"> {y�N>",��A�w�#�۰����'Lm³����=����_f�tr����!{��]�/{rA6?���^�񮞳��s�?/�����p7^z(�2�g���}�F�S��}Ut>���hyw�γ�Ș�3h�A�<݊�������>;� �~i�x.����'�dW��ǯƲl�!&���Q���7�{kP�)q���j����\�#ψѫ��zmc��9�>�B�t�q$��`?]�)3�k��Y1ǵ������;+�閺�������_�q��%W���&�'���I#�G���Fz�a�k��֧�zۑ���X�h&�?CC�1�K��v��ރ�d�)�ʨ��xD��'٣�n�Y㫠��)w�@:������gR`񕚤u�Ow�~������g{==~�.@�3���]^̯W'��i�~勽�S3�Z:��vBؾ����R�Ɵ^Q�c`l���\X&�MD�3���Y�;�K���H���<�;f�_��º��]�dR��{C+H#i]�!S�2�Wԯ#�3R�������=���/��G������Aˣ���P�ԡ+�Ls�D���ھ����&m~c���褆w��)�[+cv�V<}:nh�Z���2u��f00�9.b*[�8��z�T���Z�ru7ݓjy��O}�D#�� ���z;D��`�_�����sk��q��#�����L�p��='&��4�
���T�i�b�l��y�o*��>�"�[ݚ��z��4D�|��#ٜ\�S|��L�og��,��z�5���=��$�9���t�Ӈ#M�zO���1�t�IE������]���yO���s�W�M��2x�K~��&�i�����|nܜ��6��aNA���ݟF�}����ޙ�j�n��MG�c	��9�Wg}�Ɇ����C�t��U�/����S�Ue.#Ʒ��Lة=��{Ӷ7jI��wLp���'ͽL,o�� ]'�Hz��w��ho���R���>�]!��{��_���zBs�my�{U\���EmK>�_?]���7��cm�:�ǝs�~��C����bڧ1�Kf:�����ꮋ�O�+M���|J���Q�[7�����j��$�c�g��y�#cg�~�v`L��ki��ײg���,���]^��VL|C�g�Wu컽œ6_-�֩��W��nt�Wv�b_tt�;o5�Q�y:�ŗ[���ޜ$���=�7�d�Q4�z��ި,"�_���v�td�RRK�V'��R�s8Z[��)I�ծ��s���8s�}` ��v��J]���<?lɃ3pO;i�ӽtx wk�	7��L�7��̢.��ꧪ�^��E�l��c��=��N?|z:�3�6����R7&F�9���:h1qB{`��9wpx�$�+۬�`��U��3�����ꞎ����6��]���/�gb}��s�l��:�G�Y�ݩ�m�sI<o��G����r��v� M��a�Z��ؕ��rD������'�t��=�'�>�5z�	�3�Mpzz��^��WmV	^.�'�>S=�Nw�n3޳rh�s�ռF��	�:^��S����&٪^�f&8��������s��^��w���S+�br�[ڑ~��繍��	(�s��z�E^y��^=k��3n:�Ք�+wq��/~�&F�R����^�H��q���d�E�ݱcj�p��nN�(&��g�JOb$��af^&��h~��&�ŉ1_k$�v��/���v���1u5��D���:i��dɫd}ä�xb\�IGZ���bo��J���k�^�3�3��k��6��{^˨����6NG�fV�j{[F�6~j�}�嵋g�C7��\�G��5�ok�^�u�7s}7�ݍzf��%���an4\����Fv��h97 ����C�|�u�}�P>d�V��'����>�F���0����(ۢ�OȢ�{���r�.�N�eG2z�ŵQ��5rV��>�^�����+��V��A�c���&\��!;�{��d��*ٿ3W��A�*�c�o�9�k;������$�ߺn�;���Q:I�5 ���bs_d\X��2�QZ��k=�^ھ�c�b<_Ro�J�qO����H/><}�S�0z����G�v�����^��7��>:H���ρ��{�E�x�/�}w�sg�n��Ŝ�	���z_�C#c7��������P��E[a���T�Vv�9+	���X���t��q6*5�ǧ�r [_x^�d%�h��=�+��n�*�s[�;�����ލ���i�ۖ����6�_^�@�8��H𞹳��7R�n��S��j�'T�1L�n�ֹV'�{�ӧ�1���Kc=�.<!�~�q��'mg�K��)��G����Iݦ�R���o���zo����Yw���lu�����{Uj4��}���k�pqf�Β���9<0�H�ƨ>�|G��b�<� ���_,��0My��_e��$�A�u���l�_Z�{�ܮ@����';z��Օ'�;b6�Ƚ�����飦����b�d �U�:r�>�����k�Q�E��<�z����c:����E�G�\�u���s`�E��!�|��O����I���W��z�&D$$v%Ϻ�|�4��.�dY�ޮ~��{r�m��})�Jr�zuc��w��S�7���}K���P��U�{�y��5&���өr�	n��^�n���{!��m�\��ކ�&���T{U=�η��v�	
i�l����q����7^�q%��ݙ!Gab�mմ=iw}�s���������OQ���U�s�SW���2�C*NQ6�:z�CV7�w1�l�t���w���쮍C�R�3j.TK�w�Z<{M:.J��O~�̇�t�X�"�H��Ls;�S��<�Z����~�g�)���9��J�R1���:]��9{��Op��Ԉ�	xW�=����LQ�+_K�=ޣ��K��Y�í�7zD$�4.��W�*�\,�A����-�{՛ު]
�b"A�6{�4���s��⊧�־�}�w��0�y�P�L=ܚ6H�w=m-\��D�퉞�>�R-�Iz��{}�6y�ڌ���7�W���(�N�d;l�#xY'B�R6`ݧ��g��P�$��&�g�NU��#ǯn��{ڳ�7�)��4��1������z��|5�5��q4Lq���9<�ū}'\�]�qԍ '�����(OT�kD����x�I��x�G4�q':���oT���>���Wƨe*��.���A|�w����Y���:�qׯ�e�p�}�z�o�������[��DW��(wҘ=C��l��G���m)�.)�#V�]5��_{�ʕ8���.�+�Lj�mښ��<��&*�\�x2k{uȻQ��wM�|�N#��Xg��nE�bE��E�{�A�H�,��n_[�e��	)'Fz�c�W�D�[�fl���^wD�:���s����!�;�,$�q�n��ζ�ί}w�맹��}���Df�"��;���P	��cӦz+t^��[����d��>o�~�+��)�n����)+j>���S�~߭��~�T�la��4iɽM��=�v���Pn���Eد�8�ڞ��qۑ��z�{��OM��o8���x=���bߩ�x�k͂q�X������ݍ�D�^�|��K���,��~����t�2Py��^ڗr<���w����V���퇯C�3>n��߆ymPg����A�4���ڎ�'7�A��|I����(����k�+��vN���%��a���8]���ݞ#3v�+��uq��ʹ2�{}S�s��ğ)�}*�Ǎ�6��]tlEG.b��;W�s��kH�"���,��aU��y��ux��S�rɠ2cd6�9^�L��4 �Sy���k�S>�{�ƺ�Ǌ�R��e���42��F�m՜-R�cz'G�z�2��{�n���b���pc3e�����t�c=na��ow�!51��l�Vh�{4�ߣ��f�Y���žC,�k��};�
��^�lG+��|1͛���Y�߾)?��/��D
�gpk�M7A7s6n���Xh�py%����綠��e����n�rE��=�]J�ӫ^��#٥����6�^�C$�|�ͯz{m�Y#ڐʕ��0�L�gg��y�I��߼��=ܯ>>��������^pM�ٿ]!u�����xdW�<�#�����Xd߫�������1�||���p7^˨� �����-��6��w��S~�[���'Nz����k|���-�ݤ�`���1t�<�=b��2��;�)��}8�~�!>4=��~�S���wo'{^�&��A&#��Pߟ����9����Z�)��=荞��a��̖=	�K�2'9{����W]P�N���:�ze]V+�,"\�#Σ��y���~�f��a��)��3"��j�<~�ϋ������{޷���7�[��{����{�{����߳$������}�#47�6z�ǃ���ˣ��E��{���nyBͣ|*��߭8��$n0c��=M^��xr�D��1�W�f�`֨�4+�ގ�r#�-|�F��l��:[0pѽ��;�^ 7Ԁ.��ژ�$0�Ís����"w;&��!e�V[2.�2�/>P�K�s���&K���ꖚٺ6����)�L�4�Tla�l�Pb��1����IwN����gF�Q��x�N�6��K7onDd�j�;����bG�/-�u�һc��������Y��$�J�c����ࢲ�yV��^��Z'�z��{�W̏o��ӘEȥF����,u�Tc�L��*���Л�5<����¼1{u��� ~�U�~|��Lj�y�hx��A�=��n��v������Ɲ���v�n�����k��)�+�p4R����.������[���b io7�1�C�sT�!ywd��袍�&ǵ�͑�Ϗv�a�u���ax͔�Z�[�$�#H�z��o)�sҳ���V�����`��]��,�OL]��25ه�P�x���}���A�[��m���Zvuj.��Ŋqifbێ��wv�l膮"��v-�Yz�f�u	Sx�M�N�	B����kJ�XʚH��A��^�p��9͏}��E�w��ް�̵}r*f�Y���q� ���@F(�o,���s�p<j�s��W�JL
���>�x��?>�)��Ԧ�dl����͎|�Y46��-0~�ţ��~��p"�H��p�k���9���Md�y��R����ro!��`z
���|�!e+1(�_�Wݞ���K��Z��@(�n�Vk:��9�ch���z.Aj�.��'k����c�s�y���Lj��dU���;�H΂z}�|��O8��2�p���r��]�\�� ���K�K��cFx�nā_#L�aכ�w� FU\uv2��ܲ(7φM�9�6�mP��������{��А$t7�1���ޑUBm}���Ce'D�9]�)Bڊ8+�輛�H�Τ��q��">ѹ�ɐ�mP%m�̼��m6���u�Kw�0
wW֮G̗�w@�ˬ���ԅZ�y1v��7�	���v��6����C�9(d��oT���s��\ lo`�5�|6�A�v�vN�3zo�_n)����[r�Oμ���<`A"�
���k�0�'�4��UM������x����ǻ��}zW,����t,�kv>��LZ��_*#l�ö��m��L&�w0��s��=N�>��
� C�@���Bד���1L��\}��|Yћ0T]"�޹+��iӃ��r9�<�4�n�\0p�b.b$��.�RFw_c�^�A],�X����a�G:�v�)�R�{4V�7�b�QFmd��X��z[�W<n{��M�y[��ӗ\2��EJ`�����S���
��7��uLDј�(�4�&	2iaI!L�CABA$�b1�!2I�$R���CEF�P2%3� #IJA&a��&E�%s���Q���:�u�I�]���4.����s�黝e)swn�us�u�;������]��\��ע ��Ӻ�>;�z;��ׯ\Ѹ���w]7sp��G.������n�2�κ��u�]uu�n�\���wv:����ӝqܙ�`G9r]u�]�ܻ����������ݻ4�;:p�ú�Λ��SE�oXw.�չE;�ҹ���.1�q79�q;���w.��9�2���.\��(渉`���o}�������n��KyM�=�C�k&���1�úIx3E�{�gi�ѱ���"���wRj��{)����`٣Il3�G�=;-ۼL�\[	��NF'Gg6��oKW(H= �����%�[�F�S]��~�8*�{s�k�I�������}�hdB���{d�-C��x��oP��4�4/���J�!^Fd��W�����с��j��/���S/�8� �斑����s�OF�L�PEf�;(2Y����'SsK;雅X�5T�n����{A��oM��ǻx]]�`qm��\��_�U�J��W�x�M�=�n;*�Ϲ�9�~\7����[/g�{TgZ<���8�oV�^���P2F�(	����E�� ����=����dUpE���ܱ�DP��Q,��Ji��4��#q�gOMn��J�.͍��MP�2S3a�iG� ��<�%:O� 	N�@�%t����/��i�~��yw���N����$TJ��셗�ċL��AR��=(1�2���q>=J�r�)�C�E*�\�Ǟ���KbՍ���xTk.;zoay�{�"�@@��9�kӳ���t�R{¥�l�`:��~E��\�4�R�J��+o�z\���� ���1��~k9Ĉؖ\�'�i����Z�E��y�����G*�c6���#ʕ���kb���[���qR;��li.d*���2�,���3��t1��<�ەܬ��o	p���`��T6+�@�=��bl3�6���M�d�mIR�9FƋZڳ�Ջ�E�������`��+Nb�E���ּ=%ߏ��z��u}����:A�wn|gi�!�;|���|!�?�+�\����X9�ļB\C\ o���}���!�Ϻ�wnѡL3�H������}��w�3`�+Oח�7��˛��\���X��Oշ�� x��@���� ^�����v]U"�Zܕ����,���:}�g*���)8$�i�����⢋PO��5��0뜑=����k=];����h~gb�<:�[;#Y+ޠ��:���4]��f ���}-{�4�s[�!�v�kMn�c�iռ��W��K�CF�sO�L/��>��������q�`'������{,�B!��̍y�����!iL5[ֲ�91?��RL`�$���ݟ�NS�EI�wU��!؟��y1���"�p�k�����%r�P(γ�l�*�Ξ|9��=`����}�y��z`�ۛ�t���O��;[���u�8��V5r��_��	�8�%t� ��[�VT\9�p�oB�XfGJ�.S�����AAqk���#:ɀ�uϽ�-{�'V��ʩ/8�yzk�.O��E����:K��)��E�K�}.�9-�>չ�'���^+;k؛Ǥ�<�V�<���SH��KkFT����X����G�ʁ]Z{���	�J1`f1N���,-�>v:�����.�4{1��9�s7�Xt{��2c���/�t2*��oqŸ�������k���9�������� &�D��4/a<&�K�t�?�No��Bժ��[y�Qv^���M����`�x/VE�*3���i�H8}r`��bGa�m3L�qx	����De�U��gb:��_�<GS����~�/��-����$ ��g��!9���a�,�YT�e�=��E�*�2��[vZ^�w��l��e�/ސ̴��v@�vng����]؆�|��N[ƨ�ǖ�lk%���N�]=��7�'XJ%s�z��/6
�Ƒچ��I�L=���M��ۧ��n����ΩC[i��Rp��j�I�d�,�j�y�إZ�A{�������0uшwdݼ�īL`Zؘ9mg	�(���g�5�P��pNek�eA/m~������ S	��/g%��Y0�h�m�P�TDy��
9�@|.hN��k:�jR�o�?Mc�0�:��;��v�z~%�N9�ZR
�o��yJ��b���} ���4Bax����쓫ޗn�9E�)&C�`��776��B�@e9�d�.����ϫ��������hy�D<��s���|n�->���g�4	{�:&���9K�п-�_����0����xi7�5o�i��1Pr���c���sX$��X�����{,2�ˠm�C�[Yࢵ��B����o�gH��$,bS.�h��q�uL�6��#ݭ�q�f��������u��<z�������f�ސHz �4��>: eC�m����(=��"Ү�_N$+�Uk�5���t&�6k��f��0�z*�!H��H��t�P�:)���f�ou���9Y��7q��3L�$���K窣��UK[W����xaT]
6
��z ��]Zl���Xˈ�Q�(�x�[�[�~-����TzV��x}�����2��B����m����ɥ��U�ƞ�������.	��g�}�q�^��HM�x���<��Bdޅ�-�����7'{��>,�LPR��ɶ�5N���|mw��[�:A��	냂�9tGWe3�I��#s�~�+v_����K$�9��F�
�|���'��}h�a�$D&�\�a�}�|��g�����N���l@�[%�Y�N�X�R���c_����<��� 갂��Sk��4=W5K��;pYf�PD&��*n�i;�U�=޵��ʂƼ�L?5'��|܍Ȗ�{2�6��;�ט�PaP�� Y�}n�٤��Ͱ-XNP�Uz��e�)���okmE�A4R�	L�<6�^sԺ�b���}��^��o���Yw�)�P�>[ǡ�U�_[����w��*Lr��K�갾>�%�;�I�����yV8���갂�Ż��<q�xz�jmu����}\��jT��bu��G^e8��n�:v�����>����6�2����Ⱦ���x=�#�:=í~oP��mW=E�|��a��Z�U�♋�]h����L�Gf���t+cZA��moWÕ��� �����h��cƎ���7���u3CO�S;�3wgr���K,w���C�'��p�W����y�P�`<{D"�<�\	��f}�G<U���׎��O.Vd�ce�����C�"�*}�{>�,��Xh�q'�/�oei��+w�����1����E�v3]�g6�����^H@B|�T0����?7��%82 !�e5R��텡���Nρ��f
y�Y�=�`��xsf�i���JWA`ÇoV-O�iч�T���n��[���E<1h`ZZ|B��Nnj}<�6"��n��:oU4W�Gjn�92�;>�a~�Z��w$:�l�zǫxU�)�08���Ϣ���株q�V6�����l�<u�gu�v�voM�����R�4��t�y�/x��O��[�����&�-���p��
�DG&�U�/��ow���Rj�!8��ȸ
SL�Q�����9�<��;�?np�����K߿X�8>���16��<���֌Hᷡؠe!����J�������FI��E�
o��U��M;�����|��P�F����k�/3�Cy;S���Yج�]/�[:��$��Ti���g.T��{��67g�r�}����S���X��އ}`~���$�tD�I��Ju���&��ny�>Eæ��M�1���������B2ʹ'e5�2���B��T�ሤ�s@��s`m5D���1�ږ�P����3P
������D�?�o�Xx�WӦ՝,ז�]0�E����`�JN���Qz^���y�@א�� ��#�������#��\?�\�z�w��g�9%����\CER�F^�9��z�>���C��8�c�~~�BrD�\c�O:o��ݗ�.�FA����o��TwU�>gL��׈ɷ��>�S,ٯN�ۻ�Cs��ZyU>����2�+��z��'�t&�ӚMVJa��5�:=��&+��_�?��C�s�`9K\
�f��7+o{�u�cL:lש�t���Gw��N��i�H@:S�2	�[�_�׊�c)3{
�Q����!/���v�:H���c`k$|7�?<�u	��h�P�1`Y2����^�o�辵W�3�L8U�,��o�ȗx<y��[�<:N�b�)����i�[��G"5����~-����&n�����:g��W�, ���&�j��=��Y��jСi��-{t�O�j��	g�ޘ�xUNZ��}�,��Y<�Ъb�=�@�0_q�4��*�J�7)y�!������Ң�B�*�-��e&i�]9=r������k>b����?��8Q|�R#c������^Fa�[�Zz�<���l�w����B1�=Ų/sW>���/��s�B*�ų<�f�9���d(YT58b�VJ^)N��l�*�c	Ο�]��!'U51���bS�Mj���1D=�(Mu�^@���'汆OK K��>��|j�x�sn�3E.9ڢ'��Qq�3egP�)p�.6#����#\ɯf3��D ИlZ1iՅ�B��U	�4ym�0VhD�[KLOZ�y�1�)�(z��D� �K5З����f� _Jb�D&I��Jse*��JJ��9d�\F�c���r�t�Ǧ�ΜoD�#� ��lʀ��b}�fL�L��'c{�|��ӵF����%�V<��x�7�����O4[�!�!�O�= ����o]O"�ƍ���wn�s-�GQ���91��3l���9�s���vk��������8\�!�n����j�9�cgUMM���]��n� '.��u&r<�Z�E��T����ȟ�H�;�>Aa���f�ʴͳC�F���2Ԣe�Cӱ\��&�Y/�V����] s)�J�����}jތ��o��[Qi,b.E�{M-z#];�t���[c���,�d�]٦=[�9�VƼx��t�E+:Oc�%�i��D�!]Y*�⫞����k�1�)�V��0V��o�gm��O�*�,��@�p�Ԫ��bu�D�n���:�g;���v\��������7��5��`��ʃM�0k�9���L�[���?JװT���P��^��Fb��^)�6�ٳAc+{�&��d5�����춳��桅*���8��js�BM
��WuO�wrf���K�z�-A��2%߁p�4B`��o���vI��z]��5#X�y��˘ؘ4�0���l�Iv*�G�iD[��_Z�.#4F�C�|o61�òc<m;97{���@wS��ȴt�$?� ��Ca�ʀ�xc[�q�F�b��iV̆�>����<��ME��Xͅ�Y�Pyj��@�r�"k�"�)�P1p��\�ji�,�5Y�q��L��|`�I����{�1��eT��yr����ԉ�
������I���y��b�~�ط�m���
�����ӂ`��q�>[8�Xکnf�!6X���ɽϘ���a��^���ly�m7܄ۡ;�B��׬z���{gh���H|�&B�|Cu��#��K�h�2��i�6D����L(JE=�[���z [���<�t��	x'=u�����U���g�n��ڒ��@�ֆ��_5��oq�a�ݒ���SI���xNn�v	ujkY���@����8�R��gcYT�`n!4W����= ���ٻ�K�59q^G��_N�J��ێk��2&1���k��ܛfq۽�c���}���L�)����>����2S� �K$��]%��|���+�X�֊���Oϲp�<������@M�5�"D��Hyb��ʥY��oL7q��-N��drr����ٛ����X3cH� �G@LwУ�S������֢��YY�,m�~`4�V�e�Y�r��̺ц���p�N@s,#�-�"�n�٤�S���b��F�Gs�WF73f)�S����;��sn+]x��x���ߘtz:okuN�6��Z�X���&�J�m�T6�?n��u����(�70ͱ��d.��c���_�x��@4�E]�[Ɗ9���\m�R�G:��YGS�(�[�fy��3�؟�8D"�L��-�:хn�GU���x�r�f�v��K��I@���ϰ�i.�:Ļxw�Obꋋ�&�n� C��bT�=�;��o&�)t9BA�!za���q�':ʕ-�Bߦ{ro_���
a��g��->C!�V~U��`b�`ޡ�}���eg���T���R�8ښwi�}R�;2�c��P�݅,�3�g��Joss�}ӭ&�S���0��"f�"<�V��{��s]�#��ws- _T��}��98��JWp�*lϭMT��J\�T���|_�%�QǊm��4+��E��x��p��������Z/�G�{�����m;��]bȁ�f=TU�.�?�P����?����^�*}9U��5�S77�[��5�����5=�;y`jW��5�����I���P���f-�2/���O
�UX��藸8���׈\ӷ�]�;���F6i���X��ߕt��(�^=[ռ�,>;ǐP2pD�Q�M���=RO�=zE��u�(d���'9D�.R�d}(�kw�{l�uފ��;��9�@�Q��mQ�y�5@���B^�/��'�Iz)�|"S�P%�i5��6���ցK�-ݦZ[�X� �k��+���[PT�m	��Ƈ��W�*eC���T�ሤ�g��RmC���n(�Mc��a�J�s@F/���ߕ����>��g�3����.�1E�C��1%��u7���_��[ތ�y������9�sL!p��Џόxr��+�Q������Wp&��9f�,Q�/�R1������C��$X���t��ܣG��v��*���쎵���Ә�ܠ����)?5�2m��O�D3e�b�ٶF�{˿���ߛ�}o������{����{���~����OOef���rT	-��<"d$v���x	6{!+Ǹ��>[|{��������\�]����q@d9(�h ^HVk;�e��u(�K�N�����'�UL��}sJrwD.<����?{sB�E�S� �ueV���Eu��C�������go��{Ny�-aC8-qPY���2�S�^+�[�FJ�X�v�����Hd���l�2�اga��fZ�[m�7���Ӕ~�� �[@�a�u����I.T��B��w����"J�o>�(b����;����ϸQ�64.�².���M���R��̈dz�cr�ӕ���+��=�E��c\�Y���*���e�O��WK�;0&�������J�vg����~�� 7_+� �wr'*�#Ks*�=^C��'P4�Y������&���,T�7pMqT����!�����6�Ǧ@�ER�P�Z"��E�S?e���{�z�c�d8C��ʾ��&X��*}=��R=>�r^�|Wq~} �i�%@���L�#�����0�l���\ݫq5έ�!��r��6�۫3Vb*�,Y�*�7�qjb�4x��䳯�^ٔ�v��+��V�xy�ol�k��ui�֧�`��
���ܱN*�\�w<�V��)4M��vV��;���$�����4 �N�G�������@Un�Ī%m�kP}�v���[�b�{�篳�4����.z8&�	�;�Rd�}9I�ƟhC��һ�����v��}�Ws���8����޿Y7n��[�y�v�Ǆ����}*V�Jԓ��e�ڷ�R�b�V�d"tCwE�� ���z��m�
�oC��Ա�ѹ��i:��Á����Le�7�Ů  �"���\�lWu8�m*���bیs��Ж6�N+h=�u��w:�e���3 {�?�C�Ĕ��s2�ۮ=S5��AU!�������7�sV���}�B�.��*��Ř�u�Ȁ�/��]Ɓi�=k��E�&��������.ɭj���s.�]0�}�9���HX�i�8J�n���ޘsN쇙����c�l>�&�9=8�Yz���p�<|,�����0W1���on��x5AY�=�<��S�=X�b�����vC�3�_N�\��#s���<0^o�k^��v���lr�_ٴl��T�v��䚐:�V���v7�;PWS���[_ij���gLE�c2�޹�ц���d`_=\�5K����ki���B���8SC)�a���S��r�k�
�Zi�}�1�:�c�q8/:M��7���I���
�.O���L$mL��ҵ:t�Y;V���#݀�w�V�X��(�ymGew,ٙeVc-NV���-�R͇xR�r��ĺ`��^���>Թ�P��zF�����Y���������)����Y;���"Q�]�K1�ь22w]�n���$j"�K���aE!$4d-�h޻��n��Q�V	3w.�Q$9���c�ޚ�b,QDXĚ)���%$��I�BPc!(�h0����2b�BDPPH�MvV�(��PbMa,3EDEJ�t�h��A5IbA�q� �Z(��=wѨ����nnp16��k���!&(����I(�]ѴF�mD2��2ޛ�)��X�K6��$���!����ʤ51s�A�H���ۅI�d��Ȃ�W6�ѱ�M�D���2H����;��n^���ޝ���ￋ��G��i;�����ho�=��&�.gy�^�����X���1�� �k]����i�2p�`6�K7FV���=n:kr_Ŵ(�Q(��
i��� >�&��g��ӹ��r�*e�iwf�<�����hZ�R�u1������zLW5
,#�?�u�v��*-<����p{SZ��t�����:}��hGa����0V�Z�5�4��5m��Mms��#eoa�@/��s;G�-"+�+�܍d�z����\f��Ҙ����ܺb�t.��,�������9��l�w�C@.9�'Y����s��J�(���5�j8Oá3BћP]�)�A�1��Z���x46E;�gܘ4�	��c$�,���۸0����;���nn/[�Z՜�,��� Ũr�QFu��f�V@�t�9���q�Z�=PF%Z�E�Iސ��yLb{`lMmV6���oA	���	�̭�����;��G;�u�j- �i�v�G��PfC�R�Jq�ħi]:şs��c�yN�Z�R�yUݾe��1���j������YQ��W� ��(R�u�xIڅ�p��ŷ�$���n�TM�r��Boz�v�K��8�ئoM�N7����p��2�/�����f
n�>�n+�"ŵu��&���*Qe*���0/�WjW+�{��̗(��f��F��������.�܂+X��Z;sEѺ�ZQ��֠&n�#	�(�썛湜��o�c���e�î��sU�җNDP���웟�������d����~^b��I}�]>,�8^����xa� ��l9	�:�!��l�i��}�>��#��ͧkS<ߵ�V賎nK���ٮzw�~yp�Ѓ��%�9���I�zWݝ�����1�S�I�ʺl4�U���Z�E�ʒƥ�aI�ݚ ��lc׌�
Sr�M�z�U`\���@L��<�n���m�o�O�������Q�:1~1�F��-ɯ�6�K����0r��	�tm��BՇR��Xeҵ���U3=�g3.��m�}�%�]�^/a�I}�A�ġ�k�?/T؏���h)P4�Y�gL%�� �����5�l0;IT�5�e�Pg8dK�ƈL#ν3���bt.��r��n!�7��v3Fy�bK�0���b!��Ƈ@�r�.���3�0�
8ۂ�6�%#�)4G��:��o�=z.�r��#L�C�*(��O���\�Os���o5Y�1��:�cݑ�N��! D"��@N��{Qx�כ��l$Z��諐�y^k|�M���8���)�Za�j�W�y������/j��2c�ѐ�Ocx��*���/��ݙLd�?e�q����$�N��Q�<�jv�mg���k��]�{'�b�ar��x^�2gY���u�珯���[���Gp̣�]���4�T�.��j�YW���� ��=�x{ͼ���si}o<C��S< ��ĸz���U��3M�\�.s��"�(Q�z�򹱎�S56�u�f�b�Y�/�n�"����p��`hG;-�d�mT�5�%6���Zpwr�D��;���A?O,T����$����F�E�����N*1��p&���/8�|&�3/i�;woe��F��1)͎2�&��*`D�
�{^��=|w�!�ǘt��v�s0��Ro3��.I�x�Ct;ا٦e'Y�]zi�:q��.����\ �s	�_[wt��h�U'j�5fa�I��^�a8D[f���1I��R���LV��wQ�\�4�	��g꜐������7ϰ�8Ѕ�74�"u	�	�a�la��*���z�ƋO�S�3|6�=^�3��fo���z�7�5ƈi|O�����^:gσ��&��6��a9B�8�0�N���;�lV�h��QOR��.u�+�@/n;`8A���7G�8u��'f�TAidR�j����U{3���g]�ȰCsg��r^�υ(���;@s�O�
��'�����~>8����!i���~�y���
���s���k����-�p�#9���ؕ`�Y�鑯#?�-�u��J���Iɻ.�>#L�I�5�^��ˏ�}܍�Ęˊ���6��W��iw,�ViꝪJ3+��]�숵5ů7-�*�v���4Ɋ��������u��"	����K���llAT�ߙGS�(�[��3�GnY�z�p�fp0#�QVUڭ���,��zg��7'�¾u%�{����l�m�/����/��"�#���M�b��!؄F��4�ͬ)]��F�7zY�t�N��S.�,"îp��ƽ㥽!����
]t���ꆜ8��N�ƺ&�vސ�M��z�c�TEC�xĳǐ���c�v�I�z/��`��Q2�����,�g���vɽ���+Ϛ������X���N��!:g��s�~���4��(�z��y����ջЙ����e^&�(�se�U��?��J�,�a~��ӄ�Gz,SÜx�W���^�sN��eLt�������Pd��i=���XP=�Bޭ�[�y/]٥��oV��S�|g�*a�	��+$�7;��o(�E������n�oqa�E~I��B�{n�n�){{�Δ���
HQ%ٲ��0U|$>��%��)�|1�^�ƁF�[q�vt��P�;S�4��؃,����
���m����3n8>=J�|1���y��·�Ƽ[c�����8*Ylb��w	���S���V>�f��f��6��.�1N�N���%L���D�D�ܐ�ny�x�{����]�w�1�d�BwN`P��5:3�o��T��<�c[�2S�:�i؛iO�f�R�������������>��-f����3�|:�����j�Ȳ����찋a!b6���nΊi/�T���<5���*����=J;��C�{��H%�qyH�0����c!��i�9�F�2�w\�-j��k̸�����n[f����M��j��⣹�'�q��H�����k�ej������s��6T��M����RsbL�ePM[]��WyAlԥ[́[>��e�(l[�6ϵ�w�f��(6P�msW������Z��;'I�z�hg*�Ba��1�������g����+����$�����;��;t�@��xAb����Ӱ������I86s4�ZBA��p���n�{����6wB�^��n[����v|����H���nvF�V7�?<��:��֙I��E�hõ9e;!�,��	��tE��9����{A�4h��D�N�l�o������Z���d�T�������R�i�oI�j�S��R&a��Z��E<�.�0��C���-��S���c.j�SW>�y�Z؜��fb�
�A�1���6ʀ�Ο�]� ej�4�u\����x�;pg��s.�y�JX���B��Y�޵PEk;3٢�*E+���趗�I�u��+Ca���0%�͹�9��˲I<��t��6�����Պ�aR���v���J7�
l�w���c�d)P��:[ݳ�s傄��W�����ō�3��~���ϡ��+��PFǶ����7���׆OAd	cEw��<?S�Uϑؔ�������&�ò�D? �3:͈�q�&'��.�d�.z�e�~����D�j-�J��QE���%��0�C���T\?W�1�="zf�����^�7	���-C�$�c�t������X*�ֈGyu>_�*��]�6m��ȶ�C��|k� _��|��*�ֿS��oa��/f����{w�2���c��&*��"�ג�@�t�zw�xg�O�d{k�!?^I3�z0��VZ�Zո�����N�fyF)�9E�sJ��4�O>��?<�{b%i����y��xܛ�ӕ��B��!�k�آ��&��,�L+2<�j��IcA�a)�ݛ�m�YN�z�zkK�m��O����b�!2w�_�W:�&�Y�bN8�ϓ-t�)�U�&in���GwY\W,�Qa����Ö��@ni&5���C8еaԬq�t�xj�K�e2m�3q���?f���	��q@�皹��s9���3!��B�sɿ�>��U�# �pw~���sاg��ĸ���u���O����Q��K�6�I�fTJ�Y�oK�v���]FV�[�����g�2�,�,������7���4\�s�uȳ���R�(dD�	�Ս�����YR:3s[p���$n�K��
N������믾���M��������B��٬r]�3��kz��X1���2%� �`<h����ߕ��鸥m����[��K��;�s^յ�(���L3v>�:��g/���	��崅Z��5��zt���y�ʌeݽN��쇜� ��
��J=0���\�OJq'Y�Ӈ�9a�5��̴l	����$Fd��5�my���f�A�� ^�W!
��E��n!X�#�,�ZoԻ�{R��P��[���
����ل$��"i�^�{}�R�ԹH\�]\���ܛ{���l�s��B���u���H���5�L�:lk�	��#��Z��K=�Rť���b��&3+�Gd��T�{6G1XdJ~��B���cռ55���b�S�!��b�$)�M����"s]GI��^!���-AA�XbS��0LB��Z�V���u�I����G�#4h��J�oZ��f�v�¬0�4s�| !#�פi�I��d�`�cIL+ϱ|��a;:�G�p��]0�s��Z�^�a�d���О�J��H�^�I�E��酎U(��x�4������޶�C�r�2j�i�~�n`���A��n�;�VYx �׽
O�zc�
��+@���˻@��<*�O�gC0�x���> q�89ǥ�2xo��v{�a
��ϥ�|�u-�,9�R�ȟL�w�r=�J��pd�^�⧃J��2|���_O��ϟ����[m��6ڢ6��m�m�ZصW������{���_?�~�_2�����p�Ђ�li� �T�ư�
60�{�r���='ֽԊ�k���ۜ�e�Φ;�����L�C��v찏w�6�E{��u�MW���Մ�����f��֫�w��ʡ���eH�~ _9jp���!���0e��;4ڦ�6���g��u�-Y��l�*in~ٶ��2�)�z�4��A��m��l��0g��<A��u�qйb�[
�α�;t�i�Mό����g��9R��Q��|�ӏ^�3�@�f5�ؗ�t���lȊ�j�-���X6|�" ӻB|���t�C6C�Ⱦ�_��zHz�"o�g���,n�s�u��X$���N֪%�Ck
>'
,�	��t��rsk)z� �F�:�lv�ۥ�o���2�-�<�5Վ���>�1�����9�i���5��7zY���������u�>��l.��`\dÇ�/&���xiזx��斐�����l��5>��&�XX-h��y�؍���:�ם���A��lP(�͊O�ǫxU�N�=�ŵ�E����k���xv�lC3KTe�]龹�9�M�:%�鲋G�RBB�)F��:�4�P��"����0��;�,���K-V�Z��T���2ET�3_>�J_�љ���[2XGQ�L���2�������gv6��h�MLt�&�&w�U�UUU��m�}��{�qΏl�9`��h]/�����Q^�7���c��ɨ�i=�]:�צr������8�E�-~�K�B��jd$�`!�*����yD�/`�4��MvF��Ef�FBp�Z��ѥ�q;9t_�H01<'j��S��|� �rK�'J��'V9H��l���֤Rk�yw=]����2�<����������}	D�lN�{���,�H9*H=J�x�nz�b�8Y�5����Yoz�dWPk�sQ1e�>G�|����Bm���ݝ�_xX�u/9�v��'A�{7���lcl?���e ��./#�f�D����������@�d��bO�,ͽ�ã��4�Sw4�c8ֵ�[(�ځ�a�}�^O��ûs�;C`p�-ۅm�k=�{M�|�B�u���Ȓ�D�Ơ����)?5�2m��)�*�f�طvm����F���j��4� �`˃�:א!غ/Bz�s��]�R�uy�k,{G�շ�1\�J�o:E�;j��)m7��?����0g?3��X��^��:}�3��i'1�`���=tl�?�.2��[�H���t���8���}е�8�w74J0���-L:+E�WGZt5�t걯�;�;]<R�������A�$=���\�9q�[��k_�j�`�t9��Ґ�J6��OK�IQ#oj`bS���qA؝������UW��_}�F�lkm���5��F�F��j�)��{��R߀�t�^ø�v}��~����K6C���h�0���r�{.�asz���ٮv*�h&:��{�n�odK� ���5��I�jcl�͗[؝���t�Qr��>��T�44��j*q�dLCh�ִ��y��CW�\>����6��K�����'��x��J�f�kP���ˠŊ�!�Fu�6/��v3���*�[FJ��9�Xѽ����h���|��z`��YA+��V6�[�A=�%�kY�ˮ����˫۷|Rn7TK�T�C�8fH(6"K���v�.�d���\��  ��(���M[{:�sqse���y��ڝ�aM@�N7K�:ˌg��C�A�k�xIڽ{ާg/�1�;dHx����Om�#{4��t2"y��"�UE8��Dgc��s��=>3�~O���,�t!������y嚾fA��Ɇ��*L���X�E�.4�N�|��� B
�^U��3��������̿:�a�c�a�,�*���$�Ͳ.���sO��++��O��O��o�������������~�_����}��O�=g�~��e�A�v��I=��2�N�.�8�l�Zi�`�s����7�.ŧp�o���(޻?7zѣB������\���ަ�`���f'�]��Ɋ��k� ǼIn�k�j��٢=~rѱ���%}sh+����|��Ā�ŗ`$�Li�,؞'C=ֱ�,כ�w��:K\��߭�W;w��q���ZaNu�Q��^�X�$إ��X�f��e���^.��3|��i:dən�4�6vJZ��ھ|���)�?BZ��EmsG������+���L};Q;���N�rY2�9j�Y8�.LH6�k���pJ���lX��rK�oe�ף9c��Jˋ6���M���P{�����o8�G)���]k�_|�6���v��Q'��f�53ou��T�b�N�r��mkf�n�"X��qh�)��1��f��)��-�]#��]��9�^M��n�>�m��������݊���5����ym wd/)t�k!����˃�p��^Xq�kkG:�<iq/7'i�#zv5Օ��vU��T땶;�mH:v"��c��싞���pg�ɢצ��㹥�����?�d��Բh�R�u����N]�*lӓ���唶;�z�/�W�M��.+ V��M&�N�3�{����c��'5�����������X�����-�Cw�����|��	Q������ݚk>x;NDhJ�W�L����F������C^��5��Z:����k�0��Y��x�F������Ҽ�J������us)�N�ܡ)�Z����D����@�zM�7���w1]�e`�^d��;���'N��4�uH�X��%��`���#��Qu<�@61���_m�����F�Ҹ�)��e�<�i��qvɗiz"��3\��������鼷�t�Y�r�BJ�S����I^��{}����5#Y����[MA�]��s\Ԕ���V'�$�4��8l/����/y$�qX��܊�h��V`z1NCF��Wt	��pkABnN3�{v�b[�y	���~�엥]��9nE�i��EX�ۺ �;��!��@�sCY�w��������a���;�X���Ԝo�2�a#C�;�У����V�������Yu'l<�3x�6�	�~�@��S��)��$G��t��^�C�)��$��{7���K��jV���)c�Ի�6B�7NS�Ҧ�+�b�4b����I�.oV�s�d]����y����Y�ã�0#��a�Rc�F�w�Dj�4%�.V(�{.��]� {d/6u(f�=��5����-Mw���3r��7x<R�L�R��T����,�Ӥ�1�,+˦̳û4��ďY��l�o�l�X�کx�uUG��W)j�����ݢ9O�E�gM�`�p6��z�\���ݍh��ܶ�pU��(aJ���flѐ���>��{{Sjw����1N�����~����
M&���
*-�-���$d�9�lY4�Ԅj(�wW+�
M�Pm�Ѳh��ۛQ��i"�H��AcE��*1cb��,c[F�6-F�A�b�2Z	2Q�j�DmE�F�ĭrƣI&�h-X�h�1���Qkk!�R[cZ���smt�$�1�[Tm��w[�"�E���MFجQ!DlE�NnlF"���5��U�9�� � �~�}�9�>��n��wo�J�du��jNyzzS�ْ�1XV�pB�ʘ���z=�$:�ή=O�|�(����������_3>��a�}�ـ}�kEZ6����kQj1�f���?<|N��
[�`pq�:y�OE'7�;t(��I�P9+�Z�\��~*K�Cv��*��N9l��>�(wfS�����)�-��7��u�Q/�Q%Qa^��̦u��V�N˝���מ��lO���ۇ�p������� (LjzG6��4-Xu+w4cS�)FZ&Ơ����1�ۼ�����P���O5��p½�<��� >'4'e�oer�bw6v�휣���d/��StM��f��0��z��^�9�"]�p0C�wv۶����\��T�֝��������$����v�|��;L�v�{��4�lh�l�����)��ጭ��t�,�HB�p�]���l]��v/"�y��A!��za�l��^74�c�M�\3uL�5!p��@�ӌ�fJO~��Ƕ�����	��f/E\�5�����L?l��~��~���\t0{K�����{��0�_l��3��*���.R=�8��]�1��3��}��a���N/%G�=oM��y�66)���ӂ`���yڗN�@?�B�`��T��K&ڞK��A>l�h��y���WZ��t�^LΡuE&2��o�f��H]�@#�Y�ՆY\ը��{�y��;���y��xT'	��̩˃�t��LN{������t�`%�;)D��]rs3on��F�tY�`����0R-��=rl]�_��}����X�6�k�Qm�m���� ��iMՠ�e��[~�'[[ܜ&G�a�I�vH��u�cռ4��;B-�!�=�c!��*n	e��_�P�6��2�R5t)�/	�x�LPR��FM��m�'�|wW�絒�w؛~Pr�i����uh>З��=|  v���ԫu��K$�=�Ƽ�����Ld�����#b%�V��/�l���" �]�������i;Ϭ�'L,r�E�{�)�+l�v�z��Wp��}�
W�~j����G��#�&��	��Уc'qUeWC�ͫ*�bm����M�|�����r]&���p�\>��y�kTp�n��.��f��XأeNe�����Y�5f� V�=Q��oԨw:�W>�����!��a��1(��/Y����~�z��v����Vn(*��zV�NKԹ����6�����t�q����ۈ��\�k5�/�l+�P�]4�C�ǯ^��WRcl���z-��kv��1a�v/3��R3��E�cƭ��������S�x�t��6C�ϯ�oqh���D�/>>o9_�*=��Ү#�~��K�wGj�����zFZ�D���4�>��x]��^��=�z��r��"����YON��w�˾�!S.�Ϛc�kUO?�T���6�r#���	G:��g��˻�j�����4ݢ���g;�"+��:ܮ��:�F)��-��ڿe�3[T��X�b�#Ufj�+��������皔��Y�<4�;����������L3i�F�؞��Kdf�0R�� �-D��9��E㍺�������꿢���b�n��}�ǃ�2;[$���{87�ss�v��>��W�q�yf�&iC2u�������p�{6���xi��#�Y�22���� �|Œ���mn���Cٓ8ի<��E�Rɶ�v���'��x[]�`qm�ڡ޽�k�(nQ�Zh).�\zHS8��]s~�(N��1�{
�u��|��x/�c�D�y6�3�/Ѫ���a�Bd$E��#!O6�B���%�{)M1�F�X�ŝ�?uG��R�N��q��_Z����S��'�%;6T�&
��D�I/])�|1�>���N[Y�s�w�h�ގ��5���]I��j9�ޡ��8�a��҆m���f
NJ�q�����T��O����t:"���7H�^�\Ú�	�/^���a��B=r!6����\�&r��M�����4�q���ޗ�<�P���zNI���<�������-��ύ���Oӕ��#�찴m4�9�Z�IS�ai��-zQ���T�P��=�u^�W6�r�p)ڮ0V*mu�OL��Wp�[v(<���m��Q��t��Ȋ�`��<�F{;�7���jX,W���������VN�r5u��j�Ǩ,rqK����UUyTV��h�(*ɍh��*MX��}}���߿?_��]���8<�7k�'�i��ֻe��#XÔ�Κ�Ɵ��;s�;�2� ����r���գ��q���U]b��ǣ�[^�I���6�b��TC3{E��a��Ы�9�y�x^ߚD��d��������z�����4-[�L:��5�=�z}��2L���y�Wz��;q��|����,D0-+���a�|�/�p���;��E�Bl����_����8�׷D��(���LZ���s�<������zvF�L�R����\w"����r�DȔ��v�q�b��>?2 ��~U�Z~��D��h��Y5�L9Gb�ɛ�-]�+��.-�>�Ǯz�i���S��PD�5��'�y��["��D�o{9]����u�N�,�����{VlN5Z����,UB��:�^͛e��6��ɥ�(,��{���փ��I�!	��0A/0��L�k(%��m�oA	��;0iA=�9X�����Ǖ��1~z9��������VT\:����8��Iq�����M�2=?B����{���G���ߋ�@�,K󞾋�^�6`/��Wz�gw��嬡������~o�������/�����w;L�YQ315k��YzP��۸�o��J8���#�S5v�!���t+��&z���=T{_Q��q� Æ���Ũ��n^c�e����Q�g��2v�;�ݻBm�o�vh��ĀH'�%��E���X��Q�ME��LF�0 +�n���}�'������8���\c<�-�Pe��]�$���F��30Z�'�5#r�&����9�W[K�1��)P�`*��]�ٶ�ȶ�]8މF4�t��8i�5;1xy�!F�cFY���fA�v)��i�I� ^b�sȢ���׃�[�G�tdO��p۞0��q.��[��"��v�_����|.!��*���jRy�f�X^<9�-/#N����Qm���uMe����9�Y��52�wd���M����
7�4�U�����/6T�7# t�M[[�ɅHJl����-s��oÖRD�%k�g���� &��=ήMг`��.�%Q`�o��d�(�˅��
��zm�=�}jΌp�.1������LrzG6׈��-0�x�FtL���E�����qX���PK�\�E��'���FsF�c�3!�Y�jur�M��{a������\���*���=�a�v���z��^�90!އ��lk����b��!�M��xo��+`�#����v)Ս�v�$�%㝻��q��i��~~܀�>�}���H`�(<����I�w�����Ϻl�$�\Z�O7�
T1�o�����W�&�]��w�U���zǁ;�+ҟ�����Q�= ��Y���5l���P�SA
���IGKX}-���^]MK��Ϳc�i
U���Q7�l���_T2+����몺��lŴ�h�����foy��oy���f\jiw��"<�yO�(F�����/�y�4�$=�醘��<��a��R�B�M�/v6�+�o��5�P$�����l�Ľ[�w�as�A�z� _.�����C��.}zv!B�O�\e:n��s��x��Xt�H��������誩kjÛ�/��"�+֖͍+{w��u�W�e
6Up���=s9�>��Z��9n���6l�ǩ�[l��u�nc��K&�"Sm� �H��$Q�u��흠[H��{J�
�S8�Tu�B�=C�!Y� �;�WB�Xc�YR�&��B�"�����	�ś�ڇ�e-�p^�:5F(w�ñ�:!��	��@"}�k�bu��Y'Y�Ƽ��|�M�ݙ��d�sU�ჺ�saL�O�0���	
�DB`��zcB����w����E���?I�wg��KF���-ܹ��L1J:��p�����A;65�M��n�2��̊ʧ�ަZ�j�]�ʡн�/�S�+c���N%Ýp�~a�`鵦8F�T��u^*�vzj�:�~gX�/w�y�y#ُv
����
j6�<�r��P�y�-��#m��a^�Q=�c{���P��j��J7�.��V�IS`���?��u��J/P�MI�3r^7C��0��s70t�bf�`;h�.J<�yw�{���}{�w�߿ϯ�����Sh ���>��>���\�`�߿��K���������)a͛�"���?֣���*�^Y��������&���C�,3]���F/vWU������1�V!*��L�{*	{��Q� �K6���!�A&��3e�]̋����Aֈ:���Ld;n=^��U&6�:�-����c��0��jƤ�06��+wv�L��0����>jj�+�����l쾔_�?���D�9s��7l�2(���tM^�ͱ��	^�-̀6!�Ϻ%�X@��\O�T�{���`�A�l�.���� }�'=M�X�_��/��hwP�;�3��-��kt�P�(��?g��C�$���{2�|�a�}k���Ң�-�5e��f���èt���p��^ͧ�y����,�b9��	�-�G�'�Sx���J{H��e���z؋eȺ�n�2�%�L�!�l�zǫxT:E;�s�[�+Қ[2�e#ӳ��)�7s��)Ucoj+�7���|�M^X���Fk�?W�r�߶�(����7k�Iyj��>;��a���;�"�y���A�����N4r�d^�Ji����nk����@���0�I���㘶\��a-�Q�vK�� �W���x�h��d�~�y���WX�_I��6Gі�L���ODX�Wfԗ3��WY\�ّ�Y��Q<��FJ�צ�I��n7P���z����Ѝu�C
������|{�������m�&Ѵm��<���M�rZ2�m�Z��Gc�W=���=�ă$(���@K�`��7�Iz�%:Nޖ�v:0�e�.�=O�a�M�Q���s�O�p�� f��JY�682�a�`��F®�OzBݯ#.+&����"����(�a�y띭��C�	ق�Ȅ�q=�Eq�h�K�:��V���n)���.�ft=b��
.W'���ae�@��ь�"�Ӹ���'ލ�6k��d!�N$FD�Os�4�u�nZ���BԍcEGs�|w>%ݶ�����oB��)�D�wk��l�����B/P쟍zr�s���Ơ�����I���o7J}ϊ��΃��wv���w�\��7Sӻ1.���?0�C�y�mt^������V�S��5�w�g�L��h��Vj����^�w�':�C�l/�Ph��+C�<yLZ}���Nç��"9�b�E�N�hR��c���můk��!�f�1\�_��b��3��~gn�D��4�c^�mT�x�{�B� {+u	bV�x?<�u	�]�÷1�C�:"���x5�%�!��홽�f	�s`'.���K�>�gEj=�[簻��]�v��E��o�X�uj�)]5��X�0���.�,����r1]���*�4������V��r�
c�����Yi����r��q<	�h����#�六ӵ]b�j���2�)q�����&�6*f�c%~~���]����_jC,o���N�ӳ�������i�k�d�8�5L�M�����6�o	n]���D��=��{i�5	w^Ѱ&GL =Ų/bj��ٯ�kN�p�� Ũr�QFu���V����ct�FFM
�溦4���zw�V0hI�C�0���M�EcR�A?5��O5��Y뻔C4�P�f�Y�+���kkY��|j*.׮3��\��Iq�1<�5�=��O[,N_Y�kE��D5Y�E��i�JĪ,)��ra������N�7���N2�b5�pj���n��e�V�>ʽ�L�!�<�Ԣ$�����(*��]�ٶN�4+u�!�V�_]��/�|.�koD*��z*81����6�����J�,/1W�"��\hӅٲ�9�zp��۳�~��~彽V�X����BzB�	eeK���W)�E��X�/#���lvQ),=t������V�4;����;�9y󇶏-y��z�E��'@�I�P9+�Z���^Q�p��r�z���	y5z>��g�۴ȟx�%���(|m�[��n/�z+�X�t,ى8��T�>��ݓ-���=[��Y���Q��:f����M�x�]�/�7��I�=8@u���	ɓϬ@2&a�{�Լ}=2yb�i~7F�nw�A=���e,ݘ�Dա��u��s.���ÃU�hSY++1۸����l����0�����?����꾺���ﮭi��==��Ƙ~�%�ߩV���A���H ��Zx	�O���tv��{K1�i�/8�a}�HO �N8����ze�Q�$9a�+Z�>~�����(xk�w��oC�9O�]��uAat?)�vJ�Ra�XR�m=����f��5-�G�Yz�{���v}Gf%�����W�m�݌A�XC�+}��d]fö�a�,+�ėj�2����fN��#"���&YQ��3۪yw��`L�#ϡ�>0�ۜdw��w�"�y��A!�Q��B����ct�:�4����V���x��j����?~B<���;?a���� ��܄���ge}����k����n����C��5�K��z�]�g����I����y�ƞ2�Af� �-}����c /:Gsߎ��Zl�F�Ty����%�Mz��O���?�J��w�����(U�6՞f=؅e��+fa����M�9HL��
O~��B��נ1��E<z�Nȍ�or�u��T5`���	���}^A�v)�=(Rd�t�JSԥ*~���^�g�����x���?�������������;�O�a@��XmՆ��uw>9�G��5Z��m�f�QG�NU�gRK�w6]wZkx���7\�^�o-�1�6Q�ÿ�>>�d�-����YgI�uW!���z�35�u���yv%���WY���'k��W<�CZ���ۀ���הV��Cx{˖��H5�ݞۿ���p1���R���>�TNf�Wh����IBd�	�j��swH[��]���'VQ��A���W�T�y�¢�,�v��7C�c����������a�g��#`�<7%8w'����.C�g��tq�]!�:�]*��>,��z�=8&��!�X8��S%"j��h.x��]u�}*�>��w���Z�xh%2��d}T��!(���7[De\�C��C4�brsIG�,K����r��N��\������I��Pή`�TɜL�<	�?{�d;��EdsM#ԗz|����[�3�UݩJ[��~�0��r���+���'�����K�C�h���K$�$�ۻ�-%۬�7|�����]�Ű��R�zk7[�!FT����9AP�\�f�ɑ��QΊ�\3�P焽7�xA*�9�����)�� �w��(�Q��g��Ӭ�<e��pj���!��!ÙUv\XUt��Q�P�	z��*�(������0���������f�Ǳ�5zl�ԇno��u �����xb���b��'{ōY/�z!��s�����^d����Vo�:�҆H#>����q�yx�J=�}�5Ŵ:N�Gе�����d�r�3��l���"�c1�C��eq�7�r�X�D�J��{��,��0�;��4�^��#}n`�Ρm��7������џV� ����<���B�[�Kf\�y��ed�Z̋a;��z��X��.Yo��p�)!1I"
Z��wu��X��=�a�:�y���}�";�7y�c�&�C��9
�sLXw^F@���_8�M�������9��d;7�n�S2k�t�,e�iJ.��\�x�Pd�V�3��gۆQ���G;�����y����Ws|=�H<D��ÃG��j|{�n��%���<t��#<'jcF�w���w�I=�R"�ӔM�{��X�d�5PshS<#�Ù!Β*y�t8wf9�n6'��d�SMۧ�畸���mg<s�M�f�,��#�2��p)s�5SRĨ��ԾG�)}��<Ԃ5<ެ��~^!�%���K:�B�ynzO>/� D:0^ǭL��x0=V/n�q��g�R�52R�1,A٣�7��݇O/pL�;8�b;�;��R���3�U꭬��Z�zf����.�Q
�����pC�wK0ㅝGuK~��� �FEFW=#G���A�.�.�=�O����kku����+�=�}��zw���������߿^�ׯ�_?KF-�j(�4j�6����#����6L'5�wv-3Ii�sF�cF�7K����NvѮ\�Qc�Y�cEF4�Nnj#wu�뻭���(����\�TN��[��a7"�͍�`��Q�k�'9���Ȩ���9����2j��&��͎c*�ƹ[�r�.�\�ͮQ�+"[��cI]�[Inmnm�Ԗ�9\�6�؋PFلmΘ�h+Q�G*�b9��-�t�Qn[��ED[��AA�ѬF��1���r�-zZwlV��r�˚ܶ��1m����}�1$�O�
ΥS^qx�!��o����N��U�7�Y�nڢ����v����f;M6;3{��`��}�U~�0?	�)ٍ��~҂;�XK��g�gw�~yl��.�$.�h�N�O�9���П�|�x'��v�3):�]��:�x�3�����L�Mm��s��A�/\W��c^��ց!C6LB`��zc@a%P�I�l�'L,p�ܖ,��G8�9�;}��������T7Q��-N����@AC64�M�=!1���Q��35�1fno������~<wQ����C��q9l���a��8� ����@6��#[�A��Tm��Eda���j��ɶ�aYBV�����w=,��ip����:9��L�6mø%y ��|�ɦ*��&�N����{�PKܽҎi�Y��^���n+�zޱ*�>���22��^���>;����S#Rc~eO�Ǣ�x��GV_eQX1L/�5sɛ}9�I���3��d����y��]��ٟ46о�_l�zHz�c,���+�x�A�����{��-�6!�$tK� ���xFÇ�_=;��F�����/5���.�E�2�7�����i�[�v"����	��-,���z�'>o8��ʊ��0g�Fz̻֛9�ڂޕ5i�`ݦ3��gD���L��]��2�jv5�txa��V�x�5x��j��˼��v,��ޥS���.]%�沛r��q�z,�VsCw��nfc�m)�ҋ7�W�B˺/rr���e:��bN�,[�G_t����$�95s��[��49�p�4����7YYA�C��ٲ��6���yg��-Ҹjƾ䮟�	v�.{dB,��\�������\T�jeK"�����h����~`���T���X�lvj��D\zH��=X�,ڊ��)��)A�R�~�O�_O0�/;r��1��л�2L��N�k���[�y'�K��Hy]���\�3�PN,������ɞBEa0Ճ����y��~�,49Y~Tm+��d����B^W�A�$���v�v��"\�[h���t�{�[%Ω�c�Mmb6皟"���@.�mP��mzvx2-���5��$ޙ{β����:��%�԰�7g���RS��E#�d:��\Ú��/^����[A�T����Gd[�Go����!�{�R{�¥�l�n�E�?"�A/ZT���`y���[E�V�k�	�o�t�,/����s�ǆ:�	�n��Z�~;(�թ������; �ʡ����H3t�ʽe����]���|�H`�ٓ��OP��B�FE5�Vצ}b16�^N	W��u�ΩJ���y�V��$�<���F��|ʋ5=��w��\
hߡW
Y ;Y_�{���>���Tt��jy��!*�]����џ�����: ��Q��dugNA�yJ��k%6q�u�Qu��m"4��0�.m��y�/�x��h~{�ۙ�A�T���/|L�u�ve#��~a?�v�E�OC��Om��?]<�]��Lg����Y�?z޺�}[bTW5���������x"v�����t�w�B�5�]��SK;��i'���0$8��8���׍yXH>L��5�����W�o�ڽ]Q�pvߐ�#~ޠ���9�&�3Eی;�Lq'DYz�tT<���Ib�+�l���lx;.9��IՉ���u�ޟ@��L�^�'����A�ș��}kOzoe��aSU�M��H��2�J़9C�xC
ݟy\��W^k�43�H8�0�������6\�d\ū��]�NvC��Xγf�k [9~iw�a@�!'�|Ǧ"nA7쨬j]'�)��!Z�"Ҋ��o������b����k9~��T\9�\d��>O�NF���O㙋W��|���c2���tv��OpCn?'��4)X�E��ypy=i��A���}���}�1�Rg�lz4�Vʲ�%�0���Bd���rWH�g}\_�ؤΰ�ȶ��Ӎ��}����>�H��u��m��pUnN��I��rw�.ʔ_|hL�.�ݑ��~O�U�O�����S��=۾����܉q3:��^�8�'Lӽ\������I���}�)NK	����/��]����R�Jm �T��;X`.hDcu՗�5/w���'��89y�ɝ��nCml3po��HiRe�����<�/Iq�l���;t����Ǡf��uo^���n Dc;����/X`K*��}��'���E��9����,楫i*�8�n��u�����f�}u�lC��Cs{��������
8O�0�پyn�՚���m�˸6Sq��V�{� ��0����������:nw	��s�:"Mв�cLTK˺1Q�dMbg�'��ޢ��G2�)V��y]q!�F�ZA�����?���ENk8�#&+0m�m�%��B͹��:���k��4'��hN�5~�:�k�\]C����U=#��tos�oe�~��v[YԘsPi�kf��q�nj�FC׋�g8`择3�%�V`�w���w@h�C��+�	�v)��K�a�,	x�c�]�^��h�k���-����n�A�W�}�����^]� `N���О�lm�29�N�/"�y��A!��^n2\ݐ��Z��x�ry_K���-��)Ꮈf�\G"ˉ�����b{8�3����|~���w%�ǜ��K��q���_�ց�kT�(��lW3��ѳ:��|���dpU�d����XA�wX�����{������n��ʬ��B�ӑY��t�wٹ�������S�U����ٓ;[E���g��������e�OT�hK�v�A�}�4`���ezQb��&�N���zd	�	��PB��ךE�S����u^�x����I��D��3�߲��8�|SkL>ŝ�C��YU-mZ���rvPeanP�~�G�=ysX�!�tK<h���k}|�Ŵ�{�9�â�Av[�pکnnr!6h�!2�,T)=�Wm�Ӻ��V���І���0�����s�d�hQl�G̘	����y��	L��bS��RX&�BJ��x��֎�2���U�W�/`���{�[��6��(���]��z�������L��x�,e�0T>�k�9
��;W4��I�>��{�����3d�!0\��C�*��N��=\�~�sJZ�OmHߗ�XY�<���[��6�� c��Pw��P͍1�tt�e�,�+˺|x�l
����Co������qV��?Qi���,h.��5�\<x��a�2mk�iXU�[m^��-�]N��HM�'��	��NP���ը�s7�J�sז@������ڣTl)��60��V�1y��0d�~��mW=E��Ql5�J�{�~1��|�h����BI�9�g�7c��3��oj��5�ǖ�<٦���T9*XaC��V{i��������E�a�*�_s٥-��#j���yѤ�c��<�@c�J j�b�����T3`��+Q�#{�<R��G����U�Ql�}�ƌzUc9Xd�?����^pz����㡃�B�ȇmt�ۏB���X��1�2���ϧ�c�x�
��ۜYΩ���6�1a����f~ƈE�����[.��ے�}}(�@D���cf1=�Tp�l[1٭���f��b� �b�:�;�x9a��Se�N�k��߮#��АF��蹭���e������L"�$@"|OT4�_E��b*���ZZ@C �����Ÿ�,�����]ع�]Mŧ�ޕ��#{U3MfSA+��#&=��i>yǆ�yg�ކUY����%�'�gv�n*����B22���j}<���2䥛{��dS�Q�Y�i��͈X�u��gG�Y"���a�;��8Z��	l��7����d�b�O��:��M��k��n�V��x��O��X����2}��.Ǽ��ܕ\�:!�U����sN^=Pc¹o,j�Y�i�#)��-��r�cD<�V�y���D���?U���[���,�h��sq)��v]�ۡq_Kሔ�ƩƊ4���ny�ϑp�<�3[H��
~?h���?�~�3��xE9(F��=�������X�v5����~{_����J����g2��Ҕ���\�\�ϽJ쳴���a�Ý�]�1e�S��
��m�+ �^,H�W(6�62@���X�9Ǐ:@}i˜1��E�ʘ��IBg�B\]�c��-o�9C6Y�����tҤ���r���X��sP&,�>G�g�"�5��K�^mG����ȄƧeTt�R{�.�,�n���Z~XH%�J�Ԍ����3DD�ů�r�ufb�l���C��$FĲ�=sM��q��^<�K�9���q����lQ��K6���R�P�1TK�k�;
l�?s�;'�^��\��&E1�dյ鄟�<����\���'=�?��w����l��_n~m��$
���� �^�;s��'����q�j�d��q�5��2�hs����a+͑���	��m�LW5x�XH�P�n�����tŬC�a{�C�k�"�+;��k�'�(fu5�4��i��
$@�8�sQ~娽�q�}�����3�~A�MF�P���Lrss�5��oP~y��@��>��2�ZI���,�9��KnJ����9Yʨ� ���!���i����ә��s�s輳L�Zd�Ql�#����K3�	L&Awɶ�t��j���֥������H<3�D�r�ӳ6+Z��(Y��y�J��c+�Mud���Xx�U/�y�m�:sӜ�	.Tk9�Y#�)
\v��̰�L�8��eE��+-�WZyl��T��٧�n3���J�T��c9�A'g�^=n|�=���tp��*Y�LZ|mV��J���x�K��侥��<=���K^�{Rh\�<�E�����g�ٶU�/��{w�`���|��za^���ʊ��;K7&�W1��F㺈��Cv8��%�Fq�@1��Օh\g�
ȱ\e	��k
�]hU(=����swwu�n�,Y��:u2Ǳ�):��Х~�E�5�8���^�+��6���	��$�.�S�����B^9;U��!7�X��L��xNx�B��U��6m���Џ>�W�p/\�ƽ^moE�o 0��q F���f!�v��i�I��c�E���7�)h������۶�V�ʙt��Ï�!"1��BzA�TT�5(��)�u��Xj�Yʺc�|jd�v�p���YO!W��sם���mD8Z�!�n�yNvMУ�S	��ӵ�V<�!�Mw��w��9�F�Z����x�,i�ߐ��D�LkL�~O�����U:+�Z1C'�:�,/y��g=�wj��8��RX]<�eN��^�>�58}`����!��s^�l�����\�걫Z�����BՇR��Z~��eA/m	�ז�+�u6e]w��< �Ԣ�����V���OcY��/-�֟`��!����.G0�����qg޼B�{C��=;a���p@R�I���^,-��C�]�I[ԝw̨;��̕�-v�el��o����S�\���u ���H�$쓷��jʹ��V��):�7�;�gM��l����(-01�xN˷nt��0�@�	�kf��ƥ��zew�ӫ{FK�{ߕ�|���K-�@g��.�8����!0�<G[���ՃƝ�{�yE�]��e۵��<��!2�6'�Gfj�����[���C��`L�/0�>�c#����/G_+ '��kݩ�S�9�Oԍ�e:��{�0{C����-3��(`��W߃�q1�):���|l��um�[dC��4�*��<�_A�T��\e:n��u����9aBä�U�n�q�v4�kwf���lU��TkQ�������\�]D,�o�Q�@oM����s[�F�O;<���|�z�յ���^"`瞀�]�˧Yu�T�5xto���Td�Ȓ���3]�魏+����F�{qs��-Y�xd^��<A�iN%�p��}^!�sh~BS+c�YRX&�������>��������욐��d� 3�]y�t��3�範'݆�:fRu��3�/jEe��rw�5[��Mԑ����`Wq�U�Ky����~�C�P�%G��&����v�{��!�3^Sh��/�@
^���7�'�'�x�^$F�\W��S�[���Y|,�揫����y*�.@,�5]f��2ں'w�gLj�2e���3n��ijotp̜m7��/8�Ù�ngn9���x���<�{ݧ�l3��v�8s�k�Qw�y��ܪQu��Lh-�u�u��r��sǜ=2ٱ�GM�L9��&L��1U��p��C�ˡF�m(qT�]B�Z~k*]&��q.��>���nLՌ�<KnN����i���!7P��No�f��'(]�*�=Z��3b�祀@�^�< n�c1�lV��r�}�yH8C�c,z�Z�Bvi��Ijd�M�H��r���S9��E���v��2oe^�n���!�:�~/p�}ۏ^��V �Lọ��ְ�����5jT���^��_L�P]r̫�,3�.���s�y���;��6C��c�`�0!UUDt1Vs�q�sǥ��mq��)�uv9�.�1a^��\H�Se�jL<0�t�d8�_o�]/���6��4�0Hz�����H��T?W�%��塚�v��T�%�r�����He����z��^=�{z�4���l�c�gXu���dÇ�{6���o�g��P��⮥�v��gZ#ZZx(L��d���G>���.JY��A� �m�j ���o7o��~���~���{ߛ����{���W�>y���щ��u��v��r�jH�h��֟�J-�y� w�8iz Wjz��\�0־7��C��J�c���`Z�x������H�ѣo5�O�ߨX���~u7{��,�ѝ���%��
L\�sq�j�imCÓx\�[ؠ�p�굘:�>~�z���i�#��4dR����i狦��N4�A׈d�%����z�����]�U�I��:�����aA��~��A�����ҩ�nﯢu��u���x���(z���'Ց�2�������qy���+�raJ,��f���f�m ���խ�N����rGxn:�l�3d�s$�A��Hk3��棕vw���ٓ�G��v���d�9���Y��/p&Ηy���=�3A��5�����(g�zây������'MV�y���2�c��kFYH^v�+�
gZ�8���@J��4s�;U��=H�|�YyFjm�F5�O+�s�e��u��:�����T�{<&p���[�Ƴ��K���F��QiyS�2N$�1i��t(��B���2Q�^�:X�����M��Œ���[�3�R��ok�7ď^�L��1��l� ��b�uohU� �j&��N�_b��Q1���ڭu[��ө=Zm�Gi�ud�ܗ�8-��w�u��Nd��ʟ� �K�l��s{0ޗ�������IN�c|2��f�����"	#���F#�t��ΚYv�e�������wW��Hu�o�%�&xg4t=�9N�j��{�lGXU�2_��Z&�]�^��.������\��k��\���˱��<�K����a-E/:�����8�Z>�yO^(./&L�p٦�m9њN;�,wL���s��^:��|����he�9Q����1-�)b|*���+2��=g��5p���,9��,h�)r�=C�P�>����!��H���六֟��2������}�o�ݿ�6�k�7��(L�kq]u�˫(��uv�$�͸�2=�=�N���!ɾR{���f97E3cDC��ãjeX(^ޔ��X���ٮ��5Щ�A㛗�j�͎�wmX�:�4���(VvK@+���w���8�Օ����;�@��^u�pH[e[�uL�Y�RN�d��7����N�2.�BT.�V���]��9��NR���4�e��4M�얹�r��Yih.-���=�h]dN��+5��U��-�$�U�qBdݐ��}�4cnOb�;��1<=�p�?>�U�لb'!�(�C��U��d����3�1/��Q�.���{���-�}9�=�9�����[aq"��"�R�����O-�gs��I�J윈�[A�%(򽂡�A����Zñ�gm�a6�������ъK �:��:���m�w�˙�� ,o�2?l{�(t�1��H5~�g�#�h����rr�Y��S��QΜ�����In~���>��I�O�jMs\�&6�[�5���r��[�h��T��cG5sh،m��\�[.\Z�nX�h��ޗ�E���X�+�6�݊�T]-��G64[j�EW6�[����G+��+��Xڹm]wu����nk��.d��6���ۻ���-�F�ђ��snlTm�TA�j�ɨ�mi)�i4�&-�F"�Z���:*�6�RQ�mͷ5snV�llm�+k�X_�>?X�5�e���t\Ļݟ4�
d"Szڰ�"C;'�WU��ቕX����{�7�Q����I���?b�283���9z]�<��u����H2��N�[P�����dzM3*�a���W���ټ�O�rV�ʝh�*�p�b��~��4��+gXQ�{i����|wA8��33z��Ѕ�	�I�(d��0�sU�XR���.f�)½�n�)D�2�&���C���ȧ�dE�S�vk�}`�Nno;����k�u�U�]㜗F"S���Ɗ4���m�5>Eê�����S�����F�٬y��]"�3j��|�cfY��J�4�yZO�"��Ob�a�^+�q=��<���V��c�f���������(`���Am��A���6�_
�n�:/I��A/Ary�_�j�ȩ�����ͥ,��9�l��_���lK.{�����r�k�vQy�R5�=�c�GP�골�y��c1ܮ_Z�ƠK�@�F0��!8�䉋���V}�����z���o�������j:w\���ړo6�}5R͔6}7ͺ������v�E�z�{�:A[K�1���2��p���(��S�+}����6��a���"�`�����|?�}�|��]�n�{��#���2�-B�(5Z�Y70P�X�X�eun$�ٗ26���5���y�k�)w���
�\��%L�k�������P������S��[cě\�uw�V��Ŏ1��v�Y|{�!�d�f�,Pº�_��l����C���)ܹ�2#o���s4;x��h�[���w��.����:�YSj^HR}j.�+*	�s���;��pЂF�LIv�2�ZI�$e��<�x�)dp�Cv�*��Y"]�`q\&��I��N6۝���4�5�O;ʮ�G��	���y�o���/x�+�~��ƫt9��:�E;�N!��Ƚ�\���lV�P�q�\1�^z<�}��y`ke�۝\��=fͲ��-�<��}p�)����5���\�J�>����<G#9{�3=��Y^���w�('�' K+�Y��:��T\9�����X�/ᝥ½NnQn���ݠ.�ï�LŨd��?A��ܢ��ZhR�J���˃�٧��7�;���?��v�;?���᜼T7��3Z����/e���,[C�&I��NJ2))�.)�)�Ć���용SE�=��
:ޏHB1�C�&F�����COa�m2�2�^b��IwT;��V���Ymn��F�;G4������e�����B~��A{��YT�6jRy�?�:̩���2�j|SDGG,jg��o���y�8�Xsv`����3��;��$�n�y^37�}�O3��uyc�k�f��U��.�㝓7Y��7j��x�(��W1���hqs�{7Z|�@�{6�]�y��L&ky�l��:K`���v/���G��Y��vY$�2o!��j�<{51��j�%�r� ���!�Tk��*��ܛ�G-^@m��:6d�.�y��E����yk T"��IcH�C		���=�����CM��7�ӯ���N�{̛"���MS��гf%c��*�
��̦�V��'��^�\0g>�n�1v�:H��r�ؘ��2��P�+Ӳm�BՇR��X	�V��ޒ�mr��H;Bu�s�w�w��E�&�Z�K�{q���(ƕ"zׄ�-ΒÛ��@�~�Ǵa�v��������u��3;����*����n���~��@�xD&��br]�u���Qa@���%�f3>L�l˕�/�-��6��fA�ʺ���yw���24F�yO�(F��#���')Xةj��s0a��FC��F��� ��].���U�:����q��)<ƴ�d���p�3�x������u��r˺9��O����~*� ��6���M]1p��x������|��̉{�};!Ip��SI�UF5+ʩkj���`� �eȓ�Q�[�l$\�C���K�l\���v�r�پi����?/�y���$�Үp�Z�9�[�1��l�vv��*:��:�d�,u~�p��է��0&��� �Rhb	�7�0���';b�#��<;e�ʚɺApkq-	^���dT��$��;JK�2�9uJ��2���f�qg;�7�g��!5��0�a�'e���mT�5��%6�)	� �P��%vо�,��F�r�2�*kl$׻
u馞S�;B
-��Ġ�S! _W�i�S�A�	L���Jt��Z�
���>;t�M���Ӽ�d#uP�������z��;ćɒ�/ ��/�'�׷9��e���֕4,h����m�<���齃�)�$i0�ؾqOw0����X1�l��.z�C����dKV�"�{��Kwf�#����j(�ac�J.�s�1�����>t��?$=��A�_~��]����*��o6,vUӊ�Hʽ�=�sb�܂Ɔ�@+��P�ʮ��Qi���AcK���W�q.��pˌ��O��Ym�ww}���i���ǌ��+���'K35�k���c��V���ʑ���6����ݩ��"�ar�����Ÿp�F�R�ǡí~�٦�~����қa������O�iE3��7�cm�����YR���`�zCp���;k���v�z��5�V �ai��ٖ�Fɻ�׃��>��>�V����,�C2נ�ǜ3��x!ш��|/o/���J�^[��Aqaĝpm�?�'7ݯ�Y���D֊�G$]��:pq�16�D�����)�|�´m@C�s��+{����K�=;��w�A)˝����������]1d x,���t��>�uI��HK�,�]�Gv���{��4x�ڟŧ���~VJ/��<zHz$@��+�tE1jb���]�|Æ��\\�3�$N��q��ک��1_:����q��F�V0���	A�HB�42m��lEC�Ȗ{ō�ϴP|��ڶHӔhdB��l���^=����{n�����^](#&Z^ͧ��"�.I����/��wT��!O,��id��No�S��ٜ�˒�n��PeAd�֎���0�.�L+ݫ�b�/���Y�z��V�S��,:/".=<)Uc�mEz}�D�ھ}w��lE*O�Z��hӼ�5�oD렫�Xz��oV�^��N/�D��x�����3ɷ�/�c��5WL�F�eqk��(�E�Q,�t��"7��<����a�^e]��V�uv:�d��U��o���
��&ˊE�tD�X�b%9��E1�Q���#ny��.P��\M]��8��7!e�i�z
�c1�0�0G!C��J�|1���t�8��sq1e҉�fX�O-v��׽{ϋ�"�G�"=D&����:)�>��T�t�/�ŧ匤��O�ʓ�`/��3���A�g��g���<%2V���1�|�|=�����E"Uף�9���^{{�q�Rp��t��C��}����b��qs�˷�b�e��ֺ\4�t���;E����s�޼[�=7�T�d�L�Wn�����}��1s�������9l�����ji�y����)��p5���̹�z曬�[~v����Q~eQ%����5��7wb�.�/�s�	��t�����C`p�`��������W:�X�e��K�BbV�~��qıU���^#&�m\���6_�-ݛg��~a?vmt\�ڜL1�j(�:j�8#�_1<�S��0�%04�5���#�����@�������h~gA8�W��3T/��{�md!�"���t�Yʄua��	��C����^/�ܵ�#�$���5\$,�S�2���8Ɛ"c�{�^ӿ'�u]�o�i���r����'i<�1�v-���o5�=녔��m�9{8�������m�87�זe�t��j���&$F�U܊u�A�<�Ī���y���4��P|aoql�ؚ��u�حeL.��.LU:7���	Gudhb��Pb�c>�ٶT@�t��N��'$����n��;���C�uv�q��j��'泰�H71�WV�ю�ơ�j�3:
�?��2B�g�����O�g�G�<�vM��H�:�U�`1�ML�5w6��i���q;U&xTY�S�:'cDv���/��B�w�Q���3����}hIŽ^L5�}Jv'CyDǝFJBu�`���KӚ�њ�h�p�Gd2A7�k8V�y�2��W�{g�Ƀ�9�x`�a�3�.���MY0����-~O)���B�),%�\[w����@�ؔ�!�D��P믔��u���t�]/	;U�p��ŷ��$�b%9(ȤUQN-XX�2�⨾B�#�������oD�#a�$F�����Cv����&X�LV�E����]9ɸ����#�ׂ�T̰����.%��AƟD�O�= �����ʗk�|��v/�)���e�I��m�{:m�u��iy�m�\���ώ�<p����z��RreS��n��z���ZT���ևr��*��\���j��*KGjJxwf��|v����pv��^9��#�P��ө���箅�$㋱�QaV�y�ߩV�Mr[=�x�3v���xc��(���8�y���	�	�ϱ�hZ�J�i�V����'�Нe�I[{��-P�O9�����"<��(�p�\��-��E�5
��'3X�]�0�6�tg����ܥ���V:���dK�p0�L���s�쓫��������}�������U�2؋4If[�ޠ�������~9��k6�~R�����;�����/stF\�n���G�����y��;W4��.V��y�'��(-XY7pL9M\�F��������JѮ�V�E��sN)�s.����M��*~�Gv�2��}y�T=��{C��ŕ�5K� ��3���yO��&nq���u����r��vjv	��5�����%v\��lM�1���`0%��tK���f�RB���Z��Qi�:5��ym��9諐�"k�>��t�������K�4�G'�{�����,:N$E��=�F5m�T��.R=��R̡D�:��zm�O>m�jqf�ԝ�7[�*!�yg^BcH�1�>��	wig-���ނ%6��&K�N�%>�_�����߃���ާ�Ml`��O�흸����I�逐�}^!��O5?!)���r�=����[J����G��S�Δ��IP�2s����z�w�!Ŵy:A������B!�)�:�8����o/*��Ws��,���Li#I�y�b�Ľ��}ml�a�&!0\�:Y�S����{Zv�;b}I�E����E�x�4�����m��yO}����yx+��Z'�\j�3S("tl[&XnD��I�UYU��j-?5�����a��p�����һ�fd�i�ě��tUD���[U�J���i�M�G0P��9;L��:�=�`㈹��n�̍\}��++����ӧ��B�0v⿫ģ�p ˷�i#^��[o�^��T��&l��gu�њ��,�I%c�0������|�j�}i�Sjr^��]g߲�~�^���n�٤�ę��	��I����҅*�dghI��^�����q��_�"�^� >��a���Z�S�M�稵�t��j=+^����U}��Aȅ����~�z`���[�s�����h����"�r�A���A����(�����Rm���π�zfy��f4Xgc �ww����<��M�KXU�J����������n��C��V?Yxv`�C�u��q���LZ�X��0:%���������U���p�y��f�88�s�8�K�G�G�ќ��k�����O��ﭺ+��Tu��z9�������`��E㞱��ޡ�#73M_Ia�T�4#&=�Ow��s��2��[Eu��V][ͼ2^yh:!4z]źcNlMO�����5yrT��0���Dl��1J��z�9����
ek����'�z��]"���h���ǧ�yUc�^}�*��1�����rk��f�T܆l�bԱM'Sь4�ǫUi�Yİ~��08E�Ǽ�~�`�,	^�!~Lr+EN��A}|��&�~[ת��78'{Dɲ�FĒ����k+k�d������;\d�/t,�7���E����Ei���VSϷ�j
��#�ȫڼ{���:��l��n�����s����L��vq۽����;g�ow��L��N4r�d^�Ji��F�[���������Vײ�ÊSΰ��*��b���p�;4�x�
�𐄋�%�������"��e57f0���h~��N���B��WH��~z��]6}c��	��6؝���0ZJ�4Ҡ|1���(��\ÚߗL7k����T��V�ʙt�s!�[A�yЄ�Bvx7W��ڋ߰�v�M��#��K횉�c*_+�5wS���-א���0�zz:�	�X(֘r9ā˞�=sMל�Z��F�h�g��٨���t����>;��b]�:1��!�:C�y쟌t��Y�r�Ή1#:S��7s�%���k��NZ�6���n��ht[�7k�j��^�Ń8��]�t����z�7>S�;��0���a�Ʋ״z}[bLT����Hwn�����9H�%]S�{Ѡ�:���C��z���8ȎᆒpS�	;hq���nZ���%�۹��;���H~��Ƈe�s�M~��l�^�瑇:��&h�P�.ŸxO������x����o�����|�|}c��24e�F�p�0�+��o+���׶M0=wXuM��w�����^w�>짎����D1��!����n<��.�}j�$w�/Q����ݫ4��,>��% �}'r�#��3`�����G/�%������B���GOc՞
�����|6��}6�2���c;i�g	��wZ�Ʀ�R�M�s���˫��fD6V��������ڽ���|0I���۝���B�b}�8�x1��C��;F 2B�&��(�	���	b��1��)]ǩ�̨Y��ui�d�W�����H�cX�ER�ͅ�d]O��veIZ�9ݱ��v̼�%��bv���K�'-�B��8��n�9O�Fr�ɦMӎq��<k#u��D��P}���������A�)tiy��|C� ڽ���?1$��˳}��n(�<�ݞ�:u�T��V��� �܇RY�[+�ܸ�^u�lke҉�4ܷ{-�L�+j�服�M���]�5^\��ҭ�C^���a$/��櫸;#K��M�m�WD;�o>x�D��NU�LU����Av\�����gS��`cU�t������L}k��b<�&1����ax]cn�av�S_(k	V����6��ӽ�Y�A�f�����85NJ�.-Yj���@����t'a&�o�X�$�7���v�����812{v�ڲ�Wu�һ���R����[�	�ڟ�2<�uw�syf���1sg �Ϸ��S}�]}\5�v��ת��믯��b[-��B޺"����T���i��ݧĻ�e���Th�ݶ��R�7��I�5��Y����u�[f�_á���$m�}M��9Fh����f��woL����ξC@jf%�d���z�
����+z�����-�b@��{wc�(Fc�!�c���0�Տlf+�K����iVc���4�Nj�ڐޡ(��`�}}qC�b{-1����-یe�[ś��,�/ن7q�E�Npft�[���
PC�ݩ�N��],N����(5����%���T+ZV/9 Ok�Z�]��5�[m<k8�$_X���l���z�w{�E���p��b�ΐ
���.{�o0䱶mw=�ŽU���=�[��H�����ѻ$��z�7�g�׆��Y�%@{=�{ݚ���`���AX7�ΐw��s�$���^�������>�ƾ6"�E��P�����#����/c��k�Mf�P��;	��KV�:�y���.�L�3.�Tz]_b��R-�u�N���-ϵ�ls21�])͗!�6d��ia���[�fy�γ4�ַ=�2:A�3w�J�9�O��}�Պ���[��{��g.�_l,�u�46�lǣ��,�����p��5���2�ޯ���k���E?h���%���ټa]6xA�p�H��5�h��9�{a��s6�c��Y�v
�q9=��L~�4{�Y��n��N�����qX�:9s}J�`�t�Lӡv.R |��C�	��ձ�m��֋nZ�ڍ��[�Ti-\�櫛�wmȴj湣E�E-r��k�I�nk+�-ʹl[E���!j5�b�]ݶ�֋F��\��ʩݶ�Qh�[�D��+W,m\���[�Z��\�\�sZ����lX����6��k��}�����ש��^h�ꟶ��1T۟�s1�C����d[;)�"���R�5/^���0�˵#�gޝ�4t~ղ���zNu�Nh�'ʹ�o���#n�iP6RJ�=�����X7�Iw?�q���P򖟫`�?_`#�>���_��m�oH>i�ʦi�Y>L/�=R��������۲���hbLCm���k����D���~+vy_Ү}]�e���dN>����<�2 <W��X��AFu��l�*�Ξy���;X4$�h��TD�+����v�׶
'dq�2���t���;'��%�$�T��}�=�9�0_���ma¼��H�ݬ�45
DD�@LIv]ɴd�箈B]lG'��j�(�TXSP[���ihz�x\Ь�}<�rb�� ��(R�u/	;W��p�/�1f�L����(е��ʕ�wVqb��`��[�5Z��v;/�t��~�5��B�C*��COa�i�J�)SA��u����Z��Y��%�V<��O���/A�-ᄍ���>�!?T�׆��1���*Z"g1�F�-��ܝ���*m�u��sH[�#h��=;�?<�m8Z�Cw=�ůݶ/;J������{���]H�C:�
�2����/6T�4��@q>O.�ݎ����<�Ru�`)��e{��n��go[Λ��1��_߱������������#/zyō����>�G�������wgޫ.���W��[L�bW��<F��..�Z��lɨ]�Y{��2��Sj�F�G�{�2z�q�plڏ:;�5ˁGP�L�Nk�U���2��5���Mв^
�@�*谯Z��S`R�a!4�8POl���ߏ1S�55*39~����`鵤��m�2)2^�����kߊ�^�Ĩ�	�n�
Oӎ�f��f���i��U�MA�Q��Ѝ�h�����N˲��,9�
T��y����/6Y�*�ep=ɚJ��nj�Zr��"]�p0 �	�;�\�$�z��ύk�w\�][��s��V�nėj	K�k׸��I�ƀ��r�j���y�4<�5?,"�Uvc�eWf�u�{�i�C������W� ��8A�l;tE��tM�1�����/��!ԗj�z�%���!b�@�8B+�'�5�m~͍i��<����\�("k�"�i�WL\:]��q��ؼًՎ�T���82N..�ߪ����R��)���A� �(Q�Up���;7���M�/�l���¦*K�=��&��Y�?;`[8�XکnjJm�R-�f�rS��4M4����Bi����Ӻ��O~��v@���C�z`$&��Cv(�^o�}��\I��P����^�}�����X�E�������ݎ<u��n�{N���8�&r6G��u�Zgkю��TI�܎�0]��&,�5�_|���ߖ�u�M�P�N��G[}+8���	|���/wW��>�grv�;F�:��dwn���>�dO?YRX&t�����z_q�=z���[G�z�!����-��P���=Ϯ���W}^��Ju��YX9☤e0������OZ�������Sn�}���]���7�!m�O����0*c���Ƽ����r������:�k�[9�;��)k���Є�zBcCУ�S��*vj-?5��.�̳z�nL>5ܬӛQ�8u�P�%��8~L#�ͭ��>�h��.��0,p܊ �F^�Gs��b{hђ�
x�n�9��B����Ӈ�p�Dk�ã�*4-~��mQ�Z�(J���Rٵi�^�`Q����1���:�g��;ʈ]�� ��s	��Q���"����$�
!np�����X�G,B~���3�ǡ�g���cF,3�.����y���9.���+��[���}��w.Vl�m��%�Ǥ�$8�q��:"��Pwc��]ʀ�\EDh��:�m�p���!踘�7����h9��X�A�$=qhH$�4��o��y���B2��O��]K�5���W��,��������`V3�5y;.v4�Z�n��^�9*Ž�z��_���Cݹ[S]�=�8�E[�6����H9�4H��f��yx�C�/ݻ�w�&�mγF�yQ����z�=�a�m]��b�G �hG9Z�&��p2��J�{{�d&�{d��=�g7�sf�i�}%�QWA	4��r��_Hx��٥�1�r;�C�^����xkזx��M->ABi���6��x��K�������{��w_<�����{y��5VE0�C����6��o
�������������F��S�p��,:�e�5C�gr��g	�}�2�&�5j�O�]:E�ս[�z��  �f���{-����r6)�?n�P�u�(�\��!8��ȿE*�X%m&��h+0u��h��Q���\��\�kP�x.�j^�/��7�K��z%:O��Jsz�S����۞l�wC��vT��3�����u�C��/H�f��K6קg�0���q:iRO�"����Ee��γ�Yy}js��0�K��۽���a��<�9�jc�l��y���
�ia7C��ôm�3e��t6W:�Yoz������:��`y��0�`d0Q�"�q1��L�䜚cu�^I�g+(Z8��ȱ����^�Q���v�8�c�C��:|B�Q��w�������5�ec[ݽu��>U��zȇ�c'�w%q��^i}EI�|�'i9��4����5R�Z�T'%�onX�;�SOT�Msp���;�n5� �f��K���J�����qUјxc�Z�����G�œ�J��[��is>ӗ[�<�+�wF뭝��nP��M�e����ғ�X�dڟ���7�k������C�q}���7Mr����3VY�aW:�;X�'a��:�ҡj�Ja�Ʋ׾]>��I��C�mCX.+��b��&g�֫�������x>���!�bx�t�|dF�0�N
c KC���+�^�b5��9�3�j̭�]��VVy2�߃�����	��^��aΡ4	�.��lh���؅^�Z�隃���� ����t8��-=sͼ"]�CF��i���\��m���>l�챞u�2��`��z4U�s�a����kmjO��m����I<bO��՟�S���d!�Ji����m��^<�z+Z��A�Y�� U�E�|ئ[�-�<�zw�`���s��e
�sr(>Wtn�
K�i���U���j����vOAd	cU�л�d��9�="§=�749wԳ�֠�`���N2�%;H]:ū�0��e�~��XU
V�,&��9�(���!�Z�b2���V�ϒ!7�(R�u/	;W�e���&,��tD�;��r}�H����EE�r�ٻ���XV�(�p-o�QW#{�w�<ƈ������]7y��¢L�iT��T���i��&�z7._/�3R���X֊0�۰���9�Ϣ�Ž`�Y5�����w�}�uwv����>��&E���x���}�'��;�.���*I���P��}]����,���L??��xg�~����?���k�HW���u���3!6�v�C$��r�կ �\�$����t�zw�xa;�A�C���OH ��9wHo]<�����C��fk���Z�)��M�.���>��yv'��������x��e݊ivg#�oQ���ۇ�ֆ�u�s�ɺ�a��}xe��Q��*�]��a�a>O��r_)�قKB����ެ�`�_" &I�y։7B̀bN8�*K�]<�n�k	Ot[M5Ў|ia=����s�ه��p|e!��~h��1��ͻ��Bպ��:�~��eA/m7V���&f��]�evc�K���Aܡ�8�fp����N˲��,9�aJ���p�äR�ђ����v�,�]���L75��e���3�D���D&�m�X�쓧-�.�v��+rX��X��vrv(U�,	x.��2����f�z>��1eyiiW��$hy��><�>�V���~�3�lw)�`��/�y� �rT@���>:"�WD������U�L�Ųjz7Y^�̇5z���JI����W�V���p9��]��3��z�[��80�Tw��t,������}<��(PP�=3�{kW;}�⴪>����5MoZ��un���;;g'�Tg�|KW �>���
=����w�҇��es��
�i`���L�u!���C��y����SQx��3cZ��-��G=r�"k�7N���w��]LU[��Ӱ�P
)�XE�%����{��j�*���r����� ʂ̡G.ְ�g
�.���V*�Q�ٶ똦�V�)���8f�cA�3��?�^�C͜��M�yb�5f�W&���p��rּ/�
�Gh]�Ӻ�1��i흐/l�A{�L����C-���e��Ĥ*�s1���hN��1)Ղ��L�)�o���xOm��$8��� ����ɥDD<��a4Ny�Z2��]vM�H�0%'E�[�ƒ4�W�b�� �s	���xM�3Ο��;��>eف%����5�l����s�r���p0��yL�w/��ѯůi�mP+ÿNqj�������ni�!7G@Llԉ"�S���*������T*�7&��97ը�����Mq�hD��al!��������٢�S7���9B�F_&'7�>[��i�v�����(WP\�sizp�-�F��a��k�xN�U�E�=^�������{؆�!Z� 枘�'T�=��zl���>���Yþ5�km(�}�-J�3��U;C�F<Xܹ��p5�D���:����n�]�m���K��zT����w!h�wZ�C&�����h���/�i���v&����B����w\Y'u��\�)�y��PK�<��50͝�l��0g��<Dqwf�M3�T��,Uo㯘����3f��I��Q���z-��k�f4��K�j�`=�fWY����=��%�{�����!�5������!� v�y�L[�X�c5�LY�(���8�gh��wu���k��Si�N�mC$�x�s;8��D�,D��l��83Zo���J���g("l�si?VI�gl�"$V����x5("��<�pm��û�	܌�آ��Z�;��y���OD����Q��Gr��	�7\s����#^(�Hͥ"�O�YŃv����ٛ&�w+���;dm����>م>�B��	Y��w꺉s���]�|ƨP�\c5�e\+6gz��B�.� V�h�W�q��˽V���X�r�oD��}ӛ<��}���s�r�_/��k�F�<��Q���3�M�᷿����~u�N�m�������D���Y߆Q<������Ѽ��o|�sO�� �@�O=������Ϗ-����s�������l�3d�c]V/jz&*�y��Rg%�ᒮ��J�鞝ޖ򝈷�p�KL�����up�t B�[]"��u`��Eu:p�y�V��ܼ/�S�\d��o|
�OL���W�w��0�ە51u���+�j2ُ�Z���ò؎[�k�T��c3K�����dM�g��㋵����V�Ӱ�n���0e��鍕����\��Ju��sM�e=�t���.��}�B���ww�$�$�QY��sUuH̓'��J�`��%��f	�����S����]F�L�~;�B��1Q��D��	'����J����[˺r�;Cs��o�w/�/v��nL��b;�m�5���}�e�_�;69�Kr�yY2b�����gtI��!��t6�i��x��i��ķ��7�]����x��v�-�n��rG�^�����xltS�v����UyDh�w�-W�wަ��j�������
[k����8@B�y�����XR��}��w�~�)垕z���1N���CO�R{U�x"���<X�����ݲk��5��g0��58�G+D�J�l�B��s�,]l���"�Q���'{�G-�&�r�+��Uς�Kȍ5��kl����}��8biQ���E�P2U! �ƑyJm[��f巵K"�m�Nd�w�cs�u��ʨ�=�����.:��jM��꺢��ҘD�;�GX�ۤv\���L�qb:�Dp������+��_���=�Pi��|�g���ђ˂������Ĺ�*���Ȼ�HH��
��&�4iI.�n~���{~�P�,�6}zk��l����{2�1��!p��.^`+#%��._�\�>����zy�*��ϒ��o�5әq�C���x�Ϋl�����1��=������8�	Ej���:�[ϲ�Kkl�Q�Y8�����Y}��p:�e*�S�7���.�����ۤ������Z���4l�q����o#��C	1�����>�[���i\�w(2�Y�7��m4<V�m�.��=UL��q�oU@HЊ=��WyB�����o��������o������������}=��Ż]����XK�����]�����ή�]����Y����3Z{�k��AL�,��Jͬ�i#ې���0 l_bSA���H��N�����({��F�/-�!�5�t�¬B�v�^᷇A�Y����i���=��~G8ص85��u<��s`�ma�Eǽ���]7�i��p�F�o4����u��N��{0SMԺS3�kk\�1<]��P��kǏGG.oS K�Т��:�fU�Z��s����z��$���˷CX�N�ZuDý�#�}�H�5�Ա_�r�x,^�ޗ�����IO7��\֛�-N9�ٻ��B��;���u^����vޑy�i��\9⁅g��,�E)��P{tؤ�� !�,t#-�/jt��v�������H@I�i#�F��	�3-�N��]s�%"�<[��x�����_$�@�[J�H,:/,��`e�Up��QÊō�-���m�$J��u���+X�k�E�h���@��l�;��ݤ�۵�qK]}�ʵ�ڤ���ϴ�j��<nb��3����TWa�o��5:l�t���W /T�b��s9�ju�����9�7Zg��n�T�-�Tׄ^��1u�|�I�+�@�)�I��#�p��ɺ[G%�ź�����rc����'y���n�#�U���5��H_�K���u0��w~𛍤�F�n<�u�bM�e�Td:�6�gnm�U��H4��kj��do���Ϭf1�bc]և8r��Ld`���*�e��\g��x����-Ro_`Ls�\�t�!�s�Ľ]�O��5�M;�;[�^��*~�{;9�y���Auۼ{f�VhK[U�PJ����3?��7�,)3�;��E(���$����c7)QH�Gsj�v���V�
Ĺ�Q�����C#���Ⴤ|K,��aθ1�(b�˜d�\�9��!���Ê�{iE��]��-:ܜ;Vm4�Vi���W+����$JP1yݙ���J]铚�\3۽�s�eY��;QK�e��Hl�ÝtN҃qG��ݹ&�n��R���\�HO_�?����Ѿ�O6�W����΄��S��w^܎�e��D5++ �3�f��"´��W�hħò4����k��Ât��u�ҧ�S�kl�:bk����Z�tVal��sq<θ�mb�h(\�����C7<��]���S@��U�oK��n�E�Fj�2�R��U)��.n'�4ޘ��̸Z�{��QL�f�bR��-r�D��F�J[�}�G&����>,��̭���! �olK�q>��d��s�yn�-�ƺ`�jC\X8�1�ݎ��L@�f,�t�[{.��g0���ۋ�<��sӪO�{3qh�\F��e�#��� ���B$�����s���+�+#�8J��ocn3���йj��a��xRw��B70l�vObwtծ���,՛�Y�PV���PH�Кo��b�sG:������&�6���K{ue�M�z�6�?H����>�r�6�F�Qmnl[nnkF���W5�kx�oMk���ͷ+�wk\��d�lj���ccm͊���ܱ�ѭwt���5�v���.5��s-F�k��7Mn\�9j+���7&Qn\�E�9Ͳ�k	W(�(�F�k�˚�-s]5sX�F,����WwFu�V卋`�Ӝm���w��9j���\��P�|~_'�5�<���o����=}��@{�\�%��	�f�+���E�r���h�d^�3um��ę�,�ro��&��za�޼�L��ky^{Oa�����!����$^�=ȇ
 >�.�)N�w�f]�[�H�ɺ<#7�pv�&�0�����<m�����a���y622��J�����׽��뜪{U���nga�lK,��)����#{�=��*�e���n��fZ i$O�HO�s�tS�x͜[�qs�D9%���/h؎�=�/s��݋�DMq(�rc����ٶ�߭R�S~��o�,��	C�ɡ3s�6��PR3e�ת��؊�@�^�?w�'봟����L�UA\�-��vj��[V;Vܝv���;�4g�xNݭ�J��Q�ɹ��l���FP��I���8�4�s/�W���7���2��BZ�uq�rN��7���'�s��;��Vy�{��<���&������锕�����=>'���}-t���]��ٓ>̻����AyGX�G���.����X|�v��϶�d��w\�ɋj�@.�7oxvc�xw9t�أ������7�L4��	h�[yW���v'�d��f)�u;�$%��[��t�tMg��wDq��n����&�6_��<m<
�%_�rqh�/7+5�.3����[ܚgi܋��	��C&0S�1�;b7��0ܚSL�Z�(�^��t��q5�n;[)�S��vc�*\Gkl�-��"6J�D�7%۞�K��:\�	8�������;�mt���!���{@��L��el=�C��
����tƐ�����	s`J�������6}r������%��O��NN᦬m��<���^r�W���S�8��sƃw7Y�M�¦�[٘n��k�> � �w��f�>ϯ��/�E;g�t�裾	ɣ:mln�Ɠ���ᨉ�p0bC:��V���u��ĉ��;�]*b���x��_v5�y�)�s�[,�(�f���~��}���"f�En6kԇ�1G/���{�^]`\K�VR>觋��=���	G��M���G�����1v�a?K|}
��a��{����'������O�C1�8
�|厚a%�a�Vo����6�<kv�Co����������Wb���,N>�eq� �eʜ�����'85�K���@��J�4B��N�Vt�:8��=83��8���[Ï��4Q֟�R���m�|�#X"�\tDD4��������1�7�[\�R�&����/W�4�j�P�c���a��r&�0��}��$ wj.��@�P��JU\j���lVcر|%�5�e��϶��6���\�rU�Dz��gH螉=bʣ�i>u�g^������e��>��k����[$7}�_���e%���(w�吷�N8t�U�{�{��M��,-�\9f7�M�Ij�U�����e�5ټ�	ŻM.W�����vn��-�9ˮjb��N7ݐ��m���=Li�*�a�kL�]һ�a��A��ƅ^���v���;8�4�8��꒜A�4��oZiA� m0֚�P*��tZ��מ:- ��E����ңu:��t�I��_�b������)�:ʳS��̃_RKFX-�Gk9���Y?���즮���ƍ9�@Ƴ�����ѹ�H��-���`�f�ЬT���I1��m-�-l�DV�Ė	/Y6�o�;��W�Ms�uues����Kt������Z����X��gS���_=ɼ7�f�̗��t0C��E��}�:ؾ/�e��*��[��j���f��U<V�]�8��:{E����G3���7�é_����2�L�mc�ډ�C�7��$�"|pr�K�o����g@�{E�y�%��=���El�s �����v���Γ��#<{�-�^�3��`�lN�]L�ہ��mպi)(������ߗ�Y���Y@�T���yJ|,'�T�rU74�ŕOݏٰ�`��M���Bfɡ�+�Z�`���$���F7�]C�L�}�7:�'M;ϩ3��uw��5��}΂�P���"�ŗ-��'9���)���]�:i�M3���PEȄ�V��ժ����I�F��,7Q�C;�+�q�{� n[��Ȑ�<�}![�j� ���R�f���Y����.#�h�$��L�.2+d5S���_�{��݈���u�j����D$ɱm�ȫ�����.�-��yk�{S���m��;u��ʍ�l@1i��#�t�]��[�Ĉ	���s͜�%��<鬂�}�wB/�q�W�:x�n��6�v���I�{�jd/��3��B.9N�}��.�O���1�J�J㬏�� ��n�3�	ɮ�危���,A��K��9�S��UB��T����J��oK�&��t����}�v-��XvC��Q��4d�����)�e,r'���Q�j���u$���8�`������c;Vq��B�ﴮ�]��.���=���"��R�G썞���7�s?�e��=�������ͬ�z���G{Q�=���n�Fo>��6h�c ���皳.����i�7gmGU�^��ȼl�[ܨd��=ql�eE[��X5�Wu����jƜ	�6�.t��GGt<U��įy�3,��$O�Hr�â�gT���jm�k6�nM�	��^��"�;��o!�<����9����;��q�a�Ğ��s����ed��x� �UA�~�}�Q\}5u

`��qO�7v*f��i�����^�k=���
U|t13�+v���ӯ��7�#��Ϥ/�	/�dW��1B�*^�OU�n.��M����k3zJۜw%�x�f�� B�!ج�a[�o7۱R��/nԲ�(#�F���=ٮ[��9��N�����9��!�:����3��wU��{oK����PF����č�v�؞��M�ɵ����d��,R�B9'n榜ղ�0�X�0s���l�*��Z�s�vgp�p��JB�������wI�R�T��(�akw&nЋz|������!:Pɇ]"�|g�e%e�,Q�	�)�^�5��çD����ծ��|�G�����x!a��3��|�c�Ns#�0+�'����T�W�˿Nf�\0�������:�Ք�V��k9t#nzby�07S�u�+��q~�e��k�����p�?O��wi>�Ih�,��P�J�gx����ݻ�G�� ]>4��c8o@a� 8[ͺ�V˾'�����ֵ�*x���~4�Kh�j�m�S����m>�0;u��XTY��n�8\qR#d��R��l�a��N?��@�����(K�gh�(-����T�:/������'�کЫ�S-��9ߏZQ�Z�=�Dݢ����Ǧha`�+Yz ��)����$R���+1yR�M�ר����z�:�>��s6�dvbyci*Mi,��.��Z&>��u1��}8�.�\�6�k�]�qݍ��-ɗ�L�,�H����5�ȾO�|OP/�kĎ�����cD��*M�F.{�J�3󳑪Y՛��f��Y�ǅ��캧V�QƷ�;9����`�;�FCЅt?$�:��9U��u#n5�>�_sf����}w��Y�"^eBm�s#%�s�AW���
�%F�=�i�&����wQ˷�5:A�r q�J8�m)�e,������=��D�����3��#�Jz�aT2`����B��V��w���rx�W6�ʙ�|̼�iGu�h6���А��m���C��@�*�������!3oy��Ʀ�؋4�Ԋ�q �t*a�T/G�Fu�5����c��v���i���ڶp��]t�M�+͌�P|঴r��\K6�-;�FoC'N�ue��cF�	�Ǭ�f<�+��$+��G�����~����3���E+�n�&�V8�lu�fe�ַ�J�{yݵ���**��?�B褊���zj��uG����MRޮ�q���Ė�Lt�bo'b��$��bݺP@��
u�^��u�������v��l滂�G*.Nҕ��o[̸�㔑��VJ����W���
V�/�5�<J�w7G�[��u��R5����{;��h	�=B:�U񞵃e����+�B�x��mu�g�j[n�ȋ�O'/�V��î*j&t�r�\ԞJNgB��������U������i�7��^۰"<�E�@����5��@�\��]�8�S#�m5�����;�P����e���]>~�h�[7ǽ�R.˪��6�s�T7���ٱ�֕��)��x�A���́HgU�"�%X\��ű+5�S=Oo_c���<�}D��@�n�\K�:(��c���x/���n%��A�S?g�ܷ='nZ��K��eOJϥ;�?#�����i��0�l��i]�-��:��vWT/;g@в���	+��"�}Iه����%��m��PS>x@���Q�&n	|��\���|mI�G�l�4��P�y��������,�,��r��u�:����daͷ/QVª[�	�Մ1^�ő�~��.��/�˽=ڨ]M�(�c��m����J���;����3��9ی]s��5;|�t�j��q���t���o��{6�;v���M����[Rr��<ؠ��Gh��}+�@��-�]#���0�d)�OyYMv�dn��]Ӵ �;��/SL�@�("�+xMY���43Av�ީds�/	P)"�e�����uy�!cO��=�GU�-	��511�l��<e����΂M�4K����T�Ff�`E���R��T\�����A�_)Ue4z��Z�q������;<�zh'�gǭ���ÚwE�		s�=��5=|���ԩ+����ttH1S/WZ"z�oK�*8�l��a��oW�d��FAκ�7�(���h1��e�m��½sU0'JW;�Lq��7���`\.qڳ��W(�DV��p{�(�����������R�]{�ul`w�Cz�b�#�o���Cok�4q��g��n�Yѓ�=�ɠč�Z}ީ:M4s\'|aQcS�RU�H����#��8�	�F[q��N�h��W]X�>I��u�3�Y�A���A���з!��R.�$�"P{$2��[������Y7�}�ZA乢��puՖ+�oWE����c:����lfL�
A�$j�8�WX�ϧP�b�^6Ej�LŶ��*ټ������M�)��\���N�ʵ����J�/;ů��љ��~��H��V���,U����u�+���Q��R`\4>ɜ ���d�f�f��"0
㯊f#��K�~�r��v�H4y4�R��?��C��~��Wsͮ���,>b�ɡ`�'w����K2��ƛ�W���:A~����)�+q�������=1x<�'X�W���sSNd
�p���ř��1������N���U��(�|z|܂oH]+��DBJ�>]��)˥32��E��������ca/d�d�)�@|gL��x�%�;���s�/�h��M6��A�]9�`��b���>����$��)�bw�T���i��^�9��Y�-��A{���]{PM��/o��������{=��g�������}6v�6��9'�3�B<B�"����ƴp+z*���H�3՚��@3��A��/�������˨��2� �Y�����d��>��ӵ��ya� �D��{�ߣ<!�醟g���۞CD߫FX�4��].�e�5��'��j���tM)�I�߳�ƅ��p��o�)+�Q���|�y����'��M�Z��M�7�X��"wE1cz佝�Q��F��	��3B�Ż��eJuc�j�h�����������ǳ�&\���m�����%�dX��>�k�p�.�.�(�H��Sn,�� e��u���(���ɠ]�x>;*n`�Ҷ�/�"����)�T�u�W�h�Jn�4[��uD�l�T��r��ƥ
��AU}�R��4�4�+O��㘷�Mz�9酓ar��6�X����\�kTS��ђ�R�4����B*�ꊓ���:��)���}���ը.�&�9�z5�I#X��Y�p����Ų�\��"�x��]Oh~x���Q�[O�
I���Uo7���^ѐ7Ǻ*uNq�W_Y�SQCE7ٖQ���h@b�l@Uۻe��u���-+�«����UA�@�Y�eO[:��������<$�]�����BS���J�:/#d����!�ߘ^"gv�=)ܸ�N���1�z��#��o��M�v�j�f�aw���HD�/q;lC�x���iPҞ�f��A��M����}���hS���R�~S��&�����;|:���M`�4sKlO?=x���(5���J�������Ww-tβٹ�@��y�5`9�E�,����coào2���ӖZ��p��'3)v�ہ�5q�jv��k��N�/ky�Q=#���&����{��nxǋM���a߅��Oe�<�+&ol<��h���W�g*���C�̹}zU5j�%��b��vo��c7�A�x{Ys޸�<u�ߴ�7�E�<��du���+ٵs��U���\ t���|���0� QS}���xg_!���C��Xc��°o��ڄ�^��sze�����Qk[�Yὢ]ʕ��x�O�c��N��-��CW�eW�:��@ț4jm��˩D~�[�/gR4��7)�&@�c�Üb}������<�u��Nx<��Ou^d��������K�ڸ�qP�Gz��L��9��`��K͌���N}}V˟eR�V4�3�
�u(�K�'��5%�<i��v��zs*E�����hI�ϯ��ܧ�:I��DNt��;6�j��?@%y�K���tpQC	��+�4�l�*7�z���vK�((gs㶺q�-�qc�~�:p�$w��C��)�^ν�U�'�i>��EN����l��b���.)��SL�ӵ�����	w��lT��aI���S��6��ф۝���t�ހ��|���+鞑��}1�N����þ~����F����Z1����X�W.��Ƭkss�+�r��.n.�]݌[r�#nQ�v6�r�(�`Źr�k��;�nTn\�ӻ�3�ܮh1ms��l�]�l\��K���۔M��-;+�h��sk���V���(�K�����;��Q�ŋF0h�]ݮs;��s���@��wmrń�+�0X$,����"53�5b*#�oK��wk�� S!��&9¤*5�Į\�ˡ��ӻ���>����/]���|b�ѯ���6�͏��H^m	v�ޞ_	t���� anǃ	�	�JX�_��i��W 9nQƉ��e+�.��r��H���NFd)�Q,�gQ� ���7���yw���~e�
&B��(��:�/���~#$����i`۳xy�sC^�R�����r�F&�s��6�A���oS���a���皓�OU�1Rz����t�<��QR��9I�}�T�"C����Q���0b����b5�'׽E���w{N\��F��oކ�[��Ӡ�_�Ы��M(k8�L>ٟF2ɽ/����5�Go ��>��T����<�Zu/?~*���A�]��v	%�³Q��f��8�nw+sg��M�����׏Z� Ȩ�cD�X�w
�~IPהEM�HU�-�3��p �?f�)��;���	����.w%�5�nx�	3Q�����^��/�gJ�^��\P�+��2�����6���P�'��s0x�^�Vn���PS��=ܕ9��Ln�4r� �߰q�T^_�׿�zh٣�g��=x6�S�l��{$k��f�S({��e�^���n:��rV)3��=��+CX�tW֤Fl�b��n�
�p��8�f��z���#��'��-�����ؤ�EGٻ�r��0R�*���W�fV��.����^IQ�r��{�U��ʡ
�;�.�n�Y��J4R�8'j]�'���{"2������}�ߪ��NEH�EW�G�φ�E�nC�t����za�v�n����h&_y�_�Tk�QS�`k�]X`u�H6pW��ȭv�sd��7i����r&�s���5�= �]G����H!LB�!�#Gz���^޷T"�,qq�+KW$�Q�\�'�	@�-�%�uۼs=�^���W~1���������V���񎥐}E#ww�c�.���G=�j��/t�n���2CF(���Χ�'|`�Q䦖�W]�-f�<��*����%��CP�`����{��8���ziP0WPe�z����[KI���9��F���6GPn��o�����k-�|vcE�m��m�Q&܇�f��꣏��������lt3�ρ8gU���M�3���;�C�C�Qe�\?@�wI��6��o|OAF�Uih[�<�4����z-)���p���rT����a�P:w�� ����}9`yd��$�;f2Q׶�+釥)��hU��a��n����t�W ��9��Py��Tw%�[����n����������tQ����t�f�l��f�O��d5��|�Vw5]�t�
"k����M�ޘ`�[M�<2/t6"(��"����P����[>Đ5e%Rp���d�Um�(�Nk����|��/A(z��oY�1k�����L�+ro �Ql�;��ʩz��I꧇5���W �w��ђ�K'Q�Qw��5���<o7�ٓB���tK��Z.@�A�'�םlU��rK�L���7�>.�V^�
J|c�S�)ܷS�̉!M�A`��ek�*��艠�tr����lǳ�̒K�L���em|h<	ۘ����i��w�_W4As�1�t�)Ue4Q��ڥq�Ef��y����"�����>�]���$� O����f�OU�UVW<��~?{���>�W��f��.Z���4�8���d�H�vƖ3VrFe�b�����:骷Iss�*�񡺳WVڲw�-��$*�C��4Z��_��L^��i���.����"'V����R2&��Sp�*t����촱�%���"~����4�m�t��)*��I�c0M�{����Z˦*����͒�9�V�++�f��A'�/�}�*��B�U���`���5�`WLgj{�]焞?�RSb~�%{L��}��L�'��q�r����St�a�����*f�o#�|��8�j��yc�ڗaHד��.�����6h`�����"q��z6ɭ=קm�Ʊ9@xW�������1��Gd��@���fG�3&��+;�M��({U�ѨZ��ThF^#{�љe�i$H) �脩ʋa|�oٺ���;ȻY^?��$~�_�	��d��ؼ����pc��#�݄��h9p8�>(�r~��#��f�ǖ8w#���?,dWC��:���?LOf��U��u��[mW*�_��:A�k⮹��Ս��3�TB��&#��,<�!b�P�I۹4正����W~���'n��f�Y(�󾺾v.�ɂ?`��ߑ���:��������ˁnW��b��9*�Pm�Z�2��Χ<��O89�ge�:���B��)��aP��=��{�)+�"b��ƶ���la��J���ޡi_IQ���뼻����~���*��|�r	к��N�����˱�M3�}n3q��`����!ʚ�D{o�24�J��T=�{7���z:	|拉kܪ7F�c���kd5���\!R䭍�γ'ƙK��	Y�
��0llM�4�s��<��7�g��Y6ǃ
p������;}R��~=~��jb�����ؑD�\_�#/:�a|1�&��ךS����x�¢�vw'v����²�Q�K�c�Wt��L݌�!�u��zC	i��Z��I�X�<�z��u_��%���T��s��2��]Z��³jX��s<t[�9�1��7�J�A\'����1̃�/y۸�*�zm��f�!�\rd9��#}���2����=E�O��Y�S�p�͚x�A�p�"���Jz�k4y�gVn7��N�ｙo��O��BC�!�K"\��#��?�zO���>T.��yw+鳎S�L��]�d��tw��Y�;G{3�VK/�-^n�$x�8��l��6v苺��F�{S�岔��lYK#�w�b�Ιs�.��6E�nn���F�Rw`př�*D�N�W�Ր{�`�#b��!�d+��$ϨZx$T�^���m�w��ܷ_oY^����$y�YJv)����DE� A������!���D�U{+�\�q�J�bm)�� ��c�����!��G���6bU�#x��9 �\uz����.�2�8�z�u�O�i�E �Wb�H�[>�@��(�g�ߺ�ܡp�Dh�����#2g��F�u"��p�R!�U����!�k���'_2E4lt�ݞޛ>���*OUW�j �Z\X��	�t�=sD��0ֻ��}N�n�U^<�%c�q�5�����e�4Z[��	w~�Uck�^���l�+GM����ErJ��6%���<;����9�8�F!�]��úv�P�!��>���c��O[yk袑���v8�������Rkj��{��d�6Wn��V:����2��Ǌ����kA�c�Wb<~�VKm���y.A2Mw/kťո�P@~"ga�S����/��/u���c�֡ɡe��Ԇ�=�&-�nR{ʆɮT�Y��k�}�C��Vn5�r��(��Q6}?�Eca'�2!�@#~���u��5dq�^0n�ǒ��b6�u�;��%������/܀Ad��)�z8f�"���#�NM�R.W,�'E�$Ϊ΃��ٽ���UBt���7�Xw�H�0!t?b4#Ykl�L/4V^dٚ��rh�o+	�/���_{'��y�G5�
�'�K̶�m��NGU�V�"{5�7�z8O���%�{Ez���Q��ns�0��]����a?y��RjҼ�2�}'��D�����(26�3����m"��� �p؂)G���M]^щ k�P2U!DUג���Y��,��
�������6�*	c�OP6z�LR�V����^þ���Ŵ�P���:Ǧ�Q.dagA\s��qm����x��}���bf��)�fW��l��:����4�4��@Pa������6�;C_dV5��SM����m&�("�{��S����&|ln���<
�P6*a^�U�r^�ʯ6���s�m3s��{��c��J��ہ����lb�;�E(5֡p�]�@D��/��]9M�iH�C�oB� �[�ML2�&i��{���յ���#l��E"Α%&8�y��r�Ofl[���A���Yxd��'�;=|��Љ�I-h�w�enm��lA᪯��Sk�Hm�dy��#��ʲ�@�)V�\u����f�A�^�Q�����:I>ܒd��Z=��?���w���U �?>���剰ƛ�����;Τ(`��l�����ޠ#W�=4v��)��194't��wv�q��]��(�*bwt+����q���
�H��ͽ�`�kb��Y���
�/'��/.Ք8�R�+���M���0~�'t�24:��RwA�чlV`=���*����n|�oF��:�0ɶ�[�g�A�&k���=������µQ�U�f
�Ɖ�$;'�>K�d���W�5;��\]V�&:,Ǟ���7ve��Hp��o��i��FkKS�h��#�8`�ME�G��w���=�c�hЯc��/k5���
�4;C�`��+�}ѝ���u�Iz�M�c��聛� 37�uD�w;]VRe�8�ʌg��%������i�&vɥ�}e�(��Iî�Λq�9�q��^���A���t���g��3B����1�恺*5�"��
,�s�I>����XzK4�+��$�o@�w�>h�=ɯ%gE<l5�%��sH4C��]m��ugwzꞎK����2]��=|��L�YP9��{>nʥ�����#��7�rq�� -«&#8��
FM�5�=�ۺ�sӮ�r�/�{.�Xu�+XC��=�!!�D�.��h�4Q�@BJ�.����/{r0G!{�|*���8��$3!Үf��)+�xK��k6�KT��8'y���yy������#Y��[Bw��d(6��a��Tz�O]�G�;�Ԑ΢W4y��},[c��?�A�pX����y��d��K� Υ͖�W�dc\+�k�	����;t?].��v�wV���P��=R`�^�y���KF��](�~;�mq�c7��p��"�J�ne�p�e��n_��|�N�Β�U��q֍�t[������Υ��|h���A�<uX)�iN��;��a���}ڡ9��0�vZ��Ta�F�%�4�$B�XO�L"Qʼ)ӟ=ѧ���[�;�j$"���;f����W�yá_�2L�m�ٻ{Ճ-0��I�5dt��F�%�
$���nW/rG�����m.lJ�n�����a��[r��k��݆�!Yх[�;��rc�1`�7r4���53�f�	0�f}�&����<�jf�4<=ս�
�wVR�vI��������s���7�Xj�����_�e�WSvkq��	DO����
26)�FC:�
�	�s�W11�4�7e��v��]Z�j�:jH����jKଥ kEA����N��k���xTv�T�z�2W$&��4���l��4l�>��޶qmw��n�bB�ǀ{�T��>K���.��*�uH|ɭ�q�~C�զ�#�{�������5�������j�p�u�)u��zCC�L���o]Z�=Pzd��V�j�� H)�0�gl�[��CvM9����lٳf͜����w����÷�c�W�5w�ua��flj��E\7A[ܫx�B\��d��የ�Ĳ�Q��|��}����P(���G�G�Nz���v����`�ѫ�@K����v�좳���7U�ZC�+� M�JG>r�XΥ8�9R'J
ڵ������5�.`��Û���z}��+%�O8f7�'y��FV��`�^ܲ��x�^�T(u!:wa�����V��A���Vحb	,���3�=��	Ր�s��F�Þ
���=ﻂ�i�ص�}����{��BzȱN���b�!O��{�����r�O+���� O�~'"��K��5��xC&��]Nz��(���y��(.�eڷ�K�nݻ��,Ԧ�Jv����8��)�3����r�1��-�}���g��|��m�4c�p�J��X�Iqk�����U����ᔉ��̔)B]��e���>�'b'��2�{��T�d>ţ~�c�?c��H�қ|����ǩ��F�=�774tj���<!@vvux��r�>�Y2��N�B�-^"��g�¨>9-�if�zr��˅��v���n3qvt�lD�����]�O�6w\#1f�������cB]�dVKR7M$F-�h=�u��W�U9�!O�$'D�,�n�ί�⽝=ꩠ(���;���DO��{;X��}D�%�1��"Wًi4�b����6������]�"�狮��1�Zb��C$p���7���6��.u�u	�r,۽��8N~�y���˪���uG�`c��� �TZm���n�޽�AU�g>մ���Z@�C	}C7@5��x�^^n�N��a)���-�a۬�z_Ϸ��?&�7�t��Ӥp������R`+%���;�L�6ۛ+�4{Y��|w9(�T,�a�����h���Ӯ{k�s'@���
�5��S�E�ti��K����ټ˫e��S��`�iݛժ��ԋ��4LFIá�U�aņw{������٦a說�	�{BdC�������i
�)�ٸ�7g���+_de�Yx��Z0�r��r��2u�>��7����b=�Ŵ\ܛ9��ś��0�A*����w@���G��ɼS��=�	���e-��ѧ<���S
`�v���e���پi�z���j�ۦF���!��/>�������8cWgn����Nps�q�y|Et;�Ա: �޶8��
�*�\I��t�	�g�:ƨOv���hjI�޻�R4R���ܘz�f�o��zOv��BS�{�)�^�^ߺtWt�x־�f�s���HP��:�+7Gwq�q�ތ�<fw=����{��E��"VI���1��Ea����Ϥ���)ޔ/e�'^㜦�i��k(R��ξ�(Ի�sN1��XƦ�t;4�\0�L�;�K�:u}ӟ\{"kX�RfX�W�v���s�s���q�Th��]ۋ�W+���Id�\�b.j�ݹEc\�n��@&�m�I��.��,Bd��jdfR$W;�2�L���(�S4��\�I9�1!����C���l`��(�JX�P���sIl��Td2c";�l�S,�]D\��3D��Qr�	&���ѺR,�j
����(5�ۛ��;�4Q� �D�b��ґ4%�X�!�ƙ�1�ݫ���b!!aE� 5ع�QBVFD�6����D��Y����'up$�	��H$��|a��i쾋�^�z%,�_�U���j��vk��L�����-^l��˚F?�|�{�&\�ܷ��5���=r;��t��AqH��gW���q��xUP}���Z\X�
�E�o+|���N4e��6�S���RW��k�������I�L㥲åϗt�+/O����dF���R+�ErJ(T�XO�k��NA!������jmĕ��Dz�0z��ǿ���Ut���Ɗ)�Wu�X!�|�Q��a�+����aق�p�t0=xȍ�Uh�0n�P��O[�6XaJ��S�7�3	� Ԍ�a��z�o8(�ve��.���^��w���W=��ܓ����I�hl��7w�|��0]>~�]�fu3�kt2�2�C�k�4r{�/��/���#�o�߫�����}������vP�oqs�D�yWI�C>���67�������4ϸ��tQ���mh�CLT�V7?mI�f��A�~(>Փy�2�}'A(�=��_��1�x���%q~�D,��S���7���z]~y��ڔ+��
Q%�<�`���co4sxV�\e����{{�ɷˍ,�z��k��3�6�چE�4ԧ�\P;�:)���@�Yt.w�:�ʆ�$��4j�{+5�u���F�h�Â�U�4P���s8��MV��sQ��s!@"�]��59�ò�Y@㘋�i��C�*j37�d�W'U9ΖX.�=T�3g�&(TR�16S�EVdeGWޜ>��dRk�i=T�氳�qb ��Ӄ�}�X�q]���8��,���&�SL�tK�L��k|���ڃ+oz:�Ĩ� 
� ���I+�J�M䋓����|j�C�8J��cR�[��2�(�7�Eؼ�}AW8u���=�JjKZ9y.*�V����m���F�6��3��-��:dK�Ѥt��ʡe7z}f�j��)�L�n?u�ul����r�v����=0AY!�.��g�jz�)�I(y}�` �Y�w��۽.ޛ���x�:�!�}��ߗ��X�߬�3��֊�<!a�o\O?s��"��ʅ��+vU��Qn{��i���y��_��o8�,:�������l�s�%��6������d��ݑ�J��Wz�����*;B�5�6䧶^�{Ӊ�m�}�s9�ۮ��b�x���P�$�8��6���w;���6j���޺����N�fE"�F�i\�/M�Q���WU�/W=��Vd����M*t�Wj�W������)����U���[+�泽7?y�5���{esY�haHד�ާ�ލ�^�o�Bަߨ�����<���WTF3��}^�d�٭���v�2D�;&{���Ab�_�Oվ^�{���&{�u�g�.CdY���F����0V��-�Ra�j�g$w�m?��_�mw�7�*��M�: !e�+����z�וSbڍu�;7[�'ս�4D��&��R:)�ڇv �P��qA]��d��������l\��LAvd��yJoH������>��;|$?�/{^�k<�tPD�����3�YG�U�Uz�����!�����7��P����Լ�NT$#��D�.����y(S�<����M^
^#���O����6��"2a�O���s�e$��o4��P�fɿ���4�}��߱Pcȋ�����}�M���d�g+bg�m�=�g�>��@% _��x���){=�oF�����p*hv˃��G�l�bk˕g�3�i3�;��)�x2$׆i���$.=�X����5�F\����Yw�?P}���u#[��tV�r�oz��~WxZ��V�Df:�cpeE�C���YO%f���O���aN���ȼ�CU�l��^�9·w�JrU<�V�����>���x[`0������1[I�U�t����4@~�q��]^�*�J14��������m����/�5�F��w9���|UzDl�z:T�u�҉��L%��z�q�2o�޽"�?I�!�q����ܐ/z�9[>n�qMy��Ɲ�&����܀���:WP��w��h�BP�LcnO�K靔����sq9�8���vwU,u*���:|tQ����vt;�#~xVj;ν��5H2~��'-�j��M{I"�8{^ ��:��N`�;�}O���(��Q�js�_s�5�:�6���WDE�;�h#�@���*�o���QO�\u��;9�j����Wd�?��.����G�%��~1�[��i�A�F!�c�<�QT��Q�ӂ_�+zԮ�!�����:�j��9��N�g�sW�dpP�U�c.}bt��*��ڞ��P��R؜�����Ŗ^������^�J�r��"QƜ^���uϷ��)a�מ5M���
�XF�ɥW�J�c�v��$n�z�ّ�}U�0)9���Q�G��%��AUP�����Sp��xF�wUxZ�'*���9�%VFϵx�*�#2]�޷B�[؀SU���eT�b�Ҽ�s&�pp"�vK�49��{��ETj=�N��_���{���l�㣵��DMttք�v�i���uƆ�����Yo�(�<�۷�n�]������t�j7�dW&��r�ȧ�5�'j��CLݷEP5F�q�j�ل�V�<���-��oO�euGS�/���[R1kn��4i6&�Kt�uA��x�m�����u�Dl�~2t�����Y���X'%]�y{]��9۰d� Ԍ���f�#z���vW�ѷ��4қ���'65�mPg��{��v=�w�ʖoS�WNy�s�q��!7����lK�p�7{����ֹs��f� ���p���﹇�0���M��ߤ��.�{m_��!V�4#{�-����ͫ�[ˍ���ҁY���c�I��\�L��uG�>2�}�'�&���VW.��z���O�0Y�w�������A��_��g "�++tYG�l-��� ����C-�2�J�V��P�#�5�贊�n�7�G�G�tQ�w�z�=Ҟ�-�F�;T;
#�Z���jѿf��Cϴ� F���ލ�G?V_7\q��̭�����@B�D0�F�yU�ó���݈p�}m�ë��z]��X���w��&���F�,���:�l���6�0�i�NE�訞�� U��_dړ@�� �ED����Wa��d�B�a�7�y�"5��s�����[.�?��erF|l���j��|:i�M6��~d�Ki��$m��45w@bDV�{gu�HE��&��LF�b6e���y-�w[8�w~>�<(PY.���q
�!���t"y�Is��g�R�8���t�o
j�ذWL��e�biQ✃���R�`isN��tƛTf�w�7��O1l	7���F�h�k��:�wƜٳd7mZJ�{��{D���D�mitO�L����I��qf�"�C�p-�V5��c��x����j�[k2�s4d�Gr߁{>5K��_h�0��X�#���Uy���FR��Y�5#/���>V��wXq�I�}������@��	_�����d��j-��8��:�'���4�x��<�CO�cd.�淊̎[�!�-{vg�]t��u[Ǖ]�!n���_��l�#xs����r��v[��Đq��V�*U�J�.Քqq�k��٦�!LV��8��:/KonK0&r�pT=�\���^����=��o�Yνa�PZ5�Ĵ���t�see�� Y�#}B1��l�+W�5����0Ц��&�I�#���zu[��C:�Y��F�/�l��{�P��H�s7�{�-ά��U�?�{0HR���S�Y�
#�,�RP^�t���虣�Ϧ�wg�����B&��2FܚE�)�E<l7[n�7�������>���ks��L<m����2#����zja�Qu�f\޷M3Lzo���n&���[������.nz^�_�"��N�mC�0C-�O���Lٙ��h�}�\Qp��KX�U�L�5paO�ʕgO�ܬ���:q���2�vg������OOP?AY �%���]�v4��R�9�0g��/wL��af�`��f�uJ�J�LFr���T)TT�/��f�f��vU��k�k�f�O�����%e	��$_.���������-2n���Nk��hF�|����i�uZDc�W\��8�ڹ�g
+�1�x��ѣ%+�׸��F�<Sd�x5ӭ�TEmN�P)&�j�w�Ԯ�	�����V��L��ܩ|�f�����C�aH!�e�(���lC�a�=:Xh�"1%Xnz�meCΚ:�����Q��u��X�f�p�֟L�/{�ۻ�aZ:���C�/�ݾ�YTJ1 R�ywd\����mo��7����`bۆ�(���^��/�F�%�1!����߶���m���������0"���n5k�m�z�+W��\nr�"�6vӧ���a�Z�ќ6s���5���QV�Δ"�%����yS���n��p�==ęI�n�����p �Bs/��ϻe:��T�z@$��Ko	y0�^i�Ǚo�4���*�ǹ<���A���y�U^o�-{�M�A�ga�T��l��K^k��_�d��P����9��`>٘�Xҳ_��v��.+Z���66���_V#�y={��"�x�puq����o*kik3w/yST2��i��2���z�kl_Z�I���g�1�u,��^[�?�`�F����o�l:ITu�+�U�9�g��BB%ⲗt扇vdONc�������*�DtG�U���������:GJ'z�ϕ˯Oݭ��-�u����ǖk��{�4�����FDzP:��d�y1c�S�>��[�5����~�#��ATP��<b��z碲�A5�y�����ኼ9J4JU)���H�S겘���A[T����?Y�{�ke#��<��49��'�ESl�]:�i�a��j��2ƍ�:�]#�����?u�6�B2s^�I_:�C^@������_9�r�������"��VU�_G�F���m�O��m�s=%�yX����"׶�>SmRëgj�x;ޖ�g4>^v�d�z!�T�@ӧ�v�.����n�5�Ǽ��l���zM��Y׵���ۼx8�N�DomI�������$���������[NB��G8 ՘3\�(����I�����+#7�<Q���}"�T�[������� F�ꎩ��ֶ(�h��c%��n��a|��_.����q�ֆm��:���G)U��'8���;�;����#szh�b�%A���=dfǈހ�o4�+�R�{[2:��K�]A���]�P{��hl�u���F���}�d���(�F�Xˎ�1�|��C
F���hGw0�1��du=yw!��,)�aW��,c>�p����W���}%�@�o3�l��)b�ͱ�z~�h���m�Lb�/��	K�Z7�c2�y���+SG��4*�#De� �@"N�D��o����_��h�����:G��Jր���Lqv�6qV�����?��[�CN�h�U�T�3
e9a�/�ɯ����  +���k[ko������k[kc�~����Y_M�z�V�Y��[2�el�ٕ�+fZ�kfme�ٛl�ٚٛl�l�lʩ�Y���ٕS+fm�6�5S+fmfkfm��l�lʩ��+fV̪�Vf�e�Y[3m�[3[3m�[2�3U2�e�Y�����fV̪�_V쵙�3Vf��V��Vf�f�ʳ-fZ�ՙVf�c-fU��2�f��Y��5fZ�ՖU�k3Vf��l�Y�fZ̵�VY�2�el�Y��*���ՙ�o�޾m�j��m�e���UWe��3UT�US-�ٛj����[UM���V�e�T�V��֩�kS-mS6�S-�S5�S5j����UTͶ�3�UU�m�̶����fV������m�-UM�]UT�m�f�m�m��ڪ���fZ����fm�|fյٶ�f�]�[m�6��Z��m���m�6��m�ٛV̪�����ٛl�l�ٕ�-�*�kfmfm��ޛֶelͶelͶf�f�2�elͶnn����j�[2�eT�ٖٕ�6��K����]}?��u�mX�j�jf��ՙ����d�ygo6ж�ۭ�����
؏�H���(�?��:�EUQ^��;��c�A��.�m��U��[���*Jj��_�m��~Gr�UTW�����x�M 	f������K�	s�a�$Doa P�k[lkm�����6��5��Sj��-�ٴ��ee�T�-��m*����m�Vj���m�m6��f��i��d��lm�U��mZ�����Ru��7����k�v�������j� � �9/����pD]�B��Yn�  Yl��T�SN��K	��{�f�~l���(nv*����;�\�FR� *�UE{��@�A��ڵ����[z��j��o��v�O�IJ/���"ay�����!͠N���6�m�����/��=��mm����{�@�Z�w�R���0����,2  k�~痢��+�*5����9��A����\������m��[o�}k��������|�������[����oᵶ�m���]_���
�+(���>�����b��L���c"��� � ���fO� �k�x(�UT/Z$�T�h�J���U�@��)Pl�lҊ)�T�DJ��JB��
P��*kkDkQBD*+kM�\�c6�mi&�fV�*ڳ��t�F��lƚ��jj�+f*�&��Z���4���eif��gQm�X��e���X*��)���S�KJ&`��e����SJ��d�֥#Q�U��6�d̵��̴VT`1I��@�-��e���kcVTٙ�i�նU��Q(�M��B��ֵ6�4�x  ���we�s�N�Zwv�wl U����Kn�����CvN�iw-v�V�]�ӕێ��wc8:uݳ�ug��+l-�R�K����N�"�6-ckD�$���bk|  �}���P���P�}�B����@����CB������T�СB��H����Ѡ
�����@m���d� ֩k�����+�&��;)�*R�}�ӭ���-j�֭�ՙ�I-�*զ���5��зirؐ�gr9]�\���ݻ�Ҕ4��rpt��M7\q��]��waSl��mt�;iѳ��%m�"�Iε��B��7T�*ƶ�i�[0j�f&�������GA8}y� �q��F��k��gh��.�Xf��^�ݢ׼���ѱ����@���h�K�t�+��u֡�t�;[�;I"�)H�ֱm_׵��@N�pV�ڌk@P��λH�5+��\��>�֫�n5�n��J�V�)�A�v�
WG1�D����R��V�V��]�����Z��C׮��kZ��1�SMMʻ����T�*��۹X���w5k�;j�͸�_Z��\�ƴ(+�㝴�7WXڵ�#m0F��mB�e�׏MW&���]��P�-`�j)wsl3\�@aV�*����v��u�1�|H�S.�)%+��s�T�*��楍��cf����֭��4���ϟJ�
Q�ƺ$�M1ŎE.�T�������R��C���c�o
��Q�� (R��+zT�NXo^��J���*��U�%+�xZ�6l�s���[5f��I�  Y�*�J3����tkܽo<JԔ�^��T�%�{ۀ���y;�U7ou�T ;�y^��
���x*�-�z�yD�<��l�U���DZ�m�na��  =�=�����< R����@�U�垽�H�/�"Zw`���JB�+�x�i%Vu��(����=�{�*zhWY�Wr+m'�<�ʒ��H�)�b��(�  E=�&��(1 ��~�R�   S�	�T���B��S@ '���?���D��S������]qXE�A	��]�����,��y�ÿ䂠���}u�}�h*��"*�j
�+��*��APEaE=�Ͻ��G�������V�肛Wy#� tQZp�ңo[�]�&�?9����JݖV��U���:�6����В�V�`[N���jr�Tm��hl���p�oM����Cr�7�KʙbR��1#��Ku�f+��f3PH�սM�7-�m��Z�]�Z���w�.L����ʠ�����%pls��M�XӢ�TH-�e�����H�u�B��)��E��@��k�����WP�4�g$�{f��8�k�I
ݡ�(�@6�h�r�h��d[�b�yt��aD��*��!��¦�!2�yQQ�����&�϶��qd�)�Zj��GR���r��c��]��2�)�O"i��<fk���f�̅�ڲЊv���]�Њ��C4�H�����1q��� .��AYP��tr�[�AM���76XԬҡ�H�NJb7�3m\\մѤ���0�=D�
��S݉�$�6D�̻�)���*�K
A��T��%1�
���55��1L"k[e���-{�4T��/*hy�D��Ym�4�]\{���ۆ�(a�t��zq������lJQ%�Fj��I����bA���j� 
�a���y���3[�5�Y�����&���ua��
L�i�-�v�mAY�R�!��=�0<��ov���R5��6�&t�^�)��P�ڗ�@�Zqڔ�h�R"�B��]j�am�,���%`�N��N�ӡ���]h�'l'L5����� A�4ЦS15Qڐ]em��<`�5y���d��
�o"����=wu#�Rav�ƫQ�Pwp��R�#%lͨ��vb��S�m3�学��f���H�z�GkY�+4�M�@��Q��Ha��[�F����B�K P,��sd�v�<*�sV�ǀ-H�?h�k�B��2U鹹���I��$�r=�(к�)�n*�S��W%x�^���o��!øt���6:KN�6���1Z��m�WoN5��*�M��4!����ƭ9O4mHJv�w5��\܍�F����h�쟖�e7Mܲ��"Ӧ0%��TكQV���b5{���u�G���p��j���3Z�f���ZT3
���H�k��*�Jځj6�	!u�ܛ���N�*�Yt�e+��g�-���1-2��J����Q�WP�d��0�Dvm�O�D��4q�D��KM!Q�v�1��H[F�[ǅ��k�mCv9���f�j4-,��Vl`����=��Sw񛮜��v���K<���n�!S��gB����ֵX��;��W �iɋ[�E]s]oZV���L=���b豺�i��q+묡�Unޢs@�t�@Ƕ�ٴ
��ldѺ�ͽ�e�5�K���B��l)�����ddMuYz�3gX��[,	Q݋z����fMݬ�t	Kvf�Hk�	1]7����Z�+4%;�k���>w�dς@���;$�k����Gn�M�x/��ҵ�ۣnؼf�,��#w��J:4`��"� Խ7�u���[D��lL��Pn�4�4�� [Fm���gI��fV֤�����Hұ��X�v�+�v�M�#�nJZqg�Q����4Ï����o&�6݀�{Z9W�V=��h<RJ��E;�����َ����ޅ�I�]��e��|aKV�
i� �Z��X���NG�A�[%F�XΦ�z��KV
[7Yu�n0,�r^��&s�h)S���8팭d�a�����z��(�+)�+6I�f+vLO4�V�ϵ���oe5��B��lWF�!�[&��4��b\8��ʰ/o2�z�%=�X�(��6)�-�������cE�5�q'��Wt��ż���]
`)�5���2)f�-�)�x6m*��r
r��2���$"�h̬�5[�x�8U7B]8V-������9�\pf[��cM7c2����,r�Rc@[^�*yz�Y.�$c�1p
��C��q�Q�cm�ЦlӼ�N���MM�L	Ssw%Swn��2´/-�z�/9&�T���t�kknl)P�Z�y[i=��7@���,LU����oN�4vRP�ġ����*V86���r�jÆ�e�����5�{���ܽLw�覶� H�
	�$��*^U��b���o�,Q�j�H5����[��9-����Q�/ll���[��3��.�\
�,�Zv�f�9-��������Ke� Xͫ�6��zͥ>�u�ܤ)ň��un(-����w*��"n%,��j�I֋�T2�UaI���[;1����{��$Ż��l-*�l�Q�JXwA�#/t���<�.I�$�u��"�u�oc:*ڻ�b���`ɖe!�PO)��\Z�C�66Z�'�Ab��3V�Bh-�צn��(Q^�U��Kw(�'2����:ؽ70�N����X�^��_ul�$Y
���u�5��[VvTCoa1�$sH|M��z�]����eU��z�9D#W�+
�4�B�*EZ�E\�1�,|2M"�@�ܣ��`M	���M�[C2��!���h��H�%%ީF��pn\�zLL����Z���vʠ+u�YVl�&)�k�˪�C[c]��H���1n��ʁi�,n�5#'-����Y��,�9�5����t�vEWW�,3����t��L�{d�5��KIġk��-L�#�Bf��Ƌ2���j=�Y������5bs�p��q��B	kA�Yc@�2��t��.)a �2�z�֭itm��'"��VӸ���)U��G)CuwN�P��6�@����OS�ו���tӔ�UR�ʖ"-˂�n�
S�V�p*��7�]�V���Y���ơvQ����H!�;"��fP3�LK�`�uu5QG@�gp���íV���*��k5��Q�PX��U�D�j���2�F��i1����{�!��@�R���c*#Zۺ�`U��ma�H��4�"��J�D�[��M��HA�R�so�.,�f3PZR���%m��[)0 1��,%e�����iaW�C7^�Ș�6�5w�X�˱Z�h����4��5m噺��^��Rȱ�2�ׅ�.��a�BFC
+]է(;�j'�o���� ��"�)���%�oT�0�0�n�w��&<�/1শ��^�|��ܗ�0��-F��&�J��I��SX{6�7�m��G@���]�m�6jL�n�AAU��r���m-���+i�M�,���(䁺;�\za��j�����hn뗉��Ga�v�;� m������Xl���}q=Mt�7^���00�%L�C.m5�����Sh�O+6�jT^�iV�ݍ�((���z,-*�M���Iܘ����T廻y��kG�E�J�
������;V�y�N*�I�䎅ԥ�f�ʹ Tv��\���F���cbQiS��ɗ&���;�XrA(]�݇LI|3wp�[4c��u���8Mr�ZE���l���L�E
EJkE�1yB���eF�j��x�]�ݬ��+N�ê�`HZ�ց��v/`�л�Co�Y%��B����AR�oH���sD�hmP�V�D"j�J�"���qj\{W�n��6��/]x��ݡw*d��B��GH�����Lڭn�M�P��#�F�9*Ye�����1nm�9�6��Yʻ����]%Q�����/F��c��(��F���ZE�4�v���G'��s-F���L��D�uFu��h��ˠ�4�Ê6흼�l�65���f��K�]�4b[���b���iP6�v�\ј�����裶��ܯ�hm@�8�źL��7j�e�v]�����C�]�Rbk�2P�u,:����MS��R�죀܃C���pǮ�ͧ�+��4��y�+2�T�E�J��Mؽ#e�V[R��&�åd�E �j��V�b'a��e�Y�3B�b�Vo �k;v �PK���al�(��[��u;lS-��=6���6]�%V�f0]<�:�*(�O]7z�Hч[�4ѵ��cbfdƝ\�[����ӌ��n�FGH��f�s�����v�bQ(�����Hu��Z�j[��d�5Y��=R�=��Ǵ��.:R�d����6@�(�$`��!ѧ�IIF��!זGe&�\�!�� 4�Bm� ՠn��j���Ԥ�@����z�}5�nV����n����('1�Ӄ,��XL�K۩+�p�KU��c:���+]`��%@�2�M���x�`�lAY���6�-#q<�-N�	N�2B֮�/1�X�q�C�v���ڇspe��6�fd�g	#��ݰ� ����n��a槡�`��0��%�N�flǩ���fتʴ�a�S��#��͛CG� lV��9�SM�t�U8����i%٫v�$�������Զ��7e����㴀yd�7u�$) �^IO�a(���J�
KJ��&�3��E�b��C����;��.ʰ�E�]���Ø(��L1,3�����k�N��:���:w��:Y�[GU��Z\�0D���`���V�f��%���Ȯ��CN�k�v#KBy�B��wk6ȷLZ��9Qڽ�S 2�Lkn1.'a�%k F34:l��A��a
����a�x�-?H��eK���4�/tb�N�o4�ʄɅ���MD�0:�7�:���Lй A�zS�0�v)S/^Zw(̪[�M%�Wm�Z �]�[�FenT��64U��@Lid��-P�I ]E.���fޜ
�J-��DR�\�
a����)̀Bm��9��ܲ��Ř���8�&�m*�>���6��o{�P���]�o(�t������C��"�6����D���6�f�($�:��R�wY+U�*�-��S7V�愉�B(����eܖJ�p�N�2�]K)����a�Ƚ��%�]��cc�m�%0mVR��e�")W�?�7>@���;�B�4/X٪�W��a�&TA�1Mݴ��1-��t�i*���֚�#Iǿcv&
�r�SCX͖T��n\x+,Be�Vu���ݗ�䷁h9
��X��b�dXB�m�.1��eJJ�H�P�6�M�Hɷ��t�������b;T��&=��{V�릨�.֊i�4�����1����Ӥ9�e��J9����AiF͢�'{����M|D0��-�u3t���ǰ�����՜2 ��,����1��cn��A��A��S�ݪ�!���u���pfJX����E�F�����f�*S1=����mǯ5t�`x�&#{X0�3,=�5�k^�4�Rbe��K�k[�Ffa�K@e�y��'�G	���v���cBn��kt��0�lكB[��5̬�Dڻ�wP���Gu�j}�.��[t�E�kR��I���8��[,���JEY�׈��wO���yJ�B���U�����Zڥb]X�
�-p3SV�nRZ�mP�3kP#i꼲�C`��d[׃�~�JfjT�+��/���J���{�Q��,S� E��c 9t�V�(���V�X2�<o .@�$�56��`2m�imG�F���P����v��%&��d=*f�&A���s\W���Bm^\�"��NQ�r;��<�T��t-�p�������@�@�v�Ř�1�,���� `���f�wZ�J��^��cs
�,���kw{+5��^��0�Ԯ��Dr�� �SK�<���=K�hY���۰�ҧ�kWZ
�o���A<se\�D�Vq�i*��)m�#�&�k .��1�f�!'��TᛸV��K3]e��T�Dv$�`9���(a!ֲ�D���u�,wt�8jB-�Qݺ&cnVi�l=���vƩwY���Ա�[zk1�͜2���(�d��+��^��z%�����["�(%�fj9t�I����r *^R��Iv^P��-e���5��I#��V�uXK]�����43.�a%�b��������RQ9H�
K`�t����V�w�m�ToC�tl�H�;�}�"Φ�o-�'3u���F�УEJ��w�n-�U X7��n�@�c{�o�#�^�W�W�naA(#�da?hW�4U��� ����,���tK��k�Cr
����s�f� 6t���7�NX� �"�>/3Z�!"�]�-�lZU[`Iv쭗�j��� h��3�Sr�=T���Jqc9p�6��i��[��۫�Qw�=�:��XT��W��q���X7�@Q�/�v�e\�����ѬW�o�[�i��ma��Mj��Ğ�nTO*�!�ey���E���u�a�z���^P���q�@����Li�)�E�5��,�24�.�3���j������j&kf��*#f����]�Z.���2�D���FacO̖ x+j�TZ*��PT�6�4�%���R��E�V���E�7�zsS]�n��^ce�[�7��N�,�Mލ�-�tLN�4d7�e���-{����6�E=����ݍAWH��M�x֛���0���<�Mʍ�1ȩVfB�ҡk-��u��IS^$��2Ӥ�^�WY!�i�O��ݖ1��,�B�\�imd�q
M��h�D�2�֦�w���f�����30T�{���n̽�p,Eа#VT4�1'-��t���8�\��9PVb�ŢK#e�v�
����ek���!��c�ٰ0A*�95m�X���8�ڊ�0c���6f�fT���l�8,�r����%�����E�&{�W���[v7e� �U�`7E��H#yHl�Q^��E3��t.Y��T%]�5pn
ۘMn��A���hQV�'�r67��S�����ѻ����[GZD��K�7��p��Yw����r�"��(�J{Xm��-��|�l�xd��B^$����X4�g�􉹔݃��]�9�j3{��0�Q�!��z�V�{��W��jU�����Y4��}f�)��Ķ�jI�������V0q[�-/��3D��0�i��3�w��&�����8�V57&K��/UX��aⶀ�U���J��A0�W��0�9�ːɔ�X�T㧲�L��N�l��2(�TѻΤ1�nF��WVd��K�G���µ^����p4�B�� ��5���#����	,��j,vp�@��U�a]K�+,�]�;+�*��h[�CA������,����yI,�{�e�R'kV"��ۚ��<�\)��j���ޫ�Mc[ə
j�����W���~�,�U9�;�1����m-���lŻ�`*�})w9�N���9ԂV��%�蹿�42�C-.a�:�ʖ)Gy��{�(�]*G9\qm�i��Kx�Eb<�*v.L�e�7/#z���|�����a.Cln,I��b쑊��=�:݊�7x�!Ŵ4�:�b��M��؆�Zr���v�q���I��KU^kn"V<ZY�BG��dm��M�#�`'L�=�Yjin�)
<����Mqʔi�k�:��G��&���^��[�ΐ.�o����wen�S�r�>��k4O7��i���p)�-̴�;���6:��VWRI҆��뷮4i�kC�Gv^�R�1�� �F,�z��M�V��An��W`ll��ީd�d���Ҝ)��m��wڞ� ����7�(��5ut��oKaIF�S�p�1i4ޘs0	p�&�������%�[Q�:L�x)���՚Nk��-�Is�mhM���u�x����R$�aw' K5l��j���^qP�%b�!������ʫ�<�q�.�n�lyD���8^#m����k<�:�a�S=�*a�R�x�*�����7 vRN��X��Ӫ�m3+"��M��GHc_!ۨZ�Ҥ$�!�VVDwtL��n��
<̹��h�U7�pj�x�pGQ�5�.J�a��֎7�=c�5�����Pū�����n,5�)�"f�d��p(�sj�FY���zk��| 0�`�usr�^�/F�X�L��K�Tz�VmK0�)
᯹0Gĺvw`�r��9�o�2��gr��%wwY�޺�ד]���m���$�U{�k �u-U����N�+У�7lR�Gz�����ɘ����oRF*�HI�t�m�����[-���v�O1ֺ�<��)�:K�C	z3x
P=��׵�t>9ZD��� ��%��e����/`�J�ld-8'-�
��.��X�iы�6����H���1�{|N�:9�[)H���Mx�l��v�F��i�'҇c�m! 7!і�ǳ^Rޔ���#�4��x�� N;*�T�")�;��]b�d�j0IIۖB��v���шf��$lrxH��k�FX7�Y�VRN쫙y\zu�C��
�6��t�Vuդh�S�,�4n�:�ki��̹]0[:�z�Λ/��u��¢��|�rW|��ly,V0�BE��4�бx/2WZ�n��T5"c���D=�G!��һ�OPo�Ia�.��O>t
�\�N��Lp�Z3���W�4C�Q������;��*x͋d�GD[[�ؾ�F�:C���b��wbd9XH��tc�e���m�9U�e��!_'!0b�E��r�-�m�9��k:�J�2B.�Hs���ة�8/�Csb��5�yL-V�1rj{w�Vj]�1N��v�6�L'��6]i���8���h��05v��s*q����ͥ��]���PI��E�<�@��}y��+���>8־Ӆ*$�pz�ɮ�g
��PQ����}gw=�ɽ����R �Y�.���ȩ��z	k\i��S���Ct�'a�v�E��n_uh�|������M������uZ8u�鸥��7L�e��l0�CC1���R��Su����V-+-!� ղwY��m
lլD��l� "�Ʀub������,����}�ϲ�d���uނ��Xݱ����6m�7�y{��Z���Y\�V�e�L��WħP�o�&��� N�؆�7s6��.,<�Hu2�㘍op��F�(�v	����W�̩\��;��5w�m콣}�({m:�ڴs�+�6q�T�CՍ� �u¢�m�,|��Y�$��)�>ꕜ�-\]���짡��\�y;�肺���m���)�WRV�Kf�P:�F�R�C��]�l��<6�WRK�0�;/��Y.�h��j�t�Nea��1�.�V����A�N�0�kf"�p�i��y������>�Æo
xskUe�e?��E�����L#�Ʃ�N�,��{o�X�p,(r��@j3���SC��^��-�*�7�����uk�C*��md��;���܊��ZEJ3����2
/z��f�G_-�����!F�+�2%�x�[�����|�ߕ/AC9�؟YnP��L9�t	m�Z�%����M������놕���Q��.���v�r��K��
A/�k`�|�9zj}A.R#η+:a�v�(�N���ۨ�E��>WwP�<�ū&WNvT��!��:U�B�"���e�b�ӽ�u�A�ԛ�u>�.}�v��&���8�;2���Q��x�Z�ֳG�W-���EÎ+ig.���9I|r�=�e�O��잫b^���߱V>�(�R�{+T����B���;�fZy661��[�쐲�Q�F(�}�n��;�A��]�7Z�ٴt�&�x��=��[|�����e������K�v5(�a��]��;s��=�Z|2�
��wz�!z)���hTvNq(�v���]���fkD���f����Q�0����Z���)Ҝ{*_|*.ۻU%�r�6֧ilWY}���Y֋���b9x��ԻNeq;td����4��+Y�Q7B%iE1�#aϓ��w���2��j>���s�;�7`X��8i�0̒kk(��Z)�I��Xb��j�R(�՛�uF�}C{Uqڏ�Nsɵ��]�<�YۻR�ea���TQ#o�F�j=�&pVJ��U.n���F�Tq�Y�bux�d}9JhI}mj�����`�s��̲"UÖ��jw0ܹ�r;�Q+�鱹S�gf�K��S8�|�	���`��8�������4�����0�εVhRK��h�F����p� jZ�ب7����m�R�b�w@Ȫ��5�4����_Ad�ۻ\�3z�g4�`�������Bw�/ITm^9�hhgg[��U���R��т�u�)�Y��1�R��]B��]���5�Ml�s�.��[��wF�˨O+x��5E��Aár�;�;���͍�|���_#�}G\��CM�b��L99�O���:� ŷ+v��E^r����ڃ%m�
�)9J�&�����.�Ca\_�E����Sy&��_]�q:�en]�N'{��amw>͗�o��Z,�`;�e�G�l�R�Y�w��6L�M����.E[LN]����|�q��������eg#��6���L�i���;�͍�u\U0r�l�t��)=�sg�_.��t(�����A��V�ӯi��5��ܵi��7�qPf�UG���;XKq�s��U��ʴW>�:��A7V�i�ݍewp]Q�XEFh)�U�����4(���{�"[f��x���ݨ�P�4fKr�����m����%bT(��e=54�B���pf����ܠ�=��v쥼ؽN��@�ѬP��!���h/Mѷv�1�9�M�7��(�o(i��7�N��j�FH�(˨�-��lklB�j�9���*:9A���L��F�#��n��um4E5���H!�ҽz�K��w&R��'�����c;��G��&�[t�CE*��KY���`\uzxr���y� ˄�W�a֣tc��(��A�Ҙ\M��]��+l��o��$�+�Ҹ��Զ�X����uo�^˨wf���u�mf<D�-���������Z�W+ۧ1E�sh����f+P U
��P��ʹҫ7�I%�<t���+R\WY9V�YGo����V��HV�p�Mn�ֲu%Ԇ���]�E�ٸu�ä��e����i���"SE�|k��������=3~+�:�-���;�ڣr�:��u��;L��ߕ$7A��ʼ�Y��Jw �~��W[�]�Y[�b�}�+��=8�D.t�Q���x�=4_O�f�ePO�7 ���+R���1��C�����h�	����s�hu��)>d�y��1a�-�Ѥ�Cv�ɷ)� C�,����W�U�ɫ���� ��R*��k;%GZ�O3\}uӲi��,�_q��b�s��DޮLHӚ_At��H^�� ܲ��d�Ǭ�;"�-��N�^sa���p�ý
�qe վF$'q�)���_�6������E\.�Ma�@Bq�n���4U�؈���9ݲES#
��j�ܯ�wM�����K�Aچ��{iJ��v1y�[�Dqκu�薁�zP�%uE�74���J-�w"��s�������&z}�nӻ��f���wp�Ŭ�믰�0�4�"�h�:����sovFwj�)�樬�+�����O��[;�ײp�����D��ԭC�L�,h��[�Nө��"���Hr�/N:.��O�ˋU))�����_N=ţv�j�6�m��n�w֪XFp��0�I�����x�[��'�T0��e.��sk��TA�l]ӆ��f= ��:��r�~�]��m��k�r;�ZH�v	�Ii�-�4��יj\��]ĵ}յ�Q��G9�����)6���*����֓���.8��&�Y���>Z�/raކ�&�n����9]�fjo9����M�%�(� �{���4�m�E�0���{�͎`����e�N,@��a�J�e<�X�[�h0 �-5ջQSK��
�}!�;�f��ܻ�ݖs�ܭ�5����N�c��CS	ۙ�a��V7� ����2����L37i��Fc�u�F�*�۾ۦ��	�Vc+YX�%Z�` ���@�9+��^�wȎ���!�/s�;�t�ٴ�ׇ�&R�g,F��CF��UeV�I]�� ���T/�i���8� "[L<��v�'�Cc�O�J]����8F�C˜[��O(�	�$z�ab�$��a�up-].T�u<
'�F}���i�Wx��o$=g*puڕ�� ��6�����Pk�HaΕ1lw�nHffd�_S5�N��Y����U���G{���u��q��1�i�K��F�kDSn�^��.Z�mD9v��^�mQغ)*�]�q!_,Ź�ݸ@�Zϰ����٧yt q�ȫ��(�A�_��R���7o�'`cv�S�M3w���������E,=|�V���P�a�ݡg��p�I.�+��@�F��n�k\�q�Y�����z�b��Z���/&��3(���XT��n�Ƀ(�l����+8]�kq��R��4�R���91�y}0�:BZd��yX�tr���E&��7Z��m�
S%v=����u�5ڛI�
�1m���K3��t�x!n锢��u�w�lA|*�FZ��R��1#�M��9M�kBk X����vf.�w}Ȟ]6��Rݮ�Z[R�/,:W� �!�����u�*Lš����mX\�.\&�Ԁ5�����(T2��C���L���θM�ьsr��Z��WL��S&8^���}M~EAww:��<���5�Jʃ.��=]mm_7���'����7��-�6Z�v�p��Y�D0䖝h�Y
�M�i"�T�b̢�3F���	7��]�.�S"��M��$��ei�I2�aY�s-�
b���za�/��Ӧ&5�|eq�%�_jϢ�գΉK���o�
/3��6�u6[�[���,B�! Mڋ�ܘ"�]O��cZ&[V�yd���&Zf�uڞ��8r�1LrQZ�z�Vz6Q���vgQ�����:��-6%�%��70�R�"��3��:�ս��K�Ɨ;��v�v�T+��Ϋ��ӜKZe��"�_Xr�~ �����+�Y-�>�==��[��w�>V���J�1��'/�tm�����t�Q�2����	3_ۯ�9ܹVr��e�G8N�W6ҙ]ȶ�68�E����7�/1/?�mO <4���Π�"�j�OfQ��c���H释w2�m�#N���R[ب_9�b�v�N9Yݸ-Z+D�i�v���J��xc��{鴛�ӫb� �[[���u�]G�]�|�s
��T�k)m�Zoe*�t��vJ�n9��Ҭu������܆�ۈH�NfI��Sao;�x�:�z��z�ʮ��s,�<#P�	����c�6Τ�M ͧEٴ�����h��k�QE������^� ԜN��nl��Ů&��$"�{���I��;C&����耫ʬF���ـS�i�Q�`��#��(��t%��֮t��+�sh՘�1��u�yP:9!r.�f��&�흥O:�N�7�Zۉ�T{��s�����!t�O2�ս�3�����n��Զ�ES2�7x@��c3�ʔi�\�6��땕���s�^9���t1	������6�{��GUHo[�����gauJ�.ob��r�����kX)94�eĺ_p���(ff��].vA&n&�S�Q�d���Kܥۥ�u���:���9��)΀�J�q�.������'-kh�yˌݙQE���Nd�����"�xH�3R�)f�)Wj�����3ka�1�V6T���KΝ�A�f'��洭�dr�M�<��[���}�AE?�
�+�z�5v�r�Õ����Ii243��E��-u�qq��)��A��#������Q���$B˗�.��4X�Ջ4U���ք]��A��PI
v�^�VXWi4i9���xƀ��O=/2�\��j�w��6L�g	b��sv�_m,T��6
y�����+T
�d�e�t:(�i�g/v����%�LC�Wl�ɤ]�r�r�=���5_BU٫�݅k�\S����g��>�Q��ں�b��dC��1��b�/��ĴC)̅��w�#y­�;)lid����s;��A�zi裇���B��*XX����g��5����l�k��̼����U��AW$�YE���!�����!M��cU�׆s�u�l]:��k�|�SՋ]��\1�0	@`c�����*S9.��V}����ɫ��Vo�jK�޺�Dm��[���v�s�
A:����-��f�V���e*�9`z��e��f����
à�j�nr��03Z�n��݊�b�4:l�]	}�3�ɉk&��d�� "�;�g��+_<�u�B֙�P�(�v�e$����Xj P)�u���4��b"����
u�-���Z��v�'*�/I�w��p9Xej/s1'{P�t�H�}�<�Y��r�L4��`|y��mK��9WL�f����$�􅴳d��.����1viqJ�����]yf�Rܣgj���ǒ��ʤ[�W{ק���v�t#.���W�W�o��J���3*e���u�+e���Ţ���8�n���\9�U2uι�Nй&��Vk-mެ�=MP�xm.�;)��[t�AZx�E��E;�㰈��K�b� �WwB��<��}&�,0�x:$o2.O���������e�a������|&�oh��e��Zɴ�kl[r���Os��M�h�k��T)�ʻ���.��j6����VQ�����E ,���3�m��p=5�ij[T�gA�)�vr��'�4���&��Џ�i*�a���*u��/N��[�E�)�E��Gh|���ՄȜ��ۘƫ�K'(h�\]��#�AR{�qq��̭�T/@����MS�x�+7:��7��^�ڧE�w9f�HͲ��s���6���p�.qk"�CL`Q�Nc#�v�ڜC�Pǻ-R�8���h��y�*gq�*!|%,v�`��[�o,���p�Du�Vt@��
�v6��
L����'���k����A��1u�%�����p�7�n%�yQcjeQ�F�U:��%��b�+��;ȝ	�&ami��[�ۉ��yYrq�3MЧ��p�JU�*��q�-��޿�c�֒ƅ��h2c!�t�����Z��#��"�.R�{�>Ƚ"��p��t�ٰ�:�|��|~3�P̲��N��i�����p�+^���,\f����KHU�݋��\�����Y`��^���)��b�՞2c���Y����h|�$+'1V	D)����y l�)�\�S2�):��tkr��X�6ȓ��aK�w;���S�EҪ6/�}kC9}�H�]u)������b�΃J}��LH�VQ}+������*���ՕU9��sJ����i!�]�.�X�R��n
��l��Ъ�VdB&��^���ͮ�L>cqwQ�mt���^vJw��[��ˆNG]n�@|Z# ��������+�T1���gF]<�C��-�m,��.�[әB��̧f��ec˜f���Vx���*�*�Oe;��q�g��k&�	�Ǌ��nme�����%�)�Ѯ8ʳ�Tϸ��+1�bM��,l ��F -���M�/2�)�M���y�٣��ۊ�"v�1��IS�7S�m�6��y7N�T0\�D+�j������&��Q� ]��`V�&�R�f��zl<��N��Z{:����#�t�P%n�G�wSS��%k���s�
Kv}9�f��
Nu^�R�l�'���T�,k���,ʺ[�L<.Ľ�\c�	t�e��ԥKy��	Μ��uÔ����֋�i�����D3x�O+_�	���.�ФݺXƹ�6� ]�l��Z��n��)�|&�c/�zK=�(��u�.G�q=���E{mh��N��v7�t<u��c�����M��_9I�4��+'��[��`�Bu�o!/q��Ki�a�f�˦�Uƫ*�`8�5A��+nңb��]z��h��_ ��@�Y�J���<���� ;3v�N�-�hEe���;���U�����B��2���B'7�{���+���hT���9$6�e�#���i�6f$��=]�4Ru�7"ʗuR�x����x&U��&�X��F�=E�1bf�����jX��n`�݂�-�-�F��S�fξ`έ�s�]�&�Iիvk�#�H�k�{�+y_rU���e���źF�<:����ۧEf�Ӄ����%�ʂv��}��*�]���O�l���φ�¬�^�4M�l��҈�L�68CEc��Q��w�����KqCD��s��OY;J�'�o)gQ����8d�N�+��Y��(-Ԋ�.�6~S��k(��
kl��wI#�\7D�%5R��!���M�*(�/.���[Fo<�7+&���:;MX�)�
Bѝ���dҹ|���Vsw�X#�,ǯ���삷fԮ�,�'
�:eedze�q2�:�1VQ�����-ι�(AI�w�Z$/�b�Pp�d/�F`��Gk�9�V~�ZPqk�j�ѽ��
i��T�R��`Ed�HJ޷��ȳXQR��\�gfR$�	;�A���2S4�ڼBKG�N/M�o��S�[�����Kp�\`y��$��%�1�	X��|hљB�t f^^��c����Yy�jf�j�٧��6����,��OY���[��9���<�n]�Zjuf!��!̂��M�]&�3"i�}%��40�!�]�b�ݰb�8�fu�9czj!���(�0sh[�V�ͺw��f�3[l�Φ+mS�Z����)��-��3#M�Xtt��Sv���v�P��']><�(�a*ﲍc��Jרv��y]if�9������}�+�0v���ޚ�-[�-*&� ��эjr��o��&/b��.�J���Թ-�n'�� s%ԙ���B�^
�]µ!���/th�$)K�d�v ��B���O6ۧ9`�k.��7/!�\�	q��i$�
�+���nPU�BD��p��5սW�G����I��\gL�۱�-��4-�S;G59�f��4�ή�6�I(oMXk�}}�\�Z�CL��#aO�6��;���ge����8��oo*��r+ ���WW�&&^`��M��݆�b�{6�,WJG�c��y;(YIsjQ����{�յF;�ké�̭d[��:{�����MH6%ԭ}�3e�y��\�J�N<7x�5Y ��+�w
w�f���4��W�Jǒ����{���9�f��v�6u��-(v�ch����+6���˾��Y��S�?��*e7��n5
De!���*���v	��nk�j�X�ۼ��N�넭h�@�����Ô�Cm�M�C�6���XC�@��+>��a����8e% 4�p�H�����at͛���VuC��7����1R�}��:�]����\�U7eJm(MqR��4�Zݷ��`V_�+z�GNe<� S��de4�g;�C\�����E��H�AH t|��n�刔���f�0���{���<��R�ǻ�3��S�'�_P�}�b�@;6I��|��S{֐r93�oB%p�a+�w����t�1js���v�&���+���Ӣ\wj��5���rƥash�`��E(�,m�<�Y��!Z���peo�噭�Uu�5���哮��a*�Xk�4�l�!�>�Ӛ .鳏��B��5�Nμl�*��f�G�è}�I�{��f��0e���O�Y��V���N��YC�g��Ct+���76�fd�i��x�q��-T ,����:ֻ.���%����D�p0��u�m��ͳ�jyt�bo��+Z�p6�AS��w�m�]Dv,,���F���Ս�;,cȠh��ve�CJVe���Z��V7��b���I.ϻj>���F_��F��K�nr>�y
�w7t�ҧ�-'���i�qd����W�u��^o����/4�^�S5c��y�;�w����W[Z��izۤ�έ �:��n�[����P�Fwh�qc�0��r�Ĩ�O�;`p�:�;�'D)N8�t*��qHNgܐ�4�� �Ʉ�'c]�Q{ܧ1���YĉN���Wf�JӷP)\��\8����(aҶ�[6��ؠ��2�P\�W��>f�\���Y�Y���7�T����%�)w-y�>p;uuvoWgR;����y��|#|��apW5�{�K�ą�Df��]ձ�e٩c�B��]`@0�ܱ��<��}ǘU/��yy;�Q�U5��؍b��_Qm˝��\�]��k��M��%�[O�V꣸3����:m��8ZOm>f��bamP�E�2���W�H��u�e`5,��9rHVv��C[h�y5��r��B��z�N�q���4�Z"����b���޵XWn���8���ͭ�]ݰV�_ڧ@kF9��X������hD�^5���ژ���rYÓc�ȽL=��Nei��������@�K�;�x
JL{a��Λ{���lٿ��u�s�kU�
8��!J�,�;��iZ�)gp�#i�7��)�d*����VHm���뾬[�V�
�V\���:��}f�Pi	���2�����m:ww�]t�{Z����\�ڭ����]:Om=
�Ѵ�23mCdF����0jb�7f����31���ڭ|�+�r��ݎfi#z�d5�m��(�n�� ��[a�c+Y	�2��-�;�[Y�Tɛ�S��so�`7�kiu����
��%�X-�������Ad��µ�U��w���mod״��3Z!-�fS֧cOV�r�lT7C����닮v��&���1����������J��:����7�`�zF.'5f�!ѷp1-���7�v<.VP�gju[�^�4>Z� ^Nw��n��ǽ\8-��D�m����p���۹�I�51��Gt�����޻]�H���u����O��h��"(��� �Z�[���;���;&���KGhܽ�\�?;75Ӂ��>�Y���[�]ys�6�ǂ)�mv���p��6�Y]�5+�k޺�}�cw�M��	�� ����`�I�N�':�h��3$��]�+u�T�+c�&��V�CX��gr%;�#�oR�D�0�U�2�W{�[j��\wc���1`;�r�)���[!�f�'"U!YLu^h�[�s�j�B�,�MjoN�����]��@�!��4�R���h�B�D�P'(�4��Lc��<ߙ�
�&~x3j%��KyФ5-��yC5��{���AG�PHƘL�o1�\�ėnĸ}9�F��k�����vJ�,��u����M,�-pb%dZ�y�����5����tzl�Ѳ�B�w@h��gU=ph�I�̈́r�*CY%\j�J�զuT���"���]WB��Z�A}�:���i��-㵮�@h�� �T��ή�%�;�ԡf�Ձ
*�1탴VV�*�v��{{q��g��)�Ut
hګ8��m.Pg< ��F��+�AHV���D�2]�=.�
t;&�/+UJ��Ɠ{�U�m�STh �]Bi.{�s5��������]m��u�e��i��L�1�-�a��.��,�UY�g2S�MR�� ��suvj,ޗ���좬�Ƴ
FKg�|�b����^S��W��&�'�Y0�pϸWD䊜Wc�e�ݻt�X�[*�� ��wZ�A^fh�wv
�a�+�m,5�K}z�.(��s^5e��c�[c:a/��Y��$"헚��M�{����+���Ú(]Ֆ5�.��h�j̛3�r�}�8T1�L�:�biv�,��h�.�Yi;�����RVI����\J�Y�M
*X�;��˵c:�մ>���x��K�ї����0y`Z-��w0U<j�Q�t�/A-����N�,�ם�g:4~T��f�4��^>��؛�z�A�\K�n�b�֗K�Q��ԣ�Wd
f:�)*�u�͎�H�-�v���mY��mE����Ts��2>}�[M�tc����M�����vX��n�O�*ƭ�7��{yԸ-�Ðn��p��N �&��S�e����m>@nm#P���:������MUۙX�j�m�o�@����J'�M���85��\l�59��ج�(U�Y�veC�z�d�y�(������P359t�E�L����(�oM��*�뭤���u�K-]�p��5�+�]k�4��|X�;��Qb1yø�4���'V*2�s�3];�9j�����MY���6U�&�@ՙ8��͇]X22H�1�1b�5��|�mv6`�3�Z&,c�
j���H�	����}��{��2�Q��w�
�',)[��!��.�����to �:ՌC뱎�K(g'c
N���l�i���@��r�3��{�L[m"b̒���:>�Je�Cv��r�v�oZ��qK`��n�ɔ�Hb ��F�&m�
E��9��<�&r�[�J3fHq��R�5�*��e�@:Q���ε/3�(����Ȏ���V�3�C<*����QZ���u|�Sg��F��+/8��ny�-u�G�+HW0v� ����pe�K.T�dEӟ{����ȯ�	����+YW@"7zt��L}��:p%�z#��G������<�nܽ�B�h�������3�X/\N]���K�(̘s4�a�\_#��j���7�U�j$'\
�m�ᛑ���1�����kc�m����t�U��+(��f�"֫O�[�����|���m��s2o�(I�-so,a��Y�N�K����NE6d���)<C
�Y��X����S;v�� V��������U�Ty���WT6q]�bl���֡)��g����鴹�T��������;6�b-#%;{rܵ�t4�J͎^+�#���M2Z#��&���<�r���<�%N�iƵL%�ށ�-�8T�8Ӗԫ}dU��R�:�ƨ��)�)Wm/���op!f��p����]�u�]�f��WҬ�:���!ne��nAw��?l��d��ZE,�:�[�k� nQ��:�(
;YK�M�l���CH���i�튻n��=� '`��u���0����\�{�gq7D*ڍ��hZ������3j+#bg]�V�=�<���Y�Q�k9Q���1�_"��H=�F�/�t��l��ǣ:F��V����6��;K���W��/���)�v�$zv����m�����\j�:��w����e�eT&�c�8Lu��R��h.��|��U�Єt�n%�������5_eݞBծ�a��*�9ދWNu1tw�p��G�������&��(�(��
�!�j ��*��"�"X�r*��!����Ȣ�
j�fB����F����	���)��ib((��#3
����&"+1ʉ����h2L����jf���j��h�b���������)H���J���� )JJJi(
B���)h"��Ji��b)Jb
i�� h"�hb�Y��i�bi�����%�b�B����(J��(��)Ji
�i"F�)"i�`�i�hi)���Z*�*���$)Z) ��i���*�����)h��*H�����&����)J��b)��j)��)"ibJJh"J���� T��}�ڪ�6�uą�C��G^�yT�,i�ep+fu�)؊.6��W�6��cP��A4p���\��O�,�Q�I�%��|6�WcP�u��b�*�ۍ��
�gU.���h��/~"]ܿE��Գ��5]���c�ș�;�Pv�5o�וO<�D02�csOA�\)٬e]l�u=�%�=���
���^�����؆�+U���z�Y�#�)��h���t��<�E@�G�J�gI���#��T̯p�N{]��?�V�o�@+�k��Ń��6�����\�I7�_3�Y�r㶐�\0��+�#!��<�cvT{:�cZxPw[n;��`�l���k���$X���6iPX����W���I߅���e*��Vt'5�4�EF�U"�-uϒ���y���tC��Ԛ��@%�9ݏX�䊇���m|}�����c�-Z���d�鶤�ͫ�V�U�3�N�FqtW?�-U�]i��f����\�{Go3⣝�⩖Y^��GM��f�cz.tux&&8�I��\�z:믜o�xeu�>%ѫn�=a�ۼ]&����uH^�����/�D!���&�V�ƺI(	��<�Mx)K�c�?�5�"��Ҭ�f��(�(�,�4��W�eLZ��閺¢�[S���ڥ� ��uW�^9O7K��͟O�:�'�0�
JK�	�����n�x�:�f���[q��M�.��&�"Wr�-��Ov�����jB[�cN�8ͪ�r!ۯMC�8`�K]�w��*������4x��$�^p��ߢ�"^��cy))!Ɋd���r��FtE-uÆ:j�pl����<��N��,�xGe�D�gsv^뎧u ��@�BQ1>���t��LZ[P��1ˤL\0"W6��1�l��n��Q����g\H��v�H�J����t�z�+�����*�K.����&_S�ʍ��P6�0�B���T��t�~@��tb�Uׁ�U<u��C��%�^|��q�bK�]��ڪ$Z)�'�7@s�g.���OG�YC�PJ����+�O����I�L�k�5�U�MWbN��s�M<�'[�����< �f�t���D�ݐ�}�Ue�
��GZL^l��f��/���Fjt����z��a�=�a�C��y�k�1"fl��$��g� �rc��(`9}��z����_��½��a��C��&�N���[x�5���[<Nf��xk�*�D��
�����@	�I�F&4�p˳�ߢ����|̸�źU�\�`r$+�,R��O�Xf]��^�t��_���ʱ�qt:S�zueZ�ݗ5����FO0^�y��>��Js�"A���#���R��52���{����X�U���J��1^��p�sY!�%�/8�C�l>�_
�v��ևUz�3�|2��.��QO6�f��Ge�zō�.�k�'^Qmgw hq4Bb/�p�1\�}�xVf��X��A-uO[�U|37e��@�|8�j6�3+���2$Ë]^w᪘7`2��r�YMߺ��阎: �$��(	����q�)�c{�aW�,8�U�,�_em\�	�B�lz�HfA`3��M\>����2���6�{��*3y�J]S2��˦E��h�F+�.���B�Ա���h�C�8z���T�"T<���U�ʣ�1s�9O�ԙ�'�*�n	�ef#^�P���\:w.�>;YJf&�bkF����sb�քK}0F)�%T�q #��h7Ჸ�uY���<�^��u���suA��S+�t�lΈh�{X�w�]y`���'��-w�� �;�
R��V��N��`�վ�Z�#�W%�[Iu�-��(.q���S22��S��� ����g�
�v��9�����1q�i��C^s¤�$��-��}�]l�2MGO��3��4]�M̽�մ�Y�=��Q�0�ٍ�I�f�B;�WZ�m6������6
U[�d���;�l����F\�!�2�.�n��nW
��2:�J��4��j폶p�+u�i�V���f�t�W!��6�Har<B*.M�q����������Emg��Y�{�PW��!p���q2�Br��^�s��Ζ�á�3��.�m��c���,N��G,童}��lh�6X�uLE�'A��3nvbp�Q�.�����X<\B4����+����7Ur��{��`����,�ѷ��G�zv���r��wze���E�����/Ew�]t�p�ѿ�_K0��pR��M�7���u���-7p�Us,���ߓW��Z|�Ŏ�'\L��g����u�^���L����(�Y����jr ���b*!)�X9�2����U�c�!�M�kc#�v����p�Ă�����4��R�鈴�3���
�Y�ߗa�,V�Y�$��x���_��*>��������>������|&ˇ�C�(`�5;w:͛2�O(�W���楇b����+bǟS��Y�PYq�Ϫ�xwP��]�IɡO.��#i�٧}����Z?MߦՊ'��N�@L0�W���[43��q�h1���Y���љ��b;�H�\�����t�LV����M�Q|3��6��U)&.oW97�S"F��pin��T{�}e���)�;��et�e� �'X��Y1Y�xB�ѱDZ��v�Rۋ,��������ݧ����ۮ��.��&Z���X1TQ�Q�������1�[$F�<w#-�#5�2��"|�=���#�d��Js�w���������1�{�Ô�l�^J�์P߲�U��y�q#������.:]Q���C:�[��8���By�1�����x{y�0�rՖr	�D�f��T�&��Wmc�p ι�����*�LL��.�dD�&��W���A�>VC�z��%L����O)^�ͥ	��w��xs�X���]eA Ub��P��#��j���<�K����Cj���m�iF�u36fj��ր0?gKOg�ʱp	��OT�p�}�ԁ�VF=��)Y��"ٵ�a�s�ֹ]C�w�9�s&{�D|���&��{Ij�z�Y��c�ҳ�׍by��?^]h��o�f���\�o:����<0\���К�j���lh4��j�Kr�a�����Ov�޺帱��*]T	E��H
�ֲ�uJ�ȇS��{��f�YO����{E�\ۢ�ώ"2^�X� �bǵ3�sXd�����V�����uM��U���|�tdO�,��w���\F�L�zr�i�%���w����O�w���$:2��Zͪ�dT�N�ԫ�5��弋�͆M���/�d�G�Ͱ��Q*o�oz#�'X��/��
���M@��b���7�&���P���\Y�g2�ܐt�c�lơb�W���o�����K s����'��Wu�oj������]FK��~�MXm�x��'��U����'D QX���h^)�f>Ւ'�n�eJ���A��ۄ�5��g�މt�Pp$�<�=uӍ�2\��AK��\�C����u�h�ib�ֵo�CRY|s�D!���P(d��'���-y1<��X���wwFe�=���Z˧>��9c����Gc����_�º먁�D�Us#(��oK�ih� V3�DĘ�$T����3�*���5~��e��N�����t��F�ν2x.��4kܕ�8���7΂�h�Q��A���t�C���D��P�9��4r���\4i={8�g����������!.��m��e��޽󗴃t�-�b�Qփ��F9lƒ�]0V@t�. !`J�Rf�:Q1@w�ы�G��w�U<u���>�*60�0aVi�yˏxz��?�鵗V�2d�&�y�r�p�$�t�=4rP�׷0�i|/�ZĖ?bi�.��󮳻�]�,R�n@+4)�+F�g��F��}���]�����v^�������-o6�F�Yg��]�6dQ�e
9Q�楩��ؑ[WV.*5�b<bEƸ��n��K��G�)�V���든�R`����r�#w���{�m�g�Y^AM;QT�&�s�MC�Bu��<���e�\�k5�mf��v�%J'`ƍ~0�ਮu���6Pw4,1|��FF�AY�ǩ⼵Z4�rL�P������,{�v�g�a�����0�� ��Pţ,�3��s1i��:^�w��α�7��]X5'���]���~3D�ԭV��0*��gw�Q��~U���w�k��/�>�,��a�&���+ұ�YX8[TO1��T_d�D(�W�%؟�K�v���\g�>V}c� �1�y���0���cGz�nN�RI�'��3�N��8��)ژͦ����	\�?F�Г�ו�k�0vz��Ȧ��"����R���<���庼�'-���6P!���r�E�QF��P���lz��t�g������i�r���T�w�\���^!6Q'j �A\�E��H�b���;�C�K-���c�8z\��"L$T���n�71�9Ȑl�N�X�,��>�0�Jt��c�Y�׸T-}qW��}�U��綒o.�q��{r��R��n�d	��6rQ%$������m�B�,`_di[��<����,_#^ ���C(��虡��\�.�Op�Ӕ�dB@������	ޚ��s�ېT�T���2��5�u�:�b.�Ɏ>�BH����'v��w�M�U����#�� 4��Əs�lj�/H|c5�<�؍���njj9�Β8�tCg<^����؃1
d��IH� l�{�WzF�#x��jZ�;iγ�8�)��Ƶ���s!���/��ҙ��9fc����H�5��HӸ�{�|]��5,�Z��)Wt�7�N�;s¤�D$��7�F��5�ْA�"�l�̩r��9��O����c{]f����\�����'�ۄ�s<��$���F��NK;A6'��{q�]E	��b���[��K�0�8���Ƚ{k�1�Z���]�8��r�#��[��r���n���S�JE궅`�n���\�{�-V
�sWx���΅G����T��&y����gt��hvԅtעq�b�b�6~�4Z�ՉiU�~{�� �o�����6}���}p�%W2ɑ�l&��q�zhC�yS�0��XYL<*�}�9�n�z>~�=YgFDt�;,qj����`{xN��V꯻�°�Z�i�����*L#� �d^�Pݛ�ivV=_XT�Y�m5�9��wsp�U���Y]��\�Ļ�3.�p���9hښS���Xd�*7
��3d}L���ed�����ьq�;Qҙ��t�2�t��2Q<�\�:v:��N��e5a/�M ������lu�gFBQ��"�\�Hk�^X1��{=N�>Q�m0t�D�[����B�9�x���8ǲ�V�מ΢,y)UB�sw�=��������Vkq������M�N��'�GIT2��ڶA9Bhx�|��s���EChL����Cu
��*7��p��z^Ćr_N�Y1� �Dp��^�h�=W1n�G���;7��n��CZ~�q�S0�i���x�F3(�$�8�D�!���ท`M\*����,W��9H�E�腽\;!S��g�͖�f,F�n�r��3"��JS 
U�g{'a������^�D��8�hO)�3��<=���C!�VY��Wף#8�Oq�=�ڷ��z־��դ�����:����lwR���z��R�k�7=X��1�61��eov�1LttE(x�t
�ϱ���U�Zy�[Q���ԕ�#l���{g ��΢���4�.hC�ᥓ�>�Zz|[����{���4�v�Vh�{)�R��Ɏ����_)SZ|1�if�R^��m
��+���-��N��5X�RR�r��-�[Y�^��ǆޫ��+W:�8��lN��9��R�u)^ȹ@�n_Zgc�'u3�����z$f-�(��k
Q9���V`�6!6���N�r� m�m7�c�ɛ�h�r�_�d�o��rWQ����3-{�w�9<���a�^"�����5���C`�`�p
5�3/GWy���q��ȴ�BÔ6�(���d����z�C����;�f�K9
���Z�)ڎ���9;�q�x����Hxg���ms��`�_+L�Ȥ��9���\Mu縞H�
��q��s?C��Q��:n,�)_�������Ƥ�{mP	dwc�1�"J�gL�wpԉv�*���S��b�pxLV���������s���W�i�
%!�Td�+�%K�݈wMŰ�-84C.�&b��Sjtw@6Lp@��2����V���tqCK�-� 혰��0Q�X�5�[�jK/�i�{��d6�6��_�Ș�64�l<kˇ��sl��q�ϖ��<�צ����-v��r4�,z��aSv�b��N�΋�0�� ���BF�*�5;��gDR�\8d:j�a���{[���C}&W���w��/�
�h/CL�%�`k��7O�kw���J�/m�ؠ�A;�p�`v��G�rS�ɲ��ΠoNi�0����d�|��i��U�/���i�V�7�1�=�l]:�Y��t�7X�Y�bƼ@�gH8L�0+�%��@��N=o7kR����e��Rŉ���C6����B#�7�*U� �����ᖆ2E��r�g�	��o	G��4��㜪��`C��j���uN�c6��p��#M���ѕ�E;�&<���o��*T.��>��k9R(ٮ�n��v"G����n��OC�C4�ޡ�V�]���G��'e��%����'uU����L+��i�|!G��� &erfl5��+uŖ���Y���AЩ&��9��!�Y�q���2lJ�:�4�ᯞ��j+�e%��A5K�v�䵅��dH���*���e6V��Q�eX�o�eX����q:����h�e��:|]��k�l���{�#˖��]�eվ�����h��Y+9��m6^p�p ս񝜚z�q�k��&��`ᾀ��>u��AϚq�=�2�r�������gR�u:�ω�_�<�v��g\@�MV"@u7�
͎/'tʶ�	���딹کqm�(�U:�L�,�!
C�ںs�2�^2C�i=�
 �u�fӦܻ�}k��V&��v�A�ø����n�1Krѷm�c��,�۲�foe��C�����fĽѱ�����Ʈ�R����<�h������3z�P�V;n��g��ȺD���o�l��;�>\��2�@�e�T�7"�q��R��uM��;(����Xn������Λ�kJ��<�q:���^εO	��� ������P�IM����7�3~�Y�v��X@��?�^��R�Ꜷ��:��m�:�<�[���	ۤr�N�ź6�,&�A\�����U.��4��\���ɇ�Zy�jg2�9���w����w��Iz��)�
Ռ��NLثjm,���S����M��yYʱ�I��*�샒�qX{$w����I��5�*s�$�0��U���W-9ۗ�`䕮���&X��r���(G�g;*qbw`��Iq���*�#���x�Q���;M��m�1f�{������f���<u�RVm'�Y�[vr�׼0l��e��E���#���W�0A%Gx%�)s�C{N NJX󙛤L��ӗz�����M95L���B�ig0n��4ҏ�i���u.��u���uo�ۊ�}Յq����Wj�[x�:�%C�)��a)��裥C,{ۻA�W��:�����:�^N]3:�T=P-��Ǌ��e�� `�žq*��I_L��n��Z���M�=�_a�ѝ�n����9�7>�U��l�OD�D�)�̡�`�����j8��E-��J��L�� ���[6�ΚXT�&o�^�Qn6n��y�f�}��QB�DC�D%%%EST��5@U U41!BRP�%EQBRE �HPSL�ED�-4MCQH�HSJR�E �P�DRP�RP4!T�HP�	E	J�4R��%4�4�P�E)HR�S�!I@���4R4D5T��@R��P4PQH4�MK�)#IJU4M	BRPBT@R4��S4�)M	E@D4�T�T��PPDSIKT��D�U$KKLLQ@P-MSJ�
P%5A@��U%R�]3}�3i,���H���e�W8���C���.�ǧ&�������ur�n�ʟ|0��Y�.��`����u xz|�C2�����W
�����E*RP�G�dPd}���f	���f��Q�Jټ=�/^����t;��\����P��>����t��dt{�6�]����g�������hw�Wm�J���l\q���������!�\�Q�������3`~��S���%�Z�}���U!C���5���X&N����:�C�jν�n~���{s���%S�r��nG*���j�@�5A���;~��z0q��[�5.���#��\�<��s]C�2r\�2�ϴC�?A�`�N��u��RR^X�\���jz�ɺ��޳��:��9�οp�=��\�T�$�5n���PAUc�*����������u=�};A�%Rvs�l:�pd�f����[�W�sK��L�#ۗ3��z�%��u_�u�S���%�j_cq��u�a&TWX}&�U��xj��~oe�G�>����.u����:�����>]���?�ޖ�C�:������)�O��sgrw}�+�kKE#Pj~~���'w���h;���ԇg��瘺��5UO�7[Fn�ʼq�v��}�����K���0�O�r�ѣe�jK��^�>���u�;y��?A�%�^u�]��<�=������)���mz��M?O���B�^῾�̒�qe�a���:>���d|1�8���p��A��O��5A�z�n��J�����%���p�#�uN���2K���������:��uԅ ���[����A��~�Y��MpG��{x���1���Do�7=K���#_�4���HS��}��7w����ju�y٭���?N��Xr~��J��xw��C�����<�Q��f�@}&I���ֹ��Mh�$����+�W�UdN����:��hK�俣~{ͿK���w�'s��\����������C���<�?gf�����9�#p��?�����N��������m�5���9�;{� }�Spj�������}�˒�5/O�i���]s��{滄�9.}�s�5	w����U>˒�y��ݩ�.~;���K��FK��\�wW_�ߗ�9��D*z�,+�]���={����3f!A��K���Y�̥���4b�K��<0�:�mm�_&l:��J��u^f�ݮ^��o`rf�%�uӅ%��a���lU��;Wf��re����g�ރ�wH*ۘ{F�����E��P���k�"ϱ߸&O�8�������n������ݩ���9�����h7<�5�zsz�#�j9���b���j=���A�%�ޱ���Hl�5�G�!\>�
}_,Ӄk�D���V����θ=I���>5�{-���3���P�/�;ڹ{O�h��7�m~�:��&G��s��%�����l}�� d3K^�j������tE�y_�{�=�gpj����A��sPj5{N��#$�7����<����׺w�����k�:�������g��\��3��kk���.O>Ͻ K?}���p�_i�T�c1���k���u>ڇ��}�0L�C���0:���J~�:�I��5�0(
(9������26k>����u�3�y���{��Zz���s���C���CACH��1�}����lD}������:�e��O���~�/e�k�y�7���t���:����}�����7����3�S[3K��}���\�fy���ɨ�>]���i���ٟ�����+����#����<��A�%O>�ǫ�>�R�y�;�!�G%��s`yO�sXw�5�{��2r;�&��2F߰�n]Z��5dn]@}}jr2Jr\����߳�o{}y"c���|<�U��|*>>����j!�3��i��rufy��#P��\�ݽ�'pjC�s[��2A�޹�7��j5r/�7�d�}���wn��hMY/����}�ƞ����|�w���=3GS�\��0�/ӓ�r���>�^��:���K�~�-C����u�'��s~�$�w���������ո5g9��G/��]bn��|mq�������˺�|ǐ��Cޑ#�jk_bW�5	O�~�u�pj��6{/U?�����GQ�|�=�y���_��>����P�]��6��}`�7���1yn7�^��_����=���}�z���g���;�~�[���%t}����r�:<���5&��:s?F�)�=��A���Q�uw'pjO^��o�����=�Gp��%����.��?���3��g;37��ז��kZ����N����m���F[��c��y{ԡz�nTV|tX�3�r/�o_�޺�R��r�lvħ�a��8Y���7[V�������д��u\�wx�,:Zu�����<�H�(4F��9�@۸w"�*h��y��3$({���%���|�s��.@j���05%;� ߘr;��ܙRu�P��A�J��L�`��<5��yBS��u���y?A�{�S� z4D�{~k{�.�����J�w:%���>�@{�.>���|<w�������;�����%\��5�϶=��%���wO�r��#d������7�f�N��ZCP�=ځH� O������h���}fYUy���~����5!��Z��'��5}�����h����l��.b�w���ې�亍n�)똺����4A�%Q�v�o� �Fas��O�r��">B${�${vʿ����fi����y�]�C�{%�T�����W%�5�	��]h�^��Ѹ?k���`���:�O%ʀ���ny��乬?s����Q���Z}�BS�y^�"���nڟ���d������9��Z���[��������ѓܝf�>K�~�.ӭhܹ��
z�?A�d�Z��y͇Sܹ�y�nJJr\����#�Ԝ�*{������8
 ����O�^�N��r����߾��\{�����f��#P�u�����y���U&A��l�4%� ��h��@}=�y��:�m��r]gPj��~��:��2��}�"Ǵ{�xo˘��������&G�_ӓ��9惨us���u!C��թ7��2}�3�rj}�K��:���jM_OA��%R�F�Ñ�������'S��:����܋����Y��vX�E� �4��x�f1��U}�6�{��C�=�A�Ò��;9掠5��W<��w����}��uR?tX��Q�qmNK�����x�5?K�����w���� �������f�����ԉ��G����y�λ�L�#�5��6?Gp���|�j=��5���O!��?A�sBkXy9��^�7?������;��S�sY�߸���!(�(8֔z���K�|��"�x�y�;�������9����5'$ʾ����5߼���'�>������B_�i�������hԟ��:y�r�-���F�w%�`l�^��#���e���ޙ[�-D
k"-7�-X0���z����&���ӎ�4�Z����@b�m�c)�ӈn9����D�c���f���b=�[v�|{�|::kN��˽ZC�WvF�gh��[��|$���s��N�X5D�sv�o����n��X��*��0�7���s9/���\�z�K�tK����0u �b��~�ʐ��}��A�`�'7�C�ܚ�F���i)�'�|tT�מ�cDQ��G�=Cg0:��	T�\�A�yP���]O֡��f;��S�؝������+�z���������e�OS���>��K��~�s�rA�o5�ר�G�D ��ʯ%��S�!�1p�G�(��^g4�~�3���Z�BSܹ�o�]M:�*��j������[�2~�$�f����%=o���y�jO�^i7S�r�N����;���0>�����xA���q����\ 2����.�ǩu���'%�f@t��nA���k��bw�r���Ԕ������jO`�35R?G������x&O������#W�*�)��v�ŉ*���q����\|�
��=��k��>؛�<�'���A�%�}�l;��e��Ϲ��2L�[����擸5	W���h?Gp�C����K�����Y@r0���޳�w��l�9��lq�߳~&�$�~�� x(\�]C���v{�[y�����=�5<���;�{P�K���B^{����}�c�q:��)ߘ���`��>���\�Pj��9\�).��PWDR�V��z#�ďzjz�k��2=��֧�����7~���HQk�5r]F�����վ���|>�UBu:�d7V;�-�e�a4vm��G��ו<n�3+�a���QW5��U �`@m�̌���J ��]�@�ܬ�Y���I�O#�$8�k�T�,����مGY�5��� s������	�=�����w s���S�����������m�2�q'I�(�?���#k+��x�L��z�6!.��`(o )�/y����)�I`����%>��[ �����р�����cY����Zr{�����ޑ�t�ȕr�H�h;F�|�;����(�Z��n8t�z����h�Gˉ
{}*K<y9�^���52P��WUBp9S�!�j�&b�*c��u���l�U�<	:O ��܍�3NU�H_�m������)Uq�3��4�&�Z��<Ԗ_��6�u�M���d�A�2#^T������P��H��3~����ٛg���Ӗ8`���Gc�Z�g�����MYtp��V�19�]c�RQP o`�"b$��EA��P8#����5~��,k��V�M��8T;��HjW���\N�ϥϸ���-&��y�o�A��.���]�X�ٛ�龔Ӡ�[�ͼ6]"b�5��.;��0Y���A� ��Fx�vȐ��;�XH�g'��:�b���?%Pɦ�p/<0B�ȅT��t�b L�1qf��ú��.��}\�8���h��\Ry^�mT��)�&���9�@yv/�Y&c���mP��NuʝI�K�hC���Q+�';m�͘Zj5^\,�N��s�MC�Bv۽��[f�R6���c�i�d��ں���4�0��!�<�	�pv��/��镟oy�5Ŷ�M+����$2}��h�4]i͘Hv�C��c�U���hgq�O�V@5�����^^�{���	��z!{���/�k3�bS 	�3��{��0��.jSz�O�l�Z�.��r�;�2�W��fs��ZT<�Q�3eM M����.�9Mr�{~+�*�B�vT�����A_r0�[U�.�����	{�^��33h[�@�{9#t.vwN�ʹ��h�Y����iC�n������
.�$���W)Ɛ���Ws��e@���d��0�6X�{7�W���znLHDzˬ��~����MNa����5�������!񸃲°Xd�y��-ߘWG��mםAzZ8Mf�h,�g���SR�����L�wN�����ak�.���,�e��NS+"��h��U��p9�lS���Չ(�82��� vz���좍���+�1����ș�C���X�P���w36���z�e�́�*1]Av��
�R�;e���z�$Of��:��8�pfe;6lچ������/��4MO̮/��D)��f%m����T[�Oi�p�9O��t�����	��2T�>c�R�c4��1�����NѾq$F3^{½^I�GΈl��`�� F��I\oƥ#��ee]��ί{�U��ڎ�K����"*Яy���jḇ�/��UԲ�]F�VN؜<�e(�Z�v4��>�lՌkݔ���[oS�.`kHJ����۝dYl'��!M�q�b���XA�,za�M��o�\ۊɾ.�@�S�"*��b��ߢ#���Db���@��*z[:7c��cx�k��l�,�>�� |�$�L>r�q�Ǹ[r�d�Ϯ�}�q����y�(���/�Ҵ�s!�s¤�$��-��{2�H06��A�ɜ��Z�jw�^�Y=�}�-��߲=��Y�|��r��d�,�N�33�[\4q�5M6���.2/ ��X>�Z@�j�1�U���?5�T<+�*��(���M?7һ�dCgN�T�^'A��u��bD뺑�(���3gv�\Ee4w�9�^\����y<n�>{�,<S������&K�3��y��LM�E�	�s^���%Y,<�je��ݤ��#�S��f�  �*�>�5�ɯ��v�>�C�/
5��ki.�ueC�0f�'UݫVg9�Jt�Ζ�gFU�=�*�� �f����n�2���͔���G&<½�L�k�����T������Q��Tm*��4��,X���_F��[v�M6U��څWk�?WW�VCO�5�������*>������USa7R{A �V��0i}h#E��X�xw�&�y֤�59��G$c�ǅ���f�L�ڜM�)ìZ�4�dPr�rLl�i+˜U%�%��(gB�9$��fw3 ��9;�\u9�7%r\rWrp��X�e�!�@�0�7��o7��>JK��QY3'�ꯠ�oH�ׯ����a��o�ߞ��։t-]CĞ�c��7���fd�v���Zx�;�XG���Ϸ�}ç��k#�n����\����@E^��ŮuGbv��a����P��.�mX�*���Y�<L!�R$F��n�ˏ9�f�L�"��1`�1��sp"�e>[�=�v�g=J2���q�R��CP���)tه ��G ��ۨ��Ђ�eǻ<��M4zw1���Č���$\D�]4.�T1��<=���A9j�,��eۚ�h\���K'�7I���r�qq:�U=FY��tyg�����VCɰ���W7/�uC���vi�b�O0��@�!:�#�'`�t�5��1�ڿ�P���q�%
�<O-����, �e���9Wu�>�P�	����FU�K���[��A����$���8c�Ǥ�W��k�9;�9��T��>��g�9~0�p��V��6ew�ur�xs|�o]�g|�c�<���~32�9�~W�5�a@נ��������y�IWu�FE%�R��ov���
'˒�{~e�g�&�
�S�>��$T���}��3��u{�E���g��1Zʵ���8��ʍAa^L��)�Db_Q����M�ǑRu�{�|Њ�����?�2���kMJy4~�z#ވ�����p����1�cC�8��P�,��v��/Z�c<����u���狳���t���k+l����Y֖����p���N��5����_\��R>�=�e�)+��^-k��;�f���v��á!�{���k3'=���ɛG1�¡q�O)�=�C�Ú�*O7=��V�1Y�����< фO����R���}�Z�n��.�#b�~�5����Ξ�!����3�S�u��Q1p�$�lR#x
��M�[���=�S��@0���*�a��s��X�5վ9Ie��>Ci�\!q�*���]H;�{ݒ�@�~p@���Fo�e#�6�;u�,p�p��H�#p�|�Tujv0ZB��t��[c��§�G�Ԣ������C:��n�qZ)���y��Ɔ���k�.����ͨIU�8-�rWo�����~UƇP���I����~����=�b{���j�=s&��%���C!ˤL_�)��7޿]'F��F��i"�v�2�luiWCSV��RB�����eޥ�S�Z�6��=�cvF���ysAÞf�0�{l��JH,�o��Љ]C+j{����pK�^ߚ�F٥4Fc��&[�n�έ�\ �U�K#z	Z�y�� ��Q��\�V^�	|)b�n�]Y�٭� }�������f�Ӎw�!1�ʡ�Pۮ�L���ʛ�o� eX��^��i�����`�Vkx��ntT��9Gt������j�TZ�ɓi��x<�b�7ѵ
&�߯��fM3�i^�ł�mL??N=�/6ai��yp�'v�k>d����^U,��d�Y@e>ۊTpq���f ���F�t���A��A��:}��j��3*�i8���Ǯv*kf��I�w�y�c�vNư��s6��ʨ�]mW��x`95� ��Ŭ_Am��j���hze�fq��bᩡ�r5����iT<�����ϲ�.�.��QSSݕ�yM7|��UD�����$e)�ɸ,E���j�E�\�7&2"��ƫ2p�
��v�ʳ{{�<���n�QN�n����A�aX,2j�e��y}��==�z���e���<h�7%��y� �76�����ٙG�n��Z��1��-9L��n��u|9�q'���r�X\qB��$�*�p:�^;s�u֩�맯����� )���=�=s���P��F�MG�t:� �m�W�M��1�Iq�/���\=�X�]m�6��V���l�W�.�;B�8!=�7:`]n��N�}�/wm)�Y*g�����g�;�hϞ`nض+m����u�Q��9}��b�7֕)�pV�@S0��n<�/��]�X/�Rꑛ	Wu�����]��$Nh���8R2sy�k�F��
Fn��i�]�2E�A����䥎�.D.���>��RY�]�䙤N�Y.J�:�����|�s��v���V�
�t�t �^ni"�+�w|	-f������
<k9L�C �ОP3[I�2�R��.LT8� ���C�`6L��h�I!���4U��[�G�`7|K�SV�ٌ��7v!��C���!+IQQZ�|;8W9�bU�SZ/l��tR��v�P6��c��KpfV=Ֆ.�����J	��cr���;�� ��'jelZ��&%x�&���e��:�W9��+2��cmM�l�ꊌ% ���j�E����b�)El��7%N��d�۩�..m���J2-N�g��/��N�1��D.ܖR�2�G,�O��4U��q��ʰ�)�t	8��V�ۋ�쐆���u��;ZC��H]�:�u<�X��IQ�s�0Q�2�޷#�Z�Gz5\o,����Z������`.�N�K�ʖ�Ŝ�组wB5�x���hL�b�R�ړo.�Ɋ��)V���RW�U�{������%��w#ڴ��u����S��Ss����t��⮋�ذ���;׊Kf���B[�3��FEYFc����C�ݥ������*�F%2&$p.�4�0 ���rǲ�W�b�U��-b�\�0� ���b4����\kS��u"T�͏mNױV�uM�_�K)�W�{�Y�ޤ��sWIe'����t�i(��Y �0Y[�5��u������i�$�(P��	`��b��055_�޳�P�pq��!hV�S��&T,���n��_p�Gx`}���b�=l���Ϥ8��wη:�a����'��!��E�d��6�!���`&�мǯ4p�����crVk[�X�Qn�f�7�]fpDo�]�X��.�
KVI�dڗv�<�vt���N��R���\nO4F����Ǳqh���p�(3�!(�eʖ. (/v�����)����x�Ռ\�S	5�ă��M^���5 �=}1:{�����V��x�aZ#�ܦR���|Ƒ�w�8����a�rKU��:�����Dn0ʴFU�@^ӴJc�"R�f�gt���P{��Π�Ɍ恵�����D���mW	���DYVE��}��PϢv��nvV_;Ƌ^���|�̊.o�Z)0��fYq�+@�"�݋��z�wv4�(�ebƛ�t�u�*H��ݩ�a�!�&]r��oF)`�Wu�qfR4᝶M뢇����o��Jii"�����h(����	��Z�i�)@� ��)���"�
�b ���
 ) Z
 h��B�)�)�J�) �V�*����h���( (ii(���
���hi�JQ)R%B��F�h)B�(���h@��������O��~�,�e�l�]7�F�M�3�V1O��r` �c�9nɮ�ux(b�ٮ��q�s��fwV�sP+w����`�k�U_U}_V�E���z����5��C�b�P��Q\�d�B�U�o:��v�ı�3[Rݗ�R�a�7i���p��9�*U
��F���0�AJ��#�V�1Q�{2Z�w���Z����u�\�q���>;��M��#\��S%O 1�{�Λ<7��ޜ���V��"�ǖ�RN�8�tCg ���7z�͈(�W��V5n)sG��)&.�|]׼%�ǞaZ\e3~���5���71��%��{S���;~���F4��U�z�u`�sH�h���+'2:&L8I20l�=)�0�n�uFd�y>�G�m.�8	�l��~�J�L�h��hW���~@1hn:�����M�o��ڠ�"�',	5����9,����$>Y��ĺ����,)V�X�T5�a���щ�fV:�M3']Ԉ����3gv�H�Sُp>����kJp������f�vձ�z�S�4TCWQ9~�����/��\��6�,~+�>}���k��Ωq>[��\��4Tт��=�@;�M=�����!~���k�l-�qd� M�U��gCm���wd7�4Q�Tx�&�c�|�V���8r w��w$:b�e@�}�ѐd=�K�X�,�Z��e\0O��u;lɠ>y�{��z0�7n�����#�����o7)b��\���eV���J9f"{\2��d����&���PCōV0gq��o�rt_�+��z`Ö��_q�����]Tux^�^Ҟe��鲳#��|q8�I+ҕm���V3(98C�P��t�~�!���TY]XX5׀��4�\ѹ|v�d�����]�3�����KK�f����-J/)_��cU�H�.��l�r]��c�hE�@M^�|&���!�~zn&�GE�#�$��1��Iȡ�1m>0o�3
���X�7���K1/g��v\G9���!i{�#Ϻ��@f�̾�|z%���Y�8��0�T*�j���V��\g�ڙ�;Nz�#�-�#.�3�ӻ�vr����g���^�Diƹ��w?�iL��q�-���
��c͖�As(�yԥoN��Q֦h�p��P���>�e���5�����9W�J�=u���S���nީ	I�J����S�pϫ�*h
�Y�VQ~#+�+I�~uU��݆�h�zjh���)���k]<2����z���<U}�5�sN�
�W.B���X�3�w� ���P�w=�6�U֪酝�S�{�#�Q���˿��ܯ�����Z�ī�f�tB�y"��M}7��i����YI�D�Il���DD{�R����Qۤ`��Q�JY.@jtDX�A��Xw��EJ�������7��t���C9Of��;��5�)s�a�5F�  �9`ix�U�v|>eU��D���T�\�&ǆ����ߖ�°�a��H0�d��b�s�X��̵p�r �ʟ�7{��e�y�ju�Պ�4�=C�+|25Н2�.��a�^"�S����5�foyw ��V�\e�A��/�X6P�b�0�d�WS�}Bx�r㶐�d1�uJሕ,�XA_��=����B{�=6��b��;U��\
�<S���5��`�/�[(߶���R}�5l~�<~��=����m\�ܩ�A�xϬ��f�����L�r;��ڭƪ�sK��<[�J�z�19"�O7=��V��q�Y��H�FQ��ۛ:�X��6�zWe�ĩ�&�1���w<9�ӃD0��Bf:T�d�h�LgM��65�������%//T�l�;�唝uR0�+�,�2�	�j�jK:/ч��Us�R�i��"�ݗ��V,9ܻ9� ��f��I�|NƜ��/��; ��q&�l���3�;�0.� )�t�Ѕɒu��1G�gc�7M:-N2.6��n͢�8i�w
0wG��")�w׹�E�t�N��ΗE��F^Yn��w#����#���.��ΞŨ�?�� x"|�E<f��G�j���n�5X�,t��}�벙�ɇ.�qJ�#��<=���^.QG��̅H�i i�咸��k�)�����AJ-�f�W�]�p3:X��t�z�'M��|�x �@�&��q�qT�SJ�w�Zרv5}n�rp��+�4Tsj��r����Mցn���,�P>H��!­Ƨ%+͘��v��5�6���r��į�T>B�yL2{ͺ�^L��ªRsi��,>�<RqV�����y��"����\T�3�n;�qI�{��Q"�JdɸM��<�Fʤ��M�������r� !ZY�w��">�tG�]i�ѕ[ɪ���S�C���?O���EȦ*��+9X��^ٶV��� �0�`[�
��ZL\f���_Rnk��;p�:erû�F�A�^����U<���n����b�a��0˝vPtr]AN�![��B�8̷:�>2/���ۺ�w҉ݲ���>�����:��Y���|�_#��Ӥ�t#��g5ّX�R>X��n�25��k��fn��<��_�'Kgwi��s2A��Ô  �n��q9�!�]�����{�֋�6�"7��;�5��t���/��r\�W7�Z7�l�ߎ|G;�g76K̃Y�y/��DDzˀ����`��ea=�a &;<��Ja�nof㚮�tm�䘪(�2ico"�w��z7��Q�I�ɿu�CF�찬)e�w��������s�9��-�������^&?�Z:޷����yk�(�,�0xo��e9���[���3�{;���!��tA�T䃴e ���Tk�nc<o�S	���|w��wv�blj�3y��d�L�چ����g��B8OI�(�dd� �C�<�:wyA.��;cE�IO�
'E�䶚1����1��J�E�(}^���
�s�Q�7�*�+�}L��7�'������nㅩ�|wk�|!7U�TF��|�H�p�8�*�n)eN]fe�O��Z/H|yo
�NR+�gD6CɰSu�?9��Jt�hv�ұ��\��� d�� 4]�#�.zW�e3cx�k�ɶ�8C\�%����cg���Q�F��t'y��tW'A�QJ�_�<�r�ָM�=�V��ߗ�2��qmy:�i�]_���7Ը0UL��v�ǃH����]qū	�N������`���#�WZ���29رN�(Zz�5&���u�C����V)��F֐��6l�ꇔ]l@���t�vT8C��2������&�#|��\��_W���C���g��!���U&`�;I{
%���C�C�ծ��_�9�M��ױ�/$�&S����F=����/�v���g���$׹�V���Y=C&X����YPZ�9��D� �K�q��ϭ&�U1�N�2�E��׍ ��Ч���@؞*3��a+\Ym�yI ;+�[5@w2�묵��<�[�<s)Ϛ+�]D����(O����'c���(��U�q�t��M٨98:ⲫM���%�#��Cq*��NE�v�W�ʣ
B�H������$���?zz�@�܎��c	}�3�~/��,���MC^Jy��Ӊ���]��p[��摫)�֘�S|b�g`C���@Δ.(�b*#iPE`�V�4��Ap���n�1:�`�Br��~p{��}1�7_Y�+W���EG���C�������=�����J���އ�����ӿ=75::���G �3��w݉�$d��+����r����T���Q,��}E�xy��b��Gi������7�PD��@��3�5tGb�z�>�8<���9O�b:�Ҹ��>�WC�;^g]�TD���A�@����BD�}xt�M�7�a�,��̒�I�%��Q�Z��բ�n�f�oH0�ϻ6u�$˓Ef����:����#�!l�}�����}��}Y}_}�Emcse�nP�~��F��BeZڱ�sЭ�����S0�i�nH���nŰ�#[ﲳb'xy�d�Kr{g)>��D�A���"bR�
)�#!�5�\;;l�@9����A�e(�7{x��Goz�r�S2)L���j|�l�2y�пW*�5�P燵{um���͓�y��o�hq-�d�J�k�1ϝ'�%S�e��GG�t�t4��uz7�Ȟ �c;��2ϫ�"�f��Q�JY-@r��DX�A<Q;P��;�����>~��h�u5���r���L!�{�E.{l6���a`,/�ʱp	�K'��a���a���猑�؇��p�ԁ��cc�/��WQ��:㓻��zX�>��T�,�=ROI�vɧ16�5c�
wR�v��}�Mþ�4��I��4ч�{mN�=
��؎�����>{n�~U�i�l�d��A��
�(����8�5��C^��ꛃ�����骕��OEӺ�V<^����}OS��kO
�
�
�z����`x'�	��\�I��YwL��v��Y�S�>�lC}�P"o(�%[n����g��'���֎�:� �4m�Q�V+~:0y �׵Q>�@Y���sr�$�����m*�Yp\O1i��n/�mUы�&�ax�e��R�I�ګ��E[v�$z"ֈo[MO�}��W�|��3*���À�U�d}I;�C�l��pP���n ~"�hg��u<z?G�;F���[o����gB���;@v��b"Ғ:Υ:��1
�W8��#��F_�@�Z�V���+}݋��ǔpXS�*a^�
5�]������yq�U�����y�.-��߆�z��t�^j6��0���S,]0���c�jb��kV��RY|sO��{}7{2z���ޞ�8{K� `��k�a	%#���ґ�-��qۯK,p�n��Ӛ5��ȇ3}C��e��F����:��4x��@���!U#]���{�����hǷZo�y����ӣ�JU���e��']��=w��K>B���Ai4�󌚐���o�.�v�	�H��禣�0o&�r����&�@�;wF1� �#�'V}���i����=\�"�_��Zk��^y+����S�ۮ�t�-�%U)3�
���*q۵ƕ�>r��0EY�*|7gI��Q����{~����w�G���c�����ʳ���Y�,BFX�9a�>M7�D.�td�����23&f���7�(��A���]>U�0�AGf a28�y:�u"��ZN��bZ�� 3G�W:�?Ʀ��|�xӼ���h��н�W�bȍ���̖�M�������:mw���c��LG��KA�
Oa���<*p�i�<L�쳠m���û,��܉}�=\�^#!Dc�gpE[,$a��Uʴ��(<���d6�`ٳ����+���l}]J{n
�y�O��{{Oݹ�� J�ޫ$T_nW�}���Q����%�]���dH6��D^��/��8̷:�>2/ܟ[��W�V*C�
M��=���~�ʙ;>:c�2�=b;<���a�Cm����u0m��^����z��Q��+ݻ�r@+���	��Uz����ɯBS̾ط~a\9��
B�*�9��ϔpq��~�$����	�
�j��_��	1P�הk�C��3n��ʮJw��7�06����s�����P���A�Ep
��k��\�xεL'�z�@(ihv��1�V���, �]P��ͳ�#��qd��@@�s q���n���V7m�[{��o*���(\B�c�[M��p��ʠ8]s�]t-,}^���d][�c��L���l��m1�ʓ�P{ߙ�ᚩ ~�/-:�{~����0�@gEn{�Ԯ�w}��O80�/D�җZ�(Vc��}v�
���b�';��0:��������*3���<��b�)�����l�5M��̧�z6�%fC;�ɯ�W��UP�����^s;���Lf��O�r��n����u�C���k�BqL�#\؜�Cc��fk�3g�� q�q�5�C��"+8��>ԝ$rΈl�{X��@��uT��t�"�[�ǹ�Cݘ`���l� �6xA����)���ך�r{ƥ׭9��
�~��{��w@�P�:�����*�U=t#�xׂ��04(�7�=�~K�1ҝ��բ����ɊԨ�p��k�F��6^&�@�g�j�x���Λ�y�!O�+�#��s�i Ǫ��Zn��L�3I�O3c��*A��d��]t�p��Q�F� o4�eTٝ:#��[.0�.�b/�̬u� �u2!}��c���^T��a�-9�n"�[�wYI&0E����m�cͧ^h�WQ9~����
"�������$:�ˉܮk��sc�,1D퐎�YY�3�pcMQ��y����
^�p���xY�1x���W�c�]B+�G)8p�/Ϻ�i�ц��i`5r�t>��Yd�`����lve�_+⵬u}�U�NRT]�^�qQ�J}J_�5���p�ͨ�d<gE�4�wF^�^ᔠ!�M����Z�PDh�ə����ջR�b
�+pW�|�3Z���vgr7;�<kE#;4R�_�/�z�<e�.>q�e-G�����Vf[f�Q��<s�l�Hް�M��Ht�r��%+콹�v��
ǦF�:�"��F@j$N�l��/�۠�R��l�,���?.U�:(d��,sL�I�i�=r�=��3w�Z�AvE|��j���H��oOoe�Nbc-+Օo&!�WL l�r�jd�,���b.��e�˛�Q���y�Z"�A9��9W�
sy�M|�9�M�ގ�십w����8s�[[�<�H���hQ���Y���[N���>\%[�+"���nc
�BrYjԴ&lZ/$���8اJ��n�k/Vͫ���j:�G�_>3�0�+�r�qh!s���V�X��L�4�;�tu�Z�I�~�lW\W	WOMr-�}6�~�U��/z��\0v������y��_b}�h����ӭ�����Sq^�f�w��h��팏5f���Cl%���=G����T�y����t���ĺ�˻����9cB.+x˃2�k���1�D��`e�x��;-Eu������y���kU�jq����2}[�{ ��H�b�-a^�Y�%N�$[$Ү7�Ը�ȶ�����Y�Ba5FV 6�ޔ'���=F��Gd��R$��]�ؖ��74ґ�`��D���#���9;8$�].B�ZY�M'f	(.v�����Ă�«/����\�j�'�Rx����u�hZ�Ǩx���E5�1��aQ����K�v��9�K��69�sE
!}�$ܔ�f���YR���&�,��9�%*R}}�o���v�����hkcFm=�D��/pS6N��
n���V5����jy�2�He:m5�cr����i�I+�-(��AWu��+P�7��:�+5�Tb��?Nm����7�\���x`:$-�Z��̤-��JZ{/�'�u������Ŕ$!7���ْh���^���ː��k2���i�O��6�pm�ps��:ɜ���K�r�Wyq�f^+�N��V#ӭ�u��9uf|�f�.�ަ���:�`�\�&0_+ ��ZM�rn����t�cHӏ�9M�Ƕ�y�h) M�Ò�[̀�K�׹���5���sm�_i��D�o�MJ����Śv�^��KbHr�,��.���ե�����9�٣cXd1H�=�o�N-�8��R<K�a�JZ�x���Nu}��	9�ens���\����=ߠA"/��f����YR1
������E`����)�<���!1m@�3������`6.����?�Y��8*�o��=w�~��3}y�o��P;�
) ���
��iJ�)Z
F���
JF���h(�)���
 �J�Jh�JZ
P�*��D�B���F��F���R`ZZZ
�
hJ �h�(�
J�JV$��)ii���)F����X��� �()F�
A�����뺪��PT�S4���j�
��^]Z_#g;��\m�Pr���� �]�ٰL޵�n2���(�Y9�v�yض��}UU�}�QXF�{88�۞=��[��<��½��+O�\��?T1NL�r�q��-�s�K�"۔�e:���1K���wJ���c�k7}�{_0���>� ܹ�����ӻ���A�-��#U<~��7�gL@�Q�=�8X�r+w/�z�Ra:�l�]w͊{>K���3�HX{�z�m��%Ӣ�n3s{�;W��:Jn@�Q%�0W���\���c��5�g�`����;���|UE5zG\��eCwT��2��A��G�K�
S�ce2�b1�k�z���g��+3��k^���{;w�N��4S�JwK.c$�&��3"�L�����P�"}'�M	�0�r2Ø�ņJi<4�j;��v�Z��x��J��_Թ���u���
a��:<��l0*&Uq�g3����WY�q�p�Y_��>IK%����(���"/�Q;^B�`��y�*�Nud�k.d��m^��^\����] �',/ʱπU�-#T�l��=�P�i�Q\v�R;��(��+�6�C��X�v\��3��"��ԥ�*`;1]Ǹe�9,������/h*O��u����Z008L��k��w#�n�]�m��ۀ��!"@�ۗeK�.��˒�]]��k��	�&�4���z��r��՝5��~�1fc�^�11�$�J�tӞ%��=�~ɕ�>vٞ�P]4W��i�=����~�Ij�K�d#��ݴVz��,��Jf�����=0��h�_��ZuSU�����5�����[cA�B]�!#'��|GM�m #)�ޣɠRUx�5*ٞ�B��{�����*t�# f_�>(TE\�}���a
<efZ�K�A�C��E�̌���\:��b���W:+7*t�D���?�ʕf���u�6f����(�����Qn�K s��nH�Y<��źb��ƚ�tv�H��u�S]=���X��Ґ�L�+�9>8c�q�(��w
9�¼4C-��f."Z�8uI�M���I��\�0l��E�NצPມ\WU#b���H���o�CRY|cuk�Ɋ��Pqܳ(οp�]��*��x׺ ����͍��f���<F�g,8e�pmh��a�궏20��c�P��B��� �~>d$k���:��i2��^P�$v�m�A*�ޛr RT�6��Sw�,�yg��!��)��EpW�f�3�}��bu����c� m4���Z/��X3M%am��	�F�R��
&W)N\�����A��e�"F;5 �)�8Zĳ�ƻ�ǔ��w�Rs��}��g�N��<;��M��5~��e��N��z�'xK>B< K��>{k8�L�tVs\���ܣ(��L_5� h�MZ�.�1a����h��т�uU�$i��;.��p�k�Ϳu�\�2�*7��h�璿1^|�F�*�MCn�XG#YB,Q��V��c���yb�rc�C�z��S�Zy5'������d�+g�[����q��o��\D��H j�|묫���#2�W�=5SN�w'��՞���r�? �b�S��K�u�W�p���.����vhp�,*)��%7=8�(k�Tlp�T�#5:�����V(W��N҉ݳ>p3'r# \�n��|�u�%�.;m */]C�e�fr����rއ��iya������z��b�!�S�g�J�����^6cA�L��>�\�F+�l���cپj�Ag�4}��å��7E���W�D^\�a�3�
�ܞ���°Xd�$���߯�Ͼ���)�|���+,�$s+v�a��L7mbHf��s��E3
ۍ$��v��ю^�q�Y�6xSFܼ%�3��B��:�,��y�]] ⺊k�WB�f�l�͆�>/f��]:XS'dPˠ��Z0KCSb���E�6[ٕ�������+&��y��pxZ6M~&a-=m��R�&5k�+���4�tnu�*a(�^�s
�c�,8I�w�1�t�ق�є��!S��,��QGGb�	k(�O]S��y��wD�q��\.��,v�5p��>�
Ã$�z� w9����p��uz�
I�De�<��}]}�1h���j�"5�ˎ:�B���S�8�]C��W�VBuD����p����*�;��)���t�~{0F��$㬰��b��N7����2� 3���n�+��_��^�I�G<�tCg ��
P�\����u��H��7`?)��%��5?"pǄ+��2���m5��ȩ2�\M�UY**Y��a�\p���OdX�!�\hiTR���<k��|f�4�D+Fb���������5��$v�E��*L$�-��M���x@�(��>�ي����������u�sS��Xm��ƾ��	:��2�',	3�_Ϋ|����&�5���?fS-fj1ڔ���,�GL��zb���̠WARZ�'!޳|p��25K��&�n��k�o#���:�*+/V������b�56�wwR�ng���Q߶L<��`�vB��j;�Z�jRH�1�y-*7a����(oe2�fj�}_T�|Fs����}��l*�eפ��w�c,52�tF'A�Nb�ìĉ�wR#q�Z�)c�k��\l�~F�wj�SFD`����f�[Iv�z�4Z���ǖ�$<]��.�.$�6����Ɓ��h��'�WSs>4ec'O����D�L�o��Y�d�C��;֝��_E
ї\�;��`u���Nӳ�*N�Bd̪��OL��n�.���X��;�	�X��T��(>B�.҄����m�K��ǚ�玑B���Xyᮼ���Cr���S�|cbeJ7`����g�u��H���3ܓ��7�{�=�.ϝB�v!g�7zZ{D=���M��K�hàR�9���J��鬓���cj��+]ĳq�Ϩ�Os��m����22A�c�_��]n�-^.Y���&� >����a��(Ŧ���43�� �[�i��)D�u%�.���!mW�s�&�є.י	w?��ǅg�_lpM�{WZ�ێ�<	��ʓo���m���\'ts�vV�
y��૱0��G�Y��f)��'����S�v-R��n�\�k0J�p]g}�y���zuP�F�;0TXW�%�Dmӆ���A��y���5����*n�����k�A�r3q��e�Ͼ�����S����1�v���{�B��*$jGuW���F���BuL1�M%����l�u]'�_P�<=��]l!��,�A1����/����J����kRպ�N S����x4W���{Ӭ�.�>�IS%�,rP��Q:��w*��ؤ��
����-N��ن6�j����jj��, �Br��й��CU�rf��z����gY�ӄ�|�4R��u���w�Lh�ܜܝV���*Zv��<�J�(yD>��iZ�4��W����=q[?pG֜Y�l=�j��=�¿o�}RhT�T����zX��Cj
6���Sυu��.��GΈ����kG+��W�
������7��y�+�#"\�=�Ս���1��t� ]�y�����"�Q�����{;w��NPX����i�I;�s-��W^�*���ʔ6��C��u�h]%Ü��|����S5&�o��Ý�����Y<����1	��c{�u��)���Zv�"���<��Y3�˲��pbA��<0Q<Z��5�
�NKLVpf�!���	�����-�8[5t��t<ҹ��JʭrZ��p�}f��6�e#�Vf��Y�6�s�KN�y;"��,'v�J�]6���y³�&�`uc���n7A��;�+pnv�&�>,sL�V׫ӳ��ij����=84C�/
9�|�R[ �Zv�v�v稼����c��%f�WU#b���C,P�j��ݘ.�@���5{��o9���Q�p���E_��x�GA���*���v�?X
O�����z����Qݾ�,!���i��#J��c�^sB�%�prGD�ZH�C��c3��|Ĭ���pC�z�-TC��9�HW��b����uqԋ{5{����Y�y8�.A��SSͽB���4�!����TBo"��7+mu�v�NR���\����nyv�roxc���o���k*��!�CKI��s��őӄ��6w�Jܚ��{W�j<v����c_l.��4�$+@��Q�
�5�-��__��gE�4�[�B��,�J5�+�j}����Ú��v�ʨ׆���O����Q/0���5���Uv�jq�b�E�@�˟9SA.n�]q�� ��7o���1͉�wa4l�K)Ӥm�C�H��2�㝤�))`"�W�5|�^_t�8ؘ���\�"��&8�0Y\	�q�]��1`y�4�:m=#�tI����kZ�23����i�/bq�>��G��O�+�M���#>z��]�84�G�W��~�Q5��x�y�j����tj�D�:q�;+�,d���n�����܌J�nr��:�1D�b�nsb�/�?Dקn({����֍�qߜ�Rd:�����PՍp�cb����ї{C�a��òIp��j�j�Q9QH�s ��f�iAT���0�0F��/	���o׊^��}S��科e4C��v��O��XǱg_�W/r$��ї��B�Fҩ�>On�<�&���"��"��;�WY�:�Yo;Ĵ�K�ֻ�*����9O/�k\�^�{��&��]���͒mZ8��D����p/tTMf#�����Z8�[ܹ^~�m�ڒs����M��;�����R�P5s̄s�з��M+�s[�3��T�K�&�V���\Y[<=��˩��O�"v|���hz6mcIR�T�(@]���{�)u=����~�I�
u����-��h��]͓ [Ť���O�SN̚rv{�i캘����Y)���[�d�s����9 �|3���,c���ۣ�}�^T̢T	J�h%>��]���=�r�İ����U��Y'��>��p0�T"��1xt:�sSk��.5�yX��\�x�.AM�v���I0i����k�'܆ȵ��W�WP�,�^�нP���r-K�߳<g�ơ7y��1���yW<����r�k�qz�{Y;��qy���i[�>��z8e[�:軬-٪n�Hu�>�]�s�[�z�f#o��}���>�2����'`=���غ��l��)��I��.�#�e^Y��*c����g4j��!×�����6mkMw_^ͻ9Q�fW�Z�v5�{au{�5g]�����^��j�s���A.l'M����]�{g*)_��r�(���JGu$p����qRw���/ѕ��5��lR��[i�|�����1�f�z|Y��7	���/����R�:�Z�ܖwr�s���i�0���Is��[I�ְ:=b�+B���kj����S�{V���=�fm2ӏ�eL8���y��������:T�KR�N>i�=�� ��ָ�y��ѓ-��\ǐf�d�wc�7 �	Ֆ�e�>�z���p�{������*��R������\=i4��o7w�#�X�X�;3�"��w��A6���.U;),�t]y��;���Lr�[�+���Bs�qÔ�Oyt��0b5$�oR��P��il�щa��=D{z�}��7��sz�y�2�S���������#�5ɉ��m�5��Q��i\3��@{��g)�+������=��+Wv��(�h;|��Zzy����Bq�	���H�v��Μ���[�e=��Y�j�{:M�����>A��vL;��k�n%; ��`�I��w���	�5tώ�e�'�~�Z��o�\Zp�zq���ǲ�钜���]�}�߶2���Gm���/f��Ϥ�u��_Ӽ��5����VflIߜU���!Hs���:-vD�Qo+�hۈ�Mz������S�N�H����εz��c6��YZ��G�i<�����6���������I��X��_?���Mot�wP̨�5B�]>I��S
�si����� �`�k�K�g�M�0R9 )�Ԝ:�	�jC�iM
�s}���頶��v�0�k�b���3B6,���i�}8�C�ë���J�i���Up^�\T���̆�T���@���n��yx�_V�;�ف�l���
ǜ����W"�Ѓ��c�bc����f���EJ�F�����{xD�����-ڡ�Y6�1k��3M��%K�Pz_ݦ�X�Z#0X�.��C^*��׹�CrV�.�R}N�K�� ��#vqH�U�s�]��:,�u3K�[���;j�[Bf�ƅqv�I��;'(Z���;z���Rh�8��C�R�qp�$��g+��!����	\l���s�X��N����>v��(�C����	|���}w/%>��pуȪ���w�̣ܦ��栖�h���	#K��fN�ui�S8j0��jp�;��Fa�>�&���*K�Z&���F��j��9ٓ�{\)��E�瘳莍ꈐ�3F�RE��[pn�[��x&�s�w6�]M\\(�A9(�=��Z))�h>9{O.e��{wŒ�T
�^��aK�Z�7+z�vA��_Y�hM�4��h�gH���s�d�eΦ�O���̮�����o��YbK��`&�n��<��Jxy2���GbB�����o����1���y�mğ�qY;MM�ӻ�*�3q�Ƶn��a���F&�y�h�ƺu�:�i�#v��{b���Z���U������b��Q�m�t}��k�{Y��v/�i`�ŵ���t�^��/�ho���dvL�ΐ�G�	u�[gNN�5g�R�ڡjs{���t�J�@V��pR�\3�[�vNo�M#�jGa�4��+�=�jmx�� �:%I�}Z�5��7Ƚ��gWM�:��n)]
x��z�F�o&����q
n�y�bɰ�wA��vŨ��,n^6�>�F`_�u���hᫎ^�},�39�(��;c3J�U'&��k���ebʩI��@�t����v����!Y\�����yq;ضDiU88��T����"��{�r��-�&8v(��*&%��w;G@0�&�d�GUሻ�,(��0B*0����oDy�լr�vS#l�`G��*���(6�����kr�|�Ĩ~��Lvm:�{5�A��3����F�ܥS��ܠt�߷��K�7V5YNl��n�'0���S�g��H���Է�uBp�`_L�[���i/�WRlaW�3)L�Ӗ��nv��h�p���A��e���SV`�/xĵեK����K{ѽٕ�	Y���Z�}ج�|�#[S/fP6��軬�wKi:5r*Ns���J*��X�M��f��j$B� �R�B�� ���(�*�R	@���"��PP ҂RSB�"�%(���% ��B%�2����o�sMZ#��j]P�nظ�"�K�ڢ�s�ٺgc#��������x� ���m�@���p��k'��-���q=Ǧg?���N5���v���AoZN�x�m�|Q{K������%����Kvd]�k�S<�ȗ��:ͽ�U~����z�:d%�Ǻ�o��:ֿek�y��K��ډ.X�|�7�\ط��55�aXQl����ԛ���w_o�܂�zw��m8J��Wፅ��(��5�~y�������)�7��S�B(��;z�8�Ϡ���e��PU-T�kx����K���P�����ǧ�%$��-���ق��ʧe&�K�N��8��4�(���wv�jJۚ#>�W�#\�mz�-�J����*�cRCqT6�Y�A5���j͕����%�v���[c)�U��wg�
'v�r=!�o3P\��0��g�Υ����J��O0;fۖe���X���̈#z�ef4��+~퓽�:�^��7�I��?3�W�{�Ԧ�����En�y��7�gf�m�VN�/ ��#�Ԃ#�6&���cw4M��s/b٬���ؽ�l�Ǵ�zVE=w0q9��՞��b�8Y<��)`�n�u�V0/���6ѓ�֮"��]��F�JS�^�	���JU��*j2S��Z��2��Ra������o��g����q�5ܝ>Ck�3P���>��!���f����p�������J�L�;����M�ھ嫝���M�↣
�tS�;��_66�]��Z쉎C�Z�t�{2�qk�OE����H2&�c�I ��j�v������j��f�X���bW۹�R��g�/��ŝ:�g٭ׯjک��}��N�L)�jy�>��R0���x���o�9��-pU7�BV�QՏ�x�7�[U�~��Q5��KLm]���{���[x5T�^U���o�ƹ�<�Q/�ǜZ�yUٮnr�4�D��x�(�߾�s��XOq{B�^��zDlN�hpܼ��9<q� �z˜���s�׵�>/(�;v]�~5aMŞ��B.B����r��Ʌ�~'��o�}s�,�y4��%���{>���@hQ^�z��-���D<��s2�o�*i����O���䴦�֨�:�,%U�M��;}���N��+L�7:�61�3[F��MK.�.�yu�oI�7=k��>�x�Z{�BhT0Zns��Q���ږJ=ՓJ��Ӝx�J��]�ٱ�6�xBWtzlV��ذ�N+l*�N��s{o�Yq�דOD��(t�0:�F�On�fc^<�R��49�q����Of��yp�������8��{HW	�H�؜�Z�_�������f#�^Z�Y}��s�w��V%u׻8��[mu�ͪ��k��>��y)��KE�\�<�u-�	4��w�7�m�-MOb-�.�a�N�]30�]P%(�pS騞]��❍]��Xޚ�[ˣ�'�ѯ6�;p�1J&}��Πu��E�IgEM�s\g�����f���5���P�T�$�5��k�n&5��煭���28�tOy_jSů|'.�k�/-�=�jOni��M��w9���5s���m�C�w�\�^��=�Q<��w=���w���'�{gs%@!�ّ d������ki�r�u�"����&�W�J����^��佞=SN�X��o����b�j�ܴ�mXR���Õ���r������K��Ҍu�.�vk�SJCN�:��Vt�t���԰3�u�qM..[[X�3��%7��N��͕�)���#�V��pl��V����P
e�]R�|�(����=u��uJ'�`�FК�I���M���}���eAw0>Ņ�f~���kռ!y�&$�q�8�|�0����eh�~���U��:�aMc{}�x���\�j14�Q�
G�Y���c�_B�;ke�����W�KR���0��N���<�}RR�G��b����}n��Ǎl������i�8�iҮ�!j��Pͨ���ꢔ��9��=�����Oy�7��2���KV�Nf�|����L����TN�K!]N��Ai������C��SSDt.x���õ�gK`P��邠��t7���^K��cq�2��{{<�e����.�s��/z!�8�(����Z#SV�̤v�.�fz�C�\F��~rҸg5�pSl�C�f��^M8D �ݦ�:��5;�.%��!����|�����x��n&!R<��;&y�]�>�:�G��"���T#V��Έ������w� �#ir.��cbb��lOP.�����g����L��j�Ք�T�f�:pA�U�^=���P�����]V�*p 6e���Ծ��ԕ�KC@��ڶ�%\Y�z���O�],��)9{���{UǨ�M ����M�P���|֚��N� ��)s
�N��2�
�^��+d~%!~}n�#p���9��^jڅ��j��ӆH�^mLʋ�S��u��^�F�
���D�����ꈗ�:/$�O�]��+�v��c�u#���\����r�z���o*�ẍc��:��
��}\ˏޮ��m�펉�ZN��Q�L��9]x9��;�fTw���������8�^�GIz3�GV4�L�`�{Нf߶�m��B�k۵&�����^.j��N 7�s�%�끊/�g�sb�7��]�j�H"jq���"S!�b��G��<Uρ�u���P��k�q��܈����7Y��*�����}��^�2�L�U;,�+R�P1���@���V$�����OS��ރ{��rB�ԢvRy�T�v����q�,랓��.j������O5[�,����NN��P@/����Mm���g��rJ�ס���u)�mC�^�j�x�J����]�6�f���:�(*����>�5&(��̮L�a�w-���,�j�!N1E��<����8�o���:9)��S^h�w��9�|⼑U���P�-�o���5qs]��{�.m��+�O���ı����m�e-�C��:��՜�w�yX-�ּ�g�p�M���/�k�e��c�{��3����6G*��yY�\t��^��B�{5:��#��o��Ҷ_l�.��8�Fz;,�P���そT��Xt�/dV(E���7=��-m8��Ô�+&L&T����u�l7�Tg�"f"p�Ty�c�R��wRv��U]��i�]�{�k��q��,���"}�v}f-���>�;^0�����jj�&��׵��N�k�+�����^��Y�9b�'x(c3/|ԓ��s=��n�j������_/>����(�JJ��c��Ӟ��闫�CC1�[��gj����V�o���4��ᶬ�����Մp.c���U�ya'�Ʉ(��@ �Y����._u �z˸U�a�R��V��X"��I"�o��S��o;��١ΈDnAӉq� hڶ&�WbaV�	 � յ�x�9��=b=uu����PgqZ�urvp�PdYu�7E�����M����w�D���lQع�:кͧ3ju㦓�u����z��?v��ZV�σ���Aި�tkiCV5�#��x��]���M��ǜ��O9�|�x��������y�KW�����fZ��V�^]<Z�2�k����<��i��Onl�v��@nA^��Lۻ��ʤm�EvS����+�:T�k˛ۇ���c���{f���K3�d8 �q��3�.����Zhjj�P���9O/�k��-�8$�25~}��!�ٝ�ߧ�~��R\�����g�Υ�����|�����a���/����)~�amB�f
}�J	h�Z������]=d�v9f�Wv8�9�d�)7�����%+_	盎4�\Vh�8�w;�ϐ���ݨ��q�¸�)@9k�����u���^V!�o�
�4sT��f�Z �B�Ys6�t5���[h��p=����3b�Wy^�_��s�!��/;w���g1��┏,��m��T0�L�;q�B(������.�kt0�=wQ��9S��_sb�ٳ�75���I���K�A�d�g�W*��Im.Yڙu�T�$�5�^5�^"ܵ����w<���b����:��-f\�=��[K��$�j-8e{�9?v�~�����Io�m�L��h�ohf"��yk��{^��m��#ζ2]CXʆNL��t�_Y�
�au���2E����T	X2�ڝE�s�wL�����Z�߈I1����߷����y܏�TM�A����/��7Wb|��;���
���u��!5�ջn�9��Z�vPU0�>��:
p���]ڕe�p'!�b���ؤ��n��c{�-��g_�[�1����/C�J#���ǻ��Yg=�Е�t� cb�`o-����>�[b33�ϧ.Y�w4�N+@S��ʽ;<]�]�^T�X��ކ�އ�,��D�״e�<�y^��i��;��W�#�$����:k7���^3�^�O�YÝ%����ޝ��s�� �|���k�Ԛ���W�"��y��F׬���Lah2�<jU8�5��;e���*��$�A�Xz�ƞ`�OJ�h��T�7o�TI�Ҡx-6eԩ��T�{��d��;D�+��}�c6qc��N��i��qB�Y�)JU�Oy��$�z���vc�t�u�̮�NL��i�]��Z�-�t'��r���{�b ���j9�{TV�v��\���8ӎ��u�i\3���)�r���"T	H�U����Xު÷�����MN��n��ڎ|��^W�n&#�͵r�Nv������E8�:���Mzmv��ro�}	����q�ʚ�����k{����L�Ik,ym\8"�5��j�V�.x�S2�f-֐�� W��0d�:�aR���oZ7U���:|-m/s��Y�y��řɅ������Z�ꮸ�N�yG)���Xn�P�����b�ޑ�	��c����~�|�'�/o��k!��e��s�u�fQN'2���ㅞt�v�;ը�K�=QR~�QX�D�A���	�m���[���V��-�e /g,��Q��rl�h�o{l>��G���秌^�泊v�Y*�/sM|Jv0��pD����a�J�fG;���}	�Z�1��G�l�I�Q[
]�������jk� &�|V�)�e��23�s+��¯�H�H����9V��9�X\>�Q�ؓ7+��I���� ��i�O:\Q�x�\��z�O�\���][*CV��Y��);h����pr\&G�25g��.�������QM�X�`�{k�<�y�c�)�W+��$�D��V�����ϖ�vR|�xTKᫌ�S�y�W)���MkOm�ko�ި���Dl�W����%nz 	�U%c�ް��.�v���}<��_�ֻ#\g<f��T(!�������^gsѾ�p`G_h���Ȅs�k�󖕇����1�9�����ҧs�����s����^�\��^[�k�J�|���@�����	rzډ_�&�~��E��*AZ��쭎��!��tTƜ�9z�l[�:��.�q����(���6bN�u�[�S|����8�E�s8^���[��+�3&�t��wT��Wi�"�&:�� �\n7hpl̽��Y�7�����$Gz܄�y�vY����v!�v�E:��9хfTu�^6�^�V9ŉ�mE��x3�)0�B�e]Ӻ���&N�kȻ�%�ʇ���	�­�'�9���5� �ģ�0M2����S�(�ه�lK�6�8(Cz�t�}Y#u,k�u���j��Z�ò3ZS�E悤��N��Sn�Z�r�S�,�Љ�F��WS�Wn��!��A���;{��L�@�twU�)č��V�EFP?X�xJf���}��#n�$y+|���d�A{o{�<��Ҋ��;�R��qkJ��)i��{Yo\k5s�j��KARt�b�ع�Z�pf/J>g+� y+���l'Y�퀮7�;���3C-��c��ZKZ�a�R���fƻM�ڠ��nQ��E�y�Y�mn���$��yB���]brJ<���::��<{c�R��:QEp4��&��qU����b:?A�9�^@��Cӌͷ����f�W�K6�����eV���VZ����N��|�=��@,��c/���eb��b�D�(%�MWl�x^�λk\�@�i�VN�F�9�NXo3�V�Vh�]�� Ad5i髍b��_N#f��\{v"����&�B-b����VӒ鋏��\���wlz�,h��^�k�P[hf��k�gM���{C(�J�T�n�)��,�hW^�zyM��g#�R۲ͣOm�Qٹ����3;z�2�O;�j��*�j��p��V�k�;5�.��J/U��]b�6�(��}�OA���Ȁ���-Wծ8���
����^�h��:��@���t���v�{�J���ہA�,1a����b�]�).�f�գ�vh�CU�c�5#�I�� ���iJY��"�AR��mDA���BM�Z$��p6�V�Kâ��jW^�MwG2�om$z�(i���2�6t�����l�[}��L�#]����4)DN�����orv��&8U��gk�l���(i�����Po�S�
��ߞ󺫼:3��wZ�[�N|����ȍ\(d���6ڨ�\���$s�$�-�,FJ��K�5�����sj��l�CD�U��X����3�>
A��Bޤ-�]͒���6�Ǐ_F�Ɍ�\�xS4:ZDf J��'E}u�h�,PZa��5�����X�ӾO��t��d�����I1dͽY `���Q[6�q�R��M���8l�방M�ʹ'h�&4E77��ӬT�3Nn�����;8ÙF� ��ܸ�:�+ͮ��9LQ�6�,��Bc�y��~��!=��G��nL��I�ӥ=����xܗWG/*�	K�f;Uuܡ��Ec������@�A�:����S|GI��9����e�cR�q�wM>�-s�G\;l5S�I����x���[wB�DQ'���캢��
iiT)T(E�B�ii2(��rJ2E2Q(���#$h�)�i(hh���
�JT��@2W������8ҹ7j*U�dyh���:7����{cz�2P<��p�eb�kM;��)�:��\�z��ɶ�c�Ӏ�2�a]�)���;MTע�`�n5߂��DLj>�A�'���W�jSo�u��
]*m�w*�y˫�N��k�5~9Խ������Ug֗��1s3�M�wW�+0�ћ��^ջ�r���k<��e�b��ɢr]�O�N8\3*���m�z�}�&+4K�y�j$U\�uH��k�/�uY���nժ��m�b�Nʳ޸��Q�>�N)���y@l�Ӟxk�8�Ƿ�oun����{��K|˪����ǭ{�cGe	����)��%��E4պ��kUE�[.�|��(�SQ<���%�_\�������lS��\&�[��hjƈ{����M5�,�~�.����{�9�G���B�SP�������SO8�Y�g\��[�2B�i3KK����gwjT:{5Sˆ��ȇ�'���ov�C�&<�Z��	I�I/r���ὣ��%�l4�M�˘�r=V��J���դn`�#c���sGKO�t1%	%������fi�b�F�c��f=�K�6�u�/�]4^����9[�Wl�&hN�/oz:��hYꏛ�pu�ϙ��ַ��Y��ݕt�y�^KF���Z�j��"v%��.l���6v9�]��~��î�O%01-5s�G9�Nĝ��fJ�j�sj9�V�kx�M�k�P��J�y���ocMw��N�-���i���l5��o���;��%J�l��E.=�u��y��Q�Ǽ�����ڱys����$�4ۍhTk�2�qۮ�Q��Z���V�6�ΞZRZ�mjN��8f�pw�&/dH�1q��8�����{�Op�ohfuz^ezyk��{Q{X�������Z}��9�L�cP��ҜF�;J�}��b"���ϊ��<��͛�n�|���/[�>3�2e�Z��Qϫ9�Z��.�}��nsj�{I�*�jSQO��y�"�.'ݏ��)��u��[�{6��s�V;����Vf��-�$T��ܜY��oT}]���0�Ĵ�G�$!5�W����=�0r(��D�,
�6��(o(�C��wǎ�c3�su����ԛ/+P��Ns�=X����T���%}�u�R	��մ �9�T��A%��:0Q�����Rɵ��mo.d���%�V1¬-܏޹����kH��;���^H�n�Gx0����=|����[Q;(�K��V1�P�7���y�Ђ�)�eĺ�7�����.=���g0�c�9]a��Cy���0�-S�,����m��x�ۃ[�(t��%A�|�Ӳ��W���,��y\�D�;;���wPޝq������Z�ꔫLw��ѩ)7&RՌ��3��Z7���M9}֎>��q�^x�W��>D)�wIc �z�a�����a���g9ov�)i\3��x=�^m�e�D,��޹y:t��Ff��j�����q<��B-��Ϛ�2�;���@+(B����2�#���l���6���^ͬ1�n{��qap�a����:ڡ��\�썶Į�'��m@v��9�\f��\�����)�{Բm�g�u[/{`���ư�tlʶ6��M1ymϗ��P[���'�`n�o:6F�x�(Ď�2q�v�Scb>"����W��_k�s��%t�i�Z�TkB���eu<��4eHl�B�t��-k{�K�����M��"����a�������k�#u���7�Z�}R�*qk��dl�n9�ܻQ=\�SZ8]X�u׉�4�W�ʯj�u�L]�O��Y���fI]E��¼8n��~{�g��yQR���Ƶ����F^O;7�]�R�*`$����v�GRw��m`~�jS��w
g�/__������x�헻�a��������Ne�GW���w���͋t�-��9�
���W�R�{��[}z�w״s"+���U�Q�P�1��w^;�*��� |[֜W&��ވ5��g%���ʧe��PT���ͳ�C�zn�ݫIc�L&��ho-�}r��7�P(w 4(����s��%Ff�cŀm��H����>Om�kq�΋|�J[�C�;ϛ�1������Z�?L���)��츇/��ֻ"5�G^�u^]�S]�8���[�H��~R����Ю.��ա�O*e��պ��r���T5��t�fZ��"/R;z�<F�jNP�j�qa��y��mV7�[���U��e�7w���?�+�ܸ������qn����c�i�������g>���2j���l��:��˳�REf�?N��Qy�rҰ�^�=�-ћ9�2�lb����mN��C�w��	�Q:��#�k�UNzB7�����_4�ý�zw|�b��بv��z������.ڸ�NA�٥S���ϣ�'�m�p�c�
�}
Q3��)��+rT�0n����C ]��I��N���~>q��MZL�mƻ�3����6`_n��޿j�X�z׋PqQ�b]��MZ�V+�I֭p��A��V�5��Sx�ԽQǞh����u�����ѷ�����^<N9���xK1o'n�(�R4���Pki�uF`j.�ͽ��^{�D�c�v�5��r,�=޺��y�������w7TAd���C�zs��ʳ޾�Q�Uz�jK��g.��~��V�}�&i��Gn��h�>���/hb�?�e��s-�ʊ
=�@Wt�I�"�#�Ef*�CU#�3'&�i�涮i����w]CH=;ᗼ��cpi-+f�M*a̳��UαaծU�n*�sǕ�Ү����(/�-NT�V>�q��5�����9-y��ݬ���3�	�G{�No@՝Ef�䩷�¡.or�j��m�L^�ʤ��yp���n'z�,+�ߥN��R�J��)�o/К}n��5��xգ���<�y��s��۽��P��-Őx�Z�͔�j7��5���&��sB�c�y��9����]:i��1j��G��1�u�Aӧ�NS�kZ�\��EF,�Ib�qsõ�gK`PS�}%y-y�B�c�>�m�FIڋx/$��\�jѕÔ]Qu����S�k���W�Znv�׽��k%y�mswޯOHj��o�	��t̢W��^(n,\#c��읱���RWvdw&��T5��6�8v��%J�6���5�7�f;xTn��w��w%55k����W0�ٖ�`�6�Z�
CX�s�˸�p���u<�#hk���/�."q=��Z�n/�����⟍j�Y7-��[;Wz�yN�q�"bъ���0A�O�n:�2�6�s�\��]����ۗ��A���K���(��������aU�re��n�|(v���	����Г�zTQ܄j_3��̒qsm���m�"�c~W��ۮ�O�}ҵѭ;���b�����1g}p���ne7�v�:�����@�BT������a�_4�\�2��͇s1���!�/�f-���%`�C6�m����/��o�)s�T������W\.�����4n��̨.�ؾ�LTKoT
�:��ts{��U�U�q�D���2��Z�5��{n�ds�%���2z�}x��+��
��wb�j1��-�K��M�®�U�z):�TQ���'��q}�.H�c�U~UzvY��P���J�1��7|�|�( ���t��n���^w�/ʽ�y������kT.��o5W�{�N��r�|�.�aM���������w�P��I^|�vR�P�����ğ(27��n{���Y��bzמq����>�*K�W�Ǘ�k+���J�Z���:}4��Z8�S��x�TC�f
{�Ѫ�w�)�F�z�vS��ƍ�+܍�gUe<3��q^*E���p���]Y����t�7�j_���$Mz0�iA�7;�޲萵j�&-r�<P[��)˝��]�.���i-��w��x��M�g/{�Ҧ��(uZ������+�ܝ����~��=��#��%�i\3���)�r��=y�Tp�yVwwTu+�\9J�}5<��D"�=�������s6�w;r�8Q7�%(��^��g�@�Ûh����ڛ����P�Q�bO*�#F�E݋ւ��-��zFBtD�r ���-�Ȝ�q�#��6�v�%�=f��qˍ/56j-8f�q����xD�1�-m�����;�j��
�Y}��Z�S���Y��u�18f��W���f�Ѩt�OqUdǢ�gZ_���V.����nW;*^�'�>��y<�ܗ��	���"%oOk�k�d6s�qڢb��3͌����ܮ.�+�R`W_r	w8�g��]�@|�&��:����}���e�]	�&���7k�Ó��I��=H�;=~k�UXSq{F�-�!���3�*v�dVJܺ]��~@��Z�2���X*wv��Y��)��Ө"��I�hX��_&��:9E�ā�(bX�'Vq�4�V�z�P\a�OE�,-z��n�d���͓W]�r�m7h�(QK4�QС���s,ċ��8�4����AKGqq���X馭�>�[=�rP�<��^��f�u��ݘ��쥋\�\[�v5<�=���z%�����(t�B�m)R�����M��=2�K��e>a�s9�|�ߟ��=�|��%B���1G�I���i�E�OP�*�CF��1V;t�j!��5�vF�Ψx�u�`�{Mt�J+{�;9�70`y��7���9�_oD9iXy�p(�0:�yUpp��jB��C�9JY�"����P~Y�b�˪�;᧰�U{�����^jJsr����y٘E��*����j'�mS��33�-�zl�T�1�oP�3M���v�L���	��G��]O`f��p7��}�𥉉����V�mB��U5�I�ی|��f�KB�N��U���^��:Dqz�Z�Y�9��ugB�ē���Ps[�T)����cv�{s؍Z����Q�>�a�Ʀ�~V���jܾ̬x!K��
/J�6U]�P\T��^�����|�y5ZL�vhd����c�w���{GÂx"]�t$6G`��"�ib�_a�6�ڃb
�v�R�q��uH�B�DAZL�rݼ:NjF��͑70X"VM��ҵY��)��3yy<�m�W�n㜽�N9�-��Bn	P����vyj`��<�m�����W�>��|Z��q�����N߳��Ԥ8���sMM���ۣ\������T��@��7MC���P�W�����z�zY��99:e���_�hC�XM{���=~%���+-3�z�����T(���\�����9��6��7�m��X�"����4_]��p:�,��AU�ұ���<妟9O;Ƶ���"�Z۩�֏>H�H%�r����+�*�J��s{o�Y~�ro��꼢kp:9T���W�O9����EG��d�}�{�ڼS�ɛHCj���Ub	J��k�uygE-��y�Q^	h���b9�S��):���L���B[/�-u���<�hx�k�e������py8�9'�n�YڹoJ�β�Sq�0�0��"��q�Zo��hSyV`�|��hK5��V�zf(Kn:D��8��}�g��.��c����G���hoh�W%b��F��8Z+��v�8:�E3���B���t�q�]���=
��!|hC�3w.��kofƵ��jhՐ�u:�.�Kz�M��fL�Bjw7���W��w4+���sNH�ԍ�v��CR�@c6��7ov����}Y������)��e��ߴg+�ԢQ�)rb�!K!/:���Rՙ#���tH����B�-���L��ᗕ�6��eS�����W���er�:컻���r���%A���#�.��iԵw���gQ	���R�f��»�Tފ��
�����ٝ|#^s��v��=$�:�WXٍ���-R��i����Mڽ��4��F���k�XF���Y�ֲ����S��b�Nt}A��ҧ,G؆�cU�F�Ҫ����I�ZѼ^�A�ռQ�&��'"ie�WZ�EԲ�b@-u��-�Q�Q�݋n^;�f��YUf�1SS�%�(� ia�+�k���lЧw�PC(Ш�G�������V+}X8�IVRVs[�V�es#�ji�)qc�:���a*�\I�gs�
<��J:�9Y^�zh�:4�b$�H�5�\Y�%`�5�+�˧I����tE�9����{ƭu-�\�C���cy@�Vr�L�E��/��t�tW�JhѸ7B!VK4����j=��>�>P
�S4e�^^|e[�rԣm�Wlgt8�}M��T.@�wLYR5��d�|�LP&�T�k�
��S����4�Ӳ�
��5]�V�)�E���v����*�6�
��^��a�ӳ�b�Y�2>�^U�ڌ���V��k2l{��_#���f����ZӅ�L]J�B�]M\[)���o�}��X���V��2*RM)�'b�y���.���v<ɵ�q�
{���[w���`��[�L��i}�K�kbY��[p�vN�y�o��6(T�OWT[����#vӁ��v������1��Zێkݒ���[�	����E���L�QØ�� �2F&�j����Ub��k��34j�EG2�k9ʲ��؎Q�΢^��
�-�2�\	�j�5wxcnq멇EnP����X�,��v$)fN�>=Z`����n�A��<0�i륒��8Tp�^�/ul����o��p�{:p���-��|2�H��?=˥���4n8���&p��fgɹx��⃮촷��`�z �����+�Di��!�\���ɔ�T��q�������F��7�Νj*�d�V��vU��65��{a�,�-�Uk�5�}�9��:�0�9z@�h�Z��7�U���5�V���15�}��"�iqp��zgt) ~����}_p������
��@r����)(�(JJ(����������J����Ȥ)��j� (�*�,�bZV�B��
�)���B�%(
���ZZ�Jɟ�v����v���a:�Xg��˺��Z;��RUclN�QK�k��:iX봴�{%�|7��L��jc�b����M�_��I���o�	��t̢AJ�dfl�W_eU�� �����{��:{�y�m�v0�+�ˇlY�]+(�����{���-�w'���m���rڅ�:����L�n5��Ȩ�v��Y��a�{5�í�ۣ~��.�r�}�:yjS�{�OfM�$V*q\�&j�L;�/���%�Q�ϗ�ъ�k=ݿc�ϩ�"�-�~�{�O
��+�1���e��pʷ�v�κ5o�Ҟ[}�zGd6sPe���3���I��Obܞ_q>v�oE]0?��OpY������Ë42��W-��������^��%6C�|��Gf]Ӽ+�n�-�M.�G�(�u��j�.'z���c�Q��P�6.7�
�w���,l~�=�}:z�Y���g�P:��ruBV5Ҹ�x�P�)ENQ���СR�s�E=k1W+��*�]t���u�]�u��Å]Kl M�<[#b���eI��#���x.(�΅���:��$ȝZ�)��L$�t伓.u,+��f�2��v��R-��թ{�6�VMn�d�ف�pl8�A�1��͖��u��T&Gܩ�c��j���9�P�lȢ�ٕyt��go$*ū����%o�C��i���^��.�	C��	!�Nw���S�ٯ��+z�W+�4���BN��ֽ;�8}Ǻ��>�#�`��W�&�_qy8֭Hpk�[Y�_OC�܅�΄�:��9^r��;��z�N��S�����w�; �t��YO�R�zC^�;���؆��D�`��UbW��n�|�]�wx4<�j'�=�[�=�Ϛa�p3�e�4��0{�'呥{�L�,@��:rV���]�qܝC�O���0ً7��-szk�q�¸���6|
��
�˜�ܕt��O[��F���J��s�i����8e7���ׄs�������,��K$��m�zTۉ������r��9:�NP�T5�Z��j�9��dY-`�Wp1m-P1���RW*�"���)��z�Q����-CO{����
(�"�i7�Y�]����+uZ{��Ն��6(+ �,�)�m<+n��uvw_�>ݧ��u���1	U��ζΧ"��G*B7$>���Qqɭz�&�a|���W)�]�Ƅ�"�zuy�]�y*�^�K*�z����p��';E�:��1�9�y���QX��u����k.m���4k��Ԙ���L������zs(��:���Q�xA�a��U��f���|W_�k�55�~�eGml�
���;��	�yr_��
�0���<f1h}���SM\:��w;l�4s�@<�Ƨ�UnN뇸��}�GQ~��-�ݷ�����i�ؑ����c�Kf9VB�w�ʶyCOKo<����N��'��X��ڷ�l�I�����Z�R�*r�*��&��T�Ƥ�1V;�O��׾����q��v烻��7Y�3a��6ԵB���wI�-7��G:�k�r�֦@���]Fe����`T��'U8���>��IJ������AӴt7�ޮSད�<͚���V��*�8>x�\�M�G
�OǤ�T��;֨5Ol�9(��Q��l�'���\�KT=�U�;��3M�@�1��-��i�c���1F�d�p�#��9�vK}�rT����	�qϚ}ڻ/�v���h9)rƲ{&MZԔw�ZW��B�{���{bJVhE�"^wnok��V�g�\��s7�t�:��mr�j!����]�+�Q7�l���QV6Z�m0ok5,X�gMM�ڸ�[K�;��MZLm�񫙋�-D�0x{���	Kw��4�}P���ʜz��um.�W�m�p�(:�۽��ED��#1}A4,�U�Sv��1��M��v��)�V�?d��[s�=�xy����;��%-�N�2�&r[y�5V�e�������h9�`7��wm���fu���q�jڬۍ��vn�����Q78���^z��r7���o$��/�t�-�Ty��ݱE�j��?�*��9E�ksU�Ų��ܣ[N��lT%��DSM\:��w״s�{�	��gv�q�-X��/��=���F������Q��a�p�|�<�#���
i��ظQ���ݳ�Yap`X��8�J��a�Hu"��KZjn�-�V�b�o-;��d-8Y�8+Z���ա�ٸX\���.̳���7*Ժ"��&��ȴ�OGDԇ���Wtm��V.��:{�LlB�l�� �fi��-V�T�V�4/nA:vz�Y�������j���¯*U4���y�k6_A����ۉ�YO$�����g{���O�"@�d���y��W�s4���1�<t��f�Y|�.����y�Χ�r��^�y��Z*�Y4ŕU<9�Ô��Mc�ͬ~Ժj��Gny���e�B�w���U�'%�4��S��,V�I�C9�xm$Ҷs[��7��ȯ;e �ٻlmob�qD�rJwV0�-�<�3`rox_=r�|��;��Z��Y�Ƨ=�֡p�����k,)�h���ٵ�5������z$���7G6f���Z��%��G�@k#"��-e���D}ƫ:yiJ-�zye�S,y
����������s����:b���>'~��;F
�\5�X��6�yM����ql룲'/��|�bukp{0�۸)d���ʴ�s� �5z��v�fౢG��=�Ƅ}��nf�\�����c����xh�l��i*<����;F��cB��V)˫�����u[��g
T�ݕ�Y���Th����֭su��y4���zA�\�c�dt�w"���r��/%�˅��^�;�2�-�B�9_^LsF�:.��5Ϡr���~y̴�.���nr1��;>S)�����=���Qy�=��4[�m�.ޗݣE[SqMDJ���O�6������5P-��z��B{QQﷴ�q[�a`�xoؔ%c]+����mZo�t����^m��5n���v٘�O�8�;,���ɩ����V<G��-��qEm�z�z'6$o{�(>zN_�TH�iGpH��'���6����*��gZyp�kn��睔�(����-�髫QӱІ
�qθƔ?Ą�_�k§�^r���ۉ�uC�r�ʨC8�m��~.X�Uy��<�]r�H�����]�}��w��γے�Eh�᫽�.�6��C�h�n'W=�T�ѕ���7�I����FƑ� �^׭�j�v�l-�ʬ0�g�(_q�vm�Ǖ�u;��$m|�>J���/�ٿ]
*o6�G̒�������R�8H��{P�<�)Kf�n�r�� ���N�GM0t`��l��B�p���r:�SU�ɗ�\��tva-ۇ���e��CYS`� [a�����o��Z��"���"�$���Ϙ�Id��&7�+�� o�μ�[��e��#��o9zf�;��E��f��6��Sޥ�Uݥ���ܾ51>��X��"�NM��.��GI{���.{Y��f����������Yc�r�$�z�̫'ۊv��ѮS������E�W5�}Gd���z2p��Ć@�V�	j��/C��j�y�Y�����k��z��S�i�/���Ǫޒ㲱9�a��4��[���e��+X��t.Q�##F-w�]�������w�^ls��[����e��mU�c���"���u�kM?S/��]�nE4Ӟ͇[9]���[�B���M��$���B=�xF�S�ݪWn��7v�}r��7�#�����-������X�Cv�wWZ.^m[��S�݇�.�;BwHp_L������NK���,U�2R���Ǜ�r$�"�����EG�[u�ɳ�p����c��ˍ	����'!v�/&JY���FK6WwT�M��j�C\�1��V���Ot�ْ�R�m�z��7jvS��*�R����W���O��3˶*����U��˴�.T>�ApGs1�.�T��٧)嵭v`�}�ߋ�o���蛓�9T�Wm�\dʽ�����+_Z~��sڋ�:lz�r��t�;�'z����s��'�)�9NGDg�����&Z�"�.���*���"��yU[��lv��#5��<Y�zz6�"�W�$ND�R�4|�a��^�m�K��{���=�"��\�|�bFP}�Ѡ�zK6Zq���$r�JB��-S[p�VNj�﷥%�㡚zyv��{/n�����:���(ws��e����p�W$�-�y1�}���%����-�!u�?,��W�����_����C]�����*/�6�ߢ�L|�����{�W��4Xk&F���P.a��^�B\�Ƅ��<�OC���&��a���l\ɠ��g��o5Gc�P��v�']ʋ����O�F� ���i��eo�х��U?�jl��=�]Fqa��H��I�W(5�pHO�tU�Yv}�/'+�3k���6���ر�-���4���윃���fѹC��]�����9;��v��p弟c�N��L�7����}vuty�=����I?4���|��H�T�$cV����|}A.��}��r�����4V���Ʊx�������_���L�e���Y���,�Yƣ���������'��$RŹךo'|�4��=.�Ū(��7��:pk�u�O3�:��e�ޑ�q�=�ڻsㆋ�f<�k�ш�FP���WU}'��g����o��"�×��y��S�P{��>�Jg�`����T�$땦�I����94��s�y��~k�C�[�s��h{r��y�Gz�?��!��ᰩ�9I�#DC��Ý��Y�U�,,�ؠ�wǦ�n��wo�].�
E��z>�#�~�21̰�6L��5%0��|�����^����~��OКr�t�6����F�9Q�5<T�Px���w1��wg�髵x�K�>�MԸ5>.=��{M͑��븋��e>>-g�mȼ�eD���ԾzVgK��1_r$�_DL��Ez�W3Ћ8����i����,�7���2F�9��R����5}��9�q*��P��<a����W1�)�_л̺՘���N�ڵ,�`]��T͐rD������S�9u��}(�l��}M�F����	W�;
�ֺ�ﮥ���Q����Sr�d��l����� �����X��g�U��{[��Hޱ�D��rhM��űݎLt>{T����9�>߅,�C��Ŀ5����`��\�JY=P>4~���}[�=[+�מ���Ú��g/u���`�K�fy�07:jM�Qs���z�j+�A���� �v �����{0Nu�S���ǝ8�MaoWa�y^�����s���[ː�Ԩ�4MH��Y�����<B�z��C75��O֒H㱿z+�B����i���򶃾�/�X�Y�o��/W���X1�~#f���/��R�8��6xl�RrN�4��o���>	�?��w����#2�w�<�v���f��Uw�����?w+M3���P��ñBq�a�g�!��������m}I����o]kɝ��N]�n34��?T�fh!^�VhQd��P�0q
�y�F��LGu��U�A��q��J��j=;���o8�x�a��}:��S�?n\��'�>2�`⅑]5��{Z4�b���b����/��v��;�7���x�/���C�K���x+�l�^R�&I`w��1�he�@��;T��I��5�ȣ���}�3-�Ir�H�2��}I�!m7av�泡<��Un���O���D��5V�e=ѼU�,�8�oq[P���G��u!u4�)�g8�j^�Ȁ@c�q0OW(k9.٨�T������ǭn]�qˬu����̾�E�&݃X��c�;6���`ӹ�>����E#�H�k���ȴ�Cx�@x���{gh8�����^��c�Y|X�p8q���4�^�	��g9ּ�.Mwk7B�9�&�Ur"c�i�Nn���Dk��T��bT�s�L��V���i��ʓv��͹%4���M���]D�ғngU:�Zm�2�Ы&mA��0;�2�bʎfS���@&���oI� �g>�&D){�� ����M��rL�u�S�]�e�@�L�����u�(��w�wwD��f��ZtMf�p٫S��5.��ͧ�;�o����7���&�m�(�T�K��9��p��.⫂e9q�z[�:��(�38�ᩀ2�$�V�j�sT����2Lڍao:��0�s�A3�vލm����S<0YXu��[8X�E:g1vR�4��k�{�>�|�h2եi���92WR���D;/���L���3Z3��'o]�#���B���;�XM�;7�9T�=%u��ۙCv��c���͝�<1qդVB��#�+��Z7�*��K+��g��z�/i���
��:����u)��f
99�����Xp�ڱ3y�$D�en�hP��k/�m+q'��r_(x]����v��G�$O����_=s�2ƭb���EV�IDoUŅ�2 >"u��y�4rk>3�(��k;���8�h�W"@YT@�M��r� ]��t�#c�KS_.T�7$�f����|���I6i����3�̴�Ho���mU�qj:PZ1�]�G@6X}�:# ;vk7��vI ��;��Q<�zX��.��e�dѻI4��ߕc��щ��M �6a��[�5v �稑�;imK0a�q`gd9���ggN��ޓ�RXg[΁֤��$�a���*-)V4"�J�B�V`D!Q�q�/8��oBs[�+}�7:�ō��6!w�3l �,2^�a�S0a�I��\���A��q�u��Xu���YP_Z��īa��X���Z�T-�el�J<�7��8YioYׁ[+K���8��7]����u(�q��!�ķ���&��
�0w�f�~�"�AW�XӱOH�\�ک�*��%�Q	��`*�;�vW�!u���tf*]�����wV�f0�Q&c5.=�j�]��\C�{d���K�I��ۉi��X�pv�"�hh<��+��ޑd�x��*p\t�߲���� k >�Ra���v�;|���F�Z;S��V꾠D�4e��)%-]�d�Hn-��LfU�M�;V+>�W�:�L�A�
h
F�(*���0�i������)��
��*�JJ�b& ihh���iR$���)�(��
���B��)�)J
,��!��(hJ�F��h���)i�����2\��)�iZR�
)H��(b�(�J�����"����h&ZY��
�{.Q���luqO)9ln��4b�k�E�n�8:�S�=�	���v�VY2r�a]ǦS�n��s�55�]���{���E������~�uԦh:r>�e�,�x�~����W�j�C{gc�Z�N;���)�|:t���(g�]k9��B������[�Ú�����M��
��9c�s���x�cԏ���n1A�F#���y����Zc����ί�}Y�:!��:�:)��s�ۯ4��HV_K���<in��11+��7]-�Y�u�dh[o�ʫ�,��Ǒ�[~��~~���놽Kf�=����g���Y�"��~�q�����������|��Ω}�ce�z$wbh���pXi�G��7=2`��}
Z�|Z��|�����rZ������w-]��{x�k�`7�Rj�8h�71�7U�>�aɗ�����S���g�;������E֮����M���y�i���h���U�4�$}=��3V�k;3��V�'\ZP2p;���Щ�������wN���s�{���ء�Z]~��.|�>����Thx�}� ���A�������WDDמӉ�r�2�LX�W�����f�9���k�k哰�#f���~�Q}��'/����KȤ{��ra��l�6�>�t%½f�P�|�_��esT�j���o']�R�.�r���#VyJ�,���E�t�Pj�.���aj�%����؋5ԱSV�"��3g��G���,�t�^�&��6�@M��������w*�Xo��}r�U^��Nv�C�{֢���Ѱ�C���8&{���׉��/��.��]��H�T��}��Αs���8��tɿ5<����J�~�ЗNI�uȓ����,˧�m�ffL�~�b�Z��Ⅻw:j:��\P~E�f�k���K�`��׮r�0fMoq���,�9 ��? �X�WR��B��fݺ�W����!�1q�H���w�:��~��M�z��Lv�
�#��tΘ��t@�֔_�w+��R9u�1Nyע<�L��?]<�[�nMȞJ�Y�YϽ�iOf��P��F�8�*�>1�u��8�������`ﰆ��uU33|��f��<�VŎ^��{��a4��G�@��'�?��B�]�� �7�����b�{�{��<�{�B���bFV��4�7�k��k��dE|�T�9"r'��է(�́��j:�~X� �Ί�)Sg"���k�2����Y��N1�t�D�S�(9'ǉ7���m�=6�oP-V����Z�s46���΋�L����d	��s{�4�lڽ�Q�g;���d{b��Tux����}��7~R�%���Ġ�R���;}ܔ�ÿ�+���z��^	[q#�u��ff<Il�_s��jKP�fK8jc��;K��g/��~)V1�a��-��kuw���!�{U$Ww:(�i����(�@���3V�+����w������:O�-�-�$,������3Vd�eCWzo�0�s6�J�EEៀ5W���߆���~z��b�ڑ��V�\��>����4'W��et8�f�(�׀�<ks�Y����fL�sP�p&�atT_��T]yq>�#Y��܎V�����"~E��7y��u��c��j����xs������=S��i�5tW�.��φ��<�]W����{V��s>5�H�9㲠R֮ �Q2�G\&�9b�c~�@��%'�6gR[����߂���	8u���C%�>V����.�:ˋt���:��g���:�]&�yf�Z���4c�򥛋 }����,_����}n�7�� o��"ޏ��٧�xF�"pa����;z>�ڎ��"��;>3^"Fz�a�<I� ����S�:����v��d^`�d�*��$mgow�R���M�X$���s����!�J8da�NO��{"~^[�MY��b�P�U�;���7î���7���Q�y|�D��i>û�c@ח�[P��x�ޡ-��Q�u���N���鱓o�S��$s{�`Qw	��n�6��D\��qWI*h==�~ݜygJz�	��nkԠ�0�.���%�\l���t*M�I�Y��٤+{jT�I���3l�K3U[��}"X��~6'�#�J1��0�Q7��MI@l|��>!�=��t=Uy�sk:����.���5�����t�%�w�^�~r���S�q0x�|��a�QG�6Vc�c�g�*H����cN3�{�{Mvl���븋k�O��k<M6�x�nx���VN	y;e�����(gTd�1�TT��3�WC��h�P״�Soh����z��Y����ݵ�y���"�OS�#O��$5�/Y�]���d���暴3��E}�m���l:����P��hsN#�q9�(25q9"�2��zϧ�Yʹ��v�Zr�Lm\��b�s�qc���W�b�t�q�_eX��jA�?���	�뙞��L�ŗ��	��6#���e������1r���,�~���K�����EL}�W�ݸ� �ڣ��y.J�������xN����mȧd`�r�/b>Wq=~�Y��ΎLF���̉۽��-/���C�N��M���_���+�h8��<���Χ���� ��ӷZ�A��TdN�a���TKY8�e�S���W5�5,�.�jjK�.�V�f6���lᗈ�]ggPNq{��_ K '�X�f�J�99'��r�"��Q�j�H�U��.��>�˝ ���v)0��鐥\���ؘ�;��[U;7�V����G?��f+��J���y�Xإ�|D��m|c���Gd��mƓ�'~2o{T��ߴ����K�7KáFvT�,����xj�C��T�	Θ��(�Ɍ+���r�\�d�9e��N5��m{��=��U��mT�.���r�<H_2�I�V.H+o��}��}&�qoP��_���_��z�:�q�VF�'d]���۹�������֭�����;���J��Ǉ]Jf��5�����Y�6�9O�P��/~,n؅}[-��#rj�-����1��N!G-�F.��c��̹kE(���4d7�[Gc���v���u��$�^�Ln��
�ٞ#�)tDF[�"�����:�>��C>�������c��/�%R�Wq�n�_��x��t�M�8��t�wOа����4'iy�2=Ýff2%;xʝ���l�C�}]���ף���s��?rM-�26zH�K�����at�O�\t�4k�u}#x��2���4s�]×�X�reN�K��Dn�5{�&�Ed���w��EY�v|��u�'Yf�t�����iܴ2��7��VV|ξ*�ՠc�>s.�SsSZ
A���J1%꼔�&\w͂�ţ�+���Gh��Y�w1��j�vw�'&0w�*�Z�(��"���;�������?+��E��;'�"1�=]����Rj�s%mDy�������눍%�Z�c��pG8�f��J�E	��qV3'��ίP��uZG���vv�j�R��Ģd{·X�זX���� ~�������s�
��	����U\8�O(x7[�;!z��zgnfR����f���X����*!<��q���~3���Ⲿ�%΃�i�.���D��ʾy�WpU\�^[�%'��o�7:�X}5Ôr0[�Qu����:̂�GT�Ϗ8���R08�z�͙���=�s$�Ց����_�ykh۩�X�ӱ������G�~�TO��#�_����M�=흿m�.s�H��b���M|�k/<)��zĽ���ؼ4��Ҹѝ��>���M}3�ׄ�=2���*�j:��/Ȳ�w�9}A�:d>Hɠf9Y%�>��}�����~����XE��u+��,ʖmۚ���N2,���ّ�6�
l{�C˼��q��: ����Y'd��_A�iE qwr��� �t�"b-M�������͜��i���T��g�3;�%]�������<���cq��O^�ܘ��{���,�5wD�Fω%Q 2�}O��Ք�5����I�g�1����k���L��M��aH�k��F��6�{x�ncl�!K7\V��-��g\��H���Y�ٿ`�{��V����}����t�Q,�B C�(t t�1�Y�U�G���k�m�Yt��|��gvК^��OO���a5����B�O+b#�Ih��Lf8�y,�`�x�j͸׻z��q~�2=��6$e}���i^Ϛ��m�DPj�S��o�R^r	�4��
��׫��-I�����f��x�1��G[OIf�^d�ʢ<�S^
��\��e���P�|qO�!�Q�q)�fb��wXݞ�]�L6�fH��Ί<��{c�RV{�G��=�/1�F[�:G�r�(���䁓���*Z�ў�u�Ȏ�c���_���</К�C���9���䷏D/1���?J�8�;"-���55�>�]��c)	�K6Rr�Co�va�d<��l^���c��[<����v�'ʌ��N�8�n�:|�����\���VX2��n&�zv\h�x����k�a�H^�]z'�n�tj5�#�[����O��k��~�qYU��J��p��{A�K�hO&�_���m����Y�tL�=�؊�p�7�������}ݕ�ƪZ7c
��ww��V�+\�g�n��ݜ�(���n�X*r�l-�͎�AU0K+b�g�[;7;���[�O^�|-bӺ[���=���w���v���x[��3����;(>�\-`x�sv:B(��g۴��rR�ߜ'G��ne�x<��vxa�C�#O�8�.�e���y�q�z������s���J��s���>1Q��:h"~\e��g��_I�u�������W����ӏc-�I�����^��G0=��땰��XE.ʔn,�:��?�*X��?NZʂ�0�!y��ն��L������8���M�[�0�:�xL��Ȥt�x��Á'�P��S���-��8�{}i`�rkޙK��Nz���_/p$��j��X|�� |�}�s�L}��X�U��]�;��WK�8�{{&��S��.�Ol���9Qy�S�z�Β"���|����+��d���v����c�����Σo� ��M����D3�g��w�wy;�[����������rZP�W$atR��X�B���g)�+�����dm�V�����_Ub?���q�M��
��|N1�E�����j�rD$5Ѕ�D��%ɡ6�qV��t�x75�xm\�8%��h�f.�U(����v4�1�h\D�wJ��r`��4]�=��`J�I�?��En�$8I)d����>D�`��bD��I4��Q�B����pˣ��U�Z�v�au��h=O���)6�>�f˼]�7O�[�SDnY��)K�����ƶs��N#�$ı���K7J(���{�Jy�"{b�NE-�jlJwP���]3r)5��o��?��k���[}5&���5�\G���梻��OĨVb#Ƒk��Rv�y����9>��p�>�O}y^��;�VsQj�!es��V�iZ��'~/2gF�r��.x����l��Ⲿp��	��<�}y[A��R�E��:�y�PYP�v������C;	9oP_�v�����8n>(���g���·qS�tY�_�܅���׶X�v������z�b��z��ލ���n}\^9������b��;�N���yP'�X��\D���m|�[���v��=�n���zJs�C����R�۞���u�2��
���^c�^Y?$CX���Q�ˌ<k���>V~��	]�x5�f+������C�3�ь*���*=T���Q�^��1��/;�o��;�b؞S�rK��vuP��_�����o(s�:�q�NFЃD���p�ǈ���c|�	2�Kb�쑕93��xuԦhNj&�����Qg��'�����7���1�}��֫<�IP(?z>P\E|#V��1w��V·Nv%�;ﭢ#n�p>�������"�����n�@��чu��ǤL�ڒst"��� %�l�w�ݺI]۬P�ǧ6�0�F����ai��ğ�d4�7yqB������]�]�7I"��29}|���Xư�ٵ�U�#h��^NeF�-/e�,V��f�W�e}�\N��a�,� %�~�&K}$_�J�ΰp$��A�>�L�3�O'~>Zc=~�>�~����g����/\�<Q�#LGt�XHK\䕇��@����SP���V���t[��>�5����:K�k�Ķ��`v�)�Kj
��@F����&�Hȿw�<��z�K��v��h=葔7��4s�]�\Dc�#�3ȭ<NAb�_ۑ���V����%���~�?:�S�������~��7�Rk��̔kﹹ��1uB�%C�_C�q:��]���?ђ �!��q}~.�������Zrga��^���g߽�KD��tR͊�����J�v%}�׶n!��p��U�X����:.��{zX��m������փ��(U��8lfm�{�۝1�w�٨Y_M�čw*�'ޢ��}�;�n^.t�2#�Y������Y�pm�/�
{��t_�2�̯7:�[���-d[���\O�E�?�;g5ӣ�����-��z~�T��Tl�yo�쑔�6��)�g��v6�ۜ��V��R�\z~쨅z�V��_�����wn�4L��9��ԾZ�)��^�Tшj�^ĩS�GV(�dp��
qVhFf^�m�d�/6*T-u���y�,V�5"�0И.Q}�:�Z)��Ԋ��)_U�I�Wv)����ݒ��\HX]�R�=}@����a��E '6�7�ʎ���{K6��4d�"�kie�u�iq{�&��4�� ��H�L,�y{�M"�妍÷��s+-�G��F�e��Ĕ��`���:8*e���Q�5fk�`��p	�V)���M�..�1:�u��flx$�b�R�@�"���4R�s�ӡ�w<���e�:��WFWQ[R�f_*7�F�Gf�t=��P��o���9s��(IX�.����� lA�j���&��(ࣽɬ�{;)n%q)g����e�(`�Х;to�G�Zw��m���A�{�%�j����[��6�`���{�r�V����7��H�Xͮ�I�� �93E�G�mA��w̛X���*�\؎���n`fX��LL�[ٛ ���B �5�\lX�&+Wlq�b\�ςF+�Wԯ��
�-;��`�OV���@q�_<i�:��/j�&�O����h��[�bW���Pw,�n^
.�I�Hm�	���\�.�����T��%@�S��U�U�^�N?�W.8��{8�
ԕ�g)^b��5CmD�8���%�د]�^ʛX(-Kl���9u�ڬ��s�R$�o: �[�T���g�+g�4��ù���s ��v:�c��x�r�Ef�)w�1��JF�K�oV"�Tʰ7r��'V�֙}u��
��n"W,��Q�f����8��ui���M���Ma���S�ξwB�&��(4#���֔v���c����t!F; ���{�꡸�i�@r� ��-�O/�e�]W�t�Ёwgn�R{1�+�pv��].Ʉ�"��ڸiA`�9�r��l���V�\��W31#���N�{޸Fs·�k�R�?;p��<�\6h�5�gN�sSw]���D�{%زw��� 	90!Y�e�򻙁*�h��D41��U��ޔ�)Sw����G����9w��v�O�/�� ���X&YV:ծKh��������N6M9|��u��;�������Xֲp���#�y�w��)�]Jus&ݞNȦ��S.��;0.��=c5�u�v;,�"�;^j�\��*�Ү�mGf�$�s)��p�ve�,C�n7Vw�0Q|�Ӧ��^B_f��ބ�m�Cpfޛ��]}�q8�R�Y��H�]���n�;@[v._-f�Er��z�ѩ�Nl��6:h��
�.;H巬�or:��f�Բ7�.M[�'�hQ*�Pzs統|n�e�Qˢl�r �}V���T�����c3$��{t�ݵ�=��y����îf��sW	�7�����ԪZ�7�:8|�}���� �"���B*B���$�����j����*��J���J"(bH��b$(����h ��`� ((�(������Z�������
���
b��*���&*(����
j""�&����(�*�I��f*(�"(�����&����������"&�� ��������J�*��h��d��&�	�hf) ��j
*�#&$����H��f��*�&
I*��b�h"*)���"����*
����jb�`��
���������*`�	�d��b�$�hh�"�)�)�
$b������s�/Z׺VյO8��:}��"�J���c��O/�v�j?G���N�& v�4�2�ÍΘ!î^�A!��Kr?�eT+�]ɺ�P>gO��ߩ�@>Z��
t9��/h{/���ޏFr����c2E����󓢴�{�@����-!C+�*�sQ�pu�K/��k�ٛ(�ѝ�S��cݾ��l���2�|H<��bzUOǼ�*Y�v��5�|4gM����������ٛ֜֌wǜ�9A���ʦGTR:did���,��z[s����f�|�'�u�2�^oh�y�����q����B��L&.K(-3L���H�T����`�tstLb/_TW���X�9���RM��T�����s%� �3�|hE��껻w]����]����t!z{�{��wi^Ϛ��m�DSV���@j6׏��؜����7y��g�R���`�-�Z�O���a�Č}�����Y�י.^	�l��5W���QR���C���Y�30�)���<��}7Ӹj����Ɇ�������1`�O�;Z�/�p�ێ��.J&ƞ'$�;+�Nȕ���X�t�5y��p��~R����!�,kx���$�ݬ<�5���_K�Gv)�q+t�qk����K��{ۦ�tEc̩���t��L��p�d��[4�Tѝ�-��fJ���G`Ū:�Yv��|D�y��x���crp�en�8�@z1���r����}�;N3�褼��D�7�Uڻ�͋Ǒ���U1B��4�sN!e���Ҡ���ًC�x��.}�Go6�Z��u�\�5���ߺ���+c�ǳ�mƴ���Q�c�<����Qc�Qt<��H�q��¡Q{^�˟=�7,[z}����O��&��m8��2��z�>��=u��i��o���:|^���?A�D��q����'Y:h����k�Yd�ճ��G�uē���h��V�>�av��|#��z*�%��9.�D.P�i�q<�����\Bbܜ*}X'�w'����
����ڍߝb1Y�+ƅK�+��=92Ѡ2�c�\c�~F��%���߹*�Q��_�b�}�|7!�O��>�k�j�F�$���s2V�E	ɝMFQ�i��F���U�����oLeu�7��k�M�Xy&W���qZ����+�>$�*�AX�!D�-F� �(D�����;�b���.��@�_:yBi�S�"�e��L<4����:g���뚭Xǩ�d�ϡWo����
��$�z�/��Ϫƣ�w�]n�&��m��J=��z���ͬ��me�� w6���a�/+�����zF��u�Ef�c�"�'u��Pb�Y|;],�eY�ޞ)	���]�{�� �Ǜ���C�!�iSڂ�)�9�:����<���P2c�Lx
�-�淰�\�!E��fܓ��QXH<�D~?�����끱��,kO� ��M�qN�����#ޥJ�opg(}W��r_w�͠�C�YQĞ��e�ţ�T�N��9��8o6L{�Zގ16ؓ�6m�a���c��6Z���b$ut�:���v!e�{��6�qVB���q����>yѮb߷�Ê�R��,�pӈ�|h\D�Pg�\NH����.�%�}\�N��3y~��?rā[Q�����S'o��5\��av���*�L��	�;����f�S6���q�N�C����HՑ��)3�e�����}�D5���^7��"�^H�U����e.n�w�C�5㒂�:z��j발7�\����J��/yγ�ٝ�L}O������շ�ʭ��_���e�g
�NlL�?T��S�t	S���]L״L�	A���B���ܳh���jq��sQ�y7�M���CO�P(u�~E���|D��հ
Ӕ�M�?e
���^���X�!��o'�Ӄ:��؞����r2��x�x��
fJ�խ���V����>F�9/���1١o�j�>�|���W�M��N˽�[��əLc��������a<W�ьz$����Cf���d�ǧ/��:|f���ĥea�u:r�׽�J ��G�F����YPW���;�y�.�b[�����9^9%�sG���-�˿g��u��ta��k�Nz_Ϋa��ʫ���r�<Sv��f��u��W7W�}�}٥��C����5������X�r�^˾�z��K��S��\�+�ڲ�o��ĊsO4�[�{��'X	8�ڇ,K�8�Nj'K�ר��^��~�2	��X���U^��|��e[.����_�����Y���Ĵ�b��w����7���������*�������w�rY�P@J��DL��H�Ҿs�
D��Hi隫K�Fodl?�_WE����=�w	���/�t�x�����:
J�]��D�il��BMŮO�_��4��7��:��ٌ��}]�����q-�q�AO$��;��j]W�_�������~�a���4�l�^�f��H�햋|�L���u�S�rd�ڪ
�>K�ڛy��z ����q!fO�hM�3�wOx��~���5�Y(���F1�֦S�����=;��}K~��#�2i�2��r~jV�Z���/J�w�!�U�n��{�CE��y#n���ö���5�W\�&'���RPڷ9V�8�ϔʌ��q��1Ԣ�&��v�);8�jb�bO�Ft��b�Ӛ�,�(f�:��Ri:��GA�o�݊�u��B��ye>���[����3c�)$����}�o*>��ef�K��㡙��������^3U�Ac����L5p6�;��N��n���ަ>�T��?UeT�B��;~�Ze���������P_K؏�X���+��á��/���r~�e������ڣ��Yt�~ś?P9����1��W׿߾��y��;'�{>ʑ����;+_�ٕ�pJq��nwvg�5JϢ���7S-���i�)kn�X�Z�7�u"�+_N��,��V��aI�h�����Cv;oc6���Y���	�0ys�T�8��������M �k/=N�3�%�fZ�k'�dȺ���{_Fnk��4����$���ØK#�	ɖ��2�ar�jc��pX~���9@�r�(�������i����k<g8�=�Q����XȱuԮ~92���n�V���?}Xk;Q�&�����7����A�Gg�)3��vA]�֔F�]�ad�*J���{�`ߧk�t��=����+�'yӨqD�����3^�n(|��.cssa}�9�?:�۬�j/�U���!�s��=��C���~����.~��TV[*�~K6�����4�3��{k3z�n���j�\Q�VEvD �Y&!9�z���n�G7^�mt[���Q�T	tD�����ۗcχv��_6�;aΝ�s$�Ψ�,o-� {ݽ��g=</>#����U�sK��u�T�����p�]nNE��X��q�;��w~g�䉉�\��H��j5�LoB[f�J�}�Y>�_6�"3�ϲx\H��h�]�F��~���D�Vq�&,&�bV������[͉O��4OIf����Νw�곻�{a4�t�D򖒉��MA����X*\�ƅ����iKҚ��}��Iケ�VE	>{���}�$;���b<�:G�btQ3����š�B�*Z��:��6��~޻N(�#����>��:�������桥��B��~����Pg'E���"����O��{t�e�:E)H�IW�C�ν��B���9��2��U��N��:J*���f�s2.�?a��*o�^��]�a`�!Л��_O�����hg�iŎ���/r5�T���z��S:|����3���N�������4T��ⲫH�Q�9.yo����Ydܵl��]��-ox箖,�~U�ѯ菫�/&t_���ne��	�
�%�Ȱg�+>N#���75sq,s]��}r��*q��_���v:�b���M��'�pe��x�q]U���!�]{��j���`˞���7��[�^��]G3�>����xFm]�g�ʍu�T��
Q84L��Z����^�W��}��#��A��QP"�n�ř�Q��9���Ǯ�N���18��%�-gu��
�'Kԯ3(me�$j���R+��fU��W��Ϩ_�}L�8����;K���U�����Tx���3�FU1z��@V�b��ߗb�7�N��_:wP:�ku跐�>��a�s�>�s�X�(��(MN'B`��Kج����o��`�����l��d\�H�[=e�E��y&�J/L�w��:F(�e��Q�Y��z�5�QqCr��=Ƿ�j=��������y���6p�bE�;�������M�Th�U-E��Fĩ�(!S�2�p6:_ō�gQ�|����lķS'�4~�uMNf�����,��&�s��_9�TO${U(wP��5�[�Y�)�U͏l���m��[�T���і�s�u����,�-{��P�ut�#W����<�%ɗ��
M��g�z����8�ڵO�z=�0��R��L��s�B�$wJ�'<��ԧ����`�}r�۷���;�s�r��;Ǳ��1�}5&�󘆨s���R��iA�ip�`��+6.�I��,�zN1b٣�p֯Y��|��t��^W�m�����9�k���!c���
�*��??0��՗̚z]�(L�
	|)%�`P�[\�qӘ��PH���(�'Zӻ��j���,9փ���GT�TE�Ǳ{�@�h��P���e��pq�����:jQG�K��Y۔�ڢ�q
&�Iڲ�\��h���_�˶:^��MH��᥿�!�3��Q�9?cgC�Ee|6���x߱s5��m�/�xm����q^^�3y�q���w�2�*������K>^������r���J��������Bu���J�oo4�\6L��:�go�r�GS��áp���ʳ���V3�|�����u�'�yglﴸ���b�Zʋ��N��ή[��;�"o.W�E�O���³�uo�b�u_˞V��K�T�Ƣ;�1�@����|�����L|��]��YueH��s�}��\���<7�����D�-�%d����42��ƾ������%�}���Xu��Uz<81I��skz�3w�_�h�H����q
;duNL�'�L�jbq���x��Ѣ�}�g(m��-q�����gXΜ}���_���4��z"�j�U}��E�T����H.�Ԙ��~���w�.�:��cQ������B)24��.L ��b�8��v.��'5�՛L�e��y��{���9}]�S���;���΂�i���x�z'���B����OUA�X�%W��N�_:WXu��wi�Ϣ�М�f���;��@�m�"�̍
y�r;�ܯ�ֹ��K�BDO��cɠ�Ѻ�_2Q��A�]N���cD(7�ˍ���XiG��m��.�U�g��H�E5r��󻰯g�H�N�*ܔ����DW���������/��.�G@6���
y&�ӷ,DhT��`ջ9�Fߧ7o��|Yh�mt��N=5�C��ϢFW��Mm��w\Dc�����	DW��P��,�d�㪷H�<�ND�l긔�}_Mγ�wOx�ݯ��̳W˙(�O͚�=������r�Y���q�˱p�ْ�2�NKc���i�qZ����O��9���mn���ɨ�Kua��y�0=�%�A�t,��z�/�Y���vDZ���Ȼ7�ӄ�K��"���Vy��śv>��
�����'?u�ߤs���UaeM�čw*�x�{�
�B��1�̻�7z���G�-vZr��?���.�+�i��˯2���=o���o-dH�u#.�wXɞ������n�3ORj�������:�*��L��Y��[��o��[F�H��ƾ���Y�׽�~$C	�w·��Ru��2�&x0�+Uܛ�ە��,*��L���3��=�}�h�U�q2*2�ŲU{Z�weK�w�Č��U�D����A(<�_��������8��v�7t�_�F�@ͷZ&��O���f�l?�ش2+Ffs3�t�hh8����o'6sP�"W�=�V���DH��N��v[�6��Ƅ)�[7�ǩR�<�jɏ9�X�#�t��Z7��7������6n����sۅ�:gK ���6%�_9,3�V���fj�3��w�x����*��u�Gbܐz��A�.+�\�reK5��/k~�swZ&��~j;�
�_և������g(}A�L�N��K$��
�J]x�ݣV{}�%z<P��S�:O\�fT���ys���ON0�O���HN��N���B"�Xzj�����[e��_CA������^�1���hM/oc����9��O�Tz��B+�@4�.��`��Ƙ�mI�a�p6:Z?n�5��B��?���L��:~��f�;L<�W�YQ����?9�3^S$������=$L�ԅJ����e�A�Č}��:�e��y��4��ͻ�l��̝�7#��J$i�	�F�
����t��%O�� ��z�7��B0M߱�����U$Ww:(�ͦ#�s��D�q9�;(BvD��W�+(�kw�ٜ֦��{,o��]�c"���70Ҡ9��]\L{�~�F&N�Z�2��%/{]����v�rG���`N���v\z8^W�ōs/��s����;S��E�|�t�s�Ty�����"��N��t`)�zү���,�R�Mެ���(%�I��9vd�fM�or���G^�r�sr�YV̡�s�j�u�WI��u]t�ΉNe������f����Uсe�M��u�o3���\V�u�k�%�aMc0�U,*��ɕ�P��Q����7�ֽ'�ytNV�r���!�{L�IT��R�C���|�G��ov-\��z��9U�A$RL�V���b�(�z�u�	.�yk΂�݁5!���f��z+X��y����!�wP�&�:��3�EG�Kr�^]�ȰW[����R�͕�7�f	i����r��E��Y��K�C{�7*.N�gBS��L���7^�}�oB4��E�[}P�[7�e��+6��s�.��(낙���G#��=;�,��»Uø�(�|/j���)j2�w-	��-�Չ��L%mlV7i�09mִ��:>�R�i��O��e��Ջ���k�yP2�z<��{�n��g2���Z^��h���TrM�TT���3(�f�v���s+�7-;�T\G�l��kW] ��t����1��m�V(��5�&Cti�U�R��:DE껌�Q�La۳�k���	rvŃ���s��ڽB�������3m$u�v��������]y���f:iV���J�MZe�J�l�ݬ@�z�Ϛ��΄��̼�j��!Z3Rt+^��Zq�+�8HR�ݷ�Iw2P��w{"�FQ6�/4��Rh�O^[�lHQ�gQ��swi��z@�F��*ھ���5�y9��:�'9�pN[��&���KZ)��ވ+��&�щ֎�;3KG�����5��[Bq�s�	�g5ɇ���k%�Owz��x`�6��t܃4b�"��v;C��a��]9Y�Vbl^)|Lz5���zY�(��fP������ɨH%�ihN����/�z�N��	ө�u�፭��WoT��JU�xt�9�[���H����2z�$`��n�)Η9%��anX��ed�̃��*��Y�"I���jJ � k�Ф���S���YV��F����H%u��T��ZFޔ�Jոu�ef/'g?'���q��d	���Kw<t���>��.F��G����"���;Շ\�OU$�ֆ��b��_;�c��ԣ'WZ�*V���ɫ���ާ���jꗧ:%���I�O�����i��,	�JOnNZ�T5V͡��a��a��)�ηos{�^���0>��
4�H�/�����kU����mS�h��PbL��� �Mf��B��NH՜�/D��r���fh;�N��~v�R�� :��ñ\h����B�Y먦�ƃ��ѭ�\�В7�ε�7
��^�sy�	&��Ώ����j��o'�I}��ڰ�n٭��8&�Q����ݧ��]p��6�N��#��)VP1V���j����"��������
���̢���`����"ZJ���"�"$�b���"&����"

�"�*j�J��$�
**����2L����&�*�(h���
�*�� �b��&� �����*I�* *d���*�����h��	����0ʪj�** ��"���a�&���"B���*��(�"�&� �i�(�&H�����(�������	�h�j����h�� �*(H�����b)(�f�Ġ���"*H�"Fh���&
�)�

�&22�h)("�JbZb���¡�����j*�R������J�������"����rߗ~Y��7F���-�jMH�O���z����Mh阱;��^(Lg�.�ҫt�ˢ��W\�y�w;�����6#:vоjj��Y=�����ݨ��+�D����.�񡞭��2��r5�ꐽV��}39N�H��|�4�K���wӒrܠt�]�yz:���GY:p. o��g������=�/t]�k��8y��	�U�!a�%�����۪K����x	r>r���=W��eg!_c[���X�N�pm��;c�hfX�"o.W��d���e��g��ꯤ����lК��j�[[�#����]|�=W��9�3����ye^;�+MQ�NO�g�
���Q�����ǯ]�X��V�ӑ�ې]����#[�E�����I��;c�97<��D����}������=�Ѹ�̡��:FT��=~�Y���	����ϑ|��I����T{��.�Z|V�R��]���
&�R �MD����nKe�걨���*�>��#����8P����2�=�V�Eֳ�[�r5�fû�B�G�"�[��K�����6�R
[��t|��;��L���է�������x�m�^��YQ rE���S�@� ���������m����c���\'��_VWRJ�bd���uq�Q�5{R�ĺtU�b:GrA��v.�a�Z�&�s�3
�YՖ�"f��y�i}�����HrR���Qj#y��wӦV9d��]G1�ʜ��3+UZ%�FE+�f��8��h�w����N����Ћg����,�ůq=lȱ<����Ʉ��r�<�C�\}e��6<�k�,O'ث�t>{�a�=�Q��,�`CN#�4."G;�F�'&zЁ�V�ޗ��ۨ�,��_/Y��k9V��a�w.47�Rk��1P�N#�1���R�ݺ��q�t���A��*�ql=�:�7[/���R��g^�,���㑯��r��3N��4=%�[>�������먮;䮾������#���ܸ���'�3B��~R�xsdf���xvm<��:�=��?M��~��K>^��q�c�����证������<i
n<��%yy���b׭�辙�n��sCsQݑռb�>ʝ(2s�}~E��I��%�L�#&�َmy׋3s��zz"o]k*.{]86�[;bzv3YȯRVpQ�~I�u�u�V�Ċ�Ů9�ʨW\ꑩ͘����X�����׺��7����7\-5��1�}Q���Q��X�y�XI�(�+du	�-�]�vuP��_�����a�z�����}Dy³B�b��e�V��z$<Kd[spkG^ �E֒R�t��Ԏ��	ݬwdҰ��Y�=���18��i�nĒ�'5�vq*�.u�jrXo.���.��[f�}�m�Rg�9�b�\�U��Hژmmκ�%m̧bc�.�N�27L�^ʍ�Z~��K�l�P��I�	tB��:����N<>�L�Μ�M}Op}}�v��T�|gʪ^pߏ��K<�T=Fq�`�(�( |��'�����l�����6y	�E��>�.\�w>�*��э����w�4��������v.K5�P@J��A��w�����T^���K��߸Ώ�}h!��}��5��s�M?:Ɯ�
x��t�{�A�;2$�[\N��~o�O��Qo;
��~��G��fٌ��y�t[Nt�pף��۟DW��s�~�<c覕P��5���-AP��-=������_۴9�{�#(om4[k`���������v���͕���{�!���T��r$�٣��B�D�ZϨ���5�k�a������P��}�*4�>
��ɓ�jt,�n�+�Fu:�]@CW_	[�诫__������4�P��U�2�,=��:�H�0�<�B����_����܌�j�ևqS��i}8�.��bo7��{��i�>y��P�U\8��{b��s�{�V'�k
_eN���ݳ0��@6���?ҝ=�pre�����$'ߑ���;��9��}�&V���70��������{\é��_TgkO/\�)�g��A����^gc��3:,����4��Dy��2�`p5�0t|�Io��+��j��{wY؎�fD�rĤɝ��?kϋ�ϋ��t^���=�:eיM�g^���e��t�R�ݿ��y�H��&���`E����:��Ui���� -o됢)���mԋx�};��������D��|������rJ�\�~~����g��}w'��24�g��H�/s����7�X3S��»�+����=�*3�$��I�v�K#�re�+쮘\�v9��F�%��0�w����������y�q_;��7�Q�2�Ź �,�X���s�MC��(��m<9�˝Z����Պ����C�k������eS#��tΖI� ����yt�Y�f{�^�d����� �.�&�7>�|u�6sC�!:n:�b�e����1����S{��ѿ�A�@gO���^�5��>�\U�_,C�|�l?�&����ixn�T�=�c�j���MB~H��F5LP]����h���j7����������9�r*.�#�	���K~�~�|�@f�3�d����l��"}/�B�KGF�#<�<ؑ�4n�jg�?B�iq�Ѫ�&DW��� .i`��0ST;�6�ʽ�a7�b�J��+�%FU�!1!W�Dtol��$Cs+�toc��Mdtn��ޠ�F�AVJ�]IpDa��R�a�+5rH0���&�ݺ/w+.��cV���$�'rk� ���������62�"��x�6�z#��8�3!vx����*�Y�	�+M��U�J���#n1rGקW ��?.u#��3��[,G��x]M�<NH�C������ʻx�/�/g`��l�C�N����q��U���U1B��4�sN!e/�E���jA��+;nN*$_��s�;������%�
��鸥/��a+�p�g^ۍi?棊�U���+9�6|+|�� �E��Ǜ��~�P0;�X��	mx�7/L#�&���>��p��x��=RT��a���\����ڬ���awT�1�,����4j�������d
��v\
[��fҋ埠��&����b�i�X�V�ot�f��˴�5���K��BYS���Y��|��{�֡Q�(�Q�[^����E8�]�t�.�O3�'��g+�0yr�h
<K�+��AXz)z�����<��ܕt�ͨ�F9���.P�C��s��s��ʼ"w.V���q���S�S�B���N������j\�`������z-�&Ϭ<�(s����,��xP����cBz_�d�W�cC�sV���oZ�X���=c�Vv�:�ն�Y���]f6���YU2V����@u�t4fiI��c�X���aw2�F���ư3kp�Q<�h*�8�,=[ ��M䎮��K�Sd�GnU���b��?���3D�T�l�u����U�񵉖~��J��C�NOq��Y�O(M=O��/���a�[�W	�}��sҰmއ�ӑ�}TÁD�� ���$7_[-D>��y���>��"���2���P�kw��i�����9Qy�jx����ʀ[?Q�n���,c8��}�UESk棓�����1��w��v��M��/S�eD���@��&:�LB���9� �a�lb��7�Vy�[�ͣZ��tXi�l׸��dX���)�W�	y�'!�a_z�ɿggw�im*7Y/�ĩ���쏅��܋��|O�8�wƅ�OÝ҂���J�F٦Ի;3���M�AQ^4z�H2}�s��_����ܸoT�`_9�j��N#s}���u����v�X��>���r�T���
���7[/���R��g^�&��ӽ�n)�2�tfkR�IkeO��z���~ٜ���F����++����x��R�v�ܦ�{�����?F�J���c:�d/?�~3��ga�W����@���"�(��x�]{{H��@�Dj����aҲU�G<A��tp���9>���Tk�>E\��;A���5�ss+)�C_��K��S��;+���ޏ3��5j�0�ĥ���w)D-�E��J'e[QfÎ��os���̢r+��9��YЧ��9&ߜ����4tλp\�3���f^O���r�kᧉ��:о�5�Eϯ��e����7��ՓZn}@|�e�؝�������R�۞���c��'�˕�G��{����U��z�g�N��3���P�	ͪF�㘎���\y�1A�kk=�9�}:��y.�o��JaX�{�����ʎ��2N�2
�@N)h�R�\hvuP��_��E���o��W��s�c�q/�NR��g�o�ua�pՂ������]��X�rq�u)�-LO�FB�^O�әf��3�c^�c؋/��K=�����)�6
5
*�,	
S*���м2l��~r��I��=�U��O�x���bi˭�E�c���j<v��@���aع,ה������u@��w��={$}ί�v�
�}h!�W�����s�M�Axӗ!Ox������tu]��m�u���X�%�ź{<�F��������~�O�>����@;��0$����M>�����εr²m/1G28�~����R���%p�7�i�h�nv}g�#\ɍ��#�%z��T��^Z��q�J�9WZ�=a�r�ɡm%v��O#޷�Y�)���(�ͷ�v�7��R��2�ݛG1������Wv9�܍�/N��-J�%4��;�+YZ�M���^-N̸���	���.�Η����-�U��eh
�Ch�Н�Wx���z �����}&iO����D��u��=e"���*Z.t<.Q��#�Zssp��,��(�j#�x�TV��uO��FT5p�*V�Z��ҳ�v���3�]��^��/��A��괏s	���/6��r�G!���Z����Nϱl������[��*��#��\�9c�.zf��s���}�����X���)}�8n4�wil�w����+7�n��X�bd:�nw g��}{��"���_�2�̯ ��/>ucx�d���0?��JH
-(��G%v�k(��cl�R���+*��L��Yg�#}��F�-mu"�(�YQ�JU���q_�_�>��)
���;E�lL�5�9#k���H�R��aq�y�&ڵlǡ��?wo8����\?��W��{=��/���I�Ka��GP�-!C+�K��gs�x�6g������r���_�����}A킯�QZg���+�H?"Ñ�B�ʗc��;ikŀm}6X��<\�1>�t�"��s����a���>�f�0� \�j���P1�.�K����T��1��lVD��<�!�m=��.8�%\;.��yǌKm�ʴ���J��C����6��ۚm�&�	�ЖCk��NZW5o/�JA)�-�o��@�ζ+��j㠶.� �y���5#���;���u�/��-��s����WowE����p�M(�-�߽� �t�"b��E��'�V��GJ��i	�~t��������f���Җ|d������F��XᚍF������bs��=�RNkޅRf�B�u�^tVU]G`Չ���ڤ%�~� ����-�p:Z?n�5���*:����X��*s ��)�}5Y���}�0�^O���u�j�R9"{MM���"b_ԅJ����e�~<��vλj|8������s��#_6��͖��v#��8�IF�,)cUE�3���C{��~�/+��������?���s��oj����Em1��2/�����ɋC�`�H��wo�+w���>��z3ժ����u�Wz�|�+�|�T9��]\L{�A��O��e�m�N
��\����:���5u�/x�_NϼV����q�y7.0k�xo�s�em�U�������䰟���F���ОT�g���8>f��C�VW����|o�����VӋ3/G�7�=��G�C}��ɍ˓�o<��v�\U�
��ټ���^����p�:�ӟ.�ze��k忭iӝvW������*�J�]k�>26�N��y� ��q�I����\�ȨYǟs�w�|��L��83s�Y2���EK0��zLW
���f8���ԛ���KlB�y�M�x�����}�KMJ��q��כ�_q\��ڋ!�;��K?T��=���參g/�P��Xr˴��PK��BX��G���6H��$�����j?
���]��t�?����VSW��Q��K��x��WE��,��x$�F\�gV�{��bV�Nc�X�sQ�r��އ.=c��;r�a��7Ԗ��Kwi��������n:$���|d�r*rg�S�����ku��g��L<�=�V�iX%�O.�d�ny�5����d��Pb{#�NOFн��/$K].��|����d��gqD������s����ꑷ滛p(���$0n��t�^>��;�\W*�S7+�@w���F+p�}�w��ҽ/��|v��q��3NdiA������1��X�#����'uz|r�J�[�c����r×]�[^�||Z�M���eD�G�٩��Q�~�쌢giɱ���Τꏳ�<�S�o6S�A�ь�{N:-��Y�o���"~��
F��C�}d����5�v�/�s9u���Ļ1Q)ңqY-t�BU���N����Z�,Z7_�
�+�H*�� *����"�����PW� �"�򂠊�PW��T_�APE�A��*��*� �"��*��APE�
�+��T_肠��TW� �"��T_�1AY&SY	��>߀rY��=�ݐ?���`�� �R�kEI*�i�D�B�
"�ڛn�W5lVڊH�l�RAKC(�[`�qt�EJ���VX�"i��Sm6�*в���,P0�9a�P[ d h�M4�j��fkV��*]�PR�ۀ� Pd  6�7V�6X2�3f��pdN�����٥��h�Z5X�	��P�6��	��cV�f � $ h �[h�� f� ��  H �  m��ڊ7 � ��  m�	 6�� � 6`[F�K�7 �j��
Y��iMf��d5MB �h�uJ�P�J

� �TQf&j��
e:1
(�,e �hѶh��TQ��U@��p˭�C@5@�fh���i���      �@iJIQ� ɠ #@ S�)R��&F�0L109�&L�0�&&��!�0#�ԪQ4i��i��b0C�bdɣ	�bi�L#0	4�DhLF@����3Q�=G��a�<�����ۯv�m}�~����� 	!�?��HHHC��J5$� {�$$�0���D_�Q2I$$!��������G�O�Y��P?�1`�&Đ��Q�C� ������0H�4�Rd ��!����_l������|~���$�$!׶I����`g�B���c�A���)�,�i�9��M�K
X$_�������F���K�kyw�u��ue��DX��ɡ�t.��,mVP��i�:��*�y�]֨�=BΞZ�1`�^]�8`�DA�'PB���HJ@�՛����2J�=ػ*�Qv���~^k0^BVeو��/w����b��(�������yoy3����&�����_v�V*��^�\����e[���)k�=�&�,Vo�2���wv���-e��)�
���f�Y�v�W��0�x���@h��.�ov�w��@�к����"��{�^J�k�����Me%B�w���X�}w�VQ��`.�h��)��3�Z���B�]�v�º�/k�.{���
4��nvA�Bo��f�+�m3~�'	�V�M�VT�쑇3MA9�v�wB���-�OB���(�c< Υ�{	=�7�XҦ�91�u*a�z�(�����U���(������|nZ=gon�4��_SYYF�F�o��=���gr[؋(%j��c ���]��W_��]�\�]��SE�9v�W��&�es��|��8;R��P#�nR�$#�;D�'c^j"�sL_3�e.�9V���6���K��c�&�W����¾�5��D�=�y���vu�Ձ���:��@ѫkO=yj֢�謁zӾ���U��+�<l[x���{���:��X�K�j�&yRJ�r7�,Z�����Zk��x��Y�V�5��u���U�)U�XD�U��x��sf���E�]�y����-z�l�An[ʁac)����%�� r��ق��ˮw��J��-�=]N�Tv�s��V�X�F��:T��/XZ0�FɵH��e���RN�b�V�{ƺ���:��z�-�M�h������ز��E�1��<��\wj��m7}H�ˮzt�h4okn�#�����I���U`�'V�٦��hg"2������RͶs]
 �b¾VsE.:�]��C#�a���v���F��W{���&Ռ���R�3
���z�4����"�^rݰm+ۭu�m�����r�[�:+9.�haC$],|j��z�+~D缕�Ҷ��:$�b�jڿ���-�/�6�xº���T�WY�ܭ/�mgV�D�]\�s�����ڐ���39N��ǈ���	&r��'���F^��$��K��Ō9���]���6���eb�G���K'�������H�9w[K,�V�;�v/�@���J��<�.�ԒhuX����;zo���:Ih��xeZ9hr:�,�{K1���w��C�Ǭ4hu}ܰ��Qź�h����uuw�֨�}�n�m]Ռ�����m���S�@�ޱ]A� `m�&�W��Y�p�]HS�Ϋ�6��q�uǐV�f�c8�L��Z�����v�h�
�>����F�zj��b쎣���ֻi��M������9WtX\m�'�I8o���|s���͍5cE���Vg�����ͫG��<.�w��x�9C��ùX�(:�PJ�-?&H�b�b�\iP�,��3����[��>*��&�`>Ѡ��i��\���v;�-m�dQ�uzC��Y�'ς��v]�kX���D|��Z9�R���6�
�[���ɷ��Q[�V����~׋��93V[y�2�9\���f��|o)$��z���Љ���y�ɽ.�G7)��ɲy���� �D$H�����A����j��}ٖ�[]d�Vk�7�<:���{E|��M'�(��#�C�ʲt�U�N賜��V�I;�61�;�#�1Mg��;�OoAesV1w}�����z���2�7�h=`�y�;�������u����cA�C��M�C*�R�,��Cs�^Ғ3��VY{KwkAeu�;k9���-
�������qЮo���5Yd.Da�v�k�;�8$�h��~V��}�Ok�ݧv�*���=��뱝�����1�f��v;�B�W 7J��j��(�O�M^g]����x��t��t��m �6�*̽<z�s�"�cy���3��i^�����RH�>]Α/��|��Zvf�>.b(#�i<��5�V1�]3�f�-c��Ь��G.��x�׫��i��dݜ�žC5׉��&-�8)_`ߒ#s5���XJuv����,v�}����&�]*G�R;J���B�`+p��ݝ��C5���۲���
;�n�Vf�u�0ko�U+�����%A��sk���;o�B�B��Z�&�/7���7A];+���W�m5�ٷk����c'n��|���C�\F�U�w,��d���TD�I��W�I0�(֮��y��9��oR���Z$m|�Ѷ���c�I�4GGn�K6�0a��E��V��4�w}t�,Y�w�~�,V��*�%�FR���&�vk��wh��xޒ[���o�p�R
�;����܈�6B�WD� �Ν�k,bšm��ww�p$c�Xn�%{��j��čvn����,g0���C�c�%g�����k���A#2|�<{3<�$�F%��%���&�$:?p��ͽ�؊<L-��R�U��zY�9g!G�Ď�v���`���u�e]NW � F�����
����&H�*�$���ˌ3�[�r_�'���)�f�0p��]V�Y�d4�m��Oɥ���M.T����Nŧpdk�B�}Jpv3Y�7�7d�T㥔N0�����f�xW'�nH��و�큌�yM�n%jD��S�%���!��Z,+8Фo�=�@K7��=rMYl.GF'-��6Ŏ�<u�FӮKu�εY�>:R�Oj:xq�0�Y��OR\e��R[F�pY��gE]wWpr��$f�Ǎ}�v/K��v�x�[FP)橵)_ov����y���Kw`m�����eLuV��GU��*fo5��V�����k`w��^!�P�םܨ�T�=,��l���/Dd9�Gz��	���Rx�2Qֲ���i��	��C��`�^�7�����ed��Ҳ��,,C�+K�on��y0�Ӳ_:8B3o�F]���J�)�W�6�h^�	K3���y�g=g6%Wr�|�X������\J��n�
��m�����{��l�Y��G�.V�1���|.�������0�[ő���O(�cy��۶�F�Ɋƺ{}��H���%&��VFa������"K���R�w��l�+)�s��d����J��ߟX*S)��}}]M�n�_J���g=2�K��R���1v�U���4Unt�`���N��"Y�$l�9	�X�a��P���va�oQ��\�Ի*/�U��n'r��m f�6i�8�Q�w�v������ꌘұHopu&͠[�+����@���`WB�_��;Ǖ�i,�'v�#)u�7\6w�;9�e��=�(1��v=E�zq�s�(��	g=��ť)�a��\n���s�HP#2��Jm���kd�n�17rK�[@h:�V�j'unl�R-k#D6�X4�������uy�{;�3W+�Fv�H���e�(�ɇF�������SV��#&m�qsP2ĵd��x�>*�s���fﭪ��Yֺ�]bm�+wF��E��Ε�� �d�4�g�X� �o'�8��ay�7D��G��ǜ��
�T��v�u�E\Ճ+7m�!,�K[Wc^V��`fe!ҝf;	[U�O��b�ԋof�o��r�P9	�E��������$br��(��Vȵ�F�p�Yia
I�Tv�}�B�VD�7������ͣ̕"%�:�H:�Ŏ�O9Asz�Q�G+�݇�3F��s�`�@������)�˪±Ԫ��;ew���NC^]�Q�̢m�� ��䖁��/s{��н��������b�]�u�|�3���|Sh�@�F\�tPeʸ��ozV,Uz���<�A�d'ql��}�E���Vֲ���<��8�n:H�&EDO��R�D�)�Nw0��&jJ	b����D�@�zl�0I���]J��+�ǖj]�8<�4_,������)��[#�jeX�3�ZʜSx�JKq�A�p���΂fV�i|]��**J��)y��R{�����,}a��"J�ց��Y2�(���h�ر�7�Ee�dv��vG��hc��3Y�:�s��.L�iw��>o�J���NC�b�+q��&��&��ƌ����Y�v1v'\w�7�orш�z�B6��`�2�NLȩ�˺���:ȥ��#G�����*Ē�L/����jm�c�\gT!gwYtqy��uj�x�^3��,O.� �r�KY'b��i�zd�w*n;���SNq��*\�&���]k��w	����L����u��u��8��z���m��f69WN�:ص7�(��3D��&)�7Z�2�,0K�9.�r[w���ĸ]9�l�����p@㛼�N&zR;��ף8˕�U�z\���*K�p�G%bj���H��ޗ"I%�$�I$�I$���`�ıl6LSz�mնܘ�oh��e)-��t��g�l��<%��w%_8�>��ғ�֜8�D\�h�B�gX�/���5CYv��p=7�L��2̻��$pu1�NGV4͊K�(X����m�w
��B��f�&:����.R��r���l���%�S��7�0
NKɢ(5�1JL�8Xzξ��6Hh]��,`;�9td����[����d�3]�����{����s�6�#�XyP�]�YV������[wz�����ۉ�Ky��ǲ���L�]��e���۾Z���յP^M	��W���*H�n�k:�C˦�'�eާ�A�I�r�9�®
t��6c�g]��+GJQ����M�^�n�P�eV�Ń~\�U��P�aV� ��ev�=��c�M�_ؘk�yRNvV�`Ԝ�X.�1�6���OS*ٖH�BmK��*T�3C2qX�OGbز�̛�L$Av55xb5�m44�Pۣ�5`C�N
���Ml׉ͦY����f���G������^����o�ש���BB�	��ֶ�!C����������>�MB��gG����W/�=<GG�ou�cƸ�z��8�ve�նB���!�+R��utO��݌d�ލ��\�M��v!LwM5�_X08Ki�NS5|�����
��̏b��D�:1�Z@��l� e>1�4�B;��q���l�k�{��9%��G���Yhu!C��0��gH�c+7S��k����j��c|��)4�f�(��"��^��K
�6�Jev`܅�3eYk��R���I�ݗ�H;�&�
�c�b������F3R��8PE���%Qj6m�y��5hlOk�]���w׌���+c.��Z��F���L*<U��17�U��wk�C]�Q�C,��IZ i��o�C�mӮ�ܼ�\B
ŏ4������ēj���iFU�����tP�vY�����<)R
�u��c�;j�#\2t\if�a%K1��^�70�K5��T���P��1�w{�
q!t�X-�����h�ʔ�pt�Q�fW�Z�ܳ�9t�F��( Y�+p@�hj���bt�~ib�q��q�"�rY�4�^F�ǽ�E���2�D�]���n�}r��wV�W�BV�<r���A1���[5h����ʢEe��Gc1�DZoU���}����6��܏g�ö5r��y\VU���x�b��H>�
#rц�=�3;Ь��l���6�&�R"Բ��SD|`@�y�yv^�Җ1vyR�DϧJ�G��5�<���M*�SC.@P��].������V�X3v���s:J�t�fҷ`"݋[N�F���i�&'|��X��E��H,�"|L4fre����'.݊���!0p�а���6��k(Ѻ����M��:����\�Ftk�i#q��xÈ�
#�*Xɬ*6A�.��\LKb��3�T�SM�w4��>`'���v������*�ÓB7:� �U�ܧy��	a��e�$#h�L��&�<���qhd7�ew��'�n��f�U>u���n	�9v�8ʵ�I�68��h�݆�[�}�t��.�+�[a��XJ��o��o>k��~����s���,���ogk���¥�]+��Ië'n;��iB5P����S^�M]^d)���X��(fڣ@�۴�sQWFn��B�V������qk������]ֲP'm}�u6棢o2z�l��՛�O���&i�f']d7[�#�ýJ�;;�\-��2��0v��f��AV�&�'.dG�5b�}�Z<�.�tew>�y�H]n�TWH��61�"<{mgo��X�����9������t{xY�r��YNZ(޺��9�8���h�^� B�M�Ys(U�ե*Y���aŚ�kP�t۳y±�\yM�Tov�W,dqN��n�T��TZ�c��N��Ywy�Σ�Du�SVqއY
���r�9{d�A[ "� vP��k\vEG�&�y��w��UCL�m�Y���u��Ϯ��yP�P��V����^	��ZЂ1n__"b
:�0�	UaPs�u�ʖ�ӑ&1�~��V��L�9p�!΋Ż�V/�i�c�Lڷ��l��>l"��6&V732�u� Wޣ;��:��u��=|�����yw{v��H����d��ܦ��꾫:-;�)j�8t�Nt��^����TR
�y]T�%�o6bA-�Î��p�J�h���t衦�ce;��ɭmƆ�B�_Wls�%��D��ۓx��[ �)W+��u�ζ �8�e�luR�yL����n.�n
��X�,���į^E�s��2�k�]|^��9v�
�F�]�d*�aJ�)^��됥sW�w^uwg~"�{��(Ѿ���.ڱӺ�b��m#c����N��.���kE�gԮ�--�����L ��E��i���+�8diYm�݅����upv�Bby�]�7�ty׀!٩�͙y:���h�®U��V��1YM+*����9u�V;�Y��`�4�����MP�3.r����Ę���]� \M:GZ�o�j�!7-���@��!��E�q�&��);C'L�p��ӧt�j�wg;�/_}�y�N�-�F�|��**�ֆV�t1�/��N�+����5AF�+��Y��_S$)-H2�m�k"'�2㱲�%����hdM��F��2��fgn�Zl
�Y-��V�E���0�������k�/��T�Օ��;/��L
Ź�
 �G^m�n�^��1���S';6�;F�
i�4z�&mh�B�2;�T	����Kc��Kxp#Z-e�����^^m�!o���;|q5D���b��[J�ꤰ��"t֔����x�Iz���[Cw[eY45D9�G;��ٵt��he��M�h�ہ^ڈ��R����`Ǭ��P���F�Xuo$B��jѺ3�����2�Q��]hӽYg�J��if���f$�=r��-���}�Q]�l�^���v�:/�EgӨ8&�L{�t�mm�\�Ȟd���E$W� #˺d�~^�FCIN<�7�/s�E&��#��I�x8������Z2Ʒx�x�,�(����ժ�u�q-����yط㫣ȥ��$6�!��V^$�������]�wy���s��ة��CLP�6���W�Rvf�iq��9��W���fƉjܠ0���t� x���y�s}g2P��&*���6԰s+A�{^�	��)C��iF��FK�9ROz�D�M5�7"l�̀��J�yR��gg3�\71C��jo7����w��V��TPb'yqu��Z�q�f%Y��SI�P�
*��ss0f�+�QZ�ՅX�Ă*ZDf������YY���Fw��:J�ֲ*�bf��4�q
�(#1���YD@�L���f-�*�LvI\�B��*;$�%��1��I���J[&���m�#m��X�"��[��U0B��Y���
f�,�8�Q��;\C5eQEb�@�f5w��?��7/	���!�[�;*�).K�U-�<����K��[R��¥���?���}2�$�Z*�a�I�t;r��z��o�j�3�WC��.F�^���XZ�
�U��P��*Uozb�Gx�*yI���[��Vsq`O>�F<t�����S�eU�7X/Nn֙�
/�� f1�*�s�i�{�;�{Rχ��_ǽ���V|J��e�"����x��;t+�v��C��V5p}[���IonMyk�j{`�j�F�rT���Vk��]����{�"6 &ma�?y�50�������V���
������r�fv���D]�zX���=��s�1��;5{�L����Y�/k����жT�����v���0�"E@B)�^����k�,�M�M+�Xn�n���-�zl��{�6A9s���ipP!���6�
�kFx����Cˊ�z����	�ٲd�����1=�'zJ�F��h��|����3Ξ�)1��zf������p�5�P����v�$�7�J��.׷u��i�6���]/y���F�4Ut���}T�kإs�~ '��Ji���B�����!j=9�DyJ����m��,ۈ߸�}ѽK�|1��)���w��{�ĳ���
���~��cfm׈m�;�A��qCcuM����*��$N\ݐ�w�[;Z���D�8ϼrD�����4��Ƕ����g��m����xؚ��)�O��:���tl()��v�ư�H����ޡ�������lZ׼�v�&�b�/�<�0r�6�F,�w�v���맷���rN�"�o�ߵ�Tp��ս�R�c
�(��3�ڬ�Q��ԩ�P��S�f�8���!�U�1g��nE�u3Q�q��}|e��Iv����՝س�E�G>G8`�wPyGG:����f�ݐ+��!�\����C�0���;&�[S=��Q夭{P�̎{��,4��)̍��z^��$j�T����^���#Q�P
�=�2��[�����H�����wC��4���gx�Gҗ�z�H�Mb�:����6pgD�ib#�x4M�(����a9:���RG��!��2�v��z���������^�A�}��F�nc����}�ҽ���$p�1�zz�����iIxS���X[ڻ�X��}��%lC���!Ҽ���e�P+{!Cy�
>�}]����!�;;�,=��9s�>�(����_Ih�-�ʷ��Vr���ŕ�k��y���� w�*���x�Kf�De�%M����W�U��v{�΋�gO��ǟ���C��/Tɱԫ��c:3U�VFr�{ٝ��S%z_5 T�A�omY=u�ޖU���0��5�ȏ��6�5�]��&�(zA�{����򈚕�v(���Y�3���+%i.�y66z�ݏ	΁����i�7�
��+��7hv�7g�w.���`f��8��c0��.��y��2f6]�:���1�����Re�C�.r
a�#�����lE��<��������/m�[�E��Y�o�� x��C��c�{�
�byuna�"z�Ý��K����t]���{��6�f����-U�y��ʭɾ�0?,>���T��&�ܶ���X�q�u���8��|�S�|)��F�Q=��H�Tg�pG[C$ѣ��|~:_	[\�dqt, �J��L��֩��U�$���q���N��Q<��B��VKTЪ0�y�}}Fo���M^�
{�_-C��Q��Wmm#Y�mz�7���{����4�y� g��o��Z௰TX17��^,�wHxhF]E�y��{M�WZ(�|@�`���ǩ�=��$�gA7(Bw�������-�m*�!�%J�j���4��Ps�/��(*��֧��cR.���2��� k48�m�q/8f����A�-�
2f¹������;�A*�-�Mx/U�7\p2�F�(�����SMp���y%h�>��^+|9��JDu�mN��s�E���N�Oy�=X|��7���M��������ȸ�
d]�豙;ԗnU�����ݣ}#��8�|?�|��_�]��PS��-ɳ�൪�ԦM#5�$���,�b�0�T� i�$؝x����ۇ��b*I+%��Z��Uʉ���u�mIC�8�+I�Zk2��7d�wE����D�>�����v��'H����G0v�3rk��u2ۮR5y�I�ô�&ޱ�y�}��F֍��*��>Ƙ��:����+t�ϸf��|L�U27j)թn�BS(��;�x6��*�2�q�v�P�lc������#,]r�Ԁ�����:��]o+��.�Ʀۈ�W�OBȚ ��S���\+2���_�y�= ǳ�ߦ{�v��:�a�#`�+݈Um+�L����F�*b���;o���u��o�X3��ݵ�������L��Wj���!%����9w���s�V���v(�pĖ�Lu*�����Yl���1멨
1]�e��r
ӹB1N�r��-ٕ�=�4h�V0�81��ooD�Â!��ˣ4պΊ�̝/�(�v��6�e�$d�#�BPNK{�6ԓr"���
|�
��r��v_2\ۆ�i֨��w��e�:E����-Օ��(v�
+�4��Me��M��m���.6�ƣ����Xp㖕"��+*�m��a���J�l�+\I��]Z
�"�l°�$��v��jl��LUa�J�ea�NDL@�8��WVP�)@Ċ�URJ�d��j��B�E��CLuEFЗT��R�
�T+��ߵ��B�~����.��i�c
�]XR5����L~F.�5"`GW�B�oX0���IF-��d��Q}n�+��|>�y��O�GOW��_~N��P1��uz����]��"�AuK��i�봻v0�$|�yf�d��kي4��� P[{�A[4�:��.�LO.��c���E��ZݍΕ]�����d���G�޾Av�ҳ�|�m�'��g��R=63�~:�W��CR��Ux��9+&�o�z��T�H�t�'h;��VW!�v���벽�S�09��'VP�fC/x���}���$T�`�~�m1�@���_b�,�3�~$-�qZ=t��5q��l�옉�f��ܭ�/a�-+Ҝ0U�f߷1*������Ke�K��>�g(�!��:��r�J�Bi���<�۹܎X�[l)Gu�̓^I�~'�M�d��r��7G��TrM��x9M�mw���4�~ya�I�, u���^n��,y��ǻ/y=�$̋+�8�7f_z��XAi4�9�h��ZI���~��~��市��H�'�yg�j�Ad��a_!�,�^��л��y�<��恬y�z�.�s����ϛ=�f���Z��d�]*Ι���r8���3��)��?^�yz�<݃��a�{��������p���\u�O�������f��U�J�shg]8�5���O�{)F�����=ۋ�:�u��I6dၤ�Y ��� sύ��:�~$;d6xH
2CI���T�l&sH):a',��2�u��5��\�Ô���4�!6H��NX;Ӧû��:I6I�u�r�w�]���ӆp�4�n���$��vH]��Bv�鄝 f���!
Y�ˎ�2�\�Dc�����w��R����M���$�� �x����S��"<<$�{�O����|*@�ɤ:ByR(t�1�ڞL!����|���&���'hI8Bi ,	���CfMН�Bl����v߭�㮉v�oM�C�VM2I�L!�8@�h��]p��|���qH�݀n�vHo�$������O
�6C��m��.�uߎ�[�퀰3jvC5H�ë<2od������C*�]�ѿ9��ߎ�xCL!�6I!� r�xd�v�B�@�$� �	�@��[Ƴ�y��d�� t��I�N�9�B�Y<P� f����RA`r����ڎ��xǽ$2=�6���x#���6�!�g�ݙ�$/t��!�	޹�l�\x�Hu�&�鄨,�2Hp�M�t��p��Xe���ۮn���ل7I'L'$�!�$��	��I�&�	��^/'�w���#���^����ghb�oX��G�y߉��j��6*M��x��;�
G�<sל��wㄐݐP��<0��d�g6b��!�9@:d��8d�"M��:��u�^]�Y Vl��Bxd0ހ)��3��)�X��� �&2�^����I=$�2ABl�S)!���C�@�ÆS�jt�:`r�X<�<^:�v��p��$�d&��C���$ِ��$��,9d�w���|�\�Ѥ!�44ô�rɱ�$+$d�v��	��ā�!�!�l�wz�dC�,��6OCc����Q	7d��Bi<&�$.��~tu�����R uŐ�	�ԁ��T��r��wHI�B�lo�:׍�7Iސ� h�d;`,�@�����S�XMx��fH��s��ַ�~I�	Y�IX�8f���0�:I�N6�����n�
�8d��7��{�$:�Ā��fC�@�4�R�P�j�p��{��p��ﾈ���Ho,����Xwo�Y��m7��X��y~keL6�;���v�AX�7��������!9M�I��́�I6O)Փ�#�~0����ٝwHIf�����tJ=M����5�*]�Bc�\�"�ٞ̌��]��ĸ��Z<�v3sq�7PfPr64��,t���P�Ԭ���w6D?���]~�B���y��ͯy���^h(*iŞ�[�'*E�i~Ĳ����X�����o� Й�����l���g��w��~!��d󛣷lZ�����G_7������$�1�rV~-UՔd\����x�����:���p�~�<�XChrI9aN7�
�˺Kƚ&g{������zƏ�C�9��s^�}�u�������Y����^��ɿ{ֹO^�]�6�F�o^�#x5n{r/�[q�VRo{�Mk�EC�]���3ah�A���=�{�g�R����Q!�' ���� ���F2^�s{z��x{��WZ���.Q�f��M���{Ԉ�Ӛ�3�M����2��ʩ��]�3��@�>�O�_!�^t�w��G۹�����B���;���{�^��}v��7A�|wo\&"�o��՚���7|Q9F/=���:��#i��f��t���:���]��߬ޟi:q��	ps��X<���e�F�UE�W�E��qيA��ʰ���=o�x{�uS���*~��6�.��z��
��(�3}{9ß�}��}	�Y�A%򯩝��6y����� �t�yk�yW�'<��O
�o$��+��w�zbg��y�9��u����^Y����t��o�@�hc�&�
fb���DZ��nt;[����~'�|}M�O뉙��j�e51��0���H3EZ�P������ܝ��ga�N+r�s����R(� �|%����P���M���پ+}3Z.���s�7q��[.����Sؕ����g}���zcMJ�Ʈ�����\k��0�bХ彺��V�U2EZ��W��}ڵU��k�;��/���b�pRѐ	1�����jFG4+;'wN����tU�}º�f`�ۑ��{�c���pU��]\T9-�V�a�w���6n^g���q,ͯ����ˤ|hd�nf��b�D�q^�S���ٴ��ú^����#v��c��]�U�8��l��t���wr��ql�ك���*5kY��&�E�w�)(:n��	���D�Քu�DJ��%�U���N��u���,��o8�
��Z;�n�֪j�\�����0çz�,{S�,���25�F�l�?*�Ͻ��^rDL�I)���Em�79�E�B�!^���'ou�tQ"{F6e�����v�[� _��=���������QB�VB��U���q�:�i�`�!Xi�$�@�AA��Hf\�E�V�����d�VV�!A�TU����5�uJ��J�E*cVM[&(�HVG,�HQ��0IQ-��� �"�VLJ���A��Ŋ�E���Z�k
��"�#��`�LaF
�w�'�.7�S_�\=Jp�J<݅���J+���a���Q���z�*yR�����m������cn�8��s�j���O1o���A�����z+fSZ^&E�G@<_�?o�-�4�����HV��t�{��:�r��׳	�Γ�7 ��!��y��T�vݶwU��;�v���;���Xdfe�\r����*���\w�%����:��kN��4?$��wys�=�c�+mN�#�.(�������=� GOvE���n*goUI5�P#(V�����{3E=���37��̉��f:y��B��jN¢�� [�H=���}W�'�	�YW���zŎ����{��^m@�C���ÿ́��}o֨e�n��u�^\�h��]*����pst��[\M>[Z#�l�Y�)51� uJ�7�	?�`��Oq�4/um�=s��昕��o���(�埐F_@_`�� �G�/�C�G!�Qw���PA��Ϝ]]�yJ�ێ0Սc�U����ҫ�C+�ی���x!<�`�/*��q�
�.װ��FG^�C��f��ݽۊ�2��N�$Z����**z��V��˼��[<��/r�w�\���?ZDH�ڻ�1���H��L�b�`Q�n3���F����6���I1�(݂��Xb��V�9��f����  ��3�.�6n">멆DBv����<���Mea��'Ґ���y��]
��f���5��Yze��cѺҵ
�(������&U�QX�,f��v�r��(پ��A��7�҉��y
�������r��{����@�FH+���ޚ{ӂ��3|���<��t����s{���c��}[4���MQŷ�t���@q�j�F�q��x{�x��7��~PU��ݶf	���N���+�����N�����Ӌ�n���G�Y��aR�Vu���9Q���U�~k���`�0A�3���5�zґp�[㚸!Vx�h��zHG��ٮMb��\�|+��6�KVon'陖�����^��0�&>��O�\���1�݅B-���!�$n�7\�\=��e��-���/���s�31t��u�n���x{���Y�U0k:�9+7_fW�5�g�hw�j~Wɵs	G;��Acv:=����X�'f�F;������h�
���5վ2�q���:F�ׅ`y6mS9WV���Cr1;�L��O
������,c�.�q�^#>'k~��cB-{ǰ+�����F�w���<��޲�>�Ŝ-n�sZ��)j�� ʾ2I�������w{ȑ�̬���n�vp�g��ݿ�ߝf]W���E���h���3��j�g��g�a�����ko2"��)��cff� �kǉ�D���г a�FsV����8k�y�ҫ�5=��C}溞*etx�u�^����f8��{�q�h�>��F�u��X>K|Ժ��L�����]e�IN�mN���k^�grO��������z��lg�TA/QO������u-ղsAm\�6�s�����w���n��5�P�m�+M�S��a>���龯/:���9b��,n���gHV�kۥH͹\��Ѵ�pf����~0{�8_Tޝ������� 'jOE�4Q��Pm?_�4x<vP���y��d���5"�q�o�',��,*�1)IՅ#E��꯫��iNտ�+6dtY&Q���-:������<���V���~�<�~���\N��@Op�7���S@>����o|�"��-Q�p�u��>���9�O#��a��WS}�t3�3�v=8��:�M�}���ɬ�M$g.�*��`�cT���O�L�i�;� ��k�-=üq��1�Щ����=v�\W���$�2�׳9n�Ӻ�c�o[��9OWgȩ@�D�z]��1���y�naR�S��󪘻�sS�Ws��_t�E�9K!\n���M��Z� ^�E�/KK�Q����	�dD�4���ڞ�G�M�A��7�9�b�흟���}X4��b�c�fC�w2Ɗ�ݛ��Ч��y�o��8S�r��:���@m؟+J4*P�fܛW�MU�8�8Fksl�{���!A��t��b�ըR��E��_9�5B�Jr��Bf�j���j��$<iZ�ݏ���M�U������
r�ۘ�6ޛo	%U݇[@��.�''Y��ʖ[0ǚ�emjn!\dR�=棙�t�o2n�m�]
B����/�`��p�Qq�e�G.�9j�i	��!��]q퐉���3s��R\�F�[�9g��mt��3��*���6��qޥOnۨ�x��Oj�B�`.8t���9�=]�V�{��E5�p���{��� ����k�\���b��ź�D��Ƞ�y�p�ˤ��5}}�E�k��]H��t�P@�Y۴�]�	�{�xw�7a�K3D-K�軆i��]�.Et/�p�nd�u���FA���nq�|�̰Ž��\�Q���D��ɎF�nI��mpcgOd��7u�����v�X�͇��7i��� �Y�k
�,��ET��PR*�%�X�eeam�Z�bc�


�&+Z���T,��Ģ,���`�Ȍ��E@�Q�(��X���X@*�a�A`()ULM2b
�ETP,�Ȥ1,a�k�=���>1�ǳx��֥��\�������(�>Q��]#�{~U�]�fd��s3�S����x^7�={�gjI�M��ٿo��ӫ�8\�F�y��m���dm��y�]��5�=�<��Y΋�l������K�W�[4�`~嵻���Jq���o�r�1�p������*�[�U�F�]{��UA��/A�U��\u�HIYL��r=�#f��*�d(�kVI��ua9�x �g�]���9�#�{5ܴ%�j�LR�C���+�^�s�ђ�1E"K݅�^�z�_ymzb����&7Aa�A4?���{n*���>*w�tΘ�s�޺6^1<%��j��aQw���^4����(�'��}�F�3�N~(?Q�ѧ �O���8P>��\�nq���'}��X�)G�����a��\ ����������������R�_�~|�L��N,w��ݻ�0���ќ�*L"Zk$�}�U�2����(w�H��"{��mu�/5�^����~O|!�v����^��v�.ݤ/�k&�[��H�ս4,X�s��&��.@���+����E`�*��9�w�B�>@�ͫ�}4I�*���.�WI>;�k�*�����&�l�ƻ:�{������+�P��F���*���]vZ�֏Ŝ�95���8r�U�ͪHN.�ը[�ܺ��De�Jg�٧er ���g��o��g��#\W�h�	;ޚH�3�ف1幹��ԋҺ�G@u��ӄ,p`�pܮ��.�(���ZЌ@����B��˹ua�a]���`ޜ��u�q|f7�Q��>'fgL�,)|�p`���TV7���tOvU��]Tq�C�brR�����ҫ���G�p�6���P�&�	���ڭ��F�����O��l�vWrz��ɩ�΢b�>��Y�|2xN���&��@�q��Q���t�Y�_[��O���T�4c��);�k->�R�A����>�ל-P�J��vݍ+W�����_"�6ʝnk���`;mG6Hԓ��W�Oi�[��;ڻ��O���bI��e�5�tf$6/yz���^�J���(�<U[Zs(�E��n����V��Υ�Z�4��е�ߓ
���k.{���q���H����_e6-�=aq����ݓ��Q9]�g�<��y<��)9�l�l�y9�>��/uG�x�]1Y��0�|��vm��N�YU\u�h閶�c�S��{���{��.����+��ۻ4~�"9�]�r�)K�\$�Y~�G�������O�t}/g�0��Q�G�ٯe� �{��-n���9����{��O��#u0��˭�Z���;^�BH�(��"H��u��i��f�r}� B\x���6p���[��O���#Dt!�a�4�sWB`�X�C�=q�A�G�C!f�dcZu�09k21�z*�w���{��>C� �iU�\�ǉ�j�bSB,raj��rb�n�(���[����S��}��?R��!bfV~HnH{^��W����r�,�-Y�]��s�����ǈtP���$(Bf����hw ��4�6�O�Ѓ�"�SSG��(��]�i�� v��w<�'��2�" E�T�������*s"����qp�p�!�i����W���>|&B
��ӄ���T\b۳:�z��A+��d�`���j�5x����8�� Z
E!$�	!���֢U[ck]o�����?kp]4��qP*��ٴs�B�j턓�)W�H�r~�ª;����DZ�'dX���6�p�4l���oV�Q$B�iD�Vc�A���*�h���ϴ�K�@�D�4�Ӈ�S�ަt�AǨ�:}���!T�*[ފ�FN!��K�E��$��Ω���@6C6{��F�$�4@�C#M8ݙ4D�{`"�����H��6����*\���c*�@�,��_=���ݖAa�4)�D;C)�f	�IUݳ�� iDqS:G�P8��S�P�R���\<����^�i�v��;kZ˚�/f��1��{��3ݎA�|F�G�D��R��p���E;�D O,jH|�(J/,[ի�0h�:=m3C���K�	uW��G��q�#�;h24���U��d�C>��[�
��D�����#nz�h0d�p��A$ո���)�5,Aa����.�'ΐ��=�L-:I��ә~��	����AQJ��$Z��WU@�B`��qt��#�8jh��+w-�4F��a�C93��}�\���4��Q�7�kzYʖ3h�L�8������\�c�P�	B��vz(ۦ6">j��RWh�X-Iy�Zr^V+\�i��n��o6�*�Bt�jo`��Kd������+����툮��\�wM�R ���V�����r�����#�ܛ��G�3�ݻL�K3��C��й�W�8�to{��%#�G�8��.�m"�U�\H��RΠ�)v�Ԓ��S��h��+Ő\��"�I�F�ڈ���z{�U-����T���睛L�ʗN6�Ŷ�g�.�����An��ɓ�����ݵw�&i�Fe��n���Qz���uc⢅�bƶ-m�p�\m�q@I����Im��xJ̰�;��܍�(8���s��hNc]��p���6��X�;����k���IHrਵ�S�=�ϥ^����]r&�Ix���J)Q9$�����m�7�@�=�`�0�5/{>�^4�V<��xe���Y����/a��"�I^Ƞ�� �X�"ql����B)1��b35d�q�,��
B�����1ăl�
2,��@Z�D4Զ���
�Z�b0Ƣ�B�(fP�uI��
r�)3k�*�����]Xy�eV�}�[:�;�z�VͱJm��o _Mv{�!b�C d#�څ��j-G�3\M%FQUٲx�2t�9p#ܸ���"Hõ��f��:#qPA�4�Q��h���Ξ��=����6F("	���wm�0n���&5xllyIo9�u���تP�BrYg��p㎦^�,��F�<@�]hV!.��)M�s&�zG#�2Fj���0��0}J�R��"�����Ym���Y��a�s��iJLH�3j��8b\	���>��;4]ċ���'��˙�>79ϡ��41▙vn�����F�vUZR6[��H��w����c0���͓M|3\�uZ���[Bq>�@�<l���"�@UF��i�*�,��.Z��F�ș�����R�@�*#H��K(�fv�z����f���/
$�Y��������̼L��zH����2�N޻l��$���8F��}�	2De��'{���Q(��j�ax�U�ed�*�� \Li����C:cL��j��y�/���f}P�"�E]Z��p 7�������:����ay�A����^�^���롩�M�E�i��q�ET\�4�q�xx�U1^}'�'�	�u�8�e�!G]U�X`�>@���!*�G$�Fwjr�:�^� ���@p��}.�}-"U�i��qf�|�h(X`�"I>Zz��Ћ�*&�afz�����0����M�3dC^�H-6D^�e��f����݌""�>� ��	zF��Ⱥ�U{�e�(�F��K��(����Wq�}�E�I��C��$�cܼ�Ɋ<�9d��(���܁����0��%�3�}"��n���tW���ҕG'��3t8uAv�3��I�+x9�{�:�}��(q�=@�B��š�����_*�y���4�;V��	�@�WH�F�g	u�9���A�OD'��r�]�t�,�e	}�*c��A���W3[:�i��@����D��BL�4k�j�0�Cq#D/V�AQ�Ou����.D�����y_C<@�����y�l��dA�RF�6h�>\�Y�u�]��X|Α�ha�dh�;�77���o���(�E��@q�T��-��7�:����k}��Sn�-j��]+���q����md��sOe_ۼ߀Ne�#~���'�(Y�(�.��O碪c�q��օa�%�A� �?.~�U
��܎9�ARӧ�t�!��(ѨQ�;,���!���4�!ŝ#�/	�/���|4�A�'�8��'�ɋ�s`a^�Q��#���@�c�4���vہ&�d��C��HA�21O٭lE�:-iɘ,�0�$�b��/z���7
�5��Nj����A�9`�VB��-��/�5�!�Y���ofE���.�j���׋\\��ˠ������G�$2M��|����:͖+\��Y�QZ����ˣ��y$� ɣ�>���B�R��1��<�zf��da�ZbP�bV�էga�O�,��AN��4\�	<}������4��eI�q{�g���֚d�C�zZE�D�AQf2�Dt��f}�����݁	i�O�b�!��;M͜"B��`ip�E�֑r4�V[�E�A$!� ��Di��RO+���6Eb���>g��Gxgf](���8��k�Y�D^/Qh"8���^h\\�*
Q��9�l�|�+77��"K��]`���_��W�XC/���YR5z����~�N@�
�:t�A�#W���<��DAU,>�@���3���B;�:2q��En�4Q�BZ��#M�Z�藗��C>��"JH3�0���#j�cE��n�6G��ȓt�<ofH��Q�Ubwt�������R�dm���w�<M�I+Z��`RA0�&5�sܽ6�����q�E��RIުj��	(���Y��_!GL���tX2cr�v�i�0�턈K CVDJ�gŎ�f+(mi({�����[C����h
l�4mf:'2��y�󶘺x���c�/�����Bu|:��>�O� e"}����Ր��7S:p�D5��"�4F,�T/r������
$��W$E�n �y
��6b�ŵ2���Ir�d�!jӳ�6��$�����@p��� s "����O���&� �^h�8w�8A����r�*��}��	>��Dt�n L�Z_m\@����� �G�*c��r5���i�숻�E�7W��	|#�3k6$��d".�Y�$r��^�,��=1�vP%��&`�M��ʘ�ػ	+�?a&��Zz�i��x��q���{z��Wp@��_6r�<����~@N�l;����ܼ��U��æ�ZrDR��#)>�8�@�l#�G� �vQ6��FZ��q�"�]�a -Ŗ�9]Fg����:h��7K�E�"�U:�`���Bwb��"O���,�M�(i�0�a��8Ql� ���,������W��A��By3 �;�mv������"u��z�$	�]7���A��I�d6�F�Gb'��nb�r�q�[�MHsO+N杜M��D�s69�?�/:��c�>��M�P2�)#���#��$Yh�?>GTq>�(�<DD5�կ���!��е�q`�e�#Ȋ"�H3���|��0`�^��'�����o+ �DBBJH�p$�B�L���n�ܾ"���D�B"L5��5dH��b�,�y՞CH����<`���c�=9�"ϦW�Jp�G� A�L(�6j_o�����
�*H'Ӫ��%ۧ]��jl�T�^S��F��ir��y�t�#:��8}ځ:s� X���qq�Czrz�9�L������sK3�3 �h�vJ�^l�eV�� 6/]�8�xuJ�rl�J'u��*Mن�\�0�(*9�΁�(<������u�ͣ�`F�4mg,�KV,�;X.��K+f��{�@�D�Mr5�#HQ��]�)j�Ɂc�^,n�}.��o\�|1rCk���'�uAES�ٻ(Qa�Y%�)J��I6�n�ʻ�x���W1 ѓX_'RH�Y�U���.�.�m*Ze�אѾ�w�&rc6w�6�͸����>n�+b'��[Շ̏^����9�n�i�<%�ޥ��Y���/sW�����b�w5oJ�X�{Q @����w�}]C��Y���blZ8/J��or���0���Sh$9�t��$�f�;���	�V�W{���3l%��X�[�VE�qqR�7�gax�9�X
��G�nb�+w`�tFD�O��Ö��q��1��rII���c��ܒg�Y��+��観7��f���l�N��E0ıx���}�
��b
+�����%M�XbL��l���e�3.�fXj�IPƣ����0R��b2�E�Xf�puq)�c���B�j
��dA��ҥ ��d\nk
�呥��1��J���H��\�p`fQj]�Uq���0QY���`�f����o�����L�yk���n,,p�K�8��}5tui|�p��Nȏ���O!�ZNL��뛸t���$F* �8��{�/z'�j��s^�B͟i�@�D�&w%����C���Z}s��"Ȓ ��y��X�OC�GNi����e �6�=�8�E��Hr�G,$�Z$�u@�RX�%	jA񭁰����6|0��2TD�ꉁ�1	���6��2}��D�Ax��C��C��،�+�@"�>�3�daa'���jp%LL7{9�����[6�-�\�t��B����i�$'T�����U������p���V�ר�� ��z�N}�G����q�H>\EZp�����s�!�2,�&g�af�aE69S����X���Az�DCM�E��$G�hY�x�!r��$��2�>Ջg�t��5<p�(0Fb�DQ�쬂r������GR�<H�}dY�
��i)�2d�̖C>�x�:r��^#Bf:�F�Z�BgŬ1�Y� �0:-w�;�V�h� F( I�4�Cr01\jK�W�!噇"޽	� _ ؙ(I[5���%n��NX�KV+����;s�
�M�o��==�$�l�`�:`�EF��jDA��L
�wу���<��a�dq)�=��s�;n30i��@�Bm0Dg@�cT(�	ínU�<�E�������zH�����@�p&֘�e��[�drc;�[�򗨌$�`��������.������s^ j	�>�dm�6�0�
�d鑻V�:GbKê��E4E��$�$Y��.���4]�O����;:�^t
<d�AB�B�lA�����*v�ۍ� �ۂ �0x؇�{��{��T���ɟy��f���նƱq�x���q�sK�����0���Ǐ��Da�#^�VN������Դ�;�^��G&J�y�x ��$�ᔣ�q�2���*�cݾ�0�VF�G�z�I��șd��r�l�#O!�:��#�HCwo*w�h��&H�\h��#O�׸DM�ޘ�F�H�BN�0s��	��7W��q�M��!�E���Q(8�b�X�]W>��Q���$Ŧ@�T-�k{Q�;�#r����x��F��%�>36�%n�l���/c�1�ΥE�R�z�C�'"
�el��:���'?}��g����>�_H����#ƥy�G�^n�)�D���t�<i	 �R`���m���RxM@��NȨ
��YF� mtp���GA���>����	>z���9a��T+��a��O��"��Ƃ��@�v�U�����Ĉe��^�H�ȡ�TB�4R��y�f.6Q|�k�E�>�x��C�݄��f)3�>�X���dyRE������"��q�.8x��=(i�G#+��ğF����+�J���	�����˹X��ں+�,�p�v[���;�����8�}@�Ah��fFc3�=��A�ңQ��� ==]>�7'�̊3J�B��U�WG\蛳tYY}G�D�E�L��8�sv�&��&DB>�$��W�*�s���"�-- ͔|L��"�\�Ј\D�&����^��� �ch8w%�9Lz-��H�'�}�=����}�a�Bg q��ƅ7i�:��Qg�p�>�H��CW�Q	�������P#X��"�	y�#-Z@��F;�m�b�g�ً�B�^}u��הJ��'e�ϵ�q��q�[��35%|@�z!�+��+*�!��S��]�%V7��������4|4�*��H��^�0�ETҳb&>�:� i�C!z�_��!��Ӷ{v�։}��z��h+@�t�!`Zi����[�;�G��	<E�5� � �g*�V8�8�6t�-a�	QЩ؂n��ֽ���M
�:��a�A"�qm���T�"����:���(�[�!��}�$	�9�3Df�d����$Y�rb�VOg��	񼁸�ɲ��4�7S�����$�]/Y�YHa㶼6��/���u"������ͺ�6�+�Ʀ���m膦�Mk�@�Cu�z
���o��z:'�8|5��H|h�#�H#`���vE������#-z��Ϫ� ��oHڊ�0���^�f����<l�f���h�HD3g�Щ`H�/ ��St4+��q�-��Pg���CN"�C#�(�DSL�F���/d%.�Ϥ�/Y$y���8��3R*��FWL�,��E�4p� ����w�;�&=h*CN�F��2��p����\DL�#�i�L�,,�3��_L��g�o�p���6'��;K����f�BSښ������$�I����h�J�B�0z��+�&^"�l߰� T)!D@�%�#53�	�y;]�d�28�@�'ĉ4Yq"�g�#2�ETxid�8}ذ�c`s������0�WH�^R�F�,�.��Q]5M�d�ٰ8UT�(���{�R�ʠi�;52�
����&����]{Q�����b�A���N����m�l���4x���0�.�d2&6k��t3�da��'U}��"�ΞTb�~J=)>����*��f���A�Y�lb��۶�Vۀ�Cb�Z�;*�)#.O�W�~��Ԑ���(�5�=AVD�Q&j�}��H��8����c�"�z�k8�-͜�
�dR'# QӇ�:C,t�s�}4��M�$@��v�0�f��Y�����>ƀ�EqF�0Db�}��J]��Ɏ>�\�(��)!g�{���B4Dr�XDB�h�L.�*	�s���@�DmP V��
6|'���c�:�
∐�&W���!<�DJ�5)��n��/�ɡ���5�E�6j��q�,��ua��-"��`NdBE���vg� nYv���,�XT1���9dt� 9VyD�z��ʙ�#��7�lR񹸜N��S{�zE�H��E�bZ�Z5
�U��sYbl���ΩE) sb��"��l���Du��I�H�s:���X�1_ ���e=�B�,֟�82jG0�����g2���=i���y��Kׂ�Ҙth �[=`���h3[a��H��Q7�V�ڼ<O�w�%J�6�	������������;��K�*��3x�����F5����W�h*�-�@�8s�v|�JUv�K��ށn�H1�������J�U��^�=
bD�j�w�o�GZ��P��q�p��u��U��>yxo$d�S������#Fb�B��6k�u+�JT�5isՔf�9+�3ZA]ʵ���/B�m �(J�'��48L\:Q��ڋz �uԚ5!�O$�=�.���桅�ԍ�rD"e�qD�?��\����Z�Rn5�:\Ṣ�8"2��>��ʙ��P�ΣJݛJ��maZ���(���bs1f$��gYf�����[��ڷ)�qkq�XZ�3Z�4�f`��T�\l� ����rd�qZ�i��nc��&���h�\��\ˊݩL�m���\\�����#i\U�ܸ�6���͝9��E-�&�n]զ5�h�aEt�ŭm�ع���6�UO-^���w�s�E��ZD�S������ﾋ���$����>(��9#8GQoN�>�6G�q!����Ad�z�,��\�`�Vh�#Z�!�Ϭ��#l\���������t����r=DQ��2�D�/	$��.� �>�C�s�]���Af�z�8GX<G9�rOemtV���4�Y��V�p�� ���j���R�	�$	(bt�@��M:�h��Qg�����B��v����#-z�	�i�^���=}]R���e�wY�d�P��}@jNsDL0��w�sa���r��j<z�钳����諭�=���r���{G8#�������ǆ�z�rq^��k"o�n	Ķ���؋�b5�N|���o���/�h�\2��=��m�-i~�u�6G�O�)���n�"{����=��>*-^]Y���Z��X�׷�3ۉ�bMgwƽ�'kjg���j>^��d�Z�zՋ����t�tn�"��]E�h�2���]w�i���2�!pjb�����9�UWپ�yo�_���"��R.~�X������S�Z�x�D�kRS�e{�<ʗ�ǫ�`�y�3vHO�#��Y�^��X4�iQ���=5,�O�x��5~NYB?)�KSK������n��}�6g����X��R��=%Pmf�Ƀtt�nL#�#Q����I��Ӕ�MA]`p�̼������Qz�Ex�:#@u��8䟫پY�;=�G����X`�6j�>���o��]�O"p��%�Օ������	�m>��]�u�
:���jݬ�ϴ�n`��V#�ו�<)�m0�[���2�q"��yz&r����x�]��\�b��K���T��J#7X��V�����1a���O�g�v�C��ѕ��:�_�|F���If���`��c/�V�YR0��������'>Yt/��r�0c�v��z�(n���]0��t�L�Y�{�����t�+Ş>�=�!.�IOk����E�Ae���x/�����;�ŉ�֊ڣd�tR��rx�Q[FY;��[�y���"�>���;v�g����`��P��{s}�;kW-Ӷ��p��!�?]{�O���5;n��Zi�h5Il�u���t�S�ǭ��x�U7��N�}���y��xyj�]k�dRr��B���OLM4(D�{��s���1��k�Ǣ�����]!�[Nʤ���@6�z]�瞏�.M��əN̬����:�{�ٰ�s��0�QyRj7�}�>]� !>��خ�[�	]v�Cg����g���TЌ�`�Ģ�rJ�K��#�f]t�ums�b}wx�(	��}
4���n�	�۟��ꯧ��]���O�T�e��"#s~[P��v�OW^)��{���{Y���v3�	y��P�Q��w��	��l*Q�������

�6��Է2��6���������*�V�8τr��z�y^��Ъ;�_vVL��:�V���=��Ҋ��]o7����"+�!�n��ʯ#��uj-'�ǜ��Mk��21�ں��m�����GOv����u�\�4�Rc�����眸J۽t�=�Gu�7ŃH�Q�h��Ӟ��n�f��v7_�՚�'��s���XkS���Tӧ@Q�:��)D҇�l`�>��� ���7�F�J�x�7��IߊM�y��=���RM*������xr�P��$��!{��7z�^�}�C|���TV��(>�k5��փUaMk׭����������}���F������{�3�z��O�3�;��2�P�N;1�n"��}2t�G���/p����=������],]��|h,��=Ѥ���A��!GD}�n`�:��@�{��D��ȹ�j�$�w��Dm�w�׶�ţɲC��� ��k2���#_��vX�Ӵ�mJ]on�8�xᓮޗ@ap�@X¥VQ'����7�X�;��=V@�9[/�밵H�Ww+4E�N���]���w�}�������t\����a���z*��!zj!��/q�+�]`���F�x8�V�&T�5�^xhO�̀�s]m2����'��N���.����ߺ*j����y���p%{�7c���߅����]��������^]n��,EK]�n�����<EЍ��Vw���ifX���ʑ:&��Pm^A+S*W��1��6 �i�Jк�4���W]ը@����X@C���$7�� ]��ŦܶD�.DtZ-(g.]ݵ����������͓�-�z����t�w]���A���O��]=m������X7y���7ȅ�x�}���b�h�6�ݴ�̲�$lS�b�=;_"�5c��%�2���mm���s��Jb�����	��(�[v� E���,��Z��V�T��>J�u�/I�o�H����/V�9hьDaIS�V�m�������I��<P�vZ�a�eV��Qu�_%�D���r�⺏��A}��W����m񠾙�u��[�^7L�L��)PK��QYk%G�'q���c����Y1�JmC����҃��N�%
,c�1`f�4΁���cx`��%.F�h�#��2[�7*)%�諗pM�2��.�
��WƥMݭ˼e*�aݮ��!Z���
`�6��բ�5�5GZњG
-E�er��S)�"���h�鮚:q�MH�բ��ʎ���ƍ�5tf9��˙M"��5�h�4�&�6Ec�L�ە��\35�ɬ��ʕ̮���a����-�R��%mr����
�m��ͮ�h�\��Øg�E���N��*b�j�@�Q�}_U}~�!������Ì�-Wm�p���u������y'Gj�&O���Y�oW��O_�0����k�=>C�(���g�(�H��$q����{z�{�1[���a�b�`S+;�n4��x�7��j����}�j���LR��}=´����L%u�p/���
B��H�&�͘�Z����Ճ��	"D�$M�5��ԡ��f7�����{B�E�V�ף����d]�F~��X�k׽0��2:Lm�z| 3u�8w1D&�d�MkP�]��3ă:ܚ>��d	X/��&��h��f����R�W{d�L���륜�����-��o(�Wϫ��f[���1���G� >p����e��=��;���Fc��0��B���؝�yk}Ξ���{@�7�L-T��E�[bN��	��r��:ϛ��)x_�KE=����7	���Sã�[O-E)~)'ٗy5	�
U�5o�J�͕>s��RS�R�̋��b�Sn��8�񦎬7"f��L�����P��P����"�~�+0���{ɞ�{B���TJ��k������}�r�r������Ҭc��p����%ð���[����ֆ�O` �*8ܕ6t��*��ֈ%���N=x���
��<Y]��S�/i�˳��`������rE$���������epý
�4@}���2x�]؎�ዪ��xWl_��Ў!7����׼���a���zLP�
��q 6ϗ��{i��g���-�jxV3�~�(�o���Z&W1&t� ��q�+�s]H$�OXa�*P��Iܻ�.u�H�N\����z��
&�v���{��]=���kã)�RȮ��{��ʤ��7�r�͞}vzhW��kF���e?um����dU��6�[�~/���G{-%\�؝�h��b�z��4r����ЃyG	�ty��6��/�3����gi�Ǳ�%���20K|��PC_�,�8Ɋs�f�-հ�"�9�=����f){�� ���Ux�R92f�C�9��8/�g|o��ߖ��6ϼ1���cüI��U�z�>��י�T��9y�ɫVW���*m0�[Wc��.�N{��$߷���ݫ�����M�_x�,��=S�UBy�%���"��Y�m�ѽ��x�<�Y��_u�͎��F�0Ow���v�؝��vo�j�~Fo��uu�۲f�KN�R�"7����(���T��c�B�xpk}}�9��ʘ���*�wӼ�s�M���{.l��{�8�{Վ�n_5�4��lr-G��������9H�N�9g�LV�Ls7��#xb��l��r�ݜ{7A��#�q%�6h{�J�����.)OQu��N��o��jF���{Ε<N����q��x�պ}U�P=�f����뾞�7�j��0o_[D:&_����V7�+����Ғ3$���]R5@���y��F}yט���"4
w�E��!��*.���?[�m�9W
L�L�K���s������aEdvH�{����Z��Wt��>Ts��������~�2n�Y���_BA�+�f�p�}	:j��/=�(���j��,V�ײ.���Z>�ԯs��_w��n5K��7W�`�Y��ӂ�V��֒��Ե�S[�e���9Y�6����c�3�ig�Q��kg�QVh���m����4���#�T;�Ӕ��q�ɭ��pŅ͠~��^*�h}�^����<y�U�徙I�&�\�K�U6�w��{���sF��pk�7Q�ot��ս8���Ly%u�7�lPΎ�ŗ]ݘ��
����};��֧�Ҋi���/��(��]ٻ���Ӣ&�CVvi:7�M�gR鏶2N��^�'nwD#�֎����Ӹ�[�/3g�h{�n�����']�k��q��8�ծ��=;�Ɋ=��Z��~�>�&�A�����ga���|Ms���ئ~��wS�s<i�T��6yJ��C�/z�hLT��3t�ӻ���3��U���t��V��%�Ǟ߰���u��2&#��m꽅f�g�ެh�e�GY�H����p:I�\m��WR�;7?���\]�&�s��!g����;���|%'�@^��n�&k+PE->Z���i�=0�5����Z���l'�tջy5��-��,U�ly��c����f�w��P���VFs:x�Rj�������ã.�����[t�0�OO�G6�S�*�aQ̖D���a���ob|nA�
U���r�Iv�˔ٔ�5s���!�^Pσ�k��P��uƮ����e�.����j]��[۶�$dml��m-������hea�	��:᫧[��oU��+7�M��IQ
o��:�R�)wt��٫&斣��Gvaݣ�,�ef��d��P��.d�a�[5�^�V�Q�җ��9-���ǟ6�u��������\��k�A^���ҳA��f��)mCnFJ�9!
3%�cq��^�ޙzi:]�G��S5�g:9�6��=i�J�\o�󶜮]`u���Z�0Q[Jխ��ֵ-cz�:�����U��--R�5�]0���h���Q�K*�[v˵���0D�ҷ-2�ūn\X�P�3K6ɘU�i�Y�r��Z�ۉL��r�ِwS��x�t�M�yhnEV�Y7���䑹�6C�W��\�{+<~\�����_vĢ��3{�<�sg���;�v�H��٫�=Ӷo�l	�Χ�NѼS�b,�>�����7�CEoynFk5��	�%���ݙ�ս>��>��V���b�����&&N�Ț!S�4-s��˅���Ȳ���WVG�Ƀ�f�S*=�g�dR�}k������V7\�o2����筰�K��B��˺$c�{4��/����loGf���9ޮ��;3��Xs ���C��e��1��w�D��[��aXV��0���>��P�l�S��YK�|��n�n�G���Qwޮ�7���K�u�hXs9���-�<x��t��}�w���
Ǳ�X�D�'��I��e��p~�	�ԅk*�d����u��۽6&z�MR�B잷�[��k5EmU�#e�3�������3�%��f�\�P9�ra�y��]���e�og�U�y���	���WGm�1R5�8��g�>� б*;��2�(ϵ6wq�@R��QH5;Y~n':���%o�G�Y���W7�b3��ׂpN�<��b��=ܩ�d-���SkA�,
6��������g�nk�r�Ճ����j`�L����c��v�c�4�5|#j9*l�x������C��f�E�E�P*Q1��7�,�Zc��펷b�Ll�6�c-M�ȭ�T0��+Fp[�#e�-b36�(48uF�u�-��
��{��#�G(�����
f���	UJ�� �^���b���{%�{h{��Ő��|��t��,珈޲�9�ʧ��|��5�r������L�ӄ�>:::�E��W���)��s۳�ns��b���s�I<�o#MǐN�
�x���<������Ig�ʦ�9佊�O����~o}��>�ݙ}��U��{��Xu���׉���ϩ) ���������/���ϙ�q��֟I��c�*��u��z�Ǘ���0���P��V��Iz�<%{�u�W��j	Q"`������-Fr���t4CF��o�}Zgx�z�C����L'9��$�z\&Lൕk����`�b��|6���> ����N/&F�@w`:��]�n��q���L��{c��=r)s�Λ���8�G½���^yf�w��PQU�2 ����8�`]義��=\pg$����J��cTW~>s����^v=�Y<$���N�qZ(^�@��"��)gL�2��=�*��f���lr�-,n����� �pq�$�7��g�;t���*E��Ջܩ�����qX���j����0�)뱄�����x�|��*��&����)��g��������g(R+�0ؙ������ŝ�2L<j�w�Xx������ve7�ahU8pZ��|O��D�{,��G��/N�f8��ߖ�M�طdR�R��K��:u'yРͥ�BR"�%)���h�6`���
a���w��Mm�;2�ntr�Õ��S������O��e*�/ELWS�L{��� �4?G�ع�{j�[A`�^S2��y��3$�ܧ�3����c��ͥ�7��ҵ~��Q���Z�u�OC~�zYdp|X���Z�;�ov�|ai���<�̾��Uw㚝�O���G9����6�F�ťE;<�.����6�
ww>�j�drT�.�;d)���G�v>���q��g}�YC��>��u<����҉�{xU�8��u��[�z���[C���|�+s���>Mm�k�D�h����/Z��>#���������=���y���#�uװ�񃽜a/'�X�#kΎe{�d��¬j�ں�e�1}�%5&b*�H;B�d��o6z��>xξ���6�����؄X�(n2�rW��c2rOD1�#(����Ⲹ8����nGs��T��T���
���i�*�vlu���vM��U:�=j�������yy�3]n�v�6g�ܫX�6=�d^Ç4��iq�+��;7R��K���E�X�<�[���BkXNE�����N�*�c��P��b��e�Dcݦ�����:nc�wh��t�[\����_e�ɐ;���E�Y}j�%i�X+s[�R�[{N�!g��B�V�sl�}`�7�rԋ����)y�@L�]�)�)�����b�E����}kp��a?`�w,	
���ݽ԰]s�r]�u�Ec��R�o�Ȧ>
��|�u{}��k.����"���p��@4�#̮rn�q����L�'R��M$���9��ݐz��;�|�NǏ&#��dJj�&�ЖAS$ziL2\�l�ff�n���y8�&5�bކ�P���e#n�$\��$n�/Fr��R�.����*I���U�=3n�;zfT����	A�H��-�e�'S��tk���u���u���Ն7($	3�V���ܮuҗ��� KW�,���̸8ة�����뺔,��)�݃���i�U���S*��0�{�0Y���D�1�#���M��I�F�	�$��=0`���p���Mx1 E����nQL��k���s�f�0��_rUw�L��U�4�̷(T��f#�U��۳��m�M�f�]�1m*��
��ՐҳV�vk���
��`"2�J���Teui�����n�I�c�����i��(���Lh�U�����GT��V�f9�!���Q��"�AE+F*2����II$�RD�:/n��'��2��n��ZJd��uaIN^M����U|3�N�@}�y��>�F�&�!b�ǥ��<.yvx��@Q�*މ�;l�{���;ĎØ\��Ѡ�����+d�<2j�%�ݐ'=y�9���b0�yl�7�]oP�bx*-=�ݠ�˲:�l7-x{<�=����"�{V_���zr�+�&�x��G�jW;�u���|.��}�Kv��5��y��Q�P��� ��q��;�870����i\�L�*�����J�3��,[WxW��v��Ϯ-9��%G Y�l�V��KP�|�*yӒ'o�iZ^���l�ׯU2�-�����R��'�U�^���,w�*';���&�v�������-)K�0ײt�<v;ݾ�#=}�<��VL�*8�ӎ�̱�mu�?ɯiw��F�X��)jL�� �U7���bG�ex<�|���Q���w���Tp��:o&xye#�n�m��(��ki���yhy��P��([�~�qm���[��ػ��@�c��wް��)���ˇb�@�/��T�'���swV���\g1�Q,Jˇa�ٴ!�>R�14�>�|-JУ}M���u�Xy�&L8�����Ӳ�=�T&�D��%�U�H䩻!���������o���$O�uԎwo��x���Ex�/���h��gG�[�ֺ������[�oB��y��cǏ�\�G�º"C����w��V�+�Ӆ�Ko�>�[���[A+��a��u��MP^rD]�c�Z����t�w��7��w3m������u�}�ƒ���ݦ��].pe�9���[l)GvH�q�|_]"��y�l�^���~>�_�Ȫ���Г�Y�RN��v]Bv�*xΰ<�c�/Q8�Q�h�xA�e
�(�6��<�V��ωF�:2�'H�5�����{B��]��h����1��Ѿe�O�ѐC��q���^@"va]��$j�X��oP�^Q�~û=�T��<$�*rL�4>��C�E�����obIV���*H⒦�/c��K��k#|n:���YB�\�>R�>p���d��z�^�{M]-���پŵ}Y���Gv_ݼ��'eE�(�lg:�z�����Y�a���M��6���΋Z����wͭ��e�{����{��1#~���q\�H0�<vjyz��sSĢ��K����_��zq�����vl>K��Ԩu�r�F_,�q�7��zk4��r��z{���*�+���G��C=�s_�y�����"V��Be���Y�v��G���c9-CiK97tS�xTwn]�V/;z�1����D7�[y�=��j�T�y��(;=�w��K>�8�r�43�9'��B+;*]�!�[�SFf#��H֞�ٵ��o��9iE�{�mH1���ƗbS�*mvS���;��JU�R4[��@��V�T�}���g�����4�,���g9�O���WY5������:�1�5$J\���#�I���}W�$]�w�צZg��N�f�^T������4�wn���+�ƸR��v�np����wb���oU�E�]�.2���RxpI�qд]�u�R��V6:�8'����Y��5����:T4�g3�I�a3*�H�lݐ�g�l�P~YP���;�ތ8��P>���GR�bn�6���v�jJ�r�~��衳J�V�S�r�\��n��A��W��N�%��Rl�Vg�oݛ��v��,�3����cy�]Yw��m�K@ߚ��o����U��eV��ïY�P�%O��>��[�ǐ�˻
�4W���ŗ��مe]�����lS4�'u�ݼ�����C\2�$�7�z�Yb�	��/3��X������i�"�����9�u�hd���s���	�;=S��]G|�YG3��k�V��U���;Բ�-S�ւ�k���>����$��v�	��P��H������PY[(��N�G�^�T����s����kgFsή��'�{��$��"�������?6IHA�O��$�$!����I!	x��?H��<~P�`�,32g7sP,4�Xz������:K$�M!$$��HHd$"O陡f�h7�&兂oaHy �2ʐ��A�Q��W΄6&Ĳ_��HBBh�|�N����}�����!�������DL����{t!��H�4XrjC���<p�g��0���u�o q�J���q�A�r��?�!��|���>u` �q �$$!��I!!�!�$L>0����̇�C��$�{��$?M�?��?�Oy���6��<��>|���!�$?�2�����H`p�����O�4$8������r$��Sc!��K~�7�0���>h|�������V�M�1~BO�d����ձgq�n��c�����HBB'��>�PvU�:ܖaC`�)�!p06���<M��w=^D�sc��$���=Rnq@��n2���ǡ��OO�S�6�ŏ��Yԛ�?ZOl���='���������O���y�o����#)BB|�dgf���7>2̓����74����)�셐�����~������.�zI�'���@�A��$��������C��|�!	z�{�F>���x~��i99���0D� (����B��&���`��IHC���'�B	�;���4��C]OĔ<�I���ؔy�@?"M�< 	!�p=x�,I��>�H��9'�^��dؠlN d��{Cy6!�ˣ�'do��(p<HN��d2I��ϲLd��S�6����/��A����`}G��i�H{d=Đ���H�A�D='�� �#'�~�)?�<��"����'�T��>P{$�5H� �0}�'��>3�����Ϻ�g�9&���
IHC�|�޳�� E��-, |�����IHB��l�0y�p�~�t��?l>�rz�<��2g��rn1�2~���C!1�P�bCo��|Ϸ��Ã�!���?�|����!�:;z���y�IHC=��Oi&��o�3��#��~�0�O��Q=A�<�!=G����y�߽�rlCR�M������HHC�B ����>�d�H�?��#�u�@���> {��OH2nM�nO�xm�w�$�$6�>́��ln���?�d����Bx��O���"�(Hhz9o�