BZh91AY&SY����߀`qc���"� ����bH��              �C�d���-"%%e�D	(�4�((kUT%Jj�-(j��)* T ���&m*�J�JF�%TURFVh^ڮ�$��"�V�P�"U(P
�Sk��m�E �"��
$%U@�Z���Z�d ͭ��� =N����z5Ъ��]i&��rZ��À�T��R���lp�v�*�f�'Av�e�ـIT�� �)������((�����ͥ��E w�Ӻ�ݺ��Q�s��Y��s��m�s�Ui����ٶ�ei-"ʻ�ˋr6;;4�
�ws�u��ki�W��=v�L�cJH(i�V�4�$y��R����t��)<���׮��WRޞ@
\z��)Dt;������5�R�W�ĕR���l��UH���c���P�5e����m�`�7����T��X9@�u�i+bR��`-S�ҕ%(yk���)D�i��o{�Uz�n^{U{{g@��<�z��]ݛy7��
Smo���_m�z�;��^ڪT�9���%B��F�<P�h��缢�/w4�"]�Q�
UT��
R�����E]j�����P�Ew����YQF��y�ҩ%T���������Ю�R�Ǭ��j��̸^��)Uޫ{�v�@
�{��J�5��'u"@�*�ŉ$m�M�ERT���>P��2_=��UU{ k��{�ؤ%W�gO<:U=���G��*�k��*�H���w�=OB�u[׫�iUOuW=x��Z������f{U)�6�l"��JR�w}�BJjǎ�v��\�5A�P�]޵@v¶���v�iF�F�;IÀ������;/p )�2 pEJ��储�������P o{:>�P-���S�8wuKqsZ u�{ޞ�����8��wl� ݔHq�)U@%��)lb7�*U)@� c}� 4�ܧ 6�uX�t'.�(�.��P s�#�P*�+��K �ra�@��*P@.����!K��J ���/�5� �;��҃]�8 t]�^�t ��P 4�: �:��*�0�'Y�PD�h@�JR�=�o�� �Wq-��p�����
���Յ4:��p�;�w��<��M��         S eJ��      O!�IRT�     bS�d�J   b  S�I*R&��=A� 14`�)*���  �    !�Ԥ����#I�!�hh�4zG�H������Ѫ������WM�0�2���x�d���>xy��Y���󿟰
 ��w��*�
� �(���E_�"�*�Pt	������1S�j�����U_�t"�*�`�����������/?�����1�,�[�1�c�m�����x����3�cc�1�cݶ61�8�1��c�61��c��lc�1�c�����3�c�18��1�c�q�lc��c�1��g���zl`�1�c�1��c�c�0g�g1�cd�1�a�;l`�N�e`0cc*cc
x���������Ș�̸�8�8�����Ș�����+�����D����T��P�^�d``^�G��D�D��1�q�q�1�1���T�(c"c c"c"c �
c(c�SC�D���D�D�<aLeN22&2&2&2&2�0�0���)�)�)���������)�/l0�0�L)���c*�*�)�c"q�1�q�1�q�1�q�q�ddLaLdaLa\eeq����SC�E�Q���@��D�I����D�����D�P��1�1�:aSSS`fA�Q��P��T�@��W��Ș��0&0�0�0�2&0��*q��D�Q�� ���d1�1�q�q�1�1�1�1�q�1���P�@�1�q�1�1�1�1�1�aq�1�1�1��Q��@�@�P�P�@�a	�1�1�1�1�1�1�1�aq�1�1�1�q�1�1�1�1�:`��D�A�q�q�1�q�1�1��B`LeeLdLdL`LdLdLaL`zd1�1�1�;`LaLe`Laee1��SCC�LaLa�C\`LdLe`dd�\e`LedLeLae`La�1�1�1�;aeL`L`L`Lg�A�D�"c
c �c�!�	�)��T�A��D���Rad\`\aa`da&�U���D1�dLd& 1�q�q�\dC@� xʁ��L�2��c
�(��2&2	�U�A1�La�\aSD�;`SdLa �� 1�Ba\e\dSP�U��Y�q�q�q�q�q�<gW�"c ʸ�2�020/GG@��W �*��¸�t���8�8�l#� c �(ݲ�0��� � �0�2��&0!���*�(ȸ�t�0.2���2� ��&2!� c ʸ��#0��+� c��2�GGY�q�q�L�E�1�q��fA���1�q�q�q��CP�E�U��i��1�`�q�i��q�`�|q��Lg�Lg�`�8�2c60c3����ǎ3��ǌc8���q�g�c8���`�gǧ�3�c=��c8�1�c&1�3��ǉ�c&3�8�1�0c8��8��g1�g<`ƙ�Lg�1��&�`�q�ǁ�c&3��0cx�0q�1�`��d�N��1�c��q���1�c�q��c�<1�g�c�q��li���q�g��1�cƜxc�1�c�1�c8���8�1���1��3�c�1���1��c8�1�����q�lg�c8�1��8�18��q�c�q�c�1���1���1���ݶ1�t�1�c�1��N<1�c�1�c�1�q�1�c8�1�c�1�cv��1��1�c�1�c�63�c����=�1�g�1�cǷ�1�t�3�c861�1�c8�3��c�g�1�lc�1�|xcg��1�c�1�zxc�1�c�3�c�c8�0c�1�N<q�g�q�g�1�llc�q�c�1�cǏ1�c�<c�lc���<{xc=61�c�4�1��8�1�<��1�c�1�c�q�|y��lc�q�c<1�g�<c1�lc�c��1�lbc��1�c�1��n��:lc�q�lc<1��c�q�lg��1�c�>`�9;����8_���%��c��b��KY
�p�[�pY�M����l^Mn����76,vX�w%7]��4�.by[{�Qf�����f^����isk/�\�M㻰���˓}wnG��1\@��(X"��T���7f0�YOU�&��wBmJ<�x����e6�fC3l*���7��,��6 �N��q[��Mxa
Z�ͪ{"�� 7����/�a��v\'!�F��ţf���@V�ņ�� ��H�+6�m9lGn%m7z,0�ǹt]˸�v��ҞT�N��%�<�{q�,�N���,s�UڥXi�rU��N�nL�;6uָ�����Z��gz����y�uFꈑ�7�i���|6{[�.���^Ҡ/}�����2�۰CKqi�yzcd���x��0�.�J�B��`X,`��I���!;��	)F�����c��nCr��D �Ka;vv��8�{��)gC����HЭê��%���T`uN��mҳ�m]]�j^7z��Y��{���z�^��e�$
nB<���l�oE����v�d�ʡQ��]��UK�tC�0N���=u/Q-�:�L[�}p��oq(�A�֗���^9ɞ���z��
���勚�kjf�b֚^��=�y6�G�PPm��]c��S�TO�Ԩܻ�:똇V5kS�̔��n�R;����F�4h��+:�q`��`�;R ��m�eB�x�nkQ����Ⲟ�`ǯ!�@{#�p��F�-c������k%)R&�[�d�I=�͝n���N�d
����XR[u���с��~v���iU� ������p��@h��إ���
y��W��ɱ�fcW�h�с(q�N0�!��H����0�3�U��/����[���]O�i�4�٭6j����٩���ӏi]�ux���B
`��;�P8+EՍF[�B���DK6��<��^�I��j�s�w%e��7Wl�y�暆����U0���96��X�e�0͹�"36��f<�$W�gKT� ��r��vojdU�6bV<Ri�p�`��;;J�;��e޵up��i,��Of�]䠂�coujڱ��u��`	�aGkC[RU3 �2�Z�cH�jf�ړM+0J�9�Kw1�I���.��JԼ���%lQ���Q(��S2�7Y�!se�K�/(���y�~Lɔ(	���-<� ���,x� P�܏ �H�ٛyP����c�%�:�H�"�L��
���>��yl퉗�C��E����uER�V��v����j �-<@�Z�H�[�y`6�D��}�U9��T�2�:B ѹɮ���D�����@�K+&A� ����0�74Ap[��)1,��{CR�T3�bS��\��
���5�uW6�q��L�$�dh�V�m���r���D��EcvXNQɷV�KJJ5D���`�,���:��v^PuAm�.��j��j�}õ*�α�Q��ien�V��H;�۪l�e­+�h�[�T��#:�-%�e��M̕nɱPh(��Eƫ
dL����u���4�d���	t��Fm]��,˒��N��F��qfSr�ͨ���������eڼŶ�*��Lc
������ki�[�v�P��b�
�C/{�Y���OwYZ�/XPU�b��(v����4�1�\��R���j9M2`S`�G2V&nTh��v�ܹ��j��hDn�*ZX�y�U��B��i�Z�P�)�F�[t���nlUY/07��M�+��5��B�GC�WR^��"��.�@�"s@KF��5�kV���#-�N�!cGVݙ�&m͌Ս�{��WdY�V2��̈́�J#ڧw3x�ݝ˲$��r�M�/�ɒK@�9���ͺӁ�D�����Tɹsh�۰/R�2��AA:�{yE����͛x��[ �nź���q�7�IDKy���%��صM�e�7��t6���W*��N��f��G)�Q�Ƅ8�wY/j�U�ᵼ	I�������b8���^�6=͇W�ƍ"S��rit��u.hB��yP�,k�lOa�ڊ���&1Wpc�V",=��
e�"�ȷUɔ��
�4ֱU�� "�v`!m��Tn���� n<�aF��x�ݽ ��Jm-�E���r��EVS#ǁ���M;�f��V�WҲ%c^���
n���Sjl("���˛�kI/CbìB*�V�ݑG�I-����y��yJ�����HƑ���
��-^e*�/L�cm�bʫVh�ܬ��ō^�uYQ��zT������+�SH�Z��THҧ%J�j·M�WQ��J�(�27��������m-��y0ށx �M��YJ��e�w�V`ڙz�\�FFN��D�%<e�BQ���V֚�뺽��
�7��@���`W�/NyMY�i��P2-FofټQ�R���-�̰�f��6�l�<E�ѭ꠯c��m,ܖ��wa�����KӦm[�H@v��b�/B�,��R�a���SJ�Ռ�f�K��Ȁvn��76]��e�ڱ/u�V{-K��Qt�˙��$JJ��d���u�J�TUc�l��ߐw�4�vOJ*�I(�7m�PKu\z���$���3l��3M�gQ������5����҄�mAUh�Vn��5��#ӆ
���$�1iAʗ4�N��$"�S�XQ4`Y�;zJ����T�ɩ����Y0`T���Niƴ.Z{n�)���n�;4�(%��]�j�r8�6m]l����R��F7v��+��55&����E�D��8�^L^R��S��#^8���c��V�W�pˊ�Q�%E�ǅIzm���
Ē�X�h�B�e�hK�,x�\;��X��ճd��$�Ӹ*@�kq]�Rue[C#��n��3Zݤ����!C�1��xŋ�y#W�n�Ǵ%(/�YF����w�4�6m�x���)�"�Gk0$�@�ۆ��zP,1yN�� �N�d�^Ԝ��Kl��`�2I����@��D�%s5�͖Uv�i
��]�O"@YJ��"&���0��][���B1](�)2^Z�h��h�J�WGt����ۅaʠ���Y7�Eq�gu��ۜ��y�m�x�;	�BBGr���ꅰZ0��/D1���K��I�j]�T��h�40tn�;g�9.H�T*�VnԘ��Hf�'���Ė 4�GC�@]��	��C1՚��M�J����ٶ�A�l2LDjv���E�+��TK��2*�UzR�)�0�w+1�y��,MXEV���#ҡ̿`n�l��e�-���ѭhA������21xuZ0��cwR��JY5I�C1]<��QL�m���#�˩�\4SJ�;:9��%p�i�33f�&��Vf�D���tP����ƣ;�����FE���سwvvm�ka��*�Z�%���ka� �I�ňL\y%f՘UՍ�aޑ����6ꠡf���{s*e۲Ɋ�䠏�v,�]�J��F�i$k��pZ��9rQ��/;gBØ�w��!���������ifL/K�|�O�+u�/aso@��%�h�-�m����aY���F��x��)�Ƴ�Jv�b����TcP8��K&�F0U�z����̺�ZQ��`˸UÔ�ȭ��]b��F���˦�K�j�K����I��p�q�w�f�+�6����ڭ�W�$c).�\u���(��ȉ��ΝZoղnX��qb���N�K���{{ֱ���U�]l.�ymiя��w�A�(�sF91�]�Te�u���1���6a�CF�g�0 ��ݽn���T��jֵ�lS.�D-�H�7)��Ot���
�������cw,k�m'}���Y��p�yq�[4rd��T*�7KH�]ݏ6m�H�&���nF�ܪ@��	��:�g5�^|�x�rf�unF^d�,6�\6%Y`�Zn).�Qn�i����r�r�&���T-ݳ&�V�n�f�D3J��� �F��v�j/��el�1�R�B�ɵ�i��[^J��ĭUn:��Ķ�/���;��Na�fP�x6�4a4R�] ��v��d�bsh�<hF4VT-C�A(�Mݖ}Zi�/0T��� ̅���cKm�nP�hVHJ�5��Ԉv�{[ARy{ov�(���z�4��m���7*Vk�3���vW3!6��6f+Bw�D�#^7KiJ.��X ��zP�-�F�b�^]��F��@�A�b̗�w��n)7ݭۣ�e����Ӡ�w��u��p��=���J�e���k؍䭵����8���+6LDn�a�ў�M��3.�A�����S�q�Z�gen"Qu
�R����8�[.�v���� ����'*ߴY��w
u�G9ޓ�k(�ٳ		�k��pC��'��<��|)*Ѵ���kJ�"*��S}q���I�tS�wh6��)Qܻ�0a�fމZ/n^��H�0�Dư��VUY����Fރ�0
���O,#;C�[Y���L��t&V�t6��G�FL��]�I��
ݽ�
Yl/�Ȇ�P?�~OE���VDi&%bV�qd�B�jBKy�L��r�l[�x4��#!yOb`67Zu�v�ī)7JÝ����u�/����([�Jb�*�Dm;-��qB*��N�e��9�lʻח(��l"��Q�.m�����*ΪK@JX�,^���Y�{��Z�@,Rl�hǲݝ��V�8�\V*X�D�sh��k*c�Q�k2��6�
�ۊ���*^J5[]2�ۧW��	۶]�WI+,�F���(j)�1nmo��OcWg�eF��3�v2�M0qn�˔���E�gtf��R��Q#&Qf �ދ����$�Z2�U��Ŏ���^<�Z�Y)�
�%�/5깵�Ko]ۗdE�%��R��AKN�������,%t��wwU���J��;�ݻ�H��B�u��%�Qu�5ڑ@jٹ�Ey��!䣕�݊���I�9v�U��.�[up�ɗwYd)��L\J���Y�v�b�6)�M�#:���ꡠ����
ñ
�.�iju�ȸP�wJ扷��e�Q��H3X[��t���N�J �pX2*�̻5�6�f����V<��)<Tp$$O4���:�Jv�д��jQũ�FLkڷ7��U�eP6$��oUc�b�\�^�ΪÊ�T0kј�J��ٹ�r,�3���q]��f��n��⬫wi�G��P.E2��D�d5~��06fB��j���B[�I�r	��48�q&���^4Y�;FK6�V��*!	d�N4ħu�$���҅���wuc2iE�/bL��X�Nۻ����2͜T�#�덖��M������:���ؔ:.G�����X��9��V6H2˧�j-�� ə�Q�w]�T�v����0�3Kop�hGgu��f�f�ZK��Q�Տ3Ǌ�-R�seЫ���P9q:��msJ�'��d����<�J����,��d�hF4R]��ш�'�,�(�%9kT��T���`�W��X1*H�$�"d�(t�f>?q�7	�d��/3Q���.��-绩gv1��ǗM(���Ɂ���G��e�>&�oDIE�+ۨ��-Q�m:�U9W@.[�q��wx],�Y��#������f�{��$��#CPy�|n]�t��F�]�����ĝ�j��d:���7T���n���RثUb�G�8���=:[A2����xi{mns�(k��dV�8]W+���z;���D�Z�l:Ҷ�z�C�Zcw��Sy=/{|��3J]��ˢ�뙪��zw8�ڬ�������ֻ��8���Ey�!�B���tɸ��ݝ4M�}�tBf��vm�fÙ�޴Q��W���=`��6�aA+�I�ɧ��ev*��/����j5*��riw�Ȕ���n�M�ۉAPaN@�<�arW	�M?ym�j��"�?Jm$�q唙.Cv�Fk9�q���k�׫�����vn1�LK�!%�LE�͕n�'�]�:�z(7�Jכj^����L:����`�܉�XR�;�3v�J]:�5+mԛ}㫫�C�h�p*�M�v�3;�RR>���8Æ����6�:v�'jM#��Z޻k��D?D���tV���
>c����m�dx��\�f.���.�.\�F���z���?%�z�z����6�&�v,�ːI����w���h��KT�g��!܎i��5e�ɯp퓊tlfG�;/\�kcD�38�H�����љ��ٷz���b��ݬ}��Mb��t6�Ԉ������D�%k"�ӧ4��+��);V�n*t�0�7��v�����t9n�66�Ñl�K�� �yZ�����E�r��LJ�R�V��Fg2�9�Ñ��곸5�]I�;S,P�N�]�%4)�9����B�&��C�R�G����2��(V�����U����)A�\�l߬)�E�P����:=U�69�P�ޓ0Ǹ����n�]\Y��@�2�8E���Nؔ���;x;!���s�����,K��l�vA@BͶ��Mw>��}x���mvM9:/�7��|y!2�"b\_g*F�03�zl��̔�)N�n���fD��P�뼨��V$$Ku^n�j�����J趌nFw�\����a�\��{i(%��-���#9�}<`2��U)�V:�}��KUL��,nE�ɦ�5��p놕�[Q����Ku��^յw1$o	s�>�ـ��Ҭ��x���[JwI�t&M�x��56��ow�ԍ��%DLzNY��F�È���p�Ld�ɸM�ɻ8�B���C$�y�eY��I��-I.��6�WK�>[�8�N�P�J2�!�#�gp�J�MZͲ'^�h-�y�z�e"��F�dh�%�H�Q�m���:Q+	�ٴA&��42��aH�t�I�I�1�e�-sQ�jj�{�b��(�j<���]�[#��+;�[ߐ��C���>�����G}y	����[=�}�])r��:e_S����*���R��M���-��q�vHo�����Aӫz���smv��˝�;�Uvȫ-�z
p����Kec����k3uT��W�
R��dSk_s�\s:X���n���P{:b,����]e ��N��P����#����U`v��D�J���ؕ��_ɑ�[ b��H��U,`x�/P�h�2m�"���Y��%�����ʲ1���^;k�,tz�����]�[��o�J96���k����Yl:� ��ǵJlk�O+rj���.+"3�"׺",%GP0������^g(r���iӆ�B�U`vR��bi��%<�3-���4�T �m�㬇!��A�7��U�VC�7:��|/{7_^'��{Y���=ܘ�KM�U��Z��Ȏ��"�쩬Mo�L�M��a���6�á"���5�ҹwI��gH�����ʀQC*�\�p�MՉ�8NoKz��.��3��0���ee)f�0�ٹ/+]���O.����v��Yvn�
���c�;�+��]q���U��ݼV�QsOf���/���/���N����FX.KB���
d�w+xU@t=�ͨ&����bC�a���i�aYy�9K�Т��(�!�鼝n{����~�(�;'eڢb�c��W�b+f�O)��[A����'%���.s/o��N�t)+��j�z���WDm�E���\>w����%��Y���Y���n�'��wƋ�_��9*�х��.����gP�v�Qn�\��:�e�t�m�n3���xlt�ō��Y;�]�}�2:��Y1K���*֨Y�[�sz'a�f�,�S��t�!�t[9�xI�'K/�}wx���l+V�:��z��Z���]���5��&
�l��D�q�[b�y:�\H�'��U]���+��ky��r���q��<�`��z�w���U��IVȓ��{��!���'9��.�>뗎�[�+�]�Zzd�v�oK{���Q.��A,|�_f�0��A�ͳ{We7�;G"&b�u�51�N-�uB4[�7q�M��|�k/����$C��8T��i�6�S��i�ȷ݁�����8����#8��g ��8@��|�t��2K��+����E��9Q+�!RJ�ٻ�kC�6���=��R��X�aV95J���5�"�.o&����I�y`<�R]v��/o��aګc����co���B9�9{��6DpD]s�R��
�Vݮ���hSr�o
��r�R<�KL�<ٓ��z�oc+r�(9�EQWa�bHs0�v\���|����:�Fs�ZԙzK�֔�[�3�N9z�`<�[���J�ǫ�n�rwq��:��j�ΰ9���ܳ2�#"��`��bU���׮ei�bT<kj�T�s$�:I
є�̆�u�˽9�;zG�k��zCc��Jq�9N�<����:��u0�,͘�J@�u_Zx�J ���a�}�L��Xܸ�q
���y�o1�BX넽��ws�Ԉ�W�@�[��>̲��&RV�^	/75Z���.�ŋ�ah���gtI$�Վ`D�I�kb�&�����&�uw6�bk�L%��X��7zc6�d�#u̣9���zXޒ���%��]����4��Y���k�[��3u]���1n���/ښ�v��=�L[f�0�h-ҵ��hp�����h*Z�Kpvh�u�lL��d�|l�QG��'iS��ǩJ5�U(�a��&��D�ʃS�@��È1�p3�k��5|<�����4Z�/�.�7'w*W�C���Yr���e^$�b��&B'��mQ�s���a<k7�lɜF��z�E��v�����T*�Fl�F[�P�*��''P�3��� *�l�q˸�zV�Z�p�'g�mޅ�ḫc9�;5�&@��a��h����u�˗�~;]���;4<����y�ȫ���K�q�]��ρY���݂-�FK�.�m��x�2s����R��<��Ӎ�2B�۫U:��:�Wtuf��$�Ux)��k]��\��x-B`鳎ڒ8�����*���·���3Na�y�c�7�l��t@ֹV�ݰPY�}`�B]��Θ�]��"�"Q����tZ����/��ν��}��$�8�t d���1�[����bm�yr�	*��C پkO6^WT6�p�ϓ��ڃ�#��yVi����#�{swss�&���j�K��֣�;D��1Z��L(�Ir����j�ˍ���wv���K2)�V�S��xk6�}��!��
ۂ�������4���h����*���Ksd��}M��I��m��\g{�����[���q�Rm��8^f,����r�K���YyC{��&K�8uA�2�N���{;��zi�UO����[+j����u�'�c���[a\�.T@L��w�&�'Tl��U���\��7WXnQ<C��:}ӰW	CuWG��ʼS��)�58\�z���H5c\۽M��3m�\u�ر�y�m˞Mk/E��,̦��U�l�+h�2�>���\E��s��i[kKt��)���s���s��;p=��=H[!��yvJ��h�o))m�ݮ��Q��Ѡ1lnRVU���Ϯ��4ǯ1���w^JÕ]�n���y��MH�A����r��*�`p�T������h�8.kR<	�Pg�¾+:E݌�3X=vMpj칐J�yL�ȉ�5p̆7]bb!*�0䱐U%
�O�f�
�6���vt+G Z�'j�`�{[2i�V�U�v�)��V-��3X��մsn��V�]��Տi�����Dso�^f$��PuN�BT����m�mo-��y���ʙ�e���vv�i�9�x�so��Lr��a�����)>�٭.ci<Dj�����v2] �Y�!�{0��������yf�A�c^��p��)�i�1�O����)�<���QI(�� ��$qVq,�
��]�[�i���bxpJ�}��f�R���c6F*�o\_#��c4�]������F�al�Ye��J��8�۵r�ajK�p�A���ޮ�z+U}�XF��^�uB���E�&��_w͎ɜ�Y}��3S*a�MG{��Ubh�λ���B�]�v�F���n�X��&$�}Vw��&:�x��~��Z�mZb[��L^��wL7�?$t旦�nݻ��f-��glo��3Xz��R���O��C�u�MXt�A�٦c���!{ٮ]���X��̽�:XZ�0�}x2�8��$�79[%�@h���}��5C�t�O&ʚ_wA���%��q��\Vf��6*��&�js��n��q]�Fb�n�q<��	���+@X�{���Q��'8C:�WW[l�9e)}ʄC�Y'VT�:n��(K][fL��e������6k��rI���8��n[<����p���)q)p���Zѥ]�tsH\����1*��/*)c!k:��7�'\�G_z2{uu^ns�*�8�z7*1�Ğ������2��T�����5�{�Pq�M�՝J�Rɠ�e=���m4jΌ*>�F��(M�Ħ��]�MK�4[��*��Ѽ�z��e��[\�@�̂ݟ6b+X�h(Z{��a�vqC�΀5��t�#='"r ���h�_��5
�v�E��$�.v��R`�n𝆨���e�C[e\��V	/c���F�9�2k�ORg�"�%)�Oj��HQ��<�y4�21K���v���qj��Đt� �۩�\�G:�!��8��Dꕜh��A!p�sV��v���᪺�Q7uȌ ���0�1
��V9��̸ۢUh3�Y�B�A�z]���"Һj�)�˚C�tqf:�/��YYm��T�f�5�;�������[�&V��ʛT�9ZVs�dGNY����>}*�m�Eg�x_e�6��w�n�L�z:Z�3���rFt^S&����Gv�հ��ݛ�F9-m����`�Z��kz�����:���dX�c&:�2���,m�f��5��µq��5�+%��}�ڝo�v��mty�"�CO�&[Q���b����r�M{]����-�6"�f����h1�+32��ўZ1i�0�8"�nu�,�����"���+S�z�[��u(f����)�z����ڦ��b���)�f��N��	�}kc�ʹJ\ɡj� Ѕ�&މ�F.ڮT�P-�;t`�%�.�]u�N{�ۼ���3Rg[�z.ٛ��<	�*n1ӇM9[B�	��[�9{|+u�rr����u��V��;�xl�]��X�oU�(P���L�\���,Ơ��F�S1I*���._��-=Iw3�d�̾3j@���ݛ���3n���D6�c���XB��ї1�
z�\i7��Up*�#8��`G�M�34r�S�����q��x]!%���/Yc��,�E^��R������Ui�[+/�w�[X�k��׵$sw6�;5L{i���5R����b�.rM&&�_v����q�30�Y�ܙ��]��.w�<�3|���
��=��v pb���=��a�G9*h�T <��+VQBb��Y,�S[c)��������\P��qԴb�n�f�uf�R�n�.��r&����<��KWw��v*�t���v���)��"[b59G^vq�����Z숺���?��Mx�wK9s�gβ�a2���~fV���h�*���Bt��Z4�>Y�5�o��n��{�*L�JJ;�q�vi&��%����(�׈�����R��N"��>� �ɼﶻkw�JG[����U�8�)ʵP=Lk��\��z/edv,v�I	}wmӹ2�T�B��q��^|�Ş���k{ggsx�`�B��mc�v7}�]��]�3��9��9,J�'�ov�+]���P��B��ZzjR�z���ƒ��h��pM�A#�@����+b�ض�\�!*���W����땳�x./vp�O_LN�Cp�Ɂ��p��=8�[���������5V���c71�(*�P�	<���={���+�m�(]�ݠ�ކ����&�b�M�ɰیZ��I�LM��Y��P����'��xD��{U\  ������N�����
��騱��bd"�ʰ�U��kz��QC�ʷCaխB�>WVt����;�q�eZ9����L��k��2z���"�D�*r��H���.�u3h������y��_�?uZX��Mj# Uwo�v�.���3�Rn�#^��5�}�Q�u�Sc�5���^����:��⓭��6�[����w{��fa�:�;�.���(�Ք��O�\k�\r�(ٔ�,mS4�o72����)`�W�"A��R��%�)Z�{R�W����|��3x�|�[��]J��5A���1�X&��cpS�/0dL�8s�
��{8�E��0�3�u�Q�&�Gr�z���S�C3sݚ���wW�\u85�U�� ���wyA֠x��A_���`�4�Bgv+�y�Y]���uxi���p'��;q�h����a����*TE��j�����Y�WO�5.R��Ӳ�]Wۼ9L��jZl�\d��`N5R:1$
�),�N���kd��M$�ȡ�+��î�� ���N�	Y& �JH�n2�B� hA�OB�LW�Ja0�W/k�C3�PQM6��,�3t�gT6@�®H1G,��N&	����	�MUS_L�֝x6T�jko���U�L�B8Y6�I��nYM�&P����M4܈����g*'r8�JJadWR�e�aPBh��5i�i�LFS�$d�O\@�	�J��q��IE��B(���1�nq6Ze�$� �b��M�R>�UM�$�.�uP��a��H��H�����K��G
iD��3��%��N	
�U��I 4�)��r8�#�4�'��|�<Z�|)u3�(�q/x_~ty&Iǭ���$�*��O<�I�b���@J��Ȕ��\\�� �I�
�`CHq%Ȭ�t�Q�
�r�pB!������ip}�ߋ+?���|v����vw�����@�T+�8%�`]�Q<	�*A<�4��JHH��$LT!�IH���0��H>��vTd�ׂ�Դ�A@��IQ�d2��c�@�6�l���2Fô g�E�Ps$NA{�C���g*"��H�I�-t�$[�˛�zwof�U-�!6�NF��,Ia|t�e����T���|�(�nYM�&P��)v[0����y6��n���� �I�˪0�C�)(h�PM@ґi���m��
�! �@�":�4�BFb���1�A!�謗t�	)��e_K�H"�<����)S��n2�B�9��[�L����{]>֟'B4�&C�,�I�� ��>.��S�*�����5{�� ����=�*�'����?opS��������?����/��G�~���������ߟ:��O����/D��Pb�Hi�|72��j�uJ��';��k
(v˄�R��|n᧺����kT�ɇ�Y2�rᛶ+�$�1�AC;.�u�<��c�ew���.'UU����%Ɂ�N/����Eś�����\v�$�$���Jnb�Sl�к�2)�Y�I]1c%vA)�n[cHF���K�=2.�.j����֬`������yIR�Oy�3ː���/� �Z�M+�:
̔^a��B��9,�K<�.���'��^��|����A<�*>����xJh"�=jQ!�T����V������X�Gq^A�>�G���q�y�n�}�l���KQb��͡e4��R=��o� �����n�;{��Y��
K9��sll��L&�s��cH7�:��U��e�
�]D񒄥�,��N�S/���̘��;I�N��O#�\�j�p�w[](jT���N�n���ol�0ݡ�փ,��j��Ĝ�_Y#<��خL��2i��]gYt��� ����vȢu�<�X�W���s$Xݠ �uLbU��b�:�cu��v�\B���賩m]�}�������������^�u׎������ۯ���n��N�뮺㮳��뮺����]u�]u�]u�]u�_����Y�]u�_���Ӯ���뮺�u׎��N�뮺㣮�����n�뮺뮺:뮺뮺룮�룮����u�]u�\u�^�u�]u��]t;Þ}���6����SX�]7n+O���aV���i�gP�`���q���7M�Ȗ;�,��m왘�u���Vug,^�%�掊�;����@��Y��x//k_v�6�������ز�`�VE&0;�<�U�)^�f�7���X��͘�����u������B��۫����s�@��5������zP� �OP�Pʴ�92�g[Z�=CC�y!sW2v�qX��sdJu���Qk�����4��+3���ᓗ0Ķ���À�ݣ���m"ٗ�<7�B��;YJ��G�<��4� ������C���ZP6�	��u�c�w�-�4@�6g��y_:l�	�tR�>��}W�Q�Z]�Ћ@�{Y$��s6�9#�;4��=�U���@��>����b뫻ʪ��\��Z�%��3�}�b60� /++����믦E����{Skޫ��A�SW�满8��?c���yah^oL�}���[�1�<�㕦�kƶ�'1�FYҕ��UR }��)��[&#5nҪ�xi�>�j��3z-Ȭe}��|S��$�i�f�P��yZM[���MZ�C�d�3�qZ�)�G�|��wI��7�d�L=�N^P��F�Ut�D��r��|�%[�L�l�ﰈ]��n�A�mr���#���oy��sk]n��A14��y�p��=&��\�2�d��#ڵ7�n��Fuʹ�"^U{�E>|�B"��?���?h\��g5`�s��9�w3���㮸뮽:뮽:�����ۮ�뮽:뮺�뮺�㮺�Ӯ�뮸뮼u�]u�_��κ뮺���^:�:뮺��]x뮼u�]u�]~����n�뮾::�����ۮ�:뮺뎺κ뮺��]g]u�]u�룮�뮼u�㮼u�㮺��]z�S���k&��$I̹w&�^˚(s���`��sH[��婄ovN����(߽UvĖc)��w[:�]ª�1� `5;yX�o�wZ;���B{y8��prgH1m'(��w���o+�Ȑ:"t����1���r0K��s�/��s�l6��ݔ�����ģ�IQ�r"i5o��V�}�tY�8e�  }[5�#����������0��'	�d3��j�������0��0������V�5�>|�W/������#8���]�1�l�)<�xdM�P���=��8�ɠ�{�q[Pw�X$F��P�Z�������R���_$�v8�Z�v2�@e��"8��X�n�/�a�KlV��4~D�IIUI�<��3:��ߛξ����;.�-�넦�+ �l�D��ǹͷ���1�.�*�r�a�˃}�ſ�v,������Eh�G�KAϜ��{�+�j��޿���o�V�k����̰���0�=V�o�tN`1�%8�[&�)�Q�>�,�`�r���_��4ڄ��]1���|	���z�1-m!�RsL"Z�|>9tDx)2���P���Xkm��ܓ�uj�w �m=ٳ+`�ی���t@�'�,��l���d���]�mV�*��R�J��,��^Tk��Ͻ�Qz���1�*��=PЪ��3�lm����)xzW�������~�κ뮽������뮿u㮺뮺㮺�뮺�ۮ�믎��N�뮺㮺��]u�]u�κ��]u�]u��:뮽:뮺뎎�뮺�뮺���oooon��ۮ�믎��N�뮺㮺��]u�]~:�:뮺뮿]u�]u׽ޞ�\������׹k�;Zz�+Ӷ�Τ��mѪ�j�H-l)U���bӣrT,�+F#���ȼ��&�T[�6gF��Y�ά�R����/*�@�Oу/��w>��e�n�<�\�M�6��ɻ׉E�����Z��ur�l��*L.�`[U�.���dFw�u����Z�����u�e�����]�q��Ӌ4�*�yiU4bG&h��+�:��o��Eax�[ٶ��>K���{��k[�Oۼ�%��7zpG���㾴�sݶ���m�2��u��N����z^f8�6g�<��Kd�V�k2�৯+��c��탥P�i4�wY{����Y/Ѹ����KX��.}~v�X���zٗ�c��1^�:-�f&v�k�R��W��N:ܗL�{��w���e�UU�lw�*ܮ��[!�+�f<ȖYݼ��-5���
=#�7�*6���C]�w�������c����.�	2I6��Y��޽
��YC�<�X�r�*��]wF�����z=��Z��ޥD�l���Wu�]*f�+M�q��(�l��/�<~�ғ��v�ͮx�C�����|���\���|B�\jTr�0
�JK�Bgu��fk<+�������﮺�뮺������뮺뮎�뮺��]x뮺뮸뮽:뮺�뮺�㮺�Ӯ�뮸�뮺�뮺�::뮺�㮺�ۣ��뮺㮺�������ۮ��㮺�ۮ�뮾:뮽�뮽:뮺뎺��]u�]u��뮺��y�.v�ĥv5Y�cd:b��b�kb���;;��	'8Cx�0�C���ܭx��q�5^wI�g]\��nj����8�~4:����u_�7��Non��֏G�@dpyG6��K\���M{Ab��2�b���V�5.��&v��5 ��V�=c��7��~�L�{"#��N��ue=Z�]e��tz8��쪛s\`�Ǌ	�U}��\�	�(����w�󲱃��ޘ��� |�aX�C�x��I��l;�yy��\����Oss��E ��|�}�Z���v0<Dm5GR�E�%y��U���5�r�J��O1�3�����` c�:�O8C�f�2��n��Y�R�*���+���SNUz��b��oj�x�C�{��ݒ�7��Y���G�����͍m�㛂`�䪖���p#�Y������ג��D��Wu,�cm>%���9(pU�"�z�jwճM� $zsA���� �q��D'35پ�ȃ�*,v�ѱ��uö�bM�W�P��t8WY��Y�i��S,7+����ۯz�,<
w��@%.����3�.S���p�B]�p��ƯP�x{��:�~��tu�]u�����ۮ���G]u�]u�]tu�]u�]~:��]u�]u�]u��]u׷]u�_u�]{u�]u���]u�_u�^�u�u�]u�뮼x�=��{u�]u�_����]u�]q�]zu�]u��]u׷]u�^�u�]|u�^:뮺��>�q���\�T(Xci*=[���ۄ1giv�ݐf�,T��j\�$�3��b���v7.���-W*�"���Y32��1M��j��b�m���7��m�˟U�ިٺz��X�̀�Wb��4V�9u6�h�G�'���t!�_Z��u��@9�� ;W����3C�r{�u�u�.�Ed��7L���+���^�>�r+��{��;+OV���������wn3�B��A�䮝@�I��y4�eh*�d���9��lH�J5�nśn��݇��c�U�����8εy�/�9FJ���n�}�{������	���;:�'���w�����EAػPu�]�-N�E3��&����۽�;U �=5b�eɡN޾-��[�R�����J���S��nsz�gw'$C��l�Y�2)]��lT)iC7+j㡂��S�ܹ|��!�we�sBɓp!Q�u�MW�Xn�.٨m�sHmk��%�|��V5�4��7��pʐ�̨�����W���v_5tƉ�Q�杖�Qg���u�r���;d*ƨ�R��Q���g�j�{Ҳa�)�댁���&�vc����t16:ɛ�Є1Y�S�յe�ظ��[�����z���~~��']g]u�Ƿ����]u�\u�^:뮺��G]u�]u�]tu�]u�]~:��]u�]u�]u���]u�_u�^�u�]u�uק]u㮺뮺���u����{u�]u�]x�u�u�]~:��Y�]u�]q�]zu�]u��]u׷]u�^�u�^��rY�̲Ȝ�]{�you�<��N����R�����i���b�y6��寅1}::�_�fb�+��ɋ����q�'P�I�`̬��09 �LTGR̜��3��|;�ޒۭ�ՑJG8t:��c�%[�y���/��>*�N�,�R�,[�.�S�"�k��׶궟n��m����s�xk�e ��KW1se:{��.�u�&ޑ���W���<<(��CY.���� ޼�}G^�Cm�!��j�bW<�Âa����s'_Cf�=7�v��צm��ѕ2�u�uek<�j/�V��V��{0uB �w������wD�r���{YN>N�j���sg����N��:N�f�;��o��"��l��7���N�9ŵ�-�l���^��}|�}u�YE�u��Q��a\&��o�VwU���{Yr��7h��
U��T���rVN���l���'�=O�b]=*�`���T��.�������GaX..
�s=Y��G;�v)�\�v�[��5~��X�[��R�ܦ�]��/Ul�k�q��]0��H�x-)�M��<�H���N,Ц)+�[���[��u嘃��t��8:�ز���F�������B��!n��q����pPޣz�H�3̔�m�: �uI>�؞݌�)gcE'��j�f-�K&��*�D(�-��b�����`�[MЬn�%�Z������2�]Θ����*��i�����U6N�p+X.�l�H�G�z8��7[�=���^w8����뫯ƺ�W�A��f`��Y[��Og��Q[��v�BK��:>F鴐mN^�̈�F����y��E����W]�w���䞝L�����Md;p�X��N�w��`�r��<�7W@�h�ܰ�))�z��Z�yZg�Ѿ���j�[0%Z�)o_���a��J��,�����	b�&�%��e�L�h5O�DM��b�ue�5H]�z����f�O�Y[v�
<j� �9�9+i[��+��`������_R�Y;��}E��0up;cܖ\������Y�/ǀ��S�{�X��v�:N,�P=��6�U�b����nl*Y]�t92���u��d�֠x�j�q���&�e���^'����V.�<���)�_�UR����P����2�6%Z���;��a���x�ܻ��;@N�|��u�{���c�H�Z]ۚm�1�3S��u#�f+��f.J�d����s3�b/@m�'@���w]fvl�K�m[�[�;�A�꾂�����m��+i�]u�{��*v��u}�f�U~��ū��%*pI��"�������Z�t��YcU�em�7�IWe��8�0o��w-��,��\�BL��Tm�����aSum�|	{�8
��ظɗ	�%5}�W{'n)q��)��m.�C�U����Z��o-%t�3��~s/6!W���s�����N�ᦰ�l3��f[{J爎3�X��Rj���ٮ��V볹0���nɠ�'���e3AX���h�,e��,�"mw�:�bM��1�Lm�2o>JVxي�'DT���/@��qF�*|2�\ާ4���O�TGwF5!��c�a��m����G[�g�z('u}p��mm��
��.t\��jpL4ɋ��NƎ���Ϭ��7��m�a���s��7r��{i���
e��gB���AGi���!�y�7n��Yl���c]���A����#�s+�v��ב�v�Ջo]r6�Ip�պ�\b����f��y�{B�~��.H)x��R���E�%���k���n�v����K�:���ʧ��<�K�>����|�a�M�'��h�h����n�R�a����ŵ����q�t���l�(�C��v�kk�������&����q)VlN�:��5��^����nM4C7����W4�c�<ۺ�q�=V�+��)�]�i�"!a^8�'-�Ш�4n�]����m5e1׭k�}Jr�+/���M�9x�ëNۚ2�A�\�5V:��}9EI���1��0U}�����a�
Y�����K�����ee�$��6�+���3ܒ9�uv����*�72�:S�o�IZ���]B��T�ߺ��h�B�l�K]�.���'v2�;M��Q�$�j��[�)>��7v�ܧ�6����Z�k��;���Ѱeg�w�wb�=��Q[}���nq����{˹%�;`���*�ֵH�*P����}ƴ���+�+�&^4�������R�{�,p�¯m#�pX�aCf�"����ˮ�������G޷�o���∂��#����?�������<�� �C�Ì?�/�	J��%(䈒B
Bc�q�����?�|�d�)��`��
��M�YJ�a�Q�2�I��I��9��Tѥaa:*��eIi
HE��p�j���iG%�'�:�ȍ� "-(�0�
Q��C0�ڌ A��E�h�\" �hJBr�d�A�Wl8�}�V"U�_ESQU-\��Csyk���_rգ�X(�cv��]�/.^�`�3;�G)��cp�l)��%5@�lgP��+���3W<�\O�������(�}'��6R]��ٷ*��U�8�-��oI�W}�fR��s6�m���s�kVaI��9m�i�����։�{�8��3Z�dg�vT����C��j��n��6��y9�%�ڝɋb�gXy��u�٬/��r�#��d)�س���eaę�äE��`�C3g;c5��u:@��z�L7����z.�:�C�U��o��(�$+),A�uKElt�+�"��qN٬+zD,,�έq�>yskx�!.kY�ʖg�~��̆8���3�K�����Y��U���AVWX�ϗ�9[�!�ڰ���p�ܦ�Pp��8���7(j�2�|-vN����H�RoC�.r���W<�.�/�.���|����n-��s���=S Ҕ��Tfu�Y����ݡ��
�՛J��H�A��SBQX]�n�m7�*3�,;a]�ڬGQ�0m��f��P�����Q!U�
��F��"�L5�If����Q��	1 bC�&���5M�A
�P>(��X���t�-�4�:����PQ��2n�A�{����K�xH��N^:�aI L'6��)!e#P9m�m�O\�"�V�P�L�5A��
���E�"�4�-<TIhH�0.�q1w�DBA	p�'����J�Pn8�(��¹DJEF�p��H��,���ADQ4��(�Q��	��\I���D��:�	�-*16R�FdH��C��LI�K���.��6Y@�1i	ZJ�)��'*�\A>�i:�<��v�_ד�P�j��I��A��>>:��������Xw����Q��ED�d���h�0�QD��D�-���J���Qk�糀�s`96�O}����K�Εx��ԡ]B<�i�y�Ce2���i��v�F1Q�\�������{|ݾ8���~���뮺��*�+��aI.6��"SÌ��c�a�;I�`�}*�(g�6;�q̅���v7T��˻}vA��LB�E��{��	`[��@L��`s������mz�|��B��#�����
q=:�+ǧ���Ƿ�믬:��s���qD��f�\���W�ミQ���Ͻۙ|��Z��2v���������՞����U�d���_��|��[�}n�_]}a�]u�������:;.��#���1��	6�		H�sXu��;�#����݊�YH��>O�L}p�~okv���O������ϯ���Btu�T]��}c�yx�t�J��!߼p���L;���w��c�k�?�����=��pS}���{}o������}f}}}}x�W����8K��^f��Hn�|;��g�L�G�d�O��w992�L�W�Ϣ�(١BM
����!d��ЅS�6E���a���q�Ai�F)�O�}q"��
(�i�9"��NY�L�D�K�uR�~�7(�4�(C"0�~�~|�=۽��s�}�<��R�H�(�~ �s���*�V�n��t�Υ?��ww�ﲋ��&ty9b`�mqo���;��N��i�3-��*4X���-ז��wqt�{�d����������CF�m�t�" %QK�6Zj�(�$�?�4��7q�򽉣0�:���(�9�w9N߯|�7~��U)��7�����j���W3<�X^9�O�ʗ���{��^uq��{��:��*�fqn��<��}#׹seQU����%�_�0�M��	j�rjIM�c�s�F4��~�͗�lğ}QϮ9Ƨޟb�4���̜�|�^���e��=�ѝ��\�]`��{���ְ1omsۯӞ���[����Ӟ�?�����=�:��eH"9������o 㽾�9$��7�[�oՕ��A�ٹ��i��{C��4��r�����g�'��ݯ�l���;�Q{��wXjf�����W��2�z�S	R��ZI̹��ؓ��|X�q��-�"��&��W�s���~�;�]
Tyt%�Kek��.�ϭ���Ml}��
�U۵J��s�Qp�,λ���:�W�c'9�.w�ƺ�b�F�{���s�׊,(-wwWpwU���]ĝ>���y��Y����|#�v-UUt�	L�^��Q�Oz��^�v���9��ه��{��{�<��y=ƶN������;�z�>C�|8�Ζ}~-]>ؾ�	I�V;�[�&wh�{�}�L�R[�[%>�������3�=����e�#�Ȋ�9����Gv�nl[��`�Fr��G�����M�V��ڝg4�z�O�]�{-���������%z}�r�Ϩ�2Jlp�=]�}����Vl��k�W� ��r���]=�ֹ�g�H��r߱�o`��_TR�Λ~{c�^�����7_GQ^أ+5[(��g����1d�D�q �h�$q������S�mɊ������+۷W�=#%��0G7.���{�	�ܳ�j#�����~��'%�|E#���*������������ޑ�c�jY���_jbwҗ�*�w�O}�j,Vk?�W�$;{^Ps�>=�5�������L-�n2��vըm�W�S3�^��!tec�C�:�5�!��J��L7{[��{+��^������[�Ⱥ�3P��n���m���OIR���ho%�S�n�\6�Z����|O:}Ԓd�b��m�@���> �һWn��A�Px< +�칾��?fA��1]in��4�D'�^��j���������fR߆W/o�E����a:ù����"�&z�Sv�Ooܗ�.�j���7��9�[^_Z�n����oӎ��,W{�N76��zh��ea|g��,�U���fuaa^�c܂6C+}������3`%E�-�{}�nG���������ɞ�A��#�t����z7/��gp��}<����5��^���m�Eg:���wW<���G�a��u>�H��w��f�e�(�Z7N�+�qS)���~I�Z{�O���W��N�(^��1��g84�zb����g��~�cy��a�[��6��A`��~�I�Z+�QlW��z^�/{�N�N�䒲�������C�m�޲��z���������
��O�R_t��d�e�����{�K^�C7w��C��%�=��P�b�Ҙ-_[�[U�s���CqV�k��C�<dOP�6fb�)�*�޾�)&m���{��C'�_�q�i���kzf������s9Dp���^�fl����a����b����w�x��Ϯ��s�8��S�9�]<�B���D��<��}��������_yv�~�<O�PJ���ۚX�0ui�Z{�u��w]䅠��6�	Z�sۮ�}"kv��}�,� Q���>>��_�۳���o�+y��e��WVC����[��ZD�vo������?]�5?�qq̰Q�X�?w����!��K����iQ���	����3��7x2n�/�ׇz'��y}�ئ�����۱���|]m��};� ����4�N0:�i~������zE����1�iz���� g��^�c��X���a'$wn��߶/�������@n�g�,��'������2kv+�>�bx���:q�,�ۃD�AɎ̶���&�0����}�/}�z�Z��T}�������i�	�5�U� ���ۮ�����J:g���¶�Qxvw)��h��z��o��woY�&ι�ꚫ��l���B�D�̨	�DH�p�	yOz>}�oɺv���ĽP(!�c��,�\z~{J�W���貭:��X��Dv�,t�ᦆI���Lf����J0�T�<,D�B0y��P{G��k.�b�r>|�m�2�0��@$���������[}����l�y�$:k��}wV<٪ֶ�77z�A���{6Dh�af�sdm�7��^F>Ӧ�E���~�ES���P�Is�@�R�ڕ�BP������_{U��<4W�g��.���
ܟ5�?q���%�Ar;A}/���;��T�a�S��R��H�4�l�?ndv3)�|c�R��w+z��e�>��_���K��w����H"w��{p�_Y+�w�w>�v}r���4&�*���ݞ]ϑ�E�_j�+���l�w-��&��׉����� ������$N������Y��h��!Gl�}���o�.���s��]	�|��fi�z�v5�e�N�{}�c�}�s;�����+�*��A&BS����X�׵�J�6��5�m�E�w�a��-��9m��uCp�qY}4k�=��TX�g�L��ϟ��Ɂ߷?��̭��]��To3����ޒS)|{6��ݠ��u؝�`�aYZ��|r�����\�}���������	^ަ���	��N���C�N7����̾RJ.�����[��g};�x:�Fl��;yo���w�]�ǽz�HE\H;�7v�st����=���mm���F"Nm;�t�-��5S/M�?q�G�g���{��}��@��sW�^b��-���~=��es�,�ޕ�]O3�9f��C:��i}uJ��i��b�;A�����/��&��}�٬⫆K����"}�H:'`[�!�����/4\Y����Wf�뻠L=�	�W�*�|w�!_,X����K���L}�;7�o��� ����r��޻\͋�2^8Q=�3���=�f��	�g��I��Bo�|���o��/n{B��v#�e��]�����8�Nv�����%�GW���߲9|�*��oA�z���h���J��Ƅ��J�
^���9����Xr{+�6�dʚzR�hQ��m4�];���5�o�^6��h5�o0���!�	�.ٓ_ۨM+���@���KX��y����[�:!��`�!�x�g_J��U{��z�Q��f���ݵ���5�{��v*@��Q��yh�5H�I+'�_a������g���T��89��۵ j8Y�x�b⪛�����I�۶�q]{�Y��v4��m����uQ Zy���ް���K��U���;���V���xTbw���^���>�/��=`gzJ�tu��u�;�������R(6�Mi����H�+����+�i��{�s;c:�艖ူ��|n��r8�FC[�7'��������j��0���$��Myפ�s�����+�Z~�zyό���=�W�'���n����~��O���d�d��.���̱�o�C=q��ʓs��VJ+t�ܝP0X�ͬ\����9_87�^?zt�ެ�O6��;�|�Y��!��,��7�o�ۨ��Ǳ�/wobb��]�~�4߲!�Cy�P�Nҝ��N�zf|��W�v�9��{yt�c��0o���/8g[0g�rm�L���OL�Ӯ/]`w���s�폅�%�v:���[����v-�¤�]�Q`�q�W[0{zf<�.T5�R���J�p��u�y�+� x��!�~��3�뱜�n��(o�������%��Җ������:�տ1���^o�R�z�����<X(�����|r�����Uz ����22��G`/7�%A4؊v��v�}_R�Z����ۿ<��?_E���9M��0����]z�W�M���GHΎ�zݠq��k�v�8��'B�]�J7�̬u՝�M���I~�roG��I��ؿn���$�v\�y��1�Ơ���W�&�x���b��W_H�߮Û}̦j�U;~���sӚ'������^լ:9]R��}��.O\���+����F�>��r�,�,�H��t~��F��	�6j����4�I373�g�\w=�@s�k\�9<QW���u�_=��{�'��U�lvr	���s�i��:���y�l�,�m�)o�����z�`�u�`~U�r���|hcE�쨸�h�"`���%L�gH�x0podln�Β9N�����/��j^��^R�.�]�+^i{��:Oov�FFQ6�$�4��dRH�h�&0� �R&�O���y8!|D:�d�-�
�cY���o:v�	�CI�d��w�����گz��n_��g���� �>�^�'teEr�0�囟O{���f�0۾��=���A>���6ﯗ8��==��po;d�O5�T�g��__{��4w��@�߰p��8���&^L��>�7�.��~|W�/����<�����w3j,���ߙ$�����۲;�v	Ŝ�|e
��]�z��Dgz��/��M��Yy���m�9�d;�|�6/\�:� U�����p���,���U�>��=j޶p�X���dc>Խ��~�]hvL8��y��ǠH�I����8f�H�fŰu�� 
��{ݽ�� G	�k�/�p�N�*G9��NH}��w�W�t����K�N�������y���vu���ڿ�E�ܯS���`p'ӦUW���͕�lW����`���"���^�˗v9�MԸ|�^��=!�<��ք%��o2��,=�6������ߟ׺��s�������|v�f�2�k�;�NM����9��
����=ʰ�<�)t��p��K�m��!�I���Hyk*p?+� �Sr�s��Ļ�s:x-'��fC�\	�/�t|VuD�v��s��a��j�޷rI�Źo^�$=~۾�T�;�V�%Tg��Y�`���fO@�|�$��s�E�'����w}�e<x��7����n��|���G6>q�/��������t�tc�����f�� �fh�&D���b+��vl�=;����sn|mA�^�]�N��87���"�kǶ|��U��s�������{M�1a�r�Q>�'�����]�S�XS,����7��߳hLdQ��9�x��%߻C����zO���9��7C��i};=�+'������0/莅�H�}�>�t�e��s�]O6�8,w���~��4��W��z_�y�8u]�@k�����D��y�g
s�P�����8 � �߅�jh��2���������F�f���7��\b�ڦu�
��ʲ旴�75T.����VN�����#.򓳇a+7����ᨩ�M=<f=�*lw��wA��g	,���^`Kϱ�%v������vKl�o �X$���)Z-̧�=lP6�`�T���� {h]R� ܲМ8bv_>}!f;Z(Q3�o5�*�1���"��qn��:p�aE| \�;���I��P�s����߯����%ʓO���aCHnt3��c�Kv�*�NuIt�:x�i�x;�uٕ�:�UݐWe|�uq}/.���c؈�%֝2+�C��[Db���3rm�vA�d�Zq5rĠS�J�0g#��p��O5z�w3�n��5ˆ���k+��3n�<��$V4�&�:@���层�5�c�]3���+��́���y%w"���V�^U��p�)j��.�`_A5�2O�헳���ܣr��Q���2�Gy���w�q�W��v!���ۖ�1��Æ��N9O1D�]��6��։{�����y�+�́���U{�zZ<�¥����R�*�`�n��/��H7/�we���'[�ES]�X�z�9(�v�5����R�q�]W݆���ЛƅH�RњL��%s�;���܀J��^�hjL�F�o�������v�2���H�sVn.[}t�G�k^,r2��u����d珇N���䨵l��N�V×m�m3j������e�f�DI(�)
<=s�:ԸCGt����¯r@lV1X���E�2���HJ's>�$(W� {�c45��/v��q
�{�1m�m>E�����(�Ћ�(��/�z�W����fc��{n��[���L�]
U��	�DGך.�Qw�ԔA��98[+9����� �&��'vf2�49+Ce��Պ�p�[w1ȹ�'u5�����#�׍S1�V���w1N;�5��Y�y��On�\�GGwCV���9��za��r�92tOh�{����e���e=ڰ��/�Y��]q��q(�8t����'rL��fՈ/���Q>�ڸ��]�ڦa%o.<�{�6��ԕ�b��[�(\�r�r�*�@|s7���O�u�跟pV%�&L���a�sfJ��ȍm���o�szp�a��sM�'��*����ldB�ξ���OV�+R���I��� v�tk�㹋-����\[�x�лxc��Y�����s6��g^:��ÅTO��]�\8C��j�ݨ������,)'�#�T��{��x�|5cɏ��c�f�o��١���[�� h��s�{���}+b�]�e��s�P�%�,s�쫣�Fœ���z�9�-D�,�
*8d,��%��{�D@��7nݾ�>>��]g�}x����ˢ�.u!ӈp�r��S+U5�If�r
��T9��o==�������>�������u]��G),O�0�9E�Cq=���
�6Y�?����}o�_�����ϯ����w�Å\��Eg[���˜��U��9TW4�"�G.q�^��:���q���ῳ�o������5"�(�I��5e�j��*�G(�p�*뇯�o׷��?__GY��o��p�2!օ�C�UQeEq$ ��E	�"�ʨ��Es�׷��������ῳ�o����ۨDfAF���i�Q��2��.�r���T�RV�sR�z�DTTC��.w3V,��<q1Z\:S��T��D�d�ҔL�$
�TE�D�B� �Ad�,ҙ_��E��Q"�]���W�I?�(���\y�����n=�5�D72�+����\k/*o`mK�j�l�����W���� 5�7��7���a�f�I�Ͻ��iS!����׈{����W��	���[��S�^p�x �� k�R�`<�6ŎZap�l�Z�mc�����r�:�>>��c�??:���Fd�@��L�����ѝ�8�s1�hN9yrj�V�d0�5q�y��ݐ>H{������d�-�����=	�y�Fl3x���4C8��<�%Hx
���tu�t�CP��'�:����N�ɿ %!ɜ_Cÿ~���@��6m�{?6M�dksr���������� �N�6x.��L<mW�#�T�K��
#���&��!ķ�_�.|��5w)����K�hC�n0������_@ŋz�İ�Y@
�6z�ޕ�a�j�7>��qG����t�U9	 ��0î #^;��lbŽ����ꅩ�)@oY�^���v����!L姈k�eT
}�`��2'������"�[��%�"�n��l�:�&,m����5��W9.��,�&��]^�x���\ )�@x���|�����]���^~n`d�d{�=���TE*M�/=���ozp=�ѩ!�,����=�b�|�Xx'˥<'���լsI�W�0���ށ��q�����r��~WdX)�r�c�c�>i��������$r�kާف�n��)��U�*�=��	<��17�=-���4m=yy�=b��]g��7�=�}�-޽h�1�݌�H����~a�����Ofz�0��}����;���\��Cd�m�NPv�B8P2��1���Gǻ���5A{�Q x��E�;ܱKnP���=W��u�？�C!���=��aY��Et仫�	S�����h�Yl�8f�%$8�x~�`��>4�[�z�?���|'��pe/�i�WQM��6u�������������;�G)cC&Ǣ���Ƿ`�v1�H�G�|Ǽ��RKN��h���g�P��3jg�wf����ߨ_z|�l��v��\�F�-��,5^F�KU2�MW$N.l����#�s�!��C��Xj��E�$ϏǏ���_>>h��p70ܣb%��7��׹�42�fז~u��r��P	���á>�D���<W̦�E<�:�����	�j�ٓݝCAp�� �N�#f4�tw����3阇�y�ّ1�S�R�n-��ٽ�@���r���j>1m���y	�cx]٘G�3->�Ҟ춸'7ܨ��\�>�
�M���]�W�s
������Y��Ր�x!�ui��B��D=퍩���^������v��1~�_���ȷ�Y��:��})p�:>�B�S����;}�Y�n�h�	�D��K� �&�l �v9�;���0qӊ�s�y̴,��9_��6ڑ�C�î$�V�ЧS��y�j���Y4Ѫm���h�2�l
N9�o8w���3���'��*�θ�|FWj����X��D�A(ᑂa����o�W�A���]`o��+�lP��ߚ�?4��J.�Rٍ��;7b����� �A��ѵ��8�',�2�N75ٺĽ'�.�J��3aC�Z�=����^�ew��*f�Yh3=� =��{�5Ӷ�u�	iAשcT�;8��&ԝoS&������\���C�=/c�U�v�e��3�w		�Br��I��1��1s���:*u��� 3�E���*�]<�A)Z�Ӂ�o+�%� �B�*)
�66�8� ,3��-���1{�Fc�q�J@��s�����Ϡ6yw�q��m�g�%{*y���<d��w�D@��Q�hЭQ��U��)����f�HZ� k^�/�Uj��K�b�­��{ h���7%�S�C'�����L�9n,��[ij��-����no����wwH�:P7υ��� ��0�-�p(z�,��!���昴f��>��\�O���{RӸ��U-iC���8��
��(w�ūa �	'�)��T"?,"����S=�8�/?g]��V�E�;_�w�Ƕ���^w�F�m:���dᥜ�-ܲ�x���8��%(�z��3����cT�(1f�X�3klR�2��Ȏ�΅�Cy'qb�P�3sB���C�k%���n�{�+���ަ����<#��{�7�ܞ������&6;��P�Xzx�-��⊵�xt��\hHw�D�č��`���A��r�~]$����1ޖA��M��0��ᱽ�gEqY���{C���I�E����5�,a�#2C�{(�|����&�
-p.�FE{�����SϦf����d�' 7^4c���29��*)�R�F�W6�Т��5���r���~׺�>ܸڝP	Y&͛�F�Xm��������+���^�tK1qL�:���MkSs$M���������S�Q�������6����|J�!x�͓s|��[�)$J$�	[���7�S����{��>��V4���\��o�gW��MH��	����W�R�ϙ�t�m�}6��Ơ˶n��ּ�,)L�&@�]핱�Y�gh��,�k�~����׃��{���|���w�A�)E��M��J}mJ9��X���P�(�b�g��cw�ʺQ��W��?�n�;7z퀃猨b���T�_�r�/^s�Xs#u�H��^Q���l�Cn:�2��h�g��\����i�J��"b���;����w�[A�Xk̝5��~ܮܯ�$H�(��O�30M�o���w}]��b�I�zv�<^Z[�Ӑx�&�o3F��5��P����l] k�3�0�3z�}��}���z����|yπ�Ĝ+��	��k�ރ.C����,~�4��-��V#�4ڡLT��2sw��\����}�@B�\��X�%`=]}��9�@E5|[Ck_�:@���y0E��2lA�c�у��H\�W��XN��s�j}2'Iϯ��]�ͷ�Ӳ�*	nɫs��Grڜ!@��\���m����������GB8�D�?="���O�~7� o��D��,��ꀓ�{��0�t6�cY�6����C�l��f�ga.f�a���P.J�|A���)���ю͔hf_� <�3��7��0��H�֒Lbcտ;_Q-0$�@U������S}|��4]\�qp�<}�z�w
��nLz�j$x��=i��a�ڑ_�el��!��~�վ\�=��g.�,����&�����b��K��DyG3'�q�W�2 w��sU%~T����\w<di�C	��S��`�=�e�TSN�- �2cU��T�+�;�T=W/-GL�5y���, �_xs�̓~�M�)����>�͖��wt�OE%4.=���n�����N�v��ѝ�oHq�P��&�ѡ��M�N���H�Sd���I!*m)|����ۍp�%�������66(:�{b(�1�w]�]칿p�ϟ>g7���>��0����ߗY{��>c�聬k�S����Y�=P�E1���=�N45㾺�E�:V�'/�'�^^΋mj�E�^g�|`������R��0��*�&�k.���[����g�^��܌�&���	�������1<"�a��%�"q����̗F60��K�}���b�b���2��k�����rn���p`Ša�/�|�����&~0V�F^�˗��!T�#4��)]���al��k�Ŵ45�����w����_L�݃��<�f6K��+ђ�4�h�/�([!�O5PKH���~�M>����ts����VC|��W����;M�<�n�ש�82�&e��d��o��\�pg���=�L�3Ps����f������M��x���u\��#!��y�K�����i���8��m={>Z���bm��^lIӠej��D��?q"m����f�� ��ֶ�<L�ת�4+\��tsK՜�\�3�]%��|K�bD�s3�@x����W ^?Kd��Ng��U���)�S�9ٴ��w	�w�j�\�_۰K�����|w#g��<r�m}]0T��*�r��K�ʷ�ʒ�R��
�T3	�`�=���NDB#j��#��wI���=>�rr�q�MŮ_��Q=���2[N5���w��4�kqdT�.��	�c�����{D�q i��"2|y;�]�{������"e3��<C���9e�Q��#�ڲ�z��a�Ӈ��a�R���~07FO��ϩ1�5@�����*S���H6)�5�.����;�7�:� ��>$�hzLz��{Wy�S��z �Y���P�x��HSE���q��؋�Q��ΰx׽�m.��iU��O�qc�/���:�F�"�>��x��}�|�V� [LtD|��^\)�<v�nP;c�]"�j�Ǚ_O���inˬ�.��]ݭ3�y�g\��c�nS忇F�	jb�o�ג���7�0�A�^�"��6�.a���^v�h��7�u� �G�!_/��=�c��>�&�M��=Ԧ�+�
m�߅�G3({��/��ΕR��^���81�3�L4��8 N�<��K'꯬��?u�L���wF���'�Z�dϔ�g,m�3x눌h�,��ㅊZy�m��*|�u��Hʢ�+����gJa;0�y����)�tsu�lz*�O�w�n��8��e����j2��D��8�"��
���ԧXT�8�֟}���9:8ktRU�Xٽ��e�v뽗T��;w59�7��w���rLq��ՙ�V馳C�ۢ��]֎��⾶���P��R�=�������.q��v8�/5�b	*�^ci���>����l�#��n���S�qd�ٝ�k�?�� �3"�Ҟ^K�O9w������w��2aEG�=v���\M\����/�T�Y1�F����R�1�fW��2�fP$��m�X/;���w�3�����j����8��Ñ���R��V^��Lb���~G��G�}�ɨA��N�a濈@��ux�;���߹ުN�͓W�m��:�1k{�<����t��	�����k�'����'^j���a����St��9w�����,����px����P���u	0}���Um�p�CyX�W>��8����k�8e�`]�d:�p�U���E���	��}�d����9�n��>ý������$�mjL%�Qq�}�% 9�[�(u���˴	C��/���]�0������f�EK'�,�Nҍ�}<v�0Hs
�c+��)[��\	�鴉vw�@��p��nٚ'������;Iq�t|/����u�m+K	6l�? 3����04#�\���c���'N�o��sk���	M.*�S�����o#'2����R�?i���!��2l�{��|�+�|�g����{�nt��ߣ�
(I���Y��A�B�Y���̷��'R�V��u���7��B�<$ ��	 \��ڗܘ���gu�E@f!�r����C�T�ɺ�.b��y�Wk�e,�u>WY�y�N�y�7�y���l���a��VXaxH~M(ϙϝg�=si	��x��Y^2ܞ����e�g%�����7��F��O�u-Sֶ��."·eEoe�s�����<�4z�#^�EL/޽����f�+�)�=��m�@��~J�<�O<�&�u����{#��c')���;�v�Ϫ}�k�>s|�{�=k������9�
��Z�J�ż[�W>����J�p콉�WCG�]�
�69gcb��	f��J�����9�d��cӉ.t�@f�$eԮח���=f�a�'��=�~Ն�������;�
��h���	-=썞b��_�~�� ��v�s��v����Sc�-��/�C_�(�X�Ns�W~`W������kK]߷Ku���p&3&��?�j�\���|��>��-�;T���Jj�#P�;|�]���K��.�
E3D��]���Mx�y�Zz��@��O�[R�����b���w6N|9_�׏;�i�+�<:��9��/m�0P���C����"}3�;8zř�V��޸|��&z�.?H���z�ug�f�o>�\H�M�_�{sMs��C�|��Y��̞k��:CŎ�1����a�`{�ˡ��r�_f�JT�,�c7��%[ڇ�i�V�@�Ѣ�cb`D�}0=����ה.�R�d������}c�D�洝��sp^��Q�e�GV��g0'��u2B��t�ݩ]Z�����������!�@�z�TW)��e��1oC^]�;����&f�7<�"㳿X�4����2)����S\��tmj��J��!��4�uuD�6��<�8
'} LG�fУ E�OSQ駚vc�j����N�[�;ث��ګE(����R_3���>l���k�k��P��vۚ��� q�Ǧ�M����X��m�֕�\�<�e��J�,TFy��Aז7�c�Ť�?���YT��N᏷e)�xi.z%���D�n-#fi=Nq�r�\U{�/*�ZǵL��;�[��4a�	M���cK.k
0Co�v�v�,\���߹�����O�U;�6>]���<���5 {�j�:�ɀ�9d2(r��F��w+��u��XCﾁ����[�5�R�Ѷ���ss��~��v/��E���2a�z�����oV�����������7�+�vQ/��ga|}?i;�t�l�<wDe�F��w��_O �>���泬���@��p";�q����%]L��pe����ϰ���UkQQ�-j� ��f���xTl��FS��'r{��'�G+�
A� ��Ƃ .s� 8�%����0�љY����9p���ak�ҧQ�y��c/�5��$�� �F�����V5VR��{)�e��e��*�2�VK����G��s5��%�K�Zr-h�m�cЌٛ�0�+{�+*����s�d<�⌆�֦W!u�eE�G��	�g3DD����\�U���R>�ƺW;�.a�\u�]<\�9����G,-��n��7;W�|��͈̯=�F�VF�e�z���j�O�{d���k��R2E\���EFR+iaׄܩ�*�y�Qx;��X\Fk%�'Q�9�{���m�]b�6��*�6����=C���]�nGxBu���=
�Ul�w���������0��x�-����r�tk7ws�u@PS�.&��@'���'V��լZ�՗�f��u�̮�fq���]X��S9F�(�
�4l�����o1�^k�F�`	�q�0Yci�K�����:�Y�ZiP7����:�k��_5��[�TS��e��v�M�mI�2�V'U��g�r3+`U+���ЇR�냦R��S�Q�V�gw�T]a	Z�]�����مg.�kvn��������6��i�R�0׊�v���{=�b��V�0[��I.�c��y�4�r ���v������t���6��7��e�m!٢M��IqC%���]�`J�a6��V��L-+�A´���Yj�ɺ*J����`b�JL�xy�3���U�W#<�����Щ:ի��B#Hu�"�m-�Ȓd�i���G��ʁ�l�h�x�gD�~q�$J�PY[���i��ݕ�Gc&s�=�����d:S�w+�A��*;�B��-,�L��@��Ym=�2�!Ʈ4J�*]���}b��仯7��~��V^�`�S�
N��}�Z���b��>�����ytɓ��[%k#�[��u�^pF]:/r��2>UE,��;�UJ�j�.I��M{�[��k��*�^K��T�݈�1(�x�\M�6H]*K����gRx:��/a�e�9�Zs)�˨����6�c��ޚ��v���b���M�t�L�!v澬����Q�`ތ��)��w\�|��0Ź2.�����{���LP��6Ƞ���`�7��Ӫ����j(^BG�jΰ1�f)�Z�x��\����*X�鋮ǖ	��΄_cX�78v^�u��ӭ��!�:%$^΋.��1gOu�uC�f�]+����Y}(�|��x��_f�6�O���§t�Ǣ磲$Y���^�C0�j!���*�ɶ���Wv�N9x/P�4��Z���]Wz�5�
m��Mdm�r��;�ܣ���o5uoj�w9������mu8��8�v�޾�}��/Q����3���+2�щ'4�λ���h�Uu��Nԝ�,�ˢ(�5$[#�(�E��;��N�R��Cr
�&���H�0��e�b�5�!�#h��y3)r�����"FM'N��UL�uB`+.��"�;u*�@�l.Sͮ8R��d���],4���%�Ҟؤ�{R�uM}���ޔ��V�/���ק^�q������>������M���Dr
�������t��$$2B�_}�ۮ�G>8������������������<�9ʊ�$�����:���
�̿�~o�����߮8�~��������=t�A@A�П�;�UADkY���-U41R��\��׏׷�8�}}}g���׮��<�G
T\�"�ja�"a�NW��,u���"��U����O��q����~������A�>s��rY�Ԍ��Ux�I��P��p��#�X�O��[�����___G�>����=4�u�à���U�$�$� :AGg*�`�9>�w$:��5�����DJ��HUw�w?v�ÞQ�Y	���Y�6e"s�����""�tV̱+-&ʔ�Y�CSY�g��W.(DD�G0"$<����h>� l�d%��"I�$$�Hd4���{��;M���C9���k8i�~/�8�ecZ �m����2�d�f��Ӡ/S��w�����Fq�	�E@�!M@Ü����r>_S̒�ۺ똊Djq��I�_fD�9eI�p�1ԃ��e`^�8(pdE��Ⱥ�u����|�~fr��<��wj#*�"�K�F�IEI��v��pxy��W�5�y�U�7 ����q�i�O��{��c��/+H��R�✱F�eg��B!��G�U�>�	� b⁏�?�B��_AS�?L4����S�6�^x�/�?@zX����nwh�b������%#v�{]���������IW����Vßc�y�a[<�_ o�#��p�S��Xx彩YM�>1�b���y�Y�����F��0У������Pe�t_��SK>�Mp���g`wϚ"ݻ<���^;�f��L��i���
��ۙ'�3o�DG;97A�i���<�?������������	/[js�o�,�l}�}H��$����!{�#�~���`T<�)q4�?9��r�`>�܌�%���T�
�2����=eFj����k��L"��U}N}߻{�o.�aq�)�$_m4��G����g��=�EloJҢ�Ǳ� �y x�
[6\,�B���э�=3���Eiwx]�v��,�{���%�:mu�<�=�k������պ_f�З+jE�Zb��a`�]1<ɴ�s���,��,=���P�ݳ��o]��n=63�`	/S< ��|=ͱR��8��L�������"�f�L6�+�����̆V�M��d���Fmwj�A�ǹҺ���?H�2�v@pe�q��
3�OqkHe9���G��w�4�_�{�w�E�cA�V�2��~0t��2A��X{��&�ai��K�e��5��%��Z�Ly����ŗ��Ɩ�%O��T���h�9%(�=�a�;�MY�~��&�5�^�ź��5B`�h�N�ƃ)��KP��br��th�[uیh�aK�7�b�0s���z׏Z3�6c����d�\�h{�a8��[f����QS�'���.��!ȸ:H6r��!vQL���j.oo�Z�zx�������{\�}О���uY>ϗ��f�F���u���eiðQ��f6����-�[�9���(��_VݘиL^���N��t��ׄ-�W�5=�:f�׸� <H;�+����������{n�ϟ'צ���
��l/F�z�>��:�o�m�TO�Mk?*�������A�@�w��ɾk������Xo^vך(Q�wL�����	l�[�/����}TO�φ�g���ȗ�l�1�[nʖ)_@�&��X��A��'Ͻ����E��ώ��`ځ�|���oM4�ę�s�dk�!4uk�,W�v���gFT\�U��X���*KXUB��!Nokfh����ʅ9DB4��拇j�W{[
�Խo�>귇���Y�}��8���b�WrY�[p�7#wB����wMaI��Nf�7v�?�8Ä+����"p`@���X`@�J� ���_}���$����D[�;g��&�txd�^{1�SM�6|Q�����ci�C�25����-WJ��	.a����oCلsh"'��~ �V����+�edW�C��O��l�����Z쥏����
<�]d�M��!�P�l�av7iR��R����ކGr׿=����q�t;s�`��ݢ�Ü%�a?�.̪D�p��"|u�\CWW���G׸'��ADA�ڐ3��U03=}"X�1��2ļx�ZVV0��nr�E��5����܇|�=O����<��f��<-��[�c�j�w�D�[�<j�h��ͱ�j�L֋�ճv��T a-�3�G�l�fr#�$z��^�f<������='�kߒ��(?5�`q�����p9��ڬ�2.��2vvmnfǯ'���)���k�+ܧK�..���a؅94I����-��B����y:Q�-^�Mc`+����>|zsoX�a�m�����ps83�5�5Cà�6�y�z	}m9
B`cz��6���Уd�������_��.S�w����W/�oOe~A��W�µ���ir���N��QN���u�gb�;�o���h��#9�>��%>>��8������͸1>I��A{.hN+CmV�=nkvzeڣ���~��ξv~��¬2���<B�(���N�����w�}����l�k����e�1qo��c`�Pw���ǉ�;P��aS���t�^dgc�C<�G�_m��B]2OX�Qy6�}������б�Aus��� -< fU���]M��1}�1��^�B���< V�������,�ه[��~��Vφ�l
n��xO��g�d��_�d�,�����O9�ݴ����]�����5˅%M�3v��>�P/C8-��q\��$2-
���N��(.3�5���U����9
��\��[����9��&�e�Y�)��c.'1s�l���͒Ddx��
g���ռK}��&���=zj=[M�䚘P�M���r�S�^��'�۞�b_�k��C	��F���|��1��Ȫ��x2�2��\:/g8��qm��f0��1m8�?�G��X��8��`�&�T<5��r�z\�@�=�m���Њ��d�Ȑ��+�!|ՙI$H�;ҡ��O,���E��L|����\o�!4bj��D���?������|��_|�-l$)���,Ʒ�y��)\�Ża�к�wyf�U09c=2*�%;�St���x#�:l�V��L�ӊ�޽��Y{܆v�y�n�����[@�!��%ƌ�B��bS ����L̾���>��p�)�DL�(\R�Y�/�e9�m�)�)BNe_[7|r��{ã��t 7�]n]�e`25���QE�@�
U�y~�O��Xat�*��r���#�u�_(KQ��s�yO?�5tjQ�M�
 c�ۥuN�$���u�0�?���*u{���\�����[p��{(���A�z������G��tl.z.���spVr�lO]`�b��@bQ�馴�\\��xp��oΧ������ߑဂ��a�άǑP��۾	�^��#��z!�1�L�a^X��Ys�^�c��\��"S�8��]�WPY5zy�c�יּ|GGZ�2^|V�ſo�[;�g�dqR���E���
y�s@�2*���^ܞ����z��=��M�<�6ݺ��_����qE,6�f5��`sϙ�T-R�Q��������=�)�u�H4Bx9ڢx�wn+��ix. �3Ύ��A��z�'�0��~�'�	��a�[�"�u<�<;���2g�BPM���t;��i�I��7!���|_0��?p�~�d��޿=��;���X�(iްLc�`΀��,�����sn�<��� �勼�'$�/��Ce�U��bxo��΋Wx���~u���R�9R�4{�>+��Y5x#���LL/_�t@�9�ݓqW�%RyxԻ����-���Y�����ӄKT���\�x՞���U�1��e��_ᗝ�L��E��%w�q�"�T���"�I��_��y**��%1>y/qa��F��3���l� ��tI�]����� �0�"��Q!��(P��_�}�޿:������:�L�B���?��ä||^1��ظw�q���k�#�	�ޑKy{��W����L���gK{�|!��Th����Y!�C;kswuH����dn"��^"�������2���1��\cə�~��C�3��$೟4=�e���W�UG)`6����S�1��YPD��'g��g�kޱǤ��$�� ��u���Wxm���q�w�{��'Pl[�Exn_�,X��٨o[㸩�!s>1�&�M�	��q���9m����8n`Y�^�� �`�9ᖾ�&|����$��Es���{lX�ٙ6>5B�`�cwA��`���� ri��)�2�={�4]t��e7���m羨L�.�n�%~��l�SCQ��L��9�Ջ55z�N�a���c�= �k�S<���3�Z֨���q��[8K�d�s&|�ʦ��Ƅ�n�vo�/\��.j�"0��H�ǅrN����oi�m��E?`�}t���k�e9����BI9��٨w��O6{[%��t�'X�;��0/�Oz,UG'�yd���؏1�n1_^1�����/&m$�ɴs2\D�դ�(�w��u9�sG�o����GH�k
e���Գ���Pa::�r:��<8�q���pds+k��v��_u�b�ke�K4�qeK�[o��tεwλ�Y��_��D� �¡
�B<Pԑ�u�  ��z͌TU�@mA���NEY|��P��GƇ�X�3�K|¿"=)�[=�T�ETD��E�l���߸�W����z��>{�A�5��^a�^���k눨3y���@z��@~G��X6w>�gП:(2҇��zǉ�}<g�1���kt������E6ť����sbm�3���N?'�8��Uĝ��餼^h| ��@�Г�L��Sk���s#z;x3�8gh���ri�_z5�L�6�D}��W�~�x�w�ضxC���栦p<7�	�j�7��hC/]4ý�dA�y������&�"�R!����S������:�wD%t�uZx�!�tд�	Ogz����d-����}4Æ.ۖY��8���H�$#m�v���M�O�x���+E�6�����<5��ϟ˼���X��)�g)�?BE���ʶ ����B�b3V5��1x�M�6@׏E�,��
e�=��ZVV_�X�)�2����-����Ttb�K�	���hD7�0�-�4xU��Lv��s��m�f�+�� 7:�f�o*7��E��1G��;�V�0~�Yt?'�ݾ/ĸ8e�<�Kw*7��uXU��ꐯX�@ �\>C�oi��EU��5�3U�}���Ү�u\�f��q��\*^�$�h����2w��k��&H�1�s��8Ud� } �(��	d��rA3z7ϟy��~�t����Y�lЛ����ALo<�/v{�P[)y@�0S��>�h�M�e�`0��L�Oj��t9�	��Z��v��Z��yeD6����1�B�og�4�sx^σ��`!*'[#����i�vf���A�c�ImL�u�%��Q0���p᱇&hs�*��
�n�n�Y�h���OC�BM@�-��N	QC�sr��QM6���^�#��0����{�>k�U��D����J��D/zۭ팼�>z��U��>B>|��u��=�mZ�"Gd8a��`��w�vO}�9�����_���6F��X���Gk��{6�;�,�ه�cԹ�/vr��(Sy��ӻHI7(-���2�j���}GU��[L�����(�U��s,͂`��}V��^�y�HoN�L4*ɖx��������jpJ��f�#2�:�bm����"�xz��^��l/ce6 &�wG��#�t�����儻�8W'��`[j�v�E���Գp*�V��},̆��ux�K��=9��@�5��"s�k���-o�|���0G�O_r�K��yիvr������a�vG�r^eq��bӑ\|�D̨���u����&۝uj�����*b���]2(�X�cQY9�a]+qc�s�X��Ӷ$��sQ�N���]��z�����J�}��
w�x#��3�ˡ�Ii�	6�GLD-Ŀ  ��ex�B� y azP!�d��*�s�>u�j�[��n��C��*���&H��S���r~�Ovq�W������{r�|6q�.;��kO`�fvnS�u���K`b�d�k�j|	zʁY�z�!��}0�� �ާ6�P��76`f<ɯ�:��Qݰ�8<A�?�2|`��}� ��;�uE0-���z+��R)���0��'MP�U�{���^�Ɇ�1ݗkG�LSm~���B�=�{a�n��0q���[a�XC���]}hV<�o���`�r�P}6���?�J�~���Gx��*f�f0���d�fX�'�])��o6�E�i��nTn�X���@�Nw��	�����>;qk&��x�ݾ���P�mm��ʳ�O�ak�p�d�Ix-}�@}���W�A�iB0�lw�͖˵δ3��F�K�{1����YC��S��.�Ѽ�.�6���S��cE67�_����,$�t�Z��as9n��1��j�#0$0~	2��ɖW�]�~y}2*�����ܞ���_���Ճ/�O�n��G|C��B%��h��'-B\ky��E�~�7`����}��.�C,OC�Lf��uע�1����
��z���K�!�+vU;X��Wj�"m���;��0�\�jV�^	���ӥ�Q�N]�.��Mw��h�\	�&{-l�yrB��]���ʹ ��0�N�1��T��>��A�W!C�(0�,2���Da�! �������翜�������3u��� �:�'3�t����H�=
��ǒ�H�c�2z�/��y���G�]f����[�T��Oq��x�'7����"�;�Hn���N�̰�1ʝ�B��[QS�4�`d_y�d\�;�Au�.��C8m���s4�Q���s������{�oD&���_`\B��U��C�I;����׽5hxty�ż6:����eD"�|��)n��/��jZ���cݔN[�v�'!���9���LD^���]�WE�(ϰ�k�Y���O�j"�����?~�l�(���l����y���#4	������(y�mt����}��mlH�4��u2�oʭ�;q�}��(��tvw2���{�[�Λ�n�f��^)���c�.��0��p�W���7�ۏ>����u���}��� ���4������x��jŧ���+��Kվ;��=F@��8���S=P���JM������_8!���dw\xkR�v���,��ɟ)Vr�؝5�Qm�O���{���
|ʦ��>g3é&�I6��`\3v�m�pR>۠EL��s)�K;�/7�t��>����:Ds1�;�ݎH�3/�MֹmM3��]]Mwy�rn��^ܲ�cI�;6s��ܻ6�.��㹬l�9R���:ZCK��@,�+�#0�}�7�L���ǯ��V�c��!a��2EE��XS��1���]�Oh��Z ��b�̙\"�P�41s!J���tbެ2S���.���^ڬR�SXj��p�w� /�s(��A�ЧB�C�C
��%��Wp�Ϋ��h����rWև+����pc=@;��K�=�J�;��W4	
�GV\����?u4~\�����S��	�.�2�RN��<�Yak������jhc����B\����f�S�*�����;e����=x�݉Y/<���#�K�̹�����9Ao>W�����	A͝�n�IY!\8[��mԭ���K������wF�G}CU_i ������s��Y3t�̹e�H��9B��Ż��h����s��S>ؐ��4����F3��Cp�©e֦]�ܞb&3-�I=SC�\�s-���c�n�s�e���L��c��c��F7(�������{)W�i��ܯ0�ĥy��y��5<�t�tK��C/$�ySG5�AV��	Ŧ���p[��G�G�2a&)��ŹNn�t��]R�GS�������Ϣ_f)e���Y��NIS^o<���B��yY���ޔ.7dG���:{��"��#v�O1F+.��
�>�i�:p�����U�|s�ގ��I��o�(��ћ�lɼ�ש�՗F�^��7�o*싶�d�o+c�/g.hd[�zB�����y__E
n���Fc�9%L���5v"\������Nx�Gd�]%����!d\���8��n��bB%�N4n0���9v�m�3�o�zN7�s��G�j�T�m<K2��2�u76�%n�bGSK�����:��q���1�ذ%�;j��M��[�d�b�U��K׸�r�f������[j�����&	��R��p	 7!��񵕟B�ZS�C�ju���qu>g�,�(7����
�U��\v�Y��+zZf���&;�ړZP�o`�P�+�t�X��Q�z��^�t*�.�P�4fo
</3n�!����c����ݠn���ց}vڦނ�n�,�h�襓�Giɇ&o۹p�5��#]2]�x·R3�˳)�o/*�>��"�B�o�Xǝ;��6��e�7�����Q�e����!� ����U�TUIvN�4T\�t�x����?}}�����4s�;�ʯT��t���)�� �+��W-k$���R�՘/��[��}o�������o�����o��x�*�(w/��^d]~}{ʞe�3���33�rꏦAr�T_7����}o�}~����}}}}z:��}p�q�Ӵ.W8Dj���E][��O1D�,�b�%>������q����~�����Ί
��:�?�&\�oZUR*�6KB�P�dDE/�׷�_�8�믣��___^=DS'$�H�UEK��D�Ҫ�''<)�V��on�߻�}���}}�������tp�8e�%W%:�U\�'�q�<��I�̮˺����$�F�ӄ�B��+�~���M�
���Yˉ]P+�s�
�H$��L�D��DUʰ�S"9UEF�����8Q?�t��J��Z!�11
*E�\�
4,���ŵ�W������_K|1�ڠ��8�.������z�oEv&k�w'T{Z%Z��b�=$+�w��~ȁ�0+��
��!{
�{���ߟw��c~<^���&��4W8���a��&qs.�tZ�����( -zbq�AȠ�q�����/��,�M�f2�1�&�|�y.�J�v�\����F��g�Z�$F�=vl�]�%�H��@v�0Xb�5{�g�O���Pa����r�:�}�^�<��R����WeR���u�:T����sע���ގvO��f5=e@�u)��E�{X[x3�;�R��_O>����]H��֙*���>����}��@��w�|���<�;z� �����L��m�=ʍ�}ϵ��N�nZ���M1e
5�ϰ�����zix�y�=� �@���G�����H���f��͑� ֭�_%�?0�l�煄� �(o �'����)��V̈vM��7�(,K���De�p�A/ϾBK}� v �i��Xh%�4@ክ;�a��Wy�i{�_Ƕ%���5�㦀�N?�����j��)߲�5�41�����W���iḃ�~��KL>�1�͖��S�t��H��p���t����K�i�l&���'w����-6?}Q�اP�wݱ�>�O����V�㾤��f���L��j����
��y8�
r�w(}g�G	 �4�����qbyF�+^�v�B�}��hu,��7G��ok�gף��S�aћ��:d��*�{��xW���a�d�C����s��)ש��?�7"�7F܉�W��:|5��#k�%��n͚ϟ(�h���>�����&��'~�P��06��[uC>��J�/��Sm��xRœ꘬������^S���<����Z��n�1ki�˞�H�߸,�U������Z�=|��S-�켲Ҳ��0�E=��2��q�f��k��w-=����|�A �}P]7���-tV�ϒ'�r���<�y�˦��׍؝õrh��H��E�,Qٶ%���`g��`T�<DW�-Ƶm��G���q�O)tqf����0Vt�w5S�/v��W)��~hN�_�ա>y���}g��P�+駝LV��T�*Z����0� t�i��N�X�07R�nb�s���|aҞ<�鷵��1P�!��7i�P��9zZ�׊�ig�S��EGx���Q�ii��271�� �Uqu�wZ�d���-�pLW�������c���y��7X���^9^v��:��-�9�0��6Uv�x�z��ákd�Hye���7�a���%���=�a����f�O�g�W�����h�b���!p��Kln�<�u3N�F��H�x��̬=��0���IH���zN��a\��iڼ��<�dm�l�fZKC)s�P�j��Nu�:g�����,�"i99�^AIė:�t��u�uw��)����6�wT'��%�uuB%�ǖuW@�2)r6�r{�{�
��;�㍏�2cd����/$� ���1��P�89�b�ݿ�}ռIN2OI�� �d��'N�z�'����4{X�>y���0bl�5��T�'�Y��]�˽����lbק���7�L�`��_\�\�{�:�h�d�tc���|����.ƞ0ּ=�O��e���W��^SSG儚8~�+�M2a3zbf۔�l<:�r���~�<��<���^�Ag0���*<d���8}Q�`�O}bu@��4��}��]��ͱi�+�S�MG�k&�*dz<�3���^���?m�Fn{���v1V'��2Qd4ּ�]����1,*�/�u��p�h����ϡ���XAӲ�չB���s���s׻Z�9 y���lm1�`�_ԅ�� T�҇�g_�c��ɍ�h�2�����ꢙ'P��.S���;�"�nŰ
k�>p^��ʁv�%�Y��oh{���Ͳ�	���w�3�j&I��|���@>y�O�սB�1�kr>�y}����aS�/�w��/=3L�c�U�zclQ�MR�;�k��
,�r���g(m�3�a#;�mF���I-d�-�ګ�忯e���(�;tǥ��	�������n���6���K)�mὸF,Ϯ�?g֧��#���i*ٔ����%����Ō���J�����>���]�P�Z�2(Q��wo�E� 2��D�paC�N�R�����{�No����=��@	��%�ʏك����TTv�w���X�9�=�1�s/**���Z;g��F��`:9buH��6�w�WP�5��S����e�c5�9��u�>��{��q��n��w�u�����ΑZ��]^�`99z}~ү���X��W�^��������� �9��0_:�zy��B�K^9�Vc��6��u����{���W�%�9Rkj�NyB�Q8�W|���~��m!�$4�d����V�qm��m���a���t'զN=s������V@d�@�����[�}Eg�s�G�.����7ߒ���l"� � Sv�P̛f�}��ُ��_������-	�^]�S�>�/��ڨ7ם����.x�����y1#|��I9��}Ie���W��!���b䗜�Sy�c楠 �G��N?|�▅�c��F�y�^U�i��c��M�vt�mɾ��g��|7%� �k��|��n�lT[H	J�c�-h(������o��&��\n-{����8[�*�&��޳����O-�n��U�YZ���m�/:F�=��Ć�UA���9��fR�g'C<�:U�ˮݾS(:I��Д�}�/naF���X������v�,���T�?a�HnB'E�!�9���˽�������s������X��zt�o��W��Z��v�K�H����3a%=c�����qi[��z*�K8׶8���,v�P)Eۊ�g�L�ď��]�>ӳ�.��J���2�YOz�ƙ��
u��!K��'�>3���3�/�ܻ�ÿ[x�O������/�����*l��D��M��C]8�_�50P���8�hn�lf�dy+ۡ�b�*z�����eSz��u����'9>*�	t��������ib�$<����-��k��Jd��h�rN�Ę��n��+/��hi���f�2�q��6k����$M���ԧX�0'�Hl���3�}��M�sL$���Ѓx�n�0(!?=�	Y��Oa�I��Ob��ڽW'N
��{�Yh�H�z5=BN'��XJK	k\�P�f�q����h�K��jxi�l�ty��suo�>�4�U��f�Y���A����y��4��U�9���S�-�᷼���6�ڇ>|�)��&u�=J��H&����g.dV���:��_�z(�pv;U����Bص'<V.7�r�s&��v`�*���4z�9���@�٤�����;D�X=M��_�WE�|��{~�3l�S��FaΩ&�]f�,��u[�����k_-���a��R�/^=��z�ÀÇ� ��aB�9T�����d �qp��ӏ�>_������D|����Ă�M}�n��L�@��̋���)Je��oj��.:aI�{|�>�&����i��/�~�9'�yPb�*�quq�w�ņ"�����'��Ӧ��*d��9�P�c�4ˍ�ߋh� ��+��9�(�*ͨ���V���P*j,�X�r���lJ���W5���s�=><'�/����[[���f��J����	�&
��*��wx�㫹�ጨ�.�qT�����C���G��ܾ�
���b�M���v���)q`I��
W���o��f�����0�FF&Z�|�:�\y��b���OE��	fX��Sh$����k�'�/��9���=:�6�^����PE��U�9j@���{�L�*oecű�*��:��c�N��]���,����G�����¼�v�k�9aAL�L�L�H��[�����S���C�`Ŵ�=����`�2jj݀�B�rx~�����zU��j�u�z.���qPq��R�9��;`���]G�3������:��ճ��}�0�i�����üH�{;��-��m9Xz��Y�t�u��D����R!�����}v�	����l��ڶ���6�X�9<�K�P�ĵc��A��W󦳾�.M���>��l�\C�òfL��V��펆�8��k`�� ���.2�$�)�c�H�Z���i!M8'�9������$�(z���d�pe9(߿3�K�w�g]��ן}��Y:��%8QP�Ü��Y������ٯ4�\f����kjxw=�vt��u���l �������|�gv��5��U�l��R����Kg������?-�R�B�o8f���;�uX+m�	�N��<�[��wF����X��߽���t5J�������g�@x�Hs��*숗��-�Ͳ����N,��hO�!���8p�_b��}c|�	{���m����M�D�U�tޯ-��kB8�H�|=~!�Xc�~[�@cZ��]�P��%�<�<��ޏDjl��*����_��9�/�^��m�v`4g�gW��y���k�m+���U���D���`H��8-�p�# il�ʸ:�X`&r}L�����3v�}��yml�� Ve���v�c>��?����ފ���r��"V��:�5���n���s{���ř��X2J�6� ���;{�%1��DK�s5�漻Ůn�@�ܦF�Su�Y��������7 �J>���}����Cq���.P��u|D���w�^W�i����>�C6���E�8J��~�F\�R�(T��O:���Xvmf��J+jž��-�a= :]1*�B�F��X��bZ�h�[���f�:��Ca���8)��h�/NL�R���vc��%�ori�9Mέ{�� O �0��C 0�$2��7�� z�{�����	��9!$���&�g���+7�u��+���b��׊knn�i a������HWC��"�Q3���VL5㾺� �)���)�-��m�ma�b�&�9u��g��{�.u��+^Ӗ�4-R��ܩ�Y�P6W3�|g ̛�߾o&�*�VFP̊���cT3���/I�m&�iVn��n��'��4c�DA2y��&�72�9��ߓ�dv˵����N��6�Ȩ��ϒ9b��g��"����D ]xqLl�=��6��9�D>O����4�Sko>�@	�W�t�����6��:����,����f���ޥA�M��3��ü�ހu,�h-e����_��E-5}��@�Q��t�ܟ&��?mIm�*�I���2W��!8s���d�Q&sX+�">�־7ȇo^��}�
����3�uǿU�:j�i^�"�Ev�su�Ũ��N>4|�4�}/�h�ӿMU�S�ePeFtՋ��C��Ɵ	�3��H�?I�!]t&���4W�����\�U�_XN��ߝ�@Q��gw�q|ڱ�VD��!z��D�Y�����F�[�r��+|x�KˋKU�_�/w�.�R�%�a��f��|��W�ͬ��;���a�[���/�S�i:�yA��5M�r���;
&���9�p�s�_a+(C 0�|c��f��<��A�S3P}e�͍��aCӱ�A����C$�	2�M)�ji_����d�^�����,�,���E���+#�J��B|��s��~f��,g���yʖ�YR�����B �����;�:��0�1��B,��~fh�F���'!���3gAwgE>i�����s]�{��c_s�Po���}[y���A/R�R�~`Q�'W�'Y�q�����wsQ�Z
j$�^HAfώ^������s��Y��c
�rAw���)�9N�u��Lf�����0��x�55{��׏/Xh�uXV�����
�YP�o �F�1���ݽ~F�8�;���Y�:f��b�B��a5��l{���ޥ���*���|w���ǘ�n��~�!9:�:X`����=N-��%_a�;�}�2˟��Xz|�Y��������hV�9] ��ܘ^.����kO�9���s�{h�d<��������Qm��u	<b��,�h[�Y]{+sV{R��R���Hk����ꯐ� Z2$Y�.?PE��OONc0�����>��Ԏ6�х�mK�*Z���G�yt��@��o�w҄���n�Z��T�e��Re��K�ysKʁw#T.[�5̱X�%R�'����P��sOJ�7M�r����_�ޥ��T�}�)!��@J��4������??�7��=�=;㯤~��W�g���R������ِ��� ���J��R�n/uT՚��t���ߣ��=��8X@��4�WMΚ�$cX�gJ�����'��>��Y�J�w����a�L���<��U6Ꭼ�`5q���������O��,`����O�;�iE$fG����>��}�.Q���ߐ���<rǪy�������@�1�q�:9oj��J�/�8��b���U�a�[O>��m��r�_'��h��X?�p����[HM�>����xF�Q�_g���a��� �{�р#�]�h^q�LO��Q��/���oRv^�����ޔ_�sc]Q&rzB>��1rL|�y�
��U��~�~m(�}����^.����ʈh)���k�w���z]�SL^zy;�K���V}ᕇTa��RQM�ϱH��������:�L��jT��lٙ�΄����z��>������:��r��|`J^gT�ıo��:Vc�/eL� w��� ܌3*����Ev�ghn�֫�� Y<��;w.t�v9&E\"J#�{��e
3-�:���^�����=ܷ8�6΁7F�"��u���x��K�O,�X�ݡr���7�ʓM⼰���eSnp��V>2��W-�5�g4iOn�.^�z^�#,*;��R�1��쇹o��R�4Z;�chvG���^Ù+A�a�I<���VWv����t��H��;�us��y�uNtQ�{���}-��	������D�+�sF��<��:���T봤���YkpQ�.�.3�j>4\}4u�\|+�J�J�N�홑���`/#y��|�X˥q��y�`��.�[km���M�YW����Z��wPz�w#�}kr�U��$۾��ɀ�*�x��m��r�S���e��n%����į5�9��#˚`�	�d�j�S�r�����(^Mw	l.��f���L7�Q��{��hw���>=�> k��ӭb �*�M�y0�Knu�k��n+��ڇ��f���)u�}��Ǯ�l*��5��e�.��ou�ѰF91����[�f���s��Y�J�]WD%V�,�8gM���R�i�b��2�D��m�w���}��h��:Q��Cy�O3��=�]��$��e����r�ߢ��o�&4��˪Ve��A�ңj����#HX6GVh�zh܊;������̨NU]䔭&�Nell"�e�-2��*��.� �/�r���E�*�Щ*�.�S�̢�y�t�i�Uɖ9�]��c���L�9x�fP�{��4�qMר��� �	��B���@�U-��״	�[�w)H�te��S�kԡ��.	�9�ev��#[{d�uCHi�W��>R��1����L�gm��ݝM��G�6�V�p�����;2Q��w�g���Nٝ�z8�_Y��5�)_owp�Vͻ�]�x�}��V[c��������!a�I�uM6����硃���c(��!�:�*ƍX���+�����n{;twU�8nv�[�v��5^EP���1�7�\qʾ�ǫ����9C��Gx�n�&o�[Jΰ�9m��05ȳ����&�}��]SO\��2-�<�\ELg/���$�˹�dR�+-U�q���S�Cv����Z���x�+v�oD@�V���ƞq�jxe���)���H-�l낧sq�����Ռpʭ��l3L헒��8��H�;��OR�Q���S!sZ�+;�S���NM�:��ڛ�s���Ku�:�= 켃��|d��z��#�+5�U��6��#ۖ�R.[jV˂7'cic��=*fث��U�K/�D�knl*.,�ce��Sf�Z��KJ��ief����	#N&Q�*ܢ��q��T(�Q�H��c�"�K&��-FJp*T�-�%�a7"��tB�wn0�Pi��� ��.+�P(�9�R��YY�]�]�!Xb�%�D���$�QhE� �=�z������������_M�
��4�$D4%Ǜ���(�U�oOOo�����_w�M�|�7�p�[���Y�Br��F~�?�x���
�1-qdr9��v���o�?u��������K6��wO$�Q�S�I�0���"*�$�ÕW�oOOo�q��������|�7"ti��H���k.P\�$����	R���.s�O��ߎ8����������{;�@p*|��ET�MwÞ��L�]dh�|�����~8��믯�___^���9¥C퇖����s��%�w��� �f�o�OOn�\q��������ם%�ϱ�B�*)}2��I����
�QE�ȮDG�β���DQG+��8\�9W*#̪"9CٕD9!��)g(�3���
J�^�����|�9r�!���UQ^���6�U˅&{�����(��%B(��u�S��G�G��&�h�\M�����Tf��7^�_uC�KDt��2_^�ܳ͝iGkF\guu9φMw:yC���̩t�-��N����42�̺'������^��C����;�wfkǣ����Oz������&��-�C':��C�"� �gTpa{u�B�)Q��4�p �oM����Tl��Uc�0*�G��,w���f)�19b��j�Z�������ͦ3]���Î5#+���N<+<3���T�p^=�\/1����:����`�km��?!|fTמ���U�8�xͶS���o���pq�PW��d<O+}��M�m����ʄm��K�Z~n
౮R���Tn�!;e�y��ork=R�S;����[�g�55h^c<޻�hG]�߱���#u��������AF�<f�ò��n����{����mewS-�`CX���lPS�i�0�Z#oO�7s�����؆�#C0#-y�TR�L�$R���ѳ��~��~G��c{����G'��S�v����4�l��W��s�A�q�e���}C�r{���i����j���ϱ<����qmg;l޳ւ4J4b
���c�S��b��r�m����H�g�� k>��g�q�R5cI=wr��[��Ը�:���{�{�HN�6:��0�j]� ��0���������:�Ƭ�<4�|�����8��w{�����:&e�����%�Wb�6�i<�x��=�6;�,hy�r���rJ��x�����|��������Ď����,FyKnwg�Q��	�!6�%��Y�2-L���`ed!���7���F���Rm���#���t�	�އ�>����z5��ia%d>']M�(%���Ǻ�Nܸ^+d"c���v69����o�K��hUΫ#�z�
o]Az�f���>�h��~Z�&�>�oSǯ�T%>IN���rÏY)��O�K�og�\�	-�s3���KWj؈^פ��MYa{�U;��Ќw�X�_|��nC��,NMn��9�Mg���Xܻr�Vlƙ�u�	</1R���A��?�eҙW!�nԧ����Y舸D�W-b�n9����,�S��Ɲ�V}0ȇ�x���z�o����{�7��-w�J}���wpέ��(�q@���,|���Y�j�V0��Qr�Ǫ|�l0����� �Q��_6��t/�f�P���ږvq<�S�确9�Y�M�=�	�ֲF��M{�#�yV������9�u��gbRrɦ���E�;0���Ȩ1ѭ�����K�)���R��a��P������`��y�ເ7���5y=��i��Ǧi����Be_��<���5��c�.�탾@�����S�POd�\�3��c�뼥0��)Z����-�p�W]�ø��:v,�i㝗���0���޽�v��Y w[� ��꾡��q�vѭ�c|��ξu�|����@��!��0���� ��g�&��Ͻ�Z�Q�`�gQ�	��dA����G���~�FZM"�}����P�v�4C3r{�����QˣK�ˮ=>���r���gwm��f�3�匸䣵z/_�u�ϛ��W��N�^^�Ŝ�L��C���O��c�v~毉`�OY[�:E��Z1�h��5��| ǒΑ���(P�{�X�%�x�~�f���s�qA獺�a�W����=S���b"�E$ �ἥ��V�@�t�\h��|��yѺ姾T<��|�f��9��ɥ�c÷�k�旫���	�é�N8����Z=8�8ݎ���L��6�^�mn1�,M�&{�dvjy��cFv��K=��əHQ˝�����_"�m��Z�!�EE�6�m-�6[�b���y{I_=��Bs���qp�?zJ���z�'m��؊���&�K&���8r�[<~� �R,�/��E�ѱCo�����%�R�f���,�]/��ѷ@���
�M{�Lq����ᵴ5(�Bf~�l��V9�����=��:c��tk��k���e�b=z;ï���As[�xK5�Ҁ�����R����1��>����"��wF�ʧ��T���y�a�(q:(p�;ՙ��͕�cZC.�Y�x�����KU��<�뛧�>G���+�0���w+�!�̻���z�����C}�o��1l�`XȂ_-G�uz���j~��><��ʢ���iը���Y�: &kq9�q��t�"�<��s$�_����<����2̢iO+���yWoG��I�{Lf�<���u(V_<����d�'��!�_Ja;0[y�����n�Q�r��_uJ�c���>�ڠ��we��5k�����|�s��q�m.��\.�)�r�^.�<��L��߸���ԟC	b|ПsW�Ss�z��)���-�ԹPk��0�HqT*�����\_�`�0�RK�b�,'؅εf�������%��>�m&m^:��O��� 7�b*��GG��c�O�cTƘ����Z�l�S�؍����pi�g`S��^7�q�9o�E��+����]�^���{g�ϛ5٦]�7�����С�nv�d��t�~hńX6{/��"������c�k���כ��~O�}:b� 0��{9!a0�`o��!��U���Gb(w(����ptǏ����vh��%�{.��{��"O��q�'A2��M�C*��N�+Wq�1��i5���W�&2��c������p_��6�1��U�=���HBŹ�K����a	���ca��۴����P1���I����!��63��K,��n@�p
�kl�	#!�!���?n�p� r*�_o|=r��a�Ƒ(��a0M�O�ɟ�KK�|����lzK.��u4Bg(zDk�����rQ6�\ �Jz�2��^�=�v,���h�wH-���H��g+���P_� Ep��cM��t)ƵLi���ң�o�@������rŝ�h�#MDC���i�{��S����)glbv7��*�@f�P���~������oM Mcx�K2ŐS�S�S����|���N�%G���z���q����g�ۀ̱��*9;�ȫbw��InӸ±���\��uQN��ԋz0������ך��h��'�cCn>)�V���ڢ��l�l�;��������,�^"����=>�R��Ao�>+�3�V�!&�����`�b��G����Z�Q��T��G4�o�����j���ɵϟ��W�vgxA��[e}KR&������
����	��S�ؾ�L`cs����^Z��p�7պq����bN-��,6���a6��6�;榫]6������9��P�Ј���1�:�}��V�t�T�*փ�!�w�R�e�NR���Y�)�gku����ó}�-�m��B>�ӿR2��x�;����r)�n����f�Yg����cN:�b�qՕ6f��vi�����5�®�s��;�#����x�����d!� �����<G9ǹ��d}��X?��𱿙/SފwMR���y�4ՉH�|n\W��W\J�w���Lj��/j�	��̢9�t���@z�|�R��*�@|�����'{,��+v%MD�W�F����ݻ���q�'Msp�
@��;Ϣ"����a�����7Ck��4%��gZ�� `SsK�Ӱ�d�Z�b(0��G0�p|� /�˞/~����wn�7��̔���zפm�@M����4���+��:i�1B�{c���o|Gʴ�a6�టAeY	�&1��{�E�;E񐘆�a��o\��{R��w�r�5��B�1}9��u��D$}Hϡy�bj�أ8�����ʥ��|���$��� ������O�[�Zˡ3��ɻ)1ԡ�9oP�Ϟ�fI�]\5�P�az��;��%�[$<�4?-���'\y�47o\�䲫��1M��H�~q�6���	=B�C�Zb��~�!��7�]z�v��>���_��#]9�v
�hi��e���.�M���������_��O�6~�Ч�Qf$~��!�p����Y�B��o���ك1Rv��t
��6���֏�%�1D#]|P�V�'��Ժ�V�P2���jy&�ŵy.t�Nt+rǖ�˽�ۤ��cWs1�-8��X��������9�0���ex!�0 m#b�y�*����q�݃~���i�������f�%�l5�����F��=��D�ɉ8�A���5�dI�p2��"�5�E��3@I/Qno&8����i
��m�س��&M<���%F��e���ԅp{`�DkKp`��,�ɇmk�fŁs���o"��3���՘�eb*��ouqq���Ú��<��{�<�j��F�ׅ�&M�jÝ"Ħx���O�m�H���0}��\�h{-�Wo��=�)��������NZr󕌮��
i�8ҬtXR����gg�C��O=�R�OS�D�,� ��<�>7ȇ�;��6��G�J�;fkq����T�΋��;��\l�$ִ�b�Ř0�f�`�����꘳�s�Hw��((�
x�G��!��_VP�k�yѬA�D����N{��;w|U�|/+a4P��R2�f���������?��Ą�A>x�-�1S��fx��I-�}�(��v����|�FF��^�*�/����C|�M��F���j�eb���;������|��TUt�����6&u=�3o��ܶ�#��u�غ�K�dT��u/����)0]ncPBH��)q�v-$k7.�c��4"�.��R�]gS�<]��Xk@r۽ӷ�J]�n*��_��8P�X`|�2��rU�z����������S�]�8��S^��ߟx�S�q_�����m�5������^6�8����x��A��}��iC�B\B�5�]�6�t�*�,�n����csyBp�}�W����|V�D���W�t �A:n��]
�W@k
l5�P��7'�Ƭt����b�j@tby��ׁ-4�����p����y�P�E�;j�w`Sv�C��/�ճ7��\�U��"k�Ś^���`hȂ_/�=˨Y�ko&Yw"��x�;]R�V��jٕ���b��q���:h5��-��B=�.�):���
זZ�x7�������Զ�<��q��N>�'//>�.����Z�ͮ?� >���B���z�����\��:�uܖVc��O�p/�h��ꮨ�����|	�aeb�.�b�C)�����j�������٧����g�:u'al���Jc\���O�꒫Y���*��׭��qX�<���6o7�-�{ichSُ`���U�{	{\��dKr��*����%=�(����#�ך��^lZ�E�	�}�h�]�AT�94.��⮺E}�g%��t�n;��߾Jv���޾�:mt�$}׺�K�|^��r�7�g��-%���󵶟[��Ǭf`}��B��"�P|d�Bp	�%*���p�@C!�/|	N�00ʯ�_#��G�,�����Sb��p��(^���9<C��C��\�l�zF�T2�O>B��5iT9���5��0mj���1ڪW�Ҙ6�����	�y�H}l�4�,W�|���F}���V�4�/��j�":1V�
��^�"GP�����޸(�52~VE�Vv�xIK=�nmz
�j���/��Ca�s2��LHw�g���5g"}Q.e��0�W�iο|��L��Y갡��y���?�z,0%�Y3�W2��W���:�.pXzC�����z��S�XUh%m�&�\�.���X�_�3�+\)�:��e�v�<n�}���e��V��X���dn=K�j�
�^sPS
��8|P)��]o���<�'v�!ށ��ݞ5�4�v�w�N���-�h�kW��sO�3vF���&}�&��p4�p���:��A
'{�=��0�������mA�����V�1�����j�����X�u������1�\��:輲�M�a^*/&�<�vk���\���6,�j���<
��m^o���|#��3p=��,�3�Y��2?*l�W���\~3-���땳4%�u*n���)�D�x8U!DW�q��Tc�=���������}��u��B<�'k
"x1E��Q�;�j<"�;x��>����EH{H�� Ä�8@�������$20�	������'�E�m����)���J�3Ǧ�#��,��*��NE�����Z4*�b7��eǤ<����P���>�O~������8v�zh�s�h͚��d`�s(0��9���Y�K�6Η�� �*���z�w���'N���\)���[1$hn`W<z�M�u9�}��D���-V�%�8��l`S͇*��Cs�{�a�7l���C5����>w���
����ر�����K�ذ���5:c�J4k��K"a߹�\߾�Xs}��g��߹=<{�1���Ѭt���!��,i�*�_(�����~���Vś&ꫝ���gb ;��Z^��?�Ռ?�z��d'M�`%\V�_?{�Xc�~^FI_zZ�Vb�ު׺�d\4٦ �½��K�^�.`�tNٗh�8  ����YI�����׭o>����Yv�Y��D!7
Xa��c���V�z������`��A1�1�eɂ�b�Qæ	;O��S��9�<���*s~�a�����N_+]��b��A��/:�i&�C��{� IfF�ƙ[O��P9읚�ȜJ�����:ʫŽ�Q��].x�Ҷ�b�!Yh!�Pv����ޖ�4�u���9�Cw���['ڵ9y��{wҕu<r(#���b�
�/(��w8�|E"��X�v�t^� �a�@y>�R��D9D�{��n�,���Ep�St��b�rW��m>RB��UM�O�w������YPXK�!ZՃ%q�4f���m���v槎���c%J�������9X�j����%I���z��XY[%�ڒ� ����͢��Y��mX����a7�Z���ZaS��u���۽���S�{p��>�H�۬����F.<U��5ݓ�0`���y�
_!C�9U��Lj�����H9c'C��!OL~�C�+�v��կ*3U%)������(�Y`��=�i�Fk�|IF��];h*7�Rڴzb�[<�Ua�Ŭ���pfi��^��u1"���u�+���ˡ�lj�[ҥJ���ln����<�gj�p�3skF��T�&-��EGF�\�h:y,��5��B+�M�}�Ĝ�J�Zn�IN�w)b���oNk娠�P�&Q�㳙�ñM��M#�R΢��Wdd4�Ie�����C9�,��=�]U���d���[Θ�5u�#�����H�r��<0�=C�(QCAG�N���B�D��,��ז� � ��yvH�^<�$�w��nQ��T(G(�K5˿3y�> A)�G��N�i��:��7��	szxC֟Z��K��BBd/g&>�W��Y�KJ�nnˍ�7�%�Բ�Վ:a�P���7���-Y�����qo���+���g��[Wa	y�9��؊�q�������G.�w��� �掱��ykDRh)��}�9��VG�u3��9{S;�÷��3���[L,�:�Uֹ&U�ܼ��N.β=���uNI5�T��W����J�#�e^����ح:_A��o�Ц�c9��%�(n�Xj�����X;o���C*cv�*z�@.��X^c��w��WHi�1X{ֻ�*"��w@�˴�+�0��� r����՚��hu�T�o;�gjuq�yEEF���	��y���[r��0�BѲ1���Q�A��-����㸦����]Z[��?;N�IM!2�
n����3����l޵�q�*,�U|0H�]��s-w]L�pDS����>���gf�m#��{���Wg�y�qŷVFS��p,��&�i��j}�e!�
�;Y&n���wUvHW�t�� n��e��+���U���A���jh�5�^���A��T(
�Q����v\�}����"<��O��\�����ߏ��}}}q����נ��
��.�Z"b&r�:�W�)D*+�r�j�}x�����_���0�����쪖Hp�:\�4���s����"�M���kv���?__\a����뮮Q�q&�4}��93�UU�LG����Ȋ��ϯ�߮������>����GME��Q
����We)�)D(���K���淞��8�����>������8K��rBDB�r���$TAp�_6��^�7������{�z����>����t}�"�����|��[h�XdE+N]�Ð���sZ�g(� ��3�(H�Qg�V���r"�ݡ:�5J*�$�9P�QQ�uk.]Q�@TL����G����8U�YY$��~�(".D𥉉���kz�K1t�ۨ�.�3��9Ns�<Sb����[��M	w��&����@�F`!��^�����Ż��'�'�L��:��Q�v�yP��S��Ͻ8�t�2W����;S����e������'Xo��Y��n�J�X��X�؆�1�+���[;&��l��E�,u����MwT�1(t��Z��P���rD����� �n��| ��4��jnP��znb�O�S�z�O�xb����Uެ�>vQ�H�p����,����F�������:�H�#��A5߇�]������ƈP��'-��f��YX�Z�������>Q�酕kf� y��s���Oix���\K���μE"�k� ��sY����AI��x�0ϐ7��i����8h��C3&xi�@��i~�J+���Mj��.�Pv:��IESF��̖7��v��m^�v�>�	�f5"��#�����R�z~a���F�V�z����8�V�WS�ieݲX�1�eCz:� ��XJ����X �S��(t�)�h~}|jf�ns��C�7�~V��ʯݜ�y��`�5K��N�3b'����?#���*��~��wsE����wKHz��l���c{0�]|��z%eܘj�P���M�`u5��Nm��#����}�PK�=�we����^!�����J�r:V]�(���G}7�B�y;� ,��3z~�{�0��^���&�}? �I�@�7_�/��kX|�az����� � 3fn���'�V#�_^�Gb��D3\@P[����PگfӒ��έ��T)]��4$�i���a<Zf7�����0��)�oAu�T�S�fo���>#�,�-^�M����	�c��/����e��a����ڮ{W7N�F"j�TK>(t��g��K;��`y�x@��jm����TŪ-����yO�I��~���|��K�|�;��OQ�c!*���qmC.������t��-��̵靴c�pk��X���|�)�q!_��S�#���U}p0F�7�Q!��ru&���H۠^�y`*�v���v�V��pѿ[ml�Ǝ�f�/�����5ѓ�zc�Q-X�E�Q�斐)�v=k�sB�W������±<�&b�6��׉�rh��{j-����q2�Af������K�q�:�ش�b)���AH�'�����ɩz��5��o6Ҍl�M�p|�g���e�y�
yn�i+*���ќ�g��N�w��e����n�p�e�{ʅ�эP�4[����Y_S�s�"�+lUa�H��l�	�#.�W�O���Zby`�#���L�vG�9TwJ�r�jtҖ%]��_��澺��A$��+����"j
%�1�����J@���rÿ��4���Rw^���,������W�ضg?���퍸�9�V�	�q�0�p�kA�������]���0��Ovg�7������{�2���Ԕ�q^��|�'��S��uCN����0i�k���JH�t�q�{���S�(cY+�H`~�V@���Ļ�4<'%���O�3�?n\����/W���#nw�Zw�Q�G7��XJ}� ֠35�X.����R0e2���]�:����f��3^���Kd�zF%"�ے'��8��^*�1�ѸGU�>��C� �kzR���Dt�ۇˋ8�x`X���]B_��3l�8�oKc�K��<�.��1Ü�CI��<j������a��i��k��> [P/'��&�2�坞��@�C(�/�_��NRB��+�I����[��B�(��3�~����B���.��tF��(�_�������1�N��1��d��=���3k%Ki��MH�/*����,9�������P�F��a��cP���UI����?�i�ix�W��6�:���9`�]�O%���+�����-|��1
�,2 ���/�R�s����X��o)��#ũ�u���r�3���
�%꠳�9Sm�;8����@�+��C�=̮��,������ϟ5#f�����y������XΑ=�#�s��}��ne�G�2MT4U32ۚ���8��N��;,Ꮸd���+�P��1�K�=����ל�g��P��0t;)}������-�^Ô*�n�]�|�諔�!DD��!����������g�@�.�ϵ*���@�CfX���6��N0�&�f4ԋ�d�m�3�z|�6�`f���*/6��aa���<�4L4s�v�I��=yb�n���2�k�F2�,.�������WwcgL�+:d��3�L�K��p/M�����IRq���v�q�uhk��xS����^�N��Y019	$Ϲ��3�����}4���_ɯ]��r^s#u�(ƿ1��4fH���Z�t ��׌a����m	�/�[�G0vxfxe���9��%��u�(w�Ρ���\�)=GK�� �����fq�0hNoϺ�)���x@�͕��]��	���8`��.�����i�*o��~1��B�#hߘ��P��"��g�)�U�����T�L����i��7�I�]��7+t �E�B����(�y�ys�cEp���^ij�r�g����i�F;��
=d��[U�v��^�D�=M%�����z�*.���<*q�|�b�c�(J)N��('M�&���6��-��n@}�mq�뇦���k�q"q��"k��"�������q�ߍ�~l+D�x�}��}9�����"[�����<g<��I���P[V38�l/�#�:6�vB,�,��>9h��|$��@�3��t<^� zi�j/+�/.�Ӳ����^�}>���/�}�fN�>)��c UY[ݕ���Q�@���R�����Ly��u�B�@���2j������n�z�e>7�bbj������S��,�v��i�J]oݕ�]Dh��.�*�ddNo��5M�y�8P1ꫯRxvu���F�0�7��������mXt�)�l��M����5�7O������$�<�W��Q6n��	t�}���Gc!Ũ�B�XJU�᦭�]1�ւ�lϛ�)�z�9/�pg�vJ_�F$.��s�W�+?��`j�k歄Z�o	��2q�s-�4-Pu�Ս�W.�hc���i�[������>��XjQ���55ljIN�5�'�9�>e��>Dp{�^=���/1/0���~��^���$|�K�-��緶�;cB�g�X���ۮ��6�����W!�}D8{=<�������C�����ԯf@W�*jA� SZv��6���ޱ���� жd}<+p��U���O
�P��n�Q��~_�ՄD�.�wD}G��_������	�ـ�Vv���+X�����O]��nZ�}��)%�*k�C�iwI�G�;��	�91�Wi��{]��6�9?hjr�I���;��/K_�餵�	ef�_��X��\k�<%�!�5�B�i0���w��&��]�F3�4�p�p;h��L�M{��6�7t�[�(n0��W���Ӄ��k���`����`\xjLOt=���-��}n��.�5��J'�����tl����F�x��+}��H��/�z�s���	X�u\@���h��+�|�B���sy��m���91���x+.q�0g�bU���xf7 �3Y�)�v)�������.�AM�t��im~o`���4l�M�h���#B�w)^|-�˸U�_m�F�<.�hg� ����ߘ��蘊���;bZ���l]N�{ud<��Z�s��t���E����[��`�WK؝,@�!k���:�(b���*v�0���%e��$\���Uy���[e'�g�}�Mcm�n�l� n���0�Fr���I8ۍ�B�[���P)��8`�\E�N�h� E�ݠdr*�����ba]6�d�a�x�JFဨ�x��'�g��;|���=�o�ᆝ�#�5�h!����v���x���u���q���� `��D���Q�1��6o6I�ɾ�#�e�@��sB.-,���=я�nM��8�M��S5�0�F^w�2}ݞ������W!��
��eۊ�ŵ㻸�~��^^�+k��Wm�L�OT�z��K���j`B��B�~�U01���LsgREou�R�H��:l��8��S���;P��j�u��w��u�ڳzU��S�;��7H5�L2�v#�P׽F��z׈�נ�F�`��}�5ve�����Iš9�ߧo�ʺ׋���z� ��>5w��z\�yZ=��]�����}Պ�vzup�~���h�x�戵�����*�g�������a>k�&��k�X�U���:1��D�}�&�s��zi���:=�vS�wr����l�~uY�Xʮ��h��Uݧ)S�F�@� *���hI����T���֯��}}���Gs�v���0T�,��b�$��yjs�B��YГ���e׼����FF�Sf��{�,=ѻ��[&I�n��v�Dn��t6{%�oG�+ˠ,5KoXOǚ��۸3/o6z#֙VKoF�t�� H.F;u�/�hs���6��1b�kZ��z�ƪ|���c�4P��^,grD��
��񼆸A"1K�����cL�rB0�Ϣn�����x�Ȉ�1��u�S#�9~���{D1��/�â7�a�v{���3+�]�[���On�B1��r-�:̌�V]��x�jT���9W>MHGj���qc�ٓ�wg�<�D����{���ԁ$"�
�N �=�N���&mS���]�T�JOW���uM���g	1��^�� Mt�7h�|���]L�f}G��PYސ�.gdVt�%/�@;.�{��y%^�'��[���}��g��#V�8Yp��s/׬�"KXȘf`����<�"���1��[��5� ���Y�W%����k5�ܥ�a|� ��1`�wy��\��ʂ�Kڏi�_3�Dޏ��Yޫ����"X��r�4��̗���[�´-����xz��I��h��uv_c�ͤ�S�w�{�nk�e�� C��x8����f�4#-�eYPc��|�M���"�9�^]+��<6
����O^�����;f&�?@~͐�`T)7$��	�*�bYu�;�az��xXf�>��H䈅���s�/M\5mS4U��wo?n�5�Y��~T��Ӟ�m��6�Q��L�K�q������Cfcw\�s0�0�P���1��'�ٽ}�+����:��q��������M�����Fr����s���dl���E>�Py���C]-��Y�*�J�V�N?�d�{���1yX�����i/zOkI��j��p�D$�TU��j�D�1.���;��}=��Uy��9��������ʩ� W3j��sk��
e��'�1�33��0�.���o��l!��iMX*pG,��$�P�����WJ��R���V�u��ieͫw��-���[�ܴR�=çnV� 6U�6�c�̥K�V���"�9er�e���ܮ��T���ݧ#�{�$[�6iӷ��,�(�GʭJz�����Ux	5P^�:8Щ�oJ����|�"^���>�4��t�Q�������y�նo\�0�
�_'���d�'B*�� 	��g>b���{
�\<ᲈ�x�D�������Z��)�E�{־�&����nY˪�A�EIl���U�����"_��TmT��Xc��7����[#Qg�f5������Y=[��{��6�0T@����="8@�����[�Cy�Yݎ�S��j*p��	-�\�Sk����z�!���c��E�{Ƌ6u�ʳX��Q;��~PVH�g^��4
K�b�2�~����}-�˽31@f���"�����c6�}�_pD�������I�M����鄛�>�0&gL"���i����ҕ�x�_nqܘ�jaG�����w� ɻV�1�����t�{� 5��a;G�߲+�P$�jv�\��T*�˓�f�qW7����lLYw�Vb�g8Г�����)�iء��M'��<gJr�z�v�W�qƬ���k^�,�qݾ��d�Ӵ����Of$�5|I����V<�m��4�1k+�/F�K���(	�˴�t�fG���j�=�t�	��XИ�"ə�ȴPrB��oBNn�4V�V�X���^���%Z�V�r�����hF{�u�LN�81Enq���W��M��|8&��=�N>�x�E�*�m�ێ�2��8���g>c�L-
��f�Y�WOE+�66�h��%:u�&���[w�n.�ڱZ8���>b�@��[6��x�viC�]YL���y�g��6�p���F;	tS�9�j�o���WK�bI���Ӳob�g�b��XF���KA�RZ�<#�K�3��Zrm��Ҝ�%+K��s��#�Ҳ�C�$m���X*J�{,���{^����3e����m���􋾶�9�'a}˄���ɘ�D�$��j�Y9��+)&�u»��+,��;l�wR���8%ѣ����Y�u���!�HɄN�2nN�
�t���J�'TX�SzURM�8.tǙO�c���ɭ���W�c��iȲ�.�aނc/��f��t}k4�؛Y��dh=�#�a�P�|�Ċ(b�ӗR�M�'tAW���١$
PKʅ�`%�f0ub�g�e�m�50U I�WN�mA�u�E��bJuG���I�PS�2��c����@��\�`E�n��rU*�g*3���#�����A���w:���j���Q%�3����n¨��[��ƴÆ,&ftzCT��=�y��wZN���^G*�>+nB���]xubOEKKe̻�]�HwQ���t�+,�'c�%�`�C����")^�T�wj+���m,�C1n��	�K][��̓����Vw�t�.G,�7wU�ޚ.���(��tU�>ܝ�։G�S��ֻ���)����������s*X�L���iĕR�E�u�v4]1��~ٝk���ۛy�Z�I@Ȧ�wVEpyM�3��S2r�-k_Z�\�l��F�k�	��̀R��-\2�vw+_e��qe^��x���=�+|E,�tvoi�3H�	�H}*�R�G��X��M���u�*���%:�1Jٖ�*?e��{#6�2*�f�׹�F۵o�[�F/��γ�ؑ��%>���ٚ��V�K��`��ݎ�5'	�t6�8�I k�s��>�q|X��+C����s��g�N�x��E��䳴�`�k��uz��m�,��wƨ��h���:'S]������Q����H4䇅������FdA�0�r�\H�0������ �)�,L.Qm$I!Q�U&Iȏ�2\�bUjE$)9A1����իa�6�\m�@1�.�;$�d�7y<��'s[�{z��\U�"�����o���p�OC4*��'=.'4TeÐg��9�%`Us��7Oon?�8�������__^���ys��T�Qe"%�:�&)9ro�2��UMP^��������믯o������rz�y]�xAp���˔q׸bw�l���"�9�s"�+0��
\��9�=�=��>���������>�!x�TO���9��A�l�8Y�G ���aE�6O>s�eȠ�dk�;�o����}u�����__]|N�$"�y�9Qʡ+W.s
�(�:p�W-����Zݾ�����������__^wID���)�E��!E�"�Ar��(�$�s&�s��EJ�����n�[��|�7��{|�3�o����)Ց�y!z*��t�)�����UAz��L�C���"��(<����U�*T����TDUq�eG+�ّQpt�d�IXTu,�UA_��DE�%�s�����A9�eEQ�$*��D�QE>���ʨ�����$):�?>ϳ�����Ͼ���T�*AB �R�Q�����*f��e
e�*�/�2�ZO:��eHm�6�.��^M�l��r�B��,/N��jWR�z�BI�+��5P�4n�hD$�Ӆ�5A�޽�rMp�ǽ���;���y�9�O��5
A�.$��P�p�S.�%�H�{��;a��it�XE�KM6�"Ԉ?���s�,zO�/O�R�����-v������Q�_q�~�~���/q�����}�`�� d���+�b�X�tn)���M����:_�p�ׄgK�,�Ѿ�֮��N�e�v�'���YE�4e�Z�s��P�_�}����쮈���0�ʏ<����x�f0&~O�����������y�z�t�L-q|��A���K�ͮ͜�h��D7z�CR�&<U��8XG��4y�6Bf~Z �#��J��}wS��1�q+����׭�qÇ��6�b�����Ok�T�����/%�ޠ�Nq��<k��S�O���]h&��`!?�.M߼��	�2��n�~)]�W1A�97�E,�y��y�ы5�����mg%��)J;�=6TC1uq�O��>�f~�w�Sw]�#��Ku9��&�6���v
���_�_K���}�\�^�h_��T�-e��>F�粻Hpt��(�u��/����V+��(����t�
2�/��#��[}r�ˆ��z��뽉�+]Z������x3�Ѻ	�Ba�Uk�zJ*��4"V*�+ܞ���*�m{K�wd�s!@��S��h�.L�0��;����4o�D{��+��3��䴍jU+<�-[�5c�}�l-������!@{�-��`�����M[˲:�G�UH�k��������&<�=�5X51��{�q�w��ﳿK|�~���{Ͳ�1�;,sD
��w'�zz�awL^v�Ԙ[s00Xgv���9 ����k�n3�o��%��Lڹ30$���<D>0�Fa��6-@q����Z�^"��8;�ꃠ�s<�b;E*�0s6<��S^S|k׾��Fmp���v���f{���7WXӮ�x��ߧ$1���\��*EVǒp,�>E��D��4�~Sդ��Y{N�k
g�N�y��`�5Czi^����H|��1s{�a���:F������e�JN-����U�l[9PҫF�X�
<jN�G�*Ӏ{�neX�6��M�	�kv6~�$��T��mLYF�uW2t�.�!	�^r�ZZ�sΊU%�a[��-�mշu�k�7D	x�9�8G4 �泜k�x�v,�+j��kз����U�F�@}�U���M��#ŏ�6b;oraW�Q�ESϧ���e�L��2��V��MU�i��A��c�` ��u6��l�q���jLgD���s�'����m�$�FhrZ��h�X�%^ҍ��m��q;�`Y<7u�_dK�DĈ#��P���/>6��׆I��+���l�����Q-�\����&�������ق���={,���@�����A�q�"Xsy�y�l�R�І����������0;[��� �o���~hR9�N��I�U�ӗ"�{����x�W�{ٹ��kC1�1sV�񹫿k�nM�����n�������H)Ϯ�3R�i����U�U�^���0O�7�{H�x��9���U�"^�I���b^�nY��NUͽ���������n�'�2�ȷC�Q�����h��Ǚ���9
�[?��XV}���/'��;Lߵ���z���]m�R*���7��k�ćot��,w��9�	v����_��Y�a9S��K=��ve\��3���:�j�����-Һ�;M�R^w�סS\��ʟo��~t�X��!�.k��z-�}kw���o���pc}l��6��9��88�z9r
��������O6�C��ѝ��]nt���fZff]�Fz56�e�/YETT3_Sțƅ(�V�7RB}=��h#�gj#0�Ǯ���:�5.��ӱ|ĵ/'RoG�tE�kD��ܨN�M"�+��V��A��]�^ͭ��;�u�H��6�<��ޏMǯ�/���Ba�j���5Z�ƞdI����ܐ�p��c��]�E�=h�>d�����]�V\��<�\g��LT�v�՟GR����q��}��e�(�ފ~a1�����:a��ѯ��2w�{ ��#֨:�g M����S	��wt�r�E�*Wf�*�M<Q��+�!:��;]�{[y2��{F��~ d��(�i�8W9�pV���.�^*���,���Q�A�e�&�w#"����ڶ���:��S���[�G�w�z�����_�U��Rsfs%��6t��3n��II�ޯr=䫋��p�{޿�0~��� �����,�?h�i�R)ho^�������*&�ʔǟ���8���2�Ci�&n� ��`���Wt�վ��q�u��䱪dߛ[15AE�5��p�h�=ٮjt��ݳ�j1�
�} b+)�U���o�&,m�sX�M��J\v�奄�o5���/��6�a�f&ݦ�b��=��l6�Aq���aaz� >^�*�w�/���?����g{S߻W�O�ϸM�/I���v����.wV^�M�5>g�N6/��s�s�K�T^��[���4;�9S�m��m��V��;��؊3�9�UgV{���m���R�oR}DE��0�����*������Y�I��<E�����_wpQg!$��7��<;p� ���������K`�]�r@K�Ǒا��O1<z}�&�I`��̵�Sѭ�Pٓ뮴:�_����<��ӛ+�s2��G�}��_�Z|��[�c�Rs�Bǝ�XR����s�,$���~����K&����]�,f�WP0�$�qCk4X˷�{d�'t��%���] �:�1vVoV��$�6k�Ô�d8�_�^5U� 8��z���3v5T{*��ZO��m�ÂD�v]޺�:��=qG=(��U\M[*�3�l�tUu;�
:,mGn�Jj��+,��)[��7�GLW�Wy���7�^��9)����t*BH���n��Y�����!-�D�y\�>�}v*^�>/6�.���u�^!�&��Hff�ü �^r2d�IiT�e+�%�ݢ�jէFK:��o�y������>����BS�mJ�O�޽����g��f����
d��O��*��${����Y8'K��u�ڜ�%OM�y��[ݝ��[�{�`ocz��6�ÿ�ʌ�{"��SN�	��Kun�U���3�·����;͐��^���ǵR�c<���q�����\�z�Sz�ͦ7o�8���v�Ozfs���7�=9l�芊�d�����TlO�}���o�m��zf�6eT@�9�ҏ��&�����{�<S�v�L��{`�M�^�Oj1�갅&���Qvs��0�֙�l�	7��*�zyX��vt<���v�v�1�O;�LlZ˷�[���Hs8n�Nޙ�kgC+��e��������K=������}��g��;�9_hV0i0�EE5��f�ip(��]�����f9���®���(ě�о�Ş_Bl
�7���~�-C��Ùwon�Q���ܪ=#�u2��`l��u���|'���y��_l�L0��p�F,t�Fuwbڄ��K��B���'�M`�%�r��74nO��z=�Z�C{Mt�b?��x�e���4��kD�&�4��gdu<�G����D�����&�m(��^<�����t�:z��³߬�*tZKs�o�u0ԣy�wDJP#��k���'�ղ����ѐ����`u�:�ڄ(�7�%�ޛ����ܲp��̫��{9���Om�����f-ۿ�t�5I��F>��<G^ݺ|6f��h˙/�s�+y���Y:[s��E�<��9�������]�d��P���:	�3w�i576��,�f\8�BXc�셫p�{y7:^�-Q�������nf�_JUe���y[ ����Kj��W�� <�����M�q�ܵ��ǻ��k���w���޸	g���]Nw�~k%��:Lȁl;LW�;du��Ųy��BQ-N�VVo
v�����uc�L�dEUnT�S��H������f#^�y�6������
X������ƾ��!4w�AXu��J`{ْ�;X���on��~�m��S��n� W
8q�M�F�7��Ņ�y:�cM�`��N,��w#x5��'.�ۧ��Ǘ�@�KHM �\�{غ��M�����j��;�?:��-�*&������!)Jm�q��,��Y��S�^�c�O\ܱ'�*��y���3�H�x;���v��xfC�7���)��[3p��z�詝1"�l{W��<x��tnd�눞��]˦��kz��hխC�6A��z�Ǌ�v�yA5��#w���*l����%��YG2�b��ys��.���)Z���<U����-�FnL���2>s�ݸ��l�a�r�G$�0{	�Tb��|/�@�I8L�bU��;�����RFV���/���c��ESŢК�w�Ңr��<���&�{���u��uAIK�"Z��T
�d���)R5s�ΠA
-��ԣs��ߞ�x�=-��l�	�u��2�7���y���)�C�u�ϯ ���z9�uZ�z�3��}�}�ԃ��=�-�{|�r�"�J�Ig?FgH�xy�Y�8��1Ժݒ�� �)꺎�SS���^�*�>��O��w���d����瘃o�lė.ݔ�K�v��|�vx'��-�Y��Bi���99�6�UU�v8�j���Tم7�7(���]�����`V��L>�-���Og�!ݰ� ��ѩ�\�Ɏ9�COn��;f�5�fP�O/�2��4�|��@n'�]ٳ[� _�/R��3Œ�k����g0���^p5|���l��3�M�!¬��Z�#͜��[k��/g���@	�����.|�$��Atv�<�����e��#��
�P�R1+;�\�s0���^�Y��Y�}�9�!qba�l�ӊݸ�hO�M�؍ó��0{�.�]yHo7�t'CE=��4�G��e�:/X�yWZL�#�k�E�E����:��qf��omΰzAq]����<�Q�w�'o`�!C[�'M��́��d��5;���UG��nQ��Z]��4��y���;=����A���3���ם��~o�_+��>:��6�ݥ�s����o��f+I�g�� #ցv��>��h$�����1]k\��nOp��Օ K����`��'��;g��&��=a�D��vu:��rkcv��6o%���nMwf�;2�Y��7n!U�������ٝ\���׼���
�q>RU�����xv�=����f�8������[d���K=�L�q�R	��t<;�S����^w��4�=P;�1p���h�5��o{�5��Y�cV��k$�;�Ҕ�-�D�t���V&�5�Z��b4j�*��?��nju��^�Z�=7�w<�)�v��#���Ι�oO^3��,����j�O�����j bޤV�8.�폅�,�2�Gb*�����Gp+Uf�8ޠvc��r�!�=��L�+�w�������H7eU��8��u35�������Y��7��B���S9Ӊ�񵥁�#����gRA�g;.WE�Z�CP_ryw���.^���݂=U�v���Đ��ξT���*S�b�V>�إ��Z�ig��dՉ𱺯�8�
*œ}�z'��:2��7��X��m���&�厥�ōk!mW<��a�:���r��4�R����A=,9)�{�Ws�i���p1�֚�y�֣�]�;"ũqp��c��v���@�����.������	��b�j\��r��A,2���3|�I��U_t\^_��f�\vB�͌w�cuǺ�! ��1�1����;�y��w-
��&�EjZM��غ��K�.��s������S���~Fa���,7Xy]�|I<��3*.疱��]��Y\�Fg_":�nU�C�V)2�J���H1Cr����8S�L��C���l��ګU�(�/�,]Lzժ�ҧygw`���2��1��+���{��z��V���{�s;��z=�2oP�y���q��s�;�ܪ��:vN#�\í��rY�t�E��S	;ko��H�T���R�U`d��HDiǹ�E�c��|��A��wfr���-�$"��(�"�D�_[G5&F���P��=����@r�b�����>�9��S�����w���ki�����\XhMf�;3�1�qf>�i�nޜ��d�.�ᴖvؗC���[�	��ѻ�v��]�a/U5�*�7�\Y�s���d�Ҭ�4�W�����;7U��u�q�u��r�Օؑf��[�&�nt`Q�}Ǜ��ee���Ч�q�u;2��irQp�}Tg'b��������'��х{_S���u��s��F^s�հ*w���D����FZۘبx5:3�����$��'�����e]w2�R�k�^#�+��Q*������pUە��^i¼Q�92Zۨ��÷�4��qLk!��{�n.�ʘ��\�:I��I*�����
�V���Q�c�>ΈAu8-m
���҃����j^h���I��kn8���i��v���ъߋ�V_5��ͻ՗�ժLˎ���e��[䳶�wu�ނ���S�����'����nAa"<(��}�4��Q�|B�r�����8�WMK��Hm��9q�upN�mtwn�d�о=�L�޵�!�����w��zps���F���q'��� (q�Y�n;�B��a�Z���;BReF�dAݕp��֦��X�f�oN��p��ط���FHHU)�u�f��5qHp��A�RHQ�t���z&dS̏P�ݹL���._�G������������__^@`�y�4DUT�.2E�)�Ep+̫�uYT���nߏo��������>����.��G��QDTW�"(����#P�Z!D�������}}u��������w�7���D��e3�e���a#.T�G\�Q���ǧߏ���׷��׏��{{��w>_ZG.tZ�r�C��F�:.b�Gg��g��ߏ���׷��׏���i�&�I>�O2z�9Gs,�sև�+�Yw,����w�GS]\����==����}u����|���n�z,�}���s=rQ~z���Ew6�z��Dw$��䲎���<���^dRer����X��=H���Ȭ�\�Q�/�w��"Z��*#D����(��K�x�z�����me>�w'��V���o'.Q9���>U{�|�y�2��~�~|=K��[�l�˔ ��_x�:g��P����Z'�;w�ۮ�P�pk���[ٍ�v-�T
��p9Z�#���	�{���$���5<�����V��=���R�G�7��ݛj�Jg��cz�^GQ�u�_��yN����`�8*�79�Z���u���9FQ~���]��.zO 0���tT����+�ћa,��g%��gU��>����c����fɶ�Q�����M��Ll�gxww�C5��:��s��8/��h��8ўl��!�묥ՏX퉞�5�[�7ʄc
���Aphw�=��]=�7G�d��u��w 8Pw�o�*��Lj�Hz���_�3ɋ����O�)qB��zU���&"'�G(穩L�:�z��jֱ�1�8�3�!g���o�Wj����m݅T��FG=�\4�w���z�	��<���3ƭ�:��5�s�%�����I�z]�������⃦Ƃ���Z��@M�߅3�Nl}1��r�]����j����.��#���'�s��G���KM׵�UQ�V����ub>�A��z:Z&0���f�5�*<��:C��z�X��Y�N�m�����4��|����]g�9o![�J�h2��Əm�Q��s֨Z�6nRY".��z�*9BVxV'ly�R[C��ҭu���ݽ+=� U(��F��3Hmp,ѷ���o��� ۾��%wM�mu��ϋ�@��gk�_oa�+ݼ���;��wa>���s�(��%��a�������c{�^�Uo��r�[�_�u,QH=�l�`�X��`�˷�ᮠV�]ϴM��R|�>�C3�ݎ����i�v�sg�Zow�/c	�4R�n�ot,�Zo�l��lU���O/�����tn��ܾ�V��ݳ����^���K
v�iQ�����b�t�_g�p������=1ѝ���j���
}������w9+����������N�c�L��@�\f�Ψ*�����P~�R.1����
g�V/�B�e��q�������2�;�������yW�d���ډqW��5
�X��n��Â+i��Dp���n�I�S�q��ᔫ�y��rt�׵(��txQ��ȗb���݉8��[ܣL�S�s��c]Aj����:�8���؞9K
��B(V�wm�\gÝ#�����f���	y�,�V{t�Cf�0�A�$Q2���m�I?s��|��7��G}�e�Ğ{�PޜY��[U���ѧ@U����*���Y�C�\�
�<3l�,�^���_O��e�k��ή���e6�jTO�jR�Mp���}F�]W�ճ�{�1�-�^�^��7����^E���:�h���g���h�y�_6�"��k7�ȍ�+{��U�hT6j��W�_3������!���V����To\z��oNB�R��9\�'�Mh�	����H��73�ǋk�珙oI��D�)�V?R4�72�K�>��L�<��(�ɝ2�ok@�����@%˷R7^��K𙾉�xD˺q_�>�<Ώ�W}��J)�ޖ�S���oܞ�����v{�{�X~Q�U���J�|��1T�}H�}���̙D{mG��]S�H�^;����)I���{�v١��2�ܼ���*8f�L����j&hNgnۣ�����el6|8?n#���mR��`��;�xhϻ�y9�.]��w�Yv���������uԖ:���I�;Jv� ��s ֗J�ݳ��@��|#�41{I�^ۊ��E3�d����h��>�E]�u卢7N�����j�]nxnn���yi�h�6|�z����6�6V�a�Ȳ�ȡ�SZǏ���ޞ��k!<x����&�4C���T�\���h~����Ɯ��#�sB�9�ƥ�[���d_-D��Q�9W{�ћ�������T��x��F�Ѣ4��k�L�kDn�+Q����7o]��5���'�z���^v�}�7�h�
��wgDAS��9�|'�6e���N|��3q�"���M����'���򣲦��*�!��"[��͵�@f�ˇ��ouL�v~��U��
��?
���⏻�_���N�a�aLյvf.��9S�qR���n��|��ݬnW|��8ںޥ�3z�c��@0my7)�K�7��r��z������melEc��n�Do��j��3��t]�7㌫ĸ{���,��_tvZ�����bK�,ݽ(�I�l���w���	ʓ��7��Z!}؆�R�Ht�YT�=���:S�Kp��-veu��f󷹇z�ٝ�]��0�j�@q�?��~������C��c�rtό-��+�.��5z�/�ޜn&vq�/���R.sH�p�^wZxxS���gmt��g��]�+7��+��q�p��\1�:���]�;��]�ȝ���6���s-�I��9�ʵ}EA`�������w+�����3���i�g0K\+��Uk�����:�oaH���! S����_��φ1Y���Ǵ�ӏ��(����E0��ͮ�U�Y>�s�x�~7MHk���zG\���h��Iq�s�ib�^���U��l}����_t��8;��GCႢ��%�392�v�����Uϙ���v���s#<�j�i���3�ܜ�5{3-�up�Ρ��J�"���,����7�m����M�@���w��:��K�;e��5u�`�}W�7o�����:?�K?goîɦ�������*9���'Ƕ�=���q�.M)�6;7��M�v��z,�gR�ш��K&�4	����4�p.G~��]��ô\����� z�T�q�ݛ֗u�ʝ��{C <�����ٲ�@q6]�6����R	Wa<R��'ϻ̷�|�P�s�i�fz'A�{0�%��zC���n������c�
!�k T��"�Mj�E�s<�VN��Ms �����U���m\�x��)K�<��t3
�d.��n\]�kwzՠ��>˿V������#S�t��<���a�ES�F�20h��UJ���j�� �4�5��]�O�9 h#�L�����x3CK
p���wM?�O�;w`�
Ep͸���PhIn�7��}h���[+���u�K�q5��v��}�}1� baE#�e�8�������o��[�7)��m�m%cy����0�sSm�,�vCw#5$oD�nR�$彻~H����k`�����uQp��&�n3�f+ӥ_��kMR�����\��ў��F� �!�a�|0����B�kXv�;��0�v�'\�V�(F�h���/;C����t�җ���B���k��,|}�b1"����})�.�l��	�,<�-WR<՛���q��4MpMNi�t��u<�mY�^��ܓq�Yu�l���}n�3��;�|d�&	2I l��m�e��%R�(�C���G ��۷�Ov��������#���PD��K0l��A1�oFwo�V=���͸ٷ��o__[S�}D��1|�˽��1�?vH�0�}.)��W����o��z�fz�#c��̕�⢛�p��q-�V۶��6��p]�mF�b�)g��uAh²���ދ����7�=�������Y���{^��	����V2�5ڡ�C�kQ���,��?���v�3��C���G��l�
��i��G�g��܋�ޓ��Y9�1#�v���i�o�k%R��6�V�^�d_#���������Dǫ�������*����l���gS��i����@}�] J�u���ې���||���e�>�_���c��OD]���"5���g2���n���''\���><�Ĭ�%��5��>��:��Ou��z(���2n�)��o`�0���� v�o �;od����ɩ�ƜTҪ=:we'UMn��l.�.�&�dl�w١�ާ�G���V�gn�F0H��9VbF����3����y��͎� Qy��I=���î;n�tvtV�	�͆�M�2ܤy�AJ���"Y(ު�+־9Z�7��٤5β��;G�S
{|��c�/uu4�����L�]��N���j2m��Jª��H�Yvȳ�ioa��T׻N�<Û�|}Mp��/���o�����a>�󪮕S:����E��iv��b=����0}ޡ:��M��뾎���<tm�Xd�2�])չ�b���Cp?��E�M�j��J�΁��w���:`lF�}��.r
w�����pt��rl�n�U�ZQB����P-x�{��	缯���ב��X�'������E�B�0:G�Y����@ۨB2O&��3Li�We���_�hmx��d����>�����"Ԩ��.����r�Ȋ�j��7��k� e��V��h�p�M���s�H�T.o�n�"��&����)�'�ꬕ^}�θ8�έ��&�T����SuҲ2g�t�3f�T4�j��.��3���uye�l,��'������k]-J�g��{����#�A6C!�G��@���[�v�I
��^E�A�u>�sL/��VU��2"�NH^�_<�	o"3+M�3.>@�>@|G�a{����o��6��oO���ANY�z�
���w�\3l퉩��[���wi���[ԧM;Ǻ[��ە3��'s3�US��j�[�	%�z�L3.�,}oH��L&�*�>���4Dɲݠ��t\���~^��x��єUU��=�[�}�a\8�o_7]-��>G�����B�pf>�p�Y����t���wc�-[ui'7{wV߀�4��9�H54w�S7����e2S�����[IJU�S0���ǻE�BQ��vCW�	� |X�ؘ]��nG�-�
�i��wN�"�e�F���;����\asݧw��MdJ}�H�6	�VTZ���;t�t6)�Ǹ٦o����ouZ��!hN	7�O���U&4И�,��s�<_6�e |�'���8�7/r<�8W@��|���؜�����v>3��m6�¸O�R���ߝ��=�b�	%Κ�ǹT��å��&���eL��8�]�`B��]S4�c���E��z�+�Ipa~w�]�{�[C�F���\̊Hwm��7㜼f�μ��M��Ss~َȷa����v>�G��F��jf6i�W���+���j���8X`�&sM�oG�s�Qw��Ѐ	�fwr�k{���z0Q8V��H��PO���~�[1>|����`λ�Ò�X>�ʮy��e���ܠǆ���u�ch�tݤ(�W�G�Dߧ��=S-�a7:+6���ܦ�ہ_�����:3�}LEL����ƽ� N����e�eΗ�a��r ��}{����ܧ}��oO~�� {��$�X7�{�[d��M�ΏYB�Խ!+��+�R3�eS�xgz�Cqu-h�홚���������h��:�=u{���v�N�w����q�s�����׭�so:݉�6j\#Z**��o�	������͕����g��8�o}��T���Z�<�+*`�������A��|>��$|W7�O�.�n~͂W35���m�ńm���v���*�Ez��N5���4)��X�[�/p��Q���V*����.�Bٲx<�諸U���$�ڗ̴ֹ�B��%���_N��.�(�	�`Մ�;$𼺔Y^�sNj�o_p�t��B�&i�3ͩ�5E\n�Ծ��:��]��;yݧ ��w�v/���ϭ:X�ܔ�Ƀm;篁**<6�؄RM�R�?;��.��ff��m3�ܹ�w�5�D6j:T��m�u�V%�Ԭv]U5�X��2��8Av\5�㺇݀�:��6:���Ek��<����S�`�qbN�KJ�Y5q�_c}w����h�Թ���i=�:��U�m
�G[}��]�.�;&nn�\�4��z�J�5��e�o��[RG�nVc��pĄ����rv����Q4/C\J��:�u�qZ���t�9<�{.�.4�~f^&+jx��X'�Q�g�&�^𷛼�b�:'n�+w*��7E��j���\ݙ��ڍZ�T�H��7��]�����[�d���d&]`S�Gc������[�nX꽾4^�=,Y��z��w�;#.򤽕��↡�x��R��Y�/+�ً��0�m��1n��v�s�U�v���$j)4r2�[�$嚻�ɗ�蛽�{Se��
T����f������%5�ͥɩd �]}����K�k䕇u��2�[����ު�Q�;4�9�7x�\�u�	xIU�ӏ.%F�:��˗㬸m�Q9i��d±&�6*F�a���P��>zCc6HD��ZY3�ԁt�vCgF�Q���gq 1ph[�	�i��+�0��>��	
oI�Zv{/��O�Vݘ����IjZ<����ᴡ%̰F�ݪ��l{� ���9�*�u]3��⏻��rf�oh�2sƲƨ���X*�)�*�p;�����=Փv�U�*��V��+q&�Xj�h��d�Ϭ��}�w-���4vx��L힮ҥ�Vr�_"7q��1�u�����e������ض�i�n�ټ��9DW ��l<;���S���Q�cZ�U:�	�y��H�*=�[�zLD�g�O�/7w�.�]$��&�=����:�(卩�֚*n	KJ���k�{W�/��| 56��2�-���3��;^�̓fsb�9>���<�uJ�K��ۣ����,�hoo:o�q֤�d�jtԴb:A#*�r1�B�W��� V"/���2���h��J�Y��뎉���s�(����?�v�uX�j�=��Mn��ʙl'/�3U>�-`����䉢��d��_q��3�9�4-�OK�a݆�<��E>x��%,NB�3~U�9����ǰ5�����Ũ01�w�6�n���ĵ��N��^��ZMME�L��	D� |m+˪A")�q��6�k���n_q2�U:���B��$g$L�t+U^�\m�W�afqC�ve�*�L�m�2�HpF�;��9ŕ�=�J���}��0�DAB����0��m��p��(�B��#$w�9Ǜ�^lrHr�tԪ�����;ۧ׷��~���������׮�����\�ȼ�l�NN��w}��y��6�WR�,�	wt�]�%6^{�Q��oo���o��|ݾo����{�ԙL%JNQ}B�J��J"�jC���z���W����]�^�(��kv���7���o����|���oi��a�R9By�x��+z�z�#�U�N����)��c�9�^<{{{}~����>����>���Ύ=�����e���(�.A(vp���'��}zr�*���]]z�߯o�___^�___^�^Ý�E*��E䓢�-w\D�q)�'��y�݊��˗�p���G(��~g[�}�o��~����|�7������}}[��<K���7�{��'d����y�]u( ��<�e��+�\s�¾�/*:�{�Ay�ޱ�<�\�iP]����˧�/�+?W��r�K����nr��=���/�oG��ץ!�ܜ��G�$�����.�'*�q[��%�Hsa�Ei�x�89��NK	�$�H H<�.˶TMpș(�Fd�L��
���6#m�8�;�t䙡l^n+�v��H;�6:�����c)[�C������=�P�n�^���^�[�ѝ�a�S,�/$�wp%�{�:��U�{���S@�P�A$C���m�T�0Z�ed-�qP�s�� �.D�V��ΝYr�o�"Qm6վOWν|{�񈵰ړ�9�ӂ.C��NG=Vm,�i�l��u3��+;��w�8�����}�b��L�ݱ��wz�
��WoMY\wJ*��ަ�fF5��6��nu�8��{/�j�pҎg��Vt��yʊ�+c�O'�ui�:��^a�`���\�!����5*��F�ٯ06��b����;�7v��7������_�gN��>�fM��l�@Ctcbb��y�-��R	{vk����LP/��6� �Л+�z9��7B� Ng^�.@Ε�3���Q���Fk	|4]�� �i��lJ-������=ct��쥛NI )��W~���h�W���_�G��^�=6�K��O�zt)�y�TQ����{1'�ɉ�zU�17V�}�Wx���W7�x��0}�T��(	��?Vн����'��*��Y��H��ތvL�^Y|=�P[��L��ݮF�6s�n�G�E�A ��Y@�O�|�A�=^��s��A��V��]����ݫݲMT[8�\0#r����w�U�/�;�s�p�O4�0�^�3Y�Y�zp���{U��^WV��@��ct�7|�9^~�ۃz���m����3y���ǘĮ3[���o0�u�c*�-��U}�Ex����S��C�ާ�b�90:�6����{�\"�� ��r���-{S��t�B�-QP{�M��բ'�;�V�E�I�tC��H�ވ����s}������(2{˕�ڍ7[L�A�s3.ە��j���:_D�H�z��y�N�Π3�H���F��<�D1����/��ݭ� �D$��
�9�n7H�݂��(�v��N��I̼0�Z��{�/+z���p�}j��ya�g�M�F�uB9�h��馆֭u�/���c!jI�Ɯ��v}��a�#^��7
9��.�K��鞣��F�>f��&���ܟ6��0p?��}w���i7�Ӷj2X=�~���Y��~�\Uw8�k�>/'#��t�t���f�K�vmn��s��=f�iE�%_��<�S�Wܠe��#.�9
�|�d�4��j���u�";���]�"�kI1њ��<��P�Q�y����_L^�kͧ�LGv�.8���e��.Y���8Σ����Օ+�4���c*�zF�]���]��Pاkw�C-ަ��x���tM5�6K�]�S��g͕6_X�Y��	bmy�y����{N���x'jܟM&��j0�)�Muм���=�=��O�7�#�;X�u�jn��sf�;Q��"��}�!D��������k�R��Q阮R#�&rQ�~�sJ����i�ǳb�վX'�;���l���l�}��>��"�c��E ����j��ޮ��g>�)9D���wv��O�g��My�#�j��*�v���u�
��W��g@�P-ʺ�ʴ��GzUtP���X�:y��UG�X��7�~���v	K�G[�����9Hr�[$� �W8jv+py���ޑ��|����劏C-�rK��hKQ�t�H�,��������`�j�R��.ze��S~�.}��M���g'=��B��oY��	M�͓��Ô��:��TV�q��5�m�6}7�c�4�N�ۥN� ���4
�z���0t�:��*�I�y]2�Sw@?W���M	���z�����_mh�u�z�ϣMJu=�\��P��ꆚ�ZV<f�;���nu�R���p��ש���{�{l�uD�
�Z��cz_�k�p���T����X"�'V���Yi=�9#Ff	m�7���բ�T�k�Ģ��U��9����@6���;���7��6��\�
�GmR�5�7q�g)'Ռ#͵�a��/���T�}������U<�k��+7wL	L�t[�v����}P��б�j��ލ��EG)���rt�?N� �������s�~����6�n�f�{�9���������Lr�75H�_>��I>}����g'�������>���Ʃ����$�"��*B�|գ���E��KQX�A��Mhqya��X>�*g�5қԺ6�#� �酈��+�oݦ�/ABp������>�Ј+#�3����3Sя�}n�-��$�|7�j"Zujq���\��M�n��uF�I>=���4��)T�Y ��_<���M����ۘh����uv�t��z�7+o+-���;Y����z��dbHU�K�O�����w���ȩ-��e����O�G��F_��c��uѲR} �~���[ē�n����+K��Pi�T��Jٻ��[�.�ͫ��s���&�8-+�H�����N�g$^�[t{���VF�ORvۯnkDf0��{�*%���X/�s�f	�;k�]46C��3rzɷw�1������z����mV�7�V�DH1���\��;���q$�Һ��s�Z�n�G�3FS��L�	�B�R��M���z[��n�K��	vO���?�#��g�h�(U�^��:�b^~W#����X-���Hi�)<zP��L�C�F��>�7��ˡ����X��r�׫鑉w���m�T/&8��Q��'�+X.���U��	6�ldx����{	}�#r�,��W�0oO��'!��=�_H����;g���,�I���~�8�^�[�l�X��gN�rI�k�'[7f�,v�wV�`���ݼ8��p.�¹����2�4B�������y��2��/�X�y ���a�En|�|�Q<(������6�r�͆i�ogG/^��<���S:�_��*�u��1q�[r�2�W���h���8���u}�8�p��K$�˽����"״�Vag�w����F��$���e�^נ�^z��SUF܀ۜ�t=q����N�OT�(�����[C|ˋ�0o3j�R#���N�qm�R���D�H?.�S"��Aݍ#��A�ʏOg�﹕3O�@�N��猟�vӜ��!�wD�0�Ї���J+=��Įg�zk3\v4T���s�Ƕb�����;�������E߹7�\�n?�~����	B���?J��$1�,X�oD:�V.�3GL�wES�[-�S��f��.�7F��ʳu����A�� j��*�'�����9��+CXoK��`6sh]n��I�B}UՃv��!��+�譑��zeT*��ԣ�v��cn�f�vkx�n�F�32)8U�����ޡ��n�n4?u�.l_<Ȭ944>A��}�\M��������>�J۽bq���y�#��Pf�ٮ�l9So�V3�3�gB���x2��l�{"4�U��{˔|9����}F�!�&�ۻ ��U89�wES�n��EN����7`��<�	�=�l۷F���u�\�[�]�^�`ޤ�n�םqͬ���6�9����0�݀3
�:v}" �1=��*��ѽ���Q͙Ǜ�j�
�n�>1�]x�Xр[�8�F��h1F`⛂ͯQ�v��Q�/x67o+e]��\�%�u��88�;=��pi�<�Z9�ff�m�:�f�ݴkp�36=m3�Ćy����Wz�Xa��|L�23���^wدE�69:�`l:�;�¡J^yܑt
�K�����q��I������X��k1_w�Z����q�D=���>���]ԍ��Օ]=�Պ���3]m�{#��o��k���4�Q誻�{I�Qk!���y{�7&��������i��<��k�}�bC�2#� ���;����q�rrq�/-����ݘ�p��N�����"��g��ou��*����ܡ9���s}��4bΡ��Dw��c˒�Oj�S��oǆ^���<�L֦���a�~¦����0[��<l�s˵X�^v�U��El̊��Cjɇt�^�������	�O�n�y}��`����.j�V���O�%.���	�	�!+^��o[at���|�6�!��K�'���q��(�:��cn[���
z���*�����0$�n�P�nM��7��(���I	Ck,M =�l�P�v�0�pWl�wJ����&Z�a"�`U��tO/]Hk�D�Kh���2�攑ռ���K(v�m�N�٥���$��5�ؖ�?������9oJ��)~q��ML�\���>��#]gJ,���5x�݆�Ưf��(��ʚ�	SS��v��[·a��"�qݵi=��_�o�9�����y�
�$����?I�y�b(�OK�@H�W;���4h�udo���Πїw="%�o
�������K��͹O�pok�5�b5�V-�����
�������p���<�½�La��b`���fE����@k����=X�[�W�D�?S:��ɷ)���9}g��
����@�NZ���7�q�A.�٫]f��U�w�r3k�+) HD"�H a��?�*4��M��"B�������1��+X� �a���]�Eռn���[�{Z���1�����۸
�滄i4�m&�%Ri���x.¸�4*�$���/W�
D
7Xץ�i]��b�`J�Pd(��J�V6A>���?0^�_@����q�f��},^��򺙤��v��L{R���R��=��fz��6>�]���'��8��pCZ� �d,����������I�]wi�3���>���j�����d�oz�Cy*���M<��=��'e��KZow;��<��eF�'[�|�m�3]J���9�E����
���;ʮ�J��+�{�7j�iݧt�j��<�Ԡ��6m�t�(��Wh�mT������:s
�I��koko�������,;��������7�5��z_@�iSw���i�ўj�I�!y]�=��{%E�D��d,�hA��A'A�L�Tx�;��r��I�L��n]=����� 7����=q�x:J�ҽ΢�7,�ѾX񮊯ts�}%1ܿ}s���w_]E'ݪM�}���t��9,�B����pb�l��Wq���=ۯ�a����םG��z�L�e�y/v's}z��%ા�E>-��t�U}+z�������r姝��}�n#rΈ{wB����������:`m�zvn�	�s=~��4�^¸ËB/c����Gwd�*��i��������X{�צg]u��2�Es(J�r�7^c���-��u�����}GnTy�c3���L����̫�E���}~���_� a��ԈĽ>����� QK>o�{��9B�ɢ�O�{���Kic���,�@gA�V�<'�}ˬe����8%\�/��4�ozۡ��_̟?�����sh����	;1�㧒Mi$(���WK1!�h�[k��:ܫ���[����ޗ�L�[8�)~滆%W�����Wk��߼�y)~/� I�>�=�3�~X~ؖ�_�ސ��$��p�k\Wf�p#W�R��l5���c�T��MM%���|)�qרjvX��쩬��̻��"(+��;F?�=����N�^�w��fm)����,�}<� N�j��e�>�_-��]�"���gPC���/�t�%G]f���ɩ�\8��sW��ؖ㡋��wh�;&u�-w-ޓu����h���uWN㗺M�U
��,�<�����b��q	��w�t�=V.�t��J����/����`
�+mbU����w�p�ܾ�{��S�Jǃ43�H���ec� ��f蓷{̣���f	�Ϙ��5w\7�����íx9�í��AKz�b��j�M�|�(b��:�2�S��(]3N�.7��7�ev�B�K����m���P�m�edȅe���:��sfDŌJ;)�ӽ8^a����R���J��Q�N��:ɻ����ˠw�*���
�\]+0���N�6���ﲋy�@N�M*���t��GE��--��� G������W,�k)�k9f˽�4Q�Y�"*W��RƮP��Ek�HU}��wTwU�ݕf0I�F�,ڤ��u�2V�k��U���SE�f6�V<�8��{O�9N�a��m���l�F�|u��=�j�F$�E��n��;��q\R��Լ$�ף%)�ېwJ��Ӿ�;��m�s�>��D���#,溩ݫp������q�Q��%���6onK��h1�k!U���/�2�<Q��&�r�5�BIG�gq؅�;!n;=���(�;��C�U�7�:����*��-�����ֱZ�菖8^�K�|��e��bv P����2&�v�"��{���X��۔;_���a���Rb�[��Aڊ��2�$�k�)ӣ�][���Gkr���s��N}[�t�	���:��x�O[jnf�
m:XЈ�-��N7٘��V� �}�w&�G;-���]ٚ����;�@��ХˣY(TR��9�Eyn�}�{�oj�����.�����=��>;{`z������a� H걚�*�}�!J�Z{�*�*�h���P�@�ok,,�J1w��/��'y�4�j��j�?)�������+6aXpwm-��i`=Jum�n��F���q`��Ն�j��[�k�"�W]56��G��m][�!dSY��k�y�Û�՛ޭ��E����!0`^V�V�݅Y���7$���zQn�<�����'�:�{�'mm�=l�%�Z/9�U����*��n@��Gn^\o\�lX۽ћ�r �1��ә��ˇ�Q�ܫ�C���a�t��,��[�'��TRT��E�U�N��t��8K�CwF����A>#��Ǐ��s�w:�RI�QN��;����x�jF�Fݚꫤ�Vᔯo����{{|ߛ���n�7��|ݮ�ӵ��s���u\�]ܼXRwV�xd�^k�y^����y����v�����w���n�7��|ݣ�x��n��=@���u��qù�x�5E,�S���W3���������뮺��������p��A�s�Õ���齏w���f�#���e�qurP��wwi�Eî\9�����������_^�___��N��n:.x�:��*ga���=n�Y_�^=�G'���������������������C���	�����V�������͝Ⱥ�Q��n�=�ϯOn>=�]u��������8q�dx{����S�<�떑�N��Hr��0�q�)�ղ�"&BN뫒N���f������}ý��wp'\��wR�Ds�/Lw7P��"�]Ĝ˸WWwd${��ݻ�ם��(�u#�G�+���.���+�x�������^d�eN �d�8m
��dO$�G��~lK�a�k*�v�ƚ����ۨS�.Z��$j��'7 �{�V8֮�:��v���n��4�=�'��vǖZ_�[s7���&񀌚���
�[4�:���O����-Ӳ�Ӄ;u�����/�c�t�mt�7k��O��1�i��+��ӏ����6�6�I4�pɴz���s�ni��VotA��TN1��}��S�ջ���5<_@~��sg+��%����w��0�4��+���NnY�.��J f��~_|�̇�ye��j7��}=k.�{aR`ݙ�v(l�(���;11�4�(ս�a�;g�|�e��w;�<)l�;QoD�ʉ��n���K���&7kG�i�O���W��A��K�:v J{�j��w�����\�>�<�u��r+���q��O�����ŵ���V�Wztܗ^n9��3:1dy��y���5ݸtl��rޑӣ�K\�|���~:֚Ҹ	@���rld�y��ټ!wl�{��3��>R�W96�*�n����O#�\���ۜ^�7���]��YO�M��1��i�M��ښ�T>H���Uq V�0�2�t��
�]]�ξ:�O�q��`�����wYw��I'��J�;�	���TB]�w��� �h]������_�v����$��ʅL�V��D��1�_��r;;�$f�P[��{Cd����S��T/r��ݖ�X�q��8zn��`���:[	.EϹ_�6������a��[�����A��yn�` ��Z�veII���vP�w�<�����+J��u<��+�~Oi�.�n+k�n��
z�]����J�z�G��m2���Cˮ��|�c�̖fwpˮ��������
��r�VJ*���c��.�/;=Zˍ�Tm�H����r�D�cI��ffF���J���m��y:vO��E}~o�������t8z�>m�	�hGO�QRڸ�>�{M�7��ͯ���:OurUP���0�&�ێ��t�4L��V�Lq��pYwm�z�M$�o&9�ht�kݬ�qo�:i3P��2���tLy_*v�����*}/v�GΧ�
H6gØ���W\n�U$���	��Za��	1G�
�
�T0�Y�i1M
<d3��ʺg�s�Q��$d������^������%�ۂoq�����o��о����W>��#{5�A6��>���憿 �R)�
A2��1ĕ8�|d��Õ�@㪪	�|`�+�n���Jĉ���Q�>�����`�{��Cg&���+ue�V��p��o�����;�B�D�%ݦ�S)LB��>��M�>k�m�~�1}��@S}�w��{<�2�Õ�К�m�
��Z=�c=�n�ϫ��� �����B���c��� G��Q��A��X���43b�l���i�������]Q՗�����������c?��<~�7�Jk�Si��7���3��[�����v/A�q�`�����b��_3X�)�QQGۮ*����ϊ� �A��ۈ�f��f�<fT*��X(K�^�&L�/;n����d7��g��Th	�d���D4����Ě��R5=}��Ą�)l�ԙLC�g�˥��5ꇚ�ޫJ2��}�w����#,WX~W=�Lu/J�xк�jM �7�}}�7��E=�s�ᗵC�&ԑ�tv���/���By+���J��<maYՂ����#V��rv�h�>�[wMA���<��Vu�������}�1�kB��3%�����D��m�MgA�{2��D���7�����p9�U=��[��r��좭⭉�H���jVN����J(�ː
쨃������5T�vx��Y}��2$��U�M����}�w8��w�#�'\Fa�ĺzR��%�
7�y�ug�`o*{��}��j|�(�9:_������9Šr��s����#�����g��Y]���V�!�k*u�؝�l��-�\gթI;�_�w��@v{��t�ko�T�C���og���zΜJ��Ssv�f��@��%闝�NuA"^���C:�G�����8���G�Dy�2#Q�M8�q�~y�B��M����ѳ=��Wfy�vWF�_�dv�}[�
�\U�)�V����ݎ6&�p�l��w�i���>rc�� ����`M}0wc�����횽��m�z�v���jG���_v��E�����.�{�V8�[9>~�V��I�v)������Su�������+/��d�u�:n���n�#ݩ��T�׽�J�lԳb���f @P�VR�3x�<�RNwp�y��վY*��m�Dq��C��5�/9)�<x6�uނ��C��MlqhUÆ·��^��5M��������~2��'Kb=|�to3����-陙�Tp�":�@0%3cNuٟPDu��y5���]�B����
&�S��؉t��w�b�T�:��^�Y:a�%���]+�9Uf�ק�9�ق��s�~���w�����xڣ��BKݮ��z�B�3��R�]����٬�n��C�A�1�F(�"9Xhǯ�.��f��[�Uqْ��k�11y=��.oV�ߐ#�����r��z��.��(�k�F�!���\�cg_d�i�6k��8]x���kTy���^�_V�r#u�K�P�v}�9�8/.��d�m��k� =x�҃�Y]��:\�I�\:��aw�'w��n(�'ï�����
m�H�Ɖ�
.%e@05�V���K��/�@��A+��s&�f�`�s��sa��58m�C�R[]�
��u�Qk��I/1T׋9Sɥ\�q`�]*��]	6e�p�*�B]�;�og�2��������mϾ�0�y��B�[��'7Ŧ���+�����9>ổ�/�QZ(�����\ژ��dY6�׻=*^6���Ȯ�1��dɆ`Ɔ�d��C�{ΐ��G��D}����!�]�_�ض�85t�Y�[e��Qcw
�=�vB�h֜�!��aޅ�N-�n�e��_����@?�/pS|྿M��0HuP�3�7�����痟�9f�׀1O��Nr��L��m�F����7}�۴�����<ٮ(f��`������!�x�����I���"����:��8����:F�v��7�n?��aV��GR�m���o_#�����AT�oCN���W��S�Fw���U3����m��:���x���4�x�]���7^=�Kv�?�5��{h���&��nv�7�5&ޏ�����i+gW���[�<�u�HԾ��W�јϸ2m�����N��h�"��<̕B�~j/H��9^�~�[Ĳ�^ѷO޼��U�T\I2>Q�o�yERJ�dE�3��1��6�o�hHr5|3�)t9��l�+#�0Em�7�[/t�K:Z�KO]�9_�������9Q�]}��:b�)4a�u.US�N�&	0,~��9���XL[M��L��UU�=�ހ�g��\<M��R@al�1�0H���츿U�*�ob��g�_�#ُ�$��ڌ�h�n��)�9S'۩H7y$��w���F;�
��%09[,�`.���h�����%��n?�4�0`Җ�qT&��K��m�T���Ύ�Q2F���a��@I�`�ԩ��{<5� �z�ew�����nY���[fV�o�H{�v�>�Y��mMЬ�w̺�k:{�����&#��צ/��ʴ�]mm�vK�6n���Vy8�]��0o%w~���Z�UⳲ����O�;g9~��h�������~��� F��@Vd[��E���/
��ن;0���Z����5�3���p�=ٲ���@��=�z�d��冽U]A��v�2,8G��R����:�D���v!�9�~�R���4~��cXt��d��o5f܇��{� �'y��/*�:��J{�xU�v\��Z@���������]���kH;��e4��}�f�/�(�fV����d�иwA�[���vB�Y\z�71�T�c�(�f-���L��|8O �ā/���+ϹF������ގ�W��OS��S���h>��[��u�lP�!���q�&=2r�zHg�;�*�8�y��3�/�����_;��楗�MC>����:o�n�)�a��\���F��4��u�v�za>e{n�UP��������(���Փ�F`���z�/�Ց��I'vf�k�Z-�O{=�a_āT�r��]�=�>��s�Uy������&#ĚP����s�U��w���Ow��7d��Z�[h�;�30b
�`}*�9wl�\��F�����u�ƃ��p�={&�G=K����1ao_&�Q���b�= ���>����z�j�^�nX�톫�Tf�7��O�zb�j� �%Ww<h,��]:z�Ku�_	#X�wftf�68��A�z�J��ތK�tұQ�ט�|��̧HYL��g1,�|6�\������Ol���b��G���۟��i��[����ϹD�dW��1C��4���H �"�<���rLNvq�{ߜ�{�˄�C���n\z�b�U{�IRI�[��ZV�L��.�0���Q�䷲�]he�o �<������^�CyT�i"3�;��85�~zQ��M�|{����7^n���]�k��wOO_�d0�lQr##]����F���K^�	���R�=���[y� F�w�P���o����a��%uHC�ɉ�3[����Z��>��Փ�Ǥ�^���͟p�~Ѭ��_�����~,�J���[��"E���v����:��u�o/EV��B�=��.��O*��e*�����Dj�a�I��d�O������~/4����M��s��;E�8��F���V:���?S`F4=I�C�T�����L��c�&&�(-������w�m6�����9��fMZmeƺ���+@s�z�o�I�J�aX�ݘ�lv��)��5�Vº^�#485���\��Y˪ϩ+��j�{�]-OXܩ��<k�U�� �V.Q�,�[��ĆB�긮�f��	P���/_;�4����&�ՑR{����V������:���}h��v˒��\�mY�5����YQ�#OM7��BЇ�y����~o@'����=gS�u����xfx�[�VǶ��YxJ�����iO����T:���!ch�g����]r�	�n�r�i�k��p׮g|�jn����o�5"I�~W�I[Y;U��jcy�+�0j3�AW+y��7��6[sq\Ğ�#z4�6�Z��̲�D=��"~��Z0[�ߎ�1��P��t�-�ɷ���Ӽ4�������_�YG{�I�;7�bnm֞�`����\��n;VP��e ��3�83Biy�ʹT]d��87Hl�t�x�W���3��O�ưi�[�v���z:��N��woѸG@g���W�*�0Y�~�7�J�����K+@�=��k�?|�5cG��π�p�ὁbڛ�ߪ^��"�<�� �x�9pm�u7U:'s
���u���\�07|û����?�����s�З�@Q^�* ����y�T�����?��ttB�����2p�!��Q�V�����XB BTa	� C�7 ���@���J�2!*@��!�H�!
�@��"�@*u����@��	�ܢ!�BT�	@$@H� BD�R$QN�� T�	UR!�E B T�  TH�T BQ�	B	%D�P BT@� B%D�P B@� D$D�A@�!�@���
B��)��BDy�@!҃��###���� �X�X�  �  BUaY !	E� V���z@B B BEa	�% �$ �  �  �$W�Tx�� B�C@Ȭ! !!(!!
!*������8e�ࠪ- �����}z���~|����������|�?�~��������~��G�������/�
"
����_�ڊ���o�TDb�O������?�?���O����?�D��a����/gM�����'��o�����������\�A�PB�"iV`D��hE��� �
�`X%$X�iF$&P)F ZE��E��FI�ZU�``%�hFH�ba�fd$ZE�TH	V Y�X�a�bU�U�E�`Z�Q� �Y	V Z��iV X�
U��Q�`XIV`	FBAd�Y$V	FBQ`�X�fQ��Y$�a�T`dX�f�� V�b��d�X�e�` !X�d`e�eeYH�@�A�b�aP�b��%YXdX�deY�`	BQ�U�`ZU�E�Y�aIFQ�V� �fU��X�YQ�	!X�bE�V�b�$Y�dYV@�b��`X"Q�`ZE�%�h ��dYV�R��X��H�XY�Xii �Z�D���ZA� 	
A�$��FH$D��H�**��*"#J�:���p��?��'�*�4 � �4 P
7�:?�����������t�>>~�Q^���?������	�ݧ�Ï���c��Н���*"
���'����S䢈*��DAW��?��� *����z��Q\���Bp?˴<���p8����'װ���QU�d?��g�TD�|J?�7������������p?O�H�> Q\�!��ڨ�*��~��v��~$��@����?���@�>�	>~�_"	>|?�q��`~��t�|__��W�EA�����>v�������g^?�����?�1AY&SY����_�rY��=�ݐ?���a�����}U%J�$�H��!P�E!�"�)R(��R��P
H�T$�"�J��)T�J�%RfUJ��DQTT�$$��
�TH�)�RH$�DJ��
�H���)U)G;B�$)P�HUUI"@�JI�**�T�HJ"��R$R�T"�H�R�U@D��� A^   ک� +T��UB�-QUTV��*�m���(5U+b�ClU%��VkX��ER�e��Z�T��3Z�Q�4d�	)��)QQU� �(�@(P��va��z�(�-� [hRPh5Qm52�%�41�Ф(��-���҅)DZj�A**��  �]�F�J�imI���@�*�4��SM�"�F��Fb� �ZUJ�4��P��AT� ��Akh�kY�QX��d+F�BPh� �mM �UUF��c���ET��EB��  �
�+�i��5B�mU�`*�L�@h�J�#kAU2�P&��Q&��R%BQH"��  -sT��Kd��P5ReSlThiQ��,@����[ Pf (�X aUPI)*���� n��je0�a@lX  F� 5L6 
�,E
b� 4Y,  ��B��
�H.  �( 5`�!� �lP�Y� # `�� Xc@��0  �j�B���H���  Y��UQ1� ��� �� 3&� SL�[ j� ��
���@ ���i*�� P(��  8 ��  6lC@�#2� U�` �KTlh�1�@B�� ������TJ��B��~�d�T�0      S�	)IR�#C4���E"d&�S�2=A�A����!�JU(       �A&�������6�dh  �	2��U h@�   ::����Q�3V}x��;39�qg~ʘ�bg���w���_����M��{}�����]*R_��!Q3�!E��3S�B(��1bY|���Ǽ�$~���D �@A�P�
���#4�,HF K Q@A�Ϊ��c��6j�P@A�C>%6�MJˆ��/;�,�A5��]��M�*��.����8,Z�nU��i����21�[�^7ĤK,Q�)�+r�2���Y�Q���jTR_�53t��>��W!�n�Uټ�@��ss�c�%��(�g��Yg�z��8.�,�W��a�F��q��ļ��i��kͲ���[�W�f,�_l����B�֔�B��O�6��a8�u{�ID��I�@�*�I��k�qa3"��B���X�����VX�� �7*���F��+���O+1��X&+Kk)���I�0'*]��P�	b{n�$^�i��c�nDn�g`�DS^^Z�#ҹ� W�V3G6�5�ٖ��,�E�h�h�u��9Y�H1bb�
�l-�Iu3��6�d
*,֝�eө�`�6n����9�NU�+Na &B��Ѫ���=�z�[�,m%W�=޸t�p�1�t�ŗ$��ۭ5x�=P�JՑb�m���T�,�%f���t�ʷmT��x�9i�CP�ȨXѯ	�9`k���,:��F=ۛJ@���F%Xeǲ�Vi�zܻ�.����/n��օ�j0�[��F�A ���6��2��2�޲uJ��f�M�@�ٱ�r(f7�E݂n0I�r�l�U�z(�~g2Ԏ���Dʃ6�͖"U�������M]��r�ǎ��f��[�xV�����&˻��0��Q�O�r��0[�C
���6^,s��R��_Zj�*6�� ����"<b����e��V`5:1	�P�����ǰ�sbl� �-9�p&kƂ1���#�"�+k)�f�I:�l�Ô�n��^v�p[f��J�b�	k�Ӱu:"3V�j�Pէ�F]ó1�%�A�uq:I�x��hc�M�b�6�zMZ�Uk3$TMnԎ�xvЛ��%y7lc�y�H32���l������R(Y��xCɡJk���f�T5�Q`�GNJM[em���v�3�n��TU*F�^�יZ
,N� b�j�2�9QV��*�P�01zwLi` �xeأZ�'n�C�N8fƙ�Mk�x�Tr^F�Y�mԓ6� �n[xZ�~M6)��a�B�z��m�5ʹ�X�TjlM�L�Ɯ���geakk-�1�'T�-<2�dC�F�Jw
�u8<�
�S�֚����ZB%P*A4�Ȭ�Q�n��aU�h(����Z��ve���՜̨�p��G#�Xp�j�a�jք�%j泱PC(h1��.��l� �!Zõ+Ek7#k&����ʀ�,L��iAB���jhК*�:���K��ݙ5���E�o���C	�H|r[�y�$�Z{�iШ	��d2`�
tĴ� ��ǌSX\���t6����[jnfn���R
��+̵�ӛ-�v��u<0U��%�^�EP��p��|��I䩤�[�����Ff*����ؽ�H������wL����b���$�2N��\��F8�9�-퐱���]{�4��'+"���t+��eaw���tLZ�Y��H�Dc�@q)���!O�MhO��vA`d��y`k�u�썑i���WGhe�f���X��V1���J<�*6��ǀ#y��[n�6ȼQ�u���D�n���Ĳ�UͲn�*fY$dԫriGC���$h�&c�X4J�Af����=	�76-`94:͸�*�1�L�8 Tk)�0��a�T7,����Ҵ��	IƤ�e�J0Q�"���� ����{�EsOp�	�˶՘@�Z��
*V�&Q��T��J�2T��d_=8F�Q�{M�rC0�0� [[�71���̈�+'�ݛ�r](�`�Y�F�n�e7����Ȧl���t�\�������Ԫ[�lཽ�n����!
f����ŧ��lC����,�c���k!�c%3Q���'�r�lbq�N��Ӽ��K��[��ҥ)��G2�y���i�gnE&�x+i�3U���22ٷwL�K����\�%�p,��������˼���I`��7�V�+iA"���߬�Ak��ne#0�&��D^��Un��dV*L�C�X#3M�*Zk�Z�P�3r�hT2� �#��i�z�P��O#���Ow�{�ӆ$�)��t~`����IS���]��V�`�mn�if�	�H�z7E,I'z�Od�r��W�&M9�{�r�����T�"`	2sV� ��5Fe��&|��%���k-���nT�:jC �Lȉ�إ��+��W`<W�p&hawxL�R�cF�lُPp�ˑ�̃��K�[P\5�eY�LU�.�������ұ�]E���qJ&R��ye��;�z�!Vk�uݺ%����g�7mT��sH�sBӃ����2���8Yw@J�R���Ymn	g�0��!ٳ(��r��&�P����J7Il� B�7UG(.+���S6+i�9 �X+ȕ�Qo&ErU�HIAQ�%���"�v��Y�PIi�:��ƶ��ۛX��䁴����'Z6��$�)��R�[4w�mcz԰�kYx���;� �	��Q���@GO2f�͍�R�s6��T�R�����Q���Т
�9�%�$��)hB��\�m��+(M8P�)���50h᫰J����3
���*�7�MT�CcL$��ϐ��B��D��f\Deӫg���fS�e�9�jV�
;7Z��a|�j��w�c�޷�*��q� c���7��	����p�q�sb�l��R�`�z�A*4�9g��ܧ!�1C:�A���v3���{A"\��ۭK	�/@pػmXb���ja8c�XHZV6i��3v9,�ly[Ӝ��jo=�M��L��f�y)iXז�P��Q^䊈Vh�b � |V��6��!�/^d{��49��fbx����kL���o2Hv �I��M@F����Ic�d�*���dn\��D��a �b�`� v��vu����+��ۄfb�V`�ʛ�F��8ȴUX-ӀTҎ�P��l2)e�ol&�:*��i�YH�+�9���L�J���&м���LZ�C %y�G �dՠ|�nQy����+�x��4l
��ֆ��&v��nJ+,!BR�a4�'��*�N�bvf�!��ؔ�Y���{��T
htm{�@��x�7t�l�I0��I:�B`��X$�WD�:�dT-�u#A���a�^�vͺ�@�SѶL+4o]���r��U6���&�F��vafb�(�;�Q�=���L���������݋(U�hSn�2�R��s��Nœa�b]���J�I1���Y�: ��;���J��Ӕ������V�L��JaQIc,�W��`���=˥���Tu�����7�*T��a�"��p���Q7*;�et�52|kbT�]��K[�vo2�Gb�&m��W�+Ia�OE���6%���U�ؽ�*�^S�U����ފ8�v�VU�ZGM-��v���jVm�u!`���dT^�5�x��k[J��nq���E��e6���cj�-�	Yv	�P�Wf�&���4�"������X�l1�֕ �19)�0�L��f̻ܺ�B�* a,��5TEZ�`7��v��5'Ұ�-3Y: /s��R������ �ݒ�^�[Y���Kn� 9�r�xh�f�6�QHR:q�`�Y��j:(�qQEt��;�Z���{��(�:�T�q����]IQ��±nn\Z�[4! !̱;���l��-��en�F$���%��z�$r����4��-�ց͊�Ѕ� <47L�cf�:�8�j3�J��L��^��`�*XPS(�hf�+���P�w�fdn|�(>�I���x�u�X*��r��^Znਃ`k�n��$Ч2��a��:/1+�@��Cf%@�5��-kZ�Y�얦��Y�3e=�5fh�3��6#�KF�����ee�V�4)1��w��`��#��ga��֝��d`j��<�+��1�<[\�jȡ�f������b��N���C\���*�U2<%�W�a[-l:�)W��s.	ݻ`=�:En\�YI���~b�u��bWW��-��kU�^HV�j���&��$�Z�wn�˴p�ƩL&��t����5�{�
�xE��Az�c��"!�Y�Ή��;3hY���5�i���Wy��E,��^�0�B!ڸv�ǌ�sA��Xu�+�t����42�0I�='�m�R�Fk�)� 2��h��6��e�p��嚴���;N�7R�|f(U.�f�M����^\�H�e��J"µ2
!s U� �2��k8QFښCŸ�ԭѧ*�+�;�/w�SVYy�F٬��R���г����TmnU��l����m5u�P��z/[�6Z��ZӉ�{&n�Xu���w�l�t*R��3��*�g[on�rY�e�K��R�˥� hl�Y�ۆ� �i�&]M�)W-A��0���O���V�d٭� ��򋔚͒�U�f�
F6���O*��툐�B��9W�UX��Rc)���,�F��n1������'Ut�:q�@I��T��n2	&�Zb�]�REV�Hj�S1Q��2��I��͹)�(�(1Yq�ݢ,�Pk���4�BS�0��Z�K����M��j�v��i���à�d��ݫ`���F<���]�ֵ�k��95P
��nVp���҉RkZ�@�J-k���5 ǩ�vťo9�f�-f�Ly��$2�=)�Y�+d���3t�B%��/tU�*7�*u�m�
�(>�q1�q^��J��T���-Hrd"^Q�N��D�d��5�sKf�i<i$���q���7�f\݌=�m��SfnS0�Nиr~;Y���&n�de��U��"�Ssj�S1�d�ޛM�0��u67�E��o_f+h����fՀ �Z�ƛ����F�)�BlǦ�L�Z�)IQǆ�J�
tˏ �F�����}"f�6η�e*xE6�챴�̠�$�7if�nT�{j-g���Q�l*�ӎ�?����KY�3U�g3�٤mPth�B��jN�<�[.�e���7QP�:�0oq��N�KtQ$m<_H\)l �3*�D��k_Re�Ti�ִbwR�Q� +!ƣ@�ӷ)ǸQ�@[#u۰�N��,�:�L��wĥ*LV����Fӗ[��j�I)�c �i�u$݋2=XH7.���[2�v�=����ԡ��̫5��cX��"�1�i��j�V�Qxl�O����#M�r�e�`e�p\��ȱn�$��e��+#ᴅ��}����T�7h�$����l��-�b𘑿��{��zs�d�pm�ʵ����ff�Z�:D=�Ku� Vqk��2�B�Cr3�����+R$�{S=����	y�dCebn
�I�a����Z����0[���j۠��F)/~�p�ti���@w5j2Y����Em`��57J��sY�x��hͧX��A8m�U�Ƌ��Ѳ&d�JAti*V���X��ۨ$�Q5f	6M���2�C��D�l)1�k;o]��<�:�(�k5�b�ʫ�T�kT��\�wn�.�˴�R��B-�V�t�sw���3Y�Qk�3,��_5�ժq�n�ï{��=#2ˌL�{ze�'Q䌱&��6��tq�ճP�T{v�����b��˰��;Mve��ՠ �w1�<��7Sk�s�\��l�IԱ<[ۗ�9��;3�Q{��g$w)�4I��]�6���ʽ����944FQ5U�����ά�)Z�2��t����8�[ ���j	+���|oi��]A�)w�!�@��-��e��6��{��	�}I��n��ۋ�Qmg�
��P|x����H�r��i���>��b�F��CL��{��Nֵ��������aX��R��W3�'�mnK��z�u�z)b�����Kt.�c�̸9���g�X�겞�|�z�f�2f�j�X|���Π�>G��{\r�ѷ)R���Z����Zr���f9��n�}�}�y�hb]=G��د3v��;(�v�}6oj���U��Ē�*��!�͹ٌhΎ+W��3 �t:̻�)��-��
+��Z�u�����N��̋���v_��AZ�m�ū|��c3�WR#�mo44�WƬ�3 V7^��/�P,��n��>'置�7z�&57{�x��N�ų�0!"��ŉG��se�^�Uӂ���G�0u���nU�X���>�|�#Slf�_W)N��ǍW=���s��Q���b�X�(�.����ʯ�Ia�vA�.T(tu��t�坕�8��"O@F�d� ��J�rb�J������{��c��X��{��;�W�Rut� �������#E�&����.��n+�1yF���.˅�*.8�b��ݮ-�rH�vuӁ�.f���nƣ����p�[�FM�R��{QTUt	�/��"�e���u5�������K��Ȓ�%�ՠ`�,�G2��}��M;^�����!�=���N[N���oU�d� M��J�l�k�:�YMwU�]�oS=Gah�j龼*�l`Ԗ<!4�5�|���C]=��R��"��΄�(;�r/��·>��/�1�
D�:_V��Μ��I�+z\K����4p\�jdԸ#KP{Z�s"���(Ӣ�݁��_^/�.�#����csR�y{\��D˶�EGxa���}�5(��N�\T����R�.O�C���P�+*U�[�*����K���m*ʀK�e��tmV
@����Q�
�+D9˹��(��u���9�B�����C�Zs����+��Y��ʉ��v:����ޗ)�ȫ�$>�:6j�܀���om΄�����L��q��ǆu+��<Of�`�Ɩ��w]^ԕ��#|e�����6]���N�{[j�E[��&�o%��1�L��z�b�g]�=��uY}��آĬع��X���H�\��pt�]�L
��*�����)�s~FmX")�W��o)JV�޹.�)^�b.��3����F��X�Y���O�ͫ��%7{(w������r��)'�5P$�����	��u|���IaB���x��dv;�#s�|f��U�v4e�����e$�tò��k15Ł�GqF;&_Pb����ɺ�*t����T�:��;K�n����
7n�8(�V���Z�W;1%n�)����s�IQG%r\4n�ǻV	TC�K�x��k�xdAգ]G���y�]�I7�i��V�Pq[r�S�b�Q�*q��l�V��\���c0w4t���*=|ԫ��J�ae��v�� ���IY�O^����V����6R��e�6�U����O+���	����ZV���3y:�6��G����Gw�{�R)��Km����ʁK l|93��|oS�\�4pga����N�Mt��j
Q�:����0*�Z���(6Ez�nWw_q��A2�ա5��Q�����^VM�e��9�G0ކh�]}���1޳t�πv��bˈ�dpx�@�׃)wU�^b��a���ʋ�����2#o]��KvU�S7HT�b8�bke��m��\ܫ{u���@���OML��ҽ��]:�<�۰��ʚ[#��Gf�h^�i૦��kl�Mi�`�4!1�f5�����+9�u$������"�vs:�+�xB��'9��\��L���&�m�7�z��vV���ז��vj�Iش+p�6y-�B�T�G�oml�v���:\V�9�!����i���Sǚ�t֊�"�:#̽�!oMF��(
��d�Y�����2�;g*����u��f�5\60x��z)��k*uvi
��1}�\Ӥ���Z��d*7���VW���R�$Ռi|t�%6;؊������[ܮ5��u���Wk�!V��c7N.^JCmv��}5���GAc��YՆ!��a!���pܖ0ӽ�_1��3rt0;\��53L�WqM��������KN�TE_�wKiz���ϟ��zZ���U�k�7]ʢA�K�N�!�yG�M�f�1�z�f;l*���"9g��lJ�\��W:faz�9�ڜU<�r�9w���oF���unDe�J�˧�r㜬T<!�nr-f�o:���
����x��W�����.��ӢZ���AV^.�M_���1���+C�
�s�p�̚��7�4��u��H�&��k�Ec\�\��9���v鐤��ܫ�$u�4���qt�s�>�2`�+g;��N���t�F���]�d�$��9n\�{r��d���t]Z����X��`����tyj�V���ՙ�8�I+�u6���ˊ�ub%���<��V�$�7"�ռۦ��K�Q]F�̽2���`���۩R�ǝڔ��^<�Z��d{yj0L Z��Z!����_%9v:5{���orZ�<E�%|:K,����	�Q�¥��a˒u����Ҹ�&��C���\m�b�z�k�u,7��g2m�$|s�o���*�\�q���k�8���M�X��5�AP:oZ<%��zp`n�[�%��v����,�Dj]�'�nv'ׇ�)g3h���PE�jT5��$�i�,@�*�
\p9 Ox��n�AWN]�`ۘ���|�P�[8JЎ�4z�v�li�P�8J�ZRuw)g1f�_T;y���uS� �
���%i�L�Oۜ.��Y@gm�u:'?e[''.�v�n���R@���N$���P��S����
����h��ZV�j�{K�*����
�ۗJ�
����O:���=���8������]"�g)��͕aTO7��D*l�ٴ>	31̜�S���z�vwg,��Y�E��\떶�,�[r����G˸��v�ݲ!�Ľ�^�U���U�WK��r�/��;p�vn7��MmaM����XU� ���qݥkޮ�/������|�`��35ѻ�$����C�Q��9������f�:����G���T{�c��{�˻�8ꊻ����W����K����f�p�w5+�Y��}%���ne��N(A�e��vVG����[P�6������Y�N!���'
��Pf�-��mbb�oV5��^va�,���˓�G�'jN����W8m�{�H�kqT�� Dm��A�A�r�^��J�=c�s�Ty՘�f_�&#�}i��3|� �^v�C�6���^j�F�c��*�V����n
� E��pd�(P꘻O
��io~�8F��^7���Q3���ج�K�e���;S�Muӳ�H��R�U���V�/�����5�g�`q̺��a�Z7�Kw;��:�J��E/����q#��ue�O.��7P�0н� �$e=���Rc����8��5yC�mM��*���!�w�T�]�r}�؟q�m����y[u��8�|��
�5V��+���p�VR��m}���8�	��NK��F�efe*CF�����������1\�N�ӗ8+7��Gq�70�zO	�Y?pwU����X��|e.hM{̇��ፓ��V6����אQ�f8�m�"�k.�mrU�}�>��A��up�<P����ڂ���o �}��q�#n�������d���:Si]<pE�eڇD!�oVT����u�������J�b����]wgU�d�I�K��*E)�.��Y��%�����`�M�k�=�C���u�,�|�oe�vbE�q�˅�ѓ+�pɴ�l˲#�"��JX�2%�G�D�}JsH��	�'��1ٔc� ��yZ�^�|��<f�i6�;W����R&^e]:C8d�B�s�v��HM��ܮ*��kY҄o�rSI6���Xh�lC�v�V�EuC�g�]뭈��Q��W3���U�]����<;Ť�R<h^ �Z���2�J�J�÷AV��d�=�W��� �d�L�ٌ��q�47��9`�i
��4��4ٝ`7Ԫ��h�
��\�A�VZU�F
��mf�P2�Kӈ
#�EWt�]Z�ܞZ�BH̡����7P-=�u&�k:��t��׆�E���p�!l:V^��6WTT����]7JN�8A/���zw��K�xJi�*�&7���)k�������3�PT�9׺����2�}n���;���M��j뫅�R��9r�Sx��k��{���6(��f�v�5�U#wY��--����]oo*v�R+n_v *+%M6��n�rt,^��u�Ez;���g��N�G*�p�ʽ�ܬFE���}����&�/���c9~~�����-'E���n[�k1K7P�Pr��`:X�iGh	��&alA���xj6��VX�w�X�}h��lo �є� M7�⻘�����G3������\��i�2���ql�?�9YO/���^Z��Li"���k�
���d�3R���xG�h��gΟrW+_rP^Y���F����Z����j��%`��1RDI�
M+���!Q�Z-�9�k�#q���h���ҝ9�5�u��tZ�DV���
��}�t�vk^����2���j愙h]<4p(�[r_b��8�(���|�������;)��fj���%�1�����O�e�ƌ�#Y�,
�;E�y]��_����jŪά;X�p:sP�g���t�����k7�]�8����Ǵu#����ݠ�P��p,�aH��'���*u�b�NR�L��%��P��z�r�c�v8����i��/�k^���S���8T9��f���q�V6h��+��15:-����6�p�KEJ�=��ӚB)o<��q�:��.����5@^)�2+�e�XS��p��T9F�<_nBj�uf%A�=u���6s�ZC,����t�)�㹹�S�mf-�0VЉJ3���Ա���R�4�����P��f�l��V4���]I�y��Y"�C)��&Z�qea�8�\�C�9�W-����Nid�K���s ��hA��$�d����w�@�H�LNQ��e�FN���fܳ����3�=y�t]��[S��K�(��Ol9z��8������r|aG�,�+A�B�\r�Cz9���D�'rth���;���sI�4н4��&�m�sge�A�Ɔ���`S�O>8!���y�/lr�E��]�����[۷�n���R,��1��tҫ��_&&��hOU�Hj�],@��^F��xi註oJ���P�ӫ�v��-|�Kd	�}(^���w0�t�"ԫ��e#|�M�v7�}\�%[]7fw�Ɨ^-6�Ș�7��pyyK*<oo{:��}����I{Fsl�էs���Af�I9���݃z�D�e�Y��9de�R�3%��"���:QA´� nKN�逈;N�����a�ƪ�Ÿ�g��*����-S��Â���ѡ�4�1A�c-ѭY|�J�4�5���lҳAY{z�X���.i���Si[̥����%���=�w(l����h���F��t&P�ybe8�λ0-C�F&�w:`8x[�j^[q=��
H���Q�Z
�M܋�v��D["��߳���\�W��rf�۩r|�u#�&�km˼�}Y�E<u'�0�Xs�Kד(��p��]���o�R���έ5n\}�s��ɳtk�g5�U�.ok5���Qw'Ys_S�&î�76���|P�)��_f7�S�m��fp���eճ��ي]��o;����}C��h��N��}u܂�睪�W}}�r���J��!MBk���)��!���kn�Z��Z�W�\�`lr�|�I�.�0�k3�6-�h�*8��å�ݹ�]7���Ћ��TWe[���IM�ͻ�E��AI�a�_Z�24�TE�Y�D���A��Lea"���4�oc�N���Dc���li�Q���F�i�`�0*C�Q?oj�P6�Yf��ZXL]G9��iڹ��d|��WR���(�j�V1���v�q��/�!27�$ưԾ� �Wr��zH`�������g_@���7V�Ûʰ)�uMYӏ>Z�ٜubl #N��	�Y'�;�jV6�x֍�4V�g4h��y�O����Y��hӗ�����f𫇦$ ��Cn�.�=�L��c+��@7��Fc�.�����N౴������^�l�ln��Z�k�韥�8ᥢ�<�@*ީج�S���+*��ξ��t5�	:jJ�[L:�WLb���.	���ÙV�q��B�����f�y���y����/oiE��,��	�X)�J��rĹwAe݆2ҡ���ir��G{�C"��LZ�ӊ+@ǻ\k�ae����v^��>p�����mrrfyyHh��®�	�D�y}xf�&�C���ۺ�)X�\I�d�}�K��-����v+5[�L�Lje�f�q��4~xp�{%������e�����;!M��4^et��-CuHz�V/���^hQ�Gi'9j7�iUt����Dv�T(�̈́:?\���#]C{�
D�Z{r���u\ȱ�%+�����t�՛��5P�4��̜i�/�R@u���r�N�e�!-�9��e�V~�:(�=�X�4�*=|���
<~v�	�h��Mֵ��v�N^a}D�SA��εҌ��ҋ��a׃�8�1�Uu�ˬ����Vh�Ѻ-!u��U����ۂgy���`�Һv�6g��4�<%)C�I��qxA�T���]Z4&�jafCz#Z���(����r�;Uv�1$jU�CD''fvXC�:3�6�j� ]K[�Y���W+a��̳��pr�F���mr��]©�.��xA���J��Yg;�k�(9/�܎�p��-f��@�=N��{��ʻ�t���G�`�����M���v��z8�3��X;vG�v��5.��v�o:���os<�Jw����+pP��G�Z�GȺ׻���d��;��.����Rg΃s��\x�v�h�0�8Q�z��V���D�]S�:��;2�x���W��d�O:v%6�Mv3a�9ԝ
N��Xh��,=w��A�&���V2؜q�p��⥶���(���:�v�i>X"��ہ�͎��A�B��7�x�`kfYJ�#���H�u>˺7�2�%֮K]�ԪV�3�^�:+Z b[ult��tN�B�a��n�iL����8w,��T�r����<˽@M���ߊ��[��?M�[�'==��tY��SWQ�.�T��F#ӆU՘l�7�o����.v'}-����%��>�e�ܑQ7>���vZ��p�6�%E^s�2(M�fWt�L�/������˲�����5èhޏ�,�m�T��0��x2I��������3W6/F�f�R�'�����8���p���]!
���N)]����I!ٵ�E�5Ȋ[�a��l�Ȍ:�о)���:,�k���wg+;Pmbh�	�)%�6w�TZ��7:ے�#l5t�Jڂ���Ᾰ�.�B�a�xoIh%�]��u^=��R���X麏6kyB��<6�
��zO:��>b��s��X|dz���CủJ�|L f3jC}I��\���'�R�`��®�*�|�;r�n;�u�f�n�x�,���V:���ճV�,�щP¨f�.�9�
�*d�f4�͚�b��.����׏�]jfA#�cK�ӷ�]L��5 b�)b�{q�5�"�b��� lзm'ڳxk��䂳eCC5mryaN�[�b�t�·^��𥻽[�\$����R�����][��]wwN�M���[�RT���8�J��A]��4OQj�~}��q#��Vۙ�+]7Hz3(�װ�)��*\��7X�=Y���㫮�nP��M�Xo��"�­L��m�k9��[���AW�u�W5ۺ죽�)r/�x�С�^��d�?�^��m��NuM�՛l�E��S��`�N�5D0`V#��rBɷ�/l�d��M�4�j���S&䖝ru+�Q�����j84��5�-��k#) �u^T#[��]b���F��-l�讣vh�����H�tvP�廠I��S}���������o.��(�6�󰲇ob#�ˋY���l�|��jq(�	2�p����A�ʀQAH��\��I��3`G��-,:^����)��UZZA��]X�>�-֥�.����6�
<�,l'%Hy�8-��.�ל�\�:��}�),Do��w��&�ͨwM\�UfN�v��v>��F�p��]
�-�1e��J�R�����;g��\[�\���i��n�QW}�@-�ut���|�ǆq�B��JG�N�*�P%Q���4��{33��>j-Tq+tS[�GGv��˷a�ξlN��̊��5������0Y�2���T��6q�%��eiq�P��v6AY�wt�=�Et�M����]��CW�]V��:�Wz҄)pª\�2���9��I�V���lF-6�S#X�<�z���!YE�w31�İ��.=7��.�=���Z�L�zv=7����aa��\��9�#�@nR���۵�$��^H�V�G>Y��w�z�hv����IwV�۩�V��� Q�2'��7C�u��%b�wju��oP�v���(�K�k-���ț������#\�n�M�F�C^v���Q��Yzk��,��lo�:a�G5�s�7��^S�+"��ZY���y��f���Kh]-��#8��j�EW��d�����-�'_L��3&��Ɍr'x����īrH�1�g�����L͔tmNv�*X��3"i�n�J��f02r�.�������h�.�RP�r�P:s#wˍ��ˑ�Z])����*�m���]8Q�j���� a��ՑR)�ffU�/��L-�.��eX�,2%,�mݾς�"4��&S,��	��ęK�əj�NBe[44�V�{|�Wsc�J'n�3j�����s�Me+�wK��e��:'�6��[\�J�ÃCvJVܿ�\�k��6�^Mj0Ӗw6�)6��1�s"\�� ����uիf]ZJ��Ͷ���K��m����W7�����e���6��R�ދ�HծJ�I�t�$$���3�S�U�[���`���g�˓��ܺ�K��zFf*�+R�]O�^�iۢ���ҭ�Z�xV�]cV4��^�����.���@�y�[q���L+<�s`�ܦ�k�N���t46l*�Y�鶪ӝԳ�o9%u���ܦi��"u]vK��:j�U�Q�]d�C�fp������+�%��&���nz&��wfr�8a�{���9�C�J���x�\V0"J�٢�5��/x=�6��V�9sw�,+o_l7��j
Ǜy7���Oj~��:ȹ��*��j;�������Z}1[�8�ܷ7�!���8��u>a=�x�9Q������r:�:�G�{(�ٕU�����T��ܽS�����������E��펹eThr7�s���e�Z!9U�^�%�i����+����*�a@�r�ț�3p
#C���4Շ�]]ZA��+y��Cy��mIF���y��/�G�=6S����}�HhC�V���Q���c
�	Mi�<h���+tvҤ7�����á�Q��'��G51��i�ܺ|�/��P��?. ��U��r�M\����0^�� �We�X��R�+���Q�<�7V�]��.�Ѯ���[L�0�;W
�R�01Ւ�ur�eB�^�Ɛ�T0��4��_�H���7�i1�)&��b��َ�9��4�t�j���9Sz�rN�i��Ʒ�E*\�fdє4����C.WDf4�5��9.�J�g[t9M�X���=�r��kb1��HY�Ɓ����+���K��%.ۄ��r�y}|MBz��y��pT�:�AՓpil+����|��Z�h����aD{N���Ya&�Vm�����q*}�q՟s��:̡$��J+�n�� ����92���t�E«��SL9832����̬w*u^���޵�c��XE�'}�T��P:k_6��v,+��^B1^Q#���Mk���W}��h��ח�Eԗ2��M���<j��&�P���#tr����ݭ��U}�Kq2�:�^�QT�N�U��uLte���qZv����]�dm]
�j�L�ݝ�m�9K]���:��8��ź�ӏ_P�em.����Ȯ�1���$�|�bmj�o�-����H���Ƙ��21�k���
i�o3�#��UΕY�l.*ㆰ��=�P�Etz�uU��0�־C�W�lY�
��a�8)�[,��Zڴ;�����Η��
�*WT$ -��ͫwQ	��.�L^	��ӣC�"�(a��ɮ�:Y��Y�=��a�Uh>�W��%�m�����o{T7+��t��串v��7�N�zWlCxM�B�͎�sk���z5F���n���ݛx
c��5�[�����R6�m�ِ�ܜر��s�f�0�ioTF�ma�'}�^Q2mgΥf�`�;�
�.���9�j��ľpɐ*ok�f���+6�d�u�]��J�dՂ�[�8v$k&�a]?)����lCLbV���M&���aqګ��!�%�"�&�/���_^���sAs���jdk���ă�D�3:��^Ny�X���V6g<��9u�?�Y���{�������X�uZ�r��iG�j�@��.�2�m9%��5)w����l�������2�P���}HJ�8l�X�0o���AS/��̇�
�
 �ط�x�����t�dM��:����,f�G7c����4�P.�gK�i�l��?�
vm���C�hEN��n�.hֵ��;��0�;s x�T�ӏ��I ���
WuusU(�5�+�8%XF�0�/����-�]vi�i��w�;���:4��W%D�;��=�^��z�b��K�:���Y#�8�/��U��MLt���muYF�d�ƀ�𚽧]o
�*4EY܆�����E�gZ����0�+cΕ˄�rVr҃:���'	{�����9�m�脊�wċK�}������H�  �A�����ģv!�k�ߌk:8Ūf�Z[�oE<X��ۡS�[V�ʼ;z����s��(���W9h� �����x��Зd@;۸
}��X�	K�X_[4�s�'�gp�VME����0J9��l��DE���4�P�8[F.Q�FØ3j
��՝�[�쿐�tX�l�E1V�Wq]X&���i�˱���f�lo���M��mkر^����]d�[��������Y�HB��)Z��,�V�;+m�SB�f�pZC��2A��݃���j���b��T�]Ն�Aێ��ޞ�|?ߕ>�WϮ��T��痂Rj��qb
���6S�{#�pYQc���h������qN}���]�Kv��ײ,��J7�j�h.pwj����N
�
5�
Ĺbe�b̚z�[I]���;BSIH���wF%hI�d��C��.Y�,g*gm����*��-X�)�vjg;ŦZ�}���#4�������B��oP��@(���5uc8��Bf-=5t��~���^���<5�~�]T, �ʋ%�V���<Ñ$�=�t��N�ny8Q�$�ա�y�`Lȫ�"u
�[��9!��;�����N����=�c��7Pqu�8�&IaW�║�u#-Z�W�J��f8P��Rs�*9���#�sB�E��r:�	2�S�Q���;��.VNN9�8��I��G�܃F�'��*w1f�'�]#�t�r\\"�g�\ۨ�O1rD�\t']�u8�{���9k���';�<H�3��X�Z�����F!y��"�Vܨ
)�2�.���uȳ��.�������S�r�DG�N\�Q8�I4�q
%U%A!$�.���FT\Ԋ)Zˤ�eFe�I˔�*�LU5e�hBNBw �,�d\�9�QQh�S.�fqdkC��ʝI�$��ib�_�J��������:�(�r��p�, +{�6](�@)n��A�C�2�j�ُ�s}�o���Z�h�a}�Vl*���>�������yJ�H����Bk�Ь|v�c���r�*Lw����F�0N}�3?����������ˬ��!Y��aV�+W�P"���}�r|CD��� J�L����HB�����lI�1s'�M���O�O�j�������Q1;��.@^�� ;=0n�^^�B�m�a>��,�<e�5��=*���A�*\�QHI�*������p���B-9�~�ܭ��5B0�B��r�O�t��/�)�z� u?;��`#US��G��l��*<,}F��{N
�i �v�Y�	�S�q�ొ�A�7�q.Ě�k�Kf�D��{ё&��x�/�y>���,�
T8xG|����X���[~�����j�덅ݏJ���Ҷ���M����'�������/�fW�g$'�k��Ur�d@-7X��|�v�~��I҉��X�@큇Ϊ��Ě9�/5�\�IS%��E���t���+%*Q����e��u�8�������j���p����וa0a۠
@�Ku���:�e��"�+uZpKl4�v�=iV�J��s���
Є�7��/�W�p����
4߬n�k[S��6��6�\��� ��,���\�3���Mg�=�N_ט4^)�]�7��S��@�D�T`9����u�Vr���8t@iA���8���(�����V��#�B�b#:�~LlM���ԥZ���k��-ozc*��������e�|�"̱ j��<t{*����&�s`����䬭^N�g�Y�+镳"��@�7L\�0�;����� W>VG�3闛:\�#	�0��?at�\D��SFT�v��%s
�P&���y�ٕx���nk}V�"�AR����&M+�Ο��i���^T��������������*`ؼ�IG�
��/�g���w� �R�]|���׍��5���չS���ZZ�Y�x�u�a������\�������v��sU�inp��MX�81����K':�ϝ6!�~YS�cjL,������3D*��,y�S�ԍ
Ǜ)X!�J#������-"���������1.7��!����ۼY�{1x�p"+����T�����Qڕƪ��zT�yx�9t���cwn=`?�snD<+Ñ���t���"�`����Yȹ^f	t����k����H �?O�*�
�w�W��g��V���]��z�@0�uo���Mo6�=]c;��Ѓ&Y��i�
�������	�*ࡦ�]��]���z)�f��֔��+�eՁQg��Y5����u�tR�֊u�8�ӂ�Z_�/ocSݹ�� �C����U�M��i�KExG����E��asw@��f-Y `;1�\��|�Ǝ���y�
��n�ڸ�k7n4y���9Z�p��d�,��ڌPWVP�7�/$*��b���t�X��� �v���guz��r�:ǳ�+�>-o�#�-��F�xܦ��.�!?b������R����b(B�a|L�N��<��O�s��p�iw�0[��<Y�'Et<�� �\�cڒ�V��#G7�(�2{.m���4-��>}2Z��n�.�@����<���d��� �G��L�=�j��MX�줹�ϸU�{�:Z@/S])�7��3uvЫ���^l
T�<����!9f�FJ�a��ћ{z%�l�n�g({���	�zg�p�Sh���A�"tzCr��EZǺ���>Z����Zz���"=���MjvR)�=�WH��5oU�h��}N>F=�[��b��C�`ǕSl��]��3����%_�D�L�.���I��-A?K&�7UB���@Ճ���[��
�#�@p��L:�D�\@���|.����EM!�����k��\d�3{,
� ǥ�0/Jr��8�_l�@��"$��g�9��d�%��|�Yj�� Z�<PB�B�}�6$pB{y��]x��E��xnW�Һ�xU�{}l��8�[�����\������Z{W�/!�Ե:y!Ml���.}JkuБ�SK�8�bZ+<P�O03��L��'��y��+�U���}�.���r�0
�B�vHNn
*q���c�6��cwu�y�]�p�<b�U��m�mǕ�9+������?]��`�`-SR̗�����F��0���wj�6b�*�7��ۭ�|j��Y�I(����*�Ln���b�zc�sjO?aez͎�t����t�} ����X��[��hｆn+��a���z���J�L��L�U��Ux�y͍�-�9s�M��>c������r��ճ}��r�~`�����ڍp��q��EΪ��U�O��Q�w��yF��K��oь�a�D��:=<��Y��z��m{2����?Y�z{.��Uo�� ]����M�&�6h���q=>��^�I��|�O�y7HD����+[�����s���h�Vw��&������Y~�/�J<c����� E�`	�[�fΑ����8I�y���#:��7���fŏ5B�>�a���| ��1"B�/i���3����o���kq�c�	j.�Lb�����ȏ"��HI�"ߜ��w�>m*՞�G"�Xtv�p�J�0�f��Q��n��O=o�HF f�̖�L�mY�MG�dz����e��t��ª̻T�R*�3�MD����<�f�93B9�Fj�)EQ�ˁec���R�B�Υ�WfG�����j���[���B�u�L'y���XW1:�)�u�f4�t�nR��N��l|��,�덇������Nm��བ�M[�<�[�l� VS�������J�u|O%�<�AW�*�Œ������U㞷�= ?yW�ʧ��}��:�n��`��S��u{%t����\(��'��������h#�����R�j�)	��q ��ł��.oJy<��;����7��*ҩ~4���Lu��{fb���eK���@=��أ穹Y��1:w�.`�/�kx�=ƞ4f��$����`���g�m��]��B����}�2��8��u���=QV�U��^����z�E���U������n`��p�$)�Ɉ��������JZ���i�U߻���?�6|'/�5���(̧6�9b�
�f���P���� �;������vg���`d��Ͻ��E^Q�i�9�Q���^������Ҕw��.��V�g#Q���3X�@[�̨:���"Y��S!kj��X�`�D��r��34��+2�ty�V�4!�p����i��j�ӗ-Qik}��᫫���*��b`w�n�V֦��z��Me*�k�*���]#���|�u�^D9�X5�Wژ 9����*w���׬]/�K"��A�l�00�0F�d�ׁ�z����ho"R��: �uƳT5Z8*�c�ԏ���}����k�7=�w��=?8���d:=�ȅ^���10��uk�/��Tn���������hp:8�x���S���+tK�k�:���{6��og��:.E�{N����B�l�#1:�����b��0;��zjhY=q�U����,��K�aƲ=1��:��S�!ޕS�ƣ�E1���{qv����==hp詏�V{O��R�x|�{_ǆ)�������-��E
w�Q���C�ZU�ĸo�Wq�Hw�kEh��B��_���y����X�?7B���U�tT��q�0��ՍV��R�8��ծ���@읙��3VR��1�6їu���N�C�3gp�Җqy K$�h�0�'�$�اQU�y�g�N[LՋ�b���$��_���-Nӌ��+�Y���ذ������nWE.�|d�ƆJ�Ǣ��1��N�c���D�͠c'/4����`��ƴ*�O�h���4�-_[<2�d�b;RMxuq�MW�xI�o����;���ba���7�1��h�p�Dd�B5��^�����Z�f7�@�Pqf=P]`b0B��SWE
D�2��a��#l1�Բ�0E���u䏻����<�)���T�ȩ���ǕЪ¹�8W  ��'Ŭi���u�:8�<*�V��{g����Wq= w��(�]� �̩��7���[�8�A�k�auZ����`}��4p�P�a�����BQ�ɽS�4b�l�� ����xGH�ܤSOm��Wl�Zj
0��_;��J���{_U�I�p4)�@ft��#�pB�1�,�ZF~��i>���L�R�a����P�>�|@�R�y��W�0/�G�����=�7w�����0�}�R��
TA��f�Njf�:(AZ@�|�"�$�H��d��F;>36���7�ҋcw(2-׳����5�v;9���T�οqa�����*�g����2=���q�Oo��T�d�{}�w�8�u�h/y�82C*���Lu�u��i��\���`aj@��W7��$�9�ؕ�PV�Ά�੥<o�#ݿZ??
���yw�<GɉyMr�KJ �y���حUr��b�vx}R�� �Q,yN}�t|�N���nZT���֎ͅ^�?�Zv��f�f�T��hΝ����q3�ut�T+����mvL��5�ゕa�ݧ���
C9k{+n<f�X�kj�r�k��7�1��8{��4��PS��ĳP/��
�$h��(t�<��yAX�{�x�W���9I���w�ZعIt5=��h�~�\���qu:�\��X7�z{�nb�5=��.h���ьd��:9�X�o>5}f�`���;��ѕ{�u��}*�Q�Q6Fi�F�=�&�6K�_^���W�	�Ӓy�v{�ɽt_Ƽ ���ވ~�<�����!}g|l�՟!^WW�0�W���H�C3�i�+�Yg.5~�^we���q�YХ��K;�9,S'{Zo�4��W�F��e����鋰 �GgL���7|����_mmwY���E�&䇰n�)ZkAR�Xz�m��z�(<�)v�@zR��K,��ch����P�ds@��j��:�{�Y}`����G�����{��/=^0�lhZA�ޘ
`�pX�K� �$H-�.7E5U�����[>	�LP˚b�}u�P�"A�.Y���.�Ɋ��~�G_UY���^?r��C�pT}n�MJ�0�e�|�(�Z�S�S��]�ڻ�[��.���Qv�I�<�KP:�R�t�8M��u�X+���p��2�=���	׶.ۀ�]�?]���'�էpӮ,��}��v:�1r)W�ꋘ�8�~�y+����p���@�W*�/�yXu�l�uڬ]�o�'��?{����x<u1k����FF���Xk��o�{5!>�\6�3�v�Y۽����PWG��\�Wr�h�и}��U�Z<�}�x!�a��}��Uv�EXQ'�����s�{�U È����EL ��Y�4��Ƈ���oJq?R������O߇х�~�=Q���hs����V��ӹN#��A�3��2:�Q�'X���x�F���U��j��.��@�l"�҆f���A�մI�#̙,4Jw�*���De��V��,���K�c �{@��]I�U��z�]��y(�|�1�z��%e�t��U)V��ه:C�l��-sV�K����η��2֊��H�]�f����ãz"Ϲ.V*�3���c��h՝�,�r�[�� (Xý|p�S; *r1��P�ZOpt;�՟���+5�MZ�İ�-l�H�{O����ڼ��B�,\$���Ml̿�>Z+ �̪Qo�ݖ�_Y)��e	���8n�{����m-窹������]�]�/GL�X��\X�gK�NS��j��M��<�ևQ��D�O
�����	S�5����k2s[�reLĪΊY/>W��&��5��%_�U�Pm�7]�o�:�Q]ꭳ�CAL���A�&r�}�h��Kጠ3�vtv�\%^�(���	��(�Gts�f_'���n��Q#v�۳ʢٰ���h94��}�;,��Vذ�G�aγ]Ft]����,E��9�� �N��]uln���D;sR��JhH���v5���6J�y��V����~{�!�Û @6s�gj��+(��q��zx�
�(;:��B���Z��aA�vq{՝V��c�՟X�8�t��"�QǻJ���\N��r���b\�7�������|{9�G�mx懘��u��,��KTW��Ť��T�o��ψ��.�֞��.���j��L%:;}�ڨ�a=��Ģxn:it
j�[�d�0�&< l͙�"x�}�p�Ù�>�㶔D�L�\:�:o���а�[}x�R��-ܜ������,1H&��%��D����]����'Q�n`�?���,��{�ܑ��־�7�hG�nLD�Spv�eH����͹0!�����|R�L���s�W������垱V9`��8S}����{h��5�����e	]���7x�uL�\#�|{�sZl5�u�N���U�����ѵ�3(�x3袾V�Rt�y�ks��WZ�e��0Y��m@�Y�m�d;��@VŹ�$���}kDd\��]��f	�@���&�+�PĨ�K3p���,&H���(U�uԮ0YՌحt�;�f�b]�I5�=؟r�in�V_.��S�=��--qͣ����L�A�
΃��ځ�F��Ć;��c�fbl��}Wd*�t��$5��?�K>�T�$�>#�� �'
�BT �jT]d%Q�L�)S3%:�,�#K��EL�HU���.]!39T'
���&�Br$�ˤ�Ċ�$ˤQ�J�/���*����Z������1(4U"�*�l�r�J�!b	�(��E$�I��D�FJ	����b�ʬ��E�j!(�4��sV�ΐ��(�"�J�s4��+h���Q�g.%F%ʥ�1P����E�i�'(�X�Rt��SI�IT��+S�\�R&�LJ+�t�()dQS
"
�\(���!	bb�!u<�n��?��5�Nt�십͌�V�V#���#�5��p�} |���w�ϝ���yL*���&��w&�����d߉���ǔ)8?��=��P$��G�<*\I�����0�����W��$��Sxw봇�ׯ�$+ޡ~f��tEB!��@���D}�N��u�������Ƿ��0��~���o�*���W�q�?S��탟	�����S���y�;����>�3�B>� ���F�����tI������P�L?�rr
av�}���ސ�����(�w�i_O�M�	��݉�����wߝ�!!�9���<e��
������W���������$`��ot7YG�}cw;z�z,}D�=$�	ߩ�<璘��<&q��ro�N��=�|Nq�'ӷ��iӿ_��y@�����+���N��HI��~�r}�M�>�"�>}��_���_|}�����?qΝ�e�I< J�~��7��	�������C��)�0�ۏ��巗�xL/���"o����?M���������j��>�DDH���e=�9~�Z�u��4��.$>�Ǆ90��������0�}O>�pzM;���F���J��V97�'ӷ��890����}q?_I��]��|yS~����\��{7��WӅ+{T�F� ���진)!�5[����yO)�S~��yBL/��z��
aC�iɽ!'>�x���'^7�����y���Ǉ��9���＾?_<{^�FƏye����DCA}�B����i�y�xW��~�܇�����}�����<�����奔^~x��O	�]��A�<&��	���}D`""�}#�b�/I�+� ���^���ϴ܁��ϖ��
���i���}B|'�n�����NO����Nӏ'�'��	]�|����7�'ۂ������gt�,�����W��n�_�]�{�r�Z٩�P��38�Y�W&�ӹ��`���|O�r�����@�����J��y� ���=��]�{���94�.���NC�iS�w���i	�
?}��/k��W�~��82���Lx��X��.ʏ��G�]SE��
����j�}�m���Z;�-�.�\�G����L� ������>{՚n�%叢M�sE�%��C7k[H��3XU��M��Q�<H9��~R��H񭬔n�g�*I���L8>��>��ߐ���a}~��o	&�y]��&�_��<�@����v����>k�ސ��y��?�av��7�����ǅ�q �v������>��<ݪ���et|�D`��xC�)��>��N96���o>��]��~;���8V�[3D"N��t�$��[��˽CM���ooe���)h|ji-s�C���KD'��߫w��Z=�vn���yo^Z���R5+w�*">qoʁV�_>Y�U�����ʈ	�>�ź�E(m.�g�l��Is�@�5����U��3A5�%�t�>OǷ��u�ՑR�ܬ8t|�+Ϟ��1ά�;�����S���J0y"zs�x�Z=𩇂u�T�k���c��*5�L���úY�z��]�y?S�H��Z|�`i���߼�TL�COY��|������n�.���W {2�x�^t�e����Y�ls_w�]�si_��7fn��`k�������(d����*�B��*�֡�7'�5���ċ�!|�<�[:ޥS�.6��Dq��z�-���8/:�� �M��;��d��:��QUҽ��)-���t�kd=,g�������jǥ7��*��{�����-m{Y)�l� 5�j}���4�,r�o�%�Sn��\T�Pq�o�ً�`>�߻)���x�8�4�^��:���RS��L/zu�y�R>�wN�P��B��꨺7Q��24��;q��%���y�'�4��֢�h>���_�w�p/�X
R�~Z��o��yN��$�����2��s�D�}�6D�z����,�����Ge�����~�z�g��P|��s|e��7��|�a�u_�)�I�p|���=��������Ε6G��ͭ7�h��;Ş����fq��ֶ�@+�Pήt�h�4|�/WsWޢEh��|{������Ϻ*}�f+J�z���ɮ���HE�eb�Z7��r�/;$�͔V��p�`F���1N�5n���o�D�94�)���=έ>��C��@j}@P,��qb��S�o5�θe�II���AK�����E���!M���Q�[X<����P��:a��3��=��S�ڕ���#��O"��6o���W�+���%�{�ӑ�v��U5ߵ�>W��3=6�p��Rf�T5nMD*����ھ�*�X;ܯz8%WM����G��ٍn`7bS�Q$��慁A��_���;y;>chÇ8Ɇ��8xJ��a�L�p1�(�rw�V�ǫ*�}��H�zB-�0�sNI��=�J��h{�)�����$��ٜFx@Iߗ��ۘe�FBa�)�TT�{|���ͺݷ3&5!c�Ҫd�b~��lN�|��j����̳�y��՟R��+r�Lb�s�����.�h�]]�\9R�	ǡ�yҨk:mm
YIJ�1��q���r�t��zn�Z���>��
��|I�T�7{:����S�0r:�ٚn�p7��gL�i�j�Ѵ-V+K�ݏM>��l��LG������w�����#b��? %nN��{3�y��e
{�0�P���]��ȥ��������q��	��߁�ƻ���WO<پ�����^v����2Nq@�[5��]������T�cү���^h��s�����\��gw�{Z=p�T�Hy��}�.�U��b�<{�bk�h��I���:.Fx�^y��]x���MI��Uc�sh�=�7Bf�[���#��R�m�T}{f�:�+Ʉ�&5z�,�����>V�=�x�^o��d�	���V�Q���j�b̓���n,=����J�@f��boH������/g�c�&��	���J���TLRb<���"ᢺ�mgV}�Wa���F95{�a�k؇��+����ޅT٤;�ʛ�����$q:���ae�_��_�jܛ���XlZR�qr���	�H."�;�?yf��Owm<8=v�i�$���.+R�ZU�+85��m�����ܭ*���Uw��;RU#y�u�'t�?U[�{�f���fo��xU�"r��ڕď���,�n��h*�4~��f[܀����]Y�`!j^̉���Ϋ�/X�Jz��{מ�yݎv�݈ϭZָ-�����L걳Oc���b5D���X�w�w��`r�ݝ�`L�^c�圅��;C�JR���!O�*w�xE���䊬�a�Q5q���B_�&�z�{!��}8<�)?];8�K�o:A{q,ó�������૲�g��:x����h1m���Ы0�O÷�Kf�k�YH���+zd���C(V����5ٛB�z��y�/ġ��0����*�����p���{��e��'3��2{o�O&�-��c}���VWp���W�H�
��b���%ޥ� �$����<r�wr��J��Y��$-JW}��hO=��˒(Թػ�3>���.4����
��0^#Z���v���c��bt�z8���r5m$��89/|=�R��}5�/PZ�׭	�>�nyd͠�.��i��{�8W�o��kwr��G�bf���w��꾐%w�N�E�O���g�Q�u�СeΊ�RA��5�q~K%V�p������	Ֆ���/k^�\{d�Z����ӌ�5�%�����kk�O�9����I�{��'�Wz�c�N0���*q=13oZ'=�;d-Oh[�[�N^��Õ%:^ V;�]9ڔ�ަ��X�7���]�<uQ?iP|��}��\����g�fX^�qw_�~l�=�X���.4�J^~/���3>eI��NzR�!��jCg�<�i�|��8yM�©]���Q;gkr�CsՋ�(t<p>�zh�C0�J�j�kӐ{ZI/��XDˡ3;�8�Mo�;�w+y݊s=�X아�zz']!S�`����@�U��v�G�71$sHpiu/:��N��ت� U�S����>��;S��]��Yy��U+l<��.��?59*U�Mv�ڞ�I9yVr��3[]�.��������k�Q=�������e�ץ@�z�_ZO���^�y�5��|8V�N��%��}�3��}H�݋|�^�$�^����46K�ߥQ�[7��\�'ǖ���T�߽��k�L��財�p��j�F�����7�ڙu9�䝪^)��2ߤ�~��n�y����65T@��*Ƞ�ᶂu8\{�Ϩk�
=�6�RbN�ڀ�����/&*=Sj��'��qz������~t��Ҝۑ��-�3��oZ�7�+���ۡq�+]�4�B0�3
[���1�ݥ{���|5j���h�����z�w
w.����gmt+���G"�Ǉ��� �v��ŗ%0�~�=��R�(ky	��a*C�(����Һ�G#�;���4:��R��Nď���_f�Y��L�o���cK���7��6����޿�֠!����W7��噵=sj��L�Ѻ.���d�"Ĥ*,Jj"�����s��+�9ox{=4�J�+��Dj�۫ڳ8W<)�-:�{�9C����9���vV��Rb^��ZM��C�dA��j��N�j�!z��^��>p�,�M�w�g{Ϥ�*�<���Ϝ���w(�x<	�}���V�����K}޻u��}<�TyV��@�!n^S�KG�w�n����<T�֫j����O-i�<����_VL9�z�+G������]��U�9�O�W�דCQ
ZbD
�z�V1ū+�j��N�9ew���j��m�-�B�[��\�H�Ca��/��zRٴ�H�la�W\�!�ǹ|̛�'`�jS�b�S\�9v�\2g|�V�v�v��ĝ�s1V8�]Ӹ��/:�5Ώu��8�EZ��ʓ����7÷w��T�k5��+
�Q��&S�PՉ��3ڜ`�0?<�.z� _m><h1V��G�1�B��}��닡��t�Y�.6�?gFTLF<��v7-��(�+dz}��~gɶw ��By���J�z�lN:`�`��g>x��e(ew�gP>����n�=��L��{j���bN���l��]8���kA▨9��3*�؇��5Z��eZçfG�~��L�=j%U�pu�a�0�^axx��������k�hߤ�ϩ#��VT�ϟ��jf�/N��7o<���EW��p%o�����^�>�]��9۪���onL��K�C���x��z��٣�8���g����v� r�e��<à�̆�D�f���9����������H�L�%�D$��r�w�����V_r��vaёG��'&���7KW��a��b�^\��u�CV��4�k9|����WI��j5lbĞ؊�m#�A���U��F���+*E%�yr���U2�Hm*V2h�A�b�W$�YFt���֭����+<hiX�¡l�O��
�uÇ[���?t�����A�IP���,�ݎu*��k����D�`3.L�cG���NR^V��u(I���7�J��=���c�k�.�\�u9=6��l���6�S��%�.���D�Ӊ�:�e,结���+ �R�Oe��K��}vt���̝
�p#�l5|K���';�+�F�,��	��.����s�1�c bWM5+��y#�-f�<�@Z�vk��9��֥̔6���0&�=�J3r%�d�S��d�f��%�V1����!�ߞ��0VOٔ�ـ*��-�%j��.��(X��XR�}|��z�3$;��E���k�Ve0�`d˷�'���<ෳ����y] 7,ӝ{��E7(�`���S6W.	e$ȣ�5�Ė��r����=Ի��P-,v�²��.�t9��w,FAK���&|����\�4�N�J����'����թ��t�kDU�;{_���-6�ʮ�JC=�T=������;'cޣsXmԀ��h&�,&S*�{�@��1q��8闟v����H(�f�gU���7%��Z��Q��}�z�����	7���������$q̊�[ݣЬ����#��n��"�ƩR��d�HS��i��;77�جW�ɕ�S:�w�v�¬{���O*�:3K�悙H^�������gɔ��M���h��k�5�_6��VJ 5�O22jB]��n��v��i��)���.6���(p̽��qA]�SS;���M��ݣn�:�������b�S:�%�AS��;Q��d6ŇX<]��f
�p�+�����Ze��lʼ_mRo�<�(�r��uú� �����������]�53%o6B����9��V�x2�/%�Q�Qf��e�. ι,��|
5vh,�@J�Ź�T�GZ�!�3��S9�Y�ʤ�s��PF�,�tmkN��]FK���{�ܑ5����`3Q)t��q�5���e�t���W[v�S�=�+�>����������OG��#J��I՛���Q3L��GM��g5ZPUDA	�ja$��ijh�����b'�J�$թ,�&aYr�B-",J��E1VS(�:���T����
X(RdhTh�g1.���(�%��%)�Ha��ZRd����%Vgkj+�J�:ba�"3T���2�ʬ�,Sm"��3br4T�Q	E��S)2�fH���HhFV$�%tT"��6�Z*Ĉ��r�*;"��QeL��*蚈b�]QCmZ��h Vd�I�B�����@�Ve!�R�r�1d&�UV�(��t��?�qSK}�J<�������ݙ���g��/E��F�&�R���7Ct�M���밮d���}U��x͞���o��f�	�X����ʋ��;Fz~RTY��x~�$]O}�@��x�՝1�6*ѵ������z!=��sس�z��3(?�1��zT��W3[�C�E���?+kf�ރ׬�vf�]&TWm��}�I��%;Լ��i�����~}�Sy5Ȯ�UZ̝~�^^�50ȱ��UQ�:�����z���R��3梠ߟ�bu��9��f&��UCh�U[�̨z�7Jːt;���C��yS��g��W{6{�B'c��,f=�k���)���z�D3�T8�e0\$�Lɷ�Deڥ>�j��xf�Ղ�zbroY��i�*Z���K�|��nqW`x�5{��3J�y�[JA��!�+5e]�\��bk��e��FԄ�V������ե �4s2p_L#�Ӽ�ʏ��X�YĮ'�L�5�.D��Ͷ2*�ƃ���4�gs]��̠��}.lc������t�-�h�?_xM�e�
3ɇQLy:���}O�_���x	2�z�0yИ��:��F�|��jg�mj�K2ٖޜ����P���\�ߟ��H�G��S���(z��W�Z���j���мTmʸ��j6�=lL{|M�����Yz�SJ�U��KkB�{��#>�g���(�'�=K"�Y˰�Oi��3f�U���m�^����'�Q��b��
9��["��<6.���/�bcwʦ�ͯ39{�����>�-�O3�	�|�Q�����צ�]<c�{��e{�Qg���~{�L����z�8f.V��݄��Q�z��ƛ����g�=����^�huvlؽ|v7�f턔�.�T*��P��v��7U@uR��s�������w:����x��]ٜٗ�;�ٜ��γ/�����j����&NǼ�5��#�ui��k̢�j�[�Ε�؝ėﾏ���l�*�Z�Vt������w*8{��>Y��?lA�b�3o�t�ˑLj0��eP���nb�1S+�����R����G��8��ݼ�w3'[�;������]^ 侖Mex%[O�wi�T&6��^gr��F��{&�F�Z�D3��M���AnAN7p����R�`+�ƫ���R�����W��|)���󙖷ǗUL��޵>��/�����8VO��5����k�Cy���ϋ�H�8��B�����jsR"$���&<���BV�-r<+%�}�{^�铞H^��f2]��b��U��F6�Iz^#�_���w�׫yi���:>�v�����8�~�?z;�aQ��rW�e�
�H�ދ��3(W}��{���a�o,�W�g)$r�
�S�Z}܋ǻt�Btۼx�AWCe����o#�,\����q�]ˬ��IЮT+1��|w���y��7�Xs6:ZŨ�%��꯾���+�wzN�Q��iv3ƃ�<ᾞ��
��!0�����|t��D}�ׇ��*�V��Qj�����2x1�~3*�[����9И$���O=�7�R
��V�NA[A��)�4�w�rz��x��ܗ[u�ӫo��\�m�s�U��n�x��,���LM��0�����u(��MCU7UR�C`^Z���o�� >��V����mN�����I�ι>��xNv4B*=��(���;ۀ�llţ���_�&u\����Lo���wL�����|���^N;F�}�P�Z��ז+����	T�*L
�a鉓�_g��z_S�����e�{�r��/�5�aKU�h��b�<w��=J�&hnr>�K�-rx՛��v�8L���5h�n�%��ěñ���>�{�fr7���1�K���J�;��Rc��̗J��p��jmQ��V�\��/�UE*.�Ѽ�3:���t#a����yr����_}�}�ո �V��э��|S�Q�k�Bc��z��ѡ�\0��.Vz҇�Ⓥz��_ڱ����&<��F�Qr�=5����0B���>��rϪ+5��4����O�_T�Y����׏kl
���=�3���P�u6u�����"���bi���������D�f�4��Z��j�s���w�'����z.Vߩxmyv�̘x��J�5I��]��S����V��M]��8o�w�-�*�ό�9���� �������4�p�S'5}�Eh}{C�F.:��O���m���O�1��>�U���=�³�~�
++E=���9NrOW�p�{����-�C<=�6�ڈ�-�F������w�𳀵\E�W��3̜q��i�v�B�:��F��,��y����#�R%���Oe=�����j��EN#�����߻NVu�<}Y��wv��Zy��,��p���^lfߧ���>�����T��H.OԙN�+���_��!�U����;u���8%{mz�Oo�����϶{�B�Vx��YI.��t;r��Br������̣�!��d��xL-nF��'wGx������:V	�F�v���x�?�@o�J�=���(Wf����{@ms5Rj-1&��-�ʂ�f�r*ACx)�q��e�C{��Y�%1�+w~(�5��lo�_����
�yv��˷��+ێP߿+�+ς⎙C��꘼���[�xz�"�:U��Ey�{OC�]�Ю΢���c	���4&9�u���Za�Z�T�p����yWN4%�<�sS/=N<پ94g�W�?8>�������ʇ�tl�}�����7�������-��מ{�q��Ki^�[��M0єf���nq ����Zj���\O.�ݯr�x����Y���xzm,7�؅���TuC�6���U����;�a��Zx�6I¦�]ڃ�_W�U_�'���Vъz�"�:�;��^�Y�u�r�"��K�w�o���f𷇽^n�u@���oç�L�|]����Gi��8{����=r����C����X�;쐗��K����?_�Ν�s�{��m!��.t�r����nט�Խ�.��s��Bw���=Tv���],���A�JT�& '����@�F��޷0����I]̼{3��n�Z+�¨�$LF%t��4�"a��Q�mި>	x=��O�V:�������F��+��ً�$a"������0��
�e��'i]\fؓI�Uv���5�7Tg��Y��W�����󙖷>�����ʚN��R�c��)dm������l�J��Ι3
1���F��X�8V��yFʩ&�y�wiשl ޒ�����+ޝF۹bu���'F�5�hd�{���ڙo��`�|*���%*<���H�WN����������%;Y�����b�{G��C�dZ�|�_���lP��9���s=K��R�e>����S�����\�n�ʾ��s���ۧ�r�Wu,�������3���T�axVf����DMþZX��/
>����>s',56�Z����j��^]l��W�5�SҬd4�ᾞ�>��͊s�o�e��=]�/}�⫺�jd���[Ck>�~Oq��Wς�a��|m�=�۵{�L�*:�G���L�M�a=�����<���F�ʧ��A���Ν�ew����Κ;Rɽc7�a��H_�]MN�}����RC�
�J��ڟ7�g�c��f���4��ᄏ2�)m�CTy4#!�+QQ<����TL���ܖ4t�,.Ǔ�[��N�����Z�"�3|߰c���^�*S�cFt7�4Ʃ�n�p�ĬN��J�k�.��Ō�F���Q�RȺ���ش;��;{cj������}���kҒ���؟��������5���5���/�cd��뫍��{=)�q)Ê�&�*4�.O�d:f���р4�����g��G�_)[�B���$�8�z�/a�L��{j��%��ɪ�k��k4�ӡO�*Y�w9��/ۋ@��[�7�:\Ɗ6�އ�|[��J��0П����)h�A/IRįc��i�ϩN���}W	�TˍەR�͋53��mB&u��j��J�����J^��޾�x�CC�z�\2C �^��gQTvo����ޗ��hN��1�<	+�q��jjf�3��ӛS}�v(ֳɎ?T�w�Et�z}=س�������26q����5�v*����������e6q킶hV
��9y�\� O��J�o':���\�t�J��U��%�>��-l[{�ּ����Bp�g��z�a;1�*{��v�j�/�ï���?k����gޑ/�	�N~�ﾏ��'r�u�zc��?�=�Kz0��ڡ�}�]����]����5���G
��߄���h>}��_��!z����ܶӱW�3��K���{�]K)�=x���4��*x�>>M{�7�gr��V=��j���'x/<ӆVt[dr���{���+��w���s�Q��8u�2-R������ž��qןIQ��l�& �Q�'[��Hy��ka�+}O<5�x8�F/�|F���_��qP��d+�y�v+V��k����Wb}[&��Q���p�j��1�}��^Vu��ɞZ��]֚4j��s�]-�P�y��枿Z���<���Km̔���;wq�Q5Q�D{bcK������˭����Z�zJ۲WI�s@�8.2SV��]u ���h�č� }7㱫uas����S��;��˸T5/�[o,�ř.Dr�#���< �HT��//�{[bx2�!��9Ԯ���݋� �Z-��+]�.�����C2ږ��.�tl���}j,�v��*��\>�K�btoh֣÷�X�,�/]s�8aޝX{(Q��ڔu���t�9�F��E)��{����jf`|�����8�Ry��M�&R���e]��~��g���p>�+M��c#���zxd�o�+lt]&�{n���t�ʖ2o攙C�~o����(k}���;��Zh�q���>l��88Ř��^(Fe�Cw7�JwMv�!��2���s^Q�2:PoU2�!P�"�:�5��IEv%N<��h���f�C(���h��suf�8urf�*P��V.U�Xq���y�O:�tHrM����Ml���
�Q�
�W�r�]zֆ��!
ʖ9)X���X.S}�v��aRR�W,ÐN����v��;K,\��Ea᧽	k��./G�:�ʚ[S���Z��\��X�#�Ev'Ӫ6:�����t�,�4_\� ���KP��ƫ�m�iV�G]��6�b�|2��xN�q��	�P-�g�Nג#�>7;�.ѡ[e�벦借#c�xs�a�ŝ��w5A� �'C��n>uG]��J�����޽8�C��i �Io�Ze��DÉ]�i�0�Qﴬ���4�nei<�U�<u�����U����bL�+��?3,Ө)�ٜ�,���oz�J�~X�O�J�SH����o�\��.��E�e��y1}���2�ׁYx� 肶6�X����&T2`��m��8M Ec��8.��vX���5����������R(wpQ칢a}�"��tv���.�QF=�բ��wH"���Uv��M��:�/#�����3��=�A�V8k����:��Y��3�L5Y{��h��i'lǓ���)��I4�OOb���!�so��
��vJ����y�<��5D*��u��Ьޛ�U�����ӳ~�vw�}W�A��̮t�z���kT�v����k�a�$ooȔ��Zn�3�`ᰱ�V6�t�g<�Z/�~{���|�(��vDQW(�������QQ)CN��E�ir��gS���E���-B�D�&q42͚�dH"�C,�Z�SU.�U\m"��"�ID�ȭNQE�@��ťQ��
#3�gCB�4��Ʃt%:�UY	Qr�J�Y!�D�Y*��dar��Q\+��sHU�˰�Rqd.I,�B�E3ZUAu0N��M"�0����$V�L��*�Vt�F%QW$�����.L�$:B�b[T�.Ps��BJ�*��0)�T]����>�q���s�ߏGݞ��e��D�*��6?*�`�:�E�]Nٵ;�vI�rS|e˹Jb�o)���{�c��W�UU�F4��?V_�zN�a�Aҷ��r���#�FQ��{�Xp�֘[Z��P�S���������*/,���nkڜ�笺�
§�c�=����8���v�2�c�����}�[o�������d�^�|䝐>B׵�C&|�+MU��=+}e��4�U�u�A�����:noi��X���>���z�jc��kZ ��t�=��&-:Y��3qN��g��ԓ_lr����i�=�������T�Wr+7�.[���:t�TߎS�=�f�Q�կ=�vRh�\#o���R�M��d��������,���]
ōxrC9Wq���P?j����ۊ�Α��I�'sW6�e�e8�PA�3�c(�k���B1W��1��'��v���t]�4��yi�36�~�R��Ä2�b�����7
�˵nH6�J��ڰ:��M5J�u�=(C1_e��B��s�}�}�]��8Qu��{a"mu��ϐ���k?Jq�kި4���M��q��ș���Vx�+���?k:V�j��\�'�8+�r��*6Z�����P�{S.�o"T7��k���܈�OV�{`�'�4�h8W�Tcɓ���c�����\�,�ud��VB������z���ӊ�WѬ6Ž��~^0U�P��K���:n{��^�wO��.��)�|g/wUR�����a�E�CROo�:m�8�r�m�V<Q�b�]�|�eS�йv�a-��XN�n�/ն1��z�y�/lԩ���Y�XS{4h���+�^��C�gG8o���>�&e_�)����;��._4��ջS%Du�B�������à���Z�ĥ�<�؛������u��F��59hmIF\�ab�o��ϥd��#��xn ��n�;&��Y*@+���sw����Ǡ�w�sC��������H�����#�^��7�Юq��[���u��L�t+]����W���T$�=��ŖG�צ|'��=�t��]�(�z��sm�=�g�����A���C�?N��ewXDVU�^w{���)�Ģz�����{p����Q�{�d���.^�q��L�0��O+˞X]o0/	N�R��=��U2+B6�S�{p��Pal=c^{*&
�&r �ctfʗ��F�}�;��kW�~N�R�S�Z��}6�׳_/o�y��(Z��y7s��=Qhn�
�t����l��PLC�z�{ii�e����߯\E�$ֳ���C0�g�-C���̖�)^fk�ѿ[Q�{#u8�9R����|[�x�e�4'������rkZ����ת�/ �F�>��
#H���Ծ�O��3���+vzר%2V�싩
���j�4]λeC2��W������z#����Z�X�{]6�_E�n��ri��nk{�����d�t�7�<�ms}�����>5o0^��g�љ-P��`l3�m^ŵ�<����nI��V� �^���1g����(�|�>p��1��=���SA��������g�93N9�X���˯��M��*j�r\P��|5G����ul�G�5��ؑP`K���&h�4=7aEL3�Ur�Dap)�p��9-5���*ER�w��g��t��'��3C���슉�������߻����<�����L�Y�N��+C5�Z���(�D�;��˕\��7��t?��p��!ۧ�N|������7�Z޺�f�C^��(�i�����Z!+��p^�=�~��ɋ�\yR�bR�����Wӱ�'��f.�$^^�vԽ��>���SHvP�de��F���>���;%-K��x�y�@r�-�Z�כx�VE�V��%v�Iʘf�d��b���E���^��m&EC��8*Qõ�;"�4���*��z���D�b�;�1����7G`Y` ���}UU����{�*��۷�-tYc?7�S�I���j{+�m?l���Ӊ�I��]��9�x�1�p���^S��^>[	n~S�Wi�hߘ�W[��TZ��*k�7U�q��y&aP�^��Mk��o��'�M���5t�v�zL�˒������؟#k�e���n�9�H�4�z=�4�iT��lƥ�4ҕ�QS��:��̬�^y3�,Q�v�⼜��\f�K5�iB��ܯjNK�
�8���Ӱ���\FL^���;a8g�Z�놦����;�����H�VlCә��[ Pi��ܼ��Z4'��܆/�Vu�g�B
��tz��.�>"�>ը���.�(�Zܵ�Yà@�T�1�޹���|���V�:j�Y`���(RVcI��:�#�y�B��:Z=���A<�z'&�+ꯪ���-}�=Z�wqFS����r�]���i�s�*cC�ŤĹ����ʽN�3��)W�R���j�eV��=�ç���{7�+ZG/LM�VF�H�N����5�z�=�(Vwe"�S�w(�	ד��{ݙ~�����s
Ę½8$�z��:W�*��Q>C����_�$�n|vK����}.%��S���J���b*�Ш�-�)A���5W�Z�îP��р�^���ڙw_Nҫ��6���ʨ[�3�[�9��f�KE���:�0�L������^>2o-�+O!���X���]N]Fc��N\i�袰x�9>w>���B�K"�x���#�G�|)ug�V?N��Ak�R~ڷ(���B~�mTޘ��J9�RH[��'��(Tlyɸ�U��њ�o(x�ԩM�mؑ��Dd���WYr�R��XO;�ǖf�t�e^������g�e�;�W;D�ݶ�����
���|b�g6�4I�n�������$�yY��`QWp�K:�B1���F��~���rܑa�ۍz�����c�;�x����^�qxQ����ML��5��ɾo������#g�f�
����V�C�7��-m��,/�r�m����s(]u
�5N��>�S<���/~�g������8M��SxQ�%wQ�c�u2��|�\�5{ެ"��.��ъ3qx�����gN��V����������{�,�ô��}��{��:���ʿ�����~>k+�߻��>YO��Hv�,_}o�M��|0��5{	�p�r���[N����=���Q%V�r����6��o��񝯇��TKq+[��bq^�f�Ry񟚩	�"-j:2L�,Ș6WV�_n�\��<K��CЭݜ5�M�Z��`�ط���	�C��Hu�S�=�q�f�K6�]���v�-e�vs�DY�^Ա�O��̥"��k��b�i06�d�(�9�8<wȍZ���JĘ�h�����KT��k:
��ڽ;޷��ds~�
��a�.(�דLDx�^�Xe���(�[���:��n��~����8�ϫ>�St��3�.0��7��ɻ�R�ݡU��J�O�B�/?M`yRO/d��ыC����곻`��
�
���)�=���e��1��.L��)���q;'�ݚ�sQ�c�w6B���+]�t������7��ߣ�r>��3���`�q��W��נU�^ELQ~��_�����GL�����ϯ�-j��{:��شp��={BF>#�輯WguV�e2������M�!F��7�䂍��ʌ�링y�����i��i�
����x�[N��ו���gX��;�вf�}X� ���z�l�i\h�|vȢz!�͞��"�Ͼ���� =໼�c���n��|��nn���E`�C���]�k#�g��W�E=�ҫ��eM�6�5�[C���S�>���MM]���P�g0QyȬ05�����~����e�Y�g�>âNo��������u���d�룑��e�6�݅%^	��[����lˎ�%��R��8;�����o��"�u}2hHx�,vm�^c��w���å��s�s"�	�7y��>?��]�~���7�1�&��ŵ��f�,>g,j�x����h;L��2ZC�w�U�� q�g���-�7��߼��?W�����Π�w+v���^�
�B8\����E�Ǉ�5�i梶�����oD�8Ǫܒ}��L���є)���nr�,��{Q�Q֦TӸiN��pf�J����.����u[�q�9�SV��	K�Y :�R%re�
�.аvn���,�N�k3)��K[5>���������-�{�l0�~Y����9p�8ǻ�]���K�������~�[L9���"k��s~~��N����:��}<�����|k!z�?lT&�N�s�)l�����/%�/Ӧz�<���o����B+[kzzQ�n��1(�ܔ<�m�������l7R:씆yA�*E�6��v_��o���}���ߡ�h�y+BԾ�Ա�z�0C�+�s�2��w�n���IX}��Nc��1����~���ܥm1��+��d�2��gcP������)�Í2���η�~�q�~b��ݷ<+닳�K��k�ǎud��
�����=�����h=`�쯴�}����ի�i�l����Χ���ջKy�A�-];���g�9["|ƽ	t�F}��p����\�V-V5��SI ����o2��Vq�K�0Y�^*\�hg0�!��`�x{l������+��I��Lg�����:]�R
�TS7̌}�Y�}���p�
���q�Er�5����C��ST����o�¸ǯ0�)k�a�*�2������p*�����A8����rQs�"�7&��F����1w0�g_nt{�ڱ����㱕��M�:/�*�c�J��ʳOKT)��w Zh��x�$�U�n�;��"���1ڳ+6N睺� \��2w ��^0���[O\�U��>�	q�z�+�A�`h
���]k�����w�ю=�t��y0 �Aýw�%�vl��Mk�1!��HUܼt��kQ���M8�yn;U���ù�k�`Q�'C�l`��
���ɷ��ƚ�i�����Lg��g,]`	ni��H��s��J1�,��m\��J�b�mw7H\;9��:N�9�ۥ$d,罐4 &=�>���;-�2���:�^l�DEnѷ��Ջ�f�4I��{o*R�蠑l�1)\]t/�2O�7Y6�u��<��T;-����4�>���/��Q_aJR�ӇH��s��p��+�(��h��A57:�;���6���8�+�f.�wJ����H�"A}t�AW�Ц�_=d����=
�6�w"<%,���[�����tM�� ��G0^v'�	ɣ7.��;ZYV]_'&SZ�֎�˥��)U�Z�X��"�/]mBZqVi�6,��w�TS�W.�u�����jޮ	٥]m���Vy��8+耵]|�����t_Vʻ�B�B�o��!. �"�jK�R;�c�"��φ2�E�;ה�>aU8S�%-�����x+5���&f�|�Yk1ɛ]77��Fu�.;���<sj���H��+�B�޴W*��Ae9VNs���@�ѯ	I!���u�%��;�u�-�Su�9�����޴o��4�[�zP��%rR1ژ�7y8V�)-$�uvt4���u�O.|s�%�Ie��ʕqq�:~WK�C�';�h�`�W'p���:��%�&�1y�À�����ә��"P�*FՍWo�^	����.�oc��8+�%12����ElԺu"��T�yC��,���e��c7t�i��މ��7n�*u�{MS�̷w��f_K���aì�j�Ew��[��R� P4~�    E�!\,�-�է9p"L*�F�AA��ZRA*(R�b��N�I�jD�"�B(�B��BW-YD����Q"�f(�Q,����U#���AjU�U 䳪�R�9��"dp�i�+�j�	!k*��*��B�N\P�#�-�r�JZ�@]ZQUFer�$*�U�EUEkFTvUr�ͅQ�Y\�H�"I]��*	1�+B#����#�p�m3�q&] �H�����Dr-hI4���˗T���Pr���*�(���B�d�
ّY���p��**��ȓ+����QYS���C��\�>#���Wv_e e̇�1"}�j֍˸��%�jh�a)z�:-�k�ɔY����U��-h�Y�=J��^�0���-�{Q2�iUߪ�e�k[y���eSK���/�W!�L2�'6��d��<x�e ��Ma�J֬�/u����;Q�?6���(:{=�t9��ᮍ�g}�
;�}G˨{cYf5y�*,��¶�����B����J;5m^���"�V9��M����wݾ�z�#��j|���B�/����n��^*�����C���]��N:�l=.�x��c~�Wp��^�BYw�J�5�J�Z���э�|��q{�Lu3Y��{ǆ�\k�@>zsؾ{6�n�{���)�(�pחlo�[L/+Kwշ�.�5Q*����4��c���ǳ��^t^u��N�U����}��~4���7Ĺ�B�ji�
6|�=��v���[�6���-g�Bvu�&Wnq�@=yC�q:�N�ˮ�
�ښ����>F)�]==�^�u;S�ykV@��8�x_~�������w�1΢2u��8&c����5?'��r�{6Ww����u��C�_����讻�Զ�p�n���g�E�Ō���m�h��6b�A����y�ʂ�y:�PW��<��"���Ϣ�x�����~m�cX�^e��o#\�^E�{�u��_�C��o���-ƺ�l���^��7Pgr�1�)�����I������؛�fF#d<L8i)->ջ~�v�x4ڌ�uk��N�Z�`#x֦1E��_zT��m{cZ��[I*������M�ߪay�Di��>�Փ��Q/cX'���W����R�wK%#�+_jUD.
R����
�z �󆐸N��N�ݡkn²���_.S)y�^ߛk�Ց�{�������O���[��*����yG����eG]���'=[ �W[���utR�oc�ͽb�={HV�.�k.�Y�n^P�F�pyp3�|��<�Κ��J:�W��W٥�Rv�\z���<�Ty��8�Y��ꋏi�-!�a��fd�|:o ���{Fy�I��6>ߙ��V����,�^N�:��[��Q��y�rxR�AT�Ð�g_P�<�g9�y|�o����R�=�v�עF��̖�~�^�yoT�N���c}�����d�k}��H�0�����Խ��]�'l½uz�QF!N�b7�s��f�s���~��<��8�>�[=W8*��IPQp���cqޛ��nCu��K{<�lוT��坨ʥG����{"�U�e�^��r�+}S7�*�Y�x�ޛ۩�S0�k�j�S�s�3Ѭ����n�M���d��}�����˕}�yS�]Ot�#��W>����9K�ϊ) m��<v��+��v��S�r�i����(�x�Kip�n��%jz/��a���u��*�$c��|.���R5�J������£1`�����#��7�y*/��n���.s�*��5Ro�O�{W�\)�ɽ帧]S��c*)S.QL��2ZC�w�̕����_O>�@��h��<�gG��\��V���6]k�h��M�g��|����y'+��T�ӎ�A����t}ᛛ����T�<�Fv�~=SVx�''��\՗��hl��;ʞ�2�w�~����>4�m/h~s��+a�p N�����9l[g|�M#���Lՙ������pH����Q�3��V�Wd���&ѡ��u��N���NrE՗�{u�F��K����{L)T���>����:�;�#ݾz`	�k_�Y�hב���Ki��h�Y��2(����,p�o:�������#��ܐ�����v��Q�Rd��h��Y��t�1mĊ����(�|����d�Ov*tB��ָ2p�5�^J�F���Iu�R]�c��U}������~�����~�|g���.a���z
_��O>�~h���v=�
q�Q�p<�r����R���#(z>��/o���z?O0�f�ឺ���m�Z' x�}��ߧ<ڍC\c��I������i����m���ǜ�V;G��)���ce(Q�	A1���N��jiU�����Ŷ&��=���e�?ju^y2Sj�E�x�k��x�u�3'����ҍa�Ľ���O�0�4�O+�诶����w~��|VU9X�=8�2^\	�C�w9��>�al�NMZ<�W+��3���1�>��U�����v{̛��=��/
>��Q�ZI-љ]�J����ȃ0�Ӗ�����8�� /΀��w���u�4Z����7x^�481�f�F״s�b���d�w5���v�����F�<�O+�XEHz��\��{cA4k&�j��N=�������p�U���Ls�̍��i��)����9�����	� �,o��>�5�]��"�5�ْ��u�X1�Y����f��V5=���b�0N���S{s��m#��˼ma���=�g
֨z1EN&�!������>��[�����Y^�Vs�/+tRUC7�i<*;0�x��ϯ���摢ʝUCU��g3hp�վ8�B�ܢ�hO���<���_�Dƨ�m���-c^z2�~<�e��K�0pm�?+�GY1��=b�UyTJ�n�1�1��aY��{������x�Ly]�Y�q��MÍ��߁a�~������J�1�����w1v$�k,�!�L3
Z��ɝ �DB�{�$�\�Ֆ��.��ҡ��7������^7"������Wb���F]�gBP��"-Z=�yC0ʼ�Ԝ��9+�H'�J�6:9d�V��6e�V�9��R�]V���Ԭ�5��_{��N�̶_���@/�߫�ݜ�/�auC|GϽz��{ƛޠU�p�:K��G�{���)����{r;�V�ƥ�5z��A~�۟Z�~��U��Eɇ�����T6��w��z 1t��ג"$��y�a1���\��BYAoǩL�A7�}�SĖ�9�Ͳ�Gυ<�)�'N��+���i�r��x���+�[��ү��
�cM����Tn�g���ݺ��맠��l�g�%mP����y�S�v�,�٥���r���7�ήg�~(OZ3�@�'!�;7{z��CJ��z4�ۏ�{Pi���Xb�lϢNn+��V�j�S��3<�[Ӡ��Slڈ�t3��3O�����`�%���G��s��9^�G��j��t�삝b��������z8s6E��]��u(d%s]�(n#V���s�ޑ����O��$��#xLZ��Q�AA�(�V���kt�k�*��i3
�i���
J�
P���W��V�d�����+D�(�:J�m�,��Q*<[�y����L�e���f�Q���Y�ʲ�!��5썿�ƹ��8q���l��-EbԷv��N�}[]���s���}7�yp���%��������g����A�����~��?���SMT��ֶ���ߍ�u��j�.4��r���E2~^s)���U�W�Kۂ���-�٧�|�Y7����ӽ��A�(o��p[�Ιa�O[�.��Ƒ�2��S�v�j6��dۋ�$�x���E�ܼ�.���ч��E~Μ��U�ueN	fb��3ψ�t����x��C<�\>ŕ��yWP���k��{n�X̟�����P��j��ڊ��;�T��6
QY���)����frir���sB���z2���4��y��J��b�}ϞUf,W�����֥�h�Q�ҔbQ{�fV�6�7?�W�U^h������~Ro�'�5l[g|�h@:s9ޜEM2�����|�H��g���<Ga>���d��� ���U��
�x�.q5�}M��I���Nr�l7R:씻Lr�~!^���z��8m{�u{���sK�	G�^J]"T����c��}"����#���Y�R1<C�a���ϲ��!��:��e5f��}�������k1�~��׉�~�y��}m�FT)i�ϡ*�:�q�A�w@؛)���5��֦�=��]}.����?(%t��4=2t��o�}7��=RjYRU3���5�-��L��RUF�>�:��"7W�ם8J���"ր�3���U��'�6�A�@<�(��,���=-��J�$�'�ܾ��Jr��\��y�^���hFmY��\�m�w*t7�և�R6�D�grVp�6l�[r�2��=.��.Ŗ�Wv���B���u���3�����ﾠ����Ȼ�����4Mbcٱ�u�c����&�r�p3GoT7�{�P혀����(�Ք�?o��X�dӡ��S�t���e��)ݡU-��8~��������pԕ��Oz�Z�o5]Uy]���׮fl�B�>�}�&<�ز�w;�ry�����)���w�W�}��՘p�p\oӦk�=�租t��n7�^���P�P^x�M�X�ޭ�Y�p���͝����k��������U_��Ǡd�����fS��T׽����C}8w�4���ҷ�H��o"�&��k>5��@϶�eӽ�����*��juT5�u9=KG -j�U�������PB=�IW/�@���1�>Y�(��0�Q��v�A[�ج�["¬y0��)O�&�J�C�K[�fM�)��|&>6A�'�Y�MJ�6�F��x4�����f� �k0 h���̀$X�.k���]`�U��vu`)�M@&�ǂ�J��)�4n��]�n��3F�.�Z������8:���]u�*��� ��[�H�i��m)�X�����wb�z��.�^�Ll�����@S�;�����O�/:�GR�2�:�F�۟.�s����j/������}%�E�D����t��:���k�5dn�b��b����f�\�<�#1�-���!0�3w�joÐ[��.����SҼ
�W�~�}�c�ҵ��b)>�+����Îv�����P�J��1�D��Q�����AG�+d�����%o빚78��-� ��-Z��@��@3S�n�R���[��`hWNS�;�U���#Ar鵯t� �Z.�oWm[K)U��i[u&�Ɲ��:�%HI`�۳N�<t9��J�+o*��Spf��"���*[	oR�(�y,*��ۢ��v��U.u�Nv�g�*����}"�x�����i�z�n�e�]0��b����stT�A�����VC6�b6�'�����Ɉ{P���rڤv�=��2�!�2�v�O��^��Js�'6�����$ڶ��u.;�Ga6v�01�q�*<k~�����
�6���G'Yo��.�@�t��s���XeKԂ\��sbg�4��&�U������a"ޜ��a�|��ol�Wq�=M���=��1���	s*���=�gU�ݝdWM�'�w�Q.V�J� t��)1,w��U|Os�[4k�v5����-fa��p�APS�Tw�`��]�h읦�i��]�ـ�5�OU�8�����Q��Ǔ�n��wKM�}z!�>����C]������&����xMO���%�z�CF��D��Ư]%W�1��4s.�̤7�D��f�b�>c�
:���l����2�u][�Ĕk)���*@J]h�[��*� uCE�-n�,����z5����B�Vto!}��U�I�` [�i���U�e�ūS�wv��@�w��ޕՅD�Z���G9n�����u����]B� ��Q�P�K&�T�ZHA25*���ad�ڢejQ�$r$�$UujeDU)�sP��Vl���]YU�������X�EU���gBe\��l��J���;"*�r*��
��U��¨���r����I9��\��C9We�uB"�R�ʬ�(ҥ��ar9J��]-"�E�%�-�r�*.�Ef�UM*��Ôr�l3��Ep��9r��*V�#D#f�\�dQQ��bI�Յ J'*����p�È@Y�AQȊ#�$���p١	�\���qP�3 ��$+$�)��@���A ���oa\��7��/v.̾�}�{��a��ZY�wN8+^5��_V	�U��-���gW��oo�>���wq�������V����=�ۊQm�j�y��Hў�b1��J<������d�}+:����eL���i~��%���=�?U	�Vb/h�h&�Xm@q������f���xVf��̜pܚ�~�Q�d3�a��W�i(�y���Z�[��80ۙ�����͛2�O�}��˔g��y�>�bW���z����s���$��J��~�]7A����՞Ӵ�q���*5�.W�-�T�Y����sZl��ţ=���ɾ�K��N���8d� �Л����_�i�-�m��߃� ��T];��)�8��OLc���K<�5�`����1����"��E7����D�Y�6X��M�HįwB��3�XWp*on�xM6xO!�o,��7�N��j�n�D^z��15�ӷ�
�/uiډHF�xWI��Y�t^`�+\i��ة��{�����kBn�%�F��m�D�w�C�x�n��+g۞;�~��^����)	�V��1���^z��|�ɚC}�NNήy���_|$o$�uVIúFy�o��g5S�� ���=�Vp]�
|���,Ȇ>��}{�'d�[��{VnDn�ye7	=�<���
����a��
�PZ��H�J�:��
7��ݾ>�^Ҭ~�^�QTOb��lm��}�k��b[�c�5߾��z�J�_���8��x��w�t�?b5���>ힼ;�z��ՙ�|v���߶p��c���}����=�Ը]�λ�����J����L�?g��1�5oת.nD�S�:�8�L6�d���KCM���O^ޥ��m@�h�B���.1��5�u�=��y�U����d蠺*�5���L�_v�¢�ࡣxv��[w�y��o�F����*'9���Vs�bZ;S<�����4F����q6JvF�m"Q�7��1^��zsR�]�U	���i~t�SP�3ZgR�ߧ�g�M��>�N�l箧�n-�����N��6&-�7�/<l-�̡N*�Zup��Wo�<B��'��t����}�w=G�eDv����ߗڄ\�b��lzVFB�2��Q��iG���5�={Q�Y���oo�o��ӻ=@>v���:���,����?0l]�2�K�@U��kts�s*��zN"T�]x��}��*����}��K+���P�����x�w��Mu�Vp����z&.>��Ὕ]Z90���g#
�W�;<;�hڪ6���7����^�;�ɲ�({���W����wW�Rʜ�j�FŤ3�;f]5�=�m��Lg�YUS�t�+N*H��z,]�8�� �J��uf�yy� Z]�F��Dg+3��j�zEu]�·���8�.]Jct�ڹ,�ˌ��,��FH3��՜�����1G9������OSf����ZƼ�TIU'�ب�Y�[�J��=_C�0k-(e� l=ɝ���wYoCH[�֤zGS2ʘ2��"~���]}2�8���=��͜�E�׷�����Y��m	��&Kt��a��� ��^���|]6_�2f]y��sf׮��y1�=-�zmE}�6���l���Z�j�@k0b��o��η�U.���'Q�s��ug`��"z��s&��-�7?-��*�C`��V�1F#��d�^���Q+X1���U�Y�AmP[F�k��Rv��x�T7�ǹ�ߊ~t��y-�k`ze�nkU&�����E8��a��$|��me#9m���8���~T�B�\�:J�X�e��y�ʆ-(S�i�S��˪��8W�g�h�4�&�,.����B�Xm�	�h�RΜ�λ�8�ŏ���L��s��g_t�}��Q��2�l��r3��=]�Q�/�mo8.Ow�M[6v﹯6q�;��~�����
�Om_J�5�H�8V���0D|�\W��D���`+�j�O�z�;�ԩ\d��K'<�� ��
Wń���9��ö=����S�xmz��cK��*��э���N�rr<������i�����:�Һz�y;cK��ݓ�Nf��(S�Y�^A��)9���IQ����^Y[�	�ڂ��?{����N��Bv�u-۸�e��w�/5;�\m�n�z�Y)�l�R�����H��Sk6�g��gQ��V���xS�m7s-����g�.�ɉ�'j*n�bӵ�7������t�����vy��<�����$D�.5��	2[$����k���@WDqFWm�զ���v���C�7�W��T�e-r���.�zwPTʼ��|n��Ւ��f��H��#��6+ܝC{��u�(n���$-uY�,��[�!>�r�Y��F��/=[b��ˍ�@z���zTӟm(i?�o/k[�y��E�w����틚�M3��ҫ�J�2�?���'�H�dpǽP~MS�����њ5�y��,�>�X���h�C�^{�� mz��d�*��sĠ�z�!�B��V�q�U����z�������Ln���|Z��VZf�K����[��|t���ZT��vl!�|<&2�)�z��}���U���kY��߽N~v�a��ɼF�B�kz�`۟u:��!������Eu���y/��������]�j}U���1��H�
Vp*%�3��JW]q����~(z�<z�W��}�[��C��=ub�^�\���8��R*��J��7n�,4�O��7݅,���C���a u��J�>��'���¹���қ��XG�&tU$����Ѹ�99�����5�$�!��m�[󅅇-���܃�%���n�L���h�V";dar�@8�[�R�:�QJ�mt-�HZX5D]r��Wc�G@���;�ue��%C,�th�]j����G$ծ t>�4���Cǧ���u�5�B�=�؟п��u�3l����]�U�[{}���7@O��~�Z��6Y(\T�s89F�/�]��m��@��3z����u
�3�*!t������zh?�9�����UV;7\��/{�{�9;��1�l��NㅥR��g�F���2H\̹�M̟w��WyF��	�}��Ctj���4��I��{+��\�Tq��k�F���b�I�o:��6V��*C�Sگn;�H�c g\z���@{��k�g��ػ.�A�w�u_�O�!�X�vH�����o�����V~2�����K�t@r+Ѐ���C}z�=rz4�l�M�	���!�U��/+�=X���a>f/	�Ȇ|V�]T�}�c^�<�;=�B���H���O���0��jf�F���@U�s���P���wy�z�&�/��{�g���~��lR�7����ڂ�����T"�����N���`��CHj2�K��c�Y���<G^m�WL>i)F�-�J�NVV��gk�bo��Ȱ�	��ژ/h��j�fuj�%��n�s����n�w�'�E��$ӣ�eyק
5���,��x�D���Cg�O�:�p�=��If*��\�y�{�68��6� �u9��z��ԁ�-sy-ʸ�a
�|+c/:�Bu�\(�i��q�<�f�������zfE���ҺNL-ۨ@������P�Թ�P�09�����~w�#���NW�H��ui7��Ʌ�Tu.���x{׫���І�ˮ2��dt� 7>u�#m��	�S:�??f�N�oR>~n�t{�=U�L�2)2�3�"t��_�w=t�f�Rj_��F���8����o�����_����!q��;�m�� Z��5�C�ߵol9��S˞ObB�lH~�"0��fb�è��!q�$w\� ��R3:l�;��*����j��DOV��2��j�TX�D�MC���$7&kq�w���Y�Ж�`���R+_S&:�*ʇ�M�)}3^,����#w6' ���X���9=���Oq��L�ȇ�#@~1Z��x�xߥ��M�\NA��`��"1&'��/+�60�O��߃����^݇����X��":S9aK�r��e��j'L]�k� ɵ�8�e��r	C����1���f��=��Q��iH��Ǻn��Tj�E�~�*��'ӑr����J��}�\s������#�|���#�#n�e'^���T5��^S�=�YY�����s��}>��SC��Sy<�ޒ����0\���1t�xG�7�T��Ի�3�nƽ���� ���,\a:����nj7]`�JH��g�'s�+��\�t��=b�g:D-�L���q�dӪv#	At��f���X���{����oqcnpnI��D$n'���F�_��Ճ��0Q���2��G��s�~�y[|�B%��ȍ���T�R�ħ;��C��
�)��tr�9�b��9u�U�����7)�]2��|`�LN��;>�q[J��O+��{��\Ŏ�<.�K_3�ģ�L[��5� ��8�I`ؖ��`9���s9j��:Ǜ�:��*7���� 1쒤��2���c�k��sҽ�޳�h��v�
�Ŝ����}vV�wʻ��ע�OC��R�]��8�߶�XK��C�{�{y�4�v�J�X�|��yqe$� ٭nn�̚�٨�ӡ����eq::\����A�ŚF}|&�3�����5L���s�ˇ�!��*ο�p
��FB�>���*ՊA�3���3�K����b����rz8� ֒��9��ɡc��wfG�����9���f���Z�	ڬ�W��T�r J��O1��4A�x 'Q��zΆ:I��Ν�}�O�u�04��% ::o��,WI�30�e8X�iк;�(V��\��Mnq�c�7=��:8*w�Og
_N��c�r�M`���HΔ%z��㘜���j�����F�teϪ{�� y�mG{K 'G�Q��헑4<���?i�{�1�]����tu�c+�+���5�Qb�s�ь��������MS̈́�n���y����r3'��c��f�Tpl��F�Wp�K�'����(-�C:�7�W�e:�����s��A
������@SRa/�J���Zf�H}(�:��9���Ǜk݃�z7��}��p[�ɯ�t�S�ʀW7��E)Y<�_w��W��0lz+�1Ku,.�~k��qJ���,��Ӡ�ʇtPבM�#�J�١bMJ��e��h������sy��ۓ.��f/*fJ<��ty;�H�ح��&^v�"S%]���pi��~�aTZ�zwnܠnu&ť�
�ֆ�f�����*�Ϟo�2��p
A�pv��Q�B�+(Ҕ����Su,��V�%Y[Ԁ�9�t��N� �f�*�R���Н]+���G��-hz3$en����K
���}4%ˋ��>mQ���ާ�m=�y����d+�o6k6H�4숵��zu|�b��3��V"��\�gT�ڝ�Yn;ȱ]�=�][�lpv�[Ie�neԮ\��v遅,*_ ._]�܆
Qh�#���7:�����]�����'Bl��x \�ѷ�����F�3�8�x�p�{(.���]��Q��j`�c8*{[���ŅՖ%C~��ˣ�'1�@x$wt��4���T ���������@�n��͗�u�wj��md���=��o;����)f*Ysv���x�2�b�!sz��C�S�#F��j�:�����ݳ ��5�nUi���Ï/���envε����������a���t:�mI�M��eRֳkx����� ���5}v��{v*m�Ge��}e����y�w�����ز3�p&.�se�L�'�&,o	�й�i�u�݋�]�v��uZ��ŀi�\�����ub3�]L9{�Ì�rЊ���_m�_"���#����sn�Ά�vR�
��dZ��R�yp� ��-��u�wP�������-��U�O2�\��K���*�VB�uKg2���M�V/��t(�-��6����;E�]��klt��*�e�o�MNEb[�K��D��N=�,�Zwo$݈1�閆*�,��>��P�;�W�����u�o)�h�y��]�Sef�)�m��}w#���jż�Dˤ9\�
]L#�Nߟ���,��W8p�#eL,ǒs�� v�np��(�E��][�+�7QY�2�3lTU�����Ee#��8��k�U�y���ICzG^�YL�0��Օ 1u	�ܧ�\[{O1v���x ��4]�Z.v�J&�,2O�z������VK��.��C�cԛud��f��CH�3�L�u+,��i��c����C�����8�:`��;˥6]pG�jU�A&��d�.��tuv��I[�ذ��H��wjwr�5�n<�3�(�  *���@���$"�'J$��	�g"5*�PL�	
,.Z�TQ���Ҫ�4R���.�*���DQ'XL��!$	G�d��SFQIJ�r��%(�����@G.�R�
T��"��(���
*��̋�\�
����
�PS()3�(��g���TU��Y͠�\eU�g"��UEʢ�E�B9]�r�ȹDL��jI��)("(*�(겨�a���Ă�Yf\�2)�#��"̈.*������/��(�E�,r2�uҎ�b��C�乺sI��q쓭��݂����v~+M�U���5���������@w|*��[�N����W��>'2b��up9(nŜ
�c�6�u�:_T8�rrwppt�0���Lu���xw�Q=�wV [4�p19,d��]�����秘�5�r���:{P;�u�9��骎�c�� �^P5п��e���_p��{s	������ɾcD� �wT]�@�C��@�at��TdJ����0��-�f�x^�tx8�2G|�t�H k]\f�:P�j���^�b]N#ݔ��X�!-���z�n�x���L�}�2xtt����=$?�9�O�j��]�w�+j8����$o��r�	6aoκㅢ@�g��GI�"2;zf���G��*^���}=�3�j�&��xx��HF�c":�P����a��M����k�Ӫ��U�����z�|N�T}��;��v[aߐ�V? 1��t�J^��B2�{��'}�u5�VB�4Ad����'�u�Y���e�,��Yd��0��8nW�# ��]�[�Z�^M"�g%�EÃ�kY}\*�
J��Z �4��kk�ʴ+_w#��{7��4���Xw8.�w��N+��Z�d��O�8�T;�Vvf�0��}�`��0��X�j�'�C�v�Ӽ'�|7���E��:����S�=���������d��t��	��2�^��Պ�L��8=;�헙���������!�y�
���HA9ߗ�f3��)���'� ��aъ���-�X��z�z2q�3�{�A��l`�4
��>��ʥ1���p�0]+������W_�����*��7-ʽ6�G±2��Ϫ�Th=~��7��4��d������-lX���M]��j�_��p��Vι�5����Wy=����T;�!�=2�=$b5T դ�'7�
��5C[k���=�D��t�yt�}d�7̎�/�
s��FS6+D�P����S�;�b��5ކ�w�z7�*;�6L�Ϩq�WP���w�lz�
�1�:�����Rh�X�u
����=�.6g�wH�W�<�}�f�q���^=���-p�+U�+��򝶦 �Jŉ��P�zn��	嵐�O��<�]׵�k��$�W�e]����=���7��A��ݙ;Qr�ķ�ʎ��IU^^�%�+�_-�W4$Z��2�����GoP�7zz��@������L��++�����z&�,lGz3*��M��L���==ʣ�����y����$wwMj�+��Tw�z��]VM���K f�W
�(z8�7=���֤w�P�5�3Jh&��OU��b���y|��瞻��B��|��cƳ�%m+�v� �6�\#��7�I���"��J�.�􄆽���M�������c�Y�q�Gz���_L�:�u1x�xX��m%~�B'��K1ە��ދ=s�&}ӿd�=zH~��*T�r���o�ׄz0��U��If���u]G^�*8�g���v���;���L7+Y�Q��GC����� �Ϯ�qv.����G�=�b��@;<�h4@��oip���*��s�a$֨�|��攸�b�|,w"�F��M�!"���#C,��et��%���# �i_�GnW�z6U�β��;8a�Ctvr�5���k��IL���A���{��t��j��;�'c	=��K�#�Rq�鳻+p[wrW}d3o��*�Q���4Q�v�-2���lA��{�q�����x�oɗr��I���ҽD�T^�z0mIڽ��oy<��`���?U����`���L���Nj.�����r�`��ndĉ3�o��%4��С�<x]�C�pdD��1q,��s�*��ꋒ�v�}᦮�l8yr��cw=v�u�@b�T�+$���^�fX(g=��7^u>���8���O_���l�5Q��4r���T����,R�P�3�f�A�]����},�R}d���"H���;�#vVL���NZ�}�QK����{�n2�ǹ��UM3�����0{zh�\���Wd*����G���wp2OC��T�:Ԟ S�=5�q,Ɔ}�3D����1FǕxv�y�թPz3�lVM�{�n6X������U>���<j�CV��(j�N�ܟs�z�W��nz%*�;��:2=�no�q�{Q����w\�ޕp͎�T*y��>��_����U�VJ�����\+�X�T��*F�Mdy6VE��Y��8(��!PG1f�EWa�����JY�h
��l^�Ҟn�w�,���[��b@�����������cr���u�EaY|}镔����Y9ӎ@Ծ�#���{�歃��1Q=.�z�_-���Ѣ��Wztͅ/`�ǀ���;�,TY<5ϦPK�ӵ3}s�m�{�w�ӝnM���ǯ�@S���KNR>�]��-3�o�sQ[�a^|�'�7>3��y�����ܟ@�G���� *�����W�!��� �3�k��ʹDa�,��*����ϯ]`��<Y�Z��
S=R��F)��f�z�.�}]t=d���e�Pڋ8}�����9t�����Й�![>*��UmtgC��@��z���.����ٰ����p�������Vk�����{�o��p�E�w�n+��$a�n�\�ز{�@k�~>�w�=o�/}���]�=��< ]1-t��48;��h��X{�$�F�6z=\z|�KÕO:=Q�T)qt�ǈ_ w3�2�t�PMS�ʼ;�s��o���pZ�RRTB�yW�IX�83!� �03�k蝘�;!�K�S��ȷ������=v6����5S��*�v��*�t�i���d�����o��Y�{s�ps�����U�j�_!90�=�JJ�GR&x�>�<:��_��"���.g��'�����ղ�>ʫ��c��I��]q���S=<xK�|hD�-��S^˅3=Yy^G�.g��\��jL1FMJ�<4�� �5����_ȹ��R���U�ܻw��=�6+��\l��^159׷>�U
�d��0�;��?��^]�J�=
W�_�ؐZ8)��p��<�}L��>�~�'�o��0s���9��[��ܵஈ]@e96�b�(\&pV�T�5ףD���<mz���9ژy~�v�/_�]��ﴗ�sd���U
�����q��b�u�uo��>�oF�,���W�b�L��VB�����=S�.9�2g��M��6��Q�إ>s[��%Le�l�R�Uĳ�����9��7�N�Yw [�ӹ-ʸ�V.��X����\��lŮ�m~��j�k s�E�f��I�L��C�t^��ran�u
��U������엙g�6�xmיĸʓs��ۆR�]�X��/����ݩ�G[���K�	�B;�:#Zi�u�P�w��ٹv�9�ۃ�
N7
y�������sX��I��X;/8�R���m��K��l�b��(w�Ƽ���Dw�]?Ɍ�I�;ڔ�]��z琺}��6��%W�8�n���	�P�E���/�,\x�Nw"+�#�͊���96��z��8w�2��<1�*�netȤ��xz,���TS�+�����W�n�8k���6[,_��S�P�<x�D�P�7��@k��"EfR}��B�ظ�s2L]�뎫6$��(b�3a�z��ݺgϞ�G�K�s�T�/A�O�H���C̕X!�ۥ[��N>�H�%w6�_tdZ����Uм���G�Pfn�+A����yP�:p��˪ɸ��d�/9Tl>y���6s���R��c���qŉ�������=��}���^�{V��?d�Mg����.@6{'�ƨ
s]#Ȱ�ULa���D*2(S��� �׻Nnǂ�����{Ò�������Gb�w �/�E)�Fݘ�N�)aɘ���:�P���M�	���m^Z�Z��P��H� �y�)��_'W�S��_[k��S��%�w[P���K�q�J��|�/�������ڪk�o]�7���>�8��	�t�:�Y}ڃw�fa�yG�@s���Z�'<`���H�q���/5lǣVTn�W��G���$j���X��ҋ�2+�}�@���(dΩ�%�ٵ�F�azP���
�#��v��{���2�wb�d7]6��q�4��ip��Y�"S��B�f��{N���B���҄��ȍ���K�@&}RFQ~�+�o�5����/gk͹��v:'�{�c��xW�+�zlWS�˩x$���s������
�o��{ǱOp����)k��ם���	sq���,�b�e9B��+���+ �����w�m�"�u��ŋ�t]�A�q��0��P�+�G���k����r9}@z'��`���@G���V����,]C 0}���D��^�El�>�[����}�{�f�_���Wp�i�#�R�K���T
	�3�xF��r�s�ݤ�Ls����ҡҮ�/�T;�̩6VL����OE�b���?0���y�đk�Kv�9����N�}�׎�}�������ď�n���H�^�6m�I�����Ó�.�_>[����k(�{NP�v�F�q�#ͦK��@�g��G��v�j̱��?C�fP�&T��'��2x;a�!R)�Q���U�z-�.�x�wջ�yM=���Mzx��:Ԗ }3��,��Tz\���X#6�Fc��ˊ\��U1�4�D)�q���B�p6z���/�����Wb'��Q�O݃�(zg$9 �5��c�v����ڎ�m0tx�����}'꙯.�b��w:�f"��`Js&^Ӹ����E��7���8z�z�eZ�H��x�t��oA�8:��Ⴁ3�K�Q�
^��X����%����VV��-��z�Zp3�~�o5ׂ7��
|8T{����P��KNR>����H�h��[�lH�=�0���v+%9����6ta�9Ȁ�T2�����J�Y��	e����׳�[��Ɠ
嫥Cg���ÜY���T�:��~��~���y:Ș��] �"��z�똴��+8�
���7��j_�]q�t��^=7b�LG0�*v�H�=֭�P�����g/�)\w��#P�׉��ZYz'=�67e�;�q�pp# j��J�E��
�8�`kk8�Cr�|/o_ǭ-���Y��ˮ*�r�z���:�0��f���������A�T�=�Ղ�M�����6%��1��us��oĀ�8bb�]P��sv&�Kn*�v��m���T�4�����]�@�C�P8�];荺 �P�z�7�^[��s�gDL�棲森8���	��t��d\x̹:=�5LaX���A�K�'��OX]쨒�[&�����C��D�}�̞ w��OI�,_뚯U�����E�s3([&����
�q�Q�c��8\%R��g�F���ɚ��&6goG;��{�l��Κ�_�;1�*"�����xi��F�b�{+��{� �/sݽG�vޙ��68�w	A�Q�L�ԯTMκچ��B��3�����K�t�ύ��
�oe+��9q�7��{=�M7^
̋z�12��ǫ+���}�K���D�چOL
���.9�Y]%�Z�9��!�r�C�i��}?ҳ�Tx��k���S̫��~(�u�t'h���V��j�:�*OtNޖ`�p.�w�����44��������8%)j��s�DL�%.�L���2͔�´�+P�f+�bRwvK�P�*+�f���o���4����H�-LX޳��kU�ғ� ���0*�I�4^�0�a�obJ]�ՔtRt�D�����fȔ��ų�A�вuk�ʑG��\z�����,�o���>8��@���)R;K�"��K"��ryw�^���^wfv��gh����@&BH�^�fL�K��-@�L��$�Y��^4�e*�3������j�gTHS�fS��싆�iuwa_��Z��o��G2�!o-�ô2�T~e��:��p�սʴs�#<�E�ܼU�pt�̦d�G&o:p�\+�$�kK6d�Z,X��l���5�a�"y7wv�<JGm��n��!�u���h3c���L���s��㸝`B�jwl
G�e�Ӥ�Y`-��'��ۊ��r,	�ɮ�%}��6~�w]C^Vc%�%��2��T��o  ^��p�q��j��\��^�k+z�@8��n������s�}FG�WJ����vʏp� ��M,{"�Gt.j������'F�t���[8��@�A�r%]cV�0�L&m[����r��\8{�x&��Ö����e<C�6�VG��j���].��Ɏ��A\�7]w�IVV���G{/i�]�˭���(��M���{�6^Y��U��Nʊ��
��hZY�YT(ٺU{�q`��h7������;�`����2%� S�� }y��g�;W�.�t�[O:"�ؠ:���߫F�m���+�'4B�o�b0.cݦ3F"V���-}N�d���+D:3'c�G���ev�N�F�6��=uc�Z��ԱS��+x�d7Y��-�=R�z�iZ���T�����+�S��$ɏ�R@H�Ьj|�VRIr���8�SG�+l�2�V��2�5/�����V]<9֥�� �ߥ���[|��q[�|�	Xz�[�#��_Bq��,8J͵�]�kT�.>��	x��7ɴ�P���x�*�/�3Z�K3F�M3>5*�f���ǋ졭n�����b����МR�7e��,�{;��q�!c�u0���q���27_>���b3�V��M;�Ѹ��
n��˥�GSB�
�����xr9]�W[��SV���e�'��0�#�8ZaB�,�fW5�;


.ʪ�VmR��K)T+�XYEp�q�A�¬��8Rt�L�I\�Ī�C��WwG�rs��('Gw;���(��)"'2�֕DG	2��B/P�Њ�]��r��Y&j"Y�QPG�����'8�L�$$*�UE��Z�D˔r
�E6FH�PU�Є���UJ�YP�̜��(�O2�(�TW��I��Qr������L*aF�H�"((#��{����b���OIك�uvv�M�b+N��Ai�n���+4�U�Σ5y�2�s���tWvf���®�?�u�Ѭ'�9�C��U
�z��9��ڏ\G�a����b�f�/��g�[л��VVM\�2e��M��1M�>r*�ڜ���`q#��hR~��ez:ݿN�7� �*�
�et��-ʽ6��|+��X�)���Y������~Ώv,�B�+����q�P}���+(
�ҺM�[WP������f��Ҵ��w6�
*�N��I��|d'�����UB�ui:����;���c5�T:2��c�Tj��T�
�.�)Ϗ:,�6+*F��q{���r����7�\�� }8�ï�U)��NdT&@��d�H�@jM��v�u��U��`;R�:�
s@��{�2�p�u���.x�����@�\�a�"��Sζ́9�̓|��\Бp��j#
H�������ŷ�·s���������P���H���n	��̈�X!�fT�j�+��{5�f�NKU�'�{n��t��+�PQqy����j��b�7�]�Zqq��&�=�Y��u\8b�=����hJu���"k�2���N���8@���:P�S3R�r�w5��l��Vd7����m���\�
�Y���ʙ�	��#��H/�!Q=�����7;��鞋��b�a���R�Uc���Z3jE#�zk�2��z&E{�{R4T}/�z�r�W���/*2x3q��.�.7��E�t۳ыj�E��6����
�WrV��XG�f�k��b���:$vz5��O�E��k�f53�����y^���)*��3�lN�u��÷(^�R�d<��(�u�����;s�/!��GE_���ߌ���&/;g�}ioV���چ�u��j�,�}�>��l��b�z�w����t+�2�~�Q��D�T����|�¡�A䯽��Ǻ=����b��|0WqB�Ɯ�"7��Ȥhd��{�¯�r�����gf=�z=�]>2�c}4=��C�R�$���x��kC9���'˼�.y��>9V.����U�l�c�/�.p'4e��%9C��vu�fw��B��:�s��<>�"o�5ǔF�y�mf�����_j��VMQ퓕2�^��t���L';�χ���4溳nPΆzlz�V"�G��JhכeV�h���87[ê6ӭ���Qٓ�Xsb��b���96NN��E�+=~�3Lf�X^w鮜�G8�c��s�o���V��˟k������ +�WK��[�;��g���X�d=�T���MB1&�������<��wu����J#ӱƪ5��uX�FB��(X�J�z��'m!|�����3S���t�z�]ă���v�M���eH�γ9q�P������8��3'f�2�B&zk��	�s<�1�4A���.O���ED�s	kH�rT��dڔ�Q�`���I`
�ULU�ƃh������e"�:l���v-uYc�t#�c3�вh�S�㡁�N�l����g��k3(eny��GF�
�q���K UoU�X�����q���`	�p>�[΢����Iz�����O�<ly��
��{�}2�TL.�����<@��G���J>շ�.���yǝ�}�t�X�ς�Ϊ8��=q�+�;���T�;Ю��_�z������cvI��â4	1n�Aٍ��m�;3�e��\�AZ8e�j.���ӧ�.,um�q3c��F��r"$����E�f��F\w����a�a�5�il����bZ�����X�Y�e@��MU���NJ�J�c{��JuJ�n����lbcV�@�p�5έX�{'��=�Gt�ޣ	_�Wa�g�lO����+������v�7��N��P�^[���]���Ǫ�Xg��r[���6{N�fǣ'rk��(}~����,?����݁��U���銋N�7Pڈ��L��>����؛'����S��#>���tee��;��邅a��{+����ub�el�A��8��
�Ҭ���<tO�!�vۨc�e;�|���1 ;�t���J'�cU��/�wV!6���E�ET���Ed���G�7�� ������\�EPr�����v���Dí�X�9�zp\L��F�0����g�C�溸��Q(]q~� 97����8�{�C�ч����K�z��0����Y<:�gq��=Co���l����jH����d�j����cy	5�eC?~���3��O��F�H�����p��)�(W[�>v���\$���m��:W'�W+��:�L��������"^.����\OL��$Gev�,J����ǀ��z��"E���/wv�*�r�\�=[��IT��;fwt�w?wt>���`ۨlʚ��Gf#P�Eѫ��3�N��U��9~��1���7��k�eL����Q���Ԡ~�t����7�ez�-�~ N��������l�V�ݾ�� ����Ӝ��zU�6$581��oj3������\6�x�{�-�<�C���\�xe���+���)jP�s���HwW����S�'�×���������'�c%�ҶH~�F��HJS���ꌏgMԈ=�}��Ue�{=���ed��R��-Og�l6v����*�9��ؗ�
.�U�����+�����a������貮@�+�r[�q����38��t�j
�"'���b�ܕ��}�7��zt�c
��J�90�����FMuy��v���ñ��ׇdJ6�1�w�h4rd���Ƃ��U�OH�+'�]O-�y}7��*6pKE�a�)�9,(��ַ���V�!��£G3s�����6��Uυrl�3O�mKa՛֓�o-X$[F�W�*�P�61v�ꮓ!�[��%�r����2I׼�^Hq-��.x\uh�L�f$�;Zw:H�*&�y�qѝ�1�X  �����pM"� GL뚇�|r�M̧2*9� �8�1]U=!��*S�X��Yҵf��=Uv��(�T�#\�@�G�W��!q�3�'U�X��x;����¤�}Gt��t����!WyXN�≩a�(����y�Jb�Ȑ�}=p.A��P:A��؇vc�lIQt���.�����9��2������!�� �:B��Qޜ�^�w�U����ܤg9.������� t���s�Z<'����O#b�4*F^�+��0j�#������3��7z=�NOG����2�x�H�X�Móa��]H��b�U�����y&���z�X�@]Dq�M\����#��l��k0<��P���f3�[��Q��ϫ=������ׯ�x��÷(\a>鼞R�d<���j�9�ݷ�������z�=O}�1u��VN�o��j���;���Z[�ZL.ͨnA�޼��P��GB��А�����"ۡ�R��Rݥ�p{�뭫%
L���T�ZE��V��q��(t�v��]��)�6͈2������wy1���������rY:i�I����-w�t-�| �\{>�B�ۢ�{�\z���:��j���˕Ü9+����ܨۄbb��v�+������b!#K(�"����O2U�#�Fe15��kT�������N��?/-]��}u� ��Z���F_b��^��wr�+��������O�`N*�_��a>.�q��]�&��=v�O�|��~0P�>��}n�X��t]�A�q�fo���zx��j�e�.�s;ݔ�-��ٷ_\� j'��(v���N�*5��Ǖ!�x*oЃ�q�%�o\�J�z��t���_����&5��#���R�L��iW�/�K��c��]�jWH�LwMOs�w�t�2hX�YP��6g�a�,��n�z��茞�YP�Q�	zx}=���_�ޚ �:��O��<�g�y��փ��V
����y̙���4�Gd),]=�_q,}V=�Bܰzw=WlT�Å��^��uk��LԻ,�mj��(����������ˑ*��ھW�I�����fWu�j����p��P��ib�ѽ&�64l�����}W\��W(J�e��p�|�ADg����>�J��ݥ��3bP�9Z36�Bɠnr���� ⷐ.'��E���B�tJ��;���GG����s�`�&�����a��[��~���em0��z<%35�s2oo@�@�w'z!������X/揀z�M�cl��dY�7O��s��{��t��c��['-W�xz�P�pͅ.�\ +�<ru��f�Uں���>�İ�#]X�:�z7
��ǯ�@S�j��s�t��������� :/��\��bzxa��ͪ2S��w�cD��[����>O����x�Y�Nΐ=�b�)Wr��7-θ�`�N��|���U~�ev��^X��J�H~��sc�ժZr�b�B��u9hC��66e��a��9��������/�-�pȉ}P��DĠ�u�CE�u`�����nL_xOeծZ�u�Y�_J8'�T=�PǢ�w��� /M�B�s�A��c��"�uַ�!�"��jQ�$�X�-{�Sb�����
�)n��Ӹ0���Z�G���5gݗ�WX�N�B).䝯�lщцjʘ��[�o��Az�}to�|+7L��Wg�N��U��3�0�xp�a�7��`�0�v��Hr��X])��y�~�WN�9�EQ�aN9�q3�5�/2FGqt��T k���.�g����z�ndc6:	����ï�ÂO���5/���t��1P�3ç�~���9� �̫�@7ߪ}6/�}E���*�xl`�#�&������`;�t\�V_����*�qd�=$z����3Ds�S什Qو�1Qtj��xx��x@	���y{���o+@�g�z��c��#b��6*���&�5��?Y �ȵ/�G{�}I\�]�� � g}΀Nk���I��eHǦ/ئ@�K�������E��z{��1^'�\y�5�m��4����
�ʐ��Fz)Iw��@l`�w��=_b��ɟ33���d��q����;�`�]͢`�~]	v�C�9�gF����*�)aa-Of��m1b����O��t����Ł)����0OEfӺ[\-:GHU�k��Nc��%!�Ӯ'�e~��*�^����P��F�����]�\�R��,jss-�rL4����'Y���Z򠕨J��*��D��k�eq��x����n�˘��`.�<��g�=7�7w1���5��u{��S��þe��LTƮ�B�������'I%Q^��_��O�c�8�)[��tz���
H�u�C]:�Өj=$6G�F��4<�K��"�+7���P虿2o�0��^T{���*A�2Ǩ����GO�Ι>�z*�L�O;�Kb�������yؐ?����U歾0��!�d��[o�tVt���Ғl�w�GP�%9�Q�͂+Y� �.��O]��[yC�ooz� %>2��fI�y�u�TY�!9�nP�|�L�joS����*�k����D6l����T��G#pMTvgҫ<��	 uc���=yY��7V��b�j����=_r���;�܋�e=��0�+;�>6}ו�u��5=����K<��E��zj:zd�#b��"��.^}U�z�QW᧍A�_��@��TeZ^=P9Ɠ=�l��e9���8��]fu漬X�ּ������s� c��ȬU�rY�D31vh�У)9uʓ���DA��Y0L9-Æݱ]��a��Xggv����k��ѭ��v�`֘���da����v���n����Uq�Ƶ�_pz�\ξ��Y]D��h��}M�v��{���L�f��:f�1D:�N��wVv�y����R�;���H�9�G���� ����Z.��Y�̖�S}J�m�\n�����U�2y`c���g���`�z�sz��Ywx��o�Kۦ�ܝ�e[P�ܸuoTvgw+�u���Lj��U���mf���2�T����O��y�5�`TbG3\〞�@H�*G�=��gTh�;�������e��
gq*Y,�+�˴~:Or�jr��(�:�n]&��x���.;���FcQ�X��5�}+f�ڗÜMF�,���kт�ڹʖ����~�e8��QH���b#�WR�4��;c��i<]ʌͤ)�n[ɏ��绬Z��u����л"��:��9܂�`Mm�����J�Iڎ\yzày]Z�V�g0��}��Ob���#5nԸvc�NR��qp�-���9[ܯ/�Ӂ��E��Z'Zn����E��T��2�8�ڻ���U�1��YT���J���%\O��9�v��2��Otd�$(��F��@mN�k:��:(Q�{70̍���15�Z�R�t�Ӗ��|e]C�ǥ��I���3�S,tA���ՄcܭT4J���=z�nt�Tpv\��O�S��vwo:��`)��3)��P��4S�� �� �;�+�1��z��C]�z@��D��v#�ge�9i�� �e���ꭆ��XqN�5i�e�`�M9ݙ�E��7K�5i�/)����PZ�Q�(�G��2ȷ��#�Ö�c}V� �����}9�,�������B)l�-e٫;��u��)�Qj4�zN�!��0��)�ҺT*X��j� �cF��Ai�����{iuu .�l��m-6��N%�\�P١��`Fos�Z�cn��+p��u����d��1�ӻ��Y˳ �� �+��`S.*���洈�b" ��J��L� �ʊ&TQGN	"�N�M=wb�.�ʪ
�Ԋ
�d�UI�p�(N�E;���TGP�2�ɹ�O%]�L)�*+�z.{�
r
��I��Zs�
���9�r��R��0��( =7\.eS�T"�dwsz�;�Tu*ss*&E��\�ng*�W;1
#�UWN�E����\w\�@�șL�PPFMܱ;I:W
eR��.Uˎ�G��R��
�PS�r�Q\�Uu˗��QEQQ$��9�.�.2�d\�%��a\�����ӝ2"�#�TQE��,�
#�]�P�;�UEAQܤ�4H������6���k���&v�=Ҧ�{��E3�IV^ی,{e#���-�w�5v�c�����Z5ޅ���v�nM�?���{��\	�o��LoIx���޸[��篼v_F�y'����k�a��o�f�H�\k�}2*�#U�.a���7��^R�:7ԅv��K+�t{ܡxO�o'���$?i�B����(�_t�O�Eo�us���V��*N$>'�?��xO��SxK��kv���w�mv,���6*;ǆ)�;
|#؝F{�
�̰�Td
2N���ژjV{]zӺ��C\�m�U��E�b���Q�P��(�K�@&g�Ե��>��9/gP}s.E�9.*�j�s��<�a������w������V-�񙺋��|Z��<��'�w!�ld����x�Vpc���;����Nq��q5��v��:͖-�Es�CG�iܭs�!�J���aQ3��b����u��#���k�����r�GN���:����S|`�۞�E;��<+�%�F.m�Ow�$C��X7c��A��*��t�ﶶ��*���r�
ti_tH�7Z�Y�ި��X�&���u��ܻt+��{�g*k�T��B�b�G&��D���V7+R���.��lL�2�#/z�	�a���
d���k7X]� R(�N���]�h��*�쌞�P���ٞ�yv�%��{���qu�&;������Q:��EOx?8=��C�Y�#F��̨Nx������zi���1��H;�zL�����۬��U�|�	�(guV
����e��j�1~޸����zk�%Cp
6;��N��j��&fc��:*��U�^�j_��`yS�=|`Q����p�,2l�y~��AN��;�a���|��Y߼��ڎ����<λ���u⇠��|}/��4-��5�6�ɖ]@�yE��Ξڷ�7xf��O�).s�8|��=q�r��8�s�>$k(͏K���4E�Fѿ)���[}c͹;�V'EL����PW����T�ad�1�X�� �W�|V��wfנ8�g���
�Wp*>�ɛ�!��z�%~Wb�%9����gD�:�8(���r�oP�jg�Q���jbc�V|2�{y�~�׈�dn��;�H��\]���f[��K�N�S�۝�1ɤ]M̹��7B�6���^7��
4���db[��.�q���%%W��⹠��-1ˮ���"�
�i��%C���p:�N�ά�� mOqtҪ3�n����،>�qL+1]m�*�<Zp:��ͶE9�Ug�{��ݗ�!��l�d��4����Y���bkc�]�7��w��un���躆;�뇞�(Ta��{+����wV ["_��n ,�����;��<xp�����P��C ����� {gѕ0��&	}`v]�7�<���D���Lu�d{)�E�n$��uA��u�,�S�\5L>�^�ZV��^��t�2<� *�B�aW�P����� qS�m	�}��r�����=մ�(e���ÂJ1|Md���*��0�'��x���D��8*����!�����!��?�	?�"hw�����~���yy���q:�oݮv֌���膍��Ds\f�bܯ��Qو�1fMM��xi>r)xnT����J���5��,��=3�lq��l:�R�׵#�Qg|�ׯ�E��-�Q$��ߒ7u7�M,oLt��4��5�`��,��~�w*t���<���o��[�]J�2ze���u�I�|�e�Q`ޒ�Zzk���pD��p_���o��@οW =Q��]5ӎ{ҭ�ɺ�V]C�q�:~�{�.�v#{}�n^����\;�'��zT*<O��: �+���S�6
g=ESRE���M��$�,�=�ߪ@��yP�i�\Mz�	�1q��g6Hu�[/Q"ԧ;�\�}�^<��uF�����6|4�G]�*�ɫ����Z��6��,f��3���K�(��e�<7'��6��]1��B�T�V߀�U g��鼖�����T�>{�0l$|+4�����1���p��I	g��nA$`���xo�z�L�<��z���z�v\��L.����N�|�C]:��N��zHl�L��E��J�=�a���P��Zd�a��QxaQʎs�_�R+�˦*,����})��W���z���4}㟩�#O;��7�/��Q�����Br���&�4:��w+�uȵ"�P��d�N简�4��xe��*,�Y��d��{[������ T���n'��=4pZ�VƦ�y�#Ģ��x*W�r���a@�K[�\j8��}Enٝ����3{��r%�x]j`T�W�7C�L�lF�Ci��7Y�@b���J��3�&[�r�#,�d҈�~�z�{r�X����-�R�J�3�3�w
]\d�������u�ҿ8�!w���p�c'fm�x<��ފ[N;�0��Q�k=����� �p��29�j��#b�eD�˟Rܤ��V'7�I�W��.3�_9鞯����O�$���HTOz��!�t����YJ�-�b�/���dڔ�j<X���NF�\M�y%�a��[����]G�}# �1]ݷ&�����oe�0� ��o�\B,{�ݘ�P�g�j���}��u�{�R,[�pm�UjO���1�dy���;׮�/�!y�wpyU�Vn�����|z1�Bs��V}3e`��N��a۔2g�;<��i!�G?S�(uÊ"Υ�׭S��c�_��qǁ��Uw�
ɹM��g��;�[	V�����������%q9Tr��ެ�.�ehc���ꍴAf� �AF�YH��ܹ-}��f_�L����������L-�*�������`�=�4���BE?f�H^�n.�t�d�f?U[¨�ymjT�uP<
�렳7�`�9��U�%��58���*���'Y����2�"�V+Ƅ��9텧U������)���C,��g��E�KM��aTk�
�%zcA�hS��jrE����͵S�Zh�ɞ���B�hV�S�O��*�l���ɗ5 '�:<���/G�r_�'d���v,�����X�:��򱚳�;��#Ն�x����1ӥO��x�P�Y� (������EF����^��IT�
�ܟOD��d07��p:j-�P��&<���`Gw���d�z���GvV���tX��P�355��&;��g��H>��`��]�N�v�U�U��ǒ��1��Q��R4,�9P�j:��鯟'��<tǕ�Q�ª4U�}ټp��t=��� �^�/�}Lyb���zP�&�c��:Ԗ }3�v/{֙�����N���O]������S�U�^���;,�p鞍c�1\�d�q��+�:�`w�V�C�yUưV	�F�<�{���me��g 3�W�]���vT��,L����-�<��_i�/��U3���-���7'�Z�
G�p�Y��59���t�c��c;q�'�:�c���{������S�J4E(0���:V���$;�M���woq]_\\�C|�K'�ܬ�q��V�|#��i�5@l��iH��ލ��L a���d�����K`�iV��&+'�E�+ 	}�rw=رnM߰kU=�7�6�c��=	�`���φ
L�,�cڎ,38I'G:�y�
<�w�X�Y(oNx�񠇔�S���8*��Xf ͮ�Z���Ʌ�=��TZ��r�6$>��1��P1r��+&��.���2jec��]��'&���w6ʠ�R���@e�����ܬ�ٱҞ���5�dJt<=rΘ��TɉJu�@=Ȯ���w1Qi�𡽕3�{.�)�x��U���c��t��9u�)N����B��B��#���n �9�6�8u�b�V���:��B�*%��!T=�PǢ�w��s�����y;m�:��y���۪ j��0�^K����|��e�7�]�@��T�7��m{�ئ6g���w+c�C���Ģz@�g��@]6x�˂71�򧼵+��>)r���ǈG^E���R����i��uał2o���krM�{�W�,u=���3�F��ꉛ��J��eӓgvu�u���knv���n3ǈR��T�g*��ÂJ1s&.Pu�B�US�d�T;Ү��j�G�Wq�	�����#�O�(��e��q��
�>k*6$��t/S̞UJ'���K�<%��";��h����5ި�ϑ�b̚���g�)��y��ݴ�T�G
�Z�u<�S��%6l(?L�ug1Xp�,�����:���ܟ��h] _{���@]5Ҝ��\3bA����ʑ��#���<u�G��}�; _GW�:�	�>���x����DZ�4P�oI��/ג�7�?u���H]�	w]p�UC�F�b�L��e�$U��/5gʞ��:��fOFx�w�^nP����iλ�*�>�jXɖ���l7���v�u.��8�7�A\����ƻ�H߹M�ocxk����]��l5�3WF;O���Jr\��M��Tb<2�0ş��5N�a`����*���"��T-.���ѭ���d靽ڡ̧˺-k0��87��]d�� ��N��xCKMJ�t6Ȝ;���%"w7:����5��c�k�]n"q��=��t�;�-�c�sӝ�w��zQ�f���	��'��Ex����90��!�lv��P�[��-�P��40�c��ԁ����>���d�#:U
�g���.�E�
�Ts���YE��W&3�{��/5�W��"�9l�H�c�����F?�����'|_�U歾5�$5Y��� z6��	��M�y<����F�QR.���K�\����D���+�2&��+^����^1҈�n���Z�� J��;MT<��q�fă�g����NB����8���TT.!q�$wX�棜���Tc��U`�ٺ#5�"�����ڌ�^��rĚ:ڢ��˞s�=�!�$lv���������ߩv/p�����ts�� �ǆF��E��	鮞�1�#a}���\ߦ�ܭ=�t����yQ^�T0f��zPj=*�Q Ǚ�!L[�OD�v��:�n�D�fT�u"���
e
Rrhvq�dy��#�z���%Ǎ�?V5p��."�\���tKy���2>�t��o$��W ɹ�^A�/MͰ�����@ϯz�@j�b�׽�F��[{9JIh���p᧎��;[�v���7�u4��v���[خ9Y��	���̿�<�o�Uw�����SYX%�@g�0������yKq�����0ח��+��#im1c�,�X��syଛ���_>_���ö�C��}H/s�:���޺�����϶����lR�C�z���:��QT��TP@�twaN|s�ۖ��׬t8�@�:�ф���م���W�1����C#�4�޽�D繴�3Px=:tӕƆY�et�E�KM�Zχ�W�*��ƣ;��sK7���>�}� s��:�O3�]X���r|=Vck���������/W~��}3��?��?"S��=�q��^�`�7}�ü��ht��{��)'�~c�e���S��-�:��,\��=1(w��`A�wQ���]�^�Z�]β=E;2�.{��r��`ls��wM@��+�T'���^>��ӵOiF��UFG9�MDd�]@�_y���lI�� _.� �>��r����f�M�㉓�^]"��C(�Ml凳����qMB���.!+�*j����5κu�̧�#��f��'Y�H��DVN*q�#7����ed���!���I�쐲v��ǚ�L��ҙw�ײ4�J��,�(*�&Z��Vgk��ů4\t�ݝ��� �4�mB�	��f*��ˤ�go�e�]�^w�8���Qkp
��N��ъ\ς��Q4W_Ř%�o���:'o�Tγ���G8r�$vwF:�H�0�,xv�
}6^����P��גe��\�SJu�+�}�(�i�*�������B"�
�6�Qhgl�J�����ur]1�/P35V�9��:o5�]]�ʹ)K��Bv�Yn��;(�����ӄ�3�C���*;��O���(��+Or�X��!�;u%��Y����GĢGwE�:��B �1B���Em�4O!M(4n=[+�G��v5%Nv�*	���g�ۻ����y�t�!0�������f�K�-9P�{eoH�V=�5���W
(u�8�UtY��9�V}�.P�M^:kUtv��r�n��L�ٯ�te����#ѐ�=����L�M;�k�u��j�\��:'���aΤ��>�b r��n�E:�xf ��i<��ĳo0`8�l\a��5��EL�҂*Y�+R|���w���A�0�}S*Pٰ�:�`�[vɋM\�����F�n�s�\��ҋm��º'��:Yț�J��q�+2���\�P��Y�̽q�Z�R?[�Kqhaf��Nk��������xt�|3���+,n����u���EM�L6���:e`rF:�xBq���*V��,���І�����������9�4n�Z�w	��;>�VF��1Dh��+�`o"y���G���V��oet��JQ��*�"��0�6�b��V���֮gQ�Y���Ug;��6�t���`}h��:�gh�&��%a��Y�n`�G<��Wm0p�͖o5�-�K9��(;���-֎�q
���=�7d����;����}t�[/݄���9�E��ـ��������NV��̹�//�heWbw����s�Ӊ�!P���wP<
O��& �����淕���_w���M��\�M����I�]G�CV�����8��c�������7�pt�:�����R�h6z�.?t�>� ������������/E"��艘X�:�h9;3L�r���̳_h�O��*H������Ź�J���gC��5d���
q��Ir
�����.y^9;�]tIWuɹ&�b���J5e�Ԩ��U3��L<����=#p�6n���^y)��pX��Z�T���<B]Zy�=�/-7q�g��f���HM0�<��u'M�w/�l�r;����[�����à��N�Iu���(��WBD��C���t�t5��.v�FTN8e�R^dFaWN�M�3X���ZK���y��N�^�+̵�CҜ<%�9���.Ty;����;�]��Is�������F�2�U9�%	�U-���G�"rr.�g������n�h�Rt�M/<=�����aj���TT���5�v�:�n�����N��{//0Sܕ�
��\�f���p널[Z�9Qh��<wp�v��$�/�Gi��;6l�LK<���5�HC�r�3�K�-;é�a���%����Q5+Ğ��T(ᕱ�ulv5y�|ӣ����l�v[��]���q}3�����4]���Tu�T�=�&�ʅ�Q�X���O /���U�7ݏ�{�]�Փr.㎎�pY�?TҚ�JI��@���%���Bǯٸ�n��9�������=�͖/v�B�6+%�v6X�\������K�0;z�M����s�j���''�6*�����{ܫ1�T�k��f��]��;�Ԁ��n�J���[8!+�CGޙyN�zK�}ϻ���-�קx��}�y�zd1��j�7�M<����W�-�G.������O���<b���,{�'����	F�X�:�{p�1�]^$�.��>YZ�B��ׁ�T;�5	i*p
UP*{Yy$>��Kʨ{%9�ʙ�u'S�ܡ�~8gc�s+���w���:�)O���W��K��۾�W�{����y�6ЎMV�y5�W��!q�
R�������si���3ܰ�~R�.wk=�g,b��Y��uCXb�)�v�OVS��^:LA��k���R����ru�C���'ܡ�l�N�t���8#�S���Aܱ�֭��jfun��Z,���Vz�w��[B��[�8��,`�S�5s��ӸpfT�Тb|���h�e��,>��;�g�[lzk=Iu�5�\�np1ㅊ�pKF�*�w���eb����	�tw v\uA����S[�	�s],{$�ϥ��c����m�S�iVNc q���Ƃs� l2�tนW5
��^uB����9�^��������03��Α�R��MS�μ;,��#2b�_:�T���*�~�c�����߿Q�"���fg�Uc�#��������f�}~�	,U;��ЏO�������4Es2���Qو�0�G+��U�u`�nq�>,F����ȹ��68�}���hc�;4��Tż��<���D��εq��{*�F2uǩ�=���z�� w�T3bA��#��u���,������1T?F�7��L��΀:��6��b�yܽ���(�t&t�c�� �Bt>���P�է;�%������E��q#�������Ma(��eVu+y��ۭ��q�s,�>�'�N���<�y���#諁GW^�ذR%����#X�nP[C8��g�����X�������~C�>\L<��1�O&tH{���Ǡ��k܃��m���1�Sޘǆ=��)�gF�Հ+*��b𖧭?(�Yav���X	x�B���>sQ�Q��S����.`v]=���?~�es��پ����R���jz�Ձ�>(�y'��E�.���[;�%��S���{���װu8����s�.��pW#��
,��w�z'֕ovs�D�8{I�NW�5T դ�#.���
{���
k3��v����չ��)�#���R����u<�I�8d����u�ʥ=UW�n�5|ߎL�7��5��s#� z��\*,���OL�O��)�k��1O:/cf0�mx�q�˨GFw�R1s�<o��N�P������h�ˎ뎹� �v��N�-�s��X��{��jfy����!q�#��:��T�r9&�;+mYχd��ՠV�5u���V_F=�vb:�ф���ݧ�CV�{���f���3C������e�Z5lF�C{�t�Zx��N�ɝg�����g
���^^��F��cN������:R�NN�~9[uvG�V����t6pI���u�1p���s�=Ȑ��#y�6A���3�>�]l'����+�?j��H�����5,����#Q�=<:g�W�:��`>�U�ƭ��?�2+�T�/���捕���oe�N@��}"O�׫��Nx��bC�ѽ�Z�{ۥ���b?��M}r��.<��7�G{�[[j�(��QW�=�����28+��1z�x,����ؖ]�ܡa>�yWУ�feZ�W�Ӓ�����`�̱�1M����]��[3<|�t�[�稭�2�ے�f�a-M�<���lT/2���>�Q��S!����� ��F@� tWSa(.����U���G�GqCo2G�q]���U�F���|}L��H��t���E]ڥ�\����a�]YYƷ|z)���������͞�T��� 78Ox��O�62|����६	�[J���1��F��^�A��1�4��%fV�N�D9.�[���	�_,4��9:����_rGWh �ҷ$𕒷��;'����:����h�y��	���1h�0s�K�m�����T<�:!wrR��t���@��(ɼ�����'fLAt��a̧(o<����׮=V�ŋ�t]<zx�2�)v��o�qw惡޹��2�L�=<mKm�8�� <��=1:;��!�P���x�S�{�V�v3��OR�a� =g~2��� �(��;�3cDN��~�cV�=�D*�!U�H0���B�|�+��no��c�r'�`v�N��gc����~�V�s�MeG^eHвd�FT'<e��L������鹞��34r;���ۯw���� �7\���Wa6�E
�����% c:�#����.�~��mr kFvz&xeD.��=33�����3 ��6�?۠�7��_~/�?�)�q@x����c0.!��1�#�؊��U�^�l���|�C�.M�_������ީ��@�\mGz�� ~Z���+a������X�ɗ��ʥ]�u���g��d��@צG�oTMS�g����I��hj�MQ6#���؏gR�m͍��樈(�N��45���2��v���z`z�'���@~�>)�u��WK��gb�1�hJ��H�Ae�����	c��K'e𽇯��5�t�w���:]��I���/a践VS<�p9xz��b����E��\�A\G��j�|��1��}��+�/<���n�:�����G)Qj����I��F�+�����H��R{��S,~ö]~:2���`t2���m��V8�V�S�ܷ:}u�LF�<��o��h�6#�����5���d�*TSS��Ǩ��]�L�w?��}����&Vu�����8A<0WN9����.��S�k�
��Y}�hx�fe��<��1�UՀM;���b����z�1�_\���NU����X�<�T��mQ�O�A>'ߌ��B���yx#I`[�.�����UO8d{��|��x����;���#~0Y=T*�Ψ��5����w��w(�����<Ytzh���^xpI��9�l�e�~x1E�X��}�gW(<*<:�q ���zH����$�*�F�S���r$�y���Y&��ҽ����A��7�"�_t{q���q��P����k4��ҡCfO����7����C�e�+tQ2�Ȟ��l��_pα:���K8�a��*��I���~��ο�:�T3�ƺHo���q�!�R;u��ݾ�W�ej�Ԕ�]���&������@)=1q���Z.g�hq�����M�<\��r�߰g}������5ʚ�. g\z�����K���!5S�L��&ǹ%�۽��w*F5����
�p�g�w��1���@Et�.���+��K�ǲlP[6;s*G4p`��]q�Wp�	�1xz���!�7i[�̪���z����(��/̑}+�zb��������o��T]��ֲ2�ƺg<k��9+���6�Z6*w�<�_��g���]�_]ߏw��3U����{6@�����=үM�+Q�E��1g��G�u��?B���Wwj��_d�z�`���)ɼ0��������ز�
��Q�],��ܻ7���z��<��3��@]�"�����3�I�0���_��8%�ĞQ�y G?���d[��喝��%�K74�g�*�ɣ@e��0d�ǲ��	w��.�?SL���X[�1�\ݝ���R�g:vJ�½���Q�\}Dʘ�1�YV���k_X��-�Ph�}y�;F�t�E��[����|񑎪yؐ2w���z��v��m�]\�S~Ig�y�N��G 7��
�{�\���WN���<煮H�0w�>��y�G(���Z`9��e�?Gq�9�L�J��7�C̈�q��魃���~\{��H��,��fc�v��q�$q� &��ԇ�D��
�^[q�[�k��`���*��M]!¢:�L�Ӟ���Csq<hoz�'=C���K§�<��T���0�.�&�e��}�����d͹�p=#2�韣�ײ�}ڷ�Ow��;��dx)��7���e�d���;��� d���%f�2 q�K+��Z�D��:3eT��U�Ȃ}�
Ǣ�rx]C���g��,�[��e���ʻ��t�ֳ�Jdt�Z����fM	e��÷(]��1��}�ǨomO}��z�I�<({�MS�7&*ӯ�M£�f:��m#�>�ww����=I֨;�:�g�����ͪ�>�����ܾ�`Z���KǕi�L�[55��n۳�Ï��xS�-���Ǽ\.�d���*'DtN��[Z�lfv''�$F���yFV��gN�Y�����Y�3�73�y�CsZͅ�B��Z�>۝Q�ތ���o�o����C��w��z���uM�a(.���
�ʠ�h�w�`��1�����@��έV2�=Ѧ�k�d4n(��#<]�
�\&��%��,¨�^�yψ]QWw��f;&�*�Ђ2��l���EuPWՋ�)�'��}�� ���~R�ɷ�]xTt�L��J騺,T2S�3�r<%��n�X���9�{֩�	a�3�����D���طp�$��(��x���/D�Ί0�vx�"nuz�)ib�J�=rT��˃,��.�Ϲ�E�!+��LT�&g*�#��!�9���D��y���� .�1�;����*�;\{�9��+�y܋��V��*9eC�23edɨʄ溋
fzr���5z���o\�rz<O�`��G:���_��%�������<W���_���{���7�6��Z\��;2�B-��J@�O���X9�4B�^r�W���Gh�]�~��S��{�H��&� �+�1�}�l:�쥹�K�H����2��6��ǫ�{���1�'C��X�{^IX����TO�	���OL�q�X�zff=@xX�mV�xlVO^u����5��z�����<�J�V��`_Ⱦ��1ƣ�؆�fnvQ�0mI�S�](�����e���{�덨�i`��)������ϒ�X=9�������o3����Bs��҆m~���� j�#�f�C�@�t*�|0�R�0��rAn��B��aKߏ\xUP�L<<��x���X�:�d���vr�j�%�v0^M�����ѨKNE#�*��
��8%��0��>��s�;~ܬ=�=�J��B���\�1�%��9�
��@=*�=���Jx鳞w�wk�H,}7�x�<��ެ6�����T��)����W]\s���1�O*ܻ��/ǱLvf��՜
����c�}D�v]B
S�x"a����5���/mnW�}���%-�	D�w��Gy����Ɩ�V�h���;��1�t�������?��s`�`����@�@�U�����Q
1�Aec�+
T�D" �
(�0�T��E�L�D�B��� *Dd@ �B)����0�Lf����`=��0��bo�!>>1���\<� ����r�B���&f���7X���\��k�%�ռ�6Iؐ�qe�aV4rh�W�n�=@���5U~�1	%�����9&r��_���:>:gw�a���Q݋�$o�,���2���6ŭ�>�"�E�T�.��/�� ���z#�E��G�TY���a��_&"���3zj�YO���jM@AzY�aZLq��7`BB ���&��� P@ ��DD)}FD�W[)ϫ�CaD� ���t��(�/�F�܎Eo]�"��(���a����K��W���A��wKǝ_��`5@�@��P�Br���G���;y�G��*c:/�JвM��\%�w���yDִ��r�=8�J����<[MGA'q]�nш|��4K�h�2 �$�N��@T.W1 @ ^��̺�4s�%���=�ť@��`�B�S��!���#T�>EÌZ
� �BB���r:B�aW�BwnC�ÆB�� �܉A{��KDB4�k�qI @ ��:3:N��ؙ�1g��6���������F�HF�`~9��'M�c����o]�pzp�N���5$��o0���B�y���l�@�� ���X\�Ԉ  �y�+���ϟ4�_����Й&�X31��	Z%�5i#����	��|��N��ׅ�J���nȎ�O��e��YLzh�  ��fP/��D��
�Fw` gF���n]L�5�v^9d�P�zP^�T	"с|H;#���2m�v""��oMIP�MCn�ZQ��[�B�ϔ�3�
�$ �<��]�Z찿�w$S�	�ǣp