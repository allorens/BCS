BZh91AY&SYi��h=�ߔpy����������  `�~>���    :    �  Ϡ�j��*���@�`�TDZ�#�  0���� �    ug@(A�ww�۷Zn������u����ϟ}��z�����Ek>0{�y2����w����I�lL��C���P �5�o���ms�>�p;�Z��v���<�a���n�]�o�k��M���o3�u�u��:ז���M� �  󾻝wۧ{�w����v�/\�w���뇠wM���q�o�{�m���|=�����zl���� ��{�_v�3pb��[�c�{��/��;��xiJ����|�W���g6�V�{��;���{��}|  /�޻�z�k�ֻ�ͮv�����w,�g�_}���|��i����㾾�ٶ�         @   jy�*TFM=�#L�	�`=4�"jT M      ��P
�F#``   �%UF�� `F   D��@���0�Sȧ�Sjm	��l�OD�2�U�0 �  �D� ��P�IY�YE$dD�	dQ$BD�}���  ��|�\F�T%|�?ߓ��H��?" ����K$UQ>B������������c���d��փ�|	�p�����"I$E�T����1�m\-?�� $v�v�,��c��I$�5>0���r!�o���a~����o�߳TJ�+D��So�J�W	��Q1w.N��fIل}j��]}�P2Pd��0�B���KA��[h�5�Z�m'Re���E�O��Ȁ6�(�Ġ<8%��YX3X1�H�Ib�Y'�MV�]$��a�f�aA�>e�D�%!RU%�bC�A�c�����LPS�)Z�4�SJ))�UR��*CT�
���?2
����2
K2��)�i���%X$;,=2�-YH:�>��,E'�ϰ�	�H.�4$<,Xvdk80[8-�d�ZK`2t1���l:���RԘL�$ �~g}��)�P�:K�+vVr��^���ĻJV�M(��%�&D���
����2��/��2��M�(vS�*vS�+tS��%/J�oR���z����b��thc�I�+�����N(2n�6��*�4�ƒ��cC���T�N(�X�@q�4���MEzy4�� �J�[K�e1��f2�l�r���k%V,D�[��pK�&C���D�D
"�C������0�J�!��Mz�/�ɰX`�&1����)���wH9�C�`'��k �A���I	��J!��������������L���r��.��.��jM2��0ȏ3��HT�A:J�]�A�a鄭�L^ZV�-�W �)�ԕF��I��Hs	5ey�?�AI8�,@l�L�A�����5�T�LE�1^��RD8ezC"C"<�A2�N҇�1Ki^��f4�T6I9o
a��`�b$0�+�W�	d�d���K�&C���A��B��D0-�,�,�,�P�j@�B	�0�y���w���b�N2dS`�4Sh~� 粉�*�Ƞ]��� �I,�_��j�c1�Z��chX�`~��~b����}+n��+l�ٷ�k�nn|���4�01z�VA~,
����b��S��Xbރcch0���H�Z`��X� ;7с�b��A�C��%�cX{����\l��.EXR�2�"k�1x-��n~�Q([F�Z1�p�-��N�Sl�f$j�:+J�5&����"Y.�m�g�i[7l��^�2�V�����R��):�ZAE��哔.�9�	e��{'܀F@9���NH��s�D��3F��`7�(Q*�`������r����%���?6H�$X� ��C��&A;���!�!��C]�00�Aփ��$݊pM1N���-&jp�2ɺ�M�F2L{Y/C�%��[�&�6$�&IZ$�+&錔Lő�23:s6�ٻ35IM8)��1#}���쓨�$��N3�-:��i[4�[�U�92���5h�/-+A�yeS&�-�KW)9��J�%D��-QF�izҪ�V�vIfrA� ��TR�.�vq�L��I���$ƣ��EV���E2	'��Q�5D�)�vl6m2��������1e�Cf.Ɇ�h�EZ1��Fq�9�xI�&�Ji'VT�ز�tI��d�
�ZibW��*p8:�2ɶSGI�j�Q!A`��Ң\��xsY��ݝvS��
�u2Q���e��Id�K��&ɪEX$<!�Vٛee��Va7e]�vS�o
l�5:L�Y,�&�ٻd
l��-I�IƤ�
Z^����U3����:H���d��Jlղ���Q�7grҷ�cԵ�OI�ԥ�	dBAa-IQ4a�,Y0�2$h$a7A"JD�S���u�ιIE�����h�Ej7��G�25�MKĖ4�h�E��4�4P�%��RnyY.�5Feܕh�"���[e�2�ݢF0��CW�tb��� ���N�3Q�C�gL�'�F`U�;.�Y��$i%"�$�q�)i�:ɦҶm���Jre(���bm'x�����$�����J#Q�)��v	�i'�Ɩ΢�AM��%��+$�2��&]��㒙:�-&{)=ER.�S��(3A�LشYWf���Gl�l�p-2�-�)Y�,+C���l��u�Ģ�h���t]�j����IU��ʛ9P��ih�K0�KM,J��2q�[4q(l�F��j�@�	Ӭ��U����7f�벝�xV�Y,�%-0��E�tq�[$6SGI�j�@�	zSf)��I���	�*�˲�xSe"p�K'I�h���A�E=)�l�ԜjN5'R����oVˍ(�� � ��A���қ5l�gq��n��%�q�[4��)�6Z��!,�I����,i4�2$h$a"�.��)�-�X�IkIkET&�+Q���8�-p�	Ab[��I=E4[IcIcE9:�&�+�I�ౄ��.M���l���eM�D�YsE+��Q��pXxX�Θ
��J�p�v]�>p!i�Q??��\N�vc���6 ���9p,+�)hKB�B�$���+M�ѯ�j�,�G��`�I5�^�L���2f��fNĢ�ġ��>+SP�g�`ׅ�M���p��lVQf�+�v���6P�����@(�|Y�Y����l��ݫ@�e g�,n�������Y_}]<t
4@(��Ś0��O;00���U��G����Ϗ�����0�z�Y�l�7UAg!�]�: |a@n]h֪��͜6L�>*���$�L|z�fN=�$���?\��8B�ou� (�8X<p��u/���a`X^�!��n
�J�N���5�gr�4C��,�E�e�k�����G�J�Y �6o]�UU=ˠbzrvi蔢QD�: %f�<(�� (�ӄ(�(  !GJ:|h����䫟�兜6g�*�F�?k�0l�C��<s�)����:;)NĠ'E/ѝ�+0��t��!D�*�<Q�� P>:4/��� )��`��F�/��ښ�� �骰/��Q��"#<^�����]q��I�F��4N!�g�,���4CҀ�n����&���ㆄ�ǽ|�]�����UE�^N���v��^��!��}�6qo��p����h�!CF��= 0�9���������l��.p�7��Q@Y�l�!�Z�X0���ߵ��d�8L>0!�O���]����� C��a���gj͘t��r���� 0K�}�6U����ĝ3�~��r��4٥�UJDVkj���Hh�t$osU�b���g��� ,!t�?8e�;���@Pp�:V+��j�{I���@�PY��4a�Q�MQ�(:L,.���(��CНQ���� z�F��D�?�`��6t�+	����_�O3<Y`Q�j�%3�vn���s���#6\XŇ���Ç���Y����(h��f��(���0
0�>��/�Usu['��F^W� ���ɋ&� 
�Ut�U�Q�����u�o%نr����,[֪�����4 ||hϷ�9�@&��B�ug�l����Y��	�L揄�f����� w7VttQ�gC=Th��p��ٽ�Ν,���x�6t�uuTR�ށ�tj�`���3�M�� �b�������ֵ�{F��{>0}�UYe�� }�+�y�9��ѽ�Z�p��׳0�0�l�GHh����rV�2t��i�I�ʨ��َ[͝��ek���5�f Y�xifO(i���
7�U��cE�!�ӯ-OM m�҈��e���+���f���uz0�h��3��0lɬ�S�8�tɘ�Q�$����rJ*��wG���#
(�+J'BDƃYժ!�bkG�p��U��(�%g>8PN���m?��f:kY
�醦��@>�$��r�|g�=xhê���_�
 Q���t里Rl� ��t�֔�4�J�5�r�Xl�j�] w5��/��8P�uI�`f�TYx��W�uvP�JPn�YҁzZԀ&�l��R���_�Sx��U�_Y9�&N�1D0!����*�;�����D� 6r]�M}��<Pp�����wg8�����W�� ]r_|�����uE�Y���:����g5RU�,�&�GƍL�X�<pob����(��[�^�<h��@{}�6?-�(�g
_u^�3�e[3�Ƽ����<�0��3=��"b�M�ªȖt�CO�&�u|,�U�l�S&��W�Y�Nra�S+�L5	�@Ἴ��K�K�r�`�Ø�A��eL�
!���ڠ9� У�K��@�h<���U���_M9��.����>��X{~��Y[��͉>*�p�J¢nDP���Krb�$)��L�I�wݢ���\[�:|Q�l��ù������Ɋ<l�~:|Ne�ݚ������<M$Ô�y�ų^�v�[fD� p�,KBK&�6=�-�z��M�J�`;�, K�6|p���F�?��M�]@l�{Q��xI���جK�\�<.��]!�E�9yA��gK86�ad</��Ѡ ��XK��@X� ��х ֮5�J<xW��� 64��P�!�[��($���(^Z,��Y�(9��)�R+�JL���zc\�3�	:�	>���'�]�������M����R���r~��!��$|͐�Gȯ����>��H�J����A��*�ԥ�	�GC\0X�JF�KnKȒ�%@@v�HJ�E*
(�"��� 0�w@����-,J&ji�X<(����
ӆ�P�(�(>pM�kVj.��'��ϵOfű%Z&piP�]R�Ԩ��و��O�ٔZ&I��x�DB�\����� �4׳%ֈ�T�n9]�d9&
�rA2s��{��6��T�[�qCI�Ҫ�wj�jB�#��Z8���J 3"Iyn<;3��V�$bky�	�cͣ�H'�P�B9��b�B�9�����e������k�M�$���o�&4B�53��%��S���dQ���Il�'�Ɲ`��ԩD�2�3v4�湅�0�H�5��T.|Q�QjO�Rݥc�v�1JV�V�`�� 5K��gbT�W���Ȇf`"\�IS"r�ՎX�w����|�%�Ѫ��T��<X�}a�#UR��T@wGp$Eq ��h�1�`����}�>m}$�*����Cφ�����d?0�/����K��>�����	S���j����w����;2�n�n[-����m��ݝ�Z�m�-���j��[m6�t�-���m�޲�m�m�m����6ܰ۶�6ۖ�t�M����m��0�m����� a�H�������L�m�A��n�m�m6�m�m�������ݰ�n[n�j��6ۖ�t�M���i��xm���m����m�nm�m6�n�p�n[m�m�m�m��m�{�<< ���H���Pۧ��l��o[M������oun�m�L6�t۪��y��6ܶۖ�t�M���m���m��a��m�,6��[m���m�m�m�m�M����������˻����m��m�-���6[owNh��n��-��o�����n�p�m�m�m�m�m��m�l��m�fm�z�m��m��z�m��6�m�m�m�-������ou�nm�a�ۦۖ�m�����m�ne�����US�a��m�-�۶�6�t�r�p�m�m6�oi��x�6�v�m���m��a�����m�m�{�@�(��oHm�-���m�nn��ѻ��x�m�m��B��ce��oXm����m�����6ۖ�t�n[m�[m�m�m�m��m�a��m�m��ۅ�a���'����D�����}C�UD�	$"���}����G� �
���G�|ϙ��2}f�0��:|�;i�m�񷭛|���6���v۶����f͛Wn�v�Ǎ�m�M��b�lٳm�m��m����+����e>>6mҶl�����N�mۦ�z�m�z��f�VͶ��������ݶ��m����޻m�lٳj��A����P��A& )@���H.n![�bf��l�(��5٦ }� \'�N��t]]�k�S`��n����	MQ��kFS\�m6�_~|��%���]���8����k���=�Ŭn%B���F����]�*�iN�B:�G[�\�B�RR��lb�e�I��ð魆�32�0�1��m�����5��JG1�
%2G/Q+5d[6�v�h���M`8��l%TV%�ThYf�R�B5&� ҄-�	c��eT�m��Ul��W�@�ee������RX.l3��������˴��h��Fنk�K��`��mw4��k�1�m]��c�a�RQ�fe ��=���koR���_>����b�,]^�
恔E�l��5F��ĬT���so׺�2�0Yip��t5n��~=w�[eXk�e�44�32�e��dt�f��jM��
�ۂ2�~��z_-����0�ឤ]B�[��u�é�x�-`�s��ԳV��_2�_a��m��	m��V[��!�e�ۆ���mh%օF�]�SMuz��र�����+.�h[Rls����V��,&�V��Z\��[�C\uBJ�F�;av�4*S0���݈����ul�(�WZ�5aI����iK,��ZL͆ٶ���G��*b�I��]�Qj�0�z�ͺ�;j#��V%���j̺�<� h��DC	d1n�v.�4:�kk��6b���`�kll�iH�A�eCB�m����4@H��ʒ��X+��-�n^a�m)��X���\`#��#����ۑHbk�j�Ks�L�n<��lW��o jWYn�
��B%�h�w�cp��
�R��lӼ��ie�i����V�]��|ƭ6����t4��h7 n��
j��,�ҁ���1�l�ݻ���t��Ð��w���HR�D�Z1��]v��V�Y�[j�����鮽I�b��ɻM5*��ġ\�Yh8n^��R�pҰ����YD���x�:�L�R���������6[j e)Z�0LV�4�rJ&��K��hv8�@�A�[�Viq�Y	�6��+4��K��{\[n�0fZn�Hl-�Rgi�\����ֺ�-��E��anڭ٬l 8����� E�0�[4э�\�t- �Gm�*�Y�XA��ɲ�RJ^/lR�c�&��Hጹ��]M���4��ݺ,�L�	Q�
]Q��+����ZL�F��P�XlD�e��E���6�K���h,��R��l��v!Z@2�kl��ĳ�ɭ�օV٬�4e��X�;�u�Bm��˥��Ml����aF].�+1%�Vf.��J�>�鯠�]h=k�3޴����Kv����̻��j:˜]Md�6)��1�a�z7_\]G��Yf��e�%�G��.O���x�BY��q�:�K�h��Ҭ�e�wn�]n��r��m�f�E��U�l�3{iZ�l�דj��1�,
ôL�>����� p��P����33������oq(p��陞��s��s��]u�\"C���s�û��g*����ĩ<;��ffpx�N�*�g��2ߏ��a��~�ם�N�I��6ɦ�� T����7�Fa��-�7P��E��#Q��1ɺ���Y����i�e������f��v�h�P�:\X�,\8�mv̆�[qE���s�V���t6��v1��b+�\��it$fڡvvҸ�v�/WX������HRf�cj\��1� ,ك�[��mH恲�m�e�`��Ji���HU�ۢ:۩��@�f�G[j9X4Ku��F6�
@�D2��&f%��R�ZM�j���X�m#�J�t�(�cZLAD�$NcXJ�5nf�v8���7`�R�B�"*�I�L̶7��!XH��
�a(cTE���3X8��c[e�s��XU��F~����gy�	�����lrD�*ING��G�(�bj�HC���:�y�Զ�o(��)�4�f��"��t��J�B{�4��FUx��f/g�l0����z�T�S�Dx�i����4��������Y��'9���C냽S�Q�kk`B�a��0 B3�%I�[k���G���V�4�1���1���I&f���өC�3��-�����&�$	�j�؁K*(TNԶ�C]��l% r9�Nd��i������4`�!C��M�:�:�k�銮�4�1���1{ld��%�L���8�(��TJ��H#s���\�;��v�H��gd��0�*�&#m�����p�i�q/5\�.��N��9�2�v����a�/]�M*�m4�1���1�V������W�Th�iP*��RZlht��*F�C4̽aڮ#ixdK�%a���4R�$�V��K	��%�ba�@
]�	fB9MaU�b�>t%�� kO|� ���=5��;\hIb��	�1>&��*T��Q��w��@�LkMR�b�SC[kϖ��u�*�BZ呔��qWs��ղ��O��_N��V�4�1�d2PPQ2BX�c`fH�:w2oZ)�(Æ&�\L�H�q���&���g��R	�}�)�M�K�� ?i���0݈@�MZ�K�cZb�շ�]L����Ƙ�:;;a�2�J�8H�'�n�`R�P�׉v8c�Ii:i��M��o\&f����q���^ӹ�����B�>��a�̬ᴣq��
K�����/��>�z��b�����@��BT��0�6�M�4Ye�Y���1�VRw:�f2��3Y5��2�=	�N2l�u�VR�$ dS#����u��#�[\t֝�h�h�ióN��t�bӆ��������i��vw;��n��brx�mVf	�+/��Br��KӀz�$�԰wQ�3%�M�8̌n%��)�&�T�[&��� F &���6Fn1H�`��lJP�X��	�@e����*B B��4[{7��uZ��l����iO=ԍ�J�s��Ig�w�􇄖ڮR�fV�yE|�jʲ�j���䧭�Ye�Y�ә()�����9:�}]��[L9^�-[�ǮGOOZ}*V�]��Zz[�h�!k�<Y׷�ȺRN*"��(��[kMs)p��ƣ��kOꋴ�G�����'�w�%�ah"�A����Ap<jIh��E�7�\������'�`���r(H�p��x^-^�qs�s���9�fg�3�s�s�2��f/�-^���5򸽸�/��U��m^*���1\UY�Ζ�*�j�Y�j���x�8�^/���K��\z���x�W��g��Lb�j�-W�g����W�q������*��U�\qx��/q�;W�3��mx����������!�� D_(�DE��;�L�M9��X�v�5�F뒁���F�Ի���kSKj��ͭ̀EE��^yc&�H7��E♩��`��}�M���%z�W
��7��@�s�%I����33����T���S39�z9��{��fg�wP�q���OA=ǻ��fs�>EH=ǻ��g�&K,��0���[rt�U�S @�V���S�����'�ǲ��Ƙ?��_-��$��ǩf� V�Q���7�W�ϱ�@�H �5**�c�R�4�H� �q�JH�JNZ\y(>��,q�|u$像�˨�\bpKi|�zD�aI�GĀ�!�:-=!���Ґ���e�Ye��Ǡ�I
��`�x @���1:�1)�K��bSä�,�;d�τ�[B�`�֗�5ԥ$&��������BCl�W-յ��CPms_r�E-/5,k)GZX�H�J�Ej��R�쯢ǍFuv��aq���[z:a�Ӟ���nu�H�<=,��,���ނ�$*t6N�ټ�k0�֖�����4��Z�IU��:��\__�E�(�MV�	�[,ff��K�Ég�����[cGks&���>IČ���6Ch�낓�-�UQUi�ONL�\�<�FXі�1|)!�%2��#���t��"[������{]��h�Rq!p�R��_����X�)M:J[<̄�>�2q�y���u�tm��"�#V:U�����&ʶz����I��N�Ye�`2tJ
l�ss���컸cP�����\1�2���D���,S'!%&B-&L����bv!a�Z#$��	��g�.sK���ҴBL/v��Yu���c�	�M������5��Sm���b�DN�3�zæ(�(!V�`��I�M�R�ɰ��Ve��Y�mI�,d��J��Uq�2����=2;�����c��H1�^��(��e�Yn�O+1Zc�]ٮ�U�V�$Gipt՚#��ipL15��wJ�Hr4��F����_*k��hjؚ�ՋШ�H$T*�E�R��Ɠ.�6�s�W9�̵��<t����jOe���<��S�:�Tt~����i-0�RUT�+���ȞE����&�c��q�֚i���x#%�%����Zо�p@���I	Ko<��g;"�1�	�Α"i�GfO�.�e����`�0���I	]�l+	]2��1�4��,�H���F 6�a$���Q�Co�Ί��9n}�d�{��{m�oQ�cڷ!�I��|:�$��Q=)2���i��i����a�+Lc����������t�p��g5�I�a���kء��������Bbl�.���N��M���붍��-��P[i�e�ٱ�c�b�D�K)�M�u�.��"����Y1��
K�O����	��l���Y�(��M0�K�lG��UUUEQ+I��E�m c��K�'m)0�N�L�pD���T�'��0u9	MS�l~hL�F�0P���U��A躁��˾xX��N5�j6��Or��$�� 4����N��1vY�!$�����,��e�Yn���+1Zc�yr���g���N>�K6���K�e�D,��I#���K�: r9-(�7��9��)%zxۦ5_X E��o=@u"�1IĈH�������J*��UƼly����lѩ!i�">�)b��>j�����@RB��S��D=!D�k�#b�%C]^A�B(�uc�&F16iǬctl����3c]�֫ŷ�4�Ɨ��:��k0���� ��):�$m�.4&�\�$�5�(H��&�331�'S쏬~��*��(Ԭbi9I����
���)-C낓� w)5��J��UwY0�$]�7�
M�ᢓI�b��TZ@)�+�ԟ�O�m6�1�GǏ���0�lrţ�1m�r�WDzB��W�@�W�i[[j�?���_;�o�vN�=UQJ���lk&�}�E�hG%��qxp�6�f��
L`��Dx����,a1;��Fu3L6�d�h��_'$#��P;`��>BF�éF➤��6t�M�?�o�C�#�[�����:�B�cB��ph�Z8/p,�	����˘��<^;gK�Lq�1x^�e^���=^�3�����<^v��x�i��/N2�����x��x�/�1��x�����ܷ���ʮ-^��K�Uqj�-^,�Ş1Ƨ�+��lz�^׊��q+�8�?1�t�Wk�zV/���-^-Wx��V��ʫ��}d���g1����8�1Ҹ�6�+����g��Lb�j�G� �0��B��X��P��!�B3�R�S��m|YO�Zū2�$���2�O9�	Z@5�2�[ �������W7��ǳ -7Pb��V�!]���f$�&rf�D�U��\W�(F�㯠���rv�ȶ&�Q����$G_�Ll��٩��}���o�w�[>V����ڴõ�"�����	�8?A|5�R*I����~*ff�|������fxs�W�S��s3ß"����}wU<9�)��]ݗuU\9�*Ow.�˺���n��4�����VO��k<W�R�F�#�r�f�[m�7���ea6&;���R6-�LkuP0�7�6���laJ9rm�L%�Uu��i@v��+]��j�J��+�i]M[�+Yf0m��Iu�.�h�Y�Z�{�O'
���R˄H�J�H%�ٛK����u��DZ��Q&&�p��t��[e҇��`$���.��	iit^��`�(p�en��Km�< ��]���i�3�qNs))6�\K�\CB3�U��!+��SM���ch�88cV\D�k5�X�l��_�t/�U:������3,З���-q�e�í�H�6U��%B�f��T��3"ؙ�,3	*62л2:����s�0$ C"|���V]��������K�B�*�M>&-æ�Ǯ�M�k�LY�҄��I	�:S�`i�G���e!zJF[ADpCݐ���i���HM�g$��[w�O�v��.X�Z�x��9�:ڶCgd�+q,�Dc������Ɲ<V������d�IQ�H\Q7ბ��RU,�i@9��������8��$�q���E�$$�8����2c%Qj�kQ�ڬ��꼨d2a��ą�$g��sJ��TP(� v��Q��Q��P�m�*J�!��$b<b'�'+��O�`YR��4Ժ;x��1�g��´�
6D�A��	+I*8L%[�,�!rzB�͐ܦ�OS�B�@]i"�L%:N6��'���\/�ue6;+��
��D:γ���6D�$�s�.S@`�����am4h�H<� Z�����/��!�)!����6��HC<r�m�<�8�2~X�X����Ɲ���FBYc�vgg1��cy���8&Ȝ=M:4ݼ��4FM��#e��$��u��P�.�F��TP�;Uuur]�Ǳ�:�X��Zf �n)R�X�t� �oi�%M�`Ř�F%�g��ZH:�v�M@��JD�1�����T�4iL%���@1�2�[N����#f��wז{h���1�:;=x�+M1���L�]8���qqFՔ*"on��Ջ��$��<�[��\T�MVmWVF�B�)M�f��R�i���n�����f�b�����Uc2��+d*U�R��=��#��i2¹ՠ1rI�,6f0�:���;*��8�iL��$��Z�qN`MǨxbBI0��Y��	��$�wm!�A�|�I	�o���3O[sր�`�o���W�VK!v�HC�	���% e�zqr�.]ͼF��*�i����2����0�\���.��e���5�e��ӥ'X�<�KM�I-�ޞ:��sy+e�imbL�O���G��H�m���Ř�.4<ϕ5�G9�j�QC6��3�瑪�ŏE�dmF��O�b�x)H���H��(l�24zګ�N���V���~*!������M�A|:`��^`���*= ����1�M�����bDq�I���n��B���軕We�1���@m�4��������?L�w��]�:�=@'�I	`�τ�++7H+�0̠խ{*���]���_|���!Z�l����l�!��+8�O[#ؽ؜��qQ�j�4��y9�d%�3�8=�Jbc���&g��j(�S����OS)�i݇(�9ry��ǌ}(�-��gY9�:�I�c�wY.�xڦF����� �*ˍ���(
#��it�!�8��W^�B�z�)��dp�Ԋo�$��|L��B��X�H>&m0�����X�C��a	e���׶�8�j�,�9�n�V��evoԝCg�}�m�$��ie7J[�S�]�Iu�\P�U2뢅��jX��s)t���D�fSf/^R�e��$KUB
�J*�E!o��W�,C���-u�Śt�Km��S��N�,;YōGQ��֪�NO�z�[�z=�л������q����&���J}�I�v�u݆2���|Jn$yD$ }�r���k�ś�]�ٹ�͆�R�cc9�}�+�!���g�K����rt�l��m:;6�XV*�vC�F�TT�tǛ�Z �-�bG&���)S��qr����[KS��v�}b{�$a@=��l8D�S�Բґ�:��7S��l(��:��\ݜ���d��'Q�qnHݲ)I���&"4�(k��H~�D�8Ӷ���ܻg��������<Âb��M`�0p��F���C�c�`�аr<2
Z��:WKƙ��x_��x��!����r6��`����< $��xWVq�c��x�W��mq�8��U^�W����-]-^*��YŪ���1U�W��8�/J�x^׊��qgq�q[^�v�s-����~+����)�~Z����*׬W�������/����Ǭ�g���mx�+�t�[W�W�z�\Z�Y�/�O9��Ի�c)x�d��FԽr��s;V�$�PK����Ã��KՏC�����uU��rÓ��JЗ����c�sQ̉�  �D=q�����Y�3�f��<?,@�h�/�>�.꫇>E3�˻�s�S=ܻ�.꫇w$����˺�ܒ���՗u\;�%���;�.��]�Uvӣ�׊±Zsꪥ ��JCw!0��)L�)7)1cO��.e̷C�Z�dy�;���1��la$!�I��%2�8\wf�������Q�>�5"Zi���B(E&R�''�VJ��Srt�;�VbP�MI1�Y=�J�jq�x����Gg���.���W�]=4����.�3d ���u绾�(���T�$�Zi���5g��v�oh3����D�D�BH�%#��_�J�N�]�@��=���'��F���n�)h&�9-4��q�U\x��N�O�+
�iۻ��]��Z�2B�=��]�b��gZU�p�3���H�i�^u3�c�u%:�4K�ln�u0퍖ƽf�&D��U*�:m�X�;V5�S��Kb�$�i�h�Ӏ9�&�
0L�f���Id�o�moi)��ӹ�A��� B�$�8�H�q����ξ�'7'2Y%�QY�9X�߬��Uca�M�P% ���9��@ąU��VI:��ك�FKM���ҫUzӣ�׊±U�2��h�X�b-�,��ʌ�2	��Ioi<`���M��y��Sn�>�T��G���9�9��Ox%eHQ�X��xN�J�)SV��}�q8���a`X�ª�,�@+�O�}|��l�܃� B^:b.$�lA��4��eJLҵ@TYU�p��ڕJ.iRPQ�*��S��wf2PA���捲����uR*"
SyQ���=M^�%*������mD`�w!P�^�J�"�n�t��S�H�V���D��F���>��|Ϫ��_^��?��c�lmq� H�f�e�}	�����m,��y�'&��U�SE��Ke�(����C��}4��Oaќ��ee˗��}G���uIҫǊ���;V��-�ڢ��.�����`�My�p���Ѥ�� t��RX�kuu�qY��6�,eTJ�&u�ܜd�$�}� �%�] ʵ�:{��
�G�!V��Jڏ�y�yO���������D��.;+�j��;6�X��=k����ut���1Wkm[�IE�nI�s����+����ٻ@��5j��q�V��l{��m��mM�=O �ZߛkI6X�2��cZB���nU\�=�<{���]`щ=�4>m-���Ӣ�0B,4@��rK�h(�t�UI��4U�w��='Ϝʉk̡��k�ů�wR0dv`n[S��M.ۜ��t{k���E�H��L���f�6��U5f�2�+ج4��6C��{3.�컳i��ZC	���z�C���$=$���%���@i�/�! ��WG.軨���%��3�S�~�2�\��h�r�Rf��m�q��y���2��M�a�4h�|ҫ��
�{>��5�5����w��]��ۭG0^�Ͼ���'8�t���o;R>Y��'�����=7I����TWg5\l؄*����8Cƛ_^�ƌM��m���R��� x��'})��ϟ*�|��Gg�Յb��G���j:؝6�Z(��\�I$%z���@x@��6PV�	%p�]�w2�w���ꪌ'M�"a��N�Z��I!��\��MP
MRƝ"p۱���$�@e)�	޿"����8mڰ�V�~��W�6����|*�T[�M]݁��uw�
�)�X�^\6�HK�����It>)AN ���e��㽸\���G���oOR�B��ڎ��g��m�﹌�/��xp~��ph�C��h�X%G��\z�8�X�~q������q>g������qzq�^.��3�p�����|�+��|�_2�/N3���\i��*�3�W�8֜gK���g�U��̿2Uڪ��gm��*��]�c'����e�x�����i�W��\^��4�{��q\o-ⸯ[�{\9���՜��-^-^)���U|�߲گ�_e�4ϕ�zW�����8�.��巍��W�e��.��Ux�y-�-^�8p#�����D!bp��a�=�x���,�0%f�x�H� �yV/�TO�scr̒��R�!ؕݼ�!>��67��u����[E�Q����7�a�l�@�F�&�A7Y�����a���T	��5�^w��a̫3��`��j� �Ȩ��̄���}YwUû�Z{����w$��wGue�W�Ii����˻�ܒ�����Yw\;�#�������	�c���j±]|��i�+%��h�1i3L0����%��ٍ`Rm�*��V&K��2��RGQѦі�Z55\2ؚ'=x�6�lF���`%�`,ݖFX&��鶻�X�népG��0��z�ÆkLu/Ktu�ͦ�M
��F�m!�5�VSA�p3Y5���e�l]bmsan���2ᙹ�2�k�k��ͨ]6�����$�̽���6чcb\r3rk���pk�rC�,��`�P�1٤Ͱh�.�0�Kf�e�cPˡon���Yx��G�u4wԝ,��yR
msl�ٍ���˫���K	e�T��eH�ŕ%Ҧ�P��cU:�ͣi���3Y��kY�e f^	��� )o�Im�j����H��q�f@�D3F�NT����m�"h���r8�	WLz�W3��S����3��u�W[�#�X���~y�.3��>n}m�q����|�lc�|z�X��Z�z�B����*,R��:�:��Q�Sm6^�À���!,��>8x=e�{@z�p�@��)�^���,�	��7�w-R��wU6�y�r��Ko�	�GF);}?O�;v�1Ə���,�`4� ���H��"��#�\��:G'RtÑ��a8a7���eZ�7�$j���Z.Ni�a��ppti�c��00Ǯ6�$2<�獘M7�I����T�HHi�N,yt�t�1��zx�1�I"�I��	⦳��:�T���0^L������=  �{�������w�k��bI�(��Ҥ�˴�t3ddل������e����p�O[e�m4gf���f�>���W�u���ch��P@ �)�"����آ�H��H�����×����c�6��WV����Ȓk�+��y�Q�m�5�&��v���4�me�n�۫I������j1!-����X��e��W�ܧ$Kq�e*�e0��{�ՆD�Rzu:�|2L��e<:�6L��-��
ϒN'��7ǼD�@�縒�}��p�WRf�fY�Z�nOOݽ���g����1�Z<<v��o{̶ׁ��� e0��~���a@l��w�j~���}�q�^�k-�t��k)����$q��N�{;����넣��yi���4zrB��#T���WS�ʪ���������]��V���n���uj�L�S%�M����d#�Xm;I'Y�}�q'�L;�R��,@��
�XX��Uw8�g���y'�sf��=^���<}0�1d!	�3�R�P$!iD_�o帕IU�����ָl�:o��Ʋ�2�H��vY�����6�������l1���8j}��Β���nr�]k1�˪n��r���*�&����t.�BD�I��Y���o���M&Ҍv�z�!�w O��R�6�;!^vgN�Ux�������c�	1VZ�+�[#6*j���A��|��3�$�y q�W����D�+���B�̴ldb@��Ub��B��8׬eo7����%�	-kD/Ul�,�W1m6��A��g�$����p�OgL�������y��b��05f=M: D�lua��Q�9!�&�|��`
�F{,�Y�S��nFNs�����l���A\q�+a�������/�kh���ԆC�G	$# X^����J�����'�ͼK���H��6�O<8��6^}�(���.�)���c��D�l� ~�0ZzCn:���������ݶ�ã��~��8���l��7����q�������z|�]��{���|�������6�|�\g�ǙoN1����L��xW����<_�Ϝ��>�p��>���XO��>�`KūǪ�N/M8֗����ʫ�W���UV֫kU�խ�WkU�̫?-��j�Ux��g��t�Yیq}q�/�ی�W�����[W��1ūūūŏV�1��o�WՕ}]/�3�/K�_���_[c���;]��q|\|歪���j��x�x��1����v%1�"��:��TP�2�R�^(CpVV��'׸$a��f��媌�{"|��I+L@*f�Uk���6�Ȯ��K(���Ah�Dw\R�Q����ӈ���窲�wGwwOUe�p�<��˺��y=��=U�uø�����UYw|;�,]���UYwb�x�U�➞;a�5�{;�~�����h^
�Y�T�O��a��)�r2~r���+��T�	�O9 �)�vZw��a�1٢��BӶKZ(���&B9;��.�.�!��T���b��j��-�z4��{;�#��u�-��~e�#��lzz�8t2�тBzGԱ+}|L��4�8KO:�z��NM�!>��"]���&	��x�]&L'��V>Uvz����cow�u��Uע�$[�iUV
��^��%i_���]!6s,7i�4
�i���B�jCA��R���܋�GbP�)M���m�MX�f���3j�+ڄy���,�X�t�:�����&��01�hֈI$�a�C���KB����x2px��HH�!Jix�Jk}%Y��U�V 1Bm�Y��bI���<6�ӵW��xx�1�w���:��m0s��r�{�8J02GG����P8b6`��(^+Uw`��6D�"jP�K���6!i��� @����mP Uզ�#�p8�Y(ueY�)
Л�
x����u'>��UUj:�Q��ϖ0��U~��;Uv�U��<v�f�z�f@2�pm6��|`��W|0y3r���<���ds�I��9��ږ+�\�uֵ����r�<�_<���ic���0�5'���@H~��O��ر�k��U^4��ڞ)]�e�\ʮø������s�$�4���u<�T��mUeeBQC�@���Q������Ҳ�փ�	�'�	�Ņ� �=��nב�G<�����6񧪯�ʯ��{@�@"��\�6bd+�sw(əG���{��w�����e�O`N׮�dtC,�
�QҼU�ۈB����=tji41��iQ�43��f�lhK"�ǍZ��[jWʇ�
��Kk�.%�eu�����Kä���A�kY�V�
 �qw�F5`�K��Qd�}ھpu����T�dm���UP�E�N�\��;\<��!�%Wn�6x�v��V�u���<vi�ha���5���H4�M��O �PB�j�Ux��\koI\��U^�a�u��"�b*�lIo������X�!K��Q����ʮ;�)]���zf�cYo���܋^�5�`<{�� n��JLɳd'@/�=�B�*�  c8M=t}KyEU*a2��Xh�u;�!�f�$��a���ͦ�ڮ�[~U|���J��߭����w���d�}���$�[Ji�]e�Jmi,,"=���#;�{�a&��	)������n5ĵJ���
#����MkhZ`����/�� )4��=���3`N�
�ı�X�ԍ�ힸ����2ݾgϙ��m�Vק���<^=�x��_����k��x͸�׍������[ӌ�\].�t�8ʼ/W��|i�/���5�y���:^.��1�2�ūÌ��Z^1�^)�j�ګܶ���ⶵf��U�*�t�O�t���x��1W�8�q\_�����N/�1�q�6�Y����9����ӌ�����x�����̷ն��_Vz̽?4��������8��c����M������s-�Ůe4	A�H<�8X�J�y�
�W=n�M.R/Z�}�R�b��N*��j��*W��b $�S
6��^b��VK�����5me���y�w�cLsR�ȕd�Ы�a^H݊�qء��MZ�CXZ�$��Sx͍*a��A BP��3��U MTΑ`Jh#iL-fW�q�ꪬ���yZ��˵ø�����UU�|;��=��33uÇq=g���fn��q=g���fn��+Ǌ��O������WW1���q�B�������m�`��T����bJ��ͳP$�cuրL���n[>�޶��
���-;C0,�U��Ш�sIsnfe��e�"�b��'���+ָ��R�{-�	t.�R�0k{\S����tŰf��*��)͍���[`恶qS;���j�{v�Ld�-��RC[0��`n�6�jg��^�֕���l�-ؗK 3�4�P��T��K645�.���4$6�4�͡	�ke�t֮�<]M���ؙ�;0�m��[rd��$t��:��K�V�X�]�D�t�q�7F�e��F�W}�'�_q=aŌ�:�kڤ3֔p����M���sŬl%ՎAt�aX��MI]��Ci��V��eiN�k3UWW�8��=F�z�q�[zh5�]d�M���&�'�<�ԒT�`D����L�X����B�j�4�u��v)syt�ie�~w������v�}�銯^*�v=<R�~���C@�'����x�������&�a'q�4=JKs$��D�t��P�//;UyNj)Z2��d�ֶU��B�&��ҹg�C^Os����-�Ƙ�)ϲI�q��WOU^;�)]�}�֬����1&�:BHL��i�^  1�^X�t��p>E��KE60cd,�Ex�@���2~v�<Ԯ�ѕ��$|��nOM��Q���b�#�[i��r>����8���W�c��Wn���X�Lx��s�?Z��R�ב�[�bAD�IG � ��S�!����	��|�X+�pߒ����Y��^�!7�:�8�ޞ�Bi�d����1䁖v�o�ggΟ1�|�zx�v��Y��]��#m���J�]�|�,����)av�,`���-�ν��R�nRc��	k ن��ioj��h�e�R6��b3�B$��F��AJ7�����<זRp�zI2J%&�ZY��۫�E]U˲���iC�Ԣ�2�a��u3�������E��]�);m3Ex֙��i�}��)��sv�������ɓl���t�[Vʺ��1�1����燷s���mB�m8��2kd��=Jrp���2I#4x�Z��kM�@ֺ��m�řy�K��B" ��j)�K����Zf�>;(��=��h�a$�a0�)����1�����~�s�e�&><geQEh�Y�ۄ�R���2]�{Z^V1o�ګ���PR�R
����X1X�9��s��Χ�I!ǩ��)N��$�i��I7�))"$ 6�K'�4%��e����e�\�fZ.�(W��H2,���T\�kJ�h-�R�˙4��!3Rf,�J,�
���Sww��6k�*�cI����R�Y&6��a��-�V+i\�ɸ���읪�r���"�ܔ�j��	��n�ћ��v�*�lډ�/4새��T��9�w6�J*�D�\��n\�J2��pM���ƪA����uV�Z���:��D�$Ĥ�ޑ;��LtN	1%:S�$��"xj��Zk3e:u#�'K������|¾��^����5���C;!Cڑbݯ!v��b�JbVZ����S.6iɔ�qL�&�x'�;cLc<)Z��C��$w`�%���2�Il@b.n�
�6.��t����%,���6FA�XAYIS'v��e�u���=��vv��UII���G|a!g;sLv�Og��OS�qM�4-�[�c�%�-����$�����E���L�㔮�m6d���]Ѳׄ�V�9&���ZYV&�x�[@��m[s*s.�t%�E��B[rF�bQ�dcm�ur#F�1�D*��$�	W	�ݻJ6��OZ��k��UT��`�� �W�  -�4� ����B�R����ӎ9ϧ�Om�%�K��XK�M���gfW9n��(�El�!�3��2.&��!&J��UGKL8Hu0��ZD�g$&�a�'R���)��˹d���D�j4Ӕ���E�KL��0�0��YgN<m㏞�z�o��O���x���|�O�|���<z�m6�lVͺV͛+Ǎ;m���<Wm6�lV͛6l�m��m����_�V���p�p����=6��mv��ͼV��f�6l�������q�n�qێ=�v����i�6m�M�m������	.NS��X7����	p���(������<� 55�Z��n�$ȓ�[��px; ��OCid��h
45CZZ�C�P�TjQ�TG0�%E.,��(������P��%ډA��K��XՉ8?vJ�$j��]n�7���+�ݍ(?#P.;�uD��:�#�7P�؛*'�X'�%$Z���Ws:�*Y�h�&?���ff��q=G���ff��q=G���ff��q=G���ff��q=G���ff��q=G���ff���a&<x=<R��'Lukvڝd�<�ǩǮ����TQG��Y�`��]ELכ�#e��,@�{�<�Y*�iv�K�_a-3��!��e�V[Rj 8�J�8������:v<<R������5��~q�nXE��N2{7%�|��yZ[E�j`{U�u;ȒN�u�k��JJL�be�K<r��x�|�]��7�V�ɓ2��ϧ�\c�1�;'rs	wݷ���4-8��r���'1� 饕�#EJ\X��3v�j&��Uu�]46J,L%�c�.�"Y��j+I�&�����R�.,�nQ[6�տ@ \jU. ����@
m�Z`�8vq:���i���u<�	�!9�3W][��7u�D�L�M������z튭1��ޏ�!�n>B��14D�GS.����:\@ŷ|�Jԭ̠����}��)z��<�¸�pUH�ҋO��mk��<{q;�)Lk�We
�E#x$$�k���|Y��� T�y #�m��;��mkڹG��c����J�י��Y��'Qg�Ӽ�9�	�޻��Z���D��݊B�U�f�.N����APW� 5/�i�{� ^kn�Z�hLx�W�x�1����J�'?s|s�����Q����.�m��� 2
!��-H�,��D�'Y8�hq�'�.軻ӷ>��r%�Lu��Pa;��q�N��Q��ʫ6�2�N9|Nۓi��i�FHCEE\X��ZBC��͚���X`�&��	��Ƽ�Ć����&����msj]3�1L�V��ݣ�u����[�MN��j�<M�x&��va��d5ne� O؟�td�r`��է#G�Ӹ�'-.O#���=��m˶�؞1`M�=��M3��'/���2�-#D`X�\�9�>�&MOӎ�^1����W�YA�03,�r˰)���TY��dqu��� F� .wkF�Ƿk��Bƨ6����X�,Z�JrUATQ�THT�Kt���6����H'��.�J����~m=Ux�_�PѴ��7�BJ���i�)�P�Ie�j5�U�cQ����_	��P�R�4֣��,kʗ� D$��Bm'��e��2���Rq3ܯ�BI��g��Um��<v�*�R���p-��Y�b	C���#´jϞ-��z�f�۰�h:I�t��2ۤ%�H[V���ju��=�$��ǭ��n�9���E�����~q�oϞ6�맮6��<t�"�1���Ɔ41�C0H��6�lV͛6�[W�x�׍�|�Zm��[6lٹ��m6m��p��������8p鳎q\m��+�q�m����Sf͛t����;x�8�����O\m�o��Ҷ�[0�m�mӫ���.�M�E�P�r$������,uD֭�;��K��
��(��L��g$�d�%�c�7��]]�°MQ���72�
"�@���õc6#H�y9��Z��.�=tx4�k��)I�bX�DL��P���~2I�;��337���OQ��陙��;��=��33=�;��=��33=�;��=��33=�;���9κ뮴�U�1�t�<Ux����8��6�Q|��-X�`$u)szX��3�x��]H���F���њ�L�H�bےǴ���k4UYtuk����?�4	�V�� �}nͦ�k�X[�"��tbaƖ�7h�D#*4tZ��b��0��ⶠ�r�``��r�h�i�s-m�i�,C�d3�ب�Mnv���ơ�l%�����.�iM�T��%Yr��4l�R.eM�m���eк�e�adԷ]�˥�2ʒ̛\]�T����.�/C��js���b���n�р$��pi��3-:+̳Y�v��Y�`�Fi��\u��fs�%�ru;|���ދ��MIw`���%5�ؖ� �XF�e�M�0��CJ���(�k-�Q�Gck5��jL�34ݭ����a&�����h]��U�1*bTe>�si��4�]���ӒȘ;��TT���٧Éi�$��i8�#�����SI��磜@����4�̘�1ٌ� 42��.5Mb�|R%R��!R���:|�Ux�{������Y�t����y��NS��Hx�+���VY���=��}�=ө�KH��T��*�c0�������Ɠ��u����am��^t�ך�_`IymU�z�1���U��N��X�@,�����G�� ��Z^|�&4*��O���)%GN�ƶ΢�ی�:��y][�d~r5��~-�Vw>�F��#����j���c��Ҽa[��m�od�z�5Nj}�����H�l�9��l�s۾N9Ǐ9nb����U���f2�c����P�- ��N�nK��{МW� lk|h~V$������ֽ��i�V+�V���kIiB҉��:*�ՙrf�,�e�{��N<|�P�?%6V3u�붕Xe:if�.���-��k5�1&Yj�e�i�B(I�R(��^t��$���u5�I!��l�����r�}�82S����&1�� Zkꮵ���n]te!��:jb�%�-����;�%����w�&��(�.�t�1�f�^1�9j��[us;�{�xa(�ᦓ��UTB�::�6y'9��d�ru:ڪ������)R������׏'>�K�ON2�ff���+��N�_mZ��ڪ�cLc>>Ux��ۓ<���6KH����(�%cޙ#��(u�X0
\g̞C�=1$'�r�I$�Q�<N�/q�jY^�����H�Lsn]o�oz�^7�M���;�ڦ��[k����%$2��=�'�Q����c�g�CEG�j����	���yK6�������?b�71�m�
vtn�!��d����x�Nk\�I	��%�M&�w*/��%� :�ע�c \h��c�v�{�G��U]1��co�P��23����o+���̙��8:b�<D�^q,Jk�iK+�`dЅ.k���e�#\��wf���E�v��d�,����if��-�WbV���Ac6u�N��~c�����J�u颓If�t�HB�BI&�j�`�h��⩢�OKH�ė�;�s����!�̰�GŠ�K�eumRˬ_f{G��^����0��y��.���ד�]:j���$v�<�QxOB�m��cti�ڦ�=ح�EL}ƹ��q�"rA �$Hp�I��j��W��u,�m|t82HI4�',ѳGOL�q��=m�ͱ㶝6�o6���m�o�|�׍�m�F�m�ٳfͫ��<m��ݽv�Vح�6l�j�m6ڶۆ�>Wf4�o�շ�v�c���z�m�z����ÇN8�O����qێ��q^���޻m�l���6����u�F�z���Z� D�X�"��ҽw��zq��]�է���A���t6��IY6����d�DD�@�7˶Ȧj6 ���,�Y�+�F����ff{9<;��ff{9<;��ff{9<;��ff{9<;��ff{9<;��ff`H �HA`�h4PPQ��3 �x��ΰQ�m���x�S��zS^3i����w��,C^ef�!�n��;����cn�Q�}����ɝ�O)�g�B�ܸ��{�⪴��1��<<`PQ�a�p��Cf��=Mi��I#��2˕�X@m��O0!��:�	7&�X��v���A$R)�Ѯ�j1{�w:_ki���˛�Bd٢�G
(BƁ�X@ �:`,�7!RPSCP*L%����r�����j�T���Y�YNm�;k��'[R�D�J+n��Y�e��\]�-��Y6�K���`a
5�[ջE���m7k4z|�� �8�eF����D�AM����6�nf��uU���ݍO~U���X�{jZ���؂wU���Q A����qgӓ#�>b��;c����c\��evN��ֺ���}l�I[q����l�hyϻ(ܽҶ�S��O����0��#�D![�km��Ɗ��lp#YH��[X�a�g��v��e>��nI@˲�:��i0��K�{9+xҫ�<c���ƨ��J�VˆA�r����.G'3:80�k��)6�8Cv^xߍ���Q�k$!	�&ܙN�M&�I�U�ft\i}=�u0񪭱�Ǉgl0Ǽ{��w�]��5j���ĴýW�����?NQ�KP��e����3�1�޽>ef�Xt�䎒<0\�(�5�w}O2u�[ɴ�4O{�n�2B(�Eh� �B��Y�����U!U��ț0��(�L����<��Fœ"H��=.��m�E�M�Wit�Yx��4�й6�Z�0l���J�cM.v�^��hA�1X�r;@�m�Ӗ?$��}w�^���5�Kr�!$B{X
k\F߷���iv�Z���m|h@
�
�&�D6�KH���ν*�h�WUQH�����`���e��q+I�.�B;c�1�����ϵ��k3O	��0��O�^��f�y��4{8��y$<���K���'Y<�<�im��������Ƽ���ҋ�=P�1�T.5�u-9���0��n��6Q�E1���1mݙK4N�9�}isL���A���w�mKk�r#�)�vK�(T�V��YQU�������������5�o�-ݧG�r"a!��K\h�Wl|�1���1���u��s%]�$��<V�>�溪�}�*�1r��eˢ�����X�'��<x��V�����Q�Q��197�l�fn$�Ҷ���g������}� �B$�T�I$�@b*�%��_�~����O�{���$!� ����!D@$29���7���l��B���}A��R}�bIH��"R(��R*E"�T�J�ȕ%H�)%�*K"RX(�RQD���T��Q`��E�(�Y"�!E"�EH�Z�5"Q`��QR(�XJ(�Y%%%�T�H��Qa(�X���E"�!EH��F)�E"��E�!E�(�Qb(�E�Q�a��$QR(�Qd(�QR(�Y�!a�#(�Qd(�(�QR(�Y
,%�X.R4EB�"Qb(�EB�"Qd(�T��������L"�
*E
,IE���>t����TuH�EB��E���EH��Qb(�%B�*F$�Y
*EIEH�����P�ȣ��,QJ,QH��(�QR(�J*%�d��%
*E
)Y%�*(�RJ�����"�B�E"�T�*E$�X�)RQD��(�T�T(���
*J*EIE��*EB�%$�QIE���QR(�Q(�QD��$��P��E�(�TJ,�"��E���
(QD��QH��QR(�J)(�1�Q(�EH��XX�*%%JIb(�T(�IEB���T�`ɘI�,P��(�i%�P�B�,R�b�K��X�Z����K*),�--�e(�-(�,P������2��Q)E���P�D����b�R��%�����)%�,Qiib�I,Qb�Z,Q-%�,Qb�)h,Qi,�,���Qb�RK(�Ie,Qe&)�K(�E�YD��(�E�X��(��(��J�QeQb�)%�,��U(��S&RX���(�(�E�X����X��,Qe%�%�YE�X��Ib��),�h,Qe)*Qe�X��X���YR�J*�D��R�X�{���R�K��)e,�(�)e,R��e,�,��%���U�YJ�K)RQ"�D�Y
E�R,�"�T(�%
��%"�Qs�R,E"�R,%"�R))�B���Ed�E�H��"�d��"�aH�H�H���#��Tr���O�	Bh�;�'�}�T	P�a$S3�J���?��������^O�}i���C��x�������w�+���_���p�e���Ҍ�?.|t�$�/���M������s�!!��|��,�߽?��O����>?Gϸ{��G�EU����������փ��?`���/�0EU��VP?�h��s���'��B�Hh�1(S���d�C���|�=?��d>���? �?�EU}�T�S����,$���-ۚP�V���#���'ښ���RRRo��(�@�٭o����������_���b���w�����#z)���|h�l@�TU[,(Q�b
+p�*� ���B�X~qZ�7�A*鿿�?6�C��c��I����(�FAh�B��KER�eD�%��BDK���M������hN?�k������C�@�@<]�����R�?��˚~����("��%��hQ-~/�_Ͻ�p��㯟�?#�~�ϫ_�Rd� ����c������&G�����0?G�_'���埬�����EU���`u��Y�����?!ޛ:\2?�~C��'���UQ>���~����,����Xek�8M��IᴛH	F��C��TP�Z���?`�$���G�-�(�
P�����e�C���;����C�R��l�LO3G�����.SN����� )\�__�!$���?G�3��_1TO���C�I���~B��ň}�����������gҟʓ����]��c�	��O�~���g��H���?)�@�h�!<L"��|��ϋ�����UQ8��}�6~���w�'��'�����~ |���t�2~���L,�hg��7_t�����O�> ���ǺϿi��ἃ�����DUQ4��O�~C�т�Ʃ>���?!�� Ǣ|�~��?���x���$S�@���͙
P:�'��?:q����C�O� AA@)�{�>��>���ݡ�}?���}���y���Ժ?�6R|�rO��
�d?:U Z@b'}M����.�p� ���