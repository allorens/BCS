BZh91AY&SYՕ]Jt#߀py����߰����`�^�     B�ET  @Gk0��       �
 � �d +���     c�ف }8� ������֪�ck��1��5E���Q���۶m����p�s��72����^�8�F����v�/ZU��{�C��{δ:{{�U�=�q��7kp�c#�   �,�#��l�f^�ǻ��wތOc$�݆�u@��9��
��q����]�iݕ��n���aϼ7���ve��� �   Y�[�����x=�ީ�{b�cv܇a���V�=B<{�ͨ6q��O;wv�j�6��;����������  �sηn�ٶk��n�v�\��rwk��c�:��·�/��+٨o��ξ�u�z=�#�����^�a��o�/   �z����n���ֻc�V�nwX����ɣn�o��^P�n|�A���ZuM}��=�9��uM�wn���Ԁ      P%
*Q"�TJ��      *��i��J��� �` Ci�5?B"IU  &   LL )�$�Pр&i�FL0&��MDU$�I��F Ih�&!15=2eOSd�mSe�&� U5$��U*0�M4�ɀ&ѓ���a;%N�!U	�ǁ�� w���*7 Q�Q���8�
!�\��Q���W�7�����?�wB*�TU�Q ����	RI?6�;�?B	�I?��� �	�CQ��|�=�z�z{����pg�Q��Ϭ��s~M;�G���&	N��;����_5 �5�4qC��U'4h�jJٺ4܂o�rq1�:��I߹�%�\)Ԃc$Ć2LNS'4'4���J��9�����ޡ�0Xǫ��t:m�ΚtK(�nO�h4���C�ϡ8M�h��4ɡ5��ԇ���옒���O���q4�i!ߓ���D�lMv2P��D�"w�&	��?"N��t�'XN��Ɍ'L�:�,w�pp���0�$rG�S��Z �����4S�}��DN�"`�	B_Rt��d�� �%4DDL�B����L�D��:N��e�'��DI��D�N�$�M��H��DzYA�D�"=8P��-�'S
/���tO�"D��:KI�'��
a>Bp7I9ĉ������s:Nc�|��,�ZH�\H���h�4W�DN"#߰��hX��H�9�P�����N?"D�u'�r�f��'���l���""f��$��:C>��}�b"�O��l�'�	��>٭�M�D��'G�#d�t_D�(m���g�m�H�N�	,�R'�N��:u0�H?\�(G��L�3R�LN�e�p��Hi�rr����b;�1�)����7ʉ���o�1���0��0�2�!L�~�϶#Q�'Y�֦�s�no@�؋!�!߳��N�p~d���h�Z��nU�e��bbe�9���-+V&#vW�dџQ�H���#�+��RL���2�h�Z��yu��pཀྵ�މ~�K4���{�~���R�%�f�p��L�O����Rpk�pG�S�Ƣj�4a���W/ir�hy>��a�8X��Y�p֢#�DE�f���N �e�d6#9Qfi�AU�DE�K�S�Ѝ�DG�Q:2'ML �|����7���)��N�P���Dl�8VH#*�"gM-J����ȋ ��L+c"av��I��d��	������r�a��(Nq�d�/�d62�":ʈ��R�?H�QŐNN�������R"p�]DG9QcԳF��D�ȉb������C�bp���]���7r?H�QŐNN��������h�4Q$��Q�Ș,Nd�&���/�/�F �w�}\4^�%ѽ<�`䣴!L�|p>G��t�]�v����!ϡeH�͈�*=¸"��lJ����B9���eD~�jt�D�v��;�}��I�J8�GC�gN�圳��hSJ��ub'�=�!l�aL���969u3\"?t�$��85���1�Ʀ	�58j�pދ�R'rX����a��*�}�<�9>E�RX����sH٢�b��f��M3�gx��^�ԭ9W������w��/���>l�k3	%�qު;�L�G;Q�Vbt�%*5C��b�q�n���uy|�O�6VI�B�#	H<�r`�X�'w*r5.��&�q��u,᜜+R�Ԕ�Q��J�ÛJ�Q�6&{S��L���*�iia�9�5�O�`�t3�}f��rs&cP�{>���*�	}������wO�t��V|���{�D�jeMP����/�|j>�}��c����F}��mf/���}�ϙ�K����]��������PX���*����_t�Mϙ��d�����LS~O�����.�*z��[>�Ϭg�>�T����-����a���×k�nd���T�ȉ��; �Ӳ%�ѽ�D�hJ��fɅ�W�%�9���I9���}8C�'H:j����"�ؔF����R"'/�6;ܭ�n$����,Ly)::쯟��f�SPD�$D��6A�Dy-ep4c�KjW��%~�Ѩ���D~�5�JDy쯟��lM;���r�r�h��H��	�2�я�:&vY���Q�&��#�(N��%7)��MT�9����M�bhy4=�����q�"'g
:������ʳF��V	���:�RhM}�Q��'�D�pK�dD�jU���DЊaFƉ��"P����t~Nrlr|�"wU+D��rY";�E����l��mD�UKr�����a�z�2N�U��q8%�&��a/��&Ʀ�H�Sf�����eh�p6HjJ�<2�uku�-j��Mv���K���gD�Y\5������9٭Τ����y8�b?a�5�c��-�V	��t���M&j�:=�a�A�d+q��r#S���j��Uc �%��Ʌ�`����N��9����9�̓S3��%w&k"d9�g�_��pK�r	�N���G�;Q��x�Zߴ��-����zl޺����+�V�d����qp�e��~���ݫ�P�!�K���N���g���� ai�ý>����2��&=����9�78T����ly>[�7�7��Ʈ�����1�tj�ڞ��z���o�wإ��ۙ�\c���7rW<��&�f�'rD�,�$�buzI�I�Y�&\ΚvN�q�6o�[�sBc�sF�-�7�3� ��a,�+aZ*$8%&ZN�ޤ��O	���zN��u�<(�>2�1��gf�@�92-E$%~�堅�Aڨl�������J�9�j��gfBG�� ț���-�+���h��7[5��K®k\{�5��vO�u����^�]�Y(t��	�v"N�3(/Ou�!E���va���˵3`��{��]6}g{�+��v�dh��)�7���v��żwo�M���}�ާ��~Zs~�o&rv�3��N}�)� ߺ��~ݛߑ;辺w;���۴Лp�]����G�����G�wN�-������zn�ϯ��'J��|�6_gn��w��]ȩn�����=���٦������f�vN�s���ܚ�O]t��ϻ�3���{�{5u�wWa��f�����WͭN߳U�of,���>��=Z��vt���7gOg��5~[����J�d���٦���a�=�w�{�������߹��j��<ƿ0ɯ(��_��OOߟ���'�*���W�ߺK�ܧ{fO^�¥Y ��㰆U�xo���w_ԛ����t��X?>��9��������z��w�>kǰ��a���\�]ʷ(���5}���:w�ٓ^ώߧH�����^�{�-��)�fU��83~���|�y,���F���v�����>���w�7�+��h�;7��]؟���������E}�M5i�b�s�}�!=ܿ��{>�����;�v-�wp?W$pƞ��x컆��n�����z���g�wnsux�Mn]�7{����T��2�1����a���{�易�u�7v�f٥ǐ��a�pm5�湼7/�g��z����3�v�0d�՗>]�t<�u�pa��8��W�e ���c�_�.�/})��g���z�����4����쳿PZ��v&Ȝ���[v���_L��zS},��iM ����N��e�} t擤�M�S�0f`/��{�t2I"a�����L(����` ,��� 9ހ}(~���7��t������S�};���/^��5��ͿNT�����D��~����;�)`�j��S3�½~>��s�-1vm�)J�s�M��X�߮m3t�)���>Ve�gm��ģ��5�uX7�`���ֳ�dlL�I�$:�6x]Õd%����;�Gw3g��6i�T����tz->=��v�P]i��}�q�e��g�`�2�q�r��n�Ym�^��d�G�dMf�U��,��>騊ů%>��D���c���?٫;n.\��?M�v��L��]���"����o�{�{�Gd����[�<�_5B�9}�w-�VK�xv��b�ߍQc�^�v����~.1g����q���o�b����~�ǽ?c>=�>�|g��>�L~y��?7�ǝ�٪��n��y_`�)��p7
�nV���5���3��H(ؾ�]�>�b�|<�}�����ݼ���d����÷&lY�݁>�SC;W�}�o��W~��~�o�"{�0^~������Ͼ����^�<9�3��G��_������'�F��{�W[M�/|�BE��G�߶���ޒw>�n���5�o7̮y����y�W7U�L�����y�Ѫ�w\�����^̌,�n�)��j�W�o5Ǚ�v�W��W�}��Z��6|����Q�U��w�g��f��$�{=7����+i�q?nߏ��w=�����}�~3uN��v��o�����ﯺu?5�{���u�k&�ِ�)���{,�m!�8���~�9��{>� �μ���Z���={�v�wO�̚:���l�������WY��V���b����u��8�oN�+T�+�7���ɭ�3��_���&K�;��P_{.��ھ��ٛ��s='~�������w˳�����f{SmZǤ���!�BG?K^�!=�7���Q�o���5��w�=��2�5K�$!18���ڳ8�W����d&��OeQ?w3��0�I�v�ros}�{�����Nu�>��ݲO��5�����t=�wyr@�!�ȳ��'�/��7ֹ�3'f��]�g1��7��S�O�����N����$��y��`Jd��?c�×=<��^�v{p���ø0�/��ȻF�d~vq����M[���t��o׷2W����`�Y�I;1���������L�[w��t�M�ck�����>̚�؛�._?�����N��Z%�L6a���Y�N�˿���C���t���_۹��;�{�`ng�\��!7��/^j�W�ٍϵ��vt�,��ٳ������G�,�3غ~�w�g�vc���&�r��NO�N�S)��!��S��g�ﱌ<B���S
����Uy��̞|�z�l����)��/F|K����w�ߍ}~T�z}��~��U�\}��݃��ҵ�g����}Ґˏ����������U@�I���r@����y��,%�>����)N?f�Oޫ�5g5�gc����k����m���e��c�m��x�ٝ�:�e��I�^-�#�zگr�{���5���{W�������@�a���>����OE����_k�����3�i��f��:�ٱU�'a^fe�f�1�<i�3&,�L��Y�7&a�y&��[�5�s#�nw�W��Ӝι���ᾚ�yy���5�׵�u�Nq������������x���M{��r��3zu3�M������k�c>�?�R�ǳ=gb�?
'$|êQW�}w��r�2��,���{|o�>ٚ�j���LϷ����|�k��oV�ϱ�����տY�w2L��[$�5igVi��5闥U������t�S�T�Ğ6�؛��"l�w%ӽ�����w&v\����}����tr9���w~�rl���uI3~��l0c��y7w��S���sv�FgpgG�I�};�J������{��=��^�wp���Dd�ݘU2�d�g�����^٣\���r�ל�������`B{�f�gvΕ�����$߿�����}D��=p���!!~����קI���|�2�C�������Ic���&h��'�����s����7�2K���J�r�$$�8E�%j� ��R�\U[muZEk���'���:�d�|d�r�Q�"�[P�)#�`Z�\���"�1�D�P+?�n\�n�X�4U��YJ��e��E#�j�R���u60-��E�F�\cyr��M�n���7*������ �\����Sx�hҲ^0e�kM88�m�EZ���v�!��k�U28�u쑺a]��U�Î�eʁ�d� ����Yxr�7m��X�W��\�Ij�ɘ��5b��
^8��Ϧ_F���11�8+�Q����o cj����1I8LřSj86\N"Y}��X��v�Vj%ctU�C�F�pB��j��+M�gM�a�
��mcPr��C�Q!��\��d��G���un�Q�겡`�hª�
�v��(܈"'�C���&슎ES�ڶ����Q� ���d~9�Q�j�:�"i��iTRH2Q�_l���&���V����"'
�pj!ZQ[���EZ����)
	"mV�*`�
r�mBrGB:A����]g!h�m��\�!c,u�ꃔ��+C	_-�dP�!q7(��B�u�eC��u��(rP��������̫Ԉ��!%���UQl�(ر�4T�Z&J����f�#i���s{:Z�vK$d,��,{նm�*Z�{���=<8�
@P�,���}��x��l�J��
�:��X��p�V��o,�	9j����M��m�)J��m�q��YS��NI,Rr�I����p���֪=U[�"v�V�e�ӳʼ*�Ƅ�E|~���]:1�C�G�Ñ���먰v86���9S�R�C'k4�@�\P�r�����1ŜaP���R�RϚ�Ybj<�)g�UX�v���[�dE�W��a|�\h�|�<���/�7�m���U�l�UJ9��_���Q�L�R��b�3��="zԖEZ�5E�Gv�nz��cd��yW�m�8�J�&��q�tO�ǌ�2x�V"�8zK5K���=���B�z�s�T�u@W��5	n�:�^�?���7�T��z�0���]g�~}�h�B2 ��D$�"Bt�w��߾MkZҪ���������X���J��X���������X�����lWJ�j�UҪ�ZUW+�kJ�������UW�Ҫ��UW�Uz�{����;׵Qd��(!L�"j
2*�H*(@��! �"ȡ �H�"j*�:��W�Ҫ��*�1b���*��*���U^�UU�*��*��*��b��-*��*�UmWN��*�U^�J�⫵V�]����U⫵V�]���Gā��$��@$Q�T����A-$T�����AVDY�����U�]��UmUګj��[V�U�sK�\UҪ�WJ��]*�t��V�U�UUTUUz�Ux��]�v�Uګj�j�UUťU\ZUW��UW�U�Y�� �|$IH�H$�bUfffg2e�����UqiUW�U�U[Uڪڮ�U�U[U��*�]*��t��U�iU\X���UUTUw��Ҫ�-*��b�����������������ާY���A`B
HIc$�L ���RA@��и��jHjV�AIT�	@G��u����QTI���w�V�����@�gy�x�<L��G��N��:&	���"%�A	B&�D�	�0KgM��Bh�	BP��b'D�(A(DK�tD�bY�4i�6P��?2|� �!�Ad��:X�pN%�١4C��aDD����DJ�L:"tL,K6QЂ �	�4&��B%��>㙭���}L8�K
�r'��!?�-pyJ��ƈ�S����֦9%u 4�N	��yu�bN;"���k��Z(��(�XO��X�H&���J��u��P`�����h�Lt��yq�88�&r�MJ�%E��B4�"c_Lbx0�VJ�� r��q�VӍT�]�d�֐�u>4U��ձ�Fq��´�h��O��<��W"$��NV�A� 2E��]��m�6�
d�`%�G���$$D�RB��n~��O��g$�<�)0�b�>�1�ƈWe�%b���ȸ�#%�Q��RV��WÀجV��HAHct��ȓ�T˄E�ӗ2�,-LLH����#s�h��S7�>Ƈ��G6$&(��&K����h��$uRH�T�L	U�rTjI�ly���%nءYK�Lr��Xe�)d��,��T��H7Z4K�mi�԰Q؀h�J�4�«���kW�>��گ�Un���<U*�3333.�ww~���wyJU)333���U[���}��}=�{����������JUj���qǮ��:�V��Ӥ8l�c��=F�MU�d�k��]���$b0�q�PدN��"vT�rES���aek*�M|�dF���"g2E�X*Z�q:W8�rr��8KK�� 	�!8�H�i.��B6\�0���}F@����z�TӾI4ܺ��n]2P�I�n�.��}�Þ:Y��WI��tg'�vH:<b���v��OI��{�/�^Ba���6ڄ�����m��\��%��t5ߨ���x��L�=�p��1��9O���ç-�un-Ӯ���m��y<�G��+:UY��`��ƇR�!f�[>�n�����F�j�L9,��tQ�Q����.֚5=3
��EsA�����ne�Zs*��b�0Z0�E1T=��B���(�F.�ģ+m˭׫������Vϴ�.��H�X�jMOv��޸ۮ�պ�p8pM�,љ:�7p�,��B�U'xFe+�v���̌�Y��8�J�^�ۉn8�SZu�4񍟠ԣ��`��5"AK��]ܧ� �eek�t��Id؍R@�ݕ������tDk�aڪ�����]�.��I�変��8�C&L:x�պ�V��:�8���I�j��T��Yr�ND��x�Fbg���w��()�)nu8[	F�]����Q�U��s�Ä��;��3�
��;��E�F�c�E�F'��54�f͕;�&�m�Ћ4\0wkf$�	�:�^��4t��8��[�qn�um�mo���n�D���""�e�D*�u��!����ۜ�ִm��%p@�x�39�̍��NM371f`ņc ���J�-�|�[\ERڢg%,*����r�ҜRĲ ,e1XF�M��-T���X�e�]�V&'
�9���p�Oi����*��Å�&q9ҝ��lIɹؗ�Z��S�ԯ��(�N��@%JÓ��V��6q9YCCD��Y�=��O�і�r�-�k(��f�P���,���K�h��X4M�Bjt�L9q�؛>6a�m���[�qn�um�k��I&�DP�T��Vja�d��ή�S~����y����kb�MjCIxǒ��O1��xQ䝝1�Ӛnَ���n�+���b�!��-�VfU��S���6t��݆����Ӕjjde�� �"�$*��`ԋ(h��<&͞<t��ӧ�:p8pM�,���(k-��U��UY�����cO�p�`�ZI:��I8���'�2x��7m�l�gL,���P��>���n��2��h�$j>NjZ�ܜ_/��9p7)ܛS�.e�I
K�#gFՇ)�b#[��pѺ�������WՇ�C�$���1���X��[�t������羐jU:�r���|Âw*�*l:6%�%51;��ԃ�G �K#��]����ڊ������=���o1��b���F�S	�2�1r`a�FeA4���l�k5��Y�d�~Z�w�ggw(�n�-ŭ��ո�N��6��^�45��b��ǊݶD
�����6[dd؆�n:�0��8N�7d-�47�8���G�+�qDӒ:��`&�!w��� �i���U��/ ���b��uD�u��c�Ɲ+�tJ�^�żM
�y�/�d%�.�*�I�F��A��xQC�:'��"�b$� �4Q��;=;��gE�fsWQ1��/�|F�Q��Mʰ�Ec4l�af}$ёY\MҶ�Q�B��;h�MB�xª& �' ��2+Mu��]x�\q�V��[�t��j-X�|� x��Owɜp8�N�1�֚ʪ������rcj����vfpً*m]h�4dǖ��]=�%<���8��ukn�OWO�;¡��`X쎡��ؐ�,^T��0�c�F������l.������u]=Ѩ���<��h�!ki�b:�L[Q1��q4ŵX�������Ʊƭ:�cךLLLx�1�m��>k�|�&'ε����<k��'����6�&%b��a���}���VG"��%�|�K�M[ly�����ŵ���a11�xƱ1��1���&L��w$֗�d|f�T���Z��V>.����B>|x�����D�D��1���M�Ѷ5�Ƙ��
�CC���\��r�����Ʊ��c�G����ƣ�Ǎc51���N�Rb-11m1�I�5�26��=LO
d��:
3��|�6&�P�O�<&G�`�G�k�G�u!�9����=���_c�A1�����w�[��}���a��Տ5��lk�=���[�Ofn껾���W�T��ƽ��S^,^�,͟��S���������ӨL���q��|��'�g��V�^��rY����>��>�/���Uw��j��{^�������[���_}����g��ޞ��{�����k3333/2ff{���ٙxS���:���[�u�����?8��$�i�Ui(���9D ��a}���a��jhI��}M��d��됱	l.憋��,�&lQ�3Tʫ$8�Y]�d.�u������0��0!�>�庶�<�9��Z.�hK4K��Ǧ%��D�¤�C��q17��!C!�7��x�g���Lٺ�>���*��!ܓA�>�e%6�5H�d��U�)��b6��P��t���`zrT7��}�i�0��$@� 
�'`���˳�>:c���n�ŭx���'�Tڪ�H���;(����%a�a!h�M4��De&K�/��tv�IUQBYd*U�1�qs9�e��D8b;�^bd�H�qȞ[Z27Y�q�|=*���)0a(99�aN��/��pAJ�Q�H$��O�i|��H|��=g�Uâ|$�FJ����YA�tH1	�!���&�Fs�ĳE�E�I�� �pf����P`��I��d��ǔy	�1o�1o�:�V��>[�:Y�F�'Ygn�Mݎ�dOK��= ���֛���V3�WJ���kw٦�&�sV��E�\o�x���s1N�g^�17��0��R8�F*;I#��vc�*CHe����}���m���wU���*|s�����0�5�8��%�J��>L�!~Q
20D���0�L���4��X$�����	�0m"ϧ� 3P�BB1g22HҔ��K�t���K�ȁ�	�8������bm؆�6R+xe�˥: ��Q
K�I�eC���\13���}%�M�2\�qZ��`�>�(�	�����G��:�B��優��Nv-ظH;D؄(�X����0����b��铔Pj0��ڊ����c�-�un-ӬxN�pÆ�]��Svq�:Әjb��TP� a�r!Ȭ2��&=���hi,�ɢ%DȆ����<2U�()!�$�!rP�a=~�uM�����B�c$�FICAl�U46��RRK��rVI�bCB	ڐ8 }�Uz캪h���C�9�9E��E���7fJ�f0~��:�4�d�"�(Uj�vr�\��I��	�hd�0�$� �r�'HP¬�_~���?%�fB�w�� py"6"�3H醠���"B����J�P�wn����2�Ԫ��� {[��<[��u�-�Z�[�]cN�������^x��R/�u���UUD=D+�*����60Ѕ��bK+���!r	��K�l%y(Ѩ�]";&�����M��7h����B��xf����R���\%�K=�v4���9b%�����H��xL�*"z	:���a�)�%�A4¸��u�	���܅7�eNJ*��&���k�����`pGa'5`�SF@��	�B�B��7촊
:��(Cq�Y�NX#I�!TQI�K�C��˚:��[���ַ��_4���?yǞf��œ�B�`��J��J�N7��*��v�T�"W����'�e��х;P�))�<�iQ� �Ī�F�R]%Q��h�?�d��[ˉm��!N��L���\�����T�%�bFr	����OD��0���fJ�Z~U��paʱ���T(8!�8in ��$��P�`��,�JlE�1L��V�Z� � �03B2a�[�fB{{j�&���EĖ!0�IbCq��� �l���5�y��$��f���-�q�-�Z�[�]cN�a�5>�|G2�r2�KR\KF��H�%i�\h���¬CWm���D�d"�Yl��J)a��NX��h��@����5e�dQF�
'��|�#,p���m��Jfn�%���r����x��do$j[������������`r' �"9fV�0-�Ᵽp`z&��dռ��a�&'"z��zr
��5Hd	�pJ0ŊQ��آ�\.'�ÌgL�]�b�XK�-/)�b��JB�ʅ�4T��$��Е��$�}�c@�"5RMu�����ÌQ���2q����>bI%�P�A�XTDC?d��8!���f-�w4n;9*r����q��t[���C�1}����R�)4d��u807����eC�u�۬|�ַ��XӮ?*i�D�RD
Ny8�vH�����m���+���ф����%�x�CTx�Pj$���"ʮB0�d�.�v�%�rE�NaCvؗb̨��UW�@�ó�X��$АD~���"\�a���#}�͋
�L�3�g���5n c�ؓ�Ɂ�E�)�;�n�0@�߳���� �Bd�(�mbVbc^2n�t]�I����9	8��`�@�D.|T�0;7(�9�uMU��!bn'(X�v����M	�j!��FqE��˛������r!2'g%T�)�o��m��uk[�t�>:p��ѩ	qUUQ
��$�-˓)�u�z(����D~$NC�I�Me'�e��d�/����E�&DHi*2y. ���ff�	C
7
=M�W3���.J\ V�2�,�&���E�␳�M�e�����jE���e%-тfA��ߕ�X��<&�w�P�Щ����c$��eYv9bZR!�-�)�K	���Ҧ3��^�TV�p��^y!��+��c��-�uk<p����8`�_KR�L���^ed�K.������5D�uaP`wgE��k�d�~I.NC��cv�%�c�ɦ� �x�4�D'ݟ�-rK��rh14��Ӆ�R.��}H�(����0.<!���h�q1�.��#!ȈȌ3#!������j�l1��AK��=�͈��1�a��ED�tPd �Dc��,1�`����D>7I�H��w"c��f%�EҊQ60�����ƎA!��ȏ��	�Z�Į��?��1m1n�b-1�=KLKcX�ƭ:�O�j&&&<c�Lm�&&&"�kI��5�b<cX���k�5�Ķ5Vtx�����/������|8�,��>k���珓��mu�^1�Lm�&�#�5����k�ܑ����0�L,~&}"\����<Y�r�Z��*���>-g�|��hO��ΎG��>�%O	��28	������t�X�N1�-�OR��ɦ���bc�y1�M��L[LKLF-�8�lkBdl|(�Q=�3(�r���DȘ��<8�
�<Q�	��^��>G�%]�w�����ib�'���u�7��,�eǻ�ݓ��>W�v?��{ѿt9j�f_�,��k�*>��رG~{0y���k�fc��ǖe�9>6y�>��=2��PC�V�9J�m��55���R��X��*� �:��8��ٔ�O+�ϵ/g{~�&���U��A}Mq�(W�g���3ڭ�<�4����Ɍ�:'�
�ģ�n.��+W����L�p8��CP�� �,A�[��/vL��۪�.�{x�+m��e�(�㕨R��a�-�suC.�5]˂�` x�{��Q\NB)BEr�|w+R��w@œ�5kݴ��i�������-�uG�sn�&��O��^2-�����ۜ�4��L�����y��?��4�Mw^(5�ң��}��nN�͇<��
��:|Rc��`��`�*����P]���3q3^X>̕D�ђ�zv�I�L Z��l| ��V�����9��ۥ*j�B

7X&)�r�(*�c��TEF7��t���i�J�加��̶֕<�*K
)k�)��s�(�v�$eB갌���QH��:�ꈕE)��3���<«�fF��G�B$ݮ�TTn&��(� DO�n��mC2�PE/��(�:�rŊE��V�彏�*W�w���>��k33�~�����33=�b���˽������{����V��9w~���U�i_s�w�{�Y8p�8�1խn-Ӯ��q�{��~xGE+�,ɐ�D���i���j|l��1ҷJ�x:�$m�嬊��3qI�u�U��$F��@�B;��\
�QX227c�|��m�%���Z`�Tt���CTD�l��2��\��2���Gc0��rDd���0��Ӆ$D��FJ�b�dJ����}0��ﮫm�`�*"P÷*K� ��� ���L'�ʆᔊ�ʆJ������f4g�S^QJ&�B�+A�����*b�K�Y(��jQ0�e�F3閭~��̬�A�ȩ.�w�]k;2����n��]��ψ�?��"�D��_��z�N4ۯ_>qk|���Ӥ8|pÝW�˅���qUUHZR��N]�K��@sɈ�aZH�%��+N5�r�V�
b��������_z������<Q�1�$0Y�ЬB�/Ѩp@�%&ɣt��+M�`"\���R�֩(��uWF� y��o�2��0p����^f�)�cW]�����=4T������4�|�Wm8�gX�w5�ʅ�`!¦��F'�XΚ(`QQ���p��\?~��c[�>u��c�Z�[�N������ �I�FK���⪪�%W����N�tp����3&� ��(<P�ޠ�$������1e	U�Cиh��@�u���Du�˺���ꢄ���(�pb��No��>}C��[�_sI�>j����t�S���֏��W���F*\U�넆f��p�.��`�*�ľ
�"4nҪ�5��,j}rpƄ��02+�M9��a^Z�߉���������(9GP�L ǩ^�yuƸ�����lql|��::C��;�5S��"ѳ�UUj��Ul�{[����Ε7,��}As��7O���'tP8�_���r�B��Y ���p�H۸�C��������=�1c��s6��j�1!�0�p�3����D,�oF`c���1=���6d�� �@l������u��a~��*��fPj!l,1�r��3�s�4�i��"B�sr0�(��`�4`e�1���C�l�UIWv��3
�M�MTg+��<��c��J�1��V����b�8x�t�0�_l��q���o�R27j��U].#2�D���v���d-�hf^R;ED��n�O�'��Ij$���2�X�V=��Z(�$�-+q�����#�Uk*ZUU��"e�#]�����wa*	vT�f|Q�ʼˆ�T( ]�\�Qt�Ś2���Ӛ��aSa���'&~K������{���B��(�~��12���Q��E��n`���|��Z��{�X,�%Gf�kG�˯����fg6vz��ܸ9�[K�W:��U�UTѣÇ)L�I	$;`�1)(l;���EkQ&�����qh��A[J��*<n:*��S�[U�ӯ+�u����qkb����!������ٍ��.���UT�er��a�<v�l;D�S_�֍Q����I#@�&�S��ɰ�B�p�s�`0�Ұ�R��·�{;Fa�\M�5VhQMf���׷p|e�&.A�)����9.5+	Lf�%Q�w��N�8`޼:4h��}�RVd���598v�67�ca�pIIS�9�er��N>u��X�lc[�]Gxǎ~�xI\�����	��?U�{���ܕ��_�G�!�AgwZ��e��D�`�pQ�\�tѲ\(SAȆ�!�Y�(Hp�҇�]�7�9�i.���6�e�cqIe�ƴ�$\�7A�U�E�p�>00;T2��:������W��տ��a�U�H`� �p
�%��ۜ���a�VS%��B�E�*l��&@NLL�z4`���Jj�)�ޱ�ϟ8�>[��ӂl�g���4��v����7
K��Z�
Ԥ�3SN�UT�J�ώ�mٹ�ٓ`kb����z�����/��֊�0[���#W	vK��Y�^2%�}�ˆ������a�g�n�D�a�0Yf�5�����<�a�d�Z���h����!tz{"�ȫR&���4x��(���"RP��hɨJ�����Bi$���9,��g�<|h���ϖ�1�:u�q��{�׾����<��� �ի�y��Q���g2cj�c�1L§r�F�U��,�r�$����ز¦(�q�)x��c�&��N�Q�� u6�H�UId�(��^JR�1n�8[��rZe�#s�Ƀ������_56v!��&!��^���ڑLCGOB�ʆ�ofL��ئB�kŠ԰�g͚1�(B���TtѐK�	
 ���4U�2t�;3NNC"���2}8LN�Lp=����i)*�j�,F;TC�҃1����ou��ZH��[l[��qձlcc�]GxǙɽ{�������9I�pY�rB����UUH�Y��D�v��̯Q�QTL"j1f�,�~���!f�����pɉ����NwK�!��pg>8J57�p��c�كA��k��/X��T���1.�%���.���U	t"/u��}M[�G(CE�f!�f�2�sR`�fbY؏�e_\҂��حu#�J�?g�u8�J�4�|����b�1mbZ1-�Z1"[[Ķ-�S���D�c�bcmbbbb�gH���LF?5���11���$�5rF��7&4�%D���)C��-x�X<W�Ɉ�X�j���������~���>���\|Ui|Q�񢰾4Y����Z0W�x���+�B'�^%��E
3�O#�]OS�bm11֘�������0U>):WG������bb�1��?5��3RxƱ8�cX��LԖ�����5[c[G��eI��FI"1"0�H�I��4�,J	���*`�G���f<4|C��q�I��ݛ��z�B+�7��������2��W�ۗ���@���=�{=�:����\�}=�[��u�2g���E�����l��m�ww�����0�|�5MQ�=�jw�s]Ǧ����®rT������~A�g+�����b���9w~���:U^+J߹w~���:U^+J߹w~���:U^*�o��߽�aÎ8�n1�[���Q��5�RT�וUT�ѭ����S�M��S%�j��^,�d�F?zGU��{>5E�ej�����	�:��܅˺Dd1��%��r��-n�揾�5�����sJ��`�)iѓa�vf� l�*�9Cf��۶�j�fd�E��d�|�ef|'�s�%�ҭZ��N\�ᑉ�~qk|������8�N��6����f^�8�q�q/�ig&|���5Z\�u���q!�͟;��v�C���(���`��.�z���pd1�`�(lqCU(�����p�ՆB��O�bCr��i�r{��e��(����>� ��wE��A�xQa�=_VF����i�`˗� c3���jS0	�."uu�s���J6��pi�;|㎭�c�:�8�ǻ�5�Z��^���¦�m��sr���Y\̐�<t�)�0�?��[oxH5�zJ,nB*HO��Y^f�cp��L�2����$P�|���.W������Z��D�R����I-�J��t*c"����K�a�_�UU l�M����"��)d	l�&�_j���g���n'ǡ��o�Qf&�A�;z�`��'�lj��;�I{�Cwgz�5T��w&�ʇ�ˇ���!g'>�M�4hą��PK��_S9Xl?zr���xcі���Vҿ`p�!����>�
6MĠrf�cn׹�<���̭�9F����S�&��8{�V�tpD7��V��U"�&���gp�t�8hٷθ�1ձ�u�-h�o�$�zS�.�ʪ�@kŗ]>��
���L���isfa�=5�S�j�͙p֕F�}(�x٬B��:��+���%M�d �B�һ�>�˓����2��ۢ�����WA2�ߺ�>�C����d80�ͬPXl�{%j�Q����sF���S�����N�n3�n7ch飇Ǎ��α�c�YkG[xñ��97��d��r�H��򪪐:k���M�U{�E��h�0���}^��Ѻ7e�7�p��m�e��WBQ��]�����O����7Ăm&�A��z�7k`��.��eB�^���C�C*�z���VQ�2�`|z����+g�\��V}�I���2�Ǌ�e�e���3r%�St�ν�篚cm�|�c�c�Z���,�$�R+�C��U��)�ǜ�UUH�+��DN>�3.!�+Scrt�0��AX��g�XG�2VJ"�mLEX�8�1O�rQ��p�r)C~>����;�.��&~���U:f���N|�a��s��ֲ<5�R&`ȇڒ�.�	a���2=ɨ\�TV'e�3�C��jlލzű�1���1�,����di��^VQ�'�|굵8ɂ��weyUle�f�Xfdx�5�������5Tf*�8�grcY�%dQ6+	b�ؤ�(*��7puq���x���.ן*��I�դ���,E��	�'jC�CG8r�.�e,�St�Â�
6��	�\�yV}s���S}�4�3J��f	�(�g���i�%g֙��fr���}k�Q,���d������5�T�Pc��ػ��^����q#cQ��L�.�R�8z��Wx�zC*4}G)��)��=|�o][�����1�,����Y¡(�ۃWv�'9�UU w�`�fbYa�&首��
�x�����v��=&�U����t�S��b�<pɸ&܆�������5MM��ѼK2sJ���KB������&5ib���nH�5�ln��!�6r�������V��O�U&K2tϗ&fa�у�C�ῗFD�,�1��ڹ>:x�ㅸ��-�cb�Z:��iɢe�#Q�|UUi!�Etk�u��/�n
��d;���R�B�G��[��Љ���5"U���p�>�
:z�<j�h�����!o�!���޿*�j��Z�9'$�R����lj�U\Y�)� ��D�əs���X4dK�R]������	�t�jM����O��[[�|����lb��]Gx�w�O�X�*���H+�e�(B��|�.�ZHYʻ!��[�Q���"l�a쉘~,MV��=eP�YEQk�|��7,S�*�R�"gO�*P��>�1*|��&'!�(Od�,���b'd3�U*`�E��(�)�:yR���MS�״"ok�g�G!ADY+)�y��Zԃ�9Nӧ���$���t�Z[�n4c�>G�h�m:ƚL[X��KcV�KcKLLmo1mZu?&�k�M11��1�bu6��1+k�bbz��X��k�b-�Z6ƫ�1��4�1=Oɏ�LLi�1?1�LLc]cX�Lz֞��cX�������&I-1Ʊm7&5�d�>�BY����L8? ͱ��EtP��Bxh���̌O������6�%|�\G��#�>��2&OR�9,�
t����m|y�>Lu�f�Z�ƢbcL�cX��LLN1�ɉli�Ԙ��q�ɍm+��0�#ʒV$F�:T��E[(��+�����2>Ɗ����W��=ѤӬn�m�`���^���]��L�cv�H`�p�}�3Z�F�̮@��p/En<dC�:��������j�,��S�rh�'�N�߮(�i>��b�{܋�qϥ^�I��&�\�<�=�͙��`7��N�4JWQ7��Lv�cX��7k!��ʁ��$��;�l���%�j�>�tkS}��?W�$о����$��k�7jr8��|}�(_V���Sf	Jc��Kq{BDLv�ϲn���VAb�vj͜#[��������ܛv�=���a���fĽ_H��O�����z�{S�:x�U�{�{2�{%�o|��p3	�2\�z�y�{��&���#}U]����z�����ne�W�f��dMzc;�ށ�<L�t^��XM���`���o7i��c��kw#չx��'�9s>r�="�\���QE��w��.Ǐ�3'��w��������T/�]�:)�Z�UQV��@�j����xE&F�+�Gk��;S嗒^-�A�j0�88A�b���J�1nd�d9n!�$e�U�T�8ETnB��mT1�u��ʲV)J�U#vNA�(�$|t��Q� �,e�s"�2:�*��j�*��B3�
�-G�%u��XveՍ�:U��+EhAk%,�V�G������⮖��߽�{˵V�t�~�߽�{�v�ڮ��ܻ���{��[Uv����{ܳ6a�x��<x���٢���ưF�w{q&����(��EQcU��F���,��0��Fq�r�1�ө�q�D�+�Y2Z�c�$R�p��`c�M�Z�N+SE �X6I�(��	z��UZHo{Vl*
�P� +��~[������18\�D+&�D<Y�2"&pS����5-�ܜ76}�,J��[>�������%����*� �͖':��Ça����f3��`�5rh�=�%��?]	ߺ�k�V�Z#�Zr�D�*��\�ywy��7�v_j��Oh᳴v���>�]չ��*<h��kqkb��-�N��6򸷲�$��ʪ�$=A��5\��5���f9
�V��vn8O�L�0��P�����ذ��߮�w�1jt؉�8��0|'�f�"T�Z��X==(ؚ<�	�	]>Ѡ��*%_���+\+j���m�ʟdu+1ga�h�4h[:	�6F���0gȳ�-�M!���
2G�rV�V�$��n����[�u��1l[ź��Q��#T�jTO%*#&��UV���&��*�Cq�J��	��f	)\R��T�7>�,Л�e&�MMtߡy2T����8�[I4�o7)��E�⌫X���3�ӆV���f��5*gU1oE�Ǎ�7
(L�9�P�:��O�,�3AL�وp�,D�GM�8���%�х�.\�(��N6x����c�]:�8���d�{5�i��y	�UUi!|��I]?z���%m�Ɏ]�[��cr0؇+ˌ&ؙ(�j!_��x�r��Ԕ��e�jg58r��遂X�Hw��̙4dEUE����'Ұk���fM"'a��f;�]�*}�Y�݋
,D�fn��0����ea�T�a�ʮ�ÂX�Y�s6R�3�U�4TGX��c��1lc룧Hp�gϤFn8���f9�F����=[��o��\�P���u���Z���H����y�(D#�L��8�GY�1�6ptu���r(��U��Z�GJ�c�"ل�9L��˾�UU��f�+D���ۍ�#�;���y����[4�-�h��;;��)�����2�b�$����d�	D-����dN��ǲ�շM]_�>�dI�nQp�xlQ�^���	 y���K7��^®m�����b	�nt����1�
:{=_Ǆ�ӭ�/�H2PvF4���
��QCgh�uF�:"$7�%�

+UY�4{����T���&?��8�ϖ�1n�u�q��{��qƙYr����BQ�>f��Y�E8=iL�0�GG�<zdK4�-�t��9:6'j���.-6d�P�=V$�d���l���3H_��!���-u���ݐ�#�mfa��N�5]�>�#Q��{�
ѣB�_�vE?�gוֹioH{͐���h�"Qt!d�|~�<כmߞ�x��o�b�q�b��:����6Y��}��Y4��A�|��T�1�y�!�l�=����Q���E1&��qC3��=��(��ʪ�ѓ0�Q��,L�3�j��Blm�rI��(�N�(����U�D����&n�����m�~Uc
�S�"B�MvI%�P�>IЯ��N�4}��v�!�s��UT�U��İf�T\Nl~�v���׍6����[�-�]:t��9�ү�5�B^<UUj��/݌�8op�>��Y��;,�+��h�8�%��c�#H9Z�������VqU��
���95y�c��I�93���'1x/L����!��%�1\ڵ�<�����B�d�blNC�0\�܆�ò��*���x�gN�6�>|�1n:��Q��/����I:�qE'���!&?�C0��z�I����v�x\�-�tʰ!�&ř͒D>�t��F1v�,�k�TA:�S�v�**n<N��mX�.�]��J-��k�ʪ�$9|�u��R�B�Ed���m�9eUݖ���UR�.p�}�8lJ6�S��N�G5M�0&`�����}�İ�J*bv���_�"k���S�Y�91r��!�;/g���#�R�Lͪ��}
2&!���2T�<0BT���bgW��X�QĐm2��#�>G��x���_�(Ff��|ƚ��Gꕸ�t'M>u�-o��-�]ui��5�.{�#>م�8�%V���3�/C��5�Q�.^����C���h���`�M%�hD�0�'8��+��wvY��QٸMK�4"YSpf,>4��|l�-M�>�N��bjϵW�X�����e�Sp�p���^��hH/	e�r�7!��IR~���#FD�!�L��Q��e��D�j��v�U���sN���:ź�պ�D��:'DL:"tN�pЂ��8�"AB&�N�҄Y:X��4&�١4A��L4 ����:'D�%��6hM2P�%F�A6	�AD�0؉ƝYŶ��z��Yn��?1�a�ǌ4x ���'K:Y�ĳe � �	AL��4&�K�4z�OO��6�j��vӐ����v��I�f��os&�3˫�_���cs�տw�s��qŗ]Z;�ktk%������q�kz�v7]��ˏ�N};���?���̎�����Qӷ3�ng��wp��5=�o�=��&(�����0�C^�_�W�7�P.�]~����L#V?NEٻ���o����ss���9|�w�_Z��������{�mWj�ۻ�/������~���Wm����{���ڮ�]�w�_��Ye�p���Ǐ��:t���e��u$�����B^�j��u�_���Q�f���G6$ jf��-
���e.�S��]�`y
e��0p���>�z��ӵڣ�IQYG/%�G-�R[v�cf�f���5T�	��'���a����ɢ�����ܳv7蠱c�G3��G�E1,�e��k��m�q�OB�<~m��cn-���-�]ui��<����(�ߪ���Tޕ3Ͷ�o�P�NB�7M5>� �a�bQ�/�}�Z����+�����B�Y�P����{�%����f<c����>��pЇ�a��}f��}�ӂ{s^¡�Ǎ���00���&<������"x�&a��n��!�(��M|��Љ�w���wp�{Kn��>u�V����c뎺�ɮ�Q|d�@�\�+,������0�F����e�	�� ���0�8���ֵi��X��Պ"Ѹ�c��r����S��-�AVX�n�s$#�X�ʼB)7�[m�4-ܺp((�e ���(�(�D��`�
T�MAN�rQ]���*�ek0����(O�<CQ��\�B<-�lS���%��9M��!��Q�1sU4+������#ƈ���!"1�$�Z'��?p���~7X^	u;O�Ny�מv��-֟8���c�1gM�:C�p�d;�u�Gc|�UUi!,�v��˭ꏽ"p�	_�H*�12QBx�>��1�,�������vpĲ��N���I�&MC�lMos�_��t�B<��UuG.��D�NK��I"�R����8D,ɩI�DLʇ#��\�~Vn��F����=ŝ��h�h���1�|�lZ�-�[���:ӋT_c�`�k��!��E��+8�UZH5�농��4I>F����L��K"P�%aANCpL�2k�L���
�#r�U(�%�D��(��y$� f���ГǨ׈C��G+t]<���k����D�S8�<%�}����bw�RST�97�P��_���zc�?{ӳ�x�3���̤�8
N�����\m�c屋u�]GZq��y���ŒZ�R��*�����]�!��+�]�im'Lû rQ�!����4�/#2�ĺ��E�6T<YB_�r,�f"��O��&�L�CP�FL	fl�s��2'94�bT�R�J��dȱ����Y����6x��b$����}�z4ف3*�b9:Y���n-�[�^��:Ӎ�ns�;7�Y�bVE���P�o*�񰔂�܎4��qKCq�ITS*��M�ج��XE�2�T��ԙ;�NcZ*� �7]�W+qj�P�MI����Á9B>D�'!{<�m��Я0�V�$��i��(�nD��f���9�==3��D�q���5Ye�6�����#%�+�M��t�Vr6bxɉӦ�ٍ�R��}��h�B$��5=��ώ�'��֍SL5*B�E��E\�0s%`D��9����^6��c���R:�e�яմG�qy�~}i�3�v���mվm�1�c��]GZ8l��}�� s�UUi!�ܢ�@}.S�V��ѥ�hW�0��І`dȃ%az	]u��f��f��F����p��j`�1���ڽS�a��F*<�S"r���S8/9ĪJ35>�eɃ�12g��ѱ*1�Hn�!�Q�:T��2�]krG��X��bض1n�t���e�6]��$ֶ���BW���b���5]�8&��z!����J�S�򭶛F�]i�*S7[u�O�għQ���53,��ȴ�ś�d>8r�sF�f'�֪���f��s����S&h؎�#Sް�H�QI��D�5S�<�Of��f5�L[[>[�^��:Ӎ�qu!�х2��e2�!���UUi ���k����%����=U��ǲR��!�V�eYo�!��]@���JGg(�Bh��4�����FG~�%�ut&�.�K�X��	Is���HS�l��'aYm��P�2X�څ�E;
��jM͈�'���E��%�~��?F>Gˊ�)�%mc��|������: ��0L,���4&�4 �M�D�:X��4&�6hMFH��0D�B�DM�"pD舜ı6hM	BP�%	�4A6!��Bp؋n-ǺOV���~E��1�ŭ�1׌1��1��[k[�mk��K� � �"%$fı,D�(���R�ꚪ9����ߺ�qE�|���^6AL|��ye��(<�]��*���7+a떩�+���9�-���S�ܚ���k�s|S�����rS9cW�wn�m軕v�Dս�p����:�o�C��Z�T�1�eU֫N��Ck�E|w�n[�di1�j��V�`U����Y�h���M���52JʛVG��q�g�*�Ρ�1f7�g�==��{��ô��eY�X{���4.���ܑ�j�uI=�	�^��~�oڻ����K�9���7p��{���mU��7Y���ݶ�W���0@�b<b�>�����=��]`Q��e�,�gcx�MmΗ�k;<),��\S&j��٠t�+i�袑�+���9������F0�R���8�g+uI)���V�����ņY
�i��AJ�y,�1�!S�"c��/���H㍃%(@�MʂY*Ln� YxB��h�a+�n��RG���"�"Yǭ���$"$�R��ڑ�ۭJ�B���"l֧�`��iApq�ci�렜U��lmV)-�V�4ŭz�̾=v��ww�{����y�U[���=�{����]*��������{�x����}��sy���m�m�c�c����^Muj���-��l��R�2�D�٘��ڰ�ʢ-P�̮PpM�(�ڜ��Z���Ꭺ;�����&9l�#-�@���^]ܗ�y�UV����n��VB�K��wv���k��'Y�U��9
qP�Y�
j�P�:.tX�A�w��}���r�D}�iԦ>�mnռmW7߷A�P�(b��w"!S���S*�V����cd�r1W�m`�X�E���q�!3��$�
<>>���b=Ude�d�F|����>|��Ÿ��Q֜m��{���!Q�a�z���B��ՙ�"���!�`�M�(J�zqE��A=��9F�W��{V�S�c�E�"=y���d��nʥI!�v�7[��'�'KYii�va��.�!���2�Ѫ��~	�$=�1�[��1����(6WC���?=�V�V���u����c[x����Ν!�8l�g%Z,w�ꪫB4{�}�Q���A����mN��rt��F��`ƨ���>,�X'�8_}�M:>�gB�/m�^8�N��Y�ƣ�����Kx��D�otIr��n��u<AϮIQ� <4�,�5� ��|�ĩ��N�8f{y2 �T�s�.'M>6q�[�-ǎ����o����so7�^om2�7.���К>	�����&��@IeOy_�<A������\j�Vۂ�Ijt�ZQȫmyCpѭ�*F`����d%G+��႟};|�p6`���S���,ٯ+�@؛5�7.e��a��u�3 �175���RY��c�>�1��Bg2�l}0^C&O�)+Z=�kT�U{嵭�m�c��q�uo����:C�p�c�y��j��35��˷N8�0�\ቷ1�A�R(�O�淛c#T��1f1���S�X�8��Q��d�Z�H�g+'$�VF��Y-h�Q;���m����P��J�%,����pg+��I�I��:5d�afe���V&��|`&|4r��d/qb�%T��2�u&O��_�B�����S�9���`��H,�,����U�,!����ѧ��=\��9�W
��,781��`(��e-
R
��,S1�2�L�p�a�?Q�pxԉ*q�|֫u���u�-����,����%YR<��KXa���Ȣ����П�5�����Bm��k�*���gk����ý:j�2�H)2YPC
����jpK�b�/�)/#��9"��!��r*�QWP8�� "�#���p(2w\�y�iWAf�b;p�\Dh�`9�ͱO��(�0p����康�[�ui��<ǹ���ɦ�}/S*��'�(��>�HSJ��A�sp�.Ph�}�2�ٓ�E�pѰK�������Q�DH��46�񤨡49�4�k��h43�C�3:���-�1'�?S%}^V�:i������~��ML�zE���b�V�Zz�-�:�V��q㮣�8�ƿwK��W��Q4o���	څ�p��W��C�K$��vnL�ר�t�sVVP�PR's�� �UUĺ��rE?|?e�G�����.��,,�dO�}ϋ*l(Π�P�wr�>�O����5��hᣟ1tk����Ks�'ϧ�T���<e�|��[�|Ÿ��Q֜m�I쟜��L��Lu�f4˭lw���P��n-��	Ɏ0��rD~��ؽ`�uLe���M��g]:MaݐQE�Ap�c&56�t"�tW��RVʤ��u�=�Y��^�DCUk6�n9ߕUZ��� �r���ऑ�0��*1�F5Ux5O��r�9=2r�i�=>�
55��ft��yw	%�t�t�&���}����p8f�[諼�ɹ0t��|�.���sef8P`��۲��$d@q���11���_��z_���]�|-N`ѣ'q�έ�[�ui��7�ɯ�׎�j�i��f��UV��4~��S!F�M3�UMU�\�t9;ɘrd�yj�d�O�~���l2`�C�b�rɂXY��.�+�b�T��0��"Z�1=�p�&�隇�!��oѹw\���_��!�^Q���u�X���nfʢ���5*$;��M��i�7&�|�X��[�un�՝:`�a�B$6"lDD�A(M�'D��p��%��͚D ��ȘP�$b"pM��:ɇbl�&�(J�"aU'�!�A�hDJ��N&�����Z�lc�ŭո��Z-�c�1�1��kun���޼P� � ��P�dM�_/�W�ɝz3����=>˗�S؞k/8>�s�{.J�+�}~����_�Fş|u[�/M0�����>Zh+z/��^ݐ�Z���ۛr݇E;��ʙ{�2\�}v0Z�gU��,��轎�O�~s�2z�z�_9�����������՗��]�]3����7cl+���Ϋ�1��R���ɟlL?T��2ߚ٣�k[��{��:�J�www�{����yťU������{����Ҫ��������{�qiUn����{Af8p�x����ǎt��$�g�Zڪ�G���t�"��B��p��(�>�>8IHl�j��0d7-Q��7T�h��
qB�q�X��j`�ag��F���ڥM�ѣ�ժ/R!2��
/#�l��t\�r}�f���n�W�z����z���8�n��[�:C��6Y����n}0�P�s���a0����~"d�&�0h��C���2n{��X1-�1�&1jRZؓf�75Qn�1X\!!+�����u���{$�إQ�C��s9�4�`a~�Á�'Ǹ�P�V�q�M¢�����{ERW�
�_	4|Q�u�Y�若��������|�B��[cn>q��uo��:�:}QO��_�B-�U�T�9��N[�Ly��X�|u�؋��8<�S�@��2�1�e�s(<ݳ.h���j�Zܜ����S$��⪧#���&Ʋ!�q���m�n�����B���$�+j�5�4.D�����k��;G����1�P�dgN�zD���e������1�ܟ�V9���_t4z��'5��U՜�4t+(��3�!��B}(��!IO���i��_>3��q�3�r���l]o�6��H���GQ�!S���R�~�q��|�{�����ξ|�-խ�8�����6�Y)ٞy1���֕V����!�I��ٯ<w�r�g)���곲�9�c��ep�m�����!˗��u�Ic)}ǂ��S�%�Su���fZw���l�1��!�/��>�]R�l���3�k��[�<��K����3R�����k����g�3��-�n���q��Z�|�8pN�Բ��+X���IK�mUU�4$���/��5!!�a�-�I�h��)�4��(+����cCt���N�,�D~�����ª��rE8�:J�"�+j�4MNCs��0	S��k����٨fbv��)Y�!��LC����,pƮ��x�u2��0h����q�uku�#���rM�UίH�ع��֛|��ЙZ�		U>�Y�h3YU��ұ��p>�U^�'r�Y.���RX�e:V����:O��~��]��h��a��Ѱ�$���ɓ"rT��̟LO<R��wP�Qx��@��|b2�A�T�C�6�Ŋ��l����:t��'O��:t�J�8{c\��;l-"�8rV�s+8۠�r���m6ӄQ�nL��%�#��k1\���t���&�Z�j���w�R�Ux;�R��@U�c�i�	�+UmF
��"uX�H��%C�N�I%i����m�ŋ
�(���`�)#�F �ӻ��Q�~�!
����m�>MSF�N��L��:8f�F���&�L7[��7K�%��S	�)��f�O��Y�Pk!Æ��s��UG߆��CP>�����.^cw��&�2��1�/��g9&�l�ɠ�}�~�IRO)�5)ݴ��z�������bp��+k���}M��m�J�����4hhB�G�Qg�Wk���*�ⶫ8be��b���q����&��͟V��r��Gա=�jp��?���-Կw�0����c��ˑ���[Kn��0+\�0��~>��[϶fl;�G�C��f�'t���{��u��z�|��V�O���I���W�Z�c�ʪ����OV�?e{���H�=G�͇j}l+�>�'���R���(�Cz�&����F�~�f+"���	�5%��*�S�M}=Ee�)�M!�sLOo{*vd5��sTSMM�0h.�8^T�h�|~������[q�uku�!Âp���DDa�2��
�w�UV��2����!�p�X(��bz!g�(�R�m���\��V���\5L+L5B��Y�j}K5'نL�>g�NONC��6�
Jfϵ*|��*}e|4ul��X��H���}/�3��	ߕ�N�Pw﷿LU�eC�%��5&˸u�<z����uŭպ�V��X��0L,�(�&�DD�P�&�Л�	�"&	�6&�؛!�"A��p�H"&�D���0�h�6&�	�J��2��� �	͑bl؉��Y�6~akE��z�-n���Z�k[�ֵ��-�cz��=x�ADJF�M��8&�/��5'���I2F�)�>7NW0����;{;o/����fe}�T(/	�f_Җ���s�xy�U<e��ʜ��zz�o�k������O�f����[��gj�Փ��>_x�k�:>1���p��Vdc����wc�q��`�����d����۝Sz3&�qz��ո�e�>y�+-���"�FU�R�`��e�m�"�8ЙXn,E#�q5��>5��z��s�d[T����&�dV�p�U�a{��FǍ4*��)ty�q���u[Rd̝mh��ʽ<W���H�sd3�t�����"x�~v3.L��Ж�d�*]mخc�d���{w{#Q��봋2c�0ͪ&K<�<μ���Vz\w\u�]��cQ?���������8��_����"��˗G�\�_ ^Y]��7�ӊ*Q�'�v�#n�(Kk��"��5X�����HY�2��
����.X��0#U����bn��N+�#��!4�,r���X��ƫ���9����e�>0n@�Yd *c���v�Ș����7T�$�I$r.7����A�� I�*K	mE)ۨR����&�C���㟎�J�wwv�G��{������wwv�����{�z�U���}�{����=b���ݾ��p�:a�	խ�8�������᩽n9����,�(�`�i�b���J�+���D�AK����Oƅ�r�!�'cr�U#d�@���!�%(A���vZ�DVL�K��K�&Ip�GA��UU�(�4z&�FIBȥ�r��$Nj��ΛƢ0G/&
�oV��l�t���]��H:�jw*8�Z��tj�Q��?`�d{�H�MUp�z�W�j�O_#�[��>h��2~����*ԯ��<���R�T��ɂ��a��d*N�O��*����w8��>z��8ź����u�uǍQ���rV�VI�6�u��#������a��a���EH+[�Af	w�$yy3$%�I���)��!D�YC󶭫oC0jv!e�䢔K����`�MAIeI�����a��19G��TI��>V3\��hу����0��&� �}�LK�Ͼ�T�57���+P�Q83N�~qվu�-խ�8�����f���q�����f���f����,���J�JF�K0,<g��l�D(�ʓ���8l6��:l�_��P�W��7��LPa 0@����Ŷ˻K�˂Cr����!����+�oW�����g���_�d��-UG��6M�=l�5 �a�UK�
;Z%nJ0p�cqkuku�#���<m��"�c���m�� 8��}�$��|���0��w~ת���v7���^[�"h��n��)�v�XEA�
Wa6uh�ff&e'ɓs��l�%i��+���=�u�Nr�'��2L�ð�Ærv`�sKN�V�Caw_�H	�+�.�1���ɢ�jJG�{O�*�x�:���n�:p�8pN,я(��in�l�E�dx;�:�i�""w�%��e�IT��fb�2���|�3�8��3�;�&:�oWc�Ibj(T&��U���(�%��
����| X�]�(ء]r�؇W^)�F0�TM60ta�*��nL�>ŝ:rZd��M�&��0�K�����Ls�]���ق������d�p�4l1�y����xLBb2��]��%���E�Lݝ��tn�=��^��խ�8�[��>8C�Ht�f΅�FǺp�YWTo��x�azC�ga��,�#��d�3��c��,�r|�O����s&�SI_OC��ό>X4pp|o?-Z�Rr�E���ԲV&W
�-�2� +��퉍�F� �U��l>!=Ӆ�J�Ȉe�L��0�*g*��EA�(L��=�M��&�c��������l:�:p�d�b�>ڮ��$��W�����]�4���kF���Ç���Ջm���Q{fdِ>Ca���`��I�1�$@o򻋗��	�0��Hl�� nU�P�dْ�V�ݐɳ0�,�V*zzd��sY���-����2U��#����5^�۩8��[���X��V�[a�Q�6�J���k�O4�)���U����^x��]_g
ɛ�r(b��c��CpԹ�'�V�	 �[�f4�f�]��.��Hvp2Y����-X���602�vd��|�=�QCR�J��\��Z�;=n��yW��30�}����f��-�[�Z����8��V����Ӥ:p�g�=�sw���]���s&I�1S\n�K�M�=��ծ1M�cy�ݖ���۪nnAKTV�\%��܉�������!L��R
*W�v���"� ���z�e��T�$�D2���-Q�8����C�K.w�:yS�rֱ/
Pxڱ�;����}��!_
�a��I����|�i�F{�8ܹ��a��E���U�G�h�5�a�d�
3��|
._Й��h7/l��z��뎽|�8ź�����L4p�HP��=tl�ʚ�.��E`�C��˽x��蜟M�e�?��.�!q���qf�S���(�n�!S��uW��=&����9Wm�m)MZ8�⒖���7��Ņ�<Q�D��6��{L���ᢦ�~s��qt��6Ӿ��clun��:'D�:`�YB"P��b""&AH"hD�(D舘%��6&�2h��$,DD�(A�6"&��&�6&�	��&��̟`�A �:7%Ȝ1oQ���1��u�1����
DJ�L:"tL<p�li�i�a��Z�kx��2&�М�w�*oR��K���GD�jwl�z�؂�-�U�G�gڼR���6�<�LF�=����sfJ�jfmk\�^;�=��o����k_o����]���f���}1e�\��uL�V����P��K����x�}/u��dǸܟ-=�lx�_�y���W���'}�ٟ]��};sS�}�G�w��������[��{�m��7ܫ'2��m����֣������f��}r}0޿�N�ﳽ�ە�Qp>V�/�ٕ߷���Ow��_Əc^��s[�9	��̯e�ǵ����EU���_{����{�*������������V���}�{����(��~��y�m�q�����l:�6Y��:UXnl���7m6U�{=/�s!��K��Xr�>8���1l>�C�l��}vm����o-���H���!"V�F��}��p����Y<���䜓�'�ȓ==��r�N��l�F۝{<l��UZ�������g��R�`�n��-խ��u�uǍ��g�����Cw�uUa��LL�bfL`�㻖*��U�J�ݢ[T�1�1z4���h���"3����l7��f�Zr��<lc��	L\ަa��^j4�p3��R��n�U4{+�m��[�t<����x�i�m�V����l:�:����?>�E=�n�0w$3�㍚;�m�������Tb-�al�8�6�Y�kS���<�I-f,U�9��dm=N�J�ASw	��0�r��u�,E(Dq�+[��Yb��>�S�� ⮛��%V�I@�Ct���q)EL��x�r�C����Ӱ����	�*"j�6qY|l>�>��cqL��G뙜7�J5E��s&�&�J�m\���n���!��2z�7쇾ˢu4�I��
8�Ey  %�jt���>,����-ŭխ��u�uǍ���o������I�oV�31�:l17��<Ud��}���fԒ�L�_���M��/Ɗ����};ՊR�ɻȿ{�A�������>��U�W���?k7v�-�X�`�Q��n���&n�}���}r�/Q��Oz7�}�=:MNC'#Ǘ$q�c��[�[�[�������U)��kj�0f\��e.�L��dwnk\���r`�G��ʕ��������Km.�nT�4h����M0^�f��ɟ��Sg
���=;fM��ɦ�"G+״}H�ϝq��un1n�<t��t��,ٙ�7�R�5��3X����>�}<n����a���'MLQ��3�a�k=X�g'��;m��A2�Ͷ��j������9�hQU�15&4/J��v
Ar�h�d�&Lÿc5WW�z(̗35P��rL��H�>X�����=�����ձ�6�>[�r��8C��6t��|\��ز���m�X��
�b�H�KF��+�d���Ur4 kM�ݐ�4�U\wܣq>PT��DV�uÖȈAl��
��p��̴y�mXZm����:+e�Gf�t&gP_C�
.Y���[�I�S3�Oe�Q�%�S��*�I��=�9GR�Leo1��&��5ɣ'���2uf;a
�\���\.1���4��UY125xA�b�y�NO �]C&��7�-'�t�Ϗ8|m�-ո��u�q������DRH]^p���7[UP,ǏOѲc��kg�'!�?�O	�5t�����g�5�����4_�ir6�ݖY	�gw9�7��<�Rp�F4`�3�D.��Iq�R�%�u�� %Ȥ��ޥ�Q���C�rc�l���&D�>�\��=UM6���{���ޜ�U�q��[qn>[�p��:p��l�'~���7���!��g|����1�U"4f��3��6?mz��3�r�! ãR�=3�6}3��J�r�2�]殊J	lv86�(���@ ~���Ş�v���v���.�N���uBd*�N͚�ѵiFn	��0�|r|�d��]vN	^�r���f�>u�c�[�ql:�8����S�"�kfr
�ET��� Nip5�UE���v��NNt�F%Cq�؛�Ҫ�RKH�tm8�mK��TҚ��$.h�(�&d6��E�ߨ���Hv���7T�,E�i�a�(܌�b9g�髩EYt�M;�*�Μ8zbn�5���wx�V��7�Rs�6O� ��I���/�V
�
�D��@%~S�^��'Е��{XG�t��,Cp��6�E�1A,)����*$�˗�@4��H(A煒b"#��$ �b1��(#�0D�FF"�#�H�D`�`�H��DFF �"#�0A�� �#�#�#�H��1#�1��A$��`�#A�DF"#�"A���Db0F��A �#A"#`�D`�%ԡ����Db1��DA�" �D��H ���1F�tIpD�"1��DH0H� �!��D�"1�A"�F�� ��D��� �Ȉ����� ��`�����H0DDFDDDdDFm%b�B��0DF	FDDdDF��a �b �D�ȌH ����F�0D� �2"#" �`�#�"0D��F�0DFD�#"""$`�H��`�"#"A��A"#�#@D�" ���"2""#""1 �"#�(��
I*"1����� �0F �� �#1�#�#b"1�#b$F�0DA����D`��
2#A"#A�Db"0DA���D��0A��0DF$��Db"1
I3p�`����Ă#���D`�##�"1�
0DDF"#"DH1"#b"1 �"�Db"1 �Db"1����"0F� �#bA�1���1�J�1��`���#"� Ă#DbDD�F"#`��DF$ �"#���b"1 �D�`���0DD�F"#"#Db"A� �"��P�AH�!HJ �(�"����
��A�CBR�UR�(�!J��%)PE)P@A �T�R�B�T�T�PA
��A�!H!U�(C����h��ZBP� J!U���U�U��Z�D�@IE"����T�P@�R��+UT���*ER��)PJR��
ҕ�����APJ��AAH%U!�+E �Q� �MRhD�T� � ��*	H%AJ� ���AJAJ� �� �JAJ�R	PD� 2 "A`�D (A�"
0�@��b��B2 �$%!JB�BTBR	UB�P�%T!� �A�� ȂBR�P�D"�JB��!R��JB!*�J�D"���BR��B����*!��� Ȃ �2!$%!JB�BR*�)���B��!)���yPj���"��2 �	��"�"%!*�JB��B� �`�"�"!DdAdAdA���BR�JBUB��dB"�"� �" ��0B0A� �2 �D!� �B��JBR	HTBT%�%!�	H�!� �a�$�Ab �A�"A#"�DA�A�0@D#�BT"���JAb ���0A�!%T"��%!��B��J�!)��B��H%A*!�A���D%@��J�BD � �� 2"!)BR��5�G��@`� � "A���J�A*	P�J�JA)A*	P�A)��%A�
�J� ��"B"D��0B@b
���T�RR	HTJB��J 0B0@`��W�*�H% �� �BR	HT�	H%B� ��R��R!R����	PJA)@��RBT���ĩ@!��! 1�F @bb�\@`��#�"�`���1�F �1B0@b��D% J�JA*	HP�H%A)!R��JA(� ��#`��F ��T"��PJB��JbB0aI!QA���J�BR*	H%@�EA*	H%B���%!�B1H0H�b�b`�D�`�`�b�A�"1F$b"0A� !��0A��� 2	���pǣ'S�	����2К����'��IEE#Qc �@���Z����5���mq��rk�?��Nb~�2?i}}_�Kx�cD!���'!��]�<@�$;�3�(�>'��Nrt+����rt�w(�QC�]5ܕ�o�l�r��;xy8��'Z�����:������'ځ�	�#��P�*!%��z>�K���;O(���%�W@������O1�V<��CԢy~�EPø_��<H��A�e[���oI@���Pl1bY��I��\	�|�))?D����4ys��ɷ���Fb��o}�	xa��!C�3����r����ADP�R�@�V�ET͐(AP* ��Q-P�`"��� ���l/v0g� �P�@�N�A*�M���݂�`y�S�7�#�T@U@�L�A� F ���E�� (+ B�KC!��|{��[�2n�ͰY�"@���lqඃؼ���G g���d��@����޻͟*A�*�4�a�f��}���p�?H�������9 �r��y���#�x>� |���%��$_�r�{���XWR��8�O�����TU�C�,i�����J��0hѱ��! �C�a)N���"� �=
��?hw�։���l~�	�JS��,C��h�^8*��'��%��{�;JPD.���p7awɅ`�%��P|� �l�����p�� Xc��(�24��'ޔ�`�[��Ȑ��Ӡ �6���}.���	�	5�'�"�����>cH�k�{�@{���V�6z�:6�{���O���w?/P�A������$:�<��'�}I�( ��C���H^��z?����:��."��Rt=�D��'g�ޏ�A_�P�>?��7��h�� p'�;S�;���8��&�c��X@�$�QD!��ϔp!kb��è}-��Q޴.��ѣ��=i���G��c�.60�����TU�$�������B�3�'X=c����rC���=�����I����6� 4���7M�z�n�I�"�Q��)�n�@�Gq���:��� �pg�=�9[������g3b��<Cm@0��>��"H��J
A�@`/C�C_�.�p�!�*��