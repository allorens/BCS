BZh91AY&SY���`߀`q����� ����b!_                                          � ��7��P ��   P    
(    
     (� @
  E  :�UP��� ��T P
  J���@ 
U@
���(A@PRR $ 
_   �@����P(�����qQ[������;��Dàn��P��䣐E����@. ̐���/l  ( o� ��>���q�UK��{�t[jT��=E�ԕ[hWvꇳu��7��)y�R�X�:�� :�@)�@Z��݀�s`Ǟ��  4 |  �@*BA@��@� ُO���z����� �u� ��ް^�ްP��8��y"���y�9 �   �  	��
���C�燕�l^ �sH������� �x� yˠ;��� zx  QE� �R��P��)*��P_Pf�� w`�@n���` ��P0 d� 9 �n� ���r �`��P(�@p>� ��@]Ҋ 1���t Gv ��:� � Z��@� {�   �  ���QA@�$�*��@�@�n�v8tPp �tɢ@݀@KE "8�;�}��� ;� � C�`��.u���@������Q��9 w`: �� ��H  �  ��I�@ �QJJ�  -��@��9� ��E΀n����7X#u��(p����� h
 �  ϰ݀-�T�C���@�`�@[��R��r ��s |       S�JT�4i� a0L	�h��JJ� 2h   ?L��"54      ��ʒ�h�i�#&��	OԤ��hbaCM10FѦ� Ҕ�FMhQ�a�4�jb}_/�2�~Ϭ�� zNw���:����ﻮv�@Q^ w��EwES�"��O����n*��ϼ�86?���#����G�>?��~�>J��*��������Q_������'Ĉ�
������xDG�d@� �`AS*���͐���UE_����� e 2 ���WL��EL
�� L ��C�4��i�Wf�i�4�a0�CL��@��.�L	�@�(i�4��eM2���4��a�L���
i�t�p��t�:eM2�S�D�
i��L���i�4ȚdM0&��D�$ȚaM0����t�:e��SL��Dݔ4��`M0&�L��9d0&�L���4��dM2��v0&�L	�D�
i�:dM0&�Ld4ȚaM2&�L)��(i�<et�0��L��D�i�t�d0���� c i�4��d2��L!�P�(v��� l�`2�L�� �"i�zaU:e@zdA�QN�Q^���2�:et����� ��L(�D]0�:dtȀ�A�#�Ot���"�L�2(:eDtȨ����:aQtȢ�ʢ�|r���|�Y"'LU��/�i�&6Z�&��:wG�A�������������0��p���HVsW)ה���ͳM}~Mp�Y��Ʉ�k%�\���;F�ۧT��h��6\�E{��z��[��Ͷ�5W��R#��A0��;{8���UmL��v����,sh�uk� �~��ҭ{F�������8�4>�6��²�WM/A���7��$���o .2�8��-�y��b��,^�lӰ!L:���xQ���@��^�T:����n�5	AH�Ύgp�x���Uy���Ӗ�d��w,w��Y7N���o/�Z����٢�C���q�r��z���.t`o���Hh��R��>[��˂��@���w%Ι�p ǐP�����l	X��I̎��u�]-�,�tX��e�����x8��O��
n���r�ȪwDWF±�٨ e���M�M�Zy�XY��֤���(0a��_�ו\��TO�.�Ã� �GU�l������9��
�ݫ���gCz��!os�M<guc��(Nr��e+6���f�tx��N����D��m5���&�١�%��>���8�-�~ѳ�S�tvگf�wǁ�&k5&�yFou�cy6��>ɮ�E�{#%风�CżX�a����
�Wh�#@��0�{�����lOfSu����gio��p9��e�]�<zu.,�9���;\4�e�=�IC���!V鸔�X�>�Z0ɉ���@0tK��;sM�X?dN@�����1���Xe!%c�����p�X���ݘ1hӋ�ݔgq�=�b���i�K���ATꂼ�M
`� �v8��Qn,طe��%5��}a�[�0��W'r$s6��x�DM,{���u��xZc�v9�Q&9��,X3uX$�nZ�jʃ�קv���#��od=�\V)'xm�6kݷ7�`��\s.��n$6i�lƷ:��/�^-�.źrٱ�2}WqPwNSu>��|��w5>a�ZfmC}�iw�z��u��\��v��n�˳�:�������#�b�_���Lx�`UF�P��M,��T,Xc�!�SB�q/\6�m�sT�����wR{�	��`����=�Ʒ/\yD/������̰	�`v�Yd�pN���S|�{���\��f��D{�M�L�o�K����vm��n���9�Q/m�f�š���ŐV�n��1�a�oT��w�zܽ��������tf��^���`���a"ŝ��'0��ǷJR�e�޸���rA�H��n
�n���X��c]՛���j��>1(7;�n<ܴv5��{"A(]`f�֡Ĩ������[跃Ǧ��\V�b��d�Y�I�=}Ť�cᇭ�� ;�#ϐR���`��B)I��+�gv�-���mNwpV뛃7Ǎ���<��������t���9/*=ϗǏq�1��୴�l�7�ױ;^�ܹ��ԫ́N�!�P�����Ro+��H�8 .f�{�+G�ӓ�5�r웩��8��N��1#������Hf+VLrs��\m�S�sy�}��Է�(>�'��k1�gj�.>�!�T�xj�<�\Gt��8�u�u.��g�U�i�[,�@��c��Ż�vm�-����-˓�m��靋��t��Fx��=�z��wah���VUEC��9eF�ȟb� f�VE�d�c$=�cc�b�Q��<�6���� ���1Y�+������P!C��D'�:�@�\�#$�N��m�$'�7Z�+�&������=Z��{i�'+ϔ��ɔ-a�齣I����	��;+�J&|4���|䥛��IiC��<oBI�5�D�c���g����2q�@��k�PX������R:��	{�L+�>��P��qTq�v���ޥN���ģ���N�ru�]�r�*W��r:��YD�qP��ib����;xr �I�n�����yq��Cz51�ч���Qڹ����U8�b{�a�Mc�p��yJ�ʹ43\�t3t[lC'�G:Ό�,v;;������6
�l�G6��-��t}�2�㖪����)KN�V����v�q2!f��ܳ)�z���䫋6���r��vћl!C��|�|>ҧvA��d#7�Z��9�6�~� ldA�˫�r�/d�Sz[zC8m�(��r�9l�+a��i����Y<�c���6v�X�%�1@��S�)�b���׋�Ƿ~�Q�JٰL��E��9:���]��k�g���b㋧#ڕ$.<�Fd�ޫw��2�^���m<4h�4U�#Р��MΡϜ����8gnn͹�sS�S�r	�R=!U�э�[^�9�hU�M���sVoQ�f��n�����x�fv��Ê�;���^�m��G�ڤ�+0 ��>;���a:n��n��#]���+q��l**|�绎���q�Jؓ:���Έ[xθl��Vs��m4H�>'�."�j6����)�������q�����o�7;-��^�H`��?��S�@���Þ� V���s8a�ຄ/r�=ɒ��pת�S�U�`Z��t�S*<�A#�6����ntͽ����n�����vHrոx�\Kl�_Nێ:�ٯ���ڝÈ�˘;���k����N��p��y���	�]���"��h�ޝu�y.ub�y������A+��tPg�wå��Fod�[Vn�5�����t��n�I@�puv֦ٻ]�8˭��X��0*$�����3\g�ӿ ;�s�!'��e���g��;�v%|Z��>�h8]��05��=���tn�;a��[��ň�p�;����ˑ��_ �``��.����;�<�r�B�w�hn��FS� ��ˮ\�2N�J�6���u��]��0^�/pB�j�;��7U�2�q��1�U�?��p[Z�@�}6��yW�/���ޘEz�a��۹����,����7�oa�M�WB��ӆͮ��h�e���e�a��sŸ�h8��΄��[�i�
�p"�I���8u3�~�7�j�e܂���((l����X��!1�q��sD&RT1c�/���W2��f�"<�{H\YNf�is3�.��u�`ٵ�h�}Q�{��d���H�T��+3n<ub;YʫǦ;�0�x)M����Bݚs�{U%���z��@�[{E�U���1:�k0n�S.;��O^���ո;�
nΗ����S/R&M���a/o.�f�m�w4�gf����Mf[iYw�Ig&蔍�֝�a������"���Bc.�����=ڕ�:+��HC{�=C&�ͳ��rl��d�v�6s\l
�
�V;@'OoK�âd}���4l�9J跶u͇A��B�r��nn�Co,4�ڊW@�R��d�n�c"��N��.��37V��=�p���P��6:tQ۫bt5!wc���x
��)�J�{���NR��'�Y����Z��KQ�u������i;�6�kYRMu��
�@����$K���n���� ��x4�� :]�T���f�<Qk�����P��Z�pk$��qN��٧}��6���lAE�Z��1ƎOܹ�2�`�� "+5b,=#쪆;����K�2d�&�!��5��N��[P�I�1�7"��l�7�\�d�b�:�D���H���ta5�gC�fӹRrӱsY��z�μp,�^ [�87n;�gg�]XLY7Q:��@5b�Mّw:��=V�;K��#⦰K�D\E��]4�Z�h�j5�od#/Wn��"�r��::N�/s~�D␜�kJ��u�2Ӻ7���7v-wu�>à�d�+;�;3s��9!�|[[ e"~:�t��Z����4�Ӵ᫖꩷��Z�&^��9R�t�q¥91I�5�5��L��j�Z�ݿsLjձK���z�f���y6����u켣��PY��(�Z�E���.�{����V�tͯ(ޤnN8#�Y&��P�!(���B]zw�#����u�&K�EY�E���\���*f���얌�Ϯ�'g}�=�]u�v,�f�{n�{�mǜw'qW�Թ�r�uRyd�.�i�[Uo&1ώ(Yϥ+��W����ux1�^-�O�"��˫���[�Z��4�����xKpt{�`�C266b�k��1\��}�Dv�LO�:8X�q�x˱�&h��7�۸xFU��3��3�2x��85d���ꊝ�C������iv�7�.ȓp�9!]"� ��t�d���T*˼�Z#s��R .v9�v��n>`Ƈ|upD��u�vv�!�1=�! pZn�:�V��T��K׬f�J�C6#��:��985�۬);;{U�Fv׽�7I�������U��p��b�Y����Z;8�l{��c�.ڱ5�yx9�ͫ���7�nd�1�\OKt �B��\B�o�\�1��V�4�a�0v4(/��(�u�ʡ=��`4�E5V�'q�:�1�fp�ᣙr8Ż�\�F<\l��`d�sy
uw���x��m[�隢�W��P�{N����� 7sj�>�N�>ӰF5�nD���6�sn)��X,CFu��$ba�u<׸f�I�5.ӕ�7f#�q�f�F�Z�+wom<�n�	�3XZ�����ɜ8�J!�����5�C.�k�@w[�2�gA��Y�V��^�����#w�̝���Ǐ�i�romI�_S�B��7uN�^Y��uw�FZ�jݵ�P�iy�����B���닩ޔ̈�I�H!δFXƞ��K�P�\�ǋ�oi�qىpA�Ţ#�̳K{���s�k8Q�����ؒ�t�.���� ��&v')���D
�ر�F۹Eɴ� �=d���C��W5f���ݓH����5V!��)�-�^��nGw��x�X���R��2���,qn�\���ҹ�R��}�К��������� �j5܁wlӴr�<���^�ʕ��S*S.@��qй!�-ɛ���L���5�h#����Q�B�Ͱ��]�	��׷n����o)��I�E�b�J{�ܓs8����^,���VmS��^NN�ͽ(�� �vƕ�1���yd�v9L�
���n��n�܍�h���̠	�pi\�[�0��E��L�a��fB��o.�;�wp�:;�I�4�k�Ϛ�G8�P��ʱ��Ȟ¤�f��D�㝎q��Ʉ�yf�:U���혝�ç���r�xCA�>�[O���Є�'�ɚ�A��&7�[0u	N�7${z��;�f>�1׋757���>±A�a��j��Yt\u^]�r�s�w�;@��>��(Bl�+�t�[��b���ӹ�6�j^���t��k� Ed�<����Ș�.k�^m���U���������#�c��0���9�����x8F:�9l�Ι@����$������-[��O������N�a���&P��e�3u���G9ݻ�����t���,�	|i��Z�]�5һ���n9����l֫��ӻ0��۹O]0�]ھ'�gI��ݔ9ڒ,;������dr�v�M�r����RR
e(:�귎t����4�q b�FTTU���PӸ�6��B*��k�ٯ���{;5����wc���u��:���s�; ��˄
Q���hz#�!��zg�{�o�
?t	.�(!�mXa�{�{���-|�Ǹ�e;�����b 1�	�����޹��5��L�;z��Dzl=�7{�vk�u�4<z9LA�ٌ�ذ�{��#;���l�/r= O�L��-�x�s��D��1����(2��v��ٴ�C"ձ�K��lu��G����9"�.{꺜}/\صi��:�Y��=�$�IQ�����r� ��G����FN�	�n�-��P���c63ڂNui�v!r껿5Î�[����^ow����ɺ��D���2P��Re�uc}�t��F�I�@���f���g7B��k=Ҽ=�!� qc������65��*#9g��&�{͹CٜY=�D�Ft�9�k�Z�7o%�0,=�rz^����1.բ�!�k�וжs�,nbg��`8���ε\t�ZJgF`��B�$b���,���[�7睺uc�8��D6MR�W���C�c��ξq\ad����J�Ű�X����������2ݹG=6��7�u���NR�*Z�oPv͹��L:[����I�l�!��ڛ�p�d� ��o.ź�]��aǇ7�L���q@��ڬ�%����@(��wb�Ǹk'^��ۃK��V�#��+J�+��`np8�����ݎ��t�qsۯ]�XDMu�k��ۡ�嗶"��`��1�jተ���ĉg�p����P�gs�[�ݮ��%4��Q+����U��xB���ݞ��X��<Za�Aw}�h>ۮr����D�6�}�n]�
�!��}��ᏼi����d�W��r���_^j;�$c��MH������[��-
���c�&�����DM���8+u�ݸ$�#1t��I&�'��柜{�wv�u��sԱk��$�{�;���� �O��vn#W�fʱ�2�m=����e��忼��ly���P�j�@W,�N���?-��/sԷţJ��hS]ݣ�^�;*��5��ifIǪWl\�9�?=�_ٳ��?g����z������P���JU�T�� �J(��.H
䠁M"	� �
	�� ��JD*��" R%(Ҫ�%(P�� !�(J(��� �(���d"�
�
d�d�
#@�4(R�� 4 	�� &J�d&B�d�9
�JP-(R�����4(H�d�d��@�@ ���*R%*"Њ"� d�!��IJ�RP�JĨ"���)J�P"9(	��"P�9*d")@�*P�!H*�B�J(�(��T�d (R�"% �J&H�������7���=�q�#���������iNfթ��u�
|�\���a�]~�x>N&�Ў$X�QvF�:,�l����輪���jX�[[���4���7����ݝ.Ŵ���1���|����w�zt��$�M=Ҵkfc�����7p}�'�fo��G[�o�oX���#�>��Pmw�_G�w�~ hUAE�������߯��~��K���P����	��.�L�4��]I�ĪUs&ŋ�i�/��=�^~H~>ۀ���g��g�V�˺���,p�w�x�'9o�O�E0�y���L����ø�B�����}�C窷��l�8oʔ���˲�^@+�J��9<n��i}ݲ���#��}��к���c��^�`��̰d�s5Y�^J�î��q����e�����;,�$�˞+٣�[~*����F�0���ߚ��{,ClK��g��Sԭ}�����������>��]�������s#��^r�0���.ݺ<z�KKQ����_�K*���y���d�gf��=/��ׅnwh��jd���2Ѻ}w;�ube�N�Ƃ��9�.�9��O�ȯ�*\�����@��W[��ܻ��@�������V��Rw�YZ��<'���2n/Y�^׎�^��^��i!,�?Q�ĩ��㮾�w����iە��
j�QW��<�_jՐ��/������=���7���㼧=���E�Ig��wr�8��Ht�,�����J�ݧ���=�{M�n�C �z{���r��^.�L{���)Ȱ8�ɨ����󺫷w�3+	y1
1rk�6JY��{�b�߼����޳��ף3�a{�v��1Þ�xq�=�n�u�yS�B�|z�o�o^m����>h�q�q�܄�����Wb�k�@�M�%�f��_P������N�a��>��zO�՛5ӡT���	}�bh�q���}�m����^�z!���䱿b"��T�N ɕe���,y�g��{�+�H�9�jt�(]W��O����"S�:����ù�ۃ�~��۷< �Qw��w*�oc'�7fl��"��ƴ�.�b���^�6���WH���4��s{�����佞��B��^�{��<��m�!����}�߶����x!<�o����/n����]7�9<s=_�.�����ܤ�=ɧ �#��(�v4�����s4�ףH�v�EӾ�/��Ԋ�}K�I/�NSK�6�4(�y������������5n��wS����f��E��x����L�5"�<��zl�ζ�+�[��1��{���0{�ٻ������;�Tu5��7q��n{t(l�ȉ��d���U��0�N�)�dm�u���)�w�O"��H�1��F߈F�3
����y��'���ҧܖ�~��V�u��\gۓ����nm��^]+�D���W�:�� �tw���_o�Q~�y���5�z���Ǐ@���w�&sL��˞��]���������AޣA�>�瞬{��x����>9��wk�}��J�T�Ոt��}��I�e(}劥�}`:�`>���V�=��T���S{������9^`��+�8�������i��[ď|6��$=ٗ��{�Jv������dX��g"!�,������z��vm��ì�h�wG�욲\h�x_p��Ks�;�z��w��K��!�H�/l˳������p<�h����{��F$U8n�^[�	��_�^��No��X2�VԦ,������6+�^��A�e��IdEA�B,����h��׌�����f���}�w�ogn�a�V�@'�dJ�v�5s��3�L�G���a7�O[£��0�<2燴�H�{��`��Q��n��]��^����1h�XLGp�ioL�K8o2(����������y�ۡ5�C����]]��|\��3ΒU��_nZ���Lo}�{>�h���u�,��a���\��/��罝���]\������٣���	��JU�C �Kpa��ˇ�k��X|���Sd/G�˫�s}��$q�䆛��^��}��Np��{Ö�.�^����X Ӆh�����Ho������\W &o�_l��rSt�{��+x�n����}7o g�%��}9=���c�����ݼ7�[;x�(=3��\��>��Y�G��g���g��̾�n����и��������p�~l��n�jņn�r*�����3���[ǣ�t�m��ӸO�-�Y�+vՂ��n����f�����8����� �t�{N0���4=�'�yh9*ٺ��:*6{��RƼ<@7_�-�xF?g��ܟ=�+�<�x��+vvA)s�tr�����L��]�&̡M��b� 7|���x�<���rY�vɫ��E��4��3���������;��v�3з���?$��8����<U>���d�'4�z#現Խ�^{GJA�7u@z�vǁ�#1�����z'�����ަ��wX/`^{�<\�#�}K�.�Low(7�x�^j�k�s��z��p�˽[��У��7���u�W&=@��yO$#��x�q��6`]��Ow�>�_V�����^����}�řr�E,�ty���׼�	ǃ۶�qO�T�G<�|��n7���5��y�Q�q�V,h�n���\��O~F���"2�d3���#�Ԧ��B�@ns�%gд��U��z�����e���!�F/�u�w܃ F�����xvӳ��O�w>�{�����Q�D�ܹ�U���^�	C�`ʃ�M����"��x��_��ཎ3:��v���{a�{��#�;S`|�%nl6=#z�{�n��������tև��^y�t�0i�r�C�}����S$ʆ��|��s�jp`���ly7y�C��=m��X/��{���1��Qv��zgN����*����EqC4�[�Z$�n<����}��rؼ��r��_g�<��x��!�0�ë[|E��i�z����zt[�������|�#��:u~�Ó�z^��n���N�+ e�n-g����^x�\s���5X~낌��ݵc��ǽ�VZZ$�k�|�§u�vl/�N�n87��VwM汢ǋF�
�]���w�$���<���:�����	\�2�(�{����nO8�NP�����|�0Aͥ�b\�<����oypk��{�M�-n5�,�oz���3u�r����[�`�tsB�'��Q�+��ݍ�w��o�/�ӏ���G�m�U9r#�d	_g�Mo����4C�5��c��/.���	�G�kUo�^~��W9�w�b�d�c���{AŸ{Ĵ�t<��Cn7�$�ߗ'��~͍��,�ݠ�S�ܴi������8<��X��k���n�$�G�s������r@/G �f�v�xk���z��F�=��V��Gw$Sټ��Yx���m^}�w���a��;)�}��y��x�ƽ�1��y��Z���fLx+N����z�y6�ss���$��]��e5�ڠ�i�eNI�p�3�ݞ����pB=��/�G���ݍ�����l��U[�\\�ͣa{�<��	ޏ.¦�䗴�%繯|��ٱ{ڻ}���"n����c3Fzr�3	w�n��;G˱
x}�P{������eK�����{�6��]0��O�f]��4��ryGL��3���_I�&��]�[���4=���R1�=Z6��u�z3\^�^˗�؏�>�D&^W^gtw$Cާfa�j�Gv���|�7���'J�Q;n����)=�Ꙟ���=^5|�xRw}{�b�)-%,��4�Z:x�ծ�^����&�:��$�j�A'溦��`�W}��WB��p�M��whs��1շ;O$�o��A�� D�S�Z�����kw�yD����ʞp��w}���yT�����}�#��r�^����b��<6g=��w�t�Ǘ��e��//e=�x{��s�G�+���qc�[�2=~�ob��z�q�>5�-g����;�HFHŹ�#�;q�� ��+��D2����;5{یZ�>�\ �[zY�w�R���k8z�p�N��v��Bh�e���ݾ^-����� %���w8���9R;&�7 �u���Y�"�I��RH\Z5k���~"����Ts�N��ލ���7��㫋�>y�J�9�L/G5zu��i��w|��=ѓ���%��c9����fT"�Z�xoP7�9�}N�{�C͌�"Z���2�>82N8�x�^�q_���]o���}�w9����v���h�w�սFƹ���y�����9����Zxip�F���Ɓ��e�E;�j���r"��׽�<���zG��s��8��<ўGh��ru��{7��^�%��~:9m}��,鵏2��s�8'J�k;�����ykupg�E����x�����x� In��ߍ��/#6p�w.ܞ�u�K�!��ۢe����%�?W��^�����p=�a���s��҅I�1�]��$�����y=�M�ˋ�6�e4��Ug��r/oUW^�X'�8$Hh�_|_'��2zE�(}��������</_3�D�C"6:<W�/���0K�9C#����K��F�k`��ά�npo�<�^a������܅�����g�Ro=�)
%�4;K���?�%%������{�<�]�M������}�1?V�����΋7����y,�[��S8�����>��fX6L
s���4�T��M����(N'�ńR�0y�U�L�q�t�3B��1�9���M�������C���݁o)�-�V�d��C������7��o��(ӭk�K�L����P+gE�M��+�$tS o�ɝ�Q�]ᾞ��|�����-��>��)��V��x'bg;{�6��L)�b�ë/���l����ܗ�z�,���}��{�*&�Fb��d:�{�h�3c�I�u^��M�ݾ�X� èju��;&G��U�7ęzA�^�۞�=����bul��1���1;{A���h8�f�R�^yq���q�-���律�c�;쐝Λ�x_��T��٥a�|� ������s�\�O�Co�CW��/V�띜5t~mw�fOw3���ތosE佗&?Ӻ���=���VO��t�ּMEv����ic�;�\�닗�a�:S���=�Ǿ�ހ��3�<w����e��l�v{��w�O��s�i�.Ws�`rb�>����������ٿژ������9��5�z�=���<r���B>�2D�2��X�^��p��er��|0���8�{��b��GD�'�.��{�,T�4o��W��ޙ�p���QJ%t�ݝەv"sk"��|��h��6���z��w��$�wPi����[(o꽄�6\����q1��=K5.�8|�{.x[�I��-�t��V$�t��L��l�HY��O�̖���2���=�/��^m�v���@)):`����7�ȳ���-n:�V�_�_��qzv���5Ӎ߇���y��a�/o����yywt�3��h�������N�zS0��>��Ѽ3�<_$;�)=wړ9�bȁ����8�s������x�Fz��2��8j#B��ض�}�$�6P�ĩ̻�'���;��yu���}���^�'m�`g��O�Z�u�7�2��M9Aő0��UN1<LK0� .l;@E�X}Nu�A�_�x����J'�ݼb��G�o�ĸ �<[Ր��/t2�p�}�#�\�f�{�ī�we�ә8�������@B0�Vm�����U泵�؛�ڼ�����m;Q��=9�{m�ozG�;�!z9�^�v��ш����Wj�x=і�Nw�e6�u3�~����׸����w���^ЯѶ���F}�vwa�U�+v�\O�>Y�{��H����������얤����:
��|/N<��Ы���tTPU�`f��,n�����;���{ۚ�{x��կl�(����������:�s�t�`c����y�w+�y<�b��=����wGB J��:q��;��6���O�2��A�����`ǩ����<�׫�g�g@�A)�:r����}�FQ7���&�=DON��?nMGx/M�{}ʻ��aM^/|�7��k!��f\�7��eFV��~{��<��<#�����<��Z7���5� �7�<�{����W�=w���0��̱J�Ȝ�e6��=���j�u寘��W�x�X��ӵ4G�Rf�tE���ݶD���m�C;����b��p独p=A�D�{l��c�>^�r�����8P��=�(���QI_h���ɯ�3��<a���Dơ���jDZ�jE��C��K]��QɎ����n��n�J03^?w��&����{൞e3�8���#kҽ�,^�to���tt�(�%�k�Q�!)�a�������.{ɩ�>��o0��1nw,�Tڇ�B4���A��'�(�i�I}��9Fs����7�B�bs�uC�ã�~�ӻ�&���u��?"v����Ϣ�9�\�`��>]���7�v�>�_�kF�������:����{�-m����g�H������+�=Z���y�z׏Y����Ywq�ّ4`}����/w�7Oi�6À�/e�-3^�[�������w�{��V�ᚧ���g�P�1VUm����:�N�/�ܻ'k�7�����'�[��nv���"�s�s��D��}}WI���\���ݾ��|W�܏�&H9bmOa��7��k�üxA�C�=�j�\���{B�V��g�*�np�j^V�y�S�۳��^�j8����+/d���Eϼ�{g��W�rSxY�g��a5�<�Q�;�U\;ß��n4Wu<G��ތ`�}�z�o��{{���R���g�oe��s�t�xO�7���w���Aݹ�C�l&�/?hܘ=���o��v&�.!��ɟ1�k"s!V��VX˅�ѣ1b��+Kd�7m�B_/���~�����~��������_�E~��~��~�~��~o�������z�^�����kKC�Rr��:e��,su{D���7]��nN�^��.%5Ʈ63����.Տ�\Gnl��,�R
��ţG@�:�s:gS�Wiv�  gsM��C	uB��0-��X�m&.�$�M�oe�� �v-,�.e:n9�/nܱ�j�Sn97Q!��;=�i���۩z���Mɚ��Y�x�6Gۭ�p\�J��;T,��s�ll�;�g��Zm�m�4���F�C��ݷ���C���3w]�1���0�)��wn�)�e��0�jCF6:]6��Se�!).yfW@Ϋhi��d.ֆ����^A��S�nx�l����pv�p*���v��\�g%qV�v �F�a�B	�]H���Mk�tJx=9C[�� x2�C��"���Ps�Y6^P";r�Y띲v�a�̧$hu�����9,�`��u�d�0P�N�s�ь�P�x.v�M��8��m�Qp�����n���{SG,Z�����dN�N���v�ֻz����
Eg�F�`�T+��i��A�`޼����Ǹ�׮�ڒw��W6}�.,�WgD�&��uSci�Rv;r�n�H@U�q��c!��)i��u8����D�x�^c�v�B]a�Yv�a[��](!���u�=v'g���K�l$�լK)�cLa��J��+�W]�u���sF�]����WULl��C'W^�����E�q��h���c��2���g���1ǡ��XtF�b�Gq���Y��`k��ri�ÎV�դ�`��p�^x.�2�s4s� y�6�և���x,�ǀ�;���	�Ƿ;G�!-�qmW費x�����^��K��ie�്�w;�����r������v8:厱�����6mDpfl՚�ma)��Z����/l#ya��OK�|��d��=�:z9����x�X����6iSʘ��i��wi���n��:6�@������z���=���!�N{mvsV,6�8�îj��(���,Uk�� �d#���ehmL$%R`� F\���L�C�Y����l+Q�,Q��,��l3/1(����l2��6	h�A�խ�C����G�
���l1��h_V7/]z�L)� ƺ�֔a�0QN8)���3uQO6q�s�֕c���y]r�n1xƺ�W�0��@$���:�Q���kv�q�9���<�-������[��^یL����.J�M<b�\�;�#�<����L�u瘽�w==��Ǎ']<7����Bi�pNл�Vx�W3�c��s����脮��[ֵ��[p���8#!j��z�n���<���=n�v=�ץ1*��r�m����%��Mk� �lihh2�ILk\z:�9�t=�X{p�3�v6x�xI�|����ms
'��n��x��Л�f8�vb��nN�g�.Ǫ��g���5Z��9��1lvs,x�y�G�v�C�O#śΓ�ڕ�y��d���>��s��gt�Ր�K�$(B[�S3K1X�E�m��mj�ma�p���i-�luv��:�pS�%�X�v	�^{�q��G2r^آP�n׎�;[�l�W=�Z��8s�A�;K���I�����CYC��\9��r�<us�w%��{;��\�rqp��J���2�/��p���4�7d`t���<t�+�ֹ��۫/u��\I�tf�8mWdP�I@�g;Ţ���8��a⸹ݺ�z�#�S�=#v�W[�B鳞=�(����P�=sɚv����5�p���R�����:��^�q�
�y�B�[.^����޴#t͜$����T5��ƍ�����e.M6�R�i̸�,Ը��U�+NWH&i��k;�S\�@��to��nbై�*�1e�[�xў4islsЛ����V�#��Ǎۄ��F�MӷbN49s�]�󒓨¨%��!,f4���������;v1�񞮳��2�)f*)��.���I�q��Q�>�yC��x��۰�o;{E���܄q���5���S68�:ۧy��-ˡ�:�E�<]���/$��j�8�:�E�4XM�t�Z렦�Jˀ�(��s����ua�����z�K��v�+q��qOc벵�;c��2�r�]0,6xl˦��F�����h�hV��D�����>�pm�G,\<��j��'���.ݒ�w8}�n��k�m<pv����U��9#[�-�[�\u���U'^v���<!Z� h�����ǈ{O<s�^�z��m;�����SX��4�A:�[��Hq�Z���:��F����������͍vษ�s����a�vLl��^���ۡ%�2J�,�ZM6�#.\�vۑ1d�hSs��R����Ol�Z�-��V��>��z�[q��p��ŗ��Ͱm�!��OI�g��e��l�<pͭҜ����6&��	�Y�U)ś��&ғmu�y�1i��(룳��܅�g{]���cc��糽d��2'Tq⃗�������準���U�1V͸�=�<<�nm���]˫����ظ{m�yh9��@�oF8%���N��¾��f����\����j���۝���.�C�9�_c���j��\�u��M�Zpq����]�Cm�O�73�i���](��K�+ʻJp��16�6:8�<d�ݣ7�U�i(잼`y�OE����;���Y��y�]^�y��NBS Jm셠�v:Qz��u��+c�Dv���m�y�{Om��k���]؅��8��\S�������Pkv��5�`p��[f�MZ��@�[Qem�-,v%��L2�I�]\r�<M�7R�\Zt���1ac�%0ˬb�����N{6M�	�MfV �*�h����ż�6�)0��Qm).�]]��6����c^r;�[l���cz�Ϭ4=۠M�p�r�ڻp�lָ������/6���v��[�x3��9�����r�^Gv.\�}I�=d<�u���pu��PdG��3�M��q��gs;-��/:�v7&v�R�]=���Ղ�r�9L��]�H0�f���6d���U9��\�$��/]��2ֽjrT�/����×v�d�r�٩H�^�:s�{{U�:�Ϋ8k�ݺ(�]Dg�P/�����g����c�gҙ*�'�������-�sn�%�\Fc�,ŏ��6��t��(�^-խ*qq4�u�k>�E0ZP��50gT����S�ph�c�ޞ�x���Aq�!
�(�A3sCsfl�Ԯ�����WB�S@lh�Kw1�(P�ֻh$Ղ�Cn=7l�y^k�`�|��n-=��m�u��M69��n�|��ӽ��b�K;��3����p��<ví�h���
��Y;R���i��LA�V؛$5�u(� t�[p��F�V�� �7<��m�	�u����N��ɓg\G�2$q��bz�v��:0��I��=�ֈ�F-��mLd��a�	ɽ��mnW�\ʙ����[�h�D��c^|�ᴧa����<\���������^.��&�#mԚ股*�$��Úe�K��B� I����b;�m�lz)��2��
X����ǌk)�������q u�R�q�to-k ���<8���r��A8������6;v�nOa'�f�7i��Z��\ć�b�.x2�˺���zƹ���m�1�"U�.I��F�R�n8����/#��b�CN�=���֭���gk���k���=��[�=r� j���㓭��GMv�p��Z��E�<d�z�� �)��UB8fWR�P4�m*�m��"���z��T�'mt�lr��oI�(i����k��y������"g��Dzzy��������Hh�U�#��n�nwe��|a�0�5����u�N�X�9R���; �h�,v�Cx�.��t�j��ZE��ki���&tuR�ԍ���I�`����uqr�U��y�7[X7��]ٍ��.�qȲ�停@'{�9s;	w�`�8�XR��:��P�#v[�.@d,j���4f�ƣ�%M�I��"�nR�lg��l�vn��;/sW]�b"FٓZ�R7A�R�e[H�� a5��Vh2ܒ��ι�v�&�ڼ]�����X������������5r��u�o��s�9.ػe�\��en�m�R�lqf�����v��=�J�Yܳ�$.��m�U��:����[�h����.��5"p�SC���v�țt'�'z��1�mq���>�n��n4(���8ӇA�kmXF��^a�m��lJL��4��B�[3���r�gا^�T�]����pj����P�d�t���f��O�	�s ��l���nn#���ƻqV^�L�셂�����������<�����W:������ӻn�`U���ּ��FP���+�j6�N;�C\M���t�Xh�N�N�8�Qs]p�i�p�2���K۷]-s���v��ŻU���ͼjv}�@u�9]����v�)7�u��sӼ FKB�q���7BW4�]�G:���ݠ,�MuU�&Et'];�5H��n���V;�U���5�K�������n�wc7#�Z,��C�����ڎ�6n�<�]7g���m��ŉw����NTI��	鱉�u҅͡�4AU�B�S�d+l�hAѡ.���cR�̓�4ڸ�c��^�qW3���5V�7:�i47Q]uʷi��V��ͫ�=W:�W5�ٻT檪�$�kk��5����9�,z�WL��V\�у����M��N���#:�-���V\O������wn� xRAHq��)?3�=��#lٴ�p=�8{F�&n�Ve��7s���7j�-���i�vd[��j]��r�n�7b�=�f:!�Ͷ�tD��ڳ���:�m98��v\M��m%��N��q�c[nF�L,ì��p�4�-�kY;lδ�m�c3޷y)�+gvpJFh��6����q�'"طm���D��4��2�6ӂ���%�8��gf��\3S���ҹ�Y��Hp9)Nt��"s�"�C�GY�,';-�D�&݉p9m��p�u�kj�e6�I�!��'�^��2�P�	�6��n�B��H�r ��"D��y�C�ݙ	R*N�:���d�Ok'H<�ӎ#�IYPIȊ�ɷ=s��ٛo�u�M�]�<�n#t^�ϋ�'���ǃc��ނ`Pp뜙��"/4�pb�h-5ŭ\�-���������8*㱬uj6��ON������v��c��=��E�l��م�M=��
,]{v�nZZ[37i�֮y�v+8뢣�p�[c�j3)�����ɴ�f]��� ���0,�
㳣�s�b����{���k�W��uМl��ض�]�7�;Eu���p�}Y��᥸��XF�KS��2Y�'v-ó�۱�`Ӹ��段��g�n���0p�v Z�T�B���4�3�`�kVU�3\�v&��;�u;rD�۝j�`�x�7*�u�8���#�d���iBhL�K��ؘT�q�+'��&�uۡ���W�'V�v�cY��i��ĉ���b%���TSw;�u�Hŷv��8�P�%ܸj��	��ˊPc,�tI�v��'>�]үR�0��"�籽�]';�<��]4cq��G�2tJB��6t)Ɔ#a:-�(���랚.=��g��6�Y9����jv��\�׷�ԝu��u���;r!�w�=t�c���Ò6��׌m��`ó̜��	���Z�yIn��(mc Зlؒ���7a}���Q�������X�>V��u����Ɵ3�#��PORN�gG|�Q��v�6GkU�q��b�h$=������ۃ���PC`�u�aۓ�& [�M�-F�Qᶄ���j�hTyz�p�j0z��2�Ň��U�G����z��u�&�Zu���X�J[�y��BѮ�(M�[à��狊�kν{g�؛2�F���v�GE>0q�1�`�-B�}���o�-D�J��u͉�hs�;=��t���'M4��Sa�[�.Ǜ��6�ZT�������E��y�k�^�����k�tRi.^�2�,4��9�\�\HK3Y��s@XkThU`P�e�`�J�е%!P[ʥ$Q)iT�8<e�m��$���
[ ���n9�x�d�6�ƣa`�R��6�R��Q���Xq�%����e��
#e𖑠�mV-h��#jV�����
���e`[XU�e�	Z,���T�+R����JZ�6	b�U��)�
���-c(2ӿ���/��a�6�୯	3�q� �L�8pgfVc*�x�X�ժ<I�� ���k@�r�����UxƼ<x�.��"�k��AO��{5� g+\A�5�uL�!MBY�N��ew���|Ȉ��k�o ��[�i0��j��"I˫���?�g�}���@�$����Ү�ɦ����w�����|O�����N޽�|��^A�2۳�K<d@�ʂm	��/�wxlk�$A�֢�L:��nB}�� ���x���F��vX�{�
��hsh�pL�5i��::��눅�7e�`lۋ�lm]��~K�ͫ�ql�^K���I�ǀA�'vތ�UO��(��Y�s/ @$����4��u�:`��g$B�|0H�Mhû�^����')wy�<o�c���'�u���k=�Gm����yz��?{��>9�"�~�YaK{��-w���Σ��_��0O^A9��Czwʳz�1�`�̤ԁb���� ���� >���u��*;�f�����I�^��5ⲃ��A��0�׍תB8��z����9��Dx�9;:׏�S�0�m�?���n� �N�'��`�wO��Ŷ�)���cs@'��[тH���1����}�����]�F��U^X<�2���/X��S�����x�]v0;f��Uˬ�Ϸ�!�	���qU�Q�	'ӳ� ˊ�-d���`����`{�P���%����;H��p|s^���v���x�X��`A ��ǣ��[q�Ef�Sk�hCZB8�0N\3����|0A ����H b�Tg�ɟ����VYK�+u�>2���P��C ٿ�7�'�^h�u�o��=}�����|��Y��j!h��챼�lm9�ܺg$`ux1�L&
�y��`�֣ ���k�0,\�0v$�>;�����m� ��Q�I ��� $�em�0�)N�`�����
e��"�b����A��B{؁7���Z�3���-���D�$����I[p ��d^c.j�"|A��	�ZN95%�&4��m�u�o\��L0���{�����_�n�Z1Gu��=vum���؃�I��ۏH�ûKD���+u���J
/ &0�`L�3��^��$Z�,FMkh����l���ĒL��W�Ȓ�{��񑬴O���/`�K��LΉ� ��	��q��8ib0�mz�W�$�� �[!��#��ٓ�p��cn-�B`��{��.�׀�g�@3�W{	$M��=��#$�E{G�J����n1��K��,a$�_�
��Q��m=NU�	����G���U�>W��a�F�7��������Ӏ���K0~~i�#me���`mKek�ܒ'7 @$U�@�I9m���elf==�󍱮J%L3�?k��Lz�۷�k��٣�l�X4r�!�nM�<��b����w���E/� ג5��#��	m����C��<)���o�y�����ǀ}|��KF�'J�]�P�Ъ�=���6�߄	˭�7���A�okA
,&&D����38A�w�UμH5ki@$D]��zv�N���H̭���P	^���	��;L�m1��tcg[!���Uk��H$]5Ҁg�ȃ[[�w��%�����+I�'���`���9 ��Z	�gf��&nh̍�pH}Ɂ��v��*3c�7�6����uK�َ~�,R�Od�����������c�QlC��5�'Wu��V��gQŶP��YaQY4����mK&����X�Q��&��כ0cs�)�m��⛝[ˋ�	��5����������lrʅ4��4�+!��A��uz��>9:��:K�1r�E�Zڅ�6�{A� �R��:Hx��lm���Z�$�r��5�����f���5��X=��xa�Wocq��-M�2a��2�0�y[����5��+����k���ͅ�5�곭>2M�)�l�͎��<�X`j%��o+S�Bb����P�3}���=��6�k����	y ��ڀI �f�������c�O� v�-A�x�"�� �w��Q{0 ��$��3Z�ŝ�y��m��o����q���\S]yB��:aKJ jѠ�~�.� ��k� i���P�g����w��I�m� �Z��y�B�#��w(;���뿲�]�ױpFڜP �F�lA�n͛�9�fs�PHmk��}���[��I����ƍ�Āg2���<XvX��>�g� �^*��<gv�@5<�"��|�%��_�>Ksu��4e���E��c�f��,�a�0-Ӈ/1u��1Y?|��#�3�7��@3�qă9���gEA���Zњ�0�FecǦ�%˺fr႐��������vw�K���1,q��|
��,`��~���L��d��2��^xL2���VHz�9L�a�Fj�C�5N%��*�b��k]n/A#6�gv�@ �Vc�-T�چ� ��V�w�;�@7!����/∥��p�ڸ�d�Aܛq���x����g��X4,�T��w*��������	큆I��# G�'q��lepm�"��	�}��/�&�S;��������$P����Ղ���dFDx��^���@')��4����D�8z�	3c�Q�u3��:yx�e�o��j:�Os�����	�WG?V�΋x�v�i�A��x� �Hk6ڃ����k[���I�ˏB��cEӧg	����N�7Q�DnB8��,�mz	&�-�@#m�����j���|�݁�q��N�3;��L���<FһP'�|�0�+��S.
�x*��B���7���ݹ��.ǳ���7ϯᝉ��7�X�]w�a��H�|�i�)QMU�0�۸�I�׳ ���Ҳ��ňN��nF�C*���+Ɂ� N��< ���-��ߐʜ�U��w,�HNHg���`������\��RN͵P �}�of	����n	���uF]Iae��,]�jC�����ݽ1'��nwO.�ݧ=[���'t�,+	ē��������x$j��� �;:�D����[������I9���{^���E��;̛h؂Qk�����$�lk��HU�ڀO������^23a��V���f�^���\_�!kG�����w�Vb�O�3�o �X�gKFB��Ŗ�L��Ǆ�b�AٝN�S%���A�ၻ,r���v�x�8�H&sn<��"��Y�r.VMoRh0��r���OT�j�U�P,^0�Ū?\X�/\��;:��3�J���^b0�YUA\Eh'ӭ��F�wvH]�. ��DI��x�Ƨ���e��贬�#Ĝɸ&s�<b�Y ��*��:3JV�q#��8�уu�Ʊ�`�q$�ݯ)6�k4�vVT1��/���݋�y'$'��h� �I���@ �;�D�F�Sy����z%��Ѥ*|�ß�L ��2t����{���;� �;8�	$N���R[�CiD#��:�˹(&L��"�����o
3UE�Ci��S� ��͸H
Z=�]NS�HM�3n �ּ�i*���[I$U]ǣ�꽶��u�2`���g�?���m"V��X$��`|����0�NN�>ݿ �~o �r��AU�*�Sm��O.��mH�W�+���4���`���o��S�HJ�J=�nt�?����YJZ��ۛ�߿a�"�;�>���@� ф)�ϣ�kxݞ��\s���эoX|#�c	�<�˞��N���qs��� 0v�T<�ty�S[�H��MfGeSj4��m�bR�������5�c]����*m��7����f��b#��Ӕ�v�z����!�b��nx܅Ьl�B:Cv����p�-��WW#�q����u{FFh{r�,9�9g1N�:���K�5��iZ���t@����f�M�����%����MI%�.���%�9w$]�/ ���$��i��(5H��2(����wv�G�pk�p��v'���Lް����)1�����*lZp���	�^[8�|c�Z��۾�¨�#4@ݑ�Y�hB��);�(7��Cd��M�a$y��$��b49���@�ˁ �}���kX1�)��\n�L�k:���SE�ěh��H-�h�Aʝ�{���@$3l��|��ad�r��A	^c@$����I	Xs-Ez��U@�4�SzElz*�2s\w��x�.<��f��7���u5O/�H��j�)��xix����׷�4���?5������/�> ;����Y�q!~WmpJ����+H;�����Dz	��E��kg00ͱ3�5���ƚ�1�4�Vy}F��͎� >M�~��dt�����{�0�~���L��\�il�Vc�M:��Nm7��V��@;��T՗8�W5��"�۔�8!�:�q<S@$�Q{j�rpk��9&�r��r+`A�"	n��Q���z��:���L� ��dG���q�J�:�t�P�� c�����o&pC���-��A��q�B�g1�"�V�j�Z �r3@9[. ��������8����(�T�75���c���״��z
�gڅj9�ۊ�V���y?T�ك�(!�,�h� �v*�<H9[. �����q��=���?>����oH%jpf@;�Ix����`��;aD��� �LfDA#+f
���h�QY�xQ����8�ہ1c�[`d��:�s��]=������>�t�����׬��vv�jE҄ڝ"�US��x�]S�As݋\N�<ϟ�ٻ��s[~�ޏPI����H�$�L�l�{Ӧ�+v{�w=~�&/-9����YygO�>��`�5NE��%���jE���;R��oC<r���L��jȸyK��ɖ��<r�Ȩ��y�q���g�Հ��ʧ��q���p�}�zcʠ>��=�����s�Q�������wV7T�<ǽ��<��o�g�V�E��.��U<��ڴ		~��x�֫t�s��s�ʤ��zﮊ#᧞<1�l�˷,��J��o<�w�͗��8���w�{�o}�I��<;��c�0�o����7��p���Ol��'��@��9�-��b�~�jE��g�A/�"�[��"���}�N�:�F�.�V�8��v����Q�y]�n��"N���=����3��M�rH�"�<���3����1���ֲ_l�ok��i�qw;����Ͼ�ټ��rx-6Rh��F�,S��BwE[N_�4����S�/���3��"�g��h�:�j�����b�o:��{S������U����(˹��7ܦvqe�냪��n�=7ٷ痴p���NQEǸd�e�Y��"��f� �A�v<�	;�a>쎭��Y��{�A½i�X�^<*�c�=q�.����w���}U�_LW�݅>уoyw=+/{��Wp�q^D �F��p����Бk7:@�{��^����f�ހ��7�b�v��,=�Z��Ő�3b>�y�!�'{U�����\F�rYÿ'9�aFbaIK��������f��N��(N{[c��t�#��rD�r�h%#�JF� �7^v�G ����{!��3��N�p���'Bbv�]�h�"�;n�����˲�mnIBp�Č�e���x��lܙd���b�$�
�j,J۷vV۲.۳n�'}���ΰ�m�ח�xs�Zwb z��Fy�{3��b/�y}�}2�ג�z�m��,�Cw�z̶�����]��s�ñ��<�O>'���idY�6�>�J5�Q�o{QA'��$睋mׯ^�tv^���#���@�=���9�m^���/	�q͔�μ�����F6�R(�-	yc9�/�y^���e����d�N-NC�-א��6|�z̵�o,g��Z�y�z6�.׽{�8��{8x��=��C[D���s�g[���˄��:�F��%���o������b���ӕ9�VeńE�{n���8͵��	�d&Ja�w�[jC�qJ�$��{っ��9u�Wz��I���/C�Ȳ �y�b=9}[zw���ހ�w 2R���mG$�)I�9'��8d�q��q#f���#�&�$֜؃�@G�����>�����HI����#Br"�O���Iǚ��%)L�����6�@��iapu�41�k��r �[�{�!̥<�'��8B\��"{��Ꮔ��@i���#8o�ϟw�Y�|����\i6��[�f��m�n��Wv�i1
��E~���?� J�f��wg9co8�RK�$�d�����iH�#!3�7��v���s�r��Ns|�n�9����=����iJ%��qd賰wb�� H�Xݰ��}��c�}槹Y�/4���#���I��>0$2N��|p4<�d8I��6}�c!��@��"�7c/�4C%���n>��$��:���g,Y�'h�
9&��\p��Jfb��	�{y�\��`#��|>X��DK7J��>���2p� ��m{�<$��{q�ᏼ	�����D0w���<H�&G�{�2��׺����J]d�&����<�Ҕ����{�v���B(��$:������Y]&ZH�sA��3��Om��%�pEw�p�ݯ-�;|�>s�-\����<�;Z�%��C��Q���TZm^o���<�E�>ι�DW��D!�&��.����|-�G��\s���S�@d.B�W! ��@>>l�lΠ=�ཾ���NI]u�[��@�2A�Yαx	}#"���s�{2��/�	��$��Γ:,g��A���U�[pٮ�S�cmY�
�#v�r��g�����l���	�o�����R��;�]���	��!����׸�2lÐ��{y`y8�[���˒�@Dz������	E5:N�%��#�=�����̜ːd'��޷�m��/z:���M�ۯx}��1���2=����G�$�b�S�]����@�@��Ym�Pu�F��O�~C55Ƅ;���d��y����� �\�{μÙy��]�؇ Bv_��F�۞�ʫG��w��#�	��~%� 2rC2=�:��$��^���r��`f�𲏇KF@ �"�f5㸇�]C���^�$x4����	��&Ѵ�F��ֱe)� Gȍ���>��q���GUh�U��K�`C�:�~d���֯6���x��b��hyd��Y�qy$�\�/y>��>�/9�-��5��v��)p�g�x�e)JR��9�d<9�+L��]��|�̆D�8Ј���)�r��qOA�*N)�e����v)�C�w��.����6g���Ȟ-X4�=��Mo�rӇ�rf훹����e��8��u�ә�ו��͊ˁ
��(��BRPnLo<cPn�n����t�Ott�0�pZ �R�h^�].H:`��)�����J�1�]��Vs�z����]���w][����횃O�j�̔�8�@Yj�]1��4�Rny�Vݰ�����E���Zi��\ܶ�8Mښ�nW��+'n�H��2]jl<�gS.�8�4v�Z�.^,�C�&�dF�-kE����Љ4��(\�^$��?O�{�.4ro�o�5�=�<�A���u��q2�$9&����;C̈�
r���:��xa���竆>��dNHaw�y���go�Q#Y�1f-��.𲏄o>G��>�^H{������)�m3����ݰ����Fy��k�R�H�]��|A�K�d�	�����3]�9��0�Q�Jj$�D��A�z��x�"#��ANe�� �=�[���;S�d����.��}5%�����G���@Y)G]�^b�┥a���|G%䅄_�=�3S\hC�Il�Y#�{�1�ۗ6ɹ�� A��#�$D-�$��$�rL�Z�G!�!ő��ݐ�x;^���8�:��=�}�H\�W��</7b	�9��3DxQG�6c�Kx$���y�xv6�1�G� H�qtp��=�p|!�v/O��S�NG~k����\�%�2y�d1�<����$޻�3���'��:�n���5m��GS�a"���\Z�6�
Yt�.�!7݉�΂v�=��Զp9$�\�%��]��y'yJA��Cq�%�𒏇�"�D������<�=��&B�!2M{���;G2G`��(Nػ�<$� �:n�A #�������f�4�^]C�Ǝ��~�w��-� ��y����%I��/m�۸�B{@���Ci^���%��{����Bto����}i]GK�xu����{u����/0d�)I�����!�2\�|���6�����QT�j�]�#�d�zH�<8!0H�uj׆�Y�ܔ��t���N�ל�s����2�Ex�B>
be��6��m����y)I�v�|�oR�C���6���^�֫m�0�"]à�$z��	�a{�O�u��7:�˨2R�nv��N��y� $���3^�ƹ���R����3�0}��wt��Ҟ��M G�(x�<���X�2p��z��)���B�KgrY#���6�H���2\�{μ�8�ݼ��|��#�|�׋�4Òm��s��$�d�O��8�^B���J=�:�=�"O���)�7�����33["�w*�56�n��������{g/!ֺ屬���$m���Y��"{��Q��h���-)��k���+�L�$��6ӵr�D��G�,��E��x�}�����0�����$�[s7�"�	y'��������yTcR�EK�{��Y�l�������Ba޷��v��%(�y׸�/8�a	�m���<�0H�W�E��
�M��g.�y������k'�Xؗh�Y�8rK�˒aI3�{�ͽ�:��b����w�)��N8��`!9r�s�O��=�|
�jS&"��o�=���{T�o��ԧ�!�j�_���?����}o�o��>�:�h}�!�L�	����� 2rC���������$k3�Y�y<9
>� 3�|����甥)Bu��w��D&@lÑ��F{��{�s�d�Iֽ߾#�`LzF6DNOo������N<\1��'����V�val��o�܏R�o�q�!�'�d�A�u���|=�S`�d;��'� B#� ��2�xID&Y)�a�׸�<═�aZ���<����ƪ�]d��r�b���qnE�cj�]���4�����"�`��:�!96�'�{�.�̝�`�W�$q 6��1y��� �\�w�y�,'0c.JRcֽ�S��2C:��Y�<m�ݼ���^�������rR�;μ�z@"O���W��ზgtȘ�
:fC$�F)��
cn����]�{��Y{ϒ�$��M�ڮ�<�I��3UJB���u�(7�"���k�T�̳z[̏�+/��C$A &�[̪Y8֘WI$��z�>�PIWsܩ	-�7��.᜺t�Ъt<ڏd���W�����I)�PIY�r�$�q���Ki4k!�q8�s�2�t#J��"� ��p�RǍڻ5`�Л��'�Kic���G��%�]�����A�$���S)_�MH%|�X�2�xU����K$�7�>��ʭ�f�j���S) ��ǹR<�f`����>��*z����>N����]H߄����&��=ў�=���;�7��Hv�Z�13b�]�|�=��K^��'��kNO�W�^J�Z�Y�Ivta�HX94�����m?b�%�^���`D�灕��û����/}��nkS�e9Qq��\c��3/$���2�$I���"QA/z���m���CU�(;�4F'	�L�̉���>d��	u��J%$}PtD�,��ީܕXI*�{�(�H�s�+Mh���t�rK��%��+Օ���nS������$�Yyf|��H.��^�`��_��I�l�̢gբo�"]ø,�'�T�ř����W�]-'�u������k�I��q,��w1�τ��������Ow���qJH�:{&53ݲ�W8�L�d�vɢ]p���mع��c��m��wN�Ҍ� �����Ă���S�}�\�Z�Z�r�Ž�������#�;��lz籯�Mʘ�-���ugv���6K��Ggss��w4�����\�bԲ�nw,nm½r�n�>�W�au�81ٖ��㦬p�v������.uz\�3�㍈��zNzvSÏ7��I=�si���gճ����r�rL����ˊ��[�<ns�]���a�����L9���~�������A�t��v�Sl"IF7[6�����a8轭ۜSu>���:S���hNy��vL��w�~d��B.���y�Q��7��`�I%@I'ܚ�˻�n�%q��%�T��K�;#�̜NQ-��]��%��%#�U�E�R�昦I$��S)/$zڹL��>���+k����V :��2���wi��ë� �~d����|��3^�Z9�@@P	 �y�c>Z�E$�[�)����!3�2&��L6��CƇ�X�	\�Z�%,fo$�^�I2�U|��S����]�R���z�"R�ưE�S�^L�.�ٖ�PJ���C '��U[)�_o�I�%L��$��b�J$���r�>���'����j	����]�yv��[4�<bm�7Z���=A�i�l,�z������h����e��^I%�ՒRH%��p���B�I�˱�T�(��k�)�ȗ��r�f,C��j�d�G���\��EMqW7N=�kF�4"��iE�h��7#ִeE�6��6,N]�1�-�U3�zk�U��m�ܸ�o���SǻF]�����1��=�����4ʹI"Wc�)�^K��R�H��
���OK޴���ի��L��dY����U�vCJI%׭p�$�=)Z&�r���n$�I]�j�(���p���`T�̘�,�J
L�>Gj�fȼy���Я3Rٔ(�I$���T��I ��G�'�����ij	^�H'��Pg��h��K������=���	r���&����re����4B�Iy,�k�>@$��:�e�ٮd��̍��A��hf)&θ��5"��t!�� јs#[]	Y�`K	�'4��b\�.�F�E�]�/Ǽ�Kd�)$�渖H$�����){�ƫ�3=�ݪw�S(��;�o?J&��;��8fyu<Sl�O�i����x�nĵR�	$Q���R��(�ζ�(�aW�o/,��w[��R�s�A�vEb�;U(�k��C�k�L��H���9��������4|���-,y�����=۝��&'×_+&\�}VO�N�ɷօ�s�a$����}-�3'/�:�����=��L�|� ��ϐ%�%�����d�t�"�:t����^O!_���/$���Ȑ�$�\��� $�*׮@G��Yוf<����R+ߞQFֹ��w��ly��;\Պ�:��
��Wz�2@wC�I�m{m2�&d���( t�vcv��j�`p�s�Z穨��b޹�i�1����u��ǛO>0�_~yg�<.��V���u��z�U崁)�Kկ\�BG�zx*��j2���k�i@$K��{�p���r��%�^�3M�Ԇ���,���N��S���	,�vd���ƒg�(j�~PL��О�j��P��n	!�&��3��8L�(�x��D�%���҂I#��5�ٚw(���y}cH߻��g薙E$��z�"W"����%��������|��I-Oy��ID�L'�i��� �I׬S) �j� ������e*����NU/Ov����*�<�d����+�=�8��.�?�W����<����w��s�}�
Da�=|N��p�nn|�J�A��f���͸�9�����I�:t��[-=-)$���Hw����C�[�I)i�i����޵L���j손��9�ƠJ,�e�$C�/e�~���lq;�pw;X�/[v��.�ݱ�r�4u�%Q��w��h�x������y�H��j�iI/$�kvK|�vgo5�j\��%�9mZ�R��(2�\�ft��
9F�	���I�p��ST�)y"Vk�)��(W7d�2��K�!x��㥠媱�E�t^L���fC($NZ�tJ	0YF�VKT��ZI$���A$�.�lInI�rL�3��B�˚&�=t`d���0��$�V�!���@%�ْ�AB��Ə3����&1�$��|�>����C�̙y��Y+ne�	 ���i��u���W䫛iA<��m�i�^\����P=t����==�:||||zt�����[�\.�ww�����8e��*�k Hڧ_�;�4Ʒ��C����*���wh�э筘�b�k��:�Z��w{ϱ��S��Z�i�;�|�h jm7�C�P��[�g��{7]����L潍�5���m\���n����BB{����
g?1���桴ڽ��i�<G�c:{Bv��9���=��G4�����x��w���q}��ӷ����ۊ}p�j[#KP9U����������3�|O��;��+p�9��|��V�ޝ��y�ʅ����f�|�z��E_�����Nݽ�RZ�)'���������;���Y�k>�ۑ���}����ʫo�Hz�H�b�银�g�M�^S,�����~�s����T�g�e�1w��gx��� �_��T�
�����ȓ9�Ӽ|܆��De�E�'��v�G~�@Ogx��J/s�[}�B����'���p%���2��єv~n�Ｏ�\�9��vD����92{ɟ6wvvlk����5y�paW o�,�}�L?y�z����L�3�{�������o��n���1}�V����;�Uc�h���M��4��@�ܠ�nnz(�Ƚ��ED>!*^�a*�;����ت"��H^	�|�-'�t��u>�V4t�,}���|}�0������=�	�g���G˯�1��)���'��ڊ��G�|f�Y�<1g?r�����5���{��=�:=&�ޔ\�=�Ǐ��9��Ww��)��nso���?z��jھg�t3�'.����a��o���{ώ�T���%ke[l�FY�ju��7�	�c�PE�m�v-����:͛K<��w��#��v�I�m�����@�}����^^K�Ѿ�E�N�!�N4�&�mӳ����ēm��ǵ_zܧ�E'B��n<߃;��E��9(�y۞�o���|�t���iI���qE[��q�em{ݝ�$�H��u�����y�[K��y��.NY��ט�gA�p۬��X�nZs�bBE[�H�����A���II�yמ^���q���\r�}��rN9��GA���3D��Y�(sn�:v�ܧ=����̲�{w�[ol�'���ȤfR�㨊�rH�Bs��#;'-���	%��'}=����o}��U��Τ��1[��6SJ��
��t7E��;�C����t�k���,����5B�L䰯&���G�� ��V�륶�tc�66��d]-x݇����<`��lt���9۲�LR�b�D�n�(0�KHW*�syLG[���/w�-���c!�!���=���]h^�X�6zm��7>޶�u�я=tW��s�m��;v�:��\�m��L�kR�[P�p�^8�ظ-��|<k=�S'h��ۦ���8�w�d0K��.����\���}�3�ӎ�g�w,Хt�����%���h�.�n� s��2-P���X8��oD܇v���cm�x���7Q��Y�Z�4X{=ļ7GZwb��qu3(ˬ�;�6��C3Z���6{(�ArV1f�v��,iI�+,8�[FغꑍЉ��,@�86��8Վ�C7����n�:���uZ��Spw�ty�^6�4)]�;��������Z=tp�l�F��-�L1�T�	e��XJ�H�8���m�aK(k�笾�^Ӆ��!���Co[��7��hWu�/ ��J� 
#n����l���GP	Z��;ϵ�wW6�q���=��\��޹K� җY�D]%hC-�h�59�շ�(g���zzy���ϱ՞�4�j���w	��n�gx��d���jy�V,p:c����f���{q��vy��Y\u���:��uu�n<zC<��I������#cˡe���g:�z�' ������l:en��cˍWn�9ۘvq���Ԭ�69Ý�b��ݷj�b�a1&p���]fx���h�mi8=q�y���S��h�@tN3�c�沮�1g�u�\��*qQ��ϞN���
����\=�
N��p(��Z��'h�z��<�[{g�͘{R����ƗU��`��&�共�֎�V��*5Gk��.�3�ҭ�]Q�9�9$��C��Y�-�1m&��Bǆ�C8��"E�뢵v|��7G�����̍	c��b��p�L����g[=�u��=f�k���k��������kg0%{=�r�ktٛ\�܏c��Pn6���,i#u�Y��ɰA���w�;s�É�b�l�Fx�sV�nҤ��]�y)�!���G1�]��m�s"準ɪ�ߎ�|��f/k�M�U��ۣ�`:ꗙ8����5�;Zg��wR�����V�3[��?����ݯ;dB%\�"C�A$9���|��ջÐl��|�+M��J�&��[vZR@�]�̘��&S6v��$�/M>�UqgW;�m�a����[��ςH-l�i�W�G��v���T�R��/H�+���07r��\��$O,�h �H$ ^��'���|�RI]��iH�൲���9 �֌`�L�t	{6�s\ѳa�6�9���R�%�$�
��J+��F�������>q䗧)�Q3��7�BD0p��;Ъ]t�J �s�Zk)�����j	/oS��O����L��Hֵr�M��\�by�~��s��D����ӳ���\g�z�s�m�-�Kfi��S+�%ѻD�̫�u;��$�3C�[1������DA%��A��IW=r��B�9�ތ<��!��JI$���<Җ�Ήb��رy�K%���($���j8��c��v|������Fnv�˗$���� ��C���,�ͣXb�Ɨ�\�V�T-�Mʁ4*)j�u'�1=(m{F��xF���B��T������v���̓s�)$�򯞾R%kC�N�Gz+"vT>��Z��LɁ.Έ($�����dY*欖�A.��C�;�l���ī��̓[�)�RIV�r�>oU�
���y�:L�~vحǛ����w�PI�iL�RHn=j�	 �w6B�le�s����}[�O�l	�v�/���PI ��\#��y��Z�$���I2���z�"QI.�|�!-�����=}�|��~��u��f�!�WsiK��K]�����9�z#���Iv��%��K�����,38N�$�R��"�j��I).�l�K]�=�ZR�.�*��S(�����A��*CS̈b��g5�2A)z�H��d&�]�)^Ie�r�dQ|�*BH%�]���N�V�3ҿJB=�M�NI	�b��%��RI.�k�d$�����e������Cі�f	���{z
#�SN5�U�Aev� ��}�����<q���oN�D��K<�P�4�HO�Cj����Y���=� �F��^W�_)�����T��Zz�fL�&w �d��ڙ	G5�_'-�Is����$�U��-!)�2�1� %�tv+h��I
�� Ǫ��i��Sfd,�3�K�$�](��F�H��w%Z��I&knX�JI���&�B}/s���Q%j@f�u��O;J�g����׌u��Rː���s��}�� ɘ��{�t�L�� �J�Z�C$�	!��jg�gʭ|f�����zz��@%w�r��-�5�B�p��;Ъ��S) �o������2RI%��r�&B�~��Qx'i�4t��Pr}�L���H0b��P
1ṁH$H�֧�R�I&h�u������sT�I��u��"I�磒��&��fN�3�RO�Ձ��f��@��y"{e�%�Ey �E�� I.��Q��-#}��K��-��	�*1'7�;`�Wu~q�bO�|��&&|w����1�U���Dd�\*ZKኇ�[4��� ��{���ډ?e[ܩH4��3;8%��(%w>�$�K�l�i�Y3W*s�D_6 ����RH�����K�u�Z��6�k�c��|::�_��=V����,��F��#ۭ$a�0�VݶE�qb[K�ן,���˦r�+�[0�2��Ko��RH���jd$�pR���d���{��z�2M�fR�{Z�I�;^/D��
�i����a0󦛧"�"Y�U�fR^Iym�Z�(��1=bi�S����T��{zM`r���L��]��1f	2�n�� y�͘ku�����oSF�&�H.��2���2V�je!#���{S�	�2uT��u�q�c�2/	�%�ي�IV�je"z��w�ㅃ���}^) �^%H��'j���y�	>�҂d%׭q,�dvk��v���I���	���m�>�W�[|�*R ��e�!�.]4ߞ�#-�D�5����J�ӕ���(F ��gv�3нޏƌ	��,Xe)0ƪ%Y����O���?������|Ǖ��ؚ�0�`��8�sz�����o8ˌ��$�Zsf"��҆2��e�6���x� �7<��6�#t �*��ڲ1����s�6ݺd�-`��Ԗ���@�:��8�|1�R�97$�g����f�t>F6�a���)��Ľ�"���9�G8������ݲv g�v�8���WY�*�E�T�s6x��r��֛�xq���ķn#������28iF��7P�{���=�r��g �`�c�)��	%��r�I;|�
R��~%Y�Sq��Aܰ�1L�I�l�"RzD�&v]0t���t�lϙ �46��9��\�0�ҒD���RL��_\I�$�MwF�8����{�JX���L�u��d�ZvCJ�H�:�%$��̕C�3c��_1n��^5���$���I�mɭ���w)޼*��y�"u>TONn�K���4��I�ؒL��[��\d�Fj���	����C��rr� �b�fB^���$�	^7Z�MI㨎�ԭɠ^�L��	uּIy$�߭L����ͨ;��A%��!x�K���;n��\��lqGK'��t��<���v��t�-���3�b���I��'�) ��ۭx��A.��Q)8�w����,A_<J�E��tI��yFՂ���g �4h&ǾS)$�nΦ:KC$��bu�&�io2��X���F���-�!�S(|�|��{ܦ����ߟ�:����_⑚݄$K3�u����ٛIh�S�P��B�
E�Af��II+��$�L��ǯ�)+�8�0a�hn��Җ�4q�:΃�L�k�]]/2D���V)@I$�V����%��a^���*�$�I����)R�k^�� �|��^�=�ڵa��dA����Qy�0b@`�lz�3䗔y�7c�*P;'o^��4i%�_TI&sd��仔�B��T��H%x����X^f��P����	EVD	W�9�p�J)%�޹L�qU�smFo߾�f�����d���`��g���ӝ��^i�Ae��ı�uF�w�}<��[�_}�z��d�^J񫔉K�/%�����c�2�;��5md��
|�I*׬M�˞	�43;,�T��O(���Ŧ����K��E2I�^�L���	u�rey�V��1���L��j�$�[z�vwpY3�X)2��9H��I.��Q) ��>����;kt��)$Z�Ϫ���u��W�VS7ǽ�g�J'��X����`���]Q�k�8�z|��1I�3"C���m$d��E�� ��>���D"�)T{מ��W��|��=j�EK���JWci2�t��b]ª�������g�:۬�5�J@$�J۫�e%���]O���UU䊦�W�Hj�GRA���$���\�e�BD��\#3�t������Jq�T�H����@���*BM��E�7v�`���Db\&��Ŵ��\3%[q�7a5�rj�d4������~����`�kv���=��{�2�D�����$C���HI�#�.Nƛ�3�O<ʙEy ���JB��)O���0Ϊ�}湖I%o�gc�u�ضR�D�SecL�Jڞ�O�'\�i�g������h	)�I�q�y5����o^�������q �S������]d���-��Q^Insܩ@$#I%��	vwpY0pX+6�_1]���<�oJ�Q~�$�J��� $��ǹR�(-��@G���$Ip��o��f������"k�!���_�X����:;Ju̶�?^5Ai	hl`�M�jh�3P�jlTւA�|�μτ�ER�� A(i��(Z����~�2�τ�f�t��b]ª����g̐H�����f�|g
�}<��Mo��RA*�k�)$��~��X� �k�ù�{�Q�~Ƹ�饃��XR��D�4�4�1���6�y�CS�&�Is~y��<��[�u���[-Ҁ��I%Y��1�f	 ��~�2�WpD��d��[t�6��(����+�H��Z�\8p�S=
��mKK�ȷ~ނ��n��ke(�Kw�$�D���L��q�c��Q��JVJ�[8.`�� �OA"@�n�"R	 ��z�4�  �rҼ�2]{q&BI%����B�n�'�	Nŋ=U$��@�zN��Xiz�	���>H�	,��S)��W���][s���)!W�d$�u6���&&Sc��z��A&W����Xc����u$Aw=r�g�%�}m>���d�u=�|�o�4{���G�~oW�K�f�
p?�n��;���ӵy8��ʱ�����N}nr>G3��+�~u{}7;ޱ�D9G%YS��3��� {�{�����s��s���v����D��1�Tiݺh���y�<���&;3��`[Fù��&B�ѭ��h5��ZI���B�4���2k���Is�he�v������n�睐��nN��)��\�>���8�qd�x��q����!PmfZ9M�@Mؗ���^[)��X�\Ӭ�u���v9n6�6��\V��>g�K��$�f���t��{L��������ˋu��6���ڭ�B�ڌ����e���?S��똗p����ɟ2K��.ƽR���L�͑m'|�/M`G^�N=����f�c�(<g��I��:�/�1��ޡW
7�������}h�y$B��ԓ!$����QI]�ou;�q�u<�^��Z�8p�=
��mL�J<���!��ʕA��Zu��5;՚�$J�|�>�PIyk_[H���:Y�p\�3:��O��@mgA�|�&�$K��h2^I
l�i&R]m�-s4�wd�v�Ƒ)t�6ƀHp�3��vs�$�ZۉuW鬖T�*l��Ζ�	 ^2�|%��n�>i�+��1������Ush:��۱^�ڬ;�k�u����dzHz��Ī=w���%k4�=�?}�����nW��HJ��,KGE��U�V�[ncA2Is_[L�V!-�t�U.�,e#�ꛞ{���q�Nk��~�ׅSeW�f���5�)��/oA�>}����-\���$��i����&��uMH\����iY�v}�����@@H- �"�ȠP��w�����9�fg�k㽃��3H}�->I��Qd�r��%/j��&Q.K�^L��1���U���I%Ej
fG�u��ϐ�6�)!��rҒ��At����g�T��m���q�Sert%��CD��Kmm�! �\���G7ݬ݆�J�;Ze!�m1L����>fuE�uF;���	Zݶ�JZ�^P��h3<�I2�g5¿%�b�t��>�ǲP}h$�ؕ�1�`��� ��!�\�5��İm�̆8Ch�Ĳw%��p�c�K�b��x$�k�䔗^�Ĳ% ��c����n�Ӭ�S<������q�_̙$3��T�%�ڨ`d� M�ڦRI��c2v��^�yI �ƸR�	 ��O�]�Z`)���o+�z=�)c�1v%�+�]P� K$�K��ԉI$���W����W����{=��W�����l;Z�<��6���_9��ܧ�e}������|s����a:�ƻ�|�y�i��{٫}�r�R<������h��ػ�����~'r�ح��<^����#��gl��V�kq�[�n��oQ�8��sY'BN�컸���E�#6�3�7�VYD��q
!�AHٳW#�پ��{�ݼ�ܻ��!�9#��=����W���O�a^:
��x�^��"���P�4L�
�y���~�,��xq����)uz�����`~�y� ta$Xy�ý�)��4�1^�p�n�{���k�ó�%4���iɋ|��˒��{|5���}��H�{l/�"X��i�{��)���6t���|6��J�v��9����;���H3��e��
��#Ė�-��b��7�:�Oz��8����	�,�������s�i��iΞ�\$v��w�����c��(��n������n{��a��Gg�ӥ��J05��^��3'ۗ��oi�7|x1���,P�q����l7�?E��zM�0��ۺ���ɜ��`��w���u����;t5A���9؁�����o=�r9o���n����bn�r�j��&��Hk���G�٧�{!��a+������d�����x����[o�_�Ѿ�f�W'���ˣujnm�fv^�EQCu�8����D�Q���[<j����wax���R�*�%Y<�E&�7.G�,�6���݈��qwj��{)!g]5_"�fxO(Y7��q	���!�'l
õ'*� ô�b��qY�ɼpjطo���uQ_^�E�r�D��)��t�t��q��k.�!Î@[gw$E���a�!9'm�smA�I'6�H���;�Υ8(�:9L�8��:�����)����i;���B).:�q.t�"S�8��(:#�!�@R[[��mm��$ ���$����V�G�%��D9�ݚI�f��Nq��Qq�ĉ�q�tW��w�a���(J;��o/q#��7Y�ն��<�y�k�r88�[u�y�b��d���T�@�V�T�D)A)$��8㽹��32C_�@HH�_��jei��$�D�t�x3�N˘V�jR��N]����x$	I$�k��$�z�}�zr�ǳ~�30�ۉ$���;�D��4tV*��P�3jk�y��l���n�S31&BH$�����GU�4�Sc�t~��g���țXQٮ@ҫa5�(�.F���%�FX��Gk�&��re������t.O��wW���̄�H%��j��.k�i�%\��c��mc�f$�>I��j�I8ƀ(�v`��'Ʈ�Ғ���Gu�?[ƤJI��R��I ��A3�+It����4o� ^�a,���Ұ���Ӱ��_���a y-la�orZ�z8�I U�֧ҊI���e!V&ؖ���v%�*����y�p;m��$�UmT��I$�[�)�$�Kæ�$�}�J�~b�)�<&^����	��Oy����#��<�}�{]KL�{^�7mZV��r-5n��f7}����5U��Ѥ�d~�����R� ЁB�@PH��H��̜�=߿s��3����c36Q.�^I=����H%u�<JX�+G:��.#���ϛ"e"R�{�"T�0�f��tI>��s���^�f"�gL�.d��ێ�V)�s�md�L���=p�\��+�f89@�A��K$�N�~�t]H�!$W�]>i%�s��(n���4$i�(���E$��z�"Rk�f������ԀTo<XI��ս�ȓP��3�R�y���h���Ht�D�e)���<�{��6�AH�sIK�X�v`���'��@D����x���I&ȡS�L\ku��H�5r�g�!ӝd$�馴\Սu��v��{��s�מ��h ^o�6ZRD���d$�AvOH�Zs���6$o�L��-RL9ˢ�K�UG���y��	u�@�S��{���ǭ��释S) ��OdI��Grz�>>>Mw��������^j�6���M�
�[=�~8��{9+��À^<s���=�i�
C��Ya�V0��Y1y7%�PC>FR ��r
fq�� |B S�0@
�(P�HD*QH �s�^휛�p�[9�+�9�#h5N����c���.12og�ü!�fH��C��gRuÊ�m�Xū��큒�����M�Q&��ʵhf]�e�X�^#l	d���5�+s��� �Hg=b�p�	Lk6�m��-�]T��ݪ�F��l��Q�1�9�U���t�{q��^C�ڋOc�waK��_l�k\�tFGeyn%͛��9����Qv�]מ�k��sY�ܶ�ϗt��U�(p�t���D���̊-�K8E��%��2W�y�2��x��	���s3��o�r��O<�e#�؂LϮ5h��ؗ%ܒ�Şv�Y)%-Q�z��b�����)"zw��Gq������F˱��4�R���3qw.��|�� Ӷ�>Iy �W�ԦQ(�71ol��JC�Б(\��� ����2��@��'z�V4�Qo-��e�	4�tHd�I%�ǮS>I$��z�-��qΡ�a�Lat��O<ʐ@�K[NX1g$�Rd&��R%$�K��%�I-��u8��;8O��*R>E�R=(�$�c�)���%�Gf�S��2di9H�݊f~5�sʥ{v�@�h��M���.m�IC5����>��,Ļ��]X�2$��[mX��RI$|��W)�����,v]"��}�L�$c֩�ƴk"�y�A��K��T����H��R(�d1eժh��3�U�#�"��nF���z�������v��p��������~�k�O�[�PYw���x�>F� �[9>����R;4\'@4�ψ�z�"���
�
d�h(V��J@)hR�)�
J�h�;�n��M�����6��D�$J�_c��	���&Us>uGCn�y�1p��ؗ%ܔ�����jǙ�%���%#�
�;$s�dɝ�%W8������Q$�5r�I���7gE:$�w��[����[������c��f���z�+��j#�/$�ۡ�W����d$��J�W��� !8v`����65t��PK��bY.l7n�� ���>	����O���IvS��K�sM��X-��:�X�I9.���]���P�#{j.r��R�;��0�۬\��ٍ�]w$�Pz���$��j��J#�Rۧ�D߉�FB-��\����-ҊIv��})
�F��%�1.�UP]Z�2���U�Z.�u�\����X��e"Pۧ�RA(��9�gmu�D�7JB�h�E3��y2��l�JI%YM�,���� ��zd2���a�P�^��1\,٨�̱3PmҳC!E+�Ӯ�q��5���_�b%��K��2��&���b�g�{�S��}�g�/��� �D
D1!CBҁ��#@ȩH�@ �x	��i�$Ao=|�J+�}t�B����Xd�]�JOB�˚f��.[oXD]4N�d%R��J�I �����D]��x젊87y;$K�~ᾟ�8,���������	D�v�L�qf7&i�I��S)"���*BI ��Ƒ~��:��soGU�-��9G���g�É���h��ŖL��Fo�'S(^������>���%��a�Sߟ�v��($�J�b| A%�ۍ HH�i����N�M����ΉD�e?J� ���ߺ춵��/�}�Ǿ�=�E��)��
���٧�R�H���Fʟ$�Z��	�q���vm���,��QЩvE�1.�UR�֙�I$噍"=,�@$����"�)��F$J�[,L����ƟJZ�F�(��,�$L���;�p�/ئIuY��WJ� � �IS^�L��G���x��MV�v�g�ޒ;�B�������˥{ߜW��h|�����yd�rt!J�˳�sgD�3ͬ���������wI��yǾ��9�~{�<ly��~%P� � � {�=�{Qԗ���Z_��69|03�'@���Ъ�扶��M�O�a�z.1�Gc��^�I�Yu/)������I���f̤��sx�O�&�8%&=��N�����М�]�X,�*��a,K�L�O|?-���v$���az�F<��ۍR�I ��y�2��g��v�2�5�rz�y�K�<�-� g���v.��{�ݤ���҂W�3��0��܊�$�̋��RL���^qA2�],�)��-�V�F-M�vf%�9%��>M�f=>�O[e�i@$��D@~0-1�Wc�Z�ɠ�����"QA#��JD��a:싆b]������E���Xs��K����D�fl��S>I$����X"���0�s�o��&}+�`�E�.�$��'a�o�$���@��b�6q��{b��K�cLϒA#\�jD��-��ko�� �/Or��B+M�2j5<fC䲈��L��a���������{���m�x�q^4����L��i~��yٰ̫w�w��-	�����YZ2����٘Y�� ��"�- �s�?w�patƭ��7B�6�[�1ԩ�(yv7q���T\{��uCj19���U:G
p3d��3p���X����{)6��=p�X.H1��)�Zƛ1�^#���q��
����m�u�!a˸�m=�#,��og�0���F��r�zlz|7�s�kA�F���+/<����pN'���,4�{�w��ϊ	s5jy��Q�o�F:�<-��s�a׍�H%�3"�T�gN�?����]�rK8d����.��)%�`ͽf	&E-�������s�h����8�2��W{fRO��ڙ�;2 �g3>X^�f1[X�r�Cݚ����y=�D��f�6fBH$�k�����-�S���]!�g��B�Q��Ļ$�U@$��r�^J�VÙ$;f�4h�j�,�גI ��,ȔP�f���������W�]���IAY��y!W���(;Ce�Iy(�{���dp�t=$J]}�.$�k�b��}2��o�q��p�]85T���ϡ���y�+ұ��T}����G��I7\�L��)m�H�+m�Kو��̾��W �C�zW���4m��3�n$t,�bu��,�[�@����C6��}������V�y��a�|�$��u��|�Im�H�	-k鋘���C]y>�I�J(%��a�$)�h�.Θ"�'�U~n��)$��[R�E�G�.�{���E�_��E��9vvz��{�Z���7W���{�������� ���X��A�N��}�㞼獸7���A�JD�\���R�Ix$��kd��2^I/���G6%��|����͜`�O�ͮ�;��A�fV����I^v@�) ��Pǋ�ʧ��s�	/Z��y	$���"R�L�a��vIު��g=��p%��V��I����� �}�$��2�:$�q�8��V��ޭ5䗱lܹ2r�r�������H$O^=�g	�̬�wi'7!%����Gq���T?9��B����F���p��ʴ=m8�ul[&�s�,"�l��Y�����'<�;'�Ӄ;�Od˙	$�� L�A%��je-�
��U^�����	%��"e/W��|������%���RX-Y�1�_m9���K����z�D�H$��~�>�RBcU.���<��I�=��t]���G�*�H�17��M$��>^j��V�N��\���H�c��o�1-����ʟ.��`���l�?H�����%�u}�����1r�uUM��X��.�;fp����"�aS]q��_����/9`�]����v�ͩ;3����^UK_L���c&#aڮ9\M �D�2���HW?Z�1�3%k�������O5��=f�S��[5r ϧ�4���N�N�vln�iAW��&=[	������Xp���ºzkƩ$���|�2��Tv�B[�\B��'�\.,�LYK�l�DIn6ގ.�
���Ź���b�T"0�Yi��7m���0d�A`t��v�2�	u�\���T��^R���s�x�f,ȔRF���7�:�:p��pj�،�If����8��n=��I%��fe"W�[*�y�I'q��	{�R���a%�.K�(<K�g�RK�a���BI/$�ыR�MK�㼒$�E����^��r��zӸY�8,�QzzZ)Iu�oh�{�)/%Wϲ��$Mۇ��+�u�b� �}	�~k;�p�eSU|�3e������r0��.b����)�j�a;�zt����9.w�o��n���דz�.��*k����o�Đ � �� 	��ĐO�ř�A��'f��!��J��s"	x�b���N�Ol\B��Q�o=Fڙ�I$9vܹ'�R��~�>��"r5_�EL�)���3�b�ww�a>��=;�+���z�m.)m�ܬ�A���r���+���;$�^����v(���{q"H���PL+�a��E���Q'Om��I�ivrŘ�rK�&Sc���NWP�Ldd�l��$�\��^B@��߱L��]فC���/�ĥ�s��̙8L�85T��lȄ�H%�ي}(RI�k�ʊػ���J	���ˇ�$�Im�b��w�	d��]�A��]-at˸�I:r�0BI����RI��L�ם��z($�GT�����{�Qb�'��^�ߕ�M�	 �n�iN4[�qs*�ڸ^I:{�rg�%͝�"Uy0�]��Ux�������Ο_ޝ=���f��[omw��`Z�{�V��K�1�ک����^*���X��N�<J��Z:������[y�kfw�]S��پɜ�6��};cc�nM���]�ɷ��w���X�f�Z[Ǭ��y�G˞������ܼ����ĸ	o�!��vA��7�)Ssq�C���>�­��w�����Օ覟v��L�I}�忔N���O㸧���Ǟ�w�7�/��|5��;�sL�Ͱ��^�������nI��t�Ɩv�G��C�/J���};*�Ν��љ��ӈ�W7cwzV}�_,����=��F�rW�#Y�9�#����
{���`���l�o��C�N�Ո�u�VI�R����Ьc��o���ph%�~��{�{���I�d���ҽ��h�v����Z�~�۵�bߙ��~�a���ӹS��! ���y������M���N��~F{&��� �k�ŉ9/z���ߦ��t�o�{K^o�4��x����O��z�y�YwY�210)ܴ���� �B�p� ��B�LaY;i�Hx<U���5��|�ǽJ󕳷�L[��ou\���&���<��.{�y=޽�#O1E�0R����T*�s��5T3c2�^�qZ��������{�YL���h6�>%n]8 �۽;�����`��8}���vpu'�b˞7�ֱfZx��W�ys'$���t�)Q��V�@a
�u��㜰���G�{ ��_�w���ޣz�����=<���o���wQ���1��+�\ ����fA9�O��:Bȶ\h��K��-���㥝��?2�̢�8:����n$Ią�A��H�>ՑPW�v8IG�V�qI"J�Y\A_o;ם�rr�۳��*s�����JH;mq����@�M�w��FZRQK���v�ʳ����)"8H?An@I8>�j9�rJ�tRE~,芑�H㐄��H��5� N�*f�H�9%}�r��:$(�8�-�̄NE�@�\�����8������*f*6}w���#3��߭����mu�Km�n���`��ƞ���I�e5ҘӞ7^�k���{�lԼB��(�聜��GW��QɮL�e��Gb��H��0k�\�b&��cF��2m�y��s��68�&̋L�wi��V��e1�!r�f,���i����X���Ω�=�OP⶛"!xE*� [tH��]���6Nk�i�I䕕��k�ͬʧ.M��*&��{��*����0�Wch�����N�PuǱ,7,�\���Za��N����K����؝ծә���a�|7gU�ޕf9m�[y��y�]�#95u�vD�m��:�N��x�0�5�v�Hk����R/Eq���Q���uNt������Q����n�t��.��ې���9 A8;quv&�,Ɓ��β�v�����&�f��K�+����,�ik�se..qZ�q�A���y7� ^G��rI�X2��A��ݲF���kq�z �]�B�^3��<��F�.�#m�.b�VlM	ds8��k�'��5:���O�ţ�(D̛O]=q.��{1����rN.������g���^\�I`wR���.k4v�J6@F�nQ��p�P��S;0Q�`�gK��r-Ь��)^4�i�]U:ٌ$��:Vi���jʹ�h�F٬B����Ƽj�..]�ݖbE��5�8"G[�pf��6XJg4�
���5����r{��+�5bt�8I�&�Ni�nj2V �t��cJ�,n]�M4H���x�>�w�.��ۛ���̓c{m6��ݭՠ�5`�X�H�2m���bK4�`� ݎ91�s[%��7<�G���q6��j�A�Rm�C8^�uv�][E�q5N�سX�Ӷ; nx��+�:�n������y���I�m׎7by�ݠ���m�rM������M�������ص����4IKkzP�"FtA��l�ɖz�Rj�����]-D�SbjjsJ��iv�6�,���0@)@;��a����d�`v1�6Ƅ������5��
�-B<���㶎�4�kvű��ʄ�H���1zd9���m�甁��Ѧ�D;=�7�'.�tl��uvwU����b晳��n�=
/��;kX8��k��e�0�D1l�Z]��Cvz�s�X-��@0�k����G���Gs�����Ua*ܼ��j�X�M����k5V��˻�ź�7k�;�^صݻNkn:�8�1.RLh�F���^{��e��v%w��˙�U�n4�K�$��|�2�W:��U��{�y	�6f4���N�vIު�e�m�I�T�.��̝����I*k�i���<�m�QA-=շ}�Z��#�<�o(���3"�������Ͼ=�x����<���7a���~���^I.k�n���!���>���������Q�A��'�e3f��6g��p�mL�A��Im�i���HR��}�5�Q�o~H���)R���Y;7��(<�K�ƴO�'M�D��/C7�>UK^PI	j�i�fo$udSL��IZ��y�X�N�v{ҡ����������@̀Q�>���1�Ƀ6�ͱ�H�s�R.�ؒ����ǅi���{<����֟H	�1)gL��H$�ut������"X�U��i�i�	��S) �v�ff8!��L�1=2"[���t�۫�a�z/���� �������Qy�����4�Z`�h��8����-�-~�|=��ʱ�0��w�<ve�5R���ES^��<=� {U��h?x$���~�2A%k��\�cFWk�{'�koa�R�L`f��:tS�N�T�v�ʔA*=[	�I�L�u�T8lu�g�I%��&}(���Z�ZR�L�ӲN��
��٭\d�e�)mL�ӇBD�S�,�Ixe�t��$��k�-�c3vp��ӈ�d����7$7��;Lz��N��c) �c^&����z��=�x�3!%䗷Z�Z}�fd�sf�����$��q���)܇w�A�d�3��kp�\�64jD�u��<i��k)6�����'�N���
ǒ釳�KmVĺA$�Ϙ�@I7;Va1��	�W]dJ$�*�i�Hw�����ا%��^�ڸz�"R+��	YOr�wf��ǔ�'�V�O�0fAo>b�2o)�`��EOod�S��e4�v�vy�ߝ�����ƃ!$���\�j��_^�R�3���GO��ѧ�����݊d��o��m�,hj�zdw�fì�<���z�V^I��-�dĩr�j{�����}�I�.�[)$���1�ȿue�kC�E;$�w`$��y
�������J�UćI"P��ƒI�-΋6�0�N���{�/;�T��*2���3�);�X"!O�k��2^K�^�)�D�������$��OK��k�)�������[���9�����/�B@6A��&�6�i#p�]�N5��n�T���ڑ2ʚ=|�y������_���:f|�$��l�2��A$7:,̭�Pz��7���oG5䴄�H.��R%!�l�43�7��L��a�T�����S1*�'ΉIZ�Ɖ"Og=���L|ŷ+wZ
燾�9q���/?�s�"��'�N	{�ֺ��D�%Y�r��S|2�z����2���ts<?5��AsgcA$�[�gҝAY�S&���D��=-���;wP[7�,i/�N�OS0I ��$�Iv���b���w��=��e\͟ԙ�3�����+���ơ�ȆD�=kӾ�a^;Q������-t]B��$Jk��Yt]K$�����Ly;C�|��}���<��p���ǅ�$�|�!I),==��B�m%�̴�#��FD��J�OK�8<]䂕���C�Y�u�c�Z�����.�n��Oh�>ԥ��}����8�KHu}�?=�{�$�q�B�^I
[=/>J�*w�p&�k�	�%�]�d	UF/͠�;;�t��iA환K�?���R�-\��)VsA�$M��Y�$V��^BK�;��l�����ǃG��d��bؔ	8���J�D��	$�\@�HZW�}�N�M�%�Y�FD��F�_C�V��N�.?��T�][������(�I(�{��$�X��\�	����QmS��{6�c�ߒ^T��){�EwLP,����R�U30�	o;}+)�u����fo�'`��$�fwa�$I;}�"Sx�{wNέ'W;V�2����$�K�*��c����;����< �2{�9�a�<�>�w�/w#�=;��]���cFo��MCŌ���j�m�͔� 3�$3�����U����7e�X!��V�ly�Ț ��������0ۀn#���7g`��IIR�Ij�1�XK�����QA�N����l�\�w^��]�{5l�F��6�w&�ȇ[�O4t緫�0Z:�:��lN�Mj�A�b{O]���V�2���+ڃn""秶����|룣����j#�g&�T1e�4Gh:���cl�9;j�3ʩ��J�鈇���%�3�c���3��#Ԏ̵t�߽�y�*\������ǹR�H%f�a̤��]}�2<�l�e����u�Zh~��	/j��rd���!�	���)6v��IL*�;�E�9̾h�iI$��W��I%���=(��;(;�gE���ynx[*.;̀��;�t��h(9�.e$���x2@$�{=�;;>31�uD�����I�Z�А�tB�]؇t�&R;�v�A�>�wT�$N����$�6�4�K�$�z݄6k��=�������^@I�0�\2'�yvZiX��H$oz�D��#��&�f0I
O}/)�Yϸ�J($��o[̭r����w�HG�g��g���)ƞ��5���F�&��٪���Z4���Y��K9���e�c���D�7b�J1��<�˟��S��L;�JS�3-�Od����� ��H��=w��5���Ȼ3�����}�D���Ou���h���Ǩ2+��b�Z��Dm�6s�S5�7F1�n?D\������u�����cs�7��~8p[^8�۽���LP���m������ Y�fRI����($�y�vM���12�^�ɠ��r�p��()3�ݱ�	2W�ٹB)$�I��ؗ�����IU�a�tŒA.޷�)M��7���������̐���t�O8�QzItc�a
RI%}��!$B��K���kT��m��Iyt�a�#��-Ļ�.�Ӥ^L�v#'�%����o�a'j=�˶I#0�w`D���H%W��(�M[� ��Gg>�v�$���~���Եخg�>Ŗ�׷-�n�@Fx�5و�, ��������'|�ş�܂�8���I� �͘I&���dzn��P/� ���x%�J�.�,�2b�#^'�@"4j�{a:��$E_K��w�ϓ�_;6r�b�w�Jj�E�vwg� �m��I�������P��C�&:9��"��/$���TI���dA�,CW٫��S�Ӽ��R�%��J��,�o#�Ow�<�b�a���RDK� �2�,|��+�ě�>Jڻ�MLu,r�p�䄌
�[:&�&Q%��>~��U�2I'j�;qyi��/�#�g2��󰐷ݝ��&-��	 ��y���wm�z�lK��D�ߕorfg�<�Q䶯�D�榌}�<�˧%�L3+a,H�.�-Θ�48�q�&�����)L߾|=��c�d]'�!�9�Ĝ��� �6��d�4k梈��P�h{ �gsfMyy����;rϺ&r,�u�{�=���zjr�gē�m��A�8�E��l�Y��Ϟ$4�Wn���C&/2:"vD����I$����"s����3}� �j��H��)���&E;�y�F�M����Xi�w�$����}{s�9�o>>+�q����B���'W/A�_.����μ���;^�1�P�퇕e{=�\o�kys|�*7��fl�C��v��������um��!��X�;���)��:fH>���uwڱ�z�2�WW�$�s��d	���x�a��=��.�����3�B���V���D�42[��1�u�"�lk����Xz�K�r��|��<���}�M��f|A�ۼ�@>��x��i�ח���1�2����7&O��Yn,��:L���>!�6j�20]��A%�y3> �޷�Ij������RnwL1�6�U�����O�g@�	j�$	$�/!�]1�~�n�f̗�y���]}�$3��<T�YΙ�N�&/�x��̡5��D��䁊����H$�O<��t��y�'u�[�+�7d��W�Nal�)�N]4�Tv�'ƺ�bL��cwe/�X�n�E^�L�	 �f<U[� Ǐ�i9��h'ȨEOr�1�L��СW0�ʌW�35\rP��O��K����7���ǔ�nn�7Ak3��E^5����H�&�HE2��%"������^��lr�6F,�,f)��AӞv��K��˶�[6Q�: �h�*W@�պ�G�>2Ÿ�g49n{��2it����J�	Z�$Rb����2�<'n3��g��7�(��av͜�u����݈���X҆!imY��`�65���\p�Z�ܵ6ڍ�����&Vn֦ܪ�Ì��"8z�}n���u��|�w[�6G�i׮2ӷX��'��I�*�S%��G;���vbS��̚�s�C�w$$w�zfI>"�� �I"���M����ȁ�0+#r�r/�	j�Hk�������:dIkݏ7>�0���/v �H$�f<IU�2H7�5�%flF��]x7�>ƫ-ɘ��H�t�P"/j 5W�'���N��A��}Is�?���3��Ć��t3�)���'�^5Z��Ή��r��^OG��H������k#Q���,�g^�	[%]�LC3�Y��������7�(oD�V��mc/�(��U�"I;��2_3o��!�Ajt�N���7���c�-FH�[9hJ�X`^��i��ܲ&����`郳w6_�A�&��bA �Ou�L���\V����x$��Ι�3鎥n�9ܐ��+��$�tef;ia�j7b�����Ѐ�a���Z3}�K��o��'S5^���շ;ǡ�0ͅtS�vT{uw����Y�r�R�]݆��r�赏���*�� �D{�_t�$�~��&W� ��i��*�n�F8��rS+Eݓ���)���3$�H=��2I �d�sn�5s�W�gm�=]�$�}�&��+Y9f(�t�z$���	c�ٌѴ�i�Ȗw����$�I׾{�j�:cf��Mt�[�N9vA���y��[;"�!�XW<u�1H$�]�H$cw<�*n��=mC�o�q�dH	���v���K��z�C�%v�p7F����J��*��~w��}�X���o\Ml������`O�8��~��L�N���6kF�Gx��w�$ϫ��W�`���˳U���f�R��z^�b�$�����$�n�D��<w�#L����7��+�r38!#2Wdt�I�7l>$��:y}t��������Ƿ��On�宁b�]�/'�ߌ��e�R�X՞<�e�v�'v5
��7�w�Wy���9��To�l�#�����=`+�܏7�?|M���]�qw���/׷���շ������>�?�� 7��G5�y o��(�&�A��J�W.Y�e�ʵu�~�=y�} C�^����#�^Ob�c����=��R����e^������S���b�n�2i,���p\#sTg]��G�ٴ���=�P��%�I��
�:��\ǚ}}B��Ȭ��8ɬ�[3<�I�Hf:K)���~�y0NI��e����{9vd�Tbz�|�d�@��a��
���A/z� �-��������Q���;��8��/�{V�vl�����Nt�1��
��=�-�������Q֘�x��9zE�n/x�^c�+{��<��|�<���=�缴��x�|Ʉ'�{��cK�v����Q�<r�>��<��yg����=�F������,EK܇(&Vp�Ȳ��Up*�z#���fx�392'6��(���7����
��<8}��#��r!�F�v���y�Y�(�Q;Ĵ5���>�=�-�ǬR$}R�B��K�`�LiBq	ݚS��X�a}z�9�_۱m������u�׬)o�\��7[�x���zx^�n������ڧ`@���rs�}��{�{���E���'{�3��Ƹ�P��G��L�.o��I�=^�$����Y|p��3�NzGB2rh��Qs���H�����w�X@�`| ����A���NHt�9I�s�t�t!��#���k��I���V\��I�l1�dhh8�J��:#�I�
J�S��.�"JR�)��r�7BS��r��}���8��%3B9Ћ7'E�Ii6�N���I�G�s� q�'AY�gZ�*�Vֈ��աGe��]�u�g�ʒD�:�.,�lm�ٵ��'whR�:M���Ί����I��u��8��K��VM��8���t
�(�()�0��Ivx~�ޑ����̷��n������&�Yݓ;��T�{Ι�|Y|�pH/{s2|I"��4I5�1�vp�^1�8�'�':��}lr�e�L�t�Cذ䌚����i��{�.5��Ȼ�P'��h� ��:�s��2:=I"3
p�8����v�7��r�dj!)�m�ז���w���b×v	���5ޒ	8c:EMwL��b�3d�˜Ϸ�4��|�Hf��AN�$�31y��� �r���3�	��)�h���
j�^:��n��ٍu�6$��T�9`�ŝӳL�2��9�|CU��3��F���$���4x�S[�%�ۺc�	� �� �헶x�5v�ф���!�$}sY�$�|w{,������������6n�Y�尬w�w�ʶ�����^/G�R�7�Kg������*z��V���~��l���X%�Q�ɵ�[��q#�� 櫔��Yݓ;��T���	� ���3��H�-�no�g��R<ݗ
.�Z~�{��}��{��1JM��mh*J%hj�mLS%ōvlĲ�ƺ	1�M�~y~#�Y�X:O���prH;5{A$o_\�0�6i$�(y̺Y��	'�5� ��6���p�݂x�<M섳����A�qh�r	�#&�|O��޾���Bm�����`(����<��N̂	����I��E��0+mv6��F��fI#z��*��.B�Y˻)a�:��\�Cx�[v�$�B�m���D�n�O׊�Zp`�}�����wLC���)���2I�F;gΟFy�	�N_�s�}[��7��3�/���>>gd-���!>�>��B���+2OwMt���\x��ͽ�b��#v�\>�cҧ�#&c-S�4��ɩ\�{��@���Xj�?q��6r�2�5Q
H� Y��h��r�A�n1l�k�Q�Ѻ�; 9�h�'Y9�.�Nϳ�A���4FS :VH)��G�vtVܗ�NW�g0�����a�.��:��0�\q��+S��.7V)���8�#+3/3��g��,a`��K&ٍb��pT^M�b;G7�jF���n]��@Zj��ƻv�t�VN��2�_��(�Ny9va���
�\c�]q/=$V.��.\׮}�x/�vGaP���yν:���I �f\� �O�GsAR�. J�u����k{.f���Ȃ��A�x���93��^���Z��/�1���֛���4 H���{��lC��Vi G��	�vo38r��P�.�ܡ$��=|H2�e� �8�ݓ�	��ɐA9�<�=�J)�NRd�/":�z"޻�v�y c��}� �O�a��$�3]Ңi��'|�t��H�Йrvb�]�L��h�A�/+��� к��ˊ�����g5ǹO���`��ށ9�\��Ծ��n����9�{���V �S,�B�B])c/4Jd����Rb�y���/5��B��+�@�	�x$fo�d3�w�¶7A����Nut9�|��hL�ɝ�3%T��L�AL�E��fr�\9�o�ް=Fo~'�����s��z�=���a�M���=�g<���v���#v��N2]YZ��8��rL�8u��Ct��ۯ.� �=^p��;+�O�kzd�m�Цn7lb���,	#=p{mdANY"�=P.�� �	;5��I �f�c&�l}S���O�j�B	5�3�|ۘKc���d�D�z'-�av�Z��SE඀��&<C#^D
m��H;�Y<,�m�������h ���f�tK'��LmL�����ztC��j��M1�1��kԽ���5`�ݕ��Z��v;��)����v�퍶��:b�%l;m�����ߔN��M�jmW>{o��u��]vN���T@rI59�3�A$����vJ��,�K�h����	�����uݛ�Jg@�fA]�2$��^��&��^��o$D��L�Iz��H ��5�gV�2��|@\��X�w,���̢^�6g����yq^!x��fe���"&hP���"�I=���/O"�K̗O-���if��:���_k([�~$[|�'2x/L�k��-�6��ˇ�zy��q��~x����$�~���M1�A��'D�I�@.^�nIn	�,n�$����9�]3��R�ͭM2Gv7�w����8�'�Swp*�gљ���@��p�}�=Y'Ĝ:��K�l7[�R�Y`��ɐI �Od�>'G4MX"U��:ML�B|��.P	Et;Lv��V��;8��e6+1=�^�m1a�aoREˠK'�َ�����I����9�mi���"A�gVD�zM
�!9f)˻)�=P�z�=8�S$�Ȝƾ���>$�md	 �]\�H7�}��2��Nh/�'ټ�t�
�}� �h�ty�|��DM��3�״ �ά��	ŷ��{f�,���ٙ���GN]�5�ef��
�����=���+�Q�<�z����f-0�+.}2MI�w���EܳV�٫i��I�(��X�M�{��^��0^��%=ƈ����S�#�6q\����%��'��"�H�<B����]'��FÒAɮȟ�(9�1�B=�s>'ā�o� $����&�k����b��̉M��ݥp��v&��F���v�k�WM�=�]�	S�����d��$'O��{�UnP��|vWt7����}��0�e�T)�8==�"A���Q�@<P[�����꽓S$�>҅ݑ[���A�2��zB>��I<t+����B��m/Dȩt��d�;��ЛU��S�� �J�#���bH�@$��t	���]�rɝ�A@��n�"{������A���@��ɓ��[]��ũv��{z�[#�^�֎�]�N߾�:����^l��ƕʵ��6�$��Ι���TB����a�\�����uS֢��Bޗ]�ꬣmlb=J�i���n�Cq�n9�!�)���׆{7K��{}�V����wR�҈QFC^9���ޡϲ�ѡ��G�6��6��1˴iXb3k��b�cM2T4.��b�v4t��*hi�@�ܦ�>��ݽ�!�#�..�d��Ǎ4�Ί����;i4�a�q�f�L'=wR�Y�3u�㮸9��J<�&�b�zgf�\z��(�`� m��n!�:�I��l`(��5h���+�nݴ���^�nk�8jugE�Y�<�3�\Hi����f���6�p�svĻ�!v���[����]���n��3)R�3|�����Rin�����B�d�d	'��{� }���a:x���O�>��ɒSnk`萝?�=D�@�V@�vuUN�X���s� ��ھ�Hy*ި	������гfy�X$(��q)/8rK'�ٍ��A>7�Q��g=<t?pi�1��O�N�Cz@@���@�(p�:�L��]�L��<�N��z����'��$�Ǎ��	 �ͨ�A�P#��nԶ�?�72�����wfY2tQ>+v $�7��zj��ۚV�VQ#/#&|}׵�I���kWC�}�7�ν�X54-��X(i���ڼB\��mT��3 ��ic��j2�����Gj.ȧ���p���T⯺ A�6��6i�3������ɒ@'�:r �~TCcAA�.�L���<x�'��V���b�iq4*���o�H�CM�B��2ne.���Xf@PKA�7���
f�%D�dɫk��Qt���)�_<
�:�]��O�\�� �ި	7tei�7�����^�&�����"�vr�$��<���̩ײf�+xI۝�$�}{�U`�J^p��O��WWx��Hk~��e��w�zs�ruᲝ�Q�]��]�#(��n�:gvb��d�u8�O����@�C(��l
LE[����S�	7��%����߿G��vX)�����n�k�9�x��5��������ݶTz�����f��䅽�������8�H��-d����4��=�':�A/.����3:tYL����%�]�9��mw[Ȃ+�@�z� �|O�o�d�j^e��U�WD�J�l`�NI.�!����OMvD�I��Q���zB��`k�$JS�&&4�w��8�r1��:�N����Ԏ��u������O�]��V���]���t�"~�l��H�ߪ�}Kcqc1NN�D��i����� ۊ��͸@$T�tω ���G]�3���4Ux�>�2�i%/3�C��鍩���]�tF�\�xHg������ �I۞�Ax�IԊ%���a3�	�'a�ڒ�3�/���B���Qu��UY�o\i����d��N��3�1vu����|js:'��	랈 ����ʽ��� ON�̗��ݛ���rC@8�pDy0ˠ�}|q)S^�؇>7�|O�r�gĒu�H�K��0�(�)�:�{�͈�w)��p�+9�0�yr�x�ܪ�qp�Y��N�I��ٟA랈>����x����2>?c��RY��͝�$�|og�<H�{���5ц.V����Z���k/�/`��g��'��{�Ǌ�a$�;�\L��s�:�Kۻ��+B�jdӾ]�:��ӒY�$�-�^�f0���z��H�\n�f)�	��^=;Q�۔�Mo*8�̄��&�gdO��휏@ �}�Z��&��E�]p��;�̝��e�ٶ�"kK5��$u��֣g#ڭ������Jd?pm��2	����A;�P �ص����wOC�!q�z�	$�n<
�^5'g.��gS'�����ge�+�h�m{�w@�H'c:=s�= �Zp��w�8s�����rX8%�AM�I7]/ I���Ǜ �U�ϔ	$�gG�7:`@�vu���.3��Uc�dHCJe�$��@��؈!���꺁 �EoI��[�M(��艊���x���4H���:+�$x�ⶬ�=8�q��1 �[s	�Ƚ�o��8�������g����Ƿ���G	�Y��߼�aP?c��r��痑���$�mi�}���}C���.�yo{=�/��j΁{g��m5q��gb��|�k���YS;�^m�9f�&��|/w�{�3Wb�1�q������wy�m+�׺*��HkaW��aN��N�e�]��i�fc�w`=�x�m&-���ﴸ����o�r\P9,�=�9염��#��O-z��Mn��r��� ���=�����C�`���'$ќ}�]��d������x".yq�,�,��9�|/�Y��7�<��u@/7��<-��P�G>^tǖ�89g9�Nhҽ��Gx���<��AY{�Oc��dm�}qv�����*L.7���1����7�Jz��]y?*��p�S�{�'������B��2m�3}��g��Oc]���z ��pOQ�C��
�c}���[WV6�ܥ�bDOs��}J�����:v��GNl�8~��s��3��I�
��|�o���G}�g���O�=�x�[7��=|Ƹac�9���yL7eB�&^�m��(�޾�X������5���t���<�j��' �[��<g�x���sü�k'���#�<7����^��&�:���ϜDl�θY���Ɗ�);/�|=�R��n�c���wE�}�׆;�yg��/o�;|�y{���vt{jG�d�=�����⇬���Ǡ�q���Խ��+��N@ՏuG�N����mgl�b�o�`�7�
'�e�Zثyb���}�5t��}}q�&{NR���b��~�2�ŕw O���\17�
���b�L��7 8wեc�L���w/`���Vd�'8�'	�Pddvg-��R	�H�#���:�kG���$Q yf��8�kG[Yʋ��O2ëM��Q�۝��9Fd���ⶱ��Ӭ�Y�v�6բD���q�㸎;mY7)����e��ߊ��!��;9�m��Zq?�|�;�6�ʲͷr�w�Kc",k']����촢*͵�e��flƖQ�{n�:���ozK���c�î,�������u�4��לVVq�\tڲ�fD]f]�����ò-m�Y�\ڐ�ku�Q�]�y��vi�nYݶ̋,�����@�:U�q�qf�v}�ze��sh������vs���mm����rsn�8��0!yo9Ai�^H�Y}������k֋�/\ٞ�׬Iw�7�ְ[D��3.����u`���T�Ƃ��Q6��,�^�Z�4���\�Vⶴk��x7U��
��@|m%r������>o��� �l�,��dԂ3bWL�V�e�k4�1�^��qM����C����kz�s&��F�����6�,�A�(����'O���G`Wc��'4=��ɐ�[�������.+��@�%м��4`(��5�[�q�RsVmq�]��P���5C�*�Ca+s]��N-��n��щ�m������D�ѦǦ�:�T�����籇F��u7���qVɸR�i�r/\<\�,����C���\08�m�n�k@�m�s/�s�(v,K���6��1��͡a���歶���۪)x��ŶNl�e6���;nI�=�Sn2��-��bU���:������cn�l7ln��d������j+�;m&��q����!9�9���؝�v�콲&��'����9]��hx��Wme���W7[�M��ފ�����!!���L����JYMq��ۋ�Mi����Z;�8�8H��;vguGQ�Ύ ො5���ڨ�Z��l�v����uh�v�:���[n�m���톽������lһ��\�^t�nn;7d˔�k�K�K�v��p�r���9�m� ̖sft�-����%��퓴��]��Ƴ,���OW���8�-�pm�[�ۖ�8���-�F���;:��i[rW^k�F=cۮ���犱OV]���)�#)ֲ��)�n�i�������f��'�\t���Wiu]/4e�
�iFi��� &7.��<A�6kL%�;u����nޘ^�b������NQ{�!!�:�%�6ӽr#o��r\��k�G��6����W��ur��3�F�n܌����ZՍ��"�bL؉1��k\p=fahC]r���mV�Z%���a̦��l,%��]8��a9��ݫ�oK��]�d���&����;\k�
7,v˳S�� �{j֛5��`�n���N޼��ǚ]ִ�/F90�9:��#a�7<�Gb갞�]o��kԬ�:B������[�yS�N|��A�#狶pF�:A��� ��t[jFݙpÎ���$B���E�b�6#�ln̗ڽH�2�Yg��4i�v�t65�@otvw='K���V�ڔ55�ז��������6�3���k���z�����d��Aٽ���HV��E?Dzo%�B$��IL��C���LuH��'�	d����'+f�|:o�D�^W��9�����A��bu;3�gEgU@�8�S��$��G����R^2�$j�\@'����ωϦ�;7��"���)��;Z0�V�$����^A��4��I>'Ǣ�l����t���l�8L��h�ױ�$�:/"2�m԰���.��zAٻȒ|O���C���?�ߓ������_˥�k�����)6��,s	���M��T�J�-�1��^Rm2O�}���f�雸��� �rkr$_�k_@5+��s��U�m����fL�����g�E��;&lG����&��ء�j6��\�g/�iC}og�?soƭ7�]���Q���{r�'����r�-��N�}r�/YB����F���D5| �l��L�O��G���X�=V�#c}N��I�I�Ē̃�!����T� ������
Xz���GNvL�I=�D�^5;3���������B'qkl�q�n���x��\I MGtA>��5�:�ER�9�vd:&vo3�	�-2Sn��+�U�L���ڜ�bz:�d�㱙�_sA���+�\���I����?1��&0g;����mc����3��t�X��åƎuڭ����|h�2�h����tψ'c1���Ξ���y��}�I��ވ3M�vY� �2��v�� �w��rSw^�n7MFH$d^�o��s��If��{��}}� ��dwjd���x��ü���W=ݭ��>깒���zؚ2t;5��g2(*�$S���x��u��s�T��x1�^�^F�Qq>�&����"x���[�N�w���v)�xS��^���$O���z<E��& $Ă�%`�b�ؐ���LuMq#q=1>*7�A �O�-��$���m5��
�c�Ei18�����NY<O��5@D��NgEQ�ݨ���i���J���I#s^�O��$�lx��݄��ּs��Mϋ�֤�>�cR�F�*[Cq,9U�0�J�iIv���~��<�a�Яr�������Q�O�;5�2Uq�O�����ȝFwyP��2�=��ҀD�Մɇ���L��g�{�Q5�O3�=U G����ߗU�EL���0�U=ez
�W����)���l�$��d	�$E?�XZ�e��A3|�cď�މ_p��KÇ.�tFk�n�6���L�`H��ْ	��8���ۆ��j�#dc�M<44�X�)^�U�PǇ�B=�m��j|-�E
�{(L���L�6���K-�Q-�s��ꣳ�k./� {%��%�J�>!��O3�S �s:���^G@��y����F|�VETe�a$�ި�Zط\�'@�АJ	�"�����At@�tۤ�ۗ�r�I5g��S�5Վp����}1�wb��O��_ajs6$�I"�� �V�f��F�l<���od�m��ټȗi�n�L�Tw)����D�1Y�$�ޘ���}V\�A��+��=�c�!ǉ% �Y�	p���L_�F�����(��̎��g��$&+:gĂ+�`A�5N�k���.S���'V���QΖJ׋� �r�b	�$;y�����`|[ɻ�N�uL�:3	vw�]�9p�nS����)����M����6�I �Ƹ�w9�� P�󶣔�?#���P�Cާ�kk����x�������E4���*���}�o�Z�#��ΎA��b^}���͟�����U�:�\���%sh�o%�y���k�Ä�W��tsű@���{����x�F�1��r5��Zi���ehX�"S�����g�F�mlv�l�˭8"�v:�x���R��=��w��v�"���S�u1�-JK��Ymrv,�Kn��[A���`zɓ��:C,'h�s�a=6u�D�J-L���,���l�F����w/1����,vP�s���X�'h,��B� ��p\����c��C1�H$vs�yI3��*nAo;2�g*��I�&�z!yV�թӳ����O2[y�<��SCC��O�I6z#���u� ����D2��/������8p�@�m�$��V=��:��3t��ǝ�	@$��{0e�ks3;����h�5�t�S�iDXxQz~̀ �@+/^̀O�E�GFa��[���|�@��G���l��ı� d3e�H;�tL�sA��z� ��ȏO���ǈ=�2V:s`�͓4� C[���38.ܗ=i��͹�	�:�m���D��6���q~.�9��<'v:��ܨ��k�� �6/zE��e�/m�up�;�ݏ�!y���!ד&p�'��2H��b��ID�z���j�f�IKX)ȡ/'���G[�O���c���,ڊ���s�O[�����&ok��6�2L*������_9�����`�N����"��@%�Tw=��H��K֧I����yy��"�3�I =�-B�ΦМ��@ �7of	$t^�ω}���,Rw%�L�w��Sya��00I�ֈ�@��C�7jI$��+-���<�Bk4q݆� ��<�mfgp]��p�TՑ�$�t�z7�"V�5̖����oF	�#"��G��[\�N��M�'`��1�E���΋\�-�4�`A	p-��W(�rkLÁ�*C[ �o_lY���K��{�eۡ_+�$�z#�o��6��(�{1�I��wL�u�1�SҒ�
s��l��.y#��ܙ'���O@�@7W�=���SU��1�C?#�C�'L��O2�S$�Fd�@ ��&f���r��^&o����?	��U�x?,�8╺��%ɔn��e�=�0�X��}���NcRuuR+�5}�@%��6d	5��zq/X��wdRfI�Am曘��˥}��7�z$O��\�A$��{9u{��YLa�-����ː��v�;��N;��c\*W$�E����I�z=#���x��z���/
������`����EMRks.�����f���r���q�ύ3���Y��t�8f�Ml�z$���f��AS[�Ձ7�>$�r��	w��-g�!˳	�z]��06E���#��eŽE�۞d��� ؎'#�k.�>
�F�h$lfd�`����A��x�"���zB��j�v�&�u� ^�c؉&��= �:���;d�\����xB:b��UQ�i��P;����Ē���$�{�z�8��Wz�BU �7S���-��:��!a�|��H��O�^������ˍ-0�/��ڙb�.���F��}YOc!$���Q����h0���>��#M<{0������)1d��}���_F�mdab��S	�E\����֣d�O�/zd��>��~����X���'����6�ss�4a�;	֚7k���λ���-9M}X1�1L�-�o�$�k�"	 ���5�w���#h��v�c��>of�Y�HU ��d�ӗ	�4�^GL�e�h�D��Vz$��{0=�"L�,kp�勂nWgT&6O���ć)�0���,"	��ȟ�(��9���L��mɜ��v[��5�FF���N�҆t���_W'�.Ll+�vy�<#̼H&�{dO�&�7��ۙe޸�v�P�����R~O�� y��#n�2���_$��I�?^@�*;���s��Z,�'	㮼�c]��&��f��{"�x���X�ˏ_���a�\�t��̎'��3v�#8�ǻҀ�03�kq�:��[�<$1��/����K��͍�#�bX�Fxئ۶��ڳf�Ak1�t�ŭ£��m
�ls��	�϶lݎa<6E]0LA�-,�`Ė�q��Q̶hM�r\�h��O.�xIx2�ݳ�����t����7���FzC�Ƿ/�%x�h�͵��uN[��$V��Vn3��v9��E#��p5�x+K،۴婖��]����f����&��㝺��#��^y7��FmF\g���}�|�����{��޳�|I���H$TwF��Q�ژ'�hsK��|i�'ć΀���ɐg�N3�Az-駱�%,���m�5b$}ޙ �|j7�z�NO�]�d��Ok;2t�p��vd�	4���$����^9NloW�$�O����X��ė)�L�M���{��E�x��ӱ>$E���"w�0�L��S��H輙��Ì��������_TA���k���S��f��7R{��ȏwkY�����������3����bR�,�-��H���E2�lnֳF�]Q��s�(ݍ�Ϟ_O�.Qvv.Ⱦ��52O��Έ>$��f�4G�x���e�L��ѻ|%��	��;&	b�f�����}u��v��go�_��:L��(�;t�����<�/nH߰nE��q�j�# ��=A����77tv��}�uy�"�@���^�����tW�w�$�'��=�����ս=�?t��h�;}`�ݐ3��1�]�d��|H7��DWg�k�q����>H>̎�w��<�ĵO��t����e��$��[�(5rO�>�z	$��{0H$k�t��)���p	=1�1���dK��$��`��ّ �6�{QN��Am�x"�ZȂG?gL���܆��/��I��3	b��gL_�=V�N�]��G9Q��f�[q5��ؒ������+��P�����@>�	=z��I�����-��p#	��{�켈� �]%�t���ܗ��53�AV6%��Q[W� ����f	�<��2	�Ms�6Y��N�U���$�̜}j��[��rԘ>�;;>�����}t���������wy7x�2T�7�u��������[���-���ӫ�W��n��o]�e���geY���~	_�e��^��l���{y���m�y�@4�I�V�0���Y��v�W�^�������q���'�jg���`���y�~���3�*����S���C�̬� ���{.�F�
�V}��szn\�_��d�o���[�&��5��;���K����h�(���������ݐ�yx�YHy���������w�p�fy�@z�nB�%�ׯܧaZ�yv����tg�3��}�����1n�qyF�*�f�b�g��!����/#�Y�{�
xfv��y�F������﹠�cw�m��
��l�D;�]��S�5i�a��rw�;�"��'v;��F�:{¬Ou	g���>�Al�S��^����|R���c�׸}�|���jۻW=�a2��3潜���{-�w�;��l�&y#�4vk[���|��绰��\jV1�FM᯽���H'��@�ͷ���x�.wvu]����ݏ�_�ǊL@�TJ\�m5��g/n�6��zR��b-:m�W�N���9�\��>�>1gbʅ�e�w{�qe�g�7�����u�����i���h��wb����tp�O2߲����V6r����{}��vL��&���mRk�p{Ԃ���� ���3���Fr'��\�+�O}�1�xG�m�B����G�1��BÅ�`�q��0-�\ `��B�w$�{a�l���d���ε�d���]N�Av�]�[�Yٕ�V���'iV�|ʼ���+l_0��h�6�ٴ�.�4�۳��Vgdsh��"����"�,�BB� S,���!�e��{6���YQ[k����nm�Q�m�,��gw��+;�on��2vwi�Y�w������m�;4����mgqw��k�;mGv��ѕ��Tqf۳,��F�Vgy��ݗy��l���s������(������Qsۊ��hv���x�Ͳi��:�:�6�
{xw��ｫ��d3WȬ���춷F۶�m����/:��,��"6%��e�֤9��y^��(�������Q���[n�)�qGm���*�qE�����Ee׳�}v^YKn�-�%�'�e�q��+<�έA![@�<;9�kZ�;�~�ב��2s�L�$�C;�f��ݸk���a�U� <��`�K]fL�	5����7j�޹d@�����I�S�-�3;;��2����H>�2`�8c ��|"<H��2	�>5�όcy���:�Guz���5�ͤ[R���*�:�*�W�ci�Kd�fd��e�w��,͉n�g����������&�M���t�����7u��|�W�g�Gg#�H�F`�E1��0!�$���MF��
Y̓:w�'ȐEGoL��B򭎘�`U�i�;h�/Is&gfwE�y�jdH2: �	�p��ׇ	����I ���V����$�̞�ǰD��zL�n���f�	�>'v:}�d
�6�?C�*q8����&��q��f���S�s/��Cq�Ogno��|�fJ8�����&؇i���4���wZu��Q����9�^
��剺��s.�d�Ր1t�Yܻ4�f�A>3|�e��TQ�{�{g6d��tP��� �f
3VW7�����M㡐�[�&���1W����Ӫ�=���4ll�f%�ߟl��ȹqM�_w�2O�5ѐ ��o���7sLǱ�=D�te�@^cp��A`\�a2a���+��odT������I���	��=� ���Y�h��ь�0��0!�'�7* ���p� ��̶����#x���� �79���V%�It���ˇ��驅Z���l��XK_T� �@$v��	�73�[S3乮�!���b��ĝ�;�1y�wa�<� �^tO��b�Ux��e����Ι 7��ӑ��n��2�4��Yc��+�J��dgl��{V���"�����fp�ÏU��~���,<_۸�Ǭ�_�/�Ǳ����(�nl:�,+p"[��t���b�0���]u�L8���kb!�	��+�G4�\��[�Y�̓�nx�v.�K���]B鈤]4v�s-ή���	5ۉ�|��9����i2������$��֪���7mt�8���x:��ݳ�0]\�Dծ��;�UV�\݁������t�,F��d�����\L�5����vU�.���Z��O5�j��/@4���ָ�-��$���?{��pg�>�n�� D�6;:d���1�)�o��|�F_�f	�3�'��3;3��2��k|�dLlDUet��y�QQ^G��k�|O�7:g�]��j{vֱ����#
�j9&~>y�:;2$M�W�醭�5y�I9X�`ZGgw�OFhX�0���y�$��s�����t�O_�|v�<$���� �[��Jg���h�qmf<��V�铳9p�8�52H$�GD[��\�`�_�>�w� �M�[a$zߢ;T���K��,�[�u��t��gDDمA�4=vt����e@ ���te�\�˾Oߧ��3��E��2ݧ�A ��lI$u�<�1[���oK�.�������#|��e�����5P-�o༚��,�z1DJZhE<��;ܳ���{��h���J�[$Vx����ˋ0�a��!�1�T(�
�o��Fܹ%�
2�qI�Q�cWr��ۺ�ș�Dm>�'�nz#��_X�|�u�{��?�f�E��b�2�U�ǎ�$\��'��P{�^�ٯ �e�I��O�s���,��&J�l�3�,���/5�����NY �W\HV�$��@�H��ղdp���i���y��$P��G
f���`�h�UT�FzP#�Z�-�i�5c�?�5�ޠ�$[N@�I�g=)p옿\���D�F���;�����p[���V�z�t���m��#.����jߟ>���l�ˇ�w{bb�|I&�y� N�=�׎�&�lU��}"A �OD~�<)�'gv`R,��i�M>��]m�j&(�	˜�����j��4��3d��E��v)�]7z�&�	���{�u��֕�e��PUF�t�<B���k�U�K"ղ�b�}�R���m��y��tFs��d��o{L��1���A����PL���fw��I̞q ��|�DyG�OD��b�YJ�~���f�ǦhE��� �=@�	�5X�D�ޗy�g�v�{�@4�0 �^Q+���	�Ndd3e�I �_dI�õ@��,)��|3���"��A��3=�����w=\Wb�:�n��e<���7��E��i��맇fd�wf,���#/և�ǧj=ku�� ��ޑ���݅�
�^�zd�	�7=��2�ćL��ˇ�g�$��Ez�5�`��z����c�����ܡQv��P�O�����c��)�ݘ���Z�FgD��L�
��m�Z�=SI�E3�I�ף ��ޙ�=��3���t�L��~̈́#�4�3���v3:$@-����0�j{��J����}/�U�M<�#���!�n���5ʻ=l������/^�%�=a�VY{��ˊ9W�;*�t��hb��9����ľ��/��N��Iw��1�l{��|z� B~%��ps��^�j�$��ޑ ����GL�;��!��2�3[�a%���Kl��MCnk��y	�h��H��S��Vx ��,������>��^#Z9��d���yC��E�nH���F&^/-�"A�ʁ�L�b�����i���|I9�2	�[�Oa���Ǌ�gi�ƅD�ئn�y�'fr��H�52O�>9�� �������Jz�T�AW����"��]T9R�wgN��<ϋjꨙC6�����Đ_{�$�O������R�ذ����� �ݱE��AؗN�4��~����R�"�5d㲪�O7uL�|H=��#�ۜ�|+��!=���CW�|��-������!v���&DF�SC��m�3-�N��3vL�h�(]JD��|�״�|O����w�Y;+n����#�߼�)�wuj�"�Q��̘^��ͽ;a�@��ʱ�Z�n֘�%�O�cv�L�rv-�g[��	����uɅ��v���C�#���7�j\Ag��7���x�;E'&�^H�X�w�ʛ�e�Y6ԥ���4U�Wѵպx�F\DhP��#�!I��]il�Tk�[�Ƚ���`�r	�1U��: nm)16��t�*+O�SD�3)����һ���q����%�w�1D�ݫ�v� u����[j����p�\3����>ձ� N����	�tZf�D<t\� ���x��Y����NJu2y�� �=�+)B��D\I tc�'��k�R�9�-&'�Q��������DO�nS�$�k�I&�{�Pʗ����q� ){�^� O��sm�Cy�'fb����ak���v��> ��z0H$s�t�lksE�դ���49J�wb���L��o���Ή��Z�ގ�o=�q�S�G���� �{c:d�t���_������P:���!�Y��h�����뛮�7Bjְ]u �٬�4T������͸t黁�|�>"���	�3�MF�8-��tTo	�ǳ��\�pC�v.��f��B>oW_,9��^EP�ɏ����&C&yn�n�7��R�-���Գ]��t�γϯa�i��j��e���9N�j���H'�v�`�|7c:D��ޗΊ�¶��O���;`�.`����m�A':3"|A/6�9�K��Of=�'63�A"6�����Ç�t�gV��j�p����o����#/���A��W����1o�t�рLdSk��t�٘��犋$�Η��8�yZ8h�qo&<H'ٱ�2O���ToZ n��ȐGu����EjX�>' Ÿ�[�Q[g��4b�h^]�f�`�}�3�v2~�y��$�n�:d�H��#��
=��-�����"{� �>{�H�BbX�S&_b F��s:�Z��|����&|H$��	k�����v�,�%ܻ�V��`'���O��_V����1l��"����$,���[��B�0C`0�aޫt>Aǚr�Ftۤ�۽�}�'O��3(��E_zG�s�w��b�"ﴎ'��A$���\� �,���L�WKg1��	=��6vTP/�����υ�J�bk	�U��P$7�;y�����ۇ�D��TμA�֨<�uT�ӹ��b�q���f|!��� @$�cрn2��_"p�>�y}�������a+�lrْ�P�R,�3�;���L�Y�Mq4��7&���5��\����;ɩ�G��m�x��z1�x�x�y{���dI&�.CޕM���݃L�׏G6B&��~X��6�auEή�(W� �u�A���fA �m�Գ+�����_L�Ą�Ӕ�� �tD��@D��\5<���=|�7�޼�|H9�o�ݏFv�,9%ܸg�Kc�K)��C���'�9� �Iv�`	]= ?�W���\��-H9�������x�_�=�ˡ�u�y�F�����q<� \�~�ۆ���h�q�k�:k!��`o�y��ln�,d]�,�[#��q�q�`7_36�+�"	$�z0I;�2u�\u��Q��|�D��z%t�t��h�l]��pc�Nɮ�{lۃcD�2���1�x�v\�h~�fz �Oʇ$���L�9�����=3p#��]8����,���:y�~��$۴o�/6Եd���A�A��x$���� c���-�w�؟>�V��3�`�'� ���>�M��D�I�&��O�v�$�����龙�l���������'���C�E��DF{0�B���@'�{�A�T�[В;:�>MvP���vp���6d	5�/��G�������d<D<A"�s�O�����e��8��������wO��OOO���F5qq}����)B�j���6T��w�u\�{<���M;�p��K��J{���T5/4T��Li�T��� �F�RX��!a�-X�� p��5��
��|Y&���$�_yw��=�g���wʀ�2��:�îx62K���=���rˆ����v%��Sk%=é����Ğ����u��E>`�'���{��7�;� ?B:yvlGh}�s�@M~���v�/Ls�x;�~�����)��3#	���$��ו�Q�y�.�ʙ�B(Ĝ$.�+.���uv(�]y	"v�7�����W��z�/�ޯq��Ƕ0{P��zw�ɨ�&�U�Ǫ͇�����`�0�ܹ"���x�>ŜZC�c�޻W����ދ�R)����sNwwv�5s߻9Zٛ�����ȭ�r����6���26�@����b�y�wNj�qn��޼�V��u���U�v���8���j��:����4�����F��3���K�_�i��_w�*�< ��06��.g�^�jRT3}\3}ɽ=��A'�W�7�����i�Д�#�U�e..ν]��z~������z�^�IW)��t����Rgx<��ϱv-��o-�q�vjZ�V���;P*���l�[W��7��/�|���o�/f�>/����=G�����:o`�=%=��h��L^���J���MLP0M��(O=�����T�V���[���{�{�gC=���,��:��9�7�7��C*ŒaӘF��"<�#Nt qLzV�`��w�g���e��r��&���{tw�Y�ͻ��y��{wYF]�����ˎ�mee�vG3�����{�������gw�۽�w���+;:üf��/�n{dv���9��u�n#��2췷[j޷�7�e�g�|��m��W��7��������w�[6�p�,���䢲˽��Y[h�1�mee��N��lvu�Y�C��,�����8��.N�Yv�vt�i���m�k��n�ݓ6�Q�vgn�N��ΰm_z����/{w��Y���+K�33��q�[:-٫�ΎB��NN��[n�>�禍kc�;3n�]���u���۬+s8���۳��!�ז�k9�:w�=��ۖ�dZ6�9:s�O/mygg���z��۵��#GM��fm[������}��}�=�w�٦$ZW�ݸ�{V�0s���^���l�ɤȠ�>���ͭ��&��6j���מ�λLZϋ'U��l`�y!�Gg�Y�ri8�n�A��]l)��7%n$��H�	��x��L͑�*�^U�J�)/nbeټ�7n ��������A�6�P�:�[�Qř��%�	Z�,c�� �̈.�%�i�2���X�[��ǖ��f���qd_d���6n�5	Y�	h�6�b�*�hS��Yt�q�F�e*���C�m�8�[�0�&��pZ�U���
�;܂��s�Z[]�8�^r��v�㵲C`֙�j���D#�i.I�˃�m�s��΂�n�����Q+qx�� �j��c���>�<� y�s��ݶ����/73y���$�l�jb&���tкH���;�� mM�,��9��Z��qļ�n.��\"d.t-,��rSm�5n��D��������M�ݽ Z��K��W���q�3�3�Ya:�/v �M��iIg٢�J��n�G<8��R�;��ڸ�crqr���<g���IӢ�o]�_ڝ��l�)y�:9�Vq���p>�8�.�=����4�˜f�;-{u�h�v7�z�͵�����[��6z�C�9�!��lā1#c�$��0L�k�OQq����+s�֬v��6�t=���iq�7.h؎��n�5�'M
1�1��*��BZ����C����/W.r8�sν�q��oW<q��[��'=e��k5�4�B��l���3zn0���@�lm�d�m�k��捌G�웋M��`����;�x��k����ں�䊫�L[0��v`��c���8�m�k��ю�v��KJ9ݸ�и]e�4X�T]�pܲ�j3��,�\rt3�B�S�M�<t��n]=1bQ��x��LO %vf�nk���\�|]��b	����,)Q�m�-�����G�k.ݶNsOx��Ct�oW;�q�`\U��Ӯ��5r�t�UZ�Uh���{]t��M/k�o�q��wMFa���h�m����4��u�fۗ=����8��m�Zn+د��jʥ���m��L�j�S1t�\�&�%�,�ҙ-�[,��
�э�3-��(��kh�k!�!ΪK=��v�lv�P�u��&�&XJ˪0!D��h#��5֠'�۳����ۛ:ȶ:�LPWa��ӹ�w;��3/��8qt.3�����m�.�y�pkg���rؔ�2b2u�%�����r�E�N��QY|O���D�I&����ZT�	昙�+f	�5ӽ2	��c�' ��X44���NSq���wm+�詉� �H���x��Ǡ1o��A���]O��kb���v#v��s� VtǠ���י���GR�/�	 ��$�]���mwN�0I�Ă9����,[�e�sͽ���>/�}	 �H�� {����57�s	�93�|��!�1!wA;4�8� E��E���o��Nz;;*�O��= we���7/T��7�l[R��pi'iӸ�R��qh�	v���b�]�ڳ��vE�.�!��ȧp�]�s��L��@5�1�$�{�����N�N���A�/#㭓�#��NbA�Y	;]���zyǧ���N�������&�}��)�ݙr�,/S]A�܍(��ҖILF��h�lS�yp�ڥ̛�Y-)�P��j���לs.��>$����O.�h����ŸE����b��I�.�u,>��Oˇ �]�e��g�]�x�ё ����lgA�]�3��uUN��;S�S�5�	#շ"I>$j�ƂI�t�N�^�Y�� �]y�S�����;��<�Ţ�	7s�	��U�H���qH$Y��I#v3�|nD�v�f����%��3ȹ=�������K� s�����^l,&G^�#�Gߞ��ȆbB�vQ��DO����$��작k�Pҥ��ǌq��Z�!�↡����p�]�n��ٙ�M�p�U���π�	�[m$�ۓ��!\a�׭ƭ�꽃�#� �,����AG� ��ND�H$_��d�:�W��V7�y�*.�n]���U�?��~s�9#Rآ�Y7�*��j��2VR9sח�t�m�����4�׽��{���0���f��.�YbKd�GG,�a�2���1V�ad�:E�B&;j{9ጶL.���/�~=��?����O�l�u����V�18�)���Y�@�f�3�S�9��"�eF��H��m �NgN̂A ��@�L@��lJ\�]���H|���ZU��*j�"�!L+�E�Њ\�X[04o���I��;Gl����S�ݳSJ�L�|p��8 ���I$�]���t��Uߵ
v�B<H�ٟ7�:d0f%��e2qߢ(&��Kf�I�X$������>6������g[銮����σ����Y�&.��5gL��I5ё~�"^�sbc�f߳1@${� V�9�p{���	�Nv��&e9#���꧊ぼ���$�D��ȀI#�����K�;����L�7)�*yd�K*և��@f)��;�KUk������[Vm��ⷘo�Æ,�Ӂ��*��qUsTdW2�[i�JW��ǧ���:�-Ў����ʶ0�k�\3�F?m�H�'1yy0�Q A��q���C��d9.r��{�w���H,�:/kv�-<��u�rRb�p^P�2���.�-��i;�����%�ɮ�=�|�ML�Nds�$��{0f�̃IU�ᣗ�=3$��s#"
���]��'�&y���p!�ĵ��d�D�|I+.:d���f �T5��^�L
3����%�1H�wH�)�w�	��� X�;;�V�6��:�-�[�xDx�{���$SEC��1gp��P*��:ssx���Jm�CE��$*������l���紐�UT#�FQE�Y	;L���{�3"A����Y��#�� H�׳ �����uޙ'xilu�����e0�ݦ�/� ��P��}8��O{�Ogo�?5�����Ѽ�'��y���� �Q削��'�A�}>�������Gh:�G^��2gb٠ݠ��v����!��n^���u��c2'h��걷�k�z뷨����+;�X)�������ͪ6N��ƫ=tu�����p�Y�M[����94M`��I,�'�&ೞ��qc�]7����s��=e�Zf�,��&�%eRTw+XQ(�8f�&��m�c@�Tp�]��m%&����F��N�:-i�^ڪ����c�!�4S�n�T玈�a��Z�m,�(�8��������}�7�1�O�~����>$��Ι5���;��v�@$��� O��ry�:	�����Y<�����`���˃��3�zd?\��Et�c�u쪗�!H�e�����S<N-�k� |o6r$�I��T��+xn��Lմ	��ُOnOL��tI`�PA��,Z&�%�@f�|HL��oM3�G�� �̞�I��V쓼�����{��
Da�Ӈw˅2��D�I����mZ��x��p�^`%�_x�O��zd�Ml�z�Wd�}�9�#�u��a³F E ���k���s�X0R&/ϳ���5x6���~������ �l�A{Υa�6�nb�#��|y0f���$U�兓�(f2Z/���n �@o6�\32c9;�(@�@<��o �����s��B��9�Ş��,��q��FM]c���5��2���ԩ6���F�i����D�V��I7w;2	$�O8�͸$�lյ��h�m��@�wr��'��7>��=	 �dtƎuzd���@��5�� �ci��8f.K3&y���9c��'�eq�ޙ{ؑI쭈ucYʓ�7�v���L�}�4X3wt��T׎�A ��k8�j�ч}tO��vD����{�.�3�/{����m���s"�	�j�����u���L.�S����,��ǅ��<�.��<�|��v���͹�>$�[9	$��{5��[s'ɋ��S�A9ӐV��(�o&�N�Ce�&�cfcۻ�@�H'6z #{���Ca�6#�v�{ĭ$���r���C_�^�A ��� ���X���gb��T?)d��M�9�T���<��s����ӇTf�Ș��u�֘>3�n��klF�(ܴٙ
!q�q��g�-s.X��v ������w���Bc$.�9g��tM��x9w%�y���l ���f	�$;��OTCe�Jn����Z���C)�;8ftf)�M�j�"I�����,��7���c�fkقI��2ѓ�n���]��{֛!E��m��xX�Zᣇæ}<mk]q�^�1Hh5�_����&i	���n�	���#�Ovu@���9�\�9��#��\�`��F�)�9w`�8S,��2H9B�V�3A�n��xɃ�o=�G�s�gēӌ��i�����\"��L�L��[ !�^K�*$K6�o4L5�W�mm c��o�;s�d�]ֲē�(`��&;e6V�#y�9��$�ٙRސ�;o����& ���!��{w4�Į �;�����������p<)-�Dv\),^�=y���%��{a�BD����H�5FU�H.�Ξz��b�@$�y<�u��� 4K�O�v�D���WH��S\�XE�{�_i���5s�G�Ѷ�N��7%Ǔ-չЏNs�H༮˭v=�>���A�D���_v��D�W�Q ���聞Pܳ��h�i���y.�.g����`�N]:A�d�����_"���<��ٵ O�$����wf���|�O.����t)��ݓ$�뜈 �g���k�3KVH�y�yG���#}A�z ���,]�	��S��z]���5�6H-�3�I'rz#��z1>��/��t5�Do�n��	r��*�Ggey��ky�&V���a}�H�ؙ�A�� �}��DO�}^]W�[g��wƳ ��酼!t����k�� �����Y�n��3��B��	5��^��2�m��2�9�`����7_jH��<O��)��5�msC1v����:��o]�7�ە��X�����Ӯ�8�S-���5�=1=]RMl"u�4��o[��مa��ɷ/G�*,۴y6������gsvz�+�$�h���m�)G�a��^_��gm��s�Bp������͗�y�55��fיw	�:�6y�^�p9%\t �7Y����]Χc�ԒԸ��n�3&�.'����َq���䎷�-�O[���8�'.�d�>�Ӻ�N�Λ�d]̐M��z$�usрc��E�4��ǣ^�f<�'��=
�K"��1)�Q%g45�_��;j�(����1�$�Fud@o$	��D�BQ�}��/���1���@Ψ�����d�4�+�^'��"	%_@RM�Z�F�}�Z�b�"{��x�j���g.�
��l0vW���I�ُ ��j1�_vI�ĕ���r[I's:"�Yr�f�N��Fz  A���'۫ڋ������d:��{�s�w�^�:���2�O[�w��
qs�.:͍��Q��5u`�P�%���$�����_��Ys�c_�μH7Z��+7&N�$�t?5 �ف �v���4O`b�]::i�~��8g��ll�U��)�w`�^Nd��ģ�8��6Y`�߮ZK�&���7��♦񝖇ڨ�����& �l���ǲ1��2|���H�j��M\O��U��@��ɐ5w��ٚ�v޹��E�-�K�`�h�ͭ1�I5�� B�PW9� ��	��z0	�>��ɐH�Ȑ��	�:d�4��ʙ� ���w\F�$��Lzx��ɑ �z�ن|W���m6��D�=��ˊr�]�:�k�̂|I묁�'3��kע� ��i�	��ɐO�ۮ��ni�v;}w�px>�nx��.z�Ò6�ٚ�=��7�z�4�6�.U�c 7�߿�s2X��]����;\"I��Ȓ$m�Dͽ���f�N=�$F��L�߻u[��r�v��
��� ��ڱ�DCy�6�3���2A5u� �ʢ��{h�\�V�1o:vg��?]̒���"95�����ç�O���<:|zzzz�η�h�jhB�^�fzӹ��g���X7������$�G����6	�sk:�w�1]� ���S�܎��+�z0�7Z�e��]���kx5T�s���;����a���#������O�>1Ȳ��xzo�g<ӻ�-Úe����U��{��p�������g�x^�|kwZ/S�V!w�˪���&3,:p�|�G/��;�������=���&=����|09�=��k s���<&�$=�j���tp^������T�NǏ�<^Pbnv{K��og�FA�@_M�.z'ؼFy���Ow�ULi�
��	�2�xX�[�ʭ�S^<�i�''�#Y�%퇠]�SX�{�Vrm��t����P�|�8� Ztȇ� ��{w��~82��DP܋�˽��\ʼ�\���l�m;���yu����B���*���^.s���ՠ/s�v�oz3q��W|�>s�p+<�|�ψ�-U�;�wXں6����4R��N��mX�$8;)��l���z�'|�v�]�ǋ{ݫ�g��}���d�{�❾;����t�����^�$��R�7���51۲=t�}���}����3'���R^`_�����;�I;�yq�=>����V^�r�I��IT��ξ���h.���,i��D�	��Nv/�p�os:����+\˞~�֝�A��/n�%ۛtu�<����!�w�B�{�L��+w_�nxu��H�
#�rRNjy��|6�.x��w�ձ������ؽ�������Uݺr-]f�R�F �z@z��;lvK�{��B;�"
��ݢ��0M�ֱ���[���n�e�M���,��Y����8�q��嶑֍�ܳ�6�g0��8����olH�m��'4ֶ�n��mk2�&�i�$�Y�-�v���4��m�NQp٭IRq�hۅ��f��V�8����Cl&q�Bm�kV���L�[c�l!9e�2rqp��9B3Rv6��m�^ۥ9{d����+"�8'
��8�ks2�˶Zm�9e� ��m�Z![Z:w8NHq�6��޳�v��rLӠ��9�`��E�hδ2¶٢\s4��gi��&k;r�����l�$��u���T��	��M��D]��f����`�iI,�+0�J�/G����I��ɒA ��D+�Yk��3$�3��2b�!��c���|Z���I���z9����~|����F;�H�׀��	�:d�4_�]==�P��jk�*�	�ީ�H;u����z"�͖�����e��l���R�.��O�5\D�n,���ݫ�,���0*�;���jd������7��ܟ<�'ǚ� �I��2�m^�F�^n_^̐A˭�>N��;tC0.�U�k��1��{3�H����Iܭ�� �j0H�*�3�gLn~�䷞�N��K�IL;;0 �v�������;=�|H9��������t1o:vw ���O\�HyX6_b�zE�tA$��z1^Kčj�ى�m:,2���i]&�痽�RO4���S!�������K	�?o~�N�/v	꠫;�R��ӱ�<}'����~���R��֌����t�9.�2N� �l�x�k+�'����_P�k�J���I�WT� ��o�3��/t27i���f,���]�FO�t��L6�m��@��/ ��Kf&�ۋH�h���߼; ��ْ��dt$���8�H���Kn�k9X���{o��e���`�ҝ��v�ª��2O�yE�r7��z N�pͺ�>m��ρ$�μ��6�F��긞�_G[�!��@�.�2c_<A=W}A%eam�H��t�5N�$�׵<G^�D�콀���',
S�#�n��#�o�[��<�	��>��ْ|I���$t�S��\�z6La��]�؂�22*�d ��G�4��M��j�~� �n8�@&oofI$���2gNF���zORǁ��S��/t��ېE�,��D�#��#��y���O��o�����ܢ��U��d��(����ɻ�^s�m�m��|{z��u�g�Rk�6n�;+r;Yê�jcNz0k��v�3{m+�=��WI�3GE�1��'�nws�ݶJ�ֽ;��ٵWD�-�7��q��C�f�����A����b���{e��K�cv�=�.��6BW<�O�T�lQ�)�#�襹�\Z&#����'����5�����hɜKu�2[E��)7��6B�M����c;�m!�g�$y�y`�i�7���`��2�k�z�is�>~�}�|���;@��SF<H��؟>��4)���Sb�x�^H�u�fI�9b\��H3U���L'�5�؏o����H7;� �jrr��t�`��↳�,��8Q!�vdO�5=�A�c�E�=�½�I�_uȒA�������#�-�p"\��<�x�u{���y�  =��	�Y�N�s��ˬ��;ځ�z����bd��J �݋�^@�s��3m�̶��m���}3�H$��	�T�%�Y���jM��F�r]�;j���Z�㧎�n7%�GL"��̱�k�|�Y���;�fd�A�߷��\H$�o+�<H�O@��}̹���67��Aͮ�*��d[IwE��v�ds�g�Fw.K�	H�Lv���I�GZ+�{&���V����a���W<b�8�_��&�j�M� ga�n���ٸ?���;đ�Z�O�T�$�i�5�{�v����QA��%�;$�4�Ϸ�$ue8�AY�&��]��	
j�{؈$������T��gNS;���������jk�O�FD	�,H&�. �I"����c�+1���n����l�!�9.K��@쾸�U�Āiy��l̽N��A+�{/�N�u���΅dg	�0���<�����������70�c��c	����8�C3��gLU�X�	�9	��A�zr`$�Y�P����g��	���m��Έ�X�`*q�:f.\�<�OT�;O��ۡ�	1�=T"�`���ֈPI�޸�Dd��-��豍s��up��N�%r�Q�|k;n$��@�fu`:�L:}�Y4ٕ,��F����x�ֶ����s�F���~#�50���+���
�(�O���n�hT�j1�gJ ��N�8���H@&��ݕ@�ʩ,�!;��f�q��[dec�@4��<���z�� ���S83c ��[�dظ�EgNS;���"@$�ȅ���H�n�#���\�$]tz�~|���<���W�2S�rRd(�.��c���S��P�=������A�Bb�����]n��vn㒟�1��_\zA#n�+ү$���M�S��O���mȝݑ�3� �Stl=�n=lI�ե\�I��3~H�]	!T�˷lj�\�O�-@�:v.��y��,�H7�� ���t���3��$v�\���M�L5N�gi���e����^�-�A��Ȑ	$/�"$�WG�z���b_��_ �,Eu���{��0{��1���+�����t��A����U�w.�Ism�}�!��BN��b��b���DfÛkf��r�	�$C4�ttA��X�yWG��/v	����Out@$����EDb��&Ú� ΋8LSir�ź�2q�nvem�m���cX9�^�y����'p�2	m�DA#b�:8��=����1��|o�`D�M�!t]�I�D��T8�K��tKS圉訐�J<�9�� ��=��֑�gQ��|�MwH�	�ϐv	)�>=;/���A&�\"�!���ϛ���V�	>�q ���	݊tR,��t_d�z#�K��G�Θ�ɷKy-�����
�����&�Y�2!������Y�q wʬ�ޕ>�'ՓQ�}�=o{&|@�_�������]؛���Y.��H�QDƴ>�fՊ�uڧO��맊�S���Oq�}�jS1���H�c�N	mv��l�#ҷ/s�ﴋh������t���#y�YT�̼�gwl��T
�-� M75��K��ɉQ�fݡ%�N�0]���n�Egg�����W2%�I�f�l����[�X��g�ű��C���]@�F�����u���J����YݻWj�cj�[����s�$��G9���M��F ٨E�tq���n���d��$ȔK5,Yv��Q���\�R��ڳڎÙZ�3������y����p�Z�,�.�Dts���>}�x�JBwI�
��	 �Kd/m�dO���j�\_����n"<�:P�t�3�v.ϛ:6do�x�6�ni����|�� �^�O�	o{ H2�����WVsf�ޚg!t]�E�L����ھȐI�Fw4C7Fr�L	��vH�����fs��J`ρ��A������ �w;�d������^�����~"=��؉.��fy�s���$�s+��b_sS��q�5�z��I��ȐO���"��N�+��TS��Ή �Y[�\j�������&J����Cm�]�O~|?4��Y�2!��ZO�՝�My��@�'�|-�d�d�p���L($�wy�>'�*Y���t�� �G@��y��8]�v��s0�M�;S=��O�
w���=>.j�E�E�q���3|���ʺ2����{A_h\���{���u�2X�W+�#��&I ����oX��dB�8�ڵ`�QigN��ùp�[z6d|k�"!�3��
k�]ü[�,�̉�mtA�Vu[93��
t��N;�N��uL�� �ި� A$�z�"z��ź��G[d��Ι'z3���g>A�$�$!b��O�]s�nP�v��{����O�l�H�HGt<{�	3�� ��bŭ�ȒI\����"��v�xD�K��(�kcp�E���7-�e�
i�aJ�3;���%�;̓3��ʌ� J�؂H3�����۽�����s O�˼��ֱ)��w���'9�aޘ���q&���X$���^�}�$�]W	)�|�)c5�s0S�H�ۖ`�	��!�d��D�c���+�9jΦ<'�*)���iݼv�*�&t���2,B�=��??�Ɔ��O{}���P��]6��m4�r���5q��A>7�� �H�� �ć3�&N�ܸS8�:��B�/�Q}皝AUUǠ����u;�:	-�qz��S��:N��`�E�!���=}� �e��VY�"F.���>� O���`�[ݓ%��a]4�Yl��z�͙k,`�nr�K��Wb�B�Z�Eᄃ�I�&��\ߟ<�ĵ�B)K�W���9t�	��ɓ�18ٓ^���׸��6�7T�`�d,:d�Bd��'^��|H;w/�)�����G����ݑ$u�3
�Ž����	�J�lt�ܖ�;���Ct�gnD�Bڶ��}�I�}�7�'*�� A{�2O�,�3�[ɝ�!�F'�dT����h��"�a��ۑ&��&��c��R���Ǎ>�e#�[��������Fp�w��Z}_'�L�$�����c�fネS��:b�LK[E̼ꔕ��>�čw�KUHGY�&᜸S!�cf|IՑqͼ��}�d���^^EU�L�I��"1�8[�"�I�u�;�]p�I�8#�-��ҫrk#�����]�2#q������Gf#c�ͽ�[�ϻ�${\�	��<��Z7 �yv�H�|�`���|��0d�lǟЁ��n��g�8�1��7y�$������z�Z�XwKvO�m;2tBffg��U2	��W@�Iw�	*\�}�y��d���\�\k��䷙�s���G;󒣔�44A�����O�'���N�@�-��Ӊ��������G4�[ɝ�!ڨh��J�>4Տ5�2g��͊��y瞛�.�����������ػ�#�*�����T_�����`U��llf��&ٸ"0"�(�,�2���*,�0���ʋ2"�(�(,ʋ2�̨�,ʋ2��*,��0�̈�(,2��(�,ȋ��(,ʋ0"�(�",2�̨�,0"̨�*,2��2�0��̤��,�̤�̬��!,�L��L����̬��03)0�+0�+03+2��̬�L��L,���̤�0�2�)2�0����(L"� L�ʠL�L(��N�s� !0�
�2��
	0l�.2�eB�0*̊� �;Nʫ6��*,��2���*,�;��,�
,ȋ2��(�,��(���0���
,����*,ʋ2"�(�(,ʋ2�̨�*,��
,��2��(� ��0�̨�(.��;*,ȋ2��(�,ʋ2���(,98����2���
,�+2�̠� ����탎�Û��@DQ
ADf�?>�4�������wD�C�����a�?����_�����Й���?����{~ (��~A�����

��B�(������� r~���4�s��H~�PWW��迓˲C��?�:�� �!;�������a_S
�(�!�*R 
2��B�C �"� �(��� � �,�0���$�����@+����$���0�����c�O�UPQiDR����g�t߷�����P{��c�>��~�B�(����|��M�����͍��r��l}��L~zMϩ���T�>�?��~��<�Q_�T�Oև�C��C����saPW��>c��PAE|��L��i������?�3��n|�$��~�9���@Q[��I�?��'�����T��}�`w���ϖ���po߁���$��?�t8����}�<?���P�
+��A��Hp�5���&�����}���;���a&}|
���'1�=4����u���.�R7�� ���<0`|q�(+��>8��C�O�����)���O� [@l�0(���1-� tJ�
 !B$���aRE�T U
� ( RD��BB�
}�)E � TIR�  6�ԩR64�ZT)@�HT���:aQ%5��P6

փ����ٔQ�%	R"���kDJ �
U�                                               w�Jf2�A�:��/�r�>� ��{:�%�$ �T�U�b# 2��n^�󻩽R@��+�  �_3By�����8 ����d��� �6�|� �hP�����iW��G6{���j �;�J���wP9o   �         ��F��tP6 {e͊(X.`@q� 4Pf{�̀��倢���{QE� ���q�����E�A%UEx  W�7RA���J�� Ehw`�� q�71��݅�5E+ �T2n�v��@�U4��.��|�(B
���  �         ��ɪ���׳I���A�� g�� ��R�/N�R��ԬE�˥5zx �JU��J��Ǫ
Z9�  x��ۖU�1��T� wM5�͸�����"��;��V3��V�M� �͕��W����۫jm��ڷ;�i�/p�m��O� �        ���T�Ý0�]��]۵363��Q����
�����t������弌zÛ=h6W �+�\�w�J�y�p�(T�Z�i#�  ��}gT��8�R�t� n;a[���U.[�fڥ�t�Ϸ/-�fu� {��R��Og�U��j��ҥԚ�t�J���!���  �        }�M��}�*�Lv�ն�uN�b�e)�x ��*�.�t�o;q�Z��δ�m�1ݶ� �Q&l�-B��*�W�%��A_   {׶��ݰ��Z�ZS=� {�[mR�gX�l��1NvUpjq�E^� hGs�ˡ%+-y��Uz��S����� �O�hJR�  E=��U*~��@�A�*��J@  Sޡ�ʩM h2 $ҁM�)P�A����7��h��O���g�1��g��1w��35ny��H@�v�y�P$�	&��BC� IO������$�P$�	"O�>�ϾϾ����=�����~��;w�б_>椭�#K�v�0l�w��Xq��M'r�}�bś��t��j#�Ȧ]�d��v�Y�UݏOK$e��ˢY{F��H�e8��3��{�'�m&��v�1,팝.��[��Isé��L�:#��F��m۱�vo87.O���/;���٦I�+�Jd���!�&�j@�f�C���b���.KP.�;��0j�m�9�F=Ų*�Lzq�t��
*8%X +�6v��F��E�fw]�����qɣPk-b谰����nV���9S++���t<6�F�QS{���g*�*�J�7Z�\�;EC���`�Y�%�6���ǩ@�jѡh����g2�}�w�^HSa��Ƿ[�a�)J:�!�SHS�/H��,�w{�i�]�@7�?�����C׋�s�5�Nľ܍c�l�ͣ���~��mwb�D�N��Z�]S�\�{�*'h�B���l2�9��A���Z勺q�(�6�<�vP� ��u�Xy���AӪ��w�#�g��w"��,�X�i}�↴�̎`KS]��E�r�o
�i�;�P4�6�B����oF�5A�q����
�nG�p�Jh�:*�1�R/��3ܽ{��W�@�c�+m
%y��L���*cV�!$9k1�I��t�3�^�.�s�;q5jY�u8���Ιۥ�l�s\K���C���Kڍ�C^��q��S���U1DL��<U�8,�u�=�����=OW��5�%M{�s���ۓ�z�çW�����|�Rf���U9<�8�F�`���ڕ5\\�H�	���LY�������&�.���=y��n�| �{v�M�,��7&��9>�eS���=�\�^̭f�dPf^Z@[l��jGf�(��ۓ,�{n��۹&�S�7q��E��.�^�H����eNc�/�8��G���X�wZ��2hC�f����^��:v"�Op��	qh$n�{RҌ�&�7+k��n�|kRl8 ���G��U�Y�����#I����`�j�^FĀ};��B��-��ٛ,���sr_D�f��Q4	�	�u��'��JQP��%;5s=�8��r�.�sv��͖�A���*l]�&ɦ[#tl�2��۽�F��RS�jo,x� �R��@x�s���S��<�Krޡ���纡Z���V�k�㯨8����Aw�2ڱ �E��ڊ��9�#\
�"��j�Tޣ��bMEP�r@ƀl�!B��7�+��8��-�u/b��l���	@d�PR����]�u��HͿK�\��a�9z�6��nM����e��)�kV�v!�aѸ6�VK�,d8iu�+�x�
��P����Ww b|lY:C��3����$t=#.˖��;PPs�9]SPݚ.���Bf�l��<vN8f�c^Kd�r+:C�S���G�=d�5�Ԟh{�pe-��[zPʆ-��3E�qT���tJ)ir��
u�A�E�Gq�zy�3��	�D7���v%�-�9�<�43�5��ݢU1l�V��;�}�,"ԶY'F�ai�ս�����Djs�\-���8�ܮ��k��4��*Ԡ��Y:T�a0s�Ū-�v�ۑk[m��w��u��Y�)i�}�s��.,Pj���a=;���+gL;��sDխ��i���:#eo;J��)]�7ش�
v!��4R�2 1�e�WG�������sY�կT ���y�&v�֕�������
C��y��{�(a��M:{k�D5�V	e���;5�p�k �7Hܫ
.;R�n����	k���Ҁ׹3�c����x�Y�۪��1(�|$@�����R:�l9z�&U���&�د�9�3z&�B�M�	�oc+��E#�=1<�:&{l�x��gr`0��8~��2����%43�G�.��>=\5�|3sVh��t�rk��K�T��N�R-k_;%�Q.�&eU�93�A��t.,�4Lt������7��1�]\#�]��H�u�����i1��F�e#oFB��C$Eԣ#R"�
�42[�PnٛR�4��Y�l��v70���ѽR`ɢ<��W�5L���J���*:�2�\�=C��	"�%��@!����&D�����ͽ�C��HN�@�TN»�7V,���֖�3���{1P6�Ö��@�.
���/$�5L``��sm�j	�� �t��ŷ
]��ѯEv�2�����I�>}�]�7D�r�$̜�قl͘{Z5H�����F(w��#o{�������4�@��Vr�N����Cn�J���]ѹ�@S
-�%��OM�2�>����p�<0��̼�:���d����,N/i�[�;7�����6�_a��ќ7js�'Ԉ{Hf�D�}�N�����L�i��	)�o
��.F|K�Yba��]^2Fk��窟nwu�kr�w~ת�d�!B=�A���oX�x��u��A� k	 Ӹ���Ĭ�X�%FjFV��Y�5c$�(gōҾ[��с�Z������&�PD�8�NkcmKM=b�B�tUق�"�Ô�3�y�F�Αl���6�W'y�=���0�4i�L�n�-V�=Cdb|���a|�j�#�ܴ�;�a���^Z�T�y=a�����Ao�˵>'�8��;mx��M��z�ŝ{sq[�p%9zt�:�������S��ȟdU׈�f�7)��C:o1N�Wږ̙��3���h��@c�9r5iD�a��邡��2�&)lY8B��ѹ:	���.��aPʕ4�{,`7��nu�N�������3_#]����v�3��I������x͒:��P�.c�]�3f�6�;��^")�2�u�у-�r�:���R��PZ󱅯y�'@��P�����v��&n.��WJ�z�DH��/ov��70�������5���O��N���nq��²\.��3"h��������N�����l]��a�^�}^�Ak�r
���'�+��1�ӛ��8^�gf�j����{��RnG''�ձu��$����c�^s���;�k�e��3G�wcLo(���%��uֽ�`b���~����.����QǇ�{�Ԏ���Aȉ�l�y��E3�͊v/��������M�F��X�,���f����Y��a\{��t�ݮ�N���n��{v(�]��-�Z��-�Q��vc��h�꩔7yc���h��M��Y0��M׳ f^nTY��"f2�S��9�M	��nW8��f���>*滭�shg�Ub�ݓ`, �M��F�ɜ��~�'���8e<%	C�]���Z����/s��N£j�$⛝�&\�X�����C�,_7�3�!ǥ�YW�=�/����H3���׃l�8x����: �ws�U�P9�;�1��{mZ$��8\�n��2k�ᮍ��X_L�p赘�ć��5$G�w��NP�A�;�QV�w�+$]̏6ZF`�:N�G;��K�e���ȯZ�a�e��׸X3���nq���;Ʊ÷-ĕ�g��)�(R�ǦjG��ɲP�I�S�>q�b ��T���23�:5�X�гz��>ğ�x^��$��O�ӷ�1��;s���GZ,͎A���(��j3��EDD��:Y��<*��@��<D���TvL�wo>m�׍R��ߍ�!�!'�2��!�n⡠ơ��"��.��V����Hp,��8�di�Gn6p��k��p49ٺw�{VN��.:�v�Q�2�#�e�+�H���K���9Z]�Kd������r�q֎��a�ry���d�;�:rt�-|����FL����(�mю&�eX��Q�p�)9ln�5�"��\�v=�C�F9Aӷ�:Dt�\����,�7�-e�׬�'c˽��S��0r��&Î�N�%�M�\8�x�wע�������;��KsrCs��t9��ɬf�Ցȝı����o�CR�������Oo1@ou y��捺�h7�Œ�,��b�`ȹ��`8t�y�q��y;;�I�C����j��ӭ���z����	݃��ћ����/GU�OF,U�P'��ΤN^�s6�D��7W�6�r�1�K�2s)w'm��t�v#��㼚"f�$�������L�/� �@�!�õ�Sʅ<R�����zC��1scov}h�.`x[�vI�uWՎ2\԰gld<XI���9��X�D*{D�b�V+���)�����N�a��o�v=�E#o/m���y�;��rH�����ײ�h�v�cr�۱r$��E������p]NY�%b�vgs5��0Bɟ<�tF��<q3�L&]m;�S��ne�ױ׉<�6����i�^C�<#5��^��-DTz�pⲄ�G�e{݅���8�L�$�ۈ��݊{�Ph�+X��n,՜�\e��ky��hp�Σ���S;u7%�ؔ�ovؓU#��S��]��S��y>��&H�+�'e0�f�b�c!ы��c���DNs��-�/
�w\�z�X`���YQ,���˯�Unjse2N�o]\KӲ���/_�zG1c�e��m�5i�͜�q����##��;��$���۬fY�h�y��nsIrQR������r�Յ'Ɩ��l��e�����A��}��e��].�׻,�y����J��}�$;3Ձ����Fi�&.I�qR|�TGnp@���ܚ�j�$ۇqV@��ݱ�0��Kf�;��:��jE\S�$��~b���1I�ź.:�n�-uf'�4]ccd�߷��:�FJw��C�V�>Ń]F�]K��[a�[�e8�v�oJG|�u ޘyS��t��J|��؜����k�+b�4eewEn��)�ר`��4)!��]�Rc���� �Ev7�ˎnUG#���!�F��������$v���fLeJN3q�̙4�kޚ�$��2��nqh�g&#{(�c[�U:��}�v�M���g�/�n��]�
��4c���:��z)p�z��
P�S��:�v�aLd�B��m�Wd�z�b�2a�ii��l�:8w�7*G��z��򐒽�XQ��<ߢvE+��H�BrM�7�nLg��3yE$�̫�.I�%�'c(g	Xs�<�����޸K��pnV��B#�\� 9S��\��7q�hZ���A*�7-�rvB5ZՀ��s���	-Q������]C��5�vj�^o;��@옉Co>taj����'Q��2���T��DZ^��-\�a'T�w����Zy��t%�oYӉ�;Gc4���9�6[�;MU�&�sc(��a��$�����2�d܃U�D�S�Y��u��Ô�iv�<Q9�4�tՑ��Ԗ���]# ɷ4)m�I{V������R{��.��0���x��z�z+��v%�JFq}x�6��W��S�4��zF�7������Y�ax�s՚�d��3A�h�����c�V4�97MxzJT-��]��:��!��C���[+*�u4���Ujm�k)s�8�˗fc��2�')��8-Q�0���Z��8�ˎ��.�f��[4r�2�t�t��ff�pi-0D��f��3���\L�Z	���ؖ�3�W&7����[�-���Ԭ����f�m��Ȟ����n��E�>j���(U�#��1.'�?Z��_���MC��`�ĵ��U�t�����U���xs6�r��n��]z%����q�����C�7a(�x ��nD���L:ջ ���i4�CE�J�v�ݰ��P�ܗR2q5nc��B$��Dî�mn�7�*N�ޣL �����Է�.Sp]<i��&��%my��ӹpgiɡ7�o"{)�	�dY���/��bK�H�ɸ���WM9�I����X�Y�s��C���!:���dwu���F����B��g��[�4��T"sYʼ���\��+$��=-�av�-��r�io:l����H�Zs�)q�Xsp�t�W�p����vmh9uU�����9CGc��H0n�cV����a�p i�ˠN��91^�kmA^��<��q��f�����g\c�Ƨd��0sm˩��;��J톔0f�4��ό�S\43�:n�'�$Q�Y��m� �����^]�k�N�B�h�V3c�4���k1���R"X:���n���fbSPl\h�#��m���:^��&+�ۻ  %F. �XЄ-e��L���է�+�t=`mY
W(�G�8�d�(d| �@�
��u;������&Ccc+�T䳃�׺�m�J����%<�JI�p���Bh�:Yr����!�LP����,m�K��Yx��˓����:�\:Kǎ��Ӓ�p�;���Bĭ�	�`r�X�Yr�UA"�����T�7v!�{���.�sgk�A���t�t��=2�7�Ur� %v���t5;t��a��ҫ�ی�>��u���;�qY3�&��B0���d'3m��@Z'W��		�
�$XB)
I	O�`�P�(H ��d�E����E�Y"�B)  � �$�"�*HP!"��)	 �	"��@�R@��BE�B�B@V  �E��@�d P,�B,����
�$Y Y  �HB��$$��XI$X ��RVHHVHT �J�"�R !d,!*d�
��$��Y�$
BI�	 ,����J�BE��!"��� V
�����@�$�HH$�@XI%dT�
�IY	H,�P�
� P 
BJ� �$
��B�IR?�$�����$���{'����5~a�Vse'Ċa����#��U��,�;կ)�%��g�kp�ܭ��Z�t<����LSՃ�4���9�����ıI{V"8O.	��gs�<���(VVW��ec:��}V�2K���t����Sa9Ǳ'8�cz���;���^!X�G �6�%����z�Lݫ�ȡ�]��:w���OY��l�$��e���<�5��%8���Ѯ�Q�bR��*��zf��XU��Zta�R�)8�{��0� �\x��[ۘ�}��%�C}t�_;W׏E����E��m��JƯ,�0�6����VhNd	W�����U�$��H�S��۹��Wfs��M�qU� �|�L�7�nx�oE�ׁ���&\�`y��Yjħ��O����v�>|�x�tLQu��Ӕ�[a�r����"��nóP.�Y�:Ѿ��!�M-��C){%�6�u_m�~�׸��}�!��t˩[/P��=�[��|�-JgMRX"Cw�J;�l���&`��K�Ѷ��թ���Cm/�#��L��z���Y��o^�$�V/\]7��wN=|r���1������Q�Ⱥ��]Us�"r�p�E�1��iC��p�H0h�$��U��JR�U\���UTu�;;���yPcY2��s\:͛��c,� �&P�ee�^�Y�y�s��{^L�{n�֝ka	ݺ�*Uy;��f��ϲot5�7�<���l�U�|"+�h�!�N���7\�m3�� 8��p��6z�Gar�4�o�d�	ޣSN�Y�ڨ�����#�fv�=_.<зN
q8��̼�B�̷�Ρ�9�R�B��ƳE��������;�^?���ϸ���⺕�΋�����T���:!e�Yu3��ڴ�l�>���o�յN�<9�5�}���0�`�z�i�f��4��'�Ifi�+	��7�u�y˙޶D���Im��Z���}��c=����S��5Ǵ�V�>�ס5�J���.b0���5uK���uq��]��k��ϣ��ܕ�K�#�ЊP�ٸ������B]��As�FµM�Lʲ������Y�9\�>����GsArk_AAʖ��\���ͳ�|n1ד�#N�;W?Gó&.�䨭Br�!���uz����2	St��ưe���o^ۍ����;����NFB^�L�6b��<�8{]����Z�M�Gw�0J;��f)��oN[��Ɩ�ѢwV�.{���Þ��a��½��Fx�������Yˑ8�ēx�Z���ـ�y�7�Or��Ɲ%�سz[���>����k�8��ܢ0,�$L]��ef�e59Pc��6��˜����__bU��Kn����ո�s�l���7:��h��(��9b�'v7�é�I��8G`�x}��;���I���g�V�hR�s�,ɂ�;#�r��u��uK5OB/m��{�s����0�N���wc�r�Q�Nl&7<S�^jl�+��������;��dB|&>iܶ�:�Is',Q�]j�Tm�m<���8;*_qrU�)�{#e ��[/��������-��߼^LzvS�j�� �U�T���C-�]��r�l����������mުe��b�b/.x9������=�k#׭�G�* /��	W��R⽢�:ڝ6��
�b�1uE.��m=�.�8_A�Z����#:�\�(^�G;W�֕cy}���N�qLc3�k�_tߥvn9���:����YzH�R"�fN-�y�LNsC�j�����0��:��݁G�	Sn�G��P�d���p��%dԾj\�=��yxN]�RzhE#�.-U�1��.���{��RYu��P1�Qk�vSQƂ��k�I~�/F�hСﯯ��9s�����oz�u��&�-=Y`+x�"z�͖�ݑ%���#�"^�N���o+3�W��X��<����oe��k}'w��	�Ė��r�������}|��r�`�'oa�\�uk�����ၰRK;7qL�V
���W���"���u|�R�M��M�䏤`��Q�x1�u,�E��Мm]�oV{�a��l����z�_/2��H,,��ƀ�5*�cėq�)�KƖm��o���s�qs���M�t����y)$[���-����Y7�����-P2g�3'r�`��m��2�\��7<��qF��J7��Ab��}3G\&��zQ���SO��O];l��y�9���+w&7�=5$�+6@qN�Z:a�o�qGB���Q�]��b�j*7bz��K�!���<��z=Κ;���zytvh
�E���X3�˰�[�GB�f%���4l|��^S'U떐$0R�4�$��
/�f�\�����Li�k��Ç�܍�yO��x�g��p!p�;rV%Wk�e{N���aQ$�סͼ��2�nJ�x��0
��l�Q�=�f̥��I?j�'�c9�q����K�԰��W�̾=�fAۛ\;�c���5�x��c(Z�XC�i����J�rN����iG��[�{Tz�"u�0����'X�w�-C���:3�|�h�->9C35��omjz��]��ˣ����ئ���Ke��f�2FYԲ�C��Ǡ(��d��(��N;b�b��Ĳ�	Ě�rw�>�X,V^駻h���&;���)t�Ժ��`���l���6n���o.J��j�;]��o��Ip	v̶��:��EG<��\{q>Ďs��נwI�E�8.�'Q�b-�n5�ʧa�WY��紻���ݗ�$�G�l�}�ۮ���󠑱��U�`�&�}p{J񻝼�h_�Ji�67\/jm��n�Cb�E�0j;�.lÅ�}����}K';�z��mv����%�N����q��W�);�ZѾ�c�U�#b�L�d�vѾRY��$i�5�N/�by���ܪ�3��soV�䯤�VgR����ܤ	���Zk,��37z��T������rvB~=sԼ��幾^G�=fl�5y����I>>f�9H�S�l	�2ߚ�����9�|��p
ۻ�~�x-�h�m�����8�.�|xJ�u���������������ê��2*6�;��s�;fA&\P^ٙ �uN�I��V�uw��p�/^���i�u�P*�q�i�%a"�c�Z9\�/z�S��Sj�z0��"��]њ�F�Lj����,�����:�9ֻ���h���{����i�O�9�ɳ.�V{=�NE�9f-��"̡�Q�����N��u�Ҩ���n��U�cep�����ɽ��ż��#���x�9؅Y8V�~�И���h!Cz�0��_uݲ�X�CBi��Aa*r[Q	�x%X��g<š���m3��ʂy��K�T� ���f#[�I�V�^b�.�<ҘG{㷞�J��C�T`�φ᱃��v��@(��	pq*y���q����{=�]�_��t\�r�0u:��4gPZ�a�B�F�a�8�����΀QΡoz�YZ#;����9���|�E� �u�مk)cLS8ʴƎ.�rG��F^�+Ѩm�w&��4���V��뻯�u��Z����U�iR�R/Lj��?G�J��۫�N���Y�>I���m:��̷'<����{�mP6��{Gc���\8 \K��'OZ�x(�}����6
�:I�\���;;\T)���E�v�#6&Q!ԛ�eӜ�9�u�U�l!X}�3@9�����W|��1��v2�1n�8��f�\���{]�fx7�hq�e�V�,r<�i�E�=W�*����o���2+2�em�|�7�����;��R�4�$)κ�C�h���� mP{�Z8�v��X��x�X�iO�a�!�6���T=Q����Z�����e󭙧�� G�m����b�.�k�}ɮڗ;�81�0��ٱ:�r\Y�mՐ���4�_���ʇmSg��xws{L��`����K��t�8�3Y��/��4kk:j�A�˽b�Q}��bVj] ��l'�Le[��Pf@A�Av�ˡ��8�2V�*:]+b�F�>R�XR�\pu�}�X����:��<o\_�ɧ*]�+�{=]��F����2���,M1i-L%����"�s�3��쬒՘hz&/O9̓&�~�s�Ą�S���Iа�||�w�UG��ص�������kY�K�ڸ5�rb�}��hbީ���t7w3_5��{���ݾUj)�q䪡����ea<7K�t̽hvc�lY�	Ş^���B)���{���j׹b��\�+ta�Nt�%��{���v%��7j���Uݕ�JA�^���N�v}tC6�Êobe��X%]��{3'��v�i��h�/nV�E��zuy��o.L�d蛥��H�6Vi6K�d�T[Afتtcי���ܞh������1�,��ݻ�wУ�w�\evޛ��x���j l�zK�F(�x`�6`h���q*�߶.��&v��W	�&(r#���Tt��k���z���tV����r;f!��������j,�p��qm��y�V�wg{�3�$�����(��t�G.6�^����W����м��^��<g��_��9��0�ow5���[��P&:ha��ܨ3��D�Q}h;r����KD�\:��չ,6{�1��_o����;������XGI�Z��&\�fQ�!����7s¸,��R�-���]t32Xsw�r���]��K�#�j6#�;Qmʝ/��9%�f��*l(]��:#á����;�{́���)p��c����;��*�c�`��m���L6ʆ��IC���G������D}������vL
��� 1;��V�53Be�[o��ᓦ&�.�H�,^�Xے�]�5�9�l��x9��A���ϥ�7��ju�e��e7��c]����飆[|�:g@�[�������zQ���8]��s�${R	�~��3���C�-%��3����D#A��f\��*�rv��{n<���c�{E��g��=������{Lsy7$Se��\:k���mҡ	J	��3:k�ӹz�ݢ��կÍw;VOT��xGx���I�}=�3��{pW{ ����s�M9���h��٫њ�wG�Oo�W|{�=U�n���v���vWv�h:fvwfq�p=��O����f;�PY�n�Ay�{`�!�XFc]�p���.v�8��=K������X ���LYf]g;�%],��=�m�oSܚ�ʅժ6�_FX���2n>���J�u#j���;Ic��ufk5�!L$��X��b y�A�sD]$��.�_^̉����-҅n���.�:�1�S?A��X��؊(%�;k��B���)����Cڼ�ƌ�C3�8oBԔ����N�r���"�'m���ZK�(2���m�m+2>�/�	�;ow\�P�㊢9YZ2�����M��T;�zՍ�J��Ȓo:t��W���[T]��/nܑ���ID5�|��G7&a��\���Eruy2"�C��9��gs��4I�=�|�'�Y�\Ѭ��� 9��Ȕ�`� �'7;f�&-�wq.m'iOv�<��OvD�^��-,�^y,�Ǭ���f�s���}�R{�mu\����{Gw#�&]*�%eL�c��HKG��t@���]tM�}/� Q���<h�V�rL���=�3c${���ʙ���1��:N����7+��K��R���o�'֛;gA�u�cRվ�]c�A#�"o�<�J�/��/�
FЖ1�(�PD�v�n�ӻ��ק���g��9gt�ScQg]d�9��)���U��6r��޳�
���o3�o���'C	����3��ԇ^��,P�U��CS�^R�R��ڳ�/�ɛ�Ĝ9��R�R��D��i�@;qf� Qq<�Z��wu-)�j=�w0��lF�Ƣ�r�gm�}v(� �#�'�hE[���Z@�v��ܸB�Q�AVǆ1]a�����v\B��snx�E�9 sPĪ+&������/M+5�Pm0[������Z���ӛ8-+~w��6Z&-�����%��%�<.�g[o�!��;�jrs��wbt�욵�����*	4��=ݍt��
ܹ�`�t��u����w���xeܡ�?gU��F{�rU���3/�b: f}4�59��U����3���s�ώr��r�B�d8�>�n��ϗ
��m≫Ќ�E��6��B������p�w4>�NK������6�[1�3�q��e��Q��j��U�"c��͇�f3��Li��'yM�$����lʽȷp�uR���/�����+��c�K���L&�53�S�3=X6P��.����|��ב����@�%Cb��+����4�e!]>7��ovpY����Z[(
����؄1p�3��;��\"�o�y�Zږ��{Vz\��w��ȟ����p�#��^m
H��^�᱗Ϧ�)0:���J!�n��=���d��L�WaךKīH��s>N�\���{7
�:.UfI��Z&A��͉�V�d�J��V��^�h�S�2e�-{�ق;rT ����p|K�ٸ~�ݒy�+6�.«�A��p���5N%{�>���&v���D�uκQ`w�Qe�w�c�-un��cK�q4eFWt� �Ns��q�ud�s{/H�a�V�^.
�:%[�SŽ��Li�EΫ3��L!�0���Ǿ+Y�ֹ�6 ����� <9�;D�We��̻ܮѪ�jVx�O�����&Ћ���I�{{У��jn�p���H@�p�I�]pnrb��՗��h�v���d�hWu���ka��粔Y5���5<s�w$g �lqێ֍2�;��]9z��0�z.s���m��v	���G�݇�N4v��Ӻ.�wh�4��NM� ��Q�&�����˸�\�jx��u���8�����Em�,o1�B���n,&э�<ԱĶ��N^�e|^w'�����.�^Y�:����ݷul�uV��p<�ni3�n؄�T۝ۮ@1/=l\G=cnNJ�vSu뛯*����(��:�m봱��;iɋv�ۤ-��������-��d�9N�
�9�������
��b�^��6�$�]�|�c���{vp)��9.������Wl��]n��c����++�wv9x�[u�w]M���S�갸LS�����۫�<6{R�ӛ�:�<&��y7/.�rrym���ۣmnud݌C۶�=����;�G;<��c�����j�Y9����uܡ�\{���cn���t㝠�1B��s���J��cv�ju��m��c�Xμ�dqK��K��A��g��-^y�J�2�k�"���m��
�7c���E�x���{k)��)Ϸ:������(���g�D�uŷ����"筛uX�]�b���C\m�k$�:x�rI�W���.��8y�]�W>y��^���2Q��+�����p�N:u�f�kU8�#re�뇑�v�Y�[69*�Ep��+�7:1��G]��r��{{1ex�t+K/=;�:7����o`�n;!�\'`��h��n�ݬd���:��W\�XW[3-ǣůvn����í�q��lJyueu�q�u����
+n�2c�\��me�4{X�@'hQغ(��{]�<�m�e�����-�Қ9�j�ӗ*n��,V,s\n��n�����j�g���]C��˻q��Z�i8�6�� s�y#�����d�t`7�%�ǭX��L(����:�9]�a�V�.�|b�� ��L+ݑ������0����p�u�Y�F�'���/&Խ��;��x��<mO^�<�mv�ƶ��P��>2l���g"<��>u����@�u�U��n���l�V4�%7j<=\/d�Pn4M�On5�e��՞n�׈w���Zkq�i����8����=^�h�"��׶��C�훱�f{u�;b#h���f�����/ ��ӭ���٧�cot�:���Dsj����j��{cp�t�v(}�;�f�XZ��t��8��`�1���=�g@J��GnP�g���D</���/g�gq��kl^Ar��^Sl��%�����u�^;��N���$��\s��^�\n���7�lvvۂ�u��1�Ȧ��;\��z��ݎ>r灶�=�rq�׏NѮj��ҹ��I�V�F�U�r1�]��6��/]M��;V�"�]lflg7�f�ەʽ�q�[N�0����v	d���ؑ�X{�7qWD��p��۲1���n6��<\NcN���=���n�m�=Z]�ʧ Sv����<�]�#SAv;�qg��]��s�\srGR�"�g�@�;��ո�{g\8񝳹l��4.{4��lQ��:Սh��`y�l�[�+�t�ņ�]�x�m����ǩ1��1m�zS<v�.�;��-��m���a(Lrn�f�7\���+/���s@v��&�Hvݷ�ڀm��蜠
�v��m�Z�F۝t��<N1��T���U��y�Lv=X�&8���Gh�WY�*枹Â���q�n`D���sؘM�vh퓨9 .�:��[`yܴ�9���1n:s�gva�k��ssF-�I�vQ��ۤ�$!���k :"9�o;�nմBv����S��f�t�!t�s2�,>Q�y9�oh�x<v����ڶ� ݑ�s�����]�yp
v���lJqq�v�� um��NzČ��g��ݝڭ���{g�/����-ڮ7g��<8^f�gm�,�<��ln����ۡ�����#ug�M���9��kEaٮ*z�9�����[;tޞպ����GTsF��n�X��;B{>�e�C����P���Y3��咷V.q ��mV�d��d��ݮ$�k����y.�����'%ۋ<s6��d�^66�6�F�td���wA���;��=7:+�X�:w�WRv;����`7bu��đ����o9	��8J ��)���[�vY�NǠql�;�P%�]s9�;�n�o1�v��]f�C*^����R��0y��su�w[������g���	Lv���.:cwcq�=�c�e캷-�6r헉]�s����y����꓀�OK�{�=��E�F<�+�*���Oc���"�[;ƷX��bX.<��xպ�z�l�;Mjv�÷3Yힻm��qXx��8<��;r��ұ��sgx�Ӈ=�;�<���^������luV��n!���[��"8�x\�v�Z��v.�gy��=����2vn�l�^�Y�=;.�V��Tt��ޭ�}M���f6X;v����ݺvqŅ��wے�M��^�S7n�wg�pk�^���d�N݉J콎t�mt��^�r�kJ{�M�g�F�/i�ն�Y�j6�q�c%��<�Y���)u�㌗R�V�d�����e�Dv��Ck��i����k\n����N���qc���v���{��h�x��W�;n��t��[�qq�63Թ+v�NMr��b��S��F�p��vN�P9sl�.	�IxNt�K�ێч�h.5�j�Ÿ�W5O`7uY��{�Q=��r���*��뒂,�[e�#[�wg���m�۷j���;v�I�F�[e����;<r\qΔ4��Ee�]�93��Y�	�y3�����n-��>}r���g[.G0 \����m�� ����@XJ��om�
n����[����n��;��v:�϶����n��\����v1գ��ك��.�v3�v��Y=��w�9�n��ul7kl��卸.ޠ�<���EkrU�m\q��kݣ��cv��9����X3���Q�pr@+�x��n�8����ۊx���۸1��.LL�񋴆�A<�;+��-�A8�>w6'r�[�݅z�n���d�:�=��+Z�����؀���B���mX��㝇�v�v�OKٸ�v�l�����8�[�a.H5��K����٫�z}6��mcj��U��{{Ԣy��n=U��2z=������A=���ݎ�ȳ�+s]�RTʔ�gx��umǝ�p�l��jv7�،;��s�k��X�f�Wa�tY��W�Xp�l
i�5͜�rQ��qmo�`�S�����
t�4$:�<���xK��$v�'[�K�U�힜j�<�,���N�m��@�����z��r<���Q�:�),8��=�V7mj����>lV;p�fbص��mŮ�v.�;�ǐ�y�	�B�g��G�u �y��n�-�qȜ��.�u�lrvȉڏ,��7	h�*&�/��;�v����i:wV�.��:��d�G��q�ܗM^����izìYt��]�l��`"�
^z������E�1�S�װy^6]��토�@v�^T�z^�m��I����n�p��C�A೙���^ۢ=�=�α��쇞.��sve��g��0��F�n�s�#�n��#ty3�9ć:��5q�;�mn��Nz��h���E^E]�C��U.�m��x��G=��{�<����WF�mu��q�m=.y�Cv���n�%��!�^�ƴ�m1�d����;������ݰ`2�nhժ�y�<��S�xk��wn�0�w��
�ɫ���|x���A�(�m��[;p�2.;v�ݎ�f�c�trmn:���s����㵚#Wm�z5�=��ؗ��\�g��l�v_�g��ȋ�ܘ2EX�t�h�T�O9ػW9ݞwNS�^p�Dv��6϶�����pRͶ��];�ݮ��dV�s�ny����/���1�8#W�:�݌ۮ3�yRm̵C�Mٺ��9ݣ�##��;C�P��-��k�#U�ϔ4�����y|�����
�Er�Yl�i�6�ݪ�]��i��o4F�4�eXQ7��գO��r��r�#�c��-�g@�I#��X۔�:s�c��{\���zg���ص�a�c4���'F��\��:����4�O��k�\� ��ԓ�7E��z��kl��$����cWl�+�zų�u�۟Q����7:��$����v�v���2;n19�v�jP�z�h&t�������`k]gav{gc���l
����+�l=��%7Y�Eѷ`�|pcj�^�NWn8Y;v+n�r�w9�v�.����<���q��n=[��r]N��U����[u��h��/f��Y�č��'��n:).�c�'1cnNqѷ.I���cgR�/b+j^�[����s͛m��;	�[��n�����t`�cxmǠ�.��\8�������Z�N)uht�uZ��O6��d�;8&�7lc���{mݹ��;N&Ƌ�ѝ��k{&L�s�m����n��ab�'����U��e�n��D�:����9(��1#�76a�p'i���T�N� ���R��p������2�\��L9�u�6���qd
k�m�����q�l�84��<-���I���7V��w2˒-�^��d�:Ӌ��!�ssk��Ŋ^3l�i��d�l���N��]:�v����-��#썪(գd�)�v:z�+�]�>�'�u��d��A�˳L\t�M�}=H�v��|�N���z:ls�H����$���g)�iøu۱��p��kʝ%�ϭڭU�7��hx�)�ܤt>ݱ���[���n��+�s�yٳq���&x��Y.�Ï]v�]���9���9��d��[���&��p������sX�ɶ��{��8���<p'����	R��+EPEb�AEU�QZ�V�DE��+l�()AEUHTQ`���mAb���H��PR*(�
ETV11E�jUA@��Q�T�ň���5(�1X���PAeJ �UAEH�(,Q�J�(�Q�"���1b�ʪ"2*���dR"
dcm�D�QQ�R��"�Q�Ԋ(�V�EZ�U��"A�"�(0RDAEUc""�TV�AEUU ��U���"E��(,PPE`�X��RҪ���mhQB�DAE!Y
�b$UUPQV"#"�D"�QUciQAAcl���E�����PX�Ȋ�EV+�����Q
*Ȩ�UE(��cE�1DdU Ċ(�EH�,Y-�ȌUV1`���TQADE#hQY�
E"�* ("1X*�V�b( �P#�Z���AE`,QdĒH�X�p�P�c<�gnxۣ����a�lS;�-ӡ8�����G��%z�R��y�n�]"�ȧ��֌�/���vxS�v3�^N�
�e箷[3/fǫ��6��vrsZ.��7m������a�n8Ku$�u��cr�q�f+��#c�ɸy�7���;��_Vn��-���9�ZmOr��<=�e]=T��*9�i����������GHrh��=��nۅ�n����6ݵ�@���l�����
�n7�b�v���˸9#��Q�-��=�r%�=8�<;�E\f�=�/r���<�J�T�n
�\k��:�W=����x����KX�}�{%�z���k�n��s�ۃ/�+m��,�� d�����b�Nxx�;$�����v6+�3��8֛�J�����v��(���<�v�|�6��:��q�#�w����儴S�띳y/I�-���݇�퇵<v�N��m��(�㰯cg�p���6�8��D-��.��u�"7m�7@a燧{85]�u��X�g��c���
��x-Q�ɱ�}�1x�xpJ�[Q�jSf��[n���=�u��Z�N){,��Gn���wϛr��7&(�t��İ�e�]cr�nӛn.��ѻN�J�w		0iNl8�m�7LCp���j�
�c:���dt�ML;��:u��t�b�r��%�E�ހmm3;��^N��y�4��;8�g';�b�m����r:ε�oi��q����n�=��6��`�kN�.�C�q�)����nۍ�^F�nW��8�^��!�\�n7v��ۃ�.��!t��)š�sWs������s��٦[	�ձ�9��9�J2Z�m<�^K����r�a�p�N}�)�\g9|d���]��.t�z�e�l>�͇vU��c�dǝ�eQu@z�;/*�g�ƙ�㞊����x�7ic2y��M���`ܶd^��]Z�{����r�ďs�<����zB��yC�.�F*g�.��h�y����%q==�s�RCKu�w�g�zF���H�0��=�7 $P�H+<)��
.��
�����p2Q(\$�����OGP�t�34�>��:�.�7q��y�p��rM���=O%�0O1ǂz|^���Y��n�!Y����?��%H�l�B/�d���7{n|�|�.�W�ڋd>��~b���]�wv��E��"M���P!?u
?yř�{���Awvݓ� ���AI���'� ν��_���'J�(d��{%J�zM����X��a�+�|�~'����F��Q��g�i�,B�u6���Y��r�r��Az�n ���w�񝞛����b�;YO^u�$w�R�R.8n���@��{�����]e��t��W[�(��IA�c�01- r�J�9Ed&l�N{F�U���Q�^��oO`M0�c�Z+�n!��������
�����ܻ ��ڢ>!_{�.��:�:�M�e�]}B�Ʃ��:���Z�f�{�����X�z{D:��f��̎���A��"�,Gu�쮩A�������Y�r*u�Uj앴:����[R��ޒ&� �l>�g]�˯P��`�=%�8��"��l���~5�K&ą��8^�Q��yb��1 �J/�v��&��u�R���Nr��Ɉ��U����Q;��ρ ���D�O˽yv?��B��'�V_P�XN���"X�G+�y��I �omXذ�0z��$�ҁo�.�'w�n��B*o�%���V4^���_D"&P%��z�Ů��܇/G!����0C*F�k�^ѝ$�8Q��v�P�I^����	����ݵqv�w3ez����^]�H�gh!Pbp�՟���#}�mo���v
 ��g^݂Iݝb����m��jԾ�/>��T�A��0�-J�u=�dgv��>y$����exn��R+{��{w\�WG3��F�����!�1N��o\� D�o�Y�����u������N� �E�y�VVu�n����ﴘ�U��X$����d�3gȸA�c���a#v�#5r��.�VH��u� ���k�1֙��G6�n�۔_݋p�!���_u�$;*�b��ّⓍH��AY���@T)���]}ٞ�#�~5�6��8�� "G>�4�mg��t�jvZS���6�>�a��vǲ{���TtD��
�_�q���~&gT�`��%"����L��v��f����ӜK*�f��7`�vzP'8?K�X��=�޲H'�s��$DΪ	��,�!�y���}��<�ϩ�J�n*ڙ�`�O�OuAFUY�C6��w� ��:�&uP��T�L�n0��߻��vz�q �����H5�R����,��u��Oe����>�Y5��3{�V-t3v*�����{nL�δ�i6;&�sq��L�T=h�t�T�x����v ϙp���� K}�$��,\C�G�z���
_]�`�ܦ(|Hw��w^nc;�0B��F�nB�a�*���qM�vK^����9�k�7hA;�����:���z{f���� (��H���;��%sޕ �X���1���YHS /�e؛=����D�[2r"��o�$�k+HW[�`��F���;�=;8o�e�b�-�D����W��$��^�A�Y��~����A �z�h?�W]�`2�~%7`�����cOY���ך��m���Y�I��y�rj��b�"�K�����[+��r�?NϬ�;����0��5�ȡxM�څ��n�]���ڰo�F�R5��\�U�H������kS�܉��dh�y�ю��w�n�����0�eo�+�ֻ�r�ͬj���� ` η�)}��%��tf��t6ґ��D��!�J)��ۓ6��<������mv9�9��w[��nE��-�ݐ�ܽ%������l[��� `��v��6���KF���](q������::�6��|��O�s���S����{c�����u���^w%�y{Tl��̄]�F�ўz����۱c����6��nw˶��s�6ugع=�k�!���\[���gc���g��7o6����x��pt����t�ǝn�`x�n�u=�\s�������cp��������I+����w��{;��،�w������?�'��R�T���ܕ�ⷣ]�C�n�d�Jν� ������hv��y��do�RR3SEh�l�{6�P��ʰH$�j����[cΛ�̜��I+z���;��v	+�!n$eH�Ϗ^�g�dZD���%���	��]�I�Wg�kB�3�:�2�U�B�yg⚈�Y��B>�?Q�uLO���8�����}VI?{{�v?�ww��-l���,��� ��Amͅ�[�6w��:z6k@AEɄ�BD����BC��Xh=�H
F)���u}ݽt8�tYa�7-w*$�/k���P�����>�y��1�Ha�c��/�Be-0O�x]L�a���wT��ތ��iuh��^t���u�\�w�F�	�ę���g��c-��e���E,��0:���}P|H$n�zł~�֪�zP����gvL�����w�	��L���޺�H�U��<�s#�k�������	'�H5�uFXj������)F�<z��2�ǿ�5�ޯ�~�u��$��{�Z����7<*}���T��HF�tiԬ�5�@���B�5����ww�'�~3�m	 )���\���D�lȡ��룫8�7FQ�+��F-�t��&��۱�9��$8�2�7��[Q��J8�zo�������~�IC�U��Ykq׳� ��~7�hW��J%�$���Y;����^P̞��@
�SM�
��X�§mvP�fV1�`�����$.��A?��5*~��ɇМ�j�����^c4��b.>����t���4���n�td�yT��W1�;z�
[����Ǥԧ����E�t��	�۞��>�V��H	�a(�Ha�ػ����~��~!�]�$���VA����b ���G����!řL׋V�Bڌ���J���,�~=�������vBF��T	���$nnu�&�����져��j������画*�֜�Z��Bu���ڞf��:H�q���ڵ��6�0�ԏ?�W����:A@_v��V;����tŘyՃ���	^�˲V�a�u^����>�=1�;j�̘� ��?�f�]�I��7s�7�{�b���邙i>-�
M�vmߺŐI�nuX �v
�q[}�^x��� ��\�
1���,2apQ�{�D>~�C�������:@ ��J����*-�朶-y�N��f5[
Xff��'���Z:�]��y{���U�Cش�ͪw��(}�o�<�!ċ���Vj�t�|�����X�/wE�Y,8n�z@ �~3o�g�9�*|7={p f�]�I �+�m_y��ݤs}�5���v���9�҆8xq;��ӎ2q����\6P"8���F�,#$Pf���A'���,E�Tx�n�ɀ���u�ē�wg]�@�;�R�JmH���W��g�h���I'7��Y?�}L-'��wkQ���s8,����2GO{�@(T�=h ��Z�b7������O�	�z�y��Q*�"�%"�	�<�U������8����
�g�X�z�Nr�X}�p'���vE�s��-Lj
 Ƚ��&<��iB�¤cS����E�_P`���C�� ���W9��[��;������hЃ�+�_���B�Ɂ|��pC"����c��*�9���̸l���Lv����������J��ԛ��]�;���^��X��%��	��O'@Qk��"l�;��2���N��\��=c��N�
}p�ϕl���ھN��7��ۓ��:�;y��c�F�vFXW��j��z���*R���n��H�[2�<M�c�z�q�x4���-����l��:z;j69�K|�tm��ϭU��C�9A�9�g��[m��{�v�9pv�n�V\p�v��cu�p�ۦs��Z�ܼ�j�;���?U�`���ՙ�����m� �w��;5����ߤ�(��<o먄#���XFH�/;,X֎���X]om�w�O��z�c�u�"
�g3�#뮤��c�N�m$�R�6��L�	��Bwx���*�9~�$�oU�	1�u�!c:0����2GA�g�R9\=ϱ�͖�&5X����`Nn�_��G��')��$��UG�Xi�$X�\�3/�@ޞ�:�����,+OP ��I@���+pN�I��%^6(����0�q15�m���[m��#�l���Ea���Uy��8I���2/m2O�<ݻ �s����/(����>���|c�uY`W^$�-��U�����֐��/�W����߲��7yl�]�t�Ʊ(!�LG��Nw�4|���֬?{q����j����kӀ����ړV�Ђ��wب �ݕ��|ӌ�ٓ��襌�5Z�T��7����o��`�{z���O�����Wf�#�;r+�	���'�ݾ���3� �f�hٕ�7;M�g<�`|��I';���$A�W��U�~ԯ��� =����8M��h�#�������DE����p)��73�o舍�}v$W+�lu��ł�K+�6J\��y��[g*�ۮM��%�pnC�ֻ�{�m�MaD�ټӤ$�y"�) ��̽���}i���׽���s����f��O�W�Bq�S7"�S?�D��i�(���+���Tp��GR7ݵݹ^$ &ަ�mɐ]��w��$�\��������t[�p���,�ܹ�\�Ǯ�ˋR���#��]�V�h���#�b�ܖ^��f��v�\�n��כ�,��Z�^�{��W�Մ�o�Y�x6��Y�A��tN�*��CW�o^�������ޅDb�[gvK��f޷C�={�:ُ�Zz�q�w�g"�\� �7�5}<dJ��{�$�����l��B�T����Ec��t������]���3ڡV_a��+iॹ�WX��=���e���f{��y�{�/B������"�s���Z[�7��f��D����W�V�9�"�A9À޻"��f�}����-,�Lx������ʸڰ�9�Y���3Nb�]�:���u1#;��c�aKN-�{O��[o����WJV�v�o���F��yh�k6�7����u�{GD9]�S�����]d�HU�9ܣ/�ǳ����8}�=�W ��Ld)�5 �m�𗶌p�"l_A��\�G�{�)!�7n�������@t��B��/�!~��<΀�'�W���X��W��AI�F�N���*_o�z��ݓGIg�My��WW�s�XZ����{x�ugܼ}�4�]��+ٺ����#Ӆ��}F�^a�1IZC��*ɨ_@X<���;]��<�&[���ri��u���̱4��%����pŋrVm>���B��y������gi�s{4g9���J�A�4.�:uR�[���kvY6�j�en�l����n9�Mag=�_o��������C=�F�<���v]��ǡ[n��n�c�������(���`[AX�1���
�H,�
���(�#b�V����QQQ�TX����
",�,����E�IX���EX�)b�)Y*"EX���jQU��EX)"��QH�
��PX�`��
�V$X)(�IPYQ��dP��!��F,U-
�X�TPF,�+�"�+U�
H��AX��dT"�E-(
���F+!YR,PX�UD����h�KAh����b�5�Tjڢ��`�0m+"�U"��"�X�YPU��b
�"�TUD*�QU�H��F,+DH,X,�"2)UTb�UUT�����T�DE$D��,-��`,Fҫ�AZ�#���EPX�,Q�Z�ł"��Q�(*�E(,PR,U@P#�#1�W	���$�ޠ��^F5% Bᒾ>���*f47Y}^� W��l
>���&,~އ@���I@V�ځ2i��M���_�}@�/��!���o��u�O��\�������m���Jn��"Q��M!H�O8-�ϱ^�)t��u�^m�e�.�ۈGg�����~����!��mV��^[t�ē��w�:�~�=ޝ5b�ee�'�H5�n�K�%�@���BfzJ�Y������Py��VI$�\��Hs�.�'����e{W�����񕜡H�	���F�<�%�Ͱ,��uk��*rw��믘$�;�����6�iɐ]oz\�D9�p;�����pP�{�]b0�:*rU��L��tru�q�͡3	�쑞Щr��p�`��G����hS=;����Ź�X��S-��6ꚣ~�#��@3�1P���Ƥ�@\2Q�w��A�޺�l=�]�[Z��
�Z�7T�<θP�wbq��g`����\�C
O�h����C���LZ��r���qӺ�m�k��ȑY��������e�4mOq̴ ��s�T����o�a'.mKt=+>3e?����a�$((�r<�����T���-�Ն�h��@s7lY#w�����d�r,5�ұ����\EF̡Wy]��=�]VH$|C���i�k}��w�|OĹ��`{z��^;rF�LD�h�����;U������ou�� �ۛ�Ĵ(�s|��J���I�I���� �G�T��7/s&���$���X�{z�*P�?[�9��"�
K���!^17.��|y״��I�L���#��Y�m�@���QpC�e,`b��ȧ���*vf�EM�wd�X�
�2�� ������u��X,���N��;��:8�>|�(��6�ñ�+e�t�7:ۋ�u�ጽU]'��l��C���J�ᳮ��O!��ƻ�m���v�g��5�mSm�Gq����S���ty��z��y���e��#�;sZ;k��7��&��wVw��sj	��l���-۫��6{;.쭜ll��q������ۙ�3��4���e�ѵ���(���v��7nwv�Y��n�����uc���4�K�#f�#��?�?�R��L��Y$ݮ��I��(���|��0�	0{�{e�� �ͮ�$�RI�"8˒;�Fw�B����{4q�ּ�������d�I��� �{�z3fuga-o���8�mW�ş�ӫ�?O]nضq�:�޼ �=�]v���!�M&���J6eٿ{�p4;ǯjs�ګ� �k�%|IS�+������UfE�g]����4�f&�_J�]��η���j�>����������ۯ���3��Hv۵od�8�Qe:��p��Xҁu�l���&�^8�nwM��[��xݡ�O��E��	� �_e��'���ʢB���vR����3&b��ސ
�Y�����L�&��;`�����<�܊I7w/sWs+��HJ�GdY%�M�TA>�'�޺��#�U�
�]��Ւ��XRp�������r����_�e_ě��l��=Zt�'^MK8J�)6�m��+ݙX *�ʰ@#r��G�ݳli��:��IWvط���q�#�"�k���ܻ�{�z��đ*�U{v��H��|�5U��ƹ0����4��棅(ٔ+/����޸=��Ka��>�����  ��;�$s6'����A����ݙ����-�2�zu�b�Gu�%�%ڟk(����������}D�U��{guX����Qw���l�~�	*�:쐀����h��p�l례��s�Wv�Kjh$�[v�뿉"��;�sj��Il�#6�_�Vbh�EĈ�� n��Y$����p����-2�8f:.�c&U��_
4�(]��������4�oDo�Yf��-��ۏ�o�|}%m����������_zJ�������˘H���H$�?t�Գ�I�[l���6n�ml='��v��dٵ�v	����{��WW�ƒ�/.�%`z<b#�&*K����B��;뷣~:4@���9���'2��� ��]B�~�z�__��߉דF���u̍���e�Z�q�&Rm��vY[���(#���>���'X]F��	�~�@��]J �t�;��Ke�y�ͮ)�π��ސg�����M X��3�)q�{A�a��B������]����o������q�d�ʁD����H,5�F����@�A�H_}�y����󌏏��~�>H/�C��|`��\e�''=�{G�����h�&��%B�+Ϻ>�{��o�g����%��}��9�����ߵ(����k�5$� !���m �g�ε�sՁ�ԅ����h�)aHV�o����M�*e����je�j�ߟ�Ӷ�����j����Z�M\� ��G��;2��v��_f�iR�x8�7��y�l�;��%ǙK���oY���I�:�P�C����C�+�_����S.r���U������J!RT+o���pg.�-���w�_�P(������ q*A`V���j�H6R�����8�_����S��v�ӎ��DN��*hwk0h����հI�^�˖ b"�,��ja_ѡF"1	\9Ǡa=���~�Ă�FJ�W�9�d�%B�%aLo�{p�A�`���οC�K����ĜB�VVJ2���jM��)�l�.��m�7;8�Ĭ9�7�0+R�;�9���[��ލ�R�B��[{�{p4�� �������������{�>��C��ߛ��lQ�J�Ɯ��#�u�����T�B�������2VT�v�?o�ɧ�{��~8��+��Z�����t�JB�o�{P���\���߇R�1�P6�s��q=}�v�?�}�g*A_��z6ɴ��V����0�0�(¤�N����$��y����~�M��w�j�6o}u\O��6�3�;2����7�}���F�)h���/8�w�k=���9�~�������=�M�(�YdLo����q��,C��=��r	+k��/Mw8���/ۼ�5�%��4D\&�\��KG	*s�`�T�^��i^�.w���\�^�\�������z0\�Kx� w�L��{���>��_���4�Q�`dG�.<��o;`������S�u��;+�u$�����H�Z�*[�8N:��ur<u2�i�ې���D����Q����:=���v��9M�����`�W e�N�O�FƘ���������c'
�c�uq�;�u���m�OGD�v:�;�c<�u[��WNt��`��\V�lmgB`�S����9;��X{nL��6�٦�v獎�|��~GVݴ����;���M��ק�UǣjEư<������W_ڗ%�\��!Ԃ��s��a����+o���m��ʁD������r%`~��g�S߽�g�������@�� �B�����Co#�������3\9��a6$����ND
�2Vc��������O���ގ��B�*IXS���8�R
N'{�{Gq
�G�~����}e�*�}E������Pm���V�tm ����G�
H(��{F�)
���5����Ƽ~�߳�O�*T
ʘ߾���q��w����ĕ�1�ǿf�9�nG8���'�`��y����ika��] ��I�*Aa����83��@���{g�Xk��{P;O�~��Ʊ����� ��-���jx��2m|[�)�w�Ĝ�9�ND
�++%}yϴm�H?��ߟ�������IXSZ�{�q ��¤����q'��ed�+��{P2��c�|�G��߽�����oC� �Y�8�\�7�񮵓���w���n6a#����p'�2Ɉ0��� <%a�~��<`Q�h���!l�*Ai�s����*c�k�~���8�����$pd�Q���G����ƿu�./�.�9øq�#.�P�>�֮t�����^�qp�雐�:s[{\�IZ�bmK����^��sV��8o&z:W����� ��r*��v�ֱt�NLaxa��u_�	<a���چ�?�T
����l���{y�jR�B�g���+�p���چ�
�<k������n7�ĝ��~����Y`�YFJ��ߴm�HPIP�J÷w{�3���1�{�����#
�����Ĝ�VJ2�VW�����i>����q�XL�@#��׿P�P���\k�`djB��w���H<)
сZw�ہ��J�YS��jgߴs�����翎}'Y�2T(������pIX\c3���s�V�s�����
���la��!RT+o�wGq�?�h����A@��߽�hJ��H+�\��ot�JB���wچ�0+~��K�y�͊#���,H��YO�QL�[��T�̜aN�kE��s���������`�9���<����h�q��VQ���ϴm�i
$�)���$��z��}�w�i&�~���$� �Pe^�jM��)���q=�Ynp��ve �zo�4�E��;����P� ���C~)
�Z�����n�h,+*c��C��2T���޿8��ߜgr?_��P�|G�����C~L(wp�0�����i&Щ,B���~��G���$�.���oS���:��?J��;һ'v��˥�+L������P7�|3��߱Yu��W�tr�T!:�+���`�z��L�{ݮ퟿�@������?�� �u��@�� �o���<`V����-��,�n� ����P�?˯�6��:7�u �ђ�w�6ɴ��IX\k�}�q ��aRQ=���I�{8�;����n���2��c*����6�@�=��o�q�X,� �{=}@x��
5!B�?}��F�H\�?��{���1�W��{P4�*X�YDƹ��g#%ed��}�������3L���U����5ls=y巷��WV7����`t�r�7E������Í�W����u�#�jO�~�U��wA��i,B��
������d������8��+���߿}�Y�w��_{l5~η�H)e�5Ͻ�q���C�_�V�L�k�N$��h�p@�����[�?3�䟗y�I���ƽ���0�*v�~��>��'��f����O��T��hk}tc�ķ8p�;2��+k��P��R�=�{�6�yHV�+��o��ߵ��G�}u���}*Ae���8�Y�J��}�h��+
{o~..)���Lg7p�*��~�w;���;�s�2� ���3���8�YR
��}�i�ư(��w��	_��Nr]gH��&�햫)6NP��*]0�&���s��cAyw���^�,�<w`'���=[ڲ�f�	���_f~�����|W������s����W���|<|�"�r5���Q�6$��sG�ed����jP�y�����͘��C�+���ۇpaXQ�IS��}��9�����Ww����M o�[����[y}��)�:9s�r���ۋ���[(���s�m�k��c���a65��	���0��?ۭ���
A@���R���s�_�2>�yX��!�� ���[^��x��*AB�;���8�X[����)����\�P�>W{�=���)(�IϽ��=���c��q�d���@�{}�� pJ��jAy�oځ��)���1���v���P���[2mun0��L����N��=����� ��7��a��X����p��u���C��
�RX�{}��$N+%^w���e���{qf3��X�|	�z~�?t������|O�P(���c�y��򐴤*Ahs�߷	���eLk�}�q����^sc���f�J��~߽�C�J������⟥�rc��q�~�7�P0�hT�B�ƿ~��3��]�{{���R����ҠSw�l�A`p�^}��P0�wHZXc_��C�d�~z�Ln��w�)X�7x�T�y���!vB����NiL�:.��=���v2���^��ώ������H�%|���/��z�v���5�&�v�V7n�b����q:�0b��$ns���6��0",2F��+ڻ��ë�)w��:�᫫E��;+<f��lU���~#:I�ZĲFJ��C�$\���ːo��u��|F{��S�`�����8+Y�R�U�Ξp�X�NwN��A��;ݦ�˯ɕ������joV`�e�z��ņ�o��,��S7���3U9��6'iWǇ�(��6�\�wJ�s�T��<(�=�^��:���=���h�3�Թ(��U�ȉ)���1��'�&��hwS�9J�2�f��wj]!� ܕ�ӥe�Y����GB��j����^cP��
\�ފ���:�(6��ӼA*��@MX�+w��]X���Ln͌�7$��"�a��
�=�~�W��q�ip*�	ő3Y�.Qmx5�b�=����Ʒ���J#�b�V���,dT���&6�u;>m	�����5z4>$���zr��ѱ$Eh�r��7}ҝr=�;�vu�P+\S9`K���Y������ʞ�]0Jߎ�c�ջef�t緑휝3��v��k"�ftk��X��_L��[�����Y̼�����ً��{��^Ռ�Rr���1������n`�q��Y�y�����YI|��Ȉ�ǻ�a���c ;=�9��{����C�Og7HKw�ZGKs���M/l,ծ��S���O�"�yJ�EQH�� b���*�(,�[,cQb2
)�1�ڊ�+F#Ab6�[H,�Ab�Q��R,EE~��ŋX%�A`�Pc �F(�DA) �����ᕐQQFH*���X����Y�+"X�,AV
��(ᢂ�EX���X�J�Y��$XEPPD�Y���b�T���TP�"��R"
�,�V*�UE�R(
�`*���E�AAATEX,�X* )c1j��PF�QC�
��)TdE`�,���
�*
1c�PQA��E"�b�$Q`���Qb�"�QE�
#X8�"�F(.5�%��Rĕ�Q��Rq��n��#�6�x��̅۝���͋(�7+]Lm��M����&:m��8Zts���퓭A;�/j�Eh�����Ocv\r�x��:�緡��u���=�w竮�sx�ͯ,K=";�h��nݻ��`�͆��-��O���=���9��B\�t�َ��zR�c]���].5BX:��g��\]��-�V�s�8�����s��ݛ�s1�v�oG`�w/m������{;W;���08��:���R��g��Z��"��9�k6�7q�cq��[�=]����2�Ƚ���К�{Z�N�m�d�*1[����R����3��iT�͞�wZ]7��1sێM�N�r�s����p���^<�苠6����lv+m�+Xv��ێp�cм�n��u�^�����7I��pt$�S�pmN�&ݞ�ݶz�vJ髱����װn̼t[��ż�OVۡv�FQ؍���)ř.�/!vϞ�+{������p�\6�vN�ۙzҽ���\;�ƕ�n��Og*s2{pu���d�ʑ�q��7�[�C���&�g)l�VS���w1Hc+�v����g��3�Z�<%;��f�Jَܼ{>tgtjlNoQ"�`{�	s�9�y��b���r���cluaQڍb�u��\�uث�@V��Q�z�\;n8���=������=nɏV;l�.�XR7���ۓ���m�5%c��m'h���$g�[��n�˘e��WW=\4s\���k����뺌i�lG68&���=��^��Ԣ3�m��Q��5qt�z6ݍ[Z�71�n�1Х�IE�v^��w2m'�lڻUՋ�'&�7��y�kqW&��MU�$ݮ�1�H�;������li�z��pn�s�w�[�P`�v�;g�[n���l�[���<`����g��;P�����e�}���z�9��YQ��	��OZYx��c�:�c9i<<�);��M��V+�ת��e����m����f���;������O�⼛`��ۡ�Nt�nM�y7��%�vJl�Ƅpcin�vܽ�=]obw]�Fe���66k�M�f���u�u��.wg��mz��v��$,E!�qZ/[�:���������vy��n�Gnv-��C<�=��S���q��R:�2)��ٛ��٫n5]��ˇh��;te|d��M��Nݩ[�^;���<��Yn�{�۰�;g���tvc]����N�f���]�S{8��:�ۥ�e��]�Z����O��:]�ӯ��)�	5���'
�+(�_߱���d�AH,)����0�aXg[����Yƻ�ӟ��N�s߹�I�!R%�w�}��! /�Uk	3�7 l��� r%a��o����~s�����iu�@��ߴm ����w���n T��7�����pd�����g�g䧀�_�����J��q"�\b�:�H.u��A�R
J�a�����g+*J��oG���g�}�w/�ky�O q+��`׿���s4�iK����q �4����S92n�N��=����ޯ}���>��d���F�2��*%aw���p�F�T�O����Ęξ��e���;��ƺ&FVJ2��7�I����i���$M����!�������+R�>����!g��?���ސ뱁[9�y��a7*Ae�����3���d�{�����%a�����fO����L�m�jvN��cGLv����ݻ[Ӧ��w �[�k��a^u�7��������y�E�za��������T��y�����$
��w��� q+_��c>�z}޾}���gޠn�HZ�����x��>�z��F4�"��@Ͻ��m>+(�Y������uo�O=��0�K6���g�	���F��%���Iw]��/�PU�R�u���a��3��۸wD�����xG"%�VFNs;��q�߳�ߟ� C�M:�?wP0��y�����aXQ�ID�����Ă����]��k��q�i���I�$ �_�-�ͨ�h�,x�=��3.����Z��h����򐶐�����o�ǝ����o�����}�m����d�w���������BJjK�#�~տ�@z�׽�o;��7<��ЅIA
ß��q�d���@����� pJ���
y}�ځ���p�������H6R�����8�`V�?m�~.0��L�����߷�h�p@������������A�}o���]�/ֿ�Aa���~�8Ì+
¤�}�o�8��B�Q����/��Rn&�������������kWn���X�3Ŏkgc��1��\[Gn:{3/���Y,�_�0^�̊$ğ��+󿻨m���hw����R�B�`V�c���M�T�>�q�o�s�?9�,O����8�FJ�*�w~Ѵ�Ý�o��q��.w0�
�{��a��!Rkܟ~�^��~0��}�GY�KR
�}�l�"T��W���@ٺA��������{~1i�C����<�`V���ۛnDɓ8�>��Ѵ�@��d�����c&Щ*IX2Nk�}|��a��y��Ϸu~����TY5�m�/<�$���GU�j��`�+�h'>�(���-�gw������]�}����عq}@!��^����*w����Ă��VK^{ܟ}`� ��X,��ƚ),x�<L?~߹�}���y������`e�
��~�to�!iHV�
Ӟ����؁R�
ʚ�}�C�d�k����=v^M�C�I�g�ԛd.�}�Ì+qq�I�w�2��;���w;o]ӆ�u�n�:��T
}�ݜ@���Z��y������-�ֽ��x0+�����O�?�Ͽ����� 5��[[�B�Ok�����64�qH�`��	!�^G�M�b����I�����'
�R���&�&�
%af��wp�0�=���w��}���O�����Ĝ�VJ��FW����`d �_�0zԊ$Ė(�,��s��q��!�{g�s�s?��o�7���`V��ߵi��+k�q���J�7����c����yCG��_�e����&2Կ����W�~�Cl6�Rk߾��q��T�wg�m�׾����*A`Q�=��������Zﻨq��}�_��cr&L����)��^����֜}}�����6βVX�^����d�%H,.����8Ã
�ID��ߴqU��G��=�8	�x�S���'>��/gm�g(tw�6�S�v��U�1���:�۷R�c<U��9Zp61Q\�泅u����y�@���'�ʐ_�{�@���p&_g�m3�H,9��oP�AH(~�_�7�R��������`V�c?~���eֽ�u3�%e�%B��{�h�IXg5^�e�q���dB�,�
?H"e1��$�x�uݩ�*c���b'+��Jf��w�����ɕ�1����WW}���$�T��V��wGq���T��w~�Ă�����;��`xk��}�H;�-,5����ǌ
��r��q�8�L����M�����@��%g�8�$�/�oF�4�R
k>�w0�
�RT�{�h�Ad�ed�?g������6�??���I�i[�����spg4����yϽ���jB�@�}�h�)
�Z0+��|��1�c=�;Ϡe:�R�V���6�FJ�*}��G�٩�[�Qڗ��u~�@ �Lz��w�?}���*���wG#8�YR
=�o�8�Ĭ
��u}�j}ëO^c�� �X}�>��ǀ���y���܉�.q�
n$��4q8�YFJ�]_����id�������G��m����w��a��ac
���{~�Ĝ��ed�+��~���*�Uva��Y����8�^��ݯ��[6�YA=���+|��n>��}��j�:S1j�ޘ���hx���{�ǞS�K�P�4�[��������?Sﾹ�ٮ9<�M���kr�M�5/&������lek���0��n�Qs;��q7�6N[��cv�;;�l���\��0�W��H;��QC��3Q��㱮��R����6�k���9�=j�ԗ;��1v�����ݹ�*a�tv��1i�K�1�7[���c��=ٙ��F���G��dW:�8�z��=��T����m��	��-{=];\i��ʸK<Y��W��j��U�875��g,V�s�Q0�c�mm3�H,9��z��F�,��w~ѾJBҐ�`V��)�
��������Z�9L�_�VhM����q�++%A7_� x���'B��%�%°�º�?{A�I`�I���F��o����~a~�~�6�P?%@�����$�^�=�3H6��ɟ���������)��乔ٍ �N$޹�h�AgJ�J����62e
����_w��y�s�5�:��
°�*~�^��$�!Y(��Y\���az�`��qs���.6i ��7��;����tn�� �{�������l`W?���q��}�Cl�?}�#���?$3=�����q%aw���0��Le�1s�q�W�c\�$؅IP�5�~�G�d��o��������:��*�o�8��*A`X�=�>��l)l5�{���#[���eWqߎ{BBD����C��kO>ݎ^T+X�O.NS\l��u��ݸ5�>~��ܫ�3�z��?w߿h�q�Q����wF�L�RT,IX]g����aXw�;矿}�}�m��������d��ϱ��&�e������ki����?~�����h���'�������\b�w��6��v��&bƭ�Gtb������f,�-�ta�is�x��`=�Ȟ|�Ь������s��&����ѿ�H[HV�+f}��p0�@�A������g+(2T.��5�������v����>�+
c9|��櫜�\c��Xm�u�s��2��RT+g���m ����X?s[5{�{�m �F����P7�A����Y���q�`V���Z�lƌ_�x� G����<D�U����3��YY+��}�!�� �����nH,9Tg��F�{=�?w���\��~d���FW|�=�6�@�_�1�"\���V(�,�~�ޯ���Ƥ(Z���F�R�q�DM�H-���ہ��J�YSY��ڇ9*��}�i�;�=��u��{���S�t�]��Yꗊunݩ�ZqZ�mȫۅ�\�E� L��A���Ȑ��������
���c���Ib��߾���2VT
����Ѵ%`}{��5��w���r��k�c��s4�il5�����[>�����5r`�q��SbO}�~���H,߳�X���$��q�ځ�8��D���}��Ì8°�
���}�h�Ad�+'~��`ǳݟ��L��>��e���}�mmÝ�@�J����惑��H[@�����H[HV�+�����M|��Nn�k|ױ��]�/?CNFA���NIRj�%{�]v<���gԘ��E�-j�X"�k(�*K)R�>����u������G�ߟ����@�����ڇ8�P������8$�,�s�w�\�̗�w
�\���~5�_�?~�RtB��V�=���%e@�T����q �8���ߵ������c�zAĤ-,1�o��0+L���{��e��ɸN$�7�h�r VX�YY+�ch�ɔ9|{{�1���뾓��9�����aXQ�Ib}���8�����VV~w�����=W��C�c?~�=��ކvz��F-q��+]! r=���/uK��e�j���x��o�u�Q��f"��(�?��w����jB����F�H[HT��>���M�T��_�~�/{����{�ڇ�J��P�׽�C�%atw�c&13��w0�a_��sA�IP�0k�/6�}�:?v�o�����P�'P,J�}���8�Ĭ
5�F��7�@�A�!q���^{:Ʊ���|8��P�ڰ'd8�01w�������� ���j�%H,7�{c���̹γ�C��T�｣i8!Y++%��}��Rn&P(�m"K\�E"�2ǈ�#�����2{����ٯ��x�kmH[@׾��7�R��?���q�>4*���V�g�y�BG�c��joQ���ɳ墳DˡS�ph���^o3�o���i0~(���ϵ��¦��9W��]2*��NR��iz:O4�>�������H(}���h�Vc?j�s�.nfK�g;�a����h60�J!RPB��}����2{f���:�{��v~@ؕ����H,H.{��P7�A����~��ǌ
��?8�w\�{����x�<}a�˃���[��g����[��郭�Pa�椅��"��s\�NL~���7����$r2VQ���7���L�*J��g�{p�+���M�_�$�{�}��8VJ2�Q�ϝ����D �_�>1�\��\6(�,%a�s�h8<H)�����u��_�tw�����![#���P0�@�P+(�Ͼ���pd�cۭ��3��%w�����?
�2�S�
l�Cl80��ƹ���)* ��}��9�KP*Tw]�p��{�1�o�%H)��oځ�����Xk=������V��	�f6�E�"�'���h�k��������?�ld�����k�72�R���w$����}�h�N����5ߎ�d�ed�+�uu��-�Hy@�A&e�������0(ԅ@����7�B�ɮ{�����{�}�]0+q�y��a6 T��5���P�82VPd�Qw}��!Ȓ��5�{�����>�pr�ⱗt],����?7����L�1��W���]���vwR}�d�U���^u��i�ɳ6�9Q��,��nyK���{�����>��pƺNW�s�ݵ;��u���+����hψC�&l�&����n0ێ"��mk����e�y8�$�n5�q���Y�γ�=h�m���z��/[m��&���ngI�gOmv�ŕh�gڮ̼��:H�^{\�"��2��5��s�%ǳ��뵱N��8�v��������6�����I�]�g����4�i݆}]����q�tx}�]c]GZ75�-�v�cn^�������k�1��?�0�������2�RT+g�{���d�*A@����@�V�s~��Mw�s��ߘ�~�>ޠa �Y��ڇFl��b��1�+�&�q8$�s�8�*Ag3͟����:�5��|�x��>2�R���na���*J'{�{Gr!Y++&}����9�����oz��2����<���g8r\eѤ�a�o��px��H(�����R��\��Y������k߱��0��,@��������J�2T*�y�C�J�G��$W�H���N>X�|����ҋ����ϖ$�%�;�s�83��P,��s�8�ȕ�cXk��~����ߩu�w��;:A�HZX}�sڇ	��<�t؍��G_ H�Gߧ��#�
�2VX�]����c&�}�����^��|�XY߷��Ì8°��@���h�N������jM�������~]�������^0�ӓ=�����i�fr#�Iѧv�n�.�e�b������܍\b��%a������
C��~�y��!iHV�
�x��nR
j�n��g�,�����8�R
���F��J��g�{s��73�8�7
�q�4����~���?��=?Vc�jKo�V�����j�S��0+I>�vם���3�*Ý�o`�J��]�e� b�(1�uW9�<{�=�/�0 �0�������w���6�X��]�{��oT�i����hZ���|#s+�A�P�q�}�$\9\�w��&������e++%w}��@�ACbJ�~�y���kF���?Cl:°�*J'��=��8�d�����jM��
k|u왫�g2\e٤Ĭ3�{Aþ�����1�o���H[@�����HZR�
�x�����m����ｨm�o�������{%g*C�yϴqD�������ŮL�d�1�p�A~��5)>B�?��ҧ,�`���[��}$X�e�����Ʀy{�yf'wꇂ	�� �$�.ۤ�N3�=��y�w.ا��������}�?}KX���F;�{�vOăG��D�����arλ�����:J�7�uL.���DA����>�}wZ�a� ��1^���$X�ʁ�λ�Ei�U׶6t���k��fD،��e.��C�ο��IO�b����F�ܲ�vo2����쥕��Gz���-�1V� )�>���m�k��y�C����{Y{{]v~y1�6�&L��`���}Y���g|7Q|�<�q�_�f緽t�H��?9i.+�,�7��v]��[�ق��ٚ�vp[ٹ�l�˰o�����I
�[;�m�;��9�V���A�4W$��{+F���g�ۈÝ�"��s��}P��Hu��+z��ͫ�S�:Pl�pK�:7f`=8���<��;�`n��RI���^ѽ0�N�I�����N��M܇��[�������z���X6����e��Ў3ս')e�db��ø��[\ͺ8�򰈞웼���pi�N#*Wvfi�o{v��/�1q���)��u���Z�{����Y�"�F�>�n;�2@�ub���N��C<�0�J��g��5�ص������n�����w�}p�]���-�#ʕƧ��IRW}���NlF���c(u�������[�5g^�,��hU�����һs�Y��[[�M�T��y��gP�wG=C�2�I:�V-���6e��u��|S���GnZ
�<��)���;�0�u�$�z�L<��ԁ�KB���˛�,���NN�JG�m(m �MV+^vf�x:�nvc ��T�*m�V��sz�Vrę`�ܤ9lZ��7K޺C=�ڧG�1㚖p��`�����WcBD5Vf���PH_gWa�'cd�u�y��±AH�XEX�H�EU���`��A#��"ŐR(",�AQU]�|�a�`(�(**EX��d	Z�"������(�(�@X"EEQEX���
(*őE�J�@(�0X��U#��!�V"�H�6��Pm+�+YUH�UŢ�E��F"
�E�b0Q�@U�B��ň�*@���R#P`��H,F
"((��QX
1��QA�*�,YAT�
%kRT
ʑF*E�H�TUQb�F*�U�
Ă (
H�"��8J8B�T�V(ȌE�1E?��9��u��5��1�~��)���y�$�i�%_^z.��gM��9�L�����O�nu�'�۷�����wVyb�`|��c�x�!&�2��6����%бK��V@l���ĂC���Q���Qc���;]�ն�60�\���OC�l�gyD�ޫi�	�u�i�^����Ē�(Y�ki5�����C��� ����x����@��t�O���';���LD\-#�:��Rv*XJ�|I����}ސ �uB���3ں���G��$�Pr	�� ���U�O�oP�8nͯS��$9}�`���f�]��f�#1��f8�|a��ۚ��y�*��� nwz@�>�I@P���3����{pb��ݞ3<x���ޙ�����gLr�r=K3�B {�fe���)b�Έ�h��2�Kt�����iu�����ؙq���}_}$��S��}���f���ۃ.q��f����D=�Q��w����`'kz��?2f��?Y޺��w�bX�g�8��d��P�0�^��j�B
�ϸx��<� �q<��Lځd{�y��"�l3�7/6ł^�������Et,��&�qg��T�� �(��&�P0�i�cU���R��jy�j�vn ��y��d���LGxm�3QX_a�N�����}�ʧ
R@mU�z�
X}/�@%�V��9U��v�^�u��^�����~"���I&��+��B�����;F07n���� W��l ��u�븼n��&�I	1�d
6����T��W�׳��թ�l�S�hy�y2@ ��V��} �Y�~���k�W�/lR٬������
rV������ݒogk�ˡaÑU�i �u��g\c����3���|>[���$�-n��Sk���X��Ŭ.��y��9[�Y�8�g:�#�S���A�z�s�Gv���P^��i*q�q�%'Z���6cq�Ea�[�F�sk�s�ϳq=�pk�F#����'Pq���e5���8u��mGmȫ	ǎ)���v[eF��90�۝� ���˴��;z��ܝ��M���"urQuk�c��Nrr�c����ky�=&�$1ok���������ۮ6�=�lmGn��!�#IZ9���8��u�v	�v*�g�H'�]�v0�4dk+7�<;g]�'�~=e|�U����nFLf'@ܼ꿊�]~�^éʫ'�~$duʉWgW�zA�l��{�/�6�E�N�ڳʁ ��ʲ8jF����1�t� �f��U���o9��D��wm����>B�w�\�W�]2AU�۲I�r����q��&ye�̍g>"���I&��+;Ղ��[�`���0���`M]���-wl�P����z<#.�S�T?e��$�.��,�\s�����E���&&Qnx;	���Dx�-�I���I �ٷ���o��>��E.���mX%��cI�c�݊��]���|-w�t�4ݎƚ���-�זƙ��,��x�}�ܕ�'R��p#F�v�����}��eP��T��2�6o��}��b�H'��o������#��}K9Ǎ�A�sM����@�A]v�@=�]VI�V,�4Ner�A"�wX���ޫ$1��6b08�r�����*�U-?u�$�J$S_t� :��ν �wg�Z�~���`7� I�R.1��T0���WSԹ�^-���ݫ�v�cq
#=]�8��__ό�z7~��,=,Fm,�RR���N����%�A��l�eQ����s��<lpp�?�߀����J&f���˳�ٽW� �z�r�*����y`U{2�	�����
�-� m�qH��_{�~j}����T����d�w]�I�*�bW��$���BU�i6an#{W]C>$��e|�Ă���TҠp��Q~Z2��Y��n3�ؘM�u=���%H�� ��('u��/�K���٢f����M<�>��4���?B O��7�A^�]��R=��u�kx���f@�
5E��/\��M�H3�u_ĂI�T	$S����s�Z��Omn݂�U�I�����՞�� �}�~�; ��wh�2I  v����]ep�|�E� }}q�~�q�"���1�;�=�/#����vP��t��L4D�~����)���쟉>��'�M=λ#�ka�o{v��$��G�#I�a$�(9W���O݇�M��>s/ ����Z��
�u��R�盷珮�D|5�]PZi�N%FR�������� ��V/��j����GA�U� ����H� ��l�F�m��Ǐd�׾1OE�L�I=�]��ͭ����q1CF�s�l��[�u�#6�~��k=��߶ݏ]�}�V�NzD�{3.�� �{9���a�,���:.o�ُ՞�����~$�߫�~��<q�p�L���]�~>�]�`/�!b�"�!D��{��9սvP����Tѹ��	��V�e�,��Aۤ����O9V3X���5�s[F�y���w�����ۮwN�Ş�*�2ł	��b�d�\+�m
7 =U0A!V�ݞ�k�5 -ƒN1�:�~�&��ZS��I!W�d� �ϻ�C���}��cz���Y�4�IFĻ�r�_ޛ�V	 �9�7e����@|Z��� /wzJ ��j@�h7N%@�[��G�<=�U�V�u_Ă�;�����O�����nK�����
I�q���ω �gR���w+��w1p���ٹ% �����O�p�g8��.����_CO=]��הy�(���d�.�`��_J�.��݃q���:
��7��Y�\�Qç����)d��q��| �]10��◉�۷!�[��Sv�B���F��S�͞��لlZ��4������+{p^0UHF�Ǵ�C=��q]�<����s��s�#�ôp�t�(�u�m�z��:Νw[���8�D��q��Vݕ�#����l��&��p���2��
6��m�@s���n����;��usV�8�n���.�y놴�U�U<�o-v:��n���;�M�g�n�͘�̷�g�v���$���gGX�C=�r7{���&�E�?�^�eX$��B��>~��y^%�F;N�����od�P��ou�!���� a@\�vs���^;s����̡���;�_ę���.Ǧ�C�n����e,iH.��W���|���d
������yQe��8���Iy��@/��tl!OK	$�t䡙큋�4�,K��ϗ����
%�M"����B/�;�^z�I�;�$yd����a�}(~���[�m���N����vX�I}](�O�����&%���
{|e|XWAω8ȹr�xa:۱WHݝ�`p����v�:�^�p��rn��_-z
M����^�I}Y+�A>޻��˥�ˣ�pW{v	!�l�e(W �)Ca�.���pR��i��;�za���^�+Q*���QY�Q���gA�c���ٙ�7��1[���&�\����0>n�wuܝk���B����"�������Ǿ����o��ߌO7v���|Ho��# K���a�nʔ���{;ޛ��H$ש�	����?n�KU��AM��c���Z�����x��:Z�G�A�ݶ,��޳��T�y��N�<�7"�E��( �b�Q�����޵�� �*�=�����'�U w�� }�U�ɍy���KC�
7�,��(C�61*�I.G3
�m;��Ttlu��������_��p���-� �$�����oP�����;�n��'��Ņ�-��mG!��]X	5�'��#��{ُ����c��	�go]�IS�"й���G�K�s�?Jx��b-���&hw�vI{�����嗽���3ʫz��X�{$��Sޕg�N��XQ��cD�dM3'wU�;��3�>ޤ`�
�������*j�/;��ᘫ2_ﾪ��{7��H����Vv��'�7�	�1�M	[�I/�}מ� �']@�ޕ+��U�D���bJ�����e��% ,&
)��;�J zo�Y�[;�Z�` ��꿉�wu��]Aԋ�T���{��|OFZH�0J�6u����ʶ�m���-ϓt0O�dB�jBa���Ǳ0�J6'�c�u�B�ޫ �Z�dԧ+$W9�ӲŒguٌ�O?��7
���}A�^��ߦ>s���	��;��$���� ���ů=�z��Y+�q�1���Cw���A&r���?w,�f��T�Q>������?L�]_3Y|�6cj8��r��i�!�ęy�B�����P$����78�Lbˢ�N
�'���K�h|��є�Ӽ�s��9�X��}0I�`��
�6�bW�DY5�(^+�;�����ss��>P���ojd�8.=�s�#J3w��Y���B���,�S�.����$�U� �c��ޯw�6���u��4;#�7n6������痧JL���K'm��tD�@`)9	y��ԗ@ap����s$����t���\�Q'��Sq��vA/ʲ��I쁆���b���dϺ�'���U=C�KΖhHou��nm�U˛�{x��g�x��4�S��cp�2���%�wU�O��m���~�~��I~��_���W���6A	�ĕnw���FK�3-7�*n������\�˿�^��&cB>,TIn�����3l��q�<�7/彽@����S״3��W��$�b�����n�gs�����n9�@��o�����ۇ8^�۱��yglwG�'��X��&��_�@����ü؝���<>�n�<5��&�q:�ȶ{���-�j�ߴ����fk����Qch��X��ñg l��n;�����J)+�;��샳;3$��g����u��*�]m[󙹙�FD��݀]~�we��o}������O�#)�s;�\f�)��B�_e�Z�|�٬�c�wd&u�Fj�[>��雷x/�y�)K�01��w:zz<͵gs�=Y����t��\�>�5X�:�?�sM�l����G��~���0 s��[1=�;*��)�ܪf�x��_Fs��G�g{�>ו�V��g��f��
Y$�jOOz\~��em<��9�;.��aj�x��[;y�+h�y�.���T�M}��+1�f��Σ��*V*[��n�S\��.�>�38���V�<�&2cͨ�!
�u���ۗg�K�I���9ך��&g��V__z[ł�ӫa}�ƨ��Ud�/��U��`�Vi���]����XA1�m�G��d�$�oٷ����`{�1X��k�۱��|��H��j�T0Bp�ީKyVGc�ō��;�Vo��oY)�c��n�l,����,z��0����E��`���%��c��;�����X�l����7�E	}�i���A�k)���A�3�+�+��b/M��F����)s,��:ڤܙ�j� s�nqlz��^�a����Z �+םR�տB$�1��
ch�;7>�٣7wD,�
�� �Ȫ(�"�j6�V�[D"����U`�X��EU"���PZ��PX1���,�[
�E�����U��
)0«��E�(��dF,�DF(QQUQAdb�A���F+#�-EJ�DX$T[kP��X��U`��DFEEEDTb("1�-���V,UQ�X�����ZŘh��X�UQL2Yl�(��@F�YBհTUE+JT#-*B���(�F��UHV��cP�*�)(��B���X����DV(,�V�EP�x;�8�}���7��`�q�'��>��Lv��sf'����[���1�ܷ�G������hz�u�U¼7s���nz���<���xd�a�v��//`�i������e����V�ɫ����v�^���+�S��[�퐸���=�ܻG=�ٶ��-�9�ɮ6;9W��^�]�p�睰9��#�n�W;.�n�q�U��z̈́�-(�=�z�m۞Aq�4�nd��u��۶��r���[��N<�b�	�R��mf�vgi����ɩ���͸ѻ+�5ڹy�h���(�;e�_=w[\���1zx��ݶ.IuŇ\bHgY��]�6�N�&q����خ�A!�h�7k=7�k�^�S�b��לG]uuH�#���&�u�p�v�[���U���/`��uw<l�������=�/r2Y���kY�'��&��Li����	����6�vӏ͓���:�������3��"�۞s�n��Mj��8�|��W�m=���']�T��	� �c�e�f���ۯ6큓�gO��O۳�q��۰�`�hTjb���3u�ۅc�m�n�z�6|�Lp��m��lƖ-�]�ǎ.��up7li��}��r{NƗ����1d�<i���gq�և�@��Gr��6�n��T�E�ù�Ɗ�!ݎ|���SqΞ������gƳ��my{mƞL�lpn���(���]u�{=�l���#Y����\vܹ��]��W#{�:�8��h�Cۼ���� ݚ,�,��v!�gb�װ���]��/@[�]۞����<�	��L�cn�nG-����lcn�d�L�=+��y� �7�(7k��繵���z1�wM�i���zy�[�T�y��;Vۜ�#�vk��X�nw��o&��O�r�ڰ�hz�d�6[�R��]���q�um����֝��\�cj��^���'�Ot`�s^G
�"�[S)نq��v{��fا�;nBdݶۃ�S���p�;�;��k\gn������b�绽���������So=�ƛ��|*�z���gh�<s��W���u�֕��/\8S�<mNs��8�f�g����ϗRf�'09⧍�nx��w�h��K��hv���;׋�9�B�8 �::6�-�ٍ�z��]c�G�s�+�D�o������S�����s8^`�h���k�Jޑ�q�v��&�E����#f���Z����x�F�8�6s���P�n�n�Z���P�;��~f ���������H.o���^���F�0y�x^�w���п�m%�M��p������~!eE6V*.�]ƀ+�����.�*�׷��;�E�)��*6%�7�Y`Y#�7�� �>`��	ކ���H%��]�I�z��Cdj�\-�T1�UU�8���s��ܪ$|n�}b�$���뿉#o��ˠ1SY�x�Y�μ�(X� �i�L6$�y�>$��^zQ5<f�0�^�F>޻ �Oݝ]b����J ��l��'���-�u��KՎ��ݙ�HQ.#�^Y��Jť��/�s��ǡfَD�DS�β	>ޮ���7��\��u�2c	���'�s��쟟��jE�]4�hIC�5Ռ��>�1�<�O�XcW�ë7l��ܣpS��O�N��۱��hԻ��6y��p����tE�r������9u��]�7&fm���������@������>���;�@v=yv�r��7a'ZI�#���5]��?�\�H$�������~�� �ސ����w@}Y�f�C�KJ��7={�L;�&@�z�H$�m
�O�����+��J����]�$Xg��l�č�U{,
j{������Ba�&��P̽u��i�m���	�K�*ϥ�������y��
�#[l��l�(;6ϲ�G�vSc�Zs�ۮ(���i�$��C}�{ח`��}Y(�>�#�_�:OW�l9Fz�CAu�Ct:m$�D}�w]�,�zOx�U`��֐N^\�T�۲L+�p=kZ�y��� �lM0Z(v�%~"�{,Y��Y��3�MK��{�R[5���8Y�"d�3$�y���nt��=コ�nٹ=	�z̺���k[ٸN�!�5��^�0o�<C�8'z���W�������̝߈?�� ���m��-tK`�L�o�=�d��u�q�?}@|�}noI� }�}�.@��p=��A��J �7E*I��RQ�.�9�$=ޫ,W��"��݃�o.����y��gw���*�A���BȌ���sL�8�Ҷ2������{���@�v�m�A���x�1$B.��QԾ� {�zO��}���3���P����MKΰF��3ap�k.o�Ń<q����W�s	�@�ۗ��S�J#2��ؐr��Ku�6��� �Dh�ޱd�ݵ�d�%ϟ{G���0P'�O;*����]�Z}d�jH��ڻ=��p/u!�p�l5��vݒI���~$�_N�CM�ꦃ��$�������MW��3�S1�:���q����+�i�vSJ]�Z�,�ydegL:�X��y*q-�3��}���~�ٷ`��V���)8ۉ�~���@��t2ˮo�o��3�n>��(�޿IB��=s��nM�[`�Wb~g�ai$$�$����\;vl9���4U[�����(�PRH(����
p$�bo|}����mu}`��U�
�U�ܟu�\H$om��ā>|f�c`�$�E_�t���*j�gf�]V�#s�����}(A����U���J�C��P~E�Qp�.���łA꼔I'0���e
f����	$f���$���@��]�И�I3!��gnx�c���{��`�A���
 �E=λ=~��^WU�Z|<9�$QF$iU�{s% ���Jg�?Y>{`9&J�9��
�}r�W����ݓ�/v�|F�_��Mg�ٰe����ˋ�ۏŜX�N���6Z:�ˤ�����;��E��U*���S�ީ��ߞը������d�.�[&�-�{UfOgݬ9�;�H����x�wk�6u��Gn�m���{�̽�*�ݫ��{4�	�/Q�'�u���c�
��*��{l�yrt����o9%: w�:9N��w��g��=�3���v�؍ܩ��u�q���\�4���=���+&��w<�g$>ֻo[���>�lGp�pb�W�۫���]#pA�N:�`4�M�㤡cs��M�[�8xy��+k����:�El�A{{za����q4�l��o{.���Q{�Vo��o���+|�=����� ��
��K�T
tIe ���g��O����A'��(�O��Y�79�}�����xuP12CD"�U���?N�Y��KS<��J��$:}@ ~4��A}� v����bVw����������`|'r���-n�P�m�OUy�..젶���WN�=OE�Im8�����@=�}W�Ỽ� �������{d���v����k[P?X�3���E�BlY��3�nҙ�Y\kulE�!�$	h�{N�F�2���c�L{�Ynm�Y������2���vE���[�.2�l���}X	)��zѸL�g>�g!�Aգw))@u�&'7b{;����!!C��K�X�፻{�b�u��u��ͩO2�3��9�O>���Q�@5�߮�=���$�i6ȫ�w�~��At��N�,�䡙�%@ ���@|:�H�����vnE�}�5���}��ң�Ύ�0�Cb�ey�j��ηĂ�3%A@U@P�/8�ڝ�~����@Oٗd���P~E�SQ1.��P�A����\��!��{�8���$�������}��a����f�K�
e)d�������&��p�a�%�/\sl=-��Z݋��۰C��lQ1)�0{������I3����dE�F���e:����Cz���´�zKr8�A�R�K;R'+e��7�3fe��� �=��D�j�Ϥ�h�9�e�"���^��s@LEQT�_{Ͱ� ~���5BWH�2n��g���'!8�; M�x�b-��z>�u��	��9*��|Ƣ��y��/����5֧	�����?�\����bW��V����v}Y=s=��H�����E$�W�}v�g���
&)������*�w�̩�*��2 �+�i�[ݘ��%Z��Β�A[�F���C��h�2堷��� .�����7��<�qF�s�d�jH]ݙ�5���V���X�"!�pH���Q��Rnz��n^��n	�n�u�uJuۃ��9(������?r�U�!:~�` >��r$�u�٘���53���ٮ~�!�f���"m�Ѷ %(�"�=����(oVc�ꪜ�&k����� ���DD5u�٘���$Z�r��i
��.H�Q3���O��@>	��y�@�����2���"!�'m� �7�٘�����4�)8����+�,s�u�1'e m��ND�@M�vf  �o��
���P_���z$k�M��8{��[�)�,��WR�;|"e|����w�9W����M�����VЌϯ����r@#����s����*�*f�Ǘ��� [��q~w�s��ֽ�@+{\� Mﵼ �[��>�Z���x��!�颀/pn�I��Gϖ��It����D��v�ѝj�y|���G=�@��
<r~�iȂ"ow�`|�(��;�tD�+�=�V�ˣ���^��A$ҽ��ω4�Uz5��4�*O�>�I	�{��-c lZ���t��yݙ� >���� N?tʁ���I)�s���S#`H0IQ�C}��XDD.��l H3�:w_?I���y �of`DB�o[Lk�"5I#q(�e�����e��P��±A�����x�]������A�ʦ"^����ff|�^ʃ�$�Il��R�{sd��I{��F�xò ���3 ����o�@�nO7'�Wm����b�@�S�D:�;3PQٚ8	�v����Q��5��M���7Hѫ�.��6^z��ܣ�������pZ]��Z'a- �9i�n>�B����' ��G�e�e��>AE	]���=��pl䋇L+��'�ݵ��j���=f��U�8���u������r��+�����_	#�yâ�c��1�5�<+�ү��cq�k�^8��lq��݉w��]���.f��3��m��:�ٲ�.;j�;��7#0�3�q�ヌ�ӝv�]���4P�༫��J�s��u���T׳��C�����B�����t�q�u�!�g1����֎i��]������m�/�tܻ�� ,��l A[��D-jv��mK/{<��+u���_m�$��(���-�y� d�ѓg�"g=��D ���D�^��D�O�*Yխ
�Г�
��4�3D��	�sl+��� H#�Le���Щ�V������($�Sm��T�>�2I*8�b����O��Y��
k��Ȁ~u� �����܌O5�~�����>@!k�]�j�D�7l�Z�s���[A$���l����&1,���5� �u�h�[�Ui#3U<������,#(<;j-<�g�/��=c�6��p�����o-��k-��ǉ\n��I���˻H$�J���� ^�6���=�~�~��$/n��Lؽ%|�������	��pÞ���O���kc��~�#��Zj��.����Q7�}B<9���)Ó��frn�`��3�;i��YQq�m-q*2��>���!y=������*��_� 	�}c� /{� ��z_�f3&�詽����MW��Y�	f�J�Ϭ[A%�_��� 
����or.��{�9궊I
��I��Ñ6b.&�uai���s��.�u�֜�E�u��6+yڼ�D��q�#;�[�������$�T�,��8�/�WJ4��mFt{a����b��'rr� ^{n�'�G޹UgV�+����t�Z�ѷN�&��TA�j�Ѱ�z���Z��ݫz�x�L�<3�f8�M��j�.�yv��$��l ҷ�?�,���z��w���{v$��۷d����0��(dRSϐ�;Ͳ"_�B�R5N}=�D��~�m�[�������ޜ8�̏T����ɢk⦠L�X�3��I� �ϭ�@$�Y1��۞�r�~���7 �mm2��K4�������8
��7��S�:/u�5sx��]�緈u��c���\�/�ѽlq���˞�{۳oN�7Hk����M��M����2e�d[�~|��Nz�H�o����%�?<��|ؕ��N9:��9_*D���+꽛����U��2B�)�FV�U�B���ŷévq}�3c���-/*ue��ְ-�-�b��쾛7^����������9W�_ч��x�&y��u�L�Ոu��>����`�e�oq��G��ʘo�ڒܕ����6��B��*���vr�*���tT]b�97�i3S�� ���Κ�Wj��#�-U���:�b�uv�n�[�GE�U��ݗ|��.H�����4���>7>�����e��_;��,y��!�l���G�{�Xu�</k�u�kk�����L�4\���*륒���swjD ���i6'U�ވ�
�3N�%nw٣39:vM��V�;��w�\^��'v��wv9n�ĭ�m�`7��k�&%��7����s���H{��!��Ijm�xuً�t�������Y~"��W�~n6�{tX�oWea��K��<LR�v%:��kϲi�?p�Ϋ
��F�/j~{�4�|�^���37�a�k���Cm���x^�Q\�Z;�� �U�%�Э�ݔ$��/�u�so
��Ǚ�viœ9r��т�6��F-��ٖx`�KV]�v�]���1弩g|E ɤ��	$"���E�"�`��*E�,Z�V�d��Em*+
[`Ơ�"�%J0R,R-J"�E�Ab�ibZTZ���,Q�F�Ъ���X�`�

.)���X��B"��D�mEk%b�*V��-T*�h�R[ImұB��Q�Yڢ���AP`�\Z�H����Q�F�\[���Q҈1�TY)EkZ����Qb5��l�EX¥��jE�`�YB�m���[mdX��UqJ��L��2�V�ZU+[J��E�+���`�B�RڬHEZQK
��DTaZ�X��mDb��PG�b��)l*�LR�����}�n���{����u�lj�В���S���=�?E]�'=�7� U��� �� !�O:�j��7.7�Dn��_ʟe &�iHk�=$&�{'�9�<�=WWW��Ϥ���y�/ry��}����j3�T��S�4��&�5]��Ɖ��\�r8VB��u�[m��H)AL�>[�6I('�_)y�v����� �ܮcH!�o������rID�MgN�%J��i�[)&�JBwڶ}� ��2�I���@� /ry� A��'/ޟ���g�{m$wp0��F!�\#�=TI��g�X��H��W�ײ��o�� .��� �"�'��V��n��I��O�z��vP9���*�RH�wp� >���DD;���d���?����5� IG޺�m
o)3f��3h��G���e��r��o{z�����ՙ�z��E�Qe�B~�\.��U��OX��������c#����z<�Q���H �<�T@���m�[=�.Fk���p(�Ǝ����l;R��1��o9�W��d�t������G�_�.� iG$��	�˶ �n��J�����VVfd��3d_��֦8��3
LW�m�������~"��.��a� +��9h >��m�;�<��f�^�d�����y�a�ZE+�N��\���9�m�@ ����̩=wq���9� s�m�O� �h�0۷>5~ݓՓc]l�e�fJ�� <���`|��|�}����ll`O�䌼�қ6�6۱>>��)�	ݾ��'c��{u��\� ��m� ݾm�1[s����ӿׄd�Χֺi�Xf���p��m����k����nz����R�a���tBq���7�.G�콥H�:}I��@�>9�n*�pa��]���!`�����Pqq���7P���Zy�
�i6f�OG&�n�ƹ��i�\yU�4�y������NA�<���l�j6����d�����1�n-m�L��q;�A��V!PN9�]�΍s\�spn�V����������E�,F5n�'U'Y�����gvnq�M6":��{g�Y��v�Js�Źz�y�txwb��Zv�f��lM0܄玐p���0��{����.D<����F����Yoj����Tv��2 5ӺITJ��[�*�5Um	��p�s���c��� ׻v� �;��!�&W��df�Xw�j�6%A�Y�6IFg�]�}�F��9�m& wL�lْϳ�{>� �_��l ��ͦ
�2׈��&E�R���ݬ�Yl�,�@�2�BP ���lZ>w뺗�#GD���ZHT뻴�5�AX�i��Ir����� +���HM�6zb�b�	��l ��޷�� 
��iQ���g:�������2�0BJ�H�
8n\nlq�]g�j��qDi��1�����	������׶�@UUV�#;<��&=�u�]���/�5ٔDF�W�U�/�A3��,�8P��� Q`ұ*��s�2L�'/u̘��~���X��j_t_%�Y�K��y�k6�=��m5&�̌c�:���b���ǥ��ޞ�Ow��Q��ʼ�������退Eh�� AW���2��nFQ�����D�SUM�/��"��u ��zc}9��{�+��H��v����}L�2f�$�!v��(�o2�nP�s�` ���C����tY���q���d�7�m�(��e�V�Y�	A*�ڢ�����f�}/ް������������5�+a��֛ly��i�a]r��=����mE6�>Ԍ���s�]��������-r	�4�N?Uf�'ğ�c'O��
����w;��偝�����%��%�O�c��L4��ns۱�ȍ�e��*G��d@U��� �����Y�D�/A��4�-����$��h-��ЀA~��_w�����7���/?gn}vU��0A�7d������ۨFnf���k@��]���9���g^���>:�8��� W�T@�sl'���3�-6�|`��X�fQ��/K�3���l�Z|M��w>$�C{���ro+��P��Ć�ػn���ہ�A�k�[���`��&;�mX�λ��#}�Ŀ�Լr�y�n!�L{y�k�^�'7u�Q���B���$ˡMK�7\�xgtF�kEC֭��uR�se�@/'������i�Pi�K��w- ����H{z��<Q53��+��Q _n�Ѯ�P�[N(��ˣ����I-c��	�S�rSiЀ���������Y�F[�7}����4��;V�:$�ۂ�� oz�� n����.�g�"��l"�1��Շ�Io���ۅ�f�Uk��k��g�(f�"u�[d@�I�ΘD��|���9֪�6x`$�-����ߖ�1�)Ʀn�;ۀ�r
�\hJm��.�h��F���o;e��~x!Y|G��X�	J��A��r/��D�k�擩�~�O��g��;���6�DD��[V@�+G��1��=
��9Z���kY�b62�{sr\�k8� 헩����F&`dA��ͯ��3>C��A1�ۨa%[/��oa����iM�I>$�$��щ~ST�"]%-��Ɲ�g�"}����W^�Ȁ����	 V�����V���Ԥ���	5L��$�S(�8��2��A�)�j�@��Ny���7�
&s:�R$����}�Ӊ�c��$v4�{g���<}����m|I'��lJ 
�~r����ٵ���/U���9��>�KH^��D��J�-��: A}��0�����KH#x� E`��D }}�ٙ�)��z˗�ݴ�_N9�}�y'&�Ys���]�":�N�[BN��ԳC:r��>�r�ݾ��:�{�M�l���|o�,5P���	�w'��;��@A�v�:uψ�wl�:��܂���֍u��ݧ����5�v��S���������מӞ�$`�8����J��Ni=N����c�<'�cq4���d�l:��S,����jD��lv�G��w0v؎'c�>ͷk��c����u�:/[({n����A��u���մv��N���i��a �kq�5�
\�-�dn���Q1��z�۵�JwQ���}�F�b��Y�/+�ԒD�W�.� 
��٘�7�eܭ���z/��C@��j������T(M�ٝ��N`�hl!ۣ�b�����D�^�� ��}�̢M�d��=}��^?t~�L����x��B���n�%������ ��TMP��2�DFmvTG ���� @+�wf`Q�O4B�І9r���e��������$���n� �n�dDF"c{{(�+����h��I*���h�˦tKM�9�ۙ��&7�ڲgut͛�d��z�!7��H  �z[�7�U2�# �i�</n�'�i7�u�.��뗝;[k�C�:�c���@�z�w��D��J�G��i���H0�#�H�����j��m��yͫ @_��3 �~j�J�"UDUSfM�O���uW�d�s�e��i%��.�����}��+�ȏk�u}�K�bz�!���<���c�[77���3�ӛ��C�<o��"_g�π��wf`c����C�jΐ�O9wIS"񣁐~0HI7aN�w��	�s��2Q��Q�f_��H����I$��H�~8�Ӥ�h��R�;�C���I��D���` �Rw7L �����}�U���>O�3Y�OIS52*��tь�7�� �7^!����O��X]ݙ�|<s��i�/G��(�۬�i�=Aw)L�WǙ��&hR���#�d����n{s�.�"I�!�R�n",ȍ�����KM������	x�\d�H�zƂ�T�	�+j��>���f���'̕�=-&( w���G��"�ޒ�j|]�>����9ܰ 
��]�RT�$��纜�{�%����䀠i�Ym�Fx͒� �~�eDJIo	�9R5T��aЯ?u���$mL�d����$�t�<�)�zA>0�����\2�B��}���y��y{=D��g�D�5��$z筤ҦE�%��~0HI7jW{�g�����z"�AT=���|�u��`^��a�ug�yU������WEf�Tҩ��
�%��O���_os�3r�r��U��S���z筩 H/�ސy�y�Z�Y �h�T���d��샣/�mZ�����q�rη����Q�����?��MD�������6� �/� ���vf)D�}HѴe��b }om��2���̀�ݻ�$�<��q[.�߸η@+�^cA+�wf`t��":^���g����]��*�h�7��nO�A~�s� u_�L_<��n�V�C@#[�7$ '����>��VΒ�A�*������?WM���.�� *�]����� D�N>Oc��qKD�[����9�ᙔ0ϊ�Mw��m��ڂP8n�N���'�W����r�E� �)ReUebl�S�����H9��K �`�nԫ����($��ji�ș���)�-��o����3I'��|��Nj�N�e��*��)0��3���B�s�-h2�!�2�i��n���3#Q��rY�2���	^�sŀ�Ouc ~��/{Ϊ�⟾C��tA�	>����p���&����ryl����>�����~Ùр�o7� ��o� A�p�T�$�^�Ϣ���22���㎍���w1a|]9n@ו��SsW> �ovf@���m)DF�Lh@�)�J�&C�/����n�Y儚�vgc�� ��u��`#p�{M\e^%p��OQԐ�o{��H?����_A"����mP ��3�ҩ���_ڲ���o��|�#��m}DD����|Vy�r7g/�ib
�7��7��n��#��LI���-������N�{Hsٝ����I��C�D8 ��;+���n<Wj��Xp(v�S�f�`�'踵���󓢹���e(5֗������(K��V���>��=w��f��Y�蹜��s�MD���aP����� �s�y��?�랜����(��y�_�1�dPJ�>KOt}
���u��]��.�w�/����l�/���Vr��&
�&�HƟ|�w7����WAt�h#�ƞsܢS\�R���Y�5���Y#j���qɈ��OY����N/Q���~j[����}�dS��R�c�M��V۱z�)�[Mx.���G9l�1�xkUa�����{������Z��&Xj�p�߯��Gc6�p�|qQ���0\�j]���2wt7�]w��ǽ��_n��"GF����+���㌧�{���.l}�(7�[9��l�����`�}±fmub���d o��򹖹���,*�=��fr�~)�<xcx���#rN�!=R�8�5�w1J'Xӷ��R�N�<��
WL�:5�<ـN��>;4/3�}�������x�F\��uGs�:���A�����uEml����{���(���Yݚ��[K�A�1��D�7�(RniZ����)�C���B���ٕ�	��=�Ƕ��@��w�̵J�a���.[��n�c����w-�OV���;�����d'pӃ�O?�;w�]�r�X�����[���ٝ�Y{�#왩�YV{�?f*(�����Z�����EYbZYiJՊ֛���*TQAATPQDTR"(*�iVVDe\\p-������Te\7j%b�J��$mFkU�m�h��1��J4�ī�`���L[U���PiJ��)+U��mF*�Jƣj�DZ�T,V[H�J�
VJ(ؔJ1�UV��T�J�cZ%��"
�iJ�ETX"T�J5��TDPJ�cm��Um���������XQ�AA�m�V��DQJŪ0�V�
�QVҒ�R�AV,0j6(���E��i)iE��E�B�-b��TA+U�TJ��k)E��#A����+*���*[J��KQ,�
V�-�Z�
²��UA�7�8�K�&��p�wnnm�\�W���j3�d�ƺݞ���6����z�뗓�hs��8�v�]Y�A�&3tݶ���w��W�Z��n�k�\t�6�{v��g���>A�/^�����\U�^{s5��;��a97\p'=�r�[[�۫W��wgj�u7����GHQۀ#����pvr�b�h,�����Mk1�5n76�iyk
9�7.:��j���.�k�f�X��B��]Vv�<=�9���QێuW�:9NM�{s�y���H���g��=�9�xݢv^�ڜ�6$�skۗ��`����52����n]z���M��u�#�&�����͞,�.��1�k^��Q�����#v��kl���ren�����a˂�U���s��v�����Mu�&:_<籞ھ_/��=���<�v�m������z��>vî�a�pC���7	�:7dNznʚ�(�M�{� Yg�6���K��-��8�{��[����Nu�1�1�nܩ�>,�ȉ����Fm����y�uݹ�\�]��)��K�.3��7��^����e
x|eն;�{�]���0�ma��0F�p��\ux�Y�X:��u�\�.wm���ã�qFI,]�T��%h�z޻^2���t;9�����WO����R�-;���'��c#���N:�d�s�;��L�lc�t)��4n���k�F��-�]7hswM��^A뎠$��ki7O/�:��n;m��P�\uե�˅!����q�GO	�=Y�6��m����Ύp�[y|q�����ur"�KpK� ��`ݻ,=X#��g9]���r��,
; sр��$=v��J�&��W��H�c��U�l�{A�6��7ls��Ð�g.��R��-����k��o<�nm��n�V�h+o0C\�_g�����sOX�SŹjn9����b0�۱�|���>p��pq�ݰ���`-;��C�{���m7c����[�s��gR�y�k`���L��k	��Ǉq��y�����\����0S�ཷ!a�;;��ӎ{u�2�.�!Ϗ
��9���W,��Ǥ�dN�	|Lħ�*��%ۅN6��cc$���ۋw/n�ص����5t1���:ˎ[tu��v�'+`<�s�x�&Q0��j�oPWg\�u�iB�=�l���k�j�]z\O�E�v]�a��r��5�u���BF��gpWgi�Kع�.�[^�kg��:�����;���Y��n�J!�����` �G^[�@ ���4{��5����a#G�.}d߃�P-�!�ZI)(�qݑ�%�#b�w7�@i[��@ �������]"��������Iw�xRI8R�.XW�mX �0|�u|�ez`��}{�:�0 �{􌗽N�%�Bi�������콻�*�﨓�6.����/�	ﻳ'//w:�Y�r�ʘ�3�$bF �� �e2�\4���@ ~�s��{���y=��!� .�|� ;�� �wv{�%��I���P/8�{/ɑ�)>���[��9Ü4��v��s�&:w;�J�[m�^��_ػ�zT�>�TUC��mP|c�N��@����Oh�~�'�ѯ��mQ��b�Vw��)B�*�E���>��fv��}���E�nF�iҜ[���N�0�P�Խ���v���3�֪��yy���(�/��D�\y^; ��tQ���ߗu3��yM� w�'��O-2K�X����%2^�Q)�[H��RQ;�vTd�����ay�6{f���]^� _��� 
�{�3�9����jTUS���9�ͳK�V������"�7{3 	��}�ޠEWVlGUh�=�}L��N�!�Bi������K�x�\ǂ������Gz<�P����� <w��7�de9߿����^>��A���ƺ��::�����uk��;���6'8z�z����}��)����p[7�АD^{��X �x�\�ܶ�7˸�;�� >�ovf?R�\�*�M�ĆgI��K�s��2t��"�ZU�Q �ݙ� >&7�ݐ�(���ƕ,�f�2/�� �t���dD���m�D��q�@�<�{2��T���-T�ֱ�B��.JΓ2�
�c�:G��q��K�%y�c�3��.�OUɧ9�7��g��a�ȊuM��� /7�3>�1���/���Ja��-������=X�M������_kŀ� R{|�Z>f^�V��2� ;��N$��`�@�� ���-�o� ��7\�gE�w�� �o�� �&;���@�+G��7qe珶���$��(��"������<vŬ/�N;C�8���Ą�@�$��v�С)��M4�|s�ݙ�I��;�s� O�e��y�Uܹ����Ā@$O뿢������6J�ϩ_�� N��ky�����9` Z��+�C�k3�]u�+/oBH!3F,BdR5K���I)��Ŵ@�=;\4\�ph�~��D�M�� B�/B'քCZJ��	t���g����ݜ���a�`@W�s@|כݙ{���s����굪�F�C�[Ὥ-?U��ژ��eI�e�]�k\��{�;�s0�|���gӗ/[�g�����J�� ��E�Ͷ%^�Y�e�-����l�� ����a��2	��{i�Θ �|�R@�W�ݙ�7;�5:�yS�
���73N��U�x�-��P'meծ�қ^-E�Dϛ�4��$[�!"r������ο�� ��sx���}��&����ly�Y �s��^�M
���E�ڂQ�{� �f���+�@�tϢ����k���>��٘�A~��B��W���ٯ�UI"��T�����9D_���� ��^��� A�=dC�}���@)�������*7�o�A���� M���Ȃ W���� �&7���'=��� �k˶���
[`EPL7�V��0&;r�VIQ��ǭyy�FO]60_��3��c{V[]�w���wd�Rr�+���k-��v݋��u;f�gu��WZ���ueI�/�K�c�����X�֩Z�9ּk�lm_�~j8QEM�+2m�ݍՀ��WZ\�c�v���Hs;l�{gGn���)�6�Fx�S��&�sթ�x[�
>�\p����ts��y��-v���p���j.�:ӷ�0�$�����N��i�g��,vtV�������]s�z��V�%F㧆����=\�a���4&�9۞��9�wnn7m��<a� ����f�ΞՃF�������g�y�#s��n�V8u�tQK�[��bD��n� _4uxy"�i�[I.f,�$�}�sń@�Roc���u��eD�K�H	&�=���$�1�m$BLM��=2�����;1O�~�NY� 緳1 D��6�� �^~����gM��Az�K0�ѵ��>�̻:��&w�P����Z��^���i� ���1  D��6��ЂCd"��T�?��Olf�٬�l�o�;��`| Twe�@ V�瞳Cr�2/���g�%���f��T�0�p�������e��I)]>'%��^��*�� 3/33��}�Y��W�#z窤q\�X���󣍧�`j9��ۭ�Q�J��,<��Y���1gm�ND!~ń���#�����`|
�ܷ`_�����o�egs�s�0�D�;�r���J,�����N�,�Q�������I�%�(�J�pԥL�HhD������	����2u��{��~��OӜ��#C{~���^�4���<nj6�"��Ou��Wv;h�D�}v�INu3*�ٚ��9#m�TM\��<�� �'���*��T��{�A|*��� ��ͩ=TѥM�- �n	���{鿷yVI=�h=�w�U{Z�~�o�ƴ{���Wp��O�[`�� �� �(( y��I����7*I=Y�_�����ڐ�m� ���nH�>���f�\�o<m���1 �����*�>���pu�<׵]0�'�L%!@���2���F*0В!��p��	 ��yv�K���� ��J��>�N{!{�oɐ! ���i
�����6jV��X	k���T\*�G�iK�}|� ��ü���0�X��2�z�s��l��Qe&�M���'}�,�	���>����=S��ϮM4�8ή�rމ�PC-Ӿ�F+wG��ƙ��d�!e�/�����r�=a��9�:�ѕ��L,�o�v{�Jn}�H���� V������0��rF�N�Q�W�חH�gJ����}s�9> ��wfb V��!�s���9aQ&��R'�_1( Z�����(�)���4�����[r�
��1� ���f > S{.�ƮZ��GE�>"0�e8$)��J�;[O\,\.�ݭ��xˆ��ӳɞ^O����~�����L�{��H��w_��I �˫	C����0�Z���%��.�+�۽�x�#T�,�BHj��[`�{xy��q�<�2ˣ> �nݴ� U��i����ײ}�ɭ�p��\���A��A�aT��Ce7ݙ�� ����a����AՄ��t��Ò �;{3 �V�����<8���#R6��K;���!�j���}��0 Q^�;hZ�^�w�����h����S��t��meZS�͗�m�uq��7Km��S�Z���w\���g����l�����4GUӏc��-����fb�=eQR���RT���?6� V9朡_q�3薦}֍ ���f|
���!��+\�iI�OW���켴ܢT�#�	�{l�)��
�@g��q��`v��Xnm�ٰ���}�Ĵ�(ɒI��wvo�<� U��`|�똇,�W��]9K�,��f`Wo�êЄ*Z@
�*I�g=�����];�gM�I?O{�m�h������l�x{P��{۩HG)�6X1��PQ�k-L�~n�1C�XV�ہ
�|�d ���t	�� �*�ER�����+��(3���/S �|�E��6�>�5�7�
��i���%i�f����F�i�i���n�+��hg�˟/L��w����f�u���ϲХƾ�T)wG�BJ�c��NK.�9VGgY��:^�sr�?u-��.�^u��x̰����v���?h�L�(��l&b�.lv{k��d^z[��kp�v�]�;	�v�`ݰ�n5q���X�E�5���^�{ �n�K�ݺӼx8�Ǉ�hӋm͎Og�(NU�vs���ս�Gn��ɹtU�n�]u��Q��r'lq���v��,�x6��r��c�t�a;nY�e���.����S��r��k���C�X�1rn:�n;5����;\�[==�Yc7n7��.�+Ȏ�Q�g��������Ȼ�������~�(���Ma�y������ ��fb�*A��������"=3d�Mm�DűE�m�*�w��0VT���,N�z^�L �[/����w�1 wS���.�_�&� �A��E@����$�ozg�Mh(��˯{����Ex}mQ���{�HFǲ)��0U�%������OuS� m�'B�^�{2#
���w0��PH�<o�� �"��.���}�H��ʣg&�t�&�Q��'q� /wy� ��˿�ww7���e��\K0Hѐ���7���踛����s�Y�/�-d�����;���llh�ԍ�U�,垧a"k�z� ���� n�n�/h�x�}֍��v")%]���>~�R(�r"�q�4/s�i��O�\�����DK�/<�6m^4���f��D�^��{��w9Ȏ�wR~���κSϝ�xb���Wvm\#t��f��8wm�zf�2��{�٘ U��� e{���v3�#h͹�'�Z�(�]0Z��n���԰�V��ဂ�g2�c��F=������@$Q��j���� ��	!��P �箯�LԟI�h�7g�� �:�V��<V�:�~�=�+�3{��IHFSz$���JDm����o�`��+���.���u�Sx�����DTozڲ ���e֧f�t��27"Q��m�!D��SX;Ylg�3�xK��1�lmv!�����;����;�!H�D8����"������ n_9h7J�d�o2���ߝ�wfbCە`RB��x�f&��(ڻ.՞�p��؛��N�z�"RHE��	h#X��|����#`���}� �3��� �M8a�}�Y$���J��Iߪ�n�h����7rW5Xt�Ö��l4��l��Fjv��֕C����t��F�����˃���.�r~����`6)ۼ�?DI�%6���!+�� }�k�`��V5o�^�������������в���h���^PqE��9<[���`��N�Ǔ�5�tyٷ�4�n�qQ`p-�-Σ����~w���+��-�nLO�Qp'�-�����K�c���:gy��~���q�rQ��=[B��NO77���:\��=���#[�JdE�XN�bD:���A���s��Y�l
0���4�̥}�ìu���g�HĪ!k,5X�^v��.�h��*�����:����:��'g�ȰzK�pz���������ݵ�9ݼf�� ��L��/K N���^�>sLj��b���jf ��3�CVVDLOʋM�M���so�U;��U�H����������%��˭�1���ZE��]=�<�f�9/�d��\ժ�_]Dv,��^A��v�p8s�LS8�x9-� 0��Jy����v�C:���v�+��UdO���-ȍJ�K;�hs���k�YVﵻ����/:����(�U��,x^��}s����[��K89&�s$v�}�q9Y�lK��4�cf���R���m������;b���5Y�������`4.�/=W�n��a4��@>��Ldd�yP��n��5��㶀W��'f�Ǳ\�y�@���ղ./v��X��ԛ��yZ����cEWD��)���#X��-)X��EE�j��)�mXƢ��Z�*�,�"���PR�X�R��FQ������(�ڥ�KKQ(ѴQ�
��FZ[aQ�ֵ��b��Qւ�ԭE�(��Z��mm*4F�EQ��m�dQE��lj5VV����T�R��b���kR�ڶ�(�D�Q��QUeK(�m��mZZ�VYi@�TFUJԪ**6ض�KlF"UaV�[h�E�J�Ѩ���j�)F�ch*j4B�-��$EEUAҶ*�#b ��B�Ш5�j���DI[m�TX֢��F�E����ж6Z�1J�KB�[�h6(�Z+j1E�6�J��Z�0���R�XV�T+**Ԩ�AhԢ��k�o�Tn�d#X�ڠ�ι��*0arY��w^�-���LvbD�>�\�r����=m�^C�����{3�|�=ͪ��A^��"�a(%&/Y�I���ޙ�Xx� �"-gNy�C��nH ����0�����fJ}}~g���������튬�^���η�"�-�Q)$2"�Q���zDT�
���` ���''� >O����r<�@��NQN�̈hcs�?\c�R����!�D���d vm{	��q��̜�RD<���� '��f�����At7WIH����iEUT�D��亮 	go<� �=���M��do���i� H��ͩ 	-��{�	.�ʒ�r"�q�VW?=�frj�쉗�^��� �wfb�����mT\#����㚵��ڱ��+7�9T�����@�'�
[���z�gض�練X]�9X2�����]�z��W��ē{���K)岂0B�%���}��H/�rڑ�f��aw19徖�Y{\������������L^��=��x��w�v|���g==s�s��g�Wb�CaX��q��G\u�M����(������~�[��r �3w�` ���,3W�����2�t BNg����s��D�E���-�J'�0��D_��;'59 /o��1 �H}Ӎ�$��፧�f)1W���h��lq[o��  �v\� N�Jˏ{�j�i� o��3� |v6�K��&Pe5M��2Q=ڳ4vR��g��Ȋ�<�` �q��ny�L�]ś=�c@�D�O3ـn\m�h�␪j���������@7<�s�F�]��~<h}~����g-� �k�)��[��M�H<�K|����o]��7���樸���1�eq�)�3�����^����D�|qu�6���� =�,�-K�{�{�Av|R #̲ce��X��on�y���F�m�s^ɡ�p�c�σ�ӂ��R����s��r���o[��6v�u䭵�g;ۛ�v7�.�q�of�pF�d�\v��vt��G'6B;v7i���.�\�n:�a/5������]�q�Ͳ��ۢ�[��Ǒ㛶฽��n�-�oln���v���S���Y����x���'>����d����1T�o95'+*�{i|h�b�ʼ�cg����aN;F���n��AB�&�t��{�$_%}��� J�����W�z~�w�[� ~��G����$S7y<Ӑ#b4�[޲��g�1��@ ~��0�H���@��Az�����6g�1�jbh%"6_S�D�	V�˹�wK�N�:�W?<H�t忤���R	���B(��H��ם�yGmC��y�v�>��X�@.����^Di/�ȍH�l�r
�,ꘙ��c�F��Y��v�A.��)�>m��fuc"�y���|������Rrz��ST�ZQh�T�t�F �7lZ�N�g�{T��*�nێ.k&N�_�����$G$��.�yw�H��Uy���ĒM>��`��[���hW�6&fb��?�-�[J�	�&����� 
�W:�z,�N:���{7v���]��](�7� ����t��k��B]�;t���iriwïyp]�:.m��dN}�fu���~�w� *��Ȉ�]�ّ�a��uty\�G�+��PhD�1ٴ��|ӑEf�<�FJA�yq{�
��;}���"�ͩ ��ٙ����E	D��:�_���;3�L��5� ۽�� >t���{`��l����]���9����QT��;3� >@�ӖԞ�g<�=�3Ŵ�լh"���f >�~�F������ڴWS0XVT{��:���g�b9�a�C���z�D����>b栍ct$���d1B�E������|{��}�A�Ӗ0�u�L���y��"Ğ����$�3-����SUT�=���* cٱ��_v��r|/k���FF�[��<�Si��W�5]J�KI�&��{}�|A ��e�a�DPӓ�����)�k.���+�_�;��w���乄 �]#�c/3<��O�xvW��G6�Cbq�7��ùl��|*]�n�̭���V㛧$�=��A|docvz���ځC������Փ��\ �xeEi$��sq�|���M  *�<���w���@���t$�V�䗡��a-F�qRl���v |{>i���Ȼ]�I�e���ݙ� 2=���A�_�]��߷�,���XeH�j5{sd���瓭L���!�I�B��[��gq��D�5A����>�"##w-��~�c�#vsp�Y��[�ٙ��27�K&�tsΘH2�n�fBw9d� E�Ms+!���{Q��~� ��!���O[RA�x~<���i�r��v�䞢Mzf[h�I�������$�% y<ӓ�7�0�����AW7��o�  �����5�*
�UR,�(�~����|}ń�	q�z��$��Vٟ���f_�3eװ���<��v�����-�<��t��c�Dg�7=�z(M���=WZ^�\\�r)~}Cws��>�u�߽�O|��z������"�����4�;c 6�y����}�q�@31�` ���Y��&_��\���?@�H� j��m�p��u��i�wL�s��ѓcC�a�:�;vq��"�a8��{.�/�_%+���� /_��"A~�$��3s؉����?K�^��2���a�@&�?�ǝ��E���[~��U���� ���3�@;���|J��hw�rɩ��($`�f��Y ��OV"PK]��!�vBI�R���P�_w���VzIA��%G%W��]=��ܭ܈`��最 s��� okQ��'�S�{0$�w<܆\�TE�TLMS������{���g^��Y�����>�:�4�{����@|8��Q��3گ�*�Y\1�S%�,z���Q�;����,9#�S�{ueVg6VV�wW��ƾ0q�=xrӢZ䙞��é8�m�,s���P�m�G��8zC{u�wd,D1r�v��&�x��Gm�y���:�3�����n�δ�fmn-f!�cW��ݶ�������g�7���LնY�Vc���n3Ջo8EW8�+�dы��a��c�q����s�=��-���苮7-�s%�diz�p�F�@C=�]{3;��t������U��:���ۜ���y�֌��v^���m۞������\`�wg/\l�g�Q�ߐ[��MH$�L�{H�}�� $ɛ��*��w���E�����D�c3s��|��D��!Q��P]���� <��)S���ND n����zt�S �2`Gog>���#jF3Q�� �aP�����0�=u�$)�} ����Ј7�ݙ� 5���O� {R(2�L�̄�j��SÄ��Y�>X  ���@ ��OX�k(�Kw� �=&�ksq[i�H'@��UQ��)�	/1zTY֊u�Āy��� ���!�
�O6�Y�RT}�<X���e�P�L����q�o�=����=��'�=6]m*gnT�n?>��:L��H&&�#�������mQ|{��N���u�y[w�8�C�s�d���Z�"b�*�S~������˹��~���ˋ,��2�B���+�K�G��.����p�U��f�B�]/��7}Y%��I�.�+	b�T_oV���/^\aX�s^�q�-s���d�jHta��8����os�$�8l�@dd'j�w]��_%7�,''��=��*3��{z#P��� �{�Љ#�A!�J�l*U;=�>f}ٖpD�=-	D��?>��` 3�ݙ�\`�k�k2k�@|���#7R��Њ��M3p��YfQ%|��n'�v��s�)���+�9vD�=۝�y*�;���B��J��{n.v��z[�\�n�נݣ�Lt���(kg�nY1y��ͦiRO��o�;��!>$����" ��vf ������:/��|����!�z� �I�V/�ݒ�=#��9]lW�bn��A[��h����{����۳f���u��e|��"D8�bKVUx�ŲI�����("�tPV��0��tpm�WD���W�x�v�X	���zM��K�و��ce0&u��sm��k�X��Z���+�y���fb�B&iq�bl��̋���g�������>��mM��l{r���7�/�5�����^:̼�~�b={��;��r��ER��*��los�03vڣ7kr=�4���
�����ޓ	$������10(!��E��k�v���
p��([����-���ێ7+p�dC��x�̍���%ڳ���_ ���� ^�y�A[�a3u���6kelE ���]�%��9#0���8��p�ϩ^}Ͻ��?H}�i���D@�{��1@����D�o_t��E�u�>eaA����RY:�������D@�ĭوV�/!��k�&"#wof`>7�a���+U'�Ih����xgO�Q�<�%�v_�M���)TH�>ɍJꏖ���T{v�n�:;�k���ȳ�x�_�����Q��[Z���HVM��esŸD3�.�Z�g>�X��9/��M���5�ϸ�&ge�O��6�9 "0�q�e�s��	m����z���w���X�}�� ��� Age�ߏO�q���3O�
��pD?���
\J9vϝ����<��^��Cg�*��ƶ�w�������R��"2+����O�� �{��ʎ�Y���\�^G{�}��� �Yr�7W��AZ�ؐ��6Tq�V�/Nu�}o��` ���!��3�n������۽~A�𪩊�FB2J6�k�D�}J��$�^!uef?e�;��Db@|n�q����><��)�6� �-"	����d'���X	W�m�  s3�, ���f��t�������O
&�j��!�O� �9�ޙ��fm�A
��X���[T@�v�y�A�$�ǏK��|7+ȃ�N	�~�l�2ˌ+j��݌�
�In�wdP���4�f�^��ƙ�>��m��9UsՋ����nUa��;�t�ovu����>_����f_V�HX�9�w��C-g}�EٳH�{.;�X��0�U���_E[7Km�[Ҹ����B;�5�\+4�������׌V=��r�@fm�X$�Qd��fD���پ~Y;�ak���E�{=��^'��-)�;��.�ɫ]JP�a�j.ӏ<M����ˁ�.5��6_w����%T�xx텾��m	g_�VݸG���M�q��-�p�$KZеR"��WƈZ=V��6�pl�hd{�+���<�����u:iQ��Y�Z��h�;���c�dS{	�p�w���I����Dl�m�l��ۃ�}N��g$�G��Q�����x:y*9Q�~�+�7�e�.3���VD�r�N����]��"��C��s��r�"�D3��UDGV�w�P�����t؃kD�Z!�����Y�e-���7�>�9��sxB�-
'�&w�^�Ӝ�mv]�x+��Q�]���,jP�������
���C0�T��Gp��&l�B�w�]�w#�����=����ɇ��颴���shΦ�L�E�`K��͡�������L�of9B�K�b�g�K]�tt�"@֬&��^&u��qn� $pJR�6�^�C���M�;��w�/��R��{�o�禌���7=�Le�{xL��(��0nI��������y�Z���D+UKh5(ԤTYXZڔ��kUKIUE�mV1QQ�Q-Z��*�[Q�Ֆ�,����Q*6���b��E�m�����kYR���Q`*(�ֲ�bJ4bT�Z1X���hV*�m*Z�UZ�A�,k��j�*PH��������[J�EV[%X�6�����kZEQ��h�J����"���b�����
���m*�,EJմE���elk*�V��Ŷ�(*�֪0Y*UIZ��
�Z�D�J�-j�Z�Vڣ
Զ[V��*�Z�Q�,U�%�)j4)YV�B��FEF6֍TFV�m��kQEU*���ږ�Qb*�cB���j���1+(�-R,VТ#iX��,���"��Q�"��'�qʀw��xWo���e��n�p�Eخy��jkv���s�GW[��4��xQ��n'��=�V�����tٓS�vu]HzK)c�8�\�m§N:��39�q�γ��d�WDt�۹z��r޴���M��Onx��k�]�Uĸ�O�^�$ra�6��0ru�n�l:݁.gq�s2��{��3�m��8N�)�jx�:�w;[-5�ԇF�1s��� ��7�[���@Wg���:��m�.�=p�6G�$���#���1Z6�m<ލeJ��G�1{&7��{B��x�wn[�mNJ|�lؚ�N;A�=��nZ��ޜ����k;G����Ww����c8^8���Om�c�3����۬�u���æ�.t"�v:8�mn�ݷ'3�6M�l>���vv�.���z�rj9��3��֐磊�5�6v���nَ�4O�%WH2e�OF�����;(�������KY�ք���xLls�{qs����4q�BL�o&����g��"{oB�p�Ah|����g��9CP�zS��V̶z�-�[ӣX��#�e.�9�����r�r���;\�����S<�2�Φ��go��͊�scw\l���ӽ�8����.\nSO,��8����tFvIy<F�}����۱�2ݧ[0:�R�A�|nP�ճ�6���\k\���:]V���I�Wun��K����ܙ�9㴽uѶ�q�m���p�v��[s˴ۍ��ݳ��rWY��F8�;a�9x��[�!/\��X����SӴ��vx.#×#Y���7�6��ی�/8�nP��C��Ts��7&8䵯m�:QǗ�ip����2]��q&v�H�l�u�h9hz�N����شu�B�v�juF�gn�ۘ��N]�����@v�{n��om���n����ͤ���kt!�ipJX�X�:��g�h4腳��v�:�L�Ll=��Db��.P%]��sG��S��^7��\&�c����ƞ�&se:�g��2m-��ӫx�ظ�wnx/6�n�V�x�ѷ fX�b�����M]�(���%�n*���Nx{^ˀ��ge���l�n.[g�ė5��wrA��D����v�\f���4��Cu�Or'�n��ñ�NmV;y���`7Q�h����2fj�:�,�\��sϱ�l�g5��k\f{<�y�8��{8���䶮ݞ�h��r�h��v�c�r8��۞{{��u��kj��99��p�i8�U��ٰA-�=r�;}������:�+�e��d h�9�	��ă�7A*��^��ϰ��L����Ž�ݵ@�s�������@����5ǟ���=�PRW�r��"�QU��e�@{�� 1K#��[���c���h�E���A�������喘l��4�i�(��u���"�DAX_7@ f��dF oƷTzj�d�-�?��!)��M �.��Bm�:�ێ1 ǲ��>��{��ެ���gM���o7�Ǳ�+�}S�qgV�K^댘BD�D�C�澍S��wGnq�bgqS����)
Q�X��$l�o�oEBUEVg��#�f��ϰ� Zw��3ި�<̒2 ���eTb��SL
IHMM&�q�Ρ�+,�4��h'�<�Z��ܺ5�5m`�n-�+_o<YM��.�[�V�n]9�Ҧ�s������C0qLQ�=��y�Ղ6+k�w�_'Bnw7� ���t �4��1����S	@n�Tf!��睘���7-� {8q��Ԑ��N����gvf  �������ff���qѸ糁cl��w<�����x�syׁ��˔ż	'���fg�L�V5M��.Q3E\4tncv �;�(����r�Q&zM� ��}� /NzJd���M��J�`��|��A4�-G����н�Y��Wq��Ex�6!
m|"�3�����Ĥ��ri�}���I;��[�D��z X�D�|�LN�'����{$d뿋��`�p�d�=����楻��G?R����:��I=���@ 
�� �1����2���}�H	�W�!��jAf5�Y�$�����gkU1�E򰆣�v��Ue��m���FגּQs�wz���;X�C"���Pf�t(�<���㷜E9������1��s��;}\p���l�y��;TA�E{'��� ��(��Ǥ�c=���t��U��0�@%Z��`|��f�dW xg2��	 �{w�+��2�:�7�K ==���v�r�ֿPS�L"��8�`{s{3���Jϣ����ߗM��NR�t�!��m-����d�y��P�r���\%��^~��O�˝�c\�)�-�wɂ�Ǵ� ��ۛ٘�f�s�/���H�~���i�5E.ߢE�	%�	�v�ϒLқ��>�E��ƄAZ�n �7�0 ����b�No���6��n T21����" �f��";}y��5V\�oe�@$Y�M�nof`NWY��E�I B-ԟ�틃��j��	��4�^����>[��������F_J݃
Ž;^m�M��^�׻d�c\��AgN��ڳ�w~�9��Xi��T�a5���g
{���O�����&8_7M���DMDUDC�vf  �ۖ�f���d��8�U��0{7���!n�$��9u�N�$�E*G�w��� �<Wh���ʚ�����5�1<8�=��}��V�$-��'6��@$�g�3 �� �W���<\:�9��uq�}���̢MT�j�m����.	�vd�Bj�S��k�_
���! U���`D�7;�D����T��na,���H�ch"j�;�N��1`| -�e��|���gE�]ޯs�  ����@ ���7��&�z�A��P�f�Uy�B͒�ڟj =w��`	�n]���W����v*=��Y� ���f|غ,��!�QjAv��v- �)����x�E�{*-f_�o331  B�v6��W���V�b��� Q|u)~�.AMg^��q+r�#J���s�9><y����g����- Y)�{	e���k�=�wi�ы��l��`/�X���t��=#v�S�!L+��'M�8uź;��)��\��7�l�6$�M���OH�<����M�1�7Y^W	�8)��r����sg�G��vݹg��Y�ܛ[��]�R�fz���=�Kz�غ�e��y��^����Z���]�0v6��N8,�wY����oRũ^�v�V�=ۆ�4��v��ce;;к9���=v�s���no5�=]{x㮍ϴ�{6�`�&��tD��U�?7���� [��l *�z�4B��u�T^J��{�'� �gz��A�se��a����\4��qR��e=�{Oϗ�  ^��� ��z�D4��ح�(����o^�|���*l�$l�\�Y��x� ��O�� u1��F��Ӳ��u}�g�L� +ݔ�N3�@�da#$�_ge�aב���޶�@����@������+!�vQy�:R^kl5_�Kj��"�rͥW�,ZA"w=�v^w����)�;`�^ܦ� �f�dG'���t����<D�G9a�!�n�����^�;Vu�6�R0$�
"	@d0��	BBm"]R�B��6�w����ݛ٘;=���M4�]yd "��M��r�z$�$�UHm#[���H/��Y��/=���ˌk,���h��Gk:!�YW�
r�a[�:+P��0,'oD�nU�e�xj�Y�g��O���<ݾ��"+Ϫက^����I%9����g�v
HX�
:�n8�DJ�M���SL A���� �=ъ%��:����"!��������ilA6]�Tt_�q�v��M�l0?�XD����Gv<�Ϲ:V�� ���ڠSSӵ(Q*����4V�nb�@Gv]A�j3�ד���gOy�@|��� >���j�d�@��2���%B��B�FqF�HM��7�G2�zƻb쓔\�͟g½��_~�oݷE��� ���Fh��>��L� `�eKK���X=W�I^l��ee �*�f"nofb,���PTB&B"j�h���v �>����U,v���N�;;��2;����v��v<��r���p$jE�Q�BǮ�� ��}�*�GE�[K�(�s-G��ʇQo)U�k�qt�+R�g;ַ�.�4q���p�#���>�n�-��t�a5P�&����x�}u�+�<�/.j���$�����>�#�V	�j㉒h*�D7R�o7χ��\�����&{��0Gn]0>����u��Խ�^����I���$�Ӡ�t_c�h���6َ*�>�n= }��31@dwciY �����{��+�2v�\�d����%�"1@�jp��D+�&쵼�7F�m���c�T.(��=���� �����v�}��춬��/ι����-j�)�{2"#>2=��V�Y\ۤC ���nb���$�9�g�(�(Y�wx�,"�t� �9��)*�C<���{XӾ��p{O�\"($���M�Lu��4 ^�����u���L��fp �ݑ�=r�1OF���2�=��
ӎv�:���8~��� W:����g`����#�<�u^w`T�x;4������Z�����:r�r{b����O[�պ�9����K�*����C�X}�p݌�ɴ�P$MCh=�8܁���0;`��y^.�9� �.���w�0�Lc.��:��h>IP��(PJ"c%���ӕH��ιOgu\\v���!��?\[;�����pl�,�@yJ�N�w�ʢG<�KŘhܣ�=�Y��/\��]sth��4m�(�o�3)��;��������`��ט�H�ٽ�� �,��rR��Vj�]$5�S�!h�	�(���" �Onw�a$�F�K�����z殴 
��mD����0iZ"��$��fv^f�C:�E���6�  ��vf �FF�<W��ב_ ��t�1�34R$�SP[G7����o�g���������U`y�ۆ��nwf` |-�c�����y�����<!9���]ݸ35u#�ķ_=d���Ù��凫��J��	�w!�J/8����%y�&�\N��/������-�2*;�m� ��(ɸ͍v1��e��s�!ܼ��펵�����r��s��OpcJ��ȁx)�!���;�g�������d���ד��G����yޞcgI��B����wI�M�vu[��u���_`������':+�}v�p��3i��x�z��7�1�hKqی��=Sv{f̍�ݍ�&���S9��ڜ%����}.����;�F��ワ^{4;���q�=��۵ېA7�0�2" �Y��C�4n��&��D�5��yM0@|���` ���c�����߰��U�);i��������_�2��Ƭ�C����$k�W�+�*�~���� ���� �*n�`^�{�����d�q�2JB�K6���{��-��0A�D{�E_�ޗ]�H������>�cl������@��p�~�����6T? �c�"�@�����f{�gH��*_S��*�̻'���h\�� �eش�AZ�M&G�b�_��P�vn��!=�6� Ey�[@�K	���u�C���:5�Ϟ�KVč��iɌ v��s��M6G���D��	�������O]���Or�Ȉ�콫�A+g�:��O�|�s1@�Fw��X}k1YĠ�����x�BIG�����DY�*G��1�_�T��7q��jy���p���^���W(Ð=��_b ����R�͢��"���5�s�X��f�s'��I4OFw��@W���DD�I�����]۳�{t���,$�L:-�тU6J��Φ� ��2=q��v=�� ���Y�{:�@z��*��P���p�}��b,��^�� 63�݀ +s�က[�����9��k^�Ib��VN/�KͥMXN	D��9	@|��y�����Ǆ�yS�@$ζ�@���8�h۾���坷�7�U�زb�8�H�o�Pψ&���a�q�n�ݷ!���i6SB B!�f��!�	*A|���0A[���" ;wݙ��o�"�87v�-��L���:���x��F
��V���"qwGۺV��UW�D��᠈;wݙ�"<��]�k�о��mP�C�*�e7��,��i��$��<K �P���.�S+���E�k��Z]�|��^nˋ1�)k-�Ce�H̩U�X�1Ou���kgJ�R-H Ob�]ۥ���Y�����:2[̿V@�l�Gd������#-z��x���h@���<��W50^�Y�,�c�����e�A����X�.��aK	��ޣvAfY����6%��{*r�y�rS.��Ow�#�_�^v�N�>m#�);�Wd���=���,���Ә���i��*����B1�\{���ZF �L'vK�R�5�`%�pp皡�=��>�MC}'�[խ�*��lm
Je�h��V֛����;x�=��p�h�b�������+�vQz&n+<���᪊�}�����t[[mk�u�L��Ww:�ٲ�c���mj��e�n�CÐ�m�<pc�] �}�ƶ��$#`���Һ�_��T9Nĵl遱CUg����Y�����o�/�m<�?xg�m*P�+'S/]Ӝ�]�n��C���O����N�ҁG/�K������ʬK�۸����.�mong�x��/Iv��|�sH�NsZ��τ�{���*�TZk���E���}�t��єfX�r�}�|�9�qx���(m����$m̹jgb�Ң��vnSS;�*���8�,Ԋ�f�*10 u�.Ij�q��V5#3��咞�W��M���p��Փ�콴Sc��N�(&W`Uy5 l��;-˩ j,��7[�A�s=;Ú�dzϺ\�D/�5�`����7*�[^��Ե��H (��+X�j
��JTQA�YQ��eEE���b1��KkmR�[PYZ
"Ԭkk��+hV,U���X�eш��VT�X���QKaAX��X��(V�Ee�*�E��Tb��(�QPbE�-*�D�`+��Ȫ�"5�R���b)Db*��T+`��IDQ��Ш�EUR,*)YmQFڈ-�[J���� �[e`�F�m�,"�QE��%AT��AIQDE��V
(��
�mV,��PX�+X�E+EEUQDX�EV"����l�X�*�VE�,�iQEb�TX#T[h�*�+T����m��Y-J�ؠ�QE�V(�"��6���KUb�QH��[H*�U���b�b�l�EQX ��(�
w�w��i�n���/����28�q��C:���ږ�v�A�ަȈ�彾���"'�癄^�k����8 �����SUN�LI%��ۗ���Hg�*���kA�蒧���n /w{�0�y�s^�ӟ�fD��SZ(�,0�t�<k�8��/]�x�C�ɳ��H"0&�p)$l��so�J���5���SL �n��,�#��.Q3.P�[ԭ�XSm���I5���{�%i�j4l�J�Y��IW�녪�_��«�~�Ϙ ���π@|lgy�C\g>��b��k�h֠�ST�"�(-�^�v8� tf������,�y۹٘�@|lgy�a򵘢�"QQT�I%��r��띚#���q�` ��w�0>���"�2ʛc��uN�XG^N0W/LgnA�Ѯ����vy�wbڷʇZȧ-� �r.�B�Kݫ�gd[�h;��^��\ �d�fa'�ܬ����E��f	���d�$����t�j�$�wg� �G�$�1��k��d���\��
�@����l,puq�٭�)ԩ�^��i�&`��n!��_���$a��0��{��۾��H�>쫢$���ʢs ��$�vK�z_�0) ��r�R_���Ƅj&\�Me����/���n5iԋҝ�q�"�o�D4O�ͩ �"�,����y���x.��@*��[����K B\�!�q�u����h�y�@.����%}򗏮�V�pK#r��Ī­�vd���}g{ @���i�OkX�v�vf�H^�"�2\����:6({��A��-Ev�M~�d��vs�)���ҥ�/.�Q>�v��/���n�vf S#"�H�]ީ�����-p�o>;����7�0Dwʵ,��:dfd��f�ݿ� +2��� g:�����q�w���
��w�8�q�]ƃuw�ꌛq5��l���
�8��@�\ Tt��/e��quy�]���culg�W���7�����;X�hz�s��u�n�F�i�$+>.N�:����<���m���t�M�h���Z�a�/[�s^�E�ys���v�)uK���y�oa֩ݞ�ۘ7+�;�����8�զ��(=�d|ɺ
ݷv]]��8$�����]N�F7]���nA��*����ق��2�_��H̒F̆=����"�^N� ��٘�n��v�.�k}6J�$)��R:�M�����v��ga$�3��0<okݒ�0���̈h���� m��ѫ��8)u��i t(��516��L�]*"I'{�� 2�ۗ��M�e]� ���� �w;3-�M��L�]�*g[�]�p���I,w�q��nvf s9ľ���ߙu+N$_�eXJ�	dm�1��Z���ϰ ٛm�.��a��t��<�ϭ�C@n�vdF >�si�q�N�-�=��`vI��,���ED��c��[3T����ak�v�=W�xql�7w�~��S���D�{��enSL �7ݜ�`  ���l#�5o��Fz��H ���ݙ�;�y�m�#l�a�Go���Y�3�C�����I�s��8�>c7xtr�����uz-����+l�X����m@S�#Id�3�̮�!ܘ��^-����*�������ra� �{ݙ� ���m2 u{6����ε8�g�~����PASSN�_n�,� ���! �Ď�4�LL��9{,i ��fe�[�ͦ/(�rLmD�1D�W.o��츻�Œپ��I�H��K��=Y���Y�쪸��g�DN���A���uH�	H+P�:��H%��.����:z�;��>$]��*�:��Bwf���J��ĉ4�a�{v�'��=�n���pݎ<�"bt��o\�4\/}�}��35
�DPdV�����m� ՝n.V�ƕ�{�=���A!ng7�-b���U0�aIE��ʸ;�#�ݸ��^�N[��  >���o��Ϋh �/'�C��o����(��I6Ҥ�b�Q���bQ&���O�  Ι}�*OU7�C���u�Ù����¡W�1���\p��{~��b�ZQ@9�  ������
��9�/uҊhX}q�/�� [��d |�Vu6�*�jeTR*�5p�G_v����^zY��;ζ� ��h�}َyWٹѝ��D�F�7�T5�:��&�"�J&_��a���sİ�{^Q��F�1�����q��o�3]�?_x�Ƿ��Ί��y���u�=۷ϙ�JnA^ۺ��S#��(����Rx��%4~.A�����" �>�r$�}ٙ�gU1�vcy
=�z;��V@��O6�>�G(=I�A�
���Y�I��=�
�t3�1<� �d���o��x�FWv�/a���D�Ȋd*[ۜ9 ;��n"0-�xa�:������[�Q�ݐP���� ��L�a�4�,J���ߚ�囹%
��.@Wwo�	=�v�^,���F��4:����:�b!�N;�WAZ_˨�gDk'E�K���R�{$�CdY9:��{��7�V~��k�ӫ�ۂ����>W����E��89�������O�{ۘ���ҞvU�H'�n�X�����HAA���_;�+�q�n��r`��)n��=S�Ŗ6z�����{G�g���~��?�j�E�L��(|7�=s�B��'�;[W6v�Ns�sd� ������>�iV�
#�$E��|^�2��ݐH��n��Y'M�1Dn�1�9�뿉�k�p��/�=  �n���J�g�otH��u�$�7}B����Q"Fai���jq�|�l�U�A?���: �U{��SZ+f}��$^XJ�BԌm�$�̺�@s=*d���W�s�{�z�U`$��k�����w)�ˬ>���u����OT(v�r�^�as��i�6��LѺ�8�Bk�A=�;K���ü�=w��!��{#1�7���͹�g�T-����ݎ��A���]��l)����C[U`s��f��z����Z۶ͼ�ewkt�3��k�2���f]����;�w˻/S��p�.�8�Λ���3��Gъ���	�Şxە���u���5R��@�q�4tďON.��9�\/q�s�'�j-��q�����-�Pg�=��a�1��)��s�`G.�ۓ���m쀺$�p7Gknk3e]�8�r�s��c	b0D�!2)񐨠;�ϓ��!##��m���?뽯��~$.�u�T/�zAT�{{�`�Aw�(��a4Z[I���W��J���|<=;��_ޠ~>����_V|�{7�%��s}�Ě�y:��[(�$O�THY�˲H�׺�t�b�N���I�w������Up�ɎBd�Y�o��>de@�"$5u_BH*��VOǷs��Hl?;z<�Q%���<R
(�P2�o�zŐO��vu-z7���A�{��$��}�`����	���������A����5%u�l9�:��c{=��t� �ҋ�6O{�\6�E�;�/��u�� ����vW�k�f�=��w�v#�*�0'H�௺wz��~7}��T�*>��J���|��{8�\ʕ���e0[����3�`3�Vq��1�,N�C�o�}�I�R2�3�Э�b��_l�h��m�	�m���6�Ńۻ�`�n,��{��"UIb�i��#�&e�2������G>���M��GB���x�~w�vA��b����-4�2A_�����c�����
"!w�y�k}H6�D�S�V���Y�$��1U����Iw�[����-k�H~��goU��w�X�{v�F�-M��p��.L�4D�s̕���\��<��x�&��w���ң�Z��'|t�P���oP�MT:O;L��<k�Ʉ�ë�w۲G�s��7���	G�;~c<��|\�ު���dA#ws�X$��(�Mp�������Ta���FG���d�O��P�h������(�t����r���#wr�x�k�;���]�fhH��8�G`���+�L�A����^��oD�W��FF��oĒ;7:�N���݆*(6�9"���+7�P���o�@�f��DU|��H$/_u��^w��
������${�m�Ěx�0B�H�$Q�����Gt�!�j[Cݒ\�B�u�_�ą��.�=^��}���q9$hI��8��0�i���㭀�<����3�u��m�;mm���礡# �ɋ��g�n� ��yB��G'zA��^��c�����|�|+�2�1c_���.|���˲	��F�t�p�UOV~$@9W������"�D�f�n{a[��@�q	n��J��]�OŤ�OBh�U��_e�	 ����^��N=�P���0Y��_t����j�.���B�_��3e@n�_�U���pם��Oi����'�½��^�8�5��<�ލ�q�<�W>s�!�hNmx|���7�zw��ͮ��Y�јVu�g;v�{~����c��J��M�E�%��}
����rnS�sslh3k��J�λ$�n�_�]N�S�Ǿ�li�Ai�!f2�b4B���4�0�[9��;>�	��l4��;�Ϯ��z�7ib��q	�h
$���V?v�u�o��sU��q���Y鎬&�S��&��5��������O_Ug=X��Βx�B����>��t�P�z+l�1t����X�ׇz���0C#�oo�����H3�7�-�� VmՀv{�һ��'�{"�v�*�!TЩ��m�Ք?3Rtͬ�߲\� ����*��t���-
nNFP�@����:��"�R�f)s�� �(VI�7|$���Π;�]�����ڊ�����$�	'�$��	'��B���$�	%�$����$�`$�	'�䄄	'��$ I?���$�Ԑ��$��	!I��IN�	K$$ I6$ I?�	!I��IO�H@��B����$��H@�p	!I���e5�zߎ�+u�!�?���}������( P @  P R� P�  
D� �EB�D	�REUUT@IT��*�R�)U7y$UTJ�$R��Q*"UUED�P�B�% ��A` -AH���#��oN��{c��gNz�t�ɮ�-��窽�kپ�T`{����[�X�׶�]�v�C�ܣ:����%��}))���"R"�оyA���f��=3��.z�l5��@��g������5>ET�� 
Pz�z >u��#l t@4 wcv 4s�� {�O��ѭT٥r�E^�کTT�B��R�F��#f��ޤ�<�:PT��fu�7�X�v1�I
_�����n�a�R�E*��=Op4ۻ]��W`5l�����>�*	%(8�40����]���x��Q/fz �g-C�
U��!�=y�XC� �.����4 �J�O�J�=�	�"��(<��`��YW@P�gMvta"P� ��A�>����)�䛈�{-�δ�@ٕ�      j��	IJ�&�b0 4400E?LR��       fUI�J�=L       D�J�QOQ��F&��0 &��`����1J�        �I��0��(��z���h�F�O���}^��� ���&�y�����ӷ�B�T?��S�!'��%   !���$����?�jd�!&�^����O���O�4���=TPa!�$�!#
 v��	I�d����BNO���5�|�'�}߯�?�� !	:��;����\�p�K����I�켳��gp�
X#����O�����ڋ���ؒ��M���UR^�Ix�=��0n>DV�r�x�����c%�)!�d- q�
��s�i��[��d2�PZ�6�PZ��ށD��u���Z��ׅR�x�<�p��E}����I�2J�h���f����s)�-����1g79t����@4Բ�}�J��`�5�zGσμ�q:�M���wz^�v�]�lp��i��sX�q���n��uD�&���7�5��b�G�Nv��CrNR�Iج�0Jn1C!6,�˹�1ݬ`݋
"�������riݥ�N�\[������t���04�1u���\�KA��̗q]��C��G�X�q�)�Wv�:��m6�V�%A�H)�؞\�vv0�]�Ԫ1�]�Mҍ�j0X�,�Y�8U�nl裛�m眠bl�)+:���zpQ��MS 팹�>	�o�3��tLO��Y��%�u��9q$�LT�͙��q�f<4�'![���ь4x_�Atz�ᩀ�Ѡp-�Tm�5^������C��mK�vP�Q'�`]g�oc��9���ߎ��"��܇n���_l_h�7{�f���a�o�]�q�V��������Jqʥ9�X7D0N�$� �X��\;��$��?�Q�1u	5i<�q���qJ���l���=k��Oz�%7l(��f�WG��ܜ-d���"u�5����� �]kn�Y� ��;J�^H7��D�yZ�2̝��e�N�nV'](p���v��k9B���X������[^�!V�V�p)�E�B��zp�.�ge;x9�h	��شa�EY��^�S�f�7;�/�j=�..崷OB�|�e�oJT���5�b����*�6M�%��y˭�zor�U�b��Q��{l�7oDD�:��y��{���#;��PQ���Ft[���He�;��ϏH�xP�K�d�̃�
�C���҅�6�f��Y����������Hغy��{�&r�^�K�����V���
��!z�
�ɘ���G�s��"gځ�Q"�Ry�{���J��+QovBxz��v�r���GG'V��H�=y���Mf۾��ĳ{��/��함tY	D4�i/��v����vm9j/8�DR)�O,�m�	8Ϻ������M9��.�ה��Pk��v�к�+��9�1�6�\tf��s>���Njn���g&�(|�tU��GV��n��H^n�K5Nz����&Rx��&���c��V��A��WLDig��\Y�����r��IR4�E�ͫ�S��U�X��P�%�l�tS��=gV�H�����V����;�d��oc]���;)B��Ns��-��� K���k:�ܦh�J��+�p��4nv�KN���]�łN��߭�B���nꐥ���w��..�˦'�~0l{'�7������2';wVN/�E�!/!�6*��n�8V��t���3��̉*�a,�H��e2���'MnL��uM��3���`��]�8u��A�Š;9;�6w^�*�z��w�y��G��A�߸G, ���W��n���]�x��*}.��o�n��Py�$���
:2μhɅa6u���}�:0�*��!� �����A�����Ӫe�a{��ӷ d�u�\K��]!�Y����C���v��Ϙ�2#��D� ��4�8�f�ʜe(;�����bj�9e����+�K���q^�[�GwV.���3.EU�f�ɍI�� 7��[��o�Z�� MT�v7ʸ��PoP�����b�Js$��7M��=�p�@�-��s��< C�^�5��r��P#{,kZ�%�8��"
���Q�0ݣ���־"� �ދبv-:�:���/�Qt��t�����a�~s$�0B���˹Ƥ���x�J�<77O[�A2�MJ`��D+f^�v�GM�}
g ;I�yg5�J-���MH�֣�m/�sc;Nn;j#f:�s�K�	��w#r�c�lYst�u�Z�)`ͳ5^��Z#�Ѭ5����9�a�}n� VoA���
��1�������=����]�;�1�m;�N���';���n%E-2�k�����z�YJ#�ɽ�B�jb�]kۙ���uݫLl�q�Z��狶L�_���b肱��g%!91�VcY�6��l�q8�נ[�.�Nm�ъJ�SW��cRܗ���M�)"��ʌ�-�ā��h�l�uᡦ�|ڻ�w,o�� ���u�1��=�y�ع��\�`��֞�V����W�.!y:TP����wx�ٵs$�Ǌ_p�,!��ۻ��{���[�3�f,��A��~T'UI����F��Vv@i��<�ѣ���\oeg;@b��L� ����P�x�뽼7��P8%�|{v����8i�v��w�o�ԧ�:2��#K��mRp��z��_�G�i�Dp�*�����t���ߕ�r_�'q�2��5־�LhS��r�"ʪ�g_n�"�RNܯ6����Gh,�7�f�QB����sG��+�ٯ����{��o�2-�\3�u���B�����Yui;;E�z)� P�����Om5�z,4��ƌGI�1X�&��j9R����;U�<���áy/�3��6��r`:���8O���Rp���Y�^��)�� ��u���6�BqT���O|p��83o � X:?�����Di�z�@Zs��*��!F]��O:
��^�-�?���cXt|�:�A��M�b�X���2���J���=���L�;]Ƅ�Q���a�w5�q��E��wkh)Xi��:9���X�E��y��Ѱ��P�mf�V~�|�R]��QD�E2`�l#��ͪ�uNhԩ��6$#p��2�7WW 	� �Si*��L�s����t�:OL1з�՝�w�j��e�̛�F�k
��gY+�3uf��O�`�]��`�i�9�u���j3���3��[��{�����o��͝ƣ3��p��b���$�[j��q=��sc�/=c\O;������X9�(��u]�k���_ ��������5�]��Fh��`���	cv��,�:E]�����q���2��bDbq���=/,��&x�a�D W�v]�X1�6;b�c�����~�~ϭ? �����Js�����=��|x�sl>�qNv}_OϞ���	!�� ��,� $ )  �E$)	$��!R"��YJ�@+ @R�R
� ,����I,�!Y$�I"� E���%`,�) �!P�$J�I ),��,��� $	
�B,	+!
@� 	"�H$�XI
�,$�@B,����>g���|>,�|�>�~H��� B_`���pI	>\w���i;�Z�̆� �$�G�����Y~��z��sG<[�ַ�V� �z&��C�J3�y4#�/1Ҿ҄5����ڽvZ9is�N[^bw��?N�F^f��-k�r;m�r"��z����}���&��cw���/J��m.��^X;����T�	���Z�}*X+�����ݢgz�=ط;}���K%:�y�n�Oy8�8} ��zF��Y���тg��.�u�0_}羹5xw���_{�;�7^k;��xu��G��<���������Q/a�h�~�Y̱י�n�f��Z����m[���W5���\��5��ηVm��M�� �ԟ{�1n�x,D��6q٭�e���g�K�h�.N�Ӌ�^�ҫ�2%qi>��Px�E�/g�̹���^�L��vl���ݗǗ+ޅ�{�@f��yO]�}������[K$��5wf�V��Z����
�U���X��Z����[#7�.t��wlz>za�f}�$a�r]WL�b/�frW9.K��L_u�JlKy-�u W��0j��0��]����ˠ���cVҒsx�;��W\酎�YUZGi��3�GI-٪1F�UL"9�s)3���;�Y��I��|w��+$L�[���{^�2෭�'~�|.��{�4�X��x��x�+�I�����=�DVvhm�?+�9��d���R����� ��ƣm�7s�3R`i:�t�ME��{7ï�8�S�zrV^��vfݘ��x��#:(G|�c,��,��#if�{��Gv��[h��If�
���R��}�<sfqy�/@��'>R���7��ʜ����Z0 ��9Zg5=J8��ݾ�<N�2K�Є@��k;a�;�o(s�p�Wr��V�F������[M�y�X�hi� z�u�:w��&��{�]g�0�lG�����	��X�Ș��˜���#�ۓ7 8�Ԁw��e���D6I</w&;�mr�9�5�u�d-
[����'��Z{27��gCWg�5�IǋT~�,90���|@�i[��2��h�i賑Jq��|��JX9\;dT�n�0Cj���;x�[�����F��(����:���,ԕx��5z �����|"w�:W6D1��9y����ٲ���U*�ڔ�
Z�4��iJ.YԻ���!J�S�*|~փG��ٗf���̴�.�����R�Vim��ՙp�������Yl+FI���F�.'OQ����#T�jp]�jbhG��_n&Y�|��=��fO�ul�����O�d˪�-�wڲ�<�B{V{�6:G���7Y/��ީ��HFW�p�3�c�tj���S����	�őI�E�3��;��/�^��(g�j��EH�t�YL��i��_M|�*"IIN�ӍU��0�Ǆp�6����!�v���!����u/v��$�+�p�\�e*=Y3&�.�%%��;:����x�S���}��j�#ٽ�96ōz#3:LjYU'V�̣Nӂ��۴ފ譹M���=\��ݞ�i��I9��=1n����i��`D!2�9��]b+z�f!�c���ך9=������%6H+kyt~7A����#��I6��c�^��&���	2��͇�]���D?{�<u*�]JwvKz�͆��r���i1O�ʙɹK��%փ�	��}����ۄ��N^�M�.e�Z��i�V����U��9�;��f�/�I��ѳy�w�y�����[�Ɲ<�&����JGÐb�*h���^��� �R��Ώ�ĢW�7���[*�v��\c_/?����7s�4�y���_�v�=�/�A"�w��o�(é���g�	�TP1�֚V�J�,���$mM��s`��{�C�E"�i�)����UY��D�W.E�7��;.yڹ[�L˥�ĞK_vE��0���}���B.�a��4�b�;�f<�y�/��fR(t��v��4;��y�%,��rM�w5��b��{���7*_l��@���wh:7E^��;�??k��qd�B���au�@�{`�}��.��>��Q.�'���D��X솬c�e=r=(�[&���T{�eI%N�.����W��*	��r��x��u+p�1�;�&��,	��������a�y�[�TWrE��P�9�v�[�t����q+���
�U�[��J�.>l�՗[/ngdY5�'���c�Y�e�~�zb]u�"W(\�7���#u�yuD�(�u��WwaH��/���RYZ��1]���'.���Yx+1�b/�e����.omP���EX��v�Ⱥڧs4�x8\���>����&U�`-��H8��w!�^�`�1�k鍎G9͛�&=��r49��Ş+����.�r˾���K�|LI��M4�qzbG�,�No��;���U{\  ,��x�N����)8�uPh��5Bj�Lؑ��+�\��,��Tূ��rL�:��cv=ʱ�_C��=ʮ8�C�N���!�+�A�NFŪ*{ݝr�h�Y��/<�C�ޕa������K� �DU.���T�Wv!�'��ΌK��Crj®���uC,��?�D(�w���p�W&�9�t����ֈ2+Ӻ�1p�b<���]��VuT\��z�1�M����u�;��wP�*�h��xn�W�3U0t��Ry4Qg^��O��D��攭<��ُ���N��۪�.η�%�;MP�����vj�q���;�4M�UP�O�!�i����(6��s��1[���";o�I��q�d���3�zt_
���{��ϙ<lӏ�ļ�	�.�Z���6i��|n���Kݾ���'NنX�t�kXe�2"Q��㺨#޻!qJ�x�Etg=�(������U�sǏ��N*�����D$��A�;U`n&���֧�hS&��N��Z�D�#镮�i�XIzk<н��1tv1�r��x8 ��O���V�[�;{�0��C����4�E]�[툲3צ8]XP˽���c��YQ���vn�!����dմΤ���u�Ɍ,[��*"��}e��=����Fs�1&�WE���.ި(�+3�Y���/��{F����n����}�u���b�����na�ޚ"�j%̨z��jꃮ:� �/hr͔0�-Ul�"�57����V;�v8�����흠��%��8���r0l�d���'P������r�]�Q�9V{s]츧u�p=Ju8gZr��J�:���K�#�,|�ٔ�ړ{�і�+�
�v�T�U��K9���������XE������F��'��<��/t&��zߐp��ɰ����y��O�wn+\\]���k]���7��rZj�d����]�lZ��Ǜ(�31���d+	�5�u����O[]��n��=r��.z�۱�y�n�I��i�n͍x�8�R�]���:�n�*�s^���&�K0��1��������J��UW����ѱ<<�R��&�;��nγf�#-�4�BNv� �,k�{v�/Gq�Wv���,"X�R2ٓr��H4ϝ̑:��6#K�9�Z
�S��ե���	ʜh3y�y��;v��7�* �H{ln�a�6������,�ʇo2tL����b��Y�#��Ζ5�qjKn��l�e�ęcY�"1�E������iWɕCn�ͦanZM`��aܹ�[_uٮ�{c��!v�1F�=�V��I��c�R6j�`c9��'Y�pQ��5Y�liT��#4`��k�읲W��ێ��)�7u��p�r�;=f�Uz�ѳ��뵰��Ů��q؃����f�5�bڏ9Җk�������l]cV@F%͑�pK�q��8��%�b���^̫����=n�F��6X�+�]��q��l��R�l]	J�5[i+����)�Bk��+�t7=�rs�������	�4�QqTKKu#�M�j�
�İX�^�gͮ�\�}
��</kl�������nCD4�q5�c�ǷR����]�&N&��.�Gl^0���/�C���3	F[kH<L�h(^r������fk��ojKs���1�i�rg��u�])��1���'����`�c�y�e''!���q���4V2�f(6�bKgc��J䛞{oE@�\GX+Yx�wh�c���Ys����*�t4)N�{X\C��jg:��f�u�v&0l��%��ʯ�!�����{cSFb�K��A�k�Bc��b]1�{����Tr�=�iX�14�BR#qS
`d�FP���[,JUs5��+A�VZ2��V]�i���)��Z^�ӟ#*{ ��^=m�MNN-�m��E��R]�k/����!Pw��k����2��8�,����iڮ�6#�aʶ�q�2 ��]Ź2�p�n���a9�y�h͜�D;6rJ��ζ<�@x�s�m�;��P�q	uyѺ-���#
΃p�j��7 ���R��Z�du�Rh�����rui�#���s�Hh�AZզ�)K
i��u�����+��kcx���:͙�v]EZ�m ;ud�u΢�>Ǚ�T,*�YL�2۱b�뙥J�۱��w��Wc��.�ۉi�nH�	Rde���2�-�eK5-�L��[l��V�������K��IMx�o4s��s�}a��9������0�u��W[�zb�2&�M��	��p��ˎ����a����ܛ��v.���:�ˢ�5\�-��6B�4�kB�MnX�9�����b�[H�W�m��YwmQe�U���*�sbA�΄�s��7)��N�u��W1�N��˻;<�	�v3�r���D���X��m��"�t�Ƕ�kWm�aՌ�͘�"v��q���Hs=@xm3�ҝ�;e���v�CV�ՕZr���U�4���c�9Y��E���\:�`-˧�e�n�&#q�Y��r6��ͮI�ܯ�Gv�sr�;4�n�/e*�[ ���45e�I�qH�g�݇��i� Wawg���6 �J�t0�uٳf�bq�N�����i'��śc�\9���&S,oj�9R(�/n���3%�6�ak�.�t �l�Z��:,��
溛V���l�:��b<9�%Ik�F�lM���� �&�c�A��[� �Yc*�X���K��rOOf;����-�zzíx�8]l�	&�m���gBR��HY`�b�v�zT�`:�9Ayn�g ���^G^9�!p�Ɏr�uZÊ6�c��b�4�c�S:en�vrmƈ��1.��vC��p�,�.�M ��L�G9���	�@�5�0%�;gV�6tV j�R�z�(�P��ժ�a�9�y�<��ň0�����n��Ir�ؙ\�V�D�,�UUUUUUUUUUUTUUUUUUR��ʱ�����ҫ 멙��vb �d�zѶ���k���̸�]i�^�L��M�A��J����3Z9�e�#��K��l9���7\��Ncr鎺��w�#�	�n��8�@6;v܄t!�4�Ѳ��-�@��=�ۏq����8p\��j�SUk6T��0p�t�[�6�yv���(Wev�T��W��[a��l%�q����C�,$-�\h�:����k��o	 ����d]�9�-�u�b�Y�:ݖ)��tff��/f{�z�1��1I�@咰�� �Aj\�Q�R�U ����m�"�츆5�PUq1�(���ewB遤�$F-��	��jۻ���*[Q����-&[U�X��TR�R�
�q��M8�E��PYYP1��b��1D���*�������$���Ԋ*[#h%b�i*("�*Ȳ颂�H�����Qk-��*@U"��T^3(��ڒ�Q��V`ͳ�eIQE"��$�����%2՝	���я�<��P�M���
���©�&(�;gw�v6����.BU��ҷm^JA8ݝF-�װ�J�r�t7��B���lv��є�b����aR�9���A�y�x����a}���A�S��n�ya:#�x�jii3+�f��3F��ҶX6]��aC���Ee�^h۬��b�%�Gi�ӦB�5�M,�yBX�Vc0if0CaC䖚Ȭ�c]��҉���T�0 .n��:��G7����d��zʽ��]kzqȼ�Z�8_qNn5�Ƈ�w/�������pջ"���kq�x��8�6�s��!݈۞�E�#��ܻ�vz����=g�#��HGvu����0л� 54�!1b[��pj�	.f^b!�/i��X��ڕm��ښ��a��SR�>�hj۽[�T�nUTUf��v�%���1I����WI�c�;&�����4f��.s�`��'{Y;D���T1ȼ�4<��(�\�'7\Hץ�.+���W��fy�Zn��2B��GM�����(��+E1�7�\�uL^S�S���"��j������'��w�߽ܫ[R$���5���I����1p�N��.��.�n؁=��[`M��S8�>���(Ym0YP���V���w���Y�(���+k��Vr�A�0����Q�A�5����Y$No$�׀�I�	�l�A�N����^o5��Q��Æ-�ӓ���"nw�^`���I��D�	;�2[��0����O��ma]�t\+�o����/&@�	>B�է�e\�9���+��h27P`��si{P�1��6ʎ6X�PcL8fCz�0�8�fz%U*Қ�oa&�[ d��g����d}�	EI�М%7u�VņH�l��7��H=�E�y^��y�we���'�`�-�eI��|�Om0Ț���Aޫ��e��$���q��r���MY��ql��1v��wI�PmD�'A�0|��/d��mپ�gx���2���);��:�����wɕ�P�1N�ovzaʸ��0G�-_���@:��Ѭ��ݴP��վO���8��0�l׾��32& ne�ڀ]��0a��*���44��NMB|[YS��8[m���=���謍���W�_`3ɐo�3{k'��G�%O��1{H�	ן#�����'�H�<�:�o%JSQ���=�EYIwU#Dz��a�]b�o�|6���d�H�N�ݣ�%��"�2�y?⫞lG��ɐQQ2A5��s��h�~}I�0���RmXI�"�M)/s̥�j�'��_2~�c7�6��kF���X&��������C��)�	e�|�����]��G&�0�3�"y�:�[�w�kg �K��b$�gt������KA�Ǉ�Sӕ��Z�RD��:+0�vF]�ՠ�c�a�V�����K��!����������T3��w=��������Jil�Du�dk���t}z��a�6j��u�!k�fcA��zaN�\�V$ͷQo=��f�e�2j��[+����wjz�5�2ܦ2�]3Gl5#(�	H�gSA&��ɠX�$H-�X�}w��s��hQ��𲅱�Uyn�	6��"�-��L�y��Ӏ`h fب|^Lqځ(�v9%T�G;yK�	�h��Yz�K���]r�&�����������m�Õ�-�ꢎ�9
�G��[@��0�l�9{�%��>1��2&����a�]v��y|�|��7�����=�or�H
�
�D����<q-�=�<�	�5X�$�]ͶM����8޻�-�n�E��w�Ѝ�b�-��#��e*#�z�f�"���L�wP�L�0�f����kuu+�b ]��yw���L�L���oCQ��Y ����n��}k���¬ў��$��f8�e@�H4#��$��.�o�m��v� ���E�e�$�"wWP�f��
���foӠ-Q$���#1�B���hl7h�OѲ=�߿R�_]ն������m��s�o�ǖ��^ ��``���`�)}}Y}l��+��wVˮ��+�߽~�'�{�3�&�;��	�N�&�mݎ��;�����\fId���ZnMHE�r������2/�z	y�����a�i|��OlmxFܿ����ˡW��@�Ђ����� �T�2%Q>i��y�M���<e�Y蠇v>�������?I��j��a5�QCK^s����_V^r�Y��;�;y�g�sa�*�>e��Vz�4(���"������\�C�Hχ�OV�RR�%������<�+���&I�g9��.ô,�v�7l����謟��5��vI"rd���+�{.N�T6X��\E��23���foz�x/T0/!����Ȟ<���_�݆��^i�앳��ī@��d>�x���/��0�����:�`���hG�d����?/�9Go�=Q�� �v���)���[�{6b�8����82��YJ5)M4�j���VQ��[�kU�.,h���@�j���^�e��8���ö;p�Fkf�iF�G��k�f[$��b�<`���^v˓F��&n8�3k��4V%���L�j�{;5�3��=�1�9���#*����r�X�����^ܒ��̃U]���	� ��a�o��vZ���5��0g�$�=�וא�FSg���V�ە`��=��>�ly3��|�b�X9	�	A�dJ�q� cL˽�!=�z|�{���!3��a
�M�n$�%2����."�I�"�)[��Qd�� �hA�C<C�:ښ���l��:�_wc�ѬY��0.�J��p᳖ؔ�#d���)5�����f1�Y� �]#�Z�$�ؑI8;͈8)��
f^�ו�d&��;�n��rbcNꊁ��M ��`�Oo������v�Fܫ�������z�4-�bۅ�(�W��˾
.0�Գ%Ή.\G:"�'���}�A�10~���=�b���26#q�{୕�X�rX�������~L�sd_//\�6��zGl<��� 6��l��@�����o��{���]��o���z�}���m���p�ku"ř7��D`�J�;��Z�����W����q�!"�u}��X�����r��7�d���wU�H�щ���򮽼��򓗨^��w�����a�~�ӛq����k��c/�E�{������c��K/#�G/'�B��Wz:�[fo8��,�3콳�)W�ÍZ�u�+}�P}�3���e�U>�I�'m�Ek�u}��;6]J���X6=�z�T;{`�#�+핶�j������g���/y��:ڳ���h�<m���q=
�^�}v6ŝ�|6yC��u���(������g��CWK��$����>¼�{�@Fd#dl�j�wɮ:�}���l�G&�Fp�OR PC- �x�EŐ,�l�h*��0��
�f�e�T��$�[IL�D�P�Q��E"����RE��PM�Qv��ȪF*��AU@c*LʌDQ2�a�Xi!���DZʀ�I�ƴ|'�Q�������.�ܤ�JM����@���0;�ϴuÿ����@?%�?'_~��"j`�7W�,U�U�e���d0T6�9__o��D�Uk>�p��a��p�+��_��ȕH�lE`�O!4m��q��W��
"eG���1m6 El��Y�b������H�d8q���fg��>��q|	� �������
�4�e�X-
��vQ�Br�Ts~����w^9%��>\.~�H	��2^^�����І�\�ibM�]���N'+3���n�x��g�y���C]�sl�zۮ3<"nU�.������@ �b��4�� ��(eAFs���K:&�BH���p�^Ol��j�<���`�v�g59���FF�2��b�`P�Q��ozж�b�Ba���z}�nn�S�#��|���39�(t�3�����֊�V�����ᥘڞCF\fBQT��P·=n�Yj�+vi{\���NI&9�v���3]����#�b7c �h�1����(�Kib�acn�]��QS[R�����ɠ���9Yn�u�b[NI3�~�$�Jk��S`���ܮ��g��H7i�zߖ�#�����z����LH�a��[��;qw�Q���|�9��"h��1]�9�YC"U�ݾ��'�>�1n�ܵ�n_1�Q���D�uW���i�w��O.�@����Ϛ�}����1�1(�M��DL�2��9�k����>� ���q�����`�H�lk+�$�K�w#�O>���}�vJo�f���̮#NJ�c���8t�;/%w0����я��\/��p֟�.��U�.�?�ˑ�_u��$�L�B��w9@H5�Ǆ:��EH1���n�{~88~|2������[C"x��-����j����)|�b�a�Oa�%��,BX�#R�����|*�}\�#i0A�0M�χd� ��͑��Sn9�s;5�� /a�/��&����Zd�Jz������Sr����]ʿ���M�G��=ܙ|����*��U{�9%��� �/���;���.G%���p�L$��$��ă���U7�r�$����G/�V�SF�[��Q;f�&�-�/��5�r��s�E5��u�bE�_s�{�j�2;��=�8
���VF� �A{�6ʊ�W0ʻ�uݬ��������"��6␷a��s4��
���S�)�$�O:^�)��I�_0w?�y~P%��;?~[{l���o�����)�M{��U����/	��w��������?���4�r~�`�?.X���&A�2;�+�����+%e�V�J�i�4�]UQeopj9~��M�L���/)���*аv��І��_!~��n02A�a����fS�^��6�S�Ҋ�W6A;I�i\���HC�� ����`�㙎�T�ˆ&�B���ޤ�bd��"��޲ҕӿ��_6I�0@$�&g��{��bK�һ[��:�p�w��7o˰g����K, {��<�+.���if!M�te����L� ����a�����f9��"�
���ڻ[<���S��2Si����[c(�Wa�TV�j�Qm�
=��a��je�*AU��[�,_�����$���3����L�m]S�K�f#v3�(�`"R���I ��r�1w�^�bޮМJ��hB͎Wn�ւI�	=�{dv�QU��;	�dsl9uwop�m��7aԎ������څqa=3}a�lA���=m����3�Xm��l��'zq��J�@T�'"�9���E'���$�����倪o�{��,֜�L��&A�!����r{�R���oK��m|���Mл��I�s�iP�*f�t�3����Y���H�ɂ?y2MVk�Ѫb(�|��&�ѱm��$��������j/���dNL��'v��h?uS���W6���t�L��i�\_o�
��O�-턄�b�ѹ��3nug����dh����3��]C�53�V�RU�؂�<��ˈ��?_/�tC*�`'u�4�m+?Na�T��A<2-������z�M]�q�6s�j��8�]�"�N���}���k��=�㱟�Q����A���r<���}���O�y��o)ZP�k��� x���l������ok��l�Z�G?�}�}����i�6��wЫ��(���-��K/�6����mR�S�a$�3�����oa�	��$RX�XI��[���9��H֟=�p9����w�=^�ge�|��;Z��_���3{�*1�-�֍;����6���Z7����N~w�g9�u�Y��&�f�)��ðL��L�b3�_�
]�~F�Н�.,ш �Mp�8�Q3��N%|?>4!m�B�C/w/��l
��?g����Wu��6׻;޷j��F�K*�\{�mCn([p��_0w=���A?I��&M]X{"���vU`���$��~�[*�z��X_�RG+��I&sw|;��W���A�O�I�6I'y���'lt&���}����ȇp��s�|����î�����#M�v���������������{AuL��/9f�2��\t��g:�kU���# �a�[��}����G�����f�RJ������Ŷ�'��C��"�6k�����ՙ=�_˾�r�ߔ����LH���#�3�ۋ���5a�(��G�yN��;=4��|�/F.��7٫j����À��i�`�k,�i]����B�.�$��I��s��n����Ŗ�W/ �0u�,�(���v�U�6sO
��]ט�+Ʃ�.���EJ���}pn��@�}���MӦ\�zoG��΋�\��[�֎�]�(5	�k}�{&��֯���gtڷ:��@������ٯ�M�D�"�}��1>�Uj/�����-�T�*���
TZ���d5�K
ȤP��Z�P��B��T@P�XT%j���2�jɤ f�B����T�oVj�]U�HWTr�R"3,*B�M[�J¢ʐz�י�E3"74i-��z7\���-�9hl+Ee�.�n���x��ZPQ\J���!�l���a{-�s���U`�.�f�!1Zv�l�s��`�0�&���͒�9׵3Bmj.aB,�b^ю���0ꡳ*��.k��;O:�qX�8�<��Q�6F�� �>ޤ̰��nd��^�ͯ:���l箮�
˶8�t��b�fYemq�)�n\��J�)"��Z2�[�1Ykd®�q,��2P��J+׌Y�e�����r[n���XȜ�F��0�L-v�ځ��cElGS`MZ1�y��xy��N��L,niw�F��f+Z��C�VK�L\5
�1�Me�V��i��n�4e�+4�v�y2ʮ�#v4s��1(jwx�԰c<u���$-f�<q�޽�����Y;3��t[��ʪ��Ն���նR�@lp0s'm6z�vU���3Ƹv8�<��]q�T�1i�%tWZ�Kn/�H@%�p�q^'���N��VD�^92:].&�F�Ja�.%������3C��{u�x�t��g�9Q�L�n�M��1��'��o�fr���#�]����l�y�����Ͼ���2U���F�5�b�E�/?o�@\��j"}��}�vʤE��l��
bU!�k�9�\1�6��q_cv��*��Es|I'��I5�H���J/��{��K�mY�j�͈���d����q�v�q?�'(u�$����Gw��?v���BL���Zo\o��JB ���!E�!�����ww�RG.��"y|��&kC��Psl���O����r�Hg�;=C|��9��h$�Rڧ��^]�����3�*<n�����m�����HBI�s~_�h|yv,~8���s{���#��	����`�6�u���Uu�t(�^�G��A���$�d���%�
6����L��{w��[	�W��D����dB�I��]h7&fYp�a_�y��"��Z����I���}1]�z��B����:��g����=�0n���`>�n���c4��\�
����#˙5��;�P>��0בݦ�l��]u#���0�d�왓ye�{������>�_I�܊d~)��y�5���8��9G�p��ߥR�*a��E(T�L-���ƨ��b��x��]�kȢ��1#�h�6eXp�(\|��o�f��P��bʆ �l4J�����.�`�գ�)*�b������t7i�' �=��U�w ��'���[rC�I�+�H���Gq"�w�2n�^�~Ȱ�M����	���Z��Wߒ����כ���/�������ex13������B��w���s�.q��h�v2���.:ߢ��<�R�ЄVBb̅�^����q)��	�`�bŉS1r���^�h�&/k`]C�C6ר����- �EZ���
6����6/;��� +�̸`{j�����nNA�13Zg�iUCP�֭�[V�khf�k���LK�ηJ��� ���h��������}%�I3P�n��o�~�L��B���
{���]�j��S��F��d�ѧj���}��l�����^K�J9CwWNbc����;i��u��ҌPu�<�۶99����{A%]�SZ�2��;��nعԺb��aldsX�+
T�A�XEh�"��
����u[.���"ݠ�D�PI�5w�i���`w��~�1���ˬ�v����I��^YGo�A�{��/y�<mU��~j�/�%�_�l��_2[y�Q��3wuh�LL����e����v�Y֟3a>���W�	=Ƀ��1G6���6	��a,T,�_]*?n!c��g{��	)ID�`�mW]UQ_<��
>�gX���w�,��,�Z�SM/Q?��1g�Ӷ����[DC��r�v��ޭ�1�,�/��> !x��^?{W��Vi��R�����wՌ�(������&A��|�=	�
6���S��{�BA��$��2A�Q�`�{5�IX{?U)f����{ɟ��`����?=ϋ��y�~�E�E��UCA!N)��'x��@=_x��-�ޯy#��zy�r9VERbfҊ�
���FEE����8j���9�A~�ĴD������U��\���'���:1��}����ʓ�I,g�丹�e��6K�t"��q��X� ��;�/�X"Sb�=aF���d�ԾܴA{͒�L�/���Bv��"�Z�#1ے0Br!���?�Ro�؃U6A �!N�����;���Nx�ʎ��3��6LHp�`_��U�Ҳm���C���E����#j�$���2A���!�(�c*_m�I[$��[���(�1uoftǘ<�&D�|�߳¸�E�Įɞ��� X�F�L�]x����a$z�z��B�'u���UF�=ɌL��,yƎ�er-
>�~��ɐ�Ig�B}H3͕ީ@�&=͞��vE%�d�n�;H�Es�����.{1=7�GW�Q��lD�#73Ȫ�!�����Fcu���\�ET�7�(^�&݀�7�D���5t!�,�L�܅,��U;X��+#�ۆ�6b;h�=�ߛ���Xoee����2�v����9�������~����Ѭ��11׉�e{f,j��b5�2̵�	c��D�ۍ�G�ЦY��NvvI�]�8l�!Y��n�n,��Z�6mn��aVf�nJ�B��,J��#
g]�4{W��q�P�WM{EMH�PHd�H�����{���~�0��x��)���b�����O�(��{^��B�$��3ܾ��ۃvR>�IY��@U/��j*�����O�q0l���r����z�W������;��mJ�������ʲ*�`�B�+cuQ���v�N������2�PH�p��*�4E_>�{��1��y-�τ-��&W���Ey�l~=Ƀ�eX(�S�Y�T�s�|���;�I�J��鏗tj�,����ͳ�+%��|�י��v�~�K�}�@p��z��mNd/�z��ͼM�&	A� �� �bf��d�pO>x	n0�2�d^��V�e�x��W[d���f{������&0�a��!XhaRQ
��)��eH)9�I �������4�h�Ӆ�f0�.R��S_~��?b���gKz~o@z�B������� �׽�M7�Ϻl7{�Vr2T���4ĂÒ�����Ñ�M�@Ă�ǝk�<�ަ0������P9����R
B�{�Z�HW�|\\L`yG�GO�"�W�J-�~S:d�;⁈j$�+
�~�43?~"��T��b����!#�n��d�^�γ^G��p��w�����$2'f�7�<
��ˌ�޸�A�P�+��?^r���ҺZ^���xRÊ����U����k�����)@�*��;h�|�اW�Ԗf�;���Y�fC���̽�J3wsڬ��	û�m27\޽�XE�+����Xu�$n��2X�hf��ت��j�	�7�%���;��pw�`!B�ano�Өr,|�k�w��Ѳ�7[��0��x~�L���z���yl+�F��飘5��j}]O�Z��r��ݷ�u+o�=����$N�w6�x�J|�����Z�%pX����ூ�z����)"������[ۭs����G����Py���+�Φ#��C�W�.Z�c�����y�3yߴO�Æ(+�z`����qb�I�
J�B�!r��1�1��!rۘfRu�ezf�A��``�4
�Щ��(�)WV��Pݸ1MaV,H��e�YX$r���"ȍH,��Z�1*c�C�.Pm5�I�\�e���kQE���(�R�P��kZU�E�	Q�&ڈ��L� ��^f�+�%B�s�1 �i� �}�1����˳ư���x4\R
A@�g%!Z0+X:�4 VT�;�V:�Z�HhIP5�1��
Þx��ӭn0�N��bAd�+/i��t�Ʀ�
��H,5!KN��kT��Z!�u��<�o������Q��WXܥr�ND�s=���? (�2�d|	
AMy@Ă����܅H);���a�M'���4ʐR
y�&�H���	#�0�~����u�J���R
AMw����Xsz�Vp�P�*	ϼs��t� ��93��[s�)5�r!R�
ɦT���_O:�~��\�x�XjB���@ă�B�s̅t��{+=�����/p\�B�f�v�]9h� �2T�hI�*J�XS��P�&��7�3��̬�g��w�d�=r�S^+3�KP9C��#���3����d�ed���(�����물�X{}�T��P>7L0����I��+*u�d*ACI*]Si�a־uǚ��q��8���-5�r0�a�9@W�矹���^Ä��s@Ğ�T�Ë�B�%@�]ᤂ��[�� ���bAH/hu�d*AG�γ۫��N�{�4�Y���Fl�s�Ĝ�S�&��%H,.�B��
�P:�ɦVJ��ι��y��S��1�:�Y�k5���������L�HV�*AO/�� �r�R��N�H(i%@�bAa�{ץ�7�,*o�����a�AH,=���1 ��p�CR
AN{�w��\� ��5�d+�Jro��s8��'SI�
�R
y�4�H_|�{"�Xw|�T���
��ߔ�AH,�eO<�bΞ]�{O5s7X��{R�����%p֩�{v�G���*)Z��+�}�«��������!b�ѱ���^��;��˾.���GI��{W-�Z�l�0]4.�i���{F�qg�$�N�1۵��ێ��p�f������fu�;W�8�ڳ2��&Z����՘�E
���?uM� ��5�w�8���
�S5HV�k�^P14�S�y�����0���� ��uM0�
í����]kp� ����$�VM�y�w8a��!Y6ʁR�P�4�X����	)S��\P^=�������W�N�۫���y�19@����*o�!�� �μ����ޡXm�IP�yLd�+%ed���T�H���;5�f�9H,8����{�$��ϴ�)
�R
S�p$�e��!Y�o'Z�i}�v°���~�nq �[�Ȇ�
Aa���8�s}��?{1�9BI��,�R.  �5i�(�uHV��w�������tp�G��)�	�����?��"�����&� 8��}|�#�L� ����i
��޲ ������7鮃�z�2x2����I��/F�����bAa����∅�s��W��mW�Է��|�<�oM�ŕd6�r�͋�Y�j�jOg~j��<5�|�	> ֩�!Z��9� �Bw톙�J�P�|S<�{i����}x=kWZ����$�B�VVqa��e@�P8���\g�[΍���զ��bA�!Xy�:`Ty����l�	<�FC����9`^���=ݒLN{�;�I���Ad�<���<�MkY�R7C�I!m~�5HW�����u��]0*w�BH,�ߖf�*IP�y�4�X_9����֓Ɍ���Zݡ�ł�3V�ֽ���[�AH)���R��Ă��T�xi����=��S�h��HV�a���F�둷3`p����i4 T�����:�q')�P1 ��°�a��IP�*s�4�R'�sϼ��w5���ɉ�P1�q��5�^H,;��N�
B��S5HV�+X=�;�z�k}Tv~	}���M�ӫ�ˇ[������q�����$����
z�Xs~2 ���0�aN��#~4�\C��*q������ �r�ë�B�j2�T��L`hjAH[N��wz볓�
Aan� �W����������'( ���i&��|�w�~tN�x°����4¤�N���4ʐR
y�.��<o]�杕Ѭ�Mj�rA�%k�uU�?�|�~�ֳ^$]�z8������)��*AH)z� �AL��ƽ�Y�O3̅f�J�P�yM$���~�8��S���$�VN��[θ����Ă�P<���Ԃ�S�(�Rϼs��2��|w�㙰8@�TĂ�R
k�v�I ��;�������+� �������Y4��t@�{�u�f$_08��w�w����RZ��j�� �^P1 �hOs܅e.�ߤ�P2�4�������g#���;���D�[2�큛�5���O� ���G��ȇ<SI����ѽ�ָ�,9�*q�i%B�VV^2��8�ǻ�iiP.��I���,����H�BZ��A'�=߾�u�4��3��f�v1��[�,?|�/�W3�6����i ���q@ĂÆ��܅H)��o{�;�SI�L�7�&�HsǷ�Z�kg	�y
�R��w{�)�R�
�R�q�i4�R��'��B�4���ߋ��ӖaXq��չ�)5�P�Ad��<��+&�T����l�A`pԅ-;E!Xs{�T����́�r�����s݁Y�J�2T��j$�AaXV��P�4¤�T�=��9ɽ����s�G W0�bJz�W�����ë�B�5ih�LH/}p{�n	7��
Aa��!Y��R
}��i�aΞ7�Y��Z�.~�/i���d���[ݳ4��>F�S9�c9���_����>^����Vmg˒ڬ�u�YhVf�Q�F#�瓴��f�um���om![tP����)n�����lÜc7X���l�L��.W9�A6�ݭa�0�f4b��f��GJmE���ߟm�4~!��<憐�J�d��8�d*AH(��4���rsߔ�	<�ѪA���Cy�B��
���Y}�\� ��S�
�Y���I��)��H,+
���B��B���t�&�Y(��q���]s:M�q4�M�o����,ZÛ�B�����R���S�=��8��
Af�y�B�L�
��D9�H,;�.�5n� ����Ɂ��!R/�
ɡ� �o�cCR
B�w��ӦU�q�pJ_���o����K�J�`oc�_Ҽ��4�~=���NN�z���:�����Fl�g�++�n ��|�~�y|��Cj8�{_U����M�i��b#�C�m��緧x������!�p�3ܶ�\���N������#�O|���Lx���>Ш���\��gZh8�z>�ɕ�рn�֙��EI������@ d�(��fV��ħ�J
3��j��w7GH~��;��ϋ �s�N/���i�4���k3Y�V��V��σ��I��j#ԙp�#g1BA �%��Q�`�����LB�"���ad�W��PvЧVkQ�$�3���}��|�'�}�#������|�t^޴|�7g�sq�xÙ�H����J�D�`�yQd����ۻ#u��X��fͰ�"r�A�0Ѳ��� �T,��x��
�jB�M��膈�����"fy}�Ş]?v�n�B��lqQ�2�������ᷕ;B6:&��`ou���<ʂ��1�0�"I�_0Jɮ_�I:��~�檑�C�7�e���p	�LW��&nH������tt�Ǫy=��r���
(�*�;w۝�W�8���>>E}��dnkz�mAT�lI���if[�i>z���m��pcf���Ҩ0��Q���n��H�xٶ�`��l�r���~�Z��5>��W�$��� .�痽�Uz��'sW���/v��N9WDi�_3x��X��C�h�T��s� �n�fD#F���mW��!қ��� �[��ZX9���<Oڪ
O�6`�=���Zrlk�5�3�J�흚:m����  ��u�K�Xa绷���mp�{,Uoˇ
id�Z�Մ{Z�����2���;_^Ԏ��푷jP�S�p���l�m�����μ=��I-��4!3q2WR�{]������ye\��2g��q�.�^�[
��&�=��3v���.ケ.��#�k]���!�I�}i�p{�_:�QYQWof������7.�v�U�wdȰs����S��m�v��hU�O�6�CU��x�;�х�'E��yӖ�=*�Z����!���ХG4p�U��M��COE�kZhւ�pq^������e�;�Ⓤw�.���7�y��>��|u@�����IY ���H�Q@�T4�d[�iӦV��jLe@e�V
\�V���*0ӡ1P��mm3"�-J�T������ǽ"y��Y���ȩ��cU�`�����m�lU0�K��j�UMa\z3_�����a�4�3RǭnB���ͨR޲�n:ώ����c��;T�+�enm�Έ����>!}��gr�:�:1oQa-��l��깕{s����D�ۏB%��ݕ��&�x�ڀn]�=�gsCu��T�u�sVTЬM����u8�F阡��i�x��59���%���0�v���أ�q��;��]�&˺�R�K���tn�9����v�Lu�S�3bhҫilf�d�ia,is��lѷ�~kq���>�<��ⰭQ�m�pU�&�S".k7Pne�`WF�MUq����]n�����~��+��wYT�c���˞���nw<��87$Y���N�ٺ�]Q�1�<�1͐6̋�89@{[�+[Cj�d�L��L<�Np=#���]�F�Ef���0Y�V�U�m]16��f�T2���������#�UUUQPn,�<�ry�m�9�vc��^�(m�#�`�ؔ��4��b����7��|g�Ӽ0e����v���}�`�7cNP�n6���gL����@4GY�pۂa록���`�G����b�k��h�Z����6�x�9+��Z �En��k�C�y��#���D��	��L�7��?6��n�m�	�/�/�����`]���^G.��dd��+/���	�� ����y��Ï�\O��:x�O���u}F���	T����9W��.:r�/��oh������xYP���޳�{
���ƤU�F}~���I-@�I��H��QϚrȘ�m��񚍒)�Z*���/c`�P���_3���n6��q�R��V���=�Y1�ͱ�Ҫ�Ek8�������k�\O� A®8�['�߆���v�U��$r��B��� ��kB��)}��s��$�b���>��D��H�5I�N�L�G<b�5<7�h����9`3�V��!Fjg���u����]SL�Ve�f]�K�b1����cK���=K�j�۔ �g&Gb�aN��6N��j���`�wPevG�6���8ϡ�m 6c�KPi���I�K�<��D�UJe�u�Fj�|��y����}�W��͟�͑���	#��W�}ZIƘ ���6`�К�;�R��$�b�S;ʪ��jI2�u�i��4�oղ�����#^8���o ���ן6���<{���[�2=���hƗ������ܻ���$�۩�����QX5��)Н̒��s�\���|�9�#�d�>�u���v[��7��{,��8-ڦfל���*H�Ǯe�F�wf��=fl��w��ҽ<Kiq_���8~.�����9_U``��͗��HWĝ��q2��I��*}����(2��V,a�Y��b�Z��g/a���=9ǝ#qʨ�B���;�ֶ�6^�BI�L��euX�c4�hƗ��yP��羃wɁ�7a��ޢ�i�>�+�6�3�� wY?O�}�lݵ�%�__8�+e�7a��h~�T�#Յ놇��O����U�НW׊]�N�TW2�ߟ���b=Ik!�,H��\��Up�3��L�64�4��7�õd�1��a#n�m9��&c��$ӵ��	m��N�en�#�ugl��mN��YeB����Y���֌FT��1KZ˲�Q���7�(�����d9|��C�8_�y}��ϦĜO�z�}�T�'�� �`����<ձ­^�������WP��]���r��f�*Ωq+���Vy*� �H����8�p-�P��9��m~pOi <p��s��}�Y+XM�칋X�c0�j��b�8k���C���I�����?{*�}����9pR9J�H�K�:ֽ�x����]�U���f�ڨ`�����V�Z���ɥW��9�����������3)1�Ը�����$w&Gul&_kP�� � ��[J�	݊׽/�U^�]C Fv��L̩ؐE�x��E��GR��qV����� ��/�z�Ά�C>��$�_�R�D�ڍB�r d��Ç�S�ǭ�A��0A�u�j�r��bd�Z��9ԅ�GM�5G�'u��W��N�j��r�
���0��G�����Igz���nt{������s�+�d���������&�l>���nITNHge�_|��+����e�����h=Gi����_`=M��==xFy|��r�x�5�i(�s�F��"VW#\M5��ܒ�,�`mC#�ԝ/��A�6�'熅�B���L�մ1��s`�m��&�zLK��� ����޹4��p��~,�f�S����ȟđ��`���G�ܐ~��U޿L��x��Zh����{���2���R]�����?��B>�ķ$�'�M����(
�ÀU���*TU}�͏c�*���4�e�U�[-G+��u�j�+)�g;�|�-��)o�f�6$��	_z�E}�B��|e�* ���<���%�U�jżԬl)݃Z�B(��ުDlDvAX�A�	�b]�(�}��l�����H4����w��%�����[�8�٣d3<���u^Մ��E��{S��e�[��6*�i4F�թ\���s�L���:�7�!=���=�~����u[jt)�S���2:�x۷\�yi�ugf�f��� c����>�����6E��]�����q�X��i���r�A{Y��J�`�8CerK(���k==t<M�qb%���m$����~1�`�;w '�O�w6|Г�{�||�C����y�%��UQ� �G,,{�_���s�v��,��� �E��Bʆ�ܳVw�h"�$f�	sR�Чbwk�>�E6�;�0I��{+1�ܘ&�/z�:� �����V�R7c����^�s�Vv�6l���c���+3�˂q��h310A9�bi�=_M�͵�Q�g�T�^˷��v~}���,��T~F��gU����8�����jQ|��.՛O��}���)�rr2gd�͏u��ީ6��G3"��7��A��'3#���֋��u�Cʈհ�Vk�����R$�ݐ����u�}8RH�a�	+�P�Le��j�q&T��s�d�{m���pOy
�Ϲ}�̒_r�N9_J�ɹ����yQ��{�$;jez�P4�ڍ��p�Grdm�٢��^����W��u�b��S�:��\�}���,�g������P=a��ϻQ��|���s[�;�E�Z����꭪L��|���sɻ�+U,u����-	��C�d�S���n\46��ww��$����+X_J��p<-(�2���y]�#$t�
nm�a �˷H�yU+���rrT��������V��	�7j_Bj�|�~��<��<��]!��5���P��>X���}��r>ѕMx�~��Ս^�7�6뾮��z���<T�h�$�~Y�DÑ�}�J�{X:t����S��"�����i]�����\�b�ȇ�K��po�;�[��d���;��*��3V��Wc��$��+ߨ�(�+�)U��Z�K"��k=ֶ�B5ْ��J⭤�"9f����
9�E����U���WN�-��V��H�(V��F�h������0��w�iҚ�ŋ�t(T�1�E[Y�k7Z҃�QZҵQbv�ٶOD�q�)ǎ�S��!i�swb��b��k�(�cA���Tlq��@I���?�z�6��8ǟ������l&nǶ%ӝ��ٖK�l(���0��VCV^б��|~�O�N�da:�Y1Y�LP/����A8���ځ������z�M�<E�d�w�z�j�./�������.kz��K��H ݄�1��[�w[�lyC�5�U���P�e�lK^V�`�Z�k�a�<ɫ�7#���8��� ���犙~���M�R�t�|\ ����iP<wydB^�ߞ��*�ԇ���� ���a��n��~�2#zi���I;��+�tJ�&B�5�[�a(ЌE�W����7]�;ޤv�C+>�]y�I�j9iX�)؛�ܫ��My3�v��H�0!����5$s[��rA��|�93�wA�W#�dK�8zb�H;��{-�	=�2��~zbp�@�܀�܆�;_c��41�a�fd�{S;:�Q�=���e�T����!i��#�"�_�և"��ه��~������`L��^�.178B�J�e=ZܼWU'e���^z�v)�}�U5�<Vx�ۘ;n5Թ��u�ntLs]�̺3[S�AW-Wg%f汀��e��\ۛ�^aDЍy`�k�~���R�dus�����Y�#B_��/���]��-�gUJx�B�zT��s+�={`�����;����Ai�H�X���;���b|F���E#s�;É���!$b��<^�3���Mf\Z��5b��Љ�h69���fG3"��m��L5�52��
�:a�7���o�N<k��$o��{�/���k�yF8�����꫑��y=V��}&z������o{���&�qՠq��3n���].�ڭ.�jF�9{ $�ٗ��C�VIsw��j>�N����D�֙o6d¬t)���=wu�x���R���ts�F�M�d��g���[m���E/e��A�4�_3������Q�!7�@�|�L�\H�$�);sW#���' 3�v},{�33��X�"��18gު�xN��u�=�2�w&q��"��FV��n�����`ѡ�v�wzfJ��tը;����PV�HB%��7̿��� ]��y�����A�uJ����%R^; �܈����V��g'�ЧW��]�k+j�\�����o^\~�I�2Ɍ���9I�#)��s�G�m�z�'�:�@H�!Szo���0��.���H����fw0ڣ��b��"�o��=(��=�&��6�s5����a*�"n�JwS>�Un0�NW�$�$�� �=\hM�a�*ꂡ�ۻ�W�&cfG��q�NX媯7G��C�����9�y4T>#k(�R��r��`r`�ͯ@C�B�?��/�*TI�LE�م"�D�;�W��S���v�y��l���P��*ڻ�[s��N�v����=ɑ�����a�}��.{�Q�'a>���oi̄�5�q���
W��;��H$N`wnJ�hA��)�}�Un0�]s`����o�ܼ$ߗ�{͒��&t�%\-�������$�Ol�l=�}����T�qKY�K$8����D�D���,)!?8`���Ӯ���r��eK��i��ƀ5!��g��K\�]�G&�fe,�T,qqv�s��ɠ��v{<��*�����)�d���]� �a�%�+tw$h�A�%�LK�a���Bݒ��|-�`��K��:�Ƙ �0ĚU�B��;�v{�!���־P�b�K�b�m/�^Uw����#��"���r�}�:4)���A&���n�U['_��0Q�����@�&Iu�I�L���7�Z�b|g�C���(�Z�Z�~|�>�瞾����A9��w�U������D�QTF�3+��^�Q�c�K��p�6��ׯ�wQ��W[[8~v��$���|G�/����:��¯�$����!m�������1	;�C����u�oN�\��5�"9��#1�Ak���$��?�R)φ)�/k�CzX2�02г��=:�nV�4�$���Mu�JlR5USϿ~����kE����j��P�����ks�]j����{=փ$w?�h:F��fzTjd�G2��eC�]+�ٻK��3�ۺ�6'�%�nI߃�b=4���Y�߾w�/�H��#¯�$�e`�(u�������=��^�4
���q�9��Mu�9����;����W
�B0IJC!�i&1�8U����ɔ~q�yc� ����=�<D=�rצ'�u1���:��*�`f>Q��Vv(9�ʕ�S����^p���'��d��&H�k �H#���J��!̙0`�o[�9!T���ƻ��X��/�U�i�0*��wՓ������9͓�Y_���>�0.Ծ���gؘ �ou�	�Cu߫&�K�
����EF�&2�'e8�*L�<���e!�+�����7{ü��|s<��>
G.��<����_X=��#�}����m���'km�F�z��o8Uէd�e�	p�fv*;C��1���g38��N ��ɝ��f�t$U�;�`�C-nj��U̕=r�G6�9͉�V�M�ow4;���5��Ǉ��`�fݍ��1�	^C�Ǐ�z(�Fl4�I�u_*����f�csQ�Qλ�$`L����Fk��<�;/�_��q�'��>w�yX���p��k״�w�;^,�l^��{�!Wrq�%��±t�y�=�C6Q��b�&��wy9Tvkq��
��y7Ec�#x:��[���f�Qb�:Fv�-Rİ�t�I�[�>�Ayϻ�뒍>v�ww�b$+��U=��Uc]㗼TR��6�2�-��|3�z
���1c�fv�Q����svt��kdU�7�]��J��h����q�N�V��4&�v�n����׸-N�JY�@�쀳���H4������dႲ�_'�^�郚�����QaH��4u�d��U-�+ilPV�T]���J�孶1�YD��4PETs3i�4�:r܊"Z�eZ�26ҴN88��q��y���e 1܀��گ<s)���ܮ�*BE*:o��"�r�ȥU�k������b�P��j�b[n�`��jҲ�����L��rVTkF���U)m��z.�(1t��x���^K#��i�Y��.���
A�'������p��ρ�ηW�����:�̍b����W4rv��v�44K2�Xz�wR�t/[��G ��rk�Ӌ�8r��q��v�㜼����ۂx�v�+Qu#�y�58Е�d��5�d�Ύ}�o@��ɍ�\�ce.��G)[�ԓDfU���Hpb�x��tM�ak�R7k��-!el̕�d�3U��)���\��L�A3*K��]i46�l-��t��Gs��X-s6�f���+kR����y�'TC=;�F���2q���!�"�&��&��E�]������5���|`ݸ$�L�d�"G6���;���!<����c<�D�����K}$�Ⱥc])n.�e]��-#�mT�	�KT��ܽ.�9�
�-��>�'Q�f�-����ܬ�b�O�O�UUU�aջJ�E7c��Ι��l���e#q{��7n����c����t:�n� ��	"R�bY=@�nLl�P���5Df:�Y�<d��ݶ㇜���_e�����Z��D�K��ŎWGRb�h�u2�������6͘K�k�*��d��ҩ{B:�.*&�m�5�a��ڃ�)�~y�߿�ĝ��$]���}~�+�����L�o�(����7ɜ�� ���=͒G�����u�1�>�*Ȕ�re(ͬ{��˅V�p�rO&s�G1���d���vwT��& ��U+P�w\� ��m��RUtD	��k[?fl��}��g׃<�a$EHfXM��h�1=����K���2G�3��8��\�x�k�W�u�v1�u�-&�N*�'���3��D����#��w���W�~_��}�!�P9��0����W[gꮐ��랣M:�q��l�]��.\�I(�:��h�r.,˨y�6z��ٲa�+�*�T���s�B�c��̠�FfZ�w��!�ׇ,QjRi�X�c0�".EݫW(S�V�;�Ġ�b�]�k�{�u��p�l����E�*^�4�r�Or󲧁豠;�����a�b���L��"��áJe߱<�v��W�s{=b���s5QX�~�W��o~�s�1�QG:�p�v���,�s��E/	��)�$�9&gb(��)�/i�=�.��/c��-x��@�n���p60Ÿ0a�v��X"�g��<��U�>���w7񵡢�A>:��}֩Z;|�3�g�:=�F�fC��s���0��d.�,6��5S<�Ad���9 ��'c�����̗����]i�E�ك�a�*���Oh�k�@�۲�����FX�������|'��h�}�}�T?o~QG:��Uk���^m�q�&��v��g�U[����7��8xՓ����.�(���>�+��MD��'��|Q�o}U�gև,~18`�+�BJw��p��$=�2Ov�;���Q�dK�T�)�װ��5�Es>��^[b�re���y_��G�G_���K"y��͓r�������6l��D䊃��kҔ�ƍ<~#I ���o|�%ോ��O&�'�KSj{?d�'�g��F�|����!al�9�ܤ��75�miUy֍j�&�XV�Pv15t�e���a���R	��.,͂��4&&�4�m�d�jUU��L�%ಶ�6���d�)���Y�%�'��??(��������I������nvf͍�� ��}痡qJ�D��'������p�N���wm:�pE2O��#���_W{�|�}��6�u�V�N�/+�q��g�BA=ɒs�{R�ӴJfg��h�W#"���P�>1Ƒ�/��/����������_s�������;�L��D�7I���%,v_�I6m����t��|���4�=�똗.v��;��[�Y�3_�;�V��r���x5(D�6��L*�s=�����Koq�M>�	�)�ò��Y�]�U�a��ɒH6)��<��A?w0�ӨE!����^���	�^�L����=݊�>
׈�8%����nY�[cJ?X�?���Kމy⤁���$B}!�>��8baL�'O�ex��`�Rh��lȳ���h�+[D�]�""in�ԉ���`�4 ���Q»[�]��;C=qΥ`�ey�u��k����:.��?\ں�orv��5~��.��33�$����"��2�g�9��ɂ���1��(,�~%�ء\��Π�C>r�}��Y+ֆ�=�� �[��e+#4����"�>%��T4 ��|���lq������\�a���V�K���g��HA�*�E<A��R.$fۄu}��L���tΤo�[��b��������Ct6�
��س{X|�We��2v�V��,����"M50k��n(����}���y���k*)_��r�`���p9׋�ǷX��>E��\P�L���,H�b9$�_{�7!�_��ud��hg�"t����e+��]��]�^�D��Q���DT�n�^��l&����=��_�gn�]�yy���>��Ry�TN�{en���Y=ȡ�W�N����	Fvh\���Ҵ�}No#�6�~|�+��e���*����L��+Itt��X��ib�n�s�:ix�g�^1��nr�ʶ����		R+0��*A�d:�U@�TTC#�J��;��
��V��7&�6a�DM7�K��*)�tA��s�{��Fvve�	�gJ�<�����]�1�־m˫U�)�L8�������#���<���
�${�PF�	fS�e.�-�`����n��u.��j�mm��u[���|<�K��٫[�k
�iġR{pw5��BO1��{~�쯱
��{�̨����m�V�o0��y���k��wn�u�/�Yח�o7�e��|>��?n���Ϫ��Z������P��N_i��lgm���n��j�F�JzQ�-������v�Z����H����7��8�����߻:^R�$�J�#]t��m2�l�'�{����{i}�B_�ЧZ�j��K8�R���m⻴3כ/�t�_�QJ�@>_{��h���'}s�E9��pfV7��X͚���a%Q�;� y��U�!��R&�ޓ!�͆{^�X��;r�o,4珹�G�P�{}���u� B��%�q�B�q���O�b�ջ�/!�C��PT��c(�|.u.J~{���r6ӷ{Fڬv�x�{��`L��S�^�q�~^o��/�b&
��ʻ��7q�J#���g9F�L������w�ˍh��)K����_P�Eb]��qWl����W>�����C�sч���^w�ϲ�c����3-�ׂ�^�u�p��j�F��YT�M����d�d��r���&��r9��=w�wE��ioa���[I�U�X"ݽr�����.@��Q�㗄=�-�����9���G�ǎ��V�lk*�E�m�JQR���Ռ���Q�j��'�O3̧������W�<^�S��E^E��J�bR�v�`��֥KbV��J[���.d�0��@남^O��({
y����<�>x{\�y�E 
�x����'H���x��(�!��r�]!�v!J�Uc�b6Ķ��\��ee�[*U-P�pݣ����"�(�R�B��ͺX~w���.���p!�*�_��w�,���wܫ��ߣk/���]��P�f���e��*R!���&a)���-��($�a#}
>��_U�.���y!��g�`Qo��؉�@7�]�hZ�g,+4�Sf���*�_m�_}Q}�}�ǹ�]��U��}��4O[g���1]մH�S]0�Bg�Dڣ�_��ח���\�I���Sm�B~s��9�{=����K�B�T�Y����A�X�D#0�"�Ŷsþ���ݴ��Y�g\��ݾ��v׸x�7�+m��s�i�}��PQg��+پ���=<���;:�R��׻�=��u�3��{�QE��:��.m���˾���}zα��ʇ��s�Gѝ��mђ��o�7������y�Q�
O�b8x^p+ٮ��<X�M��=���o�X{s�&�@J�	Y��r�9�-�+K�� ��bz��gse��8��*!�GMM���UK��ñ��ͺ�n��ta��`M��I�����.C'U��h+��z�(�=_Ře�}�� �y�����}����Wf�o�������ȇ���5v|*�˼v�t��\@o/�q����}�(��>��3��&��3�2v�1B��`@���)�Ʌ���D�_�*)��{}wvk�������2u^V/�̓��S�q�C�<��9=v)�C{Ëb\ �����W��u�߲��s�2��k�������{����"��hl��mM7�}�O����uv�����E^�s��d̻�|���3KG���]~�I$���h�i�1."y���������G}�:�?�C;Ý���qw]�z�n��?�o����z��\�M���Kw��7.��^���hN��gl�tvnaĳۻ[q���[���{���X�Ѻ}��nh���/��^��{/��h�z���Gq�����a��n �B,��$)?�����0�\��&~;��(�\�Y�v��������_e��TJP�d^3w~��wJ[�Q�5���Q��|��L+Q�&q��uf�[��d�̦��Wٙ���~�=U��p�m�gef�᳚��z{H���쯶�5�l��{�xT��6��N#b�Ρ�W��-�F7��i�岪G��h�9�)Z{�?}�}�
�y�S��@NV=7MV�5V1��+�_Z�叭��<�R�K��`�>A�7wk��n9�D�}a��)pُ:{�;�}�Ԇ/_�RU�`NM�6��Bn;�2�2J������!W��fg��c]\�7��7����\��Y��mPb��cO�lt��. S0Zڻb���A&a�4XW&0�\�7']����]9V�m2��a7hfU�JU�In��A՛��ZJ�b��0�:�MPj��7J�n�F ��c!Zh<�6�Ω�#L0�1���g��5�~�+0�����F���k/p��9�!y{�A隊j�<��@dt�B알��1���u>|�5��̙k?g��^{N%�C�ϸ�7�D���ds�m��D{th�@�	F��JL�"m��9���*C=Wnyn����<�{�X�cC-�����}�?q����ӹ��=�^𷏖�����k���VK�C�8}x��v�sDS���2y�y��}5v/M�S\�άv���{١$�c��ey�V�|���u����]���~�w��Q*�s�3F�`� �8��V�����7|��޼uqI���7��r��A��汯6�t,2����?��-��A%^5�=�&A��r���E;ť�1�Kp
c�=��orL���^���E;�Хxǵ�j����Fzm]|:/�2^�������>ݪ�q��=B�A ����l��a��"ӉB����%2x?S���2r���z��q�8/6�|��ۼ�nc��¿\PM�^}|��O���og<n�踫U��c�|/Y��S�)����YtӰ:��C;0(��K���r;y�����DSЍ>^�L)���_^�������@��AD�b7p��d�����S^��i}�{a�zR���C�%:o$��eV��;�ᇸ���<�?!懻�v���S�Wշ�7����)}T�sw�g��r���o���r�z���;��	�lS�VnL���>�&�g9c��U$��O؜�8�8n�D��I�x!�8`5ݶy�Pݡܭun���1S��q`u�3f/Gk�.�3�o��"�%��Vv�4��b�vs��'g�G��Wi���o"��9�,IQ�жNN��yT�ǹ�:vݮc��RJO3��M�gF�6x([>�l�9�w���zS�v�2l;H�Y��2�X�Ӛ*N��k�=݊t�o��(�j��F^>������Z�Vnu�:�>����n��೽4�t�v���F:U��Ƣ���Q�U9��6u�*��<-e��[�����;x�+ٮ�)f]�wX��;�s��BT^��1y������`�x��a�uZy���9�W$�rPP�]T���bYD6B��Hs%DJZ(����*30��Q#E(�Ѫ6�-fKnL�Yt�E��L\*�������GF)�8^)T�QV��0�)AjR�k[%�B��ңJV�TT^'�Lzy�M����E�r�r�c*R�ݪ#�b��Y@��yϒ�뀔8��+ܝ[���F�2�s���IY11e���b�l�d(��E�H!��ar�mU��R���\nP(�d*֚CI���Ve�V*�jc�f#R���Y+*�[M!�#4���
�P�ԊE[KI�	V�
�5���?!�RZ֤��t*�%՜�Fr�ݥ��W"�x��sx;g�.�رsdS:�0R���e5.��#6����1hMm�a-�
�0���̱j��U�q!-���8�ly3$��㗯I�����*��:�������M{3�f�]tN�Zƚ�Feʗk�d�䭣.�#�f��af�5�mn�L[	bE�{.j͌vZ��.�3�QN����]ny�L9�۞�}p!�{u�ń��1�����!���U���c��Hl*\�d�c��m�)46f�M�7 �X��p+nک��c+4GP��X,�q��l��t��{�<���4Cډ��XT0�.M���tk���hf�L��Dx��P*:�uhK/-����I�۟B��;��s�͞l��r暠�鮉k^�*��l���L���isUUUU2�f �ڷYwZ�j�z�ư8H۴�LX\fȘ���,-���-x53�\�XĦٶl�7J�r�+"�Ԥ+"s��5�K+�8�s ��;�+v�I$ӕr9�smGK4��av�5⎋�Hjl�%��14Q6{hT����2q�2��*4��68\���՞��y�v0	��S��"PI��G��+D>��;V.��_���+����/�y�@O*�b�|o�Z�AJ%0u'�+�üW��C������s�_+��c�ۊA۵��w�2mX�{���S��K�	$��!dȢsQ�DΉZ����ߓ��?<�?�V��}�K�A�"����GaMJ��Y�Y�7F��[�Y���ḛݧg�1Cݩ޿r�`�˩�^�ϻ�}h��Op�:[��T9D��ۻ7;���n_�t-׏�q�v�6]�F�=l	{�Kn������F[�n�`;e�<���r�����_n�~��[�^Ҩh����^܃������/����ެ����~��耝�6���{�๺�,W�:t��v���C�U�u׶OXY$���_{Pᓭۮ�=�^b�Д��_f�b�)�,���F�e מuwh
 �e�퓔�!;�b'8:3�1cv�`��m�9ۚ|�[���ΰ�a�>��T�Wն��Xp�m!��t��:�E�u9}Ә�~�����q�za��Ļ�X}e�^*�PhBd�v��߯w��,�t�E�Sk�7�/b����Ԍo�	ˏ��|���;�����{�)S.R�����6��X��Q��R)�7TΫ����1n�t7���x�;��;AKQ�v����Ծ���w�һ���mR�u;��_{<���;Ln��
A�{�VR�u�n�����>��h\��[�}t%ĳh4����1�.9mW�z��6t���
C4�2f�ˋ�Dں�gcK�S�NWZ;r�ĺ9��ɣ����!��� �	�h�&�&�:���eF��)f�`fv+�P�#IqVsb��66Ƭ�B�ð��-o�OI�S/�����n�~�C8�{Cf�Ŗ�Ԯ��"�?n
�y�Ŀ����7+ԟ��o}�L����@��S�Um����ᴻ����ou�QxB���̋�iP�}���o:�}P���yc�<�iV�*��k�_~{��<����b��,9���jx�]�*���{��N�/{O�"�OF��eќ�k:�gv�î�٬����Ow�R/�������!�6�����J{�w��U���w[��n`��W;�V��~_{i��v�Ā;�`���sP�{�t����y߯zmN�1�8�LfB��]�g����7���ݒ��w�B�2�/)�ؒ޵zy�R��=~"Y�9����vI�ߦme�뾳��|�{��Ȏ&�t�j4X��3�l���^بZ�u��u�������4�ܸ{Q�v,�c>�����Y�D�J���.��X�0�-�*UU������ݿ���uwoOo���{���}#��c[��j���n*ƥ�|�x(_�4�ވ	7����u����>�,������zj���W�=��P�~��8�z:8�=�v����������0�}�w�U�$�ԽU�X��>C��{|e������ұqI#(��0E4�A���ϗ��d|�:=C7��)���_j���W�v��_�uffK��&��������?�]5hLRVe�
a�{ރ�����2Գ�֤2Z��D�����A���պ��\<�:'v�3?E�[���a~N���z�G�T3��z� ��rJ��~mF�"HUe���F[Vh�,D�5��hXu�$]V�j	+c�4Т)��T��9���#�����}2�.�������vx��0�3�gkNW�i�K� hdc&ԯh#-k�d4RKi���~�ओ'��3��������������5�Lܮ'��T���&��~�.��u�����ϵ�j��}]�w�W�)��C:�[��Ǹ�^m�=�&����(|��e!X�ʐ%F\YU��-�����חsJ�{���T���3.���:����n����R�H���-t++l䆞��\�z�ۋ��}N�,��/7� �ڋ��\��q�}:N�)��wj��Z�)��zGe�~�C;i��q����k[�qm��]"���/P��Ζ:_n���PI���vhV�Z�G>��w�y��I�_z��܀��p��zy��7���ԅ淡��]wA��l'$��/��_��Zz+�������[2�*�x������q{�zs`�-:�u�B{��R���*2���LOq���^��=����7Q|2|��?[N2Ȟ������P���i�t{��t�=�koN�T�r����$�e��^�y�f��Z���ףN������U,�cΜ����J�))p"�*.�3�W|�s���7s8{�7�8Ӭџ3hlTx^��O[.{�I�w��}����?����|���VQIf���9̦lB:�%;7UTW��7�n�cpn3;�M,��ь{���蔑�w%i��Pý.-70�md�w���,�̜lmWh�n�UwJ��5�������wԛ֙3�J��j���j�v�ʽ2��ZM���Lp� �O,pk��1*����
�#6���R)�B�Y��eKYP��	��cl+U��V9J��
�q����,��
�2�H��%Hm���K
,�Sl��J��E&�4�2�J�Q���Tc��X�4��IPm�e�
E!�A�"�Q`,QE�AkP�X,�\ea�J���mP��dU�V-j
9f��2�LEj��,RV����*�R�R
�"AH,��T�����h,��T�u�[[�5�"|�l��K����w���ި��]lNY*mb��y���<�@�Mv���m6ep����F�Q�8����<���^Y��Lv`�(Ga�S�����X�_U��g�'o�u(=�]w�us�qٕh�&j�ޭ~��l.�H��������.nt�Q��X��KԳ}���>�������s��|����m���6�}m��J�j�-؂�p�0��qe矔Q�}�1�Ϭyzz�����}���{'�i^߽K�#��s�;|���%��l����@fzj��B�u���W}����l�7�{�kȧ$�RT��@�'!�����.�.�y����a�{�G��5��Л�Z}�m�gD�K�Nh���:�Y��84�i�[�5�(՚4%	���غ<�].�i����r�YN36N���<8�2Q�C2m�7;J�l��Y��a�QYZV�]Y�[M�9\e*=����S���jQК�Z�@����T�~���}�G��W��1�}��NV;Kx���o34KT%]}T�u���V��q3�*y ��B{Ⱦ����W
+Ev���ns�� w��43��3�_=}��rm��2s�CɭĞx2ʈ7"i��M��`%b1.U��<�
�|}�'Ϛ>������k^��s/�'�/���to&^�J3Ь]�onN����;{ӑ����������g�9a�q�9U���2�����or�'T�:x�P_�}�^{W�ʇ��l�+!F�!����uֵ���r��Gќ>��?����5Fo�Cu�k���JOݫ�gп�<�K����x�Ϸ��e9'K��{��;Vb����7+i��)�r�$ۥ��>��3�������]s�_��<Mf������o��b]�(��v ǨM��xw@spp~�s�=^���en��_����$��~Ot��{�܋�4s�nrCJo���2��/� +���Á$$@z�ϙuӘd�Ҩ���@Vc��i���rM�)}:�a$� �&�j����߭
7��>^,��ыs�\ro�i&����ARTl4���}#�gV��[V������8��6l�f�j˪�F�dkH��n�u��~_7�f�F6%\�)�J)n%����T��A�>?{�˭�uᑰI���S�7by��⊸����d{98�ډ�k-7�}K�_�vg��������e�%���ެ$��f�9���+�`���u8�3�}`�.N�M�Eb`�I�n����zY^�In:jb��{w���^p�6f���/nuɹ�?��l����9fFv�^�򍫷n��u���Vi���D�:�m�f[2��ԄX��4e�L��$!.g��v�9�,e������┭Ķ��9q[S:�uh-E7��}K)uafA�l�CDJUUG����Q�h���$�/�{/b���I�µ:��T�֘y������h�Ɓ?U/�4��F�M\���xAt��C����u���Ɠ2�%3̵G�(�tA�Nr��_Z]B��^�-�.�>��D��E�&swi��}��6��)"��"�P�.5=��<�E��&)�`
�E�	�3jw[nC���%G.͛,�Ėgl�
��;z)�4�ْ]�&�d��/��9�ޝ�;f��`�y���-^�H�?u�/!�a�wf�9�28�d0Q�S]����UP���u�w�d��|��_�LM��Z���=H;��]R_j*�G*�4��rN�vUF��7
��&�̼�%�	����|�PW���
(h�b!d��F�������S`��ğ����I�A����9^�^�9v�,����|�ϛ��=��L����,���k�ֻ�{��L�[dhOF�5����W���D�'!��bhG7a�@�M��q��6�*&Ux�4������GȻ��&	�{L�_Y�a�0%�(R@�qc��`Zc>y}�k���<�=H���Z�Ϯ�nIVs�1���ϖdX�!��mR�g1a�K<�OD��*mJk��&I�3YxE�"�wuU�- ����0� �%�og�uBE�۰�����(�+Zf����^���S��Pߚm:�ۑU���N�>�
�>�O���n{uV�ߗ��1 ���c^p놔Q�-�aae�]����U����d���Ƙ����4MZ�Y]Y���;�nc�B܅�{;qh�0�#�0F��ӵ���Y�(���@J�Ǯ���/&��H�Aյ�G&L����0��4#1�/�S�%2�U�"nVv����g&��:PU8��~���!���S�j(�U_��!&4��� B�B��$�!'���#8��`P�8ɜ߃P,4��>�G�o�^	�v�La��63Fo�Z��� ,XB;-��⅄��9H_�C��P����+ n���a��҆2I BO�H�'�'o�����G��������B��8�f��ІO�"��F�r�u�4���=0�)I�w��'?8P���;�h9� ��������g�����`H�r������$BO�������_�ο"�?�	����?����_����~Sa���?��������r��<�>�""����?��a$6}��M	f���!�Cd�QM�����[�đ�?Q�!���a������'2?����Y$�!"t},�$�yp�c�5�����@�� @��#$���R{%�P�|�p07�ӮM��@�zO��>� ��)8��b������	���|���І�q�g�gd�}�L>��ߤ�g������x?����<����)���� !&�Y�>��$>G�C�H}���������'�|�����C����Ϸ�8�? ���96�C���?�|�>$�������O��d�@��@hȃ���?QC���>6N��a�`���P<����B��C_(!	L� ����O�'`���'�ش��`��D��N�@N�����C��H�� }8�,I�0~�H����� ����,�' $��}aě_�g�|�Ì�I@@���By�D�I8�Y�`$Ė��r�h�`/��A� �$�`~��?�=$>��I$H���	?�	$C�?��D�����?�>>g��'�}P��>�|�`H~_�>�>R?�~�C�}�?W���?&�Ą���C_��|C�k�?�Y$�!'�~S翤��0���� ����:��$�@��O��������� �>a�`~_��}>'�	�ȇ�����<Ї0d�~T��Cc�P�O������?/ϳ����C���/���Ӭ�$��>f�Z��ĒH�>ߴ��C�k�?_��~�60�O��Q>��>_0�G����)�����6CP
ě$?a���B�#$�&O��}D;BC�I����w����BO�O��	�N	��!�}Ԝ��u�?n@���8��Ab �>�'����>O~s�����)�z��