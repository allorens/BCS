BZh91AY&SY�����y߀`q���"� ����bL>�           =��F�tr�vt]ݮ����	��9)˕k��iݢm@���6v�7m���F:�N�wP��3�v��7n�N�Ww]��[c�Q�.�F���+��ݻM�i����$�J�
��l����D�h��ka�	�bi6d֦X�ͨ�XQ�ڭ�QR[j�ʫf�Ҥ6��]U)�ģCw$�['G%u���x��RYU��j�0j5\�U֢-ip������%��nڇ��0��X�L��n�IM����Z%)��v+�-�[6-�UjͪK��^̶�UCl�< 4IPr}�#UqM1�̀˺�6� ε���^�ݻ��خ��ˍUں��Vų���̻j4�]��u������cM�!�[[b%T� T�T�E.���x0�AIn���JR��K��U���r �[{G����V��(t��\�T�){�'�iK�y�{i�$V=N���jm�[ihf:�   �ye��J�:���C���S�x�������@=[��*y��"B�K�G�{Q���<�Ҩu��wK�4�{ogn�=�&�
�fl31�5�(-�  �g����Yy�<��j���m}��)C�V�`RS�X���
*�zy�D� <o�˦�RU=�<�T%JW������@kƻ�z]�Ӻ4�;��:Qe�f�RU8�   8��O��i�������.+�yW��J�n���Сz����2u^甪���s��W�};�}M
�+��*�Wg�,��4���Q[�;m�m�U(j�i�Z��m�  �A�N�]�tۻm�h��>�OB��G���l��GRJP.�W��U��w��>�u�ڧA�4ێ�*�Q�]�� :�/p�j-�J�j�i`ж揀 �| h�6�\��
ܬ� �w@7p����.�� h;W{�{�4�6� ls�����@���Ե�cCj�U4�P�6��  �� i�4(��}�� �X ����F��;��7W/{�� =�`((wq�z
 ��G �@{�����ƖOc��4��Χ�  �[����`@O.�]�s(i�4V7m��v�7`:ws��
q� �Os@ ���w��%)�+[f�KZ�D�d�  ��o���o� �;���}� w`nP��à q����ִ������X .�^= 4�     ��   ��2�*�#  CLL ��ъR��� �� '����(      ��	*��h�    j{H*����)�6��� A	SPz��M����d�d��6���	�>����������g��˷~?|ί��:wZy��d{������ w�9��WЪ ���*�*�{���3 �
���?���!��_����� ��:�����
��>��d� ��������d�&0����d�d�'8��2q��<`�9���O8��N2q��1�<d̜e�'8��^0q���d��0񇌼l��2x�q���`�'�2q���a�!�30���2q���`��<`�8��N0񓌜c3�0f񓌞2q��a�9���x��0q���d�㇌���d�8��N2x�ɘx��N0q���`�8�1�2q���a�8��N6g�<d񓌜d�'8��3<d��<`�8��^0f0q��N2q���`�8���d�'x��2q���73x��2q���l��8���'8��0q��<a�La�'8��N2q���d�/<x�̜a�x��N2q�a�&a�x��2q���<a�'x�q��̜d�/x��^2��8Øx���N12`��8��x��N0f�<d�<d�'��'8��s`�'��`�8��0q��񉓌`�'8���̜`�n0q��N0q���d�'��3'x�8��N0q�2q�����`�8��0q���l�8��8��0q���d�<fe�"*<`� �2�A8���2�x§�(<dLP8��*q�N2#�QxʧT��N0��|aG���0�x�L�'E�
�0#�Ax¯Q� <`������OT� <a��N0�Px�/0�2+�Px��*�d��q�N2��Ba���^0��Dxȏ� <eN2�0��Px�U��`�*q�OS�"�@2#�D0q�0#1�Dx�/Q�"�dG�"�2�@x��0��|d���0��E8A�*2`2�x§A�<a��0#�aW���C�"�� a� 2�ELȩ�2�q�0��T�� �A� �aW���^2#���L*�^0 q�C���^2 f8ȯ@<`P�Q��`��<`W��^2�q�^0��|a� ��^2�DxȯU� �dG���8�$E� � 'Q�*�G2��U�  8ʁ�Ex�3 8ʯ��eC�x��x��0񇌼a�x����N0�<d��8���'1�/L��N2q���`��ə8��0q��d�'8�8��0񃌜d�<a��N0f2q���`�'8�ǎ	��<`�'8��0q��Lq��d�'8��N0�2q��d�8��0�2q���猜`�'x�񗌜e���2q��<d�'8�`�8��N2q���`�'8��a�'x��N0q���`�'�Ø8��N0q����>2�<a�x���x��N2�0�<d�x��1�I��<d�8��N2x�`�<d�x��񇌙�g�����oA��i��?��$5_����g�]��e�$*�h*��X��+�C���Zڒ��vZ�7r��ɻb<�E�ˑ�� ���2�I�Vs Z-Zj�G��4����$(�M�gor҄�4�m�Х����x�rƻ��y���_^_4QI#ۻD�����h�ُ�I2�X� �%\����]�eT�$n�5�N����dF7v#���Gsp�)k�0��Z%��:4Ԁ��H��5��:�kfUd�ֶvz�Y�ێ�ͼW�
��j����#x»W?Sʄ�9�b�T��:XR�b�mǩ1P8v���	�b-�� ��=aZ\�՜��є��������0��)�Ur�V�ޙ�J(���jBSǎ�
�N�m�<�ё1�Vnڶ=�������/p��*�X�S0�ƚͷ"�x��-;�H^���z!85^i6m�Tˌ�Ș��\���c��ΌӓY�b�U����.Y�%��QUj���v79n���,�=��kF��#ү���K��R�*��X�NMux"�,��2�ȅ�E47v�r�V��Z7�ZA^��օ0o�X��Զ:���cZ���4ֶ��Vɹb�[�x��Ө��{�����z�����D�W�V,a��-F�@��n�L5t�]�chS^N�C&[��yB��z�
"ͬ˒�[�B�!�v���e����2;բ�uFuB�i̾��w�`���`��+�U��KB�V�"a�s���]�iR�%#�ƴ������^����� �`��r��T���.f)U�y+.�������x����m�Y̆֓�%�sa�ْ�CZ�V�n�t�������4Q;�cuF��
�S{��_�sׄ�ĴX�lf|Aմ��[G��u�ʬ!�G[��+���.������L#oM�\!)�L9iQ���\����@�H�pk*�\�gal�ôҌ��ؙ�P�^yY�cK���,�60.fm�[�v��-r�t��j�6��F��=����AaK�tyȅ�b��6�&:��`8/'�W�.؆bє�-Z�,p���CXI�-u'GJ�a�tyf������ݘ4T�(ʄ���V2¨���>���2�<ǔ0T�IY�uyy���Cc�ܳ/#�Z��j��7��.�!�����i+s%;��2��H�x�O��Y�iM�a��Vn�3UV]��rBhS��,,m�Tَm��P�U�uX�.T3Hb�A;���k3)m.���p�^��|U4�n��t��ȷG�%G]%��J�!�;f��Q�U��t���X��or� �R6(^�-�$7r��������b�ӤӺ5R�^��x���S#ą+�r���C%�;Xw��n�eީ+Y)�$�԰��x�JQ��nV#0��eG��1F�
؇sv虁�:�]���{U$��!�#��u��Xh�TS�c#���&!M���Z��͊[�N�N��oNٔ#�;"����W���sp�e9N����c�(:u!t�
�O��ڷi�L�rܱ�Ի�b��c4J+5j��	d���"��Dk�,�s��%�zr��$�ˤui��u{jL�l]:�WX�M����V��[�,j[ޡuh������Oy��ū���8��hRk0�"��	�:+�"�kZ��J*ܲ�����]�L6������of�Xu#r�'�L��B���Zjy�M����q�e�܆��<gi�E
��r�a���רs���n
sq�8�[�f�,ۑKݡWI���j��"�=���M���Nݽ�@Y�Ӧ�ux��Kzp�vH�m1w�i�1f����[b�[�%�S%N�|���ܯ��M�_;p�?�O�q�m��a��k�˧t��bt��\��������&@�����Ѫ-qJ�Mlo2ۨ'&��8��E��T�gy��NW'����	r9%M��>V]��L�����d�2^�Ae�e�z�*,jJ��	�]���f�1�y�B�[Mqfa>8��5���@�h�S��7�6�aͫ(�dRG��Tl/��ʼ�z���Fܙ[ �Q�8LGp F]�m":���'[)[C)Dì��t�l����Dni3��7��������L��BK�O��D�\P��3}5�)9���t��f'�ҭ�lU��1��$!��]�,��"��*�ҧV�����Z����ݼ^�ʼp�*n���7/JY`�\�u$����Xf���2r�m����񠵣��AE��۩�ZP
K6׀!0�@�*��Y� ���c�Il�^P9�m�� Ӫɘ���J�w�e��w�u�{/i�j�G T-4�M�@�$�[�TZښqC��䡐���n?
�P	څ/E�1�x�jQ���B�&�ܦ)ª�R��a�n�KZ;Sq�tKɴ��Άv-M�f��Y���NT��-S;���e^Y�iܭ.��#�mvͻ�-a�t*��SwqL,G�rii-��!SJ�$9�e�@c�"��e�Q;���=2Ӧ�7W�g�M�*��+sP��£%�Epf�3Jʕm��hU��5j�I�{�+ٔ"�0���ڄ�EflnEYfh,�W�sH�[�Hn�yVD�Y�eǠ��xs����lj�r����V��y��9+'��ُ+%�j��*b�H�D������=��\;3��S�{E�7��P�(@��!�m�BZ2ee��Z�L����6�t�Bރ�J¯NчDt�V�bc^���SN\�w4i��iVovC���[b!��5ѵs^>W�6Yn:�%i��Qۘ�!{��)R���,��[�Y��ȯFCx�ed!#tY�m���O��+�MP��M\�wb�m����AL�z�/*�[m�4��faX٪س`�aT/d˼��m���D}�3�����y��%c���󪌽�֦�[Aںݳ#%�\�7M�Q]ɐ��Ǟ��
'F������e�V$�Tr8��wsL�ڡj^��K�T[�2eWeIM�+x]����T+J��N%��H�F�$��ov�[�R�3*d9t5�@w �ͬwYqA��f�YUl�
�
�d�꭛��K��f�h�t}qq9b-�M��ݖ�Hգʛ���wJ�[�^v�U.�*N
>ֶ��|��M��7_n X�aY�g���q�m�5/��o.��!���A�)�U����)<���ǰh-Ne�,�S��wu��׹6�ID��&:��M^��懊�i�����zh���@��������!�8͂wu!��\���Ł\���� �YxZb�1�E�E�(��A=��ٛ�)��&������'X[���se���z��M�K'U�[6D�&�S�Ч��%B��W<VV�K,Ǡ�1ǧ�u�+n�+.K�M,���#��-��Z��Ĵ��nő/a�s%�I�t\��P�Dh�(Ż�%�Y5���<e�7�S��`�ZA�ĈQ�s#�)h
'��s(#+e���M�Q�NM�"�+�hq�n�iǩ5*�f%��l2ָ�8��{r&^�̖Ј�W�]M\ݒiy�I�r��X�f�k�lo��V#&1f������qEu*�9�J�c<މ�,��b9_.x��h���Uʲ����;���`̝A7.�i��1�*�[�R׹�۬F�c!)]<ܛ�o�[��t�o<{�=�>N�+�tF�(�\�V�Z���S��s]�6�Z+
��Ғ�B��>�dǺ�hmJґ$In��7�&� 4V�<����c{7R�@Jv��wS6n5ö��8ن�kb��Xh��ܢ�Ӡ�S�M-��1��!oFԱ��2PvDd-,�2ؓ!�R�۫�j�l�H�Ct�'�x�AH,β�)�oQ�liwXH��36�/5۹)C����oke5[Qգ�͢����xV7
�E��VwP� �f�?l�H�=7��]�/*y�w�����t
$���D����H���K[�M��ŉ3r�ԩ�u#)�a=�Z�c��S�%WRMhH֞b�y�oun[w����E*w�!�½q��j�#�ʹ��O��,t�7�P;l�Ѵ�;{{�
YWH�����{vS� ۫����q�Z�kSW�ZgK�72�XT��L�Ut��P/iK^=@��V-�!��_1GY��'���їR5*���Lí�u�����Wټ9��_XN�}Ŧt99�Z��M��2�c�b�/���-kP6�N��ŗ[-��;�7��ͺ�P�$�F�T��J�ӧ�x�[��nl&� ��cI��(�u��X8�&h8pV˻�$��:�^n�k�rY{o.\�5�������Vۍ��,�{��V�^��qm�Ռ��u�y ��N��Փ0V��W��,0�yن�GfUصr���k��Cj�wR�s���uN ��Ď�8����������{CJ�f�pu&֎7�S`s�ov��� �� ��f^�x��f���8��C4.���ۮ�nP�ہdQK(;�FYguj���k�����p�	�;;o6��x�QڴR�t5k.�|ӛ{Ճ��j���`s	9���wdUP{��צo��y������bշJ\˔ܽ5��n�9�֐�6�ݧ�д)��ds���K�g5Љ��E6�dDC�F݈4���N��Uw���X���3a�TN
4&��x.���\"�i��0 ��u��,ͮ�z�ٵz�q�nȻ=�ս�Ŧ�7)��-���Rzw����f�S�׈PكC�n1�]��� p�{��="�n��U$�z-�fF�J�܄��oa��ov�������f-mu�bQc�5��ǰW��P��@���-9;�������8]+˹bM��xMv��]��E��2�Zֹ{$WdC�M�j� ,�r�
W%��Ֆ��3ejnꈯ��,�Ѹ\�ˉi���ˆbA��2���u���<��=2�re� r�+�<gv튱�y�s�E��0�ѕW1z6�Gi�1,,�Tua6�Ɂ]\�b�Z�S��ݓϞn���/s����4-*�YuH��I�X%VH&"Mqj�p-������ay�e�T���Ä+R��Y	��g6�̴�\���oc���Y8Xj��Ena5ڛAjVPIw�V*����̚��'\�IЫ&�V���DX����1�{����yW։Omt�.��o2���o�.��p�����O^sb�[Z+Lie�r򔬿<EG7l˕���|l�+868�t3��]G�7��̽r$X��.�L����+4���e=�S`�fe����++U�7+�̶w8I��;�Q���+5�X�ڵb��v���T�k�N[���D`������'���tr�5N�ɶ��SF3W❼�d��%�3H`����m��cF�\�S��ʷR��Z��KmS͑�iq�����nq���M"Fv��Sn���7�Ry��&\쮬�1Nܧ�^��rx�������� ����:�aT&��B�#nF��Y�z^"l�3^^< �T�5"���K&�WY�t���;�^)��ʻ@��/�DR�{P�3V3x�g,��.���o����CLэk��75Z6uln{
���ˉ���!P=��(-~o&9�n��rSXi��;�yZ���!��5���-J�R�۰fM��]M{[��Sɂ���[wSLPѸ�"�zӶش�h�l�w��*�	�ǫdج��`�*#v�����85{�6��k"�:�q֭5�m���=�0$�r쨭�9r�cq� ��壯+v�1��-�i
JSp��r��s��2��NP�#U�,i����v�A֎�[���9�zm�-�6��G�+I�V��Z��N����`ᣘ2�f��U$zVn9@��7Z1�9U6���&�j�,}}n��������"0ʺm�i����34�NѨ��v�X]���&�8ix�ߨf�GtXt,��Q{I��m���+<�|��K�h�d�W���?�*tu��ㄇf]����]�rY(�.�r�0���6ɠoX�öYQx���C;���2M�k�P���'��z�5BT�^�v�����l�8D"����B�F ȓy`�@i��0�B�v\-�8��5����Vi���U�:���W�YgD[��D���Y��A��P!���&�=��xmlfѸ��[��L�=XqZ�d٠��� �M��*�K��n�k�\�K�
N�����5RB�HQ��$8�7)��
�頉k�N_�
?Js�����%Cws��ʆ����S(�6�ِS��m�F�m��9��Pw��up��%T	�ha�#�Խj�Z@�	(�B���<��0e.i%��>@��|��q�5.hQ�v��e�B�R�3�Vrp(_j��%Ԝ�,x����J���ݰ��Ĝy���qh�/��aF6I�@/8C{�X)2��ͧ���8�5 �':��a[b;J�v ɵ!��귶��+���|�U�d�ujW���6�@�є�f�;4�9�cz-�W6��y��݀�a�d2�]]�PSȭ��"ȤQ+A�L�V[e�
��f�8|v�]iV.|j:��z1�Ѷ�k�.U}���z��֎�d��[�Om�p�i������	�y��\�
�B��WTMy�<˳	�7��d�s]���K]vXn�`��u�iq��Q\�0�Сv���'��G���š��^��{ooa�7"1�B˧Ci:k�MȽ*n�ܳ�i�B�v��]2F6^Y�V�ŵ�_��*�՝g,�:��h�ª�_]Ni[�k�Fa�4�>���7/8�Uh����8(�gT�D�Uθ2D�3]�e���$8�}�;b�"-��Յ�MQ4�١T��������11!�j� �꼝�m�P˽�i|��>ёV;�}%�kI�w&6^v�eC;�2a&��|*��5�i(�2���$~�j�|[�� ��[�>���3��~j��6ͤ�C��L�sX.T:�Z=db��@���Z��Q���-�U��[L&C��n�W�k��bx�d��Q��Av��s�R�9u���Ҩ� ��OYV;S�qNNt��,�5�8����i��D
'y�2Ŷ��j�17E���vN'��H*��t;m+�AfVj�{���"' ����k8p\�M���$��ɼ�1v=i��X�;<d���K���bu�vMKtw`�*.�j��V�:w?�yU�~��f�I�F'�~8/]��z���ɺ)�O�G'�Nv9k�@��ʮt�WH6�7u�-ȐzBr��L���l�-@s��w���_+Hu����s��'i�)G�E�hn-���pA��p�[��R:�3��&����&	�kR^���Z:u�n�Sdh�6N6�Nm�R����ڽX8����8sp��ar��|G	��ڒ	������r,�c�gm�
$&��Cj��yZ��`jfn
��{|v�C"'͑8��(>B0-ݒW]D�r'ڤVpLaZȝ<�J7t���=w[Һ�s��3prG7t��H��F�c��od��bާL�Ĕ�X� f�摋M�*�4�a��.6�Ɍ�O�����kܫ@>B��K�)�A�Xfٵ{]��tZ�}A�f��e]�S�v�f�\poҍ⅞Bֻc�[ �&��d��E�J�C��_E��w�բMf�'��J��/��8�u�8�m�ɩlˏ�f]<��F�������4'ϪPޒ,���IZ3:E�/.��\'%]��P2˽�s&i��3V�V��44��>%I���H�\��tˠ�ܜp�gʴ�"f���8E#d7��<뭅����F#[Ω&��,^5
	Yoz��H�e24G�������D1E�r�ֳ��C$	
�ȸ�t�ۉ�?��0V��S��v)��1T��Fi���#��*68�F��o\9�*j��U����0��U����3�!�]6�S7��MfU�������ͯ�ދ2�(��W�q�Mfߐ�CÜ���y`C��ج��''mgY�DG�ՙu/n�^fJ�M�	��y@���������#�u�3��*�U�9ٮ�z�P�)\̲`�16������Z7�s�5*NTw�b�yWԨr����5"L40�^���^�!����ֻ6�N�ӵ��8qfϤ��)�������Q�=K`�'<�H5Q�xz���Y�j���K�ej��V=�T���7��T�>|�.������fs����G7~�yD�7��nR���㉹�5"N�oN���Z�m��r˺�z���������\֣��/nr��ͻ�g[�qt�D]�{|ڹ�p�ɥ�v���50��r�,}�hAF�-�(ov��|��{���peT��
Cz�R���n��8\?
=X�^���A�"m˲�m���ͱo��'}�wd�ʢ�M=��L.�$ԫ!rȵX��I4>nd�-gef���K;&���Z��|id��,c[��1�7ۚ��2�d���-��y|�d&�iT$
�`��t������l�[Y�!��×�A�u
����[WP3�b���nS9
Q�}��u���{ ������lÛMt�J#w�eFfYWj�[1���Rok�X�� /�*�~F��n����L<�i��;�gۮ��O`�m
t���Q�j��6�nI�"����	�y=Վ�����hI�"]���B͓�(��>�Օ��h�e�H*�2`�ܻ�c�u�M<��X�d�Vq#b���6:���1�6j�Ú���XD�U����6�d����=��L��ҽI\��Z�i�U�vwi'۴����Y�,�R=R�[y+%��4�4�릃 �F֓r�l�����ۮ�!������UbV�^�s�#Ǌ���ݎ�S�T%���PP�NT����LIW,�!�&�ilSŰD�Tw6v�R&b�%��A"�{�|�iԥ���2!|�yD�tw��5a�;����3�����<�RE7s�b�tw�L��be�9�A-�ڍ���%V�Bi}e��"C+K\�p�Z�����l\;3/�D7w{D�f9�s@ڇ�l�i���d��TB{Ǐk6�X��W#��W��z�d:Vب��]q�A��GIҵ�r�v�XKs�)��� ��b�8���E��558�u7�K��nj���`U�m\c�1Ӄ{M86k�ib��i��wo_���DD�̸q���U�9W݄��&�l!lK�çG���\�o����y���JԒS#B�\�늣=GZѓ��2�+	����dSǉőèsu�^�؝z���p�0�q��q�:+�ki�卧8!��>��V���0�ows�������p�ʅ˗YB΀�A�I�T#NEr��ބ9��+Չ�\�
���wڶ�ҋ�u���d���H�]	v^c��٬�R��_��xq���.q�3��)��4F����+%�W>�aa!u*oh�VL��M������p��͒~��N},K��틺���JzM�֪�X��7�c �#$��b5d���':����cB�jtG�xǡ't9�*�e'9�nu��V�QN�(X�݊�f
dǷ��� �t��`f�<]l��.?waY���U�X�)ޕ��%���S�2�'�Yp�&��M9��᳴��Z���h'��ht�xwc������YC+n�ܕ� VS����꼆|�a�;/2g;)�ٙ[�G9�t��(�N:��ln�ADE�H�B<��G+#q��Z�S�@I�9ڌmu��9�@V4�9Wq-݆���fٝ���>M̼�-�vX�����S�ݍskF"�U�m��@a�ZD�s��٭@�\c�w�U�7#�{��g�:eX&Me����\��E�D��!������oZA��M7�3�R��u��ͼ.��yuC�-�%{+J�M���)Gw�x4�J�p�H�B��C��e��$-$�2�g1���O���b�t�kwY��\N���=�[T�mJ�h.*o;zC�}F��aY�ۣ(����>Sǽ�N��)Ij4r��7w-��r��M�k��7#�`.�Y9C"E+�]H:��6�uH-.�U��W��#}��A�)���s��2���K+�\n.�+����,b�!81�9{lRE,�,vJ��9#ט:�hH��!5��4N���bG@ɵ�
�wu���#��]J��б�Q�0]���hk���ꋸ<65:T�QXL��O�e-�q�(,���<�����t"ݽ63�<�j�G����o��Z�)M�,�u�v^atkz��5�t;�2e-�oI�[��������%�(�*;�Cvs�V�u��ZR�э}�M�ݍ����NΎއx�g;[(�j��}�1��R��׮�c���Ջ&�Ρ؊���^�Y-_=�.��̮+����4�k�syZ,@�]���m6��4]�r�wLn;Y��ƍd��GQ�h���\T���>�/9�D*����GN�FyRWW��O5�֯��[+O7�>��/w���8���Pе=4{��wƭu��;�s��S7Ͷ}�v�!j��B��kAb9�У�IӗwS�)l�p�W��_�=��
x�ocNj�6�-� �f�d��o#�(��i��+�ǸMG6G+T89�cs�Н����IY���ݪ��ou%��6�˳i�"�R-���9�M��D,�H̘��S��t:�a8^h&��#���j�����ۂB��g�Km�k�Ǝ�ZS���kbBEҺ	-o-廷����f)��8U���i�3�-����+��Y4V�m�{+t	��r8q����YX����󵽌R�9���Wf�]�ӯB���<�Euo|���.ľ��d�7W,�m�ٓj�,*qyA�U`��*�����7�#�b�|��+��g,t��-=��`�HLX��oK�ݣ���N?b��[����u�������l���(^�˫{)k4er�橀V,�N�6���e���άskj&�T�>�}��Rڀ��14��K3�H�U�92tиe>�=�%;O)�r�%�X���k���=����u����u����lc�[u)�ʾ�(�l�Z�׺�s�Ȁ�Z�H��3rEF��kM[T��=;��n9��$r��6�i��Z����ݝ1+;	��x�ZOnSla�ѯ�b�	v�͛@��/v&%N�H��W*�&�v�E�\���d�� *�j.��b���>
�B��:��W�0�g4j1�fHr�MA,p���SU㧔�M(�Mok���(J�M�WDò3����!A�v~g��%Õ�07����W-�7HF��<ʙ0Z|����g�4,B��a�{f�s(�yR��A	�@��z������A�V�M\��e�.��poF��v�#
��-��c���خ}�ʴD�u-��o%A>��4���h�Z�r)��L�{k�1�!��r��
|��51���ќD�� ���ÑT�iफy�e�f�<�N�q��J�-��fڷ.̎����6��%&����+�����Cr��1��ʕ8-�FUTƁR8�9y3�T$�ɺ�]��u1H"�m&��0�^����V�o�\��
�iv�%�q�`2&�.wnNҝ�H�I��n�.<ݞ��s��ނ+�=2���]ț.�fR���3*�絩�����xNAwi�"]}�n�r=u�foLt�5�m����cQ�u���}�l��ŭ�kU��KV3��O5ӣ�{3J��:�o\t27YB����Sd梀]h�j��t������vSaQz�x�ږ
>�[�:AO6�mFuE�]w\�:��2>����}���؏8+����C��;�u>u��O۽V��W���νZ�A��ai�-S��6ڣH�|75k��L����7�$��-<�իBS����n){���/��p���1�'����}�Yx$2m�Mo06�E���;.-7��q�*�����{R������$2ٛԩ�[�)����y�!�0Ҹ+�1���GI����vV��;������o[�u6��.����;�;���=T�g��{Xzyl��{R1p��FwkXҜF_v!8J���`�i���2�N:��r�j�؈�����	fT��{M,������p�,_�+���J�oi�.��z�M/���]	�Wx��](X�q�]�f�5W�e:k	�U�����|.��0�֝e�8�3�S*V�qC{Cv�_ZP���6�'S���8��1�l&�+�`Y�U����GK��Zf6�n��x��*Z�b��* {����j�u;�To(N��ھ�os�����l[��{yِ[�G��\z�	�)�B@Օ�(�>�Y���{c&�7�<њ�mf�3Av7n�u&�Vr�Z1�9+
S��n{���0�G��r����ܭ�I�8����^�V��u�p�ф���[��*�6T��V� r=*T����lSV�]�aL=��<�7k0c�[�5�=��bf���.�ZTA��L�=�6��ƙq#��P捆�����FN���;T�)�jٝ�.܉
������Fib$�֪b��bgl��*h�m�O�Em��Ww6S�b�\�M��L�8��ۮ�yɸ��q�n,5-�b�-qR�車�j�0���3��3^����/4�cQN�}+�?�����u�Nf�YX�\�6��[�<�_�X�h�5s����4�k�9��*��0v@��Ν���Y��'ꀼ���%JJ#d���Ŷ�Ywi��G2�_K�7 �0�՗��/��ԟ5��#j���˨��T�:�����k]�iwmLy5̵�T���[S�S�vmZUXx� ���� xU����n��p\�1oF�C`��o���D6�bܲt֣�o-}�/�:�HM�9sp��]?��_d�oA:Ĩ��9ǩj��#i$���d�S�͍d�FZ�/nEY%4��yI�� |�A6�Ψ����
 �4}K���X�x��m!:f@7>R��u�H�RrF�I�����m�r��u��`!���SO`�vP�T��+����4:�kA��q�SUHEm���N�Eu�u�)߬X&�P'����V�/%5�(��@��
��J$�Ci&�zˆ��32���� H}ilC�4���8a�\D((��wEQ(XQT僴�7S�P�������U��)J�'�鵢�ߍK�I������ԡ6���#�tT� ��i�M�T��_�IBN�pZ�ܨ�Io�� 	B� 5\j�"h���h^�0ؖ�#-YAX>;�*�<3�J��Aj�D\��)GjCe�ݨC�	 :�&�x(d��#�.�v��f�:��=�~�>y�/`�u�I�i�����?�s,U��&h2��h�)�ۮ��'q��ШQ(�$m
E�E(ʫOb"���2�j���(h)RM����*�� n|�Y�-tuM�dPM�	��,��%c�F�����ȑ*����
l������g�r�:��B�h��Bt"u�%YH&/�q����W��F�I���p�#�"�o.�l����C��r�RP��@}H�Gd�����P���".�4C.F�H�"l�#���	�r�Mܷ��~��{�{�#��?��GDQC��������O���?���y{�?����}_o�?�~�Щ��i��
�}�f�W��U�h�v���q�X5o6�150{�:�j<5�Kۊ[�k��	q�{K�*�no8q˹at�.b�t�=���"�B�tnM���vkh�a XM�A��\�.4���VV^ؗNfo.�k��;�Úh��Ä�U���n'���4��˨2���ʢ6�9���p5���a�x��NN�GO�}�����fY9�a��[V�([T���OE��sLLv����+�q��ݛ��Mw���=�;k%�?8�Kڌh��gD����rᖲ>��������������� ��7n���,]= �V������
�Gsi���dgo�d�L"�a��(6�cĵ���k\3^f^�O�b���Jֺ�&��er���d��L���+U�LY��Qo
C��n[C{"u0r;q�nb�Ue��Wn� �zt��w-��wZv�(p���+�
�Dǵ̱-].������KMe�/�y��f�h�5�Yn�SP��3Ө-H-����(��T&��v�"`亁�؉g]�n�1^�;�g����h��$��w���$�:]d��	�X&�t��X$30G.�/�p�V�w��;��������V^iX����Fd*������}�z���g�^�z��ׯY�ׯ^�z�z���ׯ^�z�z��׏^��sǯ^�z�z���z��ׯ_�G�^�z��ׯ^�^�z�����}>�O�z����׮z��ׯ^��^�z��ׯǯ\��ׯ^=z�������z��ׯ^�z���z��ׯ^�^�ׯ^�z�����ǯ^�z����ׯ�z��}�޵y4^��� �x9�	�Lt�f�:���n{#�8;�v2w��\9)�XX�V٣��)X��\�N3W���6P-Ve��ְ1�I&�/pV*v�5�X��>�T"��= @3�l�k����Ǡݼ{ҵ�)��eb'���[-�G�����*��%��^:�NnV֝ G4qvF�����7��{��g��9��/c�N���#`]੫����6oL'��8�p�Pi��72
���8&��3:��
��t��[Ԧ�vR��'���nP铛�(,�m�����vs��|�<�NȬ�u�7&咭,�f����Mɬ(�m%��q�Fs�gK-��(!p]�-��?jĻ�3��Kv�S..� lGL-��d/�w�֚��^�(G���܇��y����[�y �p.ݮ�E�B���ؒ��Y���ɝk&1J`�\�E�kB�����U�{������;&�5Vd��ĻY�74Y�y��G�Q՚b{t�+�.�q��ݎ���[43v�pI5BkY�X0�e�̌����z�Nвt�,ů��:�;sg�[ୱC1T�rċ�e YyH�|����Rk��MjfI��!f�����nqvܸ�N�{����k��[=/��1p�UUj��}>������ׯ_�z������ׯ^�z��ףׯ^�z�����=z��ׯ_o^�|z���ǯ^�z�����=z���ׯ_�_�^�=z���}��O��_o^�|z��ׯ�z����׮z��ׯ^��^�z����ׯ_�z���ׯ^�}�z�^�z��ׯףׯ\��ׯ^�~^�z����ׯ_�z���|�ww��k���;��+z�#�RSs���.[�/U����wñm[Jd]2�w�%�K��GC�eɛo�ɑ�U�.�/4���j �3��<b�4��B]r��a��	�IYz������J�x"ƮS\��F��0�f�4:�>�OG�#o�MM�e�w��ѹ7�d�(�ړ)Ԗ:����̽�à�)��A9Ҳ㲛�nu��������?͌*Y�3TIB�qc �\jҬ��u����D+�����S�� ʽ�ZS��nÑ␉�0+yh��p���}.����p�K��f<��;���v�o!��-I�����Ȯwk�nå��o*&V�ռ(���j)O-�(�; �u0�v"��:�kf��I�3{��s'pU��
x5K9���!��xv�k6��%a�e�t��@�+�-�
�nՔ޼#�0�-;,d����|�6�CTݖN\�� u��5�l�/���C�w�+���Z��(�!�enwVF��b��Ȼ��7.!�Y&м����&�ty%��:����}-0/��̤p�a�Ej%���n%[*,�`���
��ky|���������N�zs�����^�z��ׯ^�}=z��^�z����׬��ׯ^�z�z=z��ׯ^�~�g�^�z����ׯ�z����ׯ^�z��ׯ_O_c���}���z�����z��ׯ��^�=z��ׯ��^�x��=z��ׯ^�z�^�z����ׯ^=z���ׯ^�z�z���ǯ^�z����=z��ׯ^�z�O����}�^YRέ˖������ĸ#���ivȗ6o�ܚ';��b�3-*;D(R�����v�;r5��|�j�_e�'�
9���t&�X��~��fL�i�L!.��%nma?�8!�c�^�}�F�6Eӆ�]_7a0_	�\��\���mM���kj��h�;��7,�j��F��Ӷ��K�3d��L�G��xY��X@11���ꀻ�:I�쾻w���Q�A.),�NU�'���GE��U��1 6i��C�-��n������뫙��Z���(�fP�1֊7}��3)�s�S�'�۩��QT��*;�ʶ��{���iY�����0j�x��(�\���欷��w,�MiPb5ue���΁r��auN�0�Թ�	Wr��bMa��GI4���ɜ�B{�5,S��h�����[1�����ʾ�zlu\�6�P6�����KhTLO�	��2��]�y�;=f������bx���^��{ "��L��Օ{|��6���˸�m�Z��*�N�� EX��*t�u��`ۋyX��ͮc���P����k���:�oe��.N��Eͽ�&�Ԓ2m�����6nr.�:x��eo=`e��R�X�z�zWBa2�+J�&Cf�t}��LeDk3.���X�O_����~�z��ׯ��^�=x��ׯ����^���z���ׯ^�}�z�^�z��ׯףׯ^�z�����=z��ׯ^��sׯ^�z���}���}�޽z���z��ׯ^�z�z�^�z����ׯ_�z���ׯ^�}��z��ׯ��^�=z��ׯ��^�x��ׯ^���z��ׯ^��O�����}�J�}>�>�'8vYwxn �VYh;cz(�}*������>{�Wf�]]��~w/�?^�̳���CϦ
P�|9�%�S�9��U�E	�a����u�>4�[��������wdv��h'.�${0��*�R��b���{�y��@f��U�ؑ{G���������<�Φ�!�1��1�e����NpI�X�gZ������	�}c]	��͈þ�5T�*c�|��I����ݏ�T����_U�Y+�`u�!��d�^�Bs��N��^�l����X.��^���s��{v/�vʌg�C[D�:���I�_��Ƈ�$ XA&w��U�R+Ei�g,V����-L�WT��_AO�p7�L2qm��*�=��5L��%v�	8@�����tO7[ڻx���V�+��#2��0�V+ۓ�lo 	�?=��v~��ɠ�5Q�8�v4�}���aZxw=1+K�� vj��}�Z�l���7���X2]ۭ\iM���7@e:%9� �U�CD�Х8�ln_i��"ݫ!GU,s̺=F�0t���C#�C���e����sO��N���j��l��D{�u�}��a4�3�?�ū��o�b����H����Y=+�`�����/Zp`�j)��`(m�]�)��`A�F�y`�� +B<^2���� w��pwR���4�f������e�����y��]�cu��-T�܌��ʽ�V���}E5�&1̡4B��2�frq����J�k�gl�ddyuh�|CyU���[��؂`�e9��PW��Z���O�	}#���-,5r[�?W+A��XH*�0����*2��7[���;���	;��FX�j�1�K�*�t�LS�}ه�
��]�Y.��y��,��2ۮ������{�Z���nM]1u�;�\�orkE��G��\u>邋�_tT��d���������btw\�q�:��Θ Y�[�}%�QLin�,<\/EW�_&d��7���T���i$��ڙ�BQ���q>�����LHJWb�U��O�瞭����3�u�����v�;�Z���UT��0>���j��Y�+1Mf/�_#�r�iO�t��i�s6W5Ϙ��ϥ��s'.��-��ﾶ�\�LR�*�v�v���]�n���H��1n+;`���U�L/���\�����[�{���n��:�+h$�h蔮%	nJ�lnٝ�9(�ƀ��SV��JT
�q);�U��{�}��uf�䨊<)��CVɺ�r�t�]�;a���������b�C�0�q�uCv��o��M
��D��.�z��I�	t�>\��X�W7�� k[�&����띟�/�ec��-�Jn5Wzd|�9�*�^1Ɍ���BəeG�(''@P1��9�G������j<��"Z��]@(e�^�g+��{ڭ�d�N��c�&������wod9���u�.�EK.%���P�X[Dw}�k%e�}������Sl#Kn�Y�&o6���u/�.�Չ���#KN,P��v���cP�J�[4���*�6n�.]�����,,�/{ ڔ�c�x˽���r�U���hA˷���J5�Q��\��*���Q�66��۬s�gSM���{���8N��D�	E�l���Uik*�:gؑ�V��X�%���V/����*7\㆔�kw�)LKr�.۴�k�-�ړ3��Ar���"p��K���&_&���v�{��75�'n���'-=�Zw�Æ�-�&���Yʵ888)�i޵C13���t(�ѥ��Gz+M�d�Ә ��>�hi"���&�*=��`C�W�W�<����%�dn6��p�战��������#dS��������̳��јn�6@x:��y
���Q��v'rf����A���)�+ATS�p����)��=T��K&��A�y��9B>;n]D)�0#Vn��⩎ɖw�r ���1Y�7`��<l����@4=T;�tƢ2��yE�^����1�l��x�x�9-Z�ϸ�*3��g�����Rܐ�b�e�B�Z/��K���6�R�X$�:rb�o2Y�A��ڃ97Ŧ���������n�ݥ ��+w�"P�Nʣ�=���������9�`�aż.K�Y�t�742���8���*谮1�����6��]2�+�.�s��s�W�w}�dp�G0��Z����fƳ��i��t̓+�S���O�쥬l��%9wq�+#�,{r���`=�}�&�M>щ�9	��-a�t���Ea�͒*cBN�B���wCd�Q�3��ӳi�,�p��;j���>��ȆU�ɕ��z}(�c|5�[@�Yy��/�}~Mq��A]����/*��d�j{���N����{)��e^��-q�уze}yh/���f�V�)������%9�j��V��͐��}8t��.��Ti���B�1:��I�V��˩'*]ڊ�iN�͙d^d�'A;�5�[cr���Z���C҉�B���
Gۙ��׸oxs.�XЅ�@RF�]à�X,V�s���[a�w�Z�:Tg���l=]t6�:��ܑ�f��� �*ép2:3*��3�����\�:�]��]���� m���/�Lܴ,T[H�P�=
>p_��K�VaL%�`�@��r�����˺�Y�,p{J��z�W��/��i�t4���b�R�dŷA�0�� ��Jf��y�w����3A�=�ЛJ��bv�C�`������Y��e`͢&4�8c�d+���k�f�4�
൦i�����KN%*я%�8���^nl$WL���8
.4�+&�ۮ��i2��XL���Ard�]�9� X����l<�+u��3n���&c�7��zw9q^��E�U�2��\� ʮ�d�f�)����'궫0�F��ȣP87kC������mZ��32|2�l�s��̨r�þ��GZVR$M
w	�!�7f@F��%������I�,�/�s/���Cr�%�I�9dq����y��a�A�~Ƥ�B�S�T��û�2)��j�~��&�^"�vr�r����r������!����H�7��8�brs��k39:�b2�YG.i��M� ����:N����W}H�jي�H\�֣��y�iR�׸�-4u�	z!����
��Nc�-Ǭ!�y�!��B����1�k���I@n��$(�1���FV��9����9��S�٪�U������~�.��ԙ�H�G��Z�0Z<��]+����>NV���Mu�w/Q�N�h��cp�]q�1�+^�9�®s|ź,�(�78AmZO�gn����p)�F���1���	�����*렧+�XO"��'�U�>��]�-�+n@�u3��k�D���KN�A(�/��p�s(ԑ��9o��)�%P$o�%5��Uz2�H�Q�-��u<d7غ��
Z2��'u�m�Wz/F���n�j��
��bHp;��w�*�4��콐���D�)�r�uJV3k+����֊�"��_&4,t#��c���y X�� ŉ�N��݈��&&�ԸI�e�����H�vu,7nR���� Ҷk��[�e
�QN�ܝ���i8IǏkw��ؕ�╝�X�b�4۫?M,K�2��=o�gJ���>�[9s�`�	:x�[���M�T�v��!�����݂0L�P�.��X�p�yc|��qn�b������m�c�m��W�"�)�� ��S�!ף5ܡ3���
	]+�ў�Fw�	7.BA�P�u��0t�P��b��el�Nw�#�i]L�wa�{�թ+M�A@�ܡ��s���Ǧm�u�a�p��)�)��ϻ�?���_}��~��_�����>����߰������>��=��Q�����{XQ���0"Ia���jI�犚F�襷�}��SF�@9>ܕ��y��|�����7Nl��ݙh�r�YMh�&��]�VK��r��ȴ�;�q�
F�Ҷ�mŧd��X{k�*�;��g9L�\}nK]RC6��"���G��؍��c�{H=Nm�fl"�������
�P[�omC�#�F����GX�4��W�!�{�4�����J�5�mY�f���0�@�sI��Z˧y�*V��f��[�M酗@��R�n�)��F����%Y����e�s�O_kɸ���\4�m2�bA�Ǩ���4�r,��.l����92��`]v5X�ip����U:��#nپU�k��tu�w���Ux�o'�+ "�
�D!�_S�w�[��Wxm�(�K���l}D�m�i"�,�Sa��n�-�ja=��4r�&@�=�w+ª���:Gg\Ǵe��!�q�|���N��q��n���Dr��۪�
���xc���뤣$��|/C�f�T_.��ՇePdh��	��٦Y�ݧp����bG�����^���N.���D!����X1�Ǫ�_R蝇�I���	�.h���[�U,�N�u��6lIS��ūE:=�3Zw1�w�rT�U��kQ�|n��N9$�,�SPw[��D��":Qb4n�0�DIn�U�p-�.����ͪ�����1�Nѫ���ʼ#^��Bn���y縪�[1���mf�-j�h��'m�Z��h�r4�������~������������b(��ᶶ�Lf3��ڵb6�F֣��o-^lmb��Z4`��|z�������~?����~����N��U�m�Uk!�(6�[����V��<2�V���Vg=z�z�z�~?��������B�}�^Z��FьgO��~؎F����2x�ѣ�o5�y9�M��$p�C��o�Hm1�v�<�#��<||>�o�����~?�����?��Wc	VΚcF߼�����/ ��(�j�4�<����i�_{4�7����6|�,��]	�T��'I^H'g�n�E�Tӫ�y�����J�y��x�Q���Z5^P�ًN<��̃��m�= 4n�R"9	�i��%�8ۄ"cH��H�m��xD�mG�Xxo+��h|��DS�+��<��o������$�#��p`�A6��$�B4'�ȇ��i�<�'! ���6�^iڪ�#�MpCiˊP:hA" �Eph�c� �4�y�o�k�3�*<�[��ESULyo#QD���y����A�y�f��u�Q�f(�����5�DU�Y�;�/=y��2��E�#Z14h�(��;��4���/������=r��׼1ޔ�%s,;�7��18�Ϳ,�3�u�*U��3�]��T��M��ӑ�Zؑp�9�c��)�?/��Ӝ1 �o�;��(^xt�=p-�^�'��X��s�ؽ�g�zM�׳���1Ҽ&�y�l��O�|*����;�bRW1=��M[��.t�ʐ�1�&=ZX�������w׺�T�
�>��}�x>�!'�c�����[;���"������G}��\I�+��|�ϩ���o��Ma� ��z柪��:}	 |=���WopD$��q��/[O��7q�|vN�Y"�����`\wz���$�,Qf�2����� �7;>��ޞyc��\m�o�g�W�y���9q
�}9�}�5A���ds�	΁\y�{�y��t�;��;�?2��׹��j��7�J���c(	7L>@w9�1�+�$��ic �Ӆ�m�g������Y��l銏���;FG��ѽa^�}럫p�WC9�"o���R�㓞��j��`�ׂ�'�:��㘄���6�,cs�����ku����m"v��ҝ�1��_]��h$�,33+0E[+K�I��I��:�����V�kMkϓ]Aa�(�\R����j�{�j���n�!�{G��>WWKʂ�.����5��9Ps~�D`��]/�������l��y�p�"��Ӭ+�a��y~���}����K��W3%��Rx,f��~ۜ���9R'���Y�a$(�{W�e��\�:֥L�{�o�T��Ww��(�j�ezk������c�z���|Yg/��{þ�~򘪊c��y�Sxy}��s�6������� ��w:�����Փ�+
�Ԩ�� (2���\*N�G@�a��3��䌪�9<i����
"�G�ԯ��G̎T�2��2�ۇ��U�90o�����:j�J[��Eo�^�oηAp���o�<vH:⯎}�Q�N���޾Q����6vvAʺ&�[��oUǬE(Z��w��\��ܞ�^�����گ{���wڏޑ�Z��b飾6.hU7��+�[IҖx���<T{�����c��{\��\����p;ɨԢ�el�n�{���Q���ꅝ~����n:����h�R���y]��^�1�4�u��֙��aX�ٽU[a���>3���s(q�����H�A�O{z�׾�=��GzK�o*���!G�*ݿzR����3��ld�䧟h��[��~s`��g>�hx<���:����H;��o�Q�h�W�P�گ��5��u��3s0V�"`;{t�{�wd�MlV�6��i��"������#�2kL��۰�q��JVgwd���0�(��f�V���]�x��a�D 8{���|�o_^edڛw�+���iǳ��Ves��T���@��!䰥�\��(<�u$�kۗV��ߗ�m9*.Ϲt��*�L��FW@u�+fo��9�]Jto�J�7��N��;����u+���B�`~�㽳|FS[����7��'[�$:w��L����w������Qe�emա�*���]q^?V�䧣u���Tb}�p��Y�+��i��h��v�6;{_mT23Ըc�1�ŗ.�tAR��=�F�a�.������A�.�o������G#�Fc�t�;�%.�o��i����fY�+�6��w���b�|��Cw��ʱU�' �ܕrZ�gͺ�A�����xeޘ,��/̚4�3�����3�U�w~/żo�^<:��ս��z��s�Z����\;�`iV��$�v��=��G��y��\��X7�E�rMwv��Ț/�O��mw�r����X��Ԑ����m9C|�A��P�MG��}��W#�ڨZJ�Ьٜ��ݠ��3�3S7݌g���+f�}�ռ^s<��gPkT��w&��󙛓[��#O�2���}�����0}�R�Ozv�n�rh������u=NF|����-bګc�G�OVd��{g���2ν��H�O��/W�'�Tǟw�⚻�U~�k�<���3��S�^�sY<|6B��etwt��H��S��YFRv����Y6V�sǗݳ�fy���}��L/?r�2�X$�5���Н�"�l�	(��Q�VU>�T�wJz���N�����L��[�`����{���d�@%ƭ�]Y*X�<�y&��v=��ԊitaQ8��L|��C:�m\8f�喂r�F:�gJO��x���ܨ�ۗ���(~�K�~��ALɷ����a9��̮�(A r�C�TT��<�/z�_.����՞���\ �4��·["��d9�k��7ƨq�;��8q���2/�	cuf{>�Ǯ��S�P]���X�B�{���
E%{�^`x���{<�Sp�5k�X_�q^_>�_{>7*X��u��Y��O�=4=߆}��/�t���z� b򇧮���k;�i6�߽����FW��uCM���^9�(��&�w��1���{�3I��u��<s��Ky=5֕�����z槹��|������j����|���<5�{���pYD����1°ڎ5�9���Y��Fdt��gކ{��q������ökJ�׽���j�?_��0�\�D~$Q����UD*�-�ۮ��|��9��r��.����޳�-C��*��g8� طo=�$��ε�c7�f�5�(�Ou�t��J��P"�<�
Z��+ř�mNo�5���X��\r,X�<��o���^}�yj�7b�[��+��,�|�V䉥�9����W�M�tf�};c������9 T#��\sy��V<�3o����8����g�M�Ri�7��rC���Z�n��~
2�'�Ϗ�{G���{��z�eԁ�q)����w��y�*MǗJ��|d͎Ny�o������KN�7Wc��&u��m����Cec��6D�Qx9��|�;Z^��#"%�X���8��q�
�3�V����u���}�{��*][��a�]��<�Fs�g�^�쿹u�}un���5�������Ά�����X�}U�Ʃ���Bf�??�]t� �F}�J����ެ��L2]� O�@;���_¥�^�ze�x�m�Ǫ�A� �����P�3�y�V^����i=�+u�u ���p]��U�'y�z(F�XGp��ff7�K4�o�w�y*��	
�����Jޟ��p����#���d
�o�����O0o��pf5ߦ�t¾���������ǻ��ʙ|N��4�d�����i^�A�Ƿ��;���7�^�0.�Zh,a'(W`���HO`���]w3�I�Ǫ�����<�z:���X�ڷV��:��� �k�E�jZ��v�6.ٯ�ț�i������@bɤyM+l?�������ky*����j1+����o���k���}��{)6�����ǽd�m}�6�45U]�}�T��~��f$�$����ӗCܛ��o�~��̫Ѿ���}p}����M��� n���S�E��[N�m�9>����K�w{W�*M��/�.z���d��V�I���{��'`���#2}DV��r}�����mOs�骼�(^z�Z���B�������۫�إ�D�o���zr?��7���{O�l��� ����D�Х])�����z���u��pM�}_������y]��{�=M�3����9͟$8W�7�4l+��2�������Ϸ����� S��3�j��|�P�~T�"x��+L�������\�g<~�kkj��\k��}x����;�y_`]D}�ù��Q�����Ʌ����pZ��ц��"����Ae�%�Y�O��;�Y����7�F�@��o�����Ո�7�cֺ��I�o��3q�u�2�U�qO����"j�}�Kktp�tvS�j��2P.���=�&��>�{V>��u���W��{k$�2��z�� ��v�}�h�������/�*�ܥ�}��ؕ�|���^3�~���M: f[�,˝`���+��@�U���B�m=�_�W�� �/Ɋ>��j3>�0y}]�Cl�����Ӧ7�J��W%������J<ey��ߎ�+Ƣ�5�߈s��u/��xWj:���i��=]�(n���]��~TG\<������_l�7�BS�����>��i�ͫ�]�:Jy���_�aM/��
��NO���myj{{w���sa����g�����O���q���EgO��97]�z�㕁���l��e��nr4轻 UթVc�vF� ���
���vC�|����οz�����髗���FNTe�H��r�A����iz���ct��������W=���Q�>�.�G����Ν�mZ���%Z��X:V�K�����c��Nݐ(:� rt ��i���n�m���������,��Q;T/���N�c��G�v��fe�¨��P"xws�#���]��kk�x�@� ���	�2���L|�w�VU4=Hn^�}\��%|�+��<3����n'��]9�RyM�grL��u����;���7ϰ�4���J#��8|	��f��_Ӡ�w��~^sb�O%�9ם�I�)�=�L٫��ݯ���Eh�Et��5I��Ѯ?N���}R'C�:���ur,rW��O������9t��
����=��ܜ�^twg<ax�ӽ�eю�դr4<�0�|�߯l^ś ��c�h�1鮁T��y��i̝&ww�P,Z�8_�����2M�%qG{
�r�Χ�����c7��:^������q��Q��-������W�����ƪ�WW���9���/�M��BM�O�rz5Wk!{y�X���M5�豸�η����z����u|�����.?����R���q%3��`����Rȍ�낅/u��ytL�V5����ɘ��Kմ�r�x�!��?f��dh�1*]�DɚA,�@n��$�u6�dT�R\k2�1�e,���)f�հ�-J'����Z/��X�4Q�������ż侖�'���� �{�GZ�fm���_�~7c@�@'�V�>>�W�=k��*[�g�uX�Z~�6�������	L�n�mg�>N���d5��C�ﾽ���r�>��o��gk�=a5�I�.?�??g9}vM���T�������� �}ݞ�ɕo'��臨��ڏ�wa���{��F���j#�^>��n�{<�\P����\���>��"�����Tݪ�ͯ5����2�V��<�r�~�/r��F{]P�z�?<��Ndݸs=ҫ����ڊ~ ���;��|�F#�'6��0Ne�Vl���p���[A�Ϋ�<�d
Ѱ3�,�$E�R�[����r]��Ч�@��ʵ�!��h�u1��{�sͿ^m?�e�����F�M��-q�9'L�E��յØ����5
����w������b������������? ��S&Ҡ��qp�:�9[�[bΨT��ݗR,�!̛���u�yn��}Iʽ��˂,G��Ѥ�$�Z��#JRBޱGs�i_#۠�X���
�+�8T�7o>lr����C#����9��R�q��Dn� ��)��g8_P�]]Nlq{m��x�h��6Zm��S2oq���gH���L���P���infi����|OP�z7+��;5�=g�7��&����ugqM<�u�۰�8��W"mͪEZn	�[4��ڝ�..�C@[�{��MNŨC/�ѯ �[,�G�"�GN��sO�<�C���:3�9�'g�� ���*X���}�r����-'����UA]v�C;_�I�]aC���[Z�]G��Z���R�����l����w���|���7��b����Kcڐ�R�I��7h�]�+dO��!�[U���Z��_'@���ʜ��>��R�;�|atzi�w��i���\E%���f��Ag��3�>1L_N��rV<�]�E<�,%.f�h�W�P�����iO]6�S2��rմ�F<i\��`��zQu�+6e^�[wy�e�x�+;Q��o݊n���6��X�ف+TIIw"e�7Z�8�`��������ւ�}� �tMҐpٕ��j����y���U���V�khc]�ti��]d}��@Q���6�J����.��i^�.p�a���u�g�ٹ���O�嗤б���{�ߤI�C�%�����<l��d�^Q�s{af�6��xPM�M隁K��rm3�k��D�Wle�w�pd�T���̎���P+G'*��C.1��j���bE�]���
�M��ݽqQco@M��36M�^eݍ����gA���*Y��2Un�.�dZE�J>�K�z,��uU��	ݴ.�Ҿ��b,u�,�����[ӻ�.P|�K���:��#�j�gc�<�ǖ��|�Mٗ-p�/A�@�����T�Q��梁��]�JSW�&,�*t��T���ܶ�IH*�K;x+jȝ�K��D���t[�Qu버76�=lm�Zy�ӝ�#n�	�����sg(J@��!]|�]X�;C�`#�z�B_O��4���%�si�E�/�OP*�}pc��1-�sM�)�;�S���>L-�x��:\�J*@�ݕ͞�pkؙ���f>ή�̕eW;q�!n����[���\��u�2��+�Vu,�lT=P�hc�f�s-u�a�z�9x�J�w�wp�U�Nv��v�[��V;�I�ķ���r�5���Vfv��9F�|�IawPb��/X4���x����%�!Y�Cx���v����v-�q.��1Z�+Q��}���w�??����#F���&�f$�j��ڍ�W�Qy�UQQ�<�a��[@g>=z�?������~�_��v�X��ASF�-���<O��Cy�:���mlkF4�?�������~?���������߶���sh��mP�.cU�Ʃ1E��&�W|���0x�4Q�hգcb+Ns���?�������~?��ޟ�{��pm�V�C�I}��y�͵kcl�j��k�M�lM��&���\y�3����}���_������~=׽&�i�0hi����4EZ�؋�<�l���F4j"��b���,z5x�c1!�1�64!�� i�03��DM��P��T�QE1m�š�
��d�(��F4��5���9*(c6�Z�gm�����3EF4��h�	�Н$[��;lE���|��SN18y��1Р�I��M�61V�ڪ)+Z&vͲ�z�y�;)'Z�
&�F�)�(��4�Ph�4MV��*l�L|ƈ
��$Z�٬N�����D���msG�&�x|���M��:�:v>���% �z'Z��i�d:�l��)�.��j�m��$n��U��|�͸ʽ�||�o7�����������{1�r��6@m�l3k����w�~Cҫ	���^�#/Ԙ��OЙt��k����%ߐ���B-ms]8��v>p5�fP�����o4/5�1\��S�aށ�J+�#WT���������;E-@3�.-۲}c'���� v��"W@2�L�iv����J�3�lh��@xv��=uL[��͚������������D��F��F+8��|�ElD	~�sH�n���_�Y��ytM�7�������d����U��Q�*A�W#�>UH�UY�1n����]:�ni�ܚdɽ�lKbQ�a6�
����D�p-�|��H�/�D�z����9��&�p-�&#c��Nm��R�.�-�@6��OV��)�qx�;.��8p�V
��68�g�j���<�����A2&�[��z1�����R�>�� M��yV����kW��k��n卧������������w��}���7�=�Я;�ZZ�&���G�q���n�1�W��v��X��:"��{�ܫ�H	Y^�H�1}@�?���U�/�Z���]�/�Ƀ���9���˛,/r0c)�l�ֻ۟LP��޾w��׉�C�gY;F�Nx�:������,��� 1!9�qus��ʢwku8�]m#	9��gw	�VX5����%1{��t/��2��苓��E}���5W,�VZ��M��Y�*��\�+JO0m_�����o7�'	{<� ,+ͻ�C���~&�L8�p��ͭ@=����Mć����j�{��[FV��s>�:�k_�����v�����y�x�<5n��
���y�_/�;:|�p̨�Z���ř��9�ѽ��3wv^����^���Ҙe_N�^�sf������cT��4 -��%�`W��,ojq��T��,�ƥ1��G����S��z|-��{d?Q��G�\�k,34�mf���wI�Z�ׇ��7&{�v���a>��o���.CY��m��z��c��(A��4��3@把���ng��~ �?��'7����g櫜	2�c�� �=�T_y���D�Ti�J#07^�\�׼,� /�[y����Ƶ�/����P��������8����������uV)����-8q�t ����	%�=�u [5%>�#��:�m10�!��\O� ��#��������Ý1�v�fˌX�M����Ǩ�M�)z�pe5���fy������9��~���0�>9�D{Q�7��u��
�p?t�  ��h�=H�>�dA\���_[����+/�?���4��v2rᦵ"���g-@�Z��K�y��Q\4q�>��z��)a�I�o�*��D6Jo�Qmr��y��]�]׮�z�҃�ǁ�ZU�m+��GnN�㖞Y#�D�q����5uF�����YF�������;#3$�p���9V�+{��Q�G���p��ɍ9I�(�z�?�ff��F���_����۾�T�G�3�6��D��a jz݀dED����6���yNӻCi%���le��{_��k�n�<Z� 7"!�k� y4[{i���ؗJ���̤�ni���@;��\dx�����A�k�����<7�u�y^����������=�gd�3�>4�؜���W(�*37����qr��%ɽ��0��_��Uxl���y�n��mL!0�!������n���"�����I�f��A{��0�5��6��6�b�۩�����_��Ő1�����/�n��M[M���۳�� S>9���,�/���q�<�.�;��XN�S��jL5�a.ļ�J�����7}���Ҁ�k�l;��,�'�lTlXЪ���U�����Tw?����Z�
k�ڳ����p�sޞ����j��?���&A���5	�<�y`�N0�5J��,q�{����\����.&���g;E=��{
@����������y���S?����O��m�����DK>/	��9?���nr�X����WNʷ�L�{��9�����N�w���� ? Nykvos��M�lap(K�|a>^h���~��YX��6�P��zRb�,��an��;�����g��1�Sg�~�C���V�Ϡ�j��2{_���n��=Z#ò��1�_��B_{��+j(�e íQ��
.�jqJ��s{m�j�r��[c�l��}[�<������4�32{��>��￯^�~@�i$q�l�7���pw�^4�p������.����R#��-�Z�Q#���x-y�/b�.�ٛ��}O�A����7����lPwbk�m���ͺ}x~C��~`�����⿭�� ���b׈����
����rG�����o���x�Z�E��?v��!o�߀**��L�f��G�%#фBh�g�2��(V:�ɛ!��r�i�X���9O 2�by��l�9�
 o�5<�y~��q�|�_�,]�5��Ȫ�b�3�6߱�լ=�\/��Z%�ߝ���M6� -8M�������sf�^�F=ݩ�$�zx�2|��!��2X����:��L���7����3@�W��Ơ]����ۏfs��ɱ�<����|ݑ�����)�T����ʹ�m��|���qg��x��
'r��O����� Ʈ#���L�ov�(�	g��)>���A)c�\��\E^M.���͹\�ՙ���ɠx�	�p�*���j��l쮔��7#"8�K��8[f'�u�����w�ue��8�PK>�)M�Lɍj��(�Á����]S�iu���YA�f-��+�j��Dx�m�����gy��΂��0�w�v�v�gGl�owU���E�VX@��U�&�p�{��n|�W�=z���ۛ�+~fffe����g�mᵖ8�虈!�7���
���4{�����#���8:���B�}���rRnӧk�@^�\
m�F�/�#5w��Ak�k�Ǽ��S�Ő�a�J>��_`�>�Jݜ�F�<-ߘ-����<}���
�i|N�I�66�@ևm��Ey�$�(
�f���=[op\�n�D�bI^���9�^��	|�E���h���^��o3ǁ8�"@�~|C��'��s����|y_C�0�}�AaN4t�x/HQ��*2������(فk� +��q�IMx�(����ɛ���T(�����|�^wyy�  ,Sdx;Dq�j㊊��(׳/��q�\�g>jo1Jp���e�
��T�uC�qύ��u��!��L�4��؜�si�q������a7��{y�Tw2�\��Fs����v {
DY��j/��'+���_A�R(��[@�R]�_�ީ�pҎ���ESN�1����v06�s�{K�� 9IfOA% P�\�U��(<���NY!������R��V�J����g��,+���w@�k�iƧ�t1�0	��K&����m��W�Y�ߖ��Q���S�;Q��9"�)��g�������^ڋ�5���'T��A���.�zO�����-$$��8�q�ia^.ǭ��J9=���<���6ws4{2Q3:=�˛L�G[�� k�5r��7�"����Sћ}����M�K��>����z���?�f	�`����o9�g�I��|�7�c��׀:��8��QEխ��[ ��ǻ	N3�y���#U����E���� a�㱍l��N)�`!=��b����T�� &&�м��_j�9�g�B�f";�q�WM'�
ꋇ��/w�|~��q�/�'�_��:��=���#R�`9�`��)�(��M2���^�6��z���z��ʆ��[����s��*��H  ��?W��;H������d���X�������5��k�z=�q����6��K�؀=����=�g©8���ɀ�7"y���^�^�]�1o+m�� '��.��}Pd�⌖E�a��cD�C��C���:�a"��j���ww���8\#��r]z�
�yH�� s���+��|"�}p}z=w�=k��'z���W����ïm:!ػ"��l�ҽ�3\2��6�`0[�TV8���/v )�X��1���(�k�頼�f�s��8�v�'x����>g��͋���v�Ο	�N��9܏ �Y�7_B��;
�*p(�L2�˓V�*M������3Niz�����1Ϭ6-�0���Wɟ�������_�~�W�������Һ[p[0*���(��&�x�lҒ-uL+3UD��M��bx�3���#_p��W0��C�wZu�-��ۼH=Q��qj��u��\`L|5�TzS뼵Q�8�f���]}�a�KjÛ۶^���5�_]Q�51iԒdм8�����.���uD�"�*yB
�Ww>�@?��7���;	�����G�e���a�{z��~�v@.- 7�	�����'���ڽ�0HKy���6���� [{gf������7X;�cm�&d��Z ,�-'a���
wZ@�3{��yח�>���* �֥+k�c1�oC$�{�֭q�������c~F`0!����~QP����߲���t=�4����A>���m��!�-��i�p/�cXH��[ �\ ���M�]�[q\�S=�Ȧ�kӗ�����Z�{��.ߊ³�~��5^`{�-~���1och�mg6�g�`�ˇq��qP������Ʒ��a"�/��wXh��z�=N��K�	NY���q�M^>�_*`n��TS	��B�� ?���ᧅ����P�%�0y(1_���T:eՒ !��0�f�q��uL��vK�V_-w5a��C��k��2��|+z��%j�Ik=ƣ @��h?aCh���{�G�x���z��Y�n�S&C��hh;�9������y��{/��E�sm+W�C�}�^������8��5�^�m�gPPZ��u�<�M5�ߋ�4�Xh�MF��s��Z��!�<Wv�Д�(\`T%���mF��\�W�K�ˏD��
Φ P�$õ36`"L:�YR``&_22��mk ��1��gQ����RO�U}��[���W���{���-��Kn���r�Iٜ�����K��-h�T�x���Q�﫵�|�3߼*��P��o{�����Q�]����}��X����\{v�j8��G%��(�q�Aj�1\˗=S�ON���N!�]�F��f�&7�w�0f��9=	��xh>u�oh���T���k�Jڧn-U��C�e.#��^��\=�F����wT�goD��O�y�ο��~.��8|u���;{�Ɍv�3sG����z�>dF�>)�ekG�?A?w�Fj�s�h���Aׅ�]��
S�r��[E��<�
W��3�o����F�^��U���Cx�� 뾎
�w�^ĳÚ��8?��W�%�m�[`o�~��	f�S���X�4�D(u>5�,h�,%����Bz0��W��$j4�gN5�����,ZPl�"5�|�	@;��C�	V� #��ǚ��.���]J���fU�g:�����"�|h�bp�d�v��C�H���J}��$�	�6N�hc<,����O����J�u?��Ǒ8nbiw���f��,����c�.~����Gg��S	ndLD'����]�_]�.���b�O����+�~ŕ�-ٗ0����ot�6g���Dϐg���dU�*TX��]�*�9��b��y����P�ni�����i�ҵ���9��.�T�#w��F�����c�|�.7'v|�u5`̫;�}(ș*pQN��7�-����X5`=y�u��H��!b߿<�ϟH?��s�g9��H��)��:�/*B�s�<�7C�Y�h
b��鶟mʻ��_D
�م�o������<6����/��~�-����Y�ҺW;s�t�Ft��
i�iM�Wt�d�YqX��1�WU�W�!�X��]��@{��ݏ'��m���u�R��9�.v"�ϱ�~m��c�ifRZ�ɹj[��WoI���S�d���/l��?4[��3�iO7�fr6"�*���Q͋f���Q���`�f3p�S�o�?4Ʀ�Pk_f� |k����Ѧ4jeq���F���3�W�8����_n�9����[���\�@Z���b� Bƙ��pl��� P�P�u-����Uf�7�|B݀��m�<�U��ʌn��`1�lT,י�xΘ;Ơ��7�-hi�ʷ�V�`������n��a�r��ю�^�Ȏ��cc��^o_�}��JgG�ւ=��>�4�@�e�5��a����e�ٯ���B�0���ϱH�m�m���_����94 s��[A
w�x�6�/��Mv�ޚ�5��¢1=˳�d�:�%6˄�+�;2}c(���H�h �, '��p_�e��w(��p̑�)3�w�*�+���{��Q��F�-0�خp��bk�opҝ '���V��1F�3���>_�4$��m��H*ݼ��;���s��2��FCa�L�W�"��7X�u����|�h��߫����_���q�s�3���M*P�*��~>��[~�_�~������:���KC�/�q����7�J-|�V��Ҳ��R"��Ԛ>�d~���g���,����n�n�x��׮\�w������L?��8X��ǯ⟳��"K�^t߸E�[d����ޖ��)��ń�[+:�O�E����gţ����~R���ʄ���K�lK9�z�����
�A��|d���e�u���S7_���P�7>�����Ŵ\	d�]j���6��~﹂y�>��cU�S��,y��M�Y�%�e*��})@�hi��;nιE;'�s9��0���r�i�(�ɶƸ="m�4
�8~�:'��C�鷈[B�$�%��r��z3�v��,|�����CS�^j�L������.��2��faˡ���-�9�9So��<�+$ =��^���3�m�k��
��j����~0Wt��HxyG��V��9����)�/ُG��@�l��]a����-�=��ι�]1&�t6��� �u�C�Bm�8�K�\n�ʀR`��sR�>5��Q�Ҏ>i!d��6A�������m��-3�W?T���]��ӺP�L��-Gm��
Z�'��1U�$,���kr��On�vP�}o':��k�|(WaŚ�Yr�M��"���Z�-�Vq����xWP�;^_|'��`��Y�h�i�ڊ�ڻ̡����.m{��[��

��
�8u,�����+��[̽�:y�DɷW8��F��}\��U�ӨkN"d=�1VgH�[鵓���V!��=��`�e�*鼆����V(�sǦ�)���p��
W[)�n(�����5�*�yw�w\s:Hղ#L�#x�nq�r�����J��8=G�.Ay6PU�k���������l���}(�tE��&��ty+*��7R.�Is\:3������-��W�m`�t
���ݱ�H��ٰ{(��Y�i��!��u����,l:�hYSu4�4r�0`���t���Vl����f���yu�6c��*�`��ˋ��v<��`���r��D�5&�M�
hQ��(%��vb��;��n�"{��\KǼ��4�˻�KKb�z�ݕϷd�/#3�6&��S�Q%Ө�v�ͧve�C�,�aƍkF#�ޥc6Q�z�.���6Ju:� r��83���G4�\bL電�a}ms��Q2��re��v�z
���فU���=���m�QkȄ����� �zXFU�`>�]��۫�v>ͨ.;��'<_���[_,�=1�-�K`��űa!N���d�`�h��.�N^�h�?���зB����U�~d�'���4�P��[Ai�&q3j���r��{�eS���ץ����8p&��x����I�;©��g����>�q��E%soSB3���YK�ُ�MU���1T:����ތ�C��A��92�.�	Y�^$���J3����Y4�6Q����Ҿ�|q��0\��&���e��/(��ow]&&�=�Ũ��\��Q :�V[|���e�x�����3/T�9�����:]>���;2��N
�|B���;y$��N�����2ыd��DP���ޡ:J�%���5`
v�]r�-����̵W�E�d�5�r��g���*U���Ы@����<J��#��P��{`!�/��6�ѕ�����f�S�P)-ͽ�[�la*�Ya<s�R�/N������l(�[0����͡�oS�r���R�z�>��&ó�Q�r5�-�fnc�Z�y��Zaµ�"��\�0�5���u�V��Qh�X��ݰ�ټl�F#3Y����rp���4"ޑ�R�%��%��=W>u)>�xze���A(�k'95��,��.G��]�6e,P�f��y���wRJ.d����u�*��]��*�ɚ$W=�7hLա��ЕŰv�]ݰΣ��.����*,�g�\$�rA?B�t�&Q��E�'���X���DQEM�!?AM�$�Ƅ�ʔ�RHnU�C����M߆��k1D�C���o�iRk����y��}���Q��RQ�T���y�)��EUA�Q��`���<<�N�kQ&g>>���������~?����~���:"�5��֨��(�Jq5�h5L[`���`� ����*��[ljh����������~�_������~|�TUCD�ݍj��&�gl��QG�������ٟO�����?_������?��k����j����QZ�UDM��UU孱�ЛUy��QLF�`�l�N(�*�����o^�������~�_����.⚢
-����DMDA1QSX�
����v5h���A�k]ؚ�ؚ��ff�b�ggf��#�b�N���(���*!��LDh�lh��*ua�D�1V�"�MV��*�Q��m�5Z�U٢5�*�Z���f������i�VqDձ�j+F���h�Z4blmQ0T�DTF�cmy>^1E��H�#Ad41�6� �m��iF�!��QM��Td��EMMTh�T�^�Q$yb"�O}��y��!��4�!��o�-\���+�-��̭�e�0����es�>|�^�[7:M[R�r���eCAt(���7��'Cc
h�QH#F@���� �DJ�9�����$I	�3� g8 Ъ�#J'�=<��տ9�YE}����MY�+����{��2��ҿ�g���,��G���Ž���>�/?6�fA�G��~j���b��<ƙ� ��O��졆��z���Mt�<�y&~�ӝ�~�e|ˊ���)��$^:�du�#��ssS��^k*+���=7a�&�'4su�%���M�8e�
����K~�LM|��jH�Ƀ����fhf����V���]��\��3�v���R�t\PnJ�5�hNޮ�w�OKϠg��T��͛���̈��5�]H���2�P���v�3�Z-�R�<�����r�
XE��ݑ
�@Ѳ��R�eҵn�^��j`@Rײ�5� ����A��0!�WMü��0��!i�<TOI=��cF/:e�)�döxK�zi�8)��P��^��Ȝ����5ֆ�-���5���s6䨇[P�� ���E~V��ߌ��'�����u�vE'OL2�5��U��4TuUc��g��/��r ��3=�Y�ciٍw����#����k�Y�E|(��%�l��^E��g/�g�$�F:�iU*�Uc1��������۵KmU��Ml����Śo��0���STK�M��oQ%q4�e�n�����+2N�wX��V���j��X񑱵��7����k����߻��������8A�p��	�GB�R�Ċ#fykOCu{�j�"mm�׫W���Tm!+a�}0�_|���P�/W��3o��8J���h����@�0�����ٸ�\��O����L�c
���	`��8n�nߌU%w�>����t\�^�i��F�In/�*Sm�ɽE����Z�`
�����T��v�Z_��!%������dY~/^mqU����hL^81E6�nnZ������������#P5p����C&b ;��Ӄ����P�T��]���ٽ]�Ƽ�F�}��T�n�0U�R�Y�V���!Z�x�y��?D��0��� �8���^���&V���xJ��l����5r��#�[9�pw�x+�
�M�\��U�)�ƨ���J�粓�idY���IG5ߑ��#��~�Ќ� Nyh���'�ѥ�ױ�!�4�,�l����_��!�}9A����1Wq}ʥP���|�'k^��z#�[3Z:w��cif޽>D�zq��c��5�_�bz�ώ��}j�#׬��fڥG\��gOD�.��|�� �'fJ/m��I��XKD6aȹ]&'�Be�v��}�c�T){��}���L���DH!K�+35���'\��U�uVyJe�it����8��ww�>��͒�)|8uj/`�l��++
����k�����}�.s�� ����t�"J� '?�?}�������;��}ի���k��+f{^m1v�7KŜψ|+�l�bL���U�cH�k3�׸p��\���f��2�>g5�f��	q������1i��c�楇6(��k�ٔ+��`��ڞ��2�4a�Q�9����g���~���CZ�ہ]N��&]��Sk6:��K�zi0�P*���ŕ���P��>w���jz[�m:i��;mi������#�8�Ia.������1��(��m�jm�
���,����X�C*�M*^����=����F?��^ԯ5x:��A�$�	��ɝ�ީM�}�^7XȦ�b�����uFu���fvR���-�6�oG�~[j�&�����1���ƫ+�9�.��B.ý\e���y�;�R�~e�P_����	�F������.�ҩ��Jy��Q�T�}q\G<�_Ei\)��X�H���znm/��6�:��C�m�!���ˤ(�8^���J�O�6ڋ �.b��n[��"|5H��;���fA �.���>���*¼��ھ�g��5j*Q��������M=m�JDO�[A��ӏ�5���BN�rx�?b�r���}�I5�%���sb诮�Jn��E�N��K�<�mMMEۑn�aAb�9�����ͷ��=B?TeB�s�\�s�H �"�H��Z���h*i�Q`!�������e��s^k��<cZG��u��k�Z��z1�lU�%�Nד��/��C���X.�.��Zz���j�.��*�v����%WkV�6����~�'�Ȓ�l�@�>�A��eR�X~[��$���k5l�͝�~�.zJ��{��;��9̾�Ϙ,�����&N!_��=~����`�ל7h�t\癫Ͱ)�Zv*�N�i��5J9���*3|�._*��g *�7�E�����c��n��.Y9J������0�ZB�hG�?}i����e;UȀw蘚����3Q�;����̇�Uoa����@��$#)�?�T���#�]�����Y����\r�Ф��h���[b�6��]�<���B�,u�Wˮ۰+��US���8lP�F�;PR#�]z:���T�@@;ƿ�W@-`c�������Z�KV�E6�Jo�6��&�o����j�X�v[���>�S[P��H>���'�q��k����Ɯ�z���vI��ۮ0��70P��.�u�:,Ս���d��U����@���D�pLG2)����ƥ�{�[[1���&F]I���@a�kF�P�+��D����u�q=ʝ/X��i���Q��4�Ƿ�'��7f�p��;'�L';O|PW�v]dr@�3��m1@�Eĉ� �{�(�s�]*�r(g8|�=�����{�%R㔃:��c�����nWnqǡ{aڬ��y�"��jפ�a��~��P�F6F���q.j1h�@�Qu���z���W��P���}YP�G�Ư�9P��鲏��Gv�U��84���Q��Z��*D�<�ǒ辘��H��T8�wla���p'��J9�n�t�*V&N���D����l�j��~���t���D�c<6_F;�l}S���:�˪��v�Y��/	=K�r^�?4x^��`�8a�g����KD��D����쇧d�8�p;�����]4|mZVH��O�!�y�*���Σ�D�l�����SQ�C3���#����?U_��T^��~hE��'�L�'f� ��o�.3����;H���VmUY����^k�1W���9�7��v�<E��2�+ч���0<wʀ����c'1y��l�!��߳�+|T���0��ik�]b|���,]�9hw�@C,����⯨�>z�B��p�Ђ����
��n�1q`T�����ݶ�f���O)�uY��u5�މ��Ϫe}���'q!,҅���*���t�$oX>}��s��:��I2w�9��z��/�m��Ė��HW��K²��7�9A
��&��<��PnEATcev��HFm#La��ǈ���ޯ\�x_�'eF��s�S9ʦ�Q)E�=>~�������z�a� } b�h�>��E�dLj+���yMÊ31�K�T��Z�����|��x��=B��޺cD^�)Q}Ό������+s��W��[
v5;wX�T��u@Зd�D��g�c]��Z�����k�`)��}{f�����-�w��u��Y���(�q[�m2+�^Dw���Q~��с�r��X�����:��J����K�^tx�9B�д/(R99B��4�d�E�C �h��x4X���3��am��\��`3@9��}�F}8Ų���S�F�l�q71�.^C����L�YK�C���6�\Ј���)�������UΚ��}0�v�In.^a �ڤmJ�t�,ϼ/;k���야$�P;�U��C����k��ъ|�}�@,���
���2Y������788:��{;�������C	Xz�p�5
!?�ɺ�ǲ-f��<_��z;�4τ4�V�KOS��nS�1x��S�Eٷ�cC ���#�yP��ʿE��~�\�2��s.�kʚ���7r�_@�T�Q��]��x��+^q]
�b!�Bd(�e=J�h<��Sw���V�}�os��c�b��擌m���!۟at��+p9��	�䃯e.ڳ��}0l�Y9�I�B�����}���}�_ҁ� �I���hBs�\� �P'8ТR�B��� P�4�@�������?�^V!���rԓCZxűb�0m�ql�`9�/��[��X������h���.jg��kW����}���k��U�5r�4y0��ϗ���?=����|3��_Dya��}0]��$x]A�j�w��˼0�?���M�^��ʎ!GW-CF������h�Ij�Ɣ?~1x�P�@5"���� t���R�`�x�H�h��ص�����ٰ�G:3^]�Z�G�H�ED��TF7�=�q�w!�-�;B��ƥ������٣�����?
�t�_�D�U#���[?*5���28˧G`�����Xի:7���P�Z;�<��%�+\{k��~�H�pJ&��~p?#�G�W(����H�kv�=٥�b��ӌ'�L��ګ�I^X��ʈy�f\��v��Ml�E��LO1�|�f����]�ݑ�Θp�a2�fq�b��ߦ�-,�a��C4�L�y/Jx]�	cED�����@�Y"��65��2�$睹�y8�QM��Um�k=X�Y��~���ۃ�~YV4v�f�vmJ�EwY����G�s�%���5�C��E[�ĀJ뷱^�9��k�x$��T�Ce�n;��s���,I��O�e����Ң;.�v�Y ��&�g;��}<���޹�=��z<?��4?�*�s�9ȩ��DР������ReTxu*l��kjo|�<��&h��}�	��d>��8�ǧ-���ad�|Ƅ�nNnV�l�hWZ����-Ü�1]E����������}��_7�Ќ��G6"SE��e �7��t	��v�{[5�37�>:1r��y�n<���Z��?�cP�Wڇ�\}����]H@���_T�-]u<�#d��!�����`QD��_��cG�j�)�QJ�*�h-,�0�x��{;Zm��c�.��yhhcu5����Gς�cY�)�4؞U�I5H�vo3;n��n�A�LʵMy�:k��K�����i��:4��
{����&P�'���.C|�=�g��?��ku�vǇ�L�(!F�|c8�oz�� F���&o�z����O�z���;7wlW?�~�_cv?��"�����	�E�z�PQC]�vFez=�r1�vn�]��ƮSZ�2Z�(a�.3��װp�M #3����Rڃ�J�Uk�Nk3���Q8��"z93/2$� �ޢaښچ��A�ç,�w��*�	g~$�]�X�}�؟}������/��tVD��P��43L�w�:�>��,��p��exK�n���N���~���������RD:R�@����(˙Q	5ɵ&W�n������)ѾSy.3�����L�iS{ˎh�n�O�3fn�U�"�<zhR
�,vɶL��^m�ҩ�O�� ҄� �s�9�!�P(B���m����jk-������5S�,�_����#�@��>�L���bsϖeC	;�"J��6u埳j�9��Ԗ�M�S�	j@Lxn��@�
ޱ�b�ĲdY2پH�Պ\[x<5,���oTI��u�-i�ދB"�E�Fy�����h��m���$�ߵ��bz.��m�ev���&�V`'��Y^d�M��m��G�$Zm��\?�-�4R�a8����T���������DcZF>�Z׹iz�[j��<z�Ϭ50�^S�.��L$��@���g�L�ޮ{Y�mw\q��q�p��L�}�R1�Q�^m�(�g�0(�O8�}F/���nl�;�cO!�����]p���mJ�D3�������^<�1��mih7fk?t�ՅԾ�5�'�l��S��o=x^\�'�d���BƉl��{f��-�o���Ndk �#�"?F0x�G}OE�{鯌	��@s��lO^����.�~���jvؿ�GvG�G΀���~?0Y]����Έ��u��tb�`�c8��ce7rJn�Xб&0�8i�{�[�8�y��pӾ�/�2�6�f�>B��8R0����#=�3�=t���I�?�@H�jb�9���s4p;x��;�yK׹H&���$9�y7�ܹ*=>ÈĦ|�m ��kbŉ��ǈ��t��9������}����iP C8AЌ�*�s���P���4)H�!dv��0��Q�F�2��h�,���ݘ��;���}t 2���'��͗�Ke0��"⨶��ǌ!���Wvf�#m�x���B?*ȗ�t����w��Y�(��;��]���|�I��x!֤m7F�0/|ΔT�N�я���{�i�����W<��_cV`}�=��$?���j���z3��^���f���H�5�ty�E��8O�<��Dֺ���=��L(%�Kո����d�8�,a�thȖ�]7�"p��v)������l�Y�i/��=�ϖ[�f�`��y��SW�<���=C�b}1]������+�����^� �%@�e�!Ѐ�Z�~{vbA�v��ן)�e�/�5�jPS�Y�$g��$�z�d�sa��S��Zcju�t���7dd�����T0�}�:���^�oHq�0�8�,��aǎ�71k?/�DGN�|�������B���c��[8ٯcm
]���kb�w�! ��v!O.��V����^�y��|��d�������o�V^@e�x>���oՏQ����O���Pc�榧�4��v"�dE͵�W�o�v��=z�JJmL��X]�`"��/t7R2i�X�������d�Y�y\0ܫ�+bjN�̮,�һ�J�[Vw|V7*�����Y�0�E3�{=p��U�J�@��h,V���&�:�=Wl�"R'���m�cpd�o{�$:�U4��J"�U�-黴2��0�U��8�a�"��	�2��u5ɗ��q��ކ���wѰ5���$+/.�W�W �'�y�9�k�9����r���t
�n�pV�.��A�U5���ZSY��)nV2�P��y#�m��_q��C��$�u��с��P�S�����h0�r�yc'z�R*'tbT�i�ݪ�ܘOX������	�[S�o^{]`�o��U������L�5vA�1����%�+�`S�w���GEi�ж�l����7��sx�l�4N�SOS����.Q�ƭ��6�����KH�8�u��Y��xL���xFsKX�rwcJTm�*�j�J{������/+��J��%�[C0�)���x�\�h�ˇיw8�U�-f��,��Aj�o���jm��[*m�D�c�Y���d]]^��̏���]�S��Z�܌�Dr���;��`7!����B`�3[sl`�\Hl$��앚�oR��!(v�ƭ�'�cw�R�;ul�w��k;�1���3�ොӎ��Z͕���P�O)���C��{M7�cڸ�ӯ�-)�����ڕn���X{��9�R�.�IVA}ʋ�G���pLu�_uE���!wݵ��d[ьC���U��&^��-p��T8�d���GvK��s�QQ�d䣸�0M�08ƅ�E^�0`��W��V�`ܭ�w��(�4����30%{�ڥ`�e>/�i��u��س`Ḩ��ok���ʓ{���KLBKз�B3b6.�ռ��?�er�sQ
��{��Ic�"�ڂ�_@�!�s��n_�3vRX��Y�Esyb�w���y-oLG ��h��;<1+2��C���hn�R�Y��gG�.�+���rg�����C0��L{���K���p�}p�%��S���ѕ�a5i��[���k/c�W:��0e#�z_;ŷ��%rv�l}���+��G'mM��K�\�5i�Ksw]]E)����F�J�sw譮��">Y�HH[oe��#�Srv���� ͺԮ�~�ִ�a';��tj��c�K�E�[�;w�̛�>�,C�Sv�wc>ڜ��X�o4�Ҝ��mڶ/k k,�s)���P'��bl�cELٍh/��<#l�VƠ�b ��*�(��cY��?^�~=~�_�������U��'Z�&֪i�Fמo6��*($�6qt�[bJ��֪f�|s��z�����~�_������~�(�k��>Z
<�5EQQLWvb��c�q^�jb����ŭ���z�������~�_������_�6����ͫd�}�TSUPy��͛�c4\����5IUKkP^�Ϗ^�~�~?������~������ݪ��������킊J*�j���iƶ��v�ϫUUE3yj"�޶<�V �mgɅ`�Lޣ�*�Ym�SI%IE&��h�
�
u��Q�6"�(�H�*
��(�j��E�f��#gj���bJ(�֪���CQy�h��׾c�ff����̛[cDZ��E�L�M�QIE�L�Gͦ���i*"�j#��<&�c�)��om��Ӣ->g]�����éq5];WM��U��Z�/2�yP�>΃��{�3w���ܼ�8�A�F�R,�2�c�E�2瞸}�{���~����_�W�*O��MP� �Q���Np�����m�L[��6��MKzCHf�xW�`���M�5O6�*Vw����N'��<�|���,���_�!�=;B0[y�c�y�dMٞ.���O7 e����X{�n
�����5�Xc�|��- ���B�G�	����kL��S���]��s.Ԭ�n�W���Ђ�%�(,8-j��{N��|�^n���Qz��oʜh��u��'�\A����f�[>��33Z��i2-=O�B���֐8�>>$�Y p�
�?���:��T�啤�Z0ıd#���q������nBV� �p��QP�/��._��qM��{�xy��U���l�L1!F�!���sL﮼@��p�}G�q<ev6�u�'g��Z����}@q"n5DV;c�L2!��|n�*%�X���g_E_'��j���mM���!fi��5���k�G���z߆!���Pag�&�����9�;����_u�|{��k*E��p�n��}P톃Ķ�Fz�@��)C��zgk��82���q��{d}�����X��N2�*/V����ڎ�J	zg��r�N����K��"]_S�p�y���Ly�n��[9R%_[�Y;���G�{���@a�����@��H��6nA��i�]=s����(���(hs�M!@3���Y�D� 4 � �)@�!���wϝ����~������_�	j�݊g�A}q���a������� (�`�=I~�Lro����g�㰋��<�G��}�s�1MJ���8����[Q"ݙ�;ݽ�Sh�����=6]����v
�D��?~jy�kg��C�wL�=Ʃ�{[�@%u�`<��'�2*s�)��KhO�w:�F��0���B sc[���Hu�0�6�Şi�S	�x%V��
�P���S]���Ů/1�K}�?S�U�6�������O��Dh��6_t��R��
��<.~��"��0�Q�ɖ �=�u��R���8x��l�c���.����7(>�>��S��)XY��;�o˷���z��B.VS�.%�ix��J,�����&���_b��Qx��;��'��DB�yp���6�eMh�KV����	�RQ����L�Dƈ�6k�m݁a���ʫ��g�ΕvkK�K�t��ymg�͖�)��5�P�^�;�3�j��MK��m5O��ט���S�|1��E �9�ͅ����j`cG�#���O�>�E�7~���J��d��*?��V|�5$���'���o�I�Z��`ȫsS#���~k���j�k~��9ő�C�k�n7�I�lF�*St�9v5���,�����a��`���f�y�����
c9ѯ�Q>h�����KЋ����<fwIc�	W�Z�,3��㘤����a'UT
Dp���)��93��iI� Nr�� BE
J���r|�W�8�X͌E��WŬ:	���͐(�o3��02B�/X�]����<�_�)μtB��B�se�Wi��U��WI`�%i2�A2q��.���:{-��wk�3���h��3�R{��͆:��+��An�/��/Õ7培D�ę�o�6'��	��Wv���\,�V��:�z���P���B���:�e�s%]�VTc��f�!�N����vC�Z�S(�v��']MG�El�AgW��<���L��m�o\���
'6�i�>
g%���y�?r���U_"XQ�%�]@�R��2Z��t�Վ[M�{���D���;���-2�і�+ν�tHw��l���*������>7|\�Q\�Uǳql�]��P	��R��ߙ��8�+���_����ֶr���o���c	��!u��r^�]��1����^����sR�z/���ډs�#cz�i�4�7=@�z���@§��'�~>w���X�P�G����0� �/dx�j
1f"���T5���j���/������fM��b����d�Gs:֝���O��c4���߯�鉤��*�W��(�ͼu)��.�Y<�NRf�|���X��徤�<0�z���P�д���s��#�LE�+;��|���*����r"g8tM��
�Q(4B!@P�
o3y��%oi�������W��e@���p�(���}lKn��8�x��bD�4IaH�'StB�Z��^�)ݘ�����%�Z}�P%�_K�TMǣ��yLO�e���\�,Op�R���4�U��}�硠��A��CAt^����5P��a�F�QiN�:}~n�؍gJ�룻���C]O�����f����X��1/^�-��2 ��5��"��_+O�T�cw�-ޟ!�=b4��X�;kƿyt�� ��a}�GQ���o�$���%��^Ζ��s5�!��W�����[���&8#���O2����������~�|3�X���<h�Ѐ-*�6M��V03�� ^G)���M	�]�Px�չۦD ����r]y�x?�M"8�����B��3Sqqۮ/������f��A�<�o��N�A�x�5�f������y�ba�]��V�o��ˆ�uR)��}d*����ʁ2%����Ӂ[�wD�#���4��Khk �R�`o�3���ٸ%��|)�O-V���ۨ]��8mn�湀N�8��^��)�e91�����i���8�*:p��E�P]��q�$��'h;�1�Z�M�f�<�r��%_
}"Y���Ò�O���t�Yhn��E����3����m)6A�����}����>{���?�G���9�iT��M�piU(Pf�f�3{�f Qm����w-k��3<�^�4�`�\mtK��f�^����y��U���	nyNpo6��l��]O1Ѧ�7����v���ɔ�`}�EM㋼[P�E�;.�-�j-���_¶�4on�x�Aus��fԧA��#b|X�@�'6ؽz�(R9/�V��<�4����I��̴�T�n(�naS�;u��w��w�~F�~k6>�P�:?s�Q��Hݍ�I�ɍ���R�(��t�ln�>Ν�;K��>��^Ӧ�7�(Ei��g�����T���G�j-�������Q�q��F��yz�C�۞_XC�짂�o>���y�f���1�=�ʮ`�(�+�?�z�3�S��ŭX�@>?�yC��%�%�?<<��-��O��~���#B�(7�����V'�w#�j�ipw!˭�o�q�I8��})���S�@':�ƆWK_ç��b��𧾜/~JE�~'Z��7�viW����0)W��a҇y�^D�La`.�1<,�0<=􋬍zʟv0>���Rʶ-Q�#�܆��uޜV/D/�B3�}+�ۣ��s��_0U��)Kkw�~����Ai03�x��Գ
�X�oD
�V��YTǶ��6vl6z�M��ȳ�Շxek/*ͺ˛$�.Ź(�KmP}�3v��4��ِ���;�׮����~��<?������I� 5H�"g8t*� y���x7������(w��1��z�b��a��=�h���r�B�����N?K�8[���utN:gu�xg���T�3��?�
{f��6�/&q}l��#2�LSSs�]�B�:!�g�	
��A��(�*����u�ʼ~'����~��=n�ʦY9_��ܯ:Y�gy�X"���Xe@�H������u�#���p�E��؎~Y1�ʿ����5ѼOM���Y>�a�,�=ʛ3��!4J2*�+�c�y�b��Lߢ�tc�5�2�ş�oQF�c뙗-zDF�=:�c�!MHǅ���p��j�S�CL1y��_��a�n��l]�ܮ��V;7'̇�h��g'/�#�k���ͨ�l��	؄�8̱N��%u�5n��D'�h��:�4T�b���z\k����@����7g��W�T���������Ʒ��Z��3h��SlI����n���TǸ>��ڸ	�_t���W8���˚s��3���
1[˭�
"��Z1ͥB���@y���𽦃�0����Ҙ�(}��oߡ3V"����u�肽����7j��N������T6oS]�����u{;{ˠ�m�Ob�"ڶ���-��F4���tܤ�3�v]�[��s�ڦ�\���������6��(��.��v�{��i�KW4�29��j7l+�&��a4���a�~Q�i#*2a-��ʏ��94+9ˠi�B��!(�hQ)@=���~~�J~-�y��{�j�\�U�Q��q���j�>3ʿsk�~�=�'�+2���\�\�~6>�׾�=>�a������(%|�x��}����R6�U�c��V�[Nb�^��x��bC�~���CK�r�/-�"3����Ӭꅚ�5O���='��cL�Y͋ꡥ�cbC�/�/������T|V��`x�^=w�^���i�N��sM�u2���+�Z�C6>;���CozY���-�1�A�uV,>��ڂ����w��U�HS�4�Y�G3?V*�K����b��P���_�'�O�2����yEc�ec���E���.m������#�_����o��m�?*�SU%��m}-�O��l��r��_h�p#0���sG�� g5*� �L;
d����OC��T�	��U��i.�i r�w��+�%J@���9�ҭ�:��mv����>��l�x�e3k�������v���]7��$��o:�C=�ls�>}R)��C�j{�
����Z��1k�d��تmT��e&pUCe���w��|�W�
3����k��)��/M:�ݱ(P�c�*y)����׎'b����
c�R��Lz�Fq�cG��u�5u��j�3Q'���fwq���A��q �&�q���}|�����P���s���(hs��	@!s�����W^RwK��yo�����Aޚ�1��]��>,V1�j~�X�}�~�h��y�G�{9��b�{^;"�kqY��6/�#y�.]����* ]"�}��0ǝa�\�,*g|���F�W#R��̶�#�7g�(�n6���Ul5������{a'�W��'�� ����=���˔�h	�j�
	�"��������O����L�;�������k0wU��!g�/yo�t"}|����-3�V�.ټ�H�7(����|WFC�d��[��y�_�s��t�S����Dq���8�xE�q�d�盕"��>��u�	�X�d�8b|��f�U��2/76X���wwd,��a~�ԃi�Р���T%�:Ot��.�л��7���0ه-���6�[ҳ�z��Y�zO��3��d�����I��������{U|�tg��ʎۈ0^�^�{�Z����W�-�:��>���;�j�|W�"��� e�F�ߠ��_Z�u�9�N(�
#r��~�ף#�u�Pp,��L������'�8#��J���D�� �̙���}����niі��d2w1]�VQ�z�(%�ݻ�Ae��,p�GY�I���X�Í|��_��"'rHF�xzi�1�r��[+:G�B�e[�-��:��Wϸ	|��5u��<��oK`���r������F�D��ޯU���t	9���&��()���v�y��zT,�g~K�����H|e"�������b-��m�%�q�a�*��b)�=s˾���O�u��n�fc��8����r}8���g��`C�b�(Rޏ?
#������Բ�!��rv����d���җ�����3��/�N�a@���)�^�ŵ]��0�c����Qa�`Mb-�u�n�O�K�m�=1zk!�C��}�c���{5%���XRQM~�6�*ф[����3��k(�����T�����f��ۋ%�:��uy�)����S���t�+׹P�7gX��^9�����^�Ȣ���W��v��fUŷN� ��tU�g/�޵�GuUV�-��g-�sg��ln=���!�]Jl:g��կJ�q����[�0�fڥ�w(��N��A����l��pИ�l��x3@�ރ���&]>��E�(���_�`�Ƙk\�gVen2��71�#�Ν�cX���\�lL��2�N�In/�*V�M����b�h5X����5�E�
�Ib'�ڌ|w���2�ic�������k��f�h�ֽe+�;)�4�f<��w]0��:�I�ŽY�<S��I�}�����}���oۮ�:C� P�({�Q#����P��>�\�snT6�lڝ��"�
���W�;���e�]n�v�G%9kx%Nb/krvHs���߻�?����M�!�s�s�&���) �`B��_�y[$a��r��q�<�2�Ɠ&�B�Q�|C+ߜ%�=_��6���F��nf�u>CV�ݸQ\e��u��͌NS�����,%k=N�x�6����<A1|���~ٴ��uU�5���*�#�x����ᗗ?c2�-�~�]=}���ƨ;���<4?w��Czʬx��{�ݓ �g>t*��8�" ^7� 8��x�.�
��e +|�߻��2+��6k��15�o������G)"qP_}��ʿ����V���\h$-��,GX�ʻ��oF��6���]��.b��h�}�gp�����>�ߑ�\�^|iկe���aԄ�"���Myr��Q�`��֓m	�=��q�hJ���6�r|�%�T
y��QcOJғ4U8�N�V9�Tf��d_��(m������*B�cAA���p����e�[%�C�<\r���l|,��S�)�CR	�lS\�wO�M�%�z�e����7�+������<�I`D��?
���9��6�Ww]T�Y�:&5z�g�7�6:�ia�����%�S���J��\bʈu�3����ӴΦ_�B̈-7T�w60"Օ��n�s�m��>rY����eu5����\��6*� yƻj`��Sn�#Z���S�u6�Vsb�\���څ`i�jVR�k��3��`���Wrs�:�!2E�C	��O��Y�h�ot���1*��k�w8��%d��pX�zq�QF	��OCY/����+�_u����7^佼�橵��YH��Ky�I�>8��!�K��p,�B�x���|'>aF�ͫ��*.+h[�_k��\��otk�|��kw*LSkX��x��h	��\�;��jn r�t#A�Y�6.�|m�n.�Y�8f�
��v�,U��B�tQCύ�-�U{�,���M���z��2�(b�̼��T��s?.o@�ɚ������z��	���E���ݠ���]]��x�`r��!�k��억�9���50f���t���-�s��y�b�L,��k�\��p,u�6W[��#]��v�[;w-C`�B�7�:Tj�v6�l�,_��s���V�;��Q�$)�3b%Ƹ48S�:�N9������Dt.�h��gK.�3��j��%.�󚺄����sC���jV����9��7u�:��C[�m��$�:�]���{u��$Ύs�Y-�κ�h����( ����u���G�Y`nTb:mD��V�z<e�e�p��]�� ��!Ip�~yuٕ'����߅$����o��[���"(M��u�4�:"�H�:6'�T2��J]��v�n�";ٔe�tZ�o;D;6�p�zZެ�o�%��%:���ԟjt�꼩0<��:8.*J�X�C�^-p��h{��
�,WX��Tr������Ζ���{�BT����qq���%��]��M�*���J���zn�
�����7�+k�Y�c׬Μ�1|��Ķ�&wT��ە!����-�w
�c]��u�{.ۜ �`�Vحv�Ǒ�l�	��b�Md�񙥩�u��ute���)��ܘ��bc�0*�t��|`J��,���6�Sf�^�}ָ�w.8����0�����%�QbV�.򞝬�î0��lTd����^k�6k�>���3��WL;��oH\F[��2���+�[9^�v��k���c��:S���wi�D��D�p��ůMLś�^8��q���U���V����"�f���7EȺ�c�3/�^5�c�J���+���u�Q��7��ݖ�p��qYU��IǺ�Z�7v�2
隦&����r�5�����zWAbgL���I.���6��Yz/���Q��jg36�f�'v>�u���M㦬7���ꋔ޵F�i����YU�Z�#����s#�Y�į
��Q��ܦ���0K��4���-��Uz�(m�DA:�T� ���&�xnF�R&ڦQQ\�U�&''���N*�C�*L0R�2F�J)�� H?�7[��EG6�Y�ڊ��ъ��lD�TTT�UE[m���)�|z�~��_���~�_�������~b"���EAS�ǚ�DVƢ��+VE��;�>���������?_������??�I��ִ
�%���h֊�f���(���-�UQQ��*�<s�ׯ^�~�������~���1ETUDUl��0yI�C3E��[MM1i���ׯ��_������~�_������MMU��T��f�'o""�lTM3U�T�DEI@k3^�
�M%5QLUTME�UP�ąVڨ"���QUG��TT�3AE1�f�*h����+1UF�DQIP�TKQ4F��F�D5[�*������)�����j"��"^�<�(�*���Z*��m;8�
�	(�j�X>l�UMr9yPUELEMPZĔD�E[��/��7�<9g(`� D����u�	.MklQG��s�y�0(96�$��Fc�3�ˠ}.��{�"���u�jpӹ.\g{$�&�=�"��w?�_��9�'8�$�)�Y�������Ō.V ��
��/HA)׺��@��hg0�a�#|j����,ټ���sUi}C�A6z���ɻ�l�FbU�|Q�*����s��y*�~<O/�HY�BӞ~w��\��Ό�i����'���������U?\�����^�TG��GM��o��!��Ž������F+�ѷ����%����|IJ���0��1[E��K��2��zx���2N��w*l)*���3��䧓�uجsש�u�zkmL3����\;�o]Y�گ"r�5J�l�8ˮ�L��Α2�]ӭ|��p	G7Symz�*�ޅM2�o[{�A�K�(�heAM�Ǐy��A�Y� ��7���x�͔s��營���L��Ҳ�ýܷ]u�3��M	;�v�����
����?9��O��0�����z[F�d�إ/���ҝ��b_���x��|:�����[��^�(�1T"�IaP��o�L�����#C�%�Tyk��5��L�ùC��x>��'�7�y��7`���9��DE?�a��i��#k��!�ľPipu��H|������h�涂�,������6�M5{�3��%'�[E�]hj���Y�"�P�#"�����8�7�:��_�;���:�i�>J���b�W�TI=�0Dֻ�V�99��;��}wUWT���9S9��9�:) f�f�-B]X�M>�
�P歑��@���	��!ʧ�<����?"Q�@�(�>��~�C3���\�߈x|j(^0�&�fC�%Y�|���iJ�G{�^�^�]���'z��r��˶9�� Z΃��;;�r'=��\[��?����L����]O]C��v��܀~tp������fg��[�`{Q"��	k����]@��[�!�Y�ĵy:v�e���c++7�^aWRַ�;�.�g����W� _89��~^�"^�U(�Yg^�wb0�#��e�7�;�8�lj-��q�.�-����׶Ю�Uò���1MmP�)���lC�Zv��z�>��}v�̷�2FZ19��~C��X�
�������k#q�ɂ'��~k�
N�~Su�e��L2���)��f�c�����3HT�WDLY��O�G�89��nFѹ�7`@�����P����j�B����!�a�����g��xd�}�|�Y��R��x�y.��l���r�wK-�$���D(Ù�&N q�!�j�a�'��t�y�ڿ5��q�����z�)��fBv��w\����%-
�JͿ;����w!m̦��]v��Y�������2vlj  ;X�
j,�[��؊�O������=�r��ᜟ<c6]3-	w�/O:�noMGS,-��k��fض�ӓ���H�铪.�stb��>;F?�JO��43���G9ƅii
R�����{���_�X��O�=�������	\����~��+��������<�;{��9Z�\+//P���h3�<�.�*�X�6�r���=���M�`��7�:���4��!%vo�"L+�a�I6���-��H��g�=�,z��;/ʇ�KG���O$bϠ5�D�R���Ya�{�t~��Sr݀��l�?�k���˞�"8#��D�D��-yMgS��Լq�n8�|Μh�}A�
Qt/�G�K� �U�{|��{+J��3 ����So�E6I��}���.���^Ľ^	�,-��㸻Ɂ�_��iq�⼜���P%��[E�ySt��`���f%�%Vf��<��0�N�W�#��2Уw.���e����g����ɇj�ד�l'9�.�4�(�D�;�6���m	�NE�_�}?Yܘ%�^�iĝ ��
]N��j]������І�)��-�j��Z��mz�b��v8ύ�:3`�%�q�"j}-p��ۜ��0�����lD�]�M�]o)���Пx{X%7�.��[p�c)�l���5�UN�-��5+C����%1#�ZfQϮ$���ο��v���w1[��E,��uF��/;��,%�E���d��(�4�*�O���K�������3��J�Z<+]��O.0��>�W�j����%G푳A��� ;�Oϟ;���G�=�����/�٢��8�Nv��s�Q%B����X��&S���[��@,��=���y�70pQ���4>(ߒ�6s�~i�o��&k���a�|{�
��~����~��C@��=����l�o�9ye��G�c]�`�W4L���d_C��L�e �x�����9F9F͖��hb}щ��σϷ�0���^_o�+{[z[���Z�I�\+q��������s�nᦝ����2n.��t�t�AP�����9���=cpL\%��i�}�ƾ��D�����m%��������n+��{DA*���,����U
����UTG>5������u��ٷ�ݴPg��!6wwqD�֩�'���@�[5
����ym��-~oEH��}�X� �Cޡ�~��L�&�^D�����c�eټ���&��C�~"5���Q���!iůԅޞ9~|U�=M����W{��zy�h܀��3g;�c���Zd���������b$[E��ϓ��gsoN��.����-���5��3�P+W�ԑ�}��_��<����7�����y����eW��-T��G�/!U���XY��_9[��N�ֲ�6�f̋��lj�� �2� ݞ�=��'eJ�v:�H��]�6��yL\�`�Hk�ru�	mF��w�js�)�޾Kwd���	<ˡ+I}orوۺb�Ϝ�m�p��?Ӑ�r�8�Ns�K˚��~�������yU�j�����g���+�-#�)�TKE��w�z���k�`쨩>i���.����x������p�i6������~b��;^���0\�Kh)�;�e�D��2�8v���1̱k���r��Oe�:�K�Z�\l��l�8Bh�L�ʹ-�{^���j�!�����Nݘ܋����2��<��KH�a��@JEϹ�B�jlK�ȖJ�Vܳ3@�6�Uv,����pD,�
�~���?�� hD�6o��
����8������U<���eSSe��f�a��X�?]b-k�X�K��
���k���]z &Ɵ}G(7���jL=5-���r�t�s�E�/�[R@m�4�B��J&q�^ˋj�{��QS�w�M�.h�03�Љ���HvB�v�'�����{1�ʎm�T�~k���_�����"I�ֱ}Yu�$�{ş�u=��V�D���)1�@����^!��O7��~4&x�yW'�Ds���;k�J._��~w���2滃6��ޖ�fod�
V[�|5n����x��P�!۟�3-�-L4��ol�s�4%��jVu]��L~K�s�:������T�ĺ�Z��QI�:��<jVg]m~���<>̂B#&gdO�=�4����F)/�s՚����}�_������)Q��_NA�����u��R<�x���A԰�,�.�X���ԥzd��r��{�����O��v�s���������A�d3_���H����>�x��/<顡����ޚj��U�n͎m1���w�H��]Y�^-�����+�A�"
>�����
5��<r~��W�Y� ���w�V�ҩ���A���ίPL3�fw���W羨Z�W������#�y��'.�M����r���^Qp��}ޖ�[eX�A�ķ2s� ���"Kሰ�(kH��d��B��Jߟ|��?i�'$M�vJ��sz��ve۹��p2@;_���Ŏ�����nO7��&g�P��j����R��Gd���ǣW{g��SƲ��O�]����*D��Cw��̻i��A�çUWbfX�=���go�iEZ
c�%wɉ�mU��y��O�u���x�xd�(�fU^Z��NPn������G���|Ȝ��$�ҨG;�☵lQ�_[LA%�-�>��mC�Av�5�!����0xۭ{I�Z��}�!Ͻ�T3�m3 |C~t�y�K�����)�y�\{$u_�]����7;���u����z��i����M��Qm��캽�>�0��T[1������H}bϺ]v$]���Lf����Qb��9��x�h������p�B	з�Yǁ�ke>+�Z��6w�h.�y�~�5˫�%\}�{����5A���Ou^q
�IA�r�l��B%-:�bj���w?���|����q�͈3`���EP��KPUVߌc݃μ���ϣTB~2���Z�a�H�Lcϴ�����_���hɽ��3��b�e}�g}�?��Y<U�foE��
�V��@�c"�O�EP֟
F�|խ�2-�)�b�Je��2�՞l�`�y�m���C�3W�3�&��v���ݽr��׏%Ќ�6VӜG"��ݴ�*b^����Y��k'��� w�d�7��F�NU���2 �'��7��k;U�A��� b-�a=e�uπH0? ��/����KD�E�����c"�j�:Y�͉��Ng�b�l���vK9zv[�.��s�=�R�qkd00�:�_G}ιc�Dy�DŞ����7�Z�w��Md�}Π�r�q��躮�@�<��PAS�6C>�z*]h�/R2�;���v��s��d1U�j�u�X�=>]~�K�Z��zr�0��Pd����4s��f^ե����+�Kk����/6�{p���ć�V�֜�Ə5�m�� �J`�q��΃u�WR.L�����yw��5�>)�4����)�7�UC�6�_���U���Lu���[�y����o!4N���۝:YkGH}v���]���[k�Z�n�9��gn
��iwȣi���O���nu����oka��n�v�8.;��3�g60M@u�Z*���dx-�{��U�Z8�3�.��k;;/V�\�sS�)�����;S��;R������}����벦o����~�?��7TH��y�D���ʀ��7Hmy�x퓧.��.���Kl?s�9=ב����p�}��hD{!�R*�,��^֚e��S:���u3��v�~o�&-�}>�*yT�7"o|��_\̼���c����}�8tG�ü���5lX�v��5��Ol:Ƽ&��Lq��S��v��x���8����]�o{��}SeF�w��3�����s�w���+1���U}0����	=a3��v�؋W�j	���M\�j$Dl�+��Λ�^�Fj�j�9e��D=�і����rzb�s��	��s3FM�ё�X� �v{,����Cb&��p���X���߽AW��:��Y�3�'s��syH��n���e��尅ұ�*a��kּ�q�/	��m�Ƃ�+m�zb��/2�!v��εĄ�V��d�,xw��wj�8|8�*�?,"t��6}�$[��!*�X�=��0fi���0Q�M��1���gaӔ��8�&K	Z�:Շ��#jC�8n{�?@W�>�w�5�O;g��h,��{f�b]SAa\�ru�\��V��G.��k�c�5�tO��A�Lo� #�D6Bh#%��qx�VA�>�gF�Fд-Z�����d����;@�������J�ͷ�E`evss6�dNz�G�D�0QQ��4np��1ȹ�?��3s���`�|�ոA'�����^����e����؊�|cLd�8�����bض��F8���S���Jp�g�g�),������Q��Џ����O�����|��Or!O36`�j��ٗWu^AY�0�Y��>����������2{�����x�HS[���g:ʻ����+]b�l�;��}��ЦL�]A����L2����Ʀ�|��P���`�4�����ɢ�3sL�o�C��(M�r�a�r!_)ѥ����V`��mT}a��c��n��d\[�����j"!�k�{���42�m;�L�64sԜ�����4v���`����C��"�T�Sg1`���A�	�r�cߗcȟb��{�����:`{bk/S��'�w���1�
�*���u��//z���} Y�/���h*�y�ӷP�L�DK^�~��0�zP�����KH���tL�]魧���ӄ�I�A����Be��SP��p��O
�t�X��-���ֽ��P	Fd@�ƅ�gv'X�"li[lи����RC�+aO�m�ߖ�3w����P^��ẛ��J�^�7}]i��� ��^~�_�v�7�D��=�0��t����gj�J�E�U�AU
B�_�����>���ᬝ�:98�tV�./;�K���j�} �t�*�m�Wl�AB���Z��S2�*�V�\�=z���5�?������߿��۝�|�^s&9�̈́�ǱAol��m�Sm�э��\[T��D�#��"&܄�eTB��i^Uh��~��2䇟a��qΣ�ǌD'�EG6��q�	ñ �g��?�S�5r(v���5o��!&JUk�c̄�6����t��H��28�%��s-�bF�ЛI�5;s.���\�+d��{�W�^}߉���1��!���ʐ��KU��n�RQ�ܺ\&p�U��R�H-����6�3��NL3���44d.��2���&\_Yӡ�J43���Ӭꄾ�A��2`��f8�b$��y����=�>�{���� �����l
��[����/�\���w�|���X����T�W���n�~�n��v���F�GU����P����Vs�ok��䚤]�-i�P��F�0�O�K���nyy*���9�L�`�,�����_U��N�x~fg��\f� V;6,ɏ4y�ي�m�����E��o�P0^�N��A�ZjKC�� ���q;��59L΢����>��8��,��(-q|d.r#���;�5��a�s�wN/�Ԏ�;��]��YOz�+}m�T\��++��ʷ|�XW�!mR�!�	����pI|�-Y��h������F�5�fG8������r�3S{� N�I
ф`�����h�e!ۈӜv�У�/X�.���.�W|3GK�k�Zz�9
LְmE֫�Kb��W��a��0R�#Q��2�3%��cZ�c��傗'F6������]����i�9�LŌ^QB�a�.�Z���W�u�L�+jc�"�9ٖ�P'�֞5BRk���;"T����Gc�th�B��/*.���7t%���`Z�Uo�gF�9"x���Fa�p���h��WR�3�0��3R�a�Tҭ��;�J�y�B�7%('֋����q��A�#Y���VR��|&�O�,�v&��ke�Ȝ����T#���T˫��:̘��EbT�$S�b<GU�ۂ�F6��u��<�#Zx��~�\r��UQ�uj�H.���9J����VZ�fĿF��AM �(m�/�N���)U�=�a�TНک�u�2�Bc�ף�}\G�~��᥏�X{��б�h�Z�=ZkN��*q�Ѡ
�VmYz&*�h{���q����4�7��f��(9}��g]t�X�VX�� tK}a���ֶ���ӜցD1tj���/%���u1P�ʳ�zGR�i]\S�G0*�<�\+hh�3�ʻx�� Z�x�)qrh��^��w��f�n�bt��.��h��x��,p3�M��[يb���ܵX?��}���<ɸs̋{�ެ��V���y
,�m��R@�Ov�]X.�X�8�k��\;�K6��Y�Y�ռ�/-�g(�5��LQ���fA/c�l
0Pe��<��T�2� >im�"n��2�=��ǂq�-�[B�47�)u<����|�>�4s;t�2,U�F���i��`5ܻ�aq����nN��#�L�th��� ��ۛ*fLĚ�\x��Y �u�Ƹ�RY"&�Û8�FG&�&����4�׹�A���6g@��:0��[�QZʎ�{Ԕ��ۗ�dU���l�˷0><�*�	��ǁqwW�!У���P�Y+�.��޹����ӊE�Ј�H�Ş̒��E���3z�ʋ)پ�W>�7b �s�<�r���D��dT���S�eu��wh��,ې��vz�_$4@/UY��T�MI�`� ݷZ�f���g��%zH"�!Wnn�w��Ü��^�ȵ�oo����a�3B�X~�F�B&�p7��t�1�V�����e.5F�m^a�X��mM=�X���2�P�f7,��ȴ�����	��5�3j��z�'{X��&�C�[���ծa�ŧ��#�%�A�H,�%GmPLSTPDT��C�Oׯׯ�������~�_��������((�$���Gc�QX��)��D�4c3��ǯ^�~�_������~����~����f�*������툢��U�ԑM��7�TL�����ׯ�����~�_�����~����t��������TQDEQCAA���)�><z�������~�_�������������AD�QRD�URQ5W�1�/X�AKI|�"����<�51UV�+cMD�b�**���̀�:j��&�� ��#�43W̚����j*���j��h�*(����`�AL�ED�13̚b��Q$�$DA�()�f�I��c1US͓�h��
�9�Uy�<����
o6�UERET�Urt��t������}�;����t�U�^n��#�����;�C57I�S� H�k��,�(Y���ϫ�_�~_'>\vݝZ��/�j��1U4��/SP=R*)���{�t�y���d��#�c�9�r�e1b�CZn�����5;�}����D�>�������e��s�z��Z�K=�Z�ݽȺ;o������%D0k�y^_(�|l�6\�3q4b�7F��9��cmwj=��ɜ��>ϝS�y.�["�)Y���@B���T�|c��wCAИ��p���Ǣ�����k�7P^�A���u������e'��7+���j���"v��{���K8)>��>���JB�m�.o{'��^y��f�/�3FRU�`d���w�]�c<��eP�F�l]��aJ�mf���b����G�����^ C�>�!����=zɗl��:k�{|^'˔Y��
�D��R\:!��6 �X�OT��������=���T)x�+ ���ZEto>g��I�g8����C9��[X�ǹ��C�Z�"2|aP�y���w���o�1�t���a\�y�fV\��z��Ξ�G��3�>9N?p'�yE#������������VÞ�[�u�ns���"U�#�_b���W���u5��P�4��n��}�2(��ah�׻��ӻ�݆�DQ��ir��:�wj�2�����q�J�c9;����͒����k�Z���<���)t=L�y�S�ZhU~��o7����{�ONv��l���S���`X����U�C�i�S
�&Gw��<�.���Ϭ�ͅ؎m�qOHnr�������>��3>[����T5�>��Cz=�g�Hg���4=9N(C�}U�#�D~̽�}�W�H�t��i�	�i�e���ό�(/�~����:�����68�q�a����s*���[��.�s,��&7�%�4�Ϡo�/�Gg�ߟh_���;��+�����������V���>�5��ͦ$Cμ��"c!'�Zh��{����r�|D��ec�|"<��.[a��t
Ayր�Cd�ɸw���5u��=��佨}�鴦D��4N_�ihѣJg'F��T��q'b�}��yq	��=�+>�CR��Z� Ό�6o屌�j����̎٘To���+��"�(�~o&��Lu�nE'V�hmUf��v]����9�ѹ�f/K���y����}�W��b}4�׸����k=�⸅�/]�Y�dF��y�ۺ���}L�9����;�l|�s�8�W�2����]��s������S�����;C?_�?mgU�+��+e�ɡWK��o��hv0�)� Ю�P��;Vܙv��}�*�=P�ֈ�t����ڮ򃄥�k�R����
K�Q���1�h�l��+�ː>�H��		6����4#�4�cͷ�{�s[_(X��	�W�y^��~o?&�I���aZ)~I�L47�: 1��}���s������rW��<���`���=��sn�5�'�"���>��>+{�gq\Ȱ���~y�~|sؒ�����p�z����q?����-�1|q�4-�T$�f�9�������Ӟd�n��������-��co��]�c'aN��okŇD	�K�f<b�Ŗ�z"19�l����aT*�v��������S����H|9��.SJ߄5>1ܭ[�Q����y�X_��9�穘�З�R#$��%P�=/oۅć�3-�)�b�������uM��,�{��'������D@��}W(�ʄ}�T��ʉ�Z�p�#_�ߞ�cf��3��C>;v��gP��_��s��B�o��#מ@2@�a.g������_?z^|{�������n�磘S7�^�B�Y�|���
�=��dD(�r�iǄ���>+_�-�c���i��ך�E���[q���WOg��'�'�R�=�E�����oC\sxD���
����6��
j;2/*+�|�dS`d���9�ʫ�����p�8�C	�몗��'�;����,\C	Ab��W���3
�{�V�$�����9縚��e�R�ʏ~߈4�(�y�Y=����%�E 8�g�kZ��Vؓ	6�;��gR0{���9᛫v�i�r�F2����R[cP���$���sh~����~���bAv����F9��	��YY^!�E"�G(R��z;DN=�n횁oyw�O�/�m|5RXf2+�Æ�#~��Ȇ�����9�lN��<2ZWT��)�ϿpMs�����}�%IK7"E�L��?l������%����ϑ�L.'�f�~�"f+wy��E��L�A�m�*�`��DxU���a�MI�e��kV?�U���[��v]YK�!��:@y�9.��]0�?�7qSM��k��A�l����p�E�Ǎ�f�A��i�x�![J`�د4f��q^x��I�撠��)P��xm�r�N�1��ka�m����gS^��p����_}�b����t���zE�4"����G2~����뗕 �0V/�{
���=�3��(>ׇ���,vuRc8*e�E�����/�P��u�w�5kr������eU` ��d-e��C�H�B��B^y�/_�)��LKn�k�*�Q���7=7�G0�f��������?�j{1C߆1���laao�~>���Y���)�Y�w����+p_�L?ɖ�U{�����-t��KjO���ۦ��c�EVI����X����l���KZ���҈P��1T���`�g�\��U��UM�w� �Ji&��ro�������+;'y�y��Aj9���ƌ'�)�߾��������(��a��KA�si������p󃪃y���-�\��ݛ PXL>#R��w�D�K�����c��7ӆW��7@�֧���{nFy���F�m�p�=ۋ��B��5+V�#.gv^��֎�p�f�"������Q�>3x��s��M�:�4Y�Xz��1'6�U�T�]����5ɂ��a0�,�se�?y��fD��Pſ��g��Wy� ���}��I��l�����|��'{Bb{�w�`=c
�)�j=SQL�>���/2�h5�sk�Uv?v������co��;�`q�!ىW�4t]B���` q�?���y\quO��ٻT�fwf��f��WN������^ω��ʦĮCN�\<w���߾�����6Ћ�4�����}���iCY�7���1�AdQt���Jo��NC���e��u%d�J{���6���"�CO>0��=>jJU��	���y�8xgp3Xś;ҚKpR].�P�t��Sx������&�C�d�^��s���|��mw�qzOY���d�՜�o����rw�+Tqxmm\te���`gd�3���e���\=�i[[Y�b����7�If�iF��L�{I�]Á�p@��aG�g� Q��B��Î��q 唦��ũ�^c37��r
69p�HۮV��ѐ�c��^X���ʖ�T�E��b+�x>t���30M����s�۝�?s������Ѯ��^{��2�W�){\�O̚��l���4��ΰT����ĭ�s^J�'��<Fy���a7kNr����q����k��6�!?��*=�ɿ�r���[������#d�\�W���j��	T���y����x�G��}弲)�ΚM��n��W`�ޣL�*EP���V�Z3���=~���_h���;��3@m��=f��&.��n���v���R���_E�T+�S�������fu�q��-C0hh뺆F'�*q3x=�?�^���� UjD�1l-��o���7����]Ӭ2����$�DR�3ut�>���x�q�~[�`�t�+U�X���E�5�]��{z�gZ�?OZ�{@��V_D��Xd�8��b���ix�y[��ؤT(�𸘶��*0O��ی>�c�S,U�5}��y��_>��=�O^%�٥+��|\U˫mM�f�zez�zv:�X��݅Y�.�!Uv��Z&]�P��ao��k]����� 쩿�~������o7��&.���m��K%>�.20p�F�k�}+&9�*�M�������*@io�Q;,�.5�_Ƴmo+g��໣f�t�e"����-�e� E�>2���h["r��t��u�C��b�"�4���a�Ύ�5l�k����z�򹬨�m@�Uc�6���s���ny�:����[�z�ޔw�ox�=���~�5�.)Vrb�܆�y�Ɖ�����5W1=P�0f8������,X�e>dN�n�B��,nL뗣�#�W��#\t{�SW�1��3�1��yO�.Fr���/r�ݴO]�1��0�fò�^q�4�'�nUu�`$t�s��8ϱ�����'z���)fU6��3�վO�1[_�����۹�� i��Rb�xf�$3X�73vs�,u���4���1w1�*_|�m����^����S�Q+�)�f�Cld�g"�W �zKԦ���e67��nN��hh��a�E_䇘����ož������Eoނ�Ʋ�<��g�H�^�׼\j�a�M2`h�,�ýj)��s�׼[�T�f����o���0�Zڥ���j���r�0g����T=�O8�ge�ג�>07=t�QaK�癭�0��֭EE��[fx3a&��ƍ�`a�o�|�]���<�ޜ�g��f�����7�2��ce�P,�U�M�W�����f��Ͱ�J�g�ͧ6i�H���<��	q�9l�V�/p������1E����4�Va���	�:�`uۧhN��nLA[{#Bq9]z�L�n���*y���:p��,&�,@�q�'�k%���]�ƫ���uI�PM�:J}��uw��Y#,�'h�6��.�b�iؓ�>V����h-�݌U_���������7��֝ri��f�nW�Y��\q��Ø'<�F�k����U�#�¾����������Mrc���^y�Xש@c>[�q;�]}�����L��佖�dD�P��R��i@(Wwh~��mѨr�-ݪ�S�S�����������l�z�}@P�c�2�A���Q즣��5D�QR�	|��
��Zȱ�'���r�ж81�X�iz*=��K^�6�y-��*q�ߞ��B%��C9ji�\-u,��lcئa�$�	��6���sS�n��h�r���c�!�%{�#�],�B��w��?q?�5Z�.�^Y�qԻ��k#�k77�Ƈ�#�?����{��X�W1��ڞD �n�M���1�%�׵�^cl��l��d�sWG=s`�An�=T�=��l���BQ�/�F�p�MH��@M�uM=��S�o?%��z�Ձ���=�	�	T���U[mZ�+��Ld>6����
Y�^���\o�n�:G߼%�c+��J8��gK���i��o>G����ֵjC���J4S��<l�����A�ϻ�F,��\�^���p.��P%T�&�ۦ�ӵ+R������� U�dk�9�Bͩ$/��<�]����%[�-l��/9!6#Vi�����N�Δ��F�(�mEg�c)ͱ��e[���;�y�o|�7���,��Rd���^�iOj��?AWc��(;�'������Ns���Y�ى��{�ْl�2���=���t�Ė��~+�C�"|D������w�
4��Ƈ!���CO�a�!5w��y��uS��ݔ@��26��3l�(v���������,����<��y)f�(��͋`��k��;ӭ#�5�Aé4���<��"�y.�ņ4@O&4͚e�G~�:r�e�ְWΣ k7?k�{zO�[P��2(�z?w��|o�)B�������=���o�4�:=+�`/H�I������-Ŷ6��g�{ɒA�T7���]�%@�/X6�m�a��i�A~L�)ò��MR㊊�f(��������w4
��%�֮ˍ�kÂ)Ln,�5c?o�zw�u�p�/�e�Ň_����~�N���"WKI7^�b|eY����%��9�d�C��/^.ͥ�F���o��_Ӟ=x��n��)�zۓ\�.j��Ǜ��M�))>N��k��Au�0�ZJqdϋ��U_��t�]�Y���C�I���{*�̃���y�j��`�gs�{_����ox\��N��("X᥋��������oq�1��=�<眂h�1O#E;�<|1��t�B35l��N�����[j᧹�t��^J��^RG�p���&�����j��BR:��:Ŷ�X#K8ٻ/0��y��g�6t�4I�#���{\���Z٦L�V�6�W"dZ����s�ъw���#U	w9�q�������SF�c�] �V@���+z�Lu�tQtv���/i靦��Ӱb�n��0���i�p����F ��d[�J�8���8�+x��`��C�Z�a��eu%BBݪO��V��p�s>���7����7�i��\Dsa���%�5(����y��l^��Zs��Wb�Y�o�X;	�b��/by��
��A\hbg�+�ߩ�{
����rĭ��H���'��x�=:_�_}�MQȰ�1S��ʣ��Y"z]�i�ތ͛U����Z�b='��\�%n�c�(�'$v3������p�)�m�;5J�����â�f�q��fN�<��z|�^��t8ї�̀=����x�μ�]��8?�UoK�d�}W��*�{L��l1��5���ۭs۫0�N�{4�KF*���1n�d����Z���΃冧׈�u��/���Ͼ���w|!3�'BD4g7}��R0Jݱ�r}`�[OZU@^�SJY���,[������=�8��1'
�Ǖ�a�e]�(��h��U����`cJ����;,LeVRx;��w(�h!�}��]���s�|]�+�c����%qf�.f���]ݼ)S�Mi,��m�z�KH���]l/X%���{쿝��;��F4𹷠��Y+�:�L�{��w��L��e�J�>���+j����Ez��vP�u����	���띚�%%���ꂙވ�].pg^U^�;�QB�PIL��sC�pR_Z&�3Z���V�2�)��V�R��F6!�ڢ��dN��ݏtV�7W�X��6F{]��v�� ���]�hj#�p�+9�^j�45�0$ӛܲ�X�)-L�W#��;^���o����w/�ˮ;GV�7/�М��wws(�A�,i�{q	6����$���y��Ō��[{��Q*װt�9of|���.�������a
w��r���gE�P�}���1Yn.z����X�S�/���
l��d�n+ܽ��LXP��q�%a�iI�)]�0@�"Nb����r�7r%�I+3�2��{�VO;�x�A�k�ⷚ�j�7y��T[�[q\��d�z�93+2�0G��QJc�ueJT�^]��V�F��gJ�,�S��)�DKQ��CXQ5� �.+�=ķM�`�Zl�@*�eG-��@��/;tF�ZIڕ�˘Z�z�4_>kd��K8�hAvNG��SnR�2<�|����n����\ae�L ]�gI73J���۴ә;�=Y��t)afq��ڄ��'�p�:+z{xެ�����m��+�!�|e)cMY�ݲ�zinC���4�y][��'L�O�s�g:	��f�W�u���5����7#)�Z�|ew�����)pJ���S��(w7[�=��@w�-(���y�{)Ž����׫զ��.��X�G,��~��3@ZkRsU9*I䶚��p.��J�g9�1�kwv��;ydJ���Y[%s2���W7#E�<Mя���[��4¤�`�e����rN}��I�Zl�8q�'���em9�8+�݆�	����j�_ua�+]���������\Ct�I �2U,YIĮ�u�\�����e�뇂�E��c�zy�u�WWg�ai�[��(�ɕ%F@��j���T9�h���*T{�չ�Z�p�&�f�7�	��ɐ�f�M�B��d6zrT��gH�lR.�y���v]��Q��C�c����k9T�$��������I����%�!|�I���Kp]߮!�7�gI�P��"i�L%Ue�����A�Q�b�e?�BA�C�	d���ԁ8�th�we�X�#�y��7T�eR�ҽey��%�D�˸\�@�(6�ue[E�H�5+B:�%T)o�~i��uUE3A"pe�Z(��:j(*+ͨ���&|x�}�������O�����?���$�֍��)�h��2b��y�&�'�ǯ^��_������~�_�����jb����m8�(6�&�_lS��T�ǯ��^�_������~�_����)��ij��&���Ө�����qh
�׌����z�������?_���������#�N�(���T�Fڼ�Z*�#mA1	A�8�	�#��h���$F�5>�TE�3T��EQ44��PPzF��O$�5U����R�)��`�\�a�x�y�h�ד����h����"H��\�i��Jij������
�2�"�J��&�����)��cK�����
��'� 	�z����$^s׫d4)�����^�X�9]]���{(3��k����aǲm]�G�cotڗt{A���;���_�m��������o~?��.�O+2i�w]�"?>x��[��^hN�}`�e���-[�s{�٧{a�5���><��6�y��ǈΞ��gЯ��|�P�^=���CN4	�&ӪM���Z��R�Ii�i��dG��g�k'ώ��aܼ�Κ,�dgk17�s�k��W�;(�;w���G:��[+���Ī7�6"�R�}��k�׬�Q".�ˬ�k)Nb9Q!Jͦ��p�ov(��a>���M��:�Vty���Gj�R�V��c�9RL�.��U�l�??|"�r�+��u��]?,���X��C�8���_p]Y������x�t�Ֆ5O~{�3�og,������m�w�Y>�3�L�m^m���!Љ������=�]7�}�m��k��>��S�占�Z������[��k��:��t�4^Vb۩�L����Q���o�oo����Lպ��3WUjP)��Ȟ"hB��J�m�����A���Q%� X�_{5�<g̍�|YGjY\�k�R�Ӌ������PyS�Q=����X2�N:Tk��|5 �z}�_���.�B<F*_t�C�����r󭕜h}�xxxx7�����h��3]�ʱ>���o�d�tQ1GL�Rԑ!r�=��{��_�6�[-5b{7c�pA�)8�û��f�[���{��Ff�2'@�|V���s�sػ����^1��)��1���2�ɰ�u~O��Z�����2٠r���~!���G�{wUg����7��>��n��G�������ݶB<��xCn�ď+�y����'�Wɹ4y��ݔ{F�]8���
�b����y�{o�>���(a�q��(V�ư]��#�P�^��d_����{����cy��OC@��A��L�tE�g�g�vI�����k�����/p�v#P|>��������Q-�5RDi3�5B�P�/�"����>����f����y�=w���ْ��f�W�wT��J��׻	p����b�b�q�7�{v�{�7��{Փ��P�M��$U�fC��Wl�6V�������Λ������*/A���7���\r���_\rw#�DZ�]�o]~uŶ�Ql	����-W\�^�4k�Y���D�]Qs���{܈F��K���t	��O��cޫfɶ��o"�2�Ǐ&���{y����^o7�� �a�k8�1��1���{�%�w��@虲���V���=\tU�g�now�R�d�^��k�Í �l��I]���jbf[&own���Pc2-\�{����A�
@_���~%^��l�k����[p�v���l�+4D��X���>����R져J7e�-Y]�R�xp��T���bї7z'"K��;;�6S�w>�A�@�1�!�T%oO���EqF��10��k�/Ϲ�X��vm*��9�n�_޸��Bcb:�]-����u�o����$�<G�[�_,(p���~oF&�����|��&��xF�d���(޻��칢;z�
�c>�MS�`qi�^[�Co0).�xhM2ٸ#wW7Ci9����gZ�,`�\�m��>
�sh��j|�N�޼����/y�K�HE�0����]y�o�l� ��-!��h�Λw��\ڣ7&����Eu�Ҵ_/#�m��B��f̙l�9{�:�(|r��l�U�j��k��ߚtx��}O���t��M��ӻ��k��d s�.���9)ފ����B6'�Ћq&c�a����lv���w��o7�����}�|�~Q�]�[��v�����>:�u&���i��%7�/��']����[�y��3���O�.N��n�M��]�\u�=};t��3;]k����q,�0��(�k���dD�s"�x�Q��5��nhn�JHʯv�~��1r�2X���e���^rK�YX�Tر�Y�ʳ��g�}��ܧ\�=~j*��T9�f'��; +�ݧ9MݮD���=�~<]0�����=Ω��P���ZV��7
��a)]Ό���W�z���g[�o%����Y�5g_��Y-�����ö�Ֆۣ[=��mva���h��ǐ#�u�=|�{}VC���O�_-�[���и�nl]�m1���#w#��Y�I��#���7jWs+~���V�5Esv�n�'P���HH�xo;�N?��{��_�`յ1�ʟ���7ӛ���wp�9���aS8�8�jG��sn�X�"$G���j�O��t�0��v-�f��=kj2��W��WPw����M�d�D�5m쥑��I����Qt陊�4�єּ��X�u��4����~�zq�oO,{��=��	����y>^��^A���2��I���u|���]IQ]�ls������XvW�)��ׄ6ߨ��}q^ L��=Y�8ue_k.���\ ���k���9h��m�PX��.�i��Z���q<.k����*�\��=^{�T�5�����y��"C��7��HD0�=�.aF��V�q8�m79ƛ��Di���v��ǉ��ՈFsz6 :�o���2.�}^�w�Y�p��b{��=u3xV3�-w�!��O�@�W��g����W_��W�z�<z&���*z5
)��׍�z��W���g��/qg�W3���-N����6.f������������^v�D�sX�Yz��-GH��5��{�,w�>f�v}g{颫!�"D�h���)� U����>Y���
����=Kq+�.vx�5>����*6��~�m��P��*�M�X��c��*�w: K۷Y\X�n֗��LdvӍ��̫t��ḯ;i��&r�֮ۥ0%��]Obm�g{"�)��h��u�i_e�p�v1�@"ۖzRth�v���5eMu��zo	��XYK;��[���i�9���=�U�ͺ�P~�������xU3�J7��/U)M}�k�u7��^�=�����Q%b�{]��J���i��l~��/ѳ��7ˏi��ej�}Zs@�cR/�/~F��l��'�����>�3�f;)7orn��2�xג����Q�q��jj�Y������]���Ȝ�<L�wH�'�����ۅH�t�yYX�$MڅϮ8��q�5d�LZ�?OA�&��^ɁB�����GY�䒾��X�Z�6HWiV>��uv[V 6�}�H�*���љ�\j��ʁ;V�xs^����`x <����願���G�m7���6��2�#�����o���c�61=�[�ӲL��ٿ�=��%��*��ƕ�;LG�!���_`�(:w���]����#^{�%I/���\�=�h?H�l,6�.����oF
�q1٬��{% AP.�FU��~�bxْ�+a�ώ^	�6Dͣ����b��i=,U'�$p̙R�M���w��_����f�-Q78�/�6OR���N��d��X���A��e!��_8𽜙�׏,
�^e!�B��$i�+L�9����0Zr��[�c�zz�z�]�ߗ~����fvs3�^`'kw'u���ً;6/�g�9>m1��!u��s~*�ݘAL���k��{�ـ'�s�6n���_�/Le��8s��cQ���ۻ���vS����7��g%��5H�Y3�w<ɂ�`s���v��������9۵d�w*�z�,Ӽl��ݎS��ʹ}�o*���̺|ZO�ga)냊i$+d���G���}�>������u������E[�֬��5����y�YӍ�:��#�T�����dܓV�%��x�E�q��Q��?�&�hn�����voC����!�4�e���=�9s�@l�tQgl�ƶ��(�M+��a�����Z�/y�ڗLl8;��襋c��b�⽴R���B��+�o�?|Q�L�[N����[UJ�E�/ 7�]'�o��'�$�S9��!���{K��kv����%��ǌu�����՝,�c(Z��		�t�/ �t����P�l	�b��o�c���_,X��? ȩ��n)��q���r��I�ٟ_�ߔ9l�8��� ��,V�t+nG�O)��=�:$��d�kxu�l���b#Y9)�\�.{)i9����>��?����WZRN�*�{�<{���֭��Ԧ�����F���B���jub�zZu`�y3;��q�yK�;�M�G{6��|�F��j�܈v׉������~�l�5��i@��~s�����=v��ӱ�UV|�І|��h�aq�-n>���XLrN}��3U�+*���}s������+�;D����U�oD��8rzz_<�������U���j���fn0!ݘ���FGQ"Uc����l��8���mR��]�-�6WxbQvή�GC�d��{��9��=~#���V�ҧn2뻼ڙ��]��򘛫�όh%f�v]n��iL6,�(��%<{�k�փ�����i���Iɖ�K�m��@�'7:��uP�[*cڦ%�/Uz�C8�/�ZU�J��T��ڻ�Ց0�˜7jf�/Is::�\F=y�5�M��+�ZqVPJ�=q]A�e����L4�g�.��)(�S����u���|w�QOy�U���щ�ټ�FVv��R�Hظ�m��h��F�"7���H� ^�]���C�59[3PF;�ޫ�m>��\�A}4�,6�K�xl<>�ړ�Z_a�u�ݭڹW���R�U;����*���)[_Z=��?���p�3�;d�H�Ik_d�3��N��o�z���e�Q9����#�,��s膇70I���]�DY���6Iݙo�i� ۂ�8���y�%:��g��P�n��#u�Ƌdk�����;��*�M��6�E�n�����Т(Z×�������L@j;�n���tnJF���Y�S?	>kߨ[lp�}��-�,.ߗ���>�YAq�JI�]~�QhNN>l|����]w�pf��HF��6(����Sj�ȴw�G�.���W6P��)��q�3�}q��S������F�J�ә����4l�>sC�UZ�mS:{�:��zu�o�e�h- ap�WMq �Űs����(G@t�¤�cwS9�����uez
�^����ˌ��_8+ q�{T���n��3��1�䁒d�VM�U
��E��D��8�{ҷ�;df[�z��K���MѺ�8M���ۣ�4eGpPy�ŝF��NLb��5���.��L���H�����+�y�����1��#��h����3�� ��S�K):(�H��s�K����Y�Κc����Yϯ�W��q�����o7���?���g����[d�Ç�T�Z�o���*4˩�ڧ���^ރ��[g��N��iu���ًL�Y�����@�=N�c��5�扡��)��W���=�r�!�	����/����}����9�tt1XT-@_[�l����29�~����7ޏ6��o
�t�m��ۃ*+N��f5������߲�G��:|�q�p�܀�R�i#1n�4�:ؚ��ѭ]��t3u�2�O�"�p5�r�u��U�c8���`;���^�m��N����f��+v�>�ѽsOVTCUP�L��7�ͧ6��e>�y薌�z�{�x�-�[�[�\�3��U�����;4jn�p�[>���u�zU��鮕���d��q��8(�����U���E�[^7����h�2ʑ��w��m����'��{���6��w����P�޸k���U�pi(F�育ì8���W���_];獺�l���T��t�؆OdxIKHt���%�D&m�D�1��R|b��Q�t�֙:9O��:
Wѐ��t�mgrC�@�:��%f��W۶qA줺|�U+�B�q�@��Y���#Χl,LTIrrL��S�h���X��o!c��SyE+F����ӂ�J�ҵl���UC��{V-�����O�����6��X̝�]�S��ʖrE�.�("�=���{����+D�WJ���
�Je;�����9��ɯYA�Mk&-�]Kf]���*�5{s��e�겘o2g���@�3��K�s7�E�ӣ_T��d���N�T���l��i��g�.�ʸJ�2>�����cug5\.�
�ى;@I�F���i����������
g�>g�t��O[M�1��n���h��
wJɈv�������<7C&Z晕�y��9%�L��:%'؃�]��K��B�Fb�+S� ���8�NXy�M�j������_s��A̼$˽&ؖVN�� K��{jX�q�X�,�]�1_����M���R�ۏm�7�V6OQ�u��e�j�u���]�dE:KC�ې��X��x�Ha�]ҬN�iQ5���+!@s\܈!�D�f��0��~��
d��'yzp�� dHP���#�r��IXh�rD�92$XV��z���)~Lwe�$�&+C\��f��+�-��:j)wzz����{@Ż����5����E�|��z�'b80L;�	��u<پ9�F���R��*+��dE��^��
.�
+�n���X]���lY��i�؝�V��v�Cy�������+���6����L��uu��\�U�2�J@��n���5��s^���̥y��dv']�0��oKX90Ӹ���jD��4��GWm��}�f��ѳ+�M%X�^,�!�oQ6O&n�J�4�ݟu�J�5��(�u
�Y\��x_H��Z���
��,,��F�Sz��iO]Zl�������r���6�᥎f����aSr;�V5ٻ4�v��ɠq�<÷�������%����-�˽:�6=�۸�j���V҅�ϳ�)d�z>* @�mp���9���^�ٍ.�2m�e��4)�>H�o����HS�vM�ʦ�+�b8l��,�U2�.�v�LudlM�������E��j�j'�WGw-M=�@�؞�8N�X�̮g�FTGq���oÍ
��⢓>���	��0���
���=»QJ�����'E�r�e3;G`w�9>�J4�Q��_d����z|8�OY������`x$�y�f�����W�0�r�Y���ytj��4�F�� �Ď!�D�-TUUL����_`�R��Q������?��_��������=N�U5v��3yh�5��DDPğ�j�W�/0�����z�����~?�������:DM�T�v�m��}A�EAz�%-PQ7�s����ׯ_������~�_��ؤ��%�ajj"�*�u��i��h���W�s���ׯ^�_������~�_�{v1Q�O�bJZ�ƪ���E��D�*Z���ш��T�A���9�TQW�����RQBSHSG���(K�W�*�J]�J�D?-���<Sb""��O������CBh���LMDD�dד�N
��������M4��>gnd<%��"h����J"�X�P��H���i�/ �m�d5U��ۚ���}Z;y��m�w��mEyF��[Kt� �NO�jW{�����j��������̮����#�����Xw�]������Zvxk�@��m�M���^�a*_'��6�i�V��x1�-�$��\�	�wdo+o����q�<����#���A���B��c�`�ly��oќ_��(i��1��_8כ�ʧC->�ۛ�{�| W�����y�2�{�4g�Y�^��5��X&�LH�
�G2/��/�8D:(�w8���Q�n�;�s��)u{�=:z��u�R�lcw�\��n�{PT��7@�;�3v�+��j�������w'�O���6]^�bg����R#�
�G<��1v�5����f�Q�P�����3|��)�U�kj":_}e�S���**e"܋Gj�^�۫���pPAT9b�J�S����^�믉�V"�-�o�D�ae{s$qz������@�ܣW�N�c���ں�9h�v<��S�����Gӑ�ikeh�yG�����1����԰�\�y0]���^Ӗ�@����Eh#4I���9wXΐ�I;�wj#��x�kY��J덙'`�]:ġ�����8 t���eŀi�^���ﾞy��������G���0O��ݑ��S���e�Fl�
�s0���g:���-8Ul��eЮW�t�3�9�/�����TZ��>N�B��w@���Iuy����R�Ռ�X��{sbh���m�00���~��Z���h����dGc0ٷ4�ŏ�'�L+��i�����*�l��r��*{A�l�orm���[����z��Q�=����]���5Ⱥ�wI�QP�[E����ݦ�������l�O ��i�a����gU3~O���׺�kW�Ŧ �ٲ�N�}�����1r�y,@m�0l�r�F�?��z�Z�-c4��sQ�G,͘C����w���(�Q������b��9@�ݚW���(6�=b�J[8Z��^�\q�~��e�:Yi�{-���o��Z0au���bm�:x�m�k����[)מ�EF��a�c��;�^2_D�&x�P/ӳ��*�rQ��R�#��%�E�8w�4K.�S|U,bw��j�@�]K���k�I�aYV���8s�j� �r�c-�C�-<�hw[r�{�����"P��j�p�^��L�P��9i�@�Ԗ�)+3��X�PUu�)�81�l�������҈��M��@��Q)�T!F
9E*^}�$>��w�y篾��;����_>�Y����E�^`�Խ됕�Gu<1@x��j51|����{��F�Ķс�d�%}!v����%!qȥ�+w����{[hv�5��ަ�ͩ�ڹ!�Sz��=�*�<������*�W�d�"��d�d���֓�*���i58�5��ʆ�\�VlsSd䫞T,��m}�~�2��2jusyT�Zmׅ�wHn}4ߪ
��
�`ffF;��V5C3�5۵q
r�{E=^�v���{+d�.wg�
�aB[ g���UgBnh1tsm��7E�Ѐ$�<��+ J�����u��<,��v�U�g:1b�p�!e�?��t�@����z�sY�l���r��<^_��Ahb�Y7�:�Z����`�e�1����=]�޹JR�&�Brw�79�t�٭�i�5��T�(��8'�����^��:�gn�q�L��kA�۱�8ui���� �v�ᯤ�6=�Ű�rb��O5�ڎ�������V��Wv�N�����{���f���f�O��/��0-R �%s��De��+@-�y.�\�:���HM�Fe؉�����y��o7���|��sE�AY������dGZ5��@�®��ӓ�Lj�"b����Y�M�[����.���
��:�}"�XŬ�5K<����T��~��w�]�n�UȂ`��Y���R�pׄO��X���.ּ��$v�E��pq>"AT�6S��U��j.����k��m�16�q_3U��t�D�@*������G�+��+S:��|;���7kL��d���4�^�v	�����u{q�ǂ��vl�;�8���3���N�N�$�I�HJ����]l*��T���T�(p7@�6��5P�cL�8���ܜV��~]�	7�N�ͼzi�������u�h���;��٭�������J����Ss4m��0���m\?DK�3��ɞ�x،\�C��^���r��c��+�콫���əMC������� ��W߷�� `�Qe*ƙ���6��^S�N����C8��8���\f�ژ���1۞���ͧ�n�3�[�q�I�����0^���_1X�5�����5�-X;�������j�kcsmR�{��ʬ�ly�z��^o7������b�3����_4v�����^�)�o�޴����o�"�E�V�]�$�7��C4���P���M��os%^*��O7	�0�[���(���|Ҧ#yNl^�8Ʒ!�쎈pe��	q�q�)(��>�c�,�H�Na����jl�̧�h�Dk�fl(�Nx�v��{��C�;�@�;h�z��d#�����F�M����D��3�ޚ'�ykNߨp׌���ͥ�`�W]CFsN�Z�i�5�)Ae����&E�{��.z���LkY�+�2���'㞷�|º^.�?��sĵό������l2�X�/���e�ǫ��l_G�d6U�l�#�lO+3�^Qۓ��%/�t���������x�{a`�k���=��d���i5�*�=���}���G�~�߃��E#�#�D��kP���g�N�t��3w"�50�f\�n�٨��u���^K(}�PY;n��|&%�IZi�%Ĭ�}b�R�ݞڨ�v����j�?5o>�����4��WfH��̆�݃s����(�1�kt��nv�oP2��&��������V��۪4|�R����Nˍ>N�33�A�`:��U��AɑT��vlwKe�ޞӐ{CWq�W��O���m�2��e���)M=�?Wϧ�J��w��
�\_,�PDf�;�9V���J�q-��*�+w���[����
��,'NV���k�97 �ͨ�ޜ�r�`��3R����&�A,Ǳ�œR�hs�޼=�n[y��fzj|�oD���ϛc�*Q�q�6��>��vg�����ȼnW3�Y��U6��n$V������r�{�xC6�g����zn��[%+�oT�u�q�̵���'�.�q2����iz����+�� �=E��>V�X�3����g&�ՙ���N��G�{-��I������'��S+g��m����ԗ}�}Pj���^��*�ίL^���B��?e{�N��w�s���2�Q�*ߌ%#�ww���wpk��[]�_�t(Y��GQ^�&��F�xl�j|T�����SI�OP*v�V�֑�My��Z�U��[�٣�����iԵ�$��n7��Z�X�+�N�6���ψ�ͅ^�ǩf�A.S.ȁ�(bT~G��y�盞y^p������fff}zb&�,��k�qT�!���=� �a٫=��#��?o�zs�K�L�}R;W2г�i!�k)���^��e�"0����4a��~����}���g�I��϶�OX����֎ �y����>�U�`]�7s�	����E�q���AX��ʗ��s�'�� ~���\�T:雜�Y�M��d^�B��=̮@Jݣ�XCN��@�{ko:1�luV�Y{�v������h����()�!m:�������f5���k�'p���cs/���ґ�l���r���K�$����
nx�C]�H.ї�j��Z�e�z ����Pv�̞.���Y8}AeKaf�{:+���U��s5!��]�ʠ��U��_MO�<e��k� J͝[����w][�o�,�m=�&�J��<�ږ�f��af��!��l�"��ߘ�6���;n������M9����]})1�*��V����a_<ۿ�o]�FW��`^����7�'L�0r��*]c����f��oAC9�K�k2�v��Ϲ�A��GMϬf�YiV^���Z�3�L�B��9��������y��o>e�݃�(nnϗB(�=z�n�`OMz�j��u��в<��
�|���z�Z���:���\��͕���-l���~.�f��ʍ�|hk�7'���#�����Y2+��
�J��w�T�[@3�}Y4&hq���S0o1����v)�V�G'�V-U�����ԋ�k�d�8��ֶ��	S�W�'�>�x�:s�naC0�ƅ�hK�yƶ�鉗���I�zv=Ɨ�j�8��nM��WOy��+{X�L�ъʪl�g���������s�Gf�.Ig�:|�Xey�w��<]��Nl�A��9��������i�7��~̻{k��sW�C�z�,n���|/X���D�x��.e���N�2	j�d�c�v�ƿK['v�wj��m���wK�/�b� �Yk-+H���{�ԙ�LSc���OGҷ"Xm��=���eY�6g� ��#�o�gT�$�}l(�rK+*~�潙����v�kP[]�w��T�+���W;0
IWr�J,l���\�4x�<��XWg����ӗ��9���޻�{|���|�[��fd�g���	̖v�����ײ�!���6�95���������]����<��ܮ�]�Tj��ҝ�n��˘5��1��<u"����Ǹkq����\C���۝pH7v��*!�73O:���-so�?{�>�1�h��B�G]ǹ��ax	J�ٽ�V�5U��x��t���%F�p�:��=�
��F�a�#+O~��ƻ�?{{ͰVa���,�(�Q���!��n��OM�z���p���'ϣvG*��/����GM���Ľەgh˃8X��GY��Npo/7Nϛ}�%�Ȏ\q��W�r1V�byDS<�<gv�u�W5��zp��~�;�0Ŝ��F;pZ3��%���޼��w�LVc���q�Yc���;>Ở�`��F�%�Qƽ���9ֵ\s���!��#|w<�l���d�f�1�2��C����d����|�~p����S����]8Do����u�&' ��Zҭ:�/�3�Uj8K���Y񉾭,��;�o�t�M�BiXy���8to,l5y�Ӯpp��(�\�X��� �R�b�n�o6�ݗ}"��$����k�_�����7����o7���v}�ez%>��۠y����kx�Y�L�����l's�"�&\���e���lq�ҴU�G13���<v�'#����676�ĳd2�{��ɈK�oTE���E޼d[�Kg��w��}�'�Kh�=�#fS/oS�;m�����h�ƹlWw�*�H���|���Ч���Q~�M?�����j��O��w��V�k>Z����\�ZOlV����J�[[`�>��[-&C_�~��?q���&�$]n)���y�Qj�QVǋ��Z�1�˔��H�[�	{�cl}�א�t3��,��:۟qqWя�� ��RQL�0�\�x����Q7w�gj�m׻�3R���a��=X���]��w͗�K�&��b���Tk����U�S�w�*pY\���^�+O��[>�E����>��Sx�gT��t��V��y�����tz���VO\��B8�م,�bH���	��C��Շc��%9��k��2U�"=c#<�O��mjbӸҥٗp����=�8��v��4*i�܉���X��3�A�Բ��ˎ���9@t=!7 �Pغ�_ǒ��9��c�����������'a�t.�n�xlӛ2l�!&���*����}�6K��V`eZ˻	' ��Uj.�G �@��W�nP0c�[���3�8���(V�a�7s��ӌ��e�bJ����XtS74Z�r�%� ��\���Y(4-�ƖK�3:"�i���Gp��04H�Q_=���۩�.���z��<�36�2�t����p�Ĳ,ͮ��d�w5S����+F�>A���J�cT�E���؛X�̈́d�:R�N�J������k�X̉Ǹ��[��ka�#t#D�pu�в�Q�0��q$͔�2�m��ɗ$�Y�#�3�=|<��Oٜ˷x4V`s~]sq� 3v�Yx�T�N�M�{s�K��0�P�'�Q�m�f��*d��C�u-�s�j�n�.j��:�]��2ꆮ�C�:������s}W'Y5�v� ���jD6b�ާ��e� ���E�[@(��-���^�7Yp�6�͙ڸ���b��W�4I�/�v�`gBh���6��~��2棺�TH3.$����rDd����R�<dd!�B��n�(_\��4јU0I"��A<�FP=;�6�Es�\M��<TZ1]�̏���m�#rh��z�	�)z��'�������ω�.���5v��J��PvzN}�u�¢5��q���u��-���.���9D@�^M�aW��lL��o&�7)��Ci���h"�R�6�7�mutû	H���i�I98�>��aó!h�d�Ź(^��Yp�e�٫�->��l
[2� �aЮY��A�&s�.�A��o96��-�`<4��l�,pU�M*-�:D��^�� �#�s�΢�݂ ��U�M'n�Vv�-�dk��Ŵ���B6�n9iu�{YS�^�M��3!ʴ֙�ax���[�j�ɒɗ6�ec��PS�̼p��x�-Ҽ�] �t��Z)�ĮNO�_���{a��ɧ"7cD�]x�3C����8��V_
�H��^��vcoͻ#>��ڻk9�d��4,C^E�Qǎ.�(+��o��r�!k2�au;%�]F��Mb���B��_QZ8^��7L��/;�@;rw	R��/��-�m�之{�*�.�7��r����{���۝E���ֽU�Y#E�gnK�ޮ�,6��.�Sߦ;ւy ��2:�LX/Uԫ�*Б"H��Ye�T���	,�6�?Tem٠]�^�r�mJ�"b�:��x�dPm�إF\���,$�8L(�ǄA��c��U	$n=-�4�w�v��%�H�Ki�X��׫~m�$7T�D�E�s`��h�"��
����?Y�oO^������������:^l14L�UW툪����#N�*�~�DU!]�3�����ׯ�����?�������%������*��cAs&�9�Ǐ�������}����������$W�j�����^�<ب����%�Y#gLm��9��}���_������~?�������b���𒖩"
bjj���JJ��$ղi���5�X<�i)��)ֈ�ѥ��Z[mi�4h���th��"�(�bAH�)*(��i5�������5�"��5�^ZKc����ɬͬ툴j��)���1�X�L�6ƒ��*�冝	�>T�4Q;{�
|���E� 9�.P �A�b]G���^��Sr]�=�d/�͠ �@�Z�tn5���5��ݢ�s{�����t��*�oe͔�\펌��ѭQ�&�*�ny��c���=�1^{���ff`�����Z^&�;l>4C�����y�V�l���37T���녯.��r6�N�M@s�1W;��7q�&�V��c���rt���r�F\�������f��N�rz�Ą<X݌�.�Яr8��u�ln�E�.�%ܲl�@^0N���;Sri�d�xicݣ7O�t׫�L+_|��'��~Įk������-/Y���-�X�)a�1q;�ei�/<�����7)��$6#t���Z����k"|�on�L�*�S�[����C6�>��Y�s����Q�9�r�e7����f��w��~y2�5c����Zf���q+A-ז�O�!�.��*� twCk����Z�#���:�����|�J�9���/��� ��Ӈw�
��ˣ�l��<��=̮R�h�N�p�x�h��Vݎ�Z�?WJ���s���~�f|��`�	�Vy�ө��� j0~g7���V��6H���K� 6I��&������楁kЦ��r�����ڰ}�~��Q���W_8������\u3���]�g�n�H>���*�MEI�A�9��Yx�����;{2i�g�����y�����oQ}��k����LjQ)��/�b9��عQ������&��i��x�&=-w��V9�B*�;:�GZ&^iZ�ݨ��D�7V�����7�NU����7.�6�;7�[p���]�U��g�/=��Y�r���9W&�j5ns'C^v���(�R��9:Ӕ��Z7���7���&�ya����KT��C�P�~���{SIZ��{�^A\�|�����{y�\�r��ۧ��~���������$�%�;���G�򞐌H�ؤ�k�����%����$�k�'���Ք�8{�����H�ǶY���/���� �Q���1��ݰ��l;5N����f�-��	K�iᔡ������9���~��j���h_�φ7��O0a�C��#]�������eʬ/5a����ܺ����V=,;��\W�5���m?��2!��1+�Y����7����՗�NE�AA'�B��4��k�m
>�j�Q�v�^�.�jc5�8���zf����7-�{5��f;�K��[���g�s�����T<<<*�����ǈ;����@�h��OT��9B	>���xY��~�pՍx���n�^�b�lz�a�����z|ڭ�(`5^��b9��OqT�|hi�p��^��f�n��TPJB=�6�f{2�TI��qǓ_P���ʷ�3�ʩ�7�5�~�-;�����ixN��ҿi����̖W?��ۿ���<jC��*����Lzg@��-������grf�c�t���;j�b�~���pف�c����M����0s�y�f�=�3-��Veީ����t��\.��Wˢ�x�0W�M�5&�C����=���"��״�l�&��l��x���_ ����c�ND:��Q���镻c�y ��F�A\)���8�Ӹ��RxuM��*K[��r;d��Kg%��g���4�ĸ~�j����dh�_�5뽆t�x��'���؈���I�/����{�)B^?);�~��g�c}�k��lq�e�cVWm3��;���s��4E�o�ޥ���R�O��Ul�Y3�Zfu�h/7����o0�����U�[yEG7@m�N��uRj��8)�:^��w��ޟ�i5�Sh���T�^����G7��F)���>`�2��T�ùF\^�	�9S2��P(��~$�>���Vo{���<���V�%�;#��cp8m�Xs*�f9��Q�uf�;�]�qYŽ�[DLv�3��P�}�u�Lr����e���ljw����c�R iǟ\�����<ӆ_L���ƋΘ��z�jj������{}���d�v����h�xH��h���S��uZ}oA���u�����1��\���ﳃ��Yqe�,����s�}����#�m],��Y�m�z
��Lz���̘��W[���=�b��6�ϻ��֡l�Խ��'��w�#��������-�{X�8�V{��� ��������Zۈ���A����[�T@/�Ǻ�k��8�&B�����݊����?]kivbۘ�ne�Gɕ�]g�bn�N5`�F���h���F,+�ȃ�i	Akh[IU��6�ɰ�p���%�x{�F<8%M���r�]��G��x4���m�m�(
0��D����պ�d7saC �9"��C��&ŋJ���
ê�������jg��I8`Dpn�����N��_BuV�ΨJ��uu��cz�ֱޢ���QH�ǭ��4�2��Ё��
M�8��w���G}=�����왦&_��E^z�8{�w~��68!1+�{?U.�aě��{i�ĕ��7oOT҃H�xH�W���%�e��snvb�����<>�i���d�MS���;����ts�msɵ`�ҕ7�C����w�)�3l��f�uy�
�[oe�ں��wZ�zK��R}�C�,�]�s���vcnoDBw�������om\�`�LmsЕ�>�ortWr����rz�T�
I�9:eW
=��������;}3�\��7��,��,�x?'uo�m}���A{�|�#̋���ʇÑ���3�V��V��a���9��*���j=+6C����v��a�T�"큵�����.oc���9�V{ݔ��.�}~7����|�
�vӳ�M���.�	����/YHݝk�^���&��.���������_��Ç�m[Xs݀���	�;y�U�,5��}��>�l����IL�͏V8$�E[u�1�_n�eq1�a}�����7���su���,�'����B��u#��0�����:�{%2h==�Vmmס����4���E�v�H�'��G���0_?N��J�f���mA�kv�b��x�y-��m(�=�i-y@+�h�N���j�y���/�7v+�����H�E�4�Ȫ='3��	�����[k6��f��Ƕ��O�,H?zJ��A���	�b�t`W���^���ES�`j����6YVVQ��g�����s���}�E߷��Ϸ��e��w�46ZSw�
"d?���ovY��{`{UW%yT��U��_M\�*+�g4̪�{����7�#�]B��v�1K#�-ӓDm��E��_�V�Hk|*�o���Ŧe���YΗ�-�6X�=a���eˉyY�
��j�{�2D���[�]q�/�����ꗰ/%�1��Y��=�{y�]c����������RC���/P��fNͳsW�T��.���3�t̶�:ҖUX�7Lz%��n��Α-��3�t��� qCt9���f�� ��齻�:s.���\�e�w��v�0�5sª/1�����@7����y�^��0d�\2e����y�tW\l
Jg�}�*m�LK��s�7?���������b���\6O�<�w�':}��=<��Ϊ��x�`R�կSp򮮻5���6/*�#�4�W���y���v#C%k��H�L�����&'����&��,���&w������~8�|u%��u�"��CF\uk��題��3Dr*Fah�q�۾;~���ɅҸ1�����,��V��]�:e�-Qy��b�tR1��[x�>��UĜ�U]I�(�S�y����Y���bo⩞��q7�%�V���r9M�ێv�m��^�c���q`��WFf]���x��B����3�v_ϻ�n����R �o�獼y�w��>NMK��V��Ȇ�.�%�t2E�t[����/Z����	�5ՖW�|9{����&;��g�1gLe����9�*QÂ,�;����8=Y��fp�ρ��V],�^�5of����[�ͼ�%e14�aI|&\5�t�Ev)v�wH�-ni��M�L\��fs�M�ټ�'ƀ����y��o7�n�t��@u8�ّI-��xf�V�57V^���i���>���a�dzr�����7�~��'�N�@�J�	�p�8���j��۽4��J.!��e_��j��pP(�R-������	X�N��W`��3w����=��.�\�j�̝~^�_R 䊑�!�]�N[}����0�f�����mC�u].6I�����6��eսC �#���;��! �MS�+�#!����{�u�Ŀ!7Պ��7�6`�Y���t��N?k�*hŖ&Y�Ȱ�T߼=C�+�dNe$
0��dp�t�w�<�Li�ԇ���Uy˭��L^�"0��y���P�͒(���h����>����µ�Gv��V2n7"_M�S^f�D��u�A�������We���1��A�MZi���38dO�Gdτf��w�>[o���iU������/O��e˾Z4/E�FpnHԋf��q�=Ӌ9	�,�d�������&w'��xH�nӞ qw�W�;J��?���{��Ζ�Ow~���ɭD��Eu=��-�M�Yf�,͟aħ\���e'��v��Y!�fJ:�]�fgV���ys�ܼ���fff}����xZd���j,����bZ5�>�k�z����:Ǣ�+�Yb�=vӒ_%1��'z�_����t�hR�w������b�@���N�2ZɟB[16m�|�%=�ݕ٣�O]�� b/�>�s��<z���5��Q-��)�ۙ��9p�b�h��Dq5}���U(��R�Q��ٝ�E�T�p�415�ܣ�5ڞ�h�^�"&�ܔ5Z�uS{��p��Z�\�䱄���4�u];�����AU�U�?��z�	���Wx�7�wC��^�X� �6ׂ��6�啣U-�wDUV�|˾��/y���D�ÁMĪ�� jq�
�6���/o�rf�����߄h���oT~�։X8�q5�K�z�CY�>1��n;�h��Ǡ��IaC�����Ule�}ZY�6��ѯ�"(���<]���u/޸�<�U���17�C@'�n�i�d�u	�/3g�w��u��};tʔ�z����sC�����D}�}�s�͟����oe��o�Ȯ�;VTw�.]=��|�Ŭj�� [z���+�h���S�C�[��W�]�R@|�7���~�85�n�gf��E�f#�k�E�4���N��r�a[=ϴ]���7��ēÓZ�=�P�T��J#���zC�Y^�eƟ9����r0�gR9��e���δ�_��֙�s�6̋�����ʲ@��FF�'ݦ~�z�
��>�����͗n��#���d@Xd��^��5��D�N�Kv�G����=�e���{=
iý&���j��u]ci��\8�]��\��-��j����;_3١�����O���F���b�oO/��:��i@�g�1ฅ=̮|��Gu�[��`��Ǫ��j���^�E�j�Ȼ�[G3�{��q�|�{�������Z`��`���H�wo@�7����Hz�ӕ/�=DoL���fUS���]��6��Ù8x��vg��17,{��=oR�����!�!S\�*�7&j��=����Tw���³�+]4�[�ʣs{����/'=���8V8h�m�r\8T`oZE��\@����vc�@x�V�[l��o�8��gA��6db����+^��P�(2�X��(�u}�w��^�3�8�d��Ѭ�9=�h��X�t5��7���ʜ:�qX^2o:�^�#c��q���,��f�U�d|��tRTtݚ}9���Ŏ2Tێ��K��ottU3B��q#��j	
z�[���fU���*��9)Lω��!�OGK��/vƠ����e��jSMQ�㇙��c1�5:Ph	����WKhS_M�������YZ�I�{�,�,�1A�+2�\Ostm�)��Tٲ.�"����+��{�rV���zΗj�Z���I;�6�i������z�ffu*Ժ-l.D��6Y��E��|ĲXʊ�)ݷ�mm�Փ�2r�3�d����6t2�MgJ�St�u{y�f\�֬jL�![l��%m�쩵��zq��Y>�>�R߾��W[2�@��f|�Iq�cJ�6�fդ/�Z�
�C+pb�tJ�N��=���~�_�ѓ�@�ȚeM��5��q"���;oyv�M �fB%'�/0� ����9���Iq�[�e��.2@֣�@�>š`@�ܡ�}ћk�u �s���wN<��7�]�N�n3��7f�0vTPI�����~T2�N=��O84N���"�7^�\�p�8̫�0�C�b024�&�i�l�ҏ�@���5v_�I֘����6�CX블x=;d
9a��V�u�X�t�MV�/���Ju��˳m�.��?�x��8�E�5�Ln"2�,T�c ̇��8v2�����8V9�
�}��Z8��;�;�k�� Y��c�"�n�Hv�%McN�ge�x-=r��r���SgK��1�-�3�R�K;�����.J_2��5vN#�a�{Y�N�}7Q�}Ga���X����_����	�ӿ9��E�j|�b`z����iނ���2w����:Q�.�#���U�철�����5�0_�|
U�K�SD�+���7�W!Yi�x�H��^��fL��{�bDMi\ig]�|sS�ĳ�Y	l�Xu�Z�ojgq6�H��"�7x��9�D)��EΩ���ژw��u�̐ܥ]L���Cw1���Gd�[MP�#�y7�E�~�9d3q�o@["�����E��V�}t�MQHƎW��2�d�8ˍ��}�Z���m=����6���d����nΕ���`����5EU�U#��dg=@��X���[/���u��}3]�Te��wN�܉��"F�bX��3�:�W��%m�u�fh �ly�{,N�v>��������wL�j��r�9�	j�y����uYD3�q�e56�$2V�frO�Q�_m��{��@�)\����S�<�����8�-�`k�̒S�}�r:�2����Օ��b�8S��C8F$�3�wp�FF�����ٕ�����4��r����<ҡ��k�/��-�7W��mY׋14����c���8ܷ&�P�ήq:u7M�<�]^@V"G�<�U����Ѡ)J*����rEY�}=}>��_�����������ع�T�W�5�t����&��4�Z��Z�et5k(��������~?������=�~��V�lQ�q-��[o��3���lZu�A��U�Mfs����=~?������?��[A����SPi-�ާ˚����1��Z�M �|�c�|���?���������~>��ǯ���~�i&�m�-i<�SC��lkl�))���kZ1��ƇM4'�9>E+FK�a�&64i��V˨�5�y�ʢ
<�yL�O%�<��ZMccM63�Y��MP[m�d�ԣ�X���j*�k��A��V�-r<�M�<��xf|�����!�Q�����-�5�4Z�ĻZ�����մyx�LPEExA�5�(*�����k@�hhM؈�����xkͰ_ּ��V1�1y���*5�<b���mb�h����lX�e��u�o\�����H�`���XX�$����SN�W����������>���a���J�R�f���<;������~~�����w9�?��Ϝ���)*Ѿ�V<^���e���r�z5�_
�����{H$mGmz�m�y ��ސ�	]��u�7+Q�����n�z|�k&�?
��)h̷ٙ!��u�>��/C�����̖M�]cVm���g����u�5��d��U�#=M�6d붉�P���U�yN�ޮr���δc�[W�̉�g��s���xa�%�b�_��7FW����P���GE.���k�%��!gu�m3!�D��G�3�t��������-�(���1*���7w�o[�t��;�ܰ8��9=���>��{���Ό与��]���fC���x���޿j�;y�5���-���$��r���O3����a�F�ð٧+L�a�`0�o�&���,��n�xwu��[/ѣKRx��~�ʅ#Y��Y>m� �������`y�-�m��g��"_���b틶�X�����Hf`t�svY��}���;�wc�s}w9�=��s��$�_v�%����1�s��Zk������S�}u?�����?]���|�^)镪��w*�����A�޹iԔ����y�o7����&�?}���Mi��lϢo���g�kx�M믟
zӧ�59�:�Fl��mL��g=1�O�nGR���h���y�]��O����(��ϬF���TR�ކ4�ڋu�*��Ԉ馩xj�@�[<��%�'�i#N1��'^��U'6��+w����rҧ��IoWLR���s[������5kݔ��Ԏ�\�G3%*���q�z������k#ާ�r�y�BF�˾����ێ�+���)b���W��ܟ9p��OQƝ5�r7g����9�殆�H�
v~�c�ew����ʇ��x/�O�V*�ڟr��k�h���GjSŏ�����`���4� O:эKǭ'���v�F��T���k��,}Y�/Jp�M�`U���!�� �ך�#+S�/b���P���g2-�����|�R��+�i�5�TĻ��c)Y�Q*7���
�vA�2U�<1�v�)�Td]
��ٲ�0K��إ�hk\�W,��i�О��pt�B7��H�C��j���0龕�8MsT�alE ��6����}�5��w��-���di�N���]\�'a,�qU��0���������_N���i�����9���鑼��4q��wVZF����j��t+��^&�^l�"!t�&��Ew���\��>��4l�i�WW}}��4�o��λ�
}��r0f���[Ɨ��Fݘ�Ux�Ѹ����uo�ƃ�k��ƎR�Ϡ+3`� 3�Z6���J���K>Dv���y��Z��4g���.�l�Ǣ����a�.y��J����ҥ��e�{����}��*᫹�[ԭ@kupE���2n�Gk��{I�8
}��v]���CY�y=R|��Ҍ�aX+vts(g��u���3�ޡ�c�k�x�NR�x�N�|�.��S�;�0���y�D���ؐ|��=U2�r���T�@�T%C�-M�]�^�V��`�\֟_[�
��Pʮ_Uz� �^�buҴ���`��7�1�]��(�����	5.�^Տm��{�f��opb̪\�o�=���;��_\��*�ᮬ��w����u>7�F���w��c��Tu��g�|�	vgS�g����E�X�d����ڋ����3O���y��o0,`�[l�={���oE,J��^4�>�y��/C�9|#��4�j�銊�A}�_(�E�	�ì��[z�z��q��5�C���Qo�������O]u����q}�zzu��4*ZWl��|����吻z�jh�܈���|��E>D�ꡛ(�O�]��N>VU�a�*�寚.���Ov�����*DD{��u�������f�ۆf.��
K��k�2�rM�7"�� >���&��<�!��	����8��[��#��V�w��7CB:��Y�/�6m�(�n�t!��ߧN�'ޘ:���nhd(�82TÇ�!ۢ�S�Ɋ��O�׳���k_E׷�>�{%��>�F�n�yy���v�/1�o�6�Gv�Z�O��s�s#a��hdy�2c�Z�3���xGQ�L�	�;e��_d�jh^��{�A�Vy���9�[�'Ʈ�%���A<8��Ħ_�K�	����kfM�������YJ�,�~Y�Y��u]u�~s�D��X6"8�T֞�Wy�!:�n�[�RU���s��s���m�\\D�uq&I瘇���ob����y��`9�x��s~�L����Y�-��zퟒ��er��M�K8�kǞY��Μ�}8�f�N�fd��}u"�cʎOP�>e���8D?x ��&��>��O�}ޯ4=���C�m3��UO�����1S)KA;��c4Wn^�E�ā��I-�_&�mS�{����p�y�&|�l�"2Y��ؖǩ�#]�'�%����rM�8�
��+�F{�-fz��b��VҰ���V!�T���ЖX(�ars:�����W�^���خ`&x�Gl�d�>[��ܴ�xv�\ZY 6F�^V핒�r�엇�]�}��s��Ms6aC�/!�?Uv4
���k��,C:QmƆ��Y�ݰ��ﻥP�6P�ʛ+��+�\m �]v���p��u�53W��`U�Q��Ę�����w���-�>r��騠]=\GCam���y��0�7��tL�'=g1�YM��*IM�i���/9��ICD��R�ݬ`��nQ�:���61�WB�0ȼ�6�맧�ı�Ij��\�z^ ��k�l�qŌ�wسS�:��wz�p�؎N����h4z�n�w���o0��y��nu^A��s[���wV���}Gv��z4���[<$6�Q�ؒ1�����8�,�FL?vaU��p�=��g7��8Y��z��x/�m5�����RH��� 6d85�>K�j�t������N����x���s͌����i�P\[���#�ȀTP��R9G06�4%}kjkړ5ck�\�]ikV�^�mS�i�Џ��N��ѵM��U�I�j<9���gv��b}[���7{}��(G����Sj��k�iH����=�M:)i؄�lc�
�\}��=G�ی�;Q���`Ug�<�e��Ns�f�^^xS�`\Y�ʽ�G.P���&�skiN�x����U�**�z�b!ej^s5#{`R|u4Q�씫�3 *jh�ʷ~k0�K*���|��tzl����+�����D�Zo��f����K�&ܲ;�n�S�_���b��QX�#����Ȩ^VL{ݧ#�Ф�3��#$[!�y57a�}x	"�6j��T�qz��z��Gc�{t-���T/B�(�LԥDI�9{Ifk'�ٮ v�&L��kz��<��Ĵ��HZPq�-ȔO�
���陙��y��������ק���v�궟W���錗W���BGe�9��e�휿6�ƢF=�t�Y�f�W��	̌�O��:*�RF���[����ͯ�rZ��sl�:㯗a�<��]�'țU	�ci���}�,[���S�.:�F�C�ٳ��p^w?\�iO`�nRW��62_-}�tj6iӗ���vXL��x��?5�oB~����y2��ՖS�X���FB.�Q}Ԡᶒ��z0��}; DoLBi���߷���_���_: }H�S>�\�S-�9J��[�E��(�m�I�\��Nl$C�ӹ�{��o~�̜ݣ����kS<vry�E
����}k�N6�����ESo��c�-�w����C���>�Y��L�u}"N�)4Oa����x:C�欐��3ZD ����~�ʧ��;xQc�������>�r�'+>ܝB),-���m�39�ɻÆv<�HV�p�=�d@�Ԙ@k!�����~=b��St2UF���/�̷Ga�j3�EeGF�oE�]�:T:��=��'-��N<9<��`T�yכ�ȵ��$�$�������� �9�I���#��UM5�p9��&�����íˍ ��/S�[iS0�z�LT��3��]qY��]O�CA�h��x�ی�G���;�CZOQ�E��j���U!��>P�U�{�s���I|��[WoW�q5�@u^���Χ���=1	��_o���0���,��0�4rnG�JN2�/d�a�Z�jqZ3�┈��+]Iވx������5�a��18��}��W:�� q�Y*K}�y+>�߻3#~�P625R��{���;���nQ���x=�:�^��2g�\���.s<��ل:������7����5������	�rmf���>s��=�ͫ!vM��-��-��H��<�������b7נ�uU�փ�����;���nک%�q�[�8��7�ܮܟ,p����T;�jV�#]Xڰ/.���g��Ź���.Xb�gjU��E�ү4�;�We��[|u��c�K��nm����pc®D/����s<Xs��jOj���p,&��n��Ҵ#��{�����tʭ�����8�e;�Z&�^�`c����[��b��缼t���w&��O���M���TKF�T��ʹ�#2d�Hޥ�����=Ӑ7��G{�-���]�٦]�Xw��c�_����E��}�>���xf��{쎎ytY�(�`�9;�4Û�!�׶�0�F��
W�c4����N��S0��ِ1���������QH�x�Y���I�ĉ��"&��Y�md��#���E[)��\݇���42�a�"6��jP�LMS꬀�fL�ۦo���k��{M�	��^�\i�KdO��Q!�zDi��g�3�۪�v�i{ �S����y�F��;�����7!�	`WT���2�r��� c���֎J�ԟ�*��JǑx�$7Aή�lm���Ȇ�����ۇ�<��]�]#\t��Xj��y��F	��kc7\FӰ6Y��F��+�{a���ꎹd�δ��a��m�TW�aŶ�x�zDQ<�%mr�.��MR	$���m��m6��kސ�i�8T�A��ͻ� @�⤚�2f�|db��w�Gt̙/ͅ3|d}��T��7�z�Խ�Si���R�rI� �(�F��W�Px�Q��^b����7���H�"��l%V�[��yӶԣ�N��I{�=�eMi3i�v������t�ށw�\��6T�5?�c±A�g�q��oFX.@ٙ&D�wW��R*������D�'Y>��ެ�k2���
sb�d,Ǭ����H���5���
-NN�8t����{^����q��+%K�dތ���;������e�f^�/r֭�!�7x�Mo������n���V۟B�7l�^�̝�:wZ����\}^>�l�t��P���S.�/�Z���އ~��i)�p�Vr��]��O-��w�+�֗4-��tf�|f��=*�)l{�'ͫ�w�������C{��������������&'Џ(��o�>��j����Dk>t�ǖ�q%�i�^�c`i><_ׯ^��������ݑ�8� ����
�������� *���
*����xxBS�����@2�0L
@�$4�0*���M424�HS ��CC �3�M(@��4� �M�M4�"�M!(����*HS"�2�@��42)"���
02	4� ̠M�@�M0�4��"���($3 �M0#4�2�M1414�$�L*�LC�34��$���HJ����0�4��$�L*LM10 CC�C4Ą"@ʬ���40)���2�4�0�4�*M!�*Cʤ4� 00)4�*@Ȥ�zd��00,# Ȳ�3LC8�p0��0,�*��0�aȰ2(��00,���02�#"��0���2(�°2�{ �D ��y +��@ dPTA ��@ dP�"�@Ȁ��!��@ dD ��@ `PQ �x��@��2�"�@2��U �� !��@ e@T ��@ `D�<�D����H����H��M�p	HS*�2� �0� �2�!L�HD��x���Ȅ�L
@�$*M! �2) �H@&�8�ei�dBE&��h`FD eRB���a�+����c����� P� �*(P��o������������w����g��?���)~�_W������L_���������W���y%�^����h�����U}}dV ?����@�b�_���`������ �����)}?�^���GԖ~^Z����K��.���~t���b���UP�Q)��H�		D��%!BP�%B V$�	Q � R�I�H A�I$Q%X�D�D�ID�P�%$�IIP�H��		D���H	P��IP�I`X��ID�	�I�IP�	P��@%�$�H�	D��Ie�H�H�IaeR�H�J$�� �EQTQ�� ��P+@+H�B�J�@%H�R��ШI"(�(��D��L�A �H��	!��I� ��<?�"��?������4PF�R�@(�@o�=����������À��>�� p��������g���?��8���O������� *��C���ϟ�O�( ��`W�hy�P�ʊ�.����a
�
������Ҙ?�q�{���� �����|=O��x � �r�������
���@{�/}� �_�����?�?�������p� ����������
������'�/������`�������?��>��O�BO��� U���!����� ���x�|_��;��"������뀊�.������i��������1AY&SY�R�a^SY�`P��3'� bB{�{B�(��U��R�*��TA%*���%"��(�UE�J�U�H�UU
)T��YJR���
�$RUT�$P�{J�eH�UUUHR����R��U�l*��H�RJ�PJUR���T@�U(�*�"���(�(�PT%�R�T�(�
�@RUE� *�S�Q)Q%*���!�	P�R R�(���R��%_L��UJW�  -#�$�V�eL�B"KPզ��#)eUj��>�t�4�U�̈�R�ք2��R`cld����e*�Alڥ����5m�J�IUN���)!J��x  ��(P��СBD�ۇE
(t4(P�(P��А�7*���
m����I�A�kV�ŚR�I`�ئ�i��hYU���Y�RT*IUPU*��x   �t���RP�ڀ4m�Q�T��5��P�i�Z�
j͋m�)Vڦ`*��B�"�0�Z�6��  �R�	TR%H�PUT�  åZ҂�M���
}�@� ���ݴ(��I*� Pմ
LҴ6�	f�@j6ƨT�UJBM*R*�|   ��H)�a@��2� 0Ң���v�$ցU��UP��* u�&�a�ր��j�0}5U ����*@$@�  ��HեZZ4ͣ6���fM�TCU���j�R��R������ P fVj� ,�"�JT��*�D�  � ( f�  �   ��
S0  f  ��-�6�  X   X� �T�D�P���I"R\  p  ��Z ��� t -�  i  ���
 6�  (@ -�e`  3 ��(T��H�� �W�   9`l �0 �  Ԧ( 4�  �m&  mj  ��@�j� �(RJR*@B�)PW  ��h 5X@b` M�`  mF )DՀ �� e` h�` ���  �~@e)J� )�IIR�	� "�잤�T� )� ����@��@j�� � z�"ʪ�  =5=��/d/?(��1���9�H�q�;S�pkeX�xWi��և�-X������}_W�o�<����k[oz�U[k��kZ����km�kZ�٭UU��>����a�p��
ԫX
���p�dfHrbN���)qJNh�2df�ff�!SKyQ֛f��(�rS�>�jT���E���ST�è��"4�ޜ-�
;ܱb(��H�&Z"�2��kN�[��U����ñ"QùK�*�S"Gu�'h�����Ͳ%5�-�kM(�[N����ŲD+!T��H �h�e���%A����+.MjC!7p3�-͹.��?M�8��ӆV��lo��)�n�B�V�9j�oib�K�����E��*^�0 �ŗ�0������)�{�c�&[x�a\!��Ӹ���[���T�ƍ�"�
�Q���E��DY�^�2k������"
�m�T�n�CK.ni�����n�mjSN�8F���u"��L,C-�:��!��ʣ���"�a�f^ۅ�8�ҭV
n��h�Ou�	ۘ��A&��]53jc�M"H�TǸ��EŸ[�tJ�Z�d�b� =� ��<���M���׭U��O4%BI�hÈ[��c�qd�f+�Y�	6�;R�b��R���r��K%T-��0�c��/F�v���T�v��j�B�t�R�"�m�h�J�Db�B:U���X��GEcZX�3%��r�k�d�[X1L�ۺQ���o.<;#�X9�,KK5����J��%=W%j�Mƪ6pⰔ�)jSAK%��Q'&���^mIY��D�:�Ԅ���S3>f��yQ�j����̒��ՊfZ��W�������b�X�[����(s$v�ҍ���U��B��e�Uo6�Ē7z�ͽTm݋ۂ4k%���-�D���Y�i�6���W�3�Vn��Q����&��1��u!�;�Æ����)v��d��c�2�2�`t��KBYVPtb�LIŎ!1ܹXq�)��Z�tR� `�ٙx�U�k�,�7���*��3Z��lS�3az�:C�,ۣ���XM�A��nY�)����&��L��w��j)�m�̊��m�әw�F�i�Ѝ��lY�^�J�Kt��L\��]�2��u���v'x��B2�k�!ލQ������O2��(a�x�O���	)/km�5�!���؋p��^�������(Q�ɏmi�3A[����[Obw�s6�;*�^�Wn��v��IV`#zM+�̗#k��P��oq����[���lU$��a�1 5�h��Ke
a5-�E�{��m�N4sL{XQ.Z���t��=�eAyHIMZڃ6��Ctک/�3���9X���o�H,0�ܶ�i�|I���(�
:�r`Y�Ub!�YZ�a;b���-r�b�w�E�7�������{h&�E a�����'�����xࡡP�6���@)vv�"7i'(}��ٱ$MR�M�G�^L���Z)%���� R�ǋ!L�XLU�G��j�@TxZy�^�0I�P۶o �a�R�ɱ���D�&�tA��5՚�
�M
xF��&PӐ�{���;in����]"����T�*�%p�WW��VDX��;H�.����O-�y�B*��l��Y��t��]ʴ^ا@�s6?�Ӈ��JZ��-�ؽX@u�aɚ�´6�ɨٻp��\E��A��P�¢[��*�l�v�5&Vp+�;�H�����^��YW@�0�".����hKa��c���U��@A�upj
iܒfi��>f�U�˫e2�	��'6=KV��W��ڳv�͗.�pਓrV���F҆La�E��$���_mebnƭܛ��J����@ǋ>Ie�5De��δ�1�E�!���=Hԏ\�!5�+�dw][m�LQ�ͤ�ûy5���5P�ƑВZ����	4��G���P:�Qq�J�+�K"6JSd�`0m�2f�oqm��.5D�z���7��,&ݫ��k~GvLZ�	`H�U��3AV���y
u4�P�b��2B����bT�͠�K�lbTZ� 
N)1I��7�/)(]+�C�W�n"��؀[t�*? 'fP%��-��k�d�JB�,a��շ�B!xnH�f�8�$L��lT�GE��@�Zc]+g�m0�Q�����U�l�CK4��嵖�nS-P�����L�����2����m���u�`Ts3�X�2Z�J�L"Rǉ��P�FIn�P����idH4d�r�e=KwbW5˗�-�,M��Pұۏ�A�A#Il��H������w1:;�Y�훈�1��[J�����y��Q64V[#��V-Ki��wf��dMh���n��;�b�5Xu��RӥV��Dj�����m�;���Bj�H�|��MW��)ŏ��Q�%@��4i\$�]V�g5r�Ҵ�̒���1fX�{�4Cn�@]]ՔmG^��E�茦>5�$�h�߉�4�ZX-a@��^f��MN��3f�Q*ȥ���� ��6��s!o� ڑ��y[z�|�hZM��lL��N��ʹ]����Z4*�N�=�*�u���%֌��lR���)�q�,N���NV`�Uth�ku�&E���P�̽����T��M�:.�6ra�,�FfQ'^U�T�I6C���%	7e��	�I�u�5{���j�w�g�Mŕ7�b�H��&T�����Pum�v-�Q&���V��u6�ix��Xf�HM����.�4[����S���!Ub�W�vx�a�nU�H��K+ �e�p�K�c.��ġ$L#�H�P@�^Lр�<�x@�S+qP�lT_nm��%�:��MŻD*+�[�nc�7�+1�j�8 r-��i�mAx1J���U
׫\U3#(�»h��8�5GkR�GU�y��vJ��iFF����:��1�nb�*l`6B����b���A�q*xN��wmP�yy)��#ע�Mn�x�3{�/%�OU�h�6�S��J��a��zͼG$:�j��3Fa��������^k��{5�lذ���7`*m�ͬW��y�5�&7)�W�ޠ�b�Tޜݢ�z�lQ��r�h:r&���{b�#��K,y�2���F݋MM˘�c��=���`�d�Չ:B*ʠ1a�Ê��J��ԛ8�p%��Ւ���ȴl�٪���+iY�d^�T"~�`�z�Z�ڮ@B��%�n�=ö�|Z�VҌl���p�� ,�2�U�e���.���ݥQSu��U���8e�1a<9F��D����P���[�(��Ix�V�0Y晣*ݔ�m�rC�
y�n��x���}k1S�B�i�9nP43��5���	BrT��)����.*�ۃS�5�ym�A�U���r�8Ka�j�f ݦ�xLֵ��k��x��V�N�����.���[�J��ú�mِ2p�yR�p�ЀW�T���1ԓk\hZ�{Hظ�4[����^ѳ{�|�J��i��m�ݨ�+)My�e�&�l�B�F>xuln���[$�L�a�+RZg[l`������m冰j	Gx,���V�*f.Ԗ�н�l�d#.��mTq��Y��[2ߜ5e�x爞��"e^����Y�q�8Ņi�m��
�r��VVڴ�ÓtXk���YL+�g�Y�B�?�����U4H��a[�� �4�_�� ����fW�%�F5.�Nm�V�\t�w^�J˚�R�`�ɔż���Gs��(h�j���LI�e�:Qݖ���:��c�S-f�Ĝ��j��Z/7��$Y��$�M�7m�i�d���Oh�yS^�Z߯/l�hX�)
2��h�w��dˠ�jMC��a�1cM;7n�-�֤��6v��Q���<X���RIU�ْ���C{�)��wy���Į����T*��u��웕�O�j����
����y���VG-��$�Q-Ĭ�>Qy\��Q��{�	
W�0�W#ݷ-0un�QU�v����tkF`y�*��F��~w��J��3x0������Ց��ZE˙qe6X ݣHT�BP���z��i(K� ��zu�2\`������]^��,Y��tH�eKjթW�.Ɯ�,�2h�j8�M�K��W�z�V�I�%K�D��+5�J3Fe�ռiHRT�[х�C"w�y�UL�<N3�m���7U�$�Z�V8��kr��C)�r
 ��+qT�l�kfR{�Y`l

�͹&�Zd6Ղ��*Ų~FmZ��1��u�#ؖ��uԤ�'&�zsvճ��+]d�1e&�dr� ��͗ti\��Cv���)��cN�
��{IQM�,E!���m֭nܸ07{����HF���n&�B�Ƌ�3���96�����ڤr�i��F^��x�7[��[rT��n��ȕ̽65�)�yoQو�uf��`0�[UĈ3%�-Z�i֠VAd,�Z���rѽ �Z�($�![�{S�F+�n��iȢ��Y� ����˶�Y�h�r�ZƷUŵ��$�܃$lZ�����h���E&�l[/j�d"�*�`P��u�d�z��'��r9)��CC1�8�u���jM���-��ᔓ�l���̭�dd�3A*\7,k��X�ܺ��R���*�mJy.��K#J��vrRע�OH"�%0J���W�!t�ݢ�����V�`-���'kA+��;/ѥ���������3Q7-�dK�Cu�.��%)6LF�9/��i#�r�ۥ�PP�.�ŋ��R͓Vt�7�:�����an�����(Sw���Ib9G�%�R೏)`��aF�L���-�T�E�(��c����!���q]`3��(lbXv���I��.l�U阱�݊^)[V,�a���\Uf����Y��S�m,��۠��z�����j�P�����y����ːM�I[������7�-��x���'B���Q���U��nR����k������/u��^c�Ԏ�[jopV�5��
�^� ��3vL�`W��l��HZ�iH��'Z�b��q�2����~��h�S3IW
��7%�WlR	{�{�
0�P*{�K�!7����I�X���N�XƄc(Q�4�6 V�x�=-�Q��ZjA�����7���b�PT{XA��nҘ�q4�ԑ��M'cD�t͋Z�ӕw�]e\UYIݭ��ڥw�0�5�aӘ6���m
5�gE������ڳK�Z�Sd�Yb�Y�R�ǥ��jv��4�W�^���P��ˆ�7��;�ÁM��ʹ�Y9I��#r�J4��oY�Qg%��nһ�r�zoL�ZML�5^˗ZCX2͓��Nf�%��\�V�(�E�M�q������M8��z۳�A
W�oj�f�v�09W>B�aB�Ԇ�4����×���+"��I��HGHH�yL)�e�f�"nU�SB��@̳@�p���q\��F�&��W/��^-	��i2��S7�V^��ͬ���j�řb�4V��o�n*ݧ��єt�F��r�I��C��n��YmKP��/~Ur� :;5e��x$Xȷy3tZ�.�
1�̧y׀�a���A&�
��Y��m26�5�,�ˎֽܛb�,(Dj��iaXJu��Qu
3�2c�Z�!��� ��юf�׉F�10��[`KӢ̋�Ql\���)�6��4h=�	h�5���4�;R4dx0e�ͤ�)�u��ǡ7N���ZQjX�t��I�,X�%Ա*�d���nsHu�1�7]�[�v���
�7h�Y�����(f"�;h�4M�����6,�KZ&`��ޔP�{�Vj/\�괉��j6�9�Q�G�)\f�V��[z͂fL�ͬQ���[�S���S :7�i�GJ�j<H�K+/ 9t~������-[����X�QRչ
��/~�
���b�b�LVK�*ʖ�rq�@$,��*������8I%^�Ūr|7M3���3bU��̀� ]bVf���-Q)Pk�]��C4]Vѻ�%���#�i�)���3Ppdnl��ۚ���JAxӕ��uaE�ᗺ�&a�z�i��K�Z��]�/�a\j廵�Rg�D��2�x$�B�]��45�h�F�8����#��+i�
�$T�DⳂel�v%Y>�í���$Q�hӕ��K10���쿬�ǅ���f�ۉ���G�@���`@�Z�@֚�Д0<5t�EW5�s��J��]eZ�`޺v7�ɕ�����5CJ�Ј�ɕ�Fc$Q2�Ғ���2)Pj����
)m��W��ɘ�U�M�����Y�Kl�L�#�����V��ٸӤ^deL\��p�&����v	���u).Y9��(bPn�f(w,��1���Ʊ�Z�5K,���7������,��,;&��� (ZN�D©�jI��pi��4,�4V(j^-4�^���I�Ǖ.D� )!O���V���F�k�3Y{�	�� ���[wq#+M�!e��a`:�&���Yn�X��wXF^�Š0�Rtc���p�Swפcڰ2��X��)IKb
�$�I��onJ�^i��O/v���h;m�r�2ވᣛR��*}�Zr�+#o{C�6aձ4Lo-
7a�ۦ>*���a��۱]�KP��t��mU	f���R�s����PւxΉGn�!(m�QIʖ��
�e'6�X�-l�/&�
����7Y!Y��e\�)Pʔp������3�Z01y��x��v��v/pd
��F+���X�`��]��k^,����i
W�)t�x�ߞ�����V�o,�m��2=�Jm���/pc��˥?;��i])i�f�[s��*4E�� VfS�4l�1�w��hZ����C�Q}\8lVe��l��3/#*Ƹ50u+Թ
u��6��l��۬���^V֧�/�U����>kxc��;��LN�b�]7����wY�5ح+Õ�M��N�_#	FٸzVrXL54*�K2��"�0t���s�]��7���Qy�ޤ�Wn�)JU�g��uYr`u��J{f]�W)р�؎�(����2����X�����,�enNҭ	�;f]�wټ�X%���l#L�J��ޕ9ͣ�T��zW&��ݾ�M¬�Ւޝ�ٶnd��r�hǠ���Nʆ�cD�6�]d�7�7,����(�f�x6Fa�us�zFYu������jd�%��}ܶ��%���N��T4#7,y]ֹZF�K��n�].��ঃSvnmu�[ܜt�������cWiF��0�,���
u�Od����Y`���]�o[���JΧ��[��DO*`��gI���u�q�b�b4�i�tz���ī+�V����j�C�}ζ�TW���nM����8j�X�����S*���v�l�n�#�{��u:�D*���y�]�)��O(�abw�X5tl���(K����g���(����OM!���"�v�;��`��v��z����R᫈U+v��wT^(��;�b��]�p?{���ǺGJ��V����#�9v2 �E5����
��w��t�/9�Q�q�T<zT���q��4�s�R����6/q�����GpvұG6��Lin�堼��N����`���S;V�cz������E�B7��Vn[�&��)���fdf��

��'B�Y�0��+L�N�U����:�t��G����cy鎟V�r�Mqđ  ���ޟ. ���r ��"r�DXj�U���V��H�5�C�H�mMCks��=;�Y�����唷�S�f�־n�/��U2�̾���:���P�|�L!��QK�t��4�X��ֿ�l�|�JLճ9}dg	Z�_B΀8`��kO^�'S�KM�(��n^G�^.���D�Ǚ�@��:��8�Qu7H6���P�#��XɐM���te@2���:�[��PO'f��+�K]�n�B�H�j<�t]�@ZlbGK�*���W�v>P��io.VT��/��K9��Xq�s��O�+؇Xf��sHl������R%�+WXϐnA�1���;���Y8`l�Wj���������;zr7��o5}��-G�v
�&�w.��Dj5�F�Q�[�{��!ʴ�Gd����J�; |�L��	qV��J�$�b|wq"�fuZ�xA�&J�J��ܕ�-(R*�)2�}춊n�X[k)�u򸍪Z5[�pZS�$�]��ݘ�����yk���`��!$�h)ς�.�3�ѩ�٦��	M 9���d��)q�,�˴u���n��2��e�7�*y��UppF��w$Iot��G��q���^�p�.-k�n�6{��p�v�6��<4��u�/����d^�65�È&��ws�	�@N�SN<��u9[Lq,����t�,I)�ns�VT���U^�GY1���or��b�Q�i���0����wN�o/�s���dM�26��k���fX��"�h�����R����i0bY����������s��c=��Y��2��wq�ͽ����e��/�;�h����Z��Mor�u��s�{]:�q��^��Dg}�_:��ޓ��qGb(@3P�����Ƶ��7�X�u�gQ�+�Sƛ��XX�0�ٕ2� lWsU\��ܨ�N�^Bg�0�j w*RӘ;!��W>Œ��dt�fmB-��f|fBY�"�p�K.�D�5�z����K�����P�3���#����;���Q�������<}=�{<�]PQDM�M.�V��hf����)f��@fE,�C�����*B�1�Y@��Ek��PsX�M��ˮ.�	4�Co���v��:-a�� N�sMtJ����o��㏺N_I�vƾ{iw�o�_.9����"�W�:��d7`(��Q`��m]�Ζ���+Y����qB��fH|�����E7q��vq���v�RB)f�qcg7yn�/��"��쫩O6�j���(�Xݾ!r'�M39uK(��P�*�H���c똚T����a1yp�gf\�}s�����;�)wsm�����tr���s{+���5 ۭ��@AB�|�N-Jw�uk�go����;�v�άc�x��������sop]GrdB��&�ݎ��̢�à�~-̮Z\�:��0�tlIʯ{j]�P�q�U���GGt�&e�e���#�]�N��7]��P�-����݇;%�_����9wn�uY�H�b�IF�۽�O>�Ԕ�'�Y3r�t�-CuA��V��u>6L]���R��p;"Ž��=a���>�{%�hK���:1�l�V���j�w���N 2��������r�͵���V�R�r8�$�:hg0��WL�V�A���fܡ[���$�$�o�����>����Y�S{msV*��\���H��Vk5ʋ=����S5�t�Ų��d�*��BSvo�U���Fr��:�岧'��oIRw�MՌ?[�E,/(4Hؗ,܃�(<��S�$��HT����x���E{ua\Z�s:�T��Z�%�V�-c6�m`��t�דN��o%ϯ!ڳP���ojW]�*c�j��j� �#LNv�j�t���}�u�����jŔ�4���kF��IbL���s&�r���):����[�a�
AutR��B26���߶�]��q�-(�r��Q�|���D�,M��O�2f�g.�c-l��RؙW%g�h73�b�ʵ�U[���9���wuf�렮�J���80-��Z8t��SQQ�T��7_u�=����3�cF�U��l�7o\�(����v}ە��7}#T+\�e�5��Ж6��j�~Q̬(7��� ���G��(F��V���)���|L�lz�*��K�J�0m�w�kŕ6�7i�{u�t<�Z������%�����`Ǭ�=�wu5�N�R�7`헽V���ʖ*t��a�~R	��VYT��Qr;�Z��n�L�*{�P��-:ޣ�o�Q�d4Ԡ�e`�"��h�2rm��Glj���5ۈ$䇐������e���gLSo�̥�8&�Pҵ�ldʊ�
�Q�<5+��zV:�o�-֘z��Sk�iZ�!�vLq�n�i^ŪA����Y*Uք5�������U|FD�}�U�Z���Q-���\�����N%�fR�r�9��88��/�R���of���Z
���YM�y�?`ֽ�o�^Ze��J��/A6�X �m��������h���)�ec
3�7�jw�sm���cpӊݶ[M���{�["Һ�婫���q7��ڢ;DT�=)nޥ8O$ؔ�e@�gO-Աn��ڛ�aU�!��
Qt�w��\[�]��ѣ@j7n8��{)e��i�+������ՠS�M���s����ב;�9����&J���e1Xp�}�:���r�t�|{9hƘ썫��,s΂�5݂�r��Vr$x�(zU�b���c���W����9P����7���GR�s�[<��4b���(���q9MCT��Rn�VmQ���uƵ�owk�#1�)-��
�j�*kR��
�v�έQ��&�\fV��r��_+�NY���\;u,T��.�6��2�P&Zo`���n��m(h.9�{�U�b�!gk;T|i���R7u��G0yU3+��2_CY������&	#U��8�B���pk�ȩM�b|��������f����
 �by3�0�j�$b�$�y<}���k��6$�A�#W)BR{0��곲R3�:�Ub��[�1�a�����c�67�(a=zz�k��(�De�x�����4�[��v����S.�X�-,�՚ɴ�<�4�c�2J��pZ�Gl�a�T�uֳH���)_=���pB�ɹ�kl�/1{+�Ö��CQ2\�~|�_0��,}+7�w�F�ol�݈d�
�+r$f
�Z���b��@ʳ�v|(�٢{�:,w)*��̣F5u��R�Ѭ�K�Y���ʮ�ڨ���f���y�i`!iᎲ�
N���[X�Y²���S!ٙnӢ�3{64jk#�ќ^q7#6�'�Ռؾ���ȷ���:i�o���Y|Z��@I�֌��^����I_#���r�j�a�A�[�2��gX�ӝ0��y��Tq�~�}k�ΐ�&)]]���µ*���cMT���h�,���sbޙ�p����:{����X�w[�[T��Ļx���w��F�<ǎ�_n�}�#����Ռ�CVFs���u������#)�b�;�/�>�n�͇boY0p��;�6U�u/{jj<*d�ń�����gw:�R�*�J�WDN^b�t�0��xUL"	O�{����5WB�:	I��T��|��tӴ#�6�t���ycVp��V�՚�q�q�ʉ/�G`w�;�,x�wQ9ܛ�uM�� #��G-Q}�u܎)-�����X��E��L�vo�c�%u弣W[�*���([�x�y��ٌҏC�h2���Ԡ�CsE��8>|Fs�	f����q�28J�3{��v۬kV-���!t:_U�V�U`�U�B�\�+L�z�cÉ���w+�+Ef���"B��GmL��x^�;T86,ĳ���/Y@�.�k����Y0<�$"<��t�р�WO.6.��A�T�ܧ�b�YwwMJou]��>tkB���������	�P=I���ű����9-�" �h"r������b�\u{�>2Y�@[�[/a����Y]z�*M�� ������m�Y�S��BI0v=l���"���k��i��%��`��Ŭɫ�u���h���6.c&b�E�P['l+2��X+��V����f��	ەa0ed�u4%ɼ����Q���}dYadT�ث�TaRw�l�2^��ᯰ��8B*��2�{��d�֪A��f���j��יs���q�C��vw�$󉊴B5�n��64�Dz7�7�}́hFv��K����sڱ��;.V۠Ŷ�kQ�14T����sQ�7+̻�q�hV��
�;�&ʕȱ�K�\z�P��9�5�r<a�Z�:�Y�ae����tp�[ae��E���s
�ZWi��ʗ���p���@#ͤ�]�x����A�ڣ����p�e�`:�g,���]5�[!��:�۔�<��ͬ<G"T�;u2�A��u�v�[\S�^�	<%�ms��f�1] ��51���`�oYZ��s��oLtC�������8��oI��D���@�m���ʳ�:�,��b��Y��7'8�zvi�+�o�7%b_b�\T�l�B�k�F�L�9c���n�1�W�� ��G��.���HIh��0�g%p�Pt�\�I�s	��+�d�����u⺨�_:� ���cG�(�ʑg)}�(I��+�+r�m�S��N>[	=u��v����t`��7bӘZ�(���١�`�{�����������c�.�T�]��|ǘ�غJ|�kUn[�tpXlM���].*���>�9l�E�8Q���7:�l�ʮ1�CYNLޭMGt��+k&��b������t�\Z�.է���q���\haޏe��8�z+��1y�a�U�k����Wl����-����vlfĕwd�tuRL_�K���
h��[�sΐ�ٺ�p�[a�c���S(��0iէ���dZ���K�67�s�+�]�tq�*�%�L���رW���x�����F�Z��v݀�Ю�ћgW7�n��-�sq�wn�t�7S�����2��niY�&� ܩ"�.���M������!x𛽜���C#�$^r��KU�ݦn>4�8=�"ʕ��x�M�;C,�c��
� ⻒��u��kY{�"��U�t�(Z��)Ewpզ%C �W6b|]K����*�^�ow9J�*�vS�,�N�GuG�b�dr�wx�V�k���>9gq�]�B��SR�u,�0�b���A��ʷP��ڴRM�V���ٺB�l�����6�-/�F&��Z^�FK���wݺ���C���i&�6�����k�GZ;(ͧ+��]�}�6q.�3)�`���%��e��� �G<�[0���[�d�!Cgd�n�pt�{{=���*��L���k��̟,q��K����Z����Ƈ�mg"s��O��q�g_D�71`�h�f"�h��c1�Y�y�2����fà�ه/���f���d�/(��'nB��:�i0q郶tޡ��+��X�q:�6�]b;��0䣋�#483.�
#P��9c
9t`w�'+&���6:�8�LNs�`�H9cs��a;Y��G^�ͫ���b`��;�֝�}�8�'+��oj*����S�/�+�F���靈�Ȅ�6'*U�}e9��~�c�S ���u�.أx�s	%���*�guv�19�*��x�d
t���j� �Q僚�[�C���S��)ڹ[���q&3cnV����ndg�rfmF,Vco�ዜ:�ҁ�}zV�r*��^��W��6Rf���u���᭩���w_M�
,��h�/�2��u�k���eޮ�)q�u+s�O��c��ќ]���Y��I�*������זv@��M�#oE"�g#�=e���u0V�����U�K���zְm-�%�<�`��-�s�N����]�(�L�ꃈ��^�+��S� ��۷�o����j��%����	U�\
����o=�t�������WqhVv�ނ���*�+�s�5��.�=9ꊟR���uӉ]��X���7���8h�e�� s�V��3�{����s�>�s3������������Ͼ������ﺞ�/��M*{��_�k8v]��f�FT��e�dH���q\ܵ��<9vf��ƪچ tJ�9w @�!����ݬ��;%����t��q��$.�d�$��������uNJ��1 �W�8���;��t��e��M3[D^��5tm�Gi��Y�u�k�� s�q/�>�H���� �0��A�`4m\yy%�=r��W�L�DC�Qe⇷�v�-�p�;�;�]t������V�쐁�6�Z���83�ˬ��%��_l/ �����U�Dj���Ơ�/;gt�K���a���¥�� �֚���\=�$�s�_^���s�p����e�h��-��k�5-\MLɥr�]v��M9�8=�w��힒�j֧���r�\��1���:p�7ٜ������!�V�Z�<D��I��mд�4��dR���U�]o����[P	�����8��~�{ײYәh������LX���*ѷhuh2��	C@cWR�)��򡵷��մzJo	˕A�M[���YE;�
��Q82V�M���k��5*]�|�=�1�8��^�.��Q���c�}+�k�rܶܰ�M��2��8�͆��V�q��T�{��P�.���E݆0��&\�n6.Җ���p镁ul�o0��h��0}կ�/��ID�f�: b4V�]5�M>�=�6৅��3�U�:�Nq�-྽�gN׬Dn(�ZFړnu�Kk�꣢�я�V�XܡEj[Hm
�9]�12�`���6�T�^J�;���T)�q�Oh��X�R�f��z)����B8�-�g��q�t��ըnwe��T���\6�-W;s���k���.�J��v�����:T�T޻��[�֊`��c���w�I`��ѬϹ��H����M�ʺ��/�.�%b�)	�#�����m�J9�����yr��Ym�)Y�V&�R�W�`Y��1X1m&�fnj�Y;wj�~?R�ĵ�Y�����$�x�A;(���zb��f�;��\։sj���/kDީ����|TY{;��XZ�7�1�O/hw��s]�͏C���n�W	L�8l�rx|���׺;\�e9Rv�0u�R��"M�[X�x���.���Vd�]hӦQ�2X�Y3xoگ<��&E'-����J�TO'U�.^Z5:����w�w� ao�3�Q����=6�6�),�-�niS�S�z�� �{:}xg�r��H+̢y����wvJ���2����jSu��ъ�V��l㡇/z��U�`]Z�u�pi���LP�:yK]�;*,4����xݼ�ig�3�uo\�[X�HX��(�%S�u���wTs,xs��+k&Ӿ"����3��f�t`��Yf��a2��U�lm�J`��Y����ͤRBK=S��i3��w*��wG�V�YV;*� _wZ�q�Xԑ�u��ͨ9h���cvU�Em�+��S�O�\�ʽ�xk�6�Bu晳sr.�׬j�j�e���]��q�e}\��A�e�֎��Q�H�G�v7� �W�iNH�����	n2������oSM�h۔���3g�!P|�8
�F��9b����G�����C;�p�ܘĩ$@:��(��J-�̺u���Ymĝ^]j3{�\��=���F��`�j�m��o2[˩�߹a�/�RkjA�6�b��;a���O��v(����16�0L��^�`ލ��3�F9U�V[P��>ڜ�2�̾S����;5����聖�w,
��{h�W��B��/��uM!9�J�zA�ʴ��̭��q��$EًGB��E�ݴ_<�|�:����f4���@�]��j����Aie���x9�Ѱ^��,�_;���H4PDh=Wdԫ�[j�;N�w4��F�2�l��t��B.�
�<�|���&VZ�`�P-b'X8�v�[�Pj�Y+oj�^Q���fu\q�9vzk֮O��̈q�R�齻|��yϹ뮄�w!YV�֙���;�tj��V���p�@e��]�c�����"o���y�%.��q)H֧W�d��J�T݆�L����g�DS�/1�t둹Ǹ!�X{6��j�]��&t�T\'�X�NE6����U���˴U�p�O9h�uWj[@� b�5՛u}��9�s��!V��te�\;yɐ�d�j�hcг����In*�J��O>톈��3ef�����RƇz0���rƥ7pݭ��f��M0�����m�a�ں&T2)�r��sﺴ:GQ�T+��l}d��MX�\�r���+p�P[؅euZ�[�,,
;�� �	];
�o�8p��c��V�ч�Z�-�pMEo�#����p�������T�;�[���6�����J����H�3(��2������go��{,
B�ͺ�S2�]R9�d 9�9h	嶵�m�bwtv�cz�f�=[;p�#O`K���h3x-�Pdܒd�:�[����M�g�ڴ��̱��e�:G�J���A3}�X`S�6;sK��1�{-W߹J*�f��)J�<���x���:/��9��q&A?'j;e�X���>ˬwʭo�s:0���X�3�
N�k����A��]K¨��hm^t:8�ǉ�$,}Ht�����`X��wJu�����:ӹ�e��[�6M��s:Wb���Ma���S����
 �2�&�
�62���l��)f�(��.Ǻ55tOrЁFSᵬTZ�S��W�6��ȇJ��k���H�լ)5j�v�>޶\4�j����ү{g;�x�nlt37�
�̛;S-��vԮ�[8��xo��i�Z��n��}���tG		���n;�gq��;�,e=�louX׀�37��V�ER�Ô�̈J<��巏��.���6)�;���#�J��.����#�"���ie��}�%]}y��:���A��+�`�����v_u��F�5Yζ�4 4����t��h���e�f�UA��ɘ&�o�T���WԢ�[:�,�qv�]��x�#��c��ά���OV���s�Mg.�ϝ�TL�z!)�iu������W��ٽ�
}��^�+��u��Ϩ4k��ge�n���m.��f5v�fېz�5 U�ǵ0��Z�=m���*u����B���q��SR��]N����T��A����ՠzj�sm䙽r�F��B,�뤪�b+Ir�q[!�1��Y�Њ����iT����G�f�Mc�:�e�R��ŀ�
ef�V�͸��K+�<��;�]�����Ě�<"�K;dMv��[,�g�{�a�����}|b����z� ;���3O�kdU���cFJ���-�X�Hv`�q�n��?x)�OZڇk�˚��^�`@[�(�fX�+�Wh�`��Y�����S�#@G��|2�V��ܛ:����	�ɳ��5�sV��w��^�Q���>��[���˕���q�OEZ�Z�4��	�U�;B�ڷj
��E7�Zі�雼�rGF��:��v��șY#�y��;5$c1V��'[��u�N�ڹ��,.��v�>p��yn�4)w��r�/T�'>Z4�8�vI��X"�8kP�kB��{	u��L\�f�7ϫ�S�*�w2�\9s {�q�9�{(m�2Ӭ�xJdc)��F�c��&6��z�0��ܖ݌=���١���:�GPqӊ붑�썼=c�-��k .�]�6��@i86�AgP��� `t֊�S�k�0�Q�}}�t;�؟*}��ݰu,�4�rl�� خ��)�B^K]�Dge�׺�3�'mn՛;#J��=$�±T�j��V94��x(u��^�U戅Q%��2ﬞ����ó"3(`�5���n�8J��f�qLR��FB�YT��`\m>�3P�իF��
W�v�U�oR|�q��1v�N�9��Yù�>-��`u��9X"J��WJQ�5�.};Ռ풎b<���w��EP=�3'Nʜk���P%O�_�e.�_\�,I{���U�W�#���p���5g�9�M�}��ul������{k�fEx8��[],�˺C���9sy3��c�+.l��� �i��n5���
��x���gb��._]�#���T�|�O|**R�j���s9]i����0�ţ�V�>
��]jt�M�1��B-�g�f#�Fe�JSZ�΂�Ə�г���W�"֢M��[*]o��R\s�|��|/>1$n��.02>e-�9Mj-:3im�],Z���A�wd��Bx��ovY�Af�}�e��v�nd޽�4�C���'�I�4
@>Z��iLOv��{��uiX�����+��Y�tJ!J�
��q�\Bݥw�Tmv�(������ؾ΂i�b���yL6;��T��=0�w𬖥��K�.�Lڵ�כn�ȩ��Ko�����ō�U�;z�}��w7�n�9�����j���uj�0��n�|�PV��`��'n�/������q�!n�c��3B6b�S��X7�+j��_M�9*h]9��S��w<�47XY�vQ'��q�{su�:V�D��Y����Ӿ�=����9���z�hw���)<1�|TUy��5"�f�H�nH�!�O��W��\N�4�%���6�a7��H�����7�sgRh�GWV]�"Vn[Q/�����R�QM|m��wfT�BR8�8���1���=������ܝA%!y-�)j����� ���4.�]��V���*J:��(^��{��;�p�<��4�NA.7ݻ1M�	������.n�*ᬾE�h�F�Ѯ���w�-pu�J��8NgU�%�j �0-]�N���fj��;��n;���R:���`Ǫ�;��+v��� �TVQ�u�y��V�������ެ4�<�4��+��%<��ʘ[�j�e�|��qeԿ���q������gV���c���5s�B��ڎ�CH�&�ݒ�U�iu�M=�*�GA�X�Ow�K4����L��Eɻ%�S5-Z*�Q�7l�{Ow���R�ׁi�cj#5jyv�?L]kƀf��8�YЏ:�m�m7y����rb�=���"ϸ��a��{�h4�+�$�� �ƻ����儲���>���T��w��t�1�R3�]�5���8�9�X��P�v��
W-�ԌJH�δgkF�1%ܯ�m���r�Bj�>B32�fV�ڶtC|�%�YW�B��ִ�;�۸��g*>��],�Nm��Р�.�f8�(mV�8�]c�F8 6�k�|v���a�����@��䓭�·S�#^��{^��ٛ�8͘����(h�r5�]2@�G	�(�H�}/�6��`������vѥ����_8��C�rc}��WQI|�"�o:���ڊe�`n�d�2 ������}q�R�_@�*�i�E�ܙ�r�����ř,V�9���[�WjoOH��m�������!%�Ybs��si�U����V���%��3te�;]�ѧ!�k��b�q���"[}+U_�u`4�
��[9� �jV}��"$��j����/�n��@�ȅ0��+�;��Ki�u��J���u�{Q�+�w�Arۜ9�fp[��`����c>o�|A��*�.�](�<پRB�5:u�ܱVkz�Xü�R�[%�][��2���.16z�N�n�j��n��ԻX�ƶ�5��j���|�Y|��d(�fP��Ԭ�F]\�.pZ����}���@S�.���I'���;*]�/����G>�Ũ�w%�t��8�hz7'�ie�T��CQܶ��T��o�N����-�w*Av��B�WY��A\�mwDU�cg3�|�GB˲�^��B���˻���%o�Tn�⏒!�2��=8����Y4��+��n�I���7�M���[}Rk��w�CK+��=�� ܅�6#:���O�d��ne�V�l�C���.(�t�(N�nZP���)�7'�co�a*md컜s霴}�@9���"8l6�e���})���,f�(0��m��.v��N�*��6[�xG3���
��g_{»��5�4X]�E�k��F^3�]B��,��Edel�6�f*�5�+w���������yi�9J`4�SOM�����d��#��AQ� ��ץ."�]�XށE؉̖��n�:J���N�.�@�iT���aU���Zս�����d�n7Q���:|��1�»+6�>��Kk2�Kƨws�_NZw@�U���z�D�u���[�w;T�'0A�v���]rh\>��޸ӹm�u#}.該�ʹkdŻY��j��h�󫡦�C�K	���O2���V��8��4�q�<���]l\�C��Q&&�޵�sS�}�#��|�.�rI`9}�MR��R��ֺ��oeؤ����|@�ۤy3 �x�O�z�FNd5�.�U�(�7���F�E@8��Z�E
�����Y"�794dؖ���a�3��vs�!ލ�w�(��;���!S����/�0��w@�K�#/k���ㆴ^�Jw0eq�I�B��ݑSF��չ@�:w9��J=X�+Zvp6��.��Yt ��#��^t����Lk�t�}ՆoT��q�e��:�xACk¥;���3Yz�H�r��5[ے����(n�t�\���ĉՋ��L�%Rs�{y�括ގv�
��o/o���8=t�o�w�L�P�OG>a�=�K��<8������ ��Cz���m�r�<��:��Dkjɡ3��2=�T���wL{��k/MmG�X{���h��&�>�F��,�۱${��Az�N4������ӗ��l8���/cJx��ׅC��CO�=��� ��#z�b�J��u*)0 ݑބh�|���%7N[+"w�*v�f�Ve�a
�'���FL�bj��r��1�����"�[��n�pn���k��q�.��	����:�!���l9����ﾯ��������|�g�"�{+lϣRPm�� m��0]�9����s��fWV�-�r�k�� 4�7�l�ӕ�S����	nmĹ�h�@Sx.A����9�Jss��[5d��E��޳��5|x�"��� P.��T2r-�uh|�)�^���,J�.I:�(�o;�4�rѮʕ�`9���N��ٷ:����-Ͳ4�}���ah�|��u�h���A�����52���32���k�t��Ta/�VS��X����ͺd<�h��Ѩ��P�k�Í��y��ݛv�!օ�]ݮD�>�teݺ�Y��G���d"�+����dYN*:3y�=K&,t�,�X-s�D�����. �ӝ�6���ĸ�����7����Z�e��Q݆6��=%�R����v_t�v�Jwt Mdܘ��4��.�IZ�Uj}�[R��ف��D,����67�u���YG���C;~�����;6����t�X��_n�kS�oq�����㱜rj�Ϩ��l��fD�v�]X��j���&Fh��`[�s��^8��Y�]n�4��c������PA�-f����\�݊ĆM]�����x!��⢘X�Mݣv^iT�W�`ɤ`���L| ���9b�P�Jr �n�& ��СW�ej*�_#gּ�}���<�GY����]��a�&�F����5G�	�tQ˳rܣ��Y�ҹ���F��ӻ.��s��AQ�wpi4Y6���nw;.�ø�.c��W-�.l���nn��M�@�\w\�ͺ���3���.r��s���'u�p��Q�&(��\��\�gw;�%�͹��p��J�S��˗wl�,k��r�k�\һ�G8�]�'��5˗75s\ۜ�wr�cG$��s�7.��ŝ��cq�A\�����r��+��sH�NN�wv�u�M;����.��Ar�wq\�r;�ι�.�w79k����ݸs]*��ݺwtj�듎�����Ó��Rww8%s�wv��-�+����.�w]̕�9�u���w�v�ܹsS9tE��L�o�_��f�2j���hE,�S�S`�l� Ac-�������������5�>Y(���N��H�m9�'�˕�mm�O�����C�|����Y��k���*�K/��[kC��GK�;�f��3%g��>ԛ _��`>�hI}�ty}�yWMx���}�ɨ�!B�m�Z���u��hl�S�L�wk�������|יǱ?
�Hp�U-�΢����
^�Ik�%?{:�x}~���S�N������ea����9,v���ؖU��ݬN7OhB�[���o@_c��	Y�:�]���y1�}��6jV���0!Z.�R?z�Yr�4OY\� (A�8���X��(	�@��{�����_`����Q;r�Byp8�z$h��r꩸l�X����3����
Y|�t5gk!��
�:wMK��͹��ZAZv�n�?z�×����U��ݼ�;1���ʍN�w�ϛ���Sx�)7�<�{��?}8��5��\�N`�w-:����T�J�����{ylM��1u¾�U�����TaE8Y��2��ɍ�q��n�3��:"��YHA�0Y��^��2��od{�jyB�̲��9XW�`4�Ղa�Y�i�:�Q���]�P����N�0���Q��/m�8{A�t�V����V��㝑�Z�t]M6/0�)�Y�,v\�*CF5ܷl��M�F��s���غ����D퀷�*�ɧ��LX9���L!�y�ƶS8,8g��r�ک�~�yP�vC�tk�*��3gFIe�;�gN�S@8`?/w'x�E3���]b���|X'���1�8�y�����/��V>|��t_L��$XȖ�
�1��ʅ�1��V�#��PB�����nV���g���Iݼ�Kgq =^�2�dLq�B�;�ek�6��=�3>����ݨJf3�Yj��������t]]��]��*�tE@RT�ԆP胢a������s|wH
˥(u���w�Fe-�����3�l�*v@���u<��i�K�<*}q�����n�=�#�>�ů�,;B��w����Y���b�(zP�`?t~D�V��hB�ΪZ���byMt�Ռ�!}8���#����%
�2\�'!����^@��%�&��f��W�b(�ke	�k�wR6����Z�k���.���p���ħ9W���6+��~�:����)�)G`q��.Y�2x���<8�~߯&0W�S;7H?@�X��U
-<��������kѬV��	ER��F�ͳ��lہ�XEZ覃�Xa�bѬB�'r�o�dT����*�w�X��t�ZL�{����|��̸����fM�W��M�8oY�	�����>܅�k'7��ɼ��7Ne蔺t�5q��s`�p^��=�&)P�/�9�Cd�N�d��M�/~Z�D=���R��:�n՛\`��g�:"i���Y��h�!������_����޶�a���X��!V{-,�ޝ��S�nl�ٴT�&�B0���_,Y��'=GE��M�_��(�H�KZ�L�Y�.�G4�в{_���#�rd�F�&W�2#k��m��>���|� �(���>�.���%K�����i΅:��xjfh�Ke����*�P�K
K7�����;��MO/��;~y���e��g$�3	�Tk��%�B��~t
�`:�[�Z_`j��]t9V�Qu?ٗ�A����9»���Օ\�� �\�#겑�G��]P�����r&L��gb����OY��9�@e���n1�਷j��$+��۩����3N��!@�P-P�5�	�v���W[G���"�l+����>�xdT�v�vI(���&�n?7�6�=�R��㋬�ÕUn<���Ud��}^�����NOȁ������eKup��ZJ��󹋁��Og�^�/�w�����1lt��
h�5�Cg���X�<o,]*t�Q���$>�ͫ|�{D��{6Ws�I�u�'AtP��|�]	���S�k����JŝXw����V�M*{ΐ�(fAB� ���r��uK�;7��L77�4�	�Z�����Aw+Ϋ�f�y^�|��Q�d�xO���h��¼�i�%
��P��t�J/3�6ޯog;L= 0�дת�^�Pj�=9��
�ͧ'D`��0��A��z芅�fg������`���xj,�~nDσ�q51஦è���Ї�璭�oocC�+-C#��w]U�Ǵϔ֢BN��~��dE��u���\�C�2ix��������ϕ�����|X
�"{����)Ϛ�܋a��D�R��`(���;ض�C� ��5ǆ37:@�q�!��m�|�p=1�'<:ᬾ�G=�F(��GX��НosD"z��T�w0���,U��7�@���/#Jv��c�u�9�L�2��B5�{�k��.��/�q(l��|�#���G�u҉��;Z��Ώx�i,��ж�6{ho�i����>%y͘/{���}(��;U� T��&}����d�W�mf���h��f�w�HVQV�ʅ)�/��Y��N�O�/-�]��sC�6��#a=�b\�>�t�ݞ�Ҫ��[z�w���,�1,�B�C�h���R����U�W6�OF�a��Պ�ގJZЎw+���}�C�H�\�a���ZY2�{9=ޒ���kӑ�?0��2�J�v�����(S��캦зT�����@v�[��?/�ģ:����N�1��.:>����];혔�� Fmd��IF:6f��=����<�a��<����k����|x\'��N}�`��q�L-����b�Nz���x�}tZP�߷r�*�и�+�e�����Z�b+���<�`
�l�w��:�wSrhQ ;�
�����h���v*}�0�^r���1-�F,�u�5%<)Wu�Ƨx��\0�]��܁q3����m�:/�f���1 �}Οpٹ��T�ǘ������dʈ��Wè�>�~g]���g�ʻs���{.n���xr= �)�h��Њ^�cu�ݘ(�$�M�UZG��C��iԾ5(�~5�z�F���k���ǚ�Z���EF��3����yg�u�p���~���}�*z�B;�mQ��I��ݻ� E1g�h�=�D���e�/
.�P�H�[�m��T��/���vp����Ƹ�S6��.E�Fkk;{y$�s��¥�1��]���|V�X�ѳ.���T⑓\ږ����W7G����EG�������|�[�����w��-r
bT:��e!�v ��Ԕ��4����S�u�X�w!G��17Y:�ɦ5ޮ��W}m�o��i�4l�X���������,�``�7�YB�O�Ě/�͓tuw=�E{=�%�_-�/+u!��r��ˌ*#`�1 �˾�L�Pw8HJ���Sbs���NP�>��:gݘ��+�p��J�ia����/Z��y��:��SAU�H<6�ei��Q���N��Q�Ԅ�L��Z�:���ǝ�y�Lɤ{�WǆF��W�e3�3�z!�|nZ��P�#6�儅�BMmX�W�9�ޯ""ߩ�U5Z O���c�J���/��K>ȍ:�dY�oCSz��(Gʫ���"�=��'~q�~�n	p]T�),Ɔ�*T]F�)S���Jd[��%�a�t��G# ������~R��Ɲ���Q�#�ޛ�	H�dm|�n�,4�w�F�j�sSJ��e-�
�k�rH�e�rE��2�A�0�>(�7� �;������������Ю �\f��=�AL�.^�p�\�V� ����1�\����h�>�{mL��l�㽶����R�����Gd��wu�\�k2�M#�F=7�,_Dб�&%�jU�U��_�K���`�G��Wh�7A�	�6��ܧ���Cޜ�UXZ:Q�Hgq��q�3q
VMcm����+3���j�N�3��
��f��j·F���0��B�^v�8��wG[g��T����t����Tu
�Qʝ�����鸔� <(
[.H*~���KY���8��;��E��*0u}r�Ʉ01�ic+��C�.c#���_�T�
� L$��+ ٓw}�8����k|v�9>�jY��Z�au���U��|�A�>ԏJa�����^�'�X��-��lE3���@}Y�k� ���"���;�ge  ���MSu"b���V�O�m��Bx�9�ECr
�t�9�;�Jy[qג�gDE��0�2�fl�mc�V(���	��P�FB��O�9�9^V+�[C0��Ԭ`#���vy�Z�ttL��^�Bw�U�i���[� U�$��í�_��(�,BG��`=�%�o:�T����{aB��-1!s8��R��_j���T�8�P��W�������vUgV�)5	��܈S'�(�SY���\2�\7٪�!t�1��0術���%ò�y���ט.h*.Ƙڄ�қ�1ʄ]����2�����t�δ&�y���c>�V�������ƹP��5�_rJ�&B��q{�Τv�����1Y��W��x�+�f�:�r��v�2^��M�����WZs/���a薎�vV^I���b�`�ʕ�}g��[]��-��|�xq7�ff�<�ĳI�_��G���$��N��}��1�˺�:����@Ji̠�����	����YP���D#{���;����;��_̥I�@��E������Dt�(�>���M!CO�׮*��qC�w}G	���{���Lpl_uC�:_�nc�!x�aX2��P�&���R��0�`�53m�0�'(��Xb�Cb�nC��Jb���W^5\�~�������U�ʷ���)<�\�]�|x/��r��{��u~Ln��%|�}�j��R�>��H��[rZ�tt��*}*��ܪNJ��	�x�v��'U���Z��|)�q]��+��׾�O=_����ʡ����/ˢ�Ò�v���.��t2�Wx^N>��G_Z�@���o�{��8N�Y������ʛ6�&��~����.SPy�owW�q��S(��\z�&e��{[p�4�"���s?7s|W&0Ẃ�*r��uK���h�׽X��(�=�`r�{����� �b*;����|�!�ۊ��N���m���A����3=8�9h�Qn�e�ned�]x�v�X��ԔL�[T�U��S�=Dgg�0Zc�)'`�8%������,u�4N��;�7��;I.:�u�L5��Zt�W$�Y�&�bf���XXp�sg7]�6b�V2��x$X�ԫ��Y�uz���R-�p�@�t=1��T������؞v�+����D9���i���>�h�����Ƴ�~9W�s�2��Nޜ���8k�lqIwFt,De�|��w-�+xU����ò#X�F��v'�<� oO�x�R���c[W�'��x]��1����s�Z9��#݈���7�� O]S�QZ^�kV	�'�X29S���K�ܨW9Rӣ�7',E|�ݱY�A��PB�s��m��4�G�޸%]����CZ7�XCBi�F29¥�B����/#�U�O��8���+;ն��T�5��ʉ�G��0��C�'���=�*s\�5f���:0]TbU}�wb�XL.y0tv����|n	\c  �gt��������<�fFZ�����R�T S�1�A�i��PZ5���rP����5�w��<��]�U�|yK�t�U�zN[8�tl@�]� uD'�Z�r���m�]|���tC����QV��a��얃�qrJ*,�&�i�tK�fT���s���b����j�N��1��1+4�U�Ö�@�SO��c�6_5�Ջ(u�&��p�̽�˫6M���f��W������G;�j�&��u��,l{�mlRPz��Axp{����v��������8W;6nB'�9���8��ًb{��N� �B�t���Ӑ����* �t��d[�"4_�o���Ow��׶��j�f{��1���҂��B���f1I8��5U��[����{Mf
1��Ol{!�z�����9�3�j�_j�rP�Ӹb�P��[���3_4���Z�e���wO:�;� J���c*r��}V�,`�8�w���H�[�m��T����L�R>設�i�j�5����a{��6r,@�[<�����m0Oۊ��J��jJi�o�ůgQE���l��;vY�����q����퉊��n�O�5~6:����ֺ��ڏ�b����󃤡�vE�A7?,:��`��D��G	G��m���]y����g�
�+q,�J�v��O���J���r�\vLh���1��@g��t/x�9o]0j�w�.Qf���Tw�% �V_\�X�c��U�.2�����oi����]78�q��@�f���^��:y���W�	��wX�U3���u��Ý�0}�|i�MVٳ����8;4^����诹�s�]'I;�Ѓ��;8m���:&c���V�C&�/]�I���a�O%�o�����dσ�����G{��܃���@.#��߮/����B|��Q�̬+v�Pj� Nug4	ժ����ml^��Xuu��TjΊGE�Vd����YQ9צ!�u��(Q���h����r݊v���)Mޫ��^�6�YohW���Hhsx���8'I�4f4i���]L5 ��(�v�P�a[���$o/�T��ۦ��[8ge9��"�!I���F6(�*�[{U���]�Uï#}l&��<���4�K�m�-&����d��YZ�����E�J<:���G72u�$��[�7�8ք(���{k�H-(��aDaő�%�.�lv��$v;�s���t�Ծ)��͡@��6�� 5p��3pW��J��I6ɀ����L���=�[o�`�\'��N>蕡�0�!�=s�Q]Mt*Ĺ����9�>��UtU���[J��x�Vm)b�*����n�%��v����\[O��*whC��}�u�2x'�L
%�w��ms���yW���4�Y�Nc�ms���-&�J$L�`vxD!��k+�R�f�h�s�Z7fss�B�egWc�׉��/�S{_ga�U��w ,�j��t�u����^���^����lկ�~��o�W�^�R��کѾѹ\���}P-�4�����U�V$�����w(�V	
�z�u��#z���wuN��kV�w75�"r�kO	V_��u�bv�$�|�h%�m�m���t+���2�}�i�������GR��C���J�g 8�s��=/]IY��L:Ш[��clwh�4R�m^��g\w;��+6�g+�\i}\s��]q􌧒�6A}z@#���]�-v]g,��>o�}���Y��]�oy���[�8������]i��~
�t�����W��]���������h���n�WN*�
2qf]��-�bd*��@�%e'!z��Z���n3�������P���(��9�PdW�	����Wc�^�O�V����6{9C:LKk�,��ֺ[��q�t�Ж�E��rt�L�fm�;�J���E�L�G�v���Z�T\�)JJ����}�@�5�f��ڰ��Ő��7WQ��h8g@�fᶟv���ը�`rB�eet��#��CW}bڝVȚw2��6d
eZ9�֕����)�(Ev-��Q�~K*K���fךW��r����|Ƒ؜<s���J̐�D�a	v���!9[��J��V��y8�g�]6W���1��rގ$-�2��@�tU伭��Zz�	c�
�,꭛ձ��U��g8k.�L9E<��5y�c}�8�S����h��
�oJ�;������U8m�+\�"X�{�EUy������̰0X��i���W6�a�}�]�#@��JJ�n�G�IAT-�J�f��5�Ws*�l��qW^�m�-����n:�Nr�a�I+���#�$]2��]Ut�r�' ���\��r�H+�.[�;��]wS�s%�;�w;���G7#�.�#W;�.S���s�$'u�+����u�q����ݺ,�ۜ�ȍ;���å͹Eۑ��AN�%r���I�������s;t�ʹ�뺍��%E\�ܷwnr�w\����b9b���n������s�(�I���:u�In�����t�0�W9�k���9�s���s8�s3v��ۺ�+�ë�w]w��rwGwn��:�]!��uۗI��s�W9tCu�n���5�sD��+����I]�A�q���;��%�"\㺷 wtw\"�uغE��)�\4��n��ˑ��p���r�������D�$�1�Ѵ��b介0D&AF����4M�k醹6����1�P�Pw)�6�>��h�`!���;F��:�������G��;Z�DD�7�>�ʭ�g-�[�b��G��}"G]}�^ւ���%��7�{�����*9_W���*�sW㟷��7�{U˕�~u���/�����i��W����*��{�����ߏ��o��W�����;�\7W{��z �B#DG�}�g�W7�n��ϭ^��no�}y��OkF�/��y�K���U��� ����������W?������o����ux��W�_��{Z}n{�}����}o&�xc��S�+�=���>��!Q���o}�>������^?�~�~����7�n�>�z���+���=z׏��W�����ڹ_W��]�y��soJ+���ߛο�ך�������?[}�%���8Q�uy�y@qb"��BD}�4D��ڼo�~�ow��7��������|W5|���_�W�⽽5��ߞm�^�ss|~}��ս��\���7��[�����9\�>/�o?�~W��~��U�r3��~"����R��0��f��}U��}�6=�^�<�o�-��O�_����n�WŹ��w�����Ѿ5��|�����}^���y椷��x��_<���Q���7}��^�r�wߟ������p�"f%0ȥ��vU��?��! ",k���ν+���~/������*�/w�+���^�x�����_�w��5�}W?~��^O}�W���{��޷�����o���z\�ׂ�����{���P�~��:ǔ]w���w75��e�/G��ʼx�_>~�ܮ^��߫�~��x�U�W������~-���{ҿ�Z>?U�����_��W��o�r��^�]��.k�]����W-�Aq�~��X�~��FK�dY^�/|=??�>{�~�J�x���������w������7���?ݹ^y��[Ƕ������x�����KF��������/kA��u~�K~���W>5�^(�B#�8؈� ��#�"��ARӯ_��unjS�#�b�����>��#�#s�}�����s������y_�x��r����~����ۚ��v�^�������^^��\�6�^<��^+���_�z�����|�4�W��X�>���@<b�y[淬����P`@D�>����D���w��⽪�ͽ�_���U�ߟ<����/w���U�_�G�~_}~����6�}���^����m�����E�_�w�r���x��s~.��߾���p��I4�G�:�g���V��q��B3�u��e8�Uڦ������kzm=7td酶+�#\yo(�,^��H1M��J8Wo�h����xnb�գ���+������h�U��V\qw7��7Z��C��t��=}�]��\��Џ�1DG��V����.��_w�^�u__�����o�{��Z>��}_��ʽ������z_彯�~|����W��W�����|_�Fߕ���zW�����Ͼ�|k�o���D���(,�T������G�"#E��|�v��ߪ��;^���^�^-���ߎZ����+���x�~�߿�W����~���6�o���~y�����_ͷ���%�қ�V}���g�e��!y�}"Dh�}��ܽ-�\�{��n~6��o��������sno~v�}[�_/��צ���s^�;ҽ-�\�/�~���/ϝ_�x����������[s{���������}dw��z�o�8��}����B�W=��~��~��~��W���w��[{�׵���ޢ�����o>ux���>/�\Z=�9y믋⽪���~v��7��+�ߟ��zZ5��{߾_U�^�� ����^S��W~���!�`�5���1zWŹ�������������Ͼ�=����s~�~z�ߟ<��/�<򹹯��J��׍�.[����x�~7�:��/�k�����_��5�}cwT0���1��#3�r���7�7������-������ߊ�����������Q�ϋy��~���-��^�Ͽ��6�U�s{_�}��k�r��u�\�>|�^?���x��|^?���2|EP������c��/��\���/��m�j~���o����x��_��������Ѿ+��^_����ƯϿ|����o�����ʽ9���_��}k�W��~|������W��|�c�G�|+.���Tʘ��娚�b���[��~/��{�{���oz��yzF�߭��y�}^��������|W>����^��\�V��|������^����?ޯ��}�|^��}�x��|z�����""/C�|]��J�ѽ��i������^*��ﯾlzo��^5������h����{�x����>+��cz[���k����s�/ۻ^�|\��{�:}�\��s����o���ߝO�}c�>�(G��8���㏰�ڽ5�{�_�����ߟhޛr�^�=�Z-}���_��h����=+��ƿ��׿?�Ѿ+����_��x�^�����~�J�w�k�ƹG�����W���G�0G�!U^G���#F�#���Ū����]�#c�ڍԣ���~��!��oO�"�� ��L��Ӵ����7�R�R��&﹁�e��I�O�K�)�p�Y�w2C���ro��we�ᳶbv�n��ٯYk/bz`m���ը�V�z�DDz?���U�k�ݷ�}����+�_W��?<�鹷+�����}]���~^�y^����v���y��oƮWֿ�/����/kF����=��z^6����������D�N�H��0���c�b�^�u��kگ�����zo�żU�w��W���o��߾��^��W>����^��n[�}�F��7�^�}�������Ǟ��Qo���_�_������ ;x}3t�ϩ0�����F��D��z�צ����o���m������W�RW����-V���^����+�\����Z����������h+����Z��W�^*��ם��^
�[����p�"���=\3�q��{�9 m��U�+��}�����[�~<o����~/������_���x�r�|�y������=>����KG?o���+������������_��߾���F��@��t��S����晵H��#���{W����z�(߯���h�����z~��W������^��\߭�^5�s��k�����Kr��������񫛛s���7�~���7�~�|��}�T8}�WF��y�frK��9X�;�����=�r�5����_�x�/��|��o-�/��k������]�->u_��n���^*���ߝzk�~���_�����7�_�żW-�\���Q���������	��;0�����~}�{F�������^�|\�Ϳ>����[�\�����ܽ���_����{x��ν6���ߍ��m�����փR^{��}okG�~^ux���x����ʇ�|��x'09�{"E{0�T;�5�}�{���D1@ G��`��DJߟ>�^����+��<����_�s�~_���~�W�����{��?~��m�n��~W�<���ss_����^7�n\�{��=�Ao���������h[����Ͼ����"�}0d}G��W�z_ߝ�7���o���|oJ�������P[�r����?~��kӚ�������ߊ��[�y��z^?ͼU���~������X���~=+c������z;�Enq;X�a#P�,`tӴ�g8T�柰6���tPٳ�P��3�`K�2*'�������כ@��z���I��u�G�,AΨe��k��g_moꔲv�Z���io��sB7ud�+�7�ђ�d[�����m�S��Pu� o$�s��A�Rθ�;�a��Wq�۪�=%M�w}�l�k�e�v�@��8�|h�}U���3"�&[=�"
�b��}��0�B��A�V{n�A�\^ٿR�����o$�����f�ɉЖET��'C��� ��t�J�bH��q�/��X9:V���w
�^�©��r�Do�[��>טl��\*\\ڍ7sk���}�V�����gA��P���,���X��3�_^��b0��t�OX��koë� ��
+�W6y9�R������Υ��,FE�ɸ�=P�B��k��Y���;)	���4��F��O��0Y���V����mP� ,"�в��7���T$*'3�f/����Tk�qp�?J�Y�:�]�����4�5/㝜�[�&�Fr�/��2�*����c�R��@OM"��`l��O�d��ș�2�(^{��k�^��]�n��6zR���Z�u<�8n��)�v�5�z]U��Job����,���4S�tz����{���^x0�C�ʷ��*�x�v��������D!���)�©7�d�]g ���4�pԦ9����݊*���)�������_(��Q�
�6
����o�d���'��n.��7&r�3�Ey׶�m���ɴ�En�q���=���ϝ�RZ���W2���y�f��� &��p��7`!S�u�#P����m9�� 0������V^j(������o�ɮا�,�b)��J��˳i�eqד+�k�e�P��H����лvV��&�i�8 ��~�h��|X���T��L�p`|�e�T��;l�,��վkgt<�H����.`v� ����	��wX�R~V8J���ug�~ x�S8T��1P��⏔pϜ�W���#Ne@{�UH�R�3�1��[��`�:%.�8�����ovB�ik�A��%�9�ZF;G-�U�)�aωH�w3��`<џ:���� _���T;s��p��V�Hƨ2��m�m�����e�V� �[G�@:����}_Q[H\)�e�ȗ�Zyr-�� ��F�NQ��Ց��N(%�+�$ ��Q�֍��P��s1l��_ԹJ�4W����][��1{���WR@(��f�<�ʌ
�'~`b�K_t�(p%�g'A�3N%�c�]�&�YhDn	*۹	ʹW�`�R���iV*��z9w�[�j��7G*̃�� �Q2U��V��y=|����ƴ���-�3
���*���!��ɣs���Rb�[�J��f�D&���`q^=�5���;(�[}SL���Y�������ڏ{;��7���@:��%�2��q�NO�Z�k�֫�s���p�U[�k��(�����]�畼�tM���JO2D1�
l��D�׷D��k�+�~ұ^��=ӹ�z��l�GQ����- ��ӡ��@l.�'�fF7 `��t�|�H�7�䡗���85��lg7ڕQ�-��_i�Q΀��nX�FJ��T%n��46�t��q84���sFq�/R��$w����V�r��rkޙ:Px�|���x[y����<`sg��4��:%���E��_ӹXȪc+옠�}s8��d�ⳕP���l���mD9���ns3�=Ʊ�+�>�>C;_�N�^_[��n �x��J�8���>��V��cۧ)&;~�;��/p34��3�l�i<�l)����Ғ�B͟���
�<�Y�;�=M!�M����g:N�Λ]�M�����n��$�l�H5�G�_�B[�
^hb��݊�ҳ.�U3UT�p�5}��D$�#���oN
�v��9PB�@H�09�xҹ�^哝�=ƞ>l��\8��Y�����{6���)�}��,��1Ի��A�����n����;�k��j�8+'�3��1���po�u�E�/��K����7�cM��)�n\�M��[tN^D�r���q���R��I=�s�5O>*f�S�U��Z�5W�;�x���$o���P��:_�m� ƓVW;�%ۻrX���#�#�c����WJ���GEߛ�S�\,J<��_�=�C�U֦ ��O71a�Zr�:���h�0��$
�Ѳ����M��-��Q��܁(eb�H���������)
�q%���&3P*'�@�a�汁��}����7�jڝ�f�VZ[ȃ�r�eΈ�ې�2-�( ���I,vi�������iɹ�<�==�<��·�n�p:.:cx�ݙ�É(�d��͇��M����,u��j�5�/��,>�W6�̚����|��N�����.a��@�J7d�?7tx�k�L`o�/T#�4�P��w9�|��\�µ�V�W�3�}Zx	UQ�]�����M�{qM��-f:�7�eR���q�4a���\�������>�*a�_ /���| �`���*�&:w������w�5QW�������̎~A��e+�2���:��_�Ϋ-�De�w��&��6��,Ɂ���
�a%��+5+�M�����[z�=5qP@�/���۲��d�+Y�:yR�Ӑ��=�V�rP��4.�u>����9j�QJ�μZ��1�\:��.�Wme����iI1��\Safi��2b�WjɊ=��">;+�%�m�>�U7������C��qI��"�3�*�P�	��R�꯶�N�􄋍��b0�ٸ��3�X�ʯ�Egܨ�tE+���]9F���Jj���t���3Fz!��)�&��eB�R��F���)�#�Jǒ2;&��]DE
3-]�;���*Ӱ�"���T�;(������(ugC��;H�8�zp}cUFc�Șηj�>�ދ�)dJ���<��TdI�-��7G�xK<7f?��*����!Ҽ��������7���@��L�V�d¼1-ى�d�C�Į1�
���J(ˁ5nHwJZO��C�D8
΃�����U��P������*�yY[�[
��z����ہʅ[�2���qV
�^����7�n ���O,	��; TL��`s��e���No^{N����@�ɒ��+�:;�畇!s�9p� *�z?=N�7�X(�y��U��nxp���Ąl'+����d�&MF��?\v�b�qS�����q���jc3
u�=�I���Z(7ioW.Mv\:�-D�+"<�X�U�=sE���ڧZ˧�g,��H���_nc�gv	D��B񼇺��c��T�,e�6��ʺ�Ng5�����
_qW�wuW.,^�p�{�š#��"��obb�α��[��������%@o�Q���X�`bȬxS���S�)1�o!��ʈK����c�-�B�M�fJ9�2p�j�&�B�^W���Ե����>��
˫��Gz�Zu���~��Y���	��6dj��ݴ-�}��~�6�y��*��A��m�����@y܌�Mu,֘� �ܠkU��l:����C#pO��w\x�zz������gk閬'+����@ml��@|l�Tjv�[�_f������@�fp�C�Z�6���Kd�˼��.�u�
� �\+�2gO��p�DIeٸ��W���;�eCj���Q�M��K/�tb@�.w)�73@LT�"��FL�z��Q�S8!�9���ǥ���JW��F��K�����j�����\���m�	��Ӿ*�i�p!�m}5e�����IZK]Zm�l����C�
����f����
RDY��eB�,5�	�z��h����
�]]�!���r
���������ƝU���H��M��m�f�����th�	*�e�Q	ʝȘXkn�T��j���m�MO^+��/�-�poɐd▾�r�����2evy�R�2���@X�5�vŶ����]���� �^���f'-�����D��j�Ά�k�^�KW&_7ҦLR3���#��[i6��T̜^����wu�&=�h=�7`h��tED2�"ԆP��aS׎�<��)�x�Q���<� <���߂�AL�.^�i�Ȩ�U
�б1�2�rw�| �_Ҳ�E��$L��r����P�U����'熾�*sۆ*#��pI�W*�J���� ?�/�\M�\��V9��#\,xgՇ�+�%
�%�\<�/.cv�{��m��	�k�����zJ�B^�*�׸����]��xa\d��Q���f�a!�V�1I���ś
gn��<E������D1��Uz^	�聚ǵ�/,��V+�gjn)�Ǿ���רf#�U�<�䪡��X�<�a�Q�+�I��H�f��8�|�u�8��	ON��i��5T�T)�����l�4�޷Xo���G��:r����O �q�HR��G�B��&�V�g!��U�w��Y\��B�i���=j�ȇz�ln����,B�U̓�([�������L�+�������S���glP���mbV�Dj,�'{���ǫ��6�E�IՃn���F{"�QUk�b݀���3���`� r��f�t�׻4gw;�螞ћo��M�zĉv�G뎹��5�7�-<ۥ4/��A!	��8�*�m���t<[��hY읜-M���se��q���v��杀>�#����:��zi�˛Aww"p�ۀ�yw*&��`�C&Nǽ�wt�ѥ��Y�>SV�wk].�S���3b��zE��m�����Kr�eq�{7C[��]*+�����+�Y��>�O}}�π��m]v���˔6��9gQg-:��_Z����Vh YW3�
բ�6�퓷%޵R���Υ�l|1!'
yM�N�i�2`P΀��hl�L㫥�jU�m"rah%Lɹu�]��m��+r�Q���
,�ڐ��7q�v~T>�}��t�O0+פ�RN{�|�����X��:"9B���d�W�H�K0�
/I�ܔZ��+����;:���%j��1�����NJ�^⾅��x˥��i����gT��fZ]��;�om;��O�����}�`��K����N�4�&Ҵ+ f���8���1HQ�Z�͢(.��u�l�XN�Wc��H��E����Suշ�;D�n�8���;���a�Y�C�6��=�4̔q�h�!Au5n8`�o\*F�+Zb:�1����QP2��2G�.�Q�ig,���#�Z,ј�C)��V��i�d����l�Ws���x9��w8��1naT�zm��V�Y��(!	?����9��Z�(:꺾��e�'�.GnVeu���.��8m`��r�u��ÿmDb{.��n���	��y�b��ԬW!��Xm�[�b&���&�T���{�Ǭ+��KE�/��h�V~�eXp;j����B��9����������Ęr�4��G�T!�Wc�i]�;������1݌b�ڙ�(�x�'TF���ڷId颹#��A�,l�M�sJa���A����Acz�.����rG��V�goN�xw6F�q2�s��Nʸ��T9\ �K;2]:��wHM�79ri>���;�xU���7j����*���K�n1Wj����2�e�ʼѺ;�$ȟq�PYl��bǝf��O{�a,�ʾɳk:@�*�]Z�F��\�f+�t��ʮ��ƅ�Z�cV�'���o���|�b��c�S�f�o�:��д+���m�o�Pq�³��Ы˦�a�Z��b��&����i��pv�9X2��N��Ґ+r\��Tn��˕1�z�
A.�`.�/�D�Tr�8�ҫ���H��6���K��GV��rF2
��������fv,��f��ȹZ�4޻�B� 4�:�R#Ckg+"��Iv�xYz�Uq!�7�r��=�m3���U��bv2WP sim_4w�K�����+5q@4u�Hީ��Yϕ]S���n�7g9"5�X)�wA�j�s��K��;�]�D�h,A$Lnt�s���0�s��� ιs2�\wr1N���w]s��.ss���sq��d+�κ�˴�w\nú��q���K���]�û����b�;�RTw:�	F�v;��'u̦��3�q#��L����wsn+�D��M�vw"�����ݹɕ�Ȱ����)���ܛ�Wш��w#r܈ƣ�+��"ѣ9�fE�sva.��v�&a�B��.wu҄�C(;��N��E&]�"R�U�Ld��� f��Q�l�&�1T�I]ܖ#"k��;����A wr]]�n$D��NuC@Gv�z������w~N3�����}�-}�@��ٷ;ݗս�
���ʆ�3
X�\���� �3B	��q<w����o,i��_W�Dڛ����EU��&��\7�x��B�=:����k<xJ��������(>���J(�u��SC2),P��X����E�J��!�����ʒ�Gb�~��*yo�E3L���ny���O�ћ�B��ъ%���hp�WP���EtSNg�F.$�{p�qy���ޮQ$���g�6��W�_W�Rv������v'���O���`��S�cNy���GAD��:������.1��ǯ��\L�|m����9U�<�7j����ajܽ�8�vJ�10�U�Z;d.5���j
����}�^����g{a�v�g_ *�],�5U���#��|�Kiv�|���4����X��܀P�0�1�r��k��f8�A�9�eWD����*���1�so���P:��f�%v]c�~T��+�#��O��ksS�������qb(T' 7����`?sf��X�	1�9���w{ؕ��4���!aP���i�W�j�K�	U��� "�CuL<G*l��&ˉ�x=>1�X.]N�e�ِ2<95@��^`�g*��V`b�%a	ќ�W�p����$�*�DJ��n�N"�`�5Ĕ ]V��w�"2��<�6u�^�zZ}}2�����66;7�u�!N�H�P�1P��u�� w����,R���lg�)�����}UU_n���/ ��~���KX�J�;Ģ��Tj�]C��ʽD�X(�L�0�˖o �G�Nk[��8 ��w�[X��4��΢��ʾC<��W7T�W�ʅ��j��"����v�cIXUQNa8b��3��
��*��;<%�S���ƃ�����rPpd)�]�S�<��o�,��'���%�T��Ę�Q3�D�����9˺`aS�
ps��R�$�5�%kNku5��͎yh}bxo}��)���?E�k�Q��9�] ����m�M+�%��(>9�G�Ų��cUJ:z��4��B͐%THRX�pB����5��(\�Q`z5�D�~��^=��G)Xz4��iL�����ţ�䏲�C)T���l�:���dE��ْ/%�����(u0:�i�f6*\sO�.��=bh��0����mn��
^Mi,\F�E$G#6�CԖ����	*�p����3��tM�`>$7�ۜ�v���H�&y�.��.i��nY0�Ah�l��]�R"`�L�{M\���M�9���Y�=�j��
�ޅx]�z�n�}V�k}@�a!YN�n�i]��R����|��%�!f��@NB���v����}L̈́�1��':ヌ���Q][���,�0�>���=��ׂ�N�9���<m2��f�_W�UU����T����`����O��Z�����\j��r���WN¥O����^M�V���[�����#5�&8D��[4����xX]w� ��~���7%?�3�}�r�v�H2�l����-�F
�sԕ ��Z�9���ô��R��7۠�OwD�Ap_
� ��n.���.�Ru��_ݰ���4���T鶪�0h� d��/p7�n�{@p0P��]����,Գ�+��N2����T*!��3��\,Z����t�Mz����\0�o�(+Eh�J�p��xh����^_ظ3�+o^f_f�X��i�om�GLhOn����
�qS�l�W��ߍ�WQ���o��>���+��Ƶ�  ��V�"V:�3��cw�*��A�	�c�T�ܗZ4��QC*�k��0ޜ˽M�'r�|a3�@�x�W٩�>B�uKer��ŵ!-s�y	��n�E\���ۊ�m;�q3���ޙEY,�7���U�ƅ��H���%��f�:�%��g��d�"B�������k��`f�����MM=��ŝI���6��L�o.,��஺�:�Wg�4�2����ď�c:�0Y!f�|�s�;�]��pO�zuy�e�޻�H�.���͂��ʶ���Ńs��">��&��Wi�s!@�ߚ�+��K�(	�5�C��xJ�J�{?��x���W�A�qt[�	��͎z��w=��G���p4B���g���U`�L q榺#e���&i|6::�e�|��p�v���Jӡ�/~n�CӁ_Ҭ��_�˨{.�� t����N[�l��uE֦���nb�:H�Qe�0T*�*"[g!`!������" ɽ��/	~���8�2����˚���r���Mn�+UP��A���DTE��()*H�j�(�CcyFk��f�뤬��(|�'e#��+���V���F.�\8����r]w��̘rk��W;�T6[�:��+������}7LE}{$B��R��@(gH�Yʝ��s?=&�&b�Sػޮ��P)�2��]1r�)&+�U[��#��O��Pf��]�tq.�<�Vը�70��J�1�\��m@��mQȒ���j���VaY����:���+�ý����qf��N��/�0��n�C
l����#�O6t�X�ϯ��įj�b��ǲV��2�O�5%}�/�N�A���� �x�oR]:U�D��ʐ6�F)�ߏ#�Sݚqk�����jRSol���[{����~�vI.��)w��T$kwu�]qh6����De���A[0N�ô�V�&�>�tg
�J�Vom_]��UW�_W�K��.^�����x<y.���X����k���l�٠���~W'LS�#�۞p���6^� ̄�R���u�zb1��J���	��ȿ���'���t����.:�6���|Ƀ���V0��v}*��*�g!���~�v�չ��ǡU�Ps�nA���
N����a��\�0��	�`��SY1��@\���f]=}�� ���=Y-��b�<�S�zb�!����ૅp|yg���g�	iWU�̖�j��e���h{ո�s<0^>�|c>e�S���/��Jn%LBۉ����g�GN�J7��gs(���Fs�]UGPX��v�uu\t�VSNe �4��!GH4 ��]u���Q7�89f�S�J��H����')��L�
Ǫ���<�������I��T7��0������L������3w/��	��t>5�71����°�k�vJ;R�e�=��G�X�H.���0c����r*��F��1�!5����{*��+UI�˺���U�j��k��)i��[}{m�#}�Z��E\�iZ�{J�-���rs��-c��[,w�x������(xu��Zb)�q�^L��s���@Ύ��2�5֫J׵�<�@
���*K������Y�DIҔ�5 r*j��DG�V������Q��c��u:J.r~D	Kiw�~��I�:W��=m���G���ƻou�mg4����f������I�����T����=�n���/���h��*�ul�]���׫^��\�xS��dT5��&���o�T��j��j+{�3��SOv?"�Պ*2a3�wHo�3��L�)̰�!��p�	�2_��5��ٺ�X���B��\M*�q��Uk,<R��Tqyץ^��@I��'�}���]�D���y>�:�E� ��_2��c/%�Us���$3�G���*����@a�;Qs�Ps[��UwyfR�򫄭d��Q�p�G9#0��^�\$*������>�i��wʠ��"�B�\�G]ݸ�p���k/�d5�Q��8J�Y��	WB�k<J�V��S�=��vw�W?������5�1��-�uw�ѷ��u�����g��Y;��"�A�jy�އsMu�8$$j�P�s�~�<)��j�tƋU}z3����W�&�b���y����zX:���tuy��8���'[�%\|/��1v��e�\�8֢�v�+���Fǐ[���\OO:�8���`�޺��h��n� p��\D�W���f��Sq���:�C`C�sG�*2���[���#���p���������Nb.��7I���*�Ai�Swe�W4�汸�R��I�C�"֙)���"ŗ ,��T�2�84b�Qc����c9¥ƍ4�{YӝY��SI���zZ�1��*]�V.`VD��2xD���:�����Һ���|����;T�t<o��;�L�ۃ(�Oźd��6{&'BS$FA:%q���z�el���]h� �2�B��}LE�vtn��ĉ�"3����䑯�ltF��p~����$��V#���L!�K	mZ(��#�l� �́�,C	h��1ûogVF��qK�	��#�-�ɨҴ�9ŉ�-�SG#��9������	�S�u=Z�0UL�c�3�r������p��κῸ@f2qR�W�;L<SX�vwEvU%(��\�X�ː�P�����c�8{"��O<����x��|��{�y'aL�[�{�:�
��;9-���5�l��P[f+E�n�8}���|�!E¹��p.�\9�μ/@6�	ΪĹ�ۑ�m#�m*͙�;�P�#�%���i�;d=j���v@C/|�Tٞ�Ϋ��Ӹs��$ka=3IT+������"��lۊ��ovj.B��m��F�(,�_VsXZ�õ;����-��
�u��-YXSY\�BK����^����#u�����5ft��7���0<��FCx+<3�zIçg�gq�2�V���(���Ɣ,���, u}����TG��n�E5u����Z7>�u�OH3�c�f���w�ZG{�O�5|]������S�*-L!���X���ӷ[ݔ3e��k&�2k�D�R8?���U�z��Ο�,��:K����')��ٌĂn��(p��d����i�~d>1u�bL�i/i�>ɘ��O˴�g݉͹\����<���-�ǰ�����ث�d��~�r�m�v���Ӿ<�
V�>2�4Gm�l�}t��!Ĥ����|r��5j���X�����ş.��H�-w0(����R���9x+O���}"�����]���C��q�n%.1�* :S"��7>�!��%�ql|�eaWxq�-j(��&��'��������	t�eW������*~��C��D���eb����5�9J�}��a߇^S�h�84o>��8J�\���+j��Ͳ�你7�`.r��w�e�B\�7mɯ{3�Fxv�T���*`Y�2���5�w��ە� ��6����|q�k��_^�q;~���{p��k��4�!ڼ���5�Ә����]�3�
K��L��}h4-泷��n餇P�}��DN�wV�lt��P ���\K�b2�����"��/dLwI��r����G�ay��X���o�O�+�_������%R�Z0�+�Ue��֯���������VR��>�9��|d��&�3�S��_CD�=���4���aB���0��3��^�y;s|7P+�J�h�,h��Jq��y��lW����ϧ��%y��%,u�Q��+�æufm9j&y�Z���˾}�0o�� ��!*�`Z�bx���܁���t���YV���<7Ky�Dg.Pˌ���.rwLF3ZT�cּ/���s^Ty{kZbk�.z�L����1�8�X�����NyT��lS��S\���7��4R��jg�ɰz��F"�3�o��'�|�	�yX��3�T��6O��V�+;>����7y��2�sE%
(����Ƨ��-��(�}�P\�ؚ�ֲ"�#��M�#��ҵ��A@��m�Ҟ_���:yЦ�M�L-�LJ�+�m��;	��Ӽs�W�ndvK�ȶ8��ww�e��4(��������B��C���O��|��n�˦�F��D�:�s`����3^0��nQ�^bdz���������{�������wJj��]��Ȅ��'v^f���;cx�؊�l���0�����_�_W��Ukz��>�'��FZV�ؚ�+�<�ƣj-�q�.���[3\⯠,�'v�'��'&(��ڛ�LV⤚W�;��8Ɋt��Z�gI��C^Ԭ!aO�a:���M�}v;����wr��MpA_g�
d�'����l����0e�+�S+"56cR4.V���p���4����b��^�}ƕ̍���O(�ԥ��к�0�X2�'��k��Y��T�U�����x1�7ֲ��R��n�O�I��<�쿍,��
r3�"�L�m��p$�/-)���s�����Fޅq1Μ���}�9�sǗWsg�(�H\�;ͫ�g��uR������-�<i�Ⱥ���ł2rVV[�v���-���F^z�ݯؠ�Yӊ.3�.���VQ�|����.[Z\E������P�r߂�|�W�b]G��	�R���Ĳ�m�J��Hu��a��6�*+U��|�Lj_�Oܖ=��u�g��iV���ܘ��uGy�:�h��lk��oV�΁L��EnҺZ�l�Ӻڃ4,ZK�![z��#��
d>���֋���SW�u>����[�~ܝ�5��X3B�T4��V�W:���+����3��$opE5����rn����M<�
okT�Y״��$6G_8z�HK�h(]�uã
�岚}GF�ڥ�)�]�U���&\vOPe%�y����<6�-tB��R��\��G���GH �5�6��æ�S�A��	t-����X�]ʵ�j^��5`�א�b��F�'xA�]�w�O�'{gC	[��t3I=�Zu�"�3I��;�Ii��.����-�2Ƽ�[�rP6ܛGs'=�Sw���D�pTS0�#Ju���|�#�,޽ݔ�g2J����t	���}�hqut�;�t8*j�N�6�{��)�(��`�e'��%&���s�Иk1�k���|�N�l�n�Y�Yγl�c���v��孏3��o�l����"��T4h�07�z�4��4�wz��W��1t�/wrn>-�^Բ���u�T%�Y\�$����L����Q����Ϸ�6=ܧKB���Ll�������mC��Lx��1.+������{-b�1�θ �8%a	�Ϟa�{��(�w ��gK���4y{��H�L��G���Q��C�+]���QCyX�Co��*YwK��M�H`�l tԨ�elĮ��iU��ӡp*k6�eJ�(ӼR;�m9�K��;�Ԧ���.���]u�G�j�����\�}��N�-�c[HӰU�guVZ0��Z�n�-�ظ�F�+z�����
Z�Ujұ��&��#���{j���Q+��c[�1���|�@֌4�^�*��u|�Ϋ莳˩�VJ)c9{�I���7S1���5����CF����Nt���+�owy��f`;{m̻*���j=���x���Z���t{ԾC+�����	ް�ퟅ��ՏyL��hxw}"�s�C�Jf��*@�Y���t��7zU�Q�I���F���n�2S$�Ӗq-%���l�W0&N%��Y���6���8-1y�h�%��3*�\h�J�e_��H
�Xr�v�Ӵ)xu(|�񕯡�4�Z������ �[Q�9��/��ö�<���r�6�p�.��������\��~�{�.=��!(k���a΃v�eX����R�X��+���EV�+7\�S���C�x���6����n�6�P�I�mi+3�~ړCf�ȓ�g>�5MbY¹7.�a��D����f����7�O�1i>0���d���]n���r�����[�נb��PJa�sCb�3.lK$��L�1!�IF�wqfh�BE��d��2)�&d�KJ��H҉i
��w]�w];�s&LFI	0���M	ۻ�(d�Q&�e�n�rL` ��.qݸd�w\�H("&�D�f	�[�d�&Idr�A4�#@d�d́����l5ݺ]ۤ#��D�0���2!��211��0̚T��\$� �"�he"dB!���ᑈ$!I9�F�ut��I��2%ˁ�3��"���'.CH�i2J".�%��N��)�#5�y����ɏZ��:�����;���;�R���'R�F��j�*.��ڸ�|qV�|D���Q1��C�eatql��UU}_}��i}�7��P��>�zjZ|���#�T9�(��>{�K�ug;ay򍬎�w��f��U8W8M��Jڔ�Ͻ�3U�i�9�J��9�ޱ����gkֱ��0z@�4�/,�=zk���[��r!��:Y��u��J
��}���ɳ��=]A׫���ݿ�ŉ�g����dRs
kz�ՁuuMP�3<�ڼ�|�~�~���tVm*}���w��i]����oGW�!��� s�}�2�����+�����f��wVl�tS�ia#xՁ�s�m�K72��b�T��}n5n���e^�Xz���M���]/��,Y�ڴ�Dǥ*Տⷺ��o8+�NQ�nYWa����I_S�O���t�vc|�せ1oK�Z�@O4,���Vn���j��k���e�}q3���S�qgC��Yc{2ù�����q�edu|��*f ��W����N�^]\�%�5"l��R�.�����~R�S�7sUjv&��6���L�r��Meg<gM���h�N��ٔ1-aZ��\�L���$G�{�B�ۂ��y�l;�-�T]H�ؕ����op���OwR삤�R����);��ڃ2�����i���۝���_UUUUb���w��sf{,)��?cǶ�v�U��'��5f��߱�����+˧P�V�'�|Wm|f�\e�zg8��HS�%�m�Su�V�9.�Q3���:�\[/�~8��+��^V%R�F�A��ai͒�/���p�P�i��VTs{9}cn��ʀ����k:Hkٔ��׳�Z�uY(��0��w�8���D=̚�oW���V�\u��x_&�~ń?iP�`�s��uQ�1V�ɍ�\���C��q�v�Fhَm�uA��q��B.e����}U�Xqv���>c�_z������:N���s����aM��g ����Z��\�֫�8�,�W�*k[�M5�\IVa7*S�-l���Wr���[�A\������D�>UW;�j�],��.j��U/�B��N;c�n!����|l-�L:AB͛�)D�w54��a*Џ�^����{���%q9~5��-#*e��a̚��"�i�3vG !koD���L���6���e�s��fH��Y�+T$��T��ͺ��ֱ%0�-�e��9H z��f.�wa�Y���� ��0��uN;�X亰�+iv����w�#����k�8�����E$�^�8�����a*{0���xF�n&*��4�w���h�m���}��)}��w+�1�LS�S.Wa��t��hV��!�6�ɱ�V�w�n�S��̭�ު�v*��(ݽ�M��t�X ,0��t0r�B�V���,+׬,�1I��.wP� ���s+L�^]JQ���.�.����1=�
�%�ȭa��ÎP:��x��<��	\��:��o�ʝ��)�ʹ|��_��"ul3��WD�v�� ���lR�NYS����L�̓4��/�0�wZf�0�h:�ˬ�)��~Ħ#��i*3�!��p�����NGbcs7v���vn�R@I�,ί��r�ƴ֨1�M�j�qq�U|�2k��c���?T���t��S$@��9�g#}���Q�<��W�
��88��'&Z�Ҷ��BD��b��B��\}7��prŝg��u���S7#�)���*�0�6�㭑e,����y<c)���KZ�S�7��p��.��f>9�R���S�<����U�5�{���V�ﾯ�菍����J�`7>��_7�t8���U��m���6<��}C��{xd��=�e੥����{�׺?3m�C���W�Ƿ�zOsa�N�=&�oܘ"W8�|��{���S]���BUAV�����hDC��s&���ӳN-ɱ���~Rt�����j��V���'Wgyt�yȲ��d�ͧ�FW��R�ڱۿcj����v�ƶ��7|l%;���.��4�o��c����z�?`9�n&�57�k�P}ܣ;�Ԍ�fU;������a�V��ز\�`w9X�]�&�>�\�Oպ��|
6�S]����oo*
��oW�~�H���5Q�93U������D����{D9�:X	�zvee-��py�����p�)����"�ᭁ&�[����q��z�+1�9���9�-�"���YM�M*fC��)��G%_���7X�#�0���P�U�����}
�&?m9��H�$�צ�\�E�;�L������f��ۤ;����S���Ү��+G��ʉ��$��7n��s�6u��K\f8�@ڮ�����S2=Ti=�!��nm��v{;�s.S���j�i���=���䋼����}U��U�����m�{���E1��2�F'#��k�5a'S*H������=����A������Fc8��R��ָ9����ȵ�1�u��h6���\G~�p[{pg}�V�/'+��P~y�o�b��f�Ь?���{Bin>�r�dT�v�M7��:��}G`�YoU�*�R���;�s��T�H�{�鐣��U�tN�ޞp��my�[S�6G��s��Qokg/_N�8��\��m�.i̯�⊎X�m=T����m��7c�T83��%{�x7�˞�s��=Ǫt�9>���>�j�[���ע�˯:�G���f����yY�-� ^
3)�_Y�����'�~�uzE�<�-�k\b�wv��a�����Aj�D�N�K��Rw��F�يf�� DI���rs1����!Y�\���]h�[kB�,؉7%(��joS�f�cy��E���ĪT�c��9��C��7���.�YR��n�<��u����Θ���ss�ᕰ>��N��%$����z�㖥3�d3�5�cF�a7o�����y:�(c�n��$CqD���u0_Q�B�ƕ�\�ﾪ���&O{�O��#/��8]���[�:ʸ�	`�Y�&���΁��Wõ���q}����u�T7�㌧(�Cl*�`�XC���X̚�[��yΦ-%Fl�N���a)��Ekv�����V�Oԥ��Lٮ�i�f+NSh�TF�8��)e��a\�k���5�5�W�B�}��[��b��Q )0r�U���Ú�3�,{
��-�g#���iˉv�q�P�Z,�����J�bX����OM�/���Ȣ�h�����U.�G��V�咻\�Ҋw��pi[;8�i@�Ю'�+�r�o�:�*��=���.aeO�t;��r�����h���l��s�u�mӑ�Pq]E�SE�\�wOb�R��[���/^�����Ɨ��ܚ|/�͈r/N�A��s/��gB����]V��1F:��1��~�X�s�����U歝�{ǓN���R��*-�B����K�6����툻.��F�jr:�^��� 	�<'.�d=���2�޽5zE�e��}�;�_k��Wv�
�K��(ڹ���M��h��4�dN�1G��;��Z��ٶSq-�	R]��Fq{O��M>y���}G���������z �`w.���!yuN���d�el�����	[�{^L�=�DL\7��+�z�U3�=޼��},f/�֪�+��4�rQ�fvެ֐���k���1�UZD���|�"��h��Y�*�N=�X�r���}��}J�{Ō��TN�wR�_���I:�eG���v{��K�ъ���&>n��A.�	Pj�Vkov�nW^弗V����u���x�kuR��6�O"4�W�Q���9DڕYJ���e���iP"��1۷����ˮ�����u#��9���X4��/zS�y0�w�ɚ'�J�й�0>g�?��%]�����v����2���;n�YK���&���ѻ�E���4��ڽ%vM}���mC�Dr���ٞ��yK2�={N�B�{�O:s�`2���U�;��t�I�����f�;�S�t't,G�9/[�|}y��@=�/��`[ܧ.���C*�l�mAZP<��+5�����lkR����	+��ᲖkD�s��K
�,��)w01��}�U}H�ڝ^���	==��tz��?G'��N;��tJ�/����{pW(��2^��ӭ�R+q�������u�%B�q�m�6j��+H��Q�y8Vj]܋�V2��Zμ7��������	����d�%�(k��<��k�hY�:q�z���(���'�Pg��]'P�w���f�M�x{Vr6�9�QP�*��E�u�1Tiy/��[�3��/k���s��].Ke���w�P��Z��Ai\9�oi�B��6/���x��U��cq��<z��v��MvKq�؄�*�I�L,�mN�Y[g5�.C����#����-X|�U�ҽ���vC���Z7�\��LJ��,tY��aa��z97MA�蟢�*��Q��:��>���_9���Vj�uΰ�$!<��l(Y�&�Q<���kqT|�K\v�	��S����n�3=��L�U�^�]~Gא� FN�$kt��ͬO9�˵��+����+�M!�}�.����r���8��J`�h[��0j�{|��#V��vΖ�%p�:
�xv�ԉT����IFn�;t5�ܐ�O���x�M���le�#�E�W��>��;A�c�OQ��V��e^J�0�-�7?}ws��LVhQz���R�]V��GF+��hsCy���
��SN��O�5�c���2��ٚ�}�S�Ã{��T _?�_T�� +c���O,��b$�.��ʎ68�!՝^v�L��\�$��M���>]up����D>���eʥ�9v�]�EG8a�T]edXX�u����X�U�HS�s_rp����*����Ր�X��xw��j]O=�4�*�[=�%c)w��'���������K���P��3� m��~�����w׿e㨼���v#in�N�bP�wu�>Tsn�=Od�7c�\ʇ#��+�z��r�cv��ҝ����x�뢳����o���՜�{�E�EC�qË��F��R{1���^�߈�<���"k��[�i�5]�lo}k
ۈ/0q@����{�P}�3�Y�p���c�����f�2;�Zb����vd�Y�W'踫���di0	���*�\쏢}��{C��?�*g^0���}�^��-n�z����:CY�:u�1gR譕:K=p��ğ��_W�\�]��Ç/oS�8����^}���z�����ik]��ː7EF�1�4�d�S9l;��Z�Y�_Y|�#OLa������o_�t����Z�=:���(�xĪ+�m��N�]>URw�h]h!p*�[����	b��	oJ]t޸ڇ�ݍj��Å�m�J&���]�N^7U��B�W��\�V�8i%z�ocr��>P��%s?`7=6>x�����cy{�k[�D�q˧���s}����&�#E�edjlƤ+� ��.�P^T];|�(Ðg�7��n~��UV��w7����R�;��އ�Ϣ�8 n8.ۉ�~���̿���a��˭d
l�J:�>�2�@�^��m��TI��)�>4���b�,y
�:B��j�����?rf�}���sHT��[��S��M�R�n�̫[oL�ذM��`�=��X�v�أx0�Lv���o"��t^�/�(�du�ŉG�)����nZD@k�]��͗��k��,Cr#�yS���;��Qd�����RUO�\�N19�׷�(�g.�@�[M���b�=���r�l����̠��Fw2�S�].���,�V�9!���.5{����뚻�h;�4H�*]b�2����dܬ5ի��e�>#"]sN�:�x�<�m�m�����b�Gu#sA�a�c6��kP��m�%s���YЫ�^����ݚyD롦.��N�rvz��(�18�b�'.�H��X�ܸQ���E�z9�u�hέ�%��+�-+��[��7���,K���o(�IjJ����֦�3�����S�6�������5z�f;؂�4}����톌*��,y�^��n�8XV����Wn-�Nn �=�Iyy-��)�b������U	̥��E/�1}�(��r\��n[�
�F�`q��@�.��\B�}�y����R�G}�N�w��ϡ��1��4�<!z��;K�4`v�Toz�pьTjqt5A�s;Q�{Z(2+�����/�"��jS}
��)Q�.vpdj�+.]���ᇦ�ʃ���Hh.�C�|�!�CY+^�a7!xs�u�35��J�IX���)��3����#f�����ڞ���b���B��t���S2���Nt�ն�n[L�P��F��c���*�^V�]z6�4ƪ�&P��c륙}P8R�HZ��¤6�b�Nw����:����E�a��wx2�uՔo�����\hP��+! 'v˘��N�#&�<1�V��k�a��4�9�gH��N�R����A�+^�3�F��BJ�+�*HJ�To����k�5����w
͋)��1j�;0�)(Ai�c����c(�����!��s�7{7�zպ/�<c�0�-Ʉ��d��)9�l���vlͦF��������(=�n�+& z��.��@���`ղ҈�Ajg5+�`e�犝or�vo\��;᪵w����A�K��#�Ǚ{X�%:Cx����xu���ؼ�z�wsXg=�\�q�Pr;G997v��x�V��ʏfd����\ Y(�4���tn�Y�LEF޾��s�FG�ګ��"��4�5�klc���cM�7z�������n�Q��NP�Z[r��	9�>�2A�h��⬖sR3�0�:9�	�o�	�액m�XǝܱT=��[[�Sǔs��7�9&epE>���5YNmѬΒŪ�ǧ W%ώVA{��=ה1!��-�\�0ᾷ�f�ܮZ�c;�Ɨ;�W*��j`�5��i�VT���Ŷ����v8OT=l �M��@�u�u��3Mɐ�b�$E�{�*�y�D�2`]{H��,���K�(gd;����uVgw�tM�X�O�]�P
m-��a4ke:���#y��ֲ,�vd�!`��Vs��$Fg<d�C�S��5�B���(
P@��;��n���s]������4���ӝ4'.�s�F��ѻ��.tطw$ٻ�2�2dCDc �L��0$���1@	4�8�9�Ĕde2� ���\�LL����PHc;���PR���2!0fX�����������!�9ʘ]����8!;!F�#H��d4��`˻�D�dF��'u�J�ti�"d�I���2B��DB�E"L�8�E�!J
Ms�r0�#��2ddb�wk����14�J&�JLJbΒ1�(�����h8i��`���n�LɉI 0B�ۚ*�? > P�m=X.����G�ٔ{{�aÏ�]��<���p�a@/&�u���>8��v�J�f�t�'N�S���K����}_}_1��z�uy�n�k��޸�b��D��:������0�+�-`i�{���c���,%^��՝!E-g[79����m��GeA�cL%�;۬p���V���O�o�UL��<�G��߼���%O �c�r����X�wg7muTc�u\e}������{�=�3V��L����Mھ�!��U��*�8�G.�4����b�,fY��S�l���J�vּ�Rg��EsO��49+�(�V�v���=8��r�sv��,�����5N�q*A˷7۔����7a�}�J��#MD�E��{{n2vƾ�����#�]��io.��6���)��[P�t�B��n	���v8@ݛ]M(=/Sq����һ�wf�vw��������mR�VO��ub�����rhb��z�.��U��q�r��1N��䭱L�`�Kf�p͑+8.�7�1�ŕ�sSr qR�s�Q7�LV�^�7��>�%,��(�Jєls���K�s�JSk�k/fT#��!a�d�����S#���m�X�.'��ۮz�WqN��4{y����fO��W��h���Y;�F9��U�O�]o؝f��[��y�M����R�W��.Ai�*�5t�0�5�[M����}�
�#^��-',�I�O]���F༎����[��Z%tg���iY�f��~����Z��Wf���Z��Ίp��C�!&Ls�Vle�PcD���=(ȽG�s�'I����O�!Ol����*q��\5$���'u8�@�n�S�=��8��8�y��7^���}�O�fTjL�	��i���S���w��j� ��*����_˼ƾ�S=�����On�Ln1S��MS���ԝ�}ooFZy��Vׅ�qC�OQ��Բ�WY��u}����="y��k�O9?v�%'n&緎^qU�\ⱏqF%�X��6�O]�O�� ��Q4�{8�6���}��-!�G��=�3�y���Ѵ������FW"̲���N�����[gn��š�]��䆓�Q���:P6^��B:�o,[ٜV.�xD��]��4���l��,Yӌj�>d2MÜ';Q�9��Uw�W�:[P3J|��2GwM���t���ʏU�޶���Y�{��m�]p���}U�����w<Dy��ps��4�7���|�Z���Զ肹"W	�E�9��RS�҅�Ĩq�n��_Y\�oJc������.�T�Ȼn����e�v����� 4��ۈ���S�g�]ҒϷ^��Z�&�r9���gsݷ��/���a:[0ݎ��'BQuɩ��t��I��P��R�����]ѱ[�\e9i�g�J�rۓs�\.u����b���ԻB�+v�)�{�i�A�b�v&����5_a�[q6�y63���*R��͵N끚�V���+c��],�,�A�]A���F7b�1�EqY��
q8m�Nofhw�<�[J�p�॰�FD�f2���N_sY�|#������\c�5�&;h�ו_rp�#o�0�+X�빝�G�)�P2���ۏ�4���TE�8����]��#cAuT��<�Ҭ��.���ޝ�`�f�$S/��2ػ�
�o�$��c.��BE��im�`
�5r����}���^��۬[�\ׁ+n=LTpn�s�6�C����.oc��ĭ�#{�����*�
Z̻�2E�a]��eQ���iɯ�k��<×z��﫳a��y5�u3����q٪�_�Yg�{qw�yx�(�Z���]Bn��-��g�v�?I����������^��V�ײ�и���+0��5l��9vڵ��,q���������'<��T�����〯{�d��Ε��J�I8��/b��#wTW��^�CmTr�{cv�������
yF
i�*Rpʙ��Ү~�N�,�>���-����y��U���d���Ún�6��-8�%Qv���j��/���<ݧɥ��S���2����\���ȗn��຾�'�(Y�Q;�t�U���ǻ7���M�۬��ƛ�Sm��l-��S
lI�)Ew5:�����Sd�l�w8Y�.@��]�Ҹq�*-8���GW�g·�7]����P	��Mnr�=�3@x�V�+�k}�;����5KԲ+����}ZE���t|P��)���nh�{��8+w(t� l��l�F�l3w��%��������Qrz-�{]�ӈ;U�����Z�ym,v�ކ��gD���%��skR��>,G��
B��b�']#s;Rqo m΄ _R�{X��9��w��U}[R�à����I��t>��	�vꨍ��î	7
~��n$������n����r�j�Xa���w9�N�+s. '�
�Xs�iZ6�ڛ�gP�#0V	ۇ���霥�h���%tg��h��V�/'W�>�}�2�#D/G����l��zsP��&�N�zC��3K�/E�3����^�EVp� �Qr:a)=ʌ��W�l�]�l�tU��9��(G)�M�I�J7���y�~�n��(Z�~~צ��Ѫ����\[�@�\�\U���}��\�<j�ݷ��T������v�{�4��E�3�LrL�lT�<�9D�U<�yG:�.qWֺ�E�q}���<��1E��3zJ��I`3/;4�{z���s���:��;�N&�(��A�1Nc{����z�U���oy:�W4�Ƈ%p�m
���mQ��aX:��}�9��8v��C ^��ۣ������j�A��e�<���,nE���5�:N�7���~�e�  ����۸���L��˔�P����{/�o^�,_h쵗 l�g+\�&/�7��Cwn�d��"��EZ���7�
B��U�m$�1�m�PKЎ����(of�cv�1*����;�.q�����U��+�Ժ��iO�R�Ҟ=3�m�D)�W���Þ�T-���E�K�W�mħ�-FlnT?�S���(⻯�P�q��[��*V���t�����W�'��Lb��%�n&)kw��4-���!��X���w�:y5/+h��p�J��	j��z}+��k}�]���Q��Ow�[���CmFo��'�R�SP��m�~2�7�@�������yN���wnn7=SQ�5�rtec����3H�΋��Ӌ`��|w
�|�'5�6�HS��\"���Y���.c>ۈ3KN����:[�ɦ1S��f3�N�쒺3g'��+�����o1�J��
���-�U"^������+�����]���G��~������x^��^z�ǳ�[�"��������Q��gwZ�?x�b5�Yf��%+��RDǔ�H�0S9ڹ������yf�ꍹ|*�r��'Jd/��Mg�j��#i���&�\��[o�t�C�@�P��t���t+�A��:�=L�Z9:�ҧ��W�0�Y�g�upg���9����^�����o�uUc��u3p�k~�����������r�U����q!F}�j�R��>�91Q����I��ȶ�^ӝ��6���l�=EC�s㋴���n���U��	��� B�9�ڢb�n]5��m��o^`J�����Y ���\'��s�Y�}/���DY\�J���=Oq�Ʀ�/��w\b�� A�O-I��-v ���&�[yyՕ�U.��OsR}�ڹ�Y�
��U�Ksn��8<�f�(Vr6%(�|�,��F6�#J��0���S10{m5� ܿ�iu����B\ʅ�&�
Q?ErjoOո�J�u=��Fj�S�*��"35�a���2��P\�[�7 Q��4,��t$a�m�4ܝ�jPb��&^�N�+q��؉�Hs�!O��7���q�^��'@��Y��EwQ�
��}Gtm4Qom�h�d׹I�tn���x�h�|�m��`gs��ɦ����.;liz�ݵ����]٪4
��-f)����Si�c!囋M�f��x�#n��Fpv
Hwu}�L: ���k�J��\�荹7��dH���ՙa)��Em+����m�;��B,����tD��R��sN�'v4���`�,���@W<�岵n
���*dS������jX$&q�A�y���8��}�'�*����N�+���RY}/��jҊ7���sK�n:���\���:�_>�]��Z����]K\�>��mgEa���v�nq�6j��Yq�{pg}�x��r�x1hVa���mЫY�z� ���;��X�?<���_9�q]�P*����[ٞӽ��ǩ�z��M��:�O/Q��=	��y�S�4�z�����wWN�d�:���)Z����Q��|�T<|��w�����\�"���nn��Б�S9�ī���Ug[�UVWѩ�����ۡ%pU�����w����{���P~�j��/������]������b{�j�Q���_��-$:�F�0�l%�����yz����{\]V�[���BZ�+�u�A��OZ��Y�ǩM���kwk#��j���E������\W[�)I�0
��L��2G��a����muLo�^�凵�1�Z�1yw�������ޫ��Z������q�]�t����9F��)?�z���b�\To^\V���\�\8}��ߺm;�����Ъ�P��ܞ�4d��Ԭ��瘗<��^J�E��ڢ�:i��;s��?7M�q�VK�Bh�n�{�.�N\ڸ��FN��{�j9O�]?VhU�LV��8R���� �Ю�g}Sk�2��6Z0�nI��u�ٖ�������o!H5�tK9t��ho,FB��D���~�V�Bwz�7�]��w`�LJLn��]inm.�����G.��L��K6��a�aϱc�U�/�K�i8st�r��ǆ�P��
�tG9sӵ/���,ʵ�oM� *݉D��gj����Ӫ ���q��jNZ���6B�/��ν(CN�����r8����X�}My�8�g�A�����
�����ָm\nO>|�`�Y��g'�\�?vhY��WM�����w�oJʬ�g�C�8�R�dII�^}d^�0rו`�;��q��-)��nL�Ys2�Ʌ|�+j���֧ƥtt/hx���\�/I�u))�s{��v�'Dt]u��4w��\{t�}���S�ջJ=K��V?�Wkz��DbzkT�Q_g<qq�U}��n9�ꉠU�2�k�S�מ�<��V���mM�Խ�Գ�jO+nvc���eovu��*�����my�{S�l��Wj8�~!{iuNߘxd���]{]܎uV���WC�J,����im5�:�TR��5�P���Or
���/k�({�a�Q�;���ϝ��S]�7����ED�Q�O��x(��y�Vɣ]2ҫ+�ƫZ���{��n6�_+��b�]n�zWT����H�-(Z��dV?� �9�4�)����x���nZ<Ff&��mҜw0�n��0�$!=�9B�X�M�▷x�z���}��kTwr����sw��`�q{L��NVJlƥq&��]��w��V�N��]£���41t�l���U[�1JQ�j����ؕ��>�q
^RyG��}��<Ë��\�%���ϰD�.�H��s .�8ޮ�:�&�b����0RN��o�)ۇ]�vڭ����g�,��㒰[.�B �#\��J�����Պn�m���3缱�L��FN�
q#bR�i]�m�m�n�����`7v�V�o�:�uzR����N6Dʬ�R����0`.%P�A���ILu=�k��iޠ��X�qݹ��S*ʨmN�,��Fe��Rm��_r�Rȱk���3�U4�7C�{�6:�C+2�(3B���qG;�+%ZWӔ]��
[����ke�$��S�W4w�kj��
��5{2��E�;IÅ�F�̜�����\�u�Nfos��&�9-;���VV�EDZ��wD)�����	�����X3�k������"��*�=��x�(q�v�Yc�����ut�_J}��-����z���ĨcvZ����ʄ�\rSj�.ܾёak��8��V��^1.ڛӖ}y���j�sԻOp�G@��{�Z�wI0�Z���s)v
�;hԉ�4ʛ��㫡	���m���
�6�p�zEp�������!��u8�i���iVo@k.ʘ4�syR�9�-k��:���)F��'���A�5��a#{~{�:��:�
�S���n���N�}ٝR��Y}��5�*���Q^͇u�n��ȫ]V�F��{���!�|�l=��]��q��ao��Q�N�^+��r4�-�ň���i-��:!� ���Z5j;7���);��-�X9lz�u���]MӰ��Bave\%nq;�:�Z�ˡ���7+��W�mw]pX���"��ֶ�=%�ʻQ�
�P��k���e���ݭ��uޤ�r(Gi�i�/�ۺ���ʱ�&�U1�v�)]��*��J�e��v��(���>��yoA�$c[0�2���D���ˋ�:��r��p;���f�Y�A�%�b��+�w^�!��[Ǜۭ֝�^Bf�5��)�U�/*A�����\�Lp����(�.�.�a���tw��!sS��{�S{%s;�S;ڭ���@��a��dm���-���z�Xrhs��q%XXz�%��]�6jgIZ�cw&k�r��T�r����E����2�X���.����.+�i�_WR�]Jq%[):��}�W�dؘ���!�wGu]N6��N`r�a��cP�S���^#u���(�r��i�y���a@���cv��٫����
�<�9�c��S;W���hB�0�[J�NG����g�d��[��M���On��yS��%�p	�O�A�ڻ���L�:��4F��WZ�W��^�3E�X��t3��n�ɹ.�V�V>�H*��޵��k-AC��r��ۃ��C]9�R��+�3��6!�/��5�Z��_��P먫���8b����ά����Z�3m��Kӹi�Ĭ�pu]v{��8*�޾ݱ�mֺ��m	�9�X��ci��َ^k�  W�*�PV>�����ٚ�Be�3#0L+!(�n��c@d�ˁ͓
3  a2I�CD�0QF��I��%6�FDe�]��(�EF�,1$ن1Q	L�4�1w$k�q�0�d���e%���n���P�I2�ܒCD��(�F$�Rh��؉@�M(,T�H�%	)(�R� ђI3�b
X�V���$�#��s���"����H��&NWJ1!�1D�F�����QF����E��B$T̚('�d,�+����� �"��
$�����|�u���s�A�����¸�x;����M�r��̧����G�j�S�b����z�G|gL�٪�����wm���cnz{x+D�Fk��e���M���uBvbi1�����ڋ���ȕj���<f�n���dm>����E��+!�u�3�`�5�dӵ.G@9�R�w�ޝ�x�]�
��8'�צ��/q*�'����㏝���x��h3�L���**!k;Q&;���t�7s���~�u�c�Cm��ϗo�bߗy�}P{�(����o��~OC��������גS�l�[0.:qM��2�c�9\�^��@��]:�ep	��Ϸ�V�G�}��չ�c�T5�p��& �����i�L���Y�R{Lrߚ蘮I���n�o��:Ք��K���ÿTn5��ܤ'��;�v�V��Sx�=�M�B�޿��܂�������R��lf��OQ��2�:Y����=��U��Jyx��g�������g�*��q
��J�x�+����\R���φN�Y�r��T����OY�ϳ� ����':U\Y�67|k�iu�a*vxb���.�kr�S�\�O��͏��
�r�-`a���\��O���B�K׼�Vf������t���)��\"N�wZ�;������;ht��5R��|��mcj����"�i|��v�����r��qz�����qB�o�\�`9������+�)[t�^�\�S��ڜ�J���\w+�1N��f��ݶk{"0o��[������/AO�i�vҊ'�ޚ��k�N�.lk���<S�c%�8����qX�.����k!+�os�lu����yfb��^h����5�47Sz=]��U,�q��rkݸ
�;Yu˪k��)�)i��`CWt��JN���"~P�+�4������*���gZ�P�U{��9@���Λ{��I��_���[�˔kې��Zy�W�R�c)w�|�w1o��\u-�ܽ�3�����)��k>�_<�<�;�E/iX��y[������+���	�b�=<&�������|-���"���$}<�Z.l]2��e��Ւ�����{���kfd������VݍI��m��ek�g�=>b�'�6�U�o҇ǂ��b����ݕG���|��9�]�XO����"���n��jjF�iYZ�����nG��ܸ����LjFuڻν�~<���$��p�@ƙ[�[{��z�I=�x�JSTqQ��\.���7�9���MOv(r��b�U��u�G�Ąяw�Ի~c�i������*��&�{�y���i�=Kݯh��4���vʻ�Yqێ]Ҵ�������Z���c��y5zJ��x���Z�b�T��u�5"���,��b,�����t�vX��ul��}�(�oiMv\j���A(Y�Pbw�~�� um�}G�6+^��*��g�L�mybkB�nn#��|�B���X��ö�����-V��@�<���>�����������7q��W�J�u�tXao�3KUO;��J�8ק�|�f��>�� ��y1N�ؚ3eı$[7;��o2��Xy��9f�?���2��oݏ�5~N�<=5��=~���L�J`��T9f*9��<4
˾��w(tU����!:�_=knJBj�On��v�wV�4c5j�E�n��ײ�5!*��  �ztplʚ,��؎_9[d]�U�F'(V��W]���\������h�ά^Y�x���w�^Q�֊<���6N��{(��q�����u+��лC��A�".^h��ྒྷ�/=Xf>�{��6����=
����g�K��3K��Onoh�_5ӘV���c�!v��pv��w\L>��������ܳ��Z������voѫA��'i���
*1⨆�'���m��gqaD%Ko1¾��C��YZ�W�����*7������;��i�}�5��8:�_`��ûjE�WQs�Q��c����l�tN[�ą��n�;�3ȥ"y��������f���k8���TB��ꝎvgW�Ѓ��$������S�o���7ko��:�aJ�+0u��C�~�0�(�F_L�ٲ{��#�S�)hn�>}��d�w���}V���H��쩸Y��{Wi�ТT=���uW;�U��)�v᷵
k��gT�.�ٟ/�fd�b���.&q�:8�9�g���0�Y�{��%}��˻�^f�u�v����ddf��L_hƮs6JRWZ������76�m���w�=t����+x��/�7��2��S�ʇqSj<��].�T���`-�t'g_0 ����ܔ�/z��vu.�<��5��z�l��/<S�N����{�\M�'b9�{6R��~�]5����ɷ��ԅ��y�(�]=z��1��9r��0�}�9i��/�t����uf��,_5���ܼ�S��y�\8jb���ϛ������s���4(� ��t^{����ګⶒ��TBvf)K1Q�v�g�Ԟ���#���ug$�^�~��3S���+��[.d�&A��ɋ�V�{{Q�����I��\���EM<��<sZ�zB�����T�sJ��N�|�Bw��_����vtdf�Ev�篝�]��Q����j�K`�0�w�/�b�Ӿu� ;��L��j��Uy9Q�����N��`;r�_5Rq���7���=P�2i�Q�nW�GeDWQs�<a�Zo�Чch�h���r�B�����Ԋ�e��[4Q��L<LV6�đ�ԟV�xQw:�j=��>�Ꮤ�],-<x�����E�u7�ܜ��<���&rfd-KՌ�K�4���ט�;���[�9t���Y��eH^�&��m̓
�gW5Hn�<·
��B�~��pꝾ�]�s�c��[��Ϩ"��*�e��g������2{������4���i=�w��vl>��k
Dr�f{6`�n��\c\�pd=���h��,�Zoڛˇ�kyЧ�:�͎lJ��SC��nl))��*����Pb_�H��t�|{X�#K��C�d݃�WA ʅ|���r�i��aj`��;�
���};h����p�Cbx�E��LȔ�{=RTl��{��L+�]G]*-�7jS��^ ���W�J�q���0��NJ���\}�2b�%6�Xa,�y�2�@.���OW��&LW�{׋���TV��O8,q��JQ���h��;L�1���<o������1<�X}��;�����u|�B��A�׳������Y�j���
���Py_B�bV��'�p�0�#�Ҹ	�ޣ=V
��w>���2��B�h����{����_S��ݽ\0
AU��6��9�[6X]e�L/���w<{�.�`Ս����!�oO�<gC+2���aQ-���5q[�㤔���N�%1˳��fv���-ǋq�*��DZo{{�a=�W:<��������ʌf���@�p�]�i<�s��1՞��"b�3zm���Am<3��jɎ�)�.ˊ�"�48+������D2�*����v��df�W�����T��l`�%�V/��n)<��䪏��;P��B��֏������
K�s'�c��;�%5�i��ҟژ9�q���N(�_u�7&^���1��Z�f�I��*�[�7��ƫ��ʌQ��A��D������o���q�D��O���gT��^;�wg}oj�b��e��ꉊV���6���U�*nz�޷�J4�|�U����W7Ԫ�:�qʣJ�M�%!���2��"y�Qʽ}y��v��`Ġ�٨1Z�E�U���BU��ӣ�C�6��/�nH�zw�U��9�>7Я�ur�c�9�l�M��`���UNܽ)u�Q�v^({��F�q���ZT2�h��ʃ�n�"r��ǵ��|Z��2�U���m�Ȯ�%l��;y��҉OL$e��J^��hVc|{����3��PDDe
���i���5�Vee�m��h�[za��}�<0 ��Sح�C4m��;�7��'X6bK���Δ�B�7y��3^��] ���k6{��������k��-�4ʧ�[���0@=�$u����F�ě��]����]?Vꢟu�7��8�ǋL񛀧5	ta�ԋ��=�[аC[�5mĘZ�"���'=��N�jZqED��Y�kuFr������ữ�F%�\Oj'A����ޅszb�0&i�q��yOr�b�N!�l�qڝ�Ҷ`t.͂���]�n>b���;��b�=�P	�cml����N��|D��g�����f���6_��݈�U���v9�1���t���N;��%�q\(n���#2B�1��� �{�}��j5�3�(;-����nT����c�X�)C�]}��84��z�R;:���������>�U3���4��U�:}܉�����+pg�>K7�V�r�e����}+[�q��u����1jmi�vl��,��Oc���)��nL�W�HPV�<��[��2��lб�坶��ʎ��<VgΣ�\��V�zjl�k���B��p�-+E��K�W��e����C��F��tv�Z��-��#�ٮ�{�s*g������� ١��qv��EERw�w#;b.=��0q�m؉�w+��OԹc�w�_7k_X++0q��l��|�et��i�T	���in��ѥ*���&�nD;{JU�ȇ���[x�1:n�L��.&��-�>{es�冾������6�zk���w*�L���n�R��XUPʅ�q)E�w57�b�*�+��Cݑ���-Y�]ۅt�#�nSV͆�%P��&��R��Mf�5sҒ�{�՜�W5��d)��B�9��r��r��FKr͈�a>�]t�
��Cy�mE��q��:��9����Qn�LRB��[saӸ����=�^��0$M������Z��u��.�͗���,�A�K{-iC��Vn��9��8��?�X2�N'�
����.�Y���0�)z/)��ߴ
��#@��PF�h�w2�ʹ)mm;��˭�ո����k�3 5��/��X���l׃��=���%�kF�(�KW$��i� Δ��9���)��[�*�V^+�����w}5 �9;����t� ���r�{Sm�:��������7NM�s�c�Jm�4�s��Z�lw�_wY@r5���J*�\}����Ŏk^v�Z)�o'�
U����c�\��n��)jFj�������g�Ev�篝��U7}�\��١�.X��}�����k�nq�G��;U츶��|�~+��j��7v�l�)cOz� ��5N(�z���t)'0WZ���.s���i�jr��8�3����T�)�~���=���c��[��5C�T�]����5�!��e N�8����y��~��A����T5�P�i��jя-�ї/��M�C���t�eT{b���u��&|���s�{
�����ǲ�9����I�{9kɧR[��C��c�*J69O��������S=�L��s�T;���yEq�bk��n_���(�u����������\�Xe��n(�M�
��sq�����\�4���*��s��]4s����|}5���9E���@l�ޗ@>Ȫ��.��G�����~��*ޟqWXEM�2����]);��w�u��da;���&��F�Ɠ|%>x�9��췚�=M@]3�zƍ"��w�حրv�Dd���ܽ"r��� �)qDwJ�����R���x�Z);1���y{wV�+\�x�Ʒ��5x�L�d@B*h�,�+M1��c�����s35���Z�LZ���<�y5gkb��!��X�q��k���bZ۵[{(��^�*ۤ��N���Ya�ӷ�����mns��j�g3{Ξ��7���p*��^��/�mjd*w���۩���߲�$y ���^��{l.����V���ά�Cz���6�;�QEud���4���sG+�������%��n�-@�b�t�*�0a����`պ�Qf\�,e̗ՠ�v���3#�¯�Z����g�f���|�,��>�������J�9g�:e� ��]���y)TL���L�&
�FrS������L��]�f���q޶}��Az��]ȍ[ ��s�Nڃ��V�6n�����
���vC)����gm��޷G�Aka�~��jD�i�72�Q�Wp��=fD�`d�e�1=�\��ޔ���Ù��OP��гw����
�?G�)e�!,�4��}��X�5�o@�ﳢ,�,��vMI�㑮&E�/�)uJ�p�Ҟ���%r��0��Gn�k9�	{ح-�/���b��w�Ⱦ��R�7��/m@�%ud��9��Z�
g��qn*yZq��w��D���;.us�k�;ǫ��S�;�h�[�z%���p1zy���$�l���s)2��*���Pp���K���ZjGyKT�ځ�1�T��CaJ*z�B��ϲ"h}���8�b5ܔV[u�N�$鏳�T+�����Q�.���9��u����p.���W�uT�u`��W8e�g�F;U*"8n��#Ej:9�А��#�Gk��8�Yې��k�7�����m�;ZN�g�̜�t̍Mq���v���!�5׋2��d���D�U��-i�{���+f��n�1+�q8���I��ô����K�k<;������t���rt��,[���ha��<��#�;�t�`��1�V,��R�h�0jҠ�
�ZV/{A�:�ije�v��s��q�0�"v��J�H/&��R���mNל��䭺����m��a��?�T�]���
ׅzn�j�1���9c�����\4E�M-��������8�c]�X ��ܱ�"W��b��C;i��zÇ\�a��O��jK��k�����M�
�M��{L�=.M��E�R�6GP8�_TQ.vlu�W����Y��"�j�x���VgJQ��΋l&)��S`����T�u��`U���4*�
3-�vؼބ�&��uI ��_&�z���v'O�ے ��a��;.�$W^���;d[��$��+7Fn@�˾��@�X�D�o�����(�ۉ��srh��λ#\#Uf�*�(�bfwfљ�������߿��ޒ&/nl&����+��L��@c%23��F��c܍�.rKK��c��n\��ݺ�����a��c9uF@F�r���x�;μ�E S)1<[�J��E��;��"�c���J��.X���#`�Qx�E��.+���ܡ1�*0h�r��x�1�lEx���](���b6H�E�μ���vK�l�b��	��h�ҊSs�]�W+���,X�F6H�v�^6�9n�$�j�2c	(�J�E�c����-�&����wI:�Fw�y��HhX]���!��U�
 V,D�䇚�O�um�!�ʐ�5�ػb�/ni�9ؽ�����y
�e�o&K"�b�erޜ�M_i����,��g�L�(uwV���cl�o�i��[�y����͘:���K���sw8C�ս�ğh�L�a�峙�ς���]w����.r7�;��dnY�]�)�:����1��Z6:�/�ya�)�c�*�����=8KGv�]\</���t��~���/g����7Y�̹=�=~b����}��鸮�>��z_�tvv��R}V͠��,�@�_t��u���5�*�}X ��6����x��5V�ܢE��M}��~�`� zS����à�^��ʔ�Ê��Y��ޠ<�'�P��ר��>OM]xnnV�q;�5��N���BYs/�]�@��3>e�B�s��EO���{ʛ7��^��O�Ț��6�E�����3T�9��3 �2���Zn7�;,��ǅ����j�*n=άu����1qށ=���Eq��;1���i�|l��,���qC4���H뎦�ڶ@�^������-�2�,��H��Mqּr:�M�P��Xe�,�9�����ڇy��7�@�}R<6�]�Qi���z�W��
�8!i� :�Yu���	X��tv�E)R��	KҪ1�D1Y�'�;��9:"��+T.4����Oo�	����gmk�8zdY�Ev���Դ���<�me�Åt��e�^�p���oF*�[Ƙc6iĺ<NB�� F�ں�X7}4�Q5�rf75mr�=���Æyh�/=���V�*s�,f*�vNz{�&o�X�wY��Y�~����>����_{0���+����T�ymV>�)���
Ϫ�	��\;�&S�Y�O�Y5o|��gr�jp��]�|�/�#��q�V�6�9�e_��"���j�}3@�481U�t�W{�����"=���y2�}��<e���ǫ���_�ǹ��<|)��Q�TX~�����l�DUH��gQ��)�[,*��������蔏o�a����uX��)�:u�չ�i
Y!Yp�̇齙PL�c%z�%��ͨj�o�b��R7��[|��Ӹ
���
�zb��p��N������g�a�#�.6d�r(�ʗ�� 4s;�ƢuC��K;�s3�U�d�����O�~� ;�=�E[�rE��Cŋ:%x�Ee1N{N�~9����"h�����{J�@���>B�/*�,w����^��P}~�$W�@l��>��Y�G�H�ʥ�V������r��({d���{C+�B��ʽ70ߤ{�K���^��F�����O����F�6����_u�F
N�"Կ��R���w�Z��ԫ,���d	�H�՞���^aG�ڮ�����g%����m�}�=�ؗ�u@����\gn�N]lV�EikYX��s!��\�ecȠY�+M�Q�(����O\d�t����3[Lz�M�}���#��p̳�~ʀ-=����mUj��\�"|��2���dOT>���0�6������� g�^��UE�o��z�c�J��4�F{�ܶ}���wM`�(��/�E��j�L5�ZoK���`	T�
�V�̙>[5	��i-����Nya��خ>��P�����;�V���7��d�B���,��7�\�Uf�\{���<W��󀼕4�c>��=�G��Et{�_���w��ւ�*��ɭ/�D+�=ٞ��W�w�Xv|��=��Sp���d/\	�u���Y�=�^<����\i�[%��V>8��Ԃ�eGI���A�OYc�3���2�y�!���{�?:�=�iQ�\nG��|a(�Iŵ7�륹q�4WOJ� ;�������~��@�S=�,/g;���%O��~�q�z�;�m��:_��tvj�J-⫿XT}Qꎿ�z��8J��G@��
Ex�q�����t��/�N�����[җFí7������~ܖZ�2���`{�A�-�
�����j/Þk���Jv�՛��1�7�aO�^� ��=���q�5Y�
��A�=�R�����J��X��`�t)�X{ �1+<�r�ͬ}�,���#�9;�ɆC[5���2���1�&��^�r]�V:�Zx�[��Eq[�a��؊8�v�=��+H�ޒ���l�S��U�/"4��ىL�}S#*%ב�C��zƪ���6�q�~�6_�[�N�gޙ�%�zGy�*"�S�����������b;cV�J�����8Ό=+N���W_���c��zd�΀ײ�*"�פ�O#�]M*�d�.��P#ݧ����F�IVѿ���ݟ@�2���b�zi�s���S�8�̯!y[��zO�:=q.xJ�}}��5��rˤ�e�;�^�W��.���+��E*�}����y��.3�e�w���O����}�e^vjQ��W��Uc�ssj��m{���mC�L3�T�kY���b�������φ�~�V�g��P���7+�dvK�ϯ���V����c�>nk��X�=�p�����3�{�n*���G�����	Cnv�ɻY,�㗾�7��J�bO�+��´޹�����\�^׷�!����<�ۏv���k����H�#V�3#��g��2�kJdΣ�����{{i��^�^��\;޺CT��>"�����j�WEu�.��=��N~����9�p�r0�C �뉾�sس���[;�@[�0��1GP����~���@i��oO�,G�]YB��״��s�U�x�0���e��e��-&^㼱��j@,�4.���Kx �Z��;x�/1�-5�r};����a�WL^L�73��GT�:����=�ߙOx�x�1�7&}w��i��^nUW�+�ܿ@��<*���N�&����\;��o&X^9�*�F�8��y^�]��O<���l�����n�[�(���DSXg���1M�
��'8�纖}������t�ǐ�S�kn&�y�G!���{���ߪ�*�e@���/UHɢ2r�z]P��\�y`4���)����ա�~��dw�Rg#}#M_��?�Ic��A�uQ��҇;����ƨ���ET���e���^9���/����wkō>�E�x�P/�pB�{�_\X������9�2Юb��(>��b_O��%���X�=�å�[8^W�W���-�IJ�]�7(O��-̉�f�\D����!{g���11O�h�~;�aᯗ��>[6�a>�g�.�ۋ�R��^�#��x�� �<�	��원-H�}pj�1ٹD;�읍/O��`�O��V�+�\��}Bcj=�\ٴ�@y�p{�<�y׉y�5���׆��ho7DO��r:��?���V���,�z����ʶ�ƙ��sX5Q����˹�A�W�\�}�_�wv�Y���&u0dN�(VV�J�S�:����
��M�6�V^����)��jث��ɪ)���'R��֭�T'��ʶچ�.�8�Q.K@�j�u��}[D��2E:��L����iAT+��k�����S���C�[�?e���_�x�`ި��3D~��U~��g�4s
�FN��q�X3��Ϻ�q�z�^@ϡ������Zj���8`<�b(���E���]�ooԶ@���ʓ�;P��/6kN�{e��U��π�W���@�j���O{��g����kEh�/t�Gd�YUemC����o\����xm�� fxG4B�>�R]r�
y�Q�,ٯCu�\y��<�R�e���hҦCj��2g}7��>��=��O�wGL��R����c�Ɨ��Z)����p]``���b�����(4r��wTwy�X�ǵ�1������qw�9��R>��)ի��{e���%�-��w�����Z
�J������~��R􊋟ߏ��L���ΰ;���tk�N�P��m�=h�c�ћމ��^�W۽��ϡO��U#	����u��;�_�y��=�{}@j�0C�"#i�����o>���G�\*=zd7:O@{�R0WҽKA-fF�5Qu�X���H��<�8z��T����n�?$���Ӛѣ��T+�E
W��tzl��hiZ�U.�;`�n�Z6+�C)յ��Yu��p�8��ge�ޖ�}�w8��ѹ}{���iګ(* ��,�Rԥ�/xT)@z��^�m��eX�m�>��U8�1<����__��"������sq� 'ӑFFT��a���&�ׯ��B���[�[��w6���G9�T}s����@��dT[�rE�y��b��^=7$K=�7��鮓뜼���~�+�e�a{�H�_����^�
�~�����"�Pȉ�_�yfs���G���׽��#4��:�g����+�5W�&1?P����=A� �S�.�Y~�ޅY�*�{����!?}Y��i�c��\�����m=��)�X��Q�ŧ�����WJ�|�[�s��=v�'� ����R�쉮��g�Y��׸�zx��`	��x_����FjKє%蚎���VZ���eq��uyi��!��ŵ����Ou�ǭ�\ 70O���3��RAk���A�f<��s��#�U�<o�v�п{Eh�^ڞ=�%�����[�]-~��/�����#���Nox��S�{������x���q�J���{|�C�#�ߔ�*e�y{;S�?UW���̟$oѳ>�����	���~�n��=G�sO{��;#�l�x�d�M.=�>�fiW��g=�90NE�����9���Nj#l�;m��i���x�P��o�����i�'-���ԨW���S5{�C.�����.4g8�a�s���6U1���٘k�h+v�� ̝q�/+Z�<�blb���m`�x����oc߹�&�,h��Y��:q|��h7窱	����y3��dϑy�!��S~�ѽ�^G�.}�^����ED�A
���w��/0��h�e��pSȁ_}~�����xX��X:#}�=3�{؍�*{j+�;{|����\�1�ޜ��W��9��1p2)��J�u����mC>�ep�8]�L��z7�۾����?
�K{�Ç���ҫ,��	�A��=�ȣ"�"[�SS�б�U�'}ފ}q��)�l�u�z�^��G�!�F�'EE�����.���0y��defnۨ��'\���Z|�џe�<���Q}��u��#�;ģ��z�>�7X/�2�^v+�߾�k��*�z��L4/�U��R�Ό��Zv�Gz�z�]u���9^��O�`+~ˉ�syC�ʽ�;�QKk��
��ӑ/ǲ}��#k	��j����|;�KP��K�Y�>��LŬA֚y���p�M9xe� ��5bO��5P�~������t�O���4Wʄ�*���*��O���*Z�X�=� >��P�/(
�;5(����j�{N�L>�6����������}�� )����75�'yK�ԥv��x�k�-t�ܑѝ�W7
�-��P�dx��/�.pR���c���	�b:5ҔŞ��O��lGuv(v��%Xz��1����E�us�X�V�6݋����4,�_Ӗ�q���Cy�9�U;�L���w�%�tB�"��dS����,�2�]{�r��s�t׽TǱ�5b��IG=2Bñ;,e�z�;>� �'/}�7�7O����ٟG�Q�����S��ݻqW�m�6��N�H(be��yz�5��%K� ���L���7�F�o�j�J�������*&���x���MO���{�7Ȏ>v}.F�υٜ,w�3�:���G���[U�5��WC� �:����ڮ}�.�,��N�K*Q�g��g>�N�+"�=��1]1FL�7�>	�T�;���z#�l��𻵶)��rq�;�S
��1���Af�4���8��j,	��ø�2��ɖ��o�E��{[��ێcc��'�#�x���[.Z��9E��~�)�����Q�'�n�s;1n�c�
�x�{Z�^����mNG<�w�$r5��\r7��ߪ�~�(��+��ݏ;�g��[�{�>��&��Ȥk
�������3�z���a��������U�������7���<���c�>�����Y���޾����
!��;��Ç��������~��soͺY��"4���6�==Fi�%�]��l>� +G�Zq�]�h,,4^PV�&5%�g˞o��Ml�
��Xݣ:�7�3K��u\��
�q�{O ���h2RCD�ɜ1(b���Vy#��7�;��B��<���_�T;f'���1<g�XLLS���9�X�B���j����To�L'�:�u`�J���q�_�WO����\�������6dS��7���`�xG�� ������x�z����0zǣ˪�r�@ydX W�X��耋��{o��yl�9��2�Nˮ˽�G{T8�*��Ei}Fa�G:�6���(�5U��=�>�Iuw5��Ϧ��7���;�����8���ymxMl��f��z�]�;]U>���z*x��8=�3�6}�%�����=�_o~�����ه}^��xWFN�Ӭ���_�<29V���>�7���c���1]Y�woR;	�1�8�9q�ڏe�{��p�����0%M2^�����c�{��ڮ�>�����}���P�v�О�=>��VET<5[P���{�� k�#�=�=U�g�۾��_>*ob��y��U��Z�N��{�C#vK:}(aS!�Q�����r�]3��?{@�6M�*iv�Gѓ:6߽~ӑ���}��ױ�
ȏ*�}@S��dUX
>��mV�*-�bТ�2����8�a� ;�EY�j�C���1���T�"X�e.�,�h���zF�s�#����k��=îp�V=��z\4`�qꖶ<פ#:�K�/��MW#��i��w��Z�mK[+)w���u��В��|�@�}���&���X+� �=N�7�M�|�^1xY�p6���H��X�}v���ַMk�Ď�[��#,�JX��]�u'���彍As-����!���s�u�[�J�{�k�ݮL�^�Һ�����B����Q�t�r��;���+��ŵ�^�:3��D]�R7O'Q���o5���5L(��ƌݐ5�v�|�v��Ex+1��Rv�!�e��M�_e�O���S�h"ݒ{H��Hq��HX��V
�2�A������ņ�
�Γ$��'�G2݆�s����;-�$'��iΝ��h
��f�s���y5[۸�uS�*�j���Bu�k���C�DKڛi�>a��"�:�nFPs��I��*���:���_eL�Ś�HL�}��\�N:��iu���������+���,�F阠g,�u�7�U2�B�4��q�g2�a�K��"�56
M�+��I'Z��(�/7�R]������Az*���@�c�i�Qv�p��%��<�+�=Smiy�z��2� �*k�cb��ܲ�gf�b_�����2�Z�s{R��#���sw��Z�H�#x�Y)��z�;�qf�}��|�n�!���K�N�,c�q��ܩD�m��t�֘ǂ�������Vc��.��M]���ʷ
���)r�H����e�M�B�G07��[xޜ��ǥiʄ@��2TU��v�o"�=�ή�9�u����D=���S��sR�r��&�+2��ĝ�k\9�I�O�w�[֜*r�g�/�EG���gd���&��P�}�_c��3mk�4;�?N9I�r"�s}[��2��_٦��o�R��upCͤ�ȁ�쭷-���ܲ���9J�0�-����A�ye��P�|�jĩ�݋U�wyd\(M��hS�����%Ð��7g��aC3ӎX�����9��܂�u��Z�#6���-�vk5�uð�I�ε��6��U�R�k(���I�_>��\'�5�$GMeI�pSŴ�t��+g>	m�h��� �-�����
�?�0V���M�о�gMHP�eb�_�w���$��I�q�E�:�����Cp|6�u%ǹ+��(�r������9Z���"�I�!2gL�\���.�\Ozwt��;��1.p��Ok���v���/B�1]�F�TܧVnͫ:�ofgv+�o��"q��WA]�.�&ԫ�Q��
��t\O�`��u^��&�c��ו������㖽/<"���>�t뤜W!p�Y�m4��-��p��7�*�tW1�Z�q���,Ao�\��d��uu$�;v,˛y݋�t!�d�DDC;�	��Q&��؍6d��ʂ���7�Й�y��F�ݮ\2�y瑒��F1(T��t�.s ͗�s��(�XB��F����b�o�Y��&�V-�v*"����u���;��[�/��w\���A��[κ-�nh��5�7+�TF��ۛ&ƹ�CxܮnS����KƊH��W(�7MwuwuOY
KŮlI��d1&׍rK��7��n+�+��H����snj抍d37��-s]������w������ιۃ.�l(�|�5k�˫�u-,�o(��ם���ؙs V�5Tmm�CH��w8s+�.]&Mw�%)��2Ӝ�2���y�_�G��T=�q��TYW��h��c�@\�,�-��S����U�MO�s�|/&[>Ϲ�c���5ǩqȇ��u�����Ģ��sw�o�J܊ƌ?D/
vo�K�dUHʙl�QjW�����W�({}��d��N���mo����}�o!�u�9��Q�=���*W�a�%��ن�]w2�z���^E�^�����a�ZTN{x��@�F���~�R7�z�ni��72}9da}^��KGu�c�k��X�����_9ќ}��=~V��#�{�����d
��2EG���`@���!��O�#�&r�\��w�*h�����Gt�ļ5�Lz�O��ȇ3�>����W�`W��$\���ۦ�Q�N0��ºY�?,�}s�2*5�xv�WʅC�>���o�c�w蓐=Q�]�|[Y�����gr���]]Ox�D��{sr�<>'�΃5Ly%�]G�����TC�㨼������WrY/ߠn\K�M*7���}5����0�3k�o���3Q������=&x��1ߞ�¦�/e���fhb��<����l�y.㝂VT���F������0�:�/��P���8Xq��I$5Uߗ^�V��8�%
Wc�P��_��tt�%��Sȅ"��;��}P:��N��}N�C�;SgW7�KfdrR	��^Ԝt�"�l��rwѾ���9��k�z$�ˏUv���xs�0�f�i�/ǧi��SZ#�[��x��B2 zZ�.<����7�ݺ����/mO���ge�?-f�Bk�^����o%��:����e��7�k�I����=�G��EtG�!�;�֝K�<���?0Y޶��_m� !�<_�2g\�ꐜ��d{ls�@�>~����5�+��[e1�uCŜK�H�����U`Y�ɝf�ɟ"�:d7�}�c��ב�e{�l,��F���邆*�ttjX���:��aW��U3r�s�V�� U�S8K˩�`��^���s�9��V����J�w�=μ:�U �6B~��9���&� O��QjW����h�`�����u[}�%^�wz
WF�'û}@`����d)�,�7+��`{�(Ⱥ�n�9�K����ɢk��N���K��\}{£�ґQ�U<���	�^����.O�1-�pǜI�_�C�ɑ����Q���M�3�xo����E�T;�]~��L���F�~�!�n�� E=�i�r[�x��Dުq���nE˶��M[B7Q'� �Z�C�ɴ�'�ͩ���ʏb��y�#|���(W��[�LMkK��Ѣ��e��t���8MN0�M��P��0V���o9;dV��Q�_.ܽ���.ﻭ&y#6$�T��B��G��,K�U��9�ta��;��5��C��:�u1C���n"}���u
%�Va����G�{̛�aS�$��DO���6������7�û��
h�*9z��L{�9��;Y�w��
������=w W�ߍ���P�Ț�����a秤�x}N#��D߼�5㽻������|���9���	�R�~�a�ԣW�������ܘ}��>�<;�ǎ�;ڏX{�(RL�Tr4���2��}^��ު��g�U~�����ϖ/��nl��yD�׶�Z�{�/B�:8-�����^��fs����{���Q]�GC~�Oq�Ѿ��2���v��O�o�}He�Mi�,N�����'p&�{=03�n��s�-ۊ;_��΢���ޝ���� &tǣ����,��c*2kK�;㬁����{r#��'�m߼j�=Y@z�wG{6��uW�QλѾom3��W��zJ��Y�WL\dγy3��GT�;���F]�2�yY��t{t[P���g���G�=����!�~��R#]sr�s�Q`Mw���zM�S�x�	�}u�O��҂൷N}jQ��1�u�I�V��P���Nˊn�����������l�2�e�\-t��ve�<; ˗�=��q?^T����n�˗҄�]4l�#�U��-.���Kw�.g^�fNۮ�̛%b\@����R�����N-�u�O*
zCG��Q���~��x�g���Z�+Pg���E��(�Q�\�
��Ԭ/��﫭dI�y���4o�2���a�Β9��+�F�_��_��!NQe�i�&�Y�U�.�g�Q0���誑�e��r�|�dl��"��;��[f2;�ߎ��~�P�݋^G�j,>��䜅�Ǿs�n6bP}�R0���+�3g�U�png�PO�H�7�=3������E���#y�%1>�]����p�!��3lĠ�>��bb�W�����,z�������s�u՚��V7'ه�ӕ�V?{�ˌ���_Ҩ57�B�NE`���մn4��Bv�R.�/�M@Ѭ�>�#H\{��������~� ���d
�C�n|j�1��D9ܲw����ew�k�>�N2��XT�_.�͛O���uZ=��y�z\�L�-7�)}r=�X�ɝ3����aD���=���'Y�����&�KYwp��Q���u�z�G�ʛ3~��Ǌ�y//��n�?~2}�W������ܭ��;�5����\x^�א1���=?d�3�]2dR$�ߜx�}�^�r?�YƲ��%�pPb���������4�\�T�/_TȬ��q�Ѥ/LĮ�Y<���Ej��7�إ�Sq��h�n����R��9ZL��^��+჻���r�ڹ��>v'�kI�x\��[Ґ�>�6ViJ���t���.h#p'�ߪJ:va�ϴ��f��k�7�L	�m[ M�.�oSU���ܽ�h���9���Z��i��:���ڇq��7�@�^���0J[VWn��U(!��n��9�����W\4{�E!q�jY숟V�*d1{�����Yt��3��FnU�.�����tφ�?_��o�?��q��{���9IG��H)��\-G��DQV��`w�n��辅��9eǯ&}��t�s���8��~��߽��.iTf���*f�����e��JUB�����U�D�쪰&*ye�Œ�����OSGFC�J�~�SE��l�9�f�ݧ���8���wl���O������Kd�R�]f�
�:<;���OOZ�a�z)v��c�]ѱ��~������9�p�L���fT�U#DJ�, 4}y0��ܞ�/չ�#�~�6=
��zr�/>����둱�j=F\��$�o�2:��}~���y=���)�v�f҉����@��5��9�����{Հ��dT[�rE���`h+�X��W���g )�%��^ʂ�<��0�r*��]N� ��m�����Ѱ<CP�pZ���bG)nrxf��;���D���B�6��j9���ݹ�.A[��r�O�nT�:P��^<��0�4�a+y�e��pOwqSөƗZ�������Q�Յw�mG o�a�Oj�9��Iߧ�@;�ʀ�_��H.����c�4���Ҕ(�ޗ��g۔C��V��;���*��^����C�s�s�<�V�o�A!zϬ7.g����!� �������"�4��_=Lx������;�X�2K���*��]�d�+���_k�W�������ۀ)u�To���OT{�2�L<����O5L޸��^\=�d�ZG�8�ww�=uE{��z�꡴m~cU����?�Gq�y�M���X���v_m�k�@y%ϕh]*�����oݻt/��Z��#�&tf���l���1���v����7ޛ2{�˫�oO��7}y��ߏ�����⸫�v��'�#��U$Y�߹���Ьth_���Le}�Z^�c�������[W���;���y����j)�/E���������vO�ȟmh*f�˞�b�gY�ɟ"�Cwƽ��y��V�7g��������^�>�j������fo�S7.q�34EO"��{&X^ȍ~�῞��G)��Y�}�(@�f�s;�s��N�Z.��BU�%��0H�^�����3m��|^��/i���V�0�V����W��O�N�fd�Zq���8R=QȺZ}��m��}-�S�g�:��tް�S�ꕶp�ї��UM�Pnǣ�%�����t��u�?Q�͹�숚��1M���u���f���X3��c�\}w\<R8��n�������+>UA�i���J�9d\���n��UA�;+.[\���z>�EVF�y��:��r=��w�pt_�܋��Qy�@l��������3'}����u��L��T���i��~6��j+�Ģ�ޑ��{,����N�O0۶��<�@^� {��K�ىA�VYN{�FA��;���ޮ��]na��zgz���;����˛�Zq�ܜ�#>�.��3*H���eǻ#k	�jv��q�XųRX���v�3a��sSj�-{��ˡ;7��]��~7�])쉫�{�Y�竤�z}Yz�W�����6�w�t3�� �1�����e�H�T3�>���y�(�ϫ�r����	���Nv:��=f�g�ta7�eɟmG�US��]�##�x$}��5Fϐ%�� ���;�R���n{e�l>A�絡�d�l�l���Uz�������ޟ#~�ۊ����:T}^ȃ#Du�b����#P=3YT�QQ��O�ej�j1e�寞A����"MG�J>�{}Юou�z8�ӧ���U���D�iκ9�O���/$�.㫘���-�5l���[����(��K�Q>��ZN�8m�},#���b�1�z���ǕK���8ԇ>i!�q�-"{A��}�����J��>vP�ɭ.��b��#==XK�@���g��ӿy�]�jr�R����.��p�g(�^��k��c�a>"�r��3�c~ɝ�r����`|MP:4S�sO�Tq�g
��i�|��u��hw{*Q���g"}:�Y߱]1��=3��cٍ�=�{�����C�|����#�s���=��C��
��vmI����+�P���)7�=��i�n��ӹ�e%�U�/}�״�Ѿ���/Ã�T�)�,�|�DS�������8~���xwj���������O��w.D\�9��,�s���$n5:-�O�ܯW������gy ̙�4��<sY��e�)� �>���>�Qr��5��¨�����m�_T�]����u�����F��H�8�����OI𕊗j�Ĉ��[� G��,uF΄�u�
�'�wCȕs�����gg�G~�D'U6�P���W�{�\LS��%���X��J�ȺV3s^�r����8٦}��+�����w��A�?�P�K��(";����T���y{�k��l� DE��;7TdZ�ybr޹Z;��Po6{��޾��|��T�Գ�%{�!�{\��8���e��FOX��.غy�4gJ��{�io���w6��@������3�<2��Q����o��ܸ`"up��tJ�V(�;ށ0����i��Y���dX W�e����H���U�;�����=���I�L3��2ҶK�9�3��JMF��Q�/M|�L5ީ����"\�py@Ty�zK�Y�9>��b�G�W��3��&���ܭ���f�X�3������_]צ��=�U1�^�ywy7�rnj�*�~�R;�G���z�Cǲ'���;�����޹��m0'���^@��<���i���Y�:��}�hm{�f�o���}$���/+�X�͚Ӭ����<�n�^�Q.���^3���9-��S��ɱ!���Z-{Mw��:����{��'�4�ޘ@՘�1-h7Upo=��>�Τhێ�`TZu�=[�|���<�R�����hҧ(��7D�A���_����ў�3�o����e�������~=��e��^�y��qP���N�^���N�dI��s��h7�m��ד)�^L�zr�f�yߴ�?�ǲ_�V�7y��o���5w���ܕ�E{Έ�n|��4�Duϑb�ɖϲ9�Z8:5ǩqۋ�Ho��d�+�����W��F�N���c5:���1���q��v�]e{�/]����=b���k��c �<���%��omq�s�b��S�����u������*������Wu�cqG)M�j[R��,�8�>���+ĝ����֣�w"�t�1������~�Z|ic9E����f�.�}�ET������^sZXJ����sͧג����:�����#��� d�{����f�٦Csq�*슩*%z��%����L���F��Ë~�v�</��H�ԁy�EE����x\;�L�9�ِ9��0!�85���C̓Foէ������ݘ|���}��R�xր���꜑y�����{�@�Ǖtt�tG���=J^��S;�>�^��&=P�]�ɿIQ��W�?e�MzoD�%^<܊�SR /\��� �x����#�V��wǠ1k(�5
}�1q���)��nQ[�up�^��t��T
�Y@=.K����z���e�;��Uk��]g��cc�
h�&�raSչޥIo���X��ߣ�*��ޚ���
��ɥF�S�x�T{{k4ü���O8�%Q��$,euw���<��_Zު,�����q���s�lS^�<w"g۝�xn3�P�-����<�Y���;�g�i~=7H*�@Tr�o�Ȇ��x߻v�_����k�֝��ʪ�'q�M��xa9�Bomd͓��n��.�|��9h(�KJc���ЊWQ��,������71'sn�J����ˡb�]8T��e�[_=t��R�P	$Uս��3Y����|������y�s���s]ݤ�56�Yǣ*&�n�Qᒭ�yA=7E7��8����ޔS��b9�`wa.�؟��{�w*˧n+ۡ^���� ��:݌r�`}�R�{ol�F,�<F����>8��k���"(�&%u__f�[�Ə[��)̔eB98)�ѥ+���š� ��7��鵸�(�w3hji����;Im`��%�T��]MZ�;z���f%��9��<�PK�Rf��73�s������V.�]�V;�ǣ���Y���'V����&�/�7;Bm��IJ�%ӱ�Xyf�y��"�s#k��Wz��ߗ�������*�˾�X�O��_+�ŵD�]Z]%u- ��H����V�ϯT+%K��8�x�[��V�\�^q��p�`��\ �،�޲��e�6o1����;y׼+�@-��Ԇi<�=��w��5���Z6�΢_V�w�Z�~�y�Χ�0#6���Q�Ӵ�r�wA�9ۧcP7�m��H��`9i��B����W��3|�:�j�7{���Y�=5)��6-����uc����5\%7\Ɣ=�(|W:�q�G�j������Ff���t{sx)�b�ɻ$(u�hBo`���+�J��X#���S3-gM�ػ�uk�U�OX�V)i�ء�t)�*����':����oei���TW:<�I�r�I�u4����swX}��<�y��c���<�e��]ɊS�M��8�b��Hˢ�mm�-�"T�VՍ�f�֮�
�W'���R�;�Tfa�V+����nWҫ��IJ� ������'f�|�ȷ�@%c6�șBaまr�G8M���)�>��4��W�
�+p�23�\�Աuou���=\\t�̘M�z���jŴ��;n��]�d�H�%�r��ɥq��R���g6'J��n3�w��>�L�Nr;��ޜ�h���s7�v^¥�z����+wM�WW��M�mݹπӖ�g-��钅-�لr��iu���Ј|gf;v2ZxT���2���;��f��X�N��ձ�H���Q=m��s��S��R�D�fǶR��z�d�=Ĺ�����2d�h�v���Ӈ�Ի�]t�A5�2�7�+�]�ģ����Y�S'i�ڕ��ܥ�+�߹���f>���[*.wz���@)�f
z�\���6�DQޭ���1&.-�c*�q����Z��Wǉ��C4���u��	hؖ[��{�]dW,/��J�^��KSV��t:.��*.�Y�r��ۓ�3& ���wnO�����R46s��ؙ�[S5�Xx�3���v�<zhPP��@ 	��b�A���9�+���s���#^8k�s<�y<TE;��ix�Z+��Q������nW,wcQ�E��\�w^+��;�(����us�xܫŹc7+��FܮEEG1\h�����\�#W��<h���lrb�(��ܶ�+�F�o�˨��<�cW�׋\��%�x�q�nsn\��x܍s�2+�@B�n�-.���xԑ�xw-�s0ܹQsr1�7wU������7wb��Ƹ���"��;��5s�\�����.hۑ���r�6��BmÛ���L�ӻEssN��wu��l�WHܱ�آ5��~��2��&��:�j�*3�����Ԡ��.�]�-���
�M���;�M����m��!k���4Uu]z�J@�!�t���\�p3Ǿ��Q΀�N����Tj>�MTo���8e>�P]ly��7=3J�=��};���"*�2�����'}1��r����?d
��^~�����33㊽��>w�:��@�7�^Ol�y��-�����������X�u��2gȼ���G���+3�'`�Ok������~�X�#o��;>����T��M���	��@�͒�z��L�o���j�����u������`�o�|�g��{����S��v?Q��e���&��LE7@.�Wlo����*g#Ϩ��;����5�\M�I�\O���������g�J����CsGҀ����{/�ܯ_;��w<�+��ˁW<ܺͨh��T;u�H���S;�8:"�n�_��^���u]�����
/��.��ľ=�S#
���@,-9����|�_�Y9ģ{�<[X�fy�Σ�R�O��{���=��$
N�y�0x>��e�����i��3�<=���ur�K��{C��of"�����Ͼ���q���zH*%��>ˏvDma11MV��|7`�qu@�G��ܫ^z)�r�Wd�k^�T�)<��d���:7�����yu��hؑ��;��l[����2˖��	��_u�qʅ[x%���{i�X5��K�kq�Y;�q��]�ʾF�u�	i*��T��\jsb#-�^��5^��{ږ�j�Vم_+B\2j�Zħ�c��W���c�vN���+��nĪS�5ws�����t�5Qs���'D�����%W��*	B�UQf���ȿ/(
�R�O�ވ5X=�n��W����;�[����^��-�q�/�����»��2��}^���B�,ߐ��UV��}>:�ey�\I>��X�c�
�����Ƕg��|�Q����z����n*%�=���W������:3G��	���P�6�v��3�Y�+�r7�|X_'p&�{?*^��Ztؽ�ۿG�����~�t�W�Ȃ�y��*��h>U��[K5�Y����\���:�{]Nq���Gn�z��˂���� z���knt/z���ܣ�=4���*��j1]1y3���+��WW��唫m�P3��Ԅ:����7μ�o��ë�6�}�D��]sq.p'957�'���R���O�k�o��>��^<�a��w�N��#�=�{��/�J�.�V?Q��q�7޺�d�I8���@��E�T��7�Cjr;�P�:H���x�9�|n=W����,��k�w�?';�
4�]��n�B�[&˓�����
�{S�Y��u�&Ј<�i9Q�t1X���BJ_-��إ��5k���am�a�Y5�i�wW�R\�����l�j��G:�9��)}����I,}K��Ʃ���ܕ�|�����S;i��t���񝣮�/+�̀�o���$^}.�S>f������ߥ�}C���n�M�s4S{qY���,�7�Em:����,^LKF�bX}�R2�ex�9�r�s"6|}}\�X��s�\F�v�w��������e�����wR�j9���o�ىA�͓O��r	h���xQ� ��̍ہ�5��g� �rݦ�WF��*�����p*���H�)Ȭ�{y���=�-�F/=T}�Y��`�6�����PX]`\C�Xo=r��x�^����&�ƥ���Fp�cW$w��Vɭ/O���H0�w�l���@Os,z�{�`c�9��-t��5�az����Y�M�q�Z����fkKM���kk����5�%�{��j<�-���}j{Q�n��NT����/
�S�ǲ&��͜��:'ƹ���L	��\x,�}� ��j��J���|�ۥ9��꿼�يk�+��gnv���{��5���r�Я*M�{i�w�9`��ٮ W��`dCU�+�+�h�����D�FYP���[P����Zz瘟7X���T��_�^H����m�D�s���tn��
�d��-���xֱJ�� /�i�y��^QR�c����n�Z�
xn�pI��>��#�v&�=>��ϮGtt�P�2>cz���s�7���!�΀�N����h��y�p���27D�����ҥ��T�2�eX�a�Q���G{&u�2�e��~�iϷ��Wz�3OB�;�[Eh�p/�3g��nq�,
�a��V��=�2����_q���R��v#���Y~9��WL���;ԝ��GW�^����\�g"T��g��Ȏ��,^L�}�s��-��
��95�Gz�y��O>1�>�>�������ϑ�,�c�N��] �>���-�-��}L+�=�Ǣ�jN]n��U6({���dw�)���t׽~��ϡNx�<�L���e@}�U#D�R�&C�Q�O��:�rU&�8����>}=���u ^���^�R{��p��*#f@O�x��]+\hu{>筏h�D����gG�c�5���κ��}������p�����S��N�4&OD�����c��D%���eL����;�>%��������M��O}+h�X��7׶=y��V�&'^}���"�]�w"}��ٹDz��#~�;����aםV����:L7��=,���em=W�]����`p��U�o`�X�r���w�n,�!��̱B�^�u6K�S88��7:�EoM��]�|��.f�I��r�注V|,�g\��c�0��Jߔq8e�ڀ����e���&�J֌�S�.C{������2to�N�(g�۟�>���� 'S�=F��������mf�q���u�v6��{�c��`_s]�Ż��'��+���k�38}�� W��]�����"�͆�ET�1^4������j�zϢ�Ǹo�@�H3� ��*B�UE��I����ѵ�5���'�_��:va�$k��9&�����})](���[�8}y��� �V������xOW86�V�^ڞ=�O�u~2Bկ�ă�/O��O�^V�u�KW7��o������	��<}[��#q��H��<Vlj�ᚵuT|�ԏq��ւ�*��ɭ.�g}1q�Bsq�G���}z��Ҩ�|\��1����m �V{���Q��E���-������"�X�u����/:d6���`.�O�#0ϴr�SVl{�N�=�{+ȹ�Q���񅑾Lܹ�ZI�moO˼z��qcU��>ɖ����{���.y��gރ�v���O�ؚ6�~�y���� ٘����M9��8�ou�X4xnKfpǸ���P�I��=�o����2�^F��)�f)��p}9� L��ݚfGD����Ktj�.��7��(�}�lE�y΁���R�.i�CEn��u�(�&�,1z�{���p�gx�.��n�Ź��<u��m��@m���Z"�Vr�Iol�w�Rν76�9;9�:-�a�l�y;Y��d��G��r��~Wff+Ӯ�U��VDmCF�����\zg�L�G�����=�6&Y����ō��5w�<�J�Od�;�x��GT��9����F���κ����Q]�����{ip���[Lj��	9�tE)��PZ8`�[3d������>��rc+��W^�P�����%^X�<W�צO� ו��_��H��k���gΰ���j����o�g�z&�u�}U~eb z�{f��_{ޫg!Ϩ{�%΁���O���*G�qM]�ݛ���M�]J;���>;����'N�d�Ul���BX��T|[��E���#� s�F�'ް,�����u%��|� �W��}�څy��7���F�?Wu�p��Y��'���V�1s4F�{�ﬖ�E�oWG���ŏ(䀰�vP�s��rr{K雀�1����fs����Y�F��x�[[�^{3�|Z#�>��:�:�Ǿ�Vkig��r7�|XP�����~��\vl���.��<�Ι�,��U;};~��o�AR��k����ud}T�VMic	�� k���k�1O=p&��rU�-[YW���/����V���3짮6֨�V&ɻݽ�96#��ݸ���� �	��S�2ņ�KǾ�]��n�s�����V�l5�Ǆ��ް�rV����z3�7e�o�'DLeA�|5wv._"Wdw����m-�����0b�^N��ކ�*=���؏O���hvDw���Ǧ�'�0��Q�5�遃V��*���=�J]��T��h�L���G����~Ӿs�:��W��Whh���R>�*�,�n|�گZ���w)p�޺�`�}�,/�����Do�x��{=�p���b�OQg�5��Ṹ������P�62X�"��y�>N{����*3�\c���s�>�1��t���ٽ�Oo(_6+&B/�d3q�T숪��.�r��5�,*����[fnxgt�b�ϸ�U��ܫ�6+���w�i����Ǯ}E��ٸ���dET���W�Å�����S�tiOvVk��������,g�����4��ypE_����G�O���bP}�T���Cp2vDl2*;M^Ɨ��Q.d�xN����.%�[,�������$l[��r��7�����4�eBb$��z��v)����fS�q����1�+|gã��g�����R *�{,
������� H�U��(�����77(�V�d�i��Q���4�L:�w�l�����9������j~����U Wu銔X?j�?ms���F(�p�ef�ua��7@�3҂.������W��f���˄��P�&�vG��6��m�>6�+�tg�Py͞:+��$huY�;]�}en�8^WtB�o{���-x��D�(�OBq�V[��k?����|?>�W��L;gNx��D�����z��㭕Q����W	����?�Y|I��"k�����>������f��	�{Ҫ�Q�k��q�����쁑�^�7��W�m�(��W���W��[�Y���c���1�>=���F��{��@��V�0���.����~�{�=����D���}#
Y�T<6������蕲���n�=ޅ��Y�@���#�o��i�����Gy]p���<=���;s'�Nե]�*d{�_��q�'\�@L�L����C�L���7ƾo���_w �c#�{n���8a`^o�� ͏�"�����ø�ɔ�.2g�Ӝd7q]��~=�f�}�*�t��Rr��HGVXh�j��r<��+#}DS7� �>��&"��s�X�[>Qΰ;�l�U~�L��kݦǾmC��ǔ��^��tY�8�F���<��Q2��ԯUӾ��Sǳ��<��r�c��kG���v�w�Wȍ����#�T�L5��Γ��UH��+]{�70��N��-t+�#r��:�6��Y�<��5��[he���]��N������$Еش�`]�B�ڵ]��(W>`���ĵCgs�yJ=k��쿲\��>���zb�((kr���)���r�J�����j#����W,��U�VԮb��h�X�P��噤�~��E,����,t:�$s�{��7��8^z�z2#��P�.hy�0���D�^�P�'�����}FGT�	�̃ǳ�î�x�mp+=����Yc24�)���_��`�^�#��q�W�gՔE3�s~��%������X^>�~���xB{���rd����,
X��H� 4z��~#r��D\�2+\�`,e|�T4{W���}^��vž$�]{�yN�ot�����Xw@R�ר�)���m9+�u���U��Qxlyr���݀*���8n=Az6h�+=�/#>~����~���^`J�~�P�{*n�5�t+)�[@�V�v�~�}ρ�ڄ'�^���-�zO{�#�/a�蒎_��;�uz�q�3����f}	�G�aW�yU��g���~Uꊎ^���5w�\sە"��+C���`Z�bFfyﷺ����G�L��p�˜�VT�r0�[��:�r��!u�Z
v9�{Q��q�+K�E_e>�{jGq>61uSY5��;�d2���_ڞ@YP�������X�[w������%%ov܎�:���w�Kip�:���Q��J�'8v+
qUH�������[)ASA;{I̔���|\;gT��6M׻k�m�f�d��T�OR�]������|�{$z@����o��Gu��9�EBEַ$�{��Є[N�j%����9��,z?��c���;I�Z�?R�x;��_��<�;�	Uig����q��s:���dl�*n��R����3�������9Ε�^����W��T�_V�9�'��RӚ��~�sҖ�yT�{�G��,yt�,(<�z3����z�:�]��B���P�� �g�9� ��ǎ�=����tF�P���\o}ꆡM�������Q�_���ӔQ򆖠���8�>s���"��P2.y9�dmCF����i�zB)��D�}������L������P��O��]%�i�71<�eL���q��P���U�T;�n�xT����v������j����Q�3�V}����S�q>񽘔eV1N{�FD�r�Cӯk�B&�(߯�ޙ̧�oFz'�����+��{Ӑ�ub�פ�T�A�Ƕ�ud�>��w���~�䌷s���� �F��<����4ͷ^�=9��W�� W�|j}.+ȣ5P����7=`]TT��d�M<��
���|��=���~0�;�|[����]P����+��;�E��v�[��w�Y/V$6u��e�`��#Y�]c�6��]�P!���ǉO��WlWsP�[4m<W��.�(DVJ�wyV��*;mB�p�w�rV:��Q]o��������S GDp�0^`����0��0Z/@Mv��-HzoV
j�ܲ��N��$IC(q97.��d��ݰ�k�vv�fV���F�I�{�Mrl$7�X��n5=��t�ٙ]�8��iDM�6�q�ݧq��׹�Q��ֳT˫�D�ضR��>ynj�[P3��y�y�� �e�O[�4�u��B@�?,�[�Q y��г�
�hpW��'����N�}�tT���ǇG�Y��f���.̱y�M�l�LI�:�o焝7Zm;
��[��t�Qlo�
��nb�P�-���8,��E�kl���k4�-5�t%�O�&�G5���\Շٙ*sY����f�`����R��:�]I&z2���7�j�V�	�gD�:�Z�g[6.7�rĵS�*��TɣNZ�K�-Vm�(��\%*�]F�)<]���d$�@(�n�P'�5,�r3��Ŋz0k���Z2��e����H�Ȓ����z�(0�Q�{�YL�[-:�Ȳu`�2U�R�����.A���P~��1�7'Nu���Uk�%7'$�sm��0�n��gh��\i;'6	��n��Q��.��Iuk%���Ԛ���=��{LU^�+:�����+,lӚ���m=2(Ң��D̫����0Y�L.9��%uCo���]w��������G]����Y�32�}4��o"��+E�;�8@-,Bw]̮�@IxL��VXG������d������J����%� ��D��b���8�س����O��n��t�EVS�Btl�����ۓU[�3�:���Ӷ�.��"���2,�sr��{�E�3>W��ܠt�<��\�eܶ�wf�t�[������);�tn��3��D�]���nE}j�XCB�l��%�`۔��m]��y��iϹ����ԇt�	�gxr �����Y(�5����G;�H�0+��G�9L��
��G5�IܹĐ��,�ąn��]zJ��G�b�{�ۤ㼉5-�VSt����m�L�Yٶ�9�`t5\jk�ن��]6�N\4�͞�7�%c��u��S5qW�^d'��z�r�N�^���c�lL��S9���z&r˧ȝ�'���J��kZ�=�u�}���!���N�lW���p��])ݵ��M�%���]�c��U���v�q�9R��[\z�Ӿ���ص�v�gZ\wf䜳�Z�:�(��u�`�U��y:����,bi�}��R|����
#�n�!�G�gK��O5�<3sd�w,��E:1W�eZ�o��zC�6� ��!�ᛛݜ������_bGN�'�Q|J�l��;ܚ0c��w�*�l�x��e��Cz��+��g&�=iM����xqB�	nh��=�Wn�,��x� #�3x�oƯ��nr܌nsmʋ1nU�ܮk��J���6�U�t��Ge��ݚ��;�W7-r�1�gw)�nk��ww1�d-';������ӝ��N��8F����;��wG1r�E�[�q��q]9��n��qˮ���Ms��gu�v�A�r]���+�7KE��i&��6��-�����wtDW�n���u�$��nm�k���ݵ˛r�;�;(������E�t#�ss�:F�W.��wj73�sEs;��˻�s��ܧ]q�W;�wQ�.n74wqs����Fu�.\���2wqlRcm�wk��\�E� ���p']�Nkr�Evdۥ�p��r湴i�s��2'w[���]ݷ-(��E ?P_�c���楨Ӯ�v�%����/�!12rS����js�����7�qF�gK��"ui��*@@�9i�	�(a&9H����7M��M=�O}{�`f��~Q$|3�Q��j7~��QP��d���1�����z�I��gp��zf������vrzv4��kKc�������۬�rּgqlץ\�������]�n;�N	���"�Q�_����Yϳ�g�>��>0|����]\5k�����}�kz`o�u�S��3����N�>"�wERY5�*/Ӿ%�C�� h쇝>��vq$@�H���`�}�z!��w�t��w���zi����'��������V�s�gǵWhiu�7ޡ��}��!����}�u�{c��q�e���71Ѯ���ɀ ���됳��O�i��&+��׆{��2e���F�^��~�������=C�EJ�Ӑ��o+x0��Hz��w��C��{=F���T	��)�B^��eD�t�F9=�P����8����׀���mv���:ʶq�5�tyU#*%��.P�3q��U��7�;����:�OO���ig!������Og�a����<��Qc6b[72��/>�^+|\�������ʿ��2.n�`��O$�v�n�X��_���P�x�D�e�ޙ\ϹP���\kV���sJ�^�vW�zA��=��Ѧ�g��,�V��P�]Ғ�ӑ9���$�`x;E�P2���dH:��M�-��[�w��]��s<��������o���Tu�(�o�k���x���(�������lT/Q��=�?w�Q҉`�.Mj��4*�\@�s=%�P���A[^g��+>��@w�ȑQn�@��������C���j���6�x��f��Ru���wpL<5�xO�C}V�|��� .~V�a+j�����Ey�w%�@S����eU�7#r�w��8���T&/T���@y���<��nR|zwE����q�����<����Jj��ǁg��z#e�35X�B����F��ps�9�IuZX���Lz9(��q���l����,�s�O�{&��͜�Qg�7����w�Qx�1��}.����㇣������{�Cj߷�@<:=2Q˜�yFW���i�Q�2���nfW�]��=�g�|5t�5Mx�P���5^
�ݗ����+E������s��}����Rڳ^�>`AgޥQ��z����@�}Q���NwǩG�C�,�~���[C���rR�ol�u2GzY�OV�>���3�oӸ\F�g�n#��*-�g}��w����{pZ۫�W����s�U8=_vTEd��4"��s�G�V-�'g��g|�Yu�`=�ӗׄ��7�"W
��ۜ,^#H�qڙ+�<u.
�__r-U�tr�=&�ĵر��w	�v�5��1(u��P���o+�T&ց�{��q+�PsW,5~��>�h���Y�U�7޸w�,�E����	_�{��'�"�y��HWTNW��tK�<,��w��o���ol����L�X{�U`LEO"*.|�K��6}'�>����/v�y�8=��R��O�����q�(Ư	tTz] �"�2b��)���	�c������;�,�{(��ΘU��CjP��}�}�Q~�\xwǄǫ�1+��p��=�w�Y�O��{��}�G�w**,�Sͨj縱��ԑ������~�R7�z�n�s�f���mFߞBx�$̙_�;xs�Z;F�?I+��:W�7S�����Cur��o�_W�2�;M♡� y_�-��``:;f�G|r��(���cڟ]�1�Z���].�ȭ�P�b�����7'�O��W���o+�ARGO��5��?Q�21z|7��X�Ǯ$���-^�Y]��WT=��ǡ{�'f������s�1R�AU�k��eߍ,�s�=�����0j��з��<B�|�T9�P��]��	����. �eQ߽S�{"j�ې/θbl���*���c�k�uq���Im;�DC�!ofrd��������k�ڒ�\�Ҙ��3���;�Ҭ��wB��R�qt�lq��C\�g^���{�{:v�YxP[3)M�a�N�DG>�A��e��䕉ȍ���b�j�^%�_f����
_�����O5P������TY�>W�+>������5���n��LN?f��U�į3wL�����Oz"}Q�7��U��V�>�龤 �^��^��W��v�������@����v�����=c,�#��'e���ۅd��Fzo�.�ܨ
^����q��WTͳ�sou(�ϣ}y�絨�����Ӂ)�.��}�L�.5�gA����[��s<$���b=�w�%:��}��~�Tm�{���;%#�>��VUE��=����>&�O�+��cټ��9����{��s�;�����:�q��P��UqRo���� �,�!�7F?�]q�vJg	a=�ey��do���}�W�\:�A��8�?I��X�Ɠc�����p^�{蚋�1Z�e3ц��B.�:؟��T`����îk��׽9�VufH^4W�KMɑU)\
��^�V�4U�æ�i�zB)�����|^�`p"g��z��f߮-<�Qy�@l��1)�ʙQ3�7��~5��T3ò�����&r�b�~:'r\hJ�3��Ư�l��ibc���Jer̹�/�0�q���շ�B��D:��"�>��w�tf��p���7i�.	z�%]Ww�Y�H���b��f�Ep,.K�3YRjC�ƹ�'"�2Rk���3�^�X\S�7��z=�D��ޢ����9�&�O��ىA�EV4�ta=���ж�Ҧl�h���w�����,��~��
��{2U�� W�*%�g��Ud���a�J��k��q4z�S�G����L\�҉���Y�l�s�W�w W����C�z��?N�x#�݆���c��/ղj0�>������5��>/�yAuC<p��'��܊�P���t�];���ř�eWvA����nmC͟	��ƺ]U>/���y�vE�o��d���*���P�}�*l��Ĕr�]B�q;,e�p:��Ɩ<Mi`L__�=�"}#��M�_m>��mf�i�/z��/�g���H'��G�Js�g�WFO�i��#}5\{���~���o� ���1�O�n}�*#�v��v��ߐ�¬�������[K5��<��y�;���ѥ�k=�{�����q�!m��l ��{L���o�h{#�b�-�L�wp\��f�Z����I?��_�z>��ׅ�dγ��uHcy���o�y�eGT/]��=�����>��w��9;#��dh=Y�v�g\	=q�pQ^t!7�W���Z�O�{��~T���!�$hgc;��%i"�V�jZN�I� Y+O&���m��J�`4Ubӳ+�gd9��x�Uǡ�:�	)g�\��t��Ιat 虶&��D�������5����p���SsU���x�q��a�Vv�Ŧ�T�,X�sһ!\�+���/>�,9@7=l	�Uk���!/J�eC�ΐ;܎y��ɚ�zLS�ҍ�|�}��~�nK.1���K�eT��t���<��J�K�f�FZ;T�;�2頽�����<��e{��t@�r|.2�)��K�H�W����C�V�u{�
>�/Ц��������ԋ���HQ~��*<雅�x���0P{X��R�}��u�c�
0��F��g	ogr��=�4��3�������WLz�b�zϧhRN�5�YȻF6o�/`(dq!vϢ�LS�ѱ��;�&�>�U��g�� ���C���.�o��&����&���O�˂���$>�Vɭ/O��xiP�|�SF�S�6��k7�2'�S%���� ��T�_��H���T^Vy>񚍗�ɯ���y������;x��pV©�����g�J�zc��L�����z�l{��^���?���k������1�Y����{�j�'j��E����"f��R����SK�=]��ߤ'i�$ʋھ}ګLl�u(V"�+O����R���ίI���hr껛��v�͊��;�5�Ǝ���>*�+�""5�iPN�o>�r���O&L�9�	ܮP�w�f�7�u�<��]	
�>�H	�o!R@���s{�Ch��A
5��W�ª��3�=�*��ȫ]]{�����O�<<�kM����}L	SL�Q��~>j�'��vފ���p�����\h��rT;n��𳾗Q�9;1ݎ���} o����t-u�=O��y:B���k�����yз�mPzǛڟϧգJ���VV�;���M�p73���}nS;��q6<f۪�������uDgc�Y%��,��u�AYV�_z��dι��'ԙ�2��#��"x�k�f})޻>]-��~�z�v�6��g�o��eD���U�5<���"�d��@�|i{ٵ��Ԡ�zY^�νρ���G���{��6��ì�4����W��9T슬[�Ʊ?t����[vJ e���Fׂ��ա��KV�F��q�����#����!�9�+�ߡ厉񊮮�tO���*�`:��ϸ�dF�5Q-"�:�6}���=`h�v�Fk�n3��{G����~�fB��l�	��Q/ְ�Ĵw6a����n����\
�#NV��� �ឌ�$���T���[�=����Wk"����]�]�vw)kPqb`Ֆh��K+3��eA�����G_�At�N�16��ۓ�R�]�ՇC��i��R.�*�v�e�8��.3�y��495��Li��V�C��f��T���^�e�Q~���~t<X�:%3��e?S��܀|���^������r�,c
���d�������q�7�yH
���}$l�����ܢ&)��CY��O \�������� v����O���������G�x�+�S�w&���mf��oyP��W�&���(}�d��XuqԆҚ%�J��9��yNO������	�~�iQ��O����)8�3�gM��@H^����1כO��zx��<T�dj�,�}^������8j�Ug�*����v�^�u��ŕ�ڣ���B�x��כU������ �^��3�"��
F�M�5��ζ�����t��k�������/�x�֍-f��۬,��S�9G��ۼ�,p{v}�ɡ��Oj�_��#�Q�o�ݞ���ݶx��Ԏ���X�ɭ.�g}1q�F�^�r;%�U��¶��Z����G�R�������#��WP��5o�����WEW���e�������㩯n���g��}�~+:d>��߼td{�y�e{���q����Q��L���2�ߘ�5Q�Nl[��"|��������yÙ��_���î�7��-ygB�ݝg�+��a���2٘���O�8����^��F������[ԕ�Hͧ;�8n
W5�<���YIs���+C[N�^f��[�͊=���C�Hڜ�Ryf�TU^��P�(�0=Ұ�����c���xX��ף>�(�2�#ʼʤ����eyE������/Ozq
#ªN�j.�y��L�0�����8�H�ả}lpŭ������#������Y�Vb����h#�G� �\Q�u���/��چ�_mCo�٩�s��kI��c]��/�����p�{~�=>��칠"gd��*��d@,/͟"f4_�7¸��z��-�f�kT���E��ZE��%��]�Ȩ�T��̯�bP}7DdS����n��aȭ���앱�vzl��GTy+A��S�����S��N���pv#�꺒���k��1�ᑽ���;�_���>�c���tozW��h��	�[8��=ӑ.tq�f@�Ơ)�5�^��|�0�{�WqۛXL*�u�j4�O����J��_f�Y��@��2��❮�>���U�����Fr��%G|n�/�����׏���Ly���~5��]U>7����T�^̼ً�n^�ة�g�����pВ�\�����˜��+���&�K~�����v{�^�7{�-�6!�p�L�]��sȾ����*Y>��;P�Jz����X����I��D��W3�v��!7Z-p�SJ7�k%ޡԥr�$�=�a!	���n��Ar}��ͅ��p�\ÃCϸ�/i�@G�������X����Ǥb���[�8�������{��}����=BPӲ��g�����j��d)&�\�§x�<ϑ�'�N�%/=0:�r���ݸ��m�0��{I�s�S��$�z�a�]b��2|�C��>�z�wR=��m�,{~�[�� �'�1؏er1��>7�6�է�
��Z�)!�~��=��=u�y3��g��9];��Nk�x�{)������uzߩ��5oB��Sk�䐇�/yѧ'��+�����\;��l�/&;O�}?K�I��>1����;a�^(���
ʿ^���,���N˦��6�\�Eϓ����{p�o&0z��P�z�#]�����{�G��J�߆GNQG�7�����U#+�t������g�v�GI�{
��c�z\���p?|��l�w�R��k޿\z� ���/혖��-`{m�-�B�W��O��/��7�֓>�5��e#�����;n�̱��}93�n!Ҹ��>5����*��������Z�D�T�����c�t�q*[!��<�`]ď�}�}G�����ֵ����Zֶ���k[n�Zֶ�󶵭m�붵�m���Zֶ�󶵭m���Zֶ��m�k[o��ֵ���vֵ��͵�km�kZ����Zֶ�񶵭m��mkZ���ֵ����ֵ�����km�M��km����m��1AY&SY��j���_�rY��=�ݐ?���at��y�(�� ����
	
  �A@R��@�(Q!TUH��)"���BTPJ�UEB$)Uh�UPE$��A�*���RRH�T���R$�""UP�����(J���U)S��*Q��¨fjU)hb�
�h6�$�f�P�&%THP �%f��n�$�( p p		�)V�֢q�� h �i�J( s�� )@�� �,�U�Z��	�[i  N �R�Sh5)� �Em
���T���!T�b��6
�aUI �uJ�mV5([fV��lQ�R�UF�2�%���Tlh�j�f���R��Ҫ�VR�T�J� ��Q14)UM�M��6���34B�4����fݲ���Y�m�f�Р̦�ԤbHH�UT ���v�P��eH�L��P�ڪ�p��RU�)-eZ�e5�-eR�5*���آAX��  	� Gv�%(P�hi�R�ؑh�J�����K)*Dl�ي�5����,j���R���"  � ۴���l�)J6�k@�)�iP�el�k6�)���5 D� � �I�Ҡ��d����PS2�i�	,�V�R�)Y��U�����&LfUV�l���FUI[P�V�F
U��M��IH��� 3A����    ��
T���A�h 4i� �Q4�=$�hzM@�    ���T������ 44  �$A 5S ���#����0�l�I��d�MF��4�jh= �4 ��N`����Y�0뮄��J�q��Jl�!BCN��Y���'�Ii!'d�"B�a�S�U�xD��2Ea����+�}��0���REJ��F0�	
�(i#M�I!!��2Da4�XBB@�;Hs�e����`S������Љ���&����`g��!�������{�?���w�:�P��E�����:�_ǝ�����z{3��枚Gq����0�q�����v�Hu�Nm7��ዺ��`�������6�Xݤ �S��z73"Z���� �$�]奦ܭhAB�a-��j�ļ7�*�ujٳ��_ӺNC�-6��//j��][`k9Sb	.�V�r��n�6��z�K�f�:�'p-׬^���E��ukj��:�[��H��M�Wo�)� @۶щ]X(]���	�`ʰ��)��VJc�;�>v�*�6�8j��R��ƾ���VAOc��^���.�����-(�-��5�n|LÃeZr���x�`$u�(-x�譧�YW����Ř��؝D�b���q��C�F���o���4�ٴ�$��2��yn�yX	V�v��#���QZV�P2�Mj�+�{g7�v)��J�Zs�O6�6�K��yi	Sq��h)i�^�l�8�`�4�aGaÖ�	cP���ە��B��yQ[���[�Ѻ��x<+��WH�1�Xt���Y�A�,\��T�l�A��Z��G	�vR����)Д�
zsuf����u��)2T�:eI�����ֹ��.�YL!2��]ֺ�Z�	�u!���f�Cr��MM�F��Ф��0��6����փx��G
��YVѭȕ�n����R�
[h�t����C54@-,Ia�ו��;����|��[�a7Ƃ�@��:Z>dn�fl-�e
[���J9WE����n�*�J��k$J�7n�X�WY�(�2#r��C��#ͧ����W�!ƒ����;HaS�� �/ʙ��;��-U��5��ݵF��N�E׵tj�ޤ�n�����ӋS�CW��j���X��y(d�L�G2Ҋ���'�,��(lȵ��" �鼰
��Y4�42�ͻ	M�wf��*7��Ŗe��D��ȣO�a���cU�oSw@Վr���jD^�W˻��S$p�v��#w$�hhk �dѺh�x�d�~W��e<RE�R��<�u��S��-�۬ڼ��E����VR�hu��8kjѳ��|xߝ2�.�O�F�j�l�OVճ��@#��(*t@�n*7F�����[aJ8���� �����yi2�աA](n�[m\�r�v�^T�WL^�5h0���/P�;���s�ͥh�;g>k�!B���c��z�}�����c)n\���P"ixH�Ű�k�Lkmf퉻X�"rVeL�ފc뚌2m��^"�z$o(�h�RA��nطwM�^ǘNt�v����'�LV�x���@żw2�֜�@�Yy6��`���B�h�dܻGZ��$^Q=�)��*��]֚	c��2�;��W��/i#z�n\��S{z��)����Qkϭ}���K��֫<�.�u]իU��_lzS˒�Ƴ@�Xܑ�ø� ��`, �|a�<b�����{[g^�ue��ƛiRkn��r�ޫ�b$��1=�e�4�F�un����� �B�l˴6��kF�L���pJsN衎�3A�"q���Y����-V:U]��TU�z�.�iu>oR�w���v�Q��gȀ�b�n�:�`rP*MS�
'n)a]�0�'/r#(�f�'�Qܨ��Sf��}	xq�f��L%����&Vm4��h���ʽ<m�6��cv�[��St	�u0 rS�]��7�H8F�
�?f`�t��F��wooKlͫ�l��P�ш@����Yt�8��^MCX:����Oe�8sw/ �n#Zٗ�5�=�f�cf�#[/um,f�B�0��]fb�j
�QLZ�����F��ED��(�Ǆ�Ԫ����j��[���Š]`��;fma k��2��̕��4��>�ff�(�.�M7%�s�n����n��4�J����KّP([كh��ٹR6�Pf����m��Z]2j�ͦ�X�._�,;�&�]��c�ujq�<Ri"팧Y���Z9`h�F��дc���#b�V����3n���>ѳq(��r�B�� K-�e��Tԣ/w0"M+7r���m�ˡ {Dަo,m�1�ͳX���\e��7�Qd ������wuv��-,V��c7t6��;Ƕ0R��l����:����s/("z��*��.!���V�#�wvk.�&�����vx�1���K���F��ݘ�Jy؀�ǰ�i���Z����WNc�%�5*�B]�h֋E��8�MBʳ�d��Sa�J ;�ܒQ��ɚ�8����էR�Cb,r��Ն���[ibA�)]�e9Z2��0h��houZ��`���W��I�
���tz2���p�D\��e+7u�&�d�\M��	J�%�v伨̭ǂH���)d� J�EW��Z 2���-�O/% M=�i���)5	_l�[& �^=z�sR��.�����y�QwZ��l�CAd:���Um������1��+��QYB��[������ote�2���w/D"^�
ܧ,kNHŁ�s��]�c_a^���ag۔��ډJV�Z%��v�{ylQ��Ƞt�A���u01eP
)R@F�VD+r��;�pm��#R�f�J�Y�Mݧ���tw������w9�8!Oi.�A��݂�m���!8���;n}v2��,!��J[�{�A;daA!夯&􏺸���;��+6���[�R	��u�%MÛW4 r��3Ag��j�KiS�X�ݬY{���y
�4�R��x)�tq��C���Pջ3Vn:Q+q�қ����d4�A��cmU���h��U(��j�/,��i�Y{�h�㠑ߴ�� �l�&n8D�/U�X��ڒS�K�X��#W�ٲM�(�K2��^f�Z�������]k׉$f-l�7����u�hA���#kmݛ�X#hm7u��t��S2�/%Z�N�@ef�uCy��ڤ����1^ɷ�y��=t_{��j�����y*[´Փfi��X�ǻj�JhI�q�0b���G������VIZΝ�/Y4����Z�U��˪ԁ�[oFT������U�]̷t���t��X���2�"hУ�h�Ő�$e�"=6�.�9���ڲ�Ǹ  �q�oq�1h%|�%4�e�{�W3*��n�:i�4i���\�/m�� &eJrī���K�Y���ZäDVR�Y���0+CJ�
X-*U�K�;,����@��e��͚`[z�Ԩ-�Md�WY��U�vva�X���]ob�9�;(Y�y@ ��)N�[���s�L
�su9�u�t�����v��š�U�%��QTax����8ɦ��sm�{r���l��jjX_I%�c���n��Aj)�דU�[ӌ�t5��[.a�ʕfT�dkL'0�"ԁͳ�0�,��se!�nh��Z�m�݉Y
sh��lG),�z���U���Ʉa�-4�j�c��'�\����-���f����'ǯ���aT���$�`�ʐ��u/%���v�w[��uk�r���!��v�KR�܉�h������Hkv2��5mT��fMV՝�[E�[�vF���cto���^tf�K\!t�u�C6�OcM��Oy�F��	��VL"i���m"����6�H��l��b����6�U��:h�U����W�l�����^u0���Q���z�;Y78���]i�Y�A+�Z�=XVV�j�4�f�� %U�B�]��
�ـ�)�qY�!�����7�1%񸞽�nѳq�wZ��fH����Q)R�
r�^ˡz�����{cMڔV[7�8֑���E����[��H��H^g|����4P��,Q�X�6�L�g
�*��㛁|Mw$�- IB�ڼ��I�o	!٬g��e�V�ei�h�
�l˓R+vL��j��uF-�m�WB�Vf@w.!x�#���8�ѭ��.ՙ��	�̲U��4G�I%�ʖK�5��ޫ�X�t�fU>�4M-�]�]m�=v���T0��`�B���F�ǹf�*^�*m��T#Ou��i^I��gQw��U��l&!�*�\�b�BӚ2��,%���3���D#��`�CZsF#���f���ş@h髤��B�Zs/0��Om�f7����O�²�4��r�#u6
����Ei�ަKj���r�ڤ{��ZսG� �w���P���Ƹ���a�FM�u��I�@�M��,�.�%,�:��I�iԗ6�4\5/4\1�l�0�BJÔM���el�p6�k�y�v�'����Μ�/pnkH�@���V�f#c!U5�3#����}_������[��5��5�Jy����G��9��Q*��g��ܿu~�^��u]~�c17��3�#��i�GyڋK��W�9�UrM�V�����Sv�}�Qv֊�(Cn�����'�m\:���ʙaиZ'6��
��M��7�a���ۭ7Ҁ�bڹ�	ɷ�3��5�5�V� �J�윥�������ѝd9B����,'y�ۓ���lBԱf��r����-�
/�	K�:��se���F���
���y�X.іvi8���/b�M��pr�'{v$����;V��{>���x�ӕ 6�����7^X����eM-�ãZ��|j.�]N�a�3�sz��hV໊̐�)���O@�F6�ډ=��Ѻ�%Mu��Y0Y�_9b�W>�ˠ��%m�伓��u�TI�/m��������/5ͨk��[�{(�$�YZ.,��'�Wuc5kx'R�)����c0]盓E��"����1��u*,��jm��̾�B�Ѽno�7]�G._+�a���i�n�7�x���(�BAݖk,q��q#����	�ڨ����7��E�n�}c�2�͇�+Ga������gz�@9��һjA;��YGt)��������͵7@2�Wm�+��t��:�d޳�p��w��S�	�/w�;7Y�*���M@��v�L�s)<޸a�o�>G�f�
sf��;G+��� ;>Ә�΢���+L�Ʈn��hN4z�.�F�]gj�w�/P��V�\�\�ءV>k��2;���z�O���e�n�۸�e��D:��"���J�ׄv��6[���4%\QN����\�]��� <�r����+-�f�S:���7|�x�B�8�i����X����U�i�k�($��h�`��FMÃ$ �GoofMy�5���':gwh�'D��R�WZ.��Ɂ�mtvz탂ꕓ4�B˧KcӋxԆm�2��{���36U�P��v�����œr�s��l	4d�Rf��v����S5�o��H6�j"���
�'%���f�|���'�� ��c@d�$��l�l+
�̤�&��CX�� �f�X�ޥۨ�F��䷛&5�q�k��]�i�#nƛ�{�!�o-�/]����a��{1^Ҧ�7/u�M���֊
�;�85��4VCֹw��We�t`<U1�Fw�;n*?�i��ƶ9�Ȯ�NG���`s-�}R����4'LR��mr3��-fZ\���,��r�:��-�ʋ�]Ҡ���N�,�.|�0��6dCv��m��uuX%p�� #f��h|rW(�f��R�]c蛰{K�:J͢4�������}�L���U�9��K���up����Q#B�Q:���h�5�2bYQZ�a�Q�/�n��7	�5%��kd�ټ�1�h^���K�:��sb��L�g{2ʧ�d4,�aR���̵ݟZ�Z��F��5���iupx���[Y���,�n�(u��{��R�9��h׸_C�J�W�:�Iu��ل�VWba�1G|�^���_'z�t�`�hؚr�N��4>T}�嗢Cl��ehgP�������4(�� /yM��-a_$t��ۄ�����6wDI���D�F6�mv�b��������]jX% �k8���@&�mmd��;j�oI#��;v�we��ͣ�V
��n3@RW��8�[���/�h�&|f��C�Ð�PoM+���`[�j�[��I��8�Z_B��\��i�*��:ì n�on`:�+V[2�[6�7��X�MӍ�b��s,Dv��AG_\�U�=�iokזC��τ[��xcH�b��|���qg���m�V�ɺ�	�� \��'r���R�fhϴ���/3kj�Wcp�3������q�^�:��%�>�a���uٸ��h��4�����}j1ok���]��'q�i-Y
lͣ.<wo{��iI�Y�:�˔��6d���������hֺ�6fœ�gǣ2ɒm��Qm���u�װ��^�7��@v���:a;v3Q&[v�ºڢ-U�a�Cqw^u��Avc�l5u�t�м�q��g΁�ը��P����x�+���:�Vn��d�����Q�$��!7fhĄ����WC���T$��kc�&�E[I洍_G�6��R��H�{1=r�k��H�2�04k=���Uu�p.�(���m�8��=*Kù #.
5 p���غ-��7�v˴��-���\SVۢݮ`���tm����mE�d�̝s�K�(�sN����F-;���E� ��wU�\����H��(�� �8� t"�R���W /5gT��gt�0���ڕ����X���ً���Q�s�s���=��Z��t���!<|2���+Aٹ(����F�j����w P��\֌����J��f`��\d�ޭ�������+���I6��`�3h�A��F�Fv`���f�,��7���la�4ȓ�O �Jj�N����o�����9g[
0����^��X3�u�x�RD��쥵���	��|(�
]�X3:��^�c%*���T�i�^W���f^����1���Nh�`�
�@�0ʻ����̤_c#�2ۜ�6@4�ހo8��F�̄�z��6B ��@IL�Br޹9[Nm��JXո�m�|�v�n��;�qɋz�B��nG���ϥ����{�^-�����1����,�\ %mN-\�����H�v6��Ē�®�N���E'�1�=�-��9�u��'#��\�)Znnh�;��-u�`k{��F�
`���kĻ�[[Z��%�7��"�L]�(^8�mp]�c�>ݺ�v��`��v%@���]���5�l���j��.�=�͗���^�\�Ut�^=B5sM��a�Y|>Dxv��a��t��㗇Kʿḳs����Ʈ
��,�}��
�A��ò�v$h�"�iVi��*��;JT��fP��P�IAd5xpf�س7��(���N�Rg� ]��5�wmqn](_`��=w�۾-}&%N�h*O)�q��*�F�}¶�~�0bV�����,mߥ;�B�F=�����B{��+�1!5�}��j�/B=�v4:��.p�"&�\	gf�ٚ%��g�rķOa3[:�Wu%����Ev�_-6zec��'!�����9�n9�i�wY���66�k�a�(�p{-KNn�\��4�t*0	2�12%��r��4�U��n�7j'5�V@q^���x,n��E:͙.�*n�@M��.�^%}��X胨҅���#�7aEG� :���3F\[�&	�3jV�^L�:��[�G=�:Tق�Hȣg���v[@�0Y�yq�M�Y�=�����i����K�v�tt�W6h;N>�2����lR�sm+p����Y躯;.���^3w|q�x��q[\w7���L� PQ>�:q�y���/�]�V��6��=Z���9.,R�{U�J��P퍥ψS�4�Qǝ�%�S��u�#�ڊr�yit�;�E[̸uS� N,��[��1���W1�ͭIVc�j�b[2�<oW�r/Ӧ�d�������u���b��C��JZ1�v��{���}W���b<�Cu�n�kw%��Q����)��T��g9n�"$�c��:�JU�v����՘;_ni$��Im�=6).3�2֚j�Ě-�X��+3:�[�R�uq��Ȫ�t��HE^'�U�&�N�a]Y��!cc�Eҩ��3F:�Y�4坼���׹�1L�1t�O��Q�"���s혰U檷�]*�q�һ�κMי�,�0��7ZUb��,	�X�3��3P�+Z�U*G�J=sː�䒳`=P<٨�	�J��Å�y;�M��Ŷ�|l�/S�ir<$y4M�A@o+�*�E�W�3��[J�G&�G�7-�Q�]�T�9$�I$�$�I$�I .��R���R
F�e@/���6�\�e�+t:%t�L���%��d'�����p-f�NP��b�KB��:2�k�sܝ�c�[g]��R�����W�F��
�,Y\L�d��8��k��T/`6sn�u��/b-tΦ!Ӕn�����th�q��Y��9xx[Sx@��\�{�݄�}�W�usb���=:��Aٔ���on��hG�i�ۤ�=�1���-���g�@Sa�su¦���Q��K���/��%�ҥ��:�LQ�D��69�ZH=�/.��v��
}��V���
k����R:����16�.�a����.�U�����7r�E�����`�c{+fC<�"Cq�����lQ�z������].8Z�L���T�o�qP��a��ns�7[`��r�pp�CV��>w0sҶy��Ç]�z&��e�j��n;j_�HH_\R�_NĒH��m7I���R�<��D$;*�Zs�m�w�k���V���^����8� ��`���:\�-WqY��rk3F}��m�-X6s*�,�
�c�#OVB���-�Ś��E��;o1R��������sͲ�Gn��MU�n�9�6f�y�-�;�#[M,�2s��7�ec�lh�kn���r��՝���c� +v�WQ�hՌ������;D��BR�t��ɼزax�6Z�*rL���x��f���Uo2�\v��1t�h�Q�u���g`Aa��.�&V�C�8��T�=j����wd����4'�X�֙e�p���4�<���v�c�vF�=�A�I�@4����&����,e�c���+�:U��m��7�*(NXw0
�+z�%nӫ�����/ư��r���ҋ�֤�0��2gݴ4�� �� "�}�u��:�wP-��&6<�r�Wp������:2r�Z>�Ky&���t�m���Ws�����:E�0rW}we�;��+4���|o>뗅+ү%0�oKh��,`-�&����9J�ʶ.|+U�C�HF�W�1j��U
"�-�r�a�ȯ�p�tp��k�ٶ�ʺ���q�M^��1t��pb4>I��\��B�q�'s���u0�t�+\U,;�T@6ՌG��d-�}�0�� 1�(�BM��MkK�|YcJ����ó1B�3 %H��X@N�:�>5�u}'(7����l����F��p��+���(h��V�6�CF��(L�)QU�Z`��)r�n�rx��tM@�nw�ʽt6�]+����SY�*y�n�Re���.�#tf�d��K%h%YyE����[U�9T�糑ۤ�U4L��^�[�i��K������Z�# �eۙ}�����̫6�V��XLv�ܮ��u��ks��>���%6P�Xk�ޭ�(�%�W��s�����S.��&v!Fʧ�� �gwV����/r;�c��ܩ�:�,�S2�R$��R�v5���D��uK��А]�j.>C�fu[)][���K�k�ҵ�9���!}��c�9�	�8`i�%������.����s�ф�uf5�(d�]����m�mh��;m6`�,�]a�?n$�=��A�Jl�V�7��7y�Zc�U�-�����o���dX2d%��`U��D���S�⥊�$�(�PMըj���Hk������u���m*g[R�Ji�|.���F�Y�j�V��I^��W]ܵ��_Q�%Ԥ���[Uu�q�6�S�Owf�x6�ڼ�2����x\8Iܷ�X��qʮt�dɼ�qWT�K{ܴ|^�J�Y���e�[���e����޾,+;��]8f��L�Dd`1��ӽ&� �����6��)W�8C��V��y�3�����V]�NXbi_Z	����av��X��Gi�*C�g]�X����%=4��Z��M�f�αc��6v>�q9fډʎ��ꗐ��hmCI�<�Enks�N:]��XZ�]:�1�b��F4�Totc�꾋�v0�극dtw0��s�a��]rv�];-.�����&�)qPev��%��G������(R�uʚ(�-j7�v$AX��);�vX�Bi��ٯhB+4�q�T3�.H�Ỹ.n���vG�fŅ���Ü��K�'�A��M@��gp[̾�-v;�'Q�\�m�e\�>�ZC�;�c
��/)�D��ȱ�E�ū����2�
%�p� $ۗ����֙���a�D��������s"ހ�2�ͽ�\%��ObK!�꩓���:��`*�ۺ�Bշ����[poR��\o�Q�u���X���9K�d��_U-2<��'Y��۽����	r�i�E湎�>��c�;����
AP�YH�o'9�N�2�'Fм�������k��@�s�^�L�v���mPR��wea�J\��
�|5UǢ�ڍ4�D�NN����a[܅��J��qF�Tet��F��5�yk$�SkG-��ڦm�\��(��d���»�~��/y#ښ����Ⱥ_W,zq��8�P������7N�a����=�&*;nN�	�!꼤�.[��P����\ZZ�;ɀ���Sx Μ�Mӑ*P�Vu�������Y��{ܦG��C'W �b���A-��b*�tC�m����{cN��&8�Y�*��%s��+tY�6�"��\�uW���:�MY:{ �!��.����r%.�͏{$�JsK��>���v�4PU��H�Q�`�yf�bc)��� �ku']n4ԩ�������ȑu�(��/�Wni��+�	э��ŵ�G��R&���q���
Ƴ�3}����_;��8�37)a��S�#�J�pW�*V��r��ull���^t��(�Ǒ��F��*�P[s2�+ �$YVq�GGoqZ�Y�%Rׯ/yC4���>�c4�\Y���Z�Ոh��Y�7GC��%m��	��6�D3w�_T��8sg��PCx�)�1:=��i����U�L�SL\��<##0ՔB�-g���e1۪�Ͳ�J,��;��$�����J�U����|�2��c+�'�Aٽ���n+;z�CS���Q�� �,���z��%^Cw�\[�+&s���[��҄�c��5 PS��c$"��7�P�ݵMX�|7_i��a��71;핥F�� `))�����7XRx�(u�ޣ�a�`���2r�5�6�ӵ�[Q�[uv·a�3�J;S��.�����&j�뎴ԋȕ�Y�X����|.�dlv�f����yy�����L�o][��nҭ�,737�d��rY���˻�}�7p�i�9:��$�=�ׇ���e��tjdJ��.xUL�7�E+B���L�6��p7��d�v�80-�/^{�@�qd�+����D�Ky��8�:t&�k:�PH.WV�aK�Y����.�&�E_	�񶅇�49@J%h�w֫��li�C8��歋ys���AUx�%��݀d����iU���a�s�;���e3�k�B�PY� ��oT	Wp�V�u�$�n��y��F�U&Χ�l�m����ʲ��lD���aT�S���Ji��.�էF��3	���>��"�%���uݮc�M�ஒ��� ���Vi��)�:ݝ�4ӣ�jN
�#���f����һ|MEʾ��v��C���b������.���kKZj�Ef�v�X�)�Q��y`�s���5�X��Un�s/6�S;�W�v�1	]��M�8(�L�vBz����tc����p�u\n�N떩��oi����|��i�)��*W���)5��NK��ʚ6Ȓ�5�sMG�.�ն��傉����b-f'z��N������֞�źgR���*�ԫ�tɵ�%�D�v���\��꺇�E��
"��mEn�=�dS�Y:Ԭ"添]in�Y�.��ډ�
5w�x�N��vֺU����}{�	�f�%���ʲ�)A�a�ϥ9� 2�n�iJ{@�7ڝf����V��;[����`����J��NS��v��#e֪�[om��u2�^c�V���>�l��+���vP�µc5Ʈ>�vqu�:�%:�C�}f�D��}�V�pb�=6'Ak�xH;C�wZ��J�&ܨ�
�Y�Kp�Kn�wИW ���'��f���G����g��J�+Z��6fD��]Y��V�%�9�ϫ7~5xXY���ʎ.P�K/�Q�V4hP|_}���S3~�1��>�}:�A���������ͺ��!ul���>���V�֫d�6+�]��I�u�H��{�R�W=fU�)q;*Vi�(��;*WK� ��F�8�����ª�ٕp�aj+y��غf�m<�$t5Y�V��v+){�=�P�� <�GmP�F�/Uؼ_����Y�f��q�'mu7�aPJV�ξ�kD�GhM�Z�w�KW}��Yׅ=`*%���w�*֕�����֕�u�jwm��|;kI��u��ʄ�
x��j49�g��M� ����١��F��q}f�oef�vrc�J�՗y�	YI㴩��a�7*݈2� {Xz���R��q�Z!��Ƕ�)�E]Ֆr��Q�|����D�˴�;���V����4t==Xl��P����yW �@yG�q���X:Y(e�$$˽����ވ��_7c���|<�ꎇ,D��|����>�e���zN��Z��{����=�yr�� ��T�ۛ��3C���<T���Dt�,��1;��V�k��}S<~��Z�N��7r����CN��EA���_+̳\��Y�_~��	XE�R0z�0�9���FA5�^gwJ7Z3�5��o^~x���L���*4b\]�e�X�$��6�xrh��Dꙥ_5Z�Ⱐ�7C�:.-�;��`Z�-� W�Y���Xʝ6�p"��D�{%Z���O��׌Ӽdl9��+Uo�w�W[qa�b��W%Wu�t�e��i/�])�f��(k�"+��cy23��%��
��Y� �i,��@�Ѝ�B�`�זn�G�R�X!�-�����c�*�m�*.+sC@�\fM{7�@� �����MR�����ua�Y��(�!.�Į�!��qw_,���,�/j�8� <�]5��R�����w���Z��u��8���6172e^�͗�	a<�%�2�\q�5�8V���6���#!!�f����{^������U��8�x+���\y�h��u���b�[�eԍ��hn�vؠs\������+��V-�4[��M�;!�mU]]J�}���{��7ǖ�7�o9ړ��Ц7\���7/f��7,Ё}7�����І���}o]�ם}��f{QZ�++*���o�d+�SGM�"cW,̅�ET�=���Y�����2 �WC�V�(Ŷ�E�
�l�JT�m�mE)J�m��m3
86��m����Ũ,Z���j
�U��L����BZ�
ʈ�u�`�+V��A�aX��+��wXT�X«-��e��b �ީ��Lĉ���MfAq�əVV1KlH"E�ʭ`��`�j�0U�[�9dm�W
*LqS<���i���w��-����>��x؃Nфk�g|Ot���.���n@!�;﫥�H�����}'�e�����gE]Y-V�_Mf���K+m����*��>�!��Gb�H�c�/l�T{+\�@l�+ۢ�wQ0H�\��F�K�ٌb]��/�[HjKٻF�\��"|q����/zY�^���6P�;�ZmU�y��N#�&�� �ī�;Mƻ����g�t������Б�Jx�ج-���Sl#��ڎi\�pp��滯���8XT,[\jL.Ċ�WKH;��m��;m�#��)�#j�QJ��5�}�^�W!ި̞���k��b��J�P��I��RI[�SpY���%-�[Z��f�����}k
�hC�Ou�W�ڛ�{��J��	�ld<TsTygbղ�����]3t/��K׺b�V+'V4����{a'�bN�0f`K�!Vp~�^{x;#ޖ�+��4w�z���:v/*�`2Wnk��Iu����)r��et�-�����}s�TIɣ,�5=�e�jkx�hDn�יꦲ�p3��z���VR~��O�Z���c�6�q$��_��� N�.�n��k���Z�鵚y*�Ie���D�۫���\�}�TFb���������9N�1x6h�dZ�Q��]�Кg�}�(�Wԓ3�Q\v�ڛv黾m쭢�A�������A��l��6�]N��1P7���nR�^�4O�z�=�u}56�6.�* <���������lw�)[콗�#X��%���<�]�u_S{��tqsx�F�U�'08��M~���^�x��&;���N�;p*�ݵ̦]��ಅ��	�e5W��0�G	�78�sm3��ҹ_^��+	�jL��t{���yy!����NB��â�������qH���(+i�x!��ٛ�f�hx��B�gb\�M�P�#o�	f�8[�U^Č�P:��#y"�Hk1"��<V5�����C]'�(��ͥ/�*��$"Í}l�Ĳ�|�S��$��W!k��U��	?p�)����F˯�מ��0\�o|������7}�O������â�GfE��wJ��.����"!�<��+N�^����i���ʒ+"\#�p4��1�E�I�������q�~+B��0QOh>U�٭��m���ȗ)"��3|���p��"b�1qCg���� ��ZA8��X����ٵs)I����|�b��)�T�m	��@�1��y�Ȕ�QU���=o����w�X�iE�Vy�
��C0�.�@c�y�T�77���K��b)v�@<��N�
ʨ���S�}
�9ʫ�|�}}˼�~Z}�'W,Yx�Z�T�!�3	���o���)�e��Tq�����xA�I�R��f.G��gq��ˎ��PYB��f`���rf��aA��K�o��h��s��!u�@�}ׯ`쌝\
�xu.Rޔy�/9���v#��^�t�/d��|`F�*�fy����ŒV��NM��E��i=�������^2�a>��d���gZ�U�'2v��o���Q������� ��cO�� '�j8����O[Y��̧���o���w;�z�G��\��%g,��v�5�����Np�;�QO�/�T��:�����Q,yo�T�J��v����(f	w���v�-s�����-��o���K:���,E�lQ�<���u�%quų�.o.0=QPQ��i�G��US�=�����j��K�azi��eDjV��{ON'׺�L�`��k��-�ـ�Zu���V{�1_�s��j��k��x,ӎK���{�vr,�;�3�M��}�YQ,�uJ�y7-r�yGo��Hh��i�$��СlyХO>tq7��T)�s��_&B}}b���Dz��q*55�*R:��A�%�}��|F;;�<ë�o�q�[�xM�6I�;wN�騫�sױ�`r��1�Ry���ǞgR�S"]	�*����rg�R��KkbBx��3�K��bX�b,�y�pܧ��WɦQ�Q{��g��5f��5�c��๷��<��S�D���{ɘ�)���چ8�t�Z�8��luBft��L^�}݇8�e]��h���M�.|�ҩ��3����0�Z�G��2v��<���H^]wp[�F{ �;��:
1�)�ɹ��PD,noT�}b���I�*Cfn��꺐=���Z;�:����	O�f�ʐ)}ə�u�=�6��*�-��:�\m��q5$B] \�ADy*�	nJ��Ga1�;oB���E�O�d=@S&�uA�F*���;[*��<wnVu�s����؛H�V{.H�o>��񏢈������f��	�NL�W�Y�P�\�N��ȢGU����[�) ��إt�ҹ�\���e:�KJ���#�2i��*Z��P�WvM�Q�>�32�2��#��p
�����/=��Y�~��-�ar^��V�Ὃy�o4kD��5�X��p30���Ӌ�86F���v���J*�Ҧ|�P�qp>�&���er�M��WB�-�@�ڤ%n`�a\峒�,)���}} 	HQ�E%4{��p0+o�E�嬂��WŤ�b�ȱ�@��FY.��-�ʉ�LΫ���S"�ܺ콮�Һ�-���`#�ͭ$_8���U`ƍ���������*M�L�*�8�4d�w^�_${WEIM�u�
H��	Y��o�<x������:	عd���%q�i���ڼq��]�t����j,��r:C�ⷁƓκ��HS��jٓ��J�{�ͭ��f��5:p�ط^��D�1֡�&� �v�v�Yf%���xgo��T�N����>題���Hl�)����}�������ފ��/�ݛ������Z`����4�N�31�B<��p�AB���+�r`H�Ŗw��A0�9��x���T�u��̾��n�9��=sX�U-!�ķ�(�9��AYp`�H���̸�դ�Ko���ʰţM�"��-÷lޘ��Uq��Xyۺw�d�m��;r�XǐE�ե[/]8FMmʭ�������x�9�k��.u�w��F�DZo��Z�p��/mh�Zh�Zx�ɬ�,�)#���ܹ����n��n8�0�*���mM�-2q1xZͫWF��
t��v�EO1��R{�T�=��[x����.�Vd�+@�3tH���:*z��p���q,�'T9�386���[��5d�P�x�W<�� �������$�s�r����:�B�J=������f'8y3[+�������Z���v� �˽�m��b�dJ���6s��j�a�]������k���e^�h8&����o6�t
���"�v���:�7~�UQ���x�j&26�v��d����tm�bWA�}E!���.�&�絒�c%2ֶT��.�@�>���MB��5��^N-bL��\zH	sTjJ�	ӷ$�m�itNt��ͽ�ׂ��m�!V��mZ�t�����~���b;���Y[���1y�F�i��m�}��7�pq�k��Kiמk}�zt~�>J���k�~}��]��^�����5�r�+NH�N����N���E� OHqX;'uݺ�
	�:mB��xV�pr�z֍C.�G�,�G��%�2!W<��ݭ��}�Z�������D���f|�t`��f[t��)��p
�2�)Av��{j�^��g�n�;8�܆��X(lձ�7]j� d��]�Z��f^=w�-.cV�(�Me�̻� �{d���W�GX4�p&T]�����WY�S��K�$TI�B}dX��Ԇ��*E��DzG)���1)[M��ժ;��û(��۩�M��3 �|�YpA��%�Ǵ0�jH�F��6]�������%��g0��J�&e�x�,b\0�b�Gg��ē�Y�R��p^�eզ�W���X�Y;:(��>��D�*K9sg��Vx�<g�a��mgL3(�x�\f=�5�^�Ғ�� ���y{cVQ�5,�0����Vu$���uޯ��U��ѥ������8(f[��)Pb�.�,\U-��D�Eg��:F�SI��^[wx)e�I?�+7K&
�F�:�!��ⱔ�.���*ͩ*�2;�]�Y�M�t�Ye��R1�� c�V�9�++$	��ER4��KVbxNZ���B��	e�]X?ma�4�M�cՈ���a]�7����B�P�@ĕ]8��`��h�m�w��QV.�<�`J X��f���\��ϠyBݓ*!�X�&����Y�MѬ��3J��fL�g �����y�5-a�%�T��ڡ �a)2�J!�Td��� ���o�p��D��a�s>���S�uf+L[j��2�'w��w2Ql��`a%Xs2��m��VQG��qԇD��A|�D�(�v�q졶R��v���,6�f��/~zx{�\�~?&_�QN�eg�U--"Ɍ1r��-if�5��1@�Vcuq\UJ��1ABgY��i�Z��Q#"�����VIP�QX#DV��UAMe&0Y�D�F#c*�D��TYVDbȢ�R�Z��؊ �SL�UN�U�
�J�,�EƢ�����b�b�A�c+RUY�@PQ�
�2������,�M2T��E��IX��,�����E&����d4�
T+YR�B,l��X)P�(# �����2����)Nu~�=���	�YX�G�n�h��7��kP�:��Y#���w{}�Y���t$�o=��9�;�<�Mgl���5ܒqQ��y&�B���f��:k5���U~u��3�#��ƒYA�����P�(�p�.�>\"�_���O�+t⫳��M�c��;t��Г�j_^���+0-{upCY��O�u�Q�F��w�z��<�S�n�V3�*��5�$؍44���ۢ��W%&fڵWA-i���`�l�Uf+��{q,��3X�/�S'Z���8+���a���VS�uV��	���l�����������7�&���B{��k���d[�rՖ2*��MJ��1^|h�vl�1:����v��n�5�L#���#�Ed�gN]�]�H�=�s0���^�bZpqe;�5��后T-˾��0U׸n����~s�l�@�(`�4�O9�n8�*{]2S�~�K�p?dꅖ=Ww�N�'s���c�sE����6�F�8�J�uRHx�$ݽ��"��[N􃩝i��OM��ޔ��ek{ɤ�Q���ӭ�����(��7P��!���ͤ�� X�;<���.��y��*rI���=��\I�5v�9zup�Ie��{C��Ҿ�κ���%��i�d����Y��-�YK[��~;���"�(&�ZYg%_$yo�w@�Q7xk��;c�3�
z�i��5�*ϛ5}v����^Q�Y��!�4W�u��t(Q���$�-�1�k_^����;��Y�B��J�`*��^7Z��B��,wRެ��Ψ,r��2e�2S��G��]��rm6��z����#��o+gT[L��6:�͇Nl�Œ��:\����S��ڬ�~��ym0T�SG(ǂ��"�2�z73�Ux�!s�U��B�;7�g�U�w3,ta"��d�N�=eryp���N�r�Aǥ"-��7L�ݹ)H� �����k���m�T�/)E��>��v�c/tz1�	��-�Q	��w�.�l�G6��j�C�i��0�֨b��G����s��ϡ�L��Ϙ��q?Dl��2{|d<C�m�v�y�q!�C�!�"��`v�I6�_RCǝ�6Ȱ3�	Ĝc�p߭��ы�v�u���%��Q=;S�Wg�ZT%Ձz�m�5��GqUU�2w�)�%�AO�8��S�1q�ۭű�V9ǒ�:��Œ�Oo���9�⒯��H�U����6�H}���d;v�8�z�;N�)��L�L:�Hz��N�'h��$RO]}�~�ϻ�������k�Cā���I��:�q0��>��I��|���	�	�!�ԛ`�`x��I�l*�N���y�W��{�b��z�=�|����q���a��C���x�R�d�2s�	�4��CӔ��'y�x}���������N�Hd��H[�Ci���O>`wݛd>C�z�m��$8��N��'��i8����y��־����$�C�s$���zȲj�&�v�ZI�5�C�� ��O��0:�6�>OP8�=��$6��?=p�}z>�_.�R9�����#�b O��{f&�]�=dXO�]�t�j�m����C�(i����&�����(�>O~�nˮ{�޺��6̓�+�r��6��u�@���M���͡k���O_:�&���טl����Y��>������ T6��z�z¥a��d8��	�"�ܲd�
�}�=a�����z�Xq���o]߶js������}!�B�d�!ğ�ćE'��O�&�����Hb�:��zɷ����}c���Rλ@�L?����b2r}Ƭ8�3\�Bk�t��$��b�RE'�ߔ ��dYX�m��`v��s�z����:����������Ӫ={�H�yE/�S���'1�Bc�# �v����һ,B��Sh�(kh��^z��S�K��3pq��3.	X�YW���}����R?7�}^��z��C�:gl��:a��6���d6ɮ��;I��hC���Vf�8�=�������o�{�Ƙ$����8���%`tr�C�x�t���0��N�h�Y$3��`m��&��1�W��>�gJ<��w�3��#& }퇬6�h7N�2q�̝2C�Y�!X`x��l�!�dz�f=�W�ǽ��{鈈ںLm����^}�~�N�8ȧ����43���>g��O�9d>C�zã��<d����Hg,<CICY@1&yOY'�4s��}��ӟw����ۿ~���E��N�8��C����x�>a�;g���v�����S&��C����1����Wm�惏EO��#�P���aߢ�<zd�uC�m�|�q!���06��'H|�����ԓ�8��L{�>��F��e����_�t�z>��I<`v �u5�$�Y̑@8�6�w�X�|�wHm��kw�ԓl�O���7�ooo5�{~�=�>$���@�=��Y{g�=I5h@�G���^a8�6�,�0�|�>I�x�$=a3��_r�]����������@��&��!��Y.�z�>C_S�!����N�h2h��m���	���,���<`o�;w�{��w�}��:�~��OC�q���r�Ԇ�>5d1��kvC��C�q�;:�@RL���&����x�XM�?���������ѽ�
8�[���g�]�;;���V�{Z�q�?HoUD�^o�'ebl�C{��i]۾���⸅,�z�8.�9.;����fS�7��e9�{9r[�e�7Q1��s�9���A��0ClЁē�,1 k,6�l��ް��42�OXa�6Ȥ�j�#�����]�n-��/�S�d�!�Dy2��+;d>C�(N2y~d�!Y���Շ�0:��q'�2��Ь�C��=�~6wǾ���|;I�IϏ��8���T�+5�	�C�N$6���`|�)׾a8�1!PP6ȡ��z�������^��]Y"����$��:g��j��hc4u�j�$8���&07�$Rq;�sϝo������;dYr���!�d���l'̋6��'������;C>�By�:d\�D\e{�1�>�C�cP!*ՙ����B�۰Ē����d;Bz��`,Xm=BT��v�'hs�TuyO�혌�z�F�-�u��b�Z��u�ޡ�!�O�N�|��v����ā���N0��:`zÉ�;��>C�G��	Xr��!YP�!��~^���hC�@�$���O��x�Ԃ�Н q5� t��z�o���|�n�n2v�qߓ������������}�}��>
ä�3�ɝ��I�N�@�$�l���XN�8��208�{CoM��>�Bk�{���l��G�pc��c5\�]�*ߣ�S{�Bt�״6�L"��&�:<�C[�,��Y=dXI6�h|�v���U�U�
����sҎV~e����%�?\���ǃU+6��N��
SG��a�i��5�����{ʘ�yף@�q7Ϧ��7[��r\Rm��Z�z5�ʍ�ڪ��M''��!�c��V��C���5�2d��I�!�ϒx��J��0</Y$�^��IĜHt���6�'~tr��z�^>g���Ԛ���Cn�)'�i����dݘ��S�6�ēV��I,И���E�B#Чۻ��ų�]���GH|`q$�3����f�w��!�Y6����a��N3�������"��I3~޳���ջ��������8��\�W�i$��8��N��}������i<a��ЛCl���@��dXM��~o�&���ߞ}�;���E���0�5l'��y&ЛC��C�z��ā�z��$���aĜ`q1	ěa�݇|����|�>������{����`t�����L<N��Ha��W��htw�|���I�3(d�0�Hu�y�3�y�w�}�Ϻ��):I�6��S'�5�=Bju�<I��N�RN�Vk�ԇ[�Y�ӻO���d����dOd��>�����s�{fg��1��ԇ̋$>@�� �"�$��	��x��2C�쐦��2a�qw�k���~� ,=`}�xIRz�$� �,�d=Ad�"é��@�x�8ɖ��x��!�4�I1���=�wq�u�>�w�0�����$�ι��N3=��}a�E����N$�d�&�&Ї>��b=���Vd��6o�\uE��w�p�w��N}u�cmk'�tx{3��(շn��^{p��I��}�u2�i����X_�/�S�!���{+4�U]�������{׭��z����!�N��z�a<���L&�$����'HO=�Ē�m y�;`x�r�ѿTz!LF��0�o������f#�b$�0'L;d�d�f@�I������^XM�)��M q5� t��8�ov�w�f��y�s�xbCI4��5�l�i-�J1Pf~Q��5M�|�t��������H��k%X�$E�}�o�UĆ�����Z�Њ��jE�u�^8�����Ҩ�Y)�o;^��F��"vMO0��Ul�(��[곔�&�Z:�-��{���j:g����c�L.�g�kf�)���³���>��x��xr/�Ŵ��p��w�Y�Ux�QpD�j,�9d>8��<F����١��5yu���dN��E�v�P@�N������Z�U�W.h��
�/J����P���ӄ�E���^��×d�ԭ� D"��ވ�"1�����Uחm! ��t�|QƇ��Tx���}���}�CR�cuUf���D����GQs�"cϪ�:��U̯:����tE���һmrE��!v�4
�%��;K��)OF��>����q�MX��N��[w#���|�V�Y�Ϥ���+��_*��G�J�Wg�"����TW^=5`_P}խ���|�i�����/ϓ�O8�D2�ddUd,7	�`�ټ\ֲ[�B�����nQvq��3ZKr߫�_�}W���)^k�Y�ր�Z��ɺ�� ��-=g*۪S�\�%�����rS��0r�E	Ûѽ����\���~��P^�'��^8oq��\�%9�ee��7:�~����_c���^܌��P���e��[�E����x��Eߙ#ܸI��H�iz�OY黗Ĕ�~��������W�C5	t��=Z~��z�A�x��h�b�:��o�Ƥa ѳt736'�&�Q�gƲ��/?�X�u��{�㎕��<�Wk�{"�J��N�Q����E�Y��r4&�0�;�UF#Т��wP!v�J�N�=Ϳ�-��Pw�s$�&^v�@��0�seI�}xr:�5Uo.���"��Z���q�(�&Y�W�q��_.�.������T��E�Qzh���;����ۺ�s�j�Yƍ�BG�7���#�E��~�����N����k޼ec ^�}��D�������<�r۱�̫}P�FG(�B֚2�d���;�����ۦ"�z�z5�Vj��͡K��#��r<�ɛ�$�P��������[+R7���7Q�F�ةH�K�w�1�8�vD�Ա���ò:�P跆��˵y�P@�u�G��X�X���M�
��u�zJ���Z��H�/��䯶�Etc;����)Wy�(��[��"S�w�y<��ќt��8U9��*�R�����t���s�\��WN����ͫ���!ȋ%�A��R�]��i��� �+�]����l�tǯ*�e��X؅�u��`ͥc&7p2�ԅ;�:}u��W2�6�tw�@+H�ƥ&rv�۳$��4������Ԥ����X���3	����
t3�t�KFnQU�_��t� �<���}Q/�(cJN��ѹ�dB���];b�d��\�L�)���qSg�B�)˖-fZ��++	��Q� �ܖ$�HL��a��*�,c�TlY%B83.5F�pJT$twN�K��Q�pX�^R�%24%���a�����i�e��J��wm@K�0%L@F�#b�ۡ*5g,1�D]�YN/�U����fÉ��U���k 4]���w�Y�s"�����pd�_��ZMXqˠ.���2ʁф�$��,)I�
E�C2��*1AP��B��2I%�f�2��n*i/�
mZ��``�\�IԆ	f�JU�������dF�ӹv�X(���tnLnE��Pf`$fMXM�	�Z�E��9�7��2��)5Ȥ�u��:	�����S���ǚc��J�i��޼߉�{s<�}�N��O��@b2 �d��Pb1c�J2|��,�F5���QE�
�h�+-���l��H��QC
�$0�
镐X
`�J�6�T����+"������a�J���jGY�Ā���$�d"Ȣ�T"��d��& VD`�)H"�X
,E��,�QT!��r�(B�
 ���}3��z�����&P��_�ر�$ұba�
�V{���;&c�gY�����f�R����{wWsm����O}�TuTrO�Q�����m��6��}8_s<� ��xS��dm�.)+��ŵjU���A&��,���K>�UX]���*/��pV���b3B��I�#�����D-�D4��W8|z����o��U�� �߁���3�w�X)��h��õ=��������p��i%��j�58�h��ګ���zK�=��p�4�1�Fx ��^�V�����R���4$R����[���֭O'����RI�(2�^��}���'c�ׯ��k�7�i�u;��;*���w*'7ܺ�")5�r��� 6���;�H�ޮ�n#YX��pT�}u=ݽaK��r9t��s:s�u�7k:ZH�j�׫1�s��+�=��=1Ž1��s�7v�?)���ک�]L/G�J�}|_�ʔ���mF2�R�էt�Wys�ɂ��i$��Q.:;1�)�*s���n's0�l�����ϡk1J'�T�Q�R�F��dR�лmZ�O$�v{.��3]SQƴS�t��I�/L����k#���6�6�Q�Y��#����1^f�u.�n�7���t�-.,ێV;X���!������p:C�$���;O�Q�x�[���v�.�B)��y���o6��<G=o�����k� �~a{���o��R�����ɳ�^j�*�M>IՀ�s�=�s��m��=��ZU�]&{��x�P�Ҥ�*��+���O�R���z=����3�0{?^����	%Y皛ޤ��.��	o�e������̶�a�Bq�WZ߾����~�ɽ䎅�F��U��v�s�f(���gh��m���~���sfd�ۉcs�܍R�u
�mI֙W�Zɿ�\<�ͼ��.v�kk�) _�I���&xD� MU<D.8/p��<[�sR��/r*��rUt|2�q��̖eE-Pwe�m����#�S16��m�qݫ��]03�TNC�ň����_f��K�|T�%5�n��Ň��n���U��D��i+�)@�ٸ�U/���ʡ�v��r�N��y�5�P��`��':nc=�j:idܦ̝�*�}X���%ӂ�<�)��ې`g�_��G�����IV���j�h#�v��qP��懱�Z�h{�4(�Ǿ���w��8��HN[W����G��*���+�:�Kfx�̍�ټ�e��ц�fա�Xzy��NPlZ�p�f�dK���	m�]@�����*�i�z(m���A��d���[仼�����[��ʪ���<����k�}՝V=:�wI+'�б�x��29��UǇ�#���X�|k8ci�\�-61�ߩ��ْMgA�b��OP䵴�͇��m���5���wgwm��	ח`��OX�1o��6�Bk�-�$�ӫ5L���]�ǭIѤ-���G����^
���,dn��6ۮ�w��&EL�2t�')j:J�����Dw^4�_Ue2:�o�+o�+�F��d���փrNB~���2m�l��C\����@/I��"�)�Y�SQ.~d�6s'z$���藕IZL}�*��0`��Bƽ;��y��~B�Rd+#���ilz�Q�`������k��z�>z:+n�ܤU�=��\l�{�y�|�hEU�3�=�J��� ���<�	P���w�i�[�)V���m��0��@� ag�C�p��85�HW�H��D��\��&,�O�ېt�0��<���Ţh�{-�v��9�'&�v�'�VUY�ni�[GHա�`��*��*$�.��f$*�J�D��*��k��ټ��8���ޏD{��E62��$+Rg���Q)d�T��=��E]��ѝ�=�q ��^xs�vխ����Kػeƅr����vH��CW�X]�wRt��K˱����g��;kw�e��a
)^^e��*A�9��Sk��y>(f�%�X�"*��Yɤ�5l8&i.1l�N��+��Q��3��V% �z�w��+k3�{5Q�a�����F�^��`E�:��`x����N���w�G1�&
��Q�[<�����Oy���7��)���	#���B��l��^�]t�h��WT�>r�y0'	.�ͣ.��ۢ�Kci��n�4�r�o[��,+��gc��M�Z���x���2p7�&�n��90j&I���U�{���{o�Q�L���~<ܸ�e�i��/���k��\o���7�pyQW�j�����g�T>�W�#Jo{��t��YtE�@��VM8�J2���VkB8�<v��g��ظ�-\��8��$X���W�֦<��21���)�%?gܒ�v���X��yy�`��2�S���:Y���W��Vv�(hQ��M-c��GԢ}������{\*)��H���÷.�4�U�	��5����F+q���Y��nw����'�$��nE�2&��(�]tZg��(����ԎR��3�&y^o�����9ʦ�廚l�{f9c�r7�2.!A;xӊrʵ��vVӗ�*�Ri�[�}�v�e��LM޷$�Gv���d�ټ��)klZ[]$̗��ROʈ���#{S)�{���"͞���lx�C���C*�u���q�8�E�ᆲOB�+[��3e���!���ԋ�K���hU2]\;���������K��!����C�z�'=������G��B٨;3uʺ��OzZ&�0kԘ΅9��:�3.�M��+���Vsf���z��k�;i۲�y����k^�*��խg-��qx5���m����sdb�z�ᬍ�sS(tfm����{�k�4���^��Z�YM}����K�0���i�)��6�.*͸���f����Ѩ:ǚ4��	�/�c��|c;x��[��}��U��k�l�ߡ�w�:��մ��3�������̾U+��S�J�x�j��k�Ж�]��H��%��ֵ_,�@޶�j�j��a��w�W��,��Ð�d�KG]�b\��l���32�(��DϺ��H+��%m9繺�;�1�Ɍ;�vH��V�rm�_�}�)�r�8�R�gzn��'�FkKj���BU��Hr�n�Amt���y�n\��Ou�W��ɨ2���Τ6|�K�q�y�x�6Q]���/�"l_Z�V4���(i���xY:��v�1��㺞,��ػ��:�8�d*�h;٤aȊĊ��Kw�ndzM�j�;7�;�N��%͇Z�n��\]�Z��cgl�x�O#�����K�{ވ�<q�L���G���2lP�>5���S5�N�%G8�=�m6�)Ld���Գ��.D�MNz���.cE�̌�eV=h�֧�l�i�����|t`�kx؄�r��җ��Ym�P��NȞ���P��q`���4"�U]9�t�1�<?�㻿%�~�M��*_S���e�w
S�/�BDeC}k�j(��.-�R�k�dF�y>�A�e��{Gj�W�6nS��E�U�n�g�,T�إ��TK�����Kj�C<�������eN�?
�W.�����������U��z�7~��ޛW�T�᠊��scEV���T\�^��<
G��SdOd8u*�����p�OS"�ɑ��)��t�G�jb�����μŮ�.ðv�>�JU:�����ZFQX,��9��i�jow�)l2#W�
��}�Kҏ'CIU\֜�(��O��j�9f���%a�ƫn�`�
��R!���6�IP1Q�+4]f
��Z�sǬ����P:Գ#�=�6h�ǂ�e.�WJ�k���7���(m���q����qP��/��z��z�|1��:��rS��C{�'dض{�;�J=4�,;�ȕJ�8��ǵE������J��YӴ��\(�>|˝]]X(M��X|�:�-e]�w�r�"78�����h�%�<K��Ŭ3�s��E����pW�	ܮ7z����쬚�5�VqS�ق���ϑޤ�go.�=t9��V��8k��k����Zq��d%�k9����[Zu�C�I�x�Dyi���
�`�a1���W%�ʓMu�#���Z���n�i�Ɩ,A����V�nND�g#S���i�X���;�y�5`�ul��!������������&pR��"��=L��{��2�mF+n�&�ɂ�iڸ��>2}ĘLc�U��V,WJ���a����qAvY�&�2Z-��˂�X��̖�U�ܰ0�2Lo/��� ��@:��x�e*�VZ4��1�����0	��Æ�bc�a$�|- �}�yX`4�6���X���t�t��ͰM�Ɛ9��I��˂���V\@�R���e�r��Cn�?�C`�s.����AR�H� �,48���Xi!��3�A�4.�1�w�	�̕H����Z�`�4�`��٧�,o��m�?"��eN�2h6�|2��-��u-�Gv�9�.k�xr�럕��8PUE 헔�d̠�
�P1&0�� R*�"ɉ	X�,����
Ì�XE��,	���R,$

H)+$
Ȥ�"�+ ����,��R�B�,� �QVCI
�AH����ȠEQH�`,"�,UPU�RAb�#$X)"�a��f�� 
�@�T��{����.k�����Rc^�¿\jc�۹�iC$�GF�[���l��Tݜ�S�DDxަ�V?��T!ᡓWZ@�5T���= *��*q��R@���V�υГ1^tۉ�+��ڀ�4=�
�<:�F�&��.��Ef�Ud�U��F��i�<8K(`���4@�ڗyܛ�d�J�ט�#޿?��9Ri|�>:C�kͫ�<R��	�G���;�(�+X3�� .n�A���'�¦);}ɭ�c�H�����xp�M�n��0 �lp;'�.�1<o�:
�t�%_�.��gh�"���3���0i��ќ�ዑ=)��. \�UN���*�`�G��^�T8f7�6xC&�.^���������\K�0,�/iKZ:}��*{�L�ǥ�<iHdC�t����U�W�D�#A��g�|�y;�w|U�3BŻ@{{:�t����\E�%cV-�E���P�͡�3"����Fb��Y�'�H-VVu��5ûA֟jfe[��1��`S�hs�2-L7���W���w%���ة�.j��h'�%�z"=�c7��ݶ�Y���˛����X�3l�	uQ{Pg"����%�tRTk'����Bm�ˇ3T 7OաB�[��O���֎��X���1����gG\��	�9}���-W��Ӂ�6.�x/�s ��i�`��6�w,��/�E���Z28�J���p+�P���x`R��z��xW���)��g��t;v�*�v*b���I�|�����@��D���ot}��=YG�Z@����Z:��3V��U֥\C~�s��E�
��q����2:���S&BB�zV*�v/����u��CeO{�L��}���`�2���~UMW[#�;�}S]����)ԙ��W�^Ӟ���f�sP34�����J����) J#�p�b�y.{�y!���+��j�6��BC���EdvW���^��}��ܡ?xP�4��W[��]U�>���n���i		A��0g��}U��xR��.�S�Ʋ�7�]$���ɾV����L�eY�.zkV��ܪ
�DԖ��ڴ��|
���ؗ=UU�ϲ[�Z��U
Xl�3�]9~��:�6�d�	z�KD\�,f���C�7�&�ATš׹R�V,ap��$�O���x/m��]#��;Z���9,9٩�5�U�tɡ3����o��E�	�k��kF�]Hוb��4V��F9�cu�J�Эo(�j�`Rq`-Pg�[4!��\lP�_N��\ܢ�t�U� ��
�V��r��c��;�n�tp�y�(x�ڭ���@V�F�ؚpcKDNz|��1���v�>�B��g_�l�D9gd�\�Ϸ�M��LΗ���G_jj��)�/�����b��[]$Twx��֤��!����'�Q'�EH�0iK�Dx�4��T��Q�1�fg�ݟeKS*]�71��źR@k��}6�׌�����+&�>��j�|�J���D�Aڄ����V�\�F��X���r�}q�{��+RnW�Έ�d��o��dC�*���x�c�e�07�*��i��\�ꮗ
��.[����u��AP�J碝{P
Z����O_��[�:�Tâ�n���>�g*��� �37���Ln	M�ɽV��/�t���K;f�k�FF�@�-儻:���xS���`@�SB�i��P��T�U��2��c�p�G�����*���@�0�T�(O�Et���).��ԩS���K��(�I�;3.)����)��K�T���r��t�ͧ9We���H,\���_(�����w0���<t��77I�Rڛ����J�o9.���0��B�F�g:Tuv��1�S)�b%��ӟ�W�_^�}����q�P�C�� a��J�i��j�Y�������Dh�j��^UʏP�� hY���[�ܝԯe�x��۩��3��ªS��H��U=8����Q��g3�� Zm�F\�s��u���[*�>� h֍
��q�ZM3Nh�e����
pV*��R�jp��Vʔ�ɩ�&n�OE�Җ���Cf ��X�����Pvk�t����+��]\S�6ޢ;�_�Jx�A�b��8X#g�׍j;u�u>���t�5VOY�W*�:��^O�9Ι?��*�X���Je㼓�^�h)�u�y��|G���P�H�<�{�X�^�k&���+U���>�����c��j������s =���� ��+�y�H�*���X��~v
њ�<�.��]�v)���37�S/�e\�&qL�7���tt|�ԗԫp[�7�E9m�i!BW��;k�s�o��8�\6��%ml���}K�$� �c��E�Gk�(���G���|U�#�b;�D��9�N���2_h���-S���Q]۶<���a�Er�r�.����W/�=OX��0�Gvr���$R< ��قс�bR�^'�
����<=y�+|��F��F#���h�e��J�QL��&̵B�.i��MY�쮝�
�ưh~�]�hY4ժ��^D_Y�Yo�ˆ)�U��}1�̉�;�cG������s�߱���yP4pR�C�W���S����5���Fd�c���8'�Xvk�}|���F�5��FV7�~�Yh�+n����R?��P!�׬�ߜc�j��I�ܥ����0O�v*��OU1���>F�T�f'l-�;����e��,4he*0i�x=�+�Ѣ��씖�{�\,�;��[�sM��G�"F0iT��
�d����3�^@�Z+���;-6jߗ
{�+,Kϗ��G�6�#�ja�À;�^�x ����W�~���^�U�áW|j��j�;�U��5(Dpa��ؽ�0`B
6tz��v�m	B�[���/Mu�倜F߻��uz��p��(*��:�� &~��c�k���e�}4�l�vvT�� �A(\�B`U;��]N�՚鵣%�O������G�[��л���xב�U�+��H�q����v�i��I=�ᐥ戎�X/ǆ�����Ŝ�
����K��V��2|�¸R�*sWY�;^��]~" Rև�U8��3y˙���=@��ǃG����x�{�����iZ+n�!�����S`��� nԼt��R�%é#��@v^�y6�y���%�;3-��MZ��nL���`1{�����0S�l���]��;5���=��d��&>(L�æ.*�v�57���\����ïpR;E���P���%n�`RB��*���)â�j��1B�,�y�~e��{�� c�x�íK�o�XZ�]����\��x뾼�2!��
���*Xt�"����6L��@p�v�u줒�R�hH�Z��fw�e�t�Bɮ�Z���n�U�RI�����75/�Y1�ǘ�n$!3�*o�+d=���j�i��b6Ί�����X��X�0v�SO����Ǎ#h(�����}�{2�.�*��dؔ�o�J����Gݔ���4){N}���551�1~dL�K�;1v͋m'�J\:�s6�a��Y�5��*a�D�W��5��~U���9	�S�
�olY�wbf��s(�����n��<�������נ���gN���F7�U����ќ�[nT���	n�#$�����yf��U0���2�g��,F�fֲn�j���̖;�<i��3���-�i퉃,8&У;�9�aq�8��Q������+��9ܣ30%p5>�!�y�=���w
S�&�}&�uT�Kt��.7D;���]3"(�� B�0t�:��^nV��$U������7*T���J��[���X�@�vxU׍;#yDT%��3$��=w�l�S"`zL�!��V��
T4N��y���c:�q��7�<>��W�*�Z5��)�^"��o[�S�:�]\C�f�:uVG�,V�\��#�BF��+(F:m�Y*�
��`9�Y�*I;s70&0�kBuI��j�KVw�n��谍�|���y`�(J��5��b���*4v����&oP�C<�&���=R��Ʊ�5�q)�Ӎ:��+*.�h�هU9Q�n梀��v�щ�CD���ge0��J�mev"J�����e[ؘ��j�ܩ
�k��U���ଡ�ȸe�ا��E,ڎ����΋�%5-�\tOmB.��!���<���NWJ�2�;��¹��V:�υh��L2���V-mNB�5�%�DŚ���>W����������zһ�����H8�o���bDeB�1��Uƶ8�$"��ҝq�˛���F�1���KT&v����&��]Qү�[��Aث��>�S���02l5Ç
旅,���ȖEI�0���&�B�#�*�b��&�գF��G�鷻6���0u��pѶP�B�=��w.�ɋ�v�Sv�<_l)l��R�x1�]�=�5�p�j�,@�{�5�
��e�u3�n�oS Svn���N.�2��9�iù�&ٝ(��L��7]dc.$7���mR\��f�K������sq�y�Z��~�p;�9�0É�0ED����DX�v�n�E�Że*S����M�!��LW�33�I�i�Ẻ�K������*`;H"6���v��7��\����9�Y7[�ׁ�P�o��:a,T6���֙�R,a,�a�=[s��"��Sa�3n'�u�X0�#�8�w���%�����=����nV0���\�)\�sz.VVd�B��Z:�'[���	Q�2���R�Aō+;';��](��������z�����&�
�}���2��F�Fp�$����E�g�g��=�(�~��5nB�T��7{�;��4��vGhV��J9�6h3a
��v�䷺Fѡ2����i��Zdv�G��Y3{X�SX��=Qx�|�ŗ[�L7s�5��l{�@��w[}��5�h���,�˹�庱'�sI���^Ly��v�]p����F�G��ۛ�:��:����1;�e�<�]y�I��o�;3[g��:�ϪN���t宍�o���5(2(*�av�靌�i��r��9�ʺxw="�R�Gf�mnwVp&�%ܲ���6Z�㽩R>�R��Z��C
�j�p��NӋ���ir+'9�]���zrK�<9{����"��%h+o�����^�6����"m+��6�tʎ�w�+.XΥ�!�N�ڼ�Y�I�$�ŷ�1R'.�^ٲKujJ�$�A�=�h��q�a�O�G�n�pڵ���)l�(��H��{"{؛E�b��U�C��͋z,>��Y�e�:c޺�!bE#N-�k��#�C����*l5�m�X*<1i��]�va�{��M~�+�>��
�"��%a"��AH�R*őH()��PY"��Y P��Ʊd�CT�R�XJȠ(H�!�XcL%d�ɤ*ām	P"�`bC�aXE
��L���R*�,��"�i�3�VT2�i*i%LLd1X*V²J�U���Ȍ���"�L1��$\`T�m!q�T)&!���wηώ%�z����(��c�٩m��6�?nR.�
{x%����1������?)�ɿ~´<,�ub��[~Q�^Ud���y��fO~�gz�=Ɗ0`��@�xh|-U՚�6�%[B�=ETi�����-�!��I4�ظxV-���+�����w_W��!,����Mj�]C;X�ii����	��i=�%T�my*��3S:8٘F��G4\]F��	GBb���f�*�wQj��X�#�jf.)�w"����;�+������G.20h��^��V)�1�&b�P3gI�"/i���`���Kz4�`}k��C6�p��^�V+�C�Q���&�Շ��.'�w(MML��0n���W�l��1s���kh�{���sұ�Q���0"��Y�T� 49�O�u��ܠi�?e)�t[x"���<��'��6�YDCr��*�.�:�t۹w���U�⅀NȦ�
�򎜾� �r�B��
����f+n@5�����`�~���tF\�dw�N|8{�
��ׄW�|��
���S7��
�8=\:�V8�ex�k�X�ӳ~�6EGU�/R,����I�ֆ�Sz�d�P|�q�@[ţ��PB~x���o9uP
>�8+x�M`����
W���<x�<�����іk�1 �� ��kv�4W3��/�p훘j�������Y?
3X�;���Ղ���W�4����0�Xܜ�����ƅ�4:�.�tq�{��n$)�^�>�cstQ���Y>n�WmD�T)aU�@�^Z)Q�@^�ZpeZݶ��e��f�`炣75&bU�Pff�(��x�'�qR�7�.-��ǎeM��j��&���
T�*l�L�^�Z�"4���	��[C���#΋{sq5�.a�����V��:ۑDȼ�a9I���W`��BVrT��4��[{ȯ�G�o[]D��_�jY�j�6%F�Y�E���B1�Eƾ��/;6\H��<f֊�uCE=Tɱ�𬳠3��i���wkB�T^��9�JK�����Ȑ'	�7��PZ���|^ٙY�K�5�M��O��]/g�����a��i/9x~��V��c����k�Գ�ks�FF�Υ�.7a�}�y�O&æjǶ�Z�g�W�W�f����z5���������U�]t�T\��:lW�0�<���]�yD�l��j��έq�0�h��C��x� ��h־hV�8<���r��TԻ�w��f	�p ��
�jdZ+p�dض�xV�V����J,�#L`�ԧg�O����Pw������οz��,ku&�(�׌��ȟ%���fg���d/U(��t�0�^��@]��gEI;��%�B%JY}�ѝ(�������kX��3²��W���m����7Ӱ�b�*+Ex�uVi#��\�)G���=��v�Y�j�T�`�9VU��~4���=<�֍��ۊR��WMX1��"�Sʵ�*؈�Zh����{�x�{���h�Y��+�ɔN
�W�0��y��
���N����rL�j�f�S�5)�Ue�.�O.�啖�������\!�������� ��@�{����B:`�{�P�U�ώ0��ʡ/�ܩL(X�cekc�����"k[i:�t����	B����p�,K��F�X�K*F+����We	px\�T\���1cNLߦצ.taY_-0��W�]���熫��*�pp!�K���oʩ��=��]>�=�
;^�R^`q�%��lV� ?_l������7��Dt�у�#O��HI��u��fEd��Cruq@1�m7ZP(��h�I��Փ��A�	�~}�y�=�Nױ-�6�0j������2o�[ !ҕ1��ݓ���g�Z�Rz�r��?{}1qB���NU˕`��¢q�&�p����l��Y��)�����K�(И�t�Q�*3��qP=Qr�'qp)�U��A�5'!�*� {�٪R�w��@�~��4TP]������E;4l�T�_-����TGZX6~��0_��B��;W����*��ɸ�ƃ����)V=B���e$�w.+���]���N�P��]	���O��6�F�pR���x֮UՇ��йi�T���壠�-��𲊼�.b�ɓ��jd�2<"D��3єh�/dV����I��<Â\�OkƸ	�j�:��S6�L�����+�q��o�|�&{{.g�z�G�/���
[����uv���@\S�6�j�p�����R,�LY�ٱ�V�"��XO �{��Q9y�$�WԹD�'�7�t2ֻ7+*�5��祓F�h{�`�ds�,���u����
��*���P�X�:��8�ջ����Tтͤ;~$&3��\j��T�����B"�Â���1�H��ʐi�x^Fi��<S
L�K�:cS�KD�B�'���I�.��:r��t�NT���:�"��h�������㜌9�޽i���fhVg;�*�����n���UZ�t{��^ivW�̫ޠ�� >gy�^�N�zs݊`FW�֪��'��c[�,<cl�@(p�a������o뷣��쥾n^����M>�+o%F�R��Z�1�W!EGM�9;ꅜ"�C����p�ϯ`�n&:+CF��g�X��t��4�t{r`��](�9�YC�7�S/���-˗k�{�L��j-�Kݢ�'%潭�{cc%iv���}J��ہt�Lˑ�ܘ����Y�1r3�J%}ۥ�cC�p꘹٤}<8,���|UJ+x��B���o�y���6�+���N>.����s��aj�V��}�4����<�ʺb���~���7M7Ƭh �a�:��Dv����vܬ<�p�e��^Z,�T���y5��K�ca�����������K>��VF�Y��<;�=I,�"Lܲ��,]u.b6&�"��oB�18�����GT˦(���xp�^Pzχ�ۭ�}���I v�n{�\�jK\�X�T�sp�{G[�9������!�Ȫ��?h���xk�[���^p��[���W;���9�gf�әQ���yL_�l�0�\qJ�u��Ϛ�)�eѸ&�]�z
_ W�wuܔ<E�`� P��vOs��Z�@����#&�Mf�D����j*3�*����^iJ��ڀe<�G6F[��s����֣�]j��m��
�1,���G����t`2�U���ȹV�L��+���NeClt�*��.zb�)�|K�*��0Nq<��'�϶տa����u��rϛ;v���=x��/3��-� d��.��x���E�+Ç��a�)���i���J6���ۜ��V�b�32Z�r��<�Wc�)���"�+�L�T�<��N��s΀�`�ᣀ�W��:�,�$d�Ԩ���
a�z�sKT��'�@�5P�֚��s=��c��!V����a�ɔ0R�-P��xm__9ŋ��ʆ�[&\�A��Rb|f,DS�,O[S�����쫣,�U5pDEF�MBA�^��
�d��C�U{�.�����.�J��;VU�6��(���V{f�Lh��W�`o{ճ�v��lH�J0 4U�b�h�ԁ�WNRj�!Ju�o�řP���� �U6s;���i��ڭ'��%��Xg�|�R7��G\�=�dY���,�mT����`L�R��
�E��*�A�<8|�:�W��+�X�(i4���s�c��?pB��K2��x�g�)o���]t2��}^��KP��	ƪ<[��>�^,=^�70g6��
���7����r@�V>gb���q[~��G�a��<;�x�=+5�^"���Z��
�a���7tۣQ��+���ژc�4��O3c�Y9���پ��@
�9��T��J�z�Y���L�aJ/e
xe��w�W��5��W��gʃ�u�G��F����D��,��gl���Z=Z��(�0X��A^U�
__+�^Qq�������zL��<2le.U6$<N�)�+��U�3x�˜��r��9C�Y��E>�r�R�tUE���X�/^%(���d./���\[̌�&�纡NģUUiJꎝ��"�O����2Z��V��}�[%��Un��MM�V��3Z:mk��ê�g�y�J}3������&G�W�UO3�eLdT_ǫ�Mr�*�aM/��&_��lV U�*�Å�FC���śʝ<:}yJn^X��GNL-b-e]ј�>�:7�D�?<F�|���]�P;J ��-Vx(sHu�\~���B�Vv��vLX�\uB��@u�U�Pt���C���f/{{z��[&˵7������)�h\�t&����Oo*TY��US7(h�.`�X�8:���{Xp�N��A�d������T�Q����T�p�/#DGf��*x��B#=��#�*��vS��w�p����ϰ��4�G�o�`���܇77��`�C��9Z�l�7\A�/y���eB+V��(��aK��l���W�ĵ'���̽�snH��(sPZ��Fʎ��{D*ۓ
wRޮ/*:�"n�6�	���r�~��8�C&�әmPT���Ʊ%S�{�[��$�4�WKXES|�*1���+YD�ɴ��,6m�aϵ���Y��Ei��47"�� ���&�l��%�s�������pۜ=�y��k�����@�,vVi@��-��y�9�j�hyVl����R�TW}��5o�t����]`Y*�Tp֗}��T�G�d��kΓ�<L�"�WFҀ�o&a�*�y}�i�qq�8Livv���0G���t��[��D�pq Ѓ�s��E,:^�,�h ��O+�ޖ)j/u�ʔ!��6��`��ч0
7|j)5@	��W��|2Z0�����F`04$��X?6����Kn�>Oԫ+3Pj�M�E>��w`"vE]P!�&sj��S0�c��9�&�����DG�A�D��߳��"pa[ƴ$̖�2��2�j�Ia����4U�e���5�ϲ��&�5�ˊ�Ҿ����i�v&�8����������Sآt}/w���<XT�D��T*�`	��汅io5�2��^��Ҩ�i��+����� ^GX���^����b^�̍���q��(��S.ə�:ݫ@����B-?p�����T�0���/F�JF�n�{_G��J�Y�w3���kOp֣�e0�\�x���G�J�r�y�uì�;\5�ݬ�,��C��R�j��gnC�>�� �V��~��X���
^�i��u0#�VVh�`]5S�_��#��v���h̝(��]�v���:{Q�����%��鍥�Q�щ��K�p]��B�jʕqBsYI�q��̀�-mYMnH�X�`N�{.c�S��L`���pK��m�۫%H)SY`�[JȢȰ�VbAd�%��b��+1��1!D"¥@X� J!X��BH����*�`V�`� 6�i�@�h
T*,�`)QdQaY%d4ʂ�B*1d1%E1�
�`(�T*Q`���PRR�Q�
�k ��-��RT�꘎X�,*�%J��XUA�٧1	j��AeAJ�b��Җ_O�s�q�8uf*��:�[���E�:H���#�?PU�P�)���^��eg&�9*z�f&zo�5�Uol�αNژ��TE�o��ͫ�Q�$�AZ�`��|�p��墆
�O��]�\6�c�o-�5��r˿I���K�X,xn�lS�����e;�aAR<+C�j�ʷHY�t�~5�)H�������3�بY��EX��*��ӑ�)�R��
�:��۩�i�@���E:�j���4pѶ�ӡ�x苪�0Ն!��xn(0�W�1Ӭ:���G���ZhqU���@CG�f��}�G��;Ƹ68[3�5�\�<���n��^w3����I`u`t�]���K<)���:�R��ᮢ��T�p�U�Iq}�y�=��\�Cg���"��� X=��ӱl6n�>���2m�V�dH��7.�B  �v��ǯ�J���:��9S��'{�-ҍȖ0�8w�4\m+֞۝|6p��:�rO�Wg�M���d�Vi�X8�<pU��xN:4x9y�w�Dؚ��3�����:`s#8��C���f��!�
�ˑ?��1A�=W���et�O�]0=�"Ǝ7&IZ��Ps���2�
]�q��kn8[��M��%��Ua|Q���i������9n-@�yB��/�T7GjV�G�uQr8��p�a*y��&�X_���oi#fc��x���?c��	�E��E�m�la���Ke�s=�?�\�Xa�a�Jj��
U�� �nM����1������tV�P�|��7�Ԭ�UaD����IŮJr�Mۃ~�:�׷*%ј���*D
����4Wfo2�����ޙmT
��h�������r����T�6���E�!�qͅc�x�ݣ⥮���|q�w��̮C�y�\p��d�c,���Yaδ�5y`��W����e\�۴���.Qn�ܘ:��U���Z�]�.��1��%ؙ@%6��O6n��~��[h�6�~��R�f�:z�S��h��$X�PL��Y4� �$���K5.�|0A�V���`���&7p�����d�����2[<#�Kbf.)
�x��L�T����e��Oze���n�p�]d����vW*��A��XI�ڷ����S���mWM�tˡ+8z�1k��%gX3
wr��e�;0덂�&�*�L�^��@��`�B��m�mH\u�w|�cv�VЗP���u9V:��<*����n0.��-{+���;du����q��\��jV-r�����_a;!��}�eb��W���]Dѫ>��F����Ef�,�?:2�1S�����f!����]ƬU�/�w�N��m�&��&&��h�pȐ���s1q� �\~����y�Y��$R8�N��EI�R�iM22��!X�9Jv|3��J}��h�;�\s
�sX��:�L5F$UF�d^�����^ޯTn�3)�5���o�������
�v]P"/F�m�L�uN�3�-���p�g�֏���HA��,xh|�+��"�㓍�n��j�1�A�0g<蚰{�5�����*�j��ܽN�o��ׇ��'�a�ǝ�i�����mN�b���'�w���a��Ɋ�=�e��D��񙝾6f ������ȫZ�O^Q����\�J|_5(W}����l��=3}�c ����Z��V^O5WVkf�}�O�D�~�<94S�Y�����z*p��Ud�Ɋx�}���W�;�,����F.��� ��;����n{J��b$�}ƬYщ��۳����Fh�\��|��QYj����1%u�=�A���7�z�%�艤�e�"��~|�
�׵W�ύ�A����9��o��	N$5qO�ٙpk�;=�9rg�zz^1��85y6�LL�[ςwT\Q�>���a�T:<�uZ�8=�=��r'�6��欦*󯶭1��suSuhu��5X��<xsŁҐrh��;�&rK���S�S�":�,g����S1q�79o4�j���%N��8�`�+�^e�4t�6`�0�b����C�
n�H�}MTn2!!�"v&:FS��_{O[%3�K�k�b��<+A�Z�`S��a�}af��w�ܝa4l���\ .�����JG�%V �.`��>].˭�s7|渽L�)��N��Y*�ʀ�%!&eј����2B�
3�֪=}Sw�I[�h>��ZU�����ǐOktU��0����7v�*�S7S�ȍ4�v@�� �r��.�'L�E�+����oDt�K���N��3��{�	���T��,^L��]�m�(+��U��ţ�����F3W�,V?/����L��C��;G,���e�9�00J��^5,�5���V<7��s=z��v`�]�O�,_r���[��?,��)O3OKe̗���3�&;*-�4��)6�K�}H�}:�\���u�𵯅M f�Wk��[9+�~�7N�]��F��~����5H�z�C­�C�_,o*U�3i�1͉{��ͻ�f�9�;� MI�ݮT�e&͖JJ�2���3
��U�`y�&��pO��W�q����J677�x�^A�<n:'Nzjnk��c��;㩌r:��ͧX��7[�ř�;���}[@��Ԩ�6��,��u�����&�YN�B�7X��S:a��74p"��^ԡn��Wh[Ջ����|��<X���Zt�k�iDɴ�S���͍TT�C���:y/�=r�J�@�p�b����,p�;�Cø�B�-��#���<wZ���LυM4�5�
�S&K�<P�ʝ�"�n=|ڻؘ}V ��>�e����y>��\8uM�u/s��F���c�}�Ñ��=<�1:���4�j�~9OX�I��;Ÿ=�`#^�ָV��d�h�karr�jait��"�@���Gul��j��R�z�b(Tt��c��:J��&�����칇)T�ډ�0b`rL�J�hS�/;��|����Ÿ�*zjT�`��jԁ�T����[�U�W��-h�Y����<&���`�ȕ������er�#�ȃ�ĥ"F{=>ZtXP֋�pR���
�B�\�������P:hmK��w GQ�B��G��-�y-��0>3&�ﻒ���_f2�9Y?uz�W�D��$�E��T����
sr��7��i�c�{��q��=ʫ�Iz�u���]S9nr�}�Z�%m�?>SU�L��C�T��@��ɩ�6b�K����P�%�7�r�,ї���]Fb�\��.�B�t�BE�=\���lWL���.pps����J�;����18�ҋHГ-!bn�/j��y)�U���n+2iH��%���k�ڢ9|j�{�Vdx�v�d���Eg����#I[��T�t?#��B����(���'����C���t��չ�Af��x`����Mb����+�'����o��0����#"��Nwx��ݦOK����t�F��0渹qp;3�z��N��d�m�M�m�`^�>�W=y�dHf흡�(��1�C�w&���
�u�����n,�q��h�Q5N�Α13����jL�\Rs����Z�w�tQ�舥N}2w����L����GL���v�fcޮp,V+��3�Rk˅gڕ&_��	"�L2Ύ����2�2*D5��떴A��n�W��0�x��>�{ތS�X=�>����d`�Ia	偭
Q���k�)�Q-�!E��Tf:Z�5���
���[�z�,���g�Aә�:=���GR�ɜ���u
��|<�W��R�M�J�G��nS�6���I|��1�f��Μ�\���Ɇ�FMϬTeڹ�	7�y�]T+>�lbQ�靖�����{�ʨٱ|l��C�����a�����uXM����y®�ި���%!�VA��O������|�����nv�r4��޽=���v�O6�zqIit{��T���ӕ₢�l�B��+�;kJ��Nʸ�#�F�Ꝃ	�WZ��o�ҮJڐB�~}腍s�ٽ��|�)�s�54j���M���@At+�N�{k�sݾ�f��>V���0��Z5�k=�
LػZyˑl��wk�j��| �c�� !ʕ(�)>�(
B�^M+�i�^����^�jN�
ug���>/��T�� ����O{�+�M@�3�������*�υ�4P�8��2wi�Z��̵r#P��0�Ml�sEՏ:2#�\�ed�F��ԙ(�����`*��u
�U/�jY�����Uʹ�j�o�1~�(8:��54�Іw*�{�{m>��H�{�J��3�}��n���	VxR�@��:�UǴ�|{�/�ײc�=�����>t:��53��OL.�1r�������im�B��B����sU8��Ӵ��VWj�z����oA<-彉�̐��6�g��.ir�.�L�0F��W국��=L�-���}���x"U4��������3:�%v$��f��^����!� �j�n����Q;[N��W
�Բ忈���/�l�㒙�ZA�U��������J�t+�D�ʘˬʾ*;0r�)�w�f�rȺ����s����Rpܧ/�6�d��Q6��i��L�>�.��.셷������A\2IQ7y�b5�wk#�#��Н(<}��D�T�A�U��e�X���p��`�5m-P�8U�k.����4����&���ͱ���)�˙���¸�Ċ�'��FP��w�
]�_X�b��vbp*���V��y���iTt(U��i�|�;V�R:s�t�|+q�*���$�R�w+�Qz��^�Lg�Y�.U�A�&��X�C�.���.
�r�p'��;Y����_m]p��%N6�b0ݴ�h�(�4�*��ű�1��<� LK�&F���0�h����X��m���]PL�g�UrB���/�EDjIx�Ř��]��8�#��rJ��E��',�L����O�$]c9N��@��k]Ղ�L���V;ڸ�����aL��qR�K����ᬲ��K$�@x-$�+���#c��˫��Ĳ��&|��J�$��1% ���-�t`�\D�J����l�V�E�)���Q�m�"��i [b��ʖ�F�����r�
����J�V���pJB3QV2�f[�)�&�N ��ɍ��)f}e}�`�n��fd� �ժ�c-`�l�ڥ1e�xhZ�*8
����T���wX���F��'-s 6um038��J�9 ���λh�F�����ɳ�2:0\�P�X�-B����X�aY-�EX�b�Ylh"Ҷ�Z���E �,ި�CJɍJ�`V�Ċ�)`")1
������CVJ��D��D�������ָ��iI�I,1�hbQ&2�a�*ŀ��L�(�1`���E�bc1�f\\�T��c��rҮZ�Z�LB�ʭf&R�Y���X(-F2�"�ĸDǦ���H��� ��lC,�0�X�*��T�Aj(�E�eWLZ�ږ��0B��b�0\f+R��ph����qSXC�,5���1��fùmvZ�D\or��L`Zq��m"v���V�r_V�@Fml�&�T,���PU�.F�,�������o��~�ʘ�����V���@+F������
��Ӕ�͚K"ʛ��f��m/�lBt9XUO)R�Z�y�v�4�W�b'C�>���k��g�C(<�ʙ�ΛM0�G�Ԟ�~�a�EX�Q��]ƪ.��П7�eOLʊ"��9]�B��и&�`���a��O�9V��ˬ:)}5Rg>�GϺ?no\��%�ix+:)Wp�5�88,(RGF�����4�9N]�$�.�53\��ח��[�*�Ƭ��+E/%���Q`z[Y�CG-�^u��_5xn5P*v�k����B5��3w�e���Kv1�uخ W�{9p�Ã	��j�>��Oϳ�́����]ư g��8pG���`��8y��K�mYK�F�_Q.�w|�\�:W�x���s�v��֒O����(�������u9V��X�4<z�n��XV�:b��p���<����5���"�uƵj@骲wN��.4c�����̀���^eg�/�_*�D�ܹ
Se�,vE^�yy8��%���u��AI0��Z�^f�uj�x�G��,������g�*����FM���f�=�B;h�Ŝ�s����1�Q���'��Q���7�3�2�C!)��ɤ��㊈I��b�I�x�EU�BTl����ø�}�dԚ����J\��^ҖWY��M�VHUFt��ۤ��
a���F��
A�<~F��l<8=��v�0�F�y1�=7[._p��17U4A���:<�����^̭8�9�C��	5�4@9J��-���9C�^0f|�0�C������XҞ�LXM+��7�F��!N32�F��h�vq�s ����ɛ6R�۫�����M��*��&��?�[��+CFxӳc!�円���D�?eEp��B�I��3Q,SX�c�A>�:�e��w؅���pUx��yZи�<<8V`W�oV=\Z�Kcg��OHȡ"BKe�˧W*�{)̩;����n3:*���(��|�����P�7g���:ʨA{�u��+��\wcn�6�S@�*S�Zԁ�9y�1�[��1c�iB��G�k1�tA�CX2��;ZP�]�={=SV�K�F�`u�`��*���,�AQy`y��;w z�9&	
\ND¨�*4�]C�2aϒ�4&�P�3�,N��MQ�H���� ��|x��X<���g�1O���]��S:��t����6�� �B�yՑ�^Q��#�;x��ѝN���v�L��d�w�,�;U�p�؞��CbޱXT���+3�U[5�^����9�ei)}����l��
���Z���dFJ�/+dʓ(���u�*��9��ҵT��EW�b6bTfE���h�FXʧHV�O'V-r���{2�ؿQzo��*&}l+�����y�J�Uj��%"�?z����HK:+�kE�C�`�;K��C�%֮�x��E�*�X�Ueې�k���Jj����zN���E��]!�ţ'
���Hgg��s"f)�[����I�cFK5�hC�
�Ĩ�����<:�Xuztv.�oC(y��	���f2}�G���A|xhG���g�ƭ�o��&"*�x޻��%�)^;������.�8���@�8����sj����;Dt����`�����<�:'zE�d�K�b�*�ބjý�A�\�Փx�����fef���L;̧�Wv#�/�5��������K�*���n.[��p�ϥ���@��W
9XO"��G�3��zD���p�W�"�p�7ܫEK<�Ճ��g�Vߟ�݅P��2\�y�K�B�2'�
&�]u"Dr��:�$�HRU�r��VY�0�N�����O��W�^qɔ����'ݸ�Bb�vf)�3�J���B��]��x�w%ML�meC�� @x~���Zx�P��84m+�k	H���;i�!ON�6!J�Ȑ�Tl���2�U[�f��΁(��a���&}s�eA@t񮞪���t�I���:�#ԫz��9��<�9Rt禥eC��*�fu�h>�
x�IG�`C�1�pp�}z�xs�V�����y{���oo����� ��C���;-j�?�)����FL�N,n�s�k5U�u!��1�pe��g\������s�\Y�g%u����6�E֦�K��T��p�����iཱུ+[]S.�ڕݔ
=�}E�L��#*7���1t ��~/��F�>����h��{�{A(��w��8=�
��U��ک��q��;X��N���<q���w����o88[�&zc��sn�Ȩ2d
�z��X1����j����.�^�f�a��i��U�C���pύ�|�U/��=�94�a��`����vD�ꉸaD��9
�x���Q�=i+��)�t�u��<.��@	�6��ؐ]STp*����W ���N�{���
���C�/����R�oS�R�++��\��Ep�bM�h�:*�xOH~�k��w�5/
���<�חy0w��BDUFH� ��!�S<[�:l�o��~uD�N���� �"����mP�'�x���\~��f�#nM�����C�8�r����,륇lf6/Ήu��vή�7�0{4��׵b=�R$l�@<���.m���gf�7}�W���D�)��m�Q@�ŉ��"3k�<�!W�w[�#e�f���]��f]�6����.T��������C����f�<�k��=�d�U�E�T4��k���ѿ3Åev^i9;}��B�`��k>�r�KV�o�Gs�n<�m�����+�"�^�IT�*�S ��0f���d^��㸣}Gg��c%.�$1P�hB6*����*8W��l�S�|o;��TF�T5���$�Ь+��I���Z��;��^{θ1�G�V�>��r�ƺ��+�.�D���f����9��A�@�{oCz�3���X��k�i�����[Ĉ�.���:ca���!�L?�*aq�U�p}��F�n֘�e�<��ҵ�Q�u7S�P<����\F���z�d+�#���n7�[��k�'��M�`���N�r�L��5�ƺ��rlLk2���&	ũ?+꯫����ج����@�!ʘgR"��C(�|;k�)ZvDj =��=ꂕ�P"�W�hy��T�� $���VV����(��~|����5��iB�j����
v�K����=ܕb����x ��>�V;O8h�����d^��:A5��[���b��3kbؙ�� e)Sp�߈r�ླ.7O9.��HM�C"����Ʌ1s�>�Q��f�� �ڈ[�j�h�i��j���a��(p�zl��>�:�<o|�h	Q9��Yl_����]MS�רg��<rj�&�U �c�,�ý+O�FIq�b
`sU�s�kR��r1}Q#N��)X�sQ�-/*p��}H]��X5�5���YE��S
����=��dru��vF��P����A�{�-n�
'T6�=�V�$����d�A�	���D�u�����bQ���$���������U�!�µ�x��ǅМH(����xH��dr��U�,n���b��6��;�)���#��h
�p�>�X�0<|+	�o]��0�GDN.�?��
je]<�/{�ܕ>��j�Cn]Iέ�j�C����]�XxǗȳ
nc�#�M%s>R�WH�"�ͥ�1�$/<���0cn��B�J7$T2�����J3Q�B��<�����se?p�W�k\�h�g@d�T�)2g�Q���B�%��aϨ�h:E
�k����.K| �8�V���[s���(��pɳԺ�]9359T���ˮŻz�.�ySq�/�{MK.�o���p����P+�����z{�U�&ؼ�Y��u�?%�2�H��a��0j�F��en�	 ��v�9/t�,-��=��(��:n;q�rcS;��K�\d��G'��z"1�bI����і��P�q�*}�Ttk��Zxm}�]d�}	���on��	S��Oezy�Z���u	ɇ��J\K�n[�s����x �i�f�Ţ�>K��^���Ƽ:,:*��76�4�۾���{�瘀�À���PR��DC�S50��f��6�P���MB~��i3�u��<�~�e����8�fx=�3m���D�BX����|�����4α"/GM�w�Iv�Na%��#��h�yx`�,֍R���p^R\")�����y��u�ã� ��
3�Jzd�˘2�J�&��I��k�t��\8N����˨R��q=�v_ �����|q��v�;�W[�-ێ�97�M��F�G��y���Vk�J���)K����_M��85��\�c����Q	�iΖ݁n�ֳ����љ���������X�!e���:�C��e��\E>�*Kju���t�o�X��ի�����M��S��m:��ͣ�n�i�|)VP�5���ow�����I��/5I(��j�Մ
�����}�\�����C2�;J�7s)k����ǂ��ٕ��)�x�#�� �β�0b��0�&VKӍ���\Qi���{�j�86�l&r�hԦ��oa��à�=�5�&�U�ܺqM�S�+�E��B�W���8,��KE	X�h"U�T�u&6��Z��Fū�.ǜ�z)�C ��fu˨:��
������*��j�`m�[kɴC�`2wn��U˟Ts;2���ܾJWV��khqE4~tW�r���:���v�J����86�3r�%�*�h�E�1�=DT�Aˉ���Z��Fn�]YY�bc�� �wM�bU��Ԧ�a[�}u�D=��kJ�A���Q\�(�nԢ I��TM+���̌HVe��	W�Ô�*�B��2˒�ݢ��a��S�R�"&�̆K����r�&Pww)ٗ�����W��WY��5m_� (xl*!Lr���3J:���18�#h%ϥbV�K!��b�D�p�s3	61��v��ǂ��̤��)b�3$��G�B���2Vit�о��҄bU��r��@�����X���TM[�o-,!R�XY tU�l�B�(�� a��N}�e�M�4H���*@���h�n�Uf�u	�Wp`X/�mMb��V]�D��ݦ� �brG"6�ec4�Mx�L	�R�f��Ve�w��°Ԙ�Jk����[R��V�~�������:oW@�oe5&/K��N��^�-�sʜ&��,�UЫmDU1R�c��5��K�r���q�-�r��V*�q��pUdRV��1M6"��D��D�b����+�*���AV��UE�q̩�[1%a�K���Y�+cf&k1��"5���4�F�T��c���B�M2��f8��a�+�s"�TE�S%�W-������ʕ�cu�&�J���k��uTuK�*�ikfaq+���.�j�Hc�Q��:qs.&!�Ę��\%�Ylr�����#���QLe�j2�Z���8Q/���9kR�z�g4�V�}A���ݘEE3:K�؛�-�buӚ�k�)~�=���M>!��5�Nԉ��t�^Yʘ#��hp�Ɏ<�,���1��k�h��Ny����=5T$�nza˜���C�:^�Z��\��]O��X=��~�����c��K���M0�V��y�0�Z���¸LZ���������p��8qB HEҫ����wR%�TT@Bgn��Ѝ'P�GI�J�j*��:W$pGM�d�&�@B�SX���R��z�Q�P=��Y��u�x�5�Z�+8��.ҥG��b�v~w���oV��$��Vưh}���ܶ��i�j�=.�ފ��ش�[wf����Gp�\��.��GL�$xL��� �8�O_"_����0Tr�@�#�*]b��ᢐ��x��{���VxT�J��5-ƃ�T3Z�54�Y���^Kso]�X���uyGU�7�Ɣ�d�m�/�,j̚'lZ����j��v�l,���AĪn��+���;l�g���o`��p�<��h���UeV+A��.�TM�[�c��q��&�
�v�Efܺ��\��%^HZ�`{M,$��F��|#v��n�[A��ae�Uk�PK��g�Avﳜ w`_*Z�z)�V��vZt�[��ZM ����r��:�k=�U5/ۂ��S2d��B�[�K: ��*[
��ϲw{�]`�]����ɣW�C����:�e	F�h@7(���)Ze�I��������@u��}��5{�Et��k|~"-���~�gv��/5R� 8~�u��X����x�C��}�^�e��~'!wʗ���4�ǆ�����)R<�y�r�q�F�E��){�A����N��G\ï�M>������%Z�I�P�5��M������U^Ă:-�|�����­�����xI�1���{,D;k��e�ղg��Z��J�k�r�^+ؼ4`>?`��^���=&���ʜ�,e�C0���Χ0���ѕH��W'��u��`{���g�$��)�%o��j�o�fD���	4U���Ug����o��ң��jC����O/L?�C]�q׵l�im�i��|�L���5N5S��"�����3�A�97%��C>�3&�N�ͣuhS<�Il��8:ȥ����⣠�(�y_^C�93t1� ���͉�`y*Qǭ���W��R��b��m�X[~�����s���U^��k��+/��ï���u�;�f���Wd-d�u͒����%9,]\���0���$x��)d+*��G/���5�ԋ��vt�`�*1 �e$TeJ�qr��
$�ڰx񬪨�P�W���њ�R/�^rրx��נtS����]�}<���)�N���4�ZU�Z8a.U�w�D>*I��O1�c)�@p���հo��k^i�>_I���)�����vZU�Y3+UC�R/	�����jy�`4��S�u+�x�j
���VsD�K%�W��Fz��x�G��k�3Vb�קFC�7��/`�E���o3]]F�Mmux�>#;(p�-��r�*	���R��L��x���V`u�o�h�!�ZLΒ�C0Gd����,�es��l�#v���v"j.��Y9ل�mJ|2p���(��8�r-�)����U��x��-�x�<��8�Պ\[�Y��5����W��Ƌ ��VŢ:C�0=���*3edI�I{�U�
"�|�n��UZރ�_�{(�߻�<�1��X����/�r��q�$�)P����ӻ�qp��}�gW,؁�T}᯹6�yJĳ�q(fلl=D�yc_Gue�5���f�h҃{ר����)ۉ�B�/)�%+ˉ��%t��й�O"�α��D��<��X���Cea,Ʀ�+��KMt�hW��Wt�[�`���xaю�Ά�����\��0��Ư̔�,Κ���Fý=.����ң���Ri�]چ�5��ە���hNcq!�kw啟6��P�pš�^a<�7O_Gl�r�+:�s�}�Nz�������+�Syه�
-�Sb�*�����+Qw�xd�v�{�gZ2L� ;O;8�i�̣o�xE��v�g���K����2��:��"�#b�ǈܮu{9��V0b�`P�J�GÇ���(�Q�.�W
:Qƈg����T&���-u��D�7����ф@�El�meu+��0��j$qh-�;(���hd�^�;���:�(w��F���T��fY�U��+���"��E��f���5�sb�ھM=@���FXa�(��ܛr)����(d�z��N� d�W�]�:{��/"�����Լ/D�t|.�7�ʷ��jq�{:�ee-۲{�[���U���0����%�*�WVKz[+�q���In]]@��pId��4�Q����o��o��������ծՓ)�����,�)�%�F��i��l8�5��W�.6žE�۹%:���d
�<	�u��VR{�R���D���&��:�ׯ���Q%JX��blvr"]��(d�
��؍[#�{59��2�k}��EU-�w�����uЩ�6G��6��[�����(�
��R\��g݂$E^ԁ�=G9�n(u!ٍ���;��ŠK�8x|�;&�Mc��t6�
д�t�*W	w7!¨5�v�vMC2Z��v��)BxM`�����gYD�$v���>x��_���[B��Ƴ�:\�U/w��M���uZ]ПQ�˅�coD�̉����E�5��Z��uA7�v��֊v���/X�<-�#���o3\�VݓiqmWq��*�N�<c:+A{��ʪÏ�=�Y�ݼ�r�P��m`rKe�y�z�M��m��y�
Z���cx=���x�th�"���fQ`��ѝS��և�qC���~�+t���,�Sd#^U��J��}����6vKԓ�=��bke��J���9���j�׍��c�3%+���%+�mw�C���V�m�a൤�����p���R��Q,��1��_7u ��ћ�9\�������lH�:143��3k%I)ZU{[ɳ�͘���)�Zjx����*�KT�48��n���s2����.I�y�:	�!=R�i�5�6툫���i\�a�J�XB":BԮ:=/���m9�t++t��B1É��T^���L�h󩔊��:�7��,��φ��kqc%�p�|Q���n^���)v�F6E��W���JC:|�V��x��;���糯���_�����BC�L�h}�V�����'�X4��Z��*9}���h������ť�-�[��e��i��V&�=���5�����PRB_$�^��*<b:�����S1[�i�i���=kwU���Poz�A`�gz��\�e���w1J1!���y��خI����;5}8	�2�"��󛞾�ٺ�g��eONS���r4��Zn�V'v�ڷΥc��\�\�~�&�O4����uӓ[�osMu�7lR"6}��IƊ�N]�S�56���@�4;Ǌ�\��0x����r�:�좊�}�,ndE��1����&��*��/�����QUY��>�Bh_b쉿7X��R��'i��F���~��|�'XL�
;���b�kg����>4�ؒ#�"�t���
�wj�A����.�Mh*�`���ˆ�Mb۷Ns��zU�L����#mlA�E�v�i��R����t"�4�b}׃age�C�Nrx�������wvd��X쬫�����L�P����0i�d����ݩ�8ԫ�|��������@�;w1���m*��獻���r�l�#�jYJ>ح��:��[g#&�����
�j��thk�V��AZGy����
^�%��ï���#^�f�b���z8̼U�IM�]���G�(�8c��Z�Eu�E��0V_p#9լ3M;a���3XY|ܮ��*�u�ƪ�n$��z��Zt�J�c\*E�'T���%�Rk��N���E�R�⥗Ҭ����,_v�Qc��j֭�w��[ �0w�����R-�}�
jƒ��uղR��k�.�U'u�D*,�LS�&E/!3y���
R�wR�lT�VAa���hEm|�
7D˵�*6[�%gзy�H����X�'����Ub
e��r�U���A�\ U�*�p(1�v��Y�Rg����v�&;X�X��
�0Z2�Ux�@�q#v���B�c��E� ��>2���&,��c�*�a��-X�6�2�K�)H����e$��^Gq�D��R�SH �qᲞX�+
5�YiB嗎͗V(�X���a�9R�Nb(��8B�)wN��d��лPլt�1����w��t��9�%W�RL�MI8�
�ⷩo#J\��.�Q�lpz�C��.f+ۡ�P��6Z�(P�d���|�؈�ff�YSL42�E���Y.R,kI\�2%lQqGj���W1E���S�eB�f�2�*�*"Jԭ�mq������ffZ��1��J��"c�M9�m��X�����:")J㘮7-1���3T�`�1r��Me�\Q���V�:�\�´3)�LJ��l�b�\�:j���d�Le��AF,[��%ʵ�Ć��q��E��.9i�Lʲ�n��k5f!����P\u�i11��Y����^�7�����ֻ�ʖ��nty�S�ΛҎ�D]����q��oq���Q�+�1�7�=]Y�֜=yyN�W�l��rY�,�6K��(����+��+i䩡��Q�ϸ�V�ois�k�;
&�,��9�֠ ����8��5x�Vˑ��B=���߫��9��
��@�|h�uhV�"݇�u�jdF.j�E��f��kf��<L>�%Q<�4���U(4:6�E��k2�2>Z�gy��6�ˉ�[)�*kN�$����n��K�!��Z�F���{8��nh��d�0.��3�MW�Ո{�v:���unx��B�b7�S��\b�:fq줕���[�@|h{���u�P���k[�.��h�6wcԱ��X�z���9��-����>��}6���:�WJ���4��L��a# �n�uBR��h�J�Fa*�@�_��.
rn!���OW����Qg��� �$5d��4����||g�L�t�~Y�Ӽk�h��"ٍ��ǵ�U�\� �G�<�������v��>(�ϴ,j�ST�u.�Rw�EGi��."�N�;�F���F���h��ZCk��,LƳGLU�x�f�ǋV�H�����9��wP�Rf��Yo�L��ܲ3�
���c�s<i�N�#<��J)��2���G��B��c[t&���JWO��~�?c���ML���:�٪�	��y�-+�59�r{���zNΰ�V� o���*�.�h��vJ�8��
��RE��y'�����������ma�7�.--�HM��uf�!��V&s�f�k�-ܦ����n��n���(a�,Gp\���M�L�E��K�4ΟY}��w�8fo�)6���D����5{L�M� �0�Ԗ�6��������1j������k|�����D2���1P.:��ƪMV��TzFk���s�s��U��O4%¤�z��y֤�w�A�b�횂k�S$T��QH�����D�Qg�8�z�)S��9S�Rsf�[x�IA�y��V�k�v�M�luv ;c�z4nL�1Mׄ�2���$:�5��Q�X�<��|�����ܻ��갹��{v���z&�����'�L�^�y��9]*�ҁ��ˬ�.�%b ��G\[�T�O��]�b?:��2�;������ӽ���Kѭ7�T8�QMbj-X���f��������^r�7�����m9�p�ל-��S�Fߞ�nx��\'�4&k��Z��)����py)�kt}����Ji.k��Ḗf��y��a��Wr*o)!�]����B���̗�n���Zcf{DF�I<,L]Gp����̣zڷe[X�8�)w���]��5
v�/-��2κ�k"���������v�[�;4��AقB"��ZW��,Ԭ:P&xWY���eb�p�<:�BÝ�����.E!
�X���">�l�F���ӹau$[/��q&��8����z�TS��]k��!�t�}l�t�<K����Z��x��؍JښS쉩��}�Ȫ��v����w�Ŏ'��\3S�l�m��U�9<���/Ip��4�z	��IY�ðe�8�G6�w�t:n�ꖯ�7

Smf�`S�"rw9�sy5-,*Ǭ!@ǉ��!��s��%"�/+;{�X����P[�T��f��,��S6Hcb���s霞ͼ��isշH�)�8g"���+\���#�^��1�l9�uu�<�i�����w�^��J?!�z�\B��^��k�hS�x���C��(]ى���S���&��4�+��zi_:�0-�`�)�-9 �9��E��~���41���8�qI��IE8��{���ϰF������4�����g��t�:AW�=�r��@�����1,D��{[�v
)�fC�C��^��&���m��X���G��#����z
�Ω�������l9`W���s���/q�ۦO�)��:�Jw����������l���xq�(��HB�ܯ�=6�����{hM��[jK(r������R^�'#Y�r�N����t1·$�x��R�Gn_A�4�W�Cꂊ�K(��oo��y}�y�9��d٫"\�K7�#��' [��l�e��No�8�W���V�r����>�!���g��P��T�����EPk�4۔"���c��a��dݮ��9�%�ߙ�P�5�~�Q}]��8�_U�ۍ�!�`�,��XiW�`�:�ۆ�����by�Z"_�ى��o�s[��8��P3)(P����w��j>I�=�]�H�����7���q�j�i2�t�,r+kDWpm=�ţ�Z�傮KZ�8�J|�_E��Q��F�����9�ҙf�qɜ9�N���v�>���vyK#dQ��6�#K�n���6u��]�7r�r��K�޳^��,.�!.��]��Lv>�Ղ��o�E��1d�S\9��8̑�!��"6ӑ��X P��������R�������(���a�O#���Rmbǋk��+���[S�Ɂ��Dt��u���(�0��kN��N<|���=���I��l߮����:�����i�.{F�.���Ыq�㲫��،�{�v�!��j��]"^4���Z��W ���Z�`<r��Mf�旕�92�e��+L����S=��s�s��⡰�`���h�G�urtDz�"������H��t�\�`g�V^�E���=�7��-о��w��@�;��d5�C��N�Ћ:���Y=P�Z�-�,�j:k�6sh��qi�P}W��uΟ!�l4�����ݓ�b$�MC�O���*5H�%�y�:���\���#Ix���옖�߇��wB0(�iAK�<�6z�d��n-��y���K����Oډ�#k�p�����m�[KV�,�T��v3���D�C��sW�(��6������d�>��oG�r,�J�׶��Cw]ǭ�?{(һ�lO��_OOA+a,�y�TGk���Muo^�~{V*�+/7ĩƽ\Nj�Y�E����3[��[���j2�IK��:ڋ{}�ʏ�zX�x�.�p���h��O_z�'1ޡCnD�ͮ*| S�*%9޹���Y].��x �w�ԭ=��~���.fU�w*h��5�P��$��nL��$�.���5�8�$TrFf�vr�u;�%?zN��pvpp~�MX���Z�c�����j����^���C� *��$��Y��^O�B�� ���*ʪĭ��1x����vS7�Ų�����$C/;4�īh�9]F� �e�s]p�L�h�݆P�����ۊ9X��{*������)5	����<�!3Q�;x4��sv6�y�M{Nu�b�Ќ�2md��i2�'�?w�/>�r�F{���Ҝ�����L�<^��S;FC��oVt���7����s�c��3��l�M⺐Y��H�M� �}DfrU�kq��]:������)\+�u�����S����NY!�"i�8����\�{|-�/���أ��r-�J�f��k�EΝ[[P�9W�k��y�o��ם���5�.�'���m҈�nͭ��x�S��\ф�q�S/3���g\�t�����+ǫ�f�5mp���쩼{6�ef�82tq
[�ۢ��Oaܭds�L=GF�ǌXn'��T�S��7q��l,�mN���l}կe�����U(*����	:[ٴ@���6���Ѽ�\Y��/��S������xPκ%��'3�s��X�c,gk���d��D��jڗY`�*J�y5PY����d;|5����x��9�������%ɖ	���)j۲�����`��:�Z��`x�u�:$¦�-}��v^�4\�Y7�jy��mud�ޢ0ɑ0�Q��rA�����d��	[���e�iv��<�Ǚ�RY]m��L�Z�׻D�Kʶ���$if�)f�;OM�P�k��47�[����5%%�ׄgv'��8�˛��G�`�x	�ǲ$j(*;ݤ�����LVweK�Q)�r2r�d�����˸��|�u�t�Y<n ��z�2�c� �{�xWm��muX�y�3��w������&�_U�{��\���Dӎ�Q�͕l\��	�&E���B��;J��p����t�0�6X4�m����>�-��.s2��ض ��8E9:k�o��)�;p�k����Wf}�q�S��[�3�ʃҊ�[�Q�Ċ��Z/=+f�8e$sem�j\t�Ѽ�-�T\��\�CGY벨Wo:EY��]wV�N���Ir
��{�i���J+�YI� �ɭ���
x
f�L �꫉e/�vF1it�w
68�ɴ2�w��{q�T�|B |� <ie��qna�Z��9[(��-]R�Ak�Tq����uj��c��[]a�L�¢E�\��d�����iˤ�SN��-�[i��Xb�T�-Z�����[sŴ���ɚJ5��%����5L�W�ciWF��5-:��SOX�V��䮜nJ��q��h�-m�"�Z���1��b����Y�幤����s2�a�j�Bk3WX�m�+q*kW
#J[S��\���C�
?1�7^��Y��윶¶b������M+���Z&j�p���V90������m�Gh��u�A�xd3���T�JG'�+��2C��fs�3��\�P�:3ڡ@	�(d*��JB
�.PQ�J���P��7btR���EW\�)�N�K��z���r�p�;��.Ѹ�U�	�������S)�:�^�N�ӭf�vj+�M�y4T^�{��RGgc�g�5�����mA���u�r)Z�j޴M
�0��X����f��3j�+/YE��j���温��|�%SMWDl���⺣���_��+���A�+o-�0�5v&�T7�h���0&fm�2�b�,��D%q3*�m�S��G�>�O^lu{b�{pL�H78��e\7ӌ���d�+N��R�Z���Ҍ	U�SF�>p��oL���!I��ٱWB�Od4�ƤoSw��x[x4�ne<t���Pڊ%��t��t������Wr��B
��AH{W.���y,�j������ӷt��U�Ԝ�EcA�Uk���q����8��yK6�H�J��`ݲpPM2Z����we��FC�Œ+�$�cf
�.{��ə�>j�����fKE]u�8yw6Ƹ�e�'Q�xC��N,��]�|˸=p�G�%voc���fQ{A�F�J~��˾ݔn�c�J�u�����V����+/�����:�b�^���]ضV�wŚq+��wmc��ݩ�0N8ڑ(�.I���R=3[�n���F����q����0������qSia��gQEaW>�x�m��/v]`�5�sLT��'�	��̎��U���#U�Ӱ���H����,����>���B_w?0O�F
����gnN�]��zKu�X���W>|��c�y�F�ٸ,����gܐ/����1؃��]�7L���M޲�>f��c2�@h���zuf�M�Wk���:�q�\r��ي�n+og9c�e
B8�����$|�����<��ຳX�U�����'C��M�ZV�2zi�AC���O�O_]q;��%#�����z�wS/5���gn����ˮ��DXwe)ob�ac�2�X
�%	�K�ΰ¤C�{���=6���Z�^΃��O7X�͗u��E=UD�_k��(:ST��X��\Kz��꒤X���y�ǖ�B�ֳ:@�B+������VN҅Q���R�(���+���1o<��iX��D+���閡)Jc���}W�%.�@�o�Z��݌��񅲹.��b�g�(wKf�)4ZOM#kӔ��[[F�k�#3K��c֕Ӄ�y_tCŶ�&�*�Ӊ5�f�����8�[in�kG����l�B��*���ݼ凓Ul;)��%�/z�Bޫoq�/�z���w0c�i��%i�	MChc�,�IRo\��GrZ�Y3V��8����a�>���Xr�^��[�����ۘ�y��B�v����-�*8��8/=Q>�>�ԟ��W2�f��95�X���.D���t��E�n4�\ic5�Z�1²2r(��$J�c��� {Mx4��!;�y�@�y�-�ߔ{��:3�9SF��!�ό	cx�@��S���ʥ��A������݌�3Ľ�ep���Dnt��HrB���>7���o����z�(KΫ2�A�QXL$T4d�����,m���3�ȷ풉�����VЬ��&V,D��b��Q|�n����ٽU1U���G'
���*RA�W�|���G�}�8�w-�ʞy����q<I(J�@�|�Gwl)D�.�u�r�3����ush-��~�v�7��\�)�����_^8y|Q1R��fs0� \Y�R��r^yy��n���oF�jn��/-��5��<tj(����e��M�V�{��i>�Ӗ�nV�}�Oœ~G�����=�췶�a��m�oW'�y�� C�ȷ��v��+M�����j���(��^jCwJN!��F��{gZ�xэ�usʖ
�Z��9��a�SX�Q;�h#Ykt�7甅G���zẶ�> ��,EtT�Ȩj0c�e�ozM��I�����4�,���Av�R��}��=4�_/��Z�*�Cܒ�7��e�\LŨ��z�m�����k���QR��z���&B�j�6d��8=3�(�p�5�:�J�y��bٖV\��8IN�f7���%��;M�x0��t��p��/N�x/H�S�%�,���zi,&j1̛:�3мX��U\���E��S�����.mG-� ��3�7;�p��-=%���[��zc�5欃�[��Qq�	L��kt�����Q�"����m��×I�-*pވ��1f)�3A+|��x��f�6�]�N2���@|��ʵX|�uL��d���&mr���=*�;��Y�0���P�}��y8�Y��ߞ��uw7��j����Q{�����}$w�4���t3�����g�bd�]v�j�}�]We�����N�DY`Ь�[�����_\3X�Z�w��ܤc��of��YU{%-ڑui�TMʛӺ�Z)�4���)�&׼�����Y�i�|y��̬�m�[�����I_��}�j��u���"�ڹ��N(>�ͫ�ǠI�F��׷V3[���a9���zXu�bc���}q4�|���\Y�O��bR)�z{V}�P�ܸ�-�ju\kԔ��y=E7z/�e�+�+��� L�j�����\.�6��[I$����J��0�ȣS�M���������������c��U����rm���sZ��p���Ꚇ��Q0/��l���.�*���_v�o�m,ڴ}��_V� ��	�f�3���7*m��ݳ��U�fkF+b^���
�J��4iޢn3�=3J�6���S$��:��s�EK ?s۔�����r":8�b�|JX��Kfn�ٍ�hf����yyПNpnƿ^�4o]�P�y�S8��G�7Cr�B�V�5�!���yq�R�y����˚����G7mZ{���7�84�@e�ܘ',�EBHZO�L��ɴ1�4�w��u`�Um.�k�݉7��D�����F=��oz�����4&�{�GM��ݩ�e�.�(�=^ �׳Ϛ�YM�ѝ�}Ő�	�45�q[��uKK�]]����y���0�M�6������Ro�t~�5S{t(<<
\�OJWw|�`��Q��(��d�mvIdV� �K������PϜ�!�Mfe����l�[M7��u\�)u��ZRfj�T�Gŷ����">�7�^�+)�+=&cB�c݇�I��D}U��^]3��p�1[�e¦��x�\(���bO;��Pk��z������^qB���Q��Y����ڮ�nPB�=E������[�I�gN5������=���oZf�g����,���'�}C1yՒ��z�6J��5TiY~e�^r˘��t�� �qK�3�D��{o��ZC�7��y��� �����g�/G��q]Y��w��5G�Z�ݞr0Ԓ>Jj�841�y��m��?�`�����S�ҵU�T_���$ ���οR$BC��E�L$BCY�������:�̙���=������N�5�8&�� P� �$$�!! ���EC����uᓣ��x����B�R����f���V@�B�yc��z��Hx�*��tM9[w��k-��=��%�F�Q�YJ^e&,NX(���C�D<����(y�dό=
Rw7��$��a@p����<�ɠ�$?�5}n���M�Ĕ�0�I"�Rg���a�"�-%����:�b�#��Ȟ�c,�6\�����:�N�iВ���"D$49U�w;jJR��d\��*E�F.��
Fr�/�o� ���Đ�ѭB��3�"���F��3����<��Z���O��!@OOӢ�D�o.&?��b&�@� ~�I ��?��$�J��K.���fu\��W�Fspe���`��"D$6ɔ��*�������˓{���{��-zT�w��Jbo=���<�;� z�B0*�  Џ(��� 9��*���"�KISR��yH����9����0,��˅�MP����淣��.�1�*�NbO��n�=f��$�f^����3ot��Hn�r���r���z�[f)����]J}��W�ݡT��a�D�R�!!��>�(�=΄�6Ť?Y�ks����Ox'�1bF�!䌛o����o�(,I�2`�$C��I���	$� �T��&)���.FRb0��Յ5B��V�� (>��!�N��~�	/Ik#L�c��r����D�Hj�<��G�ZG)��	
��'�'�)$����I�}��lj�؏�jc���.H��8ɱ���.�Qupw��Y�j�Q�b%�1�F;#Da��V��Hv:��p�*�H��A���F��D$BB�{12��]��H}����}��r6N]�9�Fy��x����*R����c�j�>�Pux�l�#7Y�z_weV�O���ij0୸y��BD$/�܎H�(ǜ_�$��mߖ*�
xfYMƓonk��ʋ(س>��Ca�bb���蔒D$?�T��^y�Oi�GeyO'	��ςI��'c̜"�$��e��L�q��d�%C��xz/|YH�R�Q��:�lD��g?���)�4֛