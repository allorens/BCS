BZh91AY&SY|�{���_�pyc����߰����  aE�ꋽ/�P aV       
 �m� �&��                    �        G�wŀ�����S�|   �&(���m*`5�*�[aFک,��3l�A���L�w�m� ��� (@�  �@� �   ]e�    ^9��	 �m��[e  �4 �6�B�M(� 5Z �1@��6䖱���@6Ā6�h4 B�6
 ��0��*Cl�
IN    7p*Z�(�`� l�-�M�:Q�l�lL��  �Y��
hi�CJ�`4��CJ2     fK@h��hi`0R����A�4,i�d� ƠN;8�F������6(f�X�M�
2�ؑ�` `    �`pV �m����P���)��aF��6ʐ�`8��2+0
m�Ul�4I�KE+l��(}��                 
��%H@P$ EOM�~�J�H�`L � C   �����z�0������h �" AO'�b)��)➓�d�L�Px�HB��� �   @ST�4jJ{L���~�= 4�)� ����*�jfBh�d�1��a0������Em�(Q���G3��O�o�S��Y&�����"���P?:E`�0��l0|��7�8D�I�UT ���T�>u!�E$���oRͭZV��a��!�:�z��ʫ�݃m��fޭf>�ɝ�����93f�lcw�^rtts񥳦WV8�q<n��������o�x���y�~���ў�p� !D��C��QI�N�飇z�Ѣa^�</3���|:0$|<t���d^��&!,O����<5��<5�d�2��Z����]5�|9�}6�ڍF��s�9�#�r1���Ts���7�p�k�G#��ߔ���
��ESdr��Cѽ�����f�YEwJ˘Gi�֕�9���)ϣ�m��:A�9��n[Xb���4N��Ǣy�����2�ǲ���2�e�:M>�gK:ub���ڴ�����Dgն��"j���F���#�Ǒ�qʭ�l��Mu�")�g��4��*<�P�J�l��";�GS�)>DG"#���D�ی&k�E#UQ�b#{�D�<�Y���D�R��+�F�Q�DD��e��+�rWXr}QOVԒ��T�DF�Q��9�}ߪ�"3����DLW�m��}]���Sh��#��TGYjW�F�3ʈ��+�=*��ӵ�'ި�,v����G�QM}_y�"5���J�G�5a9_O�Q�s[FwQ�+֥iL}���N�"9*:�ҩ�s5[b�쬫�|�J���R5ڎ#���}�'*<��Gey�W��i�V0��9Q��qu<���m��m���i٬:w�E�f��ka��mt:�Q�#=�"*V�e�T��UDn6�*"'�=+e�����=�8�E=�k
f#q��Q�m�i�9��n��;�aĪ�+���y^O)ﺜq�#�*1�q^g��fW�fWXq��N�J���=MF~�>��I�>��z�Uy���'����V[zKH�Z:��:���5����Kn���>��|.����,w�I��#��Xp\>�Ǉo�,w��Q�lx,<�³�p�gO��y�E�z�њ=�|.�����}���tǢ�j�����:k���oO�|{�E�i&� D�����V�N���W6[v��t�\q��=.T�}�v��)�0�Y�cZDsh�"$m��;c�m��DN��q�5b9�aȧ7y��{��a�:���4e��Q�v=�=�qƣ:k����ͽ�;ߘV�o�)H��Q��u�"}�R��2�r+Q�&Q2�oJk��ц����!�v;��-�5Y�3�k��J�FݏG]{�w�:����*;*��NE;ܹ�s(�[��}G����۵��y�4�VV��S�B%8m���93CP�r�a�V�e�f3���"=a6�0�+��7߼����Q�{��f2�aȎF�jO�;�R=�D��O�&���Ǖ{����;�yޣѧ�u8�e�#S.���森��O��S�m�Yf�"'��uH�G�a�m��";�F^�o�}֘Dw����<�1��R1JG�c(��G���cDF����q4�i�)���"9��	�"2��"=�a>�<�q�#�3�<W"���#�Dy��F��2�ѵ<۩�c1Q�g��3a��j";�Fg�a>�"#�DS��O��qDڐ�"���eԬ�L��yߢ<�iJO�F�DGt�'�L�̩�!�R)؉�ی妹�4�RaI�~�Y�iYSQ��3EDy\b6�F��E)>����Dwh�y#�������;n:�y�O�q\c�D{���mr8�*��Gc/i�}�\Tq�*<�L�T���F��G��4��y�<�\j{��Қ����TG~��v�>�e4���;�mOqO}ϸ�Dy��ZL4�2�����o����w���s,����9�q6�Ҙ{�;�G#�S�G�����.�߰S1��q1���ӎ6�akomZ��9�Q����*8�zq���!��[V�G�##�o�U�+��{�o8j3��Q�U���#�B%<�=�V��U\G�ͦ�!�B�ˌ��DWQ:�RR��a7�Ty��w�"5�Ds��*6�GT�>vF�q\q��#�Da<m�ʑ3Q�=cJEa�#(�G��I�y�YF����#~G#JDW�m�TDs�"��9Dq̢#�J�3=��:�mH�#2�R"���Q�����_DFr����Ȉ����Gx�Q>��m�z�ˑ4�0ɘ�n"6��]M)E;�4�R8����H��\DFcl0�H�G��#��"=��7UM�T��Ee����y��XG��9�і�<��aF��GN��(\}!p�YQ�G��Pǫ�}ߜ���9�v+
{(��������Qͣ�G�"y�9��0���u�b'�O��<�6�Ga�RR��y�i�#z�4�9��t�>qʭ0���Giz��Ә���)�&�Mi���0�Q���H�X�̣q��<����F�kH�0�m��[��i����St�1L*��;�cHwF��p�솶Kv�F�b:�L��5�l�q�m�J�:\!�}.�#6��m����g��i�6�Ǽ�v'�<��{�#:F�G4�4�D��eܶ�T���&�9��Qܻ�GwuQ���EGb0���{or��Zc,FZ���:�7���9��Dl����ApO
D������,V�_N�x٭��s�ҎY�(q���q�8ޚ�Gp���V�i�����U�8�1��󈭩[F��*��Ft��4C]�2����5�GN;��v;�\�3�#ڮ7�#�F^�Qӌٱ�A��ie�R�gG�!�tt�:k
�VҊ���kk��s�9�,1Q�C �2-6�L�R��Ƒޣ؏=��1�c��#;u�0��*#�i�{�IZR}+���DG~��}�'Ȉ�r)�Tq����&+*Gb0�}F"8�"}m��F�Du7_O��ˬf�";�����,�\��ˎJ��Tu��a��[aI�Do5M��F�Jwꨈ��#�QǞq��}ϹQ�f��ku�DuY�JʘEn�5ʈ�J����G��'ި�(�TF�Q�Ty��R���"0��7�T����8�i�Ez�5��6�n�#^��)�[S�TF�Q�Q�^�H�r9I��0�+*�_6�1�MU"9��;+l'��br��sդu���Ym3Za����"z��;+��&x��y�X>f����8O���d��h(�#:6ή�Ek��-b�#�m�TDO#�J��u=^i����+5L�G9�F"}��f8�����n���Wj�Ԫ��U�uWS�G�����b��W���:׫�J�uIڌ:�]q1Q盍9>�E5���S���$�o�N�)��^>��l�"1�GKgV>�>����Ɗ#{rC%>�ܒ���x�'O|6x��Ӑ���Ba�^İL=/o�K㮶Y�eFi�RJ��Ig��*d`���'���P9̍Y�؇�f6�z���~����	�%#��۫o�M�����)��JW3[�.�lx��WwJ2z��l�y�Ot�=��Z�/�S��H�����2������k3+s�$���nR���v�ZJ�d�__y��w��~��T�gO�[�I�:�`�z���v���\����nw��l��]oN�˗6i�2
)Z�3Y+JW����2�R�u��g�n� #�OtvAGS|[�'�0��J�jֻ��=��z��+�u)��ӽ��o�<j�ݤ�������ry��CNLp�M�ɏ,��#Θ"�5w��=�0����S=�u�o���WP��cy�ɞ>m��z��՚=��`��\�V�gc�c���oW���w͆"�ֻ��+�<�y{sݽ�{{����Yfvޛ���c��h��BA���<�n\o�T���,�N�Y����tt5�����k��t�_��Q߂v�6l�|q�)�B���:�^��G���� �p��qk���w���Š�����ufU�x)��Y]`��r�M�tt>��{DK*�����Yz��vl k�Sg�ǩ}}���ݺ��w���u�'��t��ť��!O��.�B��J��}_�������ӄ�����:���]l''iZs+�Bt����:�}/s��%�+`�SzK;���7Y~3 ���3s���>(;�2��5^����""��ky�L]��J�����C�'M��8��qā�X٪�ވ������gc��؋e�Г[,��y��D!쏡��rt>�7&b�{鞙A�]�gۥ5������g��$���<�\k�o�z:�8��@�x�{�9F��T%���ڻ�l,� J�nL�w���9dq�Up�`ӎ֠x�O94�Fh�fݗ����=��X-�+h.�fIwP�)���{}�,��Y.΂�X���C�"f�T�)�G#��2�~,us���8�	���^�*%��|��231�>,0�ow	�g�����:AI
�W�#�!Ix�ix�!�k(I�G��o���"�;��ni�ڋ���z�E��䓕2��^8s:����q�"����2�V[���ݶ��|�-?{q��fݥW�v�p�uǵ�W�Z��P,�Ea�w�w:��ɒ��
^yK:r
Q�κ$$α�y������t��ǹ����*Q��Wz�Bŉ�C�����4�}�Z�"�v�LmI�Cpf+^�A�rv(��7����qG��Q�Sd�&����B��gm��}���x7�3�v��ؽK(ym�� ���c ���ۉj���ѝ(��c��0ߖ>]�iE[��!(�˩��NHf��!�K~��S�f�>K.�^_�t.�g]��բ!�"��+���7������{�'�8�e9�����>|L$;�z�Z&�<}�u�z<+z�����'`��[�|����3_����^C{0z�6`����6.����/��޾�,}߰g@[;%�_\i\rF\c�ܙ�k��]�'t�m�c���ف�sniIm���st*��G�h����=E�_�u҂(a����u8��f쵓������(��'Tt�A,6�w6���Bj���լ�f�a�Ҏ�z�}�O~��ҕaq���}�}��ǋ�ɪ�&�C2!�n�!Ǒ	�dY�F�"�`=ek�J�%�
��4��o[d�&Apfy�o���;
��p�FhB�ܫ.r����2����*�f���:^5Vw�Y��:�z^�{V���}����f�̰������ޜ��b��˛׽�^�u�,���g��cq!�����k��k�#TLA�;&(�_N�1/�b�ӳ���wk�O^"�5����=��[�'Gz�ϼ�^�.���ʺ���q��hL�7qw��oWK��0��&2���cSG_�^"_Y�\��{nf]��鑫����_j�w%n�C��0y�O�m���-f�&0i����7}�^�JN���R�������k����c��.ݽS&��5��ڻ�M�1������Kbn�K܏/G;�L�����m{��۳N�	,̾��
W&9��)�ȧ��B<4)�YJZ�»�Ks���=�������y�	�?<����z�	U�0�R�H���:�u(_ӷr�d��@��5O=��s*�o|��&��=�7�}��C�;���B����&wV:�~X��c4˛�#{{j�1�ǨX��-�>ǻ�@>�,/�j�w{Fg�ӝ��B�e�L.��ұh��ˇ�R�\��_`I��r���S���c��6���GFZՎN�4�8�� e��ܳ[�)w[���ޙ�0Tzadx�^J��L�ŗ�d��j-ea���fw�LIa�[ƙw=?jؾľew�<�������E�!�n�^w2𤂩�A�� ���[3�t�g��Ha�"��+��A���k[=z��)��zo^����D]-�(y�ӆ�Ѫ��߶�zdz����V�]��ǦŲ:�y��J7�!�{r����g�S�1��r���VǞ���7��4��kM�#r�י�5W��Y��H"\&Ġ!���s����XX%�N�0��/��ɡsC3cp�Ӕ�i��X��N4���o�a=52�H*�]b&�Ho��J�C�Z������f�s���oO��ſ �MD�d��c;5g�}��]��c	u������Y��l23A�){�95���2p��[t�o�&pkW1:��	�-ˈ��q՘%�"�;l&*p��*����D�э���o}u�Z�Ƚ�z}~��6@�A�,��vJ�I�H��\�[��)���xr'�^f��fIN���&:3]�f?�������}=����_q�3�Do�Լ�~=�I�6�z�*��\�	��p���r���W����g�D+'�s��Zez�\��������<I����ң�3t\.N�0�����>u�WSS�X��%|,<�$�V8Ţ9�@c(Y)t�Y�J	���5�ୠ���v;벢IU���7���6͹�a˯h.E+��ٸ��__I	T0c�Uw>۟kfa��m}�F~�<JF�&aH-�4oڏ��&�͹�}ღE'1M��{�=�Ú��Rt��ynd�+��?Gzv�-e1�4�t��	;��fm�C>����јL钄Q.Fv��ح_cxfǄ=|Y���̯O�X�+���z�#͉ţ�_�z�k'��u<�&��1^����QXd�-�cin{���}��"���)�}X�^#~���x�ur[�E2,�9�Ϯ�(��=��������o˰�?k:p+�^;y��^����:6-!}��0�le�^[ћ�WF!�+���}�ߤz}����P�4g��{��7w���O	܍���I*y%�Ф����9h��'�]�$~������>�>���t��R8{"��v�Q!��ޕ����o�KR�,ň/�w���U�x�����D�I0#��3�15Ei�ڻ{����f��˫^�Op�Ien�ػ��&�6���7f!�q����f����s;[��@�{���N�(�p%���"���q�绋����Xa��n��U�G�FK�����i+͊�����̝�`@���}p�><��ߵ�T!���e�.�k����K�Q[`G5n]��2ǘ]��A�{��T޷Ip�л�����A�i�µ�i�X�pl]O�+���W�o�����{�6�;K��Z��������lޅ�/�t�?�A�/luA0֧��F���0pK��V����lʫ�R��Ͱ��� a5o�"o*XlҴ�[��u�&z��(�{5�OB$����W�����$�e����</�C��OD�.��k��L^�t�BN�V���}�uX��B-K|�י�!~қ%� ݚ�:7!�Ź�����y�S�;�(��':ܸ�hv��D����k��զ|<�����͝H�}�Է;��e�$��E?�.�я�{B��m�-���H��g��4��J���Kڟ{����A�
31�Q诽����{k�`�_nkQ�}���1��s����;�ݝ��w��ze�T�S͛Գ��S�q��{�t�۬kS�����	���T��}���h�j��˙�������]e �� �F�ُwr	I������"�}7�{XЇ{Z��(���-�vu��ވ���4���,�:��4�;rN���F�@����ǹ�#Ij��o�6>�gVd�BÝW7��>��(����O�L�<z�;OR~bSi�w����?#�h�)aBz��% .�j�WL�p�vSDIH�e�O{��3��3�q8�8�N'^1���Q�ؒ=�r�h�����}���F�}bI���T�aE(�R�:s`�ip>E웶��y²7�ܘ5C���ˬ��̼��_�mТ��ENngvϾ�R#�!jͷ�8;�@g��ʞ�8+�R{;Oo����~Xp��ԅ�s+\%Dnq<��!�s�q���G
!�=ե �mK���jI�Ɩ>1��>��n��wh�έ����e0C0�@��Y̅��z���"(��Q����H�K�Gs����)�ݞ��a���y�gZ,�xxjM۲Y�u
���l��3gew
DI���e��~��9�Q�8#e%`I�5�gq�6k��{��H��x��4����c^SC�sPJ�M��Q�I�ܐ� a�"�ڄ��.kf�	Ġ�x`�8�� &¼k���V�C+�ezp"	F�$�A�Dl8�ړ��������bl���O�&��8��A3\�U����	J"�!�a��Dt�j�`,�I�
I�g�d�M��YL?[���U��tɥ�3��dƑ��0�W`[B�H����V�b8Ea�4�H�c��\	��AmK3�bt����I ����C���H�IVHʅ7X��(���$A�ݮ���������D�c�D��E�T�JN��`N���!(�lh�d�"� ȈRD"DDA���)HH�J�M"�¹s��@��,&b����N(d��#t/Lw��Z[����f�BM�Rw9&X���ܜ06���jqr"ԆD�#Irb����.FrHs�'��Ɩ�26�-��R#H�T���uA��r0�HA�܂1jօF`��IqJ�?O����&\A"�-0R��W%PE#d���D��-1�E����!H�QI��È��(�(S)�U"c�pk���qn�	�A�o��
N�� &zS(�&5\� �J�˰�DDĐu�CoOy���n��B�@��b`ѷ|���So;�Ƞ �4 �x:�v6�X8�� E�ڀv6�`�l� E #@;�ڀ�`���c��{ @����{���{����i[X�m��:d6Ք*��R�um��eF*&�c��2�l�Dڋ�3�V�Q���Յ�lli�`Ċ�;��f�޻ �6a�;��������v6`v:�@�l����P4�@<P ��ks��`�pc`;;��{��`�hM��ěIVj�i����F*���,�����M�3qf�9f�X+
�l�l�PSm<sn&�e��J��>�R��C]���w$��I����8�����x�h P4��8`v�@��@��`v:�v6@< �@���6�� �hgq���2�
��V��5emE.q��FֻY�4�jJ̭-�jM��Tī�ni��i�뚬�><�����h F��@��@�4 (��, �t�@@;�`�pаq�������ww  ��N���{���0b�hlM�mY"C�ou2-M�nL��r-l�V՜�6�x�6
�X]q�&��6m�r6�۩�rr�ɶ�#���giɼGk
��l�VëAA�#@�M�i�RJ8֚%D%-B�)�nZ��:����=����&�B_��_���_�����w��%?�����#O�i��6��R��"0�"#M��DaDu�G��Ѷ�B��!S��,�4��6�#��<��<�#��<�:�"#�:�6�Da�DDi�uDE6�#(��"<�"2�8��H�.2�")�GǑ�DF�DyG���F��QL��F�)B�H�F�H��4����:뎢"6�#h��6�#��"<������6�� �S�7����^3ҹ�mg�=��_�"-��ۂf+L�04A؃!��jV�Ǌc9r��b90�:wWVn�c�9��a �.Tr�X��A)�Nؠ����/>�8�$���UMq�"|�k�6��Ēe�����6�2}By1�)*XdG�qc�N	0[+�D�=�n���<�$0Wp0lI��ap�$�a�6� �CL�q��n�#6��kp�Ѩ4,/1iU�7�a��%,)�["b�C�l��n�)5�J�	���q�\�y���X�).����v�"5z��IHd���b� �u�8M��:��a?H0�|�WTZl,� �,�u��P����gz0��5v"P��߰t����j1�(̯
aJ�`�I'azE̘�����[�K�\����f��K�#t_�K�U�z�G��	
HLy��ޔw�Ņ5�*+Q��
2A�+�{λ�vB�i8�$)KUmM�Q�[L|"���Q@ec1Ě%5
r�N���El����2�I�q]"t�y&2�/)N�L�� A70�"�0�<�iLe���_ݝ�{����*I$��]��z��Uz�g��"�wwy^��z�^�t	� �������W�g��"�zֵ>���>��DeF�h�"<�6��/<�\eS�I�Ʒ�VU4FTBN�o[d��S
`e��6X(�lX� �	d2T�.�JU�A�l��"8��C1�*AH�v���AI'��0!!m�=o1	���I&p �.��E~�":�L1�1�X2H"o�N�S�_�j� ���:R�qhᆖ���e�`�ʇ�������=�r��q�3p�K�'�3ěH����K������o�z�Xt��V]�O;�����B8o��#���ޒz���M�F�2�H�\�[�3�N��S��ZY�J�$�e�P��׎,�/3��@�,o�wǅUH�:m�-�^eykqG��P!��F�wpMܓ5y$���Y�j�%��J/���F^�%�.#9�eo(Gl8���3�,�-��޶i5�>a�7H�6Ƿ]G�C�66�4<6Q��:2�=���l��om�5�F�=���ϸ<0g��-6c
F� ,��/)���"S��$�,�oC:<��Q�*�z"1�1iuk�%�.�i������6�a��2їYy���"#��8�0��t`^��>�~��"ﻲh��p;	$�=�)�c�Gime_6[3Gh�d���M2���,���'�p?`�E�M���9��e�FF0��!&���K1�޿]��L���K\��+�T����D��Q"�C18G���\GrݫZ,����f�t�"lVkd�ëf�UC:p���4�0�AHp�ffp�Ü-����t���6t,���p8a�2�\eu�"<�#��::с.��r<��D�Iaѳ�፳�������wS���{κe����!�D%�6:��m�Ȱ��<tz<U��&��L�#�n�'7m�9�>a�MM�:ׯk��^�$[Z������8����B�<mK(��"��JYK|�;F><zF�k*������
-mQl:�.aN�ˬ�ӫG�p�gHp�͜��4l�Uǹr�I�"
8IU�T	��e��a�TБ���I�0��f�Ur(�MHS(YJ0%��A*�0QaSK�d$ĄW	*��/�a�k
9$,02m���T�Q����0����!ҩ�\�"ဖ�Lm(�(��i��!A"-5F�$�+�ȅ���I!�`m�Ct��0¤g�&�B�`m�A��ɣ4�h�A�� ���Ԇv�:���6���l� >��J}��<g;��>�h���UP�*-��]
^��@�N���jTiZs�<�%2⫮S�w��e�֋p���]��2oM�IA����#$N	(z��`�iE�cQ���,H�S���7�P�]�a����!Cֽ���t�:YM��-h�"<�#��<�X�{�j�'R�I$��,>�'=0^WΞ�p��K�n1��w��:F�5�*{q�LmDC۶tኸQ;0�c�pc�j�U���_Zrmlf:�6�T
8l�jMK���C)�-��v<��K(�M
$�E��Z2��4yJ�~�Q�=�Y�kZ�ڡ�l�K�kJ�?:U�Ur]]S�-h���Q�ad(<A�Y�e֝DqG��QO<�\����$I|o�ݹs���i$�A�2�H���)��M���aӥ����h4��HϞ}��BJ�0|_E4F��]�������VÊ���},�2r@�Q!"H!m�[b��i��:�\z'N�Ûon�c{"�f���8��P��[C3�H&z.]�-���5$�p�D����K�<8�t��;︕M���~���e,|��֡��3T��.}ί��8�p��SM2�/4�-�DyG]E<�O9^�k�w�UTٱ���gW�/��+�����4̬�a͍���=�}]���;��y�y>!�l�D%4)qSe�%� H��rؑX��+>�q[1Yd��tT�E#����K���-(<��#�㋋2n�Y���k����K8Y��ͥ�F��k�lpeC����8Q��=Q�r:�3�͓�a�it�;��ќ
 �i�y�QDG��u<�U�<���u��QX���1�=Mѱ�c)�'TN2�-p�,��KnyY��T��^ ��|)���L���I��,"TV��e��{s����c%��,Pė.�"b ��B}�X��+��՚B�"�%���$�	��I�Ċ��eA����)�$��$�3���,v��(u�A�:uMӠ�DG�hkV�,�vE�Q�ۿ׵����q_u��8ßmϳ�Xzw���N�]��wV.�$��4t�$h��''[��mE�l{�A�sY��	L��o��+X�C���"�Ff�8t���ϸ,`��ס�zxȩD&Yb�a)�\��bG��P�4��h��3�!�i��N�QAK�Z3W�y�WK���0��u쩃�)֙y�y�qG��x��uOo���;�Szֳ�U��m��'_%�jΝ8r��X>H�ƴR�ʫ��5������픘:|�!*�6��O�y��m����ȣ�%:̙G�>U�V�G��j,4B�&���c#��&���A����yG�F��)!P�`.���F��8b����嵁c"!�6]�6�p�ѣ�v�+�)Qҙ�\L¶oʊ/J"�QC�� ��@�e[!�P͍xgL!��f��x|Ec �'����~<Ckb�j�c��i��j�X�Z���Z�U��j�ao0���ڙZ3�c<6?6��&쇁��ͦxk� �3d%��DVx��0~g�-N-��^W�jyl"�����F[TR�hũ�[�E��ilEyN��p�U��[6��Ū�j�E[�3��_[iL��V�j�}n1j�-�~u�����y�����ñ�4K�?�:Q:x�<O�������D��O���Q�x~4Ū��U�j�u^�aձ�q�Z/B����x�P�4�1�{!<1��c<1����x�^xx?A���d��g�c�lEEEyי�Z��q�-T�-V��[alڼ��U�����qd����1�=c^M���$��3��>{�i�*��檽 ��1��4��<����>��_���{�'�qx�M��� ��r�1�N��'K5�$T(<V� ��$HE�L��1H��x������Ќ(�����6x�I[������~E�z{��_���
MC�n����E�3=rd�ofo���L�%�;���%������ s+����]�g��{������j��^���rI���ffd������z��U$��L��@fL����{���z�$��L��@<f�37��;�ꪪ�yO6�̼��[���<��:G�����}��{�.�t�h�D��@�\L�4jۆ�be� �a�膈��q�9X�0�l����n_�QCQ0�ց����w>�LKA��n���v�f�+�
�1��D[Tb`b�_��L��E�����}_���u1�"'ڗӡ�X~�&LX��E���\aJ�C&��������Y���ĸ11���щ���j�c�r���F�Z!�J��pFp�#�mZ�D�h�������G��itb4a��ف�dDm�ZV3��)*_#ckNJ�A'��z���K�7�e�̣���k|��qD{�#���68�1|�|0����l��ik[�<�μ��y�:��A��)��ɀ��w�$�H$��#�f.�9�v9��K|ltQ�DxL�"�!8R��ծ���s��e��<����iİ�a�8lN��K���F����֍�F�a� 1�c�(gxp�7����y�H�aa�l���Z<�%
 j?��h������>��H<0��p���6�����PxaѢ���7��h`��J�,��E����/=����9U��"c(l�A����Pa�F��Ã��A���G<C����=�1�:4�43������5c[S����H���"<�#����/��)�g{��2�d���P(L`���P	_��¸���YXB`�ͳ%U��"�$��`B(��4�fd	1�L"2Y2����W]T���G<�����JH|J����E!�S,[B��AND�B��A$@ @k�̐eY16�|b�S�l�:0��&��[(���\�#�b�r9:Xta��]6E^ϛy���-�m(�`�z��
ˆ�E�a��E��m5�a�F�nU����L�Ϣ�5�P��h�2��
5�V0�Ŵ���J4x��^x�x;I��8�)v���oF�(��=��3���8��#�?G��̉���Fm�A���������<0��ܽ��ZM#�sO�:����tj���G<�흾T��\Mw�ꢽ�ꬻ�&V5R��,��cI���m�+u�����wظ2נ�K����T[1+o��>����l���#���<t�ӁÇ�p�m�w�o�S��*x�Q�Oձ�7���u���t��H�@�_4��We�3�3C:3gO���������IX²�(Z>!�3��C~����F,�63��X��,hP�ᲅ�ae!�i�h�6�:�q�qaH(aϸ�����м�ƃL�������ѶRd!%2+)[L.ʪ.�U#L��Ç����:4]Cy0���&�M.���>���y�H��1y4�P�>L��V�����'Up$��B*V�$�ƕۦ�'.7t�VC7�%�13-2�Ѣ�銄��:�J!��ƇhaC��-c>��Jvҡ�C�p �4���Q�4�4r+�J�#8AQ>)#e��P�p�GA��AGx�6p��ƈ��":�yN����z��m[�7ɺ��*�®BHIF�dKɘ2�YH6��p��9!G�e��ex�WG���q8m�ډ�J��]#a��n$gXD����|�ԑBEH�cٵ����d<R�6@�SpM46}�b��0�	�#�!���4[GX���Tw^P��4��1P���0�8�M1���D�H�)�/(K�60���8զ}�E�A^�I��kH;���g�kF�1�v���>�ܷ.��W��zŗ��jfM��I�Ki����͸Q�YI3(��tb��}��P���}���B�6�Hy	��D4�&�QG����08ч"E��*���MC5��B��0�J�P���(�줩�3Ҩ�h31���,��(��m���DyG�<�V�=�2���M��gLx��:3�$�H$�@�q-����c�I1��3��y��H1��_F:�a������4����7�φ��u�c\�rl"��x�����$�eIڲ�1*ؒbG#d��\�Yh{�s��xgǊ%%���m��1|�"c^����pF5��3�C	la�vR��4��a�䌤�|3yM���m3�B0�C�P1�D"[�p1�<��p�7��bM�҇��0�pƢ\$8�ő/�"6ϕ*����f[>�I*�1��"�Mĺ2�RdCT�V��40�Ҵ�4lc�0/�H�Ң�Wf�q��F���0�������3L�g<�La��Chl��B���ɢ�&����s%,b�Y���+eն���"<���ǞS��0��A���=��RLdh$r."�I���M�:��%Dcd��?L�	;�/�.5���Q�F��bԨ*�Ƀ"��ڻ5��[S��8H��r�
nD�M ���q�c�C��!A�,|U ���\<6�2B2F��B&d��܂PP!��-A$A$��.6YM�(���q�EQM
�}��ɇ��(�6D|3��� T�l�([v���n��X3���m��a]$�w�c��ZA�%y�]�a�M���q"ccif��d&�\$x��x������d�j=P�ŸP�3忝X����#>�1��>M��7����^(�iX�C3�GU�hl��L��6|�6B�š��pV��(`�Z5A�n�k��
����cf�c@�����ޗ{�	��{ș��wװ���sp����-����C���(���qv��~*�D�i������8ꪯB���
F�4ǲDk�R83(��w}��c�J$P�h�ҋ��+*����P[SE!e�U��yO�q�8�/̼�����N�:p8pf��i����|q���lm�m��67��9�&�l��;�og�BHI3C��Z�.'�/�*>��)����xa�:��U��rT����k[TP�`���"��d���4=/���(NEky�aŤ�wY%�����Bőb4C.&f��f��׆bZo��Θ�e/o��5��/z�?`��(����>m�`�V��
��"����H�6�n��ck �� 2�!I鎂.G!L���n^�SfJ��^�-��Ӳ���tZ����7L�c�^����G���h"hc6���^!L�l���(O��6��0��߾�[�f�M+��tl��~S���(��?8��"#����F��~���E��BZ;�$�I�-0�o�[OE�ED��$O�v=u�Cґ|���&:�O�*CkJxt}Qe����+fK_�k�#p�J�(44i��]�T$E���6��4��B���P|���ǎ�NV2���[��唪�zrE�����T�m�P�1�'���/��xa��i��܆C�>���g��z&9f�+��/���84t�4ay��hy�a��.����yC�]L���m��e��.@�+Փ��w�|�uw���p5�A�DM��lz�ꪁ����#��H{N����������"�����مe�m�?8��"#��������'�x���C��k�~q�q�a�0׏�d7�Jr���Fuh�э�Z��	J�a�ƾ�Ϣk@�QQe����A���f���Q$y��"�5��2ZQ���(G ��8<��G�7+i��C\(���'L���g����:_�Y���aᅡ�u�<�Z�1�t�|V�80�d��WG�N7
\)�N���b=��ޓ������[Gǌ,���&P��-E��l����ᐬ6x����ˊ�C
Ok���Acf��#�uX�|��^lw�a�C΄)�y����"���.�{�|��#e��h�ƈ��ށ�4ʍ��"���|a�����c�v5�'���<x��1j�"��a�e�-�U��ձj�،1i��R*�h��a�c�mL��J��R�.��0���*�JZ���:�)m1���UjmKSkajql}juQyl"�W����х�F-_yV�-Ql"����؊y�4�)V�[[�q�R�j�E[�aT�ٵaL���j�mV�R�ajZ1j�+�c�u����N���i^SJaV�[V�ٵ-V����c�¬�el�Z[�q�[QV�����eձ��:�>"��:>!Ec�t5
>)|ByIyIyR{)yIOs�e�˃�k∾�?���2�����ңX��F<�<Ū���b�J�Z��-lZ��-ZZf��j����CG���:���k����m�A����H�k�/6N:�fǘ�T����P��W&}�ȁk�]^7�ވ��{P�K�.ߝ���k}^o�7�-w�zI����g����P]��I ��Dz���ɘ�ôF�8�Ηӽ�`iN�Cf�BE����U�#P�m�b`�*�fS�+ �5 �r��UrN�am�C�G�(02��)�;�d[�RC:>����1Ħ
�n���fH�#	i�D�l�����fi�5�Hi�~j%�Bp�B�Q�8^�ȬI�;n�BƟz�&
�A�%H�����Ί�<������ӢѤND��<��H����aC9h��q['�cC��6aAKw6:���3O�Wk�2�-l,��P���t��	��8��p��b��z.u�T��JotQE�E�H{�ڙAT'�Zel��"���H���6��
X�(W`�8`XqB��)��)�8�/��Q&����P�i7HP�[1+̅�`�6 dI�C蚎��%�j�+��D�Q�O؝-���-C%e*��	K.�Ԍ�.I�0�ih�ԒK*b��ݹ�:�h���
�45��s	��={Ez���E��_`�q���9��s� p�}��뛅�O~��:l5�w0U�C=��c@����]��oQ-Q۔<B\���%��,�w36�4��_HKý���<�Af�
(��M��%�rԍ��<��Qk�n�eN��3��#"YEd��(*�E�T]��4�(0��F=)�M��r��ZQ��c,t��l��"����L& J8XI	�"�B"<l�GX1���,�� 4���$c�S��I	�P�Di:��k���\ޞ]M\N�!^��$ù����=�t�L���y��$�䙜�١����$�$��l����=T�I�3,6f�r�W�Ɣx��SͲ�/<����DGQ��)ճ���|��z�u0ִ�Ac	D�jN�(jR�4��("Hm'L��0JlZ���	8AJ ��=7.i]ǔ�a�E<�u��hfa��1q(K�A$D�L���I�3����(��%�K�SI9 $ �f$�;���]-���F�Ҷ�#__Ň�
`����j`���b��:,ÇÁ[FS�˧
�6F��"�����C/��l�ZF�.�Ƙ�h}C ��>:,�A���f�1w��mq_p��g�]\�:l:0�[�3��|aH����۔>�KF��]X���6�ҕ��)h���tm[��8�0�y��2��|��ӌ��Ļ�(*?{�ɡ�>[?/	�QKDw"G[��I��"�I˕�]X<�x���k���ύ�e�"�F}�� ���(8{�-Qc���}�F�R5è᭨SS����m�e�~[�DyG�<�Vl
�Cg*���j�=Q���Ő�����1�B�[�l�V��N8�8�80��;��7XZ��J�80 �2p�>:b�c[4Z�R��ц��,����ya+ه� ޸�:0)�����S�gF��:'á��F#p+E1ͻM���n����=�x�h�4�08u|���7�H�O�"�ძ�}�G��2J��"ZUvBe}�\�hE c2'��q7/M�"(�V������}8\6R�[���ǴM.ac�rde^sT9(�z[[�Aх0�D�Ȉ��%���<Wq����9Z���h��#�(í��˯6���G��x��.�A˱7^����y��ժ;NQ�8�0c�C�����-��&����������A���t�j� �p�j��[��qզ�0���7ɫ��V'�+Fc)`Q���,
���Cx��̤�k��D���+a)8끨d��Y�h�m�m��t�����N�
EY�ypf%���*��*Q���c-xn��̩n�cF�`�5�&r��gU�y�8�}8��\4�������x�l���7��aх�#�#|Z��E��#� xa̭v���9����&wi�}��h���0�2ːmD�Ax0�D8ag�:[o��-�Du<�c5�+:y�����!�QE@@��4��0��v�����VtȎ-�b�o��;�׍�y���kG�*�J��JdvV�LT�p�H*i�#���yd�aT�x�\_G���g�*�TE�6=�`�^pW�x?��3���'��ͽ+�K4��y0���:���m����h���:b�0��"9��Q_>�&K����ZFˁ��L<5�5���-s��Zp�[eQ��Z��w�=�x��i@��]UU�/��G��)��uc��4Uaj�wcv��8Ptacx�)am`���l��&4�(�DZl0a���kC�`�'���Z�7"���FQ�2�m��ŭDGQ��)�c��C}�(�K���!���R.:ai/,��ے,����;$��B��� T��ȆHg;/4�i�����nMrd��&&	V�������CI�W���!q����n$��$�H�HDQ��W#do�XI ��j&�qp�#-�Z��QEQDX�`L��(��j�+%��^���4�{ǋ)��g�{����� �kI��E�li:L�촋楖�C������1����$V�*1�'C������m\pnH� ݌�HfDi_�8Xha���j��G��8x�/�y��m�ٳH�a��-*��p�����L���Z�x6���<�>J��h�C������X�1�sz$�+Q��9J�F�Q�5�%^�w�\s�n���1q�G�BڂB����� k�ZF�R�3���i�%��KU�ܦ0c־c�\G���q��:��m#O-�~qkG��:p8pf�,�!v�Q[/uI�S#)���%�76��t�c櫵���޼s�/\�8�8�0y�UXiY̢��@�Z���XthR�+z4��q���]N%��`��0�C��Ե�O/6�>;kA���J��5��q�)#�{GJCŲ �PÝ���Z��>٢͛)�Y��$ұ�t��F�q��x2 ��`4)�͗�^��Ռ�"Z�� ~��ዮ�A!�D��h�S�.�Ƥ
)w�w�RBn��|�_7�O�Z�b�����r�cC*�0�%)���A����k�Gv����̴DEї�"��`O�:C
8DE��u3�U-H:(z���b�GHQCV�i�i����֏"#����F���߾^��A�d��w�`#�t�q�A�֟��l�]�To��Ø��o���դ�0a��KV���#
%��3�+g�80�xӈ�{�J���j-����1|5�>j�<PHh�ha����[f��4`q�$��6�!�&'A��%�Ճb�CU��w���y���x|ZZP�z�v�Z�"�ˢ8�R��j�2qZ� ã@�DZ��hU}m� ��r�*�B8�	7 ���3��Cs5>�w�A�EG g��趶�G���Ո��V���`tapq�6Xƚeö������m���HWH��������2�o_c'�[J~im#O�ͣ�Z<���ǞS����3�⽮۞ϼ�}���8�0�0����"��8C��!:S�N�Z� �m�z�6����\��_���c��w�އ�e!ƬGx�(�P�0�|�c%��Ϫv�-������Kd�m�ƣd�	^m@�͈�I,��CKepцȢ6�����M�t����mO��.!��B��[6M�jM�5�ʆ�M��c{��^Ɨ��~�D���.�QmE��m��7�I�xi��Fq&��n��5�>�)��TU�HS�:0���Ԩ���eRG�"!��4P�K
(mm�����	��3�"�T��C�V3C<�
[l�Egu�}D�
��,�l���c��?"��y��ym��Z<���ǞS��w.Lk�*�Ղ�{\)�\@�P�N���$)bڹ�7ȍ��)OuJYl�2A%�k@F�r`y��*E�@�?e���-C
&�A�L|"��,I,�$-A	h�!i���t��(��"��r4Y⛘�V���z�oh�dQ5� ��!)/|�:݁���8/l�!�����hi�#\<D��>���i�k�!�ta}Pθ��� C�!�M��P��2��C,��|248�8.�>��S�Y�*X_�:R�h,c���߮�\til����RR�QC�FΘs�s�ccŝ����>.#��)��:�Y�-���h��*��P¶mQ��A�ȏ��F}�8��0�WA�8��UW-r�cQ�D�deʪ�U%B�\V�S�0�P���Ԣ��(�<���mu����*�O������0�����&,83��Ӎ:��ߜZ��Du<�T�8�����6�c`�q��� �'��
�/?t�EQE"�3�f�����`�{2�EV?4�+\��ysc�}�S�(��D��e|k�i��X�YE�aᆏ�����>��xg�e��r�U�k�}��C��j��8ܬ�.�:Z��'ǌ/��0cq
׋G�Ĵi�F��7����6�h��d�W8=E�pV���6d�pa\�sPn�|E6�t���K�z4��ިyK�p<0Nΐ�[A�q4hT+�j��(��U�R��e[E���Cd<Dס��kL�����)haz�ۘZ!���G$�ZTA�x�vPta�P�"z���i"'��dha>����lo
��U��.����6��X���xd�6QQ`�ֆ��,����+�*�Kaj�qV�mV�y�U�-�p�R�ŶŴ�mV���*�l"�V�"��i�)�eVR�x�lkͦx�D���3�<6j��Җ�il-M�����ԵuKWUj��[(���F�Z����KTY�[��g/1�mV�U���V�U�Ū�kan�©lZ��0���-V���j[�Z��[N-��\��<��Î�g��{.6��6x�<J<O�����eE[laV[�-�-�R�[6���R�ǕjEulqZm�U[*�Q�P�~,�(����0���A�6��Kܤ��(������<��xx?x�lg���Ұ~C�q���Ū*#��l~m�+�lZ���Z�\[�LUZ��V�eN��^��t���'�y�O:���T~>����G�)�F��!$LpȢ~���7;>~%�AԪ
,l���u�	���A�}�}��E�f�FEm�	de2��iwQ^�Im��Zf�#��6�5ǧya�)���'MevcX2EުI�!ΐ4�<p�y����RD���#O++�%� ?!�uzWz}��f�kCa��ƴЛ\h4Ѧ8�����Y��uӎB�+����6�=4S�r�m��Mc-��ʸKPg��F��ZF��J«bB���!�۾�~=��eܻ���������{W���۫:��e�}xO9.�V��U�ek�W�W]����݆��м����$��fXl�E�.��NI�`�pt^r�.��NI�`�pt]��n��j�R�j�]J��O<���֏"#����k	�S�-��&�{�`��aEQIp @c���5�ajʥ��f��qL?;E:��րct������v��@�5l~�:�;j�ٮc1���n�X�f�]�n蜋c�Gɭ��":j�42�00e�[�8O�;����H��R�l�rK�j՛6��d8��"��!r'�(�����6V���1h��?HUS\ѡ�6JC��QQ_p���-h������y�-k�"3������٣h��x���C�6FJ��F�R�WUF�h�i3��a���P\Xy�E��4.py�iX���J���E��e��k��l�l�Yn���J~q���帷��y������F�қ����,p���)	!$D�\rB��XܣJ����u���De=J�Z(��X�5��8r��]"9�[-�tf��Q�]������ s7�~��oH��V!�e�9�-��E��l�C���[aVZj�\"6n���Pѡ��?��ƝÛsվky���0��j�ݞ4p�K3Zq.c'"-��AC��kd���2"�t����$�9-��6uz�������/G��jх"�9}mf�RH����aя��k�2��EK�<7aѥ�)��q(��Qh���Z��(Pf{rHq�}9�h�"���D�il)�a�Yiy�ſ8���Du���]�'���$1B<��8�[�:���)�$�E�%VD�QU��I؉��!Ll�_@�&��m���[PO()�R���C�-c&(�W�����LG���1�(¡���*H�I��L!H�ƌ�D	0@"��A$A%���ɘ��)�16�HDc�Ea��*GxloVZgF���_R��x�f&7_74}�G���^��$c*Tm�;
2��`Ή�mi3�g� R�����F5���-?>*�8�)tc"��5�"���g~6t���Db����i�+�}8PQ������GJ�S-yH15����M�wF�0��ڡ|3CGǍ�c��J]��_A������x��ﬄ=�.p�)M6�8�hg0��G该�(b0�	dء����f<cM�{A��"�q�����D꣑��P��Xh�<v��k#l�<1��H�CMH
a�u�e��8��V���GN��i�f�	J�r+�հc/"����{�a�+`�V�-���mv�q��Wt��Wt�m���fu�@[̅�j�7Y1�m"���E\��4��r����TGس�]�ؐI�Ip F��8t��}u�w��o_<i�\�!�Ծ����-�<����C��Ս��qxs8�5P��(�����e��(���k�wLq�d�G�~�G8L��mł%�&�E��J"C�E�a��!���H�
Q%����[`�	D�)��4
mJ0$k��i͇2V�ڹP���G�`@Z�e���e	[	������C3��X<�F�[(��i2k�rQ���t�B�x��dq��<�q����3��QB#�tpނ�aD_|7�!���TGFf��~�Ϊ]�FC4�-"���hn8U�H��#%&i.6>Y)#xۢ�I�����̍�>>��٢�/^m�%�c!�!���~�J�����Yѥ�d)�L�QIl6�A��#���-oJ<C���m��U��?)��a�y��G�~[�Z�h��ǞS�޻�n��[l6r(��S~Π�	 ��@���E���65�D!FA00��ܤC:v�F�HP҇9ܣ师3C�3DF�2�(��:����8},���[eif!�!c0�4�+ڣCC�l��1��o���&���E�b�e�BP����*:(�h4al�4eh8ű�1e���/�,��c4�/��S�l�_D1�y��|i/ ϼC�ѢQl�F�"ƕRhlԊ��=F�x�gyH�ٙUUT������E���u��g�}H0f�
EP����\j*!�矽
��a�u�>�c9��cE&i�y���=��Z��Q,�(��?-խh�GQ��)�o�n�-̐�.�BHI	" ɶ�|��p�l�cG���Ư�D�ip�%�{���V3(���3�DE:3�ܜ�nK�H����
��	!�0NQ|3��t�Pǰ|���%ѥі3�J,�!у�܉�&/��u��>8��у7<d�'0�&�hh0f��|�i�_Vko�ʜ�<����¾�
�h����,�����3c�Q��� �4y�s�B���*�uj0���������9��u�=-#^42��1{P ���E�w�C��A�uZ��=� ���і6�(����J$tgƎ�H�dh�CF{�?�mW�S�e�u�u����Z֋Z:�yN����T�NV+��1�|G��2?VEGL&m�D2�a�(��b]I�J�
A�A	�N$����VL�O4aF���9B�	nEqϥ��=� ��(���Se#�b��4�iNP����I�:�Y�Af@r(R��Q"EtJ*��`�˩RVQ1��K�-��U��dM߮���Apiq�M(ɺӲca��GCD�c���e4o��ihh��biY��հ��e��m�.P�iB�p��0|��W
��鷉X��;�[T��)�~)�i��p��k�Z]4`׮��S�]�^�8�82�9�uk
��_�i�UJ1N.�Q�63cV�#옿$�l�I�<B�� �b���H����f�����M������<:( ҃>]0��#p�o�)���y�?^>,�2È�2��\~~ukZ-h�<y�:η�9X�1_s��f��3�l�Q��:c�ݣ�_���$���"��@�i��1�DP�D0b��?6߱��3∌=�d���F�\��(2�8�	��5����ɒSr�Sm���i�gOc~�hf��[��#ƌ<v��:A�D�9҃C>�gdK�l�tcG:4��иA��_�s�隿=��Mu�o��w�Տ��*�@�f5�X�\~����^@��R��DR3��*c〴���� cy�p�c=��ƍ#t|P�2��~�.�kdJ�[�#*�h�(�Kk�U
��C<,[^>(��f���� ʡ�u�;����^=FK0�T�N4�-n8��V��֎����F�U����Z_���(�lm�ǫ��V���$$��c��x���ח[������G0�K�9C����h�[Z(62��+|�U3'��F����:8i89����ѳ0����}E#��Ou�m��"!��~�|ݔ���*F�YJq$NH�����:6�Ƅ`���t�K�#���aGOa�G1m�64��֨�b:6}�V#�y�b��t+����6׎#�>��C9�Ld:|p������m��7��hc0��Z0�.,����ѤC���+O��0d��i斷�ukZ<tٰٱ�:n�R��U�V�+�HI	!$DjDwvG(Pd,�Z3�(i����~�i4�V���d�TF&���E�$�jC�m0����a��AeB��-�3Gɭ&��N-��1Q��P��ރE����A��Ȃ�z�ݟ#��$ �h٥H�Ӵ1��}0������}�9����nO�+cxZ8lg�,�7>0����FR���-O�^g��pܝ\�A�;�����6�p��"����{g�0���WǋǇ��Ӳz):t��OE���,���>���d'��Ūټ�1j�Z��-x�1��J�[Zض��V�y�����j��[�8�Wa�aVR�JYK+�Mx��l��xg�C,v?¾��Z�U�n1��j�N����SʵR���<�>�b��E��Z�V�[�Z1ט��U��՛V:�ql�lZ��)j�Z��e�U-�*ԵmV�R�b�jE��h����|"��p�fA�*�u�V�Ū�kc�b�J�cj�ؼUb�j�ص��ͩ�EZ��:���Y�0�%���x�Ã�� ���3�c::R�JyL)jZ��V�6�W֬�Ũ����+�U��ձj�<�||N��c���	����▨��U�Ëc��q_h���YK)j�}j�,����0���F�A��$@�̈́�/ڸf���FK!M�D(��7X�0�:uvD��2�D��_���64U�p"y�j�fJ!���1���I�k%dvR�����B�l��D0åF��a�ٸ��.�9B,���Xw��I�y4��5(�ZE�8��{�\����kv�I'f�9E�nJҥ���#(����L��A��L�:��e.vGփI:���'�bB�ĳDX��j�2J��f �!)c�	�Ɔ#���3��=��vv!������Im�N%a��I;
����:m��K�:j��"h=��T`�4ԭ�-�%�a�l�0��UcIGSh@x�p%$�XX�.٢Bw 4c5��PH�8X�f*����	e	茏d",0�J/���I^^��Y�7$C�H�,�[�f�)*���%���R	�1���p�&�B�:X&�
0�'N0T\aP�E+�Br�"x�7(JRPK�g
?-�c��jf3�c=��C����w��*\��^8g�u����FZN�l�8� �JOS��:�~�"K�3R}���Z�$��:S+�g_	`���G�¼����LB�E�����)��ɈK�D���P�Z��[d���R(���.j�$P�*1������p�hdX����,�Ɍ8x�hDIddNlA�'�.=�!lM�$��
H�f?&d�N8"�@�S�Ӹ���$�`�K�6�c��\e�T�W��w����߯7������`��˼ܒI;������.�rI$�fl�y���$����8�fkZ�^>x��y��y��mŭ՞<t���͆͌��6��T�Y���HA�A-:��<�FM��.+F��� A�҈��e��.�а�I�0ڡ!�~b���y�^N�|��2�P�!�$�-ePR.�ړ%t�f�w��I�L�-�%q���E��,�BY�"�h�gvNH���@�ɱ�th�����$$��Ѽ�������m�\G��� P�Y[g�p�p���4R���P�&�����(V��z}�	$(�F�����^R�����"l}0�L�Z��<,�C����3c�t5��Ob:0��(����f�-f@�7�f�o��#L��4d�)�W}�Y��h�JuF�o��Y�X�Z4]/�3�\.�ͦ2HD&9w��yG�1im:���:�V��ַ]:���6��Kq���h$�H$�!�5�G���7�u��#�|w���T0c8M��S��Za��g�,�-X��1i`Ə���#�鿛�3iA�S��Lv�(��Ä_,����µ�����[U���RV�4�Khh���E1+���m��tS�Y>��l�ɖ]�n�S��g~�h�e�~�h#0���/:3�d���c���;Z�� �YI�"[G�//0fU�8��)EC�/���ӽ��Y�g�{�x�3FJ:sA��-l�ʑ�i֑m�:��ִZ���xxOM�^�)[ל���+�,�+Uy�T��Ǵ轮I��Q����p���p�BH�3��ih�=��ZD*������m&3�'��������4p1����C�{�"$q�A�o����t�hPd��è��E�)K2����یg���d2�2�A����F���.A����X��(���◆|�H1�=�M{FՌ��'��HQ��"��8PP�*$J���ƺZ��%ѕ���C#�e�kGq����u�V8ZcE�[n�������62���D'7�_B�8��$Æ�l�Ŝ,���պ������T�������5[��[���[��I	!$D�G��ii1�d�R�X���j�҃C/��ԓ��M�ڵ�kK��pg+~���̓����:�J �B�
l�)��]S����	��񵁊�ql��ݚA��:�ǆaMkx>(�l���L彍`1�0q�rL=�]=� xf�T��z��wuE;��M����Q��D^��N߸ꮯA�mx����^<�lt��ewY���o5���󧆟�|Q���jΚ;��kZKC%\���g3}|�������E�6����xf�n��:4kd4b�Q��2�6Y��0�պ������T����gU��5Ƙ$���"�[Y����"T� Q�QP
���"���}�[�4�D�	@�]���(@�$BIRȬ19K62[W(��W	%3!L&�J4���	`��.�*�#�-U|�	!$$����SLNxԌ����#)_��lQ��_q�A��XV�k�����S�=OMldd�b�a�)3CL��|w��Ip��Z)Zc=�ҍ�iy��Y�ݱ�Ϛ�;D�7kA��_�\(��>�sP�c(ZM|���8>[ZZ(�C/�Zo���Yֹ���`#������G���F�R#m"� �Xe1[j	!q� �>0�o��6�q8����#��۪ç4a�<ӭ#O<��uk<t���͆͌��f�T��nBHIn���c|6�X���7���dZ>]��F����a�����A����E�M����'��'c�n?||3�&��ly����1�1@ctA���3t��f��m}�Z2�9Tr��s�y�V�3��y��Ʃu��.����*��܄
(��[u����!#���a��б�g�u4Z�;�6o��� Bϗ���_��c��7�4?+;�¡�������)����#�ᆑ�)�#4(Xϋ0���>0��:������T�:W�ǩ���H�U��7R�q�gOonWKI>�����)�,��S�~�BHI	" �Sb��m�N�vQծ#���dj4�<<���"��Vx�P`�1{(�G��m?CzmA��xg��R4,�c,���|�x���M����Bu'	Q `�2~����}�o�p⵰�����4y��
\\o�����C9�z)]5���6��BE�ZH�a�[���.����*+7��yϔd�tx���U�`�a�Ǘ|6qqN�jjA�42��C∍�>6ae�#ji��q���"���ִZ��M��)V!ԓ�71���_�A(I	" Ν�G�5Ӈ�m�n��V�[�2��2��i����:�4�_�����"�X�>/fTM,h�r$��fĻ��Ru��pP�;}�hg�kj�E��������h�+ŭ�3��J��1.�/�	���eH�B�	o��g�!���0}��uhfh�գ�S��P�4p�}w�/�E�,��t�1�4Z�l8�-{���Ν`�zϸ����k~��o|�}O����G��T(f�e��G�\~ukZ-h�]S�ԎCR!*�x��w�w"�1Zim��q�N�X�i�dAF*���LQ�rj���o
$�IL�����T�V�d-��1�O�T�Ȑ�����N���T}3�L*�`���`�Ԑ�Da�@CI2���H$�K�,":��7�$�I��e2�'d4gL+4R��A�f�ֺi{*1��g;�����B���֗L=�a��QCX���"���e�އE�Z
����Zt����6|��պ�Fm�0��5��K������g��7##{�u��j1l(g��b��޼1\4B�A�g����U(I��U�Y[.$M�r�n�:!��5�+��M�lLg~��E�W���ܗ-���߯���uM0�YmZ#�uխh�����Xq}߰�Vy�k��ޮe�ks�u�vBHI3�F?�~:p(c�m�f�Q��g/݇��1�2-��Vf^��Z7`��m�.g=�
�c4�����}ru�q�{.i`3�:3��{43]0Ԛ|6��o`�W�O��{�Y��Tra&@�@�2@�H�A0o?wH��l���z6b����p���ظ�����tmzR:16���7�/&�����C8��#���UH�	�t����t�̘`�Xa�y��~im2�T��DGQe�DF��#Ȉ����m0�!B��a��F��i�G�uC��<�#��<�#ȏ#θ�E:��(�"#�!�"2����G���FQ�ѷ[m�!De�GYB"��FѤq�<��h�6�QaFaJB�!�"2�F�e�ZF^y��yo<����Z��ikZ�Z�kZ:�6���!C�?z*����1��z����-ŀiQ�=�_4��S�D-�|�����P�!�*�B>��BW���y�i@����Uc,�!�����G��[T\D.C��c$ء-!Fc�u��b&�d��%`nWLթcp�~�
4�k`�y���9���Ժ4�T86s�"�oغds��ǔ/[�u�ޏ����]H_oquGӱ����곗ߕ��uk�;�e|
�˞y��{�a����RI$�fl��w��ԒI;���a����RI$�ftI$�2I5�kV����u��iխպ�ִZ��]S�8����z�zw>���<�J�O��w߫A$A%��#��nC��D1�le�ţ�0�Yh�f�).�422�s�[G|�h�Dl:`A��՗�U��z��"��<�Nc�>Y����cx�j��4��6C��R<����pΪ�Q�&�������x���Ct+(k��0�4|��i����}Z����A}{�uA�|x��Y����Q�AD������}	�YE��2 ���
q��O�~m����F[y����:�ִZ��]S�8���M�*���BHI��m��3F揾ٱ�̭G(��]m�3��C ��i���?��!�/#&:���xgՏ��p��3��Jڵ��ԏeb�3�1���P��C�}��#
����8��{f�ZĨT��Q�eE����5\��GFpQi���cU����j�Gt�Mwg�K뫫wUW�?.of�Vl�f�CG�g�p�
83a�-�Ө�V�Z�kG]uN��`���k�A�F��8�&"`a��H[HD�������UC��J���"H�	e��(#&B-XN/ҧ_ u��h�	A� U���|vAE��q8Ɗ�R�ҁH@K� A����!��	h�۷r�E8:e��ϯВBH�0����D���)�L��!���£�qr�uØ�p�f}u�w����15�d#3~��=��}��~���K��#��ÃD(�E�*����˒��h���L�� �k�(֏l������Yf ���t��3�c�����������m�Â���^c��|0�����b0�og�I� ����F�]hR�|r���m��=}Ѳ�ͨl���H��k�"�Q�F����*�Mk0�Ji��-��?-��]Z֋Z6l�͐��=z�����$���""Ҵ�fϰ��M�3��ƺ�'�6����xz�{�B����̼n"Z��ٳ��1[�p�,�������.:<I�H`p����㇈%ԗS\E���:2��^�p�!���R�*���j��6mGN��gM8qΣ-.~�w�Ϻm9�߷[]3
.�X�2�L	T�Dh�yx�p��5Шz��������9#)�CgK
��[��ᡑY���Z4�)�B�t���7Vof��������GYmD[�κ���ǎ�6lf�h�7������
{�S�Llm�m�1�8�ܡ���i��,�Z���r���I	!$D:h�dTR2^�4C"�2�m-@ֈQ��qH�m���=w'�ڳ���u��_u������m�N�� gWqɗ5N��m�G�s��Y9�9�L��r�I�JHAڍĄq�-��ݻdiѽl�p�kjx�oj��������4Z����h����b6:=Mڎ�?�p��X����ќ,�6�X��d=��)����[b�͏��M��x��K��3��|�f�l�W���ex�8�Xy�QƝE���Z�kG[63d4�y����ثy�i�����DB+6Q��a�7�k����F<C:ib���U�������R�F�d�D7\��>�����O�2�/�sM�T7�
:n����u5��xP��](�2�M
0x�0�è��Xl��X3:M{�%'�g1�IX�5��~[0�Z�7ť�E* 3�mv2�Ƿ$(�Ã�p�4l�AEt�8Z����,)��e�uո�ַ����F�4!��\��O�q�ԑ�0�Q��*&#���qĢ#��Qk���M ��$#
*Y+bm�GHf@�6�Z*����j��Cbp���N@�f�*�KE@Ă`�Y-5$m��	8",H����I�Ӎ���r9�m Xq�I��c�Zٝ�8�p�=c��o��.7��cm�5\���s���Ur���:���X�l�����U_s�~>t�kd6k��Jx�qs���0fϙhh��_z���63��6Z�Մj����3�X����H���/k�b��sƍq��l!�!��x��g�u�MW�P��`˙f4A���qD�! ��08xM�!e��8mE����4m[��)�f�Bܨ�N9M�Z<�3�6p���[��έ��y�T�/�T<�R'G��I	!$D;v����ܒ�<h���}��Y�zƸ>�q����aغ������ԣ�*��xt��z���t2�u�%�lm��5�e�ʰf=G�e�́�c�#��At����f�4��f�p��!��a���y�ǌ-�j��>#�߾j��7G88�-Q.��cL���/X��(d�_�Q���
�=��dw!(�M�w�1�#��-)�u��i矝[�ykE�y�:ß]}J���_Uf�4�0�g*1��m>0���7���c�����I� 0�#�,��~����,�Z������C���f��>G�zZ3F�>>��e����ki���C�i�[���p�S���ko����g�t�BC]4��F�� o�xd�U�F _�l�	��E;�.U;�I�rݐ��a�C�n&
��*:l6}��e1�No��{m�q�x՞G��F*(��Y�i���슟Y�;�W_I%3�n��T���Hߺ��<��7U]��)n�M)iPX�+��2b�I�������Ä:5Fό:qh��e�?�0(�B���2�4�?:���Z�kG�63d4z��:Ꜽ��BHI	"!h��yq��*��*1�\�����|t�O�Q�Y[Ñ�㰬��I#�
�`�
�����̭"�R�*���	���Ea���`>��N=e�a�'l��ғ6��t��Rj�~���_B+:��4�0�����E8h"��(��ڡ����Fg۪ѥ��v���}17�(T@��h�ip��7�����KG�(ᇚ�*O��氛Zf����>z�p�gg���[ao�}��E6�X~R�i��m�����S�DFQ�u�")DGDDu�y�q�!R�!ye�iF�DqGQ�yN���#��:�""<�:��B<�����:���H�����FQ�i�Ґ�"2���#��H��Ȥq�Di�qF��:�(�0�iHB�B�E#H�2��-0묺먏-o2�֥�m-�G�kZ�qm��XY��B���]�j�ݳ�cp&�j�	�bT�y!��T�#+20�D?6�T����8��]�eP����1��#�Ƴ(�<�#s����1�����-����lx�>zqU���$Aa&�c��,�,pi��j,�)\O�H�\d�U�@��,����KBC*�+n`U�xJD��	,-���FN&݊r�!D_�ґJ'�ӖT�"C��6Х��	�jY !�B�!�h�&8�A�
� �G���ؕg�P�,c��9�O�TFx�O]Сt�vYS6��%e��Ǵ���k�i�7b��;�W\�w7ul�@]h��WwP�������j�r�TU ʾ�
�s[s*�_8a��	�	(M�8t\.m��a(K�X��n���p��ɲ��q�%�#@�����%1!I{^cT�H2q�[��3~3�6��,$�H��S�|�B�JH�p&K��3:�A7琈�w�Ts���B�cS�P�O��$%,S,���1�SE�"�@�l��.\�	f"�'�F(���O!0za3;W��7[����ی���m�:���h�S��~�#XEn[ԥc�r8KO#p�eG͜�96��Bg�5'T�Y��'
����K��1�cxAX��s�q(�h��v������H,��7���F$�F��B�H����HB�br�-���淨�K$ҁl�S��j�
2��
�i��p �M����l�H�cv$�!Ԣ�D[����0d8cm@Q����j�{�}k�}<�1<g@;���jI$��΀v6���ԒI'�� �lww��$�L����$ֵ�_κ�Xu�]e�V�V��Z�kG�uN��y�y��k�{Y�L�F\aX�_"�J	𖺰�$B��TmB�Z:܆ȃ� %��"hBT��k���nWl��T��K���+�58�r�Iq�Nd�QR<5��$���"q鲞��U��$�	�nAY�x���b�cm�a��uKFՏg͹7EVpf��qfh�T7��AkƖ��1��{7p��(��z��D��1�~[_D�}q��ɜA-�;�F�����ߡN��1Q��Mb1|PQ�K���,0⣔�I��[6��G�PϏ���TiA�pEy�(�Yka�MIJ��?%��
��M�6�s���Rz=���y��S�͆�t�󧛜m��áf�a��YF\~~~ukyխ�u�T����c�u�$���"rn��ў�ٲU�
7�E�-���}��E�0�p�a�s�O<o�7kF�!�U�5嵱���8� ��`����0�a�hm�݁�W�x��^G_#
:|ƙf�~�e�'��/!�u�O�}�憚�F0���G~��J0��0�(�����/�qT�K�b齕cF>:@�ώh�KJ�|JG��6}�u�A��������ti�ˆ�Q]o67M��#Fp�g���iju����㨎�-�V�Z�םS�8���W�o)_U��Lq�P�[�ޏr�$$��k�2��<�������&t���g��׋�E��3AG)�98��;)�܄�F��a���YkӨ{���p���ۘ��������,cm���s1�����e@+a�,����Ad�lݔ��Z5s�a��o���5F�8�ٜ�q��m��\����h�������lM��i4tgoڢ���4䦬�ƼO)��SΙ->u���_8�֮iT`���#a��u�[���zvf2����#.�eL�ی�������Z-h�Ω�nS���U�1�#l���^kn;N��+=2BHI/�F{����aӤ�[��e}��>q��ˊ|y>G�
9r�7���4QI0���MM�!-&�~���׾v���
�0�gL4��Fʃ���H�5~I����Cc�ن�䎭��a���H����UU�E��=��!����gG�<�]���|���~�!�Ӧ~����ߜx�ҩ��`3��	�4SQ�Pt�`�Šk��GT[F�>�Â�Y(�Fμ�����Z-h��)�Ea�&�x	%��&S!FK~r1�Ph��$;c�
mB�9bK��8Ҫ���@6�11E��\���I��f�"0�J"T*S��(�eM�T�8@�"B#����D|g�2��#�����$�H$��V�HK�yS�F�bG�!GC�45�T4W�q,,�4Y�{��Η��zTꡞ��UC�^w�I����PYE��=�<?&�g�p�=�q8g=[i�(]Z1�'�Ǔ�*�/�\�hѢ�p�GL<`14ϸr�����A�j�6�<փ6��?zI��6y|lc�S/A��V�����U���]|sэ��٘���b�Y��<%�#$��Fn���i��b����,��,&�����;����e�2�Ke[�#�[�uh���<�Xq��8���ϰ��뺨I	!$D:}�4���6w�l�$�H��V��
8�_p�lj.�7���c��áFu�8t�4��^n��G���2��h�4��?p0�c��Qc�o��5��k���DC[4o~��yj��T(N�� O���5#ʻ��]�hlv�CcS��Z�ΓK��QF�����gA֊6mp�VmV�1�
G؈���o���3f5���4w�ñʒ�(ëo=�j�C�a�<ï̸���ο-庴Z�מS�8�7}�7�_���wv�o'��$$�����]�m��r{#����2���n�lхo�*��/�Çx�_u}�W��p,�v�Vbd88��<3۩���Ԅ�"H��l	7"$���b��|�l�3#<A�\��c���]E(`%AA���<n�BpJO/>��.��)�J7q�j�Q�c��%DG���ڴ�*�Kąq����6܍����udB�$�d1�m$���[!J %�t�%8��,4��Q0�#\a�	��x؁dDTL$�bS	d	".1(>��^~�s��:���m���٪_h���]��E�ŢS|1j�w�4p��V��f]S,4��̺�?:����N�<t�Ã8CE���f�8��F��Wuw�DA��0��Ǧ�bc#�5P06�F	�-��[�E8�ȔaM9-�1Pj�aY l����;am+i%ul#�1�*��	<��Pʡ��A$���=��Gcc�##�ʦe�҄��	S���p4p�3Ƶ������U�Ch �`��*�i\�Q�M�N��,���ua��E-3�>�9Ìl�����g�k��h��Z�⫼��W;1]���նѴ3C�3����aFK̴�K�8W��y��GU8`h�z���<��B�CL4�f�3
9���|\��:N�gy�՜6Y�D,�_�~[������-h��)��:	֌�E� ��xj��'i�#	��E�����[	��4��9y���F`P�5Hv��X�v:E��	d���I@�B�Λ}�K@w�g[56��b��"H�E��`�,�$$T��eV���PI�Ip!R�DCJ2[-m;���I��b݉�a��ƾ�C��s���{���(a��I�l"8R��XA�/6�5ĸx����L)vYfl"�l}0�lڭ��[1���;UR�og���Ԍ������������g�OԮ�ל{��/<��T��/�-���Io[Y���9����t��E?c���~X�f��&Mԧx5�Ì������kI������.��G������}F�h�À�iM��̿2��:����Qk:l���!�����P�N�ky{yG��I	!$D,��6:�4�W�Ct1�������Q��4Cae��٣�͛K�>�M�E~]oC��E5Լ�������f��PQՄ�&j�d}�0�ױ��VW�lk��\��/�Á��_�P@� ��
��E�]�d�mt H�y�Fќ�0f�|>�5_n�)�*�����|A�=7��Q��%�S�����IT����=>O����p��aי~i��~uŶ�8��DDya�DF��G�mF�FTB��#h�F��i�G�U�uG����eG��DG�G[aH��(DF�e��2�#��G�DGQ�iF��Q�X")�F��u�")DGDyF�u�mH�l���
F�*��!�Dd��H�2��M0�:먏"�ee�KZ�Z��G�m��i��ʖYe���ϳ����3��� �c���H���N��yOJ9�{�+�!�/��"X?v�A{ɐ�b����l��K<��qs5^VĘ�9!��)�6���Tì���O�ǿ�o�1t�d&��26�a���ϚE�<w2�5(�q�t���e��[��m��gh��a��WU�k��I>��`ڭD�}-���L�������v�~��{��m3M��.���aL���l��v���Z��{ q�tm�c�O�t��FO�'�g���˺ʽ�у���b!�i�������}��?�=��z�j��u�}�2&hà]��*I$�&hà]��*I$�&hà]��*I$�1@ֵ�Y�T묺˭:���������|<4ttа�q�����
��*�)Ϯ��	 ��#`�����S��2��Pǯ���j�>,"��4|��6�E����[�1�r����<Qa��۹���.�t����C���%HR�<��3C�a0�\J,�3�0�e�HE�����<�������>6��xg�Xv��4p͢eԆ�<oF���烑��a�Ċ��a���������]���o��LkHO�a�_�/�}�:�����AQ�1wl�}:޻E�x�;����RQ \��M�t�4;�'����0�����G�H璲�t��(�f�>6����QkG^yO8˥UJ��fD�~�6�>I��7�)Ԯ�m����a�q��	!$$��n�,Ჸ{N6�UC��8���%v}���a���E�z�<Qy�t��i��ۑ�$e��'DB�q#�Z�QD��h�,�u�1�������4h��~oͶ�l��.4EX��l���gG�{n�U���n��(�>5��Ó�a�ڑ8�*5��)��|ϊ���Y���"+�õ�T�)��E*6Ľ
F�T2�f�����@�f�p����l�
���"�D,�G�8yn�o-n�֎��q�w�����wR�S-Ę�P)��q��E�"���D�6�	)�"䅴���x�$�v�ƼW6�p�H�d@H`H
dj��:��ÌT�1N�J�ⅱH�SD�B+���@������A$A%��(�[hA	�DhQJ2�.!IJ���	��a���,�r[����l��u���ng~h6t1�����ч��k{0${����\;�?��c$
L���Ig�k��iug�0�t�g�.�cxYŃ"w��EN:mv}����4����C,>�G��?���7a��鼪qX�-��YWv��n�Fc#��=Gǟ��
)x��c�f��?U�^ݯ�����ctP?�R��ۋF���Q��C�u���έo-n�֎��p�Ovoϧ�1;~�A$A%���p���6p�Kf.�x����J�.���:e:B[ox���"�4v�6Z��0~�H���컵�i�E�Apz�T�s��ͣ��T�ۨ컄��F���K�K�kD<w��g�W���*2�Q��-��E��}7�??��`����f'd�epyl���
�$@�i[L��@O/4Y��,4�-ӓ�p��C��R�ш���jA�f\�C�V͙E���g���1UT�_Yܟ��ï)��e�_�����Z�E�ttа��$�2f;U�N��	 ��xۣ��&3i���t���{�#���s֏#K�����Æ/F�5ȸ0�[\(m����U>{(��谘`"��	�QBér9����C��lh�P�^|�Ǡ��v����tqXգ�M����'�MϾVh�֎��9�����iX�<�ƙөh[m��ݗ�=��#:e�2�.2�N��խ�Z�מS�q\d���rwZ���p{�)4i �����Kmp��0|�cf㈝唬i��Z�Uw��so��$���"h�s��T��W��
5ώ"�cP�o(���L�C2;UY��2Ea�Е�rZ	 �w�PB�[)u��ӣ���|ɱ��|a=�wG_��d�������b�����%Q�ފ^��7�U(���G���g�>g�϶�ˋ�o�CƕY�������PF?�p�3�G
%���E��yE����p�jul�/4���ukyk:l����EI�?'א��rJ��#I,��}D$�Xx�0�H�ZH�xvI�B@��<uC�J�`�)�X �B<FPbeD
�.!#I�Xm27M�_0F�EC�q�R���.$I��ց��b�Je3�v���	 �	.
5
�L���mI-���'n�K����n����e1�s���S���]ٳ��Z�2�A�m�,��c|?���Qf�gɕc��a���n�_�Z=��(�w�ha�o��0vW'�>Y�֫rFY4a����a��wF쒨��CXۛ9c��t�f�6-0 �:���U�,`nD��R���jV����KG�,�"(��U1����M4Z��}��a�)}�гq���y�^G�o-h�֎����.�e�ؙX�g� �	 �����������ut�(�䯳x�K����nb����vqs�p$��P�0A���:5�q8߃�3��$�{TT�<��h�Cm1��N63�6��4iZ6��t:���8zX2��R�X1������{���y̦�	1L�M�	�Øh��7�m�6蠽A<=��ͮ����s��}��Sm�h�����_�Osx��a�M�0���T����0�8�]��?,۪y��e�^Z�E��Z�מS�8�7�s���7��٬���fw�	!$$��-`���_�)R����߸a���͛�Uo	%�������9r��}gWWD����k�����\
[>��8P��Q���e�B�Pdn��_׶�g��o2��i}9�?%v���81��Z,(8�59�<�m��8�b����P�a�f!:=�P�5f��3��2�-��ѽp��Z>:��w�/s��}x0ږ��2�-o�"��֎-h��)�W�_Wڬ7��푶�l�Q��N�]Fӹ)�V�Z�]�!$$��<iEh�ke�B�G]�}���6�ꪘ���R����H~�}�?���5a��������>��ny��߾��o�w��	��ީ�;F�b)scTa��Ǧ7@ͫ8�(�X�~��އ��r�t�È�f��M]>L;���ci�ŜXa�ݝck�\��X����CwApo\4�\��Dm���u�4�L���V�#n6��y��qH���"<�0�E"#H���Ȉ�6��l���ChB�ae�eF�GQםG��Qu�#��"#Σ����"4����:��"2����G�DG�iF��XC��e�F�ya�DF��F�G��mƑ�XDaL#�!B!�e�m�Qi�u��u�[����k[KZ#��"#��h�,-e�me�Y��լ9z��~�*�ﳮ{�����2Q!�_��a&��8mLΌ$8���2>:{jS%���z�t(7�<�UW���8N��'u�Wsx�&oY'���eS�� �[e��A���Ѩ4���}V��L1 �d��2˄Q*f4��q���3)��"d���)#���ͭ��H̄��PM�E��b�"HD${��ġ��ʓ Zo����@E2i�����\S��C�����Z�w ؛V{�{���uML�-��P4J6�axR��!W�(�t(�X*&4'M����NH�r�V�H6��������I����b��2��)�OWKGF�����`���Ў�b�y�I�d��yi����y6��hk(����q�	,'ې%�3��#26�չ]��i���TX/��	w�����-d�.N/_�D��edR����L��X.%��6@l�q�~��D
X�$��%,C�fpy�
��y#�����M4�~2�(�r���s9.:LHa�k�x�QS��$�@��ع������ؚ8�i�Љ"�4cݫ�~78��KXއ�|5d�_Z
�:��s���GH��� ��!�{Q	�������wkː��a YP8��3��Y���+��u�(i$��Q����g#!l����{��G��e��bx\hd���e�I�У7��[nH�0�ll"p�0�4xEsg#�y:}P2`%��h�*�&Xp��a�A�ByPy傒��Oi��y<����%5R(B%�8ن@�D'p>D���@�~�2{���wwl�$�L� #@���T�I&b��]��*I$�1@�.��*���+�:�-��N�n"��֋uh�à��F�𿈈4HfBԅ�0UN�%*JIB	�EN6T$��0�a)�5?;�9�W���Z�f�%CHȧ���I��9��h4�mH���J���I�IpQ�f0���M�1#-6�h�9��>z����L}!����J&�������������b�E�WR�Q���m^#��!����H�j7�b��"���Μ;l�w_��/�f���/.������t�ߕ.(/4tF�?��J�h|�}k��8
�ӹUUU�2���a>4xt��E�9�q��<u���Kyn"��֋uh��)�Yr�b�Z�֞���Ȝs=�5.�u�U*�uaڈ�)����#���C����]\�	+�y�&��(5����I��.aF��m��,�;�5̿Cg��R�wdq�T����	���P�h�H�5ϲȴ�-2�xĵ�����e;��%0J�JP��	�ƚO�����KX�O���|Q�h�5a�xh�����F����	�C��<7�#�LrW�.F�*M�2�x���4�#�Z�Z�n-y�<�c�e����S�=�	�x
�"!�����N�EY�I�WEG�΄�쵳�Ӥ�f��6	��^뒎���`�ŵ�@�K|��el��m
<��o�؈�F>!+�v3�&^<����0? ��\�WUִiaE�q�3��llѲ�bg����>z.���Su��8�i��C�*oE/6C�uٚR���r�i��VDf�n������9��<-h೓�:<�"6L��6�ѕ��O�~qk[�Z,����e�SM�5�N�ci��291ݚ��Ȇ��?2<�/��|�F>���n�p5Q�,d:X����e6�,/Y���`�5GO���e��R��,�TEj&�uN�^8�mʖDU�Ͷ�Z��I��3����n�}�No�����@��5�dd�����&�^�4u;�h�R8����|sн}qɫ����~vM�͟��o�������ﬦ;�CM|oh�z�xR�7�?hk�K!�D[۹�������.��O<��ַ��[�G^yC�C�x"���HX�"p��1�A`�<ÙR/k�[4���]Ł	����ʪ�#���M6
D8ʄ� ��v�.��ȩ"#m?@��H^�Ա�tT��G�%ȩ�����]�c�*��q�V�lllm)1�i�d$l@E��(�#$j�n=88�D������C3�~.D�g�m��<ӣ���j��회<@�Wv�T�6��d>N�3c��w
e�uX���|���ܰ0g4$<�F�bPIp��=F��@������î/}��&Ჺm��Rlc���t���n���f����\��; �=�ߴd�����<�4�:U��� �]h�h����`�1�kTx�^P5y�۫��	��?��)�Yu��G�����thc'�yn��$^f�t�;��M��Ql��͘�hf���2R��E6�3˛�{

�:�o;�Cd���0v�3o�׎�E�2~�f����Y��އ��߆�Y�4x�u7�)�b��oj�����&5�avl�a����βZӳ*�7D �B$���绿1.��@��.��t�5����3HáF���v�l9����zv���Q�FD?�<)�]kW�)�4��˭#�����֋qh��)�Y{��n���Ƶ����666_x���
�]�>gK.�c�[,�gP�oܢaG#���ͅ�_%QuR��m�0��j�A�Z�k��Yq{f����wx��£���1���Ɓ�C�|�J��!�gvU+�~~39��F�h�ӊ���`�C�i��Hyݺw.�;Q�uN1��vEЊ�A�n�g���&��F��d��	j�
��$��,6p5gZ;�2�.%:DPt��h��,��n?-o-h����u�uJ)J�	)��Q ׈*�i=�A �>"�����*Ua5G�Ed:��*�FXh��vY��M=�U��;k1Ӛe��rFWO�|R����ކ#�kƛ	M�q�6
P���}̯���=�.�s�=/G����H�3��Q�
͐�2W���(FL딭a�?Z}:�-��G�}��xn9��q�l����o�o���L���k���ʬ�je��F�~[��[�Z>>::���%<2��#]xl3~�Aź�́�'�f�frR�Q(�U4E�UR�]O��!$��I�����uc���`�UT�<�*]�}fe�F�GVih�O�ʯSj�	�,�^4o���@�b��YrHA��Edq�C!�$	�w��d��,���j��\.����ږ��m��l�����ߍtl�n9;!��?0ڰ��<o�<�$q�8�tet9>�jK���Q84`��;�C�4M���䗝���z8�m���U�663آ9�����Z4{��X�F��+���ܦCy!���*�N,�*�*4�i@S�]��Y�ۋcǠ�G����:i(���7����Y�"p�QC8h��F�y���[�Z-���<��0}�5{�+=Nbv�+ä	��ޗ��X��h/9��Ȣ+ᨙ���Ε���gשUXb�:��+����\�����:�$�2Lv�/i$�]�j���y`l������:�޾-�Ӧ~�z~6�����/��Qr}��y��5��{a��KA�gC�nI�Θ�����T�G8Q�A����rK(_��>�'X�UF3e{�;�^�7���C��F⢍ͻ8�����i�j�1��\/fQ�+��p�k�R�0�a�Q����q�����DDya��"6��#ȏ#��h�,#�B�:���eF��F�DuG�uG��y#��<����l"#�""2��uHG��"6��<��6�#h�4�L��E#(������DR"4��"<�<���4�2��*��0�)R�!�Dh�G�ea�u�]Dyak-kak[k[�G�G[FѶXBj0�x<���X��NH�����eq����N�H%�:�֌z9޴hU��Ngs�L�����,%o��:��}��R�#
z�>AiDL�tV-�{�@KR0͏�؋ l�3�jZQ��?-�=T_5����/��}��<Z��L1HX73�:K����}v��0�q���%���w�|=��ݲjI$��@�wwy���I&fP �]��&��I�� (ww����^W���]iխţ�Z�m-y�<�,����'}r��f;�	����E��9�r8p4Y�(�ia�y>&p8@�����n6F�,��mC(�����l:e�8W������4@�C*,�<PT�G�F�R�&�?�C=����^��~}��l�ܺ[�>Xg=`���֋+ǐC���_XY��6)�|=Z��O]es�I;��~
�t�Zx}��C~�߾�R<�2�N�~GQkC�:l���6QU�{g]In�wM��m���u�we9o�KJt���|���Gìy��{�m8�-���v�ʊ�@�EH�~���5��:k�V3�iP������`q�GWp����ca�d\;�G0��d8"�=6�r{g���&�] �ˣ��G��j����4T	�������>L�'�ݾ�˅�lzOZUWQ�����)�Y[/4��-E���מSβϪ�_c<��<N�>4e��<P����_��F�����r�4��b�R�bp8�*�ld�E�絕�95ni��h����irp�dLbLҒ&����ӌ;dD�j��l���n��	� DP��GVP8�J��B��q���4��g��$"%�m%�Z����I$���q@�v8\�"Q������٢�=G�-�}���!��NINS0����eC� ��KF�c�E�C��9dV����Q�q�a�h��a�����cu
4_9O����d'�+h�F7c!�n�|���R �I�8�2�K������7�7�\�t����]�ܫ�����M�8��[/2�O-n-E���מѡ���))R"�pٺI$�(�`�����⯶}��Qa���ۧ)C��s�p��d�(���t�/�O&����s��3�g�\W���I\����DX٪(� ��NP��i��gj9U�le�mIg�>f�p��1�{Ep�7Qp).��~8Z�|m�?pP@Ν�]"E\�fTj
�NEJ�m��p�h����Tx.�\4N����FD�ΰK�z�ܐ<�)��b������|�0���6I���iP�Y�Tˌ���G���u�Z�h��#�C'_�%���r�{	$�,�W�Ec�G���G�1����\9�ǲl��2�ޏ�̪tI⇍�a�����=gd��j�����p�쐓� ��H��n�p��c����R%y3����� ۞6�ԮJ�>>4V��X�l�p-��3�3Gz�!<fn6�`̐;|+����3F�P����U+Z4��9eV>˟B���N6��u��G��Z�kF�y�<�-LT���o]��쓎UW{��^�m�������; �GCn.�_�
������P�H�>$����բ���p�����1��2����d5Rc���JW<i|��h�o�(<p4�#Gy���{�f�ѣ�鍖lޕ�7ӄ\�����5�Q_�e���(��/��b��<�`$�����r{>TӃ����а�^���M8��{�ݹ�\sG:���D�:Z�!��l�a����6Q��Z�Z:��[�i�T댽�+�ZЭ����U�����['$�"�v�eB�T�`�-|���!IrQ#%A QQD��d��L��q2Nh��Ő��#](d2��p�X,pAA&c���XA��Xr�(G07ʬɗl$��%r8�,BH3�D�n2�L��<`�#1}�I$��W��FHbq	ȉ"Xq�1ȋmI�ｽxP4x�&��Q�ym��G*��ϋ7������y-�L��f�zk�.K����sH=�Ə+M����i��8t�-�QC:gG�[:Q��lp��6�;���uy-̫w2�:����|Q�7��~�U(�p��Sl�#مp�h������U�rݭ�ؕX��,ÊG�~e��Z�~GQ�ym<�q������>�{͹Wm��;l�hs�"��?v����m����Gu��-�S$�D���b��|��=N�QV����c��\��HN�ն�S�=F3�;$�i�Z,�i���Ş,�����]�a��xE�c�AJ>��H�K��r��J�ꪜ�7 �]�5�\>->�9V8p���f�d��ei�%#���..CC�_���ݫ3?u���G4�#�
1q����6Q���p��Z:�����y�:�,;�lq���Z�eoo�I$_xǠ��3��$�[�����������v��un˦O,��t�C�t�ƻ���-=v~d�~�)#^f�Će��c.��]GU)Զƶ��*-��K�FlÃ����ra�f�Eє�Y�5��[��|���v(���ѐ�g,^�|O�o���d5P�b��tʶ���=����.eC�n���e֞Dq��ykyl��q����f��E11n�I$�>�'�|B�#�{�2���P�(���*GH]���K�l��|�$���Ylt�q�UBx�D����M�x�$��xGxم7��*�����
�ţ��)aJ��Fz.�p�]�r�^�o�jJ�v��I��7�k��'���~8ys��l�r���ۓKh;I���-��-(�d�d��iayD!��D�"Y_�VR��cl8�{s�w����S��2�C��%
`�@ ��BI@0O�H曷�[��m�1!�3i0x����ݲk&�b�Zn��d��M1hZkLZkB���ZkLZZ-LRMh��KMi�1i��-�X��5��Mi�M%��E�KMi$�ZkM4֌�RMi�D�Z-1B��%1i�5���Zjb�ZkJIu��7YZLSZ-5�-5����ZkIAi��-1i�5�-MLZZ-��ZkE��Ŧ�ֶr�kJI%��Mi"�,�,�-$��	���"�AdIh�ȴ�JI%�Ii"�K&)%�%�K"M�%��I,���,�-$�Ihrf�I-ZId�"�"�%��IMLZjkMFZkE�I-$��$��D���I,�I���Id�Y"Id��%��d��	,�,�Id�KC���GI$�I%�%��I	$�H�I$��Ki$��Iii-$��$��I�$�Y$���&��I-$���&�Y$��Id���m%�KH�,�,�m%�I,�[I$��Id�id�d���M�K$�,�Y$��m%�$��K$��M��I%�Ki$��D�I%�%�I,�D�I%�%�Ki&�Y"Y$��Id���$$��-$��%��$�I�K$K$��,��-)d9��Ѵk25�̍fѠF��[di���f�m�Y���4��4��dk245�[h��7��p�#Dkdh�ё�#XC�8�����,�D��Q��c��F����F�#XF�F��bͬF��b4�ѬѬ�����3�F�F�F�F��1��hѐ�g�f�k4i����m���Fp����ۆ��fF��i��F��1���F�k4m4dhhѴhhr3�F�Ѧ�Ѵkf�m�XF��[��8���5�F�h�4i��c�g`�5���Ͷ�fж�,�d!�m���B̆��[��Xж!M��!Bl����h�CY��B2d-�d&�XЙ�6F�[4�4�[d�dѦ�MfM6M��6�M�LMcM4d��4�5�km6Bki��i��bk6��	���m6Y��	�[bh��	��4ؚ�M`�-�5��lM`�f��4��[m4	�ؚ̚6��M���X�ؚ	�i�a5�44��Ѵ��X�M�FM4�l�&�Mm����hɦ&�Mm�ɉ�&�MfMf��4[i�4��s�(wM��k4�X��4M��5�h�e�5���4�k4�M6Mf��M6�-��i����i���k4�Y���-�[i���i��ѓ[i��Y���*N72h�ɤ��h�5�d�Md�i5�I�֚&�&�I��M&�h��I�ɬ�M&�i4�ɢkM��&�i5��I��&�m&�Y4�Mi��Me�[96I��M&��MZi4�-��Zh�ɤ�5��k&�4�ɢki�DY-�,�D�"D�""�h�"E�4H�",��"Ȉ�$YE��h�dDY-�FH�$[D��"ȑ�,��"Ȉ����"E�"�$H�"��Y$[D�""�$H�""ȑdDH�$5�DD�"Bȑh�BE�"�"��"D�D��F֍h����HZ",��D��",��"E�$e�E�"h��H�BE�B�!e�N@�dH�-��h��"(�-��i�,����$ZD��ij�@�B�"Б��D���FH�$ZDCYE�d",���$,�dH�u����9�E�!h��5��H�"F�DB�!hh�!"�D-2DD��B�!�	�B�!�	�-hPH�v�p-���;NEn̍dk#k#Y��CYE�B	#Y��"E�Y1d,��E���bɬ�ɋ"E�Yd�DK%�o;4��y��2S_&��F�T �zg������c2ѳl��(�	d#P�H��}����׏w�ܚ����/�~���1��l�7����H ��}FE�_7P��U� �X@k0�b�D�p�ʘ�j��u�H3NAW}�I���X���ڈ�#�xT5������PT ���z�'����_���;�@Q�z�����&��W��f����ߺ?��|����g�[~)���>���:Oa� �7�@T �|s����C�SI����M��p7-���c�t�j0��ay�}ޘIIO:\x�BY Jp����/�<�;_f��ԼO��;����;��RC�~_]���?]��8����WF�sRQV�@PUVe	UPKF�u0c�F۩�e��EI`� ,�����b��e��@Z�_�Zx�J�j�X���Cvos|������`ƠǢrͶ��-a� nC�p٘�!�������q��ofwx�幃���@C��poZ��apF�P,$�`Zv�j�_��q+>-�
����b�lz��-> �z,��: �����6�Be�p,;Bq9H~�ό�a�h5"B�36;A�A:!���;��q��Π* kC�,/���@xD�w����1 �:C}�o���كOC��m���x�U!]�����J)�P�򌆡��^�`Ш'�BPPQ���@D$8	F
:�, ��!D ��uZ��-��Z�� �d"RF������[T0�.���AH���[(@��]�?#z�6��ކ�}o��a|��_{a����w����s���4i #�xz�G�8]k�UX�!ԛ
HF\�8��.#���Y�J'4��h�Ԏ+QAPT�`��:�=��zT@���/=��C��xp8���4���3�����^8�<D��?����ۿ��ukA*1v��jq 
b�R�����1� �`TxX%��r]��A����6�
�q��@ցu�b%!�M˰�C�C"T�x7���	b����@Iu�D�A�����p����!�0���� ��� ���S��^���ԥVC �ss������p]�[�t��$CZHH��\L�/�����w$S�	ɇ��