BZh91AY&SY�u��5߀@q���b� ����bB��     }$G��k*�JQ
V�	��5��R�lhM�֩%�&�T�,���j�Md[Vٕ)�S,�(�T�ٔV�Po-���o��%AX�%5E�Mf�i��V�Zm��[md�[mKj�bI�m��բmZ��`4�k�֖���j)�4�(��M�U�
�d����%JJ�D�ʦ�me��յ��C TV��kl��fիZ�����VU$��`��44���I��V���ڴ�V�eZe���jW��޹�mS,m �  ���k��S��[[Q�q��CWn�Z��(WN����۳
U���F�m��Uݙ�ª�n��;���dmsm�$������m�   �P�r�҂�s����u��V����@((��:��ڦh L�p 
;�ۀt�
����{����
kl�m�UTj�7�  �\y` ��6� .�m�;�PYJ R�h X�(4jaХ*��s�@��<� ;�Wm�l���clm�Bֶ��x  O���W�=��T�m�����g��)E�=� A��p:� J�( {���@=���z@
6{O{� �m�kMmZ�U5m��T<   ;��: i�� �Ҵt:� �R����@v�.��:pp(R�wc�v Sg56 p�8@:ne�IlͬX�5��@H  �枀��[��� t1� �0�ئ����M�F����k�(tܦ�  8n�]�C�	Ѵ� ��-���XҖ�ERO  ;���P �����p�d�n�$.F� .�  
̬ ��p���8 :0 ܅�����@V�)��  ]� C :4\�4 �. 
�.:�W�  ;�� r8 P� (�N�CAA��#j�Vh��Z� d� )K�\ []�  �0 n���e��(`m 9�8 �:pTn��sR*m��ř���L�R�  {� {�� �k�A�4 �� jqc�h��� ���� ���7` �L���      L�)R�M 1 hE=�LR�U� 4 ����O&!ITP 4   h T� JT�L 	�   L�I���@��P��   Ѡ ��M�A�f���F��F�4�OI�����<)���~+f����s�U��,��/?>#�����x��� *��AVTS� *���@���~'�H�8O�����?�uS�`����Uz�����	�L	?���H_� _G���_��C�0���ȟ��?{
~��(|�'�2'���,	�A�
zeN��X3 u�:�e�'XC�)��"{aN�L��
u�:�dN�'YC����#��)��
u�:��`N��XOL'Y���D���dN��XC�!�P����u�:�Y���� u�:�c�:�a��Y�u�:�`N��Y<�XC���@�(u�>�!�P�(u�2�XC�!�@� u�:����� �)�^�Y��YC���P�|2�u�:�a�>:�a�YC�!� ��e�'X^0��:�`N�'YG�)��eN�̡�� ��:�=eC����ȝeN��Y� u�:�eS�
'UN0�eU:£�	��"��TS� �YN��=` z���#�� �P�
�`E:��u�� �� S�
'YT>Y:¢u�� ��DS�*'YN���dQ:��u�@���XN���`>O�D�)�T���|0"�a�U:�
u����@S��Y�*�ez� ��C��3� �"�YN��=ez�*u����Y���@� u�:�`N��YC�zez�a�'��(u�:��e�'_�u�:�d��@�u�:�d�XN�YC�!�@�|0�XC�	�@� u��)�@�(u�:�������zw���,h�ˍ�T��8l���9nhr�l`�TBYz����)���NEPU�,�YYT]�X��m�q��^Yge��#[.�#�cNťX���=Y6n=Y��F����+4]l���!T6�hj�x����ͱI�gT������!�);�'����e���j�ӧJ�kM��KD��ݩd�/0`R?��|������#�I*����;5���e$�#l%���q�J�<ڱ7&���F�܉���06*k���e�h	��hm˧#]���]t�i�ê��6�d�X:�h����u�MU�"��� ���KXؼ���Z&e�Ȯ3��:�@@�zTݳw��5�l�o,6*`wl9�kӬ�%"�!�Ԥ��5��Bn�פCH�L�N������ݖ����x�;�h��5�x_�0bV���u��#XU�r��Y@Ӣ[YR-�X�ч,���%�#b�BD�B��)�� H�H�`����q0����*�9z;4'��grǮ��AM�b.��Pv7[P�$�-��)�A�zd�s7q�Nέ��)P4�(ѷ50G/ˬCW�-��[yR�%):�Yt�5M�-L�Q�4�$µu��U{�ݰd9�I+]�x���)Гn�cvr鬴Y!�E��5M#�{G6�߱bՑZH+:�4c�5±�V��YV�PO3��*��OZ7vڙQʴ�-�80�����L��be�f����G(;ʵ�H�Q�Sj���ĪH ���WL���qݑ��=��Tm�͒@�#��E�$6�wh;[�a��Z��x����An��1�3mSp�g.�n�w
.u,�yyw�����\�76��m\{5�E-Z��4�j��xh,5ڳR�(��3ǒ��,�Gm�#\�{g|����Ӽu�sq`������1�0����6�iU���ϲ5Z7X�1��2�D�e�OU��4��(�H,����=ui�n�e���ʈ���[h�v)e�Z5!#y@��wn�ț�Z��4���Ҩɵ��;Cv֭Ȣkd�낆]��z�d�l�nS��ʔq5�j�0�H�hv��x�V�̹q����4��n%Z7^n��T��J@�
�}bU��w 4�;kA��3m%N�⫓6��-��f���9�6����cB�b�Ví�w��]I&h���;y���ʸH��O�`r!5Ww,t�nQ⩱c.��`v�Z�c0�*�����',nf�D���"N�GU��I8�F�&KA0^3�� ����zwm�� ò��Jt�F�����
B�`X� se�QuWu�ɣwv�Ua��C�U�&���ųq퍨��+�P��!̗����,JJ�s�
�f��jxC�u��B�ǦS�Ѧ[ز��cٚ��Vk%���ӛPJ��H@�v#9��t�3 bxF"����m���f��:p�+p�g|'a�Wwe[A���i�!z��vQ�ѳd�/"��W��L^�L���!f���8�B0ӽ��#w$�c��%k���e��u�ɠ5)j6��,��nʸ�oUvR �	e.tP
��������\J"��-��E�r�ZŬx�SǙ
�&(��Gd+n憩�ܭ�{j��#s5��C=��B��CC���-]�HїZ�M�yKr�2m�X�`�������Pz����h��+�^���ֳ����-k�%iY<�\��Y�g$Zش�W���ݛ���]�f�J�.���H��ź7Z��D0�:F=�7.p�͚*7���Ց�X��r�1�:�	ӷ�-��/V���`��J�P��sNʗY$b<w��[5=K����:���i��`����x�_m�k)b���nh�f�PSe�z�::�ڧ�к�N��Z����f�	�*b��r��ܴ�׬m:��v�ZZ�؝.�f��bI�l�.��n]7ͤ����Y���[ڟ�ѾV�Zd��VM��٨0"r��;�VX��u9�m j=�̷��rAi�����;�N,�y�m�v/b�l�I�S2v��u��6���d]�i�Sh�Sm5r�@f��
^֗x�)$uJ���vl�Ė9�vc�b����ɹ�"̬���kf���E �3"[U�e�av^Zږ��s
b]� $aDn*���z(%�DM��܀��u:�5G5fp�3]�rU���ӑ�a!f��k/0̢Ҕ�$��&4۩E��z�n
�	�*�y����h���&]�ۍ�	"[:v�l��t�Zdi�ˬ�ȳK���[�i�*�;�+bA�#;t�[�6eRƯ����VZ��-
���ݎ˓sp�b�yO�V��F§�Z�Orܠ�@v-�N]���ixQy��eGaK��^\�q=�sZ�n�Q-Z�v�(]���r�`մ%�����;G-�Ŭ]fN0�l�o��(�[4V�����ڐn�W��0�ɦXÛ�C�m�cR�K;1V�k[�7w; �
���O�����CJ��q�f�8p-�C"*Cn�4fɛY����(�r��C��,r' �[�jס^�r�r椨*�9t�E�uzPs�tƉIG��9Ji�V���r6G=emcj��cnø̓��:̌1f���9�����0�ls�q�����e&��9��in�l!eE��n�=��V�YIag@��nx��o@��Mhݺj�#1Ғ�]8EK��[�W���ㆳ+Tt���m�����VoL�V7b�d�)Re���̻�Ś�J1U����0�={�R˛�6��2��W`h'H�Q'^�2�xi(����%�k��[��-I<ߴ\˫�C�Z7�rA���EK8��i�d�f�͘�m��V��Ui��,��|^�-a{�v�]4㻀����*4��Nރ�������9J}z/u��M=U{y���cz�-�Z�V��xF�
�؀�[1R�vޱ슭R�oF��d�`�kQ��������6���OS'��� 'r��1C��e9sv1+w�RQ^I��V��-���0hx	X�ۘܙ��͡u��𭺙j���ߚ�")TY�v��X�z�dSP�@f���K�ʰ�&�j� ��=j�)����.9Ze�R]�EYx��� ���#wm���f�sS˛�q��	l�r�n��T�e�Sf\�6o�W�����۩��i�1�kDAHw�魕�|K[s]�kB>���D��;ˤK����s],ٵo�=��4�ky@.Z�&+-V���X��_Z��c�*�$��N�tC�z�.���ol��m�`j�x�R�^p���mj��bf0A�C��>@�m4$y��<�.�e+[&H��Row/J!Zr�ת�:�S��[n���.�2,�t|~�h^�m:j�{n�6�/�eZؙ7o�Q'3Vh�o�°�zV�]�K1i�yA IU��Xw�#-# ��kGIJ�'1��Y�f��N�l<��T�g4:��8�7d�m�%dh^L�6S�f���/N�Fd	��m�h5۬w>����J��y�f�x�P���v�j�V��5�[nbѰ�Z��f�#�f5����@�:�ЋBZr�{� �z�C�0�зVXl��&�34!���w�,��6�-����v%tn��,1;Z�͏�4�UE9�V���n�GBS`��N��`�1)d6&<)sv�l���v�h0e�U-і��nxE�$�,M��5�m� ��'I2�`��U� ��7W1��7N�Z30V�"�X��É��tZ9$�n�ٱ$����P���6��{Wc"3�į)������[��0n�[R�Kn��9�uЃ�S�D�B%ǖ7d��ځ�6I׊��m ��XF�1�w[=�9�]k�
W�:�ư�ȍ˲�#�v�V�SУW-/X�O)A���hf��Z��
��������4-��c��`��ˢR�{nm4�,OA���<�Q�u�L9a$A�"�]�ƗS�I�3	��[���[����ޖ;Q8�9Rr���31]$�ۆ�ȴP-��Fe���0�{���|�̧�ᛒ�͋4I�+�Pn��H�R�����ʌ�d�@@�7�[�Y7m�f�Nꠥ$�V�fT�VL���`%��oQ2-�}��.k�i�֊m���;�N�e�C-�T��7NnŵB"W�z/a�ޤ�thf�)���+����f+D�l�������Xk%���&�h��%^l�`׹d��TƠa!���;�^JI檐сj��*Cd]r<5��Y�^S����Ԃެ�MF!�������`��e�E�j��Jy�lhH������уt�)�k�kQ����
ͬm�kB;��7a���$�"��t���T��(�.���V�^^���7z3-ػ ����K�=�m�g&`^�9i��7v�T�[��tE�M�fatƺ�U�A�̈����׶/g���xk,U�H0Q������<

����x^3�2�\h2^�t\̙X�m��X�X�컌<�Y���V��^���L��Ȭ6a3F��܊��� ��unD-e-
#���V�"�e�)�v�j�7s,�lj*�n3n\ҙI0ѥgn�m�$u�Iw�wrmɲ�V<U�4�����ЅV�ߎ�ڸc�<Rҗ^ko�XO�Ŗ^��OW�ڢ�b�xԘF�� SD�=�)ws��1��j����3.�j��8�[��T��+�d�[��<�^klЦK��Hz7Bʫ�\v,�T���q�i�R:��Uj�_͜s,���]�JQ��l@�-]��.c��3ki�E����2U�6�T�+9����g%f-�(kv�2���z��-
�^�s&Z��<6��tK��vi���nجQ捼;�M�S&�2D��IK8.d��-�I�84R##5�0����j���%�6�M�Y1���y�2e3�gPE��TU�l�kͺf���^��=��3~��<7*c�u&�̳��Z�l���ɪ��v��!iYӮř�h�=H���]hm�K�:��g/j���M�vM�0�V���۬��͠%� �hfL�d��i���q�FM�0��3�c��ͨ5X�a��#����6�m�j�\O#;�!Ǳ���Jì�J%mn�/0)bT�R�"b�ۚ-���fm0]�����ڑ�C1�S�4��#Uଁ�*�X�$Cz�6R�9��S¬_WX�C�:����k�O�ku"p���Z+;ZX��&�[DR�zq#�F53�c�T"��h�E�+�V^ �1�n	����+ͤ^���Mu%�ӈ�(]d�4��[KUˈd�݆
r-v9@*��%�w6��(���Ċj
yf�:)V�]�-������ɓ6��Tja�[1�[��� T�	N�ЕۗL�(]�pM4йu�����a��kby��[OKu�6�䥉%d��x��k,e���5����Ҙ�V�����j�?L�źNZܪ6�3
���=Қz
�͂�ғ��4^j6��8Y3 Z!t,�GJܻ!�7e?a��M�RMP�N`�u�(Aci��Z�P�(�l�!p7�t�n·S�t��2D�I���2�N��۫V���؅n�D�FJ�ҺG	X31���h:���O~Yu)<!�lP�ǎl;�2<R�Ym��֌���L1�t-�E�̹1�i�PD�%�djY�c�#e�X�Z.lo3oF�+[�f�cc�c����{�wnl����.��e��2�kv�V���-jK(�*W١�2�I ��cL^�Vf:�W��i��O�I�f@��o�k���D#15��-�J�԰n],X�����y$'v8�6�c������oiK �U�;�cU*kՆ7+�T�E��z"��N\�M4�ٚ�[�D;F�M���n(�M
�YB���8��'1�j��$°́���iۂ&x�P�}�;AZ�Y�Ǌ˻HjX�SU��N�ҫ�wV������MK`Б�T��{W����A���N�yqmj3J�E� ���{�<�fX��P��ԕtJ9N�U�2��;!��G++up��#�1�(����ad�Ml��.ܼ�̢u1˽�f����G��EYPn,[�RB��������8�VR�����oj5̛r�L�1M:By5�vA�z,���e�m8 aRV*���G6,3X
�c�<��x�N���d��m�:N1�����lNb{�J�V�|�e�j:�Y��K��l�N��{a;�"F#pR��P�Ę��yeP����"�g��N�L�RX����{��ۍ-6�BC�e�I���u/.��U@�YS
)�*A=9�S���jue���̦�ʔ��g% "#2�:&c6}`�ld��M�5��b��B1�ͳ��h^�ylR��$��P�4Ry��Fݹ�+mf�c%�ʖi-�1��U�
8���졅M1��-ڱ	R��vvnDtmn`��C$�i���Tlf6iV4��4�(R��܇qQzb� �MGn*t!��w��ڑn��+,� ���Y@����qD�J�(�l�]RZ���%�U��*�m����Y(��M�yC2�M�Hg��9�lv��}���OMY�XZ;��`81��I`��V�1(���p���0B��Ą��2�2<��`��8�4.��(#�ی���,Y`ղM��L�ͳ��hC!�zc;�w#&.�"�����i!�9W-r�z8տs��m�d�y��R�p�@2����-��W�Է�`ƣ�f��qIFi��h�d�jv�c!gb-<N�bQ z-h�X�XET�%I��"��J��a�2��l��^]٘�K)0k�q�M*���l	%���"$�!Ȣ�=ɐ�Y8u�gt�!��jR0�j�:�	�t�pr9������ւqf����&�܊# ?����3�b��ܗ�kF���J`��~���Fn�x�����뽖�P����*�����%����f�nQt֞t����|� *d�f� �YvԦ{�V9����\E�"��)2�B��׺s���C�*!P$�pݵw��f�+�ð��y���J���7CW�Dr�,:�p��}�!|Q�t��u69�KS��6��]�C%Lt��䧦]X�9�y�\y�s-p�D�jci.���{1��4�&��C�{ff�r]ݢ7�N*��Z׸�+�S�qޮ�':S��JC��i��!z��:�ub�\�[ַ�2X]]V`K��K;S�l��*	�orG�l�m�ݥ�ũw2� �!�����6 WBK6� n<�kd�3E^Y�૔:N|�Aj�-=��=�EP�������bw�Y����wN�V�#5a9`:���"1i���"\Ln��¾��
rjãam��f*E��R�*.s��{RHcSb�y�r6�rq�z�B7X��a���60l��@C�7f�-�9���B�����̚v�'�R}���X2M'���z��ܰ���r|#9�Z k�M��a�0��hi��}�r�Vy��'V�6N���W�rp-ɢ`�I���j�n�JL��h��A�o��sQܤdCZ�NfR���V"n�&f8n;��2"�ָ���[x#��o`O��Z������L�t��Xi>�R{n���Z��v5��t��+�K��ƀ��e;�� �cˮ�yp�V�.���(��V��e�|����'�5�( �}��W���E$㢮��7Sn8 ��F�C��7�m��je�R�ܷWi�i��X*�on�uZX�ou���4s���3`����b�fd�袉���~(̇��6c�r k7�oNt7R��H�"c���Jd��˳�Nt�9���9�!߮��YB<�`������˷�Y�=J-�[���H���>�rr�s��H��YSG����e
{e�ڼN���֩|�MʷBV.��;��]�{N�0sV�\O����3f�������q�w�˦�����zl3���4�������O�9پ����wxm�G�j� ��LD❗�ݑ�NIcm���^����w���K������ʸn�R���Ӫ����l银䩅���%<w�J������ΐ�=���s��]6���]f�Jn�k�؎J�|�87T�l��u�ultT�t84)�C��}b�/��ߵ��^�$þ��������¥eXC������1��{N�v�2�`b�����ΆgE6�YAӷ5��g�����3v���3��u��hC���!���;Wh<qwM��m�����"_����4�lVq��C����c渠�2h//^cm�$M+N,������N:動kٍԫ��C5 	9K��J�e�c�f��N���y���FfD����\LS��dMd޸���
Ȇ�w�̠u1�i_P=v���[�6��U��MN��G���E&8e���&'�#WA��ׅ i�N�v�]n�A��O:�~4��``�V����=�XM�k�u���2��3 �V[��@���ث� 73<�@�wz�h����L���7Z�e{ö>�x�MԨ��K	xk7�Y�p+Y���f�?c�#���5�9}yW`���bΰ"�ʂq�:�|�A)NC�j�Vs4K:�ٰ5��^�i�9���N����Q�p�C�SL�q�zb"�o�(ɳf�u��OҺ�h(�s
߻���v�\Q��_u�[vf�#���y�R�0t�7�8B{|Cd=��(Uw"�-�ld����OGx���� �8�ol�m1,V�l�{�н��8��b}G������r$��:_Γ�kT�%�1J<����hǤ�α-�:�6��v�;К�����o;R����JP���e��ZV@r�Ђ�;��l�xr�����Y�"�jF��T�}%"/D}]`�Z���\(l��ǡ��4k��E˴3U���G��Pre'|���)�6��j��0���,Й|��gL������u�$�N��m#�-�祠`��:�D���F;�L�\|+.�U��|��8�L0�>���Y��/�T�CB�좩�Y	����޻7.)��͎�{J�
MJN��h�!l��W��I�8�Be��h4���@��Աr�2��x�*�K=B���7,Ko�����.��N/;M&9�T��N��9�:�je漰mY�q�w�l�#�6�)F�{v;6x����Α��يmt�-��Bt����R���j� �E�ؾ})�%��P��3�%%e�t*dv�7�;R��{kMG��f*c:ís����AS\G��Uj]j�1l���}�r��on���ڬ�f\{zM�urt�P��gu)F�6fdG�����Ƿc��̎�$�z�n��9 E��<�c2[���R�Blvpצ��=����+.54j篲R�<&��+�[���7�']w�����j��]����A�Mv�w�3%��<]t�[���m���dǋi=V��d:J�Ӓ���,�N�������+ۇs�U�Q��t={���,��҇�1m2��9�DС�}Pfҗ�ȵ���E��eZj�Jg{`��Jh�]^h��.��\.Bq�m���;��@��$r���k�/3/�3Dڛ��S4�eB�g�M�����r�l�<��V�A��Q2f�[u��W�2�T7B)j��B೸�٥\y)Li�ɢ��^�AΏ{�X�ky�n��<J��+A`�!nm�^P�R����ګ�]�bT�S�GŞ��L�屡 )a���*�fery�,L�ڴh�sV���]G9�h)͈��Ѧ�u�P�Gi-�/q����-w���^vֱqnM��w&0,��7wBm�&�[����v7+.WC����X;괟"�o4�Ƿ�x�5q����e�pr^-c�D���|GMyǄ��V��0���ɵ���U/�me������I�k��i�p赆�^:��J����L�ăW�q,p*훬��e匌�.\ӳ����r�mޔ6D�x�
�4ڍ��2�J�M��g�JH<]uu�V�'nh�;��;oT���v��o��+i���r�eK��Ӵk�Y��+���#<���NgR�˜�����e�b���S�XФ����|��&c['f ھ�U�k3T�v��YES�����{Hh<<�LCc�@����y�w���dei8���t�oU�9�[N��N5�&��fdb��IW}mǅ�|I���r��K�W�&��DT�E�Y܃����{��L�@�����oA�*ؾU����uS3�ok#�[QY��0�Xe���i�Of�.vCI���NR�u��*�1Z�3��Ǵɣ�,]������@��}2��S�g.�X5�-ќH�b=r;���՘6#���Z�g}�[��չYϻR�`�(�T��KU�A"��2�˻�P��:��Jr\���|���!1L�g����i�'m�!65d��S�z�4�Բ�$�8M�⛥�Y�o1SuB�\J¤oH�r`졭_d�ݛ �y2�.��%{�BFܻH���<Bwk���3x�� �<��@j�sP3y|�Ѥ��;�q_e��'�.�U�pb���맂��2r���]n,��,�,��gK��%]n��b���s�rغ¹�8q�Fˉ����ú��ׅ��M���B�+x�Oo+���uR�f�D�Wl�n�xtޕ]j�[v��3yBs�1�3hF��n>���x�g�]�Xl�tʫ<f��e�I��<3���iT�C��]�3�k��]��*	ԁ�+��M깪�W��j����A|^�J����-�9}�dVy�haP+�N=�e��1晒"'���Λ�θ����L�&�u�}�R�CT��pY��oI�[�V�y��)F�7AkQ�V��KH�|ზ�PY�̑3%e�O/pGZ�EäfWr�l�r��0�K�"�l
�r�����zq����8w���L\��+9���0��t(}ײ�����$���9��pX	����=k��	�Z�T��Wf^��%�C�����w%�.�V��Y��<�r7�4�o%�fq͑���%[��*�z���o���r�rf���
���Z�-���SL}�{T߱���K�:v�ɨĖ뚷
Gf|�9u�L%^�,G$�y=����/�#�j8��uvN�i͚��q)��4�p�	pr*9'E���q'�8,�T����Lik��9/_j�G�2��o9�敍e���1L!��P�m��B���+s���������/1�����7|L���3�'�,֔u�4�u�6;�K1Z��KBVc�d1��3�U�n$�[,� 8"�����̣�M�M>�5-Gn��t!]�Tvw!�3r��l\b�6,\�������/�7��R��U����q��9��G\u���ퟨ�ڛ�Ycc����B���l���vT`��4:�G�0���7c�U�mƎR�X�l�]��>���v��Y��]c4U�{�ۋs�sĵ�K�����{OesX���h=����5b� ��6�Pcf����<���;�e���VO���tKi�ފ�oXٴ�B�T���F���v��&���s�/�X��^ޮ�)���S>1Z��%�\��u{��F�����Y��Ҙ]_&)�8)1]�b]c*v��M�\��-�a�u�&+���Ƥ����;6���6��(�.��b���6s��&��#����f͸��\��g8(���2la9�w���g"�h�#y��Af�2���#rAx8i�x!�Fsź4��U��
��8�ip+���&�=�u�)����)u���G��˹�͉�9���R����QE�pudƳmnC��T��I|����ͮ	�ܹ`@�%e�ܬ��w��@TR��I��Y��L���nK��N��g��yy��rL�X�x�=Ƞ��\�{��ZtA�1�0��qb^�\ћ-YM	�uz���o'SX+��ƒp��W|������	�YzWM��͵P�����=�FWc��r[w��uܺ��Εcv�K�+Ű�A�*ծj2�	w8V��Y��D�f�J<ؤ3��uu|�����^`Z]^E�ػ�z)�#����	sz����6�"�'ok,�Ia�RV0�qJEb\㷜'Q���f
T�$��:@΄0e�n�^�,�r�ͧf�u�g�LS\1�R�-^v�4�s���A�����rS:Ȩ:I��i��,���{d�۾	�N�p����﷈.}
��v!�b'��,D���W���d�"�g���L��G&���W'�$�q9R�&C.�[}ζ�ou=̓@��Jq�T�x�R�#v:�>�FPT©c����˞<j<=�aFd���[cފ�V�5�btœ��3z�%��ΞD��L��=\�w	��6�]AOj�k]^���Н۩&,D!�y^(�ؑ����3Uh�yt����(�j���;)�*
GQ:��͹�)g���� 9�
���a9�h���H�:�&-`Y��%�(��Mt73d;�E�ªF�'G�o��j��.K��tz��1�R�U��Wi"��V�����=$P)��u�ͫ�\4��z��U�,u܏\[v9��^m���ά��:X����r�9�B/��:�0�kX�^k�pi������gҴ��I�$A>=)���n�r��r.�dfܺ5 l��Pǃ(Wq&w@y+��x2�=])��F�N.l~�⣙L���l]�����Mt0��溑z0՝y���0n�d�x��gGk�q�}�����!�jt��s�	�i� ̭������&fK%{|����z�p���H�k��\�7ܠ�VA���Q�K�r��ֆ�W}[������
)�t���7wO�d��ݒ\��2�e�&�t5#���"�|�@��bF�B�3Y�Q�c0e4�|Y��7{U1uM��0+.�u{gu����YC�J��շ���V�����h���{��Vs�L�6븅�-]B��w� ZA��>[E�s&JT3�eZ��֕��0r�f��@��DI��\��X�)+���6f^���3�ɪ݂�.��ląr }c�e
��l�2�р��w��$k��4�6��c��>��FM�ۥŗ+�!ry���4�l��d���5�@�nr��Xښ��%il��*@
�
|�i(ؗ�3�u�2���l\;%��v8}�-ډ�﨔�S>+���9]ͣ}�818�����@3 X29t����q�94��M
�c׭ȡR3�a�
f̖c���kE4P�D�W���>9�վ��e���_��t���Cp����N똗gE.�/K-�p�ꎮ� P*;[U{[M�ٲ�p�+�T��qʳ��BF��\0V���:E�t�I��nf�DxqNmX$�x��Y���uu-�jv\$,s&��j��Ky^pqO�U�Sn
3�z����\頾�@¹]q<��4��)6�1�Yu-@�K��]���d.��r�r0��o�����Ob���I��L��0PuF��/x�̺�!��|��O'�iħ��H�4�O�9�z��)�7����?��<ޯry��>|z��G��x�A��A�O���/�����>%=@����O�Ϭ��s�����=K����%|Z(<��`��"�Ϲ�������}�����}�?���K��̓&dɛ���޶��v��A��}�{����b�����S�ۨq�b�3tf�J�LݍHXJc��/9c;F<���4�S��/)�����V������ú9��ɼ�Fz�We�;1���Ρ�YS�t���в��켑E��'Qm�N�wrgd��\�+�ȫ6�MZ�����R��r�N�n�P��$;����ц�e[��GI��&��� �Gš��UV��=�ь�<��ͅ)�I-Z�����,i���2�>��ij�	���Y[קc��t8�/��1m%n&Rzr��>i�b ��y�oFp�Zޕ4�C:�z�VP�P��r���23�#�g�[bƫ�u��E1U��+;�Y���\iU����7�Ed�ؚܸ/9=ˍ�-u�'9��(���T��^r��;�ܢ3�p[�ۦ��)���Y��p6���)�ݎ�h.�r��b�p�f�VS. ]bx&kg���XF��m\��%6��a�:Mnު��`�y��mI�MB�&���4+e�J��D�5��óY1}�т���Orm��P���-��r��r��ӑ�V�tH�h�&^�j*�d_k��|��k�	
r��ky�^J��h���z6��T��C�E��Zʙ,d�]ܥ��n�͗Fj�(:�(�9,���ě����cMa�w(;�ɾ������Z�̲� ��Gdoc�C�o+&G	�� �������\ů���l�i�[�:�E�ƬB���}��X�ș��O)o]�e�$���iN�z�æ/e���zO,c�!B���K����H��b.�49V<����d(S(b��ݫf�b���Up��"G�p8k�>��A*��
s1�%�e�Q���:��lKn̸�f����F���=s3uq�B�v[�Ķ�w0�� mf��#kX�w�\�2&[ڷ�w:N��n�I���G(mN�6"D��l�Է�r��[��e���b�ߏVn��bh�0���*��|YL�!�v�sձ�C���>�Y!�rĭU�x��-77��/��I�8\Aʋ9��[=�Lq����r��KR��v���B�yM�y]O����t���2���Lf����.Hjd��3Yj���B�*U11D�S�F���*,�_^e!/E��zə�I�v-͎�w Zx����#�l�m9i-����lLc�қ��%)Se���Aغ��sb�ρ��SLt��r��h��5Y#� �z�Kwc��^$C۵}:��N��s�����9Cw�K/^��6vl%�T���V�W���ȝ�%�tc�/�;/�ʂ�l�i^;A��a�Ԍ��a���n�M�,�E�*���x�̸�,�l�����iWγ��Y�V�;�@����k���ϮZub�ٛu�R��r-������M-SS�-O_U32�J���Q�n�t�o0�F.��Wl׽&�����u��ҹ'lA�D� *��m���G�*�ͭ�* �2ε�]9-K�L�MIN�5M�e*$&#�ҥ�m�&�3���|��n�X��<�r�\�#V����F��ۙ3��Z�"f�!Uu��eh��J8+G�1([a�}�[=�8cWYyt9��;�nsв�Q���~.�o9�9�uHh��7Lڛà�%G����خ»=��A��z)+��ń�r��ۼ��՚�B�Z��R�Ep������ZDj}35�&J�Ă�{��X5�O5��I��5���e�wd�ʖ6	�i�ˏo\��;̙ב_'`v�+�A�e��k2dm���J�3/B�6���}M\�o�4Ż�r�����H�%E�V���"/h��i��y�&�Ջ�c/IT3�P�S�dG���$\g]�7|SIX�ޘOb}n�=.�]��vB��M͹f�J�n�f9S��h��i܅�-eFoz�������2<�Մv(�{��Bvo>�����vp���W�S`�8��mL<&�4[d�loNSk���Lѧ1��ӷ�����4u�ui�yQ`���
�Ku3K� �}K
X(20���.�vpS��;�<bA���4eF[i�.���EL����֡��^,���*`�UQ���u�Y���q�b�6rQ�yM-2,h��5���`9Y�T)����{3��f�͝3�n֜0��F3x���/J�}� ]R+������l͎�;֥b����36��H�
M�D�v���
p0�wd����Y�r������cf�3�6�\v�#��v�9��3��Z�uh���r\�-X���9o)oE�w�:��35۠Z���%�'79��Z��N��V�� q�h��ˈv`�w\��ސ��Fъ�32��ىI�"�r� c����қ��Xح��o�+e��<1;��e���Q�C�b�����r�5���p�ɻ�جz/sLΒl�-T���k�|�Wbk�wO[S�U:7�i ��)��/$�y�8�T�k2�=�(�IgM�B��۪�Y�&��<��H-��d�Y��Yķ��Z�!�Հ�̜�8�uٴ���fX�CyV��L�,+���9	�rq��v�lR�Ǝd��/Y�np���ƓM��#�3�M�����4ph��8	��Ǳ1:Zwp��9��mh���t��Y����Y�71�lYXy�0!9�YB=�¯L��?�����\�':zk��.U���t��yi%��,_�bX�]v�_J�.��N���UY`��>��V4r�s/��7+FO\�BY�h:�d����vzx�sp�޼�]�RR}��<�%\{Mڂ�kZl�Jit�u1�x��y��E`�#*J�@.vg��:Dj���M��V��+�6��m��c�JoV�u+��!#�ZΓe۠yVSu��V�e+��t����n�D�%����y�P�{gn��$��kK���/%��U���������)5���j�9 U���3�*3��Ve�x��<�.�o�alj�j����R<�f���q�=:-�(������Е�k��&mGa&�ٵ���B��j�Ă�Q��w3�ҩ��M� Qe�p�o���LK�]�ƶuh�F�ռ>�*yxrh+:� E=�>�z��y��.��j�h!]�eC�2M7nN�sO�=�չK9���!�q5b�����9��"�C�C2�C��[��AA�/��:�TI�� �v�cGYR4]��̙�,葳�c��;�7λ(�<���X��70��8����n�m�����/�,�sȟnN���K�Un���,���Ǟ�������7C���������`ήƠ�	�.bY�T��n��u�!E�C9�}R[��QLN��j�6�,$*Mس����PtB��:�339j4�r\��]���u���Yz�e
�E��G*N1��Mn��oۥ����n��{Oh���N���Tk�w|Hm�N]lE�HR���PM����,�Ky�����㷈Z�o�s��T�՜�|�]��Y[��.B$��ڎԨ�Q��c�6����s��٠����4rE�b���뫙�Y�ʟos��!�����on�u+xm
�O9�����革��k�Qwl�0>ׅ��q���͂.=�X-@�;Tf-�>������\w���ٰnBA����&L8���f��rS�ٺWkM�q��.*�{�B�[���<�],Ч7��i��S'�1�5��g7J6�G��ae�Ĭ�ot.vP�5��6��ӎ�b��X����R|�e��vՃq����I
|�v��޵Y��e��I�w-5dR�E�+�ݲ�f��æ4ʭf�2��x�t�$E{-�[w=pfb'�
$dln�(��Tߴ�}�c<�r֍��Мj����W
2�A��r�w3�$��R���w�<9Õ�m%�V�j��6:x��b\�4ܺ̔5�=̓�s5��eM��2e�J��:���m	�-���4��~9'c�9�)[}��3��G��V��ʩ��.�ч3��I�4�˓����ˠ���Z�9��rGk0��"b�O��]=P|g};oF��&.xr��f��QVD63h<�-��-��
�w ���\�u(3�SX��h��.λ"��	Z:�S����/-��}eL�=fΣk�"��.i��W--�U�;��:o����ɥ��^+�Bۦ,���1p�k�	3PJ�;�����Z�r��9u�eei�sNVՋ�rЎ0eݔU&��|�]JZXPP���ɫ:b�J�^��c�<R����S.�����њ�L�Û-����nnA���m�u�v�v��c���-���������U�փ�K���ɅXm���5*_%V�$�]�d&@�B��N�ƹ�uu���+Ț��͛�֙�f�Z���>�@���!i�櫢��S���]^\`ֹʵ����S�b����m�h�[�־Yk��dNǽP����Y�q��A$ڧ�����ة{Y��s�p8�b�=�A�U��B�|�}[j��qƦ�mU�}���/K�W9�
�F�4#L���T��պ�֜Y�Q�~&�;4�Bf�^��̸&w��`�6b�l�r�-��Yٜ�"�e��	/U��UF�Q��F���q��Jg4Q)28;v��d�er{����� A�_Te��B[��_Ӹ��
f�]��_qĵ��<��7�'��n�R�;�ͼ%�Ay)i���f���]�j��9�kabܟ|7��=�����IJ4�4�=ς��Tٳ/`�*Ź-8((*S��W�ܙ=U�X:��k����q�B�K�g{%�h^k�	���|ŋ�2�y�?�"�n���_]�r�f�J�J���B�9k��O:���&LD6����j��J��5M��[�U|U8(�+��A��r��zh�v��f�R����g�ca60Q�@pl��;�9���݂��Hjk�vq.�;�ka�b��:��3)���4��f�Zb�fu�tMZ��!2��`�҇8���{T�hЭ�b7jCjiT�츜�ץ�ӕp�S:�sL�����Bud�xa��})����VP�=�wj�pL*�2��s-S���-�)��F�_u)}G�p��N�>@���}�m��m7B�}E`(x�{p^��v�B�	B��Q�����AS ��0�Ta�+����W�w$�L��C(�͆mz
�K�u���\'��˩���J���Gp%�{�,&�F�q�Ǧ�;�U��W�m
=soD��"�����C0�m�rt
N�G�q�&gpʹ�C�F�����m����u��[Y�!��
t��ݵ{��[z)�5��sw��S����:��ۧX��H��Iob9�]�J����c�b�6'�K���C����*lmLm��t�$�#�N��m�ە��/����t�#[b� ��)Ͱ���"�pC=}��d(����1��o=��n�v�������p����ȭJ&����O�u.�U]�`�d� o�P�,�OV�G��A���՚`y.��jj����2!�8]�yu�N�ۀ1S����8�5A�>�)�zώƛ�upy�h�������]2���6&�\�ڟu��ka��'/)��Ԝ�(�OU����8ءؖ��Ys&ā�IӜS��3E����:�{Eq}{y��� \��ၫޞ�Tqɪ�0�d^aѶ�n�.VV�.��"��7�Թ́[�%e��Y��@G��Rg���n���;kH�宆�I�r�6e��i�Fc\��Ì�ո莵�eufs',��q�zz�t�F�hQ���^6�����M�@�h=���܅���j����p<�|��]���j�ed�[���N�WK�h�{�ڵ��ξ�f���Οh��4 ���T��ӣvl����n��xm��.ΤP�lA��ޚ�b�D�.����8I3����m6��d�V`[�0��'v�I�bQ��9� N��tCqfT1c�^{v��d6_M�&r�ý1k"���$T�cw�wۆG��>��ۣŞ����"���.A(�����b'��3b�m
u�um�5E��R��@�r0���ql�<M��$Z�ݶ��!zRC�쬫�����)�v���W���9+�hdΖ��*W5L�֊���3Et#f���j��-�S�>y��e�`"��]t�5��7��ng<F��b����HK:ņ�t2�t���sw4=�ʼe�3{��X��a�Sr��}��ܑ��6u�0�������搝s�me��Դ�]�Ii]�m�#��:Ժ9�t�s��u�����D�<�h���B*W��N����M�_},�o�\�}.��jV+�l�qy}��pX|�yw\�A�q]������`�%�6靿��\-`���\4G����,Hf[C���jO�Y%G�*���Z��%�8��}h�Z�A���fV�/$�7�5M��^�v"X
Oggk�P��˻�u�V��C���5:�>��Dgc���be�0u��^Cr�\9�L$a�(+��`86	��q�hU��Le���=�����u*B�����p����F�4@ɚ����)�ܮ������m#��mXZ�'����Z{v�fmZ�I8�.Y���n�/d�7lf�WpX,n�l֫i�#%��ĝ�0gf���{��ڷ�$U2�uW+��Yx���x�N�|�`�-�T
Ol�q�Ƀ5���@�Y�J�g1`.��K��H.��Ԭf��v�嘪����6�vj|Ct?��1�� ����������W�_�?'�9�����������}��o����o�>_/���ο?�j��m�nr����$!ϘE�EH�nX�|�� �*3�0���I��q����FPf'�H�,��pL$Ə���!$eKQ"�A��ށ>��P���z�H�c��ލ�$S�0󤫺q�CM^��j�4#ӧ;H&�o5'��ԭ��6yo$:`׹����;��+lr�#pޱ�1]K7b�}Fk<H���+n[�n��q��R_Wp�]�sm����"e�f�"�.�5�w���@�.�t���Z�ӹ�Lb�@:�H�8�<gR`���:6��+;`�,�of�8�^��R`n��P�{���4ۨ�e����cy�t��ʲ��
lb��uɹ���=��`�\���(d�k�@.���Z���u-�gzw,�=IR��x��/^"!Xv]s9���}ʷ..\�t��.�G����1��0���mp^!j�%�V��H�����XՒ&^hP�U-j�Z5�Kb�1v_8��;X�ӥM񮳴]vD��l�����K�,�Y6�T��b�8��1AYoL��v(����w�d�o;f��*�W�9�JFHv�v8f(wU��3FNXv�J$��;��d��3׃9f%3Vt�#��ݮpC�[��@r���	tF���0���:Q���E��y9�h�M3��*y;���2Ծd�Z��n齫&r
��}I�����"M0G9\��&k߻�!���K��6��r��"ƻ����Yuѹ���Y�5��/\�C��i��sꕡ���귃T�I��!����{Ȍ"����DI��Qh�I�!�B_�蘉$Ӊ���Pq�-4d�cR�$�h�X."�n7r)�jD�&Q���"*(�A��0�(d8�f!����d�$�>nRI
p�I3
-��ȋ%`&�q""08ā8\RO���!/���0�(�& �G<s[�2y*	��O5V�5EEMh�,s&�b�b*�j� ��0ID4Ű[LUDQ��fh��
��*��6�&��5Q$[:���Z4b�!��)"
h���4ܹG'�1�֠�� �������*H��j("�������h�Իb���&".���bJ)h��\��MT�M��M�UQ���c�����UMj�
)��"b��J�"h����*�"����N�j���5�*����j��LIM�i��)���*���T�UA�1EPD��떠��*��*"�"%�������j�d��)�����(��J�����78q"����(�����<b�"&�)"��f����h��J��LDǔ����'=^,��7O#G1�՟}bP����)�Ȝ=�г�D\�����ES�a�Q�vGV7PJ[�>�����PӼ��;o�5߸���	���k�C!Oņ6�lB���RD���6�hۮ4���>O�s���IۑI�w��-�{�WKo0<�*j��z��Nh
�[��S�5�7^�&M�5�=�C��ni����`�Ǘn�OUػ����>=O�z. ��o���l#���<K��4NT�nS� x��a%/J�ў���=b���������r{|C�c2^z&�m訲��ϗ�d}vo������6~U�r�vP���Jx]g��Ѳ�pҒ������A2I��2s_g�zXg�� �μǚ�u�L���Y�I?x���2gq��y��2t��w�d`�v6@a��%�$ޓ���Gz6�g[��[�q�E�=3O���o}�*m��u׭?���F\�n�>J߯B��OU�]{f���8|j������{Z��X���N�K\a��h���	a�.\�ͣC�ޞ���9�>X|k��Sj4�Q�G���}�j\��d���S�*>��}c��ŏ�Z:���a�|]\�����f���ǂ�壏�}��^ݛz>q�p��-͂������fL�nQ�G���ݙ���ݍ8vh��wbq���5W\��z��M�/�S�*VC=��z�|��!�s	��d�/:�v��u���xG�\������s3����6|GW�gC���2o��a�:J��jg�*D�z�q�~����˕$�R��?R��A����n�}q �ts/XI�{8D]�ݯl�_�V�$f�f��~ا���w��pc���#8�;��sȫ/w9Q1������GP� ɺ;S�^�>x�>��:���4�ʵKޫ���*�lX�aS�K���o]x�M�3��S���ޜǧ�4�G;fOm�ʔ�	�ixu�Mw���~?7~�Gg�
���X-�Ys|/�G�`�T�w;L`M3�3h1��	�m��Ⴚ6{kK3y�Dw�(tk���}��{��'��od5ә�q¡�	�-���b���'�����Ƕ��c��s��~m�'7dw_Hkl�0��x�Ki��ۯ���[)%�JT��{�HFY��y������P\����1j�7o�]:X;���'�TNZ�w�*����xF���t�I��,8���˶��{IA�����仒���Is�f��Y.�y���\�q��wUN��3&s��c:z�(bɳ�_K.s�m����7�G!Y��=����<h�=5z[����>�
�g]�Ҭ$��[�����C���3Xβב��%/y��b:��ʺZ��|_���Yt+�����dW�׺�k&��d%�yࢾ�#���+�g��̞Ԁ�̢1����=Ng�����>�<����0�iY~���$�突���Z�^��<��ۥ�ة^��e�|[��a��q�sey;��F&����[[&=��mCV)�
��o�ye���e�>t=�U�7�ܱ9)�y�N��&�r�r^EF1�w��SW]�Iw����Q���6�S���3���e�J߫�>���^t�e:��������R���
v��}c[-ڨ�z&�o^��"k��BɌz�4� �|�W�r�q��T���jv}�ﮨȁ}ŗT�:b�:�6���B���D�3"�0H���P�>������Q�T�p �k3x�&4��5���L�N���*:5���,5O[��Ѷ�Ge�_���v����L�R�}����;7t��
^w���O��4��˻���y���q]�>�su������Q�3�{{n��4� P5����c�����\>��V��*�/�;9�7��I��K�]��sb��@����3�f�%��7FP3�(�D�"�l��ō�&��d��ڍ�s�O�[���仓�m�p����S���ҡ���D�y��$�9�C^L���#�4���X\�+�;�=�c��}Iݡ��؃���[v���3��G�ñ�\���=��	�Ϳ7�m����I<�=�sd^�^G���8��ly��[c��"MOt�ǂ��mp^G��;5�|_��vՋ�}�=��W9�z�>.����V}	����_\���x��ͪ;ogy����FS��g��~N��	����!��5o)�;����U�O��xp|�U0:o�$����'�nr��ſI�c�����K�r���<�����M� �R�e_u���ٹx ̫�ͫ\5�VZ)��i�.w����)��. %�F��Z�0�Ám�vI��cON�u;s&Z*�,���S�/M!��V����,�ާ7B��&AH�A��{ջ��X,��䗸�h\��P��/�Qz2���y���{ۣt��&Jr�^q������^&�Լ�K��~��ߑ��,}ꙟ*�c�kO�����e��>��LL��p�A{W�u�9�EA^�k��+�߅s
�ޠ�]6��:��nN�w�z�z����������)>cG�튮�{қ(�+׸ۨ����8�
�c��f��;;~^�G���^�>�v�т"��Y8��1�^L����u��Ջ ������įq��A�$�\�m��#��"Y�^p�g�j�"	|,m��rW<?��q&�qYٕU�v��>g5M�ngޫg�
�E�p06ۄm�{v	:�.���]o��{����el�\�[8�3�8� 6֊�7���'dz8mhs3�l���<�o�[�.Hj�r4����A�}�}���g���*�������nJc�5�8��k$�^^�޹C�L˾��^���5��Q�Y�.�vv��A��)���8W�G�*yL�A��Ш0K��l6��q#v��C�hj���M��]���@�p��R�I�>/ge��ʊ
.E�sx��\8�ֿ�;��P	�No�'9V�����Qxl���FN�� �>�0ñ��i�'�tO�3����^S�U�l�!�QN&OL߫�ߴ���k�I{�O�<�W�i��a�pQ7HW��r˦>�I���xx����I��W9l�]L���A�3=sgy��c�#)�=�b5���z�nP�꺙�C���œF�hx߽Y��o��=�c�o��\���Z�K�Kk�k��)�g���A�JH�{��E����R[�&dTcڹ�N}����t���0���	VF\�7s���q3-���w��w�N�X?W}�t�Y��4���s���^�O�*�w`^Y5��	�$o���Ҏ�����鋟���!�U��0>�̪x}�Y9č�|A�n�����Ժ�٣'t�3U%�a�y�U�p(qj}f�|{�ou����ɲ>�]d9�M��$���.��]tR��o�V�4Z�gh��N����}Rݑg��l�ùx���2���nzb�:=۠}�a3�W�EO:��ܪ{#&�}q>6t�l3��ǒr�����w$k sS��ɰ�U�*q=yֶJ�AL��&����	4dWE��ާݢ�/AVW���a������f;��t��y�sq��da��4����K�G=MP}��:�Ǆ�G��Y~�ޜ7�¶��;�"�|����l�O3�r8��5A��@k�;^q��z��4�q���w:[&�Y�<6��c��s�����^M�I�~��{�4d���ޖF���7'��"�d��/gcL�<Ǧ���T��z�P>����8ܩ���}�־���t�,�q�kȟ��ͣ����>[gKg�7uzT��it�m�1������6�����Ϲt�{�9�
�7���h���fF}�O5�*n�j7K)}Jr�"�����1�r�>>�Y�Y����*Ӟ�g�֟/������ǵn��kp<+�*���Ox �7�k	�����W�t�n����u�kjM5we�t�m�����yM���1+��{:����oX�|��]捕w2 9;{�*�����-P0�-U7e��ׁܚ���ϕ���T�W]��-|/�{�����¶���22uC�NX�]�������ԡ��m)��B��F�c��.5rtw(��J�C=���O7L��I��˙��{�f�H{hwOTݘ�?�W���� \o{6��^�<�v�	�7���Tf�w������zd����pp�'��i�k�//{��2,z��x�}�X'�ݍ>�f��P��ȕx��a�>������p���}Nv�H9^H1���'1�ݷssO�(�Bp��^E�Q�W���TzE+w_�sm����r�t�@����s�K�g��o���A�^ζ��l���.1�#-�G��d6�h7A$��2M6�b�2�ۯi^���5~������a���1���^��$�8�kɌ9S�]�O��y�t���<���VfO�ɈFs��We	^{��c�����l���W�3%��Q�#�z������d������#���vb��=��G��6.j��DL����1���'3�F��:��*�Sw�6�i�۷�3n.�w�Grj�m�W� 3no��A��/�L���C�,��\b%�9�Ŋ-�U��X�e�P�c��u"�st���.ᳯh�����G+��W-Zd�39+ыDu+c�eǚ\ˈt�w|��`��h����Ċ�&8�� �}��3`0=|�٣uTX�Aӷ�D�eh#�k���w9����wI��ـymq����#;d3^yb�X�����#$�`1���{��I������{��yQ�[�3V���mu���چ�[G��e�����=��U��?X�����=7��6w�D<#S�|�v� �����{ۣc���}�d�8���:R��w�?n��s��<0�E��k��r:#�/��ܾU���n��0g+f�q�3Fg�a������|	"=���I�lS�
: ��vNs[��s�=� y�J��E;ǽ+6��=��o�\��J?J�%p@�uO����ߛDV0n暎"&�hE���>㗜Aۘ8Oi�6�5�ǂg�3W�ؽ-wx��z�ty߹�H|�hFF�p5���fM�c��o�إ>���:M\����G�X����f���g�:��tx���?I!�'(����Q���W���pX�!��]K��ʽ�(c�MCx�J���_G��Í�]A���r����x\�R��۩y���I���lY�TGU�օŜd�Н�oI+0���4ٔ�{%p$^�gg���x'��C�Fm�9�v���O��7F8�2T�5t�w�TڬJ�딩�S�G@���$zCo}=�C$ߛdω&Cmh�sy���/�%?<��+u돚b�J1Q���3nI�^�\������v0�%�wf�gu瀞NyM#z��~*o�E���<ߏ�������{.�V�2�l��$k��1yW�~E��^k�t'�O��:�q��{�hx���މ܊�5���tԒ�wHxن%���>9�gcz�7 wsmq$x;[;N�4v��FS�h֏�a�\��fѯtG*�*�>o�v�fQ�o˃�FD}Sص�q����*�Ե^��.�my�m��5���fQ3��'uP��۝�c�Wl���s���>���z}��/?�����{���g�������z�~>�`Un�zqN�lg�\Y��}b-I��n+���Y��r�K8̭�K��u��l16;�N�ٕ���5�:����n�^�9���y�,Ԏ�.�,���F��� ܱ{P��J��c��|G:�YV ����h�qe&��wm�^�FUL�+�"b�/��A4��^���髵5Yz��N�.�7Q�k��94���[�i��3[ڟS��Gb�z.	�0��Ѯ�5�T|"pn����B�G���2�e-[�A,����Տ�c�N0D����w,F>�Ѹ���M8{Nt�td��]Yɪ"l�,7�(����o�e�����!�Y��"[���m����)e�U��"4�t��9��٭--<YY0v��.v�����/��i<��J�ɔ­w��G�@f�i���K/�tHD��wnlǅ�8+sl�e�Rr�$fμ�ˏ`��}�]ȧo��e�fä\^�Ԭ�r��.��vr)j	wۓ2}4KĶ��<�R4OKm��q��r��a��~�R鬫��$����]i��]˼}�	(H��­��\T���sjf�h⥁�tC6jB&�]�3��u�������R^��$���3��}�1���ɸT�r�
i��ejz����e;1m�VP0v�D��]��G2t�ӭh�lX0Y�:<�z7� ��������٪h�p���P�#�hj��>އWNP]�4��u�dMؼ��6K�� @e��Qإ�k��C��� �
��Tj{;�5��qڴ}7jW��<��ۇ�YGG9�S��v�1����؆�l]�2�<��*�\��u�ù.��s�'�2X��fu%h5��T�#��Xy��ӴW]JV�.=C]����S���r�bm=r
��ւ�t���`�t��f��E^�]vYB잒c$��~��Gtw���^cyX�7���t�B�XC�u1S���|��:m��e`˂RP�Q:�'�&� ��4s�%�������@�i�[<5fku�����y�J�7e�
�����U��ù��hz�v�\�o{3+��Rj"K��k�ַ����:��v� A�t̬v�=��ӊ������K��A�w�v�+ܜ�.}ρ�V�=���I�vn|�3t/Zɓ6>[��G}q�L	�t�[3F���&���\�u���+0���{u�G(��vQ���g
q��i�B�fƲ;���v�ŷ�T��冞�Q��8X1K��32�9����cU>��z��R$+[�b��wȓ����V�ٯ��B�ՙQغ��PH�\B�S�͈ʙ���ΙS��s���F�w�r�γ��-\�EЧ5�vc�,MG�6�+��س�"PBt�`�h$p��,Ct�a{������4��4םy2�Я��y����V<��J1���ֳeo;ѱϣ�/>j$���������LPMDA3M)�`�b
h������)�(���
�h��f��`�DUL�D�IEE�E�*��b ���+lV٦j(OV���b(f(	�cT�4�Ps �j)�*��
���*f�j�*��f���TUQT�L��USD�UEE1QEDU�SD�@LW�nMD�sѮmE1U��[%.�"*q�q��Z�kcmZlK��&6�QX؈�(Ѭ�7�nk���6�M��2[Q�a3�"������O2dg�6V�%N��Q֍i�j6���gU�h�œ�5�U��9SV|c�-3Y�Q3F��Mk;�f<q� �r���>'s����F�F��clg3��G3h��56(*4��ob<Z<N��I�h�Z��j�2�&���y¨��8mL��IDm�gW3�N$�1��k%k14�Z-�"�rE�lr8�Dljy�c��u��W���w��ǿ?^w2����AmĶ�N�vZI=6�f7(݃���W�[];&_V���P�k�.0��Nn{��,)����M���<6��L�$n�0v�wA!�g��>��Lϼ�Z�_3Mu�~�MXa�XԳ[P��2��X	�=�sО�ǵ���4��i��(�px%����o&Ӂuݱ���q�釆gN3���W퉟�R�`\Y����<x~��>�z���5xjJ����Pd�)�`�:!0���Ǖ�7E��&��ǫx�"��с�מl9/=;>�V0]s�^��%67���e�!���΂��62�Ms�bI�1� z3�oV�^����/K1�{ճ�C{�h��5ɕ�3��F�d�N(r�d^�Ji�%)���,<h��>�i8<�>��8~׵�3Ιʅ�{}��M����G�<��]'�)Յ�)�$i0�#�y�ϑp�����^��a;�7+Hk������A��K02;$�����4�ሤ�`n�J����$���6<�:ɺn޼f�Z�Fe;�R��!0�p1�oC���@Lpm�����a���/\����R	p8��]D�n�T����oX�^�?	�at �`���M���@����ιM�ګZ��/8��{�<CqS:u�;@�9���J�7(����{�!}�"������J�t��f���ɲ���&\�����KZFIuyy��7�Ă����M���c�H[�b'{��t�]$͒��i�3t��)d��.�;���f_?�����#uzN�Y&��D!�J{��|w Ļ��ga�d0~�vOǦD����>��I|��2�c&o-�f��Lt�/�`�u<ѹ���9AQ� �+�H�@�H�^?}��瑙UXf�_p���F�D8wQO(r��%0�/�^���u���_�8���̂�.(���=�S��nc���ws"�����9e��w8Ў���pm<x�0�����-A9�Pw��y�� 2�[��6�g�����H���66�k%}������^�.ŧ�
ޗ������w�I�њ&����{�4�f��N?~Ys���>�!���Ov������f�������)�2�����"ߚ��E<^�P�4(a��OL�蚹�u�ح`on������Me�cu�h�[���P���Hj�Fu�6 �[�-�<�ӼNIݳ[æ��������l�$7l����i�ɯ��OAd	eI�z��Xhe;k�l��Y�gۃ�'�쏭s��qpc�O;Hݝd��<��,}�'V���R�*�
j�Wӽ���|+�e���/߇`y}.�5���%��+Ul�'(�>����E�^��l�T��r��O�C��H{b�p$c����Ⲕ�'�D�/��U����� ;wo)��pq�wsu����ۦ�$E�`45�{����4�q����ʫE���W�.jHf�Prч�L
��*N���G�;J^�~T����,���q�%g����>��@6�r;�S<(v�lj~��=��%:���j�RN-�"Pq��-jU]��D�`��hT=����#D:Añ��n�s�Gu*L�8LS�,�~,��nm�W<-�҇c�[��Y}�-��r<#�!��r�	�G<�����P�F���zNU�+��&��מ�u�%6�:�09�ع��O9Ȟ+W ���ڠk��&_���ο`�L*z��2�·��o�K
�J疫W)<�*K�GjHO��d>;��`���
���0��֭苴T���Rss�BՃq��*�
��̦º�����NƸ`�TA�jz0eT��-sqi|���1L[@��׺�smg�򰦕��/ҹ�%ߡ�¨�{�]��A`S�������M�r�&�C�K�0��f^Р���4cx���,�s���8��I�k^�(vu���9-]���m��ShB9[6����3�@�}���	���~��fM����,� a�-�Л[c��]Wz���n;Gs���u�e�@�lhtg/:����0���I���d�i�@�P��4!���!��5ƹyv�k]��S{�{2�o6���E`�cg>��헽��W�qJ�8)sV�y-s�ľ���߶n<�NF�nֲ[������1m8���3�;�����H�k��D�Y�A���.'f��7�Dӓ��?�z8���~�S���0Hx�2	A(��7'�gm:"�W����cC`38�`L�_�f�if�6�J�f���k?V��S��͎פ	x��F�r�J�!\�y���-�W�b��tS;y䪈�xN%ݚBMU�5���K!�_���u�j1��ӕ-�ZT��c ʖ]
V���� y�Tee���f�2��yB���8f���|���?�=��o���~F|*
N,��	|�������Ў��bT�U穃Hf��XAE��8�(Lx$'��CH�b�j�B����l�NK�Sb�j�#%��������T.�d�=k�{z([�PqM:A��!?c8!�B��e�]ӝ�jzx>E�uTӳ�>@���9�Q-�����$�0��qA���k`�a�'�	��Og(��j�����A���N�'(��]0�9T����W��Cqs.[]�kǜ=0۞:J*���m̴��rN�S@�YP��E�D�q=㊺^�E��)�IoCsP	ĸpÛ����ÝY��N ��G�>�iDktlIu�f��tϱ��*�����t;���$��/�k?X3>���s����;���̇,ʃq�G���cJ���r���.,�퍕���r���kZ7��¼�yǾҽ�t�(�<���&|������N��˓����j`X]�C;�=v�	���<٦�H�U����m�,�{؄�����v���1y�A�.g@q ��
|àz:��ښmW=E���6�I�\�5���<�<>�5����^gç�ձz���p�6��d.����ͮ��a�q�����zW���Q�����X�d=g,��S�S�ׯfz���c^1a����Hv����u����s�p'+WSQ�a��;ݚ:W�MNPFC��}(�A�c�ô��g���-���D��ż.f�Q֝�:%��C���v����.��1�e���z�8�I��F�ci�H~,�����V�C��Mq����~�[�m�����&���[!�=	�{9���O�7M�M�I`R�o).��ݗ1sΞiԺ�.J5�<��O�坽ZX����ssS��{3�K��n��Pd���l0�^�`�&ci� �;�al���C6o�Ui��
E<Yv�(���_���lN�U�E�t�}D���s��39ÆС�(1j���ܣ8��ݸoV�^���xA@�K��Hp2"�&̷��j�dZ!��ЍkF!�1,���YJ�]���ơ�l����ņ����I��9w3F\VM��P6!����z�_�r���}��P�V��˩���v]���7��?-)�0,�8��:r�3�f�ǌ�#@gr�;^+2'��g�cS�l�s��qs,�]Y��3'{���0��OZ�Y�̦4t�e��˻���)*����m���.NóT9a�n4��;h۷<'I��"S��7�#)���9��.7��\يN\�N��S�.�}^@h�f�����`����K0]�a�wQ��Eg����U�\Ø�,:&��`��	�)�����B=�&�rp^�j/gT� �&�z����l���b�gF�䲺|\���[�#� ����a���ߎ��� z����8{{V�?f�R,��TsrS^��fqmy]�q�X�����T?,Htq#�
"��5����}���huH�tެl�����2�6+ľ�}�sg���9�I�`\�[Վ���T$�v�;��!_���� DW���S�o+����'/T�mC'5��^�D�@�k-tz=;Ƣ���`HB�}����r��ɞ
�8�X���ccH�M��W��s��2��S���-�	��_�9o{ys�����'�[}B6��+�`���r�
��5_o�R5�w8n~pК&h�_��;��wKs�z���bc�w���bC��;�_j��P���?��k��i�5�'QQm��t�2̳C_��jk�x¶��ǅ��3ۥ�d���Y�:�G�.P��%��6/�<�9��������]�hӡ��×[��u���R�_1��]���(RY;�X�"��l9���:ՠ�+Jl�Frv�v� r�YTS��6ߩ��w0}��>�gw4�A����O��"�l��ulێK��T� ��˴��Zz�-?V�I<bO�ջ?��Uϫ��b6�A�e\e�E������� �jb�W$2F �}͜e^�Ξy���0:NiՍ�O	���K�S��֋�\��D��i�NEcW�A	�� �c�d�N3��|j~�xsB�3 ��ݺ�i0��檇Y�8�h���DN���D�l�֯�6���be�`�-S�*��nN0	��;�{���#A�vp̦^��g��]C5d�NHܗn�����"��Jui��v��M�}6j�v�t�n�*2m��r ���э�DcL:AĈrH��n;�0�;�Rd�ڜ�P׵-����!�;$�p�^��E��q9@؎�.͔��m� �cL9��S �y��	dޫ��S{�zI^fLq]�r�E�ћd]`c�qsO����ٹ��=�x �kȇ!��yy��_��4�+$6���	��zyW���O��-V���R��x���m2?�=�h�gO�+�A�t��V�۵�4�* s.zj(��9B̓q�.�TXW�t�)�u�$��}n�(U/��^��U�y4W<]�;�&����2����|�Ž��p4!����}��c��WA��C�o�W�\��c火S~��A֏e֋�tk� �[�-�x��3�؁	ҙ¬�x0*�w��c{_-C�\ͽ����*�f�ð�׏������o�{n������L�4�>2�X5 �W��mD�q���{	Ao���9��JUKU���2X��t�c�l���}�l��y������潵,�s����J���ָm�u8݊�3"3EV*]/å;\��{������W��&8y�Ɔ���^T$�_t�s{����UIu����qx��2����f]���9��l��^]� `L�/"S�x/_l^ShxJ��v��m�׎�� U3ǲ�zw�H{
��j��L��xe[���Ǆ��V"D(�����ْ0�n	u�"��_��,o���T9G����n���7�n޼gm�mt���-;W���jS:���:q~����5�WFL5�{J����Yt)ZTy÷�N��K�F4��MK�.�+�a��ކT5zm�M��DƴÈ�i[8�X��njJ`2ѐ�7�w�e4��V�j����wڴ��h_s�[��3)YE���d	�	ಣ�	��{�N2n���/����������8.n,�_�JS�P�[�U�}ǅP��� Hql� �� ��W�����4^j����}侴���)�d���X8��C ��Z�N��0��\�:��Ĵ�� �HS��ijG�e��7��dC�I�s�3�5��B�X|1k����߶���d4���weY�ӇM�g�rj�V[:��7��W=wz�{/ٙݴ������'M��V!����^����c�:��TT�P~����О���H0͍��{0��a\՛ٸ��V0�t%�c>��*�(��dQp�Qu��L�oT7Q�NZ��k��h2���Ʀ�;L���ŝ�(dE�ɧЄ�	���y��(➛�v(���T X�]&����ּ��������S
�_u�t�������):�����r��uu���ד�y�C�u��FN������U��������?�H���s�������4گ��Qke~R� ����MRr"b̽�B��ۯ=˪~m7r͵�l�@A��ৃ�(����D� -߷�NWc�]�b�w�C7qG��GO1I���dzu����k%�ы�d�f�\>�E�u��j�����wk'��E��ζ�N�6�BhgI.y��C�g��y��hv|z�`�����h�):m}�Cx4�L45��6^��f�Y�k������=� ��iW����_E�����7�lP����;KL��~B�Y�9h����O��z��ǳ�#[������}%����Ayǻm��n���Pۊ`~���r��u����OaP0%��[��~��ߔu/�WjD�=����8F�$8:�m�#(����:v�3v�&��&��S:�ӗ�Β��#ٚ�Нe���>�M�ޤc����{��BQFj�+;A[t�O�6�)�ʯ������n���L��]��n@���6�ӯ,��5*�ԁ����\��3�R�nod�(��`�31v�6Ot�ƭ���Ĝ���6����{�S�-�â�L\zxW�V0I���OB�VF\�>�n��p��^@"����(2kJ%?zQ�aC��}j�?*� �����~XG�'N�ۤ.�Φ�BHu�dp��\��'�bY'���(JSN�om��t�=���6vats�u����"���yٶ�0X�ivA����>�o&VH�IMMގ�� �s[b3��"���`.�y^P3���m0�Y��,��৲L8��4���"����E'��՜MЖ�Uƺ��]c��-�df� �}��g�Ǚ�mLpm�{<�^��0�rt�Vo[3ӫ3dk��\�GZ��G@<�y�j�3L$�x?O�E�2(�oH�#�*��?q�]<iL��v�ډ�
o�cZ!�ySZ�%�c���t�����wn}ga^C`7sߡؿ��V����.�λd��G[�*E1�*����)9`,�M�*�a�]�6�Cz�ٶ@�`�C�@p�}?O������<~��z�����~_�_������ؓfDnϙ�vC��ݱ�T�T25�:ۼ�H�K\��l����N��k��n뜺�lX8

'a%`�moCzּ��Ԉ`�rU�E��z+8Fٳ96������b���ʔfbxK:C:�mX�If����h�2���&�h���M�SӮ,kq,�?��u7{�4k-1h�U�%��j�X�S�b��N��<
��`�LǶy�'G����kif�Fq��3Xz��QQ��-PN�����U71)����o�1���t2���*nu�)͙��u���*_Z�:̘[�TD�Y���8������d���{���;�ݖ�6OO�S��D�`
���:�#M3��F��L��hLP#Ӏs�Ԯ�b��9�4u=�%��.�=z�L��5ڎb�Ӄ�J1xOx�ڧ��m��`}#�y��K��4P�8�$���n����-�J����YnC��Kd�n�bw�BKY��d)ec��� dL��bi�*`2��*�[�ٓ��]
]�ݳ��q�����{�s�v�J'HV��3��̝�.އȂ����������E�l͈vnc��_'joaF���yRV�s|A�zX���V�muu��,�K�����q�*���{-�Fs(���l��`Y���d��]Ļ9�̸/Qe�\��=k�zz�w��!�:Шəچx\����P ̱t�AyP����0�(�Tbv{y�Q�vN�7rZ��NJC;�h�"]VB��:U-���C{z9ke��Q��		K�[9V���f��]��9���=x�~'
y�A�{��};�
�V�2n��[e�X����n�|�x^�I3	}5|���<�̑
U�'=V���&f��U�X�|�8[P��-��3�^d?v�XTlVa�������^d��0������ԯ�ۈS��m��`T�w���E�ܠ4W��%�����7k9��4c)�W��a��5�k��/��D9��V%�Pen���3Fs\���n)���!�Ǿ��)�唰v�;qkr!�k.s�Ճ*�Za}�87�v��ףpk�a1�}c	�v)�*���*�A2FV	l�]�V�/e���ۇ���/��]�L�N<�҄��ڞ.L�)<��+j�q�]:��e�.�Ji�-˚�ȣn����/Z7\�(��t���6f�9O�fр��=�NZuV`���j�ﮙ��� in������Gu�[��,�u/ʵGJb��j����Z;���[yO�6�W��R��w���]��C��n<�MVm@��y�2�p9K=:�8�� ���Z��j�q����0l�7U��iks���ik����7�4.o�L�*1u5��r��X��к�F�z�e�|ӱ�v"�4����\�Љ��o+Q���_\Tc��u`���G�
�,W.�WoT���'O$����R%ϫ1���2�`�ύ����~d�
5Ci��'��"�(��.Z$��a��#�'Փũ���
<X���E�9�-��*���h�<��t�5T��`�)��h���K�*h
k�1B\դ�Z��*��u�Ns�NO��DQ4ղ�`4��T�35TUQx�kQU�5D�ؒj�i&*�%�����������j����")*`�����U:�UUF��AEPUQL1ET�̔�G���f������S�)��v30�E33Z�QEQSPL�S@DU4�QMADMU@��b$�*5����j���
)�!�
�9:�na4��AQ�`��+�yr�.�v�G�g�к�LIZ55��E��KQQ��(��Ө�ZZm�#KTtQM!Z4�RPSA�֍U'�@R�45Q5�E_��9�4) �-��$��	���>>��.����bx��ɦ%:��-m�iǑjip���5�2�k;zܻ�ȍ�b��sI`8m�g"r�V H,�9�d(T��%K�a��nG#78sǏ�ED~��_&�'��H_��D�6[��H����4�=�ϴq�m�����WY��j��z�;sz.t۪~�HpC@��|������=�C��������86��0�qh�Mz[�	��)�3�mNw -�˞ø�xgA�;P�����X��ԍd�oP~|'��w��3Eٽ9��-a�=cO-�f_�;["��h��|�'��Ac�A���|@�9:�	���s���CrYd67��n͑����jf�T�vJ)�m��O�z5����l�S��(!���G� ��|�X��B�O�x6[�AtV�
[)�0�&���A#:�C6q�8�t�@�h<��5��q~ʻ[�+���.��ޘW�nB뜊ƭ0�}k��  ���ʂF���v>5x��rު2V5E�<^�co3B��xT��.1�S1�Ӧu�Td.z�,{�1I�z��H�r�0� �hm���m�o��w�u,�EÛ|g���
�{�@L$�;���@����	�{�齖O�<Z��+u�Qo����3P�ϥ�;��0���xct��b_�e��ntCO�z��m�)�11vR�&.��'t���n5��
Qn�hU�ǫ��Z�}Q���'��.����Ȼ�Gp��
�/�ޥ�gȭ�����}�A�f���Q9o=��䈱�o����K3���U�N�`��n��7V+g���(
=/���2Vc�[4�v��������<�3z�J����t�w�<�_<�N��&:p�x;�0����>�'���#�
:.�zz�-��{»�:za���I��1Ly���y�i؝~�3�ˇ�A���#	�Ꙅ��ܧ��;�/TtG���<�5<hR�-�¨��-B��O%AbB;P�Bxwf��|y����g-N�ZO?h���S�R=$�/<�D��d�qD��
�O2�S�U�����˄�o1q*\:��`��X�`�H��1�ͺ3�I�[�ħ3�{}	=��f�2M�z�F�˘#v%5k�wR:��f��0��f[��O����d�3Tǝ��/�Z�#���m�wh�8Է5���Pg&;��h����߲a�'[�{ �ơYF�O"q��^jf$��Ł<�w�=����Fhv}@sW���7���3�4���ͳ��e���P{.;{�^�G=�B2�1��� fE��^= ����Pi̻O�^�z�m���v��[�B���C��b0�����5�m{��7��yj�AzJ�!�Ϛ�g�ʪ��?�m@��'�eh
�c7O�yf�a�/,c���-0�}�^�Z��
ػ�����t^���Rd�A�d\b���U%���i�N��xY�\��!5$`�%��1ХX���@6kV�A��V�˰yn�8��)���c��b��v�G��� }�w��Q���@�q_(W��;�B|��ʿ,�����KcW#!k߰���.�.�İO��Q�&����ۑ�����}ז{Bc`�-~��Ҷq��em�sS�	��v��6b#0�B��h�1��vȝz��w�;�fY�Tpy	�e�mϸ7pe�"��;�Muy��HE�d�-��^$���SԤ�q�x���𞅾;�[&H>*v��5�ֺ6��*U�C�ds���t�v�肝w�ĲN���XIR^p��Xh|��z��x;���gƽTx5L��l0�1kD��t;"��3��@J.��)�yoT7P0i�D���9��Q�<R�m�L�!�Aæ���Y�t��7Hƅ;JQ�=/��Z~b��z˓���ZZ�^�^��֮��^���L��y@`鵤E���ttIu�D��	�,9B�F]<�k�λ3�kW�R��o���r��K��.T=�q�T�{� ���×�_�umM6�d�2Uom��s�4RY�د7p�Vr����iA/r��q�&�Y��-���<9>�}�:����1���ޓ�n�/��y�î����C���&e�g��Vt0kM-�}uqa)�Y����M��K� ���ـb�u���˚��7����t�ћn�.�Yֆ�T�V��9�jXxi}2r�[6���)�kfIe�\6Gxf4�J��=�3�\v�U�����=��/��x9�Cn��E�K��ٕI�����F}:��fy��f4Xgc>0��Te��{Up��.��-s5��C�:ױ���`;n�J.Yx����-���`:"طPwby�|�a��fE��w��m�)����h|�_6�5��h1��X�۹���@"}�Ӳ4miF�E�[{'�v����~�魡��|����5���By�+�*��p[������<,A���i?H&���&�?����5 ���ʀ�-3��Vg���Ϟ<��ϖ�0̹��و�5�X��[e��ך���ܖM�-@��6)=��y�p���E�.=8n��h0~��w����w���]����S�*+�u	��FPd��Ji=�3�=��[�z��t�'P�ֹD8��j�z/p�:0��7vB�y��N(bY'���+��I������ΞA�����mђE^�F8="��@<�]�2a02;A;$���Jt�<b%:��)�FSSwkSxh�~/8�joW�t��r�<�3[L%,�SM���guI��RzU�==����q]�b����C�u
�V�&�ճgY�H�w��^w�[������I�I��+SHv͜(v�VF�{}v�ֺ1��D[�{e��+�4-�\ԃ��p�]�.�f���8�|�K��b��mv��P@7�&����}�}G��~�{<ƯN���iw��}8��{�<�c�l"-� �z<�Bm���[�^0L�����3�Ej��-�<�t�/E�/R	}E�����=�.�;#�?=1�BL��X�)�������`��[��8�f����E慩���砟��v��dG�u�����߱y�R��ڵ��;T�Zb�(mP���S*���5l�t���L�z�s� �K6VŻ�l��[C��;�<����]Y�GKh\���wf/���k8�BՅ�ux�k-{������e���(8Թ��V%U>�pri�{9	��	��`��h�ŝ���k�|��B;�����0�-�K�D�/|����m�b8GR,�|�nnj���x���C��_lmH�J��7>2'rJ�֧r�%M�͍�r�\��2��w���=�ߕ}�[��V������:����riľc8xO'���Mgsdp��儚f���%ڂSl�r0�����?`$�1'��xE�f���Jm��Cgn�k��zy�j��(8�Y���Y4���g͋e����=;�0����m�`*�UA��Uc�<\
��pu:��k����{VSQ�p3ײ�i]�_͢��.��ӎ<������M݉"?�$��~ē��ğ��to,#�G�ȇiT�EW�0jc9n�@�&�4 �<b���A�O��u��#Dڻa�v#e����� =����1��)���?��� C�=0�����"��j��X�'���H�3��ƍ�\�8�]:�l~�'�y�_�0J����Ü�P�9�igY5�\�:!X�LRukU
P�[����`���G#����2��u�j.W�1�C��sՓ	;nC���M���t��x6��tzY�J�t�*e'��l'�-�P���� �}C ��Y�3Yc��jb�꾩Q��C 9R�݌�&*��RzH��Ӿ[�	���F4�r��-!�wZe��Vhx�!�
�\Cn�L2�%=X�N+'�`sJ�yG��ٹ��=��+�Iv�T��;������<m�>�I��):�O*�e0� �yj�Ry�T�4��0���^w�jط�b�N�������O΃���`��bn/S�\�H��$㋰J���G2�ְCf�k����t�SD�l��Z�����YO�>�4� �c��tg�X���)�w���̕Ϙ�s6w��G-��^
����&��a.�s.�W����~^��O�E�1�j�9����u�̩4OV��tԷ����4����Ķ��EYFm���V��E��?E�#���}�)�e]w�1s3�����u��Ɵ�z;��I�C��F�s�z��޲�����kf��(R߱�պ�ʻ�cH�4�F��W����앙pW�諭��|���0�V%��z�0vf�@���}.�L�k�H����Ɂ��u�J`���Wmq�s;̡�'�m��E�,�p���
ėj�.�^��v�tE��:���yw�	Q%���3�a�r�s�z�L(�m=��;ّh<P= ��?����c��<S������t���܃6���>drx��zm��7��D[O��^��W#^�};�? ���L+z�*r�݁��pF6��a����8{��|��cW\�My�jR=�6e>�t&�V"���E�U:�އ~� ��]����	=�4�:�tS<zS����t�G;g�βV�K}��3�D��-�e���0r
O??�Ԟ��ix\60��0~�}G5XHoe�製}�����O#Z��Jei�S� �L(*El_����׭��$8�h��xF��P늆���l�T�m�送y��}��):�1,���tS*�J�
~��u�_0F<&R�0� ���!�;-�" ��z�!��@��&�dQtÔ�.�n�d���8�~��Y'Ay�mZ���کZ����2;s6�7{X�.���%�����;�Ͼ��)��w�·�*�S������Vj���Ns�ui��ZM@�CT07W'���M�V�7�½�}��0�	w���!v�vv<�ϭ+�`����7`ac�n��NV�c� =�&������HI�`�碛�p���mf�}[��`&�ƅg�֡�W�t�Qi��E6��ͩ��*�*~<�c�[g�~�׍y�c��ߗݿXA�<U��l�u`I�`X��ad�k��������or2�%�U�����4��8x܀��a�tz<�ֿPښmBM��%��0��������nbc��!˥s��ʢ��|g޻��vB�@A@p���.�9���3ow9u�j��|\���L3Y{�˼�Ll'�O[�y��֙�j=��P�Q�`�Ck�A���S�o�8>
!����^�w��'a����"�Q~���!�@�%��tE�j��k#]V��٣�n� �Ͽ[�1�i��B=,��޺DA������H}Z�c�Ϸ[���^����]��M
_ZQ��˯!	��!�ZD=�NޯOM�����Lќ��Mf�Ӊp���/h�3�a�������Af����Zfj�1a�x~�b=�����Ϛ�L(��rw���:��8� %L�~�(2��lQGj<�Y�_�?��S��:
I�Yb����ͪ�_���B����-�V�J<��nlr�'��'_ݟch��1,Lǀ����W:9wݙSi�!�����u9�,�Ѓ��^����"���åXN' #)������R������i�H
l�\1��]@��Bz�l���������
UJ@Z G��<=�[�͊9Qk�Z+��}8Z�0����cQ�7�7���xeMC���{�gXQ��z�o�[��b�Z�=�6��E(;;��!@��> q:�A#sP��^'��+��5ߢ7^6�՘�gų_8'g�I�'����sȜk�~����܏'�$���H�H��sP����~ں��ޙ|ìYFd�6=C���C5��JY��,��`�vI��F�}���UF����7�E��|+��a�^&0� �}��
A���86���Q~yN�ɝ��9��wS}�P�5o_���	�����e ��E�uf�O�z�q8��6�G4�t�s���34�h�-9����3r֮u��n��kZ��/4�ct<�w*�ćO8�z��um����W��VW"��wf�<��Qs��dյ߻�'-kL��EX'��U,�C"�ٵE:�QL��g;���!�X|O"��z�.��0_�NеaD�E�Yk�=>��j+��� ���!�e���镲�hC�c�jA�<!	�O����	�t�YƄu{$�ߓ����i��d��c���P�q*ݝ}򯗔�nl�伽��)��{K#74�t@�2���+jn�l���_|�!�t�NS��#��j\gee#)���9]��\�̔1*{��Y�����ۃk���^�����������|���Ǯ{������@���R����
D"�*��y��}{�~>�s�t�?���nn���;�gg�����X��ԍd��	���n��Ȭ��|�u�el!<bu�x�v-#�q'DYz�m�׶D���~��h�昘I��`����y��L�.֗��ي�O�,�4`=$�PJm�nF���?y��C`����'`��Zn�Py���ݿ���hzc�Q���حja ⅘A�P*�H�3�E��-�9��A 0w;��f�`�{G@���a��TM�F�"��T�Z��'����$kY�bMMX����l�B�4s��zc/P���Aqub%8ʘ�v��u�>:�ވA�=��o�Pܛbi�s:�:�ggn���;<�Yod�Q��sB�=BL��>Re���]�r]�O�%71�u.8B�;���]�n�b�_�(еaU#�0A�a ��m�ny�[zh�j��O��d����ELd�z���Ͷ~���g�}�#M*L���X�I�&A1Ӆ���o'r�n�is�,����3O'�)��y���C2�3�� �~�6Ⱥ�09�-瑴�vng������x���>>�w�����{���O���������uon�o�V���U�Ԋ]T�1j�mؤn�N�.,rĮnR�b��6����qU��{ï&�e=�f�S����)�K�L�Jh Ђ���Ȼ��eb8M����e��l��{Y,�c;D�I=��[Y���p$�,�'����^�d:�U\�F�jL�,�����*6xK<�G�i��;�̓�yV�2�꬗ �w]�}�d�M�x�D��E�m�q󔌘r��s����:�A���/2�j4o�h���c"�J�z�(<9�jE��hD��
g�*mX�x6a�I˾��( �[��ѡt�mb��^tw��Z�ݮ]/l֧]}�%q��1��(۱$S{��.�S|�o-8&C��R�׻���9ҋՓ��c婩�8�Χ�f:��<S��0|m3�)��Ҋ��;���[ �t�EY������ڪkŦ�b%�LB��=]]��9��H�S�郱�T�Xٔ�P�E�n���u-�Ǚ�-ӉL�,հ���E���K0��m��
K�`�Kl%�t�r۬�9��_�*����� (�Xu�ޚ�Y(��8��8�n���foB�9����774�9��@�7%����j|���-i�EA�%��#�!.�/g.�H]�lZ�|Y�oY�W �fg��_#)払J����;��(v��ǰJ��fw��1�=����/(�Xch��SZ�;�]��,�BŦ\�k�,`4�Hn�U�V
uѝAv6imz=��Y�GU��"��qT��AB�&~�؉h�?wz����dJ�0�e��9õ�������¨�r����gw7�3��n�2��RP������V:�	�{�;�ס�x��Ə�R���U����C�.cT��a��m���o��y!��� ���������ݚ7M�Q�f;J��/��p����yWU��kf>�c���_*Ei��8�uf3�/;��iPm27Eu��=W0���̗����je�R#�a+�esX	t�wh/�*p��ep�,qx:��}4�"֚3M2�"��J��k���cB�ט��❘���o�]���BX��u��a�sn%��n$��["������V��yհ���Z����sV��L�ܞ �ާ�c��b�\Ǐ��pN��TH9�f�b&���Y�IObPˊ�<#�o;��2����u��W;}d�����9��T��Ü��� s��NCwD�D.�\�W`ʼR�:�a�;kc�؟�-L�W�ٱ*���֡�M�(󪿵�#��b���q���W���(�ST�;�v�ܩ �n�k���eZEt�j\��Fv�fv[lø��^��1�"�٧˦����{��m��Wb�ղ�ͭ�t��7�p�,��9���R���Y��<�Or��˸��qp,q�R�1�הԬ���ۙ:�q�޾�˺���-��k���ﰢ	���c�E4�DRQTEQ4PP��J�{�PP1%�P��P�sh""��KD@V��T$T4��$T�S^��M)�-�CAMQr�L��UP����E�$��)����
��i"i�"
Y�"#Z�����b"�f�H��+Ɍ�-V�ԕT-�PUE�UĚs�AMkHV����SMS�`�hhڰ��MTEHU,U���Ѡ�T�)(����5�QMCD�QAAT�4�@R�KQ	TPV�JLSMSkDQBU�&��m������*���� 

*�65EU�N�
h���������[��xjB�x�U֩���bR�K�	�6���ufr�>�<p��I��� Wlj�H��r��әY��b��H�b�Q�JTh�
A
 JQ�C߿�����w�����/���q��!�c�R򟣌�:�aTrW<����{�IcA�a�2��ja��\6L��)�{yp錀��t��^���n�ě�f�I�d�,(Z��R�g>��=Y�Kg�ew��ڮ��hj��+�Zz|C�sH��1�ͷ�ʅ�
%c���=�]��ja��.4}�m�PS����q��K5�+	t�Ŀ�5񁅟��j�Nn��k��Iv���FF녌w��%Cm?Mk��ӴMKsP=�{�|dD��p�	���#xW�~hcF�{n�^#�����Գ$�����.��2����f]��D[���C��:��kiX%ӆ���y�"P����!�>0��mY��f3"�x��	A(4�F]���e-�>mD��=whQ;i3ԁ89����'�2~��S�VwV�Hyj���J���r�ju�eb��y������d=C���x!0�a�q".��TcW_�*Zچ�!k�P~*�
yY����sL�ƭ�t+oÍp�7�w�dT׳�tS~Nx���ų��<f�E󩦻�����+�%Ӑ��A���q�o!3���O���Ut]O�(�f�I5r�n��o�}���x��Y(�� �X)տ��y�ш�+����9��ԱL���t��wYf+cϺ�c����a���B���1ua�nE���+���ڿ�ﾻ��D�)TiP)A�G����J)
�\�߀(BSe�PX�RxG$Q��~ǫxi����[HN$��2[��'rbaUe���[N$Y�hda�j~"S�	�Q�%%P�ȫ|����{lw���Dܽ�E�-iN�F)�	�C�	�Ay�hO�z{�Rt�$��[�	*L)�Yp�kֹ�Ȑ�"��9�xu���H�f��B`y�\��%P�=�E��*�]ctS.�MΡ!>U:����ڊ�Pؽє���^���_��8Bk�	�/�
6҇C�t�B����{+_7z�ۇY���r������ǵ���>�B�t��==Bvh��I�`[���s��q�k1���m�/I�.���uJ�w?x.��v�^�&7A��4���$q�������T1	�����N������ֶ&�'�s�Q�+��.;���'hs�s�0��4���[p�my����vnr�l�1ǽQLxT��x�}F=��L�5�f4b�;ڱ�
�	�ڜz�8aȍ��0F��y/��v?f�vݾ�_�?���-�����o�Ǘ`5}�n2��2��A��WD�o�c#��;�]*;�dYKs��SM��O�ɇ����1Sò?���4�$׏����3�5q��Tz	}�f��+�,���j�� 4�.[�i:̇֘�Ќ�}*�l9���wm���7�U������7��f�E")�V�
Q\��SC�w��f��f"t$�JvD������x!�y�܆,3C�q1*l��Fk���>�v��gs��V"5��u3�w�׹_�K��+)�F��N�T:ǆr�6�&a����=mt��FƓC�*i��� �S�:	�y��4"�04��B�).��^K��r���j�;�3��~����^�mq�ٮώ��>Opl���K�q�.J����Pe^Y6�� Q�^�����V�dS�{�g9B�.��1��[��Q0"]��ʬ`��v+�܄��FPd�-���Fq��ǯ[ռ�2��ڞ�ن��|���K��\�as�; ��b�nwA8�LK$�R�er�&��瓐�3/i�eQ��j{Γ�:{lw� ��ؒ��B�ot�N&�kH"NN���Jt�<�%:ݐ�zS�yh��4��mB���������m{��yG��������0�5�k�ݲK@��t�r�{�ռ�DRt��E*msb^��#Ͼ{`��r!6И��1I��[3b�J0Y"�������M�����
s�E�u#4�Ey����Ϙ(ֿ�O6�8r/?_�?QzF-6��׹E���CP�B}�6�v��C�EO�y��/��\��Y"�nw��u
�������h�"�+EQl��F�Ӗ�s�:�N*pb.��c	뢣��;�J��7�JL�d�N8�,m��.��^K��s7�v�_� �� � H�B�("
|s�����_^�=R�N>�dK"���2��Z�gW���jF��I��5��&%ݣc�b���(B8q�3N@�0|/>�d�tȞu��"�ѓV�c�Rr��6�j����l�:|��t��k���ҥݛ%�2�����6�/�P���dR��ux�k-{G��~�4Z�;0i��|0���G>�_l	$J��$Q���׽A��%���^��;A��o����I���)�|�b�+	(���0~~2"ac���O"���l��ۚ���Pb��.�5ǽV]�ñm�.�|tW���E���A�4h�,b��.U7]��^iv�� �����V���}(�6�=$�RSl�P�eמ�>�S�<����ɍ)4���ъ�.�o������0���W5s�؜j9	?��Z���Hd�c>��2rS�z�*�Y��eȎ
���o�ʒc1�`~�Y���.z���j��^A=�%�i�9O��	�I����b�}{��^ʋ�ڸ�V"K���v�S���d.z�c��y�-?Pו��<���sʭ��1ޞ5N���AI�w*�,�fg��)��z��]l����ڡLA9gj��{ε �^��Ǣ�����S$Vyţy�4�2m��հ7���w�� �d���!�Wge8�m�4Ӆ�?~�{�����O�T	!B��J&�()�h*x�i*T6��C@gM�y#B��T�<�?���w,�r�G����@F����-é�I�(���xk�܎��z����Ly�:�N�2)��qw���Шt�z�#� �j˹x5rjg)��XUք�ܼ�Y�4����4�c	���"��D��km���o2�� 6VvF�T6Wws�n���ZCH୔>uB` ���1�3�0S���"��敼�6��z\�C���oB��X�΃�Mqwd��^S�	�B���¨�yj��O6T�X��w��,Փ�u�Ѯ4Ӻ����ͅ��c-�M��7�=ήMг`��,�%�k)m9�x�X�s�����<�+��0�݇֡�n5��G��i�����@0��P9��Lܢ�U����B�d�����3�a�V���j�i�EԮ{A/maTs	�M49XK��������1����L�Ddlଁb�.�n�A�5���3��`X�R	O�Z�9C��R�ǜY}/a�ɑ.�������]΋g���-pj�3���2��s��t�v��I�.��]�^�&e�@:"����_���X��M4K�6��b�6M�ٮ�>蒧�y�ˏ;�
�\kZ�y@yn��FrDfh���Q�1�P{��gB	�C�P�>��m�UϠ	}YZaϞ�t��ՀE��]���x�����up����>�8��|��:���5{���{���}�P�U��P�	$JT �	D�=�ן�\됐mP�b�G�Gk�<��P���c#�u�0�{!�H$=� ܌;")�P3�Qש^:\;��P܀��VD�X�@fq�ay���bq1�:����۱�7�Hyk� ��׼\�B��C^h~�^rq�欍Ƕ�t�Ú�L����8zv�)�Ƅg|?fw�/�i�N���u:*c@,��*<���ӌ.a͍tS��}����_4#��&u~&1�������u	U-�@����&JqP��(���ׯcռ4���m!��lE�M��*3V���@zSpܚ�;L�P~BS�	�x��f	��IT.�&��_q�=L�`�V�K���wC��h�D>P�����3��I�y�K$� n�d����]�Z����l�xDZ�p�\�z���c�`��\���D��a�Ȣ��E��'��n����v�n��˛[Pʌr��k�p���3cLp��S7M�M�~;*V��w*�,�܁[���6��.�A(��r��.��A8�u��݁��֟��S�E�yǻm���n��l�D>eب�����m�:8�˸�R� �9�R��wn��ᝠ�1�t�'+v�dEڭL0�p�:���XN�3G��u;a��-�X�{����f晊�vt}q�r��XT��}�z�t�$YzkFTy#��2�k;ӳ7����� �	}� 0!�R�4�B��(o{��7���
hu�A7^���
aY�q�6�����Z�����%F^�Gs����z�D1ip���y�,:<�|�|��,�M��w�*�4���#bz�[%
m��ҹ��A/t��9��c�9���3��{����5��[��Äh�#1�����f�z��V�I����\j1�׳��p��m�"��)�X{�����~�(`��C��>jj��'a���!�d_J/����!�qh�*�҇3��`�n,�9�/t��ClC�sý 円�������|��c�:��aO-Xe��6&�Elu��'�j�x���x����N�T?7�Y�-->C ��{d��=�fV*۵��K.�2t�sdp��!�i�,�`R�iGC�^��O^�x^z�� ���P������xt+wkF䭧���Kо�ơ�E�3u��ʖM�-E��3f��ǫxT:E;���eL
�"��0�L�X2��5�EǤ�
��̬N�{��Mz��ɫ֌�{�gP=�œMA��vl��̓3��&)�.{��
����� a�`�����	�ĲO�D�=|1N�|_�v�E<*���rT�Y)i�]s�)ʁ�8(]t�-Yh�}�s������[8E}�����C�-:�c4���ӹ��tmϯN|HԹ������3wCL:���\z^=�y)Ǳ��ΰ����8�գ�+(0_>�r΀ǴZ����hO�}4t��U}����$�(��Iih �` ���Q��)lŬ~�Fc�P׶t�)�� ��d�D�f���`�v4�$�<����<i�g�Ĳ�]�����JE7W�T���y����?�X1�lj�rNЏ���$~l�Ə�%]o=�j.�\��z�p�j��;�)�I��Ș���}�0�a#�C��B���r�����zSQ{�:�A�M���-?,��5���f�p������'	�ˉ*�*����K4R���#"[y�z曬v��kY�E�ڑ�a��Gs�|w#�%ݻ�$1��TL���N�(�;E��K�1~�v/�X��Lh?8$�������/�s�^���[�frc�����t���wf���A�����wf�E��k�ƅ�D�E�Yk�r�G&,����<��F��R�j����P�zd4.)���9�SZ������v�'u	�ɦf�4�������i�y��D�sQ~�Pw9�C�;V�&9κ���B��Έ����pm�-�"�
�:ztК ��v�2�Zx�wtE��sͼ��m�:�E�l�5^
V/)Q�zn!�gJ����H�m�*��Ơ4A"�.�U_ejS:שd�Q��!���;Yd��j׍R>�pB�I(^��r��n�b
{�j9xR��i�f�퀥�U���c��?k�7rED���ōP޹��>���P�X �Z�K�o ����:��]���ȷ�&'�!`�:�n�t{�̳L�z;ŝ�%6�]��D��C@~�H��~ԕ��3G&nB��t:`���|�����]��kQ�H8�Y���HjHγ�5m��j��9觘HVhE��6/tg/ sӼxX� `��a��W�M�&�TV5{T����	�3j��#��ݤ�c��� [�kJ�ϱaȩ�ԁ9�~b�<�P�s��d����S�����+4v.�訤���B��T�SW���WT\:�q��"z�,���N�ON�[ig]�ݻs��'nc�9��=��N�$hZ���qv#��O�"�t�z� c=<�:�/L!ss�%��J��1��fA�p�4�R��	�\�):D�&:p�;�0�����L�e+P'rwHw�C��B+�G?\�"�o�K*���&
z�r�d]`���1e���ymT��fv�{Kߴ�z���XP�
ρ�mx熄���4(��L(�.yn�r��uئ�H�/w�wb��Щ�;P�9�ݛ���>6�M���&(�Xn��}k�53ƽ�ȼ��$�k��%�$d��eM�_~����w��*#x(�����ꭈ4����7��X������!�e�a,�v�]8�3����	�L�u0�`�P����� A��u��*2������j���s�rc��rlۧ�:E�+z�v�dS��:
ji�O_a�K-E4AA�~�	XS[�r�ҙM��a%���pN�<����y�>���~�� �����;Q"�p�(Ĝp���簔{�����O��&��a.���?�_xk��//�8.�/�u��0dm��fJ��a�GR�l'�{�;N׉�nc�,�^�90!޶�^_9�9�����|�� �DcwV��Ⱥ#�Y�|0�LIv��]�^�3.���%�quQ}#�`Y���N~�(Z_���M?$_��������#בd<׏H$=� ۬6aglJ��zs3��d��U퉷�:��0((E��̔����_��-[����<&9�u֙g�Z1�7#Eq4#���.�W�n]s�>���8{���*��	�"�Yݕ�_h��E���!k߱B�eХc�Q�Czq���C���3�鱬{�j��*��/N������AvKg[��v���Ȅס	�yb�I�Q�g�u�cռ4�{gg�1r�Z���S�q�9����2 ���
�^!��<��Bc��N��M����b2s^�_������y{�^�w�����{�~���������ٖ__r���7Y���nĵ�n�_���Y���;�(�+:�Ϣ㖖�ܴ�o�Z9��,�5�h��;�K��}�1��ղDRڳ�n�U��B5N�l��B�fd�\����}s�|�}��g�����v��±�Ξf}�,�\M��qr�c"43v]H����,c�P��W`{d�
�ǟ ���E+��`l�c���È��"I�E�x��۫�c��%�R�Z�`}�V�m��ݬ��g�(rɩ�ުO�(h�o��1;�����+�4mhk5�b�wW���n�����\�`�H��Y���� y��vj����Һ�F��W5�F92T}�$��P���Mw w��2��ƺ��g������q���r���ox>[��/���ǌ�偲��3
2��x���Ai�����N��BSٳt�pK�t�ļ8�qa�ծ��E`#�=gp�4�͗ֆG�z�����1O1iN��uAǵ�c0��(�M*�PV2�6��q�%�uy����}O����� *
*��|"�W�jnM��[\]���ŝ8��9v��.�wr.�G����n	s��P�K�6��p<}:�� j�8qng���ȣQ�v;���u����Wl�沅d�9.v��f����L�K��sIӂ�.�
h�iAy���9�8�j�s����`͈7��_j����#�
)��7]��%�q����&�5��d�>$�����F:�ۄ��l)��;Y���t)�hC��,HlD�b��hAk��c�3#2�․��yl�R�+-���W��ME%3%;I�hu�z���HP�8�N���B��n���{I�,V�e��n���4���kda�pN��qC��ņX��#LI����e�����vĘf:o7w��Η*䦰ؘ��Rm��t���B��ò���]�b�ϱ3PK���Q�U7�Aj��-��(P*�4��E�mo'Y.�N��T��1�P�Pd��bvDZ�Mmڝ|˭쭁�\6�)>����oR�L/8k�&�3w�N��V��$��GC3R����dU�˜Ì˝�,3EA�6�k �+r+Ck���7.������ss�� ��O-C�o;��'p��}���f*=r4�i4P�mM���̴	(������j^9��\,rظ�
2�v�R>#%m��3B�8��i���l��7jQLR��r��˺�N̺.��=y*P��<���JD3}n���2�w ��7�rj��4�8��bV+ʶ�[��|͕���v�=l�S����qp�=�ucW�a���t�R�9���7]�J��j��so��x�%u�W�}��u�|_T��o�;�ז��,[-����Qâ펙���{EJ�brFB&Ik��Q�����߿F��s��P�ͶѲ��c��%(H�)b)*�6�!�T��V�Hi�J������Zj�i�j$��"�h)֖����$�
)���H�*�MSK�AIJT[f5�m[Mj)Ӥ�u�(�*R���h
J��*�5��f���%����K��"j�"��SA�%4UCT�tP�A12i�QBD&��E&�hd"�
j*����@[h��hi�(h�&�J����֒�������((Ӡ��)����i(������6��L4��LE�Ʃ)bj�x�C�Tr�B�I�E�j
Z�"�"��Z+X��d�������v�j���JJ��-��@�ACTh�U5MSM4�R�QRĔ�Il:�)j�4:h)i��R"�������
�����M�1�Z|��T�EPl'-�}uY8܌�����.�V���T���R���"N�o�9�͛-v�B��J��=;Q����`��XtNa�*���Y�e�N0\P�� Ф��)�&�.(apD�	�PK�~?~�{���.��NL�]��
֖�h��)�s�����rC�8!>z;A�k�;�Ru�c�:����5t�FMk\��o����g�������_�F�U�����sץ�n�!gey�(�`�460�5��C^�=;Fܣ�Pc�Gz���`Ӗ��@}yY�����	�&�eP�F��T�nn�\rZ�8�&L������PX�]&���w:�������kO��kp0m�,n���n��dp�]nPf���(]���זGs����s�q;/No������z�Ŏ�)r�x�8����9�6���Ԛ�X
Uc
'�s�J	{�T�ƪ��-����d\��QW����`Ȋ��b18�Κ�a�q�^��+2�1�'���F}:�	��Z���3\Sk�e��X���m]
;���l~�Ƈ��|����ֿ.��� _J/ş�_FK?'��]�Z�C����EEx��"�6�b�z%�X@��\<(��6�/�	i�B7�m��t���8��� �<�hH�k�[�����sY�M-$d�l��0�v��Y�L�fuX�r�i��LM�]\� ���J���Eo�o�:���
��j���:��r��p.���W&��9ZZ�[o\��yu�F<�V�%8�;�����l=�W�p�8WD������+�����?����f��������6�������ᗦ��BH3xf)�=�T9�n�h�/��5䮂;��AAy/��Zfj�?�>0����U�YJjP�Ȳ�T]G��O��}�3�AT���2�%�Lh(���6����*�y۷�KC�T@ˊ̂7���!p�C�h��<������	F��=�D�>�	UMV��xF-�*�%�u>Ocb�z�C�)E:	��׭���,`�as#U�hq��n��'	�d�\/v��\f���A���E�I���F��W=������c'�<��?�~����X.)�r�L!Xұ�v�l���/��:�N�.�L�$�5��d�P�p�= �5�JY��82�5�Z�՗x��]���S��L�I��Rr�@��msj��:^��y�=����s=-��2�����Κy�����ΨjNuD7��/C�Z~XH%���#4�O@~�.�Z�h��"�$4XPÐap�a�.&6%�=�[�i��N�q�I慩��Q���z�����X�������.����3��X��0��C��ƇU
���Ȧ4���,wJNZ֙6�^q�x��^T꫔6�%�Wv,�����X����}���!��R����P3�w�[�9�Yu�f��"�/�3a�gJ�	���T��&�k�x�Sh�#g.R��΃�����Vvq���H�A����0�I��gT�(�ꮁ]k\)���U}�[�tt��}�*Y�T2-ݘ϶3�L�9���]ٹ־{��hg�D�5xU0�Y�����m�p�E�����Ǫ�ϼ�����鬃��^��GM�w��:}{օ.=�����4���aW��.��i�-�����1�P*�A�ɔ�������2�W�g��:˜Zr^��S�LǷd6�Æ��]�Oh�^����(�Vr���{Z.J��iV�Ʈ�W��X��xu��'�m�ݾ�n�h�gK�%6�5�˴��Zy���1��'DS=^hQ;i㐹����M��x*�����'�Of�M�a ���,����!�B�O2v_&T(}��L�#�V���e�)���x�0BO^��Ƕ蜐M����j��>��ժr����G;F����2&��{�J��ذ�S��V�+����y��;H�:ɚk�-���Tr�͊�z�w:
!Z�E'V��U&��8���7��D�;��&Y�u�:g��^qse�[N.�T�p��-�^�Y'�b%:HȤUQN.�ۼ�"�{�����}�.^8y]64����s����EhKrq\����2��w�7 �	�kV.�n]4�,yM��}��8�iY�x�5���J�9���X�� �:m��M�4�ph��=���G/�Jڷ���tJ#�l�曭���S�f,�?�_U.�S��7��ׁ÷�e��ntC`�u*L���s@���4�����O�lI���+����0��{�#G�vC_�`�"����P�;*Jz�Sl��`s]���ѫ$,ģ���=o{aGf��;�r�ځ����z򟣻ƅF�v�
����.��Ah�A���n*�duJ8�JeH�C�����n���[Y�&y7��ubMг�]�j�U;���i�G=p1rU�+ֺy�Sa]k	��Z�Z	�<���!��Ly�?�n~m�X�u(��B���P�~1+u��+��PK�Z��hF�s�w��p�35�	�����6�'j��7�6��mgRa�GR�l'�{��v��nc�/�@�W�3���3�ҞǪ���p�wDd�� <G[��T���t�t�9E�]���v�f]��upK[��W����ü&3���,�S�Q'������)�ۜds���^E���= ��M����k�Yl���/�E�\�]��v{�m�xll�O��.2}��Ƕ��zz��{�A�)��R�� ��V��ӎ~��/=����+muu��~�J(2FZ��d��ɂ*/^U:�m���ME�QC\��&�\�8�h�5R��N�f1�qƤA�nn��zY��ϕ�;���(aɛA�śK�Fǐ��&�m���tq�V��� .8j����}x��?
z�p��Yc3�NV��P��=7���9\�(r5曌�]�������x��C����W��$���k;>s�ӵ��SvA���2Ҥ.{΄;���B��J�8zޜa71Lu���[�`���pأ���'��G;^F2=;R��:��a(cB�ܣ�,�f>�z������\�i�e�Y�2e�E���|�LGd���Q���&���)�P�&"T-����hg9ߛ�K�:�0�O���9�ªf$�Wڽண<�և6���vOy{ıb�-���+g�ѻw�4��j��"�\��~U�զ"r�o��Tr�_	�vQ����"}��d�+'^�I}`��Jca�%�͘e�9j��8zh(fƑ!7T�Mˮ��������֊$Wl!exr�*�qWK�o='�)��.��IĻ�;�|�=����k:�
���W���}���[h��'J�7�3m�����w�s��=��^���=ydi/N�]�-"j%��0�ۅD���i|�[��(����޿OQke~Jq��ҵ�`��{
��2u���߿i~�|��9�f�n��:��l��䞓X�e/�6e����X��L�Kr&��kNT�%}/2�xq�=\�����4:4aG��y2���\�b�	Î�hZwI֬V7�M���L*����נU���
WO8�<��wگ� >��7������S��򁣫�dd�*��eR���:�l#>�r�5���6�{�ڡ��8GQ,�d�w=v8g�h�^a�_��:~���"�Q~�M�����^U'*�ۅ��c�3��8�zN��-]b�<;�Xhl.Q}ڌ�Kk"�"1��u�˫3: ��A�,��$=�c�}��#<�Z�n���L~��2t66s&�'U��T�o|t�n��t'"�����;�i�*�KI](w��4W�b���*JO�%t��U�걜��E����i���sR=<�/fq��T��aEd��
;A�b��Q��޵�<햣���CpF))�����\�"���g%ӱ^�"^�eM^�f��c�9��U���r���y���V����?�1�`p���x-����[�!�.S��i���[G��I��E�]����5�F��W=����{�`d�D�f�	��v4��󮄲U�ѳ���.�^u��xN�]"�RJ�Y��d�K�����c̛0?ߡ:�C���_o�.p���l�y��X5<������Vrnr�0�i"+��5�jպ�GL��pn�&�8HU�`��A���2�<c)����S��5�3M�NJ �ҵS$ҬR��)KZ��6���Liǌƻ��7�6A�wg�L2N��x���'M�����f=��7�d�RO�I���"���9�����kz;Z1�����d�C���*����@༞�P�2���z.@�Sq�t��Qi�c)�o �u#4�Mt_k�����N�r&�~L!0�s��t9���ˮxz�
n��Z�vy�T5�=%�LUi�C^�q�g�j뫺�������x������� C�~5�ήL�c@ɫk��I��Gh���s�kv��[�H+�GUI9Z�"vk#�O�x��/~H�9o�C�\�g��
���a�m��Zƣ�Մ�+��2�����3�A~���uv��`����Bb�!������jJ������$��ONR=B4��i��
��;k�uƾ��Ƈ����O��%�f��֖UN��}��j�B&
|ٿH��I���7	�f��v-���tE��y����CݮylwO�Ѽ(	� ��"a6'�Ս��=�2�3E�K�%6�7#тN9��J//�ϝt�:�����sͼu{�S���a���e�j==�6��l$W����0���f��:�U�(X��$��U�Ji])�o�z�����vT����S�t"��L�i�^5b��퍝��%4j�X���"�=���.�F>�R@�/�3#(nD���ܠ����C��Z]�h96���/N��0>�g�0%�U1�퉯�Uzg��]ߦ�����g��3��zw�����5����˃޿��a�n��Ù2�R=�x�tDg-���,�,�3
�>ņ��vר[�������9�N9�V�a������v��}@X�6<?3s!
=����_���J���'����z��D��N����n:�\>^��;�r�Jas����8��%���2O��Jt��H�U�ߢ�u�4&f'�)]wk3F��T{�z����F�âL:v�����s�{�Rb��!�6֞��8;b6��:�����巰vp����[�����0�'�pG>x_@�U�j}�RS��d]>[��W�yQa\�j��C���LI}�3�ˇ��-y�7s�B~�<hQ���³E��ʚ�#u]��^y����RX���L��$Mv6��/ǧ͏Ǽ�)��l�Y��x<-�=2�����(��8�*K-t�)�u�$�}njp���g�}=Zx��<Q��},߶��}����*i^ڐ���4-'�n;�~��S���b�0��:�9�;�8a~q�}._j�u!��c���R�R��(�]]u����o>)�S�x��v1y��<.ͻŵ�6�]oCO��&_��՜wk����kM�!�%��*��5
m򮦥%�/���Pt���,�ݼ�J�wYt�r�T��MV&��kd�cbUiZ����j�7y��/��=�c�����]���t�/��w$Oa��]�%\c8lO��,ݹҘsp:�a?Mk��Ӥ�76��0�=X����B�b��f�g�
��T'�OC�C�7���ʌ�:��f�Q`K�v�q�n���<�Q�S�p�w�%��G�*9�kW-/~n���$��/��ӳ��;����D}=�H��xk~O�9 ����H)չ=�v@��e@tM�1��̀�4��Ĉݔ��Ƕl�f�fqo���M�E>�<T�t$Z��O�\�+܍y��-�WL\:�:)�;D�V��F4��Z誛����GEjϦ���U,h@�|���0��,���Q�o3��8�.b���gu6 ��=�y�I'%�B��@`�֘q�|�q�\�Kwy�Ȅר�L�V�V-<I���u�s�ن;x..��j8�r���
-��J|������#�O5t!)���)�P�&����yʱ�pk)mOeGb�2f P�����xO���C�h.�|�'��iP�5��):WH�ǏtJ|����d'W1�)�SqJ~#�;�(+��*���9��ʆ�O������c���6B��O{*�6��XX���ׂ���o�7Y/`[+Pؓ��m.l�J�͚���	�<��R9|��jsp�tu�n�@���GP�*��2�̝��V�BlQ����j��u��\�N��Ą����́�>�!�]��^���ó{9���ݙ/���:�Rr��5(��7E2��P�F9jw�����!0���;fЅg�j܏*nN��..Ϊ�z���ʂƼ�=&_���K��|��q[�M�j��Ս=�[��"�ϡ�r��.nL��Mȭ%Q�����+���@�^�=����.�7pƳ����V �"�d����Cji�X����X�\���w�q��~���3�.�������M��d-�jC�<y��ͮ�!ٶ޳��L��I��4z�ݐ��F�����gU�OA��.��֮>;L��`ge*1	��t]�5�Nç��l�m��U� ��E�"��iۢ"r�.�%����I4ԔW��W�K�jb���.�����xQe�֢�&Yp�sS9Y����I��c����4���� LYŜ��&]��o�P�X�����K��=W�c��o�Z��e}������C�"�'b/"�7s����T�/��4�W�Iwy�9����m���~�]{��z��̀*gZ ����Ag��u���O=^��Q䩛���Y6����w����������/o�����{���w���{}===*���dE,��0յ	 �z%H0�Fn�����ev��l�����r�����R}zn�=w�X�Q�֞�.��
� ����ӫ�gɚ,T<K*ֆ�ic)itu��U�R�[IgY��B���֨��Y�ڷ�{-M���쮬�<Ʈ��K�z�ϒ�=��ժ�{��i�ѧN�h�j�|m��)�S�c���o-��zpd�r�z#{܎(HB�X�{�4�6�ۇ�)$iQ��s,[ �7� ۺ�l��R�w�Zi�h��a����sn1PZ��vvŌF�
�Mb\�d�j1�+�ٽR���l7�)鵈S��V�!4[K��M�hIC7�43=�6"�X:�t��$l�����Y��|���wa� EK�g}���#|��������.�ʘ.�P�%űj{�h[ǵ+��P��5�l�]q��o��\\������l�cQ`x3P.�����\#m�h윛�y�;S��6�!���o?3��'���4ls6����
�R�f�7~������P����x��t�&ھ/�c��$��7��̂�w+9��Ϯ�8ҵZCU��Һ9�IG��g9Je�<,vk�Wll��̒ƍ�xG�_n �y���D�.;ϒ�o9GC����/%"s]%���A�=EN8���Ң���z���p�[	��9�\�vs��N�����@�Y7Zt��(
��NmԦ`D�ј��op!5�8s9����wT]g��aq�� ��v��r���"�6��Ӳ��}�i����� �����Xuf�#	�kD�Ȇ�QAJ���o���9<�
�"@^���h���ś+�Y��2t�ݎ�.cP�}�u�(�췝�I�3V�پu��	�	洘d�n��$4��Ѻ�Ȁ��< �f4�kM�S����X��o�Q\!(���}}]W�£e�������/��a^p��5�Iʺ�����ױю�2jZ�� �h�c��ɢ����"��$:w �TL*|�X<�٫,���q�ڛ#v��F���ϴk��D��7N�Hj
)���ꁨؤ�,%d=3�Z��S���=-�ig �h��o:�R�u�Jȴ-����v�1Y%e!\�إ��˴�.q��������Sr�+*K��Ld9ڝ,���1Ĭت����Kz~ڶ��]�����K��='�S���5��]bQ.N8��ip��:Sme���+Y̭h�LVʹ`�*�}�]h��>�[F��mC]�7y/�N٢����9�2x.��fV�����I�h�pr�j�,���ZLA�eYc)��o�b�c;�ݻ;N�k�u���NQ���5��J��\�A�Q����%c��b�N�W'/y��)XVM	X�gf����r>��bU�QA;7s��M�&%����d⁠%�Y���
6�wǙn#ֺjf�=}5,ܮy.n����wGswE!�٠���1�쑝UC3������Jb�M�b]��th���P�4�RU:ZP���CK4TTE4�%��D�LU%35E%A�AN�!Mh5EP�$Q;gA�"h+N��
i5�I��Z
bh*�h�Z��)-�-N�V��8��!�JB��-Z��)�Mh�(
�)E5cb�����ca5lQ�h4b�(%��B��ɶ�i���V�6��`��)�h*�b)�h*������T�CĚty��5��9:j"��d�����4U�'DMrJ֓D�A��)J��(�!��Hh��4;b���Dl���U�f��[&����Ӎ�e�1� ����uE%bt�@'��.~O���Ϥ2�+c��r�ڲ�9�lب�7)�^�/V<�%M��黜	3���3T�ޭ���{ܱrTc�:=��<��/��C���~56��=�ŴS�\zz���	_�b�=�Jl�eLf�h�O:�/�m��e�v���'�a�s�Ve'�`��?��d��Cέ�EF*�T¬��FEY��Q���ga���G8@��E�%4���ވ�8��&��<'�%�¿d}���	��;wa|�p���s�'�9�N�ˤS*�J�[8q�������kf�}M�njY2���d^�0]�a�wP�|1���)?��c�sP&0����&0pyv5�FS���-S"�z������{<Ԟ�:�E�mOC�Z~Y�R	}E�ul�oG]�g�~���{��B?U�_<��=�5��H��e�`O\�u��ֻ;^�^�b���Sjq�2c���U��V��~�{�D&��>�,k~�@B�P4.�H'/��2)��4�.�̐ƛQ�޷y�y�FU�XW>�U,ٯN�ۚ}.�7���uCs�˅E5w�]��ڻ���Q�,x�k-{G���j���a}Ph��h\S��ψ�����ʸ��a�9-�08
5�/�|t���W�n��?�n�f{�=F�Z�/j���5���M��IЄ�a-Qw��<*��u���)f��"��R\U��1��}9+C��j
$7��r޺�{�d�p���Rз�$�oDSf^]n��^"���\��=�`��)8%9�aC�@�b���r�z0C�gg����p�o9��j�\�=L�FAi/�*���+6C둇	�L�v�q�b������,�^�2��sx�����a3е�M�D��`�<.H���X��m�8;���f���I.Ԕ� �����8����c��g�NȽ������K�
�B1��~�N1����Wf�2�H!z��7��Sa�^�T�=��=���@s����g͋e� [:y稈q`���	<�|Ǧr	ݔ��eЇ�ܴ_h���,��A?5� ��@�T��g/��xtm�k�}l�~b����W��8�n{Qo����Ǥzy�~�x�y���eo��'V�P�
S	e��/P���꞊���w�콅y;�Kyx(2͔&	v܇n+��淘L��xN��R�)�؎�as�|�'r��0Uv�v�n!�CD����$lcH�DL�2�m˷�Θi��&@�M�?��R~�)�ׯz�r���S�f!�qx��-ᄍ������`�>��,��h�)�|��k�j�F#*K��lN��D^H�zwyf_��Eq��==�>���F��Ȍk�R��m,��R�1LZ~
�n�W� ��/'-b����{�et�'	yj��є^�"��R�Υ��[��V�m���ʛ��lG�������)*p�ԻԎ+3Bi�����}�zI2��/.Q��6K]�R�׊����(	�o<����~�<s��>5��s�>��z�OHO�3��|�z�c�!�V���I���O6T�(�7�i��k�g�/ǣc��-}��nJlSN�j���sDC8��zUкL�N8�%QaB�O2�S��ܾ�{p���I��$	�q����4df�f�u���t&��G��VJ�e�W=�T�֪9���'Z�=�x�W����T���C`��g2H��P�6��mgQa�GR�l�5�|��v�	�ne!������Ŋ�B5׹�3��c�����!0���~��0��Ӈ(��bK�ݦ}�g(�\�`�t�k�EL�n��\������kށ/�0�!�>0�F��#�,�Gf��]n��B2�k���%�a��\�Oss������	;�f����C��·1�0�p�\��Z}y���_A�%r��ךG�2�5t�îyg����Ɩ��]�S�%����ƭ����Ԡ-~�2�]
V�����	��P�<�Ϙ�,W�k���m�|��;��������r��6����\g;3
��$�8�Y#���Ev-�:}0f�g*� �:=Tq�o5� ��`E�V�2��ݴ�1�m�[��x��哨�+U;��f,��EewE@ղ�:.��fc�.�}�x��CD�iG;O��2Q�ͳ�E&�`&J̉.��|dt$��ǃ�MV��"(ĺ	��i흠��iN$�P�		젼�5�<�:���^%:U�7��~\-O��o�t��dL���0��$8�,�|�0O���3��[^�;=��*�˽����2�d�g���W�T�U�`Wq�U�H�<����?r��W�ۚc�<�������b�W{�O��7�I��*�]yd�fH9�������B
��gU��>~һp�<�Tؽ5�	�f��eC�㊺^��~n*�pK��h^yA��y�����4��.�1� �;�M>�!2�ٮur@�`Z�;�����F^��:���Adnp�{[��yc@��?��	��N ��w�������U�Qkd�M��OJ素��z����bИ���3�;G ��������d/Ӡ ��`x>�_�1^w�|ފe���$�mWi]�q�y��3m�p�G^�S�׮3<�Xu�1�c;zk�a=��/Vy`Z��>S`�0���/�wخ÷Y�!�-Eـ��-W�p.L��A���;8;����������+�^��p�Q�&�%ieM����8r�,������rm��'=(�j �p��S����bu�{�y��f{a�)j��/�����ٻ�S���������)���zK���Kϰ�b��!��@��b�Caq��%<����j�p�׼}Wν��&�������qhONŴS��"��Ȗss*����f+7��z�2��Z}m��=�k;�sH��L�}����C�}y6�2:�V�Z�W
����k��3+������<��S��^��W�%L�c��dS�Y�(̺e8��ɝ���W�L�zǫx������,9.�������Q�>��%6t��5��%�t�#��s�j���q�����?}ט\.��p��_��(ب\@#[R�~hǾʾ[��v�N�OlQ{��(����=���_�*Mn�j�VW�+I��2�y����-�E8sb�$*����m:��CSH�=�y��$�O�bS��S*IRkg�m��\:����י�zޜK��{tb��6��3C/Fl�*�A���f{$��0�I>x�S�AXt�U���9�����󚋾�|��m]��"��Cy8�#�-��p^�5'����M��r�O�)��/�-Z�]�vf�jg٭���U�E��,%�o}�{;1����h`m]��"i��Y(ɚ�{�+ :�t98s��ɚW{7:P���a07x>a���/��.�f��'w-�G��]�s��{�e�l���G���m�=�p�eۏ[}:�ၩ�2;�'�,���{`��[@�!� �˞�i��UkY�E�iۛ4[�5����nE{̛e�#��_�I�wm|gaHl����ٓ��U
�W&E1�wiNe�Q��̥��S6���nXЍ�NZ�s�OoV�|�U	��i�Yx.!�<y"u~��*� ���,���;��{�����]����������W4�����!ۧ��a��-�mƷ�a��^��3�ۘ��t��dGw��N���0�- ��@�r��`��&�׃���\��tg�}��E���;��j>�aj|=�G����!�y�Uq�B*�e �$Ђٚ-���*:� 3�U��^u�}�`��h�q�>0�B����s����e�b���G/tn�ߌ��+5���Mt�����֍�5��ܥ����I<bO��4�?���������)�T��/�'�~ ��4m.���-A+��3��3gc�gO��������y��L7Kwps�Y҉�zCvj�*�Ơ4�	�� ��&Q�H޳ь�Ƭ��sW��P,�Ǘ+XoU�Da�̽��.�-��#�b0)�a��Sśq���+��G�m�cBt//@��Z�J�%���
+=p�fȮl-���bǝ���,W8+J^�'�>�n쭹Â�Rem(f�� �3s
.��c��uM&K|4�+�D��	Y&g�WˎͫC�"�V�u҅��S�}����o^���*����Z�B��T�SRܜn��uMV�'��<e!�gk�QgC�&�{c���as���v�#�SsP��&I��"S���Jg��|�e�+�m|��ٜ��&Qmc�!@���@�.C)�l nt�H�j� \&GYVofM+T��޹�h͞ҁ�C��qӅ�;�0��@����Bs�y��,h�P��Ǻ�I�W��렝zIM�N�09��o(6��W"x�XV?j�ׁ�U��TԆg>��Z�W�u�e�
ބ0�a(��-V�Ry*R��O�ݎ����X:n[1���˲��ݦ"�j�Bv)9�O]VI�J�Ʊ����|d:83GE
1�_����O�h��G�>kjd=Ac���8д����]���Q�Ѝf�QD�I��f��s��Y�����
�>+��C��r�𹡵,�hgQa�u)��{�Ӵ�-�$��YJ�*����9[Ad��@�gނ%�A���~#B��쌟ܑ���;�X?�zՖ�Mn!�bu(M��<����ȩ�g���÷Ts$�c����g�����ZZ��u���[E���VQo3����+C���������iKy����slE}&�+kEs���c���ma)R����;���1�]@��&���@ۘ@�����2co�����v�&]�^��e�A�ƀ���KK����P������oåa�tF�9����/8�A/5�A!�(4�@*v�-m�:&��k�`L�\9���<l�������xF��^��Om���o�<����W!
�y��6��u^�y$>dT��%��A�"�z�渑�ʹy�ƞ�2�Zڽ�H\�]D,��*<����v�9��g�m��gPD���!輳�r��`��q�v1���mmr!5�#!2���'�:�Jp�'�?U�>�C��%Ggu���ᩭ��n���%�$/ò�CH�S�C�	LMK%ǖ�ȋ3=9�Y��l�_PJK�!B�"������y-�'H>T�!<���m�����eM�^eN��͝�b/�Pe�:��ʼ����0�l��|�� �6LB`��RY3>wA��m�#�ƃi�+nzvEL/�J.��)�-��0i�Pw����F�ʽOz-5��Y�rf�B,AeS�H� P�~;JU��^��~���4I���]��=u���q*&��F�f�����W������$F;���]	n�:���У*�9
	��av�N0��|Oc���Yi��3��j仂Ĺ��Wc�.}&�^سI�*$^���X�%��I�M}���zi�J-�v�i��Mu�s�S���K�7����H�#��`�g���==Bl���&n�൙9B���еΦ���rWC�(G�E5���֥[G���^ק g@q ��
C�@p�_�@�m[=Ey�B�`N��ٽ��ѷ8Z�OJ0�G.մ�~���N����t����(*���eﬃ��_އ�����KciI�5Y���O��я���W�d��ؗ�w7�DOV�!�_�MP��93�8]�u�ONW)��~��Iz�@�%����-���þ����Q�A`�c�x��J��H+�l��w��b&������$=qhON�_E��b*��&&O/Ymo�pn0Ά--#�gknO�z/�t�k�2�&�KA .��K�w�Oƙ��c�*�����N\]�lj�0,=0�?�<yK�T�>n{؊l��[5X�(2跮XJs��!&�����f�OzzFyT� @[E�E��q�� NW�%ª+�Zq�.z����6������*Pb�-��(�0<�o��o���� �f�b ���5�-�p�����T8�j�ǄA ���bMWi�����P�F�X��&_9���ƗDݜ�1�v��J�� &��9����6fi�{x�]�ީ���Fܷ�!���T�U�G�'I�P�-Qa��}�սJ_�V�rj2?�T�>���z���ps�h�A8�LK$�R�e	Jjw�x;��L�mW�X�s�Ѯ��1����Vv���@n4�'ݒy��%:O��Jt����5����<6��?Eì��ړ^��)���N�����lizY���o��,�L8��4��"���n�J��0�n��q0&N���t��6c.�u|��>����&���7��E��i�=Qi�"������4�C�,�������U��h��a'�?yY������[��O��������T �{�It�my�K�JBeEGs�|w^چ�3�E�t����ʯ�\�1��6�6�Y����.H���=V�~�)9kL�z�s�SٯN�ۣa�9� �]�5�S��l�6bΘ�L^��چNs��\�S�^5���z}]`�s���ݣa�l�Jt��:i�Y/��Ã�m>63�k.���k�ʄq�I�>Nf�P��׉��Ꮮ/O,�c�$و�����vT�p����v��Bi���ojF�W���#D�j�.ů� �/w�������{���w�����|G�����x����pb�gc���lE�Yπ��v��[|&V��hRQ(' �S2�竝Ʈ�͈	Z�V��\5�Yr.m�W,0�U�j�W;c��{�$�<���٠J��S+�]��j���@u�D��gƎj���&���X}�"Ӆ�{ztw�d�n-`K˴+��˔W;��;1Ε�!��U��.}��K
=gU\��
�S;7|�k`S�VD�w���R*�� )�*wc�I�6�:����#2�ѣ�:���)HLa]n���8�c�=��3�Nu�Ț�,݌ñb'�g9�
��bzj�{n�w�5���i=�V��\="
���`X8�iuLqQ��Ky,��Dc�o����1>ݩ���'Ա��O�Տ)so��ne�I�7xՂ��s�����Gd�O��ٯv�=8ԣ�+M�w8��T]Eu+�5l�%1y�hJ�ir�J�]M�0��E%K�u;a�<��5*���K�ԼC��7jh8m��q�RI�d�;՜��I��k���mvmYD���x��׎�z,R��аmrc�d� 4H+u)�'xWv ��&��k(�������
�"�nT�ӽ���r�(��A��**Ӯ pj���>��k�A
�;�u7��Pu+ػ6
\�����n���F����dx��.�B ��Z7Zuj9\����%�7XX@�H̫�|�HT�˫���M��a-�������]��ݛ��0� �FW`c���ç���WE���/��C.�9��x>��9��	��U� ̔��O�^wA8���is����SK6�P7�v�9��h����i+K��kc��]�2vs��؝_|�S|�C��k����ȣ��~iF�ر��eYӚq]꣺�b����"�\z�x�ȕ6�����y\��´��3������dN�֮���� ���'44Jw�U˽��ksl�˳Ph7�H�˽�J�� �dk/x�'�f�	�oWK�$�W���z�*TȗF���z���S�2����d�]L{q��9�°���s���x5T�v���z�14kW�ͳ������Ό)�%�鬬bna U��;")�bSFi}��o��%��Ӏ3�7^<F�%K�q��7:�u����1K�n:�Ƥ�68sqT®��h����깑�n����f��ԩ���Ve����789]&+*�u�R�Au3bF�� nV�����&��ȱꥠ�'NG��eV��xɂ��9�eb�J����c�G-�Ađ*�*ѴAj�q���{Ύ���	���G�f�M�d$��J���HqtƳh�	0WF32��n����soI�[)�6�s�3`ִL��T�9��-���]1�
_K�c���]�F�^�^�����.6���h �7(�����c�K�mH馞�{Z���t	�$�����9�({�¶����T.��		��BkAE�[�@��AQ�uA�S!��(�٦�Ū4δ�"�h�Z9��4d�kER�q��O�6��ŌCJS��ѡ��h
��ILAE��c�R�[cH�9����j�UlV#k��4TZlVR�ӎd����К"��)���0�b(��M�$Z�EPl��Z�SlIK�ܲ\��<�@D�%:��\AB���d��F�����G#��4�i4�6F"�h9r9Prt����K�9&��)Nb�a`����Ӥ
��$2���]d�T,"�k�Ae�c��^Q4�O�2`����b��@z��2�z3�
��Qι�ndg���H���s�Zy��BovKY%b��0o<ۃ�hh�hD�0�����DB2�`�шnD�h!b"%@[E���鷫�g�x=�&ЪVN;�ؐ�
�-R��l&��/E�3������<;k��t�2�	bwj�x艮{U+��O%�L[pl�.�o�i���o��)�0!��4�21�{W>�H[,��s9��z��KWc�3 �!ŗ!��������f�2��l��sӼz����t����3�Y�����z���/D�9/6٪O�`a��q�#Z�_���ٕh\f�q��b�ד�����:sl�����i��L��FB��2ǲb��Z�R�T�SW���m��[���k����2�ѣ�����΄�M��]L$�;���{%73s�I��Ju~HеU3)"Zz��eM��3��\6�w"�{���;$;�*�1���)�K[�Tغe����V�[
�y�ؾ'(���O4{r ��>�!?P�sȾ�,���"������ɎA����or�ET�x߃ۄf�@��ෞF�=5�Aߙ���� �k����_o�)�z!^�ڶ���T(���zR疼W)<�Ic^GjOɤK��5� ����~�i,�v�5�
��^�z�ꚣǕ����٫Nt�ٴb���X~�U`�;
���&u�Y������V�n�t���Ϭ�Up"�]��;ofG{�p��CMDd��ca�ے,i��닟m��,��*VꇧD^�j8��3������3߀z���$4�i��s��Qsrn���1'Y*Kk��M��a ���sS�̌�X)n=r��j�]�J��f��bBc^�ʹ3�KZ���_���r���>U���Rإ[�.�[�/t81�@�?aӁ-��?�B|`����Գ-��E�5�P7��5�}�t!��3�r&&���C�;\��[����Xg:�w�A��0��o�0̓��,�}�'7C��,�F�v���l*'#�;��kG�"3��W�ŕ�5D���3�0��'�E�E�o�F�&U��q����T�#בe��C���C��>����r�>��`����X�[q�L��6��6l��'�(��^���؀5��
-|����B��ךEϧ-�X錇Dʈ�'���ժ��ɼ�7�b�u����8���O2���3��4����c^Yt)X	Q�c��2����W�
�C���X}3��g!�cX�0��?;-�d�NԷ79��#!2���[Z�
��K�ՠuԝ�c�w^��V��Ol�A{k	ė�p���^!��O2��o⚸�_���f������ �=�5dc1��P�0ܤq��ޭ97�V�تf���{���Ã�����Ч�J��N���ޮT�{Y�R�e���i��͚�5K?�}��^����9n���okw�:T��v�]�"�E�N��޹'���<��S��PZx�g���Ş��2X&��q���5�վ;ć���ʘ'l�en�2w�]r�6N;n�|�pC��H�2��^'I�)��&���=��z_g�!��l-#�S�W)��Xe�V0�u.���*�(��cz(�a�aC^[�[��r��mz���7)Bo_93�,��fM>��[��c�v�iC�Ux⮗�Z�O�`�.��B󵦮8�{�����i8��������� ��N�L��M�"����~�S8�ׄ$���e���._��{�8v]~��n@p���ã�k��Kj�=E���U�/�>�:�6X�l����/�ܞܗ��K��o�������.���|9����h��g�;���ߞ��n�=�~�'�ᛸy�2h�����`#>�z��Q�b^�;3�03�:%�eL;�JΥY��/��_���t'�����>��_��zK���;h�D[��ptK��8���K=R���`����D�����VA���0��>�!����.�|v���W�����O�ԻhF�0H�Y��x������>,R�;FMh���Z\Vl��n	m��\Wv�]-^7!�5���Z%����*��^,l)�o:;�]"j�3��SM�6�b�h>��h��z��b�'a�S��Ì�Mݷ_�2f��.gc>�~����9hj#!4�{d�9��l�n�i�j�KA+�-*��{�۱����s3��p��O���5�<,Aii!Bi���75>�z��Ơ�*f��
SGFc@13�9�Y����cs!�m�ٟ�b�O�t�������8�X�}~UX�*��$���_&Ƴ7�o�V��p��^�D�0CBњOr��
=�Bޭ?*�'��������O�6D�wt1�Zv���j�d)-��N(��E���X��5ߢ7�=����x�O��i��F`���h�) �K�l=;A��<����>1)Յ�)�J<�f�Y�\�?�\�>�\'��?�$C�"���-E{Y8փ��H�����)?�NV7H��S�n��i��V�Q�yŬ-�df�c��=0�>b[����u^�5��a�q�Le�C;r̶�ػ85���~���nf��Lg��5�Ԍ�	���{`m��i�s�׆Pd9���c��Bq�~'��y���Jj�Tև�JO4-o�3(t���>;�/�@lc;l����a�q�@�!��>��;��K\Z�:�EGE���������N�ev��s�;��6$X�	l{���w]bS�4�/1��!�m-\쇯�R�t�p��(��49IeA�������A�c��GoK��nZt�e��w��_:�����b�kr�CDOI��)��J�k��)8�]<������4�@̪&�������?W�FvަjiЇnu�C�m�Bը�è�e�a�U/:��}���mv�Z�ګ�l�Ӆ�Z���&�p�3�1O�j>׳�?������1�a���&+�pʦk�I��ŝJ�}e�a�c;<�!3���?\�L�����8hW��.ݷRw�~灛j�̿Jv�EF;��ߕVW��"�52�[�>q�^Q^��K6'=��[f���w:�D�������Eڒ��H�e�A|kO��sd3?�!�縶E�nndGy)�kk�l�-z�����7��Cs%PChH�i��e]���ӼX0:6�	�ERu�4i�"]Cս0�"f����+Z��O�σTHO^YYPHֳ��q����*Vپ��c�����.f��vd!��4<���t�&��q+��eo��d�H�Ҩ��)��p2$J-Ъ{{��k����R�^��=���ޥY��v��#��Jnj��&E��"S��]�5-pk��25Y=��i�v���u}&\�Oiݠ�ZK;���bp}�+Xɰ�Yg�'�FV���S&MЧV�����U��#���AV�*0��-D����z��#6N�;�q�a u����+5gP��� "����c�YQ��`)�N�/�7Sݏy��r-��1����A��^�2��.�4��#f�n��1�,.+k2�g��\ܼ�d��J}H���N�o$�"1�C���}��l"2�=]+K�*G`�1V�CO�*R�E�1l��m�HMAu:��#6^������C��A�_l� �kN�j����f��nB�Х}��U���T$�⠱\fjxwf��|~����t�g��G:�X@�����z��Rurg����8��Ī,(]<�o��XI{��)����9����~[��g�\<0`�Ö>dp��Vԍ>u�H����=_�PK�l4Z`\�W�c��-�������H�p�38#c�D���+׵�QԨl��;��"���{V��9�ۤ� ;�R���0� ^�90�p0C��o�2��'n���=$e�`���ko�Lĝ�`��$�q�n�& �-��l��s�� \hl/��X充Uۦ�.�9��샮�V.���7u�%�c~�jJ�!���i8"�u�� 3 ���}�h_V+X�^���B�,nnl��i;���U�7[{/�Q,� �����1�f!έ�<%����2���n�Z��3�1�ϯ��+����)�u�S�;c.��ˣƺ�m{ҥt��)c��X�ل�W'|�N�:�G�v��kOo��7�IC�����昸�z�x��7cZ@��C�W������B��H��tј��2k����<C���`�a���b�k��Uz��K[jP{[�A�ʐ�	y�[-WW�Пj���xy�����d�-���~Q�~1��!l�%bw�t¸�M�-��.���h�pt��v�C[���bI�z3�i�S�; ^��q0��DD�j��)ו3�w6E!z�[��0O���6U^�(��<��DcDf�[�Ag��[�a";4�m6�wE�
P�[���}>k�R7 g��m�U��'�P�|֚��}�:���h��3�u�͍�e#�t_c���)�r!7 �?�h2�:vozQ��mli���D�'���;.�3����k���)Lim����~��>�v���]�Q�
�\R�!\�Y�ś�W[�vm-@��t7����lΪң�ܩ��ܮxֻ�*i��&��=�t%��t�;E�?.�}�U�˦3�f2`]c��#�짨|�s��b[X6���:s�4�q��:�c�A�p��B:�m.�*L���;x���zv���1Z�%C�#������1�&�J��8>���PYS���.�Q54��L��2���|�qXb8�a��F+�y5v����'��t���|9G��x�����c�y��9�baʇ��i�[��2�zo�f�r����d^�پG��L�6�s��}#�2*Z�jY~|�|��c��؎�v��Y���H(����Fَ�$O04�f]8ٸ��@�SX��x;��t��O�6�"��{)Tu�m�n��"'ݼNwBX�S_���9���1A{N4U��˫�K=��'�U#U�6爟��衘b��ǻ���)�L��	���֜�W,�l�u����ؘ�vyNa���7t�0���QAH���v�i��`TŅ*:%��i����s�	Ѫ�.7u[����T	�h�*�#2]Ϋt���|q���)sw�lq�T�]>�nغ@mH�t@�H����zی��G]
���q�)n�&#t��)��+0<���AV�]��6�����K���Kտ3�C0�u�P��(�1����ɐ��Q&^\v�qoQz��Z
��ێË'��yI��k����Eݻy����7U��,&J1�Y�7�vI��p���'l+��#����ϝ�b���q��$?������I_:�':��"�q�'h�AȌ�8�$<v�Ӊg|ُh!y�\]Ck\��y��z*2r���6��;(%I��l��]����Z�o>Bݘ�I�M�l�oD`����zdu��)(��t�v<~����Cw˯�:����=��ވ���x�p�̓^����(7T;��Kt�x҃T3e�g��������{���m��ˏ8D�OdޚU�J4ڳB=�@��mǺ���Sd>UmS:�\":`5�'�����	�t_8�qy�ҾL{�Al��+Rj�������w�!�d;��q�;:���I^�tY���x^j5�qv�.��`���O���I�s=S�3�����ڲiԼy�s5y�����HyI	�y��Z�847�`� }_�xW��u�E���,�Oc=��Q���Wb!3p�͇uLvҹ��?�M�j�<���{�"Ss�s��H�����6���W�~kI=7��s��L�a��B�%�Gx%�F���]�&Q�6���������r�F���HԖ�����̃p�ї�9)��Z��i�O�rqW�t���	p�WJ}��O�[r�*M��1{�pl}B��UD����)evyy0RGZO[Md��z���I�Ct�p�y<��q���,�:b��+�&�&1����q#I���2GCf.�[4�4΂��PE�%�n�K5��f:S0.�&V�Ŋ���"6�oj�1Ʃ��:�ّ��$.}(��w��-��yx�L����>�'����yR&[+EK��@��K���,պ�L9�s/�w��&T�{��zy�P��6���wǧ���8a&���=_a�jͳ����R Q\g��*������wO��
������ɠ�w�	��[��dw�6L��2s����ծ�)�L�f�1�uή������7���k��+�&=ڬ�J�u�Փ�����{}��o����{=��o��x��^�W��M9��:��&���+���k��R>��}>l2��ZǸ*�;-���`�G��"��61�)������<�C�Q����ن?�јjn]}+1�V#�<v0�cKot��޹[Өa�湂9�&��j.Ȫ`���ݬ��%d��n>G^»��M�a�L�9���F%c�Dm�]�Nf�OX9԰����3�jq�Ue��Ҹ��R&p 1�ddWilkNv���ض�}o���VJ��"ecb�=Kx̡V-���7�)hN���d3.�WS�§�yȡ�aG1�IVm���N	'28�v��e�k��yV����h\��e���6X
:��F#�����ygos&�Jf̢�%0�����;�e�p\�2���r6�u�V�%_Z"�|�~m���U{.���{�6�G"#&7صn|ܔ�M'4�7�Ɍ*��ް�ͮo7{'	+U�̇�1*"��2�R�m�ޮ5t~v�;vN�n�4��7-�V�"�Ƀ
�h�|�^Sd�� W3�uf�j��.*�����.���@ebI���x���@uC*�a�&]1{&����u�M�/+�GC�+�
������.�o�1q(`�����
.em�'AO^gk���xT.��Iij\�_u}г$��)}���5�0��֩��M+!e*�硩�Qӆ�5��;aw̽�'/1�Z)�W��K:'nd�\�6+N��~��:d��]�*��p�y�n)�
wն#	���u	�F�@�ޱ�T�\�T�U9����!X��:����&t����e��n�s+GoBg[�Ϧ��i�ۑ��j	\2���^�����X�s����G��j�T��K6]L2n��m*þ���$�M5WZ�>-'����<0�w�F�.��0뺳Q����{)֚�n^�%}�#�G�(��+�)ק^`j�_\<����C/&^E�N�Y 1��F��1&J��8�;�U	0� gA��䬟�_D��,&z�kZ �U�)��yn�V�5�9k�z#�_�$i�}�x����r���y+�,�<bR�,i�B��K,�s�q�c���9ŋ���8t&��Ӹ8������;Y�����b�5����3r7Ǫ��H�uN+-���K�H��y�X�;p�{���$̓j����S��hkԑ��ڙ����ހs�@^���ˏpbJi"�#�V�f�ٻVum�i.���3\2ͽ�2��:���Zw8.{Ӕ1�	n�A?����yl[9���EՓ��v�tb�`���Bm��׸��؟f��7�{�L��o������ߓ�j�f
�\Yנ�
)ab�r<r1f4mo=R�Ξ�=cj�9QW��JKlIX�<�n��/^��{.'V\C�ά3q�˱���\�CRϖm��N��A��v��8���f9!�l�RKy9i��&��v'}�:َ�WN:�:�vYi��O������<�T��kU���Ti�\���F�X�j��-��,�t�M�6V٥�O$�hq����:4[�v��ܒ�Zi9��E��T4�M�A&�-��:"u����-ibCl��
�ڨ�ˠ�ض��i*���E�шuKK�+X�*4�+T�S�Ѡ��ڭTQN�K�l�Ƃ�itgM;e��$f��SN�&Ŵ�Z����4���1E4cl��ADi΃k`�kZѥ���mS�4ճ� �Ɯ�Q�i���h6�2Dmd�����G��u�����Y��܇oN��uf-/z�	���w,�sԢ��Xqk�'+\z�`-�����jf9Ω��ɯ[�cc{&\��/{g���߇St{G�sG��a��*���U��c��g6���v9�Y�ǜ�P=>ذ׍�1����#A��ZsL�œx�ݹ.��Z8l���i��L�<[�A1��M9�m@ܲ꧆z1��R�m9W�ߨc��1���/�T�K�>�J�I"}ı�5�y~���h\��i��w<��y�u#ƮO�S��݋�DH�=>F��<��W��=p�tdP�CH�|;��qCa��Й>�B�.}�J���S:��+re�1��qG;#��yjE�9�j��0�$-�bW�&������ۭ�e���R4�J�G$x�܊�s5l���n]���y-YM�4�Ze4y�/�6o8D ���	�D�%%�W�.�m2��S��ՐcWU��W���'{���N8���lDm��IXc	R�2I*���5Ӡ3�#�׶�y�hl�b�3���J0��WS����pT�s���0�y����B����;�$�j�is���ێ�˽�_V��E�Y�q�
yD�޽K�#��r-Ƭ��H��P��4�xm�ifzp�q�tKj��"��/v R~]�A�+����<��U���J���}m�;vj�����$F��Mq��Cy܃���ozMO �ؑ�������o�Eݽe>"��5�m�ܦ<u����cp����=݊�Ԙ�`����5F�̓�Kk�wAIy�&�a�؆���oN��|n-��RQu{���=J����)s~
�`^J}Ѿc,ã�q`l�f^L�2�/`�v]g_\^���Y�@gPQ�#�W�)��1�=��_r�����*�G�q{� � ��͙�c���|�w��Ϸ�r}��+���������n�3����)@�� �l׶q*��bGq#���{~ޔcm�O?zRr�N�S"�<�^C8A��WC�I��N��tD3�3���ی��f3�\��ňz$q-���������5R5螞w��,V��}���$'��}�3v%�a��m��ɽ���������'�_��H�<��m"�̗��:�V!�����J��mcV��`N_h���������:�g;'�����jR�b[-��a�)J}Gj+7G/_�SD[����3y�p�tv��ֆP���T�H����ww�̽i%U�M�*�ͻO�]2�j��/n���l�!�V�OkE�@������D,��
iA�OO�����)y��� ��u�&����i%l���Nz�l�U(�Je0�fA˽�3��O����'xK����T�%H�n�~]C�	�N��[g=�+��f)T�ێ�|�Ou.��@"�:B�P'�s�;�%�t��י�S�Ӳ�m��n������Cf<�A�!k���ljڪ]s+���׌�9Q�5w9җxՄ��[-�Z����݌� ����ܮeSɨk�=�2�3`���ꞡ�fz�Ċ)(��t��,�F]���l[��ve�N_M��y����`�zrg����{�<�[�(҃T���k�c�WM>]� ��K��8J��8�dt�H��^1����9���u(������=~�m�1��}]�V�;�2��+�ᮬƤ�)������@��evI�AG5v����}?'�����YWW�':��`� �s�U��Hs���՜����h�u�5I�j��E]0@�^��'�mP�1�o�J-7;����n��3̼�@��F�_̶/��8�Q}��8��u���� Er�e��j����fGPe��4s>;0A�uG$��v��i�<���[u�9���C�Y5$w6��%��#���tF�t��z�N2f� N\]��/�Cf=��%�d<�ĉ	y�r�U�s:X1Py�S�M������9'�E�nl^� �!�/��J��U �9��b�]s��"JY�!π�f��3��i�"ƿ�U)�^i��ZR����R�$u��*��g{�����8��,.�_��p0��;��j�ɪ1t�r���q�7|�|8���<�x!!���r�Fi����=]Չ��ml�d�͝<�}gY�w�G�'�R+��4�+ ܷRf@�n�B��B�P����h�t�k��ۯ�KpZ�3��m�$��T����[!���c�F_���	P�{���޹����_5���?b�?l��}�S=�2�U�a��#4QKG�;p\��j:��|�n��b%�;� �W�8�bGx��h���w�`�gJ۩)�w	:��N{��>��T���փ\�Q�/�)W���X/�1Ҁ;P��̒M}l�q�a��/�:Z��da#�ՊUv��+T.#Ao>���0�H�S\�q�%��>���炵!�="Eq��ؕ])REww���ë���s����U����ob#�8k�,;썔�P`�κ���刞�}{R�'t��	�Z�X��Ͽg���*38Cs�,��Oj�gT�]ͨj���q�[U���}��ۨ�Y~������|�h�pF�/6��HY��}�D�n��v=G��� �Rn���2{�dv4���[&�Ȱt�&�y��~�#$9� V�*&H�qn�7���,u>-�i5�.���Hib���,��W��:e��� D�#�c�C����rA�ߍ�Hl���{u���G��� �Fb}j�ѷ�׻������L�0�nO��f�5޴CΙ'��d���S�Oa��BP�Mzf 鬊�H�}�R }��b%���qW�+ja�#�RRZs� f���o�qR��mGY��
�|S�\�
��ۜ��.feH�Ӟ�����eC�|�� 	�#��{��3��_���R��ܫ��tOk�p-��f3ێ�h�N�ü�����Pb����K�p�q^MM9��=�h�,��Y#{�����ӝ���=a��!n%N�KF����nnđW��è�JIb�O䃷rM9�V�7d�vm)��Tm�Tf�7n⶗��+��#>�!O�B<JFUA��F�(�c0�N͒�)��L�$p�� �F�lDm�1oBT�L�x�����e�uȾ���G-�<;�Ŋ���S�G����/#��i_*EXn�8�n���� ��ӵ�dl���$2k�"[����[>��4����L���x�L@~%�gW;p랴x��[��m�0�� ?��W�k�u��4>��No��_pjޜ��䘣�����O�0}�p��y���Ϊ�t2��r���H#wW��%I�
��r]^H��6:d^J}��΅��\]�޽L�6Xo%�r�I�ds���3A1�X�t���{��'��H�w�9$=��r�[B%�}&ݒ;IC�6p�+�'w��5�)�_)�Ee�8�y�����xq�cq��J�EO"4��]�}��f�O��r�
����rX5mM�0�ُ�Wus�7�bz���>�l\�ÁL�ύNADxUd����������$k�X��ϣ c����7���o6��Fūl���FO��o��D�|;A�c��+,�E�}�6��g����8%��K5�s+ze�Z��m0U�Vͺ���4 ����Y'�#̚�\V���ZO[FV�ģ@%paȴ
�R6)����Dy᪑p�����]���gHl�q.�\���!�Ƒ(�nm)L�e�
�l\�Ot�qE)l��*d\�ytc�iAb(.��Դ�d�ӝ*Q�|���T>n���f�c`��}F�X.��@�&Q���F:'�z���窱�"%��nf��?��S��n;O�R4��9�yy��| �f������?}�ު��G]9���$!�HW���85O�9�;	�f��={&��{������l������3��-�Z�4�g��:��MV!ݷ�PO�Q@eo�|>Ǭ����zc��cQ{���wS<��0�������oDY�{�n�st'6Q��,y���b�9�f�6]`�5�q�,	Ե��TV����Nt۩C8�Îb��������@&�*u�wV��$x����D�Dn}v���:�(�g���}��R��c�u���[}\Z�t�ݶ�:Øv_��(�L,�z�l��w�$��x.�-�^T�$�w}���.��3�{%�gft�):��M-�PP�c�	������C�L0HԀ!p����7��qmY��Qc���N�ѫ�we�4�Dw�$1���^hG��ml�>��ԃ��V��ٮ�쩩6ݷ��/�	7l��8��`p��4sPRΫ�9$��$�g�|ܳ��H����fƌ�+I,tI��������|��]wXU��Ժw�%�;_�l;)~ĺP�%e{Ҕ���ƞp��{d_?p�5!���'���4-G��v�h�.�v��/��	Q��W+���^I��o�'��/�N�p,m�3�V?�b�%�|A6�?��gc�ʱL��@�}��Bpt����7�U�&uD��=�P�p�Y5�F�Q'λoz�o�ˏ)�vO
kF�h��AaB����������ٖ��V�\��j���)�ksq��6Le��.��
8�L�1�{��A�s֖;	p�`�������e��t��hx�@�L˷����TK�L��`~�V�F.�r���zAV�d�[Nl�nY����5>7vw6zi��L��Ȼ����%�?&�n�^z�6L�{���)����#f��J}�n�vd"��!o6��\B���Z6������[Dm��#�I7JH��ml����F�.+7#d%���Ͷ�!�p��Ϡ��R{�뒵B�,R���'�����'��v;�2$�p4�/Ao2�B��q^�giU]��������G�v�����4�C���-�'`r�ޯF�T �9�9ܹ?qz~�w5Sk�����@*M�{��[	C6t�\�-��S���+߳��g�q� ׅ��!�QI�=Ҋ�;#l��t���%���)x�I�n��=��D�'Q:�)�r�FO��{�6�!��W�����!�ZcjV��MŘ-cj�����-��K S���<���.�^#8<�wi�B��O��?INoթ$�W�;����gL&���Z���|�%[�3m�7M7�1͏kh
��U�M1q�����o�e��;���z]��15�䄙�]�_�U��[_���q�	�$qn�^�Ӧܨ}��֗웪	_��u�p:��\�� �@�ڭ���;�f[X��$H�[cKY2:��ޫ�B�Gp��dbgt@"�y�)��������$Es���Pf�S-��,m�a/�i&�^_OE<{a��+���P��f	�hŠMC�{\�����Ԋ@ʺS�m���\ۙ,�
PE��W�Hk�1�"��Pn��~r;H7@�J�)T!�>�y�� H�gB�8 7]*��k��ѕ�^�D�ּP�b|_�>�AI�D���e8�{~f�m{1�C"*9�+_~�&�2�0d�j#&��#o�{�RW���-�I+7���ܼ��S�+y�z/��D��-�+������h�H����膈lxV�<��@ӆ@2m�HAn&5l���8� ����z}C�������{��?���W���~?��9���2��t;F�эl/{[�y�n��<�Twl^v{U�W�����O߷q*mIN�+����E�/Tf�s~�g����[�f�Vƞ�Ɍ�����_�3�mc��e���%�j!�QFk���������C�]�ɘ��<��o�S�2�+4T���e��g%�p�@#�,��q�c����!=׶v\ծ�P`�{㾪X�i��<��x�g���O�����Ggbg/��
\lZu�\����,U����NvMR��
׋xF���B�m�[�t|z�fsݼ�^f��2ڽ������o1qN�w�K�����;	{�(�(�i�F3�s{zh�x\�@�e�A�}v�\�zi�Җ\t���!'I[�u��U}�����1���1�P=9=�$�Ʀ�ݫܾPɤ-ڏ���Xf^��N�$*��C���6�ZʨE���¬i�5�%�x�so}�ȃ��8a��Ǚϩe��x`��a��ki�q��Q:�fh�!�@s9�Ff�u�J���כ�F������Lc�yG3\w��I���AjSL��ïE�ۓ;.�)SU;>�ݓ�J)dd]6�f�j��Q��ou\Hq�xE�^e�M�+Vͩ�g��;��Y:��֕u�|����d���\���&��$.{LS�*]� f�܉���U:�5���ח�x p��0���j�"!�N�l�i�S�tN0	�(�-N���,#F�$Y����J�]����1���[�k׸)�'5��s�V�c�W��Q<�*�9
�����s&ɑ�����Y료h���O�(.�kqÊH&�r#L�i��E��Ε4�u��o�[���e�� �}�a��-l��bb�A�V��5DB7KnP�k|�S;I��h4��9�1ȗ�p��X�o�7�E�=Q��2��w�������wb�$Uq���m�i9y�k�1:�MpMwƥ��k*���	Vxf�Q�s�D�'U�����d�5N�$�c�"Y�wk�f�U���.�7�`Nd�`l��eM�Q�,�S�$w��X\��o"��2�y�k/y�3]�S��k���5��fˡ�dy;[ɯAB�!��d���*����'��&5��N�M��)vm���F��XIbtPq�Ge�Ӳ˾��*���e��q`A<c+6KKuU�+m�7�K�}�'���#dKjՇ>��&.e�1��u��O�]wWW���8�釵�K�d�f��U���wB�v0��(\=!Ʊ��M�G�ޙ�<�$����]u��tTs�C$ӊou1��]�Dn��o��H�Xn����x9vW&��(fg6�j�l�G�B�|��,���������nt���2�/v�+*�Xyr�o2A�ݎ9�wQI��t��Z�b���p��U��K�e��ow�F�}��L��j֮��Y$�2�o-jq�z�:���t|	�@����@E
Ii]h�׋E'#E��AX 5�&
����E�ƌ�Q�1S���V�th6����&Ũ��VӵT؛j�j��-d��j���	�Nƨ��j�#��h�<�10�EI�kbj�ՌV��M.�kEX�CIm�����EA�i6�kh6v���∱V(�T�V4���լZƶ��#Zi�clն*5�j5��m�S�cZ1�S��"hѶQ�[�AF�kP8�����b��)�Fتj���M��KF�(**��c5L��T[jb�N����Ѷ�m���QZqb�TTES�#F�cM%D��Ϡ��z���.`�b��\Ś&Zd�����3�cˤ)�IF��$W2eneC�*V�U����wa�p�Nۇ�-9�R+�A�z6Mz:�(1u���}��	DA��	�D
�TD���`��L#-"Y���RLj�&�KȤ�#7]P]���,g>�~^�x��Q25��3��`0����[������^`���J"��˲�q�#5�X^Iݓk�`�q�ޠ�{��?�xPZ�j�1V:`��<�::���]i��?�d\�'��Qꈎ笈�1�i��h�,;R1�ܽ�E� 9�a�������M�-�i�Nps��&:����I�F��i�̈�Yz_k�i�~��m�6�ȗx�����ɻ���#b�v}A���^�!�C³Cg�ѱ}f�͘��������+_�������;���)s˜v��B��OՒ`���=�0'~q)-g��|�g=����x x�xUҟ�s d��*�æ9B��v��NN�&��qBt�\i��yަv��$\��w`���MۗxX�j�AM�E�j!^���R�>��=�^> �\i�]w%��'�s�a�.���>pu$)<��Y���+Np�1� ��DI��c�i|7en]y��g,�����f��{�U���J�Z��eGw�v��SN�ǩ\80�n�K��+S4u�'gfF9��x'r�s��zY+�e�%+��v8"@mv�\J�}`�P�o�/N��l�t
�L�@�;fЅ�,��5��ẍͶ�l��fHܷSV�b&� V�p�ظjD�`��� k24�b.q�v�*��IU?Tuө���,%Ԉ�D��'���3X�_�5v��'���[d�'Wg|�f<m�A�!o47S�?{[n��]��a퍑����m���R&�-�k[$�R8n����9�3�n*���Ҿ�i����݆du���J���6�yWf't��w!��{a/!{a�
e�b5dq�F�rR�::V9L3OW���+���h�FS�Ł�pQ�t�O�M*0WP/�W$�.�У0dD��t1��)���N�m����C<��"#4��=��q�ijuԷ�1w�(j}=\�Uy:K��=��:�������Ww���b���'W�f�"�e�_�d���t[��i�KE�Y�z��y�q<��F�+���#�z0-Y�qP�q-�R�:~&��Vk������:懸z�v�]�.G�ݣ�j�]������X@q����IWRc��`2�ۃ�\QG��ѧY$�o��=^0�ï�ͤ����c�y�Dd��ڍL�9TՇ�x5��|�'�}�+TfZ �"BD@y��Z��s�B��s6ёW���s7��X*������7����ê�����	p�To:8q���y��T��Ţ��V硬`����U=^��Z�1z���:��t>�P�q�c�;�#�ss��EE:��� �=b;��Z�_DG_�%�Z�a����xقcT����O���	N�z�N�{���v"K6ޫ�n������nI/	QEO�q��[t� ��s��]t�zc[|�8dㄽl�m�݄��䒶�S��#gl�s�5��xh�De�R�)�F	����b�J8_}�%j�Ķ�!o>�^6�F�y�n�H�ѯq0�Os��=P�����$]J��G��o1�%��o��S�CF��=23x�ԍ�F�c�%Pm��0��;\D� p�Vs�hۣ���1.��l��;�.]1`60M�����{Ǎce]��T]N�� 8���v��(������[�g/UtYB�-{j��C�d�&i���C�l�����ޯF�U�4g�:�+����ƫ�������Ǟ�H�J+ʷg��:Xe�#7�����N���ZM��D\����:����t�u\vF����Oy�go)ڧ��a��,�ˣ�n/I ��JN�H�������pѰ� !˜�n���b�K�f�C��>"�y�Y�d�s͘+W=$H[�|L@�л{8t�֗��sh�g�K��C���f<��M�6;�Fe�{w�H�4��a�&�\qS6�8�#�\y~���
6|��ڷk�uۻ����KCL�Նhj�\��=�k�Y�r�f���M�觏l5��	@{�4&c�>Ҝ���[�k[z��:�XĂW+
�i��"��5)�H��H{j�#vp���f��ΰi y �yb�P�W�̛�s5m�-`��Ih���1�_�7�E�JZ��� +��o�&��uǕY/;�n�;���i���LdA���^��0���&��>��&_��N�wy�ɘ�t�-�,k�*�杵,���#�R����{|c�p��(��x`pI��C���k�9��!_,{�ro���G�7��#���Sr���!��t��.�%%	K\�9능Q����B�,ۥ�x33� ����2D��mq��)+�*['gq١��h�����3�����]9��� ����k��EpP:����M4��1�\��q�۳��6篗��{7tw_O�6�
tp�Ljٽ�,�F�,�<'�st��Dsޫ"݊�jG���3U�L�E�Q���a]G��Ѵj���������;k�u#^:���H�,/ ���H4�����7�]��.X-�殷�g�a�|�	U�WTM�2c�׻��	R��g�>��Ol��]?�f�=�Z�¼��/B�8Ҥl�ɽ�E��Y�yN׉��cc16�����u��,%�0>�v��<�Fl�c,�z_o��/��w�92c���U�wr�c�KT0�n�R:�>�_��B�dĬ tb���������؏�����k�S����tŨj���N�N�J���hkd�̚Fm�	rĘs�f>��e�%ƱB���=�I��&��Dڄݝ�����si� ��ȳ�`�B:�dnv=w/ֹf��=�s�q�
̗�#s`;un����;%f>�Gv��}�v��_�y��c���<(��?c�hW@~Ia��U�2*�a�l����W\"Go#^JБȴ
�S�s#%��AseT�����"��E������TJ��{��!"��Ƒ����6ԁt���۲�{�kw�F�4�
�U����F��5�}��
��'�M�޾iiُKR���O$�4(��
�\#V��[:�@�^��z����F�,����=�-ן+�Վj���ЧEg����VZ:�.���,���v���>�QIP�~�S�^|�BC�W9o0N���[7��z��H��^�).eĶɒuup�v�=���8���b�B��{:���a�A�E�N�>m���R�l� ���;eOsv^¼�y,3Vv�������!�r}��#�z�b�U{�TQIG%��&�� i������pVZO�Ƶ~i�k��H�B@sF�1�h'8�h3sI�b�hv���g'Z��ʹBMN���B��� �����}�d!���\(/Y�~Y��p��&VY3O}������0��"����BZDJ0��H	�YF>89�W�_\��Q��3`����K}>Q�s7����>���������{��r��W�KSvh3�����)Ƨ����z$g�=�/M"�v3aM��Z{bP]�t[0�/�(�yU;�#6Cn�|����!i5E�i3z�f6�2�;�n�=Ƽ_e?�1��1�h�AܿC?�s?�.�8�-9�VNN�����������2x�#y��[��Ez��l3u�t�3m7�8���b��uھW�`fY �"BDF�h喻Rt��%�1����A���}"�{Dxp�{�^&����+E�)Q� ���P�g;��G8>�8��@�g�qA&����=Q�z��׶Zy�4�Q�U�O������z�R��bL;�h�h5ˆ�̓�\&�u �$�6d�3ʨ���Oi�<��k�y��P����jV��Ku�"HG�2v��\j7���.���hՙ���Um�QS�A�YB�]�E4�yZ�:_���¸W%�����c���6NNY$Jf�l�ιDMoj�u�z0��+���ݧ.#$ǑYMZ��-�9�Y*��V�I׫%~�;u�}�QD���(�1Ʃ�u=�J���MS��2��#߉��2�##��@��݄��A�T�L���fe�]���|lp�ß�0�Z�N4h�G�AZa`�/rUj���ڒ��z^�kY,�3љh�En=�6�$0�I����"@�2hv%U㋢[j\�ROx�s�sם�|w�O�0~��7�%�oTl��HK/�,g���k�[�GI*�w(�*ݐ�t��`Fny��`Wm]��[�Wo'r�l�ۮʊK(�0�A�[C�u+U�v�Σ����X�H})6ۙ?*џ��j%��氣GR4��ӎ�3���v{=_z���י������X��!�k�'��68[X�Of��9Vc��^�5�H�Ż	wg��Dn�9�n�8�[�!H�f<��7����m�������{fB�M�E
��vkM�<�λ�%1J�/��� ����5uԟ�����5ʹZ�`ǔ�M
l�q����` �oy[�Y�T�F�6�gt]G��:��"	�*Ν{-B.����^��׫�[�8��<Y:U9�B[Y��n�q�&����e����Zۂu���r�򅖤�6���v#�79�g�*�pdl�[�7�I4F�M�����}p;���j���Uc-l�iRHkݲ�g���*�׾}��&��5!C�Lɋ�����x�87��G	��z23�U�)�%�^-��SNa�܎��%����%��U3�`��}��(����"o�O:�S�к���%-�jږ6{U�sWeVq""^	�馡Z$fB]lE���~�����N��2Z���>�[�#M݇{5S��s��D��y+�2�N������?r[:Jc�n"_�IA�T������l�/pX��Uy��9�o.�TW�6��|�E����D�#7;[}]C�-�	��^v�И��ٚ�b���<�)o���r�(�y'vM��L7��X���0S��-���VS,��o^�T9pŨ���[�l5�R@�ٯێ��$-���Xf�n�#}������]�H��k����vk�e� }]l�]�V�it��X�c�������z�H5�[�ڻUF�*]��oHȺ�,���g��S�i?s4���|��{���i�*A��]�uy"jiWL�1|s�K=��Dn���Os�0s��8�dl�ɽ�)Q���o�:�����{�d���C��@n�L�9���2*qç�/�/��:�c5d�U)���v�刖ܑ�#ݢ��5vp�t`G�1+*���odN�hNn�g����p���ĕ��>���>�Z<tVN�?c���tl�'����|E�fm����Te���k�� v�)Rȵ\��rY��7�i�1S�7�ۥ��U���Z�u �r#�#^H�H���J�ޖD��$6�n���'���Ń��s#�ɨ����W�AH����q��ݯ�9����8�nS���)vf\K��@Ԋ� A�V\-�@�ػa�㨻訥�ӻ*7�;�5����s��O�[<�NEO�;���3����_�����{���o����{���~?���x�*/��N'^�k;�:��H�G�*rw�|*���})E&�֥�G�.�2>���W�'	��V�$�:Ьn��:���rS��y��%Gԫ�̼VX����j���*ĽZ�)�I���`�ͨ��bLdx0Pud�4M]��2��X�k��'�iYlL�\������=n]�e@��e*,�QT|�.�Q��σ����?dy)r̗��XޡL6�3;�V�6��� s��Ϥ���{�ir�ie���pm`k�lV��;r����_f�{�^���xV�j9 �o�Ԍ
pt��8uK�j� <�̭�4�V�`b�V����qP_{�j����,Y�D�w�C5�=т$�rƅ.�gU��\fYl�������6���C�A�����0c<�\��9I}\	����kA0x�5�*V��Y���4*�Y\%�295M�ԙ��Y��xB}v�;8Su1�]�V�����9��Rܡ�ter�n�`H��ɖ/�q��$T�e�A��4Ͳ�oS,o'��X4��;�;�� �RY��{�$H`����~9�����jXy�R�!4o�kH���&�<�� hԒ��_g:��"��3����YG��݈����L���x�M�#c˼v4���e���K3�ab㦶���$�{b��v���y� %��k�M���XZ"�R���
�%��P���w��>|G]a�!��]�'*(�m� ~�z�X��w����*���B�{W{:{&6�'���s�j�1@�fgrq�.����t�]u,�kL�������'������ͅsv�:�bO5�n\���(���۱o5K�E(0k㉞%�E��*,�)�Vˎ�Z:��2��=���������
�����>��s�&�)h�E��Ҏd�b�.spo���8�0:*�l�ǩ�WF�GM����`�hR#r��xص�M��u>��nqr\.c�6�<��G0��O�wt����'3^VQ��vb{�|.�>�n�=�V�S��׵[1E�lQ������Çi!^:K�3*��n$D�4���PJCx
�Gv�4pEú�ɴ}��q�%Z�2�3��Ai�{��'.�K�ժ�fĂ����K8�f��4����F3�̋C՛ym\���6���s��Gd։af�qBX˙��Bmq�9VbқZ��n�h疶�Y+��p;��-�=��5���] ��
n9՚��N]����b�s�^���@���q֙�����j�8����h�ڴn��Қܫh�J��7��'o��r���!X�L��gۋc��(M��b�1ma�ȳ��v5��΂�nAK�[��.\{�lT:�œ�^�//2Ffwpr%3����wwL|V�M;h"����"�Z3j�X�Q��ѭED�cU�A��N*4��ъ>nr�F�b��6ն��6t-�k	����q�m�ٱ� ��[E0Qb��4�E��
ˇ1PU$�"h�i%��*���LF�h*"�X�5DEZEm�*����c�PSk2DLRh4�MEi4V�$�U�TP�li��4L4U%$�V�Ik�D1DAFڂ**"&b�����j���钦�)��*������ŊX��`�	�����(��64�QDA$UPU�TT�A�Q�k;f��(���4AMU�UU4AQ2Tl����u��"���b���$�I?	 �?|���8-�u��l9(X���u��CN�no+t��D��"�؟Y1n�N%o;��q^��!��j��]�Ңs�S�6P�������^'�T
o%T�]:�. p�հ�kMc^gk���E��+ߧ���.���3�uq6t�x�m�Y;��^֊�Τ��8�`�� ��:v�풧yR�a�ŭ�{eM[�P����N����v �������r5H����Ɪ�3ֶ$QIB]׹Wvr{�c[��M(��v0�B��t:�;3����u]�3����{�Y4(̽���v#�s �J=�C6XP���C{\�:{&��1�d��Y���z��Y�"�]-�˺���2v�l�{|Â��FpOa��/�Vv�էm���D���݄��UɎ�&:Nٞ��Ch�R֍g[��V������}5p��:=f�ė#}ŻdZ�3��r�/3G�75���l(�x6�
"�d<�ڴwOfY�<H�%�O2��$�1K��blˊ��Ϲ"Y��Bd1��_���~^��mQ�3p��o]k&��'J�:&�ed�eb�u�Iv���*jX���x��A�]��^�:�a�;\kZ���x���t�$��=�e^v����wR�;�G��G�
�U%o��������(�R;WUy�����s�!-�,��j%��b�pE]l���χK?��f	O��MD�/�H��Ɔ#�V^h��<_nȁ��a�mop㶥RGZO]<9�-�,��;����oTD��Y����7�6�bP��t�% ٓ@�*;W�4�4�=���%C=��g���H��2����ԑ�^(�8��S�n���}O]������m���g�K�7Qp���� ���H�@$�n�)3�%N���2Օ���=;�w�r��H�t�k:�F��U���%V�\r�9�]�"-��̋�|���Y��d�)������	�l�M�3��ؕ9��f9�� m����E�绣�{�'��>&��`%���a���{#e)f�:�i�9ݓ3�/z8�;u[Ǖ��
s��a e�#3�l���d�4�rF5�54Ҫ�nI�L�l��8dʏ�{ea��jb�D��G�H��v�5ww���<~�Q�+��wf�Qd@��=�����%���B�
T���\�Q	x͗�S��Ei��X�m3�e�\���C�k{�E������Z*57
��:���j�0�T+�{V��V��i͹�?��w��ӹ:�7��7.¯��4���p�w.:���9CTd�t�Ӈ�����R���ȴ���)��<e����x���L�<[���i�Z�����n�������u
��H�d�`<*5�x���љl�n1;E�m<]��.�|����.%���"�� a6�����l�%���������M��g9��&��A4F�M���#�� �j�J�(e�4NF��{�rr���ؼ<���Yr��c^J�sNdl�ؾ�y+����\��^�.�t����s�Ȍ�����䝹��]��;��*)���A�a�	ϡ\��D@ՄH�]<�)=��JWm65�a�ؒ�/�ۧ3��^���ճ�V1�	G[w���]В�?�j��)R9/d5�uЈmK���pe`��eE�2Ue1��Ui곚�x�������S�R��IVH�>%b:�������κ&����t������q��H��Tf]�7͹����z9f���ȥve�m���Z��
�gp�1]��v��_���{SJ�����nS./置z{��L������P譎pAFij��̶�צ���H��#�d�FQH7J����}!�l0� �n%\֌��5uU�FY�ڧP<��@�skc4��~H��t�f �m�s���O��;�ARC+g~�,1��� �����rIF$R��	�6��b��/;uB��^�~~�>�ya���b5dt���[��"fxPo���l�x�ǝ��-S���F8�R}�PC�!��G`nV��u�s�;���#Z� �U�3��-��2�ATt�؀:Clo3�΂0���zܗoa�Iۮ�����t�e�q���ܑ�>�HA����x@Y�̙eJ.g~�3O�����__�#��<Xƞh�`�;�#3�;��a�T�L=���{f�0[��7Hu�Ў��c��WHD��4�9�WJ}�N@�.f���2���ݘ�r�3���.ᢢ��S��b���5����4�<ۂ.���Z�G��� ��u�3'P��@��<��K9b��edPxXa���]5b��3
�p�r��w���ɳkI,'V����k�C��{�4�,�ҹ��v:r��7��L�ڨ��������W!��4�$t�ؼB%�'�yyN�
���^C��������T��Sd�S���B�E�U�7{�2���Ѧ]�z���U��ˉutU P��xG��R.��/{�.��n���ףR)�IJtc˾�+u��g�S���F�8zy����s�?:y{i�HKBJ�����N�g�= �������V�J����㑓n���6��x�4�&@'WP'��Z���I@����ޙ`����F���J���J��K�������秦��.9�M9�c^�*�����^������#�{�F���"�J*����[)�Zm����t��MT�5�?������u�vgUGg��*�q�-���Tw������rd�߫��ߙ�R]S��5�Ogz�3�f���0��5}'Ы�j�i3���e_��k:�DtW	��Lt�嘠̀ڭ�<����%��� �9�+�����Y',R��c�l����n�h5���WSnv�ƹ���EH%�
i�ʕ�NK���Xeg,�?�h�=�y�L�)�=��s{��W���G��i,6�pa�;�;��]�l��m��;Y\z�/VvV,�8�w�����=�i��lt6TN��N�?���x��g�
��-��kk�)r�޳fOG	�m2	- �/ie�r-�\���
g����Q-3��4���2�y�����cF�튳��Ka�g�b9]�ط3��aD!F {�j&���;U���&�e�J�,�,���O��G��Ϋu#���PJ|�2vozh�{�W��3(�R�\�3�mY �6�$q����D���W ���Ց �"�����9��s�<J3�lɣ<�����W��&��Z�=���1�����VGs7Hd�"6�F���#e�,��T�*�=�������?vk6����P(P�DfxA
=��F�@݂��A�U�=\�o6�ܮ}�юͷ�L�iaC��-�o5ˬ�]OC]a�39浮��S�U�V�ԛ�m���ܩ����D�}�*���W�*�'n�#D	徶��F)�Q+�ǻӭ���j���kd(L�f�ۻy�M�W�1�6Ա��E�>a��ӆ-�����p���EqY���V���u����/5S��A��t��ʡ�_�
��h�xu�j�k��m�_��y�A��1��]C0+(?΍���M�};�c;��k�v/k�.4���r��IE)堮�y�v; l�0Ѭ�m��uC6�����|���]��58;�*�q�U�>����e�����t�����������ޡ�;ÖzvWʒuXj�{���(���#��3�B�kkv��֍\]�g����r�0!�( �n��ԍy?NW�FOtl���
���ǩޗ0w6�Q�A�{B	�#o}���ȭ\h$K��]�*W��f��|l�7CLo9�dj��㡝�E�uF�M�7�;q��(L�Y��VM5��":+^r��d�ӤH$��:����g@�!f�Y)�}�͹��xݸ���ُ���x���=!"t�i��#��]��p�BWy3��g�4��r����"+mu`t���U0�V���B���,C��DF-yY|�ie�2|��SP�s�P���<-,��*M�,�Lz�9u2�2���@f�o����1F�#�Eì�$M3]un�GtzQ�E�P�N-��{4�;�y��&2r���J[�UҐWcO����dۜ�!t�%�d������Ľ�cΣ��K��*�y%^�F�S!�V='vr�����@�~��J���ZȻ� j��]��y�]�A�m3'����.\�i鵈t��<��m7D�<�;�DlB��"���ٷ��Opm,ʾ�w��� �^;&I���k�R5�����[U�OU�H~�
�i��.��+�qu�9�J�T���R>��}!�o�BkC�Z-��cj�cfff�M=
�Pa#zah8���:h괉���HO�3�ڱA{�xɪa��H���f��P��;�q��]�*�J1>����mtwj��O�Me�/����W����"i�X��0*��;3��t�~��^KI&e�C)Cb�����./�k|:o�]�A�t�����#�
����R7/zV�Z���\]y�O,˅�����i���A�5���ҁ=7!�&T'X-��H����S�W���?��ޞ��ʻv��*ݾ������&'/�lH��ރ|�yFSb��wfa�N��g�KvV9�U&��oK.f��`�O:�����F����3:��\%�	$j�KQDJ"�q	?g~�잆��m[�,�"�Gc,w����wݛ�o��owξ�]���l�ѳ�/�u�h�ú��B��9�r)��j3���sݭ�8�s�����,v
��t�b��zS5�����!�NK���)_k��!�x��V�"��Pɢ6'N�n��ų�o��ݛjR�m�V�H�OOU�zuCF� k��$��h�k;v�R�g�=vg�M�햠���p���E�N�e�oOX�}���ܛg��n>ђ7��ٓsU�6-QB:�	�4�ZK1����W�E�^OlQ��K�Ur�h�*��r�u[��g�]9x1�`�_<o,�6M��"�7����^n�h�J�J�?T�u��|�-l^Ȭ�he[7��6^�@~ N�79�RWϾLi�L�uux�P�o���8���@�U�eڙ�}y��5q0T��br���U]��͎Ҕ`#���9Va��kʱ�������5$��)�<�ߩF��7��2S��Î��{����A��s`��]�E��⣻���-]��D�|۪��f��g��Ђ����;1�b��|�%Mr���l�&۳�G���Fm�m>�5�BZ[��-�Z�o;��#zz�b�-ֶ,X����D��̓�k]��N�\��=�.�Ɵc��!����;�=h�{Z� ќ�Os[��3M���Gt�J 5C6XP����
�!�x����w�	�	�U��E�O�=�z���zB}�#4�վ����O!{��?;ε���9�g�P�e�ٟ2����8��\�����l�Pc8���q��[�����[?�c�}��s�,���u�8��N׶Ig�hE���z��c�W%i���i�]�p[���
�>գctǳ,��=�yٷ����=�$<�F���x`�k�M��/���v<��Z�5u�|=�T�;cU�c2��2�Ď�k����Lj��W5��V���3��b�s�|���M��2 U�U����,� �r�(��������U�B�*̋0,����2,�22���"�0�ȳ"̣2���2,���+0��� "�!"̣00,��*̋2����,ʳ*̋2���
�+0,²�ȳ*�00,�ʳ̫!"̣2,ʳ(� L L0�Ȱ� (� L L�0,��*̋0,�+02��� ̣002���2,���0�³�2/�>G���fQ�VdY�f�`ex����e��|eUp� ��� � � ʀ� ��r2*�0 ���(�ʊ�"¨���xx�U�( C
�(��2�2*�ʪ� C�p 2 0�0��� ʪ� C*���2���� C  C*����0 �+2�ȳ*à��� L2�³"̋0������,���*�00,��*̫��2,ʳ�02�³�+�7��>����?�PEPQBaBd�_!�������P~���������뎏�����/�,��eqd�Ѥm��ܒfI$���q?@������
��H U����>���'�K�)���Z� U���;��~$��=�=��?�'π7�����b��~�"���*�@*�)"�P� R��  D��2 $�
�)
 H� 0 �*�*� *�"��  B���� �?�@ �>q����������(�"�"-@+B���@�������AA��? ��?����Ƞ�߃��o'��>�����ȟ��#���X�/��~��
 *�؇�O�鏓��O� U� ������=���~��=���*�?�����_�|��������O�|~��<� U���?������ U�C�~�`=}�������?�����>�'�8Xz� *�~g�?����
 *��<���􇐤�����p�@�|��X?�������>~BO_��( ��>(!��?$��<�=A��������tPW���g���T���_F��owY!�ї��d�Mfy?�:�f�A@��̟\�/��l��� 

��6ƀ�Rl�(( Z���
Z�� aT�BT P�٠b$�Z&��K+Z�M�F����3Tŕ1-ME�J�Jڦem6�T�ǳ��ac��"�b1e�[[6�+%��me��le���3b��he�3k2������R��Z�	��2�-��U�j�4�
�e�hY4��Z��IU�V��n�춭P�mm[m561m�)��V5V�3l[J��km���  ���;�u�j1�v-��u�[�
�UZ�ln�T]ʺ�:u�ҭ�[p:ݚ�.K����Ӯ�Fw;���-ɻ�(5����-wk�۵��2�F�5h��lҶ3Z^   ws�СC�hP��(\{���}+B������>����cB��СB����n���e��V�{��� ��ݬ�9�֧I���kv��l��q�˶�٭��ڻv3��T�n��gwi�4�9�IUI�35���Rd�   ���
�.MN�u�*��5;�7+�5t���]pʦu�T�j5վ�z�����
�v�зV��)�v����q��ݧ:=���k�ni7]\ii��靦�%���   v����+����m��F�]nkN�6�k�5;�{�{�Ӭ�uˮ�ne-ݩ�Uֺ��� ���m-��wK���i�I�5E�Qum�kJ�kkM�2Y�e��  ��*)�m�qө;a��\�4�6s�����l�*چV��V����m�薵�]\�1CW8ܠ���VԂ��$H�[*ګV�j�V֥�  ;�Vd����ᢵ�6ݪ�P�k9s�YkTv�v�UI��W[%*cQs�pkEK���ښ���E�ֶͪ�]v�Si�heJ׀  ��z���F�ٝ��]��r��	�.w��jv)���Y�kr� h�uuU>aM��{�T
(�{S�Pzʒ;�ͻʒ�T.�5�1�gFu�ڛA[Mc[f�  x�X��O}�{��J��A��ۚw)QA��{���{IPot��B�{��䢪�����z�$)n���T�Ws�Ǥz�U��kh�b����mh3a�   ���W��\=(*�+����UJ�����]j��;�-��*�[�ٔ"S��ozT�*���3y�4B�GrTPGf�Nꔉ@{]O*�hdf�m�Q1�e����  ��}ѪQ$�y7(�{�H�I֍�e�%;iW{��� $����ʔ=`]��d��U{��޶(�J��������y���(� �~@e)RL@ Oi�����di�M��d�R��  �!��T�@ h��&�T& C@�R�&eU@  �O��C���?ο�����J����;���+�a(T[���G],�5b��?W�}�W���=[�{�v[l�[~�e��e���[l�[�e��e��,��,����m�������?s�~��������(�J����BХ4�ȴ1#�/�]�*ˌ��u �n-�j!ͽ��]@K�n�֊Yv�V�(ћX�e�3����F3l�S��Z�ZU��(]�ŋ��H��yÎ:*�e\W�q�ݽn��QQj��@�I�V�%�q���J����*��j͸q9L���+�^��޺
ݬv�u��1����X�q�V2�*����ta(p;�b}��iC�����,����aZ��r��p;��7wl�e+ں�*:`�K�%5rl�˘�0,y��K4i^��ٺ��m.�ڕ���2���q#Y�s/�b�8a��P%���7rJ�R��+�DS��@Sn���Y�����L�՜z�c
Xk&��e�[%��lD�]�f��(��Ӳ��x�3Dܻo�BՅ"�V[Ee#����k�m;YB�םʖn�h�dR�	g��w� <�(-G�MaR;���a�)�XwE�U��[�_��tY�珰K
������e���w9w��]GRX���J��V��h�EP�݇�&(�/=�tA�˦,Z[��
L�b� ��E7q��5�*K�"]�N��_Po�A����Av��Q�Tֆ�+1j���r�Ŭ����s�Zu�y�����OG�ʶ���30�R���:��,��_ْ�C�4��f���*�[�*�;���,d̶���R�:��V���
��F�bѶ�k�[��Q��na�5̛����K��b9	{�����e�(
٣~c���s3pl�*,��Ov7�2����;B�U4�����/n6v|N�����֌��^1/�RX6%��e�w�VK�C]7�Y7Ja-:���Ŷ��/VGg[�c��n�r���[�UK`��v60p��[���x���l��P�|wb��,��wڙ�I��2�'�P��6U����`�oM	L�	r�MsM]��r%j��9����+Sv���rZSM� �cK��&/�0
��#,Y�":�_J�ow�/hl?Mka;r���v�jҥ:Q<�4�T�[/32f,���MFTg˸���1��^ҡW���EP`������Z��ӄ�yWe!��hk@�tb#�K�=�wt̆�ݱi<���F�D,7
,-²D�L!AK�P�x�^b �S��+M�voQ\�0��^'C���tu�K�YU�͵y.���lx� ���:��y3`��Q��cu�w�f�B8�ZX��I ����]��PU	ݣ�a\+�s6� *��Φ�.�T�y2��j���U�j)���+u�u�u�B�$���w�
Xx�.]�9 ��B��<iS����[��֬��WV:�֮�V{�d}u��'G.��Ӭ��:vյozfe�#Q|9&� �:�pK��{˓Ջ٭�@.e5��`Km�!�����n��c+���<5�,�A+H�!v+kq'���J������	�.�Й6�Fkm<Zf�e�N;˫`�QM�ӡB���"��l����aZw�g0�!�#ue��E�B���5㕺�zՊN���G+o����\m�ح�`.9�WPlօ�%�,0�[����]E��D�� ٳ��Ҷ��Ai�:��h���*���X�e����hR��i���&Ƙ�nΠe��y@�@_m
L`xp�vI���;Zx��)�C���5u�m ��e)w�ͺ8XE1�5�Vf(�M���F��6�Rv�F�!)j��;{��i�V�T���&!J�pk����oEe=Ũ�;�*�Br�`Q��I�LȤ*i�S��svҫ˥�髸��[5���
�)����OyZ�fE>���f���&V��e*�Yt��6�h�8^*޲*y�x)�f�
�GF]+�����K��M7 ��pȒ'r��+�t�AD� �Qy/��y2��`6�u��j�[�n)�f�K��),���t�X�}��+�2����)7I�R�մAв�&u���'�hr� ��w�pm��kiQ*�]�
�-
�rѦ�*���e�G
Vl-�+eJ���y
��4�+l�jԵ
X��j�E�2�^0��;��ɶ�ɕ����{�����w0�rl��J�
��W ���86����*¯����y�T�ҙ8�!�8�B�Iu��5=��-6Wx�g,ab���l[V���Cݍ2$ilb��j��WZ�,��_Wʻ7ox۵����3��;����]�� �`4OQ�2��x{{7�%���g,;F��hѭ��㤶�a��p�.ɩ�b̑��J�X�a6��k�����S�K6��m�W����]���t읎O�Qj���k��|�Q4���}�8jTy�y���56[d-Ȱ\mU���E�ܦXX򝋚�v�e%J�E�VeITQ�X�M.�6@{������T�v�a�x��W�a�l�4t �`����ܶ���Ne���h#�Cn��=w���l]�K���zA���O�`�M�p�d�G�R��Z�w3h`�w�S�bGv�9A�d��vv�A*�t,��x$���� ����y�����p���%+ ݽ6ܖ�K�w���D�$�����nҤaAU�T6,��%&L�zw-�7i�ײ���4p��n�qm�/w(I�&L�-�-X��4J��*��!`l�f6F����t(�)��̆���G,�n�r�+�U�����$�1h���r���	���j9��fv���HQ�-X���ã�G4�x@�y�?(M�9yz�B6�a��>'.liV�u��]�(X�IԥF�ԂàN�B�'H�t(@#櫩Y�-��R����r�2���=�g2��:)�[]N�([i[Ԏ�������P\h1A)�p�5���s�Ճ16��ݛAЂ��Sjfskl8�`(���6+��^�4�V3���٣ͻ�݈�
�&�<GiWn�5�4ZW��դN83^���v��b����/j�hmU��˹x���_]������V�-�:��c+�����]ؽe�s0�D�\.�5c��W�N�N�R����S*͢Z�M����"�n�-bWd�6Wn��}yz�T�V,���Vm�.:!���P�ɘ3b+�jV�zjF��.	���x��F�Rں�2�0��!��T�*�WC��l��x�R�Y��<Q5����Ыm`,.�E5�2K�H��P�1���)�!m�sw�^���[&8�w�W�:�t�G&�ƞ��P�P�K6�@�?3n���AIͤ-*q����ɋN	���ZzݬuQ�{C&�cX�i`�5x�X�F�6����d�A�E�
��պa���02(�T��Њ�I^�tL��;�F@�2���6찵����zvjV�B�=�Ȼ8r�{t6e���R\oP4����Q��:��S[�)�+w*`�e�-������;��6uk�+,�h���4
��d3^l����w^!���KR��(&��b�Mw���B��k0�y��]��$7��!��-3h��X�ƫ��¤{�i^$�`�'^�0���]����J�k�����]��@�HFg�;�#)^��wL;�
M��ڂ�� FU��*L���`Ȯ�=(��3�D@�{�Ҁ��UMOY�VDͦ.�n�]kjR�E#V����<6 ?H6��xV*��=���xhe��E<;���]��V�"��c�{@�#�"�@���n�����Y����&me�.�gFn�c��(Y�(QE
����M�ۭWzFa/r�*T�Rf%Cd`@ˈa� �=�.0�\֞H�V�lK�GOA�����˩��4E��7L=[X`�L:��ו)�qZ��Ӕ�8��y�(-��ŷ��)|�e�{cf*���ҭ�A��K~ر���:�J��W���|���S7�Y�s�"��Th��\2�e�kI(����0�v��c��ZZ�Ԍ��m��E��:]I&.:[�b���t�f�z�`9�݌6��`�j�v^K9P5S��1ə���6f��/f�4
���!�f&�^f���spT�H4M�*��[���m[V,�x�	H���h_O����:�[���c�z�Y,ش��^��X��y���$]���X���E����Y��.�&��C]�0mV�[x�R�22:�.���5��d��̹"V�pb�q�����5����a�8��ݫ�F����Q�oV�ټ+A	��CQ�F�(�#��i����Y���*��$�"����E4��Ӓ���;d`9[c�!�xRէ���9y�k�B\��wMx��3��NwQ��qẌ́�Ѵ��j�6���Ҧu��r�fe�/^��j�Yt��3��=��	���7Y���[*ɗu{,U��Q�n�˸��f��o-�f��@%�T2�"6)�@�wKon�[N=��!��{��@S��ޛ8��jKu ˣ�"1<ɻzoH�ǷA)�Ė-;�F�p�uu]�w˺��U��-�I�E<��X��lB'��lq^�6�9,�QT�Y"�=�7X5�]�r�x�����ǁ-�H��0m���7v�o4�d[�م[��v���f���.��m�c�n*lk�V*�G\c�$Є��Nkݹ�H�)PGS��(��͛kiA��iQ��y����V�v�˳U�OvQU���}h\�U�k+6�SV)\�E�C�"s]0F^�%}}ʖ�,T�&uV��N���M�p �^#M���gkQ!m�z�@��c�!��'�#@9%̉(��6��u�)�Z��f�XP
�
`��R�8&W(ؑRMe㰬8��݈Е����Lػ܆Қ
�w짓v�8��/i%�'��ܼש�z[�tP��]��Ce��{y�
mc�7hͳ5���9��:Li,+Mț
�h�����
�Zc����abSu�k4�o4��J��-	vn�ɕz�޻�����Z�) �p���F�W�7N�ܫ�r��93}��)� 0N�k
�!�n��� �S���n�s-�7[�wGr�ϴP���OV�Ø�#�[�Q/275QF��T�'���7�+�y���n)u+���.A�:�s�Ũ�A��h׵���# �٭X���cz�n��9��eY׻�7�����pA��N��ܬ4[��Z6-� &�Oh�Lc�Z�涓pN�Id�v�{�+�Ci�M��u�#7�֟f+ ތMzZ͹��@0]�r(S���bʕ��X�	*��m��5{Ҽ�b�0F�OI�,R��z�׃t�%(���H����pm�2�n
L	�&�存◕w �J'��"�P��5��p��e��pdv����;F�fM��ڹ�-e_����Gin���-,��-M݂&&R��Vd�{K	����ԓw.%7�cqɸ�;1ݑ�Pà�#T+).�mn���N Wb��o#��wXR��m��i,�YDr���=��{���V!���e^o'�i.*^��!�WrK�����ի�Tc���eɡ�v��9�N3��LT���4B�{�nø�U�x��D2�Q�ţ)e�ȍރ���B�[��eXgq����ZG(qj��� �k1?��G��<43~�n���g���%�.�������ѽ̉ɶ����ks)����0��.����	4�}י���Kf���40.��L"6��tZ\^��*�v��و���2��b&:��&�8��En\��R圹��x�փɺhą/L�J��f��_u��*�|��M�}�r�3�`�dZ���L3t�"��@�$�1�^j�����e�J�Ah��Z2�Ep����i�|-��R��'�IV�{�u�eG�n��AQ��[YE��eZGs���0Ib�ݩ�a�hcDP�ۡ�:�U��Ku�1a�f��B��[1��݃l*{�u�c��V@6/��][G2��7Mk�u��-baݍ:77"pJw35-�G��@�O5:��w�b�ߦە*��j�Ѕ��V]jĮ�RF�E��4;�%�WZi%1�]���e^�$�)�`��Q�7��{u���X����C-`�hbiպ�;X"�H'`f�R��u�bz�r��jz���Ud��m&�mgQ� ��W� FزQ=X-��0�z���:��f����\s�!u�P4v�\tYx�V3���na�ei�e����RmP�U�GB�{.܊[�WY0��K8��k,�
��Pr�CE���lt���P�T��SQ@�k�_�ɣ!)���Y��ע�	:0��
�]�cH3)i��{L�b���2���D�ލ�$խ�`M�I�g^a{�Q�3�/on���)M���찯�ZK�Iܾ&�,:�VkWW��Q��g:�Jm�l�*�{iVP���*��P�p�w�d���G�[ob�X�,�~�Z:4�Ѻ6�!��V�����4�%�"�LVee�ܠ��NX9�ہ:�.��s�X��Is[}�r!����&�[Юm)�
F���	�*(mF�4Z8.ai����A��SH����,�l������X��ߥ�h���tņ��R���;�2��ܠ�g �TtY˳kws���iu$7r���A���L�3m�B�U�aٹW��3P�X�
6� �7��Y5�n�ƥ�D��W���q�˴��(Vณ`�1�q]�z2�S��fAB��h�Y��)j[��#��{Kf����X�,;n�CM����(Uw&�]�\ӣm��j�.ݝ����a�4;
�[V-Y����;��.l���wܒ���j��?������KM�c&]�Ј��7*G�f����4�B�d�����3E��^�cѐ�����v����;h���;�+�/t��,VE��ѾdQ�
�`�
�oB��Ò�-n��r�Ia�Bj�vަ,�y���6d�h2�F��˛�]�[�%ܖ����N�9���
��Ε�VIe������:_;*m���'E_r�lLT�CRV��+�Ս�Tc�WtU@^�q�Y��Ċ1Z���4�)Cjΰ�fw*�CEt#�.�,�[�3d�����]�曢�:
�8���c�i��U\[��KD�˸�c6�ݡ�+^���njՔ���n�.��t�FL���=���ۚs��S�H�5ڧ'e�3V�T�w�F�㊌ڎ�y.��FCy������f���2��S����N��F]նl4��E��9�GJ���
ʺ�_c`ؘ�#n��G(H���3Մ<W@f���gy��]Y�]�Q�C;dѕ�&�r��j���Afu�=���`�Q�D��1]e�{o�^�	#�d�S�!�4��=�4Bj;��V�-Ζ*@����c�fa���<�C�|�����zCa��L�.�>]dķ�s���T�3���**���k:�<��wmC�u�]o3��j��Q;
�k)\�[��A�9l޻�+�|��<ܥ}��	XCN��w+��}�i�V�Vfˮ�&K�),�L�ji�ά���3H�t�u�gy	`(P��u�[AEv��Lu�������]3rA�D��5]��ݐ��EP��G�\���+�L��̙�C�R`����F �In�2�J��r'!a�Obщ`����j��'N�\�4e�M��!�9��94k�2�m3)�A��x�n�7�kZ���EQØ`(�� .QKyZ���4��Wy�e��\ۢ����ᎊ�f�)X�r�n�[�,q�~�*!�:�i%�.����+�|i��W2E�����%	�_:����E�ܐ�U 8N�]U��#�8a�b��F���[>�YYBI�D���AxխB��V�T�`{7u�W�����O��
b��(��Jq���QQ�"[��̥;/��0�Q0s0����5��RW+��S�f��o�V��ŷc-&�ˤ�9P�Q-�Rn�a,}x���얐k܎����P;A�"�YPeLV �|�� y�6��	:��8�U�k�jdx ���;�/h������p�;/�2Ci[�]�Tc8���Rj����Y%��.�+T� y[|��0f���L�'F�gb�x��e�FJ�G!���uuOz�@���3W���mY3�a��ֱ��*�9�h�jg&�ƚA�j$��c�䩗-S�yaa�H�ep�e-"�`j6ۙR[���3E�M��q姶ڹ`�s��b�o��X�(ZZ�CU��r�<Q��˭6�t��a�'w�uk}��t�X2��؎�
�h\���G�졒�r\���@]M�[ȺF�,�7dͰ�⼂�<[�����8���4�<��Ge�ʮ�&��h*��7���u�;ޢ�R �琁{�k���H�W�Jھ�����ޓ�A*���1]T�r�9�j�s�o!�Ѱ:­��3V��6mX�:�޺����}��9�a��Zfz�h����]��`tn�]9�[�.���6���$�x��-��rfw�&-�]�4���SE��qe�IGA�zWQQת�om�e,.P_Kx9��kn͵�%b�+H_ג	yL�1HP�Xv�X�>�jM	^�N��xP��|��c.���c���$��(�͛�,�Oe�	`�.3T]2ZO�{_k�%�̷��JÁ]��5kk5@R��&oj��1i�x2M�a��,�,걜.gTc�;�!Ԯ�� 8�$����v#�;9��Hlu�9Q�E�8���դ4k�ӵ�{`
]Iv�J��T��j�\�5�f��j�Æ��m���h�V���+�&)Eom���*�]��o(�E�Up��S��{f� ���w�SV�gj�HM��I.em:�E�$MX���0�9μ���{���d)p�J�8bE�"�|-g)n4����K��i���w���s������b�]��d�d}�a�o��ʱM�71t��쮫�D�F�];�e����K�R�� ����0;�-f�5V��MX��%TVv�6�1Z��edq�~G;,f:ѭ57��R�npEvԼk�����E�$V6�ib�k�uJ�+;��n�zZ3_2Ktho�5ȱ}W\���R��;x9���D��܆5B��YY�]�ǃ��d��o��(Su{!�u(�����W��uu�^v�|l�_m)��Tn�V��Anu��pM�'`�=��r�t0TL\y��js��tx����Y�;�]DX��?vU�T$��Ɂ���v@K��e�5����\wZ�X��T�%v#�&[]��*WV�>]f��QY�1<R��YH0�y`�����n�5�x��d��tՉ���9$%u�y+]�	������S�,��dUĀ�$�,^�˕��:�]7��k�Cg%��*^,>��^��qܺV)s>�t\j�K'�^�;��lE[�cv��.�i\$Bң˲7�p����h�V��*��k"�AV���Yˬ���oYt�L��o�gڑ�d%c�"�{\��a38�xt,�����L�(-N��5�V��r�;"[B1�bEJ6��{�#Hs�Ysr��8En5Y�t�i=�C��f�j�Jf��X]��C+Q�kkM�% )�m�E�gS���C{��>J���Co��R�2Zٝhd�h�r�LQ�w���F���J�q9qq���t����D�R�!ً��S>]j�B�Lv�G]���2���\��'��pδS9�-����ML#yQ����U���p���s4%x�]%	p�x�!��ԨgP0%+Q��n(�o�kҋvrK�𪷠g*4�iL+�sz�P�:�-����0�\�#.�p�f�Ի{ۖ�'��B��]`�ُjݾ%�q��4r���j���Xn�'�8,r��� ��t�i��q,]��:��u��qgr�5j�1�����*9kv3ZJ�d��啛�~�Y�չ��Dル�2o Gwm0�A��r��l���yO�oN�)qP�N/�h]�\����%���e���r�A���S�|��ȣ	ż#B��LT3D{Vv��5x6�X�U��fгl>Ks`���8�
nos����iO����(nj�g�`^���uc�T�Es�h&o�b���8ܓ�w�q��6+Y��$�Ӭ��
��Q�X�ts@ us't(��4�8�e*
��S���ZdPۣ��p�a<\,�̘V��Yc�ܓ6-4�2������
:trY�t�VNP���K���g��)]C�2��}��nVf8N���o;.��w^�D��T���[ǁ`�����.���ǅ�G��dutl�N�pSJpLq[2VC+�:~���S��,�՗kGR$��:c� �D�+��6լ�Г��T����Y=�FM�J+.JUΆ`�2���	����*q,*�=�P*B�jR�8B.#y[�l���Ie��V&e�z�d40�k�wI��;I�D�{n̽���lN��6�-Xy^R���Y�g�g9��5���rh�ި�PM��Fwg^5�jv�Y�\�c�ҥs�h�o!'��۳7��p��Ҏ,{KS���f�����n�ZQ5������S��%[�}�h&n�47"�X���q��4��u�!Z*ټ+�dT�C�����ܧ��H%Bħ����)��W���q��]�+9�Ry��[�;:�ܛXp��]��pU���v��3L��w$�o{���E�Y\�X'6� �"�6t�.[�b���\Iu�b�.�⬄m�5i�S��B53�ͤV��%���jw��ɂ�V64Ea@ΔNջg�<3@I
�D�[���ڴ4sA�8��B����Q�V�ܳo/l�����J��|�F�r%������>�v��z��3jj.����P��'�:u��Mb�-�6����b`jʷc��;v�N���[���&F� �N7�Yg(��h���6M�{FX��	��@L�#�KRV���1c�[0Q�U�I���;ej�&�,k��4��6C<�uܻON���Q���V��.J�oT��%��Wf
��Xf�t:�J椾d��'��:���3���\Ќ�t��zW��sJ讔���Z
����8�M`�a�}�j[إ˸��)�B�'GP�8xЍ���(Щ�W<�hz�ٕ)]��W�3�I�6N\��|q�$��y��b�r;7&�ׅv��KUBeܝׇҼ��t�3B��&g]t�[y�H;��޺HΜ����7ym��6e���r���*�����Pe�So5����|�;�&��+h�g1�f���Tj��ƲS�u��qi��?��ŗ��]u�N9l&��ƥ�˫�T��h������U��A��wX4�fU�0򭙫c;�`�]�s�tr_FuɎ-�fB�wV)�V�4úow@ɍ�����JZ�t%��T��5^��r���:�܋��!���ae�cjG��M.����iyz�	o��yK�*�B)�}�:_���Y�yS4�%ٷ��n4��)uvVO�K����w�5�nIūj�����A�i��k��a����4m+Xx[7Z�U�so��s��������R5�u�k�0b�Ӄ��Y�)��e,�]/�%t�$.:[dcb��:Α��M_Z�Q��WYG�3��>~�a��N�A^���x�0��ӂ�Ф�Q,��w�Zwk�{��ul�ʬ��/�Ks���In;F�n���4����۫��Juu�b:��H����]��@�R���غ;µ��u�6�4:��yA�	���%��!LW�*�D�X#h�;��T��%�:g'<c{T}j�d��`����cq�Zt̠�ZU�flۭw�z�*Z�ND�q�Q���|r6:��7�7��nY�'��1웩�\��)�v*�o��dOx� J��;-��`���[���������X߸���cr=����n������S7��^��ז1=��f9Z0�+��b��-�4ۈ�(V�<��e<O@ٝڻ����.�qܙ�����KW��G��+��n\L�K-D`'&Eׁu�u<�2���A+�]��v��/��9$9�ɮ�fq�x�6M�@�!/�s���v���j��w�"D^��f`ѽ�2�f�T���m	���5|�m��,<��K���tաG�ek�k27�3��+����Wi�q��ɨ�!B���{�8Ḟ�W^�.��+��9�۰ʾ��"&�Owq4�%�-q����z�ʛ�#)���)��{��yLV��ؙ�Hl��*�/Ee�VsR(�6�t��հk��a�SM����wF!���"�Y}���`"�p9�3�2����<�
V�بn���Y�.; u^��`SgU��t޻�Y)4�]G�+)5|�Ǥ�#F��y np0��#���-��6=�#�����Z�s�Ftn��Wqh5h��n-��\������冇�ي弬nl}g"E!��ܨz��u)\��V�V��hV0��7{ImH���:�C�����8Гr`Fg,fV�W-:��0�\�R��"$���S��D�Wr-�:�l^˔�󓅭ysZxq݂P�9Z�X$�8�r��e �J;(޾�����_b]�1.o_.���:Ko"9֬�	���qդ�f���h5�z�r+:�J����K�=p�3FǪ�p�WAK%�і�=�+k�r'���#ơi+d6.���m������-���{�^ګ�le�){���`�����<��U�̥��ʠ8|��\��r�ְ�z�`��u��.��l� �q��4��5�3ݑy,�P��ov��SN�6+`X������X�P�	Pa\��4[����o6�����1S(�M�����ќE��:/k�	|�P�ґB��V���Z{�^Wj���U�%�5��^��2m�q%,�E��<���f�nH�D�%�N���u�u ,<���5���q8�Z����ٴF��4��V4\9�oV*�����He�"dT{�]ġچ�����*�\q���f��Ԯ�&���=:��;c�H�-.�mWb��eR��no	�v*
��#���cQu�>�10�;M�BV���y�h ys;�&q���ΫqP�����6)�1�gr�K&r�T4�������i��J��.
�d�&͸�!h-lv\�nN�J�/X�W��$�b�P6)�r�����E�Ik�֯�#,:;�c9�� s�J\��Rt���{ r�#7{:�T/\�R�OiW�Z�U�WV�,�������k+9��h����\T���|�5�oSML�۹�Y[�(l�([��=Wֶj��:&�)�ܧӠȵ���G1��0�0�F�TG\[�e�C� k���N��S�L}u�cO���Z��޻�1uv��ӓ+�/�����^]���x��AgKoIh�]`"���݌�νe�a�6WJ��a�N��^���W�i<^f�GԖM�@�MaH�wJ����"�7f �Gh�|A��&{9��Ƴvmh�H"/6)7;n����lJ6��[ $�d�W�YK{�V�R��s�(}�26*22�s�� .�U�(��ìf�ʾ"@��W��]'o7�5R���\bD8�-h�Z�Td�s�p;ك����Q��wq�&	*��9]b����.]�yt�"�
��e4Y"�,L�t��hc<u���
e*)9�|������y�-�j!�7��i"�t��J�irz��9҅�E�c�N��]�óg��5�Yz��xsJP�&�$�ֆ��3Y�D&��`����Vf�o�9��q���i1|XC�\e]�_TU�[�f�
�%H�IN��EY�kJ�,F��P�ľGUv�v��n�7��'1'ffj�J������	��<��b�7�J��άj���������}_}_���ﾪ����uÅ`�-�6'7	p�sE�+u�[u�;22��4F�i�[4�We��$C/3 ɕ�n�[Oh���Zs2=��y���ǵͫ�f�q� K�k.\UN�ۅ�C���k�7v�p��F�l��P�	�b�K���q��Z����#2޾AY�C���{�5��o5w��xZA�� n�*��O��F��@�$p�y{�g>�!����j��٪	j�.��#���s�QLwr3l�+�vU���et�U���2�����PƂ;t� `�$ђ��$���(|��w��EZ�:�7�jbt5�\&��Zо�
*�au���3�Vdw�E,��A!��K��y�456R[��˶��ջ�RTe;�u�)Q����l���
�����d12Ei�]b�O6��y{ג�G���ֳ#"d+�v�M�t�u�#ǷK%Y/P�,1:p�@���R��nH�� k��p��ayR�EE�*(X�b���87_SJV�$���9AI�y���fH
B.z:�*O���	l���ʽDgHs�v�k��2�[�]��b�=<�+ѡ�[(u��"��$�4�����Q�5����M�9���g��G3#���[�r�1q���koU�R:���,sE+���`�zl����]��!\5�,�*��&V	Y�$t`Ev��90F1�:���ҍ��)���Щ����Fӂ�)�k�B]=�+-���TUub�%elZ.��N���+-gșz��I�{�� =���.*�4�j��Y��ފXY�E�'��N���-[�7�^��>3�јL��J�	д�X��e)x�cWn��Ե�/:�%�°�$��NeԘ�ٵ2�'O7-����$	�W{.�<�����*��	gw(��4�hz�t�҉��賍�-|�4͢��rXj�|j4
٭m�srM7|2�w4xQb�L���*!X�v=�s��2���-v_C������cɗr�����]��dзp�L�" I[�'v�1Z�@���ndj�3����%8T�gI�YB�=u|iBؽhoU[J����u�4��CM�
l��W!:�	vк���mKOV��j�6^��*e��o�Ɇ��BR��c�dϟN.+�:�1�U���du|B��j)iŗ�pK;Y��yY9��p��*���yX��Pҍ��qN0�L�9(�u��Ne*��yp:��g_V�K���w�f�肑��)�HX�CR�����na�g=�������,�r��+GB������]�&���PX�n
�xprF�HV�$cI����g��e�  a��0��;��Q�hi��V1җ�J���E���US�%��0�B��lr�Y�6���)]��W��k��a��J�WǱ�}Ք)��R���Z�^;�2�eO(vϭTR���"E�/5Tm`�Zh-��t����v�צ��b��/p�t~�o�Z\�%�CV�}�y�n�^�� �jZ��7�޻��-�.�-�1ƚ�摇p�*@�4�����]\�R���7���v1l�v̓:�ʻjq�w�]RѼ�b���Y�.v�A����v\Pd�KKM�p���	�*�kZd][�I�o��#��L#��ݶL�HJ˶5�@�q��B�k�k�[܍��)
�W%���5�E�ј�;�_A9��bߟbvo��31-P3]�f��3f�⅕u�NE0����NWE��e��#G<�Ӽ�_[��(���2w�lY�3�����R����+�g]wQ�o����ihKSo�ה�6v�Vd��ȥ3�N�na[��v���������`sIG&Pyy1���ڶ/IB�t�"5���ڻ��J�E�,@*U�|̥�8���H5�W[)uQ�D��(��d���zM�������#p�̦��@u2.]�uۖRĝ�r�"�dV����ӴַIY���ub�����5�|mS���tJ��i9��f?��[ʰ�E�P���U�oeN8�����b+b4b��R�Jw�Gt��uh����ҕD.Y�\��)Qi�Ô���"�S��ј����%e�\�vb���o���ᇨ�B��+n��s(�/��)�d0�*�X���6�d��t�Ό�#�H6)	]Ǫ���ط�_Q޸��1�A��
��b۠OuҠ�|��ЇWSX���8x�B����4�iE��GL�J������+�f��gu����r\_%&���Rj�f�1�p�yG���ow@(+,�}O�����z��ٔ���wn�2O:��l�)`�:U��WT�V�H�u��9�oݬ4_noCJ��j43�yg�`�C6�f�դ$�}R)���l!�$���D�1lu|� ���Y�u��{�F�[�Ǒ��q�����g׆خg(S�@��s�3�5��!Vl�4�sjS4DCd��U�Hn\�I�F�
54�U�Lܺ��kt��G	&^l�սv����eV�5�]��7� ��㛣��_XI����VMN�^7�u�ա�VS*D�㸯P�Zq�9�����d��I�Tju�*�@G]eVČiE�z��n�C45Rݾ�*���D���f�'�����hPc���3b�z�b��|�a\��@"<�\��e���S�z�h��/E�RV!�8h���G�g{����t�HΈY�}s����'Z�@f��V^5����C���W�]��oA����	�MJڝ}l ��B�����zbY�q:�޵��/�L�e3����/�pZƩ`�)��<Y�`�XV��	8��L(a�e��ör����X�'��sL]v�1<۾�]l^%G�O�G���L$����(�7J���چ *�ky���=�y��K�k���m�Ğ4IT;8h�/ƪ�J���u{e��8ydw��o�+��Mb��l���F�%]�m��ZΉ]5Z�%]�î��X�_U�]����'+kf�kG����Jd�/�T��D���0�a�Y�7�'��6���Χ����o��d6N�Xd}u*:	j�Y��fSK��@uZ���O�Bv��w��Q�͵ň�;�1l��\vkN�Gj4`mm�\����7I]DԮ�Bb�]�q�5z���q)�&�oU�/QӓD사lp|���u�؝6�3���v���kˇ�^z��f$�̤�b�V��ԉ�O�f)��6��㝦�3.�]5ʂ�:�uj���c]�n�i��kLJKT�n˗:<Iu��iМ�Els
�7�v��^νp> �ϋ����v�Lwˈ*������{���zȘб�јM��6e �!z���!����#`CKP��M��s yoGi����2���ɭ��`8���ʽ^�[6�2,��K6m��ݔ�$��f�ź�X�AlY��ԉ����7���	,ˑb.�A�T�_K�=�Q�x8�Y�r"��{�I�JJM�V�I���%�����_as�q�znt@ҙ.f�7{t{��]8�b��A/,�����ʕ**��b�AM�Ƥb�VL��{"N��Z�aWQ��Jj�ܬN$�	m:��'���E]LR/�fh�;���6�fDw��]�n��f�ޙ(�a�C �f���T}Kg�����AE;ý7�v�<1^j(:�u<\�-�y��*XV����7X���̎��m�ŉ�"n��:&,��9\�U#Ӷ��o��y`V�+���f'�7A|ڙj�\q֞8��r+�Ӽ� t�<��	�<�g�,��j:���|J��0Ӡ�h$?�����[9P7�KͶp�1�V���m
-�fdԅơ�ڥԥ���[t eju�vk�sG�	�Q�&�;B��\��Է:�n^���K�\t��;��(�ŉv�+t�ʹ]e"ﺑ��m�kѠ�E4�}������$hq4��:2� Q��c7�P����@q"�m`�T4�Γ�p�(�I���hi�s�
�M��Ӯ��7�wZ�{c� �8�+��9<<�hU�6��RIefN���K��0���[A%��9�I�;�D�gM)V�k�?Qh화�����m1
ͨ
�Ժ�
�p��/5�Z�򮙆�co�)��1�^un�T
�0vWnr!5El��0�������Շ�:-][�f)y7d���e�v�HV�|{�t�\����祺�X4�.&��/��0U���ů.�����j�=�{�1���lA+�*g�J�.f��Y\f^�]�2�b����H��+F�g�s*m�p#`Wjs߳;��A�4d;�n�J��&������Z���2��S�Jgt��-�v����ޤA9}�/���c�j$�yt�]As7ʺ�EM��J��9�@��˄h5�t)�7��Z�ذv��-�;����kS�wG1
ԧ�q�w>���</i�ز2��㗴��\�M/+Oi�K]A��(��.<�'L�5�]nՙ�m���pd<d!��=����4hV �\����v����t���I�9c(�]��H�Ywf��]ƻmS��m1=��j)d]L��[��[��OU����/,!\sIy��~k�/��+��H[cj03����yq�.l�׽�i޻��&�fl �N )�Zy�(Y��v��˓!��V�4�`"՘���X;��h��E9�:���56�t*7fP��˔[���=����m66�V�%�y��@y�6�П�sI���s��V��c\Ġ&�M��{x�&l�Η�\��v���*��R�R�,T��ڔlt� VjF��W��؃;r^G��*�YV�4�����I������hp�p9�![�i)���>�k��a����A�FJ5���������w�r�tmTJK�}�����Ao��ΐ(^ލ���t�A�����&nb$����]%B5{[����]�KF�W��a=W.�+@ki۽B���-���4a���)�|8�f�d�!Kx���Z8��v�Y�1' 0T=ո*�Jݪb�,e\�n��ُ�VJ��A�/��h���I�A.�6ns�b�_r4n#K����kDN�@�c7mk���s�Պ_!���L�D""!a:]�Խ�g�a�S2�[�B�.G��E:=H�R��NR�ڸ�-b�d�m���_��-��t�����jȢ�M"�H&R�A�q��^Fu�|9n_O���=��Mc趉�b�
U��W�����I-��(.�h˅�c*źvT�V2�!O���X�R*�VjgQz�*�[�u�� ��[�	�.�'�۳C�SW�e�;Mu��u�Zyҁ��7�e'��}����I�]�:܍]��F�M٭��p)asҴ��GoF�:�
�Y1�,Vn�E��2�V���mӥ,D�/sj���ZR7q��(2n�e%� �f��s�m:��1��<j]4�	j[\U�]9�K�W�<�ه�����3���X����CF�%B�V7����ȶWR��	�u�]p^Gh̅c��*f�WZkU�+>���C�xp��w,��3�։0�-�^��.�L%r��;��]n[���N�z��ѝ
��/Z��ů�e8�u�z�-sMԫ�{]z�K��𕚨3I���v����.E�u8];U�J�YS��������:��\��{{2hmS��O�X����Đ�ɔz*&�v�(֜m|3k#4E`��S&U�;k*��[YpZӊ��Đ��jXK�,��k�d��vP}���/54_T�Fv
�pQ�FQu8�s4��}F��o��Y�,ɩ�A�'+pW=�{:�=��n�s�X@k�wjr�Gh݈�풉%������J�z/tiD��8�/8���5':J0;N��N��Z���Zr��mY��k
ֱ�r�';.guWRŕ�6�}��Y���gg�ԛB��#h&$;y�����u'm-÷q�ևgx�1Ű2�:�;0é��Y�J��DI{��Ojؖ��I���O`Z�L)}���݃�]����D3tTR"5���m��W��k���ea]7H(LY�uցn8X�s��b���b��ݛ���g��ۂ� �mf�E.�&gH�<`���Z�,�R�4b�N�C7T^�p;N�f��(ZY��q��Au.���CsS�ZL�dCq�X��x��Q;�&k5�70
��er�_X.)n�P.�يtܥO��v3Y����ӥz��iS
4xQ�J]h�	����)��M���m�&򍰩�·�W���ق�<�c�짏B
�v-[ԲR���)�eIJ�̓B��� Ef��[vN�2�&��o�)�:V��}��r�>ʹ�$wgھ�@2�R�ćs�;��4�[Xf�r��J9F�?��Lvh���\C\��V�Rv�C�u'��[z	ܱ��I�A���;&��".���>�o3Y��G#]|QuZ�;lu�����̖h'h+kO6Fc�Wms4�PR�6�%���&\� *��f�h*7u�%��e��8^�|��u�p�EZV��@qJ�$wP�bX�%ۭ�_v�m��(�_Tʗ���p ]�=��-:����7Z<Wh�u|6ɭ�����:M�U��g��ud��g$����:d�&�q5-�m�V���!FV۹Be�}FgQ����5�f�ko]�f������k�]v<=CAw'f�QnBL�g��y��;��w&t��� �Q��:�8���ゐ�SV�P���s��Y|��DZZ��v'��__ٸ��[��G\��Ҩ�fS)�u�p��u���9�sS�I,��%��nh���ɦ�3����F���0;�5nѰn�C��3n��naRWd��;}`�ʝ��+���H*�8z��Z䷮�3��T�`Ei㢂���t��it�XGi�\N^fM�i'[t0�4pR:I԰��g����諭���>��f�>��ײ����Z�-R$6�W������Ҳ@��ʺnVM��ʋZT���94x�,���NY�ό�TӬ�+�c�:���x2�ъ�qy[�1E��\EHoȣ32}9�x>�ѐ�-�S�\�퐵���`����9�qِf)d�&.�2��,nF��Ƃ������T��Y7Xݠ��Kn�U���B��U���Р^(лq�]
��u&8�֫V�o�n�J�ԥ�n��	��P5ذb���
�����W{Jw�l��[�$�e���YH�����@nia��7.�`�b����F:�{XX�R��"�d��[V֮roE��q\��c�p�0"f���y��f�@�B�,[�����R��t�"�,Z��-���[R%���-���c��1���7@u@f\��b�:�35>I{{aV_GAn��
�|�Z2b9I$v�����m�D��jY\4t(�=�5W5�Q���^e�e�!ʜ8�G#|��� �uץ�ʮ�n�3gPW�wQ�Ź׸�7ʹ�U�5�D��w�a��9�2y���Z��C��P�2Bg��;���;����x�7.-V�kK�r�� @ll�{(�ZZQ���)��VV�C�>ͱ���݁���KeuJ�(͏U%]�X��b���ӆ�E��Uָ�y�9ve�����y��Gy��Ν#Ӵf���/���Pch  #�T(|+�~$@RR��0�L�	ss�5�	��A!��K�mP	�RA�6���(/16Ѧ���cM�i�4�e٦K�d�戈��ђ�D�9� F�R&� H����H3$ ������%��"�e�ns��$!"$N!&6��#,�y�DD�� $Sk�]bTGNE��6Т$)HHB"�D*P��H�3M���sj�5�"���"�s���ⓑY�i��.�\8�9��vh�iƈTQ"�8�"!�)Dd�(�b�3Ui6�"投��� ,B-�4�]�@�́f�"&/d"*��� @����Eڒ��E�����$)B�46��Ͷ�FM�$3Uɳ!I�m�X�i�$
�d$C�B�H�w�`��5�/���<8�h_Y�Y�^�I�Zl��9��}E*��g%	`t����]�+d+-0f�w�ƺ�<kLn���"�Ì%P"a��Wgi���e��N-����{ۻ�ǻ	mԛG.z;^Q����ՀiM����2:Y=�"f����+#�A]}��.ڲ{a2z���lF]賂5[���0<��c�uS�v4u�{_�P#k������N>��ޭ���-�j_z��X��z���"����mT~5���m.o� ��FN���W��[��n5Z�?8��	�ݮ�Z�a̪�!|�u����w=�*W���WiF�z�Nxp�j��v�C�X���7�N�X����V���
ӿ���3���ð�����;ܳ�sI�Y9����vp���?X�tB�ECw'[&�5Z$��RcU�>�~J��\s^�f��*E�UV����kHfZ��-�/��kп���B��mNc��gC��ڞ0�GW/N�s�d����b�cs'GP8LLq@��2��ʻ\k��qP�2�,��}5�z%]�F	m����!��G�g|������ x"x"�)���d���t����b>?+��i3^g��A[�h�V"W69e��k�PN],��4�XMXT��ա�[R�܇?M�a$۠�a8x ��R�Ϋ׹	hG�J�u+�Y{J�(X�^K���@��۵6d�\폤��
i�i�	a����!fkO���v�����|>�On��_MC�8`��z�#��i��{aT*J5�@��N��XU��v=	�W�8f�+�9/���S�*��>���p챩��/D�@�~H�[��i\�7t�t���M}^"��ABiU/s���*��Q��\��T�jx�a���iF[��%����O$�w]͆��
S4߸���.��n�]�\���zW"�DQ<Gc�����軖��`�x� �\,����~T���{^�O#��h���!�]{h�O�13w�H�e���M܁�T+�1D�لvF���ja�.����y+��&�ߣ�z�Wua�b�9���^\,I����%����{V�c�gb��U^�Fi����8���?Gq*w��u��eZ�K��~��B�#�r����ub�����%���TA�ռ'��$��3��9�:�;M@,�9q�hW����e�fs�똭�����37��N��۩�O�
A��s=ET��s��+U��$���5��jB-� ����'�2�[u[`�YV=�[���#ى���ʙI붶}yES\� {��@N�9���Vm5v�z����K{}#��qT�[��٧YY�Li0>�lY2�K�Z�Z>`FWG]N�4�dU�N�T��3$
�^M�{W�3�b�rq����9j��%���z�S��f���[Z<ivV���q�qU{��^����[Ԙf�q͋�����ҝ&ImOq}�/�:�/�n��{7'ũ$��<	�
I}1���{��9�-k�9�	�����J��/�'-��Sw���<4Q�)� 뢸�Q�=J-�.���5ka��=9k(�j�(M}��^�t�d;Pڸ}�q��P��	�C7����ͷf�m�s�D�̠$d����*�/���B�%�.9�4cYrW�@p�L��~Lk=%f͝jM�݄���P>�� �8�J�����VBϝ������;t=��+Ε�s�6��4���Q�Bj�SQ� ��}T$*���ǒ���5��\8��`��zcjeI�O�q�Dq�	�yX��@�8 �I\pԤo�`<"��qѷ��S��^DPޛ����$z��#).�F���i��*�*�$T#L���ck 4��yVIoq+��Vz,H��0�i�.:!��xT����f����k�1Q�F˳$�Oi��1ާr���1
�z�X4����`��a@]a%��փ:yg
����HЖ��\��:��ҢW)Qǿ
LZ�MĬQ|����PҦ܏�4���;J ��Qbz����Vʖ�]}\�>�3oJ�+��O(��'7Jd���A9�[��XdV�d�g���څ�!$��\"�s5�r��Q�p|i?n��;��O�~0��ܱ��Tg�OΗ,�n.�I~,c��u<߅Z�A��Vl"nf.�-kD�A��9����`��|���;��b��J�VO'��q�ׄR�&R~z�5_4_�T�Q�%�_>7��r��s�¹�/��`vG���Zn�{ģu�;N�ˊ*/RZtt�>x�;M&Y;��ɪ�w�������G����ѧWG
�r������<$�E4%��q��,�l���`�������8��Gt�'�����Ĳ�'�2������Ped@�V}���T[�LE�-��u��D�0�in8�YN�w$҉��Qib��f�upD�2���.�v2����e�:i�3Y��mw�'9�C�kD�h��x���O��k�=�H��w��Og�Ի:��+���7�qR$ƶ����T��U򯁢z�� >��(	�)�>Б]��o�*�D4�z�� F,�7�>�d�}�*+��+��~#����cT�Kp:�zj�}��0���@״�h���;�	����@r�d�Y��E+�>D���H�RX�#��3&lt��Y��a\�����j���7}(J�eQ{��F���r��j��(P���cw��䕦WEc8���c��@��;���2��t�a�`�&}f_q�M$&VË�����d��!|\-�����m��&��p��ۘ��uLȯ��F�T��.��kv�Rw�Z�qi��I$��BuL!�K�s�����
j�0"WC5�O�f�fb���3Ʊ]$�Y�%�Oa���I���\b�z�o����j�/>X��<"�+Q���ν��޷DR�I�
M�}��E�V��ѻp�V���6���P&��4��ۇ�KU�I��@�����K'�X� hvm���ߊ�ǠRe+�t�1����FY�=i��M�ݪ��\������z�Z{�\*���/��+�0�Ί�%�÷��E]nV���-��u�B���/�n+�Z��O\mFiB(:1bp���{j���rͮ���?TI���l�:���2R�b�gy�M�����q[� �9ڱ�L1��fbĈ�xTU�a��@1c{�dd+N�e3����V�]��2�,���=�i��}�.+\�n���YA���ɐ�����E]���*��qn(
^6N8�g����V��]�����wJ�[�aN����K���;�3)�[��i"G��!�{qq��QPn�g1a��I%�r�<�G���.V�Tmq<T2r\�O+�zv�����|o WP�C׌������ vb���B��DУ`�Y���U�wK�Y��qc�M��]Z�'KFx���+��@A&��^h��ꊎ U��{�f�(������6b�Z�7"r�t
&/����P�adT�0Ů���Ti�6��9�(�g	�I[�̆^�~Cju� R+A�x�t ���U��b�iX��6/��i��?b��yۯ������i�#O_�q������RQX=�i(���DOf��[w��]�)�EA�iN���Z놌���{,nD�l��� ��ݘ�v����jE��M#��Ɔ_B(o:���T�8͸�nQ��]pMR�H�(B�0T�����у	p��ۨ����$p,�����9�z����b��Λ7y*+������OTL���[� �*��Tx�1|�k�ѩ�wٕ�Q�>�3����	m�=<�����Uا�f��0'���èi�V�����u���On߸ֱ�.i0�}G�ٝ����-�j������n�Y��WQ-��w\6�Q}�g�^r��g�l?�V������+��WU�����!Y3�%�����[OW\�����-P%8ʬ\;6Ժ�a7B���2�f��$��-&c�a=;�T�=��+E��zj^\$�V�O��&�J�:�e�Q� �Q�M��)��E�q����ʖ��ì�․��@����:}���ad>���c�+[��J ���?)��,c�^q�XaeL=5�(�9q�hW���FY�g!:�c,=�x�`M\��]��t��9 ����iܲ^x�T=7�E+U���:.響�[�I�����b�Ǻ&�G��ڮq�+�q�1!���eaf;"�R3�!�����U�w\�J7"�%ռU@�N&���/�!���fo�@��Z8.�i|La-��o�t*���S�r��',���F��鱥�����9l������1zf8���l�c����n�[)T43x"�~���@?��*"g+x���E�F$Njv��������j��A�f!3�{�ՆW{�=	̈́U�x�LQP
.����+�.���.\����F1�g;6��Odrӧ'NLC���aW�57���}���U��1̬������\D�q�[��:ncoU���V�Sw_G�Ŵ�Zۛ�w4�.��;V�!�"� �rk!��+)�~�RkH�����-b�$Ve��7#������ �jJ̆����Rĵ\���R�Vm���@$�},��F/_\�z\U�[C/0����$���.p���zx���ق1̡9�*k�� F$1�h1�qy�Ҧ�Gj�����Ԯ2���r���/+�mހ͈8�I\lԤl� �L����4��Ʌ��x�wU�ᱯ���c*#�[�p��b๶K�� FQ#>F�31�K�ΌڬPA�y���O{`�9Wm�;1�Eg���xys���I�杚7�s��*����0 5Zt��(��0<�?��� ���V�W���g�^�p7�-?�'�f��v���I���E�(�˧�����ɒ(���c@��Lct��-��^��q](C��4X��b�S{$>Cra��q��2��;��^�@�ey��E�6�;�ݵ��+�i<���L�i?ڴkޘ��[~��0$������߽�٪�(Yc��~"���x�,����K�-��Y�(���D�ؕ�ϕM&Y;(k=p����j`�u�R��+��j#�\�p�=�<��'�w�o��%�tֱ"ʣ��+�P�W9�X8�='�fo�ޣp-�q�G�x�"j���͓ʑ	�m�S8dx��k�pmCY�%�ԯ�t�>G�y��?X���_��p�Z^de��;�LdD�����Y(�Le�-C#��4'g�\�6�>����v''XL��YB\x���'��O���۽�RJG6��Na�ô�.f��X����+�iAN�o���7������*�:b-9l�S���c��1���m�ڣ:Ez�8�U���`�@�*>Ґ���G�r�T����F}��Lc��܊���tm�r݌ f?������O���@|aN�H���w��Og�q�&����1��lmmap��ko<��7^�������q =���cBEZ��:B79u\i�',�����qW2�q����#j;���2�F�w�]����H%Cɂ^�s�m]�|R���g[�òS��a7���\��m�N[�fB$�:��cn�W�'�Sb|���0^`i�s!�े9��W>��,������q
������Z��G��J��=�*"N�&l�1Y҃p�Y\�?TsT�e�WҲp�.	&�pw`�¾���xк� 
�\C�{���:�����P�r���=Q]��"].��N޾�R�.�ܰ4�G*Ň��=,���!z���Hb�0J;cRӯW�iV�E��up��1:g{�*t���Cʚ�6�q��Yƶ.�$�Żq��h�F�#Ȏgh��<�n]g,T�/�9a�q:u^1�$�p{�2C��r��+��(��Pkv�ujlw�>ۊV]�Zr��k�����M�K��(#%8!�n�.t�xh}��g�Y��*];ρ�l�ϥKl����(�I�+�ю)�q<{�e�u����<1q��s+a���ً҄P4z#J&0��%��LՄ��'�t� NO����D�9�(��k!�uJ�rq�������j�J��G<i]n)��>�0�􇄧iᶹ��X8��i��;�[�L�ո�c0��Vi��(k;F�{<�g�����b��������*'Es>
Oy��Q!�՞�D����&�j��>�l�8�^[�k=�xn,*�m�\I�D��+���5����e_m�+�{M�lgu/Ux34�i����1r�1����&8 Iܤ�=s��g�Ljy�͇�q\��qN`i���Bj#R��9�e��?!�8Բ��l1�S�w�v8�!qР�y��r�c�����h�x���N~�r��]�v9����)�!�PLW���k�w����� !Ivy���)���ڿ���7>L��U�-�X(�GE
��L�=\�/+	�B��_C	��ޑSky����[��n!�U�A�v�x_ʙ��:��hu#YN��(s:}��gQ\[l�9��o	[�h��>�۔R�ww�:��7ĉ�ue���y���a���zuZuv��m�,��ͥ-�iXNs������&��n;@����KGMV*���-iV[y�fK�1ObNv]oQ�̦�8� �I�(Y�:���].��_Q��E�/1�ggp�.7127Q�2ܤ��؄\u+2U�Ʈ�T��@��d��Bv�R��h�9���9��<Xa춐}k$v�#zX+tT��sh��rcVU�\z��8��'L�t:��Q>�z���J9ٱ=Um�y�r�]d�+�X��]����(��l���dsB��T7D��wW��q��Z������C�ѕ�!���ՐTCfCyf���Ct�YΥȁ[�� �%b]�s*�����Vi��ƪ8m#e,�f�q��B�k����p�Y����.�9"�n
Ҏ�-Q5%�N�~6�cy�mAYľ��xdZd]�a���UI:ŀ)��#��Iq�
eҸ.V�S��AtӸa�aqr�9t
��+��Aqm��I�*�Ψ�33�c�E
�D���gWV�GU���|�*u��
[0����;.A6.�In��Ө��5����Ժ��+ݾ���o^t��l�9�U�l�*7@�Ү���]VQn��?*bA���qCe��rʔ)��7yW7{]�[��ò���!}͑�*dH'`�=����
4��H$^�w�M�Y[����Vu��;�2�F�<wR�=����{׫�4�<	��2Hm�W��MN�
��Vr3%�4���2sVq$�\a�M�ȳ&��F� �ʽ+fH[}�5�OLC��49��F��N��B~�/s���~��u3;#r��Ԋ��.�(^*[)Ja�<��&�=[�f����]�rgcY�q�+	�v%׋�][+\U{9Q!�Dֻ��q��`�
�5����vT;N����1bN�z��R�iYΔH���]�5��@Pmcv��.�'؟�l՝C��JU*����q;4�y�(_!�i��sH��t^.���9QZԵr"�t�Q�k"�ySau>��嚚\a�L�̼���N	�����fV�����&����stUcΫ�@4&L�D]'s/�o/R��6e�L�
T�-_!Sw��	��#�!d߉�Z�Y��t�yE����45�C��	�ƕ]s�^��hU�]�����%Xd���c6Vn���4����ky��lS��v՛�T���䊰-\���2��GD�}��&�9�F�VD�7����`)��^vԝo�U�`➾����lQ�Z{f��c�m�
d>�p�G0�VT�t����;s5}yyx��x�cf�����R�������Aϵ��a�%k��F��ܱ��6�hUw�NNk��&F�f�*Q"!DH�L��D!��N!���g6,A�M �!	s$R)JUUK��L�Lȹ��d�PH��"9��\Bm1"B�fL�#�8�PA*"%m4,̨����*�D��8�R)Ƴ�Nk��i��̰$�*��t$H'3]�	�[9�'
Lm �	&6�Laq	m%�"慉�"mZ`Diq��XB�$Av�b$"�d�],�0���m�`L���tI�$$D��p�$�	���"B"��H*d�B6�jnfj�˄�"B��"""���dDB,TB�`UDh�P�H��M��L�LF�\��$ƳZ�6�E���-m64�W�
D��}@P�ҹk+e���5�@&K�1\P☦1c��8"���v�5X0��a��C|�|+�0��ބ�{��X���mI�������=Џ�^���,�N�5�=Iİ'W�g�'�8���Iͭ._^$�i���'ë:�����i{Iĝ~��O�w�_���$�,i��?w��$��>��ޭ��z>��Ul��u?4���k lR�'�5�{I�V�9����;_�v��O��,/I���/�),&B_<�q�'4���if^y�՝'�{N%���$�|Oq?$���ݥ�}���dd1Ϲ �ۅ�]ۧt�t�?i=���R����[߾���-��Ծ��_Re�w����9$��d�ךN����'������x�X׋r_����?,�Y3���$� H�Y�\S]�V'h�T�G�}^$�'iǳ�yd�}I�x�'�=��I�,>K�u'izI�N�����ԜN;[Ǿ�}N�e�>�y7������{���޷�ļ^���X�qo��;��_�DB`}1��+r���ln��X^�{>�^�佽�^�k������~�%��|���떗Ŀ\Y���~'ia|Y��=�|Y��'����ui	=N�q{����洹z}O��y'�տ�'�_��)#�@
�c��'�U�N\��swl ��w�B~Iı�O�=�t/�ܒx��i�o���'w�ܓĝ���pI�|I���{�s�K2��~�����>%��<��V���8�����'b�O��iب�b��v�U�.>�}��,�}��,�:K��I�y����Y�����rN���,�M��Y���c�>w�IOS��$�nrO���s_�?}���ęr������Y	}I���uo�a�}0Na����o��+�6Vٷ�|8��y���/�'=�}���;B�?��>'i:K�i~~�t����'ԟ~Nrt�ğ��OWĝ%����N��$�{�u�:�K�N'��n�I�>�>�!WAAy�O�zA(5[2�I-��G�\� `�>��?|�((�r�,o�N�O�u|[�I�4O�����{_�r����������ľ�K�&��:�N�Ŀ�/s�t�S������G��Q����ShNk��1�݃�i�B�v�$�y���֗/׳��x�o�{����{��_��O��,	���O���O�8�>��}Iп��~o��|[Ӌ��|�9/�:qo�e�.� ~�d<��_->0�eA��2E_�f#H���/r����X)���*iq�53*�-݂��2�'�f�R��i�٩ձ�2��ӥ;N�ī�ڧh+M^��&��R�@�
�ˏp�wWj����D`��u%.�nk�J�M��X�w��n(���LW՗�g��:�[��:K�w�'�{�^8��Ｗ��������;_V�k'��y�'�8���N>K缲t���8�'���OR|K	>���O�>�����ϺL����>��$�lS�1B�Xɪ���%�n_��'��_n��I>���N-����ߗ��:������I������-�$�g����%�����ia'�����OϾ����]�)!fT�>�-�uM�q�}迒q,'�m'i2_�'^iy旉8�z��k�I�e�gSs����%�M�X�}�|<�z �E��:hy-�'i�u�:�����/�?{����u���G�����n�]��g*�}�\�\K�=������x��ǉ:_���>ٴ���x��{�BHBOS��9�KkK����Ľ���q'��rR��[�4���7������w/�}�_�#�b��~�{E]��ۦFb�ǩ���ܳ~״�?����,��:K�&}[��߽K:Kę���u��~if^��擮��x�$���qrݴ�8�[OV䰓'�i:_�w4�7�I����q�'٦G�����ƹ��Ӷ]��D}���'�rL�����}��{x�Ĝ[���l�`}�8��`' �Q���G�|�oĿRe��{���K2^'W�:N���4��q�v���ǎ.L��nO�m�U�c=1W4�v���e�#�����׼�/��8��]�}߹d�}I��'���Rd�X_������_W��Y>_=�I$�}I�{���K�N'��坤�ɖd��zN�-�^$�ife�S�����TMk.:�g�� (����N��nI;�{��[�r��;��,�'?k~����������_����'|�̾��}��Ygk�q,;��'�=O�8�'|��K�HBO����^���i7|:��H��EJ���W��`�H���N'�&_�����ٷ�N���I�מi~$�X�N��~[ؿ�r����x���~���s�,�|I�V�<���,%�&|��z��|�K2��sޭ�[��/��:T�^���ZN��o�N�w��
����=�K��%�s�g��Nץ��O�x��q?,�6�N�����|�r}I�'�w֞�����'|���y��OS���߹>$��_�w��������ʪV?���g�~8�?�a�t��K�b��N����ٲM,�m�/�F4-�븥gVp/p��q�u��])V�[��F�[�Y[F\B�|n�ꔮŐ���DS��7���Cz���w)�;IdZ��2a���(o��5|ЃfP����el܂o�De���}�ԝ�[��'�^�e��$�}q߾�N���'��;N�t�>I���_�ğ�;�s�e����|���O��X_/z�/k����~I�\� >�G�"a�6�^���Z����rG� (k��}���|!%�P|[ļO���X?k~�?�r^�t�9�'�k?���[��i�:�x�~,��%�&��xmd�|^�I�sORu���|��w�f�;٣��*��пf�j5W��>��œ��\�~���Y��O��NHI�����<I�,{��󾺽��R���''ZY���o>���y'�>%�?'���Y����N$�%�;�����w��O�>�D���o�W���f�x�­jo�|�ߩ~��{��:B_�ݝn�V�������\�V����'I7�/ջi|y.��T���I���:K��'ջ�I��I;_՜O��'}r�L��8F|�?`�DH��>��5f�b�Iyw�k��}L�(�z Q���Y ħ��w�gI'���gsiε���}I�/zt��vYϺ����|s�/�7�z����$�?��{�k��s缰��k=Y��|������8��������?�+S����ʐ��0%���M�U�}_}Oo7I?�~N%�������/�8���Y�d�ϼԖ<����s��彤�&_��:Y�~~[ş$��&K�ow����I�����=��S��[��9��+Kig��A{�&�X���}�３��&�[�>y�>!/����:�|I��,���mg�K8���{��ŜN,���st��'6���Kk;��'K���/-�>y��,/=��>�g��9I?*Xg��#� �K������q/��rN����V|���v�d��߮>O~�~[�^�g��<�v��!/�֓���9�Y;��\�mo���q$��ݴ�$�x�K��%�翽��7�wP��|Tv�{�#��"G�>�:������Vq=�|��|O�a{Ns�Y��O�8�~����}K��}I��=�Y��d�����z��I�e�_��']���%�;�i���se��~�q2��~�nu���￾d3p��Y��Fn�: Q�0>`I�������t����Y��?��끰٨}:G��� o��~� �S�c5�'����$�yg=䓡g�L��}�;Ki����v�oN�;5�R|Q�e���8~�;GD5T�sxD��$���ع<���{n/J�/J�t� ��Z�p���kt.��`Z^�Ć);7m���_::��oNʱ��7�;�D>Rj!YY���� w��4�#�4(�^>#\�6�n�rܜ���#����z<~���y��i�:Kę$�9��o��{[�~���E��_���%�&�[�{��B_�������ԛ�,��9�=K���/�şӜ������<=���9�c�|��w���������8�X�^��qz_Β��'˵�:K��s���N%��\���{��'���[ך~[�{_���I�I�d�o���kŹ>p�/g��G�DsP##/SPb^V}��?s�����㵼N~ּ׋�n���X���i��I�/�'R~�q/��q~��my֖e�>����OR�'ia{��O�;O�>������΅�.}|*a�@0>��x+`��ꇞ��3�6W)�F�� ��ۯ��?X���˿��N.[��$�y�:K�L�o�=���r�䝯Ź'ɴ���XX\���^���N,���������N���Y�l	���2 �
>��Y[*�Ͽ'Ѱ��o�}B#��>�������E >�}@e�� ��>��r�z6>�@�~���̳'�����s�v�%��^�{�?��_�2_�7��ޓ�����$�!���|D��G�Db'���j}��VˎK�����#���!b>�tş'{��K�Ŝ_������N�Ş�|����>}��2" v���'Y�kk�5�K�`��笠p��{�r^w���@�tmz�:֜�>?`w ��7�d1�����:����認�9wXT�}�����[������T���W5�J����i��+N��m��yU�֕%�?r�|&|��Ov�4�8����I�3�*��	P�������&`"N`�u�w&�N�$6�O)��~/�^pxn,*����x��i�WԈ�.b��"�o����E�N[�z\]�6t}\D�7fk�K7]�4�ˊ�jJ
�)˰�T���S5��J�b��lÈ!rV�h�5�K�6n���# #k2c7��� ���"��o�y�f�F�z��Qf^I�b�sc*��uЭU�>�����U=:>a���f.%�cMΉ>ɥP�$뤸	d�i_C�zk���S�e�t�(!"s�J�d2������|��[�6΁L[�o�;Qx�ZYYΣ@@�6W�-�#V3��}5�8`���;�F����'C��=G.���N{��D&*N���u@b�.�5;�N����hȖ��a��E叁;�;���2�j-*:6�	�'�,��o���|�J���U8�nP�Y�].�������w9�1<�|�ǪqS�LXb�&��Z�<w_A��u@?$j�v{Bג}��]�i�~�9
C=�f�	��+��Q��UM|���3L��W7ȧQq? Gx��y����x�$�q^��)���y.y��y��Q'�4o�m��:�\b�30���{��o�4Ӣ�����GӮ�V��߷9���+����N�ıJ���`5��W��<C#�9`x��r9�[&x�`1�X���<62�V��(;��������ARnncqli��,n�WZU�󻓚�Q)C��&����aٺ���U�o�Lȫ�O<��"�r�%�!rc.H��o�o*��h�ȵ9{l�f=�k,'�]��mmsC��2ib��45��s������5u-c�K��W��зf̓	}�W�EL�I����?�EY�L������0��zjG�� ��]Cl����,��**�ݙm�3�9����~5�N^�<�%b����ᣬ<��d��CU�*�Sq�e���~�E����L����a`�����8�#N���:CV�=+Qc��b3K�;*�N�9�_o�/�:����xӽ@���ـ
-q��W)����v��L��S<�.�P&+宾W���,^�岲)��n^�zv�7��԰=����a�Fϩ� ��PP`��gb�(�+��5��l}q�!���&�����s6#���B�g*���?x1��LtWBBE��R�[��_�-yx`\º��cv��S/s�K�j�$E�F4-R�V.J5>��f	��i7���S�kL��<���M�iJ�*�Ҷ� �_��qf�uHMB�*x ��1�)V��'��Mk�ݦ�>8�M����o
�����8!���`-���)�W�Ԥy����n��K�Rq
�Sl���, ��޶�q�VW:�z�{!������Yeh��3YÞ�Y�"�õ_1�Zj�Z�[%�i�����W�P�1H%�+���ǫt��qs&�\�6��ߔ*���,觫v@�0��'ꪪ�2}I�Za*P�q�Oq����L��x���[�i�pb�.m��*�)M"G2ng��j��o���������M��W�S�H��i�ޕ�s�:&L>i٣W��K�H{�_�xF*{�9��/h׼��%�0��b�X>�G��K9�M�І�.��I��wx�h�Θl��vq7��t��{��]T�����5x��*�an��Լ���W���d��7o��؋�e����DM1ꑸ*��x���,/�yS;hV&��lO;����4b�ܬTFX�ғR��s�,r=����� s��5]�F�={L�;��Q*��މ�v6T4�HMY�
q���L�J9�1���ȅSI�N��w���S�!��;5��&|�ކg�NƒX�P.�< ���j���ُB�K��r�\�b+�s̰q�&zO�w���DhꙷIc���oufY��>,T >�Zx[K-�8��4��
��:b	�N�A�U�o,��vC�~pzaY:�q�����⨨�[JB�L��بީ��?o<�����Q��+�Kh��,W������B��^nUܸ(n�V��2o��]�W��Ɉ��Ksu<Z9����I�cu��.Ͱ�1�82���԰�a�!:��U='l��wKBY��t�����I�v��o?}U��Uv�;��puM`���L1�������
ڽ�ø �>�~b����!�c����m������%s���b�O�)vw�r<kn���u��o�`�d E���ێ���7\�{���X+�8v�b��SUK��sv����H�e��L�^�9
�ٜ�6*�Mz�ưq��\�JG�cWq�X8d/�8&.���ȂoKG>.c|ۨ����z��e��&�{=�	=^H��~졨���]r�cr�<>�����[VYhu���5f]�$�j�����eCc�r;�zi��ȿ�����[\>VC 2 9�:+m+������3�m��9`k���ϓ�"&8�v�B�p_�ਬ�Z7�H�<�Z��%y$Q��%�lgͪ�1���e�?��c�~�����Y�b@/'��^���z�➩5�����*�)Y�w�N�J� */���]��Ҳg.!)	ZX2�U�t�������I�:��=����7�������̯!E�կ�w�5���K���>��3o�Y�<� 7��G�M�m��2��9"��+krg�a9M�ңń��6�]��}��$�)Κ�x��U�E�I��x�����rë%I�Ъ��<�+dp�zo8��tI4��Y��
�n�^*�t+����P�VMGo/{x������}_UP�RY�أU����kƸEC[X���`�9M|���WC��駋�t�Ӑzj���w���zE�}|�\F�T�`ʃ0��|P����T��ح3!�mV�E�Yۉ�#�7�����.����ڞE��I��mh�X�ޅ�����w#|�<R#ޥ���{�r��U��!�-�)���Rל�����C�N��O3FU|��U�Tj�B$ �5��Ň8'��4�d���]�ϸ�zt|õ�;��\�LnD�h�Ɏu���Ţk�T�U�V�$�6�`3_"�	�J��!��>��_CθB��ETd�v��m��|�����p@� B)�V����9���������.9봎�s���/y�sD@"���_=z��f�'�シ����P�v��g���
tE-u�AmW�q�r��p�u^n�U�d͍p�wp��N��Ҍ+�E�Ai4g�g>qT��s��R3_P�\��w6�#0	f��H���ńKnp���k���~H�:�K�������~d4G�����=z�*ɲY�:�d�X+]^�VLŵD�J�/�V�A]��*o<�焅[yr:�<�����k�
�����EoV�FcmB���`�\I�s��:`�@[❑ASC��+$���u�z:96��.O��F񸓑'��R?��U}�|V�R'^�7��������FZUMBn��� h�,�T��}(��	�����UW̖�Mg�g��1�/��1������Y�<ɣm��T+�Q%���PuT�Ե�m<�%H���4XU=��{l^F�NF��O�/���`���ޞ�Vy`�e�;�M�k�øb����eWK
�s5�89�I�������0x_��ϫ"�8������%��_
�O�����W3g"4�wA����WSL8�����ue#��bb���M+"�Ft�2��1���.5�}YWR.�����U�}78Ɓ�Ź���O)����`J���HE���R jg�r��EJ���Z�!�`�z�n��]�!4qgmEN��u�����+��Y5�s�e�����/�nۨ�zjN�:���K��M@sM��9�� ��k�y����{�.��&*��\it�]��G�7iu�j��d����&�/WE�q�/�] �¸_�G<r�c<m\�	�N��\9B�����	˸����N��7�h�/�fJ���\����\Z���z]�ͷ�}%g>'6!�UEB]�]V�����k1r�Nm��T���Q�$��kHUΌ<tb�Hn�BF�س��e�H��d.\�vy�i�P!su��s-,C{�K��J��ۦZ ��u2c���"�ҍ�F�}����A��Q<�U4ى��Ƃ0��5Ӿ�������Nm��*3+r�o;�b�Ky�Q\-�R��<�,�آs��r���}�hI{�۔L8����s� Dg�Yp�w/��cM�w���v����	�z;f�iߌk��鮜��Y�6�����#�uZ�G/o��0��r�6�adaw����1�b8�SX�r���b���8���u3K�Pq��`�Ջs���
k���e�p��e6ެV��M��v���T2M�uX�f�3��[�
�n�b�Ʒm�b��������[{��c�G��%S�-�l#��*��l��ԝ��v]�d���F@����AX�i+<F��8nW�-����{y*C�lJV\�D���j�j�Q�#7����c.�Pm�CI����)C��J��0D�u L]r`���V4X�j�]o�>4UsTp�g��� �E�rj�y�
��|	��S�����{S��A[vP�7n�
�Z��E�Z�,�%7[s���j4��霦3Q[�S��hn"��)ʾ�D����7��d��JY�95,�L��f��C4o9r	��㶵R�.�&��#��m�]o��D$8�}�N�¢�����.E6>�.�hL�M��tS/�\�H�;Ʒ*	�M�z�^ehw��;���t�v:���
%lU�EC���E��wn��l;���t���'�d�Ƣ!�d���V�)�[a�7�c�+���ׄ���2E�E@��L���&�#��V��J���֮u�#���[�loY�>���J�Qf(�R}[xUe�pj{�v�f��]n�9b�`�L��i�5ܦ�tM�}7N��2J֟Z�,Enr�|&fdމWb5���J�<���qW.{D'�%�o2�����`�v��-Sԍ��)�J4�u����m\��Ǡ��k"�J:��f�ʲ���(ԝ՝���*0ꦷ6�A)���o=R�J�y9�.j���֕p���9�ʮE���:����(X��#�o*+a��:v�����Z���|�Zeʹ����O���6�!w�9��W-M"V��u%jBpm�x�T��!KJ�w�yw��/K���h��`�L�rUvFFf�~�\��5�Yft�`��Fv�1oڝ;�ƭs�
f�+�+�m�8��Ģ�e�<��nv�8Z=(V�C�)*���+��9p��/0��*�Z�V Oӧn�L唩ŵ����,5���^�WQ���S�5ݪM�������r�$]�R���*.�$,-ɩ!D�H���]!f�m@�$*)�!"
H3��F4�JHBMDC.L�l�#."��m�+F��h�3J�m2D�k.�B�i�JR�Z@��d�J���-� Y"Af&� fXD�*�*" UTɤ!b�Iq�4Y��Dm1
Eɶ�����V\$B3T�t �hm��U���DXFڊ��P�HI�Q,X��ܛ`�]P�L�� ���R!jlTF������B$�X�R.M��2ah��H���Y����!D� �E\��I0P�L�$""d��%$�I�ˢC%��M�Hm�&�B	@I2܄��*.iAUp�U"� �QD����+F$���ǰ�k��O�8�|A������2�ĝG�s�H���\g�)��]d���I=�K�v����\����G�.Ƚ��ӌ��}p� �#"8pd� ��@��Z����o8P'��bw��`����jFes1��F�s�J�X�(���}0f	��ZM�1̬�yTr�T'�Ia9�P����o]��8R��N�q7f���'\����Ɨ���o��5��iV͙N�:Ե6���,9|V�@���|��}\�$s��6p���w�\9�~S$�5Q�YB�4�9\��x�;)�=<"�z_��3cx����c�0��d��� ��̚��������*��ـ��fcU��.a���j�.��ȏuy@ѧ=޲�▁�q�,����4�N��P�*8�2K�\>]�X��5����·�oPW-���&�MV"��������=AL�n|/���[�hZ�Lt1WKt�|r�8�W�4<�J�r�ff׽��1�Փ��*�!k��j�b��ى�UԈ���*�o��ʝ�CE��t�t@')�-�N�F��B1��Z�����N7��_����u���c�=��O����i�S5+��^a��V�T�
�X3Wb���|z�<^撝�Hn�,}%��bP�UW�ë��mk��&�e;����co}�^�S��]#�2
��9#���&.��ݖ6t(>�hl�\�e�)f��jCF�U,vu���!�Ň�I���������P��_�  �;gV����@��*��C^U*i2��CY�M_�qγ�!��ۦl��te����:V�V=^�p奣�/��.���UӇe ��1�9�X9�3Ԋ���nA���1<oc�n��yjb���t����(]:P�X���A�]XY����pi�P���f.חà�o��fU?8=0���Z\v�Z���*>Ґ�2��P�*\��y���*h���z3��e�������MΎ��h���O:+�?C]m��3��z�C��[z�#����½��Aj�d3����7������&\@E��^v�����oo3��*� �0>*�U���&�&�e��q�1�s���x�F3(�����jR�����C�#Ǥ����_����5���dJvٌ�����.cfD�3"��϶�&��uY؛n����B��P� �}4'��XO�<>���[>��q{���.�7/��E��-	�2!R�����;�8=f�䪹\b�z�y�@!�1�n\D�$J)�cB6_Kc�q�K,Ƽ�7��)$ݼ�C-q���Mn�g���Ԍr��j�k0J��yS@�@�<1����{�m{0Ц;�Ќ�.v�����l��r�!>{w����/F�z�w5&��u���\��cM��
�ﾪ��4eF���Ly{�OԒ�Kσ���_X	����Ch{���Zj���E�wʏ�J�W1���B�\����]�c 0�`ah\�A��OK'����"��|�7��+��GnVv$����7����u[:�]M�3a�}��xe�=�d�ҿ.����h�AgHZT.���͵���߰�k^����>?�^B���_��Bk��E�7����@ {�ϼO6i�,�����T1`�q�<N_ݴ��ֲs*����cLMJ3+��u�ϙm��ӵxq�uc�9�#����F �eWB�T�<6�0<,`�.��M��v]s���Ҟ�=�d8v��-�&Q���<���1�Z<�3��%��CJR���4�҄U����}a2Fũԧ�S��n~ϻn�e�@�j�����I:�Y�ި	b�W���#�U�,�.���?0���6b����ȉ����6LT�[�j���}w�93'h�I�%�V�S)��^
�(P�ԭ���!�~��n8H�k�|���Wn�����G�T���sܝ/e�P�w�s۩��o�$�0gw˴{�To�vs�@���f�Z��|�[|��{�z�)�+��.�mD3O�jT���:Y�vP<�p�����mTK/���ԳV���R���g`��kC�+�yr�r��h�u��_W��}�{�y���[�|W�l. d��<����ئm��ۯ��r��]�b�Ѹ����ZRT4o:�g�sB�RQ� w��-$Q��v����+��i�0���#���sVz�Cu�M�w��K?L#� %P'I��u�n�c��tڷ�
2���f�L"�Ꭷ���m�Ct������Z�Q;1����E���dU�܌g�q!��h��<�*�?z���m#C����(��0	UJL�J&!w4z�����
�N��ev���nT�h���>��S:O2h�n��PN�1��W��Q}�ɭ�Ψ�KsT��d�5V�n�>�׽�ʈFtԉ�i���&`M욦���Q|���Ӑ'Zw�m�p��;b�.�1�Q��C�����\=z���K޹�'tm@�.V��H���pڠ�,}_��x,\+ʔu����$*�������+*�v�8�5�2�=����j8 Y�s��S���	y��qӗ�� ��ʜ/�>!zw{�,'��5tU"q��g�jj]c���r�b�:݌@�����9F�(�{��u��mo�u��F���6��y:���3�Yΰ��r��	�����m���X(ܜ�w5c�ZbyN��a^��ꔰ���\N���S*Y��U-��5�-%Q�Ѳ�����������\�t+�X �
��Mzf��T��)�\��?-vi<����;O���r�-=aH�"̪�����<b=e�@2���<��u���q��K����^�8�d]��w��������$����KG��鋊�@�Z��ѥ����Ӗ�Q�Mz��.V���كc�ϟ��c
���ȃ���pt�s�*�3���0�:c�ޣU�>gw4��PzŸ��g_���³���b�_C�L��d$:;1�m��-�r�� ܋��[��i���Z�k�o�÷U�P.��h�0���i4)�.{�3���z-��!�	MgS@�_���^{D{Ɲߪ^�p�p�n!��N�	D�9@����5��5M���h|7��q%q[�'�ⷄ��rt�Ȃ�6p���z��X��!�v],o:�ܜ�'��ũ�� ��5C�tE�7C`5�ϭѿ���_�Ͳ\����ꍚx�'�d���q0=��Hu\hiTR�u�5�.U���_�����GqБ�N�g4P�T��-x%�"����ɺD�[�F���/)cHf W+J�V(\�mLT��X�|#��p�C`W��>͊��Q����:J�7jk�_�5��Y�zYFV�������}J@�keN9ute�P���8�ַ����,7(���Z�
$�3.���S�}�������Ց�Rd���Fȡ5��0� ���X��ҳX���CB�v�lS�[��,j
ަW)���n�P"�s4��$�9��F���e��1WKt�זaY��T}Iǯkjt+��VӴ4\��/�Sk]k��nb�ML�����ls/a�Mɸ�=7.0�	>+w�1�uo&0E��Q�j�ρ	�u�㪦�yz:�U1�j���o��XəҴ��~ܘ��1u���(o�1� �U���k�P�
�\&��4p�GVk؝<�~Z^Y�)ٯ"8p�ς_B|�k��YGe ��1�y���S�37T7y��vԈ/Q�t��z
hm�׮�42^�:Pʙb�����.�QS��}��@u�r��? ���"�n[=���9Ɵ�1�,P�T~�T|-�!���vOp�ġG8}O�Yv#��S��&�� ������GX�<j8�J�����`�(wκ�x�w�_g#��==N�*=���O2�Q��Zn�H[�'�~���m�H{j����G��˗P���x�@{>�`���8*6+<Ҡtx�֙��۽��V�Y����Q0^"���:'������ا�+7c�X�*#��w^ۆ��]�r����igV�K<�+�8��<���E�����P=XS�t�����}�}�l��;n�g;����q�p44V)��{�M\M���˘c��' V�g��t��V�/S�M��݉�^�@��\��)W¢�eςƖ�p�6a�zZ7B��h�á�kg�Qѹ!�&�'/�T̄IG>U?*$LI��B�C����s�쓂��u�=c}5ؗǪ� ব��LZ%[5�J�t�<���zi�:<������"��o�r췮i8M�/�Ԅ�?W��2^,y����(��Bӑ�D�DMe��Q�c������pڽۄ!s�a����2�r����p����ן<���L^�<���j�q���<��(�4�lz&R�K�����aW��n���kG�_�7[���ڷQ�E�&�n�i�Wir��B,B�mg�p���`0���3���fW��Sާ<{��CN1��i�u��F���iD�Q�a��ꜣ�<k%ޯ3^�����n,�!+��@�5�^�����x��O��w1]�2���x?���@xfVV5]߷ \���g�"�u�%���mؑ倝�5�o9pO8(2�y[�rrp���� 򍊊l//�m�g�r��=E!c,����"�ˋD��<U#��Ɉ��t�]X��jQZ�8�X.*;/�:DpGg,.;o$�*�������ꊍ�r��w��=��
ӿ���;*~HuOv�<�q�G���ύ�uT��Wpwzt���it���T>��#j�or����T������m��q'J���=nN�V�y�BՃqz�"3� �P�]����Q��^;��_��1���h�U[�m����8f��1՛&�^<	>i@*E^ʦ��/�P�:�==�9�9����mNѽo�UǾ݁�d�6� ឪ�� ��"�*ꆮ��rW�=~'��-�Zبx8֎�׏��+'/K��i�8�����s/�D	��$3�{��:!�Vw������J��%�9�/��a����wp��N��,�0�f8��t�3�2�3O�d�N�OG�'���7q���Q�.�G&� ܢa@b�&�mցq��A��t�)h�����0�u�\��~����|���+��e�UM&�y�4�.�RdL׸m&��y��ڋ0����_#5�v�{�Y�����w���r�'d�&��۠9�U�������/O�Т��o+01�(���[r���b&ߜ�KǾs&������R�Q����Җ@G�n��۵�6��e�xQ�P�n�c�f�J�̃Z$v�����^E2�&�3n�5׸yRyj�W�� ��j�ު��t��AQ�5����������qU�?{S�XW��D�2���.�xX�ML?:Y�~���K��Q���,TH�y����^)6lc��}�[Am�^ٸ}�a����Z��`�����$�HY���L^[�7��Q�n
���~��Y�
�@�u����B�
���ߞ��l��;�n��+'d�6۾ ^��;�e�fr�f9����WR/�'3`�,3gU�؇o�xJ;|�l��՛���EZJBe�fwY��o��ڮ�s���A2-F�ȽKK��K���yc9��	C��+u*e����ˀ�	e�\�|�cT�7Y�����;��i�����ܖ.-I& a_�gB��}1<���_-X=�`2��s�,/�OV�JN��Z�^�>��ڡZ�1��+ă�W ��䣞.Z<eu�w�\��F��z/���o���o�zS�3�m\>�3��B�p�,���BC:�B6������A�w�C�k6�����.T����F�v��p8iR�W�>όxc�fj��ke�P�N�����;>��\�W��Q\��3	(�Zي��[\��#P��!p�#��6�Y�})�ȀV�tC��}��L��^�=�ib��o9-/�7��-Y�e!��k���!�gc�B�J3�����n�sqE//%=M������z��q��̲X����*��|���_���.��݄�of������&"7�t�R֛E�s&5��5�ƌǠ֙gP_d/������G������z��S:�p�}Tif���"s$�"N����*zW��͍�c+�[����I�.�*{�1}cRVpi�%?��D��f�s��bGG���J�p���]�U˃�,��9{ˊ��&L6�Y�ي�Aή��YD�����@��5���/�{�8��8����A%�w�ۻ����r��\���d�e��2�߯3�n��'��7���&��_��wdw[/ᕒ��:�"�k��vG�Ń����_u]H��Z���boo���ﷅ����B��h�L��q�)���V�@!�5����5]Aˏ�s�uźf�꺮����>j�v�ق9Ý2z�1`���6Ҟ'�V�T�{��*�L�bF3���v#��vvZ�ʂS!?w�ڠ5WZE+~ ��̖��>{��8.�P}9��@+��D���w�4oTjN�ڳ;�`E�V��h�,�nly�W�ei���P�D�:�p���t:�G�P��;OwN)L�6�r*�*��V���4d�dM�K�5\�``�D���R�n��ä����zΫ��rO<(�� t�Ź̵��U��)�WtJٴ�}�«[�볏rA���Rklt:m�rj�{�B� ��\�}Qk��R�[u3��(�
ܬ�q�����j8"\�cv1jS�ӄȎ]F�J׏�:O܋^�!h�C\�k����R�+���h3;����=Pb���#���8�gU�Z�2�E�.��2^��ru�èmf�xp�������ȱ^��v�ź�R0(�ّoU���w�a�|;�_aQ>钋ʜ�xN-�f��.x�̚�=������QmԳ��F�"s���)�Y(�������Z���m^,
47])}H �8+��;8�=M*�3X�9uyk��,d�t�8�&��*8rm�b39Y�B��Q��;���*��ۡ�'k_MZq�J��P����7�h��u�%Gs��uըE�8 ��`&���s�qd*����7��D���Y�0^:�p�Ԉ���8U��*�Bw�X��;cYu�6[Kq�
pc�1�C�@�\4T��׵Be�*+7�s�֪=���1]N?gkѱL4;5�n� 0�Sj�e>B��B��#���1U�ĺ��"��b��B��|F��&�fF����kJ\  !|���:�E (���7���-�f ��JG���hv������fي��3"W][���݁\Z��1�'S�w[��1�4�*N�ICF$��Td�/Wq<IKtU*�t��{�j�U�D���rJvo�p�$��a>yDWΦ჆ ��I��n�ؠ��r�*+I�KGV�A�Q��قR���+�֓���u(�]��ѵ��0qgMЈ�t�܎WjsP�@:�7&�ݹ�FqC�����
EA��Ty�RV2�f[�f����]d��vJ����5�/1��jbe�S3Y����i�a���J���F�ǧ���|�ã�ۏzr��9VqS+�9fӂ�Q'y�Pm3R"YX�!�2�A�A|�픳Op����K�K����u��oa��bm��e�ϣ�ۋմ��Y2���<���F�3FR�Ę�:u��%d��({�i5��;�Ja��⾚a�|����e[D.��C=��'>b��ӊ��Fۏ��W
`�q�&�"�:ͱK6���Tt#5*��j�v)Uq=a6�GJO[O�[̌�{��W[������)���↺s*u��圐W&^Ǵw�L���!���BUo���j���]����d���,�"��S9�O��.�A�H����v쭮��ː$��[S+���bf���d[Is�s(V(ù¢Z�/yVu
�0'¸�Zb#:�+
SWpoe#�̙���wRͲ#dLT�!]�TDB ɮ�lRfDmq�k�	""���!��HB&dA��l��TړF�Ck� Ci�j�2]�Tɴʓ2CM��&M	�H��ELզ�$&�&��2Č�`T,m�2L�kI�f�˔�C$�b,ƺ�DP�H���TfB&a�Aif�F����M�$*	�Ԗ�J��6�2da*�DB�B	"��*&�v�.Y��@XL�2\��!"�"$f�4�Z&IBF�,�,$!I-�@����DD���̍��4K����&DT�-ͶB��M!b��E�E*	K�DD"$��X�A��$�Y*-X��E�6�E��>?   �ݕ6J�o0�{w���C����f�����Uo"�H�N���]���E�j&>��I"cZ=L��uIu
l�}��_W�gnrs�ߘiѰC�l����gZl?1�P��gJS,EDN�����c�G;b�cm�o�ឯ��P鈸N[=.x=Ed4�c\X�+r���*����)�d{S�c���/һ�i�|A���M�P{ף#\L1�����	��_�����)�ۭ���2��e[a�5���Te�쾻������AJ�d3� ��ީ�~S:�rD]f�w,��>����m�D���P��z󝍇)����q���9	��!i�w=:Lésw�N�y����'�BAJ"�2JU�)�>B��-�����m��22���8��a1��5\X�W[O���~�~(:�\��Ƣ#=
r�������2h���)r�##�����mQd�'�3_D��TMq�'n�s�=�*"N�&�W>��26��V就G(�7�)�L+֮CT�_sT�y�,x+�9�"��v�Bҡd<�7��^4
�}���>��f��c�V��_.{l6������',/ʱp����p�A�[Y˖Qp�=�P�2�;,� ��'I��l��W����ށ�J�U:CuF7���;�I�V���G�e\�Ur���2C��:�����������ٛ(�q
���
QPG�_v�awY2�4:C�S�y���r�9�[ɿ������_,~���v?X�0Gf��,�4���A]}�n�~%}9�����&�={��^����|;�9f�nX끓�7,\��'N�^��ߠ����.d�p���סz�
\�z{v��#\���Ƃ��Щ~��_��3�F�S_1�Z�Y��2�jMJZҕ�v�ÅU�FC��{!��$��5շ�i��@f2���x7i᫫�-�����%i�@X�0�b�̄g��+���>���]�h�U��Ic�2|���Ex��GA�2h�,}NFY���$lZ�J{^S�.�1�����Z�y��L:��2�c�x��^��g�X)�j���A&�c��r?0���6b�cy94���F_W�8�כ�-1ޠl��N��@�뮚\i��+�5�Bk�J�d2���iFh!��=J4o�1�}p��M���G�$�q�g>)�1Uc8�����߷d��8�����`�_\|�c�܍=g�0�*�RQ� wi�C0�4?LMz�?j�N�=7k`��3��s%K���,��^o]!�'���'�ղ��ՙ��:I��`Ef0j�����K^����i�բ�sl�[7�$�1�UϥV�wj�Ĳ�C��E�����r#�'������j״�w�����wҹ��UU��X�`��P���=��3�m_��{,n']��=w�ĳ�� %�	�`:r�\�L�s�KWv�h���z�����b��� `��5h�
-��5�͡CG���ς� �3�?�PrD���7]-��W�ј����M�ؖ ��d�]g��=�7y[Uy�W���N.�����^mT��ozW�O���ĎY<ɣ�dH�̇N��;zv�R�o]�S2�^@�ʃS���;)���K;o���a�v�z��^�c5�<��o��cn�z����<�v۽���;� �s��F��p�*���^�}[9~Ɠ�$0-�Hȱ��T�#:�ϟW�j1ڳf�����3�e��J�V�8�R�Mr��=Jr���X��;~K]ݟ�z��6��u���9��s_WՕu"����e���gG�mr�1d�hA����U��$�	�AW L�.5]���gbru���ا�=��
ϣ�����Ѥ,�,��*�>o����a��q�ɨ�<��u�}�*f��w]S�۟�);�dE��jRc	����_�*�ʅ�0�b�J{��z�r켿h���
����mZq�(=&
-����L���y+�:d�v��a�252�.%mrW��s����U��X�m.z��V�}	��V�ݙ{jMe�<͵U��������׼�b��h��#!}z�qiQ0z����4�]9�T���C�o^ι�/fvgo���� I"@�~>���V��]:��a���,z�Y��e�v�" 8��1�n�"fÕ�*�3%�[|>�P���Gj!�u�Vx��1P(|I��@�H}����=�^*����������Y����F��C�ޯ��JƃL�N��TY&轜ʋ��M���Va@T�P��_\U�w,���u:�Ľ0E�:�']���"v��:����=/�@����-V�ceq{��л������}�l�s`���:�0��q��7�z��U��<�S$�"O��& !3�GF�V�xj
�����K�˫2�6�Ŷ�wJ�Ҳ$G��/ *�*9>$:�44�jzƼr��3M^Ĵ�������+�Αn!N��	'F�Cs��F}����g�فQ��T�1���Pl���Ժ��.!'wA���&�����^T��W���b��
�c�^x�3[n�{gO(Ȝk�r��Z"~F�q=�[&Q��n���c:ۨuyj8<��U<��^N����9fT�˒�Pd��gKFL�]��,��4��%f��>و]�1j|35]�X���;���a���Ad�g]u2�TՒO着��"r�A{>+�Q��Әn�X���lh���7�Sp��f�%�MCs*:��P`�pL^�c��{���	�Z�@tR�W��OK�>� x����`�R�hp��
POAkH�������~&��(d�������(���2�(��Ʈ|�i2�PS*���W\���<���0�o��u�nU��\��˪K�0���^g��z,���;��U��P��>�7i��$���H����^
wI{Ǡ���@�׮�?�����U������gfr4w�W��WY	�}VF�_V���l���p}�g8��G~� F��2g)�������Il�	��[���3th|�z�Gl"���q0�^:m�w��qs��\�%�q��7�x�n���`��}B�����=Tz�7�������C1�1�M�ꑢ�O!|�m�ս[�$�R Nk�(	
a���"�X�9�����;��0�i��X$�V��+(c��W*:6��i���摚S ���$��l�e�}r��.��G�o\R�1,���Wd��Jݺ���+i��H�<S�l�Q�ߺ�Y��X6��lk�}~׻@mc��.^��\c�V�*�n�^bm��@�`���d�0�ӭ[��N�N�i�5��4Yu�����9�xε�a޸�@�U��&�H�}���}5ݒwy}=[Hǉ�-��X���D���8��+����BFz&.��^3ȦBu����xHmj�\͟{:�Ru0��ڲ�A1h�l�ХLM�'`�~�ƅ&n�F���t�j}	xt"Y�✭1W�ø֮C�}S�G5L���5�
��N`����\�Ё�q��6gw����.�UƇ�.��h�-�B+�\��mMQ�d9�ʱoL�y1k$nb\�oz��9�U|�H�V�l��~��Ǡ�R���.x�#�]������R28OS����_��ظ�b�o��%���Ԫ�=�ϴ�sJ�v�Ҩ�字����G5����<�L��xf:=�39�X��g�{Aj��w��8�Ȥ����s���L�ck���洄�sz����O{��7�s�A_WbI�͸�?v4ʞl/�'�vb|�>�}m���<}2/����=c�;��V�ӓ�;���6z��*֥�����F�����ح$�W���Gmu�Y�v����۞�#*������8��������wQ��{�b��g-�A��ڇ&�f,՛������/�OV��k]�ڕca��Of�tb34�lTor
�`]�Y�_f/��t_n�8���K9����視u���w'0o���0:�K�ժ����yxۃm�:�*��rJ�s�<nG�cӀ܂��ʤ����
�T�k�I�@֪[<'#B���k{((5�8z�
]5G|�J�����6�\�
��I�ݮ�ԓR�ʖ�7--k��q�Oʈr�

~ﻄ4�duuvO.Z����@S����g;k����k���c�OtW��Y@.�;䛊���}��&n�[���A�R���\� ,T��W&���ô+��C�GU�5��v�L����J���sS˶��Z�Ĺ�D&�;���M]��L�hv�jW�{]0��&ap�	][ܡa�5�N"������� gj)���E�pn �egz�%[�B�xj�m��>��t^;�QV;y�#0�����+T�[��ծ���7�_k�z�l]P3}�i)!�h`�{�ؘު����-P -wfG)}��R�ϻg<���RC8̭�̝2�+�P���؞��Y��%j;˴�dɽ�F�u󡫭u�cn!QH�c 3��xc$��bO��%v
5='���w��}F�'1V"�=#�_U}_Vn#��Cp��t_.�nV;�r�k�|��^93F���9���yR�Us�+w���=�/��Xӵ2�����n���7a=�pev�-�
��.�	3g>�絇���~�+)�-���T�8���d�j/y�}�Z�}����u`�W��uCV5����|��p�-��3]�Ck�~D����g�[9�j�Ƙ9�:�K�P-t��i3�9������lt�qF������7��g��@hQ_@|��=��ꖕ��O=_�.Ρ^�Օ5�m놳,�m=�mD�����Tץl>���V����}|�%xڠ�=��-<�x�dF�ͧ�q�B?K"$L������>hB�ڟ���Jۺ��,���k�-�C�؞`<g č��F�`V$��3���Y��L�b�Z(j�gR�\�P�[�7wF�LL�4N�CYW���揓[m���]�i�u��ɿNh�ɭ�jD�V��'n�*4�\������[]3ڒP�l�Iձ'9q�1)F1��䠪K0:�Bm�+�6��˴� �+m)a�y����ܛ���������H������M�S�e��JQ���S˷prx��d0:3-���f�=�9)�4�8tÅQǂ�Cg�y��nb
^�Y���W�o1$2Z��%�2uĶe�4��͸�a\O�艎CdZ�u9}�{������#�&���ͣ����ⴝMB�jpw�λ#����"v�)+{�2���U��c�/'M�ǝ��_Z�z��c[�ww�7#U����^���d}�����֔��絑ZN>��w
e��^է'���a�ej�5�~�J|k#�3(����8Gxm�~p֑<	|;��{y�Y��x�3�F�?&�B~�]r��=�b���&{��.ʍ;M�bc)���ˏ޽��Y[�{���Y�n��`���+�yl����J��cU,����?s���F]�7{�oe�,�!�k�"`,�!~^��&K�u�r�^��p�|��Q�K(X�e�;֢��7/v�}ᗕn0���X�[jW7H��E(��\�5';���rb�w-)DD ]���0v���wk�q^��ք{~*끵,ґ����/�&[*��Ƭ����材�A��[�-���7���fiWϭK�}�Z�����)�Iﻕ�K����T�j
O9�Yn;,9x�I{B��������������)D�}��+䘿���M�OK-�mj3M7V�
��n��y����Zӌ���9Q�g�B����1E-���d���Ę�]a�orEi�N�v�P��l�r��!qK*Հ���KZQ�~�p�'�;}�ܧٷ��i�篘o����B�{�(�UX~�/kY�W�a39�[=r}C�a��ڿ���h��������p�3��G��R'���֜�˾��WFU�ws.'ڿ�V�x�U4�ÚMƽ_dY�1>=�ǒ~M�{�n�r�է\K�8��Dw-��+;��/{p�M��,�.�1�ӭ��������:E����m�D�ѷ��m}�Ë��1n�ӊY��]]�AE���SZ�d:��xD�{�qj1�s8�[�Xѻ�-��3��]#2��j]<��4;.����:�j8d��we"�o8:;N���t嚤�J/�;�_s����� �K3"K�n����s�&���j��t�CV]�jU�A�W�>T�� �Q�5�JAj����]�pMh�۴�p�X�SE1Z�gxۺ�Ϯ*ɝb�	BO:�-Y ��!���!%�5�e�.Yگ�I�6+K]dMl]��4��z���Z�<o��[#�5a�ի)b]F�B���u�hjc�,�H���uX�ܮ�G!<x����oV��e%]!9��4����:���3�qi�<����S�t-��8�j�,(�֓������o����Sv���sR��GR�h�֤V*סE2����YL���i��Q�z�.�u��B����w]Sud�w���Q����N��r���um]�emJ;q�MڰV����p�d�8�Q]ʵ���WE�b$�2���w��\q]G�'K������mV�;Mh{�k9��*��GR|��_�!�N%ӥ�Rڗ�k��CO�uoe�h]��qn㊶F�-��@vV��G+�n	F�� �ˬ�]��:L��Q��ڗ����C0�3B6�Yu�2�&إo�R<x��[v ���O���0޼�(GÖ��0#�.��C�@�vI�﴾X�XS���B�ܐ�mA|V�X�iY�յ&�CS�d=�6�۵V	����	iԞ> (�7	��u�V�V�q�(cS	n���++
q��q5��@��Mc��j���@s����M ڶ�q��.���0�]]:��d�]Pe�.��B3�̧f��2��֋](�1+Υ�D����ԯ�f���b��B6̳�����ȴ�q,�3y+*jJ��Ok/ZZv6�`J�x�g?��ty[��� �9ń��+1�G**�j�Uqqd9�-�X�j��}V#�b�#�Te���F�e5�������1��bǎ ���*�/�ƕ^�z(-�KT���|X�)�S�y��w��n}�,�q�Y�A�.]n����u4���e�ݺl����ofJ���g�pV�fu�m��:V�գd���[�LNj�Uװ�4ś
��ْ�S�]����j�Yۄ�x��Cy�\{ �WZk.��IV�o]����c݄���T�nt*Ŧ�].��"�OTz~�I�������͕�4b	h��0�vv+�9rG�}�P�FdX(�QNk���C�gɀs�/Ud%%1��r��~]��6��\Ubր��w�N�����Fe�j����S��u�4#� ��,	���Ϧ�Sr��`?�d�,�IQ�h�}� 8��s������\��ҩ����0�;�*.Q��˻����'-�n,Hi[op)۸�>���ˉ�
Tl�2�ُt.�̋m�e<��W-i�ҧ7���Y#�(
	�L����)$Q�[�m�XIVh֬R�L�MD� P��-$����E �*�P�HT�� BD���6��*!0Ћ��!	!&aɢM$D�d�l�qi4*� �
�i��m+&��EX��!
�EJ�"A""@������,fD��A��Q`�I��*3TCD�����R��X�DPQ,ɳ3H,$PV�(�@$A���@�4֬P�*�B(D����L��Ј�J�3@�J �!	DT2`�*&] �B"DEET �(��b�$�B*�@��q �$�QAUE�@TG���sZN��Ajs���6n�6����%���3�%��U��f�޼+s�����(1VL��C��w3#m�����~��c�*�cF��?E����^]�4��-+�V��8��HC�J�;��� �;:̝^�Rz�L�c!־��v��VU��C2��9P�q?�їi��:��_�=;Rv;��;$�u��|g�����Sɚ��u)fm��[Ԅ�������G3X�I���c�7���/��j�K��(}/;2���|�]�=�Ȟ2�eL�aHaj�z[�p��s�n){�yk��ۯ��n�D����_>W%'=!)S*(@�����=gT���{x�#��ţd6m�?��m��$�&mjȝ�3*��=��%���8����_�������r�

{��0�$�l���U.���l��,���W'4��{��v�Ұ�^��:3�Y�BP�5��K�������	�v>����Άo�M+��@v�n�Iqst�5z�:�&�x@�f%|>��"��}XF;���*[��>m��]�0q�E��.(��
J��w�U}����s�5��v��fz��#�$���NV���������G��*�pV�L�h�AOT�M!�
I�3��W�?}��vez�N�޹>��*�U@�`�sQ<�j�������9M�w�; ���k��曍P��L� �VV�畿'��q�*Ϳu���I�g2H�=�n5��NV�"b9�kh;uٕ�]Hڎ1��NgtsEe�*�m���k�4�P�yox�U޷�Y�m)q�p�<8��Q]������^��_�m�n��nVz��fw��/=��v�i~R�H��.�-���Ǿ^v��~���o�}Ղ+F�Jʬiڙx�|�5|�v��>�ַ��=N��Uv��<�z3* ����͜!1��ΥS;��/Oxey臘����ۡ�e��w��	�{�������C�c��j�uCW\*�-�ٖ���*r����[<;��ô���۶���TRG;�U}_WӪ�7����,2"ږ�:�jK�x�k�w�Z��6��X����g��ڹ��#3z��=��ם�����]��S��wm�-yq���m3if���U;��,;��3�]�e.˓~P܎�sI�z����pZF&Yf���QaÜнZ�y��zs*4�`#uӱmɬ݈u�J
V�ׂ৊��;5�AH�����^���E�̥�R�f�L�S{k������΃mT@����M��:��1эb��H�ie*�=������]�k��y�)JFS	(��
q�V�-e���{��p�]?����>:�Z�C}���]S�^�`��Wz��%�A�y�5��<GLw�L	KE|5s̀����^��'���RV��u�:H��W.p`���*��]�%*���O��yv�@����r��e�l�T��ޚ���æDq0�	�Ght:�
�3� љkl�F���^��znv��ƹ�M�MG4��͸�p��k�'���]�E;cc��9n-�Y��ve�8�j��[K���j8sP����*�5�_d����|P����U��_t8��c����{Q�XZ��ۡ����۩U������q�n��G1�mg�1T���=>�g�f{�O#�U�`Ţ:emʠlvs*�v�a���k��L�f96#�]szԩ�,*�ʊ��I�H��"�kp�7���P߶���S!��'Q��u�=�>�Ij:U�Am��&=;"t)���[&3��2�8�N�����W��{:�?{r1��#=��P����.�؍�=��q��n�mna�x��Zgi�ck����{#�g��g���,��o}����{��rV��Rp�P��>l'I��䶽�=�[g�7�qz?��N�=��aggm��j�������[���{ޗT�=�oT�2���6��C}�K)��g6A�vY[�J��-���ˌp����&��5�]�}�v�����cw~�>�X${E��ȱ	<��zsbj��r���>��}}I9��߾����<�=f�HiML�����PKэOb!.z��T��W�[�Έx�S�g�B������P��^�ڷ�=�cl*փ+�u8o^�m+��0T6�S�e���᣸i��onjD�w���\��[�܀��{�*9�V���'��T0e1ﾞ'r��gy9�[��%�j�+�׳aYKr���w\.���Mvpy%��:1-x#������C�9Zuev̼��+����w�4,I��ԓS��r�l��Dw)<�j�"��X�Z�@��j$���Gj�j�
�y�sl���̟�_W�܇c��>fR?����Y�h�'=Z�m��>a8�;
�o�����鋘�z��W�tC|���y���um.z�!�SK9`s�v&M���!s�U��56n��&�kj_T�ʉů����Υ������\a��{ν��S�	�W���F���P�U6��ѓ���*/§V3��m^�)���35I]��r���izZZ �]�]o,����|'�j������z'�Ɲ��:�����M���iE*?/h�0��Ǟt�£{\M�T�����ؓ7�l_Γە۶�� VO�aC�cl+���s)6��	�끪��TN�J��W��_c��!�}�S�o��JU�v�)R-�v/|5�5��v�?eXp_�V)W�d���yO�΀���{�l��v���KOn�T
1� 6`�!򨒓��	�N��Q�mU��<k˷̴�_T��N�v1�|�ɢO(}�e��/��u��� ��؋/*�sh��3���I�1V�)�?;{�ߑ�#%X� �!�*8)�Ι(fمV�4c�n���f�\6�F�
��OCr;ܫQ�6���$���_W�	���ֆ)�{�q���k眶��T(t�ϧ⠎�v�l��b�c�����	�u��������ٮ3k��9J�PS�wQ���Cܮ*��f�zU�p9X��>Y�u-}�[J�;ש����C�{f����B�]�����H��Ӑ��v�T���|��W&�7�����ˌ���y 
a��_�e�����8�@>U��~1{c��珜���=��k�5,��,E�KS�ӡd�l�c��ȘR��AeX�?[ܡa�5���\��N{����\cę\Tݴ���sPۍp�������:S0v����n�/T��ua��kWM�I֭p�E�[��x���Y�������M���q�;�6�S��+�9}p��4�Nw����T4veG:B���k�\��PlB勽P�w
e�9	�W�u��gC(i뵒Ĭ��K������İ��0��X���W�3�xW^��I��1e����i���v��V�{u�l�Q� ���͍r�c}j���r�:`u�����]���B�%c{�w�Ǵ��rv��q�G���c8�Y���+�������G��+rzG��|�=	{�۩�O�ti�����rsV����u/�w��0��
�To�ǵ_$}^�m��I��[�kj�9c�g�'T5c\+���L_Lՙ���y&����箛�/�m�LE휨��ǞU���9�;9����{������
�Id�)���mꖞٽ��l��7 Jn�I��E+����J��9���YĩT֦���e���6�ٶ�P�o/�3��8
�]���v��zB3�]J��Of�O/�5ٮ3jq�������v=�������i�=f��{���]'鲮s1y��{~�5�@�su���7���^q�Ttn`䍷(�ȅ=�R%.��������;T{*A�U�^Q�Wˎ��+�T��z�|`�m�:g!���Cj��xkik��f�%����wArG�Ur�o�K��&�6)���L*By��@�:�,_��N/8w%����*#�t��7��V����/�ei�h�^��[B�����^�au<]�xe'�5a�G&�[��X:7v������e�k���ۧ�e��M�H�K�D�
=Ð�A�tov�<��{dE �p=I�~���7|��'��pE�}���\æ���bzq�FF�"yJ�c;B�ul�k�uo��ׯ�)?�\���Y�#�Dj3�~��T�W����"�� E�Y���Ξ��˶��Hp�)�i��j�wqy�~Eq�k�y�����r������ԯk���0/�<�^�v���e�Jv=�ZNzU��{�E$�S�jT4UM��W8�Ck��ͧH�GxfQw0=�����=�٣m��,d\�Ld���ޝ
cU����lc�|���i�-!?Y*�C�c�9�Ef�^�͢�l<������_Wbrn3o����ۉ]��+�9�S�&�>�]���ĳ�]D���'z�����}Ἷ�6����[Q1�m��ɼsSc&����s{�.��<���kag�Se-�c��,��g,:��\�\��΅�ꡩ��~r���P���h�~5\�S=�ŵ��|-�CحR�j�SA{�*���b��]*֫������ ��%�E*��rm��b�92\躰��T�f����EW �%�F9HQ�SN�BN�.,�ғ'(�[����sɭ�L��N*��-���]8T)b����b�og'��A����לoT�;�}�|�5%�o�]�-)�k2Q�pYV/9&KY��*>u=��Q�B�ﻦ
Z4�m��y�o��k��>��^V��R��W޵�kl�,�"�j�.�o-�n�^_;	���Rs����M��{���w�	���H���z���u�gy�H�����[������Nx��o�y�	�n1�Ef�2�{t�5w6��Ǖ､[V��F��"��ť����j�VN�v
���<})W1���=�@w{�[��fvբ�<����VӨ�k{sΑ���"��e������p��s�u�L}C1TM��n�5.n�z�>y����\7
�N�&�^�h�|�j���;��M�.�<���fUX�o�aX��o���sӕ��ᝮ&�7���:���n�kޯ���:?)�*��h1�75Gk���la]N,-�לs��ư��Cj���/3SbR�r�R�/0�΍Pd^7ڒ�߳�r<N߬H�&�)aɱa�n`k�4��|���iו�%ե��,F!;Z`�Øu�$�R��X� �&�9ni�_}O�v�L>hܟ��M?5Xq�y���2�Z�{r�t9ݬ�]/(�{���&��χ�m�ܰ��c?b�&���#b�7���s�������:U~^n-=i��z���kG뵕A�,8py�R����T�j];۷o��y��qtj��6�����A�����*�򨒓��j��U8����9��:ʚI=���[�s�[pm(����*Qk'y�a"�(��єо�ZXoz�V;�O�����vDk�׌��R��X&��ŀ2�[�?o���Am�#ZY
�c�	w8�;׹	���8T�5SC�2^[�d[Zծ�ޙ.!���oL�٨���p,T��W&���8x1�z,���&�+�l�,��h\�[��y:��p��N�W*v�kC��������,�R��Cg�{ΨKG��\��|-+}<elܸ��3���"�z�8�#�k��EA4��1�(#���$���r�{��O	l��}x([��jh�dy���i3�����M'�Vrj�Ԩ�t-�|�͑|o)�f��a��y��ϊ;���6�Ԝ���Cҙ	�M���o��
3F+�s���Զ��:�'���&�����᧒KN<�=xq*�W��`���]��ҥd:�]�@�<�:9�7�b�֬B+�02�Qc���E� ��/������]>9���A��׶yTȑ\����t�f�nV��>��t�-�A��4�]���*u�pmA�2�!i�4@�Է>tV��ͻ��,�*Ŗ��2e<���]�9�Ó�:��K���ظ�LT78]uͤ*db�ᶅ(& ;����q�tw���yX�q��jz�G�ebN�3��
#n����|�r�w3{��Ӝ�IW\���H�5O���1�8�/�o&T�bnwo���̫HPΖ�!���8���Q����	mQ,�R|I��6�J�`V��p)�f�] ]Sm.���	!�Vnq����rsv��l�-TH)�]Ӱ^Cn�ai�gh�U��٠��0��%�����㌧M�i�;1�璮a�XgN�24h����'�u�#+����9�-��t9[�s�]���y�ȫ�;H���͂�mc(�	Ʊ\��&�t4B�nDn���/b/���Ihh�Դ�<1��GIV�nJ��`��rLRz3 �)�
�5�w�wr�f��BU�Vº�	�q8��CV��u���,4���h�(9qڅ%k�a�=Q[�z%��=]���|�d֤hA·��Y�0K���}�&����5�ި�LU(����M�5bz(63� ��ܸ-�p�mHU.ˀS�m�]�s9c���(���t���+*�]/Nj�>t��*�Q�ƆV�sp���,�t��;ˏ+�ň��ï:,���!k{'���.���U#h�i�bd��id�V�'�ujhA�A=/��T�wM�,����4itn���:�h�dsV���Gw)p6��j?��˽ņ�P#�:���/5>3u�������%m-;R­F��3h��[w6�f�sFlI�..:�v�+�%'Yu�Kʃ��9�V���$�;S�����w [�ؕoQ(!�S��]4򉂵��zKR��-$����UZᰕp�8�/�v���De��2	-
E}�Տ[����˹�8�¸��w�$�:t���������)�Ow0�k6 쮍-0f��q���+)�5�X)	C� ՀE���W;���������=�s-��#��3�b�Hs�U���-��4���V�ӣ+HD���A�;Z�\��C�oC�q����)6H�jc��+������)�:���s���E�Ks)�.�����tqɬGK:,Tt̂�飔z�=#��݊�hu
N�/-S�.	�Vv������M\:�~U h�R]�.��� P��JE���*$mf�H�J�X�	$)�D��L��"(��%D$B,@��KIm4��B (R�����-E�E���!!6�	��ET6�%�� �������@
��L"�DlXD��#l��l�d�"m$M�E�.��L�E2�,M��t�&�l���M)I �6ʈ�f��DX�M�������i�#,@� ��H�"6ȂM�a�mr��B (�*sI�i�lU�H��&��4�\�PP���!"""�D"�jRD��`����	��u�m�<�њ.�yı���8p�
���{W��5�,��[��3H��:6��U']em�|H�������|�/M.p��U���mT��bi��)��dO܇H���ѥ�<d�|���M}��<�;Iy���=[k\9���_7�Z��k�ME�W�;y�v�C�_����q���kj��)j���3�O�W��ߗ��	�I�~��~~g�(�����<����ݵ�+G��OՍ;S/���I,��y���m�GN�Z�V�5�ꬫ7\�`Ua��*L��R��/��V���0x>/����71N�{Ѳ���hvz�_r�s��c��una����)��O�x�sg4Tr��>v�_��v�t��ʤ�v�7��M�]��˒������h��3iz�[���o��i���=QH�_�ٰ������=jt�[zpr{E�����\5��8Z�y�i��WO%b���s�sx�4I�?�?I,�TC��PZy�����͎��&��x�"@'�s��p!^TL� ^ع�J�J,`�~�䏝��.�\;��9��B��/��	`��5s�Z���O�a�iwsc{�N�7�t�	0����ۘ�SarkE��dȻ&�;�p
:��fԌ�w�y��TMj��Ǧ�ū�H�B�G������Ԟ�S��yB���p՛���V�KE@�k0,��k��v��Q�r�j�,��Y��G�D)��)��KE�\��kwuQ�#��A���+����w�w����
m�W���)p�J���]�|���T�7����y���9M�j�����s~�(}˱����%]B��;ڸ�{K�u�M}�1-�������̪k�]�ժ|��z���w)>���*�i^�otN���$�z8sI�:���JJ�e��\��8�����[�؍�3��/'�~F���9|�m�i��j�i�����2i��o���OH;JZ�/�V�ϫV�R��>�J��4�3s{��!X�Q)���9�ڏ�ͨt��w�eq�Y�������d��;̕���?�؟�w
e?Z�oy������5����ڡ�Gҳ=e�cN�:�E�
ѣزc�P����D��`�B�B��>k���7mº��a*�7ז)�꺕C��RՑr,�[]�W<L�O��|�n��92�+ �օxVѥs��+I���&�,�<�����g��O�V���$��ԁNk�
���S���_?sb�t��J���vu�����V	���4�����\��聮��lU�o/����{�9�'�g/�����sT{���.�e	2�8p6k�Sa�Z[ˌp�@4ob��\�K���t����yŴ53f��۹��ڔY��,U<�)��O{Y��8ڎ{q�m|�T)J�:{��E|b������\�N�n�(	d�u��z�D������q�_<g)�2�S�wOł0�T���ؔ���0���s��B��S�=!��T`�����3�D��d8�N[9/�og
L OoMD��7P��Ts桾|���n;�z�f�Y<�z�g
���CnK�56�ky<|So�k�a�F�f���R�B;iHG[�S��"�9�V�sV�\�=�՝����^��b�]V�.�Q-��k�1�W�rru���0pT�iV;����9�C�,�ۗ ʻ�]z��"�\���5����s�ۄih\Ǘ��.�X��	VL�0BŌ$X���f�����èI 6�0�n�;���U�,H�f���6�0�g��^�^n5�3�cb�6 e�DK̨�ů�����VcW�9"�2�J��ͺ��k�/%Nl7�\��F��-�G�1
�o ���1����q��-�K�{�W״�ysq�dC�;��~Uf��C3���͞Lާ��=m�Ëj�zZ/�j��3͌�Z����{Æ:b��&�n���>�p�Ѭ�+�"nU[p�Y���y���>����}�.%���h�1��+��W���]ｺ��ׇup5_��"zT����H{���>`X�K59�3�������َ�9_Rf8�"K�U�U�DR�Uo���?7lg/W�����o�Z{poz�P�@l�A�y��r��w�z߫�Ə���,ÊG���8�jr�Il
=�� ۙu`�ݫ�aF5��?iZU��t�j���v���x�S����X	�X��c����T�m|6M;���)#8L�p�d[j�oV�d�KEm-8�V�f�&�^�r�cp:���
��o�ֆ_D�`Hj���k�2�������}��!/���C�8��*��sMms�J�1N�z8]��Y�(�\22��]7�!h���&ſ��;�^��o5�gT-}�[Jý{��h�(/��>SW���nQ@.���	�R�������Sm1�ʡG��)V�9�w£��t�|�=P
T4��D���MFЇ��Iasl��G%�.|�.1��dL)By�S�����{WaE��{I/].Ry��rw�O/[j��sPۍw�S����赽���&�%9��!���4v��ͧ�k�Պ�u�\9��cw8���vx<ʙ��v,z��/��M�U�C���8�m%D^�;����Z��}GNVN&+��CT���l��Ѧ�������՛�~°e�(��i�)��S��#6]<Ƶ���Ȃ��W�R�^L�ѧ���v����5X'����(3^��q-L�~�J�:��c"k��u�sά�;,u�s �W���E��10��\Kv����ڽCw$IT�f��8���<�Ӷ��=7�g�n?r�L��S=���+�&�6Ѵ�;-C3K�ͤ�ͱ�3�YM������ץs���bU�Eק�\;|!R��S¶�L{d$�����ۨ��D����lX��aj7oy��E(Y�������}K���EW�q�D�Zxwm,o7���Ƌ]��e�gm�\�����lU�o-6��zyY\ևE=��b��|ǉ�a7��9w�
�Zl���X���3�����^��ި���8GZ��:ȉu�WwO{utf1"�'��}0q���T�������%>�k4��̐���_�ժ���~��VY_y[�V߬�~�Uә���|�x���#N�_��G�ި���W�`�U1��ʥ�K��):m���^�b�gR�9��or�m����
��S�f��JW��c�n�o.�L~:τ鰇���������:��� ���*����s{u��ɱ��cey�����^�����o*\�o�y���c�Qt��fk^�c����\V��ŗ.���_��)��?I�͋�����w��n�+9~�P�w���3��B�n��j��
����I������l��;�>Z�t�;�S��s�u:JK4�`^�E:�:���t�1��#�G2���J�.���ع���o(��p�% �M6M�Q���r⎶t��\Vwn#���}��G4+j���ݩ�-�ګ1�ۧ�Qy�qǪ^���H@��%y��M�'T�m���n��N�,�IN��8�um��yq�ʶ��g5*Gv��:�S/.9�k>�Ck�{6�t��U_�W���W++~Ϋ�����j��E�w��4O4�}i��k�ɣ���e�:�4�]Zc��OU��,��^{}"c�1\���<�]�7�1������\������|z�{�y��*M�XΉ/d�����}�|jھTc;����xր��j��U��V3��"�io2u�S��o6��Pj�ojOl��|(t� ���$�;�����(}������Cy��5�-�y�_+J�P���}%A��E�5�ŉ3N��T�����N���O�|[��o������yr�c��M�7��4�N�����Ig9¥SO0��oz�h�N���(��iK7$��g�fy���k��B/�uyq`'�IE�¦o�	K�FJ�»;E8��3_q�D~�&X�G�mw,��'9���[]hm��{f������:�!D�I`(��n1z�ή̛g��|D��{���9P�r��1YK+���͞Ons��n9L��S���J~Y��Sj��p� �gQ��?^at6ޮ�Y{�u3?#�jj����5˶����#Z2���^Ug+/FsoT�:H�Y��P]�{�a�߷\~��~�(�T��q�3�W)���]SP��M�8G��Εo#W����rǎ�]��5�Q?�5F��'Xv���1Vu�u�\9x�l7�Q����E�S�F�����-޷ٕ;�6�S��u���sq�>���B��o�+�ǰeK�;˖ܗ��,�}'���Q1�;�2ظO_[u�Lb��CF��יF��'yln���gu������qo�=�mJƤ���%͘}ӆ��̊K[ܬv�Owm=��;,v�9�Ӳ�҆��Dy��h�+7C��L42����K��^BR1�� '�]�y)�.�N��25�v���Z�X���v������:j��:�+X��]ɦ}�އ /���ވ�.��I�����*�'������i����5xu�� +���Nq�AO���v�	�ow�'&u�ˍ)ޯ[}r�nv����0y�U���}�*\�ȽJ&��EQ́O�oi\iN��7i��Z{f�z�O܀�*+�:[ڝ؇�z���o���k�j�g
s�iz�����@ɿ^�f����ń|֮u�C�ju�T���e;��vF��o�VK:P�4��E2���8�=����a��W�y��}е�@o����T��Y)TnpM��Л9NA��|�_�P~F����9��w�H�уX�;�_T�>���J��h6�2���d�y?�N�0�v��{*4xeS��e}	s���÷�d"��!��򡏴Ӊ�Oc��}��g���2ץ��\o-��{2��M��adƺ"c���B�:8���)�~�ѣ=��|t�m��n��]X��T,p����M�,�xR�;ʶR�Iݔ�
���4���8�$V�]�R��*ei�(U�˙� $�*��%��N��6�5 �ڱ�gh�H��B�Km�Fu�F!��N�N�]�vt�(�.ౝ"�F.�q�+u���%�͵�҆�Cbnl�����ʳ��k'q�y�����w�^������wwT6Ӓ��y��*���p����T�ڈ��2�9�cOv��˙3�,[V�T$UM�����^<k�#L��N_qs���sN��UV��p.&-�"�!浧x�j�p���:�ɭ��_e��:­�w���͛���n/k��q�c::1��Z:��U���z���<���J�Q\>���NWRw��އP�Ҽ-���7�	�Żߍe��=O8-Om4�Vo)6� ������]]U7�Ἴp�k�~�g��E���flN�'5��zD�1�����q���N��|Zx�V�#'b�K�-U�rҸ�:�z��r�o��ex1��y����2�εs�G�e	}��ZeH��p��O5�6�*���������1�LY��"[���������ug�F�K�%����;�q�F�C��:G�~=�&�K�-v�3b��ԎSˎ���Z;�C�$]"sMYn���V�����,�PT�2�=��r4Ȇ�	+��X�kӛ�c"��D��o��Q+�]���Zu|��`άL���ha��&.
�';�A����W-s ��E��h���:u����ՙ��m�iY�7IGhڶ5K|�t6��4JI�OoF��^�v֪x�1�<�4"�]��o��e�H��l�������*wfv�Au*�7��T(7}w&�K�u�0���M
u�ѝ���q8D0�	$�rт��Ss8�k�����j�����\6�1G�eX�
�/V�.I��e6�,\a18�*���zz�u^���ᕿ��gݡha|��[�9F�ovV,�WL������k%��v�=�m��c���	��;fMw�m0�ԏ���W�':�N�����W|t�����Y�;-qK��57K�P�/!�wDiv�<�T�v�é
`;�U��f�b���w��mڤi3��|��� �Ao���}��'l'tMm��$"���7D���+�~�Xw۸.�Uz(�w+���r\S�u�:�g7m":x�QUvR��[��8ua�n����٩�J.����h�~�R
d�hgax����ٔ�����3a���w&M�{{0r��P%Ws#��|V(��F�f��="h�=������[k/>�eC}�6l-��V;�'J\�aC��m�:� &.�3,P4]���t'��%��x]O�������zP�Y�ǓB弭d;�oh��ƒ�ĭ���N�ɪ����)�۞'Nnp��f9\r�L9��L���g����d���3��������I(�۾�y؊e�,vZճ)�r�9�v ���Ʈ.N����H�}K������,�ozl�Z%�3n�m�.nS!�Q	� + �L���>�"MT�a�6�;��K$e�J�b�f`�5 ��QZ�� u�nv'��*U*�l\�f���l�k�{ZUʑmϑ�����O�f����"tA��&��,��ݜ1��k@	κ4�f��rLaP^>����I�K�e�8\F�tVnl<�v�[1�4�W`,q��lF���7E>�Uə�S�������� �8�����Un3��X��DV�W��fQ�ͥ@�N��`���-p���h��Z�u9Ef�|���Z���#2t<z�<����9CS9B$���޲}�g>��ͥ��ɤ��h�Y=�Z�N�¬(C�6�uW.[�Э��Lh
��B����P������qUծ%���ەb2���W��⑸��¥<�U-�dc(l�6�9v)መnB�{�D����U!%��ֲ�Ӌ@��V1�zM���-Ӻ#��e*ӻ(L����N��ч�����t�뻺Z�zM
X��M�Y� ���"DE"!b�B$B�$X�,(8¡@��5X�S4s`��H�H �.��E�� ��)�Q$�@*�)b���q� �
H�����)Z�$E�""�(")�!!Q�$EB"QRM9��Y�H�X�昰�7b4�Heͦ�ɈVI����&�Di��m�f�a NsI�6�F�H�� �͒b N9ˈ3m���2�XFػ�����̄@m�FM-ʙvL&F��h�8�"D6�l�T�UCi��&�l�mdf�^l�f6���&�-f�m�4��fM�\��V�P��'�M@�P�b�:"�am�y�Xm�iLJ�h��9J˯��Y1���fN�+4t�u,�;��l����{����#'5���y9y[��K{+�J���0T6�1�1Җ�\Ը|^��u��|�T�=Fbs��'Q��s�I�ٴ�9�]�����.�~�zE�u���?@ۘ=�jorj3y�a�}S_sLT6����c~����{�r^���#pg��=�'$�ԋ}�$�eY����� s�u*Zt�Kock�wU��;>��c��5�/6�fK���u~J'�D�&�u]��+��+l<�p\�C1aUQ�·��ξ-"U�΋m�Q{I�)����Y�mD{ٮQ�軒��0�*�~�v70�N��Zѐ:����cM�
k��k]�eY��wx�d���3����	3Dsډ��>��{���9]�j���l�j��f�繛ط�dx�V��ծ�)R;X�V�,�-�4"�K��x+�)����W3i��{AJ��3��V.�QF�l����EB�ึcl��۾������Ҥ�8������W���߱�D���1c�W�ֲU�q'S�ڡR�)��3�`R�L+Y/$�b7�u)���:��9�5�W�����	ϼ5e5�z��U��3�/\?E!�7;��;@=Z�����sˌkk��ۃ{b*���Q���d�F�{�Ͻb��t�W9��:�0�ys����p���u�R�}�T�2��u;S�[<-]6Q�/Փ�h���>USԻk��W�T�MIS�/���{�ή��.�xW�{��{Q���i_�޻O06͎�v�*V5[�V�X�޶��zd�FOF�[5���Y��56���F����x��~�����_%~��Y��2���?B�/a�)�J��<9`�<�7ҭ49��m����x\p�A[��� WI�h,��:{�du%��(*���mT�nz!����|�U[YOr�z��ګ�[ʗ���5�BW�o�}�{�+g\ru�\9O�o�a�[�
zq���X��+�Y^#JX��o���dF��͍��R���M���Q�d�s7}����ˌ��+i�r���U��C��� �{;�����d��2k|��ۑ�,�������"#!��y�J�*��bU7��.�$ű�V���,^�C�|"��f=q��s�)Ʊ�Z�Jx�>4����R�d.����3'������͊5��<�WH̓O*O1��&���l'�S��t����ڞc���W��C\tdstU���9�%���(�Ă�F;4�k(|{��t��>ݴ����;,v@U �TK����k$U���RW<���M�o�/�\޺oK�;��;l�Rd�c��o�ә�gZ���H%��\J�Qک_�[�p��m�Ĵ����PyN]�)6��<<�H*f�~��ҽVޜ�#p�,�~�:^�C��ƽ�����3�������bϽMۭ�n���%N���r�sƵ}�3x81woʈ^�lC����{5f�|�o�\��?Mw9��ν�����Uu�܉�V��6��V�z�=�_,g+� ���v	�ѽ=s���z�%�V�����6��X�nT�}g*K�w@MR�:���w1Β�"�յ�"��Sv��*���kRt�1��}Wn�`�:�Ec��QY'�6@.�)�0��C���V��׳R[�v�V뺈�|$�bv^�sk��� ���u*<�I	Q�7w�����jp�p�_6�3����ڰ���eWr�)*��_%)���V�9�P��Ts�)�}�wd"��?X�,
EXy:�G0M=�n����So��y�}���gy�PۍwkDq�.�bQ�$J���{�&��h�ٶ�v��]X��W�9m@�������zw�M�8H�?[ʽ��ZOk<��v=�M^�;���*��أow_���c�-�Oh[U<�f�T��߳�&ma�j��?v|T�����I��Z�F�Mz�<zr4΍4��7>�K#}��9Q�師��3M�@�7:��;߸�lgε�����s��򠫎0.��5{�sgVvˉ铻�1�F&6#�7n���dIoӞj��hŠY��i�r��}
�وuDI\*�k����n��6��yGU�;�@��E��n�FJ<��sZF�/�c*�A�7��Q\֒ζ!m��ݪW �I^t�R�YѨ�p P��_@�^L�vS5�Z�r�������Fӗt{��=5e������Z)a�R=\"j=���U�˔XK���jm��p�Q�FGx��rm}a�m���,����k7����R��+R݌���VlH������+�vRR�>�Od8Zz�9�C!zǓ���9�ҝ��Dk���!�o)��%
�=t���Kw�����*�8��.���o[�Z�7����N3^3z���;�鏋�`�;{U�ܽ�sj�`p��Wܷ�l��:֡݇�6�S�f�]D���u]�_o�V���G{zj'�=��������\��|�j�������g����B��l�U �r^����W���C}S\�M��!ޅ��q��p��q�l������2���{W��s�p�{n��_Ǫe�7����n�5����t2��Ƴ�����m��M&�a�f��e�X���r�iȶ�ބj�n�jҕ�6�!��뻩���'d;xVi��vH���}7�\
���Xfh�����WV1��j��6��J��ru�g]�4Y7+��f6c7��dfZ����P`�T�9�`g��g4`��t*�S�V�>S�Z��M��C�6�Ѩ��W��W&E��9��4��$�5v�<��K�֣=�3=��sY�m{ٮQ��3=<]��;�vW_*Xn뛜!�y�&+h�l*�^{��KW��&������n�=�t}���֕ͦ��]`��~�+)�<�ؿ��{�}ӑ'X�Ѯ����mg{�z���5BnXP籜R�ڵ���K��+���$[�v��5��򲹭b�?r*���u@V��R�Ŭ��˫��kg{/7���i����:y��PC���z��4�[S��;����]N��R�޸kn1�ڈy�l�U�LwϚՍ�T*mkV��CZU�c��c�ثķƋ}��Q�3j>��^���2Ɛ�p!	ӎz=�|7����Cy��}�_m�m+��^�{�;.��Gk2g^�:��VM���(�1�5#A��f�us��,T��Tri��������2���vK���2ٖO��@=�F�m�C��
zvо*�%�G��6�K����ݳ�S;nb"Dz�JB]�`�Pbʉ��wK4_:x,�h\�"[�\��*��\��Y[��N��/s��"t{
�b��ƕ��/"��$�ɣ�y����9����)�3��
Q���5ˑ�N{;���˗[�[��~��{�yt�6�6[�!M� �P:�ܓ�^��x��T]{ԡ�D�;Խ���v6'�q���DN���ӧ�ي��{l8����V>�Y�2���'������:�λ5���{ԏzS>*����*��I/��%:EJӢ⓮'�;��C�Up�ZwC���Z�٨YZ����G��,^vu���^auץx�2}��
�^OJ�7�]V��xt˫e/���&xgr�'�B�۽��m�ϻ����v���5Lx��eN��jm%��X�(�V(^�=Ϭ`�˙��4�
�a��n�|�ؼ;�v7]��ޫG*�'b�.�FЗ3�W�c�4,�w� ?V��v�;\X���=,�Z�^:�����g���Dٸ�\�9_L��Iק�(�c��8/Se��,�p�}){��=��v9��}�˃^s�>�g}/�<�+�gNx�(b���FEs�?�;��T�/�ۢ7Vyeƪ�jC?%�~���^K���^��\�ms�q47�Jl�k����qH�V�ơ�����g�.��]]�PT̜_T��6hroX]*(m������qJ����R���%3J$n�z���
(�5�$��әܳOp§s�~;�g���y/�I��YE��۫|�~��a�E���o�;�<���K�i	��+��޾0�.N���I�`H)(�������D�<���^K�I�F'�f�g�x^�%CF��}��!:mӨv-24���
! {�	��Y����ʢ���}5��V�9��/�T�=�8�[s���v�E�s=
y#�~b#�Oţ��9�iw1�j��yط\3'F���E��$]6��5�����m��3L���4ew�v�ޙ�r�<77�V�ﶎ�D�[f�؍M�y�"�k�rk�zK>���K����⸘��Y鹎���TԽ�ܥ�|�N����)���!5�f*}Ӹkٳ�h}��C���H���'�b-莑aw1�t_[�"��}�s~�TQ=N�#m�[�۟E���5��c����7���P�H=S��R��q��ovO���8�?\TW;�q2v~�!�B�B\ݕ���ѻN2(e]8��˖/'��γ꫹ct��a��f�{�����Z������گm?�ә��8�Oٜ0�����h�q�itx���D�����=�v�;����JQq	M�����QЭA���u��98V�`DF�V�Y9����������[���֎��fB���*��BΩl��i��Np*f��S"�!9Z�Z᛼�5�E��%������C>uU�'�9���un5�p�W9'/�������t5��g�Z靵SϢ�֎h��yŉJ�>���o�=*u�M�X����6}�|^L�^'=imv�{^�f��}�h��%є%\��qCՆӈ��/����u�Χ��	���zDy�X�{�G���>{�����׋�d�
��+���S�1Ǽ#�w��pb�×��g}����z'�Dڪw�y���⽤N�p4G�~^�4d�Y���v�5F�y����;�}���g��=���lhj�7���L{J�rx+�rQ�Y%�*�q]4�t���n�N����GW�ַ�;ⵉ`.��>��C���vz�{!�0�Q+>R ��K`7^ǣ�f����S�/ʻ�9�E��{"Ks�_ů3�o�j,�;t��5<T�JEe�X�o��9��qf{|U��N���E���Q�ʐ�~��dg_���vKnB�9�T<�гk>@�<��Ϳ/g�-��Q�"�T�N��9q�÷����\l2��e�\OY뜹��w7Yl���N�2��/��<��N_�����>���,L0Ǝ,��X�7	[y,7���O���K;v�5
��h ��Ց]�E�v�[2�H��.���	wr#�V�*5_>��Aۆj(V�����ޮLb}Aa�n���S�*[����Q���+%���U�Wг�H�\��ۊ��=�ޣ.#�Wt�]���V���u{�)N��T3�c�Q`y��A�,��C�}���Z�Vd��c�ҭ28Mn�b�e=�W7���]{�����>ϙʱx�T�����`��m	svK��A�:�܌���4g��XkŁ�v����]���@z�z�o�勎/fr��`�G%�5�9V�&���7���Z�U�hNN�8|b�heu�ҥ�؝e�w��������Ǎ�8^��j��Ҭ�8��笹d��@����NQ�T�d�B�`U�G�:���;����g��c�Wf�uo���+���o��,��^T��"�����^���6hJ�z-tF��ev�~`S�ߟ��^pY�-���i�s�v[y;{�XhQd��C�d���%�鸊�@72!Vo���Tc�ۜ��=o��f��X����Ì���nRQwK�8ef��Sӊ6��,���.�R�-w�N����P����������O����#hA�vutrbe���=���z�,��ia��
Nl,�t�NNgL�͂���DD�}���E�37s`�'f�a3;2�m�J�V
݆�X��x�mZ�Q���xT��Gm �(����xj؃fgm�;Υ�R"���c�z��M�,\⠝�j͚$��q) O���G,f�����mػ���(tsY�ꕔf�Ӻ����Sx0���!�����Ln����JΣ9T���_1͒�+��>v^��!o\���}��kA�3Wb�yo�&��e���(��T�;�4<�m[ܵ��ʲ+�Ň��Q*��p�&Q�8cO�O%<6%f�;j�[D;�WE��R��R��w���7g,(��5�D�#Xf��ם�>���.u��;Z1�9��IJ������p���;a�:ңW5���&�ly�`p�1�eϰћ�\S+;�Mӛ�S��s"�̕blQ֑k��}����IyP�`%U�̬�d��a�`���Dd-����+��T�QK�d��P�'G�P��P��*�u��Xz����8:1�*�A���=�8/)*�����E�zCz3�L��N���w�S&v�,8��{���]/d{�f�68�Byj#[�6�$+�oM']�B,��L��X�:�
]�k��E!�*T[���9h�嬾����c��=n�!`�'@N����[���U>��DiL�Y(���}�	�++��qEG7��uy;�g'{�RIl����?��Ao��9Ѿ1N5ͩW�Wp7�s��v�0�R�DsCQ6Z�����-��cy�%���V���D��Z+^�+.%�0H��ӑ��[Rjly�ѣ"��iY-�rԮ�5�܇��q�ث�ΰ1�R�g��i�۩w�"v�Z���q��i*�O�4z�����O���a�-u�]u��u� ܈N��?�#�2BxQ��C����@g���t�n3��Ζ��C���]]Z�[��w=����Sz�1byλ����b��\�����Bʶ�����lSG�9���n8�m�)���H}0quʐ6�
��{(���fGB�]E�vQa������܌��f%R&M�V�"�U2A��Er�{�ϗ1�����% �3��+`IM؜��Wg�q�z�!��C��纠2�w19VC�Z�C��I�J�}sP���>gf�v�n�ax�j�]>��j�h� .U9h�ә����ح�D|qnr���ߦ�B�\������H8�&�Z�T�G��^�b�5����`Wm�A�\���K��[�̨��g�\0v�Z�����˱J�2Rś�X́=�v�v*��v'X5}Kv�Q��꺰ք���{p�v����WA����*�d�3�{�9Q��Y7w��!Y���^R�(�����ZHo�E����ug,N	�$xi[o�*��V���c9d�P����=	i��#�(P�vrf�&L#A�"m�h���dD�X�m�$��!8�93beѐ��3!�e�44�t�Lm!16m4L��]8�Y�J���HXH5iLӛ�1s3i�M.Ni1��$q��v�&n&��M6h��V�bL)��3�B�My��@i��I�sy�h�6�S!���2�͹��l��]�h]DLմ�m��5�3SU���L��Mڢ�8��,�HͶ�k�ѩ�lЋ3M�	16٤єT.h�"�bm�k�Z��p��6�+m�6̩�i�ba.�d5�p�d�l�٦�6�m�M�i�	���J4�EnnR�+0�f44�&iDɑSk�I�bLM4k�c]��ʪm�m��f�3cK�M��$�k�u��u��t���+��c�f��qS	�h�p�qX�]�u�J��D�:�(��Q���De�b��q��)jo���[�;	_g/ѿ�e���wE�v��su�+���7��j�|����
��x|{'��mVr��x�GKFn1>=���|%��Tu�q��v�ՠ�����SQ�X�W�2{m�٘����E#�F��AQ{���_+��_Ͻhp�����}�~7�a�!����+�;ޣ�}�Jn�p�s�fK5���x��^��u���C�ƾ|���~�i�`�̙w���O��yΒ��5��h6��)��S�4��Ɓ�`�''�uv���=�f�B9�����9b������&���/��qo�GM�OL�+O�`����W��zh�8a�%VVU�3h��K�p���w����4:�2d��E��1#����qŽ[R4:����R�������'��߫WS��̞�@gU���3�oc����Y_{׶h���p�����\�gw������>���S�:%9�w��=g]�q�r��ñ�k]�!��,N��;Q�+�%<�<�*pޔN홅�;��W��s�殶 �������+c*f��
oڌah�g/��cw-i�k'�mZ�ḓ5,�q�;�����{�T"v��s�f4�	E��������W=J�̨g[͖��yj�;-���e�;Qs����Z1b�|:��Րm�y[�jR��6#'3��!a�*d�o���5fd̬>�^,�%?x���=�j3�w��ڹ�y
Y;�f�0�+*��/Įs�)���;���3�-;�� �/k�-�����u�[sÒ�Z���=qs�P�]���B�6�f26t^����z͝�W;ׅ�V#4���u�L�g�b�#_��CM�[-��Y>��^s��5�u5��|-Y�	B�S:�'��坎j;�\�>j~<�q��#���2}^�#�Y���!՛�tg�ܐ}Pe �|.*U/��Qf�v��s�xhQޏOE�[�㉘�[�b����͉Oٳ�r�f��>(2J�,	,줧#��_:~Ș�<��듾���ddz����=�|�0�Ŝv��t��� yQ�p&uĎ+���5E��ڎŶ�-�ݍ�K���tGRzoG9��}��ުbY%� �I�p69m��_�������<��f��E�͉_�]�����`���_�\E5�UC�%�pj[7\2v��>�w��6- �/�U���#�x)~7�B�W�z�����Y4�{�t�D��x��ќ&	]1�?q˺��
)F�n�֬����.�49����dF҂��x�"�{�H�eY���6�uշ�P��&�U�LS�l��Xy9�$����,�vy�s��ۛdH��F��cp詚�����,��&����c�vL� ��w"�4�a�g���C2�ڴz����|�p�j�;��C���H���49�#���Dv�(c�꼫�bC��QD�<OF]�}�*Z�ѕ������P�ކ1�]���\��F�:�}��.:})��ȃ���\TW�ʃ?bd�C��+�6��7f���/ov�d`�OdS���OHb��3�^.�����0��6q�������Z�n`�5�7r:��K�)�&���T*3w�u�'�x�쮦1�W��^��#����{�-\���Û/�����]��莯nɍY�BX���BR�'M��f����x����j��нz�ƛɝ�4� �	��{���sW[,�D�Bgä�:6��<�i��pX�:˂�s7��C3�fO��]o&�߽y��C})�����)Ǧ
��_JOM	Θ�ތsQ��˗<�N<��S���G�#��=~�跸m�s���� nzV��Qd��P�d��@J[�뮠��V��,�~��u�Š1�=gT�CPy��o���1�*rx+%x��
!�:����.����{��r)v8��'�/QMZݣu���I)�v^� %�b�:�B]7Y�0�;.�{�S��u��)��[$����ʳH;��>��H�S��b��*�D�:����K�p��*�6vact�x��Y�[3�ʻ�wb:�8�4"KW63Mv.n�C��4\��
��g�Z��=nb;{*.�S��U) yM}%��7|�
ˏ
:��)s�+����h>���Z�"�ߕ���n�f��:9���ܨ�����Ags�sǚ�k<=���Uǃ+�K��@�å����Σq�!��m��>ο3���[r��k�n�c��eW�̕I��u1�:H!54'KǴ9���T�^�q��oh�R���l:�ɫ������'����A=+�ʄ����"Wd�5>]��5t7�&:;0`N1��gz�S�ׇx�O�6�~�z|������,��Ga�_�O˲nϦֳ�y���e��_�2�v���*�ٔ��7�Rhu��s_s����>���r�ΦNȃ��4mz4d��4�T�+�o��__��s�u<5�WC}����1M:�n�_����ǬA���?m�-V�gw�%�m��v�
XW�e1��*��;�������J�d{[������ߪ�ú{<�?��p{��,�3b�̌����X�����j��n,	[,����D�V���%��/�]�G�5x�2�ț�b�Vcia�
�+޾�]:�bi}��˜�RpQ��vr� �1�j��_��:���m-�w��T��~}����q=�ys���I+�sQ�M �n��ֺ���;��b�/C��Ҝ�zӥ ;urڣ9=�6�[=b�"��6a֧.�y1���s��_sIY�,����ޑ	��ɭ7R�,�m0)k��"�O_�U�ym_^T<9��Oq�K�����t_ڲ���Y�)\���y^�F����~}�8������=����{�>X�8y�]l8�K#n��e.$ᐎ�P���yHC<��z=��x\�nuP�ar��[P˿}n�z����nx.�U
X$����^����^p�=Y��	Te�L������n�W7^һ�<_�ﳪ�3���l�x%���.~]'{� ��ނU��)����辕�tKs��s�����v�f<l�67��J4�+kۍO�{%����IG� e��,��9�t+}�C�D����w)�B�Ɩ{`Y>��~��k��Vk�.B�(���酄��d�}]-v�u�ԾQ��>���&��JV��t1�6�x�I~ף����E|��)��im*;�|qK�\�z��-�`���h��O�j���>5�����&�7;��qo�:n"@3ȩ�������c�..��=���D�-ȧ뭏{�\|�X���4�2�V ����i�1���)�߽f���޽bv\Mչ9[���h�;-M)ޘ z�W"����k��[O�#֪h��ݫ�Nu���Xw^!��/T��a�B	Z�j���Vٻ���OuN����cA$N���C�w�zuV���#�{����ה}3'GZ�L�����队��H�vnr�X}>���9ٹ�e�O&���6ԭ:'}��k��|n9��<��]�c�<!_�w�<�*��i�ne�Vf�-���v:(��sq�)ٸ[�	��c�3��xb�{�m�ө���껎����9�YV�⣦���<M���+�:��K�BWM��nWDF�8����h]w��m���*�F�s�)�:�{\�f��B��b,��a���*�䇹�ٸ#����i�lJ�~�%�����"�O7'!�F����H%�ڧd��콺���<��y��;q���,��W��x������e�&����u!�������;=����7�1���_J�)[�d�4�2@��5���9�ʇc����\�5�0˳﹦���}A�Fܐ㢃��U���bo�\����_�C&`��� 4XȩT�r-e]9�\�^=�0���B��<���ة�4燢�Y��[�3�ø%<I@�:H�_����_��c�`��r��x͈�y��J(W��l��cD^݊�X8/w/ש{#:>`�l6�+���3+�����k	$NbϺ��\��K��l�0����BW:����S�֤F"�@��K@��m=�:�Oy\��Jht�1�U1�5;_U�����FM{���l^e�ȹN��:���,㵢p�:u��f�D@�0�In��=+��ܘ
P��RK�J^�ei�B��<t&�{��zs���t;r���3Ч�<�1ܤ�`�d;��T̫���ҭ]���/Og���n!Q�����}9ų`���A�W�2��{�M�d����y�����a �N���v^����̼�Cٯiɮi�,���K����ٍ5���u^_v9W��CT���;�u`�X��>��5���5��Cofd�z���q��~���������U���9��r<$rtQ3��'��O�O˶���}^�y��[Wz�vK�ǎ��uU���%9��y0�P�A��늊�T�;1�;(B�#k�svV���;�B�zd{���c#Z�����=�t����0��6p7sQ[^��\M�F�@���QЉ�;�{���3j��r��6}���7���!�W��^�楪���{�.ϑ�b�6m��W�x<��yB�vN-�3ŀulmO�l�^��>��D����Z�'ϼV?;���Q���S,yZ3�z�wT�kN���`kܦ�������N��[J,\+���<P��2A��$>�Ul������D�@� ����kX:%&���J��e'��B�5�d�����.ka�N���;���6MʹV�};.�q��jl���ە������4�Z+�;�?�s����Íf;[P�FԮ�p�(z��mtF�}Nk�e�r��WQ^���Т�����,��͚b�������Vk�,�����H���T�ўrjz�=�pxz��0*�oW�1��0QM�|w��a��;����:��?�*��R;�PS��[��>�J|c�x�s
끝��_ٿ[���n�G#pE#�c�;e�{#��0�"�-�/#]u�h�O��:u@鯺�P��_�j,�1��w���t�`�*��<����j|y��w,Yy�9iV��|�Z�ƣ>�(�z�8^gp�5r��J-��9�|�+�>��b�j�7%^[Pt�1�el�I��nK�ct9�m�8�Sfg_�ߏ�@ߢ�y�"� �k�;��ʫ3�������H�c�"���fA�<�'��F�5l1R�����5�Ww)�V��㥴���2,D����+��H�ba��_W��VK]7�r�<���uHT)����L��o��\6���>����0	�<N\��~�?.ɻ683�`��f��m�M'o�&^M.�V��#��sy���]�r�@�<7Z��麦*�[�]�7��(��Y���I$��[�-'���@v<� ����͖kf�3�����.�޾���QCN�2a\dT,�������j��Zr�#�I�<�Α��ڢ�J����T�:s�q������GN�t�q�|�U��L��|J���ت��l������Y��\$����~���7�V��H�=�]]����c��&��H7A������wY�5�-CKkV/f�]�������6t;��cn�>'�wK��w�t��؝g�P9f�Ӧ��1G�s�^r�w���������NlL�z�·qS�t]J����`+�<��R�x�shgR3'�Fc��E�Y�nj3<1��.�*�,����ސ!==�)�R��i�}�U�n�'wW��}fC���-��9ﾞ�����N�{�Xj�% a��3���H�����j�#7勔g_8EY����Uw����y��\���W�7<7��R6��x��i`׽ ө��	~]!CX���=Fs��ʀY�|�xar��0�����N_K���ӑ� �;碮9�P7	���2���I�,�Q�#jR|�N�<zyLO��3�}mG��hvn;ͺ�]���t'.�mo;�������`)^3[,(ީ�\��:����~s�Y���	:V-���B]Z��w0J�@U��ܤ;�xD�]*��=W9��q<��*�RΡ�9�!�6%,�TH��y�Tw5G�g�;��/�հ̇��M	;�b�&�ͷ�q
��)s�J?�K|�fgY��;mG"�u�5��pE]�+휌�+���|��ۏU3��f�P@J��|[� q^s�9Э��᝛H�����1�p�%�+�T����S����N�f��
x��F��	�bbW���t�}��T�:OVԣyj�fW.�8�[{d`���la����z}M��E ��)�KhAQ�c	������:�hL,��o����IK]�+6Cfޔ<������`�3."-��鸉ߑO���7`�g`�EE��	����c�,��O���MO�����hv����UI�ֹ�&�s��GL�{'=�;��~�Ǔ~ΪH����A���������q@M�S��d�:��{��i�b\��s���T�iHexV>�}�B�9�ٶ}�p�q�*0�[�����N	Nt��]�*�eP�+���˅7^��i�T����ֺ��BʷW4��'��P�"�B}/	]7׼���C��(M�u�;�=��Dg{'!�˫eX�:�kSg���R��T��,����<5ʡ��
�u��+x�xu��Q}]�g��L��i )o��B����;���۞��нKQ��'�?���`�-_j���Q1���^����5��$C�dNIe,T��f\WÅ�dN�J����r�9�0뵜�q)Z�5w�;��O�{2ʱR��b@��hV���7>��%�	��XtĺKʹ��ma�'-ںY���$TάF�qt��z����MOSݠ�d� �%���HTdWF6��;n��VS�ܳM�E�'~��Y�cڸ�){�TZ�z�)V�mD�R'o](��ln��m�Dj,#z�G��Y�t�w
Z��-f�u�*�T;�7�Y�YB�T������Wq�MKf��9.��%�E{�NuʳC�2;8+��Hb���EY���: ����k��wpɯ>������vmx^mq���l�~��S�eB�hг1(�Hy��:��� 뷃T��U���z~�����f�V)ݔ�f���;K���(���O.W,����(^c*S�YW �']n�ʲ
{Ok�)���E�5Q��ZP��RU�[��Q|H�C�J+�D�)�Rl,��n��آӏ7#�:�v���.(��=ww�*�lL��vR="����v9��H̭�������{�@j���P�c����W"��)��7�j�\��N��w���3���9C]%�X��'�Ҥ�p�cẲ裫sd�s���r���ąЛ��	�R�#2�u�=|�=�}eRA|�jaY�\R�=��B�NV8qI���b��>�~8��4�<�^dDsU��u3�} ��q�Ĕ�NZ��N쎒�TQ�:F�x^N�`�T���+8��q]���3[g��7S����>�0�ٱ�1\���SV�Gz���-���׍Rt�����d᱗o��YKV�1MWnWH-��o]\{-��љ�����AWR��ۤ8��2ѵ��47S��^5P���j�1��+tg&Y _vڂp�RUz!���:�c[	M�v_S�BZ�K]5,Pම������0Mv��3�E҅�Dಅ�ӈ��(��C`��ia4ђT�`ZĄ�y+�(�,�vPr޵V4<9΃��P֖0�AvN �]��pp�v��(�K}� ���8��;�Fә�����(5��GZ�ŋ��U;�VnJ���0ĉ�ެ�T3*�>�r=Ъv����,�Cn�:@ A�)��m��jȌU�e!)njv�v] =�b��in�v*p�H��Ի�y��O�o[`-�qV+$�M����>�o2��v:B���%�e1�P��r�]�C��j,����	E�F�3
y.|�>�b�98dz��]�ANٳ�ۊ`=��fVeރx�Y��T*�nͽ�\�)M��5��h�ň�zi�r"�J{�脯�@�`v@̜�+���k7�:E���J΃�p��*�:k��bT1\��c6�P����{�'�`)|��&_*��2�BiI>��I!\�uAne`���m��F��٭(��w*Oe�Ư2t5f�Ôk���6N�256�*dvD��ai��"iʺ�@P�.�]��nsr$D�\E���1�BV�d�X-Ȋ��L�,1"@�̓	QrM����k���Jlͭ.�͓�kLV��&b�"m�M���bL���ɑWFMk�i6� 	�X�����3C$1�Fl��bhJfm�@�L�e&�VMP�]��.���f2\��FM�`�M�6�ăi4�mFa���6���K��m[T6�M�"���HƳ#]L��LX�Mm6̹� �kB@�2BB6ĘSH&k�Ą�0%qp �@^D��f���h�5�mj���D�db�&�m&K��Mmh"�cl�l�#5&�h$be͚�mt�d��	�C2$F6�m4A3+.X��I��B�j��q9�D.�D.���R��ml�i�D��Q� ����u���SQè��:�u�&iы���\�[w)�k�0_�f�ص��R�^���1Q������l�\+;TaH�<C�5�g�g�uq[T��J��G@{e�&��e���A����3<�/Td/y��P��Z�Nf��I�H�_�x*�	d:�����Y�c���.9�]�sM�ͷ�*�U���Ƿ����;Y^҇Y��rA�2��ȱ%J�赔Y�n�U���p�l��[����w-�b����Q��a1rQ�|ITe�"b���O���d��F�3v�^���(z^��������=~�BtۧP���`C�(p�{�	�
�f�^��C2}��E�v�b��]�hM��c��KӖ9�FNܨ�s=
~�-���U�aNk�8gڰھa�]��%�Z����-�:�F��i��8}9��;�Z6��)�2����4{�O�k�{=ȝ��5)���!W�*h��
_���B�h{NMi�,�旙,ە�!�@ڴ�����@{�^$0�H&<�@��_KX��	�N�f�a���C���I��Y4���|�VE�3%�����'E_"��0���0Z��8��mwS�BpJsC*]�zWQW�yZ�
��jA�eb�z;5 �	6h��uҥmr�O���(R#G�Wd��Q�ff
j�.Ôz�wmt]F��S��bF�v߱y
�z��b70oX<}�a�"X��(����ss;7\	`)R�:�4�x�A�{�xů�-^�]����jfNm��&*��N���̙�c��9U�i�������x�;1�;*�����bD�dVnL��n��z6��a�09�FEe�ӏk�z|;�3���p�w54�W���N��x�arHY�f$�������oaۼc�vo})m�g׫��쮧�e�:оŽ�!]__�+iy/>Ӆ>�����{��Ydݟ::ⲫH	����6�P~�S̲o�K�}Ϩn���L��|�}.�߶�|��˺/�k�8�������H�F�Ѹ�+��]���ֹ�\�O]{�G�ȯ{3��Q}�m�yC3æ�e%f��/h��L����Ѹ�tx;�aӅ�XkI�{6"A`^�����;E��0ܶw�\�<��{ܩ�v,�OT��FU1$�z��s���Y:�L�ܼ�˨ްk��T�������;�����Ǹ�<|.J5�,���8	5���Ԇ��uVgT��}��t�/N1N�\��8�v|5�|���#�ӽ�n��`�*�����g{�dQ�Xz�*�w�RB�*@���/\��W���M�n�f��:5qە�J~D��9������W�F�(���ѓY����Wo�k�ڞ�(���d�.׊�+�/TS8��Dȫ�|9�l��OWr��"�5+���Z*�Ly���]Z��5g䎗w2Q]�bW5/�Z�/�7��a��ƍ���-�0���|B���E%���ec�/o�I�3�Y���3��?D�\q~,b��Q|�b�9�!�����z���,���jS���{��[�%�t�s,���:���0�G^�����r��NoiEʖ�3������r��t	�Y6�^�ƣ`S����+�ʄ����"Wd�5>]���~�4] �{�T���U{a�xg�[{D1�yULW��Y/�CN"��|����2���ޠ:pm�;� z�T��8�g�W�t�̡�k9�8o��޷15ΜF�>���r�����D�w~5���جs�9��=�0�yZ��mn�����m��O�\^�@t}������c{25
�l�j�{��U���-m\d.���:��\Z��M��\�eu�.�����=��b������'oQ`��O����3����ۉ��6t;�����U~'qu0*/|�<-K����M�(�'.�g�NK�N3����^�W^�f��'twȰ����u.��@�Gw�͗�����oZ�.b��J�}ծ�|�y�ϩ����AF���v|JVfza���{�t�U����bE��eN�ܢ�@q�>s�jU�G��j�׼!�86z���c�<����)U���w�������k)��5l%�m�ΐs(N ��am�v��hb�}N>4S���mKt~�q�ϯ��R�[g��_C[ܶd7e4�t�j��IEl�s��ݷn+s06�_Q���,�p���a�x/ND��*F�\�Orމ`U3H_zϯP�7|�+dz���S�Dk���{�g��2���7�>N/W�#}^�`#r0���^W�����D��O4�!F�R�rq�[Rx��騚�O�ơ���j8��c��D���x&6�f�j�r��4���� ֙`O�J�-�5�犏_�
������G6\[�ݹ��Xw���E��n��g��$���
����8�9ж/|AK��.^Gl����ͧ/�N2��0�nB����S�3�wL,$%�rM�i�.�U+��8�y�נz�U��a-?;c�:K�q-���<�Kk�*;�Ϯ���wY�$�[��!���P�^H�����Ⱥ��ry��_|̸���鸊uNL��gjj���{.�<Ic�e�`^�Y�q5��[9G4���(?��KҼMy���)�{蒠Fo��kk3�8�gԑ�8⿏�FT5�ꕶn.+__��wS�}����~�FW~Q]0?-�ı�f}u��	SkRon��p�mo��4�Z�Um9BWk���Wx�YO��P���Ǫԭ�v�9&��n��h�θ�jz �[�
�Gj�5	����˕om�Z*����VU���Ł��JO!�r�њ�R�z��3x�w&Γqi}��0�~D~�ߖYZ���?F����<�mE��P��E�u��wS�e�{�Zx:j$��~ǻ7�:���;����k\�L+�n�*(�J�g��������Y7ՙVQ���N_�+'g�{޴ �n���][*�9�{Z��9�'b��*=�������,ə���m�{���lK�8hJZ�X6� ��ݑq
�����WN6��?=���l����-�%Z������io��zvgJ��>:&#�˖MkYyo�;�{C2�}/z�O�̞Y}���s��.*�p�	����(Nt��]�j;�\�5�0˳�c1m�?��7����_~�<�ڝ`���	F��A�,	ȱT�^9�Z�,�;sQ2�FZ3���A�W��FK��>./�[���<
�#����id���\�"�줧��Ќuo�4n�w�yd��4ë�D�.�W�r����b�W��ai�t����B"�|f+�]uK:܃�Փ����d�˰��t��_v=�4��lx�/N_9��h;r����.$��?Lƹ��U���$F�ز��w*�KӑK��;hɗٱX@�������*8"\)[e<������6®���BB����3~������m��G{p�EzY����YTT/*S�g2�ݷ�aG���=�qh!��rIwi�,������c6e�Μ�|��MoV0s⤉�V�R/Q���*7y�q�װ�l�n�\D�����ur���{�W�x�%6�9ƾVq�qA7;S��r0i�y�ċײ�����YW=p���Y�/��@�4����)W~��k�~,]<��o'?Cc9ʇ�B��7�F�̊�;P��+����r\���d�m1�#�xN'E����2a���a����g�Z��o�Ip�-ޫck<'��E����xg�����m8��5�⢾�r��d�ǐ쯡]�Yxy��hG�k��H�q�^��?��J��o�_���oo���#�>�Y���ǽ�b�^T�������˥N�w4<�_5}�)�|[�W�e4d�i8wT���w��S�9�Fv��A{/�������٨�z�r�-�:�Y���w��u\:�L٠N�tג�����J�e�:X���Zz jP���x�Ab�~�絈�4�L�^'l�Bg���}GD�#�z�F�pg>�]
Z���S9�MA�[�ܽ���Z�VvT鿬�|����b�g��s������E)��:��	���s,^o��z��]��W��/��j�%�=�z��"f�b�(�`�m�3���)�`�;������i�*�s���2��M�������R �*�І��9o7�Ul�d-j-�WT
N���vm<�����L<�*�'Lc���N������}�[;����5�X�ʔh2Oi�~4eS<�q���oaz��ozu�ҁ�6��z�F�a6o���vW��C��呵�R:v8��x1a� n3��fj���K= E)�Ǯ��i��_'����j,����5�R6�S��[��S�{�'��$�� Jk�(	��x-���ƣ���(�;�Ak���Y�cd�z�}>�mM�>����)�Q�PB*�]2�p7�����/�����1w=�n2-O".�s�[>�����WdַA[I��3��uFI���S�N���7�9�!^~��պW�뜎��oh�����fE�����J�r�!����"S���u��.��d��/��ޫ�mͮ]��qA���������4�-������Y=�!���ꄎ�u?=���������{2�Ü�\ho���[�����8�/Ï���ܨ4ݮ�#��.�����:�;}$����*�4&�����]����o��V��1M}�n���Q׻�Zh}������)��t17�yW�8Ke.fDmj(���tb�k.暞��	��Ÿss��*���(�����L���ok�8l�P4�*����f�z�oR�睺�!��3yժh]��\!�݈JB��B�-u5&"�h��T�	n�%�+�哗
|
5'�F�n|1}J�Ǹ��]A�t�vF߶�N��R�]DM\W^�Y��~���(~�W���ToK6��N?:�z��t]5��	ܮ��9b"|+h�����[e[�et�q����3�����5�����(w��мU�z�`��=*Լ��kG|��Es�F�O2�����qrػ-����J�B�'v�<��Z�£ǅOe��~�e�.+j�����UW��"��7=����Ë��"w=*,�v�� �rE%�:���M��2V��t��b�����g�jw�t��}.19Po�f���������R�'�&P��$�>��7�V+��i]�/�-���x�U�J�G%K�4o�������A�e�6
4���_`L+�lt�Xޕ�t:s�31\]�z�ϕ����0˘�o�i��c�ߜ��KH�"��:F�C=،Qů��k������Uŝ����ئ�S��|����~�q��s	�n��_9r��3�wL,${�z���Y���q�Y��1��m-�έl�<m�t���J{&�0c�n��N��~���?b63ƭ%�V�+O1�z'�n�c�6N�JR��N�U��3�ۨߜ<f��]�U{�g���P�
+������9	��M�7��W���0^Je6�Ic'�2"�g�h�}����u�,#B~t�>�"}�=87�z�
���\KK|��Z������i�ݧy�\Y�a'��hN�5��f�o����������^ o� :�%�
�É���	�I�ΟT�g�@�����M�ПN��}��|3�P~�f�ֲh��C�9*����4��NxLz�1�}�q� �l`f��J�7
�%�]����t:n=^Cd��WWo!����7�\�����I�~*��d�ǐ�7R��I����>�^_� Ndy�}��F��3�wK���5���P����E}��^5g���x�͹R3������b���%\��elDO�o�ǇL��W5��51v^<���ң�5q7b���PNP��ڵ���^J��%'��L_bn�Ry�+�u�q�H,�{�}�5o�F�+��]_o:�t@�d����U��T.4�
��O2��S	r�P��V�_��oc�}Z����y�Wը���0NG`���Bs�*�j;�\�'�����W��S���3�B�h��P;��ed]N�C������BzQ�^���vJW
��x*�"�o4U�ѵ+�[�
��Ni(�=��vb��G|��J;O���}Q�N����b����ʈ�m��x�m�U�4y�э�)�-��ǅ%�#-��G��r���5�Ɯ�ZhW#$��@"�Ԫ^9k(���:�yTd�X��J��;�m�ldxg=�sr��<W�(�r�%W�X
D�uW��)͏z����/=�O�u �u?dLPO�\xk�|v��1g(;��g�!�I�Lzu�fQ�Vg���~� r�'��"�`t��C��	���c��^����FNܨ��B�pv-"�vnJ��GS�3�b
�&|끱����Q���*6�?[g�8��O����g�:��~U���}`~�猲Ih�Ƨ�#�/ԅ]*h����y����{NN\gl�s��+��է,�'Ki{	c��8�&7�<qH)�Հ��47��K�򗤯A��Ѹ/���I��ۙ�w:2h����<$btQ3��ɏ!�C�O�J�4�*,�Nq1��ܟ�i󞌯�j�:<s���:�ÕA��W�_�*(c�Pg'f<�e0��cW���\3F��#��\�x{lnӌ�˫��xzڎ3��z��l�QV o��L)3U2d;��1�ËWp���'�M�U��!e(�15rP��L��ڊܲ��o�NZ��Vؽ� ��=[��7�U�S5Z��'5N�.�c�>
�sWdeᚳ"��i+l����/��$i�(ۖ�P�j�Mi��w�(��<7�3��"L�������t*���W·a��]��
u
G�N���Üx�d��VF�i���+~N����_�˟��ymK��B�����H�ۘ�T��&u�w�ي����yu����9��ԩJaZmp�X��绸�����n+bm
�#
ދ��Z۽�J�ĵs���}��pӬ
�
FVy�3mh:��3<+�X��Ґ�X*�"Ӆivl^����CP�0^�kE^ ꚦ�{���̀��T\�+�W���F���$�]a]������7�s+2��I1�uډl���b�qȪN�h�cb��Z��wSQ;�Q�IJ�ǁ;�/\��Y>0��
���s�.ٍՃY	ԉ�ɯ��8S��w��ҸͣI�����@ة&f ��dn��]!��*0Z�v�h��n�A���^�0]���چ�Q��͞�O�̑YH]`���(S�4���U�%�Q��V0�W�p�֚���Pmlֲ����>�[�s��_c�a7.��i찤Ye	�!�WK�M�ûCY��tn�J��4��݅�T����R(	a�0V�PY6ԮU͚[8���_9t뉊�i����e��tЏhb�� �r�9%�%��W{���Iv�*&_i��wJk��(�S���[���a4b]�NٔJ����䫞;�,��N1�tU�ޤ�yRt[�kL��Ie�z��;1b��٨��:�9��ّIe0wl�ɵ�e1'����͛)��Z�����N�R�C\M�����V0�����VX�{WR+��������z� ��A�d駔�P���w��M��LB��Q&it���T�{:�	�-E�Q�i�i��*�)t��! <���`�D�8����r��p3U�M��n�.f^b]�l�r��]A���2ۗ���یCp�m�}��]����60�N�K{�I���(�M�ɧ:���ͣ��t�S�/<�`gʐzVh�9(�9�e�5J�a����PZ�^�Ɖ���i��ִ˰�tJ�gV�<9��5K��6��0m�/��4���4�s�k�5����e�)i��p:&�5�^'�j}���0��-�\���o�OS�H�q���)D��K��C4٘��ŏ��De�3/���Q���U��2
R���*;j4�$ebr[�b8$��zݔ�i:XƟ�V�똚�� ��s/r��Z��%��Zpv᱆pŝ�V�*>�w���[�-��e�}��f@*�W�9MR��諨�ήJL@�N��^��fe����H��<BU����.��n�p�Ha��As�Oy�H�l!9����tk�I�6"����Ci��L�3!DY���m�U(E6�R�f�2�����6�F�A���F��]�	�m����j��;Mm	R#� T��K[H�$m�.�Q(R�m1ˉP�6�r�D�� �	��#���] M�&�jDT2h���&�T�ڶ(����6��I�D&��	4ڢ��f�jxӛ8¡G6�*-9�I9���q18�b	��B��9�m��3�೛�^m&M��m5�F�m)BH�"�٪��D$6���B&��r^)I9�8�h�Q�h2dB͚�R"f ���m3&�@Bf���t'6M����Uf�HZB�$�"���H�8� F�b���["Bd�R,�T �m6�H��i"sj�&�Yt,�"B�		���m�0H�D@ ���
 �@U e�ɓ��ܮh���������-��FJb�lKp;W'wt�V�#"0Uh��Md�G ��r|��'�	p��#���{39v!�=K���@,b7�ݨw�ђ^��~.3�ߣ�t̻'�k���ö�+�X�30x�R�V:{���ژ]'{O67�ߎ,��سq�|y\uO�pД�����������S̲M.�}�)�׹�s�v|����W��ג����f��=0�FД��UK��8vX\A��/ĭ�%=�}@��wK��S������7�{)+6(�>@�y �.�|�޽�wo)��dKP��C%�F��^qG��j;�z\�0���M��s���{��=+L�r���뚄x:����%BX���s���u�k}P7�[��`�}�[�����x|��ڊGL�{��U�˩ܟc��N���@�H��_��Y�O(M��� �#�{} =+�j�K��G�t�Ρ��\�uoS��Q7� �,	ׁ�-��騽>OhM�n�����Gs3��'T��<;�szMŸ��7J.��+���A��}DL�\��~,n�:���Hw��p�j�Y��_r�\z�LǠ���6j�܅�e��26P��"bJ�I������%�]��
����]����h����|i2��Y��@��*u&6T��DL+���D ���Ʈ�י�P)��������iM���)���2�)�[��a�}�̷Z��Ӿ��m�D��;���Fr��5� �Vi�ۂ�q;��j�p���Fz���{�����1��VY�i{��dX��A{�+����x��cӚ���-^]Q�ؽ���,}-vb����1��{U1C_K%�q�C����K'���1�����޾�(�,���lM���(v�)Ǜ�6���~����9V{l��g�U��v��m�T�Af�^�pvp+�[�������BR��ݷ���/� z���0^��:H��﷑���������^�\
#F·u��J��";���g[����a��\����'r�V�eψ7�u�������^��ZY�tq�~�WBW��#��>��Oi캂�!~��o5Z�.b3�t2L��n�����}��H��J�Zx�� �ޑ	��I�힆L��e���/���꜠7�m *�ߌǾ��N�O3������ء{�Xh
,�ؿ�K",�s�U���,�Qӳ(�r�<�UW��"��7=���=���q��D;�&%����U����SQ�K�,�9���$���<k���xar��چ]ې�/5sq;[�j��R��M'�,VWD�%�p��B$�0h}{�]7��Ѷ��4(Օܩ-����f�.�WV.n8�����+R.I�ZƋ�H�ɻ�Gaw]1�S���tλa��,T\E�v�C45�Frk�^V�{��Ǧ]#��ٮ�`n<�j=��ML����s�q�X6O�K���`O�ʡ�T�sᖮ�.�Э����mΜQu��A�󳷫���p�ac��r���5ǄL8"!�|e��Ϡt�Xϵ�o�glo��>;?M��M��i��)�у��z�;�z�n��g��G��1��Q3݈�}Nߍy�赭n����^{���W_v:���o����e8��9�ӷAYi��q��" 6�#�1�J�*��^��J�ɏKu�n"�Z/�:�o���?*C�z����p6��)��C�P�5HH�ګ�W��{�=���L̿|�Dq ��QT���f��{�|d]�&�7;��qn�W���n�W�W�%�׳΀s.L�����e���/�E]e/��r����(?7�R{���T�[4�G{{9�I����c�X��#8�R��T5���T��~��?����b%�ҫw??���v��:��1��ZG�c�<!^���|}�p��+�d�W��O��ڪGS~�/|ln����>s������ƴ����5���jW��⣦����7tP׳��f�u1,�'ޘ��2�g�1;%d0��n*����ʏ�h�,�Mi2P��]l��ڼ�f.Uu�i5�J��ϕ��}J����2��H4��J���:��'KOJ����)o�PwDeY�E��_Z/-(C��,b�����$�r��uG��H����q>{.�Vʱ�w���X�9�/o*FH��&'C!^HTZ�#Y�k��K~�1�j
�B��*��/ĮL��#��T�r]Lb��� ��a�!�
��׎�����:��E�-'b�$�d�������\!����u.|M�J��{v�bV4]�{����`�7����u��������NJ[D%��)=Ag(<�ژ���r���!����:����19�ڢ�x��l�����5�=�Q�rA�,	�"��R�x��:+�!>x%�����͟z��U��ÆGz�_��q��C�y������; ���a���xg3b��x��=�L>��t��1_'ή<5ܾ;�G���aY��^Y���Y=?b�v��^��S�]���*D�>e��Q��Ws�,C~��/�s��ӷ*-ן�qQ��n�[0��;}Y�>�>�L�� �2GKu����@u��B�m?[dx�x���>6uڵ��*���;�����y�<�������DĿRR��Х�߹	�{�*���K6҃����9��W���byR��*�WKF�L����yy�S�Mc����%-71Vȕ{��ި�@���KV�Y��Y��{�#�U�-e�����]d�;z�ܾIѭg	��*��@B���J{�	W!�U�,En��Nܘ��G����'��߉��
sL��= �^_�.{ƅ�c���r�T_[��u)�5�b�Q�c�oj���Ό�m1�#�xH��v8����vP����>�����Ow�����+=���*\o>��j�c��w:��naʯ�i��~�����&N��	nׅ{�rq����E�;7f��]���q�C.��kI��������4��F��,+�;U8�}[U��-F��lG��ٻ�����K��>��s5쮧��e�:о�v�qn�r��{�vΖ0���]K���'���j��>��BR�N�'�f��T���SU}ԉ��Y^�ð佣�[�����]^���y+�Z6n�K��!,���97���z�^Y��>��z=��o�
V���x�����j�w�֣�S��|��2�T<Xuw��^T��>/Ezu��sw�Ft�w��pb��\_�9l;<W���nzV���s��BQ�����/�r�Ƴ�2���v��Ck}P7Ëuq�a6o���v7=Ή�੏A�&|��h��+חN�fO\(�@v��N�D>IA��=p�����,s��R�ZF��p���Jρ�0��z!�{��܎i�q^��(�V��捾J¶�"�/ 70���L�u*t���\_m���/TC�l�/N0��"I]Ӌ�����)�&?��$삆�GvGP�S�zzdu��_'���kP�g����7/r"s���W�W�+�Sޑ�e�l�T) 55%�!��7���]X�qߕ�\O�i|iKC�5{;o/gѽrk��Pv�E�jx�&8��UO����1����9�A�0ҕP��%^��;e=�i�k#������۠��s,��O�;�2Lת�Yk4����(���n;*��g����y�b������g���'��2,D�t�#J�r�$5��'��o���'o3��콢
�nJ�ݵY�l�7�&k{U1��%�z#����������X�7�_�s?}�=��N��t�����̡�s�ˍo����s�_s�����`S�} ���k����S�d�>�>%T����W^��u�������Y	��>��
�eMNͼ^A6�R��m�`��r�\��t�Q��K
�·q�Ქ�:z;����y����(��|8x�$���8��򩥦�Ox��ڠ������CK6��q�b��W�W��H�WkM���1��#���q�$B�ܲRu�/����7[r�&�����s�}hm�QG{?CRt}��_��w�j��0"���������Wg���szQ6u��fm�i�]�Pp�l�zs���[���lj8Uq3��}�c�E�?0<�s�}�rX렿�N3�nj3=�:��� ��	h��r��e����nP���՞\hz)Mq�������)k���uk���og�c0�7��B�Ұ���q���c����U{����(g��-R�Wz�o uP�q[�/�s޹��8����ˌ0"�ЎE�7�9�n^��C�>��t.$�|d�:�����\ ���ۅ˳�mC.��v�օN��X0o�wO��*c�r�+�%T)�$�,�yT;����"��f�v��M�R���f���gW�KDqz}���U��3����*2���x��:[=�ֆ6������Y>x#����ź�q4���ǵ��x�Y�v�+�3�uE#�F�� ��	��Ԍ�?�WN�ʲ�-�+zr���z���;`z��5s�K�!x��9r�(�Y�n�5�͋��K}��']��	<�K�t�_��k�|���~v�A�����{ӂ�h�%C�F�۾X��	���� ��G3��W��)h��+��w��ۆ�95���o�T�B�S�{�!�j�x���wF�$6�.�iGʟ�5�悒S|���������N׍��{�Kb:9loHq��k�]����<÷�ӛ(��u�W4��;��1f������X�4% ���a�\js� .s��X�*�b�w�B[���o�sB�� s��hꜙ���xW�e��8*}�o~2�}9z����U�A�����ۮŕ�y�%̗�i�2hnb1�<؃�H�U������`���i�=��3��+��N	�%�A9��eCm�q|In�YM�Ѭ.���d�;6.n9�eq�g�ӭ�z�f�ݧ�}�y8Nf'�ʫ��/<=�c�ֺ�٨Y~�7�yS��K't>�٧غ�j��7k\��H��};���nWDDվ��Vʱ�u�֦.�c���7R��XH���hN���nZj5��w@��BSج��$��m0&�'Z���j��u:ݦ��ǣ�m��<�g������;'��%%���B��R7].�����O�Į��c���fo�3���ɯ0�C����;���/#qUȓ��s	du})=Ag(<�@�O2F
�d��p_�{&�q��rv�e��_�8�;�p7�~G��7nH<�Ȱv�c�\`9������fR�u�}~�<n6�j&��8��0�����9A�����3(�r�%x�9^{	�óe��	��&�[�ph���t��]Ah������9�W%|oi��|��x�Ť��\ݬX���Í^Eu+ �մ:V�[w��ҷT��Hy�e$��S*v���]���gy%�@��3����hK
�#'Q��,�w���i
1� 
��:1,��
D����n��.�&0'ή=�����1g)��+5��:W3�;N����^��>(� .��ӄ�g��:E�����o}��_������q75>}��g���MU�^SW��Z�?��Hꟴ�C�%�	wNAyb�Q�|�F�~��9 ��s�Ve��ۺ��ozM�e��[����*yI-%���&%����T���K���n+�k�Sw�wu(c���l�m=%�~'�:�)�2E"�H&�V
�=�1>��>��j�ޏr̷�{����>r��ݮL:�T�_k�FM����<'��d�=a�vJ�����0�w	���;+��Ը�wSp�ކ3��w1_u��*�4�P�늊�T��ܫ0pf{�Z^���I/��5bwL;�SvV�����N2(e�Ӎi<;������,6��tt�7�ӗ{n�3��zTz��M�C�F�GP�zQ=d����n3�߆C��i=���^��VU�B�7R���-�Ay�w��^G�\X=�júʮ2J�(�.DC�3F����"�pO[[a-��eԖp;���(Mn ����d���]�ͤge��Ce�tޕ�`��˻��4��X�Sc�h7��(����z5+�z�����μtN<�Q'�Y�hY\��q�h5CM�cMф��=
U�s�vf�O���G#4ƣ����ͥwy��ʶ)��N��n�3��Ff�uzhY�%q��_�tzaOu>��w|=6�#�Z�;^%%\�1|�Ŭ�ڋ�pk�s��>u<�z{hfs��6��a�d��]5��<�,�̨�/޵�$v5���q��J�/ w�����pb��\_��-��;=�^�'sҴ�x]����e�Yu�>$�(^������M	ʐv���T����-�u������qpG�����{5<�����#fF�$�#�Q{#�Ѹ�P,�y"q>�gY����_�W�ůl{.y�X��|��F۪a�6J� )���&u�lt�^k��C�+����c�e/�N�F�m�̖��yz��ُ�n�]5,�C��PB*�}DLKu���~,j�M^X��26sѳ������,7��<���!�K�ū�h6�+�2ʎ$�����C�����uXu����R+�y4=-�i��à�h�ֽ����Yd���2,GO �4�����WLɂ���7�N����Q\䚟.�U�#�v+!���W��2^,�U���#�m�Ւ�e���I-���Y-�K-����d�ۤ��,���-�K-���m��o�d��,���-�K-����d����-�K-����d���,��,��%��e�Im�Ym�d��,�����%���e��e��,��,���-�K-���m��o�$��,��Im�Ym���
�2���Rq �� ���9�>�.���Zҥ�J�%Z�QE���J���Ud�*�M�R+kj"�Y�Cت(��I Z�EV�"�I*�leMQcU2�Z�e����J+j�l�-Y��5�����f��Ҵ�,��j�mL��6�,֍�-��2�Ѷ�kU�뮳���Xmi��حk����۹��Vk��j��L&�m���ږ6���T���Ŷ�5���e���U�kIF��j͋J�cm�fٚ��d6X�5�E�R�1��Zֶ���a�   ��o|�q���۶Ӛ:����ݽ��zouv�vU{�{;�ηmn�\j�ǎp��opn�Rl����^�׶���UW��wt�����ڴڭ�6��fm�m���  ��_T>��E�w�Wk֞�s�ѽ*�QEs�c��(��(�}�=� ��(�P㾽�Q@Q{��ƅQEQF}SQ@ QEξ��(�(��7=���щ��m�lX&��  w{�QA��0UUv����=j�)��AT��s�=uY{�eڨh9��tk���ʸ��P��7:5CCۭ�X��sˢ�֊̛*�����[S_   ׆��hAj�Jw�⧶����m���q�:�(Sn�����l��r�n������Mv����gK��m�֣�N����ך�ӷqN�t0�dֶ�M[#U�l��  o�m[O�t����m5lU��l�ot���ڝ�6����k�(�ٓv�۹u.k���^��vv�G=�{ww:��^�]�wv���u�ջ���w�ڋ�;t��Qfm#�K-��@k>  �����Wk�ܧz��7Z�v�;�]�mgs*�r]�z�^滵U�<.��V�֛][�knʻ;�wN��wi㇮UW�]ڬ�9��T���%��W;��87�����kVmU�h�5���  ��^�ꖢ��p�v�@�=u��i�׼;�Sm����u�zu�:�0q��]v����^�ܥ��ն���kT����ݼ�zJ����N�'�nܺ��ɚi�U�l�٪�M�j�I_  ���>����{ۺλ�:�w�����U��u�J����F���ݕ�oOi�����s3�+�����kW�/{�j����*�{���9w�G�������^�]���w]e��ٶ�Z0��  ���W޵V�j����-��wk���;خ�Yk����:V����u����7^��zٵm�=5�n�+]�w6�ݶ��wmZۡΫLڹgn��3{�u]���<�3f��6��i�RK-U�6�   m|/�wk�3N'*�j��wnwܽ{�OKf������3�۲ۯ;ޭ{l�YnT:��:�4-J��X6��cީ�ˮͷkn�3�{��گ<뽫w)���eIJ� )�)JJ  CB)��J�A�  "��	R�  �~BfUT� � �J��*�@ ѓ�S������`����~��r��?��\�W�g�9�NW���k[���y���_�	!I��	!I��HHhB���IO�H@�!! ���|��Q�?���}������Ckw��%�ȋ]|���U@�����X�Ȩ'J�!m9f��S�X)}����)��ĥ�2Q��>��1a;��An��2;������#����0��g�7t�ӀGt��[)+��ګr��P��R6���Р;���O�O	�#UF��}tb�m�$��W_�����&�����N�X�0w�r��75[ݔh�eqZ�/%�mٛ臽���3	|�D�f��u��Z*��v4�n�-Ճ���䑨�-=�rC��,��B8΅�l�LJ��k3t�D����Să���,�e1m�jũ�yV_O$Z-��8��=]��G�`ur'Y����E�ͤZ�s2��MQ���5i"a�
�y�0؃���+�ë�ΨFj���/1ZNoVݶn;��
�:(ϵ�tY1��Z`�\փ&��2�^�hVբ>a v�j�#��Gh�t����@*��
��-�NQ5y�siyo��i�)xܱ�,�t��Ys)X8�V�1;]�L0z��<sSU��lSF�JM�f���/�1Kf�֘ǩ}-�t#�n�z�,dt�Z�7��C7Z
����}Fm�	
�ڳ7JEF:�-ef[�7�,c���L�a�v�[O�&-�z��r#���"��oJ!
O8r�t�φ�L�4�E,Y�ʗ�E�HLoA�h,T���X���P�
;ܬ_]Fsv��56Z��rə��{���f�kE�o��xn�]��7`�>�9�G���Y�3srm�j���l0iH����"��JRIm�&��%4j�d�iǁ �\wz(	t�tH+A��{�G�Z_�qz�7�P�����PՑj�HKC����o��M��L�����)BO�	��L�����kM:n�M�:�C(]Պ�׋M~�DC�o�ZV��yL�JX���V�k^�V
b+G�k[�y�	v^u�f�U���HTLи����a!Vk���i�D��)ШE�tH�YU�仾I�DŁ]L(7}`�6�Ͼ��A��Ƥ&\.��b�<���}�Ǡ,7�A�W��x�v�K:P:1�Z�e����O�=��M� �Ʀy]ͭ�a�%,/c�N������OqS�,I�~��~���E��<�B}A�$1z��h1��6��O�N��'�V�^#�����pV���t\� `�Q����OMͩA|�7�ڜ���4LAQ5\��t'.LD�� h�5c���}�6�/H��+)A,i����ʕ����/+V�+-Zwzt��#2�e�9v`F�E���tўݠ��A
�	���h�e����h�y0q<MݶY=�{���%8�W�[�4<2�D����R�C�����K���;���30�Y�ӭ�ö�;�}b�c��lq�v^�#����Q):8��&-n�ꬬ��Ҕӡ���s��-}7ry-��"^#��:	�7�,�샵��ECM����|*�L�7'Q�<Õ���-��`����̢�t0f*.�Z�����7A�BD���˲��4��=��E��V�諂���Pdݔ�XFe�Ә�$��^ޜQqY���8G��|�5,�0�}��AG�&��V��e�l��ܻ�%���A65]e��O��6 ɷa�����1i[kOp˾�$�n8L.�ОZf�E��3+��->� [�F��*ȵWYxH�6�GW[Of��D�dU�I�EY��ih���Ho,0��[�VKl^n]G��gU1��Z/j�LU��7�q
JV�n5�uh���na~ۇѐ�5�=]܃�Z�R9��r�ZwS��}5XO�܏�6���R�
A�FnY�ǖ���뀙2��^Cn��X��.�4�Րc8Aӹ��/O
5:0�gn�L`zߩ���D���֎#��f�Z���7��@M�ȼ5.�+Q �BSHa$�y��qx@�)�Kb��c�uT���^ɞ-e��̒E�֐n�
)�e	�!�����\�.�͏��$P7� ����m��j'�X�C[h�CqX���wW� ��"�j7���S%>�%��;��3��ғ�1L~��Izj�@2��c�Vu���Ʉ�u��v� B���x(l��#hL%�2��ئ�wI9@f�\�;�Q��Q/['f�~�)n=�">��Jp���g��k��r,�h&�PB����'n�wh	7f;zՆF逺B��3��S�𣉜3v�W����'�/�L/�K��0�N�f]���[N��"�u���}����o�7H�-óaz�hel���l���͸�,b��NƍKf?H���(,�z��W&��_)N�����9U�ۍ�]��?L���VƻB���j'7 ����'�x詊Hv�-k�j��@::^ҋ%�f8��Z��A�&ZXp�M�
���Ͱ������H��f��׫��Q`�x��ļ�j�Fweÿ#�/ؑ@�8��uz�[�-e&6�����o���H�n�ڹu\{�-0ma\�r���<����5U{�%8t����"h��to�Y��{G�<�����\���.�T7捎.�"E�&�Y�g^]�l7�i'q�h�S���ph')m�vV��{)�f�[cO��F�׋�E�ė0�5���K\<B�Y���ь��.�C��'���q$���f~��^���r�#�U�}o�P��B��nE� ��DX�QG�ea@�˹u�ag���=��p�?��+97^n�PF:u����}�ax����_���iZ�#�Y�t!�Dߕ/f�f��9ba�wEi������B��$ZF<��х<tA�'�{)$��P��{S;A �u2옝	-;eY��^�ʷ}pd���Lmc� K�ݸ��jd[�`ߘ�����264���� -��Z�J����+�e��ݬVq��Ƭڵ@�r�O	�G�l�k"��{B��TT�����Cq��
$^SY>�I%�����.E6ki��H×{��ȴ�򋒳b
X5�L=I�Si��v�8��4ZޗΧ����ZLe-Փ*	�D��\�����Z}Vy�U]e��(5z����|�J�F�H Zk7b�K�,�6n�m�����ŏ�|&"e��4Q��ccW�(G^^�;/�^�K� W�Y�_5��q@v66;���`1�o�Zw��C<�-Zb03�GvÞ�y�K�j囎c��qM+4#�ڠ��)朤(=u�;4T�aհ���T%�E̘v�PAn�9��Ԕ#âj��*��g��i���\cm�,~�l7g��U7d<mbE��{+#��{�v:��P������37wIԷZ��*�@��ꖡ���E���ʏ�^>���y����=EP�TU���Cd5��n϶㬛�o.U�J`b�J�,���A���T��`�#��kɚ��Zj�"h@��";}�rx�f���܈R�YDX��paR���w�v}-\�e�!Y�v{l7���>�r�+Yj���t<��I�G��7V}3�uTâ`p��,ת��8����D��7�O���WwUtk_�	�]�VLB�2�͖��]I�Q�W���GQÎ��zM�hR��4K8��'B��gnX��ףe;�#��
�p���N�W��Cl�v��@gPOr������Ҳ��i �L�,�q]�ڹvE�l��͂�c5L7*���_����g%�P�6?��M�H�l��*�'��%��!�F��Ѡmt�(�3��Zl�'����֭#r'\��gfg�8PN�(��b�0"��(�33PuI��u�6h�|��kKi����IU��g�q19=�X}r�&Tږ��l���B�A���i͒�حӉ<&�"����ud��-.���agou���i�u�H]v���X%K"���$��ڄŸrLS��������y��q�tV#\�sEҰ��)kݤBc>l�%b����+T�/�.::TW���w�;X5U�*� 2:{W�Qj���D5������K.4n��	VX=t
��{wts~.����!+U�%i:Ľ�+A3d*��Mxے�
ͫ�%�H�7�A�Uҕ0¨�"'���z��R
�6��i%�|�8�r�u-��W�P�|�UMx��� � Ԝ�����6x��?��C���ZL��ef���f�<��&L���τ}r����iW��e�9��	�-y��	VqӍV�aЋ%�l7�轅<:�n�V�Y,GQ�j�������*������T��f{�'�Q�R�Tmk��}�D,f�Ѷ�c�l�IE3u�M�#�Bi�{e@a�F�(-+�l�t���H��r6���e:��N�FCS�&�捸5���M����TȲ�^ZP�����4�a5d��k��]��	bi�u]YB�r�[����늷l�E�bg\fckt�6^Aqb7�J�J H���зT5���n�Ѽg��
�uq��a���������R6!"��b=dV�E$��.aպt��mA�e�=���aHh�9gg�]�^�	��B��S���+����Si�"9ö�Z�e��Z�%�
��H 0���;fJC�]tH�����VVǖ��@��Co���t��JV9��07im*\F���Hr�T1*�sī�O�x6���6ߢ��򈑍�e?!0�7iMG�����9�,�S��gd��b��Y}�g�u�T����ܡjJ�\\+էR�o!�4�kbfjADoP<��
ۃ\��pe%	g���u���z���*� ��u��Y�2�U��ވ(�էNFT�FOd��<�7ѧ��v�׹�+�r|G�U+.9m�9��
1\�[�RmӎP��[v���8�'�x�p�����92;I�}�֝K�c�ί2���1'j9�q��~Z�;�cwW�bb�<g��VN9}q@�[�ٲLڟ���:����:�5���hX%�K���Î���Fkq���2mo֮��T:F�E���f3R�1�/V�{�' �aˁf*�\�(Q�GXM�8�d
	�;�=��I��75Ş�}7F�F;p��[6;��h^L��F'��	�G����Ǹrb22�:[�3�
��X�C1�F���Л�KÉ�8��*��c�*f��~W��K����B��oPm��Ў���fS��%j<���=s���0x����{J�Y��t���]f�;�s�<���ق@���^���LQ*��
u�,�ϝ];͔�ŧY�`Y�`����q&�[��	�na=t�L� �&���)����pV���7h��8�5��@�D�#����S]B��uui�Qn�ۄ�(��	�f�K��Ҙ�[Z�����v�����f����}���\�He�y���oջ��ɎO]/'���V(Q��mQ��]kt50�d�M�{�E�Hc��'�=y%��g��w��\;�Q�3�A�`�V��jCYZ�Uա�J��b��_���S_�"��"=���}f% f�=Q�_�a�����@;�����P(�"�neYB�P�7p�HP��)�C�9��:����]�<�	�{��F&�푼q^j���E�J�Rʼ��z5��n�y�L�	[W�6��-��U���3mh�}�����"��s3�d��у�h����c�����	�gj�K"n�W�i&,ۀJ�J�j��mڄ����K���(3�Tǎˤ���!T��e��x�:�l�7���r��("7�\��8�|0�o����|1S��eM
]�IA�_z%�.G�0�=��&���ӗG�)� C�I<�oI�UR� 
s&�C٧{�&h�3O��}�f3�a�jѸ+�ې�Gp?(�Z�ٿ8uj�h;��*޴N
J�M��iVV�^�[�΂]=X�i�Ƿ����*d�f��k;Ӱ�\{`��4)����ԖM�6���w}�^��-�lQ�nŞ��H7�e��>�fnY��@@(e;ņӡ��B7Suh���`l���p�Z��*f�7�br-ї� �Ə��>Ï#����}�����|q�� �i�3����$x<��f����0b(����0����dB4�mc�)�2b���n�Wj��❰�!�M,�Ƿ��}a���f=f�;Z�z�,a�7L���N�����1tݼyH,m֨�%p��a�d�)��a~�ںF���z�#��m��Y�U([UpM1�Uo����C�=634#�A[2��+�i�c��'�e�=hc�6�Zٴ囷B͖���J�(#uN�c�)e�إ�7.X>k)�kCһ�\8"�23VX+&]����	�a3�y+T����B(#<���� E;X��u&	A׺uˏ�5�L	�~�}%�%�O<��	~���*5�b�����stF�*��o
U��eX�ͶN&��I���$���˞��Ѹ.��7ʲ�)�g^ $I��}�Bb<�W�<\)�-��{�m������$���Z�u�2&��	�P�sMK`���B;ZL������AU���+
d6��Be�SҚ٘H�����S�B�[/\���W\U�v�2�X�{U%�� ��%A��	����_vx�������1[��Ρ��l��g��od
�۔K��[ח*wbR7;�'�m̧�DWXջC*�ST�����O�t���ƚ�2���v�ED�?{˾ʦ�ޕ; ���@���yyf�Gg@��]6�d��:�K$h,��8�h���3�L�le=��
�����5ض�..�إ	ظ�d��݆n��y��VJ�r]f5�Q#2���6&M�H�Ӊ��dKڕ��)\rI���t^� ,5Ӵ^b?/eBJ婍7b�S@��q�c��;��D�b=rlj���OvG˺�zò���Bљq�@������Q��1��	BwE���KY�K���%��n�u�p_�ε�����	��Y�v��n{�<�E׆ ���eJ�;�*g5!Ya� �������������LBt���z-]n�f�^�+&�!����[�م2B<�u�]�_<ru図[�u�O����v��.��PȻ��Ȁ�q�eZswS��h�a��:�_��.\���{G�8�e>�_�S�h8 ��f/<v�7d3]�S��p�x}�"*�v3Y� ��J`᦯�}ң�V��^_�u_Z:���=A=���O�X|=�',ʶ�[�b�Ծ�f9��@�ə�	j.SJ�ĳ�x��c54�s �qA��0�M`��6I������[`l5m���
I?'���G�H|n篯��`(r
iK�X�^ͺ��ɀOv���V0#}@�N�{ګ>��a��5+>�&�F׮�dY������Z��`X����%>�|F��~�\�ַ�|3���֜�Yj�]����_V+Dt>,�C"��2�@�������^�9��NU|��[�-�����������`���잕�!�q�`^��G����]k�\+O� �NU�\ѯ�=�<q��a���~��ޙ��
�NU��w�R��!��p���U�ͩ,� ���t�7���Ɵ6�B>e<T#,��ypT�������'�cŽvnPD����Q]eMW�YO�vd��/�L[�c:iI��]�����������}�L��d�������9��`���m[��ۨT�l�kr�od���]]�E^�ԍ ���E����a�8���WvQ�z����+�%}�r�y�T��u����'�sۭi*=#��8)(�S�}b��1�:N�����X�������<�2)��"�&n1���v7k2ŋ���/7ݫW;8����I�A�V}�(.C�-���~D;�s}|�a��]����*�zۍ���i�X�1��ޚc+ĹI���Z��2��p�`�:@� $��E�}&�G����)hKC�]L�f�؆�i�x���{�����t[�3�j�|�E�.��=:V��1�$�n��w|�'}mXȷ�狄�36H>y��e$nmi�2�Jo��o�$�Xi����Tu�0���{��,�{��'>ZQ;A��t�|5qjZ�y�/]]�g�W�N�:{H�+�3�=,[�kܜ�͡i��au7�V���k>�iT�����9��l_=�ۛ�DQ%��u�5�j��E�����x��*�/!Af���휋+���l��|���pE���J�sr ��ӱ`����;�T��
u�ﷳ�+Xp-N�+����Yv6��s�S@�G��l�gʄR��';!
��Tw��
�f��B���a ��}����8��pe��}�U�HW���;��pU�Jn�IH��J�o� ��5�T7�ࡥԜ˞��@	\DïW�|4S��|=��9(�oCZwt�2��֗&��]}dp\��̑r���yȲ��e]R����K��}��vr�n�[���vK"X�h���8����<��)�1tPZ�b��j�F����Q���){y��yH�(P4���Za�*�X�oJݽ�I�R��QN�+�W�=仗������&����ÈF���'��c5APZ�e��U�ƙ�ip�9�_pp��sR�1�k
���11��fc����}�u l�9%�����%t:��yZ'��]u�@�	��_3�E�����Z�?f�;�� ����߼��v�r��:7Xs:J�\X춪J��kSμ	�6�n�tèg*5����EkS{gnʚ�v��L[]
j�
�l��7*NPW���Mゆ�"���/%�����1Z�dI�����6�Q� �K\]ɵ۴
��f���8��g�J0H�k��p�,#.�G�X|ƪ��t�{�*� xu-�F�l�V/%����'r{.&�4�o}�ċ����#��xo�͡�.�Q;�Y����V�'�҇��|�X�P
���t�2u��5�n��H��c�=���m�k%�rܼu�v����YЎ1�x7�+E�{���uyWI�´��Ǫ�=�|5M������7H�x�=c8
���*���:Y_��q͓Mx����eK���C3PQ!��P�mi+��=�V�'�+b<E+�H^⽅hT��-��}�d�}�k�#�{�M�E[t�Ju�q6���ڡ*Àc��:{nQ��Ӻ6Oe��3�Z:_8�t�Ό�nh�'�tf.��[J���zR,�n��cu���O�:[��s�뛑��M�c/�T��nfv���Z,Jz�S�Uɵff��Ղ�sT���q���Tq�]~Kq>���
7s�Y������z��O�>����UCȡ��s������$�z���.��e\�5�ް�dΏ!��D^[x��Z����U�TuPӺ'�nK�`ͺo \�C%�Gf�'��漾s+M1^5�k�lۿ<{LL�F��+"BYa�͚�@�Y��e�N�mt}H���P���<
u�HgK�.<�7u�؂W����{q �h�y����D��y� V���w��qv��M:f�R������Xy�R�Ce�q��YiK��d���A%��dZ�[�~O3M�N!:�v���}M1�{�y�#$K�x)G�C���yw������z̜����^ӤhU�N0�k�83Z�6�6q�̿n�۞F�RʾA�/N>��;};X�oj 7sq��Ȋ�0�1��eH8�}���H��y�����v�����;U�j{w�s�o���um�v��=�42Tܟ\���([��]Ƭ�4�덄%�BӒ���v&�f��)cv���
�u7y�� y��f\2�y/� �yp��r�\��J�R����`�����|*3��y�=�G_ǵ �WFkF6� ��Mo�J��R�|�� K��GQ%W��J��a�L05��[�T�aw�У+�=����J�+�&��룗$Ґ�:�^�t���� �K9*�h�ꁟ@�Ñ��,&r����=�w!<��@����J���ϥ/ �E(�Z�-m�g�ᡚ��ȷ��
��9>�)�0��Y�m����7q,�Gv<� \֞�R���S��&� �}�=��Q�]mY)�D��u�8���1z�,峵7>���{Wm9NI�/�h6*�4]����܏�yR\�9M�t�K����H�4QX�aB� Ո�*�:t+���ļ.�6n�d�V�U^��CYt8]d�����a�����R�QL:����QR�u#v6F|�bʃ�rm�X�7��v��4o�y� m�!��!�w�.�";][�j��\�3c�tA.��y��3��;81�������ylggr�
L�G,Z
k�i��V�0�W���e�ˋHn�o��k]&+9�	�(�1ԹDr�Cyw�fuZ[1Gt;r8� �͚w��E��
.�N[���
��V��Z����R�QS������0^E��fe`j�ߣ�jX�ߵޑ|ԐQ�+̂����!��hPS�.��c����"#�Lf��9��Y�������l�7���xk�-����'$gr�S9e!43�Ȉ�J:��u�.��
Bv�ܗ/\T�fj����U�q�:�;ĲS�<7P��);�6�v+�*		�ŉ���ы%�`ߨ
�|��Fs����x�ڏxc� f�G&ɣ��=���;���E�U2���;$�&�i�٧-�@U`���M/Q��dV�U����WI�%E�d❛/��)A��Z�WS2��ގe�V�:����:ʨ*È2�X&;^���7s}�M�P:�
��^�6m�,W R-�R�Fլ0���sj�V��Y�s�8��f�ұGf}��dLв:��s�x�#�*���)�kz}�Z 	��w&0GN�u����;�dѵ���E�vru���I�@�����!}\y�\K75aξy �ה�'k��^�� -�|P^��")1�t+�&:%��x�P����_X���n.8*�r���E��Iޙ��nf�u׽@�o8[/GK�Ŋ�ۂ90���6/ ݡ 8z�JZ� ����_md<w�����ɣ2`w1�PM�o��7q!�;f�}� �a��p˅�t�Џ
�����s5t��iQ�p8{d]�NH����eL�2�݀�)��1��	�Tpv��&n��z�����w?i:\T�A��r�^%�gP���{BؒVb��gY�Ȕ&���f¤���:or�Ph᪮�MX�b�h>}������_�6.�9��{l�� ���z���9�Q��O3��1:I���,>�����V����˲��Z�Y��ʼ�y��f.J���MI�K��tTN���V*�f��X�V(�/Jכ�D�x�gP���0T��j�Y0.��zN��x���da(�-Cmm�t	���<̛o��LU�3�[R���B�;]��Yq�U����2j��L�������=�$`�Ԃ�����'P���6�>�;��6�6��D[��lE�S��t/c�ߤj��!+m��AǄ�鸴����R�ż�xњuާ���{��=yO�<iCr��C��b���y;�>L�\q��2t�w^Q���V;�2=ѷ�9=���uL�mۧ�s%�E�ƹ�U��B35�b�iC'�r�v����ૐ�$�4݂�+}$ܗ�a���Xk^��i庳۾6�s�Y:��W1He ��ŗ��6��� ��*�a�ǵ�O'�~<�)}��ZL�ъe.�豛��8�	G���[�d��kն�����%�������O,���6��Y`�
QЕڮ�o}�E�a�GA|Bݞ&���l��VV"ʱZ}Y6�W"żZ��V`M�P�A�x:r.�����y���'�ص�m��B.�D��u�o	��2���5�Jv�k.N��@�r��X�A��e6��˥�x)M 0�A�:s��3��z�N(�H�U�Z.{6wg3�t��91���X�:0��ʩ�ca9�����чl芡(�XUK]>#���ǯ\L�΂��3eaڃ�o�K��fdTxu��AR�V1���5de���\�hX�G�j'��$��%�57��e�AJ���gc������
&+k;D$#B�<��%�c����	��v����ט�V�A�9���]�� ��%��	&pJ�y ht֮.����<�o&��K� O6`К��Pj5ʊ�]�80�7�dK��jޤ���0BH�BmwҞ�=`@ۅ�T#&����rSZ0<x,Ѕe�}m�DZ�wEgY�ҾUpmv�c��gK�S���Kα�[�)����e�%2��G��k����1*���|�ҭ���<��N� ����03�j'�̔��vqz��ݏ��t�'I�|�:��6�5�N�`����u!�wW�eo���xe7��<4#��E8�Ű���X� {�m����1����Q��2���0��+rtA��&��,�=�E�-2oH���)F�c� �c�{V$��[���K=�3^���]h9(r�Ʊ��fX���Lk��o�R�e��t�K�yW:C��������zӛ}"9!����V�c�mN/���5)<����T��`��%<�^^�q8` `����7��u��a��Co�r�zlMI]9�Y�p-U(��&��u��3+w
�@�	'���ɱ��-�
-�v&�U��ם�(�t�A�����<�׶|��ZLr��uݠ������)�����n�]]��3��>�3��wl}���W$W
9� u{ո�Bv/�^d�S��VYw���Y����.�r�-��i�o%�=5����#���Ǵ���n��E���e�_I�v�5}R�if�*�u�[����13BP�4˩lvR<k��e���C��X�n!{)q�I1����lu�rI�k��Aoby�o��/Y�7�L��酏ee�sm�x��=������]�Ǉ�}$E7c�?����M�xv�Ij5�QF�
�6�{�j���/x1��a"�@�;H��hkX��S�5��\�f���Ã��V��>�pڶ�u��_}���:N�އ1��52UJ�w~�w�C}�?�RC[��l�'sR���j,yQe����[:�<��7B���8�>/y�Kg����<�>NK�f�*x�t���⠙�$�S����x  �w�ڹ@u��\�5����zh�s:VR7�u�b���ԛ2���d��0���;���˵Zz�.���w5k`\qo&�A�\��|�.|\��ټWZ�9`{�ô�����E۵��B2�R��#��!�xq���wkb[�6�d�w�!�JgBy��æH��8��������2b��5(�˗x����������)�Cb��7��U����	!I������Sy�y�߽=��b@(f�JZ�����u	�k{��Ú��C��C��i�~zQ��>4�i�L�ӳ��tr��k{-A��7s+�nka�.��H�H���]��6�z�-52]���7���t��˝�$ç�i~Uۥb������q�bϣ�ʗT]���8lº�eϏB�A��uoT�n��ulח57���vFU67�HNm�]|��j���L�et`S�˳l�)Y��6�u�O7���Q��Q[�%��v
��L��L�C_v.^��7ۚ�@c(�A�4J�Vl�ڻuK=�²Vs�y`�=Ef݋9s����B�l��Ǖ��^�w���j���1:�=5EܦPy78�C�0"w}��ǝ�ӕnl���c8b����R�WCK�Cr���<G�ò]�P�:׹�!#0��T��2��!��.��.�����V�*H7F�y�`��;��V���:����˞���G��rΓ��,�g�>�,,{�HU9o�SI��w	�FSa֋ܗB���{����#�{<�\|�4�vi! �`];�2y�G�%�]�/��R�}X ����@i5�'WqZ����5�U���gl�+gͱ�Y6�Y������2�`g��ݞw���f����饃����[�N��p�<:^�������%ц������%j���'NSUTz&ϩ�a�Q�1���ڮ
�)W3^�୘l���]������A�)b��3��Q��I��	�WJ�)�oᠶ/����s2��=ƌ�p�eni�Z�Z�!���u'���{���ϣ�d�gC���=P}h��+��YWE\�څ(7zlhw��#�[yդ*B�3$��W�:��.���#g°!�M]ֳ�bF�n��d���|(�0�Bp -*�KBV���W,QV��UASR�9eX�낎��P:����,{`�5������KZ.��L�YOd�K�9;8�9/6��^;�b
�ܻ-!ŭ]�p\�%���g=���ߺ�����;��@���}��V��Y�;GI�o���K�a��}�H�NL��nӬ�}e<�a �;:�Y�X��a������9�yo&��G����#M5n:�_�{"h�Ɖ��'��	��9ɧ��J���l���'���u�=v��5l����C��{�(T�E��瑞��϶�m����մ��lf]�*6,��u��.��3/4R<�8WQ��̗�{��0��^ �X@�)oGJ���i���I�E[��d�P��%��1�k�a�8���E\�j�V��	i|�<�[�֭���c�)AU���JӃ(�vyr>�^'��"���x�H�膙u��i\ط{������˱�dܶ���=wٰ�M�a.��^q���)S��&�,*��f�w(��4�h�	:�}F�:WJ�`�Tn�jur�+����(�@���%�$q��N}��L�cri��;w���!a�]�X�b��
t�e�^F����u��0�3�fh\����d�.���2�n�i�*�-U�V{t�^ �N)KBD�G�O�����#�� ��O�sz\�iys�f9�X�q�V,�>k�&��$�`F`���d(���}�6�/��>��hvf<ۻ1e��f4��!��Nca�U׊9��%i�'h����5�Ok�a]A��^����b�a���o'wlp^�1�����l�$�r�C8��(��W�d�4�a<�/j�e*�;�E����b�07�+}2���p�i-_nPI1[��ܙV�\8�����ۓkBg���i+��ʱ˞�����6�:^���r�*N��=��԰iK>��$(i��r�kc�[CP6�TN�U��s;�X�Џn��Cm�嶒�)�T�-�z��ttc�?Ch�pM���2���wx��0a5|�MWC�A�pTu&.�@$U��E�Pt��ϲ�XQ0ܺ	qOH�nܞ���ꦼg���`ީ��;�c�]���.��o����n'ډf�<A���#��1$E�����̌*��_et�a�A��f�|��h+B���L�j��h+�v[\��;4�)�6,#�]���<�׼Kz�81(��8��gt��5{Q��ql�rq�8�}�����=�}7lI��;Y��Z��e���j�E^wvu]m_C�_ϾVU��3�t��c���}.�����0Z���7y�<GH��p�ZFS�̇1�X8��v�����NP��NW/+���w7���Hd��)�P1L��:�O�-[��%}y�٨K�@떋i��ZΘ�2M�z�뽶.%+�}���|Uf���bsE�z|�3��U��X�����)8���z�O�*|6KL�]d���t���ŀY�۹��xL|`0(���/P�@m�������b�#�r ���Dt?{4��sA��8Cף����K� �=���	ѻ��킍���ҧ�is�=���+���m��o@ր���T0��<m�[5�R�cw����t�:��.�ܱ���α�5A<���U�pv�Q5�CL$&7���řJ��H=�#�\x�H��#�Ltt�r��rJ��Sk'TzM��th0L3-T��L�ʖ�$6 ʖ7�t��ɌW��v�r	�w��\�K����]<�ʖ����N�1kɞ����k�'j;�h���a�~�;��N��{�i�J�<NT��>|,������A��u�Uu�G�]L���K U�{�����B|��xF>&vn��<����F�N�qu�kޢ2F��3Ӏ
�
g9�{��]�o��F{ҟ:����h��ԩs|���*� ɽ��VW`װ^֊3�U�$ zだpb�/)�f<�f�&�����֪��)<U"`�n�V���nkfv- ��B��1�� �;�1���.�;����4]ő:tYoc���n�>F���-|0bJ���`G�rmݡ������=�)�,�4H��2_q��p��.EW��*�eJx+s���@�ՒVh����ޔeTr�ޔ��̋9��+�_�Zz+s���1��.�L�ղ�z��9���&�s�e�v�:i��"h�-s����PV]�
�T���VŌ�tR�6犦��9��y�7+.�+M��ZƎ�Re�5[��I��mT��;�:�Y?A87P��>�y�q��T\�E���,��ki�eh�yy�!����HmGS�E7Y���KÒ��Û㚗�஽�<z������ӭ�5�ɖ�@w9�pѽ|7k%�5ҏT��`R].�3m'��i�C��1uĮ��;ɫ��\{�J�k�ֹB���%�K�T��]uv�*�T�3x�j���	}v�ge`�9"[F)��i�7��E���w	��Q�f���e�a�/Xﵶ�sXn�4�r΁�i>��R=Ǔ���LΞ{���A@b��u^����Ι����ҝ��W"N��ӥU��R}�L����f%��ֻ���T5��)��w��Y�a���N����4M�O����(EsY�PƩ�f2u��ǡCX�քK�9,��vt���
w�o/�׆�,�=Sd��S��v�]�M�,�vIڟwk��պ�8x�@�Ꚗ㌃IF*�=^�-&֋������z�;iw��_E�e���1Cm,�b��-�Q�$��r�k�R�M�Gn#���o�Z�s~����Ǫ���e�t�wW@�L�vy��S��{^�>ێ�ᑤT���n��tR3�/Y�p�H󬖩3`^fh<,��;�*��ԍ]s�Δ�l�`U=߆���C��13hÐI���S��!�U�]M@��>R�� �Z�\Ф{�=�{��VG��-��wR�:��vOa6��ˊí���٫Fn���h�qm��z�+��+�D������C��g9J���g_8��r�Af��T�؋�@�Cz�$��>K�"�R��.{�|�0ު=�A�f��%�_Q�3��[�A#�lD�#*3���32�ep����uŭ��w@[�X�ǡ;�+5�W�S�*0�\�_�Պ��H(��d��}7���΄�nnL�צ1@�����P�)ԏmD��S��x��fi��A*g[%�8�L��!Gn�����һ�Fm&ȫ���N�B�R���m�N�8�G�����.Q��X����S.E�tG�g�l���#�����/� ����6j���@R8���YN�Uˣ�lO�J�S;�r�`�s{.���SE7�z�ۅ�|��>o��D�q/
')�B��w��
5F��zU��^Һ{h:#���!�`v�-K�\��&mo ��D��Ӳ���@:�}�3ÂҘ���$��<���@�k���(�^���
3���@�87�g�VMD=.P"�-d>3��7�6�=g\�%9u��3j�u��{���Ka뱅�\���[v"4vj����S+8��V.�V�+ov�=�b�qF�_(�b��ĩ�Mr���3jB�[]tS�ɐ�}�3��yv�����#�Eix�pzoHeII��1`!E�u�� a�UѻrmD{&nҵ�Xx>�Q�)8'��}Ҳt ֢�NWFz��{���#��֤
f��[m�P�4�@~�r���AN��wB���iɱ�L3o�J|��F��ӥ�X��Γ���D���	o:����	��2C����7ATŋ���0-�:72�i
a��[�Wb�}h��:/a=�LYz/i<6�*&�,m�d�Y����^H �y�������lr�U��F3w�s�L���m�Z<�N -�)�:�@E�Fo.�V�<��d�U�����/s����-P|C�\��˯u��)��v����qObxE�ا6�����*�u���@Р�=d������8"PX\�̫��S�C@V�w�2��n�j�GXs�bo��2�D��;�"wA���+��)y���r#|�������U�����ax��B�Z�P�&(Ze�[@=VE7��}��w���2�p���YD��;�l�ئ7�"��J�c�����}��.ppg�|�@�lL[�V�	k�@��f��f�5ݗ.f ���C����F � P�WM���<�X���٘�:�6�+rc\3وO�oi�Xj�;�A��y�N��t�]tB\i�!=� ��+q^p��u�z��R��L���������%N��Q��ҫU���<x``��D�N���0��e>��XnֵXS�O���G��{��_h��Z퀫�z� f�3��S�� ������yo\˽�v��p�o�כ9tS����,dZ>}
=���M��TI�j��3�+{���0�H��)�L{,*����^s~5���p�y'P��P�gi���P"�7�3+�e#Hʝ�Ҽ6��,umv��.A�	�봬e9h7�h .��T6 6�[�ǝv�g�@�0��\GVK*�Zv�h�B����[k@��R��Uh�����e,-�XB�wxY��������ں}��-R�3��1���[�˺�@�A՘Om5bP������vJ�yb�U�����V�	���랆s���4�&��X�p� W#
��3���/<�6,��5vH�n�70�lf�ѩ��Z�	(����q��j�^k�.{�fm�lG�.Oxj�����x�s�-���ȣ(������ǉ�?��B�^�YT�?nn�郝�HƲ^�����V���]#�\~9AҮ�VV�x���q�,��gDL	����0��//��ە�`�2���b+�y��̌�ǣ=u8A�yb^.��N��"�E�y|��:����k5��;��y$��[��vCr�2i�'�E��Q���e�����7yF�:G_f���Y��L�9��̔�¬�K�2�$�×�֣ya��k3�m�C�BInY�Nb7ɇf��{V�u�<��Վ�KVܵ��c�L����P�O=���'D0N��.O&�&�I��*�NQ�j�"h�F�Z���<��Ǵ����{r��hM�"��
�<伣�g2�R.2Z�B%+[���Xud�H��s/���׺��%+��b�*���4y �j�	P� sk@K������"EM�N';.���rWV���	,9+:�g�S�^b�A��6�Ok���������9�٬��VN�2Z��xps34�m
/h�hb�1v�i�.��ϑ(3�B�)�����[1�ח}"ͭ��>5�rI�v��~S��ř��_\��b���	���v�w$2 �ٛ�id��q�Ϸ;! ���,�ppܾU�N��E��a�5�����m��v�{�x��LT��p�sV�v�Eh��m���W-����ye�# ��W�o���wY�9m#�9�zn�SO�w�k"��[�~��t�����A>Q783���0��-7ʍ³��� �_^ܮ���i(�n����s��Fd������.�E��qJ��&���%icu'�`삘�+3������WC����h�
6Rh�M�Jѵ*-�Ƭ\� E�k���{c�o.Vd��,f�ĲIʅM{{�-�U#�
�b��&�8�7F���q*\
�ȍ:յF�����5g^���4++8����ut���+;��$��b{\���:�Q�u��f�t>��e�勏uq��nӓZc�͙�Ӹ=��㾑�4^�#vf;w0$���2�à���*�w;5*D��%E��p�:N�w���<�� ]�dv}�ȋw~]P���ü�-V�����X�/wah³wB2����zwSkt��ۡ2�d8��sZ��j�Aayp���@\�dשQ�����N���hvj1���_�5�{�{u�h�n���p�����]wf�;�Y*e�S��<ް4q8Ps��n�/Yν���8R`�{h���unq�׳���T1�G�ǐ��5w���c�`�F��	�:V>���9��w��$:�HL�Nw���r�P�yc�gW;�����f|�t�d�`�zu��GT鋟��Ey���6Jw{ ��*��X�ӂ����rX���A�e��oc�����@F)�3�/Qw�kX��|q�l�}G^��۾a���nNY\�	v���P���F\���6s)t�d0�ۇr�X���k��Z�[Q 2��LK��v��G�;����'��FK�K����J�˧�o�W\���:$��WK�F]�ݬx3T��.��2�p��#Z���w�m�� �d�����@��Sw��������GRg�{�sL��VDop�%O(�0m)e%�ǡ��u^'��^J�z�"�'�b�H4��qf��8t��(�2��:���#������v>ᐵw�#�v�B1d����XOT�W+:��̲2�wH�&)f�
W b�����:J��7�L�/EU¨�> �(��R�+��m****E\k
�Zж��*�@����L�+HŖ������Z�D-����VUekD�r+�W�,,AVS
(e*���f2�b�-�"-)D�YQD�R+���FV��J�"���*�m���)�VB�"��[i1��ҵ��VT�lF%Q���-*���T���fq�1��G,1��ŋ"��Z�
�e��%IT`�e�X��,DT`�Q��b0D*Ue���eA���Z�l�����%`����VT� �[F�dEb���
"������X�U�
�c�*
�*TDA����F(�V*�F��X�(��*"iDY-)i`���T�+%b�Q
�V
iAX��Ŋ��[e�Ub�"Ȋ�)Z�R�I �}�9k�s�9��gk�'T��^ÄN��+��~	���{��`3+�����)ێ��4��[GAy�e�����r��}��n�.�]1>��F��c4f� U���d�I3=����+��Ip
�_,��Br���\/�˶w�C-h8ʄX�(3�ffEj��z%X#z�F��{5��W]^E�.�t���]f�T4%��m�
z�(aەDB��f�)qƸ;��C_
ܓR��[�F,��\�oz`�=�՜ i�8)�Z�`ۿ���75�U�{���E3Q�!ڇ��(͛�J��w�wܩ\�̎&Wo���i�d�	Y��^��ᎇ������&?	B
���/Я�>��:�y'��,g��ǽ)[W��q^�%�D;�β���t ����1�d8�v��[Mr��q��v���+�۩%�eEt�
ˎSk!�L�`-1�3�L�Z"�V#�Y�R���|�F� ��yin4�x����:�����FF�s+�eCTɌ�C�B�}�|�֦�d1�}]Y��GO��o���^ڔ�а�W���9�2����K�p�и��m��;s�3m���Km}���]�"�-�^f�v��o}���z.�5�ެ�)G�4kۺ�$�U5��m�L�ډp���Z"��Y{x�����#�V��W
�vX[r�$�㩲�y���Ϣ-�-�4�	]|j3�$)%*|�T�8��1aÉ����bo}����.5ʭ�2�"��(u�����1E�Ɇ59C�)�ͮ��K�CUO_��V�^Y�VhUy='��a<F��y$��TG]u�V�E5>	 �ފ٣����4��G�ׄC��ƃ#�����.�X�����	����9�ՙ�a���w���vH�5����>��<o�%�^��av�$O}.�5��JtK��ܘt���x��%��{�<.���q�\�b�&��c;��ǅ\� ,T @E�q�9I��c�sz� �H�.��q��:�(p	��C:K���=�]LZa���L�v�J��n�V{c,K~o0�3�d����
�K���v/w*�0'Qk3��FÕ�%S�r�'ܮ��\�r̜�q��hti�#�Uu�B�¶��R�.��0u�I����ՀV	��/���u��}�a���."��zh����'M�2�~�g�P����.�X�s��=�+e����:�.��U2���!Nz�'˷}}P�#�O.��eq*	
�e�W���JǕj��i@�.a�>���k~��y.�f��	)4W��K8�������t��;s+�tvw�P�{uL.5x*;.��{S���;�
�����޹,"��w�,�D������]�u���]�Ш��L>���i�/o��a�̽���4��ɭ���$[�oJ��[˳�N�t��Y�&�Q�f�K2�!Z[�Yu�8i��mH��������u	�����Hݜ�U���D�aqt���΍�Vw=]F��Vy/EjP��ȫ�v���!�A�L����Z|�/Si�=�,�\��jM8��Z�پ�7�>K�K�	OR��k�\�8���,�M���{���k�\?m"�r>�p�t�~�g�%���KG�b+ǅ8�82�wUX�s�=ẵn�9eA�G��d� j[��#67�j��C
�l�x�(v|���8t>c-QAx��ݓ{�;�Օ��ߟ�'y���C�a�Wj�0��Ӄ�&gE ��ʇ�g?/HI���h�����\X����K��fk1
ý&
h�j��)�3�\Zp�d���u��@a	>� �N}i���^Sn{�dl�c�VM���V�ڜ���Y��ݯ�zo��o熉�'�/�!A�7�$,���7cVzY�������8��F��7R��<�*�}�m���|�QP�G�����
�r��>��y��133��ȃ�O����|:��ǽPt�Y�4
�c���G��t���;+"�6M�g��%N�u�8<g�D�+�^�ڶf��/u7}1�F��S�j+��!ß	�Pؘi�I��#�x��l\�4AՓ��sw���90E��"�э2�Yj��\jup_�!���N�IW�)��)&}���	�<p�G$�����r�uVf��Jچ%S~r�����Ytn�m�O��A���8Et1�,��"�i5�[9��ս�N;V��-�TW�	��h��L�c��y�^Fo��|�:�~����)��X�vY��܂/4�S�n���s�=�ň�#W1~�r�gGB�;Dd�Zmnv^�z�F�&Yd��[�4���ۮ�CMs�؝�Z�����M�n$��[�m}Y-[�j�h�{�+�f}TΥ�C��2��� f�ޞ��Qx��҂�ݰL�=v7�*d��.��l�Ѽ�܀��Y1Xߺm�Y1�T��~�A�7�q�o����x�>ۦc�V'|��z!"�^�u�F|_´R��g�b4|����]2F�-�*���`��sH瘩�K�Xu;�U�����ʇ��� ����{�u���R0�u
��gV�}O&�PN���3���;w�l�����l��Z�杝����;.G+J�/�$$�[���#�V/7�JnXc&��ۋ�)X��!W"�aCW��]iz�
��f��*�����qM۽$a���J"�J�,�L1P���0����{�[}�񝏘y������#�I�/�\�U����/k�
{��{ʬYw�uW=%�_.(mfnf��zC1�`oB���9W�R>�k+�%Ue�N�$n�f�iONO=�WT�5�:���tB�������|�(����k
��{-άV%�>��	���L�L�5�4N�OU?��:��ɷ���!��0-��2�q�	���/ɳ���CA�!d�DFCݮ�Z�\��Ȩ~��F�oN��u/f���A�cl4��,ݬ�F1�����2�oU�ۈ�ܭ� SW�J��V󘥭QL�	t�v��;W���><���!�4ey�duŢ4;�)^*�nݬ�]���@��g9�y��ǮAC5���Ew�m{>0V�p�e�@��͵~�l��a������|^lck��gC뻢 ��[~����YJZT����n�S�V�AŸhՁ��Mbټ�Po����|���<���2e>�]��-gK�x%ݬӾ9��T�CF�Gh���O��zb����ϰU�\��+�m�#L�Ռ��\1�z�%#�Qz_{��<V�^ߏ�|8�\�;�%VY�����{p��"������G6v�֠�ow +4�{8s"�I�"��rdău�t���.�z,�JQG�7ڜ^�ʦr���1�ۅ�׏�����62��s���6���P�q|x\��� _��I�O��-f\�,s��?&�1�g'yk����K��Y)�N4A�"�dV�D,'4_T��ĵ������N�����,�>�B2�ֶ�Sk=�C��f	�F�y�ގ��}�����U�O�����myTmxGB��˜�uH��U��e�tj����q(���lC��=�����޺��.�Ө�Ĉ́b����^�G)ve�bE���y���9��j��t۾'�»[ch�ǉ^r��Qu׾*�ِШ��^~����z�����L����.m��ˇx���w`�c8-��0w_�E%�l��9�	t��gH�w�3���,�A+�M��:�_"l]箢/�+�B���.:�ٙ�]145�{��=n�V�L[��o$D�;{�'-4%��f��K�wc%��X��'��h��@-����ٱ�s�G�)f$��.�e=�'l�:�Ohf���c[R���>�ZLG�|ͼW'�h���tʸ�QǨE��S���߲�gUr��p�w�HJ9�v��y|���A0�o1��_���Дl�mmn������F-z�X�Wb���\���-bhsh�ls�i�r�U�|�W��R-e�nu�s���҅�Z�1:->�����|6��CB��Q�1Ξ��m��}����^xe[|�խB��w^n�U�C]ܖ$����\�_NfE"&�"^Aj�J��n�l�����ߛ��~rﯸ��Yi�d���z4~����w����l�X�b�pp�V����C��8+�k�j�mwB�i���I�^�GӔ���}H^Bo0�㧳r�J�V%�z��P}l:'LG����t٣����y:�ƍb�N�����/�W~���=
�V�s��������2�������	[�\�N�D�{\{�oze��08��,�U����������+lںZgA�����}�iNR5��Y*й[��ç�ٰG�\�n�*T}P���s\s	*K}�>옶�zK�2��a�oUZ|��vw���Q��=�qq��R~ñ�}f�{���x���=W-<�b@���~)�զ��z�ٌ�����r|.�M�����sX��Ǯ]���u�jx�P�&u�ڝ��o��a�;!oO>�U�'����8�!��%�/D�w��3���"Y�z�%���.�A�:�ӫ��l\�$n:���nz�����7ϙ�]�lVz]�^F"}�:ϥk�� 9bv{{��ݢ��a�X��1\�W�)��SH���S��bk�2L+�i�n���n4��g�{{�f�F����¸�s�g��NZ�V��نwx�06��ᖥ��*�7���.�>����\�)z�2�C�I�ǇqoM���������e["ʠ�k=���|��.��V����x2ةˣv1��r���J:W���If�ҭ�'yᒭ�{����#8�c὇�r��u��3<a����m�or�ڶzaO#5���vr����z4{�~R>h�=W/�����9�bf�Ue-��CƠ��MN����T�2^�-#<��>^�m{h3�!��?k[+��v�hJ�y���uaqh�S9ɨV���Vn�YC2)�H���NIѳ�Ua�N9���}����,ֵ8�MK��K�&�mc�
̮�O:�IT�p��#�37����~������J�ϕ>v���}��,�{;ky�Q~��Ⱥ�����;J#VSG�� �c�-�;۞�;��N<s�����Q��-��2�#Z"g��RQ������b"�3���U�wU]3���Y���U@ބ+Ч��:�m�Y[Ka�M����D�Eӷ����������¥P7���Gt�¬y]� F����d =-U[W�% o7{�vΛ�Y�#Tto��x�n;�4S�鐞;�M�OWQ�xgs��W�u������ب7���=��ܫN�E�������p�85�����:�!�1Q�	�y����:SjbI���QЈ����ۦ���ɳ�3FڏL�3�Q�\8�[S8.��]<us�����_Iv���L(��glA9;.���2�&�9Mj!�"T��\F�ٱ�RۣOoN�˂9�/���C���ٶ�>��X��iQO�I��]�k��\;)M�X��m���37�4�P�g0��Y"�0&�wk����9[�Օ�i���t%>UxݻY���#���ː*�r��)m�V��ߩ&������7+����w�KN.�y��m��|�,��j��z�\ƕ�^�x�}S�m|�{O�;�����5=J��p�ӥm!�u�`i�y��൨��g Vi
�sb�Tw�'�7ܥ�v%})�ȯu�>�������^�]G��Q�xި�E=��E7�{s�4jc5���8�Z$plߛ�y�q%V��� rD��,��Ex���9�Vv�>1����-���p��ć��ȇ��p��]k2�m藷ڬ)|�Fi�+�ckѐ��dΩs�!�W����8�Ր��]Kݽ�J���oH����%1����J�K�n�u#/�S�$��M�[8�40d�OJ�{�����}\h�!������fe-d�&JX��׶D�]:��3V�0(X<;jΌ��[�BV�2����
�l� �i`�;����WK&B�]�xB����W��ыJ�[��0&���t���&��}�`���\M�V���><�����>J�gݿF�[�;8���*�OF��.�p��3V��39���}�0=�� ŋm��5b}�ܐ��uҮ�W��*p��~�{Vl�H�es̨��k�eB&@p�胉��Lo���5��sב9��AK]�m�z���3xts���k���qJ��(�x���&�b���n��=���t��<�u��;'�w�]�Y��ý\�p��6c&�TW1�})�I�ϯ'%��݃C�v�����R��6J�R��f�� �R�95�>�л��=���O:�5��`�E5�vz�b>��;	�oΔo �a�1�T~eɛٷl�nDM^�(�Q��*ɵdӓ2�e��=�eZs�w��۝��_B��ޘ�{�پ�ˊ�J��5��Y�|�\�D�G�v�{|)Rf���*&��X6�y�wܯ�iÓǕ�i�Jۛ`�6Jco�>�w�á�-ә�˺�|����sD��J���M�ߣ����2�U���HB�Iv>\O\�_2tY���&��v^�B-�9�-��z����o/�	vDf�"Ls���Ԥ�q����P�۲�V���`�{/��כ���a��=@�Lj�(�,t�M�{�`�}��i�V2��a�="M����=�.��ëE��ڹ��ïC9��Wolt�t����_NΔ��{��.�]�pe�0S�:5���{bU��Uم��#Z�5-��O@�� �ر��4�H��ڌi׸��ֵ�hCNv�(:dsuj�_F�_lT�����7�]�](�li�ˈ�r�3/tU-ҷ��puan�
�4�T'�n�^�n�����h��,p9|��;&B,1}��D�i�Mt!H�7	�0�u�O�6��M[Ć��\y	m�S�[�k�=a�%q��ݣ��n��!B��!��}h�3X$i��o��̱��'.�)��F{Nk.��G%�ޓ����;۷]�~��ћ�6�_���C�h�r��N��	���ipW@�J�`���(unPU���.�U�F��)�7�n9��{������u�}�&v�� Ld[R���v���&命����t����t`7[t��L@��6��rsu3HZ���h���m��\
Y����vp�t���a���M��Fs��4t9���<�����eˏܨI̬K٧�51�G�����EU%����:�h�[�+�o ��,v�}n���̼v'�vG�
��Ī�Υ	�f������{�{]���,,+
�X[b��iQdX�""���,Z«���QUh��EE��*�F �D���(-b�iB���
���
�(���E�,YQ�QT[h��"1QEJ��X��X,PD,TDX�`���DR"�Z�
�(ւ��"�
�Čj,����YQe�EAkYib�[�T�
�QE� �-J�"��d��*TQeeQF�QPE�Yb�(���*V��YZ�"�#�!��j��,J�
(�+m"���D*�eaQ
,QJ����A+�Ym*�@m%�(,V0X�����DE"�ֈ��µ
�AH�X��:��y�ʸRR�����-�jD79P�ǧ.d[��������8���NH�`.�t�.&R���x	8P��-��䊝[�]�7��UX	�г�ڂ�[�YUjxO���<�����Bc��)h�cUt6�"��{Eo]YO���!�:u��x���&�T��lXb2$6zx�,��<��j�����0�mAz�C�޾�CK�-�F_�|d-��QX���z����N����K^�z=��y�m��������U�����V�'ڔ������"��컶��~��o�����X#�lL�a�+Y촵Ѥv��a�r*Ucv�E[�I�V�GS�gLW6�P!0��e#H���ץg��j �Q��ʵ��>��}W�t����9�Z��6�	���3pמ�;{i�E靺4�){E����7���(^�k���A	�ر�7�ڊ�瞿�xl9�D</����G���o	^�,��M��a8Ϲ����@h�V*��aM��s�Q�x��j%�6l���6� ���Ȕ@��P�W�����i��/�g�f�9�x� �+~�;��V-,��&rn+�fe�T�Q[ ��Qv��4Hs���66�ܧ���}�H�uc�`��<��3q�9L��Y���FF��[�Lnv�Qz��i��I��A{w��Y+i��W-�5K$���D�eu���d>`�z�I5[	���&��l٭t>�U�DT�E;��J�퇼�E�1���]���i���XD�u���)�uݾg��5P�f4��a�dvC���Z�������4��ch�mĬ��j�7�{��ә�}J���B�5��A�y��Lۖw�􃰚r޸���8��#[�為��5�+O3X�Y�T��}����i��ԡ�Wܻ��\gL��B��>9W�R=\��t'�)W<%�:8�o��U�/��R���n��0�q����چ5�N���r4-�z��C�gu�.p�\6r�l�l�aR15C�~xr,�cٜ��l��	��}��#9��fo.2�o&%��vXLV���.`��_���������v���{μ'��ᦁ:�/�~����X@�/�N_DZ�4$�	拁���3|�4	���3�.\	*��-�6�'	��2ķ��yd�x���}��&L7P�fL0wWp��ڣ��{�sIKM/�^₵9�9�i�eV.�a��(m����1��ܓaAK�{}/�?T:�F�y����y-h7yk�;��1Ak^��)��l�8}ye����ˮ����뮽ÓF��.�x�;Y�����
�%b�����!�چ_��W��H���ط��%�eP7��|P�����{ud��M\�u�0�7:��CHZ�o;w��E���Q���+u1'�l�1x��f�=���ʮ
O���23��MA��$v�8M��*��bRzJc��y����3�1�g����O��]�������GL:6�˭�<�avwŦ�_���n�,(�\
�8s�g�7,:�05�i�z��Q����M~����S�Q��:VL�4�Q䠌A���2޷4#H�@��ٯ��Mi��gGi���U@FB�"g��:F,OR�1U2�K8�"0�AmX��h�D$���V�"��| V3�B޼��	�D���<���ۨC	�d�R�$*b9\f�ع9wsB�V�(��O�y��\�n�{J�����v��+���F:Y�/�V�B�WnH�gao��T�-�Cˌ��O]O\[U�L����S�N����r�a�u`�v��k�v�u�W�3[�-�ںϦu���:!ois�^�2�{��Ncj�k�Ln9����W�%;���t۶Y0+v�#�K#,�˛��4b���w6)�8챭ǁK���6΋�{7N�ء���{<�J�<$�p.�V)�f���:~�RÙLnX^6���#������d�p?f��u��^x|}��؟2z�u?Xu����7���O8����gY<C���Y&%a���3��2O�x���k<� yG����F�6���{�P�'�Xh�p���O���'hߙ%|d���"��,
�'���݆�8�~5��Rx��9�lQ��ʶ�-�!yz��G�p��8��
���:��1<�:ɴ���8��T<����2~����N�k~d��s[�OY:����>����;�}q�^�%�N�`Txtx{�B���<N��@�4��Ϲ��!�5����4s�:�ĨMw'�6��T<�r��2k�3䓨���>d�y��w�٤9|&�z8l��V��6����z�}S����<C�N!?n���'X�y���d���I�C�Y���=gy�d�T&��u��}I=d���u�)�_�wo�ue�29�o
W����F�X9X�?�C��2捽���,!l���')�.w���W�jGyk�.ԕ(��Oe<�U���VW2]G`QD�t��f���^�;V��.@���V�����r�Lt\�V��:U6�u�M���娕�OY�N/�]}���������h2�|βi52�2OR�Hu'P��x����,�n��d�Vs�`N$���M2OY��p}�H�h)�;����j�w>=�O����:�=tf�Jɦ��M�'�f���?2u52�0�aSHq�y����Ad�t�N$�*l=��{��\�
{ǱD�5j�o�w��Y>��þ�2u���w�8�z�ɚ�m$���+�և���a�4e��?2q4e1�|�SS� ��Mn�:�<K����9����w,�5���z z�x��a�� �|Ý�]��a�fN���M�zwnI=~d��N0�Mf�J���=ed�����d�h�c$� pSy}�����q>]�s��	���{�����%`k��x��N�C��������ߒq��O';�6�'��wnBq�2k��VI�~�?d�'�ųhX�����b�<{ں�}U�nkw���;�|��;0�Oq4�i����7��N>�(i������@�$�k��O?2y�`v�ğ�9�$�i�G|�	�}��>�.�|�[�\~�Bt�ΡY>Aa��=IԝeM��{5a�d�g�~`m��̇����?!�o'Y=a57���O|��]�u��{��º��"7��wb���,�_y@Q�y�$�7�%AB|�%d�VO!���M�XXN2|��î$�gǜ�q�;d�&��Y'�����'�&�푠��+Uڝ��9G٧U�*=��}�	�i��,���C�MN���N!���*V>�VM�d�e':ɿ���	�O��y�C�u��s� �I�<)}���Q���f�����m|2<=Q���i��&�S6����C<Af�d8���;��'RsVJ�$���d�����O�;��?Y!9�>9��**Z��i�G�ܱ��;���D����|�Ư����>��$l�y�|��5|����jl�#�%*�6������e�=�>�΍M�\8\�q��w"Ά9�kһ{qLS!;�p�]]{�u!po^ �Km����R����g�81�(�� �5^�p=q~�d����N��	�7�?$�
C���(q��k}�
OR~9���N#ֲ�������H�G��d -�i�^k{�~�߽��m�w�d�!�5�OY<aԞ�o m�d�O��d����}�PY&;�I����rz���%a��p�����N�s��|�s�מ���5�8s�>�~��+�$����:�2Ì����ya�N2�y���Oq���2��'���O��sxu�by�u�iYv��m�Ԭ8l��6�E�+i)�M��� ���������|7̒�$����XORi��C�'��jya�a?kx|�d�N��}�I�4��>��OP�o�u4�>Aߝߙ��y�d�_]�6oRg����c�0&=�y dxs'��;;́�&�4oϿBz���'�d����XO���+8�=J��Xu�O�ِ���(7�I�d�u�6�󁙧4������� mH���d�\ì���y=�d�&ߒ~��	��|�+'�$�Y1��,������Y�I�T�� ��s�����}O9����}לu'k��DP<��ϫ� {�M�f���N��~ì�	�o0�&�XOw:��;d�哌����+'X��|���N3Yd=g�N'<޻��~W��V��N����G��{��L?w8�ĬO7�Xu��Y�)�}���쓬<�a�N>������'��4sY'N3Y������1���{�k7�o��7淾�Ҳ|�L��C�?2u52��m�_�q?2M�3y2q+�R,:���6{ܐY:��w'~���_�� �Q�d{�E{��:��\F�%���\�^����VI����IXz�)�
��,<���m���)�&�q5����$۬�C����yy��':�����	��g�̛d��.��=�榮�;{�n� �!��&�{�7����<��[u�}��:��\�^�k.n�ht�0(=��m^��y�j����8G�E�у{��lֻ��(��j�\ݛ)��9D�Ae?�<��5o�Yw��QvK�Z JőTN�Xg8fg��� ���e���� 66=��5W���[&��B�O��?d�	�Y�*N �Y6���OL,�i8��P�?0�f��:��yC�0���77�}��������wx�b��P=�m(q�d{��k�'S��$���!6�2k�dY'��%ABj}fЬ�J�P6Ì�J#�� @W��}�8�O]L3F�?�����������&�Rx�s�d��C��d���d����w$�i��|��i�]�I8�?Y*T�G׉+"�1�R Q��{�v|�����r*�7���ٿ:I�'���܇2�q����̚CG�ɶIרy��I:�9�{��M�����p�z��s��|ɠ��}���zc�8�X��6��{��w�}�=IY5�R|��&�����m������'Y:������a�����c*�a�Iô�M��99܂��z���Rz�Ϸ��o߷��ֺ�^�����7�gY'�;��J��ovE���*N |�O���C��d?���O8��o m:��'�Τ�ʇ�ϲu�$��o�u��)�_x�O?f��;s�����w5u��2z���H,=d��c	���ud���$Y=|I���2OSS�d�!�^a�:��$�V�c��<5����& �-��ёtr��]���RLOڦ�>J��y�Ĝd�+�,>d�{���u�[�$�XN3F�OY4��&����I��k����<r�_]Ɠ�_Qf�Z�����~a�M �~��!������3S�d�N2�v�m��l���&�4o���u�G�����N��P�}d�.��=�lz`}y����}�u�����o�m?2|�����!ĝA|��8��4s�M2OY����8��h�u���?$�k��0��䕓��=�1���1������&is�+��&L�����m\�ͩ������*ژ-�A�j�Y��;/�V!�]�ύ�Q)���AS��+���c�3lZC;m��ў�V������$	��I�2��c:e�rd����YM �ԗѻ|��>�E��}��}�Bϒ|�{�����B������C�'S��6Œg�2u���>C��J����a���:�a:�vβo�	�w�u�G@�����{�ؼ��V:�x��ػu���~�����P��!����M�A�q��?jè)'�d�T�����d�T��2�:�G?a�l��<fd��k�Nӗ�=���弓�Jek����}����{�Qb���	�C���+'h�l?$�4q�|�SA�è,&��[�q'X��'Y;�	�rAd���}��w�5szp����ST��߅Fǽ��� q��w�'_�5;��d�3�?d����l=J���!�I�hˌ&�q1�S&�w�!Ĝe`k���汞�sl���ϒ����(��=뎏|�{�@�����'?2x��Ox�V��&��%I>g2�X����B�q��H|�:���6Ì�﵍��^j��-�8�`dx{��V׃�yl�K�:ɷ�=��u�l&��x��O̟�I�q�L?&þd&�L�9���C��쒠�3�m
�Ԭ�a����3����f_ؾF�Y� 2�=���O���\�ی����rd��C��8�<v��9��<a5���Ԟ$�Ӿd�M2|�I��!�I�PY'���ڇ��$�J'37���[oޘ dlJOYRTm������3Ϩu�I����~d�>�N$�x����d��{��&�z����M2|���P��!��]���7V�|� ��vP�I�7���I>v���+'���d����_�'>O�ϲx���N0���'�9=�&�LN�����N��_q���D��x��XOg�s:�1�\z x}�PP�'�,�{�:�̝�1�u���d�+	�l�&�`xe'>d����q����x���N0�t��M!���~���z��7����v����Ⱦ�<�Y�*�g�J<*ujxŽe��^��	�����_}�/e9������n��zh>	���t�]������uAZ�^� �Ɏ���\*�}�tG��_r��iS)h�`M�+B�h�jFP��1N��-�#΃��}�}���9��>}���&%a����u���7�4���w ��OR�Ѿ�'���k̓�57�I_'5>�N�`~
�{޸�����q��B_�g�-]���q���=I�����8��o:�m�CG7�PY&'��Y6������'|ʇ�}�
O�?{�I:ɭ��W�O;U�썏{�'2>��B]�i��1|R�߽�=I6�ϐ�������i��:�߼�&�8���0��:��o���!��a�N%By�<I�����;�=g�=�쮁�} 	[�j�շ[�U�UY˾����߾v�'��J�i���t������u	���4��({���:���ԓ�:��gS�$����d�L��� G��#�g/����O���K���}���̛d����Ld����OZ��'Yd>g4��:�=J�!ԝB{���N �h�y'�q��Y����I�5��:�d����r���㷾�����r��~�Ϻc'�l'g�a�N2o�Ouܓ�����VO�}I�����є'�������&�T�Ad�~���'PY5���N$�*~�?u�_u����7�������П�~a����I�Nfd��	���q�������&�N:�d��̂����a�=�d=O̜Me1�|�S_�q��a��]y��wW����y�o~�1�iX9�I�M����H,�a�}î�N�峬6��NwnI=~d��d�a6�����!�hz���D3�: �=��n��S�__=����I�~N���~d�:3�d�V�y��Y;�O��'X~�p��N2~I��x�L�;�!8ϙ;�²O�C5�Lt�ϟi�~�S��e�VV�[���+'�,;l!�'SS$�N'�VO̓m��q�yCL�d�;�r�'�s>v��'�O!�`v��0���8=��̔��f0MP���b�a!���G��0�����9G����W���y�D��{f�h��"��#��5z������`нO�4ۻ6��>�Ω=�ÛJ/yj���bұ�V���{OXx���i����	�.�g:]/�^�\hIl^�)+�  
����eK?xLx{�������0��P��A`�m'm��I6���V�I�~���N�2^`z�x�����d�����x���z\?�dJk�}��bχ�=��lx�ݔ$�i�G|�Y'��a*
�VN�d�IěeN2z�k�\I8�ẏc�N��i�I��<����߿�F	������/�+��yǇ�d���@���:�2|Ş��2jw��q��IR��}N0��J���N u���'>OO>�|�N�q]=�w��v��5<R����<7$(��G�xvs�xì��i��I���AC�'�,���P��]�̓�9�%J�x}x²m�Yd�'̝�G}�{�5wn��Qw��J����� {���{#�p��z�L=���bV�:Ì'��s�4��)s�2z����Rx��k'䓉7�%Ւq��~�c�;ۅ�~����k�u��"��̲m�����:�}�2x���$����L�CϷ�d������u�c��ru'R�$�'�X|�R|��|���Ǻ7p��m�m*�wx��(���e{��qaL�Y8���OS^Xi�������M$��y�>f�8���a'�u���è,��y�:ɴ��0�����{�\���%�Yu[{� �����r��2h�ϿI8��O�:����O��2�O���ya�a?��ɦN��OO��6��:����I�a�n��m����t�_
����>��{�@��5�p=a�O��zw��M�joϿBz���'�d��Ĭ'�R~g�g'�P����Ǉ��^� �����8��ߗ��7�x����V|=�8���Y���<�0�'>��O{�Y:ɷ䞚�@�����2J����&����іC�~d�h�8�=J�'��~����{�˥/;/+���V-ur�p��Ap-0g8m�Ħ���ߦ1:uL��YֆlxɄB���d޾����4	�&��|h-c=�>�wZ�	]4�&������+hmtJ����]W|\^�jg/'%[��ܧD�U�p�1m"������j����J&K��f��-M�=Ww��GRt։s��3)�����M�Ev���H�����$��m�/�w���C�{5C���dBC�@6�g��{�6h./b�l��MpN�t^�:zN�Bo�e1��uO�^�ܴ��hK��Ͷ���Ľ��ɯ��:����m
�\�#s�֍c)�]��.���=�I�m���oC�����}��-FT��+��S�`�8��&��&����z�K;��7��[�dS� 0��]s����0f�m�;bB�������+-�����jTDӹՓ\y�&f�c��F��2��1��H޻������F_:&:��A�đ����\���0C�e]�5�䄳yGn�G��B�����2�E�z��$��Lr�K�t#�J*�"�]�٠\p,�p�+9�c{]��Vyo2���jR�n�`���Bp�eԞ���d�Zq��G˽��V�T<z>�f�o����|�\�+�ͳ&�N':�ݗ�E<oY�]�� ^��<x��}�,IͬS_9ӝ3L�m���L+��-�:��YY��WP�v�u��9ƓT���zZ;�y"s�n,�n��k���a��}��s�V�1�a�u�Q��]�Asa����<���J���w{���XKmzzu�g������r!uM�%�p�J��/NXj�1(��YPV�}7��`�[s�u����.���F]�N�%lK��1ŧy�N�!��[\��f�h�]Fb:*�0 >�'9x*Ry���Q(��Lw��R��L���k�&�7�J��}s��zx��M*q�˴���xP��zj���8�Y�U٢ܷ:�L�9�IӚÁ�wt�5�N�0��T��X��qħs�' ,�IG�L�[�o��'���o��y�q���B�����t$�;��Cu���h�Z�~��G{���^`vJo�g��;r�]��|F�'f��Mr���؄��wy�e8���N��J1mo.t��h�1�a����%ӕ�<1F{����:�V������*��Z*憳&���ݖ�%�����X�Vb�T � �u�z�����ݷrP@�@ƺ���!Z�Vv�#�'m���j��MtQ+�bŧ]|y\���ʄ�ϲђox��S �݁�e�Z��V�ņK{p�oq�KT�&莘�]�z�YVJ{ʕ��.�,�cjdɚ	ܨ�9��_M�wk���%�:�[���ͣ�Κ�G�7˸.��(Ƀ�*}3h�����,�W�9��
���k���v�eL-���+Uo���[�ջ�|������[�}��Z��QVʋTDUEB��PPU"*�dTD�Ŋ-J��X��T�J�*V+l��Z��������
��dX���X�TU1�QBҢ�(�[H,��,X"(*֤k��A�D��T�ҡR,+
 ��ADdU(��)RԕP-�PUX��QQ,X�֤QE�QY,U �[i���c؈�����j�-`��UPD+ږ%d�UFF2(�2,���[QQAQR���2
�b��E���mTU��-�E+b�UVV

*���@EU��(�U+hV1�VJ�Kj�b��*҈�V,@FV�@��
��*"
�YX�J�Q��DUeB��PPX�0U�T���@��][Y�G:�����;3h�˝{s���]\���*6�ʺ��(�!�;��M�t�!>k�,����{���{��T�Ԗ>ˤ��$�UCi=A@�|�AI�N�f���N�����4�u���:ɷ���@�_�9�rN2O]k$��`~�@���8��(�9Cf�5|��os���2~N��I�f!�����P�'R�<�"Ì�J�r�P:�ܳ�Y'w��Y8���Ogv����N>q륗��Dÿ��ؒ�m��Lx\{�KCIY<I�k)����єē�8�~����6���8�Ĭ{�"ì�}C�{�'P�����5��;}�y�'����岪������{ӏy���O��d��̂�aRq���!�N����m'�1$��o!�N{d<��񓌝}C߻�
��>F�[�"�;��1�d{�=�O*��̟�5L�ܾ��J���3p@�ؘ�]���:^Z����a>WW��ʗ��>��0�|C���0��:^cO���s3����v���\�|�M����#:��p�/��{���'{5,�Kr�����h��$grw,����7���Ԇ�m�;˛Nr܈̌.Sti�:q��0��s�]���f�׋�Y=�Ƀ[y�9Ct�Gim�:Խ��M8V��wcy�R�F���/�D�5b�ˍ�l6�zձnd�|д:a��>E=��tA�t�.�`R�Yw[G��Pz���4g)��V�%��/��mK�t��M�mY-�����G�J��pi��J��N�m+<x��()-N��m�e�եer�x{����v� ��m�������=qh�nQ�ʣx�g���\��"l����OC�Bh_>����f��G\Z㕒��$�t%Y�1��xޥ�Rʮ�*�?i�y��-j����=�/i6��u�Uq�����I��݇�ݠV�.�[I�T�_�5�{�
)uT6Tw�{�X�ש���rb�.˃�Ĭ�<&�4/�8CJeS/���M���nf�R���~�=�5�ys��=�e#/��+Bpo�Pm&U>y����*�����Ӛ��5����sF��7��3:�1�%�v�+�l�9���	{��[ہ�K:���(���b��+Aw�t������D^;k�>��U��X.of8^ܳ���b��4A�b,���\0���jg�ô<�\+]��O���ں��0��C�סo���tk��d[�ՙ˔��F��.�e���ptz&�=/��
{�����[��q4j!n��#�.h<q�002�u���shU�9ջ�9q6��pj�J�\oh\�vN�ǷKc�'���#�Y���FSV���پ��0�M�kR�[�磌着V�ήب���!�zYX���t�do7{���n����Muf,c��xld/C�U��؞��v7;���Uv1�l�F�vv��՗Y�غ���Wl̕�g.O���P����K�Og:����)��ޗtʸ�Ì-��IUϗL���r�k_$S�9�8��QI��֨��&A�1��_�����u+{�1{j�XG����i�y��|ξ/y�-bZ��;Y�ma�z��n��P�dN��b_>��9d�t��;h�*��-fޔ/V���+Z�-�lZy�Xhl�"�\2;/�j��{�����Xxa��YTRYƅ��G&ukQ�M�P��qK^K[�ޞ��
9�������&��H��^-��!}��қ�q��w��wmr[v�N�g,c}�[�$��oE;��﭅Z$�5x����X9�N��>�Hh;eXvo�6�LV��=l�t^�ʗ�v�;32��w��1#T�u%��:n��;��䏬��Ӿ�4��@c�������X�y��/_ػ)���D�K3��JT/�Q�������&uw(�3�~ x�՚���]�*>�O��k/�Vm���Tm�CGӔ��׼2�����n$�3/����q�����j-O�4��ɍ+�B�j�F)�4�=8��m9�DR�g���V����T��a�-,���J��l��<m&�kw�ſC������������<W����v�>���B�^,�ұ,�]�a5P$j�(G. H�zx:�F�Zi�c��ɝ���ݽXj���a�B�`H�*yt�u�6��`�nFL՚�&)7��yfwY��᾿l�΋�>vx##TtT��E�0�;��Ξ�$�p ����K�x���p�e�+M�2�\Dꎾ�N���|R)E-��bZ��?G~Ҽ/y�D&P!0��ei)����
��ai�[�Z��R�������]��=�W�#瞓B�"`�����:�p�r�:�M���w$2 Rv���� ψf��ج�\[#��*ʛ�b
I�sKuoL��#N\�"�o_$1k�lʱ�v��aZ��Cn�Ea7:�f�c��e��;$�(QS��5��T�+o��/{'LN����.��.p�v��5�mŽ�U�U o��҅��B�%fQY�R�%��nݽ<4�^�M���w�XL�g�U�[;,R9N��/9R�ì��c���A��w�㷙�H��L���q;�����c��|�,���SR��[c}�����о�DNS};��6��P�f��4W�&p�c� _�|2��/��m�U��I�1y��	�c2g��^矛�T��(0V�����A���ږ�_E�����4�'���Zd���g>�~�A�7�u���A���x�}���F���{,����J���u^.��Z��;�O	�k����Yb��jLP�91ľ�VFx[l���sy�G�NuI�i�Ō �;��>϶b�x�'����v�`���-�O���ŵt�V�a*��7㽵ԩ�cvcC�3�.�!y:gS���.Q�p����ς�w�]N��|�u��e̮I�Zh�؂U*�ԝy���<Ur��:��Ա��\�����ݭ/���,��ɖ��.oT�6ʸ�Pr�QAuu���_܋�)F��<HT��}�}_W�]kM:�Տ��gӯg�[�`K7�	����a�'� �@�pgC4��V*��V��rl�]���﫝����o���C��-ɳ;�݇��*����V1ሜp��k�)H:q��'5�W�$xe1�WYc��ǃ��}���b�@�y�(3L��*����MQ��X�L�范�%ي�.�kcZ�AOcb0�4sH�=qh�F[�s�oC�x�}ћՃW����Z������MZ};[�hÌ�Ţ:�*�tծ�[�]׹j���Y�ŋq�scJ֠�-#S��ϗ����=��p{�5�L��N�I,J�ʏib�f�/JeS9ɨB�{�Y����E�S������[�"��q�%d/ա�}��W>�I���F=}p����\ў�����ǆLuwE#9L�_ABt'|�I���f�.��PP6��o����;�ki!�u
��b� �.�,��c�3�qY�C>G�w�.�4�1�z��GT�t�[�wmǈWX�B�h�ߚrE���Y�W�m[{ݽ��J��o,m�T���[�n��MtI��(͌�j5��Xz�!�A�MS�_}��^�.w��]�.�?�yob�ȉ1������%��A�/�+���q舘�{��b�����[�`)��a��P�B�R�d�jE�%e�9����Dg���{�à�U`������Ҩ�ZJ��VvE�a���|�
��i�E���<�\+]����F����;�B�z�<7���q��n��'��AzKs�w��=�j��n���D\�*7|@��|�%�q�R�z�W��ЪN��~y�W/�/��dy���Ӟ]Ǧz���^m�<�x�^�a�F#Q�'����nlo���xq��o��J��٦7-uä
c���e⸇\:�V�j�������5�i��]��X]��y�-j�&P!0�1��iuŢ4;�B�t�#�wc��.��8�7}o{i/o>��J��'�b��nV;��mot�����g�M�}�+n�&�>��x�H^�T��5������k8~��M�F�q��\+^5|�bc����Զ�y��E�L�ץ�����(a��p�]g���m��Zg؄�/��{�D����._[ѓ�J*3,q�fw�ﾯ��+z'�Ylį�m�>�xE�@���!ڵ�c5kPm�l)�m��ټ�՛��]gu���Pr�[�*��(ekai�G6u1�Os}N��<�$���^�d�a[S�;D�K^˝j���u�����3(�i����S���ɭ����-�`��H��e>4-��5�Ք��D�::�zޅðgCeS�jZǪ��EF،����Kw�q���D��ߊ~���(綠��l>o�/�`}���Lj�8IG�u+3T^������g��3�qA����: ��V�v����������ɻ}{�ds��eFC#y�凫����<�{@�뭘<�xZ��'���(e��f����z��������u���k5�U��{
��A1�9^�-��z�XT�	��<��[G\�4L����!j�E�C{r�$�M���J��ʧ��aQ���3��c�������vP�M|�vB��u�yu�����w�jq.8뾼�{;�@���(�M|��H2b���(�n����h�;�[��j��]ٿ�x��&�ҵ�����bY��	���:-�������|{ڵ��-ۙ5Xx��������]qK��X6��SNڱ�_����tϕ�XQwQNd=~�+����ݐm�{�r�������+�t|�@���y�v4S5��%�����=GԺ���h#g��������y�-by��bC��}���vה-���c�~��g�rm>�GE�"U���x�`�҅�V�6"��z7���9X�q�JD�]�Zر�4�m�>ˋ�+=+YQ���o+�p�Y�ƃ�Ķ���8��;~Z�z�-�n��n�.uG<�����q��ϩ`3��'�|T�`����)�L�Mn6�y��]_E.���L^h��g:�kZs��2����EhL|�I�]���,��Ë1�8�p�*��y�!���4ϗx%��Z7�pl��į�I��q�^<𬅥O.7Bϵ1C$_���ixyx���c-�x�L�{�fK��f��T%�()���	�yN�Ω����X^�����cy�@�}�U�J&���'\y��U}R� k)̻�+9��L/n:�Vc�fV�@ڸ����d�ռ��=��xM�Ěq<�)n~��^Z�7=�MA��r^�^��a�u����u��˶�Z+�v�K��>�fܳ�Ϗ(��~���:�����
�PC���9�ǻ�{�'�=�T�]p;�0�:!}�X��XC��So�&l�﻾z�񸽹����)��O�Հ[WV�>V �	��˨pNWoe�֍�Y���	�-K+k��!,�_�3�gK.�;
1�����A��=BrQu�7�d�ȳ�^y�����-_��e�+im�Rb��=��Y�۽���T���u�Z�J@:q��9�c�j�W5D�u6U�}�g]�x��4�\B��i��5F�-f�;4�(�� I��9�v���^��a\o1��3���і��eAW5����2{���v�ڮ��zz������i�����6��=qh���n����_{#Y�Ct�|���6���%v�ό7�v�E,ǀp��[a�Gu��.�����âA�y�M����p@���OR�,�w=�����x�WL��.�	�9�����,�w"g��z{��*����ݩiqo0h�&�=\ts�k�Ɯ��'V��h��]fyD<A��mI/�y��	Z� .Uځf��]m_�O�ݲ�w�3�&�ᙖ����ʃWC���K�>�6tkc�ZB0�
�:�sns���:h:�\e�
�>}��@����I-+ՙ���r�@�*1z_6�r��9���}�� $#&���:F
�J�w+`iz�zw�NvߜO��8 ;�	����)�x�{~�5:��	�� �$�J��&�6h��h��#,�\"�v�ze>8.:���'�����j�I�h��|q�ӟL���X�e,�H8�j�M�`���um�}:=t�V/�<�ԓΔ�#�V4��N������B�ZD���:勁��xsqR�'��|G��c,O������-^�p���vOK��Z1.'�_�ބ\�5�u.��R���U���6�V�W��e(�w��'PGp���üo�W�E��n|��T�iW��/�yB{r���?F5`�Li���2�#r��+��S��+>�m{�N��Ye9��/�V�T�JU��oz?:`��,��NVo�z넂�kiR������9s��4���a��?=ᎀ���$�a��irr���Z��ʽm�*	vˬ����^bwn܀��q�z-Lsw�c5/qkY��J^�}�͞"=��ܸ�ⳢV^�r���ެ|Z�MYP(��P)�(+�}3��I�փ��}ۍ�ٻ��t���c�~7H�j�+&oD�uYW���p:��^�u��v
�ۏZW��2��TJrA 3���U�\u�0�Ab\ܕ-	�A���]�&��նx��9yR�,ʹP�	С1CAg���|-JYF�&tT�U��zӹ�	$嘨���K�B�gg�.9-��o,V&��ζ�ν%<��t�K��p�&���_ k�t�q�k"�r�_iT��i'��ƣKiۆ�j-�@�FM4S8;K���u��k���J�f��.�k�m^NV�b�p�9���۬��*N�Ȧ���}c�����F�0�2u�Q�=t6�[R�ޠ�e���%Vy1�M���BZY�,�6���be���
�n�2��qb@+W�����(�ӻ�Kg4���K7
�H�
a�ޙ�9l��ʔqv�=%�(�F�s�ƃAoP���p.���ܝ��30P�Ո<t���K�w�P&��-Ǫ� ��׬v��ژrf�&����;��9(���&J��Ge�>e=/w�y/?5%�����^u�6�����`�z���r$�[��w���5`#��
�E���Y��Q�,F,QEQV1DQ��������*1cE�,���(�
�`(�lJ�,+(�֬"�ڢ�Dj*��D�aZ��PF1�PUT`�"�,eJ1�
���%J�H��IZ��QX��
�T�(QP�j")PTE�b%�c��X[b�"D`�Rґ��B��dD1m�����V�UT
��"�QU��m"� ���+
$��B�cj��(*��TPX�(V�(��T+U+X��Q�EAb������*��
��
�
�im*V���Q�"%�U�����H(��JʌDciQED#RQ�����,R(�E�X��")l,Aőb�`��U`����@$��
Zʅde���Kl�1F����QE�U��
��FڃhT�,QgpV��.�æB�:���g����&1�ۉ;�B{�c5}�'n`9i�G<�/{:����Y�p�SD�WD������r�\�j�s�k?x��o�V�����y۸��/��r\�G�T��Ds�L��)��(eka)�L�mA���Q�@�BWؑI'�bjc�g(��e��y��W�jz�iL�L��S��˝#A%���6ۜ{ٝ5���v�/^ߦ��)')�}
�М|���QwѴi>���R	�f�=�ԡ���/
<����d4}=H�3�X���f5�y�M�c�5����[�\cѽ�A*O8����6坧Gh��Q��r�fTΥ��뵽zg�_�7ر=��2��S�('K1��q�B�<�A3�ڜ�v���9P=H�5����o�Ֆ�ջ�y��Ry[�{�<�5�mx�Тoן�~��U1=�(����,Ax;��G�Xb�Kj����v�j���}F�нr����Үl�Pz��R�ᷛ�%�ǆ�a��6�Ta��Q���q2T�\x�Ʒ�ީ�������f*�93�{n��>עs�f��B��/����}�H�eƨ'b�ҹ�R��s�ھ��U���ڬ����u�������y�vZ,na�!��ۊc�s��{�xt�{��k��;�O-�t\��0JvJ�Y�@'���f��,{,�x�ֵ��%k�u>�)2�C�
c�&�Dʖ�ï{�쳷2'd���w:��{X�/�k�V��E2�L,��c(iuť�o5�t�.N����s�m:%���]�>������OŎcQz�N{e�a=�
���3�e��y�K�"ʣxZӔ�j�W1�-j;������7�o	���3I�Rej����q$J�l�����������{[�h�$���N-�����vo3"���Y��k���R���Q	+���^uq,&�T�X���oq�$�����)�%t!���kN_���YJah>��I��Ե��6���d�ף!��9#l�u��mY���5y���8ty����:cS�N9�����T�`bH
�����Y�ĩ}����N�~�O�������4nI�8I�x�qSވŷ�z�n���6[.����P[��6(�mhw�+���V�\���D�"Q�+QzndF7�oSY�j�:����3m�v>z^/��p������>�~���]��>�bFgQ�\|'������ _jΩ�;W-��|k�w��C'7-���/t!Q����q�k/Э<�5�Θ���	�N"�gw�[e^omU�9]_�ws�D!�����@_���ۚ%n`��N�V�>�&2���Gg�;p��g�|�%P�qC�ˌ���䩐p�M�כ��Ip ��?x�=��L���`2���T�D�Ttk�DeBG����b�V�a�I��k��:�����_���ޗtܜ=�2�=7�5*w��%k�{زjò;�O���9�D&PL+��J/N�Wqкh�[�mb���"6���g��n��oq}I�^T^�Ԇz&�|�mߎ�\2�]��,y��0�#�-�ʼ>���+����]:9��);�	��Lv!7ϡ=f��[�����u;�"�dQud,(��֧f�EgA��S:�i�M���[��#��~�40%y����e`=�=vZb�s}F�ཐ������csG+~�̢��Hk�ht�z�P�<@q�C����G�wC��52�U��0Ų�q0h3B9q���{��v�kibYU��V��8χ6v���"�-ֳxu����g#:��qM�œ7���>։��b�(R�[4�U3���in0^a�2�z�z�U�qcU�����#+"�xMhh_㽉2��}/���{��q�Ȓ�����'u��'�nex��@,��U�+�Gt|r��OD�e�t�1�R<Ƶ�N��H��Ϭ߽���M�c�l�a�	;{�:��nY�슛�
nv�7���,�:;G��d'�ծ�ɽ�L�fy94�2��O��q���w���\�,��Uw�{�T�	�qX��W���V�K�Sl:k�}	�O�Ղں�;�J�A�3���U�b�yn��Uj튈V�g?�D,]�%�V�}p��	���G��1��3�3z���Xݏ@�=5�Nu]=���;Y���K��޻��Bw���E5���o�,s��M�li���VwL������8�ִ'oW���5k4OA@kQ�!�hF�X2n3��1�r�#��[�J�hR�ѱ(t��,�"�^�u5þ�>��e�o�ɫ>�-�\b$�rQy� �.Y3Imr���=��Z��i��o����H�N��2�ԫ:q�t��O'k{G=u�*F�W>]�r�>lv���4��Z�[yt�x��Hw�۫is��d��8��/�E���)��@�2�4�\Z>іϩ^C�p�<8����]�/q�Y��ާ�|���i���`s��=��u]F�U;��ms��r���'me�k�N29��Z������l[���9����gy�9��x�OC;p٭�ֲR�:ذ4�B�r����E�]��YMsFv�r��sv���̊fq�+"���{��)�G\͹��b�۵jt��ym�ۅ�ۛ���g)�}�h^���i��h���QE~n5]��G�jc桫���[�1�#!�=H��w�h��x���<˾���������k{^���Y�tv��a��������C�r�Q���h���\[[dQ�s�3�$��ip½�Y�	^c�Ζ��J��9����wg\�.��j��q�����<F���:"���[;�J_@��)͵˝����}��K�U�Co%d�0Ceu����psN�鉣�yi?�V�|��Ž�k�G��Ϻ��V�w��E�*���Ӆ��x��3Kll�"96�ϵ��u��=�;!�u�ԏ��˅k���[�u~-����Z����X='�6؅��oǯ�O.��4�ևJ���~s�c�������v�[��m�˫׷�M�d�
�05GE��I�bw�"@̈́N_�@�������J��bn�pe�����+][��ۊ��9D>��5��|�Wk�$f���!U�b�hrf��0����_�F\#��Ƚ����o����-�>7��o���{�s�))ɑZ�`��^\��]T8��z��^��&�s�e��ڀ�G��?�ߥ��U��Jޗ�7
�����y�J�{|�wL�/��5���e�C��t�(V�eq�G���6��#MX��o��=.��OG+��2tW"SWf]�{�ج����o]z}���"ay��ō�P�z\1qveI��j�r�w��)�+x��q$�H��f�E��C�Qz^����+��I�5���R���q������{V�`�p�]�r8�-D��,)y݈a6��攁�k�k^�.ݝGrTK����E��D�s�{q���B�.����� &�o��0�wk��:�ص�\Ōl���Udm��C�����[��a���Oh�-��+����-`�|g&����C��O�a��?
����X�(��	��c>��h1t��K+�-N����҂K4!.
:�Me2N�\-J~B�Դ�o���x�ߥ��L=q򷯯no��ZZi�*���\�]�w	>h�
ȌP'P���8�j���kvǯ�sͿbP>D�P�m3\]J�اr$ve	��l�e������^a��K��1=,���
�T]�c��V���Q:OPtNq��R��.g��s/g%�p3M��I�B��!�:�t��~��LѸ(:�30�L�#�@k乮�:erL���J�����)Ӳ6��-�~�7Nzw}�o1����I�`x?@�[�@
�h��0��t����s�E`�fs�����t�9�)y��V-�9S�u���4���YM�wzS��{���KH�P�;Y����Z�A��,1*���!��vPוb�@SB�'�B��!��^^�5槚KH���͊ԗ(���|�J��-t�M4���ʊ终>|�EI����5
[F��Dt,�2�������s1�X��vwYe^Ҹ1�W,�2�aޕ{Ţ��p�;�ufz2*7roR�o%x{�<��ǩ�J��_����=��6�%��m{}J+>�T�ji˶^�<o�]Z���~�������mFIY!����1h�C=�؆�_���{�ś�����f�#�9/dzq���2�4Sb�+���9�F��!��3���.鑚s|)q[]���:ڼ����$���������h��h񘞥ҼG��!�l�s
�Vd��|�[���$�s~^O��D�ڮ3�X^�#\؆�l_�y�2���w)p��F.��g�Z�ˡ�x�33�����S<�rfتb[]��Br��3})�ٱ���}�[K{�&x�x]�ln��,�WY~�WQ/��W(�|*Ds�;&ly�3�x#2����4�$��7:R�o�J�ꗮ�|�<X��Z6�p{>k���N$py��,���j��^��l�ݍ��5WM�:#5��L�f
�\���U��j<�U��:"<8��4��nN��`뵺:���!l����{}����̤zU#�ɚ��K��#�ᣤ���х᪽Z'D#.��3l��fW#���g��rd�wF�4�]lͥ��jT�LYZ:��[�Z����ׇ� �J2�#��r�Ιv�;S��o2�A�6��Ғ b�[�~�t���]�k �����d�@��(���W�&0�-�J�����|�Yg;D��o�p�M�����H.>؞�l�OZ<eNs�X3�p���6t��ކ����B�ޅ�����@�����xg�p.�ݎ��,��&9`^g�G��C�8�x�W07��r,��{����>ڞ�p�^������/���+o�� 2�'�.7
S�^���夹�Z^�uP��Τv֞��Ϫe����m+l��Oe<�~|��Ug�I��lIP��`�,<��/���2�-s�o�MSx^����H'���Q�v��*���2��s�=G��4�g����因��bW"Hʮ��|�SX�Ÿ�_j��鑛��'���=KK'mY��Gz���C�n�=$Xn�ޏ$<��o���K���g
�S�L�c�cJ,�h0�;{P���4�=Vz�8}ݯt�.��p�8�Zqכv���*��u��#�m�k�3~��k�l��S5;}7��gv�<`ν��5�����o�|C�����#�e�0K�#�+�j.�V�/���dH#��E��qW�L�x�)�E��їw�T<t�u\�	��9}����в{�K�ޭ���Df�[x`3Ot�K�3{R9��:���9�o�����A,Xp��=�ڻU�yX좌�[�]<�jY���Uھ����u�<�O�y�+�z�����>ZV���X�������X9���Y�+�ȹ������
A�7��e���9.wV�|\vV��QE���e��4���=���s�GW/��M�'
�Xf?��i�^ub{��G������R\Ϸ��(�C��-�����b�(�!�F�V>�ݖL,b��ϝV�ؠ�û��!����
i-tw[U�;v-F��$��TG_]�V|���6Q����%�b�08l23��F�E�~jtk���?-�W�`�VՇsýBT3�DñH��,	VWml'=|��*�W�����+޽^�y�Ì�A-X���ݠk�\�J멗�)�`g[�0M�F�Q�K6-����l���^yg��g�OL�9�=s��� �XZI�)��_���8�RZ��1ON���7��|�s򙐿|e[Z}�Pޣ�eù����d���⮓�/v����b����7]��_8ze�rn��:v��3�%v]Q��H�W�����YT������h�Wtzb}x{��y��'�VM����5n�'+t�6�2g��u�܍[��8м��
�v�)�'E�l|��[ջ���m�'���y��*�3D��qh�{�@%--=�#�r[
�-�'{�����]���Sr�s}<��D5������Y�����A�D��Ø3X�G&ݼ��y�9W�J�Kb-c��g\���].�]�42e���e�n+�]o��EG�4&�\>L��ٻ�<��u+*7uEѺ���!��U;Fw�d}��6=�R�*ū�l��;[yژ�kڛ��ȃt�
���=vT�\�V��To�5�;��q�7��B�1ݾ��5e1y�p6�}���y��k|Q����^w7��ΐ%�f����9v0e��+���Ѵ--%p�T��oxNn� &����&q�JX���:�]�Z�*2�r�f�4�0���|�o(t���&.�3w<H���gGu'f�ݷ����x�<��!峆��j��9I�J�@��w6�c;PW^�N�=����<�b�ꁟYmO�y�j��D.�h�7�:����$	��ݨ�G�%�$�[�٦]]m�M�J�x�Q�,򡓹rkv�=�|�4�ǜ�������Y�k0�8
�0>_5OЃ�@u-r�t�O� �)t�hұvy]*�
y��ef�٦k�a��A�يf��j+M)Qٯ�Z��c˂�0�Oˀ
�Y����.�Z�-A��W�9Ə�:��@���#NSl��x���v:�� �ԆV��ªh}�ӈ��f�e�y�>c&�"��Yݹ��Et�11Vګ����%\|�/�����E�����_EC6�8����m�s;^۠䎌;�W�Y��^�D+�y�B�1��t���˅�qSH�㥌J� Mwq��!�e���X��C!f�	�������z�g$�seZ�<�.�Tx%WB�}.���w=����kLg�^�C���e�S��Һw�V�u�\�Y�ᦛտFA�+�m�.{"���� ���<��q��=�B�P��n��ˬU.���*���4�ea�O}�lՏ"�n�^Ɔs
l��຤��b�Q��:i�6�En�S����6��>Y���uWq{%d2��:_B�v�Og�پhk[ў�K|QX���kª�]ܩ�y�G{3n���ͤ&�L���p7<�k�7oħ�F�{�O;��;��2�[��|��]�J
zӔ|�%TV�4�N�i������� Ìl��||�c��+^;�niŁV2a��J�1·��و�\�n�������J�cb�\o�8!�лK2�ͣf�O{�;��B:�>����m�ы�ɽ�������孋g����ܹF����X�
�� �M�[n`�vH{�pJ�E�O�o+�[ȉE@�Q*�Ӯ���џ}�����PPSIE�� �(�)!D��E��D�"1j@F��VE�EX���E
Ԋ؊���1��PR�DF�Em�R�U
��Z����*�
ѩQAJ�dF�PV�Ah�+�ȱE��4)`���AE"-j*6�E
��m�b�b�,�1k+�*�Q����b���Q�YD���Eed�YQ`����T+*(�VKJQX�[j�E�ŀ��mQ-�jJ�Z�*V��E�
"�Pm������%d���Ud*��*V!R�E�b�V���	l�H�*V"���*�+��UUĆ& *"�`��I[b�eC(R"((��d�%Qj)UU��1�2(�J�XDL��2
�Z�A�T
�PW(��+XG,�.*����,Ab��TB���6ŕ��R�T�"�G,�ek%`*�}������>��~}�x�����L7���Lbƅ�+rpJ3��46�.܄`���
c��Aͥ����꩓ֹ)��{�����ɺw��31��k���d����s'b�H�L�r탿9E�Y�N��U�V��Z����9��)�j��$u�j�{}�>*�;�]#j\/o3�6LE�#cС�ӳ��.,~��2Bs-���\X*r]�P͐}.���Q��xmʎͫh�2O\�v`U����9�W6�K�[뻮���U=���^חb��&�uKlb����L~�p������������x�:p=���,n�[�+�b%f�O��)y�Pߏ���B�F<z�-�|T����N��B�R�ݳT�� �Ճ�\#|.\>8+u�w�pw��̰��q��"ZoA�%>�*�P��"�]�2V��|K��u���v8�]Efɩ�I7�����2a�%��RKGG�:���W�
�F.2u	��|ӫY��m���y'Hk���C�����uR^I�kj��qu*��N�H��(O,��b�Y��w�<�){��yɳLh7��+pu���2�ਏKR�m-�g�\]�;L�8��j�,�"�Af�i��6�C��jq���N�G7�(`֕30V'�cvzJ�z�/Bs�ee��:	Y��r�l�TKS��3X��ʻ Dvu����Z]]57�����Nj�;�1/��bټ7�>��L��K�|}ASym��������F�7��oV�ߗFz���c�<n �p�H��(��ǻ+)�M&TG3��;�HQ� �ݨ��z^��
���Mf-��q�Qw�L7��D��'���[��L��9ժ��q��Erm�!��Q��{���������t�w��S��o�'0����*.�/�'������g��w�`\aM�PP�2�]��i�����杹wӾ�O���r�g={�� es�_�
��U�T�,�����.�eÀo
�k�\��V�M��fu�X��Q51s�+$+�a�Q���B�������ݖ�^D�v�]�v8}��Po�V:�h�r�&�Q>��N�X��9
d^^r)�-���Mm�/+y�ӛ|�j�b��n.�P�\�����&o��ݺ�-��f��Оy*���<d�m%|�^����g���A�� dZl��^��wz����妫9�pR�_*=��⽑�c�80�2mS�h�"��@b���ߑwca4��.��yN��(m��^�O���¦.�[y�[���ݽtAj�>
���֯o���$~x�>;�E�Sl�	�w��.���������G�����hX�K�zȺ�\���[��E��p5�,j��>�����h���TJY[�> 
6o�'�^n�t���<Zq���9������C��1R�~E�Y}�o.�v�Nm�ft��{!��h��U�r}`WM�K֢Ze�hN$g�b�H��z�4��M�L�Qٳ�;�s
i����se�h�`��V#�Y��~��z���/��\^{�G���i��ل̔4��ڼ��锏X�h񰂀�����pr�i^�v;�y2��wH����H�L�᳐��k��@�b�ʧ�I�jx�{����a�ݶMS��&�q���g�!���A�ۙ5x'Z�>��A�|��Ӂt�g�;,+:ܫ÷s���ꊟ7��;)Cv�J�S1��>�͒:�P���ˍS���(qW&����vW 񥦷fH0��+�x("���yĵ�Üo�]U�<D_���'���p�ʯ9'���z1��Z݇|4|�*b`�,<���W�o�h��A�Z���F���=�l��]�����Z�B��V�6২�P�S�!�����T�E�܎�_!��w<(?4`Xa�T�q�׍�n��ϵ֑�h�\�'9�i艕�+��F�S��6.�V�n����t�����9G؉ެ�w��k!�"<�&^m^\�ѦTدmΏ0䆬@�y��陁bP��%�_����{���_{k�=c�q�_����"s�n{���?{w:�N����+r7�2&�=K:Y;aY�+�!��	<2N��י�gG���z�lb��]8�t\���cS#�msQ�3�agWK'ģ��On{��e�^�P��_Ybd���3닃��x{6����,�X�{1�%��T���<;��N�E.|��6�W�� ��_��`�|T8+��E�[x����^�E�rH{"�]OS[=b���K���9'�'&K��N�'��2k��
	���Ol�X�n�&����ZS��x����t�jd뇖R8|¨��!�:��z^��>{������Dp;��1?��f[���jP�<��~�/e���P�]��ٔ'k%ݎ�Jyɝ�ݝ�LT����R��<��=(�y��u[�=(Ot�|�w0���y�3ϻ�e/#`�2,��,UQcn��r)��(�c#�����k+��;
��3�ʆNnZ��aU�l����`��J�:�͇���'����	�E��5�'��������.������gL�P�{>(�
�.L*�e>�@��Sgo�W\��9f��mjVG�����aR�w���g�(u��Mp�wo���Z@i�0�9õ�#�@C��^�;����񚄕+c�n-�U��V�-�1��}�����e^oeR�?^�RuN��
�����Cau2�P�e�[�0M�F�`R(�[��<L�Uﰮ7�W���G�zfq�	�u!�����I���[���J���{nF\���L������@�`����i��Cz����(�uywtXX�~�8�&�Ѧ��sm�Q[d��cĆ�����}P���Պ���"J�y�L�ϥv]Q��}��7��]&m��#�;��r��f?,��M���溽s-�#��:�;N��Nk1n���n��g�ywP*�U��K�pv�|/<���T��Ĉ��Yz�q䛥��nE`^V9ٛ�!��E��0�ML5�Q�R�Rb�p�*4�6�޳�/%7	A���O�\A�� Ý8�oM���w�f9�H�2/:��z]�?:5c5"{y�����ƚ��7.�4|t=��C1o�׎��e9�j�JNX�p��Nʼ�ϑ7�t\��HUp����.��P��w1i��B�zJ�y��0ؘk	H���cĩ�^���u��9�fQ�\�ٍ��U��w�7����&�^��nJB�ʓ4�Hk��V��E�\巫��j��/�L�wC������J�z��6H�N��vn7H]�m����CeJr��5��2�Ļ��E�8��i��휕YA�R��磌	|����R�[�Uq�uN"((P:(!�G�YL��P�T������s�����7��-��`�5L��ꭂ�}U\f�M_T$�΢[+��'P}���E�:������*]���f��zkZT0�l���qGu?6:R��3����D���ؽ��`x��X�A�}�o�kN5��`*#ĝK�Dk��]��eFn�#_gQͪ�����=��a��YeoI����tR�9�@�:C��P���v���鳝n�X("���x���g`�F@���+�\��d���4O����^��S��yݦ]��Ȓa�!5{�L�;��j�f�B�tJr��4�c&��Y�c���K�6:�����f|��GP���V��0ۙ0?.ǈ�a���ڑ��ឡڠ��nb$��#��^Z)4�дg�_ݬ��+7ۀ�cB b^=����-ߑ�u|�D@N�$�d��S
8C2�N���
��.�c���k!�(���8yJui\Vp1u�Ô������U�h��z�y\8`ή����s���"1�7�4�+��\�����FZ-7�^Wgc����p�i���1y�t�o�h�,��=�5��ѕ�Ec��R�q�iΧn�F��}_|���:����QM��~뼂���'J"�QU���c�l3L��f������Q�u�����C�k"��^�93�[�ѱ�#�bz�J�~���[��W�ey]�O���[�asqd��/*��v�]���"�=���M�{����{�e�Bφȅ�G���"��~DA�K�p
��0U3�X�N�Kkk�1~�Br��3D�*�{���~���řk��>���*<����Mx���G|�BM�:g��y�Q��y�{8�ܗ��`F��ǒÐ��_��2�Ve�6t�*p˺�qu��]�B�)pT���yo���u������I�'5Q�q��o,�P�WKP��h3dm.�J��z�KWO6ی���^_���ڣ��~E{����E���^���>�H�˴x�A@n���1|9��􄘙2�=@]t�k�>��^,�{f*��
9n�z�L����}K(����5��R��Q��f�\�"�4��m!׶�j-y�WK�>W�r�8X�C��H��̬v.�V��.�kITQ�oʰuα�f�w����N��T�����/w��a�mi�PQ!L��r��ƭ�{ ]�܃XV]K&{f���	Bs/�Cxt���:�k2	�WuM�C�u�J�R�srWV��xf�jr��j
l	�^��W�9��mfK��>T��#�S@S.5L�W�w�c��s=���S�]�YϦT�0 ��\��\�9�o�]U�<D_��$Ǯ͗�t�h��;��2����`�Q��b�qB'��C>�k��댺�g��뜘b�."��7���aJuj�WW�e�/�h���OQ0�i��yQP������s2�qqC��jo,���/'�<��Fg��'�D��=K��E�׻O���϶��F�R��G=�_ ��K�����>�\��`}��9��XY�Ov��^ksG,�����LS�,N�p�����Ip��&��`s`���̣7+iLI���S�q�~�j���}|�\��m:F9����X����N8�\��jM�z�<n�c��~�[(`��;���Լ�/%q`��=tA�w�����w�C$/�:�5tx��[t��s0�J��7i�뇼z��D��
�T*�)Es�^�ҸDy��c���c
q4mV�޹�뢱D�Z!M �}k�?-=h_J��&v2!����(��+��N/�V�U8��čQ���w]�a^�pS]Y.���I b��t���6�%����V0���n C��u���==}���]�x�ƛ*�oM��&��g�T-f�f:��u,x����~�=)FF�W�TK�==vf�}�ݣtd����PdX����J���K&���yzhM�*�U�=ˮ���l���ߐ���u(���Ē�TF������SW�Q�#�K#��
��ȷ��i1���2u�A
�1CUT��E�qqe��T}���`��m9�=k���6��`��ȹ���{a�B��|��5���Cau2�3�*��ȺUs�]�V�]��Cv�+����suq����	�BX�.�w�~�������k�)�p7�f��]OE���ڑC$wB��cPޣ�eù=d��#d���y��Śj�t���ْbX=ҍ�;���Ź���Y�c�FÕ�%S<��тP�|�s�8*��~QrrG!O3�ߩ�j���GE�KǄ����$��JD��(BwhF�ɷJ��$�n�f��l\�޲tؙw|�K�r$Y�"��-���p���\X���C~�u��n��D�
�N���w4��u���S˽�~4�ѷDg�������8:�h���� +E�:.��m��f��s�v��{���?EA�[�OoG��M;���`5����`z��J��О�0`��}|�jݲ#�gp]-����-���<���0� ���^�G�ڇ�)b��j�y¬�>�ˑ3��ә��{������鄽R��Oj��(:e�{��o�^����JɺA: ^���?#�cGb�?Y��_Uң�ga�qQ��Z����C2Z��г����t՗?/����sػz���&�P��#=���P�"]���z�zK�o�X�=Ǫ2���yy����
�6��3<j�ʭ��T�5��B��63h�)�⿝ˇ Rߕ"�̓�\�*���R9?6F��R�Ғ��Ė�J�����5�����uY
z�S�u�J��ٺ��.; �l{P�C�U��K�Ckj����r��D��n%GLWϻ�V�{�+�v�=�v3mC�a�W��,�҈���^���Y���gY��m7�y�l�[9&b=�����E��I��0>�eע!rF�*+�w�H�ܩs"{�4�w���͒��C�B���^�<�}
��^��`��l��E���zN�;��YPf�j�^�e�<�7d�2��z��h&�Үc)n�A(>��a۬�	R}/r�ț;�d�fL3�!^;��k��{�by�OC�	����9�Am����; >ԋ���+G��w�]ҷ ���˽%-.���0�v��p�p38{<�֨ɮ�%����۩�(�\���7����B�ѭ��d���ԁ�{���o�������i�o7\+,Z=�˽/tad�P�T�.q�!k��:�����.�:y[B2,n��K����Sn5�:d׻y�s��f �6Y<�t�IDJ[��6[��XVCd��F���S�"'k=�z��s��<F�
�/����|0=�6�m[ӸrF�xn�A�ub��_i�������h��Dz��U��X�����7�%���;��x��{Mvb� to�;�t�6raܣ��Υ�_2�fd�5+��n����3//ֵ�!�.���tw����#p����֊n�p}���	��]79|�j�����}g,�{t�-�|f���>��4c����w�Ӏ�7���ʇ��Qe�����ME<7���/u�HGRI��^�5'��0��<7}{肕	���oVܫ�#:�C}��tX�i����5v>n���˾�|����ܺ.��a��^�S���iC@ۊ��/�(B�f��-�e�T�[J�9�b�¥qի�Y���$��*L�h�h����9�g�]����z.���<�ܳO�}���,#��g*��dsp��Ų*2�IR�=�������Y�6Q��sɛ�R��M�V�VK�إ�r'��C��v�2b3C��'ӻ-Mqe[ϛ�~�L�k:��V*Y�z�$'zU�ά�t�N$���c�N@�ޢ�ܜ���f���Yf��"쭖�9��-UǗMAȴ��X�jB�Xu�2���2H�mm�7�r�dܝ�;Km�y��QT�m����W2Mج%�x��;q�c���(6�f�T�w���]�Zx���Dk������â���ߎ{~}_mn���}��f��(�i^�q	A�P7��pY���2v�pU�Ҝ5�\���C�xot?�Q�;���,=�X�I����<��rG����Q�6�l��ج�2߄i�`��%ߣ*�Q�4h��38B�9F9�oA�X3.j~�T� �nAV��A�G���r7J�v�}G.�����LǶ�r��7�:B��,�T�ge�{�_up�ċ�Ґ@�ZV!ݭ]�åGd��צ�Ϋ���n6���({l*)��Q�K�#�eN�����RT���͏�c��q2�����}�7C��10��;"c`�납�jMx�I��(��ա�����"�_3 $	e��i`ǭtce0t.>c|Fv){�9�F�m�+q��������⋨2v/&�vYM3߼5��ݟ�>�l�B���
�[J�PE���
�D]�"�`�RVLE1Hċ,�YX%dF�B*�AE����"0R6�����X"+r�cQE� ��ڶԘ�DQEX�"�XVV��m��Z�b�V�
�1�AT,X�l��Q@Q1*�AQ-��m�%"��%Tb�+%aRDAED1��%X�#�X

�*��U�ET`��1V+d�R��Y
�T���* �a����*媤PD�-QdX�lTQd���.%b$YTb�(�ȫB)m��R(J�V�±E�Q�
F�q�X,PQdX� ( �UQT�$��nR�x�Q�j��ϥc��`d��/`��ip�I���Z����I��ٴ����<�_6�'r��_Ͼ�<�I���Qu�?�yJ��-��5�����&Y,�HY�tJr��o�<sέ���m��I�n��5����x/>s �q�g��_�Yk9a��LU�{Q׺�k6�\����Pg��M���I��GY���RiQ����|`Q�ir�CG�R� e�e��z�w�~̕i�@�'Q�U����(>�.�ӡy}�/��4e��߻�����+֐pu.�E>�Mht#D��'zQ>��N�Y!p���n܎3��nQ��e����{G��K��m��*6���T��G>3ԺW�=~��>��%osde��;,%y+�%%��^5srJ��=V��/���-t�xcң��)b5VV���vw8��pCG�ΊU"6x���/2}n�Z�bN�c*�9~Eݍ�9�x��{�	��+�d�2��k�����\8T�t��&x��s�h��g�μ.��`�ڄ�k��g���ݽ�׽P��z�-5}CҊ�W+��S*���+�t��+#��>#2NZ�%����۪���3U�P]��{�e��#~���;�2D��/Z�-w�>c�xQ�4��|��Z�����/E-�Eӻ��й�'�ǻ5!������˛NRx#�#7�3nF4�O�Ýn%1�F�0��&t�"����:�ig��C���T{\tFkydʆº[ �Ƞ��@ڞùUDR�gaQ+�.q׏{��gL�i_�b���L�CH��=�u��Ͻ�͑��u�tD�g������띏��3䬉a"<�:��8�Qcg!C��q�ޱQeS�N�r�==���Ñ淑�9�j<`�4M�Q(3H!��崇Xۙ5{��Zg�y
ک�8�F��*�+jq��q]3�4�$�p��tsԻ��:�r^��W�T���T���B}Y�C��s�y�eƩ�s�nEz旮϶�p�ep��C������3�U���S
dҧ߉q���<�1��[䧧�N�p���fUS��`�J��.*0A�t�b�!Y��Z�q-q�OO�x;0�=�Ok�$�wU���g Ϣ�+����P�4K�v��>k����q�#�Zk�,_����_h�`hN���[]
����Ff��J�{�ѳ"`ۂ��҉���/N�,��ɬy�k+�C5��\����](7�ۜ��E�dtͅ�Dgzp�
��vsxb���i�ac���Nt����D��n�b��둾�;���v���ګZw�#W8֐���*^�T39"2(��gKz5���Bp�a&C�5K2nH�aHN��m�{<�ǯ{���q��ق<�\�Ε��8�ֹ�5��A�wC}�lɏ��AP*������.�A�n�=��z�`:<�������Hߣ�m|� ��k�8|tnz�0a5��Ǻ��0."e��0�\�m�.Au���sY�L�̵/=�MӟO,��L7f�~3�G6tU�EZ��<�ƭ����۔ߑ��P�>:\I�[1Ի::P�!�9.wV�뇖R��V<0���(^{��^y2���i��%P�48@�Z8���J��3�K�q�S#!옽��Ь�ݬpm*ʼ�ԋ����{�Gx�����T4�弢W�F)��Ɇښ��U���,/��Ͱs����{�ɍ��q]v�I��Ȱ}UB$�ܭ��9��Q�G|]�٫ZޤU�vɺ�2G)��pC"QC]R;��"ł���PL��vmvS�W�͎��_r���F�|��޼7>�l�,�4Ht��:y(|K���-�����'��<d��|+���J[���(0_��h���j�B����*:�ܮ�}�,@��������#G7S��Л$؍w����f���$U���Z���i����1˓��l��ыmwk9����10J��W3�����T�J9:[�[�{���;�,������C��2�i��9��s�y^���^'�^䁓�noLd��+�1����� �~�҄L��]F��(oQ�2���z���˩㥟qRW�����q � ��ݯ1���NE���y�ht ˶p3����U��v��E���;�n�L�ʿ����S���٘`���3|���^����-):�Ю��~���]�mڲ���ʜ�c�Q���YPE�;�[�:�!@���[۵<f�ow&o��W��nW�Ժ#���C<��`�'ګD��ٷU�;�2u>�|���r�׌�x��P�-��m�BH�=}�x8�L��^�����#,��`K�ٟ"�=[�՞��.2+%�Q�T_���c�d50��c�s��C�X#����GH�κ�<�̥۽K��tE\s[�#$�d8����!�L�r٘��->B�zJ�c�\Or6�3����u�˭�X*ۊ�~f��Um��
�I��0tf��p�N�P�+��d�����+;/�����q�
������JK�Z=)�ɯ��lgQ-�и�~�y�����5x=���M*6��ڹ`���ь�:�Q�Me?*k�.��bR]��>؍˯�z��s�l�hٰ4�w�m�����]{5�h1���K˝��|�9�!gE�������uA9�z�����S���2��'v�u��:����r�F�z����{e�U�{E��ֺJ�,�qxt����c�5��fp,i���7�D���)p�.�ǹ��P�Xrq�6%�Q9�Z�a-�R�m
��1f��n��Ʀӵ�F^�z^3��++zLw�5ye�G>uH���z�lЦ�{Y����F��t(7u��|"�r^��Y �>Y�et�t�Ƌж�KK���ՋG(�����l�|I& G���6*�J:����=,�HAȫ��m��2�;K�<�����~��k={���[��Wڕ GVz,��>��gPf��6"��eUf'�Ҕ�w�1HȰ�A��',�z���Y��H�%[T�Գ�V VNC���i�	:Gl��=�P�a˶�����&��<�Z,�����]����+zݧ^=�K����m��7՝�3S�zUϦV�F����I�҉���b`�Z�K�����������ǵ���Rⶹ���\!�2��ؚ��̬��s>#̈
����$�Yx�6�/�,��W�P
\ľ�xJ��\9Nc���uQ<�2ڛ��:����T��^�^�ޔ���߅��K�e�)wc�Z�ULKV�2�ǎ�8���˙3(��'wۊ̓W(�iS�uܴ�s�\���f�(L��M
��:��wٞ�p������φ�v&<7,lXdZl=���gѡ�{-�/ϛ���R}�ϫ�v�
���_%�2R\0�<�N^���[�������2��J��ܥ�v�akP��[�i�������
u�c�k��v�����^��s�����ldDnK��g�c����9�l��#%(ϋ�Z)qh�>�/=5�S˦�w.�ºdC,R٘�b���c.��'�����f��L�{U�J����4ϵ�L����Y/%l+�EW:Khpp����%�2�lϝǇQ�B!�};ݲ�!rb��������|`YZ����$G5b��}N�]��f�l�a߻�ue��9be�
1c�f=QK�N|�e���D�J#�Wm8��v
���"b� ���z*�-��ɧ;�4ΜW=�d��O��uͬ�PB4��t�V*��eȽ�A�΃�O'��Wz�82�7�t��Ǉ�/]a��j𞩈Y������49�-+�8F�K�9�z^O��r��
oy�>۾�i'|yT�,&z�D��Ō��N�wO<���7ْ�pyJ�����sՙ�}dO<d�͌of^mӄ�d�Q��՛n�UT#J��ȇ,�ȅ�tx9)֨�t�G���3��q��ѻ��RnzXZ����nM*8�%�([�3��~��v{����w�C-h8&T"�
�yi!CY�JL蘻�1��]��|�V+]uy_�p��r�k�W���aLP�U�N=D��	TD0Fe��q�k׼����·$���M�܃�:����o;�=�՜Z`��
z���;F�H8��fh峳9��������!�Y)�e��/x�q�Nd�I�) ��makQˡ�SU��\���C�fg������T�A~�x^qpu/$�{��z切���Jw�Z��ܞ��4���!�(�j��-��8�T����o���}0GX�c�㙙ť$�!�\�]3�����*����C ��;�T��3�^��}�	~1�ys�`��ܼi���n�%�b�!2v�����E���2ȿce�V��p�b,�,tz��|�Ž�qh�hZt9 �D�}��Y����#22-�9�pހ�'����K; ��G��P���mL��!0�ysQ+ΌQ`�L7�S�5�:��g��o�;�ܳP*(�ٓ��/0{x>���|�4���k�������"N��	����:�p>����q=E��}�Q�)�{��r��g���I5�ՓS��nѹ4l6wJ��K�\!92�o)�uh�a���X�r��2���4����%�=�ضbdW�N����-��Z��(h��ʤ��O��+Z��\����:o��Hu�E�S�z�2�n>�j�5��G	f�ۻZ�$X��qq Y��촢��������o�	�4��;SX��x;��oMw��t.Ո�U oW%���4�#~R�������k��^���%ѻ��d.�������3�x}=o|p���[X5����I�I^{(��.�T+�^u�P��-43��X��3<{��ű�\��eƢC��ܚ�Ǌ��l0���	�>6I�JP��.������r/N��gI���+"�]�U,���q�z^<{I�Njq�$lcvL8��*b��جRge�jgG�j���Eoz`������`wb�ʵ�j<��
�'D0�B���``�K��>�����{�����qc����.�D�\yEQ��^`�P���B
u�vg9�t�q�*r]�]�+D��A��.��v�{���=��VJ���nc:��!s��!iq
xb��
���t�-p4A��Y�l7��o	����/�.)���4q
��>9k6Ze��zl�)>"�b�qa�瞆`�� �v���.h齂��~��L#Eir��v��Õū�ɺR�R�X�ùl���SVr�����M��:9�a|nm�ZGA�*Lti��78�1��;K���Z��yC2Z��
�8io;B���:��	�����T���:�I�`�!�A�L����ZY���(~��. ��{CĎ.��V�6o������VZ[J%�삅|(0o:�Qe2'��x��׸/-m9�`O�Բo��>ۡ�c�7�Ҵ�M���4\�h�"A8U�l��ˉw�r�V���*v��fN�1�oWh�������R%ʋEqb����ʖ���Z�Ýљ��1~�(<��!�}j	�yYzV����4�$�Z�������z��b��[%���W�\e��e��.k��aޓ�M^A�Aff7��s�0���M9��q@���.g��
͞2��E���q�zY7;��{���P�DF[Z��w�'�=>�Y0�xh�)k�8��(8�f���TvK^��j�	f�Bueҷ�It��t�Z��u\��y:g-�����
pD�H��I�b��ԯ���g����IO�$Ό+{l�,��,��Nb<|�;Ӷ�MbJx�k�ք��r�7��ay����b���9b���$\OkN
&�~�=�O0�t�-�OVkd�{E��Ի�1������<zY�����+iE��Ab����S9x�=}������+����%{7��i4���,�H�Nb�ƦC�v'�=%}�Du���R%�z�ry� ��N�s�1�1���_|�� �=~��˶ �<�(�[˰�i&x�iߞJ���*#�Y����Kʭ��z����)���*��Հ�F���� �u�]�g��;�W�v�a��[�&G4+�]��3o�m�7�E�ͺ�|;��^����Es;d����;�H�,�"ލEw]�)_��:�vd���nE�a�2���bv�N$F��^w�1"X�d�8�v��Z�{T¿[��G�[�JK�痄�o�6�-�#�eշ{��[�`�~z�n	nT�=��r�cѶlU�f�]*���b�6�!\WYո(��H�é`���..D_�҇~E�C�����p�F�Ֆ��GMX��R��=�
oI��͛�S�{ʨ��`и)��1R%�z\"é�#*?V���-C��j���QtjC��d�kr{��#)K�C���-+b���L��4���yv�*���fWSo4��r�.��ݤ-}�h������O��#X�5�	�w�Y�;=v�}7r#v/
����F�#MXx��f,��^�����jY'J��o7�	�_?x�S�����&�g�o�W�=�*:xB:��1�(u�{^��͢��Q�VZ���$�a�L�iܰ���N��ϱ�M�Zv�Pj��� ]��ͺ� E�	$�f�����!����9�C��l��)td�wg���0Vr�U�PL�(Å**�hT�J��5;��$���0�ޚ�Ԟ���բI��y�^�b`�횢���P�`����棷\�-�ȴ��@�XB���ݽ4���	��|�L2�Ë�_�"ya��!St�*��]�����v����K%H�.�]i̬�������8
�+2���`���(+�}���e>������O�822�E��{��`ɔ��t^�n��B��GA�OJVЬ�cz���P�c����T���0�b��u�Σ��{q�;�)����
�;uh��,ī,ڇ��P!h��O_�-��I��u��}m��Q��dais��Ф���d�j��p�zt�b�$WP-���Lo6���('����6�	��&�)wm��u������\�WA]�"�lg`�ɍm�w�wQJ��x^�|�S�C�r�ۊ�B�N83�����!��sǊx_2�(�QI��+Ȑ�XO�Z@�\EC�%�[��{l��E6t4}�J���E�ʒ�Ү��$�2"�Ĩ�ɽs�N����^�f�5{[����Xa�92?.�x�hHq;�E.dy�,Z�9�%�:{�$=��z3yԨ��;�)�3[�s�����R��3�D�������7eQ6h���r�z<�\�	+�D@�[}EA��cۻ�[{F'3,�����2��# �3.Z=pͭCA�<��u�2�\�.`���kv����&�89��GG+�5���l��^��BO.�x�C�ꘋ��1��Y����7!�\��3r�G^+�*v���	���=:���"ܕ΃<����$��ԉj��}���P��k�7Hc��3�^L��<`���M�NƇ���dD{e���׏�ꈽz�Z�������/o }�廃��9����P�1�w�>J�熬+�Kr1xƖ�T�r��0�OZ�&��2�U΅�[�F;���M��F��Xx�*E�:H��r���e�*�Ǒ+��;�c�
h�I��ы�0�R�p%CeK�=��a����)㻏O�A��]�����E�=�C�(��4�2h�3���<i��:r����j|%�B�]k��GbӚѻ��b8z��I�S�|��6�i5e�%��!Q�Αlu��Aiʬ.d8&Թ�֒==��Y;��I*�Jɟi��eہK[GN‎=y����S���m煪�E����J��@QTr°�TR-C1��H��(�"1�UXEV,r��ʠ*�QjJ�-A-dX���1�"	��
����0X���FZ�b$�+k
�&Z(9aQQ"��3,R�,\q� �c�bU@r�T


�[k��1JȌ��I����(�T��1q�,XbB�T�%q�(�neQA@QL��%��8�̰+*��YZ�E*��k�V�dD2�A((�V��j)V�j����eKn!Z��U�	Y
�*T�)D��5��Uk
�D�Z��Ա��(�D)��nS�7<q�u�Hc��~c9��dp�2��s����t:ɸ^�}&��y��;r�A_2[�i��sJt\��E��tZ���=Wv�d�k��v; �x�Ӆ��ل�d炎��t;����~1!��R�+	Y���<tK4M}ΔF��	q~��=�D���f�'%ܓ��Ԟ���Y�^���l���zJ�gX\4he9��nd�@*�ѭLmCz�^��wirҭ-���ңT��Ȱ�9��s-<&TłxPn���"ҿ��.��{������^'���Y��1�[(�Xj5�T˅�˶w�(e�&T �b�!Y�����S]ر�����vB3/�zY=s�t�T+��o��/�2��p=G>Pù��[�'�����)�#!OѿR뼧��!���ۑ<�ȸs�Ff��J��jȔ�+b��*7���&߶{8q�� V]�P����¦��][��D�\O��*s'
O�H���G;�y�����+�7��dXY՝0�7��|�����T%��/�����:;ץ�(����ڴ���,n �cK�y�J>,nm¸,����ߢ�p��#G/_������*�[�UU�m���;5L��ܧ�E#����>��[�&^#�b�Rg �k��z_m�wF���$M5��J�2c��WsJ�D���Â4�)R8�Q����gU���=眩����%��#8gK7k-�B;�]]5e� �䜪	�#&�vf;��K�/����_�i�l--D����}Ӷ�zm�ٰ�|����IC�矱v4�]o�2��k8*0>.$��1��;�����unN�xͅuU�>������6��ٟ{M[X)m�Z�Bբ\>�
e���U9Bԡ�_�T�9&�qO:�O�L�uJ�8z:MLtd�R��>[j"��LP�\�Jǝ���a%��3�W�Oi+��.��rL1����q���3㕆��[I��U\f|�����C��lR�y7���]����$[]l�#������P��mj�ԋWPLͺ��:�����Z��>�0�Q���"Ļ)��`���v�ye�av�DH��@֮JWBXKb�+k��"�-l[+!ۥR�	��fU��\�Hq՟�3�L�k�8y�+T�?a9o%F�=��g��R��y�
g��r�8&�M�,k2�p.�->Cz��<^yG��x�q��{�^;>�Y0�$�ޥ�_���>Z=ܮE�:�Y���Fܬ�3x����*�|+|��+j�Nݝ�b�
w���t�#��j��WN���-�+5�5�1�ܱe�2,v�`b;\"�VRZ�ݹ'�룙16��s�Wpp���]&�Y>7�m9���tg��U�r��Ԣy L�7�	�N���`峯1&�ջ��&ĩ����'Y��!�eم�H�GZ�L�ϯi��f/����Men{�/:�V�e�
�|�x����kþr��s.�ϟ�yND�>��g,�
I�������z�=}�����!����.�}
�,0l9^i j���ߗn��{�]�(�������<�퓹4M3�ۗ��u��L��,��i�L&�y�$�e�+åo,�u���p�}�V�W"����������8�+���"��u�ݗ�`u�8�Ӆ��|��x�^�#(BY]�9�5�
뽈`�Y�1�䯌>U�>��S�I��������-3�qJe!��)�F���{Q�S�-��+�a�q�--�4UC�dW=�E��<���<���\}7�k-v�Kkn��Rޡ"���Xdz�Y�{R��Ui��\f�r�7���GIs�7��S˻�TYv��>ˈI�' Է��4=�W!ΨU�K�H����}�w�d�dwn8�kp�c�͢X(��t��v�A���Q�}�z\r0J���|��ʢ�`��-,��U�rl]�!'{�߸��o:GY���ygL��F�+}�=~t�[3k�y<�W�e��B�	^Q܏ú烄�g�gq�պ�̩8Nwj���˱�8����)lU�[Z������u%I�Pо\�3l��m�:�q��Ry`=j\�o;z0�p��q*����g9sW���=�����VX���󠌉v�2�Ffu��^ᶹ���7�G����'y4ރ/�3��/g ��ƨt2y>Y�9UX�d�䩳$�U���j�;��d������t�E@�\}"�r@��!X�Q�/=M�չ��Ҳ��Rv䭞��m46�/�$��s���C�#C�&��2:���Ϲxs��*8lk�/?izx�z�,�%�����;vz#"��A�!��¡��Yґ~X*W[��3�����n�n�-��gt��w����4K�.+�B,'Q�FIVHW�v�,��wvO}sͯ{s�rtOc�f��ו��B;T��Ev�&��&��=91q��t�°s9fk�R˽�;C��nG1·%Ydf�#@��-N��S������4|�Bk����$O�=��1�R{wXt�K�l�������R�J�d[V5W��JN��(�uz�7�\��P��*f�iQݾ^4?���wh���-�%%�	u<�E�lA���E�z;�S{!ds�x�t�W>X�eu����1>�pt/�jUn��(�*Q豝zet[���f��!���V�K}B�Ĺuq0K��d���H�v[a�/�-����rY�+)7�l=�V�����Nc�1�b�I�����F\(��׾{��s0iq4��%�ܷ�{|{��x���k�%c���3/��޲�����Ȼ��>�
��z_Iͺfc�x#2��W��ͥ��<>wB=~��de�Fzv��C���j��U��Y<��VH�z\"é�#*?V�#5��	�]z�*h�f>�r��ƻ����z�N�*�<w-+��l�e����i핲/�*1���VciE�{����r���6���!�"9�������K�f�f��|�׻\��^�)S��j����FF���D|
����.��Lz�W��W�ă�h�+�.��#�����9�A����3b��i�wH�D��cYYB]x��9,����d u?Qʍd5R�ּ*e��iŚ�)hY�1`����49�-,��p������k�Z��g"�%C8Șd_�sb��]�/��gL2���2��d����z��'һF"ڕ� 
&��W����=����^W���aLP��V��K���]_���.~�B��^����r�:�h��1+_�,o�2����Ʒ�wh�q�e�Q�s���הy����C9=�]B��Ȥt��v%�H�a�Y�׶�:'�nԉr�Y�#V�����`��2�c��hQ���m�F�͓��NiH�����Pu�Pg�vI/�M�[���۞�*P.��RB�jL9���MrZQv��v�l��/-��4b4�0���s�=k#\/��*]�_���F�8�\^#&�[r�ݹ��/�(�N�8"�ά0�676�Äav:��`U�(u�zR�����������r���|%[�WN��m.�� ��P0�60<��&Z�k��ҹ�m��{`��g���ͩ3�E��|�]�{��~��v�L����~���Nۭ鷜ke�p.[��t��/L�lɠcՀ�m�<��+Ш�_����l�w3����,l��O5sw|�'۽{�4�e��}�rW�ҫ��[h�$#~��9��Y������S��7�u�a����#����F�8z��1���S�P�,S:�5�F(�Xs.�l5�bݗ\�稚>;��:��N4=��I�D�@�:8���t{�$�y+n|������x!-{ Q4�إzB#�Q�#떡���a�r�uKW��E�+����OiVԝ^�[����p̰1��:jլ������U��*�>�q[ä�a�-�NEN�Zq��V��h70EX=�f��lZ����V3��%s0M���sԼ=��a�ۨ�!o���SFGB|V�.V|�=W�&�E��u #Z��׍�g9;�M��ȘV2H�*�{Z!���f���/Z�,�W�D�R�9)��mu���lf��>:��Z��*c:�)a�p6,Mь�[��&��Gy��xU�
���"U�,����5�,5��A�CQ+���L���r�3e&��6�4=�m����a#�zu:a�]�E�3��G�>�၀(�r:�{�\��}��[��
J݊����ծ�F��*�cyZ�.5�0eWd����8�6<'XD*�¶8g��x�?���m�a�4E�J䚮V�l���2Bt�Rd����y3�|���%ߵP*�_Tܬ쨧C+S~��\O΍U���V9�{�'`�xe�7�� `�3�9����9w�h�N�ϴ����f�GN���U��g�V޸��P�,�	�w	!˧�/j��v�m��,�T�o/�x�A	�U���(qъڳ�mH������3Cv��/N�}���5���aE�>3�m�C��ǥ%~2/:��:�Oi.���lPf�8s�]��qo)�xfq�u֖�Z�x�������x�^��ئ@w����o7�-]1l��m�I��(Ó��U�ϰ]pU̹uۚ�p�����v��(:9�G3�uU�i�ƹ��i�u8>�p{�r.u8�?i\����d�C���,�p���M2cr.�fb�T�� }��ѕO�ŉ�
���&:U%��%ᄹ�T��"1p��\����]�&]d��v� �el�7.7��P0����ʐ� _Vf;�揇x��f��>~���ݓ>��2NDK�p��:��Է���͍��A�@ꠗ��8{w;#R��Ξ�N=kN-�U�X���~(�v)86
��;$�3~
k	ƻ�u�<�<����r|w�aI��i���%�m-�"��N�,S�5x)�{}�n�Lm��޽ꌘqp|=�y�[��;��R>���(!�IsS(P�ԙߝ�����:�)cH�O7���#�kñ�<d�sص(s9���=�i��s���4M}Α&����B���o+
�v�e��|�v�*I6'�f��lN��!�96�;��yn.,<ໄB��<KK�j.�p�N��ι�.��D�$� ��)�sʖ�:����e��qX5��	�P��)%])���,�+�A������f��g�*ݯ5��j϶U% j^.�8�G��2J�BU��H������L؁��o0]F�}`��GG0W!PMS�1�y}�}Y�]�I錦��/��kX�u��7No�-���������zy*�&^�ɮ%�o�V����6�mUo����Pȼ׹_*.���ҵ���^�7��#��\7��k3���ʝ�8x �΃ A��v��^V{���{�şoK��K&�Ѝa�L �\���/�<9l�΀g�"u�����vY��܃��"��2��S���^��Q`�w��W���w�=��Ȩ��>�s�[�^�oZW�JK�;�nE�a�2�6DE�+h�[OB
�wq�N�k*f��Qݢ�lti�������%�dK�<|/���Q"�x��j��ZYTP�U8^���.����{}m��E�٠n��F� ܴ��\2�ʙ�n���7-����+6��sGθ�Kۦf|�^	�z!"�^�;�VZ����Vx��qh#����{~z��6���Z�S+FT��9�����p�����5Q�q�#5���fM*�`,kR<k�Kݤ�df�:��V�+Q抬������ĜB�=�bt2kŵ��d]%ל��zzׯ}���O�L�zU#��M@l%�K�����>{:� n_�Y>"��=��ѝ�SJ:sb*��b����	�g�閏��(�����C���k�꼤^F�.���MK��gE`�iu�|�qû� ���s����`�/T�"G��J��N�8H�x�AR8�ĐܝYo7b�C�p��g�{��[sX�^�V�N�:W��0�#��24�B<<�c�V���|=u��L�ذ?fú@���D����i��
�si:���	���#o�=���p�^��でj𞩈Y�&TłxPD+2#�.�[=������Θ3,
u�͂z8�8��o�ƹ�	KS~�e��e�;����P�a)�Kw|������(�7��夅��L�p��������^kC�����ϲM��[��:�{���5��#�;"q	뜩]:l܃�Y׎tr��z`�+���yku��w��r��0o��]�����k��E��5���엵\O��7��V������\J�F*��%��*��0a�ϗK'��m�:�1ؚq�'�8����כ�w^媞��'c��\�9�@+�#V��n/rԧ�x��ڇF���y�}���#{���oW���oŵ�kJ��A�x�ՙ`v^��˲7�e�grђ���;/�'��'�N!3GY��|�U�܊�p�,.$�-���a��E/�����ڛ�t�4$���)+�n�;�1���P5�k!�Y������D��(���fg���i����e��n7LA10҉�6���;����0��D�؎�v��z�Mj�9�������
�:��w��觳r�L��B����}��A
����Ю���]Z��*�X�Kڢgh��1��3֛u//~ݻ �36�eGCj�:�+5ٶ�X��4;�]3ZQ&�(:����|7�XxE�]�d�R���銻�Z��4���,hH�o����~=�Y}��P���ci��T�ׇ�a9�,���o�f?�5��6(;#d^����tz�R�Ӧd���
ʳ�s�Mx�Iԅ��;4ܛ�\���ܴ��	��ؖryF����2����8W��@v���S7�b�i�łY����toTՇݸ�`��D���x�\�wWo<��D������Q��j�{{ܽtw�ŏN����`�ׅ��!ubg�:��B§�y+fȼ=��sE���"5G����GC%��'mN��s:�Y�X��k]Ћ����OpaڽX�
��)*�:�"N���5�۽C�ED��7k"T���q��/�pHa3����"���سd�~�-�ڰ`{�8b��7��^Z�L���E���FR�>�m+�F�i�Jެ�jK��w��H6��r�AQ�2���_��M�1�sJ������7@����儊�K�2.�}nC�טͣ�iA9�:X��B��f�������( �&�Եˀ�(!]��yo��-,4�����P��߲3��;�$��F���k80���Y�R�a��Ӌ�����s���#�	��ʻM�6���-�q�r�����:I��]��9d�q��\�sőݺ��P��:{��ǮHs
ں������ګ�β�Wi�5�g{��R5d7x��.m��:Kr>�Rƕ�'h¶�ոWj��j��ɿp����>.�m̐Ã�L�����&�D�|��ܰ����l�i�����q:N�KC�^�T;d��t\E
<�r�8R�#ࢾ���\ɼb�t��9pֳ3J<AA�hgR^{�;>� �d��G��C�v'	�{�9�t�¯h�)2��E��oнL��uT#����7�
K
��ʵ4����ru�S������.�5b�<���w@���d�����<┍����ʺ�A��m�}�zMJ�P���Q^��A�"���Z�j��j���`��0�3�������>��r���>�d�'){�m�d�KN"�B�6I7Q��/o�k;c{�8w8c���v����{��$��U�)wd�N3�b�<��3�9���{f�$�ӄ���n\���r97���>w;1��!�YxZn�ܸ��"e�k�;�2"�=vgx��v�g��б�2R��Zn��W ��=2��j���T�Z���QJ�e�F��
�QF�,EeKYFV+l��Dh��6)UAa����IX)Y�\`�b�L$����ơ�J���V���ƪ��m*�UaTB��2U2�
F��X�e�D+X-���PJ��U�e�*��b�m�R��(�*[qS�+���(�ڥ���+DEj%(�c\C�[IRT�8��R�`�Y��8�ƥ�Zf
�e���-j-�Z֭cmJ�.%q���BcQ�VT���,E�
�,RQQ[Lq�2�0R��Q�Z�
�V�2�Z7,W+m�Vs0�F[-��-l��j)Z�4o�b��� P��^���'�Vϟ�)�T��<K;
�CMx�gw���}�%�)�&���=#��4ԙa�2�)�0!���nY�;��I��'3����,�p�Q#�C�N�$# ��%З��/��f7@�qL����)�ۯ�yY���-ub{9����Ϫ���T8��(u�j$P�5[���-�뗌J_�.�w/�z�L�����Cۓ1�8a�7��M �2$���'5������\o޿w"�����<��b���Z�k2q�ȹf���ݭG�,N�t�h�Λ�3��e����L;�B��VS��.99����Z�0�W�D���у���>q��u��K��&\)��J���"ьb�^�MQ��l���!�.g�)�yX�2���]w(%}�!}�j%t��A3۝r�8&�M��u�Q��5 *� @(��;�z�gH����xD���d��8?�0�t�s��!t�3�Ks��B��T�Ukn�c�fiJh��YY~�s��o۱	�dt�˪0�)�ؑge���"Zs��t�~nLf`v��z �O�X�=��r��<�r��be�8�K�gQ"j�b,Cb��NP����x;j�G�%�mII�y�0W<�!Ө�.�ʱ�*��si6���~�WM����2�[����.w����gk�`�����=�.^/I�Xf4�g F�����g61�������2��9��y�r4c)�n����W�:�ZgzU%��)�r�[�=�K����)����v�-�&y��#8Ӫ<�\�LpN[����qjǷ����p�,9���ѝX'2.�5m���!ލI�y�9?��ݞ�w��Rc�L�;}F�Y�S� �B>�>�k3�浥����[I��+}L��W�n���Uz,R��a�|*�>����*c���E�������->j�}~���bįXV�LtK�K�	��P��������t����8���WNr���z�[9ˍ�B��Q��"�W�n��m��,�>s�v����[�n�>�Le`��'P�Է��K�LVAQVeZ�}�a�Ϻ�zN�v{�Kq,T\�LʕE�r$pl'�zQ2�I�f�����]ˑ��M��B��vn臨f�X�����M����ϩW�N�)ʞ\���l�jߵ1���;ޫ
xa��"eM���$��Ж�	��ۻ@�<C�\��9<eB�O&S��+N{�K%\�F��\Iȧ��؞P f ����;��`d�=�E�A���t�C�אd'����x��R��	f�a(3(:E�|h���$��pY=��i�z���F�<gC��t��.`;�_w6�.����z���8�dW��a�)��\]�#�����%)<yWV��s�a���VIǅE��a�0�5Α&�#��B���o+�ɽ�p���+�����ͶGz�N��=�ɿ'N�o[��x)�13΄s%��r��4��˔w܆��U��y\��X*d���c��mx_�!�ߞ
p|�gr��)��8Ҥn.l�|@a�g�1�}kA����D}Iˤ���]�p9D�9G�ӎ:�3fd�s����J^�� K�C�|��f��g�L��S�tU��	��h���O�IeX՞�x�E�g2�]߾*�0���V;�|+r]�Fm�"�hlv."x;��)ǜ�[�~����+��t����[��d��X�m�x:�J��xOg��K�끣���}�k��y9-��C�϶�W�PW�E�q��m��֭ް��Hy�cC��%�����S��?FYٜ��K�#��_���߂.�n	NT��v��qZtѼ�ܖm��qⴎc܍��vwR9j
tʰ3��Gθ�Kt��r�O5-���H�W��ƫ(�j�]�4^4
���H�'nw&SVu�:y0׺+��J7��a��au�ll`A���t��t��y����:^=��%�+�
��q[�%�(%Zds�7��Zɋdcy�q�)N��Լ�-NSm�M)n���a{0ɬ|�q�52�t���LIK�t���뮺�7�^��)�yPH瘩��GO�<SMmt	Yn��s����-kq<��Ϲ�Z�Ҳ�!`-4!�:��J��p7������n�&
�=�8{O�/^�r֩u��2\�vK���`;��>f��kM@o万i�X�v;:�4�v�[��/M��5�J�[�X�!A�JB?,�W�x.+ё����y����#�
+����������8�\���?	u�V����o����p.�ݎ���J���e���ǢO���.��m��r�Br�B�A=��ˍS���(NNK�fA��͇��w5j�2�%��3�3u�4ޤy+���{}�v3��>-�җP�2��Z�Q(�w{.4��^�R�4��[B�x	�Y�i.�-q�uz�Mp�#���C~�\ ��e������o;3���3EMG��*���(N�p�-����i���Nd��fϴ4�����}޵b���Ί�i��O�h�d颏	ZD5����p�6��B�*��mmf��wRg�����Bra�C0⡝�m��WuXi�4�IVi(ҕ%�\t�4u��v_v�Up�C&�g�����3���:w����7#V�YA7x�}��	��v���6�73d�Z���aP����j�b<�ъ���3B]n>4�D\25�b��³zX�>��_����������B6�nJy�|��K��;'O�ܚ�l�;+����3;+m@_J�-�7�ig�k\�8|w�͸j��U�6��^N����q#[�?Li�V:���p>"Uǁ���Y�v�05m5-�wd:xf����������Ǒ{�r��;���_E���K�f�3�s0�T
�M��E�T~
&K�W��lo�p��֏����şR�B�t9 �+C,E�
P�8vI5C��v������Az�����yՉ��cZ;TdhtpT3*���T8�����j�ۍ���k���z�%�G�T��a���jW4ӂ��7�FҁhG�t�x��g��7�ǽ{Fຢ=u/�X9�᲋��k���#��蠠s1CH��)#�>�S��W�^7���VE�PL���WH��/Ҭ�����o���yN�C�ef���Y��wR(�Y6�C���@mu2�3/:�)�n����
[�w�1c�<0l� :��Y�����N�D�K�L��y���x�~f�3jP
��T=V,�N�K��G�gX�&����q	Zk���u��2�4�U�Ȑu�.�D��h4(�2[�w�sw\U1���sxj2�U��R��6�����,p�auIo��#y����¹�=�ؖN��Oͷ�e	B�W*(��X���B���)C�e��}�X�	�y���G
1A	Z�ֲpV~����p��%��!t��\]{v/w*�x��T�,����x�x��k�PS�rd��	�1��C�a°H���<3�H�������L�~�Y�yf7�m�0A�M��.���V�<#�N��w�^Q��)Epu9d�m�Yw�q Î��E�����u2���52W0E�AN�N���tی�Ry�Y����\Ԟ���3���.�ϕK(p����<3���8��X<��c��$i�GX�b��l�U��� �P�S/jr:~�8{)��S����~��o��/,���h)�l�F�)��gk��M���i��w�!�Uf�J���E�X]G\)�%�s{�Uu�5yko9��4VI�e�UL�F�K��c.�g#"�Ed�aX��ST:���
��v�R$�d�ϳ)�8A�4�E���+w3!�T���C�G\*�a�:�E��i=��B��j� P��MBe@C�9�y�Z�;4l�๥�i[��"O��yv4l�� V;�HW�ۥ�� ˮ=4Z�f㴬a�e�xh�u���V�(o3c3);���z�(�Ƨ�[�QM�BKU᧳m�r(�f��}�nvr��p���8�^��9;SL�}��f�Vͻ��L�c:�l���'P��~[�3cy
h7��k. c���/<�pD�W�V՗����r��D�}�P�Y�D��'���z�n"�p~��^�d���`�C�Qi.I�a-�`�\]'I��.l�.g����3f���^=đW��V���ÿ*�_�#6hR+�*�yK�B�#�<eB�O%b�{4���>�X����:�;� ��f�m��q�Q�(�tL4Mt�4G����v{��9���z2��Ip���[B��� �o$,�@��N��������S�e#��&�1�D<N��^ns~�v�=�.�3+#Y����� ��YS&%P��'Pg�����N(�{�����Z�Nw��C��P��Gd�]f�z��E<#����+j^|�`�r��չ��3+9E���?�"űۊ�Ֆ�>h��^Z//��qK��阳z]a��kvP�K�z�������	�����tN�6ٳ]+ie�G�Eq��ⶺK�p���P��ܔ�܊�u�l\�s��7�Q��;�ܒ�	�h#s=6�%��jx�-|b�һOxvx�V�V���]�m�'`w�x�V���O�]�>�{��}����[�B�g�u�b�w���I�1K�D�J>��R��
���$<wK+K��y�qn���F�Ԉ��uy~��t"P�=����ׄ��u�I^ �Q��ې�֥y� �k���Z�Up�ʘ�ۡ脁x��rS�M�{����XW�ڢp!���KϤ�u�U�Щ���kÉA�\o'f@}{\DT\�f�	�ҿ�Ip�-���^#�jyQ<~�Zy�N3��>c�c��@�l�kB��|a'6陎����b!"핣�o�*�]�2�]�Ab�˓�W+��O*_yLH�H�z\"§�E��D�t�/"�pL�����tA����2����Mo�:��T6g�p7������m���+N�	U ���S�cL8m��|���e#�"4]����+x����?UZb�����ҷ�%�����6��:�^�k���^��Z2WFF�0�ZG���׮����/vl�<߆n �T�t^	ךz�r�����֮(E�	�;?e�@�����6G,�r�z�|�)�T;�yX�=MԸu�T��e�~S�,ɕ1+��z^�����=�9&;�4b[�qޚ1��c#�B���"��\N׃P�n����&���`v�x+�Z&�Gט�;[�w{ERs�L�A1-�}ս��ùng^B���"V���T	�i˦3�FM�^�|h9V�E�<���t6m�~lܴ�F%�)�.����3��mF��\,J�}�x'WQq����\N�z܋�N�����X})$<�Ի�u�^�z��_�|�������W���DC�gW��q���궉�$�>�TD6��
�L���T܋��nM
����d�w7X�k"�z�R��j�i�8)�X7�tXC��!�b���k7���S�=,��S��\w�>�SFq�?d�Y�,rXAb��c"�ή�O����T~��]���]粆�ڽ�I�i�^���2��}��i��,n|׺ |U�m_����(#�8a�:u���z��k���G�m5�c�����m��">����r�ǷAJ�9h�G��/ӂiD{�x��^��U:EpL�+���Y`����Y�l�t�����Փu��1�^��wX��zK�չ:�唎=5q`�����R�b�2�W7ivSU������{˴U��4��_K�T�ȷ��n=
�Wh񵦡�m)��"���=ڵfLJ7� G��A���`�}�v��ƚ��n]�&@t*�����F�r���yJ�����AN��y�J�e�A'²�lM��>G�t�˫o,���Mz��is:VЪ^�U�1!�����M��0g엓.
�=�QQ���h鸛��!NFI����e���}�~6���R���'ܙ����\mm&,7�S#/���'�yi����{���/>��%���2�r)��e�#얽��a�r�xxZ�f�}G��6�97{�,P)H�V�
	�c�/)�E�VS�����W�p[<��م]����>�)����r�D�N�_ji@O&^Цfu:S�ۄi����w�M�WxRY:)1.P�gZ�|��w��g�:�� ���Q$y�A3��)C>�-AWܡ�6��ׅx=1P�%�ޥ��.�xE-x�Pޣ�eø'��l�$!��X���eF.>��<�b |"J9	'����O��k3��E�q�˷���Vtg҄;	�f�"k�3+�Y�����n��(�o����a߈�:٤�xvoL���EXf0s�(���t˪pH<$��hn��ai�[�L��@0�
Y��6���q�7���0E[�.,k�hW�q=z�F]v>��M��d&��/4��1�S��g�vq�1��l5��SזrŖT���7�����ny�I�}�����X�p=u�����Iऍ	���l�g���+0����c�6��)��A�㫗{)����h��|ٵR���^v2lˑU�(�;�WtsJ��Tðfׯ��Ì�Vk�����s������$Aŝ�J��xݻ!.]��d7�W!n��B鳪Q�C�����X�i�E-���Z,Y��0.���5�ނGGZ)cid 7\���]z�����;R��2�][�ѱq<�]�x�f��6.��t;v��uΌ�(���gj�����{���҃��m�f������2���k���R�qH��>�lKGQ�}f�v�.�o�Gʹ
���.��
�\w)���/)|E+t�[���|���s���:FOAe���zfV�SL�p(wwW��DEKL����$Aj�n3V��_3zo�>N`��R������yK�ˣ��� �p�ȳp�+��]�2�n��mt����`��%��noɺOo�ٷ�Rv���B���7f�F�c]J��:4�](SH[��wh���xb�����ޓR:��ޜȕu�LI[{�i���ѮJv񨴗����@��4n��6���XUM"-�P�з��݄�6�P���2>W��{�)|��w2�>e<�}8ً�WSꐂ��ׇ�3O�Ľ��`~�%�.m���G.���W{�0�8�n(�y�w�z��}.e���?�ъy�4�5�j��x�۷�v�;�+��7���'i�H�o[��Fzo)�L����nv�	��Mvuá26S��;!,a�orv�][�2n"����ŕ�UD�O��ᆉ��w`�2D�7J���2Q'�sUB][��Vn�����愶�u2���Ӭw���hv���ѼYS*�f˭�]I���u,:�vz�:�Z�1����S!��ȟ9���w��9H�enlGe��m��4Y�Yᎎp�[���ci���}/q|��[ 5���}Wd���Ԩجņ[���#r��4�����j�r�B�K�T�z֝J�&��(�.�jmJ�V�,n�2t^���K-�V��C��;h��.�bBy9w�f�.�:��~c�5��0W;}u�� �[����ֲ���cf�f	��԰r�)zJx2fE�_����"��0�WEv���!�X)*�TGh���;���v��R��9�)�Nwn��z���݄lS��$�}UG*F̙���ǫ곪�ިe^�f�eR��=�YG_{s��S)ks��Bj]�B�/���3^4cA�3o� �L�,����	�-bw���6���]�gv���f����Y��:i�޷��V�eqϮD�w�5zľ��wGG	��{�F��z�Vq��l�D:J�YF� ����)�.�w���
�ݝܭ7=�_}���y�~�Y��%���m�&8�Ƶ�iXb���F�X$X-��J4��(\��\l����F��m�ej\rQ�VW.`5��`�J��E--�iaS2�YS��J�*�m���F�US�+l*�Tư�[`�aZ���s2
)X���X���B�X��*�k+��µX�XRՕƪ�K�eDF+n`�"��V1r�lDhֵ��`�(,�V-�"TmR�QaQ�*c`��l�
V��+Ub,Q��J6�Ck[h��������m�\J���5�2ն����
8�LiFѕ"�Pb+E���-��*[U�X[D��-*����X�ն�**��h��+l�F�	(����+Yg;�s
�%w'����=�4�q�"w��C�ls1x��y�N��hD����R���s����󽃑n�踘�Ӎm��^�g�z���|w�o���C��ϼrjc����+�����ٸ�x �7k���6,ykW1�(fKS��ob3C�+񒗝aup�Dr��¬��O���uy!��{eC��w;����.�/��'�x����Um��4�g��u� ��ߜُ�z����(0s��.�q:�p��Rޯ"�{��a��U���M�/��/q.��pUq��LʔO_
���:�l��o�>R��梆l�ɢ.�ݧ�ǹ�߱��*	rQ���̥\^}r�+�[���(<��:�f��PL�i<$�W-o��ߧ�U�
��w��m�he�4�$�SE*���i��.j�A�*=4_����W��v�Ԋ�����۔�)�v�x� �52����;�z���'N�����k]����O�a��+����໊������N�8y�y�IzdNky�ҫ2�\�����Sv5`�o$,�:&�r�-�	�O
�YH����w��ް,�MRV�[{h����\�R��F���h$y[�]���Y{�ڲ���@]�㍃��|��U�p���f�O����˛P�66]^�v��"�u��r�uҀ�$�C�����Wv�Jv� Z��{b
l37nO�%�\��VS<f��C��UÜاn��C$d_��3��!􍹑G.��ۙ��Pt�s��`ܤ�ČĚ�)&Y�^�z;Ma��.�����e��I3�r^w�Ӷ���f `�ɋ���צ�$�u�}d�虍��k�P�S��)*��`��Ft��}�]�j���6�����&�Q>��U��K{·��,���nA��jz�48H��yG�[�%Dce�a��y~3Ӆ�_�D?m�Un�xJ��u��ᒒ�~Ќ��ե$��u�Z'�>�v`ۮ�cMs���{-��zm�ݿT:x��y-R�W����^�,֥O	;7ْ:d�R�k�،;]����L���)�����������=]�jo�����v
C�Ce��%c��\�<�UOiH��|a'>ۦc�V' Է���[w5�"d5�W\�>���4U��3�ƫ���qՊ^�0T�*��`��GR$��\� ����B��ͭ��跅o�hϽ�f��6|�:i�p*��j=R����F&ZUp�@E��J��S6p�eku�@��z,�����L�_"(�q��H_;����?��	pPth9ԸGy]\��G4u�����v,�LP�� J�i�s{0��9�x��8�Z�.�_`x�<���sf�J�kf'|S!䨳�R�U�Y�T�F��⡝��L������tJ�^�N�^Ja����Ƨ,)���G������?��<7��º�}���8�e�>8����f�f�ac'<c�͵u���FF��
�y��xJÈ�JV;u�\���Q��bv�r�o�Bu枭�!���*��L�ر��0j�kބ5�oN�u�y�\�Zd[�Ƚ�A��rtϹ'u���NKyN��@�������f��7����ixS�]໇��{�=�:���=����rp��K�Y��=��\}2�0P��I
�0��w�����K�\�7��<^M���Mr������n/bg�ʶ�p'�yCؕDCa�4%��O��]Ȃ���7����d��fsA������ۍY�Â���,����,�#�#�+w��,c���n���l\u���^g^9�ʕȱ���sQ���ugL'M�m�=�@����{�3��J�-{�k�_�P:=k����S:�@z-#�Ac^�i?Jֹ,�O�:+�����Û������0�_\�DBȶf�梧Gc|3!��e{6�5�G�g��[�S�{�q���^�Js��~�u��s�r�����KZ��盽�OM>����q��wX������n�֌�LL]��Z9p��o���qM��4z�k�2�#]>?Ki���yeA��*b��;�q��ɓ^`r�ȸ0zEU�Ƌ����1!�֯�t[Y�z��3�8K�#���Vo����m'r���s��Xvh^���ţX�I��`�Wq���["�6_uo��q��E�]�?H�48֓]B���'�d���r�ߛЛ}8W��1�ML��]X�r����Ţ4�ܖ3�M�0G�z�z�^��[��D��K1E=0�m��ԾhN(g�L�x�)��X�5��~��P/3ѽ_���|;*����]m��r)��(�c#얽��a�h�����Oއ�L��{f>�s~>ݭGR0x���,��v^}N��ynmo�E�';�}�Đ֑!e=��gvs'L�GC2C���T�>��6S/
fXηJM�G�=xw� ����"��3ŨG&�g*���<w|re;\@��j%b�5�B�����O���9�Y:E��^qwxv|��O�Pޣ�L�w>��Y�l�5��e'X�v�֍7�^��A�E�q�pi`ꝩy�3;,�ֺQ��qʓ9܁��Va�w�&.q@��6�ogo;)�W�Dkxg�?�]��'VQ�/��U �c���*zq����%��pd����T�`8V�]s>�tۖ.����q��Q�|(�q��n����W�zu�:L\WbUw�@��48_4���5^y���)�9����~��*C�GF�Q�����|d�7ґV�B*Ù�QkF,�<�g�|�x��Z�;w����}�9*¨�q^�/�8����Z:�qcy��\�
�&D��A~+�s�M~��2B	�CՑ�	�Z6}+P��U.&8'-���ނ�<�~��j�O_�I�H���S6�$X�-�^+yg{�L�Z���W���8i�;jE����xo��3wg�����=8#����6t�{#�zm�C�M��j���ۀY�<�oЇv�崇�N�y�{;�}n���X��T;�s��)p�o��p7�bW�+�&8�����w{������k����Lb� /���-E��+w3!��Rޯ;���uq��ӄ��ٙ�;'v���,�8�Ih�O̚�	9Ȗ��:1_�N�1�oW;ZZ��;{nt���Y��
�=>�Q>IĹQh�-��e���D���őr�"j��mAz���CI�Աޛq*����$!�\:��m��7��o+6�=���W�m|��:�Nri6�s����Y� �!���ؕ�n���"�N�*��"7��3�zFA�,�9q����Q������z�=�53E�Gp�Y�AاMR�MEI�th&�Zy�98�r�0��ӉrLv)�1��ɢX��U�����y��p�v�lk�E��I���� �fZG}�@���	sQ9��S�S��#�t�i�#�@8+�٭��Y�{kHs�e��z[�ɔ��������&f*܌5�X������9K��$;�Q�.[#�䅐��N��� ����<*��`ާa/o6>�	��]lY@  7O�ϫ��;�=�;�yPo�^�����ubWyn�c�c�,Μ׮ZNRau	o@�S�.�g��e�T��规v�Ãz]$�0���2�T�]��N�ضP�^ *�{���7]+m�x:���.����n�8]��(n�p:��p����(�ycԌ����m�L�c��*��޵�´�v�h�����XI��ո�}q�H�UC�u�Z��qV��4lyǈ�3ԥo��ݺ�m�x:Ҽ2>3��5v	�ܒ�I��J��M�+k��Y�v<Lm��]�-6�[K=6��ڇO�ñy���Z^0n�7s�!�G]e-V�=�;<z��]��-ی�RQܼ����X]I+W�� ��&Sl�YN��Y3�5at��ȭ���o��nPV޺{N���m����4ط�@*s��ˌr��6�X�l[�O��rTfX������ȷo�����2%�	u9x9�'�,:+�s)�<��m���{��l?��Fv�%�6�i��5���E�9"�NI�~���Y�Jү�vM_
�w�v�3��x=�;���R���d�u�|�z��_:���Z)qh�>��AE�=��������D�$�۴Qv�q'�+޶R� �����G��2����ee�B��A������w�PB%��]��կK��{h�P>���l�e��Ƙp:��^|jr����6���\CZe�:v�����f7�GZ���d��,�Y��	�';x\��W�����e���b��}�v��/dy/$�+�!a�a�C���R�tǨ��?-3P���/�
k��+a�~-�(�A�ټ�oT�|ߏq�$ݥ����eȡ{�B���
eƩ�N�E�Nof�����K�б^��I�ez-�a$VߩvN�PEY�=ʦ̩p��㏆q�Z;�j��W]��0�{�d���wCU����2�&
�ZHP�V��r�旆��5�}�����I��²�&TWu�~��fq�»6�"i>͙l��m�N�Jw�u��I&�����w!��eu-�r�-9���� �
�s���Y�+���l�؁b5��0[�3.������d�%����牲� �7p�D��֎3F�::�����ʧ�Zr\��{����y�xe[D�
z�;bU��
��v�{N1��Y̿���Z�Ĕ�Y�'$f^��~�J��v*J�iY�\�.�O�+4Y�GawQ=��vk5�zײv��3P�OSX/������w�tr�r/y��6��(��"ك���`��7��������s��^�*V(/a^�}qpuR�Oem���f���G��*/tGьx����N�E.|`ڽ��e�8�W���w6�+�0.#.<�������?E_����_$Ѻ\�`,��6�vyf���Z�0�/�R:)��¬���h�B�[7F{[�����rݨ�2��\,w3������;�FN�ye#��M\YX��)���>7{��<��=���׆�GDX�)C�B�Q/��*ddXz����|^VZ<N�����o�{�r[&�gWvu\��SC �A<�̟b�r�L&�59BԮh18��������^�����6��c}pߨv/j¿Aٕ�RDw�����YȦ����G�-B9I c6ʵ��� �ڑ��7��8��PoH6����,�̇k���(���W�������U���3� �+��y�z��N�L{�P�8۲YAF�syW[���]��	��}�p.�)`=u����Os.�E B��& @���Ѓ�ǉ�ѓ��������P��]�VR/��Ŵ3Qi�x�	幵�ȸ�ǽ�\��V��W��T��-��C�e�@x2#c�`>u2�L�M)`?[#Oq����ð�\��τ�����[�`6��F���qɔ�!�@��Q+��υ
e�Y,G�~ϛ��Ip����WS����fx�jZ��7���.�'��l�$-t������8��U����op��,�ܜ}%���
n��'V�,�2V�bj091�&�����Rƹ�^�.#d]��[�7=����rp����7�
JÕ�f0s�(���j <�'�~�2G��"�ۿR��o��������6s�C�=���m(XޗI>�Y��w���rgv�\�ҡ�j�p��܆�Y�h����yT��U�j��<�߻��<>��Ob8���r��zQ�x���J/j���lS�/jw��!�ޑpQ�W�8U�\��/����K�.���슩���!ƲP�Ӄ��8=6���u��w�(��7Jc���I]��:�����x��!H� �.��������<�i�fZ�X�f��Yx�VO8P{�7��(�Ӡ�����MZ�hP�.�07�.�����\���f|�h���7;(�Z���
��?'���3�[ɿ��c<���oq��ة&��wq��_b�H��8._���^�P���eCUL�F�p�lce�����"��$��3�;��Տ�;���RZϥ%�c�__
�Z����s2uM����5�x��h�h5��%�#U"���E��I`|I:<��״� y�Keg���B>�����3�9�o��-K�=�(#zo�T�EP���ɟ�خ�-�Ԫ-uF��`�<����C%�3�N`�X�"���� �����k�g�(�8�$�S@�\^^M�bLZ�-]N��z��=�m�.V����QXw��M�����u1�;���0h%�E#=��s����*Ӊ`!��ضY{9/K�Z=,��|�,�2�o¢��p�L@��X��*��ov�_m"LC�B�o+ɞ�T�5�K� �B�hr�-Ʌ��O&�.+�F\ǣ+j�k5��7��ga�v%�T#�Y�fŜ[�-[��Y�L���c��组�wk]��[[���p?f��l<��u35Α~X*WWT��^�GK���.�#��9z�>�.��;n���Vư$��x iR�MH@Kk�V���m	F��lѤ5�d�5|�k/^�/o:Z���{s��SY����/³�}�f�j}p�+��4���o{�GQzJ�wHQ���eˆ�Z)7�g�W���l�OV�||cd���Lۧ�R7N�+Uf铬�p��Ż��j�����hԍ�u�5��+nH6�f�,�&a!��"H��[V0����`�&s�&^�z#�©ߛ��G@7�|����k �u�&���Ae��0�R�IOK��벙���u!3~��70%D�˚�����Y�R�v1�	�.b2F���2F��a�B� �l��{Ecih�Z7�=ۡ.�7M��e����c��Bc_�r�Ie��\�tV\�/*�@ͥ�K�z��~���o-닶�ǣC	��Ɍ��I"}<�p5��V��Z��|<�����4J��(P��{�]��Z���C��Q��p(̓��4u!"���*$]��r�b�ĵ;�]��x~9d��D�ő��Â�c�1��p>�L@�Ի�zL��e��0Xl)i�_^]����|(W! vo$�.����d�f��'�c���$+#x���ێ�8��R�4�ٗW���JU&
���̧ئ�{I|\7���sp��ax^JG���+���z6ċQ�\���{�9�k���N�bH�U�#Cxf���T�����KUڮ�FŇ�B�X.��@�n�h5{r�+�2Vs�
�qt���F˕��Ү2���g^"o�%�rj9� ���y5���)��iGG��'y��ǋ��Ja�M�<˒��Ǚ�h��BP:��D�0=C�*,lc��6o	�/q>h�ь���
aOb�3}��?$/dH��O<<za��<<9��O���)6���d*�_wtL�,��b"xS�t{zcܲ�=&�=���n����;�ˑL��A����ڹ��zV#yO^��<PD]qM��V_��
��f���/�_d[= $����U��9Ǳ�}�Mw4����2�>3Y���ör�rۀ3�����k��ͅ0s!�=yW�\9k��X����!�������E��vx�E�Θ�='e����]��`G���Uw�r��3�n^�GN_e,�=��u]�W����;�\+E��>�-��D$�ݼ��qk
�-^g�5$���	������7���F��C}�^�Xs�>[�"6�(w��s2NJ�y^���{n\3E �&�6��r��D�*~�p����SAt6bޝM�:�W)fh�S��C�[�ޫ=�l���k@�Yߥ}�CF�j#�t�R>n�>��|����y1���3�3�zٜ����r�Ӕ��^��VEҙ��Am*�Ҙ�����������L�#��$�#��|ki[lTV"����Q-+JUVk.)h����ֶ)P�"���+Zekh+B��DQG�Աh�iZ[m�e���kEV�ڸ��D�X[B��6�-�F�c-���ґJх�
b�ҴYR�5���**K��Z5l�����31DS-���6�EQZ[Z�X��K-*���h�b�D��fe�QR�m�-�QUF�-��QDX��ŭ#m-�d�!m��TZ��Aq�AJQ-�mmX�mX��AEڊTJ�R�r��1��RR�-�UU��mZ�l\�J���a���j��J���R�KmJ�(�ڲ�����"�D�mn[�b5�m��V
��lZ�(ږ֖�E)S��r�Fإk*�+��6�EQ�Zҕ��ƥ�im�
e���*"�s
�Q-�0��ˉ�� e�UX[j%����[ab��-����(���dUA�Z���������[=�5KЫ��'J2ސ�]�8 ���N6l��T�3�%��;v�|qSɶ� �vؤ+��qL
v��EmI����%nb��'Q�U���3*�/$Ӯ���!Ex�^e(ŏ��{V��v�98�:�OkQ����V�A��!1J"�#����~�[��������;]��ݰ�$\{���ʾSr��qqO�GG�x����ߺY�8r�f����a�X��/�B_�W<�F��WF<��o�6�(�<e6��7�W�{`|�[c�m[-�&�gܽ�M޲8z��ò��2%�	u<�ӶHj� {vX�f.&�|G{�r]�#i�BĎN�G���l�@�� ��eW�ł�iV1�4/�H��q��6�*���D��L���5�k�{<^�9.��3��ଵ�8�j�z�R��LG��5F]k��wc}��Wh�2�ݷju��T{\w��o,�P�VZ���#�;�l��nAʹ�{:l���gu h��Υc�S3}��&X�cL=1k@�y�;�v~��y��$E���e��Ɛ�˞$�ɗY�.���C�.�͍��s��!����E�Z���o��h�|�?Wncŗ��0��!%0�����;/���A�k>�坫Bg�3�Eoq�=Ѕ�U�Ŭ��^�0MWP�gs'��SwH$�kp���r}t�C:X�N-#�A{�\V)�m�iz�W����u�J�R�h�#�f�<p���Í�DD��{���3픹x���$�tǫ�'^i��5�ז��*��,�7��Lai�2�T�2s��Z�����[��t�WT�k(&E�VA�Sb�ð�i��w��@aQi>��W({j���B�L�����k�"Һuq��TGg�~$�Q�@g�շީk3��i�+,�Y����ˁ�<%���5��S�2��͞Fѝc\AO�����a�:����5y�P����ʶ�Ϝ�
v�Q�	��O\�s���."2�kM�oVwb=6j����ݞkG:dfoL��j�i�n�L�00 G���oS��?M����z�7���Z9��{%�W�>�2p�zX�AB��c"�Σ�su�6�-Wy�9d��@`��1�
�εA~�S�ټ�Po6����z��;�0F����w���Jc�t ���xW�)��e�F�|�+\�zU\|C����"7S�z;P.�o_.�wY��۲7 {q�0zI��rV���ՃV�q`��	�&�nF�2�AyYid�k�y�v &Qt��7�pПZt�8�r�W\B@�7y*�	.Eu�r,-�fm=�yfG��d%t|{i���@����v��R$�d�{���6�,6Q=qnH-�g�Qp37{4����pA^��)�Ou@�q=l����.�P�K7-���aޔ�~��ug���4�D`�G�X;Cq�tޖ���JP�B�:�9��T-mg"_K�S#!꫌㇡I����b~ܣ;'�=����|{�J�je*���D�yъ,�	��jr�K�(��QE���,��3�G�ؼ���>]�ߖ*�� ]J#`�.,U�e��u�Pf�^��o�ݤY�R���I�d���D��.���׶��І�u0�	�Е�D¿R!d�F�ʭ[�c�u�=�1���q�o^�[�-@av�DH��z�(����̿��SQ��SY�?Q�K�G{��N��{to���Rf�����OL�9��x��!���R��p:��sk��3�C<°u�{���Xz̩�HK�������"��u�OY,�$�3G�鲶Q[���jl����v�E���>u
o�"���rz+gcE�7��6�~F3;o|z�u��e�B�Z<3�G���3y����o�"_���I�zN��A�wE����z\{�,���-I�]L��;����޶ar�+�6�3��6Ү�t��w�)XJv�wZ����N�j�	����UN�3z�.�{��ը]�/q6���eu4�&�W���b����e-��825�p��E�o3N-z��s.���K�r$Y��9c��uR�%��X��f��V������J��R8S�!!��;3�cg��qab6}�	���*�>LpT�Y�/�`�����IqM|/�2���?u�i�뻩��l?�e�{�GA��(wg��Z�a���Y���yˎ�Zz\d#<� ��q�γ��*pcb�֮b����:���죧t�.#���w���]�7G,���W7=Ce��P+ǁ,E���X����%��b�f��nx����rJ1)-�o�e?XFH�e���ߺ��Zf3�^AB� ��E���C�ù�����P��Źg}�3�ԤV*��O�GE[�����Y���>1%�ҟ�
���&�΢[+��ޤy�W!g�~qǝ�������#67����T�K�O�1��Eh���c���7�y�E����׫X:�n�+%��Qm�����Ӎw,�a�֨�4�6��0R�sٴ��Q���m�օ���]�l�m�����x�AҖ��U ~�8|$����}�J0�5t���+�w�劕'_wM�.Sel��qMZ�*;)NK�N'V���u]�n�L[y����K�"��"�������A��il��S�.�#�;d�ٝ�VWd�Ǎ.��"�R��Poq31ֲ4f������ܜf�,����3{xʋE����բY ��fǌ��5����n�n�6�װ*q'�R��>��I����W�o+���2������~N��ݣ�]{IN���_��ēj���^μ�`�oْ�Y�س�}E�}A��*d��u�^�'Q����V8瑥�Ibr��P��IWå"��\EmS4vע��e�>���I���s<ϞڪK�vv�Ϝ�G�q^���y�z�L�<�\stY
�!2{_E���ø��[��U�ܞ,ޗEX}0��B4M�)�o�]���^}��G@����3�h�h�:��Hy4r�y�A[�mw���b����qb*&�b�ܭ��Qp�3)�uf��F�`�qOYmD�3�z�
՘�ά6�ͻ
3n��41�z�V��o&�=�G�	e?b�w�7�w����0yq�`{Ե<]��R��x�2�{]�HNoȻ��s�[�ɨ���P��2P��]�E���ٲ3:�+�R倿�0=��|�x Щ.M?e<D��;��34��T��T���"zP1X�v����{s�lN� ����n����Zܮ%9̡�<s�����ΨZ7����#��o:V�݆nc�K �2h���Л\�����s��0mnu���
�����[�9�VGp$�o}O^�C� |��xg��WJ/�SWK֦
��^S�9j��JOI�4ȫ��~����,:��x5Q�q��o)j�-rJ��:�������w�8z��cr���2ұ�*�0�d��u�ڼ��	��\�G�-��������ez���kA�%�BHؽr�vu�i`���ݖL,d炎}r��^p�=�^��p��4�;{�����,َ�4�DPݩh�\Y��]����Qk~Lr������U�\���[�i��c+;n�eA��b��L�wH�J%uLƐ,��VA�Sb�í=��Lƶ+��#�cz��t��{�n�k����ϧ�o-\��jz.����ʣM�x.S��a�'��N�n�U��)��Īg�K��L�a�I

^07&;��Mn���&����	&�n߹g"��޺3��e[D��<����"d��C�pVcs+���sw���_h���ݞ�ދ~�L��邓ۍY��=K:]�f���Э訤XT�]�{h,�}��E��J��8�R�4��p��7���:�慂:t�n�(�툏�238��(J�{��P|��T�.q5,X��ћK��2�q��Ҹ��4��8�ת���;>���T���H��V�199���tۚS�Vo�Hk^�ֲ5�xe��˿K���]L�1�>��w��"�7�=���f���֞�_h�ϫ6��L|)�c�T�W��`�S63ۙ�޾��J�H�$��_'�u����\��"X=+Z�o��Y1�J�X�t?Ki��c��<i�1�^�=�K�M�vy����g�°�06���H�m�t����yƶm�wXhK�(~�����K�K*{}{)�.Q�<yiq,ܶfs0�:$ 1�������A[\�Z�}��O���C�z"Zl+�&Q��h�b0g
P�h(|�}.3ʙ�;���r�S����R�&�&{��j8b�^/V�x)P�w��W�F(��	�ڜ�jW4+3)�Ү��4^[z�w�͎ss8�VW|��F�+��*�����]m����M^�F!�=-NP�Үy�~�8����S���*]:f(iD����L G�z��	P͢a_�mB*^"�gu>]$��]m��[�݌����W5���ڄ�=��@֮Jk���f'.}ʼ�ckI�iVz�M�JW�ma˶��ٙ	��e�t��/�T,#{x�cq�e%�o�#����x���v�w��OQWV��Y����AFr���9Z�r�j�b��ڸ2t�+1���mm<R.ʄ������Wi�Z&�nBX�rxɠ��*���q�����d0���^�\����AY���"�ۊ�ܝ��:�ȼ��B�ʩqoY�"�6F�d��Ե�"���p�	�%��f�����{�W��" <ڝ�5-�6H}';��9���M�7b���܅��[8���O;ևx_��R�ZN��|�v��3x/(h����<���e���|d��JD���!�T9� �z=pL~��n=�ZтK'M�2��b��xl���o.�X��Uk>d��g���	��y�UL���΂�N�N���t��\]u�g�P��ǕK���+1�I�CU����?H�96s�k�����y�q���'9������p�O9�S�6l��6�8Y�U��D';��Ĭ�m��³Z-��pz�c��U����Ӆ���i k���_e��zE�	'S�ҥ�غ"�9�wMؤFɲ
�(��n[3�����^����;�Q6���<N�n��R7�����}U[i�T:���P��������}L�$�v��r�������b���pQ]>��}�oT� �q��]��],7��T�G�Wӻ�5�n]2BQ:(��C6��$��N],x�,Z�kNX�V���m�8�\��9�Ť֢�>��:��pB���5���p¦�J;���+������3�mHc7��>�o�ێ�U���(����U$�z?0���j������c���2��҇;h6e?-�͍��A�D�>�1ґZ9y!��cC0��{�w�./=�U��P�,�L�;��P�Xrq��	��Z�4�\��ءAV�_}���n���b�sﮝ������/������&;֚������ћ����!�J�V�o�%�{�s�#%�r�	,e��q۹��M�u����	�0��\��¢�v҃i�b2{��waj޷�O;[��?q}�(8�yP|=L������R��1�^���r��y���EؔD��g����z��H�JM+�du+3��lY��v��uz%��e{�b�N܍��oC�c��mxc�',¡�2�Uґ~X*WV*������i����<���e�0=wIXjX�LQ#��r�$�d�~�32��}N�3^��V�q�۹��ݎj��-M��>��fo�
�L&���F���I��O��X���WJ������љW�ɣ�b1〡M(��U>G�Ox{%pC�w����Q)P�tg�J��7��D=&E�o�Ot��KA8w�;!�9�{u�v����"q׾õ�Cϋ����{�FA�o,�*�6V;0�Z���X5�r��2�3�:D��k�3��xV�q�׷+qO|�\U���yǈᘞ��?m�J�+%�|��q��~.kSB���m�W���<j^7\6�-��#\���j�T��W#W\�=���H��L+6�Y�~'��2Z{��6��õ��$'5�� �T��ސ��j{�������]�@�ʳe����C,���>��&	�Ǉ�I�9�l�{��g]B�ܼ�O%�Jw%�^"6�̹0:)"���D����R�P0�qYm������=H���Y*��~�M�q���9q�Q3��"���Gk}˹��������&�41�%pE˅2q
p��&d��u�ڼ��L�z/v���\���{���a����G5`\����W�3}�	��s�G.V�����Y�:2�׻Ǹ�ܴt�(���(���A.�Rt��:�OW�`��Uʮ��^�ܽ�]��L_2�c:�v�
�LK��c����W���S�晴$���$ I?� IO�@�$���$��IO�H@��	!I��$���$ I?���$��B��@�$��$ I,	!I�$ I?�	!I�@�$����$�$�	'�H@�bB��B���(+$�k$L�N�M��
B,�������
�{� T�
+3NX���l!����*PUP%#v�v%:���h(;�P&v� H(;�)�)��U��4n��L��T��ӫF֔���gYI%+Ke"M�sj:i&��f��Y:�f��%M�R�6�.��٩[e ���m�6k\[��hj���    S�Ԥ�A�14�&L@ �~�R�(�� �10L 	�4�ɓF�� �0F`"��	J���      �&MLL`��I��CS<)�0���6�4�S�)�����\��I$�G�4J?l!$�z�IA&@ '�@�p��$��IrF�����?�4�ͤ��bI����  I*\"��I$�M!��k�_������ղHI$@�vU�?E�cI_�Y�h9aAE��oǣ�ZD8���5&���x�&�ۮ��� �+,S�2�pZ�K�6�� +�4�)�z��Ѽ[�6�s5��4t�EB�	laJ�0���VL�Ք��."�)��p��̆m�d���T�EU�6�`�0y�U[��a�6��M�b�(_��T���u�Ĉe�lA��Ncd�h!�:�Ɂ�0Z6�&l�ɍ�F�ӄՌ��o�sq^�&� 3�p�޻ɦ6�j&����X>���M[�V��ݜ�j۔��N�[
!ViB��A�-?��i�P��j�/a��ʭ������	���ѕu�	��J��X���R�[��I]L���k\D]da�l��J�z9*�F�ʳ���-�8�* 0��x�m���{�|�JxԶ�*��X;�T�vܬ+�J�:��q�`ʔl��`�+f���x����>���f�7�6��̕5��9�Bϣ�k��ߒ׊�F�Ѭlف�x�Wj{Y���H^2���)����Ś�c�;�Q��F,Gp|��GMm52E{�V��wǍ�/�tK���7G��BD�.P5����-��K������g$��U֕��G�G��V�kM�'KH�+i+Gi�y&m��o"fJ�:�#SA�eYt�|��BC8�1M� �ͱI�)��Ud�Kf�ܔ٩Ln�r��1l�]���_�ZYq�h�P��Jx4Q
��4�S'��5�L�X�ݖ>�J���b�+d�*;���i)
n�f omA��)\3�E�W�a�^0*(�T4����c���j��,d)�(�T�Z���H݄���3�qӱ�a��M�D�ܨ��]���!Ō9�˂�f��U�rV���b	=�7I�kmi��:���n�Xk�cV�1�����?��6�n�BD�C��qTz�<��y�fʫ��[���&�k躑�dጬ\QMb��G�!�o��K0�9ܟwh�uM���9�b{���Z���6����^���4�y�n�j0�gm�:�ot���
�=W�JUw��e�Q<ٷջϚ���rt'(�˗�F�]i�i��VZ��֓U�č8�0�l}&UTJ`�\U�Z��3�l��R�Y�,Ep4�d=K2�0���$}�:�����ݎd�ρF�Kc�m��+�fo*wOc!��o��/�$��(�`�s�e	�읬`�x9�n���q*��ZaX��XО�$(��l{!��|<��ʼ̑�VBl�b��%�*�D��UDq:�݋��v��/.�SI�s.:R��teu;|��\|�լ�&�s��Qҷ��ً���zH$V�U;���f��5C�셭�1<���dY�k�W o�� ��N��n[���ӓ��.]�.Ӈ����uN���#� 7,�Imr���4m�Vв�hI��� 
,��28m�'���H�`;��        �4 #B�w%}�\�;�kr�s{)��T���2�=����M��˺�m��߽l��`lYck�Ԗ���X�X��,�.)x���^p��G�.P�[9���դ��/��v�+VN�4��M�z����]W6�[�WRTm���t�39k3p@qa���vo�S�c/��4ɣ|++�.��+v���ڕ�W[��G���.�j�d��e�0�]����3uWb�4v #� �#f���C�:���]Y�-e#��C��R}��>���]�
Ժ�.�s�o��Ǫ�bv4��qm��= �nl�5���@:T�×1î�R�{�RBN-�2����7�zs�7̫Ŋ�Ps^ۇg1���E8��������z��C���u�����H���� @儁듇�:,I$�cg�����G���?��`"]����(�l�e��
&�D>V�(�
�	׍��:-Ȓ�(u�e��T���[�����ٖH����jR�i�8�a�0g]�ku�
,���:9���2CR\�o&�Ԣ���1YW����'z>'f)j������(��)�k�;���a��b��w�]E�uu7A9�O@g-�ֵ��@7� �E[����l<��Ś ٴ��W)�������)vIrN��������^�s���7lVf*+R�C!�t�:��|0.Cg#-�×O"�\�yJӻ�!�l�=9�ҘAηB���5fV�<��o��:�DY{rV�p@���5�����1�Ų�l�*�Cb��Լ�v�-���O����G��*�pW!�x�k,4���h�u��,�P�q����b�8^V%S��)����'Wiׯid��guY��,+71�un���ju�j�A�
�f�]涪ݱ�6���V7��uЩ�QfS57���7��3S.Y��!s;.�d�����v��0e��t��nu�fJ.�%LJR
�iW���<kZ'K�V[�0qzm:�A�˔-�t�*��SM;��Ea�.��J�2��C�Me�كIBH�sۖ�Y�V�����g�wee��4��ϙ�D��Fq3�]��z��b�����R쇦;��@��A�	[Y�����q� �V�ݭR����(lG{����>/��+_��FU�0d���uf��0���I-��:(	��Y�D�.�^t�I��SZ�^s.���JWb�϶��gA�+Y�㔔]Of
X	0��2�ͼ�
�]o�^r������dPܲ�11���J�8��m [+�1	�;����0��!Q��� ��g,P٣О�}���jW^	�		$�+"�P1��^,��v�gx���)�TPы�K�]l�	��ƅ��J��4��$���Y��ot���`�سkX`w��ad�l��������S[��m��\�eZ|jv����yV\�QHt��z�qTa#�*�U�%%%U�,��&P��e*�E���D--�T#MZԫ�}Z+G�[J�����/��J>�ª����ʱA��ǧܔ�����O�2�S�V��{���߻�o���FH��/hKt���~����d!�6y���آ�ѯ�/�=t~a������+�e4f�3^V�M�n[�#���;v<�*���W�mD}�ʍ=�Gx��`ST�Z��+(]�w�q^S�Q`��R��e?\WW�a������'n���%C���vWxvĖ�떮n6˫u�W�$I����/��x�])E;���	({
�v�ڍ&npR������7�������&Je���=\5K��Mt��R3(��ԏ���wp�t�g{�����Cݗ��m�f�f3E�u�Xe'l�ц�<�.M$�b���=^�n�0+��w��Wi) ��;CS���*��i�Nn�2Wz�&Ra�oTa�^�^:�s֨�w�jΌ�ϳNt�r
������5ֳx/hSBv��38�w|��a۶(,���Ĵ��q;a�;yM�3�[�1�&s�㴛H�M:B���f�Hdb�hN2�z��I�
H-�t�Kx�6��S/��2�9������W��Q��x]Z��c77d���ؼ����%�L��a�S��q:fS}�I�[�Q��nɄ�
���k��Ŝt�hS
��^�^���I����CQ�r�d�T5���;t�Y��t�C��N�gul�(�gL���5Ξc0_9�;3c�vh��-�� �2;xßsη�Y���ZR=���L�me6���}�ɽ�S)�x�$�Xwp0��m�Jx�;�;̖�֪ӭ�k�6�iRN��櫮gi ��5�CL��u�ww�3iJ�f���:�U�B�UJ�ԇ���+ܫ��~��5s���*)�ٯ���������V�w&Zm���Q�t,�t[
ʫ{��l"��UַP�Ѵ�5�,KgN��KL�G|��,����]h4��UoL�l�:���HRq�L%��1���)��F���Ni��u�Z��VpʿV�m���ˌ宫F��k���oX�bܱi��ʆF���fSL�&)���.*e�ZN� �gh�Y�
t�3�������$����c����i�v͹IĽ�r�a���K���)&R,�N�70z'���0�y��쮻�gʹ��a���e��=/�!�����u㭆�YI��sM��{5E�7��8YV�U�x�lT]ԙ�� +�Uְ�;�z�m�]���(���%:����y��=�}M_��g���i�̢z�kF�j��-����Z�*��q�ݽL{�1�l��������5��p'D���;���hw����1��<\��Ž0�Q��Q�j�D�-�����q�bi��)��j�Sj�!H��(��&L&\ �-
dQKm����E�%$꣍L��~\���w�g;�]v^Ͳ��2˫�l��[M$��0�z�)x���4�����^gul�63(w���i4����a0��X�,�
N�S|�sB�R[:|b��P�OL��\�k����Rd�v�EV
b��*�����3��gO��a+�{�})ؔ��>�)�
�>��x3X�2��!�yp�+�e%���^����[��δ��Zi%�L-����ln���[)���c����m9fQ}��AMb����e��i��tv�L�e ��������8^����RKޞ��_N��_�<���Ʉɬ�]3��He��5GEsx28f��/u)��gn���i�Q-1mI�T��������h���I|��r��Iʢ�CY�|�S	�r�)�vǪ9�':��)1u6��]㬜@(�4Q�p� ����-���W��ί@��M4�7������FAquMѕO.��6"�8���t/�+(����P{ff1��"�y��Dzt���YF�2�n���5�7�7g�7���l�>y���W�6��z?5��io�N����Vv�Y5� �^)�3g��V�B�e��=2�*��U�Vڦ�7�*���E�N�}<o6j��� ��>���v�<<�Ӣ~"���^�Mj�����CW����b���.`ܸ�t>�)���w�^��x��D<��Q�W5���cr-�~߰P�8�?Ғ>7.'k�XN	E��U^�	U�g���߽=�jG`���,��9�A���˜���3��T�Ӫ���W/+��f��]7|��w>�'m��|�N��o�va\Ϻ����d�:*�f���Â�I�ݖ���߫�����k��L�����`�6 }�֗�-�Lm���ד�wl!�t6,2iC��2�]�icMq� �ƽ!�..�?}_U'��_n�^
�����j���d�ժj_����dM��oi%D��T�"0�2u��-�P����]����;7�����j*��r�܊ ��R���0S��&,$�����hq�I�'^]+I
�R�m��6����8��]m�_�uo�6Ya�\
2�y��8;��c����<�2�ߥ��Ѱo�z(I�]K����6���U�j�N���\1k�b�N�oN�!%rv��-a�w�.�+�����ň����.'.�-ެ���ց�:z��w���;�1��B�`��*���):o%a��U(Q��JRQUM�,i��Њ�ʊL4ش�����B��BRUST�U#R��\QLl��Z�-�V�e#MH�Fs������]����y��8뾐{������;��Į�&:uX��W{�z5�i a����B�RB�P�O	$��VI	&Ё��$6��u׋�d-$4��I!
@%!!�����M����O	aa����Il��(<2m��B��HW\�!	��I'i�$9�I
C諭�}�E��_�M�z:�2�ޫ�5�u�@��&XXI�������z�	�2�a&�Ⱥ a��x��9Ф ;a&Y-�f��#�Y��g�g��"ߜ�K,�X�3���j��3q]��V�"���������a�i�{v�,�ٽ��}�ܿtqxS�|����H��;(�q�����;C���4<�_�R�?9o��T�9��+U�ϼ�W{��G/���7=;1$���}U��;�D��r�<��$x5�M�M�B��v��}�U�n�/��;+�����!>Ka�	�<]�w�3Ϛ�}ݻ����NhL�C�7C|���_����Y�ԡͦ�>Խ/�ϸ"��v&��Hmcv�A �A���[�=��A_���;�~m����������m
��b��g�'�Mu��9�-ʰD��u�J�e7S֖I�{����"�a9A=���ރ��[�����ݻ�[�f[x��I���ci�$]�FP�Z��u�Ε~j��Uԟ�//�՘b2��P��`0֔<��Q�]'��7��{_w�꧝�o���Ոp�,<נJ���2'k{ˇZ<ǋ��=���):��l����Δr�Jz��2w[~~�q����}��g� 7�gHe�2���o�s2�=�g���I��z�5��X-%Hu�fR�K
��7���s����d+��U�f�LI6�x�ݶ�<5���ǟ���
<ow'��/��F{��۾�l lOm�ʿ*Xj�'��������矨!Oc
^,��+i;�@�:�f�7���c���ei��v����4-��}ב�D�B7Z��b��Nܽz[d�W5�,V�9Xq�*`T[۞u�l�^�˳��CQٜ�鯰�1ĜH]�|�-FCt�s8�����+�d+����A�Y����0p�w�M:u,�ӂ2��ihF�j5:�)�՝� 	{��ҵQ�]�tZZV�F�2�J�5���Z-�U
�l0�F���՗uUIL)S5BYIUU�*�YJ�@���Đ "��H�u���8���}TI��p^h�xc�����/�+��U��^*�x�R�ρ�5t}�}���e/x�Z�nLt':7l���C�ŹՉ��uME��S26(��O<k,I�Jϱ^i�m�7!�v����稳�j����v|L������W��`���
ܱ�mx���d���y-���w����.�jm)�Y�le y�U)�o��u�6�קk/��鈋��7�o̟m�����J������{/]�+���z��Ø6U�Ly�r��D]�A�����s���K��b��K�]fp�%d��fj�uY:�qSئ��=(�P���M.�L�(S~�>���.u0n��d�kS����x�e�v�?r(w�p>�=����UU,S/����`թ�[���X��~']�D��h��&+���3��M�R�A;��v!vh'�L�=o��C��mK{��Ț.1.V����e��� ��O�j�e�����N�ѵ0�d�㔢��W�=R���VhQ5�f��7�5����MhSu+���m�~��j-y�9��,�NW��INn�4��.�j� �{^Q��nȜ�(�����l���vM.��a�������Z>쌬����y"u�]y�\9��^��5V{{��W�)�����3�{5��������c�׫��7N���@`F�x�Ş��_yۄ���_{8Һ{�G�� G��Mp����Um/Q\�<[���/i�/MF�!"�%��g�b��l���֪�o����;^񮍚�����w��@c�*�OQ�����/��)�m��e��{�DʾŃ�3|͚���_qO��G1�)a��ݝY�&#<Ƨ�s'
�p 5	n���m���
�GjڝCv�|L��Σ)��j��u���&�Ӯ�䯓��F� �����a�QN��t�
��2ɤ*4�ğ��@Q�	� ���$�Q�_^��]��}�窱��wX��^�=�A��yږܧ���Vsj,W����*�����@�����y�{��R�e�=�;^!�0��ͳ�]�Μ?���1�"J�Pܯ%�W�CW,�E��Y��AQ���l�\�Y��=�S�<c�F�ˮ�w=�G��	;2�6�N��Ν?}U�����x�e9�'��ñP�{m ��1���o��L������q�<Ϗ����D}jV<�]�V�M�8>����_"���f�pg����(�e\��"k=�/��."�b���J$Zϐ>Z����S����)�����M��y�@a�޷�;���}��o����T��W�j��d�U�k	��D1vL�Ͻ��_+�d��O���L��:?x�͘����c#*C|��s������K.~S|�Ͽ_��?h-^cc�V����̊�"�Taf^B�2��*��g��}��o�a�jܜWnW���s&��Zc?�rjW߽��Z�~����{��y��6�wӝ�6��H���{wާ�3@A}��dJWD�n�La����{�7J-�b}y����l��F��̏��UL��Ԕ��$�̤�o��1[	��Ox�XY�|&NiQjͼ�$����~���89��}=e�G��_ �w�"��pJ��h�`A�̈́��ǞZ �y#��Zk�6^�y�p���1y�!�7s���{���u�?=e՟�����`
����Rs`{1�wR6���JQ�D��Wn�_�~��;�5~��*�X;�QR���h(uAq� ������W*�o�P\�,ZLTM㊲��;�/\��F
�ɬicRT*��$2I���T~B��y/�Ui�,�����Βkk[�ĠF�T�"�b�f	�+gt%�fR��M�:���??�]l��W�k�07c\e�\m�T'�0�L\`_}�Rn���&��\�N���]r�*H�VUHiUcMWf0�+�,�g��e)X���uDc�Lf�?��k]��o�d�g'͛7��u����~��z4w=�(E�e)�('�r�/1��/ɗ��u����]�FCT��ͯ^��~[7;�ǹ{����p~��������_�%���;��i
/���g�F��A|k݌�>0I��%�ȭн��]f\1���t�|����Vl���]g�ʜ��.��~k^�J:�3�@��v۰��9���ϱ*��zG^
w���=�lt��;9V���Ԑ>γϻ����h
�|�B��!�xQ|�ȴ!�Z��U� Q�0��߭.R�~�֣轳B9/+�y]�����;�Sz>��l�?P��iU�u���$�������ǭ�T�r:'���qʤEEE�g���_2��5�@ x2��~$��oR�O�*3���ͳM���a�{��T���Ŵo���D]��u�ϕd��Ӵ���j�E��Hg����,��V߾ծꅋs�I��}}%,j ��]��,�'w��k>�K��4X+�GG��ȱ�4�/�繓4a�5��1�j�C����d��)/ˬ������r��Q��w�ǳ{�W�T_1�*��v��6�F����~蛔��y�4�9M�vϲ߯׎%�<F�h� ��l|0�� �>r��!�����˴�ъ�o�.�[w'�h�ήv��Y*�=��s$��W�A���R]���06y��X�$X瞆:Q=F�Wia
�7��o3w�z��B=���?���^%�����d���v�#ko�����v�^*de�	/�T������PTy�ԥ2��9��	k���t��h��|��/�mA:�{�k�=���ʵ�Ni}xw<�*�Y}�s.ZN��^;TW�8,b).�:�o+S)F����}!e�ge�3�G��+���R�9��c��SR�ƥ�c�[f)���sa�0��ɍƉ���v�.��%{�o�VE����=�z�A2��tj�Ɖ� |�S"�GU�Q��t�B�R)���m����j4�K���H��7F�|h|iQ��@��%3���󛫧O�_W�7?1�ݻ�� �{|����@;`�����!�y�
���;�?�IZ���V�,˶;�%?wc��%��
�KT�`ST��U���̿��PB�n�L߯�[�b�ت�n���	5�{����h7dՀ�a��z��[���8�Ϭ��;3�^�����b1u����^����窱�~D���N�h�����HJ.w����P��)�U���ZUy䒻i���{���Jg]ۓ��^�7�_l������r���ss3�%�7�(��uq��ζ�ϊZ���-��^Ā�-���f�BI�]~;��W���Z&�*��i�ӳO�wﾯ�~�B�uy�5�+���Y�Ⱦ������[c4;2p�V�^�@9�o5C�	���i�_*�3�x<�*b?>)���˻�ﾭݯ��6�-eT(���Ƕ�Ȉ�_��\���7�ŭ�g�+ϻ��U,"-����,Zo�ݐ,N��E����H��O������R/��n��ߧ�(���3m��.Χ6�o�7W�1�a=��k(,�=�~�-q�*�g�W2_y5�Mݧ ��f	ֽ��[�u�6U�֛p�_Z��@���M�<L�r�j7�0jP���p��n�JT{���e���נ�������+3t�Wc��l&�7EE@�Xl�=֎Xu�9�.ެ�U�3(on:׺��p��1�y�Ve�"=��,^o��aqH�1ƹ�&��Ѥ�V��y�(i�*�2�^�K��{Pkc�iZ�"����0�
���-��fAi�ub�Ƙ���wed��p�xKj����h3Z
9x��Xk��Pe-���O���>�%����;SR��uyK+��4i���M|�����7Q?M$�]�g�����ˀ�O�H]�#�s76�P��vz������~����z�����l �=Զc#̷g+|��24"�E�Ӗ>l��?�R+BE������"��Z�wm*ZU%���#n.WWhU�n*Rᩊ�v�2�a�� R$�"�(
l�A'�D�E @f�~�?4��w(����O�c:wVl~ϕX�ֱ���*�����[�i9�f��(f7ÒW	Y�:;�.ӊ�������S/8g��}��c<i��)@c��֐Z,�`=g������x�8����S@	���e]����'@����#o�e�P�ħ;�������<�?���⏒4���@m$C���݈� CwaOQ��S��/ֶZL��ʂ.�۝�F�l��W�'ӏiqt|P����7W�&e�x��ֵ�����azyvo|�Sy�؀+(�c���)]�~���P�]O���.� Mhb"�t27��T˭�^�G�࠭9��s�q��&W`y����2���`��!"���^8�V��-o����{�?nq�����Xf�z�~�/��T>^Yk]q홛�%�A-��,��d�Cٗ�S�3����
@/N�L�I�΋w��Ώgv�~߼/ء��
Ƣ<�"s}~Q��뷈��c�Þ�E��c��X(=�s���{��nIїN�����Ȟ���3J̪�M���:'&>TԶ~�g%idu�W�v���0�����Z��14�:�gbh�F=;�L�<�Z�7q��\]:���{�BbZO]�Î*�g�ٺS|.�� m:,Sd�㽷��p����+�9�l6��7ú�*t���'r��/n�áIz�3ŉ@m��=nO:���wD���24}k�W`6NO'.�N�?]�u��N��U�!��Y�׳_��-�{D;�2��jOn�	�)��YO�ٓ9�(ۢ�)Y�eۢl�9K��3d�7%��U�)ӏQ�Y�ܷ~]��$���d��C,��%JΛ0�DVD������A͹4غ��h����(�.��AeP�`ŵ�0;��3tצU��z�!�������Wo[���R�u�{7X�����
(��G�QH�D|�d�:D��5D����h� ��
I|t�)BB)�A�����?'�s7���ԓ.MA<��J{x����� {B��dK�12e����nZq�v 0���h�o�v��k^͋c�����q	_�j�}���>�`�$f�Vb�j珨2k��djW.~׷�ϝ�dl��ْ�K2�Gx|�[.�Ư�)ӳO�rx����C�\��;�e���/�*y��{mq�cо$�(ٜ��+�!�$"뉻J�:Ozt5�����k��wlC�H��1��K=Ap;��n����1�B���G':�߉�O��P�S�'�4��Rd�X6
���t�j�R��������r(�|0"�hmߖr�̓���W
�ǀ��QV<)E�{�mjt��XF��e{}�yW�Y�>�����-^��,�s��D��ջ�^$�/�+zy1��9��~����sK|\��>}�l`���yg�AY���ly?�dr�1���=���q���{\�=V7�z�aO{���0]��=�r }��p�J���+ݮ.n�Cؖx�H�}�+�n��TtM\�_[&Jma�nn��t^T�~���B�qY��K�g
���˂<n�@�cw����VuJ/�;�\�'�p��ZV�Fl���m��w�I%YA
�UR��9���L{=
z1��c:�`����TKI���[�g�E��q��F��0N(�)s촢.�󛦟&��|!˰"g^"vR.��
�Cc���<-b�(q�+q�ˏF��5s����i���ٯPJ�|���WX�߫�?���űP,����ΏAR��us{��LW3�P0kI��u��m��mrm����
iYr�F���ԟ�O)#B��[ r�1g�8x�ѓVvS�;6BUi����]�S�+��X7	���b��-]��7��h���ں�{{�G^��8���y��k`ͭa��wQ��4�w�i�4$�� ��ϐ�y��+�:V�����VuZ��KKn�mm_u-�S)��*�(�������IuP-"�%+i���NR��F��5���Ӱ<�wu�I��gi#���莍�p��r*.���Te��m�\�7Bm�~S�����~w�FGj�Z���1���j��{ܗC�d�g$��]���I�_��ዕ����y5LP��[�����U'��	
�vew�Yo�J���t����e��te�a���m�/�\���c�۫ݪ�`�[/���;q3F�x���Ny_W��Z-[��c֨6_\�EKK��t��wj�jVNѼ�ҽg0fyъƭ� <�g����ϗЮl!��`g��X��a�$�9W�1\��ș"��rz�;��������rf��\gos/<�cB��"�6zի��tk�n�9{���:�����t����F'6V�?u��*���tV^z��������N�Pr�=ˡ��:2�as�y�N��n��
	cْe���Γ��n�,\���oPT |[EY���;M��^��iqt�V�� ����o}��t���m�k-�'��٩��_�{5��F�*�`t�������z}P��Z|������fI;�W^��.L��-m�c�/�m�Xz�&��6#n�M�༭ݑ����\<
�I�s����$��K���=��`w��T� ��ɉ2'��w'�Rdf��m�_0���&�xO�X}��㘘{8b��Q:|���$���o`���@�:I9�uc�m��~15��ըv�Q�ac����pR���w�Z1A��I���4�����{;���{�?��T��)�TU[�P��Img�I	$�o�%N�!$��'ꋠ��݅�AO�����0Y���q��O��a!$�����w���x�&D��?�=(�I��/���>���|��x��x��_<v�Y�g?F�d0�.M�~�7�yp,�^A����ff��I	$��N�ï/o�~A
�$�O�: I$��Z�,*K?a��\8z�=a�3'���}޿����O���x��G��$��N~�}��Xoz
��$����=��4\�?���&dy'�V� ��,*��׫�'��������!��#H��T$$�<��fz�zr}�7a�HI$�j����
���Qegʻ`U��y6Q�yv���I	$�SD�B��|I�g��)�\>�4Y��<�r���ē�|L�����(���K~��y{��I	$��T|�>�yk���g���2]~/�-N���'���||�Ot?I:!����<z������g����		$��{��ϯ�E��<{��C�?����Ȁ ���󄄒O����H��_�O�ARz�v~��:8fBzL���z.I$��<�ǰ.X������H  �Lԙ6 ��4::"g4�TO�ԁ֣%ɭQ�,aU�f�����d��I�a��?��\=���I���H`B>����I�����ǟ����!���}Y	��y���?������|�?t>���z����9���BBI'����d"��'���󄄒Ol�q�ϼ�ԟ�ק��N�N�@K�=ɜ��#b}s�F"K~��|�>����!־�:C���W��S��ϖ=�0��I�<˘�������۬�8�-�OGA�!����wY���̆	(>�d��$�I�"I���ϧ� >��?w�߯�� I$��>��OH�A�o����GARpI��O�c$�I>�'�
 ��&����"�(H!1R 