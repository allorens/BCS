BZh91AY&SY#�S�ߔpy����߰����  a9���  P>�     U �SR��Ҙ ����;�  ��EJ���gH�(�Q@*DM  ��(!"����@"6 @�(  P��*�  �Bǭ� ���ӪI�07k�;�A����Sw���}���v�S��ez���7x���ϟlv}+�.���"�O�����}�x;`���}���מ�EV�݀�;�ǧ�ϧ� z ���|ø  .|uEn�(w=�W֊}�;l�j���"�g͇W�{�_5s_y�{���*Z���4�� ��po=[j{o}����������}a�>����}�f =�v]�@����� ��|{� ��I6�݃������`N�] h��i����t> 3N��>��9�`rw�OGݎ���E4^�9��;�J>  ��=� ��E
5��F��h�}��;@�F�m�
/�s������
(:�G��x7/aO����OG�� |,;� ���}( 5�O���<{ت7��wn��@�4�  Aܠ������ֺ�ފ�d1��$�3�]�<�                       �~�7�R�SL& ��  C	�A����Q�00� �L���JS�P�      i�P$�Q=& #����` &����C"1&�O���O$z@2jl�� �5)J �d4�1h��4���>.E�Ym��6~C�'Ԝ'�}��z(��v0����@@7T�����U >�q6�������?�\š��o����(P�)^T@�v����5��U����*zS�c|]����[X�Ԫ���}����~�������/��=�=kKV���+����x/㩔u,�I�i�ؗ�Q34q+_J$�0Z� �|'	��g�1X&y�d4O��L��3�}�eQ�:$�%�g(�	���,��϶I/�vY�6���u.�퐽���w ��ԉ�F�J��9��"cd���m��F��D�5(L�Cq��s�Q>w��"pGMW7�tE�V+"Q�`�D��jR"'7��b:ԫ �"QOe"v��ǒ��W��el����H����,��DM��u�&��W��J-�&DG���??%��"<��rW�ݩZ�JD�H��\,�DH�R&���~��rV�#�G艦�"=�Cϧ��R�-ԤN?DE�Xlo��~{)/�o7+bk������5l���R�-�Nc+���0��e|���Yo�tF�"c�XX�����H��R'�"ܬ67�_?=��}�[O%"j�������|�Raoe"s],���,{>r'i�d��nI��"JH%�)0�A���;+Fd���t��9%�h�b����K���K/��%�SeȍMȕC���'M�����Cd�	P~{U���}�����eg�M	�%%�X�f�\/Q̕��_e�ę5D䃨�w���N�ӒljU�Î�&���T�9��]R`�Iӌ��M��S�$F�M����/�Ud:q�rA�0Ԯ��D~N��s$����`��d͙�3R��îC��5j�!�Ml�ꇵC�C��Z	X	V	]
�:�LWZO�,�)q��[Ա�K�*A�Iu����}�grYܕ�J�ƒ����I���7ԕw%o�ZN�'��;G0���P(@ט������kK���Z·�β�_4�ӝ�!Vld�m$I�Hg�#�񢖄;�J��$ޔ��LE�J"�$(�;�F��H!�n���)�'�D�E�'~Βo�I�:��"=�6l�rD۲r��r͸Na���`��U�h���*$H��N�bN�
�<&�^��0���/
7ߎ|o�!�F��'bg?=�Ϻw��ri4���oP��W�p���:����Y��.�u ��ԜN��Z10w�&}̒l�H'Y'Rd�Nh������7�Nt�rL�ɐ��>7���d�!�Hv�%p�(�ԟ]���5[%!hu!�ɢ�(��d�.�&$8<����tJN��"?pH���'0�!_':�4�C�q �a:$Y*	Ҟ�����%FLa3�����&��6P��Ĕ�2�l�I�='�	����Ä�e�'�7'FD�:=�(M�L�pf�C��D�"u�(�͓��&���"Y�B&a�94O����DM�%é�I�hJ���ZP�(���H��
�M�D����C�L6O��D�c�D�m"'L:��[��
�!�D�$D��Da�'S�xO��M�U�D�$��-I����"q6P�h"'m"tRgIE�����%�ğ&D�,u	�D��z�	��:r�&u'D8��l�m�&0�9�tپ�N��݈�GD�a;��Y
D�|I�Љ�~ßGD٪8&��;�(�(�g�~k�Nm"b`�L4�D龤Ý:"=.����%��v�s"pI��rp�'�;B?a�ʜ(��}��f��Uu�*'F�D�Ʀ�aZ�sSf�r%7R��G
&�j#����*厧ɽ"lՈ�A�~ϺX�&d�}�mT�uu����ѽ�R&u;G(�۲�gv��G�\���bp�3�:T�����G0���J�tN̣�^�.�<�7Q2�`��NT��oܩ�٪ܞ=�T�g���t�j�
�F��b���4{�w�� ͕�v�<j%�B����jn����F��ؑ�}b�LG��ϐ�w",M�ψ\ϐG�Q8i�،�DE�6[>�2�"j�"�&�j|��DG���ȜjY҇��G�Q8kQ�TD�'n�u��:��D�L�2�"?w�4�(NF��7>DY>����*'
�S�a&4;$DzH���pA]JޤD]T��KR��� ��8_�ԡ����DM[R�2|���D^ԣ>I2�"wse�'Ȍ��lu���yQGY�˹�$DM��M2	�58A��p��;%�lj&�}���jQ����A�0HwMM�y>G��,�Y��TG����N�lD���^z��k��q1��n.O�f��fX�|�}{����J2�(��/�v�s�ݕ
.Dy4#�Ts�pEʉ�58C�͕B<$N��D~�(�2ښ;q:omM"ϡ�Q:e�Iʛ��h9��Aɚ2�1\�8�Ƹmx=�`{�x<q�%��;�;���h�; ��ra�85ڈ��jo6GUSBvښ᪉¯B�[���]�О�ByOx�>�8�7>E�q������eO������������}�|����g�P�h�4z4{Z+Gu#:���j�2�:Dz�=x�f��*&�nL5'MI:��#�Ty��Z=֊�Ei9h��z�[G�#GǳQ�;��.F�#�G��o#��)��G�!.Ѱ��%�Z�W�Fg��<�3PR�B�ɡ	���C��C��x{M�K�#�#}�����:�ay�.�=��6� R �=c.m{���C�2rJ5R�F�\yǙS�Q�xj�m�,F謴x0?i�i������x���*��l�sl��tV.F"��F�B.E�TE�!�w����I������	ѐ�6�Gn��[��4y�(h�֊����37Eo"8��$i6t(��h��\�:�:8��jiAj-�(O#̅���ے",�D�H�R&�WK��?K���"QO�0�r�1�8Wȓ�DGqܔ�0��kr��E�\,or�~{)���fߢ#���e�"i�H�bP���|ԤKu)��nV䯟��D�ܭ����4������|�R%����et��C��W��+e��DM�)J����g�JD�R�8��a��J�9��}�[O%"&؜.�_WΥ"[�I�;��,y��|�=�9�+E{=��
�<:0WjV8�Ҩ~E��2Vd�D�N���l�4&�H��lp�ԸX��`��X�`�n�5"%l���N��!�l�t8Hl�A*=�!�,��[,�}��;�Oe"�1����Xo"Ͳ�9D܃��'ȏ�9&Ƣs��=�ИG}�K�tG.�0N�ӌ��N2M���9s��藍Uq���$I�Xv�?&2�̐rC�K�䃿�y;�G2Vd�R���Z-���g�g���S��#
�	��u$��}I>һ�W%u�W��J�K�K�K�((WbU֖	Ȯ�h�5�%J$�RO���]�_rV��Ӵ�3�����t�Mp�
4Ѫ7
7f�־ѯ��Ni&�JM�+Л�E���h=�aV|�u�p��5(�7g��<9�f���������a�#d���/�|u��L��=�u��6����Ŋ׻Z���:��mV_w�����N�FrJ�>=�HtSBN��v���qq��o��@}��TN��J���x�k�m���=�F�>vsG�8��9���$�)�S�tو,V����qP\QF��4h��*����fFʅ�N��GOsʛ,�ǝ����� !�8A��Y���d"�ݏR�3�N]ܳӡ1lg�hUT�Ҏ-}�t��x����ll���°El�]��N�<|/�]���;��w�gN��z���T|!���U3m�~6~6}U��,�6���鳣�i)�WF���.�� U�Ai�9M���2f��EGg���x$]JC�=,��ԧH9	m���5�,�5�D�@�zmi����aل����q�Ę�[{�n��gQ��G�P��#j��\��,�if�6Q�l�.�⭲x�������1�O`H���t+;zcm0���U�>�ٯ[n�T�M�O��wl��ΖK�����������sK�I���P���5v��� U�p���d��sf����vir�tV����̧�Eh�8������V��-7d�q��=�t�iٛ�z�e�Y�E|�6t�Z�����kӥ<@|�鬪s�)�OO�Ҙ����7X��+~	S��6a!��x|%��ݚ9�v3Ц��SǏuJ̗F��� ��q�\�d��<h�r0�ȯ/.�Q���*��w���)�1^��e:=�x�<h��+`fN�օf������&���g3Wz׈S�w��424A��OFb��ަ�y۹���/>�! ��.^�k��;y9�8b�=����ݒl�'^ޚ(��:a���4||�pẞ���I���͟��t�.q��B���ѡ�M�4F'�1C�W:t��:(�4x�Ӥ5�G���螀�́�� V����V4s5�jυch�f(�F�cz}g��Ξ�,��*(���q�Η�pE�^�d��4���w-�dЁx� �3��I�O69&�-F.�h�Qf� H�j�ŏ���I�Ν����.�������C��;�sİŠ<pH��:gJy���`(����l��9�!u�}����3e83B\�c��(���Tg�Y�QJ�M� ��� �4l��C*ѳ�݈�鳦�i�<l�P81+�K�ԛ~՞1l�Q�EF��A�^h���>�!=@�ڪ�b���!ֶp�.�X�#>��O��ƻ�Z�I����!F?��ih$Ç�K/5��VP�D<sc U��v|�u�ӈ!���7���0���A5ɉ�>�G.<�����Z8Y��^X��^��n�UC����v�����պ�[NU�ow[l&��g�w������g�C�]̰���Ϛ8�˷�S� {h�������T�^��2W�:s�g��Чv���0�=y�ۡ�	?(p����'��>��^o웉wnN�bu0�i��g�ċ_#�K̨}�Z�5oT.��0����Vz���9��l���Ǐ����8�wsٜ:Sg���s�bZ�98b�H�'�vxb��7c3c4p�6���B��LT������.�	/7�����?���nCㆀ�����ND�f��k�{S�3f�Ĵl��[a=%���g�޹����1G���q��U����g�`~�<Z��̛!g�L4ps��K��e4FR�w�M��t������&@��><t�e45��l���eZի�Y��2�66f+�t��W�U��x�}�Fl�͜$٣��3sr�6h�j��7�9tsf�MNM�� �})�6l6��:��F���=8z�ʑåcYç�CǺ��>,�������:(��p��D�d(�՟\��
p�!����]R��~0���\dѳ�� 6!�Dv�kiѣF�����m�lѵo�U�6p�+� UGa-x��ݔ�6l�S��ݜ6���@�4Q��SGd����MEe�e�EvS��%�GN�qw�,�L[��,�l����ox����n�v�A���x��K��l'���/]:y
�^��1��QMP�uU
1�C%w:$��>��ϛ'����p�*5m��P��k�>���>8ۗY��Q�u�0���<�vY��/ ��@�Μ���}��r�Z�_�>��8Q��?��#�-X�5�:M��6�ך���e��)��� ��~6t�y/5Å�o�`z/`x
�zl�ׯ2��e>,��I�jp�HS�͐�����YbS���kg/��&�Q� <~�� �?M�Fh�^%N�:h`��M�6��!�4t�G6p�}N� qx+T��6<>���?nl����GFld �5!N�I=8x��I:P�d4 t��'���D6h���ˉtc4 U[���ɩ��-��O��A�Hg�S��<p�f��sZ7��&� �賂n�7�N��Zl�Ayٹ�7�K ���Y�pr�����r�K�@��81�7�ý��:0����
4f�C+�s/�G�s����1x�ᾧy%8t	�F��чK(�lS Q&cޮ5;s��.;7UY��8I�ʳ�{���9�����t����40)�W����^�9�R�x�@�$��D1/k���u{�͐� �N5��ؒ��)��y)��5�o���Oz���h^�&�W��Z��I�6]�/M�8Q�d a��9��Ӷ�+�N5��tl�����ttهO �7M�/K�-�F���wq�Q���i��2���*p�͜ i��xI������F�W>���tζ"WgV�?S��A#�*eS,����t��yQ�U���}O���z^z���"~ʔ|Ըߩ�����U�d���᳍<a��os<�sv������Wm3f"��� ZjZ��e���5��X��A�I{n�)�Kl6��������
:x�).(��u�)�.��ˍc�e[��@]�
��[OL�͛0�.���F=F�>�2��ce��Ř]J�N��(/��=,�_:tS��o+:���� 
���溺�����A@�~?�����{�W� �D�;�s(M����3t�ͺ���π'�:���se��)�V�:p�� ;��un�Qw;)�^�nq�TN�a���C���醍0��Zm�uU���qN��l�%�ۅ���K0�f�� X�N9#�J��km����;)���2�˶�oM1�$�J�l��G��dYEXP��"�^L�gN�O�W�G��w5�d�7e(����6l��x��,{�q�N��1�=��E���qpY���z��y\�*�5�2�� ì��I�9G�F�1�78p��W�\Z�����2m�mqDۙ7o��I�'f=�zl���03o�i��>��]$�叛�4����x�7_V�vV�z�5��8��h��z�U ����z'�]�|���$�����{��
_�%@�lٷ1Ss���q�~�_������H�v?�{�??MӠ���=�������_ (e����榟�����w��u�-.niN�b1R(b�m�н��g7J�k�" ��5M	��C)�f�S%�Ճ�&�%�P�H��Y�y9sѼ[�L��ou�x�X�������C]l.�N%Ͳ����0bu�+g�����X�N����.y�Գ�[��L �bp�lE1T%
e03!�d13-y��ş~ڏ�1x���\o�1�.����ok�2�3K�$)g[#�#/Kx���J^��¹�.�Xi�o�'<��	c/qJE[̲iu�z4�jJݡ���ǀ���	�Q��1��8��OoKJ��dBf�ͣ4f�P�� bcd�D`���0���҇�.��魲%�,l*���ڨ�d�SYJR�ψhI�.@k@$	��VD��ߥ��W�e�&(<��F��*�u���S`4]4�dAP�-��ڊhb5��Pi����bu܊��ٱ>4��ݯ0�o��[�Yd,R[#mW�o�Cڌ��fF[f��iYx����+�&�Mf��35}�6�z��-᫽Ht�o"�q�։�y��
���M
LKH�W�ҫI�0J�QB529�:�$��pVɯd�'���hYm�H�k\�e�`���m�����_�#g�&c=�h��50M��&�qpKZhB�q����Ε���z[��fo-��[	f"�0��b,d��%�,z5��i��,��!�e�g3���n;����JF�tf,��Kդ��1k�@Vě�r�4í%-W �cs��JWpj�|�W�h�y���^J)۾��IS\b9P6%��@d��r�!�ƒ���hbCgz@��t�q�6�|"�ѥ7��kGZ��C]ڔ�����\o��ɼY;���{�������E�J�/��o�ҁH�.�`jM�2�N��lՄ+�6Šȣi��y�s��5�-��h�Ȑ<��]�4.�)z�*�ԇP�`��;H.s�=���!�5'R��/��[]��s��}�?&���:�UT<�k�/c��Ȩ���w=���������������}�|�O�v�PUR�CY�f�����s�����*�U�Ux����iUv��iU^�J��b��"��������WB��V�Wj�V�U�*���U^�*��t��Uҫ�WjEU\EU^�*�Uv�UUb�T�iUUQUUQUUQUUS����ﾻ�;�H�b$��C�0�pD�J�JZJP�����R A"�Ð ��!B�@�A!��W���|>>�j�������1UUQUUR�W��U]��Uҫ�[U^*ڪ�ZUW�Ҫ�X�����u��mUx�*��UUq���ZUU�Ҫ�WJ���EUUU^+j���Ej�TUUUiU^�J��ZUW�Uq0~��$��B�J �X��") �@(�J�
D��
@�(D���}�B||I����V��V*���U\X���Ҫ�X���������[U]��Uv��Uڮ�]*�U�U�*���WJ��mV/��^���������V�Wj�V�U�*���WN1v��R���]��Uv��UҪ�WJ���U��)�������P�gV4�$J�i&���1&2�57����+�Wj���Ut��Uҫ�[U^,UU�UUTUUq���V�Uz����Uڮ�mUx���ZUW�ڪ�WJ��k�k��Պ�����ZU]��ZUW�����}�]*��mUW�J��1UW�J���޻������h�H�b#1^�P,B�� �h��J �� �(�B@�J��C�&B��:�`v�MB4B4����:��v��2E�
2"9�u(j ���w+�'���ߨ~J�E�?�����H��A�>��}��3css��rpvh��l�DD����dDJb'DL0N�,C@�hA!�,K!b%�b&�N	�:'D�	�DL�`�DL:pM�(L"h����t�$,�X�8"l����,N�f���HhDM���!�D؈�"Șt��8'NG	bQ�O�A:`�*I	b&����t�ӧM����DJb'DL0N�f���AAHJ��ͳ��sE|F�>��G��H45� %-v�r�U���2�v��m.�(F�:gfX���n�a˶M��'{�6���뼞?�a�k�~M*�Z�[؎���=hh����	H�B`l�I��"��kY���j�(9�X�7X�Q&Ay�3L�.`d��̺˚��6�[�bAJ͋蹱l�l�f���%�,��H̭��fz�����&��LA��Lj0NE*�g�kX���3]I�m=Yn��V[���0�ڋi����$�0W��Y�O�-}a.r[�uƲ�?~�޹43��9�kɣ�v~�؅���hV��թ����#`q�v@��Ϧ{ޯ��_�<���2���&��X����&ڨZb�V��|_��p&��]�^���~-fnif"Ԃ��	���.�X:h6�3��zҐ�Y�]�,�d�Ws)v��`:Bi��.�!X�u6Hf�S��������	J�Y�6٬�މ�Mpm��e%�]}L���JJ��,֗HYs���vv�ԃLX�Zb]3&�&�������Ѿeףe�%��3�����Sa���؍��Q���ے�]+�U���L}��Ef5����-���1�P�ݭu�i�-\@&�͵���Փ����4�#���6eZj�#�֙�Q���6"u��ʓ\F��V��v/��@	-�<1<iB�.]Q�в�ڢ;6$t��l"jd��5�)��(Fͬ.,�X�%�-�ܗ�{z�������1l�؎ɦ��V:ܡu�{1����o�è�������k��)D�C�7�K+�M\mu�" �ѳ#i�!SWbP�i����9��L˰�����\b�j�B�Z��D���V�\��t�P0��׭}�t�ځ2��;l��z{�=,�]qC��WZ҉���{J��ix�/6�b�\G��Z	����
�hVS��{��,G�v�ѹ�֠�3d1I���A�v���ԉ�%�W2�uV�,����$D�Z�"ۍ�)�^6v��׶Z��o׽�����Rˁ�#̕��C+��g�s#�w[�QU՘K�]�J�0\2��I��u%�[�Q�%�x�{�P�_��[�#���ufnf�Rݭ��2�ْU�GW]u�x�L�X��2��flcHdؒ���.Ҏ�e+a*�T�:L]@DX,+�N�[�B)t�B�����g{����-��]\��-UT*KG]vG)9��k"j��B�oM2�n1G�s��LY��uuα����]mՌYhꩰ赳F���7�ͱh���vp����L�O(��v�U,�tm��i�:[4`�1�@L
[�:�L��=�X��J#\��@P�6V�\B,���柃���� ��d1Հ=�BR�e� �6��6�1���B��]-�͇"���Z��j&]\e�]BX�Ќ�B[Dz��2�@3.�k��bZ�G
6��Bm
鮌Fks4߳=�C�=b7Y��.�&��&�V%�M�#5]z�K�n��idٖ�u3!�8KaHj�5(�2��RV]�[Y�Mx�6'���ޤu�%40�s`@1fn�]�l�u�Ccii�j��t�^&�,m.�B8�a�KD�,�K���ڄ[��q�eh�n���3/hP�-���,\X��e��#UPE�PZMkQ�i3z蚲[l�k�։�+�����m ZYR�ө��[F�'B��Z�B�����[u�B:s�pP���,δ�B��6�lZ�c�2����V%�l!,�l�Mɩ*k��q4.0UFJa�i��	�Sy�m����hANV��ZZ�
������5U��t'���T�.�k�Yw�bp���.�!�������P���a)�ryOR<�v�q@�l�i|j�ki�F���q(��Hlk���f[�������h��l��L��C�q5����F��z[e�S�g�G\���qj�z�A�c��Ah��ӟ�g������y*���WZִ����努�UU�*�ֵ����,UW؊������i������U}����=�{�UU� �Dh�4�I4���pDLF	GD�t�g�������gH�$�URF�e����+,��@�4tK/	.KPsv53���7F�/]��0&�lS�$mծ���-�Zk���d%J[i��&�u�I��Z�\b�\]��g��V�����!��eW�J�t֒�js�Yt3��bj�m�	wZWl�h�Um�[qI�m��168Х���Y���:fԱ�l@�W6mG+����]VY�F�Mb�3i�]�zԵ1/�{�6%���ĭ�t͕���aX�f���b����U��Bݔ�WtuY�`n����t�����4��g]]tі��K�ͣa6c[�rfl$�^y���n�.t�ӅڼM�AKu�ѧ,̖�f֫lqhYtQ��<�B\���I$����r0���ܪ�R��f������s(�͖7M"e+9zUh����dTqjO� Ӻ}T5T�H�kl��)�4���;��hw�&j�J�jCUY��>'�?�������oU�qB_��,r�e�.���ɳo�y���Ѵ[�UDo��F��4��ܺ��Q%��8R)X�A�@܌�*��5��Qd�y�q\���4�� 	$bM��Y�{�uB�GOD�t��j��DQ'����2��L$�(�?�<x�⎞ ��F�0X`��Q���g��8[����m��G�I'G��i�2`���_���g�!nݤ��I��F��@���q��!@���~ ӚH֚H-n�*��8AAh���!\	��>��-���6�7e[��爲�%����A�X~��`}��J�'�D�4ZtC�YT��66�
�ޘ��$gJ$�Oi�N<&	���a�:p��T��۪���n۔YLQ	� ���,|�m�{Z��b�H����x��q�\C0�ƕ�JS���pt���&u��7�6�d��w<��[�;�Im��5�4�8�ô��#3�����9C-2N��d�6+T�%z����K���U�p�LPakKD�"��q��4�^��4��,�g0��0M%`���7ݑ�.���d�G�$�+�i����FE��vA��L��Q�a��Ç�p�^^�#��LX4
0Cq�c���[�.%՗r/!�h��dF ��\�rb��[Um�W�m�=4 GPK$�I#e-�;�\<j'�j��x���/��_`Ȉ�Ϟ|�m|`-�߮�y�^�p�0@��X4I⋘-�6A4Y��:`��bC���`��L����b%(!Q%j�5�4m�R!{����5�DF6�5��n!]ynͻ$�],tI$��]���[�9DF�h1f�c�ܹ��*Ww4-�A9��Ӭ[B�Z��)��n+��]Ks76�D.��wcH��Q�PP�r��c(C׮qi���%];��y)��txP 3�9,H�6������:V�8�:j$l�,F[�mǋ��a�.�#	�dL�=E��+Q�a��#G���"b88]<t��}�$���$�C*s4~��Kb�hgv�q�h��嵶�O����vy�$��1����TJ�~]�i�m�yV�6������t�����&	��a�,�Ƙ�5vj�{���ED�1���m�Ӆ��C87Ћy����^ɞ���uy�I�n��]��h����g�\�����)Q|F�"�Y��Qg�DD#jA�ѵ%��G�0}�o�D��R&��p��NqR,�	/я�@^I%(\\,:bgo�гt�K$�	�0L��0�8YuX�^�كm�����v`�3����2,A�$���J�
.����D�8�!&�V�H�:H�!:0]k�]�XQCPdY��u�ϣ�8J 4�E��m��6<1��]��ME�w�Z�vX�z���m4�-�k�8�4t\0���b$�$=�(�{��D#��Wq��Rp���,D�r��C��q�/��d��F��>���4C�<Y���Å����`���4�Cb�Qh8�3"�q��f,��u&+^��s�9].�&��ɽ�����xu���c�[ST
U�6h�jU"�?w��{)G渺��fp�`V�I&�d����1̽|9���\��؈
��t��"`0�IhEL  ��q1�E:��4���gN�G� 9:�K������RJ8���.�g�>�� �,�gM�8"&	�,4h#�(� �h�Z��h��]�(���m9��*�7D��P��[U��� ��~�\C6��T=[y�	yX��m<�٩�^�����­@�̩��������Ё4�s��f]����q�C-8����ٽ�b�m�:1�f��,�`�`�w��:-�`��p�z�m��:�����(�*x/2n���U��pe����HMpA��1q����,�:a�ey*�NQ�$�^qT^��1�('�Cn+ƫ��F�^������s���Q��
ƊX�B�dLA0)���2�_����)��0�Hg�C1h�"�B`���,�
:`��8!Ӆ�y;?�zcmuU�eUF�ù�`�Ӯ���������a)h�k��L1�C���@H��ޘ��B�6�0���j`;�Î87z��1�Ȯ6�F..��Ͷ��Dڃ(��$��</`�t�F��{�M�m�S���G����U1�'m.!�^��mi�|M��4:z�GJ�;Hn�:��5�:3Őxv2�h�;0�n�xr=	�di$=�'G��p�zC4��G���8i>���=�!i�o���a��/�dυeDx���G&z��/�H�gá�@Q�@�G�s[�����4���Ό�(�g�G���8O	G�$��?G���ȁ��4�Dh�|8F�G���za3Fih�4#GC4�=o���#F�xiG���:i:oH��3h�u-Ǎ#G�����=8D�F���I�h����={<GL��pzda�_-��C��j�|�*q#��^�"�Q���vdFT� �����*��֔A�H4��g�H�"#s�&<WJ���4zIl=#���������zx�N�|4�X�!�CF͆���#�G���1�<�F���l	���|k��:	DR~��q�"GxѳA�U��x���WN��V0�V4:EU��*8��LR��4,����G�}��NAu����yj��&$U�z8ve*�\iike)��LkY�����k\�!)Ř��K"YB3?UzT����L��ߛ��z5��U�M��kTQ�JйuT����!l�(
��4�UK;B%�rF{@�;T�|_N�������-Ǽ߾����?{��ފ����wo����̙�����z{�Uqn��}񙕙���g�=�{��*�ݾ>>�����{��O{����*�ݾ�>�!�af0��"`�'�0<"Cf(���h5�g�BY,��N��c�:�[:���1o�����(dD
GS13F%&A��LѠ���c* 둢���q�ԕ�'�<�5,�$�a�h=v��.�m�b��,�G� Z!�^�RyX���a��)=Q���Ρ��ΟyY�@��ƇD0�p��Sc�1$����	�A�;$l���w��I7p�L�<�s�u�T2@xK���o����"��h[4l�ַ�P��>b>)3�j!th<����T�����IG�$���IC0�'K0�����0��$0��.��(ɂ"�"  b!P��0��3$~%�M�T��%)JƏ���!4S +!����L!�~�9k2�C�F�a��e��f%9$u���"���lA���Ɠ]֘���Oxr��p��r����������/D�5��G[��T>C	�1���nTE���K�Lw6�Z�7��#pb�Eq}�.Q(�Q�,!Q�bUg�����AѤ4�2*�+�)R=��r��q�F�)���Sw�:%���͜Ób;��MRd1
(g�	>$�G�>8x���:t�$0������&]�D�d����T1j�'Zږ4E�%T�<՚ܗc6��v�d�L0�����LW^��� �	 ��8��|�d����Y�_8ޘ¹yDm��Ћ�WY�{�ڵ+�ce*Y+f̴"*�����Y�7ۋ��ꔍ��*P���;Ͻ��9�y}�]K�f������Z��_ ��^�ok�-޷���peS���n)<143D�E"��I܍�=l�&�&��$m�`��<�Mt��qƨY9��᠆3���m�(F��;D"y4)���8���Z�+)`�)@0�SRH2�d�1�8�8#h���w�I&&�:0�v`l�0���2�]�C
C7�Fi7�Dc'�D���8 ���"D�q� �"�bg�Aϼ��QS13b���1�֟F�R0v���aK�!#
s�5�DH�Q����cPv�1�3*�g̔K�%�����������`�:	��!���V�Ƞq�-��H,�39aw%� 4��<'��I&��T�!�$7�����OF�^�e�>�w$�������R��`"�
P�!��h�piH�e� <0���m�G	�	^�<�4m�� ������3G� V2�	M�BLv��$�b�/)yz�A��ǒX�>q��,|!�ͯa��@�X�h�%��BT0��Q�$�#yu�r�7��	9������b90*�H"Ɛ�d80Ph�� V4H1�O6��k]�Y�p"��,`φ�ˤ�$�A���H�4�ň�?���"t�&x�
8���z&&'��g�fhV��qm�_� �HK:��<�N~k^^B�E�zH[C�҃Jm���J�0���v]�^Ua�6��͌SrS�1y`4Br��郖S:�l�I�"C�s٢�Ō���m�].�κ5��A�$��1 �|;I�8`�5�I�8"�fK���߂ EY��]�p9�����1G��Ē4�4w����Ób7<� �7�ǆtb1�刌�bG�Mn��ԛ��FI�A�w`����ѻ<�`�֐�7 �\H4B\]癫5��5�s®���|$r�>���%P����Ը�KAA��|=yzʤP�d���<3�0������8"&�Ӡ�a���}�^�����lc���F�&je3&ƍ(���0��3Of�$"8�3Z��V��=�~�*�C$HMJ:@h�PU�N�4A��1�x��ض�ѺA`��Մ,�SI�M�C���T�2e�����qQuS�[勩@�,ͺ	Ԅ$�!*b� $�xm��tp��Aw5��!�f�1&��Y̲���к4���B�������I��)�!Ө�6`���E8ؘwU$�շW-�&hp2�}�T�3���(3� ���Kl��|8DM�$�KF�ѭ+���EB�nF��C av"�AG����#�m��>�]��ē����X2�=�Fcp����8l��ag����pDL�A0�H:a"��|#��Wv�b1�����۸�mC�شS8i]򭙡��n�ᐫbhOJK�"�F�.�H�h$�H$�@��!�-���q��m��O�T����[�oQoω��j_��۲C�t=7vUl������&�����W+�g�"Y�H	����9@���$�:{y<|�w�sl�DV1�sL�a�Rg�hvۊ��r�&g���rF ��������V���9L�A�	�&��;0�)�5۲�Fzp�D��X��i��E��(�筚)L��v�D�H$h�.�:�+��oTK&bj&ғ�xd��c�F��9�T���o�GĄ�D�%*:@�PI�'�Ȱ���9�A�4�:0r�E��D4A"��@4F��=�&1���CF�m����4Y}$6�P�0v�!�'�����k�*�;4��I(���u���4H[��Q�f)�	�9��\P���qE��6`QC:|I��<l�~8"&�ӢC<Q�F�"x���$ �IS��A$@@�ex�`>�
S��j��4'�v:|q�%�-�R:aц��8�1��ĶA32a�:Gz���D卥eI<04�*c��p�8���5�ZL<0��H�4Ƴ��ht3S�o�|���@X�P�z�|)T)X��R��-�B]�o���n
Ǥ�j��H0�M������N7%�ڄz�e��-4�|:%b'��\�11��JgQc���\�T����V�d,`���YY6�}�ǋ�B:�,DI�J::C��<Y��l�����"'N�WWɮ�(��~������```1(B��M4�M��I�%����N�9\Te��}p�)�)�Fw.~��""Eч�0�;t{���Ǔ:R(x``�"�WP�XR��DO"Ϊ�Å)
����Z>D�!A��ǌM�Q�-�\y��8�5�dn6��D�P�\�&�7e�y�WV8��$�L^H	5�㝞'f��N��,t�) x��|%Yaᅦ4N����12.e�c��@���%\%-V������sI?�Ҍ�#RH7���(Z���+D���O8q
Y
�Z�! 5p�4pg|I��>>8"&�ӢC<Q�K3>����_]c�x�3��}}BY!'�/�M�����A�A�HtaѠj��TUE�K�m)V�"�6��Z;��)r���Z���jD�C)Y�G )<)Q�Zޏ�ߗ�%�ta=N�E�
���y��lC�f�8��Q����|V��80�z���� w'�"8Cn�_e4O��N��"H 80&�#�12�bi|�c��h���:�{EZ�)֘Ã�H�ōڼ�x�i��R�A*�4(�;��vP�����i�z1ҥ� 80$ix�^ �+���E#�_����$��$g�]G�T|Ag�2��>��&�ZE�I���6�i�4z?\�#F�#G��/Hќ4����~�Oi�4���9�!���f�٩����lz63Fx��F~c>,�G�/�X?�Q��9��4x=��aHa�	G�����,�>#G�������hΘE���zi�pp�G����=0��ѐ=&���p�G����4e�Ɛxg!h�ޑM�����Y;�d3H4tI���z<4�4�N@�Ѝ4��F�N�H��z3[�<Aæ���Y
��������$��z<7�z63F1�8C�GCz3FH��$f��D�₏a�&�����x�?G�4l�4zI��#G��������A�H���ѱ�3SoSl�1�oA�6=���2F��b�eU�/몚�.9��Z��bI�v!b�|՟f�N&�UC/��Vwz�&�Db�Vd[�n�L�I�(��#�\�������"�1�}�"�+����ѕ���L]{;�e;lf���!CD����
�I��3U$�5Tr[订5��EY.d�T�1�	��0J�N��*�W�w+��R�n���Z���>��@]N]�un��T��M�uʗ2&�������BO]�\9�� ��]OQ�X1�=��HLܣa\)��������u�1E�c���jF�dͫ��&v8bH�*µ�Y
�.V�9z7��!�
;�1�v�����.��?bڽ�6�-��J�Uka���,��Qe6��*�V�]8s	B3Ks`��/�|ح�iv5ͺ�`��X��Tf#���Yd�f5k(���W�����Ǜ�6Yh"�՘�Ԧ�U�����<@�����ߺ��{�����wv��2�33���������-���32�3=�+J����=�z���>�̼��{�Ҫ�����������0�6x��0DN�]]B��qy�����G�=r���N֩����0�lүe�,̩fГCXV��f�.Ք&��Wh�,M��Ԍ
�Kl�c�V�p��K�F]2��lm	��W��9�! &f�2�l��ݙ��.!���țf&��kΤ��^�:��mHͬmr�(�l���uڰ�;Y�ʪ����.��s��0��]�\.�\��CY���cS�hZ��X�K�}](_!} L���1ZV����.�42�M6n�-��_����̫Ip%�*�]�k#nm��v�iv�����T[4&6ѐxaVۨ�R.Ԙٗ�٥5���˝��e���ͣ6�Bi[mNx%uY��y�hCb�P0l~C��Ԧeդ(�[���BXZ-�kԽ����c�l��\�!,�3�g�[j��W�tc�1&��Z���TgJ(�T_8l�U��ùZ7�{U7�iԎ���������ʭ��g�՜�"�9o�AX�o�_	�{��7���-r���N
?��}E|��6}�&O�]�����|4Ɠ& ���P��B:5|�[�\V@���D% Bj�]��`�XyuR	������n��V�&�����$��nz��U#-��/�O�iO�m�2c�XխD�6�����R��̹�%�$��bhƸ0��R����� h����8�!�:����*D��@����_)Tu��+��78Z��(�#q	m	k���-i���]R��D7�%/	��j,��*�4��XBe$@P��X�clvݣ�w\CT��
�<`�0��Ox����"'N�0�O!���>��c�$iɤ&����1�bM� �� ���I�&wN�zs�,a#G!?h�e�Y�EP�k�����uy��W5w.�&�V�:�>G�)^��%+�H�J�jᆪ��h��� �Z��Bd"�eJ)@ҡ�ф)�(�h�tm�5����#Į���
G����a�14�YQ��[�n!Èq�|�^X���Q8�vX���&D@bf�ͺD�0bk�y�@�,�4�d��%���C�H��Q�-d�Ij
�%C#b������R�&��D� ��d3t��?�0DN�a�8��lAD1�L���cz�޻]k��&%�0�:�ȥ:1�c�D�:���(�l�����~�@i4��wQ�R�Ba��M�^�d�J-J��L,a��Z;
�T�A�{��˹&�D��Rx``10T��AF��ϑ*}͚������~�"�7�Ѧ��F��q���
Y��J$���p�Lbv٥���Oiy�Pۥ,F��(�d.�!1)���d���!&a�\�`�cC	<|��Bm������ch�&A�^UF�N���&:0�9�0���(��� ��i4�!�%4�<Q��t�,�Y�M����"'N�.��q|��ߗ�h�BL�:1�c� ك�tFKq�z�Ã��2^��#�D�(*0$���CO:5��avPB]E�%&j�X�����#L��T��C�Hd9�iqh:�4Da�����b:c��3�Q�ЦB�n�P�j2���-I����T�L:Sc%�%7Ip#�C�$��M��{7p8'vCd���8n�»���I	z#46�kYWTO$B�����$m��hp��������4��f��ġ��D	�ܨ#�q4��阛,1t�C#��LC]0��n��k�1c��ܗD��9���
 ��'I>4��Nx�"t��t��{f\�sN��n�D6} q9WX`�d������#�}���O�5ɣ�:j��卤�.��c�$Д�/�7�����道�VM�N.˥i�;u�ea�5�fs�v�cʺg��\�%1M.K.�]�������fol�w {P��~���g��;���\���x)�&����i�'���5�n���6��U�n��W�1��>E���:�E.p��#
j
> �f&�1�O$���A�+�	����D�液w7qܜ�����1wk�"dm���!2�8��-(G�K%@P��dc��rD8!��BP�IӤ����#T@�A�ͺ��u�ƺ0�����H��ɉ���1�F�-U%����5�ěb!b�.�DAGFX��[���J8p��!�Xa�vx���rCѮ�."긢��B\�r��N��*" �ŋ��4�,���M�0 ���0�Gs�VWp�d����]SK��٠���a�BY�6~?<"`��:$0�<t�9��!ڭ;���z�(n�1�I�%�����>-�2$ф(L	S	T���V�*EH⏯�吆0��,��H�����#���Ӿ;fx�tL�����W���`e�����K�Lzc^:|��:��Q�mƐ�%H�	<���j�?(!5�>D��8 $�	4a�G�֍;��>�?�Hh�mب��e�ciG�1�t���b�iD%~D%cC�������LMZ�f�,����vc:5��z�_�F$��� pcI�<��P�E`��.!��ߣbfb[�s6j�
�D�@QD�x�G�?6x�p���"t��t�N9�3��f�14=��)JR�BX��k`���?o"�&��3BD�K-|��0� ��y�8M@�b�J!/���9
�H�P|4E{1�q,�P�e!�,��cv�4��
!6:%�z䴚�2#3HH����R����ϿGl��+�lg5���t�\z1�i�v���2h�M:4�]K�͚��ﺟ5��vj�x�=mv�H��5��|M��)������� 1�A�L�_0��8��эYВP�CJ��>�c���LqZ:�b;E�`��σ%�!#f�:a�A�^��������g{9�@id,�t����l�~8x�"'N�:���V}M��"q��2�N�4�i@�61�c�BJ/ɤUQ�`�j�z��R�`�,�d��T��x��B^��{^�;��]�t���UYE])��A�P����i1�ǰ�1M��ӲK��[�u�;���I̓��O�ߪ(4(�'IJ6IJF�Rg>o��v13�\%����A� d2��BjH?��XZÊ������`�P�ɩBU�Hh�ˀ-֋4�&I%����4�H<�&�4�I!�A)�3�j�D5�tg�Q�F�||p�D�:tHa�:xy�/.��m뗹.|��z��ϖ/���k��<b9�|�y��CƗ�ls%�ѱ̐���#Zh��1�bM ;�,wv�6�;U���υ7�t��c���νŎ�q�3���]ujv+d7S���wy8DN����,���֗��j#済���4SOm�:�b����;x�9��\�E7	�i:$ߺ�x�`0�D�&p��Y+����C$���G�.�qq����0�i�DA��(�9���A�у�U�Tr�ni�D8C���l��E�%d�Y�jZ�$���$: �T��5�K=��69=l�X���`'d2GN�W
�B�
��TB5@�P(V��w�T�_�i�̌?��0���N�Q�i|3��JX084�4����Ý�:����8���ȁPx�ΔaG
:|Y���M<t���h�F�P�$�TmBDr2�Δ�4Jڹ��)���1�pa�&���h�'�.�Ē�4����224�q�`ƈ��&�Ρ/�_4�$��F�]�-�5h�F!��66��{>t��h�D�N����@�*2N��N����Ď"O�$�A��!�Q��Q���J���Z����LD%A�84�:�+ (�Yn'���.OԾur�w|�;�Yw|h�	M^X" �鍤��0tA��=��m'Q�i07I��y�fp�y�}t���19LSn��SrM��Dr�^cͪ*�N�h��s�}(�ȃuACCQR5�:0�e!Q�+4�ψ,t?���2�i=&�/H���4z?&��`z6il94�������޶�=� �nG�r=M�4� dkm�jm�i�1�F�h֌��֎�iD*4�F�z8h���?�џ�����D�~�	P��D�O�$<D�Bx�<%�:CG���<x�<Y:=824z3G�����=�h�(��ǣ��f�#GM�4�6��G��|p���|f��p����?AF��������=,���Y�h��4zp�tz?G��zDoH��i�[tB�H��7=�I 4�l�n=m�z63F�Q���٣���-#��$hѣ��- ��H�};/�t}0����*�f�����t~#G���7���~��4����7�1���3F�h3���62�Hφ�ț{\��@�8�e'�l2QZӘ����B�v���9I�L�϶�/N���z �ZH�J[R�2Y:�z����m�+ �Kh�G9t"�ť��2��Fv��U�]���D���x�����x����R���#�UTpC�	�[+g;�Uu����Է�uҳyF.V�gi���؞�j���'�����+�!��*�j�8a� J��������+J�����뻿p�̼��{�Ҫ�Y�{ۻ�o335����mUx�}��W�ffk3=�ڪ�b�޵�o���a�h��<p��0DN�a�:x�r�Uܬ��1�4%�B�/��b�a�g�ÓX�A�x�<M�xx%1��c��K:0]�6f��4�$p4X�Mju�,�"�a��I�Gpa)&��6g��9NE
�)|��t���x܋��Ɵ �õ6ԐncA��ɯ�b��ϣN�ɦC ؔ��i$�8"�Q<��0�%�b*���1�O1WX�na˱3�Ϛ8H�|t�Hc�:�Rk��rCP�sŢ�	�@�4S0�c�5F�S��RIQ�W�j�}=�M1���]>�â<w��,d҃�"h��B����ĤPQ�>(�Gx����Ǆ�:tHa�;�+䅟E�K �#	�>V��)��F*#�E��bߕ�h����X|���bc-��êJ�D�mHp��a��T1��d/�*�I#[pr��]K�1<����m�߾�H�F@�P3aH����)<] P3Ǜm����C0j&H%J
���L��<��]*������_<A�!gs|z��;n
��B��*�.��f|�D����f���Q�%�!�,�͵ґ�!D�4�e&B7��|�a��"��7[�bjFj�ȘD ��)^�v����TX�(��(��g��4��Ǐ0p#F�3ҋ�Ŕf܀հ�6���Rո�C�<�5�ң&��ֵ��7t�P{��ό��q�D���WL�_�V�����z�%*l3.���	 �	/W���g�y�suWڮ�W��pg�`�F��	�e;i��P�K�+`����.��L�r��mwKw�[o(N�fww��Eiz��:L]ϣ��6��C���
|h�2���љmӾ���p{�{�Q
���hm�P�"&����+�T�B��	�W�)�PK��!(�LE��M���ZHඋ �@�M4a��g("8B�{�{'%UT[J���g�|R)�#҈E���k����|yK���R��V#d����F�\Vq)6O X��AO'ģ<�x�
�,�8�,�>!r�fI�8�,�"p�4!�F4㘞o�~MUp��F�D#H	�6�J �D"4~D�ZD��I��L$��Ni��4��<3�Fab1�r�i�6v���O��~}}�/w΂g֩�D"�,�|�)"�h�|P��ICK7��H���}q��\I4�GGj����)°����3�J�K�#ϰR `p��yB(�T��L��qi�J:0c#э�9F�p���G��ϑ(�P�ӿM�/ȨY���ū�Ww~�8E7尊�Gk�1��h�D#�=F�b>9�Ҵ�tc�Tq����)�&Pቐ�ᢋGP�E��>"�(8X�I��4��O��<x��'N�0�KI�eU�-�'�Ж~��("ޤ�OF�m������M#����F���2B2�E�B%���F��G��d�eb��{�S�gmuF.H��x�L�J:�8�]C͙��U��}$q�AQ~�ۛr�^�;��whb�#��փ&i~��;�m�*
Ě^�@j,gh��� c
jh��	Py1�T��*`��90�v�!�GB�9bz�Xϰ����GO.���������}Sʶ⦇ɍRuk^G�Y��(�cl�`��ݶ�V��""Q%c(��|I�N|p��4Ӧ�<a��t��:�2CHb���ism6�m6�4/�5�p�NM'��$�rF����5T�	P���O&{"�T/�kd]�j2�Sq�!��Ld5uHZih�EJT3�)� Y��+�{���1��j!G�
T�.�4J%E�2����U�R�3�����ڟH�T�!�8j�Q�B���~�{�ߚ�N�R��4��"��yd�L d�ωZ���p�h7Ŵ�-R,fJ ��v6�f�d�L���
	 �:I��t��O�O<a��D�C��ʣw3TN{�#��6��z{�'�T�7͛C]�B�1�5�[��A$A%���oqٲժ��U,���«��rM�'����F�+w�wUS�b$©el�]l4����tթo<�s�e3��<�u؎1S��Ǖ4N*�"j�w��6���$�uRb��}�AE�YKI�X��4�ч��e���E�>$��9#I�d"��yt��[���1�V�3��B\p�T��	�ɢ��榈�8���d�9���M���b1��<��m<4�K�a�B ��ƣ��b�>=�IX� ����M8���Cw���4Ro�]a���D.���i����+�U��~�1{�����h�
RS��Y��K��N�Q�R0��Y�'Ěp��?<x�:tHa�:w�^h�4ѡ3]�Wc@Q>4�G
0K���ƛ*�i��i���3xa��(�5R���Hpf���O&��E��&�\�I��3���?���6F�Җ� �3ˈ�	Aj�e�)*r�0���M����z�"����s�I����B��u�ƨ�(GD�"�(勵���I�|}�Dr6$����#�6��p�9h�#����q����R���\���H�j��Ä"��p�������8���X��\7�Z���Dt�9	:I|Iӆ�4��M4�0p#F�0&*���e)$�Dk�" ��"=�6���K�8��A�G�6p82���1}g�]G��DOL+�O
0Le���F�v�p��up cfH̢B�h�]6Σm�vFQE\@ȉ�
����H�qH�.-���_(�(�����MZb,�k�:DH��_gǂ���p���ѫ�t�T0�}��DA��"�5fEDL��Hf���3ǣ����Zמ�!MԦ�Q�)�*�����/��`pcD6@�;+]\F.�HXa�H:t�ğ?C��ᆚi�O0`0c�s�Pi���HH�����E�4�� ����i���"( ���H��Ȃ�v�D'�XP�cDgf	l�1�R����
�őN�П=�4��Qej\^8Ã:5H� �j ������a�z��X�"3��Ŷ�Ӧ����[~-��KG
D����a˗0�I�Ou�}M��Cx3Q:ϻ$���q3�㡃:.�:���}��13�l|d�&"��ʫr�0�Ý[�x�sᣣ��s�:5C��
:B��e�Ac��l��~D�I�q���zt�6H�Hc4zA���t�=�l���=m�����c���f�57$-M�m3FǣcZ3FkrA��[�h�і=ӄiI�x�(�A"C�Q����W�����)!�:P�+��+	���=�G:8҈ӄh��I��g%�E�/�xlc�x[���t^ �t3ƖO�A�-�� ���t=(�FH�zA����4�4f�GM#G��diƏG��h�iI=o�h�F�!q�"�#L �H(�	4�ܑ��?�!C�&|@�����/�aF�ц9Q��d�F�z8,�ђ=�]4�vGG��|:F��Q�1��e�Y3G�m7��l7��=����C��3A�Ѷ٣c4�gH4lz62F|62F�p2b��͎Rt�����V�"��U�2ʦE\{��Ck��k�<�d4�,�p��ȼ��t1*-\*��H�t�Ff���˘�*^��{�ʘU)������/���\[!G#�����hh]ܔ�]`�|��/�*v*$�ueSO�U�Ba��hۃ����W=y5*��r�h�K	)�.�S�C.;�'"��ŕ�9d8l�IR���Ց�Lv�L]�}c�4H���yP���ݪb�U4qU|�e]E#�y%�̅��D�ߥ=ݚe��I�G:��yFtfU7�(�1�-S�D�A��Q	A2������.r����@��8|iBWD�RzW\᥻�$�ԭ�����{�v5������Me)��nu�a[V��]A�TT�!,�N�9"I%uٜD�+yS�F��������j�Ŋ���{y�������j�Ŋ��ֽ�����{�U�Uⴺ���k333y���]*�V�^ޫh]�$��J:IӇNi��i�O/..%��-�#�� 9��B�A,��@5 ;-�f�7[�-q�e�K\�?�=_1ڒʖ��M ͪi�ը`v�]�&�xڲ՗]11��*�t�(B[GY5uQ� ���R�F\Z�e�k,���8T�&1
&n�ֽ\1�n�L�X!,��t�#Ńne�ӂ1qc��YL�M�V)�WA�0�-t�4XY����Yll�8���MWv ��2�Ζi�ml��C�kOB*rg���:�qM)El���Ɋ�kX�k�Q&�4�3,f���X����,dl-��R�%��Yiڵt\l\�y�ۭ+m��Y=�r4��\:��^��%�MZ�!$b�Ml���:�2��I].0i�&�j�-�#�e�������f�C\����Ж{��0��PȦ�o�*M�+uV`�7�x����W(��v&�Iڻ��)F�o��N9�F7�2V��Ԋn�q��ʻ���DX�a��D���+Uf����Ń{�����h�M��`�L��3�Q��%
ߠ�E"�Y�u��0z��!C.�E2�f@1���z`��2��Ȩk� �R���W,a �k-���b�����6{�
�p%-�܆�ƾ!!3�����i<0c-n1�ڨ�4�/h��x�Y������mI�I$��Ͽb]B@�k:���_���3ȴ�JFO]�Z$�H<pҬY�H0��I0���O�4�Ox� ������i��[u<m\�3���>�i��i���5[�އӋ�3R�YA�H�r�5�q.d�qj�QgF�nǠȇ_#��/dR��W�
3eI$қk&K���GL�:M��tlI����� �e!�e�����T�sD��&������'娅`�@��Ll�����l�G�gA��l8n5Q��x�]��E���;��]�r����IQ�O�p��4�ƚx�®��t��".�K���� �@:���-��FM>�f,(_#�,�cJ(�t�(P�\.H	H����}I�5��] ��*�r��ʪ�
�!~W��I�@O::�#��������*�5��<A��������?�g�:���cV�F"�}�i����C�)>�A��1����&F�<A��Mɡ�'y����CY��o��xgE#5bQ�_#d@@I��(ҏ�:t��Ƙi��4��d�����k��X�oA[I� DB d�nD+=݃��,Rt��+�]G#�D�^�ٹ�j��N�e�t�W�"�1̶��U5��c/
xi��F���@P�#�DQ���vj-/�tg�N��v|��Å��I���v��uV3�1��6A�;&l�Y�q��	���WʑkhØ��a*�՚M�>c��vE8�o���]G���d5R`�(���>8p��4�ƚx����s�C��2n�m�т�JI$��tj;5$�%^;GP�.��Ρ�pM�+6l�M���A$^��1�6��Jw�u\m�כO7m.ۋ�h=�6b��]ۇ\��w[uy2G�%u��w��w��_;�)M�/��#�^�}*�ݝ9	���v��+\n��WZ��s6�7.M�&�[�RL4��B��@�֝���*�m�}8���	G%c���d�X���HPɴJ�Ы�>>Z�(:1�p�DC$�o(�iB�	HPǿDzbS2�"�w�x�+��q�����L�lZ�\��QC3�|o���]*u��xd�D��¼7¼��p�Ǚ#)H�:��&UU�̍�%c�b�L���x_���;:9M��5DE��\��m�!� :5��7,
}hs��gɍOH�<A ���Q⏏�4��M4�0��pqחH���q5q8-,g���,���36[����ʱ�
��(�v˧$I:�nL����P~pk�}V�nn�Ku|;!+�tx����3)�7�0��.ts��:��@te�9vg��{��5y��B�,�#��g�QM�����̚؁��d�T��E���t�V���咋�D�C1|%+G�F=!�Ck���F��峎u��qӅ#�җ�a#0g�؈h��z�Zb�P�((��4�M4�0��p��>�u,ff���K���@ ��]2�C�fH�(�pq��^$��	�>�F�PgDA��(��ўL�:@2Q��1�1{��7-���Cؠ��n���g��#��:8N��{*��6�LdI�]Gy����Lxm����qF��1�mt�����_1�c�"�8���DRg�0Hΐ�����s3>o�qMQ�r����3�(Ҏ�9���M4�0ĸ���ڒ&b%BEvڬ�V�i��J�m?��X�����N�JZӿ���Rf��/���4�1��+�~��y�.!.���j�(B'{��y/�Z�8���fA�"\9�Ƣ��3�m�Z�P�@1�#8���Z8�Ӆ#�,g���ϧ��oS_-�;�o��阞���R)a�"�c>��ݟ[p��xp�8�T3SE�~]F#A�6Р��:Qҏt�N|a��x�O``�E�wAH�OZR�/�d`<w�6F��=<����ݥ��k1�����u���ʟ|�I�Ix D�ѯ��ʼ��R]��Ah��䰜���If�ern�Ŷ�M_A/ӫŻ��P�՘W��*ّ�v�����·hSHI{hun�Y1!ˍIwp��u�Yˡ�X�f0�T]M�YX1h�*M�!d�y&U"	�[�������D���aΫ��C�H�8y��Le� �}�:�q�!��.r�F��dh�o"�mt�n}�Čo�ѓ���;�b;��c>D��G�Z/�I*�]F#��v�1U��p_.b��_	�I@����K�#m6����E�-�iA�"A����N���# ͅ,V鄰��h$u�Ã<Aet�O0�4�ƚx��)�,�������$Բ[�G����M��M�M��U���ͯ��x���y#Vt��a�Rpf��(�B��AZ�r��LA0L/��c-uX�%"ݜ\_#���G����9��H��m��-�:�cB(d����J")6&F2�8a������-p,ce��c_R)�)��#�`�����G>9q�凔��p�z`X��"� )%H�Ex��$�O�<Q�id<���'KD�"hDN�`���p��f�A(ADJ+�&��4"lD��:&	�L�0L�hM"lL:p�DK4'"a�GA�M���ɣ"hKBh�,�$DЉ��&4t<x��4x��0L��BhM��%�BQ,� �A
:B���Bx�g��!��8t��gO:X�$B"pKDL6t؛,�A�Q(��~'0��j����|c+ �/wa'y�S�l�6�f�>I�{n��Q���]�C�{x�gP���`�)S�|V��DDK|�e���*55p���̺���VY|2�]kG������F�{$&�e�@��x/(ܢ��g����5�c/`����u<�#:�H�w-`�W=0��X2`�ײ�d��et��
��򥽙[ĺ��o�iUҫ�iu��^�fff�=�*�Uv�.��kי����z�]*�V�Z�������g�j��]�KU�["�ѝ ���:QӦ�a�i��4�38w��\DA����z�IJ(��,|7�ۀo��s;H�(��t���I0�aᚏ����#���qΊ�_��vU�\�j:�W�o��4�B�����j<����F�&�����qqV�F��<2NN|��$냢�ߺ���y�8(� �R��U����O��a�Dw?i@}�C@ ��n�l�4��4Ã�4��W�j(���4Q(��l�aZ\ � $�ψ8|YG
>><a��i��4�38^>2ZP�/p��:�[f	/���@ M	�S��m���10�����{���:|�9'�m;GQ��F}O�4�#Ʉc�`�r�&��6��֤�"�r�Ť���;�I!-�qp
����a�K�|�E��3�A����A�@A��ǵ���:Z;4�!ђg�!�+\T�E���}�C7�ڋKM>^��0���Y�B���,W���@�Ro��A�t����2BH�<YF�t��4�M4���p�����Va����B)�"��Q\�p�0Qq�	�}d�Q�Z	q�kS�/� �@^�����*�:Y�5klU`FYWk.��;�Ϳ`��]�l���0�kj���:���73I���5ۤ4�Oj�.���Y.��c�+6��8����*F%1!��^"��3���$�U��I�d8�j3���<P����Py-aA�C��K�~0������\IHБ��T���tL��«�F�``��R�-p�� �q멍�������"!}�Y����(����(�	7�|���]9t�z�`�� ��w���/ˋ� U����_��E�<���O���d�,�Δa�L8i��i�M<a��m��J�3N.���Y-����w�@ �u��}��f���u.�P�)ɺln�i���kJ�]���xZ�R:��K�K�r) Ӑ_�k��b������XjL��'p�)�x�>8��7[� �PvQ��
D����� ��A"[l�?H��2�U��Eԫ�X�HE"�U��\��mp8@�T|a��/��,��8#�К ��R�!a�pC$�ω,����<x�<'N�!Ҏ��eo�6ҢH�L� ^m��D"k�j!�C���8F�|b%J�OD�5�}1J��Q�|���N)CW�2F�C��N��i���P�R��.�dׅxa�2��4ϑÌ4(���g�a��U����y�L5��>�Z
���߆�Z�.<a���R�޹�VK��n��DTĲ���
�}�}��N&��蟃��B�(��s�3��IC(���Y:xÇ�i��4�3�����C�QTۣ@�
2�[�܂"�"!B8��s���y��3����@�5� ����Gs"��߫� N:���y
|� ��)>$,�&�j:�=����8�<��Z�(є�\��c0T|��|F:VIgQh��F��|n5��#��#�/����!\��������yx�3�t�I���7���6����c e�Y�K8Q�|a��i�M<a���L{�XZ�LW�w	KDͻ��6�P��ԍ��"�jT��- (�QE��@�&Zߺ�I�Ix!��މ�� ?��S>�hp��X����H{٬��8&hqN$᥹u�pCX�}�.�J�o�umq=�@��9l]�ܮ�P�eG���nv�w�U�p�z��t����HiS�(��{�j[iT@ܣ�aR��-r�&��-���Ѕ��w�T�4p��sg��Z��&AF�D+GVYӚ�,�Fzk�wn�	L]��顋$�^>c���K�Jt��uo֩P��5�Y�K�%�iAm�_���)��ſc�d3]�ҋ�_D<m�Fiw0�3[��f��+T,��S���Ǒ��FP2�i$�
>:i��a��x�Oa�0��`7�	��C��c��h��ԑk�u��m��&��Ƿ÷��j��4�MH�C����g!������i	πB}_vҨ�$�%&j1
�3����;���9�m�>T��'{EBA�QK�^m����⣇Ԏ����kiik�^`%��x�B��%&`b�'��/ܥ��v�s�w>Z:��]ŁgN�ǖ����ň�`�T�;��4�0�2���Q18�^H�jK2H:Y%�Q��|a��i�������[Z&��&
F8��g�τ �O4���;@��~���f1R:81��PIh��GA�p �Bjt|V�Y�<t,���D�|>�|��Ǯ6�h��BRD(:�ѷh�yg�E��JUP�ah����5Á#*��l��z��������R*00�荇3K"[���"iH�Ӈ�NR�Pqi��yR�J���,�GO0�4�Oi�0fp���4$RF����
SM���cSa����y��1 �@:�l�}L�:�}NWȓ�g8�Q�X�"s�_�LQ���--%�ÿH(����°u���
��ͭ��$�`�8����E&Y�6��y<Fp���XQh�}Q:��)b8�,�o4���}p�i�1J�ju����D.��|�($�����a���Z�:P?7�>����+G��1�yY�Yh���t�K$�^&�ƍ� �"%����t�"A4"'DN�='6YB �	� ��Q�4%��b'��0L6a�:"`�'D舐؈�tN�(D�"hDD�&:h!bX��:""a{$6%��4Y��#$D�4""`�t�>D�"hDN	B`���<p��4x�(�g����!�0����B%	�!ӆ�8x�Y���<&�D����DL7�lM�P� � ���X��$��-�e��iU�C]�fӳ��*��j�M!�m�	��[4���,�7B�i�5VE��<�Nu��<[�n��,j�n�Rt�"�-�,��W�U�^{,_]U����m��"�u�Q�`��%GiWY*5!��h9�7<�F>C�C�{P+6��e҆��s�s2�p۬Jr�Z�W\��sO�M�ߕ�V1s�]D�6䉎h����㊒6)�(�vE:-�X���}nO,M$�n�xs-��Db���e�}A�ė��Z��9GK��k�Z��z=Wkڅ�[���5U+줒w0�J���������7���S/���Qk�|���	[�A-���"q,>��1<�k��t�h�5�r���T+��e��M�C�=��K��׶�����Y�hoz�Q���1̷�v�B96oOy9��ٻ������Uڮ�mֿo^�����{֪�Uҭ�ֽ�Vfffs=�U]��V�k^׫3339�����t�n��k��0�0��O:x�Oi�0fp��"f5����\LYGk1���E�vu��/:�%��6�.�ck��\��S8�hjJJGYl��`B���Dd���(uձ����ulvx��/׸��]�����:����Y��|#YI�;MfkPoY���t��!.�nSf���㶘�F&�������SWf�Ѓ]QD��4���;F��|��Ol�&�p$��mB�-�jS-h֡k��f�K��)p�ƭ.,
��ҹz���mHҹц���I^+lF�Wd](1+,f��;]�����zf�����u�e�q�#&�.�GY�5���i�yk.乺��s�M/F��Yc,tV�#5׮��(��6���=�3n���ls`[�L��A$^n��5;+�P:`���gfP�Ws3x_B���A;�V���Y3+&M�;טE7l���m=�S)Of�9S�ZYU�Q��^�w��+zo��|2�������poB��k�'#j]�֖�_��=)6|?��~�;�`�,,��P��ke�,gHVx��㈶�c7�(�A���J*��$� �x�tXo��`ll�pD�g�G-<�6�:A+���7�O#���5@���A�� 8ag�R�}�`���-"\����S�Pt%�Z�_���Q�y��J�"�~[�u�3:t��
>:|a��zi�M<p�a��1��p�w�t��yk,��W��Ø��ga�����{�DAD"j)AE#TR��{�队b<px66��(��*�X�M�V���)Q0��Ԇ�h��Ն.#~>E�]M�i�sfl��3xb���"�Fxw���3E������Qn�V�&�u�4�1ǥ4,���Z����V}�F�X��%R�0e�b�y(>8�d:���ʠ�d��|p�O|pӦ�x�O0����3h�Ka��� �	 ��B}dC�p�N���PAըg�LZ4֜_[����uh���b0�c)qq����#�d��<nN��+�����mK��.ݜ�����G[����b�_.|:�,���-4P}M��g��,�R9(�3�W�=����?�%E�X�H�~�1.-0�I��֑�{W���>�و�:Q�yI��D�2H>4��
<t�8i�M<i��`� ��[	�4�h$T���u D"3ô�7膠�#�ȓ4P���n���|8
~k�rH�)��iԩ.�
mėu^:5�<��[������H �|b0h���5�Ű�6/�*�B)Sv]�����q�s39�h��u�R�S/S�T`�����}5jQ�t�Jf"��჆��yK�ϓ�Gk��3QH�t�Գ���>!�k�Č�$�N>0��:i��4���9�٬�����ī�lܗ�&X��˧�5���4	�B@Q��~��@%�6׉a����� �	 ��@�LQ�_�sw�ͻ�qaU��8��i�:��n���;������f������vY�m	{�jU`�+lAw�n��e�'���W�q�=�{G*���K�jZte��>>/șJQf*R�'᳅"'#��<�t(���-�s�Y+;L�JTZ�1G(,��@z���.�C�3K��,V�G(�i:wI<����:�I�N�4|R���I���ߓż�M{dq�i�ȭ����Ak�9��vG7I�a���� uo��r-�'�X�^#�G|.�<�[��Y�I��<t��:a��4��0fqDLF>8up�F��A$A%���Ibw��xo�̂��Qk����\B��]h�':I՝00�a!(��u6�����F����%�)�"����w��E�'��8`�ç�6h�a|Adb�C��.�c�X��rf.���9��a/�PA�Q��f�����'*̯����]9��|ߋG�	:��>E�I��Ψ�ѥuQ'C�C�,$��A�$����t�M<i��:`� �&���|�-��|ʞd�H]d̬�0�6�H$�IC6"�!�����:5}o���k�ľ<�����xӫ�e�P�8�ۼ1��_"�h�S����e�$��v�Ъ����׻�ԛ9Ϡ�դ���nB�������AR��>8�u-��l|$:v�7IOAc{�6����-9ۧ%��GN�8�C�pp�*tA'�'���t��<xN�0�v��P� Ji����PI�fba���0�6�5OF�t�����禔���	.�p�����"�jr�5,�o�C{�����Z��~5|��m�������H��d�r�hl�I���ldLӤ�Qh���R�d�R|�,:��Ě�Z�7�!�ؗ��q~���6Ɔ�mE��P�-F-Gx9>��E�i����26ўp�w
4��e�[m��Ջ�"B	�p���a���:p�Oi��38o:A��S�uD1\�!*?Q�)�gEVDJ�W`� b��9�rn���7u$�Ɯ`�N@��4��A$A%��O������u�)��4k�f�}φ"�-���s��Y��U������,�b��L3�RT��(��#a���SN!�c(�FG�0���_]Bn���5�ozNG�q�( �̍�c3�ҕ���(�1%:�*T���V�G��S $���"!��RL���_Ė|I���!1����<U�#��V���������	GxQg���K q���#�:41�D�>�; yu:b��6|����J4�xh�4A�h����{$�2�2W�++��*+�g9��0��k!R4��I�8��0SӇ���
0���0���:p�Oi��38P�G	f�6�m6�o_�QD.�&\��ܟ#c�A��҃|��V�����!�LP|�IxWD:��-R�G���i(MQ+T��XI�u�"�T}���9�q3LFv�û�]�ku��ĺxI�O�<�|*/���ZY�o`��k���O|�+
�p��Q�AF"yh�Y�����F�?$B""`�(A���B`���blM�� � �p�"QF�dK�M����`�Y�`�&	�`�&�D��6P�4""tD� tD���b"tDD�8	�blM���A���"ɣ�"A4'N����lM�(ҵ�Z�A�խ������D��hJ�����g0N� �<x��ǎ<a�"a�f��e � �	�f�ek�6������\�5���������ݖq�e���1#i�Q-X12�'0#�M��Ŧ���]t��
�F��n�&#,0������`�jV�5xv��Be��Y���ˡ�F�թHg+:��퍨6n�ְ��`�W#�9u'N��E�Щ�t�ȍ����/�{쯷���
x�{����w}�U]��V�kW�L�����Ԫ��[u�_������Ԫ��WZֵ�L�����Ԫ��WZֵ�O��a��Y��:a㧏x��<xN�a�p�?oM6�m6�]}�F���G���ǁ�1iK��	e��ê�x���Z��s�'�9~�Y�.����P7~� �m��L�o�)�����1ɹ^M��z�ޓ�h{(�<�_��
����iif���ˋv|3���T���+���_\̾1��	r��׸������]�7��wŚ�jԎb/{���x0��,���(�0�Ӧ�i�M<aӣ0�7�y��`4	7ؚFA�ذ� ���mҷ�u��m��)��Ľ������t�z�!�DI��g�y��_t��8*[��S� �i8LP@�8X�}���4�-	i�zM����o��KJ�#�CF�8dr�ʗ >G(ccJ�fDD����d�&�%P'�	8Bh�s�O$����1T�Ԗ����p�j		>%�i'J>0��Ɲ4�Oi�����d�M��(�K =]���
폚�L"���U�ꩆ&0���V�֞�E&6�^�K/�����lm����y�k??A �@:_�.��+-j���q��m�r�x;�ϥ��v)Z��r��-`�>w}�/Iɦ�&��Pmpn}�*f֗��U�)�\�*�ӯN:=�
�vL����ܲ��*��+]@��>�|2�E��~+��Q5ڢ�
���/���ɣ��K�}�+��ы!���l{����ۈڈrU�>r���1��|�fDC�D���՞Ȉ��R��<�G`�p)1�c=" � Ll��|>�������3MH>TURt��T�����p�s��Æ����o���E��6��F��D�I�:x��N�p�ƚxçFao-��E5(z��R߼�!�p���r	 ��E�>d�o��xc|>)|�+��hpb&�ck�!��5�>k�قSU|A#8�U�H�`u[��CG���j*��a�Ë��O�K�������B����%�fDC����}�=G,Rؘ�/-�{��5�3�C@zꩠ��h��j��ta�h��m�7G������0�"���&M�m���uJ$�(��I�Oiӧ�i�Nx�O..��q=�HX�j(]��M"��3�h$�H$�+m-6�|'ü�N4Т>��Z-x��h�zw��0���,Z�CV�m�����|K_��q����Ѫ�MT"��1���gFA�������}-��5ՙLm�l�����1�N�3���h��,)5�AiQ�et��G;�Cz
zqOF��=�8X�$�'�:|t���N�i��4�N��o���ܧ��/�羈џ}==Ѝ�G3��FT?�s�D�6;��T��51U�(m�3�̱��Q�ǃ��)�ߢ�&P;Lg�C�6��9c��8��Sd��hv��J|zZ�%�-��FKqf���g��kaǦ�K�-2)�k��J�p=��7�:�$<�:A���x��U16%�ЃI�K$�Ft�Ɲ4�i���8�q�&�p��8c�Lj�k���[�P�KDD��L�����O2��1�x䅸�%B�)�U�,�nG\يk�����~
���A$A%�p�ID�s��؊�/�˼�gٷ����u��>�E��]ea�֚�y
l3:��*��as�����B�c=Gm�$R�u���QA��L��t*�Ɛ^�!D����T�X�R����q�1R����(��J-a�Ђ��C�Q&���IR��O���Py/�T���_�,�A�1R���|�M��p�u�j�:�Q��#��Ê0�j���AѶ�A�U�EuMQ�h�Q�Pb�9cm��+�K~�$�����dM���6�Q�<LD������&�w�.�;��8x�	0��>0�Ӧ�a���yquu��x���D��kM����&�IӬ�t�%�fC>�Q�8+�m�7�P�UI5PW߸�����Y��\"W��"�ѧP�C�tjѶt�>�Xӈ�cm6ؘǈ���$8k[��R�3��W:ߜ�3��ȣ�*�:'�7ya]ChYg:�m������B(_J$-�A��|aV\\�)P�!���,�<`�?0��x�0�Α���c�my�e�d�V黄CF�����{�6�m6�}�4i��1�F�1�)WPx�J �԰1�#���xƚ<��hY����U�Z�/sH�7]Hܶʚ��2g�lcn�ٮD-]\^:�	>�����4|_��8��E����h����_u)x	!���\S�h���K:�����]�D4�t��<Id�Q�ӧ�t�L<i��:tgC䭗��4
��z����@ !��=��S�n2�GQa�0�Q�j%V+F�:O]c�Օ%*&���q�����Z��O"�)�ZB:y:]G�Q�����;Á�_���CD��Ǖ����U�6�V�1�6��4�E&��Z)w�A,�5լp�d�蘙n'|��:.�*5����a'����/Z&ш�q�d�	4��xYf�4A��0N �DЈ��0��؛,� � �`�d,�BX���pN�&`�tD�0L�`����:'N"p�B"""t��D�ı6"tDD�8&���,�`�Dw"'DD��"A4"'Lf	��tM�4X��(J<x�zC�}��x<	�J����BP�:l�Â&	҄ ��:x�<x���l��< � �x!��Q��*�5!����Y�B�c\ؼRu��	�@i]�۲�H�-e:������B_136=���%��(q�9���NF��1�����z�=ѣdDH7���G
���{�����K�P�ՔS�P��ɇ�`J�ua��f%��EVӠo�\�m�V�|�V�
���:<*Ti�q�&+���K�_^�8�h�Ckq$�R,Alai�"�����Y���z�mS��im�(�u[�요����\�/E�޻�����Yq�}.�T� ÷�ha�Ub�8����꾜Վ�qb˝u��f-��w%G��^\���!�����a�V��ľݿ�u�5��fy��VVP��,ߎx4s�=���}>cZ�m��A̳;;:��#u�]�ooz��6��j#1�B}�u��*�T���iX�m�[rY��rM2N0�I���5��P�`�m'�^�[����o��?���g誯�WZֵ�L����g���V�]kZ��3333�誫եWZִ������z*��iUֵ�>!�af0�<x�M0�0�ѝ8I����9�d�⠹�jk�t���Օ�C:�\���kU��%�0/[eI[�e�;\Ԩ5�����9��+�ul�cp�kfE{:]�K�bÖK+u ��-�m��ɻg@�ٷ�nhjnp����;+�c�CW^!2�fk��]�)4�"2����]Kk98�&�3]]�Ѹ^�-�vɮ4�lŔŬ��)*�@+v�q-�%�א̲�f���7E���\Q���2�%Sl��l��
Bݜk�6l&�K�]KS%�e��J�����sBRR��c51[��4�YF�lac��1�FǠk�l����k)I��`���\8�em�l��`f�n��m(�i2d��)[I�If�5��f�aaVU��m��R�.HeƂIrR�S�� ���K�^�y|���v�W,����OU�G�n���]�q7FX9t�CJ�T'���ʱ�k�7Y�����b�u]]��z�����z�k����P���4[tx�8�	��Ģ�L����� ��ģ<>��4�!j�"f��
dD(�Ť���s�mÂ�Kz�_��)���1�p��{��1ܯ`p�3�m��Ԝ
	V�Y�3J��:��m�Ԗ�l����1�AQTDTT�kk	8�<O�����진��i ��I<i�4馜<i��:tgNs�e�m��˸rBu:�9�9�_"���ۆ66�E��������$(:���J��^��t[\�6650a�OR~Z���u/��F@�PQ�, 7��)>G��I
p0ľ=*%&l7�!�6|�KAq�m16��)�{��4B��z�ǗkC؟�"�G�Wމ�\��N�Ȓ�(�<{����]:���Y�d�ĖI�><x��N�i�ƚxçFt�&g��%�e�s��X���-:ߦ\̎d~F#�qG.;4hs�j1Hj�1|�T����7��1E�飡JS٦+[��5�~��mEMVޛ5s8��V]���8�������g���[m�u���.��%t�����\C��Ca�|��Y�8��b��|��l����u�b0$��x���Q��i�M,�0�ѝ8h�*�e1nX��눢�MG�U�*V-����D��)�"(�j6��q�U5QPJ�PT��<��
F4!i$/�ѸpZ(�r�M����5#G������|R$�C���30��]�0˯"�}��� ��\i�p�D���$ލ{[уŁ8�;�@�Y|T6�1`�E���,�0��<x�Ǎ���0h�F�`���ս��T$PU*��J�3T�6�Si��w-�.��л�fh�v�Ñ-t�Ҏ�/��[�Fk���������C��!۸>����	&�ӧ\oJ�:�uۥX:���z�����(p��a���͕�Ur-gA������_GC���)a�%쒟N�d.h�O�O���~���X�Y�r���Ed*U	r�B�|�F����}���l�WXܸXL��8`q|x���8�.�{GzigBC9��cp�!$>-}�,�7����Qd����؋��8
`qń!�Vb$�A�C��QU.u�hi�M� 
Kix�{�2�#|��#�W��
�����EC�Y��<pOǌ<x؞<'N��umD= =H<�BnF��H��llm��Vr*�a��zt����qH���(d.���˙Q���13�M4I~���7�7����b�
p�F��	��S:�����&)�·l�'IC]m�'�kHc�8G$��JY,t��_`�/�8p�^AH-�"#�p-�D���B�J�M��hN'Q�U���|��iR����/�G�B���8Y�О<pO0��bx�0�ph�S�֌3Y��m��4��I�����!��qA%��4�ǎ�G��N>8B����0����A�����,�;���`r{�Kh=h�i֞�,n��uuU1~���H��|�L�0-b�#]E+�42Z�(�� �|���ƾ�ѳ�苹�,����3H7�d�s�Ȅur���u�yu�$��x�ĘQӧ�4�	�Ǆ�Å��*Q_J�VY�QE�tO'}q�c��w�0lx��q��߂���|�YiW��QZ6&���ʶp�nGy'�a׋�9^�Gف0�V��ќ!��i�o���G�r،G�-����5�h*�����Q�Z�&�6�����)�`R)d��!$�p��1�%�C��n�2��.�gEвFad�$�G�M8i��4�Śi�F�4X`���.�7KKe�C ���U#�SY�S�4�p��iJ��.���ZP#`��f��4����Á+Z��	�|2C*�Ґ��?�c��p�5Vޝ|8�6�|ȥ|4GL!)���� ��T�T�B��:6�Ѩ굖��krл{N%��1�/�@���w3;Q�V:��T�ʚ3��^\cD��l()�r[LsI ����xPl�F�K��G�1��IaH�:5��T�NT��p1G�>&^Dn6��&	�qsx�|~�qt �F2ױ�p��Aн}�����Ӻ�h��x#F��-A�w��1PO�`���F�ڋ�\�dL�.[�8�4�>"���]�&t>R<���yY����p�ĝ(��㆚i�M<Y��0�ѝ8IΚc��dq'������L)R�*��&��U��DC����p��G�O:1��%Z�5%��:��n�>J�<|��d��)%|�%Z��3���g9O�j8�'��Tk�ˋ��x8�Z���~����%�oV��`�Cc`}��#�b+���A���jO��0�Pt酖|l؜4%��`�DD؈��p�D�6"tD�,L�؛,��� �"C�X��Ț�M�����&	�`�&	�`���H'N�,D�B&�0N�A0J(M�'L�lM	�bp�M�"C�"lDDD�
DjDGr"9"`�:'��6t�b_	@�%~d����O<B���ؐ�8'N�:p؉�p�D�6"tD�0����e�x< �<9<^��>��"��'��O�,���5�+$F,�lIZ�
��Ōmy<��ge��w�0F���Fe!�T][�j��|�UU)��`�6jL�3��b*[XZX֚sTͥ�ﲮ�U��I��G�D�Ղ��i�e�8Q'���Z�7��nTHS!l^��[�z�aI�M��&Q$�V���{�pA�S��oJ[��b>,�#��XYU����U���9���UΝ�g}���UW�J���i񙙙��"��V�]kZ��333=�UU�ҫ�kZ|ffff{Ȫ��]kZ��0�afa�<p���<&��C/�i��b�غD�rCmG�gP���45�L�I(#��2����=����aJ������-f{5Խ��Z|뵖tz#is:R�yB$�u����
�0�>�(��/����|��	���6���<}l�J�����D!�� �x�j5����4��(f$�'�4�4Ӧ�xӆ�0�ѝ0�L��G�� -�#G럗�|��  ��0����x2�[�e�S�0A�[r�]:j*2��;}��4�o���U�ݯ'j���+l��e#�E(]<R�4��t��)��#��2�x<iJ0�Z$6Z���"����@��c8��6�+YSq��è�W�T��$��,KF	㇏0��<p�4�3U��%c�R(@Q���4����q
4Ye��(!��S|ɼ���ƢjVFY%d���H)A1���ջ-^� 	
��4���Ҟ����c&�Ǚ�yzJ�mD
�y���K���t��v�ye�mb�B�7x�!O�b��t*�7̢��Q0��Ȟ��[��
������r�-�Ų\��%��+�>9d���p�������xR!I	��\�w���E��Д���]Q�.*d�a�u)�8��`��0p|6�BB���;-��)���GK�.SC���bwŘrI��Z���1��CCTֻ5f�V����h!xW�A@A�ݟP�}p�fC%�4a��<a��x��:aѝ0�ɷY%4��T>5���]¶��^݋��oO� :��m���E,�dba/a�:Km�5�/��9�R��2��=Y�Y�EI4u1yR8�G�8���N<�>���w�,��Ф^T��'GC��.�b6�R�V�D��f�"���.a���u��٪N�1x�C���gӤ��;�mY�\�EQ&�TN��Cqȍ�)�C�jЄ��8>��k�`,��4��M(�M8|'�<xO<'L0�,�s�3���UšFԓ���^� 
h@����^��q��u8��R-}f�C~ԑ*���\x?�њ��i�Z�θ�����pM�E�Y��6�G�,D���/��8�8�q*�%Ϩ�@�y�<�gG�N���2�m�c�j�I��Q��{��0W��vJ�E��ڰ8q}!e��D�I�|i��x�Ǆ��t�a��zor�L�-3wMqn�5b��� �����'p����׋8t�ʖ�J�W��&b�s8��UMۧ\ݟa�[he��EF��R�DB\8Z�e"��Z�]��7��׀␳�oE�"F����\s��*�]_b��}��.xq<���~$h�J֮�+m�E�~Kz�+\PB@p:��i�����w�!�yA�0�4<X�(�	>(�ǎxӦ�x���}0f$��e�+�Ir���)'JZ5qm3P�)�d�0x�kB����{����M�S`[ �pt��rVT߼ �s��>�2)�e+N�9(��.��F�N��8A�U���++}4��s2�����:�(�F�e^������9_��"[[�6����+[;�5����p8py5Hhӂ�
,�`����oRqa�"�i�8qw�q�ǑԛU����-�N>��T��:���{;��+�|�1{�у�\<���\<b<�q�#���V��-�;C-q��,k�Y�P�� 1�>i�B!2H\J.�WߤK)���d�3>��C��������ihŝ���ң�����p�L$ҏ�p�<a�M<i'M:`�8J�L�fL������m���5���� �q��J?�7�@��I2���ƣI��V��ҟ�QŴi�Z1B����-[><.+%p�F��xn��/�J<��X��Q!	��Q"�
����n�[�p�sUL!�&։�$��y �R��=�ޢ�g���g�$�B���"8��dh���G�(hoWoz���(π=�/ئ(�ʡS6Y�G�?<'DO	�<a�[Q\��3���(}
�m�3Kb�m$�� '�OВ5�1�:Qc^V��4q�A��8��,�鄦����B,�K�i >+b���b&o����FՓh��,���X��!%��`��D��E�!�Y�����>�~�V����Q���7��|e��f{]�&\��������H�.�p������A�JO�IE�|I�G�ǎ�rD�(��C�&˻�ޝ�M7.��x �+@*��_u����)�B�UqB�mz}�Z	iT���["��.'��s8����+��-�x�}T8�C���X���"!a(�l��>^���8���!��I����|��|�RE�Į.�li�Q����I	A��>�(h�4�_���_��%Q%}5PUU

���S�҇�����L
���l�4]�`@�!
` �h�����Xi�ʩ�"�H�H1 ��քv`��f �f��0& �	��`�B`��&"& �&��`�B`���f �&�&
&(&	�&�`�& �f	�b���H&	 	��H����	!d�H�$�� ��Y ��$��"& �!�H���b"H("$�����	� ���Ya�������"&""b"ab$�bH��"&"$��SA�PL4�a�B	"""H�$��&!�H��""$��& ��$"��"b"� ����"!b$���"���"""%���"H��""H�&""%����	b"b"bX��@8DD�$AD$,$DI�D�$,�,DK�DD��DD�,D�D��D�ID�,ID���D�,DK�B�K�D�$DI$DDI�$DK,A�D�,DK,DBD$Aı,��1$DLDI1$DK�$A$DLDI�ILD�D��1$DID��D�LDLDLDL,D� I�I�I$A�ID1I�$DLB�I�L1ALD,�1LDL111,B�D$A�B��1I��D�A1�D�I��D�1IB�D�J��D�L,D�$DL�$�A��C$2B@@C$!$C$D@C$2A$D$A$2B�$@�!
@�2�0"�����@Ȑ0$(���2$��&@?��P�� aB�� dH
���a�b�"VD	�00$�
@ʐ0$�*@Ȑ2$&*@�00��(��(@ʰ2�	��2 �2�"2�	 0,(@��(2�(2� ��@���@ʰ0��@°0��@���02�+��0��(��,�
@�00,"��00$# @�0200��@�00�(�ʐ2� ,��#)"�H@0�"(@H$*@H$�@B�Jd�PLA �$��H @B$#�@�# �2��C
C"C
C"�0�2) ���0��$2��0�) �CC C+�$0�0�2����0�0���ʐ��C+!
B� C#��2$20���$2�2�2$2$20��+!�
J�#2�����)�)	$`�0�2C`���
D1����2C�2o�jP�C,1��1��3B���32C�C�C,1��2C2C2B���2��C,0C$)���C	C�,����2��C,)�C,0C$0C$0C$)2��C	C,1���C2C�C���C,1��2�2Hd&B�CC$0C,1��2�2C2�2C�1
L1���I$K�A�L��0I0$A0DIA0DA�A�A�DA0$�AL�D�A�LA$$A$�A�� �	 �	�$� �$� � �H�`X`h"`( &�`�	��N���"	� �"`� ��$�$� �$�H � �"	� �( �"`�&��H& � ��H	� � �� �CP� �L�D	0DL0I �$0-0�!04��2@��$�,�2@I$@2@I$�$@I$��ր��LH�$��� d���H"�H �HH �`I $��HH	�� $���f`f�6��`Y��`	���`��� �	�&`f`�" ��`& �	�&	���X��cg"&	�&��a	��a����B`��&�f	��_I(z���`u��/��xC��G��(��  *�(D��Ǔ���>۟�q��������Oo�!������o=������~/�<�_p�h�_���w��+�}^��p{�w���[��<��׸6:��_�������c�����k��* �w���~�?_����h�(������(
��"@����'�U���|�b܄p��I������c��G�>Ͻ���>�xF����
�}"������@}<&�'Jhv�~��K�_����a�2�i���I���I���
��ώ9��9���?��0(�>o�7M���Q4����~i�&$ �{�hDCB��M*⠨�
�e@�Ea�U�A�H��QM���1���ݝB���������o���{��� �
	@D*Ђ- �s"�&0�(�P �*����~��},�����������c�<������8 �1�0�ٿ��~������\�O�`�@O��u���?��G����>������8�C���d<�3�_���� ~A�]������K���??~{��~�%��O������+��z]|փ��g��`w�r��?7B{�_U 0/�}��������	_�������ր��t<}�Y���֎���p�؇��ww\�I��~��|O�@ �t��:T�#���>��3qı0��Lp��TÀ�,��;a�3��;N?t���z��H"�.��_���<E���@���q�#��������k}�>����������84���N����>��:C��'��o�� �������?O�OK�̠* {�v��<�!������P :����O����ξ��Oc�? ������A�><��R���A߿���؃p����}�{���������u���A�p�{.ηe�~�C����~����C��j�sO��x>���.�6�������������}��s��f�:���~u���P�@Q�fW�k򃣏��������>�äP~�Cd��M~_�K�}��r�I�y�7_�~c>�>�����>���������"�(H�S)�