BZh91AY&SY��Y�߀pyc����߰����ar:���@  �	�    �  (���  =�נ(iZѢ�Ѡ @��       7�=    &�
      � �@!�0	�0���   ����!���:H儗�R.���`�p%u����y7`}����|;0� ;� 
s�:%Gliݛmlr 0p=vǯ{ ����\�v 8��f�>�    #�^ ٫�y�C�>l$R��Os��
���@����v�@0;����Jyj��;b�{{������6�8���T�o�Ì�H׻�(����p
�9ت]��p������Eޠ  
 �`u�	]`+�Ϟ�Aw��P�pk���u��x����h^�=p
��ڹ���u���;��; ���{ӷ'(���Ҳ��uG>�<#G�r�P!�  � ��:��^����փ��4;pѭ9�P�ܶlu����pu�v̍H� !������2�}�$o�	v딉۹��wh5ہ.	s�:����<�π��   h���{{lD��ϳ�� �v��Q�U��9áƍ9:D7�A��{�q�a�Ȭ����'s*�����>��7ٍs�!�H=      (��         ��                        ���T�F�b dɂ4�	L$$�$��=&���b`MCA)���R�0F�# ���	��jd0��Iz�A�@�4�  H�J�4L$ƣM�5?@��y��)��U<���ICF  ��� ?Q���+�� �#�46��?�_�����`~��T ��&����L�P���@Q�@�����O���nU@���UT]�\���W�7�Y`��Q��$s�b�Ҁ�T��U�u����8��-�V��ej����k��kU�_}�	pDE�=��ڿ�����l�?�{�q?����>-����ύ�t�~�+��_�xk�9ӟ��#J �֯ƳP̈́�	���%��,ja7J�W.�0��O_.��wr#p�B�YeP����-3�܉wҺG+��N�% �K--3MLJ2�II�%����$��rR�!/L�+��y'	KLLJ�T�(�ҴC��zU���K������	$x���&�����a �'J��*
���	�}13��+�$QVu=�,�t�������0��1gJ�R'n�I�r嘙���Q""{b��FcJ7�t� L!0�M,��Oē���A"{aȉ�	��A�Q�DL�&$���������Db(����&�	1	�u�G����DKDp!�%����S��DGj;g����e��Ky�;@��;�bD�B&"t�s9���DȄG���xn8��=肄�B&%v0�,r%'!bΚ�x�Ȳ�	G��@�O����D��#�$v}�l@���K:7y���{�Bz�%c���$�:�u�L<kie��:���c#�#�'����1�:<F!��M�1�=ز�<P��z{��%�Ŕ&�a�,�Q#أ�$q�It#�g�I1��fG=�:U/r��'fK,��t�x�I$�"jh���<R#���nidu ڂzA�JKOxMG�a'�K��M��D���F	%tMH����t�Yd'R�#Ol`�cK<�,�&�����4�`��4� x����v �1nxo�y8oz�2u���2�N������{�����n庖Q.t�N�5�N���z���Ǎ�K���"w���N�YW���6�#��v��'�'n9-�m2�K�N��'��ARKQZ^F%d"�"N�����
ز{�K�A�$�R%�5���kŘPԙ�I;��A��̄Hؓ�� �b&#�X�+M/�����Vw����b5����L��B]�)F���v���4�G��,���:��:ZAt�i���M�w�:vCǓ�;�Y���f�Y)�'D�J�(�t�äW
�@���-10�����3��(�����RA<Oq:WI�!�1L���x�z#��z8�$���S7N�,�(�zBc�ZA����%�J�VD	xV	�#&�ǣ���hZ%(��Z���t�J���Vn��ힳ�{�����mm��kZ�ԯ�L�H����$#�5 �&���Ζ�i"#D1 ��7������#'�ܳHK7���&q4�RM<`�c�:'N��8��D�S,x�G7�Q�ǐD���ٸA�-4���GG�<""f�5 �>#�ٓ�&X��yf�h�J$���@�Q��h��%���I�<�c$�/�@��d,D�MI:8@��#���:<�4N؉Z&�{�hE��W�D�4�Q�KM<Q�DQ��Ν�BX��O%;�	DL�Ν:<��� ��ΏK�4F��D��"Oh���D��@��(舙"X�C���B�� �Gy%{ēi	I���= y�����	J)ɢB&�gR�:JL{��@�¸$���&��a�,��i&��i^�Yw�R"n	��BIign"�����#��Y	bN		�2x|A� ��I�:�$�""wN٧��P�m:2A<��(HD�"h�������#q�3�P�b���ĴM6�P�G����'k��*Ȳ�S4΅���x�JD�ƈ ����-/0�i(�$aF��t�t �J.�h���<����b���X�8�>l�<$��(HK(�,���E��aDIbYV"v�-�s��q ���t���簘aX��"d�#�{2#�"V&��2J ��,��H�(�H M#�#QBh��;@�J"]"F�$�Y�1�O�Y$�%��У��}���ò@��=��b&�b��<$���H�J�,�I D�aG��D�"h����e�DK-����:&�@�W�"�N���JA��"{�&؝h���(�D�3�<��(��"x�DdK:x<�"%��&	Yr&��AR@�DD�lDO%:Y"@�D��a	�&�M�D$��#�|x�x�)0蛢ixP�%D�h�w��+�s���S��BOtK�zg�;��9�/��t��� �	��:A\��@�^�L�,M��OYx@\��3�&'Q�4K4�$��:j0B��5[L���m����ԕC�Y|,��:w�� Cy���Q$ j:ODM14��ؕ� ��%"M��{��,O%�T�ky�u굫h�uϞo�JaiL�A.��#&'y�\i�Et�sd2���9���#�p�rn��ON��OD����h������I��%	��y1i|�yFIzD�D��-�d�(�O'��%���g��)0��|�!1�=G�n;G�;��R��I0�)5)���O�x��c�I�R��LLM�9|�O0�K��/��jl	�d�!'�QI},�&�3�e�DQd�G��i��Y����$QP�_n�!;g3��- ˃��v�ۣ��M3��bfZY�:�1eYԲ�Ʀ��G/��{�"BWD�	����SǺQ�:�4g>*���`�b!�q(�RW�rD�$L�7���Y�ɇ���0�:"z�ɢm�h�$	(��D��<���K<I�	c��b'OD�%��<M(�B%%ȉ�QǑxþ�DL�D}	G���e��bK��tx� x��肴H:��Ȃ�B"'�"Śid�G/����v���D��L#�,x��EB$�"%��x� K� y��xOD"Wa6a4��A�!:3)�(��ib\�#as��jvĂX���p���a�X�,�-.bD�#��FbKر1�:<L��f��"a��x�"<P�$��`�X�ŉf1�M���=��c�#��Gb�l&1g��\� ���/{���v!�n�0�(�H�;I�7S�2��DDK�:�,�$O%��	�l�X�A&E�1&	�`�YX�;eDX�,��<�Ɖ��Y�0�@�'L�,{	���[��yE�A��L�,AYa��t�&�L�����	��u����^N�%�&�Q�!W�w��D����L�;�/b�(��	و�N���7	9��� �L=�.+z��1��y����+��?5?�a�!^�V�
;?����?�Ǔ��~�f�#��$�D��vI��_�Q,6��9�^�p��1����g�����P��"�ăI(�	/^m�{� �i��8k���g)��p�s�A�J�m��ji;��A*!��Oni��Nњ^�������4�{vD�HZ�
�!1�/�vi
Rb �N���!��h�-�}������:"��[Y�M(#�8>#yN��f�шBf�%�a���1g�O:�����g&J�htG�Qg��}��^qǜ����������� ��q�D��[����B�c<3�+�1e>H3��K�7���2S�ǆt�s��Q�#��(�oI�cg��JR^2w���!æ���g�L�	�$�����՝0�H,E4D�'��d(�8S�5����> �#ǆA����
Ӽ�f��<sD҈���K$K��Q1�ExH�FCN�|�w��h�1c������+^�V�
i]�<�˶�D4Ӥ4�t���|0�:S�����n=t�:i�B��ҟ6|'L,N������p�c��2�&\�E�F�8h#FS��M]��@�3��j��e4e�5g8�L�i��y���ө��KG�p�%R�������n@��#�)��#��x|3�:"�G��\M4Ӣ4��M����<x�6곜��k�g������ㆻ�Z$��>)�>44c�28A�������xfb��+泆2�g�!�Ĺ�h�Rf�f����2G�P�ct4)H!��w~�R�4��7�dg�3�����"��8樂xA6!�v�렄C�(�ǎ{�γ:t!D!^��iciD2jļ�#)C����M(�A�=�n���P�Ki�I�9��7���:�,�����#�� �������4�)�'��wqAa�T��?�5�k%�q����E::ל=����Cw�����nع�>�9��� �3�����{�����z�oE)۴՝���ܕ�vc�{|�'�&������k�5�YK�z�f��W��R�x����φ�M�y���dd�Ezs�����L���|C��3�[��~���>-�.�ɮ����C�Cn.�I�dӜg��7���̫�D?2����W�ҭqz�u����:s������B/�T��SOs��H�r����dW��������|���M�����~o���\|5�5U����uw�������a<ͰַR,����������\�zo�׻��z����C�ȗ(<\닂��]������q� �s'|Ti1���������
6��?~�|�d�/��3��m��=,�����D����y�-�^���e��rW;acKG�����͒�.o�`-L⿋��y��B�{x��k�}OQ�w�V�^q]ykώ^��&(���!�B�ة����c�w��v�8\Y�i��<t�Tx�-��!��jn�F�حx���v�d�d�rC��!�h��LI��9����$).������y���b�5G�xEo0�){���6��Ӝ��E�E{ķ�z#Ws���g
�9�g|w�������ONr��)>�v��.�{����U���P��?C����Q&���|ͣ�H�tss��+�t*���G�9��J������u�s�tG#-�{ӭtz��؉����3�^�ֈ&��
/t�"�*�\�|l��3�'r���;8�Ц�t��:N���"����S��E�kNp��9��P���{㇯
o��i=Q�q<vX�O���ؓt��+�#d98p��9����G�7��	���YB^���🇍�^f�A�{㆗��gٿ�4��Ǜ(�4�D�rQ��K�Cl��L����7���,@���П3�8���7���	���p�:����)���)4��;�mq����w�;2���*��;)�][���H�t��+͍�1��v8M�OVԯҦ��f��e�LO�=|jz�q��P�;M?!��p�B����8t��v�"�G�BX�e���)���4�{�9�+��z]衩�q��JY��}!޲tf�1���p_/����4��6Bg�M��e���¬6<�!+l�J!�)&h���wD/3����:*�}�Q�,^rj-᧹�D��L�k!�g�hQ9�Vh2X���M��6R��<%Ot�O>�;�u��g
ɨ�饗#�yӇe:lD��;ћ�sQ�5ʬ�P[�6S�=��C�C㱚{�w1Q�#��Czn�89P�7��8p9)�{����$ExvDA�z�8R�Az���q��b�
�kȽ�:E{G�5����y��7w?p|��u	�G���zM�p�!9�N!��V�~����ޕ��Ok9φ�9ӿ�����Yӟ/בt����Y�S�1�1h�_;ËNE�Unno�^�N�C�5�~�ޭ����7��p�g��i��ZwiĎg�8J4�[�&�j��h�����S�C#�r{�Z#�۞D��ܢ�\�W�+�]9��qb��S���i�Мya�U':iγ�M�;���H���9��J�̜��xN�ŝ��2��A�x��y�g7����K2�E�}G�5��v�����s�i49N�"d�_�k�.�Zm_�,�ߟ��y��������-�1��^c��{G�Ni7)�]��9M��|c6�orЯ8�O��U�]cgQ�G���N�P������G�wϐ�9;�~��m��êA��|wtݧR#���Ǭ��7��+�Y��Q�|C��̨B���'?q�0������-�?��4]:�%+W��I�P�)�
�wCH�n��"s'zEs�|��G;���ΐ���>Vs�~9�_!�$9���Nm5�G#�cӋH��c�{xs�/4�
��nsxq��-&����ï�h���>����c,�q^.--�,ClG�w�͇=�_�P�B;��n�f�ud۬��m��%3�V�cf��&���n�x����E�q�sl�Q����ޏz?��W���㟖ш��ءg�jF��ez'��g<��=�;�R������ß�=g++g��Q�̈́�d5�J7�_����x��e������O5p�G8�9���8si�H|�ZD�w����c�S����k�w��=�p\Ep��5��z�b(�^9�n'�4O�����5��=Vz���쪣��ݎ��s�[ѝ6�yN���n��:^ު��摲^��oa-9zE=��9�-���}��*�{�s��b������}�Y㜅��s�4�s��=?�nhńӾ�u����߇�$�!��4���?��:�;.$s`��s�9��]#�9|2��F�3�;�:3�iC�V��v󎩢V�#�G��9խ�)�P�j��+�[M<�M�8����<0�������
g��	�T��C�xL�ߗ�~��M���������i����?��	#��'��[��Z9�������j]-m�������ouvyo��mpK����V�8Ln^z.��z{�]��>l�[g���a���oX�7�힫{�����_l_>s���M���w�ME��"���FFf�Y���6K.�}��r�����8��l���m���u�׵��MJK]������V���F�H������>i���g9��6g*��Kt���㛮8��.*7d^9�:��b���|�;��%�;�ظw�����#A"�y �ؗ�j���|w�K�vN�_�j��CK�K~�g-�(�C��ױ�BeH�f�{�.����{3��i(��$�b;ˬ�l�}��B�'W��۽�^�I:T�By�4Ѵ��Vqiw{�]:�d�A�G,����K��MW��e��S�-��;����`�N	�x���9zҒN[9����3u{��j���ڸ��i�qq���^���S����O�Qz��w��o'V���_�����y_8�W����o3��{[I{���T�|����o,�.z��ڵ�S\���*n�����I$9!�o��+�y�s������=�MzbuʧW;��qʭ�=��Tx�{ؽ6{��K�^o��G\������8�;����ooJs����W����s�r�}�F����;�=�U�GJ.�z◔�i�8��Q���]R�oy䞞=����B��%�M�﷯���^���W�{�4Vs�{f��ޡ��x]��x���|�ӏ����uo;6���!�ȫd^`�#��HZ��B�e�-�Rs�q:���ꜭl"�TV�?5�p��Dܞ$�aC�-Ԩ�%d^�U�E^�#w}���C�*�.&���o]pi��{ow����<����=۝Z����93��7&��J4���J�"���T�:��N�E�8�����[٫��>��QH�����[S=5p\�cW�l�^�n�t]�$:�s�ݮ(-�������j�krN���s�{�l��YΪ#֡?n�r&%X�]K���LD�͙5$��w�~y%��T!R���{Կ���٣o��*o�5�/��ٿ/���K�D������m��{e�oܫ�t��'Ӿ���7�Q�M���z���nb#7;���Սr#;SگA1�������U</$��q.wM;��y��s�=��]ݳ���Ǯ!����F9ZVgzw�5�_�������VN��8�V�T�v2��K<۟�=�{��3-���7�Ė=m9��#z��O/�?������z��=E{���-]�P��M�ͻ�s���Y�ԓJ�ry������&���;͗�/��y�,�>�z��vM�a���Q�/w}�zu)䋱���u]�����o�v��U=����2+�Y�=���n�n=����"ShI�R_n�j�vo>y�u��ݭqk^F�-�ݫ��ݧ'{�[��ݜV-�m�~����l:?j�bi3����v�}*��+���i]u+�J�ervw�Ye�s{Tޑ�y��k�����w�
��T:��{R{M�|�]���=�~��_ci��nz;�������7>�պ����G�J�?����v�~��%@��׫����'�.�Tݿ�����{�ȏ�㕴�B�q�sr�7�yu��z6ׯW7��҂�6V/s�����|Y����K���\[[6����w*57�����wW;�s��,��8vU�oz����R�q]�R��#�]H�N���,߿:q?gc^���r��J��H��i(�e/�[�������g���4����ߥ�ǉ:��]��E�w����b�'��k�B��^;9�^��;�><v�����S��
c$�������έ��K}�Bշ��ʣo��rp}�u�4��̕]EN�~^�:������߸P��1I{;~���s�F��x�fH�����|�%��Ưo����w�5����ە�3���&�Ѳ�-�lغ�8+��$JN�i�2NM��� �r��|��x�z<�i�m7dx�����R[R�!#��ՉԊH�]ZQ.7Nj��`�[+b7v�-��������lղu����iB)������,�Go����IWS�W"�����K��2�:�N�]/�k׎'�^�J:�U��#V�лuGb�]���ʣwfߦ�N9�v��}�ti��y�+O+z�Q��j,|��"���ٓ���
.����#ic�,�lnNX}^�s\��m�9���Ա<�&¶�e���w�RL}D�H�I>[5�#R#iȔ�H��4�5{���G#����qƞ�+h�DWͪ=�[�c�̈�p�6��d��֫�_KN2-hR�;J��Z,��dG�Աk��F��o-�9�>9�^R�fأ��'��jq[Ŵ�5�ܻ~�D��V%%�������R-u��)�e��c�%%��$�R&�wV����Z;6X�"\�{�9ȵIc�7�IĶê7U�$I��6��w����>�R>+UYeM֋D�#Q�奅{�f��Z��ZI;����|��6�6�[ETpM�I��vȒ�_����H��Fl��	)S=4���ܓ,��e�n�N���zs=P�����w�/��W���W���'��s?'@S��'���~�������'*��(�� ��[O���_������~���/�~�1;�Ώ���`�9?6��w��UUaUWVUuUU^����U\EUm_*�UmU�V�|���UUŅU]E|����ھUZU�VUZU��ª�����*�j�Wʫh���
ʫ��UiVU���ʰ����U[UeU��UY�����%��4T�؊�6�t5��f�\Z�K`�E)�4mEF�h�4Z��Z�mfX����9�ϫ1[W��⯕V�|����U�U�YUeU��UU�U�YUU�ꪶ��YUiWʫj�U\XUUXUU��ҬھUZU�_*��*��*��ªҬ��UqUUUqz���O�UeU�Um_*�j�Wʫ%��� "5Ilm��lUe#X�%jJ�,���f�&��V�5���r�Tk&�ɶ�lU�����6�V�BD�ad�u�o=�ʪ���V�eUiVUV�eUU�U�|�UU�UUu�UUEUWXUV��Ҭ���ү�V�UUQUU�Uqz��*ʯ�V�ꪸ��ھUeU�z��+�UqY�ڧʪ��UUTUUu���{�w�\�����HȲH��b4ks����H�L𭹕�BkF�X�]-r[�5��L��s
��>��~u�UWXUUu�UWXUUu�UUEU\^����ª��*��ª��������*�j�U�V�ꪸ�UUŅU]EUm_*�*ʫ*�,+*�0����U�YU��*�33�*��*��ª�����£�r��Dp"9�M%&ކ��KL"��T��♨�9�h��FDd@�H�V��\@�!"��F�Q ��R��	$���7�	;�E�5F�n5�4m�G\�[�*��\��Q�Z.6�cU�^?S�������@dI?�����+�@�#O�?B?B�������`����<Y DI:X��%DN��B&�"h�P�I�C� �"t�	��$����0LK0ML4MN��h��i��D��DDD�D�
:"xDJI�	bP�$�,��"H�b"Y�Y�A:"%��h��:�\qm���i+B҅�� ��$�$	gD�$O4�L0�DJ A(D��E�"h��aBQ'DA
YՖY�G�W�����qܛSŸ�O����H]�AFt��HS�ٲi�.������'�Dy�8A� ���(�a��(�p�DxGN��ކ�B���!�b(SN<E�\)�^iIĆC$2X$t�2��LC���
A�ҵ�Z&k�&B,�Х|!�.f�+qLx��l�jߍ9t�m!�����Y(s����vmd>1/|�����V܇
t�������\AYd�B��xB� <F6ٹ2��"b�Ȉ:B�D��ЬE鬀��U�F�#�)ii~����1&������ 4�3��5B�
�mA�A)�����Դ�B��ȑT�c�$z9N|NeXB���8hlW�A
k֊]\9�s���{���q��j�,�Z)D\D�tf� �Ǝ	jON�Sj����,E~��4��I�D�p�鈻��=�p�>�v��|��}�o_�I����<��섖��J���p�_o$#�E��=��I�v�{]G5Iʍ���ّ�����s������淦�&����_n��i��aji�%g9�_y��_���N��죈v"
�y7�;}7�rji�+������q�H챖�[}�1k}�F]
�J�D�d��娎�Qc�OV�^��T�'�D��ʛ�q��vm��溕�$V��B%��?�Y�q���j�m_��w�w_�߱aUWQU�����p�^���,*��*�33�9ß+�W~ŅU]EVff~9Áϕ꫿bª���33?p�p�� D�D�KD҄�<i�p���x
pq��4)�0��4Ӥ�Kӵ�Ac�U"d; �2����o(�7rR�J�u�<���\6���a&�4d��/�9x���5���Ԓ�f�1q���9�n⪱�h�+gjI%L1�~ut�?�g+6�����:r�W'��8QȢ�� �c���1�me�i�N��9�d��.��,>=�2w�6K�x�n�ٍ;�SM�2Ioz��A�L�8�`ed�v�,l{��x=v�x��7�a�L�9��ƞ�8SEJ8n$uC�i0I�&�HL7In��c����|���!�X?�����lI5]�[J�Hڟ��5���oq��n%����nI:#�:C�:|�V��j[�-*Ru�<�8Bi����Z{���o��$�9��������i�������6p�q���c֜4��Ls;�lh�9�g	,i�!7/���޻$��f]�qÓ�p�m���B:f��I�#�޺c9Y�?�p��G�u�"�e+>f�Pm��Z��Nޤ��rOw}�l�9��ɼ]Uʻ*M49�܎=�x������R�� ܑ�sz�F4 �Cki�ژ�V��j[�-*4�:������G&�b�}�{�ڒI!>�(4'�>����x�q���=Z]�އ,Z=]����o�\����&S>�Gy��g��H�޸v��s|f�ԅ��N�9i� ܦ���_����PH�,U��4��q��܃u4&,�s81�J(���>�D�ÇN4p��D-�^����F��.��=v�#vC��;� I�Z��Ys�ѧ��m�
쪯1�림8;�m�S�gD�ϵ��JP�u�����ֵ-Ku�JCΥ*k�\!�[�y�ΫF�I$�e�x��C��d���i��>��^�ݞ�HC'e��%#!G����K��[6Ӄ.t��4��4�9cA��!�7���	[�$����\����8e��׵�ᗦʅJ%�-b��݄��&���p�m�l� ��^8j�6k�f�����0S��xZ:p��;u������t�P�m<�ͼź��KR�yiR���x���#�s�m���0Tb,�D�r��4DИ��uM݈z��Q�J�J�>����3�"�m��"6i�%�CF�%H�uRA�=`�H~V�&N!T�!41����0o^yuys���:u�9�s24���n��Z.�Q�/h�u�7\UD�����֣��&�@���TRjI$�E	!j%i��Rز6F�4�$�.w�^�1�Z|֙�AN��4G<�CUG�]�g�|k>�#-�Y<w����V��"��ֳ�3�&|tB_b	!8�c�%���i4[�du���A��tvi�f��z�7A�Q�2����?b�ZT!�H\�2�!��c�4��.�GR5��jj6�X����ܐp�����x�f��nx7��ے�K7�g�4���-��im��ukZ����ҥ!乥)�i�9����H���\��ӗ6����p��2[ڪ�Lf^S�d�N�BK0��Ipܨ���#׎B�Y�y`a�nR�0�N�s�㯚yΑ�Fe���m�
=�<N�e�
���
��9�r���%M*(�HLI}�?^�ɸ��q��E�u��5���o����.���\:pi�h<�'�8\�7s�qb�k,(��"���0�KD�0� �H0�(��I;�{ͽ&�ޤ�HG����)�T�N� j`����>(�Ѯ��������5ª�����u��Ɲ8�c�������C��N�
܋.Kh�u����AIχo
�$���WNӇ��\��I����	+�$M.��=t��9���1}��ؒ��\DEL��c��ǋ.JY�����߰z&�P��d�{5��9���|x�uM׻��cr(:��=kO]'
�CSJmKc�ZԵ-疅),�p��]M�I$����.���ǞOUx�U����Z�N�'�5U�o�2I׺i΂Bl1׶0�;L/�E6$�<Hu��6�ID��#>hŎ����;�)+ʹZ���?� t�S<{<~>[�α%r��4M��ѱ&�x7_n<��Y�G	���«d��2�rhz��nBS����<m��[�4W*]�=p�@���u΍�/Hp,�6�N4��Z�Z֥�o-E(GMb> 2d�}��G�W��=����4$XR)%�ґ�n�������A����5�B4�ʴ��]����X>Jr�H̓��H��D-4�b�CM%�<Cd��S$&�I^��&,��HB�$~C<s�P��ڟ�]���:Ɵģ�6�D���%k&6�ݢ��ɪ��s���6�;I$s!��eU��ƱF�qH��u.���1�M9a�����I�hr�`��j�\ŗ�NX��:>���]7�Q��}�����V�8^�[�7̕����MI�pNQZ��N�1 Pq���v�4=^k9)���4�&$���h�[��d'Xdԇ�}o��x�����a܄"1�H2������ܩl�A��ʊ�VA�q��s�;v�;��m�6��q�����.i�ē�za���Hx�
R��ֵ-Kyj)HyWR2��dr��RI$3���s�s�I�̳�P��*:l:�g�٭��v}��$����*�I+�^�bJ=�T!$������4�?���k"��f~���D)N��^�S�M6ۻ1	#	��f�'�q�Xrߞn��B�pd��ڝ������@���i�>ϋ����0��ULv��B�IW�O\�7�6�����r�����h(o��H��F�~a#(tQOHY�)Ŀ#�q�����hJ0��1��1ļ��1����6�5�Ɠ��'�N!H�b-�ZX��ws��e����Ļ��K�x�wM�N̻��rw/w.x�wW7���bF!�%�u��H�bĭGԆ-,ZTı�"ыN!H�SlK�&�Hy�5(�b1�5�c��b1�F<��F#�Jv���Fш�}���bӈ��"_�:x'�GD�+��U� ��>'�=,}>�N���t�>��:I�����S��&шb1Eb%�'��m��KL#lN�Ĵ�S��w2w=ܹܓ��rK�Q�S�x���<F��e!�eb8�#h��h�Z)�5��[�S��'�'�ORƱıF#�"��'�qF!L!��LD#��"C�CO��^~{�4ӊu�����Oͥ��_SJ��.ڒ�Un)2���F�7:�,Θa�:QҎ�DY�G�De?��h�X�c/�7�녅><z�z���K�z����`z[� ��H�`2X�O��.*�	�'��殽y__n:���x��_{ɜ��3���y�~&=���o}y�j���{�}�w�y�:�s�ٿ٨���2�~���fffec.�Z֭��UZ��������fec33Z֯>>*��UU�ۻ������ff��e}�UV���;wswww~����kZ������8ҚSjcZ֥�o-E1iS_L(��Ǉx�����_z�t��cl����#LFp�L�#qy�N�M�e:h7R*�`x@��mU�p�tq�[e�)��'*��`��ڞ�@��F��p�U�3>�Y��lN��B���`�kT�@��P�	��r{��&	�l\T�;��zoڷ��|e}��{��ؙ_�_�V����{K���Sh�d%� �`rƆ�i l�J���-���h
 t�%	�<��v��e0�A�ψ�d��σ����ӗ�׷!�f��I��e�vz�4h�VX��3���#�Ν6 l�F�oз�d��4�
O�; 򔈝>�}��5��m
q�4���:�<���R��%�}�,���GZ�f��"����<�;�(�g���<�Wiw�	m�)��.�3���E8�P����8{���N5�A�9}7������L��؉��Aa7�W8�6 �h!��B�w�)�Kp}�l��� m�2�lDd�Uc��>��@�׸���տr���� kd�C�D�V������G���g�(:DÇ�f�JDt�ڻ���i�0��.�5���'ʻɇ�1��O
�O9u�L`}O����5�N�Xx�y�9i9σ�0�b�q�_�=#IACL��Ɩ��[��ZԵ-娥1**���dek���H�a!���PK�-�6jx*T��=Z\�a��R�5�,bBx��nYo�9��cJX9,jX����Jva�-o�+>���",�o�u�s��Ϝ.�
�}�p��:w�˩Ԭ�%YbN�1�8��8�R��r�28�t�"����,v��s0ɑ��MAD�䌙d�7�#*�Xa���E!�w��}���\p y���AP0l<̙�Y�q+�Z�d��F�V8qF�&r;l�y�l��Q��U�:d�X7�~((������9S�i�[�`0 q�����[4��x��g���0�4��[�0vI<T�p�`B�$�17�c39����}���þ0��S
:��<�X|������0�`d���e�t�2o3�b�::��a�u�H��x�wqāilx@�g�GN�,�!A*�a�Y��i�y�f%���"b���=���k���Q�8y��%b��r���D�̐��қ[��ZԵ-娥1*uˉy%8�c�ն���G�DD��F��5�y����CϑQQh(���w�8��$L��Xi��Hl��X���f���{~mp@�&�?4>aߍ��R�F\����[:�i��#c�00��l!�	���$aз��9h }��*��#�u�"���{�J��$&!�n!��2�Ah��yV~{�fg�8�~h0�11ym:���I%���c���nC�	i����Z�4�9:�`D��ߙ����4lݚ�V�ڢ]12��L����@4F�6&\:��=Yla�p�xZ���Ń��}��5Ǎ58�l�[O� lixA@�A���EBA=�4�S@Y�k��ۀ����D�A�E4A�Y�2Y�O)��:��KZ�Z�Rc�p�|y!�q�og{�'�J���PQ���a�4�Y�jn�(�*�9�x@Ʉ��no���S)<`�ǍPJ��-o�9bfA��D�p�O�}�*�~~C�TU6:a6�:��2�4S頢K$���9{n�*謅Q�i=�&T� Y�����,���D��$�1�M��Qg�lh ��c�\|��� :�lOa���0��XcX�ߚ�*VGZRC�l�Y�u�!��{�s뫽g	g*��{�9'��bY��13��㤓�%��9�,�y��t�el�ye2��L�8�R�0�3Ɔ0�A9��+}�<@�C�pǑK"��mSLJ���N��$�n'� Qr��]`�Ƅ�G�U��	���)��WK<��8Қc�8�'�:��KZ�Z�Rc�r	�w�ږ�ٸ��Z���}��QQQPH�D�W��.��	�`B;a��Bް�UR��M@>��ۄ�t�[ ����)O���[���'-$>`ָ���bm�D �a��j'��It��3H���q�H[F�'L�"&ǔ��������g��c��ڰ2��l$M������.(����*S��M�6s�ju���-�6l�j��0��7�|�N��9m5͒���3M���%&`d��	p�Q(����L�$	h(���qI6B���dA�S�>�%])�&��[vL4>!p$2`��h������	D}�%�8!li��O�6�16�0ı�Pv�p���p�hւ�X���n�P����E4D�Eǉ�-��c��!�� |��& �ST�P�'�ap	�F�e�
������1�����ZԵ�娥!�:ѪJ�L?q�)Ϻn55#�O#���n̕����
���H^8���n,C۟��FYFR��q� �x�_JAj_kr�

�%��
Ldn�|�ӄYRƒi�ah�	��H�lHL�����lǬB�Ʒg�<X�v��8�նAT!&��ݚ��K�d.OMb***	,ܭ컝5��i��K�5��ב��9�0�,7>�i��bA
�C��㌤����F[]�:Y%0d���c�{�I��(�u�H����VN���"Y��\3�*C��H�O�
M4�H���� M�e�LF̄ղݰ�|Q>�SE��7�7�_l��W��n�<B��Z.<b{�}��Zϋ|�0E�؆��m\P��BPq�idd>`��!De i��$CA�V��Ӳ����G����%��q��8 ��������Ѭ�7��\�9�׆�$���/eD�i=�HT�0���P|@�h�V����5U�J�0�^*MjI8f(�R�,v�1�(��xݏe�JWӻ:I׎�Gn��&���@d0ݓD(�4�kM�)Ç4q���uƟ�S��έkRַ��!�����N���1b��!$��4���~�}x�=������pk��'%��6�ϵͼ�N\jT�<@��n�4Y�D�ʫ���$��[l���(v�WD�TcXyQɦi�yݲ�(����0a�4 p�������p�ه��b�:7'|�[zG+���]��\�!i��ؕ�3c#�]��Y�m�	��^�����)�m��$f�B�u��7N�i�IA){��n�-��s`ܕ��#a�5�h>�$0K��6�7��fYn4H$��rc�Y��5�S�r9td����ڠ� ��M��m�4�G���Ta*�Ü����sʀ�1����=y��}���yƔ����ZԵ�娥!�)�m���n�z�M�G�EEX�HP:I�J�4a��H�	�Ε4v����D	 �~h��X�f�SͶ2��-��= JΞT���JӁ�}��,\�8q��Ǎ��:����ӅP��f�)�@�;�l�x�������N�P�MX�ap��O����afl���ʂT�J�t�j���y�4�������`}�8z31��Kу�Ln��	Xt�`�V=fN4����%1:�4d�ϛѦg9rm������1����<I
���}o�T�^��}�V=Y������m<PA�D�ʛ^��SJ��hȞ4��������3_{Y�ٍ{|� x�:�q��~~q��խjZ���R���jzH����Ms��W��>�c�@�y�WR�����*��t��!$��4մ n+��pC���D���5���a�r��zl��K,lE3)�#dҊ�����Eu&YiK�����`x��i�f�4k��
 ���#������#��=�m�����3e`1D'�������p���5�6�ߪ��Qa˚
�{yFd}�;��p������90S(& �����ǿ�^1����F$�]�%8qN�̹��>��� ۡ�c����~! k��X�\�َ�?5r���2X۝|�q����a��^]�)����Ѕ�I4�0��8QOY���Jv���.�h����F�F51��'�N#�9���I�'�3Q��u���1���KK�OP�u;��.�wJ��.]��I܄1BP�<�����:F!�11,C�O؇�kJ����R>�%�K�-8����ĭ��&X�B�NؘF#�18�u8�#��cɔB��"P�bq�#�c�b��>�u��O�c�u����6�ChJ1��1�5�b1b�Ħ؞�Q�cLi����S�M�шc����bz��GF��'L��xN��],�맋�'rN�ľ�w$_k�Ԯ�'I],k��:JI�p�!���h��#h��-6��)I�b-��S��b1�q��u��m��F"ш�'|�ܽ]��/3��N黥�K�<HO��\=g)�Y�/Ś���i2=S1S�$"��F�a�����)�x�9����\�����rD�t��:Y$+��:?�|s�Jh�n���B�����ӂ6:0E-��2������F1�č!�sj�Ƴ�B�NeIH"���܏Q]i�f�2݇�->+�cr8�ܒ�ǔ�Mʞ1T������N���X]������h�qj���m5[!T�k4�����(ɒ�c���O-�p�*
h��s���A��IS�r�B�B���G���Y��4]�w8s��v���,�4�����9�^vT�;Ӈ��2Å)A��V{zG��>���m��Y�qlM�WH��A腭S(���G	f&(�!Ѹ���^�PL��"�	��= �"kq�����[�&��z[�e�['G58BJ��dR��FT���I`�A�v1eԛ�yb��~7C�8x�t��F4���M �ԙ�p�x� ��p��_n�Ȧ��qAo��.kX֡�0B�Nz�-v���kK��������v4��'��"K�-ם��N%�$l�Xʡ�A�'"My7��͜M ����Є�$K{�Nǐ�6�p�\���"�ğ{z��k9Ώ#����Y�,���6B��ԑ[�xʕ�[E�g?�����*Ww��^�����O��%Cڶ������Ϧ��<�v�����w7o�U���'w���)_�g�t����w����w��&�9�rG���TQ
/rh�v8�\iC�wT�����"�oYŪjS�V��D�l�ĸ���5Ԝ��Ūc�dU�/'1��rsy�*{���U+�Z|����X��	P��J�J1�iqUjPLE�m�Y�*��H���(�$�MYĜ�TIl���X܍+9��	s����^*6����h�ܟ��ߊW������T��W�ݝ���U��¿T��\����߾�_*��+�L���wwv�~�U|��������|m�!N4����X��k[�QJC�m}����b^�p�>Ks��L��n���2nL���GjѫD�!,�� ��8*&��׭�a��^=!N�׼�:ߞդ&���5�Nm���9,��o7Gl ���Ő�Y7z�*L�籌c�H�� �#C��C��B!ux�V/)X��2p; ~4��ٮ��c�����|@�7ƾe�
�8h���S����a�l��z�׍�v�aN*��>pX��Pm������T�c:0�Ge|��0r	��s�._���N���n��h3�k����t�ä�&z�i���8P�qA�qA��w����Ju�̓���#}m�� �Ӎ���p<� d!�>A6d8��:����shr�Oq�m�
����������~_���n�)���O�;5��r��b�$�K�����Jo����%x���n\���
3���~�2�(��'��Q*5P)�_l)�,6)ĸ�Kio�?1�-jZ���R���)�SKc��;ͱ�_DD#�H�$ї�<s�����Ӛ�y�q�c�H��t ���s�M]K�C� ԡ������ӆ<v�/����x��d�(H�$�Γ��Q�MW404�;��\	��$�4�}��.�[^e��  p�J�dena���p���/;��FL)�ǫA��o�X���,��t�����$B�e��L�vx����D ��T2�yj�rV���u�O7��>
����n��~s65���0��)���X3�E��ϙ�n�Bt�p,�e���f-<zh���@� ������H��._���➷N���F�i/8��O)�1�-jZ���R��K|#�y����k��=��}o�����M4�@�pFy��e2���I��s9tA�<x��&�E���i��ӆ�BH`q�Ƕ��B5Uxc/Lj��CDY%�8�o,ɗ�.cnFϳ����_�c��7)q�E��!gh�i aeųH궤��2)�$�Ǯ�<|O��d��lo(��9$h��w��~z����C"}�m��m�:��05Ɓg��)�Qb�/ck�g���Ph�M�����oϛ�s�ę0!�>�p;���ːӆq��3A��9���������^������ϸ�����`�Q �(�Mz:YGm�-�??:ŭKZ�Z�R28�C���٦��T�M4�ADnd��ˬ&||���47�o��)���AOL�h���g;�����C��3X&��g����ɓTBf�MB�4j�=[G�B\I2<>t??�g�[�և��x�4zR��`�9�}�_����}$ӊt�y�d<@�@�8t-��K�ÿ8M��ǮC2@���<���G0������:x�v�v�d
`y��:�&�Ӯe9�J6t�7f�÷4���J���i�b
xҒIBg�d3�f����qRJxp�N�$���ä09�a��%z{�H�q���gF� h���$C{"Q��^wz�!������Z~q�4�8����-kyj)Hy֝Q��Kq	i:#քڃ��63��Jl,�����V�f�6��0�M%�qRW[x��O,h̥W<]è�֙���gS�IEG,aadE�E�1y#�ѐٳt�� �3�5�a�Re����ʋ2!�$�����)m�VҌ��(se�!$��ڒBZ�[n��*X��GT>�D�M4�@��3�CD�\�k���UR���D�J��!y����,3rݥ0pa�*�6�%�t���<ɬ-����g#��Ņ�# �d�����͘B��� p�"�u��@��"��Ps*�C�i���4F5:��˷Xko[i���(�Q�@�١����:z�l��S�S#��=�㬠�N��FC,y邧���hxTC�Y�б{[�J� Y��t������J��P�տC:����<1���DiO�`�n��s�R`�=��i��C����>7�ƃ�`n3��;~x᳆7E�f��	��?Y$�h��l�2am��-��1jZ���R��>8N,�M�%E��g��64}	���\K�y��Q5�a��Ԑ�_�g����\c�04xl[��i�6��c��c��t��t��:�N2�*i�6���e.�@�Ѩ��f]V�y=$c��:>`��,��{\�檡+������Sz������j�Ǿ+F;nb��l��U��=|w����,(N9aJmģ&�{�t�3���/rL� �8l����Α��" ��d�<C��c��,�CM�.x��*�n�k9��|}&�<��R�㮸�^���,�0ct����P��4l��"d���*Xk�M�Fx��*644��iӡÎ�
��Zr�e�Bx�|�Ox��џ�wX
�YdֆD�0l�֋l�a��:`�F2|~u�Z�����<�Z[�~Ľ4&����7��'<�F�y���1��@;y�f�S�}n�fI���V�$�}zc��$
�0�V5gZ�m�7�O����h8@�J�);ӧ�W�_7�.�-�ũ�� [�9#�
"MPƺ�U:lt�؂�4gd�DE%&I1Z���.h*��-5�t�:���g.��g5�2���[.�e���l\{y����2=f4���n��-($K�D�+��aU��5Hv�B�*�VH��YQ-u�n�d��w��t�;���8��3�V�\/�`�)5���b�6z�$�r=��y��C��d0�0#�;�RW�(dn�j��G#�� tĥ��4�4��Y�9���_�����[o��-��1jZ���R���-Ω;B��|�����k�I��1�`$	P5]�֊�O��k�S].Uܧ�#a�����yװ��vpA��4����/?�/�v�e����Ju�P��%6���>r`~Y��8 w�O�?�r\��M0N�4�n�+��Иɍ�sr�ǁ�S<�������t�:2��lv��}W�@���O[�#��#G̍��z��b:+��i�d��n�����d;��2"d�'��V0A��f�=��$�9'v���F[v������Ǥ�nu�ۦ�*���/
z�p6@�q��6�eX�)�cGt�0l���d��y:QR�c��ۺi�<�i�m�4���:c�Ah�	E���^��F������t���2��������6������-kyj)Hy?6�i�֠�u=��:8%:�(#�p��-�j�˦�26��p�HR�B�F7B���p� JR�yi�m�{�X�pi$nBT�{��P��e<&�]'�:�d�Sˮ7�Ս(�ڣ�J5�9d�����i�0&���X@G��F̗��b�x�b�I��m4>uOy@��4Ӗ���':I�> `�.��$n�	�$��0c5L4����Cn+��> 2��u�=�'Ht���x��.j�`21��t��G�5P�R�񏎕uxpoM�\|í����ì'�c���6�@����Xq���~m��/:h�̄�g�>lj60K |b��1,�5�s��R�{�ߘ�l5�.x�΂�16۶M�lh~��-<�y�`�8����Ut��ڊ䬸�6<�E��䃒7L�%Ϙ�ঠ��9a������{t����M�d�����&�7{|9}O�i�A�C|`�F~q�α�Rַ������]�}W���z�ܼא�9�@�(H��<y�yw���q�ɷ�7�ɢLòFg$�6�cERU�Kl�3���\<�<�d�g�#r����RuQ����<pۇ8>+�9϶:���}xo�2g<���������u���%!�^�h3TU�@���]~j�|��BZl!����X]r��ۮk{��Q��LY��'��VU��c�Ñ��Zv�A8@������0�悶����M?s�Fc�e�gE9s��?/��Ga��\j���r�6tZ�>AK�[9c��I`������}O�IF�j?h8@�ղ�7R���#���g+z�S �6a�����YC_b̰�<���)� 'O��Wk�[~�$$�	y	��6߭�f�i�HO��Zw�!d,�	(���)(��?!�%�$���\F��D�K�Lc�b1I�b-�5(�!�����F#�M#1�Z1�����z��a��Ӱ��.�wz��ܒ�]˓�Q�1���%�q��ıG��y���4�%��ib�ŧhb-�Z�a+bqŵ�'��1�F1:bm�q�bV�y)D18�i2����1F#�'�-��:����F&��R���yG�����b|���b1E18E�L�N#lN؜CcX�E��&��Z<��q;�Ķ�CG�d���|a�æ3Bt�t��>�.�_h��7�rw.�SwG��O��}�-�#�-��O�'h���?1?�L��!��'LK�����F"шű�<�Q��gS�w�a.��'w����><RM��㎲����"������Gǉ��GH=�	
H���i�bV�����dzd�f�!dK"rw��8(���ܭ��������qu(CHQe���4X�3)���U�9���xAa@�@�⼈h������+��.��s����8�"����,`�Fܒ&���&7�G"$N4��D%E$b��H�c��!��X�Yq�22$WsY�-�����b#��G����̬w~66�p�����ܸ�kϱ����η'��U��'3j��M��<����#��v���_}��J��V���g�������U�ڽY��~�������UeU�z��L�&���n�����ҽY��~�A�A���6�8�:�-KZ�Z�R4���FS����r�^p͞vL�cUID|���5��ͅ��e�d�t���Kۤ!��:>i;[gd���R|��JC�%���0�,�/�JȜuT�sqg�	+mr��h�=so�{iْ�����D��V����=��ǻ]���4�
�9.�H�\n�r�ΝG3睯�2��C���	���	BB��jͷ�M�g�C)��>>�����4i�Q�V3�ƭ���9�iâ���:��Uo!��P�.��t�暍@�|z����]2
�����}m=z��u��M5�swYug-�(2x�	�������.;j��RcNX��u�4��t־�!����m���:��Xũk[�QJC��ikw����K������АѲ�"���H�n���Ӯ�'йy*�fN�GX��E�E�<r�)�&���b8��F�˹�����x�nZ���iM�#����c�K��?2{����5"_:"V�ZB)�?����r\���4;wn0��4C�8Ng���o�b��rk�4S�O��$��]9p�93(�kt�8��44���>@B?������Z8X��Īhv����t0��q�͇c�9,m����9�{��UF�N>!�nܧZ���g�0 x\��(p��d4IUn���ç�-h�OS�"���¶|SXJ3�@j�IZ]y��ڟ�c�c��娥!�ʭ���D:��k��R�>�k��d6"��p�M ލ��eg�&��m�4tՑ��DT(*G���!CO�D��dpd��8'4�Y*ը�-G7_0� ��sMF����lje�
����M�KI����}��zz�MCU3ThIͭF� ʬ��3P��.�ĕ(W������	y��\o,�"��ęm2��/'�<����	5�z��ﾢ�>�XCl$��)ç�4�|��L�L��kFB4%G�!���QG!��Tb��Ʋ!}�e�	�<�)r��1��֎@��h�T8�D;�F��49
��O9|jdo��x�Y��I�dri�a���pj�0>�G�SׁGv�X�8C����D�:7�*W3},4ǌB�n�D(�i��&C��yÇ�SƇ�7�´H�1tC���]>��&)q�#����䢦�%��C�SG���}�Ps>"�����<t�����p��
���%�-�2�﹐m����>��|h鴴��im8��_��x��M�88Cej䦈�T��Qt�H=�p$vA�^�w���:�wB���$����H���������Uc��,� ��|�<��^ԙ���
P$�Py�ny��QQQZ7�^�;;/����[�~t��p�p���S�����\���>|e��Ki�Qdh�|��!�WN���P|�o�8~;O�!�5�긣Q�JEĠ�N91,�
H��d��Lm4�29"$�䉐CI4����R	4'!��,���rFA��m1K�\T�ȗr�,#vo2�����< �y�~ا_t�ϲ\xW9�KM"1�Ԏ6ᮉ;��3����.s@�m�DpB�t�U[��|�ӊ�v2*Q&G��0G�u�a��D)���o�p�-�|IN~�C��K�!����^���(��J��Ca��ץ�RR�QA�C��{%��s3;�J8p�c��(6C%n�??vqۧq��-d�)�
s��q�|U�Iw[r<�N^��i����b�C�
�++E%5�Տ�ݘ�S��?0r��o'Ɯ�0~b�--%ךSKu���<�1lZ�Z�ǄtZS��h�u�iOMɼ�7�9��EEEhHY��++�ײ�P=���r[C˨nM�6Czv��;jU6�)�S�vߝ��1tB0vыV���=�I�ɡ���僇��!�<M���#4�KQ�cm�`�S�N��-��M�g�Y	rv��ө�a	)$,�ꮥ���:r�9�GqNE�V���۞���C��u��H}r�B������>�|�0(��i�A�NKq`��ӈ��~��H�#�v�Ɵ�X��X�*��L����I>r8y�t��i�~u�#�}bd���Ǎ<iŔ�i>��S����=����L�xC�-��8t��0l#���J��i��Y�Ã�<�IR�cKuN�1�1�b�><<#�ތz��V4�e���clTV��p���(�T�+������x�Ò�03֖�8"m�=rp����8�C�8c��>����;$�ێ�!q]�C(���n�ol�SćJD��͏*c�P��,dxĖI*����;��;�۱�A�}�W��
��n��;`�!gwɞ�J������%cr��;~�8t�'>ᑃ���&�����e�Ɂ�d��(�`�?��Yv�T.엀��b��p����)����sǹ�C�8c��j���X`p1�S��i��	�1��ڕ�}X�H����Xz��
�>tt��q3�ඒ���>r�0tYe6`�o?<����c�-娥!�<�r'��!sH���Ӂ��6Q�Q֛�]�8��i�"�Hh�㍤ĉ�$��YD��R_�l5A�I5Y1�/��$ڮ�rqw�������G,���-�עҌ��X&�5��ƿl6�W,���m��s��TTV������,QZ.����=m#V�F�Yw*����C	��1�<��3�N(v���)�y��F������$�ޱ�"d~�'FrBb�$1$��;>�h�!�Q�a�I|��!Lpۣ5�ᰣ�B����g\�0��f�Sd��x�2d0<C�Jz۰�>���7��؝`h���lp��ރ���?Z��M��Ϙ~y��x�ӟ�u���#}��j��\�[N�v�u%T!���u]�9h���V�Cuu\���bĸ��Ι�hdz���R��?D��[aD����hB��IA+ē�Z6I��	o�O�4�V��c�ο?<�1lb�Z�Riĸ�=j���:�>�?=��T			g&_<'9���_�QQZ(�?F��C,`h���(��OI'�$����/���U8p;,9L�
!�ҘԤ��!��Ң}�E4"Y#mܒI��[(�{_$��i���� �r���Y��L"���ʰ���z�<�Z�ΐ):�8C^��7�}��]37�ns��q���[*�q�~��]_�4�ٕ:aR���l���>���5/H��%��_�����rQG֤�	��S�Ӛh6��O:t;���D,`�����2Q�h�B�N�޶�;��h�6F�|ʙp��͖�×��D,�|�u��s�L�M<|zܺ\��h Y�0m���:��c�1o-E)4���F�tj)�BI$���BBY�o9fsw���TTV���v��	>:��bl<��2��Yi��-�x@����M���d��8n��3��{��:e�$'��v�-�x�:6<4I�z�lv7�Ř�@�}�O}�6��2F#K��ыn�5�Z�D$Q�þ�K�8H=|�p�^46�����-�=�5EUJ˱��� ��uf#��t�dc\O��~>��ƾ�<I]w<��r&�p���0���.�$ːۿ��5&����[���x9ᑕ��`t8z?$�#��2��m������1�[��<�������������w������U%�T=8`�V���QbBl�d`�<q���C�	�5e%���q�ҍ���Mk�Cnj��caǉ:1��F�ш�Pd�X?t����v`�[x�c���d�8�Ѝ���B`���&�C���M���h:�0j`c�9�����w���5�ck�y����p>xF�G����a��S�,(8<4y���>u�����$:e�����g<r8{Ad>`��߶�%�=��~��.�C��4�~�I��:���Ԗؗ����6��m)�C�ƳQ3��b1I�LRv��1���'��b1I�1ı�RX�]F#�K��wK��t�����.�w����#HmF!�}�%�q�:��G��y����R1�C�1?bӈ�1��1F!lN-8��I�u���X�b'��X��E#�b!�F4�D1;F!��1�)8�Bؕ��'�GQ��q����'��<�~�1���m��b1��'�'��'&"q��8���!�Z1b|���%��<ClKKLN��i��6��G"#LJ仹%�K�%�K�.��F"P�8�G؍<�A������F1�F'�R���4��?5���O���q?���N!��%��b�뻞�s��)��t���M�K��Ą;�]y3�d,�D��T?H1���8J1�e?Zp��3�4N�#�i����.���>��jc�O��Nd ��T^c:m���sk��g"B�<4��Ä��f��!��L�C7O��Kty��I+�3��44��b����Ӣ>�goP�q�J+B6���ش���5���	*���qh��<>��5S�]�z26�~F��pi�Сɟ�K^r&^��F�a[�؆ ��tܿ�zs˙���P����h�$BL���sr�G++���~��*kS�(���R��1SM��Ko�h��Oz�b&���n2XJTRi�J^��F��<Dp�KN�u�HqT��~+Tm��BR��)6�7���p��I����f��	k�(��X�D�DT�uK`����1��Φ%K4j�D%AKa��G��A�1����5>8r�t\e�%$8��>�Vg;���lE(7чƗJ����|�#���m��$�(C��w��R���OM͒�]�(҂�5|��	w�7���N2�D��jIrU"�K�1���FG&�D����U,�.���ꄔU�Fݰ�$�tk.��`��r�����9~�]��MZr�ϋb���%�������.�毛)���6o[ʾ\����[_jJGO'�y�D�w�>��zE�/D:�l
�(�!�B�R�D��/��uu����8�,��Qq�G{,�lm$�<��$B�'�T��#k����;H)l�B��NY/U���*�+I{m{��Ɯ��M���c�Y��!��y�U����3��V��X+R�C����v˪��5�X����*r�~�?���~�UYUi^���?{wwwo~�ʬ���Vg韽�����}�VUZU�3�O�����߾�Ҭ���������HSjmM�N:�<�1lcx��8#�<$!|��7� x�BC�(�"9��㜲ؖܟn3!�h؇�(�\a �7����I54��6��K��D�2��⧹�Unw�ܾ��I�W�[VT���.��M��E��7]�*�^z����$0ٳd,�7"�1�m`�J��eUD\���ç���v��*U����
6�<v�������1�`�������NF}�v◑�:h,�p���!%Q+.�p�Ã�M�!lr����v�ޣ"{��*�%J-�n��lq���v��ֆ4Bu�ଃ�7��pw�������%V��ﯜ��2B�(5OF�X�m�CP!>7�E�ű�W"��xuSޗM�ݍ�"���/��k��,�iˋ�C��s�x���E�eJ�w� d�s�hp!Dt�6�lc�y�1�[Ǟ<�h�æޛ����^��m���� 1��+U�!�s�%���C����m��N����~�w��L<k<p��2ڏ}��e��Ǎ�ω(�v�����RaU��`���ƃ�$uc�D����+��8۰��p��5U{����\Cϋ���>9Cd>�'�������{KWU�hr@�oO��dc�r�Æ?0M��F��}�y}��Y��T�^�ڒ��}i�=l#�����a��Hd�J�̴�Ad e�����Ç.�Ą<i�t��ƃ�vj���O�:�ߠ�M!m���[~y��1�c�ǞC�}]�Mk��ϑH�jK�J$�rDdL�B<_9���珮�x��r�co#s� �g���<�|��׻rG.��;f��:z�1�!�`�`B0Ig
p3��<���R��0�#���|�pB��%=�a��iD���!B~b?H�Ȧ�� ���KnZǵ�D�ˉ�'�!��l~p������f_�堍��p��	�I֋xhm���XY5AmRr�>�䇼���@����ˑ�N1�>���#M-�`8Bi��`�;$��`l���0!N4��t?f��pL��` ��<�Sl[�y�1�[Ǟ<�0��,�O�=`�l�I��fTm��j**+BC��}]�l6V�D�IN�hhL��B�� pE<�x���p��m�?;pv����!��������	u���v�Y
=��&>st��q��X��W���޴0/O|��h24�׎:��&	�|!2�%���S�ͻ�I`iubm�P� Μ�Ʃפ*�/�˰��:�A�t>8c%I���d��f����N�m��cO�!
:`�	w�ƓC��dl�0�O�&BX�Y�x��}�Q��I�o����n�7<�-���̎h������V����~zp�J��i��0�
x@Ϙh2�nÄ:��Y��9u�`��!��mm��1�<�1lcx��u�>��Bf'�5��n�9uM���"V�2&�I��pV<D�W��s�!�*�d��t����	fLCY] �h�A����m�M	���������]IH��l֛�IK��
���5��	d�+x�/��ϑQQZ�g���'i�K%�"nHZQ�R�ܺ�����I,8Cmd��8���6U�ܭ��Z�cQ��=����~�~{��0�8��M��x���>��v��g��:[UU&a��{��q���g�B��#�.%J�`b�M�C��)4h���p�;�����p���>!�A�`Yl.ά0��)dV$()�GR(��N�q���8B��0<��m�6�[HI<��Q)ҟ��_�c�c�1�<�]C�ù�o{��6���А�M^�BO<'���}�G��aF�=�a�.G�^i�h�t^�4��n�1�:s[HL8�d�$�8T��S�#&�<��	���������8I-�}�堸}�v.c���|z��;v�,��H:�󑳏��t���1GY 2�G����b��V�Q�d��I.��>�]�M�5_Wxp'^�=�>���r�-;w�}D��=ˬ�g�����^��ԣZ�ո<yӷq��|��Q�Q�|�J����E���5�"���!���F������c�1�<�T㐙��K�����3�O���� )2)���f޺�={��~�clm��|A,Ɋ��̹�������p!P*1���d���N�p�Z|��d��˦V&M?g� OS��V�|љ�����v専(x��ߓ˩�BB'Zzn�tsT��*ȗ�;���=��qi�=�:�ϰۺ�<l9�C�S�����xt�ueZm;_HF����de�Z���nK���!{�>j��A!��2]�x�J�)�M1������3W��S�O�=<�h8�8J4QUL|�,�0��gʹ;v��˃�
2F��n������1�[��<�(��SY����hܜC��z��(���	Cڇ�W}��^T�K�Mӑ�g\�^<!�×�}��0߼4�|�tC<s�g�`�VWxpKG\�9Z{\��2�U1�rL��n��4�i�q��|j�>�ˇ�`t�'�bS��g��ac��C��ϒh6Ce��~��$�zѽ>pa��l!w���9c�ף�5�-|�,�0x�wv|�����Vt!
c�pq�����"�g�Ǐ (�lg����-|@�� ��z����<m������!�%�<��~y���-�[�y��}��RԙB�B���~;���NjчvAUK�D��Qvő�(�,CEz�d�M2�����h�DQ
#���T�!�9 ؆u�.(VZZp�ְ�;*�~fl�;툲�?�~�.N��(����Y��j�J�%i]E�����=��QQZ�Mh�P]mD��m$�A��r�D⫳#0S��r̸tXy�Q�o۝u�.�!TS��x��29��d��:z��D�rL�[e�2�+�wo]N�-�X�L��A�1=�Kp߹�I��M�C�0d�U�nX�:r����@�S:4�p���uQ�CeJ��<r8vC��?d5�V����4�4C�Բ�d��T���A;r��m��iV냪@�¨���������($2�aN��ʇ	�@�A�^��1�8�L���y��4��b��y�b�ż��y.�� �#�yM�������=���z���1�6��BϲÌ�3�zp,�:I�8wP*ɷ�04�!1�neI-�Bt��N[p;�0&�nfy�m,�B�p�y㇅��쫕`���9�ۗ��kRm�����٩$�Bw�u�G9zI����l�pH�wX���s[H�����ό��gZt!�r�m��������6t��'��~��tC7��KsC�m����q��*�aWv��8֟_�w��uO��Jh���R󭩥6��i�!E�kikZ�Z�h�$�""X�h���YBq����Ye�YթiN�-�xI(D�,L4MD�RԵ-KR֥��ZYKC�ZO�"& �'DO	� DL4M(D�<&�%QD� �"xDD�"@�"P�.�e-K[�-�����������҅�Y�Y�-m-mku��M6���ԥ1Jc�bŶ�1�1�c���q��e�Ye�~iKC˟��8��-��>�����|���)��x�4�8\��wk�N���gt,�ǱNiM�<"q�'%���w���^_��>�W�K�m6�n�����߇>�ι��d2��;s�nC o�
}�uߎe�s]u΄��d����z����]��4T$��J&,SyJ��M	.����Q�O�=tu�Λ�^h�3�fɝ���;�g�]�ro�i��Λ��������
�}��s�UZU�_33�����ݽ��*�*ʯ���~;�����}�U�YU�3?O�����Ͼꪶ��Y����A�^y�m�1�<�ű�y��]�&���mثy�)�4��SQ7S�y�s���QQZ
����SY^��m9$���!:*�@a�aۦ���t!Cp�\��|FE�����Q:�Ì�|�$ձ��oو�#�5V��sK����u�]ڳ�G`�	Tm������~�z���n�ӧ�:��My��K���ܺ?!�,��G}��nI�>4�K񍖒�;�6��r�<���SXp��5���m��<bM!r��\���G�Dt����,l)�4��ӊmK[�y�1�c�Ä8&�||C�F�ɟM���U-4I�c������v���͕*ߜ���;0�����|o��Ln-DT�p�T��,Y?b��q|YMFMU^�?:r��f�����P!�T%3�:���#��1�?uu�ˡ��y�\(���}6�1ސ�ۓ�-����l��y�e$�<cѠ�'Ϻ���2� �c�(Y�S�8�6{��Y�����8���onG%F�;6�cl5;cǦ�M��\y�m��<�ű�y�DtgO�!�KI��:L�ɺR�iV!	���l�Eg��6��"L�2�m�2�U���*QDD�T��ɐ�$lTx�7�� ��5�he�/��Y��y�0�_�"JQ�3����o[��l�R��VIZU�ʫRQD��U]��dU$�������&͉�c�rĐ��.�0�8�R8��ʊ�d&�p�4�x6A�'^o'�9�9�~����_m��[��L��bU���yn��>=}+�h|�xq���Sm9l|�il�p8.��b�U�͖�64e��m�_m�}m��B�8r��f�׮��Ì�Sֳ�����h�6��BK��(yۣr�p�GuSNG-0(��\�q;J�M���rb[6���a2m�`�$-<��N��nݴ��ׁcaN޴�^SކkNڎ��˲]hì���m��iǛ[�~y�1�c��!��4��n��R棝Ψ���	�5��%ew++��`lђM������}EK�#|�>f������2883�$�5���/6�˝�S��*�<un>����1]�$�R��������7��b�\v=R�0�_F�T���:��p����5��XV'�I����:^�|�/�|���{��ɐ�d�x�p��.	�ô7�c�n��v�88*y�к}N�'f���������lbȉ�������<J�1|t=(��Kg'�suEʖ�cy����d�t�fN�����c�1o<�K�w��V{�w=����u=ƌ]kd]L�$���$	*���������О�����.�67Mi���c�s3�H|���j^���f���T��ͿM�7�]�t�_�:I.녑�?	�x����h�w�������&�|��%�W=Rc�^y�"�+l(��T�U�׉���d�#Q��[p<~�$�9|����0M�Ɯ9r�%���Q��.�$���v�|Y&���}���i��z�|T88od�#�Ց�RY*Wp\r�G�X`x�.�x�ɪ�\3��fp.������9����qAm������c�<�J�in�����1�[��y%��yI)<�}�_7��}稨���W*�U�$jOeG�S;�<Ӟ�9=���}��?�4�
cH��B����CF����~<��C�,���=~�`���srse�T>�n��CG����Zm&Zf��N8��8���̰̑ޟ�=o�gϩ���?{_GM�1�2G�U-��Al�<t�xbN<��h!�R<;,�ǎ�����]��ױ�Ɔv[�L��Ӂ�0��(�Q��0l�ן�y�b�ż��y.�i�u��XO�DO6�!���P@��4�6q̰QGhB�V!"�MY�!,�����Ҵ���b���W��Nn3S����u����I�Z�.T���)!������z��-i�6�[J%v�%���J�-e����6���j9��R��<�(9%j��JZ����/����\�{7i��._�#�����dpv��nb���f�Z緊���N�#����8�{a���NOu��g���;�^SVppR-�;t��_0`d��C�=���:n2�F9p���Z�{i� C�LT}.�z'O]K�H��g¥Vq��<��� L�i�n�2�����6������| ǉ��"��ٙ�dq���.��$2-%X�Q6˔>�<v��q��t�~1(2p��:z�#�"&��Cs��(���8S��~y�c�-Jy%�;� ��ad��g�q�=0�G��pB����O�;e}7���#����$�t�|}ð;!6ӼC�:p(�ə$jߦ\�o{�J�u����<�[z8~k��$�x��s�J�pk�ܹ��/�&ԑR@�Ɔ���tٗ'8v����g����n��SFŘ����x��}Ϥwo8�x�2����gL6ۇC�T)����aE߫����NƝPQvrT��ŕ�]6�ۂ�=t��i�<��iN��?<ǘ�1lbԧ��]f��4Co6�95�i/�No�e�D)����̳�������@���2�IXg�I��Mr���Cl�4���z���a����$�i=;xq����5,WK;�:E�΃?�������g�}��z��E��6�;�?JpJgY3���g3��A��!�R���p�ˍ����sZzE]�"�d���r��t�S���v�ͽv>4�1�C�絠��I:WHJ;-�~m��]a�c���L�c��`f{]6RY����Y�Kcwpesڇ]����x���y$�Ӏ���6m0�%��J�e�[��Swx��`R۷�/^:�+35��m�Qd4��Z[��o�?<�1�c�8C�l������]�4��QQZ��t۾x9:t���Իn�L��׌r�����~�t���������y�,m��wi�s.�b�l�	���!7��] �vB�e����L��o��x����5]�񗭱�����j��Ï6T�c�N�8vG��t������F:
<I�m��t�d�F�1����//�(�£��爛6={��X����2����u��@�O>��XN��޲��Gae�}4��y͟=rS�����ɐ��p��0l��'�m����Zֶ���j[�X�"H��"h���	��f��e���Ye���M-��DJ,K�4��D�0LDDM0L(�	�Q�0D���"I"%"i�"iB$��$I<X�� �"xDD�"@��h�%��"$�%�bII��	�:)m+,��:Yd-m-mku��M6��i�Z��)��1�m�[�Z��1�u�1ƒ�Xae�[�T��Ii�1
>c!�ሁ���. �QÅ)�"�?�ZC���mq���!=���4x�2לܹ�Ћ��<C����S��f���T$�Gp�D��\��M<L��;�!FT3�v�DȄiqcY��i�,�W�섩��5�LI^�)ůT�3��8&��-�ei��-TM3,��Z�Mx���()`�z�D�6�(3�׋:r�����u����سJTq/�Ʃ���k����QR"�#�<Q��Ч�Kz&wm��o�,wY�/v�������3Kh�\�2�pD9�|7*4�Mx�1A��~f�9�])i���[�vA�w���80�X�^C�6n�e���b��?"�9ɜD4HC�e%��#�1�n�Q\�CI���k�MTW-ʈ�-!l�7����bm����&R6"d%u
�Mɿ	�9ѪK�7��!�5d����Ppӳ�jH����?�����1�(,N�t��U�R�#�u@wF�����y��?ג�2bX��u�U���,��}��l|��ڸ�W��E���1����Dl���7�魮�2$�Hr�hda�F.���[r�u�$��������B�z�Zq�Л���UqIz�J~7H��ꪾ�\��9�V���{����h�[z�~\��c���rq��]��g�J�.%2�淋���)/nUe�[�$H�����=�Wb�v��S�u�7�b8ӓ���O�	g�c�#Q�`���~�����uT�o\�rbI�5[tj���	��X5a�A��#*��Rs�w���j5dHR7G��vu��Ud��8�M��Ic�EmD���[���F��mn[��I]�n��R"U\���Wjk�z	=�z;��9�|�?uU[Wʬ����n�����uU[Wʬ����n�����uU[Wʬ����n�����B����Y����A�L0�0���<ǘű�R�C�u�<��}2F1p���!�Ӌ�f��� �h�Ls#��
���
,n�,�Hʇ�ңM�j;Z#KG�-��Ģ�A\yP��~{NE*��{͎�&���!�i) �WƱ���q�/�|Ֆ�F��Ȩ��	��D4(H��V�G�I$���^C!!%�O?k�a\��p�ye�y^T7HC�{#+ؙm���$�ӏ��x�l!Ǿm��o7x�4�AF�^>��v�w}g{�>�W(�gU�M�8[wz���M>~�NQ��.���Q�����#���agr1�1ƣ�'i�~��;1�M��������I)�M�(!e��� ����F�kn�?����Ɩ�JQ�2�r�m�/g߳�b�5��>pωM=m�z��������ͼ���Ki�����<�-����Ä8&ό���#��Tj��J0�,l:C�v���Y�6��/�o��`r�^;:v�]g�ΐ���>�W�k��2�k<�BB�D0x�ĩYy�&^�$�B����=t��/ÖޟB0����x̻x�`Y��.맦����r�������X^f#�C�څy1'x�f|w�x`���҃�h�N�t���B@�#�w��E1��$�F���<u�:I�2�$�xte��NS�s�6�<���u���)�1lb�S�y.��Ze}�6�B�LH@�$*�˾p��EEEhHj�`o���h��������?�$��~/�2�Y�����~ɓ>7��N���o����0���ʞtq�3\8H�!�t�{��*8^��oY�It��.�����������G��}E��ܟ��}�����3sp�f�6Ԑ�L3	%H�4��|:9��À���}�A�N�L�0���x�,�*�<�������Zx����M86�f�!<�ð��&�ݘ,��M�ML7��~����}�!���N�����c��1o)�<�Z㈔;zF<�>�!	U	$��7)�kM��H���	�w�ɇ�o껪rt�X<`�'LK�#n�l8jp���������g�`����J\r�G��k�mJ7g���)��;�N\�Љ�gG&��E͵L�⍗U*�!4��i�2����Tz�{X<�E����b]����xw5��EGA�8r����ߤf��i��ǣ~ð��6�<{�|��t�O9�C�$���d
�����#��Z��~f:e��(m.��4��~y�Sb�żxxC�l��M�xB�.�̦H#]���F1�dj5+7d5<���6��b(����͒n<ܱ'�joc WK�4k��1��7��c����'�
U��L^��^�vjOc��2J6*1"�YlM�Z�"�DB�岑9$���m����7N�����?�h惱���o~c�4�:Ӧ�����c�]��$�\k��_X���Wt���g�y�IJŕ���W*�ʳG���x$d8���t��(%�����ĵ렌a��1d�0����c�歕�N�c��=u0|W�0O�k�-/./��(��y����?#���0�$8?O�����ۆ4��uۺ$���#N��=!�O��D�с	V9ixQ�(��n�d��\"HFz��G0񾱌lt�Q�����G	F��6W'\=�}��Hi-���ǔ���1�-�[�RK�[�:ڡ�5Z��]�TTV����)eU�D�ka�o>�C�ʪ�6:�ˈHM2�:88뿱[��p�C���		���:I��^��߉0�t�,���
M7��Ɲ���<�p�*��p�!'�:섰�a�m��B����sF&)�P���j�o{:;���(���|э�g3��l!��kZ�ִ�,m�A���_�Ѧ͛7�n��$���O�48��:�?4�0>��~7GJ�uW)�/]�u�s>0��FHZT�ӭ?<�矘�<ű�yO��柑��~�#x�U�_��6��М�k�o��ےs��W_i"�`�!Lm�B�I,��og~.�˽?ÇNG�޿]_��)�`�s@Ö	���
�Y�M�y�-����$����JpɷvV�Q��щ\��G��Xd<�qA�ۓ���F�>�ׯF��Y�d|��)?��>fd&��H*22\���2g�q��AD:H~.�e�X*X7]NI)dM�ZI|�!�����V�#�H�jڔ�9J%(�=.��"�"��RN'\ly�iƤ�j,��$��Q'ݪ�(�+�X!���lV&�kM>,r+��fs���s����GpIP���2���u��!�e���`4�����8[UA�EI�.���t\᎘$˷!f�i-�4��Z��~b�ǖ�-�8C�0=�X���jjH)���h�l�8�K�!V�D����*FVD�%y�f�L�1n�"8�x�T,�a�m�E��0�!�OI%I�]�]����!��VPm����B�
�|��p;Z(��E]m�Ć	+�<z�,��L��ACq3h�a�u�5�E�	#�{^��lE�T�Q���5����ӣgА��W#�$��8�6u��ׁ��u�M뺐�:V��{5��!&�;f�=}�i�Kr�(��!o`�8���O#R��4u�׵�uK~��Lt$2��1��8��Z�B�;1���f�8��ۍ?4��-�1Lc�c�%�27H��ICzkHC�ty
Ј%ʋ�l���ZtK��
:��F�٫��	Z6�+���B@�{%,¬N�(��JA�&�o7[ڿ�}��Md1qE��R��3�H��%�U�L�� �Q(E�e�D�X�G5qգ_QQ��)�Rr���-n*K#�����Ϙ<�ǌba��4��5�f�=��!S&`�6[v4<m��2��Ilx�<�=�BHj����f9pl!NJuf��/�݅�ݐ������+���۽�Q1wp�_c�=�:�M�zXY=��&�g<a����kP�����7ۼ�.�*���m!-Ŀ4��~C�u�j�|&�X#N�o�����cǯ#��������(�|�􏞙=-�ǎb1�J�tvӧ�h4`�%�4��֥���1�-�[�R�X�-.5.RW.v=��9�g�3%UT�a��v������8֪�u�e�Z�60_�0i��&^<C_j��o'��4Ϛhn_5��3O�k�sO�����#�(ӓL$�W�@���Zc\��й�c����b�"!"�!���c���ڍg�3��	���x�Wa�&�i�Aӭ:��:��l�!r�^/S�#���J*VB$�Zl��?:k���o�UR��=��Ώ_:}9���C�yM?6ڝ~y�8���f�"$����a�HDD�DDL(J�	��A(N�I�H�B%�lF	�h�&�&��4MDDM0L(�"I�D�"'D�"%�&�"&	bH�$�'��A�""&��D DIΈ�"&	F�X�@�Q��xN�$��qB�����DK<"��J�m�ZԶ)��1�m�[�Z�����X�ia�!�af�⒤6�v���"I[^y2�<m�!��V���<��x�����44F�$�f�ؒ/�H�C���(��N�15�}+Eh��n$��Rɢx�3]*#�j0�vH; =Ò�0(�WEb�bBT\D~�� ��������#��H=��|CB��x�7ID6D���N�Z"f'`QDN���؝�L���F]�IVҨK��ȕ&;"��r�m�����$���Q�!�jD$��x�$NDG��M4�>���
�^~|s�z9���v~L��~�^�8�؞��Ș����2]�*���V��Sq�q��d˻ߵߡUW���̿����oЪ���Vff_����߷�UU��33/������"��/UY���0�<��<��Sc�<�1o)Dx|�ӄ�H~�.��-�������**+D���J�n�>���~N]�d&�.?|>ce$��}�O�=u+a�q�L{=c�ё'���a��m�i�I1F٧�~x��ӏ~~y��HV���\����%J��R���t��R��JmE����I�2}�$��������4��n<s����Q�NIr�;ӿ��S��$����|�8��˧÷��	�;�m5��Ͷ��~��Y^�ϣ�,m�����D��.����붝��&,�EYT�&)���L4:x�^v�VL7��>:IƇ��}X6��N4�o1O�?1Lc�c�:��OЏ����P����(d0`��H;��I$!x<<�g�i�<$����e��B��P��m�����/\a�nMW�6�;:���D?�!d�!�8u�D�5��ܴ�X��ۻ�K����BC�r�}���~7�I���̺��n�l�7
6`rz�d=�]��m�K'�ݏθy�n��]��T���eقǿc����.[�4S�|�&J��E���an�yC���Ӝ6�,��B4UPge������'ç<\7Ï��K�Iu%�Z~i�)�1�c[���)֖��qmU�i�0�����R�j��W���)��ұNMs�K�ǴJ����2@�i�e��{�<X��1d��H��D
Q! ��㹝��/�{�S>���&���.A9��˯^:�)��lo ƛ2�H��cި���Ù�C��A��B�!"��MإJU-M��y��_~�yf���n,ٟ���4��ܨ�M�~V���Y�t�ކG[��B�zt��y���!eM����Q�y�B>$ƨm��0��*T~��`��}�gC���%d��y��<��&X�Lsweʗ!rv�c�N!Tro��Ll~�o��O�Ϝ=�C�}�ŖJ���(o0-��"RcF�����3��~cǓ&~�iܧ� �O��ڿr/�M�M�_1r�I��wDa$�����4�8�:��1j~y�S����O�8S�3��έf�u;_1QQZ7^RR����r�*WK�V������c��j-��j�:$�9�����
2�a�v�및2�QEUG��J�0�$avᶗ�w�M2��n�"I7X�n"���MB����ۘ�m?��*Ӎ������� Y�an�옞t��i^���|��8x��~D^r�.��7K�.*��e��*!d*��\y����?b�9�8��=��g���V�pr
��F���o4e�;��虷0�o_3A��&�B�Ip�7i���6yHy/�4�O�Z�~b��V�<xG�Ĺ��ܷ�JY�]�y��b��f�%��e>�x�p&���Hb�p-�4��1:mˮ�˝i�����2��}D	��yO�/K�� ����B���"VJL�&"��RAT����k�M���jY�>^����c�i��?a4�U���7^���1�}�i����M6'Y+�:z��׷�̽���dv�� C�@�$��##N�N�ICO4�Jm�o1�c����)=GP�5���L�iw��Й:z��7�uQ?��*��B�Xŗa
��˜VdGU%'���z��m������:B�n���|וo7���i�݆J}Γ�8�L���ͪ��ݢ�Ԅ���[�Nt�u��6�6�ve��&��O��P>�m�2I�/����^(�Ƙ�/\�:�ɉS�Lk�}eUo�鿚wO��s�T�u)��nG���K6��|m�8��?���B���'"�հ�9��n|=-m.������������n�`��V�Jq1���ߟ����1�y�=8xxC�e�<�9��hbKOj���|C�F�¦ԈLbitlN�&�!��\7 �Q�LeX����J$V8;���"piBG����)"I6�޾�My�ҫ[Ĺ�݊�"�6��kՋwb�u,BN'��n�����Eɦ�Z�J7Y�h�Z�L���4�eX�k�ϡ�\�+ж�"�f���Œ�
[���}�|f�o�1�$�p��BN?�ã�ʪ����=,���Q��7�	�`>;4��m�19�O;1%&+����kE���8kN]��o�;Mp*��xj��/�:3$��0Rxz�1��E�3�#4\�!�Q�V�x��HZȖ$Ҳr�(�$9�bD=�9�z��yiv��g,�κ����~�">r���(��n!ԩ��4��ߘ�1n��yJB�i*4�n!�����1��k2��������|�aFy>��3�s8֯��Nī�3�xt�UO\�r[��8CL�}-׈K�����s�*���W�y�4�$��x��<��iӡ�l>=,�Uq�3.�>��e�]u��Ő�������M�!F�b�)(Ɨ��Zc%X�*rB6B^av�!'pI$a-�ƗAG��}#��zn�98|f��!6?[�9xɬ���G`x��2�˪����o�7����֞l��N�X�2l��4�Jc[�1n��yJB��S���!m'�b=�y>���.�EUTURi����:g��!;=:7���J0q�q�d�$q�e���gsVOcK��)�"u�X_�|��p�=�z�㳤�n�f�V0ȋIHN���SQ2#�y����fK�����I��r�>�װ���qn��]0)�d���q6䝠��$��m6�4�˦��6�li�?x��YP��$�|Q&��4^����sy��N�u(=AGx��ű�1�ձ�c����)֙^/7���{�z�s�@(*�	$�T!51�͓y�w�**+G+Κp9�e��0�F��a>����d4K����ɧXV~����?p������/u���?s���������wܿ�w��9>���������G`�W-����r���4BK����g9�I>ۻiޙ��R��^�x;0k���/^�0:ni�c�d��._}n��4�2>i�6S�90�2�a��5�	�Nqۀ�Q$[}_{u���o�J�i�mn:�qIa.�kZ�Zֵ-Ԭ��DI0M,�(J<tN �P�$��<xD�<'���0��4�L�0M4�0��"tD�Έ�"a��O�BA�i�,KD�$I<tCH<xD�M�"@��"%����o-�[[m%kJ��([hYe�Y��ZV�д8���֦�J�yǞZԶ<�b�6�-o-KZ��qn4�0�0�)5_w>�בm��w���l����CJiBb?�1���A5:p%j� �>�iXp�iWi�8:>�飥�1�:3V�3��5��!uS㬃�\�}(|p�i��d=�b��ȥ:�$PEC���#:G3��["�P$�y�ثRq��f��W��|@�D�'㛨�x���y�H$��ŃRI�|�cWD�Õ11�&.������Hl�2���ow�n[�Y^*-u������%� ��L[�Ɩ<��c�1B�M�Fl*�RG#&F�ɒ��F��2���>8r8Q��	NVЂ#��2]8N�)ʖ&���n����!��rf��hQ�RMG=�㓂LC Nin���	��83X�x��:4�� ��-���	LeT�ܪAi1-�Ϡ�.���R���F�j�("�w�OiM��Dq�
�RA�!��)k~"��B6
DLR�?�F�{M���*!"&�҈\���rٺ�h��A4.l��t����oËu%�����#Nw�]��M��M�y��8B���ԓR�N"�D�O�֢w��kZ}�QNl%���me�!qŻ�2�h�䭢6n�ضr�>sd78-�ӊ�V�� ��uU!��ʸ�.�ړ��Z�K�D�������8�/��%��:�'=u17��C�����zl��B���*��8�q^w�����Ȼ�6�cM�'I^9U��(��}힚�d�x����6s���B�,�ԋ���<���F��^|s�X���t����B��;�d*#nU%|UUb� ��Dq�N#e��9J}6���/��!�M�X�	P��B�$�tu|��>sSe�9�U��X�Y,�MԚ�4ʅ�%�Uh��ʉe&$H�������������Uqz����񻻻��Ȫ��
��̿����|��������񻻻��Ȫ��
������0Ɯi��c[�1ly�yJB���.�S����B �EJ"wFLOMwŔu	�P�n�J��R�d�UCB��O�oo0榴Tq��GG���T+�|�ěUخ*RV�m)K�LJ"�7w��3W���s%�w�TTV�8"�dlY�:��u�e TX��s-�Sd�voD����,�����-�յ���Ԙ�!m׳5���f�e�n7�ޛi�f�nX�<�`�Oޤ1�ð�3��y��ݏͽx����t���!��%y��5A��D�y��тO6�0��±AVCR)_��ɵ:-\�EF�e�w���r��Ο�P���N�O�G�)(y�ӭ�Lulb�ű�-�)
y��K-[���$[F��]�ﾎ�`�"8gg:��Z#�e=��|pfx����b���*�=�*���M��Mn�Z�Z��n�vi�!	�p�;�oz
���㒦��ҡ��Ɯ�m��ZS:�D���h�_�n�.Wn�p��)��VΘ!��Jt�n�!"h�n�oZ�E"�v\�k�x�ۣ2�n��M��O�h��;�5��K��2a�l�1N�2k���|�냤���q�W��5�>����Lim�ku�b�ű�-�)
y�9����SjS[�}�$$%��me�e��8����a��D���\��#nzq�p~z���v׍H
2p�Y4t�]�׌|}҉�.Ð��n�Fy�6۷�/س����-�M�-��-�e���ɟ�
\��Fk��qk�j��eo7a�䔲�呣��f���1�]�x���GeGN�h�CْM�Bq��M���|\��xx�$��′M6�;i������xu��|��^��̃�v�V.��B3!��.����cܡ��O���Li�ߘ���1�c�[�R�g��g&ᢏjBI!�#ɂ����珟<�|��			(�(��ڒ�l���A��e�x�Hiɍd��`�9����������.+�u����2�Rdj���$�t>1��~I%��,�sܒ���a�A��[Q�}�����ǎq��ǎ���+-'y�����dz�����t�t�GK*�@�nZi�����.���I��=;2�TÇF�v�I�EUXd8��L>��f<��OL��cѝ܁2���>aО4��oO}��=�G~�Ҕ��ҚSjS�c�-��o)HS�1�oN��4aX�
��\�.
�������i����g��2�▔P����t�IH�[cbB�`�	�"�.�I��mq6�6��-���FdR}:M�[�}'��h�J�ڝ�L�K^��ZP�C�9E��$g����			a0�3G��R��Y$ ��)#��hvą�I��a��Nc��:0jh=?��kZ��|�$��I(�>��qܴ��O�uQ<�[��$��W��i�D���XS��Ne�F��u�5��~��p7XCN�mQ��cs`�MU1�N�ѫ"K~��Y<�|K�x��d,4���}6IAia!IguL��o̒`�N�9rfK}Z��l��m�%��F�ǝۈ��/l���9��3���|����G�ּ�VUUݶ�;e1�:�.�?�2t��[1����cӤ:E6�[�c�-��o)HS�:�>Å8t�c!��'a7��u��$�Hv�m����nGA��;#�U��ƚ۰�w��:��Ǭg�*�/Cmh�n]�ی����;�&|uZh ����~���|����/���'r�Ϻ���G�'��W����ěvI���̍f�0�ôɠ���XdW#�&�4hJ!щ5/���zJ��%�86F6�9��pr�,����97���nÚ��|�w�1��n��ϋ	L)�n����̚y��n�1�c�X���)�6�-�`�c8�|v߼�9<@�����0UBW]�h0|ͽ�~嵖�>|�3�����Y*��wVR�$��9�8Q@�3�����.V۵�x�������u,�d3�K�����b�����#�O��y�ą�~~�<z�c�CO�N��?>~(��f�GF�	�?��ښ�Q"ؚ#١.�ǟ�䍦��������n ��3����L�1�����m�/�R���wLm�p
�Ca�$i֖қ~S~c�-��o)B<t��1&?��Z�JZ�bN�~��'$�]]��m0-�ќ=_����i�q�4ͅw�"�tލL��K&�`�/���͏8��>�r9
-�]I�rm$����%8�]�=����kX���c���/����!��2�Ha�O�7~v馣FNʷ��ON�bX��;L�4���~	*W�|C��R�A��4I��'à����<I֛�0�i��ZSo??:��)�[b�R���veOvm/��}Զ�Q�s��)��p���i��	�-Tu��ӱI:�8� ���K�26#킨��I�aKP�^����-8"�zZ���ed(�*���U�o�Ʉ%1����
�.+ESA�wo��F���^��'���K�(���2B()S�j�aQ���x��щ��L �1m�MW`��D<R�YnKm�c�e�ـ�8q�m�ۼ�:���N��Q*�T��wMӀ���p�2I�>�*�T�R�=c}vzZ�����ǖI��6r�Z<8W�%�񊲤�珃[q����|z�!<rt0v��Z^!&]��Lx<���$��p/�����Y!'-Ph(�9�f�N������+eUb��a�Q$�l��m�����Q]t4o�!�]�DI�4��c\zi�)֘��R��~[�-�1o)HS�!o3IqT��B��^������HHH)��1��3n�3Ý�n���
{z:�R����+ҽ	�e���~kW���o�*���	�W��G�C'�Kc�|��I�!��䇫��':I�P��y�,_}�ِ)/˲���#��ߟ�]m�O��~k~�7���U���cse��eU�T0c��~>������8��J$:ɲ�U`�?�~���%�\a�����A��L�_�O%��&��$���A�n6ن0�(8�nX�Ɯ6�,�
	u%ז�m���C:���DMΈ"'DD�M4L(J�� �!�$�xID�J0LM0MD�4M�4M4�0��"tD��"A�%�"xDJ:&��%	bP�$�I��'�O	b"ibY�HDD�JD�,�Km���!+J҅���Ye�,��kl�-պ���T��q疵-Ա�1�c����KyŸ�J�-�q�aK�o1��!����z4�77�z���.�����2�<"⾧�e�ْ	�N�O�Ɯ0�LCH(��4&zKl���i��;��%	W�B����u�y3��pB!	�`�κ��9�⛍ԩ0�HIV���L��=駢_I��=��߸�/݋���T�Ny(q�����4��>u��U��ؓ^��~��UWXUffe�cwww~��UUQU�����������UUEVff_�7www�UUY����C�4�O6���ű�-�)
y���1�6�-��c]��\�!HH�r��]�Jf���Y*��82�N��r��q��������HV_3/3m�l�i��I�L�>4�g��q��P�����Y�w�tmf�V�[�	&��uL�?���?ޟI��Ż���{�ֱ�>{���H�_�9p�>a�a�|9&��i�F���psĪ��y;'��Xӆe�ħLG߹�ﬖе4����[��ylb���<�ZShzCIN�Id;�$�v1�u����{�I<��W[�x��J�Ӗ�vɧ��!��%��*+- _��S4lRYvȧر|Iw���>���9�����o�fI&C���	-�~���qߤ$N�i���Xr��e��փ��CDc���s��A#�Xo׹��W�N���UƮQ�1�S�i��1�L���C�&ك�e�_w��A�P��1�6���-屋cL[�R�M}�}��S��[ƾ�C�Ck$��,�C�� h�ic7I���Q�E�9��k��81�G(���aKl�3ZELL�pq$��.��r�Q�r@���nT�b��ڵ���I	- �=h�K�5�,G���U#�jb�\Rs��j���%�9[�h�M%�B=ȱ	�Q�cm�MN�����I$�B��(2�N=)b��Zvh�*VAbHG�t�׭��r����ǥ?4࢞Eʸ����ӆ�e�\:t�u�Pp�Oi�^a��	>q�1���8N���ri��t�I.�/L�.p6:��Mk�{6��0�!O������b<:\�#�Q�h��[��H�ߞs/�!+��sq{9��d�Ǯ��]v�h�k�^*��y�H����XҚu�1��o-�[��R���C�q��)������,��gܒI.�$��RQ&�7�ߺc����a%ʰ�����ߞ9k�n=�p���g����^��}��3}Ⱦ/���������	�تV<Q�.����$/}�v4��X�Ζ�V����8���>�f:,���Z��ڜp�D~7>'G,Go��UQ�,ҍW���{6e|N�2g��FЦ��m�d�vs������ܧ��Ğo��8~s������<�}���
���[x���Lo�߰�hm֜i��Ku�o-�[�R���{�;��mc{uj曻�ϸ�I#Jti�7�D%����EN��b�SҸ@�ξ�=�,m��$��Zy��YUA8���vI�Z�S\�٣���������9�*��re͒	�#rQ`$��0��<'O��1�{x�ʦI^v����;>~2Y��W�����xe�:{��R�+�s�$�r�5C�p��ٲO0ӡ�y:̞n�0��Ӄ�kh��N��>�kC�4ƞmJ[��ylb�Ÿ�<�kJ֖��Ǎ�٣�n�U�Y��w��ܒI!�����-��Q:ԲIOF��l2��ٶsn_������!8��h�F�`���b�-D,��/��9���Q�s3
�wV��t����?뗅��&�p�U@��Ī�Ü+s�:2��H�a۽�:��Z�/Ÿ���M?�"�rّ1[%���������2I�ڏO_L1Z�l�+2���2����e�|I/�N��s3ជ���	7�8:�84�=	$7��
,��i�mLc�[�[�1�<�N�>!h�
��
Ό��؄i
4��D�%Q��J¼tU1��,���G/۽?�E��
^ʪ6Tە�M4�"6�X��̎d�\��ZAA�?[��:��픞8'\�ŕ��C� Q�IŅD���ջ]Ѯ�5��k�jIID�Yc�$+��I%i���d�W��$�%jzN)(2����ZBm(K.ʹ��*]�BH����yr<Y��|�:석��T���Q����i�Ƨ�<ʏ���L<tc�޺:VI.����7�Q6|�3�����3u�铧���F�t��g�ζ��%8m�Ot|ӗm��f`�^�v��L?��&f��p��ބ��JBB�$�*�49w�-�ݹtP|��~�f�x�F�MM�O���]B���Oͭ�u�o-l[���u��j��q�=c{ѹ�I$��H�D�����3�ϫ&�'��^�6Y꺗ur�I��M[��e4�%�$�p�����ܽ��%��xO(�芆�S��%��8�ӧ�e����EUV��ӆ��O�5�Ϝwﳏa��ˏ�OoLÓ=�Bn��գiF���km�Q��"m&1<��A������\O�g��:��\�w>���D�M�W���h%`�Mp��z��V�f�����z~��#ɣ��&nye��GN��O6�1�-�Lb�ҞCδ��[	t�1�����}����W3"""!���)�dӡ�9�9U����fCO�����7�J�t��{.x&pzX��̽v�u>|V�s:8�8��"/�R�R�m���D	#)�ʣ�:g�����}�駱|�^��Pr�h��m�,uD%:Ctk�ͥ=��&km�8v��G��,侹#N��l9��w�!*96S7�I����f��[��Y��Қy�-n�-jZ��1�)�!�<w�w���
;�
�����N�|�o�G�tf�u��%e�n�t������L�b�y�x��e�p�P�(!�$*Yi
�k��8ؒlI>��%�=�f�KC�Į>r��S��!���m�a{v��}A�tt�J��!�N����c����fY1���eTÏ<2��nZ)�a�0Y�Ui��N���鹀�M���|��]kNY�@��,���0h+-�mUJ!���ԧ�R���I��,#�g�`K�
i�t��H�� �����1iLl���!�," @1Ö��!T��V�YRʖ�*R�Z���)jR�YK)jRe)S-D�2��I2�Y��,�I*Rj�s,���)je�R����L��Il�)e�R��&Y��)$�JZ��\��$Z��,��L��-JY�R$���n���R�Qe)�R��)$�R��)%6U)fR�S-JY�R�ʔ�jd�e2̪�7,�e�je�fmt�s,ș$�2Բ̙K*�IK)%$�,�T��$�2eR�I���eS,ș2R��L���$��I,�JM%��bd���%��l��e)2Y2R�-nY2R�)2YlҖL��%&U-&IK,Z��fX�)e(�Y2d�ɒɓ%-�L��%&L�,�l�ɒJKId�d�ٲd��K%��T�d�Y2d�d�J���unK&L�L�,�J[2dԙ2Y,�L�l�ɩ2d�ɒ�KfJL�,�2Rd�e�ɒɓ&��d�f�ɒ�&MI�ɖ̖L�5&K%&��fK&JK&��d�e�%�&K&MI�&��%�%Id�Y)5&UԶ��ɓI�d�dԙl�d�dԙ,�5&[2Y2d�dԙ2j[,�L�,�K&L�[,�L�,�K&MI�̖K%�&�ɒ�e��d��)%2Ke�%&RɒɕJM%�Id�Jd�Բ��e\V�k+-R��Vj�ͬ�ڥeZVUJ�l��W�Z��R��Vj�f�Vj����YY�+-��J�-J�R�jVm+4��Vm�eYY�+5�]s��� B�! �	��ʥf�VV����YYZVU+5�ee]+\���V[+-�eiY�Vm��� (V��+@�U�e_�iY�����Ҳ�Y���m+*��R�T��J�iYZVV��Ҙ� ��l�bj��iYjVkJ�R�ZVkJ���Z���f�e�VZ�el��+-��j���W%k�ҲԬ���T��efԬ֕�l��Ҳ����VV�fڕ��YV�����++iY[J�Ԭڲ�j�Rڕ-YSmJ��SU*[eMjT�J����eMYR�*j�KYR����[*Z�J٪u��2�J��TեKYR�T�ʛYR�T�J�R��[M�Y�K*���ͶY�,����Ye���T�VY��[e��eYe�Y��Z��R�jY�eZY������,���m,�e����jYm���YZ�*��m,ڲ�VYme��������6��kK5R�ZY��kK5�eZ[KYf�Y�K6�Y���l�if�Y�,��Ҷ�me��eYf�,��6�f�Y�,�m5�RͲ�Rʲ�ieYe���e�m-�������ʥ�K6�����j�u�:�z�ܪY�Ym,���eie�ee��6�iVY�,�,�,�,��V�5K6����ږU,ږmK-K6������Rʹ���6��R�R�R�Ye�f�eRͥ��P˖��4��2ܹ�e+,��i�e�Y�e�Y�e���ie�fYe�fYe�YK2�l��2̲�2̲�,���R�,�fYK2̲�,���,�,�,�)e�e�j�k�i�e�Y�jY�YfY�e�Գ,��Ye�fY�f�Ym2̲�4�R̦��L��ie2�)���L����U�R�e,�Je,�����e,����K)e,����5)���R�e5)��R�e5)��jS)e2��YL��2�R�e-)���2�K)�ԦS)e,��\����L��2�SJjS)�����S)e,�R�eYJe4����,�R��RʙK)��4�SJ��e2��SJ*Y[)YJYS*eiJJ�M)eL�)+L��,������2��%2�Se%L�V��)�ʔ��f�.*�R�e,���iJV��R�ҖSJ�SR�U�JRS)e2���e��R����R��(�T�)Uʔ�R�2��b��JT�R��R�R�4��Ҭ��R�YM)eM)e4�,�T��Jen��]o<�r��ʙR��2���))�4���YM*R��U�RʙK*iR���R�ʔ���ʲ�%2��)IVeL���J�**�ET��J�U�����S�V�ee��V�+,���ʲ��JVjU2���VYZYL��YjYR�)jYJK*YjYe�YjYIK,����)���"�"����i)��Oë/ZV��R��'��H�QRPQBH@3�����k����k�5����_�bw����������v�������8���0�"�����������������%�#�o"R����{G�_���a���2�'i�G���O����)����������/��m�~�AP�U?Y����A��x�,_���P�H(
?�'�� ���)�e�r��^��*�y�����}���_�i����J��Ë�B!A�?��?���9�~L?���?�@T �~�����"B�D�a�l���H����R8��A�.$K`��T���Ĥ������@���	�{��4�?����?���,�LG,��	$���:�?Ĥ��H� 1�
	@& *����  �BP����(\P?H ��bb
2 �F*�� SUۇ_֦ ���@�O��D@��;�6����ؕ��DQ>_���~C��� )P@@!GD ��(� ��@ �E���B ��B��?��A��+�Q?��hu�����R���QD@������> �(��%�@��T���'�T'�E��/��\���0b��I���m��`��h�6�����@��_��:!��z�a������9�������������H�����`�~a_������ͳ���?Р* ~�?t�ί��r�����/��<|?��۵)M��?�T" �F�@T ��?h��R+�Ba��X��Je)�?���?�h?P�_y�]��h�`���0�(Q9F���"G��^E��R��DU� 1,�h�6��BXǼYD�����	HR�?߰]���4�6��@A�\L��]�e?<'����P��=A (]�O����< O���ڠ* ~�������U��So�A�7J�?���������������?���.����?�?at������'��������H�_�KL�C��������4v8 ?:�Z�"���~�������h�*#�1�1��,lX����QQQQQ��XѴc5X�llh���Q�,[h��F�4lZ1DcF�V-�cDcQ�Dh��F�b##��h���,Tb�#�#F��F��Dh�(�Dh�b(����4DF"4Dh�Q����"1�#"1�#���#Dh����1DF���#F(��#Dh���"�#"#DQ��#DQ�#DF��Q"1DEDh��"4F���"1Dh���#DF��(ƣF#Dh�Q��Ѣ4lEF�1��h�lE�؍#F�F���1،F�#EF#�h�"14Q(�4QF1��DmQ�(�F�F*"�Q�Eѣ�ѣDTTh�4h�"ƍ�4Th�h��,b�h�Q�F���1�1Q�cF4h�cF#ьlTQEF�Fƈ�#D[*1���1c(�1b,F�j*,Q��X�ƈƈŊ1b,b�b4Tc1�؍lQDThэ�F6,h��F��**4Th�bƍ6��"�F#b�E��ccDb�1��1F�����m��h�(ьZ,lh��F5b-#b64DTcb"4Dh�����#DF��"4E�"1DQ���"#DF#Q�#�""1��F"4DE�"4Dh��"#Eh���#F���"�F"4Dh�ƈ�DQ��(���Db"��Q�(�Q��h��1DF�ш�F�1#�F1���"1�1F�ƈ�lllh�Q���E1�b1#1�Dj"�Dcc�1F�E�F�b4h�b�b1"���b4DccE��Q�ш�F���+�F�F�(Ѣ(ƍ4j*4F11EE���b"�b�����b4F�h���E�F4h��F��Q#b#Db#DX�Q����#���#DF"4DQ����Q"1�#�#���F��F#DDF��Dh���"�Dh�1�؈�"4Dh�"4F���h��"4Dh����"4Dh���"�F�����#DF�F���b4Dh���#DF"Ѣ1#Db(أ�h���j"�"�(�ѣ؈ѣE"�Dh�DX�h��؈�#F�Q��E��F5(�E64Dh���h��E��cDlF(�E�؊*#Dh�4b4TXƣcF���cF#c4cF�4h���64TF�6"�"�1QQ"�QE�cF���F��ƍ�Q��h�1b,cDcDcF4F4b��b(��c4Dh�cDb�h�4ccDh����ьh�X��1cDF4b4cF4b1�bňѱ�1F61�F�"�ѣ�h�Q"1�4Dh��Dh���#��4Db"�Db#Db"4F4Dh�"#Dh��F���Dh�؈�b#F��F���#DlDF���#DF�����"4Dh���"4F��"4DQ�F���"#Db�����#DF���cDcDF��#�Tccb1��F�1F64Tcb*#DQ���F�X�F#Dh��4F(��F1b1�F(�F�h�FƊ(�5Q*(ѣF�4F�h����ccDlcE��,h�F�*(��1�,b�TF��j4EE����?������/�E�"��������~����֧�/���8����-;A�B�B_��c��%h��LV1�"��7���p��~C	���|��?����A��������	��@�o�w�&�@��O�X� ٳRJJ������ڸ��������=����)�����4.lȚA�|����8<E�������B����1�m��,�ô
~���>�i����PD���x0��4��Z�h�����1�?���o���$���J
A��b/���=��rE8P���Y