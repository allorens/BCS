BZh91AY&SY���ߣ߀`q���"� ����b#_                 �                               @
( ($�` ;w�6ö"��e��g�� `I@�+b��r%"  � P @h �,(@,�B�
 (U  �  �{ۅ A
�H$P�EDAUJ (HDE@��� IAD���
�T�(��}�z��= 5�.��
)T�J�V����/{����=�/' t�'�&@7w��Ȼ�Х�UQ���E�   ���*��%V�����k�}ޒ�<�4EoJ��2i픠�����A��cɡJuy�a!� ͏>}�T{��S��&�zy����}���   ��7�IR��S�!UJD�BAIN��*o��l}g��}�^�G��>7˟J���|�+纨+�`����}� �����: >�﯀t�:��c�\ ���_  of"})J���x��Δ>_;;��@yM�����*2o��`�4���:�����3ﻀ���좋�����`Q�8�� ��` � � u��\�R�R��U(B�AEِK}@#�j�`<��;�:f=��P<���J֯Z {�<�rf9� ��� ���w�=y@P ��R�J�=��>x�{>�>�>���@�y�7;�����C�:�z)�J�y��9�9 �Ӑ�   xuO�*� `r�EUP�ERJT��	>{vv�����A+�� ��#��;��Up�w�{�  /P%�@+� �w��c�ׄR�k<��a�@b���A+��v �t���y :@   )�>�)Tz�H���U #lEW�`���{��O{ ��I. �� �H7`�v 9�. ��0A�( ��馂� vw� �<�^ h������� y��zng��rv��g��        �� ��) �  4 ���T��   i��*&$��4     S�) R�� �L�`&!�i ��* �     �Hz��R��bh���dj�S��bz�5?T�S�??�����˫����e�ü����ü�� ��wǷ�܈�*�"���� �*���$TAV:����C�����T��U��\���� 

��}��Ԑ�EA�����?��g���c���c��q�q����cccL�ccLc�61�c�3�ӏc�c�1�c1�c�1�c�c��<c�1�{xcc=1���3�x�Ìc�3�c�4��1�cc�1�c�7�cc�1�lc�1���1�c�1�c�;q���1�c�1�`�63�c�c�<��c�|c��1�cc�1��c�1�c�<q��1�c��1�ǆ1�c��1�ct��1�v�63�c8����1�c��67�1�lc�1�lc�1�c�1��c�1�oc�lc�1�cllg�1�lc�1�|xcc�1�c�1��c�ǆ3���1��c�Lc�1�c�3�c��1���1��g��c�63�c�q��ǌcc�7m��t�1�c�1��1�c��1���1�|���g��q�clc1�c��q�c��1���1�c1�lc�c1�cc�1�q��c�|c�63��1�LaN���<eLedL`LadL`�1�1�1�;aLaLaL`LdL`LldI�1�1�1�1�1�1�q�q�1���D�T�P�1�q�1�1�1����"c(c"e&0�2&0�0�1�P�D�D�D��1�1�1�1��LaL`N�SSCCS��T�D�T�T�D�P�����ǂ�2&2&02.0&0�22�0�=<T�D�T��1�1�2�CC\`I��1�1�1�1�1�q�1�1�1��@�d	�1�1�2�CSSC(�1��&2�SCSW(�1�1��\dL`L`N�1�1�1�1�1�1�1��1�1�1�1�1�1�1�1�1�1�1�1�`	�1�1�1�1�1�1�1�1��)�!������(cc"c"ccc	�����������gCCC(�<`L��P��P�@�D����P�P���D���P� ��`N0�0�2&2�0�0&0&2�0�0=0ʘ����&2�0�2&0&0�0&0�&0&2&0�2&0�0�0&2�2�2&2�Q8ȜadLe`La`LdLedLdn�C(�1�:�T����D�D��Va��@�D�D�@�D�T�P�D���q�&�P��D�D������eLdLdN�SGS��D��1�1�1�1�1�1�1��1�1�1�1�1�q�`\`8���8�&0�2�� c
�
q��E�Q�Q�@<a\e\a8�2�2�����*c�(q�`\d`�T�q�q�q�:a1�q�r���T����WW�Q���A��A�1�&��E�T����@�GG�SS(�q�q�r�GG �:a`\d\e�WGW�$q�q�q��W0&002.2'�@��8��`�T��Q�E�q�q�q�1�q�S��#���+�������)����T��Q�����1�q�q�q�q�&GGGN�aea^� ��Q�����1�d�ǆ3���1��t��3�v�3��8�7���c�q�gƙ�1�c1�c�8��1��0c8�(ǆ3�c1��1ӏ�{c�q��x�8�l�8�0c8�ȱ�1��3��8���3�c�1��<q�g�q�g�c�1�1��q�c�1�1�c8�lc8�Lc1��8���x�3����q�g�1�c1���3�M�c�3�c�g�g�1�n��1���q�g�|c��1��1�c�3�c8�1��q�g�q��q�g�<q�`�<g�q�c�1�c8�1�c1�q��g�|c�q�c17�1�g�ǆ3�q�g�q��c1�c�ǎ3�1�g�q�xc�1��<q��c�q�gx��3�c0cc8�3�c&3�����0c3�c�1�c�1�bq�61�c�3�ct��60v�61�c8�8��1�lc�1�n661�c3�cc�n<q���1��g�0c�q�c��q�c��1�8�1�c�64�1��1�c8�7�1�g�cǧ�1�cv�1���61�� ~f�ިb ��?f{I]<W�G<������>�]�����k͝�u�{�dz{돟X���t,���@��N�\4�T���B�G�[�w�#iԝ���{������b�_���틄z�r[��扣���:�{\�^�=:4�����U��˴ɗSs�LP��0���?QaP|��Œ>�5�BdD퓵�tꘇh�Vܠ]�ݧ�ǗM��n�o�v�}7pvSx3�[xQ"bS.2��
 QǪ^t���W,���� I�I}٠�����Z���e8���,F�h�u��	��哈���[��Gl�sX8Գy#�&��l��"kth#�L�f⋲#n�X�9��/un�{s���;�;F��=��b��R�w�!��[\�����	b&_��+�!��	��>��BlX����������Yw�5�Y�n�����خ�/�]�lېnm�e�{f ���$���u���*�!�\�Yxw�Gj��n�E�/x�3�dS��hf������ǌr����o�ǁ��$�ָl�J��3��nɹ�L׃�pj)������ۯ���3Eg[����	�f�f�׫~�Wi���z�=Y���Ye@����G0ss��f�ĄW����{&3�i�Ì�%�]�$���^snn��G�y((_�UU9OR�LBL\<��P90�%ۜ$�:n����w���^�. p�Jggn����2�R5F��;zs�IL�n;^��+������Ö�I%oV���g�{�.���n!��&̣��<o=���s�f�60y�ñ������9�{��4�b\<u����ȯ�7w_IU5�q6!U��z��L$�8��4��F*	/L��pw���^��Ƴ���'$M)1��7D�w�n��2��&ԯN�q�e��S�1��������q.5)A���܇�5�]�I�Ƿ���ȧt�x�$�D���;����D5�8�X �xX�m��n�'i�w�I:�9�I6���!�{��^��{����3��:�}ݷ�P�󒙄��9)��4�9��s �׃��>�ӂ���|7�rd�����K��������سZuV;��j(rs5 ]w$Sٽ`�{�F��7�5�{�N�Uh��x���;c�۳
�I�O"���ձwL�Jz�����e1(�d�q�����w.`For\��mv����[�^3��_C�]��0�n�C綻of-or���;B��9ٴNZ^���]��L;ڤ�����7pvkr��i0���J��`Wb��x�o_N��)^K#���C���A�W^iע;����j�h�A;f��_js�t�a�6&V
�1�Ο1�x�߬�N�I���z�>نWu����6�]M�c7�t'𻇞�Y �c�r���2���[�����'GٻgpXdj�rMo"��F�#z���x�%�R}�n4o\�lJ��p`P��gC#� s���������{�b���B��H���s��f�k�;��a�+6��qd��ǭ͉p����8����A�o�(3����Kd,�3}�J��29�d�2=}��R��O���1��.�F4�ׁ5Ϻ>9P��=�Wiz�jD�Ǔ��%�9�е�k��s�+��:��,�됙ڃո�ev��zC�бQ9�fj�We�˻@Z;waLv��%|�ñ�N�2.�˥[��ڷO.COv)U�a���E�� ��3H������D\ܦ��S�,X�ܓ+�Z<�����Y���'�0d����[L�v���#{�]zu�;cqn��.�D���ɳ�ʳ�gT��Ke�]�=٩�SL/{7.��c:J���cŮ�d�H�� ��^�`q�#�S٫c��=:wv�Q��V�Kt�0/�a���qt�C	���P6���K�A�ٺ�n��3��z��S ��K�O4Hk���&v �Ŭ;I�Sh6��\�6sBѬ��.iU�k���{/Cg�V\c�J���N���Q�c��w��DC@h|ηO�����
Ž�}\�K�n����C s���7�\H ͘�Z0��Wc�xs--Lr���(]$4�w��gx�%Ǉ=����:4�zX�3V[-0`�7��c�I8�Β�����+�:��L��*�mC���:vI����/(�'$EX���T��9S=��ݏ&7L2�d�&���Y�Ќ�Dg9�M�.h�;��s
r����2�w@�.鈧o6B�Ǣ=����	��Sx��i˨��(c��.ͧ��vMV`��3�ö�q^��l� U�otȷ��9��;XΪb�e�}����Sq�eglũJ��g>U�p2�\��J�t�H��w�n�nn����Qy�jF�k����k�o����޹͕�{�T�X�	�t�[�>��=`��"��t�ʫ��&��5�p��Qt���U��Ճ�NƐS	�&��^�v��aZ!o��]Gchl_ww\����\g���1�,ꓱ�WE+��˴U>��:J��̘	�,��x&���=͘��V�՛e�՝��H�^�^6�<@�8��ۻ�M{B�X"w`ã����FШ;��2J\�/n��v�{��w�=�����׽Gf�%�i鳝qj�-����ڲC�vw!�܉��Go�ۜűZK{Q���n%Ћ�xD����[�������=�E����*L���Hu�	���}�V	1��R{�{�dw��p$���a�s�0�ygZ���#�5p#M�uL3cz��`��+y�d6�:,ѽ�>�+��5x!����#���nɣ4�/1�D� �:Q���jʙ�5ۼw��hjw�9�H^��h]xpx�!&K���:U���7����'x��s�H<�.Ó��@���Qm�[�F�w��c.ͻyI�1�)�r��f���jg�h����w�Ty�8H�51��+��!j
#^^�����n4�7�W9$U,��ܼp��.4�ëKE�U�V.�j�{�K�G+|�>n��f�K�j��&���!�����v��SC��9	��-c��vA�%�GX�{^vp��:�����\ӹ7C{�q-�ϟi|z��'v>����7a9dv��%�H���V�O>��h�r�
�ntG��9��[ ܃!�e�Nܘ�HWڶnF�����>�R�z��卌KV�:�ӻ�`��yƋ٨H�9�gc��j���x�^�	��P�Q���F��7zsS9����Lӛ_=q�����/jYNn��4�/7�-�w��^ف�VFQ3u&۫� ��!�)90�w�p���"��-�Y��|)V���br=S�w->=���ц͝�~L� %Z�7�Le���.�P��n��vw�9*�W* 0a���@9hI<��P�ƃV�>I㷕�˜�:�Y�]�@Ն߶z�K�2���D���e8�z��9��Yb@��w>�~��������tQ����S��qE�j9���.[r拹gE{Fmû#��=��^�i�G�a�{y�}�^����*�v���`�e\�������o�����S}�|�VA�sO ���D���)��i>��)lI�@���N�� 2n���V�V<պD����{*�Dg7���΄�$�v�9u}��K	��A�n�-���.4��v��j"q��f�nK���v>���,���X����Na��7ۺ�C8	U�fP�zv,Io-�.�m5�Ë��P�i�ۭ5�p���Z�v治��،�����;�q�|9$ٙ;�Ν��G[�k+"%\�W]SsS�_A��ͻ9y[9i���;�q���bſl���@Ot���6 $�:�?���}�x͞;���L{����۔/�ǈ���F���UҴ�hߩ��!=3K�v]�1���u�. �s�r\����5X�����;��-Q�V+r�Agn�s�FD�1�:�|wH�0��.n��X\�V�q^��v-�-�աՏ]NE���wUX�ws|�lS�EC:��t'���8��n�����޼��uv�h��/	s��8?�<Q�b��(�D0l4��"T�Qd�;�@^��3�.7iZ�Q�zoe�.��FG�%ǹ���]K㻌f�����mL���r5�|�hr�z,�'��m� q��#u�,�,�ћ��#c�²�w���E�}���}ر����K���Ɔ��e�I�ܐ-�R��b��z��$�qE0���1(;�r�H$���Ҋ��m�|^&\�&!���w3�ȇi�ѕ�Ք)�<�W�wU�b�ɫ	\w��"��54����}1����K��.��L�4�/ww	4��CGQ�5s�a샇q
JK庀X�-����l��b����B-�;��Y�4��$����7x�=��8�C�����}��$j"��m��D�r�5�/��l��;`	��4r�U7(�.���4��;����I(���AV���g����X��v��3��:������q��w͍��1ٺ�0m{sY#�K�<��;`沪�#�wS����Z˽$�����5j�g`�*DW�4�M;���p*%v�.�Y�5�f���zಫ�n�w�9�g�.$�f8�<Kgl��3R�=�³W�G�.>{�9d�7�\��,Ǯ<��4,4�W^Á�F�ou�8�e���5G������^�B�c�x��D�朷$/�ý��q���{Z������urC&�X�2���<{���3mXJ�I������r����G��:�sD����ú�
 ��u.�5Ǡ�l]�p�b����٣UҶ�n��<gwf�E͑���m+s[¶�ķy��,+�����86��Z�l�f�=�@�1�td( k�𚤷\έE�Dk)}��y��v-�'mAof�R���f�'ov64v��f���;���ۗ�{9���+1CRl:�0�3XC��Z� �aa��^��Z�E�����3 �^�]�\�n�����vq|{_�w�2.�+��e��DJ^�-����n��&��q�f�3f{UWl�0����iue�k�j���ǟl��l�,�{������F,m���Ϯ�C������6t~�ϖ��[<Nۚt�C�t暂���OG�`��P�cf�3s�7��(eX����_g��[���$C'V��%I��
Tj,��4�+���?_���m�<�*4HD��ެvn/O�a��qѦUԼ�G��h��i�K����Lp�z×�ih�6HS�E�<�Y�_�9"H�~�Wx���>`̑>�A{�!&8~����Cx���o��rʋ��-pqPt�����J����+���ʺ����<�f��a~:�����O���/��=��ܬ��r�'<{� �aK��1~-¶�1�E�l yv�G��n_+a�!�����;�{��Pl�ϴ�q�[y2ۖgr���� �z쿓}4�q�y�-G|��VI�����}�^����ǫrb~�>�ջ�Y!��g�g�������y?�5�qn��,�,+b�͒�^��os�w�w����Q"]������T�P��o���^�������ً~����|ܔ�|%�$ˣGsi�8��ԯw�2sc$����b�&���T��͒e�O�雥o������
���7�^�=��|����;�cg��o���F&oV��͵u�3;kю<�T�o7q�Xx4��.6Y����2�'ܭ���߹�5�_<���4w�ҷԝ�{��������,�w��M�����FGE�`�
e�ڞҳ��~����k�9��8my+�V��8,�|jOcئ{�����ٳ�N��81��$�.��GGl��ou�w�M�Q��{�+��v��#=y�d�!g�C�uQ"�߶�e���ׄ�fn惂0L|�᝴�3U~D��m!�i_��x;{O�)�������k{l����R��M��Ѹ}�n٫N�5	���N���W�����|a��� �0OW�xyw�n�q�RL�߷p~?�H. ���ԝ=��\�,�>i�I��ِ6RxĆ�ꌹУaz�}6��HQ���
ttgl�}��{gz��>c��ǎ�!�le�#l�	a�k�*q��}��7`{w��o�v�^�3@L���q�.�;���s��;�p�|�ҫ���&Z�{uv{ۼ8P3�h 
|��Th�8h���k��zI���f�����p����;)ę�����{f���"N�_��<��'Ž��y����[���=������}Ѯ�xi^C���5{���ޏs��/z�r�h�����h�k�(�Q�t�wѝ��7ǽ����3���{ok��%�~���=�Ӊ��b�6���ݲ�O^�����<7/ډ�I���ǉ��aN���t�_�V��ރL��##�j��)ݐ�ݞ�#<���v�<Wl3��9~\�嗜��q��5m�s}�O]�����R4q]*�η�F��Q����u)Ei:�Gߴ�d�)Sz������ �2 NY����K!�n�1d����Ѩ�$�紁�#�v����>9����i1;��·q͊-:��Z9~�&{�&l��o��3�!����J�Ws��)^���օ�Dx�⤑�aa�%�r=�r�����Y[�dD�K��W0�3�l����S�?4�B��`B���ϴ�n���0�]缽)�K��iLN��Xj!,վ�_y�n���I��4�z�:bt�Һ�6l���rA��JC�>����?;���O߆n�I�Ҡ��:�T^�ߩE'���=��R�-+�#W��֩E�G�R?'��1��ſ8����7��D|�k�(T��()�iTP�E)hQJ
QZJiT�U)UR��P
��J@R�QF��B�Z)P(J@)ZZ�hQ(P( �ZiD
Q)i)D�A(U(PV�T�i@
E

DJP�P�A)B��V�(ZP
iP�@��P�(U
 F�Z@��(�
J��A�Q
��hU�)D :I:����[/���'�� ��A��~An�+B�;�6m!V�K&�N<+�?�G[)��#k�V[���p�ea 3,}~޶甛K]���3f��"�c�	!�=?f�}����s~!��ېH�4y[�Rx����������<�ma�����(����CH��Q�T�	1!��u��{��4UP9���%�� S��.�&�0���wCp<��v�6٢�Y�	�{�7`ö;NK+i�Xd�Xɑ�s�w;J!\x"�|���˦	ދ&i�_��G�2��"(��~~����bZ��X����7�t��X�4��G�����qe+��>p����o[^�o�f�İ��gý�*�$���L�i��'Ԝ��n��F��Ę���`� ����ː�1�!{N�ˤ3	�0�e$cg,��ln��<�_t�)gb�u��vS��k
�YFX��&�:b�t6���{ѾZ����
0��h��� ,	�	��XƆ�u��hQzMޞ/.$����X�S׭ٺy�[�b``�d��]�Cu�����;�f�FH�³U[�6����W�]-���.`���d�8b��<]���h��c���:0Ř?`L�p!��]�҃ ��\,���5#c�߸>�'��,X�,�4_V/e,�Vwv���(�^嗛��7Mn��w0P6a�H����u����o؜��&��rB0#C�oS%_�bԗݢ��0�v[ӻ����}l��x��7�-X?W{�h䅟 �Z������MBO����ax�����Y,��7���a(�'�a����h!�:���!�ත]&��Iɾ��!<x"�c��b�w7�cm?��>K:o�r�^�d	��=�6�)6�%��G��2���8~�^�$�V96ηl�����J��{�n7׾�>���+�<H��1Y��%�1M��x���G`AG9Zn�C��Ic�>�����9>!�����m��5�c�	!��;����20��8� �2�����#��\$ee&�e�kwRaߦ�4����oLY���}+csX�-��-�6k�>s?�TE?���P>��#�����'���"(��������O����~���_�����yw��I���)$��� f||O�X�b�g�fg�l�W@���E �^�|w�[^�zm� s^�.Lns���y	�^qV���l�,>��g��񦵓J�*.lr3��Y�g���C�7{~���*�"��x�7����;3���g� �}��VtR�l&�S��@�W�6���iO^��O�J�p0
�P������qq�!qS�rޖ+������Ђ��x����l��9�����ܝ�6&3|7u#��vac�K`�	^Į����3P��no������g]
�����}�kָ"��h˗�>�{{+wS�\��y��7|V/7���Y�Չ��3]�J1�\�����t[�N�;"��u>�㛗����I�*�z�z��$����{�m�K����E c|7�WgpO;���v]��/#{#���v�o�� ��}x`G��ɐ��
UŬ���c��y��[�Oj\�B��"�xf_�*.i~>�|��=��O�V��d�<�g���u���>���Ͼ���A�������cJ9�''!�i�&�vֆ����֖��^:뮺�Ӯ���뮺����]u�]u�]u�]u�]~:κ�ǏoN�뮸뮼u�]u�_�]u㮺뮺�:�u�]u���]x뮺뮿N��뮺뎺�ӣ��u�]u�_�G]u�]u�]u��]u��]~?��~?��]u�㣯n�뮸㮺��������]u�]|u����W���b/[aK1>
�����OV�w�.�	=�S��{���9wY
Y�,��W���kFm�7]5�^���fwX���g�G:AϽ�w���< �j�J͘Y9�ٽ:�6�Gyu��6���}�
���78�p<�sD��ef�Qͭ��s�T������n5�Y��d>�ݍ�dZ��P7_�j�;z4*�z��ɻ���u%�����e5|�p����h��j�����8:]oz,�>ʇw�6����}��ɕ��\ž��)L��e���@��W�����'�pf'x&ַ7��A�Ϛ���C��s��g˰��M�<{K�`��fd��{�vhy� �Y�>�uN��=x�%���|�zec}#����>ϐJ9���aM;�l\���]鼀��',�mKQٴ�:�"X�`���㽝N�;�0/m>c��i(�%���ֶH7|�0���s5���9��!���ܧS��yq*q	1ֹp�/�1�H�,vSb�DP�YH�TXR<�|s!�_|���)�i��Y�5��ڵ����̎��>��ᩳ�ٞh���G]	2@yA��j���j.�3
�ի^\6����^�$�f�0�wE�D6� U�{��f[fbԸ�MU�A�P4}�"33���.X���c}VA��b-=a�gN��3�B�	uni5��M�`�4Ľ�#aĂ,�md�����뮽�뮺�뮺�㮺�Ӯ�뮸뮼u�]u�_�]g]u�]u�㣮���Ƿ]u�_u�^�u�]u�]u�^�u�]|u�]zu�]u�u�^�u�]u�]g]u�]u�]gG]u��]u�\tu�]u�]~�u㮺�n��~=��Ǐ����]u�tu�]u�\u�^�������u�]~:�Ӯ�{�џ]u�H�㷪�U]j�L!�2Ӝ��r���W��
��jOd�L0a0�"�\n�JD��MRv E�`�yqZ�F;�b�K (�R�Y��k`��rj 2�|"J��Y���������Oa�>K+�fI�7��DǟfY�aս3o�E앰����b�MxN�n�Tb��p�(��0��E���d����c��]�{w-[�k+$&a��ܗ�X����+���Y�RH�o��eg�\�cתg��[�j��k�+�꠲,���~��h�k�݅P��NDiW:�w���h���o�q}�מ���g-ck�H�b|�f�#>˹#���M|��yDn(�D��Ƞ�v�N�t �p�CyW�'���T�؉V*��12�m��ӱ��f�z��>(p��k#l�y��|�>�?^��wɇ��r�i�۾�����%�����o�}�%��=����.�ۍ��W5�#�~��7��z��{��$1 }rd�7��&+&�ʁ��۟�35�qe�������kt�obX�n�������o��oy�_<3jo�|�b�
��v9+(M����xWI��l�LBb�Y���z�f�����{0%�a�FC�������e��$��>���~���L���m�A�;��>���by瞣P���l���#�v^�&6�i�ש1�TR�%����C[c[[��u�]u��]u׷]u�^�u�]|u�]zu�]u�u׎�뮺����O:뎺�Ӯ�뮾:뮽�뮺�㮺�ۮ�뮾:뮽�뮺�㮺�ۮ���]u�]~�u�]|u�]{u�u�]u�]u�u�]u��_�ǧ����~=�u�_u�u�]u�㮼{{{{{tu�[[[[[[[X��ܐ��@� �E�}J�r��p�?���z��̪e���q�}4=p.7�gvH�˦c�a�{y����%����:K$зz�W�y�gg���^yyn�y9���J�1������,@h�'�oh>��8}�o`~�6��uov�on��a�<��L��03���o����n���h^^�'�^���|��ow�{^�U���R�j�S�uS��r����`�)sl���Q�'<�9�de��k3�(z'�����=�g��p����}�nw8��A���d�o�<��ax�t绱���N�V�i��5�VU��N��n@�|�+
�>���lZ	~����b��,���7�wn�#����K�3s�w{B��M]�6��Ã+`��<�޽q��0y�����J#���.�V��.�N�Vn��)� �h�3�����샼ϣ��}�v�ц��byayp���|�Q��v����G�#G=�0�|}��;��I���_]�rr���|}�$U��j��I��FZ(�5�\�yvIڅ�ga�+��z��]�<�.����x���8뮿g]u�]u���]zu��]u��]u��]u�_u�^�u�]{u�]u��]x�㮺���u�]u�_�]x뮺뮺�:��]u�]u���^:뮺�:�N��N�뮺㣣��뮸뮽:뮽:뮺뎎�뮺��������~?u�^�u׎�뮺��{{{{{u�u�]u�]~>�}7���l���}�|��*�۠!O��߽���W}7u���ǡ���@]��0b��<8�}��_���7�`����:������l>��=2=����Ƨ7�cH��˅�1͙��?��Wp��$U�v�՝�Wrc��z��Y��g�省�`0=cċ5C#5��,m�%�Q���z��v�ĩ}9��ߖ���n�J��p�uWzA=��|��שs�^�w�y�@=���K���1��9����3��v]����]�8�8+�٤h����g��>�s�t���m*u�����k�þ��Ai���x.O���膿q��]>á�����/�ϸPd��^��-7W-įh��� =3>�hw@�����Kc�e񣐝��T3Ǜ�:|��!U�,9�)sImo���ȷ#j���︇����c�c�y�oo�+�����}�j�� �=��6�Q�$�ܵr���K�x�fRU��񶺧d^�gg2���3����<L7��G�]ϰ���3>OfG�!=��:�C�����9�$�A�}�w�p��O�q܉�,�VA��p�`�[%机�]�����ƶ�����뮺뮺�u�u�]u�_�]x뮺믎����뮺믎��n��Ǐu�]u��]u�]u��뮺뮺���u�]u�]u��:뮺뮿N���]u׷]u�_u��]u�]~�u㮺�n���]zu�u�]u����������~:㮺�뮺�뮺�:������뮺��kkkkkS��U;��]^I7�ŹinL��B���ρ�\�����{�T��3�	Y<g��{�{��ԋ}}��U���d��n6���z��,s'��O����3����U��&���.W�1D�	:���a��l],�5A��u��NqV�����K=��A�L���2y�.xN���g�]����`���A�oD� �K��f�m��q`ū��>i<"y/H^ e���p0?0{Ek�aTc�{}���ۉ�2W���0(��}�g�^�md�t��}�?f�È/(��ݧ"����=��������A��{�	z��Ǽ���sw��ӕ!|�ڶ��/R�ȫ����Fޕ�����l�hw��FM�U�D����*�"�j+�c�N��8��^������~��K��m|8wm��t�LQc�6Pp9��s�@j�r��~�Poz����zg}�K�V��M��X��!|PG�w�e�V{��wR��5���x��6�w�]#}�>��:��,ϾnH"�}R����k������������ķp���/�	����C�>��xl^�����[�կXe��\
1��kS;&ֶ����ֶ��.�뮺��G]u�]u�_����뮺��Y�]u�]u�u׎�����Ӯ���G]u�]u�]tu�]u�]u�G]u�]u�]tu�]u�]u�G]u�]|u�]{uѝu�]u�]u�u�]u��]u��]x뮺���~�����~:�~�u㮺�n�뮾=������뮺�ۮ����}��6x4�7�J��D�[c����רu��{5��_eؐ�ި�����=����>��]^���`���6<�ޘ�ı9L�ʔ��yn��s���vs�{��(օa�ݯ���8�S�q`LT� �Sȱ����Ç�ySvx{;��~��ހ��G=�w�ֵY��[�i����zy{o���ͼ{�E�y%�<���h�e�H�ܓ���7���{Wnu�Ӎ���Q�r�f響�i��n�e��������טm���|_����D�Q�b��Z��I�C�0m��۹��������`�Fs��7����=�$^�wV����1�>�B����a%�/�Ǻ�/f
��V��L�~�m��3379i�{�&>ZrK�D�PT�/I��ҝۃ�/zs4�uw���)Ӝ{{�՗��us���x��0���Z3Qױ�s^�e�Br����L`fڄ�Y���x�O��[�f��mNn��}������������q������.�VH�ۺ�9�8]_?	��5d����!c�.�}�BՑ̈�-ΓA��	��>�O����</����K.��\v�(b����z���kJ|�����ܖ�@83I�r��тU�dصA�ܭ��5Iy!�-[t��Ǵ����.��j��u������R�*�`C>�9x���e�E�6L�$�sB�������� ���۫�C�y,�<��3��[�_m����5��*'�	SwӅ�}�yD�w��?,�}��x.s���o��}2�G.3��q6>vpS�z@�q��=}��= ݇N���S�-��������LN)@��m����N�N��{��0�,c�y���Aq�0v�it>�j>��٪�(�K�8��Ł�8Jv)k�T�`�s�h�-�H|�F�.�Z�v=�9�AZ
�XUƝ��n6�.���F����zu]����VV�X�_�.b�U"���SW(����8fek[a���<���6M;��(W��j��#ј���wa�B��� ;�}�ʟ*,��k�c����ż��wsYP� ��{y�THѽ����/{�;Q}w>�����g��/sw�zC�o@�nR���c�p�y�*u�XU�ᒔ�7�|I'��^ر�ʬ߲�}�$��}*��=�z�|�����d�8�y���	�X爫�6��C� �ղG�1�{ٺ���q�V�n�[��m��uዽ���5ո���D�}�3�HQQ?v�j�������҈9��z�熝yf�{�Y<��Ǫ]��;�7}v_I�&s�|�;4i�����@��7�<mc}gdY�g��;�l��
9u
y�45�4���m�݇-�/�9���8t[Hf7ݧ{���;��`��_���n'ų��p�lxi蛣垞���<{1E��|R�-��ɰ�yz%Ŗ4ї��Y|�s��n��8a����r�^��\rp�>`�yx����]��&�7��f�:^�h^��Af\f�ƙ�V́,�> c�<Lt����q���XLهmds�h�k�sj���U������j#��d�I��n�&��esq���Rdx���or���{8��k>�w�{�,�x��]��</{*�cV���4ć�h�����ѻ/���x���r�v��k���6-����e�qf�����sF�R�{�����*;�n�wT��l���־��D�d�sӎ�-������MK+�o��[�+M�����u���voi�m��>��_{��#7�7��m���c=;::aC� ����,?TF �<�(��a��
�����p�/��/����s�|��z���S�� 4;��=f���j��;<��2�����d���JOx�;;���yL����%S����XW{`�)������يn��*�{'٘�g�d.��bh%�c~�*_8���PP���=�dڤ�nF�j>�9s�O�,v��t������-��>5�7q����*�F���&��=��;�74�}ztx|;��k��o��+t�/���_����{S���{w�B�/�lP���dY��ϰ绻d�u	�Q��Ȁ�6�VU]X�T1k�B|�B���4�.]����~6�͙�s:4?9��{G=�����44�����#��¡�hp�R���A�ry�q�!�7g.?���@{Nq��{�3��!�+�槔�i3=ɘ�7zD�.t�u���Gۏ��L?/k~;�S����kg�y�;�]",��npy����1�U����Y�\w�t�n� jFy/O]V���ɳs�嫑�?m��&�n����<���**s���jx�6��Tݼ���Г����_�U�e?ϯ�?O���M�K���������?ͭ`�Mw�v����2��_������__~y��F�����IK���ڐ]H�	C�A3��Hۦ}��,���/����#Ty"Ha���S�,�����D���R�`RZ�8��f-�4ɦ#dfZM%^�5\���91��h鶵�2�0��e�5ʇg64�L��ص������e�-�jM�Me�p۬*���U��/�`�q,֜�c`��kY����ڙ]bdBh�Ή���T�n�9hK[����.��bdH��6<��fh6�A�b��3F��]�63Mҹ:�c+Mb1��,��V
��Z&i2L��
��.&�m�ԩ\�MԴ	�UL���qI�嚘X��7mVl����	Y���D�q(�&�T��[�b6�)L�Âco��׽]�mZU�.�r5���s9�x[n��ctJ�QɁ�#�Q��2�%crLٴu�q�vb��֋l�9�,�Η.ŭ˃^!��q��k�,6���]���h�q*ZY�ӈp�f�j�3�~({�k� +���������3B1��k+���� [ˮmlm52A�ؚ�q3q�eȻ5G�Y��].xB�5���y�qv�A�a��x�Z\2���)a1K,`Z�B$�H�4���f�i���m�4`@V"P�H�!C�8B�Z٦��X���] �H^n��LA�v�4�,*!��ŋsͶ�Ѯ�<	K�9�҄w)-��s`�նQ,"��5�б�Ga��:�:�+I@smM���jZC K�G��2rX0M�SZ�hƑՃ[x�i�[2��A1�ˌɌ2�!��j�34���1��h�I\�@o<2�(��Q��9Fƅ��u���y��eiU��\�i�ѭv�
�˱,cpnºS6f9%���`j�V�+�.6��8[G4��Z�T�p 3i�� ^�c��n����&ØY��m,u�1�ЫK��kt��*�lCm�k(s��:�
l���Ma׶�d�f�Z�њ���h�4v��S^*�V�-[��tnȎ(��4�b���U��e�Gj'.*K)�B�a�m�T6�B�,�ґ�D�@���u�b/4х �+.�M�5�Ma=V)�JA�ښ�&�iu�:Vf=��VXL���[H	��ݜ��ڪ�qQ�!����������l��r���=�uN��Ș�kb��M�R�M�[V�� 뒀E�wT����uL6�4�5,��%�ͣ �wb�B�Q۴�s����9��f1H�m��԰��.�f��p������0��YHG���0���#!]4�Aub���5Y�K�TR�e�#��&����&ejT�h�LLmւ��a4��k��ͳ��0�BV��u��%epp�m�u�!�Ά�j�̷�Y��]���x|O@�00��a��hiw*&ib:k^)�B����]�`m���w;����6�t�;֞|M@��k��m&2A�bn�B�Ye��⸍�R�f�GC�M�VYX<��0�l��CM�6�f%��V� �-ɍk�� jK��' �A�*�lu9n��Թ���h�b�c]��b:��ݴ.�3YD=�ǯ��G��j01�&Hjʸ��6�`�eY���գ4�@5��1�0�]VXB�i��t��u]��X-TH�,�`@�gL�3.�
��]*���؏b��n��Վ��ҩ�\��ep��(�(���-HB<����$b��m�B�&���uɓ+ɯ-fk)4�^r��e����5�M�X�Yd���^�W�]jĥ�"Mc+���̵�n�����0سL^.`XXFˉ�20첵��L򲁒ֶ��ؚ��au���ڀ����-�֎N�ѕpCe�F���MA-�&%9�vty�K�Na&�Ǝ�R�*��K���(2r��l]	x��t1M�Vc��&f�l�Elij�a/*Mk��$��5a^6խ����aKM�%�nl�m�٠�T�A�ϗ��]�{%�u ΀�6+����W<#o8���f���x��$�؆vn���q00�`%�@�����mEvZ�aJcr�p�K)\���\�6�	JMPfFX�Om����D�5�XJ��%�e�l�F]�� T	M�m�� ��ۗ[�5��.(`��1c-�£Ś�\P�U�RLM���jl�$6�yhˬkR�D,y��͠�hl��4�ѡ�`������C�[��ӌ�FY��h���%�°�kK�$e�m[ō��������4�δQ	��)m5e#L6���-�����i�XB콊A6v�	4-]���ڑ
��m�b�H0���4�(*�.��a����G$����N͖S������mJF��]MF������k���5�P��\�DulИ.��+�]����)��7X��v�"$�r�n�kF�R��!����t�crf�Er�[)3v�ubYv�m�-�I�e�2�6*�d�jQ��GI���p�"��Cm.��&�kX�q���F��K�vݳ�&l)��7��\�@�q���	e�m�1�q�р��X�`�9�8r�l��w/^��-5�C�lB6�*�Id]��@ݑ��sm+4��b�cky�K��	`՚��43dhL�M�4ĵm��%#�7d����MM-3V�Y��n�cJf�R����7c�<���4u�0ܻ6&\�3�6��*�B�iXSHm��q���.��MlD��1���q^R�r]H-3�5v����lum.�3
����6��Q!W#1�,�XAɶ�54X^�S�
٣tl�����l%a��Y^`�q�5ViB1+&�-ann-�[��S�1�GFk�sRd����,d-%p�(�0���-��JgF����:ŕ�9�Pu�ˁ3ey2J3��v�ZcN�`�U�ڥZ���hUjdpѦf�mlHEo5u�l��"�Y�*`�Hm���h�]a,�-���خʗgl�6`f�]��W�jIL���G�
�E��B�L��VWU�$�Ͷ����Vgm 2�,ɠ��X�u�mF�R�:��KGc&Qw�g�Ƕ�Qbn��l-�L�����R�S]�$#��4u�چ*%��h�5b�ct�hX������֣��,(u�GGV��As���Ò�(�5�C�vpJ�vњm.�k��f��l��֛im��Z���t�J����"͌Zl�e�����g$����܊JBeҕe�c�f��.	�����v�l5YIu[�� n�Aԭ���ݒ�cpҫP�2�]� ��9[.����l�ô��mK�� mb�Nt%)�kJ�M��IzZ�������u�� �-�4\�,&201��������n�z�R.tv�B���Ƭ@V���m�j�����6�45�u�]-+�B7�c�˴��i	�k�y0�.��t[�XB�sF�hf,�bk�Ñz�oWX�!����ƈ��e�ԀU�!�m3)[�8��V^���Fb�.�Fi�BlM����^CDu�.���j�n7U�m ��[-̶�aK���Ŗ�3ErKc�%����f�M6�/lY���i��4N��3Xe-u���W�e�1)pY��E&�٪YX!�Ҽ ���n�ؖ��]2��y�x��G��`�el
�\�G8�� S`�Ե�Z�˱�U�šV��ZR;��-�,�R���v�VdPق7��;�SX�r0��ƒ����M^dѹ�a�#M�KīT�4���	�2C�ї+�fp�c1)]ph�!��f+l��X��4���Jl�Ʋ�^Ħ�&z�)K�fk@�ei(r�aF-i1y����4m���Li�h�����Q����V������&ue�2��L�t.��)�Z�њj+[qr�R�­�U%`���M������
gl��Gmbۦb��8e-b�F�Xl8mΎ���٢ՅRg!.�b犰�������
��ݖ�p�WL�r�8���gjh+l2�ɳD%��P�o��zI;!�t�����rϐ��� � sVo}Jp���o#��in�k6���o;C_�x}%�z/���{�oC1�2"Fb2�%��0'5p�OV(y��LѺ�Z��	Z̑�
YhHX'ƩhYњRژ��>���w�f�ގ�����M	1� ���b!��[d���G�A)!
^�׀�*����3)U�AVT�V�j�x����,�jvnnjjjzN�'�����hc��X:����U�PD�	�dU����
Z$R�	*@+ (Zذ"�%�����k-��YB\� R(�Y6��U����R�
y*P
g�O\~����G��׌�}}�*���hR9`E!%H�$W�djUd�I31 �$RJ��22o�Y�u���$OC�+� �ԨJ�*B�H��
�B,(�ӊ�H�(X���BВ�9x���(��3%��NM��MMO���},e'���"8�ٔ�[�m�M�n�O����ab9J�EF���t���IE�LC&K79;77555>'������ϓ����y��У�wj��*�M& ��7�0�cG��Qq�j�����O��ssSSS�v{=�L�ɑ�g�~��Z
Ue
�2���J���V(�c�U-��,�����������^=<g篭1`5+""V��R���MTӤ��)B�����;t�"ʪ̴��mCĢ�m�����"*��ʂ��mm�ֲbu1q�2�]��U��e��,T^��$TE�F#(���k(�R��`���j��j�pe����%�No���D̺{J�9�հ`ͭT�&���ˈUM�#�%Zch�tYu�Y��"�ˇ��Eڶ�W1�1��r�Tl�
K��WXiI��h��.`A!u�O˷\�B��hښ�����
Da43Re+�n$J۳c-�c���ы,�V�Mī�嵰7E��b8�&�[�����q��B����uvT��j��)��q+s�#���5 ��m�+,���]Y�Y��n��GT����Z
p�l�
B�
��d)k�]���یhgWK-Cj۠R6��[Ԏ�Q��N��X������6mԖKV7S�+�aB���(͂�5�˶��F-FZb#�`4��f�%҆eݳ�m��=�v.��W0��^sR\�0�K���2��U�v��[�⑗k��uU,���H��"EH�[`j��ʷ�V��ƪ�aI����c�x��k`u�]en�!C7-�(�,ʫm%�M7Q��ԉa�j��&e�M�m[x�3L-Ź�tv�bד�Z��,3�a�Q.Ν�ב��t��f\�rv�K�D��`4m�8�Ss#e���h�l�:��c;׀٪0b�'[[C0��V5V���Z�݈�КTYMM+1�Ke���C3T1¼Ҧ����F��bV`�
�%jS\�*�
��s��ܣlKmԡ�hF-����8�R.�+�ny�8ܙjap]V�K&Hٮ,Υun�)ac�n��#sic6�@<��nٱ������s�y��b613vV���[��Xݪfc��:����!�'o�亊��i��B��Q
B��(ڔ�)��m�H�qN ��[YmcJ��#-m�-e�[*ج)^4���%�-yW���8������-E�T�IlaH���2��e�YbE"5�d#��-����_�>V�ܬ�gB�ia]�\ܰ6IWAZ��M��=��/��a*���}�4�޿���f��:�-m�D=&��>�P&ty���0�7�?{�o��IK}���8�\�}�������+���݌澻�,���ε;ë޸�z�s"��V�L�y���e�ߖ�8�0T��,����|&�U���|Q�kj��M�e�Wb���m�,�P�P@`�]�hxhv�]�P5�����̌���OBϩ�4��C�E�v��}��#�6�M�a�������}��W��9���ms����ᬻvwYC��r����-�@{2��=7��޼�ü�bokfz�T�ϼg�-�g���$���?/�}�ym^�x���J�/��p�$�䍓:Y�4w��p��f��f��.�q�U�9T�����D���0�T�<!$c��>�y%�[���ִ�r�$�|g�B�S,(L�=; &��g��G_�a��j+_�|rL��Ӄrs.��Y�ֻ����{7��;�jj�
�^�H�ǆ�{%��-얶���z�+I2g��Y���l����1o*��{��]�VzؙM33 9��T�m;��V��=��\�P&�a�V<8�֪�2�Vlgl���c`E4@���
�V~?h=�b��շ���R��G�k���nnxN[ǎ�U���PH$5S��6bH����r�w,��3ڡ�w<��p'��/R�槭��
	j�v�ߣ�/���3���i���}��!3n?�&���ڻ¶x����1$����2�[����Fq'�淏�:x�b>�=����O�N$��'9�o{���[���E�S)���5�S���y��pyڈXp}��,���:�~�����,���8Muc�yf�c�yq@pA���TI�\���
cL;@�����fA���5�gEW����VFN$�M,X_����S����ٺk]�nLm6�փn�z���D�1$m��$�#54βgaE<罱�u����ll�C���hA���WC,��ؘU 6���62�'Qb�ݎS�ݹJ}5�O���	1��f�[y��= Sӛ$i�!�Yؘ���ٙ7<cך1�w|%�M��BL�ƪq39Z�~�zgэ�&��V濓�x��Vx��[Nz~��ߡ��M���)�|=�0��v%<_KxZ� y�O�}�W}�=���pHݼ��Rn���{����RF� ��%��h�`���2`�h�0O �78S%����S��0�R��*�C�d�!��"U>F����YE�,���g������P��<_؃��x*c�߯��>�����a��[ ��gh���L�m�dPxt`$�MS2�)q�`}�������I8lH[�������� ��aUL�ʵ���i��P��$!��ӈ�(���;���k�o4��j���&pˢA�E�q3�Dσ��|Ȼ�z��J����^�Z��a��!&d	��I�M?��<��iED�`z�`Ǎ��b"�S��>�i�L��m4�S9&��6<7ލ���������u�՚�/<��$���2όAȗ��"��`/(�א}լ@�
f��Áw��^�f�O~-1��<Lh,�ڝ�H3�����p�.E��Yoq}�n�y��H���0b]�|�zY�@�Cu�$�Bl�;�$����2��r�m��6�+�4���ui4LBl��2�Y�#-��k5��.)�H�;f[Vi�-�-sB�#e#�@K�ݨ�e)VlҤu�b0@�%vf�glfSRl�W]�m�e�
�U��K���X�X�5��������4�K)5�q��6�QU�C4�q�e<�����t������
Y�m�Q�uj�v#Ɗ�Vٙ`�)c4�<��>ig�,��f�o���x ��>�ɟ^N	̕�hj�v��~������N=�b=1�v�p[ֶ�ԟ���W��F�t��b��b��(�I��,Y�T��)�=�Okrϕ�y��z�]^!�&�*5Q0��i����{@�ʝg>TD�3�x�:����<4 �l�nV�]TxO�=���i˘>��'�����O�q[�V�٧��w��4�3�- P�k3�&#|��3퀼�G��������u����u΃\W<�X�n����	�� >�8���=Y#;H
��/fz=�P��������e����{x�RʲP(�
�[yʩ>$�)Krcm��#�����L@��F���돽}�bN��׾ߺ��^q~���4��Y@I�ۖ-����wI��>xS��vs;`*�%�_Ȑ�K�Ijd���ibf�=/P�r�W���hvT_��Kd1h� �7p�O�**��I��Θ�!����T'�f��0�N��`���y�����҉���p.顢��;�����f<�vɜ����r�i^�z�&�C݊n^�ًxq9c(eԟ~�>�>���c\�X:���Z$e�u��i�M��������g�<�x=�~��o���-7�=x�CvZ�OTH4]�j��q1���v����S쿃��MמM��2YU�jM��T��Fa���T�������O��n�C�w���y�r������ԑ�������y����E�p��w��y��"�:OI�IԖ��_9�~v��Z�5N����i({r�gM:�y@���OJ�.A��稿�44QpNUSJ�>��;�A� c
 �ֵݼ�X'e�/fny�O���Mg��q	"���E�wt�$�`�@s1�dL�@w��G��A�5��`[�[2�hgm�D�:1���S@X�C9d`�k�V��,�:dʵ�j����I�g��0��^�!7��ԵFߴ���#u��;Yy1/~e��W �<�����e�"�	���d�{Z� �e�d)����k:"����M?�W�����O�Y�Zv�x��B��9�]��K�S�U���[�*3�Y��^b��V�y	G��11���/|�0�'ě�法��i��f�N{D��t"�k;��ȟHۗ�����w͟YɄ
8 b@^���-,K��dg�����y�p)l�kz����➳�H�Y��3�*�'�r���|Ai<4�GD&&��g� �d���v��1#B���׳��6�rj�ir5�@�"�Y�k�[��ץ�>�U��ܑ���ޫ�r!��$	^j@P�"��N��}����=�|!���?�#���$��3�5߽���Ș� �S��^e�f"�NJ�xk��[����g�硌Jo7�	t�i��&v��S�J��޶������SU�}��;��<#ڄ�P��[�˥i�$9$�/��T��}���v������c&m���M�V{�/O�2��k��jL���3㙞��R���/E�۹5~���\���v=��kN�f��;7y�J��C�X����&o�&��0��/ű���Űcb�y٣z�Q�HYe�^ZXJݵ�&jB���o=�2Y��9a5�O*�ʚ`sLT%#��К���@-\� ���%�m��7Z2�Y���Z8eA�(f�s\�,�1�6���v��\A��K�!`��:82�T��1���3VhE���5́X͊�I��$"Fb�j]a�2ܮ���Р�f�����b�1�#�[TH��ɓia%�i�>g��f�1���X�!ue6TT5e�3��L2\1��0��#Pk0�e�'j��7�b��s��N��oF�үzf|�N�X;h��M��.���5Ӵ����[:<�sS;e�SVv�U���çJRC�H	i�����a��@����2��qX>�E�'�5����qWR	]В]����<�i �]�h-���'ўsU~���h��0�Ɇ7n�7�*2p���v����!�ܶ*v@�Nz����՗����E���_��*�eׇ�	��<A���]e�jDwi�j��@ѤZ�P��P9��wy�ϼ�vv3�YJ��#{in�#8(��R�g�L4M~E1j2���lV��{�Ix�ڷ���~Ú��C;xn��X�8�!�S�i�{������m�b��"�[��<_x/h�~�Fw�}��ŀeo45�z�]F�MU�i�+X׋U���q�v�+PX��R]M�i���b�sI�{�(��D�k���׬�b#�ə��}f��+�>��j�i����ƚ��j�.�V��<��xU���S��m�z�; '0W�3�-T�}��wY��sO�����U~�}씦K9��T"^<w�=����D	!�v�gJ��[�y����>������њK��v+6�d��0�-�o��������w�;�U�Ǖ��9�����wA{�=t���K\�1V�"Z�9�zG�M�kuګ�u��3�oH �֛m]�����Ԡ5؛�1�*���&`�� �����N����n�;���/V�ee���1J�Z�KB��0��&����x�*r�=�7L[��8x���}�"�W�o��j9�t�a����]q2ߋ�<�5�m��r��,�ycS;t�]٬ߛ�ow�o�R��©����bs�C��Pk�Վڙl�X!{}�IX�qc\�ݫ� �����ә2r��x��yV{������ܾ!��rB�y�W��̓�L탇�Ñ��g{@S5�Q�g�[��u�[����4�W^�����~<�wv���f�L����7�<�P�Em�f\�|6o������5yo�C}��8�{���RЛ�_�t���2q|��w�v\�=���{%k�!����ױ�{�d=������Q�҃�zbe�Y�A�����W���A���g����G;�``u�f��}�t�t��щR���.��@���@F#����>t�z+p@=�/�7�����Ơ
��9����Q�ʇ��ٶ�>�g'BW�x�}�7���Ors/���4c3�_x�t����;=���[� ��%�~�����2gg��4��.������l9*�w�^˟������@�8N�g�b'O_P(�8�" g�#�<�����i��x2_s�8[��6���W�2FS���c�R!�Y1���>�혆j�`y���1�8cP}�����$ўˉ2��Wr�䫲����<�`�7JѭQd�(��\�e�i�(֊�pj����Z��f*k)�,fM̝����������XϦF3����W-W�
��r������L�f�!I<zzq�������}~>�g��>��N�X"?!�&5F,Qh�2؊8㊫m��Z�kKǄE���Oo�O�>>>=����_^3gџx��iĞ�J1ADDEwz��1U���Z^�
�(�Oǧ������G]}x�Y��ȯ�`Q��) ��qkb'�j�V�3DTAf�f��8�oo��������}h)����YU��q�(iU1���9��������8����O���,�3ߏ������J�Z��5*5�Kl�f���
*6��QY�X\j��n��YKl�bF#��Ƣ��l��*���TDթ4��(\�X'JD�Y��.����Pkb�R[(-BT0��4KZ{�yf��-�V<Jŀ��*��q�J�R��3L̢֬�v�)PAZɀ�5J��_�]!U��5�LULj
��^�mm��f�bF$c1�$c3c���MT�<�~�U~�0����� ����2�R���f`�C��hd���������|��5������-D2*�}0��,�#��L� �`=~��v�,Hg^�p�k&��#FD23^^ǌ�!�q��tם�U��LXsF��i_#�]�'=���Dǽ��t0�� p���u��Ҭsc��a��B��;��9'Ͼ�����ZU%��8u��`��d��У�v,�X*�_7F���,q�#�)4!�(-�y�{�UM���> p,*:=�4�./�&���C"�ܰ���6��%�p�Dw�Ԉ�f �F �<Z\1-�=U��f���~�@pvA�P�� �F��`��)�O����1.�����s3p���C�)����`��DT�K����`k�G��
|&/�~/XX��Xvh��s =�,����)�@C;��앐i�H
b�Hlg
���fp�3ڻ���y��b�<�-ɂfw=r���^�Z�$����+�z���Ԅz|Z-쉻��Ug�c4k�{|�ô�����l,�IOs�V�w}���	�1� _��n�R�����߻}m�n����jJ��,�	��d���ҢƳ��b��&��Šw��d�'�c�%9�LChS��a���х_��Y �`!��N��?_p���X�f�Me�Ƌ��Ҭs-U�4u�6���0�2������Xd������2�V���T�4�X��WV��y<$>dߔF��Fr�Q��Q��l;j�0���߶��J��r Gրu����p��A�@U� ��se��� n����M�v��C�i�{� o��!�G���a�S�v�\��;���3S�� �l��3�.�1 x� #Y0��؁l�>�ݦ��"��@Z� ]�v�n���8�����Sq`A�sVֳ��{�Q�%��fFn&3�)�p7�M��P�)��eH���u:�`y�+�^�u�T{���JaÙ�@��6��G�4��v��zQ�x"�f�*��E�����fw��g�재���t>d�t�&+������v�~}{C�/���s�|�A�LE�1 ��Sؙy�٧��Ғ�#�FR�\R,"���:ٙ���Q����2����$c?�e��ՙJ�'��Au���9�KyiK�l�&e�2X��qN)��ڕ4!��JV��Ìn�`;e ��Zk�c�3�m�d��d.4[P���sǔ�i*jțV@�C��E�:��٫�61�XV
�G��,",��5�BV�kl���V֖ZL�WaKK/638�u�>�~�����Jk��4���-e�3�K	�V��Tѥ5����{hd��!}��;ݘ����N�������f�@q`����\��O=��,}�2�,/h\�i2YC��0@���?~�Y���ł)�C� �~�g�un�@�"�n��!w�C飾}���L����E<�v��A�^I�$�0,qۡ�di�J��``�;�}��XV���ٞǹ��<�ǁa�����~fC�I����C��b���3��]�g"�o"Á؁�y�(b���Xa��ݙQ��}w�3Sc��v-�y�1k+:�������P�CO?PÛ�Z�P�!�.<`��HV0X+��ءuK�v�����j���$��[���ibRŨ��L�hd��5��	�Hg�I(����G��en`!.�.�`M�^,^բ��bJ���V~I���O�{^�@�CX�������`={/W�����O0�#>��`-c����HJ��r���oͨ�/�0�$0��GaOZ#�30��r�6I}F�W���2<r���H<����l�(N�g�;ϴ=ܻ,�g&��z|�u�zo鑜e����3FX�f���i��;!��k۱�b�ܵ߀�\� 9��Y����Z�{�G�pnr�x�ҋ,�/���v}D:�ۇ�<'�O�	G{�=��燘ߋs�
kAذ�!���&>mMA��3�Jy;�/ػ;˟J^R{3¡>d=J��SQ���߶�w���W<D�Qh9��x<����x�@�׏,`c!pY6B:�1U�����w,S�k	�4M�r=4��������'��/n�Ʃ9�"m^���'�R���LJ��,F��K}�hP��4le[0��9��� jMu�3��4����x�0��w��"__X�!v��{�[��Г�Ƶ0���)�zr{e_�����vv;����*"�܂@�NAU�|��j;�T�{����oZ�Ξ ��J�
�:4{�ɰ������2Y���,E�=�$�B��F��ٮ�["����;��_����Im����'���Vn�c:����R⛗?�,��y��5�u����H�X����Ȳ`Y1d ����{蹥������_�h߯#�����{�ڕ[��NJ*bx��V&�5J��$��SYB4z��[��O�'��pp@.փ�b�=�x>N7�݈z��amcv��Ո�Aq-
��V�3΢�t�T���=_D��-��L��,�̊A�K�_Uz������" �p����t�^�1�Ns���)�\�����%5ɝ��z~O}^�g�a�čTň�%�$Rg��>��|�c����;��j��=j4�Yy��e8����yIH��M̂�Lϵ½�a�����;S.<B���*���(��Z�H��kI�42e��ޥ��=��'"����3�]�Gt3��t��^��Ԑ�[�G��]���Mmxi�Ih8 ָp��Z�b.�V�Y����.z4�#����0^�9c�6CP�3��ϣ_ݐ�b\|���cU�u���J��r	P�ͅM��WC��~������uY���L�;++�ӐK�F9�`}�G1����[(s>k�O���2�VX�2�{ᩄ�B��`,Y��?���;�3�5�ssm#HXc�E;Q
v�3he݀���xJ��u�\<����Ŭ�`Ey`DӰ{b,�cou��be����\�x-�h�����J�
�3��X�c[]�aWΙ�D�]�H��u��� $��A5I�O����ɝ������>y��H̔ =�!��]�)��G�x��/|�٫�U�he,];�#P�.�!n�]�	��]���g��-M��1n\�:�h&1�S8��%��8 ͻQ�B*�.P��>��:��څ\*�,a���1r8�����o���m*�M��i�~/��jRf`VJ�Xx����I�{2��}�ײ�w����{���;,�8�Q������i�o�k��߳�8��>L��{q��W�����d	��Py,�Ls9�Fg��:���|�.����^����z��v˔{U��L�BU�-3���L^`/�z5�qN�E�<;G�����ك�23V#4E�~#/��z�B���Dp.ō%b�Mn����������1�N,%���B�R0�"T"�<�E�n��:h���Hfi[3ȃ�0�X�(%8mD,�Ve���f�j�X��hל�u�T��lQ,Ri1��[��7�g�2�eIR%�Us5�XZ�y��Bk���J:+Y����m�fVu <2A�9v4��yu!�E*˕n���$��,�Uu�m�Լ�h��V�.�q>~��ܻ$�t43.�Fl�B۝K�[6�vi�5rK?�)�B�>� �()�6B"�9;�=]��k�W4�8��Q����oiA�p�g]��=�F�"��rEy�yy�X3I��~̓���u��U�+=�ՈSb����v)�l���=@�I���458���Q	���B�B&����N˼A��Y|!��#��>�D�L��V��*ӀA��Fz�/�cvP|d�ñ��S��>�U�5��Ã5��2TY�q����#d�g�R�4�N�	|Y0Xu
��Z�b�P����0[(N纤�o�q�}L|x�RڵÚ(���v
_���X��PL-�y�z�&��u]/����g��Z1M�&T4�h�)��+�)�aMc�tbBϟ�����N�ءHK�V��yn���/�f&�	��]���D2/1����Yd�2
��RI{�N�=ޙ��w�ُW\�3��y�s�_��}�1 ���N(�Ll�_�_ �iU���������28��q)��O��C�OH�(���!��GVIm������=J��}��`��}��=f��w��&�,FS�%زYyX�2����i��A{� �kP-iI�Zǘ�RX��i��/Ku���k�=���"Y����8��5�
^oɓ1�0̔���y�����}�Mj���W��>DD\k�i�u��O�;��̐Z���W���w�'����{���Z���ܸ=�b\84G�2�t�3
!�0�A���o�v�OY��Ƽ�؈��r[��*�0�=���`�{�}$;�N�E�x�����,�V#�e�iubk�#�4�3�I���l��+���/���N�~��T��W��ƽ�c��v����{͉�L{��I�����Ě�rC�'9L����1�f�}gK0��I G���D���r�v�F�Q[�h�~~ɇ��8�}�ݵ�8�v�O��?N������£|�0�cos$آ�
!|����OK�wB���ǟxזɯO�e�L'�����3�{˯`+G㽦���(���)��?�����i��ʭ���L=a�n���{s��5�>Qa�a�a�a�@<��b�g����N٪����	��C;��67�!�U�F��`���t_.[!�ɖH�b��ܸ3߽������<x�^��A���Fz���wb���*Yi�����niu��טnj'l@;F8rV]���wCZX�M�O}������&��\]��rA�$1�L��ҭ�uD]�����	ܤ��c�8�O�O�&1��R��܋NթH��
Lm2gz|O��iгJ�v�Q�Uك}���'��w^w&���ؿPu=>�D1m�Ꚍ���;��w)�*�{)��1E羳�&��=�.���F�=�D�W�����/s�ݜ��n�p��P��w%�a��ҧy����i&[� �W��y���3u9$�w@Aݒ-e���=�V�U��X��td<�� � �S�H�d�L��ӹ,}�A��y��=
���FrrA�9ҏ2�%�����=��z�Wp4�/&pH%���3��&�/s�חJ7��?�"�&��DZ�@ƾ��<�z��[Ry]�|w=���&�Hר���Z����f�b�HdR ��80�r��P��%
Q��}�bj�����ɖ0{g;J?����8��#X�*��쯷�~s7u��ˋ�'��O��9�����J>F��ž�z�N�#��ז~ˠk��]��o_��{p�f��͛V偒��"�VL���SJ��Xh~1y*ꕂw��Ns0T�#w�~�#�=��|z�k{�ڏW��v�ô��D:�~ {>�ٺ/�s���H[Q��������{����HD�;8���[]'��sN���me�n`3��U1�� ������wo �5��<��{rny�����m�������ম��ǃ�M��Q5��uر�e�p�xz�-u�<�6����S�7�ŉ��"q�U�����W	|�w�;X{g�GՇ��G�s��+�����17-^Z���f��":��s�z�g^���n�q�����X�&��e�6� �j�Y��&�M���b�u��gut�����Jn���ٓ���f��Ď�q�&��Ͻ컴������pz71��=��O��9|VvX�=���/2A�Ot�Ǔ���]�m]�_�5��5λ�uz�SՏh96�5N�;4����׻4vš����:�`O3�t�>�y�^\S��R}�Mx�USy�t���bvg��?
_>�ZM����0��,V
���Ӝ'W����>�qڟ��ɺ��������=G���a螣ą}7����W������-	�^�U$�>t��xm�:��*��(�Y��M���q�r�&mb�;�=zz,�/p5��˳�cg�9rল��h˷C��,�x#�J���x�-�������q��l�[V����5�+��̏���[�(�O{���j~2���Rg�:�H�]����j�}}Xx�8�����I��\�A<�-5P�m��}��x��6��o}���Pu�\�jo�:c�~(��������L�@�����L'���#޷���t�����i>]���!��q�]�/��'��!�s!�����At������43x��BYw]�L+A�����XX)��W���?9��~��kS(�zg�����yn�L��myr� {�9pW�;y������ּ�k�1�,�WP���FX�g+����i���K���HԳZؼ�������/�ߏ�Iy��Ŕ�1�ݛ]0~㑲
CF�(`�!�����|�y[OT{	gQ�ɍ�1�ߦ�w硝�9��}`h�#n�-f����	�.���X�����������wJ����P%�;JB�t'�~KY坱笻�H%HEl�X�CAh3��(:��m�b���?BwᯁÝ��:�nY�5�JQe��,A��kw,���k}�Ϳ;��S�	!<�� ���P��S��n�D��0�>�\k~8���3FcSM��Q��C��{�$��XW� �
�C=ֱ��u�D"�Z�e�c-4�6՞����q���������Y߁zĬ�,�MZ�?Y*,i�aU��!Z�QMY]���{qǷ�q�������ǎ���f"q9)E{;�d<�Yk�A���|L�����W}t�]�ǧ�׷q�|}]}x�g��O��`�me���}J���bQU"��X"��0E�h�7�\�<$�~��q�|~���},��c>��4G��#��¢���H�\5h���'-+<|}{~�q�|t}u��ǎ��~K�̦�I�A��o�dQE#Ab�_IwlR�J2�x�>=��:�>?C��>�g�O�jW�+m�X�����ΰ��C�q�d�0���R�m+65��@Y�5f���p7hi]�UD�l��1q�*TD�%��kN�H��a�����2خYTI�����|�CAIMi�0S{�3MQ�db�yh*ŋ�^ۋ�!��7��w�R��6�#7)�M& u�ܫ���4)�6��s��a�M/����lY�&��e*9M!fS�B I�,ѵŕnm�l���XJ#oZe�4"�\]
�.�8�*����l�\�HM�2͍�҉D���V��.M����9��,u�i���3�B��S�%�W�(nz뗆D-,Q���[`�r�d���jD�奩Jb��MnM�f�Ptu�λn7b%����H.�&qaln����scۍc���Ź���q6�5���Y[k3�У� M���99�-��#H'U��g��O_�F"�l�[v�Łv	{"g6�@G,L�F�V�Z�9���ai�hX���u33��1exݩ\� �� ݴB�+.�y�������#u��<B;��jX�L�δ Yl̼�m9F(T��P��a��rƵ�s��(7�m�n+�2�4�֌%a1�⛨%�F�\¡�*XЄ�-h��ʰe�Y�i����Hde�[Hݠ�	2;m��30��3I�*�++��8ٕR��֙��M���s0k�3en�u�fi,��P�v��k��F�J<CF��YqEP��i�H��b��ba2MÜ�帲��h�Q�l��R����0�K��'b-)�j�Dp�$ �&ml����0.i��AJB�=l|�3u���t415ؤ�6�r΀p����k�A�ʦ����7a+��:�P.�kJ!�ik-�Y��u�Q-�m-tZܘ�˚���vK�	An�Q��1[��7-5P�Q�U�#�\�A!���==��yXl��K)7w[�S�(E��3�O����� �2��� 0�@� d RO���-̵s�U���Í� �j��jŶ�S	,�hU�����vh�x�3�`���S�y5�2)��`�f��֌Uv3F��.ٖ#�.ìa1\��4���(\B�6��p˚�Z&(�94CM����ִ�ĺTX�]�f�l���(]��2�ڙ��1�XRh樝�9�������UF�I��\-�-2`۔��n93.H��ֳ1����O7r?L��e+��"���*O4;���\U���ǫ�5߼��d�O{�R��o��6#���j-�]���>׻}|���$H�Zb��Z
 ������x+�����ǩ�H���{[7*��!�Hk$��%��h�<�D~�4�|���X�Z�#�=o��U��������xq������Q��'�d�Ǎl�D��=��2�E��mwrA:B�a����N�Cս����$Ԙ��;�}�z6�zD�k��LI#���6�;�D�(mܒ�_����6&,�S�}����x+���k�2D��w$;  ̂�9j�<�f�>���#�%������í�|�={�����Ψ2�H�]ekn.��݇5�sWI��>(���qP�MU8����|�=f�X��=�Y���W�'ȃ�Uk�iC���k�x$v\���X���}���Oz��ry��W=�g[p��b��7�}��k��u{o"K�'o{�6�km�>��~�nRU���Z�;�E�yml���Z���C��D�� �Ay��8� �A!�CB�Z�G����9���=)�W���u}�����!�����84GS�>E���8ע�@��.ó� �ÖN��.^�G���;�#s��c��RWY��8s$z�'bC0:B$L3�v��g�$�#�|揬z��c/|#q�%��y�x��كk�^�9�������a������D��)�f��Y����3<���[F�d#�~8Y̲��������<�]៷6��f����b<�� �;Yv-B�Bh�xt-Q�� 9I�D��Qw���U��(f-��S9�ܸ&mU"�ٷ�܂?����S8@�8pEYd$0;�����~�z�VH��;���~��%�cw' ���٬���M�ϾQ��H�yLa���3�!�gV�46��L�u�}�^]��/u�;��(�7s:b�� ���]�,Wa��`��@b���%;���ک��F�$�ʺ�9q�2�l?{���l��C���E�_�����\�u�m�.�kn���g}8|�m�t=@�����K�ɺ�v����#K9X d�9��.I$� �" �R2HJA��	8u��!*�03����|8]U��S�$V���dH�p�]ă�x�L�����F�S�8pE�A�+���p����p`7��Y1�	(Pz���Ÿ���9�6���n�Qbd��ѯ
�F�]oD�V��P�8~���ݎ�w]�XW�9VI.��k4�g���@�A��2l�h<�d3��r��c�>M��:�.�n��6ڌ����P�l)XX�S3>����)7��g�-T�i��,� U�����Y���ѩ����eކ�B#�a��>؍�w���Nrh��_)Sj���;
�]-E;�lH3�w�}�:�V;x�!�M̩�2�ȲɌ���id0g*)��U�<'�a↛0�2�(*�ܘr��{�:p�w���?eNL|&ivwd<]ךw��d�X;Sap䚷g�i�PH/T��ݙ�]��t��Ej��-��p� =
Ai��*yW{���J�xx�$���ٱ��7�?<�������O�C�Nc��������'�trY���~�e����v��gA���!�D�o��+{��5���}�3� O�2$ R2)�G�(��81��t@�@ D�4(P� O��ٲ+cO|Ѣ�w��ѣ�X���c�����7Y� ��2���}��g=���d��P�Ŷ��s�',b�ܵ~>�O>��� �:��k�M���%�ֻ[�Ē��Փ	cf�4����f���#5������#�R�Ze��)��sƣ�w���w^i�rc�z�/@���4��S�o0�Ra�C]�o����X>�"e�w��R]���T'�%���RsLXfJr%FwO�U*͑���,B�A؈�M�R��;���_.O	���#��l���w��"��0�/�_!��B���݇N3Sz::�������7W�iòL�RslP5i��lm�����ss�փ��A2��0x���������>C��4�<1Lt�X;�wuV��!y�B���ж�W*X�nS�`셻"f�7&�W�I�Wq�:��T�7�ǈ�L��rN�&0�Q T8��pW����F�C����i�
��~�!�����rػ��o�Q��%�;�'���3�+\�CŐ��=G��Z�#�[�5.Y�%.8ֺ6v���{XF�/��0�N]�]S�WZ˗5���D�����y�pe@��$�H�� ��!2�����VXFim+t������di\�%�U��0���4�pjd��l�6�3�(�63W:�B�He��i�Ria��LE���pɐˡiM��.�4��6@��q�������/�թU�K�ע��vmp�in�H[UB�R8e�N-v\b�Æ���U�[
\���}��d��@��#L�0Wd�rͦ7j�^��������=��N$�7�����V�O����D����\�����nwn���,��_=���h�2SLsT��UJ{��T\�F=�0mt"�
�z}'�=α���Z�!3 A�p�Uv	ݪ+�CBPd� ���PAx��C46�7Q"ڂZ��-׳׷��\io��zLf�7� O1�9���	 ݽ�V�<c�^���͆�oS� ��ci���{�'�D���;v� $1���Ue�GL��@�ͤ΅��ǟ�+KM�l�wۆD����7���`�;��9�z�����E�9�"؈n^ ��e�/cW�R��ҙ�A� ��Ƈ^$y˥l&��י�s�ܕFv��ذ\-��E�����d>�����`D&�vUI�ԧ��j����w(�x<��=�Y��Yٵ[�c� �9b�(�]��ܒ�|�h^p������u�{s��Y��j��D}��{S�@�??5o��ZGܸ�>���(C5�~��-7UBdiݺ"*���y.M�;r��)���AF@� ��J�����{���@��!�!���\"�)��D���a���3��D�����tO���Ŧ���`���K��x�u��snʺ���j&��a�8YU8j����[0���k3���b��F}C�c�^(�/,�ʥ�����m~j�VXxO��x�ƥ�� ��t�(�hd	T����������2�&h�6�E�0֏8��q�� ;Ik���K� �k�r�e]��e!<��z5�"�}���<�r�\Ac���K�f[�f���������k���S�� ����w��w��O�S6Fۚ���i�#�pZ��e�\k�o��O�#�g�dh����UMמV��{�d��5�h.�>�Κ� ��LY��A���v6D3��Ҕ@*"��Ahet�<v��čc0��n]��0�7�8=�܁5Z�l��#+��ӗ�� �#����F���m���i��\̄і0��#�cG�(�Ch;��3�c��}���M>��M��E�֋��4�/jDM�L���׹�=3�e@$>T�>� $0�C(�0
C$0r(�hU������z+��{5C�����8C�;ۂv[{y����?p��g%��viG��;����*]�\9��a�;�O��_>�o{	����w0����H]�"�X��	Wn����M�k2� �^6�7�p7�����8O���+�	 �)�k�۳g��	�YԎ�,>��}��Z*:[���m7+f�sW8��Y�e5P�g��g����:쟮=ϟ!"��zb�E=�{�>�z��X��b��k�H d�	�x� f�.���2k#�o�d��)���a��1pG̝���A��ʕ���dE�5o8$Y�$�ބ1A��|������|s��;OBn5�>}u�E߷3��D��r[��n�C����?���dψp@�1�l�1^݁TI(f��"��u�T-����5�y��G1}L�f+�N��s�w$;p�w8�bN42�<�T��D����t# �.�i[������{�@����4��ќ)n<�晄̛;��=ZY��� 4���! �H� $@�E�)��9
�@�RT���L�+?�������8�<��M��Y�&�������������ߑ���u�\ռᨄe���qE;�ʯ`�����
��F�Y��j\2������ۘ.�;:fɖ렄L¶�F7rУ��r�t����,�σ��CS;�A���"�8|�9Y�"��kxx�z`D�UxB4��0� �x�t��7��&��8�<��7ovx���z�1��9�{:מ��w=��gB�KC j���9+{�b�'�$`i�����\9�$����:����#6z�f����<]��P�E���U;��ɖ�(��.�6O�.�'�+�1{@n�!6��B�z�B�4���q]�Rf��6�^w�t��wny"-��Ǧ�p������P��l�9OLi���;��z� 2�ɻޭ��Z��;����cN��,����(��Dx��O�obT�����6\n;ȤL�+M��<o�N]��g�z5�~�Z�C�B&�X�Ю�g����# ��\ ��~G�o=�LR!L^LB"$Ą�A�a��uy,�������޵�r�4*�ӯ�Hu���a	PN����B�Qy2�	$�A����)�WN���晡�4)br�&�{uɮ�[e[GaMs�V��#D�1&��s��k-��	�S��\�ޖZ��5�b��i�}�����iK[)FhM)��a*�v�^������kebǮ�qB;gI�!c4�-�����l5.����\��!1+���.m+XK����㋂�t�&���9wCQakrT�ѧ�t��q�w�}��N �5N7��T��\�Eg����&����`k!6���+p���h:�X��~bA+�LX�v�p�Ɖ�/��x�0f���);�8w�'�x�:9J�.S'<��$y�����1�s!��q��
��"y�;��ȍ���z�k�teVU�Z���n�o�G�\D|K�{ۧQ�o(w�r!\b�������.Prg�8#
n�`m[Y����\�Eg5j��M���C��x�6�9��Z��C �U,���Û! f��<-
��bvӇ�'޼��[��e�Q��q ��pE��_<y;=|���+�>�(��Z�_Ԓ|~��`$Ǝ�J��sT��;�k��1��П!	~pH�d1�6�7,�X�L�o{�t��;�jl�c�+>R�|�̂L�pcPJ&���XA�A؉�����]7j/n��	��R �m���������*�*J��)���A�^XV�qO>ySc�,\ee-/-�)]��5�� �c�H���e9<� �½H�E:nԡ
0 )$Y$Y	a���I��F��`�Ε]��,��'y݋
 8�zd�K�3��'�:�x5�T��V)`@�(�'X�1l�I�8@���`D�R��#���fTLe���t���Ňv��D�Qd*�sK!wn�_ҺCY��\9n�A�O�}�f8t����t�ez��Eu��R��BR��,�ܐ]��7i�"�8pEq�|%G��?�E��U���#/���;&Zi��qW�qe����V{5�#z�e��nD�T�'��ό>�k ۵�.Zf ���(1�:��A�!:3��xJp�CŪ�L�w��x�У��7�5u�Ԍ\�����YV����q7Ƙ&��A�w�y�k�p�P����1�8B뵛��Qæ�����2v"��96����@S��<D�S�!_�r^�ި�ߨw�ݔ2<@��p  30`Gg~�{��8�n��]���|J'���h���r������6��p�=7��fɏە��9q��>RN��o�Y'e�ќ�;�d���]�^����S�u'$ͻ���<h�sPte��^�G�S��Ρ���*S�Tx\}�7pv?��g:�YZע�o��Si�y?{�9�⢎ws{�����y����!.�5��=���ȱA�b�%�HC�uL�h!�*]c�~��|��A�W�LԳpz�?3�}��Ɏ�g��4^w�u���v���\�dk}��e�/o#G"�#��/�� �N}㳰{��2���`{悜��ѯsZ��ݜ�s{������缇�����79��c��]p�&��D�U$��=�S� &���܊Lwl&�խ]-�~{~�ES�?m>\����y\�=e�cP���+�~5���!��ȿ�I���z�����RT�{5q2��x�H]�2��w����E�uG@��NL�v��t�׺qL\��|1��|�p*f�TJ�5���v�_��z����J��P"� ��k�4/R�m�gAy!+Ȉ��_�2r(�P	��]�՞�h*�ᳮm��g�gE@�����{'����q���!� F�"K RF�(N�G����r������u�޺3��E����6hӧi�ʬ\Ou�э�un�6���3�D��I;|���9���H�3��36%�h�� qE1�ԙ��83�����ٷi�A�wI^&���^{�f�4��®L���y�q�y凩�o�ʧR.��4¸���ܦ<EFK:0؈"qB �2H�rX�`�C$��ى�z��S�|��}�Gk]���13��q����1�E�*72b�h,�*�*���TX��O�����3��������|~��Y��?�}9-��S��H[b�X"E#l+Z2,D��R�FY�������������^3�L�������L�H#K`[B�TQW�Q*��8�V�2d�rnnx�8�?Y��?�oy�9���|�b(/��fݡF.١F���(��T�4�23&MM��8㏣���^3�Ob#�yyʱI`������"��!I���r)J))*�������_�8㏣��>�g�?����Z��k`�;h咤< 2Q�1
��ԕ8r(
�{{}q�����?��}�3��||�݁P���k�3)�V� ��UW�IZ"1jQR��PE2i�D"�J3O���|�d�<�b,�
%b��.RUb�	Z�U�Q5KF�Xi�=@�R,PuJ'P�,I�˿8�AUT�R_8<Q�Lf�fس-��������§�2� �
�,2� R$�+�Y���o�k����<�~��o��l~�&y揦�{�3#�h�H%n�P���|��k�pZHFu8,	�)[�9^�[��7G�x!L��A؏g���2b����BN�`[|�������/ܘ>Jm��칼��I{ϭ���g/E7�d��B�ٷ�]J8t����M�1��<�"�1���I�}*�_B�}�~z�*�ռ6+�.p�a�e�npT��54�.�*gaЖ~Q�@6����}*�]���~�"�όcw��` Ϲ�&����y�6��k�k1�O;`����Lm�f�GΜ�uC=�m=�o��o6��\�AQ���V���<��ϹNTZ}��KO<�"<�A�_U֞-�l���M?q�}�f���u����zִ�	Z�p9�[�.;e3t��o8aj��3/i_���2�N�榆�0��9o����O�}��ߵ��h��������iI��3���Ǻ+�4�sͰ�d��zT��r/LV�,�!P(��0
�����$�C"� ��0� @�u*�H'Ƿ�?O�}�a�k�rP�<��/A��\�ͳ��bXcjp��j{��GK�����'9U�
��h�z�>���&���1<V��M�_�}?g��~%��,hFm���Z�e�Mm!�K��)��{?��m���#R	��+BȲ����%]�i�:��g����<| y6�.!��L�8k��ڲ��y<���"���ǽ��`_�1����p�n��]WӼ�� ��i"�O��z^�J��.����C9�����P�^s���<=[0�7�Q����*u���V��2��B��w. [ m�=޼ٽ��`��c�s�Ju݉����{�=��>�^.>�ANo�<)���!��1��jH'؜�j�A��0r(�߯bX�Y��BF��m^�*~���i�n��NE��L��^�ջ�ꢑ��JU
�[ꩲl�ŝ^������|;���=GW�Q�,�s���^��*��8��S$ヨ)#p\ù�'�V�*��B.Ȅ�Lg<]���tc�!f"V&m���q#��>@ݿ�8���d�BR$"H		��a�9)����
�y�����tl[#g�`9�����T`Y�*�.���9u���BRh�u�6�qW�ר��5y�bL����s˦&�A�.���:)3�=a��93RWl��ڴ�ۜ�M�p��
�Z&ŷj,���k��ٹ���F`q)��G&�L��c]�ٞ
�"dl�$����xQW��������n�9M1����ہ���
6�XO<�����År�A>#Y����N*��^/:{������d��xֽ8�[0jt$r���& �;"��>kP��+֮�����t��g�bb�Y�{�=k�>�1p5��������V�#ѵ�5�K�Wv'NJy��R`�f&� ES��^��Nü<s:׳�N��m�lP2B^k!�s�3=��g:4o�W)c���ݹ����xBsW�,*��.>|���'[�=9��A��ᅸݠ�̇g@�]\�?}u|�ϵ�����:jZ�z�X���9T;LDk �
v��V��=y�^g�Aږx �M����ؠn�?���ڨ\9�	�� �|m�m�e��m��h�-��bb�n�F������/�1����,ʩ��=*�=��^[�X�\5��w_����ffDC:c��F����}�Ϊs���e< .�����������i���)>�bB�w��`��yb6����r�H񽴉�a� 
@���	�U�C'�R�@	��+�}�~�"C
ș���	� t�V�
B0]J���p~�|�}���뭯�LTg�*��I�p��qs�I�\H�il��a�l���9N�Rj��@�_m��s9����{x�A7� s[@X�U��N,�!  |��Š���Ad������$�v!�6��ֲ�x��t�Z3��E�>[�(h�#���8�I�|9)�n�� j�Aб�Y��)|΅�6��׷��q�3�����Y{�ʻ�V���\��z����A��Űc+A�3ԯ�>wU7���X<?�'VG�g���B}�3q)�G]�Խ��=L�kl�vߑ�-Cz{/�+k�&.3�"Y[�h9�ሲ$���Ls{u�:��~O��>�F{��i��N�ǉ�3?��������[�n]F�M�a&�i�Ǝ��M0�4	�� ��Am�ER�.��{ܥ��������8�u@��66J�"�Rd��b4���Ă��w$����d�ä���33G�� Q�U���R���J���w����Ec�"�s�v�F�x?0��і����K�S��yo��5<'r�*;�7��ڧ��0�ӷ:��<�����^�R=Hj��K���7ޡ/���=f���ǚEJ�#S��f>G�eX`eHeaH` !�A���t����]\b� A�A�"��1�(�2
��o��S�����r=m�f���f�
�I�En�ܥ�������@� �r+�9W-�g-���]���xY��a�a�Ǔ~x|�ۜ�yÍ��o��*���W���C�:�!٪^�ĺ�o�w���Xkn�����?~��>З�s�����dcg��j榪E��4d�:�h�����&��w�@���P/���ʝ�JWň�!����"�����ra�<J��p�ǽњ���1?f�/a���0�zA��\W&�ZK!�w��R��r�:�qLE�������Ϊ�Q�0of�6��,손6В&�v"� ���sz�:�ng�H﷒UӋ�;���;:�7�C�P��+A��E�n�\e�[�LYt��� Evvy����+���1��B�z���|��v��f���7��s74-�	ؑ�p繛e��$L�C��v���mj�}���Y���1OI�x�T\���b��2�a�!�@�������[Gl��O=�G2�A���"w�`��߯3�����gd�BmL��}��S��r�:�qy�x#ő�NAcv�<Q�/���@���HN�@�{����>���[���sE�e��H�����*:����G���>���i��J{�g�����<� ��)WN/4�;���cF�`6�g����gh��� ��18#���������%�����N#soѕ=�%\g<Z���p戡��TFM�N<�]��,h9N�B����˽�z��ϳ���#���ש��bg� j�LH`j�5[=1Dsf�F�3cHx; �� �H@��>��t���v�y��K".`�kLk"��Sbq[A�L�h�F�D?)�9/l���UWӓ��3�8&�A�g�� �P ��úƋ;�
b!��ݛ/h��,]�7����T˞��<�X����}�orv�zxią�ص�khP$�����$���͗�{��%��Ɨ�j[hya+2�'dl"ac5�G�ʼ 	�N <��#|ԥ}��{m�����G�ea!��d��</��p���I�3�ЉJew0s,c�N�n�j�ivlqc��\Q���)P�":���Ka�\��Z��E�T��:�K�G3@P���u���и���f���q�i��VˢKV�!�`��j�Z�G���
u�lj6���V��4&���B�V+����|���?Y���!n�]M4�[�����f&UQ	�m��ݟz���G�X>A9����nቲ�����DGa���\{�<����}H=R -�r��:� ��dA�Aᐋ�~�Ctkm(
0#<��tt_��UӋ�w�%��{c �w����p~��;%��ec �'!2VD��lǆ ����V��.m
��g�f23xE�g�9�r�v�B�,\�(7s��q��<H2c��Z����n��	!��>@Q.o����c��gn&㘜��Zw!5������~�&�9,��G��߿�!E�&�,4��:�"b���K�ʪ</{�UӋ�w���ЀES�bh�S��^Eu՟)(���ѡsu���ɉV��V�[t�8���2�OP��j���y9l!��0M��_7k�1���.#<��~����=�9�!���86?��c��{����<����<�]��N �@�;�����ط53�C�`a�z��l���K�Ar�;�up*�&zK�WQ޷4wy�A�^�3*?����$H��#8��d2�K�)�'���n�ݟOA��Y����e�ݯ��Ú�^z�x=�?�嵩���5Eǹ:r]�3����A�E��ݛ#("{h�03?��ý��WN/��
"�T�1�d=j(�	��������($SZ��kٳ��q���l#�v�t�4D�-磉�~�㷑�|����/9������z��4oe��"<�*�/:x<Wa����q �����n��� ��c�)\��J5�t����>������[0Y]��R�+��ā��lM�v���#;�_aϸ���9aE ����>��*�NsV�8����x��c���L�B� ��@U&��s��
P� ,�s�0
�[ޯ<���C�g�,	�B���G^d���������a��]�R�i7k��~~�q��ޟڤ�$Vt�-�<��6*{|jn`*�������G-��e�9��g�02Ү�#1�F����c!��2��ZD,�"V,�dH�W���[����O��v�n�X��r�L��9�"�q,��o�+�W���-��X�q��Q�A���J�NsV�c��@�7�}s~�}��������e�/��"Nc��&I��HNͪ��� Kc-���V\��O���p��#3���D�Ӱx4�3޾�˨��C���a��>�xNB��E���SMd��4#��inԂ?#��.[A��b�eÑx���e^������f:��q{u�-둹�؍,����	��k[=1$ �{A�h{�z ��i���z�����*��j��E����Ȼ�y�_��x�����M`a$�r�H,o�nBF�G18:����s�ƫ��e���ޣ���<A9(9a6��!S��\ANM�^����H�i��a�K�:b�<Ԡu�߻���gn�v����vW�c�^��@=����wx"�����"	w�D>�T���.zլ9�yOݰg���<��B���y��u������#�%��C!,�����T*@��O�N�B1����S���D�y��?��}��P��6t��UQ���.���xc���ˬ,�߶<��>�����.�.�_߭���@�E�
��Y�Л\ɂƕ��\�4%������72X�ai7h]��/;��w�w��y��6	�n�d��dk�s�0�]�q60�*��D�DL�qa��ݦ�ű2�]{��ªxfd�{��jn U-�Z`0�O�i$��-:��r�8ph�!��c�z>�|�I�f��NbN^���潆vh�M�9n��-��)8)�!X#j�c�.��z�I���H-w������^���Ci-lG�f�^�o��[�ik{`E� �6�"��S�UO���v��\�v�"�36n�gª:�gn��T��<��@@-T�3�0`<�*��jL�Y�z;���ٺ���]������Y��xs�/K���[��590��#'��F�j�C=�����Kd�4��-Jt�S�`�0\�	���)��B
�v/v������z�ã.nq�Y��y&9�9%ǽ��J�:�i����݆e�����p�6������F��/y籖0{*ŝ�_D��GE��j*o1q2��8b�(�x��佻)7�ڊ-7����1����Ü�C ���&-�݃Q~��<�d�k�^+p�/���#�z����w��1)��x�[N��(��v�]L�\�I�p�ϽI��AG��xf�w] �ٺ�2��W�]��0���u���9`^��2��kU��*�Bخ�򤯔�k�;5��;�&M66-�;��'NK��(�se̪�����wg�{x�Y�)����� 6\�^��n���W���aЎs�v���b�}�/�oΎ����u������	Y�ѝ�G�-Wۗ&R�p��ߧT=}����f�?#�3z_{�������7���1iZ����:}3�j���HKt{���w;|ȸ)ь�ŪT=����iZ�0��xjT�zDFyn��{)5�v+��ݼ��u�����Ҥ�Ʊ�Oߗ,ʺ��S��jV�߷wu��C^�� i�	��^�sc�4u)��a?^Y-�D�C' �Iո�������m���vS���[\�T�|dL ۨ����lD�v��ۣ��d�_$2�13eudg5(M�k��8�=�s�9�B�o�߆<4�I��c��J��I��L���{�D e�p��G���6��w9���q�U\a�e>3Me��%�G�g|<�k.
|6ljw˽��o�},�&ٶB�B�W����g<4�ǉ�w��Ő �"��K$ �g���g_����&�
|y$�6��o�Bk��gm"��E��T�!���#W�i�
�ڞ�_mt�1`+?ON������q���Y��?L�>�%`�
��D_�!��H�)��A�Ԙ�$}�d����n<|}q�����>���>��>�3>H��(i�@�]Z*�,��ĕ�t����&��鹹���t~>�>��>�AD\�Q�	�,��d��&!X"E�_�*
t��P4��ۏ�����������~��}��d:���rB��N�2����ņ�f;h�����n>>�>>:�::���?L�o�VVcU��r�E~�����Q,S�j���k���%����������q������q��9?Q�;riՕ�
��J�"VJ����@W-O��VbWH[eeM$�B��&!�
",�E!R[b�LCƳ�DPwJ�ʕXJ�i�*
��VH��T̠��y�
bVno0X�U@�-aPDb4o�bbG<���y�	pbcT�iY릍.�y�i��P�qmuV�w��Q��Ը 2�n4T�UvWFiIaL�.&��5�Q \v,-lpK�cA�mw��%�S4 ���!� ͚��כ0X�F�3��4�H36��l�jiV�A	,9�f8a� T�m+m�[�e�(�Uo���#��u�-f���4�H�ͳ��b�к�V�=�.���V��6���\0�1q4k�bJ�m���-��n��.r��1����g�nL,r�+SRcb�+���m��+L�2����+DQ�����&�Q���Ʒ	����f�n��2�jQ��ڴ#*�c�fnnq��b[oa��^Bz���ZL%�ZX�i�bf�ۦXh�2��dɬ l�4�t*�WY�j1����X�Ů�+����3X���[�쮘#�.B��ҪX5�1-��@X��)s�&GVsi-��LD&y[i�,,B�Bm�Z4�fs��R��j2ذ��ֺŵ��R�Ţ�G�B2�fe�����m�1)�R�,���cV�M�[Iu�QEk6����X���汆"�,�#02��vS)%jV��[��e�M���q��]Lqi�-���3ID�4"����8��4�nP��g6gF+6A��Aΰq�6"��k0e��ɡ�)�ر�1���(.HCv3ūe0�ۭ���Ғ̗
��P���Za��8%��r1�I\7as�B�S�M�KQir��S8Z�*[�@��\c'bi`��]	���6�w:��h�u����V�V�3��-��-'��w̺�ezd7V�E�Z���7�4����"T��1&(R3	�u���x'tǾR|v?V��r6"Tk,llx�֭*[.f�������C�Y�x�$�Yq�m����<.��B��԰Xj�kLӗ6�Ѥ2��PLMKv Q�a׮"�[�R�h�l��yT����h��f�F8�gK3�f(����2�)��.��ڣF�%�q�F*69�g�?}?��p�5tnj���h�[�6x"�S-���ʏ��.{w'}�8=J���r	nܣ��=/o9�{�G��'8^��x���b�x�3��Lܡ��"�w9)���Jǜ걍BW�ALu�%~������"�8am$�l���"�Ãd{�>z�w^��T����P��R��$���܌�詫�Q=�=������y��v<[a�v����هпh$�1�!@�.���޺;��=֕N�ns��N��Qi|F{C�,,�~���(=>�H�v���=�p;&^��՗]�U�^��C�g	y@][8m�"���ZY�+���$�xY!���)B�V�d���Ͽk|�����-ƛ� %e4�U\�)��aKt��K���:	�&�ծ5�!���ZdNN�t��8��"j|{�5Kc�#� o��U'}��:b�F�i�,���y�*UTw`wVM���G�7���*��4n�Hp��wtk�e�����z"�}�	����j�q��o��^�k����R $d�JD�$I�}�&���ه߽���a������9�HD��U:���1���k��N���#��c>��l��\�ILUl{��Q���[�o�8afP��2	��!s8�$h�8�������K�7ť���J�E����t𪊾۫�el\��� sM{=����������Z��P)ƛ:���! �����'Տ?SϷ�H>�02݅�ɱ���ڙ�6�̼C�b���،�v&��5�i���<q@�N���#�v�0X��37Uu,*U��iaq���3�]���O���r	��N]�3�g�S����}���o��A�]�d���sQ�? 2����Ʃb*�8�HIDl����j�4|�g �����}�1w�;us�NX���V�U�4����Gu�!c���v�p,���x̺�j%�����:yٱ�Ws
���=������{twg�{��,�Q�蝾Yh�����Fl���L��Yeg�Q���"O��e�fҌX@`�&a-�;Oxןxڙ���F��_����s"��g{lL3~?����ܜ@<B=��e�Fb�3zw6����[�6�{C�λ�;������LO���e��g&�0�R�B�|�'{�Kh��x1]�<*b��=����!8 ��5I�i]Nl-�I���ww��>��l���,Ĵ�nօrщ��llcٹ(륟�Dp9 ߜ
-N��wOk�u����>�qU겫�O>��a���A��h�ނH�ԃ�Q�N/*��!,���N=���M-�^�K����i�fb�����}�V��b�t8�z��f2�Z�46�O��Y9�gc���R�������X�ܬټ�1w�;5p ���U* ����K;Y��U��Sfja��id�1 �w$��o�������d��(c挭�39����w��B��v����^��m��}�j��+��)���}J��~Vw��M�L�F��Ğ J���Ŀ�~##<i-43�������4����4�c�?2
�j��z������oZ����}\g,��!���gh�zA�g�A�\'�r!��N�՗�ޥ
~�5,��@l6�nM
�ڡq��@6s,���!(��g�HqÀERg�{��z�xTE��٫����8{��������x0x��]�w��}�ᾨ�={7,�vy�����9E�p��D^A�~��9ރ�fw�q6����Ȫy��s���W��F5&���}�lA>��A��P�R��޴�O��9�j�/%mhS�x�gg�Ec���4�O�Q<0�5�Ѻ;�yb�Z��o���#�1n����1�����w
���ۨ�Ǐ�~�UX��<��N �'QE��HH KR�i>^�l4<�z�3��zQ��m�g�ҋ�S{�ֈ�h�i��=Ў�ն�U��yEz�T<�Ͻ>�w>��K�{|ߓȵ��?]������=QM?>�^x��`I<��X�*A��/���}/d����Ƒ��3eo��{K3edb�&e��a�w��Y��bf�b~'�$C�J��FD�12H���vS+n:0���D�%c��swM�.&���o\#a
ʱ����M78�,k)nqcVl�Ɋ�A��8S7R�يǬ�[GM���z�R.�ڣ����Ѐ:	e0Fd-�����4�	64'%ц�
Q���,��3gc��g	����`զu�֌Ұ���b�c2@���ϲ��v����j��í�
�[i��˞ڵ)��b�П����#P�ڙ�,���L����z7f���Fͼ��N��<L�����K����D�0�ҝ�:�2�|7�|�c��>v'KqY]��R�}�;usA�N�x�5KZ/����!Q �z�����\����gs��7n-�V�����=]ܳ ���2��;V;4@V�*L�R��&�Ѽ��(bd��b�8z��zc}~
1�a�XT�pC����w�L�cI��m�4��a	؁v����6��m,�u��	���Y#ۨ��	b��qD( �O}ק����qkDG߷�n=�\җ55�#f��^���ٜ0�s5���m���3���`�~�#�q�A�p�+�z�{��UN�V���{nn��y���0O|ɑ9c��t�yˌAؿ�|8?�q2��r�����{�8���<�<|���m���/�t�mS6�x�y]/Z� t�??�Č���)�4�'ι�SW��說��������B<�N���&�Ch�v<�W�i��K�L?1���E��iXo<���{�|&_g1�۫�Y15�xY鑨N1@�MF���ȑ�㝍�8��ccd"�ۍ�1����U;���k��5� bp[S+]; [&�X�h�TŲ�> *�z$W���GsZ�gL��ވ��>x�1�; ߟ��̆c�׎�������9H��%R���_�����ݴU���B��]��.i�l5�b̩�����lG�pʙÅ���X�E���gp�~���n�#j��N��y�Av*�C8KJDԂ�I�9�� �m����l�ڽxݟ /_�@Xf����T�5o3�t�)�B�Ñv��>�e�)e���N6��	*�1�[/1��c� \:vn%P�>Q�M�M��F�yb��]��<2���L
�5���������b��9��/�a��k�h�`#�6��6�����K<j.]q�GMJ#���"�HĈ��br{|��y�\��Y�0��S+���!�Y���p�NĂ\[�ցW��<}�	#e0pGjg��cެ��<�9�����&lk>4�����UBm������
����_X�DI�A�5���G���<�1�"�^��UYͷ�耎���)�k�b.�8�13�D��ܪ��Ƞ�$#%(w���_���m��;gb�ԚF�M���X�0gEȘz�x�Jr&@*���J��_k'ޘ\*|0������z�51�s�H@�n���
�H4LG�ǝ9	����#v�;ie��W����g2�jn	��\�@�dڛ����v��y&���G���ה�O<��d�G�������>Uؽs9^��>U�ۜ���3svc�vv�Y�x;�$�JmkL��M��Ӂs�_o'ޘ\*xa�	�A鐺3����_����	��Y<��M��pm�]��w�+�{���BoF��F�1���Wc�+�N�x�=B�n��f���ғ����$fI
K*�%�7��ҰNy��s�	�H�(b�.!���~8[,L�g�W���r�8�ǘ�o�"��j�(ݣ��HѤ�W��/]�I�]����Z2�}�1�鈡]B�ha�uɌ��R�8�Yr�0Fg��`��2<J�Nf{��k���xMVsns�Z0�ﳋy�Ƹp\0=0�&�M��1�N��H,F�jޒ�Y>���Sᇘ�Z��&�"�d�;}9A�5�ިL�d�#Hs,P�q��lDZk}�������u]�����gf�b��g�dn��/
�?�q�������B��n�8ƅ2��ý�/��>s�5Y�6Jps�1FD{���|-��H�v�dj��MRslP�Ȧ�yq����:�;2��#��~Z�)b�/��	�<0�c�C 2ЂӇ6[ �n3/�b<�ͳ����g:y�1NeG��L���>�pO�St%ƾ��&[�� �B\�{� +[)5�0�F!�ӪU`�[Ա
0�3�u�[�%��#s�G���W�7E�?��R1"$D���Bf)�Z�������Q��&�k+D�eȃ��	�悊hK��66JJ�,�ֱ��e%�q\c�u�0��i���
3;&N�jX��\Fkj�Ex�gqKv�bՑ����M��+E�J�
��)imm�v�1�k45�{Q�΁v2��oW�3#kt��M���C�R�_�����߉H�ڥ���IMfv��Ci��U��жd��a� ��D���
�gj,�7ۻ��*2k3�W3N�pmf�U��g��k1�6F$�]���s15��b�D���5��?l%Y��C��d뀘�@B���z'��tp�LU&�	+�I�{C����b�7jh�o��/=sx6�T���srۇ4B"�0t��'���-�J�KyE�jn$&�B�W!��lgnnw<�ʬ�f�6����'	�����������|��I�9h9�9����5�C��~��ƷL��?����m�8!w�p�qLFe;��;&�RǻH����ޥ��>���t�3M����&ۚB �3�mLjѠ���\Zy9`y23E8 �j�����W�
��8agm�?En���tX�Awl��c����A��̨�4���b&�j����v��[�ay�O~zY���.�,��C���n��y���ʣ/���c�"��2"h,-��qo���*E%����}�R�%'(�upv-	��;�7{臉���m+�s8���/t߮0ئ;k�QE��;n݃�+!ȦV�d��z��Tz�6a<Mg��6�x��"�3�dj��T��Kn+�B�ɂ���'T��X�s�ÆUW<:_L1�AŲ�&�q�q����9n�Cxt� )����tu�Ҝ���W��t��e^{57���-L�2v�y��\�۔7c������{��u-�������7s�����&Z��v�0�iqe��x�Xi�u�6%��Y�_V�G[�ce� ]S�v���ouBx��m�q���{L�y2Ц��복Zg�P��:pX8V-��������V"ı�MW�j;�]��Mp�t�c��db�46���A1asa�vZL�07͙�nL�!�7�߱M�G	�ʻV)�t��t�U>��r�J1$O^����Ӓ4�
���/�һ�����-߬QV����!��	��$��f�crg%^�"\`�ëld!�{��q�
������:����;�hs���yy��:�&z�8�(e�6�m=��!�P�)3ݽ��5�L��2���=���;�78.5��]t'�)��{�����N�C=���{��d�xtr�5����Ӄ�gz:'��G\�تg�o��+�������BwMi��0������1���빴�{:zJ�we�8�	�;z	��������8gvv�h�E��{�G����/w/A�ujl���9�~�U�x5����{i~�Z��i�*	�>7���yv�q ��ڶwOk��LM��ފ��8G���ro���d��=� ӥ���Ş}�T�/���VHd�o��=X�����mXA��_U�B_��N��_�}��ۇ�fd�~-��e>�ߟo)�v�����1>��C�A�3hN�+/�|�{7f��tW{�얜��6�������Ǝ;�(.�o�`�g�h��63鴝kz5��.-9�|A9z)�{A֢ܓ1��c؏���0E}H����'��G
�;�󯗵(�զ/����pp�?a�4��E�X�1�F)f%қj�q3+�PU}��vՇ�G���!��$����z9f"���IBFd�,c$$<%c˦�N97Y���я.��7ޯK1� �d���Dm��W���]���z/KǷ^ߏ�����㎏��ϣ�>��E<HV*�C���TU�M�&��
��&�E�U��,�������\q�u�g��}����Y~��Z�6����,PEI�+PYV1@��,�}>�>>>?q�}u��q�}8Gەl*}��i� �(���U�qz��Y����������G��3��ϡ��YU*�,DY(ʊ
�J�\b���r�X/O�__�}_Y�\g�6>C-&$-��&��J��cPP�!rx��
�[E��99>�>>>>>:��u����Sۜ�.���!�Ř�,X*"��Xb�Lf{aL�`�+ <o]"�MZ��Ib��n2��ŏ־4a4Z�QdQb�QE&�I<�����#lU��(
�	YR�FZ�Uf���v�=-,�����33����C��sU^��oLEN]�n�� ���5��6�YCVY^�3�8Bl���VEV�׫�v��A��;N���T��U���8 �Du�ߋ��ʕ�<��[�h��oQ�yr'P�/����nT
�,i���z�Tn�w�4G<p�d���Z����H�wN��Y�ңc�5�k�z�����j���1e�fz����٬������;�|��F^w�Ov}�{�!����w�!L�OV{{��)�/4t7���~�<��%��%W������C-�+1hd|��C��ϻa�B�����eotӽM_ Fo�(��l�ņg�q�xxUHs��yL��yCA��8��Ε&pj�*B�nfd�yx�ev��5C�ۈ�p� &�p�Y
J��=z���B#҃��<���!��o�9�2�Wթ�����=�K����>?�<���=٧�|���l����;�o�6w*�������w�о�y��X&��_�~&��r��RZ)��\�������=��p����`��d�>;w�����}��:�[�鷩��9���j�a$T����4�}�{�R�(�(��Ď��-ثh�.���b��̉��,k�jmj�M>�O�[���rd4��k�7h�gm��WW�>TW<FQ�����C[�2#��Z�"Z ��c3μc%ϻ�^e޸ͻ�G�&.<���-��W�s�Y�5f ��+._<��V��h,wS�o3�_v����p�,���=@���ޫ{�����al���|A؊��C@eT��Y�����R�CHige��&);Wu[�{��*+�.��6ǷS��Tz��oQlb�����8 ��EU*S��S��f�=�����n�-������"�u�q�rC�v����ݥn���'?6n�૽�'&r'ϧۣsKؓG͞}���Eb�B�԰�� ���>�������'c��'�XM��D�����oV��c.�c��������7��Z&��Z���N��P��!
K������@����Y��K�Lq�QGms��\����v\��h�Lj]v��m���.f�EJ�\��fy��jE��
M-�V�6�VP��:�̱��-q]�$f�r����ڠJ�eвV�%�tJٲ��M�{7f�4Y�R`�fY4��l�V�Q5k5��tf��nw\����#V[��0�Z�I08�`٦֌n�cj�ca".�eǜ���3g�L�}�z���}��W���Ǻ��m�x��z���q<��3�Ӊ<��&�g��9��/�)$
�� M�pi���P����� �
���=�[��Q^xX�b@wl��#�]���D�����T�
�+n�m�1��AL�9��m0�s��b67�k��w^�[yۋ� 妜M �'T�
.
��w]]��nbA�>��T� [86��g��gwV=���n��l�Xu�S�'�w����Zm-�A|���g��� )\iQ�v)a��M��������TW-�- �n�DES��y������JYO7��(Ԗ,ӳ���5��iur8+ZJճv��Tt,6��hGY�g�����H�!�8"����2���}�]tb���\F8�ײ��-kT��I1j�4�ːA�A����s.P�p�ޜ�=��n�
_/M��O/)�����'�&G��ND�� ��3|��(�?^�?w�ܽ׏�;۟h��z�Tv�G7�F{h��M�������).RX�H��!�h|�eZ�ǯ�Y����̩���M$�p��������X���E��( �#��d� �R���ko�3�Z<�O]�:x�2ڃ�2N�	��+!Ĳv."�>w$�P7i�ϲJ����nr4�������Mv� .�}Ü�b���M�-cS,b�q�I.�c��NZ-$,��v��d�p�i�:���/�ۢ_�nls�����ۈp2B���������������m�K�0�%��z�vٺ{�-����	�v%�����ٰ%t���u�&�Qr�����o���'),y����:�#��ò)�H��l.��3)y�+CC���̅�E�FL��.��#w���`�;{{�9�ŷ��CX��� N���P�c��������@�BX�m�"N���[�&}���M�{]�?�6�E��;}����{),�+C*+Emd�Ux�':��'��z�A:�t�w}
��Y�9�`����A#-#JE#���2Y�ܿ�g����S���;Q��S�e�v�$h�Rq�K��LB)�>��.C�C�'�nS�e\F���dS�0��PG1b0c�u�Ţz^�F�#X�w�U;�h�Fث��]�Vu�_oJ�pv<�n�=y��^�[y����X�� �ڝ��-m׈�t��]��R��⼅�F	��kx"5)�a :�{��}�o��g9�MY�iv���Z5�63-څg��'���f �;QF�T���m��>�����Ϭb��{=NF�.�vv4�]ۨY�4qsN1;ΖD�/�L��}W�uw��ᧁ�2��> ���"�I~�`G����ypA�]���gLsH��UU�#U�OD�G;��m�f.�ӖKc�gJ��X�'Z�t�����]SH��0�}�{H���̎�vE<�m��Ԁ�k���Ub>�M�����wr����|E�C钋������<�~�m��G�����U�ڭqH�����ȆD6�|�m���Kc+t��ݦ{L�R������ױ� :j��3_��Q\��v嘃�Fۇ6B�B�
h��ē�2������k�����Y�Wm�XgdL<c�Qh�vh�6���v�)���P�όF����hf ��&A������ng^�̄Ͻ�b)�5�19ɑ�&j�-��"T2'1p��P�V1�j�̂�|c
�:=�u�O6�3��x!��&��u�Ց���'�eܺq'����~��9�4�+�U!���`:qf��#��k��[�G2���!�����=��G����ݣ`���y��v6���t{�9�nY�{[
hc����[kR�8��K�v"2�7VvB�����8yd(���>����8�z�Lww�&"|�|�"
"u"��X��\pME �m��=��B��ӡ*޶�<m��PQ�^�y?a�����}����w �)�� ��0���~[����Xp@�_�DPJ�B;m\`���
�K@0���ep�[nt�1�"5B+��alWA�-����u$�D'8��{�զ��\i���1fs�t�F�f`ZRQ��\�
^9�l6��[S��3�a�k�Q�.�Jݣu�KRV��Ͳ���Y�&]*Vk���׽�X�M�[��10�q6+��6&[sC%��5t�����
p��Y����V#�a����V)�E7J�a��#��z��%��*j3[�k*Q��ٕ#��6�Sb���Q>п �el�
{M]��0��\⺊ގ�jj�4���Ȁ�]���چ���CS��߿�r����/����P�kc�C��<^�oOD�����\8 ��M��ݪ~��.hQD ]�5K�w�f��z���f����GC�P��30���T�h��\�nu���6_;I��N�5L�Qd'���1{O��4�&@�X�T�����������a��� ��.<v5�ᙄ���b<E7)��Wɣ.�I��c~�5��#0��G�[ikʭΎ�O��� ��[i3�LY�R� �K�8��<�.[)A�����~#W���;@���̤f��T�3�v�T�qQF�~��_�8B��兕��6f��LW��f9�x� MgPH��MzC���C;A��)L�|JF��� �W��Auz����&��z�����gp^�<���=���~��;Ԃ���{����qdWG4���w3G�o ,�ٶS�?����T�Ċ2!�� ;i�N�&>�Wl;�}�|L�xiln@f����gcI������[!�흐�9�S�F �bi}ܷ�>*#r�=���3{}��N�pu�H
� �Rx�ҝ�O�@��<h�-�Їx�m_ ��"S�v���L{�}o�|��D"�l6�f�C��&C̳Nbr�@�.�в.�:��a��t���~��^�gk��%�Pۖ�TZZ�.<�}�yP`��r�����A�&7K�Y���Qt�1 ݅(h�%Ֆ���qv4SX� �� �e>�BiUsCE�U^�G�����]�>C�"��@�q�d5��o&�V�n�i���"���A�j�GtǷ�n"c�������]�D�X���Uk�FA���&��MT�X��%��+ֻ�v�r��]�w����X�d=�[ĳg��vm�`��s�������)d�,�0�\��^�j��N�����O�"��v;�{�߉����՟�w���'ek2Z�b�U ����]��1{W~l�1��'#�]C>6[�N8��p3ݎ�w��r/X����
����Ŀe;�3�j�-F��yϜt� �cTB@��GiC�߹o�~p9�v�M6h���醚<:����t]҄I�}	��S��L.�W��cx������h���ܾ�MC8��
Z��z�2Fb���ɽI�ksaz{�b�n���+��1�̕W�~�BhlV�����J��Uk��t����K�GN��JɎ��c��v����A��T\c�M��mm�5��Cl��v�������n7�[��VE���r���m�{;Ǝ����T���n����_�^�;p`]W��P3�xK�z�����ג��r�97�*$��XQ��`I����H!���s��(�����;Z�D|�_NNSs�������˗٫��Lyg�&�v,s8�:�|��YD�������0�BlQl�1�#f�cA���Z�6�-�'~���g
���{&:s�l����c����n����sHKQ���<��D�/L#N��h�oB�i}��7���;x
ge��o���P@��uD���tX�l0�h�̇��y��6�0*<���s�9/��3�e&�v�B�����%�&Cg'}}]��,0�L=�L�j�=���l���d��p1\�N�����ۗ�$B+r6�ePJ��,[d8��=�����
շ�H3ךa�� ���e�wE�f��ٌÂa�#�uA�}�f��=�=-�Tk;=������k���s�dc}�1�C\���w��Iپ��ٛ��yL�0����w���O��c��kpN��.����g��{ ��'n+ر��vT�^��yz���'������(�:��+���U���P�3�ս��]�2|��ټ�Z��s��G�����0M���.��uzL�ӉS��¬��>#�h�斞Ǿ�s3���C���ܩzaQ���Ľ�w7#����S(�}�c��J���T��<A�U�_c���uƯ���M��zm]Ͻ�ݗN+5��!�v}+d1��ˋF�<�t�V[>cX�6��t�DQξC�jr^�{w���r��z���r�,����5tҘ��s�oyz{���s#/��*���'zI4���>�w��s�ߦ�e{�vMŏ;��wٻy5���K�z=���o�V�&BY�%�pnn8u�^P�ԭA\ɯ��p�|��HȽ;����ѝ�x�':+��ݓw���w�oq!�C�P�����C��o��@q����͋����顫{s���� %��{<s���lb2r�j'�~xk��T0p���r��{X�p�u�f.H?�r�6�IYB��'���i�`y�|vK�r�$i� ���ᢱ�W�G�Ÿ(��ۛ��j�"�yv��f=�8Wp���<)m7��B��Y��9qB0Bl��i<�gv�DaG���;N\6b�7<�ܐ��}.~� <
=�Q���p�AC�rnecfV2^/�I˸vB+&���&�Q�B0�+��r\�FK���"̴Ɉ:�f���N�?�
��0,8�.@��`��?���йDg�z�m��|4�O�Ǭ}})��{�c�K����BY�c�Xͫn��u�����gח�����ǽ�`�g�N���uè&,�]�C�'�6��N�}�t[,|���&�{ct�ٯ��>$��M�f{g��Ү�3(��8�i��m}>gx� S��Б1|��J$�۴��K<{~?\~��>�3�?$P�R�&��g�ִ�
�יESiX�+�S��������_Y�_�=�)�4��B����(5�XV3&篯�������?Y��G����L��AH()Y�LeTd��������}~���o����}���D4�*
��-DIY�:�u���I����������������g���7�����~�>�^M*��t	Գǧ׷����__G_c��>�Y'�>J²���q���mE�b֤Ir�S2m�N0/����c��)a}�I�U4��8�ɗ2H�����(�PF��5���`V�4\��Hz��`��{�c��h�Z԰�|����w�h����U�\@]��,��V�ֺ�v���pMfKX��	�1lλ��U!Q�؉p䙅�	��GY�&o�+�q��k�BR��8�0�둚�n���6��n֡E����m�\]��#)-���]!�X��j3&�RV��6��3�fT�k[��K���m��Sa&l%�#���B�̛�8��!-���.nt�\	�WD7KqGT��A���a(�,`�݊�%h6%iQ4�@�Iqdoj�-QB��4&��bXcK� ʶ٬�۴L�<f�3s���)pMThhĚe�26jCk��њ�B	GJ�2�6����k����͎m��ؐ�к�hB��\b��PVTeM	��a(��ʛWsVM+^Yf�0����ef�K^��XB]��bh�l+�a��lj.7li��k��I�V�l��l�He�+6���M�L�8��b#i�����y���+�L�vX7b눶��؀i]Fk�j�+����gi��q��E��1�i�	N[�l.�:�h�\d%���	��\f��cCM`�e��.v`���v2X�Z�l ��,��D`��\��c�o�6�1Ej�䆥��X��qY��ÖҼ��D��@�j)�/\��c�X6V\[�a��#�Y���)hl�qO��G��d�[1#�r�ZM���v�)-f���4HRiD��gMgZ�5NQ��ʘA�بL����m\91Cp�+�Q�i��vѳg<b��+I�h]yKV�\?��y�[���Vf�h�����lU�]��3l�����@��{�k�I^�f���(��G��o<uܾ$��m>'-��t����>O|�.�!M3���F,S\Mkkl�G��]0��մ�ie�k��f0Rn�t��]��ֺV�3l�*R,a+,ڍ�i�eJ*�(��Ƥ�G`�u�j(Cm�-
�s4ۜ��*�ѺhT1�c�Q0U0�h�l��em���Y�&\��V:6l�Q�9�*r�i���?-����]���.���KtV0S1-����m�V`�߇�'��<���T&�O3���WzLf��od��(���ȶӵ14����2d�i�l��'�=7�d���[F{ԙ��۱S]�y����9j:�Ut�
�G5t��xjol6Jv�wcHVlO��|x�^���{���z�V6<Nw��ݵ�MT��S��˹�Vն��؅z���A�{1z���l��ei��V/S�[Oh���H ݖ-��[2�bxM������c���nf{'�ܠ�m
��o����W��8�Jwp]9z�H�D`�\��ғ�]H�M.tY��Y���2����y������Z3|�/�}���d�u����l<Nw!,X��i�]]��g2ص�ދ�+��u�GN�ѓ��oV|���M�R��{�up$��OP3ܮ��c�����ݸ�|6��S_�e���L���HU!�T���}��f��e5���U�u��y��5��_�d�^��`��/:�"z3�M�Od�kI�کKy�������5eMS��1��H*����qݢ���sͧ��
�DۯL�Aq8�ҢA�41�ӳ�.y�&�b՘��m�=>����w�滖t�h}o=׾��������1��OE��fm�f��j,��.]EqxvI9wU@�ã=l�j��������D����C���f��b��t��͖8V�6�Qj����/��g�=i�;��w
 �p/"Ff�'w��Fm5l3� �������ٙ�X�]��jqEC�f���_2 ���u*�Ckw�	�1'��j}����v�9���3��yﺥv5>'�!(L�@bC'��޼����n������]�t8ݶ-�F�^��@��0�I��yѝT�{/��n�^��)�[̩��$[Cbz�=w��]�2k�jB4�T�^ñ�np�e���T.cv��o�*�__o��5�"���}��tWK{\���45�6�@��ֽ�&p�׆f�����M�O~��z�Ry>��^���}ɻ�\n+.!^�����֎C7���h��;;��q��ϾM�M]�/9���N��|�	��H�}}T*d���k&�C
լr����л��w���F�:��x^���ͪ�g��d5d��x[�&��7�N�����9˨�� �����Wh�7�c�����Ti���h`7��h�ӇY3�~ؽ˼q��j�������j��**��������X�����[1ݏ6��wbM��"2{�i��g���D���w���D�Ӫj�P�7ӡѬ�!��w��>2�|>r�6�n1UѲ���A�De��G[��msC���dӼ�n����e�lG9��-��V6E�k�5yy�R��n̋@{n%�"Q%�;fH��*���1�y��zn���|ȶ��C:���9�4"Bb�$l2��ؽY������N�c�?��/{ԗF_�Zw�� ��I�$�m�*�>�`*�^�
���|ZvD6c�n�{��;�U��=R�
�"'�*tg�s�@�l�!r�z�6�^�z!��${f��Ώw�̌��M��{������e8����CN.��S;�(�1{�GY�O��ֽ}Y>��k=����Z���-��/�{5p__iC���}�(�9�|2В��Q��N�T�k���FغVa3dZ��(J+��-56?NI��,���w�`z}�f͡�Nn�1�;�K�X--��"�ùDV�A��e����e�Yp��2�˔�^]�;m����	I�3�]���F:vZ�l^�Q��ԃ.���,e���E˱wi���A�],lQ���/7JnBЛm�PVR3`�.��[��@�h�38�x�$�0�;�w�5�����֘n+t�u���`k�����D��}��S��;]�{Ny�ԗ@\4ox�s����y�e�%���]��"�4�(�2׼�'��'�u���s���׎�4Z3�F���ɳm�w$.H�MUJ�:k��E��iJ���W����v��U +�[���Ќ�{����/�U �㽂ot����t;ep�Y�	K�.㺦eo�)\f��4��,�p ���-l�ȻYę����U��x�5=��hK�.��vY�c�9�U>x�y 	e;�ϞK����s53n��R�Py��,�=e36i�򌄠<qQwd����^�|������W�+�w����mZonx^8�g����4���@���FǸvɘy�F�.Jٶw��=FsN�^�� 9&�~�&0u�m!gd�7D��<�K��o2i�3e���f��fe����U�	��q���o�_��]�
I��B�_5{�T��$�yǚ�۞2� �+�/e?��x�m_�T�����|7SCf8L��6f�"=Q;T��Jcŝ�U*ڻ�>��#3��g.gJ�{�������n���UW][瑞�_T�����<���e&�,�*�o�F�b$ą�,�d�\�V�ۄ���C��A��1�����M`�:j����B��)�B.�Čl�u/�ށ���0d���ϫ������i��F!.'���ޖ�\�ّL����'ݖ6�*��}��)����K��J�k�^s7���<;�[z���ƾ!MiU�,�}����/6P;��զ�W��3.��l��2�z��w��*z����g<W�^e�vk	i5�����ʂE�����$&��
��y�p�G��/�"��R�w�`<� �����V=7���w{��e_lS���]&��g����ho)l�3�ZI7p�Fb�בk4���r)��k{�{�|:s��NeS��1i3�lǦ�>�[��1
�pP!��Q�A�~@��qbij���\X�ܚ8ưD��矿O<=~��]�Mw�Po���z�th��qy����zY��ǒK��]�宐��n�Ǳi��Ǖ�/�,�Xɕ]��b�͇ō�`�w�=��L�{W�ݝ�Q�����n7���t\�V�U��BM:��&���ߙ�D�#I��E||�Lʀ�L��xb�BH"F@p���a�j+�.�D�n�bw4�2c�t����9w�VP�ײ|���Mp�W^b���2P�;uȭc7slM���(H���Q�g�Z���J�ꝛ�\�s;:���ў�RHvB��ǖA�;�c�/�Zd�.�{p���R����G!`����`X�/bS����x��:��7w�~�B��dK߻�~��i�P	�B���ZZ��aS�Chc �(E�d��J�F(*�H�� |�sy�S�`8 1!���s��U���s#1�U��_>���u��Y��`�ߺ7�)�=�͠[����U=q����!J���K�� �ks(�9�ؚ\�,.SB�J񊣱dMQ)���8n�mkN�.�TM�(��YYY��^�*�]�$��fku}���J�XK��;fy��Y�vN`�ޮ�9|Z�5���2D{��9�w(�A�C��B�1aw�׬��OxɯFi�5]��I�ZH[]�8	9��+���@|�Ԅ�j�2���I���"��[�����n����+�d�6�o5ٻ�w��ta����u�����%���cF8��8�B�j�Z�ޡ�5ûx_S��Ij�j�yp_�y���\*�~&b�b���&#ݬ=�U>+OG�o�j]c�Ww�Ŭ���~���! ��>�$�������y��{��p],�Jӵ4�k<�Rh�B�f[����X���f�Wk��:O�9 y�������U�F[.l*�Ja#��%��RlP,�a�5��l6yɪ1�4������[ej1���b*;q��5�����K-��1J���]-�e ��L���Jȵ4�����`����.�0�[�V�����۵�"�A��4���66�6��V��\ioh歈1��w��{���,G�6�l�&�l���r�I����Av������_�X��
�������SU�m��'�xKi�5�aij�0�M�Y�qF��n�M�͞ʗ~�y��F����z������6	�.�Rj�i��yD��З��0f��ǧ��n1� .Ƴ���)����P��{��`�5��-�:4ܼ~�5U]���e����r�h��4�m�k��PR�M�-���Y��]U�浏R���{��O�l�g76ޝ�(f!xUǣ�_�s�ϐ��h��y�)�?f�c����Ẍ.��ajTV���1w0a;�J�$�t�iC���U!��oFw��:@��l��p�Qn2нI�U+�"�p��z�W�����]�h.-��<2f�E��p����=����ӗ�7�|3��%�h� ӓ����r�ߵ��ao��?$�4��R8�?���M��U�=�����U�ᔘ]S;Μ�|e
�������$f���g�׷d���+GfW�!�������T1����y$Rɔ����u���.s�AWt�Y&�X�\GF_�m���F=���{i�{ŕI �}l�$��V�w���<��Bu��f����j��x�v��Mk�����F�K�H�q{:�z5�s-v}{������m���D�mQ�˖QiuHL�+�\k@0�(��vg�mh��ӳ�9��S��a��o����n�V��I��)���i��a�
��I��1�s���앯|�e�iĘ����/'�o�ƶ�x��.	sQU�m�̞�Dl��ŷN=��1�޷�5!����dȱ�oo����&<t]�)���L�D��ۓ���Y�R��<�5����0q����J{緘�qL�?w��״������L��w�{�B4�▿<M���<}�J[�b훞8y��:�<��y{�n�y�����{����fv�z��gE��qz�燳�읹�@aw�5��9�;���h�o_o��Qڑ4ؽ��/{ۤPװ[/^�u�9g�rK�=��܎o���c�:vU�����%���^�/��=)�v���;j�� ���϶����W��<�z�A������wV/�0�S�^�p��z��זy]���O,>�`|G��}�*i�gf� �����{8{�9�i�ԧ�l�C��y�����,�ɯo�M�"�z��)���W�גw����j}oa�Y����ր�w��v�;�|���|���p�PSɅ�X���!�1��=Y<v����w/���rM���g�e�ܡ�w�,/G��Z�g�Mw.wi�:y�������9Շ��s���������}�/!'�������w�����ml/z^�����lb��ws�j�'E�m���$I�*n��Y��������}��|�flI-&?Lk���FÆ!�Dc�1=�̊��s�M���g<�鴽�kut�+Y�X^�M[7��w�u��Zk��Π�Lg-Qj�tR���1�큤������k���1`xͥN��7N.YSiX-E̳7�M�ΡƧP�[FQ� �0Y��@�^�x��{�ӝ�ބ��T�y�u��hm-�t" �o2�z��b�&02�}h��:xu#ǧ_�ooooo���>�=>��%����Z�QeM@�B����vA���>>������?O���3���| 6�b�+
���Ieb�0L���PRQ3
,�L�O������ӳ�}>�fO����r�J�G)��)KbZ�W=*A�
���ŋ*|��Mg.E0h��(2̛�����������c2}>�j��>`V.�aZ�����5�,�4�Z]I2�!I==�����������3ӻ���f��5h������DCL��֐>�N5�[[z�{s��^��_�����N����#�8A�s��Pq,��Z�nPQ�D�>e�kF/Z��*�ke1"��[Uj�E*UAdFE�\��rX,�F��%�4�ũU"ůd�h��Wn& ��o���Z��(�X=j )�t�p�Q@V ��[d���U|����|E#�Ć$58`0̀w���0�������PB�`�"��������׻�*�5RȬ����q�s=��)�^������mh�lb���1w��2A��|���J8��y��?q>�*��/�`�YN���&�}���}��" ." ��Ao ]-]t�::U2�������:���3�����|�韾��U{����L)���Mt��bb7Zoj�X��m奮�;+��/���6=Tf�=]�	���f@v�Oz�Pre�KL��g�J��bqj�1̚�z =�>GeZ�z�{D��9}�D�h[Y榁���女#һ�v�����������i��{+;�T�S����x�G�΃��m���������~bypk6~H�8�et�XSjvn����~[��?g��Q�vl��!�8�;�|�F a��/n{f�y��f��I?���H��d�E��݉V�_�ke;f$��CUT��r �6��Q���r�T]���v�h˛u�A03��>�&�\�X�}y)��ܲ�f6.�C�3͜���:m`��q�K��|��s7cOkCS��ٝ�p��{�*�9|%�fn���pɲt����N�`�ȴ!v`#s y�j��*�3��곀��2�>���Ԡ��I���-�v��dGElӘ����j}Qw�<ѹ͐�B�+��l�R����?ji��N�o֣������t�r-ohڸm�hj�xMmw	���������8��s7�T�V{�1m�g�̆���C�DO�~�z�;�O^�f�%j�i�p~���]�*^)~`���8�'��gul��*���FI��v��оs�t�fC��m�8���&cA}Nta�6�\!�F}X2���:�l�t�D��^���P�e���D�H�i)JNz������S��x���4�bݮ�f��݂�f��r:V�,����K7Z����r��f���k5����M)X⤴WK�c���Q+�kep�,U&���Y�lXJ.ұ `炒�B�ZL��#�x7sW�G1�!�1+jC7!�.)�\,4�i�ۥ8p����t���`#�����P~�̵#����W:1���GA�2��MR�f"��}w�6��-w,�~���=Yu�r��q/l�B>ɚC95�m�k�+I�f!0�3Y�qwN�=Ԛ��3�^]�n�\�O�r��Phd+�`��V�<>�Έ-~v�kg� �=mY�%5]��٘�ݔfȗ�K3}�QuY�6��Z�K�	 V6<�G�IC�ʡK����bfW>���es�k��;]�e@�=orqy�jAa$�fB2Y�;Z@P'�m�9,G�o1�y��K�K�r�x4�j��W}�}��s�?����Q���dh��>��>_��b]�g\����/��n嘔��� �-{.>�{�o����ٝ��.뷦�>q�Pg�bA69�t�}lǦ����������������6_6�����<ÿ�[w+�z���w^ԺP�����g��Y�(9�1�/��
+tm��r0������nw\��k�OtB$����,��q1��S��W9|�hij�us>����w��rH>�d�o75M,k�w�sҢo�K�J�/tRv3j���5l���w�g�p7������������k�h�}��r�w^m-����L�{��c��R���c��,�
���5����q�y���-��[�C?bk�����w=7.	/�Z�p��
m�V���lY�[e��-Y�l6�&�>z?P��b.�Ǖ{oȿL�q��ᴣ���ԡ��;�q�=����Ҹ��\�D�-�B�՛0e�y˃�]v�N�Ш�a���k&���My�n�[@2��6�9������^g,��9OIS�8�;�<���7PaFvo �k���>8�U�!��*R`�x6�ʅ�����s����U;qɨ�j��y�j�P^C��p|��ML��v�u{��_�W��ww8�=�;��X����$�v���OU�ZQ��'M�Ї�Ӽ2-�y�T1}�9L3-�5��WAA(%>�p�u^VW[7��Jg6̖lb%q�o9"�`�W�: ������h[��v��^��u�z�:KĹ����s8	�<�M-F�@�Jںi�,�.��3k���[�3�-6�Wj�\��xfa;�z��j��ihV�m߶�4E-8;&E=珼_&/��T����.�i���WF͛7�t��qT�b�C2.3N��Γ͵U�w>���q�c_�:e���g���^�8�~.z���2�{Xt���^_>"�7��_�4����|)���J�S����
�e��P-n��
�n�������F!�.����l��KT�zE��{	�#�<M�B$�o^���>��s�U�]�LMSÍ+]�uTO��wK���%��ދ@��Z۲m�h���c�C"����R��nup��>O���~y4s��l^q|��gc�r�Y���y�f��(��r
�b`L�C;fy����kM�s�_���Γ�e0�-2z�例�wg�oD�)��cN��LφD��e_"�������L�̯O�@��K�fAX��nd�;x������d�x����Z��(�!÷�}n�	�t�#"�N8P¦�Gm��"a�c*���S���誜�8�ǀ����4ʪA��Ov_�ܨ�l��7!\쬨�E�-G��=��K�����4�,�c��'���6{����$��2�x�����O�!ذ�[�4@���%FW# �ۖh�Чkֆ����*���>rp����<	��i�Ib��F۴�bƢ��0m
��4�����e�5��L��֙�w"�f�5�n�2Ө�PR[Q&n�ѵ���+�},eZȱHɑ%�f�묹������B�����l�K����J�`L�\�A�-y�cFR�.2)eюڷ�����ys@ʰ��0���7������X]��V95Td��U��k���	�T����ɯ�Y�ߟ��A1�<s3<W���r������	l����jh�
B�����F�v�����V��qYw=�^��v��{재 E�{a�R�>��/�_N4h���X��R=����Kg�L�;S	�[=R޾su=�s�y�<�TL4���'�W-�jbӏ_z���ь`�GZLm��ŠV�H%��6�K2 �}�:T�f��J�z[8��E��W6;!Q1r�d���F�t�� �x���=����'�d"��c�\f��k6��e����5g1L�K/��<�����5LE���Ľ�|�9���z*b$�6�k<�e�$�ij/G���xG�B��S���욛��mT.��~�ű��6�fY���ަŝw�$=���)�p�^��Hb�����ʍY��\'cÞ�����gnjv�l�>�W�l�q� �� &\1������}" �>p�EY�9WR��,�MT�)	�%�������7��� �T��7�Kީ�Σ-��)fg�����Zk�5OD
���8��i��n�Eٛ��NǇ>۷0Ԅ�D�(<����ecŰ�0S�� B!	�;�=���ٰaW�Bk��em�3L�)6�$�c���}�V�xD�C��z�V�Ƚ��ݰ&|�,�En��gc11�����*9�e�^�/ܗ�UO�G:���:#8��^:�u�@��[Sf �ʖ,x�^����*(�ӓoњTh�X`+��JPڽ��xL^���d�5�r�M;�x���Mf�暒�^�w�ڡ�}�>�r��e�����3f5G��-d�F�KKC]W��o��߶y�-+m[�`by��8�|�=�f���u�&�9W�?c���#�4��5 �F$���L.��ʛX��R��s�2�v�+�%'�%��~���\�G��\ݰp`�2ݨBU������~}����(c�>����:v��s�:)�����l����<	8����wx�Ѭ:�ᮜ?T����.�}�-w��]b�nd@ �kC�F8m�3z�$c�bs���/��>X�.�������d��Cl�ai����K+�#Z�^�1�!� ��VrY�3æ��j��X�e��E�J��J#uҜ6��*��ص�'�I\��}�ߵF�%�%�O�,��~+������9Y<|t{��J�K��"�D�8����'�W�(�p9�Y�N]�y�|�R-sG[ow"���o�ު@L�?1���zg�e�o;�K_6�T�Ri),�������e洵區��F��*64E�$H]Z�GTx�L>U;E(ݼ�����ꥐ�z�\U�{��t;;�K9��5�]�Nw��C�x�C<��Mn�W܅7�6��3/ؖt���Z�g	�+Sa�-�۸�X�R��!�f�s���x�S]�cF_oQ�*e�v��5$"�I||V
�x�"<�1��x^���^u�Tg��� �1q8Sm�Ar�'[6�6�jgo'\_Y^�Qk�����&xu���,��!5U�p*�2�5#A�p��C��o���|��1�w���� S((D���9�!�Nph����A�W�&�jt-*�p5R����*�� ��j}լ�',���ث���%�{�����#�v��<��=C���@f�i�����x�{e:�-�.h9<�op�������<����>��췈��wy{}=xc��"C�����V�����m�+�D���Y��%�w���jKo�q��h�  ��K��67z�bϷF)�ϔ>ȋ��ݷ;n�~���;(�
���p�8����x �y��t�����VS�)�+�.���n^���<6�l����~ȹ���:]بm��3�ӺQ���iq�~���V����2z���T�w_ x���̩yz�Kk��
'����sr��.SL�X,ʻb��x���Y�Cms���o*��b�n�K��ط)Z�]�=ݬ J;3�����ܦv#�����W��K�ŏ���ϫS�re��B9c[�����'ډ�^@�{Χ��c��x�Z�qjEg��+���k|:#�D+� ����(U�ˊv��}�����u�(�Ł�k��x�������.�=�Y�t���{�t�1F5f���#�����$c�üp��=����~5aI�v� �4�<���9a��閲'ڛzkJB�J��eD�eW��˻�F7���6	`7��Ṹ�e˵��{q,��p�=$��~[�C�|��e���D�m�ŞY�;pF����Z�������Է��)���[G���i�u\��U�L� � 4�G��4�m�q0p=`�P��sq�y�K�UC
25�m�*��Y�S�gk3�|�H�g�@��܅c#6��&��-�p�M0B'ƴ�K5D�Q�"O�pv�5�
Ԙ�XO���`Y�.�r�m(��m0
��� 6���%V�	�i!0e����X0%�{s؍����im{&'��z���.�yt"��,���+��ȏɉ��i�B��9,���Ƿ�������ï��N��}J��325�ZTD���X�t��aY
�!Y��de���MMMMMN�'��}̟}�h�(4lU+S�!����QR'�������������������c2y߽>�QdQt�@mS�L��"�%UB�Ef�Vj��zz||{{{{{}}~3��3���ZD�Z2�AI�r��*(ꅊ��m��Y���jjjji��~3��3Ө{U1Q[��.JZ��e�PQ`��(��xu3=>=��=������ξ�=;�3��ϳ0uES�pT*�F��Y**8�[l\�Z�G�����U�)XVUb�j��A�e�+�e8�S���E�U�PGE"�X�0h�+E��1�[P�X#{s(�F��`��%�D<��"�ZX���0H@�+���Gm�c޾��������%��ߏ]�X\�Quj��1�-v�֘.�ִ����ŵ����Y�V�d�ؐj+u��h�0�Kv���.��6R�h
�m���caa SWh%ALgRQYtÍ%o!a����H[s���k5���Kfe8.��GM��K0��-rM��+,$6Ś�ЭW���(Zu`Y`f�U��gR�%�KVݦYR��m�drpKac1̻�k�B`�mUj��!��h���-�X���(�,�9Y0����pk�y����p �%�ͭ�.
6�Ȏf,�����3��u��k�����k���21�k1�f[q�nu��v�FY��8Ҧi�Y0ٍ��C8�tG�P����/b0�1�-�K���4�b��尃Cg�1Iw6���D�IM�6�;b�V�]��:�˫��ڠ�2���3,{�4�Z�@�Y[����dog�ˣnFh͜"�b�6[�CkK	�j�ՙH� 0��gJ^�.:���2ћ��Y�)x@��v
ᩇkZ�\�Ȉ�6�6ҕ� �%�����⃱�sM���c�%��l�����d	4U�a��cX�XS"h��Cm���K���M-F���e͒�B��S2�öxMf��';�R�j�إ�-.�H]n,�A�� �WXg%�ciiz��6-��4Jb)���@4X��2*(�5Ki\f��e�l"���n�S��%��ݵ���H��54u�6s���V�5�kqp%im�Rd+�Z75�[m�����8�t5#�e4�l���W�e�2G�0˯��w�<�xv�e��鮯Sn��{DC;�&Jo�14�mr��<ޅ���:�T�*���Y\s`a��&¬h]��h]�f�X�RdH�.�A��B��Q�bdo(]�m��6M.l-�`��@��̱۝n��H�6���&U�jvl6Տg26Ű�6�%{@�K[4n��V���E���5�X�s���Y]	Sl���<��/�e�t+��XEҔL�TUh��j눡���qB�6� �\Ŏ�9"e^幭�Ml��wc��w:�w�z���3�ggz��3�ӻ��U�a���C>S��`�=���y������{��HO9���7z�&����P��.�C�B:�����׸;d�$��gu���Z��Nɷ]�c�����r�W�;c�0O��o&4��0c�ȱ�|���S!)i)��	�t=�Û!���'�~�U50��i��D�g��c���C���Y(X	����]E4m���sm�aUr
F�%�Zu1�&fch{*�r����{��iC�.���,[�����<��\ݤ>ꆙ��f�*��R���s���RC��Y���3��yb���8�	=��F�N㪹{7뭱p�^S�k�< m!�C�W4zY�/��ϼ:�Gh@*���/�,( �^�A�v����K���o��"oj����n����K��h;L3����a�Tg3��+�0$ώ���yO�o8d�;fTF����3ϚzЫ�� .��S^Lk�kCX�z��zjwT�]�(�ci�BL��d���z��Vhz�~/ߖc1�kMp�嬪8�����e�֐{!g1H���,��ҥD���ö��5�<ۓ��b��I�LΒaDn��*1�4ݧ;Zzp^��~�y�d{cDM��`�P��b=X�Ay����1d�[b�y�fF����7���`�N���#8�x<�T����{�_���O��^b=˷��(�)�r����HHb�t��dq<+'x�ɏo4ҷM2�vv��/�Dx�����Z%���5*�oJ��7}�5D�scM�@L��r�{�o_:{��u!FsULS"Y XR^����SՎ�^m �M��O�m6c��hhJP�7�~����5u�
�J
�8O_��������c͖g@ZU���e������K.�y��1<Y	�VI0�Sn���9���z{��#�n���?Yj|�$�@Lj��i���B+Ă��m3�4G���S��42��iN����j�-����l�VyMO��U fK;	�	�����f�1���(O�/3���R�Bd��eeQH,rq�������!]xs�˔��6C����=p�L�7���~�ݛ������۔.��='��v�����]#���x���c���,�X·Gt�]`���|���'v#�9�٭�A ̇2�����O�g�w�4Fo������p+��v36#F�[�éL'������o�@f�m͸�\�3�]a�8����7�k�%�
9���uشˉ=�"�����o3�|'���i��I�X%�G�b��I�9jHA��uy_�l��np>So��W6�d{j��+5m�ìR���@O��S!Le�P�����F{�xD�wϩ�s�K�	��8��l�P*����>���*P��}c����c4g�Gt���َ���ghTLMN泖M��5 �Jص�mp��Gy1�6�#�7{���a��.����5�.�����ݴ>�]e���q��=���Czjǽz*tD���/z�0�^���S�gB�Ч�=�}-������C�Dd���k~=�:���͡c�
&P�30�ā���Q%��-��7Bm�^w�TT�tKI�vp'|q<�6R��M]d��A]2[�3n1�+6�F�ַ7n���`����2�k�sm-Zq1U��1v7�Sq�ʫ�J\bgB�gj��Yt�ɮ)Fͭ��Cik19�v���9e�W)�lJFY��J�խ0�	���e��&�0�ѡ΍�ű!��GMwƣ[�7�������/7Rה5�e^�adh]:�Ἢf��ߎ�g��7��d��N5z�h}��}OC<[X��n�a��;&�%�Y҆^u�o
�?����f��X:z�.���
��ǂ'�J��N��o������y�_�0�w�t���B�6���|���"�i�f�G����T��^��ϬZ�R�RQWc��wtjx���=6{��{,�{�j��A���b��1i�1sJ{o���{4t���Z=]Uyى����6W�|��{�~}6��,�W��O-�=��f��.Ckn8f�.FU�W�dMtn�qf�ŷ�8�a<����p�,����sp��z1Cɐ&+"ek*qT�`�П^u^�8j�%�P%ť��YF�R��������3���5K]飴O'���gGR����2�d���{ss����S�+� ����0�6���9{��u�\
�1�-��eϬw`�n_Z���(L���d���!�<v�ܳƺb��s5�p-�=$*��G�A+�O�S=N_��G��N(b�V�3�O>N������%�N�X���C��<��w��D��Ì��2
$��%�{�^��Ջ��''<L�W!$K�����j����f<D��0��_��-�%�)k���9����a��aᣒ�&�AJ��G�cH!��)��p��w��s�]���\O����K ���B�l�����������_MS}����ӺR���,�v�*��NR�������
���Ϋ�>��j���,aا��A|��0��֮6Ok��.Ð�S����λ���>���U������e��A��Ȇy������q�H��K,cؚ�UK9���]�U�����U���55y���,�S���H��y���X�DI��S�N���~7��9>��e���B�i�Mx�X�ٮ����a-]+��ߜ�5��Gc8���d��-�m72�����1S��<�]�����8{ν��8�.3�ƹ�kژ�8�OM�}gݲP+��Mk�ݞ{m=��(��`�Ϳ?'���	�8f;0,f�� \�C5��b������1כb*�3ѧ!fD������/��0����L3�)	�+X����Ye�Yb}h�>z���{��q�]���O�s&�B��v�A��=�ѐ����=�v/5�R���7�:/�Q��:��Ǆ��7�����-��\FB�f�t;�0�70�S� ���jN� v!<I8�!����;�2{&���5{���|����y��*�8�ۉ"fg�7^{�n�+��'p�ﯗ���Ѩ*]�73��fi*;:�K���
�n�e���l ��o;��'�����0�۞��Jq�u�4Cp!�B��[���M!��e��ί5t+#Խ�5�u��:�L���N:i�+t�<ݸ�Wb��v�$��v�e &	��s�.r���z諱�*��M�z@SH;E87;��Q��ǽ.,�)g���ȼ~;:ݔ4C���Dm���Zi�i�SE���ϚM���Y�[KlCޯi�?��Բ�s��yb:ЮpA{�^:��q'���>�aMj�|s{He��x���Uk\�=�7B�j菼U���ȍ�����N͵w�nPc�Ğ��KܾޔF0ha|��o�z}6%J����t���Bi�I��9�����
�Q���.�Rm�� �fJfM�F���.�3Z�lT�"،���]3�&m&I���Qf#D,[�L��0С,�F�@f�3,���-bV�K�u�.e�;d�:iN�6�m��H�M���Xe��l��["�i��4��%�]��+��s1��M)
F#�=����e�KL����j�`���T�PN.�Z� ϾO9 gKs@T��`z��K���l�RZF��n��J�ѨL�nk��z�U�4��v�,��ͽ�'C�n9�1�Ú���Q�]ף��J�A��3EsS&5���sí���7�3���,����K���Z�ٞj�)�c��}�י#w�0�OU�p����������r�Z���M���ſL�>Kα4���{��z_.Ll�	�a�0k��9Oݽ�A��Ծi�����lR�X��Yx�X҇%���<rP�ec;v�v���F�#u�ϗQb�*uB��l2��o@�Z��kl5�F��ա�>�T\��C��.��yf1U}���.�sV��:�*;��Oל��s}=zl{�ŋ�QQ�hȢ������*E"�<%9<ߓ�-5��/ջ��z�41�S�C%
JC���`X���J��J֪�
����&���;)����h>��ȩQ2ɜ'3'C�WY���o;�q2��lfJ���t�2}��	������n����FV�q)ç��"�aE�20ܹ[��9�=&�����=w�w��v��fY�Pu�]�ڪO���u��+�s)1.P �/���>���gT҅�ԅ�hJƎ!3b�#R�Rc4�yJ�������"]Vz��7}������-hVG������Drzkp�1w(=K��#-H 9�e��4/�_<?fS���2�b߶6�X}�2��gYۚ�hFη�����d�`��x������S���j���L��9Ç*�wb�:���|�Q�|��-w�^�� <�
���b#��ד�"�����׾>E����~K9[�u�X�@��i���p {�Ѵ�	��^�viY�|,͂�o��j���s��ѥ؎��a�)�^�M�1��qٷ���{�HDy����\Ӹ���M�su�i�
����vF�V�l��O
�����{����&c7<�v�{C��b�ݤ�<Ҏ�c݇���r{�}����x�*&׽��ײ{�t�{�}��qW��\�����$���$�=��N�z�u{�?j�w��C����E���{vw��D���f�*k�'�P�/O�����ĺ!4��^�s����{���x�y۴�کd�`ox�<*��;[����:��X	*�K*m�볷wH�����p����:�R]�|F�����7i�'����{p�f{@�8�`�9t\V.�n4��L���N�]'���S����Sӵ�6�
n�o��{d��6�M�s�x]ʽ��RWr�{J��$9�k���2x܂��n���|�č.��wxg�F�,��`�Nj/)95$X�.{5[���>�S�1K鏁z���U��ݴ���\�r*�l��� &h�$&HI6�t4^�ٌ��Qx�nrp��V[�}K0zD�A�0 ��j���i�Qq%3Y0V���[V.�x�~��ڊ�*��(��g��ӏ�oooo��>�}\�z|�QkYQ�*��UghQg�V�W�+�{���X�ho54�4445��md��v�yb	���U~�|�\DQD����"��UUQf �i�S�1�r��x�믏ooon�L���}zwуTT���=�mj�*�Lʃh�U�ޮ����1�2jnnjjjj}<��Y�>�=��f��KJz�L+j�Uۈ`�1E�1�l~�H�E��=��>=�������\�z=��4��Db*�AL��SMl���Qm�j���0�ٓQ�����������Fy,��L���<#E)�eX�e�n&�i�h"b����9l	YAX-�*����B�(��j�V�	�A�UQ�T�ki��Ҍk*�>����ye�DV�p��_��b��P^�պy���c���s<�F��tdGCv�P��nW�\�"�YUR�#E�DE�+T2������Կĕ&�����}�^s�ΛM$L�82�m$���#-��d�79�mhoS�M*��sU�A��m|�����I��[�#�%�Rf^��tߒ�oc�������/}���"PhIi�rr!�L{�ؕ0�p�XVz�Y����ˡaiW]5#u��9A��$3�����Z�R y��MB�����Z��}�x����^=��˃�\��LŐ�S1k�A�����&���|��psھ�xL_p-Je4Ϸ�>u~/���Ch�UV�Iq'���~�o�z��R�u7쥞h�=�s�����T��@�ײ'2���dנ��}����y�mv�pAݷ[��_�fB%��^��w����p�ࣞO�*���>(����{�#�r�^��̨��L�n�ܚw��?�E�|ܻ�W�����l��E��{@����8��x��������ʨy���K�x[���	�p�)m	N^������q����c��m�F�FbqC�0���D��:�s��j:��I�n�::_e,���f�#G�SRPǫ�iM!�L��"��T��zk {�;6�i��y�,G+�Dn�.l�o\�k9�H c�-oM�
Т*����.�Q{���tx/�θM��d8���I�)�Ik�����Ec����"qs�qwT���5�U���*�n�d����,�%��\5����UW�y��4���k�c����0Fi4ėgtnvx��j��$��ˢmbk��<�;��Jc��/����yH�ۅ�Xy���m�=�~:�::S�e9����,X�+"C� #�rQ2`�F�i�9���em�2�u%)����i�~	�A%ͪ-��¹�I����)1si]MWh�2ש�/A�t&�;����˶���&�E�j����9��)�A�c ��&��02ʖ�6��mښ3˕�nf�eq�Tj�.F���:<�8u�J9�QkI�͵�2��a	Z�<qq�d��Q���k�F*�ޥ��������C]M��"�n�nds�%+Sr�p��:��$g�э;"�b��V�tg�B��̙gf9cC�a���K8�����T����ɰeo?�l�����̎؋�W}�\Kg��%�5v�%���g���}���x�
�2NgN��]��j��Ά�q&�T��d�E�R<�G�mϳu��l�=���ܻ�W���3��1�{��|��56��@�)5W�6���{�G{®}���Wu�R2�C�����,��Ļ��ڿi�t��}���Jp�"Pu\(�"m�ĳRcT33�K3���$��
"�lh�B�˱;�Ѫ9�]�t-Qy~��:�tɈ��t[	�����oH����:��mna���s�;�v�&iޘ�����������s�ŋ�w����T�v����y5��o�ֽp{���Z?�z�āc������/D_zJ���dD��9j��mBl�q8-3Z�Ʉ�n��7^�c�ϑW���g
�óX�@KZ��E��>��Gr�k-�)3H�0�o4�����}R�u��ii��m�N�sּ���w�d��Ml�zq��@�g�r�<fl�:����)�g4�j�[����a�o��ۘ�q�;�h�M�#����$�#���4�%�K�@�t�1w�ר��r����&2���0AJ]�������w1�#2LC�^��Mڤ�D�D��"z�=9�\m�B.��4��X��c��î�;^p�F�E� ��6�/*W�7�� �o�A��dHte�Se�>��I�w1�sΦ�7/�t�t�gT��R�ß�N��?�'������]Q������o�I/Q&�=R�����b@bτ�WyJ^7}:�Fx�H) L�Nm��H9E���w��n�j79�
vL���2�q?nqOW©�Ջ�x�z3d��-����N5�y����C<[��~��Ns��܋��u�xu��M�y��������t��r���-2Q�,l��p���L=�/����h�⛁W�,�3�m�]��ٌ�$���O�#���la���
�U;�E�o��}�K%��ރz����$ܵo�@�x�ݖ�5�#պs�t�u|m�p�y�~ ����������gk���\�=�C{+1��z{����պ�<:�󄁊@"e
cU�qb#����Z�6��ɽ�.y_V�}���^��G0�%.29�x��M:u�iD���_����uk�{R����O�{��^~O�{{}t���R��]`q����OA�FI�Y�?����0=�igrs���o��+3qr����a�vT�������5[o�����^B�5{i m�]���_�O���X,v`��l�4c��E��\�QH�v)	@�n<�
�O�C��c���]w�YÜy�Ǯ<�L�>@E!,��I�GG�O�Z �=��7Fז�d�S7����jS.*�	�ky���H�ZZ���MZ��I��-U��U#|;ϔ���tO6s4�mi3�Z��������gw�z;ލ����[�R�Y�@����D���1k;F\LvLֽs�gI��a4�(�e�TMU���Ǘ��G���^�'���K2=~
&�5�S0Z�f����ծpEFtG������g�d�N|2�jc*�����"6�}&pFɏL���\��G��n�--�1!��D�k+����/!�D���X��2�u9qD���VH�8?'�R~�4c����F�h]{U`K��+I��si
J,����)�dR��'<��yg/7�O�8��2ʹk5��3j	������6c��C��Q�e]��6�FK��vP���u�Z��[`1�`&��J�&��F+C6���X˝UDc�V�)bJ�s0h1v�%n�)-�)*�H`֛ YU��5�]oeKK��c: N�uZ�&Ñ���!��F�m�[��?}��4��K%I��٥�����p��!�t�%�U�T�2�1]\�xr�����g����5�y�g����U6p��C[i��kǝx<I����l��ӷ���z�^�@LI��}SQ�E�S{���q�U2��̻X��ٟEA�9"�i�7ء��}$�­\�+�gl��6<_TB�dǇ�>�q3Wj����jg���M�h���nyr�P�>��R��!��l��{@4�3Fk#��Z��LcUH��\���� �M4QI��s�ܥN��c׬`E������,3uBm���������l3���]�v�`F7kiK�5�da��{.�ϼ����ꅤe�5e��Ǉ���'���r/��'�Z`���]����KL�L�O�9��ËR��0���.���i�1�%�Ԏ��3��G�R�z�<��cX�znm�Go�=�s�컡�Y��8�
��$��~d+v�̳�ҿ=to�7�9�'��[������~�w)�IΎ ]�2��ۓ�z�uEׄ��]�O�y��m!�6ZŠX�U:pA�S��0Nq���9�ܗ�en��k�M�!]߸sE��Yi�=�:D���v�Lj*��s���U����b��{�=��n��Z���U��C�=%��D���ˈA�	0ۦ�h��i%�:X��[��۴�=�6�*��=��iwz�~�����P��;�S]KVñ{k.�i��\3�7�����#�8�v�T,�����{�����M:Yڨlvfi*��<ۭ�x���,QRDəq�,Vz��D˟I�t3=�i�8�Ft�U�����K�O�z�w��}�ݜK�_�\��V|ݽy����W�E )=ֵ����SQ7�sN�>�6�N-��������dWSGr�vXf(vm���]���;`��?{=����@��ql�B�h��S�� �6����=Z+�o���MWe�F���َ�O�3(�&��t 䔠������/�V?S8����m�E3��kFʺHi�(�bN�uM�����0�	�O��V�w��L�7�ۄ��ɴ�o���i:�E1gd��K��FU3�[C=:<��0�w������C��ͿV��z��Qg�,� u��ǌ��������ޛ�3=�& P�Rc&e[�#"�\ʙ,�6��o_sԽH�8�@�-V�4�r�L=�d!ksC����'�Ɣ4����O/���'=7ov�1a`�v�w�O�:�� �I�$�Ds��Ho�g{!1�*��ζ����!	�������3w�Zd҆���쳧&T��s����Fz�o�~C���UإS1R(�a�pC��	y
����ֿ �B�m�-���{�q��{ҫҦjBn��<�P8�ۍ�/wR��v���q����=/5�,k��W����p��\M�TB,nЪ]�gɝ�����b�1t�#f�u^�7��L�fR"fص{�6�O#��v#�L���ޯJ������ɝ��[P�_gS���z�!��M@�PɊ��3c��B��<v���nD<���շ���UY���w��w����_��#��Q^� �*���G�∊�*"�ރ��EK�2p�!��0U�U�	U��E�	E�	E�	E�� �x ���+J,!(�*! �X�P�!"�@�"�@�!* @�
��^`!ڢB!((@�(	�Q���	�$@��!
@����C� 0!"�@����H(�! �@�����B(!  @! @� �@�!
�J�p�  B �	!�  �  BD �P A{`C��( @�! 	�#���X���X������q8 �� ��(���������²#H�!(0!
=u�t���������������������@����
s�!�%!%V!V%   !W�s��A��2����(�**�̨�T������������������O�g����g��������S�����/������?��"�
��?������
� �_A  DC��h}���S�%������Hz* ����?�G�{x������A����'��������\+���  FAZ@V�B�F�Z��F�(UJ��fDi �A��h�F�Z��Q�Ph�!	�bDbA�!E����FF�fQ�IQ��bQ�d	��iFBAbQ��fQ��hFF��$D��i�Y!%��ieY%F$%FH��hFB�!BQ�F	D�h �YFaFD�!�X�`IFF$X���E�$X!%@�`�bE�FD�fQ��ddX�`!Q�E�A�aY�`�a�eXFF��dE�VF�aFF�Q�a`Xa!XV�FHFA�eE�F�b�dY!dZ�e�fA�Fa )F!�a�`Vae�Qb�F�hF�bQd`F�hF�ae�bPb`	F�h�Xd�F�a�hP $�F�B	�h �h�PA��`p�?������UT�DP��QR�@o�t������_�P}�������O������TAW����G�~c���?����������������U��!������$AW�D~��������܀�����=|	 PU�����C��I�a�P��8_ۇ���a���6`v��*������?�* ����P����������~����O���� �
�
��a���
�*��}����)?5�������ρ�O�������$���U�?���	>|?D����~A�~����~��O�>��"�/ؿA��
� ������x�����S���e5���{_^-� ?�s2}p!+��  @         P       �(                c� 
P�R�ED�P ��(
(QEP P(

� T(�	��P(%EP%R
$ ��}J�P����I�
(�*�IU"�)B��U)I%DR�TE!	*ET����B�P����  ���URUB�EA4| 3a� ����A�� / �A�z <�@� L@����@�p*BRQE
�   �
|�:

"��: ��D�^ @ �gE�h(����X z2 ��EA�#�Ӟ�z� ���
��
�  ψ��R
 �P�R���. c� d��� ��� �	��� ��B�  � s�H� wS���¨R�A[�  .)����G �u-�!]�ws�I;۔��܀w���JStTf� �t+����s�҈���(��� ���)�PU� (���\l�P�U{�t(ͪ�Ww�QE���fĪM�C6UnR���rԁ9�@PP�*��}���o��\ڢ�Ñ�v�Y�J��u6�D�P���W���J�n���!���*� �(�� }ITR��*
$JI$�W��  ����=��  �uT%0 ���@7`A݀�uDQ� -�y ��(��� p/�㳾� �*B� ��@ d� 	� �EI\ 3c����@�v 

PN��1JR�D�Q"�EEH�W�'� wX@��� �TW �: n� �`!� i� � � D()AT(Q�  �`!�� v�)Up m��>��ް�� ��T. X���w�+�`��� 5=���4� h�"������� =�L"��  l� JJ�F L%?R�UOT�A0�h�j"f��6�P����~����߿ｿ�I�Cg|�α;A��+uǳ�q4!��@!I:Q��H!	&�	$��!	'��B�BD!$�BC�y��}_ѿ��ƫ��U~<����ɽ�ɵgT����n9���m�v�E�zȧ�pJ��k�3�ە��NC��ٸ�GP���c
ݲ�H����.	�g.�I��zU&�P3��"�a�cvL�I,<�┎5�!aZ��qn����|����M(�� ��~�#����݋EY���v�J~���pPE�U������/���������:����"���r��68ۂ[2ܫ�Ѥ'���s�m�����c��5����a�\^�P���^!��'������� q�6��ڂ��w]���
�:yHs�w����VH�ڂ�fv0F���ky0=<����Vlɻ͙Y��I�_wu�u��
�DƏ��W!����r�l7,��)�Ѯ.��5bc�� ����[�ŦΞs��#�Y����j�cԙØ��5��a��;�z��2��ܥ���;[�$��;n�[�R���9Ҿn�0.�ܛF"�\߲M�&� KV8q#_Bs��+V�
&��n��n�8����z�z��a��7�Δ+�T�hG]=� �A�Ĵ��܀��FB6gnp�ΜՖ4�t�ᯃ��oBt�<�MZɻ������7���R!��U6V�"t�0X������A«�p��Ԥ���>%cG��O3Ku�'qK6��5w����t�L���vn��޻��gV�^��ue�x��l��iը�g@�ss��i&uHpg�$�ؖo	�x۝�
 H5a�|�^��)�lw\נA�$8�H��k`LOnѣZE�M���M�>�z�����z]���>ݕ��8��x>��5������!3���U��f��ж��n
*���I�8.!�ަi|^��j�r�p^�[�֬laFX��Yj.�v����*��0Z�@�q���1`�)�e�����T��M�3�<X�zf��K7�h�^�X�ah��j�~��Z�D<������gm�6J4't�Ï���ܙ���k v�4	P|�vƤW�\AG���~���9B?r}pQX[	�s�&GF�M�G6�Qg����㣹V
�V��6�,�En�߹l܃T���°�=7(w�]�nk�/[�vx(�C�Om��:�Q飃:6wh���[I�ۍ�=���v��B�lV����4�BD��224�]qf��Y�A�5tn�\)I�	y�=[�;)@�5m1`�h�b&���X�NF��^Z����ll�ܲ�.kY�-�kVb��jIZVsCdf2S�Ną��� �M��/0�tY��GC��7�!�\w���q�j#:
ӑ�ۺj#��Z3r>�^�po,�E<&b��r`��9��Ghժ�����Wd@n�)�:O\a��=��ɺ�s;B�0�a޸m«�@:��ǢK]��u�dN���x,��H����qQ�/T��.���j��v��2��bYM�G���ҵ���Y7"�eQר5�;�F֧����3�&�%�zgi���ĳR}���v��ʚ�B��� ��	lӷw.�3�g���SU6w<��Ϡ_�_v\��כF��ۥ���JfM�$,��d*�RY��1��I�;�p
KTJG�O�s�ꎓ�N\}"S{a�]�R����Zc\ZE�$1H*����-�sp�)�\�������2���ʎ:�ɜ�S0RFk���7�+�%������=�����wu�~܏fؖ�a�0E�v׽�*GL����d�`����f�b��ܡd9�ɜ�7ݖdҨ���P]�5l��4�+�Y��9���Q��i���Ղ���5D7uRӠ�Y�>�v��Fs�)0
:��Ng4��c�Pq�n-Z�N�=Tj������]�oD��шNy���KN�;#��S�BӢ:h����xp\K���#�Q��Z�L��N	����u>�S��W+�`h1�xK2-���x���١V�2O�o;�&ǁ��狍����w	�N٥ �Z����Z(�*���-�s��������F[�2n��sD����	]唝A�x��1;��ȷS"Qɰ�4��7 NSۜK�w
W%��C�M��`��l*9s��{n�P�nv���x��l-F�'9�v���,s�M0k�gQ�f�]i�r���(�,�,�u8�' ��:H�8�t�v�q[9Ū��ò��7ElI��;��Ugn�$��0Ꜹۢ��Ú�V�@�{�-ڇS�� g������O���U�ճ��<+]�d#xώh{��ݹ ޥ�wu
�}4Q-�yH[��B]����Cjv��W���
��/�_&fFū:cN���0 �W�
�&E#x��$�<T1(��2��g.8�m�cT�j��[w����y�۝D�ú5��O��l��2wG�D�vWM!r��A���w��`��S��$�W`9Z�{^�%ñ�C�~;�ڎ�'(>������g3�}�o�R�0䗡_C\&Lޭ�Z�.�q%�o^i����=���A����wJ���c��cA��i�6��R�(I�Ty�z����r`�T�);��sίm��o���U�ڰ̩���[k}��G.-˓��tvrP�պ����Ņ��+A�&�KU��kx:�+��F1�Շ{V�7���8u���]�V]�on�@�'ZBM#Q������'��E�8�s��f<.ڰֳ�qr�|�Tqӥ���}ǚ��^��A4����P�_^�ӻ�֒�L��r)u�:\]�^YR���#��w#�(Ρ�r��gV2�;�#�{��8e��7���
�<��s�� �u�|��׌�-��z1R�����a��T�;�pN�<v⇦ф�B�u����c�q�i#�u�˶�ыM��Ţ��܀{X�boZ'�ifϏL�ɇ�0�0��jv���r���]{����@[�T���cK��b�-ywwI�\��ip�� �-�'��o��,�*���t�vn-�~2>��m��Fz�6*�	�*�:�3��xc��٧��S��p�6"oUy�=��������Y.Wr��G7;�V�ѭ]�M/2�:{,(�i���8�ӎ�Ň-�WY�$8&%x/L� ����v�*���nC���wv��B���6���̹'8�~��ݭM
��v)��yKX�p9/dc Z��^���	�z!�mz�:�ɍ����Y�ȷFu]��֤cv�],�٬n�<rJ��J�\`����H/�ն����ϵ���Μ�U�R�:L8�t22����7�Z������t!�p���^ch�ؕ4��V������wY-΁�d�7rvl�L��Y^ Ǧu��lS�]�u\��޹:�R5�ӃCWq���Pё��RQur�{��6�eZ�Aι�q�P�EA��YX��#�=��L9c�+oct��>\�Nf�㽤�ˬUJ1�Ka)&#9b�BO�2�X$�i�Ӟ��1�K%�"��5��Y�dd{f�#�xZR�6d3\�sb}&�*�7w9b�<]V�sǦf�㋻t���-��a�qnk�:Y�Ik���e8���>�^�w�3�ӡX4��[���1�ZV�������l=�9�3z]g6�/bJacN]גn> ͊��i�A� �)���]m�N��ǂ �S��V���R�ف���p��i?T��\.d9�QL��w4�YW�m�h��A��������P"���%��qn��v��\���i���t�{.��nj��[+FU��4*� r��<zj&���1ø-�t�Xc�'[�~sn0_q���q�ҸRQ`TY�Y-������8��ɔ�&��#NT3��Ω�[����܇���PbX�l �xrǧ1���eoo\6_�΅��h�E80�B��T���������Z��\�s��[#q8�2{�;�7�-�1�����&Q	���٦�*�hx#�SŢ��^�7�R�1�i[�&�.��:F{��)�u��{�:'43�7�h�a�&��"�ع���m
8��4P-�l��t�\;�Ro{u�@�k'��B��/Ju�叵iJ@�Ջ��[k���,
�x-|�rE�h��]Ӹ!���=�j�J�Pj��jz�d���S[�-�ro7�kڞAF���R6�;��Q����y�����3�qm�&Gx@[��C�����ξK�,�F���BQ�-RUt�3��P��#���tU�lW1�e3F'+�<����K���{.�:�ef]��ɷ+����1�5�ol�e�s�
�S�gl8�+��Q`M�B��d�Orga0vB\�5IA0��{�n��"uT'0�;j<;l,j��)TѤpR\���Fpj���O��U=Z��{$��$�`,'x׳��3�{T]=��[ݓ;�;1��0=�ӧ�k84h$��4����cY�GmW6�C-Џ. ¨�1�J�r*�NL�PR�<ZZ_�\�u��6Z�>��/��X��/�� r�	�bH%��>���P/o
�A���\�6�e�����r;��K�Wl�M��$�/k���/ ��NLQ�vQ�9"������g� ��%+˪G_'_��!+��4`����G�"����	��Fݸ�D�nn�ݹ���Ss��� -ɗ@(��z��nGT�K��Pt�x�$�ĵ`�n��s���Q��ڷTӖ&Vj�ܮ��"�fѸ#դ3���wB���sNs�����,�9e4ժK��d�����-��#�����N��^�'pGp����\�	��ŗ�cs�����/6�Ζs6�7l���5&`:#'F��y3t�QU���g
~i�ƾ��;L��8���C��I�Q��ܣU�u�UD��Їcޜ�su�"i:���h�����7{�E���<���}����ɤN�V��L��	_>�sA]S�W�a�<J԰4�������ʻ�6��ǌȃ�n�rj�9�cf"��w�('ʊv���F���y�qqwz����R;�q��XQ��r�fG�M�6�� 6��.�{)9�w�o)3�(Y8���:��|	ps��^�������Έ�Ж(�}�-��$�wf�SZ=/��jb3b06����c��Nr�>��J�O��P�f:��2��]�v��:�F=89d˼�r��J�5)] �;����%�n��x�p
s���:٬=+f%�7�t���I ����*$�Go[���]�H��$��	�*C�i��׽0�a�ǵm��J�
A�^{9r�ؓz��MC8��si��㝏��j���F�Q���h�q�Jp$��i�H?)�/�+pb[�z�mÛ���&�h�Y���Y���e�^��8� sM��ͱx��v�����]�goa�NS�Ү<�x�8uZ��5-$U�]��x���%9�7���MJ1m ���TZzQz&9c��t��A����h��VεBX�u�s��0 3^p�T�rcnv�U�[�a��$�A��"+y��h��=[ȾCUA�>��"��:
dG hv!����]w��Y81�z��o-�X�\t��m��`�۬^ޏ+Ciʵ�m�C7m:5��	D�m��t�Z�����7��0έrūtpk�ֶ����-�t�SO�U����ya�@��,�mj:�r�m5�G}��5����zt���(Q���b2<v�����8�:A�9�ˌ˼����1�G��R����)wƃʺ�-�{qdB�����ݍ�9A]MH+`�Ҭ����9�"�S]Q	ǎNǩJ���;D�6�|��ʸ�l��6;;�Jgwu�
��G[y����8��PY2�˶ϒ�J��{F6��{&ղ�#������#�7I��˜D��[ۉQ��gK���}٠���{LpL�,����,D��QxVh�v���-���l�e�0�ڷ$��q���OwqI�`c��ځ�	.j�2D��ݐ.�&80�>U�l.��wn�
�׍���4�&��p/���L)�mY����׳L���O�`)cͧh˶�w�owi��Nd��+w��#�ˑ��r��Q�cQ[y�GU)v>;-�����C�۽Ò�_^�8N��t�����Õbeˬt��F���$�.L�8�;.��j<iך,���ܗ'Ut`��2i&���C�:E�\#�r�G%�)���Ҁ����udUĤF͇4�t�N�Q�P��I�j/���{�sgf�:w�0=�W��7�{k��t�\ܙ�1^��,:��t��s4W�X���@zӺ�3`FB�j��;ũ���+.����/��zw)��֧n-��]cx��]��
�.6�)����8�8�K"°]=1
�&�
�S�:t�v�Fov in�s��tF�s��3w@8��C���]ꪰqGq2&h�δ���������@ �N
9��m���G
ٻ�wi����y�>A`ɇo��l����0�a�d�	���ù�NN�4N%7�`<_;,}�g]3$�.�j���E�nhۛp�7窽���s�������T��z���>ӓ�\C�L(�i��ۊ]�6�1�Q�U� [��;�rqn84f�0>�FԵ�4�G+��� ��Vq��Z�ޛ�ӌr� kN6]�\�6C�Z����z�I$P������$	"�$�,� �� @�XH�a	!u]Eu��UQU�UtU�d$"�
��!,	 P,��@ �)	!���H)	"�BE��$�B
HE�R�	�()"�H)A��,Ad�
� ��X��$ @HBE$I	�!"�B
HE X�B
A@�)!$R�I!	�@�BE		$Y	 �$��I I$RE$�I@�	,$�BH�R,��Y�	H )$������H�)$�,�E ,	'��$�HH~@!I>��R�DO߿?i*�V�
�J�z(7�ng$�<u3^��ĝڙd�n�ڔ��w��Gj��C�Z�X���h�'�Pxw-[���h�0l������s=�mwvdEu�BԽ��y�o�����Ҙ�@���r�g^��S|h��W�sRWxZ�u)}q�N_y���Q��-�j�DR.��+>z[�Т�L>�E�����,�5��v�� �BC�TwCܣ�n���C�ݓ������'t��yN_z�v�]��I4�1T��\�з5[�qk�A�����'K����M�;���e�ǽ&.���7���$��׍��F�{J�������u�wn�}Q�	��.��W���Ϲ-)=�y�~��c�y��$n*H�%J��ʳ��£�i7ئ�-��ꠔ|��$s�;ҝ����F]��wG35Ԍ�$-�ͅ����Ie�1Fu+P�TR%ֹs��ˣw~l�c��s��r�����n��ӓ��u��uJT\P����\�kFR��fx��u��H�|��Ӈ��%��&�-g��A�5rx�O/w��@��n�)co,�x��g����&2�&5��c%�ʐ�sP_f�ķ��^���6=#����:���q�z�'�u_[��ph�Cnr����ГL�`�n�
HޞI	6`�.Pge������|�e��>����{��X{���{��Eƭ��,��c��e-b��ݕb�qE���Fd��A��֊i�\{�@N�O�O���5K�[;6L�Nn��o"U��O`So�FO�A�]d[MԨ,�/'��#�u��s�r�����S;�p�QD�#p�ԍ���t�}�jE�{�o[��q*=3j�j'T(�����6D98��sZ�fnJ͟mʹ��NQ�Q2&�.�M�5��z��͡����A����q�^�7�,���KW�kv�X�2��:*����4�6��L�O*�2=�v��D���D�
tE�����+,Uڷ�������];6���7�������t������{�3�T�e��q+�*>���	=����#�� �Ŏ���Y"O�����j�
���M���>�-^Y��b�Oxx%8����۱�ޓG;�:�.�Ԍ��o@��n�#T`�טp�j�@ |�q���7p�2�ﯙ>��*7ۤ�F���y�W0�^op�{tL:;m��w�����w�����99�1�O,���Ί��ɧz���������8�nk�_tԅ�1�0��ݚt��v�{�O��S��O�yщ6��μ�{����yNA�+Ffa��������F7�S��K��t�5�F�%��[�ɬ%�D�r�^kIw~��Z&��E��� ED{��뚷=��R޺o�����WNyy���0�J�ʽ�i\8e�u��B�vL��MC3]ޝ��w��CtO{��q^���}s��v�|;���z���
�ƂZ��ӎE�c���e�o���
�P�g���Y�(��������8=���Y�1��]��S�����.l�v�Y�d�9Y�wr�')#Le��B	��y!�l��s�&��u��m7��w��FU�&�T8�{�ݺ�n�Uq�w��y�#��#s{�A��^�E�U0�u|�ɋ޵�Z�~��ԗz�ޫ��&n��6�sP:(k"�:
DX5��^��1N��Y�J����{���&�pb�,��q��uǢL���F��DbXs��6gg��4��Ӟ����E�:gz��{cV� Ae��r~���n��lNt��/A,�����{g���!�}/���^z<<��dx�i�E�r^�)0%۝��Pdנ��ˁ5[R(-�Q��A��h(���Q�hUS��q�fg�6^kG*�aD���2[5�Ys��ޮg�P��s��.7��B9��]϶���R�)�<)�C*׹p�z�|��\�V<�;��K�z<"t"߭G�e	��)�/�s�*�ٹ�}�<3��s��{
�3�Xc�a�F;����NⅨ�T���e�n�.c��ǩ����LOO{{ik��u�W�{�T�"�؂��sv�e���h*�ur�5'��L���4_�}���#]���mO`~~<��]sZzpc'��1ʘ�	�G���]{[ɪ�O;
<�oh6��Ĳ�э�)�lޒ�<�=�KI�g6�ܑ�TT�b'��y�tݬ!�v34�(v�@��W��0��i�����{g^t_Y5k�rH3��V�T��P�y�|�xE�æK�!<��]����jo�œ���g-�����S_*�b_ ��]�o����̡��<���G{~���z��p+����z^X}�҂�UZ�-�j\݊۝��T�-\E�F�{��!L6�ɚ�+�}�f�>�v=ù�1!������*��2��t^N�lN�;�.�.eْ�A~վ�0������}��8��Q�����[sУ��η���h��h:,��P!�d���݇Ӯ�o���w�Şk�ۤ�q?������f�k�����B���꽆�Ht���wf8�}�=p&���r�ܦ����G��5�*0=��x3Nw���>#��2�w����
�G�d�./��
�S�&� �:��Z.���Χ��/vp`^���j$�ݾ�|qq�(w<'��t����s�9eYl���������O��_rn`�3¸��}�6v��懚[z��'0�����W��nLj1s}N��!+�|���0��A�6t@�ۺ����vp��ʽ{�0H�ȚS�6���Q�={���ҋ>�2�˧�6`����}|��7�T{Hn�����}��^Z5����HDr�Z��C�th:�?u��U���Bg �g�C'z��������|R�5Ou�^�9���8��e��m���~���v�b������D�CE{G_4�biɳ���:�隆ŎQ�(���Qo�`�����ˇW�	�6����A��ə��[µ�{]��宸zJv��
&b5�5�n��e{��Ə�`>tL��H\��V��ua�����D)CRf�E��L�%�W �*�j'���������N��[�<��t���f�V�`�z��
B݇O^էiݾ����קv+�˝�]Ji�^��[��w��V��8�����{�u����FXx]�0���3Do���6	��Pܫ7|gME������z���+�ж~NOI]V��_!����|��j,���{�}͕�s����ͻ��,��ɜ��X�'am[���3��rf
'S&��[yP>�(6�/gw,٪�o�}�w�.~�Ӭ9s{�uU87}�Kv � ���<}=��N��b��߹�nU�\�X4,.�t�uꋴ�k1"�8���W�\��eQNh�8
i�]��ם<pSW�ڳ+M��.�Ý.��<���)&/��K RY�Ԛ�mg�{�����N;ny�6Z���4��I%i;+@��b@&�w%�2C���]��Ŗw��4s"�Ev��kl{��'ݲ�;H'� ��P�{(9���み�k?Q�ڶ����]ך���(��H��Z��޸7���v��z��x��^���]*H]���q�E˲���]��1<��Ru��rv�.V�� ӓ���!b���v�}90D��MPI�t�Te���O���E�'���<D��+��])���f�I�ó}�}�.��N�S�"���Wf�$���o����3G�cԅL=��Y}��oڇVfl�:�W��~�;E�5gm��ճ���b�c*�[�.H�4C�n��]S2����)���⃗H��j�Y���=���2U�R�;��X�eS��JPsKM�b���;%���e	�9���yw"���OK���:u@��	{w�2M]��qU����v�B�{پy�'7�֯�D�Wp{<n�kn���_��}��"U��{3Nk�ɋ7��Y>��N��%�\�o���<����!e�J��ri;��="ܖŖ��v��W�4�^�����0�#=�����Y�!��$Y��	�;��q�=��_a��A`��c��ti� q<��`�|J��n�%������/7��ܧ�����U�(�Y��f��yn9��B��3�{���]��=:Lc�ܼWcx'�/���}��nϣ�X��F�Y��k������2��qltMb5_'��No��#U�-E��
��������VU��U����ݝ����s=�N��l�ǁӨ�`飷"���]R��ԁ'�������k�*�σ䳟�5�HvNn�v��¹�8�O�X�C`Q���]���������0o������<���|]O���3o*��wx���:�C#W*6X��Zs~I�qe[�c!��,;���c��_vB>A��<|� ��ȴ�H�-�̷����p1�=G-��̩t͝�C�@�~�� \�~�Q���>y��ky�q+&k�
"���"�2�����`j_��Fn)�
��'QX�,��n�1��>����7pf��ڶ
4ԥ3��9�с��}���[-�S���L���ٵ�/L����sv䣾~w�5���o�b�n�T���|{��:�Tb���>9`����$�q]�/g9�6v���N�����}[�˯OG�#�夁޽��R=@�Bo�~)�^~+O���-�x�z\|���p�^�l{+�.e��d֕��z&��N���X')��v�ʣE<е1nK��4])��5�Ki)r�cef�)a6S�<;Au�P�ײ9Gn�ci�2R�x��"gOWb<���i;��7�,x��������{ �:�c��G{ؼ�^z�>��L�B�!Z
/y�ǻޘ0=�#����c�v�V���G�՞�hͣ{�ܮ��u�m����/�om��fa��6���0d�JaiB"����}T�}�ET�C�F��8��)Y
�5�ձUP�3s�jh�!ˉk���=}��KD�j=W�1�V��u�|\���t�n�Jy�BNh�_Y<0%��9㋅�Y�z��ܔ�;�Q.�`{-���f�3�:��7=���S3}�=���^ޠ��\���"�jQ�:�ͷu��5q�����x�þ�8vW��x����ګ�
��1گ���Wu�%ؼ�xi������Ğ5d�ɯz�
�������a�<0wn͹"�D�(a��D�1a�:+����t�Z<��<��W��
ƃ0��ᱟPOYz�:�����z�m����l��Ǖ,�osԙӺ°mԴJ�l�� ��K�v[����i[V����mi.��)�zm`�;`�.����2V����= ��fQ���{ˆv;˞-�k�{]".;�,ד.��tLv[��,S��s�B�&�ny`��o�{�E����s�d�Ɔ�`�Ai��4��ب� �V��5i�k���G�(H��9�.��>��8��
�$ݑ#w\����.l��M�3#�ok���{�t�n�n�uG�I�4��Dȹ��x��]�Kw����W�����+b�i��9b�xz�IW{a]�`�₩��B�j�4�����%빸���&y��˜�)qX��>�}�w�\};P���Ӏ`ɺWW��OHWH��!ܘsXc1�+q��^>�r;���q�����Q�C=(�߇;�|�xa�9vnv����p�I���X&C�Eo�7����3�}�%���4?[ʙ���^s�y`a�s�GY�y��~V�"	�s�B�+Q���f6`�vT�A�q�Z�w@��l4�`f��97bo]�7A���~����qp6�x�]>�x����m[&�6��&��& �*	��X��x�<M�ɒ����)G�R�&cd2��p5;�87��s&����jxϽ<���F�l$�B~,XB�tM8n˛��*Uҥ]n���g�k�sL^8Pk�bHwQ���P:X��7��a��O�6�v� ��X��K��X���0�[G��rۆ5��
���'E��E�8̍j�}��L*w�n�0����91�	�f��˽��L���Ǧ)�vy�})�ф{�$F9f����g}��@��Rɂ�*�tT�O^U��:7�z�\,����߯���~~=�L S����Uܕ���4V�O���ٝ
����a��\靷��^��a�=k��ݰ�՛>�7[sn
����ͽzq�,=���Vz�x	�M�l�|ɲ:�[�C㰠� =��g"�m���Z�.DIcј�L
RmDP�ȕo�U�R�b�WY�0|�.�w�^��AO���'�[���[S��t����Z�-�z�v�⣏�|Sf#7�K�y{�{A4R4�,ن�THP빷�F�$�M�q+n��/^A�56�ҥ��dY0��ϛ�4-���A7��i����7!�j�-]^��Ʒ�Þ(�_�1�R �P��_w�rAS��t)E���I�)�Υ��^OdD��j�GwZ=�'�Rx����1Oh��2)y�<Ō��-��A�]˙�n9�c*�<)�a+�;�oz�R��w4z�Pu���)"����� Z�,�x��۾p��/p�W��Oi��z#ܸ~x}i�;�ͣ0�e)���c��[�Sm!���ك�yO��@Ӣ����КdR"5g�?�^ɽn�M��D~|��i�M/'-�
���]!�{�ܜw���h�Yʥ�FzW����׈��4����rU�v�3�-�m�o�I�A�!tEY���=�jW����>�%��5 _>J0n���-�@V�ޘ8]haA��ܲ{ٰ�[pp�>�S=��A�i�RsK��
/��S=��9i[rns�-z}�777}�~[�B�4�g2��:��3�iP�+��n�X$��ص��R�ءO|qyK���Q�Ƈ˸�,����׆T�9����Fo�v�>4�����o�u��������� �p�^�탐J᥅Ζ��3,)�mf�1x�G[f"[6�q����l�A��3ci*.�%廖f*S�j�\�5��E�@ٚ�!�\�.3
��x�w��sٵ-���v�G1IYf1)	@�v�XÛIf�A�����ZTjK�:#���6���Ř�L��ic��D3�7h�ᚳ��Y������Q���˫�7 U�]�8���O!-m�1���M4��R)�R���i�Τ%�\�A�h�cZ3`�^@�L'e�P�Y�jX]��M�f:#�i��Bc�l15�F�)i���ں(R��S;@�1�5�3,�c,�瓂k]E�ɰ�FYW��\ó���lB�;��훮v3��RUT�!1�%�,\=YK�օ&�7.��5����!NMM���5���oYu�m�hК�Db� �梤J�%2�6�t����i��VY�ɉ�����BWv�YKx����a:�hL���4�0JY)-��v�[���(��g�U6�on��R=��Mc��-M��tة0te�ŕd�Q#&ګ�6Z���mK�-6j�!�ظe��z��1e,P+n��T�R�L���xy.֣4�+�f�֚����)���Y�(�Gmf�Vm�KE���d���t5�A�-!Ee`�\�KP�&�)�j�Տ��	k��ai.��0��.��բ@�n�J�n�����r�y@�A�K����V�Ջ�(��l���Щ�˄�iZklRز�5+���ha�B�AҌP�ir�6���*�3B	�S1%wY��4�uM�%���]�at��4CK�R.ճBj�4es��[���YV5sF1�h�k�	f4��N�Mz��a)i3)��f6��1����5�:ƙJݜl.3GGD��C��3h��9�#ZjEDz�=DJ�����	R[[-�
T��sa]1�e,r9�#n�XV(��v�g@tl���Թ�@�Y���e�C�$	�۠�i����#Fb�ĶU�y�����&��à�R�X�!�A�"�ki�����:�0���[�v�g��V�m^�����a��-څ]��sK3c�7��d���]ˆ���]\D�6�ŎdK��e��U�8�v�iA�ȝ�mH�>�i䶁�N�R�Y��)hC*Wd��V��P�7P��X�:��&���X�'�x��.�Y��)�`�U����x�9c\�[�]P��l�]4�E[WM���mv�cV�l��7Z���j�RhmQ� ��-���O�*x6ǋ�n�ZJІ���I�0#-�5H����L�jL�ۻ�*��F�i�tk�
�X�q-i�e���4 =J����� �EN���BK�MD������`ie�\sf��1 ����
c,2R�x��̬�Uf���Xv�ՕnBݜ.���iR����@��'�:5i*�f�R�M�fK�C
�17Lꔙ�`T��m���TWd��ݰh�lm�
hݥ��tԭ�l�tEMAE���7bԴ�H��X�E44�&��gY�f&3LBX��mk���X����P�W��f�fҤy��5L�k\�+I��� #ar��r�0��ݴ��P��n�Z�e0]�Yh���pKP�;ljæ d�#5|��!��H��=�cVb��y��֧ik�[2�k�ԘX�5��5���%�[��4	M�[b�$��[�6%ڳ��cfu�b�i5W�0T��c"�f�1�p�k*�mv��4C1LY�g6�i�@��,���J�͌Ԧ��CZ��J�1MC��͎i��R�Iu���P&����E�Gͷ�0Y�L[5�`v�%1� Zܲ!P՗Jl�����!b�H6�n�9ܚ�ܸm�Uѣ����	���:2�eq&ڤMam+1�q1��;V��GCki+�0K
�ѹf���6�I�ģ�)
��+�U��k3y�x5�J8#ef1�� J��B���J������:��1��,�5k�EGl��E,�.�HYn�"e�:3BҚ��Q�����֙��%��Xa��xNc�#Bh����͙���j��JH���)i�o:Q
��@��z�a�R����a������*�]E��͙���\u�������f�Iu[q;WV�ʫSb�[��k:��0�6�Yj�3V�r6Lĭ�W�VV�M����0�=��
割�&53 ��n�`�e��XBa�l[B��-0Ct�ұ�M+�m��)�٫�����Ktu�j!)pP�5wQs�ѳ�(�u��ii��� 15���`��(�
�a�V+n%��^��X���Z��P�G2�]�Bm��R�[�X,53\�Z])�5bU�ڄ��S6X5��� ���A�scp��"c���T��u��B5�-�Х�[U5�,�c\�Su�]H�Kq���Ck��2�1.�c\ Vӑֶ6bZ\KP&��69��M�T�L\AK	��ic�������aCm2�(݅5rkK)�/Ut���݄)�누A�14҈��ɲ�T�"�v&�3Q��b���pW��4ғ]��i�n2cB�U���v�aanu�Z�h�KK���We�u+���I	@�m��ô�3YUٺ�Z馘�8�9�e��&se�4��̄f���cY��5�kE�Fmxt�d4���4��Y]A�(3X�G+c��.N	s5��a��a�f����I[mIQ`�b�j�1ih��v	q,9pj���\���6�1��蕛@��z�Ĕeͭ��F�v�A�6r�&��7]6lC퀦��i-XMk�J��G;X�]0 <pMu�Wa�;�UYt�hY�+��u�����]*	,fe��]�6�������9��m���3�[Km]��l��-�35�|���������I[2��e�lX��.��x�B`<�:�Dl�hRB]�K�fT�MK��-7easm��
�S!IqK,qr�le��31���^�+e!et�h��R���G��j6�ѱp F͡Y[�;f$k�Ѷ��̀�%cE�����/�M� �{[����*��D��3��b�K�3xea�ּ�(D�]7c-y��2�:�)���@��z�1�k��F�JP�4R��F������)iB����s��0ķ�L_"���Me�j5Y�(���77-&��6�lU�*`ekKfm�6[E���ҹ��.��A(�㘚�β�ѬıQm֩\��m�a���6�H�`��h	-3ɣ���D3\0]Ʃ3MD��P^9��.�l<먻V��B[V�5�������V:��%���T���u2m�!�L[��j��%CZ@,\X���.%/�U��������V]G@�ܾV��� �6�<ʖ۲vbj��X��M�����A�45��.����%V-���aj͔SQ2M^�\����ť��ԅ,�lBR^�l��MfB�5�Nf6�;hL5&\�Sk�Rm�BR�+� [��mAbC���|q�151rM��
��ԚYbY������u� ���a�����W�]���VxCkA�hT��"35�2�(�eH؀ͬ�[�If��f�5е��ݮ �2	�R'm"�
it ���lh��SXpZ��Ń@�T�ᆚ̠◃L�R��TL.���'��7�4�,#l!�]lƥ�2���5!�y��(i��bR1V�ͭ���j��H��cj��Υr�Z�b��Bf2�V�vX [�r����l�0[E�m��r��v�r�JL1f�5�.�a��7a���]x!��a���,�-����5d,��b��6�r��L�6X��6�ɦ�Ք�l:E+�6c�re[�f0lH���e�h��Z�2͂�:YMU��J�K�藙�e4B�ax��v��
z�����8MneX���,	��]�n�j6R�	���̧]��԰[��D�\�6��
�]o+B��e�f�cc"%��GR0���Mm��%��S��
�i�-Uh�]�K�C�|�O+f�i<l&����6��1���iH]�P��j�ۈT*�ճp���S�"ɵ\��YWm������b7	gf�wU9�I��m��R�)k�дe4 �8alYe�ǋfR`�͍6�d��3m�j�p�:l�ٸlP���L�q��:Z �Fe�M�uM��G�V˖^��f�4B5�3�YX�k���ʭ۰�m�Y�:褥�K��#��)n]ڵ� �aK��J��	��12J5�lwf�%n2�u2Zk���5��ф��L�p5�iks�HV�l�	9���F�av͔�i�Ҏt\Lc��8�s2�m��k6iK0��UM��3㵞2x�q��ڹT �.��A �L�n���ݫ �,��7W$��\���B�b���׮��ƫ�^��h:0��mbZK 	�ʺ,6��Ik�J�5@�͌6Ȍɫb�R��i��z�`�1����b�؅	� 5ەշR�l	�V�.4�&b�gU5�(�A��:�V��kM���i �6�^��&��t�nB[K	e����bM+�X���������t�F�g:�بR�0K"���$ۑ��H�1��Yt�2���9�Zɇk�=@q�8��Mf��eM]��%l+CE��EٗmbJ׭���v�e3J찜2�<��hD�kwV��2L(\�,��BJ�\D+P⸎5��])�&��2���n�k�����(51M4�e�@�tY�1�u7h�f]iq�TqW�^̾XW��d�`�ЈA!�e3)Z͂�s0�e��@��R�q]ai�"����b4,�vb�9��Ws���nkSB��3�i�eɲ��j��:ƒ��kòmX�D7[& ݢC6�'k�$�*2�5���h�YZ�)l�0��G�cbZ0 �̺�&s+�L��i��&�,0sZX+c�u��]���4c�\�g]�\�UUUUT+�u�UUUL��
��UUUU�Q�&��W��F[�l�j�W*����8�!���y��s���	�'����!D-mV���lJ'����)-�q���Q���"Bn]�Q�!(� �-��e{���������6�t��GY{c����Vs�K�DPAY�'8��;�����l�8��8q��N;.m�Bp\�I"\VV	�؇{]�n�	�+�Y�	��� ]98S����E=�H��ي���μ��X��X�0�����*��Q$�=��2}����9]���{5�iA�i~ol��':m�W�Ȝw� ��|�kSL�����n�&_mÀQۯm�-��_[|�:$�����y�r:Rq#k$8��.�H��$N������+΍����)�;>gu���+J�}��+��֧�{�$����ґ�,��
�Y��!6�K8�K�L�9m�D�����i���3.-n�+�֤dnJn�8-��p �H]..����j��jB�S@�LA��Z ܶ�eFWgB�M�܄b2��]����e�XB*�u��Y]�-j2�D�16��0cB:l6�g�h���0���er7��%ځ0s� ��9�f�a�[R�L�Fn�֙��qf���aA3��Ʌ!D3��l�Yt�nB��)0�]�k��� ci�Wie�&�u+c6��WP��JG%nt����q�L���Zh�(�!�N3g��Š(��[V�tcuqRfk���ʱ�<��W�B��3d ��	�B�:\s,36�W�b�*�,���@f)1��5�Ƃ�ũ�2F���IA�Xњ��,�h0����,&%p��ɢ�FYb��Y�(]�dʐv c3`Yu5r�(�te�F洲d�BK���r�ؖW&n�4�5n�#a-����v��v���1	�3+��IRPa�4u2Ki�,�2B�K����)�^c5��4�v��GXk���<7Ű�� Me/l�#�c`�2m.5�:EN��cU�.3vV����M�S�8:�!2dvZ�ͰXк�khڔ��"s2M��Q�u*\��"6���%;Y�%���.!X�9ѹll�2D�
[�hn�a:�WqM��7��%��+���.-�5�.�$�W[rQ�%��0E��Cf�.R���JP��9ys���4�Ȑ�Ē񝫨E�ʹء�%f��j\�U!q�%KinQM:t6�]��&r���#�m+2�@�K�ѥ�L������a�PB��YdkT�CJ�lXa�������Z���b�tH��7%cuu�5ib�6�+[�)�U�B\D�h��m`���0v�BmJ	.k6��3X�#���nYh�4Mz��k�F�\R�(a�[\Vf�s�KT6ʶ�����W��F�@	i��<�lP�+-�%�j*�a[<Z���a(5m��2fy�o^�7kw��$�ޒ���-j*Ք��*���6V�TEl��m�V��6��1�J�i��%��-H�o0�y�+-(�^m���R�4�ZI[�e1 ����2Tk.�JL�ʱ�,�e����} BG�9�8�u���(�mKJ�qS-a��-"�4C4�-��o��H|��IJ=v'�ݡGQ���1.,E��Y�~��8V��AIЯ�⒡E%4A&
L�M�t�t��3�M2#V�����3[��W�l�J=%=cemN�2OM͑�q�J� ���� ���Un�]��kw�]k��DU�!���.�E%4$#䕊��et���N�+�ȏ�4 $�R�靖�p����Z�"��G�&݇y]���`v��Jt�QT(����oo-����"�nC�}�M���s�ֶEx� �� ��ٷ����'��~l͸��qq9�����E.���wi��B�aX�D�1����ϛ���� �`$�b�꺵cu8�`�s�����#�bg�)l�+T�� $���JE24nT�d����'���m�Fa;S��g�Q�ī�w\��'Q��{�h�K�{;+�`����1��T�Wjۊ�i�U^�6� �>����Jj�;��7�x��S�z�]��ٓ��~[*��Ӡ��U��
")ب�����q�]�q�b�rÜ�P&�ȠB>���$�h!Fʆr����Ҁ �t(�0�J�b���)�˚������@#P�DMOPϨD��(��AG��%=nq<����AB�����]�k�����W���<��}���T���331>Z�G��1��v���H&J�lcS:���2�C	�2g2�H � �u��>DFZ�}+'�!جL�Xy\��HGrfRy�,���6AIP��A))�.�bٸ��y���3/j:u52�g;��DF�@��(9�X����4Dx�}@P ��A
= ���AIP�R����e�D�\|�.�������b�cN����7�
=�{(�r5�v�ɪ[�vo�K��Cڵ�+׻MI�\j�m�qp��^'�Y4/U
!R,���/3���E� ��(Q�s@�
"�뎛���v&7,9ΠA��(��7�y�={���՝�(�����T(�pM3��{�Kc����O`���e��؇s�8D A��x��� ���2�Kl�D���&"���L��Qt����!�%����)�$�.��D�]P���2y
�9A�AIO�R4(��4�>�m�mx�>�F���Z]N����_���J���x� �o�琞Li���(���7� ��a�u�"�!G�����UJ����+C�^P�4� ��RJ��⒡j�,D��U�B|�L���x�]B�IMxJ"	*+�ܦ�f��wr`�6)*�c��t���k�� ��4��:������`���;3�eg�(��n1ǸNtx�5sT�C*#7"DB�P�&khW�H'}:F��n�'��gMv�B�q`v�
Jk�QIH�����q֨lO���6T\7�G:'rÜ�@�J@G�
JhRT-���Yv�:31&bd/j�Ѥf%�b��b�%��LxT�Ys�W1(Wb[.�t�<����L��hN���{�^}�`b9>*e��؅s���D;�ʋȐ��Zs^ �Q%b�%"�]Uw�q���fJ;z�;n�7j86c�^'�>7j}A��y����f�ţ��1e
)����
%>�D:!�;�����wi0�,F�9#�� W�>IM�|��@(�t��<t�K��!�W��)*3�O&9L0��}�a�*��y|��l_�{4A!$�
�JEADG�Jo�;�܅�����
���T�����
��= ��4!�D#��*6(����lfs9��ť�<z;t�m�g���6G/߫L���;hƄw@�vБ��A3���/w085��:���M�ʑ9��o�wBR�kM�&#��6�uff6�IuK��.�ʱh¤̺�b
źVQIGs�j��GbT����*�!�B�1XYv�iZ�ۊYr�;�*�p��#c�0Y�.�;9Ѷd
�,�P���F��Û5�h�, m�t��F��e��RR.-�\f�t\�+֎�d
K�Ŷ��sp��a2�SZX6����'�v|���@�4a���`��jC4̙1.�e3km�i��U_u��I����ADF�zc���&E�ܰ�;�6�b�S��R{��S��y%B�G�
Jhѓ��%�24���B�4��3��*�#b�8D@��(����3b��̑&H��^MȢ
�Sd�	U�t�|gn傩[�f2�jE�F7�ބC9�4�i���F���������h� �*
JhAD@P�޺���L�I��!gW�l� ���;���s^#5H����%B��;54�Q�K�JC����9�r]�b�| ����� �E�<��2.�x���0�����lM�qj�&�������k6��j�T
f���o��~�a�����R)E�*��/�����A<B���L#�py:�>>IP��� �� ����q����̐�Œ�nٛm�'�U9�pL���sbٗ���{����<��D�P*k`o;?\��M�Es��u:8�sD�#��J���MS�+0B���� ��
Jn/m��`�{��P�E�Ϧ�!%B�� $�E��Ww�����GC�]NK�lF����5�(���D��Ϥ9�Yl�uE�rd����*
��ӫl�r�5H'��Қ�jIWz{g���0�f�]B�IM |��BJ�x���r�p���T��ip��L�8প8J�����D��⒚���K���d��`9$a��]�tf���(ց�a4E��9m�!*@ݦ�kU�N��}�A��]�'{����銖��ї�b2�C;�n.i�dLǷ��M�+ϕ{u���∂S䔍 �Q�޺2����]4>ԨP)�ri�}�^ O	�S^ �t(�:��|d��F�У��G�D
J���Q��ţ�6�WpW=��[P�rW">Lt�!x�s���7ő�5s%��QKčnm�k�{��Z�u	��'-��f2�'�YN^�eD�p�fܣTgS-LUK�,�P �����@))�A�J����jd�[�#2�nYg:F<|BJ�d��t跹��a�،���`Y���1�:�� �@I]RR(Tz<RS��`u��Bˁљ^x;&)S��`�^ Ox�Қ���䔅��-ӭ�(I�U&*�Ma��ya�2�jԗ:Q��hh�Z�ˇn%S	�5�Rɔ�w����
))�|�����gy�S�Q*�)�2�s�fҐ(��j�$�h!�)����R2+�Lt��t27x˝Eod��wtc.x��E�RS6Z/E�A�U��"��k�^ �� RSDJ�J's�t�����b��.�99{
�<A3[5���P#�$�P))�]ϻvTݾ�Q��B�J}E��Fw�r���T����fȯ��w\m�ۣ��5u�'������!R�Mڛ*�99w�n�4䷓j۞ܔ�p�X�j��"�Wt+��;|6�#u��2B�f$VV�g�A�4'Z��{��!��F�u�|ᾜ�9|P,���D�L��9��&�A8D99u)�":v�����p>Ԃ�]i�����E����L��ֲԅpm���!�`@��=?�ɥ��~f�^�I����)*���b��nT��,�", 낭��5��u�x��n�fψIP�����'�L8��y^Kx�{�Q��7��٪W���ml�!SuvvV�ў��]
# �⛚!%"�F<|���,�$u푏;�]�D�ũ�x]��e�N %�+�%4A$�����o^١t%�H�A�Ai�x���0�b��v��]�-��&�f�39Bɳ�oZF�ڔ�%4A ��
))��tཱ�����gW��5J�B��Z�A�AIM�Tq'��HBsQZ3�g=Ң�zcu��n���p���/��#Ǜy{��k�V�y�?��p�^7O��#1���{1R�$���͐dO�d�C�Gf�[����"kl�`!U���H��/8�[��Z(�Қ�U�x�*��;+\�����	��f��Ѽ��e�i�ok�Х[��Q�ֳ��3b`��a2�LZ�������rC��sڐ˦�Л,̣pLJ�/1��K�Z�����m+�4�i���B�5�k�4k\c]Q�����V-���N�3��z��}�vT�F3=�X��9��S75o�&�h�\���c����l���x����ޑ����u�=�ty^o�.usS�b�����8�l��"3hP=�k�Ȁ��W�R+�a�fw_S��F�y�˚ ��^L<��O��&���M^��#U�ٞ�͡GWMqAIP�RS@�Q�����z��h��5©^7>���z<RS^ ��
#C���P>��A{� ZJ����a�܌�<6��6�"�S�_CѲ�X�W)��"IU⒑D"Jj��
��4W�z�\cf��{�	��ՠ��Y5�Az�W�D	*I��r,�yP��>��TDS&[t6��Y�1�-�n��vHXl"3:$0$cvî)J � F�B�IMJ!Ǩ�s�fX�W����,�#L��L�a�9�
J�x�}))�:��u��٤������;���l\\,��5��.Sk�x;opw��;�-F�`���V�A�ĕj�+F
�w�E�;1u
�Ƣg[�F&�\9ʍ��}�@ ��W�S3w6�N���a��U�NEx�zIMRT+8\vN��Q�c(�KI�3f�h'�&o&����|��$�AS�>������B�w�k���磨�sf�R��*�W�l���ܫ��wF�^*�h
�B�! ��MRT(Y{/��!�����YB�^��+{�*f�\)ʍ��a#WP�⒚��b�՗Q�u�jf*Y�!�3�";GE�ΠW[5˯$�Y�iu���pa3ZV��URW��j{�l�!�({�ބRT(э�S��j�Z@�X�F��$��Z�;*rk�3:����$�H>(�"g��zv��=�h���ձ�������*����)G�����[���t(f�\�$�Q�>)*�"���Dl���a�(�Xn5�"XD�Նҩ��:���.F��S�K(�{�øa���<��5yQ}�q��ӓ�b�5Ҧt��%�� U��f�Ju���'o�55��1l��	8�y��5J�D��Rf�����u=���(j�(۽�W�"V{�bb��ڸ;.1ip%ԣw�n�n��<(�S�L��3%2�ɧ�4����fL�q�衾�숡�����m3C�I}�.9xȧ��x}�C8�s�U�9;����</3�H��&i�y��څC&j|H�:3��\�u�.�5�*�~�1@��Q�$�kW)�]�綨��7�Q�F���A�|Ǣ̀\~1��7y��b��3nu�B���1�tmDK
�v�����d�HK�N]W�MA��6`~}�7�f��y/P��R[����{:��N@{���vKٴ���U�����IB�>��
j��{w-ې�bˍ'�{Y7}}"��E�C����){˸����ڀ�
`Qs���y��ץ�}��}��
�=�f�ĸ�:`���]�:���V?#j�����Z,�s�Z:#����<��ѵD�{�P�y3����	�tt3���=�j��{h
�y�����r�����1�������"	�:̫�,S�\�6�=w�����v?Fr=�{!\<M��Su}�ڵ�e�y�Y��.G���>r9T�7E�{���z���1����'��� ӎn�[�/`��n<˨ � LӴ�9����������b�l�NYwl�3ˮo�|���tE*��"�
k�yՁ�a�.���׶����\'9 �[��IGY�yc��m��I�}����QEE���
'.�?}��r8�"': >vDSk�M��"EV��tS5�e坝�Di���ʹB�;��~ݢG_+.�۲��N��y�Gΰ���,������\ugwol��m������^^vyn]�����N��eyI�9s��.∣���)��V�����/;:���/0�:r��N:6�wu{�������Q[h�@�{wgI�wB����:�ʹ�wD�	���*�՜��.��[nʿ+���u�X[7$��$�	QW��q���l^�E��Q�Ԝ�j�Ä\vvfAͫI<�9�3��:N��ooq�A{n�Vp\� ����q�A����O.��\)���,�%d�'�@���^U@P�����$�)3,�M�) �P�r��iI�fXlv�Ro�wѳ9�=�,�A�!I��p��Xs=�i�FJH(P�fY���eg�U�^�Ͼ�׎��CUP���)����L��) �n�yҎ��u[�R��P.���h�g}�m �`RfY��@���\���bJH,*��m ��
@��4���zg5{���X�Y:2����]�8T���\�Gj�G�>�@�����3�i �RAk.�) ��ˆ���I
C3,�Aa����ӿz��镞�A|�v1�[1�1��x2�˚J��z�SM/SQ�,V�|��N��'�8����)�sۆ�62�
ϴm �6�Ar��R�̸m<	����~ˋYp�>�@�E���Y����~���<j����XPk��6�Xm� s��M�RAd��r��iI�fXn;H)
*���4�w(�$��ߚ�9������`):�L7��H)���X�<	�-};��]$����b �RAH,<�.d�) �Q�}Ѵ���Iʨ>����s/_kY��R��ۆ�� {ܳI�
H)����) ����6�Xn0�̳I7���L�*�(���:�oo��WVNܯ�Bf�j�G�>���AH}*��;f��!I�.�) ��ˆ��d�����i ��
H.U��$���5�~�G:����M��
��6�R
A}���TAH5P�ˆ��g��������o��v���/�Y��@���^U@P���X O>�.�_k(�W捞8�;p|�R�n�N�QNn��7�{+u���tC&%�ts,ڱx����i!+2fjZ5�Z��7�m�m]js����x,=aH��i&Ф��C)� \JH,32�c�����32�$�
H.0) ��p�&X�:"Z�{�z������O'
#]� ��F������!:��䔀h�F_TUŢk�]EDM �!2f�+��:�m����Ҭ����")��Ն�f��ΓHk,�}) ���N0) �>��Ci��RfY���Y7N0)�����_W+��^��ǩ���>6G�#×�En䯳k�Ȣ<(�$���R�)�}�ᤂ�P�C3,�Aa�0�����
J��p�&�RA@�7�_{��|~�H) �`{tAH,>Ϯ
#�����p��̅Ur�>�@�E$�ϣ%<`R��
3>�6�Xm� fe�I�w�迾�<H,�O�`��X}����U��f��!I���R�
a��3q��
fY��©��>%�w�2qR��*N��e�����L|0������.d�) �P{�Ѵ���H.0.肐Xw2ᤂ����i �o~�Q���W�w/�d�z��8	) ����Ci��R>��$��Y)���,�o��y��?Wwu��z�Xf�a󴂐��<�٤���RAp��`��ޚ��Ă�X{�ngY) �Q{�H) ������
a��2m��P32�$�I���^Kk;�
A�<�m �����>����>r���o� _|�I�@���)���%$ϮH)3,�N�) ���=y�b���c�8�k�w��e�u��8+{�=�'�. �_�'Kgw�q�5�(�g��3E9�V�3&�k�xj�����O)u!� ��Y�k�Ck�4IvG.°.K���jі.,4�ٱ��un�b6�6tV�05���y���A��k/.ab��Z��Z ��-�H���7(�4�`5��c���XYmeՖ��2��2XX���y��#�:j�t���Yx3��e�u���V��԰Uк�b��1�e��B�78&�`-)̵�!�-]dI��SQ������������sF�N8f��Ti�K,��5X̪%�]��k��+����:OO�'�m �s�4�vQ
H-{wH)h�3.f�) �Hfe�H,gܭ���﴾c��=������$������������V��Ϯd�P*s�Ѵ��R�T �*�p�Aw���i6�I��NU@P�%$w�Ͻ޽��U����4�XtaH�i&�) �P�r��g}�w[�?q�����o�Ԃ�5��i!U@y��ItB�S.�),)�f\4ϼ���5��U�$�A@�=�I�0���T0������nH)3,�A`u���T�D��3.H/{�^�}�M|f��7��w�٭���� ��)>) ��JyUB�RAaGs�Ci �fe�I�) �S)ʨ
AH,32��i!���y�k�k�}π�|�I �'.�),@��.H)�32ͤ
�{�׮���}�̿7y�=H-U�
H)��ˆ�6�H(��&|}��9�tĂ��i �U@�TAH4��ᴂ�`RfY���Y�Jr��R33P�Aa����i#�*�O~�Y�H,�e>U@P/�������}ϩ����o�Ԃ��;H)
���H;��\�����fe�L�%$)̳i���[��ߛ�|=y��r@u�nq�[ffц�م�X��e�6���]E�X�W)fο:Rt�d�t�%!L3~\4ɸ�H(}�h�A`m���T� ��p�Aw�hx���mlnN�_x 	y"��$x,�������d��T �}桴��l)���$��Y)��T ��a�v�R
fY���G�1��W�e�F��k&pBѿ� k���$��w��m�vw=���O��d�\%1�N���'f���9�P3�3�H3]�oOyX�27��~@R
~ S���L�%$)��"��'��?�W������._�G��P}�RP�0�9p�&�I�{��\���{�{y�����oZ�XoYp�A}��{f�b$Td��
��
33P�Aa����i&�) �Te.#� �Q���t��*w5Rɍj!�7��Aay��i!R�;�4�R
Aw�p�� S̸i����P�̳i��RAr����8�u����x��Ρ@�@IH!�O���M�̝F��|p�;��ز���(��>dA	*䔊 ��RRn�]ьޫ��,Sʯk쎱]k��0��OA�ɢ�@#`��%@h��D"��W�8=>�(Ԋjf&"H�f�|C]X6��6P˞�d�K�L;m��u������<%������>��y3�TGgm�[�/{�lጀ��d w)D�
#�)�=�s�r/0��1z4�0|}��T3�>k�ݜ�HU¹�	� ��RR;�L]��3� �h�O]P �)*= ��%By��&z��ڮ�sV�PDo���w���P}�o�٨�]��F�d�B@��s���?*�Q
#^ҥ�peV�Z.ո��{�k�z�;O:	�v[�&s&�=t7�䔊))�Gg�<���ח)��D�/���t#��!oW�6@����0qMdW�<�׈K�P! �����^!���^b&�q�8�<�w��M¹� F��@���>(��3������=�޾����6�i���
,5��S���eܕ�2� �\[t�p������3PC�AIMRT(�z]�v︃7L6	�<���V��S��P�8��IP�RS@|Q�'.
�	�n��ej�P(��/���t#����GݑD(� RS{ڴtiX���ղ#L A<��!%"�F��T0Qxr�:�}y.��5�W>�p�!��E%4%!%!"������v��A�q�/T�$���t]��A��� �5sDQ|J�V Tَ�rƺ���w:g.�P���SY�^E16�YwJ�*IT�Q��.��r�7Kk�d.��i=���^k@!z���F9��4=�ni�@!%"�Jc6D����5� F��[ג�l�m1xP ����IMx�J�9Z�{7���T���Մ��P&L����L�	�Q�U rjF��g6��`�&�6Ī�@���� i��R�x�s�*sP��s���^^
�W��h!Vϛs�ADA	*�JE*�Q�)j���^l�#Z�o[軮n������^�B1s�w\�\AW��!��� ��#��
�IMADEF��5v5��z�#	ٍ�!oP&�ȯ�����%B�F�[�73�ݹ$�O��@q��T�<}��؇S;�EB���"���Fn��2�G\������$�P>)) (%+h��t-��#�XO�{����\�72i����Y4-*F�R�1���{���í:j1��T`�F���i��M˺rF�N�7�(/O=�+Z-�1����b��\��/ksD#/�x{�fT6ռ�e�?[)n̶d�^�L�M�����KymK��k1M#f�٫�K*%����q�����i��D���E3���ۤYs-+���R�̡�4�a)�D�ZIA)�.6a���͚��CmG`2�M����	���UP����m�;=�����+`T�؊�:a�M�ʘ�ft�D����FS]]�G:!]E��ō4r��~����ڤBj���h�˱�#u���a��-�kL"�a+�k�f������BII��^))�J"���y=]�z��z�sOj�.��	�͐9ǣ�w���
#RS�}x��Չ�`@\G�%@�C�����gu�W=�#k��)j�ss��hA���@�ϤQ�$��$�v�L�I����a���]ާ"酾$q���JF����
�IM GV�{lq'j=���hQ�s@�B1���Lge��騼�!o@�kdW��݀�T���n����! �����
#<s'o���zB�������L+� ���}^IN��Q0=O���߼�����>KNi[��2�h�l	�IX���D�ZE��Ħ̔B�:4i�����^�2�. IM���C������>��t��O��J�ky�l� ��8��JE�׈ � x!tᎫ�R�s��Gt��Wz�N9��^��.rY�7^MҼ.�le�d8�K���r�F�A��U�����iL�G1���}����g�54 �!u�|�3��T�T^[��["�>
= ����3�����I�����<}����@�`�% ʊ[β���m��y���٭B��N ���Jt�Q%"�R�8��2�YG���A	*�R˥N)v�a���x|g�*�a8V+��2'x�i�������z�"w���{m���.���DFvV�1�ݑ.������%>I*�>�.�C6Fp���~�Ͼ��4�q٠�\�� mCb5ڐX.n��i�l��V6�X�R|=B���~{�"���T.<c�W0ad�!S
�ͳ��L�l���@a5B�8�h�Q	*�RR+��A��~�Y�D��SR!4a��Qg.�Z	���4C�"�B$��K1W8�y���n΂	D@ ���)�A�Dlk�/�u�3��`ڝ�gd����w�2�ә���/*�PV=VӔb������n��1'>�6ed�r'AD�B�j�Q�FQ�w���V��o��K5ylCυ<m�(��� �T(�PL	-�
���D9�C0|RT+�#���/�D,��*!\��p�"��C�[�����x� ��P%%"�A
=))�bg3c\y�+6D4���km��� �mO��B1��T�hҍ��3�c	�k)H��x#H���q�d�k�&G]�T
7\cUQ4�x�l��Ȳ��>DB��c+�q2�^[�b8jL=���d C>���$�l@))���Y꥾���Q�F�>��W��-q�O��yYhTB��	� �H�RRX3Qrov���B�� ��ې((�x���$�L�4�D�3���b)(���F��X	�	�S^ �T6�	*
J|�B.���p@~��V􀈿'7܌Ns�&Y��bw�odW���ei1j�q�˫٦Ny�L@=���s�ɽ�[����A=B�1I�M��I��K��ȩ�J��`�P�:�dQ�t�ôUb���
*�VB������w�}�@��l�%>���@�s隱8�w=�[��-���L<�Xj!\� ���}B�JhJ �v�3a2�sN����1TB�c�����3�����۴Sac���@�� ɖ(SR+���%4A	*�	��+i�@�>�چwS��&�U�r�D|�hНi���F�w���HW�r�l���ѯ<͒��`�S^ �Dyu��]g:�e�f[�G�"� �����������D# ��k�� ���T2�ʪ��qӚ�<�Xj��"��@���A(���Χlm��=R0����-��A	*@����C��� �f������"�顠�`kr(��E���E%5�b�C���6�S`��u�˨̶!_
�"����$�@�3vM��`��ۆ�W��h��o��Jrj��ِ��1�L��g�f�Rp��i�~�$�X��������xf�����Ks�3��%+ZB���Y�y�rt^/,ո<����ΩJ�/�����ؚɕ�-�6�;&"�x	��s7���5���h2�:�Z*=�R�%go�X�.UcҼ��N�g��W������g��]�����3��`���&���h��"}�q����&��{�F�6��B�:o����w��.�ܛ�::�,`yڑ!g�!���|}$�CLR�ܙ̇�L,NB+ Jq�y���.�����b�uw�H��ֲ,�	q���?�����=��=vp�"<#'W�w9w��G��.���Mt�i�vǪ�ȅw]8;������.��	����PE��M������o�Q�i]�VA�p�_��vk,4*���Ӯ{s��*�w����4L�X�Vew]v�t8:��W��ޔ�h����	�.�So��F�9�z���=�Nf����{�m�'��HV%~"�[��Q�g��nȏ��9uf�Z��u�g���h|=�;w�	Z������^hK�J��鑙���w�&(2E@TF�i��%�2�j6n��
L��*�0��{�dn�{�"���7��s«�Gh<�����v{S8b��T�h%�Y�'�ų���F�8�J�G����gn���M�B�x��;�S�.u��s�'�C�}>�I�7�E�EK��	 �,�A��@��(:�qz[���1��ȫ�=�z�J��N�m�ۊ���n�y�E�>���{dW۴y���w ��gsڛ�yX9�u<�Gq���#���*;������m�:;�]��Y	�r�+#�Y<�p���������9�.������/N��՝Gsj������X�q��d�;�s���Vwy�.�Ӭ�(�avۻ�j���e���X��,�wi��@6�ϙW�Q�{o�^���m��Y=�������k)���t{h�۷W�}��$) �����RW�ڬ��ܺ���:.:;����+"����^g��ݶ΋�9.mX����\W��N��]�S�9Ύ(��C���;�y�
8䓠���v�Q�uE�k��n�(=�GN~y��]�N�H��.
�t�C�>y�Y�SA۷�Qt�r��	m��&���㔵ˮ-D�S�萖l�$v��nR��X3k,RX۲؆m��m$�[K��v�t��plX��ʫ�r��P4L�nV°���"uv�^�����i��,ܚ�mĈ`ģ�X��l[�U@ش�u�7R�$��͂W"[kS��Y���/!RX�b)Wj5iWP�Z��)�9�p�P����4��`��v��w	H�pF�S�G5��:�ڄR\'[���L�x��D+��Ŷ�%0Q�icB:컲i�]�iV��j���3D�ŭb6��D�\���r`l�4094%�� ܒ&ٚ.�$lS�\]*冺!&v�4���qt\%n�հ�c�xt
��A�K���P`4�+�m5�Q��6��z�:��@�L��Crl���styh��-Y�Π����FR�����К��7f�%��N؅W0�+ye�B`��,�c�"��,GiXʓQе�$�cI[/,W:+J�g0���WA����7
��SԎ(��qh��j�ٳ03�qmɖ҅x�4v�)�۝�L�˅:�.��4cvWZGe&��[���-`@�.ű���� ,^�LV�3mp�陭�̉5�ݦe�����h�0���@kcc\��3:�gK`����.$��o#���������b����6�!���Hj`s1IHi����`.�Z�n�]���Ң��h:����&����]�����.zJe8tf�˦���(Ț`6�����׵3��@R�SMH��se��0����!�,3P��p̒�l+Wģ��|7�Զ�QO\��K3��M�A�U���j��V"�lI��i���WZDtn�ʶ�`�P���[��Ő�LǄ��$&����ʰ�P�f�36e��bm�س+X�\�^v��0�$t�ͣ�ڮ�C;]kiKB�pX�[QΕ6�!�l���EuQ+Hua��b-4ãI�]54X�6ʻej�������'I'��]	M��L	.�2�j�Λ-�$e�(�0��
�3X�3@�+tdv�˷[,�� ��m��۪@\͌kD��Ѻ8 �8L�,�!�5��8]�Pɵe�m����A-8cZ(�$�@4���f��i���F�rl��6V+vߖ�y�)�]Z�ti2��GQ&Ͱ�%��.��G6�i����V�CYB�P-n%,Ԙե�&I ͳ����櫡��s��u�qHK�ݦ�R�ƍ+)\X��-�CA�8�ʶ-��� y���H��⒡B-9�P�{�úY�P��<�tt��[�|E Ek�G�ϨD��E%"�\�Ȕׯ���q:Q����Ar2
<}6��箅1|����~Q2=� 2,R(����In��++��J�#N�v�B��/6ETz
Jh��
 �|���D��h�#JX �}B�B0|BJ�Yӎ��.�.��e7<�ΥC�r���;�0� �ȀBJ�@���@|��
Jgbʝ�O`���Wưu�bzE�OM��@��l���t3�[��}�7qt;Q35�$�����:5ˣM�ex���7:�uH(Mf]q.��E+_޲!��@��� � m'|%�s��ӽ��
k�7�]�j��ɕv�P ��G�n}I*F�J}9S��vja��p_~�:�D��Q{�WEs����i�w;_��޲�ۋ���MA4�ܥcrި� �z7������QL\f"��� ��?/�Ex)�������R���*nxN �}B�Jf�ͼ�X"c���+���6Dx��E��^!G�Ԧ��*T���[�ث�VK�О�p�D� �f�h7B���	*�Jt�9�=9\��� ���r����;�4�F�����\(�dW�OL��Yݬ��))�5B�����)�����Y͓�������}/�\V�̬���� [�
J}E�����2Sb�"c��-�*����[��Pp��*����A;@t.�#{�^���R�)*w��N��uKʉh�x�c+]'1��x��N���IP���� �D��a���fJ>d@
��v����J��G�"� (�x��eR�Ϧ��|BW#A`A�S@����T0	��o�O;0%�k���XyB�\ܛ��7��k�˽��p�	ɯ*�����:�^�X�l3 �&��f0|��=�'v�K�k/2J����1��
Jh|F<BJ�BnHn9#��8�H�Yq��R(p['\z��h��r�h�0�j��(P>�����9V�N5�9�Q�)|�浝�#K���1���.��xS��z�z��Ȣ(�%6A	*Th3w��]tS���L783���r��2:�6e?�k���h&��h���(fX�S�~XC|�2��_�O(��
R3��wR�ŗ�%NϝЙ����}�דS�!!%T))B9ÜnE��nVf�M{z�dq-��GG;�����͚#[�^>TɈ���h����H��� ���T+�%>�B3���Tp��)�wy��*�)��E" �S�IP���T�d���'���AY�(tG�J�)�M���e��=�Y�˔�X�=t7��� ��v��cݙ��?,l����]-E�Wd˯b`�dT�����Rq��kj�������缭[w��<�H<ߛ>s��|����IHQRS��;�Gݗ�Eb}#
�	���{�.�)#��	�٠A�
 �����l\ֵ}���T%4��HhmŶ��([l�u&ȴ�ԭ&an��ˀCCT��L��vw�,�3��x����T��]�p{�i�J���z�.��(�5
:2@�dz<{�k���@�}))�G�����]}��`rr+�FC��멛Y�5�T�� ��-�
))�� �h�2@��XuH�* IM�R5`w�4%nҜ\N�t�LU�RD��v�}Z� ����$�A�K�3:N��5�aohW�7>�
".싻�zM=�W�u^)�[��B�6��˚ ��l�
Jk��
!>�sE^�^�
R=\�]T���9�M� A��%("X�B\��dFd�H��U�7,B�Chh�wZt(;���P`B�p�l����3w��j���H�U�D�ɘ�Qj��BG�x < t.�&NK�Rs��Vi���t/mv��ŰW#��`3F\P9��$�WVk�E*�dGPC�S��4���+a�n�\·k�Bl��L=R]H�UQ�k!L$f��a����Zk&(���afR�a�k�ךǔ��qkl��-�sJ�n��JS[�66T�3fE�h�ŶJ@cq3][��P��EW����R[KR[e�mkV�C�6��\�}�v}����.�s���쑎HXX�&�
���Yuł"YVޕO.����l�'�w����v��`�5�s7���7���=�0E9@�=�РB1���%:A# �ȑ�:�sqs��MH�
�싾��M��W�u["��"IN2�i�nY�����P>q ��Mx���G��T0�Yʑ�杬7��Gfw8wQY�b3
��w��� RSD��T=AOVd�I;�`��G�I�����l���nf�R �p;y>��L�{4�-F�7B�IM(� �%B�IK�}��HI�H���βmc:M��w�O��#�))�IH�k7;0O^�=�&�Keq�L�Rԥ���n(K�bPiU�i��i�Q���]����y��x�����⒠�k^�����v3
���.;�'�C�D�E�E>�D���JE"��<8�Ł�3���{�>ǳ�1��MLK5.+;��6�$�˚{U6�녎F_fnGqr��Y�gA�{�S�   E �O�/��[�5�C��'rR ���4#S�D#^��tg�7T(�s@�Q)*�Jt�
#2/x����a)��;�b�d��
�W��* IM���^! ��j(��u6F%"�B0||��AH9�6�O�ӑ�U\���Z�A#
ڗ�Y[�D�	+�AIH�B>�RSՆ�we��kV�Я�B���5�����A< �5��B��%Y�|�_�����l���"u|�ø9]Żmue�Q�fl���+����#.�lԩ�6ł?�� �D9�RSC���K��o���3x�^h�]����#���׼�C��=-)�@IP��A%4Cy���/b���a8�ʅ)5�����pօW<�k�
JL�\����=��q([嚑�}�B3�*=�oH�*�j�95�9C�Y'���꿾����ùT�K��Q�e)Xn�m]��w���:����uU���V�œc&�ehۯ���x�k��K��������yzD�sF��a��S���g�E�)^@���+ť4A(���]7��r3x�^hS]@��Ƞgo����n}A5@#�))�A	*B1�3.�ێ�@F+�A�)�I�Mu��p+��A��#�j�RS@�
#-��ŗ_�cj1�b��j�,-	K��ԢJE�B�c5��G�P��jL`��@��9�S�T0�-��{J���*P	�����M�G;3��-*���*RS@�
"��[۹b���CĦ��"'WE��g��b�y�Mw��EB�@))7g�[���͠�A9�h���@�`��%A��sv0:�Dt�=q�5, �ͅw<A���P))�|�	+�[�J��;�QX�`#�))�RT(d0�ќ��t��T��N<�"�n�ɪp��Ȧ0�"TEe�%���"j"5��Mm�,�X�8�iV�ɻ��эnA��*6W�w2�*k|`�C��vҹ��������x�0|Ru�� �D�T(���oM��4j1 " �]��6y�Y4)��|^9�z
Jh�����=1��$��f�+[@�Kt"�E��s��/��M<�f��1��º��C50G�H&~��w*F�J�)
6�j!�G/d�Ws�Je���sz��4A(�$�QIH�/g��ۭ��}�ϫغ��-٨i�N�Z� ��&�#[�
6!�k�B�xo:j�"!%B�IM�Eקp9f���_o#�F`Z�B��([�A
 IM�R(�|�}��r��}�g��hP#�)
#bu=0��d�h�����%�\�Yw�I[��#���,�!%B�))�zIN��	\���8F�
�C%Y���-�Y*A=�A8�}Cڝ
!��	*vy�9�":f6r0����
��NTc�![ʪZA�N؋Ȫ��f�꣗ђ�2��U�QJ������n)m�a�m�[����Įy_�$�5k��{��IwE�^�Қ�W���Z#F6�u��3C,-�n�evQ�d.�����s*RRlqs��;[��`���m����6q3�3#,6sK�s��,9��LҜX�myp�RZ��ax;�-�K{͚�6��Ju�Vs��ڝ�*�p
�3�c�ڙ�m1e����ŮYGsba��K�Ŗ�Be�3n.a�n0���h�_S��))��[љ��jIf��g-юb�����1a��R!t���꒩4W{}���/"�$�H � V��|�
3׺�z�\Vo_iN�Nrdaǣť4A%B�����I�kʙ�Z�q�`�0�>MHQ���������@���W�Ja1=-;R�;� QE%T��@�����J�d���]��v�лus.x&�Ml*�j�>��W�F�IP��� ����%[�t�)]y�;�A���^�Q�FXZ�B���r(���;Y����C����F�@�`�IMRT+�#V/c{�x��ޛ��z'W8�tW{3E5<A"�R�
J}D"�t�1�hr��K�>Y�^I���Y]y��숸f�L��һ��-ɗZ����麽*��驝�DR������+"XJ�]R�����Hm����沽����Cݕ����Dbq��r/�q��{�� Mm-��P�ѳ�8o0eMX��F�)��\��/S����]͟��Q�4?/(�c���7N���ͧeW� ��,|u���ε�=߹�*���tB��r(�t�v.�qF���WH�����"��#�nϺ��:sU�q7��UT���
jxA`R�n���nϤvm�J��A
= ��n쌘a+�uZ9�UGUx�^ĀD�'�͞�k�HY���ݜ �� nȓ���z�c�PpQ� J����yj��k���	O$Qc����q�h:1����4*���x�1r��U�gka-���LG"��[�SD�jmt����c�b3��'#�Yg2�'Sx��.���U 0��(�|��A�"A�sDt�#v=��3�.�́K��n_����WP�eKE]S�g�ڪ:�����$�5:�4�Ό&۽=�y�Q��<A,�nǷvs��Gf���ULDp��y�{��}�Rp��վi�k��8��ۧ�4�X�3����9�Z�*��%1�^~����fK�Z їǰ?h���I{��F]��z����P_��I���oOjzT��hM��X�aH\�t��ۜ�����U�� ��7|�s4N������5{M��-�o)�*�E�@�1uur��ݖm����<ܗ����vlq)����l��~x�A�M��lX}�&�p��2 .L�-+�9���:Gz�K�vl��ډK�c�|�
E�1W��.��wNk<�$>��s�g|U�)��[Sg���:�̘c2�1���7�����"��I�(���{ɾ�W{t�ý*#=�~��3�޼�>��*�Ԟ��=F6�����*���I�;�R�q�TѓkR3��b���y�E�e�tʜ��(X�r=�7g�#Nt^�����:���1�>��[�S)�op7��ݬ�X��n'^�h�q�L9����`�$��`~�Zt��~�q*ʠm�p�b���Dt�$R�5��������Z>��qu�іnxM<йӳ�hĤ�z����V�m嗪���U<"�LM���ݰw{nD&����=v����'��
������E�{����&��t�@���j��Ò��Z�u��ό�Fi����N���c ݓD�&-�J�o�>�G���v�T�w����h�fn�e�yP��a�w�&q�3T�Z�
<��irx�bd~�/��oo^u�{�"�(�3uJB$����$��;���vwW�n��"����N:)Ȩ��{��w'eatwDtV]���y�ێ�;���u�_���eqQԗ˲��v)vV�����tE�YY�GR�:�ˎ��ˉ8��軫�++��Y�wW��D���j�a�y]�n�/lQE�,����˾we]�Z�ն�I�:;�Nmu��W�w˲�{u�GQ��u�:�;�:��N;�r*�]��u&��D���^w�pgaq�u�u���J��!��9;:ȸ���%y�����;��2�∣���G^ۻ���WEGv`�r\wߙܔq�qםdGD�^u�n丿+J���՜tIr[���6�"�� {�򳙞g}�qf\-{�{U��}��;�$n�#L�^�6}�_#��4� n�Ѯv'W[tiW{sbª� �dA�Mow3��߷�Aġ9�,^s�i�S�V��e1�������ܺ�<�ʣ��H��'�ks�#۰22�NN��I���Θ^[��p4q�vPPcH3\�������,&��W�h��y�}�����������w�nS|�ZY��t)�!	"Y�ɑ۱�E��\z@��}��៸6)쿉>�{���������jw�R��m�`SS��`Z�>;�5WW~�񢊉��j癖hF<Jyʱ7-�����f>l�W%jc��tKo?�@>8�H#[�G������b�c9��	�� ��3�l�wr-�Y���B��U�ʊ�7-B�RLDԫ���T����\�s��u��h%�(�f١�����f�X���D医�o�Z�G�{'oz�(x3�/���O���=����؝
>؏nđ��(�x�Lq��@ȟfK��_&1Uw��0)��H���R$����:|���x11e�
�baX��K̠P4�h�T�%%6�2n�Vؙ��g����)���Ȣ
�A݉�whP���J�/���)X'��*Rqj��vIc6"�#[�@�0|F�;�4}�Ac�P����4%�q✮�Gy�̝Ǻ�U�F�@v9��!�9}B��D}��'9�4�hb�{]���+�&v'9����)F5<AȀAH���D�@#v}#3��v�ػ��24GG��đ��(\�#R�������>��B���E����A�tG�R$i[���FnZ>�����ɬ���7!�M9�}�7����{�O	�r(� m�����PO߬� ��,k�g�=��z��_k�{S�0M��ۨ{7�q��{���R���^�r�ܫ���d&ʮ��:��ޖyZou� �}9U�{!���t4̷Eֺ�F��K#�%V7�	�-��vҒ�	l�s�R#�-�\�,-й�ElW����D��C ܜ�ˑٻ8�j=k��l�DLP��\G�l̜Jh� b�`�C!��JH�Zf��HW�Cc�t�WiW�ڝrK�%Kt4U3M��b36	6`�5m�G.���v�VRT��K���Ԇ$G������Ӷ4L��Zln��Z:�VS�Ǒ���e��Zh�,�u;���7ˈw߾�ý[޽Y�P����amW{)F5<F��7f�̈́�;�.>y�Ї�h�y�Y�%��v[��5W,��{^��q-TR��'�ť^=�� �n����"����m�|B0݁ ����F�x��X���m���i���{�LyR�;c�wb|A��� �y�V�_TR��`�;
 � F�
��emu����� �� ����h�s9�j}@"ݐ$wvE}���݁q��s�JvC�B�jT�e�O�[@�p8�H��P#Lx�v���P���=��`�G��G�R�ke-�mnk�	�K��f�V2����n��-��}��c��OyeǞr��(����v��K�7)����1���qu~]��>݀7a9��7O��֣{�3��].�H����-Xѯ�o���s/�~{ΐ}v���颌�`�j�;{�*"d��̚f�����]}�G����*esem}de(�U���=�-�;Fn�����ʀ�Y/�f�� n荑��M�U;4�!m��ŭy�؜����{wg�z����A��Z~�b��D}=6�9J}k?za?��@�sC=x�-�Ӗ�|���o���3���Sl��J1Up���n���ۜ�k�F��Sb�LYFMTH��v��b�%n��ш�*��ks6�n��\�~��{��}�v�v}X�����,j��8$ЮV��gm���w�֏����)k6!_XK�S���}����{����>���ޜǑy�k�wK������7\@�wD3 �g���Ce�r��L��x/˳��.����~}�׻Wl��J�3�Yʵw�쬾P�%�:z�6�_ =�x֩ɟ�����eb����p7vG�`f�SL1Ok���\r�7vE�)�W������./�K�>xs;�ׅ��2�mh"]ѳ���W�W�X�}�s=ߍsΎ��(~�h��y
|���;��1Ʊ ꑶչ��Hgf�!@�9���:Z�d�X��l��5$�9��n�ݏn�{jUKm�_�&��|���K��"8�Z-m!��b|l�^9���ʺ��~��ӎ�̀-9�C�l>f�ྋ� w@������S�N�R�n�zҺ��/��ˑ� ݏn���Dv�X�KOw{�g_�^Z��oVԣl��]���� �]�"�<��SՎe��{1>L\��ɻ���Ը�Q�(�`��˛��t�F�$��:�4vzn�9��	�)9.#�{��[����$���2�� �T_�>�>�݁���w�ep�B�Z�g'g�7]e����V��;b�li������_�v��o�5$�:>8@�>ѭ͋���0�(��떪�0���]��ɮ�1�?{���~=��#ve�eu;�z��f;�=�A���{��j<��ݽ��X.bfp�(�(-Jr�<�ԣNl��.����
J��gq{��������V[k<�&����/�7[eJ8�����?�Fc��g����iOEE΋���۰f�eSwʒ���\�.c�k�9��qZ����v7v}�-5�o.�]ki�Vu��w'Wx]�Owl{u��z�'�'*���/|Z7'\�.�ە>O���jUЀ{�� p������+��,�5�
�,�y
ܙ��vL5*�����������\F.��d9k!��W^5-h�%�Q�L��E$��J�T B���tcq�[��<�n-q3�飁)j\�U-�LS�9��+Q16j-5�h�d]-�&e�B���uz��2Xi�g[�5Π�����Jj�WU�XF�4a\2���q�!,,�hd�ܦC:����ѰC	�,�[�Yilk�bǳcXX☥�qSl�͝��s��~/+�JG��(KhVJ�X�K@ZX4���	kz�k����������[ n��Բ�-_t�<Ǣ�_U�"�T��V�/�V�vO3�h�i�-?=���ף� ���/7U'|���9���۟p7g;��5<*f��%��ݝ�ݨ�T�ծ��Q�F�m'+$fy~�1�w�����2ш�o�zZ��N����4�]ū��y����nD�n�휣����Q����-[u�+�w�vU��<�����ޗh�w��8�fz�E�.�9���i�R0p���uf,+�6���X���	�R�ۿ�R�x�0 �Ƃl�+�O��w��n�Y�W�F��Ң�\��j�9��{���h̶��S�w���ڗ�3�^��;pv�D)�ζ���0uˀlY����Ϳ�Ðy!����G]&��m�)VϢ_��g<�g���=�>�� .r�%�n���g��3wG���F�I��n���_m�����lxn���wi�����j0�]����plZ�s�Y>{v7wv�M��1y]>�=�=��C�W-�9Sf�qUp��%��\#�j|���#�v7s��K��CWw��Q@wr{F�o�&y�8�������J��~��e��~��K�ˣj�y��nɊgZ@�h��d5ns�\�h��\z~��û��߽����mgvg&�LR͇�u���Qfsl-��ݝ���{�rt."��ν�tkVO;�n��2��
��q��"ۆ)Ed �Ϸ`���wNp��
�j�e�FUsOF�Z��e+��;DuV(�G{u� ��~�����.IYz����n���iU�>��\�1��Ps��m�~����c���Z���׷�cv=���f�y�7�oK�Ͱ7cv���u�jt�"��2��[�!KV5\W��~���h��s-~���CA����ꧪ��\Z�2��U�	���ۯHȸ���߰�l�(��W9����pJ�ıe�����&Ȭ(����
���u�s/�_[L���6��랗�j��^�����9C�i�p��m���#;g��zug3�>�O[]�ݩ�Q�\�e����/���{.\�q�fw�i�}j�����# 7�2����Q�7® N7vG�c۰=�8��c/ω�w��S��_M�OK�5T{1b�Ӈ�o.n����.*a\qى�k����u+Iժ%d��yyTv��F��:L��{���0����a�v�d��G��^\��8p����+�����n쁻��؁��1��[��K��N�����Y/cv<7v+��'��_���敆9��+��n[��q�Yn,f"4���4�&�̓f�g�u�}���߿��d��ڌ;�C����vo��Pp�=Ί�{m7��݁����ow_w��eD�8�9��U����^º��.=�ۧM�j��Y��~~�����p~��>��%x�=�z�$b�����{v=�ݑ�v<�Ȫo�*��y�݁oQ��Ss=cݳ�6�Dw������h�����U�1��������c���F�����;������5�K��؋�~��k�f��4�UB�t�]��L�;LG�Z����Zv?��ɑ�O/I�={`�Yw?-w��G��i�K��(���,���LG�����=1���cӊnv���hp�$�fK�-���A�U�w�lX�D{Ѯ<���:�©�.&d�i�ЄHb%�^"���p䫭G�UiS$`f�L�	�P�&�0�de9UZ�w��h��KCB/�=5�n� �������lb�w}�w,��68)�޾�)U�'9���z춁9{ئ��<��9O�e�J�Țy"��0�2�6��'b��ń��xe�ʕ�a=��x�c1�rE���í,�յ���Iհ�(>'<��Ç���1m�n�+��ծ[��������{�qWV�eV�&x���߮��耸%A�X5�y�<��Y�$����L�}��ydЇ�<�9�'�ϋ2l�2�K����t��&�tQ�U�%��7BU�%�M�g�ᓬ�s�z�|���qKЉ^ɏ�(������+��j8<
�B��`�;�$�|�����Y0�=��!=�.&�U��C}ە"��Hf���t7=,��%�����ٯ6�����?��÷�h��p�����V,G��6Y���r��]��;�N�sP��諭�Q}�d[���n�:��ĩW�騗I�Z������@���N��3x�n��Qj�:#sӄS	ū�2S�O���r\_so4`��&`U�]���%Ve���A���v65B	Y'%DKg�Y]�z�1�͒�2A{��q �Wu+�q'\E��m�+3��*���+H��
<��̸�䳳:ｳ��� 룢��E�_�W�Q��)�㨂����ˣ���8�;���;�_�yQ��u���y�Q�e�Wuٶ�K�#�m���wy��[��~~��:|�qϖ�;�80��+8J,�����^Y���^WC۲#�kﴉ2��|����p�//:��8��i,���X�j���\�|����@r���QQ�Q��˳���s{��G�Yq$>���W9�gW�R�[)*��`�m!B,/��FȰ���(��3rU�������;b�i���3Z�j�є�fh�t�2�]�&0�[��%	N-4r�u��2�6�Ln�-l{)����Ή4��G�!d0gk	�`ô�UB�%��f,�6K��i�]�=����o%<,s� 5��6:��ŕ4�W��#�M�.e#"�0�J���m4u`��.PJaM@����uH�����c(7�h�e�)QҚ�ˮ44T�Zl��Y��*݁�%�I�Ɣ��6�(Z��]v�,70X�&f�r��[�q{5Ց�3�U�j3�6���[��
b���KH�t��ER15�Qe�\0�%̹�LA]ncf����叅�$|X��u33Y����L��Ìg+v�	e��Hu���tD��ՍW6����-�My�4�ڥ�6��Q�����tЀ7[��ZF����<���R�SG[�����^�u����L��cdLl�2�Q��t%��������Mv�U�4�!v�0�DV4�Ʃ�0\�Z���L��]H���[K�Tm��[!+����R�$0�J4N���G7C:��&Lj,� ��`����3af����9j��ie	U���Uqj�G).�il�3LeV�������h#a��2�u���LDuٛ1�B%Y���e*��7���-�F��Iq�[v8T�K.Ҥn+�s� X\WKe%N�".��ιqa�"�9��YfcsK�lYD�����dц�3M���IU&"gQ�,/0�ɮ%�ѫ�E�̉���caI�#�S�m.T��F[n%5V۠(�ŻKQ77D@#q�l�0��٘ �e��1���0h�h�k��q�s�:7U.�&�*�hL
IP��\��A
�Fˍ-���+�s�F
�K��a4��ccb�Xŗ�љl�v�D��m�]Me �PƆ����,x��*�Gbl�d���V=S
Ѻ�;8ڪ�r��]U���s��-�Vk�C8ю�Z��$�`��f�i���J�Y���1�Ķ���cC�|0,f.�d!Gq���l��lGb�v](f:�K���1�&{�ZX�-;M.tp����v�)ЎkG�,���P�*3f!�v�7�1[B�ԙ���n�Թ3)5��V���Ɖ)�V��ڭ�A@3���Ѫ3,��m�MK��΍�M���������\�F��kc���;�+�J��XfV�a�d"��(�z�?��z{�{ׯ[���v�{k�9H�-�<�d�M{�����ݿn�nKn�|���:R����-�.��nb��EG��r�wl��v �ԪI�N�D�n!(<)��+k}��k���=�JS�Sç�֌�Ǵ����)��s�ܹ���w�Qv��;���-��i���������e,~w6-K�s,�s�.��v��WA����|g��OR�XK
P�E�Ɓz�J�*����&�+�T�(�c�L�jz=Gߌ�	����~�o���7��Emo �ekScsf0zWO�F�ݑ�W��e�K6jy�*i��h�T�sje:��lև�澯j�ďx�zj���
ș3�>9��-���3�Y��0�F���iT���3S��y���mc�|�|���:����s�Z	�rOt��kF���7c۷�7�nヱ,�l�N�/��N)��?|���i̴e�i����+�f��@} n�n�
+������]��e�o���ۙw�c� ΁��� n��	o���M��w��$�(�Ůx���7`n�8P�X��D��D��vj`@ڄ�l5�3`�D��ƾL�cn�	���GJ�`��%@��3F�T�.6"�4�����1��}����s-Z3-��1�3N��c-��Հ�pV��ywG�w�H���R[��L��y�ݍݑ�⧧]�ŉ���v�-��gɆ���0��Ȑ���D�mp��v��f�.�-�k����{���*��Z�6	ة{2��� �9��\�iڈ�X����Q����Omh.�`~��ۙ������	\5L[��ngCU�yu?G�W�X�s%���~�E�|wף���we���Qzr�m������n��{{�<s�;I[�٤�Vh���S�RV9k)n̤/[f���͚�����h�Mj�?|��$���g۰N�I۾i�n"�c��Σv�����P�#v=��,�XN��5����c�K�����;. OwTjY�m��#�����3�8�-[J�ÿ
;xpgZ4\�O췆~�ʺ���z�O�`���Ƚj�+}f�{7�_�r7MVsM7�o)�r/f��ѓR%��[��K��#6��|�n��{�u�^�_�ܙ��@���F���jr�V�0M)5nT3W��X�NC�B*��T��x'�O�ݏn��ߍ)՟HKö����b^ڪ���p�ݐ7Vѷ��_Vϟ���5�1�͆ή�kX���Dqb�ҥr�-��p +wG���_;E��|�|��l���U�v\n��U�2iA�����F[M�ޒ�vO��i����wzy�M6P�X����{�]!�������|<�~�'�[M��WI?��D�ޚ���;��lN;U0ў.<���=��3��)������>�7v}��`�*�_g�)�����=��_��m9��=�����Z��G詮�{����gV)�� =�n��������W8�o+y�n�3`Tt��4+,��}aYtL��&͜��+��]�e��G�~���~�ȅ&y���6c�d_le����3��k���y�Ϥ!�7ƭKe���պ�B2,�Tn����(���p��L�jumƬ"Ж�@f�!ue���a�Q�4ں�9ѷ��e�H��3��m�XdҐ�Q���E�a�JV	+Dׁخ�M��W5��1�ۍL�h�ف%k�\��ֱ0�K�[�4���q���f��cv�ؘ�q��d7��	��J&�Q��eֈ��J39_��'Ϩ,FKsF��G�m-6��Ty�.�����\�X�+�C%��[ԤnǷc�����2�ک����t��];�7u�~��v=�� �o��t�z�ͱ��wQ�k�٫��.���N�f�.���U���xnǷvF�z+�4e��g*L��䖥�J���T��Fe��4�t������0	�����B۷[�2杪�jc��]M����ٙ����Q� n��n�c�_k�Fݮ��T�h�ý�7u��N�{o����?o�f�x��%�H	4GR���f�cu�5���˶t8l�qh7b�ι����>~��v2��t�\�ǥ�K��[�\�S�1��8��P���7b80�@ngBcΙT�d�&tʠ����e)��.�jߥ�� s^���p|�մ'��z��Sr���� ���x��nG���Bܾ��Ր��T51�ˀ5n�kټ��:S�W�>�����n��£*���z+/6$f�eG]���v�Ȁ�u�3�G�� v�ݏek��v�lk��l�����"w��t^��V�j���ݝ؛�\�}��x�OX]YԘ����T51�q�Q����ӽ��x����~)ZD�l�f�.	�;X7,;(�v�l.vmWGML�B�pa[�"q-1s?gp�[m����͗Č�̨�O�e���s���7vF���M=�q���uv���tR͞�}�7o��m��=ш}��_�k��)���rt�A/��c�F���Pg���.����8�N[���Le�K&jaHT���Q�ipܩnQF�B���n��

K��f}�.�\�������9+�mƭݿn�݁�R��O�.��Zz�}m9m�?s���n��?cc���������j��rі���Ry�)�\n��>�u�ݍS,%�<=8��{ݍ�w��|��w�0Fm���L�hGa�� ��(�L��A��,pb�l���T�����K�=���� $��Ϭ�z˚٨rW�#yj���[�Gv�j�ln�׷v^t�f�p�s8�=�JF�������gr�����l��]_M��j��U~Y����ݝر�~�K+��U�v�La,��	� =�����ݏ	�n�е2��ؚw�$�����3�U�ܕ�r��O��Gv��E9�{Ή�l=?I���f�ɳ'J�ƃ��iݭ����պ�(���)��d{/�$iQ��'��Lଭ��uP�c�ڛ�� (�����݀7vF�飻"{�y�q�-��a
X����ˎq�w`n�霂�;z�����M�V�ⱑ��;-�og[��ŏV�������H[���߲��-�-����]��F��<8|���Qo5����v7c!�0�R��Y�`%���v[<��m�RW� j�7vs���&3�M\=q�����۱�wm8��f.G��v �����?cc=��h�mۊؖs"���� n�%{=ܞ�Ob��<��� \�c�q�x��v���Q
�<��^+���j�g�ҫc��V2��iϭ��j�gf��?�X�۽bf:��Xj,T��A�֭j�׎�;b�yoCn����Xg�Cs�w�݋�M�1?{��q2LA>�N)�B�jໍX�
��iB1ڨ]��6��&�C�.�[��1�e�,����f[*�%�b\L�/,�h��T����(��h���5�H�j�fZ�R��[-�Ҷ�S
.�G�te�cY��
�]��Tש��*�ڎ�B#�	-"�4BQj���Kq�\��a�I��n�m���؏V��o%H7.�A0@���a�S��a�5�i5/ZU�]0�4n��v
���#.Y��}Q15���jF�����ݶ"�T�xaU�pW+���&=]��������d��:7+���r����]���B��g�)H{�˪�c-�'՗��^*� n�o�_{\���{{E���{�g1x[NZ>�~��}�������z���mw�c�ۧ3�
�ˎy�\L@ل[&�o^��Ϸc�ݏn�[��ʮ`;��/�v��pa��<%){�@n�67T����d���,a��Ů]�l)aL[�V^�tɂhb�n�p�&��0Tw�lxbS���E5P�C��6yo~�*�] RZ���ᗸ����ȹ+Pg�O�7���2�Q�kZm��K�y�X�eњ��F�����r����Z�/���ٞ�������);D]�t^P�/����n5�����?+7.;�P�ס�����h[�둻����9��6�Ck쭗�=U�Ɇ�l��7cwg۱�j�U�+�mnE�o��f�]*+���{.��G�Lӊ@N9N�ݑh�?���8���a|g9w4���?�~������F[�����h���6�v��&�5!�s^��[��2�;��-x�"i& �E$�I�ݾ��wd{vs�9���R{t{�S�3H�)�`�/ь��[M�ۤ�=�{�*�vą����E�P�����U�+o��wx���!$�m�n׳T��݀7u���4��h�T�yB\Nx�Aq�I�v^�����o�i�p����w��}|K���g|0KE���n����V������ovoC�#��{t���h�W�G�Ї]����Lh��IQ\SO��o��YP��-w-ų)�P�~b��/�%x2�{=ڽ=��"n�@�pxSW8��ć��P��(ܸ�4e�D��*�4���������.�^�����xj����шB�1l�����aѴ��4�����OnP�SV��e�g�'��p� �4崯gQ�A|��FרS���.,:�`^݁�w� ��7�rd8	�4������qq�oz.��stޖ9���Z���;���.�j�i�볝�k��l𦍽���h^ŋ��Ғr�z�	w}��&&u�,&�ע���GX��ĳwCgP5�`5:}Ⱦ'�N}��z�0����O<0�y!��S@_Mtb��DJ�7��i�ؚ�jW�n�E�[�����y��2�:��\�h�7d�/A��տy�l�QG�%�b(g���^�4�����="����s�0� B��]p{�=�roҷjc)�Z�Mcٙ��=�Bh"|����x��[4�wLR����З)FCZ���l��ڡd�5��fs��#�O��OEu����v����������f�G4�={��N�5���-D�v\|����'�X:'C�'i�3tq2�T%�J��W��Snx��.��-��g`ݾ��T5��&��LN
���vZ�f���u���f��IL�i�����w�Ď����#���.+3ӱ;;I��oz���}�����_��kk;���c�#��
�����J:�y��;���{]�G�ɟ{t�N�����5�!�H$ĕ�I�%l�;�i���wӾe{Z�ս��8���������~u�|�e�;�E�۫3��ggtiܝ�t��e�w���������2���Zw�̨���^'t]>h�.��=���o���u�qrPe���k�}^^we�ү,4�.��;���g{nzݖe���D�q���W�j��V�wߵ�ԫ�v[m��
�(�;����e R
DS�B��|_7��{��M5�xU@l�ǆ���b��N�u�#v���;9ec&Z�S���!��N`j���y5#v7`�ݭh��;<⪛�:Q�jK}�&�j���Yأwwn�7.���YQϰ���	"�d�5�l�`������H�El�1��k���[[��<?V܎�������]��p�r����V���zX��4�{�-[NZ1~˅	��
��e��f��s\���������~�����x}�;�9��xe��m�~��.o�fp/B�o�߼�m��t8[O�m�W��/�_]��=G�Ӄv�v�{%�[1�]j��Tt��W^�X�iZt�~��8��w���C�a@��+ܱQ{n�M���:iƙ�gշ���<q�}7q=w�=	
��f�Q�� <���7vF�xnǷv�r��;:�q�gٛ5���n͵���%)�і�w|X�5��'w{I�Pӥh'V�6Y��nR�6��M�h�>9����,PYk�s���7���v ݀�����*�jj��0�j��8��y���e��m�
W~�+�j�=��.�:Kp�c��4�n��y��8+�1z_;E����<}��8���]W �s������=������ ��;�m���݊�ݏ{��Į�u;pj�I���LV[�
��z}�Z3-��e����N�CY�=�����]�	lGS؊��v�[���^rZ�A�'m�[�e"�j:��BE/b�wy��3=��/c��w�*о[�y�.NX㴢+����\
�,k�g���Ӥ�����%�'�;[tS.BGK(ce��)*H�׳���������F�rR��Mi,����4�u-�/l	[�IGE��޼�$hcGj�[�U��=0̀mz��i�Vj��6�s�n!�6٥��f��Ksk[.��bSZ�AjWk&���;j���t+
��h4�����L[��Jg�sr��ͱc�R������u�&
�%�ZW� ��bͪMz��s#�s��L[���h�b.�_���>|;߿h݁8�:�b��a�����r4fH�u�I������[M�2ћ���g[�yĮ�u�,UZ���P7w���9T��^ǹG���n�݀7u��ǒ�U;I���+L�g^�p��{�n߷wv��-ػ�ݶ=� J��4��wl1���JH��)�*���I���Ƿcwws�LF��=�1��ȭ�7�Vj%a��{�wd{wF��_p��WĞz`�ylf��aśYu�crw"k.��f4�W̪Z�#j����r<�����Z˪�l��̆�#���t��M�X���v����D�AD�6]�Ѷ�2��mL��e_w��(}��] ę��@ݨY{��o�:�淫�#= ؑP2��8e����7�Q�z�nϻ������Y����w�T��wt�gA.�6)
�8�mo_X�6@*��������������{r=�7v}� n�x�(sV��6	��r��7vF����l�s̆���JX�s >m�m���F[`>G���6o�o��jy��npxm�Zc���z�G���m%��v�{܁Ÿ+�]��#�&�-6	��@�u�l� �46!���e�S�`����V��v��P�%ݮ�Ĭ���Y9}�;���?e����j»��:jCp�ݭ鞻�h���u�ͫ�ߟ}��{WK���?O�E�۬(u�3�E�A*:gj�)L*�KV�Zz����Lb@�[0LP���^��)ڐ�,}�z���ݡz�`xKo+�"���6I��x�);�����ƴ��x��������G/.���&tg2���*Q�}���ڳ��zX��\?��;�h��~�e��	�?Y����f���"o�������n�ݵ����נ�~OI�¿H�h6MÖ<һX�3����&)��.v�fh �+�ܺ뎹?����O��ۻ>݉��.�8:6�1��qu:���{�3`�ݿn���{\�A7�װ;��+����jLN+;�n@�wX���t�c�����{5O���xn��-ceT��k�3|0��8]@��67`m� ��fg܄^�|`��?e��{�/�Ì���Zc��H�a��NI=��{r>�p~���x8���������{����U����߭�)��[�E.=�Cٝ��:7Gz�9��w ]����:~��}���FZ-��?���g�H��_����}���(�7��Ή��i��Ώ=���m���H� �DjZ	�3qB�jfJ&��)sr۷inepF�Ƹ>�f��;��{����zs�Zjo��#��xdH���D�)�m�-����{A��z�Xۜ���N��=7�8���Ֆ��O�M]�v��������=
�V[���=�Aa7��vr�i�mY�M���RFK��3�7w6�����M��� ���<2�f�����F[Ne�7cwb���Om^#}z��)읔)��N��;ޛ���v=��g6�]D��je���[+q-b�ٲ�S*�L�,`Kɥ�_z�9b�ov_wwUt����=�e��N�o���vm��v.Œm*���N��l�ں�����.���@x��Z9���֑D.���Q �!kZ������&bj�����]64قM6,��!+	Xj���KtKr],�J-��a4�[�s�,�0�l[�Ic�h�6�f[Ý�X�û8ȸ-�/Yf�mM(���5b�`�bY��tX\эX�a\5Ԭ�qBgx�5̦�]I��t
,���)�%����L�.1�p�]��������PqZ�l5�T�w6�e ��K*�>�w�_2Ɗ�4�4���s���s�t���v���o8:4&u^�e�˥�w����-�� n�݀��(��
�r���9�^�se���y깎�;�?[ �(���<�X�e���-�-�&0�rT��d�y%��N��;ә#ޢ�����D6��ߎ���(s��}�����ӳ*�	bDΫ+����*���
�j�}�Y�Fe��h�MG�������F�=a�B���fxU@�.���3[�����P�in�-t��]Z������V$*��a{U�!���vL�l5.��Qf�O���d���φ��r^�I�8'u�֘�9��4WT��� ��7vF�xn����D�C8N~Z���?[|=�Ȟ��p%�i�>��M]a�(AƱ;���)�2v�=��˛��n�D��^j����p�S ���ybu͸׳��/���(��䢗ճ*��X�3�����n�g��;�Ħ�_����[j����f��4�cb����W��Vk�*���}m��4C04
�l�o����zOQ����Zc�us��)�!�|?����F}m9o�/�f��_VL�]:�����(@�>INR����~��un}DϾ��	�2jLɂI�r��G�]����6qF�Y��T�Wj�d˝[�?2��4}"HJ=!%B�Zs��p��_agU���vTv}�,�������^���)D�BJ�@��I3�[�B�ճ@�ԉ߾�=��?O�[��K~?H'/&��HK{���_X���ﺅ��Q$�y(�(�{��WFB�%j&�~2h-%=�����S'���3K&�=���Ԧ.�0@p����c�S�����5T�iχP�L��b����u���j3��ʾ��ȉ���
P�s��%"HJd^oO���#�?�O@�� ���JJ���;}��'��+�.=�7q �EF=��W{�?�|BJ��@�R� ���qS2�h������|g�-�ܥ������I	H�$�U^O4��B����UG�T�x�0I���E��(^CV�2M[���`n�ma+��S,�Oߺ��j$~N��H �����WR�ϡё������ס���뤮�c���wH���x����	@�RS@�+�߳��H��+�O���Pձ���udO�!�W�\{�wA?�P)Emd�Vè�X��/����$��IIMx��<�t]�ߍ�ne�c�O	n��-�D� �̚�D����j�%=]��8>��ڛ�̈́�E�H �R��y���v}LT�)|1���I��ăJ�'�����V��ϼ ܁��=���nW�)��Ȓ��e͝�i�WhDnvm�< �wL�1NgF�S{��g���? ����N}]�$����J���Ң*L������ ;�����I�����*����&�$}��B�Q> ��v������o�����4�`M�^-�lEk�搹���t�*�M\d�=}��Y}}#e�=�� �R'_��l'����zi-�D�$Hyv�Gu=��K{����B�|'�$��F A(�<�&7��"+�@��'��<���m��e/�9�P � �p$����ʧ���>l��Ă_�hJD���|RTc�=�Mw�l���j��d�.����A7q�wP��I�HIH��ln���u��:�H��J�G��=2�|"`|k2k�Jar���A��$�q��]B�J$�
Q ���)Fٿ��J�6>�3�ŀ��{I�}��P���G�l	��$���!)=?|�_K����ڥk���Nξ�u�e|i곺	�%�yn�,���E�Mm�5�%�W��[�pWop�����k��ad��rf{��vރv�������pg��B��́r,R>�ׄb�.��0�t��.��z�5�� :N���a���q��4�Tx��.pf<vW�}��h9���y��yn�أ&�a9"�e�#�{9�v�'a-���/dB��{.��6��aG̚*)��pUd��n�P�5���	�N<����]���`�s�l�թܶ�����q�KJ#�	�ܡ�sڦ�L�2�(4Ӎ1�����Gu/{3��g��O��3!���q�e�70���s�w]\E��JAڃ&u�^[��)���n��\ڥ�ϛ'u�XY�� �f6���G���G����'�{|u��6��t�b���w��Zz�i�Ѿ��Sk���8��c�.x�z ��
T�@"����E���!T���\~�����OK�^/G,^w޳��of���8��>����#��F�������;���=_Hـ\Q�K2�kfJ3�82	�5��$�|��b�f�|ޥǻ��ּ�^���wc霺��p�X���Fx�đ��ӽ�{�ձ��Jb�fxN��$���gԽ�]�*٤wjܰ�[�S'i��%z�{63�yr[} a�گ$�(���ٽ��k~tg�E�9�i쳾��-��y"��1��yj��&oh7H��NԨ)͵Й�jE�ś'#�ÝRΪɓ�h��Y��$���O�\x��Tہ5�[>��2����o�����
�7G�y|󙰺�x�աi-UD�R[�;��wq�]�g�u��Fu�k�������]/�e�]ֶ��d�q�[�"�+����z۲���+���r�.�mQG~u�~V���<��'�-��;����+�;���yg_2�$�}��üΒ�I��w�v�����ڳ��H���/���e�����ݕ�`�ey�5eƶ��/^ם�縇<�ߞ�y���W��w�^��[�q�v6�F�{ݜ�V��֢/�y�rwm�)�;:��+$3���[qM۶�q�gVY�[޼G��;��枢1�L�4�Q�F+h̓C��wj��{(61 ��(ڛ��mjg�=��޷F歺�%Yx�����C*�a�p���sn%2����cJ�K���Cb7uHA!e	t���T���{7��� �5Й.�k@f���st�f"���B���.���+R[(S��32�\A���N�*5ف@BR,�k[!
�g���JrMԣ�G�[.���f*�҅���gu�I�՘0彊�JԻ=�Y���Һ3f�YjkR3L�s��G]��L�EH���[̔�\+
�a٪��mbj1�[�K.�nĲf�U`��)c�ILh���i��\�t���5�kh�IFf,ΚY��ٶL���	�U4 -�"b����0���ieٛT�C0�"KL�G4��B�]�����B��,l(�&B�Ҁ�1mԃLF��j�B�K���q��;�,4[�-b��HlM[5.��n��H�<�fͼ��[�u����fI	�����ݭ"��3����	4��J3X�D���S�65��bY�v,���c���"K����u�4��Jb]�ͥH�X��������U�����\Myf�i�K\��5�,]P�d"��êгË-�m�rۣ�ĵv"�ᕩWM�6�5��f �d��!���r�R�^��e������{lu&��,.Ћ�⌱1���2�����Fkfk��C�:��G�m� �M��@D����@��Xje��-�&�ݴn�p��-��L��֚�ūjn�M���iIL��.s���Rg��\�\�3���g5
,͸���Uz�b�J�\H��%\�[��6�LZ�[Q�4���s�NͲ`�kGs)��T�+�&%�B���2�U��&�,Mv���TX5�4m�Ք0/l�ji�s�6 l�`cm��C&��D:�Yf/�O	��j���6]��5`-��b5�c���
��[��ء�W(K��M.�u����e((@useq�5��ʷ+���.�_�u���n0�+��M�	<�D�]��ҏ4*�)��r�%�`۪��g*���rW���ek-b8r���Jc���b]�e�T�9�(�7bZ�i],k�l6h�%A�K��\7���k����b�i-�t��4�]kh�9m�9�]1�2.:�1��kq������c+��'�$��h��@8�۱��Mɣ�g��8���� ���}���l���6�K�mx]":�V��X����\Z�Aڕj#���$w��� �Ϗ�T;ӣ~W��,�f��}�����}[}��߱G��^� %��@��	drcD.��_ ���R'��Q�u������RτO�A�&� � ��|GĔ/���yʅq$�'���%A�J!Ϸ�s�[h�Y��~�b����~��w�IIM�	%2#㑰�B�z2]mN���GtϊJ�D�G���r��w�\| �ǯ�X��}�!Y?w����
�S�g��H))�����/j7ԾQþ��_=�+~|O�"���� �̚ ��D�BS>Ԥ+ė�������hJ!�"����% ���fe����x>��&���j��]o�߼?.!��������ZQ��/�}s���}�!֕�	o�$��^��!)�RSDEw#�'�_VU��#�PE�I�(�J���&Y�,�a��컌��(�ݩ���ɊQ8�>b:�/��F�]r�hm^���#y�#�QAg��/��>}�(j'�-�����*�9������A�%F���b��� ʉ!}�@���'�%AIO�)-������ȡ_?���[�	_�f���� ��BS>!%B�Q$}
�6R���?<�> �j�x�%(��J;���~��C~g���@�(+X��됳s�9�;��s���+�|
Jh�	!&����j��LW{=��+ۤ�9�v{�̧nc>����Đ|���H>J>�gn*#�0�M�X�v������JT%&Հ�Kiq�&npb�M��dδ]ۯK��hc�h�̢����A��|�=}�̼������)�־u����۽��Yi��.=�th��g{V'��##jv3"{�Y3���H%��|�}�����VP߃���7�$��H))�j����^�ˮ���H�;dH#ǹM
R'�%>����$����E��_t���n��
�ŵ\{��ӂ���4K���ٺ�Oь�� ����QP�Vg*�j�H�U����!^þ��v�3�\{�7�)D��
Q$$�P�+�q��}��p�#.D���h|����)�?qf�\BW�g� ���"-u�ݕ%�R���O��B�J$�(��T(�I�l�ܾ梇��l��K��oY����������RS�JG|���e??^ �ݻc�-li7H�P.e�e�=����EHfٖ��֐�2a65��~����XB�BR'��*����[��ۖ��g�q�.��)VM9�9�N(��}B�(�	J$��^)@�����c��z��#T	���iwG�m��U�*~�|v�h��D�L�P���M�w#��j�Q{��zRT(�A�}}?7D<���[?P�Uk�f�qa�S��o IoH�RS@|��!(�f�}w�Ñ-���`��$r�$�g��?�ӹn���W���q�	�W�}/뽈ȼ������v`���[Jk�G��f����6��+�`�Ǹ�z~ml~�¥�=��f����>J;�����}�$��
�|BP$���{�f#"S|�{&D��LKy�|>q�V2��S��[�DR$���J�n��ןV��p��������'��VT���È�4�4NմP�B`v5i��f]�ҬB�2c�'�j�|�` ��b_|~�߾���\����P|��FJGG�=@ ����iϩ)��H%%>s�V҆%֚(P#.gŷB�H\\|>_p�v��UǾ�'�?�E���R��}ӱ����+��$���%8!)��W_E�rn�}Y�G���U��	�3&�<�O�Jg��*R�j���#�ؘ�(��e
��R�����?�7�po�^@>���֠��5(Gt�%"A))���$${u���'Mgo���%�(n���w���N�WM�H ���E(����b>���0�υ�2\Ӝ�F�Kϧ2��E���g��ӮJaRݗ^{:g&v`��vM�3�w��srDL��iCk�ꊠx>�g�����]6�b�� j� ����XĶ��%Û(#!A��vH$Ջ�ic�rжt.H��۵��[�(.�[0cX�4VQ��B킴��\L��Cs���R\;L��C�d��H����͎lt]5l�iNS
�\C2���*��YH�YPܖJ\�],e�]e��&�,u��[!�4�M`Mi"@���[�YT9��lZd�б��3e_��e'�B6-��JR*��&vTD�^�b�t�f΀@҃��4��������?�>�1�%4>JD���:y��2q��
����^/��p()K��"H��|��E(�)D��%�Xf\l������J5'��L���Plo��	 ���䔱 �_p���H�F�"A?/��A�RV'�-Tb?M���C���'�ګoh��pT}�_u
�)D�	J$���o�O�Ie������N	H��|:�8}e��p��S���!E��nO}7Sw1I����J'��H>IP�R������B�3�l�^&~�N����(�]JJk�����{��_��m}����V�MS[�3�p�!�Vu�F��)�i��K��Hֺ���w��ϳDR$����T\���|w*������v�E�t0�ϤP;�$R�$�� �At��iO
��ɮ���;��.�R�/t	K�&6���$<��]�V���im��I;�+r�z���iQx2ئeI�����������
�c�W��xU|$r�h��D��K�5����G���I	)�Q�(�q�_.�"��g�z�8B,o���(yH>]"JJh	H�BP)�Ȉ�R����.t�5H�Cq�IPHK�����yZ;n=�5�>#~Rغ����9�>>�	)�P0�	%5��$�"#9�*�s�=�/���l';��H'3'�9H��'��*�3yW��t2��بM���k��ua�����]b����7��ճcM.��U����8�C��������AJ$bO�U~�?J�E��8��l*��Iߞ�*���dY"|Rs@��H%>�JJh�T}��0�g�4��g�|��I�r7��)SՕ���>ˉ���@�i���<�F�ЯxA�Ϻ�S�%)RS@����k��	Ug��Q��Cm�U޺�	�R2��XN��b����RSې�M�w2��<��1-ƽ���#�����LF�ų4����a'�_"�u�Æ��a9_���H'3'��R$��||��E(�&hm��5�A�T(�|R���u�q�U9b,/�EH��@�'3E}v�|���!�j� ��׈J��h��뿳�Tn5zw�^���Nl�����������Ց ��u
(�)F���쿬0~�	x����5 �a����6PH�]ƺmu5J��qF(�ɯ��p�|{ p,��!(�Ǚql}���0�?�W�E^\������s@��H���䔌(�%��v�ި����Y[%��m�<��R�X\&8	���D�ر�]�,BT�o@�~��)(��%Be/��0d\�N}��V����> ��D�F��(�H ��I	*�;�G�V���W�;�r'�;�A)>��eű��ﴩt�Q뫟�\?��G�H��5�U�S�?���R�������\�}�0~!pl��'�#UW2��&����3��O��w�QB�Ge��b�{�w����РR���Q$U䣆T��[����n*�>?)�.��럽@�yH}INx��]��]�Q��&"L}�5^0�rT�c-#4������]6�̹�T[�M�~����ϗ@�BR'�%B��#3~���z��h�(�ޓw+���5W�3�-D�|R�!%B�� �v(�I߂���|m�5��﹎e���K>
�?���A/&���!%]Q+�8	���;^� ��|AIP�R��Z�ʁ�}Q�A=N~��W���N�Xs#�yH}Z�%"HJdU�ߦ���_fO�� F��J��E����|��:�Gڣ�J'���u���M������p�H ��H!%B� �H!)�RSs��W+�卨;8p��z�|;_��̚ �9H��>IH�ʍ[�u��%]Y�~���*��
�O^Y�/��0"�Jhsή�~̽>"�Ig~�=9�lLŌ��ݺ�Aق%x�\������� �*�����^��ŅaP�� ..�݌ڍl.�vҙ�ԉ���(Y�6�HS �`����kf��W4��+�Yv)��Y0��8��H�kh[R�k�JSk0\H�)[.�����pKq�������as���F"���.������Ŭ��
�:`�H�aF3KB[���U�U).��)�YF��M�.Ɩ����%хq�cMA�U��~����`M�2�K�\�MF@�l�]Ivr�wZ�\$n�b�=������ߚ~����%��U_�{���&��8��C���ߝ���ktX��s��=�'{p�����#kۚ��������t(/����~���ӭj��A�H ���R�|z:S�����}�� ��H))�
R#���k;�G6�7jEGۑ�z�s4�|2��@9�4<�I	G��*R� ���E}�n�֢����^�ǰ�1.\�����U�a�\���� ��K����)��7��V)��H%AԦ�)H�BN �o鯮���#��v��ޗ��#�Z>� J��-}B�R� ��]�T|������rR�:���5T�kgU.Ku�]� G��t\�j�ں�+��Zܿ��HG>� ��$�� �)����>�-|̼_��W�5�0�S���z}� g�> $�P(�R�#.���Թ5�rk^����;�n��W�ōp����+G���)��LY���5���w���vV�Yo���ف^����칏� ��?x�$|{�V����ݙ�*��8��>}"JJ`T�j��4n���}�
nD��A���P0���IP�o~�}�j�p���\���#N��|�Ă��B�Q �(�U@�����5�A�"A�S�g>]%�t���_3/�+� �̚�mg�'�cޑ��]y(�A)D�
J��,�O���n�Ȝ�������*��8��y H}"JJh����\�q�����>|)��묦�	���F�i�SHj��*\���k5"0}��~뿽:�����	*ɓ�������'H}�>�P���	VR��?F��l���|�I	*�JP��`����什���B����N�&���z�_	�d� �R$����<��{�e
�݉�$�T(�H �� �]M�뜸�?f�y0*�=��A-#X�
�oA�T��-P�&֫a���׊ѓ����y����d��w|��*��-�=v.�X��
|iya�n�{��ق/Z~�&�]��n�{��z��X�Sv}�i�������{�/n雛���Q���2�w�=�_����.͐a�^wH^�k=���F�b>{J���s`EHS�ޅ�O��;'6�i~���;�`��&i�p�Q�2�,h3˫����={G�㛜��|=�\�R��y�'%ݯ!�e��Q`�\w��d��(�%���T�ytk�ܳ��XF���c=�w\������)�k�.A�}�B�{�t=���8�������^��v=�oDm��}�&��½�c�}����[�����,��D	�o`�}<�Acr @S��m���aѰ�ՑG�x�Y�I��׳
�v��WXkT3VH{UWk5=.$ԙ��Z��3Jڥ5܌�����]�)~�wyqӾ�� �K��8{͹5��2�ݹ�s�&�u��xb�-�`�޻x\7��{�S7N�Zj����cxG'���Z��HQ++j�Mc*��5�Rw�Mˊ*�U�5!w�N�u� �ߊ�_��qO{T'{u;hg�J燺E2��=B�q�l���^�v����zr ��|
��z�=�p�B����쫘�n3�C��[᧏z�ޝ�$�d]�{ͩ�����Y�xJ�O^Sˑ�Ɔ݈���87P+(���k[�{��1È���^�a=���m���w��uO��̿o_P)yt���37޷��ׇ��M2�"�R5JV����e�[��������N7.	�6�f;,�����{�ݔ�_����R�X�����=��[��v[`����ա_kw��N;C��{���)�6���gqs�<��o[��치�d~w�^u�7��e�]����.� �[���mdط̂��k�3�ie62����ی�;lڋ%��~_+��p�Ӓ6ڷ,K�l��#-��Z���|����Έ��h�v۴�2������[X�ͮ6�661ͷrq�k��l��v����|����/Lw��RU��QB�%;���e�?$�r��sz�=��{�\\?�����	 �H��� ��O�JD��sR��EVU|�͝#T	!�"|BJ�sd�w�|��ƓV~[�q$G˺��Txv��؟A�IUR�$�O�JO_@ߴ����¢��f�o\T�N)��+�'�y4<A�'�%3⒡�<�;�6}Ze��T�eZۢѫuCzoUtl�m�줭��P�珐�p�m	svbJ�����?/H��E(�A�J���/�����pw?P���3���;�� ��7��)BP$�����SC]�&3�Lp!�����t(/������ۍ�g���>4�@ ��
 ��5�qv�\H#mH��	 ��O�Jh����s�2�N��U�I�3�osQ����5�6��A�ɢ7��|RT+�(��C��ud�1��u���>)D�M�	�gʓˋ��w?z�9�$�|~�&��~������0�۰8���BL�v�>���P�h:����K��A��A��η��8��a�wnժ��h��MlF���fo%ʏO�
��㟜�3��-;۱{�ޑ;�,D������m{����rj�ۉ��q�q��^J=�)B�w��b��ꯢ��Η�C�s�B\���ش�V�.�T1]m��i՚��u�}����X��X���>JB{��g�M�\��6�67}�'d��L<�,G�"HnD���
)G��(�`+�;?"Wk���-D��{�o�����|_�	́ _H������?����$��'��BRW�> $�F}�}Q3��/V�Z���zs��|qĐB_P��H>J$��P���p ��y9�JD����������o�k��d�#cJ����[�dO�9uD�|
Q$$�QJ>�\U�\]��	�}��'9+���7���$���)H�E)�����U�\����ώ��qAw��\��d�e�2^��>�D֗�=:�x�k�b�B��,�7G4�N�XD��R�KwP?���ѵ�ߤ�w��S8E�SMqvth�b)a���l(�Lg��]��Iu�Y��F�V�@4m��u�#+��]":ӌ����A�9q�
S*��靣eآ��P�dM�j�v���\Y�ph����m(4�6����� �iuk���M��d�m�Fk�i����Y�1UL����l�W[T����&���&#!lv]����֚+�ר}��/�7S�jֲ˝Zd��#i�������Qًv��n��"M��@���0���O�JD����[���c>_z����q��	�0���~.4��� �BJ�R�$s�wP=]��:�� �����w}��c�St�߂��&�s�>%���z62+%y�P�� �q$$�QJ$�
PEV��������y�n�Nr/k���	��$>�%%5�JD���G#1�Y+>��l�!����C[�|���Sx%�n>�� ��S��ʎ�,q$�<���I	@�RS�z�>����+�z������N��mo�W�	y�@�p$���IP��9��<}������iz��,q�l9	lmv��¨�ul��#�4CU�=���!��WB���^)D�A���K�_	�n������9�7��7Dn���� �S�JD��� ���D}��ҝ��=)E���S{�g!�#5�~ĔkFg����lԸ�M2�(	�sB�k3mJ𯩓O�=1gT�uuZ��J���> ����7��R���_zRr_��� ���H[�y(�b����?B#�
��	JD��׈>JA�N�f(J���v�Mɕ*m�|%}>y�^ �r$��|RU��=b �U��$����(�%5}�|*����'/k�>�o H!�ڻ�(?�h�7�I	H�JJh���,b�������y]C���UJ�ғ���=�[���(�O����M>��`�=x} 9�iI1z��Af�v�5�e,����5�G]�BQ��$ɩ����} O��
J}IH����w<��LBSm��N�$)�hr9u�(޵��+�O�ޏHIP��O���U�'�����pÛ��(I�>y���w1���{>���9��
J{r��DD?q�7��� ����)JD���|���wV������=��CĽˀ��;����pK�C~q�
�=�N�H�6�LI�&"���
�8m��$�ڇʳuIV&&gF:��9�J��D�r_�������QJ$|R�!%@Pۯ��J�7������ ��H=�5������w{��I0���p������@��>O�bA#��ޡE(�	J$@IP�R���lq�V��?E��fp��B�m�.����^nW	��P&��A�]"JJk�%/�eW�I�~ܾI�b&��;��^�mi0�vN]�
�t�6���$v�!��y4A�H!)����
ߟ(�����9����|Aݫ�:��.��G��W�}%(�U@��	#�l��2�fM�*�8}��S@��#W�G;Y���J���?��$o&��HKOiG��YN��O��
~����	*�Q�(��~��q���&�;Y���������Wo����@���%J}��w3@;;y����ǧ��%B��U+�=��9����{�'�ufB�;�}Q�d9�3[c�7B��v���������A���
$Z�qS���Cv�[�2����r����y̤(�=if�}�غ�����D�O�$T+�@�)O�R��^|2�EI�Ѣ܉]�Y}}$��S���H&�MyȐBR'�%Bc��Uh�9�~��=�O���#5�gvbJ���6ci� .���y,ў�!.n�6����� ?�q_��a���R�,y�n��oɸ����Wo�>ώp�YX��t �Ȑw��!/�W�ng͹�F�P�Q��O㰶�Y�>)�
	>U�8����FF�����k�}B�-�}��X8�G�7(��7"AmϛrYD���L���W�H�#Sj~_O��hy�ngŷB�m��?LeB�o�%"�����[����>�N*���{#��"�����:���뭜�
7Knh�܊7�{���4�����}����\��������q ���nt�p~�����t�.L��xf9Q���1����tq��2/�m�]�¦�랷�W"�ԇ�̓�3��*ɀ�i��5��r��Y�B~�Z/�����YG��{	�D!�e����\���H�ar-��BY��Q�J�]Ast��Y���F�q�����ٸ���W��7�MZU6�L`U�
��
��.�m�-��0�v�%6Ti5��Z^כF-��a���������V`Q�ք�fE�Yb�PK-��%	u�<��Sg[%݂�*WW�K��3��{)]m-��P�m��U��D��h�_S�=�/}��0�U��c\J�]4�H�T�K+D�p�:�]��Wf��ޟ�~~��~������y�B���=y}��RmO�k���Iz�����@}�����mТۚ ��I��������Y_o���� '����}�ړ��ݯ�V��N@��$��̉sgB�@_`�Am�[t+�73���߶!�$�M����Ӻ����ɍA�-Ͼ:�Hk�ɹ�%��uA�~���H�}�Nx�۠��]g<�D�E�����A��ɠC���a�;�,�q��}B�n}@��r(����rs���^S�����I��;���
�"�ϤO�nk��ۡ�Qd{���z�1�`��l5ıSZ`�j`Z����]�cs[�u �|���>����ߨ���6�P�N��]־�����������QҺcA��P�{����H!�B�ۑD0�`kq��_�C�ٝ�<��x�xx��=�D�I�ٸY�+�Ub!�;-����Eb/��[v���EW�}���]����.nh(�|�!}�+��1:��d	T�iG�k��� ��B��n��þ��ʅ��@�yĐCn��� ����OY����o�����F�z�Y��k�P!t	�>�۠�H��Z�/�f�FT����>m�R���U��~��u���%(�-y��#����t�1�S�>��t+͹�m��5|v���V�;����O���Q�k�H'�&�|�������S�oF_�Tt���BҚ������6���e�6�6P�j:d��&�rU�L�������8�!��������oE������o������ETW�w_b���\?7>�$�P!@�$��]����l�9���Pu�����ݟ�\JE���� ������������g�����yD���(��Ex����8-��۟�Ѫt�-�\u��u_\Εr��9�Ҁ�{�=���;i]�iW�}�s�V�ZO��&`�� ��d�}�V����IG�k�H �d��^!��ۡ@��ڥ�����]��(nk��Bk�/����4oV_ë>�ⳤQ���{��eﯺP#��W�nD��[sD�
!��[�����*�*����N�F�$_ʜ����!��6�||�p����ט�晹0A��jE!IY
E� ��%�Ƥa,�k�f�6��06rjg�����"�?t��m�Cn�G϶]S}�@�V1�?	߄�<�$�1��ݿ)���Т>��܊�4|�y��������X���}@��>_�>�߶m|��ڿ�NH��gH�D�[s��i��~ۡ^#>�H%}��� �O�mЋ��1��/�꺭KO*�4�*s� ��<�H��� ��A����4�����}�R> ��>?.���B����uM��qV�|'~�O^O�u�*y�?�hD	���m��!�Dm\�_n!��_!�gn�$O�\��Ŵ������}��ҽpSUۣP"\I1B��M�ȹχ�=:��@��%���
-�y�g�2���������u�l�_:ۥ��
k�Q���9�mЭ�}������DH�]��7If�
3dh��Ġ���i�jS9`�5LA����A�s@�>]@7��t?���K>*�5�>���DX�큣0�y��}}����sD�A:�n@�f�1�3�{��6�ׁ���:�u-u�V��p��A=�5�s�D7�:s�~ܿ/\}�
+� ��I6�P-��A-Ò��5'�+�}��ͻߵVj�˕����7� s���5�CnE�}�?WH6�'eG��
/��۠��T�ڳ�򸳖S�N~ �uG�{����l:�_�jk��7>~=�I�[r(���H)��?�;q2�̜��������D����++J�N} �}��΅�zCn����}hi�(GC��'	_T��7_��u�X�k�@��=�L�֦�ͦ�x�\�o[��tc�`xV�s��|f��e��]ξ�ǉ��L ���^�|ظ���,S�.��(��=��%��eKKfVm=�x�D�\i�wX�״y��^�i��5���-��g/���ݜ���c~�P�/��׸a
Lj������4{��*pz�qQ���w��;�����٧�kYy<)�7�M�����ŭ��g�-�z̽@򉨊{sE#y����H�����ZQ����W�p��.C$�v㫷{z�v��XC�z������|�r�`ٰQ�G�{s�L�3m�G�8d+Տq�f-��Ŭ(���*�N��s�Lξ�8�*ᱮ"SmIõ��%�5�v�j���ʹ�D9�X���N������a�@�Ѷ/��`✵�|Ji�Y�A�1�c���|;������:�=�Q��ԋ���Cp���5P��&C��8Yٞ>|��}�w9�{�g[�(U��;Y���q�`��T)�,����4��ۼ�}�gE�n��Ѹ����t���J���5��Om�H!.5�º��z�H���hsi���_HrWo�.=�<r�j�)��ξ7�}�#��.���\��{7���T<����|���}�����7y��*��/u:�a���<r_l,��f�@p��^�t��s|�;�mH�V�$ZMն	c���ZU~o�a�t�{��!���*�DH��
��ED*r��+�ޓ�ﲩov����/=&7��!Nh���3"V��^%��M�������S���/B�:ܐ	��%%�+:G2�̞��f���kI���o/{hu'����Y�ڶ�jm�v���y>�ry���[y�K�{M�� m��{���_@죹Ώ0��������Y��;۰�ؗ�<����T�IBC�VX�B3Y�d�:"��"w�^b�[F�6h�{z�+��rpp���Z��쵶Nu�{c�ҏ����2˓�r�������ۭq�޷����F�a���_k�݄��e�f�m�4��{֙��� ��PIו�|�9 �!��1��_n�;�_{^�RRm��q�ٚD(G�V��m��.�3v֡Ѷ�)K�i�m�� �l�@�IKk�&������H�C=�Iq��aґ����ֳ7��Z��jEm�QX�
��<@�M����n�/i���]i�9RŃoU����0�skTݴ�\4c��yw�<a���
��M�#�pI�l4]khJh� ms4̤dĹeѴf��(�Vc���TR�\��	q]0&\,�ı��1�3L�+�p9������ÒL�	���4���E�m�񳹣�J��l��i]��30�hZ�Xjk��n��&
1�F�ۜ�̣�3Z�ց�����X��k���-�����E��n�p���[k�v�T�fiHD��m��`�� Ffp�mf������R6�yXۣ6q�B� i���k%���(]��4K#��M�q�4�!1�֧-�4�M�#T\TF��Y[����B�b�+�AR���z��F\M�n����u�,�d��=�v1P!y�2�V��[ԅJ���[� V����[�5m�se�����0Õ�v��Yb�D[ѭ��L�F�[�B!��e�r8P�7a��C[��KH�x��U�1�ė:4�bR�ժڱ�\grĆ�J7R�1d&�*���gM.&u�أ(��^F�Ԯс6�(k���hSj0�=b��t��=e3�p��J�g8��ј@�HkZ�����)i�q��Z��z�A��*@��T�И���H�B��b��-j,�����mH�MHR�֑�eJu�aL۲r%60�p���U��il�n���V��&��u �T������Q�d &�(]V�0�c���a��i�v5��cm�c��W�R�V���[���,%��9��f!F�bl]�SA�VmB�͊kCipS�p�n#��d��4tԹ�tB�a��"�ҩs����\q[�Y�0�%�YF���%���.��+�M��&�1.��L��؆��sL&�����a�&�t�M�mƍ�$�p�]a�e���tft���F��ì.a\��V��c�9t�0k�#nţ��6�����(J�.Fۖ�9	H]���ٹԖt�XM�!���e.��-Q�ַSdr5�ا\Y�@�d�f��C)�������\˦�̈́e퉩#�BjR�lp�:�;:dbi�)�E��#���Z�+�K�i\Rb��n5%,������5��Y�u���lFChbh�I�2�5�yȍ�k�\�%�e���h�_���g�6���⭏-Bū.��q��eDGF��g��_79�s+0ګ�����������׈%��<{���~�;Z�Ʌ���
o�MB��߻g�@��$����
!��Am�a�Ϧ�s5�u��#���t)[TƯ��������5��qD�F��E�=��R�=��0���
nh|ۡt%^Ӿ�#kz��U冕p����ɠA��@7�u���R='%>F�}B�-t׈%��i�'ٙ�����L;�t� ���
_۟!0��5����QȐKnh|ۡ@��.�o����ޱ��
�u�b�[�Ũ�z��s��b|A�]B�m�An���7�G� �;�R"	�f��GQi�҉f���X��D�,5#1�b	3Q53��C�H�>-���
��-��_B��*�e}"���__N,�_�9��О�r�33F����#�X����T�/��+�z{DwiUu�{K�B�m'j�$��a8zV��Æ-Y��[UQu�=���t�	����a��NWW�k������q���}���D[�������)����w�鿨�H�nD����ɹ��12"�	74!�B�nG�͹5����;�弝�z�7r�����?A���P�۟P-Ǜr#m`��C�S� 1�"N�5�mС�O��]ƾ�Y�W���fMQc;)�WY��|	���}B�n}^-Ăr(�����[�����ٙ�S+~q��Ӓ>��� 7"Am��t"OƷ���������a�>O�v`-v��
��X&tY�n��.
l�nPfȕ����g��hC߿�� |��o��!:qՑ���J෽���>����&��~��7���� �Cn�܊�#���*W��������Mx��P����-���e冖|' |{2k����Q��Q߳�!%k�z��r����6�͹���S_mjoG�r����'��M�p4�kr��1
�k����t}NaFOwl���JWt^�-�w!��"��mj�0f��V��ڔ������2���ӳ�#�Aȟ��6�P!�����k��S�_P�C�g�ͺ�Z��|s-\8{�c��}j$��u�������MAG�y@���W�-ϛs��~��W�!C+����/���t�04��s��d� �΅x���ۡI�[k��"�1�
kú��qb���b�*�k+-snv� �$�K�A3U&KR��}�C�E�4A��OWϳ2�S4㿇N�(W�ufWM>?o�~s�!�~���#ͺ��O�sD�O�&��lzW�Pn�OcY]���P��Ft�&�H ��P�ۙ�#~ʯ��P�W��}�}!�Ȓۚ �ۡW��V��I��y��v��K���ד@��΅�Kn���\�:�quy�N���}z�s�̿�F|�ͻ�v�7�"�G��v)��_�F���1����-�2���V#/뷥����ְ��5��{���I��Y�5�J�d9��J"��xrdL�EM|>-�4A�P��%�>m��D�޺�r�E�
/�����/)9��Ft���I�P�۟W�q];x�>�b�U5c��J�����1c5xuv΍ƺ�/*3v���ʧ��H�t��4A����)����e�i|#>�J���Ơmmk�7���Ϗ�t(�� ��H ���Ҩ'�g�fϫǺ$^�\粳�+>p��ԏ����� ��3�| Ƒtz��ה+�vH�|�� ��B�n=-�뭭�����М�=�ᗔ��ߣ:~��Đ_�^m΂-��۪�oa�����9��n}�mС�﨧���Z��6��F|${4E�Nn q����n>>��ۚ ��|CnEx��.����M������Ϯ����+�=��@�y�(@nD�۟Sn�h��*(M2dԣ�c�	�*��H��@��K*At!��˨a�����AG��,�O�V�AWw�h��j�?uP�'�<�|���f��C4�S5X�-�G�
�.S�Ü6����c<!	��mq�*m��Ů4��5(щ-B�j6JD�-���P�;4�-p�K�@ʤ�0J�]]H��#��Il۶�U�у���cK��L��%5J�fғ���t��E���uCLñ�iWdAɒ��W��m�.�*�l$���m��F�jZ[�%���}�|��[�4�#(.%��qV�l���;$n[�1�.�k�n���5u�/���>n~{�@7��6�5.O����������O����EF;����Χ�^ ��P��}E��O=@�ۑD}�d����_�@��C�u�~޵vm��3� ��4>t(������e�~3j�{4 q$�
-�����ã�2�Wlnͽ��ݺ�|�ޠM�(�Im�ۑ^!���Wͽ��3�@n=��T1�ձ�®q�w�7����c�k�kb9���w�h��!�T-���ۘK��ز��~�<>푱�f��{z�U��k�d�U��@|�����_8�.{����:8�5$�W�$H�������j!1�5�hmq1�y��7�
�V[0ګ����@���}�(���֣���ٌ�L:U��H�j,\���8nH��H�R�n�܉�nh���O���E�)�����ˁ
̋�^��t6#{f�4��sN
�Uc%d�`r�Mź.=��7�Vʹ}ﮡ�@��ڼ�dU̓�">9�����'���z���۟� �Ă}�
�1�7�nW�$�y=�P ��E@nD��׈!�B(w7V��L�Y��C+���;Ww)����AZ� �:nD���P-��*�a{Y�GwP��4>��mj<�}�?V�a⯃��
�r+�^|w~�Hp1��c����>��Q��۟6��{T�����٪�fӓ�!��n�S��m��ױ$w�H�nh�p��ﮭ��֠�a���v�KD�(Z2�l�6�L䄺ֆ᥮��-t��j^0���o�|�ﯺG��1����ۡB9��Lp�~�{w6��N@ϯ����^/���Ak�Q�O�mכs����Ir��suTN^�ښ>N'����c��L<U�{_z�6�@��H�$9_Bod�T���$��-���6�D�&�����ٸ���o��:w"#\O�y�%Sl�v������Q8��}�=Nq�e&I�r�#9�o�J,Zjj��UB8���2��Ӛ��Q��)�cLt�:ߧ��	��� ����ې�6�}����XV�H�-�����
O�2>_A���M|&��JY5�����~�u��ψ���׈>��|t+ŷ:�U��]X��CO8��Z����6>ĩ���w���H�Cp$��-�}�V^�Q�wGk��^�K<�;�5�X�!wU�iq	�6�LSB*�Ԥvun�����hEj'����=���C���X�܉�mЦ���/>�S��qϹ��������� ��s�܍"�2R����śܟ.���p��w]��P>;jh}��W�nK�b�1ҽY]B��SD{��ۡ@����;�I�"�}7Y��7��KY
�k�+ם"�'"Am�n��"u|�J��������h���@?�|[t(5LN�}�m�ӝ�q����������.l&g�
���F4n��yi����[�=V����%����� �D�c���y�"=H>�%a�����nv��ٻ���}�u��	_G�r0܊7mΏ�;��<����T��6�����9v��e@��4A΀O'͹�p����g0켘'�SS0f	� 5�X���A�::�â�����r�Φ>�ާ�}�$C}B�[sG���[�����1d;P������p��V����@{�$�t��ۡ@�� �����FG���>q���r�X]�?���)��㟈>7��ﾯ6��k��XEx�h#7�Q��
nD�ۚ!�#�lwƔ`0�V��깝�w���m����A;nh{�
7"|[t+ŷ4E=�;��B���_P���@���k~����|�U�[
�k��t�/�f�ʯ.�LO�O�w�P����͹lW<���I�[ϼE��
̾�1]���4�N3�N9�|oc���
�5������M���U�Ⱥ�ؒ�bş`�X"w�\<$�ugu�(��	�cM�2ц����:nWe��cWUa��݊�&d��	LT�f�5��+�&ABF�S�tZ�R&���weh�I���P%l�WJ;4�+ZG5B���
��LhcF�𡄻h�*M�%j.�fQ	��D��G�Y��mns��f�����t۲�s�aSPى�De�:�ښX6bժ�&��¶�˵�;a��y[ncT���SA��&h��Հ.�"]����n�F2�[�G`RZ'TY��6v�}�I����M��e�5��4VŁb�h��9as.���+�S~�{��>~i�A�%�4 6�W���î�}v����Fڏ��|�}� �n��D��"�[sD[� ��=��y�{��%t<{�|]��W����~7�"� 7>m̹���U��66@��H%>� ��B�n=!�B�OϾ���
H���M}���o'ϧ���ؐA����� ��H6�\�߷�����>ݑ'~sD�>�p�|�bbvq�	���#���W�	1W������dO���Ss^>n=>mТۓ��l��Eg]Є4�>�����߾hj�X¿���P&�P ��[s�mЏx{����C��p�`��+
<TXAT���^�,�h��ؖZJ��z��}wY~H��O�R+UX����Ҹ�7ң�hN"L�H�;���*��� �[�!�B��mȠD��\b���_#g�3V�>�jŜt�Y*�&�4^�X�O�-x5ׯ�)����o,����m*��������[2��)e��ݧ��*7�>/�h��Sm�u���5w�E@��9�A�
!�@�9��{>J���4��'�t(�׈%���Ǣ/�3�~_gԗF���Jq���#�y�(Cr$��6�Q̈�?d��j�n�ﾛ���@��=!�B�5��3K�q�i�����-��ꊯ��U6�X��}4}�!�^�|[r(�� ���F���C�dk}h}���UB6���\��O�st+�73�t7�hu�6E�������)��Q��s��[��#e�t��S���Z�+pm��������h[s@����wݽ?46uN����>��|[�cT�H�A�9{���#@!�nh��� ��+3wF�����>����	����TE���4��xډ!��͹�k3����a��$v�)�!�n|ۑ~���U�ْ1剃�Ed��o6U�Y�7j	���1�nۋ"n<|W�Ύu�Uwvmݧ�R>���U듳9���Y=ťz|p��-�ob��7�U��y�&Ao��M���D�І�����3nk|��0�=��f�\��F�������-�<yd��U�p{ٽ��J�ȍ�'d��^��nS�i;���nMx�_=m�娗���h�c�V�"�3��o�A=-[9�5�e�Ɔ��֕���r�7j��������K�;��,��x�p��3F�ui���5�G�m���h��iކ�_����K��n�E��'�(E^w��}��ǜ�'��W�
i��ѹ��0�,��x����wM>-%B�T(�ԙ�~#��&�_v(�>;���qu�,|8����Z�Ό�ҝ~�L�߳�$F��%��"%^䷏�����]�q3�>�Zs����L��Dwu�'}�M3�n�md�S92�.�q�1U95��}�ެ[�2^������<�r^�5����vJ��iX����.���n���I���oD����.L߬�r�.LL0uQ��ql�4}�I2#&]bj���j�����*�5b���q���.{��t���7rX�ْv��D�7�'yB��p���������\鞓���E��JI~�^\�U��#�^�\���x��}9��[ǌ�m��uH��
��=�cK��r���	�ƪ7,C<s�����0͝|1�f�OM���r���f.^��xm<c=y��©X�������,L`�w76���l�����f�V��݌�BR����e��n'/����k��	��)\��_�s�ݛ~����l�nt� ^�n�����ü�"�;���N5���{i���y^�	�1{[�������"	9' ���P{w���;�:'/;
|�~Yy��p�f{�����)B@��{����4��;o+��z�'�o�ڲ$�߽�~w�aģ�F_�\�ט���`�ߞ��n��fڐ�8��޿}��k98���:)�mN
!hI�[3�mR8V���q�m����n���N�X�q�i'|�ҀJ��m!O�������L�m��s�\���6�����XGm��v��NR�����N�.\�''�m��K����Y֝��n��+{Vq϶@"\�R9!~�$�@$�]��3U55�U��#~�|o:h�nEx��͹�ۚG�.���d�5uG��΅��-Ą�{���_-��Z�߃��U��P7H��S�y���_J �_P��%�4!�B��w]L�C	{t��iЭ]xb������w�3�?M��Ao�Zs^ �[����i��T����=��|���9[1�
�k���[���Mh��+��V�b��e�=0���z<B{�n|ې���l���MlUk|#~��m}�I������W��>��
�m�An<�ϑ��<�& +�(��}G���߻��[��Q�=�vT����Ds� ��z�aS��e$Ɓ��G�@�A\��ۡD7�����J˸���K~�ɡO�K��AY����[sG�Ăt	�-��{w2 �"N�4!�B�|w8w��յ5��#`}�}��Z4���^��G�����I ������1��}���9���ӽW�Bˊ�j8z6���Ê{f,�� f��˴^�|>f����y�>��Hۡ@ܙlfyQ+�Q�jz�����dhY�<�r��z���r'ŷ>m�����{�ׯϣ	�?9�ʚ�f��)��]�ܝF.�m])5�H�r ͚�Y��~�o����{�=������ۡ@$�W[�~����>���p,�ɻ�t�"�A��:��:>-Ău@���P#>�"���4~�����}B�_(��;�*~����zA �t׈#��@����߮�{���{�� �q$6�P-��A �\��WT����}��=9����J�P&�d�0���t(��F,}�k�>� �t(���>#ͺ��1�}_|f[S�K�n> Ⱦq�3��}tr~����H6�z� ��P�7>m�O�
�o�L���Я%�������ѱ:��#���t��'B�Cs>mȟ�yɟ�aШ���uPa�H4�ļ��1��[�^�w{:PQ<�KfL���i[�F����p�Q��1�ۀ��gc�w=�d����v��$���]�A��.����%�W�[Y�1�$����p2m(�I�s�Z۲1��0���3�v	n&�23"�,	��ę�k4���{bk�`\MT�X���S:�mNS)uy2�.���26Xj��T��lB�b����0�K���5st%q�&�X\!ls����R�YxÌ��**X
�3/R8e�a1�:�lg+����_�5Kk[K���#��Ò2�^�W%C1�T�
A��L��EL?s����zC�6�H%���{��/��Z�߇J���܅�ge���>�D��s@�ۡ^!9�Knh�s�>WtUk��>>��P�� �_�_|dEZs�S��[�Ho��n{����Z�Iy\w�\���E[�%�4mȚ��G������y3�kUB���|$o:hy:��y�B�[sDF��������������<߾���9�ְ��J��	��D����b�XЛc *�h}�Т� �ۚ �� ت�=N���]������ݵ�Ƅ]�9�<�����o�[s��n3y(�sk���bv�X��4a�i2�b������pԙ��j�Rjj}F8)�(ΑD�H�[s@�t(=/��]�5���>�t����:w>��O~}B�����[s@�[�Gfk�mq�3���-τqqՃ��y̩D��D��k.�z$����9�X��i�u�,�\���%ˋͨ^lɒ�sz�q��獇���.��of� ��O7�m�߆赬=�t����A�t��.lb���wl�u@7�����n�x��|Cn��~��a�ʫ����wi3b�۬��O������^-��A�n$uB��^�7����l�>�$���B��]��k��U�:������#yt�12u�@e���
-���n��勇Ճ{H�C�H\�|���_�kX{�r��^�;�O�m�n�Ws�����~S�]6��nc��H%-UEspX[�5�]4�ѥp����T�6]��ҳ��:���D��Ѥ̏HmС����?���ػ��>���'���B�����.��M-����P>-�EW8�A3���@7�5�7B�ev�ut�#�U�8���ސM��РC{�����2�/�їt(�}@��6�P-��A-�����u?!Dd��D�`z����WU�����vk)B�#����R�<>��qx<�%�'��F밍�IW�2l��R�۽�UR�+b�V�Vٽ�o^�eh��{�ʟVd���%�4A��Cr$s�E����ӏ���Ӥ�B��'͹5���S���j��{?/"H}�q��D�ښ����,�
q��
��Q��nO�w��m��H���*}]?��N�'���A��7��7"||ۡrQ���g����?��=��5�,.wf����2iaVP�ܗ&����GLgl}�����/������
�5�	N%5�~�{䜭ڇ�+�Cw����G���D�Nk��n�x��|ۚ-kk_�r��� FtzC�B��q��>���U.}Og�	�A��W�nht��f}�n�>5q>!�T���@Cr'ŷ4A�}�k�+߱���N���J�g��U���9:Cs>mȠ[s@��������Ty��@�sD�B{�_}��[��[�{�s�P&�dQ�r�T~�ɣj;{��ùiX�^�o
���f��[Q�e�{�u<�fNW㩮���KnzOj
��R��TC��To"�B���E��ϲ|��B�!�A�4A�mТ�x�!��3F�^y�_enD��ί�1U[>��� �q$�������=}.����`@;Ȼi�3s�cUZae�2Ya�΅�] ������1��̍/��K�H-��n�e�����OR����5��.*vs�
�S��A���+�/�||ۡ^-��	n<��Hq}׽�����M|~������붵�wO~������ۗ�C�l�L��5L�[s^ ��Qǥ�Cq,�2��˦c\\��)󉩬��S��[� ��
�4|�I�2u!�W=��~�r2v��;��ﾚ �ۡ^l��R���*2������k\������̟�q?���>?.�E�5�	n'��t(��Q�K-���8�D��M����om�;�߃��W�vE A�ImϨ6�1��?�i�VI�� rѯ/�LW��)�,�E�Av���;r�I[�v΋Z�4;z����`��׌m��5��G}/����9q�ܮ�7~@�'j��j�j�02�l�[�"7��x����cO���W`�T�n"�!l���n�-�ɫ(f츖6�UeɍZ����x��C[M)ti��f�݁�͘%�]r`o�j�r�j�	6\�b�a��\n��&�l�uJQ�1�J���9��.�m���uтG3`�� �Kk-�����l�ybO�:S��n�s���3��=�t��h6�Ƶ��6�.�E=f�G��)s�$��ɫhK�p��QF��{��^�4)�
7�6�k�e�Y����Md<��V�c��5��+�WMx�n<��P>-���rT�*Θ�cs�Y�ɠ!wP��_u)}	��K_£�Z� �t(���R�fH�}�D�-��nt@-�����=�nc�X�7���˺���~�7�"�A�ImϨ6�Q��c�w�쮋_t�� ��P#�O�t(k��]Go}7SY>����^G���]K�cu|ٻ����_{~�@�]Cn�͹-ϛs�|"�xL�9B�~�Y����:��u?+1�_�b=8��99Cs>!�B+jR���>Ջ_��e��.��KJ:��\��3D�,b�f�ZvG )[����Ye��z�>�u
�m�-Ą��v]o|Җn�7�ӿ
m���[�j�H�
�D���A�n�nۚC�tu�Cbk$P��;��⇁�1��d��&t�v����Z�E���5�Î5B�p��R:�����pw_.]}B���ܻ"|W�P�t����{ꛚ�Y�r�|yA�_P�۝��E������>�U��Er$���A}¥�"�%����d�n�	��B5c�L} ��5�� �{t(��[����ǹo&=�]���;�	n%=��]�[��*f�~;��@�K�<�ݧ��wT]�X\w�^��}B�Cp$���B�Ch������;�^�;g鿧��c+)g��~ ��$�����%�A�����I��M�Dl�9�Xܤ-v*[sj��;D0[������SiՔ֛����Џ�{f�C>��̽��
�L������Ӣ5c�L}��W�Q5$9ܟ��A��(��>!�^m΀A��&��b>���{�QZ��8����v]��=T����:vG�7� R�nJ���b0P�@���	mϛr4��|Cn�-K��3$v��9M����r�
�g�什�^������@Ƹ�_��s��f��̈́��~�Nz����8_M}�<1�ه�H+ăe{�S����zRϫ��>+"H-}B�n}E��CnCɌ���dU�JrF��]4Am�O�>K;�1}:#i�zA5�h�u��Mg�q9���}�>>]�
 ���q$�y�W�g_�9aܺ������������/��Vd��.� ��6�n�[��=�l��z��ﾢ�F�Y�RmlѰ.��Bd�]jM�+�"���a-c�m�^�l��=o}����$#�tx���
ݱ*��_Q�x�>�S�!�O�s~��"�P�Ϧ�Ÿ�Cn�@�ۑ^#$�l��(�:���k�ӡI�a�y�Q��h���	޹�{��^!��>�>�;�.G�����=!�B�nh�[��ysvv�?�>��k���M^�ö�|��@������nD�w�{�Kje�[�vz|ۑ���V�?�D�[y��?AY������O�Q!�Z��ʁ�ף�_�gR��X&��4�R�߭�Z�4T��j�w�7:�FG�	��Aq�37#k:��jr�����e/�۪ŷ"��[rf�����G�*�s���Q��S���mM��P!����
�������6�Q�1Rj UDT�GmG4����:�.��[{.Fg��;��v�0�X�;c�?zM�{��nk��kޏ���?O4�M^�����;���w�P[��#�A�%wMCn��	�4��9��gd.�>>��W��c�����ok>���JȒ��Qm�J_Q�+]?wFג(NE[�%�5�m��&~��4f^[��Gъc�D|$�4A�
7"|ۑ@�戟��쯫��+�}�in$k�������W&kw��_W�l�"�s1�u�^;�4#�P���A#�����4&g!��?o�]}]����;��W_W+����^Ox��I�$=�oPE�k�BI�PBO��$�� �!$�!	'�@�!$�BO� �!$�`�$��@�!$�BI�BO� �!$�BIPBO! �$�B�@!I?�!	'� �!$�BO�BI� B�t�BI��(+$�k*6�@��
B �������������8V���C �J
   %4&���z@6���   �S��iIPɦ@h4hd @s �	������`���`4�*h%@z�� �@ 0	����L&i��$�A�M14I�4z�M�Q�I���V@((�sU �~�hGDGZ�����T�����������~xa����q@T��i\F� �"2	�T@��j�an��۫���* eCo;6�M����G��<���E@�7�F��J�N�]T�X�?���Й1/#��yw!�+s2���Ɍ���M�DVQv����MKwqX&5AT7�Ja���i�L�wE!p���Z4إr�H�9Hbf��sX��w�&�4��|A�������sik9 �*��K(���A<"�H
�w���s�i��t��5ς /�KjHi{iqAM��ȁҙ�;�q<�g�ʨ?A��X��i26�`��7�F"���B{L���PM�O��h�Ҳ ڂ�m�≎�=�ڡ;"��U^W[��UP+�� �x�Y�f �$�!a�&"UMVL��D/ۮ�	,;n�؄(UD;,e�@<��Uv�]+nQ;*n��@5K"�J+jV�+uZ�
�*�Z �)eʛ�p���"�%�d66���l��3*`��I����!K�E�����rʥqҹkUUl�-�Z7:���{����'\�"���&\���]]�6���6���H��`���fM�w�YkL�]@5
a��&��;��VH��I"���u\ý�e�a6����\�5=.�bv��1:6���FA��a����+n(�9C޳4��x���V�P�=q�ۥq�2�V�L0���3;��|���2/Z9�9����Uq�V1"껜�� �[�<��bjl�UO���	,G
��u�W��+�c�}oc��$-sՎ�]e�uZJ'aId�&^�.Q�^�����۞֧��P�I�R���ش�/3��o3����r&��29gyH�>(N6)�%�\�V8� «^0�I�m;1�U�M�[��
K���Z�If�}L�y����c��v�]�2C,sEVe'��bSZaf�i@:l%��춂H$�H$�H0�2	"��H��ժ�I�I�I�I�I��R�R�-R\@n��.LŠ�ӗO�L�n͜�Hݥ
�� �鬀3�}����!ݡV��f)��+��'�W�i�].jKw���������e����TV���Z혶.>X��<��L��mr8�����̀��$��P�iM���al"�	Qz̴/�24�{�U�JI��FUfEToU.�#������������"<G������)��eM�K(|�9ŷ���1�=H���J�R�����K�����22;�D�v�s҇:/0�6&���:ߍq��Ia��&�iB7CI8.(&�|ã"�^��;�����'����'.D��x	��qL�@Q�]�E빉Y�%LH���h�\�����DׯI{j���tk�Sm�UJ0�g��k��P�|���9Xwg���� �ZZ�'���ً�{� 4�i&N�u���=��T� �L��Q�rv�{93��S���I�8炷�h��9�Y��9\��ܖ$�E�Ch( �i�N��Ä ��%�a���ʤ���QX؁=�e��s ��p(������b�6�P�%l�G,�}�v��h���A��F�qTf�r��S���zn��[E)Wڡ�&V ����P�"h�|�f�T�JD�Y*��lT���f�$�X�">)Uˌ{�\Ŕ�rD�1��nwۭl�Jq_�{k�xR��(�� �)T�iG?����S���
=P�7�;�g����X���쓾LQ;Ajv3 ������pBrP��, ��ʝ���l���-k����P���&�M&�p��u�Xpm��G֭�^�p%�+&�v�c?�U����%a��ve����_'�T �SW���f]��  d=� �A��(Ȕ�9��ý8�q��|����g��:��yw�k�Q����J���� ���f6�cb/sF?���.�D�{Ak��Uv�#}���i�^��Cxi�O���h�� Z��	իv�ؐ� ��Xh��"�b4X�v�Qj��z��8M��遬�T ��0k��zoo��a��>�pJ�u9��쁬L46�W��0�{ϸh���-2�q�����@���Yw��6�؟������L(�aю���h
r�ʻ��������M�p?�јx��;�}ܼ�{���(���#3���2?O3e�<۹ؐ�)F�S��]���r�����s�N�*R��5X=̋�k.>����贒��6&�	�3�$TE�Cs"����~��jI��T)!�2��,�8���J��"�0��A� �h�;x�ǆ��N"�C�F	:�8��?���5o6�5�t��'>\fϑ�&�z��{�Ȟi�!�7%�\6�P�I���|ރ'�U�?o�3I� ���c�����=M7�?��ݩ:c�C�۩1�dGl�y��X!�i�\������נ_`hG������gc'MA����m� 9u�K���.<R[mv`b����(�F���jza���2�Ƹf\0�ܗ�Xn�E݂�7 𞏳��r�׵D�x�� bl�:��qovb��D/����b�HHPC�P���#�{���ܑN$���