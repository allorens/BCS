BZh91AY&SY�GI��߀@q����� ����b<~�    ���VڀRJP 5�jдʩ�Z�ѥ(6j�(Q�J�m��m���%UE*ZR����٩"UJ�%RKMSAf�i�ڷ�޽�F�������H֒�Lm�mm���mccml6�U�m������C#Z�Zf��ʶb̪�![,6�J�J�d�G��jL����%m�l����֚�3kV�#Y$�km4������T���m�k5�Ԗl�UV$�&��[[3�ŵ��U�1�`[V���y�6ű+@�  �>�U(�]n�WMr흷�+v[.ѱ�c
�J�����(��6c�F���֫����jcq�PS���e��kT�-[@[PV�x  ��M>��o{�ƔL����P]��p� 9��%@+ҙ��PR�v�� )��M���z�+@h ���� �8n��216��fֶXcc+�  Y<( �X} A��p: c:p� ;H�
T�p:���CJ 78�ǡT[�`�w�=@w]������h-&l�m$V[T�m4>  fy�G�׃� _{�q|�>�����:
�V���(�u��t� z�\���l7���C�T�-�h4\h�(_e4{�ͩ��Y5MHd֙2P־  %�l �=�s@ s��} �ynС{m=���A�� ���[=�ހJu�sW4�顦��8PcM��e
�K2�l����� c����N�8� s��p� �ӝ==
=^� t�q�{�=����pJ wKt  黣����ݱ��PwI,X�4��M���i�| ,W��  ����A�@�LС�8��� ��0n�m��ǎ �0�� ��� �*�Z 3�q����֬El���ͩ�m�6� �  6�n _oz��d` bj
 mF Pgn(��׻oU� �b� �v�T�V��[[mMfA��V� � ��@׶pu�YK  s�p nup ����l�p)��� s� vN���iVZ�2U�j6�Ux  < �!� �UX� ;� (�� ������ �  ;�8 �B��   �  S eJUF` hi�� �{F��%J�&�    E?!)UM  i� ��R���      ��M5U�@     I� =T$���z�&jb�'�h4�	�����'��|���o�l�|3��)���v��ub��?������}�>�����U[m�umU��j������U��ѿ����m�u{V���/�������_��U[l��p���U[m�W�6����k[o��?����������e[�����V�f׬��W�W땯��י�y��3_9���W��y��lڼ̵ͫy�W��y��2��7�V�+^f��k^�Z�5�2��6�3Z�-���f��Z�̭ͫy���ڼ�k̶�ͫ���ͼͫ�ּ�j�6�3U�Z�sU�Uy��3^�k̭y�W�j�6�3j�6�2��̵ͫy�]��5^e���y��3U�[^eV��[m}e������Y�k��o���}e�[�5U��[V�*����o2�V�-������UY����Uo2յ�mU�Ͷ��+U�ʪ�f���m�o2�V�6���Zf���Umy���3[Z�6��2�m�Z���V�̶��e��*���Z�eV��V��-ko2���UV�6��f�my�_9�my�ַ��ky��[�6�o2���6��̵�y��W�k[̭�y�j�f�[y�Z��Z�y����Vּ�[k̫[��W����5[^fյ�kk^fּ�W���5_yU�m^f۳o2��j�ͫ�ּ�k�ڼ�k̶����k2�3U�V�ͫ�ּ�W�Z�+^ek�ּʼ�Lڼͫ�̵ּͫy�^f�̵y��3j�<ʦm^ek̭y�W�my�y�h��#�ux}�~}6�v���~��j���B&�4T�$9�������s"�z��aM�^��rX�h7r�$2Af�zү�U�!��kAbC�y�r�90�8�d;�Ⓐ���
bŷnU���;{M,J1�;s`;nnhd��h�iCv�����.�QM,V)���uup2��B臘������Y�j�9���D)������E٫Y��Y!x��&���-�X9c�wz��L���lnv�F�{]q�A���z���Z��[�u�1,6鿦[�9W(,�c�y/Z�b�%��]e��
b͗�_L�&� ���T�[,	�j�7{�4n�2�F�$�V�Hϴ/�deIWE�Z~�r��)�cK��mn�5�������ZK\�n]�eM��O��Q9�@���Vy�#̳���P��ttH�TJ�)�ɸ���DL�AГ%9�h���`P�DI����&�P��.4&}�pY�Ñs\�Cr濛��*Œ{��|��1mKs�n��-��*���: ��̚u��5�O"8��r�	:ǌ囉Ju"�j��'+50��5���7�N��j̹Z��VPG�,ީ�;`bԸLY{XkU�O1h.-�{���l���P��df��bѧ�*��٤)�W��s)JֱT�X81����:j����YE����H^�k4�<��:^�$�L��*S_��u�;�*��pW˚M�^�f$+3�C2�:�;�I����Eɮ)\����UTPzd�(ȓ5`R�r\Id�+!\�r�ei#Kv�M;�˧SE���e
p��7[��P��z.a��PRr�F�,�m�(�bpJh'T�O+4ѭ�TgR#�)��y���\�bjX��=T�^#��S� �0�N�V4��l�6T�&h���i�m]$*��46���qhy�K+��8��&c{S\i+�S�İ)���(��a;��;L[`�`r=�a���Xu�W�r��yC^V�r�J)�]��r��YӨ]��%��bņ�4�X�]�Y�ET}z�e�u,��8�N�[��B�
ȷ%jN)!b�h��kN�����.cW6��xMQ@��
��Y��[YF���.-I�:�wr���V`ԱlnR�ajX��Ԓ�ݥ��â98�b�6H���������J��eL�Viܨ�d�Y�%e�"��L��u-jܛ�A�V���ki�f�$�x^j��f��4�`��/a�m�M��+֩�N�+aɭ�1�DI.PO�Fxf��vb��^&ٙs�e+Ϩ$�_gQ��l3oC�1P�4(�R
˰ꂊM�7e]��N\ڠ���'s����bڲ�gVf��E7��G%f�m*�L���.4��j�ޑ0
K^���Q�y�`A�N�j�T�u���m�ob��7AhV�[*\�Km#$�.�݌f��0(T?b�����3a'st8)��wU�f�Eu$U�ͼ�.�s��]��(X��RWIм���nE�v,/f���i�.�W���K�]���E;V�o�+n��6����ɩ-��EZ�mqk
� [z��%��K]��F�]´@o24��ǙS�e6��P�r���uN��q�3vm�����9�2�2ެ�F�B�z�%u%5Y����z&1w�XwQ3 y��c�R�t��5/�2Jl�C2�����3p¸no[�S[�Ro�6y �oob�V�+��I��ȱLZ�`[.��ɟH0��m��{ZU=�ے�4�j�1�f�A/P�ͽV��BHv��vpL�-ek�(7٪��jЀU�n�f��zc�9R��l]�ͭ5K\h�[cK"�T�OMe�(4���a+d9V^�Xvhsm+B�еYXp�l=��k�n6���7!S�Y�8f��2����Ά�'[�`Ĕ�N��׌*IB��X�є�J!�+UoR��:��Y�wDV�u��7��662���*2C0I���V;��� P��70ïU%��qa@��j��o�f��p�%��E4uB��;�������T��M^�+�{4��AM��>ҥ�.�9��,ٛ�����h�M"k)�PLs+q黵ѥ��kX�b�޺K03cCA4햭e$-��F��wm��
���݂���0@�"�Î�F(ڙw//\T&7��xĻ6S�ĵ��z(=�)�Yz(Mʺ��2e��7�Uv�S�� $��G35��rY���m�������d��u��H����.�
O��j�s{AY�n�����)༭��V�:7pF		�mԵ�V]MN���~��͛�N
r��˩w��u�iz�uw[A ��(�ݷ�"PH1�ŗy�P:�Uh.*����0eu٧6�b�tӬ�x�S�pc�ɔ��@ *�wZ���wn�ۙ�Kzb�SmF^�
�KKi���c�E��ZZY���)���cb����!��k��+)%f+٫i���ǥn�m�+:�e��ut`��C��S"�&���M81[1ܖ$�{�f0�n���k�s�&���bb�Bi�0f���m�Om
���2*�7�SB��e^�r3(�{�	�&���i�@��DnƝOr�d|D����y�sv:�B¡�}�MT%�OH[�����u q�	���f<�HnGZ�.ć�F�����IӒGi�7,l,��966F�����ȱ����.b\�Q�V�+�v�ZKG�[��N�^6�͈j��ɑ`�̫����u8EYZ�U�Y�ģ#@9�P��˫����hj;HӦ�D���Q:ͤj:ٿ0�o0V�r��RQ:�ܵ20��nYA���`�smn�m����{��X��6����ۏ(v
g3�9���w{ ���5�Ԫ��,���D-;��]ۢ��{�yc"t#T"tiR�5�ŵ� ʹJ�8c�6��smMB��ݍ,���*�+%<�L�f���m��Ub[X �@��5�eV�z-����on%�[y�c!%�0V�`mk	�h����P�K��e�B�I�3wt�l�e�5�����OwU�*9��Cn2���ӓ �m����,ߵf@�>(����#���fPb���)C�FSp�J-�5pd����2��V��2���z0�eÌܦ�ZWr�X�!B�h�Z���)n�b�xS�k���Ur�n����7��A��ai�1l�w���F�xj�Kw(QW���-̳2�Fn����&��%P��!�,h��J4@��5�7 Tb�E)�P&�]�˛��(:C]�4��%l۲#?M���
.����[ș�hh���m6���Ny��751�־t0E��[Ϩ�6��/r�:y�AW�Ř^�-����'v�x����DGGT��MHh�Am��eچ��լbʛxeS�+b��&���ٵ�����]v+��:�W�*Z27�6�̲q��O8�4��m����Z�͙$�J�t���ڽ?��0�z.V�x裩�T����;F�s�ic���t�	Dr�ˋF�F]�f��L��
�Qڀr�<X��n�Y�S]��΀}J���]�4M�&\�Cs"�i�0Ub�-26)�H䣿!iMF���02�yY+	�6%��l�TCR�7�M�*|S�j0a�b��!ʔ���Q��U*;2�`������. u�E�)	���d�l�EL���Mف�m�Q�m����n�ky�RJ���o.[�	���Axq$��%M�H��CT�T��mS0��+������l��/L��7��*�pJ�i�^�h�#X!ј%"�5��a_�Dc�;.iYg�U7-h�[�&V��U�{z"V��P�m9���&��if��	�Ou�m�ԊL,k]Tp��Qpi�X���s@j�V��S�^Qx�݁���n�C4�!'l��܂b[��*S� ��1�0=Ӛ�'
��E�:k`S�ףf��EP���&V�;,�P&u���1��s-9��Y�L(��e*��Ś.�I`���YWQV���V�`�r�c$y�Ň[�#��r��hP2R�0j�3Q�e�V#�Zh����%��Wkl˻'I��)�h�i��6�1��D��ءG���ʸĪp,�\�����"v$��4ءcZtE^漛��b�)Z4�m� �'1ֆ�Y�9�=�WyGT��S"�Uܑԫ�w[{�Bn�s^H0��
D�Y7kv���5�����W�"ĭL1)�s*�o2�t�䡳LQ1��m�3�4@&<ǦLx�B+U�ʧL#M��y�V�b�O����z��l�-���l�ṙhel��Z��$�<�Ӧ
�6�S�jD�]ȶ��/2��]���dՑ^�vm�СE8��4ޝP �٦�ӣ1c[�R��kN�-[`
Dzr\M:��n��۶A�������i��N��� 4�H�bI�AkY��S;vM�6�j�8S�h�yad�ńR�R�Lj\�2"Mbʧ�*5w���ŀ���OXD�]��굋ׅh��W�lx�Өd:��J��yi0Z{J:]��Q���װ�Jel��' �@�;�a�qXʹ���UN�1��g%̭���X��(�X���F�6a�TW�'�ֵ1���X01���a��]�X�)B�<�eK�\�ʡ��ŲXƶ��^o���D�-�#j �%�k�h�c��
xo~��ij�h.�\N�� l�	��t���2Enҩ�z�P�q��`�0RR�I!/2��Z[Ej�m��y���՘�('�V]!�n���F��t�u���x�֎R�庉����G�8)�0��B�^�A���S�z��|wiY�vQL���wu�Ay��4�[X^ť
�sHti�nP��7Z���GF��R6N�
�ǃ[���YZ�A{,���w�k����ڎ�9o����T�����Ǡ�Ycunjܽ9{��i��vC�y�2A���U�Ov'��}]CJj�R�	�CN��`yx�T���]-{&*Dv�* ��oF� ٢�:27zF9�edK+:ň^ƭ�n����K�n�0�h�'ٹ�A�� �&ȉ]8Y��<Wc%��M�K�H�y�eB.�E��i:yh��\���0�ibL�r8��.�4����Qd��.m��,˩`Y���cτ�*��g&ҏ8-�@놀vL;�2)���	K/eϬ�5P�v��L�J˷�ڸ>n`ݹ
`��L^�\��<MÈ*w�e�N*�x�[��m&���5���M��ƞ�5LX�7LW$*�'�Sf���͒��6����m�@�yL.�&���d�/Kx���fԃp���{%�`��Su���
�ȓ�]5,�Ão_!EbIV���J��bQ�c�{��i�Q(�����L�ͅ�]������u�[:��.�+#WngP�����1L�����[1]��-}z�6��u��,EK���ko�Z6�ƃ�6Z���d��re
V{��i����HT,$�n�u��7Ji�h��*�7�J��L�$���"��++jPwWB`L`��2貶�S'^���o&-գe��Z��0n]/�s���4Z�<���C�\��LBww^�J�X��[�Ӆn8�%�x�����4[s!����r�H�:â:�w$v�&���h��d�&^}5���77P�'*K��O-��ڰ3�0)�7)�,ВÒ0QP�Z����-o�Z)��8	�앧��ټ�했�P�-�vBZq� n[�v�[7`�w���^��FÖ�m��K�cRęwR�'6�n
]m0��l��&S ���j)�����m��Z��Ԩ^�k��T��7�]���xY�we�Xf���X���Q
�7N-���������p4�(�������%��U���5��[x�H+Bx��Tz�SsJp��$�5���Vӈ�H+/m�],ۇ졨5b}tdr�R�\�D+`ԨD���r;��kK�T�KtK��g3*�J��81]P8�!��2j��褢#F3�t���R�����kWQf`G[���4&BT�J���DfꚰӂU&ڂ�\4p,2X�����E�9��-É��,0�ґHf42�V7W��Ǵs�Q�1���@��V/R��!�X5z3�$���]UXx�1>�.��7�[�k3QM�k����'OD��
���:���a*"�c�0�^�u�]1��m<����h�i��>�R��w�1Fpi��ar�aTar2T��v]����
�i����LCeK���s3�Wi�KbY1ٺ��E%H�f��X��)
��4� V�xqX#4��7��Cw>�W��i+&�h�cM��b� �ė�V���@�M�!��S:����r�"���l��m&��:N�V[�K�	��'3݀��I�6���=�6v��ku���6��wb�t*�M�L��0`��fۓU���4<����$0	�kT�FP6�B��)��n;��Yc9v=[�Q]�\�X�EuqZ;cDx�b��m��aO(����Ӧ�9N���4���PB�F��.+j�_ne�TP�\ߥ��2���Sf��l�-���U�ѐ���'unڻ�Ԑ/�6<kw��kW��w�s�t�?���(m	��9��L��e��$����:���jR�RY%�YvCܕm�cA�ys%͵u6U�or�Pl֓��;��*�m �-WCN���ђ@�T�v���ȼ'�*�fn���}��� �җɭf8YTN�[�4������[+b<SJ�p��+SṮ��Uk�ƵmK2Z�xa�>���t\�����&	�z&�3�����bl�S-��h�g��f�N���o�84�M��5s:ޠ1��>Ɍ+�4�\\���k&��G�掽�If��lh��8G�6�$d�sA���GVf��:	�%�e.�dX��Gt�h�'N�Ȉ^�@Y\W�_f.�щsY���/����X��G���%/M�I`��G����/��m��iؗ�~���}�0,p�e���U� ����Ӂ܂��C�|��>�Ց�n֎�v�oӺ��p
��^��o��V���:a��X��9���f<���l�:�kk)��v� �He��䬈л�Yw����ٛo�ݙ�3N�#ْ<�3F�f��d]*w����k�fpe�z��hv�8�Z����,S��p��u���A�o2E7r����B���Z���"2Nk�2SM9�.�u,��Y6��({9���\�H�>�7]�׽+�bf�Ę�:�:R���]1�;Q���T��9M1�(,�b:��e�ķ�
Be1�+Od(|̼��G2噱���qW<B}3�D�O�Q�Eq��{���	�ɢ��\���d�1ʂ!+T��6�Ac��ݵG:}��Kw�\��B�pt��ٝ:N��S�硍U�[�.oT��ڞ�����)��I]>|NaUp�c�[6 Q��Q����ܻ�C5�z�J��vI6�{����u7�/�m\%o/��ެ��1�QK�0����0��	�`)�ۤ3�'fS�C[2�sZW:ma�E���u�K���q�1ع�i;��c��� ��34u����5�=����O(,�j�I�:]�g��mo-��[���;3]6�va���w��7�\�7Y��mn	���v���F��61t�Y�	M�)�b����.���-ϯԫ�Wfp�d]���_͍\ս�uv�sRT�]�wa�x���0 �U��	˸����T���ɫ ����q�M޷]�Lc��������U�Ge��G"��jp�����M7���wvo��P�>���ֆ֛��=�k�Z9��S�D��{���l�ǩ��lB�).VUb���na\��N���Y�ћ�G^�l��7���ҋ���[0����"w�SvL3F�әn�w:iэ�Y|#U��a-ʥ�dD}�3پ����{rm3��H�,R+U�
XY+d�K;Biĥ�V�	����L��J�a�SKZÜ��iXeǽ
����[F�m�= 7{�N����t{K�7bTyO�q]����v�ij���f��%Δa}�d�����2�7����uU��6f��E5��Ŭh�9ӄ�NZ�]�o��!��E	�Գ���le�J���.��P�����P��4�B�y+�,\6ܥ��@��5e���$�C�Ī�wO�H%�8mj{v(>�'<h��F��iQ�3erʻ9�)�A��&�Vj�p�|�uw�������^ʽGją�C&Ϫ��m2�D����D7������A�)��"�AfS���C�|���#2��U
s0l�"�ѻ����]��(�w��]B�u��C�M�k����b ��U-���ND_ F�/.�(���33nL=����۲�D�Ka�b��WZ⁨,�qX}nL�������o��ݞi�T�V��}>��iZ�a�\����X�[��S΄��-�Y]�Ia�f�!�OP��ī.Wm*�`�Yg�EӖ���p���Bn��e�$�>�75��|�,[9ql.��YY��/"����#�ͽ{*L��Hx��g^�t�`"��f�V�x2\�Љ��KV��3�-����.��!iб.����f&��%o.�^�|����,�v{�I �*�*;��[� 5�E�)O��}���fb���g ����Y7�c@=w���d5��R+y�tWH>w��S/d�U>�m���=�Ըu���� ���:]A�6V��dk!�nIYr�^�-(�P�z��W.�q�S_<��qCe��r:!�o�W��9}�uA]}��{ݮ�ّސ��.i�:�٤�>���#��L���-2�a{�*��[��.纕��q��v�A�U�!ܩ��U�v�eBV:�yQ�B��ѓ0�s��
u�)`kf�oh�����2��օ������S��u$�9)����_r�V��%�v���@ؕ�p��k�khGz��L���s
7T4��N�J��Ǉm���"��'J盩�B�L&��O��1���+���c��s*�m,L�{D EHn��u�{#�_\��D/#R��2�w~ka�gEep�-��A�uFsh^񣓜��+��mbv\�Qu�4�n���A$�B�9pI�eԖ���}��W���ɗ���Ǿ=p��ʂjo_d�n�Is̻��.!�u�������>@l��.�w[<�M̬T���`�d�F��P�L�BEi	�.T4n��sz58)�BGd��t
x�|TZTqD��32�;�D�Ӊ8>�L�.�e7W�R�n�<�]��]�܇ڛ{�[��� �}��4�4]SK�Zu<�F5h��lYE!miv
P.��}��.��q�m*�ъ�ff�v��/gUBG{"�6�(1|j�ۜ�L�ψ�6�8K������pL��l���Z=�R6�V3)�=�j�ڎyx�7�*�0q��V���',+��4�073������G!K:#Rq�ghgo���G{%��őzu�Rmr���MQ��3 �c]�v8�oU��r�\`v$wh)AКtb�E�2ج̝t/�bŸ��ot�/%�������TQ
DV��ʂ�H��V!;Ȯ����sjWM�0_h�4���U�X�{a^��n�L|�i��дn[;w���(dʦtY�5��w�H��ub|H,kg�� ��a:���]��&_�kk��БgM���"�I"��8��գPQ�>Mb�r`���f��P���8m@�)����&Fm�@@t�U-��.B>�@Z�<8�_�>�j�����o˨��na;� �YM�J+M��y2c��[3��M-6��5)���pk滺�kU7B���	�C�r�*\��0֑��Ht�z�+�t�}GU6�+�q���l�Ȼ����k�U���o_!*d�O5K.z�s��p|3JJ�]�P؇w�V�u`<!�6#�E��%5���K��vE�,��
��׭��f<�HJ��� %�VWT�A7r�â���(!���+�b��V)w��S[`�=:Q����+��)��V�u``�w,Фe���M'JCH��<�ȸ���O��L�ד2��La��Yĥ9y�D�	�֝�j�[ᵈ�9��.fȤ�VT�id�7�LO�n�v�P��њ��eY����s�Kz��De�jk����ݬ�)�����{'C}Zr���&t��󻘩�Sp��aG"!o&!�6�Iݘ��T�L�8f���u3F���v�낻�C�������a���e,�ѵ��D���KuwB�w2�dV[���\ ��y�V��+zJ��Q��h냎D�2�l�<B_m�"�`� H�~9�b���{-�n�xL������oZ�C���.]�.Y�V��͛[	�pb�sD��P5��W�0;���u1�b�]]*T��e_gSn�9�����eԂ�WA���g�)wV`��b����/D���^�J{�i�Cm]��m�+u�H#��S���06.+�ެ��8����t�)rDnJ�b�$��Kj�e
�"9�c��U���t|#L���2�]��ԅ^��WV)�����ś�)��t�oM	�hՒd��*Aen1��HM��̫�ZJTmiu-̺��c�]�ݴ���b��M���!;�X��z��	�����T q��Q�,�(:_IB�N}Z����p<���7ʉ	��67Bk4q���"��ӣ_�\��R��2^�&�(�v�=�vHeM櫐��''0w0�ųN��;6�s��0��ȩ�l��ʷa&(�#:���Ư�8�%�}��GE`�ӓ3�_A���^�z�h{��.�Gy�Ԕ.�E�2u�5��[�Q���긪�Y9<��=Ad5*J�l��oT��=h�dc�tHN���ɶ{['��K6YOS�f���Փ����3/��d������6�l��T�r��Z��o1�a-�3��&�SR�UfH�r�jO�C{x��:�%;k�X�*�.9m���Y�a`��u0Ĩ1Յ��Nͺ�U������;3m�ԝ.$\R.���>`A����GaL��Gysv�ˈ:�bV�1���{i�POrJ�Ç��[��r�[<9���)nQ�%lӇ,�q<ѽ�w$L���X&1�AxO�C���4^L��E9�(2V�U�x�+��i��o	�T[(�|˺ߙJ��,h43�.��Uκ�a�q�aj�n���O�R���W���>.����Vu�[w�X��b��ҕ2���ǥe 4̤A�]w��U9��4��40���Q��8���݌�8��ڐE#����Y�VbU���3e�8���bɂ�f��E�ɰj̢VX/L�}�'\^�l����1<K�ν�a奆�F)�	��Wb�f�t��z�c�-�Z0�Ԯ�b�N��ۀ�a��t\�5Mr�<J�g7lJ�N�ҠAh�P6��ӳ&�����;�6l"��/QrR�ƚ/B����p�wL��}Gq�G)�\���ܮ[�����(5��/Y��jy���u��VkBĉ����K:3�&��r� Y�ݾ9�n�vv+:���=Vk�_G\���Cr/��u�hu��M�DVh�Y]bӬ�g���'92�=,���{O���
�uں#��kgA��Z9�а����9��eVT*���uX$ͽ�h����v��xU����Qhs�3�y���\Y�������#8u
U�xI\���;Ó��0���}��v��"�#��hmKVw`������Υ�M���ih�Ý�s��C�
��s<�8��Q�S�#����Mn�\�z�p(�;S�nR� �ͮjv��uNt8��O`ҭ��I�m��\�{K�kot��j�g\˘�ac���n;@6����:uc/��c6��:V�8Z���ޗ�s��Gb���Sr��H<�.�N���2WkwF��>���Lo��L[&���쨈5�Z�n�ah����Wt%����#��B6�!� !�ǰ�<�52�;���{����7���8��E5^��V��:8T�+��چjzxd�6�����.���Q��_W*m��9ȏ)��xA���yr����m7X���S3!�de�y�ޫ��t�!�rf�3�o��m�N.YƁ�'�k�]t��Qi�"�Dg>=i1l�;�u�∞u9Q՗�Q��I���^���sy�2c��o~*��q�z�Q1y{��kM[��ᕙ�bqf�6���ˍ>��}�Sf9҅PX�0��/�T����xj;D�5!������l˱
��C���������o����Z��&Г8c��1uv��,\[eɢ�	�c��G:ъ��n;o�h�iP�1%u�����$m���3���m��w�w��Z^��æ\WY��;�
3�.�c$��w�'0Py�"^Y`�g/��pM��kN:C: ��v�o^���2��F�R��3���wiZ�s�/�YF��E��zU>�[!`/�,��,Z�|7A�	��x��*w��Hu��/�6���u�ȴB�HxV�3oK�&
����n���z�K��&M�W���w)�[�t��J`S:)���Y���.nJ��!;z�{̙Q���w)v3�$An�vl����(����P��¥y�C$�/o:�EƲ��{����A7rQG�;4��W4�4B��7���n�ξ��i��.]��s�����*jz���mE�0����*n#��3N�۰V��}^�ͺ_5+8�opB��.P����4��a��/2l��⮝�t��\��b�OV��̃�n�]I���"<Ț�Ym��]p�e��Q�(/f��YBv����\��)^���K8Nk;>A��PďFE�;���	�x���vg7��
�'<�x�6i����֜���Y�d� +�Ug]'�ݱJ��|d��_[w�eϕ
"VÈ>��j�6���g*jB0�G�o �%s���h�wj�P�RJu;a݃WӁk��$Wd"VL�F�y4:E���q�v��R�i3�\�:ͭ�m`ΧF�ڌ-Kbi�����{
ȸԺ���Boio��#�3�r��|m'��X�[�;%�׊��eL��\��a��)��:�g9o��Bx�K�6�j*-�c:)������	���ҚÎ`�
��q�7F�w}���֦�`�p��e��]h_KZ�����nSp�JxVv3P�9�ؘ/�^���b��Y���9��p�J+SYΆ�Fuge�[3@�H�����qҴ��_2Vs�V2�H;��2�؎��� ��_�6uek-C�V�:u�]sU��.K��}��B���]5N]ڬ��C�ƻ�U<ޱ��S��=eF��7�c02IL�%WD(E�5v]r�l%hP�8��1�tH`'}��d�qv�����������ă:��4,'��1y��U�ʘ1�yj;���m���7gf=5g{����$��š[\]`�7�2;6�QRk�{���%A�c����5��h\�\4-Hy�P�Z�3{SԲԽ��)w�e���Tf�N�\/D���As0[�9֩Z$�j�T{��{��|�LɈ�ݕ�t*td�}��|�cO9Pٖw�[��16E����o6��wL��=�v.�2�����wK����K�K$:%
���k��.�i�X$��z-i���F͔���Ωx���۬
�^#��s�6mNr9��IԻճ�9��-�I�ۈ��'$��)<���}����%��4���J_	L0*��"P���:~����;�ׯOM��Q���{7�s�:-޾F�  F5�/�:h�E�� �/���G�$����a����ƌ��o\���{�1��v����o��f�{+�z{�{z��ާ��m�kmm������V�Z�������~�����*����������?�����%�~I&P�OњS1�K�]�_g� �3&\[0��_
A�����U�v�u��-}a�`V��qy�U͢�0h�wx��snsn�M�p٬�B��X���̿����L���o������<_\��j�{H�R�W4����te��4wr��!�0X7��<xadw&�W-�fα�_�����|:չM���ޚ��W�]!���pk��!���gS����j�+s�U��Ԏ�V�O�����&��Q`��.�j�eD;��I��T�z9v����7X��R+�E9[m0H?.��G�\&+$jF����Z	��R��Ŝq���Z/!7�8*����Z��Rĭ��ۙ��~��݁�!�Զ�qp�=J�f#r��6��{��$�����Y6��!t6��[n��D��ser����WW���E<���E��S�aUD�֝
^�6���gu��f$��*��� �嵭�8J[�k/:L�"�S,ꗓ��FڨV��k�u*�n;1��n��8�sor�5P�8//UAj�yĈ&D�����@������w��ۈ�H;�^ǌ"4��VZv���Gq� �p�q��,��M�e�����)�I�x$26�`��E�����X�R%�w0:3�z�r��ٟ5�b���B��qBZȻ�#�}�5��cF'yS�2o;�+-^X5��޶��To�%�8;2�r�!��+��!��M��sd�p���v���2*�M��J4��:K�����5�M뀗��������k��0w� 29����v�w-Jq۠˲�)M��t��4�6n����G��9�t��FjlY����s�aWD��t��*�W[��e��n�M����]V�;	�|u�7�+,���\|1��"��N��	[`.R�],�λECa�0��38��Ov�W1���&}��S3�C�.�R��@�5�u��'z�.�/�s�a	^��F�S�:B�w�@��L`ơˎhXC wH7u��;[�������e[�F����pՎ�N�o
�պs�\�s)�%�7�f���P��Q�ۀ��ڏo&�1[�n�	�n�1K�1Ч�wOd���[]E,
%S��ag�׌�����1�63w����ܝ��K�˰nA��H�R��nn��e^�kR�+:9��ca�9���:��9f���Y]&ӈe^-0E�\�!1�G�6)��b"C=e@^,c/\�X[�b��,a�I��U�wu��Tis����*�AM,�';������q櫌���E�q=A���r�P��j�M�G�D}D�	M�Jp��B�s����v�k�ѨZT6���ۚsF�}z(^V˭��9�T(�:���^�Ӳ�j���X�,�a���3����z�>t�P���x@9��v�tږk�H6�_v#Ì��~b����B����Z{5Iٔ[+��ؙ���z�L�Y���V�PJI����n�$xl�-$�idXY[tZg�E�ݾ��p��.��^�6�pc6�Z
��w�<��}�ӡ/��\�R�U���5�ڙ�����7�duj��M��F)4]*�ٹ$��s-�m+�2�g$��X&�S�N���ú��3f�vsg]q��-�����NVw�ڋ�k3�}R� s),ꔈЯ3����/���V���З[�:v��a@Y�Ru�K�n:,j���p��ླ�O��될Evb]pP�8�e�)�/���f�Y����v�6I�B�����cob']ǜ�~��e�����IU
}��!x�.��Z/zqfBmTh|�^S�Ww�;�.jn�*7�qldCkL�zI��t�k��A��(;�7o$�˹�(uZ�fl��U$.`�;Q(2����\�9��yHMG�R�Z��� �r��Ǜx29�n�rʎ��-Ũ�6��}����D�B�g`�l�M#�bo^�GoLp읪�靱�bv�1�H5y˗.����Wi�(oJΐ鿥I��_� �X3t�r��6�-_R�f�gB8\ˌ_tݫ �3	j�ublL�h��}�7�ю���U��Y�*,C�d]��ch�Zr�!|�ǼD�9$5Αhխ�h�]�n�[ǝ��jI9_b�D*����Yd���>5a�D�"	b�oJ�0h�H�XZ�Nj�7��q�-mZ�7Yk��K�g0P[��C��c��&��CW"7�w������T]w��96�ܨVҾ��a�G/��u�J�9\kY5��q�͇C�M��V�W��"�imn�#T���՛�s̛���X�RCH�8�4��\��jH�X4��//���P<�+ط/{
����%@��8h��O`5�������˦m�-�Z�Ωէc�mh�^�T����[��ta�^gA�W���1��� �ƀz�� �;���ʙ���j���M����,o�W|��!��u�����S����u
<8\	�6r�|ICN�������U��t���n]�.�v�AX�)72V��!��v,ڲ�J��n[�n�Z���P�4'�m�"�络��ݺb2:�ٽ0��p�����'��*����_h�)
�Qi	��A�<�쩵��]쮺3��<��/l�&� ,{�0p��$G�+����{��pӽ6z�=L��gk)v�Kv� �1"ڹ�܉�����U�u�
1�}8�VUM[��2��@�J)�o�ӫ���H�c��x`�ې�]u�g]n�V�u�gx-n���c��VKsC���b�}�I��a��,�w��"�K0D����q�=>;z.���� �a:
n��ke;�����(����8S�u����XA;��-��䮚�F�j�3��BWإ:nG��UԷ��$yB�����'�=��+�#/m[��Գ�0*��xd�����1���1/0*�����&��"�4�9�\�+9��Y���<�%��a�ͷW����F�x�ѥ|3%��{D��ܡ�6nLx��I����}xt�'�-;��7tkYa�tم�ԧZA\��/�]Zl�)��/�B
�FJ�j����)J
��n�����eˑ�[�X��Հ���A�l�4]��M�F��z���VXܡ�2H��2���Y��K)*��p��
skK�BB�Arܘ�zq��K���2�U�ʹE��@R�	��h�2�B:u��Iy���p9`^੻DT��%Ew�ᷭ����Y�i݃r���lMm+5�w�����׮+��MD���^J��aG}P�=�4A���
+י�N͝�hp��8�:�nh��G	���w��C��T� R.�0�2����t��0�]ɴ�r� %=�1�㦬ɰ�\�Q���ͧ��֝�F@ޅRHo�=�\���z$B�L;`I:�jJ9Q+�̛yke�)Z���e`�ձp�WjAdC�{�ͺ��D8�d�%�;��^��nG��3)�����**�D�9Z�VLr��e�٘At�vZ�B��Ww�6���)��B����Fm�c�̭Ѧ���_*�b�v���G��P�Vf�v����aj*<�*Lpڧ@G�3^JxJՁ�[Zkw:�=h�\�9A�$걗���B���p!��J��B��[,��K�X8��1mGU�ie�۶D�w��A�6�DUK�)c�!
Wo�cXȵic*}}��	�aI}@�t��gp�KCh�4�Bj�b��oH�N')�\p����R�����Z5R�z�4Av�K�����J@6[53w"�W�e*����Ŭ\L��HR��Z�m�[�V4Veo^J�X�b�8L�J�X\�}��X�7�dt'3g�]��.��wu�u�ݾQ��o4n�Π�0��'�͸+��.g B���7�4K�.�4�D<rb�ѩ��S:�%��P؏J�
������f㛛5���"���y����#a�!P��6��u�q��U��R�S}��ӗ"r��c|s'3R�+�����v�\���I
Ա�OQ^CH�����c�Vm�,@��a"��hԦӤ�]����K!�7�����ݫk�<7�t]��LXFvi���RL��Y�}B9@F��k��v��������m�`�
���
q\Y�/��"��� $N�g��/h�Ci_Y����Ti�շ/�p��C�_\r%�pK�ݮ�.�sz���E���]pf�2=e�A�b���YӚ��s)-��"�R�������>�	����/BX+FAf�q�(���s��cq]_pp]��j�u�h�\�z���8�i������;�r���8�1Wvk��5M��W[(�fIZ�v����A^�%赡ӫ�S��g8�}���iآ�\��dR3�K�trۂ9������o�NT�N�YK.<ܦ�j��p՘�%3��9�U��T�n<c�\b��Z��ۈJ]]õ��|��Rpv랽��S�9RAm
C�e�z������=�h[��:0n�h�4��N�뵀��i(tR�^��1�5�X�\��뼮;Y:);$��p���$�9.����WV%�!��7xK&ᩙ�B̖!���м0����Y��]P�ffA.]�����2�d<����-���r0E�u�J�Jl4ɓ&��fl�S�b��_*O���qճhڭ�d���"u�ob��.��u�#���tʏ1 �%��oQ�� �M�рo]µN��m�6��t^]��r(�w�wy&n멄�Q'��#o,�βVlh��-i��^�:21P�W�є(�a��j']}���jLO2L��GY�A�F�Ը����)��t�����ܚvY�u�f��:���n�W��"�l��Em��^�8�r���36yҝR���˹�>�H(I��t6�d%��z��F����;}΋�k�F�r�C��%�DYτ�oj�@ՠ�t�ř$׭�wo.�>��zѭ��:��*�N.=�*.Z�s��Wq�M^�鷎�Ŵ:�В�]t�ũ4\Aj��lN��JD�[��ire�>����ݚ9}�zX�z�Ze�Gpw}���:[u4Q�|w���u��Sذ���̣wE�֊��̤il4' :���K��mm\��9�-�r�.\�S��x�Aʅ���[�~�]��,<���5�N]��E�ݜUt��f��H%�-�"[VMj��t���g�#�Q���v:��z��
���C~��fv��싎ǳIc*�#y������vG��<�z�AAzu�5hft�
�19�9�	�U$�����lkc�HU��>�O6�		0��@欥�;y�������S4�{W�n!���9�)HEK$Q���J�ո\ցy��u����@oK،�z����e�;��v�us�V!}�2zP�3L�;����S�ȶJ��;�¢=�lh�l:��4�sY�I���eFNr��r��'t�	��YSd��2�urRUΛ��|R���P�8��)�%�D!�Ɏ�y+��d4�m"k���t֬]��itئv���΀�7iV�<�7���-�л��U�c�Cܳ�+Y7��ks�)>ͱe�}gWc�y2���f�r���g9���*\��gI��pѩ��%�����󥼔y�$+X4n�=�tҡ�QL����vb�IM��Vl�N���aݑ�Z{RS����j�TW��ރX���ꃍ�V�ps���WQ��.Z6�y�Y7�)��Y]���U ��֨�S�דe<����HXڮ�	�j�Z�R���6���^�sU�qT/$Y2�ѓycV�Po6+`��6o�J�r����}��ټ��ܲ�4���B��rŒWz�a���nƏe�v�����5�Dg�TT�IDo�N��@dU)��<�غP�ȫ���&^fK]���.�:�e�*k�:I��Z�����{�h]\�87��)6o �ZV��u�&E���E�a����`�𠶷n
�D>�!^�,���b`��+M(��`O�.}t'ϱ�1B����c5)s�9�Ю�<�wd��F>u���ok�gG:�VH�e.��1�y�&.�S���9�+H�7d�o�[�i��A�6�'�x���2rH��N�qL�K���{x4l�um��/���&�J�fi�ߥ�O�K{DheG84��f8J�O�m�U�,5�ҟw���l*a�joׂ�L��+���cQ^8h,�Z��IkV��㗔u������őD�f	���1A�Xvݽ�do�+BWY�8h��$:���jS�|�Mb3 ٻ�[a���DP��6��|�+���U����^)��Z�����'�|N�t����{x`�clfsq\����� �Lk*��{+i��Xe�K!U�r�Q�V��*�:�Ě�O"�������Zs�	H���@n���ӂw3(
[J"]�ea��c����|˴�͈��Rޑ�`q��%a�	ʠ���
�	#͏sF�<X�sC��+6afwno��,m��f���LF�Tf���Gv�5pˉw	�P1�H��di��w>�g��\w!`�Ǐj��㸃�S��`r����������E��:k	�B[y(�	u|�G����6�b���7J�S�1�i����C�u�<Z��A�>�����8-1�-�wr^a�(��p'E�k4s�2�C7M�l��&�(����V�ΆT#��Y{E۰i�OS,�ޫ��1H 7�j�F�:�:��V���S�d4�ݞ�.Z�+����d�P�FV��>�9$�yR�Z��[5N��6�E�/��fb�9{�;U������װئ��Y/J�g�J�j��x9ޞ��RM&�t�y'L��ҫ͂l0&.�'�od�y}[����}��Xk��M6+�%U�&�����   9�s��@����������~�~{�߿~{���~������;�|���o��>������Y)&�B�-�?7Q%PH�Dc�LQPIB(Ӏ����E�c"H���so�_���wT����t$X(�R�B s�n�pqx]��<5��1��I]ܳZ�m�oi:zj��n��%�v�m)3�u7�f͒J�s��Sr�T1P#����]n�]�8s\�K���dɸ�0X��kV�u��/'7�/�<��:雫�_"��Ų��� ����R�iL]�"bwa.,=�Hs�j
��	��k8��F�XЊ�V_Wv̳��޴O�F3��ɇ�A�p�Iɳ
w�V��\�2>��\������{g����3�˨�a�F,�h�2�F���R>�l�)�>Q�9�S��J,���(-y:����x�M�&�Y�:2�^=��l�ʷ�����f8\���  n�zz-����.���P{��8�:�}����9y��0i�z�t�z��Ճ&�f���]6@\�_K��u��);I����o�i�2�����Cv�lۦ�bq+���	ܐ"�y@u��I�ü�|��RB����ř2�uc��(�5':�^:��Dr�>�[.�b��P)��1Ү	���{���Y���0ͪKx�g'�x(�z:�N��	�Z�s�āA�r�u.[<�=P99#`�k3�uZ�u�ޝQvU
5��3�q�ͺ�%�Ҍ�%����	���읳<�9���3�u2�m�#Euۜ�d��#�6�:����j	 gI!*H!��!%��.|������e0܈2�h2�A?��
*)F�*�[:	�� A�eAF��)�R(L�̂%Z0F���%k��r���]�(I�v�i��NQ��#)أrr쑠�SPh˝��I�M����I\�i9�7$ƎsF	��Dc.�L �DDl�s���b) "�wuݻ�@�4E���RT02H��	�J1Qb�QbQJ)�}��d���2b�ӗ+��s����1�%$��H�	2���RE��"&,�.벳�sL�QDl	�JAd�`"����e);�$�$�c2�˘Q���lR6@2FI��I���� ��AЉ&H�Y��ȓ$�� $Z1�$�	Q�B*��h�Aﯝ�^��ۯ��k���李GX�.�cm�b����q[�Rx���w�[{�n�Fv)�i���J�&��ӹ{|";��ة����R@�Y�B,hJM���cXc�8���k��s�����4ì��d�e�C-��ލ\�፦��K�Vq"�ل�ɍA�<M���]vծ�'|5�Dٵ�n���%s]~��L����#F9կk�I/�n��u�`�q'\w�A�w�3��X�oޣ/%x���"�c����7����\�_u���J�K|�M�]\*Q�yz�ʛ]+=�z�׏��/�?;�1z��z��,�l���a�K�E���#O^�!��i.�!>��B��?�3�m:ĸ��?ce�|�]�n
爙�{�3twH�'3�����}�[���]'����{[u^�{P�	�TM���P;��bt֊��ė�þ��5�&�~S�nM��v��<>�=�*_J{5�MlY�R�I�R���=��C���~~�>F��jY�gV�(��Gcu���\�c{�V7�u��쫊�b�|�!+����PoIXތ=W�PVX��i�6U��&��Y����~�I'`���㶨��ڍ8��v���v9��-�;N�,�˵[	JMm���*Kǧ=�!�w�P8m�����7�{�P<��N�,`���l�8������ۋMH����o������׏�7����<����^�����x���?\�ͷ�9/�nǟ�w��$I ����?�(�l��́�|1��*Vx*ժ��g?5�{��]+6��k�~�w����/�!��U�o����k���=��D��d\�$m��6g�[H�b溎i����/1Z8�K�Y�E8���"4O��42cw�� �A��P�tf��v�i��ss�<{h�>�m�7^��	6���r���Ƀ���y9����5^��h#�L�9E �[��s����qY���PSn�է�P~Q������3����������ߝ��p{Թ��Qx�����I�,r�t�"�tz��tts���u�TfWZ�;����t�w@|������y���4 ۭ�JHn]mk�$�+s��V�tT���o�wcj��j^t�����ם�ؽ/��"{F��W��:&�`�/��r�9�#����o=teHVP����;��w�����d��{I��Y�T;��[�.�^uw}���op�)-o\����^��/S��w�3����>�GM�=��� �����]�9���w��7§*�^�T}Z�/kZ�Ms�&�z�����=���Gm�n�͵܎xd!�|0�F�@�-{�����;��:�� Δ�e���{u;~��F.e�����=:��q�ޫ�T�m����>�ߔ�������U�[]�ڷ���S�+��Gg�2���T<���k��E��x�l�|Y��#�t���Y��5�����DY��D�T{�C'�Kӕ�����+jJ�RA�Q��� ﯲ��;�TG�^���J��d��>F&�<edq��x����|��ܜ�}ns�,Ld��2Lמ ���
��S����8H��G\��������8��H��TZ���}�O�����{�w<���G`]���l5�U���;>���C���%cJ��/.�"H˗�U��k&��\;Y8%DN/�:�̀�Z�m��S���ڍ�;��ΩL읿�ߏ�Μ���h���JDc�w{.��"��f9s.�=9��o��#�2]�j�8K��D�
�C��J��4�o��ɵ=�g�"�����A����n0�-TN��ܔ纏Fܿ��A��$�0Ll�s�G�X��w��~Db�G�1�M��xO�Zz}�I��=��I�ɱ�Np��"���'�r�`���>kG��v�'��#^L�w��Ck��e��S�b���K���֞�_xh����ǽSzg��^Q��a�������M>� ��U�\9އ�ڋ^۷��y*��{�&�U��Uk�=��{k��(.��#���܊��'��`��k�0��`9ޟC��O.p��Z�|�z�>y�=T;�K��|�þ^9K�����'�cv�P�+�ޫެ�4/l�4��E����r��U����!����S&�q�y�M$�wM珴�8�ٌc���Ǵ�ٺ�\�=���~�7Ǟ�ꇖ�f4r��@⩐Ѯ<4��ڜ�Un�w�+Iםq�B�!��X���9��d<��z퇰#C�Oh���_y�
�-?E�8����BA�.�Ȫ�j��	�t8���Z��ʄ�lW^�.^��q�*�Ԍ�9HY<���J�,��3�u���H�"����VVӳ�z�'o:t�Ϝ�E�]�5���]^���������=����9�0_�9+ݹ��Q���?G�ӵ���'�n�Z�9��F����M��_����uFp���V���ߞ�;�OP���k��Ed��|6YŎq@�����hj�s����\�ቹ깋�t��_7���}��W��Ú"˽h�[g8��Ef���6H��#�,��Ѽ#��<N�7Ƈ�wFx�u崫3��V8�=���P�-���+Nι�9��H�.�|�u�� K�3�>\�Tq˭ȶ��g�e�������\����iy��ҩW{���{�Hk�����{d�̿@�q�9;>����̙l؍���'T�6���r�\u����y�C�i�r��ֽ^��׵}"�|R7�T
gsǠꐑS�����X+N�˪`2��+n^������;�k>�h�u�;[]���p*+�:��'XO�yݘ����Ǒa�D�}5>�R˩���3��wsc!P���Vgu#�&��nU�tZ���	K܉l��<�ǢO}��Pnў`�||=���/K~E�Yt�V�6�k�L���O�z[�ޠ��ql��!�]'=>ng�����۬��ze��"��IӁ�Kށl3a�v6c5x�8|k��w��?��9�y�����9wi�01��_���� �go���S>3=�j��$�֯������d�]VF��}��p��졙��Պ���+\�U���v|�,�#'�\1V�[[�d�j�7��Vm*���v�|��;��c��I�T&���y�嘟$O�@��V4>иg��d��U� �����oZ�v�^��DMol�h���v���.+d�X��w�p$���v�o�����ѿEFȭ��$m��7�ǭ�*l�Y�yF��N�o�h��e�]`Ԧi��3���=�J���ƾ�xx����LJ�n�pJ�G���\�T%ԕ������Yof�{j��d�nqGEy�L����:�]6(D����]xjy�ΒT*Kj���
�a�s���w�	ٸN�)�ˤuj&��Ks��#]j����ޕ�t�X)�R6�N��2^�O9t�֠]�>� �=��K[���~�V�7��	�p�;� ��C�t5�]`1�sxY���L�3Ɔ[�Ǖ�Ut_yuB=�d�W�=�3z\�jT֝�'���CT��}��B�_�b�(�o�7};��y�ּy�z�7��;�4�;d�c�Oh:,�����ѴlalנMgڎ���0F��Gk�����ax�:�4��q�|��q�^EC���uhO�{��Z�۩bW��F�S�<��~��zzg�(�@�]����	+L�f�w.��7����לc��f�	��=A5G�*��W��q��u:ވ]e�g�p����tzZ��o��Pzw����ҟ4�{��ڿ/"���T��#X���?��NįC����,&ǒS�>�~������	�3��ǽpI�:�?��<q��c�~�̸�x)J�3���o�u����Eݲ�����7�.%bp���J爑��:Q��:��]��*�#� t)^������%��nkm��\�8uaB�I�[0N�2'�S/1��(�\1�EULQ��q�X*G�8pr���xJZT�ڜ��ʽ0g��Jx�v���~�emT�2���j
2]q$5�R�HW�,s�&�o�YDש�+��ח�6�}J�8�jx���o�ņT�"'�����9��՗�9�{�,U�D���ٲE�w�J]=k�������t���T������yFn���8��`���Ě6M{�z����,��1&�E�^������|u���.i̊��
�[����CW���y�S.W�k��v��,J�3�=G�3�'*�lә�c�I�*��^��9�ᝄo{ܠ��	�`��ot}�:�Ͻ�����n�lD��؉S�@A���_�d���^�4'�()^.�/��{ޗ�=Lo�?P�X ���'Gq�E��q����u��`��"��
��`�ftY���{�ۥ���}�ޤ&D�ض��[��G��~�)���MȾ�����;M�RĶv�iS��Qֱ��"��CF^��F&<�S��O9�o4C\/*���u�&��#�ԅ��3i�g}���0� =[\`�m�{�wT����࢐�{�==[bͮ�8��+��˖Yj�p��ͅ#m__CMJ���Nu�7�ӴmQ�ܢ��V'Nv^�h�q����]��m��ay`u��D����y5+��f����w8���|C�NzUi�s��
����K�I�!zii�j��O�f���Z����"��׃�z[M��rx��:�p�"���8��xN�#��w�����F7�8��=�o�x�?^v��s��f��� O�����K~@��+�YL�Y��x�����5̕|�mS�<}=��q��i��+�h�#<9�����9/ݣ4�}�X��ܘ�
��>�G�����}�|I<{�=��>�7��VNL��co���:Ǫ�o��gl��C�Y<l��2�L���́��bPO��*Q��⑘����������pO���������i2F:{;A���o����I�л�Ҽ}C��g�Vz�ce������Fz��0rME��r������
��n㔕IY�/
����-S���kv�wȮU�{��3|ƌ+T̚����+�q�p���{j��w�N��ٗ��s闌E��;!RJ�kF�p��j��}�8˨�H���E��ǶҾ�dH�2�%'M�N�~��+�`�c^]R�{�����;Z��s�"�6p�����J�V��TY�юf3��*�߽����u+(�+w�^��׽��y�	��ne�������2�Z*\�c�.<�wk\�<u¹�H�l��W�^U��i����="ζ��cp�\�.5����������'�
���﹝�4�0Ϗ���W���eШ�:zKյ1'��'��\��Ͻ��zmb�x�C7��~s�o������R4��o�w�m*Vb�-��e׾�t>T��u>�ab�p||A9'��q���>�(�Q����o�|�׷��?�ӱާ4S��}�lc���Y��FR'��s��nt�s�<�����tqX=����x}�.,B���ѭ|����t����VWgW�<p��ܟoDv	�A�]���}�z=�����x�x�}��g������7��[�@�6�N�8_=m��8_v�S��N�D�g%���Mc�zb�b}r�8�:�鐻��%���{�����Hdgw�&���;����W��M��AQ�y�9>���sd+����X�TӖ�P7Y6g�â���H��(a��ڑ6�����]ҙ%(��>Y��� 7�ɣ�o^����
"@�ʊ5O�޳#�{ύ�(��7H��vĲzJY>n�7���33�l�O'2r=7�/ ^��K��m�Go��υ��'gsUl�e�؃q�[�rf<�#�Wnh�#g�6X�j�N_m�m�y�SƵd���P[��eFo�ޚ0�+k�mG�`�j�y�颮wl���/�Jx6q��%�������#�-d�x;Rmֵ�[��K����"�U�=��cd�3��	҆JF���������v�{�p{��2Px�,�C�w�ѓ�}a��3t��C� ��g�2��A(	BK������:c��sV>�E���0�9@P���i��%j��ݿ�{�$��F����Wܛ���T<;���{�w���[)��Gb�W�䜱�l�u"�e��F]��+��� ��R`B�3�"F�cd�H��ݺ�7&�ݒ�����A�Y+rJ1\����&"���;}N^���r���[�a��$&c):�f�.���["�Iw��l�ҙ��uo_Ƶc����ͽ�0���h�b�ͮz~[�!�+j+L[
Q�\5��h�q̶jP�%k�S��bP����]��=�Xu���u\&�Z����������K�.�!{G��9�VcB�|�[����N���tjJLz��ז9qӷ��H0���T��ѣ1�UR3ʌ��#d5�h�h�p�cM�<Ȕ.�MJ��ԅ<��o��6�rkD΄q�o5�jj��p���ox)y�k
ʻ �Lml�ۑd*�,���-⍳ճ6��H^e�rn�%|{׽Ĉ�EHͥ�`١m'��{q��Y��Eŝw53WnGq�C�7Ǝ^��z��v2�*c�jcΛ�'U�+���ijba6��i3bm�y�LR8U+�w�j�j�F�]�+8�&N�3t�ɭ����z��[�Å�>9N����$r��>k�;cH����wip��o	ȴ�r�=��ʱ,a��{�C�OP���k �qfG��3!P)eKY��,�34����dJp����]��@�T�%��_o@���6����zU�=)�����ըr��w���jWKxv�gIը�^�wZ�,-������M���9%M�TE�enk��eo$y��A�{0�%z��?]l�A<�ι5M+_U�qG���s`�mgp���C����Z<�aѫ�(İ���h������1��3����Xc*wv�2�b�y �\ZR߬�qq��j��k��.����<�Joe#��h�H��)ׅQ�յ��`�~ �G�|I$�0C��1l%��R�a��C#IH��,�a1�����M�I�(4�B1LR��A�e"�h�ɤ@@i"�a)����D���#���@��B��ۨ�D����s��/uw����\�WCu�ws��(�K���w��w\�;��]����tw] ����.qι����]ut�йn��܇w.�u)v	�ݎ�u��p�Ӕ�p�N�9w8ݳ���wr�n���޺E�;�:컗��qΝ�æN�Ν���7tWwc���\�����re�ݹ9Ӻ�)����qԝ2�uҎ�w�
�nK��s��s�9�()wtI��SJ�����ݒ�C��W�T�-�F��� �㧹�v�;���Z.�e��m������&+���{^�Ug�E�����xSv�zk�N�Q��c���3�X�K�F�p��P�I}��I�αX#��M^N�w��ޝB����{4.he�
H��E�OE����C�sp��@_Iaԕ�B��o&Ӂ���rv����+�������<L���8G4��	��e�����O���fq�rT��vPej-�` ��m�ܞf_5��x���A�ݗ�A���C$Q  ��B��<�ǧ�U����H�"Skz�U�ee+����V����MW�:�Fu��Q4W�l��S���To�#t� ��e���{T^�|�[����C"8'�bY�R�ej�&�Dm�5XF3���$��� �<���E�j>��O��+M�;P��C4H"�}�%:O�"S�P%�{���~vk�<�"��{�0ej��[
���s[{4Yf�B9K7T��3x-e;�ҥ'��NV�"�)��z,�gs��4-;�B��wF�G��0�o�!�pt�bvx7Vt�Q{:�l�n��Xu�� �|	p��]�����h�n۸:�Z�ogQ��rj�{�]��=���Z�� \?��lN�G��Z�~0�����f�ն�,�bi�1��p#kh�F��v����waڊ]q����pl<&��+lZum��n��\���G"�W��8��
�q��c豗�K�nA|��3+�.�:u)n[�d�M��(��%Z�ȫh���!�\�dh��Q�O����q��"Z���$���1.��;C`t�~�D;'�Bz�s����7�A�<�&�ظ�י��Gs�g���}^�1ꐜ�Dc�� ��i��o(;s�X�\�֍ټ�w���w��)>>����,51�e�~���ۓ�^/��r��G��A�x��;��߻�M��5��]���喽Nç�ʄua����s4�YM � TQjO��1j�=1M6���{�[\6�5�gDF���M�10�����KzC��ÝBI�.��e��.a�	Y�ظ�ktt�uS���%ռ�y[I�2��|S^��d�m{���8���]�� |%is�Y��韲]��3g��q�����7���~��Q��1'߃��g������f�����=e�n,���u�k;yЃ&��!��:�Y�l�dgO>�x�`�����?��W5��D�7��������@�t�y�@'�0�z K(ְ@�[�^Qp�ߤ;G�P1���8b5j��*fo�W������N�cY5ív���e�:�(���O��3�%��E��Eé��Щ|D[�6nڣ;�͐'�F�˨��"i���an���������;���=R�"���x�׵^l$u�^=)��l�=��.������mh����j�б�7{���n�vt�=8�HԒPL��tp]l���I.�2�u�ؓ��zy�2Mp0N����#�Zh9o#Y���'j������	�{bS�)P�j�'�Q�B9���oY<��:��-`������_�8>5äLlʅ����i�Re��ɋy7�6]�h�O.��A�5�v{y��Α�:p�;�0��B�G4�r��/Xc�YYR����^OB]Upy��u#�+:m�:�^4�瑶vk��ퟞ\=��&7���_�c�[�x)���dI[�#
�UY��j��Ic^Gi����D����OO�Xx��>��M&F3��m�wm�u���N�'V$�o+�'_%��y��*���>�{A1�@��8o�䡮�y.��ݛ+L�V�b6��
*��͹�E&P�Ƥ� -{*	{k���'�
����OA�v:4�	y�����W����3��G4���l;-��-��XR�B�}�ӏ��A���̦�4�6�S?Ys���,��|�j�W�ނ$�����)�K�#ҷ������>�q�'A��L�>�t6CN��4�%���"�����+�Q&?1 ���|������0~��>�����Q�ƕܼ�^0 �֞�� �+�s�!P��N�k�s��s���c�����ۀ��m	��&u��!1UL؛������� 
SVb8�d����)�|t���{tb	c�g;�����)%e�޻�7[�Gx�⁝��ٳK�|oަ�.�UG�Zd�PdLC`D[*�xc���~�`L�_ã�����E�!^�˓��5���W���vG!�b�5��t�:b���goY�-�.��Y|�����"� �\L]��7��Q�]�0���!s��A���'ATu��E7���Y��'�+q��痬��C����A�Ɯ	�G;J��J��[���D���L�֍xRp4*<u�m�Ki�Ol�]AΌ�+�{�/���*$Q�0�j�D�C�8Hh����@aRZ���7�HL˹-�t�x��U�Q�����l�h]�6�t���
��R�e�]�'�/��bN�]6�B��Xa�;;w��\�s� �K"�9�
cA#I�>��w0����zA�l�D&�tG�4?�K�K�����3D�7ҝ輧L4�s��ܱu;u c��3x6��z`.�^���{tFƾ-1��53�r܄�ʀ�t7�p��qT-mt8-E�沠��R]��'��ɷ�x�M!��z�i���<`0t�cH�ku;4�\��>fj�r��F�G/U��7��o�l:5Z������K3���=����f�S�͌�a�Dޗ�9Z�f�8��n�,ٝ$���K�׾Uu��&���Wf�]P��L�&.�;#"�S��8�|*t����Хw�sj{b2m�z(N�]����Y��=5�S���:轸x;� �s!�G�8u�ѱ,��������R=+\	��̺5]�kv+��-��n��"�Z��]Bv��d.�ØL���'W�#��^�������GF��{|p:���X�l�/������f#�N�'�<�}>���0��Ĉ|�jj����Z7��Ʉ[�M]���=�.��@��_��zK�����C�W�LZ��!��D�ǐr�6x�+dګ��Ps�z�X �x�z&<Ys؞��G8�s>ͬ`��t���&����q�P�޲ՆK�tx)�&-;:F�����D=�O@OE����ٯ�.�5�Xi	]��<׻Vݘ��6�o�df����L���X~0�8y�1��^�S�ʅ��5yrT�����=M	�3;��*;{��Q��:�/�������E�"�Xt@y�a���u�DmEx��ču;�f��Yz�u��x"ݹ��i=�Q�����Օ�VY+F��P5�7A"�;z�D�㷫�:-�!)5�@� �Q1,���	dU#�M�Gc�y�¹Akb�����2{���Y��n�F��̚3!}�����!ݽ�D�ĩ�B�n6�t���gX]��e�֜�٪�����w5a����8��2�P���]bFw�8	��S��ng>��:�_:L��b�	�1*]ڵ:�}�;(�Cy��%~�n#[+h�;5�8���HB}}(�;�t���~�[�F�[ �qͯ�p�/�f:_��7���{�nqn��GC5���f��A���z��wƕ��S���Q�U�9��:���G5�L�w�9���S��`y��l)�4�]M����Y�mEΨ����u�-?'����Ow��jBv�f�]�ts^GR3L"A���1������}G8�FĲ��n��Z����4r_w�5=D],�܎�*��^�ܨ~X����<(��k��W�vOƀ��\�5l�f]��i�O;{hc"�[]���~l�gm�TyLC5⤉��A@x.!��@'��������n�:�3��w�u��t�BՀ�S�1���ȷO�nLW1m����������SE芄,�۽�S:�����r��S�����Ў�0�O�S��M ���PO��0�����kX�&zZ�gL�Ĝ���`H~���qF�ᯌq��6'dk%�!���s�Mq�.�	�b�'�d;{2�nL��1w�C��"��'���a�`x ��o�?ߗ�0�f��d��c��g�j?�s#��S��`�����J�4����Kp��L���/P�0�6tL{��`���Q����m3r��Y��]Inb���P0޻58���W�D��=c:�;��i)G��C6p�RC{�7��[�u;����1��N��}����n��i�$,�w�UU����Y?fԞ�3�HA"�^��v�:߽�֛�����["��HF0��Ƚ���W?���s�h������]���Y�(8���A�Y[$5��=fͲ��l�瞝�0���p�[hv�j[���n��O{���U�0*k(��m�Ђ~ka����Q�g��|jʋ�4.0	c(���3�,����٣P��'�e	D�j���l:.]�c�z�\�2'
�6����d� �=�u�;8��<�۽�<�!T���Dky:�k�K�Nװ���Ҙ��L�ߜħ6J�����h��SUj�Nk�r�^��a �[Gtc{$��q1�C*��bE�i=J�&�y��c7�{�t`�mݺ�5ZǑZ�ǍqӅ�;�0�h��A	֟C�o�= ����od	��l�^3�Gu�n�v[u=�7�m�u��s-灻�vk��\W(VX���܀�^�A�p'R�ɣhou��E�mH���a*��a�-~�Qy�r�ƀGjHO��;!��66��_]o�mz~�s5� �E���Z su�آ���6�N8��E�����?N#�+���+A�u���X�%��(��ꤟ=X6�Z�֩��٬Y�
/s���Y���P-�Nns��v}2�1`d��(r���¯6��+����V<K��`�N�df+yW�]��ˏw(;�c��{nbS
�[.���!l=Z-�G����=?��������BB���!�X:ni�Ƨ�smg�:��:�~��~A/m~������Sgj*���1�=1��csPw��#�΃ls@��思�e��XspG�ߙtݸ�]��3��HY��'�;e�{R�˜Sy6���d"]��t�������'Gz]�������17n��94{�[�ȝv�*����3!h�e]���חx@���^})�7��֢���vڀ�|OGUL�bP]N��쇜��Pi���tE����v{+o�<m���?~�k�:c�WJO~��Ƕ��<���8��VHB�5�\e:j鋇M��t0���K�T�#��=1���#X�8���O~Q�]c*���(_���YB��G\;{�s�lt�>\D�ں��no����=}�L�>͍#�g`��Kg+�کnj~"Sm�d&M�{j|�.�4�F��k.���[Іc��H�Nk�M<5��;@@Ųa>d�HH���|����fu���r�C�1��୭c���P���/D�B�9�k�����&Df��В��s������~]��Z݄�C�r~J��λs(�!j�,��b�����u�W�oe�I��78�d�@U�y0��Z����[BT�ЍҬ�����ظ�2��ѦV�T$�;�ժ������s���i���_5ɴ�,�F���΍��xf�����}�~�e�f�*��(G�+5��3):,�Ⱥ\�Lh�&��+���־�	��8���i�o�[o��kP�WSG��A��"U�N�f):a�aHs�1��̎ys>�j��Y���t���o[��vC0L�a�ZD!�:c�n�;JUzʮ��Qi���T�(�C�\Ol��i��Q�y�
p��<��ͭ0�kuN�'V$ת��ԔP�uz���s/�����^u�A?�5���n��f=y=�x�����tz�Z�ڣ��2B�o��V	m�嗭Io���b@t~?�^׸��3:�M���M&�"8��k���v�p:y��IL���j����m�[����Ṷ<u>��>�z��j;r�K�gc��;G�p��
�m��yd�+�Er2(�{�8���]˕���7ҋ���IC�D�m��*�¼xE��6�(tK�b��sٯO�QSZ�m`�-��f�g>OFs��C��X�K�0�t��5P���-Ƿ��ٔ�KΫ�x��]d=+�g�ZZB���|��ǳ��9�p�4ﯤ��J� �^���岭)�x^�-�뜺��{���O����С�9
�:��s�x����]v-Y�@I��✸d���ގ� �X�1��>���|�5r;��4��<��͉�w��T�ms�QHJ���%�n�'Yfj���t�to]�����ޱ՚�FC]8����g}�<=���v�d��u��p���_����L_��x~�R�ʟN.�m�_�����0c��ʸ鳓V�	g)k2q�jNPz͜OC��WL��	j���ǧ�U�Gmg4C�۷�v�̹�=����|�H�ڌ Ɋ�4�����馞�;�
N��-����0���-m!�:��VJ�j�qDĲ.R�daS�i�"7[����=������l���s���N�f�g�_	O���s��V��34��-�4���ry��0uGWM��B�U#ϴ���8����`�fڝ����"̧p�TJN]�?�"��m��n�=L�ih��;9KdE�l>�a^q<�1���Cw鶢������$?s�L��"6f��� �Aqy��bXA��F02Y��i�s��_���r�q��Yv;N����~�ͩ��?c�'+��0�]�ظ~X���/�aC`w���������T+�����j�+P��L���Vi����#&�eG�T�6Pطvm�`�~`�����z��^�o�����}��/!��q�D�a�2�~ �a�h�w�J��̀჋Kj�L�;9Ǩ'z�uׇt�q+��D�;d�s�t�'Tհݩ�F�,��"�`�F��8��Jj�[�ٿ	�2�u��!�Hrם�7���̮�֨�#�����i��ù�^P=E��f�fI�X�[Dk�m�h�0���1�G�MXq�1�d����C#�L�bӇ���m��;��f�/]я�j�C+Fnt-`�Ņ�����܃)󵼟֔�At���k��W�oܶ�-Q�[¹YJz�2r�z�I����;$zmN�\�~��ù���VES�5��N����,�z8�@���s��1N�Ǭ��0kҦ���M��7�f�jŲnn�&�3wC7�q��eǭ�H�8�,��3`���EW�q�AQ3�H)�#��ق��;�Dc���g���#	����^1|��2�U�������Q�s����"� �A*[o����z gJ� �k�����lJ�����(5����"�>m�+9���n���s�ar�-��i\�^�;PF�pQ������o(��� Xp]5�Z�삤T"���S��S���l�f�Yҵv��W8���P���v&�T��;�]d2t�\d{����SI�#V8sכ�:�r屬%ry�g:=gF��p��C��2�A�h�/�+sz�7s
���3t�3���2v�WM�˥��v�#H�����;�֋��*���N�I��=��v�(>��<�ko	�- ��2��õ�ځ����y����/|Op�~�+���W�����N~�t�P++tqs[c�u�1s�Q�V���`���E;-��w5��Y�U�޳ō�}�qM��-���L�wD�e��CM(���E=^���@�2uQ;��yv�^�8򄭵5�;��j�棽�+7 h�ՙJ�"E3M%����2�V��&�/���)���U�U�B�,�ئ��D��9r_b��Y�nw]���6��"R�:{1�����5J�]wmڢ$y]���srV�������ʲ释������b;�J��h��|��K�}FI�!/WU�f���l���5e���Q���#��_C6�:�*<{#A_D ���e�	}��1��tD�=�ua8����Z�'9"�Y����r�k޶F�\��Z�HLsgT=�Jw^sʉ,|�p�RN������[�v��[	�<;"�*�'e�C-�3)QY�4�aǕ��]��f��Ū��^�BZ<��A�������B1�I����
|E5�;�ݛ���WW���;*]����Q����ƓT��M0���oݼ0�e9ϮA]��{pr0˖kl-�`d�4Fq_�`�c�P6��nF��5�E��t�V��Lι��`�D[��A���f�Aeq,�]�37l�/U�A���1,;7Y��:șȪ�NZ�qkj��{tAL��DE5
���D|~$�I�$��I.���%x�+�tb ��t��Ls�CI41�RCt��.��tM1'9���!#D	̉���M�IfIHd�"��hY2��&�w&4X�����Kݹ@I�Q&����:j�D�F1#fm	I�Q
k��PA���E$(��l��n[��� {u^��$�(�2dѬ�Pd��4�hؙ��HcA���M4Pd��6(��X���	I��%�&�ɑ,�H��|n���~g��_I)�g��.g�ƃ�*w�o�Y�}*ov�ux����D�Y�.���v��z�t9֛ocS���;�j>�{���'�zK��iP�0% 03&!� �]�WI�*���Ր;gHlD��;X���t���R�R�p/���]>��&+���g��;r�l\`�M�2�vS�Mژ7�t8Bb�!�ax�t��Ƅsaq)8%9�`�4�
�-&��y
i�����&xA-�ļ��{�Y��,��`�ìs��5�ސ��odI�4]�������D��ۘ#+���52�z���_�r���`�?�^�$d��):����s����T�0�����{��4���(�A�q3m�]���+�w�<�_�/��?����Q��2�T�U�-�W�q-�֣��q@� ū�d���� ��6ʲ���sӽ��#��1Ԧ�Z�w+r��A��C�z`�k(#��m�zOͅ�NV@�4Q�g/���/P�q��?5ɩ+�����fD(��q��5��nu�VL.z�e���tV���a,b�cN�5���2�g�5�[!u�\c<H�o@�A�k�%�'j��nИ���L�ߜħ1b��K�0�QZ����C�eV��í�p���H"1��.6eW��CM�`+˯L�{ߢ�e�Uo{�a(v�'�7Nc깉��YQPe
���yV)��z_%������Xw^�G���̹�c�d���IL���]r�<��Z�KV��-�m]�����sŢ�im���y�*Ǹ�<8�8�H�aP�Ɣ����� <*h�mΨ;��kg�ׁ�U��y�:\d#�Ӿ[�	2y#a�O��.�l�0oQr�mE����HS�P��5)<���X^4�瑴�s�w�8e��H�F�bBz]��juhoc�ח���4�N�c��jQ��
�2����/7⤱�v����wf�vC�Ѥ��$Vy���"�4��lP�LG�d���W:�R(�8��qTXU��c7J�������4%�&�v�d�,�Nc�����X?74�P�ק�snq�K�J�a?J�)�ze|'�n�;5�Q2�X�r����{�L�<̆�5@|NhN˲�΢Ú��@���o��+���5���yYu��z��0��L磾���w#={D&�o�=9.�:�W�F5C	&���dVƖ�7�^�5�(]�q�nǡ�f|tE��b��L~bhY�nR���w�]V��z�'���r��voD<��	E@A�0���U�6��\3JS�t�؍�{�C�N�ld���!{�"�^fR/�Q��ٮu� ����+$!^D�����S�� ޏqY�7L���av+]ǩ�	���(㶥p�W�6m�|8\t�ᤆ���`�������L�����-xR�nz�ڽ�A�����}1z���*T��	D��{��|f�72�;Y=*�%�nuثFQk�S����l�NHsi�T,�)v,��8�W���ӱ��>��< �g����I,�C�9/,�y,,1N.-�h��F5u�T�5.R=��Z�K;T��2}�/*)���%��`�b���goGM�8&H����2W�R���Bl;��D�U�v�F���!����C����;�fY���f!8,��k��&Dfѹv�D>�׻����ʇ<J~��S��%P��d�=oz;^S�>����c�? ��fil<�-�=bm��R��p@3|��4̤�Ĳ.�=�4�#*�0hv7�S��'��қNh*�>�6��i�]���^��a!h�I�E���)�] 9���v�:��WR��uz��K�d����>ߐ~u�lBvmkDsuzzBcXn�iC��YU��j-?5���r�Iq�n;�(�ˇ�~�}RӖ\����Iĸs�|�����~��'f��1LY7"}DqVa�ٱ}�15�q?���J��L��Gw����(�� ?v�q�[����ֿW�f�U���{e8�����xݾ��w�7yc
͍�E?y\V+��댝�D.�
��0���(:�7儑�P/����	�s�Hf����R�e��s]ۏ9�n4se4��Y�}b-u#���o9����W{�Fr�
���*�k$� �)T���-���Mtv��[h�)N�!u��xpJ�{b����)�o�$�!
T��
�ӔL7�xJ��Lc�{> x4X�$��Nٯ��M��Kqg�{�r�N��m�ۖc@ņv%�5p0�t�I<�e.3����wh.q����lB�I~,��G��C�W���-��C��O��Bg5
j:sf�3� 洆�.�X"k���O����q����
=1AH=$ p�MC5��b�Jѱj�e7v\jq/�w�{C�Y�!�������<sս�9�p�4����>�;y1������/lq��_���7�_�r����L�?�����R��*}����h����ֻ�
u���r/�i�A�Z�`Z�9A�6q>4��ΑN�Ŵ�ȋ�O�F��5&�N�tv�S�,/*��!6o��5,3K}���E�1x�-��5����(u�D4d�즊�yT��p.a���H<�͐�B�m��W��d{)�V�I��6���;cEu䉗IA�3�}�67��;�B��Ivl�/	�����GDJt�D�65H�4���̷u�yӋN�B6O[�V�{[2s��y�H�fƟBR��'��T0�0R,�w4Ҥ���r����y$|�{���˂�6��.>�ne�t���7c�+Cz�����Ώ�E�
�w�Γԇ��yr�`~�	���g^��u�\)���¬��%�n�yn�\�N�N�VzŶ��Nv��ˋ�De<�"i�'%��ŒNѧ�W9�i�[&���ū�j`�P���|+b~�w����ĕC�{4�[�z,�>G�d0�a#��	��g�u{:m����m{�5���G;��'9�t�^�I��qyK��D���>a��?5Ñ�5��:;M�/E�/h^�s�V�b�Mk]�^+֤k�ߟr�q!���9�D?�X�]�;�}�"�����+;+0�l~�=B��L�e^�j��L��׈ɷ��>�S,ٯN�ۛ�����Xat���N�l�Z���z�����q�j�Ja�ƲǾ]>��I��BS��%�X9���{�]���Ýa;j�Cq��<!�r�!���	�v�m�dGvI����0E4�n����w;O\Z�sz��
[[>�Oa�G;)��8��������lM�O�����@ÝBcl�q=5v����4��SN�2I���=�ߕr���l&?z-�LL$�:-���g;�l�Uus�:cb7\ �ƙ���� T� �36�֞�<����N���B1�^M�3,��-�}��=�j��К��͊֯-���!-Ed��Fu�6)�� [:~iw ���<3��?~��|H�6���ځ�r�-���TA �Z2�љ�����X��\�-P"�`���3Jʍ!yI�u���7���1X)�`��h��eo��xP��{3i�H�M����Yr`�nM\h#ܥŌo�x��W-{����M=�����w�M��{���.�;��'�w��!v�y`�k(%��m��'�Xa�@�4Q�g�u�4�^�w����V�^�z��T9J3�����\eLO;H]:ɲs��k�F):���$�I��[CTX�M=����1�5Yh�0G���~^�"��2m�� .)0���)�r��ܣ�d5�6��2�y�+��.)6�{"�F7�A��p��2�},�6�|w���D�mRP�;w����̋8LV�	/Ż�3xK�K��O:F��B>s��W3ΫXڻbu�z�=.��݁,hOc�r�fy�zm�u�/�}��6��s�s?> ��X�z�J��w��k��m]:��آ�H���I�U�\���W(�ߊ�Ƽ��0�������[#Q��	�{�O΃��2��t������W:�R(��n(���­t��)V���T6���g�OUg2�S��{p���:�e��sL	�OH���4-[�X�?Jק�I�-�˟2�4���|d'cy�A��e�;�"<��Cc�D���̨}u.��cXy��4!W_��/������yٮ������B���d�~͖wO.����V�b�d�S�-H�
Wz/(�(��v`C���zm�;��t0�Dt��m�ѡ��ӗn���gL��eA�7���<��Sl�)(/���\�Љ�*�������������Ӆ���R��:�ϛnk�v��5-�G����{�L�y�H�`<�C�]�b��c�VQ3/�n���m.R�vR0���\e۱�Ì�0{C��B���5D�߇��?:d[�Q��Q�׽:�y.�Te�2���,c�b:�$=D�1��ˇD��k����|@ͤa��f@��2GzQqQ�+���Ƕ��\��	����r�����CF�txd�4c�����_`8���
g�XE�)Ĉ��/~��j�ʩlj��!s���A�6�\d��r��Z5����H�Ww�b��7��X��yL�:ll�G;O��2W��w�I3�S�S��x�v'�x�r��]*;B�ǧ5���V��=��x b�S�!�$/�����3d_uwG\��+3�]L���Js`�LPRU|����xOMn�$8X�b�_\�sͭ�ݶ�=�x'��	�W�L�	:,�ȺC�)� ����׬������Wl�9��oY�w;P��#�S":�}�w<s��ȁ٤�e�:a��Qu��Lqt�sz��:������c���-q��3m�������I7���А��]-]�Z���8�t령����.�l�e�����P�2�al�[������ �Ե0�k#Jh����ʵ���w7�h$շ�P�,�$�y�v	�%��x���"�q\Mh�:�R���}_��W�Qj��Z�j�UV�����H�h��O/��w���B��Bn�=!1�R$��$�U��j-?4�,�D�B��mf����u����<rv����~�ψs/�L�����^_�z[�0��s�{b�Ղ�9���8�e�_�̡F�s�q\����`8��s�Pp�_�N�6��ݥ|�"����[}b�b�aEZ�T�/b�s�f����Wa1�戮�+=�~�Vн��Z��3�6?2�t;$�/�m��)�	�e��>�����m�}�@���ξ�g�$�/�v�^
!�9�BK�=��t�C6C�ϯ����!�qh�8�zA�ůM�J��=D�M�hǚ����P���{C�A�O�T�{���Y�q��#6����a �`䆖��Ʀ���E�;ҡ�>�J��uY�����-���|���y��7<��^��\�豆�uc4�wv�����P"�L�p��ʾ�-3�S�����/ �� �z��Ou9�k�$u��n~v�zY�x�ʭN0-^H������O �_70!�+��\���5^~�A������7�9H,>���3z.4�,�嵌r��gw���� ⊷�Y���� ;��f0�wq���V�7O�\�d�����bZ��h��4����7�6���H:�ubWM��,ץmt�{�i1Cv2u���2֓��ӗ���������Z�Ƶ�����?��5��ﺊ�i�raԒO�?O�����cj+�r�mA�P�{�TgXW��0�\+��8H�|� =���p�$/-�q٣P��%����(<�vl�+%W2񈀜i1,�ߊSL�ʕ&���|k[]���ī^��=��>�g�F=>2O��N͕�xL_	M_8�^��Jt�/M;��S<nC��3T͍�7��w5�\ke�ܒ͏M�nΏ?�f��	K6���e���h�)�N�T�����J�}��KJ�]s�ˡW���h��ǘsP]]����"�BG��D&ڝ���M%�Pc��*E��G=Uz��y;#p[���b���'�K����]4�$��������qJ����İ�ɗ���˙Cv�]D�Y�Z�c��^�#O��~}ʿ,Ht�9�|��C���Ҹ�Ǩغ`��<�K���}
�סغ���
.�I�Lk�M[^�I��#&�lR�G�L�el[�6���p�[S����Y�xf&�C���ٓ��'���8ȥΥ0�c��G�:LW2�/���W1�a��|���&�.,�D&Ƒ���v�0�n�Ў���pl'3Ly����o6�)��p�<=ݷE푊v0���V��{$��׳��-S,Y��<���Y�7��ѱp���F,ػE��5�G}x1����n�ChN>�چ昵N����՜���1��r��/h�Xm�C�����0u�~��{��__?~߆��%��6�ֱ����­��.�C/�^�s�N��q���4G3�
LL,s~�������~~,�p����Ox�dhf��wv���G��B|g���>��}1*�-?V��CF��g�Iи]��a�z���Ҽ<�U*�K���yf����<�TS ��L�M����y��]�(\<�0&cyQ�8-�J��z^zޗޭ
� ��=�\���lV��(8����CW�3��3f�c�gN��N����5�w*}���l�!'������PJ��������0�	��d	cE�w�۸�4��0ݶk:��m�G���Z.Ȉ�h�.�ZCEa��q�p�_]�c���N�{��˹�R�q�7u��!�s8�Y��k댇V�ςDkz�,�R��f�7Ҙ�V�����Xf��j�\�>F?R�E��ȝ~��Je'ѳl$vE�*8ށ �ƟC�Hق^Q���|���;7v}�2�÷�k�L����h�	q�lGNf�xa��:E�W0v�Rl�I��$��Υ��T����ʖmCH�R���d]g��搷�F׎�sӿ3��y��W��������}��o�����A�k�z���1��'"5���S�A���	E�Ià�8*ͥY��0�K�UB�=���f�z%�eb���M���M2B�Kޮ9���Q�\]c�}�βZ�5�9Q>�R��"}ʈ�|+�״K�kF�r\����N�W0%��x�n�f�p��&�Wt�xΎGJ����p�Ղ�Nk����6�u]I��:�F��Q=��z��y�)K�m�:�`�6��Mv����3kl�r���8����C�֡�1��"���;�T��Ln�s�e:��K�X��Р.�m�s�E���ˊ�h|���c[�+��7J��h���h�G�Ê�몸�)�CF��&��l��7�=���cY ���g�$�� �]}G{���S��Z���z
��u��;��'Lĝ1�twR���.�t'=lĳ�w]@4(G��K6ۻ		gTiA'���^�f]�A-v:��a̕�,n�U
 ��C�+2k��m��E;��L�rNDW+���M9
��z�xV�(Yڗ��F�m�7^lFq/�4Ŧ�m�O!�N�*�fv�9P7y2�u�|�f��S�p��x	�Mu{���aN4���:�.ʹ:��.�p�wtw����ty�fF�Pٹ%��C��6B��]-b�楋�5�+�����гyӇ,j�㣱ZfR:�)���E��Wu�:����-k�z�N}n$;�"&��6�;y���̳��|,V�6�^��:I��e��ԔS$oM�]�^^���X�3��W~��>~����Ri�1f�v��0?��D��Z/*W*y����������
�W�2�tC�;}�]I�WY6�jzWb�Չ/�[p������2�}Z]���@�M!l���[�6^��YFMTXu���C�S���@g6���v��:Ő(m9����f�JGDJ��\4�s����3�W���w�{�S��b��O``��&�;���_Y6w�y����ML�ܫ�9�B�q��Tv鞟P�������}���t}2Y+��Q��h��6Ǧ����I!�>�S�_t\��-�����M��0eY����#��^^e�)�o�fC�Q��!��2����w���PXmsɛ5�ئ��Q�[gd��w��5�0A�Bҽj�[z�-ggi�{q��5�}���}Ok�;�ƺ��T�L�7f⒲\e;$bU�˧g&mY��맓JP�ڣ˭)���n�r���*.r�"���{�f.���BT�K�[�M=޸��C=�'�N<k>e�M"�i����Q��!�m��[��`
�oE97�j���V<`�9��d�Ip�ݝN<q)��z�9��p|&�IV�gC[�n�S2�ĳ4=���n���Ti(F.��kQv�S�Kz�`�T�㜡��o늤BW^�HP7<Ўo|9Q[���z�г,�B��oj��o�7%���er ���o^���KE�F4Ph�C#%2"�"+�E��TccRT�&��\�!(�cE\�	�l-a�dQ��	0P4�M252��+��2csj�b��I4h��A�m��cPIP\�(��Ӗ,D��b�E��I�Ё�"4g@�!���HKEI�,�!�QF��Q��b�d�HU͹E3;�TVJ�D[���`�5�s�G4� 2��Q;��&��Zf.j� H���h4nr�sn��F��sT\�ݸ���N��ۉPQC�����d�b����ښffک�i�;�Y5d��GD�f���׫�������X�r¦���*ɇZ;�ej�}�>��=�w�ߎmm�j����V���m�����?>;����/����~[ˣ�0�1�=��lA�o&B̮xj���^l%�;0òZ�f�e�������"v�����F���U9�/�гa̜qv=�QaB�O1�N#emz�;�F�!����k\�,���>�`�����k�T	�xI�[k
��b��V�2��ɛ����73oɶYn���:	{k�})8��Ũ;���'���69���sS���*xdk�ݜ��������.��]o�ݢ��R��1~U�`�y��p�	��yݥ��Ձ��D�܎8��:�|Bz]�u`oK�N�C�瑯���C�#3��P�,�)�.�z�ۑ�-ga	v�z-V4J.�	��GG���`ާa�,��= ��T��'������]���{�=�L��hD�!24+dHM��&�����\���ycn�?�B��C�L�3]MQ���Rч\�B�!�����Ú�|XU�IďE��x�ƞ��km���g[wD-���ͼ�hByg)k3(Q�MAV�� ��j�_߃�p����|����H��*�8��Z��ɬ�US.:l���$���Tz.�d��m��v��+xѝ���ndz����3Q{(��Oq�Ps����z�4��KɆ��� �80�k�p��WR^J��ʂ-�W�����,�&rIs�*Y������{�}�~Z��Uj5�b��U&ՠ�b�j�m������Q�e=��--���ld&T�£�,�^>��V��)흕3�q$>dQ둰�	�y�n?_m!�fϸ2�O5t!)�g�犔�5yIT.�&���_q�=|w����n*��I9������f�vgC%ס��g'��|k�4̤�x�E��Ƽ�����,����:S;��M�Q�͍ �5�D���ƽ�H�fS�يN�r�E��)��C�����v6=�,o�;Y}��^w��8(f�PDCv=!1�a��/���𲫡�/=�-uF�ht3�j�|e��L�t�~d�=��� 0�����kZ�\1����pW�n�N�z/�����K{2nv;�w���bZ��е�fvFa���^6AC:�@�0��I�{�?���~�	��褼>�O���9Sl5��~*	{��J9��K6������8wM�A�\��g�՚�½u�v.�Dgza���d�+��1L�/{��}:�8��W�ܳ,3��#j���V%]%����̈�"y���^��:~��!�d_J/�Ǥ��-���x���!b��ߛ��E$E���n��p<:��S>s���8@�P4��]_dpӖ���w���?������W�v�B�Es,� 29�Mz�'�d��z��S:c<�d�}:P���*�Mv8%�W4���-�m��ܯ�ufRW���koŴm�mjJƨ�Eh��T�+h�ض�������NtY����T�x'+ `�gO������	��z.$D������t��rsk)zF��u�9�=v��NF;�|���i��o���T?VD�ǁZZB��'�=�g=�C�d�f��a�\�j*/2��DA�=�i�z�a�tFAoג�*�-3>�
v"G����d�s�yGDk�M�}�-����W��8�JT��vPeA�N0-a#���8�h�y"�Lqy7܀���toKZ���glcV]���@*�`����O���ڌ ɏ�)��Lc��x���;P�v\H7m���{����n��\���*d"�`�*��tB	�/��Ji��T�Օ�Mvެ���5==��Ξi��Aq��.͕`��&y�A,�/�}��xO�$�=����E��#�܇5!��Z���_"��ty���	K6Н��2���q��!�v�S���y�f糗s�tE՜�(�*����e���<����G��M�;<��*xM35\�i�(~ͥ-e�i�ia7C׹E�����Ժi�O�H~��
9�����n]��Uܝ�6\�tD�c�K���?1�,f.+��/o��1Y�F��`XK��92��M���+~M~�_nݩ�%di�u8ΒW!��!���vz���7�Ӵ
ImN�*f��Y%Íٚ�m�����bq}݊u�c6\�rw&﫴+��L}�W⪍h����Z6����F��-�ɢ��<�<<�&��dMe⥃�}�=�=sL��ʵ��E‵#XÁ@��z	bC��9�D_���r^��.���(�A��y�d�P��\��&E1��o3öR~k��d�͊Y��m�ס�I/6�*�wg����ܲ3��!%����z�����"�:�Á}eo��}��Z�'��(BՏ�բ�6T����4!Β��?3��^9{�=ѝD�.F����\M�4����T���TQd�)�i{�9�4G3�`PZDL,sbvF�\Z��]�_(��b�NƖ��9|���>�wj �f->&:E��'��"O��^�|_�fyvٹ̨���+���SϪvq����>��,�z;�2D�4�}kO\�o����M���l����|Ŭk�pj�����ߦ�}�3bq�d$PY1j�Y$5��=�6��{N���.�E�u��l��K�#�ُ, �YA,��V5�'�����,z_��w�fnuJ��F4v�"Ό+|j�_�^��38�Ϩ`��@LO;J��MY0��tB������^���{��S)�_�pYb�"��TC3�����/4p�~����֞{�p�Bl{UV�<���V���hZ8o�)rn١���S���j�*��ꛣR���r�Hi_�׽�����<��$�n@�RqT9[S8����ݵ��ޝ����5��>`��`=��o{��Qm$Tf�Q���m��L�m�6+^M�E�zX��e���B��U �S-���z�]�g�弜�5`�����:Y�ɺ�[����������ZYlF�OnbS�*�*��]�ٶ�MN7�A�" �b���"�	�����1Y��CO���H�I�����I�� �8^�K-2&�bO���GEu�/٧z�XR��~�N�!9��A�P�f�'�f�Y��9�ع�i؞sqfNIx��Q;1)�95ϫ�Ӈ���k�9���=�ߤ�
7�����o����^l�,F�Тv�tY�V��Sz�0A<;���Xw�������T':��箅��oB��2ʾae�`,T�9�V�þպ�Cr\��+������� A��;㧛= �cS�9����T������L۽[��;�j|�G\b���%���*p��s��$�`�y���G4�|Ng0�%�^ֻ���]���v�Xs,)P6.�Ǳ��(5-�@�/EX+��� )>ax���Ȼ���<�[�ׁ[�)�������v��G��^�.ݏ^�3�Ap�eF��>oQ�g#4�?[��j՘ݶѱ���.r	)۔;��&V��_jÙa<�CG)C`�痶����� 2��'k@�~�Ep�D#��B���gN/�r�����d���@�۽Vڐ =G�{�O��z#*�}z3���\ �_Ǯ���}�~V���-�-F�ثf����^�>}�5q
�;�!�<��2�טyO�(ۜbsz��z�,��= ��8A�"f���M�f3�>u�9�����xl.�d\>d$�&���]k�l$Z�r/����'U�k���d��q��0-F��*.gC�֢>u\�+��R��ƥ)-��|i�*���]�d"�LNE��gn�����3`�Uk(Q�
����6�sרk����p�0G����/�Xʸ��ݥӹ&陆�NP��h�L����vGNk�M<5��O��/-SӲv�.+R����#�>/L����|��z�ȳ�s�J`����]�M�׵���E��]�;MnX�+�qc�!�cϡ���O\�,*�@r���<^%�u��LR2�^��1J{J�n=�Q��YN��Nxy����6LB`��zcXD�Ve;��0�ʥ[.��[K�ˉ�iA�F���hY�v�1��;�׏8zh(fƑ!7P�����t(�;JS��Ri�"K�˫��ۜ�^E'��C���~�1��a��'��x���a�w�6����{o������,��'���`k'\L��͈���-]e���v׊��l����Lsq�>�	�@�J�u�{�]zd��«S���Kc��rݿt���Of�7��{uʑ����Օ8�n`��VҦk��ۋ�	R�ZM��9��AzgHy���AxGsm������+� �(��m�mL�h��_P[����R~ڨǆ��e[�x�e�*�=Q��lR�祐/��ۇ���в�@��rN�5��ħ]��^Ko(,��'��+h���J��=�PK�V+��댝�vB�:	�d/�ϥz��{�ӂ�-���kF��^a�:i��mǫޛcb
��3����>�z�3�v����j�������^3���>���N���r^�<��{����l��o���x���Šv�j�������qJ�"���8��xE�eAݷ:%�X@��\<(��'c5��-�g6���S���"miQ��%�7�L�t3$q5%�[�]��"Y�r����Agkd�==�~��{'�N��>�z�"=o�u�sn�k�7ި<?~��AK��I��
vd��Oi�*��cL&/����f��&=��g
B.�������[�
9A�6m={��WH�}���D�d�����hBYhs�1q�"�V0J����!6#1e�i=�Fu���͒��V��3]f�g�|��g�������'�r9�X"X,�&BA�6m��n�qCK"�R�d�J��2�]�g�c2pJ�~����*~��sU�#T(n�������,��kzf=�)��Y�$�AY�B���]���!�⧽�ޙ���"�xX�������X��Vg^���΄I��T$�*	�;�-Fj�W@p6�[Kt%�*����i�SS�n����>���_'�oŨ��Jљl���7�눵<Y_A-��ơ�l��On��
J�.͕�xL_	_A/��l���-4Y=]s�X�`�����,��^(�kgێf��u�q �5��Rʹ'g�*��,�>6"�SL<fE_U��l+��a�u����Rr�sȣ^�\Ú���#ϲ�-��@s>iM��^˩�ں�@��f�,�b�l�Q{�]��&�z�(���'�Kח���i�H=!�@h�L��3R��eY(��F�͢2����W��Ȧ���|g��tzZ�O���ܻ��>��lx��S�;����V��6y�=���OP�u~�"��V����WI�f���z"��F�b�(�t�E�o|�u�z!3w�E��}?C���|��wf�E����Ȥ�Jj���;�����.�{?=�)"���������	�������u�Nd���0�ŝ���	�t��dG�L�*�Kj�^�Z3ܻ\Z�٦3��/:_��4�����zp~^6�yM��X�U;tNfD_g-�CX��t�x�oX��GG�	��懧����?v�����ؠ���R'���X57-�by�<���3�1�︢���*�ۻ�es!#w�gVvZQ5����������}�87�0� �Hz���A��%��׈�AȊ�4��b7h:���Y�wJR}��$`�8�q�4���Pn8E�篧� ~#����O�oxo ��a���xި�K������m�f�� ��L�@��v���D�6��Z��<���x̃�5X�hE���"�#`I�����'����f�kW��A���*��+��i�<YҦ����76Kf��*�[><���`�ˬ`�S�>��
��߲���:	�� �3�e�@,����^|5x�=F��l��6 ��8=��qub$�ʉa-�Һu�d:�'�L�%M�7l�I�g8D3�^�\���B��T�SP[s�C�.U�3ǤAoB�,�B^v�dک�ژv���9vb�U�u�f!y\��.�v/	�x�BҙI�tl�'c��WL?8=>3C��<�6�)��wqq���Y��&e{�6�)v��J�"��y�K�~��.͔��\P�_]#�&�;5�gp�����?P���z;YP8��¯(�gk����,u��*��!�#�������t����� ���z��NnMУxi0�0����//�p;�r���VY�pG��߸g��hW�I�؎C�:n������\�ě�e�q_�={�b��rm5��5��h�<�g;��+�(�X�,{S8��Y��U�	�.�A2��wov?�Z���z;��A��/x2&�����(�}>����"��_wMd�l�#�yw�-�v����8������й��ۓz�`P8�����.&��֒�ّF������ﾫ�����f�W��I��waY����ZD��OA^�AC�i�Z@�i�tm�w0�� ���_G��CJ|���?JװT��%G0��:�9�:�@�����ᯋ蟞<��Wi�?]_Vdv�v���_�v[@a�Ú�L���z���ܡ�s��y�����Pg8H�{t�3�A�M,��t�7�5��u��@x�o���vE��;wa�,+�Iv��G�W���������׈]o��fU�F��̾�2f::1	�	ᐌ�lj1���v�d<����X*{��e��h���!��?TgJޅ����L��X��!24+�����f�5�^A!��K\�T���5�x�^4�)��$^$ך�%�`鋇U�g�X$��0:N&.���cQ�#��p�;�дA��E���ᐹ��aUk(Q���CzY�k׮�~�|���O�(WTG;����nf���`�we�8�^�KsS��m����I�*;B���{���7%a��6u��+zM�k�ݸ�"P|���y�QͽJ:�^)9�T��L������^�����|�}��o�����}��/w��m�p4J�l��9j�I��!�&䢏u'ۮTR�]�oW��)gWLN]}����4�p�؂��1Y�@�8�=�Wr��4��"�p����ʼ�ڻM���cCi�3pN)�ѻ�U/??{��g-��]����957��O%��l�P���ὓB�����N����S��-���C��������4�v[����۶�V0���w;n��"I�I���nm��;wQ������6q9r4x_02�w��ʛ�x�Km�̻��6��_:�4im����,r�]�|2�pWk�飓�]nm�ڹ����[I�X�kZLu�h��I3>9�.�n��isu�O�]:+���9��c�y��gr�-����y.�R��ܹ����Lr$��zE:Ż�F;y�'h8�S6cK�l�
ȦE(6�^�[��,�J��d�����x.���j4�cn䕕7
ړ
�hw[��t;
�d����:M����n�S�����ʳ	�'�փODK�B�]M@1�k�z̓���E�+��K{u.�,�g=�=���:��Y�Դ� I��=Uǜ�1a�L]�EVFx�(�P�S�L��َ�/j�C�oY���1,�ݺ�1P�yq�'_1t�{�p�ځ_B
㊀Tt�kP&��3��7�:|�f�d��#�S~��z��2�(�,.��{�X��n�d|k�3D^b�x��ki��/#���c���s*.fl�F�d,�BpTȲ3��P)�C����	GWݸ����o���gX�돦ltoe`}ݜ�Tz�g��kV���T{4<��� T�x����pQg
�Z���a����Z]2n9P�նm;����/k��ݕ1��B�*TY���+X
��B�˘Yǃ��J���R����DذjǹwO5��,F*���˓v��9!{��d[ �j+q���!��i�;M5�Pf����A�Z�n��(2e������2󡬍���خ�#�3%i긶�H̍�'�W���].ټѹ�M���ӂ�2���'!�v�.4#@:��:œ,X�,ټE�O�
쳝6�e�2/��,�H�Z���U/+�`-����Y˖�*;H>R�J�*���b��Z��"�bmic�F���;UL쿜��ؗ�WPls6��L����>"Y˾���Z:���*M�cf���'J$	Jm��4'iV��p���l�d[���3��py�;B6s&��ַ�㫷ٵ��u�U	t}GrK���h�:����{��{)��Xw�ufWU�4���p�n�6�WV���y-Nȷ�L�ن�m	�!���`o(���n(.�@�Fګu�W��_e,Y��KD̔�!X���`�]^;[vLA<�]&`�U)-�)�&��t�u�^�+�>�����Nˡ��� �S�f�����E���r�:u|��qre+���{z�ׯ^��]{{w��_}�HHca-E��+2"(5���t��7I�ݣAhƍFѰX1i&lb�ZH����زc�ڋ��Dت�F���3IF
�6�j1&#b�Pb��KIb�c5(�J�F�+7l#h6�Q�\�(�ۖܶ�,j�������F6J�6"�X�b��Bj"�1%N�q*"��Q	m�j-&ɮk���i��Y(�lX����F�&����"�cF��6�A��l�") ��,UE@'�}�}xqZ����ֽ�@ܺܤ^K8@�m@>jZs��ԓi�z>ȶa���Vvb�%b������	vs�wfo&��Vd��aԈ��e�ˈ�!��� �+�U	�"��8�f�!�<V-�'(>P��B{����5�L�N��K"�<S��ke۬����F�s4w\-`��\P{��}ml�a�&!0\�'��8D[�m;ױEc�+_Z0�%�X���Zt�{�~(o�0�?/B.xM:�:�AQc�������:�՞�l�:XR-9�TUf6����8� 8k��'�)���t>�N%����G�:mi����JpR5x��<�_&�UϨNͰMY�(]�*�=Z��3b�祐9��8x���;V��G�����!�;��E0n/qq-�6y����R=+^�PKܽ�Q�na�pt[ꛉ�v3�`��R�.�$n ���p��0�3�n>z���̮
��3���U�׾3<�Ʉ��$�6�"�oS�:f�X(��������?�P���~]Y�;m�"��/��2��`�k����\�m��=���]�{�xM�k6!�9��,0h|&T�{���t�A�*m�-r��Y��y�ǘC%��IbH�Cz}�F`��k���Mup����a�1x�j�����ӫ�K�� :�i\S-��J�8P�ٰϗS!}�k3�n�.2�$s\�3�Op�~pt�x�:��{�j�n} ��Aڙ����Z\ZrT���C{[����sPOf�ً���'+!ӵ�J�$6V��I�*ѻ��Z�h�����:7RO��*��������,�]����B��E���C����L�9�`�'ў{u��V�E�T*u~��O=�E��S7XeV��+�C��6�z����,�7��v�S�wRhC��)��;��8XUX�+��W�x�M�����i=��ΰ�#z˫�dbS������*צ�U���[�C�d��%���Cޭ�E�\��A8�LK"��pfʮ1s��wb�,kC+h�ߢ6��=���]��z��N͕�x�
���$_I.��=Ci{�j�͚9���:�؉�7�M��#)��;'����tzvkj�m��������-������+�����#߳��B�T��yNR�G�n����}�E��B=k�vD�C��,���w:�.iS��*ΛjOc
�i�	���~D�	z�R9tK�?H4	y�����[r��K^`cZD:��Ĳ玨���r�k�2�Ũ��Q�����\l3�6Q��ϸf/��w��c�;�à}>`�D;)�q��άI�M�L�Za'�C�o5��0�#�[���3������f�G��m�_�y�Yfr��\�^y�)��[I���Z�Wt�L�s�PqB�u�#���P������A����¶gRB��j"�^f����V��0d�V7���	[�\�}�i]7g<��T��bq_�5���}�c�Qn��}�����O�|��y�mt^�×��"�R�wK�>+��Y�nu��f��]�>����[(?�C�ot0g������iz����ɓŹ�K�����nt���vR�
ә�Šv��q?o�^>4�)�|Qx?Ak|7a���g|C��#�����P���+ޠ���9�&��h�Wv,K�88���x5�%����h�X�4pwmu�k;3�-��2��������u��輳L�@������"fm��>m�lno\�n^u'��=9CT�ůd�w�d!�<�Ƚ�\���b��l$P91j+$����gv
D�}M�Y���E�v*��W�g��3�H9-�(�j7 ���l���Ց���=���͕��aKq�P)м�-ę�r�Os�츘s^��P.E���(	��iC�Y3
�e9mʹ�JZ/3c���mw Ӡ6 �Z�䢋�j�J�RaL��� 8r�f�3ĈM�0e��5�=�4��K��z'j�d3������-]�'b��)P�aU$��b�u�4.���y���%�ܫ�w�>}P�+Ehz��Z��B�(9�ڎ�u�I�+�:�(��w����z�l�.^;�=�4�U�sL=��
p����CSu�1�+.��wP`���Vr��k�l��ۊ�_�a�Q:�z��*3]�\����"mݼTz��9�k���G�7xm��o��2`�T�����.�7�Re���_<�/Iq�_����A�[�ol f��U��@��c;���\��	eGCM���x�2.�x�CK�R��R���P�Zk�/���Z]4^��g�8{h �^a�n�yNt	7B��&B̮xi�vh<�=���b��U�(f�eH�C	O�Ʊ@�a�_�@��{ʧ:��箅�H}��%Z"z�bI��D��;M-t��J����A����<k�����6�5�0���v�t�������h�1�o$QNec���+^�T��*9���&��v�����>'��瘪V����[������7��;.�hgQa�XR�m�Mc�(v��1���Yr��͹K�h�ê�:�0��u�j�#`<!0��
߬NK�N��v�9%��.�ވ�*�H���ܝ0�m��~���i�;�B��D�4j#�?Η ���<�;��!�H$:�T�;�s#f2�T��_�� ?�n�`��g�9�L���	<y	�
�Amn��+f����\<�TF���f
��gd0��[_D�%�Hm@��>t����]�v3��
ɩD�: 6*�N9k��`����	¤�D�ᖮ�އ��뽫�j��7���vX�Sepu�,n���/�ըp0��p}��(eu_i�b�c!y%���o��-��X��]{�e�xY��K$!A^k}�M�1p��L��XXd�\]�j��H8�s
�gu�u��c�ʪ[/�~%HE�f��\�:
��*�Ȃ��L�~�ӝ��<ƃ�:��l�5�]��w΄���Y��کnf�!6l��d����9GhY�}ǫxh�]���:��p����[D(�, ��"��CM�j�BS+�x��ʔ�5%P���'~��u�v�4�2��;h����
L�|~B�T��Q��������}t����g����п>ጩxr��9��{�5+�b��y��־�zA�lwL>	�!�a%Y��/�,u��(�-��'�3�9������~��ƀ��vTu9jw����N͋ϾDKu	�	�2��Wpȭ]���M�[E���P��Ut=Z�O�eAb�?7�A?ka�`����W<�~^�����&��Յ͈N�'W�&m�j�r��Ra�>���T;�u�9�K��v@qת.*������.j�s��Э����p�:�;4ڣ��2J-����`r�^��sH7Rͱ��')�=�R�j�
�#�_gMv0��f��Wd�T`��EyOU��m���6�rn����vN���c�&���zgR"����-δ�4�O��Tzk�3��P�:�Bm�؅G)d�Ot����Lt���j���d�2a�����V�g��1����Ő��G �߃�(��j�i�GuU�M�0�/:v}���S�ך	��mlu:�F����;�B�^9r�Ԣ�;ᚸD"��:�^��:~���}��E��������"i��q�;۫�A���b��:"���!��D��Ņh|.&%M����t�n��?P*6m<�vl�h�Cu(�7��\��0�f/����T?PȖxBK!�Z����*%�L:�kQ�d�)n�Bz-=�ޡ�9�i�h_Iaԕ�B��E��z�xiזx��~�s�1�����s݁sC B������|�8���S9�(2�S�P(���6�$puк��(���)�+�p�[P���b��V0J���#x�M��5yb�O�ִL���k���x՝�VV����;aL�(���dY*����$w�< �{q���e��E��ޚc~T�5�F��P�t���r�]�!�0Y�� �⮤*�ԟ���F]dD��|"D�7��P�*T��|���ȸu^�����YK7O��泲3ӵ�"a!u&ܲ$�����[RX[a+8����k�:7@8K�Jۜ�-�`Cw���&0S飖�#}ib���Mc�y"[Ҏ�`�Htޚ�<��+o�t�[��)���!�Kxm�[��Y��
�h��b}6�r�":+������02;%C�2�'.��F�*������/��!�?x��5��%A�{?-���Bn�NI�gM�'¡۬�n��Y����<����#�t�;uJL�qw�L�F�}���ÐkH�C�H��e�Q-��q��^��P5�=x��y�͑+(B���s;E�������v+J"��5���ܣG��>�r���>wM5i���z�m�ck���#	�5�LS�d���'(v�;�
���~����1���w����<x4��Nk,�E�+x��{	t��$�u���`H�B]��C���C�M�[����ݴ죺�����ȎXi'ә�Šv���\|xR���a �2�k�㟪{q����څ�ݛׂ�2�L�Y7�?<�u	��h�q�b�	���;�^���.S�M�3;Hnc�B���9h;�8��cH���ߧ�m��{�,�4��<�@��A�"f����cޖm�9�[v��d�v���O��S�ϗ��`���^&�}]6+Yk�t�=�!+վ�k����q�խ!����V!���7߹":���y�3�2X����\B�3<)#�h|(��#�)�.+�%2�]�}ӷ2\|�����@��NR�v/�\	eEΑM�S���A�Ɖ�L;�ݖ�N��ِ\׷�?dԝ!�k���}}����L����8h�c�9an���U!�t:T�4\�q��<6��C��]U�F=��/��l}�d	c@�@k=�|jQp�3��%�T����0ieQ�]���h�k�,X��:12��Z1iՀ�P�~UI�5-�Ʈ��uB��H��N��\��ie>gV���L֥�'j��d$_Jb��	�|s���P�aU$��b�gd[B�ެjmu��N�>���#�cL:!ā�2��bo��oJ�ˋ�LU�y^��@�4ʸ�\�StP�5nʹ��m�p�gd�xOH ��H�V'CO�Ԥ��)�u�p�t����OÞ����,�w���W�������Iq\�AY���u�����ě�F���
 �Ww[D�']�����F�xjʌ���\���D��D���Xw����?�ι�C�IuN(��u+'_m�BW��qvE�]<�lz�k	�a����<xAWW�~���u�����3ɔ��k�#`(a4-X�c����k�PI�_��|�U���=��T��#���D��1c5���A�������ײ�C����{��Xԟ���\�o�{���>FPS�8�X�;�,��R�@n1m��+���l�`jpɡ�Cz+�����L����ł�3P��	�ހ���.�̊���mN{�!5���]s�����y����/R���7�U��������}�;.�k��XsaJAbm���Z�R��z�������w�W���
��I���'�>!����%�'[����9E��$�Pe۱�u���3AS��Gt�E���P�v���
����Lxy���P��P{s�oDG|/�(��f�)1M���w
͉��u	��2<L�H:"�s�<1̀��	A�{�I�	��{l��%5U�lMM��;;��{.8���r9����My�\m�*��3���`3.��m�J-�c�u�.�SQ�F�[r���:P��*��}�0�F�3�6��O�䥯�ۺ�n�#�l�k���v�V�2V6�[�����h�L�,5�Iz0= v���5ȉ�	�Ryw�Y�[��<753�6-�A�ق�$3��6YS�^�BS+�S�J`��{"Y�`|5w&F4u^v4�XEf��*�f����4,��!Ŵ ] ����/�&�קL�N�n�MK�4"V��ǳQi�ůܑ��r�\� ����Z\d��#�*�]$4�!G��\�l:rtn�����*���>���}�1��o�Fy�.t�J�����[�(r�b�#���l�X����Ώ�xǫ�J(����C����<�Z�Vd��贫�=��t��/����ޑxљ�e�'Y�(iٶ�j�H1���*��ć9�CLo0���{v[��n�]��\���T��<S*����u9jw�����#�&�[��j�`����:
�t3n�+�*���{OI��~nK���Rq.<@����}(��f�M�����`'�>�n��sc>�-kӳEՉ3lW���w�Q����d�T;���ťç��5ʝ�o/����8>0�(�Z�s�M�稵��J��J׿�]DR�kK��f�;��?RE��6���|d0`�(G�"����a���^��#
S�O��l,17]�ov�r�[�Dk ���̨�Q���a1���MY�	�~]Y�����v;B=������ت(MJ�K���M �q����b�A���9aC�p�������������٨��:_x.��}�X�|z	HC�}�S3|C�Q?}��W������0G�\�����L�o>�X��ĺ��Ǿ��C�@��L�^��ë�+��0a��-����/Ft`�����k�������M�w@�֖�&���s~��O=z�g��*f�eT���r����>^�/o�����{}��o�����(_�	"w�@f��.��N�����z��}cIj�WJ�,9f�nȴ�R�!v�T**Fj�U��!�7}��r,�+^�ȦsU ��Sl^8���Ȓޛ�Rj$^q��ˌ��kpDe0� l�����A+Nm� ��i�t�y�)�V%�(|K|EJ�E�����4^�SV��-0�/nt�[�;@���cXy�Y���d$N�O���Y����G�]�W:Ucxt��e)0سI�&�R�6͍�D{�s�{��u�.���.s9u�� 6���!�FvO�v�mt�&���(b��>u�d��-��&��:ê���G7�1�ھ�/h����U�/��#뤂��q:#�
�,Q7C�F�[Wc���J�ɔ�9��q�_kWS;�]k]9����P|w�َ'�6ɾȮ���E�l\�;��Hq2Y�6�K���f�lL`�S����(�n<rv���[J�"���c
�������y$�)��sIs-�����(;K8�\��wv�Fr&*]H2��g^7��S�ѥ�]W9��ѱ���ԙ����K�Zgn���&o�)���c�9:]��k]��Ԛp;w��H����h�كz�ݓ��3d�5>8zn,��쨡t��>*��v��}����&b?zQ��^-�U�y� �Qi]��v�<D��Ah+*��nؿ�nS�{
�&Sْ�də]�e���B���p���R�˒ܺzrԬ�ՁChfL`�yl���|ZW�կ��.{���h�wZ�k�%ɕ��]ҽ�\�=f�vO�.RN�!�qU��5J��maZwr�ڡ)�@�,�ge٪��hB
ճOWM���S�y8Zt2���XVQ����vEM�����[��]�v����\���9V;!u�;�+E����C������n�cJ�5�Y�'wr���Q�K:S5��iJ�FN�P�4�T�"�m���D���"��W5h�S�3l�BT6r�����`E��ޱ�r�U/1�[w=Vۮw'$�^gbֻj��� ��Fչ��]j�TW�vj&;2U�뒶���O�&���xS.���gqܩ��tN�/�{sB;�P�8e*˥�g0���2[�`|��nl:���v���l{�B�ͼ�ؠ}h�[�w���Iku'L��rS��ݨt�[G�:88��qQѦ�)(�}�j4�d��U�s��^쳼/��ۊ��_!e�0��=�im�c(��,V�م��5W>˵L��	�0;���n_i��e�+.MFe��t/��>�5[��\�پf�(��C㩻�S=�y�l�l!H���9A�d�a�Yo����iҖ����N'�h���t2e��{汍[u�)�ws��˴"&6��7slڙ�is�;����41��{�7z+t^E�v�"�4Ņ �Z\�\��;ne�����w���ǿ���D��k�ۭ^��b���*-3oK]�m��h��X�wv�@���Ѥ�65�B���E��b�jMA�并6��#QV$-��,UU�W5F�f�cFحT`����sh�l�Ff��AQ�ŴT�E�k��Q�J�+FƠ������WME�X�V6��ѵ��F�F��ƨ�V�-��Z-�k 	� ��+��w����T)���Y��vq����%�Π���+MU��<���&c�t`�H���X^�3"y��Iu�l�Y`�������WN��|�
����9B�s��M�������RV6��;�Jm���ɪ��r�8�-w���_� �G3�!����}�L+��}o��P3��DC��nJ�j-��g��E�m�1]��[�"[y��
e~T�5�F��W��<�{w�\e����B^:�3�:C!�Q�zۺ� B�<�b%:O�"S��SH�kk7'��"��?���kl���h׵�mi���ɚ�����M3	9
f�T��"����F�W0椌�{}�?.��/�w%����A����;(7Vt�R{¥�@�M��='�By���r��-s�����׍Ww��7
m�:�̰�#'�s��9��W:�����݌2��Z����Bf\����vF��Ky6ta�#��RL!�����P�Fa�,�:�hOP�urdS�U�w�@����]�xY��{�	����O����MP�6�
g!���]ٵ�|���Jz�F�6Rm΍]���{���,
O��G�xO�q�<������9�t*}����㓎����_��֨=���J��������� 먎�T�XH�����\Hݰ�.�������WT���ZJ3�m.uYJ�A��?`"I�Ռ����3s��ݹ	�-�������K��������I�v6��ͭ�kE:��6�;q�j�R�}	k'r��xOV>�f�ۭ���N��	�C$��Nf�P$@��+��)�h/a�@���<��(E�pGs��vCB��"ac����Xޠ��:����\eش�$����έeC8��ݱ{g���<U@�t48�Bߚ�L$����m���>��,Ӏ��v����!)�q]�]T-�ޅ��^='�xT6E;ǰ>B1���E�j���3b���A�u���j��y׶�I��KXl����:�Ϲ�q�L�P����L�٨��r	�O��튮�N=�n���:�ݐB~k�A= ���Q�g/��ٕh����%�]�'r�n9��I&sn�..��lj0���!���RukU
V��
j�ۜj���uyθ[��zo2�mKx.o :�]K�N�{,�M��-��~s��J��2����l"f���y�m����+h��8މF3�!bz�\?��V3�����ӵ5��ax	��y\��^u?<��y��s��@�E����[��F3�	�== ��v�8���O3��=S��������0��Nw��,>���Y�Xd1��|����T�c*������u���;�Xrl����\���L������{�X7|;T�w{}��X�9�p���|��S<w�i-�MJ�C{RI�5��wx�ܬ���Zr�C^)���XQ��.9	r�*�_���-���JR0����̫���'��e+���m�er���S��??j�5�{�Nu�z��
2]-�Mٛ�}�Vm�,-��f�'��RX�-�a)�ݚfza�C���`�D@M������3��������N]V�c��8�,*�O1��n��Íg�8P�*�Ǩ;��v�?~R.���ڧ��q�[V��[�L�\�V8�Oҵ�r^��Q�'�hN�xs�w�l6��<NUz�F�"<��?3�IΉ�v[C:�jR�m�Mc�wh��R���w�wI-+�1�f�-����}d&]��g�D��A@x�	� �o���vI��;w�(��q�.�3Y�7����C�ʚ3�z{��۫٘iD[.qL������%��0��'�������F��ޮs�'��}���w��	I@A�0�C�,�xc[��d"ˉ��I�r��F�C�뜇	_ά�]P.Tc�@�i��DD�^��s�+$pDϛn6�o��ꌇTS<h�`�5�%k23�����˄"��{��j왆��.29�A���Q�[�dO�:k���o�~OѨ(��Bջ2x��w�0V�L�}��IrL=R����!甛�'���!w�W����R��öPL�����՗Bq�^MjŸ�#0��Af��wv�� �)� �Y=�_`��۝%_�]��×�n*Y���bu�fy������9jo��M>����2W�R������d&U�Ф���̨�ɯ�|jT��&ȧ�ã���
N��B��E��q$>C��z��CM�nt!2��)Ν�W0X̒����,)��Ρw���5Ξ��ՖJ�ZwAu%4/�� ��Q��ei+e���]��Τ���=�����-��s�1�Q�b��+��*V�d�o��P����[��F�Y��K�n�B�(��yN�r�\�x�T�S�o�<z`�v����@AC63{��km��x�7�ns�sJ���gT�Zv�8�����Z�O�S�%t���!��kr����`�����7Y�Ż�F�e�^`嵤B�hN�'A�`ZɹGF��9�J�s������D�RL��Kj�f���r��`8��9��=k�N�6�z�[+�c
G�k�PKܾ䝅����ʖ�g��}���]K2���E3���@B8��v�M"2��{�l�ʤƩ����u;��c?n��Vt�u��L�Qۖc@ņG��0J<�пy%�z��Dֿ- ��%޿zif~��l���+.��$�++R���l�x��"��k�����V�{u�=����F�գɣQ�CBz2y�V#"��SP��M#Bw<RSʚ�V�K��Z&S׶��y��S�\͚$�W��I��j36P����f��s�~e��'^� ^=$?q٣�W�LZ�X�c���r�=��{��y~Prڎ��w�k����q���m�1���i&����[�}�Ց,���K.;6/�S6��vz�.hd4(M>��E�OE��ޑ����L�}�%RHɇ����O����(4(k܈���׳U�sTk�!O,��9��.�##)�L{G��{[�:�F��� ʔ[h��YK9�5\�F w��u�7�S���ht�w�-��ȋ�O

�%{Q^��D���m�1���#4�����0
d�Ms��M"��;�V���k�?!���.6	+�AW�4�׈^]�,`�nn�C"8'�2/�)M2R�5;�=��3�?3	Uu�Y��1�|ke���R���7�����$5|�xw��?�Nu@�<Q���#ny���t{uJYNZ��1�ٝ��i����r�n��!�a�`�B��T��/�i�E��4���5�/1���z��\�����^~��G��Bm�N��Λj/c
�kdڟ}گNkd{�9���TH|4n��-�r.�V�w[����{c�UX�������\���w�}���a���v�btza���i
@���Ff��X�u�S�,��w��s�6�S��]3�v���Or"U7���e�%ވp�;8Ԭ�R���[�1~vʙ��.�a'�?K�X(֑C�|�e�sV;���~�_����PP̂}�+��#��tLZ;mn�Y#'�RL!��u���!��r^a۟�OP�u��/�l������\ZLT�sDq�˰���E�x����16�b��<�e�({b�ٶ@�`�~a!��ö�/hm�lJ�oN-;��v�Er̦E�Yc����O�q���/�Ph��(�Z����o��V�e�m��9e�Bv>׳��i'<��0�D�b���nX
/a���G ڱS�nJn�ּA���E�xc�غ���٬-Z/��(oJ�e�/~���Q���?����Ej]��j��a����1�\>��S�(�I��:a�^Ϸ�ח�L�t�#|c�=Ȟ�ٕ&�6=˚�V�CScW:�o�E;ǰ>B1���E��W>��f�kb�ڎy��ʝY-������z� ɨ�i��Fu��l�,qL����l��|��L
��ͳP�X�n�uZ�~ާ�7��EcP&O�~�4�p(ֳ��{lʋ�4.3�>L�9�Q3��+v*�f ��)H�V|�	��F��s�'5�zVY�;�\���GPѭ5}�Y�@�˄������ʰSs�`l3i^�i�%.��9Ho$�Z�s�5}�L���-oB�/��e+t���c3�M	�;_��� i�K�jJv��=���+�6ߜ�r�Ͼ�k�1I��"R�,%�T[l�C�e&ڪ%�wr+!���Ō�!7�2������xgK6��ū��'b��)P�c�N0P�C�(a�xELmk�v0B�[B���H����C*�f!�z��J�&�x��V�����CV�=�FӠ;4�78^���H܁!�!�O�'�_�e�8���1ڍ��Q�UU�Ś�u#�7�M��/�s�6���R\W(V_���Q�ܫ��I��?JZ�s�m�ECȋ�D�n�wV�!e{:�
�2��֮Ry����r�v�iؖ+��a��wy�o����	|���ۼ�C�Н�N��n���8���,�t��R�a)��W=�x�t޴cCf��v�ѓ6�EoV�m���֘
*���c8еaԬq���{*	{kTs	hN�.gv�Lܣ�;9�3�����p?�3��ZD�思�e��E�5aJ��2�~N����u�`Ȕl�*2��r��@�m�jOa���\����~��vI��K�s{Q`|��Y+C���`�*�p�����xuQ���gU��u�f�!x�s:Ԧ�^R��es�D��1��C3o8��W��+�S��o7d
v,>rf;���c�!�P��7���ϟ.���oP�w�]6zJ�%e����߇���y��i'5M;|/%����3'C��ŕ奥_~bhY偩�a��Z��U�ͼ���(n�`�Tq5�}@��Bp�o�3 �e���63�0&Be����+�O��ikc
���_���g��ZE�[���*����4���M^鋇T:)�-�%���A����0�ǜ=TO:��cW_�UKc.P� ve^��(�*��z���r�y;�N�����C��g�!��0L&�#��l�%cj�����M����ekU
�9���a�Q��m���`���/9�C�ᩭ��Â�K4���C�8H_ex���<��%1q�^H}����YR�f�/hf�0-AIT.�&����������!��/����n�EU4Wi܆P��yy�3�� /Ⱥ�yc�L^y���O���A�l���s�RM&#���k#D��G.�\�ղ]�Ȥ酎U(��x�T1u;ux�S��CJ�E�J�0��י'�w�MN_�׵i��!1�; ��7B���ʇBʮ������PX��0�Ʉ8x�x��j�R+��r�?-C�8L9&.w�'-��=]�Z�7w�ݜv���@�ܛ���c��4�nXa^��<�	_Vb�r�V]��ޚD�+w:8B�š��L�`;9hG*r9YX]��XeI֦.�Z��++>�U�eu���n���v6�\m ���>t���B5�6%:�$Ͱ-XNP��F�Gs��T;��ri�ぺ�mޥL�+�Χ�t��On [�{k>a��k�N�6��Z�\%X�Z��}�2Y�wT�łt]q�Q+"��k� ��'k����W�9���^a�]4�ۏB���==-���b��x��PE����V���?g��y��۲���'�T
>�0�\<�h��z����Og[.�~�nܭZzS����f�Q~���!�@��+��tE1j���D��ŇD�`�+�Zvf�mm�
��&W=��k��h9͜a����I�Hq>$�1m���˗�H�1W�*qih�.Έ�ii�
5��'�zǣ�#@k�2�'��Xuy+��0a����ˡ���l�Q����4S�/'�{hj&||�11�笈��.J����A�f��2ǥ�/ū��;�z]�ѣ@���+�3򩢝�`qm�����W���$Nq)��A޾�x�i���nF��6bK�Fu�x�^=[ռ�o��
H"XBkޢ�&�m~�~�w�Ŧ����5X��`e�0ǽ���>��w�r����`]�u����oɥT���ۙm�x����ww��%rvvﲎu{�V���~�bܜQٳ,ђ�#���ҩԃ۹Ƿ����E㢭�!͕��-�8�M�A�Ŵ���4r��|�]q3���]��.�	I�j1'�K"�(�ER��b#m���Ξi���0�vT�ޖm�6�ʶN��vk�r��z$!7ҋ��N��D�7�E1(�jn�;����=E:g���/U�*��ӥ�ٛ�s�[(],�S���2���q>�J�|"���}"�����Y�IB����S��o�c8��<��
C�zM�;<�:m���R�6�=Qi�3��'%�-�F� �����\�<At�s�;#Џ�LkÐZ���'\��������Ӌ�U��<��j�`����ϹP�$:}�/�C������D;'�^�+��?j����U�^��ۂ1�*���$���W_����'+]�N������>�S���F��xQp�v*�Τ������N�a4-Xu)�}eo�cӤI��_l?��C�OC�w�Y�pc7�44mf�޼���	��r��S���w�O��'�s4��㳍�+X��-�$]ޭ���5�%ռ�l��	xg�b9��!��>���oӲ5����#u	�]�÷6�	�{���_����������o�����.�V�)m5���d�΀��82W�)��d�S+J���&��ԟ*j��H�ټ����=�{�uY}J��
nU���'t��v8fX,��y��ȓ܍' �"�
�rG���r�����6^S�T2�C�t6�m�N�嵗R�	0�Y��=�]UL��䖂�uɭ�S>��!*��:��]*<Ȇ��Lٿ<���h=5��
�M��A/;�Ꜷ+}���gT��&�J�cF�W��́�j�^Co����t�9�տj?J�	\ ̙#�'���c�Ou���i�;��wY�R,=�^.�ȵ�9�T�K�!�n�Ó`���İ��c���u]+7Ѫ\-:���Gb=�K뱘]hu��[o9qkVb���s�d/�)o��i��$4I۵ٿ7flg�VM��s�jl�2��X��o�]��Nv>��;��M��P,0X��//ma�j��B])rc�y�o˓NdT��Q�R7��s(=����s@f����\;��sH�����e�6R]$�q�@�$��}����>�5v���̚��G���a	w�e��o@'	h,f�Kw���]�s]���1�;Y�S%ܰV	B�!6d�-�6��=]�ru:��O�[�!se��4�h_&�WĻ��u:�r��;y�uQ�0�n%1b�TL�q��[/%%X����o����d�Mu�������NF2�Ua���7�oi��^�h����f�r�DWh���EM���S�T]�����mܕ������B�j����@�i�&���6�iR��;tR����|�$r��o���ɩ�
۰��3k��cf���M�os�EmB9�
�g=���\�U�����-V@�X�u�0�lB3:��O�I�v���Ix/r",vS1vYJ�0��]It6xB'5�a�[F���(ocN��kTY챛(��G��Qb��zrl;/&�����cv/�e�R*�.
g@���R�w|E����g.֔G\�ҦWA9���9���elm�]��W/!ys/6U��n�?_h�A��5�1&'�ǥ�U��/Ygv��Γ��(D���ٳ�@����W���ި�#n�Z2���,+�̺:��X2N�i�����Gr�1�O�c�X.�t���"���* J��&�7E}V��_�����RWg}�wn�~�����pXA6�s�}��j�gV-��Q��� R�w���5�κO[W�upߛ�@֓F%5ڛ �g�d{*��ʂ]M�����Iwb�����PZ�d:G�p�;��Ύ�z]�&��XI�s�Ny��hM�r�K՛1��[�\	�]a��gK2�nB�wA��-r�9��rؒ�r�n�ܹ��\�c���Ƈ������(h�3*άD�V�A8�&9�jM�y�-�r�0ʳ:�Ǡm$��gP#8��O���r!�'�a�6c�"r�5���}��C�Ί�U^aN�pqc���S�)T��ժ��U�u��=da(�7L|�� � #[�Q��T-�h��b*hƋE��ە��Q��n���F��U*�E�j���W6�EDmr�6�B�kh�ͭ�c*�6��,���5�%��墣X�4[Ec�lmצ܎mnQ�b�(�IkX��JK%�k1�h�5ͫ��nl�sjD H�}�殁d[��-���>bW���b--euf[
D���Ր��t�6�2�!�k�Ȩ���Tl�5���J4�ǵ����v�;ǹ�]yU�5R|�DD�3$���
�]jjtGv�ՙ� ��&x����W������J�B�:-dO�ӷ9,l>���T���d=���o�~acn��%���v^̛b�&a�[�Z~h���"��`0&P�aql�ߦ�}])�0ö��%;�Lv�yce�� rb�\�
3���6�S:|�x�`d��؎�}=֮1�:qu���
&�q���^]'�0�	�� K��>��|jʋ�4.4=�̗�����y����^��qq^��t2��5�E�e�a����P��S	e�ٻ�/kN}���{dƺ�|F1�'���zT)f�g��[�8_Jb�:!2Of"S�)P�qCvј�V�q+9��Iqo�Lȶ����H"1���2��f!���z��T�vLv�:��f�o��ۻuj�1�V�$�7�����O6�bF3�	�:ϰ��B6օ~�k������'e�S�b)�M�.���>��#h��=~g�C���-y�!���Y��kA�[zm:��?�n��XU2��֮Ry�T�49m;	�4�v5�|�ï��_��ʼkg�V���^��eк��ݾHT�cU�Nj3m�����W�T�g��\s�3G!������e�N�-���'��`��;X�h�Z�[����]vJ *c�n�)��q�.�����K5>�y���c�Ǯ�]�֕o}� sw�N��Vf�>����-z��.�Mв���Uk��͊U�%=�}j�=�v���5�ܶ=L����ѩ�P`ȇ��`鹦�Ƨ�sm�Bպ��:���{*=����R��W�aUv�� 1�5橊�C ^ÿHd0�!��F�5z�sBv]��΢Ú���5a�Mcķ��`h-��w;�/%���N�u������{�L�w�\=h���m�_��$���ۡSr�B[�����͞�Wݪ�!�������#3�hv}\ŕ奥�y�`�^a�>0h�\M	�{&����s�ꙕ�J]N�/"����ԂC�PdLC` h�e^�xc[�q�Pܣ<h���a}�����A����~��T�3`�p/#�yj�9ʸj&��q�髦.Ue��n�E^.��PΈ�a:N&.�ߦ���UKc.P��A���(�'?�ߏ�N;t=�֬����-��0�T�C�<�����:g`��-�[U-�����h�L��h�ꉹqg&���0~�x�I��!��[5����W�e�b� b-�	!���HO�+�4�)�^oM܀�W��d"g��~�@�3��S�R`�܋5V`:�]]��S�V��9��$v�u�> `��aQ��t리��@o��nں���u�PCI��ɵ�wNz':N��]���\.���Xޙ�]µ�o�b���㷫��a���7��Nu���A+f'+���ǉ�>9�R�&�%P���Ǡ5��c�Hqm	���Q!	s�f�ԑMU��w]AY�I3):,�Ⱥ\�Lhi0�a��� {������>���_�7M1,�S��w\�t�8é�� ʆ"M4��Y�N�r�E��LkS�Q��-@;����e�%��m��Gf��2 �6��BX�OHLha�l�(qT,��{OI���.��{d����j΢��}��W�G�L/ù�p���\t��=n�'f���6��r+x�0�-Gs�`��6@�O#�4�Gy��q̓Ӈ���ý��p�_�N�6������%X�?�-c��V��;����%�^�~|`��'yQ������&<yF��i����)GM��yl�-������X��αI���z1��kv�׌Xgb\3P�~2"F�E�>r�r�3����;[�:��N�6C�����`�zHz���������c���G��W�$J>�\L��[��u�z1nu�X���q"%M�����`�A���0��z	D�H$�4��-��o>��g���[8k�M�۬�Φ�Kn�P��J\�|v��l|]�Q|��vI:�:�s�8G�y7ݱ�Q@��BQ+ϫ�9���n��,�w���eyen�'�y�S�2�D+r%R�����'=-�V�ޑ��g�,M�h{7��B���l������?���x ���L=�OBz/�oP摛����J�0�\ԥ�-��?���}��4�d�U�KL�eX\[a
y��v6�ߦ��^��q�.*�����,����Y~v�s��3#���q�5 �]O�zh3VV��J`��:�>&�#���	+���I���S���/7x��%6ߑ�5,SI�Q�a^=�m4�_�;�
`xarY���(�ʫ�������f�C��FB�m�N+�K"�R�dB�������l�z([�̶�1�o��J��otb����N͕/ޒ�_��O��O]%�|1�ީģ)��ѷ<�\Ҋ�~�9��]�Z��K�<�3[O�t�mxN竃+�,�HY;$i�I>�NV�"�j�%����Yj�Y���|�v�â��������Wf�"mLpm�{<�^�.�ft�cj���3�C�0��C��٫)���$�������t��G��9���/�v���������!e����E�E>�E��x^�#YC�Q���qxwn��v� 0~�vO���R�'7�@���	�f��ٵ�[�d�������S�A�c�F\�x���ں9�J����B�U�%����<�Dq;��1��*�VV�C6�ҡ�Ӻ�b�ȝ�s{�Tbi��0����]'R_.�r�ڕ��(U�)t�*�JF���*J���݋+t�̶�����'&@(=J\����#�[]�2��_�6�*<�dލv�;4���6]�6�O�~��w�­wf�8�v���ԦY��V�9t����sP/��P�nP�F��>�*or��}�;S��·LZa�azw=0�(g�e'��i�x����7{�<�˖�E��6r�!?��Ҋ�,������K6C�9�&���06 ?��U�j]��m$�z��?��*����"L~2�/��?�Չ���s�ޟL��d��K�n�v:7;�q3O\w; ��� Ș��}kO\�o�E;�."��aql��YX��򡢛:e��&^8�حj��H88�1nK$��g�b�n@�t�9���R����`�6�ek��
˨zOL.�ʊ�\�'��0�z�	c^(�3ю�ơ�s_�)zYqs!֫m��� ��!�e1%�B��-�럝�e�y�KU
Je0�Oу^*�4c�5��S�/w2�1������Z;VpT��Őe��'l��n})�P��=�)�x���Y��]�4���<���q��Q�M1�cCIQ�o"�`���rUv$�f �{J�_�=�g�b-@��g�^�r�녠�va�I$�Ɖ�*��7,hrl��*_P��Nd'���\69����e�9[��J�S�zR��Vn5�!�3���v���%c#�Ї\��8�#f�Od[B��oH!�Ez+ѰC*�,�E�l�6��s�d�F&���uף6���-lM�9���e�$�+�t�vl��������0�'��/�1��������v�)���.�fy��m�tY�7{4��vk���3�kd-s��[;:m�uw��z�0����	Ȥ�:�J9)��B]��j�'� ��f49m;	�O�ݎ��f�I�^Y�u�����)���2OBz+�\��a̜qw�Qa^���fT�OtZ)��4�K.�c�Y�ʜ:���R?74�P���m��hZ�J���c���Mز��#j��H���p���%5x���@`�G���-^��\�ò��,5�����[1��Q��83��o.�t;Nў;�b��h�z������M�X�쓪�wf~��#���[q;�V�^�F����m���o��A��j�?��H4<�V�����=.K�$Y��krV�{~`�r�<\\0�{�RzA!�2=�2���˞)�y��m���$~/~݃�TH��k�*��ᦸ�i}�����ڬ��]�@`yot�nF\��43�1�~��r:�FL]���?vmE}��Si�jI�1��E�E7��e�S�4;�8�j�l�e���]f��bi�l�����������D�^r��}oJ�&4��?V~�Y��>d"�5�my�F��[���>+$!H��M�Ӧ&u�`��q�LQ�r���yg^Aa��8���/sQ�]~ʩle��㰃+W"Mh���;ʷ���!o).j�a71P�)�����Y�?;r��J��[���!6��fvR�mx��&�~��H?�3�>3�?k��S�
@Z�1m)ė�`$'��CM���Y�6yfhs�ۙ��T��%2��)͂�0L����x��o	���L�����ή��T��Qz�7��׳D/��4̤�Ĳ.��X�(�`����w0�_Ϭ��6��N8sl��m��(Ds�Bvi���.��\������<S͑�ѭ̜!��EABŜ6�|�x�>1�7:p���3cLp��^���װ�
6v�8���]B�Z~b��=�9�_�#}3d�4v��p�y8�s�m�{�ɵ�8F�P�E���	�c�������0�#������+Ք�^�8�*AY?�v�9�����&�mQ�Z�W��s�����q�(�O4�n�4殆����f�z��j�#sy�H��Sh~e�;�e����X��z�A�n�.��;ާ{2��7�;կ�7vL9Zs�x�r��u��2t��O��~������;23�^��^�\����q���6�Us��������ٻ�c
͍�����{���eK7i�`�L��t4JS�7>5���P��L��n��{z"��k�vl�2�1��:�lr�N�3<�j��ņv2@vp8	��NգS�i���]�l>����^5�?p͐�}$�X/���xv��˾�:�R��tH�[�OK�>������m�l�N�}a!ָ��6^�;�	D�6׫kCH[�H$��Ɯ�i�v���U�4��q�!/TS�;P@�e������y��DO�x�֜��OV�y�i�N�ST���ڛ�ת�b�6��l(X���?~+��t��;��ڵ^[H^��;�b��EF�G6VsN�e�X7����v'�4E�&�׳}�ʌv�gEC�(.�()�&��* ��=�9�k+��ӱsV&�A�ʭwF+P�������-����*ʜ5┪
x�>Uϵ[��t��n��oGF�m�b8�tp�b�_	���<$��VF�EP�"���
����+�f~MwSx���Nd���ո׻gc��
�nLb��1�g��Z0��L�sJ9��,������������ۗ��ro2�Y/�w�c;ۇW-Ӛid��Qi�i�[MJk{�v�#|t�pƭ��k����yj�euZ�m�}�N<dd�}5�y�o�J��>�[kz�H�H8���N�y\{A���������c��N�.��Fc� �� ��_��oI�|��K�}�W�u�x5�z��J��-��c���w���F�����>��KJecy�m�{�<��5�.��"��gs���`㱱�a�#x��(Q�4��mOݒg��	�mp��{��ܛ�������QBJU,m0���z����U����3[Ӣ��	(G7e镾rWQ}Y^��]bLq�7m̭�Ͻy)fk�,Ýay�
����ۆ��e�����!�J�Gf;1*�0�wp��eᨬ�|�s�F୓A��}���Ќ:��wz��`�T�=��46��VC�4�͉M�q�tI�g\��g@�h���G^Q|�ˆ���gh��ޙ}ԅ����DH=�KisӜ��`�!e����kJ�[MT��)|�6��o>Ȭu�w���WPq��L ʳη}nz<>�/N.Qw���٠�+z��Ur��������u���,�_3#��ǻ�s�<	�ٙR�R:�t��V�z��{ky���+��)�'{��!�j�+[�jڼph��=�:,��Ĺ�n\�<J�Y��� h@�JȐWE��+�������h�h��fI�����v���y��<Y7Z����4�Rh�� ����9�ho7��~�����މ������
��Gn#^�]̂�FQ�2vMt�4���\�ti�K�@Q5h�궿@]
�d�֎Z�顰R[*lf_���ZDNO��ܡ��<HG��u��ȐF@t���!H��2]H��kzc��y����`7$U�sɔ������ә�p�r-�n�uYc5M���&bd3��"����Q���S�7λ6�����+ldUCJ���wK�V���2#d�jz��W<�T�P+�t�$�$�dE_[Z�l�u�����gG��K��r��Ӟ���ʅ������@mbUV���؁����gd4�a��#b4���7�V�gR~Y>���>�g����{}��o��������ᑌ`s�S�d�|�up{���_m�$�e<��'�%ԩ���z�]�R[�C�5���qd��5�,*�A;L��Ճ�ˑ)���Vc���=3�U��R]w-���[l�`Fle]t��f�Sd� !���j��<#Y�9��&�R��|����u]�[���r�n!2�v��tV�Q\���)k��Egީ��;o9�����%��y)v`�/_�rN�CZ�ɗ���b�����#l�n;������������w/>2[V�Y;��.p��v�['e S�k�-�Ƶ�˅3��7'i��coDo7���jG�Z�Xmض�̪��@�@-����3L�-ۍ�%j"��r�g��,Ag�8m���lpbe؄�R��b����eK�qH��bQVv��\��w].����
7����k�I���
���<����7]�A^'�a9 ���h�r�� ��Sa!X�F�P{���5���7yw0<\Crb9�5��'_-�*�t�\c-���ݕ6����paU}>yh�CU�I+ϤZ��v�(tՖ1���l$��j�X�f�����fK�js�e0v5��/��hq�-i�ڭ6/2r�
M�{+��z��k��b��N��6�n�V
�μ˱���lo"z�P��^�1F1�bZ\��I����q��by�!����n��ݾ��Nݖ���Fb_l����2�;�|X��N����yS��h�y���Yov��s�V�=V�셒�
��L+9u��L+BE�a��y�u{�Zf{Ew�sͱ��m�����}�ӸCd�Y>��woGs���2�V`Zs1i}���gwD��G��Bl��D�J��:�&m`Mc�v页u�������y1�Ca�5��mm�F5�n	
췶mv��%Q8<�]���s�C�<��"++���	�ܣ���݃gDla��![֨(���n�cquog)�/��K�=Ҧu;���cRR�9�0��R�6�`�͊B�= |v����o(X�n�iV{ �X�s�͡j��d<�9=V35f�b�������L,��t̪�IS�n'����'�	�{���Y��x�(B�i�o��:Y2� �,4�ƣ�3u۬|ƍ��,XS�0�1Ó4Q��ܣcB�Z:j����K��c����MΎ�Y����b��+���ȸ��'O���A�V��a�v�oY�l�jl�Z��S*��������gJŋ�%�qF]�J+g+պ�m���w�>V�m�+����Rh@��j�*�Ӟ�N�P�SRocα�_1ZF�=Q쩹�]h�� к�䎲[���kݚx�v[�E�6)�d���[58lG}�ӷJ���S&�0��ۡa��ƽ"SȀ]�M�uj�P��913.��F1ϫ��:�� �;��
�ç,P�����8n\:a�vs��o����O�_ ��*6ɵ�KQ��E&"�mʍ��U�kr����1m��v�*�Ʒ1r�6�-t�6[�h�U�[�snZ-�m�r�cjū��ۚ�\�5EFƱ��mE�j���sh�N�kL�MQmsETn�M��j��EN����iݷ5\�6+�[�ۖ�\�s\����F��si��w���y��������������a�����.m�;mj���or�|�=w�7�3b}R����0������>h>У���u�#b,�'_����Ѿ��oG�b3��Y ^�����z.J�x��rی���y7C�E�ѽ���c��|���m6�p}z�S{�Uka����yk�>8���2D�n�.�;v�s�ځ�pU�˵�|��/ݝ7�צtU��$#/X�n�^Z'��/ �>�=��%����3�gx�|�`��:.��*5uٹ���F�0�&Z0�6��U�Uw��jNFk�
�{�g��,�p^*;�\�����.��D�=��u�7�B�F��wmѽ�i���϶Y��yd����(-Ĳ��EȦ�=���u�xv����)9T�O�i��ǀ9l���ZW!�x�X���Y��7:���q�!E��]hs����)*��w-���<����nU�WQ�Z��l��h�A��EiXJJ�xE_���2���k�@g�7ᢔ�x�e�w��җV9Jcde�d
EwP�Em��B�X�ui��_*�Ρ�d���H��*P'��4�qc�ȶv���t��`��`�Ap�E!�;e^Z�H�rP��Dj�[�훔��E/��&�JzJ��ѵ�6v[#[.�({bQd��y�u5W��ɶ�3�vo�^���Wu	��"�)�WI*�R*��|hZ֭�v�vW2M�;�V�N�х�w�|���@��GA�'�+_E:��j�e&�ݮ�z1ۓ1��{�ͻ|�N#˛�0�,��q�S����&�ɨn�MH�EX̽-s�\��7z(Iݐmt�L���`�C{��-��l�y]��T�K�̥ը��m�q�ٵ^+���qr�jl���p�r8��Bv.�!S�\Qz���;��/S������9ZT�1�d �n�ql�	�v�zq�m��o1�r<�׵�f�>��=E�H�-����$��o:)^0z�����5G�l4�q�T3�<+5x��wz��I�D�A��_3j뉪l�؋���|�(��M�9!�<��m~k�?J�:*d�$'�Ó3X�<��cے��=���"A%ڲU��s;,�1 4n�w>+g����;k=3SOJ� �XOn�MZ]���y�Z�86�3���)1mYx&�o&И�l��æ�&?A�z����k��_�L7�j{��w���o<���u��ۚ{�pk��L��f_$�;�q��v��q.A�LǽLm��v��}����nq�8Wms�w~�>��6�3F��8ӛJniԍ��n�"_"�`��k�f#ݻ
x�Y��l�2cgy���+2h�b=W���l����OV�x�EѴF�W1�@�	�[ k�U{�z�פ�H�O�=>ջ��1S�1c����.�G��S��@ˏ(B�W���&F�$o��z����.��ؖt�[��9��2��t��}�O ��Hl�7��|
���L���u�V(N@̍{�(���ػ8�;5u�g͏��[���]ʒ��
n['	<�~��s�'tn_�R��U��4�-����S�����0[�ޛ�g�3 R��J�q�x�"2��r��U|y��Wt��� ��� Cz�V��ڗUwKGwt�^�/��/�9 FO�Th���iK�ֻ�(IP�FN��uym6-�E�L��3<GQ���$f9�$^�T��_VW.��c���S.({+���Տ�΀wJ���=;����@%�k�1D��!ŻB�_�in��Q{��h�t����XDn�y��{����� x��J��bnd�7��Ԕ�����d�z�ʃ�GV�pΚ�Q�QL�������o{�����=H��Q[�ќ;��z����W�,{]�2m���í�,�ٲ�W���x���T�uV�j�[��m���=A�sC�9����f�aԬ����5p(�`���|�2�w8ے&��nR<��G�\�C?�1/�<$�S���*���{��:�g;���D<4x�"@=��ڡ�ndl��/�������b�vy�2wL�Ѥ�W]���J���+"}t4��V��Z�Y1� 2�<&�wz�i�pʎ�{�O����\B�����G�1Wa#f���LC�j��ʺ���ӓ�E&!��
�� -�k�+����׶��u5�;{��f��h��`ޜÓ����4�}V�~K҆w��
�2�sp=-g*�.ݎ6��F���RII�5Ot�r�Of@G�����53��m�p�y��]s�t�v B
��8�cG?ȫ�!.ol���s9���\q2�U
Gݽ�q�4�;(:ɸ6�d^�IV�5�o9�ڽv,G�,�</���Ϟݍ��4N�*��u� �����k.��B�^ڝM��k�Rr�	t�����j���sMNy՜��t�rQ��c��\��G6���P���Ғ���V���Ue4Q��T�7�tdb���ٿ]$��+��|w;��5�ߪ*�8#��@��#fk���Ԫ� \�)RTWve5�%�U8r�r�h�Y\[e��l�p`0��:[�#e'2pY����^��a��,j쵵u��eLk��m�AS��7�u�՜ew��b\����d����O\ہ�QOR2�[�ey�=��?h���q��+aBۭ�⚻3�{���"���^�r�E��oa��߃$p-�ӡ�3�Wz̚b�
]�y��{dF�3x���2D�,�n8�{�Oi�9�oC�|R�PM6؊���k�E��<U�ˌ*=���b|x�>)!(��3t�.ۍ�����/5�dQ���Y���ѵuٹ��gwܬ��sk_nA�'y����;Лnm(������%ow&�c�VE�Z����~wk�O�S��:D^w߸׎����h��T)j�w��+��xd�Y��o�H��惗���k��E�<��/��Sn�{Q	;}�P����¨R�N@�a�k2���ӫ�9��X�w*��`|q\��q���[�M�U�)�}]���M���q.v�����ĠWfe����y�-��.�=��E��#JIa��l��sU�g5l��`J�x����&j횙�C՞�;����HM�t�L.�%*RUW�*��L�M6�TJ���S�&rc7���o!�s����OBK�/�)3Ǌ���a���������+�z6���8"���z�x)�QM�J�ʑV9���|ܩv�"1�/Z��u�tQ �m�Mp��,�#5ug\����S�{	��>rE=x�Ӝ��W���翸�O���u�<_C�������ѷ�NS��K/pY�������>8y�s��k�a��og�oC���N�V!Gu��G\t���Ux�|�iP�.�*�E	Nf�R}�������ӹ�Z��k�M؜.8��c��@���>�*w�����Hm�w��%�t�e����ƅ1;m�6��M�4���`dՓ�����zL��Õ���tX��~ܘ�2I��|�p�n��θ:��wa�4+j���o yr���3��bru�<:���G8p�l4t��Z�8|z�F�	��oN�M��
ITOPޑ�7Kv���*\�t��G��PD~u�,��c,�z_o��/�x�f�1Ϻ�f�I
�j�ᴐǛXDm�h#��ϕ�sѺ���6c <Hr�N
=�i�ӿM�KFz�x?	���
�5���!��t �����7����vr��f��/����F֮I\ ؉y��Bn�u9,����E\�4V�g�~61�7y����Vd��ld�P�ևO��h��>ͥr��	j����Q9<�R�a���ú+�q*U*�hF7�g��-E��;�b=W���:�!��om�j�{������h�ڦ�l�t
��Q�
�*J:����;}�^3p�U��֚4��[X���EO��W����d��A�f�>,_�n��;�(�̒~��'�~���S$9�+G)��tUE�=��,��Z�h�����>��5��� �\ޠNl���NBٍ���w�#R����W�<r�OEɅ��I-6��G��N<�^b�M=Ppr�{�����^ԡ�lѩ��Wt�G�
����H���OxǱgHgF�êWvd��*of�ʂ�t��7�p�}��P�u�����(��\�b	CR��毺������}������ ��<���%�i-���!d����p�޵u���g���=�׆�j@FJTKz�Wb��(���Wt�.ǂ�m�&��tv3������ѧ�WuÓ�l�'��񌺭)M-�$�P0��Y�v��Q�:+;:X�Xću�Hτwd��ү9+�>��9w_�u0���5�XU��d��rF�oTm�RZ��w���C�#B5���(�90��5��3�6���Y`�GI�3��v���u]B/��M��ڽ"�(���{�8n�v?��D�5���[��Q���C8@�{��^0�2��;U��^wNgm�E����㬞�gޖ)�|����������$�r8{��sYپZ�'<��>t3VJ��=��}3S��S��U�0�r���U=B&�s����䶅�h�;���Y��y��l�l��3�TÖ
o�l�Z�wgnT�}�7�����h)õ�༫��IĜ��y��34���$!-A�z���¥�|�y�E�� f�O�P䜻F��gS��c#z�7V�}��ل���"�i:�ӵCraV�n�SY��f*���=���y��oQ���M�V؃�Z7y���^�����.nN�����y"�gk��P=y=4�&��=A"[�^�V^ǥ坚�s��F�w�ۭ���h�qƷϖ��u>9�!dH]At�|��$���׭V4Zcٰw���|�R㡲�Z��d�W��*jC���#>���0Jy:����Uz�h�)P�+��6�����q�u����{l�<�`}5ϣHa/�,n�9�S�ؕW��y�IR]��$��1=�vZr��t2J83�|���|[ϰV�����\�t&�&���S�n�s�ݚ�1�u�:�?���Ì0��^3���5��C�(֥��Z�c���?Yއ���\�H��1�n�Lz\b+�:��q��T����z���$���5=o>v����������!#)uI��e���T��5�hW�\�Ya�xOt��<��ᗹ��ҧ�J�+��|��s�g.�Oe��\3��\ȭ�@�W����vs�B�����n��tDf_l.�=W���!����v��f�CE�<��k��hn�%�<�a}����T}��{�
�����<`�[�x�{�Oi�$����`���G+�[���27��s+e�7���bA�D��%ݶq7!������Qu�65Ěy|��1Y��J�n�5���	=gWM�N�㹃v�鬘1��d[����f��on��:J��Kz�L���-������ũ�[dvm�v�.������]�#6����,�B��0�)���WX�={r��;r_��1x��4��\�O�ڹ��5maS�3!�ӽn�RF�`�q�m����,��G��I>V�W��>˂&��Ȗ���y�;�
�>�J�;���z�X)��x���r�5s�eM�V�����$7S���4Ty�[�Q
y2Β������ӂ�%i�ƛf��w��omt�m�� ��O�5u{:����=���������=��g����{�||����0<!��x<�Nؔʧ��[6=#)�����b��f���
{�$����}0�C{kݐ8z�9�g�Jebk�9�%�� ��G��s&�6��2�g {�1^�����<k��=�9L��$Vs&`��/r�Z5ٮg�q�E[�3L)tN�g�+'y*3Z̀s4���#���-^̱�;1�ʎ��72s��+�TY����.E)u�L��1��@���"�&N,��p��o3m˚��X��"�4��R�me��j�]�[y�<4e�䍋2:��Y���)+���ngN8+�#�WP�w)��h�VvLz������U�&Q�-���I1��c7pm)�����"�� �֖cI����+V=go7��G�����-�"\�4������[�j��/��� �����:_3ek�)���nI�:�1�7�eխh�N��l� �|&�KF�:�-6�4���%`W��DTG�*�O��{ֳOv!�1�I��Yp�c�wu���ʜ�$�7w��y�W�M#�Բj���E)�u-;ͥ��?]��w2�&���-i��nv�K�#I`�h�Է�,e���.buۼ5��k��׳.��}6M�$����Y��b:��\�8��P�F�m૫�y�-��$�p�˙F�썪�$"���C2�=̭���Z+��L�-�s�{���r�4[��3Z�GKp�t�uݦ�l���Dv���e��bڿ��n0N���7��k#+���e�:�MP%l�w,�Cmou�͢�Hr��[�^��MQn_=;�c�,���%�9ʹ�_>0��pX3U��9l��K4vf$��4<��fˣ��C6,�j_wSڶ���ESRu��\i��fpu0����wmNV�����L��W:�Q�̀�E����ض�o�p�u4�VzM}@���P�N	T�'��²i=%E�!�asĻ�,���֙�h�dʹ�V���^�1��>0 7
�f��ei���F�7�zs�n���U��)_�"��]�����1b�m!���cǋ�x���Gb�h��
���gI��3i�i����A������CrwF�76�vby���(�S[���w[�T,��YJ]3��Rr����q�}p뱖�h�&�t�;)�Av�N��H����>{�i�a��������T3G2j����-!:���E���*{t�S2�y�f�h\��S鎳�`�$W�v��͡����.�h�.w�*�r���
���w��)u��NB��7���l��͛��ɗ���y��Q�]��J��[q� ����v��VOAư�x��I�	j�X\�GT���*rŔ�r�n�a-�z�_s@wt4��j;m�U�l#������9N�U���9,�����ټ�� ���ffe�֙���\��ϋy�/��V30��q��:�����_�|�F�����\��ֹ�3lm�cTZ6�:�+���1WJ-]-cb�9�Ms�2�˔i��]ݹV���-�ܪwb�����t����-���WMn\�4��͊M�p���m����njƮ�Ɠ[��Ѣwj(�5��\ڹ��"�5r��ѹ\�k�scN�h֣h�X-rŹ���QQ��s����.W5�K�p۸W彾|��N���^�oQ�У���й,���8�M	J��>6�4�j5/�̴�9ن��V��p�����`gf��`ŅȂHLt�A1�.��"�(�4 ���"�_ư�y�������fa������*�(�\_�e��l0��G�-��6�3N_u5���\�kb^�9TJ/4���饤�8�j���!��q���5F�j1�.�,�Ρ{���Dt�g�CJZQ3%9���s|�00!#3'hB�٪4m�����ۙ�ޢ]n�|9ZT�q���^fe.�i	�n�3��9��[ҙ����Ŷ��1�^�������킠�P�DT�Q�Lb�+k".	ޕ�'R��5�߇vm�Y��Vkl_Y���zxD4��wLq���͢i�Ǫ*?��5���]�$�Y%�)��fZ��C+�s}%����;���U��|��;�}�����y�b��������{q�[�%I����ևI6�F�Fm)�a��U�hD���e�.��i���{A�{�4bU���o�()���ثǯ��+�ݴU3������6#4�l�ы�/������g�j��{��WM���K��[*�Z��S���wx�`���i:�Hh����ԙW��L�.�Eg  F'�����+Z�@��;9���8�\�L�:��v>ke�n��)�E���D�s=V��i~>#�T��D�sʆJ��CUR�x�*6.��i�����70KvtOl���~�k��T�tU��/��k�Ldܹa�.�k5��ދ"�WRIM3�tz���i�EӤ8+���}�Νޔ
�j�����q)��<i�z@'WQ8d6cߴb[��`�ѝ)��6l=XA����:��
�P�K���5��sty�@��P�t6��娭��C�*Dd�Ɪ�5�^JF+�@]� ����c�FPT�v<���4ǘ.��z��r�9F��uCJR-�i���x���\�*��T��o7Ӱ�S�!�I�|��f�J���}X�l�"puN��ξ�4�]ۮ�� ��u��o� ���e�|vMJ"��*�xUf��g����^J��g�;F}���m�����{\�El�gE��I���bu�1��92*q%���L��Q�x%y�F��&��|�j���<Nt��ظ�V��J����P��[�X�Ev�v-�"�#�MR����iD�W.	��E�jg+xl�.,Ӣ�&���]P�zhoIr��us#Y#�jG!�M���=��s(�fF��;��`q烢��1������G��k�]V�Lh�gοF^�y�Fn!�xID��mWE�ת&�]=ʎaս� ��|x�{�,h�<
��iTM]^�-H���+"J�Ӊz^��y.���ֶ�g�j��_�d�V<��=T���ll������H����W����;�y�2�CSٮ��ߩ&�{���tň0���F�W,��j1e��Gdj��z9Rz�sh�o�{g�}/'��&��n���S���&���"so.7v��8��M�H�I+�% ���S�n�vdHYX垍�5q5�qumv��K%7��l"o�"�sɕ�{j�{d�nQv��e9���Z��+�G�t�;�H�R�YM�)W�J�c]\�]m��-aw��;�v�Dnoh���%�B�d?#]1�Ī��y�I?�ϤB��3ߖM?��c��Lnw�iF�:xBګ�0�= }(��	�+G����G���E�����(J����[��Ua֡x��ߦР{^5)�1��\u�[.S��޷F7�ڤYR���ݲ�{��f���w�oLv'[�ԙw���2��#��������|��o>AO��Y��P��m���=gZ��R��1@Jݕu�������ޏ0�
���4�n�ɊZOZ�2�pq�g���wI2�����׺۷�9��W�9Ce�
j�.�h�v����k[ڍH��x4���l�5�a�5������h��w��1��T<��G@�lW��x�ź��a���ݛ{��U��[��C?�s��u4^2��w��1~��D���R3ak�S��r��to8� t���3�L��a6�q�*�w=xH�8̅�c��]-W�/�;��̢'��i��#��]�ЂP�MD�p�x-T���ę�;�N��a/��")Y����UD��d'�A�8�*�{OE;v�Ş��n��ڂ�RTT�Iڳ꺷���G��6-=?����u֝�|*I��o]rE	��f5��>��4�fv>Y:=��f�dAFe}!W��ؓs����Y�t�u�ф*����m�q��N�y��u�d)�=׫�
�yB�\}���R���4U�����M]��ݛ�^*=Jʚ�ބ������ƌ'F$�L�W�
�5�� u�/�O��R=�P�R��U�ʶzh��mp�`m��{�K�l������� 
����IYxK�;=�n�N]L;����щ>Q��O�5��*��6C��3���9�Lq6{�u�^��w"���ϯ�dv�K&�)�8n$�]C;���`�}�i�g+��������_�%q~�e��ly��`?Z�z���j����V`��x�>���8�W^|)g<�ݐmq���C_��u�5�,���6�_K����) ଑<�:SwI��-����Nf��O������jiZ��e$nyA�pJ�ۗ�+p]@S����v��65�Ƙ,2�L��t4�>��:Co&@�m�q�����G���M*�&�Q��9��Z�{�����tJΠ��]��Y�Rf��J�kh�vl�MY^�b�i��g+��p0k��y{n*i
���WN�b�S�;hg?\q��ķ�a;ʝA[]�K7b���+WL��4��G(�+ho6���e�};,�O]����m$"j�IefV<=�{:C�5��,�R�Tx˫�����;����KS\�C�.l\�wj�2������(�ا��g;�+��$��k6�S���vw?UL�wbu�;yqTA�t+)k��l�{�t,���2�]�ZkEѤ�*z��bↁևH&Ѣ�4�6���[��1�-�c��-}M>ې��T����*Ĳw�X�()
㧏b���)�]��Y����6��ĽP`F�V��v��[>�@��)F2����]�F-؎ދ����W#U��U�y�E�r*a�*��|���a��[=V�3b���o8|J�RS�}��S��l����&���;�Tf��q��ކ���
E��IX�\h6�O����o�-.kr�u"�W;�X6�3��2+�ErJ(r����`,����w\bW�������r��t��=Q|�bW?Lvv)�Z�(���Wt���?���{������e0�ڝ#K�E�D����Y�l%4�N E]5�L�hyB�ǖ����w0�~���N�/r�4L��ze��v�j#�9ٚ�:��K��Rd��5��3 �*��\��G[+�(�$�]n�S��������ޛ7'v"*�F�謪��&��>��{G}G�q�^�W��F��iJin���_�oY�}A�����j^MN3���އ	;��������n,b���ꮛ|��c�~��{ʪ�;Cg�A�=�oo��.������!�B��= ��]�F��#_o8�^At΄Gd�1����2:��C?�s?�Q<,�9�e7t�Ι�3n3���"5$���}:c��6��<��K�Cn����f�e����О��rS�YW�o,��z|xP(�$���@�f�[��ս�f��|y"���2)G��5uB�쀵 h�R�"}p2��~�~Z�m������UIs��rc�����^���U��^17s4p0�ݨ%�՝-�;\@���6�8�7>������0A�;�,��kl�ѩ�0�y�wz�� ��I1�wǯ'�4�L���Wz���DcfQz�a�����۳���-�n�꾢��sjmɝ�{]o�L!b��j�O�k!	|��a���*��|��~]ғ�)y�N9�%�3r�78�3in��Ք�=�%�_`n�
:���/�pc0��K�\��U4��E'ՊG����yqc��@�ʕ�r����c�����%%����R庞��T8wd&�RƌDj���!e�"��t$o�"���\d6V¼����&�wE���ѓ}ӵN��!���#H��E��a,�+�����mA���鶘���7��Wdo�����~��g�h	��J����CP��),Z�����t�gu�<�B����0Y}[ϰV���C= x�k_n�s��gr�Zq�f�wHۭ�E|7�<:0F�������W9�d�g\�i��Y��iS�r�VP���,��lG�ߴq̋�`1�7~�[>���t,^��ˑY�Qԍ]�s=׷�{�ƨ���]�GxCٺݞ}�~�}��
�����+W�"@�~��Ffj��6����Ѵ�%��A�o��p�q��y�Q���w��זbA�Dv�4�0�9��UQYat�Ӄ���u��Z8�l8n�lw`ʗHf=!���.�-���r"T}��R�$���/��12�,*:��;_M��(♗y)�D��e���o�(�`�z6�l2�;�V���Q�M᝘zs��w�6;���nY  �G^UN���wx�!��h�ח3|����B� ���׫^�[�[%�^E��+ö���0�ou&�O"A�M7������t ���A�9�Y��{�7U���s�p���z;�.�u>�jA]m>��"��,�P��3��9s�0�
�B �{�1�B��ulr3ثj��4�s����L�+q����:�R���":��˧�:auq)R���Tz�ud�Wu���:�G�L`	�@WH�d��+x��I_��+;g;z#z�>���=�3w�>�Hu~�C\r�-��
l�Sh��^�ɣO��+�k�^Β����gݵ���aH!!�,��]�ǅ�!-�0��D�^l��y�P��+{^w�18��'y�I����a}�c��ȸnc���z˶��U�>{�hF�U��}����q<���k���c7��y?>W%XNE���os�pP�#�h�ēط <&ꆸZ}���V���-A�!�A���;�(m0������Xم�9`��$��+�j�v�m�x�u��o�{���jn�(�݇59ƀ;ǘ8�͠Oc�V�	�y�<�QV{���辶�]���g�ѰO�מ��!���Җ�Lz��I�fp��"�e�ff�/:g;k�?!^�Ё,1���^�"�w�iQ��U�2iwx�ʚxn'�qR@ܳ�w��#S>�wb0�e�V�ξG�n	�@�Lvͬ"M�h��SUmظ�zCh�gwFY՛��IݤAiw~�R��U❅��n�er�$�GsǢ��M�e��P�F+д��P{��6�v��j�e�jH��:J�$"^�U�b���c��<�t痢���\�|`�p.Uv<(��1rCGZ �D�my*�1������Җ�jxi�n�n
����z��J��;�-�"��+��|̋��r4�C�5���5�dp;ѩyq/��M�s���Sp�Y�f)��+�d�q��/6x�F��N��= �r*D:*�G{|��O�������{=��g�����\��$�J�T�
�x]Y$|�Ax�k�5ڦ]0�"W^Q�qqSQ�K�2YW�#7`s���@c;4=�֑)}���8NmLH _B*�P5����9p�=:��+���`�-���e����� ڈm�uؓ{c�ڶ��KΡ6��I��0�{ �Z�gㇶ�r��c] �S����V���s���Oxw�&�����0�16.CEHE�4! ���e��5>�%�`�{�K�:��\��e[��݌�K��Gk���%�䲫)M6BFjoxj��jFndZ���tCq̻��/'ϧf��j]$8�ڶrc@ty�:aP�c���2�u@d�q	�����{cu�[n�]36�|l��������L]t�j碞[��V��H�wy[jic���A�(�[����y�.�J�{\��� ��5������l�3�����iŐ�=ԣ2��|��9W�h �
x{2*��c�X��ӝ���h�/u.�\a�{�ڬC���IV��̽}��|�'�5R�"0�mq���[p.�{��Iq뻩����������S��D)"&�aYR��f`'7��`��۬<��<�ƻ2�\i6*�t�����,x	j�7�n9t���4+ٵ�Q}o�ud�%�N^�5� ŷ��ʜ�:Kn<���tʆgR=W���lf���c�n�V�|��%Z�(�jW<H���~J�/F0��9�|��;WP�»{І3>R��;Մf��)����W`�X4i�:��דD|LYոAm�X������ma�K�������ݦ����޽�|g>�31�SI��-����T�b؈��N;����c��2!rd�"Mc�,����[�݊�)V4^⽝MG��q��Q����8���ͳc\*J瞺�i^ࡧ���Tu���VOr<w� �X7�WU����m��]*��L⥑:n%#+G19���l��mj��¥�ph������VI�z����$�	�t/�Gx�<��`���.�]P����c�[���嶹�7������8���W>����u'WJ�S�6.���d���ÄD��f���7s��ٵ�@#�f���ַ����1��!}s����h�����:2B�o4���bG�lX;��W���wb�����I���L��r�x^:��\�R�B��#V��	sWE��op
�S����K��ʮ�˜c�̾�i�"QzM��2jN	�yl��w��L��{���i�(;�'qb"������ۭ�΍����֮�q�]&��$���f}vM)QR�����n��RތȦέ�AX��d�\��D��7v��p�fgh�${���JP(P�ܮB����
�`�.����2\��:TW��uF,\�(�p�����sc�F+�1ӧ�2;���X�d�]�k��#�e����D��`�SI���x��ȋ�Y��*K�$IS��U����sw\��sQW9b4ww]�bѺ�ݱh�71;��b]�Ҋ6�ӻk� ]�7"@��u3���9��d�s�k��jNl�hѹʍ%�w.wd�˘%0bH0`�wD)s�Qi���K=w���&(���(㹜�"Q�E�Iv�؈wF�1˓�E�fFE˄"��Qh�9�%s��1�I3�6���3ID� �2wq]�(З.��;���`�)� b���nnm�FC%4fQi��k��h�d���H�B47�y���߿��{{}�||��p]-`�����]���-n0�G�e�و��$6*�!��e��og2x��+���u��gޙ��p8�T$����c��t���%U���W�0��P�TU�U^��۷��f0q���L���q���'WgCf<��Hk۾��B{<�g�?ϗ���S�)�
<�P�K��>�Y��;%r��9�Y}��(5϶�XS� 9�6WTuOv(��E%Wt]+i	�T"-�2��5���Y`��l�!����3:�G4`�iK�1��H9R�{,F�gv��AjH����y�̀��������j2��	L��O\M���W���N�}>;Cg�7@�o�C�"��e5ikW2ӛ]��mx����z��^D_��������c��h�,��e4Uf�Fe�ՙ
��i�zޗ@o7G��i~̈́�<�tQ�c
�Z�kk�s��o1��
}3�C�R��^i�ydD�<$W�������!��1���1Z2EY���q��l���QR�!�j������G��K�8KM_D���:�髝�N{K�l���i'Ҍ}.ˏc�r�G\�qd��ކ#yzn�mX��>B !���!KFKÆ�NS��|4�d��ד�3O|��si���ׯٓ�䫋}B�"�U#�5uxsV��M=c5�7f�"�w_��A���dj�RK=����=T�Şѓ�������T���������T�(�Iꊉs8Yt,Af�0�2�jz̹]G�r_�Rt�5+2(��3ʫǯ$t��� y�󷩢fÞ�J7���n�0H��b��뤕��h���U�S�n��(��|���2;��- GO���e"�"=\c6��"�s�K�V�����&ḓ�s]ó��FY�u!c����9]1�t���*�i0��+�3oU���n!�����S�ځ��flp�P+,?�#��5=]�Ubj���/Yɝ��X��!��gt9�����NhHa��a���,_��u{�k�E��M2���Ӣ��횗e��ǕZ�1wB��Lq��7��Z>�7��~��+?�d��ڶ��n$��Ƙ�|O{���e�E�#�:���� '�wf�Oe�'V�=�P�U�kV�4_�C#�p��}�X��굆ps�r��{l�]F�3;	����@X�j���oO&�%�����J�	�b�k{�TGl��}��z,VVoLQ#Ԕ�� ��?���iS�r�VP��J�+��6��n�U_y��5M	-|{7�Bd8,����&-�P��4u#A?NV��ѳ��d���8�]�=4�?gJ�\�*+/�-�����L�<[�TJ~
j(�L3q�뙊�؋�w���;$n���3��y�[Te�6�u��B�lλUu_�/�v(_�b"E�tN�?fs:�a�'ٹ�f���ۨM\I��N�wh�o�[� �"@=ɧכ�UOC��I[���Z����G;��q����/	Ky.p�V��l��"���`����Ɖ֔*�iy��`틅$R�J�Ɏ��<���ʥ'�Z0��⫶q���q���w�X<�F��m����$'�H�^.�΂�0���6�֯XQ3{C��n{�WGQ�s���g��Dc�V+���2zRM��Z�}�-]�h�U*z��n�]5�`�1|E�����S�ك(<�6��.�y�Ƹ�����p���\~�0=�ޜ��k�th��\L<�޻�e|6ظ���um�k`��a;�u����.�^�;��1��&�����ק�I��	MJ�G��|K�\����/'d�? �<���N�Y��[Bw��d&}X�2�T�#���w��N��(�h�-n�mt��l� ��d5!-�FCr�s��;��"W�nMv'�QZ󦎤�!q~���v����v�H7Q=W�4�56���r��_ev��\Qy����;�mt�L:a�fD��D`�O{Lxf��8[ϱ�t�~��Җ�D�T�De�j[l�\��Wӎ�R~��:�1��m�ޕ����s"���3ZV���?%��ɿ���V��` ��3��Y"���
�Ot�twd�n�ή��B�N�)�s��32�3���C�7��ÆZ]�^�xn���q�b冢I(c�?�O$�����`�;��ڂ�fV(�O]bf���/����k�����!t�*�Љx�e)�<ޮ�J���A�[j~���O"1��7ɂ�#�]�nm��:.u���U��eM8�sO)��
O�N�y!���^��Z1[�ra$u���&�:�����=�y��@��a^�Q_�Hp�����bT�Q�ȷ��������WΏR&� �W���Ԃ�G�z�4��v^2#�p�G�>��^�O�$$u��	�J6�sa�í�U�7W�3^yU5��g�p,rk�*m.�Ln�5�U��n7���%�p	����K��iڢ ���ߠ�\ޟm��\�y���������lWgp�W��)T��ʹ�n��l��\'"��S�n������w�ص�m�t8�μ��0�GƟ�IUځ�N�K�]�t)[!�acr���Ϋ���kBS|� �)+뎴v N�=g[ �S|{��0a׮���w�`�
<�v���/�Hɣ��(�ʗ+O����ȃ&��Vv`g��#Z�st0������.�S�;ϫ���)(k���:�8�Mi�Cm��Lh�]�Z��]��t ��Ϊ�p�7Nq/'��#U�%��;�o1��9P�Fl��{����we{��i��N��r[.�u�f��B,����q�����i
�vBW�����B�m�GOa-q���n1D��a��7N��Vf���gs�]"q���G�BV%���ߐ�o��ү/-f�n������sd쾳[R�<���t :#6^fqk�J|�3���ʓ����T ���7�7X�6��ճ�JS�x��X�s0ʾ��g�	�)�U";'�tz@;fz��;-Raƻ�j�2-T���ۊ�V0gc ���e���n�7�4�	y��y�ON��4@����y�NQ��/Z+�U_��:U�ڴo٦����Y�Us��n�oC�YyAE��V@B�=�5WT/�H��,�AuĆAr�sg@���h>~�YU:��{�M3ٽ��=�ti����V��#����o�4T(�O�ꊉs# ��btq���sWNuo�|�%p��EzM<��^�OM���3��ˈ[pԼ9�]AB=ZD
�5�J��%%��T�K�'���1����6������D�������D
����=~x�l�T����٣��_P�9(v�����K鋸N�0#|��򏎑��շ�����&�{/�pڗ�Ix.���&��4ev��{��f�^�f�>wz6�v�5�������13}wZr�*�H!���=Y��ӎ��;�4�W�5uC��y�3/q�{WU7!]�˽��ʷOb�G}�r�T�2���tƑ�/����(�NSX�`�?7��)?'����6���<�����@�n���٘�Ȼ	�
kh}ܶ�-Y���08z=6ˌJ�y��`�q�o�H}[��l�=OE�;����K���F��w��;�*�6U��u��#8#y��ahim�9W��tO���i��(:W!v��Ǻ���I�P��;���^����s�pL�G�$����)I'��Ox�i��Ḻޝ��u��wX���g�YH���<C>a�/�F2R/ V�4	�3��j�j��M�b��]�Tk" ��3����@��1�E��۸�N�Rf���9��o7�_�F�p�W	�:&���_5�a6�����n�\���H����|v|����l�ӝ&5�C�>?V.�/I����[�?��6�a�xӗ.:���3r�ҋaX�`�r�:���w�6E/q*43���L�]o>���(7=[W�C�j;Φo��y&ui1��5�j�������S�%�zQ���=xٶ��-�iڮ�ӷ;)Ҧ�t�s-Z���3�o�.s�4l��7�^t���� R�%u���-VM�����n^)���5L�������c�\p&G	q*& v���H��U)9�!�/04n���y]�w7�Zl��uV��:�NT$#����:�Z]sK���&�꜖���w��w�R�Ϊ�|�@�e4��#/�0��#q5��];������Nn�Y�Xg�q�>�K]:�o8"�:+cx"�(�n�SS���0�~����%_*E_<�����]!�o�PA�k)ѥ��Э���v�s�^�`��IgT-�������H�\_�x�ۮ����ۍ��w^�?w7`\���:
!*����s�Qy�s���eaM.�e	g��5�,�[Ѱ��3����.��l�)��收�&�g�6�������9�g{%�t��7�Ý0d��m��J�������e�����9b�m���=�2�5�G��t'P��3���y�ٔ���8�[n��/�G����x��t�\�-"�L�D����H[�+f��d�D���B�,��X\���Aؗ\�٧]�a�Z�u�6F�$��μ[O$���w���d��e�M�*<�*A���k>��k��M�{�^���#���,��U��3t�U�$���:�����-٣�q�'�5{�|:�-����~����{�4�q��^{�1����[c���I�A �s�	7�OӐ�+dN7��h���z�5��#Qה�g=]�{�V�%�2���a�pEwm�����&!/\��u �H�tv^�H\��C��N�ii�{�q5�K)-�-Q��s�Y7M��qA]�Z�
�H����-M�2�$�j;�`��b{\I�6}�ب���\ә�*�
� A�]����Bپ�u��{��M���)D�	F�XDj�Um~�\'"�C(#&"C�횗��E�3���7w���)*�ڀ:�֘�w�؝!���N��4�_H���#\[:/ȔtU{�L���ǰ�{<����1��2�w�3�Q�&�Z���(ٙ��r��קC���<qi-����W��P�0�;�1��/.CNZ�ر��φ!B
��s]-���a������Bt�4��r�-̬d��.��+����ʽOP�@��j�KL�^i��٭��N��nn7}��������r��6k�ټ����`�m��=��|vT�����C�ޟ�\�1�/�ȮZ��[uƱ�I&�F���^%+��`�m��`�.2#gUG0��g��]�=��#�܏�R72o�~9Yci��� ��pQj3�9vӾ5U��o�o<U�yF��]I�e{�u9=�����w���c��T��z�)�/��e��譡�o��]��@�T��1�d�CW�Y��^�^�����k6�ڣx7��p��R�����m�g7x@�jČ^2�{��9�ƛz�X<?����d3��S p·���������"O�7S#yB���&i(��M�]�Ncǹm��}��,�(��/S��O�w�.Zk�U+���������>&Ȑt8��8m�������y竽����������v�������m���k[ko��߿��n�ֶ����*�z��+�/]�mu�Y��5�6ٕ�-S+fV̪���j�m�+fkfm�6�5�*�[fV�+fUL��[3k2�2�3k3[3m�kfmfkfm�6ٕ�5�6�5�6�elͶf�3[7��U�[3k3U2�e�Y�����fV���ʮ�Y��+fj�ՖZ̶�]��5fU���k3VeY��k2��ٖ�5fj�ՙ�2�el���Y��+fZ�ՙVf�e�ʲ�Y��5fj�ՙVf�elͫz��׽�^�m���m�=����m�f���m�ej���S6��[UM���V�e��f�U2��3kZ�Z�3m����L�U2֪���޶��{-U]�UL��fmUL�m�5UL��f�m�j�oJꪦj����f[m�*����fZ��j�f�m���f���ն�2���m�f�����mUL�m�+[3[3m��ճ+fUL�fV��̪������޻zoUS+fV��fV��̭�j�[2�nn�fkfV��fV�ڦV����fj��>�+��]|?��j�2ڭ�+kV�3_������|�w��R?����_���|�{���$1���
��'��/����/���U[m�/�_����_�kmZ�{�f���e�u_��e��~�U���M������ѫ��U[m���_�~������]����u�_�����k�ڮ�?Z����mV�m�ֶ�ڪ�T��lUUQ�U6m��5UM5UM���-�UMR�m��j�j��T���l�Z��eUR��m�-UJm��յ[���[[ۯғ��������MV������j��EU����w������~��y����yW�_��Um�W���~����/��������>5�_�_����~���|���:��~��UV�~U�j����E��k�U[m�j����Z���˥m�km���޾)V���ޥ]�?��W�{m�_�����W�����_��^��oj�W��mUU��٫�?��?=UU�߶�tU��|}���/������_~W�_�W�M���u���o��_�o�j�����~_�~�^�k�����k��T������W�w�����Wᯯ�k����U[m﯊���~�U�u�W��U�_;y�}��嵶�m�;{eu~7����ڵ����_��;���Wj�����d�MfSy���f�A@��̟\��>=��>�
kIS�m�B�%IQWf�łT�j�@R�U��$��$����
��PP
V�%EI����B;#U�m�������UY��.���ّ�n,m��[lVoc�V&v�hkJ��wm�MۮJf�5��)e����meX�m��u�j�6Ƥi[j�Vّ������"$��t�S�U�lhՙm�i��m���i���Md�i�q�gK�F����l֦l�[T�Y�ٓ
��s;7n�h��$�:�t\۶廵u-�����ݍ�  ����m����p��W�YF���޷�v;��et�����ZS�nŷ���Sk�yyu����{]�:�6ݫ^ʫ]e�P��N���u�Q��hw��Y�Ζkm���Y��ت��  ;�=
(�2<ӽ�СCCB�7���С�z
(hq������{X������v=l�Ӛht��d�Ov���[Cuҕ���ڽ�<7��ht�{ݛ+S�w^���Wm{�����dF��5-�I|  �����Z�������@n�n�w[5�i�˦=ۏOOJ��軭n�D����X\�i�S[��====h��ݧ�JzW�S�fivu�\���ý�]��w����m�KkU]ػU�| Ǿk�vOMy�n�δ���oW�:�s�ݞ��j��LAzn������׎��4-R��{��Gw��zb��C*(�`�U�͵�w[��nu�S���f1�gU���ɭ�����Z�Ӛ��J���m�h����(��N�m�֟N����b]��h;c�����5{n�N���VҫmL�ڵ��5��N�o�q�CK��R�ճT��&��UAb1F�U��s�T�Tw�����V�]:7vָTL��f�:�;U�l�ֶ�����	f�B�ωb�7�N���r����Yu[4�wj9J�lj�(��6ö��k�� ۓp@k��� 4����S"J��6���h-�π =�@��c� ��M V�p  # ��  �j� �,b�N�u� ��j{kKM;n�����P��%� �� C�sp6�
�� V�  3+ ��V�;`c�  ��ph 7.  ��� �z	v�kY��)����k'�  ��  �n  ]&  ���z � wa�w9�  ̬  ����@u� ��&� |���R�mG��)�4b��(�  E=�&���   �~�R�� ���J� `@ B�	���@ j~�?����W?���:*xw�kx�EV�\Vd���{�Z�w�wg�����
�+�_������T_�"*�j
�+��*��APEeE<���=`���/��.���_�x��^��p��1%�&��e��"�I�ZֶQ�J����c^�4�aUԼ�dȲ�-R��G��x3)��3L`)��T���3p�[q����T�a�2�"R��0��z�;P|7&I@:��J�L���Q�0ңy��U��ӧa�!%B�H�-���D7��d�$T�A%���\���?�����k{9�Zs�ua�VrZT7n��/T���/+M�  ����R��*��ܑ*9.
xa��p*����a ��r��j�^k���Ħ�r�*IW�2Iz�uu�n�
���6*;�-,�	�K�37!;�P��(���ڢ�;7����N�-�A�MіNє�;�9P� ��f�y��7p^�c)D&��5���X(��㨲�7ORJ*
V7A)p*�@�����@�\ܫW*�oOt�}����3-8B���{B�.%	3�Y"Y6wX���v�VQ�Ҩ%�ɮ��|Ւb��^��ú��r��4���/i"i-��ϰ�nʋnԗ�)E ib[YHѤi�j� L[��Z�"Œ�O�Z7Rz(1J`Râ+n�T�Ǒ��V��Ơ"�q�P+��!�K5�憜h���	V��Pb���ܻN�*�@ֽ-�V��`��
�7Y&%h�f�^��F�$:�Y�g�Q5sh��c���k�y�հҴVb��p�.���15a�V�&���3����;n��	b���)��Y�7���	�kt�kr
���[��ͺ�Z��p�iP��F�.�U��4�tsݎ�0'Kb8V��(�gJ(}�A�:T��Y�|������X�]DA�j�jB��f9�1���sql�u7b�%�B�(/ _
ARx��t��$:�㳛rЭ��8�8K�����-�[Yf�*�tXi]�X����T��Y�ym�T��4�B�u�"�Ej�\�?���k��]�V��R�4�ȃ\ڀ�Tҭ��mu��V�$�ajhF� ��Zȴ�f�H�tmbzoO҅Be�vpM����F���	���d��RL.� @�fb���Nk�����m��F��SM�'z����TJ(�5⿯3.����Y�`�j�n6�n�QS��+H�5x~z�30�,��kB�K�k��/4�����)�%���� F�Y.��(�ߡ�31���ut��i�nm� �e���i�q��.�n�Mv��V(LtD���3@�{��s4ƛL���n[�/Uj�;������^�i�ZȽ"��� ^�ħv^��^e
a�x�x���C#`VV��y�mX�B�6,�[�rƽ�C6�3P`�3v����_oVS�r�I�B;�+-\�����q��r�ݦ�i�4~�.�̭��Sz��N��P#*�M��d@��Tqe-B.��M� �-����n-і0��q=��N�^���Ѵ�M�i��j��'���%I��QIVٓP�d�&����|+�$Լp�z� �x�̛���kܭsw��y�($ E^jH<)��<�T��T�+��8F��o �0�@�e[���7Au7�,-յhf�a�T���E4������t0ZwZwk���/�D;�7IB��PT%�=�鵖�­����9�D'��^����]�Tk��*-�E�ܲ�}�,(Vu��$�.;��Q�_ ���F�5n��t��%�b�蕤�&�d�a�F+
��@`"G��� ����B��X�j�$��k]��.�=*��e�f�B- m�wD!��c6Ig
��C��t^fs1M;F��C��F���l1f�Pӽ
^��(�u�ތv��!ՆQ�	#[V^0!�f��٢�$��a]�@�2��%]Т�X+owP�nk�C˥L7w�v����Y$Jl{`nދ�V�X��L�8J�u��^"&�F �Ǵal��ktd���n�A��n@$̒Æ�6���5uo$�ol(K�.u�E)zՇ�f��hqJM�5�*��֦�w��W^Rی&ueji�g4	��B}{F��vE��a��`�a=7�-kBG�[%*� xsP�3^D�a&��jd�:u��'o�W�ya7Ovl��%�[30�B����^�bKNVi]Z�rTZHc��ʺX�3�!���o*|�·2�F�ͦ�Րc�6^m�����/^�ڶ��3TC7@j�oI�[0�Nibĭ�#w5�pLf��^�z��b�/q��WJ�on���]$a�,��(�NF�GCCjR�
K��2�ݰ;���[B�&��F��l�F���]�|WY�������ŨMK��V�D�@H��n�	�3�^��Q���C$����i�WOUܚ�([%T���F
't"�i��I�]A)��{N�fT�4lqȷo!C|�IQG30ʛ�X�5��0��c�w*Yb�=C�W�c4��%ꢅ)r8Q.��$��87sB�	�+s�Q�kF��dB]ʻ���.f%��d=l�!��Ҕ2�[� ����9wHS�çr����T�/D�)y����tf���Zƍӣ�
9�/vn��`-lh�a'��T�-�DT�z�)X���'�����Ӎ��I��Ƭ��TM��� �o���K��y����(��,���Fvq�\R��x-��M�E\�wf�Y7]�G'.�6���Dr4�U�[����/#B�Ԡ�YFk��w#WW�_:X�+^�ԲB���9Lm���"Ǣh�/]d��b�TR2�8+h�lڎ����&YP�Z\������e�]��z%�d����Y��*�ָ��$( �v�fPt�Ya-�zkpAr�8���l�~71�Ӡ�3~H�[{�vAt�L-�F�f�=���[P6�w(tD��F[�/@UiRZ;�%R����4܈�'�v{X6�`�)��-�*�U�͵mU�*��FQq�Sm��޻îU�m�4K�,�,�b�iG6襆�&1cnmeV"K���st��H�V���J1�]iM���!^���#su3>��!���gf�%`���1����d
o�5s�Kյ�ʻ�'Gh!I��&����ĥb�u��Y
�Ӂ�hح/n��D���V;���C��F"⧠�R�ɉ6�Q�-��d0�y1ؖaZ6�L�M�L�4���܆]̎�����㧛)�2�,��r�2���I^˱ji��P��Ff�Q�V��)��^L��0��v&�2ad@�Tt[)�Aj­K���X�k�ϲ�.��sA׳Mj��t�l���%�Elye6SO3`����m�u��*�I�p�)J�f�úk6����h��e��4q�[�'U<�)n�C%"��aS+&*ti�c�;+5��BJ�H��e��,L[i��'�S�Z�����SH;[�i�b|�M���,^n��ImGw(��R�n����xF|�/nTkq��Ҟݧ���a��3�qD��2;�4���ۣ�,��X�(�@9�f�@���ʙ�hW[��COv#�L�ê���׭KR��Ö�E������ʱ���L�6� �B37d��mf��/t*߭:���,�YLͣ�%�� �{�]J�c�uۭ�Qܔu]�oA*�]�0c�5�"� �m-QU� EZ��[��mFvlxR������bz�;AfЍ(`uʀc�;n���\B���B�Ũ���QK��Ef�u}t8���q�w�Y*v.�4��J݊�t��P(!�jo)�D��5�B���Q�R��wS2��z@�{��U��%[�1n��W.�zm�ȡ���*H n���6��gSΈ��ᩢ�d�"�p]��-�H����r���C�Yd��֬,h��eٰ��ś�j��Ka�n�@�iє�N�f�:�J�H�gw�O~���Y" ^�բ���Y��6^�ùI��I���:˘m]�n�-<�ڳ��6�ZM��!�l��<�c�t0Ѩ�ڭ��ˣ�r�Kp$I���j���F2���vT��":w��R���;4<Q�`I �^��mhN���yK�I���\��\IL��r��dغ,�u�Sj����ʊ�Wi��c\�b����̵�3A�ˇ�M�EP5��iU�O6���ې�E'����PL���[5��:�����&}��n�����f�1M�Y���嬘��(�ݐ4�(���v�!�zlMÇT���T��l���7ccj�"��7$�X�#\���^�����u�H��XM�^Kq,���Tj�Rj
��{�j�UZn��3 �b����(S:�BM�z��L����%�`�aC`3Rr�����Zv�kJ�JڋZM�v�XyZ �Q�@�B����]ZG@�6��L+u�&6���lR�ab$/>HPI�O-��ɱ�AgR�2c�[y�w�hR)+N����.��2t|�f]���n����5kD/]RKe)s�+i���ըZX1I��.�H��(�h��=X�YԬ�W�J������(��R�1�W�̂���m�{�f4�S�gjb���클����1Y+0�a�(
�B�t�,E�jV�Y5�����cAƳ�`Yj�^�4g�R��Aߤ03���k6�:D��=ԚuzX���SL�ܐ��rmm#|���D�]��1�սZ�T&�Z�fDwP%F����2�p��^���ܥ������J�v�{��=w)h�Z�2R��k^�0��f7�K�i����,�2�yE�2b��mZ!)�1&U=Gb���lHˀ���w��:5�٢ڤv����mK0�n�Ͱ�l��VIJ����Ah���70��<����rƕR�U���КЩ�b7Y�ݥktM�E:
��1�2�"���FU�j��@Rؘ�IiJ���n�ʵ
$�����۫����p4�iչul<Q��Q4qaP����C%��'�l�V��bI���0V����X��$H��yzg^��A@�ZK˙���JV�f�<�ILI�y%+�
[/���i۫&7�Zۤ�Jz�ˀ��@��Lkw^�6����a��,�r��%!��(n\)���h_ڋ��2�"�v�-U�R�n�>ef浚�I4`QR[��qdu�����[Y{��)I���F�
T���E[�^بrbO.�;*;R$<H�km��N�ø�h�B 0�lQH�T��e�7��oC�Fd���zց�S�U��)}�jB[{w� �,�ɶ���jhkw���q<z�0K�Y�Ь��1 �^d-�62� n�*�DMF���nXw5%;т=�n��)j�Nb�Zy�5|�Ql�򲣸�̉`�Ty��wgCofOR�L���*DkiY)�w�.CB��ڷ[U��0\3D��̕�Q�^+�E�w4nEt�s[�wc�ȱ�N+r�
��$�8 7*䩩�D�n�0�Z[�Aⳣ�J޲��Yj䣨bƃܐ��,TA�w+l#	��ӫe�v[J�1鼱�����6��ʅ�<��j��)�hL+o�A\ %�mUH�CJX�=�72��Eۺ���U�Y��ˎ32�%��S�Y|���XW��1)} �Ћ٨�V�p�Æ��J�Z��1`��D�,֥��1�e�F�,��t1J5���۴��i�(nU4�\�"��:%�W@=��LɚC��夛ԭ��7	V�:�"�ԃ#7Y�;���?eh��]Y�Z�X��V��t����<��t#)h�n��һ�F��3Z���n�Zk8�1!ulKܠ�5A���Z� "�ӻ��**�p6�nnܡ��6���rVY��%�����
���Ց�  �Ev@5y�m�K6���`�L����E^Ki�y᳭�RTg&�F�cqG���B'6�X��x���͊+V,d�b�f^T��R�U���H�[*l7H@v̬˅�B���a4n�t�%�9)a�ӆn� mz�:w�^d���6E�ML1�,����F[�3qʂ�{	� �S \a��4ܙY����mB�4N#�V��, ;)e������1����Q�A��n�ga��P�ssVRe�c�%	�ݥ���D��f��]�(V�ִi�
����E;����ujn�Bf�&��!�w�i��M[*Z�{4裔��֛��p���:@�)�e;l���gR�0�z*\�ȡ�� +X-D��5n0��5�6���Q&}{���K1cR�͢ʷ�p��(n(q��iѱ��Ī�1�ƅ,�N՗n;�ԣN�u����@�%$jP����wǹ.��f�Dސq�aJC0(���
�c��F^'�kR�B��F6�f�jV))��Xհ�A�����b�1���U'{.�_R� @Ҥ���.͑V¡A���6�fü�Z4�� �sl��F:T�[i��0R�Y���Ҫ@��K�����T�l�������c
�T�a�^e��m];���s�N� ����͓њ
B�R���Q�`b�V�W��O*��v)�����0CQ�k0�F�ঁ&l�mN�˛ˬ�
P�i��4<��TI�"��,��w�p��,�a�9G3m/�^'�Ȅʲu��ת�А�:'H(-�u�ȩ���mI�U�2B&K`�Y�B�ɀ��٦�;�4��`Pn��R��j�Df��j��3)ǟ!��`@bz�D�bȇU�N�����;�7Y�*�WK6$².�����4ٍ��3d��l�̴)�*���b���i���Ƭ���JJ�ea#�QV��@b��E�&:Lbb�D�F|L!�X7V�	y�x]i����i��X2��.l�ܛu�:%�H��M�d")��r-IP[�2_Js�ʌ���Z��Y�g�O��`��zQ�6�/:�Ȁ��J���w�]M3E=��|��Ud��e\�9G"܂t���c��a<7�,��G}����'wh<Z��1���I�L-���ۨ�]����/B�#���iZ{��n*]�=c�q���w\bה�)Xr�pG,�=��uת�I�� qdJ�WE��ab�3_���6�%F�>-G���	i�*��Ǯ,��ե�����83)]��%���ڭ��K����Ϋf�W} ��1�b�0��wxF��[���wW-
U���t��à��q�����Ua�=V�-~m�`W,Wѷ�;b��o0���J����R;<�t����@fL	�m!�䘶+�d�Ŧ�)r-�Δ�\��m��4k��*ɢ+�E�b$��c��{���'�eε�+ph�a�ԷI+���y�	��������ڴ�T;ԃgb��ՙAn��٤�T�5�Nq*�wCzƠAǵ��r����CU�q�mc?E�ޔ�%qy�s�̫&�U6���wIe�{Av��G��0�G]B������Fi<��\ߥu�]��H�,�u���J��['m��Tn�(��*šӣ0/�[7�g31�$nh{H�p��WyP����/Vih4�.����,���ؓ�e�ޕf1��ݥw[Hr��㖝�M!��J�	��E� zU�[�j*���Ǳ\
�j>��U}�و�1�ze�y�)����Ez���U5��L�jg�u>� +�X��[&Mk[N�9�)1�g������T��j�M3��H�(;����n��T1>�9A���0c���RϺJ&Ҧ2KEE����l��֘ԡh���K�(ܑ e_
l�3z
��k�z]�͕{�8�Q�Tݺ�{��i8�$�w����6�ؿ���s0�Ƚ��]KЭ��˖��7A���5J�G�:��CZ;6\:s	Y�t0�v�8������Ѭ��qvD^Z`3�����Ptض�z.���b�5������lu�-�\����yekUb�݂� {�)}*K�f��������,X��\H�4��*�}������R�D	��ڄ��T��+�|*ned�.ٹ�ʂ����ȇ�(�f���B��/�8�.�`U�f2pжV4;���b^�ESR�d�m`3.��{�j�����*�zh�S!�������bz8`;N�ȇ1�n�WR�h���p�\�i�m7�Y��E;��f/U�t�yȧ8y�F�J�,Um,�jj��t�PeC�J{��m�;Ej]��M��P �K����&�Q�b��X/�v{�����Y㛂����Ջ�ZHY�*�jsd��3��"a�l�N�\fWYu�V1>C0���uZ'G7}MqL:f�h��	NW�)fPV�j��q|�����h�+���Z�DR�������Z�%Qh�]
ά��Tl�LS��S���9-�3-�7���yia�G��(�$j��T��WTӭս�Hm�p�V��{Q�򱂹hԃ��o���jmj���/������ o�����U�e�_)�ޞ�9+���n���ˀ��@��2�2���iD:�ZU�.�M��WG*�+PLnv�m�\x���I��7��?bokQ�+g�\��V���4����.XWɰ�	�M�n�*V��\���+�%7ʔ&�&�����g1ҹ�-Qrƃ�d��8.7�6<�P���]r�o~MV�1�p
b�ÁS���ҫ�/ip}���_Q��N  K���-�\������	u�u��:@�������+<����༫ý Ʈ�, 8±�f�	!q��V�	��C�x�qr�eE��;A-�n!X�L��h��PѸ6�zb�t�"�{/��9�&� ���8�7/v�2"���׷7���8&�%��+t(��z%�ͫi^D�;;3#ja̠��qn1���;�� ; c�D�9�p6+4*d:���zL�P��<�����͚�V��6Qk��0����/�m-G��J�a�M)$l�����j{\CR;F���eX,7���{.]Y�T��]��Nta�N�D�z�$�/o�^�&�]�ٱ���i�]s��9H���z���%᣽i�2Ď�+�%r�I�|^�7z2'VbW��du��5�'S�L��3�-��Z�W��,39Jgo�ۄT�[Q��ˮ�E@U^.[�_��r��1�b�7��4��[�0r3F!X�3��Vwf���c�)���Md�3��^vdE�F��7xs A��6�\p��Y3��a5ԋfVZ������/qWY��7W�q4���C���e��Nآ9Cv�Ewlg� ֫d�ȋ*��{��ڌ��W�q2wUی����j��x���H#g�j�i�_WQan�W�C*���U�/\g^�NNe0��u��z*���o���ĥyz}{����|������N�F6�MQ'a>f,���ve*8�[r���Uܢm�h4ҩK�x�>���]`vK\&PZ:��^#�#�D��[�V�ya�5��}i�Fv�0u|4-X�S&��x��W$�:���X�jw1뱮)u:lֺ��o��kȫZ��J73�<Q��V!�I�_�輽 ���բ�|��N���U����E�(�
XR��p�J�nv��1���a]]��0����i��P�kIa]�ݡ��p�;\9��z[遻�WD��-D� A�n���h� %���i&�;i��7�wj��߷U�t�܋%�
궓N��N�o�@��K���2cq�b�N��ɻtj�y��c(�\(^��]a%�����b�+KsNæ�q�yKD���M���5"���&7fwl�&M��YV+o��C���#�����-ۨJ�W/�&ٛ|ё�q�K;Ƚ����hW.ɂ��d)ipX8i�Q+�pJ<zc�n��t����
E�n]t�����1ЩKyE��wׯk.�j�L"^#r�T�9��3mVe8�Z��1��+㢷��t��Z��΁WD���@�<�՛�ڼ�D�:��4����p����4���|[��*�h4�}�0n��,_vH��x1LHd��r�8ݪ[N��Q��#�Eq�������8gNM	V�//n�^��v|E���#M-�z����]s鄐R�t㉮F#:Q�<֎���
 uLw���U��NϠ-����ےo<ŗ�l��0�fm��f����ZޫM�"��ޙ�-f��6k�������ֻu�;9��	�W[n�%sy�l�Z�d�Kh���KhY���杷�Z{r����Hn�a���������3TgA{5jm�39h?��X݄�\ˊm�y��J���Յ,��Eeug_5����I��&#ջ `=�����E�B�+�o%͈u�BYׯ�7WM�ci�k�6b�����kj1��	y�p��ם�f�XR."/K1�u��Z'k��(沕gEX*dN:��
�ڱ9� ��ڛ�{�u���{
�A]i�f����d��rI��G��w�WzU<��ͨ��S��׹(�jk��kZO�w�S)Z�饅��
�X{��)Dv��5@�W3E2N�VpQ�:	[�OZzI����b7�h�R�ݰ��䝷F��@z����A4+�eC�*,�GZr�E�[-����,�e�Qw1�2ݬp�^>�ε�r�)���aQq��
k����=Zs�7w�h�7!���Ir��74F�b��%� �q<�;�U���\�cn��B��ݴS�4���gp�n2�j�����m�B�L�)_F;��u��W��,M�/����b�& ��y\��2���	J�;�1a镥e�W��*E�<�3��U�1�D�v��T�D�gsB\W`�ʟS\��Flv�f&͇�a���gI-uq��1��#C���>��Y�fn�F=���U�9�p]cO�ȵp7�-ݴ^ޮ���h���}S{�X���ZW_ݽ˚o��Ib�Q`�_Y��2���U�n��.h�/00�1ӨqmIy��m���/w���rtS�JW�|��FݚD���oV�W��ǝ�4�x��]�6Ш��#(��(=�y*Snȧ9�4������������� �fr��Z����ox�j�7m� v���i�0@�75���E0��N�j��;x�m��*]��LА�\)�59EN+�d�jC�k>�:��v��	�I�j�n�)�2T��$�<�NŊ�.�͛M��&��P�M�9�ԩ56���2�K��>(�n�[N�Ⳋ��I��0>�� y�D�B�KH7� ��SfϦ���R5�سlkdڬfK�\s������R�n�.?<� wG9�f��ߵm���H�ƛ-nܥ^Y��2����������Hs�\rU��1|��fM��N�]�;�����I�Lt@�����Ҷj�i�|�Z��N��ǎ`���,����p�u.]�k�v��]��Y�\,��R�a�듷��)ecQ����sX��br� ܜ�*���0'��mp�|��X8��Y�*5����&�qqn��Ǟ�O@����ue㣵ur�wu�2�A5F @�]Ȃs��z����l;E��<<2�M��9��ʅT�ɲ� ���VmQ���-��O;llt'8���(��fh9����U
�QK�:@���r�gc�fN[婑;p�w*�\���w�,�]�;��Zn����4Τ�ѕ�������b9r��N�x�q���i�ݺ(���&�a�3�TȪ�Mea���yÒt�<�,K� ��Dˡ���r�=�Ā��;B���H�g��%F�Dz�\�X@�CEksG2\WQz�F���v�u��g�u�P6U,�ͬ��ʔM&D�w���Y�mV����1(V��a�b��U�W��:Ve$�we��������^ћ\u�T�ڗ ?L}�kY�Z+l(����X�ݕ�9Χ^��\��$�����q	����L�JK]����� w.폷RÆB/�B(���W�UԨN�ۋ��sNH�<ȳw�}�i4W	�q=
����Z^�7��ј���F4e�{���/I�:�gU��h1bogo$�v�0Ve�C�L6Q��ҽ�߀EOnz/I����������n��jh��Y��:u\��R�gp��V:�v��|�oQmuu�*�^�r��W2�%��ކ�2U�'s�=*̪ոu�"�e��a�@���2�b�q�˼+7�
�0B���Z�ϱ����j�fs��C�pu�(���}��jں��}!O.nHh5T��7sX��Tz�n��w\��s�X��u���4oe�P��<�;j :"s�Z�;�+v�U/h�J�VZ�A�-�°e��❧���2V����)iuW���7��ܸ�IX&��A}XDq4�%��<�v�M� ��h��sa��k�X��n�:����5��6`7qjR�y*EA���wl5M:�JX{�Q�z�_V��<�Z�1g#;��.�'a�r�ZWq�S�˜�&eb$�]ñ�{S�u�VU��	�Ī�Z�Άճ>z�������v�핑�&�=�̻h�;���5n�L�[�_ug�.�V��񼍢��k�2�_!w��p�m� =��s�(�o	+;���_<���)o(��S��es��v%���J���w4�����9�x��>��	m��'�+Y�F�Ȥ�و(u�O1&�+2Gn�.�9�#�V����h�I3�t]�#���[-C�S2���v�F7u��J�M��Vft�Z��M;.�wF_��);vJ؂��=�����^rn��FS���.eZw���a*��:��m��/<r�!bW<�*��׀8�ƔnT��E�P:��I��W�rm*]]9n��=X-Q�C�����K�ٜ�5z��dQ�6/:��)��ss��ܸ�'Κ��M-��������u�6b���ic���Iw��n��1C�j��.U�.�;�ۍ�Ki�9T���7�(���t�X�J�K�/n�̊��q���<Ft��b�]�:�5a�����8�:\�-��]�*6V �[F\� ;ӵ�{�Iv&p1]>��a���:A�r
��9N�����Z�E;j�CywY��+�ۉRc��N,oK���x�D����N����ܖ;�7,��ճoD��D>�w���Λ9�m��7i6&��%KP�}8]�����4
�t�n�ŵL�[R�o�Y4x�N�+���6�ZV`ͤ~�ּ���s
�M�limD����z�IA���H�Gܚ]l�ݜ]��κʴ�5�o�pC1�rch��~���/Q�NZ
b��q�m�$��5�u%� ;W�"I��,��{I�\:.�]7�dRJ���j���<7X�V���U�To'd���9Ҫ�'��gfE|�Ʋj:Y�9͆]�O��?�:��<�J��Id�rV֐Ml(�$��Y��c�x�k���R� �k�w*�	iW[e�,lXx��nlu
k��J�.(ڷ
���΅����/"��@�tŘ�J�Xx>޾�R�n9���ۭ�0/�����3�	�7!}��*��[I�o�XK+̢��ꆥݕH��|�v�8�&[-���Q��/�}��k���`��|�41!	'����U��g<�R�rԌ�[&���0'[V.s���5�9���.�t!���ݤe�=��G�E��q�}f��;���6�E�<�5�6>N^⼝�u��#PX�t,��_;�9�dÚZGte|�噽�vXX�KFݤ��B�K��8�s�����ۅ$�7����\KG�>L��?(Z9ɀm�7뚗J�]�@P�w�==��Ҷ�7#�эgV]���%`�޽��L�o�~��DU�h*�[�~yƇ��ZM��J��u���T����Io�9�ޮ�u9/0BG����*�;a�4.��A�6��h�o�e�J�q�6�e���11-��}wz����㭫�b���Uc	�)�p�@Վݓf�N�R�;r���AK���/Qr�YvشR�kFB�k.�ŝ{hz�:֭�p�K	���9,�BKuxY����]ڠy��[ILcZN"R����ѕ.�5�j�F��p&�nMW�����ne�
��.' }�,��;��N���ݽIX-j���ͬ�E:��; C�E�a��.����2�<#�\LĴ���0�5uv��]��Ue�f����7N����XxI��.'�v)�$`����e�V��v��F�׏��z0�Q��e���
Y�Q�ua�PP� ����Fm"x���`�p^�R��l��d��&�[�B��ze�ޢ�(�������e��%�j�c�<Dp)�����g���r��f�n��AP	�۪[W�1��R�l�%�n �ӯ�����.�����	 ��^_J3�{([6s��O�C�3���.�GB^��A�wx�l4,`\���V�Q��0ԮD�[�f��Ɉ�mG�b:k%w�2�Qur��LY�M�pJ�)����X��ҕ�	��"�� ����k9T*�z�
����S%��S{��f�hUrR[�.�:UcO(-d$��+�6�{������L0���7�A�[����1+����A>��#}e,�k�����E�S�S��U懙�I|��+��{u��y�-n\�gU)wQ��/N@f����bR�|;�i������D.�B�c�k����64a�n�M
�f�5`��u�.&�׭#���[q��r�n�u�L<��T��[�c%S��6Xd'�w�ZӍ�י6暲�v6+&��+҉ؓ��O�a�}VpMZ�I����l]�X���$�;n�*t+�3.�ݵ��4t�2�wI�3n�VU�f]N���͜Kl�.W�д���խկhe,0���ݧ�����٬:(��y}s���H�+s��^���m��N�!p��icx��TA�w3�K���b��<U3�e=6cqې�
[/3'>��.���h+�ү�g�h���C����.Ȁ�(�\���.�{2j�z�*�9R�޹*1�t�4o��d��nU�=2\�wr�m|�D�\�D6V�����ipl(۴m��o���Ԭ|n.
�s$�T|k9���i`���ϕj/���a|�����
eޝ�0����͆¶B�n&�)B�e�,6���=ܡ[�9Rkw�����6��]m�aTNl�]�Fbĭ��G�ŷ�	|�o.v��g�,�cOV���f��큭T{�)](��J���"V�t�c|�K����RZ�x�B�����
���FPuZ*�ы��J�mMt�ڭ���3a�����:阨�-vLbs��ȫ�^��ʎ%b�S�n�tau�����]J��6��7��)�&"�%7Z*�Њ���*�Vuc���ORSt5Zv,|t�O��m��4�z��Sh��8�Jl񫙦"�^��;b�:0Ko�9^!$\�HrEB�wD�VQ�n��;(*N�)���dLtV-����)8�˷4#}��ik"�-n������=r��`V5�;/RB�u������{��YD>�}��.���ᯉ����l�gq����e���1X��uu��+-�{�ɵt��x�1^�1v��T(�"��h��@���-��� 4�v�"w5���ڨ��)PJ��m�JՇo�f|7H-���n��h�����d�8rF/��6N�� �te�6���U�άAt*���ݲ;Ȳ��LZZ�]�^R\��r��{C��ؒ�i-�n�wA�����z�|�/oy�`7�Y�mg:QSN���f�v)z�}�c:k5pv{�^�U���sd)U�c|��fҶopڼ�d�Du��|��)Q���A0�|��}ܢ��q�z��|H�FTǃs;Li������A˱G�#�IP=�Y]� M%���<�1W�T�o��l�#LF/��� +^t��U�8a�qf��b���������m#i�}�X����V�k� X� y�����O����]$iMZ-��@��'z���5�:$.�pN�?P8M���˺{ջku��ԙj�3����q�If�T�l��G��U޺r��쀋��`8�7S������\�c�q�?�Y��gt+20�Leг[��Nw�ANfw,ڰCT��!�´82�'zt�����ʲ��AC��k�rv�QXj���C���̚�oN�l��[cU@*�%�e�����Ayꮫ��ʴ"�%4�7��j8G[�l�%t��1� [�׹�� �c��L����뺈�MP-9�;��nZ�K�C	�v�>$:�V!!�e�2����\"��b&�W�1o�nĲ�ı��єr�qV�o.P���5A�:HU�*�\���9F�ҴÜ��;O��n��4b���A��u�l��@ r*%K��{�b`�������HdCB�B���ָ�L�����G� �id�lR`'�_woY�b�@�6��׼�e����_+ZCLj5:�K��{Ѫbp��Z�.۵B(DBhi�O3]�1�YҥcDn��jD�+Ƌ�oi�jq�W�.�E�����[-p\��+����Y��nr�B����4���v����ٻ���'o���a�vr�.�f��kQ��P<�����rj�;�sꈝ�}�P�G��\�]nb�(�=,��4����
�B�oy,�9�)^�lX�*���0�G�j.<�R�)���E�8mb6�;�	�VWq��ʘм$��Q��b��.�:w{�s[��aLWiWU��r�.:�D�
�owة��OF��`���ו�к�|tn���/@�NJ�F��t��
4�jh��+hd�N��x9ha��W1�ގ�l��M�L���ܡM!$4���1k\�X5��/zU����C��V�؋
9m��h\��D�;�e5P���x��XP�Z���ҹۦ�����K�ٽtKt=zl*���l���YɆn�K�� }��k$G-�8Rd@(V_.�r���5�eڭ�ݢ�l �zBa�s�ë��Q�KL�\�݀�3)f��y�m����pc�'T�&�+*��@ھh�w=-u�օ�o%Rn�v����9�Kk]�|�p� 2.�x:�%�����+�bl��bIKff��}*,�{qP�H�ۺ�aj��Y������H
3.�뤞���u��߉��w��2��@-��h�{7����xJ`޽\Ue�.}sTuu�P�0���v���ds�n�H�����Z�ͫT����!xW�1�S땗܃�g-��q������X8�N�(���G��w�7�D���0jU1K o�W%Pu�Pp�=!/��P�R�#8\��0Q���#����5��]��W�������{>ǻ��Cسm3 ��]��9}�RqL�Wo���j��IaRr#P��ܧt�
�wa���V�G��"�Y�t��m�sm[km]C���%�A������Q��A�S6�!Ch��/�/ ��,��Y�\ݽP:�;��҃ʝSpX�P���y+��h_+#ʕ���%�^��~���V�ue�eSMjQp>)�xG<�D��(�#[wܰVb�T�Ev��t�G���8
��;�����Cw���0�7nVv+�nƔ����*�`��k�:����>�򛢵�:��w��4��6�Y��b�E���t�[��:b)q��7������V�q��nN�AG(��zC���#%��c�#�{�F�ʍL(�^�\-��X/�V�ղ�h80��NT[�Y���V�"�����i
�Q��i����R�>��R��Y�KQTku�Sc������c�3����*9�nڎ���y��WG}pZ��)I�gj���^����X��(`��;N�@Wv�(o��k$�nokSr�+��ݵ]y5�!�j��O���N0*�,v�ޘоY�ҮY�^V=�2f��Q��y��(���)x	��z����Y��ܝȦH��]D/2�;��5�\��Y�%s���6�����(��e}�4�M��38�g��
2]�}[,�j����T��a�s�&�l�8t�b�ܰ�f��<��=I� ��F0�Ff��0m�Cu�w;�Z���b `z��ڛ��������/dɹ���8y �yi�D���ь:�Ӌ �-E���oN�"'Fd�n��g;)Y|�&����`��P4�|����w�m�B�Z��[�y�!�&���q�O��+�TM�[]nn��)�^#ǅ�N���s�Ѕ\�m�ɫ��i�)
�SdY������3���Wx�M�ݍ;��B�Dk�7,U��`z�e���a�n���f�ە����w!z�Gi�do�q�]�!9a�Ҏ��&��m4;a��Hz��ڴ�3KTZ��2m���e�z���R��J������k���VJ����ډĸ1*'%�`����Ҷ���~t��v���u���\7U�F-��sႁᛢ�|��;�z�M�"أkF���c� ���>0�N
P�Vd���Oj-���.�
p�־Q�t62�[�:��v���c+3:s�,.��;k;P�2V�!T���L�o�nLڼ��ru阣u�F�5r���F3#u�6�L�f���kԗm����B��;M�����"2�_F7�ns��yޞWW�"a�	�\�5��Ve�Ǥ�ö�̅�kR�����	2��p�˳W��t�E�&��Q@ɴ���1�R�Y��H�>2Cl��$V�Y0��%���@T|qޣ���{�J����hq�w{�w�]��;������Z����V�:ka#�ÍJ=�&��K��V�	����s�ݦ���J�[��y����7u���B�ړ�|1��PT!�%F
��5j�:Uڮ��5�>R�T������@���i�Y�*Db6)�6�dTE厷���m@pN<{�O���2�X�C�����VC��\�Vi��oQ�K����=��d�z	�n�K{���	ٮ6rH�2���3�v���zU�ƔKJ4��Xku���lh�+gf�U'b6d'eu�N鎴_2�Kn�eھ#;.j�[��^h_Ga6�f�cg%/C4�vqH�W,8W��vK'5sy}����*��?
5#�(�ˇT�Հn��hK����h����G(�
2M�9��Q�q���Z��R�s1���]&�T�֝�zஃk,�V��3�s�
[u/���i��YZ��՛q^�a�U��7�ٴ9�θ�&Ah��^ean��r�/�*��P���,�r.����l�����Gt[�i�iL�W"l�\��=ف��M�{r0���ysG[�΅��K9Ft�iXF��$������t�;���"i��Kכ)�;и�}�`��g�Y�Z T��3�Dn�P�eɒ�4K�C<�*��Ù���ؕ:���^�m�Oz�6P�_���7�W7�����r�|�,J��t_U�+t̜i\Is�9p���ژ�JPZr��qf�;#[����\h���F�m⩣�}�;���lm��5��˺��,j-aM�ĸ�YEVn���\�� Ro5Pfo\�d�s�p%�e���e^ټ�A��W�(��F�n��v,j/�[���n)Z��A� �BلY,u�έ�x�����n�:.�u2�h���5_G�kzf.KK��c:-)���t�J����_W�[
������ֶM�f����@3M7�/QEl��;��ހ�����a�p�9gx�ZL:���Bd�t�kU����;mP��v�$SkjdR����k*���j�M̏�J��whVfM7v�9�����ka�_,�!P��{��Oq�5�ܺ+)3L%
|kH5�]:Xv��{lݪ��J�R��o�n�Q�G^<��!��a�S��oL�(��U�L�?��ik;S��}����E:���O�l�U��m�K!����lX�F˾�@|���V۽�E\�[b��Beb�(-��~:w����%'(����Q�ns�W6,�DuCˇV8�2QVH�&�)��OSÊ[�늲�dٖ�B��W��7��o�B�i����ŵh��ej�0�O�#�6�yY�<X�w
�`,�>�&"ͦ7U�M=�ȵt�<Px_-Jv���z���]eu��O��AZk���ĒfO�5ءR��Nr�l����K���PV����������\��'Y�L� ��^���ov;ζ��<V�c%=����)�[��L�-޹ݲ��;^��ʲl"�E�t��#hPaM�ՃTT����I4���+�^��`9T�ob9���8�9Knf�D�I��8���>.V��� 4�f����VJMX��f��V�ػe*X0��ܺ�x�^��w��X�B��3)��c��t��G��Ԯk-�թ}Gp�X�W�wuP�{'N�#�"���m�$Kh��7 ����;���w\��wi4w+Y���w��r��@�(�ևz����}��;�8ojuΏ#���G��Yn�hw�P��z*^�{[�k&鐪T�N}wJ^�����V��􃾶�(�ӕ�o�l��.!���&m(y[xhۡe�0�[ƭ7W���pGw���/o�����zWL4�4Y���a�]���7��t�*SGa˰�V�j \�a|e4�6�#&4
{؛�E�xm���j@�;�K���N�d6V�f*t}�����^�yGPR�º�v`�5n*���{�*�Z�D6���g�Y�Z��޽�����T]/}��^�w�[��B�r-��k����B��FUv��Z��K�� Pɲ�w��o�p��&��X���![1�+Md�rr���p���w�GM��P)3I�{�voHQ����tj+�:��چ���+͖��.���j$2���U-��R�`��bIPl'`aa)��~t7�g{q��C��ѕK/H��0�5&��/��U�6�Z�k ŋ�=�C%�@X��_Z#*
�x&�}���kY�R�9�
/j%:mv��4���2'@�����ٖ�Z3z�Z�4L��Ѷ�_of�4��70��@��ةcĕ`tÜ�$S�GwC{0�� ]bKt2|d��p�����U(f��k�>n�����ѫ-�S�a��oC��֡��4�Su��9#׊�ҰA8uM�⡋�ro7���ʧK1�}gv5����;��_v"�X��B簔ʙM9�t���bKl��Mó_i�v��n�Z�Ň�����;��km�]��ɣ���L�Z\�zm<�U�ThЩ���M��@U9A��+�<��5v�ԃ�P��\�ۏ4Q�A^���}z8�p��dXE�EĤ���M.��)�;F�ur:�����0W1����,��;`�re[�.IA��`[�q�A��3cg6E��|�BV�x<�&I�ݍIT�`Υ���`�7���h��S������(��(��j�����"���
�����)��b��� �d�"B�����	(�1����������b�")j*h**��(l�����
"��������b**b�hbIj�����(�Ē ��"���"�("�V��J�)#')����)*�Z"
����h���02*�**���"�"
������Z"l��"(��p�(����(���0�"��(��(��"�ʤ*	��J*jbJ�� ��"��J�hj&��(��b��")�
��*"�h����(�	�%�*���
���������))*�
�"���(i��*&��)
�*�("
*i�����
i�`�"Zb��hi����������{�f������~n![�!��!��[$�cT�S �7;9���2NK��`��*�`'�&Q�qs�������}�.;0�}ڥ_�U����J�טr���ASU�$��TY@ӳ9�tW����9���,�\Ltݥ�V%���Y�

�Ϗf�*]��2��:v�;}�g���@9S�l���]�&ohׅ@�6�J��j��T��L>�)^��E�ML��)���_����nfoӫy��%��i_2-V�#5�ҋ��/Z3��5Ւ�?8���뀫ԲȗN�ϥ�3�����1P���\*��{���y�L|�絷����U�a�[@1cb�_3#>V����s�}�#�.������@�v�_�n���8#�V��o����t�y�ݏ�7$R����1
v�UN>�{oQ�$�Os]��ޢ��M��> h�"p¹��j�����]�y�J���:/��z�Kj��щ��&b�*cr�D`�4���'Z\�����ׂ�CǗ��U0���M��^Y�Խ��>�,�94CO:� )��<j:I�-���12O8���Q�a��s��EN6w�k,�Q��$�5��i��z�|"�-^W��!���>���i��*��P�Z.U��nP:-9;��*�yГ2��饽q��s��%"�lޕ|�:�ovbq���ܭ�vQf�J[�U�	*��2Ӽ�K�Z���v~���-[��������-��ђ��NaU*J5��m�]hi�Z����˷�"���:����ڿ��,gCu�M��q<`��%L�D��
�il>�#��Rj���!d�WLp{��b]P���1ˤL\02a�w�ц��ӝ��	�<��Ĉ�`?y��Vˣ�])����*K4��^y+�c��OV��yd���|5��Ϲ�E8���#�_�/��x�U<u��t+�|/��$����*s>��ԦL�܁��b��J���C
��c�S��V-�}��z��X�X�5�.G'w�3\��3��>����PPy�¨*����T�.��,�}/��,K�N
��ZL\f��Ѱ����ac���M	�s�>.>����q+Foyz�N��`�rc��(�9qր���FY���xW�Ln�z8ߓ�G�G;�Zzr�j����~tQ�yD��=�	� ��I�F$Y#���z�d�r!�t۬{��t��؅�rɐ�q�Q�bw�5���}J΢F�Z�զ�0��k�^����eE͘�]u�[�j�ӭ��i�]���M<G:
Q�C3��,�%�۬��sl�	5i����oB�E9�����݅Vh�æ:p��xH��L��n\M8��L�^.�TGo>ZY���zڢy��w**��2*�=pٸ�K�1�z��8�Q��lH}��W�޸��OU{*Y�����$Ң`󠖎�zߒ���f�;yģ#.�r�CJ*hI�	���\�y�^NS+!ۿ����~��$�2��:᜵XT������W+�~�^�9���ͫ��5��l}p�:C1�v�W^��^e�Ի���""L�G�͛�X_�x	�[s#���|��%���p���c~ki���8z��p8t*��G��-����u�t�F��\�c��!?�I�&9���}¡k�r�8#r��)���f3O�ʛJ!k8t�+�'۪�ȗ��G5$��� n��_݈S�q_v����B��ة+�w�.[��}�KD4r�`-��9�(�W�R��`��q�aZ^,��u�[����_�MXܣ��p�[�m�p�,��KȄk �J�$8Pӟ�z�x4���F�Z%֗��)-$8��a�Έv�I�M��.#ޘ��S������i��zX�S���	$%L77����/��o�֬���"`W��~� r����)qV�q�Of�ʰʵ,�7vȀ���>6��ȳvm� �ګ�*94L���J ��f��o���]�d���W@�F�u������ַt	�ǱC��^�Ës�W�W�=*0\⥦��CkU��\rwr,&B������ʞ.�ۈ�`����(��R�2�X�+EE�ć�����ϓ�Z*�s,GB�A��3]�r�S6sy��w�������1�R#&�P�x�ji��0
뭾�Ñ��|29|�<̖f����]�/���]D���~TE��c�U�[���4��Qz+�9yU��`-:����I��z���U̲r�c;i�����Їf0Ts��D���~����t��-zP��紨�f��s�e��f����,�t�}�,R[1G���j��כ�-�ܪ��6��R�^���d��˗Eo�u^��� k����`t�6S:��pk ���8]uα��)���B �b,�R�].p]��*Wb@��C�a�Oh���GN&��Mޟ����6���\0���:���|��'Ū����(�R�9�nu�u=�Lc�͠�lHg%��Y1� �DpT9W�::	����d^�����Ť���lT�>�A�j��)��FF��{j�s�)O�51T��z{_G��yr��	)#�x��c�צ]��'	���Ɉ(M>�n�Djh�Ң�W<��k�:�W1�`:��V�\1\��Z�ˋ6�X)�W�.3}�S�����N����iD��� GU�de��f�L�(��>�c��j��6��?{��M��_z�vD*v��^�E|\��~�K���r���n|�Ot��'��u,�A�hJ�1�2øs���C�e�c%1?FB�Q0w��C,��kٛõ�n���P]��#�"ݯCN�R�|��.�?W�*d��X�ѐ��廪�n�
�F��T���2�Bq�YHu��G��t��ݾ�za!�:���q > Ec�������U����'��d���Q&��>)��1��J��
n����[ލ��mr�ӑ��T��l���]��/e`�
�M�����j߆2-
��|1�9W*�s��x"��`�<���q5�)w:�V�Wq*��J@ѽ(�ʃ9s3q|C��gg�$�y�ټ'd��J��Φ^���K�p�d��{!:���YƲ���Z!d�'9�Ol�����UhT*x�ݧ��/�8s�x��i����6w�ۦxX��h�D�-y�)*{o.geQxؕbn��fq0���P)��8�;=��7�9᩻r�KֺZr44�NHŨx�b�}'�s&U���fy�>�mE��ݜ����ҹ�=�n#�[f��:Omm�	+�(��$����Se�ę���I86M������}�v���^Fڠ���}p1�"���bTNA��b�i�����L��0�ﾚ��H�X����qexu,@��n�����1�Ue�.�(�|���.���;��=.|��n�u�Ȱ��4V��
몑�!Z��ݴ2�z�X/�&�y[�Ie�ȁ�ڷ�\H��l=  @t龴�s�'&��Z�{���Ӭ�oj��v��e��]ŵ'J��׮aU*J%�Ĝ"�7�F�t.���^`�@,�Y$ľ�шZ����lޖ7"��n���_�z��e�D��/b�7��u|=P]�Bt�<������1k�\��&��.�1l���U���P�9�r��\n�jW��%B��#�ʈ6D=�Q�WKc�޹���H���<j��xr��ޝ��}��B�y%ɨ��˒{��҅�B��w������#�;!r�(��k}a��;�+�	��jS&M��y�yv.8Œg��P��Ņ���X�Y�������� =����r��a7q�d�æ�N�'�TgyÓ1V��5Z��]�*�2�����mk>���CO�~�Y��?[n��r��⛋��.�ChN�}ִv+�f&wn"+�����Vd�_�n�H�C�s���۳�͍��a9�(�k��V;b����^\,���Ƴ�%<�g{��mA�

���2x?;ܹO�ņ���KF�>f��@V��%�h"6�.9��NG����4$[u���7!�R�"ܩ�p�7l}��r�^�A���@
��P������s��ڝ�M^&��Y�8���W�\1'��q�eWag��t�VI.�3(*���{���u�����Kg�'{= %7��U43���;�]*���`�=m�eP;�d�D/�5^�1����Zy�ks]�z'9�b�,"j9�2��}�=<�6�Q�of��L09zSM��bx6����gZU�ˌ#N��u�t��s��Ӕ��n����<z)IT��[�/|�)�{�������������]<�*��g[u�A���W�ͳ��w_ʢ���ɗ8�SB08G�*��$�d\t�$V�ľ���/�R�ki���8xg^'���s^Q
L��\w�(Xc�4�����;,А�6�
~����E�}�4�(e�Nރ��t"�A}O�u�s���`R�j�hd4�+
'DT��̾�Rfl.�Ԃ�l1v�CT�>�,�Xb9����t�WV�:ʵGz��RԵr��20|�=ҷ�{�0K�����7R���c��a�sx��DD"�(t͓2�s��p���~��-�<BW��jXy$����Qp�_J���b�z�Eޠ�YE�y�fZ��t��3�9v�m�qpA�2J�f�#pL Bg�+��&r\�����v>U[h�HE��6���%�!������Kc�6�eS!h�;��C�%iy.�ԍE����yf���Z�y��nxT����&ۘ�w�^�fI3�Q_�J7�ޅwKq����'�"s�&}U�h��V�Vt>C{�-7~��BP��?���"eb�7/���d~�y+���^@�ʎ�C���!{z��c*勎uLGQ�YkLc��p���!$6��/�L��@�YyJi˧|XW<ܮX��a4p����.wyr���]�y���I���|Ѹj�'n=����]},1_fO��,��s�� ʒ>��� 8xx�ObW!Us,��1���j���4!هy<CQ=n�S*�rs���S�F>nr����R4�d��u�t���V�m0�1d�ɔ��?:ͽ5�{������.��<�V8k�� �,���r�M�����X�R\;�Lun�۹����N���)Q�ז�-�R놽�]5ش��Ę����jPu}9�,_u�_>}�v'whIx��ui^D���#�7z�h��U���Ԯ�������Y�8FFҠ��sA(��*!`t�[r��S��T��7��.�淴���gK�wK�%�K�e>����S���z^�]f?��!v9	(�#U��p�n+t@c�� �+�1QQFA#&����Z�2�7��3T��_N����.��m�:鷽R6�U|�I=� �zJ`)�>Б[��TPN��7/ci��[W=ǔ�1�r�#�-�#/��O���ǩ�6�W�v�w�"�񴷦����2�g���Kz�vB�m�ρ͖�|\���D度d"JR��1U�WU����1N�>�U�,�D��\���a�9���]l �TYp�J�f����=[C�����e�kx���z�����0�<�g����5�D ������ʜK:�U61� �rP�����",	�"'�'j���ƎFR�Y^�w�Ժ1���9y���^"A�Kx�J�\�8��/�( �Br����ŏY�*��L`��F&?=Ҵ�>��j߭C��h3 ��Ƞ��$9��/iT��Euo��ndR+F��N�)򵜒�K����:fڳ�O7���M^��;�z2����q�)���t��@�n����.l��B�&K:6T�:���;|fX���>Q��qS<�΋�F��ٯ����~~*�_�ӻӑ��\��l���]��/fr�1�P<&P��b+zG43R��_zо���'���S���ҙ��:��jfI��^��ǣ8R��V��zO��9
M׎vg��J�=����X��N^u *"���2%Ӹb2\�=�Ս��=%9슢�8�V���)��E� f2�+��n��t_0<,`�\�(dB���C�l�e�vH��w���������B��ʝ7x���`��5&�� �wc끍�x.ڝ�fw�n��&0'�d��Y�^��ֻ4��]Jˋ���K��vc�ZCC7ܧ��̥P3��b��J��"�n����yc�LźT���h�l���'k��~f��(N��Yɡ��3�m��`q��X�4�[�Ie��!����\@S�-W�^Q،�W�g�e���*�:�� �Nq�e#�ɛeR��Ö8`���Ga�:V>�sB�t{69��u+��yY�<�2v ����L-$T�ju�9k�2%�_�ޖ7=�!#��`}��N#�e���a��N�#㓓�����!�{}�U�A��Ĝ���k�p|�op�R�xǣ*�[�QwIcf�ӭ0^��f]��7���9R�>����;u|G1��S0$k���L�Q��l\�r펏"��"^)Xɼ����a��B��6>N��wG������4f傩WKW��JhLY탥��D�]в����)-#v�WF�LHl�n��7K��F�W�Vj�E40oQ��7���JMN
�w^<�{��(3V���-]r�=��A,-�����k���7hI����vRVh �qNp�	M!u��E��Gnڟ&Ȃ�Y�)2�Y��)�0OL<|fnR��骻�T6�+s"�8�w4fu!�K�q�ԂB��Wt;FH9f#x���M��)�&�.X��P��r���@�lD�N�)V�#�w;z,%������Z}@w{r��;��"�щs��tr�y1�@��%b�Z�J�%��1���@���)]3H�黕��>=���=L*W�o9w4�[�-��+����B��;��R8\�#�=����14)��i�#t�S��}0+P2�O��@��f��|P�^�7mD��Ͳ.S۸�@��԰p������o�e��@�R���μ����ߐ����m�f��GO����p�3q�¶��t�)��X���N��:�5 ���F�2l���=ے�`Dp�e
(HIuv�B�`Hi%X�����G���l�VQ���)������Lu��V_nu<�}g5�6,2�$���aֆ��rM�p`�r�<�{�<Nd�#W���{wz��#:G53|^;tH�����*q�:��hv�Fպi{�y%��I�k{�/��"p.����9�m0+*���5ҥ,�E����%'Vr�u��7B��I%�oI	��9�*��2)�2�lR�ڔ�GDgN��a�����	�yB��9*�R���m��/�9}R=7z\���K��[�|,j
�Ws��Ki,�ڄ-��1�4��6�J�u��o��Zk� m¤����`^8�Kÿf$F!A3��A���=�#B�Wl7��.�S��:;8��{����8�_g��j`ѵ��mT^��]�)�YFAH^Ҽ�ps&����jr=�ֱ'D�t��9*�[Tb0=F�r��fv�����l�L����'+`@����i5��@��p�-��&e�έ"D�W^�;ץ�z֐o�+n�֊�O�d���(7�����-�����z���LP%�e.�
��$�gen��k���jB.M�a�Mՙڳ��p�@���Kp\��:1�ud��RX�;�k�hL�@Q�ʻ%p�$�j��U�Bl�z��f�Z�=�����`�tP�eK�g\]�kW.�}��mb�-M���(R�>8z�	sk�nmM�j�K�œ@ֽ4�K���@��h	��e�LwY������]'GUjL�ec���> 
�"��(�&@�)��j��i�`� � ���(�����"(�)hbj�����*�H�����)�)�((�����D����Z��B��� ���fY�h
���*�"�X�Jj�*���*����j����b�&����(H���(*�Z((��)b�h�i(j�� ������H���)J����(
�&%*�(""����������H�����$*���)��*"�J���
"(j���*B�����������J)������Zbih��*���h�)B��b�(
(Z(h)*����j��Zk�������8�w����Y��siɬ7v�b�ݽ����!�ELMW١�`��Tk�ۜr�q�(h>�bz�P��]6Mw#n�Z:�˝3�T����ܟF�����5	T~�"�#�j`��2y}�����5	Z�y��pz�Pxu�u˜���٠�������NK��#﹥��~� ��}�duei�K��ǝLϡ�}�}��NC�r]F�=�:��.f=����%;���Z�}���5R?}��#���	����&���޽�n~���{s���%S�r����ߵL�ӆ�Ū_�DC�b5���1.��9�GS칬y�s]C�2r\�2��h
�����W_`�N��=�pZ�%%��R�?G#S�용
L��Ѹ;�:�<Ϸ�ֿo���cX�}�K� }�"��",DX���~���gS�Ϲ���U'g9�èwHu����<�Q�r�����ɒd~�\�����x{���]F����7	}����u��]�}I��/M~5��N�ΣzT��律���">���#��T��4<��P��]~����Rt��{|��)�O~掤���+�kKEѨ5<9�|�2w~��惻������+�~��ɚ�ER)kY����C}y�}�����>��s�fA�K�9'fa��%�F��Z�������u~�Q���ؚ��2����w�d�\���t���!)���6�f֦�c�� }}(�!��*k'OnLu�9sל�u��G�1��1>�B>�5>���5&���5��%S�6�j�O �%����G�uY�ѩ�\�>Aߞ�����s����
A�������?A��\�u�}�;���+����p�}Z*�D}@}��1���|�ѯ؝ɪ���x��Pn��5<�S�<��ƴn���ut�O�u	T��;�p�C�����<�Q��|sz�>��$������1��UN�w5S�r~�hB>�DG:�C����uw��.�����?K�ф~����.I�y�����K��~�Z��gy�����jz����%>��Ñԝ[�R�����k�r���7��|���� ��DH�O�����5͎\�Q�z}�N��b�>�����*�K�����=�!/0�=����r]�y�7˻S��އ�7j]F�6kP�\�w�oOJ�o��l�5��訌�E��{�=�땯�V�i[��;���ԳuoM�;�v���a�i��,�o�e�l�8 �^���Y;��t�x��.��5k��]o;��C��a����sU�U���=�s#��Yՠ�k�����:��+9��Q(��7L�w���o{��#����x&O�p�������n����`������6�BP�~�s�sX��ީ�䚎C�j�����䚏c�a�BPy<�5ԟ�Ԇ�s_�2�|����~���/����m��$��{�%��|k�-����7�4n_mC����������R:��}�� ����#�}������|����>��"8E���}B[k��J������?��5	G3�2 �6~���:�Q��:5��>��$ۚ���<�����zw��������-�%��|���.@u��Z��r|�'��i�"/���D}m���Z؇sp�θ�c��u?�C�w�/�L�Cݫ��O#�J~�s�ܚ��P�PPr=�f�/�L��ϯ���.�Pv�Z}�.�����i��eξ�·�0G�,��l�v.�qˊ;�V�s}�� �.I�w���=�����s��~�Q��9�7A����N���L��_`ox����t��s0~�5�0�	A��}����5��~�n~�dЯ¾�5���������}@}¬}H��� �%9�6=_I��Ǜӿ�r9.�9���:�%�a��k���d�rMw�d:�>�q�uk�`�ް�]�}}j{����!�{�}�IW�w����8B$}}}讚���?C����i��ruy�݆F�)�G>�os���������dw�h���5�f&�;��#��;��ݸwt��5d��S���{�^��Ume���=�����
,Dx��u>K���9;�/�I����{=�K�~�֡�>����d��o��N�P���h�NGrj��������˿���K�C\�ߗ:��vN(ץL�҅��`b>�C�D�B"��b��J�BS�s}������=���%��7���9/�S�y�zJ����~����P�]��ͯq��>�>���O�1B(G�*/��۱tݾg���}>K���Q����.BW�?w��ܹ��w<�I��N��#p����oG�?A�J:w�!��A�;:�I��2�{'����#'����O�|�}�U��f��n�V�VZ�~�7/�\P�G�6����?^���=��A%���I �]��/pMSt�=A��N��-�X�\�zR�Q\،�wW\�>ѺW��fu�w!��G��|��.�EnP��J���TW�X��p�А_6�����*��H�����̐����FK�]`�<�E=ː�Z�9��)ܹ��u�reI����5��:��x&O�ru�����Ӭ|�����z�T>�G�"
D��2�\>���Q]�V�������5}��/p���7������nǜ採*�/Ѯßl{��Ky�^�s����l�S�ܝ~�p�k��u�!�~��AѬ9Zc�#�>j[�*�ף��}۶��1�>�cR�z����Ԛ���_��Z(7�l��.b��֞�ې�亍y�hJ|�.�a�0>��J��~�]`��=3�w.�|�:t*b���}�Z��y)]��o���H��_���|�/d�a��HP��������5����Z=�����n~��y.f.��[i�P����`jy.k�w�:���j=�5֟cP������=F�W]Q���_[Z�O
kg���vK���}�y=Ö��O3�!���tkp�OrQ������2�a�s����֟��2_�}�៹��{� >�3�7Ԕ��t}�#�Ԝ�(}�{�P�������a���\��UV�]v{�:�`�>��p5���9�����<��s�5'}�j��2��cB_`�f��pFOg_�u'Q�ynO�]��J���h���@�������#�j^AThZ��}��[7��?}��8��|����07�ϱ|��ΪB���թ:�^`�?�N�I������MF����J����G�j���i:������eF� ��~�xfs=]��x��t]R|��\��%Q�����>A�~�ZÒ��;�����_-\9�G�������Q�HP��`j�]F��:=��K�����u�S������}���`�d���x?+W�f���������xy�]�&O��MG�w͏��%=Fk�MG�{�=>ލ������>���`d5�u�9��Q���������G�nw.k2B��}WuF�_�u�X�lt<tOԿML��Y�߽����K���\������9����5'$ʼϴC�{���{���'�<��m�A��$f=��w<���|�zu'�d�<�P���
�ƬU���(�{Q���0�7oGc�kXb���p�j 5�6kX�ɑ�.54�}t;3h_M��@q-m+rZe>W����v��"�Q�ن�Z�u���H�-��#&5���N���H%�ݗ���b�R��C���O;P�\�u�a�1CPu��qo`ą���]s�9S�M����'��i�j�>[�k��%_bu�r7����_g�����~��%���z�����^�oݹR?��}����g�&G5���5<�I�5���c�$}�oP���~կ�kw#u�G�R�s���:���G�]�֡�����)�؝���5	];֏��0w������e�OS���>��K��~�s�rA�o5�ר�I Dgyܧc��������o�Q�C]F�ż�S치��nZ�BSܹ�m��SN�ʃ�2��������d���f�r#�Ju�ɸ��jO�_����9~�������/��u��M|c��G�[/�go�T��V��Ͻ�k�x�.���sa���3 :~� ��Z�xg�O �{� ��թ))�<����jO`�3U!C�~�GZ��w�	��va���G���U�l�fx_�ǿ5���z�����Dw:���5��͉���=w�Opu	{���sa�w~�P��Τ�29n[���N��%_��9���=���s<�q���F���Mgr�"
1�Y�=�^*���w�^��� B�v��p�w�s�z��>ړS�j<����'#Rw��w	T�����y�/�������c�i;��)�����0A����Gr�{���6�)Dt��k5���:�s}T�+%�O�C@y���Sܹ�ì��F�B���A�r]F�ǳ�z`W��y�wAf���:������n�V�j$��m��rcz�x�`�3|���W5�J�с7���
ӿ������֗G�!<����
�ٹS��Z���`i�5������;W�Gm��5�<I���:�d_�>��^�����q[�M��]�$�#<]U�D��$d&X�J��{��s�M&�.Z��6�[�L�Z���=��V>t�*y��<����?+�gF�ɚE�
SS��-�����ia�m��t�J�2r��JGK;|�WY�+�J�E�s�@�%�J��Ҝ���h�1�g������n�qC�^m�YؕE۰�����n�;"8�zph�_��1�s�7Z��a4�K�E3���7�N�;�毻r�����f�b��>V��RY|ph�6�T ���e�g9�����q�hpO!�fo�����c9���P��K��p�^c�X�YԆҩ�/N�^~�Eo�T�)����(z
���9݈d�z��m_�ޖ6��7K`\�̌RJֻ��އ���x�>>����<$�B�/���8�oW��@h�����/����;��b�#�R'�,2Ss�7n�h�f:��#Gd��[N��t�zջC����t�`��Ns����*6�*�M6�x0�b���T��"~8��my"�׎��cҢ�!θ�[�4���Wx"7�<Ğ����,��2_ɺ�;�b�<a�7H%n���E���iP����~Ȝ�/"��u]B����\�ɨy,N�'{f�ȉ~;�pZ�w��AWpգ]�c�
��ZL\Fl���\s��\���P9Y��I�^�%F��[�q���]��� �M��=����4�ڕ�e�r��j���ts���2�A�ƞ�~6�iіbϬ��!�yJԼ�ǌ��Q:[�*U�D<��d�*��ڸn�k_�=F�}�AH�$)w^MB��RCz��e_#9���UK�u��ٻ>�;f�\s�����O�A�0���3� ;q�1{q��f`���L�>r�BGt˄������iz�Ɨ�J��7W��1�Cݟg�yD�d��;V���L�V��:1@�^��D���of����uΊ��rLTQDz�	���#O��A����䑫��5��r^\�&l찬5�y����9�x�4w�{7'ڒL2�к��ֱ�=0�oTwj��12úuNf:��0������e��2���nV�88!���=gG�[�.Wr�a󈃏�)�@��K5�%�+��5�����:C2�geTv兛sw�=�Kp�g{�*�~uA�CĘ�|�H_�(H�ۨ�p��

Kc��k��������y��;&L�D'���L&�C>�2_r��v�VeX�����N��G�N�����%SŮ���Y^�jXr8I2'���u�b�\>pa��8;Z�}�NW�z'INl��`����eL��٥�q�=�JJ�guK�;���R�䴕dM����ѻ+l0�h�0%׆{ݟv�K���s�R��E���x ��w��j�[���xű��8zt��3�M=�cX�򝈆���}a	gE9c'N�1�q�}� z��t�Z�FuԢy��Is�.?�ﾩ���'�/M��x����+���S,oP�[�َG�<O���r�I��;���'�*��늜�����Lf��}*c���h����Zo�Έa�1��vd�Cs����	y��)wӯ����_�j��ϑ�E��u�t>CP�|����������D�5��r�T�'�F���\/�`�ﱠ_ڼLct��~؉s�g������-����is�'O�!^j�W*x8J����5����Q�%o�eE��+�Z�n�9��1���n�%|tH�.*�#����<��ڶ ��L�u�Fں�ڜ���/J�d4w��>yK>R�N����f0�[%٘���j��*��'"(�3���ߞ���^�]l7�+�������p뉖2�?mD�+:3�N�R4��P�W)�X9�3�k�n�%��]:M,��N5M�%��tÈF�G��+��(]EDm*�������
XxV����� ����;�%�Ò��֎�*ᮖ��@j?w��*>O[��>g�Q
�؅P���f�qW"�TP�r�^��p�d�Ee\-��*����ed�Ԫ;a_&r5�K�<)=N�}sk��9�������ɓ��x;�T�/IH����F���*�l���!�I�8'$� ���w3B��Y�^�_����}U�M�Y��[�����|��{7=77::�\�Tp�u����4O��t5ꗕ���5�'J���J����m��G������K���� =G��\z65͸��z����t�`�F3ֶ�o�[W=�n	��ݑ�i�P�f�WPv�@�R7��}�ƞ=$?�]|+�-#ơoWR��h�b��6�'VD�|���J������\e$�^-}�5��19Θ�C�m}u��-Qd�Ӫ�ȇ:�=^�sV����+蟺�D����l����b���H;����ka���o|b��y��J�~{��*`kQDE�)�����༨�ਬ�Z+ԅ4�`��U��d�{`�h����MMQQ���NX\+�����>&e�itqX���vZ~탗8�N���3��Ne+5�M=�ۨ�r�1�~Į�8��g. ���b�w��)9F;�.ӻ}���+%��= c�������e{�l�/�/M�ɵH�{h�dŏ��@���{���wo)�v��:U�f���ӯ,�fwwt(ӌ�&����K_q��O>���'*ԏ��	 >�9KJb�l*����N�	���w�4��GyB�q�~�h ���c�N�����L/��b������2��67+��u�G#|'����ﾈ�}���,P��`2C:LeD��'��r��x2r�3�z��
%Ӹb2\�<��GJ�r2)�jw�<18u��Dbʝ(@`�!�B�*��|��8�ι�"�J�	��1��>��,�����~����7��:]�<쟭O��:7�I��&�[*���#�����H�.vjhD$��ny��r�j�U��ț��;n�eܢN�9�2�ۼ�����.����9Dh����뻅�]=94C/�w��t��ț�]h���7<Ƈ�Ͳc�F簕�g[�@?��C���FϩLXbD�T��%��4CQo����V.�vӌ=ys�v��0�0-�	%�0�3ce#�ٛg�v�鯜���Z�#�ԝ<�^���wV�yy�:D>�T\*R'���I��ZHy���s�C���G�M7�o���v�Ṱ(s�࿽��� ��29$�|�B&{��\WLpz�š=�͕f�����6�\�a02ju�\<w_,�P?$_�Q�����oԫ
�ϞF��<
2��d���\{��ڦD�e�uw"�����x�0(���n�*	���-��ɑ�Y&xXj�f�lV�g #��D� �t=xN7�W)��'3΀�˕���@^�R�A�S�9�Uѭ�*8b�J1ނ�:qռ�|�ѐA����誔�cw�����Bw�����Pɦ�p/ :`E������QWs�zV:��pq����}��P����h�����Oo����)�&�7Ws���J��
��'�X2'�t�P��<�E�N��ŇQ=��{lX��N�����%=���ey�Y֨zT�A�ϧ��RpnN��z=�0XU�b����=�*��քf�y�E�-~>}H�zkf��]|<�WkH9(�hS�Tg��q�6i�9�j��%���Uc�Tڣ���:�ms�wmR�H�Q���n��K�Vo%5q���x�3�7\�4d[�����A�7��1�=��U]���v&c*�G8vn�i�%10��;�)�x�>~�u=�
����b4��X�U���%�M�'��ݴ��3�]��1��P��S̾�w�nxC�_{*YZQ������z{%@���B ����(��L̼���\t��s���NS+!ۿ��{"�3;0��'2�産8���$���!���,�_eo�W1Bj!s�>����[�}N����SN�J���+�Uo�u-9,�Ye��u>�q^�M�{kZ-�X͍�6��e1\��-
��x�ژzl��t�{E,7R����5+xnݫ
�qB��o�ٮ�+�E5F�!:�˵�_���WeV0>i̧���޼�@vwB�mނhV\5)������!�B��E����r�hچ��䬥Vk��j�Ԍ��g%H�4S�^�F�}�:�a�9v/���1c9���	�{�V�R�`\�rֲ,EK,M|h��}�&��]t�J�f]�P�GTu|J`;�Z��wb�֬����!�1��U�U�l��\���� �[�#m��P�O�ojT�ɥ�A(PP�}�X�t/���%���uȝ��݋2ӌ�I�<̵�����OF�ܡ�V�w'J=p��Ƨ�Ե�
���\�葸A�i.��:�YSy�kn��O�ode��e*vh���&�g3+lU�N�N�Dq\�[\Vc��r2�j��V���
QH����Ŋs��|k4M*�\G1���:��2�r�W��)3���iݽ�u�l�\�Yt8�����g!ʯ6d+��]�@�}m4�[�//2�jb�-�B�	���ub��v�r���X.��g*t��R�*`����3h0��ٛ����a},�(�ݚ��R��Z���%_>Ha6���W��{c��&6a!����yN�&�;�b����#A-�&w4 ��*�k���f'V��.�2�V�����P`[����k��uj0.�m<þO���o5�j�/��q�J�]t1�ܶ�B���Q��6^��W2�k%m���{���]�[�K����<�F��|.���N��gB�a=)��`��me����(sױ�6j�J���I���y�X�u����Qѥ(k�-���l�s�&j�l0{��$���+��KFc�r�#� վ�P��Z�7�h������ܹK.��;^�ڳ|��ǍG��f7���*Nr=�*A�ĺٛWX�o��u�qJ!s=�XChh���}��e�B�jY���ݸy�����u�@u,p_�눶����恙�;L-@	�p�ƞ���]w���f�WKz��5&���2���3�rei�q���[Ii�k�]	[�r��jLQQجXvv�4誻��iǉ�ҝ
��� ����9����m���dvfպ|bd+�{B�ԭ�Ԅ�0�
u�p��މ�GTr���](��Z<Y���c��0Ί4{�Xhe���oS�|y�x|)S^�
�����=�_�uȰ
�O���)m�I��}��84ʽ�$\0��[D]��vV��V�Cc�8K�g#�f�[8vV�5R�Mj��)�\�J�մ�7Z�Gfw+�Ȇ��[0Th�dc�jژ�=��M�y[H�e��T��t�Pu��"�Xg�^�w|��VP�u]��F��{�Pb��=v�6k����h�l��W2������*�U	H��J�h�)V���f�)B������&���F�d�""	��()JR��!JB��i��R���"J����(JH��X����"Z����� ��J�
��*���h(B��
*�%�""���"R��ii)(������$)*���*�������h�)�J
��j!( �� 
A���J)
�)��JB�����B���i�j��JB��
R�Z��R������������X�}�_�߇w��j��j��峣e����M �e�Щ�i�g�����@�V�-�����bۼ���J���ֻ����>��"-�a���MG@ҫB��g��
�T>$�W �<���Wq���t�t��
����5����X���a�Y���#
�Өq@�_G��@�hmO�u�G;vz�����ϯ�i"��]������Z�q���9:C���04�,�H�p�8ҡ���K��@]��F�E=�nǾ����^}�����x�:�Έl㝬�Z6 �$������M�ʋ����]��& #Q�=/���2����1��[�m�p�/��/>E���';�N{<��z��Gzi!��a�X+�SH�h����Zms�<������3��T��u��竽������?��Q.�����k�S�_g�'Zk�r�y/��8�l^���ڝ������C�L�$�6>Q�Ə6�ٮ�����0u׶wk,'c��;���jڹB�Sp��f�ʘ8|(����hS�<N0lO��듻ҹL��ck_[��q�c�Xx瑸͵l`!♿���7]D�����0Eq`ٮ���
��6G��) �2wBy�3Q�9?���\2��:*�����j�������K���/skA�1�b��4���9�V[ɬ�d(J-uӴ3�&�uU��x�Ù�z�t�M��V������aqX��&7/J����:�>g�ԩ�,+�ﾯ�v>���_�&?|Kzx�4�z�}�1�\<�U&Y9��v�W�q���e9if	[��[]ƚ����S(e|&~u;N΁*CR���6���S̰q�&z�m�dѪ�q�����ƝVz2�[�V��(xS��"�k� k����Q�f�edp�'*�nT!�DnGUN���7�)vT�v`�?&A�B����s����=�m����Y��7�UU؋a�z2	�1���_{B(��h�3ꃀ�P5����,*��rX�h8��(�1����vo������������SÐԖc^�D=ꑶ��P$�����{Y�U�م���ͭ�w�o �)�A���[V7�|����2�qD���N@���n��sHιZF�9�ʜ\C�A�rE�U�)�# !�j!oWȅN�1��-LX��M�Jq5��0PX�e��hΝ�������e����A�0�*���{����Ϯ[Y"�Q<�g}�ݻ漙�;���Fx�u���ϝ'Qq:�U=aF(^߈x�AX�ο:��u�a��-VZi ��֝�N�ɵwEҥ�.��~mi�Q|X�APwX�v�]�m�k�{�b(������/`N��fS�&��p�&k�3��O����d����r���d��P�	�-�v��\UڞX��w:�gn��ʄ�ˠ���B�={��n�e8����_}U�W��U�۵:F��]��2\2�֢��w�Pq;@��=j���<bn�^�e�>^�.�d�i�E4��W���X���r�_���O�,��姣���Ut�wm�]	j��`�*+&;J͎�ue��9�����g���}��zVL�Ð������ne�yB
��g�9��if0LOF�3+�+jO�zn�E����1�*:p�sԢ�S�MX��؞k���'.�>�Z�c%Ӹb�[��O_��	�ל�NA�����U3�Q��{PU�顕.`C�U�a�J�b�`@0��B0���L�Uc|���2+n��l�B��t�w:��ܩ��a�d�j~P���(�o���Z��/�j@�qu؈��\g�fמz�/fK��+>3Vi h�'�:�!�Wxĝ>���^��0�_�����GON���pً�үZ��&G��^S��=�)'!	2�t	��B��a��0��X�/�=<Ԗt\�Zڎb�D�Ⱥ�_>�u��L�\#���b���2)���#�3I�_t��89�E�=����QZ�t���t�n�m("s���MI�fT|&']`���%a�.�u�v�M������k������'�S�xo�-n���[��L��{����W�}}Q�p5���>����M}�@BI@H��f��G녵X�;u�Ӗ8`�K]�z�kck�a���EsN��gG�]0�8�e�@�uA���C�Tl�����3�*���V�v�t���z���޿��o������O�,�(�Fc��ചJy�n��P{C�����{K��3{��h�G[�p�i�C�Dņ02k��h�D����qHH��{�����C9{��o�@����W����U�m��� �#����≈�#vs"�U�������	E����z��r��o#{��ކ���2x�9�u@NU����cV��y�hon&f/Q�<Ꚙ~,�;GM8�X��{>�ɤWTvi��k��b{�qGg�O�����AWp�Z0���Pa��<�I�͔��a�Z�rc\����f���iZ��Ӡ�,}_x�0籬7��ݺ���su��{K��5�AhيV�i�� ��1h�:��u�ŵ43N}�?[��W҉ݸ3|Z���o���1BvS.�
�⥣3b~�|��K��?y���Me�2հ�[Q>�ã�������{�5)**��W�L���L��,B�����x+]{&��.#���FV�/�Wv���6��=ĥJ��U����/$�p���v�?W�}��U|K��?(�ϥK�@��y՚�vc�y#)L6M�X�{7�p��:�E�1#�����PN@�e��k�OuI�6���u��M�\�4n�
�a���/TE���^PVo�@v������{��w��+�GG���4���%���~J��|Ę�Z��t��0xm9L�7����).nB�pڻ9���80A��Ih�Ab����g"�(�p�b��.v��E�&���d<���ѫ��:���³Ʃ
���&?��'���}�Q,E��ӵvm��M��=��(d�,?��h�D>�����¥P�\�c��a	��ZLc��E�9���+E��J�.�k�5�
Z�✺�ܽ8�:C��s e:�%T�1���<�7�#���u.��-Ճp�^蟳�|��}I:H��gD6Yɰu�|6 �pj�ΌK��x�H��׹����J<�����F��e3cx�k�ɶ�8CC��q��n~^���%71������+�p�Ҩ�^��G��U�����7���_���8+�)��H{D]y ����0i�u!L�E���WY�Qb�4�
���(Eԧ+S��i���,�����C;uU�z�E^>~�AL��d�N�p�'���g\�G����E�֜U&I+qCgm�K�:�F������W��"��=;6~�������wd�l��&�Vj��u��:��(�����v`����N*zo6aB7��;&��{�}�F[��Պ�w�5+�2�// ��r����j�1�U���?:^M���f���6�w��z]gz��2�X��T�\-t��Q`�b�vЧXx�t��G�׸�y�*`�g��*o��*�n*f0F�Q�j��C�3p�|�j�'7�^��Ll'�&�\����<b+|��U�K(L���ʭ73̔r6f"{�y
�2ɑ�jj���LUOvK�s����{���}�Aq6o>�C(L��;NΌ�*H��j�1�y��T�\*\u��An.|T����oH�ahyG��j�1�Q��VҠ�φ���4*�F3&�����0�>4l��L�C���|f��.Ƹ��f��G��EG���qy�YU��t�k!��Bj1���݈��ތ��a����/m�?_���W\+�����~����n��1��'�9lT�́DMd=���*����C�!�{�#:!U|�I<1�D�#�w"�P�n23Wb:y�Δ������e�F�*�^�M�*�-73��,��"�4s�@��W�JRN�mC@�r�޳�����.�3 �p�Q=��=�o�{����%�2�[S���	:!�oVDُZM�&���ۏl�W����菢&{f�O{���I@Hل"�����cxⶮ*̳�n�1�r�#�۲2$
�1�e�^u�K6L� �jeTJ�&R������5z�vB�m��6Z;3Z 3 �Ț�:�S�z�W��]-��${�G���"{��W*�5�gG�����!���iBx���>�KyKvY�c%\3_C�1<0��A�C�W��X�6Z�nn������_A��S�c�����K�X��PDO����2�/*�#��߫ۋ�񃙆A��^���S��1ͪ�7���健�9V,<?	��OF��C��m[�k'F���k��Q�;ҊCh�lz�R��6���C�S����~چ��mն#e.�f��*rդ�mԳAq[?v|Vzه�:{zS7���L;1�:�T�;�8y�13I-oD���ή�by¬G�P4t2b��~8�T���ɼ��@T^���[����9�c��JQJwA�r��7�cʝ7���&���J�c`H��:��jssn�{y����v5'�}�m���MZV��t�%:;�p�L��Q�:��s/���9sz���݆}}lA�ڪ�}�t��[�\��okJѴ�ږ�7���e�{�Շ�!���u:�봻�0e�@�u`�Mԧ=�着���sD���OYո��!Ru�P�;�
���j�Fm���<���v�C�yj��5����o�y�R\]��wc��crE}jy��yLG9�a���n�eI�i89m���p��ӗ�.~�OLpTB���OU�,����!�����S�7Z:'i�y4�aCA^�s�L><	9Q2����q�H��zb��ϕ�9Ie��!��PQ|��N�l
�k���8��l*C2:����˧�M��H�kj��v��,p��y��y�M��e���ΧΎ-�����*�%���B©_t	wT�
��g��Z1|g����R9]�˝�|�xhq:��3zX�n��z�'O	g� #q@J��5��YeJ;��s�+^���9�����W� ГT��.�?1a����/�;�����n��ˣ2�Q�:E��,�3$d?z眳Kj�5�ju����4!B�Rf��pLL���f4����5@-><�Gu�v�Dv��J�i=��S:ԦL�M��{���]�!9K1�lS{Mm�b�m''��Q��#g���Q�x�6j��#��n�̀��H6�63���o����ۛ�������S�A�c��m��&�˯�t����8d���ɘ3	�p�z�\j�̹$�\C�uG%�菢#﫱Υx[a]�h��a&aL3�0������D��bƅ�m]Gk�(Uc�R��T��g$�a���vK:�-AA�

���F�*�N�>��N��S��������e���$ޏ*J8J�df�AY���4$_<��iD��A���>���s �S���U���k�Qː�@�u �qT1h�:��7\�4d^��Ż���+)��t'����ro#sZ��o��*&e�=�	� ��I䌊S��y;�p����R�ȧ�.[kM	�@���;u�c\��Pe�u�;�7�\�4l찬�~k����{�w\�'�m
Ni5aJ��U|���)�(S$���J����R�&9���L�0x^,�T�s8��s�{�����!<���߅:(��� �+�T�p:�^;S1�7
�(H�I�Q��vN	9p�w �x|��S�9���j���~�#�I�P��<M�Mw��H��o��/m�73��ő8�[�/�R����1����s\��_�����訪��F �Eڳ@�ҍ;�z���q�ul����A���S 8�;�*��k���-�oVff��)���Qr�����sk4�1K���j�gI�p!�����g*��
�27�Æ��H<\F�e:�;u���h�x'A�"^�*D�G�W�}U��*f���aI�����F��P���9u:!NS��%c�*RJd��ܡw�fȼ��ޤ� �c��ۭ�l�/v��io
��t�Ɩ���}��{� �۠16qfD�x_5S�oYVxAnd�F�Ԧl� �<"����F��e3cx����&Ṏ�	,��{@����d��sD�ۙ��9�v:�a���1q�+J�$=�n�w�n!-Ns��8�k���F�����Hja�g��G���}Q���t�۝����Z�yo��x39���B�ж��-'w"�	��S,	--wR�OhɅ�wOʳ�nf��9Z�N�,�\S�!�oZ,e\�|ꘋ��3=�yՃ�׍ �}m
��ܽ�(f�\�({Osc���ƞ�x�4�W]u�t�n3m[x�o������N��� C�]���2W����?��VP�	8�YU��g�(�1���S)�K�1��B�z�4�|����o{����WŊ�k�����.�_G���:3�/�jp��چ"b ��d�/-�}�L߅eۧ@V#P�B�u7�Rtܦ�bI" �v��)rц=PG��K%k*0�n#�t�7�{�oO���Y�:�DYr�ɹ�g�i�i�� �w�q�6��V�SP�qM�����:ģU|9n�W�M೔�����FR�[9���+0Z�.�Rw�,ȗ Q��X�M��`b�Q�n�E)jwL/]<�[��e���b�O-�i�	j��Lk:�f������{�e�̎�n�̌mn��+�S����q�<r�e�6�N��420l�b]��S�
�=���^�n�pR*�Ʀ��Mzom�ƕNo&V�`�X��9Wr&[�p�v���9Y��K��7X���h�U������)-���F�K��Z�,,��o�g��&���ܭ��\����xP�C;_}�T)]<���Z�U��O}��V��Ѩ;1mb��2<U�)�J��I};��M+�\ׯ)C`�ŢM
),���S���\p�+�1+�t���_gl6[�{����i�x-N�`@��V�X���E���p��Ӻb=���}��r���������!3I��A �D�PĽ��9Ld:B���P:u�mt�K"��m=���h�9{u�+"��G����HJ;�!Z��6��l�+Z- 3�O>U���^�<��c.fM�R��5��{4�`�'����wXt�]����AFf[�C�����=Ż�v�gE.7Ϧ�z�py����������!N,���/2=��@����ve��#���=�^�=k)��qN�$�T��1M�^��;z��XR��v4:��k�Q��똤�Vm6j�-��;�2��47��X��|�n� pHR����5�)�E�+ByJ����n�]qџ���Dߦ���7��P@��j�C-oc
�r�4���ҧ3�KI����Q/&V���n�1�.iu��aQ���^D�	V������J�J�뵚7`�e�):�,��0��nݣ��l�HS�}�.�N!۝w�:mH�YvV'����cn���
�a7x����{]+�TUn֘\��y��؀%wN��ax�^�6�@�C9
w�t�򉫡�݃�Ml�k䙎3����C�t�Q��_��'dtN�	��b�S�8[��V�z ��vlyۊ���U̻f�S���;����Ed\9b��n���~�ab��_7���x{z�'�;93��5tk��k�+�G���+�c�����`�{4u+G�B4RP�� ��w�� ��5�C�ҔN����~Ɋ\�@ș0Z]hBT$+��V~��s������eB�N��:�x������gN�	C�#V\}��qF;���=(
�,o>\1�6'Sod�7��o+���45'*��p+��އ���'n�w|,�V����	�t� mԶڼ5�$9�o:�OGr�cR�������,+Y�����
����(
V�iB���)����i�� �
"��)�F�JR���� �
���j�%Z�iZ�)�h��)A�E�h"h�(V��hh�(�(iD�(����H��JR��"�X�*�( ��ii)i �h��)��(�(���JF����)����J�Z� �J
J�)�(�]�˿�~��<�֒���h��G��Ks��a���^TV�����I9
�U�K��k�+�O��բ��'*��ꪮ��)��2^��-/��,R[P�k�F
�r�F�lQ+�6\�;����w9*�3��S�����u������3��5��0��Q�0h�3f^s�<�=플'{M�U�b^�����S�v!`��C�a�Oh��	��Ш�ۊ�T �2%8��I�x�%g[�M�N"��+]ĳb����SÐԖcm���鑊g�z8O�$�;�&�G	�@��`Hs}�"�Mҕ�qW�g�ڙ�;N7$GFʰ߯^]yJwL	�~[=}!�{�}�B��9�����5	��oW�N�1��U깇7����x����[*�!�ۨ���T̊�S%)��S�$\�}4'���ar�&.HpҌ��s�#�cv��E��J��k�\��qq:�	T��S���V�J숾9�OryS�˰���pV�Y[=G�IS%�r�� E��A1��\@�f��W3�dj�����x�5:���v��2�*��屐ګ�xX
�健�#�b��HU����b��䄠=�.�]4bW
�Ou1��N<&	dM�FE�����F�:�f�y�{��hm_V�.�]c��7]�7�,}�j󻩕����v���3*�š�ri���HZSt�L6#���±A��w�g=�MR�]�����ٗ��">�*z���X�P>�|rl9S�g���S/M�V� ��U�*w�G��U��L|{ޔ�����f���TFׄ����b��:el=��^_p�(hiG] �V['��}�d���~�v�j<���Ƃ��Щ~�8���ON^u ��g�='����껌%R�b3�s��'V7�����֛�4c�������<0z*il���-�ME��p@V��d5i���O�UM?$6n+?r�n�������F�!O�'�cr��C���q�_u� �@�v>�ܑQjy��yLG[���>����X����k8�w��0:=�=�OD�����82!j�_=wp�����a��lźT��A������=��=�qp�5�����+�aṆ:S��X�5��o�5%�Ķ���KO۵������Eӄ���G/@W�p�G�%� Ҙ]=�cF�ܶ��n�����v%�oٔC�7�[Q������h�Rt��%���sB��#��J H�����$3�{���||�w�fZ�:�.�Q��c�]�LF�X7K���n��ǫ�$/���\t.��Y�&��Y����g,���廉��')��SN2��&��^�c:+.���9 Ev/� �H[eQ��n�c��������n��0.�}��.S���(n�����v�dc�l��suÆJj�b����wp��O��#� w0��z��5ج�5yb��=�^��a��f�U��E$ա�]"b���Knp�x�&��f:��d�<£+7hA��:2��N�5�F��<Z;|����&3yT2ju��r�� �h�n�Q0�ͯ�VO8�zg�N.�_Ձ��T��n�]�����D��)�&ma���rz	�[�;ʑz�UJ��S ��!��]eU��������^�W5Q�mNA�ڿ8����Nj�#��B�@=^���ߧ�h�=��qB]0�a����1Us��mY�;ۇ���kn!��6����{�|+��|#9f������n�~����oT�\�3�\1��J�z���| ��U\B2Σ9�3Mӑ�?[��W(��|��agp�1���w�w�FE��Z��^�̠��;�r:��d�"��5:#h���R6��c ����ѕ8�2+� mU�`;���s��q�1�����S̾ط1Umb�+ψݔ�՘�6�����AI����oD���٭N<���rО�N��]���#Ql��m��k���Mt�H�V�{w�;��T�;U��ؒw�y}�s30*��*a���C�ҳ�/��6��@#�[��-���淹��;z�TQ?UUWՎ ��96��V��11{7'�nI1$�PN��[�U �oݾu�7��˥�^��(���m&���yҙX���"t����	iLB<���'k�|u���W<9!Ínj�=z��E	qձ���:C3�s��m\>�3��B�p�,�|W �<�U��s��[y$�IU�t���@��4�>������U�ي*�B�}]��P~7���nN;�[ϲ88��D�����T-}qW�q���>:���V9�1̡6)cz��������}�fx 4À���h66W�~�+�~ߒt��s:!��M�wʺ0e�0J�Mf%�Vk�p��H��k�&�#�`���tn»��l�[���bմBÉs�Q��O�����w��=\��A�QJ���x�^1|f���v��!���m`"*[�ڷjh�q��1_$��7	�F�S��K�a�g��"�_Tby�@�_F=�.�.[���s6�}w��T�L�2Ӗ������A��Y=C&J�Svϋ�M�`@��C�ZcY7jg��
� V��E*q���(^l����G6����x{�����Q�2��d�ۑ��;�e�5��WuԄ]ƥEρJ=J�m�ح*�:��@RA���蜇�n�;�l����]w�;��l���K�3��}_W�x����p��?{���7��>Ϸ��2�X��T�\bt��Q`�f$Lk��3�P=���Vwt���ӄ@'�;^�kұ�p7N�[p�����@.&U7_4Z��ƪo�]���;��D70E���O�YuG�[���4��x�V�T�{��������e32�bU��j�=}M����B�g�\�;ʩ�`u�	}R��:0�cܰ��a��}Ҟ,ׄD�n_mu׾o$���3��,RV�8��-W��r��D���Q+�76�d�zN��`�/W���Kxm�ᮾ�HE�7)��u���7�*eJ4 �?&g�zp��`���^���sq]T�N��T��,�7z[�#��]���m5�X�a������������ջN����N��0ه;-�ˮ�Y�{?o�U<-�b�{D=7z�i��t��{76��{��}�"�+�$܉��(�Z��=�[�;�'�p��+��TuD�R/��"�Ͳ2�:k�|�"�T�!���
�s�:���xVU\�b'��?%����Ͻ�)\�w�qE�Tn��!�:P���Z�M�z2F��zFM�T�G`=.��n˙��+3��G�[E�Ty����nJweA$&��Ȉ�����=9��1G�f�ܻ�oKu�q��YE��tu5�Nӛ&�ִ���>���'�_UP�Ay<��ӝ��1�:Z8�cT6�'nS2'�~�CQ�Fz&-�u����j��FwpUm��{E=�>��.��rՖs�Fx���R�|�8���z�����I�z8��j�h��])�b�u �+!���?W�*d�e��Q`J�*'}^���\{W8�*{����TW��n��ewٷF�t�}5E�`)9`ih\�eVa�k9�W*g:�nE�}lp�>��fߴ����z�`�4#TBN�N}��\�t�5l)�۵�Ӹ���{�J��J�^��B=qU[?v|Vzه�&���qy|"L�_]o�|na7�I�IQ�i���v�j<�dZ,�FTץd�wS�}Rr�d`�!O�mȫnmV�n�n���}.��Y�u9�������gN���Qa	���ĸ�P�'��ݸ��MC����1���
ӿ��Ω������Gm�'F���ޣ�Ϭ�Z�[�6�Z���~w��"Z�ߧU�n���-nu|򘎷U��ț���ȩ��.l�߲3���]����FhB��]s���G��Oz�&��������`�b�%��� h�a�v���q�(q��p��m��S5�l�����ͨ8�R��54��X��+y�B�,�</
�HB�s)9�˳߾�w�sr�{�-~�`}'2�u�x3婡�]�<�=^��a��lݲg:�Q=W��ݚ��![�,&���$�K�T=uӍ�j`3P�%�e>5]@���L�fZ��k�}p��S���G@��
<���H�qj���ې����Mb��+�d��k]�u�:V>��0�*%� wTAtA������7͙q��!�{9vkĎ���gݾ�|2%�_�ޖ7"��^����Y�~�b��b��Y������iib1�q���{4�'��[�}�|;a�pݳ@U������`p�gnH;b7���5�����:|���y7���M;�}������m�+��m����r�X����f�#��j?w�އ6�>��6�����6 �v=�)=�'��徽�߶�6w��Qy=Ԥx�EӼ�4����׮�wjU��2�3�]�U�Af��]2��ʣ��kt�;��3;RZz�AH�K��__�j�4e�����K�2�Z�w������Qo��'��Q�8�v�wVmٚ���+BWh�,+,�Lx}�.�2���i��%�G��7��u��ǹ�3�:8a�蹦���s�ᣘRv%z"j3cZğJ&Gy.u{V��r��18�����F��<�B��8���8��0���l�#��Nz��{�����~|յY�{1n�ʎ\j8\�{�I�׼��c���@o�&�+�)���(�I�:�q/�s[�&z\7D�t��<�B�ˈ[g�"�<��Aި�tvT5�j�6*:?yOdҳs�^�ݵ�����Fr�k�Z8�v�?eXP!��#(C���C�]�\���ʬ�|��P��i����ֆL�W>�1�z��v���`U�WZ�j1j�MDo'��Yp�=m<�6�@����jRy׍�aNb��K��.#N>�{E�Ξ�|�<���}z�{��S$��[�z�6Ev8���N�hPԖB��Z�k�/��}��h���[�K�!d�J���%�#W��-���2Ψ��1&��s[��I�;��:Փ�N_�L5�r�7Yu����
�ov�U%�D�����M�]W\:hU�4#YƔ�`�ƕ�����j��Z {{KQ���/=��-z]���[.�\ba�諍�&a��d�4��X���&�j�{`>j���@�|Q�~��*��֧���jJ��`�.3y%+�<��8�w=+���@Ir����<Sb��vf�T���A\�;�n���c���?��}B/a�64xl�=C{q's5r�r\F���4�`�ɸ�pD����CdZڀ�t������'�x���"�;�#Q��{�ᚄ����#]�1�|u�qiM���+��QfOU�F�q��|���G}��}��}�����ny�O1��vySj�[���˅�$^��_M���`��N�k�x�C|ҭJ�3��(z�I��Z��)��S��}�fW���=���;�mʏ�<�v���~���H�Gs��c^{S�6Q������mZ{�/����}]���/s��>�'7��O!QN4+�|ؿ��{*��W״s)�f���6go]Vp���<��-Sܡ����K�cYm���Y����\���{�ly��yd��55p�6��%m��2Y50����@�9$�>����)��E�X�E�V����&���q�����L���R��v�Y{��3٬�م�uq�6�jX�έCP�s�}��;v�uqN�X�QL�I�QP��P�*�����V�̟��>�UD���[�ǡ��i���x����c$nIx�����9�pC�S��U%�Ξ�|�<�h5��=��Ĩ���MV�����y��̧�w(�rz��jI��3�W�����hK�T����Eu��Q@.ﻦ �~)h��̀��(�oz]R��k�s�=��I�֘�gi�2�]_	J�>�P��#s�yO+����f�sG�=�sJ!���3���xueT0g���~�U�#^M7�b4��,��.&���;���4�N��a�n5�7	���,�b�B�7P�U�=[�rR-�]AX����[W�is�ڙ�8f�MƺjR�g	�ԧyFgr	7���,�\?Z�ϭ�<�/�����[��s�+��0C�ia�6�5kѧ�Z�N&��j��{��s}Ʊ�kyOJ��U5F�EU��]�t?T�����I�;����x5��M��7�kEZ�=Sf�v�Q:{ɢyѴƍ��z��g)|�M�����|�>W�h�ޚY�/T.��i�S�ɹ���MK��=��ܔk��wi�loU�-��)�8���0>5l]4+D���5�y�:7�f�^#/^
�Sy�W(kb���A�1ˬ�+J�cF�pQ�1�es/%w���p��Zҭ��]��Wm�D�;W����k�PR�J�HG4k)�e���.R��L�Wp��S�k��Jۀ��$�F������m��Oz��*t�"���8Mh��U����2�5�A��v��|l���������vH�V�u�(I�S���>a�|3|9a��(�B���%>��u ����I�w�XVC�9�T��Q*���ʔ�HJ5r�]��e����O˩K�U��,�Y54��*�s0Ӕ���1�k[�u������dT�b�#3��G"h�@q�сVj�,C.�(��
Fr�}iҭ]R�=��:��E/t)�i.��z�[][}�E�aӮ��rb�ӥږAv�(E�y���n���֏p�����am_#W�t���Z��gu&%�/��8^�VWN��N8�v.���G�#�;V�ZJB`<c��E������4=7ҺTq����@�X;O0��vXуz�x���v�%�N�Աe�l��f�y!K-F$L��!�{sz���[�
�s2a��L��ܮ�|c��{u� V�5�yŊwÛ>z��n7�;��X�.��M.��mWe�r�}��z�Y���%�X�P��W0�q���)�*\��E���u-h�{ v���'P͕�.�jۮZ5�ݦ�L+�ŵ��B�Z�,�����F�L�0.	�KL籷/��8���M�;��qO�L��h���B�喲�p��<��r�I�:��34w.H�p��TƦ=����6&	W|����-�	0��9��ZPvUʚj���yׅ��iS'_'���k�Z0��i�me�(�T����]�G�Y��� pZ�FK�5r�Zg,���'#�@k�U�|E^�#a��n��j��[��`��P��Y�a�T�����U�n(�^��)ST�՛��mJՅ�a������Um�#O1�\Gj�]�	z�}�pS���}��˼�C4V:Ӗ�I���B�':NP�Ψ*�C*ewD��|�)t�Q�e쩤��vQ�5X�hm���`��˜�����JY ;�'R@���zV�'V���Hؓ�N��2��6���k>X(w3����x"���ڲ�\��h�ō�@�>Z�V5M^:6��Z�3�Z�b�l���C;�ȪDNv�GGY���e(,_\�z��IG�]b������Qn���� ?-��_��N�A�@�v�W��W;�ӇZR�wgz_tܻε�Vy����h((����"JJ�*�%�(����
T�Z��((�� )(����(
��JB!J)iiX��V%��$
 �)����
B�X��@�ZP(B�F�bAhD����B�
@i
R��i �A) ���D�A�)���D)~b$�P�/����o��Եem��>�ON�fX��=*e���u��u�w ��ӕa!]��8����v�n��>�N�t]����gi;�q�>�����Ag���|;������V
�2����=K�V_F��\�|�NZNʔ�ȗ����>#]9}Ƅ��k��]��/qwv�W>=GOOT	�}q_.eN��ު���5gڴt�j+S��g�B�w���C����w��Fӄ��Wk��I�u�xCF��o!�Ca��r[]��Ge�s��N�'T�U+�-���7��gU��!�"�)<�������T�4u:�֮�c�<���S�T���q%\�
�c��n�n�X�,w���������5m��$i�J��)⃡m��n��lj�j�MB�ؖ5��ί����*�Aw���d-���W�V�H���-� n>�/�k���׹�}��x���Y@){��2���j�εu�|����f��\��P���M+�_q��o \��y�7ps*�l�m�@Պ;�u����w���eJ:Dc:��bBZ�Xv��ɉ��E.�g�&c����{���r���]a��W~�z��v�%�3VR���k�86k��m��m�ƪ6�'rm��{�R��aK��]���a�եKvV���vjE�^���&����'��P��g�m\w'_>Cj9s5	�/��̜k)	2�u�ʨW���S&~�6`�}C��*{rNs���	0N��7�,��x�����l��k�F�^�v@��~]�6o��9���{� q��w�W�g)�
�M&������ڄ�]�����k�1L�ܦUJ�o�SO?��<�)����w�Oc���N9���z�˙�f�����k|����to����ؽEn�w��;-�)���|���f�m�K��'� �'}�&7�<R�WKo(j7'aE�Lv�Q?v$ͪ��ļ{��`��v��9�<�l�{fj�Ļ�D���f�x���X�
�6$s��n^1%ʺ�&���!]���O�vmþ����� 4s�
ŞB-K�o�,�/��8��ʪa�+灼����I�����=QHG��=; ^R�K������O[��@��WK[�,��~K�)]��9܆������)l˺9u��f�������aU�NJ�ܺ9WW�ɮ���qrE�:���JӶ�Jޖ������r�R�1v�����V㣊K�=}�݂�u�.Ĝ��}ۡ��|p�m�e����OE5��Ls�^]m�Y��U�}#���m�	����U2{��z?;��CXm��b/h�X!ol�f.
����p`%�7�������s�=k���۹Eh�i������^ǌe!s�eU���Y�Q���s1;�I4�d��:��U�t��]�fW+q�pT4�)�(�%*�h%>��yv�}�5n�vE���}ӎ�g��^)�6j|�0��n%R&c���uYZ祪�}'Mh��A��G�J���=P�Q�I0jq��,��tD��lZ�)�;��^��'	ڟ���~���oCKy:5i�5�n�5�Q�Ȝs��j��ř�� �n�f:�Ve}<��F�ڈ��w�����=ol�&����r)�-�꘶L���{��o����9�_9�Ź�\O���6�<��e��7Co�����: x<�$moV�Q�ߦ��-_;�X]�4���5#VT;:8�p��%���8ᙥ���؂鮣Ŋ
�D�^Jp�7�����ǯl�Ԉ�Cq��۝I�Lt��A-��IP�j7��M��&\��y"��@e?��~��ʿ�X�����V����6�������7
e&2"^�Mf�^ͻ9\�eAW0��;N�7��e!ۚ騪�N 7P1����<g��--���Z8�~dM0�'~[.jC�M����6�8\ut5it� cb���O��>��v��1Ӹk]��	&����$���yb#�,c̐���֭�=�㇩��2�xw�m�w[����`9*|���+�ܽ�r�[A�LHU�,ʺ���{�9���n�=������P�>�=fԒ,��z�ï��[K���f��s��X��v��r��"����R�CSX\��aF�v����q��3���V��Y�
m����0�]_	J�hܒ�4E�\!���.�O%�>՗�.{�k�{�j�|��+g"b#1Q܏��D�W�iP�߉d��Vk�&�MwM��#a��J�������Ń�'�Jߙ+P�p�̱/���>�|��=�+l���� ����N�KG��\Nmv��Y��&whG�j�-�7��8�y\�eL�F2���]��O�&3�6u�<r�z��#�}or�.����]ɽ��'�jL;ƻ�n=|���!�8��w�gӖ��p�Ur� ���+�+s.'9�\Fjڅ��ک���;Eڭ�|��r���*�7Y�Y_��h.~׼�n)��簛���\h5�>����:���B5�q<�ޱ�]P3DM�<�d���=EZ9�w��Դ� �T�[���1�jrT��&�j����������{#K��C1�te��M�����ݭ�F��n�c����W�ݔ�˞�=}�����79Bv_�L_.eO6��Ofo�P�/Lq_��K�qK�-�]�~r��u��P�@�J1�KZ��>=jGuͬ�-:۫�q��r���m���R�u;>*'\'_7.����L�[%��+�wH���1���=��(w 7>*ʧe'��6�l�5�� ̹ӕ/AS`A⋽V�Ò�L���S�i-�����,.��f�Uf�ؙ�˖5����7��a��S�c
+3p{�w#��CS��ɓ�;G�<4�
��f�|�a�$-4�O�y��B�$��\�ˮ��n���X�v�o;9d-٬Z�8����f/w����C����-��(t�Ϥ�0;�ϔ��:�V���)�^�﫡�T>x}�}�/I��2;��?.�A�_T�N����VpX���:���b�If#�P��[���3����e��FoKaj���&�m�w��9�`��k���r!KxbO���8v�^���*��7�B}�>��ޗ�{��R3V?C��/a�:����?�xKĘ������fI{��\��k*9k>�<j��]������B���.E�5�S�7�;�M���q�Ѻ�xD�!���j�'�8��F�$��z(Q'��F�;6��[]=^��7���|�Ϸ���f��h�֋�abp�ܹ�ʞZ75:ɦ��/o�N9���	��3�&��JVwT㱽��l�A`��f3}����/9D�[N��2�o�jo$Dښ
c^K���}����D<�,���Y�t]EE]���i�1�ͱ��UK�@���o9l_lI#J-��l,�HHO���n=��4 3��.����������b�Ik�؏"D<��;���y}ܩJt3]�G�M�9C�s�זgV�޷��:��Ft��C�9�M��y��n��\_[ꏧ���a�.�3��t�i�}/�O��O%�����Z8�_��	�V?V/qJ򸁮��%�r�<ںR��W!���4�"�}n�6���휔��Q������l�Wv���\��4�u�[w��}:O�l�v���=Rk/����K���+��b����3K�ۇ��zsi��ڨ�C�C�ʮ�N\t��M-�W�V���9���m�Ҹ[E�:{5�9O.ֹ��r�n���r��qC3э�^_�w����!-y��:���_w|�>��%hֻl
��Tt�-+����D)�)h���g�gTB��}?)dOdn�;�o�9�d3�y�P��_
}'�fGq�\�=�+}ܻD�LmB\�}����q*�3�l�x�Պ�K�`��n{��`��J���o#؈<�T�s-�Ck�9��z�tr���$��E��:��Gk�C�,���)���K*Q-�a]�n7��ۛ�*`K�T;j����f���l���>b��k;mT�	�h��V�.�%����G\�X�uBn�3���*lr&Y��Н�rQ����W0��5	&}	��
�\���nC�g0TdZn9u����e�8���jڈ]V���_Zp�&��5�a'�3���a�74�-����Ч�khf:��z/'�~GQ�o�����������o@x���Rc��b�^�;*�좽3�9�_s�:���?BB�Lx�g�������K�jNlz�c���y���#g2Oxu�m%ZԔ���x�9��y;�\�{�+������:�m�ʎc0*�w�U5t��7�"���nȼz��bz��cc��C���U۶��/l��X�\��Tos9�J��(��CW�ұ��������<����tgT˩\ ��O����"���A�Q;<]��eR�J9�x���
]�MUdN@�j5=����Kj��O�A�D줱]����%?yVnTY~���y:�R�'�F�K(
���ܽ�nNӮφ��D���ʈ�d^�.ׄ�x�4U�K���p��<���dRq�T� Y�G��XɬT�Os�^�n��՜�u
fkL&�4󯕒8k0^���VWe��hGǻ��8�ӗb]����Bc�n�wf�2��8�&c�[�J����3$5f�U?��Q�����$ڈ�rTw�`]�+��Uk���*\|q�b�g|�Ψ����eAs)��X�"��ORt|���t�5������{�&��oZ��6�T9f~D.�����;�wxL��Z���R�=�E�{�Z�C/��gW㔫���\�`��1�a���=��)W����M����� ��5	&�n5�4��;(��j)�-8W}
臬l��Q\���9�j��[_B��U/}'C��ïϠ9��������'�������U�G��g=�s��NuHE����Lb�4�/5���m���*�흦�٬�:E���b���k�+�gbn$+.�m���p�:��N��Ĝk���V^O;7�]��0�ycq"��D_<r�d����)���ӿ�=�[>};�=�V���}{{%|荎��L���Q�ӬN�}��('|����d�,tn�H9[elX)��AzMeu,������d�@쮵��a���^��b�@xK�m�P�!�g^�-U�]�����U�zOVۋ��8Dμܗ{	}.�aw�R�Ӄ�Ź}��olk"�wl疟��_zg�C��[�5Z��ߪ�^���-�ZMp!�{����&�I���Z!*����(�,�c�c���҉I���'-x3qr�q:�\َ�9QH���~�yWӲ�}:�*Z�+�\03�0a�0��s���q�s��}n�ۈ5�B�O 6`�?ʾ����
av��	\��qm`B�S�����|��j-�ۃIP�����(J*��m�<*iyL�)=�Ǿ����c�O���˄����:���(��эX[I�@{Upf��^�-�y��Ш�̈G9k���׸�h�xέ���f�M�̳�t�5KJJ�9-����r�Kxm$ҿ�|a����u`�s�.VV���Q֌��P=����'Jt�u'y�pԹLIY}o+����+�ȿ�R
�7����H�C`'�:��7�)�v^�OX�*ȝH��f	W����b�����{d)N�<��=���bg���7J.@��%�#[���]u�0�75��]�yj34�ې��r���t�¸S+Sް �\KXn��h1��$Z٫sn��f�L:å� N�`f����(P��a�[%5�<��tY����	��6��C�
9�TOE�ưW*{�1�8 +s��*��gs9���FGʻu�x2��x�)ܳFq�d$:lT-}�.���+�]
��\^t51��X��t�C�;�����o� *�b���37�P���{	��N���}5��%�����4��[�� a+d�@��3�J�hEfG������]ԇl�lɝ�7Z��ū2*W+cPG����O�f[�B|�b�~ܜ����ˡu\��W�R�nq=Ak����ϩ�"�� �87$�P��ʴ7s�x#�¥>V7t曄#!ܧ���ԅ;!�˥Շ~+c�O�ӣ���ٔV��\�w9����R�kz�-�� ��/N�Gx�k��RL�Qf*�}R��C��
���WeNL�$I��LT�IU�s���J=w��>nخ��%�i*U�;�WG��:�gd8�$��j�C�m��7$�x��q��-�N��~�\��y?�,�-&rL�A�sS�p�(�ZL�X�6g5YQ���܈]J�JE�mn�*ͥ+pjW�p�ɽB��X�5���3v��Y��#�ʑ-�鵓����LxU�j��o�c	�9i&����`Cn�)���d찞�R-yӭv�;<��
�B���%7q�x��V�K�D���G��%2m�N$��S.����{��u��n�l*��ړc�n;���:�.ޥz�{W�1�5��h�f��ʑ'A8�jޗX�vY��UbgP`Qގ@�
��wY�2p�� �"8`0b���s����fR��Ҧ$ۗxt^���(�\�uN�{�.Y\�ƦQ�OWtB۸B���@Wq��˭-������N�RX�� 6�v�]<E+�(������jeggv9�8�����;)>]n��C%���E���_q�N]}7pc��u�
lFEs�꣡�Z7@>�l�2ve�0T� 0jҶ	C�zL�M����&�ƅ3/T��ۻ<�-���p���yLo+ε�m����,g�=�T��0u��{��i��ݭ%�Wتǣ�%0���q���4F�DtA�Y1P;.۳� �\��7��{�u(���ήm5��hk��A�6qe#ocqN��/��]���dY�
W�ۄ�]Z����-�
I��N�lJ��q��Oq4�D�����$�{\�u��Y��0(�l��s�c��.���T[�&�$&R�NQ�Фַ�z��W�{*f}g�	Q���$n����]`�ɔ��+w_i�|�n�B"�'����ʱVۘ��۽�݀p9Q���v7)P�vS4j�X�R(y �*P �%(%4�R�%*�H Х B	B�P�Ҁ�
R4���R �@�� ��@�+�"�ޘ:���kcw��}��J
�� �{�D�ǽEX�iߊ�RRhY�.ʸ�{k%]��)�bn�W��k2Lf�Nu�?R~�mOC���`�ɸց��dO!�}��F��%SuL�7��-]�V7W���]V�����N���s���k�g����c�;���p1mDOfz3c5:��w�^�t��y���ʯ+7R>[�kғ;�ޯL,Wm��6��(�nU�ڧ:�5���o��E�ۛ� ���{y����{˔��u��9�N�(��#�qU�����k�˲Й��nR�Nb�K7����Z8�~�BnXL��J�q������WE��N>Vj)�Ш���E4���f۾���H���v<ؒ�5J�6�/R�T\]t�z�_�[�7����>�[�G�����M�f͵��B�Og}�7�D���/���Z���Ci�h���oGmt�x�sc��\�Fwv�*-���r�U��to��c��59Ss�Y@�����'KMe!w�(�"��,���n\�<ɹ�+]�9��3�e/�טR��J����|v��
��x�&��O�s�}ks�^^`0e.ԉ��m�Π*�X�P�A.��4�yr�{���ns-�� �̫A���G��#��������.
* %��o5��YԵ�ӗ�L��'�'A~h,ǉ^r�+W8��m����(�%/�Z(j�gBsR��<������)���x�V�kle����;fc�B�)W�4
�1�y�+W�wjP��g�p��s<�������HO!��<��ᴖž�p�E�����#��|W��W0�!>�P�`�ɸ�
�5�&�v���Å���|9�µ� �f_Ӊ���#Q���5���g�A���{��mN.;nw��{��B�N�j�nU[r���S�_f��٧̼4l!��?��y��o���Z&��Ț��>�mOe[p���pN��<�0��%��]"��F����o�1گv��C��OpY=m�#W����q��`u��Zzҧkkw��Y6�ȸ��ĝ��Sc%����V�9Q�7���C]��~)KS,W��� ��>�Ej�wH��ǃr륨�ݳO׋7��ȳK3�Q1�QZ��ɚ�3�3q��qV��9�Ƅz�.QY}��=TJ��p:�b]t��]\E�4�1�4�[y+��Ԉ!l����;F�7�w	g���OCW*����͋��{p��B��_��vbG=G�]���C٫��X�pv��O�P��F�J�6+偬m=s�H�Or�Z�}u��[K5�Vv�����D��=���y=�6��iь��F,R\#�oo�5�_
� �ʾ���+���مz)��ˋyl^:�c5S�����{O��2J�{O�<��'�թ#z�$�3�Qվ��)�dT��UC�g�ڃn|�ζ��P
�ﻦ�Z�el����1G"y�~�=;���j�m��4��i@{���r��0�J�������U|����Ϧ�'�=A���P�5l��a[9��;���U��ُYV������m��j&�mw&� ��)&�u[їB߇\��j�$᥾Ck)��Z�����9������pk�R�����e�i�h�#�ZpK��ymC6�v}2�q���H��{�U��l-��Tr�!�	ά�BB�/9k��Q�lL�������m���0T�k��,p��RA/]�;�oSy��Ԭ��>)L�A��u�eԻ뼏�r����I�u�G=�qjqvq�.#�C5�n5�7U���c��o����q�����
Y��yw�;�
�����u���5�<���U}�֫u���L�~�n5�+�ignN�9��
�1�o:���L���sX��W�y<��}�fK�F�,�SY���c����78C�y��r�vT��D�]i�n��B��V$H���9{�YN��>���*E���̩�Ô���BU׹Yr=�+;�or��ژ��9<o�\���`Y*9V���.�A0����OL����E�)�L�Y�~ʰ�Ş�P�tĚ��t�V�U5T�o��F4��'����P���_>]�L]��VQ���ԕ%�n��S�R�<�����p����4�|(w|���|��cG�(p3�%p���ΟK/�Rֻ��۾����]��i���ɫ[���Zԑ=�T2y&�@�2��|��Z�ұ"tGU%�{S��L��w��������� �e�t�wF�8�l�}z�WB��闥�;ӛ/vQ�cRA���i[��V��ٲ�1�k5�Ov��D��bK�4��}|�[�Gd��<;+9v���%���o5��#�P��\9i\3��>o�R�����\t�X6�^��IN!��Hs�5#A<�j'W=�z��?I�v�𑣾���ɯ�c�Qv��i�S�fg����j'�mw'��I���N3Z��K��ާ�T�q��I��}�J�L�0
q�uC��jt8�Їt�+���OwG���>ڈ|��6�j"�`�&�Z5��ִ��R�nC&љ1�N-�����՜��歯�U�Ns��iヵ	�k�W��"��	�yn*�s:��	����%fZ3c5:����9{q�sX��l�ھ)��wG�gSd|���e�A�K蒰fr����z�`N�Vª�-���Z��._j^��-�j�A~��&�_��(�}�o��z}������:�DXˑ�[��R�������՚�q�/�p퍃|@���)��i��f�R#�,�.�m���gE�u}t����xu�hڻ�y��늴s��C�,�eÁ�X��M�Kru�.�;�ef�M�Xٗ�岏V�{�YA��q0CJ9�l�u:�8w������/��\9p���f[�uwJT.)8�F67�|��OT:��w��rP�y��Y�%l��lfN����9<j:��Z�\lS��_ͧ���5��m�?Z1ُ
�̗ڒ� ��9mN�u�JT�|��|��=�m=���SV�!Cz>�V��u�:�RT�~��侇Of��x�5�w�6=E���5�y<X��R��^jcU���IP~	h�毂ί���[��d�R��q�Q�Gη���(�.��%��cV������������B<��d,�H���s;OM4������بv���]P%*��@8k��R��K�`�;�u��h��3M��hTgʐ��5�B{C�v�@��t/[N��OU[ܡ#���T�F�����P�`�n5�Y�nQ�pu�T��)+�{�o�{��B>�ΞGk�F�6�9=�3��MY�Qu"d���3>\��]����5-�C��3ʛ+�@f.Ӕ���T!�sZj��y�v�=�6Rd�ɝ��l��Wiހ�(N���+Exʒ�>d�pj�A�V���E_VEIc��i�nݼ��*]W�`l�Ҵ���/�ڋ�'/Z�5n$E�^�[n�Y��/>���������Em�^i��Ԟz;s��G\=���;��vn��|� f*�|B�y�bz���KO6�^��;j��L����oc�i���n}��2�{~�R�ǋ_^[��I��a��I����z�����绎|����o~�1�Ҿ1nwc��mD�����
�69sa:Onv�¾@M��h�,�U�%���
�<e�h=ϪFT�����6��Z���Q�5���ӻ�������Z!>�X'��X�D�k���6�(/:a�s����M�CF�f�ڄ�ۃ[��O܀邠�ʾ���|��|���<�Cy8�ܱE�=Kr���%<�H5��=��r��P(t�Ϥ�?��Ư[�WLئ���]��*�gVr����#���ؽ�r��!O}�}N�)f�EW��|��Pz
�Z�ta4楐��#�W*7��8�������#�I�j�����'���=���p��t[�\��@�~b�I	Ǽ�o	�#y%�'��ŝ���u��+.R-��k{C���xgB��*|�Υ��e4��jXIp噊��6T2DOO�r�p.2uP`%�s˞�ڈ{�i�j�e�w�	J�����o*��\��Ç\f������64u��^r�g���Ah�3�n���f��toZ7��3�O�;r�Ȏ�Þy���I���V�=�۽jzs�Si�<��w�W���S�!}�eƽ���f�o����߯�ov�N����kj/j��I��F'����N%N~R�}{*�JE�"{ܐ�t�7	Mˉ[������e>S/-'�>�՗����������q<�	t��:C����շ��"zڧ:�S^�*{޶^.��6�˞��蜗���_+*������D��@���&�s*y�\�-Z��k~�x��;qr�q=���Vj��������^ �2�ګX�-�e��pOf3<᥁��ml�w��,��!�Q�{��i��w׮��>@Z�]a�w��U��۔�)*NJ��v����k�`��
,J����tYg�#��n�_^;Jt�.Zr=�u�=����:]w��尢eޭY��%B��Y��Z޿7�垞A��X��H�<� U�ͷ�G�.d*�2����b��MX���n�Ʒ�Cyq�>��'�w�P���?�+p0q]u�ǐ�b�j�u7��WEӧSP�=|Ŏ�[�R�=]��0MT�SK��oj��Y�0f5��-�w�M|��_�k]��u}m��@�B��[R^��t�Ą��L	-y�B����rҶs^�R�1�V�ٙjso���,�K󖢿jA1���IJ��G�pt?D�G-�G`�ю��[\�ɏ��-���E;f~E���J�h?�N8�	ڹ�O���u4Q]���5�/�Lm%̦�4�hTdB�L�!���u��SMXbrb�0�ˤ���\Jǵ>{K�;mT�E���MƴF�"~�6����e���<���rz���q�k�yDc;5��=^�P�S�k^�Pg��1��MY�c�ʺ���%&:�.f��s�Lޅ[Y6b�e]w��m��W����rRG|8���z�<o�R�˸�-��ê�\���Z��`� n�ܮ�t�5�`+SQ��&�V��C."�Pak���p ZO�^T�Qvn�]H���}{|3yy�F�f�{4��j^�'Ѫ�g�M��/w����܉�Ac���u7̯h�v��E�w���>���9�&y�� ڏއ��Y[�~r�����*Jc���f���6�Ѩ��݊Kܝ��Oi��Z8�~놭>��paV}�u��$�&G�5T�կT7���>or�}n�6��M휨���\�E��E�[�ݮs��J�vzߖ�V5�Oyp�}p�>�5�lwdƫ[���ƿA�g�Q�s��F�o>�\�s��[��MqP�Eq��:��t���J�ק;����N#�hH���Eӧ�NSͫ��s�U]26�5OqE���1ƦHj��y��*��Cy�ςΣOa_�&]�S-݉�Y��eK�k��}��h�lc(�B!Lw�C{��_U�^��M�t�e���cq��9Ҿ�ݯjX�����y�֞��x���b�t�3-nH¸OV�)۷�PD�9�V���}.��=[��� x����˙v�TW#S�S��2ѹ��jm\���.�`���ܬ�]�R�C
ɮg��*�����|a1v���0�{��mn��Ofe�D*��
�bW�gP���
oZ�B��Я�^�.�p��t�l[�!Z�J��e��F]�4����2} ��w�4�v�`�atySISzF0�bj��؝鸩!#&�$w5�׃����Yg���Ω�M��uuk<�WK]�cgm����٭�+}��j�{6���s$��䒣Q�e�%�NC��U��d�ɫf
����J���\&c�R�L���-5�m]#5���XG;�Yg�YZwU==�E����}�V���3g�J�^�ܡ�_��@���3�6�]��9�>N�l�� CE�I��b����	nͼ�9k#4N ����zƮ��NBu�F��ؕ�.�:s$V��ac��)t����
;��*��r�4dW�S�r����Q�7�ȭ��Yi��G��s�{�O���MKR�[tO	@vKfe���5�Bޜ�WW2���fc��2�:.ʩ��ӬiS�Fvj�,@t�5{��B�$�Я@і�qWm�o�V:�LR�Vֱ�4�Ƅ�qX8!pѵZλ���Z�n�V��9�L�nFq.O(+�K���R�w�w�5p��iQ���n��ɖ�����ш6̈́��BI�F��r�D�%��y��7s��;�D�V8D6��h_EH��hS&��ai9�Ю�Z��+�.a�e���;6h-�TU�������4�#W���ӏ������6���ҝ�u�K��֝q�K>���G����B�u�O6��4�c<�'MC�;,�7@$�N�;N��\�,'"S�V�����Bu��H#���@>,}���c�WM�}m�u��<�Ex��z�2�`ތ3JW ��7��P:����L�V�ľ���Kn֦o��/m���N��0,6�ha:c�u�z�k�޴6�;F	2]�����$��Q���,�M,�G�JaaW3Ӗu:+�T�j(!���p��(��(���Q�ow���Y��m�mu��<n�r��N"6h�P;��� ���*V�w����«;hBQ�C;���-.�;��8��;�O�:02Z]B�iWGO�i���n��Vd��Ρk\i��*��l8C�6$vUX]�.��(�Җv���æ'��0����S��(��n���^�ﴔ����-��(�s�n����A��Û�!����V���Գ=aەj��	��˷	�5�,�F8��j�8�N�'Y�u٘t���w@Ŋ��Y��\56��<����U�9�t$j]|�������T�P^�sy�h(u��f��43�����{6��^���-���*³WN�.�:"����ڵ��bP�H�J��H9
�� ���d
P�@%
R�
҆FE�ДR��H�+@�+B�HҔ�Cf*䔪�R�RRj3�u�����i>��_���ѵ~��Ǭ�Ӽ���=�o�w�r8��C2wl�JMΫSQ��+S���|,֥r�&@�"�y�j9�]}��ʄ�V�kx����C�g�B�)�Bڻ����,%+�ԯ��t��3x�Oxm5��6�;�<a��meC/�Z��fDa�ˆ��xy��XL��ʡ�Y����G��~�x�&&�]T�3�%��;'�����m�W���<���J�˜Oj�5mB�|�k�nٽ�6���%F���|��/�z�U�U�Ƿ^8��������֚M�=���rG�A�}����j�D�����)�K�����|��-ΌVL+X�<���.u��'je࿚����;����7Q�fW�]�>�����%�糩`��OOT��_�\LGcN��lg�/__{�(�{ꙛN���S|��Ӥ�V������uV�	p��p��.l9O�-'�{�nBB�j`Zu��^�D1ZTs���k�	^�J�cb�9�}���3^Rj�V��K�m�*��R�V|FL}����r$/z�t�{�5�S�t�bj��H]Y.� 2jü~Y��'�a����Գz�7 xt��:5�ԣ�k&F/4���T�F���a��vwKk ��K<+���5�{�ޝ0��$�ܸ6v(�9q�|��_9�P�Fdq��Ŏ�p��<b�k>�K~��TFzyh)�6�˷�	B��$�ԉ)x�S��_���qOf�S�����=i��)T
?O���e_��l������B��'���q�����S�e�w�����u[cyq\GX����<L�ˣ��H�}��N4*����ow\ҿ��k��|>���W�C1[�nko��%�6aJt4�˦�'�=�[�{�j歗��C�^l��t�O"e�йZ1���G�9�:s�Z��m\w'P��3���88y';s�\���H+��k�F�a;"y��[A��[�s�����H����ڗz�}at����j��ӆ_{վ�6��S�*�X�� ��j���}��r=ik��{_^��Ns�8`׸�2q?)�T���N:������ί�X�&���<��8ݻ�����:�cc,m�z��ow�+��t�u|RЁ��ڎWg#Dwwh�s��ro��R�:���;,���[���0&����6%��MR�ӷ�hO�cC��-n�;�=Oy��ѝ�����F�f�{)�]�(������+n0Ec
�t;����5�Zј7�?aE��D���Q���T8��n��A;�5)�C`Q�����'��Y��3ǭNt�c���gR������Y��8��m�HWh�՝;��W�{g%�	�V8�A�eIp��k=�B����M�ʒY�dq{<��j�kG��Y��1 ��ni�$f�k�w���r��o u|�Ҹ����4�C��N�H��ݳ{b�c<�м�������D��
躇N��'��[p�=����)p�2�#jc9WT� ����ܦ�r5�ԕ����C��N_e�Z�c᝘�:*(lזӄ)�<�޾����zQ�*�HhU�r�Qy��G:���-+��Fl����ۛO9I����ݢ��:�8�S�%?Z�~X~�Pt؝e՜
{��B��s��vWQ��.�q�t���si��nر��!E�ɰᙆm��|)���Ew;va�mZ�g)���q�{����2��[�e�Pw�$CE�f�ܜ������AJQ�F��ʺ�u:�jN��Ӹ�X��:gc��N�-�Ӕ��sfZ���I�^/���m�T;fQg��R����ʑ�X�@�53���F̾���_G	0ӄ�TC�6�s5�o���q�
�T����S���F&@+7����i�.�pZ٨���W���<m��\�q	�ց�vDWN��ɝ���AN<G���u��;u=�Q8���j��K��q��/�F ;Y�2�Y�N|;���y> ����^Ψ��^eO-���ڷpԽ��ԟ���w�:{�6��FB=��N ��[x'���{t�v�9՗����݌y�)��'q�5mVm�m�۳u�e|U�|�&���{��^q�5-)�d���=X���<R^�趜��=Y��9(;�*��ǣQ5u��X�Q�����q�8��Ot5q\*�cb��{�����f�򆪖��T�g&������v=Bi��g�m(*��W[x�z��|kU��V2�t�Xs��iU���){4F��bц��
���LV�i��U����v�[� V�+�bd|8(�C�i!��%��a],te]ҹ%����q)��^���8���"t+;c����[	�kd�w�F����}��I���ɜ][+T�͢;�]���U�,c̑�Æ���ם�u��e��*`��ڎ�E�{j�:c���wu��=���v-�=SW�[��5[����^�~�5L��f��τ�W"�i�c��Z�r��7³�M�Ňi�}4��_����O�[b�EB!Lw�O���.�r�#����r����֟�u�����V�ky�
���P홄B�z��,R�.u^�Q�^:�bz݀��X��w<�F.�[o��v��3�Ց���i�kU���S��?�j&�m\Gr�\ä��$�+��j�ժ�[4s�j���L֯^���S�MZ���4:6�/����1��۱��^{J:�ŪH���}�M�͈k*���L[P38���Z��Aב���p4�m�,�*�q�^�؜3�h滙��W��@�u���re����gռ�Yt=�}6��Z�Ύ�st+#%�z6�^��{4��N!���{�)�[&�W3��]��d7v���M���ö&�҉ݡ]�[�<`v��'%Y�߅ ��m)z�uM֫:y_Vc�Ws�F�sI��GW�V��S��u�*��&v[j�v��g^�ڷ�d�O���|�e4K�j�scדsF�*�؝�׻�3U5^cu˷�@յ78C�|�c��p�S`�{����e�vk}�����]ڄ�,����-g\��p�����p�=eE�t˞�8M�%��Qp��~���A܃�9��-W@��\�9��)�I�9Hn'ڟ\:���{l̠2`󁽸���o%��`�ލ�D�$��	���ƶ�M=�5�:� `/��8�s��c�����՚���e����G��_'���X�vT+J�P��C���\���󫖯�C�5�}���S�/�,}��Ϋle9C2T�p�d�� ��p���KE���q���_u�Ҹf��'�śe�����K���"S�8f4�1�F٠��(�Π�U9_���U��,����m
�dP۽�4Z�f���5���ow1�Bϫ��F��R�7��||��T�:E��]X0������\��p��Q7u��m���ْ\ʲ�����栣i� ���N.�]�}j*�0*�mv�[1ط���o��Im���=%��=|r�&�v�FT�������`��}\;�kӫ>�� F��B���;M�Zw��c�[�[a���V�?��)&�7���T��:��-���m�����Ls��.ʪ��U��gb�3P��w��k�'�"� �������t/}��^�5�׿T�+zz���$��ALy�X�٨�3qُ1_=AG'�ԮʞZ6��N�^�9yi8���B�U0�@���*�vңU�2��?�K3�<�g(춝�R��^�c	/��9ūi��,o�O�#7�+����Q�y�t��zV���'���n��3'��:YQϷm^�^��A�RuN::u�;19alY<�zQ�2�{��K?&�]E���i��WeDRf4n����ӽ}�3���:\�@u���n��g���x�-<�A��7��ތе'z։�j�-H�h�������
|i����j�x	l�E��ZhT���,.�/�W��J�\s���X�m=�PŚ�!>��a�WRqgQˢ-F�������MC�K�8G5�^��=��μ�K�gN�;�\t���ET*U5������|~�q&v�+Z�V�̫��sO�﬌���
���f���m:r�i�yp���> e��&���|}8A��r�E�ٷ�R�;�H��~�/[�ΣSێ���9�5��׎sU�X���r��t1�\�\J�3�}���|�@��ٜ��m�.�lLo��m���<=�mx��z�����2O
�2�����j�#�K/�~im,ЯR���R�}�LoDy�����O�����16��3"�E��/]�0at[׳u1htb��އ�)�S�hи��O��T��C^��Ǽ����o�d���{>f�v�Q<�W�'��ͪ�	k�d�3��0����Oe`��U��ަ:ڻ��~����=3�w����Ę�T]*�YU��%�vh�%�"���P.a���0���n��:=��ǅ�^_�f?hRd����]�=���y��st<^}����B���e�v���Q2��<��'�2��}�f<�4+�/�-�Z�{K{�[
���ųTռMp�N�Z��Vp�{��A���p����yj6�YHm̭n�����Jr6"�U�JZ:.�RĹq�ٴ�%1�����5��s����S�e.�Q\(F����2�t�g2���a]�]��-~���W���P��Φ7�n�WzrNZ����xh�a�}�ީ�O�����,��ۚ�y���O�Ҡt-n���2��s��&�9b��Xl��O��_^E�N.��e��wg��^(u�J��<�y�;>���^���^����7��#�����c�|f{�1��e�Q�`:��,OL�N�[�;�Xx7��E��z�7ߗ�G7+�QX~m�w�'��R~�)�ӛ�q��ω1�Uએ�~N7����ʉn�Ѝ���ъu�G�.G����T4{���!����qȜ�Q$���=�a@���EN�E/UD��FǞR�}P�*�I������vS��ӿi�>g^���7�R6�S�ɟ��=�RP��Ś��Ⱥ��뤏�mt筛�к�Q��W~�ZG>����:�:�{�Fߦ��s �JEP�b�7n�Ѿ�w��ۗ�w�z_���h�n��7�F�7�l�G�z��Ǧ{I���q���
��n�n乼������NǨ��+����]�����+#��5~~���>��.'x�S�Lk����ܾ��ʊ�h ��u%�\�{^Iaβ�5���_m��P����v����}G��s��Jv��
$6��]�1Gq����MDDC��Q	�y�0�뇵 �Jg'-*��j�Q
�aG,�n��2[��5�\i�r'ܓ�˛�O�U�_:C�c�%_��i�G����iw#������܉#�_���z���_�t�+ȟ}�(Y�w|�w ��Y=P6���y��!?���Vmgz�~|o�NN�F�5'�c�鿟��q�<��ʐQ�+A���مS��7ޏ=5f�E�	�t��f��{���U�o?W�����q쨞���B��d�d�|h��{mW��u��{���J}����D�zN��R�o:�ǜ���9�VC븞����k�G�����ށ����^<z��w�=�Ύ����rN���^&��,�w	�?g�߫��+>~���Ä�C�>?��8�<i��d���T�p�'v��\���q]�9i�q��:���Mz�
��/}2:��K�@f��\\�{R����ɉ�۩�qg����,5񞨨��zOS�Q}v!����Wy����+K�����%+�r=�c�=v��5<5vT��,����A��O�>S�������eʟ�/�l��^��,�}^��'�ٞ�Z}μ;&낿��UB�	3�,��(kxm�{CV�S�^�N�V��(#k;�D[��-J4u��61`!-�ʹ;f�r�j�����%�:���LL��f�Q�pvb�k�3��friO��vo<��9���51�Y;�Q}�����-��R�ַr}w�$Ri�Z�֎�2�u �f�vj=�cN�̨Up�$n�.!f�N.�����12���~A����0�=xh�veN�iF�1��r)�Ԯ���˴�`O��d����� ���:S�K3%fA�K"��V�]��tm�	".[���ݼ���1��+�\���u�fu_g7 �iP�@֩*�N��o[[]��X�mb4��]�֖���n E��2N���UN�hܼ�f9I�h`�k�j<<�Qpj,��(l��S2��Z��u��@ S0';˴A4r�o���E&����( �d�@}�fb�l��Yt��'[u*>f��PT�Ǟ]�J��z�8��g�G��èk�m�Y���q��q]��H3�BM�V��]�N��_>Dn�ƉX��Wc0��g��K��#�P5˲`Si�2�n�'u^G9��h�5AW6�����V֧�6���"���7�n����}�o������Wմ�&��J��j�<�e��ҥ�N���E､��U�H���J�+xx��ќWX���2�2Y��m�f�`u�'���M��Q]�+��uH�T�X�r=��Ky7�ѮR���Q��Ȉ��ɘ��u� z�IWP��f-=��̶ƶ�W"]k��O��V+�U���.�-��QmH��n�w�W��2�Vt"���:y(���vf�Y3��0����Et3_0Օ31��o��9x��v�B�.��,��	�Xpӽ��VyK{'H����Q���{�u���,�]j�7H�G�Awݯ[�A���־%٩iI�_�9u.�W\][R�lᇆh#v��
G-��QJ����d`t.����H9���K�
��c�6o��&�V����f�L�����q����򓴝^�-WÉ=4+E�ŋ���DE�[8�؅ˋ_:f�n�lc�l���)SxT����4^o�z�.�5 MT��J��2�j�e�����`�g���c��5�;����W��pf�"T�*f[�4;ѐ����,�&f���[ �,�b�+D�3+��}�\�]f������@�$,���z�F��4��/wv��c;�L�5�u�	uN�jͫfR�S���*�k��X��	�^�-쾠��p&�oe���J���-w9rS��vor*�G/XU�9��cg]�"�p����J�U�����[�y������聮{W�ej�����KqI��bPy�״�j�E^.HTB�:fH��C�wh�DPl��>ͳ%nt�l\ǉ��0��[��9�W�8���1�n]�^]�c\���7�,����	����@T���	��!C@�P%�D�P U-1HDI@�4�
�4�@P!H6b��U@��!B�*��	CB���	KH��-4�KMQC��%+@R��U-4/�^�yu���w�u��~����N�U��B����d���e�uZтpP�,�__�U��˷EgО�t!4��ᓴ���$�rsk�^�Q�R����|o����|�{�>+O��|z�ڮ5�e�@6
.+�<�j�����Wnr�`j�@G�4�PP��Yȇ~�+��B9���;�Iҳި8�Δ�^�1�gۘ���l��,��u�[�"�O����ֻւ����_�׶'H�𨭒u������Dgu��Uꉯ���|�7Bx��^��<Z>�&��Y�Y�ݸ�۾곔G\^�}KW�qR�^�&���)۸��2�z���l�ė��7JZ=~�sq�n�U�{�Ѿ���:���7��7��>�����C5�S� �t�tQ�^#�����~09N@~��ZjG<=�=�|v�{��n��{>�y�Ѹ�>���|���=�%D�cJ�j�H�a��o��z��63�+N����7�鿡�����w�3_��&��j!��*.��Su.�څ���>G�U�Ɏ�8�T�I���oS�λ�^�nF7���#���(�M�SŔ�'&���]�D�C��S4oO�ݿ��u��ϴ�J������i�s�Q\��{+J�^TeqV��o�bY՛����¹�����9%Y���>���T��M�Xq����vUgK�
_���Խ���\�W�;����(�eY|�ۗ��s����q-�D�k�в��}�y��嵖��ŏh�<����T$5yք�Y7�jf��J�	{���Wx�~�������	?��1�C���X�4!S��`h���t��{�M�T}`Gk��FC�^����=6���d<��t䝸�d�T�ѝ�^�����=�^�yռ�S�>��p��T1�'��^�����Y��E_�K΅����Oiٚ0�'�lzծ��s�
	��J�S1q[��s�7���]�C���u�o��.]�qyѮU�	����P��G��s�|�ԯ��K7�X���_��!�c�O�z��⭁��V_v����]�ƿA�f:��f�D��'�/L�=-�ϟ]G�=^�=/Ճ����8c"�����tu{��|�*��|�T+�rQ�� yW�~>n��=+��Q��'�����P�g'ֻ�t���>V�}����k�!�߷�#o�Pg�2T� %#Ď������6z{�^����=ƭ��oˍ�3Q�߹
��o�����x��ׁ���z�s�j`�̐�)Z'�y_�q�L6w��G�y�qN�<1)~7�*:�<��M����<|3ɚ�*!͹�W�1*O��۹�%JPA�f��s^���=���]ˌ
��f$�V�A�4v~|-е��]��QMmm� �qcy��ޯ ���n���1x=�7��c*�;��u��ՔQ��9�����"[ǈRy7,@w"z��OJ��(\��K:��irT-�Y(7�3���-�r~#��̨o�`��46+>7�%O��ת=�*�0��>~�@�]�o�c����o��^L+�G�g,�<<N���+TOe`��{��z�놮�1�	��:�\����z���*�7��xtϣvX���{jE}�Ī�s��S��;�G�7��^o{���1*��q���]��N���ޡ��=�bt߲hT/eH��d�@0�h�T9����tdt���ݽ���Y8R,z#q��s3�s*�����uq�Z+�9'`�͉���
L��|��[���}=T��ϑ<rϠR��,�eqJ[=���劳�
'G�r$��̙�ow��l�e��|;+�ً��9ó��7��o��x�dW����F3F�f%蚌ټ�zy��7�,�ݦ|<X����&��nz�<���-��xkv���}1�@v;\�'8_����錈�ʞ7Q'���>T��uR�NB̨�p���m�􎑌i��ލ+܂���G!+�s�D{��c�M����,���P$�TWӲ�V��O�u^e��N��xpJ�<�����`�U��%���؋b^[����Wc�6����9��^W�d҉f�U+�Zܱ��K�]k\�8;�-;곶j�u��iu���hs�Y;`�Հ�� ꅹa`-٨�V��"⮟�8C�h��N��<����@��U#m�0�&c��5P� �U
�Ϫ�Х�仦ރ�Ӿ+\�"��QN]wG�w�q؇�Я=�#o�L�C��ۮ�{�Y3-��k�ޤ�È�G�s���@�h�l3���*�o�ه���;��o������M�\ɋ��l�e����#�zd�50�c���r�������<��Eǽ�gǕV�?z��}������y���s�]e~U���1�J���[������)��;�mz���q�)�>����.�g<���=��o��;�TX�r|��ƾ�^`��h�Hw�VO��u+̝�{V�O_w���E��t�NjO�����W����b㽕 �ЧĪ��gfg��W��N EN��~��4Ϣ��}��^\\s�{��H����*'�=�C���͖��}��vh��O��J�l�C�R�]e!�J�����~7�n���k�c>oԼ^�]į�z_�c��>��i\�~��צh�ǎΓ�FM���R���j�E�G�K���3������^���9����w�)��j�#L�,�V �鴞��.�6
�sWe(Ʒ:�"Q�#/'1�"�I7r�%��Pؒ�jLG�dO�l�4�S<�@�V�Z�۾U�X�u�(\�֞���V�p��3跶���.F<rӄ��"sV�}�C��Ռ�+�Ө�wn �<��X�[W� Ӡ<���)�x�<���62�Y3]��Rρʞg}��'�FvT�,� a��=P��rz����'e�{�oz�*5�~����J����LydG���Y7\)vT���<w�+Ơʨ~w|�=M����ǧo�u�����(��UG��}�>>��G���n�;&낰l�P��O^�)
ٿ,r���)n{�:����{Q�UM��g���O�=>�)>/�{����T=�Q��+�݋�=��#Iɾj�P��A��A�|��f�t�X}S�+��B���CFC}�h�yIҷ�l�xG�W[j��^j�}ze���_( %E����H��J�`�I��2'�v���n��9uQ>�dKY�~�s2��/}ʗ��D���b[2Y�@nzz�WKGݬ�k������_���Wq�\�<S�8{���ldz}H�g���7��������jϦU�!�pzH��_W��g�3��*1l�e�b����w�~�L�11���I���Hg���{"�Թ3�Y<* ̿��!)1��?Q�P�]oB)�c�K�r;��uk�3���<@܍˰@�-z��0n�[�~��;9�3~T.�?A�C.��# ��ŎrUh3���s636�gWL\>��U?�ms���Z�t��eC�����[3;a��)���p���
���=g!)���mǽ�UE}�_��?z��g�����>�\)B�c�S*��y/E�D8����ԭ:.+}��{���j���~����>��;M��/]��k*+��g5Y��ќ6����W�,W�Ts�
���`>L���:��/W�!�Q���^�����5��{�ī�k
�<�á���az釵��2\�9����E�f�䜸����gؼ���G�UJ��wޥ��άof	����\�N��U�/���z�xޔڋ��f�.���n�J1Ւ�K {��F;��I���k���H,�ep���;qr��ۉ��*.0��\yͨ�{k�vF�>�wrU̨=>7��{��x��/��ey\og�Ш���:.ׁ�ڕp�v{�U�L��AT	��ʙ�� �[頽��W��mi�z_��:�v��qE_]�&�A�^����Ͼea�5�A�2���c+�\����y۫mz�8dG��1��7��Y�~��\�Q�<_������Ê%�|I@�.K�"����>���ǯ�?-��Z�7���ܨ�ԑ#��Q�������KE!����f�)�~@�����S�̳�"��hA�LKl������w�Ľ7@�e�U�W�!s�κzb�i�֛�a�ݖ�]\]��ۢ��ss�&�^��.W��Rp���"�u�n�k��7_!6u2j�^�6G�W)��Fg��B*��� tۧP�\�j<��10[�&������q#Q�Lߧ��p��gV1^����+��^X�|�k����!�߷�#n=TĲK��@�A��j��z!J�N���ywN{��@�^/wƣQ�|�G\7�l�zgx��b��{Հw�<f��-�iÅ��4`�z1o��>�*H��HT��:5�}�*;�W����'�x߉�`A�vC��u�w���bʟ���*�_K��u��J^��^�=q�+�1q�Y��f�f{�w��
��MV�BW����Q��a�i�2a�Y����ek�q��cW�]�b�EC����G�VOGU��>��^��·�_����^�;�2���U�}p'tº�n��/�����Oi�����Z���U]!�:�q�~��/=ׂx�̌�eHˍ�N�@8��چ�_�:�������R�h�*e2t�o�3q����ϵ̨~�^s��u����nM�t�t�v	��EVX��33���#�K93�~��"Qò�TB�;�dL��&�ϼ{!��r�U�gﻣȳ�|���m�WJ�ws;%4�m6����|��SE��\oO^ ����5��]��+��\������,����0��yl;������e^�X������� 0aǉ�[�o��#Jq���"�:�̎�bڗz�j��K�+�DT�������$�N?����_�F�TO��{+��x	r<�|v|���7�t�|E�߃O�JeD|
{ݽ�t#�RV�5�-{�Vx�DgeN���j�2�W��'�}'~�tqޚ@�W�k�B�n/X���v�p�h~]O�g޺C�����3Ơʦ.��O�!fTK��mP����_mʛ֪��"�<�z2	�����j�z������F�d�Fa��>U^d{�����SWt�J��J������n��*�N��#�O��o�q�j�C�a�6J�R �Ʊh�@�c�[�Z�������/#]X�r+�Q��z�>'<V��0��޲6��Lά��X��+�X>�Ô�{A��W�}DO��p1����9�n*C�׭��޿3��~��C�ʽQl�d�ol����p������A�H��_�Ʋ3�9O\Xuz��i[w赫��R��|��{Wu3)x�����&.�uQ
Y=_	�^�=�*_W��d��y�TǛ��r,_��.�j|F�j�܋��x�dO��d3q�?]H8��� �|o�쨨�պv|�������CF%
d�͹����݀��8�+�3���	 =GY�6�V`��h���Z�y��*.ֽ�,�Z���p��vM�����荙�e�kp�QfetFQ�T�2�,���]�Q�ua�n(pNmv���|�t�-�VT��Ftm����}�n��p�ߗ��2�\��~�=/��4���ʐj��@�|d������dI������u����0�4������7��Ԟ�J#_�J��eD��ۖ.�����ۭ�^�۷��c`��.P��gG�%�/Iңz_���n��L�t7�^/c��%Gw����es�����~�?����e�����=P6t;�����*U~'uKE�G�D�~�4�)��T�{�ܛ���9���;i�S<�t���KFW��~�ץm_�4�<^ �9J��1��f���s*����y�G��~>����R���L��
���P5�0��Y?$A��z�o<U��oj����Uxp�P������+ޞؿSY�<}7\*eH۹d�5W��置���mo��ǽmN�����rmܱ>6����>�i�t�n}�����z�xvDM�p��_pJ<�*������`$Ϣg����C����^]O���V*�<���yI�|s�t�����ۯF�����_+���=t�A�2��W��å����^�R~�Z1���Z�PY^ZߞЛ��֌�C�Gp��Cʅ�D�%;u{N,����=R'�0.�%K��Pn�Y��[_V�ma�]�Yt�q�����V�n�i�.n��)�c�R<V��\���5�ٲlO��ͧ�źЏ��
$d�Õ�-g_>[�kfZ����~���V���b�J	TQ���H�Ҽ�w�gB�}�AXQ��g�������ŵ��S��;ޞ�W����=^���d�_"ux�+��r�Z>���K�[0�U���>�}X�����z}H�g���6���.=~��s>�V�͞�4�C��Y4x�?'4�w�DS����j��ߓp��I���Hg�=^ w��]ӓ(�xM�u�yA�n`���S>�
�>�h����Yϒ�����{>�����&��@w�˱nF0���g�;��{�S'��0����_���ԭ:'_W�����ˇ�'�1��>�5��w�����.���j��_��ٴV��q�� d�Q����>Ӣ⓮'�7��_ѝw��כ�*<:U���W�Fr5�K�9w��:��ʬJ���B�{*p�F�N홅�;��W���R�Aؖo�9<�n��+�� ����ϡ�z�����S��>���)d����yL:�u�~��,㕻j��v�->�R�>�����d�w+ޓ���Ҽ�(Y\+:rN��'�j"2�`�_��~*�a+�B�	4��J�7��@�(|^�ĵ��讷M�Ϯ�{{E�YҬ���'����\�wbɎ{/u����VK�7F�'��c'*�(^-+�}����2�KBgAL�[��lW(QY+��
2ͻI�Í�j��=�,�gQ��'|�ؘd��)XPg	�`�[a���$U�7��_#�t���Zk��׷��+�ڻ�t�7}k����m�.��M����z�ŜF��̣ٛan�net�o�I$�u�[��N/��gPe��i6�m�Ɣ�LX��4����rȦ��Q�͔.������^Ӽ#�r*�t����2^Wu�uY�ͬn�Ƒj�$��V�kOR�i5�Q��Zf�eK�f�3Q��E!�*��p����3T�ڑc�VUuٗ�M����n�]��b�[��
�6���m�*oI���m`�5n%ƭY�IwT��ֺ�CbZn���-��7�N�AM�i�|S����Y�
V3pܘVT���,�d�F�KLR�pfL{�2��sC-�"I�L�� f��Ho ��g���n�I�1�wv��`%����)9�Orh޽��魓u�a��������B^q�{��xj�oz��e嬤Ӧr��yMu�5��K��[���n.G����w�*�� �o��Wձb�:����	��s�����W��a�q!�\ml�B.G��7i���p���Qe#R�,6��e>�glX���ͦ�sB���۴�i�E�
z �XX�YՀ�1�ui�5N��E
?B�gж�e�,�X�.+w:Sܠ���C-k�����a=*�QF���<����Q}����1kH��5�Jl�f���V�6�}`�tL��T[9�P��u��/�[��w	N�v�s�/&�[�T:���E3��),!2��o�IF��6����iW	�Q���̼��: {L�\˂�V.X�wP�j�l���!ɶ+6��Ho6�l���1n��˜���)�����_d];N>��,��J�ui���O��j��c���Z4p�%V�3EZ�2W+'(�gW^p�;�v���J��y!��]2:� �jd�v*���+w�c$E���S�<;.�F9�Qh7E�J_K%�ޞ������Uv<CS8��twPZi��<�E=��,N}&!�#mJ�G��6	�M^��Lk�r��#eکfn��ϕ٦1��g.�����X�O6
��q"跃����7�Ư�*�̕�n���m������΃�#6bN������@1��GwoqCf�QER�*�WA���y�Qۙ�5���(�:�]7�7 t]v�˰�
�dٲ��J�[��"��{"�^=�f9��
��L�kn�����!�zԩN�`�ݭ�?�e]L�ܿlۼ�;}�0V\#"�u@X/J]��Τ7�oLT4��ܶ1!}m�`�[R���|9ŕF�gط֍�Z�WDґS"SH�IE@�C3T$Q-AIT�!@���IM4D�!AMJ�f`@QHRDEU@SCCM%U%QER�AT�&Y�!I5PADIKUTU%TBDPUT5CHRSKTPS4QTM�%5M52QUA55DR�T5$TPU4%DPP�̕I3M-U�TPPU1U��1D�HDMUE3�e�4٬|��Vb��sGa�1���zS���9`R��%*��`fX��y����o^�9GmJ�&]>î�\7����;bt����XyK'��*�xu>���Jex�]�������7��hz��g/P��*U���W��<=jI;_L�ug����L��\�>�Xx;��o�G��r=�~+~��z����}��q;V��v}�m�fYط$�@>E��+�\�嬢˧4+a�_�������+_�:����|zߝǻ ��ÿ��F�U`@K�#:e�9��},w:��v��e��B���]��({i��dy�y��Tt���p�P�\�j<��/��q>���kj�}{fi��f���a���F�y\U���r|��O'���H��SP�K��� 7.n���W���&ף'���{��z}��n�����Q��Tm��l�zgx��{g�{נ\zs�v%=�;b�{��Q�]��3�ƥ�I>t�J����F_�����5~�o��O�|}9������?ɦ��;�_���!$zg��31�p`,���t��%O���#��+�1Ք/�L���]T����9�2}�������}�I�E��&\	�����dV���ަ9Jt�x��v<���<R� e��"k����k�	x�0P����j���P�[�{����n�Sk�@��=Tܖ�<�yH�!yKe=��5�{Y��\���l	�>�Zٽ��cܤP�����sn���A��+P����k�m Q(�0k�Y��H]o\Z�s�ϸhԪ�{�zfߧ�OZ�h��ɐv#�Ī0���;��^�ҫ"��^�����_��d���7�ҏ��~��c��m��y���}�4��x'����\ȼ,�P�[qzD63(�=攪�E�)W#u2��9���g[�3>�2�1�O���ko*~,��߄����W���&� ��ߺ��f>��V����<��p+�ws+��ώ3���qˬv���d���K7��y'�B>ɖ'l��S��:::s�g�8�W���x����ζs�ۊ�]��qs����n�=X�TgeN��>'�̱�2"���n#��e�ýV��a�(�u�N�f�V�0����¯Ͻ�~+>��Y���*Q���=Fa��T��]T��x�
��y�-�v�v��6��s���!B~�
#�'�;��=��[㓓�E������#8w �GE�K�5��,����ۉ����*����r#�O��F���������v����ye�5c:6���{]��� �>�(�K>-���ƣ�;򸫏W�"���D?Hҳޢ2��sŋ�vL	2<oF
�7�3�j�=�{�X`�K��c,�9�7�p�E.V�:荆7{*�����#d�Yڽ������|�q��_һIt��e�컆��B]��[C[2�+Ċ��復�=}F5��.�.^;�X�Ř��.�Sowu(���ge��&�?�@,1���G�.H����n t�7~u|��^��x�W���M��3����P'��|���>�;�'�U3"��jnL7$d��4%9^:�f|=~�dw��qG&oхmI��:3s;����}�ݖs�;�^G�F��n�iK'�L����0_O�͖�m��*��E�Y�ؾ��W����yUH�m׉�@���C7C�\�JY=P��ϲ���5	_}S���^Nx��䏢���^o\{��^���~uro�M���>Ϡ<��ʐj�����k.��*B��_���gZǋ���1��y������O�|u�@����vTO_��c�m����V��R��Z�Qν{3^�<
#
`l�s����<r#z_��[��:����oԼ[��p�n���JsK;�]�W�V3P��7�;;s>�l�rrN���W�wT�׾yS�8����󔣖&��*��?U�쎬��ʝ6�'v�3 �6���ύ:�sg��Q7��/}�9�����'~�;^���~=���<��S�����0�������N؅�=M��=1n�޹3�FuWkCK����)N�бµ�j]<+�J.kobӃ�2�7�,�x�T��R��F��Sq"w^�®�Nj��729���k:Y�),����=�11Q)e�����/�b��ld�cq�@s{� R@�[9��k�wߝ_z�Cφ��E��W�=�=ު�ƚ��23�r�<z���d^p���[��ޟZ ��z�ғq�(O��wp�z}�G�O��>�\{�r#��ò"n�*Y$(�z��H�!���>�{�N�g�L��uSs�.������U����s�)>/����ޛ4�)��kw���q��q��lj�,	
W�������=~�+��C��Ml�w�<�gw*8��=���g�pw�,��%��A!�"��-����:����#��L�{&�m��t�Z�=�ο�����\OO�'a�,� 7P'������;~��\��s���qr3�Fי��q�XGo��ȏO����n�\����ә�ʿ��ٴ=}���kf������W~ �����G�*�������5~�~���� ;��`�ə�d����e�,�̹k|�yz���ͣp\ਉ�VRg���K�5��D{��2�L����+_vd��7�]�N-�=�^{��'�9�4rX���i�u����z�j���1�ɟr��	ʡ\�F�\�����1}��!ȵ1�^X9z�}7h��"8��uh�+~f�qՓ����U�p�\�e�R��:�QT�e��{*��:��ʏ\U��\t��.�3���Wf�H����]��5��pv�˽�,����Gv�z=�}�,O\7{f��L���W�j�mhwS�:.):�{#z����ʚ~�N_���.�j�>a�7O�5�GzS�*�*��P����ƖN홅��a�e{�躁(�����'c��	.B����=�߆C���3��/�ucx���ʑ��s7�0��zr�dUT�^z��u\{5�Gў��D�"W@����ײF}NW�'#�Q��y��
#:rN�pgvU�g�7�f�і��o��艗�������w&�}����v7��n���ؿm{�M��t���~�[���3��gy���A�m?U�D��/�������)��>�Xx;��n=�|}��]�nK�Vz�j�K�G[������F��$��,	ȱuԮ|i\�z��^�6=��@���W�2z�J�!��,{�U��>:��ǻ ��ÿ��EV�����G۞���@���x�g׹���������(\*~�}^eo�Tt�����t��.K5�Ua�7�}���QȺ��Kzo�O�=;�Y��ny\W���P�k����!��}23�,K�̗+���X�n�/�w�\MT�u�#>���Ѡ�:��b[]͠K��.\�P����_b|�=a
�VeJ�Ƃtl�oen�r�]Cؚ 1�5ɽ�FD�6���,�x�v�����y��qh����v���*i'v̓#��վ|�-�5J/���I�Y1y��q���Y��& .|\�w������F��	����s�;��;��V�q�z�o\U������V=eם�zd�f�Կă�J��M�~/܅G\y�����O���޻����ه:ę�ou<�<'=k ���H?��1:)W~��5�?yv��r�����DzP뮕%[3^��d�����WyяGo�fM�?O�w��j3���(2w�L>��1Q-m�s�7IS
�"Ǎ>�S�[���c1�Xa'U#�c�L�C��	�^�/��ԃQ��U�}bwL,tg�'hU����g��?�Ҽ.TƇ�y~u^Gz��<�^	�q��{,����t��˃y[�^>�G�:����EL�Iӑ�_��u��s3�s/�S�}��(�ֶ���G��V�2�������09���]Z=t� w�xÒ�T-��:���s���{�(��g���*��m�vz1��lu�����Ӥ�y&x+�+��xdA�C�F� ��}~�O'�pc!߶p����IZ<��x�C�qݎ����A���Xʀg��^���2����D��y*-H��B����X)�_V��m���ҋ��λ����6�{螣�Y�����"|drTdԦ���t�\��u��/�j�f�.��V�m���܆�._յ}�v�;��X�\�+�n����S��r�njʕ[@%��7�\-m�*ѐ/���N�*���������h�xnG�O�z�r����R�I�3Ơʦ{<vp��E{�'u+I���s*%_��b|�z3�'�;��=��[㓓�X�(�ȲJ��萲�z}xj���,p�
ɇ�t�o��|Tz��~�~ӑ�'�{#}@{���U#nS��߮�籋��ޚ��aS�w�G��5��?z������cQ�~Wq���s�3�+���+&��nH���Gl�9��S�;�)�f�L��JETD�"e��c��c�Σo�!���ه轝��Ǧ3�^���j�����L��~~���ό�I}*L7$dI^SB�:^<������^ƙ��K�=;��b���������Y��L�y5Ә��K'��^��`��Q�K)8b�l��>��w�.o��^�'dx_���E����<|�C7?e�5
Y=P����/у�o4��G��8��-�i�>Go6��W{)��ԟc����}�U��̃�{�Etz���{w3���%�B�l9S�}[>��w��7�yp�?]����ҧ=�Q=�=G�k�YVNȮ�G��]$F�sι ����-�O	�*���1����l�j�4��ҭ2���S:��dwH������I�-�ңk[�Up�7㫨��A�e��ʯd���FG�VP�m\����=WÃ���%ezJ:�r�����g?]��m����RS;����k3�g�F�O��:Eexl�|N��z_��[��D:�����L?��V���6�Ǫ�
�j+�]ī�՚i�38m����6t;��:.*U~'r5Sp���U��تfr��\�]�4)[�����cc������7�מY��ֳ��_T��l���n�yE׀���:�}K�B�k��s�OǱ�!�s�£;*t�d�q�xQ�p	׎�c=�ߒGў�wrU)�@�]�y}�"��+ޞ�e1��<5M��254��.�:c�}ܒ�a&I��uu�JOQ�z;�qޟa�������9�^��������8G���n�<D�	;�@Hj���]T��l[�>>�M
�u�>�)>/�n�뛘�Q0���]��<_�;���x�
8���FX�R�f�t�Xϟ]o��҅+�h�R��������1��B\��+=ꃝ�a��( %G�A����y���N]���vֺ'7�m�/����ZdD�;c=9����.&��������2Y@��1�����o
��;��NT��T�$��j�l+����[�*Cp�+���>'@�|��Yˮ�qmk9���v^u�iU��5q*�wT�u��fR��s&�������<
���R}���:�'J�g[s���*J���>�Ӳ�X��<���'�;WNyQ��x�߼j5�>XG��3�O�����_�8�~��s>�^^�M�eGN�nF���rM	g�I�*7J|6��������IQ�z�>�������=�/�7J*����s���&Q�P����T�/�Eme/����6׶��Ux�c��d��<���Gt�T�cW^cT<�ٓP�<T�,tx�r{Z��/>ާ��ˇ���S�:�ߌ�T�j���ޘ�$�'�|'{޽�q���q�*0�Z6�9>Ӄi:�{<8���jz���z�-�c}�;�d?W�#"5������6�P�^ʜ7Xݳ0�BsL2)�X�x^�_�f�>K�;(�o� *7��U��gޞ�O�:��z��̋JY;���z�	jh�Y�U�z9Duq�Zl���m0&�r9^����Q��y�K+���H�v���md]
ˣ�
s�%;�ʉ�f}Z�����,(�,��)��0���ޑC����G1����'�O��W��#m/�0��P���1q\�7�V�x�tQ�T\mPRh?�/�ip�i����y��;�e�9a�����Q���7v������'`Ҟ��R�e�L�5��^Գ/7�]k��t�U���'9�r�7/��H�Ύ�����n:�E��crɇ�wp�#:/$�ˌ�{�c�=*z�*ᑗ^�%C|t�>��_����� k���ed��X<�]J�ƕ�ev��^f�/q�\���wN�[Tƅ����Q��~w�3~0�\�iU`H)zdg���8�gۗ�՚���]�*��T�E:~�}^eo�Tt����˘}�H�M�[�SS���wR��z�~�&ϥ��a��E��E/�^X�9��=�ԇg�Do�X��ӗT{�
'�;�\�^Fg�" �4}$LKu��å����Q���Tm�߭�����>��n1����w�(��Z���ŭ����=8��t�)���f�=$�B�KGF�F_�����5~����7~������y�ݲ�|�8FD����ۙ�H���w����?.��Cy]�Ѓ[c����bԍ���V��o�;�1|���7�O�w���>�$�Y=_@ɇ�}fYX������\SV�7�[�m��5w���O�r1�G�T?O��^�6;�Rt��a�f��]���XF%ꄽxb�J�M�)�.U���_�G�W��ޡ�O=ׂx�̌�eH���锜�é� ٘��;����D�x�E�K�W82o{KY6��`�,��է� ���@�ML��Υ�WW:�rN�-g=!�e)��������80�2�������ݲ�!zc��.�ŧ�fj�\�u�K0���3�^�B1WJ]Q=֘p���۹l�O�������=:�S�&I���ea]toƭ%GPۈJע�]N��&)��Ek�v�gXG�~�w�.yӆ���Y���[��*HT<-.N��C�K�saQ@ol�v��Hq{]T��X5��:�J�O�_>픺�$C�㖳%�1"�'>��	h��}�s�]S9�XF��㵻�Vfk-Py�Ӕ�r`L��_hY�{O|�y�
F�N�x]�]��=�{,��)e�W�e��_;�Ϋ�\vra�"|����'!ދ�������Э.�⎋I=���wA��Y�yv�쥂+_+� �'>�Yh^J�5��_6� �\l�����oYF�]�Z�>����ۭ�S�V�h�T�d�6V���K�Ʉt+b<):�y���u��{�.��\dJ�e�']׊Q��R���e��mnRp^Y��(���a����mh�����q0�͝·y���E�0n�ҳM��MP$.�=ѓ7M��T�9���M$�Oy��;��}1w0��7\W5u�����-%��ۍ��ٙgy�GH�?t�NR�K��"���oW¶��t�!e��n�˃�L�V�Ң ,�x�j�����yB�pD%Mx�4�0��/9I��mj��+���<E	���ń#X��R3v�(<i���s0M�}_ku�Ւ��l`�q�{�R����r�Y���dm�b�U��W��X\�2]q�ЩL�Qk�Ia���S���0E1�Kj���(�D�u.R��Xe.�%�r���>��_7]�9W� �):T�D���yCM'��`�ZU�F���B���J�u�G��i��� �]11���-�&�}�:�)���(�ܙ���1��P�b����l2��#��[���B���3����t��t�yvM����I*�)\����	�ػ=D���Q��B��:�zVmϕoCw+��Ew�PIV1%*�Vs���-�VV��dp�dRӴ����N���/��*�q�f[�]����uk@�,N�qZ���#ӻ�D����S}C	1���o�蓕��&;�����Y��Vh��`&OC{ϫ���&��)b����������㣗�v(ep�.˛�ġL��or�Q��9,v���i��ʳ�[�W�؊��<���ߴ쑮7J��
T��k0o�6].��E�ѡ�tUg,���ƴͣ'e�V0��4uBÓ�����iv���kk�>������S!a��j�ô��n-}�^�l��kh.��&`Pٽ�&���g1��,��A7)����f:���|�tKr9�7��:�ʵ��9��(_|�_$�DJT��DRL�IAM�DIQED�0T�EDTDRL�QT�L�UUQDT1UM1344T�TMDTUQIECM3Q%UQDTDQTT�E$�TUM�QUUTQUD�DLE%2DUU��CD�E&a�U�U1RQEATTUEE5154D4PDUQDP�QUQ,TIE4TEM4QMTS�DUUQE�UCED��TT�MTUMHQAUUD�QKIQQD�LKL�PLTT�LU4FYE4E1PDSQ-5D�QE�EUADMS@��AKܕ��kV$YD�]>���IC������:)nK��`C�hZ�S��nFen��}3�M7��!��M�z�w]��U���p�Aݨ��d���Z�������U{\���yK���'bkϟ��}��مY[��;/�=��j��5�;~,��:���[�q���/���R&'�����3y�#���ݥ�;�q�>�Y����t�,^	�
z}G�A�C�F� �~�_N˷�1�>�ٯOUc�c/�t�X.�3��ڸ��u��FvT����P�b몽%wQ��KN��SX�5^\54;��xoG��}�~<�=t���1P�*Q���<?)[y��'s�MM]{�-�rU��bvg����*'��!����	���{��u��Ǹ���W�(�	�-t���n�Zu�ν���P�1쮯2�]��߯�qW�~ӑ�'�{7���{UH�������P<��;t��zGz�z����������o�ƣ����>��'<{M�}8){^�xTWH���O���FyM34�Ae@�� �:�t�7C�F�|���語���O�r�.w<�ǔ�3���}�TN���dT9���A��㤌�����'Kǩ���B��n�z	��.U�/з��!��W��E#u^�2SBן��@j��|=z#ׯ����pS��3�b������s��u��<j��ɐ��BJ
 ꂋ�i� �y��C���T��޷0�v���n�g�0wl��%�hH⋸�5�x��a�h�s�����c#��g�=3�%�F��n�Qd��&az�Oa���;���a�×�J���T}NW�o>j�=q����]�mω���b��؇���{&0{�iG����q˽�쨩��t�l�z�����m�c�x�@zn��q�@yV*�f��5��xsS]��<�����.��gg��[��e��;�)|o:��'�8� 9��O2|VZZ���v㐳w�9��D�C���ٜ��|
5��a\�Ⲽ6�S�x����o:�Ǯ��U(��g��{�j�\��O��{߫4�?��7����χ��i����m����:g���}��'
�>�/S�c���<׫|S������1Q��h�wo�0�O�b�v��e�*�5�x���W��Ҡ���1����]�`���������geN��,�|�������lO�ý]܋�G�UG]'w&�Py��]�x7޲.1�����Lyg���쉺�[����8��A�g�w�Q'MI��*��WMzOQbYz�F�^���Ѿ�~R�z�!6��ģN��_�iSDk��
�b�n"�u��[���!k�t�fIM��pG���c:Z��c�n_�{M^�>0�g�{\/K���u>��H�.t�=ԕM!�t�s��t��}(N�9�WE������Y�=��6J�m�t�lBD�5X��ϴ#R���l���ٖ��s�-ς�wG���[N�ƭ@�ފ��V�ڜ�x��;��������.��<�`XR�f�t�Xϟ]o�ل�Q�F��:S������>b�����羧��N�{�o�U3�%�P@J����-����>��7~6w���oo��{A��}�A�:a�s�ý��%G�����ꉦd�H�߱{�_k�����W,���I�O�u���}��F����ߕ!�O���%�Ӏw��=�����ݫ�G��g�\T�Ƃ�*��!�I>�tn)KG��~7��G_ɫ����Hg���z��L��L��d�=w��֧+ܑ����])3J|O
�̶l��_N���^=g!)|m�mǳ�y�����S>�n���S>k��3�D��R��˱|}�&�S���KcӁ��+N�����{������@xK���Z��o������>��;��^���3g~��U@Ɇ�mhwS�:'*�]�fa�fG�bO��%%<�U�=���ϵ������k
^ʜ:���~���fW�o� ���ފ�+�76J3Y�c#	�gx��;��"ss�/W��X���zJ��ZW��{	Ω�b���53DDު�pG����^��&*z1�R�qn�#��S�p��|�4��{F�nV�˒���8#*��D -s�����[����ڊ�Z���s��3�U��gޞ�^SC4��=�#`]j}d� �ܓ<����N�3����
�*��/ĮL��\�g���=u�W���vo
��>��{3��V{]>�����|6�^zadWz�M�\�gO����p��ulO�]\�=#�c��p�}n�{=��}Ӓt?L�K�����~J��~ayz~L{�m��D*�wƢ�'6���_�>�tQ��x�z�ǖA��_#�e�rA�X�bzUO���3�����������+�X���Ç�����,���{���Ê%GĕPe�}RdFg�}X���%FR��5���dz��N{��}~�g
���dy�y��G�*����t���ͯix"}�vg�ɢ�_��S����;�d����f�Q��Wq���1�ב���߽$d℻�o�X3>7�"j�.�t�zD�=2zj!���rAnx���0�5��Tm�7�l�ޙ�>��,�'�E\N�!��������3P�Ih����zH������M�~.#܅GJ1~�W���k�����:s.��3�m,�Y��>��ݶ����8�v
@g.�X���V�.D��[��ã��W+��8+V��eT�>�]o���S��ȁ�fL�����i����!�| �7���	㌼](U�]$ީ7��it*�%!vg%t��O���Y����f�
snfED"�M�^�
�T���V��>�3Ld��S��/;�BΉ{Gy�>��	'FO�ޟ@�d3Q���2M|�'�d��>�ar�5WwSG����^��!��{��oSm]�c>��w"��zf��|���h��ɐw�Ī�����쾿A�lcZ�}�'Y��;�b��>[�Çm]xw�u^G>}�9��'f��q����⨳o��T�y���(N��7Uz<���/i:r�T�η~f}�e?T/9Rޘ�6�6��$�Y�U�މ~�[�䜸�`����N�93�b�W�GˁP����hw���nv��;@�w���=��>���{";�U;��1������h�D��UY2�d�Yᆝ9�ow�=���VFov��r���t���Լ|z���;W����ʝ4>\e��x�n1����+c�ذt�G^���r}j�>�ޫ��z=>��~+=t��|f��D.ʔn�$���㡸�"�]��G��Uʽ����J�J�Y��o,C���џ{���s�u����iS��8TB�:�;8&9����W��������0g�߄�m/�����W`D�nA�.@���o"߅{h%ݑ�����7��80��,�-Mt��pcc�Ѥ�*�Q�c
ʈ�YvmT���A��I��D�<�3Y�:	[��pdy������$hDD��eL��˙��� ��z���u6[ꨟ��\U�z��N}�'�{"7���>��d�RK���}^�54�CIH]2��%� jvK`7^8�Z��cQ�~Wq���iydR��z� UCq,J�����r��\g�dmǦ��H,���Q-�_��9�I�9N�D����o��K�)����l�zw���{I�{���d�"L7���������7מy>�\��.Fi�)�{ܬ���W��}���zg|Kϼj6;uP���&a{�����[9�V�~}�=�`�=GՒ�M�TǼ����܋m׉�x��f� ��w,��{W �_��/Q;�E�e�A�ÿV�g�#z��k�^�uto�~�=7��8�������ȆjRQx��fg�y�T�P咪����
��V�/���R��g^\,O�|\� R�B��Pz�x�bе
�J�.ʉ�or����g.:|
5rXW�������ۊT��9��k�C�tu��v���g�t��1�?R�~UQ<��Y�����|vv����6t;��:4�A���T��ZE)Gv���T�j� ��O<�
��x??rV/�w�^����iK�_F�m�(ca1���"5v��-AJa�}v�S�Kd������3�wAgWT,r)��_+Yve�u��(!�����.�k�v��s���F�T�B챩r�&�'^�����%��x�V��~��Y�3�3�Nb�0�%j	���sX�^���{�'G���"z@� ��N׌�v�~=u�u(n�y<+;*t��@�'�o=<j�E*k�w������3ꎞURw����؇�Q�z{~�e1��<6U�+�Q�9�Ώ0���޶��{����
��<v"O���ʨw]5�7�,K/�T5�^Ӟ�>>�"+���}O��PM�t���}�_�ÍO��)	=�,	�yT;��n|)ԟ��X�˳R�mx���\�BRQ�q>:�ڮl�
)Aʠ�~
W���l�|�c}������b�ண��[���ߩ
s�C|�z�;���*�=냷�a��B�T}D^ν�31H�b�Ky�l��=;�;�΅p�ւ>�3�Nu�v�{Ը�����~�TK��!9���Q���{�J����K&&'�]F륢�b��o���;c�҉�x�d��ՠz8W���vj�e�x�Ը�Gޙɗ ��8��/��n��z����К�I�{ԁ������ԫ?{���)o�n$BC�˪ӫ���|슓��\�rCtS�&7p�;q�Fṭ%�,f�ҰŮS�w��NVӻ&�.��s��P�0�r���1��}+���j���c�]��n�TK�M7:���%��è�et<%��}v��Q)��];^ SΜ;3��&@��o�)����3/�#c%�h���^=g�����x�gT*��]p�N�.�g�[&Jn@��.�\��0ʑ������ꕧE�Z��.�}BPW�� ݈��7�o,nj�}���~~��_��'�|'_�(������ށ�\��p�"�P��vkV{͖=^u�{zP��:��B�{�3_�/K�*�+fČ^ʜ7���\���Ʃ��~���G�s�^O
Zx�4��.�-�*#s��1�z��߽�^/<������ї��3���j�>��	�_�W��wA���*�qYU�I~%FK /�7쑑NW�'�1oe�W{�s}����'�ϛ�����<�ㅑ�ר�1b�Y?$B�.��=>���Nu���]G��߷����*H;GW���~+#֮7�=��Ft�nI<J�<�uW�b��	sDk�QĪjfW�R�ڭ�����z��O����~+=n�ݑo�|�a�i���|��L�6��Q����ط��Β�NE�QF�~�mz�8dyS���ǻߌ;%GĔ0�uU K��E�\U�����	���kkPWeJU5-��v�y]�o��oc5����N�p��X���뺟l�}�ȾV6Cqč�E9(�5l)m�-��*�X��4�ٵ�K�`j7r�|��KER��l.�aʈc�ޓ���X��a���������ne�8��'ޯ_
���g�}^elyQҮ=���N��T*�?<�羵e��gpu~2}�"U��u���^/v!��F�}�qW�,C�yߟ�'*s�`L�9U�n��_�K��/|ꐔI��" ���H�n�-n�Q��Bc9�[d8p�{!_Q�e�s�s3���=ՠ�y���2KDIl�$��SҸ���2�^I����p�B�<����F�_��"|\Nx�d3XC�s2)zA0��V�x��g��ϫ�����I.�e��=��^�=q�+�1m�Y��@�&j2�}�I�E��2a��P�J7>������ף"�Ը�F�1��Wx�O�r1�G�S��	�^�.;�R��봽�%s�W.�A�����~�9������;�Q��v�xh�m��b�W��}�4��btϱ����)i�_�s98�pJ�E�K'h�P����2K�p�/��[�uU�s7~UM\c3����92zߩ�wp�ֱ��ő�>N�xf �t;�������(��e�߾���߶�z����j��9�p�o�>A�����l[! j��b��+��]�$�G"�:�b�k/���n�c��ʳ})񺜀d2�rm����Nv�:ڵ��KO5[�:��=�EtĞ٘�$�U�Mq"3Aݎ�]�y�v�լ�-t�+c�����]8�!�~��c�9^���~w�VB����uߑӷIxc	A�N?�`�������a���7ԔU1n}���p7��m:^>=t�{!ڸ�sh�FvT鸋,�+2�D�ݷs�W�2�:���!��(NL�������U��7��E����܏z�����@���R��/n) �g����Ic�L���]p��S�腙Q-Ӻ�/z�dG�O�w#�D{��c�r�0<�k;ElY����l/|.OGğQ�p��ϫ��-w�~�u�\G�ߴ真9�f.vx>�T�E�=�Ϲ�����u^�%R����X�n����}41���WO@������"�,������;�r4��=�#o�L�C��PB*�'�Anx��X�1F��٧詪�3d�r�3��G��ٌ��_��>��o�������E9��٩��uJ�ۯ9�ƾ ]�n�^�Y�Jh{�J��x8�+#��_�����sĵ5����R�O�]4��<��ݻS���:���js��<^�>�u���G���!���3���~�ݝW�APE�A��A�TWT_�A��*����"��
�+��*�� �"�����TW�WT^�W� �"��
�+�T_����*��APE|APE��d�Mf[\���~�Ad����v@�����o|<J��� ("(H��(T�&�))P�j�`���H��PPE	 Z      ( J  e���i ��4�mm[cm	(�2�]�J�����*��2��  D  ���P��مZ$��C�N(�����mPA	Q� ��. rt�l�!�ke�lS!e��@2 %"JW`�  � @� [ f�@5�b�� �R�P ��P��H [����@2��h���� �25f���,�Ռ�DQZ�DUT�cU6���T$�kf�iD����܀�-� ض�e�Ԅ���!��(.1�`�hhkfҫLT$�-��*�ˀ     Sc*�R�  h   )႔��6�F   4�ɓF�� �0F`��R�M=B`20�M4��4�ɓF�� �0F`��IM h$��524Ѧ�43A�|~r��u�}?F�������k�����}Z��a����(
(�Ђ")�M��?�diDSuKo~�������?��v����!I��M�U$��N�Sԉ��6��%PN!>Ï�=o����}�o��{T��/�uƴ�!�1�c��������~t�>��}&�׫��N2��ϻ�?֜9���޵�д�0�8�#��K�7/n�ȢN#k�kk���̬U멌�ck6�M��v¼ݹ��*�u-Yb� �XnP�{T��Kwe���%m��lKz�6�A	�7�ge��ZWv7]�)+c���?#}I�	��G2c����hm!ś�?j�6�Y�����[���)0R[�-xlP#kH�Ʈ�6;ZL�9wΈ[�e1���2釪�ۆ���F]R;z��"F��e��������zE�7{E��!��*�OwU����ulu���Yb�*,����P�ȑ�h�fɛ��3�n��B�s,U�1����gr�Q�&�f��j���2�	�Z�t��-�JۂK��P�@�;���mV�ҩ�Y#��aԁ�}wB�@he!g0�����hw�m�<��N�U�|~���f��6V��(���1��F�7�od�2�����r�7����l�&��f�+��7-�b�a����Y���3hޑ*�%�8��x�j�ٷ��l�-DhL2��Xvޱ�h�B�.V:�Ҟ�6�JRʣ�Q�h��m�9�Y �l����eF����O4*)uݫ�Z(��uok�!\G
/�O��Th��h�H��Y�*�ܚ�5%�����;#��B��Q�0�N�*.�rݤ�Wf�,H:4�PӜٱ��Y��bܽ�Z���0e-����;�
�Z�uq���ќ��ݱ�}a���zX�#�ζsQ�o7�c�ػ۫o�s�h+t~Zr��,�U6��T��j�%Ș��$[w[�гe��W��X�����օc�O�2�c�z8x�����RԂy�e���n61&1c V>�A!���Ž���ն�*
�@�˕N��vMۣ�\��FI�vExeb�snb&��Q���qԫ�3`5m���[1ŵhc��R9�#H�PDӫ�]�C5��1��b:
W���pl��͛���L@ࢶE�,��U�.���S�D9���ql9BV��N"R�����Uk2Vl0�����KlT	9�(�3M�S��|{��z�`��a�����/+��koD1I���N��'u�(Q��a��٦M�m� Vr&���"���WVX�Vd�ﺱ��b�+ hX)O_^�;��G��xsM�4���&xqV�)�JA�ƙX�GI��$�;��0f�l�.�b�	��Y��0�8���H�SK	L�u�ۆ�S�PVA{oʫla��{�&SS�)em})u��T������mG�H�.e]�̬�+빆"��7FT�F��|�[6f����:��^��t;y��ᤖ�g$����G �Q��e��fR�r�1K0�R���~�C�h{wZsKQ,�����@��bS;pV<����C2�T[SM5-]���7��g!݆�6��l(#�vEDI����a�y�
��oX�\�46~ʺ�V[F����KM�x��͠�*ĭ��O�݌#*�ww�+��iK�쑍5�9��q�(���1���i�18�-���0�b�I�M�RA�J4J�T��������m:0����)]�ż��+��yb�]�v�s*�R;b ��n�~ŌZ*�ƓŠ �"��l�:��5���&�06V�2�EA���U�˼�yu�:�V�6�{�Z����Ueɴl��2_�y�� ��f1*�����uk�@5�3�z{t�汫�o*73D9m��]��$ӏ`.��U&]mr���6H�k.�)�O%�eUA�X��[��yP:�YƮ�����|Y8��qົ�T��V0�-d��[Q�_� n�Y0�#q�/MG5sfmh̬ݗ�T�|���p�A�(;�{x2�ˠ����i4�!���wC�����W��יz�;�E+:Q+o6����=t񅏨��_$q^�����v�â���Z�ӸWϴe�XN�W7h+���V��Z�L)�ͽ��hũ�bh�K���R��3뻕��.�V���acj�	�ФC6�R�SK��L.�;P��[�K�ٻ���Ls~��D*e�w|������}��v����o�ҫk2�z�6�%|�����ua�h��4�f���إ��nQ���ђ�]��K�1Е'���{5���8��^\�t�����T>�uL�tT��a�����.I[��a�����Y�Cv�[��V�є���~E�45d��4&����0��Ttmݥ�\à��&����ęZ(��i�����rb��z)��t�������YVi�cMxI����^1�q�f���S�U���!X�vE�%;sj$�޷WA�U:�H��(�ɩu��.^#(�XqfK3ܗB�7K*����)���~.�!F��ꭆ٧��)�	n�M:�,��b^����UnY�G���_u�lUƏ����_øQ�D<�y��x��@�8V%�K9(�#^�����&nR�B�rK�%�G��J�D��[ګ�V�Բr'wL���t��m�	M��J�f'N����v��P��x�5ٹ�tF�u�k\�g]��'�?�l����6���֜9HgO���{k^�Q�'�n0�V��ޯ�B��?���:ZLHf�<�LHB�7Y�1D��+��̵}NfZvK�$nHQ����b����%i���ҙ�.

&�&��B�8^�S�gܴ��٢0	�o9|��ˍ�,��.�ty�ϕ'3��`Y�Nfú��.ƹïG���<���BEH���=�����rf���N�m�d�8GU��7�5P�a�� ��y�Wgxi=Zc٤c�V9y*Q�$�tt��"�h,��F�'\�R�ɢ&*^%�Vq�]W}EK"������X�>Κ{i*�6�j��Wܙ�<'<���+��fpJ�,�HY|�gcɀ��c-���n5��\�	��e�����[e?��]��Q4�A�(�� ��(�Qn���!�n.�y�U�f�T'wÓJ0Խ�C1S"�]ai�Î��Eu0�.V��dÍ.N�d�KSrƶ�қN�r���&��9��ԤC@�3��6�����J��r��&⫴o �ھ`i̜��p�{.�����6a�:] 5��`6`ݻ�N�"�S�vu׭��N��r�D]B�T��Q��vN���x�7�b����r߼�=�6�On�6��V���v���S�ɖ	�<��l�\���b4k>�=ǖ"sv���ܥh�l����vH4�.�&�����;��&F&|���D�ޣ��z�{�L���2V�^��(�C���q�����wJ�+1Wݒa�����=�����w5x�]��~cH��W���f����˝��>�6L
�(����"�Jr���Ԭ|*f��55��d�
��XZ�q����SR��>.�-�ä�
�7�X���{���|C�V�+\�MuQ��  AX��7�S�hvf�k�^��,wt;37���e�9�Wf��y<��̳{,7�����4k]n�dJ����S{\!�i���MF\�]5��U1���j��Q�Iug�η]��s��7�a&������ں����a�I*�y5�K�B���8���)}eLm�|���(�+$�nѠP�������ӳg��3�t�^�y=<��*ڧf#�<��Ca�g*r86�p%�'�[���i��ڼOif^e���@�#X$N��C�8z�3��Z�؟\��2Έ���^���2^���T�Nޑ�V4+��\�b��i�k]�蹼c�+uk��w�G�ˬظq��R�Q�3��s��}���=S�ח�����d�4+�)��s����zfI�����2��R|N�1	���<i�Z5��Y���f�wo��ֶ���"T�.��Nv-�Gp��ܸe���`��r*�M˚W��MTQ7�қXs����`R=���)`�\��ge�^��/f�y�"�W�Н��w:\�e�F��12f���]�E!x���PydU���:���4`��l�إ֜���`�9a(-G�:�n�-�]�����j����$W9e��[�˗��{�ڛ����B�{���-3�il�Maq���m)`�xe'�86�5�kJ��D:����Don����t�vl#R�0��fup���&��F2�$:������ꁫ��ӭ{6���CS�n��$�u;�ر���}X��-=_7ב�����7M�Wz�e����A-��ݭB���b
N��|���<��n
����)��v1�Gk�Z�eK؃�Q�
��%�Ïq����׀�b,�a𦳪�dK:�sۚ��Q�"GG��Je���}���W'$�W��x�XKXǕ��J��%�2Ų�چ��u��y�x��s�/�M��.��0@����Q;��hVi�9�썭�6�rlq�Ǳ��J�ڥ��$�5ý@�8�̺�;pL����C��dnK��G$�I$�I$�I$�����܉�����"R���۰
�\�#m�z5vm?�uN�R}�oL�΢oT�]�1���2,�m����"�d`��3����0���%�����Zi���Zb��\�ұf���Ø����UF	vْ��dd���d�I�;�6�G�Q��vg4�#����7z��$�m٤����*bi�ha��.���UT�����[uu�Ӓ!wFԇ��N���+.�>�O���M��$*m1�	��u,�z�w|GIjjN�CL����ґ\��mw�����m1���!Y@�"�S��M�@�b�]��|�$1\��j��2��k�jEb�����2��Y�WAئ���E����#:��֖�6�{wتp��YA�ƅZW�M|�r2�~G8a��/+c��#q��1K8�cC
�Ȳ�j�CH7�a���=ח{)�9�Zo�t�Zh��;څ���wU]zQ�VRtH�y�DQ��6�}�(�7f5�l҄v��wG�~ �K�k����S� bD��|R &\ݸ� C�_�����$����F�SO�x��_f餂�)��ִb�2�л\��G���TuJ'R�J;*�wL'"��A;$���<r8PCSP"�ާx�\�5E�F�����������ߞ��qǿ�t����)�d�7�{n  ���4*?P���#'�a O�����4"��?�����a��'�lڛ�,�nT]hY捜�����s�Ȣ���4C@�lSK��Xl��a$	���x��)�(���H���.�.�\Wu�SəL��	���Z�D�&,m��m��wTec�4��B���A�THe��n�1Bi�v�h6Z�(���%����w1S-���ETГ%�0�n�V�+��Ʊ圴���*��b.�pN���D:m�uB5DF!!6���_Ռ<Y��sUt6���E)q
&���P�I=r.[���k�f�r�4�L�۸�*I]�"H?�g�Q�!K����0a|۪���j��Q���8��s�R�;]��kJ0���P4��4�gE�`�L��oM�D��т�]�/#�(��J"|���(����~#]�\�s���G2f\���1�.֚�)�j��f;�03�ҷ״���m�$���X��U�\�L�f	x�m#/�E^657T����`��(�T��廫���°[��?�Y�weu�y�kc'{/6�j�#�K�z(��I�TH�U�VI5U&nC��ʴ�t���nRS,�
#�Z�WČ;V��h"��B@K '�u5�(j�M$
������pt��Q��e��i1(ݫ�]��4��l��vF~e�YP_F$1�!&��B�����$$Ebd�;j�*�?Ga�#*+8�N���h�v��l�<�Сw����o�Z�2WM�1�1"�j�l_��Dm��VD�.��C[Wؕ�M5��Xd�Q	!�䳏���=b�f�����(˻�T���bL��-c�Vd	P(N�ҮܺQC =s- ���N|�Q�����bH�G�BE�d�Z����΄�D�-�}��5iB#r�~�W��,�W�ܷ���*;Q8�*�v.�bEd�W�M�ɒ�:q�t�]�y��w�4u6���6!T"v7Cܫ�Eih�'e�q\hܺ�����:��ۗ�A���Lۜ��U���|W}�m	�.��:/���U�������AZr���]��h�E�aڤ�<�D��M(l�:�.��-uƁ��5�d몑d+E���[��w/1e���"�?M�r�C]d��ZՋ��٭6�	��*0/;\�+m�u�P*x*}��.������1�zt�ެ��!��K�K+�����?�(�kx�e=|�o�7N'�$[YM�kR�H�y�oU��i�lA\#�����]����Vô�C��H�ʵX`6��@�nQ&"<"G���řh���d�5�l3#5�G�m�G�mNtq�uLZl�I�k�\#7����A�@��8��R�>����X���,�@��a�5JP�(<mKT��	b�	G{��V�&~ �XR�d�����>�����B�0!^�<!�*+�E���A�?���@�u}K���z0�㥆N�b��M{lU���u؀8o��თ7\ү�k,/�W��ȷte�ɔGn���|�%ڃ?qr�&B��t���:`�х�\�,¬���\O)��CK��׌0w����S����,��t��.�M�/H�n�2(@iz� m����ᯛl?���kO]
k�^�eKPb�L��t�-:�5��l��v��cD�������^�<-�*tF]|��Z���6���#_ƶ�ꋍ�,8�R� I�Oj�yu�=˗K*�)�JY�R��TF�H�5$�w�B��³\"�=٪Y49��Dk��a�U�J��V�c%�x�f�l�CiaG��5`��7)�7�W5�us�?mF1S�#gH���2���.��J�&7��VZySl;�v+NG'�m�l>�.0�m|�ܿ�̓�E��$q,�Wu�v��=���&e�1`#t���V����
�Ă��Y��lh=כBQ��Ce�ȄNf4%!nͺ��&�YsL=u������@�"�#�ZR�(���%~F.b|;)f����tFZ���n��8ɦ�U`NEg
R0h�<�j<��"ٺ\B|X	>wU �p@M��_d�pB�q�G,'7Zx�Tyf/��q�(�j��"��C�Dq?��T6~���ӸU>ʕ�[�34�%�]DM6Æ��Owl������F�ւِH�+��5k ;c��M�(��b�q2t�+iZܷ�3.m�6T	�3��+�E����đ'�U6���KFiv��3P�E[�-��7gn��ցhD�\��P�B�L���|nۥ�_�NpӺ'�����AF��BE�U$�M^"���52����A�X�^�3V��.��n���sg �(�A�z~��j�Ch	�^G<�C>4��J�uf��r�Ԣq%s�e^b�V�F�FpJuH����\"�X�D�w�>AeP\ML�w93�vF_I\�)_�Ѧ�E�Kg3�k��6�U�*�����ְ;d�I��0��FI$ҹ���+��nH�|�,2�`�OS�*��o��߾��~w��ͫ�|=�ܢ�)R58C"K��Нtthp�ўQ"���q�Ǵ�K���Us����9��^C3(�;Άf_M��z��ge�-#�뷓oL�w�k���)	��V�1͚��A͔��;Nf΢q��r�O�m��(n;v82fM���	���1��_d�;8mS[	S�������AR����01�µ9{R �`��/�f�(�`c�7����wTb�7#��܅�7j�8�Bq��� 	sL���q�o����\h
>�>j�����X���I.h��6x�ꯪI�9~�y}q���I��m�54R��	��H�@U;�� m
j��R�"d���P�<��>F�\s����k�u>����:�;�*���JG��Uu�`����JX�u�YN� إ{�M�
�������
Z}�=��yU�-j��MNl�Y�@�?SW�Mz.�fR�Ln�����(�p�x�tT���J:�ɭY������	���>�)�7�w�G��c�q� �
vUbv��W��ݖ��*�#j���%�����������<�#;���cS���R�:i���&k��s��Мv0�L��va�Y�f'�bS=�>�����kP�o������!y���.��\��R�}�	`I�$ml�__G�����tȍ�a�X5�6�-��'Mc[-�����oǤ母��`�������j'�{�M6t��TS8ɭ���4�����j�G�gW#�^.��/�1+��M�Uʮ�Ԋu���NG�V�4,Z�G�.�57�S'.#��8䜐k^>��cZ�P�k�TK�:KVx{+�o"�8鵔U������n<`Ӿ��=7��6����tu�kЈ�6���3{�����Ѕӷ��6w�:]`L;��5�Lרr�w`����ӱ� :�X�K��(m׺Fs<{=okL��Qp;З��{KY�k�:#jb�ZI'�DM/�V�l$�~G�NT'��r%P��j�]Us����/y3�ݕr���#7�CK�P>��wp�����~��l�ۂ�Qx�_��=	��r�M�2Z.�嚹O-�^j���L��J⅟�K���w�n��<�v��$�8�G���[]"�%J�+oSJ3Ͻ ��zѣ%�:s�zK�^Mt���VΦ���Pװi������'� �6k�A+����N >א)B�=v#��*P�"��V�ʈ�zE�S���R�	�������M[Ȩ= � ��ֲ���74�*xYK��%i����`���Z�M�q��n�	�A+�Bom�F6BMx̺~1�R"�sk�+g�)4x�^�#�ā _K�T�[S8�&�_�T�YS�EvZ^}Y�آg��zA�p��Vp!��|�r��.����2��lqN*|����� �J.X.lg5F;jk�="���+��.\}��X�7h��K����)1v)E�(��Ɔ�m������ה*��gWiݐ���q{���ʤ�b��0��m�#�L��M�I�7�A�K�,��=�IYY�����t�VvߕXx�o�ɫ˂�,O�ۆ��=�Z�l��3d�VC@(��]ǡ��p.�nB��}�hK��;��W:ȳȵw�-sQ��J[�22NlL�Z�>�s�®��T6�a|w��!���;7en��%��ܪi:z��5��)� .�ۏ����^���9uyWy�d��P�+-�����ᒣ��\��M�wz2���_5"�J���˲�z�o{�:�aV'W�cP7���X�u�8���I�����ry�����t!��d^@V�Q�w�R��[�p�6\�h�ֻ������S:��su�6�mC5���+��<VT�	g�D��L]K�tQcm��ۉ
������f:|@�D܍�s����)�
�|9��\7�>���v2k}�Vj���(9�[�F��g�;��v����R�)H�f�Ts����%�h���M{����G^˹��ɴ�Ư�ڷ3.Ck����g�LXN��S}��jw���DҗSsx�س�;yƍl���M���/�����y��zA]����~�]\�x���,�Q�t�����O8�G��&WCZ��T�_rii=������&����W,���ܛ=m�X���(�t��X���_� �m�h��5h=�pI��T6�u�kz4u��.�k�e��gh��l�/tO�Y�%�t�x������Ɛe��?F|��/��T��|n�����w��ٴ0O���r�{�K��R��ۗ��JZ�[����rJ�EG���Wg���X(3]�����o�ZCH\��J+Mq�*��\o=SZ҃1�{y����W0o(���`T�T-�Ly9�m������zb���v��-{��nj���Qپ	�]�zw���=�*�;z�@@{�Hw�rs��s�cN�{�1�(؄�q���2���f�$��섌����1C��n��w�D����o������q��q����pz��n9�<�8ދ\����d�n�5	\t*�sؗ-�ns�>��]50:��V\�����K�� '5��²Ӎ��o*V�EV�:ia�{:�LN���i���6���te��r�:�T��[�uj:�V�{j���r�/&�MR�v�`Р�X���vN��%��;����<�m"RK�$iÖ/�m���:�h�3��L�	��׵����`̢g\�C�N�ǯ0��-k��+,��3n؛�V>WM;�QE˻��NIr7mPK�u�Kt�o�T���v�Ax$ ��+$?�-lu��юt�XԸ��V5�Lo�rfr�{҇P-�ۼ;UA��NNOU��}�ݸ�k���2����"P!���s�f���p�03�OA��)�\lk3�x]c�D��7Y9��p�X���y	�Eƥ_C�n�3ld��(�!�ۏP�±>rR� FcD���Dɲ9#�ݹ���\ӏ4pQdz6B��G�Ut��!1��Ȅt�����<��/	���V�F:�CvgN�p�s����>T��;�ը2W!ȥ5 �F�������"d�)�R����&BR�L%�i�"T��vNy��ף]��{�9]j�.�!��]��'<�'=V.���B���{���P)�&9���:�#��X�?&��Q����֗����S~yl�Y�,�զ���:�2��4}�
M��-�m
�����Ɨ��p��3}���X�W�{��yz�$T��\X���lGTM���/CI�Z!T�ø9rk!+���'���I9�� �����3��Hf���驃]����n���_��zӤ����]\�N)3�0�y�ڂ+X�a����v�gGh�:�K:������稍�.mq7�0A��z�H����il�^�Cx��S~x�u�`瞂�EsiH��^�n�?7�4�=�!�"��p2�dY[���5<W�`OQD��kZS��硔��������#3rk�=Y&W���&�%s�yF��#���Gv��AŎ� ����ã�;f
�z[�s�ΙӮ��-5ȹ���{��VSJ�y��Go2k>�������ڛ;��x��z8��ٜ8r�CB��.�䞗R�ϊ�/��u������'}Κ�/�t_�/w��2E��ub~���h^4���&<�̆����y���h����}1����x�X&�2�Iӷg���Bd��6߄\��(o��.^dʹR�����t?W����m��׫S�G���F���n`#��0��:e�Kں�������e�c��T,�|�=���*Fyn�;�!��uFT�i��c�D7C�7��uDdB����Ꚑ��Z!c�9^���M�oi�|?(Wyy���%3�2�rz�~w�<���:�(5�"Q�z��C0O$u�	Cܺ!K��^���;�[s�\�m'�;C�������sRGz�5���B�;�9��ε��<��Α��8��u�
j:���1N�:��� �T�:��z���z��<97�f]o߭���;�ؑ���}~W�e�o��~�i�U�
�u���Ze!G���Iu�����6�M�y�&�:�!G�]����s��ԮӶ�z�=wߙ��ͽy�hq.�/P�Hd>���xB�R�q��S�z��)��&�����o���u�@s#�q�ʺ��e7�B���ex��C~�ͯ<۽��~8��$(��;���8�8;�z�ԻJ�(�<@����W�=F�q�fs�z��N �B���MJo/�:��\�k�(��;H�z�m�n��_#��u+ݶ�;�5�)�������/>`R�Na��<�6��� �SyCԆ�/�;�L�p�lfP���S<ΡJC�k:�6�q�^�QԾJ��	ġ��<HP'1Ϭ�v�;�9���G}��7�=tm"s��z��:���]�)�Syz����J���]k~��w�~Ȝya�G�$2�N���B��N!^��8%O�on'��{uW��7�jF�����8N��G��[%h�����֥Y}s��=f�y^�ũz��D�*1���ꇉ����u]|P;BI�^�z��9���N�۬ �T��]�:��=���3c��o�K������R����d���M�N�=Hy�X%p�r�ͷ;�6�5��;��:���Sh;�6:�6��7�<��z���� O$;���;6���]o�0�2��"s ��x�Gx}q�jSh]Aܝʝko5�s�wٴ�)���w� u.y�'2�B�F�`���&Bs���s�ל���[��jAġ�6�P'�@z��z��!}@�+�dm�*[��m�z瞓P��<��[�<C�d�C��D��8�5
s+̆��Q�}Hx�;��=v	N��uy�[➤)������PH��w��#9�n����a�y#���@��}B�'2��y������|�8�3�W�to����랕:�Ԧ���;��P�"oq�'����;���:�������w��Nτ.:�;���������*쮩&���<ۺ�M;��d���H�����9�/�U���>yUU��^�!]�8�=@;C�w.@fP��J����]�����j��J�z�<��#��"�)įPq"����}�S��~�����i��I꾟��гO�WtR��Oi�9��٨�������s�c)n�������T����CM����V�Zpp��vC���sE�#Uu5tP�ăo�q�B�5t%���Ⱥ#ץ��Q�~����+���̢R�W_�nS�?>�j��|��{1�1?%�t�B��<���)�f/꾪=����x��/�޺a�8/ݡ���C�$U��\����`�]���f�¯o+��|�F��x���
��0�>�I���{�KB0��,����ⶍx����&x��1#��p0a�ˉkYTz�
��u��s�)2�w����E!��5��M5_��jڂǺ����#V�0��b��x�a��%�Ï��H-k�tpU��Sb\��_W�|�O���	b�=���ϫH���{��H$*çY[�EMRkK��+�9�Y�njK��Tg�:l�����y-ٌ����􏊤�;u�{/�{�Y��cRZRf���X�^v(�� }9��0���뗜tu����˰��k�'�z�\���2���o-�8u�M��Oo�7��������/�B��͇0�������^��5�	��V���}s/�_}�|wdj���x�k~S(w��O���' ��f�%�m�o�����-z��"����G�%H��.VMA�<v�=���غ�b]gtK;��tT��dk�xO`�c�uY��3Ge���R���/Tݭ��Zr��Y}������]���7�"�����2O� �����C��c�����̓�:��]`#�z��a�+9��m;e�uwnw2�#�c��F=ҕ���(�+̾a��9)$j!*�DV�0�m�7\Fnf;�)�,	�{)]e�b�PHj���+y�9��⮭�4�q����"F�X��Q�w���q������佛�M	;�S���9�j{2������RN�śtZ���ݣ��v݁S���9�u�f1����V2��x4�KV��
j�T*�,�37�W
�u��������+V�!O���/ȕ�ͻ��������7nv��-8�Ptn(�p:�Ϥ�Z������d��(���W��'ei|�:v��CV��Oe��wz����3vݬ-���ouY����t�P�-��P���啧U�m��E���I�3:�.�>���%�1e��:m>,���oϭ�%-�wE��%�sJ[�-�D��O�I��8v�AWG��ww7z�)��4 ȧ��@t gV����� ��wV�(L�jƉ1��3�[mmǳ���>��
N npMAF����u&KER��d��թ,�' C�QA�0��i��	�P�Y��u&AKY�Sf�j�Օ(�M�P��\̠JMZ�)ԁ�E�P��$5�DS@PY�����"*�)�S�'{qy@�?��y�I=�/���3�4���-��#��_}_Ugj���C�v���`̮�O������oح�J��Ɣ��n��k]�e�fq��615�!E3�3O�����cN"g:SV�7���gܦ�BO�\�r���6D�X�G�����щ��~ڻ�*�P�jѾ2���ao�V9pԝ�Jd��Б��yy�M�]}\뗷�y�,���������<��f�Y���
��=I�ͼmZ��3�Ɵ%/v�X\��ꯪ��3����W���ާe���Wd�r�o�}eYW��KP�پ���l}�����Xdtav�w7���:���|]�U��(]znWtr�u����eO���#^���07&{,�����٢]�w9�2�Q�	<>t7L���������3t)osuC��0\�ۦ�i"��U���lS6��X������>pS�K6��Ӝ�cXQfH�_W�UU����?��˯�߯�Y�~��Y�N�sEOx{�52B�C2�Oo��=z�bm|��[hexE�i�,���>���g���/'9�͒��lQ�U�H�����k��0l��:������b�{˵ҁ��s�zK���˱�U:��	�X.��,�`�]K9���g�B09uF�l�d�#��2�<Y���9����aXOL�k������^��45>�����睊`ѝ�?=�7���F��}�������#00�ޗ�<(K}8xmp60\�H������o����e��c��ϗ�Dv�z��nI.�>$�,efc�lz)��,kU�R¥w�xJٕ��z������)�v�P6�˺�ظ��b'���N���lY��T}	�y�<7�k��.�g�������h�t�o_i���,�v�X�kd�(�������JO�g�Um�ǿ�������&�.->���s���zss4s~���]z�!��3 +�΁���nV^�\}�� /WY����7׊EC\�"�1Xج����_1�w���{q_��-���W���ꈝ�l\�Dm�ecOw�.��0r��n{kޡ4�}g��.�w-��Io�ĕ^�<U��=�t��3ޓ4ӭ7B�rh��rM���}�W�,	����acG>�d�߅ LJG�e^Z�}�s�ި.���2�u_'��Ҩ���[�:�4�{�����::��߲��
���єh�3���,:�:�
({�<�����X�Kb�Qvm]�H'_��/|���Yyh��hrW��w�39���S�g�3���9�w����<䦀��&�h�m�m	�V�.��eJ�I�s������퍯���k�b��3�=�#+�6e�Ό�P��������{��bG/�̩�KȌ	'�uz;��x�\"�n����?/.���5�� .�{r���rJ�Kv��yvi`ƛ�i��=/��*�C)?s9���_F���(a��<'��i�R�=U���:ev��c{�^�U�:�d���y[NR�K���3�r9�>A�$�Fv*܆�����9?}U_}\���Y�Z��!2:����R�V߳����YIMso�oh��&f�g��P�6��{�>�죑v6
����������]ڋ���q_�X�O_�_�L�K��ʳW�>�{����%˺���x�}ݞ�P*%9�˔+5��(v_�[�.ܞv�eQ Q��۳o}�u������Q۔H�
���p�M�R��A]�$oOJ&��49�P����U�|W��q���k[I��ժ����:]4�S՞�x��7��KL:mP�u�Sױ~�%�H.�y������#��J#eC�o��7�Mﻟ��S�ui�&>v�^������;�;�_N�[��=��C��MJj}"VT5�΋^�:�������qI�nYp%]�kƓ����S}fT����+�V�y�f��DzK���_,����49���ׁ��V�5�fxţsh��9L��<���S�ߚ��$���C|^�Ϻ�E��"�y����E��q�����.�gi�1'sӃ\�r��Vݳ��U�s��=�
l��^�kܢ�ͣ��U�l�]e_����-����u��Y^����_����T'��k;�۵��� ���Z��6�}(p�F�c��A8bm(���}��8�!�ErR��3�bՉ��Vv��e^A�k��2�4�oj�\Oq@�p��Y�-�f9�=�6KwTR��	]D�r�Ǔ�B��ǆl&�)%�/�^��b1;��Ƈ�����o�pA�rBj�m��Z�	%6N�i���ego)�6ue�yR�'3��"��`y�t��v�sܬ�z��q0W'����uNs���y��EJlɡ���t����l�J|����C7�]nι��I[a�IK0�������ИOl�c�;{���җjIiSM�G"K���v��=#�m���Wŵf�3�����dV��cy¥4o�I�;�WS;	�̓vHV�ν��)�W�s�,���_��m�g�������IݱI�Hp��Rc|;qC���7�oC���ʋ��8k�e�r!.P@�o�B\!Ir)#k@�z\9�I-:
L�w��fY:o
��I�EȆZ ���-F�2H������G$���a?|	 ��� L�i���r��AZ��d�dd�d�T���P���eNCYkY��H�
"��ȣ32����!���%�d�df8�	��I�fX�Y1&f:�U	Z��խ`�Y���FZ�V��ʀ�Y����NT�DA�cU&�Z��ce�3FI��'#"��r�*�ƃ"�#,��2���&��k-fY9��d�6c�FX兑�QP�'���yv��yҍg;�vS�V%���}U��|�_��Ԑ��#g��^���֑������J�Y�]��=>�j�F�sZl����{L��~}�M�!�!W�u ~pnyƻ��A�MX�۞������}~��,�|Bu�TW}��H�`��j{�*T�[�6Ы��=Z�ʍo�[��v�Ϸ���,L�д�}7/8��sm�G�<��=LFٗ�7|���O�b���I�D�U�ù/>?��k��ߗ~���q{��k�N�Q��C7�.�9 ��ڮ҆��c���56(�Wl�7�J{�W��ek��V�h/��/�١����:�0�ҡ#׹auꬼ�N�NlmJ>�=+�����:�q�Qy��&m�{�J��
�����)i�z��Ļ��M����u۰b��-c����;ُg5��]�G)5Ԓ�W�UWФ�6w������%���%w�`3FK}��7�Lu�m�m.����=l�7<׺Re$���T����C�~�29�֮�Gf�]�n�mgNV��~L_f?4��l_ԅ\�L�N����Ƚ�^�.�X��bz"烔=��7Yo1z������*	�\��_j_]Pw�;�v}����i�6��B��7�yPK��j���]���Z�S<q��cs������z�n�u��}�S�#de�t�־��^�����3s��O?p^;!zτ��9���Wr"��&���ꝕ���h�R��\��N��z�.Be��g�ע.����̜D:%�Em��C�D����8�g���>�f��5�+��Z!�^�B�ِ�0ڞ����y4\?9�yա��Z*���Ε:������1J�t��+�����!��/e;6���;�N?p��o���z pE�{�2�{��
PI��&m�f�uf��
*�+F��ZU >���c���9�$��/K����6����_�����!�8��\y��]�����l��`��L8	1��������q��u��X<4�Mއ�$7���=���������1o8�'��%���.1���m`��V�(6Bs��}_h���a��4w뮶Ѻ�4��3i�yO|���]�TfOyv���"~�#��=v2ᓡ�����Z�^L	"��_��].��}�͜G�"w�}s$)�W]�w��;EL�k֩���}����#ғ��Fb�U7ל�G�������r�����<�ٽ�:vF]���`��Q ���=��r� ����C׮��Zq��y�֣:M��%����� u?UUUn��3��o�~����.)����T���+�������p@��ޙ��2v�wd�C�~C!��y�2�xU����Oϯ՘�A�Q�j�u
/�����e�R��dB}�g���57�,�vw�N�Y��뭻��l�ńY��f�o��x�1��,�~��H�>8p���}�'BWB���Zx�~Cy]�U�E�c�(�q%Y�3*��(�#���t��BqoTo�f@�P9����}��-{�ǖ���XS;��wk����rw��Z�}3��=���b�V�\��G�{�8��z��<{����(C?j��y����^Z~�@��儑�Z�!V���?<P!�b:=0�:@UWu����a���0�i?[C��G�yk����l��i�A7���6��+�yކmM���~�"�k�㤴���7���7�Z��?�eD�>O���U�{���yj�*�A�?Q���!�2OC��_�����u�	혻5�|O<ŷ(�%�����r=D�3u��XRGe8}_}n��ÿo��,E�q���#��"����tܒ �p��e�|��՜�W|��:9�9���\e;��{�Ӈ
~�w~̘~�_B!��Z'�|(����C�"(��b~�B��,���$�u���	����q?`!�����+���R��:B���I�Qt�P��֫���e4..�^ k�h���"t�zL��m� ���B�6D?A��r�r7���~#��AR��x�C�B�Ude���/�k����ƭw��9�����ul���ku.��$52T�kc��Z����g%���~�?��B>\ئ����7�+ު��	I@���O�@��im>2]f�!���?��4��I����|8Ma�!��i�Xl��4�dC��Iޗ����r�F������*C־�B�K���Ў<~��� 1�q=]��;g�|a�@��h���t餇+�W��0�u
����D!Fj����Luu�m!|~�>hc��W���h�E����<����O�Ic�YL�B��4����C �,=�;n��{4�mR9�fcPQ�&��]�q��wN4�-��l;����;t���3:�������ե�@���JRN�ʬ�/s��6U0��MXH�7�Aʎi�&�	�δrީ7i��z�퓲>vu���oϞ���ZM-!uN��%��M����}�f6��+C��<�YD��N�;x؝�u�ؓF=wܰVv8�`O �T^�yd�W�&�/m����j��Q퓽�-4K�\�w��}�]q��*�t(���;D9��-9�!Dɺ�o.���Y�>�n;��}�%M����dK-�:+M�K|��:&������n��oWr�x �zLz
fald�����I�2��ա��SJ�<�/]5�^=f�z���c��i��b����n/�=��e`�C}O8nx8��&9��O�"뺐ң�=%3z�0�
���l���%HM[�T�7#nG$Ml�:rip r�PQ�L��s7��x'�&_ov�t���s�N�	�t��W�Fc�n���nٷ�e���~ Y�QY�U�fVDU��Z���s2*�̌b��1���3)��#2�c'-a�N�̣,�fjrȖ(,���j����,�*!�&���##*I�###$�ƨ�jb(��������-f0Lh��,�[#�(� �i�# �ŋ$�$���
��hh�$))
��L�3�����KDTD,H�M�2�&h�*
j�$�(��	2�����J�r�0�*���	

���(*j �(�ְ515�����Qd!fd�U�2ddQAA�D��CNfEL��BaADdD1d9dSNXTET4�QFff9�4�ucSQ��T�VbRE�Y9Pe��6`�&9C1Cf9aM�T7�{ßx~��ۡ#��/�)k�{y�Ʊ����� O�v|����0�>�9!��e��L�����ڿ���o��[�~AR}n�q��f�N���?G5�1�GN*���އڴ���Δľ�d2'!=�������8h�~���/���D�OR��R@;]�A��/ˏE�a�kζ�#I,�hi��G��v�j�u��'t�����b�gOD0�*S����fnϑ�q�4E�)�$��44Z�w��F�H�Z�G�C��=�fè?%*��<u����ۮA �u�� �̖jJ^;C���=����4533�o\� 	mW��g�3���	?Y�����߷�����@�<p�yǾ޼� "�D.!-8D����DiK�"u_���H�ZM4F�ܴ�F����J�������:p��H��r����y��a��Z����dYl��2{��o�.!<t�P�
~ȁ �B�+���̨���`��MXKC�f������j�(� '����:A�&�O]1�O�|x������3�u�#v?L`���������9��W\�� cAtX�uLy�.��� ]�֫ِ�_������<�Z��C�f�O�k���C�#�����Bݿ<��6�/ٗ>�C�������'�����z�:��/
�g�??Š�E	?c���0"��Ln-0�E�Zx�#t�C�_{tא��$��8�Z���}�3W��WZ�X�!g�<��j�K��T(g-ٽ�x�G�Տ�"���c%�DQ껥�����Dx�d{�HC��ט�e��{��\�3���uuu�s��!�Gx���ȐӱRÖ��n-%!�n��{Vy�����r�&�A�[����X�L�I�$��������A��>G�`:l�$�:����]^� q_�\���	��@�ҍ�7�וr�ha���
����Q|�`W���Ml�Vڥ�G�~��'O�H�؇�q�S����n1F�~a�Q~$??�	�!Ăȯ�f��30�ܻWЋ(�al��5}4��'԰�glk������K�D�u�7k!�����UHi~XX�8�?z#]w���3g��5�j�da	�/��-��3&�s4"�h�G�� q�X~C���}�ۯ��>-#�l�k��6��^�ɵwW�7U�9(����:ȡ�R�ZJi��=�]sϘu�8o��8�Ǎ��6�w�]X���s�����a�O�X�jG�dQ�����?!�dB8g�p�hcXB���]�]?qda����|Ǐ���[�}���??!hKB!�NC	ՠ�'u�D<1}F� z���+���9{I]��z�<F�:�x����q�;]yx'cӇ�P��~��|��!n�~����a�_U�p�3��(�{�W�zP���922�1rˏE�#ל!���w���ǽ}O%u��nw<�2o�tڋx�a����9��֦y���q�wN^�j���7���oY�f�h��c�^�WV��|��;":@�v��l��;̆�E�a5����$�_z�P�]�*`1,B3S#���Od���uX�Vz���S�gƉ?G�]j��:a����������2�&��Y�p(Yc�z!�W��|���#I�sݍ���>�"�Da��)L�Z��8l����F���g��"G���f�]쾣�lY�Myid^/�Ԃ�6Fq���4���K�G�e�U�_�˼�"�йr�tF.����SZ���(9I q��d�"�g�!�ӵwheu��ӧ���4�� 0�n�i�G�҇�	��ㄟ��V�Mq�����G��ve&a���c����}����^��c'�F���_\CMr����+}ו��D<~�!�����8���-Ú'���y�
?
4~�-�k��%�^�'��DC�!�`4Q��X(�=�?ghЕm��P��R|�C�X~�N�Y�|��#�q��3�k��6���c��=�gR{��ƀp���D%�?+#��a�/x��k�x�^a�kZ:������~������T�յ���Mdq;�|Oc��b����]���{[3�[ޣ��Q�猧-��֯]pZ�ͼ㓛N���?��K�f"[_v/t.v�r�B�/�6F����ʩ�p�*=�&�t�|�>!��HZ��!��Ђ�^=��w�9]ݝc�\�����g&upFE��w���r�8Cŧ؁8A���b5]�Y�"�A"��{��H�����{#�[���S��4|~@�(�Xt�t���>�W%n���¥����G��C�nq��Ό��vh�rF8�. Y�j+�i�[�j�����w¥Χ��q��V����!Wn�tGvns�a���( ��,#յwC�]PO/l�>3��?x_t�s����� j�Qt٢0y9{v�W�E~�ֆ��aBj���ڤݾ��یF��|a���qV�nz�:��E5��;��HF�t�?�Ż���k�:�M}g�hV�o�"�B/��<�����c�"j�|D8t�0��G��gW{�G�t��c��/�y?a�*�8���8~$^����0�=�p�c�˿K�#��O�#G�m
��{,��Q�*����u�g�	A���̠E�M]Z�?�dw�S�u��ܠ��T�[�T��}Y�/>�#Ə��?#��q?
!&���nY|z��\j׈��Gb_@n<꭫�o��Xag�_����Dn��z�����1�bn�q�Ȕ����.<~�Y�0��t�E�(�&�m
/���Q���qk`�]��������E��C�I�+s}=L����� TA��Gqp�B�k���6���S�a��O�;k��;ף��=)�~sE~���x�}�_���S�������KO����?�ǿpվ~S�I�.��x�J�=`����ؕ�Q�z�}E��>�v�W���
�nιe�O2�^�@Fp�
|Vw��X�.�	�e��Ő�"iN�dg*x�Yx1��s],�w�IJ=}�O�N�`��ڎ�T�j告�>�k9	�q^�0:�p��s4M6��浚#��r�+5ɜ6huo[����U�4�TT\pS��nIK�ѷ˭8�ox��ܢ\��L�@n8!X�]�]{ص���m<|{
�`v��ݷ��@r��gt���7lf�u֔�ﱹbr�Iе�׻YY�K
넜/�U�>�]JJ�k�����31Nl'��ǟG�[*[cb�ָ)����G���u/��}Ǆ��^�oq��k����ۼ-Ta��t��\��rB��B�%��ʖ�8]�&30fNu���C�a������:/m�fP|�vgG>����;T�!�P��x�n��F�]p��)�Յ,��.$�i��4I���<*�"���w=�2&� Hlɸ����sQ$�Cr��p�������$M,K7ֳ}m�m�������"���,ü�"�"�FP�e�bd�S$�$L�198TTēY3fS�e$Y�FMD�a�E�33Ec�E.��Y��KM�b�IYTD�a�eAFf4D�Se�5��UY)��UfaT�eEQ���UKAF�&�fgĢ �JYkfh�caU�d�T�aDADEe��d�T�YN`٭8��j
�&"�ch2+Xa�fa�X��������~�=���Zv�5i`!�r���n�,;wF��to�yGy�~���c��弟W���!��Z�4I�Pa��D1�]��:w�Å�;� �AZ���"��R$��(οeÖ��C��8t��?��-Ӆ�.]za�$��C�Ν>�8��u��{K�E����C��l<��k�ͮ|�=�c�&�
�Ѣ�!��a��N��>vT��l��(���HM_\CMj�j�On�s"�� �Dx�{G�57�w��QB�Z�?Y@�L��� 3��C^ew\�R&��qb��5�f<y�u�\��j#��r�k�CQ}�I��Q�L��]~8��>����Uyh��0��Y�Ӕ�T��vǹx�=��(�l�"��zo�xF���(�$���#H�O���<&U�x��pC��IsoP�Aya���ԽU���C��B���~�(�������g���z�l���&Y��"���1d�v������Hw��H�����O�=�г[� 3�<~�t�9�Ƶ��&@�}�3�|��~���}dy��04E��ʝ��Z�4G;����1������L��>���GK��4�l�B�
2N�R��#У��15g�ge/��UP�U�F���c��_��W��Z�sy�Ѻŗ��6p���k4o�0�G�U�~{Q��]7�y�H�>�u�~�7}V!�:��:��D	�ھ~���m�t�@;LQ�f����|���#k�^�����֑�+���*�0����܏��<~�Ar��hk�Ճ��b����YW���L����8o�-l����)��=~��Ȋ��6o�A|�F�}�Q��eI����x$A?%lW�?QD#N�}F�ς��"��l=˼�C���������>Pז˞�qp��xOs� ���~� k}����Ͱ��q���sdq�F�J|�{�`:x����h{���C�\	=�ۣr�Ww/�#>��yFeK������V��=O�ZE�?C��}li�+F�����h�G�"����~_
!?絽u��F\v`�;��Z��8�3̋���t�=��.��K,�/��=��#u}��My�6��Cp )7�8�}���j<{��[5��>�A����!\Y��Y߼�W��?2��^<./�n�Z��喇��Ĳ�\z1�1w��h�١~5χ�$^[��0i[^�R+����S�U43s�UUP��W�p�?E^���D
��0���=�Z���ۍ�h��?��2�(A!�<��.��n^HB�<r ��1�f$���{���E��v�ϟ!څ��j��û�v�c����!���Ȯ���<~ܼݭ���ֆ��В>����)��mٞ}���_(א�P�56D:p�6��/z��8Z�G��~�g�k�,����o��|@��D��|pח#�~�o�=�c���<~x�(~��L�+�	?_lwH�[���r�t�h>�٘U�&��0\�L|����,`ɯ7#⺴�B�R}�����TSl��O/Ssη��5kl6� ����~�x�<G����FD/���}/�{{�A��(��(��3�A7^�t���u>�1�aט�
�?	����o��J^"��?��b�����Ň�j��"���aݾ4Gy}�p����;;�?�am	1�9�Q��]꭬v�wG���x��4�d�qT��ʜyv0i�v��C*<��R�Y'� e-�o,�N���0�6l��~�@}b�(g��r�F(h8U�<������Gx6gN�����c��X�x������u��
�R£+���W�S�>����X�I�^$E���,_*�'�ڥ�ި���@a�0�`��N�cZ��H��/�(f/�������}~�x�J�L�6� �H�5�W���؁8A��b�{k�oq;�^A��^h߬��-��6�~4��/�>S��h�D
(�j�v�}����0�!��Y�Fr�j�@��v���h��F���!����j�Q*�eW��xD	+�t�Vzs�_>>#��j�W���I�mS�F�X�0����t�~��{�]s+:u��\���ə��1;����pPj�I{��sk�	.	p�%Cղ9:��B^yG~ϬeeyQ������6aE�}.�Ң4Z��+�>����S�&���Y�l��_����7~��[©5GLH&�6~6�Nl��gw���\F.c�9>^!�:_��7��^#�w�0�^U�&���_`��[۞�?C��H�Ծ�&!�8�SK��zAIZ>^#H�x�4p���3���ܫ�#qdB0�.!���da��W���bچ�Xh�:����}���#�3��/^xH�\��mN$�6Y��)·a����jT�y�J�&�W�$7s7�L���MFZ�V\P�^"x�6^���!"�p��ɑ��3�>F��pj��v�h_<��!&yТ�q�E(iH�_�
�$_?2���YgK^��{wH�}�^bƯ�S_xѣ�u��]^�(��ȏg1�@T���H�7�U��X#ԇ5�5x����P�7�/�zJ`y#՗R��}�+�~�CR����l��l���M�fh���5���3�J�?��Z��4�h�>�A�E��Q�z���;�G"�7ޕ��p�?v	�5���4�JLhi<����o���u&tpT�kD�H:�$Da��(��o/���g�9HL���9����Xx�li�N?Vc�Rr�q��0�v�>6xyqz�2�,A~��}\5��"��@z�T�8�7�c��ը0A6@��0�Q	��C������mq�F 3G�/�TbBb��/_o���h�t�8B#��QD>WVZ^ڮ�:�G�.���wF�C��~�(�G/����Dg���C=�g��~x绶��|���{�!˞���P�����n'i���b�V��wպ�p.�Gj��.�+�co�-��u���됌v�8/��m%,,��;�k�݉�t�V���3�R��#�٩�{��#�ކ�0���Ѡ������.��znܾ���!.Ŏ­�Ǘ�,ܤ5u-]ʊ-t˭:l��Q��WS�\��!��ؘ���"�]����x:X�
�\v���q�:`��A;����3+����J�:.�t':q���V�L3w,-�q�"]�:]�\�F�AuxU��m��M]���;��ͯ�.�S.�Q���k�s�d�f��ݥ�I��+�݅���ɸ�5<�� �΋,M�Y܉�6��^M�
�Y���݇c�*����=��p��9�[��-˼��l�;e�W�V�6�:�g.����h��8Q5)��af�c��K�V��+vGZJ���l:̡�C�2�ךQ�_"U�6,�)Jq6�M�$����G�6r9c�|k��Ͷ�n�0 �Izp٦�n�v)�&��ހI#Q&f�o�{��6�@��z���I!	$�i �h ��2���0������VU�8k#�#2s,�̳��(��)0�"���ձd4�Y�d�AKKCIB�0�F�ɤ��bB$��%"��V4R��CE�V*�W5���>�J"��j���"��Z[�CG�A�#�"I�<Xa�<G
��[f��0�/��C�}i"�<oP+����=kK����T�0لY'�<��N��
�%�6|F6t����֐ʹ`�O|�!�~b�6G��Eb��8g_>�����D�C��x�;�h��l>���߳B	��bg�j���s�M��e:�e8�>v��a�0�� I;��9���@�0<t����?h�=�*�{����鷗�h���	^c���M�p���������^��⺎7���iܳ���۲,�u
�H��a�5gcs�ls�h>1�y�U��9�p���nAX��z!܅^��^����^��Y��Ց���!��4@�ھ��+N��`��@2���qY�9�|�﫻U��`O/�C�E=K��#\�w|+�gV~�l�Fr��B��д9 ���R�՝Z4��z��,��>˷�h��k��쳡 !�@#_xѻ@���
�-�:�{~�ӆ��l�m
ԏ�UI�s�a~�\F-c#e��_�n.2�[r>��ղ�m{��ye�a� �N����V�\`�]2�_��*�����T⷗6�j����[�9'�����&ҮC��v-�!��:�ۧeX�Ӏ�����G���F�]�x�S��I	:����&�3���1���mǡ(1z�,���.uݼ�Ɵ0�z��OB	O��osNVz��%,����ھl]������˶��<�g@�n�
��7�U�s)�3<���u�n2�s�!k.n3Ι;y9���)�5o^M9ʯ�ǋm{l�R�6���ßC��Fhg������r��W�<�z�Dt
<-<x�Zg�����DP����{���:��HF����]��}��Uj�Aؙ���+�]��/�.3m��au˟X�=�Q\3=�3�L󩛊:{a��K(l�n�˲��u��{�Cy�X'���m�,h�n,���;��ze�xq�N��晙FQ��8xq��d�fp��9%�2��qy�=2.G�3:1�t��MwPvJy�a�V��,J��Z��Cl�dA�Y�腊y���gr�q���F��h-3�S�W���b])=Șt%<�i��\���n�l�&��ɉ#�̢s��,��v���6�e�����!�t�;�v)��K��=�4e��\����&C~�+.7Sݭ�����WK:��@`@`lM9���@{NZ�b��%����	,�Z����6���!��T O�2�fBi��Z���I�i˯���o{p��35��}C~6d!����6�F���k�e�Z=O7y�C�g�Q���y��~��w�9{�{	̘z��tD���=@L�\��X˧]ݖB��t+���Uk���2ĭ��c�>�@���c�Ν\���//ɟ_VΒv�V:�hq��"�rQnw1{ ��L�t)kr٢k���J��39-��t�n,�|�:k�D�Ϳ������3�N������,5�1ֵ�c�fЃ�)J�DB������r��ގ�L�\����A�{�����3K��֋��%�7K¼��]�4����٦��Շ���R�ƴ{ި4��:�o��C�]�՞/>Z�K�:#��<�-6ӄu'OM�f�^���z�z�(��+�)�c��3q�ps�tm�u��3df�a�-Ќu���1^��q�n�5�/���i�д/%�����%oL���h�
'�;�^n�?5�!o<���"/�s���֢�ڤ�p�*䠞��R8id9�R�zR���}~Emj+�BbrV��3ǖ���ȗ7iO�^��QM%W�lRgs6$�r�鬯z�r��c@���Xd(�K�4����T^Ho�x^�7��r:���J�EW3Rd)���=��h��hT�{/������*��`x!��Q��M]	|6��ZVf�����˼��z����޹�J���m���.�j�`��} �&���U��Q6��t�j�Qկ[f!���~��W�L̖�+�GB��|	zg�������ܺB�`&�ں�Hޞ�n�7�f�˸�Q��ق_|��%<2�w�C��mc�	0�</r��H������w�Ƭʰ��z��_��:�fnEbT�Ư��ٖ���O)�)��4�ZO4M���Z!�ڥS��";"��=�$W�r������ҫ�[;[]��eM{��]�&�\޲���ս�y�;7,k}�u�A-������
{h�۷)�=<�������f����D������,51H�Ɯ�E.��5o�i���Nmq=H���:�r]�]�N�Z:��	f�r#Z�AM�zꭎ��6���֕�{�25[u��8M�7u���7Q�f�!�\�`���Qov8m�I�nj�2Vg]ͼ<y�)	����T���F8vi��j���v;z�.����[[}�s�f��xN��֩����ڸ�G��S�4��x�{71��v3,�	���R�]9
�ьۧ��'�v�a��8��қ��Al54c��{��2�/5h\�S��[w�J	mje*q�C":i�dk�ʽ�a�7a�>(,g��{&qa^�T��E|���l��:��U&c��������˗J;6WW4��C�����VInIF�E4��X�)[�FP&4ᕂ��!E�>�6��ʻ=U{R;j;f�b�����k��TA,����ʮN�e̎�f�w�+)GZ�c�q-K��L.釵�ԥj"Lm��I"��l����#t�18�A8��wb�9��e)�@kw��7�p����H�;$�n�#!�3��GR"���o�I ���%��9+ID@dfa`�Z�AF�(��� �(��!�2S,��5����L��zׄ~��N�޾~}��_wg�����#�+���^�)Ej�*gm���T�X�MJ�<.�� x�Aںx	Z}��(�H��~ח$]�:N���v
���qͅ��-z:������ةF�Q쇺p�9�F�[6�uZ���O5lW�	�G�SR��5Dx];[��{v�ͧj�?&Wr5�3���������9i�5:����N�s�퉺��m��f9Gfp�K�9k�$����7���h΁]��^�S���@Ջ�e-}V$t*��:L0�^{�y�L�����=����N��:�%�>G䏥����Kq��@ވ|8�g�۲[�l�+c�u��n���_S��X#%�C��d/x7b��}S74��N�o�ۺ�5C���u��aszR�8��~N�N�bL�`��m�����p���j^���_���:���Y���)܎'�����"�>��R(��*{U�==�����y|�_U��:v�2em_��VR�����
Ga��i=�W�r�/��;)�X 8hӷ�#+r���~N�V�P�^��j��N"��Ͻ�cޠ��C3�m����X/љ�>=pt��U�P�*��|5�x���\��k�2�Um�ٺ�;�.�W�gͰX�)��s����y��wf�Sl�]�G���I{l�^7&Q��V�V� �V �8<ՠ3��/y�Q��Nԑz�=YCr� �s���p��Q��C͔���Ѯ�_��z8��%���/ɊWV�����Jm�V<h�<(7���dc˝�jE:ӿE��m���W�x���榰�td����� �J�l\��P��"��7���s��+v��a�u�F��^i�_��\�̛�ojK�NSsV���EGڜ��#�J�[+�&��Z�{4Ŝ���K��U)�����3�C,X���B�?mwk�F{����ӈ��]-��1�Ԭx/pw/o( �~�u����ǋ|�o
u���f 2l=]�}�t۬�X��q�9e#�6�aՙ�,e��=��7Quԭ[���(LYZݯ'6b޼[#)}i{Z��R+�鹔��%�Wx;�h�ötǒ�Ds'K��(eI�:��vk�.�H�s��)jv�����vk+�=�!tPJ�(���g�_s�Z�eI�%�m�W��}�(}��.�'�(�vb �~�!=�n�[ɚ�	Z9���kk���)�	7y��T��\�7�k�x۲2^��ٳ�[��=�4��P���}֓~;��t�6~��f�m��k)�%��{F�$�y���C��E�8�=N�ͧ��F^F�v�d�)�[�7���r���z��8L�X�Sڸ��y�nWNxǜQ�����O�5
!b�vN�{ע��pəjo�Dw����&)xݥ��ЩP���r������k6zrl#q�6�!�tY.��f^Lvw�zH������,&�X{vt4���B/���	��t5�u�������\�G���$��pCR�T&���C�b�3IQ��;N�J+������r�
�~���js��QD����}�^[��󷭬�U���/��z��U���O;{'�M�;r��F����ز��r�,4k9H5P����鵽�u�	̗��;���S�6���!�˓�v3ꃳymte%�{*o%]u���r�a_�������"�<�#���zrͻ�<r]-.K�����ʳv�@�3m4O|w7��V��T����s5�{$��I'I��Q�f��g�_8�BɎπ�b��W��v�Ǻ#�#�F��~s�kۏ�7���l]���(��p����C8���/p #��l�C3�>�D��t�a���<:��F��e�ך|E�"��aPȶ����	T1���-8C����"^���F��4�$|o6�s'�E��֌��NYb<�y���&-{�U��)��Y��L��z��Xmܹ�s��̳G�xγej�<�+J/z�Nſ5���Z~�l�j|������h��f�5�\Z��
:���L&��y�m�)�]u��Z�{�\r�k�@%^Y���B���*m1���C�2:���L�v�Aԅ6�����po~�>5=��bb�SH*�}�bΫbܧ�T�:X��/�c�!�+�b��y:j�5X�v�0����9��������Ƚ�X졷s�S�x�p����d�yvD��шӻ�����*w�߂�v*u��`�z5�";3�y�X���RV8��@�C����d[���<�Iɼ�ҹ� �c�(:��XY�ᆲ�49�]�NV���O�KuM�s�[�v6"�_�~�s���.��4[ߑ�;h�	t�k�IY[:q1}��9s�)��-7�Bq��W�j<���'�)��ͮ"]:���w�\1����R��B*�u��y�oK5��`��HWe�\�o\�7{��.҆;�m�5vP|����nk��������c�N�N�l�w��nn��'^ޗ��,wƱ�p�4M�6��Wzhe��YfGM�у�u����7l�e���ч��Z���=ň�0�z7#�����s��J��܎�����Hɱ��X��[�F�oU�^M�QNt�>R
����j����9Mƣ�qUC/y��pՠ�r
02ʦ'1֜�5���dQf�fAkZ��S�NN�ZĊ��,2��̃�D�6�|�sN�~��k���S�G@�7m�Z��
����b��*����T|:��p�S4�Ю٠�V�o�/���V�+<���ޅ�p>�����靆��\�䞿r��*o�W$���i��Q����;���d�H���c<|�˥��Ǔ�(���:�z��k��ő=�q����y����~�8���z��^ﹻ����������\�H�#��{!z�	s�bֹ�w�k;b�L�i�_��t|��X��wu9�Ё�LN#W�%^�+}��9�U�=L��m�o�D��^�w��]¶�D��EV���� ��a�1�U�f�Z(���Y���6L��Ѻ�i%�2hU��0q�w�]x��-s��a�����`X)ݙʯ{��{
�#�P�Z+#s��6�[8�[�vsP�wĨ�"qn�"�Վ���Y1�2[�h=���JsfaxxAs\"y1���$��4Mj�=�MZs�yZ&��)+�l�޻pi�ۤzv��jk���xd]����]_7ՍU��sܗ�N1��V���3J�'��cm����C�y�O�y���W��׀��͜}���b�2���>66Z�-Vs�Ue*��'^�z�"pt�=��{�t��5r�qH�U�;jƼYAS���V;��V������2��v�Y�KtM�ǘ�dx�o�Ћ{��f�h�.�JGyb���p�����a�����Kغd��d������+�H:��(y�{��W�+ʳW%����On�f�c�����$�� 8�w6u��	��=^�X9�)ꗑ���wr��X���K�ՙ�%���5�������B_�nU�ޗ���2c^ �����zi�;�)�5
�"�m�&���~�X�	Tr�f�e�`�镫ϨӞ^������y�tI�p���|m��f�g���h&�H�Z�6qf������gԑ��(N���(�Τ���ѱr�xHo�#م1:�/��=���߷*�)���lY����g�ZS+gܫ\^3����b�
L5����~�P��כZ4�$ڿ8�Mbe��5v>U�^�T��)�*��6J���A�@ZJn%ev4����^�=�5���ŭ��mp7ý|8x�B|EM鶑�ŞOQ�z��m<�����3[��)��Uк�^'nE.ڎ�����WDO��"�^c#ǥ����Sʮ�9�k���ۻ��jG��U}^�ʊ4U���nq���/-m$^�yM�x{;O{Chz׍���q�n��c`��}u�-��o-WM9��pj�!ɶ�g�~�Z5�{���y��s��tp��W^3�@���gB��H���[K���|�*�� ��ɫ3ka1M5�q�!��k�m[`]���
NiC��b�U��b,���/�Net�����Q����y�x�-����f�7�-��6w�[D���Tsƕm15 @���v�j�yYH]Hժ별Ox�Ջz���i�}X)��hh8w������zj���7�PF�hs�؄��:'^��!N:����mo���:����`�5]��0pR}R��j��'�ݛ&s�zlU �����4��m���>����#�� �|ߒT��[��ۃ���^Ȓ�ޒ��z���~0-:+8��?��J��oa��Ù�/n����ڣ�5�kC��,���{���-�4�j��� ���Vȁ�[�4�J�i�N]ϳ�qL����5���Q-�$��=\x{�{�>ٟ�c�Z]8p��/�v��a���du�>��H�F¥��<��Q�Q�|�f�Ns�_U�ח��
���|\��L"(��^�M���Bs��]P�@}�5o�v\�����UԎ��3np���I�}��]/pP�6��.�}v�S�����}���e��'�̮~�V��|�=�����&�v��؅�E�D����"V�\ֹy�����<�x�߄���i�� �I��K5M�Z��xS������;כ[������Y��E�P�>��V�.�f��Ώ���әZ�ߴ\k�Ҧk~�7Z���v�\)>��M��{��D*�㉬��iJ����%�5x��K��DkN�������ԕ_�T���G��g�:�F���k�rn�s�ËE�v��L\���WAu� �X1�5�w�����'C�KšF��;3��F���K�8,G6�&V(�.�ʧ����.wPq]���79nG�b�t�u��B���ܣ�>Ҷ����N[�7{E>@�4�d��O�
��zQ�\�:ԟ0�On��3��c�O�o�nY�Z�\K��E��Z�t��H܄� �'H+�Y�i�7)�v�ԃ֨]bzfl�����2e�x�.�� ʈ,�%ʽ�IV8���T�.�S\�֍�÷��K��fr1�n����[��͙�r�&�
�xuMU `l���Ւa�6���Ms:��kr�.�*�`�Y�Zg@��X򁼣�@t#�w�c��U6��_wAM��ar�䃵����PO�5�td�V��5�.E4f�Y
U�Z�uNg���t���]����rF���J4U�b1�b�Vwwn$LYd��3������y\8w�����0CQ��R��ֶqq�U{\�`�JD �#33)̳1ʙ����ֵ� �5a��Yf�ET����!"��Z̳0h
�z�my�����G/c���i�0eK{*Ea陈��U�q�6��W���C�����9Q5w�<o,5�m��Tk�*(�S�|�L�|H��dȬ˘�<__+0�N�F�-r¢({��G�7gV�È0�������{^�����c�r�D�d§�+�{�����P�*t}Ҫ�XO/ұj�Οr�Ak�7k)o��������;�����#����ڜ,�P
7�q��YZ+��4�XA��]o4P�ҿ[���ʗ����4{�K�%�xm��1q>5���44��<W^ �)�O���:��r�bs*̟ENH����ݓ&1x�s�i5�*euX�G�q�J
s��d3���0y>2e�ӷ�j�sS��:�[�^�i^-������¸{bզ��r�q��;oy(�|.��ӗJ<��`z��T�s��œ�Cy�D�qn�qg\)����w�7���u�k���p��c /qb��܏��
��ݡ�c͚XȊ�U-+D��U���t��z�')C��׃ry���}H�Z"h�}�X֢��r��ʑ�j��=O}zPGh-�\�6��2Y�K�6���GQ���7m{�F��?k~I*��b�{�;�2�1�ѭ�&�����-�w���I�컍�ܔ�l�y9�%��}�Cye���k\��8���}��#Ev)�!#�Qۙx&���?@G{\�Wޥ⮅2L��s9qԎ���{J�ɯ]Ӳ��ҁ��������D1��q#
�
��3¸-���m�2����}�U���&c��G���f���������k����!7}�7��g�5�&/b�*Q�����ȯ��97j7Z�P��� �lq1�z�2�]�dI��j���Cw:�IA�;�K"��K(����k���}�����/C��9�'oc����;���9�W��ڼZu�K�5�kW��l�h�Y`�c�z��ʭ"�z
�Q�F����]]�i2�{4_<���h�����.�q�E�t`�he�)[CkF�k�˕g_�7�M�3�?d�'(�s+�n�s˼�q�٢oP�L��Z������M{�B���@��}��ڽ�MY'��SgbUf��o��CKfm/u��O5�M}�U����h{�w���a�v����/�����j�+��qI��&�����sC��eAS��?b[x��{��P? %�Q�whfQ�k5-�pɉ.�/6�ݔ��W��������l)v��f����֓k�쵙 ��њ���]�\�J�.�F��uʁ���U���yf�\WV�HU�O����w�%���H�ڥ[��a�֩��5e�r�w�
�Y)ȕ�����^^��QN��0�q���Y�ܷ��|������<���2ח�U�����!�J]g^Y��ok�+����BU�Y����U��y/}z�V��2��dP���:�X��H��)�9�\�w��7k�m��>Π� ͱ6�+X.��]�ކ�RQ��XY3_>��uFS�P�mvz�ʴZ�N	PW�ݴ4*�h�y�X�yô��Uu-'[�;E�S��y$J/���4�i�=��L5$<V"j����r���d����`в��U�0�>~�F�Ϝ���s�v�پ�yA�[�p5�[�tHۻn?9�{3s'2<f��3\+<�6�QtU����eM�JP��ә�l�i����{$�rn�\���Z.�5[��iU� H���[�&p��ot/�7������'>�o=0(��}4�Cl>ɷ�ͭ���6�4�7L����Y;�^��}��֫��:Mp����Ȼb6���R��g�whW1ֶ��i��B�,�U��٫��6���|m�
�'���[ɰ	J�����m�
�ឃ�\�t��������yv��7j��N�yy���bg���X�ue�q�٩�r�py� �=%K=ϥ.�Oo:�֦�nX`$���3F�t�*�(O�`�D���2��Lp���H,^��^A:�B>�?h�[7��x�L8I^�t�2���՜��E4zU�6{|����'&j~�);N�6����ٸj�+��Z�T'�|�̃��K�1>�o�1�tH��(�������	��ң�YSES�%���������
~��L�U=؟͒'������`�֎t���M�3������xG��bJ(��kQ@������bv5�';<p�&%Ł!��&{`���gٝ�r�b��b�O�>h5(�
~D5���v���=!������Di�w7��~ ������?��p��ӯcGA�~�9^~	�Z4�MÝ�v| ��<���k��׼�఼�} "���
)�(|Q)1t}�����Oc���������~���4�Q����>���a���UAN��)�s�h>��b =n����	M
��[�F�'.�Ï��`��!.�����3���3>�\+�7�|����I�=�gߠ����E���~��
GG�sw�Y�x��pDl
�)�~V���W�����F�ăh4����.�|�z�6=��PSܼ�K���z ~�>'�o��?#�n����~�{���'������?�p�F�����?o����~���0�}�?٥UAN>C�>�!�ܧ���D�!>����h��0�������b��~������>��>Ʒ����������W�x���~��O���U=�}D�]|O�`���=���p�4DX��}]	��)��R�}������?�	���0?}�`�9�6�����~����p�Nv�@E8 ��RA�i�|�,��}�r ")�.�.����|C���^�6���e���\���0�W�!�9�v���:
�]l�p��)��������)�S�QT��>��!X>��@�X��_a���<��p�Ο�x��)����_cl��� �|���}��)?D�u��̦����'I��?��AO��?�c�| ��f }�����/�PS��8�B�������`v ��/������ t{��.|� 郔	�G�|�ؘ�@���>��@o�����v{A�r|����?��W������g�����}���EPS_W�'�M�M�����6�ݟ_�tG��a��=� }�O�L �0���>~�����>�I�@� "������@���'p)�_��~����>ς �ؿA���!�v`�>����v�0^����?ks�=�LA}��0S�����y�.�p�!7N�