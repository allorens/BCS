BZh91AY&SY׭���!ߔpy����߰����  a��,�   (�      	 �P 9� (UD� � 
�	  �P/7�	QEE*{g��a��:�.��!AE ����:�]d��.�<��k�^�9�mL�ޤ�K��s� �70��>���O����O�r:����I����@��l�� 
 �%n�3�ݹ��e��N;�.��=���nvr�i�=�z��\ ������u���C��ݜ���ݻ��9v��]��{�s�\�ΨHG�:��U��{����m��n����Ӈfg�s;��Gf���=��������)Q��{ۤ�=]w��^��G'v=5u�׼Os��˛{us�v�i�  ���#�F�ڜ۶����6^=vc�wWna��uм��ym��zn��^�9WvrݷS{�g�OsN����Ͼ��|����Um�Zv�θ�*.  ��΂a���z�mzn\�;�ާg�Wn�oZ��5�<�z�.�Ĩ�����z�������w��{gv�G��η<��u����A�O{����         Q@(          P      	SИԕ%COA�@�LL�L��DI*��&  	� ��10�d�)�T�@4      i ���4C �hd�1#L �SU @�4L����M�=���(
��1J�C d�	�12��G�[�$��&,�����M5��?�:os���t��׫�cm�[w�s����/�f�۱�6�zp�����?��e��9��l��wf�\�}����p�����w����5���̍͛6ْ '�L&��աo�&��$��	�!�HdUUU$?��Vm����>�1�}�|�|>�����{6���~���9�Yv�<�G�ھ#UH�挬7WG��,�ʂK(c��2�1�I�H�c$cʕ�=VX���ї*1�3�f�����1��1�Hǩ�1�d��1�mQ��c:<P1�@�&1�f��et��iь���1��3F"\&1����c$F&1����J�Q\�eJSJ�)J(��m��C�Y��֐2��,c�c4�����c���A�J1�f4�1�`�1�c0�Lec��Iь���guI:�G�á)tp��걐=R=L(�H3�,i2��f��H_� c$v��ִ�
j�4`�tlC0e�MI ��2�H�t�d��� �X1�Յ�}J�a��0ޓ��a|K�!�}Lc7S:aD�&2ǉ�ҚC c�c�Y��>��=L��'I�#�t\$�QI�da�m�1z� �q�X�L��c�3��7�e�d�dS��,P3�FҎ�>� b�I�3a3L��e�e�L(�BcC��0è����a�Y���L���L��4��)�c��iP��P�1��V1�:�1��f�>P����1��1�b52HΛ
�1�e��/���!�cfbcP�1�c��P�Y&1�P�Y��9�ä�X�G�H������vFM��`�#Fh�1�֐`�A��3	��1�����C�3Y�1�eRe�c:[\C�[�ę1�����e2��1��1�>Jc�3c�3Y�c6S�3ǭ+Z��-kSm�C��q�j)JC:6�D����3F4�c2�<Hc:HƓ�1��c&1�e��1�x��1�2�	�e)S�6ʕȥ)
qX���1�X�3���1�2�%� cr��1�-�2�P�1���&1�cic�1�c-�1��1�1��2ǩ�H�@���@Κ>n����1�gJ&h�U��;�0e���(�K�1�1�2Z�1�)��F1�
L�1�Ѝ$�dBcΌZ��1��z��tgK5�I���H�i��&�1�,c:2IgDm&2Q�&�x�k/�4�:Lc���4��	Le�aHe�PtgF�$d�22�"�Lљ��،���I袈u�1���L��r�f�Pȥf���4����䍪 �L����1��LCC\c�t|c1��1�v�1���e��q�cM"�h�X��cΔ�:w��#���I�Yf�7Vn�u�ie$ΖU�_K#,e"$�2��.Jhc)�X�QE0�$^a�$P3J�Je��GY�r�.x�.d�29$	�GX�gKf��q��$Z+S$e̱�zY��Ҍ�
���C4�Y�4��<Ld�>1�9LC�C0Lь��1�>Y'J0�X��J�,�`��ii���Y�cF1�3yc4єF�3H�Ȣ�%�	 `�hY��2�e2�P�C#��v�1��� �tD��Đ�����H�ä��X��S�q�QcP��U�2F�N�$E�b�#&2���a#��k2
�Hc$r�ь��2vc��$c,|gF3iY$�ǉ�2� �V0f�SC�Va#$}]�&YGx�3���2�C�1�>jdԘ��Hʴ�2�-� c6,���&2J%-
I�c���TC��$Ƹ�P�[�>$�шe�fjc,���H�3���2F1���Yf�c��$c���1���e1�ш��I�cѵ���2X�1�>%�c�2�t`��c�2`�4��2�Y�i,�C��1��V1���S#8Y	���|fc0v�#��1�f��c���ec)� `��1��K(p��1�gWF1�=J1�f4�h�!�c�\&h��z���	��>2��1�0ckH1���1�tBc$ec3�f�Ӣ e!�ddіiD�3H/F2L$|�Hh�����J�T��RZS��!M)��S�J��q���3�R�yJB[�2ь�$c�:>1�P�2��C0�I���1���0��c;��0c�P�2�c�t�I!b�C�4��Ӹ���iB�l�
>2�1���P1��0clc:3�+L!�P�$�����ff2�dq�e��e0L�������4�8S�ʐ�8�JR\=JeM)MR��%M%�ԥ;�R��0��&`�#,��1�(t�#�cHfb��1�b�F2F1�kD����3�|fc3��K(��Ր1�1��D�d�3F2�KL�F1�i�hHΏ��2Fm�!�gL+��c�C�H��c�c�c c(gH��1�3H5�21���I�ZB����2� d"�1�f�c$e7�P�)�b���)�)N)81�H��H�1��c�D��)�!I�6�JE)JR��I��H�c�t��1�3x� c,�c���@���cΏ�32WTc%�>�1���$�1���1���;1�3�2�1�c,c�$cLc,c)� ��2����L��c6�d�����1��3F��"�C,c&�2�)LcC���[�ѐ���1�c7�1�c)�c�jC1��2F1���c3�f�`�vF1�����Y4�Ɂ�eK��f��c�X�2D&`�α�ef$�A]����(�TE�w��ȥ?����̚�Ц[��?�A4~H�I��u?�_��������ß��rzR	_ѿ��y�JMmJe���_����kk,��?�9�Zoi�;�n\�gr�W��E^�f�}fr��<�+��h�ޟ��|_O�̔�����������v�$�dn͒Y���2���g5_Y}���6I�~_9?JS;ޏ�7��0����I_IC� ����<�Bf�'�{2y�O]�+S��*��'�@�;$����{���P��;I6��pa���do�{�x�x�UW�vY��rb�a�kǏ??s>�S�����j��)�
�8M��K�ߝ��_}��/�ν�)�&��ߦ�Kݐc��}���˯��JC{>�z�,���{߳�ǂaGĔ�_����}���ad�q�VwM�{;��K�f�����{<E{�{���F����P�WZ�"z���=�^��鑓�3s�ُL��������
�~1��d͝���:k���fn+�7R�VFZ���NyBq��]�*E�起��wpѽ5��}��M�{rX����o����N�{��{W�o���J0?W�0���QI߳N�Xp�Q�y������/s&K���;�X�O��C4M�퍧���n9�38�f�nC���kj�۠{��8����v�����gGܺ>���W����{�e�[%���1���R�%��|2�ϳ;�����f_FBg.!�Ň�Y��w!��8|�z����ެ%�-ʜ�Ksw������V��jb�A3$-�.fVA���N�V�2�|S��l����p����<夒��W���I��w��+��#�'��s��H��M��s���ż��Q?w?*�%�z����Fw�y�u�v�'��d��,�ǩ��{��ˋ�U����o�{N����K����۞έ�y�`+O�龌�x���[�'{�/�f������/Vwn��W;�N��Z��	����n��)̨�lۊ��Ow�ٶw�K�K���՘�Ew�ؙݾ�3�絓/���?�l�]�O��������"���ٝܟ=���g/���y�SU�8�+5r��Vr`�7h���5fT��c�T�,*�ϟ���w�}�2�>oo4v���F��rp���y��r����E� {����]�[�[��;(W�҆6~���c��ge���3)�gw��;�g�n���7��f�}���o﾿i�0�қG�=��	d_��'N;;gw� �a�g]�`RzV<�\SXi�������$�{|f�'��:.̝�Wo~&<�2�I2a���<�NO�����㳙��d��}��#IW�K�7}.�H�j��ww�SQS�<{��RI?M��yw]��!u,Nw"��ժIj��C��n$!\��ʉ{��̥�)ҏ.��b�\�6vI�g2?��r���.�+����+k��VQ�E�C����a��MH]����*K=�6sp:���ܹ�d{-W��c�?�xv��f�_�3J|3���&�}�d� J5ߞܛy�rU�	��ӆ?w�!�Ʃ�nܘ+�G�����|?NiN�9�}95l濔��OZ��c�oM��Wc�e�Q�4��r�[��,����L��ݍ�,������7�|��)�ۇꧮY�+���M��T��Fx�����n
g���>�|K]�s֝�#�s�aw�>�?L}�Y�I=�����{�n�����ISɉ��1��gd�~�Ǚ>%���f�{�B��vȧ�Mg����F8rK�;���3�.}��#��2bnO�/�����[U�#N�����ɥp���I�ͮ�K��[��_o����u��g��|i�:���G�d��Ux�
u��v��0q�	d�]��G���ξza�꼄}V����J���&H3vjג"X��
Cwo���[W�vl�y�l�q�I�;����>�;�2��9��9e{n�]U�Wjw�]s�U�w�e�{:9S�D�|�Ǒ��>�0���ό��'�96|�j{��g�i~���}�1��^�&vS{s/~>���9��5��9����͆}�__���n>g~���ϥ�6�gn�U�ɿH}~����{�;���\�5��Z�������Ƿ$��ui8x��ɿ���M��z�\�[�b2+),����s:�Y3�4�9��Y�znoJ�v�ۏQf�>��׼���ӿ��,�bر�"���;qR����nw����Ω�7V�S]�ً�3&ں-{T�����2s��w;��r�5
����t��O:��J����^��&�U��%?_���'��~?����Z�o��d�n}�w3}ٹ<��x���Q��g�;��ݟ&��نo�w1k���dY}n���d�4�0�RR�vw��TX�j�f�4��.Q���V��Ŵ{Auw+�+mO��ǒMjO������g�ؾ����'ֻڳ.z3�b�~Κ{��ݔc�$*?~w�o��,�y~�/��q���owrwa��4��a��4��Ul�����wg]�<����{����p��۟_�[�)�����Ս��Z�nY����p������z����XM�K7s�\nl�;��;��?v��k���]���L|s���sEf~�_��n��ϣ�g�(t���Gi�0B���ޗwd�9����M�@o��|�1�u��ҕ���U�{���$B�Nw�v�d�2�;IՍ��@��ܿ9�;鹡�|}���s��\8�R���i����s3������y����hX����AF<ɝ���6�bv�;|,�}�N�ٓ�Oc7V�f��C����n&
���ozm�sWh��Z���{�w`���5�8��_��j�_�ՠ?j�b˷9��vm[t��s0�W����֞��餿^�<��n��w;��v�qZ�~-��.�SL������{ݜ&�דl��:n�{���+�*{f^�+�m��9�nveϡ�=̝5�f�߄��z�3�1��{��njXbe��{6䊾��1����LM�sK��.�\���4�欄k��g�ӗ�"�H@�����qQ��N�[yDS�97�]���Z��=�����v�;7�������G�~�2��;6�MD����K�.�.p�����R���f/ĽϽ���ْl��{�.�ٷ�k_�y�y�?g똺p��3f�������\�xz���ׁ�õhwۿ����W��n�C�]U�w�3�NȿW㗧g�[5�~}�{��b���������Q��w7&�=s��bW?)�/���9p��I���;�W��*�;.f�_��a��?Us���B?�)��S������G����[ݾX랷o_<�ۣ��y�-��$�{.��/>OS������۫��wJ��Lc���:�c�������Ch	�mq�� ��m�ԉ���CR\����M�5�&���9YYU�8�AX��]��[��K��Z�X��4H����:޶B�+F:���Y�4�L\\K�b���Gl܉al&����f��l�0���if�f�cb�&�Y$�d�L%qv��Q*����Wp#�qؙH'* �A���K��p6�»[*��mm�-� j�m5�r�v��Bm3o;�B�Į��U
$�b,�-)$ej�
�ɯpkf����Y+K.�hꖰc!�-��4%���l,��/�u�IS��ˎ�H�Y,�y�R����n[S[Ɋ\�m�m]��]��jB(�H�J�k���L1�Z�AFW��Մ%��Q!���	(M�����i�`�X�e����]c,���6]q�cPUI ������c4�Q��4q,�k�U�k�3z��\��E��%
��j�	C��kֶ�M��҈�m6�|�@!*m.�BP�g��X�(�R�m���@�6��q�nԷ1aM�GLB��[6f4�dI��\�i�#E�U�?<�$Ő%+q�6��%LB�6�u�����!���qc�p���͊�6�bX�1I��׀�M���J���e����;NEm�k���tL}����YBZ_��a�b�w���%�8�J�B%
��ݺ�75����)J��Ģ��8*Պݑ����7e��}s[����#���b=	#n�Ѣl�M8��cL8���,.��3^��d��l�p���
	�,�NE����r�(�:�6�ƀP���!$n�H�B��2�l��F�B�(�Q`�Y�mڅ�<dz֒�Pkj��tob�p"�	��h�+	���u-��m:ȹ�!�u�.��'y-�����ˋR)<�T�R����m��j�c@;v$�����R]Զk��5b�%k����-ĭ�=�-)f��65�f�J�6r���[�9���*X����3W�aͨq�!Ybx��Y�a��
	K���+�Rj�6��s��N�9��vѠQ�X�dlÈl��+�T�s��߹�s��_�oc�{��rⷷǎ���/�^W���<Y�ݻzj��'�3��z?_��=�3��.8�3�.[qc�8���%s��/��ߛ����r�m�����m�m�m�m�-�ݶܶ�wm�-��i��v�m��o[��m�n[m�m���}m�m�M��ۆ�t�6��m�cm��֛m���p���p�$s$6j°ڛ
��H³e
f�6:ٍ�emBX�6YV�(!⑷m��m��cm��7�۶ܶ�m�p�m����۶�m�޶6�m���m��6�m�i��m�M��x�6�}m�m�m�����UEUVꪆ���1������� FRE�s�s��vۆ�m�nm������m��m�޴�m�m�m�m�m��۶ۖ�n�M��zۆ�m�nm��m��z�m��7��[n�m�uTc��0T0cь1�a0�#V�FPKm[P�g���AAb*"+�T0e�ሊ��f5QACUE�U��������l�f�$���������~@�����o��>Gg�����|���tw�Ԧԥ!JR�uN%Hyǔ�).��2��(ʐ�)JRQ�1c���1�1�d�QFԥ)O8�)M�JR��4�$c0e��c$��"�1�`�:iei,���1�@�Q�J1�c�30d���ef�C:1�c(c�tjS.)JJ�eG�R�ڔ����Q �1�1c0�	0��(`�X��c�X�2��2H�)JyIC�R�R����<�bla�Lޏ���_:�]0�sKi�T.
&aH-u��4��e��H��Jڮ �v�kt�XB�i��m�Kk�:��.��Rk�#T��U��i�j�#�� �Z��G@�^�Ը����6���y���̶X���H�WC[]Tᬐj�$�!jw�\c0���c��i�V�k.�����ev�CU<��5���M(��0����  ��b�$e��-�.�[�aI�,l�Y�5��[�].�0�J���[�x�O�gP��˫$��M�/lY�1��H�,���]vƍ����sfr��G�l�j�JP9�����q5�˳l Kn�K(u �;m�*�HU�]��a3���b���9#T�d��@�f#G��,g"y*��W�����$�24��Y��1�T�#��$]3ո�<[]�q�[�8�(�Mv�,.ى6vq��a5\E��kp��)���_*A��m����1%-�h��[�Yj���Sr&햎����5p�<�<��^u+���Vf����1��U�1���au��셲۴���&�;���p��L[�H�A�V]��8�hD�Ս�dԤ�6SK�(�
n�C���+�"�ؚ"�N6���`䆚]Y�{2�٬z�fK]Ӯ���͢�eyб[�,Gu�!�����kr�0�*�q�G��hu�)�VK��i�mXl60�G���G�_X�h�9b��-��\��fk{`Ƭ�t����Wee�%�m �m��6p[�fIu�[��-!˶%;8>Rb��e*��Vy6�A��nEh�j�i-&vԎ!�L�س�m.��O<�ƒk�Jf8Ü ��-����m����b������Ux�0�"����n����W�1�Z�Z�ukJ�R�R�4�4c�¯�4\����'�*Y��)��@��n#av���kqe
�6���ṋ�×\ce�˙K(�Ѩ� �t��)3a�6�g�� 2��k��$�Xm�����[]R�r���S@::�2���-��K	u��oR��V:j���&<.�n�г8�@�`��֩y4��'�y>�t1uDٛ�$pQf�Ww.l�W���\�n����j���nh�l�22#��C�F`��Q�,�m�(�H��	KN�d�ntШ���N��ПxY=FVxu�jaM�qM�d�kH/˦��kV�ҭ2ii�STi�|s,a�:va�\P�@��tAi�+�� f��Ōf�1�2�4�4c��4pѰ���ʰb|h�)��o�/wў�rj��7�K
;5�-��:�D2���єY�)��3�������P�Y���}�Zsn;����x��KIj`dn<GU��� �t�gx���/����١�s���IT/=�6�$<iC,��4ь�di��1��a�;�<h�����X)T P�"��ɾ����gUh�j6�ҟP�Ϗf������t6t�p(�yd/�J�֢��nM��"S��h���MOJ3F�ͫ�+ma��VP��J��'���/���X`��������L��U� ��mź��J)O(�4�M�a�0�DR��\4����1nl�F�4`Q����������Ӎr�Z�לע�ȢU�X�U�+�j�aaK��|j�ě{��τ�iG��H�(�"P`�_0S0`������t�\W�R,G�&�EUv�=6l�t{�O��L�N%X�W���%�-.���j)O)�4�M�a�0��vC��D�T��X��ə�c�R�.��m^0�hD�ቫj'�x:�)������0�;�����n��N*�+��	cQ�qF�vQ��tׂ���3]���st*�XjCZ�Ł�������� .9s��O����e�`��b�o���E�����f���SuE�33�R��/��������G!�3�u���q���)�4�ycc&��5���gÁCG����F�җ{�J[n$�Y�@��5��߾�&Δ�CBY>�����/�Vd�T��Z�b#�$kk�)���.��8{2t�P��N2h�) e�A�J,e��F0c0e�i�h�3���!4��,�L Y�Ua��Q/��YСg���D..���xD�9'/���,KL;Kber�T��m>v|s9�ק`��0Ja�	�ẅ́
�kf��ٖB��#N�)aN�D������!p}0�C��
C����hN2a<)�,�M�!�2�$��4c�ON���̆[0Ư��sų���6���f�I�=�Ԓ��4���ykm���� �$+����W�&��MD%����L#V6낪������fNa�&X�X�a��,�.��4�t��b�Gy�hVD�{3�F��0�Q
���33Y����Zx!�'j�7�/�!�ҏ��ê�-�=,�|4PCG��c��3Y��Y��c4��KW� ��]a��'�=$|�c��ɓ�9�^����]�|c����m���ŪgvGO�EV/yU����ag��աi}=��=H���鲘z'D)�K�9�v������ѐt���a<�J(�JN\��!p�s��2M=�$Ob	�U�J�U��a�:��Ba�\K�uJ4��K4鄘Y��i�0�.�.�;G��������ە5��B��r^|<a6��RhZ"��AQ�_L�uҘ�@72��˄�up�6���Lk���Vdnp2ݝ��֒�,��k2��k,�ŋ/ڴ�����%~gEgޮB5[PQ��L1n���yL.�:}���Xh!4Y����m�e5�n�귺�ta��2zY�FO8$�T�R�a��K��ȡ�N�u��Г����ߊMg����am��5O'}_d�#��DrTr%���	��H�Z�|n�6EST��HO��5U��V�Ż&���ϻ�[�^�)��<Y�4��K4鄘Y��i�0�3UU)%���(��A��e��\��U�Hpè�=-M��.-h{O4:����Jc�+zus�$#�6*\��܈��,=	ؑ�A�&�FQ�Z�{��ϰ�_��}z}b���;�<�d��9��������`H�bB�����h6!���+Wӫ��|\$��(5�)yq�UT��3y�A�I�+0ӱ�s��8�,4�xd�,#����t�i�ڋgK[T�6�m^b[.��D���g��[l�%Nb[0�a�eMiE��-�-�E�ҽE�(�"-�E��f�o-�-mql�)�t�x�6�V�m�z��h���ken3n�֑�u�mo5m��il�-2�V���FѦ��Ǚ�Z�m���)!�m
CHZ!�#��E��"�igKf�ĳ�-[MZ����3H�>E���������>[6�z�ifm�ml��ͺ��l��my�f�qm�)l���3e���բ�̭�ZZq�6�m���[V�e,�<��yx�Z��,�ml�l���kj��][V�i���ZٴZ<��gKSV�6�mdi��?A�<��p�_���m]w��������E�7��=���5褹��i~�vA}��L�N&жn��)1�1�W3Yk�c�u6�'�YPS�5T�v������<���'��[辗��]G9��o�=���m����{޻�����[������UL�ͯa[�[έiZ�u+u-��kZO��6l-���m�#%:-
0��!��ѩgN�kg����w�|���v|fI�d��K	X`~�}�M���E6��A@����Rh�߼򷐆�K!�� 6!�&A���	p���d����(���5$� �����#-���f-lі�7
:5�$��	mm�j�N�Oy���; I�'䑉���T�e���0�7ȍ�*��qPO���$�'sd��N��� �qb!�$�&D��Hl�&�LkC�	�0D���(c$�g�#!�Bi����K!�������l����'��%�h����q^ �1h��)�(�0Ҕ��o�|��J�Kiy+Z֕������]��!�a�O�ID�
ɱ6j�/s�~��ֵ���ޜ|�n���p�-��G^�m�3'$:��g.�o�3m6Ku!.߀�D�'�Ɲ���J���������P�¡��E��k�2M�'}�7	�;��F��62f�+�:9�,
�;e�腆��u6$����
06p���MBa��[i��7i�v['����r-�G�t~��N�@�1��%��	 �h�XD`b��&�e(��� ���Q�}�p��B��4P�,
�s�j7.f��Ġw�A���S8�p�N3���|��[��%�u+u-�)Zִ������y� 6s��A֮f�@�.k��0�9w�ڡIq\1����1����D˙��U؅�5��؉H����_G�@k&�-[�.r�RD^��Kv	.غ���,t��^%g����N~k���ɶf�O�.�Ԃtv69�0�i��j��nh���,���$�iE��Eèb�W���<#]#8�����Ȟ��%!��Э����St�� 2��Ɉ�5��CbX�8~B�`~���I频d���	�j�"O��B�:l�I?���&�,��SR�,E� T����:{��[�����,����F0� �e�%�cę��# w�
-���L�T���Y>�h�|��%�}�"���RtH|yI�ɱ2p���"OD�'�!,]G��dK�AQ�PM@�L�[67 ���:j�23�H8P�6!���$lS OI��q�K��+uo��D���Ҕ�kZ^yi�{rۈ��0�b�g�$Ѐ�(pH] 9(|&������sP<�&ϵ��6��;6�M�l�H�kk[�n�qc8&�&�H`�B���h���>��I�4ÍS�9�͉80O>ԭ���6��ta��	�M&q��y�ф�yĄ���G���wM����$I�i)cJ=�����̑����E�%�}�d���9���a8&`R!0C�M�AH~��Z���'
���d��6�����LD!��IA_De� ġ��'�.��2QRV�$���/˨|ۯ)O)i|�]K�-��+Z֧�[,{U�gZ�ۈ���&Jޮ�'�H�>��&�7��3[�� ��Ѳ�J)����ɉ
�N��D�F'�U��1�ċ!�&�A!�	$�EE�;�n` �M�'2M������bFId���4A�6}�F�-R7.�g�&�a�IH�鲓��"T=�(�P�a�F��{�D	X;�b�/�w̷:x�<�
D��?��7��B ��'D���s5'�y&!�Q�>z4�f��O����KɆLI?�,�����5!�Ad>a��jd
�LT)h��X\�֚yǖ�|��K�q嶔�kZ���s���B�."#3���.�d��:{�K��42M�<�-q�ц4�!n��0o�u�T�����;�%�����]\5Z���>w�o	4d�X�`�1�6�-e0�P���!ѓ�E,Ht�b8xe���Bo�0�2`��6�Ov�I�d(�"%,���6p,�6��`�ؐ���kcC�:0�I�D�MD*|T��$�D����pԆ�A�tdؓH`�F`�a���:Cf#!��;�*\�L���>~d��� :3ؓ�%4�,����%�Є��A�yd�(q���<��,�R��6��kZԧ���[m�R�$8������-��ZAVȉF�%ܹ���uU*l�@�|Շ�LwS|�E��[qdT8�c0ˠ`��K�!�DNF+e�v4g��8`j܈���ڌ�b����b�=f(�!� >`��w4��qｕ�������Z�j��ǐ��1�bS8B
B��2k9�@i	����g����Jȧ�AC��B�D:2O�BF�9&��I��?)5C�!�0
'������	�!� l`Q6  �~pL�i�`�h~d�� �` ��:R�D�a=��·36l��������	��L8S_�b$g�ICs��9��2�7�ŕTƝu��+�M���8!Ԝ$�C�����L2F#����J0�~���bb�Q�c,�m%/���%Ը�ͼ��kZ���s;��fy��X2O}���Dd�������9�M�,%q?	�S#�~a��0�g�!�o^Z�f�_���d<�� OJdd�&���K'�hO�<:}�\�T����	�ِ�aDD�KFCm2�!�6�*���d�.����q?�ѩT�TYȳ��}��8f�<^W>�2�uNe�~�|8hDO�E��l��(hFn�ѹC@�0�s�S�P���
(� �F�C(���O�K�q�y�kZ�����4'�qҬ~�ۇ�%b?��ÝTÚ7�B_�lLO"~�z�tO����6�}�n�@�Y'�6h�A��N	�MdC��kv{���.\ZŮ>%�����! ,�������u�~�M��'��_�~����	�Z��4K���h6¦%ա�8'�Aa>�=�/�6|Sx���Ne���2}����QC�f�4q?l�������]B_:��yo����L0�<3Ǐf�%\T�!K��*�����">VE���g�b�b�"(�TXET�:!�Cl���/�]�q4��W�e9 5Ր�G���m��}���L6��l��%�DY��k��ۚ:zt0<>���SrǸrr|w���g������Ύ���g>�p=8����rFl��x}~�!D�>�{��L׃�����>�)���^��8�6��n3.���f�f�ͭ�Z�J,�[6�m��J�f��(Z[6�q�E�1�م3�-,�[6�E���kfVͣ��"-mZ-l�����ѵ�kfͳ�٧[{[6��Y����kg+^�ٷY�ۨu���E�H�4�)�D2�V�6��m3�Y�ml�6��S.���<�|�+F�|D��3�!Gȅ���h���Z8�z�E��۴-�|���)mZ2���̳��~|���[?>C;E��[6�m�5h�ٵ�h�yn�jf�gK3ճl�kq�[+G����x�6�ڵ�n����K2�R�x��Z-l���l��[6�-�R�mm�ճkg�g���[6�6�[6���-�[6�����o���^�.�tS*�s2��ޕ3���Srΰ��]ǫ���9	3qh�3dRId�����̱ژq0,�d&olΩ��Է�=�#�!�yU��ߵӬ�R�kO^����X{	�)u�����Ԥ��'.��Gzl�M�q����FMļ�5��6�_��:>u�S8�ʶ�b�L�X�ӓ[!*g�C��t޳-~��������Y0s��Շ�g{f�ք�층�uS؁�s�q�t}�^LA)m��m�o6��u��케k���㑁��M����]6��W<ӄhӆd�.K�V��iT�φtTfk[�nW3c�W7�U���cgX�TÎ�v��u�wo�͋V>���|�7��y��iז���z�<����;��0($�V<�V�3]�����)��߻��:�K�v��Pm�}��}�{�ngp�7ӻ��;3a����͠�Q�Ss��${w=��:6��͵f�%?(��ps��ݦ�n�k�Da�f�%�d�ZQK�*ڐ+T%�4�ab�x*L��XRi�-���A��Ƽ��-�	�Y�^�d\���7'm�l�f�)��IuÆݐ�$\�ZϬG_	h�dl6��U��m�AF�9W�f0y��.p�ܸ�9�����gU�V�GJ�8���r��/��`7��*��@���i�S��Y$p�}���Ͷ���i��m���o�M�ꪮ�����eqku疵-e,gL0�<3Ǐf�����H�*��'�VZ-��C]\�neV��c�fȑh�YJQ��T�Ұ��ufu�Un�[��-q6��\G\���GV�L��na���t8�m�Zv�@�p3]j�-qF�"͙n,4ѰŹʈ1v+����lW�+�c�q^2��r�0@���컞�V���������K�5L>��-��ӿo�煴4�w2�{��w��J?' 4��d}ϑ
:M�s���������r�Wh��'�	�&�����:���\c��6��}c���A�6yҞ扰�b��7 ��'-{[�Ū�ާx�0��r�� �� �C���3QR�TȤ�c��qT�(U����~^\Z�
o�4���̟�L�{��m.2E�
i�Υ�O�S�q�y�JZ��{�L�\���1��� ��Ɣ|>B�$4)xe��Jfe%$r�X��Δz��h�g%��S�pI��c�Kql�fqS�s��8�;d�u丗2�^o���K{�!(���r�wպ!�Yuth���)A:Ya������M���p��Fj���a��o��`q�|�R�֥��T��6��Z��)*r!��n���j�A)�����v�Q���q5UE�8�>��|`�����suXC��Y��ۼ]jh��D��bj���s�H.d/����U�mp�&IQ*̘�>R�>X8�vjj�4rB0�b��������L��vh>T����-��ÇAQ @�(�C�G��bTW�{�#F��(�/��������!sNeg�D ��X�YǴ���:��|꒵-e<��o<��IZ��1�Y�f��!��>�����),^������QN����nƩu����j�2b��`�a����L;�_+�G:!��g�����������Δ!���<�|��֯������>;6"'��X�(c? h�G_��̞>,�D�x������|[$C4�O�4�c-e<���ykR���{Fy�m	�i��1�M�є��2�{�������e�SRXz� ���4�����G��,<F�TWjmQ��m��vո��2�$��8G�Q� B��&�����g��mnK�?/&��lds�L�0��Lx��b�z��MV�i���M:W4��@��~2i�ek��U��
�]\(�t����ĩ���r�4B/�Y(�n�*����vy���5�P�>uNc�J6��(B�z�!ś9&����6ns��â"[�^�n���(��˟�凹Gu(�da<��A����]r
Gټ�3)�<�HmKu.�Z����J[y�JJ^Zc��"1�zC�*�"~�0��~i�B&�ي�������Y�\�yhbKꏑ16"��|�>t_t�p�"{�j������v~>c��O���a��}Iw�}��
:n��$B2�Dt���6^^}T��1���f+xŭ���=���'�~��ˍ���Gg��8�}-��9��{�����>9�{��|�ԾK嬧��ZQ�<1�i��^�I$�!
�劶����8[�S�;��6"j���xjr��:h��S�7��/>���BP~��(muYe�p��
��,T�#�U��9�7qgT�Dሤ���g'��`����D��a?��n���������6�g�"h�	�?�5��3Ӈ�&���a���<.�$���#1�ո��yjS嬣Y��i��f�a��l�/�����������u虝4}�ن�M���,�?aDNg�/�8���Pӈ�S31C���+�vX�.e�����y?KjB�KF;ȋj"/1�Т^��s�n�}�,C�t����Ҋ,B0�&I\�����cG4Hrۧ��9�P�b�GqW9�kZ�99�T�>�4�C�!e��&R��iZ�)hS�u)m/-jRR����ڡ\QلqFv1c��M}b�4�H�S�m�"ʣ� LD��K��)�c6y6-e�U�bh�[�5���{��V:�r���˲O B���һ���좟krFsX���Ȏ��B��}�v�}w�����L�k�z]]hԶ���飧W����gC��SNs��x�DG�H���>���v���sf�艔��~=��X���W��3��1xg<*,p?��"��xH>�8l�����`3Za��<; �d$�a1�pᣱ�"l���ɿ��������������X�D+�t\\��&~n��a��G�4aDD��������읞�vji(S�yĭIR����:�R���֥/�5mk�Q>�S�U����t�JJ��32%h].5+��F�F,��;���T؈Y�M=��t�4h�"|~O�l�z�'""s���m���s��L?M�"]]�5H�VTF�Hrv� �\�tE�d���gi��e/�5iTAG#x�B��g�I�$��\0D�%9�ae: �7��j�8��n��LG��6�mŵk�Y�u�-�[8�m��ꚴKL�-�Z%��h���لm����h�Z-��-�E��Cȶ��ml�-l��ղͭ�E�m��ٴY�n��-�[=E��i�E����fγ��kgH�E�h����j�h�L�l�յh�m�|����c����-F>)���|�F���e�CKf���2��1l�l�l�)oj2͡��H��j�ͭ�[>K6[6��Ϛ|�1�?>S_>gO��Z�j�[T�]F�g�f��V�ڴ[����l�"-���[6�ڶ�ԥ�D��u�l��v�m��kf�f�ͭ�e�umZ-�=[6�m�mkj͸ͭ�[Ku�[,�1��Ӊ�&���y�`A���;�p  ��}~��؁|`gb�Ǎ��L��,��I�ge������uh����4���Q��f|�v���a�"�9,ڡj]���v@���D��#]����kL�ϳf���^��E���k:@Γ���x�����^�~��m����m���uUWWz����������ben-o-+RԴ)�:�����))y|�eU�æO�+7�^��M��L6����æ�D�ԓ:�Xѓ6(�p��҆!p��%٦����}ϥ=���K��%Mu��V++$��	�Z���/�żł'��ϑ�'G"rC�gPRDH��B�ݷ������0�7�7�b>�}��-�8C��m�>^0��>-����/���
uN�)q�jJ[�s�U8y7)�G�7��}��):�b!�}�ڶ���UJ��
$�n���y�aeX�BX,�^/�z?�,B��}�����ã(%2�KHq��6h�i�|���F3����T��h9O���{���_�p7'�nt���ۦ���!NJ3�$��Ǳ*0A��jRa��
�J|�O�8���Zԥ�hS�u-4重<3MϪ��5SE�ݕ'�s1��/� �x�T�.�ڱO�ydj��cFly14�_���B1���Q�!.��*pn��J�r�A��F� ��լ�~�����³���Tⷒ�b�b�bf�;�U�5��&�'���GC��A0/��A�=>�Λ�������~��fo��@�xuW,F�*%I��	4>�#9�9���w�m����,}n1�1R�'�F��/���`I�n~�Yr(!F�+��p�s
<���Q7����{��B��e�i�K�-JZօ8�R���ҵ%,�q��v�A�9�:�:us&��9�^tpʩ��)�4GFY�y3�DWR��	$���oN>�4���D8��4x~?8��mo���������e+��%EET5DLr>bҎ��C���0���mR�gaD��y9�AD�#K��<v��51SDՖ �-�R�)jRִ)�:��ǖ��)i눈�c>}�g�y�7�?[����z<��!�4`vj:�(�=��_���'�����\�5��9��wj�\�ې�lh���Z�A(RS��_"-.<e`�LZ�B�U��> �/������XQ)�ve��:h飇��"4~���,_�����l�d�b�_�A������� 2��v'D�|xt��-kJ�JR��JԔ���A`���*�/��S-\}���&��M�߆�F`�������.��>Gڑ�RX��i��M�K
Q�j-�&�x���_˫�s�_-T�pК4��R�Y��
R��0���hwy�t|5�V�}�K7���^:J�(����2UT��(,�dqw³�O4�����f�c�����L���0����i���T��KZ҅8�i�L<i�i$�ʅH���e��r)'f,X�Q
�y,�16���P�y)M٣�!S4q][�6-���]q��Y^�b뫯eH/4�v�]3c���Z��3�����B{�3��O����ڊ�"������sM���_ub�:�������W���-�񮟙�Klp�1�oj�xb�+��n��G�N�|�;�5'C�>z�q%@�?	���lЇ�98>O6y;@�Ml��Ơ{6����t?�|hќ�Hr��$S�MO�$�����5�u]�����9U��WO���Zԕ��j(��#ꄠ+���!�Q�ZT�-KZ҅8������w+刨���TCE�C���x��v0J���8I5T+0?��G�3K��3.p�a�Y�3g�6&Oƌ�N�h˩Q���Ķ�����ǟ-�<��}[�M�-�i�f�+�G2�%T1{�}��Qv)(���L}
	X���8@��.I#��X�:I>D9�ٌ�9�ux����>Rҥ�KZ�B�S�J\yiZ�h�Z�d@�B=�<�O�*D=��)L��'$�q�丙sG�������4 ��ӟ~-�uM{��X��)�W��uD�C�G��b�B�j1Q
���ݯ-#3�+y��|/�ТY���.ff\r����ӟ�E���r=w33|��fP����YA4l�6D��ᆍ����F�i[���\JV��k[�[�q)K�-)ZR��+1�5�Wʨ��<\�Oܞc�}�W5_yF�<0A�xt�{��i����"Wޕ�,���E�ȞK<G���%�����Fu�{h�"1�i�mA�6�3�cKV�m��-(���P���"{�z*�<���.8��n�x���'~i�el���(d��)�O(�(}#��xc6���:�mjR��ʔ�8���4�8�yJS�6�Rʌ�qHB��6�)IS�iHR��)JJ�2��eJS�h��1�23�,��J�3H ��E�e@��2�(�)����4�k-h[*J�y�)�)�%�R�B�R��)�%HeJR��:�R�-o-o-n!fֵ2�ԥ8�:Ҕ c�X�30�,��d�����e�c0`�X�2FX�2F1�Όc(gF1Ael����z]�M�7,���~��ɲZ!�y�b$ۓ�8�;��P*��8�dʦ=��}&:*y�L͐+�F�=�`"�Ů�Y��s8	�����{;���D&���wt�$k���~��_�����7�����%�eF/GDU;��3c���I�kc�n���Ó]���;���GM��Moc�۸˗��	6���w�(��|u&�q��.εr���}�f-�4{�����,R�!R�Zj���ٷ9.�͛O��b�[c鑙�b�䮕��QU�Kٔ@�pD�]���5�8̵�C�-�k���=5f�5��(�=e�q��F��˺�Һ�U�9m��3u-��b�%�m��e�2�P[�i\�rō����ktf��.+1n�;\��m"�2�9�ͭ�D�`���7WZL�Wf���au���]����
\��,��a�YTU�Tv��ҹ�S0���9�[�[`��0a��Hݖ�Li���dD�2�X�+�Ǚ���W[�R���Bn1؝�BX[+bd�.<K�Ν����m�߽�-��~�m��y�uUUUuUUW�,����kRַ��ѝ4�N�x�OiR�#`�)��سV��*�[pb�Ae�eԷ%�qY.���,�L��6���mΥխI�!%�]-�:V-lIoP��v��5��㬡�,%�Ǹ7�A��5����L9�Y��K�������G����cX�J��!5�Kkk|!ber���� BS5���7����-��4���ȣY0�ۊ��]�ˉ�%׋Ӳ仓9%������g���f�Ř'�%�C��x����!hOYA���e�4
a�ލ�56w�?o�/�gaN񎏴Q��t�<�����Sp���B�ݘ���q�A~HZ����J����	��K1̒��^G^'�q��C�n�QX��ߚ.k��D <�E����e)M��e8p�T]�le�N�����J���}B�S�J\yiJ����,�����Bq]ɬ]|Obl>�t��ޔ���=����,��
���7�z�5��Z"x�18p�c8-M��-���d�O���K�%;N�4"Z`wx�k미�������36����$?|�yuU�L$ &jGe���K��(<F�Q�h."�"�AA��%<����I��p�V򒵩kqkqN%)qiJV����zq��F3�l�GO:Z舚�<��&�D���Ӽ��G�g�7�!'��j���l�Ҟ	��D75��ճb}��a�}��ʎ[ӯd�mB�lu�M�/����8Μ�o���0���Mc.��4k*i��^8�w��a����DFB]Gx�($�K�:gr�g�����$Y u�Шm�J����D鬵Q�`'==�xz'Y�#�o�Y�R��KR����JR�R��)y�c�3�AB�-V���Gy|�D�@�1~!U�'�!(����#}%r��|��l�V��d�����ɬ��R����?`��c>�)�Do6K$�Hi���ޏ����ٳ��������� ���e���6p���;���f��C�E\_�&l�ym��̥n^��5��|����%���p��I��Z֥�kmkqN%)[�JV���zu��̙fc�;H0�dkU%�Nim�q�A�D� ��;�2<(��Q�̰����ܰ��1ڮҙ�|Ie|��*x����,����ȋ� BX��9�ߦK~���V�o1��es�5�MB�������9�8��QHjRS��Ӧώ�-<6tɣF��x�#�j߾Z~���6~�S�"h�,i���7ha�6\K0A�ƍ������4♄A�iM6{���]Uj�����.；�� ��X�J8�k�r��fגf;���k���}}�4m(��c"�5�R���i��,E	���r��5)�8�L�mN��)jZ�Z�S�JV�R��*�"=q��i&�}���@��'��L��%J>,�hp�F��+ݛ6R`I�J�'M(��(��4�.O4e�\�'O�Á�kL��a�
x��?��R��r'�Ye.\�ATr���2�q� Պ��'9�Mg�~	/��%3�F�I����O$�x��Έ�I��E�)KR����JR�R��/�)"�IϕQ=;]W·5��ϘT2��U�F��6�l�a��Fa�(�촇HKߏ���8{�j_�5�.����Z��䨸a�5���h��o�, +��Դ�tЂ���ǎbf�3^���P�X�JڱN3�#�4К��fN�Dκ�7�����bB1�O�ξuiCku�jZ�Z�S�JV�R��-��z���DB2���mt�y��������GF�ꉥ�����O(&Őq��&ev�c97=6a��NB�C�~~��^]&�<xPCwv��*0�-���n��θˎ�h���Y�܈�5�B���" �i;��,���A�=��j�]jԺ���?aO�t0����(�}�iL�����ֵ4�����/<���/"��q�`�U��Gi9ZO��<�BDk�Dr�J�\�5�Ŏ����ط�X�\ֺk/Z�:��a��r���n���2�3gn��_,}� !)4�c���Wpu�Lת�Z����������,6�P�k���eG'Q&(���ٴD��+�^0��14X�l�a���o��9њ,Lf�E�ii*'�$�C�Hű��r��c>)M�Sf��P�J�6q	���P��_)��m�0����?Ot8~`k~��@����_/�����MD�U��M���(i@m�#vYR�y��iƷ�{��N�> ��0�\�3e��P��c��F�2��6����|�2�����ԥ/--��C��Y�^Y1��d��4�%^s�-����!��\m;ogn{M�>0��6�jvBN0 �B�����Fp���n�O$�_QJa��0ޗ�QL���Z�p~)���b3@��=�B}�V���n4?��Q�k��Yj��vޑ�-�u��[�7w��:�!n���!3�3�$�LIL�,�=$��*�#����(�r�ic0�֧O4�)JS�R��*)JJ�eN<��)Jy���QD8�)�)M)IR�R��2�)JS�)JeM4ʔ�%HS�R�ڔҔ�6ژ���ʊ)HP�E2�1��L$ä��x�<��qZ����iJRT�ڊ)��ԥ)N)J2��1�`�@1�c0e�ee	kZ�ӫZ���eJAJR��fa�Yc�ΌegF1�0c,c#��1��2��b¤�S�L��O��K�.z�1F�>j(x��4��w۪�K�~����!����f��t��ϵ�Z�Q6|3ϵ?����a���`��V���Z��6��b�|�r�)JT	�>70��ܫ�T����M(�6p�O��i����[O.�˝%G���2bj㳽�y���m�����m�6�~����m��߬E<#�%kR֦V��R������vuT���;�����s치f>�lD0م0|�����H���ڥ��/���:&��:d7��0�O�r_v���ݫw�h:@��2��k��ղK��!~R8�ŋ�\N@�f4h4Q�{�1-0�q� �8�Ze�m6��|Ne�Nç�������$��a�Y�á��������M�[���8�Dq�#�:�Xrb4�%-o%jZ����JR�������K�L$� V*��ʨ��S1��F�����J �~*e�Ҝ0���1p��m���T�!e'N8��]���b���E����=4a������_'ۚ4p�]}ڹ�5�����=�rpؔ>ߛ��t��,鰕�x���,J$�Gxt��߫j3��a�t�߫xp�ύ��>�O����bc�(�D�=#6��)jBҕ-JZ����JM<i��a��#vn�%Q+�U"B������Ц,��\�䩯'��1��Ri���Bմ�p�,�c��l5��ڶ�ư�v�����7J��l�����aP$dl��~ �+ �y~X�:-B) �f�;��X�s&��
K��/�"2�%�
/�܂�Y��V=0C��6l�����KU0�M�~?Yo�b�ç,�x�ԓ^/p�6|*S�OC���ۥʴ�g����#�d�$��G��e����4ۘ�o�h�3�4�D�{�?�Ud	��+ihYd�n�A���Of���!��R��-����0��Z�)KZ���S�JV���N�SXi&�UD>���~�x��QE�!���2���,��`h�C)`�xQx�V��C�N������&.�!�|�C���5�\�&x�2~)f�~����Dħ�<�;1�#��NF'e�N!@�V��Ge�d�;n����bi��Q9��a�~;ixh��J��s��<,����f�˦�g�g�RvD��i���疵�KR�Z�p�M<2�4��Z��ܤpU䒈|p�2�D��~8�Ұ�E�C�!L<���h,�"�qc�r|X`�Y�SBjj~�vzp�����,>s�-�r�.�B\\f����Nz-����p�4��F�w狘�ƹ�u���P�(rR�s�YE���A�UO�LL�t�!D�a��o&͌�&���1��剂e���=��@g�dE�Y�i$�BV�[�JԤ�hZ�q)J�Y��a�	DD~I$ ���L�3�'�Dѡ�
�a�H�:Y��	��ن���3��2����mn�8�4���6��.�>�FA?Sϝ�\N��+�0��xxpB��0�w񢚞M�h���g<l�Ź8h�!u��؇�}0)K7�~\�I�M`��DPC ez�͒I\7�i�A����wѦ�yԡi[�R���ju�M4��4�<W���eB����:�J����Ȃ��De�-���z�:#k[3f������ٙڐ[�Jsan���Ū��j�ɮ�/XZ�Ǻ ��~*��{�=�j�|�+-z��u�b9q�Ä�����.�c����Kf�j�s���p���O
PB:{2.b�*���H�I%X�x�� �29"ç�E�/^%i�<�c��>�����>����
"
zXY�����76a��ߎ	�٣�2��V�l�CG��s8�V2�Y�˷:��՘��e7�^�2�D�OCF�?Q%��h���1�B�Ub"��%kZԤ�hZ�q)J��R��Kc��oCF0�%=���u��0i�`�k�L�>��R�Z0� ����0��P���
�.�xi��>���x�B#�5� ��L6%2d����~�m�ꉃ�ѕ�rQ�l`����X-�TMw�_���r%̵��T�'�e���D FV�Lht��Κu�gF|h�u�򔕭S�%)Z�J^a⤮�$��ƉH:$�G+�$K:&-)��lJM���ᲆ�p�����g�
"y}_�SV�P�[y�T���Tt�O�'��2
�q�����/%,$���8�K�=�)�ьAn0@����ߦ���vN,��y��0�JV"��W�B&t��h �!J�e�e�)hu�)o���hZ�t�M<2�4���� ��Q<�HA�D�QEC�$L�W������0�b�hІ�Q1m���ی��	w`M mI6�
�ލ����b�f�Tse8Y�2p��XP�`��L>>0��������JR����<;>��{�S4�ng,Ө��4�0��x�ɴB��I��Dt�� e�:t��^E�d� �V�a�'���,��H�<�+ik|�%��>R��)�d�e1���t�`��if�Y(d�1�e�C4c(�)�)M)JSj)Je�TR��(�)JQJiJq�mE!Ji�TB�R��i�)L�M�K͸��]e����Z���\ejRT�mE�R�R�ec1�fdc1�f1�gH:H�H�2��I��$��hZֵ�y�T��4ꔦ�1�2�2�1�0c��1�1c�2�1�2�x��.�V{ٙ�qa{��gvx�Fv:?,��m���Qdp�,T��5]�LxLx���mVvIX'z)aɽ�w���a���l�0�.'7��\O[�If\�3 ���56�-�˺�)�7����Q��S�=������w���_7��ϴ	�ń����ő1}{eŗe�S�R
�`��%PLߞ�n�z��n��{��Շٮ�LS�8���=�Ǐ�Lv�;�C���|{��b��L͊B7��&�'�Y�d��m��N��d$�f��d�fba4t ab��h�11���rծ-�w^�3ٸ��M��c�/V�Ɋ�I�bkZJ�Mc�۲�6)��5��P�&��l͕����%�MrTeͻ��e�m��f;�I��9��rf^]xkOn��r���f���w>ۭo�#������z�g���5w/�Z]O��uTWy
��N1HZe�0��lM���.ؔ�K��Sa��k��	ZJ2ͥ6e�hU�&e��&�+sL"�[J8��f��%����6�͚�Y��و�n���tf�s��J����j@���̡\lh+�MQ�v/6����ZJT�:B�h�]��m�4�LV)%ʂ
S��E�N��7[m�m���{������m�{���m���m����B�ZV�)+Z�\JR�:�����G���Ѫ쒪+����X�	�R�K��d�L�KB]4t��nf�]Eg"J�5.^�#�.Å���2«�[���{Ym���(��cL�YMq��h�lz������K�*T�k�v0��>y䏉��:����6�;R]�u�T/e��l�-�:�E@�H1�mb���?�%~�O���^�hj6��N��lރ��u^�7A��fd�Vw��{ز���Sܒ��2�&C�(����H��"k���ɩ��a��6�]��C�QG�i_\|!
W�Ks�%
����:&�8}-�{�M��~4o،wc�����a�F�4t�C�+�a���8�pЇ���>f��=�dL��3�=M6�9�Y[�Q_-Â�ֵ��=[4pل���6��c9�S���P�%�JJ���:i��f�a��d �������}����[L';���xzp�rH +�82Ĥ�z%�W����ϛ��2�l�Q8|l����p���D�����C�nS흏��H�������VPp��*v�UJ�I�	�:D���B�%�y��gmч\�2 e���M$'�f�a�âW�t���f8��6;��C��ZT�o���Z�\KM<2�4�4��(�\�I+�2~�um٣���[L4�'KA��KA��H�Ji|I�AD��K;�D<�R�-�J�Lum�Q˙៸ja���0��=���!A)�%Α�4>�_4ӥ� �Ϳ�D����=� ,&|�$�*��
<<���;�[��̷�����)R�[�c\Ɯ|�/�-k|�%kB��JV�R��[�b���5��Ut�#�w�=\̝:xt��}=4|&�R�p���U1,je�jf"�4�����V�sȥZv��	��E��V���~�FJ%3<)$��6�OR�{�IDs����_����4�a�H��X��+�E�'�X`��f��0�"!���ή��C�K�)�/q��iO)jR�Zе:�R���M0��ԓ&O��gj��צ��Ԅ�;y`o����]o��,�I��q3�����#f&v/B�ź��˒�m�Q�'�cE("�U$I%�$�}M���ωw�.z�ʙT�Pw�%Y�,y�ڱ�O�y���Wٌ>]�;ڧ�;Z)D���<T���#<�(����������x0���٩��8hؘyR�Kl4}�)����3�Áy>���O�<�~iiL���k:�:�Ay�8�4�l��N���&�0��[��3w9�*�iӔ * �dի��S]Yd�%�4�E��:�┕��4��J����-N���ju)y���<�q�QY�I��w�TC��Npu�n�BH�s��Л˶͖c���͚(�0��J~�>0�V���M�D��|)���P�$���;76h�ҖԴ_ǧ<>^�W�a��&��G�q̸��q��<l�$v3��//s�2�4F>��ir!�ˏ6d�6$=�w���>���D��K�SD��Zy��i�Jԧ��-K:i��f�a���ɏ$�d����s��Ҭ׺�k�4rY����w��0�>;���(�F=�6�,�$����تF��v�C�VT�q��d����V=E-r���BH����=�vk���Ļ��
!��a�ܕ�]ƥ�M��A�����B�F�vHC����8_�f8�V����N3C(zcO	M)��l�AO��x�|{�Ma҆|i'�<�jS�Z�\JR�:���6��ä�T)�Vjح��UD4Qu����l����BQ(0B;�(���(Aߋ��d�T����iV.*]�]J���=6|�;h��CG1���SX�Mk��Ki5��z8p8 �P����BϿ����Cxl��Cx#�zl����L=B���n�~(pA7~�߷�oa��e�6l>���8e4e甧ͥ�-JukB�S�JV�uyyuu^��0c�>NWU��q㼑�a�fUm�[*K]���6���Fg3-%�텰�ٸ)l�i���q�v�lѰ*���s�ı�A4ԭ.VIU(U�	wu٣z�F��f7�<Ǖoנ�,om[[՝��9��g=:Y���}�ٓ���)N��[s�s����I&��� �NO�Y"	ލ4>9Q-*$�'N�$�x��oj���i�,���pt�"3��:GD�P�J!�,GJ}��sM�3M�>QH��#q�Vue��"���K,����� �Β!�ig�y�����օ����O%&L����H@�)$�JPI��(��7�eOq-=��q��1|�E�to�/�[��G����7=�,�p�
%�O���$��!�Q⏯�ټ����:��!��kw���3�M7}i4�^﫽�n�m�Pao���w�G���[T�6z ���ý�$$��)��C� �I"����ɘ�)��(��t��K�o
����iJ]R��+R���A���dΌf3`�J��N��Q�!JR��J)M�JSJR�R�Ҕ�)�YQJR��!JR��)M��q�1�A$���eIFf�ͥ��ʊS��ҊZ��Z�R�q��IR�u�SjRc,c#4c�1�1�3Fc��I���1c,��im�)Jd�)kZR��yo<�ҵ2�)�)�6�)�)
R�b�h��c�323y]p���O�bjL�U!|��ʠ�K��}Cyܕˏ�8c�-�0��F�\��5���h��V/u��V��)�
��M�[�1��s�\�	�n�i�EGG���VE��ܫ�b��ałR4$\��$
�1�S^x�o���F���Z)F#[5�iFkY����{RN(U����R��j����m�6߽�{�m��~m�{����ꪪ���fY[�[ͭ�JukB�S�JV����N9Q��-:I���0��ʙ��� E2���s�q��!-<�2��(ᤞ7I(�b$#�,�$�902�ja�¶��uT3���E_5UP���"|`h洭���
 ��Jz$�K�ș�c���z*f%�:P�"C`_qI�WFH^��0_&�0�1m�E���>yO�S�|�:�h[�q)JԔ�籒"1�f�F�HA�AM/��D����Έ��
�H|l�gMp����w���JZ�2'm���R*���:��T�S�@ ސQ��[���3���@;笂æ�|��9%H��J���A�Daj[���-Զ��,8q���p��B��Y���Q��A�/�u蘈�R�X�a��}��%��)Jm��JukC�Ft�M<3M4��G�Y5J�<��ĵ׭*b�-mK-+5u�Z�<Y ��>HJ
��U`� E�� �@4T!�uJQڱ�j�inI�RQ��lML� !#ھ���3�}�����~������x]Wmd���!͝T�ޣ.�vhQ��8�0b q_�{P���(e��s�A@����pAٲ����MiL�07��?)Dï�[��g��Ņ)즧\��#���c�2��ʃ�i2|����ߩ|��̵�3�p�Yqt�U
��i����M�@��>Mr�$+�q�阙B��$���tiq�-JqkB�S�JV��/<'H��`H�Ī �uϕQq��bwF�<���'U?a�٣A��bs<�_#�J�b�$:"L��Bl��)|��f���N�Ӏ� �����~6tFa��&��v�\n9�-%��6����3Bf�J0�Լ�;����1�G��-%���b�3H
> �/Dt�j4!۸�F�JR�K�)��օ����IJ^{j��"!Hg
a�y�9L�v�l�zz~/S�0<�9�����ffb�:hg9'�Uj_����Q��&��^&���;��z^��(hV�3MySa37�Ʀ3G
ra�~.�!�����m��p�-���R+Z�V�����4},�%(x'��&�į�(�{�I��!%C�4���L��d�.":Y���L��օ����IJ^y~�绂� ��obʠ��jLZ�b��Z��p���DiDZ;��%�
d%����!]�����s�qO��fA
x;?z��ş�!��糳�GǇ���oN�>>��D�>h��������٣���f�2�3j�����U>� ���J�	(�bA�$��3�H|}b��:}�ǃ$��[ju�Υǔ�JqkB�S�I��i��a�K��������RLS�YDR;ˈ�u�yb�v'�,58���'���=��l�mԚ�cq�7� �Y]3e�%�9�+�������#�߶���s3�\�k;c.l�D�z�C�j���v ����؋y���9
T̉�'ڔ{�Ξ�C�H'~��"�▮PI�\����"	g3p�ћ%>pZ��l:p����rlд��g�����Ds �6�"UX����Q������$N�@}��;��ೆ�(��t�/p�s0R�G]�Tr'ʱ1jՋ�+��
���Y���T�n<�)N-h[�:i����a��%�&���$�7F��|��aD9�tܽ��-M<�
y-����a�Ŧ�X&��)"
�(��%�ڦ�)NsI4�g�;:N'����l�}u���Y���(��,�	�Rg�B�ڃ�قϦI�%�۶�&��d�z�-�ϟ8�T�8�h[�q)J�i��`�up�U֒H@�GK$X����"����_�C�C��
𴣸@P����O��!�x�촆&L�[��q0����$�����S"-&iN���e��͔58��b9���||š?$"�ɈP�B�8���u+3�3�陉E��3DQf3,g�SkZ�qN%)Z�������갊T��*�ϊp���\���K�'�(@��&�i�+���Iy\Uq6�8�o�1V��̺�0�0a����͎}�l��ه'㦃��k�6��A���4�]v����q7b��a�c��&L��i�(h��}��f�Q�Kg9��_D<R@H���0=��x���fhA��1�f2H�2`Όf�0c���y
(Ґ�)JuHR��JR�H�X�tb�2I$��cC���<�6�q�R��4���1�2I ����2�YF� `�ad�0`�&,��Zֵ�˫(���2�:�#0c�1�0c�1�52���)�)N��)-!�T�2R��<�u�T��ZԲֵ��(�)�)L�JR��<��c4c��3	#8vn��*n2X��i�ȋ1\v��V�e�����"��b�y+D'���Z]���b���9�;~�f�cs���(�gf�dYjĉ�RZ�'�_fg`tV?�X�V�]ٕ�_��5�'�����a�bet����~p��TX�F���o^��?j[�m�c��if���et��Ź��V)3;����o�v�Q5�E폳������5��Ć/#��yߎKv�"��,��\���(-���8ϟ�~�*m������G�L���JU$��Z윗��m;7��)UѼ�x(UO��+�-fEt[���>n�nk�q�q��v)��; ���;��Z��5=���BA���BMrv}ss0{���OHMk���3�wF���dU�8���&.0j���\�]�L������L���]Z���i�[,UG	�]65�-1p�8f��)q�ٺ;e#�%���g���e���T2ˌ"��Bm�Z�nEF�R�[m%�K�v�����+�%�ҳG5�m4ͬ��-3���״&o�]�x����,H�1�u���,��&�v�%�.���B�\I�ͦ%W�﻾w����m��&߽�{޶�m��߽�{޶�uUWUW[k[�yխJmk[.(馚xc4�?%��<�3ԥL��ִ��[1�k-��d)�-����n�+��Va�b`�v��
$)a[n��:�4�k���#^&-��,�lG\��X�3MUk��KI��H�����bҍ!5�@���.u���s6��
ː��W6;]c6�Y��[����eb���UDK����_�b�����[����M0M8P��-��n�yV(DD�ΔIDГ ^(:x�syf L�t�N0G�/�Օ��⏐���%�-��+�gԷ�݁F� '��Tn���D�zY�t��5�S=3�ū�����qDД嚺D;#���J쏅V�S-�e���˨[M@Q)�*�;h�4#�K=�H:af��T�)��l�ڒ��JK�<w��o�TC��h��x\����i�9��ϟ{j�����I��h��U��(�y��m�[�V�(��}2x'SB�M�2^�f�4��͠�\�D�יTkG�M��҉�I���T�ٳ��8H���/rFP"��I$�"�QgN�H(��a�ጣŭ��R��IK�/�F#z��ʨ�m~�[�����G��Z��[O-wR�JO(�O~8Y��0ÂSgJ9D�a�|����,�R&D�㩧�8����8}9�4Hx�<��P��Z�<�bl\��N'gG㒉��H$՜�����2�dGB�`Pj1�6�a-���uiy�-Jmk[.)ĥ+R���C�'����v�"����n	������`�!�]���*�4�/��ߚc�����V�]#cjĢ�%��:���=ʿX�$B,hP"��:iz):#���"҅%�P�@���)��
��BϊQ���tng �uu�K�6@�h��#DiD�|��* �K�+�Q\��\��$te�1�,��J��R��ֶ\S�JV�<�����l:�i���)�Z0��i��k|A�c0��Uw��^�M亼ޚ�Kp �[�q��&���V�M[3
<W$F��r,�tKn�c�[�eV1�f�+�+X�b�f� �������'�~����ܗfp���Z��l>�jqѵ�x�ܒ�Ι3��t���ՊX�0P�]�z��A#�H�P�p'�2�D�m�G���p�\0Џ��tgq��ܼ<{�CQ��x��'���vber��x&	����o��������Q)�~?|����-����q|�]WXgB�(�Ձ��3c��,���&�j�;uث�p���PQ��%p�\;ԑ�(��.(�w�t�O�3uO��ֵ��JR�)��{�Ub ���p�e���8&�o��+�E茮ihT2y�4P�.�U�6Q?%���?&	�������x�������I ���[�%�HԈJ��_�y�u���<"l�$i6"h��^3��rͺ�R�֗�R^�!F�(�:YR_$�"0�3N�uKyjSKZ�q.%)Z��^y,`�0�``����!r�t����DO4����R
|��W�"]614'�շ��0�0�G�����թ4,��G��{X�Z�ԅUފ����p�zQ��pX<j�{�E�x�� B<B��ό(Y�$��s���\��g�RtO�OL>���+���8i�q�!�6�����Ԧ����\JR�)��X�cC�&�U��'�O��8'g��|�|���x��G`Z�d��$Q�Ҕi�QI�5~P��P��ΊAC,�k!!G�v�X�� �i!�ݙ���J0�{�DA&
!��lDOnM�E���g6z7��x{��H�a��(�dæW�D+V��I�����i�V�V��)M-keĸi���4��/D�^�!���).eO���mq��1��	#h�cr�h� �y����k3/�Ɏ�2k22����I��.�bj�c���86��� �����~�i>q����=.I*�u���S�ތm<|�=F�[�F������^��Qo����M~Bŋ�7���}=�6'�cN�x}���i1��q�8��n�Uh�Fq1Gl��~�(�΂x&��g�:�K��I��]Y���t^3��D0�}3��Q4$-B����7+�6r��N� ba�X����/!0��N��"t�y�	4�ũ/>R�Z�ˉq)Jԧ������C�V"lO��6S�/�����Wba(��za���f��=��®_�@�=�6V����F�X�i`}=04&���uM_5��f����0��m����e��Z|!��L󇌶��g�JhKPR� ��М��4d�S�;���n�K����ǝZЦԥ)N%C c,��2L:3`�3b`��21���223�Ό��3��IEP�1��T�)�)JJ�q�q�Ԥ)�(҉R���L��)��Ӧ�Q�H3L,�Fc c$�Z�Zֵ��VYM)JSJ1�1��c$c���dc0c a�2F1�33I:!�c$b�a�I��2�1�0�)JR�Yk[kZ�Zԥ)O0cΌc�fV@�.,�#T~�;���`�%���*�{�*�֧+���,�~ۯSz+�j3
���3���k�SG��^���o��>g�������r��at���ਲ਼Z+Ck#Ӕ�4�f\*e�q(���*�_(6k��UDV��(��pX�����ۅ0��;s��)[$"��k2��DynEMϫ�:��m����{����m��~o����{m�ߛ�B�Z�ukyjSJZ��R�R�)��j"#���jf3��F:��GN�N���:#K �iF	�j�-�F��0�YJB��4q�<+�5�G��as�),�h�7�Gi+NA�Ω�����"p�Dd	><0�-/���6&���K���i(e)x��!f][��R���	�l��㒐��/QaB$�>��JRַT��)M)kC�K��xc0�L2};>I.�J<Eɜ��|:=�!����DD���/z���6���ڕ�X"�S��qO|O'4!�k��S1&B�͜<��BG�}�Ы�k_a�L$��\��}�Y���!E٢oc(��tN��w����L�����&ũ}\H���2MqN��ϔʔ��ĥ�jS�^][Ry�Ë[X,0`s ���)�cA�M�p�&�'0e�X��0J�,Vh�sTۧ[�TMQݬ�M�|�N0�1�DD�s���%M�n��ő���X�1���N�%jIx�ዠ]�L�;J��Ի[j�,A+r�������}{��뉟a�tD�ʦ!T*�T��㎺I�+���fX��{mv���=G|~i�C����x���L"3�D-q�}���3����B��y�9��Ţ8=�M���Κ�O��/N|4����e����׎�	�n`��o�����)_z�6��$C����cmi
ךĤ��@�NLh���/��<��J�[N��[ϔʔ��ĥ���a��Y�B<�\>�0�[�m�Ȉ�C�4���U��x�-�����2�����~4Y���.���[yE���s�ѱ|2�{��$׳�����g�����w�<T�CP�4sgu�oÎD��Z�ӥ�HA�w�'�҆�j��А�ؒ6���J#���d��>S�[�
S�ĥ�jS�yu(�������O`|a���RQ���;�J+���B������?s���p�>ق$K��O��X�r�X�v7YU�x�E�fat����X	�����*e9��g1h|O�RjkK�4O�W�f=��76~7��b"'��݂͓'�>�2��ukqN�kR�Rև�4��a��yIk���K��Z���K���B
����$r�t_[j���{%�$��R��1yy}�������̢�$C�C�ͫфN8Ǣ<�n��e(dO�|�?~�t���Rk��z~<8tF�ܣ\A��5�㧌< X����s®x�A�<��� ����<����<4���V��E)ku���jS����x��}͹[P�3s���ʡbU�-�呵J'��a��ef�:\ݵ��QtYQ��%Q(,P���քbz��y�4�PNo�'���8)>+����g�W�0��.jWc+��'�L��ġU�~-�0Q�,�	a�i<;��T�a����N%6�n��k�Ч�G��:��:'��ܦ��u|���v&����#������6�Q5�����L�9�"�a�:�~�;�+e�R��S3D)H�Yq��O�f�5J�m���ӆ�k��Ġˌ��ƈ!-�RT�ԕ��-n�����JyIy���u�>����Óg�4���g2���2���A�i �	�2&d1�e�I�8~��ke�-�|~V�OO|�~�'S_rT��j|�\�=�m�m�y)4�l�*����R�}�jt0�P�0䦸)���<��y4f}�2����D�(���[RR꒗�)K[��/%+Sӧ��D�gP3,�T����-/��X�%EX��ʣϕafO����'~T��4�����DfltY���-�Cxt3{���f��t~4xnp7�֟�ֳ�Y:����%WM�&�����!��E�"C1�y�}iƾE����cmN4��Dd\�U��UK?cL C9��b�%���fI�k�%-ze-�yo6��ujJ�R��Pi�i��a�R%��努�KS�%�{,�9�u`y絨���ӎr�B�9 F|��-v�zeH��[N�*˔�%(����$f9���J�O���1Gq��p}��3�UҖX�hO:t��N`Y�)=z�:y�H���>��ݟs��������M)e{*+*��fٶ�Ç��!��+?>w9����ߙ����;�R������,#���H|k��D����T ,"�A��D�DY-�-,�,��	�[kD�dME��-�kdE�",DE�"&�h�e�������ml��,���e�H���"Ț&�h��d[D�dB&�h�,��B,���&��""h��L��"h��&DȈ��6�"mE���-�MDD�mD�2-l�"�H�Z-�Z�!hH�%��5�H�"D���4B&�B�e�H�,�,D�dMl��-D"Ȉ�%���$H���!dkD��D�&�dk!"�5�h�DH�M�""�ȉ�E�hY�dH�"E�D�[$,�dHY�YА�E�"�4[D�4Y	���"h�M-����D���4Y	���BE�DE�H��8�p��"h�b",��l���"DE�4F�l�D[DDE�H�$E�Ȉ�DH�$[D��Y-����$K$�,�I-��I���-�Ki$K$��I,�,�D���X�IbkI-��X�D��M-���$��4�4�M-�$KkH�Kim&�,H�m"M-���	4��i�4��"[I�D�M,�&��$KkKi%��D�D�Ŵ�D�M"Y"L��&�[H�I�K$�,Y"[K%��%�,D��&�$$K$I����g���$K$K��K$�%�$K$��"Y"BY"D�E���$Ki4�2D�$K%���!,H��D�[H�$H��&�&I�Ki%�"X�"[I�K$H�bD�m&�X��$�ĉ%�D��9F�-"Ii$��K�D�Y-$�-&�H�-�K$�m"D�I�,[K$�-��-��X��i%���d�YbI��I��4�Ybi%���Œ$Ki�4�Mb%��4�M&H�-���H��$�$H��"I�$�-�M�Ȣ��E,Ef�#,F����6����8B[m�km��ְK�f�[m-�����!�����x�KkM���i��Dac�,��"$������ŢС"ȑh���������H��>6ܲ"--����Ɖ
�!h�ˍ�"�Y	���,p�"E�"!h�m�$Y�hN\��mЈ�&�YŎ��MBD� �PӬ2dA"��ȑdK8��-D�����ۄ,�B�"E�Gn2-E�"kmdB-D�"""��E�h�Z"&�DD��DD�D""Ȉ�e���+pDH�-�E�ȋh���$MD���#��"$[D"Ȉ��-��",���h���dH�"",���Y�"h�",����DE�H��D�b&��Y"Ț-�"E�B-l��dM��"D�e�E�i�D�""��m�"�,�MD"�"!"h��4B&DE���-�h���M"h�"!�4[[&��Ț,����DE�dMDDDE�e�4[DDE�2,����"h��""-�h�"��DD[DE�DDYl�",��E��������4MD�4[DD"kdE�4[DDE���dMBh�"9s㔭��""h�DD[D�ɢ�"&�4Yl��h���"e�h�$L���h�D[[&��h�"-�h��l��DE�4DY-�D�dL��h��,["&�"4[D�4Y["-&�Bh�-l�-	��DM�5�Y����2""",D�m�4E��4[DDE�m["",DD"dDB-��E�4Y�"D�ȋh�,D�d[D�4X�DB,��"Ȉ�dE�"Ț&�h��DD[-�"�Y�ml�-�"h������b"&�h�",���!DE�mDE�dD�m�m�ȋ4[DD�dDDL�DMDD"�&�h���Ȉ���4M��E�m""h��DM�4YDE�DE��DDYD�mE��#��b",DD�ml��DDE�MLDD[DDp��dE�"dD[D�m-�E��"&���"h�,��"e�h�,���"&�"h�e�DD[D�m�ɢ�-�"Ț-��&�ɢ�&��"h���h�Z$Y$Z%�Б4j$Z ��8�q���=�{�/�9�7>���=����с��2F�3%�T��ǌ�ї����wu�ݽ>��{3����������t8|����{������u��q�nm��Ni����]�܏���^��v���\�s'�r�9�os����w�v�2�_���t<����w���烇��6پ���<�W����w�3�rm�l<Xٍ�H��|I�6ٿ�q2�K5�7�}����\�p�ǥ�c���K,�˖�l�����M�OS��|w�֝!�g���3f�4{3������D�׫9��mɽ�xfz�~�t7�ރ�nMlY�Y�gs?��Y�q�~v~�9��q��׳�]��ϳ=8�ǣ�{9m�9Κ�kVV���q�vy}.3����q�0n';�3q��E�ln[�86m���M��i��K1���i��36��:8����#����3�G����WG3to/s�ϱ�n���<[lln��D���c
%�Q-���6ͩ�f�D��˓��c�o��x3�n��u�7��fE��g�ޭ�7����;a����O�����}����u��vBm�m����N�CӾ���uv���~v�}�������7S�~��s7�G��-����u�s?c9�Ŗߵ�ON��g�};�<>[����S|�6m�zq���~߇�h������8�;�����}'��8��ޮ� I��f�7�=��s-���ίͦ|��-��#�<?kr<ۦ�ý���N���p��y�ͳ�雏Z+-KŹi��sm7�9��lF�C��=m�f����Mn��tnMq�5��c�����]��t�n{��'(��o�v��9&wi]#�����m�n6:���T�?��}O,æ۷��6ٿ/���]s~��Gמ��6��[�&=��~��������g�rɜ�x�=n\��;��z��|����M��ۏ�9d��o��F�y���y�m�y�3�dM���~���͛lݍ�u>G������;�so����=/K<�9��~/�sg��;��v�Oo����[�ӟ�9��o�r8}���C���}>��G#���}���uξ,�ܝ͹w�{ή�ٶ�e~[��ͷ�]��\p�=���f�o��rg�ky�oSw��<]ۻ<sw�1�p������;�<����oG�z�������ϳr�0�=L���g���f힓�����oI�s���|�7u|�uu�87��:wà��7�+O�88�F��Lv������H�
��݀