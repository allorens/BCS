BZh91AY&SY�:)��߀Rq���"� ����bH�|     �S�`1�����֍���6�hj����U��l�	j���@cZm�֭�m�c[�A�f�J��Օ�l_N�� =ym2��dj6��6��Vڪ��cmMl�22Y���ֶ+��mA��Q&[kmYb����U3f�ֶ5*��i&�mleJ4f����h�m��޷����m6�幵5�UL�W�c�=kZX˼�y��͖�#&ٴ�V&���[Uֈkhj&���l�mX�kkJ�Yc��kB�m�^   \����յ�cU�V��h.�N�+�H�*�vi\�:iӪ։]��U:h5�`��wY�V[v���l��kU�#a͘��f���lm��'�   � ( �ޕ��ۣ�z�{�B�
oK�8�
��J4�ӛ�p�(*b��U c��Mw&h(Phonzj�D����Q�ʚ��-�I�   �'֒�����tl��K ��v�MP�����A�
Gz���-���=	5^�w�O��x�7_`6�g������Vͦ�EQ_   ww�9P(<�w����kA����
}}B���>�}4(
�����R��s��@(O�G�}�
���>p�
R�[�o��G���R�
x�{#Sm���D��5mh�   	����m�l1�/sC���w���iI�>�}>���W��@w�����ȥ�s��P�{�Wl���w��|��Wݱ���TW�;m��&eY��� ж�  ���ڀkM_|W�= >������(vQ���� w�l���Q}���Ҩ��ꛏ/�J�j�=կ��@S�y�T U��GF�)zN͊�ƤQ42ڵm@�6��   ���C�4)x�i�J�^x*��gz �ۻ���փ@=j�t((
w%� U\=�;P47�{� P{ݧ  ;:mi�5Ib�I���F�  ������p�t�B�;  s]�
�. 4ά� �c��˶� ҋ��P�����D�jR���R��
 ./ )��� ��� ���6� 껊:(:�� {�� �F���먠�ma�X�Y�1kT���J_  �x4Pѽ+  wN8 [��@��7L�@ �K@�ui@�iX 0"��;�  ( (UCS eJUM�14� �i�ɑ�C��i�R��F  h��S�&�%R� �  � ���J���      "i��Q)�jM4h�I���#� b4	%MG����OM G��F�4�2i��~/�&�������~]���/�yT�r�_.2�mV[̴+��r�tg9�{��H$����U����9�"�*x� ��"����ȓ������������������_����?��+���UW���U����!'�����
"�������G�o�?���W��?�����`O0���	���Ẃ��̯�^`0>d|�����G̯�p�\���<���<���� y�<�d0'�e<�9�<Ȟe0'�C̡�� sy�3y�<�e2'��	��+�& �y�<���<�d0�a0���y�<��a2��C�!�� y�9�2e0��̡�P�(y�<ʜ�`L��e|�e2�C�)�W�<��<ȞdO0'��)�� y�̌��a0'�C̉�T���|�a9�3y�9�<�d2���G�L��̡��"y�<`O0'�	�� ��<�e2�W̩�'�2��̩�A�*�e	�� ��S̢��_0�s
�AS0�>dE<ʠ��A� �� ���Qy�S�
�QO2��eA<�"y�A�()� 0�DG� 0��e<Ȋy����S� /�y��)�O0 >`E<�*y�T�*)�̢�2��L�"��U���̪��EO2��`D9�C̀`Q<�
y�D�"��U̪���y�<�0>`0��Ć�� y��+�̡����́�̯�_0��/�_2���W�̡�P� y�<�`O2�̞af@�(y�<Ȟ`O2'�̡��y�<Q A�����"Q�_?=)]�|���d�>�����%�*�eKU����%g
��r\��;t�oiu��;��@�q�,L�B<�(�ʖ���S=��I���Y��Յ�ۃ�d�p�Pvl���T���d	��G2�����c�'�b�˂
���U��pKp���8�mC�\	���ZA����E��t�_�Y[H���jxky�|�d�
��5]&� �	� �1:���V�w+w7�8�X�>�ixu@ga�Μ(�i@�=Fk��&���1��/}t��<��&�WC���er�+ǽ��dsi$Ĝyۭ��a��]ܓD6�$�,���fk�a��/1�˱�Yc�uצ�L9��CilM{cx�#�&S�֔6�;m8ژ+�����'�a�s�iiL+��L�w���O}��R�Ϫ�+++�n��U;8a�n�,�\�,����ҵ��mG�!ST��Y"��"2�z��|�b������Vn��zBНݝG%L3�O[�݇UE�#E��5�i��@j��u�8J1�{�v�gM�xk��+T��|0�ػ�6t´ �fP�:|Z�N��j�	߼���ݤ"�:�-Mf�^��sEkB]�B�)�m�V&o�،�i�J]�"�2�iŊ���gt�*�R���TDYK;�f(��f+������q $�״���cyn(O�p�	&^3�U�	q����yݔ����݇2c�Jɦ��B�Rx.�^���$/��/���{7A��i�H%�`ǧ�܈���$�v�!�8�zE�#�A��n��wz.؂0�A�K5�LrPJ;�Jɴ���:;����~u���PoXX��բ�c�b`Ŵ��@;�{���T2���w�L�(l�a�ڪ�r5�^f �d�K���]&��<�o�:��\�+T�W$t�܃�a}g��V���Ӊb����19����r���Ha="5q�VPw�ƌݎ��nk��ScV��21��fJn,�k�tgu��q���#;t�ΰGλt��W\.ƀ�!t�"�������?�:2X��3ToV�>��'$�n�.��e�CǛgk.Fe�jr�[�p��X���67RX�˟k�";��ꨉ��{�"��\L�u,�z�"��@��׎���� �|�x�b�ywb�/����c�j�Vi���jFr�e	����M�Ntc�$�6owB������7^��Źv[К�-�ZX�{���I�Y�0@7�F3�sᑅ�vNvML�f�xbgztx7�
�^�J}��R@Z��WlA�8OD�]�#���r�8�h`�^�-p�&�v�5�e5�s�ɍU����bަ���v�Ƿ��ovmX�v1��n�]�YG- x!l�]�߃��ɒ�CΤoi�t-�hK���_��V�<�+��J���EfU룅��Cv��{�T���'-:[��l�:[!k�Cx��.���q�/.r���p����2:�ś]��0��h�#5ݢ�f!��f�]��h	l��z�0%X�rZ{�(ĨG�(t"�*��ǄE+���*��H�Ryܭ+O����H��fC�)�k(���v��av�x`�c�1�C������vC6v���:<㓻����s0Ql�r��R�ףFSE�-Tv�i5��;-�5,�9���}��Ж�.����I�V�~ڲsZ��G!`�f���s3F�6A��M׳F��x�����Jv�1�����#Y_C͉�p����AUӺ�N�pRc4�A��cfHW"�0wt���u;z��@�H��J��Кy��Ӂ��%���yc�ʢnQ�ҫ|^0�Oy�.��<h�dl���7Jb�/2P�T�@�B[<���d�ū$_�T8�N�YOj��;u`g5�[�5`5���V$��|��xu�2��y����NEjouAޖ����z���xƍ�u~z߽��%Jc�
hV���M!��-��Y�0-�f�ŹĢ�>�>�٪H,:���,s(����0<lf^$��F��ȭ������^��_[�m�q�)ǆa|d���[Roh,�ZJ��M;(�/I3	�oQP��&�ƺA2#y��>��i�/=�����30�X�V�]챧cܕ2�����������Ԟƹ��fn� �vc�ΰ=�L@fw�`:,�IWQ�͹�fY���8�������5vͣ{�xq��$�ރ:.����;s`m�Mlݳ��K��b�f�bI�Z� �2�m�n!݄C�&�^�cȆ�~����(.����S�s�^�	MG��M퉸J	l}�:�C����"ԗ�R읐��+���y�C�s`1�7�7��.72bO��O&k���bS����5	^w�:�P;')��,����\�+��	��WA�Q������H�TJ�첆Zjն�^<�����D哲�Mgad�W]��)��^$��2�؎l F���Y�O�y۷�L<�:4�Z���/����V��ł�][�#�k<N�Ѯ��j\��~2kj)[o%��O��9tj0����dx��dK��p�S�r�)�cDҚ���������7FwΪ�;su�����jG.+���kS�J.u�V[�8I�W:]��#v��2��^IL#5��gH���X�5o��8�͍��n�!�Zi��f*��@��kb�:g���c�a�e�/���	8��5���8�9��{RIz�˺�T䓖��
K}�P�Oj�#:'����c��p*U��;��x<X^v�}Ж�Y
���l�����E��*��\�ok>��oӼ�Ш�W�4��^W���--��e9ۚflQ
엨0���V�X�B��Z�i��X��(UؤF¯G�k���"��&]Po�5�N����sRD�.ȣk�����'��lΑby� �:�L�zt�x5�������C�W^ ����Zz��4�����\�����GG<��nMë�<0��0dZAmGuw:��2���/dgj���S�J!`����#SGpF�!�B��7��7�]�3b�]�y��t�w�V��d�Yk8�OF�����mۺ:�C�.�*V�.�k�{��O��[�l��p�v�N��	�)u�v�y��9[���1���EB��8փ�ʋ}�+Xƽg�m4}�f�$�x4�$een��Ѫ�!.r"����=9׎w�I�x����:�����
�i����(@y�U��W�۽�f�g-!'�Ɵ��b�~��׼1�K��5�pP��_8�Qe)��tH��z7�r�kӭ�P+�iژ�7�FX̤��uø2d�u�5fs�%;*���}e��,m&k�J�ls�A���}7$�+8`�E����r-�#-qNlL|�{�+����T�:�9wn�gIɨ�WE��{�
�ܲ��D��3<4�zI�q��P�j�kJ|��Q�T�sz豝��CcFkX�-�J�����2N~tq�D��b���1ʣ��#̼�v�ko,aL�c5��D3Z�n���.]�,�G:R�T�i��zވzS�OkoNV��m)p�,[\|Y{�Lsd��DA^��V��3oQ�p�{���W��4<4ڕ��vw�:C�ovlX�w)�����P0����#z���G�t���=�@W�D~4�����.��`�HL���e���a� �n�դUP\��UB�t���/7����f�ͭ�;���v��և��,1Bf͟�Xm��972I�ŝܷf�^�Ω�+CpGخ��v��c| ����Z�$�z�'݋�s�k&�Q����M��A {��r�k'�B�2��o�"=h==06�_r�KGI����)����4S���;T�7*�E���.Z�U����7hԦ;�q'����͎���

^��qd�9�q�n�ۺ;��*�v�XF��A��Y5k�6��j��̚`���lA�J����sFt( �83�#�i��jw��+�N;����W��4��N�������4��F�Dq��k(���h����cI�A�i:���	,��y1Lل��^���n��`�WvS^��J��@"�Kҍu7m��V�'�.�N�Ir'�[�df����Y�ѧ+��MZ� �]e�i�XZOK�صp��W�e���P����V,��p;��T͚@#7R����cE�#��yq�>x5�ַ�i	�ǧ��9Gb	Vu^ix4�fA��ۭ�\HB�����j�d	�;�����  :�?.�A�&�sC0.��L&`�6�H���'`k$���P��W&o͝!�oF<K�M>Y��� Z-��������C0��-㶮̺��JnLűx���Pх�t�F6d��k�r�ث���^o�:]��1�W�,2)D �����&�x^��)Ō�I��c�jo1��#WŦ�$&n���~���
kG,�Va���6UnFf4�R�2�Z	C(K���ѕ��lXp�T1�Gl����vA���mIr5�����Cc#��]���K��R��+6�����v���Mm��h���y��3�F1)����(����ww<��	�׈ø��p�¶�;��x��9�xu�:�ǅ�­G����T�<�M��$D�-�yFC�v��b��ݜ�/s��Yt*d��֋�z�Fa���Ę5<xsF-Ѭ�!�n'��H��ІXи���iRVP����O�˲�*�&o1u�X����OR��óTG^�Oz��+&�����L
�0�%�[F���0��)4౭�3B�u#ҭ�:���ׄt�6�I�[&=M�$F>K\ٰ�ݪEyciv�tn��ECHm�b�Z��5���g��kg(D7M��j���
L��d�9F���m�3m�����r�+��|OZ�zk)�=����������� K��v�b�נ��V� ��nU#� ����1V��摮͊x�f�,�FE*�&9��bm�镖6�.d)E��\�.78w\w�4����:x�&u�]Ǵ�����z;NI���_%�
��{6��٬í�̓��u��mN���3���M����L?�-�ݶV�����u��:N�5Y3U��̤�7S��1���%�2��+5�����<;%��M�k׻R�1���^`21$�aL]�#U;%jV���f택xl뽁�r}���wwF�q�2.�f1��-��FRAOa�dP�Zy&&T��D�B��X���������읯K8����SÌ.�r:�I��W�w7[`㙥�,y�[y֩�7��q!�qT�|{��S��p,���M��W|��ПVS�a�G(P:)Kb�j�i�	���!�a����:q���Z�d�N�'[��d��Q����
���K���c�@'��������$��..�4e����Iv��s��&������[�,�Gv��M�Q��*�p���T�n�wM���N��Ú0�J������h�9�T��1��{L���0�)�]ƪe[��v�����@��B�(=�zvI&u��>ߧ-E^�kA5��V�iAp�d��N��Uv�t�M��q�k{��5�+�Uͧr'6�$K��NY����B��
+((>p�w#�)t��3�ۢ�Wd<qlF����Uv�5�\�͌K��&�j�>s��Z��ħ*�r�eTI��'�2���)�j�)8��)qi@Ƀ�CsOEj�bҗm�p���F:d;c!�KkC-��K۵h�6f�՘
���
4-���j�h�Z2K� �c�d�rmg4�6�D���ɥ	�sֺsF*u��0�TH-��n쮚*^��+u3����V)ïn����4M͆:9{R��Va4�eI��-g.����Eȑi�آ64�5�`\3��2V����� ��]���ĿJ�B`�b�$�Ӵ6Y�`���m��Q͗�\�8h�����&��U+ق��2,���ս�n^��V,r��]̫zG��u��C]0�P�
��n�ֻ��@�;v>l�9��ñP�ݧ�O9E���D��r=��dѧ�q᙮�Sn�v�橙����L��ㆩ�x4cݳZЪ��6U��bj� ov�k*Exy�$���S��V��$û�6�;�����-g #�w�NN����Fn�0��i�n��v�⚕d6�j���-CDn�(�5P�f�H-C_n��y+��X^3f0r�l	�/v�ެN�A�j�s����+���l�4��S.3 ���L�Su�`�Gr�}b���x1���\"�@�93�i ��&�Q�K���n�192�{^9�-����8�h��+x{f�GjɑÁm�z�{7V6v!�wE8��W���Z&>�C8�u�poU`SlJ��l9�&��N���>�F���F��Ф.�! ��t'i� 7�Az�6/q���_:��Od9�6��^b�nl2pR����*r��
��g[�ׁVv�p�k�Eqe>���8�{�y��DQ�	Lڑ��b�B<�\�;�~zy�I��B"X�-�ff�Nz��ZR��dy�6ȼ9@���&��x"1���]�;$AW�0 <��<�s��À�(l�έi%{ae��Ѡl��oyr�(�"�BU؅�jLd��s��v ��x��,���V,@��_D�������6i �i�a$Vf�j>?,o*��;!�Ҩ��R�s\���:��Z�{.���/�>��E+�pi�0���W���J���9�|5�r��۴�;�_Ɵ!�Ƨ��T�?���;�^y��}�{z���(�0��c��m��s4����u��[�h���޻�t��Ds7�r(�`����wea�n�o%��s��=��L��<$�H������_]D:�g;��a����ac�zVʝ�����	W�k%��@�k1'/��z�yv0��tm�Q��O�%;�ր��p��������r�]%�U+�ڥ�TPs������U���I:����Ycm��)($�dZ�u��[����Y�̭���E5y9Z{ƽ��=Z��b��(����{7r=+]��%}�y+Ke����JUp�[ev�VD:����`\`��&+#R#Fܮ.i@�܍�7�����vr�������������A�waG7��s||b�{!���!7�q�i�u�%E����(������K����;��a^��I��7�]�(AG�����pX���;6������ �E���^�+FR;�y|Q{�`�)����E]+��L͂p%en+Y�n�����l��t�n��ܣWw:���"�Z�)Lͻg"՛t�&+���q�6�Fd9��(dV��YU�+��"���b̀��#�H\<_f�&�����[�ogma����s=��U��<�l$���<��K3���oi�Ļ˴l�1b�Ԙ�U���2�;-�Ѻ�D]��f�Ybq��sd�(7������vn`c��b�٫N]X��
�]h)�5iKj:�A&./�N+����s2�����7�3Q�������.�'���N�U�v����?xj�����P=��U6��:��M���5��ȭ"P���G''i�OVvZ�k��N�)�e-xi���p���Z��-c�Cn8i=W':���"Û�:��8ݍK�L9�}�D4��B�:�sU��#�f�'VduX.�R�wd'�,��9�L��mK�g��Q��ڰh�,ܸOuof�
����Nhg�����.�:d��dI�M.�^��5�V.V#vt��w]�����i��ȋ�fR����xJO�2�Ջ;
_m���4�&�	5@gs!��qQ6�Ǿ���v:c���;ؽ�/%��^mp *�d��.�#]���Vj�{5ÒO?{��������p�av��w��PsY�\'J�ح�3���m|U0�u��+[��g@�I�mBj*푦͓r�q6D3/i3-�b��!���Ywn oz{��L؞@��I^�c������7d�BEM�9h�/rwnպ�LqSv��2nuEq�?YeQ}W��QX^6g�zs�J#3��C�G_,bW���I4I�+e�
�Ǚ�'����H��+N�2���"Y�a�W��7�|8M~���5�E�Z7�����ׇ��r�q�cJg����<���5�=�
�����U׺��ҹ�V�寴�_:9!�<��)SC�jF��C��؎\�Z���S���~����A��x�i+�v�YB��6�W��}��]\d�Ƌ'kF� ^-���w�-�W����]���l�G*	�,�]-�3�io&���r����{�Zۓg �l�w�p����wʜ��-��H�M���� �$}���.#6�hzz� x:��ט5��/1$���K�
�Q�2�̴���}"�OS�]�	�D��t����1�SOܒ�ޜ�=9�4��N�w+"��ֺ�*���+��Y�5e�#I�%���������:u�{�h�ѹA�X��:�:ڠ6V�8$z2Y.���g0k�ې'�nm;�X�p
NQ<��qy�bt'Et$�F;��.��� ��ۘ�o7-6��b�¢�����Js����+���vjֳS;�,L�j�^��7FJ[�3mK�����n��2s��D�$��T��.�ĕ���Ü�&[�Z��˝ڍQ.m�n�K�w&(����*G.�s��
A�7�)���{#,E]�;�8�N��q�6�V�ں�+����GS;P5aG�1�,os�ٰA�<n�X�֍ob0٩�8�^�ٍf�yk�h�z^j$	�ܮw�x?@i�Ӓ�K>:�{7�7�/y 6��w2v���~x�A�������_2�ͫ=ڄ��-�6'nW*Ψݸ�>�땪��*�*V�]�v�\�G
:T���7e��E\;� �qB�Cη0!�o��:g����H�n������5��]n��nb��t[��5v��V��j'h��l����.�u��n�ۺqpD����rb�]��i�wVa��kV0��ު�dVk�bn�:���*�Gm� �v4�g�;�Ӣ�J�m�ܵ��'�2�kR���`yAg�6�͡���B�LԖp���a�:z��u>琙<�܇$y�1��	ܧ���rn�c�
"���rj6��^h��n��m՚�tR󈀼�f�ף�g
<Ͻ||�v��u��^}	���tru�/#�2+�֜"���\���wo��i>A���s+�%�*٫��:Ċ��gB�C��V3��%ɻvŸ9pu�=�H�������+����q�ua/L�N�ˆ�)�PYiu;�[L]2��d�x�ˣ�J`a-޾?���-����kN�35�B�f��"39�J���.s�a%��Y��WA����NF���ٺWcY'e��L�];]u�Y��$^p��3C�"G���M��w ��4�1ol�J����񳳟��u�܆hK�(���]�sB�uf�'iQ� �W�y���:e5�O�P�����0ӻ�Ի����%��-l�d�i2�`{�VR�ʹ-: �]�{�2��++4��ff�Z�&:�Nvm	��_��W抭�"����u�EH�ʺ��y{��Gn�̬@�Z�azH�;r-���x�����\�5��ɪ�ѓrs�_���݃J�#�q��5�(��f�]�5׬Z�h�4��3o��i�Mb����L7���;#]\Y�����i���At�Y��멧<��x�76����O�j,�x��u�;k+kB\��^T`)nvNwʠ����VZ�.��"mPc0,5��t�w�s8coZ���������.��vnbUzlo��mu|.�'
���>�yVU������؞��Y��f�wv6�F�{q=�b��q�vz����|�e�	it��~2��{�����&$A�Ǆ%�b} �)h�b"������x �)�ىnfu��5��Fd�;B���;>Z����_s,>]�q��r/̍���,��Jv���V��լ',s�����Z�Ψ�hT��Q��G��=�F�<�,���E���h���oY���4��u0�8ܥ�G\��h��۔�?)��X�x(nIuҮn/�1���JNf��#�c�a����jMy{�8�e��;�*Iɫ���f�����=b�i}��s�3�����<Τٹ��{�o����Az���'���p�����@\o��!ɏtLٻElo��!#/,_XP��on���`Y���[%����;��@�Ks�JËz�	c�ce������l�n�n���f	j�������Z��J��PQ��#���1U�-g22�_iW��UҶ@�����ԩ$�����X�D�!�N�'.�a��oiU٦��� r�p�|d�gǽ�Qac�"�8v�I��}!�vCg������0�!�[�nI+z;9�O�ګk巍��j��7Ճe�S>�q�:H�c�X�[��Z=f����z�`Ɋ�g���ɰk86jr�����'oZsy]��5f�,��㊓�,8���h�����-[{�-���g��U0���t��+7�ș
��o{9vT�� �XR�170X�ŋ�Ig��!�W�t�1'�e^��U�^՞�k�tg����G��z��������9;��%�����p�=5f�*�LJ�-B�wiVqpZJN1�ON�(y Wg��ΰ[�8���^����p���Ӝ!;�,c�s�C�=l�o���k�^�|�K	�%cJ�چ�xsU\t�K	��_1!��k(|�嗄�/v���y���l�nv�l먈}�_;6�K�5J�7�������^j�s�-$�����ne2�D��jSw޶�{ՠ�{Z�x�M�X{�/������n�������/���+'��̐l�q��-T�C�|�bT�B{?��옰B�w���4�b���陸��y�xjOe�X뚟ݖ���k���n1�S9WI����,�4�r�n����U�pNW�_F���d��	��g3i᛼#��֊<Pe�/6��b�Qa�J�釸K�CQ��y1ji�����<�����������߆M���������]-soC�ocw�(��omǔ5���)ޭ�o�c�Ë�>��B�\�ڎu��.�Avk�_1*�ƴ�<F�pb���w��JP�Ӽ2�i�(��å ��je'u�kB�uN*`��0u��1��WL�w%�u�����F�b�3��rJ�6�;��N���X޵��\��6p��E�]��kT�nJ�c4���Uԙ���t�a�nJ�|��8�&�fe��P<z�C�4=/����>��C`�Tn�-7�T���c��n�Y�^���*�.Ƿ��X�a&��n^���U�E����ӱ�����y���Y2��-�"zN��>L�É\e����3�E�#��Ky��$�ף�泙�&�%�H�d����EN�m\�1w�$L����=K�/٣�(̬�yv���9v���^�1[�����P�:���$�#Z�t@�}z?��$��ջð�������Υ��=V"��R�Fe�i�',s���<���m�u�ei�T=�L+I���yW�73��9B�Y�'�
��zwӕ�ȕ�w���2��Y�ϼ{��`}�Ig�18c���u�p_�r�-eb���)��z(���$sY�;#��*�nH�`�]`���LFE[�m*K��,Ӑ@��s��<�x,өA�W��0g�Auy�^t��z�3�\�5i��s)>����x]hҝ.�H�zĻ�~+3�oUA~:��ǃ���%�|��Ϯ��wӒy(����QZx����ev6}X�,]Z��wNu&3��Jz����m��;���Ƅ�rl�F�-wf���u��O,�{{R�Iq����4�nwa�q���߹5�ŝi;u3<���o8.Il�3B���}�f�f��	�0���%ɞ�/��b���r̈�y�}h��{�Y��r�h헄ڹט^q�p(w3�j���X��g��߄�H�qI@��{�FL�����=˲ň���7��I:�����#�d����#��(n��Kz�v�,2W��N�Cf�D9��=����/dY��a�H<F�������	���p��~�[ށ�,n�nƩ`6��!�K���fӷݑn��/�9[դ]֍�(8 b��v�m�D�$���L�b.���VftG�0u#禒=iP����0}&-̽��;a�B�������J�^N�ӓ}������"�d�8�\��#Ǹ}�����51a�]�.jrZ�ɕՏi��h�fd�*��简#�!�+�!םw�R��f]²p�JWkDwƈ����:P�Xͣ�WKx�"�"���k��C���۱��m�7ô�1��������-���/��������wh�=LF�Dc���_�f�!(���]4�r����9�p�ё"�8���"�u%pր�:]���E��X��=wI� CI�k! �0Zռ	����6TC[ën<��h/WSOn�vKEݾ��K���7q^'��TӻX�nF���\B��O��{��ı�o����}�y��I�]�E�!����ծ���۷�G0�0p���[>��GL�E������]��S�Y��>n�+��뮍�|��3v�^��>~�����bq���(Ӣ[u�_ǖ�`AӔ�F��o`����Ԧ���ᇮ)Ǣ�_&00�9}�Pϳ�m�2Ӎ�蕷�>���`�A��:H.G���n�b�V�c�8b�NР����7�;�N�V�C�k{�Ӷ�n.:��Xv�uz�{}i����&2�hSx��c][̸i��go>
<c�]`�RT3���B�/&�:	,������"n���f�N���ބW�۽%7�c����SLl8��I
��w�ܵB$�P�`vZ�G��jWCyЮ��u�xC1�y����Ӊ�03+l��K��Y�b�wV#{nH�[��&��}%ŧ9�m�,W8"�qj�+j`��#�=Zim������y �l�S��.�K�������+0�� ���6�u�F-����N�h]s/��j� L�7%�MK�#IHY�B�b��Mf!f�y�fX�#bS՝���Zr��9���&8�6��-��T�ݿxd��k��z�h�{����!��!9���uaf�&��:����sT��\��Ĺ�t�͏�����r��}fWQbvG)Ft�7��]]�z��æ>ɍǬ�&ͦp��4��R��� :�Kۊ��2���E�?E2�=���ۡ�c�x6�SR�qt4���eh�5ɹY��"3V�g7%��z�r��}�{�pL�O���;��v�]�)*õ���B��R��Vg�g<�D&ml��w�z�u�n��L`���٪��[s�I������B���!�!l�KH��$�d�#��Ԉ��HX���S&��BO�(Y,&/�B����QFR?�B������E\����ĺ��%�ST�-�j _��D3��~ʈO�4���5��{�\[c�H�4�8��i-��f`���B�7L�QA
����)"��2"�I#�#EH�
r��ܑ\!6�,��0$�F� �?z���NjnA*�X���ǽ{�6Ǐ{]���	oG��?w��$�	 ��T>��=�� ���}@ A���G�>�����~_G����]�w\>�st�������Q/l�㗹������+��n��Z�{�����)t�g� >,�^������.T������j�;s�`���*{`�^ɭd�^�G{<{yz'�1M<e��jY`Ǯv6���Jq��:egG��6����2M�\��6���j���M�%���YG���0Jw3U�;{������3_j������xq7���mi/e�j�H�h j��K͊����v����5�5�V}�YY�EIl�_N��(�d�Q��S�xg �p�v��-b��t�K.�y�f����o�rt�p\��>T#�#�*��[�=Ɩ;'�.z��;�3nXs�E,SK4'�
ݽgm'Oo��w�CF��|�i�����3�GL��(<=�c]�_5����ÄY9�'�B@��b&�����U}��6t�C�KK��Ù`�DiB��v��wQ�m��^E�Q���l�w���H��Tږ1�ԡ{���Rs���#׏@5bĺR�b�s�<}۹<�kљ�Z�Al2bj�w��љ>f��ts��J�V.�V]gJղ�9o����ĈJv��(��,����z}�]t{�y�[��rFo�Kr������ZN���qI*�vە75H�4�m�&}����w�/W����(M����}��ӆM�88p�Ç88p�~�_����s���s��~�Y��~�_�����8p�Ç�=i�XV㝤�"�J8h;=�=�5�ps�&���M^`�/t�����
��|:��٦���?��qz|j{�>�q޹�}���'����ǜ��X����O���l�ꛕD{��!�m��\�%���NP�[��r��Jr�ˬpף��4O5ɓR����xy
�M��Lmћf��WN~m����8��DV���!5�+6"qͱ].MY��Qg`��pȻ3���z�2�
����{��)2u�� �6:��� �_ٙY��A�O�#�v��Z{a�X�t�]-
�%���)��P�k>���H1�Tw&n�ʑ���8�5+���墭<��]A������A����a�S��3,�Q�˝��Y��k�W3���R��F��g��+�ᵘ�mGo!��2��h���57�t9�Ŷ�	?c��%]���܅Phe<�x�H��!����VV^�3{mn-i\���m�Ws��̽��Y7C@f1�^)��Θ7�9�>���W�<�����	�K"���-V�9�6�F �eIh��L]|���}h��)�o���P�f��i�P���ւ:��N��~�ssW��w�@Ivzv�4�G�l��tŷf��������v��Rw�#9��w�p04bG�[�O2��K�4��uw�=��{�������}~���}��}����{�?_����~�Y��~�_��~�_��~�_�s�����~��~�_������~���~�_����{�]û{�?7Y;��,����׫O]�;%�m
s�[%ާ;��*��VJ�T��.5t|���M[��n�\�m�ru���զj̖zd�ЀǾE[�<�$��Y&y�,Ӳ9F1gp�{���}��mS���c����u��{��|U�>yǖ+�J:���hq%�(Zβ��Տw�.��
l�L���0�vei�nXX�Ka˸֚
���k=���	�gv(��A���ހ�h� ���?hΝ0[<��CIx����d+�t����G����Hi4I�%��ʅek��t�rU���D�1�}�>��G�*	Z����F��=JŔ)lR�M�����޺(0Dл)��n)c0���~��l+��{ԭ��Rwe�);4�Q�׆�͡C��Rd��Z����������QN�&u������ʜS�.o4��郀�&��#VS*^�:������[NLYx�~�؛�Ik��,�g���TGa�]��i�t4����5�*2Y0��2
��D�de�nV�k��ޝ�Ď��{�C*���-��������^M�����f!������+,ed�������U�D_u�V���t}5v��[h֍ꣲ�d�T��9y/&ޅ��a��՚��oq��`��F����k�s,�^���-�-a$k�!�f۬[������8l��g�8p�Ç�8d�Ç?_������~�Y��y���~�_�����p�ÆN8p��Ç2p�n�9���E�[I��W8H9�U
��X��S�-s_L����>;׃�;,�PӍ7�_M��tp����o\]ϖG���M��m�����4�'w�{
�>�}ϝ� �����/�{��,��"�!��py329�G�t���8��G�]f( kwg0�1�� !1�ʦ�#��%\��5�&����/rj�gah�5s�i�x����=]d\�*w�� �.A�{�	�U�J>��oV��� D�-Z8]�[x����|���9{X�d�-#�y���2_N;x{��7��"z���'�zf�r"�k/i��� Î��-�3�d
[��+��6S}}+�.����&�^>�5u�I���ʐvAGt�;0��j��x{���{���]	$��E��;^�J�u�����j���=5��O8�q�yhI�ĵy�� ��|h��ue�9��Xj,�c��EY�x��Ŧ�\*I}s�%5��ٲ�i��N��!0�L�*�П{6��F�3.A
w[+��R�wnU���s�4ʏ��:�6�{�v�tI<���J��SB�T4\ܻ�U��i�oATx'��bD���<�����k��(#��Y��G6�Rlp��O��6�hl�lzK1b{٪�ç�b�}�y�Å����B�w}�~��=�vgq��_cH�Q����8|���C��Z�{(Ge,G��X�0��i��r{�ѓg����6p��~�_����~���~�_�����~�_?_����<��~�_������O�럯�����~�U��|>l��1մwN�f��Ù�]tYqd��G�d�QLլ�����P�3��g���{Ǐ�DÙ��a��*So�>��τԑ<�T�5�x�P��+h��kH�+�ʳ����H��P�����Y�V�";9-M��QJ7'�-j� ʹ��X0H�i6gj˼ڑwQ����K��v����E�ٸp�ƙł�����1�1$�`���{9{�hmr�-�mE���c�˖�䆼��-����K6�wHl��,u�r-$Yo��)��0�[�@���
���/��B������.��.�8c�	Y#���}:���΀º�k+�R�9�u�σ�Z2�RJO>�*�s��F�7;G����	N}#_p:��y��w��S�����qd�q�gR�(Wȷ��MǍK�)a��*��e�c��@�8M[�R-M�6��N������X��B�W��w=P��X�e	,�Cz�n7VF�pTĢSL������Uf�'fj��*oS8è]�"��0��ʸ��!��Ʒ�L�*$�y/'��<q�m3��QW�~��_+�PɡI�������^K`Le�X�������S��kHA�U��s�N�44�����zM1T����q��2���^yh
�'�7S���<��b�}qn�j�7���}��c+�q�"��d�E��Ǯk7H�P�K�<�mM�;��`�|l�o����j��3�0�={��W�	a�`��y��Q՚��I�{V�v�׏��@�+�հ�d�)K˷%��%I��&L͡*+�uaL�0Q\X��A�+�{[O/���7�vk�$ܵԯ9hM�,�}�iUYVU�9�Q���ю�����Z�bv���xh�2�)�$_A�cK����wS�3t����\Vt��*�tH峝x��k29�]W �fo5�mCX��_W3QsC�,k��SYDɩ`B��#Ԏ�u�}��L�k�o�wܢ�$�՞3ԍ8���w���vы��>1&��J}�P�ק�^B��*��h��i���q�{[/4-]3�u9�8�b\�cwqb�X1�|�;�Gt���0�خ2�8Y·��U�-�|A*��؛�B����7��KC��J�5�+1A�����M��j��ڂ�EA����]���f�2K賵޷�;G!ʵc.�󁙝�4�1�4��	,�׎�,+��*��ŭ��ְn�L%&�yz�E:�$��U�Y�-#��B+ZF����:����+%�i�i�fsL�T��L��1�0���.j��h!�^��i���ύߛ[��OF�}M�n��B$0��<j�SƎeL���0G+[��tӭX��U{k�����b=��5�y���e���k-]O*s=}F˟l�n�۞�n�ve\eţ��ݝӃ��g9�X�$q�żb����毖Ǟ�>�C�7n[F��_%��ڦP4��4���rV��F�n<���IM	�&:I���/s�X2�2Ұ��-+�1�V����	 E����`ĉ��b�<���ɕ�����4����9/�M�����~9�3�-��=2�H�[i7����n�^�cq�9�nC����OdJ9��>;��k��\�~�2�j3�*�ؾ�n�.����:�5��u~�C�O��̒4���@�A��rJޭ��[����g�{�C�z��u�,̛W���7j�8e����y�M#���t�JI��%������c��l��fޅ��\��|%�*�r{5� ��<���>Ih��������w���6ќ:P/��a���b�w���v�_Y����7;.�YG�-���x���)9��a6���Đ1����6Y�&�h�b�@�3�����a��9:�thS�G���DM��Ϝ	s�+^�6x��բ��t�.�`ꗘ�"�,�]�و�y�����
>��g��"�J=�ݽv����}7d�c�����<���(��.m:5�{w���b���e9��us]$�˪��{��_V��Si�qܙb�娻�XUfX��b�dT�{����S��X�Ή��SkN��;�G�iZ��u�}W�%]Pïl� ��C2��q�S�Lq��s��)�F�J�qԔ��qn�g*_$���hc6��$#r�JY�q�j]�J��Q��H��Q�n���E&k����;��.�y0�s�X�|w�ƕ�S��瘘�>Wh�fE�}� G��v=��䕍L��*ʗ_:{��4��]s܈�'��������y$<�z���5G�G���4�)�V�pY�/��%�7�����I]'������G޼���T��}�ݮ�Y���{��!�?>��8x�o�!�Ou
��9Q�2��uG���plW2���|lpշ�o[a"��6���+��K�(�{w���rI��|�7eInD�x�F��P*�`��+>W��=8��7����-V�<\UcID�g�y�J�]�q�	���i� �e�C t�qn��ǌF;E,��/��qWub��5Y�r���ɩ��5|��\%��U��;�KS��6�����8���<l>�;_�_x>`�So��u괣�?^�ݯ��sP�3��Ĝ�J�v2ݴ��:-���퉾��Y=���b���1��PWC>;ՠm�n)���C���O����.��Evg6'mz�B�4gns+4<1�z郵v�+l�8���Ƈ�v��' ���@�_Զ��ľ��&E���w��G��yw�K<���Գ�S:{T�Stu踍�`���u�T�K�����������K׹l���o��f������fWs���+z��]@n@y1m�7�_7���fg'�V�5���]Ԝ˭�At/Dr�n��Hb��7s�eq��Ht�s�,����k\u}taԲ���P�z�ݏM`s�}�K�V�� ���z�M���+M�r�l�sɾǋ���u�&K�s+�'S����wxTɡoW]>�ț�;	S�m΃��wFL�E���J��__�+����!,n.�ZDg�L��#�O��؊a� S7ۯ���W��|��rE�wà�<W��Y�7ɓ��EI:ԉ6eb/B�-ӑV�Ks�͚�c�4p��Q_����T�g�Z�\,��R��H�S�Ë�d�8�'u�ͺ�$`�����6�>N��֝��'���>�p�W�dI�Y���MU֓Ւ�7Q����X�5s��u<��cT1Xa��3M�є��B�(maKz��3�qe]љ��W�Gf��G���5�����L7UO���b�'p�fR.Z�N�+$2VN���z�	;���U���LW��mG9*�K��ؽh>׾�9�o��䉘���c�
y��κ�h�ЃlJ�4��I���{*�#4o������)rF�9�4���t��]Me�	�t�^���-�ȃg����[X�}o���Z��N84�,�+f�:���iַ�,��ޞf��&V���8h��˃�l�x�KG�2��OW��[仇j�}�$#~�z��p���][��!ÓQ��Qt$��c��
�xB�Wgu7�0]Ć��9o�����Wx̋�iv�����.UAU�!yݖ\�3]����V�xz�l�ݗhǖ�	�i�';��ⷴ���hf�;G^����H)��Y��q;eN��XJ�D���*X 9>�a�g�{��H����[$���G0±T|f�K��]���M��n�����&��ln[�:���0ބ/Lu$ߢ�a^FC2։��Iۋ�VJ�������S�.�q)���^�f��Ү�u}�b�]�KR7�o^A�fYB B^��}1�}���ak<�w�<C�r��WxՓ�h�CY+#�8o��=�|.h�(��S��g�>��Y�v���T�PPɘ��ST�ޮ�X\�;�t�����s��y���^ó�ӫ���R��4���Uvb�G�8��-�O�`�F��Sv�	y|����zL�����A��}��1B>���k��^U�Q$v�e;�4�� �B<�b�.���N�^��SQ�on�
�-�%f� v���]��.�Onywv�$���O��@$�IER߫��������?�G�4'�>0��?8�s�d����F�:�D� �����no�l��r�{I��s�Uksh�م����ቿ�������W8�5�.y�u��Oϧ�{�1���~5v��$�l����ɽ�q{I�!�~����=κ�=ZR����<��w����$c��sع{<�P�s���"~�Csޑ�7����:���i�=��M�Z�/���;� � �*վ�n�!O�ap���m�U�������ѳ/���v>�8-i/@إ��57wf��2+g���ުWiY��),$rБ��� �ݬپ��~�==�����{�������0*xxzQv�]�P��_/n�~�}��^,�4�5���'\�-�E����8��N�m]%���7t�&()�V�xHu�r��K����%��l��L:�#f�����}�غ���=����q��N�����3D>���'���^�wG�����(�h�'~ζmb$�	:1:\m�с�N�obYk�hp��t�fCV���	L5�BA�+FZ�J���hgT$[̄�n}H^��ë�ǡ�s7�;�	tO<���)�N�n�!�C��j���gpv��GJ���ń��7��Lʛ�*�op��njR<U�#���J���]�wn��I.�8ˮ���{0rz$��	��t܏8���ټ�t|�X����j�nH�YM�H"���(�w �WͳJT.UQ6���v�&gߞyO�H%�f�)�m���?[s�i'�F�v��cF
ѡ������o��[h����j�Z��?8�8�M�ݘ���gc����֙����~?*��v"zqۻ3j�ճ���h��GDIGII��Pv��h3ϟ�����'��d���ئ`�E�N��tb�5K�4���wqv��AO<����~?>����j����F�R�uX��hյP�5v1qݵ�΃���n
i�]iZ��Mv�Z-Zر����b�ۺ����c���(8�أ��ۣF�.㮺4i�յ��AV���.�4�uwlQm����kN;V�Uv�Mv��c�ݻ��1]�h�jq�RD��\tq3kAE������1����E�b�e�ln�wi�m��틭$n{�(��ӎ��0�[`��Ѯ���3�u��Ѻ4GX�ڵ��룧�m֨��:
v,�$�	�m�K�~�!�Jy���ǯAI��N}2�k��y��KUƚ�2��״�l� [|Ŕ�P9jkâ�+��M����������N�]�c,�}�t�d�qg/�VL;NN�Ҥ�9�d����Ӿ߹���Id���)G&3�r����~+q��'�z{��9才-�!�b�}^�n%��� ��.cH��tr=�Gmk�I�<kV��M�c����t\��~����EW�����=�B�͂M��	7V�i�^��v��;����@��6m���f �m{ڸm����oo������@�s�S/<=Qd}ؤ�1�kɭ�/�1����{`~�vi����<�4���w����%�h�y�v�\\_�����DWa�F�=���l"x��֋Ӿmh�2�{3�ښ�Iڜ��nm'vM�t�m��N�I��6�\�wv��<q����+�g������}��c{{N���$���1�sY���	7��Uk�{QV�~��qcø��[r�a�w�^_{CW��gz�=`��Z��tB����,��1!d�B6f�o����o=帿~��-��[@)���H~GbB�\�|�F%v���{ǉH���#�`c
�؎��oj>v��Nz���ڽ�|R�- ���W�sp�Wa��*bttvm�=���5�6���jߪUөb�zX]9my�+X_�ӵ���f���3՜a�</�\��NA���e���^�.^�w��DW�>�ru�{�0g{��p{�_��L��O�A��KӖ��/?�<���>���%�~ð/,����#��'�� ���l��س�N�ݡ9���!3�������ˊ�����A�����/,��v�Y1�ҿ<��u&@���Oxڣ������:0��d@����&̙��v���g?������C ��R���=��)׻:���=�p���sW�����Cv��Q͝;&[6�(��.x����e��3��-��n��W����K;���޾x&���xξ��k�ϵ���5ƅ��ӄa/qŻk�6��:�/�ǳd�|��תtٻk�}@8��Wx=�Z~��˵xn�;�/���N����,l��x:�r��{���� r3�%u�r[�C.��Fy���T�� T�//9y�$}�>J��E�j|�Uэ�)C���H<���ռx�N�_�M�[��Xڛ}�t̎�ENC���Q?��It�N��y�����\�<�Lg�7��+���y�NO=GX���^]E���-Z����2zz���<6y������L7S��;�y�q+�YVΏ0�`w�lΚ�L��u���t�8�YK�W�Y�8�������Rq��9�vZ�|��9t�S��>��o��S�آX$�]m
��~hҏQ���3Y�=�y��U��}+��z�/w5�{�9�ۇ�����ކ�7\���=��͆�1b�S��V� ��g���:��3g��<~N�N��:�%Lq�EFO���͸�ʽ�'2�������>��NeP�?|�M�1}zk$u����H#֙��"ʢ��%L���ԥ��*�X����rO��;�1k��8��ʯJM��G����Z�[eZ>y�rg�������.~�g���4�s;��Wm�؉���FZz>���HM���Xd�7q����wuÓ�h]�,�3��ځ_>��b'3�7
�J�e��y�+�{,_X�K��Z����՘�>����_PT�����\����-	��G5��k�J��<bP�馝O�dڞ}{]�
�}Uڇ��_ʙ�Y;k1��z�꥛���͗3|����i�x2hA�߼�����=b���N2��j��y�^��V2���f���[��k�=�Krt&�A㞷z�m��6���SC��y�n��*�C�1��2��f�&��x�G`'{�1��v���3�8�1w3����]���\�N�%<M
��#��.O+�o��q�o��.���k��_#��>�yg�S{U���l1{i���a��)K�İOo��G+z�o���=��8�k����9ޘ���~-��"�v�q����&�~�O���~�Ni�,��������8~�sɇ�K�f�^Lu�i;Ä=��gp�����.\s3S��y�W���j���u;3��ۍ\7��GG�i9�>����f������v�_c�]6D>��n�Y4Nn&لB�f�I:ݹ�N�����Zֽ��b�[Oi��f�(v䧓a�.�q�b^mP���q�5#m��(-hac���#M�6at{�"��S��9jݴ�Z��:�W-b��<��j�v��T�%�\�s��u�뎉��Q4b闝�
L�t���4��6�,�׽❼��G�RS�~ld��/n��)xߛ����(���נ�Wl`�q�=t���c4�W\g��A��ʧ��ٵ�J�q��}cb��X��+��Ɉ��ot�=��[IӼsE�ˢl���j�=²�������&����N���p�ݚ��������OG{I��扴���4-惌ʍ��Ѧ'�CAAf�;�z���i�^E���w��<�5^Z�D؈@�	�'���z��I ��$m�m���rW���$Ե�aM{�׻����;���^������=��D}��Y���=`�:�gfE��Κ�9d�d������2<g��m� �Nw,@�lN�Ѷ�op�.�Kqֽ�ň|�b;$��o�N���}���f�K��.�;��-}}����*�an7����UK}S~��撔�㪅�w�Q���y�����OVa�.j��@�M��t���$h�]1n�/������3���85�1g�+�S�F�q�7�����x�ms��{(s��a�y�w[��ʶkYS����w#%[���1�3�A]^��`��{yo�;0F��uۑ�V*Qҫޝ��O��.�Ϟ�mr���<R{�/{�UM�Ayz�� ���~.��+�S�ÆI9���L᭞�F
��3¤������9�����3#��ޢm�}cZ�އ`\���<��y��CF�;���r�dzT�;�x�3^߇P<�4qC���Ր{e������s{����6R��}���Q��\a���|�k��c��e�5`�Ǿ�&d��+�R_���\�b�Vԕ+>q�}�CC�f�T��*���9U2<+�&�N��ط쇧�i�\�Vm>�j{��mzAyE1��j�Z&6�4��Էv�ݦ*v��C����>�\T�$e����{h�OT�{�0��$��������-���cz^⁋'c#7��I��q�p�f]Ũ��o�힊�*w��x柦j�zv��#|�m�^k����\qFF$̤�nYS!�%��0��hfMw�_��&<�Z^�����x�)�{�v�l\�y����>ǂ�Ԯ�ڸ��E����:�y,��)���]�SRcʌ���N�n���_~�L~_c�?g�fa�%*�Ҕ���{���s!��{*7��u�ӗk��B��w����T��J������t����-V����:���<^��)�ƨ>���=ۙ�ةEB�OnZ� یf�Jz)�b�D*Lv�����y��#^x����m�ھ�Z�:���^��N������~�+�k%,]=�Qxe��?O	6��|zxxр�ʾ�;�μ&�`���Q�P��-Z��k����d>^
m'cW]�Z��2y�2�=��t���R�l���8;��uWt97Dq���؆���{�۬�9'������;]���b�Sʔ�|)/�&�yA��Y^��$G1u=o��̏�y��������e=�o�񪉁V%��L�f����ڟ�y\���'��=��C~��[�s�Fk��e�~�b�e�����9Wra��s9ci[^�S>�t�ގk4T��O��ƌ�a��-��z���E�{wcx�u�Z`zډ5P��!|	�傭�����c���^3���֬8���~q��^�sʞv����j!�0�[�,��w�V��������b��*sel�2�w�Q�$y�O�uӓ.n�;�w�X���0�2{ƫ#:����R:���fn2�8�3�/5_�3�*���O}�{��T�`5�h�j��`fEώ+j�_=WR�j\%�	����Y���.���hy�3��$K�_����XD����{�g�h<�t�ϥOd��ױ���&���x���X�K�{R����>�R]���hmёq��A��$�8dǪOT��ؗ7V�XO���~:=ۘu�V��,p`e�6�s��j���M<g_.bs�sŤ��8�S�6��;ӆz�
��vJ�^[n���{Π��cfs��<�\���3����`�eׇk��>��{_A���g�z��^籐vrY:WF��ɂ�Gm�{7�v��W�	M�f~���x~k�� �����{�4���|�N��Wz���(z��:�6^�̮˂��� G��m{^�}���@:�\���rcN��W�6K�0�-[�$�M�q�,�٫�V98a���s���9��� �������S��L}�t�{Rql3���C<,澸z5���KI_����������2�;\��=5�o��gv����X��wR.�Գg�ݾ��0<��Ug��=7�ssN�eW��{tW�R����K����bȗS<+Ry����y3W�������]Lռ绲?��Ww��!��}yQ�'�����ǽ=�A�˭�w �z�b��g�r�{�_�stM��v$q�ϡ�'j�hf��_`s%A; ��|L�P����~��w�~�i�
�j>c/�Lxsz3�~�ʾ�߼M�烵�{	=r�9+R��{^�;ا��: \�d���e��x�'��LuE�r�U���w�� ��dlS�,��VK�4v ]ǚ�+���q�pܟ�����;�E��z�^�Owl3�ަH����'f�j����]�鋝�#��z�d;�9d�ɍ��~(i&M�5�;��Rf`��K�Л}:�x�K��I'+׌�m_�R�,98,���]D6јl	B?�f�2�U��+a�aUн�%����.�t�τ�Gv��s6�-B�fwq��(�
՗�j&��)3m!�,��I��43n�����or�>���ئ��1����Ò�O�L�FQr-���6����x')�2�t���[�R7 jg|}��7g2�ʲ�����������
X�����x�C��6}Hc���{=��l��W��?�-��폇J��w�6��U�ц�2�Z1������CL�65�歟�g@F~�xx[r��'r	�nweuv�T�$�N{E�g�������z<�C��9��x�bt�b�u����ۨ��'��ɵ�"砞���{�u��*{}���d�ͽ��FW �a��y�pó[ӓkg�у���_��N�	�W�}��8�ɶ���4^Trݞ:5��8��[�h�o�c����ͩV�����X��>ND�p/Tf��\�W�j�,#-�=[�Nt�ϯV����D#m�����:���7'�#�WO��t{a�ς�|=>��ʳ�I_Z�g�ڷ`�r�m���*6&rD�0Nu�,K%�tu�s0�贊oc�f���et����|� ��ufw,Y��*j�o���{���\��W����*]j vX��^sn��}eV����� �B4C���I�:��lh�>y^��ͷ@pv�	zo�y�����8\�[5��vz��|�3Z^��v���q�]wE3:��[	�لc�|�&���h�N6����	z�f�⠔�7ҳ�I�d@nl��Kܞ�8���>���y��Mg���[�4�3'.���3�-�|��6�D�Z�9gBT����)���9l�r���z�c;�{B�r�5%Z��ϖ����%�c
��+S���v����\��f�G��H� ��`�ב��]�[;����f�ۺ}2u�m�E=���ǲOy��4� �[;�}�_x��դ;���%6�����b[慭;vf.�n��ٱ���^^��m�1�j�|�4����@�y�_�'�o[�9�%�ҁU��գ�s�UZz��%�9i}[i+a��-�����h+3��{�۞U׵h�^]S���k�=�c����(�q{�=F����	*����ܣq�H�u���C�,�j��y�3�c���߽�>fwg���v�TJ	Y��x���-�ԑMl������qs^��/7�YZUq��2�ͮ��h��F�����2)�}���E��@h]γ�+���1�XޚNէ6u�l"�m՚Au:��Ƞ�yY��X�����|���m���w[�}�n�v%�M����V�s��Ý���_��[+��{u>M���EM�+�8'ϙ\5fU�9U�P:[�!��N̘Q��z-ŭ����O��{��-��(EB�>�k�{�^��g`Z���pe�8]MI���WM{��W����ػG��,\��&��@Sp;�;}t5��%�6$�\�ʱG��m�yӀQ��=s��<:�֎��0��t��u���Y�F]�u��iz�QqҔ��5��b̡r3|w�lm����J�yk�Ԣ�����n���]�������aIq�������9ӎI�<zl�W{�q�M2|�L���pof��Cڞ���/�W#'ޜ=���$�?��
����e�]��j�M��2�ƅ�]��q����M��twp	Զ<}Y���$����a*0ob��9�/53Q۾��C)ptY�-�̏�+j��yu/J�E�|޻���z�ACܸ"/ֶt�T{`�X����a�w��=�������{n�!D��&���dvIʎ
��[�S�Sgb�ql�V�7Zm�`�i°S:�*�^۞��˜���`܌��u\�A1�;s�/[����d�����j�)�����H��p82�,oM8�;�L�H�>�0hW�T�p����R��'�k���?���f��V�7�v���SE��`��9�b��QF��W�g�TT�^�n��>o�����v(4_6"����zwfgF�4TWc[V�w'M��uݢ�����[z��Rs����?���QO�uu��|ظ�n�ڌ[۽�MG��lb���cщ+ӵ�v�W�A�>~?����ƍ�? ��ch/��Ѫ�{�[[q�����\��5MPEOE�;�j��cK>y��~?����_,Q�:���Gc�me�#��^�ݪ�Z4t�Z��V���*��g���h0\\���\�ΜpX�i�b=�Nuwkb{�q�׽ޏ^�cN�G{�ު*�<]��]�wv������\��O��|���[����F��6��:�N�h�jܸ7kk���8��\�ݜDn܆l�k�+�wb����Lw<���[���u�pc�[\�Ѯ��������pΞ?=���oΏX��ִ�G�1���b��{DTG�AA�~\z"*,U�A��w��tx���b�Z�1�lf�ێ]�j�ͻ�n���j���{Pj��vWd�"+}G�E��9�����oQ9ՙ[� ��s�|��-��rJ�qY���X����&:��3[Fe���� ����z2x��&m��eF'G8�s>ͬa���H�D��v-��ױW�%����==�ed67�2B�a�z��M�װ�αm f�i���e)0��^ͧ�͌�
\��
H�^�V<g�[�<� 4�a0�|l�M몏O=nL�P��m���*'~�W�]&��j׾c�ze��%C�zǫx��0�{��y���l����U�
�دH�BSgU�%%�����ǎ�;`��U��^sj��|��u������0f���,-�s�[�[Xrz���1v�kgw��l�B�Ĳ/~)M2�e5tF��W��<��w�J�.͂}�l�#q��L�]�*搄�I��X34���1�.�,[�����[_�vO5y�.s�ޝn�/hG<�]Z���rf�y�f�p86�vK�S�&HޣI ��I���"����u��/�������$������#�{�#XX!���smLpm�� sQ{:�E�M��8ŧ���inF��E�alC�a��ǓS	��P�CN�U��L8@m���Yc/y�����|=���	�e�[�����f�w2��]y��j�P	g\9:�U�K�9}9~��1'��{��TO][���҇N2[�H^�jQ6�>�WR�7��O<������خ�&pH���s��v׬�AiQbX����9�S����Ղ�/gd�]!�.g9�FU|�]�z}����j�8��O�� Ļ�{��@C`t�~����C��s��S]����UD�B%f���V����<��z9�M5^���T��b'�2pZ�o)��ȴ+�NJ[����tt��#�wŝ�-Xs)�:��X�8�����1\�_o?����G�h��l�o&5>߭*�:/��[z���T3y6�q�Xi'���0�-���j�[�X�È�L�%�?eUd��
g�z��������#X�oP~yÆ����^�'�y�@��x~��vp�g*�tj� g5�&�_ ����Qu�&7^߄��m���<��ti�k:x�aE����{�*/�խ���y��~vj♖mYa�7�����	��a�-�{Y�_g�b�Ʈ�۵m��t�r։���+�AFr��˶��Azw����?�P5���PS��Rʓ�տ	Qp��Y	QV�W!>����y�X�5����z�9q�̂q{�%�h�SWe�t�����㝯�s�#jQz��,}��XZ�R�%����i�p�DJd)"3O��מ��/�î�Nȶ��Fǥ��:��??2����Oc����۔��'��y@�%����ETko</ ^����g3�6�If��R�@�'�X��V'$~�0�b��W�����Z�J.2�h֔��o[ *��&���}����3���>^=<}�b'�`�Ľ �	��s/�^:�v�@=���R�u9��v�j;$�5tBd�����"��FU��Q�[�fr�jٮ��MT_}��8,6��!?�Ҵ���mΈl��*L������p���垾��kL>� m׳�����e��F;�	܁fƘr�8#�; K*���`�fg���4���ۂe�!yCvm�/�P���6���PK�+�+?>�m�n熄�$U�Y�nD�^w;<v�	��T�UZ���;p���%�;0�Bxwf�}��!��ej4P���)�g7;.��-�n):�7B͇2q��qVXZ�%�X�Z�5���[9��Ƹ`�p=u��y3'f��a}�U�kq��
��=1i<:�=P9��MxZ���е��%�J�`�Dk0�(G<�R�1׹Y�۫���`1A�����\�|~p_%-��u��)P6˦��;�X����ߓf=��8�<�\����3L�@�z���'��&4?�i��� }���z�K���d����N��1�������~�B}���9���P�,����Q&;�	bhY�O�Ona��������7_5��P|�>R���!)�s|1)���Vl���p3������n�D!�\���˽���9�v�.��$a �	�s���t�B���B�WY�ͦ�_]�=�#�&Y��*��}9O��{5�~��#�����WC�-��� �H��O���U�5���	A쿅8�E���u�7��5��<�.�TZ{k:�N�f� ����#��Y!L���i�������Nr�d3К�6��F���A��b�i=�F5ld�Sz����B��A�,�l�<����d�l1X8��;���>ʸr�������3��GCY�d��j[����`q��,R%���^�Ʒa�$)ռ{w�v�|�n���4l�~;3��H|�&B{(x��v)�{�	L`v��X���yʴ�[f�:���,T"�]��1P��g�X�}�/`��;M�l�#�ū�zC4���l1y,�\�ĲoX�ƒ4�S�_8���OZ�� �6O������J�}3���w��W4�U{E�}}�0�U(��rt@�oÒR u>��D$��6l'x{KZl�[���+Gb�(F�И	��ؠI����U�]����n*��0�ԜK�uyI��D�v^YREN��r�G� nf[Z�!Ƅ�㮘,h���y�\�זGs��T;��6ĮίO}���?.��J�fB3�k�7z�+Jо�7B�{<�͊�[�D�>�|f�}�ͧ��yj��=�#[�%��������J����SM�<M�m���:q��>��"Kr���s�M��8���&R�s:.�Y)��v2G1�����7���b!��z�}`u�@�3�P�{SM�����P�qk-v�U��t���}��Xs�6r8�.�[���w��� �a|y ����[�^�c!��s#)���U%���5v�i���&}8�8́�^g�t�l�v2X%p�	���򁩨��gm���f;�V�z[�C����I/����H��@����Űu�v<��H9a7����P�7\��{6#H��?8Q5%=�j3\�k�̌��ӽ��#�����6|�����%��fw���+�������=M�-�yM- X0�a�=OE���oP���f��{��VPB�FL8|�]Y���_qH֝ϻsӗ?����-3?b��X��KH �i���7����ܙ���S6��M27�ы׳x7%��ڳ��f�O�G�����Ze'�1с6�?/c�o�?��災�x��BV���ufN��>��ڏI���M'�t�ʭQ����X���0���B.~�x'����o�.�R�jk�ޓ�6d���,]�N9<2�C�)�M�������`�cF��mxRt׀�gN�>�9|l��wN���G���x*�M�H
|�ѶH�],Ks��V���;v����3N1���L��M�3��5��1}��~�c���+WN��۫z��]��幓4�'�Ҋ�S8苆/�7���sa�m҂��T&��;[�T�U�{{:��C�߅�\���t��l�a8�;o���%�oO�1���\�8C��>)Յ�)�$i5���j|��N���������뷽;��HT;�P��f����}�.�vA��eF"����q'���α�^�/�Т��Z满Ң]:�>y�!���D&���gۓ�EΨ��ft?���9�LZ�2��-+h��}���|�S�z^G7�<��z���`d0Q�>�as���\�&%��uW0pc{�Dr��|�׿�_��+�}7?o�A����/�����Ѕܠh��WU
�H�M0�$o������pyD�#�[]��J~kL�z�S�Q�ޱ�n��;��n.�F!Xb�g���i]�ɥ�]C'U�ڨZ�R�è1�e�~�J_�����#�9�~���'�rc/����v�n�cpй��BBm�;&���d�YƄu4��~df�W���\b��-�{[)��'ZY�M_µPw�^�s;BH0q��H�J��x?<��Bk��v�e����|8���Qx�wL��ލ��x���i��4���	���i�L$��m��{�yf��㉆���Ѽ){�2�����e�����o��;���3��w�,]|�ޖ���W-��_i�.�b�<v�H��AJC5[��Y!���y+�v���k������!��L��!�ޫ�2��RɎn�TL楇��d�$�E:��@��z�"�cO�o��<� |D=�5�ytA�)��6��1C��`,鯖~���%��:�<!�v~���eַHN"*�"E�3������!� rbԖI@g�ٳl�n���	��
�`d���`�$�-<B{�e��5備�ci�:	���j��Ռ�u�5�m�1Q���4@�ST��9�>� ��G8�Jt�񡑮~wA�>�N����-�L�������{�Ce�|����j}���N?���fʘI�r�ᝒ���D&I��Jue*�*xN�R�r����j��4��8�}��_�ύ�A��qp�2�6�ۃntC`ޥI�ݞjW�v��xe���q�mj�υ�Ɓ�����O6�`A�v!���L9�<%��,҃�gtQ͕�si�PݓW�Ͳ.�Á��j-#��]���?0/!��@!י��C��υ*t�4uVDմ�;ռe�3�3�����u��]I�P�9�D���Z�� �v���������cv;J;��v)�`�9�.�[uԘ���>w�d닾*�
���W1��\�5���@�zL}b���H|,u��ĕ��I�j:���m�bTǍҏ�jQ��K��Y�zW}�H[ob��l_�@T�Q"�aK�6�n�`��֤�G!4��R=+~?|����2ޘ0*���25���1>����D<�n���@{��Ͳa
�A�}���R���@Q̨uH���4-'��;����{*	{k���@�E��!�1����ž:䛀� ��\baw_�0̲�Kc�<��D۹[��O?]^U���:��N T�����rL�w���x�	�!�6߬eK2N��z]�lcS�YT��b�r����o*`���D�7c�zF`���W1eyO�T]���á��whO�(d�L�m�d�����-��݇aV�\	΁�� ���L1���:&����������[F�ʧl���}�#�<�z:���T^=�k�h��C�W� �p+�d�
My��i�WL\:ɧ�ճ��-�p�E�C7'gHBas���[Q{Q�]s�-mG���~;2��B�����y��&����[�����>��P���g�#�9g`��6�K2Gӵ-�C��[���{��[ŋ�qN���V���:|.��{���6=�uP�V�������Ip2�7̐���أ� B�Uo{KX�����nz5!�άIN)0�Q�oT\�����>L�!
\׻��n���5c)1�+�e�<;���1�o����S���`�[��8#JIˮ�W��d�&��R�F33g��|���$;#��+e���1b�����1��.֎ޣ��AΚ��&�{��9νe<V$Yu;1N���T��m��ѹB_�o��;=y;ŭ��	�i�RS�����ƒ4�4{���>G��ʂ��Ǚ9�����Uґ_�3�n�p�"�	tH�ơJ�u'y�E��R���Lh-������A�7;EgFӳ����������f�B��*`&���;JUYU�"(Y�O�b�RX�����z׎k{Vϝ)���
K���W��\t����O���<Aj�v�߸�0���Ɣ�ã5C���y�8��7h��U���SӇ�����tz:���mE6��U�V�V��3����8�r'h�A��D�s�=K�J9�P}w	hs�M���a1���~i��HɆmǩ��ݼ��Y]<�D�9���uJ �,�I�Oԃ3\�Q�N�a��=P�tņv%�����|�-g����cq�y�YP��f�vپ�\�� v���wX�c#�]�F0&�+dc5mO'���B��!�g�Ѭ��{�GzC�ͬa;�K����Kz���|p���73f��}%��|��`߭�i��/Y��S��f�3������Io����4�Un�i�s����d����r��}��vz�˶Ut/:����<����hI;�;�z�5�:��Hh<�0V2���u�ZhG4��gY[Yo���P�.[�coCy\�{�v���hB�o��@��D���v/[�W�}���w{֗oz4�>����3cT)���^6#ɡ�22��ǣ�7&m�rTͰ��C5\`<[���D5 zq�n''��ٳZ�_)��d�7 t1J(=�f2���!(�P��M/Oq�{���>Ab͜aL}iM'�]8¼z/����q��O��d"�y��ρ�	Yk_}�7��Py��B<��gA8C�K"�R�?[�!����$��M�VWʍ��o��N<ʨF�O�&�2���f�,cEy���&޺"S��N]�:>]"��e57Gd�(O<�r���{{�z���<����
��B26��S�.�Od�q;�i'���H�F�;U"�^�J�����l��i��,,&�z|�>����3y�t�bc�l�ry����
��* K�e���`���ĲoP��1ov��%����f�H=t!��|����_��U��Q��l�@�5N�Q�����Fe���v��A��w�r$-����J#����!w<ò~7Q��2�w��l�+��H�|BrE2����6g��'浦M�X�#�L�f�H��d��qhA���_
��|���{�����6Ou
o�z3���#�J��Cٲ��j��⤩��P��;=&&���tA+q�Q\t��c5f*�{��gM�����2��ڰ���L�/5}����OLxo�9S���3G�͢�����LߵA�B��{�Ǉs��E=�w�EU#B��f�f\�zGHiC��;:�cUh1�����=d�-Ѽq�����7��K�q�L��x����t��*;ͫ
��X%`8o�ǢWK5�t�L�ؠ��;��8���X�c���muN|fĸ���ݨo�a�[4F����U��m�'����w�Wz�h�� �%���U�����w�.p՞Cc���z�y	H^��mZ��'hIl��2�d(3�1�1I0�Trx����(,�����:d4o:ok����"���C�,����L���oW�1y#/�2��S�^:3aN��3� ���|��6�}ad�A�>ϖ���F�؊��J��;ztb�C�ă)�N�0����9t���Ts�a9u��9d��7V;��+u�(j��r�3�ա�����&�M:ǻS�jӱ�d_s;�m�٠�#�S�	�gC0.�]�Q����)Ҋz��)�n���;��{�������x�rб�Yܬ��h�b�U���j[.��u.��@�WwvJ�pj�X]���T�q��IB]��dZ.il�F����hy�/�,1KJ������w�L���]�5U�U��C�}X	�*�b���7��OϿrs/��oI�M��7�_��ǘ��}O�K(�6��0a�!v���`s�;銫��=�Hk�̝oKxfǚEh?��s�{�lP% <si9l׽z�GP$ӜK�t����{8֌�	�S�@��R94z?xZT,�������]���7��I��]�r�\�L�=ʓ^P�>���-w1v��2��5���Tr�X�j�(�(�{	�����*`3��${���AB֛��T��.
��x;���'}X�[WM��V�M��H�ꅕ�o�����q�r���:�݋�W��k������+��v�}�nt�{��2ց�n�y����f�0���[}V�多V(�֎����7���0�L;��5������N�/r�6u��@�i^w�Uss�}Vgw@�s�1n嫜s�v��0�:`dX���X��Ȉ5�V���״����r=!q�e���e�w}˽��'-�'#��ΜO���tY�z@�K�sVG�`%kB��\r��4�9�r���Wux����N_S`�lq���ݾO�)��A}��_8�R�ĻVs"n�Ӥs6�
��v
��=�-�䰁�/C��A�+{��8�`k9/�<���ͫ ���;�)7����@T��5)q�C�ʙww[X=2U#FB�?�<���aK��%�9	��!�˵v�6YK߳H/��v���+�c�F�փ���TӯA�:M6�`�(��`��s����{pc�m���s�����>]�tm�V�j��[4�5E�w�1:b5�M��ѻ��4��%��t���;���?������%��Ul:��]m��E8��u���h��Q������hձ���Tkn�'�?�����;�`��=۬ml�1Q�TSF�b-���PQ��׈�iӷ���"��6�D�����~4|�j$��l[;mD[;mh׮$:k��m�Ն�h"jb�Ѣ�`��
u�*��i��F��-<TSULE[�ZH��T���;`��bt����)����	���M�~���1���ƻd����V�I���Ls�[E���؟^��*��f�Q�3��uM7��W�h���IQ�wuv���b�Y��&��t��TS��Xţc�� �� �/�"-T�^=�����u��Ũ�凟8(֒�m�X{A��^�{�^�����9V.�P���ú�w'��V�kk�T��)�yr�h�n��0r&Ch&_�v��}�b��v��aD�A�k-{���a[~�\���Hwn�9}a����ץ��0dzg�(Ani�&�zP������I87���0��:�q��ݢ3]	�J*��ξ���|d�ø�vy,퀹k����7�#Y+ޠ��	�3E�q51[K w+�5��ۉ�Y��	0��R�����$�����o������m�;�凐MF�;����ݽɚQ3�ڒ�d�&a�[�Z~h���dS��(#��["�7˨B�c0�Sԥ�=�^I檎���V4��Ppq�nn+$���͖~�(��r���1���ϳ�K���f�/Wq��;W���DT���Jl]'ֳ��z��Ɗ��z1���PQp䎸f�1N+"l��y����s�3/�2M���LN�'rmj�"��F��u�):��|�R�*�
f��s���I��[2���u��%"��~�v�Z²�����]0���;p���� &I���3I�͹��<B�k�I�������@�F�!k]����~��A��!��B�^�.�<�:3��݄���{�kC���M��n�h-Q�g#�nI�)���Ϯ�߆Jr��������c�vp{n^���Cn�!O��� ��:�gf�(9R.�ס2��nm��)���/9/#��{3_�oo�Ӈ��M��x`�2b��lnLu�����炖��d�t;#W5�8�'Z����L��"j��>��dc×������Umf���"�jF�q��)�Sat�x��\�6�;5�^w�~y��B��/�q͓�b�"{n��T1Լ�a�H���&f<1��^�JK�;P�Ja���T%���Dj����2�b���Ƚ	�u`�в�8�*y���n�3���<���5"�NU}��ow���
�ߟ�B0@0���͵��B��(��:���eA����|6h:�j��ټ�.�������,4%5���t8G��!��0��Գ-��,9�
T����)���dS:�ݮP�u��yU:F�(���z���Ɂ��D&�#m���,�:�:��2�ܱ��)�����b�Ó�s��'�WzF`��g�9�+�~�1'Dav�JsBʖ���|+1��G-��EܦGz]��zO$i�Hz*:��Rѡ�tM�;P��J�]KW������ƊC���2�2�|Q��ٯ}��f �ݎG9W ��My��i�h�F����
���)B�$s-������ZÉ�g��!�*�oV���A,j��YF��-�S|6�f�Xe�.X|=�u���EDY2_�w��{�j1[��r鸯
t������V�e��'PU�lj���',Ք�������<����i���B)��K�9�����a{�۞YT��X�Pٯ�w�-{;2��B��׈�b%��-�u��}ܞ{�]8u�q���*k��Bli��0Y�?;b�d�v����Bk���e�8���������V1���bC�Y����Br�1�6�~ ��>��r(��p��)Kϧ��o����-8\���i0MP��o�v����z��C�h.�|���ι|a޶Ñ��K�0� S�\����L��x�I�7E1�/�__�;�(+��U�Jcj��t��]���h��j"�n�	�A�8�%P��� _EL,r�E�s�1�b�v���m�-�S��`ȅY��t>Π��p��((f֘B ��7vt�(qUeWC�zO���,N�ag�w�SL��;�L?2�K4�a�~!���B�� �==Q�/�g��-cp��*�;��Z��*��UC�IǺ^����q͠�8x�d�Bu�Pp��m�M�!4�D�n��`����گDqf�Ŭ�a;��Pq����^���kv��<����{<p�a��!�]2�& sJf-u4����w�rEڱ&��z�f>}�;rh�#���p���b�s�~�=�;�$��uL�<��¾�2κ_��)}�U�Z��
����>�s��N�dR�h��.�,O�������S��=�Xz���6矯k��՚�C���n2'k{>���f`��pԩ�7&h��v�WRcl�����E�'͏\fy��f4b�;3�0�5�cT����E��4���T2~��!�g�ҋ��1�/@�~J/��M@؇eu������Y7�[�u[��
Ò�DJ�Obu�5��4�ͬa;�Hz$@"x�>y�a�6��K�h�j3Y���Y-��E?����ȖxBid�Ų�'�'�Ӛ�x��9���5��,:ZV�(��{���Z�f�!A�}{/�r����LX|a�|�8ǔ�b�~��nId���D��~o����6�d�X����R�^a�7�x�o
��)'�.���o��J�>���V5/l[de�Q�k�T�5J���"Se�R�&�Ji=�]8��ս4��}��%���M��ɺ&6ԛ:�0�w�o^vG
�TZ�!�(�E���\�I��m�s�:{
�\��cK{;��q[��Ȓ��Bc�)G\=(�^�b'�'��N�@�=�&����� �D2BgfՒ3�k�Բs��bC5��
�m���vK�]�a�oQ��E'*ܘ��kӟ��檲���3il.o��yX�������{���z��U�~�_��+����{�B;��أ�W�{Џ]�B%i< �JcR~0�X-C�X�8]<��:�5��}�J=��]�\�U�����[d���Y}5�2�nzOA��A�G�o�V��X)a$�RC���I?� ��k�]�C�pmt}��?�5���Q���u
Ѣ=�|3Ⱦ� (���k���
ceY��݌��R݈�C�nE�<�^��ˢXa���3������?B Q�W�@�Euq��9�U�X��-j[V�\�c�񉠲F�����^8���$_<(�>�Br�\O�Z�Z��W/�G&��B�'V$Ȧ.L�VoJO�koƎ=���L�g=;�n{a�lS�.!֜�����Y0!��C�:/]P��C�еaD��,}���ۓ\��_h?�ym�T��0
���;[;Z�`�т<!2i�����ϴ3���I��Fi�q֏m-A��wƶ��f�7��;:2�9���ţ�>���h�-"&9ف��ޠ��{=Bs�w2>��ߋ�=^�F��_�o(����W)i���c��/��|dL$����m������Wu�ϳZ{��L�%ki�kzO;QS��R&a��Z��E'��)'������y�&��6!���n�Y���nt}oP��՗����岐qx�7g��[4��yˆ@�t���N���c^T��Up�Ϗe����']Α�:w���*oY0{�s��� �Y�x�$"O�;û�n�ޔa�TǛF��'�o	�@����@�! ,B~�7�ó�ӗ$��. 6����]��\۾qb�/l�ރz`��z��(���ʽ���ō4�=F��_!�^�W�rFtc�6�B}k��A=P%�]6Ϧ:��K�^ڤ5X�E���e\9��9�!b%8���󴞝dՓ��!Z��QI��"PCW����5#/3eN^l��YQ^�u�}OD��Y��e��L$�;���{%75�L�������k=�n��l��m��iq�j���6q��ȶ{�� �4� �D9��ۃ8UtM�t���u������Dn�w���R�c��&*�<�/Iq�lGNc���q���<3�^.��'��tr�c�\c$�ڃ�u]YWa�k鄞w�f�X^6.hr'_����\=��ٜX�ϢWp�W#B�����R�׺�
6�aT,�熣�)=ZRXבچ�ٻ�TfQa��j��I:�˧�s�[o�7ٸ�u`�l9��.�E�ΎcF�k��KUl�D�ƒ�gVp|�Q�H/� A_�O�!ks8N��R9��i�V�V��cҹ��NY����:ձ�����)��v��W�XK�(p�_���|�Cj��O�ґ�`�x��2�{lf;�#/;)�����^����c�Ju�G�~�m	�S��:��l�6���ZI�9Y�`���O71����d5���J`�2m����Q!�j�Z3�w�>��?,��5={<sѹ��M��}�EԳ�k�Q��W������`��D�Y
�_J��5�c�a���ިx���-�W���1��'�$O�Hy��7���N�[���y����3E�.�vS�(��1%ډ�nǡ�fN��5�-���˺�)�ny����/��;Q=�r�~��ۇ�����]A�V����d���L�D[*oi
z-r�:ͨ�'LT���A�q��:^Ǫ���f���L"Z� �z ���&|ݝ�Zj�g���;sӆ�`�yL\9�S>S�a�p��%�UFW��2a��r���� �^ں�)���.=fK��_�w���(5]on��c>���O��~�w��6��)�6���j]��.�z6���YPX�R{�M��;�@z��KU�3��֜I|�0�7tնz���d��l�^����:j 1�jx�u~�0L��o���	�y�}A�68��k"�d,������ʘ'����ثӽ2��/�:�ǂF���`@�.-�&�"�v�cæ��7Z�o�5��^B����_�ݍ�.�/���ʥ\�,{غ��k�H(�/��yy�;��p�ۧjFӘn�fTt^`*�����j���w߷��?9��z��z%x����Ie[����c�*2G&�tuˎSӰ^�:�d��.Sw@����q����{��M��փ�����T.Nv���z��E@f���v�"�|�Y�5;����lg��&�"x��(qT*�{/I����NlKo'mv�Fkv�"/��4^G5g�i}�~/�����
����~_gT���Nб�94;3��15r��5ii���w��q�%��_��P�z��ť�����^n�?�ê~��4ڑ��"�[��w��l��A由n[*�������+������'hs�A�#	��������cG)�{���O|bg�Q�I�^��.T�$2���c�o�fy��f%�3��c��j�;�M��{Yy,��K�b�=���k��܆�k'�3��� vQ1^:��9��G�6��,X�\��w�-��A���LO�g}/z�4�ͬa#�%��^�֐�h_w�ɁN���r̩&x]7
/��uC"Y��Biidv�I��3��'KM{n��W�=q~�Чs®�aKP"��L8y��OC�m�k�<�-(_������s`UO�[4�E�\e��f�Bf��Q�m�vPe^Y8�̚ԝ��3f��ǫx]]�0��X_y_�>^_:�}�^[��$�K����z�<O�y6T X��+A����W�N@�e�E���"���"]�=�� [�n*��>߈$N4G���{�mN�~�:	]Y��xC6�;U˘��b����ٗo��oIMK��E�]��)C�~}����?^�����*����i�&Ba	�Jhe~~{��������{�Ȉ�Pg^zٝg��
دL��)6���SI�ʺq��ǫz�������z�0�v̩��JB%�O���A=����'��
SL�ҍ&�}���w�ـ��;�8��X
w^��2LO;6T�`�����GDJt�������7�����ͮӬ�3�bv;���C��<�������숏����/p!kx��Ε�Ǩ�͵�k���4v��5�/A�<�!��BG�";���{�ᨆ���]���:��4˻�;NZ�8��-?,O ���ˢXg�@~��-��
5����5-���Tk�F����f�X�l�R�(�,���w�|��|�!��$X��|5���dE��DT�-�Fm�V�K�!ڟ������,tA5mv7�W�s`
��z��S,�Cb�ٶS�kk�b�-l�QA��p��(9/0쟓�����i�i<&��k-{z}[~�\�����]�ʻ�q���� hC����,��ŧ���_e�>��4#�$��bX+[[+�Yr��_kݥI��ez���0�D�������͢ה�ꢳ<~FB���)�>R,���f���,�'j��͑yv�@�3�vy��ڑ]� ͼ�p�##���n��}+Mr�N9���^��Y}��U ˞����/��~{��Ͽ�ۿ�~�����d� L,���+BҕH��_?_�������������a���^\-|k��re?�X���O�ac�R5�ސ��&�#�I�����(���r?N>H�H�m���+ho�"��Ӎ�Ȗ� ԋ�=׶%��+z����OUWI��|@�^Z�i�]�N2H���o�i�m����	�ٍ�.�\�tJ��Z�t��O�~��z��J��na �B�@�Cb��ٶT2����2��v�|�*�n���.��wlǖ&nA1�/�|��"��B	�8�:WT�����V��<of�s�ެTj*k>�	^��rĞC(LN5;�kW�����-�3c������JƓ��ѕ�^w3�l�!����SW�nL=5췅?�?���M���;�;%77����&*S<:k����d;7S�lD󢔊P���|�`��Ы�� �4�t���9�g��g�a�TSS��5�_���o��Ɉo���|��L[��<
/^K��_C�[�K7� G��!8���1UC���η����z�C���تE�IO<b�K��i������1�O�8�܌�����Н�,啬�K���/V���[}�g���;��	]��E�Ps�h���כ��5�w"o�~ra/p�]�ch���˩�bB�VU8r���Yc�7��`����k^r��I�M^�w$'v1=�5ݼqKA�q�}�K{#t#�y�uWu]�������0c�����qY�r3�{>ϰ+Ͻ����3s�z�W�ɐ̉s��<v�x�{��{����2
F�z⻋�K�����NC�#T}<({:�}'�c����]}�r��*�)"׺"D]�rm�����=>:�z�\��=�Y�f�N�kqf��T����˾���Ŋ�Wð9����<�zNV$�g��h���:��]��.Īg�>A1(�6���p�5:�`gg-9[;���L����D�$�ڭ,w�͓�Bۑ�YW'[O9�C�YG��,�4p�O�ެ8B�Y�F�;,���єSǬ�drz8ݻT�M���&�t����O�����A����]�a�wI7��d�:f��:���/���9L2!�g�D���+�uw�07�"3{�lDF�#� 7����E�]&�Imt����gr�l'�R��SӹM�K����Q������H���,F�Q�+��:C�v�>ę�M��S�6.�֝�*(�Lu��x^wX�{8l�e�'+%;b�J��ň�*<�R@a4or.|.V�#���hk��Q���H���@��I�=��2ِ�]�u
F�9�g�5�
��t������8	�ǧ���q����%����ɍ��ĺq2żf|��E
:�m����(�g������)+�Wy�l9l�N��K����EԔ� r��eL��~<�/D�[�|1����M������%��S�bξ���;7i�'�B��	��u�g1� ���F,�B��/E��JD;��=��Ő��J�u��7리�=t���*8n��׽ב��Z�J7�LK�;�16��`�d�u^�C���ge�3O�a�����{:���H���#	�I_���������Uv� ���_!�;��0�H6���c��EEc�i�Z��t��@]lkw76T��}��8k��V-D�T�/u^���r��#V��\�'&� �",�	�#q����1��l8{@֧��W-�F0q������.�x{Q��5Ԥ:�A4�V"zfui���6f۶�9�,s��eÕ�++(Z�ǶZ��bS�U�̡J��NE�m\�XK��k٪�p�|K�=oڞ����٫aNN�ݸ�9�ajL��Nmef�[�sf;��8Cٔ]#���D�^�g7����O7%��qI^��v�$@"t(�U�	wN�Q�km�B���b��dj]�i�;�O�W�^a�1�{o׽3@d���j֤#����
�q���I�d��E_����U���3�I6[��ttF���F�nۢv����UT�J�7X��?����~M�k��j���QQUA���Z�lE�6 �k8���0T؝�DG�A�?����_���<wc��ؘj���h��t[j�PE�+b�1V(&�:V�����>~?����X��m���mc3lf���
b*j�7��I���:��6�$['MUg<�~?��*&���-�cm***d������Z(�X��[X�A6�m6�^���
-�q�61QE�
�j��6�E�=v�PZUhɱF��;��Z֩���NѪ64cqh6�V�E3P�kADUAL5U;[h�E��5��(�������c�Eq�]$o�ON��_�b/m:�JUh�v��;bi(����pSV1� ��lD�Ճg4Qc�4F6�Z)-�h�ӵ������LGF��O1ku������ml���X���kQ���mV;��[j�cW���Dj('���m�2����7�S��E�е�m��|O/gS�5�OԥNx=C0%:���TLw(�����..���UU_ʀ&�FeH%a P1vi��k4.o����C$�%�?W��
6v���es�Q˔���Æ���ʆ
��tp95<6v�ㆉn|�ݚ5ޝ�(0r�>�	��Oά�гnd닾*�(,��4�1�ѯ�w̖��ݚ�����M@��}`����[�`(Lk�R9���4-Z�o-������f[
��s��v��`��B~a�[Bi�V�@����%xk�ϗ�j���)�R��!��?@�{�Fmw��8n��ɘs 'R�l2�{�ӕ�5-ƽ�_�����$�y��?�zM*���UnQeM��2�{��b_���ۧQa\bK�,ݏBQO���p�Ξu�ߺ�����3;���GY�ѨaZ�K�
�8��K��z/'�d�6�zf\�{e'l�>ñ�h���ŵ�U[�j��fs��U!�H����T^=����
��r����@���u��߷���A�-C�1p��,�0Aaä�}sE�1��&�)^#3r��%���,���7K�R��F�4y��E�˘�s[�Bli&	����Qv�r�n�q
ۨ�s������|�ʲ�q���vx�_7������	9J0�nxq�'�utc�ggx�{��ι��Ѕ�G��s��X_B1�H��R��i��4�.L7|ҵ%��ՕKo^��&c������U�⭵�a���:}��}���f`z`�	�R�G�����������oϟ����!<�|d&U劅'�+��ߏN�ױ��2��_����	嗪gg��9[l~U�͕ɛPz
���H���Є�%���R�&�EP�Ȼ|��6<'�[�d�E4�^�a���>��U�`�[$���������^��2���x�I��44�7=s���;8_�Ζ�龵�����'���x��	���Z/�y&9T��9☮���i�[a� �+Iƌ��k4�7�CK��a҃��%��>��P;�(ߎ҇@⮗=s���d�`�f�WW�{�ݽ�3�l�l&T�y�5�&=�-�������==B9䫪K���+�a�Dܗ�UsI��s1:g����uWJ�s���^�<v@q�"��Dda���1�*��-&�<}��Nܵ�.g���*�����A/r�.��_�ʄ�k�����  ��L,�͓��٧t���͑�u�v�枘f8��ޛd�JbYG?�2џM��m=r�h��ƮG2����&^&so��O�3 �@x�<��yO�����6C�ϯ��c�^�;	y�X��z�nB4]54T�4_o��a}Gn޵W����)���h����P�kou>��~���t�%�t4�lz�2��2�Ec���x�ưS�.;�x葒���6j^�{Vt�#�s7��U�muo<`E�=]{���]��o��]߿������c��wJ�������2@�
R��Sw��1�d��k�mk'"]�pr�Caqq*l��Fk��h9͜a��Ly��noqѧtVent��4�v�BB��NŴ\{��tdK< D���-"�'�zǣ����k��p%l��n'�5{O���3J�3�%�F8}����sN�r����Zx&���B����*!P��sj̞j���׳L��L�`�,�`[|Qڠ��͛OC��P$�`Ḃ��t�
����ϟWq�]GG���0��v+Ӽ���P�&6����n_�x�'�qDo��v����YWxw��;����i�L@�|l�(d��tB	�'�E�1,P�i5���S��A��V)��5}����)ǦV��^|)��G8�o<'f��L����D��z)�r�	�j�`�msl��s�� Z׳�&���j�p�����BR��Aj�?���7�����j����i�u��'"���\�]��	���9��av����aA�9�a�6��3CZ嘇��6��5�t5)���}�-?$�	z��D�M0S����{��M 8��e�M:��H�����4&���M�8/�!��㻝�,3}u`U�4��CÚ��n��b��b��^j��0O!됓���6����t���r��/�<�*Sɇ&Gڶ��O623F&�9�V`]V����T�i�ŉ��j"{7i�
���� $P,PR�2�2,��2RPĈЂP#>��v�3�"}�xd���i��ڞ�������i����^6��M#��#ʯ7:��y��{Zu�4J\���ΪάOH�5��	�j�oJO�kL����|cKw�w���俣��5O���!S�p�a��K�7:/���kݦ���w1���=>� f�y��nx�=��غ���N���b ��iO���vόZ���F�u��i@��#����I`�4�
>�-b_��j=!����P�gh���ìs�mH�J��3s=I|&:�}u�P��4]���1bW40{C�*���C`�?���-�Y�v�uj�h��h���Ԩd_#�ز����eo����e)f��'����A�ș��з����6�ht�w�n����B��p��)HE����=����@fʹ����Y75�CQFq��f��8������R#Lk��]�x��2pAN����3r	�ȫjt�X렜�P%�ZcD���g$��f�����k�Y��/�.3��%�T���|���\:?�����Qm������K�,*�J�V���F�e&:Edud���ֲFdƆM�ä��;��˞B+�<0�g_{��y�P�_�����8��I��ZznՖ0�As܉f�GCef	���q��&xEx����T(|�U��7=';y��B	:P$P$�L�Ҥ��2�@2(R+@�B���������>�_�G^��
V%QaL���T\:��g�[Р�5�	;nC���)��U��o3�������xN��BՉTRa�� ������
�C�������GF���(0;M�]���h�'�vA�n���J�,�$&*Z�KzG��a{��$��JP�0W�qZ8d!�k�8#�d	e�fo�Jy��m�u��i�o6��:���>�ȶ\8�XT��_�u�r�Aޤ�g������������4(�;I�P�+��BO\��7��Wk,�����ٳj�;=ǹ|��SH�ԱZ~<y!��.���V��fÙ:��qTXms�**4]�	���^ʛQ��[�]m~C�9ZH ������01��^}Pq��е�P&.��$�<�/�6���4qf�[�
�r��T��%G0��'[���s��<��!ߚ�>'%����u<���P��3E�vQl�&�4�AXm�~N���KsqE�Pg$��`=��,̩���@�Q�xl_�gx�+jY�u{����9E�q�.�	�nǡ�fN��4:���o�*9}^Sw����k�;ɞǷ�Q��Gԕ�;��Hv9SG`2�eT�|*%r�6MWq�	ʉ-��$Y��\��~]�z/f�����yF,�T��h��u�WͶ0�V,S*^K�ӳ��� ���E���}��E�*J̢� D��*% �"R����������Z�fջ�p&lA/0�P���'z]�^E��ey�`*��#�Xs-F���~�l_o^���}G��&s�`���IE��	>���{k�lcM�Z� �W�
��9���������eh`��P
:~?[�\k����
��F�����qY�����w���c?�p���~�@��?)fP���%�>�[
��s�]��^7�4#������-R�ͪ�%oȳ-���RŨ��/��ʂ�B�ܮ���z�^��[�H��v@���\e4�%��u�J���:P���L��CW���WB�ߋħVR�&�EP������xOOG>��X7h^3)x��9q8�� ��-�����Gc@"{{z!'E�(7E1��&��z����X#���8bھ��Ả���9��7�>�Qx��'������u��*�]?`Ż/rv��r$mn�g��Z�i�cJ:��y�8��P͍1�uL��dI9*IVهC@v�SG+�S�r�u���ʂ�tz�t0N)�@~�C�����?>OP�y}������"��K�u���������yك����3��m�����)�e!�7&�fŎ����5QqW�+K �Uō�����	Z���ҭ�䐔�j,�$�_;[�����w%c+fqv֪��m�t��&^�t^b�,�R�E�i�ͼ�K-���ntPS��33W�(L I�L(R�0���,�	J�@�Ȓ@(�I es]��9�/V1:�1����%�.�ER������=Js��`N�a���H����o~�a�������fSL��ML�J�aǡk���R�E�k%�,�C"�?OH`��<�%�a�b��^��Hryݛ\��L3n=^��+��1�Q����kկ@��1�b�����J�v5�C;Z��,t� ��y���6���{6C��B/��=%�Ĉ��-%��Z��^^�"����~�c�x�4,�ϥ�_���ƃ���Ѳ�T�<�Mm�4M_J�+i��@"A=N�_E��5��~׆{Aii�	��'�=�df��WbZ_�ue�k"gme勩�hvIa�=�P�o���-���R�0j�1a�y	��zi;/�$��:��Ŏ�:�����E��6�y*f�;(2��q�j(�C6_ʆ*����$X�^���?k�:�1�oM���A��\殳u�0���W�o)��J�҉O�WN0�x�^>�lz�t`�#m�"ǣ�U[�t_��``�an���dU��_5��'Ĳ =��4��%��/��^
���_�����M�<�X9���1��A=;�����vq��;�~��G��U}K�_�{~��pwf��B��ݩ
�J�;ۨ�>7��	�[�m�d�Wg��${I��+y���τ���- 4dlG�����u��}U0C(L�P)2�J$�-2"�%
����T��n⩧���gހ|j�r���bB��Ivl�L&
GcH"}�'�=��'��{N{1ګݞ�Xٶ����)�I�����Z�"�����٭��n�����f���f:ۻ&�ߖ���6� Ү/��Rr���(����F����[����C�	�y�-FR�cT�F����Z��jO`�i��M���1i�by�E�u(�50���!�������D�d����+G���8vvZ�����v���(�P$k)zGs���,Ht��o�[��K����:����僝y�;'�C��s�0%��5mw�*���6�b����G+\ײ������3t~&��i�D��~/>�mt^��>����4-Z�,8�X��cS�bŎ+>�3�5lw5�/My0���ޱ�d8/��D��}l/C�����A�_9�\�4�'��u�N
�i�q׼b��p�-���cN���F����U=W��y}u��EuS��l�;h:y�.4ة1%�I����>hA����O��`�?�͝��~x��Z��zY�9w:��:rڗj�S�t�	5O��rV����]�1�w��dz��J{��;kۺu������=1fď/P:2O{j���;���3��>s�w;�vnG8�K��[֨two9�RfP.�G+�;���Ͽ҂L�P)2J4!2
L%*R�I � o7�� 8ڎ��cP�˛蘢�bL�m���>�/,�4֙<�^N2A0��ԟ=�6�Y��&�G6b���6���A�6�����y��Og�k|�A�(��sPd��Q�gSYΚ���d�r׻�M��+nJ�������
y��zap	�9�\�'� n�'7�>S8��xS^�v��,��c=o�^�v��-�P�|��y��#�=?��m�"4�K�WEGl1��K�y.PZ�R�J��ܜjꋇU�g��^Pe���v2j8Ue��l��=ś#�1Ib�b$�D�E)��E8�6q��E�*8�� �5�V��������]w�U�Ï@p��e=r�CN�m�R�p/1W�"���A}������jQ�Z5��0�b�z�5��BsS �y�%�a�n�{����6Ⱥ,㛆.i9���>+��e��E�\V(# �>v��ׁ�U�wI�'N�aU�2����\��[���T�j�Eh�\{5!zjIxwf���!��l�t�17�y�[�j�Ycp\�Wg����fjC�|k�IY��`8u�tj�M�<�GhɓnCWd���c[ݽ��nK
�v	���=no4I�6C��C�3�nv�(�,}p�=F����;W���LPf�/h�[��@]_V(� ��}S��+	tsl��7m�#�-�7���UWﮪ���E�U&I�H )P �0�7����<E ��yo7�����b��"|����h&5
�i�B�� Lk�G6�ZJ�;�x�9��砃�bV���J粠���Q�$-�:�9XK��`��,xk�0{>g"c��:lh�Ȳ��	�a���T����oz��I�5{
T��{��C4�q�nj=��V
��#�:��j�^v�b����tj��ax�7r���67�ۧQaBxvi��d�6k߬5P���+�
�f(�U��4h:ըS>:��=>�`J��y�F��#�.À��/5�A!��9������k�����P�؄[w8鸖Z:3��@�"ˉ��I��Qx��lcM�YX3���V��]g�p��7H���Ӳ���M�Ӧ�`�CzhtS<{a�q9,+ٗ��^�z���ޛ{fgo%���L3X���� �ߎ��fP���p��l;�1P�5�O��8g�����2m������ц�]�t�.�ږ��B^����a4Z�B�ܣ�.�N�ױ��}Ol�R�����^�&鞭��q:�	�^A�v)��B�	�J`��W���1v��C�@ ������u͊B1�i>�;C�2��9�#[�d��L|�����&�ç�Gd��=�XH;�!�GF��Ybk�5�]�a����fZ�����}~��]g܍�`�)y��1���K3Q�>@y��|�~�#�Q,�=�ū'U>�r$V�ki���v�Cy��B����p\-$Q��ڶKx|�f��G��b��}44��[稬�%���|'�j���vo��8�;tNG��6�ҦP�rw���Dmr0���oGe�(�tt*�]{(s�����2P�mjc ��i�����Q���9���G���,�W���
�:�������Ve���ǋ*N��V�R�n�C�`��wֈqɻNJ�Ea״�4v������n�����77��&S������E��S�pF��"��)��4]f��X�ʽ#�#X)j)]�Q�w�{�"�a�I�ն��=�4l�g|<p����&��m����Eل�sfmʱ�g�֘�
�'���+��d�*���_u�U���n��OnW>�Pv� ����m�J�ۣ�z�[Z����[��뼴3XҩT9�q�f�1���]�l��"KՑ[�ު'+��Tϱso�
��;9f�r�g�t�s�QU�ӭ��j�*e���l�)I�&��i�ν������9�o��(��-��u�At��$��IȻ�n�**/a�~uz΁��u�Y�:�pD���W�s�����{lIKA�QU��2@�OV\Jz�TG�Z�Ln���Ƈq��:\������F��������|��~��3�j�v)>���~�����jMT���o���q1���9..-"�/9tV���N����E�7H�
�(٧���r�8��S��L~����ͼ7~:x�65*��)����n15o������r�m��|���5��~��Y�����feSܴB�6$��8n��:ƼQp���P(wn+
乻}�H=t�V�5^}+ȇL�`�q��w�]2���g��k8q�{��݇42��k)��}��Nُ�t˝.a�� Ss=X��N�}a��4��س� Q�wޖ,���yF�M\$�cD�������z�5u�vS3]�"j�����|U�U��$4�B��(��d�Û��֏��پkοr�:��5$z3��EZfv i�yH�����ؽ�MqN�vp��M�I:�{�-y�|���R�<�~��5�|]��2�OOi�&Wh���v@��5��6��2�F�.h�#w�\�{odG'�9����_٘z�\�QB낲]�w�/�L���M�a:F9g�9dTI����w���L�dW���!}k��r݃@9na���))gj	u�؀����������o~�<�PSN��$�,��ȼ��Vk�_5���N�
�ӕ�d�����f�w>�RfM&��2%dpAw�[z���2DB(&Id0BBDQ�&���Bp%�'���/��-~�(����n��MuPOn���?1�ֽ�:o{��kZ�v�Eٞ~�������o�-�T�S�~�˶6l��؊:4��6��d���
(���F��Ǚ����~�ƣ�{wQ4T[9�J������5UR���EUU�UAAF�TU��j><����~�{�5Q�1�Um4�U��8�v�Ɗ�Z��DM3�UG���SV�JJ�-�R�D�����?���O孱ht��Wa�5U�6�A[[;'ѭ5њ���v�Z��;b��kW�`��ƍj��CF� �vִSD54Z�V�kb�f���^�lMPM��8��T��U;*뮵�N������Z�:�1�P�Q~l{��M��"*�*#g�GN��X;b�ֈ��E�TPF�^�%�{������DEl��1v=΢�ݸK�F��"�Z�Z�(�:;oF���UPA �O�1C����krK�K�ނ�0���`���Ʈ�<�cNI�q��S�3�_!%t�̩ԙ�tP\�G�m�>�������( ����Ͽ��id�&	�&@ �MI�/f���&�5�ĿQ��p$8����pB|� ��5����Ru��K$�s�lؤ"�.}y	�eW>o[V�?������?��,
ɹ�����K��=�"U��}�E���������T��q�S���ިn����k����@C!�3�BxBj�L�=����K�F3��x���qd8��WKаXE����/87'a��-�l;�����j�����^|����c����TvG�;B�Ê�K#��]*�^Y�KӇ�������R�ɦ�A��jӬ��h�����c�:����*��q�\�⠗�{��Գm�`�yIu_%�$�������)�F�u�K�쟚FL3n=�E1�AT��(�|�#>�}�2Y+��¢��	p��k��yωχ��G���I��{�so�;���܆�Ed�~�1�I}�-vݙ��e{gZ߸v��Ej�^��-�WX�e�ޘ�����bT�{j3],�A�u�;Q�h�z뻴�i��D���y���	���<�Z� �鮬p����a�o��4��&��5�x�N=��W^����ﳝ����o>w��T�x�D���a&�NW�*ޚ'��@� ���ďՎ��T�0�$�4��IC�����[2�$�ްwN�0�u]�\�E�3�;痪*������9�7jSŤ�����Tv�Ff��  �~ 	�B`D������`��� ��'��������hsf�i��,:��^f��)>sͼ4�ڡN��y����������ں{�Z���t�f��z���8�rTͷ㲃%�l�!�l�zǫxGh�>-� l�w7L\��5C�a��9�Eǥ�`�cϻ��H	���Pd���{
�q�F��__����+g�3ݣ��1֝�����%��@$<�v�#!O6��A8�Q,���x)�Ǹj�V)g&}Εmq�8���,4++�R��c ��"r�i�����vI���::�G�3��Kv��<�n�"y֨Ǽ������������ �5��JY���R�_�=��d@2�2��K\뻶�a(mɇd�O��Rr�y��-�a�^=]��y�s]��	A�F�̯�y�,�[8GXP֦e''����0��0���q�O�(q@���#�.�a �g�:�*F�3u��GeE��cf��
�
�gb�gc��k���ݦ���E�H�R�Tts���v�$	�Mɛ���ߗ�����we1�;>���p<ò~5�B�Չ2)�&���7�|���}=j�O��˙*�u�F��|�/����w��X���wY�ݡ���N�6>ͪ,�E��= ��>�k�ݸ"�����;F?�f�ɒ�R��׸^�Ci8}6Ƀl��T�/j<ZD���V?>sg>&�V�f��S$N�'��1��D��*�ȋ2�@� � �g)m�ݕ��>���Kk��'�k ����]�:��:����q�85m����!�n�����Nƫ�%��gն%W4���B�v3�~g!�����]��c-MA?�r�6;�����Pi'��Y�^��!/Ş�w����|�Ph|Qc���w[0[�>��m��T�\�,yoP~yÆ��48�ba���$�,�sͼ���Zۘ�=F�:���ٸ�����BEų��u�Ӎ��=�>�yf����'���N2��m�����
��$ȵ�8�ȱ�~���ۄC7���_>��ƕ��q^975�C5Ocd�ĉ�Jξ��w��Tΰͱ��l��9������>c�
7 �����A	��Zg�:�u��������u��ƀ�.:���Zhe;k�l�|<��a�!�#��5�oh��e����3�3���.���^S�媅(RX/S�\[wT\:�xS���c��M��緻�׻�o�S��ɛSӲ��d'ry���L��xY�]⪅��E8���a#ݑm
�q����>��x�>�]�ť֎Ė[���s��Uyq��r�E �.�~���{0B1�q��f���
T`Yҥ�cSސ����q�?iG��{����rՁ%�vq����q^�n3��(y�8���R��;8>�sT[�����2��뇦�+��e	�Be�&�Q�� h�Z�����7��8�Ct��vA�۝0�7��e���_<�/Iq�o�Ӆ��-��bl���Q�k��]#�����Yv��}RS��d]ax�1:a@�5%�r�ō�$^Jњ/g�>�<rXt�hcm�?�z����"N��&^�+�"f��yӧrk��w:�zX�2�Z/��ٷ�a�`A�|SB�y>S��=WB�sDV������.]���Ar�Ν8��l�E���1� �O��aVs8.��K���Ʊ�\b7Bv�!��BՂ��6��z�O���Ts	m	���?sp_��A5oƞ�r�8����c(\�jY��u�R�H�k�C��{�KsP=˖��Ig�X�涙��ŝ�gP�t��{XS�+~�2��'V7�ۧ�r�
bK�,ݏ\fa���c�s�)��ݯ0c�������-�����*j|������ޤC�w�+L�C�]sz�����ݭ4�n��f~���~�-3��	���;c� �%'�zǦ��Ư
pI��X�tU�]�<����������z�����=}�B.yj�ws*?ϚǇ1m��h�z�����epK�Z��֫���o:JR[�I5*r�8t��go���_�br��a�?:�;�����0�+d�Cu�pfH�mީ��v���_�
A��D&I��?>W����?���?���(��FC�|�Ε�CQ5曍�MC�.W�)������w4]Bց�\��T�%ZM*���j�R����Z�㰃#�B��G�=�Z�!��g��si�M�Tw3�g��}ǆ���298ܣf�GB�/���b�)�Wm�Ӻ��z��a�*��+(�(�Rɑӎ$�P���W��=x���Bc��Ju~*SΊ�K�f����3=��زkc��k�3+I�(���Ќp�8^�W�5��.x�K�]�s��'���9��x�}�b-k8�aO�|��`�k�@3d��L=�K��=�"U}E�j����f"p<���Q�Gb�~`��O1�xn�چT�zܳ0nv/��2����u	���d��E�2�9�T��gx�Buj�*��WK՘���T4�L?5'�`>Ϙg���M̰�Wϣ�u{����_����ħT����h]�*�=Q��ʰ\��z��.���w3���	Wc9ج�����X�0>��S�����%���XO��|���{�(�W0ͷ��:��Wn`TR�/�z�Ag�XV���,VsmCV1>�s��[e�7���V��ogX��ڨ�u��/�_���7���H�~ȧ�@"��p���B	�Os�ӛ�:��R�l57k%*�6 �K0oɆZ-_Rk��j��k���Xp7��y5�+�7������@�P�0�0�0B��x��4y�Pg�T����0g�`;�%���O�a�q����9R��2����3��~�7��8n13�<GN�k�e��k� <1���p����<��{P���͑~��Δ\�u�<�ۈ�*$E�R�XD���<tE�j��g�]�,#�C�p���Y|��f�Y����:�ū#o8m��A�{�)0��i�C��<'��R0yh��n��L��?g��|,V�.��g,c����w�TQ{�᪇6n)f��è���d��3b����:��h�v.�����We���g���Э���� �##)��z9�nL�.JY���A���rC�E'k��m�UP����Sb��7#a]���|���R�A�<����U��;���x�M�9J����_��#��b�k�^�G/�st��}����|��I���$�>c ��� v�#rUsP���}pݭ�O4׉GKf�-��.3L�MN�om�L��=�C�02@Q%ٲ0]m ��e�'	����j{O`߸�/�䟖��y��V5H�4������������l��3lԸ�ʜ���xٝl&��s�ɣb�P�=FMբ�������	x����:���Xvp<7��=���oY��4�
Aq�K��tw`�h&���e�Q���/�b�����z�����̋�K���uG���)�y�j $�}y�Q�lֳv��>����д L�R,�"�߯�z�Ԑm.��_S�]���7�RO��zY9Y�"�ymsj��|�>�h���Vŷȴs�3kû�u��߾P=9Q�܂ҟN����xŧ����p]4�c+y�DS��d�z��
�t��/01�0�s���Z�6�i��Us^E��d�iU?s��h+:�)ޝ��ڦ�t������"[PGSCE�垖#%����<��L�cB	�k��)?3*��]
q���^\�'<ݯ����9�ƦY�\��$�d<���)�4u}�C��[C�еϪ}9�6��W�Ѥ5j�����?�:z��-��t	�4��cB����9��o��,�s������ݩRܚׯ�U��pl23L(qh����~��~���H_&V��9�=��w*cF�\�D�W�#Y+ޠ��	�]���c�ĝe�y���0�Cw��rR��;�3�[� ��9�X����YU8�nw��/,�4֙<�EN2H���l�{k���-7ig??j�-�dS��(����Us��ͬi[	rnh�M�����s��l�	|��k���c;���]�yOz��:I��ۯ������+��L뎁��N�e���#yn���{�����BNֲL�x�=Y5���O�OUƈ����ݜ�^X�,�a�K{Y��<u��l�W�[aQmpz����~��S�ee`R`@~}��k+d�n�ݽ��͛n�dn�(�,54k4?�S�Y���.z��V~�5�/,�5띪h��!���Ș!=,�,h��g�c����j�3G�"�<��~���M��s��W�T�[��=���ƛ0u˹��<�(-T)\�,���.מf�������<ъ2��?G׺����ھ&|#ȏ	�><hs��=�)��-N2��=7E8��l�	�d[B�辄�dNȺ���w���!Qm0�!�2��.���s�w�Re�/1V9�QzK�Ye��-���=�np�5}%���H́p�i�!?T�"�����xv��꒞x�2.�VC�>il��~����ׯj��X�Eh8Z��Cw=	yO�Q�F��aY٣���)�4T��0�ڏ<2ι�������d|RD��k,;_�6>=��ק�yг�k�ꋩ�[�U�[��Z}�:�����<ƬR�`������n�`�C�w�[�v����]��t���]HL�v���<��86�ҹ�rUO�>�O	vs3[�|�C�|k�ܽA�9�X�!�#'����X3�������ʲp;*�<]� /�r����{�]���E�Ӏ�	�'��RQUR�d�I����R�#�x�ў{*����p��y��ػ�޻G%���4����d0z���=���������7���k���S�eY������㬭��cL����S��?���΢Ú��Vy����;�^�5-�^=˕.��QЮ݋ܽz��ʾ�[�r�Bu0!�42��<A7t�#'�ך�e_\�7��{�;j>G&�n���ǘ�v�|;y��������[:y�� ���k�R��>�k#�ާax�^q^)sW�eS.�k�N�p��[(�4-�4�=0�tE���6�Ɔ�Hv�
ȡ\O�2R{��Ƕe��=1�"q���wH�&rղ��\[����B�My��b�4��u^�xX4�S���q��G3V���FK��-[0�ǔ���2�,�l�����1P��3�!����օ�]��; ��i<�5�}�8���KsPJl�2%�D��+�����vQw9#.j��s�t�*��\���0t[HN$�W�BGex��v)殄%1�10�YR�'Qs\u�|�}k�i�{��/՞ԁ����|w��ځt��L��hH�5�脟�K$V#nU|�f��fl��������H�aA�/�5�B|�֐]���Co����={/�g2�*�C��7������uC+�N_�������{i.�lY���U�^^	�^7�۸���fn3\��dQ"�U;(�G��,�A��ڧ�����'��)�}ޤj��0�[�)��B�x���� ��Ǜ3}��o΃�MZ�on5	�D׾w׿����>�Ʌ&D�)�?�����?�����~?���v)?0�q��#i��ިn�c��PwQ���N�|w꿈{*$���ޝ���k^���ɇmN˯Y�O�~*]&���w:����=���8�]���,�[Tħ��J`Z����%I�>�Φ�P�z�&#��ۇP��v�)�ӣ�󤊝t �s��އ������%��)U�+�J�
�^��8�<����t&x�y�����)���[�~�s	��j"���F��Z'�e���r�O��K(�{��̹��k]ka;��xwb�㠺gZ��e@ņv3���?��P55g��~]x�9�n6�Y��Uod�i�݈��Q�נ���Kϰύu�����CB�!�{巼�ar����sz���ʽ}߁4������
�����Ԍ��Є�t�V9g�9hk����J�'ņ������=1ש1x�sz�4��v��d�U�CQ�E��z�o��ɛu}���}~��S~�|<�0f}�R몟�*ܙ���*f�eTN0-E����<�#>���2�� ��\���V����p�˦e�ە�b���썂��}����&-|y��7'�kg�U.>^�=���5@y�ef�-�`�#�"N��w�łh�ud��G:n�"7 �j��o%�u(�Q�NEk��h.��]��'6�ta��ʤou������bi#.-�/,��l��jx"ʥޛ�@�e��o�十�'^J���B�y�4����	b�ͬ���-��Xú�)p4��m5n�v$�]M����v��� �K�	'2Q��̗OL�g���=�51+�{%E�z�Ǵ����ONY+:m�����B���՝�q��dܲ��;/��Rx��5{��Fݞ��f�;�4������#��4����co�a��o7f���2Y�f�R�b�9f��!�Yf�4שּׂ�3�0s������"j�i���,�m�r����r��+�Dٚ,��z棛��"5�+K��$v��4�q���G.��wE�\5�%�[Ʉ��Z������º��}skpd�ojX�׎�IgL:9�gw���5˸��-� ��k�8�jnӡsWh�p��:-��ɣ��p)�(��,��g��3|���]}�#ټ���(o�nDף�wuQ>�<��ϘC7�u����q�\����>������;,G��B+�
�3��?3!�ቱ������ܣ���zoU���xa��7Eˡo��EGV0<���ؐ�dt���"ҽ�سl��-��᪲Rf�n*�r���)����Ut$��0��A�]J���W8����whWq�J�βhG��Ԧn42wR�])u�:�C�q��Z��qAm�$3闵(�KP����+3����Rx�ʦEvꝸ�F��ݸ���; }����zn-����$�Z��[�$8��z:L*֊�.Vw����G���^�j��� ����#��;)�5���QQ���ܮ��Eٙ��".Șq�1�u5Ʒ�OjL�+u��O$�ûL�ܶ�"�cӹ' A
�poQA݋5؏Yx�X���4�1�G-�Qe���n��{%Z���� ��ku���*x�X�U�_c���<�¦���U+�D��0�6ۻ�rv
s�ŵ�\&�_�5��{���d�l����� ���a��t�w�%L;�]�jqZ��]nc��X��}��o�pL^�����k��HS\o;����<��b`rn���{�vy6����B�Mbm��ifg'��=�4�����!��dV��J���ݹ��B�<XN�:h��v��\\��;[�Y���:��͊%�4ɩnپn��ڵ�~�-^}扽�C�ؙ��)�>�9giVITmY풍Ŗ� e+r�]=�I`<�j&)�[u-��L���θ�7v�s�aZ��K��On�����y7�/#ِ�����߶_�eU0�G�ثZ��환���ب*��DUETM5t{�:$�ǟ?���z>h4[s���*jn�:Z6�F��T��g�ϟ���>i��m��1�U�E����Gm֘���d�u��m3�����G���ֈ�&x�-'Av��E~X�mzz�:#d�%$�y�~?�ȣ��1lb`�hh��EU�v;��hݛ��{h�H�"(i�4ӬTD�D��n8ꪨ�**�6�Wv&���"Kc^��D@UZ1Zq1,S5�ETGki&(4h(-bj�ӈ��&�F��&"u��$յTv5UGZblh�TA8�!Ulw8�Ʀ�&��愊&+a��^4U0�h�;�����U�M-����Emi��]tP�R���|�
P�z��ֵ7f��a�2������w�q����+e_b�n����;U�`�R�c(�w���� �0�3)����;���Y�Я�}�����"���`"��y.==^UX�+���sE&�⫃K����J>��{��o������o�$e�S�|��i��:6z!M�<���"�Us@�|��kۋ(�gC��\9�ۅ~=~kƶ7����N�t��<t܏bx.�zϥ0Wu�����U+3�͏ʼ����DIt���tuH�4�����ܞj|x�u>������x���q�]-ݛ��c�jBa]��vJ�7��O�"���J���gS���GcQ�
�T�N׶�����O0"C�"rp���TCS&��q�O�<�%�j-#�9��1������2�F_B���,���Y���xr�����G�v�\n�E�de/VSEJ���
�F��%��ck�"a�ȴ�ь] ��kXzdO:�X�յ�NW1aU��ݻ�d#�����z�S�U2͚��͸5�W����(����u3�].�G�ް��l�]�z<�ĦLcYk߽ǧ���=\g��_�Ph�������x/���a۹�ǝ�3��;������rC�u�V��ʶ�s�,m��7Õz�H�k�˟�+�ck�ݶϗ��SS4%�(	T��F3rf�Y�TA[\�cUDb���gc��=:��aX�P��b�'M�(ⷵ
���5�廾��������������L�L�0�o7�<7��B7�i��nR�o��2uڤ?vI��ȁ4����A~��=!�3�ٔA�}��J�6�u6������`�>����{=BP�J�0�X��q����S\��e9z9*$ޖnּ�5d�w���t�	:�=0�Nx��^Y�i��O;P*q�m"8��q��B@y����LGoB�@c����y���%�ǰ((F0���E���כX�] �(|X���l�<��j�"n�L��$��8��z͛e�)�?4��'$�ُ,,L���+�IN�>�ƃ�^�2[ֳ��zd	bWN3鎷Ƭ�����dd��X�N2�.13S�ʫ�+e��W�Zܩ�����F���\����R�%���nN5�뜗W���.Y�P�Z�C�W��=Z����n��]�r]���-���r�	�"�U���L8�����e���8�=�^��}��~��ٱ��_W���&*��Qz\��L���{z/�i�i��
�9�A�-��@��i�!?W����˰�5t�O=���A8_w���dg}i�[�xs�:n'�!���i�g���¹�}}�$��)����;b!Uۏw�yQ�"��ė�2�ݪoN>�xs�����b��N��&�ev��|�en�A§P���ڋ���7�grtN�ݛ9��[olU����2��
L)0����[y��+�maz�R�O�Z}��׶W*���~+,|�T���%�?P�p
6��F����}��K�;`�XA׆^9r���),Qن������ ��!|v6>=�~�g�4>w�l�:��K�WBչ���w�<�����m��Z�B{����1����*cU�d{۱�Z��dքZYy�T�m����MV�V��zW=�����*+��m��{��]�[�V�n�'n�)�	�3��g��:��R̶�u�0�@��6��P�9^j[��n�g���Y����й��u���6D��
ǴBax���ʖd�^��t�Qa��^yY/����^�V�����_�"hv~�(��^����~���5>XEV>�~������7y�13�C�q�^Q29I���i:"�P�xc[��>B,�y�c%'GI/��[�ӿkI��:q݃?4��LW��'�f,�@J�PDךE�Ӧ�z�\�Ͼ���77Wte;a�LI��\(ۚױUԮr���.R��>A܅�B�Ru��ޜa.:h\\�q{�����K8ZNm;����^ދ�_���^�(��e�X�AO� PF���]t����b=&U�s��ÍL9t��4tf��l�ښ.�$nV����sv��Ǫ���`��3LR���P<[��p�Ro\���;�e��5�;0t�OK��������ȢEHOio�w�{7����F,l���q	�qN2V.���s_A�o�H,�)��vз��h�|��{yiڎή�����ǆ�|gh��m�!w�w�! � �殄%?��x��G!�mD�?���n�����ũ����y 5���ʘ'�v ��v�]TF*�&��Ֆ��f��nN??�]�h[�Y�z�8����1�N1�U1��[� �6\B`��n=ݨ��{,�ݭ#��ņ�<ي.�X�R���oE1��P�@��-^w������5��;ǩ8��m�[]Fs�HP؄�L��:�iC��qWKг���T5��a��'�uך:�Vp�ͫ�#�Ǻ��7��P͡=�3�r��uI`X���Uz�Φ�*�K s5шm���JyNe�.�z�á=�z,9`�_��ֿW���U�mų[+R�Xq�Z�?sԼ�r���}��y�N��R̨Űu���8|B8����d;6���M��AT���*Պg��:od���v\�3�ǡ�8�-a�d����;)������F����˘��ؐ�K�'��/���8F��k��>����;��s������y�^ً\&��,������2h�Zb�!+�XF��s,ZۜI&������Úȁ��k�gsʪ�Ed�a�����0��[:;s��{�5��Ʃ����N�|�O��� Ʋ�	qv��~��п�#232 o}�|�O�����������}�����G��!�^�b�'D[��>��O�Cyo������u�(wc�I�u��2�3kCHނC�"ǩ��_E���P���]���v:��gt�C#}q�[c/!q�>��I�z/�oP摛����$���YO�B��pl�sLm�f�)VP[�t���xihgV#ZP0�c#)͊�����Ͳ䥛BMŰ�5ģ�&f�fS�b{za��3t�C�}�5�ur�f@��t1J�7L�?){`�zv+��BkT��K=�qgf.���;��3i`jd0��s=�A�z��[�z��  �d��an����6N�F�iL�6m��u��Vǋ;�b�C�!q^�Ƚ���+�&���|�=��:x-bPy���N8<����������§Zh�y�tD�I��Jsz�SH�kgێm�p�<{$Z���
{ +���������������N�愍�4�ሤ�g��Q���9��a}ľk���]3ZS�t�/9�(�b[�op}��<�^��0��tڞ��-?,�P{ȁ�:�}�y�ܖ��>���2��0k\Q5.��5fuDjs8�n0Q*=�������������4���{�讀��X�NϪ��(%V�����#X�K1�����C���gk^̧@s4�.}F��Ae��{���{���-d+i�e�\��'J$"��+� ��=\hf�8�vt2��M0���E�^O�p�0�~e�Ck����W5�E�mP��Vf��mp��-�]yl$�����$_<(���t.�ߪ3��WU
�W&E1��� d�a�4�>�m��75Kb���6�b��TC6k�D�� �ฆ<y@��������j����f��
�C�ƅ��qf|e���t�[s���`_��Ph����Vj[�Y�uvYE���v���<��A��I����Švqy���-�W�د8�=���m<U:�lF��p�(����~��ڃO��́j���{��2��6�\���K��~k�k�����yy׺�[���V)⨘�{Bzq�����/,�4���Ԏ����4�k�#7V�@9ꖯN0�l�֋x5��)&<���<!�n��RS�:�Y͂˼����+����։1��W��!�g
��O�,�C��Pr����3�偬Ǧ����t��2͂����A��X=4�\Ɓ]Z�@�[�d�C�-�n��ImE�Po�<�����׆���i+�뱌����@~V��eI�YT��Ϩ�{<׀J�cP/�b�����T��:e��%d�}��v���<>�5ӝ�l�y��ڌ| �#qe��-X����ƒ@=�Ѭ��m�,��D}�SX�+f�}�~�{���ؽoGoK�0�#23(RԘ�0���|��s��bm�F�欘\�:!Z��S��D�3�%����t�C�mۋ����2kqY��Tΐ�����n�wd���	�{1�X)P�r����3}��^-���[��'����샞��|�6�<�7:3�*S./1U�98/��*��$e%�o�6�gAX��/N�o�i�!�^.���;����@)��l��x��.:8vB<�fۓ��G;��q�h{er���P ���U�k��*o��y���yt_<�Sr����@j�¨Z��G.Rz�Tߋ�G�HI�O�,V�ð�ǲ}��+k����j��c�<�+Ʈ��d닿"��X,���>�G�+���Z	��|�Z�����ڌ]�|4�9�;s/@�Lh�9�i�i<b�,zW=��%�ң�HhN���u�E���:�U�]��Hw�PX3B�𹭩f[C:�jR�o��Mc���r%F�f-����ҟjF�g,ߙ�|�b��+zz����?�a7���T'��7�=3�^#>m�)_-��`��8�4�8ƭ�P�fge���1g���sN�Ky{M�������'2;8����m���$�s��=�ƪ�~[7�].;�eۣ���bí͘�Jv#!��)��ã������� �k)N�KT�*pDN�-z�}���>�i���t7d^E���������
(�� �#˪��n���7�j��~��#3��Pŕ�5D�G�k��g���{g�W�nq��8f�ϑ�f�GYi� ��׫y�C�����I�ʹ�L�P&�`���l�ܭs껠�F�k�/��ԗBj-=��i��[���*��5��׮v�5wz�%��SDN�>,薸s&8.��Э�A�8�sI�1�lNT��2���R̡Fң�z-�u�2�`���g��s쫇(�)���7��'#�z~��g����Zd&T�P��x�T[�XϘ���C;���>�LՆRf�YG��g���$;'�7Z�nJc&jI]U�+m��\��oOSf�y��%�j�U���z��	���(@>�M>��О}��-��&����E�W-nѺY�o�Y2���d�`n�c@$i0��p�Q	�k�D��1	���;$���r1��S��\�%W��y��N���ʥX<P﷣=�ϩx�@�aL�m-0r�W�f�Eh��Y�>6!0wb�'N҇^8���1i���AcAt�~jN%�G]>�X4Y������1m���L�rz���z*eKxk<���l��ν��yn�Ժ�`�K���f�f	�6��^�� 9�Y׹w�B��X;�����L��ϔ]��^�{��$�=��h��T�� ������}��S7��f�����̺1�;g'g���{���y������U��2�N�|���9li�!�BbS��K�t��*�=Z��Sb�眳Y��S��ٛyzU��3�*A;��-#�������;�I�F�ǥs���ެR�.�W?sg{ت/�e��\d�s�A�Wa?���!���5l�7k��n�G4���-um�C�תX��
�,>�~1��z��1a������<`<h�]�5�YGU
��+�T�fԙ�4rj}^���Y�_�1�Iz$@��:"ص��z%�r�$Z~x��,�͋�\�4#�&8�Q��g�d��Ͻ��Q.A&��c����sWa�I�Y���7���3j��r��L=�'>�Q�����C�sp�4�Aa�
�R2a��Mg�eY��=X���9��Ы��� ���
v����X�/`���=nL�.JY���A����ǎr�j�xfo�E�{���/�I��D�`B˰��ǧ�Uc�N�{1.u��Y�:��A��I�҉N�b��x�oV�^�� �|�CDSw��,�,�"�l��3�:���{���� =٣@1�x�CI��|P��S��x��⟲	��bq컉-ֿng�Oh(vC���F��AR��ObY�����p9Y�N��)'�
)�U&v�Xk�{��G#�vD���= �� o7��4�ovy ٓ(`�I��bN+ÔK"�R�er�&�-�F��P�t�)��$p����:Vn��ɾ�9t;4�LpƀFvJ���'�b% �Ʃ�XPH�lk�nO3c�:��Z���D7;�5[��v�~���2h���OP���vD�Od�q;�i'��NV�"�-�a�Z�{���(���v��Y.��<�-��!f�yЊm�0�kq��Q}��[m����n~�6u���"w莝���8�|�B��h~=4�A��E�3�
5����xeo^����U�{D�����l��K��5���I��s�}��/�C�k !w(?.�uP�_y��W:Ր���D���(������d�浦M�X�>��e�+b�ٷ]�W���?&�OpR��Fr9m=�ܚ^1��2uڤR��p/����O�o�k����X����rυ� �1�����(h\μ�S&���'ݮ��v�X���,��\b���nZ7t,cB§o����������(��P|Q`|&��ԍd�z��ϰ�5�3Eؘf-����N�o���Z\�VGO8�XJɘ/j��XѾ�=�Fj�����S{l�xJ23�]�y"�u�h/�.�o-�d�5	f�͗�(�id�������<H׵d����!�i��p{Oش��"�g���,�%��~3�ǈ�7\B�͎��s���x�� �����X�uE����x0�/oU^n�R�꾽��!)�!�<meӔ��G{�<� �������V�R�V m(�P=�b	mZ#/�Q|��"�BQ:��ҡ�K��5���#�wuն�%����j�}ί�l�@]
1j�,ܘ�L��#�߮.�ȸ�ӝ��[κ� Re�ed.m0�ҙ*p�0A���1���q��s<�;�ڡ��z���k;�W-������|������F��V=Ӧ�P�����s�ܕ�6yη��bV�\�k�+vhI�y��.N��B=�/qR�J���M��%�g:�ƯiY�����
|ߝɻ�8��֙ӛ�2*��Q�بW;} [�+W,��6��S��z��iw�@�yj��H�=�>�l��-Ou�1�=�ᶟ%g��_��@�Ȩ�D^f��*�{�0-j(�����L���	Z���@��C�sނ�1Ϡ뫦+=[ʱ;�5y�d��v{Rx�5���b���Ę �Q�ō��MM���<r��\���e�	�՝�̙��5r���^�y/��&�b�A���Vs�28�|�Y�r��ho���t�����L؀c�tG�=�(7�5'��}�%�0hU�gx"�I,�K4m�%W@����h��7���F�a=�t@|��4J��Ÿ�臹����p�;���q�	�-Rn��c5�un��s�K��<	u��-�lׅ�
�z=L�$��9v��|Q���F�Ho�D��~��\�l�61>�%"�Y0ڽ�>��Gxbr��6*j��k��{���j��7��TeWCs�Mly�J��<�.���ޏ����6ZO:V�X��؎�ۺS��3��ݱ����T���:�i��`zl�Vݩ�C��+/��r�����o�01F��x�\+}F{��X/4'9&Ug�Y�#�VMT�͢k%#<@�֯��m�v���]�F�^�Ӻ��b�Wc��	dq̻����[֞��Tb�����Yؐ��q&ve�n"E�&Q��e��Eud�"�'{�!iS�&;-W'�U��=V3�WZ�]�quVP����R��/�6�M!`_?�=5r�VB�w\4z����^��(XTOv���f�5�g��讦���Q�j�^ѡ˟^NAK�G��[��37)��1擡�^>>��Ƕ�螷�v���K�J�h ލ��h4vi	rgˣ��~��8î��R���=��n��B�|�x��ӗ�Yv��6p�,���{{Z��ˠO>��1mF�+2���skr�vH�k�	�agW��j\9Q={�$e&y��*�۹�����/gӻ3�0Q[�v�c^�k����7���Qt�3'�1��n�-��v%\�̍Q6bL��`��p$��$qD�&?f�A���j"�:����1h�PVآ*	�^|�ߏ|־L�Ulb���F"��4�-�`�#�bj�g{&���F$��s�����>E8�*��;��.ک������z���u��Ӧ��؍bӧ�{b=j��]��9����~|���3�Ӣ*��i�mU����ئ�kquq�̟�u���EL3�����>6�3��b*5F4~I�UULTE�稉*�j*����F���^�gElk��"��I6sQW=��0kv��ثح5�f��v��Qh1�b*�����b�qFǮ�^���(��M5��{j��U$TQ;:Ӫ���j�w:��հf���֍�;k�z;�gPu������;��E&���G���~q�h"�w��ⶭj��QT�Qh�N�63V�!c��u�D[jJ��5GZKݹ������*��$A ���#TȰe�P�?wR���~5��^�/0k�:;��*΋��ܽ�`Ӿ���gE}G)�ɪ����-k7;uvĹTKA����"�E	�	���;��ʹ5�PǨ��P�-?�`�x��o�q�_�et��s��=��M4Qng���WR�W(Ӳ�8�5{��i�Z��E<�����$�<!�v~��٭>�<Bܦ+�����V��+Ҹ=�3v��Ax&ɒ�Fq��f�c�gO����'���h��}vבgSf�7���c�鞐��"����t��|��Euk=�;^s0��!������=�����f~��ual�F�"PB%>���U;H�Y6C�~wA�:��Z�B��TXS-�������IDn��9*��{���#���M3]����fK��Mͽ�'�)Ք�Z֚��z�yMa�Χ��j��4��v;/����~x`k���m�@�۝���T�=+�CU�B�7ұ�m���/"��Ɓ�8^�w�xa#r�i�'�pG?[�e�4e\Q�����r�z7X������T��eM�.�y1���C�+���P��C�R!�n��&�r+�ZV�9\Cj�|W[B���XUz̮xj9r���%�v��	�|�D�Ʊ@�øn����y��X��-� ~�g��ũ؊��w�庀:�7�5�E� �z�Lt������y������Dn�:&�:�ߧ�x�>��>�d�Ѫ���\b�����>2��ýV;FS��s�-rɭ�i7�0�=S�j�}��u;5է ��R��t��?<�o7�y���{�������?� Q��U��5t,�s'\]�TX,����������+AT�B�8~��>�v�_
�A�/�)�,ZFHS̬Ԃ�GMV�V��cҹ�r^�ʎa�����.[��ܾfZx�yŋ���pcD-Ƌ�g��=�,�k:�j`2�},�=���*�S�ؙ��62=��{��*���&4?�)n���	��7�ۍ�;������[۷�0AtIv�d��@w�f/�Y��c
�TI��y��g�5>XG��TW�/����>����s���@��/5�A!���L1��~�9�L���V1�a��=6���^-���<=��}��V��3^����A�VHA>j|�M��'�'e]*d�K���ߝ����~!�ڄ�ܮ@X��=^ܩke����PY�P4��p��{�3�U���������(y���)��mc��È�i�8�\�K	���,q��P��rʲ���}��yғf<�^�x�Z�L�Ԭ��<����C��j��;�g�h��Գ7�,�S�z�z�ꅋhz��/tY�3z��a	�*�dq�ʶw��Ӹ)���=3L�Q�#/лЛ�N3��p���"%]O�͌����m�L�#��S��{�Y�����ެ�*W��B���1���k2�������1�_��W������΅q&�C�B��r'�_���3��V��1P����& B������!C���*��͏�h����2S�/�=�tS���Z��a=q �5�k� a�9�:n�p�"�	tO�B���]0�0yγ�r[�:���-N��{b��qFᵍ�2
�aD&4&m�ΡJ�҇)�~/I���,h.��؞_���r^��gu���,0Q�g������ߏ4�=(�����nՒ+x�0�-F���*�.LX,�v-s���"]Y��Kӯ4H;�xP�a�ã�k��M6�T)��6®s!�ՖDc�-D�h�]��u�0Kܽ�c�l��vB��`���S����(���~U���LUȔE����6}�"���<��uK����[��c��9�3�O��(h��/]�;�Z��8NUѾz~Xܥ��z�:��C�����lc�g����	�/�����`jitg;�X�s��Uh\���p�I�罨�GzC�a�a#z	D�x�;H/���&�:g^47��ܲ{�P�uJ='����L���e:}��5%�!�]#����n����N�C������ɬ�4�y!�q��$�Y��)QU釘w28�ހ��jpV姜Pw\�z�\]�ƹ
z��o/"ƀ���Km��^�NHw�Pwgg��y�����x��;�6ګ��xr�S� B���T�՚��W^�oW�,�4�d��e��7f��dҼl��ݼ�,Qj� sM�6S�<ZZHP =ŧ6*���^ܙ���S5�\&��i����n\��&�ԁ����N�z͛O@c�:��)�,8o[�d[����QL	�0�R��T�s��dA�/W��,By��A�U���WN0��Ƕ�x/L͈("�_��y��=f������!�cI�f�C����'���D �W�D�/c�)�W(Ъ��Ưs�:y��Ё���q9\�D���/'�vn�,Ɛ�d}Sd�����R)��&�}����D)i���b"�-s�T�,��c�C5��2�0�O�ܻ����J�|!1W�"�lM1~z��nZ�������h��T?�����`/���; ܑ%�L4�@�<���t�vn�v���
��;WyA�{��p��at!���7V|G�x�A����'��� {��7�P�h.]�-
9^�H���=���ǫ��mu��*+Cb�q�=Y���p	K��<��B{����x�!&L�5��O����:��3ۇ���a���g�t�c��vF)�M0H�k��	�P#�bEqf�����+7/��Kk�	�2K��{׷r�q��{�9Dw���<Ȇ9g�^J��1Gn�7pב;Y�U,�����`���a�D�ב����4Y�d&�c`K�����&
�Ξ/V)O�T�6kӻ5�v�Ai����N�����oe=�_�.�@�'��UVJa�Ʋ׾=>��;{�����.�N{����5�2?<��<���1	[�a�o>˲}�24�I��]4¸���͎��Q3��۷U�����r�|d�w��-�_��H�`3���ʐ�+ޠ��o���S�R��<��m�k[��,���t9��.4WٰE��|AB�!�_�k�W��s���X����3yX���v�&i@���IHA�#� �����6�v?�ǰ>B-���E�Z��:b���Jݮ���C�n)��#�q^���[�����qL���X08�n�b��ފ<�k�!�ޘP>���N�[Pބ�X렜��%�����u��y�3�E~;9۬�w����=�v@�2GDM�*k[���P��dG�B{nscR���+��S7n\�����wqWg]t����mJVS�z>Bn���V�pΙM�C�"�ϢS�Rw�����/�g.LV�x\#��H��%򹇷a��/P��;��}-w�=���du��B��7���a��4�P�2�k����>��7�Q�̟d��|�������ZwA}w4����*�RKv���=X�
�F���+���������}ø�����B���..�'�q�}C���>_|G�����w۝#�����L6��ɚ-�z�r;#W5�5�s%c�E��Р��A����@��i�I���{��e��dv]j���F!�	�ijJ{�b)�uC�3�}����RO䁣���9v)%�[���ѭ���T1Ժds�I���UfW<5x��O`�,ir��8M����Nr�+S&��������w�ЁL[��2�ͨ���q���c���gG1�S��{mm���@�/���w����������4�]���Q+\W��eA/mK1��Tª�l��pS��N�w���	MA=����І�4�|O90̲�k�&�)P")F>G_(qA3t�EoewC��j%�(�UKsP=��/a���8��!0�#-��'�mWxK+gpܤD?Rv�劓
��%ډ�n��0M��,�)�$�cA�/�����}��T`=��i�w)���N����t���\�OL4�m:�O�22��'������"����l. ��{�y�N���ª�l�t6Ζĳxf�c:.��tﱥvJ=w� �6� ]�|nh��I.��2k4�+��0�������g��G�xJg{�� ㏹"��$��	�{�&���Ԛy���3�;mMCo���>�3y��f�xbδ�9](�Hg�E��	<�E��X͍i��"�f��������My��i�4�T
P�m��\��n�랗�u�yg�X��8A�z�`��>����	4;*Z�Ț[gPR�6��u;00؜S�4����7֦�v�E=`?G	ŉ>>�4s�
���=����Ls�m,���xv�DSS����ɹrDj�_m�rI�*�1���w��c\��0MJU���]�S(L��n#7z�C;ǆ�x��m5�kI�b#/��JJ�^���IxY_���5ө�������ò�v���<Vdp���6�����G���&E�@��M�%C����>Y���:���vCrcV��Ox�S�D�Ɩ����m�w�>ĦۊT�^��[ˣ�����S���;VǪ�\6Ȟ��{��s�����=�ȡ������n�t�ϟ0K�U�@tʧ�2��jy�6��|���XH-<5�sk)�9O�Do+MS�J�N��H^g����p�t-&��y�)����F�e*�m�� ��V�/�{W�ؕ�f{��l]�aiZz:���]Ç��,��A#�⡪��a�#�}��+�n��/���P(�^��W�g�)��1~.]�
&��)Ė"�3أhW��8��`�a�c����u1���v��?�݆�(�c� z�{�6�;��:�Ū�L�W�l~)�Ε���.��Ϻx�6���7���zd���1�U�:����Ncw����̹��=&��
P,
��$������D�A��J۪�h:�/vӾ?_��Ǘ1>���\ �����:�N�U�~��ǌB��1�)�՛eE��ܐ�z�r�v)�CP��L��=^��lſ���5�ʘwQqZ��pn�ṃ�F�GZsiM�(�j�07�0�M���2�:����(�Qqx`ą��()��?�^=y7�{~5u��\J�ޜe25v�����ۆ���<DaΑp�D����
�R��S��.�j�V�"uܣop�37UV�8�9L@#��Uķ��zF�F���*O���j����7T�<�w���t1��\$1�2����,[����D,1��!�i���?�����L�7S?Y{�}����7�~!��`S��vЄ?N��yD�n��N�*芜�7������Չ�4L[�^�)���NF ,`;�iWU�E6�~��QE� �>������1����l�bq¾t��)�ns�BE��n���8m�ͫ�h����I��L@]�[1��B��["8lm��Oa�i�P����{z�z[����R}�Z�3�2�sW�����B�5j�����ͅu���㗺uJdPL���Jh����.�>�vmt�ly��7�e��;��o'72_8�w�S$ף�M�xo%*�zjJ�H͖�]{G����vFqƾ%$(��o��p��p:�x�Uc�$d������W[��s�l�'�����	���Gaٲ�Pc���[��s�z��`��)^���V�W��:�ʿ?G��d�J����pŨ�a���z:�����w[��F`wg�q���Z)e!�h1����K�yE�=����e�͍g|���:6Ȩ�H+Z"F��% ��-��[�����Q��R�l��׆��W�v_۸��o�oB�T风��������:���sQ��Htd���2�t:H� X�}Y=j�:������(����9w�H;/����q�����{Ճ�X��T�\�Ir��Z��\�DZ��Z��-.��3)���z�����z�c?�[�c�5�U�X���#��"@+����V��Cl���.x�F��F4Q"L=T��[�2*|x����Rh��U�l�k���Lz[�9�i����A��T�r v�42WO:(��قz:bIn��l;�-=����k���8!t("����ku�O��	6��\z���:���e���jF废̑t�����N�\�]���w���n�2I�'xd��U9̿ F2\��s�]�-˼�"����k�׬$ajWf���J��㬏��d��Pa2sʲ���WV�qZ+�Cvatu���J���E����'y�v�s�	2rˢ�/zH��n�0�d��!)%�dY�ȪY�f�n��z�JY�f��]�����o�	Ck�,3�ګ��`+�4������G�8��g��x_���~>G�-�K��d��֣���t@=l��|�<�n��t�cμzl�A!��\g7a�������*U��d=z�CiϷ�I�0kư��H�p*k,��#X��&���5cԜ]���b�'�Wt�˂bZ�ķ�L]��No^-[4b��E�Y�N]�q}pū���"����>�n+_�w��'v��>�}9���C6�8�Z)c�'N��ؽ}
����?M�}u��$���z����W�ށ�X�ȧ������Q�;��
N70e~@��gU�pG�/�7f�̂�d���gN:��v
S�TR���VU���u印�3B2�T񗯏].�^�@���M��X�H��:#�O�����93z_���Ϛ�)�d��g/x�D��:��W.�t�4ȳF��.���ǹ����S]v�=��+��ҏ.��z����S����Y���`5�Ή�Fu�J%����WO�R��Wj�A*�d�_`�0�4v�r�V�o&d�A=���'I���M��)�wC��{��m���\��}�#޾$9��3����Q �s�<r�HE�O�c�v{y�,D+���C��i�����7��&���㲁G��P��L�p;�HV���񺶉PPD7���9+�*m�2\����-�1)Ӌ��1��a.g�λL�/f�]��+%m��'�*7�׻=C.�&��f��Lo:�����g���N�ޓ}�!�7�63�Q~�gn,,.��%������{k��)3X��6z�3�ua�{6�X
t��Ķu�4{�B�W���4���/�m���f�!h$�*bK��c'w%�%�l�jE�!�Tnn�9as�]ya��x�1T_bl�y��z�u�(t�Q毶@�Ǹ@���j�?vME�-��G4.�G���ˀuQ[�:�[�1\���yl�!\�eK�)�ҕ��g-�9��V�Ļv�k��6�ts��}n�K�T�nL҄d�ގ�Ǉ		���#lUŦe�m��Uh���>�A�H+��Y|�S u�w�N��n�V�L"�d��wN�n��F��9���z�/f�7F]�������gs\wUZװ߫0��f�؍�)$X�}�&$������y+���#O6Sͤ
v��tp�-G5n���aO��OvŕwA|P��w���:�w�5Ӝusz�FjA��#L�玀�5�:�k�)+Z�3dV&
�sGַi�v��LTU�e���Ə{���YB&%bj��#��D�W��αMr�'�>���k�I�E��*=�R���֪u���5�y{�}p����������Z�6fT��F��>QLڜG��)yt6�]М�`��n@�|{&�Ę��`�8��=2^�k6�WJFe�m�����������ŒA �I��Rb-�Q5T����Ō�1E��Dl�QAN���>O�������&���ED튪�(5Z5DwwS)V���T)"'�L������*����DZ��g���v�j���Ͻ���Z=��EDF�v:�'�|�~?ϟ�����F
�������4�1�(t����k�����ݜ������~|�|�ى)�������ӧݫK���Ql�׻�(�ݪ���Rb:\^��'��+l����`��SO�i׶��*
=i;۶t��>��E��=�i��RWAK�}QM{����DUm�q��}%un�]]�4Q����7����	h��}�U=umӬx�h�t���D^ي��DWm��~o�15l袢n���އAF;cg[X�8�=��Z��ۊ6���ݣ��m����tu�ό=�m�}Ʀ$�	�3��i4PH��j~,��m�6+z6۴U�G]�=]cAN������m����tc��ƣ��n�K��jz6��D�A����|0w���x��.��#z���ѩ��6�=cy=��o,o�ǭ�	�ge�}bH��/s�AF��'�{��7�����8*N�����g�9őe���c��mH�s7kE�] ��9��7^��7]�Ӝ_���0C��i��w�&�ӽ]��۽�*[��lcսʇ"A#�@��'�6�z�2�Q�ﮬ<�D�s�ᣵ�5(��;��yo;�O��y�G��<7�T�3�����9�uPg��H1P�L���_�v�"$u���ȓܚB��\�1��mewb�~���x�m�@�T=ܚ����>Z��:���y��\6��m[��3rHݍ7���4�Fש�-�#���|1d�+��C&uѐ�рV��\gc����=��X�W����SNj���E�rChӜ$]�4⭕�#�~�!H��E*�>�ٓ���=�L��(�ˬ�=tMZ���;\B�06ۄ���%��*g��7W
^�|����1�]�Ӡ��d��#�=�Ӂ�sNIk7j��ݹ�eL���AN'v�i�\��oA?0�{c����X�u �Yof��s�}���Î�4��l�X�|wo��}�e[�"�[���f����X����˴��*�Ūo��ߐ~s����jH�}G�x(l�����h�H��!f��=u�������+xe�\ɮQ$7�#V��I��ͭ��un2�ҥ�-���]�l�H|kwwny5����ha]���w+#��ݫj�yO�g|��r�y��{��w�wd��4���S�{����HٯV�|A�.r4�gv��� �ݧφ�i+h�j(Jpf��O��#��:ez���+N��|�y�Ӷ��Zo��\h,��r�Cr�������=�����[�;����)IM�ے�h�$I����$���7���ݒ�> �f:Rz�#v�nr��+�8V�c�vHԁV�l��%��]F�"A ���}��Ֆ�w�Z���9��{V���d3��!6�T#�(�MI��2z���ưt�W7�V��	�^�U�lS���X耂p�H��Om�6H`����O{�;� ��Y��M�nQ�&�y���)0j�m��8�3�P�A�4�w��Z}7����*��$hl���P��"��[(.��L��]+��n�;We�Yk�w<$��b�q���+5Ŏ�@w����x�̭���5�2� R]FM�J�ݵ�g0��a8xH� �ml�Yt�6Y�p,"�fm�ɱ8f�]�����Ρ�[^���Sr+�
@�#�ڠz�@����/��fu��7lme��Lhh>"O��=��d��Aw(\�R�t`��� V�]mx�׻�Hu~�ا�bT"�{q�Gb���G���*��Ҍ፮��e�ڻz&�~���?H՞�d �v!>SwN�<�It҆��3�v{����f���=ݫ�ǰ�lǀ6� ��k�߲S|=���xg�9T��^����4�Z}�Z���d��n���Ԃ��5�9kL�7W��韂~�*��վ5��:�֒��]˱���8mp�Ɔ��.fΦ�ݚي�c0�/]�fs�G*5�&��cy)W�f�%%P2��c�����F,���Q� �P(��==��V�`��������U�o5�\�0 䶭���+�7�9�+���]�����)*u�2ԓf��ۆ��;q]$�̣�B��yq���P��J�+(�J-�LP�؜Ú�i
�Ռ���P͛5�f�C8�S���/��#Pu�r�\��%�jb�hٳ5��Y*P�^c��gbg�^Wp�萐4���<݈��[#��{����fi:Y>���-{:������=A���0'gU��IX�תK]U.UMU���nޒ;c��᫏>du1��p���|Ζ£�4c��2��Ξ���������H�xID׿r�U�ndhoX1�6�Zٲ���_��6�9�#�$c��c�7m꼬 �#������ ���j�V)����n��v�w��a���;+�U*�3}Ϗ6�,��	�����eH�ݳ��c)G6Û�=���k ľ�&@݇X���䮞z�	�J|i�(8��}5��N5��>gMV��}M�;w�ޫz��0.D2A��F����b �\����"f�X�#�wR��r�RS��P{�;��GfH���!u(�݇
%�˵�����S[�mY0�ls���7I��ϛkEK��dz<��+�/E�B�U
�S�P_d:�zv����7�qt?�*����cT_�<{:J1���e>g|�b��S3�D�%m@\�b�eo�=�Ψ�.M�8����}�����b��oa�J^�prhP[��|������tĥ=ߜN�pۮ�:�Tv����<WIU�2�޺8��BL:���x}��m����8٣I
�\��@�3��v%T,�sr�����t��ͦ�2��U��2�X #Z��;�tw����L��ˀTw
�y��^������U�`�lͦ��=���iW���[���p��k@���0^Cn�A'����V���S�}�|�9���&��d���W�f�(&|ڮ��C�J��B�]��ۦ���@��#!?@���W�[)��똢.A2/ V�*�$O�s�1��4ۙ_��n��Y5U\��D�����:�F^.�����3���$���|U��>�G��,�M��R�9��G����Y����ں������:��6e��x�:LNn5&��zY��.��:	5������Z��7�
���A���<�~�w�z{��=�{+{��k���
p~�}G\�t�/n.̢��Z5��ܧ�N�5ځ�^Y&���!C���ЋЗ�'e�6V;�b��p��x�ݔv9t0g�K)T�,�33z`�썵5_gc�v^I��3��PJ��P������{yjni��7��?
ŉ����Wm���]�x;���ۭ�,R�Od���SNg�l�@��j�l`��zm%�_�YWi��	���s �q�hy"����nd�2���v-v�N����kB�����l��Ғ��T�zI������]�+���ݬz���-�Sw'���Q��_69-�H�h;�T��?O
���{�4�7��'�U�,��ks��h�.4L\yt�0�s{r4M��oM�+���#�./��ca�g��K�{����+��㇦S��xr�3/(�<�p��<mL���7�����F�:�`0�R�q���E̙�h
�Kk�e(�br�	Nf��O�7�æT�;���t�n-w�#GQ���>�/zV�+Ga��S�1�	� �n�?�G�ߏ%�?]����L>$��SfYRP�8�t��u �f��v�Ӊ/p]�^9��C��e��E���olj[�ܸ���ך�$���T��z�ܒ���b� U{�E��Mڌ]JZ�nHa[3wC�Y�y�2�YcFwZ�_�������2��˕E����j !�9:{������dٓ�O/��z_f��Ǧ{���F�����N'�ٶxw8��q��倛
��J�km����H�,5���+*����k��v
R6)�;W�wW7$�:��lI��t�!�/���Hn�����X��C��{Jz)���0B(¤&�4�C��z�̝檍Y�^���$���ѠQ�͕������x���	Ȝr-��Φ<�A���p��3z��0.Ae�I�8���ˉr5N"��b^q�1^v�\�#��tؕ�n��5c��C�)F�R�B��:4U�F=ݚ9���]��z���;�
���ñv�\}��.�۶��cͶWq�}�F��Uy���́�N��TpS4ڤns�Jʞ�{i����nL���F>������!�۠��r�p�����J����%���*ו H�c8o��ɣ�,��컵�M}����Vs
|���5r5nS�h��y���7T�l����+�=�d�}*��WaX5֏* 3�-��=Ŋ�΍�s1w<35�\K�q�X��f�m$-��_IKp�i���w�A�g�~�O�u�|�T�7z������u3�ﯺaa���JGN�W��rןu���Wr�|.���]B`�W<�#"�����X�N������ftЎTX����w��`X0��z9��j)�o2�x5^���zG(��
7���+A��Y�{���2�6*Q|-�xk��y6�v{�����s���g݇f�<\�mj���ews�_f�@�,�Tt��>�c��h�|	��u�$����@b�[���	���m�q�4n��q�:$���d3�b0_/z���V�R�V2
��ݑ��~�]��*��Y_Gb���y�k�KE�n6i~�̔��c�ҥ �iT�]P��X�u�:AW�|WxO�VR��|94��wYb͍�����3^x1�`�z�ʙ��!r@evdjO��c+��L���(�wä@��iƫEnn(�V;�r�8���9V��|ۜu���x
g7ʊ�L�kآ�H������R��2�,j����I��s����L�;2vMҦ�ˢ*pN�#���k��rL�� Y���\����.�r�/�S�A����a�w���s7"d3���V�E��:�ѵ�Erzd�O�_,~��U��4��c���rY�d�݄Xw`�kl���Ԋ����o'��^).x��S�n��$]y$-�+�4j���s6�kx6����"2�5�;ΒW������+EK��ڼz�mWC4T7�q��(��?��*�C]%V�\lk�8���sK$k(��sMI��<a�tqa��(:�t;�Я�#��W���[��*�\�һ��X�l�+ T�k|=�;����B�#��-�z��NY�]��I�D�MwS<,���]<;���N#S�`�l�o����`WH����1_|�}���r�U�[�_|Mfa�ӻC�u+�жF��^��s:L�����G�_����nG�|�J�ԍ23��/y�4�F������5���$}�7s�m�fa�9|o��e.�S�=�������yHǦ9�L��ڴkȊY�*b;�f�Ye[�
�eϻp��`Q�|Q�x�[)���Mۢ���ǀ�JZ��At��_'�ǧo��eo "t8�z�L�2��U��#�6�vGteލ�ᣑ�&�P!)�wǭ\k��H���1 v	��n[���6j���Xd��t�^��k0�2��n���C�p�ȑ<y�E�LX���s|�d�;�na$��6��P�,,��O�sٛ�/	=gc�֠��f)�O9̶7�Fn�;94�����;����w��ܚ��8��_�����'O�rp(+�!.ƛ�R�9������s����݅l���:U��ə+;;9{=�J��o$���S�vj�i̊� o7&��}U�p{&�œ;�[��~"<�p`/���Y�
x�4):*[*�Yu�S��^�ӏs�ą�H���u���W��\������V�swu��w4�[5�p[���"2]�r]��{-�Yx�l�\��e&j���{��«3��/���t���ɶ
pAǛ��չ��h�} p}�w"%�=m��a�͝3���nGe���k�J�ԙ6�^�#��/�IӊQ����3������д�瓌&�5Od��}<�q�&��,4
���˳٧;�)��,R�g��hm��R�v����&b�i��kn,]m�Rcj�£)Ĳ�����*iK�g��Viś+l!���
Snܠ�^���S��كN���`������l�<�N�qێ˝��|��E��W�d���P�/�L�3� U�dgol��>��G�]�q}������ ����J��GC9ǧUe���6g>ᗑ �ܾbvW��4�<<��`��a�*ͬ�o`w�� r��~��S1{��s��F�L���6R�qFfnө�\2���1=8&����\�<fV�3���LQ�#�h�Z���"&yM'�m�	�m֕����oL��E�Nվ߈1h�D������B5Ɓ]ٙ��07?��fJ�S�8�]�����vX:+��tp������ڬX�U4c=�� ��%s�_e�2>{/vu�Gi'm�U�S6��3���޼�%�;��羧$�^^% ����ה�sۓ��I�;]+�5r⮶��)%j@T8T�X'hV�)�:�m�V�Y��X�|oxX�}�<N+5}��d�O�����N��c��Ո�g�4sg;����A�ƞ)B��"]�J]<��o�2��_{�����]�익�s���|hƜ�M��y� Ǒ�n̽X~k'Nd%�0�����Hd��/^5�������ە�7�f���={�N��-�v���1_<8'���yY�{�W͛	��x�����x�[��Y�*�ձ�D"�x]d��5�<k7���K[ �X��`�0���۶�l��O���I*��l�ϝ�[h6�8��<�r�V�
8+�{|EMD�TB{3���-��2a�6��m�l�wj�M�
'S+��=���7u�-B��m�G�+S^�����v��d��C'{7�(��N��V�h`q��W��C��$��)��b=9+A�Q�Hr����A����b,6�2�d��켉�7�%l��.}ԛއH�`᝗ILRî+r��!]7��3;V���*U�Ƹ&V(M�P������B�b�;���qm��yen�ۨyrD�P���V�'�2QX�KvҤ��s�V^iLl�\����<$X����c��m�wFЈtu��'�GL�M�=�Z<�~�QM�x�X�b�+��ξ���jE�%M��3h�J�W���l��f�C�a��Z�˴����q����"ն�Ï�opd/<�ʼ��bYmV�r��޼ؙTٜsr`�^��ͣO��)��A�-i]oMLVoK�VH �)���>�Β�ȅ�z�Cкr�/	��/o]�H�Fe#��t;b7��m�ɫ��i�6�[̚Cq ���(�R־�RG�ۮ_Y����b�!&#��ـ�`�u
@����:e�P( Q6A%��m�.1�}����C6A	Z,wm�D�p�8�uv�f�=j����)Ս�Z�OGF��]4�>��~>>7��?7��q�;�p[�mj�`����i�n��N�n�q\mT[nݱ���矏������h+X�(+��K�v�V�v�h7�/w��l�*�z:���s9����?7�v�j����=n�0�?���)B�K�m��6�P��]���1��{RhӠ�Bx����<矏��������ӣml|�i{1���ǷGn�Q�������:��/Ti:�5��kt֝����F�5�'F�ƍ&��b�*(��+T�I6��C,��C,��m6]���8���l4U�{WK����E�=/��$QU�Ӣ����I�����V���U�ӏov|mF�ZJ�vM�j*b�-��{%c�*
Sыwp��ulod�E���ǣ]{=�qm�������4����=��X5G��J����lsv5tn���t�kѫ�K!`?� ��0�RHB�ߩ]7����O{o����eC�2��7�u��ȷ��m���F��ݠ���U�#f�u�)m�C����d.V�ZfI����[:����W{������Fl�l��3���ܪ��S���������j[T9"�K��&�{���{����y�nߝ_����ŗ/�Ä=�S$�G7u#���L�	N��)>���"޺n�U��y9�ƾ$�=!�y��:^�LV�S��3�F(�^��s����v�[�+΁0�g ,�/�/��u=R7����C}��Վ�i�f�p��HY��A�k��сxVv1.��m�}fڰC	g���ɫ������I�ݥ����t�~�]~~IPהm�{]���_kZ;d��3kܺ��4���Z���Y�tB	�`ڹ����@'{����|�{��/��\��	h4�]�siM�-���k�~ӻP����Glэ
PB�]�z��u �+ķ�T���v�x���T$Ԩ��~����e�ȷ&Πnʯm��(�Ƈ���%��Q��wp�|j�û����,d�5���9Å%�4����V��f�P8|T%���{��y֣����2os"Յ}�^��\�Vfn����ႚ�K��|�9ظ�I�7&���^a�|�R�p"�S��p�ڧ�dk�U{��R��­�����P$���{����z���OH���A�9���ȩ�"|����Νt�l<��� 7]g�͝��8ٷ�DT��T�p:�֛�B*pOM�f�;ɨ٫�Ɠ�u;<�>�vj�y� �]@����A�!lAC^�SN4dU���XQ��#o�+RQc�.W��ֶO�S���am��o]�HU���h�!רk�B��S�ئ�k�ZJh�+��a�����g��z��{�EL�Dm���:�1�������V��^�MIW�h�M<ϫ��u��D������F(o@p��p��7"�wy���3�xG$u��8�`�_roK]���6�n�w̄x��b4H['��l�n�W�{��_O�*��1�d�Pc��s`S�x@_5��HXՎ��'K�W�ڼ9�p~�W��DR>.j�B�?b�w�}�垹�s	�Ǳ��[��A^m����w�) � �J�o9�r9W�X3);�#n�[N��y�ƸS�K���)XW���\2?\/����1n<A\����73��kr���h��`�D��~��w���%op�<y�g�Lq۽A��_Ck�lD�Us�K6��7��/;/5^Y��%f ��[j�E���ȱ���.�V�T�<: H�{�ꙫ����X���>���k]�kZ��m���(���V����a?�U=^6y���䲇a�7R��Vcz�t�e��]�XlԷ3{X��%�AV�X���B�F�J扼�9g��r���u��=�d2hA�T�tK�Sy�=J���QZ�]�t�t��%�#,=��tQ,�p))s�*��-�u����~��|C����;u]�v�HC���n3�+9�;�t��7IK������C��)�|�u9_c^���}6ڕ]��J�4��z���ͨ�A�������]�u�n	�}��p¸.������3�ؕW��y�Jr�U߼�r�4���;a�A�te�%I%S"q�
P�BkD>}��%w̺�5ж{�5o��헻�$;ceϡ�R�eW��ػ'�~�7�O=�n��G#�<W���Fn}�2lZ�H�#I�XS��:�ӊ��a�c��Z��>�>���t]�{��;�,mW��*�2M���ey��ln���޵h�����3BV�{��qCq��� 0��]#'�b�b�h�V���X4u�8�j��>�9 qӴ8�R�+�-��:��o�h�7��Opb���y:f��a��C��3��D.���s�>�6ha� C���{���b���)Kh� �P� �
�A����#Is�#�OC��z����{Mn�GsV�|U����������;��yo��9/�9m�1	�3i�sw?�Y��N&���,�zJ}W]~�ؼ$G!}�'2�p�{[�$U�Mmh;ܚoiOE<���@ �]����kʤ��[]�L�	���t��ve.Ƒyj}sNd�t)�b@�N���r!�MvS�M��*�\����Am��rV'�
{�X��3�f��w�^�X
��`�M7\|ol�;%Tx��������W3r�l/ GP;v�%߶�&��z�o��.)�e�Ҳq�Z�T�!��
�j���z,PL7����7=���|ζ��%����I�qi��,9��Fף1��5s���8``�4u��z��[[��,����m16��ԅ��~���g�ӈM���:
F�]ĤD"����.(ɨF-�#{FE^�~ꛦr6��+�xc���eq;Ғ��yl�
��:M��ɷ�����)7��s#Y�
dV������͎K[��l��Fp�C��6�p��{�\�ݛ�;o��o�PAۂɍ[��rj$Jc��>��j]ͯ�Ӗ��@ޣ��O"�Ҍ���a]�2�G&i�~xu�9���s������M�GN�{�/*��W��{�<i�cJ�k!Q�:�q\�zي�����!6��䶂D�Дe��y)�L@Rt[Ç�j/�m����O�>#_�;��
�����V��Y��9\c�����U�&��E5,�-�c��t����� �>ّ�H�/�/���K�����<�����ltZ�Z��w`F���K�[W��Ə���~N܁�taJ����%���OY����ߙ���@��P�����iQ1�r��w{JSp�nɓ�߄���YkV�w�C����y�2�#Սd�d�����g���&�X����K?��,�eq#^��(�.8��5����w��6嗢��yB��"|H04��ôY��s������&ܞ���M6�OMWME���"$�]@�B|�s���:_M�}�q<$��3+s���<4��ܩ�*�"�rBz�3�ѠQ�Zé�Y'=m�f)���U���i�;��X�=�ȃd�\fz���
S�v�[�S�qH�~�?�k�0��
E��z��+*+�.�>���k��G%�^��B�:�"t+�,��5DF��e܍V歮p���EO��b蚶"dgWP��|�������Y�j1��c���Ti"����]:�nxĂ2�#��ܻ�.�o;g��٪�]���O���q�J�θּ����ioa��xn�O7ٞދ�B�2�V���O��q�6�ǫQQC�&�+O���;%O�����;�WXn�#�����0��T��϶zz��rןu�������-7��1wP�.�4��������c�rk٥�������"��l�u��:�2h�f����/Yy�ꑥDzچ5�.k�#� �k4G��r�Z��d��^�`N�7�Ӂ�A����ʲ\�E=��o���+��={�����'~��]�z���壟 7q���^�4X��=�*�I͕�!}Il>��=O�q?�ezk3̆l{��y�Fz{$nE��ͯ���2=�s��vwrܪ����"Š(;�&��<��ˑ�+|��{8�ݸ���C�N'��Z��:A�=!���q�������
���NMfs!Zq��.�٭�Y�#Lp�᧏>���1�����O-m�ܷ�.::��B��l�M�h��7�Di:(���x��z����Bt�6{X�׽�|>�c�v�L��^\,$u�:�Eag�҃/��{���z��||�W)m P�ꧨL���dT��c
wє/��=�V�������r�I�Rh=�'�D��,���&I�d�ꭝ�Rw7����x���I.F�{y�$كpuU���O4ԁ��]B���TBȸhm�P�6�E]txx���Q�˙]d��!4���!��.�.�M��Ǫu�<��]�֞�ز�+�u���	1#���(�����#ON�9�c�dr�۴���Y�m.}�������LƊc���@Y��K�訋I�]^`t�[5�s釱r
����Fp��^�I/	� �5��n[����Y]�(�����OV�谐�:=���$lt{6
6=ΒV��\e����#wg���͞�c:3�Ү|d:=0F�ٕ]��
�*��㬍�g)�U<��M�nކ�fv@a�K��q�.ǆ�z{GjUV��>�]KI�}ζj�l��w=I8J���T0�l��\#ϫz�AS�`����2�[���l�� <�k�c�$Rݕ}��=����:=�DQ�ٮ��\7{����s��r��1_T��4��{�\���F�St�a��.!l��[;��Y:ˉ��sY�Qԍ]9K��z6Gi�h1�m����y8��	�'�%���¾���^6@�<k�d�GVq��l4l���z�ӻd�~�7ʟ�?�<8a��j�m���tyk;� ��,��jU#Qi}�Fi���{<ۛ_�8e��zGw9��'��.��6;{�,i�-��X����۲Q�n��)?��d������?g<(����Mf���B�Z�*�IaG�_j;�6\u|��9�YT�&.���]���sL���;h��ܚ��a~-�d�[W��_[�X�o������7�~ �M(�ں���N�D�A\9�E�V~�ݝ��d�^B�4�{Jz)�a�P���r@�jBC3�Xq[T��:ET{/(s��GQ��]�K��ז���5 �ss�6͚�h�5��7uog.�dg �
FM�*V��f�ȩ�0QL��-��[��ꋜ�C��Sr���]�s��i��ĥP�|��iE��;�޲u��S��7�O_�?�y�J=��F�Ғ�^]�f��G�O;�gQ��?_Ht�X6譯N{��E���]��w�:����ٗ=�;#ufN�������m��m�0�/p����UM���3�H���i��b�[l��6s��<z���oU���3��~&,
�;y���o�C�3c_�}��/�s[����ܙ8����������_ú���=�B�����(��O2y��{�^����H?iSb��{]��yl�O�d"bW��ul;�&����
�rD�[�C\��wI!\{R��3:,�CQ��	��v�G��^wv���5�����`^˾+X�bBY۩z����������,���N,ޘv.!)Q�yx0��j�ٝ]����jD���ܮ75�z��	�*J�翂ߴ�n#�����#p�b�[��s�F��:� �����^w:��f���n�L�9ݼB0�g ,��>��|�C�,M{9�i4ϥ�N��j���;wC)�~�F���K6�GO^r�l�3݀�m�*$iDH$ӭ�$�ا��gp�t����p��wC_�>G*�Qv��bU��Ǌ�%�Ք�b��9,SKCe�ٝ�J���F`ל,��XjeI��!rBz�3�Ѣ���ҋ֨��)�����n#��+�`�w/�N��q:��z8���t�48$�m��qx^�p�v�KGoE+�s��h7�������B�V�oٰ�X8kr]Oz�Rǳc��o��;�\�a˽T�=V� �NEO�>���̗QW��%��{i��v���;Yz�����qv�T��
�ZfC��J�M�B�iGF�Y�p"I�6���N�p��;8�{-SC��$���W�s��,�##��A��yHA��zy`ܭ�Jc�4;�t�C2B	�[����r],^)d�o"sL���IK,^�`,cia��٫�a��^Ʌ�f�u��S�������g�ï7={�Ҫ�p��TϏ�c���(";�o�ICk8%� <�<Wt������S�|%�bp�I7Ǐ�����}���c1�y���܀��h���;���q�eԽ��W At�4k�p���i�b�|��/��w�Mr%zT�p�,L�z�7������Ƙ�^�I��[��yk$�{�:W�c�8�zm�6f?r����o��.]��VP���C&�u��~��C����凷��G3 �g�.Nw1�j��r�\�F��_��W�)�]��}�EV+����qd�r��˭+��
�芹%�:�'�\67b�l[p]c6���m�D"�N��dS�۠���;�3o�<[�F����js��ʳ�	;���-�=�U���k^�x����)���}R�
�}&ׄ����-呵��)��$b��	��j��G���vZ�Ø�s���w��@�}��;�N����u��wa�̚�$��ǣ�爫"�R;��}�����)�1p����/�ਆ�2�������
���9�A���jv�<�($�$�k�?׍�N�� �	e�ľ/ί7hZ�..V�)��%jӫ�*e�΄ Ȩhw��5D��d4����:C�YL��W��(*�NT�-���L{�M!j��=���YK�8��]\�|��sn�R�Yrcmt)�>��Z&]Kؤ�ä����<��?a�a6�
�׆n8w3$e+����u�ֺ�]i=���R;��Q�"��g��&�y�"�8�d�ɗ��U��Ş����=�q6:�T뼁�Fc�����n�u;�f��d}�M�.��I�U�3���3�`æ���ȶj,��y��f������2g����#>}/�=��'��m���^���v�n?<���Ᏺ�a��!�ҋ�n�]��.�W+ER*w���'v�w�)K�'�$��y��"*�����e[�'/m���w��7�G�h�l�ֺ�t�^�Ƕ��#$j�6�9�ԇ�=�XM ����Qki׹���/�gwЊ�b��r��Y�<SNq���J���׊�\ȅt��l��q���5G�t��\ag�pV ��k�F�9���n�<W���Q�f$�jk���38-�zT��b��9oa���n�ŝo��P�G�j �eί��(
��������+�k=��ﳈ��-�U�ޖbg,M9��q�f��)��x��~��v(�v�>Ol�v4�c�ܝ��6�����.ɣ��3ϟ�������i.۳κ:�����jj�8��EV�Ѡۣ���#��~?���|���M��M1[:ݺ���4R�tн=�q��$N$�~?���%|��7�`��[�N��-i��F�Wl7YѶ�"�k�9��~?��f+mQ��b��`(b��Bhm�Ӡ�{X5�n,Vރ��Otupi��Dh+��0�ѭ����WcT���m���wX��ѣ@v���]=����S�F�gA��F���իUWa���������h:��f.��8�U֣l�-��t�����{�K�X�t��P=t\�GcU���{�Q�h�TV�ƈ+EkGG���c�1�+���B���?�-��?���5����[BX%�Ր�F���6���hG�5#�w�ɬ�gT4���ة8^M�׶�����+U6���u��_�)K��ٿs�<~��$U6��ө��l�k,�ΐ��2�"�F�'U�N1�$6��'Y)��/zRWθ�מ��uux����.0:�n�Z�� �]q\8$�7&�p��c�o�J��.V�c���ؿ|lQN[������x����u���0���ϣ��!v����2r��IO��;\N
=��X���;��s�^5�}�^u�Dl�~ Ibjs��m��aؒ��s/���H���|W����}Җ�Cz �C��}�i��������k��^�A�՘�m[�Ǻ�AӐ2�����üB=ꃲq�F[&k��3x�*�6�Kpz^��"���;*�7d�1��g�@���G���~2��ԙ�<��h�4pg� d���y�<,ٟi��4�xE�cy6]�ޜ��39M�:�Ly�t�������ȍ'��� ��h�l�bσ���Q�s����U�G�ⶴ�3t����<�δlJ�w�����u��G�������U{}]�"5�HY�̋ ��ԝz�hÂ�v�y2��I�6i���p����8T<-�u����#eJ	����k��.���5�Ez�w|١L�-��&j���a#���`�,��.�gsu�#7rA������Ch�f�$�Q�3g�S���Y�ʶڶ��x;��f��p;p�X2�4
�i��3T�dag�
�9�~�LK^�4E,��>\Ť���Y��&��s'��&��=�f�ttNwWt�����qD��vu�D��Q+�x�x=ڑ�n��.��,��s�7�3{��r����E�pQ�� V��=�
Q�I,n���͔����vs��r�����_�Tc�����6̪�/��$��+���V�zE��J��Y�9V_6�vz|���d��!wY��Ĩw<����Z��Wt=v�����Ǹ�:�ޗ��k� >��@32�{.��6V���d:�9ZO%{�*V�{,/Ѹ���do��bl��Y�)'���6�MYOH�n�����SKܓسh"���_!9�R���(!�'^�P��N�x^ҋ�,�@t
��ě+O2�K�Y5�}9�"m���q�6E�/v�VNnB0�f+�ɡ9b�w�|�K��m�k���O&�1k'FX� `˾�
k�7+D�n8rV��W'N��8�R�+�l��u7F�)�鶫�<2+3����V�݊��@�F�.��.��}�v����ڜqpŋ����d+`55��o}^�
�ej�Ì�>$u��y�1b�ֽE�M;:[7���r�5�F�/ޏ?p���\Uc����k�t�h"��A�w��<��:*F��H�� b`=$�7=ՃzW^Vd���8L�ˤp��}�"|{�O�is������	c���+ ���-S7op:��fb�*@�)m�:�^Y�)v4���T2�����].2cPW��惱] �$ǝF���_��B�RT�)G^x���?jb�*��Ώ;�z	2p�V�c��h�[a�����$4���R�;��mL.�wu4��M���n�4� +����{�����gy�$���4��7semZoF�Q�D������"��K�2��J窈>t��7!���ɏ�nn~9���-E��������y�SO�Y��kT��݋��]{n-�5�����}ۈ)C�ˏwOr������O�a���9^ﺴ�@{�dd�̛9�9v��Zw�Ha�O���Z���Ȯ�#�u��̧��)�v�eX�N�9o��q�Z+<�Y�<}�D6�PC[��f��D��[�6����I��ol�ב�G��L���O��X_�;�D�<���S��Hv�����x��FI]C�mqE�
X^}�vM�2���o��k��s�s��xT��Ô8Zd���tʟ?u���[IS���ې����.o���k}�5���2�Q���;�J�r�[�ٲ1��	ض�Ǭ'�{�& w�o+��6|z�t���g���ǃ���2ܒ�zU�Z�]i��v���T�6������Ϯ·t� +)<ʺ52*$K����Ԫ��e��Q�7�H�$i֏EG������(H�p7z-;�KÏoc�P��]QڃyF���tDO�pz�X��^e)ا ih���mvi�ڦ{�=zoaO'�Ye}�%�>��5L�Q��M�e��%U��q�5L��ݳn�ɽ��L]��Y /,����7������۸�BV16N�v&B��Vr�rLM�ӣ�d���!��C|���69~��.�*{���^MoyI�ފ��C�DP��Uf���ۏX�b|M�^(�/Hv���}9]���[��};,�Ǭ��s0����\B�U~qT�3�-rD��_G�ξG�g�vө����bڳ�Ds�^޵�e_pW��7���J �)�F���Վ�U�����ER�+��-�k���f�����v��.x&�F�*�Ϸt�t�<.�*�&Ұ|/�A�:��u��؁��i�Jw����{�:��'���� 6c�l���J9�{�k�x@)�FD�6�Ҫ-<
�TW\�'�����,�p���N^]��ξ���Da��F��DG�׶�z�b����%4y�VZ�*K����.�S�W�Lr!m���W�X.dm�5p�4X�����ʜ�[֢�{�{���H��ʤd�0q�o3`z��^����-���,�]cq�������J��@h4�vB��Vaƺ�Z#��ߐ�������sS0�e%uf���Е}��Roj/��fШh��3�]v��a�t�=�����o���E�.Gf�U����i|�蘫��+�;�6d�{���g�{���x䌐@����1�]��r9��a��h'�šr��Q�c���E�=�j�϶���}2�x�W�0��eSn�y��0�ӵ�Q���f�i�;���x��D�B�3f�9e�enf�Aֽ��0�((�-�b#��ڴl6k�7�DH�xH+|C�nyvM�[�O]Al�4�;z�J��-ԍ�
�a�ш�������t;Y�(�x;���݇Bn�I��w�@����G�u3�ŉ�Mw�8z(i�aq��'��������A6��]� �SÚ�p���2"Le;mhg`�,D<���,�������tW$d2j���tKצ�)���ƺE�p��LfMhd����i���r��^�RR�v�Κ��x�1!D����7��z�H�H��!m�}67�t����o��~��oX�8b� AB)%�Z�sSZ"ݨ�w�kt�n�t,�4�<t�F$�0P3�N�mn�f�r
U�R�٢f�c��l�5rW�����a;B�E!�L_h̡!{���t����pi�h����bXus���R$�_��SS*=�l�F@�v��+u�
i��A��S*�o[Wf�d�DkZZ���c�F���V2�Et��^�6H��2�#k��q�}VD:20�l���z*���t�@�3��p���)�u8��귍Okt���y�I�����w�@a����ռ��́[1���w��F/\��ʡ�yR��0�t{��F��x��k��~�R�]���Z9����G�v�T���V��er�`u5{�O[M'��v�5���)���ă��lz�+���GR4MF�L�sUi�\\�4ԏ���ץ�U��r��&��>W\�^6G�j�\d�C(�Su�0d�����{c�A�V�}��:,�xTj2��n�ji��F���f�R�m!�5�۝����5p^�� ƨ�_>o�~aV�G�:�]f<ޚ��8d�OM@�[���;h�d����`�v���(P���o��5��̧��o��ePgM�nV�M2�ˌ�o�CFؤ7�aX�G+)sq	kNd۱�����t�I��p)�z
�j`�r��3��� �8���Xgeͅ8�G=�X���<Om�k[�p_:���U㫕����y�\��ud9�y^�.R���)WfR�i��74�0�*�k�w	���{��sY�C���<���J�F?��U�RT�J�=�v���s����#&�H�g#n;&������΂��K�9Θn���xK��B�ƛ*�[�i�@�$FH�[co��c���D�F^Kqd;#v�Ǎ4���<Ux���e����
��8)�۞��F�-�::Z1��\���J){�L�ݟv�Hb�aO���{�ڬ��ӌ�sWu=ӈV�g�aa���>�2N'�+_zN��(���8Y�C�[��=�Y����6hE0�n��)��swi���/<���K���=�|��E����}�,�g8�P-�ٝ]����%��{�tA�WX��Pw��^����*,�Tr�2a�##dnnq�.�Z)�O��=unw�|��g��o����:��fƥ�6�-C��\�K)t�k~u�},��yLPBb^��US
.������[8�ݾ2[�ȥo���UF�n��Ė�������[�:R�k��.�7�|.�=y�IPތ��v(M,�9�5���ĺ���
;��"�䛔1����n���������:m��� �`8fFHYCǁ/yuc��B	����>����y��z7�OgPg��!�X�D
-��'�o����}rOP�m�}j4sF�i��F}�O�2�V�O�6�H��뒯G^Q���]3��V��K��������OT��r��o���bI����d+F7�G�#_���ȹ\����h���|�j�����0���_WH�m���(+�XF�2�BĪ.2w�YҚE<��73]����������ysNW�Xo8U�u�x.յCD����D�[3��I.F��(�JUB�����U�p@��R��y�Z��1��n�y�YR̄nwH�H�<C��IT�pK�Uʓt�=�vM4������Qգ�'��@�d�s�����h�	����W�ȹ-�P�6��2�B�f�}[,PZ�PorZR�K�5I��}Rp��M�#��r�wZ�����Yo�;ҟ:�_M�&��MU�;�2��8��WZh�*�0\lǤ�x�J�c��Mu�]�z�
��E��pa$n����4s:orV��Y����%�Y��:s~���á�>�pdm��ZJ�ir��V�&N�l��czq���m6eH[�0�ל��u���݊7�~a������I���}M�V &�^\���,�}�ֆm�
}�!q�;��Oq��W^���C��:_��R1G
>ޥJ�T�����x��������`@��>�}^˃�\>�ߤ�����; 䌑�wӾ�K܁�;�/v��l�d:�Td-��,����sԟ�S�'h�Pc��6��j�b�ivp��d8SP��;P�Do7E�3��#ۣ�t���p��%��)������&�
l�2�
#�:T�V���"4�
�e[��`��ݬ�k1�7bY���9m�=9��B��F"noח���*�D���Tb��.�I�DTi�"��@�狜����_�>C�gO� >_l�'� ������T�����"������8���������0L)2�00(���
@��2��!4��!
@�"0�����>S�i�@��9��A��*���U�ha PhbdUa��  a@	
aE3('GD� M2 42(���C�" L�0��4�2"�4� M0C�L(v���Ą̀!3* HA0��2H@ 2 ��" @� �ʪ�� �4��  C� 0� t��UV ��U��U���  ` UX UV  �����U�T���Q��"��!������>n����hEfT B��E�� ���|�/��`c�������_�Y��������`�)����� ����}7��m_aPU�����?_��� �
��)*
��H����+������_�q�}Ο�/���~��?�?؟����
���O��������~��~0��}��HD��?��Y�`$W'�[�?����C��/�w�	UE��i�ہU����(��A��%IU �Va@	X�U�@ � ���Ud� %d F  �eU`XUXV �` @ ��  %Ue� $  HUX`_đ�*�0 J�Ҫ��B�� � R ����bܻ�}�_����E�6� @ (7�O���}������~������ �W ���7����������)�>A����O�7}�+�G��H�{���y�����1��x����E�����P����� ���
���hTU��ATW�D?���~�������E~���������J�����?�''�~�x �pZ��C��C��ό���gӯ��'���'��"���?��/|A�����$�I����I�a�=���=>��W�t�s�����4{�}@�HP��"�?����?��w��TV��?����E����?������i��C�_����`���>�=�u�B�N��@=J���/����Ee��C}�����@@^� U$T�~g��'��P�8����:���X�O���?A�� �	?`����p��ڏ���2���@���e5��Sb �M� ?�s2}p$������>�B&ڥ"l�}i�R��J�*����
��U*T��m�B���T�k	im)�6`��Z�
�DJ��$�Z;9�cZY�[S1[mR֕cl���J�V͚��YE�T[l�3[Z��I��m��c��jR�Ej�I6�f�Z6ֶڴ�5�m�mK66���]���6���šZ�fʕ��֛m6h�jMh�B�[R�(����PU��Z�mH�*�VY���R�c�Km�RͲm��&M��T��vb@�-F�  t����oom�n\:���m�x�t�ׯ{��ͼ.[�����w���4�]{n��W k�u�ç{�Yoa���^���li�^���q�{7(�g{MףN�W�ib��Ye4�j���k6־   .�}�M�ж6�v$>���}U���lm��l]��w�l}��4dm��m�>|xt(P�M]����ݛ�{������{[�v������p[��u{�����U�h*��vݶ�z�ǫ��{�������,Ն��B�n���  W���_v��Gu��yv�]�o^���޽謽w���^��ַ6��zy���ݚ=޲�����f��Ӡ�wsS ֵ�Fj�v��Ӻ7���^�{�S���[V�$Q��m��   �4{�ܬ�wo�{Ӎ�6��e4�wv�]��u��lö������սt�ޞX]�OWd�c�{t��/77-̝HP��{���K���
�B�r��+md:�F����a�m�   ���[5�
�;���J�cJ
6���;6+N�܎�[a�8u�ZԮӛm��1��b�ٍ�����U��l��st�k��Kki�4�W�   v��mƛ�}�]U�g��.�8�Y�k�2v ݹ�+�=����u�tn��+���
%�[t�T9�q�-��Β1�Y)m�|   =��Xz�`mZ��Aܕ�3U5�M�Wl��W*5ѳ��אm�  �z��  θ�(
�����ڭ���5�m&�[�   ]^  ��z� z n+�z� ��C t ��  �ta� ��8���`: Q�ז�Q��8w�  =;����-�efS5mgn��͕i|   w/� ���z �@ p�nz  �h��^��ǋ�� �[��)�����=��l�  �����z�e���U*�4))�   ���]@{�w� :�ۀ�����] t� �үp {�p��˃�����  ��o@ � E? 2��@ h �{M�%R4#MhE=�&���   �~�R�4d � � 	J�  �J�ªF� ��O�����?��V����ͼ��fV^�|{�'N�#n^�4J�-��>YB�����0m��������f�`��ٍ������m�o�m�o�6�6ɍ�����G�?LG�L�P���B�&�؊ػ���Y�vЩ.����3E�k
��:A����
�j��T�m�he�	M�++�8	x7(��;4�+�ZZ(S־hPG��U�h���b��W{:���g���T+�"���آ(�(!��6�ݣz���yɗH!!Qi�5���f��KE��M��I�M<e�Z�[���ж�B4naR�6��f��d�cr��ĭ:Zx-nad<�/XqTNk4cj�n���v�I']t���э-[gq�S��d��U�X�a�ڛ-X�
�<�dգhn��SY��"��"��D�z��P��&+��#'r���nPxrQ���H�tºJR�8.=u���h<��)��5�@)���)f�\�͚R�10\O^�$�2���P��5���%	m�M�ɒ��\�@A`R�)���$���N�Б�q���H��T�V�Yref��
/sr�^-.�<H��^�J�u�:w26aHR�$�7�Rh�W�w+Z�Z�!W�Y9n2T�X�$�4�6����m��" �eaŲ"­{F�®&�r��Q��w�3J�N�PA3�t�YV��f�D��n�H��5*㲍@ ��v9ETj��J�����ܨ �w-f��[�D#��ĕe���Sf�t��%e���N^M� m�d�:&��AJm��h� �K4�d�rf��ͱ3�H �&Kz��Ւb[@@j�D��J�Qi^ыr��0�@�����B)�(-���z�=�(����lK��b�����v�	c�pT׭�̑*�� ���ؔ�a�N\�%@ҵX�@Qɡ]j���z�Cn�+v<i j�5����p�N�	,�)��U-��f�.��[[���v�(��QȬ������:�pp�|��ф��ХA�j��v�z;tkϬ�k2�m�!�Bw{���CV���&��m���q�j���m�
!Y���ئ37@���c)��4�L�Tb�v��驖6�R���8tb����cd���f�����1A�#E(�aP�Gsec(u��wg^ZY�ĪkV8��P�)�r�T5�4*&L+YjJ.��c)�5�����X�F�n^��0"v�õW⎙iM泵��j�j���n���V�[�Q�]��S[���ݧwOZAi%�J�vg��͑�zUwNE���%srW���YF�¼-��ءN�v�ɺ+J�H3�Z2�B&0�]q1���Vp�.��+g��Zta���ɺU���c�S/�su8@�0�	"�/�&�6��s#4��O?YZ)�֖Lz^�\(��N]��e��Q
��3M��&���4d����U�]L�n�8�
9EX�  6Ctpv�i�0�̻�T*��2&`�Y!��;�A���S�K�Jkc�B��V�8h����pnЬ	��t%��v�T�L'j�EX�7��ͬ7C)cSq�7(5�E'Lz�����U��R���3��J�8��[�`6�p�v�d��kw���f􇹭�gw)e^DT����P`v6�l-6o�!��YB�ø��IJ�H�Riʱ��(Ŷ� )i\x�����5��3vT���m���J���JR��L���Vn�H����x��v�8�Ğ
��Y3�85�l���d��DmD邊;���TyCC�0�Z�B�P6�4���'p��b�$t�X��9[�3�P����`���ӬX��3MB�^�+V����	�ݔMk�-���wln��E�.�^����W�2m��%/ ��j4�w�,�����*�R���`��R�I`�P�R�����"�3x�y�o[�#6��F ���m�Ì�{��m�{v�,a�,��c��h 1n��،h������W�P6�[��o@$�w��Z�V�Ռయ��F�5�sfF�or��a���V��g[�7mF����5ě،����ƬC����uu��;W�$���Af�m��<"�6���׺�4��1�{Jdbp��q�0�[�2(�sF6M'�}�Z�u{��<5+��4BB��pЧr2�@*�ǆT���O��� ߲�;lU�
e2�Ti�n櫼�X��m�ZF�m��
!�M*�ߚ�Y��l�͑�Ĳ�̀ӳl����!-����م�+r�L����:4����n��nء�������i�0n ��f�ͱ7"��f*kv�A����` YMSN�%3��|1KW�%^�)ʽZ�oaD4,
�]ی�i�Ht��$�ԯ4��7V�t`�(�wZmӦ�7t�ܡOjX��{� ��2�&4]Oe\��Yc�9�뒵9�S��ۤ��۲���<�����ϊy@��ж��o�̉e�4�f2�I���xS&���"�^�w�ִ�NMˋ^8�E�/U6��
�$�ӏ]K�R�$U�L�Z-�vX��\�R��bS��1-�[�.jv���aSEX��Z�V� Ood��E��j�8�h��l��)�i	���iJ;W��jډۤn5�X��b�V��P��o
w���$0b���WrfV���,iB�q�1�SK�n����Ha��OV�F�d��W/XhLX\i�!%�:�ڙ0��ԫrnǈ��X�J���LE��������WGp�,(�e�6���;v��wZ�L��oŗ�U�b��i*�@��Mִ�ʱЖ�"8Qu�s��H&�*��\[���NJ�6��0Wy�JQc��Р�j�Ѱ�聻�+�o4_Ѻ�@#�N�L�������jR�����Gn<5y�ki0��{PQ��q�%������a����V�c�M0�F�,-��F�^[w/o$;��c�Q�� 5�*�DN@Vh�
���#��n�kX��̫,��q��zc�/vL8$Em�:�&]��:zՀTǻ�W(J��W�F[�MNSS�CU֛����P�ںP�HS]����Kr��Ċ���@���[�wZΧ�F,į^�;1�vh^hR:N�t�lVje���&le�LX,;m����P"�����Q��%�5���t�n�̩TM��+t����Y�n:b�ږ���bӀ7j���˅�Y�th�j�n�\L��cE5Rݤ�2�lG`Lv7�z]0<:X�'��[sXH��wiw���t+�
���ՙ�)�/	V�m�ZZ/i�
;�Ow,�+��]�T�V��m( �=N��ǖ�\��\+7-�i	��
{�7�k�	��-f�1�'a��	�����״���7 �Ȟl,�"Z.�ʹ��[-��6tֆ��(=�%��'�[�#��[�S��-"�Z���3^�X����-�KcJ�0�tȲ�.X yZ�b��{����cJMҶk{j82����3N�kVŬ"(�1Rzv�I[y�������t�&�3U�-"�$;X�b���n�(�WCe+uZd���Sݝ�\���0b�m8[��2V=�-��O 3`���
;rRٖi��x�A�5�pEj*�peL�xb�vh�݂�5��Ɂ[:�G(c1]��(�W#���ë��7��1�S����ի$Ӻ$��n	/6ĵM;�O�+�Xu�K+u�8-f�tꠈ�i��v�PY���j|wq�ܸљ����� 4QJ�^�m�shc��Q0�NͦKV�4��U�\:�n�L+|wEV�.��0\���*x4EnD���e[J���Ĵ`� t��'�q�b���c�&2��Ch���!lޒ鈀���T�Ra/���I��.��[�x�zH�����z[��Zq��u�V��6]�"�`B���8��n^kR�DI��[Yc.Gy�����TjS˶b��uo�C�NkyNT�[�VV�7O@�n4��㥧bd�� �Y�&�r�n�S7 �z\U�`Y�24�����+9��[����݁��6H��l���`V�4�aD"̂�����hH)7�-v�����u.K�GwZH#��f`J��rE��7sU�ПH.���l$i�v�{.ٛl��sm���P5*�R2U�̔0j�@�QSy��Œ/��v�A��y@H�[�{t�Ҭ�]]�[�lf���ԗSt���ȝ9��݂�ۢR��m�y"�`Tցo/gh�kiQ͆���K��Cô�[X ����HBA�8jKsl������U��0B))���v�nՁ0�pM"�dw���f�*+i��GwNh��9��[�D�[vu�$�9O�ऴ���n}e����Ly�J�^�/pw��:�mgt�P�]����<����M�H]}�b�]:�o/+p�J�sZJ���1c���� �=��T�,�ݽ�b�4&�4Yh�,m+�:�mr�|5��JU�X����܎��w*;l��P"3jT*���XR�A1����Z��`���C0b��Tl��M]�m��;Z��K�heZ{H	�"2T���cU˜����^R���6q��	��0��wO/]�䣚��&˘�ҁ�q�,�p)��W���,ӓ5�wcVj-�ۣ����&�\��t�W}�>C�hObĳ1���7(n�k�B��XL��R��ѱKb�҈U�wp�震q���6u�. ��M1Yv @�Y�^AN��r�sd�mE�,ʬ)�V�HM|3;�7��S*��F�C�T�|��#K-Ռ���`��e�@�1;F��`��7V�c	]fnʄ����i��n�]��N-��1�����'�YD��TR�tñlB�֌���@�hlD��;��R�v�­ŴA!�z��pۂ� ��)nb�X
̶�ܘ@z�!���)P
����]��՚wF�݉�Y6�V��1II�Yj\��F�1g�0�m=z�8�-�:#+o.I��E����1 �1���|�%�،1���*�B�"ZޣI�x��]�ޭ�l���N#hfE��Dp��?lӏ)�r���%ͺ:T�i@RѼ��;��z�-o�"�jh��n���o!�Q,͢�%�Teج�D�	95mf){�Y��P���5;	�v�����6,S֦�Xy�J�[�����[B��u�n�^�QL�Bh3��3*ݘ�I[3)#5��mYx�j��5@�j�X�Q�\���c��ZȎ%�$��42釧�Z�N���f
o��G&�Ul�w�t���];Od���KC�!�٫��B6Jh�ninJz��8j9�&%vR��kQ�5˝gp�/k��97h���n�yz�.:��y0U��SaF��D�g�wv��:v��U�;�<�n���{�E?��d�#c�FS4��:ci�Y�+q3^ټM�pMկ6�[5�-0�ͥP]LX�6���b�nml۔���eD
Ѓ!��JMٿ���3v��PSf`�]�%��Rۡ��>)̂�:�Ӡh�3e0��X���6���mw&�?:l�Ul8����5x�ks�Q����`�dK�[���5�^3F����� �b�,J�.��V�&(��YC.��(���iy�K����*+L�v#���7� 9�� �a��lS-pփAVb�c��mY�J���Ay� �혍��h���~U[���(��%���U��ƑfR�ĩ�-�e��j��]X�*F�fM
�n��͍J�E��CVŚ86�ZI�Wz�oE)+5z)T��Z�q��]�K6Q�ۚ�ӥ�t�U=La��#)�[N�ݸ(�AtP܆�A�%��:Sx��-��2e�x����8�om���ʗST��]�a��Ⰺp��	�@7>��
�@�R�+u�h]��غe!��r���m�b+�i���\GM�#aG .U��zR�OI�+2�S��W��m<%�4֫#E5Q05̇U�0�)��5���Z��bLǳ4�Ka��j�$kn�W�����Q�������l�dǒe�/VAm�N�����(h��F˦�4ׄʲ��d6^̺oA�y��g����!�8�Qwt3li���y��r�VX0��J�×��,2+�W��U�o1���oC���%ޚ���4���5/.��T��;�5SdְQ͗��^K�J�4�9��SiF�֪�z71�$K�����P��b�h�W�:�.�0iOH�k�xVJ��KF
�a5��ni���s�#[jhY�f�[xfh�v�*�U�ZU:)S���r�].SC;u5l`&�bJ�I/ha�F�l�g9���1�A�\�Hf[e|��ͬ&T!]i݇3\���n"le�A�)�׻e�dF�$ȵ �0Bj�W�][���^��q�&�!�	L̦�H�Vl��f��������P�J��Ӣ���
B��F�ʆ�5�JM݉�h�AVj�[>X���n�"���Pְ��\�p�1-z�p�3P��`z,�;��7�E��*q���6Č	zma@dC�z�{�w,��o[���Su�h:Yb�]��h���fA��+��^�21ouV�Ô~2��+1@���2'x\[�����H�Ό������x�w��U�l�5;���pI{hm^]kZ��lU�4��J��Rk`MM�X�&n,�r��a��/]�th���79M�Ѳ(>D;�*'Y*i�N�i8���v�V���W#a�X�;����Jy �3 qcz�W���YNJIc֐��D�X-O�:�m͠qQ���t
�SU)�g(�B�b�W	���c6���9(J�e]F�Ʌ��-ҭn�k�������sE(�:sh���p;XqŊ�����p���Y&�ԩ1��LS�T�ӫ,Ӏ�Rn�vQ��[�((&�h�d�T3U/�
�:�on���"3>D�.�����mحu��OUE����1�$��b��*q�^c ���7�����A|O�zNi��>�-�:d]@�@);H�ͱ�A�we\�Y���0��v��8��	3;]�pP�*�bN����􄷕����i��=���u��)��p�蝃��vk|_SQ�:��C�ؤ�ia���Rr���)�
&�ӭ�I�жr��<��h8��I�JwE;���AXDb���ֲ6%��350��u:��{P�VmӠ�*^Zv�QO�9f5CK�f�V�u���=�8X�����k��j�w�e#{���.�L1LjW��v\5k3y%w��(� \�]�Zǵc���}��6.��Lc
O����Hy풣�;���Kh��H�Vz�bQΐN�Q�u���N�[� �d�� 
A���G8�����s��n&�����������pn��T�ڰb��<�:�����Ɍ�L�2V��>e�������]�wTNjm��i��D7��s�O�F�Ǖ�JQ5ČJ�M�ɾ~RC���u-U�z��p��C%>yit�: �tgF�Ö��B��s:ܰ�h8��x��e�����f���5���DKT<͸ji�[I;�W㘢��i]����w��"��/w�F�*5�±u�JU��+�+*Q"�!R'P�~۱�ܦIuѡC.np��4u]p{�`�-q҃3��Ɵ���x{)���![h:/o+�{_E@�>;�&@������� l�"���t�b@o���S��]��r�Er�Nb�D�͡m.���T�H38�5	u4��.َ��/�c��@�*��n��@41Q�o 3�Xԉ���ʒtS��m�D�S"�Ф]u�ܗ��9��#%�/1M�*Ѥf\��V���ͥt֕�p��ta_�K�g[�=����R�+���t�U�Ol���!x�h[,�Gzƈ��]�^�5M�A!9���R��lH1�}ѻ<�ե٬V��H8.Z��
��2N��}�36NYx�0k��.t(�©�O���c��I�$�X����tI��Ye�L�aX�JN���Ru��*�A�\+a(q�M>TWR]PKA����0Vq�ħWWJ��*�v(���8�7ٯe$�ˤoOh;M��׍aȊ���*�z��N�6���`���*�F��~jC���w�Sc���=���S�ܱ]�J -������vNky�(ퟭ�%�kk�¯	!��k�Q/�9%�m7]a�32�[�F�%�j���ʤ�u�׋]�����^���,�i����*�F��kԘ�lW̢{�qp��T��v˂�eڐ���ۤ넷>V�ڋU�Eŗ�X�:�J����)�8�<+~-�)��}Ƭ��Dv��XńZ�ոN|)vaV'8�+�-��g`W��`���e�'�*4���J�A�H4��	�B󞺘��C�S�շMo���4�u��\�RG�uR�[�Yd7W�4`���e��v�3�L4h!�]h5�~�;sZ$ChĘ��.LZP������gw�G�u��m[��n������f��j�)�}�s�%U��תc���~:^�W�f��s�n�sum���2����1�e�JT�C)>�������j���mP'�jY���R��U�os�@z;5]��I�뛤S9�e.��fՑ{ږ�4ȋ�3v�!î�&�����z�j�i����E,V�Y6/�v^�)\��q�W������e������Y^��ﻢn֪�0�4��]jޗӫ�"�=��-g
�E���ӣ[˪uwH��v��3\L}�U�ΐ��B�L������-���W��D*vw ���I�=��n�9v*��:-*�[�N��}�2ք�2�T���{ز^���W�f�F�����é8�)���(uj�S�X�X�Vyϸ�mP��J@��ۈ�,T�XU��p�]�|��+Q��s�#�/V�Ӛr�Ѱ�'��D*V�Ǐ�9�f�Rƒ�C{j�f��;]`U�|^E� �lD�b��pmՃmjם]�	*�_a����i�������sd�����&jV���wM99v��c�F��[u*_d�N�2���B��ۉI�����]�%;1R�[xW3�2U�+'P�����w��h�8u<����:IWJ�S���@���i��hТ����#<͸��I�ޡt�yҬ \����؜pۗ�њ Ԗ3���d�����鴆S9r�X�֠�����,���p�$yy,.�*x�N�`���7|F�W'3�.�(M���.x��4�-��ÉQ�Y�겄���bz�2�£ۉ�`�p�($���s%��5Q��A��{�"`�6�Ł�]}�tAR��DH�\*�_!�`�:�t2���$5�Y�AZ:�t��VS�����\���B��X_x��b�SNpF�4��r3C5�au�i��F=!v�M�;;{"�*�LQ��i[��v��N>��Շ��gG��X�c�=���
�8�*��^��-R�Fe<�ALo�%"���59�U�B���V��}�kW�E�S9A��k]w�Y[x��EK��koQJ���f<ݭ�@���E�7�	hn���g)��Zq��Vq^<%��kY�u��.Дf��ٜ/S�_BSΛf� �C-�/EbvlX�hJI�I��<��iSxA�+�-��R��{��ޔ,]x�h�5Ce���1}�x��ci&pT��"�k�ִ���銍�F�@2�n��mvE�4ksl]��;%5J��UȘ��ie�����e��%Z*r�ea�{n^)� �h�S-��p�(�G®t�}'|����I���M,�aƀL��$�t��:��
3�y;f�)��`��+��#�uՏ�� �(�!�0&K[+Y�b��l[���7f���`���DW_dA!�t�?[�w� �7v��u�t;��Ea)�4�ҕ��G�>�ٛ�o�M^ns��uκE+8�+ORY��z�8Zt���[se"U�s�yi��6�\1�#o���43������on����;�ܒ)9�7�H%��A��nmC�֛�|�V�w���؊�����eG����v�-�sdB�]l�NW>�� �qT\�?���w��$�^nQ9ci��/�9=��;z�w^z�V"m�%&s�t��[��`�ޙOX���Rι,��TIAzd��(��jQ�1إP�" �i=)���:��g<��K�W@�D�{!լ,}�bὀ,�4_`�1�1��ۼ��e�7���'Wm�N� ��{�eڸ��x!�U�Bڌ�f��"ݸ�n�������9;��\٩���ؐ�Yj�<7�h�{�}D�o��E/��CN����^ݦDoZ�5�V#�#�^��Z��xf�u�l�=�'ܠs��,�#wYޮo2Z�� ��Y�¾�)�nV���]݀d/���S�����*�/��#���T�ˢ�K�������x ���������a��suQ�pY��:@Ԋ�cj�!r���y}{�BTy0s�	�Z��Q&@w�JZP���j��ZȾ%*'�8���L��d�Ӌ8��ᶨ���������_3�;� �T]�RH,�L]մ�,(�mU��a�Yq�����t����$q2I��M-�T�W7Xi�ױH�+MǶ2��36)���fiܮ-�9D�!��g{)�Ѥ:��Z�1dDx��wv���_,������r�D�7�b�y�V�g]^�YiL�ux��Os���E�[7m^�|Λ�7��>N��{�j�+[�����r�0��)íb��δ���0�U�+�ۤ�n�1���b�X�"�<w,��d+\�A(���m�Հϥ%�7�NM<�kf�ѳ�Y�ԾV�WF�w]V�ua>�ѻ؀��oz�KwZ�O.B(er�6��8hl����\��a�Ƞ[wI%�_7GZDrW��T�8ˇmǚR�H����S]��
����.)�QYu=������_uC���0��&苚FEܺѮ�)o^�W�	Y����a�y8�\;�Y��)Sk���8U��ls�=���>ү��ƣj�����ܗ;�@ԶSM��knūB�k����U��s�
�+��vwh�{����xB�3W;��U��RL�9���"�y��h��v���.��$��X(=�-#��d}��#��+5[�^�K4JOylu|BÒ���A����38���+Z�]X���K|�0�ю.�݀�Ñ�=7���m�B׊hT�
}tn��S-m��#˷����f����xW]����wZA��A�-�[4�W��gy��s>�:�� ՞Q2�54DBH@Sbt��lC��P���zY*�J���t6O
�ukt�
�:*X�����r��E�Zbɻ�n]]��j[[�m-�J�b�]h�Xt�vCw���	<)ͺ��|�:�HM�Q��4���T�Z�a����&vuY�%�otw\Zh��+�3J���L�}�׺�9;J��zzX���Q��]�76޻/�˧�~{jS:&xo��v]4�wf�ˮ�k��\�D�0h�n^*�9ᥨk�r����\� ��!�M�-� �}$y���dp6��}����ө�W�D�z�Rծ��Kͮ�ʐ�2dN�*�u�4T.oaG���>o^�VKy2u-x+�e< YTq��)���jEP�ju�w8n�}�
!�n�.�Pj#a�����Z���T�D��y�:� �9�h���*���J�Z)��KS�����C.K���'���82�<2}֡k!�ƚ�[�}������ӫ[1�-;��M��F����gV���b	վ���^�CWu�����S(ò�L�j�!ٸ��*Xw�$�� ly����G{���C�ԙY�}h>�i��ͧ��w��F�qf�B�mc�TD�ei�;U��K���T�.^ԅ* b�q$7�����bdy!B��Vhh�wu�$��h���]���4+�^r�dV�[����Ĵ����y��u�Rq�_4���B����ye8�j�仪���;[�ͫ��KGE�a�	�cv�n�i�� >��T�&�m�r��+�:Gj�1y\N��(ԭ���V����n��Vk��N3Z���	aK��n�:���pwAܣɠ�������F��1i:F���Xkm��	ưS�����ӷP4sC�v!���� fA��pѸ��Y:9�뻕9�u�40��P��ڊ.�sG M�1�rpz�ա#���ٸM>�a��;�Jk�7�"Zת��$�n���"��]�Crj�����M�1p��w�d�K�^�FU���`U��D&��iڻk����e��R�Ƙ��]��v��F��@N�rW$ĭ5�H���(�}��v��>�|�F}ƅ��B�Me�0�j��:�6z�@Y=�9�k�C˷*ڪ�ﺗVQ�
��t;�d�"J��D�:}�~`f0�LS���{�^�I|/TIѭ��({�
L���{�n���V�}j���<�i�׍��u;e\f��q���}��]��Ga�����o�*�p5&.G%�+8�{O����>�nK�~m�P6��#/:�ҕʄ˧6�V���Sxwin�<,5̩OjH��֤�Ţ��sr�P2�*ۿ�-�`�W�fiĤJ:�:�lH��f�)@��)���F���Fh:5˔��t��8;{h͢��ͥ(I��D`�!r����t�����%���;º�Z��v��0h���Gi�M���[�DĪK�;U�`���S1���"�`�/�qJ>�F��u �aP�X葱�	�t���/vR�Ի�y �7���<�F�e��M�;�0ĕ��{%d��ik�-<�ک)s�x��3��i�~�|e=<�[�LR����⤢L��T�坏���+�wh�A��^�Ze��v&4뉩\�I_%o��M�źxu�"���ٴ�Ua����M���y�4¹r�Z��F���fc4��ݦ����Z=��eYj#eWm�C�3�&Jgz�b��ihk|�6t5;neɸ�(i�U�bj�B��YM�L�H9U�"W����!��]�i�k�o[g���)���md�',��@N+ ,���+1��.���U;=�}e�tl��}�F��eM\����!w]؇f���X"�5�IV'�K�a�Y�y�WS-Ӣ ۑ�Ղ��'�Ǖܚ�b�fHL�Y���t�;K Y)E�ƚ�lv�#�{���U�A�}QP��S]��mc�ִ�ͭ�����HU��ߓ�;-����w,�\+I���ؘ��#��r9�і�9Wt�zo�;�u���I�D*����r��s�ۼu�fᔸk�,�[��b
�����FC������Qȥ�
����5��5x�������آW�Y�t*�wnH�eN�b�|�a�/���L��!�{�60�p�m�-f��Y8]�!���Z�����R�����꼋t�.:d�Cv��l�����! F�u��`a��?8^J/I�����|�s�/]���FlY��ڲE�Wd-�T�SM+��΀k�dͪ�(9l�{X:��`��C�e]�����T�ɋ�Ԏ��WQ��ݸϗ�s��".����J�s]yP���ŵڨ!��,G�ɏtñ�t��`���]��M�K������qMK�*�^��)�a�8����'�V-�3��<��=6�����s��c� ��F��Iam`�'6�@�e@��t(e����N$E�I`�0X��-`��r��H�E��7��-����Dڻ3�d���m*|Pܩ�9N����ԩ%�/;�r�J�T��U���oO7/�o���;� ��;���-�Z.u��)�S��SYҝm�7.\�_d��X�z�c��"�vT� S��y���p����,2� h{u�)u6�����r���;���p��k���X�ַ��`���C m�`���6����1����_P���!�;���R�T��wUcӡ��ʗ[�*�s��9i��\�9�x�ϲ�N�?��l}m
I#:�����T�Iuh�y9\ͮ�ieuY[�V���	l��oIcEbk5=9�u[W3]�GrcJ6z�[J��R�.�Uj�7л��I#��l�t*2�lv���l3�CDI�y����\wo8�f8p<�H�ajs�*1�aZ�^�����(��5���i�:�Fc�4{����U�e�t��ȫCg�'~L.f�v���od�wm��ݷ#��L�-V�ˣa[�^�w��D�-��+�MQ�8�X1�EN�!̡���R�kNC���1
�FPsM��.Y�eMٜ-Q
j�o��I��&C��ʍ��<7wE6^DW,q�&QP�bx@EƳL"�e��f��ֺ�Jbk�8#вT�9(��En�[ `1`��.�Y:��i��M�[Z���Z���&ե[�i���<�sN��C	��桤5�>�f$0�ƣ�{�;��U4��q@j�e䛉��S�Է�U^��Sx�-��#o��FsQ�����/�V�g��c��	��};��=9�z�m�wM+_h\KזwC>��ʟ*�{W�qٜ�r��SV<1aD���P����+a+@�[`����].�k��]Q���G7Ҹ�(�Ãq�SH�6zp���8,��KMC�>�����h"e\��qV�vE9JlN] ��%�h�5�|��)^��uhG���V�o^�ޖ�t�5�Y�-b�B�o�n�.��H��Gr�j.�ٖ�R<'$�x��Mp���B�4�M�p<=��*���sivC�.�F�J�N��ư�i�<qI��R!ݮCE�c�9,k_��9ٓ���22��7�6Zoe�9[R?-sm>,��uU�Z�ʮeJ�������"%U�X����B�р�ky+t��^m5��4N�`���wyHD��(X�i��پO�c���uj���T��>�;l�6�W7�s�oh���iQJޅt�wP:���_F:�kXe�h�1N��H�}�$)ovB�z�-S��u���1+��P/% �KQ��hSZ��EA)�������˻n��#r��fӒ��Kq��#N������� �9swvk�X9O�c���)�:#MAvQ�w�[������mNn˕d�s����Q��ؼ��Zz�z���t�k��3SsID�-��_b��C���eӳh6�Z�b��D�ys��
/��.��Q59Br�kot��c緝*�{1+�Mp%\�`��廲��z�f����e�a[u��t��ؕf�+��ˇ�j#`��n�*[n�t�1b���7�wqkW�|4�y!�N�9�⊅�N�tr{k��NH�N�\��uɀH�7!�e��!<�T���9<.��b�f؂�������|�q�2u����)B�j�}��ʹ� 6k�Ε��1�c�]2�؅��g�5�p�����c�2�q��m�w,�MJ�1t/'$�s�sj`���P���ՕZ�޺Aج��S�̓�7�&oQ�}�s��!�z�(�:�8N��JN��Ӗ[,+N�A�����'�j���眯�9�*��b����	շ�VྦྷV���b��u@+��R��DQ�Z�����t��ʝj�:~u�Vi����y>z)D!�^Z]�H1������/"r��3�+{��p��E�d�C�d�0.{��>b�3�k��w}�,TE�Q��k�+����7����X��*vT��"У�X�fڧ7Zd�*:
Y9S��i�� ��w;��2N³�8��Vw�e܇p�s��M[�}�W`�K1!B��s����=6�;#�z�G��,��$�D]��B,gf�ucыj��:]�EA�>�+T�n���8,v�w��h�b3�sj�c�tw�ň÷֧�L5{X�b�@�]���	�U���1HJ��N&,i�U�u^hZ�0i���
�]�U9l�Ւ�;��;(�1��B'[���R꼸�k�t�ا�&#���WP�*�S���)L[�=yj��4ڼ!�� ���N�n8�
B���5ePZC���Ψ���� ���MB�#�^��U��Vz��%��K(Qr�t�`���9����K+���N]�[�Q�3�(j��T��.�����9�d��l�[3eT��T�3$-Q�Fq�Sv3���t�jZИ��ֲ�;�q}�;ݮ"�u��ՙY�tJ�������)v�8�%��w�;p�Aˬ�}e杔��W�Pk"�z\��M��[{n�7����2�zI깯F��n33�lMíP7)�K�>#Zͦ'I���:�%��\�WY�_[��ҷ{�tn���͍u�o9����)�;	�Fe�U؝B�Ϗ,���i��;�R��\�ȯԩn]�y�e���3�ԅa��%ֿ�qT4f���[�5@�(��26�-�*�z�tC�흹��k�"�.���Б�j��L�[�mћ�m}Q�xS��ě��L^
��YT��@�NL�����e��֊��;�bL9��ړ����^��n��(��!�V�ǜ�<���M޺��RN�n�k��ʲ�9�kJWW@���o.M�.�+�� 3e��Z��^�Y�0��\��_[���C��n�M*|r�&n�s��ރu�%u�ʚ钶�	z�-}�&j�B��1˱�F,>|�si��L44L��.h�rUj�9�i�ڵD���`����Yz�T�tWy�u8��ZӍ�/�m�ѭ���?5�8eƺ�������kq�.���d����;����hb'E.���]�I�M�!o�H�ݻ=V��h����/Rl�6(�vlm���5e��cvkJ�휀sY��k��ʇ:ܻ�V:�h[�ޱ��'��5&r̡7yw�OXn�l�������a,��ɳ�]0,dO���/�z.�t���B�f����wcr`g;+�B��oU��ؙ;�gL��r�����y-;���9w����7�>z�x�E�}�m&\�R�)��V*�Ɂ&�!4by��M��l�;a�˻
�!C�m���M��ݹL�[�[@2�9Ci2�+E����_Q�I:|9#��(S�4�y6���t�6���G��;D,���0Bh�<��K�P��S�s�����h}�K�99,����(�F���J;�;0�v�6��n�F��v��y ͏z&�˜S���]s�/9�T�	����8)���8�S�!g�ì���b��Ր���R�F=k�-��г�9ܵ�Q�w^A�n�(��a��-�\JѦ���,K�%�`��7䷛+k�8���]�F�/��#H
��i�ҥ&�F�c�EJ��{أ᪄����0���[t�z�97FG�r���.��nl�j���=�\7�yz���h�a'�y[6o!Kt�6�i�X�,�ǽ.Z���>固�U&`ww���3E�(��B����
Ăۜ��9}�LyR^�EX5�Os�����-�RΠ\�mT���I��a��ھ��L�\n�.��5�0s�R����5m\�- �t)�aV�@�X�f�)���׽i,wc/MG0�7�T!j][J�ة9;�������ə6�&�4[6�Yx�ҽ�:�W0�n�B�2��կ"A3��[�w�xS9j�v��v�4/-1R2 	b��8�n�YcP��V��:0�la�f;�B���]ev�u-pJ�Դ����g&U�_a[�0�N�E�������e�Ѥ�ؕ[1�.dM�k�ޡ)��H,��.�뫲�������H�Xl�Jʛ��&�Q܃��܍`� aQmspp�����Փjb��uj
�,������[A]�y��Mn���wz@�`i��O{OXn��f�W%�i��I]����7[�PF��
|�u��d7�6�&^oM\�B����u�.#o�!p�ǲ��Ʈζ�˗C�64d�����qQ5u�����org��2v�hB�MOK��ǔ��qa�&�(�_WK"b��@�gF�n��98�I��gi��;k3M�ʵ��}VyV�q3��|՝�Cmb�Q�RJ*	hU�E��n\���ytGn�@�\�yP� ��S���36�i��C��ٵ���֮��y[�J1�Qn֧�4/����\��X��L��b��Sp�yb�z��.�=dܔ6�@�	�����^��ת��A(ć�S�淦�iA�xP%%���R#6�Ԟ��iwF��5��������n�r�(�"-y�R!��5����ŔSF���Y��u��kY%����RA���*�ǏBmiʵ� ��«�ѡti�vn�bۧ�菐Ȫ�4�oh6��]�-X���$q4NݥZ����9��n�f�o/n��}&1{�k�S=�U�A��J������\t��)M��2�#+�Pf8S�
{�[2�Vik���l�W̼n.���6A�Um�g�bK�_2I��>��z�"��c�S"�YoK޹-���f���H#=5ٺZ��X1,��g�+cC�&eQ��ٝ��;���f|�~lӥ�)�A��KK*OsNZ���qfґ��nҧ�K�-__;�E���䄮�m;U%sŮ��l���
��[�4��Ժ=Q.�(J�s'�'^+�-q��N��V����S�M����nK񜆒b�������鷀���2}(-W+��*6���Ķ��nuH�h[��Ê�T�
n!�m�CN��n�3��Xy����x��p�n��+�qw��7�kr.�H�+��������u9]*췵}Z��RbE�[���:d[F�:�{�2�h��HJ��J�R�cX�j|�
#{qe���<��1�����~�_j���]m�q	]�������}b�<6�U��^H�B�=�})k�ӝE�U%�yy
�3���@�����.��N*lNi�e� �]-���F1�v����M1F�u��N�L��[���>ݚƎ�j�৬f�.��V�	!��!)ۻ��O}j���t�F�4��֨��1>R�E1�;�>y�Rj���F�e0���51[�T�[��Q��J�Ѡ8��ʵ���ٷ}J0YXt\6�"p�jN-
2SCK˕ya�J����m��U�]VLz�Y�X6�i]ӆ�ĸ��Y��j܎ka֞�YJb�'�lL���FË���U�M�m�׷�uoũqr�Y�`�s����p#[؟r�8 $�ۼU�6%�ƴ�%@�ɘ�R8!) �T�B�9��,å����3(�)�tqn:�v���ƥM@U�	�͹�b���*�r�h�ԟ_�������{q���E�{n�
L� S�˭��\�la͡�S4��]��T��CA�Z�ܙu�*�ޫ	i3#���i�G��ɹ�A� NU6�{�i�n�}s]���;���j"Z��[�s���<p�;���з%jN���\��"�����"�R|��!r�NP��QP�V@�w�N�c���׈1�.����GrD���WAbZ�Cv�X�U�%H�+z� �����T
{�6��Qfu@�������;BEjQ㪆 0ᢚ4�gVސqs�a�̂�l9c��Ճ�J�b�����H�cyY"��m`I+����,�q.��l5�7XM[��k�M�Id�͸y�Lݝ}z��C+lř\"A5�����v :�K6'b6���x�yFW	�ڹ��0����sNW��]��iv���tm�ŷ�b��D�%����
V�\����JܸW�L�mH��zS�+A�z�9yR��аQˣ,�j�-8��KR\aՆ^��0�՝G���@u�U]�/��n�C�%!�u��5��W�S�PB��}�/N+(l�+qN��\k��k�T��Ѵ�l�P���]���Y�E����:VT�}%�vC�
���Lږ;\�k�.Ds�ͥV*�B�@�ZV�+$Ψ��vRWWt퉦�&I�1rX���N�U�'kq����G��kh�<�M�[�%���,/�ۈ�70�ʙ�F��+x5q;'*�.����D�nm��4�3km���e�o7���=ų����n^�Xa��O/�8�Ǯ:Zâ�K SNƹ�t�D�����)Y˒��t*} ٫�+�!
]D�i�M˶�S�����`¨R��u�0���ze_˫+�#��wY���\�U�������o�J��JR����Ċwf�6��
k?v(\Y�1^�
��!�f7��4`f�<��^Z���ZtĴ��st�Ujj�W��>E�gss0HF����Y�:�[Vŭ | �< ��wZU�]�l�LnM�؍�4:K;J��Z�[	�N�U�/j��5�rHWmZ�혆�w]vG�9ݲ��j��K{]�K>�JҜ���pa�}�	|���AE����S�hV��u��7e,��Z[�-0�YT5��\y��/��)��Ś�87���l���W*0�׉[��H�jc�����rW#0�լ|^u��ś{�Z�x^|F��^�;���+n��<l���]p��,p�->�Վnt�v3nM��gZ�<P�6�<�X"����ʙ��Q������i[r,���v�ً)�$@���r�g\�b��we�2��iѲ䨔
\�a�iL0.����#,����҃;�J%���|$�5}%��t�]0z���2=���G�Dh���A�B^)��ě���v:5���,�����G��nR@�Y���Ζԇi�:�rM�@�/���ݫۡ�uwR_C�9kԁ��4�L��a\y���+8'L2�ه_Z�F��Q;}��v4��#�z	�!��˿����L�.o3��*����<
ëA���=�;�'��:�q�h���J<�":ҳ\��[�ŀD�ו���t��\{��d��,Nؚ�!�O�
`}����Gm�˾cǥ�j��{y�Q�@|:�]	W��W}��P��Ҵ�ɢOW�vɭ�Hl�ؙ��k�,�\ǵ+���9P:���b7��A���7��딹qSms�k���]B�HF����aRu_t�y�ͺ�Bv��q!d�W�N]G/rI�*d|jIY�7	��Vq/ną�V��T.U�A��|�����l��ѓ�&@X���oqK�6�����\^��\���lTQ2��/50��Yggu�u9Ҷ�On7�ά�)Ry�tm��	��.�C`�0��d�y��[F�	��n�2�Rg�F��˺�|�<�-��eΥM^����������wύ.�]�a�|Ӝ��֦ zۤW,k34�*d��7��t��sL��-��"�z��F�es��Tn�J������1�ɪ���@�����I�_�z̒�xA��`�+#�'�Sb�5�.=pӷ�:��h9���j!��`Yw,�D3ۻ�4�a�SY�ɨ�t���Y���0g�߅���b�����B;V�ʶ�v��4i.���S��S�E^:<3,��p+刓bw4ګb�V���:ݸ���-�'kn<Ĭ���P���XEO���>o�=ۖy�s�;��\�ΆZy*��nNBE(�$�O@����x��:�'/=֘tM"��S��R�\]�M̍C�Vzݗ+�壡�.k���tN� i�E�'V���"�2�r����N^\����������BO]��"�s� �ҵ�������a�p�	������w;�ո�Sww/n�����r�������Q�Ht���2��v���%�J�H�U r*��< W<��$���ե�P'r��S�y�"��w=wt��q̧E]K��K�B���:B�@ram�D%Ҫ��=�@����=-��P�Q�E^d�iY�/ZN��q���Γ���9�z#����������a��b��2]��9��"rY��L��8�܏X���ʋ�Zr�v-���:���%B�y��~���&�޵%6���Z7(1�r�[:�<��Y��Jjo�z�i����Y��J܅�#ʅѴ��\�hL��S5��̺��l��	� AY.�%5AK+��5'���l.��~����1�?v������]������%S.�ɫ�ֱ}Y�w:ѸC�敭��T+����\Ul��Z=1��s���/to�ԁD_�FW�R�y=-+\u�9�"�V�H|�p*�BI�Q�Pa02p$y��ڝoVӓ%5�Q��8Q9�x��8�T����'��v��~�#��(*ﹺ%���E9aɽ�꺃�)��v���p�o��23�i����T�܅u��n�W�cEb�^�h�͎{�T%�!�N�������|/o��c�g�����J{a�1��7V�mP=���}�n�w7b^�V��T����Pl�(L_r�Y����>���s¢�k�h��18͸l�jXΌ�_��	;�L�'���]L�\G\�Dާ��U%QAf�,�RU�ﵳHЗ�}�#��_���k�K�M����� x"x��xR���֓+84�ԧ�1O9i�A��g&�*)Wn��6���c�vٽ�]�����k�yT׽N��Z�&����^e=g�SV7p��F��*�u�5��@C���zԺQ�M`S��F�֖\:�_k�a�:ƛ�C
pb�l��w`�":��a�.Z�䃌���P]���X�E7_������;�F��װ��Q�(�t;�d�jU��U9,��NP"Q!�zu��
tEbu�FKj���P��:�&�z�'M�g��'E�vͦ��Co��K>�EG�^&��8�f��W*��o]��&��-�&. 1a�t��َ7j�҅ν�z��W��+����y�ڬ��#j���s~����5�􆽂��iJ��mTR�f��&{'�6�E�%Ȩx����,����0���w��0cxfQy�Ht��'���y�k,���%
{�	Ρ� �!)'�U�*|-ʞ�����>����n7�=Ʈr�q
c�ֻ˅�	;�cO�M<�v�mj��C`��m���F��ɖ@~^V�6���J���Y�l(
ڤ�_�a��S��G�����W�8s^·(b��y�痢c�|�Ն�u�S���0��@
�q�1h�:��u�ŵ47OC5y�*�S��}��W�*�E��'v��<!��&�0S'�Z����q���9DU���3[F�i+w(�=�Z|�	[�����\{�G���'���B�=��� g{���}�]�m�|��gqTK�Uk�H��u�r���y�$�cX����[�J�]ݦ3������{WqZ������2I����v�W2���е�����1��ڡ�I�.���,�7�%�O1�@駞́=ʯ@��\ۨ$�2y�G�l���|Sj3��eq}�/�9���޺ᐴtm�$Ң`�	h�iz*���l���3
�\ABL8�]_;ҩ�pX�7	�e:u�q���D9�����t�y9JF�Ǟ�T7Y`<�n_Ԧ(�N��\9Bف�j���~�B8�+^@���W[��t+�>AY'Y�c�Z$Q0���.�),�"�T��T��p��6��T��~�h*G
>!�h����:kk��c�,�ܲ �8R�J@Hg-�c��b��C��q���a��O�3��������`�*��H�p�8ҡ���Z�]�iY����b=jV���'��K�V�|<���TQS��d��Bp5�-�,>�pL `&xED��:7P9���V�C�nw��P6�h�1����p�s��g�>WĎ4��*���	�b�ɠ왼;�M~�B����E-���R��Rb��f��s�ѨȨ�xd��(�9�)o^�*�1,�%��S��h]�c�-f�VO!+u
D���+�V
X����d�Uw����6�9�Χ�pM�s�u'����B�v��9jc�C�r�8m5��壂�Tk-���j	Sa��w�f�hD.,JI�[����\߶n�ˑ�ҕr�\�C0�݂t�k��4+(�e;T\�И��ڍW!$��_Ȱ�e�'y��1��TkQj1±T&��w��ޙ��*��k�U����ף��mU�g֤'�Q{/��kmT�$�J6��1�1ɤ*���`؞7Gu�_���Ū�3�e}�}l&XЅ�d^��QX�!��O���F�^����Z�-��p����p)ɝ:j{ģ���S�7*ޅ�h{�3�f�}��p�/VOv�d�t^)5�S��!����t҇��M8�[nK�6&e5�#F��ҡ�sfP
��1���@t�r���U��BZԕj�#a�f5��>�Z��-^�������TY�Յ�]|�r�sr��wR��V6���с~�9���>y��S�~�*���&C�S,}��T��\L!���[4�CVWj��a��Ψ��tשB�b����'`��!���۵�DC�BC�lCd���R�>���-p�L���6�D �MP�^�;�g&2c�s<MC�)�N��|/����甯]����>=Є�zp{z�9="�X�mp��ep�Bn)]�AR�P�$�'5�vB2j����m`�2Y7���h�r܍�u5�Ʉ�m���@%���6��<5���
����L�ɸ�q��5wrE�|se[]p�&�sv����mvN�I)�y���o��9��H�eܐ"��!�ȋ���Ԝ��/r�x,Ѽ�J�U!�Ʊ�p숔� V��.c6�&��28��|�~]3f�\#:����s�#�C����}P��,0��o�]l!��e��b�*ٯ�U#X����N�!��β�%��:��޹Xb�$�rk�\boz�z�Ha@}S�4����e��ֻ�\��ً�ʦ�Y'B�@=�����P(M#֫)t{�Y�2s*�����6���k�¢jt*g��[�������9V,<?	��C6>�ٶ���6��ǠRe+��� )(l��,���Z���r��Q�+�sJ����W]K?z⪶~�+=o/Su�&j銻���kw��TJ/�r����vZYk��3�=r����miT,�O(W_��W嚶��8]=�}Ԍ�qS�~�<Q9y���Ʋ�uN�ȟb���o�~�j�8��7+)���~�G�\$� e�>�<\��Ӡ��	��|̌V����w����ۚ:�����c�b^w)�;��{k/���Y{ ���-����U�[b�۬~K�xΙ׿���i'�h
#��m��((t�짳r�O�\��fn��z���E:@��=m��OI)w�JJBac"���s2������&CQ-O��c��q��'�ߴ@$���4=x����w'0M�tH�׎Lb{�l9�����zq&���\7)v_�-!���$�h�W?�#^�ի�b�n�uxܺ�Z=�=Z�E��j�����e�l�jXΉ����P$�D�~��L�l�یLZ�iH�(��q�:�=:�eicD!�:��m`�J��Mӎ]�x+�Q6�ˁ���c��r���l��w�F���3�T9�!W¤�#r�a9�2��ڧ�$� ����D�;-��
tF'<0t����;�Cs�븗��p��鋭��@b���M���4<x
젴�3�3�Q��U�95H(-�&H�T{����Эb���G��Wqd�]!��u�Di"�Vӣ<R;}�+��֍F=Ѿz�5��,;XZS�e<]�;���E��s|�u���.�_*1�yoÈ,����c�{�p���ʽ�.#�u�q	���y�F�t6&F��{q����!��'L�S&1.���lv��	�}����*�apU����}��W���J	6}��3¯kϙR]w��Gͩ����WWƷn5� 
��ĵQ�΂������&�[�;\�n�5�'r5�KU�䎶V<�ێ��9����C��_i�U�M�P�,=:���?8��h^l��Z�.$�ь�}?94�u���v�����&��J�5~�S��9[���)�4+�:�� )%����C�*}������|v��x,F��7���//�gj2Ǡ�n����a]L=4J^u��c��u���)�n�>I����զ�~~`+P{���9{�O 	o�*p#��k7+����! /�Q������*P�ݜ��`{�~sJ�wd�^��8Y��,5.�J{�����d����n�+i��I��{g������:MG)L��y1��n�s�B���踽�L�ؙЎ�{�2�A�K`����]0�mP����#K�`2��Br�Y�m�B���c���ai��Smj/�k4��L����(!X<�9}s�\i���\k�Hc0�m\>�8���y�}�]��������>�W��+�@�H����K���J�H�K/�SF3\��
w��-Q�"\��R�YB�L��.�@,;8�N��T��[C]����}G�U.��J�s�S���7Kq�]G�0�^�l^]չ(�CeӬ)d��|�� Y �v���_NΖ4�C�u9�e`G%�6vc�@N'��k31;gi!�'gfISE�X�n���y�$�e���K6��f<�*�]�ԛ2���Rfo+褴�Gd��Lwt��V"�:�%T�q #���A����ߤ��4���cU�cN�KBv<]ʏ��U��8!��^Vm��ds�	ƻ���(}�,�$o,"�4�C{dz��׈d�}H8=H0+���m�p�.�d�&�؅6��2fc�LmAi��[f��s���i�va	���������C�s¤�G4�Җ�p/�T
oԝ(����bC�ZWKe��Y8�9�jVb����8�鼏��7UW�l$��_Ȱ�',	.���;�4t��7�'�0}�f4���t��O�yf�Z�^�?1����}����+^U=�:{qH^��/�X:_r�vЧ�'bx��\��	T0Ӻv�p���b��r�2|NB'�J����?F#9Y��ڭ�B�y�(��E�s��(sq�K�����B����6��B
�"5=P�V
�{ܾ����>8)۩�j��l;��gVV�R7.,mEg��n��4�.�ٖ�5EG)L�q�6{q���jW�l).���^�ȯb�5ߌ� W�xw�0�"�2�G��q�.�P��(]GFZ���s�vww'���nI�E#g.�*K�;v7]�j���šֆN-��41Σì9m�m��dp�7���K��c{�-ݠ�jr���݆Y�:pE 3����{j9��]��%�S<"��VF�V�?�j!�ʟ{K�G��VQ��r�0�,���=1�5�ia��h
�G��TT|.�Re���%ة��<���pǽM�Z�9O&v�j1��-֔+9le�(�%���c�*e�zMg�"!�
��W���f�]�x�0��^�%I�-�".!�L���0Y1�@D��U�O᣸�x�.���6�P��H/�jh�e.��,w�1�z!�"6��p摔H": �E�@�.��c�G�C�ח{�o��Ke��=��vJvٌ&��p��Pۨ���S2+�2QT�tf�ڹ��獩�ݜ���ld�?I��R�c!��5FnO'�ar��l�(`�'q��C����I_�;�����"*�jr���hrr>���&��kW!����攲Zw���ہ����z�́���ttE(x�t
�z�e.�t�VگI�O�<��k(M�>�V��Ѱ�,��R6�h��*����X������X� Gf��>)+#���s�cr�.r�*��^��aK�S��ׇ���2l'�����ѡ���d�(�9��aԙ݃o��i�Z9�\W�q�md@@59��{�Vp1���:��X̹8NtDbmT@�4��P	�k'e6�	�k�^�ׯ8�'Gn7w��.��މm7��!m9���m��cCޜ�9��9� ��I��˱z{Rˣ\*g����i	�zȼ�fh��EH׷\���-���W��0�Ŷw�[���Z�BJ��![�a�C�Q�W'�}��:�r��%�N\gRq��:�p�q����s�G�q�1ХJ�Um�Y]�E�1�U@�T����<7E���p�q��;�-�܂!H��G�����׸��ϣ�W���A���!\x����w#���V� �*H�pb�m��ji֧}��)�S�����/��.n��%jg"��]� ��V���bǰ]jأ������U-9���Yq��-Sntw@6Lp@��2�����b��X�kbvEf�#G� ��
44&�R��#��_!��p��ߠ�@�B��q('S����|�p�S���;�꾪L�Su����봎󑧬�?c0�-��Gr��*7JM7���yлJ�٦* ,�?LK똮�9ქ�\|졹	�q">���1&T����y~I�FD��;�+gV���ޣ8�ۛR	HW N�6�p�-�kj&�b�q�G5�S�s:��m���ԕ�z9{Y���E��wEp�ADۻJ�a�hgtV9=^〧}�9:�Y4*�z �v[ד%���oIݫD+��ݐ�
�lt�Y�۩��Vs8ͻS:��X�n�He���
�Nb��R=�/���8���x��-3��fފ�N��5* Ϋ��R{-�`믅�ɡ`�a�W�d.�r�L��ՙ����]ea¤�I��^��t��Y�'��ٿ���Rs%[-�s�M���'��R�]Eɼ���&�Z�߃7�������K3m;��V�4���/{�wl�)4_4�-;���)��d�bp}�����c5�j�� �(#����7\���iAf���;%�\��Q�Gme�9p( ���kj�Yoc��8
�4��0���������cNj^e�uN3*Rq%�.m���3��w5,�7����G��\��rvEz�r�vV.ӰW7�B�+��Ce����s��,Tta�q�q��"��a��8%�2��9����)�M�gD�sJ�.Z`5����j���d(��j�pٳ&���z6���
�.����I���	m���7"Ÿ���;[�]3�
ė&ֆ�z�@wN�Oi�4i�kϵ�7:B6�N]!΢v�Ҟ��i�]Ҽ�V���*�R�p�ne�ץmMrOGv�|��"M���e-x�V��]丹���
�]��n��+لʽ+��db�6Y��r�]���Q�m�o_`���~��ݒ���t�0`0�g+j�%�7$�lT�2=��^+��Y)�t�XǱ��⮟q얣 �,`��o>�e��ñ�pܬ�b�T����<��
�@+p��`&��`������(�y3%;�6����
��R����sbz���yMu����k�ӣM`a���/�'L�<�ʬwŌ��t&�{84Zѓ�޶��.Cg�h
�K���T's�����m^�/��ƍ��2F�R����	�79b���)K�β5�C
ɜb4�D�v���R���Rt���vW&�4Gc=!�z����=Ȼ,*\��a��ĠV����s���;m�q��ωF�{c��Ww�p22�j�[{��G�r�wV�v��N�fQR� �'M��ܙ�����Q�.�׊�m`䑬g�6l}w���ͼ�IY0tAv<��(��i�%o3,Yi��2ml���)���$�6��ʸ�q��-�3(p���p�f3�\��T�+!"��wʷq����&-��.�Dm!���� �̮5r��v-�!��d̼n��� E����M=F��<��P�w4�!C(q�Y",ol����ҍ�s4�x@����"����`!�0�;r���`�]��t�1u��mK���x�vN���Xem�wR�rQm3Z ���`=7���[���.�씵q�l��j��V�� 2��ě���(i��P���p�@�h�h���H^y�sw\��s�wp�\�\ہ\ ��4��)�Hq�莥������RE)��i7awSՆ�;#��p���P4��g.��B��y&����	Df�g�yVlw8��tND�aDW�듻�8ᧅN�I�����MJ�*�*��fB:����J�4f���V�5ayȳ�L�Y��E�.kN��'Zuku=ݗ��EDQ^���A��T�g�5<�qܒ]N�:�;�p�w1��z%AUE:��r��r+�L��YUw9MԹ�I%wwn7t����,��r��=����=�����8Q�%ćDI�Ys�r���x�y�J��D*�ng(�'.�W#���Y$�3���IE)de�9��ITgN�+B����I�)��p�(�HNTP\���z�$��G9r���A ����󣿹{�޽{����p���Â#4�3z��;��j�f־ɥ�.'x3o:�M�į&>[�+sV�+��k�b.�dT�a�Bl�2g6�~��0%����)� 9	$G,r(I�M��[.�����G�۷'&��>~���7�9G�\o
��ѽ��)��}v���.�i�I�'���0|���~|G��/��q{Vz������?���;rr�}ZM�	���ߏ�y1��ݪ޷�?���0��N7眻��W���9�ݼtbw���=��yNM���þ����oy`�� >�+�5s��__/��Q������0r��ݳ�� �9f�/���������o�N���{�SzBI�1�/���!����rמp���;I����y���¸u�a@�J =Юu��LP}�jr�{�y�N���rP���>����r�7ކ���XP�@CAz�>F��'>]�����xq8����~�7��P����/�nNM����~����4}�U�w0<�-�YMٺ�t���e�i,Ȇ��M����X-��o�ߐ�[���]�7��{�緤�]��߿�����L/���6QC�xC��~��}�];��=o߸=>ݽ'83�d}�?}4c�#%.��м�d��*������ߟ�{T��p)�L>����� }O�����;I���y}�rr�����7�'�~<�/����ף��>v��O�������6�F��}o��X�#��x{ݹc)�9�Y�����̥��,�� ���C�s��8����]��0��8�\�8�C����<&_��ې��Rw���C�|��7�'N׿��<8ߐ�(sU���>b"G� 8��9V��w������n�y���.X�h9h,Ȇ�-;���1�Ǖp.��='�<&�F��;��C��}Ǆ��;�'G�}C�aWrzC�!&��>���"+�iU^G�G�E4�{�{%	��ׯ�y����B>�DG�w1����rn}|vS����x����o����c��]��q�_��m�ܮ�O1ɿ;�M�������S<�9�҄} |��f<"��a��Dy_{��QؿGk���\��@|�!#�uO�>�.����n;rs���{xw����7�{��ޓ
��k�z���a�����J�ӷ����ӷ�������;rr�������F5������~��m~Pk��r�[�_����H�"+����:�^�T�܌�y�Su�}syԷ�@�T�[�-n�P�ݶ�T������Ҁ����WJYgk��
c�[{�f^�������m���uq��Ě����S)u\��m��e=�,�����>��1I����0���������.��������}��˿;]`���N��O����_v���r}O���?!�0��ރ��\{C�>]�	2�|v�Lo�~���C9OJ��^��<KY�g#ΰzvSuoh�<ts���o��=��:Cdk� �dDކn ,/��#�o��;��0����<o�x�������s�W3�e���u����[KY�`H�@yBM�	�n�����N���8�x��|~;rnBO=��oi�<��w�<��;x���N�� xK����ők,ȵ�'ɛ�9��T:������h������F����H���|�`x��ɿ�!�ߓ�aw����㟨ro:�@QC�|w��	���'��7�۷'!�wq�|�m�c?���P���̤_zCi�`a�xnhF}oJ��jהZ�� �>����OO�"�p��%��{>���o�O�nN�~��Ǆ܄�'��ǔ��1;ü�`��۟�����N���_~v�
}��{v���zb(|�!�H����0*���Y�P��6�y���8�r<7� r�������������߻x��L���w� '�;]�~��ޓ{Bt��X���rx�÷=�7�9�÷ }~�>"������"�����h)F
�j]{���r�KX4[��<C�0�^�e��xw�?;���xNL.�C��������7�$ߐ��ޣ~C�����ݏ(�8������ۅ|�Q�*��#>���b��v�wzn{4y���02���I��-e����x�:w�i��P�[{w;���f��ar�w�	�"�!�����NL/���>����s�C���o
"#�xd9��G�4��9�}��o�NS�o��|��}"$G�LDH���w�u!�0���Ѽ�ɇ׏���U��ӽ?�S�~v��'�{�I��>ݽ��ǔ������y����������P��#�Q�Å��Т�v�����$�Ar<Տ��"#l|��˼;]��o����5�����G�=�Ʌ=��ɼ?�?����]�`�/������= ~I��ʁ����7���j�s�jԏ%��+��/�eu	�6f�J�4��x�E�v[����G;N>�a���uzaq����/����}m\�<�+B\L��	ٲx���܆sPZK%ۜ:�I×1E�|�ރ����� LS�
��l�PT�zU�Tw!/�l��xn^j��mԋ Hovt$"���i��w�i�o>~���w�i;�yOI�Ǉ���97���?�y+�F'|C�$����]���N�����}�k� ��U_h�3��s?b���-�v7����G�mG�5�׏1����ɹ>~�	�~�{N�}��ސ�|_��Ǥ��n�o#�x�ӽ8�{�	��u��k�뼼��1�Zc�#�>��+���}�ᷕ3�������Ï����{ÿ�}Nq��9=�+�������=&���|����7?��;�]��۽�����zL*���?�|C�>>cӷ+���7ʪ�
b���}�'S&��0��dڙ���o�܄�8�G��7�y�/�o)�щ�w�>;y��?���q�;�F��=��w�iP<�Ͻ�7��s�;]߽p]�?8��������]�=��z~�"��@�b�O�¬vx��/
3+}��E��E� 9o�� _��<��w�
]onܛ��y��?S�w�ߞ�P�׾��=���ޝ����x��p�v�!��aO������~����~NC�y�W�^<ok c�z�c�jg�Z1���� � ���S��������8���+�	7��u���7�;��<?��}I޼Ǉ��ۜx�I�~[o>x=#Q��?���Ql,ȴy��n���e˾d�)R3�Y���	5�E���)�����7�<�(w�bw��z|8�|Nv���\rs�~�y0���{(�����Ǔ�s��b>���jܨ�@W��MU1�S�ۜ�UYW��x5��<6�k :o�x<Q�ە��z��(�}v�����SxB}���)�\
o�s>]�;��Ν����<' N��1#�>��� �����i �B2z�7`�"- 帳y�f�0E��,���7��]�>����$���9����~8�C��x1㠓/����x������G�<y��nM�>�;���kS@rf���ڃӞ������]@{�^���n}D!�">���c��]&��7�����_���I���@�}�u��.;��@��9�]�!�����'�߸
��	ǝ������dP�D�g !f^;�Ҷ��9�P�b���4 ʹ��5�0h����%�)@�0>����ۜ�뫧VV���;i��J}�#W:��+ј�ۣև9o�U4�ܫ�-^>V����rt�� ��q�N�f�3qv]gwt���p39��v�;��VA�ž�@�D'Wv8oQ�I3���S������yC�a_�<�~O	�	ǈ��o���]������GoΝ�~��ߐ�[};������w�����~B����w��_N9ߓ�wav����Hbs��R������׾B>vQ�}����|[��9���hzռ'��z
<|���&ώ�۵�7�9�O^�oc�+�;�����'�o^�}����ߐ�E�獼��� ��۠�庇�ɟm[kkѢ#�;rw�o�����]�������&;T}C��˹�T=|�ɾ��h.�1;�{q��q�7�yL.���yOh{C��v<+�&�n<'�߾=&�G�n?k�ή7bK������B}�"?�w����y�o.ܛֿ�xt�}�'���7�$������ݏ�<�Ӵ������<-�7��������ӓ����Ǩ���?;��4D���,_{��6po���=��\�����s�;��_���
������!�0:�Soz �(�fr ���	,`��>��ǔ90������'�ސ�{B�;xO���t�}Hv��<n�;P���(�u��d����,ġ�������>|B������}M���$F���?����{L\w�����uR5�+lh�O-r̠;��GKs�_ZB�6枎H�����4�]�9�P�(�:�cucx�[������+Υ:I��B����D��I�^�W^�
���"T�ň@t_+�db���R���~�ܭ�'լ�^��e	�>z'#���,x��~bU��(_�|���[go�;W�|lt��dΞ�-5���,��5�>�{�]��}o�=9kw����.��7����|�+ט+�$��\�w�Jلc|-oZ?.�;.�ܣl��-�̾���u7����Q	g�`�/*(��*_L~-�T����2�]uY�SL�W�o;mŲ-P륐�6���J7���)wU�k�i�7N���ҹR�r�ѻ:Q�V8-ڨN8�zt|µ�1q-S�����i}N��
���w�|��u�jN��WE8��c�ù��@HНJ���r|cD!�����m`���S�kx7���v�c ��	�'৑�����g����l���.+��#O\g�M=�����4������5(]�L�~f�*�5;��Nt`rڿ�;��z'�B�v=�Y]����ܐ����
`;��ҥ<�7R�A�U�Ѫ��	uK��;Zn
�q�N*y��n��"b�XD�6�@�x�$@��>��^dG�c�{ce���)�K��_ �զ�/�uM|����������"�E�������(�o���k9�.�4i��m��P�=�'����E}'�4m�@s�j�G@��i�Λ���XÇ��=:�w^���N{����^�Rʈ��ڒx�!>����@���l��vZ�R���,}ޝ�x��5�N�C�!'m��Ta�v4���A��_ܩ�FD.t�W|svU�g�Sj<�t�!� t��}GF^�r���t.�ej�<�������|���[^�];�,�#��,�-��ʴ�胼�ծ�@.�ޫ��WGd$C���-B.ǳ.�
���7
�K������mc�ᾮ<�!ϻ"��8�A|'�M��ڛ�8m!�ٟ��*a�%/:�q�1�]o7u8d���k��Ǹ˅���FFa��k�㶅�E���]���?�+X�'�Q��ռ�j�j慜�H��;��W�	\~sJ��.�{�KNEe}����IvEk����q"����ONk��nb9��P�yek���~PV��]pu�Z:�OӨBt��==[|���p&XWS<�/�BLbs��.�6X�7��V;w���8�i�5��ySF��y�X����H*��&B����r�(�t�(�N�����̇0�[��0�J$E�@��]��ө�N��ዒXV�bF�k���p�r��~�u�Gn\�eh�G��6y
�y|̧c��a��U���t�Ap�bҐ��[Tv��I���`ڕ䛘&��b{N�������~�Dc�7�>H�u�*=�Aؤ�.�|���C��r��9���?C_W'I�.pCg��o�mށnpA��=����w���f�=p`bPg�%My
�$e�Z�HĄ����Ô2vC�Y����˹\��l�g����-���,3y.��1@��]�/zt��v6��$g������y�w+�)��s1좯�A���c��e�U�Q&o�5��U�;
SӨ�݈)����s�tz��ŗ8�y�_)�H�s1=��÷�7.�4��\�Yc��H��a�ޕ��5:���2cc�vh�'1�3��΋�SU�,\�ю�=�I�E��;>FǴQ���X�ᮨ+���n�/jO]��y�l)C��mk\�Ry큉{u��[�KP��r�ߒ�HnX/v���%Q��u�׷l�1^�ʷ�����w�شLKE{��x��yՃ��4�TvЬ���3pwj�e4`�z���ft\f{�Q!�y�ݾ�2L���?-X7&܍������J�l����T�`*�q�VҋR��jS%������67�%b�Y#�e�Ft^)������e�^)ؕW[~�a;�fA�O��.g��=j\_�]xS�˙`�;��d��b�N�����gc��m�f��b��AFd�fOkK��P�TY]XY]|}j!	��q���O`�糆�����f�F>9�5Q��QQ�iHn�cº�uخB{�]�N׸�A�E�>��|�_T�=�[[���>�K�Ω�7SW��2z�2ST��Y�!�9���2����l���[ݾR��"F�ɖ��9�7W�s"��g<29S���(�jL���y2����9Gg7�D�qxfa�����^)����Wm�յ�ˢa���[���ntu��ƣ�$�~���¯��G���c��<ĭ^2�q#���(�=��Ի;�s��m����lho%�h,����< �x�V ����z���QB��z�1U��I��%����1�q�"5��摔H"e�l�� EhsUW�$�4Y�����_S��\2�:8&R�_�k>&��p���n�rΨ�ǚ��'��nS�����K'�D��P�BF{������
Xw�|~ʈ���[VX��eu2��ue�/E�)��Ր��uP�#��J��)��#�Ⱥ�]+��w�\�2al`S��LnV;�8�k��mt�[Ӥ����JuD�N�!h��G#)Ez�4�j�Շ��v���<�b�8���A55Ed+�健�sCC�𘎖OP?-4rls�=��iƅ�l��w�����L�u)��Q��'w�!s���P��on��{3��:mi�vJ�ښ&�P�(�C��3�e�9��o'��5�~�+�)?z+Y[�Wq={Q�M��,��wZ�YJ7���,R�]w���L��P�A)͗W���/~Zfn���X�WEm�^V��@��!����s��r�{l7�-哰�m�O��ǧ��r��N�i?A'��.�f�T����ں�'Yp���j��s�f.�fq�.w�T}_�aU��,��p��:Le�ᓁ�NQ���d���H
�ƲϝS�b9��er��e�8m*=$r�;S��*��ƴ�q�3U�|+��n��e��1]vj��<��\�K�^t�+<p��lw}~�2�SO܆��]�'�7�$c>�4�Y�P��vn��GiY�n���T�E.C2��q���Q�Ss�򘎿�W_�t=��NZ��@�hd?��02�S�m�9^�(}���.���qt�柘Yc�l�ĵLnNV��@��%��G�/���'��y��c�Aۭ��\j�ń�{���T��94BO:��m���Ɨ^�NM<��כ�
��aE�J��S�I�/��2��x�x`�z�#��i�v�/^b�N�Oˊ��,�t;� �
b�������DTF'\4d���ٖ瓶d� @T9٧�z��d���ؖ�@zX��3�@��A�
�9����q�P���}�*pe��ܨ����u���Dņ,"i�Z�Q;1?wGQ
�k�*b�-Q�Kۻcy]Cd�Ӎ�U���:�M�+�d�GIU4���N�f�B=�}S]�p�f��<��5�8`��c�G��j�t�����U\\��7�����38Xzz8Ov��K��U��2��r��ۃ#��-���1U�م���ը~���;*m�/�^#�y��c*���&�x0�F,	UJL�J'�&F��75�~녡i��]sHm���!BCg(���7���m��Q'�4nt<����b�2��q�����d�5-$Q�e����*{����b��Zj5^\,Iݣ��Jy*���=¹)���$'oɸ3ak�hwWk�W�Q�	�
�<8*:�i1n��h`b�S쇷��s�.����b~׽hS�g��tN��"Pz8��?x�lW,5�}n�u�� H��0i�c��=</U`�+N��ތ�$v��}N�Q0�qjUV��wg�Qw�C����:9�)z�=�=mv v�Y��'����5\"�k+�1�)���N˔��<��\�J����pQ����;!.\��S/����[��s�B�:nN�?Ŗ_�<�hN�����h�	p�L���Г���K��X�)��(v��2�%֞2�ꄥ}��ۺ=G�,k+�/���J9���>T�����k�Hc�衔�r��U���62rf�F��� �7�S��;V��km_C�P���؎�V�R��� ��8BQ�t��6%&�F9�K���#r���@�`L�2���[N#���uU��j�;���-K�; �g@�����4̻�H}vZ��[z:�r�d5���`i�����6wr�ś�F�(5��m�Bu7ц��ʈul��q4���qsD���rt��"��T�j�6�*�*�X� R���#�v����Z��-��|s=H2���\^������'tĜ`ꕓnɆ=��C:��ꖖ�������>w���Κ�"�.K3~��ah�+#z�v82���w>g0훏�,��� �0�&��7�k�ojmcpK���U4;RI�S��+��c5��t/7N�%���J��Ip2���ϝ[�yf����ӕ{�V��B;k~gq��-�����ݫh�aL�l���tJ�E�Dw^s=ٛĢFk�TRQ{���%=j�wVh�IA�b��e#FtJ��8��GK�B�I��xT�bԻJ��J�r�;�b�1�gf�DUF]*���R�|����vTy��wj�X��j�dW��#�P�K�
��ۯ�_!Ǐj��xR�0��W�+��ґ�/jJ5bͨ*r����gY�Zk-Ԩa���(�g�h��'�h��3����B�����k5�֫Qu��"�^ښct�,uҮ���m�L+���=�
�xf�ͻ�漩�htJU�=IӮ�Eu^��ّp�1�;�-o���D@ܤ�p�ׯ8�Q�m���ru P��� Y��6��X��g���9U�16��2�Ft����"F$퓑�q`�oӘ�*�I�;.��[7�rU�Z�ѕ�{��WhK�%�TC�C��Vr��k�r��|�if��e>�)d�iRL��a\�ە�"��'u�Q&o�3ap}�QX��p�S�|Wl;��4,��8�(��6�]mM�)!E�-h�3V2�c�-�}*��_o}�����=�^V<ٗ[�j��_��u��v�9�wtz�+R�l\h�+�!;P���خk0�N����X"�nj��6��ث���%�I���v��Ԯc�3��(ј�h���n�%2�������Q�#2����26�(��9]�`0� ��P.rv�f'xe-�6��cFWiR��`5�Wv"�v`*�Vۤ)���_ �Er�i=�dW���t>7��Yv)4�ͦ���DT`X:��K���wk]ݤco&�m.���R�����S����T������� ��}��m)��m9(�9�wq
�闅V�%�^3����4c@�誱�J�|�}`��L�5��I�\�U���jW.�Hl흶h��
��+��Kx�'t"z��Xݨ뮆�Q�������{��L�V��K<O���jQq ��+Z�Bq�w
���B�!9QP\"+��d�R�E)GbTA��I�;���I)����#��riܹ�TQBV��A
�Zy��z�"pJ��wK��*/2.XWՅ��\rT(*��t�&R�^WC��t葐�gvU�qJwh���I�C��+e���<���9��
4OR��9bS�����r��$��ԣ�Me���g��e�=���Ĳ�H���=��H��\�{�:��\܌B�"T�����y���/Q��3B5�rJ�B���vQ�g�9z;��,�M"5��甴��!�aS�x��V;�ud�E�^�%4"+1��Id�K��7R�N��J�r֔�wq��D�"��
"�)}D�
v�1C��u�]g�t����{9���^�Uڜ��K!WD�ζ��۰!�U��+���˼UU�&��}Gak?������9+�;n�����a�g�B8OI�2��! x�C>r�[��� ��mI��FŻIE�;nw�?��ö�85
�B�.�C��h.�v-)	���.:�wf�!Vl������]q%��]�C�]�&���#<���O�@i|�ľ�۵��q�\�)GJ\��m���e�/��3���"���l۽��3
d���r�!D��IoMt^�ۧ%pH3�!��������bB��:=	�p�. ��K�k �1�k�%<�oԊj�d�T�/�M`&��G���W�τ�W�v��$=�P4i�4��Ș��V���r��p��O��1S,*��)���c���`��5������Z*n�/
,��_]��b���8��?����i9`I�l}�kʐt�z�TN�!����u�ng�>�QsK�u�j���Pn��ٹ���1]\��K�yS��X8��lO���In�(λ��xU��0h
[�N���En�[zM5LCE�������]>fϝd���|�G,�P�Ky����Z����W/��W
�9��&�݊������{�S0�ޙsfV�P����h7|�ڧ�U��ꗶ�t��V 3bk{`5y�rQ}�)N8��Ks�tǔ9�:}$�5d�[�[2��U�# ��B>��֚F���yy#s�Gy'���}�W^�*A�zR�
_NLTE�P��j��ps�GV����B�$��΋��:�Bj��Q�lfww�1��7�KF?�_:��G�TNF̠�����S,�<n����:Α���}:cS�W�������W�H��l���K�c��<v�!���p��������qTy����y���w\����F����QQ�iHn�c»��P�F�o��G@�yjg9X�q�+њ�a���;}��K^�KZ��N��D��������g��^#�J�e�K7Ei��G���WO".!�^L孨O�� 3O,Ӻ��,����>@p�b*���V7�DRj�ne��e�1�r�#j;���37{c_��S�4�<Mv�Ez���2����ǅgÆB���q����:h���N��D}mrB�y��w;�S���A�G���"���G>�Ja��(&_���[by[����x�q��ǀ� ��g�{;(�@���C:��!��:�[�=c��fYx�3H�ܤ2�|Ĕ�X��C9�t^h�P��R$���~�=]��wj�e�k9�wS�΄�(���b��ML�k�TD7ӣE`ۖ�q��#́�P&dd�V�l4U>Sn�`3���p]�M�!b�;.��aE�d	�?ĜV��#��>�{�}*_��ܑC�Ω�%,���9,N���(��d-7�yQQ��k��	��D���ĸ�wۉ�ؐ�z��=om�mUѿ�2��4�.hl��?t�z������cfxS"f҄jg�끹UY��oǲ���b�Vλ7�̈́ �w6i�H[@==��Z|�<�:p��C{ቺ�q���J���\\촅�:Ж�Y��^��,�'B�zr�x�f���CasRT���
�8�i��z��_�'.#:���C��ح�B�H(���=T��O�s\�-�`�����!0!�B����q� ��@j�midc����Z<ڌ�Zd8V��.%�gs�u�i�o+������F~��W�cs���.*���K��o�0M˭��d�����1�x1�n�K��m�Τ�#���_�޾̎�y�BT�������n�R�#�Q[�#h]j��qYc�l�ĵLi���(����'4�ڒ��wo�%y+P��[K�x\�E�F�֥o�2����n8.�}��D�|�y�h�����R���WmY**��wl��[Ow]��#jDhvc5�o�I]���_.L�w�З�wp��Kᶝ�*bY���JQ���v˽���
�scVy��m�lD�:i	��:� ;/�7�ݵ���|����<������}���g��˲�~��_( pC���#�G��I�n~!��mN��������[��N~����Fi�W*�\�4x�D	@y]������
tF'<0S�3U�䘖$��W��E�ߘ�����=��N��,�0�T"�sI�<�9��P{z?,e��qÛ�Ե1i����ڤźD��b�J;�,����d۪�8b9(��z^�z�M��.+%�ל��+�h�e�UMD&�x0�F,	UJL��(��������z��ޝPf�������v��J�|�_ͩ��y�F�t�W�cV�;q���_��%��;���U0���/�fߨ���΋}{Բ�[ɪ�]�K�:������J�	
�f�ۥQ���ʼ��F���v�EI�`�k�p9|������Z����L2x4�il,�`�)�r�^~7O3�s���Z��p��~�[b��h�P�r(���{����թA\ q˪�FY�e9�a}MӚ���ʺ�{O 	mPʜ�?t�ײ?e�8����C15X�n���w�uսg��V��ڽo�>Rҋ;n��p=�������b3�c�Δ�{V�ޡ.�A�gJ�x���uy$G�\y:]>o�f���,EB|���q��-���DV��1K�l��d=�5qdԙ����`�vn�3��B��j[�G /�Q.a�[��t�Bj�E�Y\&��Ё��Zd����Z:gp���pOp.c"5NK�ڭ.p%˒�����k�xK��
ݿ���K+��H5(/96��{�Dtz�"M������i{�/�P����C�+���Q����t3��>������
,e@���A�(xW���.Z<e>T�oz�>oE����U�I�"��랥�z��dvRz���$��.VbF��뮠�H�K�*�)���J�3�[2��=:0_,��f�v�s*aE�����~)V��-V䇖d��2o7���[�_!X�\M�Kw,���w��u�TF:�|�'P�8���Y��y��"���s�p�H(8�#8��?o'I��6s���`��2{g���99U*��e��"d>-z(�
j.�F苼tBj綝F4B�d�Փ]�nq븫�v�o_Պi ��ED;�:h��;�X*%L1"��,v���Zu9��9�Rb4�c2���K_�NU"�>;�)C��"6#C� �muoU�����
f��z(�M+3p��yv�K�bIЄ�Qq���7��Ά� t� �q7:�@a�כ�1�H՘��,�GX��SA%��m�Kw��m�DkWg{�p1p�����]�&5��nŊ�U�}�W���&w��.�P�x�^H�����SbԲ�k��U�Y��o*��T�֮���ױs���Î�wB�`)��NXj9��+}��x�����_�n����.�O,8kR�Y��ƍ����+%��T�Z�A���E���:jdF����d���f5���p�f%r5�u.7�0FΔ��u0�IjX�����z���8:0EN��P�:/��SP�oL9T�2W(꣏.��(|�P���뇟*�L�dF#��j��6�s�2d��ӹ��������Y���+T�9t��~�T����z,Ը���r��+��Qm�F�R1r�NF^��ue�)-�5AZ��@�׮�#%�����z���7�C�n#��V���i<�U�ɨ՟�<!�-��w\�3|c���l����*����JC~�_N{�\M�wz{y�M	�Wu؇�S��8�R:��n�n�,��r@2�6-Ik���Sޒ�ǎ�S}��Y��{�q�ެ��2���Mv:�6s�B��<�e�����b �oJ��ti�u�nj;*�'.�x��4��3�~�i�<�Zu�ni�%���HU�_D��@R��������t��-�o��
(sb�t��h�|
t�7[�k��>�e�b-��x:��jQ<5lu7�`ʆ�8�h���	�U�ٝ�����ﾎ-�J�ikG���8�2a����#X�2���2�q�.a���"3����9�z��8	o>Դ�ɐDJ�U艔��_����5�.��D�m��oJE����e�����@�d~�e���P��\H�� l�G>�j���
Xw��%���	w�v���h�Hhpy�,������Uϝ'
�v�U=aL4F�"�\b`IU���p��q�˙ܶ��4�]r��?kJ�-��֨���"8"sA���s�*�D�n'l��R�q�����\�7�p�Tj{lcj���d,/����OK'����jk<��r�����k=��+&R�K�u�'w�!s�E����
�V�x�^;��#�t���-�V
�3��~�+=mE� ��H{�T���8״R���ExD����Y���J�y��B1`��ɋ�ᓁ]NQ���d��R��bS�@�;�0n*:ݤ����������:�S�*���_p����"*�k�TћH��OX��:��.�ԑ��f��g~A��K��l���=�i��vf�擬û��>�p7���b��R�sGH���Is[��T�v�K��k�S'�;��m=�|e�<{�+���Ӫ�L�e�	��I�z�1@�����_}_}�oMPe!i�������r鳸���-��͹�=e�������t��j�ݦ&e��<_�j���d![$V)M�o�)��3��Su��R6�.t����{˱�KN'��n��7��������Ơh��Į�pr������f.%�cs蜭���m�[}�#M�[���H�i�ID�.uB��eb��(��	�J��r|cD!���5E�*H�yh��=�4�N��M���g� ����O36
G��̷?��%��ZmP�l*s��'c��#������ۘB
��GA��2�����b�������׃���גo�UXA�%Xw�����q7��q:n K?.48�E�T�IO8�j�tV���$�����ąoMFv��0o&� ܢa|����u�[�q"1�>H�9�M˕~v����b��[�����Q��UM&�p�0!�T�ɖ��74�$��'��5�����
9��oJ���}ͪ��y�F�m��Ԡ�x��D�Ŏ��:jr���.ݤ�tۊ�,��n�U�nQ�~�ZPֲ����7Y�3�K|�*�N.���r]!(zs)n�f�wE��/�g`v%'��	���V]D��f�ݗ��[��^=��E����y����Ѽ�2�$'ˀ���r�K?�4�q��=[��*|�N��<2�B+�ŇQS�~8���0���W�whQf!��8�{kz���V��<�%^%]�P��
PU�5h�EVi�]y�n(P�d�y3�E��2�0Wt�㣆������\�#W�k�+ʜ6u*�d��
�C]�p�&��fE��vs���BAO���c��u���VצHw���x��ݧ��eN�&'�������ubJ.��91���"{$� ���E���%��l�&��5só�"�� ���α���9�������	��GDj���M��;)r�f���k�\�MǞ�ޫH����Z��Vsj5�u/Ԧne u/��ͣ��c�H������`�*Έ��@�yXM�5��n�ꩾߖ�
(;WA�|�:�P>���Ϯc<W@�\�J�ej֒�]��:��`#�wl��d�ɡ���rK!��.
�H�P�����UR߄Ӡs�j&�
q]��EĹc�<��f�v����*�p-,}^���d�f�x��\��q���RdT}MN�aãfUq&���U�S�]Aҭ��&c:'UE���v˕(�M^8��M21k{Qy��<���j�l����%_--^�F�r��L���ڲ��x�&��^Z��IG�V;�<�q�yv�+{x�VK�U�}�|]w+�D�t���
pG\~�>�ފ��-�p��Nti*��ꐚ�2T��l:J����zں Y���ڤ���+H|{������6r��o�����Y�2��ǧ��ė^p���ؤ({�)Q�XD>>�c�zx����[�p��b,���y�c.��;�}j������<���
��3�G��U���>M^��w�����GI	�is{I�f��0��]f��s�ѡB�Jt���;\�P�}�e�c�__n-�3<�X:��<� ��뿐�n�S)���8>�s ��'�d���~V.��nƍ�҈źԎ�/nxB��cY,r�b9ַQ`�lĎ���Q9�*��������и�:��D��;:S;��C�j�!��]D�����3�o�m	�T���v�5��U!�ʅ�G�EDZ�P��j������˒r+Uܑ�ds4�sp{�����[K��)���:k����c	}	�80�c�i<`U���gI=�6�����M����g9R�a������|��|a&��E���S��kj3����Օ}���M6 FZغ���J����%���"�43B:���b��'�u��1S�}���ܘ<�`��� S�Chu�V��Hj����m�iWwL�v
v*,c�pRWE���DN���XNI0�qSvjH��n��0}��)oZ�!�3��\ì��7Y@��������4&�����.�q̬�����zx��\#�$:}@U��*P��F��I�\��FX�5c*����m'b�%G�%���L����hc�x�ݖ#ۂ�ھm%���v�Jܲs��4/�4+1�j��4��5�3�+Xܾ�ҟ���s	�׻j!9]�G����X.����֫����s��h�6�䮷����VV'g�;��m|
OAҳ���_8�I�e;n�l[B��8�=����~�ͧN��miwyI�^�:Ս2ܢ���{T�4ق46[NU��oh���L˝L�f,fe��cH`�T&��_�r�ZV�+�j�N�T�3N���:s�c�Ч�WnZ��f��u��v�}HˎZ+��I`.H3�y"3{�Om_gjR���m���`.츳e7 ��'o,,O�2[֝�z����h`0Vnh*�Vn�O��+�x-t;D��bx8�{��.�VvS#��!K�nQ��#�!���-�j��v��>�Lܴ0ݫI\R��Y�<�{�o#��VQ�.��Ү�;���(�+���|��p)��K=V�K�5�[���ѩW��OqM��g�59�2�U�|���]mL����%2��U�6�w�CC7s^<�B�z�ו�S�0��c7R�F�
���󾩘UJ���#)#�����8µ��5[Bb�D)j�Y�0+�o�5�E!���D),\�8U�z����+Y,� �gT�:B��"䲻�Cs�KV�o��k��kΉ}���N��tlo�[F���t�J�8s�� v^]]�u�JWb�f�;�E���Ջ�R��8�Wu��#��:�[�!"q_tF�m�WQ��.�埧54R5���bRu���^��OY��,ծN��_G��<�Fm!��e`�h�;�7f����D���sU�dƝ��JY���a7GHz����ښE�[�L˜U ����Ki��A�7r�aM������n�����[���]GL$j�x8ņ��rK-)�����!쾡6�s��Jkp��mΝ��%qaY�XŰ"�x��s17r}������Č[k���I�v�ր[��w��os}vkz�o�G�F�9����ɛ</k:P.��%��:��&(>�L� ����x5��@�鳋��xڗ$}>��>�G]�̜-�uz�F�r!��|�����;��ӄI۝��.��h��#Z~��WH>��k��)g���nڑ�a�����AA REx��*��wp؅yG������b���Va��=ȒQ/	�9ē,T7]�$�a�'���jHP��:#��ia�s"�wS��v�"u,*��]�tw͎�$9J���jJ�i��rVU���䢩�]J13\�EUR�HEI(�S���t��I:���,�R���&����
S.De%SR��b�{����i������+D+tYz��t�tI)C-1K@�M�d�X�Z�&�]<�8F�b���if�t�c�bR%C*�Y����wh^͑�����j�^��tMfQ�t����FQ,戦�Z�#���"����2�$N�&'��ڑF�u;���f��J.�t<٨�S�)�{��TU*��R�.��*t�T25��xu�i8�'tCIu*�y���T��*hJ�� �$G]Aе�<"Ni�
'D�j�f�eY�T�$�--D�N�.j^xR�'�sD;�H�(����[-B:�;9J�{���!���w�P���4-Y;`�b���ǧV��ee%0t5w]�ޒ��iL+���_W�}Uꞔ�����٣�R� w�Wr���ja�t݉e�� ���"��V����(�9�8����=Zu��C\i��
�������>Ϩ���tƸ�Y�+G��eG�G-)�|(���P�sk��4��J�B�-ތ�\L!��=��w��h��'�GIHe]��9NyLwv���!�C�6��'�YYS!�9�Man�R��s�\����g-LϤ!;��k��u�F����8��@�Qx	����hH��X�2������˘c��rn�e�o�F;�۾w[r�SL�$�G�TDĥ_
���B2Ʊup�N�!Ԯ�ٷ�)Hp��W�ϗJ�Ub�]�t�������\��j!R3�1��xd����U���6h�`~NV��l=��{8t���\���[<���s��\��J���
a�H��.�k�z<�Na�#/9j��K�ήZ�(���攲Z�e��>�# ������	
,R���B��y�[(%��R�=[�F���Cj���d*�����5W�Z�NP�J�W7��Qt&Ӹ0���]NU��
]A|�p�YG��+��6s� Uj���`t�}ץFi>`�+2�s8��&kz�uY�{fZ+T�$���W�Q�'&8г���o0-@��k�wҜY�qGBXR�7�'SޔhO���y{G`��&d$���� ��s�,�Y��w�1M��*y=1�v�譗ţ��Ɗ���q��\�F���t�jwrk:��HG�H��"7�"%�]u.���l��Eg����H;��6����.j3�M�Cʋ�F�d��"�gṅɸkH��KZ��i�4�:��j�>&�> j��f�y1lE�{D�V�5ֳ�t ��㶛�PT��֛�4c���W�ବ(G���A�o��O: �}~��DS��%Iϕ�٦���{�S��R�3����s��V�x�t�MD���j�K>�T��;�R��ה�u�:�n|�o�=9jP�z��C���r)}�'\ζ���b�g�Z��fF����u!��wx׼*VzZa�5
=��U����iB�6L �'r&XT+��a�����5��9�2��T��އ0bg#�u�x"G?��� S+A�x�����%��XP9��ȍ�B;����A�UӼ$�-[$��۶�ǟ��zʹ5G8�6�Z�s-���������FCu�#M7q4�fh�n_F]��ˮ��g���V�]p�>g��3����!�ץ�UųO�ެV,r�s `�s�"���sZ�ჩ���xmқ3%��d�N��ZZZ��gd!�Rx��Q#h69�XzN�՝GB��}���ѫ�HU�)�GwN�����:�C9:�&޻��p%���q5W���P���CW����h��q�E�[0�܆j1_�j�#Erj�Ȃ�"b�4ۭۨ�0Y�v�ɜ�y�˚��-���-~���{�}�'��b��Q��C�I��^@t�.!�.t.��"GD�SA�>����1 6n�����!<q�غ�ޗ���s�d�&�=��������-F7�i�;ilm�$����0�<�����s�*omN������&���}
b����BU��yj
h,(*��k��1�Q��Du��`͂=ە�+���
��He��?>����9^g��;V�<,m��?xՆ�um+�}��<���̐S\��D�W��0���k�PV�G����~�/X��i��*X�x�|)���EGa��X�/q3 W:YQ�׼N}���[Sл�M�s����KN�1��m����!:/�%�]��o��KU^�z��+%�O"�z����g�v�n��Μ��͍��✟p�(�0z�^J֨���u'VfY���4�K�[��]v/\�%�؁�_EP���:qe�L�V���}�Ru.�حU��=�/��R����+z� �sw�.��!8	C8*;S"T�[遞崁2�PۛT�f`�x��9��Eg��#�
ǗZ.�Q&�0y��u��\�au���^�L,��Yk*o�D�;����F�y��N�}�b����E) �@L� Ҏ�i����˂0e�{vq�L�o_�T:C1�u�P���?T
����,+I��%��_&���.!���U±�;�}��1�ˡ���X:�V�D/��ۗC��t@��Z����j:����}W�+�O�&廎]���p�o�e:�$O�՜���̇��<zt ��̧Z��\^�"��.�����f�$_��`6�#��juOilhn��:e�t=S0ѯ�@�.�~0S�C�v�]�u�Yϩќ8��!�����m�d`��Ԯ3��+�C��GK)T�Џ\���1�Ҵ��u�Uz�/eC���-��o��ҡN�} j�B߰���c�j�]�4�tu�-`�Z�{Ճ.1{�\�R6�6�]��ZN��>�u�^<�|���/W����T
�.Q��{����R�wr�L\�s)<Vr�w8�Q�3�$B��Y�Vй{�9���y��ڂo4���搧F�{+��C�谜���:��H�k�9뀁E���'i�r��O*9Bu���%�������ci14J��33 "��,�5�.�7�����=ﻭ����b�Sq]j����3j�D%�]��n�-��W|[|��u�(-#va�VSF���Q�)���a}&C�n�!��]D�ej�7�$h������Sk���v=�0E�`ـ=F�/=����,���j�n�Nv@��x�^ c�3�ch��a�jK��wR���e�sb�K�ΩRZd$�n�
�ho�:�d��������kX�B�ڌ��7%q`�l�A�1�7z�^�K��R����ixV>�r���짏pdZ�r$�G�q��
������Ko?r�1���y� nT>�������ଘp�6�a\i�-���L�7F�WI]�Y��ё�&�{Dv�y}���ֈ��K�w���Ә��+��ҡ%�����Oܲ��C�l�PR��9�f6��M�ީQ��AV�b!I@�Sΐ	$|���X i��v�T�#E�	x����D��c��Asv��
@�w)b�x��y�0���f�|��R�D1��s�V���S��!y����IvE�c7-���Z��9�@״~G,Me2�����GeӇP���(YQf	y[Nq��5�b4Z�@:k�s\2E�n�bu�.ҽz�����p���H��[�ء�j�*���b����]�l���aQ�'c�L�%9�>�>�"E�G[��Z��	�W�˜Q;�԰�Nu%����H���[z�8-�S�x�Ha8+��_s�a ڢ�\O8f��UΓ�W#�T��2�.���ߨy��;�^�sdT��\�bo�T��j�1a�O�)d���Q�JuD�D�Z���=���2_�N��ߪ�����<�ҷV�jz�U5��c�g!n����~Q��g��zgE�_��nU�2���gE��Ļ5�<^���eM����بQ�޽;3�1mW�a��:-�@�U6�h͍��'�u4�4o7��jk#~��/N�̄~�r?C�J��D�_t5��j���@<(��c�I�4��RPU����M��oCu�z���9\�`Up�1�o*���{ZK�' ]Y,m{�~v^9/rH��_-���z�����ou�[�(���\,j��ډ�[*�2����Q�7��s�:�fBة�)9ەSc��s�^��!`ŤD�����̙5�ծ���p�	$�����0��5�����@0+
�2�����[����X��CS��N����ӥ��[q��Ӿ��x�����4V��5�[�l���޾�ASNtS���rn�b�x:�M�30`oN�C��w=;��]��)�a��3U�UΓ#C��p�_������\pB�����N�uCVm�v�}�&	=�Y�rB
��sr\;��yiӖ��D�ow���js�̚�}誏Q$����E�X�6�;jN���ԦU����5ٮ3j3��CVne?�υz�W̞�5˷m�6)%���>����-��gB{���8�8�]�GkN�d����M�+5�:�Oky�#��qڎM(o�A��o"���-K�U��oi�����V�@@��s_O.ڽ��Z9P�9��a�ǥ;�)c6Mͩ�X�k�5��V�Ll�
q��"�5��f�S���̿n�[��z�Rda\T�u�>���l�|���Z�ʿ/eQ��}���wIQ�z�[9Jn>��3�eo[Z��k�/ߛʨ׆�X�B�1��{0-�&�����IV�p���P��Z��Cό�(s�@"�ȶj^t"�u�6�3�ו�K^F]hof���J��زZu��^Z�Ku^�RV����y��{`�M�/�ng'a%-�B��׽���otL�\���.	3�G�#����f]�k9���#��.�R��}���!{�:ܬ|��Z��}GkUB�7_b�y��G�X��M����O.}������<�s�~k�ʸ�m���з�[�g��RE�kqg%'&&��x�c)�ITM�T	Lu�˅Dt���u��5�c"L�n!u�ج��Fߖ3�hY-�	������#iCW������e���L�U��G���/�R--�:��F��YA��M��iB��2u���*��]�y�OOrQ��7cV&޹�q�����%A�>U{�����v�o����~Q4���kOn5�Yp�-�m=��(w0;
�v/j�]���+y���]t�:�KM��O������1�d��±S
�&�"�Z����n��mf|v'�7�
��OtT<g.mm��y�;��y�o�����+�R0R�CW<�G:�q�M$�srb��rp:�ϯ���w��/8�_'����yV���Fk@e��\�q�J��d]�s��^1�"2%l*jR�b~���,��-�ˍ9D=�y�v9r���,e���Y����h�]�H�t;���)�s�vMӫT#�a=+�lh�"��A�lD�U?� tw,=.�ׇ�{;r)[3�!OJUA�3�c�.�<{�r���bb܎�'pk^�mt�v�l��(tu#�9�R{i�X��c�'+�1�ڧ���V�I�MsLJn1�#���������g��n!��^�n��C�\��_��-�ם���ic�4����r5��0;�*��g�K��}��ӫ/<2F���-}��nV>E�-p��Ʋ����8CK~o��������^ݶmN��~+ҢV���r���K�m=jQuُ;�]c��8����)��m:f����T�t'�LuS��7w�+۷7kʝEɿc���ޜ�?&x���}�MϬ&k=�BW�Y��⡄���3�d����ק�TsM�-�B�ݶ�gQ݊c���7>���odtL��u�9w��e9��z��B��v&ި�\�N�m���އ��ފ�T�i�5x�� �t\�j�/
��먠���4�s
��5��+&3�{LBb�mu�0C�'JK�gz�0EX���s[f�*����51��¶;�ިa��rʼp�U\����t�sEd�i�-{F[˴�ʊ=��\P�W�_UQK܉��`g��3����)*Z��cб���hjf;��v�h֢g6��ry��<�:J��\��㮋�KHI��8kn�����g�/J'd�&�'�g��nc�}0T�LPԕ���}�`��r�#��@�:߱�[Fw��A.濛����֧�u�e����M��MP�sr\(���J����qޥ�l6�2�"��y���Xr�k��FKͮ"r/Ws2��5*��\Ն�;�V���*G�;��\�o)Y( ��-o�%0�Qf�<W��y�?zOpˍv�D�d-��9������9]��B���c�~���erٸ�յ����B�
i7���ٰ,�*�S�蜃3�r�y���ʽj���=�:/&�Eq��͸�����=�V�g�\f-�DO��4�K��|���7�Y�֥=*�)�2�ׯ�ýs14��=ؔ�B�Nƻ�<�Cj�Z����:`�'���*MK���xCwlW�?E��J��ES���EP�z�Y��LM06�7��͍�Z�Ֆ����o��+L��6�j�ra�:�M�=RvS'(��B��L��)�*�"�;k{���q!HRF���P8û'A7F�ݮ��5�X�%���zU�9��U�B�q������u����Vʜ�C^r�C�1B���Q]����TP�+5� Z�)]�<�^����+YtI����E�X�V�bVZ�Q�1t�koMݛ9CM.}g�l��NeLp����]�^cTq��h��w����.�������v����jQ1@ig�v�.]#�Œ�^��)�'q[ig
�WY}(t�xB�b��C��8�Nf��;@���oB-{�= p�;F��J�T��C����y�e�H�oGQj�t۶�V���@|$Y(D�P�0�'x��8e�'�1ׂww\�����k5j�LD��Bw�:�ټ��vQɱ�v�e�)����WD��|u�YRo��Z��޾��4�˒�zhǰFb�w�y�NNo6�61n�rP_^��*fM�JU�]�tMŭ)K�
ۙH������z~��nm;T�w$���`W9Gv��1�v�T��Ł�)��5pl�˥Yl���M;LcT���_<��6ڇ����Ø���:)K�_��ϳYrژ��P�ln�]�Gt�hX�{:?��pck!���2룊������KN�/mA&)�kC����w�����7hM�s�Nᙹ�����e��Sc�H>c(�K�վv��֊5�I-�e(���f����$5��粭3�ۛK�Z��4 nc�R�Ҭ��\ť���A]
�]h
�xP;�>�b"ո����^XAb8�&w!����l)l�����Q��*�]�-5��k�cF�Df��a�AZ���-}���uoV)H\3.u��י�Ġ
��'0���/�.����*�Xզg�ǯD�uq��zL��&�X���� �ՕG�V<
�2n�U���6CVcC7�S3o���Z|)U�T���K��� �(�aG
c��tI�nR�eJ��a�4GGjr+w���.������E;��3�`�� �t�G�fT]�ٻ�������}�(�R7�ˉ��������5{�lVh�z6YtE��r�������8P���B9W���Ssl�G~s -���h��]n�Qu</���2�E�����Y���Mq�ef�̅����v�9���K�Y�R�K�4�>p���g]Ih����s�iܣr�R-��d�*M�R��l�=��$.*:��a�$�����C�r�>F1�3����L�������W�����onⅽ{��d����A���|Q�Mң�mC��w�:�}�b����O��ʧ���W��!����u]Ҏ��=ܠ�R�%:(D�H%t��]�9DGC,�8��䔹;��K.���by�:,�
�L,��MU
�U�R�RL�f� �������
ĸ���T��KT6�;����VBeI�%[u=�55͞,�S)�q5f��J���\�����:;t���j]XV�#��/T��4SB��FJUHHZs,�B�Q�7%ى$���ջ9�e�*Y�
�T�T�L��f̭iY$r,6f�ΙI�,B�u�31�<H��S�p��R��jF���d����ZT�Pr��-3�ЉIܜ�Y��%DbmȢȵ���jb�����ք�&r:r����"�VF�$�e��2N(V�B&Zde�(��ܽ�mLᴤ�HI���i�,9TU�B��TYF
��bQ��HUL�J+J.Jn�l�Q;�����姓�JF�Z��E6�f&E�'��!)�T���)$�@�� �D,N�ȧ�Ym(��ZY9������f�ʎ���H�K��Zź���w��X��J��:㚞�� .������}UU��S��B�5���N��'�C�;��M}iu�o��-y�U:j [$����{_1�Bq������)��ȉz����=�yS���C~[�����f�����G_����Q�V}�;4��{�I���o;:���Gu^1��"\��#SX�,��V�{#i�Z]���7�����{rY��ļ�)/v;%�͓�N�o��V��9�yW�_P�%J�����,����u�뽋L��%������
1��*�"{�uQ����^ w�IzB�8J�l��'��q�8���j��y�>��>��6��m
�Q��Az�jPoS�������v���x�S���AO��t�a��L�J��u���t���fwd+�O��iXw�q=�_<g*�(���]��Zbcj{
�*OM�M��L?bn.�:��.4�7�ä5��o����ގ��qZ=O�g��F��Q����c�5~������7�,kGo�h��m+q�+8����mEْӌ��������79�T�)y���'%�J����N|�.P�F�T�v���#�����{�ej�y�W�����Z�{')�05�������/�&�w�2ךV,V|4��D���N���s�M�b��a�5�i	�tBp���c��a��LLG1���?�7<�w��[_jz�9a�[.w3�o�i��6�\n._Cn5�#9Z��S�UB�X�����v����(�;Y�K�[���i�(^�b��n�ָsO�o+]���:`Zꁘ�s(1
x'?ë����k����ܛ{�)}k\sX��~�q5�5���3*�^��m�{�7�;��7�P%���Q1��ڙz.9�{Q��N~j�Ok:M�Ĉ�8��hfW:�����*&�p��aC��fޣ���G�GJy�f��D�|hM�O~�cY+���k��j��Wm��eC����q�N#m��]���sЍv�?e��<�#(M��5��G2�D�@ՊR�!�Z���*�5��m���+��hf��YBP�8���s���3�b���S4+�S7	a"�t�"�b���v{�t�#*4#�lљD�ɷ�E>d��(;�ԑ��U�ܕ��2i�-���a�!-5.�G�ڸ�w�1��S��]���%��"�n8𽃙՜fw|گ����_}O�`�zt��0���d�P�{z�zsi���� P��FVE�<�0:4�-��C��	�09o]u_JZj
O/�5��f��8�S�&I+�"f����v����է��5�������ۍ����'�����N}(�!O|�1PR�P5s�G:�0�9��NW-��������1�K�tw,��f!�:R����O��yv�|9>�z+r�ݱ����qٺ�N��t�ɾٶ�	�G`s����kjw�3qۄm�z��j[_ke�}S_sLM|��h\g��Cb�u �s3u��Ko�}���	N��y�(���zg�c�)�9��^pX��v:�[�b�{�D]q�i�>��{����z����r��)|�Õ(��yu�U����2���͓���x��-���g��a^�Vy��s�q~�3���zyޥi��G1�-�Q��)��5���>Ŕ������νSWZ�z�S���3Ǩ�}{z��2rIY�jt�-�f��t��p�{�r2�[�B�M��/'c�u�6�:1k�I�]Pc�;F�h^ljlک}\�`�t��e�4gL�?W�W�_W�H/��Ϲ'��!��r?x����o��ϲ�/*��q1���@�i<����Z_���������{�*�ٟ<A�O[wت�������Gz��=�-�R6�ras���[�$طM�®ݺ�{�����&�Ǡ�t�v�)�<�fG$�����6��~�%���}�w�轓��5	j-�kj���8�(y'�P���;�����eJR�Kyq�ˇ�m|�z&ά�U��.��n[}|�$S�0:`�?@|�J]u�u)i��jz�ڢo6���9������}��票���ࢂLPԕ�b���S�@��H��xn����VƽV�5�=\�{�:�r�����Z,jk&���i��J��K�N9wm�[J��,��7㎼�Uq��%�<"xwgVXб>�ڟN�M�]�o�\Ն�8t���!��ՇU� �څ7��4�Ohb�K�g���i�8v�$����"S�-�y[���HL%���z��F�'J�ye��
��J]������{���J�!��*4uDٲ/��	r��BtM��epW��E��Вe��d�+b�ycL���)RZ�3�_UU}T��ٮ���C�������}�o'Z�t�T�I�l��p�A�/%����N�c���k�N�-0�ue�e�sٽյ��mT�|��יgE�dv�]�I�~`��!f��j�ܫj4��G�Iۛǚq����kc�֞�+G���~��9�yJu�����߅�����t�Q�,/U�`�9�ǣ��ə Ԥ�}��0��_q�A��*��&%�2��w*d�\�4�N!���r�4Jl�����̧�<��ݞu�5�����z�zS�āAT^����f�9/~��%=x��u8V�}sh����q���R��� �s�J�Z��ب�I�ϝ�՗ٹjN5��_,O'qi��Yڭd��R_WӪ�JUF�9�om�%�eH�=ᴮ{=�K�Ͻ�_��b(��PC�BOb��9��b�횘o5�ڿ:V��*�W�˵Z��r:C�#Y��LQ�<��2ӱ'4�^����W��Է�{KGճo̈́m�-����+��s�*����9|�gJLM�)���uG��7[6����I]j�]A��f�G��bZJ�1�;��w��ﾯ��4.�:�}���6�J�[�q{��Cd5f��Ͼ�_p��=j8�,�͎2WjJw��?��4[��v���x�S��>�w����7�-lN�ڗ�U��1��(v��gW؟m�m+��V���x�W�Y3�}x���l�7B�X�kP�>�����N�z��ZqriXo��H�ލ�����s��ܷ���:��Y�|��V�j\h�'<iz5#�g���U����E3z��d��>��T��{Ά�=��Y~Y��s���6<��uo��iO|�8c�Ķ�#9_k�&9�������D�r����[/�>��9��8ѥ���u�\9Q��5�c�Z�NM�gF<ʇ4��q��%uά��Z7u5T����s<���?N��!�q�A�U��aW�x7hU>ːѸ�l��Sk`�iN�ק����>電^�)����5��n#[�M�V��;3�������Έ�Fik�eov��h�=�5b�O)Su�G�>j���z���x����"i�M��Z��Ò5gct��ylm(�(�Iۛ�t��h����o�}UUU�{���<߇3��7���F�Ӱ���=��:��t����	�۠Sr��g>��V�Vb7��Z�M��Nf��D��s�	��2��+��Jӗ0�Q&u�QԯKiFn������v��s�Q�gk��6~����>i���F��i�vMy_(� P����Ҙ���Yp�}n��;��zP����KhE�}Z�U,:}��x��9��G��$�޸k.���{pm��P�.�=�'������O��5��p��뮠�R�E'��O�k�7J��z�ͷ��Úq�s]���/�A������g�gV'Ơ��p��7dXl&�l1��|�N��:Α��8�p�S�%0?AKE|~�9��"�Ş\/��Bo�i�J���m�,�so#]��W)T��Q<�u��VӍ۹��S���I�ӕ�>sM������L*B~�Gj t:��[���}mC~T&0�ԥ��p-*��fC�R�d�u���s)��M8�i�g"䧱2s�A��m��nѽU3e�*ׇ����)�ɘ[R����f�-�.���+��z%K/��nh�[S3��A�d��gS�;wL��*��9hκ��~������Ĥ��sfg�\�oR��S.������&�Mƻ�G"u��!�_ w/G[T�j٩�~�:�~����mQs�7y�*uw{s�L5=�	�r׊<�ٸ�H��}��J��qx�{C3��Ϻ���x�r��)|�×]�ugL��7o;C��&�ƾ\����*�Y�b�_8�F��	X2��N�\_��azW��34޶�B7~��}�GW�fӤn��2�����U���@���JZ�c�3հf���vosH��Q/W[k{�u���3(��w�!���IGd&����`M8�*7�GW�[�b����ܽ��z��n�iW��m�f���QzU�[B��#+�~C�%��ul�����gd�݁h�M�C�[}:� ���0";�v�R���4��ᬸz��M�:�6xnK�򱪓���jͷ.�|%
�8k�i�9"�'�˃~��+�E�u �*�{���.u�Ǉ���3�wmY��%K�����@}+�5��cλ��b%�5G#��kE�5��WM���9�pXW.RR�[3J�}��d��#h����`��IWZ��k4���k�D=��R��J�:���UUU���!Ŗ������Vќ�A%e����(}W'�ڒoCΆ� �U-�2�z�8���W2���v{.��\ur���j:퍘� ��ˤ�*`�KCMi5be\e��ݷSJýK>0Sl�C�P�H��I�\5�X�J/7���/��y	���r��;�;A1Q���_9���H�\w�I.h�UX����5�5�5��D�t�T�4�wˍaB�ș��u��酫���^OE�OZ��n����ħt�Ib��դRw���x���%+b�Mo��Sצ�Mϭ�������NU���\���R�?qO}./W�{��_{ۓ�c�\�����
�W��`��w8��)�hڐ����nW;�L����p�>~{�؂޴��:A/mHt��U."��#� Az�ζ��=E�O/�����<��x�ڥ���jx²��&P�l��Fh���;�y�+W�7˥���ӽ���DSZ=4��
U]
�}:�[l����Sfsu䲴?z��E:d�G<>�2!��KiV��2���fP�����T2�nq�ɷ>f��ʒ��P��MG�ru_B`V��LO(�+4��}}�}��pv��� F_���JC��넬���Y$[U�{�8 �A��p/k:I裼g=O������Q.z��%i��6:1&��A�nb~�����zva~�Eų5��B%]��UaÃ���U��v�n���J��;�ֶ�j�q��/}p�=�5�Q�O 6~*|�$������[�p�xu�ID�O�<��Z�,��-��
�>�*&'[�t1Sb{&�Jb��I�����e�ƻ\^t<g*�lܩV�/BZ��]�N��ԃ�����5��gW؟hm$�܄�EC�s���cg7Z�=4��Mv���}�F�y����Z�q��Ҹ�xrP�W���E)s��H�ˇ��E���E�"�T���;�3ڳ�����f�������y����q�Ѹ�HLN�6;�W��;Yœ�}�	o�O��R2��mּ>�7c!Y�ؙ�X�1u��ʗk�v�p��N-U�Vt�j�z�8(J`��d�w;ve��b�鳖컓*��V�<��7�.U�����U�����8ݳHo!giI{��VҩL�_����K�6�Ρ�.��w�MތB��H��k���z]q��w�p-OH�vū�Z�o�0�em޷�iۼq4_Q$�ԓ���Z.nBkn� �b/�н�t�n�zĴ��ӮDi���5���5�FAqo�:3�Kc�֣ǆZtfAr���w��z�m*�X z�*��xpCH��5���Ht&;�Fh��-.����Ǫ��t��{��ׄr��&�d�N�O�Ԟ�@���$Daͦ��2H�_}��aּw���o���1���Y.�^���[�b=�J.��C�����ة9�h�AAN�Ġ��7�IwS�j��p�:��Xa��۷�E���)�m������\1j��ق�]mn�
GvI9'1��Z�wu:Νr���ْ3�*�����9qϳH��9V��j�K�'Že>�gc#hl|4\�XT6���}�$�m��ٓf[޺��lwj�{�Q.(�C݀�̮X�ZNV%n9f���z(�ݾ����u��<FQN`���ۀ��4L���6:��������J�f����	Wf�2�o8�˫���2M�l�%Z��*qـv��\a�~#z4o�VNeH-R=����$W��H��!�Xg[�]w�&C�.���:wYNw�0c�����!J���F�Wv�n%�F�o#n���tU�uyA��	�j|��c�[�
ŖwMR�X9�J���N�8�x�:/� �X�ֆ�Q�@"l^����D�4K�w��
��֓N�o{R:I�ثu����|�_Nդ�7�������<��>y|ugsN�|z�賳�΁� �i�l��$���5���e���@��,�;<�m�:w\C~���`�1J'�=۸c�.}�
���ZM���vh�v�Q������X+9�in��e��ju�t !���)����k�Y�m^����U٤�C#�@�v9�٫$d��YWKp��؛��.������2�
����W����-��n�xǋn'B�p(1u�x� ��Q�H�l༃�r.��VL�ckK��I}4勦`S�GKOr�d$��S4���u��F�wQ���5�nU�1�76��zP|�NO�犬�f�����-)gE��)�YU:��i����Bջ�<�^ە.a9G�[������YrL/Wt�3b�> �/)�tJ��oi�|DFS��`jX��O����\M�i �ʵm�N�7>p�*�j�1��j˗��KWR�Ktވw�P��&,3n�/uۺ)h.5KSv7&����
�=E藘1��n������6����D��y��Qd�i �5����@���.R<�ZAe�'�5�er7�����޾I��#�w>��O(��eYZB=�ڙjT���U�r�ɒE����fYТ#S6a��*���
ۺ���
!ZAIR���!eH�����H���z�����k-1,��D��(D�"Is<�T$%h$(�R�ڤ�b!M3��UVhW(�/q"��J8�m1�Q��8G�:�!HaGQw\����4�M#M�TJ(�.����B2�a�q�<֨JfjE-�-YTfu	4�%�&JU-C��k1�)���D5%��U-Z��)L������EUT(�-6�!A̱�'CR�V$F�ĤJ���*��6&ZIL���Q��T�aQe��mf�����TBa�I%P2:��$tQQMS4�%��DM:�Մ���YԈ�5BӠDm!��) ���β)l�D$Y���\�҉-*��(I4�	
�.RuBBȈN��=���4�{V�r���WE]/oxgS�R��iC��N��z.~Q�l)����\�y&p�qY�{�Tմ�����h����W�JH�I�{\�/��JmOC���ׅ�����^<�O���v�q5/{�q,�r�q�N�Un��U��u�\9P�A����vk5�����6��l��-94�F^?�w��OF+��_\-q�d>���<��1���&v��Ͻ���m�����/n՞vӝF����V��MX�N̡�[�y[���{�Ns*� ��[yT9W�2��=늘�Us��Ed{Ag����s��9M�T{=�Nf��G��|Dܰ��=��+܉�1��r��C�n��������M�x��|�7�*�:��ՠl��U�U���' \�o��)A������᬴����{������Ǖ��#������W���k3X�Í�d����X�,�m=�GV4�Ш6R֩d��ٻ���y`l�W� $�zC)a�{���5u�1�U�I�w��uw{�f��/�N�� ��@���YC�?G�=gս7��	�������E��X�k�,�*ԬQ�x�K��d��?���JP}wx�y�)�m���N�Ӧ�%J�Eq���e� ��PR''>֣(n�?�`�Ob]��n��AO|�(����o5���2�z���C�0�f�ݕ����G���E,gYG!�;䡊)h���g���8���ξ�xkԢo��n9^+͋��m�TC�f!��(�q>�'5�N֑�-ws�2�3�֛qϜ�;�a�#�*���v����u
.����Ik}A)�O��S�S�Ϋ�g4�5	��#�:�"���gb�P^�y$�o}~h�ss��v�Y���%R�ZN��8SP����ٺ��<_
�� �}I��Ku�V�U��4�^|ߑ���Ƚ�!��<�2X\�؁ZN�򨩟k��y��,�-Ҟ[}�W�Y�2�Bw�n`�Q���n�����og���ֳ�j�TG�f�:F�;�2����l悢D+���
�j�1H�TL[\�)��^���[��z���G1�E[�J>s�]y�f�&mmi� %��k����$-A˽�%g69v|v���6�[������jeb�#��^?O�ɘ t��Wx�@k�Z�j�R7W�W�or�ԝ'J���"m(-�y�r���u4�:� ٜY���
�:���Iʟ�U}Tz1��d��G_��F�]q��TaLTrM�t��B�ݸ��TgY�vu��vݎ0���a�X�,��R�=���-�$_B���\�es}Ҫ����R�Z�Χ��Sf
s";�'i�)J���^8k!9v���=�d��>�z������N����TȄ�z貖���w^�8�y!��f�+bmR}�����1�d�����邾I������ί���ޗ�A�G�HKu�o�>N3^3z��B���~0k3 �=T�bm��S���� ck0<��ݷ�M+��,06��9fQ	H���Y�':�!+��Qt���qa�nk��\�v�ێ\�7���l� _����懾W�����-h/U�)������y:�Z.����íy�n����E�Mkc���]Dr����L]���f�QS��W��[��@���4i�>�3h"E$.;7;Z���WvƤ����cq�z���w�d˽`� woP�f��zÑ�,��$Jد��R��N�Vmv�څ�9v�R�#��&�+.n���Ee���T"��.K���ڟ ���V���B_A��W��s�"�jf�Ͼ��SI��q�ƻ"y��}�/�^aŭ��g��t�۞v�������|㛮�Z��<Gi���7�5zڽY{��Zekr�-�e/Aaz�r֥�iq����Q�̄{ݓ&�^f(����"�aإ�j��Ԛ�м�9F[�ЦZ��n�o^��+g�z��zuv8}�.ٖ�|�Z�z]aQ7˅t�B�vB��:��Ԣ�^O�^OW��-�UÕc��]H��W��{�w]&��o��Iz�'�9�n�2/x�O\u�έD��y�t�P�J�\�P.�9��gV���Qj��۞]��I�h�����B�E'�O�h6�\����+�����놩�Y�9�l��6�ןw�~O|wq-2.~��6&f�˩�KHI��<k�5�k�HMɇ^��J�|Þp����&�[�p^���6�۱R{/�J��r�#�[�li��d^`���,���j�9���ӻ�*;[�K�,ӧ>���ɻ��Z09 u�>(�M���of�Ĺ�:w�{���>պF��ΓI�e�k玳�j�����}2�:�^��߮�#�����g�gW؟W�����OtV�K6�͚���3��ʳ�\����yW,P~G��uAϣ��I�2w��aU�"u�c��U��5R{����U�j�����S����;k��Z�Ӷv2���bu:S�]5��z���HO!��.`eI�r���k��s��(v�W�7���[Zۨ�����14ۍw�"����^dH���nB�7�-Q��8��n�um}��$�8R����V�,M���	Z#kJI!�_�m@�u�*:�m�[��㔾�Z���6�f
�\	�����m�3j^U���1�h���2��[�je�g7�n�Y��)�."�ֹ��s)3�g���P�o�x�3ש���G�B�;��,����Q�:7��]p��k#�1}<&?�Z�v:^C��C���{��̦����R�v+:�l��\�Y�-$��[���O}B�nW��@mߦe�>�Pf�:�:wn��	��s�i�?JX�*�ׯ��	Й�P�n�ϵm��$7	u[9�ԋ��Ԑ��]�J�=��䓚*j���	w��*'���W۹*Sw�G��Q��%x��1Q�6��[�7�:��F��y�S���:@�+��!/zV,�����7�-��P�&ޯ�<�9;�wܸ�����rV��()�ީ=���=��v�5�BΆ�ި�����8�=�s���bEL.d�1t��]uQ)i��������T�86k5x'��8�Z �m��`G3�1��+k+{ab���,o����GZҮ<�M�l?���������Ԯb�)]ͫ�d�u&�;�-@Zr��JýK���v��!qK> ��Ƀ���Rܕ�t�.m���$���Ρ���8��r��!uz�郞ӌ��#�-�zuB�V�~)����5�ʾ�˦����j1p��}D�r��/?H��{z'�{UP�T|����~Gi.���'�ީ���F��ӎ*��`������l<'j(zn1��
H�9�Y�jer8f-/@�3n��2֋�Q�z����F�rI�m������#є���fs���p�'�����| ћ���c�A7v%ua��ӫ-;Ꜧ�k�m7W�C}]�菻%j�[J(���Z[�o֝U��q�%�w���Rv�+��w����R+�$R��)^�v���x��k/\?�j��.��������/�RVDs�kPg\oSWKۆ�����}�fӤm�*�w��|�7��%��#��$wzx؜B�tM��je6Ž��F���*�Wچf�H�Ś�5��p�9������¢b/��b�7���m�3n1�г�{���c���r�,���BW�z�,�+���i��m�p�t0�`����3�E�{l��1ʨ�zb^�k�3P��P��<�J��|�U�.�N7V�6�Y��܀Р��Gs��X@ux��D�$��z�����f��(km�[P󲕥:��L�09ܮ�OE�]c����P�W�|�[�P[��o�8����9NT��.������<�Ɇ�*Y��V���*�o*���ܘ�о�r�p8�����Z��0"kmB��u΍@؍�]Ǫ�5�2��'���]v�|��?���Sl+;F1%c�7A��`��^a�r��v�����w]n�2QQE�@*Y�f��X������}f�߽�ջ��Bi(�Zy��gg$��.z�f�mb�O��S��\�S���jИv�518&K�9=Є�U������B�TՇ�h\^��jw�_kE-sB'"�b��Xeunr��o�h�ث��]�ce���~Dv�Fy��r؜��ؠ@�=���M8�i;��}���cSP��v�λ"c������3�$�\#U�k����۷7��w�-p�x��s��v��{��O�02X��l5*1�ģ�Օ��n�k��u���7�>����3amU�y`�����%�h�g�~��0O1���r�4KC��]p�f󞂰WkFmX��o���~�����Z��Z��/�=J�tc��B8�:R�ԙe'����-s�Fwi�EC�#�yk��+ݣ��a=;�G8.
74������U�il&^���:d.�ým�ݔ��4�Jm��S�~yزT�:]u��E;�%ISd�7pՏMě��4m�Z�	���<�e(�ĞF�Y�LP��5M��5�{H[�J��(a׮�l���Ѣ��Z��"��K�\���~܇m�î��}P���V����
�%鹭���"�vü+y�I��wSП}n�M�r�q���܀�*6Z���z���躞�mD�I[R�*�{��7�᪇�q�y�fEf����#���:l��Uc�pB�!��}N�ZBN��5���a�A��<��/����ɮ��q��� ������f@Y؟t���X�Oaٲ�����OQ1�����Ǘ�48̱��|�z�~F����s��g"osU\�#��u6�b�cw���P�ȯ�����bL�v*����� ���;�[B�RV��I��NW>r���oZ���=ju�5o
ޡG7Wp��=��ٙerٸԶ�Su�MDs�}�z�����o��ש�&�B�V�8y0��v���({tjp�J%3b�O;�&�5i��s]*�351Z�Q*�U*����oxm�a	Rp�}� :z�n��"�ʢ�I�蚭�0å�l޸�y�w ^νە��Sbj2��t�vl�����ck�Yΰ����tϦF�be�o=����Y�{\x�J]ī1���8�z8�}9f*���d7���͚����2ϑ��s��;ܩ)�K�y��;��_	�[�I��������i��#VR�5q�d�s�T���2��[��uKы*�O7K�8��]��4��3Ǧ�΍._q�6�4�x�i.9��)풲�9������Rn��T{=�Ng�7�T�o�����+1��V�2��h�f���[�6��[�ݮ�:�������I;tˮ�ἀ��+��:�6�:��q��Qj˄��.��8h��K^Z1��]MM��[�⦀���I���M7v�����ko>��vM��V%Ru
�FΠ4tP}%���uQ)i�����rl/[�y�c��r��1�d����_����\F,॥]��4ܸ3�&���S*˃��a[�ϛ�x�k�g�#�Ҽ�;�^�x�S�nè�V?�`8%�ջ�-��e�a_ �M�"�-"�N�(^�ngQ��c���A0w�\�ܷ�Z�X�V,�:��9��IC:�c˽�;W���Bb"xU���oq;�V&���S�ݲ��S�e�A�}�YF�X�t�+`���%��o�.yAt}��T�VsƔ���Zp���܃7�.��ʃVG�tz�wWW5I���@%����N�n��P
�����3)���j���G�\���#5:w����:��vm
�(vQ7��jԥl����]�4�742��&�OjQ���r/8G�L�N�F�+WGx�z�(�s'y�am�Q�P#4�<�R����`�.�l������P�Y�\
����y����;2�",�!D�$�-�`��|.�X�Kk�סQ<w�Օ�C�yK�w-�z��rkXƦ;��HFn��`ئ�N��,;b3Z����6����{-����dl\����b<5�a�c,��#��4�aym�8GU�=ĴC�Pl�%x
��Vlj���M��ݗ�E��,\a��&�4���sa�M��Eg�3��s5�Q-ڙ��s+K�^;�JE/��Ք��t�:��mZ�[��F�Y����:�\��7�}&��W,iج�S��u9��v̊��
��H+%�pM�nk)��5i���Nv��] �L8ܹ��wB���ؑ�oVΣcF#;{3�hõ�Ҿ41�;l��j�K�9ZZ�w�Y�Qd���N Ż�:�n4�ǼV���uyN^U�n��1�MT�Q��M��9�������P�5,S��!+5�t��a68f����Vؒ�X�� �}��}#U�z#��.p�jV\q�ܳ�"�%
����@�FT��}��_SV��!�:�]h�x�} :�����4DdE�fJ��{ի��:�	�Ι"E�g��wv�7cb��	��a�+5�x�	@�ݏ6�ݲN;.�&{����k�k��m=*��\t4��ˎ�@k�cn�u��70���*��h�"�镉Һ�}��f��g�5�b!Ʌ�4֚V6^����qX�[����4X���_dVd%���d�Z�2����4]���he9��(����֓�Yѵ�_U���H�@�7��9^����|�������_7Ƹ��Т�+L�<��И���V[��Fuc���g�6],������Z-<��L;I�ܢ���:�:�%)mUԳ+�5J�����]U2���̺���5r:��*�fG)֝9Ƙ�G�Ԯ}sЮ�坘�D��\�U�qύm�΍��Z�SC�i12�#�Y�����V��#Sj�̗ٮ
��k�VA}4��ɂ���P��D���h�c��䡮�5S[֞4}�̀gP��ZS��s3^��qW0���k	��n�Q+����/�C�̛M�Jm#������y{��+ʄ:(�,�*Ch�**%��B�����Qbb�)M�EUU�PV%�VF�4T5$�**3"3���
eQvEaE��UJ�L+E0���\��jr�0�T�B��\"9*F)G*.f�f!JRUe�Q�JT�M�%H�DаJ!:�U�!Ą��**��)2k��l�-
�2p�F�ȮQ�@��KP�fZ�t��@���.UBXQH(UYsR��i���EW(��E%�Pi�gH�VVY�2*��L��"�ꥁ�$0�Y�[��*�Tˤj![LȊ"��6ja\��(����D��ReW.�D�5"��j�TTTZ�Y�3,Z�����b�s��a�Ka���SZ�aTU�
��dp�H���j�l(��U0$.2/�o�h��ѷ.Tg)�N���n;X:�;��:�/v�dAv+ulْg
e���K^���ڰy�f���8$�0'��Y<��hs��DҸ�,g06��</��!BVv�
��%�el�掁\\�r��ru��W>m���͜�T�ɕ��pt�,+*T�U� ����X�s�[�7�}���L��?�q��[ud���P-!IOV`X���D�cfl�LA[�s���os�+��H�N%fT�2�]��|�3�jvx���%)4�h���yW��w�;�/>��s���E<wĮ�s�S�������!{����ӗ��N��h�yYo.'#s]B�b�u3jBqϝ}�\�/6z�>���f�F���`���]��W�$Dv�r?u!<Yt'[S�iOO*�{޷G��W��+|�>x�ݯy�Ab����x��X�lр�T�����Q7Ɋ䟯k��[J���z{⟙[�lb���X�̎&ZG�6��Y*N���r��Ü{�\bI҅�����̨�g�����F��I;�3F#�%N�lc�h}��N�w�QA����yDµncS8��,�s�.s�vm6��ru�/d���A<�r ���yuR�S�q��l�+_���]�[��ɨ�xvi�N�`S��������\�p�"��SD	w���b����]!�k��"z/���I��j5o?�tr������ޖoc��_N�����#'�R���u��؛�:ڑe8��:��p�(z;_�g>��1O��K��D�X6���(�"�q�*�J|h����jqx���ƽ�*���mx�Z�?C��i
��u�}˶�)�aޤ�ƶ�5�����3�f�[Ϸ��!ʍq���٨�\�"S��o6���G��BѢ(����<j ��\��~�?C��j��f�<��q���K�;�܉�zٵ���pVˍv�D��<���u_�nME�=�E� � B�c��yg(�{uZj��g1)�Ɓ_k�9��_mi�Ig_炵��^O��nA���^�ڍU��u�\9�x��w9��:rr�5[�$CfF�U��ȮLī`�&^��kҎ^�%�9xz�P��޾�YXF��$�c�{Թ4<}<n�4��G�ևg�JR��16rK��ݩ��A4j�R�w]1��7oggu�%m�ηf$$�7\�;�Z����0HД�Z�I�d��9[����{��L�Z�Jx�������\k����c�Z���[�eP�nF�ޝ|��M��s�o�����i��ף���r擎�˴j,A����ط������_�aE�Y�\Lu㵏��]Fo7��`)I�.�gs[Nv�r��4��F�l��2�:��aF�v*��*&���Q{�Oh���M�M-~�k��h������#��&oZ�r;{�����1*Z�M�fs��55	�g]���^ć*�0�?l��rs�����R�Z���e��-�{������Hq.�ԧs4��{,���;���]!쥦�����]��5�痵j̓�P�#3�u�wD���@���}?%�����`YՉ��susW �EV�W�Ovm�����(�!Lw�H`�KDj�}�<�[A��]��5�i6R�u;�ׄs����,RU(}�8�gC�7��\�wDⷧ�!c�_"WJ���F�����װ�v�u�z�/��
8�L.���f�KM��uFF1�Y|�
�����2է6�Z�p�:�}[�ȝǹoe�srVa)��ͺ|�1<�r�W�(<�P�ȧl�"P����L��@J^v殸��3*��U��W>sP���<a�7�	�6`t��E:wJ��,�$��pwT�E�{7�����o�w�bi7�!��dI�/��P�n��zJ��i!B�}���va��gM�I���L��8�̭���<lm��#��pd�W>%��؍_s9��L���ߑ����q��{W�O�R�Y���35�~���LAe>�mOS}�zeY�m9��Q�*��D$�ޗO,��ogL�嫮�`x��81o[yC����(�J힞ВSk"�+���1H�TL[|�)��oE�{��������Ek�fϖ��y�t�M%���k�*^XS�6.7��ݿ�ŝGw:�%	��f�q����,Y�g�bCX(��ߐ������\�E��;H�7���fD[z��B�(���Ph��7v�-_wZ�X��������&�m��u�����.E�u��خٹ���b���O�̜�&����99*�$)̡�IQ6��Q��N��	����޺�l�^5���>���R2��h�}v���UXp�l�b6�6z�e��p�L�.hZ�tV�k�W�OV�{n��uA����EG��Nt�tO/�$B�ߡ�ʙ}�����[��ӛoBלoT�B�wϲ
�&(jKU޹��ޭ\�[JF��k��{���u�����C�r���W�wL'*�&��M!c������M^��khOI�_�I��`���r��!��Ԫ�5�75�i�h�[���q����p&�#�|�����A_��e-�oohbQ3�a�o��m갡���^��Lk59�K�x׼��CI�e�&f-�p�:B���Ƙ��0��tB�ӯM�ܫ�4;[T\���8���o���f��Iנ�oS�O8�h�Tk�9��Y]�/2��Z��T�κ��ri'z��پ|�u�p��ӉS���-��f��;+q���������쀡�L9���H˥0+�]�"h\�\��\'tK���J�P�+�����~דl�ܯf䝤�}'e璣įW� ���˲:n�el\���wNqq�iT�2�Q͈e�u��c�ݗ���uF2�c\|�mLY����,��뵉H,/"多˝n �{|�kY��G��N���3u@��/$�������p-uM�P��\g(��|�L��D�]p�f��Kd�gdnFԓ�8��R����U�㛝BS폰����3p�6���<;��8lvh�4w�~x�����ZW����c(ʓj��tIo�k׶�V�xQ����{m��:����܃�A�R_WӲ�a��5���ć�{S�����9�z{��CX��_KO���D
�Ȃ��|����n���wY�����^�ۢ�%�5���m�jrۈ6�D
?wχ.LB�P�����(��uφA���O���[�E�ˎx�g��6�3��y�'q�I��B�_�n{� ��f
U'ht6yf�X�m�ҿ��Z�`b�]�*�&`�K8ݵ�g�)�(�=�R4�f�is܀�Wظ�ri�,ݼF���0zU�S�?sa�HΠ̴v�n���G�l��+�����%d��$q�E��܌���к�A厙�T3�����N���u��/��E�(��U�n�e.S��u�]=*�N{�d��P�ƫ�[Տlɼ�M����Of���E;fQg�%6
�=+�v7�QV*�fR��E�P��uZS�]4����\k���R�����3/���Q/�EC���}j=z[�H��.��N_���;m]�Z}�h��@ք���d�:a����S�1fcV�K�T���~����tN����wS�s��y7�cz+�n=����YGc���7�=�pA��=�*��6���au�6�z��t\+u��DwS�۽�yd>����V'��߼`E[�S9�5S�v+����b��o)�N-J�S�x+�:�T{�貮�g�1�W��|�����&vA.M�&=Ѣ�����o�ٞ�&3M��@��A��s���G]o�tZ����rV���q��)_�Q�>#Ъ_zNS��Ӊ���mF��EωCne��Ez��5��<�T\^��]�>�%ﴺ�)���q�����֮;�{q�F�𸾒O���l��?l��=<e:`�C��GJ'�+�S+f%��k�Xy�W��H�x_�g��w�3|i�(�Ea�8�]���Tů>+�~����,fI�Z�����h���r�V�dt�x�I\�ݗ�U�R��f��)��b�a�OB��<�1i��)�0������qmY0o7α]�$srlS�	�%p2dv�+�8t��b[-�b�Ӡ��������$R��c?�����J��J���X�������1��,�y�{��F�����Ot�o�g������IZe� �H.������."[���^��*���Sڰ����EoK�ޯT;%�D@�-�g�x��1��~W�z���rW�M�������{��er=��É����z��d�9���Anx�-n]��<U
��~��Z�q��F��{���>���>��n=�^��~3��Ih�-�ďT��<�����=�;��6}b��m{Ǉl/���#Q����n=��'� �w��"��sl�Q���ר�'��W4dW5��R���kD��4.2�.5�r��㟪G��Wtbן��~>��_3Q��0���yJ�=
r�z�>�r2O��]|2c�b}�*'�oFV����c�9��c��{��\]޷;�/��ѱ��k��U��䶤>%l�}bwL+�V�T_wuxh}���Ft�bR��r}Vw��:�����K=ׂx�{�V.�H��e���.�v4T{T�~��(}p�Ļ� ���M��	���STpu�ݾY-�\3(����G/ˎ*�|n�B��W*�C�w�ҳW�N�t!�b���"�w��1��tNa�;�Vd�h*�L�g;�%��Bvm�尊�ij)^#���#G��R|v ��F��mnZ��@2�*J�	��ğ���?L�M5;q�s�¹�9q��Ӥ�#���~�EG����Y�<���Z��j]C�G�����}GY���%7�Ǯg�^��v�]�c�N�&|)�m�ģ�d�}R��4�yNl�^�~9~>���<�Tn��z�f���e��~˚���w�Wzt�D��2��,]L��ty��a�F�W�����?W�U_d{|��Z��P����o�+ݕ,ݟz��0�ARĒ�论�����<}���kDx��;Ñ�Y��3����d���޶=�>��
�\�iIUa���PVZ���\��]���g=%h�|���O������q�!�j�p�w �*��<���&u�}���۸Q<�41��2o�uk/�j��E{��o���"<o�i��þ���m�i��2* Ej��qY����p�h��j��ԧ�G�}u�n����7�R_��״��zgt��=�\Ozg�A�u+�E������^(��S�� ��4%9^;�?F�\��^W��G��ώ}�d�yCf�M{�+_�+icR��(�ιC`Es�Wc]Om�b���+��Z�k0�U�vMl���dvըʊݬ��'�:<z9E��g��yҜ�Xe���7��,pd^5]�S.�-u
��nsE��W�5v�e0��ֳ�)�����T�T�d�36H9>�T�������=�f�Oa��}^�q�-t�}ʘ�����y]�6�٪����L���k=��8��C7?e�5
Y=P���>ʁ狂+'���^@�}-T�]O��^����5Ec�y��g��X���RB������
�[����yǄ�(�/ۉ\�h�}���m���O�h�>��7�ۈ�ܱ����K��dTJ�nwd�=�1��H�Eu1��O����{iTyD��q�^�Wx����~���L͓(Ԯz'�?�U��P��̖�q��0�r��f�~�_��~���W2�=걽d�W�ן������㿕����:n8�wo�1��X����pi�Y���������{���o!��9
��S�+�t�qO%�Ҭ����g �T;�U#u���5Bz�/��s��]+��X��wO����^Y�Có�yh\C[R:�x�Ƥ�TǸ��a�HR�æ��C��MB/��~��}�]ǳ��i�������yׂ��X6O>^��K�u}|�������[���/e�y���>n�}���27|�w�U�e���7.E��a� ����iB?ozqf�sq����K������ޡ�2Y������Z>T6dō6T:4��l�Æ�����|�EV�
�ڕ�V��iP·+���;S��h\�ȂF5��Y��
���e"�{�w�μ'��/�e�Tʥ
�Af��ee���G�^`n[Z�%H����}o�n�ѻ�z�u�*4��^~�5�߭z�o�{@Z��+�f��ً剌Jp��r���N���Ӑ3ה %Ҹ��WZ�㴰���s��;�i�]�^7 i�J �=b���L�n=���5�b�W�-�'I�a�P�d��@=�T64������g2�=ywV�E��CeAX���@�l��2��UV%]�v���}|N�}��p�:�EpV���MƢ�m�d�Z�2�Er�D� �fp_B��j��z
lV����](W=m�>��蠋l�t]��ڏ"pJ���HI�.��Ό�Ր��Ԛ�b���V�B�e��ǖ���-�۵6e�e���֊�x�{]�ۼ�W�X�M��|w��������9s���X�sN��ʃ	�fwjN՞[��@#lhݓ�WX����X�2�Y&��3h�GjQ�86�5�sF�S�$��ԣ��c*�ϯ�7�n��P�㖤K$]����p�%��v���W:�b�~0�t���Ҹ�g3�����9��&����s^Xq��mo�jN��x�7t1U���λ�ڸ���,o2O��T&h�+��,�`��m;��uPӻv�HlL�0x��M���A��YBv�b�][]W��!S���B�ZTn��м�te���/�n3�k/͔��o�њ��zS�J��i&�x-eQ�d[�F��pdU�����F��r=vJ�*�]��!L{��+jj��.����������GFEo\�k�Fo�__:�L�5Y�FM{WX��\�҇5���V������ ̚����%T�&Q�D�:i�D�����{ٯ!ɺ�9k��ci&0rR�9�j�+j�CrIf�P.v9�d��6�K|��%�تg�[� K��i�c� -H��G8eF��rxʾC�qؖ��ǖ#�p�L���攘Ԑ�1��7C���W~���D=���2�������\٧�RTq��Ơʫ�"����+���`�'��s����3c�pt��W���rX�u�*D�N�뫇S�kY��Ӷ���`����CZ�=uQ&�X�cۺ��u���VIDp<��F�{ʪ�q�v��ov�(u<�Et"�J����o,�)v�BYDb��%ry������emY������-V�%@y���=f�׎�vY����"��&_��u7K���O$	^S4�@}�w����{J�'5+4��jI��$�ՑWNj��TTU�2�G.W"����H�*�T��:�*�T�H�HG((.aD-R��
���i�H�*��D��"��9�\��J�U�@��V��&Ά\��LI�D��#.p�)9����,�I �9s%:*,�D"#32�HB�,2@�%�%�Y�*Pmf��BrKCS��N��hV��RZ�U��ZVYʹGD���Rr�L����L�-a�l��[R���*4�EI(Y�P�1C1R#*(�LԥTJ��
u$"�B�jI�����dj�GYaR�b��J��+���2�l�3%CN*��w6mT�em�UJ%]h�i*dt�Y�E�
��.DfE����G
��f�������<���(�ȏDM�RV%F�����0���Buh�h�mf���v��u�:�w�1h�x��v��jX(�c(�2!:}�L���c$g��iėr"�eo5q㆞>���87%d���G2{ ��]O��ubo��q���"=�Y�����gv����v莿W��s�S�X�Z1�3}�b���x���o�E{Ԅ�O�hhϗ�����H�����즠2O�~S���„���/����8 7_ ǋ}$\��;�΅k���"}�l_S���0*kxF%��k��O�����Ϧ%�YP���	�b~���7�-v�G=j�`~��S^����z*}��b�h��H��=8>�� ���[��ʰd6nI��EQh�{��3=�}��Fo��_(�g���m��Q�{ԁ�Dx׀�f�
�t��)d��*p3)�O�9.8�ɽ�;�sG�+�m�g��/J�~�g����=��h�����C5B�8�&Mt�=#�]z}�-��SS�E�Q���������t_�Z�ؼ�ǝeC��v�c�Ez���{ެ�eR�]p���ݣ�N��I��s3��ǉq�<�ᵡ�EO��T�������mޏ��p�z���ʄ��Y�s��2/��Z}�^��C�;ʜ7k�]�	��ݡ�O�X��ʺk��L�+�XÝ�{R����K"|361�[�~T�κ=�����qu�������v ��%,�{+su�h�o�B5�7o62�v�H���v�9��r)r��M�p��8�lޤ;�˾�fBTQ���kY�9C��z5Cj,]P�Lu�u	(fuE�ՎN`�������\���F}�x��ǽ��ŰJY;�f>U�*�٩~%>�O��f��噰f�^�QO��5/YJ�.c;g�����B�NI�>%ٗ���T,����^�	�h���r�>��p9�.�>�'/�ݾˏx��֮;�{q��S�x_��I����>���3}��mT�+�7���ީ�s΁����Vq�x��C���z�G�A��Wg�Ec;�hU?cR�֌��$���	"�Ԫ^9��7MՉ�����w���纋=�QW��Q�깜م�;�=y�e֭>Im�`O��H�R鿼�����󄋖�zR�S��՗:i��Z��o�T4���'M�u��f�<��8[�&�=+��9�D�D��wML�ڹIV�N�� �_Nti>��ꑷ�bi̗5��>�s��rAe�:	���>�{��Ϫ��q��n5�Q��'�l�A��x�d�=��@��s$�D�϶4���n�Ĭ��Ɣ���w$w�zV�R�g�o�K��#Q�ʽE{��O�N��16�_�
�-�o�~g~���k?c�q���������j��m!{u���ƞR���F�m:������<��<ywE�.�8j��\�,Lo0uj�Q�E9@w�J����3$��ee[]Y�r�a����L�i#��ѝ1�3�M`[S��8��2a:�9���.I~A������c�0��M{:T��
��R=~���h�����ss���^��u�أ�G�>�t�r�X)�/�A5��k]{��u1���C���Տ,'�y�jz�nk[9��k_�^K��E����|J�0�D�W^��j���J�4o//z��G�મ��畽���Iޑ�]�����yR2�Y;��;�r|�lq\��ީ�>̍���u�~tK>^���J���q8�Q�N5u��s���rN_KN��/��W���_n��U��/�����GI��^Wȉ2�Y8�|��~w	g��7s&tb�y>��ax����=,e@�a\T�:. רyN��K�.��t�|�}��j�е�$X�J|&v5����1��t��>%+3��3ŋ��|��[����֟W��������������L�}'/�Nt��6Li�O8�ʇ�"W$������	/M	�;n�m+���~`�ߴ;��5����D>�z����
��F�I@À<�G�e���=��z�Պz����X���v\���1KM� ���<=F4u����c�����u
��mih��&���zѕ�7y��k0�!�P]]�}3�뽈Mת%�W_*��cmK���e�ծ3GM��Mz �ǜSÌ�V���!����u=:�Vu,�/[��i���<?��O��N/H���Q�ǵT��uL;�%R�����~��#���ֹ�5�OkTez��9ǽ�ƣ�O��n'޴�A����I���\��gâ��]S�=2�6v�"�zҨb��'(��t��)�1:�ƵHvD�[f0�:�>'0�����󃹃��-�-��Zw(��ş4����d�}
�;��FD��4.����χ�|�F��3�O�������\�f��^�턯͊���CS�����|�/��r�[5ܩ�_y܏ݏb��
�Țů��z��:D����n4
~ːQd��2>ʊ�}[�#nW�W�z��\�����2k��r��>��u�������}@:���}��X��ԃP�Ĩ���Qڛ���$uN/s��<g"���q�]����}��}�19�y�X�/fr�X(��9�.h{u_Q5��^��;�6XW�VSp�����/���j��.k�c��/c��'����=^��S�\�zj����uEsH,��:|����A��gG�*r���*�;����W�T��}:�S�K�u���+�\ɳ64~���-ut/��nʔ�9���j�Mq8���TJ�`�h���;�I`�{d7m���*"͟�f��y�w�횷�����i�5_wD��h��@.�Q[0� �����%�l�2V~�A�J�U�| ��Cy�ܻu��7:�;*�fM-=����!����1q��:Pd�i�yP'ȱqY5�K�<�4���!�?/8���
v1UyZyƽ���l�C�C������*x��)q�xk�=P��(�[�3���'�.GH�aK�3�#pn��R��#�^^�C�TD��-��qsĞ5%xѕP�8�BC��􊋍[ �o{��}��o�n�q�{NF�G�܈�\{�r���dD�pW �*�K��W3�Q~���U-�ǵ�{��늙}(d,���n�M�w�9ޑ���K=~�p��/ϐ���yMf��fNm
���yϣ���Fx	�9L�ql��]�����Rs�Z1{}m�H���&�v��{��w[��U�������Yo���Ҽ�t9Я_��t�r��Ky����џ:��{��7Еwo}!�H�z�'\�j �@/��|�C%�v�Q�8\v��јLϘ���T2ws�ސǾI�`{҉�x�D�#��h�\MC��ʿ���Hȗ��#b�c�|}��w16.=y��+�E׵\&{��c}^���R�5�{!��)�93_)d�2�h� G�LN��:�����؜ڽ��sjZ��w����5���R��/iݿxK�봽�CA`� A�b#������u��[�v�v�7ㄡ���Ӯ��j�,5���K {�3��S*;|�^Nu����6T�dCzg]����P�3a�dr7�==��^]{Ǩ�G)�������;�/J�4W�����߸�&Nw��r����R�_��g�Hz0������*V�������;ۇ�߮чމ�aP&�b�'F��L)~��O��֞��䶠d�WkC��87�n��ϻ��\v���N}�����*���])z��;�y��=z�E�w�8o�,�ۃ0�P'tú��4�A܈�l ���1��:����l�GL�k3�z�����#�����T��,��3||��eV��/*UxSsї+���:%y`
����p�Srr)�j�MΎQ{h_ڧ$��o�/��
�F
���OA����B�eV�W.g#�}ޟW��������{ǽ]Q��S�x8�V�Q�0`y,���B�I�L��e�T�Sޠ\�k�Xy���n3�<^���������pJ;��o!��>*����.�s8�����z��	�|�*��Z�,�Suby��4/���cf�p����uY��7q�5�~W�4W���=�g<a���H���`\�"�K�ʦ�)��"���~���ᝒ'E �c%R����>�6Q��@u�N۝��q`F#YF��
�J�[��إA[�q�#���N����u���4��g��sF�����6w-*���t���w��ʎ��27 �z�7J<�Aݚ:Y����.���K�����R�1;w^�ĸ�z-ZJ-o��C[I��w�i���HN�t����" y nx�=+���f����}R.��>P=Ͼm�����X�ey�~�M�}R7�,K$�H����!8���®{�7��+�����聳���Q��F�j:���G�����N۬����2KD���7���beziE�6��V���X�R�#ö��q�F�o��~�~���N��16��^��4���'L���o\y耿��	�s�Հ��4.��4�S�q��#����f��jDv��=���LaDwG.�5�;~��-��V�K!�`��g����m}�Lw:�8|�ǧ�
��֎-t<��z���	ވ^�.;�R��=�;��z�M¹||��c��'�Բp���Z�P��W��/Uy�ޡ�K#�x'���V.�H��d��x�ه�끮.&��s~�@��2}܀s��jy��Y�/��WᎪ�įLk�M]D���8\B��9q��ӱ V�p������/j�-"��ʭ6j|�G#f\
�^Wȓ+œ��̧�Q�����=l獛�UQ{�	�J�U�@���7m�ޮ&�=8q]uh-Zr�!ٴ0_D@�Ʀ-75#��AlZ⠠��sn ���Ӯ�Y������W$gn��H�[\���զ�����c��\�α��6�c��in�]\��\#�r1ڙ���'N���x{*]i�򜍙`+�.��t�|G���ޜ��
`X�GEw�'Ӿ�~N��.5eO��R��g��L��ty��a��}^ >��;ї7�~W�O�oW�VG����3|b�vT�vXFa������H�T�X�8r2��s���;�;�������{'ޞ>ĥa�	j�\��d�u�P���mzk��h����K�Z���ן\M�-ߴ���<��D>7��T�s,>�%T) yH^����:��3��NR���� <=u�o���k��W���ޤ����zN�����zi��z�v�Y�ὺ*o#���}
ӵ���N�/ō�ujP�/�ٌ��:�;�~��Pv�����#׹�[����*�2*�Ly`�"~��2*'�s(0�c둷�[^'��*��4�V���ՙ���:��.(����d�q�%
g�B��k���Tǽ�}��;ɚ�sq�{�U��c�ڮ�\6���#�|{>f�@�~ːQd�� �|G�c%�n�ڊ^�y�0��^Wn����ݬ���F�N� S$d~	e���_�)�7�r�4w��M1��V5M��:��lI���54�aC֙�b��U^�V����w��sc�з~s�=��m�γq�O{�i�OmB����N��[p<�H�؟YF*�[9�Rgu���שs�"<Omy����{ή��}@:�~����U���Õ5���G���+!.A(/5H�+ģ��WS�q[>��R>���X����ޠ=F��u�yt7�ٜ�)�i�}Z�)�s�=���r�X������6���P�~�;#����B�}����d>{�
���9Ŕv+ڻ����?���6�;;s?��:��iW�wT�۞Yꟳ�Ǆ�qD(�.�s�.{��+�����o�x��ѕ�5y�^���pi�Y��>�s�:��w������f����+j�}�x�D;�;�G����C��q8�P�������evǝFGxf��������q�Ss޹��8���/-�dwD\�'���8#kd�Ϝ]C4{W�J�W��2����p:�T5���9�/s�q�)�����_���vc�72���fF���ޡ����1�B��n|��=�X����q����t�z�����Z�^3﷓�p�.'���-9���Te�!J�-�2#]���{Ԅ�O�hh�����(E��U�s�F�]b�Gi���75�b���c��T���%9[Yz�#�$j�^�s]��is��k>IǴ�l0���W���<V7��&ViǓ����sj0,xD3��(�]�tȲ#����a�6�T�R@lШ�/�Roo���wz�DѬ��^'���,��	Q��-��g�y���΅z�hp*-�hb��W�V�5����NwI���\N��z�j��B"px���z����-u��U�;�`L��t�@�c�k$h�^��(�8���{ՠ_��Ng�*��=$�ӝ�gQ�����T�wGѷ>��Ϲ�?��5pڿQ�{ԁ�G�x�ϡ��K�9�O��b6��n�=D�WsS�7�(�n���tV��I��Ƚ*9��=��p�W��~���3T�o�<*ig�t\W�"��J�_�L�1�O�O�Xs��Zpmk���|y�T>o�h�>�W��Ku�ѵ5FF/=z}0%{��{f��p��*,�����T�N�Nx���c��w���%������U�7}�{��΂���׾�-�T�,��3�wL;���4�A����Ǣ�g�yQM�Ԡ����2�Q��^���;�H_�yRj@���'J/lS��[P����B��3).@zl��S���P�yY
JnJ��F����pY�y�z�$��ωCk���clR�X���H5����4��:WH����Y��p�0��pYb�,�n+-%��Ѡ�N�Y�Uw[�Sͮ<��c���w%��u�%�t���K�����Fvu%;&L�Ȗ�pc����.��b�,�̺�Ht;�e(�b����7fj�(��-�#!��R}\�6���.��>b�&�<*�L�{��͌*�D�&��M�D8y��Z-�y�S�u���� �xI�_|0����.����.��%>.����ʛ�@���R��d���� �s�4��\O�(�"v(��[���d�;�|r��\�r���Zҝ�7�o*'t:���#�`���!� /ޜ��)���α-���=:����`r�E>-�%�8���N�al��Ժ
9X�r�r�]���_o�a՘-r����{��Y�Ʒ�Wa��v
����ef�����S;��ֳ�4�����UӢ8𳙉�'׉-�GQqd�zA�fm��<��b.CXt��k�R��a��'�v�cG=5�a���\(A�|�����$;u�}�Q�Tk��6��R�jp�س�>��;�i.�lnݣ�~e�/���&����Z뗋��b�K����r�;q��A�	��d��q7`K�ţ+sq�k��v�ɴC+I�����/2�(��y��u�>D`�'K�AP��3S=xzoW6�̛bO��+�/R�Y�uԡ�Q̰���68�YKN��3���-���Y2"(���C�!B��2�N���_����B��K۳���;;ዔ;�մ�����U���ٽR��w9:�yE�%�j��v�i�#:s;Yk4jt�@�Ө=d;��q������lU����M��2���R�T�nB[V:�C�����
��	����$yu��V��<N�-^=�T�Y}Z�X��2�Ԁ��ù����Kf_�v��W�D�eܗ�(�{Oi��[Bp��h�rͣ+htYy&��h̵p&�KJ:M湑3��o��Ϻ���f�oMK���]�DH�W�r��H��1�Sd��(�c�1Y��o6f�I����W�k�ܭ��s�Q�w��7v]XiT�4��b�	�6.>�qd=Z3
�����iI,Q_-[1N�W�S.�{9N0�-�Ư����cK"_�;�S�j�S4q��N�]��"9�Ho.+ut������
K�>D.'��̹�u'S��9�.����ї�r���Nh�S,�ʝ�qVu��g���.��|��9<Ћ/l=x��:ڔ��j����R�Sf��9���(��cP�l)y�wU�P�����e>�6uer�K1�n�U�u���ƹ���V(�G��,٪5a[��&<�W�r�\�s�J�(N�:����2���<����ą�)�2wN@W8..�l�M�{{�����H�_]=:���8��u��@��9��#����+N�R���~ϊ%濼���=�w��yZ�t���j���s�$�VFh$�A�C!+(:Ӗ��F�괹�NZ���A��V�J�)LH��(
<䄇2�����-GOO+u��mKWwnWR��L/Rp�ZQ*���;�ŉ��j���"WK��N"�i�d��.jB!̰�MjYt���u���u B2���0.%b!j)Q%)aVʕ7A��b`�e��FEFV.we�P�CC��	'��Q*��,�
�\���[�����J-4�����H�GBf�*�Q��Qu�
�\���HKE�	*��sL�k�3]�X��Yd]��e��5N��b�'"���J���iY����%"EBUݮ�x'B�s�Z X�)F�Fhr��<=�)����T愞��W���8fn�h�
��ؑ��EeC��߰vT�@�S^VZ���O���w�e��ʵ�kj�-M����)@K�{scf-p=B�fJ���?��T<O��}��L��>�i���z�=��֮;����w�$��nj�/�3��'Ei$��x:�L�wS>S�As��A8�>��������Bӯ?s�ޡ�����h��s��5�F�ܐz��'�|�*��Z�,�sBw�~�����Ux��GYQ~����E{C���Y���Ǹ�JZ5y%���v+u#-�y�0��֓G�P�ٹ9�J�ne{�D�ף��+~�P���'M�u��f�<��8��iofP�
dY[���64ɵܕ��^x*�f�}�q'�V���+����p�n=��~�bi̗4���K�Q�T�̿cm���x�DO���R�}��5�ƴj:���G�����>��n=�^�G�<gѵ̎���x{��U���%q�A��>�&W�
��T�����7��m��Q���ȟ�����}�����h}w�u��5k���G���30�c�}.{ƅ�[�Ʋ9S�|�R=q�+�1k*�lzkȊ��U�9��9�@��5!��Iҍ\�Cq� ���qF�_G�^wS�!0������=ё&�=1�D��{@v�4�5�����AԂ�SZY6�NE��6�F`�����[��=��gԷ����8�6�R��X^6�|��΢�q�f�@�B�7�ep�))[4a��v�Z�v<U5�>��llڽ�TUd=��w�v����eo���|��_�}A��?O���^�.!�G,1������7���v���d�����qx߶�i�=����ϸ�}�4��bt�{�V/�yR2�e���8�U;�}��۵�;'�˳<���ei������/��m_���i+��[WQ;z�8Z��9^�e+��U���zB�I\��gdEDZ���j�N�
�t�d:�~>'~�O2�!��r��G.���6�?I;O��Z'mO�@��_tT����ӡ�:K-.��O������e8�-H՜�]Y^��q݉޳����,Z�g��L��!����>���ۃe�NuV�w�jzݍ�1�l���Hya����F�O�,tEL�l�\����lo�f~?��_���%�#�?V��'��G��}{�Ǹ�ӓ�X�(�,���8�7�Ǵ��=�:��W��G�~���t�\M�w�9�#�{#�D>>�23�S��T�]�\yUx{/�Z����z��6}��F:`�����ucQ��Q*}�H�Nx�;��'O_��#NF��]����p�j��Zy\+���މ��vۧ3�5�LD\�ʲS�_w(+��x�:Z�j�(r#+�48������~�n
彮֡��#��+�W`���8I�����q��t���/���[_�ڒŎ&{�rO�ak�o�v����O`8�[JF���X���P��Q�p7:_��@s��kT�d�[f2����w�C��Oj:m��^z�yQ>�]q=n��E|�K4�a��#"J�I���|=q�W#l^��,��^�l��I�#k�h�GKVY�L�%�F��v�&��]�}f1Y����4}��o�@�b����{5�f��+����\�.��7>'����C7D?e�5)d���*+�6}��xR�R�qzh����S=Y�p��?u�g�����P���i�g*��{jA�S�W��Qq�qc.�7�j�>|��3H�c}��7�������Y�'�rz����D�Ǟ�(�>Z���ԝ����g��磧�f�䰣N��Y^j��<s�_��m��d��q���Ew��[]1�8.p\���\��~����Ǎ��������_��(���9����W1-C�yJ�c����s�W�}]\������Gz�����"���	�,]d֛�N��"p��7�e�mw�{��jW�d:~��u��wHHs��|7�(X�L�EW����TB�Q��Aл���w?4r�_�V��H[z	��r��+A��{�pZ®n<G���]�&`���,�o��d�c��۪ɜ�gj�����9���U�S��4�"�*�η��_�2�Ք�
}<K��u͐�8�uȄI"%i���G\ŗΊ=	-�8���*����j�+��d\b����+��>����п�ڑ�sĞ5ֻ�n{k�=ҪɿZ�>V���Oz���`���1z��7�<^����S��^���mն�NH�=[�JW4K�l�$��g�HJ���2��+��e��.9���/O��v^j��D��ͻ�t\s��w�6
5( yTA�"�gKe��u�9^�!7�Z){ʏ���{5r�B�+5z{�݇Д�=C�\Nߪ��b�J	W�@>-��pzW��:�����x�*.9ow��``��C����?N�>�TNz�Q5̖P���J�u\��w^��Gx�Qx���T^F�o{Z���������8�Q(�3����O8�ؠ<�l�V�CY��F��=y�+���fc��G��@�#Ƽ �g�ցN�ɞ����0�>>��I$���f{HF��їI�����~�{Ϊ���&���P���9>����dub��ƽC����E��'G	uC���Ӣ����H��w���07і�D��<ф�eϋ��V�t7��Q1"b��/%� 4͖���e�Ov�9�m���l���`��x�4�0�T�}g6W[��/��B6t�7g;�%����2�#kW id\;��:Ž�K�kq)%�7&K���r�:Х�p���RV��9+kȏ�Mg���{ڴo�z�Җ�������!�j̍��K���)�Iګ�sI�켐W��l槕�C��RY����yU���`���l�F�N���^���w��6i{޷��&ob����b�����U��W���������}��*�E�R�ݸ3	w�%�m[��=*2{�U�����pjS%h� :15d\*�ܜ�u�s�� ��m�S�yT �pUs�}���5[��C�N��J�~w�y/�}ʛ�KZ�y)	���z�=�ޮ�������b����&�z9�����$���������ʮ+���_������7������*���w[����+�ǻ ���2�ےQ���X��Kƕ�g���1�ro�
���bդ������Ln}��\{�{('�!��Z���	��n�`"�N�W��fp�{�$}�A�A~����������{\�;�����Өw�P���PfbR��z���c�;5��.^�|vu��1~����,@z������}��H�L�;�.}͸�+�s]�gՂ�'Cjm��pN?f�����lE�_Y˿�дx�q��\����㹅�����Oo���3�`��1�����]+pb��^0SEɜ�WW��z���7Zn��r��[����}2��S�r�3�#VG��+Ŵ9J�������6�9;��l��'0nJE���5�Q֟���}9��;�Z�޽z�;������o�����.�.3�'����Hϥ����T�����|�F�*��O�>2��� 1פ��hw-ZZ�w�i��߉���U߬G��)��y~}ʜ�����[֮����,n�,R�����"�L��p7��X��N��J�N;$��ED���+]{�Ћ�ҩ��xR75��r��w��ކ2�wB��������O\/f����Z2a������0��55�r���#����\��[	_���oo�9�qO�CƖG��O��ڱ+ʑ�����~͔��t��J<�G�.>���]e4nO��9�_���j�2U{���js殢v�5�pg�_���R�b�
���(Y^Rw�)`�ۈ�xj�����d���oؼ�=�:�~>'k�̨wcNO!D��lVv���s�w�ޜɝ	��6&Xʁ3�I���)ȍ�`+����a��=�#�oъ�6�gzl�>ۦ�d;W���1q�*xݟ���2��,\Tϑ���Y��3/,ߎM�0L������W����v�$���a����5ݜ�i[�^�ly��,/;�m��R�Ӎ�p�7y[ö��b�Vы���V9���)��(;P
�,�[<���
��"��_3�L���0m:�Ѽi��8�<������t��GW\�w�w��/z�����+�({4'�B�Cꖕ�,���O��B�9x�m�U} ���s�ʘ;�,�#�}�ћ�3����}q���9��E�|�$���2|��z����`>ef�-���;�C�~���e�s��!�Q�R5̰���	�}{�on�=ڗy��Hvj$�ޯ[-k��DS򸛉��#�}9��{�t��&� W�/{6�ֹ��gă㐠�UD��-�������7�!��m�����c���1��U}�{q�GL�m��z��^2)̖jL7$d��4.):^=��z:�x�E8�Z�N��W}E�zgY/#ƣ`TC�Q5 j~u�!���H@���Fs�_Eg�W���~�sY��kU!������x�dxπ�d3q�T?e�5
Y=P�ǟ{=����3|A�F\Y�┷�������VGuǸ������:�7��P���i�g*�{&A0�.�7��'ՇRH>'�1�F\����>�)|o���dB~�E��Qqۨ��(p���eϴ��45��v���I����W�ˡ�{P?K�[݆�7�AMhV��mT"�3�1G%�W�\�h�64�.�]��}GT��S^�Fӓ�2�Ꝭ�w�f�{�S˭�����{Y������8��Q���G1CQ"S�G��or2�C�i{3�傍�p6t9Q�r6c�,T3����dyrZ�+�n��O�rb�s�S��}q��]������g�>;;s>�·q9G@�?�͍T���a��7p#ϴ�_��5����SY�gӬ�����w����ʝ7\<����?�z�3���Vy���o{����#L
���x��v�~�>��S�t���.5eO��R�3-�4���yD�љ�&�wн�Z]9�ƨB���b����|=��hxvK�B�}�	�g)<�W�1t�V�՝�ݼ=d�^��X�j���W*�͋��T7�<^�F���S��^�4׌�p���vW.�ld
&�����3�'��P�*e��ϖ]K7�X��n��#�#�����n9M=�Ό��������3�.�( yT`B+�s���c]Nx��z����c�>D߅��e<�n�(��]�K���#O{}Q9�a1rY�P@J��~��H�Ҽ�Lf:vk!^�>��R���V������}�lv��]��}Q8{��`�r�<Lg��5�d��nI�L�ƺۄq��Kz���
'�\�Wov%�$���;���{]�'�k��XM[R�i���.ž�;M������X�9�vȜ�(Jh��){��0^ ��_��=� ��䆉�J��%��l�Z���
7�$ͫes�۶�*&Y��7gB��tF�����=Q�������3��R'�Ӂ��zp�g�&���e_�q+8e8S�z��+uy!�+��W��r)O������y��mW���R�5��!��6W��^Ǒ4��3T�k���gђ�B�3>񿊜�:+c.��Q�R��?uǲ��zW��Q��5X��I���"�r�0�;�P�ed�����:ǧ��Zt\Ek�������?g��|��'2�$,���O��D>Q^�~�p'�޽���f���*0�[�����t\+u���_��d�XC��FR^�j�w�]�C��#>}���ʬO^��X�yS�C�f��n�8��,�ˊ�y=!�r�g�ki����<��W�����������H_ѷ�#-K'vc��I�Ŝ"Ď>B���G�i�U
rgN��2VF�`
�Ցj�7'�j��� ��m}���ԀÕSld����e��t@�d�az�W�nT/K��9d�r�κ�l�|͡��ȥ�<�w����x^��<.�I=Q2�� L�w3�1��K�~�	��x@xf�{��=�澕%X���J|k���2;�X�0;�6�/sAT���"����5�O���T���M?[��WKǢ��O�}��ܒ���|�l��7��;��V��띛L&Ƥ+@�άN�2m��,�@�e�]��lq�/R�Z��z���ʑ�uۉ-s�м?|�{�z�G�ґ�2��nH=Pe� �.*U/�YE����luxNU��ߵ�\�O��V��q�c}�Y�yT=م�%�|IU`H)3��RK��x	���d��)}�}���z�H��z2�����P���'M���;�rY��D-nƊ��G�������Z>� :�H㨼���j:��%}>��2���k�p�n=��q�%�5+�=��ٱU��m��*}��4\�_���-k��h��ޞ�K�X��k�T�9Òt!r6�Yۿ~����s�ә%�pj3�&"_�B�KGF�/��o����^���2�Eg~����c��g�@!���x	���sl�_"�MA���鱟K��F[�Ʋ#�>=�r=~��^��}֚��H�F^�����P���=@r�b?�:Zy�0���}�މ�*c��x,�^q�V�'s��o���Gz�C߮�=�R��|��ࡿw��>%l�}[7�vPU�Q��c��l��WS�j��|���m��bu^E��x�8�^	�q�mXUd������~E���{�k�K*!P���wql�k:OL��c����=Zv�kN䪑�i�$Ei��y���x9u�[��uK/a�p��0uU��5�{����2y.����(�S/e�E��*Ţ��%�(��6Ջ2�l1hs�v8o���%'�Ͷ����gH�u� N��H�94l��|z���O�����]%�J��ޤ6��N9���ML��mޜ;goctP}S�«���ʳ2���,�٩�P�40^U���z�xu��ueE������h�ڳY8TT;���g_5���X^���+�-�8y`��͕�{zu��ѥ��q!W*;�sa�/-E��+��sR��ow1\1إ��ʍ��6��\�ʹ����{\[X��q��l�,I�)<��"h���u�����L�����{o3��%�v�V�i�[��ئ�q���s�u*����èj�I_V2�}.\���k�=阒|�|�j l69�f�<\.m878Za+�75<V`���^9�Q�h�P�;!�<��s(Q��k)��ja�Rl���G�L���YÂ⥆�a���e�˞�C��&}��5;4ʠ�kB(<���]���-)�=Ӻ�)ZU��,
\���Xh&K6-5�Ӵ���u%mB ���Y��U6m�v۽��^p��{{���5xq�f��%3���ً^��9ʵ<��6�eN�`C���}�v��(%G7x�ͽ�
�ý����7�\�؎r7�k��VuH���<Ѕ����<=���I;�0�\b���/l��Y����Yw�j#,�ե`ޜ�4�>ś��e�L��C�Ժ���m����Q��=��ںO�J�D�t�Ǻ��9�/#�_8,CbRa-gD&�w̧�.��֔�\��}��:�<Nrs���C�HZӄ��2��lT�WWP�K%���Ϥ(޲^k�M�P��}R�ˎ��P���$��p�xq���!�6/���N�[f�;#��*إћsP���k����µZ���;E��M,��0>�}srr���M�S�ޮa��K���.^d����e��I-��ͼ�QTS��D�����v�x��Zz���
��1
YYC3k5���  +�٩ems]8���nc��M�.,��v�ڋ���|x\=���p���{[&�i�`9����4�Q���^v��b�u[��܄�������a&�ʨ�9$��&���v��0f�c���<��=q#CK]p%\����z��3ua�sL��Swh���{q>� �ۦ{��Bk(���5��\f�rvvǔD���<A��˒�2�9S�3��e��.�i>YLEgcO�2���
���@�Enp��=�u�9v^j	����(��6񻂮�����R�x��b�ya�C��#��I��a�/x�a�̾(iQ��u�fe��n��m�{F��r����b���G���*�77��g� ���;QW��z�}X@@�-EsJwSӚ�#��Xd�BEjZK�.�uUs����u��)�r���1�
Gu�W,�<�ʷws�k]����u�rH�r(2�jdT��BNaq"3���xQ^���KBI''v�TjE��E^�r����f�t�H�"]��W0��Y�
��G�r,�����%�%T��(̕Qv[��9��IH���7qwu��H<W\�8{�8TQ蛺����{��'��DR$"��(��W:��w<�wO:�R����3tY�y�wT�M�***�u�w]Ȋ�3p�ŤhJ#�9�G"�iwQ�Q��tr<S��NE��V����j����#s�"�ۣ�Eh���؄^J.�BE�')]�w�eU9�y���H���^w'*�%V�)�K�) j�h���!%-�S/r��'Q�9d�.�7�\٧��-u��Qp�K����tv�5r�z���B&+ O��vL��2a��'Y{q��ig�
�إ]���G�J��J�^�yH˝�uU�%zc_J���tG�w{=W��Z���ޒps�ը���4j�~`�?�*��ƥx�sf\
�^W�SO�����#����t$~s�w��'&�L~�7����:t�/�qS�:. ӡ�92�^�L�	��14|Ue��J3^�����]{Ǳڸ����Y��YS������,e|�bI�'[z��t��͋��k��|^��ǲ4��"�z�܏z��R��S�!�.���rK!����іl�V6��;=�Q)ВV}^������z�dF�'��D{������9���V.J9��h�5�ݜ�cn��\����f2 ja�Q�x��w�[��n��>��s�������Yw�.��z��Sk���= �9_9 r������x��j5ՍF_�D��z�9Ӟ+�z���ԖƟa����x̕�u��sL�C���A��Q-�q����Σq�R�P� ƺ�`���×q׶��Mq���Ȳs	�{޸���Ux�d�qT�w�������t�{ڟ/�q��Ӳ��W��[�b���٦��:]�1�|Jr�yD($���M��G ��o�]�]��Z	uց�QY�BRܧ#����W}6k�
�=��-��F4j�ͧK���V޳�:�#���f.먶�7��04���vv�+s�:��t�ܮQ�2k�����Bj�m�+�c#��g� �u��<j29���`Ho��� �6T��3]q�����j�>�>۟{��9����q����"<g�w���*��R������*���yr�!�|{**_�t�m�g����_G?u�g��o}@:~���\�ێS�r�՚�J���^W���:K����6vp+�V�/������ۅ�'�q��Qp{���ō99rէ\JŗC̽����(��a\@��6�]>'�}�/���ǽPa�o�uo���v��>zW�1��+�_�TN��Y�����8n���|?o�gC��r���ү��	��?k1�w�<�J�q��{��
e;`��\��z�ogz�ڹ�:�'v��ʁ>E��3}����{S3��z��:�i�}�ּdc���>��������m!z�����)N�n��{��✬7U��C��1��UL�9�}ƨB�-��Ss��������/-
�S~>��K�ҽ/�7�]Q�sp�%�������?��.g�[���}^ӑ��G�܍�Ǽ���@�yr��]��vɋ�L��p63�[�%dF{5��e�&�'t��c�UCf����J�
�y���뒈��':�����iS��YR��GY�Ϻt:��T��Q��4륧V�{�����%DB��Zۘ;n
���ɝ2ȩ;��OK���8?;���.�����,z�e�#ʡ�L�>.���n�M�sw�&��ѣ��h{��R/�g�3�wO�����\>�8˿��Q�*2���x�ql���<}bEމ�.w�nyn�2��N�h�������H���\N�ުf�.K5
	TA�<�!T�^�R��h�$��u9�:������Θ��7���MǷ����ꉨ�d�P���g��R�|No����涧�L���e�kY#E�'�lzQ>p=87��@��g�&��ї�#���y7��C�&w� �|o�䉕��7JZ=y�+��w��ۆ�������� 7֥9.�nz�fO�{Nk�5���E?/�����������<k�fNO���\{#�wtr���ȋn5i���:�ۤ�����[ؑTU��������=�mVo��jC��h�����
��S[�;�V���v�gϽ�7�z��R1z�ґ��lq�,n,�Z�/��:^(�|2��B��3k�K�/R���ᐝydd>��{�V'�}z,[���q�����{FK��P�"�u�����wog�+&�'<�e���"�Ճ�����f��R�v���ѼT����)��n����yc��P©��O+���Hz�/�^��p�q�"� l�i@���gY�.�5s�s�ָ�n����6��:���v���⦊ģ�&;�V��f�h;��� ��<��!�z��~��N<��q�d���d�(V+�N\��q;Oa/b�w<f;na���_��i�+VE��Srr�j�M��є�i:F�
�G��[=��7�$����ܻ�(	�ȏDj����P�@w��W��N_����s]�2�x�j��D�=��b��.U#���Z�,�iB	��eP���)��"\�~�{�i��g�F
S}C׼�j�vF���~�x����p5�~G��7��X�>E�*W�1t�c�xc̚���^,�)*�=�^z=LnG��=q�;�p7���F��%�<6�t�?G(���B���S$z	֦��P}t�p�r߯F|���V��i���HN��N�����Q����ڷ��ȉK&�n�"����3N:d�����s��~Wq>��2���l?W&���n(:�}�)���O���}�̟MB sG�Dķ\�:Z>�f�Q�֍G_П���Ӝ}�i�OjD�n(��}9+��{��u�s�Y$�vKf�=$LK�!W��ö��{�j5�x��q�!�LTb9���^����M�˜��v*5[�J��nl�c�X"E������]��q�]:�~��d{ծ���,G��G*�(�b��8ȧ
�8m��a<��v���TR�r��f9w!h+2t[���[���Xb�oo5I|k\��u�(m�\�)�&>���T1�H����h�p�w��"��sl��=;f�V
�\����K�!v8z�:u���3�z���GV̅�~Wtay���>���j6+��d�E��2a���^�9���"pKS�*w���G��>7�>��ކ1�]�{��D?O�����E���� ��>%G���4:�Rj�>Q�3}uW^��p�_-��Å��{~�W�}�5��x'���VO{~D�����Fz#���:wj���R��:��ܮ�C��q8�Q�M���o3ׂaP�yr㾉~����Iˎ�����ng���^%%���Ƕ��oqH���G���\�L�>���e{ΣyB��7��Ĵw�p�ᎂPu�_��t_��k!S�ˏl��pg�����⯁�^���r=u��v�;�޽f/�YSŏ��J+�*_��B5*���W�3��R>�ty�V}���F8���ޯx�T��Fo�TB�F��$���\�^��;�J�-���>�9\$�Fz���ǝ`��'��Hz��c�r''�l4���~����w6T�4�p��ȭ-a;�0)�߰��
G�����]`2��5��R�\#��{�`��η���f�2�e}��K��8Y�Ĭ��	S�}E2a�vu�x(�6�Oq=���;�;�oKơ��S��M�Dw%:w(*�m�3ḋ5>�]�����j�[ '��0��ll@^X)����n��!zG��G��|J��t�z�_(D��Y�}��Ϋ��6J���<���n��:[/5ՍG>��q7>��}��I�^S)�	�4��|缴��p���m��f�̂�(!_D����끸/ō�qg�"��v�Y�voj�'���%;L���6_�ӺM�޸��ό�IeB���Q%yM
�����������9��ø�+����0��ώN2^x�dNbP.N��!���3s]6Yv�C݆=�N�Q�]��_y܏�y]и�u�}�3�;��ƁO�r����j��x�4��s���pVTT�V�͹L�wT=+���3�ut^�@t���q��o}N�=��v-���od�Z�,�Q�R����,"߱{U�q��X���1�e`�׷<�u�6����'m-�=�7�,jK
�·qY^�_����磻4��_Yh�%g7�ogѾ�T�q�O�]����u~�{��m��h����χ�ӡ�NQ�_��>���]S�m�i�.,�q.�����Y%�0�{?7�ranXUU˙�Y�v:7��H��N"R���xB����kl���fi�q�P�R�ϊ�07ݗ������6�sn�z.^.u�ݵK2)�=w�vs�z����H'#'f�pӛ;��b���ۍdxd:���;^�eg�V7�ը�ʝ6�'v�3.+�b:��غ��ҳ��xP�d��N�k4׀�N׌�O��_�����C���������S�-E���c��ᦱI7@³�.���R7����T!\anȿ�Jn{}���z��|�}{�~���+���1��Ԏ���<H~9eT9��WK�Y�����q�{N}�����}_��������?s~�������Qy��T��O��U�e��ϖ]K2�З��\;����nؾ�5�����9�,��U��m�������`O�J�-��=}"��_'JvA�q�J������'޴4g���h��ë�o�'o�U3�\�iA*���$�I��ӽ���ܑ㳭N�s�\k���'�v�|}�lv�Wq7���鸏W�%�Y{t�J꫚������@��	�bbs���G\�_lQ��Z�-?;`{҉󏇧&���h��g�$8r|+��ͻ[]]���dʙV�f�I���R��^r�~=�f1��Q����@�yǣ�]�]��{��m��N���]��Fr��5	�傈)��j=G��򡹤uCST��m���+<4%ڥ�M�LsvKU�;���Qt�]3A�ԓz������h䮩$ݍm��x�D4���=����i,����v>앩�]Q-Z\���5�S�������f_�F�K��W�KǨ�)|o����'l�g���KR+�|ͯuv�Dѿ{�{>f�Wdɮ�g�aC� zp9+N��}~�y%�8�O����P=<}����/z������z߁|��Mʑ�֞�%����mhs~�漮G=��s�m-�>2xz:�2{;���ݷz<1:��}��OʬO\o�E�W3g>���B�!f�5�ic�j�z�з�q�묥��׫A��l[�W��}Z̨~����:��r;�H��2��q7ƌ���Z��ޑ��,��a�LyVUi�5/Ĭ�4����jK�u�g�=g�=�	�N/9~O����|�ڵ�Y#�:�Q>c*��\�?fpU�_�Ϻg��O������5��{.+�Y\�w�?v\{�z�F��ZT��_I'�C�&x;��)���B\��y�<:.�۝=w�w�W��C;�;�U n1��zq�}���=���{�v��e�0�bnx@[�u'�7nA��r���ܞ>���q����;��cr#�E����q젞��I�Z�j�Kw%�P�
��5J,q<x૿�t�6���W���+�����3}v`L^�j��j<o��Ί����c[����v�4���&�L�{QBr��e]��W��_WM��2V�Ǒ]�*�t�����'e�+DT�ǵ6�)��j	�b�
�O3�)����<��6H���p��]7�$_�-��b�י[�z��HN��N������*��ֻ�Q�q7A��뉿�J�{��j7��&��X�ey���ĥ'& �3���n��<�Wm�o�?C������ 揤��n��t�}�Lb*5�Q֟���z���Q7Xv���O>��}����z�s�Y$�D�ʃ�DĿR*Z:7����lFh�
W��3��:}йڣ~���<s��|�`��"�zj �����.{ƃ�Zjt�{6�qp0��/;څ署�s���ީ�y]ы�y������|�F�}��2J��0����ٸs�t'>A�Z�݆���W��t��� ���y�:�~�=k٢������q'%T
�n�"=L���{������z�M��q�؄�Å�m��d'U�s�ޡ�K#�x'���l�����U�J��g�����m�H�R���l��;��#pj^��Q~.;m_�:���ό3�~��4Fz���S�M����:�{\�\�!�XѪ��:EeW5+ģ�lˁ��U7�x�S��<���#Y\Fy��j]��j�6���pκŅa�Cx�۷j�?�7���d9�����,��X�;��%\�V9�����HQ���ǁ���w�9�x�	�)����9�i�|�Fԗ3����J�;:����Ƒth>��1��E��$��g�_����v�<�ϣ�w�z�s:6��ۉ�a(:��3�G}�*W��WcL�cM��xYa��`z���7	���9�x�;W���1z�����)\cY�}�7.��*/�jg���V����Ӑ�Q��a����ǩ��z���Hyg�f��.ʔw�#g�r�1d��ζ�Y&|f��=H]L�n��
��,�<}�џo�|��{�����l{������>W�˝��͌�8j#�ĕFc����2�O:���M���Kw�9�<糲lG�D�����`��������ꑷ��w��H�jKCu�lt�^����~W*�E����z��V�������'�o�Fߦ��H,�U� �<@�~,nclM0Ɇc�A�K=KTc>��!�ަ�8>ζ���ӺM�޸���W���̖j!T�q�C��	����d:��}����懶�^g�z|=q�W#SU�È>����K���P0ç�>�� 0��Zw=�7#}����',�N]���oL7��b۪�_4����\B��?G�}�m��m�m�ᱶ����M����m�m����1��Sm�cm��m�cm���m�m�m�cm��m�cm�cm�cm���`����1��������l����1���`���������m�o�m�m��m�m��������PVI��V��#�rv` ����������ꎚi*�EIU)E( �!$REJ
�
��E�T� �))( 
	*�$HQR�!���6m�6��j�m�����J��ۭ�ܮ��{׎tѴ�]�+n�v�c���	w:�͓s��խ�c]��SM�nܶ:;��1ۺP�ݽ�����]�ު���w*�(��ĪZʶkt���+���m���թ2kT�v���5i��l��ٝ��TV;���ak4u�cH�2�nf�QUD�s��nv�㓴�K7]��  ���$�����V�lh�6w�zz[T��=w�U=��kn�<��My�]��[��u��T{e�������=�����˷�wc݀n��������-�:n�N-�  ��*�������@s�ݵ�uPv��=��>  |q��
��E����   ��c�(��(�����   �>���4h ���7 4QEQ}�^�6Ɉj�Y��Yu���|   {��`���[s\�T5��x�՘�����
UW;������w=zPm��=ǥ�뢺�w��4{���z�y����=wn�w4�3{p�4�[�wm�Z�  k�
�_53�f0��w�������:���L�����P�כ�J�׶���B��n)�M:�6זz����45�5]h�h"�;n�f��1zӕevc�  -{�n��J뫸\�쭶�n������M�Nn�^�u�t�����n��K=�V���:��z���xz�:�w��@���5�ӪS zn^{�˭���իnu��V�6�|  ;��k鮴�s�w��+F���ָ�ڀhA��O]�ڔ�W���+.�潶[������YzY�k�oW��/m0� �u{�^��u-*�UT�*�-�n�U�X���Zm|  �> t]�c��w��az^��ȥ({���^�ݎ�����GB�fu����R�0�=ty����xW���7�g���ꁦ��@{�o\^���gv��&��;��cj��|  5�C_U�������P�����V�Ӻ�n�
z�ޮ�@�
:�L .�i5����]hWV=�ڲ4{��nkq��Z�E�������l-���.�e��V�ֻm�  }����yqu�=wm�۝k��2������ Y�<��h���s�{תV���<s�� �틽{�d�� �w{�Wil�H{�v����h]�G:�e�32�&
��  -�eMS/�n��5v7ws�z� �ޛ�zSK�7�c�Ez]v�W ;b�۳מ=���v私�z�N��������lw`4[�T��̪J�z Oh�JR�  S�6LUR�3Pd�JUM4�&COe6�*�~�   �ISѦU$��bhzj~�������s����.<�?�Ğ ��y����WI���}�ε����D$�	'5��$�	&B!!��IO��$�܄��$I! ����\��^����|_�ן�e]�aw���a
蒨Y!����cvp`�u�i��ӖkH$*�(D�Su�k5ӭ�'��-�*Y�ſ�/-Bm�,�HMj䦵�O���]'7ScA�v2�L����/-k���O��d��!�J46enlBj���%�-��C��цar������GF��p������n;�v�)d�Q���E�͕�K�>r��m&�#$OY7Vr�n��`�.ղF��ǔ�0�� �
o
������,�ϧ>��w��+����ٖH�����5)�ݻY#�s�rd�m��T���M��P����7bX�8�-{U��������4�ȩ&9VQ�h�+^i&;�wn"XØ1��R��v�xE�(L���b�vn�ڡ{�L���Y0F���V���Z��4R h�Õ�1�H&5�%]�fLw��G��|� _�0w��.�<׻�^^�֌��X;5f�ʲ�R��#A���F�.K29o2&��10�2�.VIK
f�ݱF�Ind����.�n;d2]�i�ѕ�ÿ3�r#6� �����;��-b;����;��wQ�V�$�\'��i��
�[J� ��B�hƦ�A� ��կV��'wZ֭S����7S���.%�8����Ƌ�LCe���(!!����� ���6�G2���uop[���h�ɚ����6Id!����D��޸bڂ��hDn�{�C[yH͠��T�]ʹ�^Ҽ,�,�R0��V��Ԧ�x)�ںu	.�Z"��p\���&������ڳ{���&�	Y��P��H'J��t�6'VXR�7G��cMR$cu�VdY�	k�nkM�,�Vp���ѻ��� ���ʁ�
y��&�	��+(�෌S��S�@b��Ŏ*E�k �b�EV5����h�[3�*Yz�f����77`c(���t�W(f
��n �d��-��Hu���n�@���&*hh۲ݚ�)PV�lc˻�0e�P�F&�8�piفkH�sUh��k#٭�ulX@6A�7�vVL`e���a�k2�&�lmč�uM��7�ћ�f\R�coi'[W�Ȧ�K+A4T����Vױ�zL�c�\��Uq/S�F:�Pi��
��:�if8�P�$.#�2��kmJyJM5�+[�U�B���CMj��b�S5pU���M:�D*�y(9�Z�su�1����#xyOMn�^�hҕt�ډ-9��Q܏L7��ٲ�ѭU��M���NVAcp̹�B
��Mb�����Kb�k%��z�k�,]�Ձ�(+1�2ĺZT��Dcz.�t�Eb�E�����ɂ��[LYT(��GV��d�ʨ��+W�>,���)4���]\Jiv*y�Cvh<-��k%!�� ���!	ٚ����v��#�������4ܩv�0TN�;�r�K�7��&K9�XM)a��Kb�n=C�1�zkE�GUe]�
�����o`��R�y�Z2��1���W����8�Vc�i5a����R��`�t^S)��^+n�[]	*𚴩47�Lø�����Kݙ>9G�[
[R�!�iis%B�xٸ]ڳE9���*B��n�)\Ym�������4�mh���S ROo��ɉ-����].���t��c�4�K*�z�Jҁ1Z�%-וd��cl��`$k]�#�w��r�JbWtp;�.�"jŬ�i�j�dU��F"7�(
�H+]1d�y2Ŗb�J+�wFGr�[zq�C)*ŵh[؅��U��M��T&�w�.����@/v�.�]n0���+��{EA�`Ȁ�c/ҧ���cM�����c>�9�l�i�k�긞��(��@�b�zvf'��4�'@��)�c�ӭ��&�k��k�Sk!
���-d� �tCV�drv���Ѻٍ6J�h^�&
�,ANE�-J�H��L(�;���E�f�*&.нO�eLQ:«
5����� f�Gu5ި�vA�le������2Mхi)й�J�g �[�Ҳ�����{K��esoE����b����iT7+��90̑�*�Mb4��n;V�e`FV"���	Zk��fdn���%7X�R��ĦU<n�ي�i��6�҂�V��-9#:U5�oE��ZV�)nX�#�Zΰ�[�Rh�.��#��:�ΰXͫ�lfd&�ݸ�ljձS�K,���Qj�S�h3"\�t)�n���Pv������E�X��A�ŗ�h�{�ʼ7����UnnV����j�kA!��:� O�Y(�^�B�))��.�RCkN��b �Z��s3W׳)PG\WLЍm9f�J�<��^��	JҎ���t�&��ԝ�5��N�Ue��V�A�_���S�hf/��mmAA.e�U�e�xi�a�B�Zۢ��$�ow�!���g�fKR];�۰j�	aÒ��318-�B�Jx����Ӯ����`�נ,�(�j�@2�F�M	
q��&�S�p]��ysq��]���6�	�PCX�2)���v�7�#��B#U���rnVZ��`�^%o_�o@��q֝���z�Y[�n�y[�Z�JI`�A
LS4ZюxݘJZ	`"�}x�Z�7�����t�m�H�lS0�M�1�ص��9���n �HV���"��X�"/F\�Z���,;��:���da�4c�*�k3@?X�E�[nly(1�����PJ�;�v h3f�}��҆�i���[)�r5�nT�7��f���S�e�[���l�6Z^�9&�^l�A��T�K��O`U�*m�:�.�3�dwZ��n����(]�FiJ!�R�):��`�U��o�Qj�Q���f�������i��6em�W�g���F�́T����0�e
m�{v+\͎����ZGD\��$�k-��TOt9Aʛ��<Ì��KU[�h�#	۫mY���2�S%�#vn��n���C,���oq�t���wJ�j�6*�Q�#�ľ)]�u-�g�v����7��SM#6U�l�m&�t`��a��HE����^���u�Zv$�ֹ����0,�
�Q�{Yw{y�U(�Vv�[ځ��A�(��U+V?�v�[�RPi���1 ��%�]��A�2J��S.H���b��1�Y�F],bjw7ER�P�1J�v$n[R��oi�X�a����m���I�&�l�SJ��Tc/�+��Jݺh���Q�j3(�T`�@S�BV]d�7v�Ԕ�vH�ͥdZ���,�qM;�m�	���a4MEW�X�%DZU�4�:.#aǖc� w(!9[��r��DpX��6�E^��M�¨�m<�K:)*�.lX�Z)ekT���)����eL�j�Ux�X�m�t��-U���:l5��*l�5�Ft�$8�T�R���yL�������m]��V�9�d�;7]�S;vec��RS�Gی���Y�h�F�R'6i��x����N�Q�=���H颵:�1�e��M�Z��1��VM,�E���V'I�Ɲ��^������,�lӳ�]��,��)b��B7�n�xJ{�䶶9���靾JO��l �� e�&s�m��7�����"�RX��@PE'A��gE���$��U�bum�"V]f:���H���S(-��C]1�dД�+
����wg6T#5d�n2�yz�R�]bd����x��߮�M��HS:�^ib�OVj;�`�7��qT�WRd"�|����dJek�Z��wAk&87 'Fwr"�Q@Wq]ˀ#�� D��c�Kц�Y{4�+��`���ʚ֛5��D[�b����QPlg�9u�i-��pJ9��ñ�X{���n�L��Z�����+_dnj�u���LU�Q���p���saq��w6��oK�lA4(�]Yh��ofD�n��[�Y��<��DF�^��U�uf���9��].����8/iU�E�:U�٬�m�t��`ձ�v�<��G�ՠ�ܙ�o)�*k���cv���!S[m̧v#�伱{��+4��yA�x�����L�&K���8%�/T�n��ӄ�)ګ�ՙlB�au���y�êօ�Q0�T�M�a���C%��K䚎���Z]���
SVͽN���Y�q �Z���k��֝-�qfa�۔,e���S��Քb���ٍc���Y�@3T��@
)V�����m�U���t��4�MKuaߛ��Mԋ�`ͧ+eh��zgf�MX�Z͗g@we"�5i6���##fL��Z�E�D�Ja�B�d�A��M���w,H,n/�!LOYe��2^n�z�8f�"̽��d�~?^ŬZ�h���kfS�6�ފ��v��ыZʴ�;���D�X���ͺV^���1�U��EJ �4cl����!�.�Z��	%PT�3�d�g댕h�:��Gۤ,Ӫi��P|�)�8(Q{F���&2<���6�F�h�M�ZՊ��h�!�0�B�;J�����e@�rJ9uQ�ɷ�\��.^���7J*��������j(H�E�y.��v���:�y�h�p*�]--ޥ%F�0ĕwm(��M�[VR��O	�R&`L���֚9�(������mM߀��9����,a7�1|�<0��5��P�Q$Z�{t�f�EGm���TS��fSٷv�}����kAB��rbC5;��V��Ք�In�
Xԥm�,Э	�Ae˽��~ȩ�μ��b�PL%b�wRY�֐Fd��kwJ�������Z��,��_�<����0�vBT�v�X���.M5N���]��u-H�bMHn-�*{��f���zt٨�ch,#2��n�+#�����r�͸�՛�@̻�y)KɄ^t�ۚ���dv�Y�"�!_K�rֱ�b�ܙ��S�6j�rnٙ��N�t���i��(K$m����b�Z%�\h�vڻ
4�e���n0Y+5��-��1E���*�]�QL5��P9�d���)��1�w�Z���pVE ��Y	������i 83NR�PK�jb���"�'p,f���E��k�Pp�����\�{k!��<HEd�������:�e[m���|���)�e��-l�C+uٺB��Dֱ�@a�B���T5km(-��RSz��TjY��1ɚ�H�C��V&;�V��IR�� �4� �@2��6��0ڥq-x�QN�.���a����*��*�FA�6�nC.�Ce�Lћ)�#2�,�j�Z��5>9�Tiji� 屙p�;��=B
�W*J�R:���Kwwp�����"�n�2m^:ؙ%f�{�Q�[M"z6�5���k&:�J���6���H������Qٕ��mb'ARו��vȚ2�a�4� @��3�Rm�$���Ii�U��,�36�̃/6�5�{B�b�ІQ���ݻ���
�.6���)J�$��-h�$���xɘ�Lт�K{��V��x�ݢcJ�5Q����F�e-4��c�ඝc$�dWoZI�p�.]�69���u�M8���Ǌ��4	5kl͵��tQ�@V�!▚9�a5pj8.�UܷZpm��`�Sw�U���7������2mk	t+Ub�@,�,��Q/u^��]lo(�r♕K阵i$J%�2�-��N��������X�i�x�軪4'ef�P5����꩹>�~�����+Bb53a���]��p	w�a�D����5�L�Z��J��%�ۿ�c/h=�5�k�p���`f
�e���r�QfdT�����j� ������EHI��	\	+U�LY����۽;l<h��uG�W0v�h�f֖�Cu��*l@�&ۻn֝iZ�q�v��:V꫙g2�4�i�=ȓ��ej,�%�e�r�(3�J��˥4��J�����B�
����FD(N�JTK7T`T�Z����ݽ��Kw��J�N�1�cqIt��M%H�/u\�b���/2��7��;b(���eL����+a��@1JJ��*�:BՕ��34f�{Vҭb��\�[�Juf�9�
O(����z�݊��2�V<u(A�a��Rf��E2�Kj�1sE���%+�T#KsE�e���6�����n���h�.��P+��"�-�0��kʄ��љ���0��+�Ě�wXx
;�"K�kT��1�ڦ H�V�M�b:oV2�]]�b�A�,�Xi,1[d롭T��t.b�5�\�a�i�Nӫ�6�Yk2��SE!�х����[�5VZ��X9@�ZP闬]Yf����l��9L�a�˥uRl�Cd �����i��gm�g-[�Yr�&d�X�2ԻF�Y��=�F��֬ݭ�]�bȅi�v��u0�V�@�Y2K�dj� ��J��α���:ԁ%���VTq����:ĕ��8qT��Kɻ�oY#Q�N�b��n�+��
�:4����rY7s^ b��(�w�v��.�m3�NJ4���?�X���{��(ޝ��S#6�����pk�`��_]؜*[�R�O$�Z7q欱(���۷P�Y�L9k+t�=�Zi�a2�ƲY�5�c�\�̩e����饭���x��-F�75��I��	0�\ܼ��NV,��� wXYt�°��u��p���/���a�&4(���ũ�Xe�kd����e3#K&4��i��5��ka�1���#n\&��O�(�d#[x�Q'�5Vh��l>�ֵ9l�3����a���E�D�J85A0�5;��v����
����uq=����렿'��5��w�YP~�(Y3@�^��H�E�)�`��,�rvN�ߴR��y��zO%�w^��<��m�R'�\�WXh��ە>����*�q�j��\>Z.T}q���� ��;����&֫}�!Ԛ���Ɩg*�?���A��`
3S���SrHm�Uj]�דܖ���}o-�rHh�sQN�ӱ�o�����j�y�;��v^��l<ͮ�aR�<�C�=�3:���ބ�#�P�ԯ�fv7q&9J�azC�0�VU)>��Jj��\t+k�h����W��X��zf�u�aKܓ8Kzvms�1D���*E�[|�l�V-o��s�����hw,��WZ��ʾ R�v�Kub���F�����1�b�����������I�%�b'�%t�^���퐜�"�����O9��B�Z2��ġ���F��c���+3.�9��!m��M�_]�c������Y:�:�B)X� �3��f^�u/�HTP��m��7���S�)�уH`�(ޔ�n宦%�c�����m�G�d��i�� �#��;�}6��R�q�wuv�w��m5`.��ɵf�!��B�u����-�N�����s������R�]���Y)�}����"��XGg�OT]NX�S�ʐCI�B�B���M@�O��'����Y��k=]ъJ�	ڵ-�G��f�X{'F���+Θ�N�oy�ƪa:z!IPX ;�u��rE7�n�v�}X�ǝ���B��Q'MOY٭S}����穳l��\�u�+��M���;|�,�\�>/�U�Z�w;|���qE�W)�;;ט�P`]4S��@㩊�V�ż��Q���)���/�3K�}Qz�R(��˝��Hf�ݻ��f@V�ʴ��g:㻾j���K�-�F]�Y6�\��+�<�ѷ�$ĐV�gu�]J�f� agqc�s���d�5�w	����Vb�S4c�o	���"���-��.-1���֍���b���w���!˝9�a�ObҺ��c(Q	Z�	�8����ٗ��8�kZ�*�]�:����R��:�5��N*��d��ً�a�"�Q�o�z�(\p;��o%U��w2h|���0��&V:�*��9��-�+N�Ap�El���w$ru����.Y�e�#�7�`��^��W�VM����{�T]q|�Gv��^V�@�U_-+a��aɚ�UY�)��%i�����4��iэf���+U�S����ʳ𦬻ځ��"w�y>�r��!�6�ZGM1'6�L��L[[����Q1�k�/'��#�����-���Zz��}��-i�f]Z�xż��������Av��`ZF	�zv��*��SUxh~y���r�f
��Z1���U�:�R����"�ﶦ�5�8Ό�!=��kYq�5}��z��R\%LjI��N�s��G9;G��Uq!��F�}u�B���*�!�����W�=�N�al�6C��iѢ�kn�ћ��N�&�3&ov"�j;�P����Ɍݎ�.�<{=�N ���N�r���4^S���l������E*�W��%m�<���y�j�W0�,�*��Qԯ���2�}��R��0�LZ*�Ci�*,n���:���H=�hk��Ven�WB�6Z�r��Z^2�tJ��`�z��q3S�[ㆬ��+���j��L�3jU��V:9�+zv�8š9�����V:�m�o�4�n�v�#�Hɔ1���]���l�q�&��y�hc�m
F�Uv��tȶoVe�������������x��C��Z�h�#��`�}%-�#�a�LL$m�a� ^YnZ�0�f� �ȸuW�P������Ƀ4�����s�V�����)���]��	k�&=ۙSm��GCP�>����z��/�cZ���x;�U%�-� م����U�uև�R|ƌ	m�w�b����l-�SQ��ں�p�6���=������޻5�Rr�+Z0Q�Y6�[@�6-V�m���ݘ������S�w��ҏH�:�C\1�J�׼�f���9kb�}�\A�g<��z��Ʈ���e�zBA��A��V��Z1�b�k4���n�}���M�2%��MJN���eA�$���jk����Oq��C�H-' �o���uk�,Q���4�3j}4�����㬂>���f��Pb�;iQ^o�"�7��35��g�@޻��nqY�H�#悹�(溵�XKJ�z�Cr�T/
vq��;1iq����F���[8��k��q��
 �_�}SUIG�o~î��M���N�d.�O$^u��]�"��|Q�}�)��tTu:>t�\�s�^�Ox�p���2�m���̎֜b�{�b���p��\��;T/��0d��z��}|�齅�:�"�������݈�*E�s>��^\@��~wun��%�x4a��:�+�O2/.uF8/,�A���)e4FkI�+�:�-y]�I*�����Ng�u|��4�:"I����rg]�j��:�`�ȕ�Wx�/'�2gE��0W���%��]ɔtřR&r\1馴9�K,ooov��Na#V<Y�l�B9v��ة����}3.�����KFs�K��mu�����fU�&�ܛ��l�:���9���QÖ����\���ly�]�ogj�������2�!�A��.��<���c4͂|���՝��㥧.G��2�k�$C�����7�7����k�s�z4�wA�5xH��4�4C�y
�Y�p�G��N�V�K�b�< >0܊� `����ÿM����)q{钕�l��.)1r���*ڶC����Vī�x�Z�5��Ïr3:�뢅ɾ�]N�͡�R����=�J��X�޷{]�f
m�"��/[s_i���|1����6>�F��H�j�ӹu/�!i\�&8�b�w�wU�*6�]"�Ձ,�^���n���7�<�v�X��K���1��8k��X�v���MC�Fg�w��q=h�l�-�C���B(��y�%�J�O�Zv�sq�u=�'�p���Z��������N:2���OC��rБ�af�-.�F��{:��U	$w���Mۓ�g`6�{��&!��t��{^��Y��䴲^��}�����g����a���݆�B��>ׯ�V79��23�]e����|��>�i��#�����;%i�¦OQ���j�M�F���/s�5���*m����ci���Mj,>�f���dB��cU�݂�63˟�JuN��C�op�p����ǩ<횳k1��)8.�1�H�B,�[5���vk��� u��XD�G���j�)�(���v��J
"�`�~�;cjv�Þ��٧8�N���N
U���NjX�u�Uvc���c=��T��v�.M=NΧV�g"��:��WK膮o&�C�����v۬��A&�]·	t�3;B�J*1�A�w���ƹ�0!he˛{��iRQ)�.�]$�l�ܷ���,����It�2�#���n����by�>�,#����;�v>���]���7��s����m`�NG���,�h�<���:�H�z����%7Z!��F�kSG:��J�ݏ���M�O���j�ӡ׫L�V���s��������i�n,�&b��H���Ì3��J�y��y�M�3ާ�=���^{��0S�ː�B�9c�gޅ����[MZ�����=&<T���/��{zl�ޒ�����:c���6&��]�����xS��=��ՠ�]v`Ȩ�!�W���U���+S�.0��+��BI]-E��7�z��E�5��huɕIx<-�?�����n_fG"Syd�gkee�s x�)�?I������j̖��D��뎆�����$l�I1�:����Qp�734�@JJ�꘨�C�=F�7�c7+��e��������J�(�[��A��[�㷜բZ�Xv���>f
1��>]x�oݰ�qy(���rP����G;t�U8Vh6���b�W(��64�<����)6z�N���p�Q!�Liu)�8���ƭ8,�:��G��JrGN^�㛚�LqQ��/��e��ԭ�ؾ�G��]$["R
A3��R �Ҧ���!��o�����'ѐH��s�[ʮ��]8��n�w4����]�I���oe�o[���ڈ��|z��w��%G�A#���4� ��k%�[f8��y�|��TE�:�I-t.���@����O�Y[����ύ�F�+,"(C�ʎw1�Yڽa�,�� ���/�3E�Ƿ2�DH���9��� �w3o]�^�Dl���&����q�	N�ͼS!
���MҌzݑV�"������/�������=�gym�r�-WS�N�V��T�5��`���ӝlh\#m�o��)kA��sB���j�˦�:w+:�mR�<HL�꒭%�> 팊T2h���6
5�z�g�p���ueh�I�Tw8>�-\��³�7Ӭ�l������,�U���J��F�h�S��C��2w�o�;jh֙�o�P�f�K��3��Tn>3^�7a*nF��OX�@� ��D��屖����H�vS�Ҋ�����Ȝ��t�:'�\Ѻ��2�����y���*�)��B���d8f����ql�1�11G�.��)ň)�dm��6VÌ�NS�+�[E5��X�����ZѤ�A��bCwgy�{$��|g3noT�2���YM���[� FڜD̢���JI��ە4VoVJ"u�9�MU����kL{/v�̀�#����h�*v�l[��ٳ�\�t�AT�rG��.�{�l��K��D�ޝY}n�冄H�2��w|�\pb.]
��P�������Id�0V�w<]^qI��x;!��+�+W%Ĩ�!.�*-V��7�jC�xNq��S�N������5d�.�����̻�>�5ۊ��m���v���\	ٰ5|���ޜ4�+\�X��!|�-z��c����ћ=��z-D_��u'����G��S\�����6�wZ�|!���7oC��7��������;��.no4��8ʬ4� �Z�Ξ��ĿWD�6�@���q5x����Թ�{���|�������<>�wJ�_�G��E��x�����;;��W�V1�I��/n���qi�-��]σ1GلK��n�b�o��u�N�^L�Wh�G�;G�ݺ �1T!	�@�J�M,�t�E�P�ݰG����������� �{"�=G�V8��
3��)����}��׀�(,&ИU�N_z|�����6PP� Ԉ�g�Y_��a��}.SWWO:�Ձ���n[��#���.T�l9�(����y�� {�c���ڥ�|'��xh��ϛ8!� X3���Fj�kv�ݯد^��,��ϫW V�!���aS7���<9����1P[qofFV��Pm����|w�����~�j����!~7Y]�=E-�]���`L�^�M[�q�v=���C7=	u���)�a6��帤���'�*�-r�>y2�fY�L�y{1�Ml�.��2��78�c�u;Pkj.*�����{j�]�+zrT�_�ߘa!�����4n�~F�R�l�cl��۸}۹Wh��V�1��{q�ֲ��S��m�$�i�WB�C�m{o��E�`-ǽ�ܫ���ܝ��bu\�Z���m�7Vu p�Sl��-�`gm:n1���B�uL�',�u�[�s��	����چV�"J��3��Њ3PҌ�)��N5}�n�8QG9��9X��'�h]ip��m��?UV���G��v���.��/���4����wxgX��l���[^[����m�ۋ7%f������G��o�$ /f�y�HI�7����a����tS� �ٗ �f��8���	�w�"�Ɏ)K�'�R���r{�ٳ��w�e����x�#+9֐5%���Z�C��it���oR�}u�b4��*�e.)�9���mg�}Z>Gϓ o��P^V����϶��vNL��:i�vN�Z84�;����.{���[BI�f?n��Ʃ7�[���,L0��K�E���LU�;^�e��S���ͦ��y[�s�՚Y�ڊ�e��]D�^դT�WB��@�ԫYC�*{+� �����Aщ-Y�:��7��ge7&�+h��%ͯ@\y�!�ղW����kn�by}W�^3��e>�ʹ�r�JpX��m�9��Ԙg?6��Wf�%H��\.m�y]2��݄)�1M�F-����w�VB���㬭����''U��h�V�1Ӭ��A��� l��i٘a�a��*��#[�o]��
��u-��Wʰ��IE򃐙��C��%��X�q�f.e=�G�I��3�JiY�@n�Ջku�3�-ؤ���2��Ź5�����M���}I����~!d���v�Y�H���r��!y�n�Ξ���j��)���B�G�Q�J%�ղl�.gq|K1��t��Yܸ�I}lkVՅ�Z�k�a�r�g���z7DUw�Ag�V�F��M��v��+ߵ�n����0���v]���4Wڍ���7�|�,.5I.Hw z��=Q+�us�YP���N ;+Fѣ�q�|��ӅAr9����8�>$�ͮ3�V���a��m+��<����oj�-W���Th�O:/}���AP5���C�椟o~y��$�BC�!$ I7��{��Z���~�ՊF~�h�as��n�kn {4'Ap� ��c���a�S@����Db7C\����[���[0�ޚ�z���Q������J�g�y��]e��e�gm���[�	�aHR�W��ݗ���*����m����&�T��|�.�u���Pǚ%��h��Ս5+:��5��1��j���7՗|�![��6ma���0��Ã�y���ܴ�x9����bf��sݚf�a�t�
��OMۉ�YC^��{�j�a������{����GC7�lL�y����:�#���(�9��WSv��P��M8k.�<�4Ff�X����Ղa���쥛a�����.�n�ˏ-���ؙ�V.��Y2�)�^�ޞP����z�[�o�]����ͅ9^)��T���U�� ң�u�qS�ӻ#i6�sP�w[��Jsa$p4�w{>��*���󳚷sZ��K�yC��P*�v������Y�d㺘�]v�[��e^豂d��r�~�qR��l,/�w4�X^96d��Y�Z<��o<��rk&��x9Ϭ�w�
ͱד	4^��w���[�>飋'���z�j�P�u}�Vˬx9�Wݗ������k\�#9���vS&of���o#�ՊyF,d2�"����]�V�8r�I�k|W�1�)&e������}��_{ Z�ŋ�k�s�@�����Uc~����WǷ==wt�^�[�Q�mX2�tc�S�t�EJ�*R���Yt+�f�����z�Rn�����X�j[���.n�'�/�hWcfR��'�s�6�w�#��̱"Y�ūL�	��Y(�澏P��1�m��t�;PV�7��PwvL[���f�	5s`��Z��c�^V��P��fn���|6<�Qp�0:�.�o$����ר�N>���s�z��sc��0<v ����{����������|���4y�&Ĳ��]Fej��w'r9J��BVv�t9��^���4Ⱥu����$��nn��6�4��+��7u��	}t�(���W�+���˭��8�]�}(N߱�KY�VM(�Z���\�P� �7z�V���	�L�.g!��c;�##j�#���$�lz�{�)9�H��VoyS�gB�p��EH�[CNmYZs�f�Xs@�C,j]Y��3p��&.[�V�$�$�c�V�/H����އ��Ս��Qʎ�u"l�-��_��'����v��9ׄ���GwTo]`��� +�-���^ŋ���>U}��U/-f�&��3�pC%Z�㖅�t�mf�X��7�p���;5Ztܶ�w��9OX3��;.NQwCZ�9z�_$�0P��+Eq� S��h�3���|3p���5�&Q��/nϠqK܅N�A8��Kj�oJ�<r�ַE�V���ihE���˛9e�Y�]�� Yh�KK�!��te��e]����8Eae�������[�5��y����h�y��7S7�S�N�f���3f��~�d�&Ba�V�AbBz��Gv���<���g	7*�|*�G�rB_!�\�skK��'e�/�aX�;�1,�A��M��g(j�e��{j���.��Кǹ�Gk2�:&�gC��pFWibD �jj�[Wcc��뾽$S�^�72�Ҭk������x�qW!�-P_�w5h�~ۭ�X��@�Y�����(���]� щ�X-v$�%
Z�Ǆu��-j�|�]J|��|NK��Bj�dV{ۣ����-��ԗ�eÔn����:T��Z6,�\��.\��e�H��dT�)�$��AP7���Nz�~h�a���j��������Í���'F��-`Tf���Ė2ɡs[ת�u_;�է�got�{q[�Sm�z����������w�g	���vҔ�YZ$�[Γ���[�M�]$7���9P�f�*{���]��yO3{-ЅH*��૮bp���ǽF-�T��v|r����R��R�,T�����&���1C�V���'}��j+�� Z�Vq�]M�"Ve1Έ쾥���	�;���ὁ]�i�*�c1��l�;�M�4� �v�,<���̲�֗$k\^Rבj��k���48=�D,-�Vl�$�0�{�Ltf�����X�G/�-��K����6P�݋r��T��n�Mn��O����!4 �����
��n�鹹G\�N����\ɧI5�eEZ�j�2��hB>@�%4Ŕ��3Z�(����urr������M��� '�a��&�*�ε���Av�xmҨ-2�5�F#o@�L4�k��]Hb��u�ُ�*ƚWm%9�u���Xo����d���rj�8M�ڻn
���4to;պ������4���d�a۫����CRx��k"�^i�6��$����m/���E�`�]Sd�g%�<^� ��Ñ�q���j#�w�^��ŹOgR��1��!=Nw��x����{����JL$)h��ۣ�<��6���W65�*��yQ�8۪��}��3�w�Tw����H��|�`����vz�86tC2m�ܡ�.B�� �`�m8�Y�P�+���[
�T�K��^n�{pz��%@�J�-°K� ���5U���3J[t��5ohZǭ��+@�D����E\|�{�z�x�lRw6eLq3�pk�7Tǂ����L���ŃrJ��:X�si���H�k���f��e�h������؊�ڀ��}��k�`l�:,�琢j��t�*�VT������j���=�\W�i�7���,��Xj]�hG�z�3�Z䉌��]�[����n����(.����e�`�S��PP�b�����G�����ei�Xf�n��q�ݤ���L�����*vL�\Z�XǤ]�{yq���x������\;����=�7�����ń-ʜ-+wSaZ]�����or�	�"����U��כ;ۤ�[g���;��j,��=x�Nz�w��[�G��06ř�bKak!�|�����Сȭ�!)ǙM
1YJ����#;Nn��m<��=*	�
��f3d
�]`��~.rIv�k��ו����}Pfq��z�0)�]�©��I�HZ�k��]�s�g�|uc�����e�pYw��gz�˥�nF�݄d%(�[���>��L��R>L+�T��#v o�x���������K���5QԎH�ˌÕ��y���(�gM�"�r�a�T�/{5t��2u\��]�ĕFpZ��@�r0�_U^��	����Ґ S�Y&�ڜ]1�&�R��!rD��^�<�`���c�1�M6Umoo���"f��̵�-��q�뻻0�k��
ǩ�����w�0|�\[%ڌ�ȂŮ���Jh\����,u�R��:�Y�z%v���_\M��;1�z`������F�i��fU�{A��tl]���S�>%��%OA��<�B�ۭ����uժj�	�'^�e.��v;��*��i��;�8��lhyY�;�4-ET�g�[�*�;(�ѹ<���I�[�ɵ�ؖ8vh���|���	5ofq��i\E���;�N��������*�Wc����8�t��m�WQ�8Z�e���'.�E�����1{��eUpю��7�_n9�NQ�|1�'{W�}�B�y�cL���P�v�����5�cfn.�w�8�-��k��^غ������H"�p���J�_lI��m���6xо���(jP-e���8��z�Uu��s\�^�H�?���:�{��MUjz�3��̜�x��6" H,TB��/lU�pY	�'S*�/�i������F+�C�U����7���ûHٺ�sm���,rZ��՝�m�z/A��ݖ�7x�06ym���7z�F���3�xg�7C�9�3ܱ\�Y�����b}�%�������zs�$��[ݪ�8�ν�5������D��+w��+��7M|p�%ڈ���g�ɔ�󯝫�BQvH{��<+1YY��܌QK�3A���6t���#��=GkOm�Hf��R��kC��ufhֵ��9��{T�wxx���r���Y�$�J�����.�4����sq�
��۬��n�:�f�r��I�M�Y�����J��Zd�#z��4���7{&EG�u�Yǩ`%o4>��\j������o�K�̅j�Mvԣ)L��#-��eV�yp�2�I���M�Ac�6�P��J��������	���&5[C�Y��)�.�m�Q���Ǯ1�"icG`��ø��ہ��,�4>�`�A�Tԭ�M��ucp��N'ԩeu�V�nDʳ���<i�bM�[�:�ۇqV;|��]YC!.��CS�9��9�:x����pRi�T�W��iS$�EI�S��T�T������_>�atc��GN�[���R���lt��t�i�Z�}˫"3�=�V�\����q��H��� �,顐2��.6��\/����Պ�#N�쾭'4�Rh6=A�ܬt�M����rͤ�h�-����8��������RX��C�ǫ�JMYJ�Ux�Au hƱQ4raա�uL\�{6�R2�WKJߔ cV�<�W�J���u��o!�ќ��J�F��w��`1�Nh�M���v箫�p=U�;r:��L���/<�w�_�uf�2�NDy��:{X��~�#ۜ�=q��(��-R_UWGʹ,���&���ZHfe�V\sg�ڭ]���ȗt������Tz�����Q�4Y�Kdw��!���|G���nU�A��5��}�م�ksQ�;����kt�4��ɺY���� �H�Ҝ��"8أv���k��|Ll��,p2��Y6��`�S�@�YЕǷMu�dv�.�v�,�5}x�qZxUk
�t����j�u.��mq|�~�����E�K���69u����3�3d�!��X���ln1��[Y�b¦v.�B`������ItUq`�N�IHf9Z������m�YVIL��t�.y{�B8n�їJ�B:��}α^��)9����s�O]��tsq���7�Ӻ���0+!�$+h��nնin��qS���}�t�+M6�5>/����x�"
�S��/9=f���Kf��	)>e����ZT
�ۦ;��7�6a���j��F���s#������[��+ʃi�H�<�a���Q���[(8�OR�xv�ݒܪ53&����B��#v$�<�%��ZՇ6θ�ڰ�n
��F�ϥn\���J<�|�.38wi�oԖ�^� 0��l�^"���r�ڈ�M�U���R=x���u��9m&��#���u3���iŕ֢h���n��J��In�R��/F�Fޭ�-T�\F�4�1{3/w%��P�L���$���,-�E�T�B�	���.�%"�y��`{����:i�o|�K��wIv*ن��i�Y���YX+vRF��j s(fÖt��ss*�ه�مY
��]N����+����I�4�^�B�e=[]Gi�;��g[���/-u%�J��v�Δ�d�L�OSb�R����8nB�;u�U�:�R[�ɗ)��T]G�*+�|���h����;������OQ:�QF/�{����g����3:-�Hf����zn{�
'u��P���,����'���{�a�Ҧi31IpVX�3������4v��g��s;�pٕh�Qs�ʰ���R���s�R�
��
�������9B[wE�aG���}�N
�"�L���B��mm���]�-�\ٛ�V��u��
�Xm�|Ky�F�Y{��^��WT��H�s�P��gL�Ӯ�Y]&ղ���{G�DUGQv��x��Y5����)�21�y��lS\�~�@�*.��C�Id��S�i�rxL�gw,mE[�E���<+��zoRw�8�5�k���n��k��S�.R��xm�q�W��#�NW/+��cüz�h�B��7J�N�U�\k�u0��U��6JEL�y�s4�q�5p5V��[C2��wP.��J�1C�6�'�E��"����ſ8�T�5ť�]���bb����fV똷Xl%�o_J[e[��tșhL�]�ӥ ��b"���`���n��Tp.b,�ŭr�2e[�U`W}.���I�Īz�\3nV��ڷ�����M��i�9l��Z��%�L:\�p�ʻs:��Z�L|A����b/ɗ�@�/���FS��J�Ŋ����9���:J�9Eai��nV��Ҭi�r���U7ib�B��)�lTikr��h��#�|m�.����Ã��ZUd3{�GvF��=Ӝ���k���L//�tPt+�\�β��Q���Նnc�I[
*���� ��i���b�W�B6[CI���ǜ9,�� �,�7�[Yu7Va
z�=MS")�@ׄ�����S����݋�\�)=,<s���,�C�}	;j��ؽ�{R_Eyl�
]��������(T�ם��]OtW�9�ۂv�fӝ��~�4��������q�G_kW�H��f>N����y��������E�H��g�9�2��+�T���(l�Q��V�m��r����p���U����e�o0�
"��.��0��VӍe��h�V��'JB���ہk?[�`�B��z�M�ڼJZ��@���ˮ�y�rW	�ލ�+(�t����
P��л�Qϰ���ٚ/5p�	��m���R�X�;�}O��s7=/����ϓc��l?k�ky(��GP�����������[�ћ;;:߭�[�sn����]���j�		�4��RǾ��o�ً;��e�n�� ]���/8�ʊs����Pt�v)0�t��|�"��\O��<��Ȕ�D�~��X�޽P�Z%s3�D7�/A(
P�� ��o�XM21lB+�%q+���g�짭�[l��fm%:6��b�4э��knn���UK\�,~�C�ɽ�^�2i�a��&k�H۞6�����RR7G�'p��|���rM�n���ߧqB�;���L=n�N
�����ti8��Pԭ���(K��%���Ec�N��d�B)�=�����p���W�x�m�F�^�4�x�r冺_l�,C.wٹg�};)�u���}Ra�#��0��"���T�,zyQ��/Խ��=�z�n����OG�A�R�ڛ{j�c�Ei/%�p$�ˊGM���A�r����%$Oj�v��;��P��A�����;
sf,JZ���0�q%6U�3Vt�Vwevl��d��:/��v6`�+��XZ�;�)p��8wF��vh5p�1o3�W>�ˉh;uGɅ�T�������Bܬ�NR��9�n�a��&�2��t�>�ҶӨ#�.0h�`\�����ZH���}�G����/���ٯ	�N
.ƚ��GL|���{"�iC�aV֮Ei�k��¼���v��x�c�����������X�R�-����k*e(�
cR�h��EQ#-rʵ*F5�0D��W-��DUTLe����T�
�m-�Т�[ ����X�Lj�KaU,��ڦZ�YQ��*(��D����X�.�"��J��ʄUU�ET�V���eb��+,��b����J��(�q�ETPc�*��U\j
֨��X���J����.5�"bQnY����R�"Ń�X֕��n5r�"�-aTb0�����(�±L���j���"���W-h� 8R�EƲTFVVTYr�.R�b1e-�Q��J�8�,2ʣ�&5m�ĩ�E��(�E�-�Pe��X�Z�1.Y(�U���
�Q,�(��6�ZT��Qd+XѪ��L�F(�EF(�)V[
�&e�S2�m>n�5$o��J>;��v�5��e��4/$L�����K-}�/o�3�_�ܪ���zd�m�}z��:e]�g�x1/�y��{4#S�ҭ{���D����p�o�u]�vNoMy�*���n��}q��>�_��脥��P��(Kyi!_k+I��oލ߮}�狹�o���|�Pg��<��w��_EV�9!���!��TD3د��N�g��t�x��y])�]���u�]Ι��`J��5B}��Pu��K�ohͶM=��R�����0�a��k�GEh�f�y�=�t��CR�
�î�W> ����kֻ��<��ݓ�sn ��~�mx��Zah�e2}~ql#�v/`���}��,p��e}�|x��I��p`ǋ�*��#]��t�X���]���o�S�jG�<_9�����=�e��dn;���Ms-�.�ђ����u���09n��������Zi�ז\�Lu	g�L���z'3�Ga�&���FJ�UгB�;����]�s��^���u�P`��*�-z����brǎzu��Z��d��t��P�\���+xl� �/ذ��f^t�}Ս���TҲ�t:��;$2�N!QS��u�W����Tz�7��؞f�i�再&��n&x��7u��ÜW��{�"�ͽ�H��b���҃�B��)m�y�	V���˪vp��x�Z:%���8��˚�X{J(�,�x:�웷p�����+R���BbϨ�y�̃DP-	�,���M!Z־�`,�SQ'����(vC�^��0mq�N�1x|a�`�ȔP��j���b�+���߱ݗ4h^�Oox3|����í�m�^ͭ,�y�xq�NY���"D�H��@mu2ǆ�
U�nX��Kyz=����m��l�%�Yީ~-��>�38ߧ���p�:G��c>.��7�A�O�G��T�k�m����M�Ic\Wx{�j�.>2+�j�v�h37Rh�5�mJn]��wuՒ�*�.��.��v���I�����Y~�+��}�~D,}��g�g	�����C��ݗfƑ���V)3��|��]v��'۾�I��w-q�٬�������SfcJMp�%���z7�*�ѳ�
�G[���]�x�;t�ݾj��Jot�f�ya�Ii+య�,0nJƵ/}Ҏ��p�Ko�ݭ��CX�� ��������V���� �c��tZ�ѻ���R��^w'�++��(z������%�v�*齴�>�^��'*ڜQ�_&k����z՜=-~�/j�:��ye9�WL���|(����w�ݖ۫o�~5;j˄��ʽ�����=�Wc�i�������$Xg��|7C�����x �3�Dh�S��6��'���!���_ǎڑxo�����zf⳥�v�v��iԣ��U5��l��<��y�N>�=^И�Io��,j���v���b� ܶfS��Hq?,���<�j�Ҙ�5�Ś��K����
ý	��c>'�	ʞ�J��*���8eQ�S���a�1d�j���8�*��뚽�C��G���ݴ�4��[U\f�M�P��=��kZ:d��n�v�|�Q��L��oWh�,kXm��T�R,��-��o�q�oX��;�[Vq���ܑ���M�e�=;����1S�	��XTF�y�M����W�y�I�������d��Z�9S˾S���Y4z��?N�%�e�"0-W��W�[�tý��eR��O��`$�]�:X��L�sW��p�ߥX�$癆d��5��Gԭ<~Λ��7�Վ��`@*�D@�/�
+ƃ��;�x;�5��W�*]�c�مF�?)�a����D�{1��)|kb��:�i۰�*H�+jy���\�m: ~�e}��=��,q��:�ٮn{ԟh�s���7���(8v��$�\���R�c8�>9�F=�)��V��<��{L��j�����c���b�^�����*�i�4�*�K�wr���"��i�\�}��ٻ��4_��;ǃ�"�q�6�`r��¡����Ћ�e.���e���T�^íg.��^�9e�8;���/�`�r���a��y�z�L�<�CF��S�O q��b<����aċ��lL�-�Y+@LƉ�!�I�#�}a�z�W��z�꽹�~M�p'�������C=�-�����C�_�����ȼ^�=�N/sk��l���{f�Y��[\~�� u�5�´�Mu��QF���uZ�;���.>.��[K���W�@��=�)�<o��oޥ�%�^R\0����u;d�ȴW�B:;Ӂ٦4�٣{y�uP�PW�0o�2ҹ�~�*v�uF�XUf�]��b倹�ق~����^.B����	��8D[,��n���9x'���xDOW�ocy�b:�wtOE��,����������ٿ���L.?z���2�ӱ�x��jeH=n\T=t�<�kЗ.X�S:'n7���V�����ݳUaջ�]��d��&��(�x�mD��1{r`�U�fp}�����	{;��O{�W�����=�vn��">�'�V�(ߥ_W4]LC#NJ�=Q�:@-N�����~��l��3 ��f��<���C˫��Lc��3��G�\'�<_�K�;V�q��<W���Й=!X��,�G����z�����9P�y��Lۊ4uw�{4�op�i��d���?mܙ&]N�˯���>�:_��r�F����ד���x�]� �~�rgz佬�.İ��k<h>dؤwj�d�6[��C��������}��<��pI/�K���	A�.b�a|Lw�}ޱ=�ڿPE`m}E�9��p��$��ELX��$����$$(�,�ܑA��ywݗl�L4&��=1�}7{�wBq�P	-��f�׹z?kG�Z���ol�� ���;=���~��_S�|jOK�]��t���%�:���t���f�_���q������S����/>Qz�����/�)mG+Q��X��zd嫱LU�v�ˤ�jf�v)ɪs��,�+��t�9u����U�[٩r��0�X}sKh?V=��T��l�ȭ�vq:Z�|f�	�A8
]�g�ُ=D�Q�b����筫�_�H�k�7��߼�;�$�~Z��
ݡ���<��ӥ��Z������{�Q�Z����W���ӌ�9��ouެ���8���ఔv��_<��:��,f�W�}���rӗ��.N5��� �*��N�K�F�>�Q鮵��O�\�A��ٿ7��;����.͙�����c���5����³��C��[.�������{ ��<���&���vv^���΋z���1�{��漴op��;�25��u�;c�۞̑�Bgk���`�_���Ύ����<�9-�*��\�K��;ڲ�'����xl�7����t�*U��}^�4iW�9*������{�Y����s�����z�q�x\�՟L��4M����*����f=��Wq�����=��.��#��U����%h=R�F���I�Z-�CtC��[M+������q^@O'�'�m��D�z��d*D1F��<�e�{u��_dZ|E�*�+�ѽY�.�a�VZ#/�"�Moo����T'�4�rL�Vc	0w��8?��*��\X��3����jҸ�>.��W=�����z��Cx�.uz����1����`9����U�9��q���^����ۙR���{,'������ʱ�����*�s/=�|�ݓ>�ܮ;b�Dg<�qމ��`����y�z)�U���בz��$�o���B8��&=9�z�u/����#�%��<���N�t��ڝ{B������e�p�8ؓ��y����� �Z���s�{o;�9n/�;��r�jO^��K�^����O{�@|�u��xo��w���@w�ZJ�a���x��|� ͷ����}�K}tt�ջ��;�Y�G�7����������p�D��n0s����fk�V�{�����:v�˓������|��gV�rױ�d�ź��`=:x�m
��a���QΘ���u���Y��'�S��xoQ�ۃ��*㍒��-��u�w�	�#H{�o_�}�!�5��C^S��@]��wH*+C��%��#vfv�fQrT/���'�ۛ5��p���}�ɩ�]��k!n�d꽼*ק8�UjL�I�H�}��{{v�Cd�܌v�=1�|�ک^�aN��Ğ�4�&�ǽ����bz���Pp 0��2𥮭�3k����]�3nd�z���_�g<�t&<NϲZ���'v�3�J!f�(�t_W��>͸�j��}��y�їXt��Y��S��,��w/k�U�Q�
����������<4ױ�cb����0jw�./��;^�9}x.K�a�wv+e�43�3uu���r�{}����\y ��9|��>�q�T�>pV�M��S�P�{/��W�����f�Q�gy�{�і����Hû݄����L8���y�Kn�^V{�{6K\�^���Wys���;�5���$/M��MW'z|p��}'�����;G�o�3�O�^zc��ۘN65�_�"v��ý[C8^oF&g$���^w�/z�>9�J�r�foQ��4��;�Q����#�~�0��v �E-WS%ۭq��v���=�>�~4��Ii��XF�����^w�~iH&M�2N')�Ƕ��-�e`�|�L��-a�iһ��7�kb��`\���Ѿ}pD�*g�;�Ѕ��>[����(��骡DOI^Ր�%�쾮Jn���y��v�=aS�*{��)m�i�.�בI��n���V�����f��sw�[���-U�\�ߛ�����L>K:���<��vL�dA�v��d�m�a9sN��{�ؽ~�������*��MM�M�w�Cpgգ������':`.?g�;�y��<��Ƭɒ�i���˼Z�TB��c�I����6`-���}#��o_�=��z�m�<����O?R��6o�݂�t=�I�&����W��vN��mJ��k�F�w�8|����F\U��Ϧ}� �P�=$5۹� �:��痟L�/λ�h���ϭ��eQ�;듙���|�Մ�N�ƞv|��c\��%z���ϻn�ϮZ��2��x�S�<�S�[�ކ^J�ӳ�WE]�$��%�_�`�Y���KZO�0�a^���+W[u��㡎cÁcW�0h�S�7
��M=���m6�
ܺ�÷��uJ��$L^m��8��<�rUɶ�V�(�π����xT�C�W2�n_)v�����m�]����Z������!j㤭���̉�*0�m�|xړs�IH`�c�^����.��%��EL\��s�O]����jvJ����&xp��ԣ���rk��o�ʝ�y磎!w����fW���uZ���W���=|�����.f��T�w�}�z�{������bĞzpt�_���q�ݞ���-��"U�Z��������̂f�>|���Kk�����;=�޿4P|AZOKWu���D���ȧ'�E��^��������8��9��{��fi�ϧ�{�y9�+U��p���]��5����L^v�s�-9~����;�p���Ͳ-��վh�<�"�u��'�8�+D��f�ܰ��tKn�����K��5,�o��)㘰�:ϓ'g
c��:���~�	��[ֽUrߧ�cl,�s����b[�
���b�c'_��]>���Z�W��״�{)M��Tw��u+�k�*���h3��'��CQ�^S����Eٺ��( �j0g��)��-�w��	ދȔ
�'��(w9��w� ��ܚ������}M���w}�����p��6����)�%tͪ$G��F�p�1�+���i*y��9nAR"y����K{.��Vl�e���0��G�/�y⩾����	P�Ɛ��h�U8�d�h�!=|Rǫ�չǯ.��j���m���%��i�|�˦t�Ʊ%�ٯR�Qun��x.����ީ�UИ��DL��o��T�t�ٽ-����NA]/.�tB�v���`�4��q�m~�K<O٢��W��F٥���ʑĀ���x�/V!ĩ�JT��R�^���6�+˘D9f���ئ�El�`�l�Kc2v�E���yW�ʑ~ik�8O�7��w]�r��j[�@U�������jy�O���˛�%_�v�9\g�+�Mh�K���hC�-X��-+NR�-���N��oQ���;�5���R��S6���s��e�����<��-+�]3-�e�/�3_^�(��+4�Q1�"F�6������lǌ�L�x��q�u�ڱ����副�.숹�V W%�/��.��V��]s3�p��V'%��x���a�˨�tk]O���ʎ�{WvW�!c�f0Mu����J�F�z��z��*�j�q����PM��>ݘ{�EL}�+�qͩ\�!텟Me>���L��^�������ׄ��J�ĵRrhNl���{7�C�tbR���"�Ӷ��^Ἣg�N.?4�h;WmOq�p�=���՞��u�ru(�\�OR8{S�)pZ�a �V�ʊ�Q�%�)��KI�:�e�,�ՠ�\�WX!��ۄ'��H��rU�r�Ig��ǚ

���D�VͻդE9�m���9c�ITHI��Nk7\IpU��Ts�3ۻ�t�A��r������H�W��Ua��q<�f�}/M	,sB�I�j"��pL��$�k���Zu��]���	�Ĳ�\9����u�B��o�H�%($���6 o5gou��;c��K�Oj����zxG<�8Q �u��,�P�hfj):��ئkv�Oa$s}��)^ 8s/'g��̨��.�2c7.)iWV����+'ZL��ȴ�f�X�M�0��"�k��U�󳹗�K��M\�i��r�^�jǔy��*�'=\Õ��'<u��u�{}�h���g�:��}Ơe�|su:Η��SD��fr�vSN�^V�y(曻]0g+����8Mp2Kh�j�|�ˢ��x�$��l���TЏ�gi� ^����Gr�c��9�k�G�]�-*��� �nӚ�\ρ �-���W��
�5iBUE�R"((��RF��Ŭ�EL(5�q��q�r�Z"�QaKK��d��c��*�-s+��-�mC0��Kh�se���F
E��Җ�*
��ER��Ah,F
���V�j"ZU�ဉbU�P(��Z�R�`�7,̳�m���Qq�s ��fe�D1��K�,sq�2���`�Z��U�mm,JU$�SKV4�B�Q�s)��)r�b#���1bkA��VƖ�X�*,��\�.Zf.8[\J$��2ʪ�Z�������QQS-EL�**ZY����fU�1p��\���j+[%��2ɖ�WnV�Pr�L�X�2��EL�I��ƥIF.70�GR,QA��aRa��[1�V�k*�EĬf[ZcE�e.f
�r�%eB��fJ��h�
ʕKJ�TTR��fQm�P̳j�ڣmA�������-<��B��E[C��"en��lW=+y�`�lǱ���Sa(�V�z,�~�C\���oL�E��$vg��������3f�kgk��I�3`}r��tv������kL�g�{���V_�)6����{�f�޻w6��#�FDFz�;P����qs�s�ڮ���E�|^>ܸ�r����W���y���d���&Uʼ��7�A,�1�i9փ��^�mt�׀J�v��~.��<rd���{{�J���Xu�P�x�s���[}1K~�r��H�g.r�Փ�*S�9S�t5�ܛL���{,'��S�+��kV}�KՔK���m��������Ň��t�ÎƉ������|.�l:���6�r}�;'���3����1%��޺�;5�0[R�{od�=ϖN�Q�>���M��ޢ��[��9�Ę���7P˜qi7S^������o���uj���6S �߇���;�6��θ6�lr��{��s�g�=;����]��㙝42%B���,�Y�+c�Q������e>�H��&����P�LWn��i�,�v\6��CA�x{%�kXHy/>1a5�g�����E�B�8�U՛`H���ẫZ@5�O����R�9��8������6�ki+�m���*�	�gl�۞���z�I��~�W=�ʡ�,�y2}�ci��'3=���y_a�/O��#�s�����c}-9s�����sf�Xr��4��v�^7^�P�S��2��'�y��1(G:a}[ԟ���{�j��j�{����;�'S�Q'�)�����?`z[ɵ�=���'J;a�3���9���5\�dl����Ϝj�|j�貮d�P��J�;-^T+�_�nKޛޯt���\�j"Ʋ�r�C�_S������xSo#dh�A��*s\��u�f̼��]��:vB�x�As�9|_��v9���7�]��l��ߣ���R�>r_^��K�7����b���.���V}[9�f:^G$g��{�EQ���ゴXrm���˽}p�_k�+ ��ۡ��t}���%�4�v�.���/>�g����K5{�d��ʕ~��dc���r��N�{g�j�)}���/B|�+N�u��V�k���4o�v�̓��JM;�g�GME��X�����V)���L��n/��c圢�|���>��o��r�����݄�r<LX��^�~�3�(<��vF��c��=�����D�B�d�:�����'���]���X��/W���EB=�ùuO��=�������Gõ*����x�՞��VΫ���6%����2��_�N�n��	�����9kݹ5�8��Wd���؎�N&ξ�Z�=��1�*so��I^��5��׺t>U~Br�B��zej�}<�W^[�M����rO�ws����}Aw���s��f�ٵ��S,��c�/|ٟm�s�o����:j�ݽ�����������Y�ֺ��<�v�N�.���Z7�pl�7,�L.?g��i���׵���i���lc~��P>;��ꖖ˨:��7���ނp�6����k��u��3���o�?�w:;�Gh||X�w�;+�wY��&4m�@Et�����҈�
���e�u���	����?�6c��ͪ u�I���M�h���s|��[m��k�4ۦ5Xbi����fM�a��)�{F�Ѿ�Ŝ�!)���.�M����4����d߃�=��V9�tOr���;��lvW��E����=�y3{0HXδF�cN�hs�����,�<xj�nJ��Ӫ���_s���ގz{��~���_rk4x#��tT�'v�)R�pN�^���V�ގnA��:�X�&w��{Y��w,:vC'9�e��0m�G(Om]�9�)�~ڣ-����WE]�J�*a>��{4V�^솞�H���d�rqvʱOsocᬻ���\�ELWg{��ݗz=��.������u/���D#���g����Rq�l���O�d�!�ϰ<v��N0��� ��d��βJ�����<�Y�r�������z~پ�1'�&'M�2q��l*d�+�w)=d��c$�>�$������N�`T8�?>'�Xi����0<z�ĜI��=}�^��<��;������}��z���3�'�*�0�$��i�N �6w���M�����
OY?{�I:�����$��	��'R��I��s4�_g���~��k��;��>��Ь?0���3L�0�Ow�@�i��/��a&��7�:��z���:�ĨMN��ԜI�T9��OY7�3i'P5�\d�'㹽��~O�{׺��|���a8���;�0�M�G�4��'�_a�i��P<�Y&��'P_7�$���Y���=f��d�T&�}� u���~��'���y���߿y�x��d�L���=�ɷJ]n��W��!�Cr�M-|��G�f䣅.�$�}�<��{��g���6�/���w�'V�N?�J����)#Ś7��X���:��^�h� �׼��M��ռ'Ms��I���$��1���Cl��I����Ԭ�j�Ru	�_b��N �jy�I�8�Ԭ�7�	ĝCFs'SL��y߰�'���ݾ^����׭�u�]t�&�9�'uܓ�I��IY4���'�I�'��=O̝J�0�0�� �M��`u��,���a�I�Tײ�����"��]*�k��r������~�m�op�'_XO=�0��2xO����I:�g�%a�!��6�ɶCYd=O̜Me1�m��P�	�~��d�V{�������x^�߾o���"�i?2�C����?s�$�a���<d�'�}2I��&�u�q��/�%I�������b��-��:�ĩY'!��~'�eB�u��涮|���ߨz��V����9���H,�a�����&�y���$�},'�N������?d�&��g�VN ���<�����39�������`x�?'fI�M��jé��u�}��N>�^`x��N�C�}�I9���&�4ɳ�`~I�M>w�I��&���a:þ��4�F�js���<��UW���	��N�Y<A`�m'|�L)'�:��a��N3��`|��l�����hx}�'Y=a5�g^2x�����:�2|���È{�k�!��z��=ܗ��o��W�bq���d�C�ް�	�w�+'�~2��N$��0��d�~��!֤�f��d8��:ü�Y'����4~�O��so�g�_��,�f��;���G３����i��,�P�C�M��d�C�5�T�&�VO��~�I��}�����O��rjN�qx��"����-�:mخX����6���Y���0�y��>d�yۇ�N$����c'�,�s�!�6ɣ�a��u&�y�T�&n�d���q�l��Ld8���w�ʬ��{��Ocn����m4F��nȃ��c`�QSJ"��(J����8"s�2����+B�d��[m�7�C!���}�0���ύ�7 �8�C�C�ۇ4��Bt�Ow�tH�,���i�/�ӽt4��վ^x{6/g���<-�]n�*m�}�=�7��'��M2z�9d+�O�?��u�T�?N���	����'R킇̞�����=I��~I8��Y.�����Y:���w��5����[������ܓ�o���m��2x���$����i��y���IR��=�Ad��,�N �6w�<I�M�a�i>�wە���ߏ�J��%rV~��7i~轾�]��~dXi�Ԭ6�4����d�!�^a�u�Ĝa�ߙl�'��$����0�$���u�䬆��q�iX\�����=���^n�=��}��=7�����N����d��̒�$�'��}I���C�&���<��0�����i��:��~d�!�N��7�Ğ���0�i�m��{׾�g�}}�s=��<J�w����Y6�'����O�5>��=`h��ֲ~d�ja6�&�Y�I�T�Va��k�!�'P5��&��'P~;�yϹ����n����?{�~{�o�	�O�_i�~I<C�~Ì�݄����'Y8�'��@�	룾d�����O��������N�g'�Sz��
I��=���ܿ�o]9���߿{�ƾ���4��ӽ�)6�Ԭ��p'u�:�0�a���|��y9��Xm�'���u�z�Y+&�CԬ����C�~d�]~��\?k���7��כ癟w�I�?3�$��b��>J����"Ì�J�y� �u��N�d�a�ì�}I�'�}2I��N~�q��6f�J�l���̖��3�s<�]�[�|��i?3�H|��OSFSN��h?P�~d�:��C��J�׼�,:���<��HVN���d��'�Mw�ߙ<d���u�M�|��-����|��_p��m:w�IXx�~-6¤��ആ��'R�a>I�����$�џd:��l��d�'_�}�	�����}��]��G��0+d8Vf8�eXw�b��P�c�gP����O�o��wa���j����%U}@�2z_g�J��	ڥH�����]�9u��y�5�?�Zr垺��W����&
�CNm��ĺt50`Nܦ��v,�K�7����;�>2q��|��g�O�XVI�~�*
��'R~d�':��Y'�8��C�~a8�O�`|��ԇ����K?	��_�,���~�/�d�$��so̞2i'ud�u�I4���?2p�,��~9����0ݟ!Y:����q��	����>�I�o����������g=�gw�zd��O���>d��C���L���>w0�&�m�w$�i��v���7�`)'�sY%J�a�ĕ�䬟�(0���l�y�!����Z�?^���~���9܇��|�^wWl�CG���$��<����u�s��?2q�����M��G;�:��5�0�?����gGT���-V�K��c�;��>G�/��)6��&�Ɍ'�5�>�q��{�p��L5�������Y�d���̜AHh�r$�5��
���\��C����ٟ��E�V~~��#���%ea>���d��锜@�Y�u����y���'��C���>N�x��ﳩ%eC���:ŒT�w�u��	���*��C�[�޻���@���J�Nw$+Y?��N }�%Ւs��'��:���8�<}O���C�y���'�8����6�d�9�u��
@M�牺���v_�������Q ���:��u*\�ORq�iXy>�Xz��{���u�_y�_,'�O�����2O�����a?k�=M2u��O�������
�}�wEw��}È��ϩ'�q�Ns����S��Ԝed4wܞ��&�d�hd�&�}d�d��'�d�'SYB|�ɤіq�zʞ����v~�}��o��Ǜ�z���#�������&�>Ad�{�hu'P_�q'Xk9�SL��xw'Rq���}Ì�d۴���6�o��$���?{I�#���
8�~�����wtw�m�w<�g��s����:��{=�pV��2!y����S�c;^6��øe��en�n�k��t�Yo/�^G���}7;�	CU���N˟�nao��8j�Z����4n����ŧޫ#O�r��%��"��ַ{������w���{!����&P�$�*~Շ�L?l����,��}�m2u*y�d'u��s��N�~���ya>9�8��N;I����d�s�|k�f;o�>�{�<�Ǟt��������|���z��6�e�a>B��u$�~ف�N�Hh�삓��J��	�a�9�_�'X<�Y9������y������������36���������z�����2N�����C�l=J���5��?$�4e�I�:�?Xu�����I�V��AI�N�C��rAd����ǿ��?�w�[�{�9��O�1�$��K�笟$�=�)'_�;�²M��~�+�?[R�q��Hm��5�O�q5�é��|߬8���s��ߦ��׳��}�(����y��}�z��'����A@��N2i�þ`~d�'��,'�MwXJ�m��%b�h�>B�q��Hm2u5��|Ì��þy���/~�j�]����g��>��߮���j���(=d�'Ϩs�u�l'���xɦO;���'�4��B|�d�5��'�Y*
[��VN�d���Y�;������f���=�~�����=���O��$��5C�d�O��!�'7d<�a�I��'?a�OXMo�u�O|�u4ɶ���rC�4�S��Y'|~����oz���浯{�y���T'g/T�2��ei8���c	�M��~�u����>�
퓨o�q$����4ì��Nܟ�>a�;ܓ��O�Ynt�u���v�mW��]ד� ��G߄� O��G���R��x�����s)8ɶN���'6��7��l�d�a�a
�Hov|�T��{��:�q�������{�\�k��ϻ�ޘ���C��T:ɴk�`N��MwX~d�a��d�+	���E��,
���d���~��'�}�㴞2q���m�d�~���y���o�JZ��N6�E
�~�ѵ�f;��r�w���"��gr��m �p���N�.��YT+�p#�R�����[�>���jk%뽣q��ce2$
�p�N���x������=Bhv�}��dXގ��� �,k�;Fz5�׌�<n~����H�r�g�_�|.���o�>I�	���a�N �5��*d�V��AI�'?S'x}�I_'4o$Y;���d�|MO�4��C���l��^���������u�{܁�i��y>�:�|¡��a�IS�Ӭ�A`l;�Rq&�P���AI�'�u��'Y5��%|d���Bx���0S�yB�W�~
��c�5s��|,���g�P�0��y���'�8�z�=O̜A~��I�:��|è,'�st�'�>;�ORq&�P��d�&���O��uU}�ϰ�����&�i����=�7>d�+	��O��,6�z�3G�4��O����4��(�$�d�������;�:��'���0�'�;���ݨ}��:���O۵�ߡ��S�y�^@�N2sWԘ������'�O�P�!�q�I�,�$�+?�ԝB~�ء���,���hq��Y���8��h�̝M2OY�u�x~�?{�o1�f����ܾ��OXN���:���~퓬����+&���>jO�8�e	�~d�h�8�|§�T8��?l��N��k�E'q�;_��i�k7�s|�ם���t'�?0�o�d�a��d��	�����O?w��q$���2J��ACl��a�=�!�~d�k)��hu1	�|ȧ4���߿w�.��aw_���IX;�"�i:ʚ<�H,�a��ï�'Xyy��>x��OC}2I��&��$�	�jf�J�iš�+'��	|?��1�w}/�����βV~���3Y�N2O�~N������u�w�N�`j{�:����l����|�'4���>x�L��鐜g̚����u�{s������[;���_�fw�I�;�^�~B�z�ö��=J2O�|������>u���}d<��2q����}�I?s���'��d��_�x�O{I8��;�=��Y����.��y��|�s�g�H�����{{�Ӵ=���o�������a/���4����}N-g �і��l���fsѕ�kWnk͡�J��&�f�J�٥.f�4�Bv�ٷ�]7��T^c��,���2R~�$�`/�^.�y����G��I�T��+	��w���3�6�d�ց�N$��|���j��d�g�P�������XO��߲u��G9�x�򿫯�o�I��l�B���3���W�3�N0��]�N��5>��8��sXJ���w�+'R�~�@�'|�XN2m?ȯZ�q��0��N��ì�o󆹭�[��.~�<������1�l':v��&�m��p�f�>b����C�N���N!��J����8²|����N u�����a8ɴ��rjN�q�}����m��O3]���5�=�|I��p�	Y���0�$�Zc'x���r̛Af�w$:��;�c$�ONy�T�&�0��:@�,�d��߭�cٴP?��ƿ=������_Y�&�6�M�$+Ԛa��:�*V��:ì&&��ɤ�AHs�
d���0�I�OӚ��$�M�d��$��͒�O���\[����]�|O�q���_}�	����̜d?�'���0�OM��>f�:��ﳬ��a����J���N��
C]�Oq�iXxw)����.=��1�͛݇<�߿o_A^����'{�I_O��,<}d�h��OSG�d�!�^a�u�Ĝa���f�8���0�hu�����J�r�ḡ~�fV���1r.��@�	��������q+��6ɣ~o������]$�'R��|I��0�����0�	���m4�ԝI�Y>C�'P}�C�@�~D�T�X�=m��
"��}�;;�8�Ԭ����:ɷi=�2̟2h�������OZɌ�M��Ԛeg'�S�Va���2�q����j'�v*��J���K�gﾄ?O{9�П$��a�i$�;�:���O;�8��N;I6�z�VJɤ<�����qL���'R���Ԩ�g団�S��˙#]���^c��WD��L�A9n���,,o�}�sv�{���������W���Z)�Y�Hk�U�(��:�WV1B�|�ZF�Y��%�,p�"jr�3Vn�N��f�P�(����6���=����ZI�^�a.��=��GD�+Ԣu����������~`�zD�{�1P�뙐�*�
�'nh�� }���&e�zy	�Q��BBW��^D��,.��u������� �̺�Z L&�ܣ�Պ����s��,��&;�
�4�[*gg�^�w�Ѽ�'�zV�T�bdm����{��5���ؖ���%Qj�U/��"j{����{��{ ^�6����z��+%�Ye>�dm�@�P�};�,���L3{��:�/Q��B�e�8N���W5}���5*E>����U�ap꺘.�m:�����J�0� |���xZ�B9��	I�j.�̮ l��Oy�(��O�6d�s�;E��1�ro�V�r�*J���S-H��2=מȓ��ط8�8nM�5ۅ��WR���Q�!��ggu/���ÛA�l���bR�]ګ+R�9WY`���40_���`N�k-]�ֶ⨴�Mu|�Eh#��!3��5���:-�x$T��`%�beIJ V��4֫�S����I��S��bA�9!}\���q��+����Loy���
a��ר�r���^��y�i��.�X���R�Z"�;���ky�+����J�dz�E��&�}�91��{=:��i�"Ү��8��ќK�
s��f���n��9� �����D��0Dm�as4����\�g���}b��{�+����_J"��n=�ǤYw�E�]�i>z�}׵EK93��-NGM�(�M��9�A�?���1�|g֮4��[��e�m���4e|�������?L%uA�*���\�4e��'�X�΅����u�w`��J=*���yR��vG����cn�ϻY[�(g��V�ʁ�I^���Q|��[�W�zUzr�2璘D���՛�������D����5����n:8@�p��1��=|=w^��������y���|�A�3�3�'�a��������hD�%\v����",�����ķb������gU"p�Pp��k�r��ᧃ�	��.���8㻰�0��}�Pf�\'�FTWS;��TFЬJ�u�hϋ;���n�=�<['�ۗ�� �y��bR����a�Jl�,j{_�.b�76S��o��m�C2# qM*fVs�wczg{7�]Co&&�
��dգ"��6�k��-S�C�7�� .�˗�Q$pR��ޡg/��<)=P'��Uh턨3�,�N<��qɔwD/v�tS5|`�W�M����s�;��ʰ�c�(���Z�n�v����t9�	���-m�v�oot�Q�x3��~o�s_��_nZ
��DPTLb�h��B��AQQDZ�FEAR���3G���*�\KX�erت6�L-ƸԅEK-��ZȊ�ҋjU(��*1���1b��UTU+QJ�.8յ��`��c�QX���b�&9�%TEƙE�nR�"�1��V�mDq1��J���C)El-�PF�UU�֬�Z�UT-�Sq#s�R�Uť��[F1�j�h�Kj�����E�\��`�m�ZW2X�-��Qf
���1+VUj�s)KQ�c�rʬ��ŵ�������)m�Y�2���D%��
(ێ8�Je̖Ҫ�1�b������ڵQ[j��Y�����s�"4iT*���QVe����kY��eXP���--�UE�4�q\a\R�c-�J�\�Ģ�Ŷ��TLj8؂�b��Q��A�UQӞk5��:/\܃��ЍF�5��J)�7)��שg������N�(p�vkx�O���E`�=����$���\��9�fk�s��_��*
I�O��$�
�;�Ru��Y�y�8��k9�Y����O�O���Xm�'�]��:�6��d����m+'�f���:�o8g��}���ܐ�>d�����x�����?o>d�V�R,8�Ĭ�y� �u�y��Y'Xyy�Y8���Og~��id}�e}�?�����}��w�����_=䕆���d�'�є��~d�4e1$�f��:��'Ό�!�N%`h��E�Y:���w���~;�N��~d�(~d�&ϟf��7���[޻�;$��N�XJ�6���d����i�'X~����'SS)�'�8��>g��F}��'=��2q�������9	���b}���G9[����w,�:#x���#����c����3��s�ޭ7龙!�����Nyy2L�:����\��9����ǰ7�t�U��d�W��'n�	S�%_�^�%��%��;���lzG����MAK�5t�Y��z�����F[ݎ9�J��O�����b��"^���s�q&K��w��3sµ�����ۭ���G�S$/E�>]f��0O�W������+�v�-���C�C�괔y9<r��Ju^������gxn�z�����k1���4�g|���Ժ�l1�F����R�-	��ᮏz���&��)k�C�Ϥrc��i��]c���ߴ̷�"��s+�8k�3�g���j� _^��k�M,3<�*�Ž��<�b�{o���x����|�g/�\sb���y����u�z2�S�_�n���ʙ{�E�I��[�/3S(�57��:g;A��ٓ����=~�;;���S;��N�]t�ҷ�_�2�I�!���~�7;zu)�-��M�S��S��y�~���4QZ�z�w��;�EɖgۻB��={ �6ܿ������7|-��Ø�-ՙLkFc����rׯp�jϝ�1y��ͷ/�����{>8���*��վ�gK~�*%#"�^[e�w_[��ῳ�f�':Lإ.˟r�l�p�]%f��G�MZ���3=T˨:��6<Ğ��<�M�kr�Z�u�y�6k�0���'_�����>/��sQw��]�҇Q�܊��]n�í�0I�7�X�&o;Ϧof }(�th9}YV��/ͦ��W^�a�Dr��@^>��N��yy��2��v�AѮ�|12߅y�ĐC�M6u��ۗ)fh
:�(u��xL%h#�c���<��>tf�ѣX8�d�g�j�;��DD�澖xŪ��8�Wn�$�����IKhv��D�e14���xM��Z����k�W]}X��+����z�s������|��3-]��;�K����L�����ɝ�Kک(�;�Z��^#��ݾ�̃xd�@gh':����B�g��aվƫ�v��@�KZ�����u*y���;W����(��2$��E
�p������*b�B�I=��XxL��vR{꺌�{��s'B���;�==�6��3��\=�#>�t�㱢e|�����u��{�Ěq{o;{r�~��m�긺V�w)��>�����ɰ`|0_v�������'�ǖ����+{�2�����~}�[��{������z�D'Ի�vx��z��{��X�y{N��Ԏ�u�{�;۟)��m�ya��㼷֜xef����}��~�vQxjG|)������Q쩆�f�����Uʺt�\�;�֬��L�B���H+z�ц��p0�wwe>��ɥ�Ƿw�m�m���j'�&��Gq�1����0\�����
O���y���N[����U�q0y�V�:��aU��M�W}I-�Yj��	��SGc2�I˓1���]��׬�m��+=�k&�D\;�w��?D\��J^��?��iΙs��\��=��e�{{-	w�M��&�I��6��^ko�VB�wM���G:p.s{oK}j���b��=~���//���tN�R�6ly�8����x$�6�,�'�Y�̳@�]��c){N�}ψ����������ͯ�oe��w�Gy�:���C������_��_�����u��p��S܉~�c�u05���l+Lӧ������Y��>���܅���N;�ǧm9��Y�۽�k�������%��Rz��3�c��МϪ�ܧ�#WmۭE9��K��O�=v�e�2<�EO�$5�w-�=�b�[ǒnU�P%z/f+s���uT�!n�������&��EIlzuM�t�jx�s(F���	���^}fK�;�2˫��y~��{�gt&��1�6�����sqӧ~�MX�_^{_r�ڞW3�f3�+4���j�q�1����X�r|m������s�]Q-hK����M��c�c6%�];|��8��F��+S3�ر5tR���U1��*�룇��٠��X���n�ɮ����}�Y27�/�6�#f���`'����^zc���c5쿵�N]����dwj�I�㺭Xcy4��zק��|h�C��㽛�ə��U���r'���������pv�lOzn�WF߷�Y��W�+?{����M��[��,�!�*ē��r�r��ǳ\���^�*�3k�Q���飢7|��j�fMT��	��`'.`=;�NL�e�x���7��R�I�^�����Z7�����#�0���i=I�����{{.o��ǝ������~�9/�Wr�����5ܲ�ƴ4N_eh���u�gk�GG0��kV�;�C�z�G۝)%���z�����[�;�gZ#x����9��>�_���_v߽=QW^��{��<�8>�6�痟L�/.u۰�;!}�a<����a���b�b��^eb��S��ɗq;��	��f����QHЋ��M�+;/w�e���X��+�5d����]`U٥S͜'RYݜe��3����V=���?^�:=��[݆�ⴁ|�Z��g��8v��70|������{��V_k�����ߟ.�~����x������y��~�ey�[r��z�7y��U���QJMt_f�����q���ݼ�J���� ���uI��q-��Jq��&���b������{~�������*a����U���?�pNwOl������K�%��!�z����%NO=v��X�捹]�z��9���zlϨ;�c���b�{)���mb�,y�Y��H��4�7'���7���m���]�Yg�����O^�)g�I}6��u��#���o��=�7v�3�bu��tV9���_�g��<�.3�:�z?==[K��Zg?�{Q��u�y���*p�7c��OX�w�������Oƅ��h�^v�s��4����2�sY}���ļ;�Is،Z�e�n��PG�����Gjq�3�f�+���=��<�U�9�����=e�=�p�=ޱ��	��3 �e��W�b=��r����H�
m�sP��'�k�����H����2��o.����T ��`��g ��C�8�>���Y��P�k9��AU��:8�3���~��[�-�`�;���������c{\����Ξ��3z��Vv��w�]N�Ke�|��4�L�7G�A��=������l�����K;Pޟ�\�{��8Z	�1��C��q�՞��{������T��x&ofHX�v���c�!��=��{4ʪn�P�C�)i�q��ͪ���?rs=���}7k��l�7-�P*�#�o�0cv'C���|�K��y�3����ɝ��?XL���fз����d�}���^Cl�7��U�{[�]��ƷJ���-=�M�M��WÏ��s��b��ΰs�&��Y�^��=����5�z�<�����;&n���vr�݂*b�/E�$ۗR�(p젞�������q�R,�K��}�ϭ|��9��]�S��4H^��3���a�`h��7�O�{�4F�~��ڳ��yZO�*ro������Ę�w����Y����b�'���frpsY��NZ�k��l!w�ޑ�.�n�mf��yl�
bpZ�L�,��'���Y�ԃ���~���3���P��6�����+o{-��E�X%\�:�d��{��7<R1�V�0���=C;���*�|#�a��&��ɿ�}��Wŝ��������)�a�U�^���J�s��IN��dۼ�Z鍕�D��Y{�����8�]���׀,��~�����3�^�0m�X�^���:>�*3{Y$�R�V�{�ov�y���v˿��=|)����{�Fgٞ��g�mo^Tz��s{�k�|.OZ�t;�;^�i�ll�;ь�I���U/8��
��a�s���;ӽ��L�~�[j0��
Ya{�}cdw�0�p`r�3c�Ho�P�ts�6u�o��g{n�#�Ѝ�S�2y��|{=%�N��6o�<�|'Bgk�s��noH�mq�Lތ���1��Q��,U����U�&��F��������\:��`���U���Z�����%۳*Qo�>#�ilvt�/ٷeMYD�0s��<����?m�7[R�[�����a�ݢ�1�u/;:7֢��pwc�\���٪V�j�R�%+j�ZC�"���d��>�!��OHuuÆ������G6+a�B��{��z�J[4qާ�\&t7�kM}���A�.�<��F�^Ց|��Z5�*�"�@Ѿ&��x���/g��W��B{�ا��>�| ���l�vm���9�2U���쒴uI�;%k<i9�.��,��o`���Z˞��移ڟ>f\���8+E�6�T��Q��ߖ�y7��{����O/o�<w��&��E%1�8������G։����հV_�Ýz&P	�X�(}y�ǽ��К��q��KW��j���^?Z�3����P��E{~V���ҼyS/z�>s�l����f���7��3��M�c�����3��g��>Oq�Շ��A#��k���^y��Xn^����<�߹�P��%y�T��Y�d���9ՙ�&���=��M��^=�`�r�N_�8�&����Y�Ɲ[�꧂�wl��v7�u��o��գ������.`/��99���襢l���ɳs��*w�u�V��kP-��Ĩ�@���zOΗC��C9��A��yT��'F�R��ǻBi���V�xp�}B`�o�h~
�h⟊�|�k���<���G��w٠{nq�wU��5l�0^�z������W���|ލ�؃���=�n����Ww�F�=�����ؽ���E��o�t]�s�W�w������`.�N�T�����$�i�7�U�d��;c�Z��s�g�bu�gh:;G�vK�.vuq��	��{��y���w}� �/��z��켑��;N�[Ŋ<�9כ��������W���%����Wo�ɝ�:�rs�ɒe���aӲ�N��s�+��T|�:{I���|+t��>ov*���W�Ϣ�����J�a���G	Uϧ���C�jqK�wY�L��z�h�{���J���=��޻���ίyr��.�x�J�e����h^ߤ���۰��ɞ�U������y��P��x{)�\�=�r�+�v;��NK���s_.��J��={7�3}�y�&��9+�����Gc��ﶖw�3w�z��
�mJ�O�M�]W�L�x����k��̘�w��}���Ï���x�](S��^��W����q��q�����/���w�a��~��A�E�䋠}�vy�1�{P*:��7-����2���\O�G�?���m5֭uL���[e2�O�{���x-�X�E��+|��8�k�gFVk��MWX�{��i��=84����R՝t��y�;���MYv]����2�7��.��j^}'��Y|Ү�&�im:�v���}��`[C:��s��>AGOۯ�e��y������a�C�Gx�ZTX��όO�zV�P�`g̍�����		q0l��]H*q�"�k���1���͘�Ф�>��~X�;XPX�Z�����'r�T�G��h=���Q0�<�s=[����6<ȷ�[�$f ���)��[uw&�o�c�b��z��`����l��DpmԽ��a^��/d�C|��\嫻^ �{)pT��t�1��t��f��G1U�6��YE�g7}"T�!�V����[|qe��AwC�ڧR2��|z��D�in扺��H�r��m��d��Lx���ON��=8뜼�2�{��g�E��ё,|3����ܭcr��oqغ��-�������+f������+F��w���w����qڨ�일��6V�o5�n���,��E�rL�_��u^�"mu��'���K���
�XD��`�v��`���Ә���
z�u�3[�����P|M�g u��h>6]΋��PA�x�9�y���RJ�Z^��9��ճ���u�w �F�OHC��p2�Ҧ��g���u�U�$T��1f�洭����Ӽ�� ���oGҦ�$��@{J�W�&R���2������2��C}P흊�ɗK��7R/8{��H���hm��Y�S>K��I �7�q%S�;;.�PrT���qӬ;u�g����@�ʜ/q���I�V�bf󎮍:+�K����Ǻvw۬���d�7&sbg�������ڏOP�f5�.� 庪fٻ\U-��D�5�(���ޚ{:է����&9���#.�eS I��{�ڎ�W�F�]i�gZ�^����4+��d��˫�����E=�g36���s���.<�篈�1���h�vi�ۛ,�>�V�:���Ⱥu#L�f��9��y��gKU�e����e��4�ߑ�Y�z2�5���������h�G��KN.wY�h7c�X2�]u��C1��v�(RC.����	����q4�Y�t�b�%��4by��"�}iN�����l�OT�칷Ux�Y�֝�=7
�[�WnI�h<�7w-�0��;l���t!=����$�պ�9!8��U�f<�#Ũ�pW�V-�k�nW�a�rY����w6�rv7uƱ��0��nL{���V���h����>��R�����ZYW�\���Z�YDqĘ!P���A"E�m�̠�2�FcS32#X�����iX#�V�� ۘULj��T�,�iTb���
�b�&V�,G
�����U
�q
�0��ر��f`�Tf%ciPU1
���m���1m�4U��J֨��(�Ҳ�%�aJ�Tc1��V�r�RڬaiAQh�\�r�E2�**�%h�-�Q �VTQ�b��h���n%k*Kki��B��U0�,U���eȵ
��AV��[s*2��ƭ)c-U�f%D�2�Z�&#��1��ۙ����Z%��V�i��m
%h�Tm�aq�pTQ[e-�����Jܳ���Ƶ�~�D/叹l:�#o�{-�(�.>�J'i����J�*���Y/IS��w,�s��uZ.�l�Nׇ[L�>���n��4g;����i�ؽ"�~�7;zu)����y�;��`��GQ^��λ��f�G�v����˼j�W��l`��ۖ��#7<���^��{}+ҋc�<�V��Y��C��J���g\�};�w��H:QwD�[���d��(��O�>�}sf�7��Ӱ�P�>��8o86X�;�Ϲܢ�i���,Ύ�������3lu�gh�.�a-�A�n�ޚ�J��K��L.���g�bL�8���'X��ttx��c>����޴���b=Tt����2v���ټ���=�,�D'إ�_T������{M��X��ϙ�P}U\���>~�s��&I��:�mDF!<{ޏ�:�Ϛ"��;�F�/��53����&qǾ̛������D��#�R��x��`n����=:������5���k�WB�pK�@a���+Ǿ� �vȱ�u�O��@TNU�J]�]���.GWP,o���3���V˗r��Pb*��63'�Ε�7�{f�]Kas���:���-��,=���×V�Զ-�@�Vo�!����j���YKH��������>���Þ܏ ��[��*����%�X�%;'Y�=�b����"��U¦��Q�uN�����dy1H^��I�.������I�W����K�՜����Ͼ�b�}<O�К�\�ŉ�F}A�;���_h�&������8])��0��������w�V~��wdW�S�VqI��qo�nd�c��xٛN����G9i[�_2���t~�ޤ��a���� �J�B}�.��z�}��׫/������}��m����,���b�{�r3~U�tp؞s���]����i���W��SAW]�Ig��w^��1�KN_�G��ԙ�������]^zK>;X���W��e,#X���$6������zs��zn��:���0ե)ٞ��{���T	M�bU��H{�PΘ�߆���)�}�eYRORK^tmx���r���"�ʋ˔hd�G�p�W\y|�vڑ8f7 ^�rWN6��]8ҥ@tw�Z���qmzEME��=�������tS����[�r"�_b�֤oDF���;��R�*��G��k�bԻĢ�_}U_U~���;����f�ܚ�l�<�}8ʙ��>��b���e��������=��6��Xώ�au}N�Lګ�9-�Y��*^�v��{;�̵��rc�x�F{�D/������^w<}���eZw��s֮(ߢ�m��;�侬:��a�vF�.}a���+��=��dݙ=G���M\�}ןJ�v��	%�ʓ҃�P�x�8��ǐ���qa�����s%�˖$��EOs�h�&��*L�݊m�����x�$y��Lzs/�U�w��~���N�"���-��$���5^}u�K�'f�sx�w��upO<�EG�\^�r\�����:��w�73Oҡ��L��5^�j��@�M8���}���ߓ�_��}��-�����/7'Z>������{��|d�㣦�͞�z��o��}�PBɣ~�Np�JUQ����7��(�G���1F#���h[K*C�
�KG��&�V���@��Y䷓/ ��@�p�7��r�Vr=�ծ��v5]m�R͕�s�KP�$�y���tR�L��uA-[��G�g��:Z|n[��U�W�Vq�-�s�u]y��ζ6�h��c7=��u�o�{Ɲ��ѷf��z�V�5���e�7}B�/;d����8�������+F�;�嫗��Oɓ�ͬ𘶄WW�
������ܰ�����c�k���7����䣒.�l�b ��y����^H��Wa�>�T��OJ�T��qY����G��.�%��W_˛,Ig���U�������X�*y��g���Y���,`;%��z����!�A�0쓡���_f�T5�3yܿmۑܣ��x����-ۺ�P���r�c��X;�^�ŕqD����s�ގ|���_s���u7��2<�99վ�6�߳��6|���<�}�����N�?�{�z�iBxyH�m��$�P�0��Ϋ���B�8��o9G�EOZ������go�� �=w�iK�/��{7,+���O�� BY������'o��_��Ma��UK�ϕhkZ^Az�ɡ�0�+I�=�[�7t{�����x���ǣ�m�k<HT�hE�t@��a��Y,�#uoyU�YR������P�}��(VF���}���Gy�;�*V�1�H��tM�=��{*��u�����݄��:�qAը=��o+pr�/�z,H|�>�;++��s��_9.u�/��4��Vœ\K��dr��q���#>�םl�VU�:]-������Eו{.�oէ ��'��ۘ�q�p�3ry�5=K)j����m��
43l���'�s�P�iךV�*foQ�k���-�~��%7T�������ʏ&E�}^ý��{z�|��}q�m1���fۅ���ޙ�O�=<	��:#�p�7b1%�բ�jZ��?�@V��v�}],i:�߭!�\/޳�$dp����wN�yw�,9�S���/�8����*�f��۾�F]���{G���KNt�\~Ͻm����
���3ɓ���v�7e琿u��תȩ������z	S&���r/��?w�L7���OֳV���ZX(8�Kn�{�yŋ�b�|s�y8���?W�H+�7%�g}D;$]�qx��])]Sj�vUU�jd�7ە�KΗ�W<GLU2�a�\�{��Ҁ]G����q��nj��o�|�\���6��q˴U䖹zw[�_ᙟ}� j�V߯y�ux��^۩P�g��6	Bf󼙽� }(��K�{����kVL��ۮ�ן8�3=A�Y�̏Ϧ����˒���6*�Z�Ż�z^y�fP�!}��_.}a���u��M��vC�"Y�ZɊ��KP�Ü��I�+s�d��7��s��� ��rV)t]yv�X�8<��B�{zdW�^?F'��X~�:�e©�"EZ�.�=d�`�$!����/n������Iqj�Y�;b��(���@ �72���� ��B���(a�uF?F��J�6} o�w��63��ٜ����l�v<�V���^�n`I^�d+�1�"Mj��t˪���RzO���fV��J�KV�$Y�6r�-��zg��6�,wK��Ap�a�bJ�Z�ꨫL�s³��Q-�Vk��9pwd�����n֡aJ�,м��L��u�Gˎ�c\�e@�{8�_�TW�)N���D�}Rg�l/�-�i��p��!h�=��c�`;i��{6��պ�=9��O�j�5�[-X�	��
4s�ub�뫽+����iX� 0�r�u��S5�)����Gx�3��N��}z�W^7v���v&i�r��st.��g�R�ֵLr�Y�IƦ�ku�LV��mfQ�{VK/�*O��^,~n�i���|>�Ky9�X��y1�U�t"{<�p�6/+�b%V`LtK|d��Xb�
,̿S;�7w!F�}��
x�}����b���=Y��p��p��Ն��q�/>��S���i�ʎ 2f;%7|�I�Y��F�(�9��d8��s�'.j�ڸ���0B5Y�7�{-}�n��jy�#�~Z�U3|����.Y.�;���d+��)�L��ACܵ
y_kM��S�8{vl�cC��@⯒�\��b+�߮]���ȑ϶z���Ԍ���3�w�[�\b)Я5�;�-���T�,�ڨ�5�\��KZ��
��e;L�9sQ�P�U���xZ��߅��zL,u��9����z<��(]��e#,K��x�w��T�|��I��1�9tb��/�Ί������%X�,I���$�j����tL;��D�JD�#���2��=�=`����\��Ѵ�s���T+���~�5��"��uˇN	��~��ze$]�t�u�o�Bl�RVG�_�i����;]���ʊ����"n�O��3�;ν��Z�[�c>ѡ�����MK��"�ѻ�L�t0�u!丶��� �'D�����ozk���vs������_#O%��`[+6�8�����B�I�O�p�˻�4���Gd�kX���Y��)�C���{���렅���꯾��ù�͓V�yy��ORJ�R3�>�\E$�|vױ?|��Xs��i+�_�f0O����z���h��u?v� ?��Vq�_��ٳ�UmYk˅�U�)v��Q1�-��Z�����#3���^� :�J�h�����pt�}c�V&��+�J�Ǎg��+O�m���{�&5{��Ǟ|�߷ڼ 
2��p|�x[�4�]/#]y��\��f-�Ϊf^����M-��%b�V���f}�]��������m,��v�L��u�z���n��k(���ֵs��KmZXZS���p�"�$����Ղk�_+�Zw�-*�~sƲ]5����v(�}�[)+\���=�"8<�I�<陂���-�[KuM����f"����88j*š��EEb��<�L���	ĎpQ�=,���fcO��M�	��^��Nm3�/rs*���Ml���R��>����&ZG�O
�*"�q0��ޑ���3]����4n=�����F�锏\�G��j`%�KH�i�׻�;��~X2�\/4��6��m����]k��'VGR�`+�5Z�7������5�����W�=hi�-�^M����J_��~��i=F�S:fkY�u�#�҇��*��w����Tu�<s��y�$�-My�$���=;ޫ�{>q,��'����_}�UW������cͷៅ>����g�Y0��x,����g���K�x�h��J#�I��x.Ӟ�o'H��/�
�^EF_��1*��'<�)�wR��o3b�|r��Û�o^kC3w2�}8��w�a���A�=���;�u�}//K�߃�11�����蛾�In��1��P��c$��G�r�旆�n:��1����K˅�^lU�ϧ�)ԒM����t�R�3��L%�ZHP�k���q��]�����C��^T]�_�����<{ڝ��E@�Ϣ�h����b�Q����Ɗ�WI���Hj����b��6x��I7~۷�-Z��r�.�+yFX;!��dv�ڳDP���=Fz�S�l{�eEP�sq�&����ei��w�{]v �PԸk�·�!�<���������"�7=�̊�Z�*hx9t�^^�Uv�s�S���r��`�ZE�=�=���&�����56n��U�{/x�c�dͶw���[M<�0.#*���{y׼ث����7SMID�m�E��=��Vc�Ž�\�~,P������M5��Rϳ�-�*?�޾��*��߭v��e�w�l���4Nz�&���z��| �΍�)�W]k1s��U�)�EY���r���Z��j�����>�o�l�/o����grђ�L��fŒ�q��VS~	�/�*˾��W��hw��y�a'8)��B۲��#��깵�����Q{�Kօ��j��E9D��mR���t+�[KS�̱N�(|�����{/�WH�:T1�Q��=[�vu[�	�n��[k+y
"W�	)ɥ~tb�=,�l�� ��h{`���3���4��9�u�ۻ^����C��IV������+jj��1\�k�yfH,3X��\�~r���ٞ�+�pU��3�H�`�.,���1ݛ�u�3��}4�A��ܜ�xZ�:�1�9d�u��@ՎD�@;�j䡰��y���踟N\*�Q��`�/��c�7���`�OLoV>&g�"���B��j$�E�S=}�C훑yjOh�%u1�wX��N��+���F���2�o��OȒ(u-*���K�zW/ �q�isoP�)'[k�l��d�VD�����;s.�9��w���'����~���m�p�{	5#��^��B-��q�B��`��m�����	�SL��X���f�y����qm��Qv�}]�H�~j
i����9��Gw;��b�P���ܝ;C�^f5ٲ��۝?{åDnr�o�g�n���@D�Ƈ����g���,��x�k�A���N��ħS��<��[����W�њ<qo�b�,,���䰎���
�<�s}l���*<@DKwj��U̘���8hO�1ث��zNS�B��{��\\.�^I$'��rJ.�4V����M2��D�ف���>���6��ۼI� �!������Ρ��h���i�e�a�w[}o�fа�j�I<���L��ǽ�Z����@��0o�+Bo5喎�-hwq�ꆹ���+��m^�ŉ�9�t���9�ۇ�G�w�s�>3��� a��a��4].�"�}2qo�+����X���{+邏o U����ϴOo���`���Rܘ�� � N��{p�VʣׅU�O�⼿#m�N�{�!�*=��2g�ݠqS��-ӂ��@{���c��Rc�jZ]�)n�^�*��t����F�Ϯ�J&��'Y+�� ��� d݃$�޾���y#�m���d���g���ŝ�r�B�s�ۗWJ��O����eЎK�t*b�Z�jͰbo5R�=�[�
F�u1��3 ,���C ��7���trJ�� $���_w ��q������v#Ɏ��yإ�&.�pby��9(Oޔڋ��Q�c/�p��{F�l旯p;w�ʘ�է.��p��eŝ��X��5�83p�j$8��6P�*gaSf)}�+Fjsb�Ǘ��ir �>yҠ�w'��n�g<w�,�BĮ_0{N��jj�	�*hɱ�Q:�������8����ޮ������Q$��n� ��}4;y�S�:��E�v��$�*��	�8>�	�����M���h°n����a�&i�	+mF+r��^��q�F4/vE�ֲv�x����-�bմN��r�]��߱�qP���|�mRm곗�G�5���8�kߙ�vM�l�n{Xd"-�]ѝ��R� ǄS6�<o�/��ć0*��k�c��ԩyr��tYn�kv�7�*@��C �Z���w'Ν���sE�Ɖ[�9t[���f=i7E���'О6�on-Qݹ����|�ׅv��D�b���i�V;.鰵V�}H�Qr}�&�ɑ�Æ����~�5{��^�[��Nw�{4�}��s3#b��!B���kS��j-Ij�(b�V6]�1v}��iDmYK!~{ }�A��/��/��41����n�}�k ����]��*~��9����(�� �t���e.V�Aiu�����E�*�G���sK��W�����FVvwWE6�}����>?D�L��R効r�dKLjb
��" �*�+��V�J��8[E��h�Fҵ(��k����Umi2��(���ҕJ�2�q(ܥ�R�
�"��+a�q�%���.Z�b\Lr��[)U�R�	X��fb$�b�8��V� S*+�b�0r����ffdS-#khc+�EH\�V���fJ��m�Z����r�Kh����[qTr²�aRf�fP��+YL�.�Ņˌ�q1\B�8�DJ�P���J���,*�*
і�TAV1�E#V����

�i-�U�m*jJ%`fU��1�Ƞ��Q[s*�R
�)�Z%J�%VEV�Q��Hc%�.f`Ȳ)��F[Q�Y�bʕ\b$�J���jc
�Դ�ʩX�\��YG�H}E2�4a���f����0c=�w4j�mY|�l�V{�^��%��-�/�Θ��ͬޭ}CMq|Ki΋����UW�&���;����Լs�Uɝ��Xg�޸st���2�̕y]�@����Q�:�0�ū��Q�W�=5P!H<��r���f�֡��,�pPZ���x��G:w��aB ����<'S7kEz�5�(���;���E4𻖯�a�l��&C��U�������z�g��S�c)����do��FY��y���h�|0M
��=�1���}�.��|#��3�Ⳣ_{��W{���>K����Vf�9JS.�?k�{�B��}��z��3r٘)�ŧ��5�#��ށA�
ܯ�<>X�W��v��e_+K	2ء_^���G�YL�r�к[��3�:�2`�n&]t�U�>���^vAx%e�aa�Ԓ���~`'�	6u�^h��NB)��f=�������
	���J�U^�Ok2��|�i����Ϯ]��S�;���_	Ӧ�6ְ��w"4��\C���vY���%�p6��3�/"^ѝ����ׇ�lQ�n��{D�5�󮸣w��1e��,��ep�[G��j*צ���9M]����]���y�Q��t��U�j隊'h���Fv E9�4�L���*�q�����QD�m)�D5�=q:�*��l#���.sۄ�v�z�~���꯲Bd�{�Ż��c��z��?G�8at��y$�#�'ڤ��9������H~�:y"�����=jJ���s��.5~�l�L�a�0�5ȒpN'�`S���S�O:���
�llPؘ=L���ү5�^�T�����J^��:���K�^�9�0_FB���~���%םqV�3�a��Ɂ��Ɨ���chg���˿uE�&Wj	��줕���ϪWV	��"�?x�x�:���LL^�^'��QǪ�o��Q#A�t����y޲8:�>����^%\3��Uc0��v�Ī��Θ��l�!��|�˱��AfĔ�7�J',<��� ��i�*X�e��RK��\�垇VZ���&uS����|:e�
7��x�}�gK����5k�q�g�0�W�o`Êަd�f�B�y�]i��u/��~�[���ɻl�(t���-́�9ٯ�ڽ��p�|�a�.K����B}|�W��,�`ءe�;��)��[32g���l2��̙c�s��P�L)�u������7�$닩;��w[)Z�m�5��h7]�^n�z6=�B-���S���:����b�{�O|��Mw�,��Q�r�%�-庙7��Tpg	hTc��EnoV��7���������k�_����� �?Y��o^X��T�T�睈I�L��������o����&���j���3S%�mzו��W+�jg�Ze�0h�N$py��"{O�Nr,�]w���/���O�=�tt�`�PںZ���A�#ir(l𻇍��e}��
+�5�*��|ǝ�6��V��}���4���Wkɔ�X�h�P	i:���1g���p��e���R��L�Tyj����ل�=���m]{ˇOFF��B����ybΕ�X<�j������C�Xi	�.yju�2:z�I�=��z�ysb}��eś����9�կU�݄U��iQ$��m��V�aiٵ<��ֽ//N��FZ�C3��x�+f'Z�P�Mu�;<�hs�ZV)�.�]�ݴ	�H�]ˋ�U��S�`��8;��쁋��\���x����*b`�/���A}Y�hty�7ᷪi���� ���l�ʕ����r�w*^	V�2���+�PuD3c��Ɗ�H�Z��x�TU�e$��v��
��a���D�γ<lH���VV8d>���ck����7b�!5t 1�t{ ��d�Fg��g��C&�y��t�kT��;o>,KvW*�\�\��󇨓hՀ+���%���	���q=�O7�]��V�O�}� }0~
�ߝ���^C�9�kzS#0wL	_�B���`��xO�y�a
XC5��D�~��{�w���e�����Og[�Y�}�if�,+fC��ή�O����nvIϼ6�������̋"�6�g��f�ۙ��ـ��ui�pX��W��3�5�#��:�3Zt�筜�-b5�G�m���p>"���������t�n����{���Qv�|��@�>�������X��P�VW��*yKèK(�لǖ��ol�%���ہ�z��hVN�������Vȱ���l���ʰ����E�B����$�V#�z�`�X5�:\����=�V%�A�c��FF�pT2V�M^��}k���3S�T!>�(KyD�yъzQ0�sj	����oL���=01�T��=�\Ǒė��0-��l�-���.�����V9�᲌V�k 0�,����ܩ�����Z�'ì�ݪG�E�+��>���ꏂ��`]��i�t��y��w6���W�nHA�f�Oi�"MG�Vi����'i��*�@[�����x�%�����Uh��>SJ*Mɇ&,�Uq ;�mIՎ��VӺ���JBF_Le�jѪ`�_D凮�p����Ŭ��g� |>���d˭u�9�O\9kj�D��65rP�˩��fh�iLt��͡u�%���֥'�۰zy�g�[xg��+d��o��f͂:�C��Y���e�k������JX�mL��2N�h`�,k�ҳ2�Zxȯ��#��D�Wz�5�����%3LJ~�~�|ڻ��zu��$ձ9�FEq�]����;L�0��>���(�˳�-�#����p�/�X���Bs�	���{��~���[��e�|JZ�W^7=;������^j!	ȑg�F�k�s�/ﺇZ�t�lk�·~랩U(f6룵�C�W��n��Ì�]tFM@^U.&(�w�o覞3j�,}Xh-�=�X�z�yw�̻��vy@��[�O�ۄ^���{T�����Y���t�l+��t�:�ְ�/kO��<��pLU�e{��{�>�	�'�h�au��l�G��Ssj�����.��F7-��K^:\OT�P�?�X�ba��zxQ&����Fw�ܶAs}��ee�\띏6�F�
���1�fb�;�I�FY�bb��xiL����Mi��y�jx�w�-r%�1�c}wG{���\ob��׼+R�]w[��!^�ٽ�=�>� �b�(�9�pe�����Mq�o���W�E�������o�v� �d��(P�63h�2V)ˇK~^3�:�X|�U=���ҕj]����t����-#Cl��k��D�_T$�u�Y���9NzW��j�䙕ݷ�Gʰ��~=� 7�u��u�:����.��w"G��;-�"vl<�έ���F�ٯ��k��ܳCJ#�>KR�l%�vQ.�D�~R��c�x���ar9P�܃��/;��z�����Qt�y}n�	��I,!�A-�:����[�,6�x=yz8eIzt���)���cH�9������%��&Y0�(���t�o�򑜞�{`�hq�j�r��>�3�ds�����"�z�yz�����_dĝhL?M���=[���e�f�B8|O��v��Kθ�x5����&L�+���c�뽜�|���O�a�hJ�����v��\C>^Z)4��Fx������$�|�O;��:=��_��6]�r:$h7%+.��uҶ���-yh�J�g�)v�ݩ��nʌ��Ph�Ew�1s��Q�͏�ZK��^x��y(���7�]�]��z��=N�r��r3�@�<���xm^<݇Q�&���ji&���ݸ�o�S��9�=���:��M��[�tp�$�y|�qc�\�稛�=�S��}��	�c3dp��/b�$�����%XLƉ�2N��NXyV&u�f�m,uKΥ��ĺ��s7��q6;�+qOΙz����#�;	����ݺ��"�ٜ��y�#+�u�(�������o�:�*1�]i��1��0��{-��n�=�*<q��5��,���y�����l�K8��S:�E㻀��"�aŔ�`�	P�3!�f���}Qsv�Y���@2sѷF�XUf�O�`�K��s�x��u�����gB��]�ɶ��	`�oU��h_W
�%�vV���°R��F����y�]A=��$��!���'Q�^#�>t���%>�������{L��kY2�����kƃ6K�Cd�5�gM�����qѭ�G�z��ّiԬy�fo��FOP�6=���Tk&R=r�7�
�%_%�ͪ�����߈��D{U�r�E���XY���&{�92��^��x&Z<p�SU�svʥ�4L�K��A�!�X[Hu���W�u�3�zm�Ny�^���j��U��їt�B1�w�
�7h�g�l��%Х*�0�:z!�ׅ��5��+,[��M������ii>��Ub�
Pξ��Ǫ_O3��؂����K��7���b�Y_�D]�bxc�4�Y�R�ܿ������-���pX�8�����W��٧'gw�Ξ�5�T7�e k�(�Lƶ�����N�T�}�	yzoU��{���us[��G<��؅��S��ז�4�KB�.�����5{H�(<�_e6�C��o9�����o��.��P�a	���B��\l'\e໇���֗e҆Q������n~=[�L�P��J����4�WާTC=d���� �#
�*;�����rN�13���Wr�?ny�k���t����(��B���4�(�(�ݪ�b\8���׵��-�pY8�[��G[��i�T�!C�c��pXOe�&.>X6��,�W*
�k`]z��__����9�*��8��L�,�S63ۙ�0'V�q�z�ȕ�cv�^�ydC�x��:C�:8X�n/�Ѯ8�#�������]i��P�w��^퉫g@��_uh��vG�l����3�\[�bX��U���v�uS5ݜo�#x�o�l�:�ΝiO�-���;�:����+��ʱ��*�X�2�biE)?g ���󀐍��"Ί�f�wڱ���{�2��OH�Zz�j�ڮ��20 ��������V��{�x��龊�:��A�=X����ӻů[����J�:WGբ�_[�����c��Qm�y*���z��}�o�� K�kϏ9�L�?����
e����r��CzVϻ/�ϔdhv`�3E{�cزw�3���#�R�������J�tb��L<\ڇ��l=��ݪ�$LOG�.v4�+	�Z�+��*�D������j��F+�塕�����Ij{7"�K��9�AbbY���F�����@�;�au�0.��Z�����5m�oixϜ���r�D:մHt��5�����e�L��iCr�=�4�����K�Ue������J�0K��%a��L�7�=vE:j�B�A�1��TE:�iu�5j�Gx6[�����6�wx�O�ғ�9��1�>��2�o��H��~v�Լ�'߰2춧^N�x;�}[� �%����Y�s���+"�+�pHj0�u�2,�Ӧ�o*�y3�-b�Y�Ƒ�~v���uQ3�Y�ިm��0$�IL�rf0{�0��}�eY�����͞�y���oá0�>�@� �y���x��u�s�Y>J�o|6�-���~��ћ����L�_Z��@T� ��_]x&��u��:��i`���MndM�V��*� ����׉����u���ۺk)��f���Zk
���x�x=ӛ�f�C�Ak��m��$��p[��*�.���	�8+�V���:�'����1�7r�2�`_Ӭ0o�y�&�|�g��0�j�ӣʥϓj��L���	��������߭3�^����I]?�Wr����E�X
���v��$�]��\�׻�b�X��Z��ڇ�}��bqYӞq�U���i���f����Ѯ��f6�	-�l�:�q�Ya��E�v�u��-���b��ɮ��0��O��agQY�������ԕ�_��m�U��*�&�C/E��<��L�r���ߓ��B,�$d�WrC�j�������8}*���Ė�/ � 7Ꚁ�_!�߽a¯ڹ�NL��K<��C:��k=�>7�u���K�CamB�qx.]���ȑ�ӑ����w�L;�.��H�Ӽ�zP���QC��A-K���[K��;]�acp���˿k����XS��(���l��ռ���y�(]�)��ԫ�Yj�.�γ�H��0{�[yp�?;����:�J��\����r\j�����e� Ef��zn�B��u=J��a�Vm�<Jk�����Ȗ���*S�Gjuw7�CN����9]p�BL�h�����7)� Z��5��(���숎�\_f�Y��8��]�o�9ۨ�{]�Ҭ�\�^�Y�m�������B�1+�A�.���hj�U��É'q��(K��dO�_'����:�����x���m^s��v60�mC����K0ю�ӄd�Hq3��n��*+c�r�_G�VN�0��[Ǽ����ۍ�l����t����lY���\;�:���P���_][�z���_z��y�
]�ۨ���)�t>�頑�ZT8)e�!�{�/�"9�=�Ȭ���Ğݚҹ�~s����` ��ջOC���=��p�Uck��'�	Q�Cx�t"�hΦ��F$>A'�\�����G��,gJ�e����R��v���� G�V��(�2�����q{2p}<)^�4
u��@T��w��}��qS7h�{·k�G�Vⴍ�E�*�"t`��&f*<L���Wi�逵���[dn�K����������	��}��Rn�
�7H�6��p$j��ZvpT���:�Ugl@�[�28<|�;����Q�ʾݘ���uc={�x�=����Fl�|��֎Z�x1 7	��>i���<�@�L��R���)�&��R��<���b�̚ש-9���ܺ��:��e�{�6(����ܠ�][��`
!�M����z��nRo7M�ZX%2֑�C�ʠà�\��j�&=ܹʟf���k��w>�sʿ�n��{�7�d�{ڌ����QQ1���̠#U�x9�$�ӯ�i�0^��JD<�[��)(%qǻy����	@��\���֒��{:iWK���/�+��,2�U�z�˛�W�w�^y]�[kRt����=�).R�Y�����(s�x_8�i�i-<�Y;[���2��na/=^u���d]�t�&�%���}ҮX.q��MV���㗀�YǪ(�T�����F��˸E�I��4dW�R����РegA#�gT�B+)�EP�s�9�YDQ�v�����lH`���=`�:|��.T:18Yy�g_ao	f�u8�̾����d�{�]KQI��쒅���O��7<nܚ}z�\�䓵mT��9h��5�za�ES_hݝv[7л�F���n7p�I����s�e��B��[p�ʶI|�ȃ;�kz��0���$����/��m<6lV�h��ޡ-r^B�M��ӹ��w)k^%�7w��ݍ`��<� j
�
���U�����ƞ9���F;lЋ�e��9Ω��@��E������=�A�������E�� w�&��^g�[Np�{0.�~Un����&U�}��p�p���C6<vh�y|��p�}qД��i�	Y��[�����L9p�]dq�o�(D��}:(>b���G��"�B�IU-*���Q�Um����*��(�)2�b�*VִV
(�(J�[m�fd��.a���cr��H����WF�33ak`�q�R����*���!R����#1�`�Ĩ��hVE��(�.*TJ���P�*TE��ŉ��l���QV�T��r� �+Z���k*�*$EUVc�m�U�V���Pĕ��K*1J�*���+"+��Ad��R�IQb��[b�Q� �,�e��T�fR(��j6���(�1����"-�j�V
��R�mE�%b�,kA`�QU`T*�V���-�iVز��e�aY�`T%@��T��a,�`TR��EA�T�*T#Qb�B��Y�U
�V���~�Y^���&gM]Gxo�T{w������
q���gv���7�߽�sFyo�U���oN�h��y�������>��=y�J��'��$�<{m
�������g��X�bU��ՒT��!Aذ��9�ۼO<�\�����%�AU��Dq�{��/]&�����=RL��}�!�8ޣ�����e+�Y
�؜�	��RK�E��\E$,�����M��j4�e_j���=�����\c�`�H�nJ^V��>�E��}^Z/���2e����>�L܋����泺Z*ƹ���&cD��S$�D߇�*��;ּ����{}N^�=�u9�l���0V����2;�3�X�plyǈ�e�-/����祪1�*E���c�w��u�fQ.݌��Xۘ��v&=�cb�e��޹-$�P�O�I����B����'ٔ��-j�UC�^J���w�:� ͻ,�3�P��]��L���*V��r�XD�c��9��z6͊���i�0{�)֕`c�j�T��Є�k�����C��o�g9��7s���oW�&k�ί�e��KK���}),uP���!Q������t	���J]�|iU�^�����z�ۙ��@��}v)wJ�U��b�p�c��L�s9����{o�:;��Z��]�*$y��jT�-��*� ;ٕ�BTS&QR�.LdS��5 4s��b��o���W.|��  >�QR��&t=x�l-ic��}���{L�kR�:���kƃ6�]Y�m�eU�d�zn��V��w�<b[�*��v#'�i�r[(��E�w�-ܖ�k�kX3g��7}�7�h]|N
��[��n�|��33�Ʌ���2eoz�L�ڢlAb**҂����*|�,�4=Ԣ6P��CO_�i�+fME�i���.Ny�I`���}�����ǖ]���~��u�.��҉]S1���B���Nͨꥨ(���5����R������pw�YLB�}r�,a�C�"�MB��ls�"������bg�Z�^\.�w�4t�ʄ\�B[�IR�C<�y�<Bj������;�5��>s�Ϸh�0����s��"}����pu�\~�����jJӖr�Z�h��Z�{A��¶��ex:����`J��a���COR���i��5nP��[{��}a� ��~�=R�9�}��zU��]v!�>�9-pP\����i��pўӂ�gu�kCyPc�.J׊z�[�ޣ�}�RFIk����4�
8�`�	�]�&�R�5� ;�M�C� s��]��\���0$&f��{o�|(V۶^:M9�7��ː�<�­�I�hCۭ�W8Z�
��,wﾯ���}���=vM��I����gA�0�ڬ����E��L��nd3Gz��g/^�T�rwױ�{6�х�P�dK&����i�cs�}��F�|�+�F:�| ���w㾸�چ���;���c;�`yb\�d{:\e��2��Hy`Ci���~�妵mi�6�y����=����,�-�fp�3GC��8�>��P��F�+��o�Tml�Y�;)Eݽ7ɇ��YB$ #>����L�������C5g��������������κ>�G�Ұ�����*B�;�$���3�Ʉ9�'/��ob&�!rOJ����G8�o��\l|��F�\dY�U	`UQb�����"����C�,�z������Ξ����c��"ĳCmݣCz�b���@�7ٿ�ʄV�=�l�]+Y��^F�%� ���s�9�z��X"j�D�N�CW%���yB��^}�8;�5��:�΍�K���i��Y����<}��38ߧ�̀l��!}�5�P���B���޺�3̀�v�i���E�]��͓|U�����c��x�F�����3�F�+���K܊�G�ٔvPX�XKZl�jZ�q>�/IrZ��+�xMN��4���1�f�HדQ�R�w���x�	�}�3k�V�'�ڨ�^,�,���2OϪ���*�>�'��V���N��\JIT�}%�~�cU��dW��.��%��rL��J[��t�⻔�&K�������NW��r/}��Y�G0#IY~]�^CVxK���g�7�v]˛QodXX�WF�	�XD!¶��R�.^��Qf�%rT!i�Nt�L'r:�"�*��qgӼ/o�OZ�"���*���{��.c����Zς/�Vq�9�gJ��N�%>��t���cVN��=�F�:�P��ǕK����tq�#h�R���ؽ�s�j
�^Sq�x����y�$��-�^��w,�r�^5MhBx,n�D���Pɰ^��'��N�fj�V�mH���u����0'�8<��p	����#�=�(r��m�������|����m)�!/���A�LΧs�՟Mw���.�K����r3�e ��`�_�cbX�JK�	u=J�υ�Qj,��+�3!��UY���K�uE%-��|���L�υa�7؋=),�Ih���{K�	��\^���pZ�ʽ:�({�C���ѡ���B��$�N�����\��;�C�6�fϬ;��a2n&�f�ݑ89L�U��79��`�;���}���V�`dN�T%4���m�ӾW�0�e"vRr��s�����]&*t#��r�^6�}��6_{$mi��V� r���=ɛh;��T�R%ʋڤV�^Ht;�!#�FSW���XS$�x����3��5�6
�Y��C�Qi.I�ilRĮʮ�Fg��4;��u��^7.��8*;����=���&��^���;ÍB�\�Go�v���'�ԦnQ�/���U�Y�T���z�8�sW�ۇ^�*Ƒrs���d�<��-�&������fl{�7����D׶�&����^�6z��S�\��W�Kʫ�+X�u�Qg�bD���Ǔ�M�n�s���na�h��V(˦G����׎⭞f|�|8�������a��z��>���P��O
���I*)傥q�#idP�,���r�xhNHߥ׷V�1�i+.(^Ev���4R�˰�w�$͇C����l9�&�B�W�o/u�_>9ޮ!ꖟt�V�d��&cD��CL��Oe���^5�+���=k�{�Q���V.�(�-<+J{G�gC�%���plyǈ��az����ݫo��{��U��|��q���M��:�Z.� ���L�&����{ZX/�x�[8�Ͱ5-�T9�1
�5t���ȷ��]�R�Sa��t6�i��n�N4�ne�8��`�[��\RnZC�(P|@%2�-C���e
��1�}UT�3|�~3Տ6��yZ�q}��&���Ͻy�m�gֶ�nXس�:l=�����`ܠP��S�y���K��thu���8}>Kpȗ%�/	ڽC�ۮ"wa��O.��/n�[�o��2�B��)���~v��]+4�=��b倿�0=���g�����x�����n֝$�u�e9x r����	�goe5Ex!�t`�����5s�h���i�70�W6�@_R�2%�������qc��jZ��V�p}�Χ2;�)�{��ҽ�*����DK�mR��h��}���kaJ�a�E}��f�O��Ǜ� Z��-�a.#�#��˰�
�,��~7~��)ƶώ8��jRߞjֻ<���Gqre�Ǩ�s6
�	q~L����&���A4o���Y��<s�,��^s�fK�]����#.�����]$s���cYA2+��A�==\X��Vz�<�'��1�Ӯ��`^Y�+lܩ��A��@�:E�t�ywg0����%kk����qV���<^��[��u���/B��-���n��2#+Ct-D�!Ы<�KDv�0�1�	�ӿ���(➮F\���s����ᵭL�S�u����`�sv��Έ�����������{��a�E��9J�����s��-�;��o3�{���yzIh�P��t�H������P��`�,<���f�#Av���M�MK�T���'�����3�)�|�<���FEf�U�NHi�8%v�̺��튖��3���=��ۥ�Hm`��w�+ir�x9��D��@j�Q���=Ig^�����y��}�ǺEzG��"�C�dk��qq�d���:x��c�ϵ�a]o�f_7�ͳJk�-z��0��o	ӷ�*j�����K�<=���P�'���=���l��8�î����j><�^	��޲���x+���<f�-�-�GWy~-�z�S�'��q�F}2��Gݗ�ITG���q�3�c�)������ ��FN/��v�d�y�%������*�>��"Y���g�#��	��m?�m�ޯZ>(M�X����W��3�׭J]hA�P`��*���}�{��Ʋ��뛣GI���Q�����;8g�dXtp->K�q��5������eΨ2�))Q'e3F��,�'��U�e��H�8�;��'y�*c.����v6�ZK�ާ
��4r!)(w|�^��̛Q�'#ݮސ��Q���_]BC�T����^pT��Y9w#�	�*�k��� � o*��d(T�ײ w2�\Xnc�?�z9i����^Γ���Z�x�@���Z=>�7L3%����;A���7�OLN�W�4�뷊|a��a�bY���Z�u"ŕ�ł�f_���㈘����}�W]��u�-��{6�ȸ؞�9璘��/D�"D�v�������e��m�Z}��g7Ã���ɗ��j	Z���l�8�^�s4�Y��$��~��a�ChGs�m��}�(����~|L�=�O�?-�B���iC�*�t�5�	Y�=�b�$U��ˇik6�anz{f�������!}��*�.���>[���^)5��s6������)����sE�po-�k!�pQ��6<:E����<�<\����Qgt��$a����{��,!A�1��)5�$�t��.���K�gQ#͜�P�g���c�Y:��Mo�+4{�n�Pk�·,0dXג�Ҏ��߄��l�}��L�o�T��j��LxX�vQ�y<B��]1��覟_P�̿�����y�$�e�+åw,���&}�͝�[t���gr��y�:�ύX��(1{ټa�ոFQ�6���=v�a_l�1��/g���w�yy6W��W�w�O:��3a8�M�M7^e��3�^擐�a�w�cCz��Y4��P^��H9���R�*����d`���\y�ˁ)_G��.r\Rˍ7��=W+�Cx���;jE���]x�	�gK���P��������]���[w��#���&6|��ȼ��:�I�7��<v(3��f`�s��z��]{##�l�EP��3k�=��ーk��Ƭ���߅T:�@��������
d8������a�%$��[�ʳL�N���ơ��!�V�c�����i%�1rɡ|*Z̸<=��;��9�N��Q;eH����'-���,kX�@�'�H�
��R�/K{���=����5�[Vq�][���Byd�FX���s҇5��]�&aQi.I�=�K�k�4��v��<���R�=�]KP�9sW���=�M|�׼����į���mxා$�tZ��Y����B[�ꗷP"FIk]�(t��L����^Snz%X�.N~���+���RŚ����zg���Y0�ð�4:R$�#��B��}ƃ�L���.`��*�ECW��0�阕��'ts��V!�w����90T6&G�M/T��VC:j�u㹰�<�<�jv���C�k����w������D�4F����v�Ϸ{j�}�wk���W�������y�}�;�]"��u�pX�U#T�q)n.�X�-x-n���.ջ%'��v��@�.@�j����,{�_m]�Q���)���S��׬�~Q�v��x�mh�,NY<*)%])��+~�eM���B��̀o.Q֎�!�_U7� z���+�(��ܔ��<���L�৓�U���̩d���z{g���Br�ޮ:rx��Z+\�V�cD�S$��D��ʱ*��)EXD��m�I�^� ���om&V�
Ҟ����G�PqqV���c�<GX^���u�<�wjx���N�H˺�M;�V��+V`�g�=y��ۘ�]i�7,lYLM�ۆy�z*�z�w[j�(��=�+��N��8}*��2%�	O/	��ە�@D�ouL^���y�uP�PU앗�Éz��n�ذ`��ڳe��X�3��N`H���%ܞ����9���-�Iͺf`�/�.[�qw����c���у�/�tb[\�ܨ�����eIZ\�#�y��,���`�.��g�^�-3�VZ�/ɓ�0�>�����n����gQ�g�*��e��b��:я��a�������P�������J���4/H�rd��e��j�k�}�7[Q:�.����B����4;�:��ڴ_	�ƣ����n�Bd����:�un�D��Ho}���q�b�+V������%P��� i�p6���@����Y��ʓ�h��D���[���j]v�P���1�H��=/���q��s+[���j��eb�ա��d��l&�����\6����/{绗���.(�p��]�LXW[���\\�F{�>�-�M=Q]�e:IƼ��Y4i�j��=��ȱh��1���o�JQs��V{AS�<ޚ���`�;i���Y���-.Y�K�l�����Z}���z�񱈽H���Λ����[0Q���_dmɡ�^:����E�qG���1R캀�Y��U�2�R�Y�O����f�ܺ���h��}�y��;2{�['R���z�e��62��&�yO�B'-$��:1M�0Z�b�a��wh�w�/�3I�/粹���jz�did�N�`�����f#���H�1V��|�Q��׷w��)�G/y@Q���
��z��Gn���\k:�4O!� ���Os����X���S7��ٕ��VJO��JX}ЕX<y�oc��`-ü�y�e�ƀ�ӡ��{�hȂuy:]2ƥ��j��^�����+��T�>�ݼP]7���m��'��R�G;C�-H/(�$���D�O\���\��s�[�^�aa:�G��;�GP�1���ؔe�T��)�V¸�kջb�ts��
\n��\��}#��p�]H�y}�:03��}��m4�Ε�,Յq�t�Or,�����57Z��b􏱈2މ�'p��<��Gۮ���0��é�� �l�l	���M���p`}�9e��z�$g��yKB���{5�7Bfi�
d]�x˛�k*g�k ��Z��}���Vgehs+bJ��&¬����l��ږR�u:�ۨ�5�S0	g_ۦ����X)�v����DFw�}�	�SƸ�s��+2�)�ko�:w�!�L�R�ܻ���M�I�z�È�b�"v,���u�:�<h�ѽ�5L5��K�`��h�^��e<<��]3���0v�K�Oڞ�D��y3�8�`���� )�M�E1K�ǆ1E,رRx2r����Y�5����� ��pe>~�.x;~�c���൦a�%BL6)��NR��-י��
K3&#uyb�׍�#T�5�N0j3>�Ұ�w*j5O6�f�(�;|T �Ѭ�u!�ܯ2�C�Z)��Ǣ�0uћ�܋�H�_�{��/]|�?#����f�IQ��Z�m'+WCY���{��5�_�H���W��ZkE��MENܭ[�U����f�ʷ��(-�N�+���k7O���XtAk8s���
�-�p�,~��dv�r�Ö frV��݋%�&j�v�&�����
����|���`���b��+m�
�c+Q�E@YX5)m�)*�ebŕX��TEaRX6�e`��
VQ��h�XҰ���B���Ybȶֵb$YP�
�[`�)+ �V���XV6մ�QJ�!P�ȃE��V�4��d��PB�d*���(�,�`�
c�X)+�J�*�+� ��U���E`��Q`�c!P�U*"�EE��dJ�e`�b�Ȣ¢�D�R�+R*�()QUh���X�
�"��R5�Um�@����Zd�U�kB����U�j��A���²���AJ�+R�
��)U��*�m"�b�kQDV*H֕��D++(�@��*�V*�Ҡ�-�[l�RT��P�DO5�k�e$%:�	�C�1��h�Ki�FnQq���
`sfw	*^��`�ѮwX��iB�޶�hЍ�!V���lCt���]S��䈀X;@߾$V�b����X5afo��&�v,�o�$g���(���N��N��r�;,�5�:Qx�A_ ��w�1��N���v� �z�����o^/��O���b��}���f����J$�1�"���]��f)]˪[���x�$��J���Ӌ9xOT�,�R��0Pv��5�:E���߫N�4T|�.z��j9`���Z:���`������
k���0P���I��z���.s*�>|�f��+k2\uJj�3�QyX7zј%a�����d)�<%uD#��[]�j�����fgOE�VY.�C`�O��'�n�D4y���s\E��0%~y��+,�̬d��Ǟ�o�W�P9h�4a���զ�ϼe�K�Y���0S|k@��[��@���ٛ�F!AIݐx��>�@0c��LS�j��>+��ˋ�������՞v��JϰU��'�ꅅE��MpX�|�cK�ع/}�7���#]�G�m5�Ǻ�)f�ȞhS�����aM��ٕ-���ϋ�,�W����n�(f��V��C1-�U4�m�z�tԔ�i�y{�YO�nv��Ol�����z��+�7���f��o�;��6Ԕ�.k���{c�5 c��k�!��-���I��u�P
I��՗�Ǎj3�zdGݗ�`����Ms-+�g��u�>�+��dϏ�(��>�y��u��TXCU�����ĳrٙNf����O�����eA��s�3z?{���3���ϩm�i��`P��+D�}��[A��S���zƧp��=c�������|=�ǃ��FF���~ı�J�Uh���U����<��1v]��=��훈	�-��u�:�C�l=�&c<pV�u"���I-�4�kZ����<���ކ�FI�m�@�����߼��0�Y�`�ȹf���ݭW��E�x��,�d޺���%�]�{'Kڳl��o���nmi�q����L�k18��b"D�.�5����r��z��*����Zg�J�8�O9υ`���5y�߇{��k��/UW���]t]ϫ�˚CG�=��Wp �٬J�-k��3�;����ht�<�ñ����ȯ�f�^KnQ��^�G�S��a}�K0�$!��t�]uA�����^)5����+ �����ʒx�����3��8�{���ͧ=��-[�Z7pe� :J�e��&���?J��gj�/�ώD��&E�
�G��꺽E�ܛ�?�����p���Ǽ}�l~�2wl�aSM(+�-S���>�Ytn��7:u�p9�L���LW��}jNlK�h��u�[��K���7֢�,�dv+��u����V^��j,Z�κ�u�B�v��9����Se����I�$�t�˸q���΢F,���p���sӴ�ՓnkƽY]���C�3��ZJ�త���+ԽҎ��]h���&~�{�t�g+�r��r��P��[�}��qE�_y�}���H�&[ҽһ�w�Ĵ�d�"�y��~�k�{صv�Kܳ>����+��㶤[�V`v^��'�9������*軫ڭ��o"��VR�^D0L����W��(j���T�`�ؠ��ļs��⹎FWt��')jY�#�j�}�
ëИ��Xϥ%ᄹ�T���r-EY��\&�ړ9fM���=JV�d'�?'�C��d�������Ғ��Ė�J~`\�1�A�e��d��t.�2J'aX<��E9	��z����L�A��@ꠗ��euY~W�hq�ǻ�v�{���~�u��n$v&.ibzw��J�w,�hM��];A<��w��)�p���ڲz��ޅ[m�u����Xv�s��.V@�羱.-zy�Wuo��q�i���S1H)�G}ٶ�8��TGUɔ�z�6��Qe�쎿w��f�C6�����)�X��7��iں�2r��Y��beQ{[�t�t=� �JZ	;�Ȯ=.��pS�5yO\#�,��Ky���2q1ҧۆ���ڜ���Iv��H`�\�A{�֙t�ypSn{*Ƒ'<�*��ii�ud�f�g��t�ǖL6&&�:D����B�������z��S�\���wLyo�|qtΩ^~(T�(��WC�/�d8r`�lL4�t�ҿ�S#�X!������r>P��
�"�nC�%N�C��ϥ����WcN(�юX���a �q���{S��E���3�7���k�})5e��-%`��y�M�	�yYA��#e�Ѻ��<81z��>�{r{e���Zk����5����,��a*�LƉ�2ODN��bם{w��]��ּ�`+|��=��Ȇ{h[\�n)���]�b��L��tO}��B,wg,� +���	[b�ZW�J��_���?��k�3�������z��}ck���:`��Jo���������$F����8���3��Xg]�LBf�"�<7���9>&_}�1�\�v{:�kOw=@m����"�}�bTk��x�=�B�w֍[�^8���y��Sh=���<��ӕh\C����[Ֆ�qT�L�'��	��8E�f���[K����v�=j\�Cr�Wh�$��*=���˨ş�NH����*��;��o�����0������S�)J��Mՙ���yJ͓�-�g��t��N^	�z �z�2l��)b��M]��䕚����.��o����[�./PUOi8��
D�ޗ��`��{L��kR�=:�1�>�u���R��aK�R����F&ZV��f��،����G=�)��ϣ�~f(ɐ�%�	��_]���Zi�O��Ջ�c���,��7e��k�gM�s�����K�7ӧ�k�3���
e��h񿥚&�:Q+�6�]���v:�=G�ߞ_���;o�OY�4���yN(�=P��0v,3a� k�(��T�i��j>+,��|���U�c�=^%�Y�z��K�u�	yzYq^��19r�,�<�-&�&�LZ��6ڷ:n�O��V��l/:�ر�cY/.��=�����*,!)��v��-7��r��c��33��BƼ�����z��_�_"���Fd�0����rCOH=���ļY�N̳a�s�:�l{��>,x>�Χ2��Պ�t�Qpb먚��"��y���AE�[&�-+}��ؒcy���vg��#\�أkҍ���3���焞�5kw�%�����Z�1��d��9H�g6�co���t�1��[�"uXv�'�׬��WLw�!\@y�-�Giǂ�D<�"ָ�c�`J����=Ph���_��w#�G��SR�v������C\��=k�0�\\%�9㵼f
�C�/6{/ڛj{���GD(�d�L���	�nmÇ���Ֆ�(��>Xe��YE�G��a�����>�z���c\=�f4�M�� ����^���c�\h|V䕋����l���rw���i���G�ZdE��zf	.����5�|�d��3���\�)E�^����)���d��%�ܺ���8U�-.%�r٘)�þ�똣^}��(u"n��[v�ػ.A�����h���5m`����(r�A���9��Y��󻜡���g���Ѭ�����r<6��e�n��MC0Um��R��&��D����_��y/�5+�y]��{]�. ��Cݓ1�8+q���h�+��Uq�.��U~��fF�VN�k�*j���1O>���a�6��hm�v�Z�E�+����T��}ۙ��q���������+�V֘�("��)6V��h$7�+�&��\WG�E�y.���.����� ց�7oWh��4��1�$$���k�ʷ+)u6nY�m���2�a��6�'���}��X��:��ɗ﷨~�g�{�<���رO�{��_�a��۳0
�'�����-36��/y{�BZ��=-�$��������)��-��魕�`N�u�ܦ����q]Y�����v���L�U�EI:���d^;j�e��w���d�!�Q$\]��3��Cޒ顝%�~Vg�2��${���d4����SoV�d�g{(�t�$!��b����|�xԉ��`�`G��눗��ه�ު��\�r�f��GY���2�À?F�#�]&v]e�3~Xl�΁�����С���7k�kG��*�I���$���KGM�2����΢F�8�¯��fM���g��+5ό5ʩ�=f����(ѩ:�Hq�T�^|���p�_N��1jo�����,>�d^z�ɝ�׍.:e��a+Ρ$l���O��6- o�8�d�AW{�k�yx
^ՙ�Kp�^�ڑnuY����0'�/c�E�z���H�+�\qyY��}�Z6m�C�Lz%~2/:�d{��v�Ϗ��rٛ��.�#R�%���b:�wk
뀰�<E.�=�u�=�^<��3���S&ng<�@�T��9�1/�`���Վv!�+Q/�l�a^+ƇZ�BB�)�Ғ��`�m�o���2��QR{։�5$�l�}l�`j��
��;gvR��r�n�Ӈ�}W�v��z�J�{O�	�^>⨽��S>��R�2
����o�A��)#�y��^�:�AL��9w���x�]��p���m+O ��m$�̯k9Y�q��2H�*�9���D�´�y(�
�:1\S���rޮ�({�� u`K�H�o��H�u�h������''A��~lz|����(O,�H�zw�ȇ5e����	�V��q���z:�ӷ�7��x����v�U�Rt��N\����=���+\����X�t����.��k��ZG}T��4�B�;}i�a���^��Ҟ����C(Z��t�^��a�:�ܦo��d�sC�"M8�����*!�����'՜�yTި}�)��k�2q�=�!Â`�e��}ғJ�S#�X!��;��ց���FE�{��Lo�Y�\��Ev4�mh�,NX'�Cs ����j�5��S6�9'��qW�kܻ�7i�8;�����Ev���4��������Ɠr���.YEo�i�E�7�u�9/s
��	�ր����[m�c��z/��f���v�Au�;w(��3ԮM=H����_7�t���|�9�%�FU��a�d�_j9��Wy��EV�We �-*� 1t�j������m�oV����$ޘ W��KM7\�]�7O��n��^w���d���)k��`ۄ�UV�ޘ��{�6�8�:���m&ii�)�ƽ��n)�P�W��(��鎶����zT[Q���m��c^3R�ݒ=^���żt�ᒒ�~��i�n�[8�S��,��N���o<�X�����]�e{1���^4:Ӄ���8}>KpȗK"�^.�ٺ��[>t���L�"۰��s0lP��u3��>�=���*�r��!��O�\�s/�I�YRm�WsG��ۦf
r�O.h\*p�=˽Z�<)z١8ȣ:���pdm$z����V&��9�*D�����xQ�3���i�u��t��a{C��z�ǌ�VZ����ԥҡ�>���L��1P��ӱs�4þ���o�$gnS�^��Q�M�i�v�Zjiq�#��.]�ϫ��f8{<l4y�&�c�m]�k>�p
3��2��WH)��e���&�҈���0�A.��A�N�^�#3���v�g^3�m{�L.�v�x]����V0p6��Um���M���x�^ą#�K�y�hnA|i�K���-��a����pn�|�Ҩ�Kٹ�xjB Z�p*���&�&.��=�t賆��0�;��}�r1��p3��{��l�rI.n��c�m[�kܜŊb�]���f�wH�D�f5^�I�g�������_��נ�
���=��Z���8qg/OT�,�ʘ�L���4)I����޹)���v�[�#"���cZ7>�t:���\xF��yp����(K\}2��n7�-nuz�C�w�ޝ�0X��I
��V\g��{�Y�3����w��V^EV�<��Џ�Wk�����=�����U���Wy]'�o.�B����s�FwK	B{[}�٢n����g_a�����9Y`��i�Q�>�f�6#�;�3մ��Yi��zg��k��]�y��Q���³k�BG,rY�
�ِy3�L'N��:p�.���`=kC�ZPz�Hլ�ZW{������q�ޗ;�ؠ>�����{1��k`�zիt��Y���Gnc�*��;��6�u��ڗ�����-��;u�$�dny�e�k��nJ�N�a���/=z���כ�#�Ό%a�#���<��\3�Y`疗��ļ3�;���NU����X>��ۤ=0wTRX���i�eЦ�9xw���\�l����]�m`�g>�t���g�b��N��k��:]V�R_Yڭf��ޚ�CV�`¸�r#�m0w�o!�ì�5�1JU�����w�����֪��F4WCV���,���,_@w�^ݢn�����Z��UYQA2�R�=VyA$��qpT����n��hd��B9W^ω�&z�[X�0m.��<*�Uw���=I3u�7k�y�W�	)'�ƚ�3��q�=��\��ett/��J�dlv��gg��hĎռ[��u��sZ����i�6�t�ʱ5�`�� t4�y����N*�Me�j��V��#DW_EY(�c�B�9`
�M���딏 n��^;IBC��F�f�&jB��ߤهPN��X�H^R�;p^���#(�􉸥���ˉ�nܠ��Y^߁筭��:ѹ��ov��pZ�DѦ�V�����"�j`���eR��i˫��k��s:�y��G[��v@:�	�{zf�%폘ܢ�0�csL��+����pUG!�oK
�2!֣ю���^*��#;:jޡ��u��=R���K����%�Z]�)�g�֘�/t��-���P�]a�1K? �WMo����h�5x7�W.��˗=�ׄ	�.��z��y�O�3��8�X�њEQx�u5�`(����q���X��xފ��Ώ�8�J��C&��X�T	*�(��xV��4������]����/5%,.�:����p׉����r����?W�xj|��q<�5�p�av+zd������{yJ_f�+-+˽�S�a����.��UÔdOF�e���S\���{)�:���L�e�����Ll��NJV8��ފ3�)��6�8��_�4Q2�7���2��-�`�C����Ӧm�[~�1�.��/Y9ۃ�u1v+��uc���wΥ� ���J�R�����bאl�]J�R�d:�_`i���L�dѧp������at�.����d=��ETo�_S��z_3�K�v�����F���k����-t;i�i�em|�Tt)�t�j�e��[����٨��Cr�Ю�Pܪ��LV��Nך7m��Wa������˛+��_f�\4V��}���E;�Q�ä5�3��pÖ��5f� ���8����R��"Z����ڊJ��uK���P��\*Q��;��oC��@jG���qR(o���L�u����:�= /�у���9�y��^R��>Z���!���b���);�ת��ͅy�B{tEvjЫe��v�����{�aq�%��)�{��V��М�K�2��4C��n�8��5
u'
 :��k��뛅��s�Æ��q�ђ�sV�}��+�F��}��G
� 轃������䶽�[�5��٣��o&��]B+K2�v��*�m��w�e�QN��33X�@�VE!RѥiZ�e�AH�*�*E�h2��$��Z�++��+)lRT��
�U���@���[@�-��,��صF()XPHV6�j(��+R(T
�«�,U��eEX
$��R
T�
VE���k���%J-�)iR�V
E���*-jQB�B�T+
�AT(��R�P�(6����QIiAjH�*�V�kD������eFҪ�bʁm����Ub�F�)X)%VTF�U���mQ-[@��VJ�m%h�[j�
TJҥ-�(�ŁDFB�Z؍J��la[j���+ZKkm�J�m
E�dkAaV�e���(�T,QF5mQP�T��D(�J�EX#XQj�k�����o��{�5ǰ27Oype����c��Ss�4��O8Z���nEl*��T�8s��������W^���\}q��e�b�=��ڶE��W�R8�3ʴ��`�Z%�s�p�Z��X���7 �&m���<:���s����ۏGE<mi�f
��2�"��(u�����X��lם��
��Nv�l����f \�r���!��1�8+q��h��;�D�|�j�O+�2�}������;�+�M^�F+ϲb���E�46���y"���J!��<�ƗUs����,.���)�~@��=BE�	�y��z��b�Aڄ�U�ȇ�.\��;'�ݩ+�h`�e|upyB��2�S2<u<�;p5��|}�e뒱�۾��3��"�
ں� AY���\�e
g�w�%It�5=���J��Ҝ�P�oi;bhx�?s�_uyi�r�E�C�K,$���������sC����G����J|��go;�x��g!�Ev�{�Y�J�̻0�) Y����ˬ��խ�c������j5��X�m�W���`�JĕV$�`䔚�Z:nf�����T˺6���8�G�P��(�U��n�^�G���K5:����t�a6�z���÷m9{�Xo;Q�{R�vs�ck�u���I>s�-9�=��벦�"���eN��6Mݍ�Z�+5�����o�n+����&�[�6]���jH�j���l-�{�e�QI�|�eMfOh~��`Ia�"����Ҏ�r��N�JD+���=ݾ>	��z��Z+��˔���C�v��"Όgz ]�� It�R�yY�y���w2�b1����zmx��	�`���R���rޏx*ji�R�]��;�m�w�l�ȃ���,��R]�h�6�����;ݔt��/W��,j���"���qؠ��KԸ����������ܮ��H染y�V[��bz°��	��c>�xa.z�Çڡ�WZ��΃!B��IGTYP��)��OJ~O��_�`�n
�pn�aq�
��$�xB�X7��������z��خ$�u�Y�������]�t5�6�v*��N[R�.��J�=]�	�y.�:��*�e˲�S�9��Byg�isӼ�xJ�z�a��V�C6��:�={�+%�qQh�&��DWI�e�N\�৮�l�i�ya���U##/{jn<�����9>P�N�:�?q�
[Ϊ=g�.^����3�i�u��Q��!+�P[eP"N�Ԓ�%$�:=(-��W ��\��;_Mx7|�͵��"Z/F�_x!��;�����*�ڪ�����4���^�J���efҰ�+w�8ɪê댭�

��H.�sn�h|��]� [qLx�C]0��Q��rz�YP�g��K�$`�.y_�[9�,�lL4Ms�I��__�Pq^q�����3��(�{��l�X�ly�*�P~�����L]�ɐ�:&G�M/
�GR9����P76.�߯G�����.Wz,����x��Q���',�xT7��I����>}cxM��'y�D_Rł���!��)���X{�$���bU0w�(��o�( �>=�'�]���)�Շe?yh�U����ۮqp��}�� �y�r�qXY�Ǟu��a��D\��}l�$�(�Xܫ �Z���R����X�m�kە���u(�c0ۮ��N��n1���#��^/RΖH�Z���u�xdK����-�������ݐ?��}g�Ղ �����^���޹�۹�^�����5�����7�}z�n�8���z�C`�����+��j���9�7�T-+�wr�}|yt��x˽K���Cly*�v�iï�+�
��ɡ|)�py�Iͺfg�����~LDOW�ɳ_e?-�3��ɢ�V�h����4�Cf�[�rw5ӲtGq�C`�7�|^2��V���:Vht���J%yA��X�}a=��<�ɸ۹���7�x���׬��O��Ao'A)�����'Ǎ;pQ���,X�uN�ڃ�� ܼd�wy�<�ԓ=WJ� ߰-���U�@j�S��"Y�p��X���p�1����<5�c��j_}�`���ZhCdu&�=wㅖ����o��Fs�z�|��m]�S���s�g�{OW�'�}2��T���$��9��CV��R^u�L��}������̑�0؞��	����y2��r��(�����{��f��Mx����F��a�?�_f��	���i��/��yp߭xTr��l3�\�Ѡ���#�&vX��4o�b���NZ��|�ؤ�y�����;�u�K�Ӏ4��W�(�*b�v�x��n��:�?N���xo��[H�PWT.���	v3��LƲ^\/�]��	KA�xض��M���vLǄP#g�����/S�2��w{�i�]�tR�5�����=z��/�q�>^���6��X����Bl�"d�<8Wy_ԟ-�����g��t��1j䟒�G�W.Fx���U܆��#�
�o�Gvў��tϘ4�u��Z��l�y��c*��y�7�����3>F��l�	��$6��5�Ӗ��]�]n�şq�!�Ӯ�����h���2O>�ugT�SZ��K(ΐc�Mqm4��/�;�O�s�G�~'U�^H�+�G�lC-*٤����h�ӝ���oqңsO��uw����S6uz��̀���.�O����,�X}/X�6�]�ў�NY�w�N-�v�eCc=�����PG\E�pX��m'6�.K�-:osn$UV�r7���@��m!�봼�X�q�:��%Uǃ�"�<��;#s��(Mr�P��Ef��is=q���'��V}�R���v�T܊�Y`��q&7-���>���{#ݚz������g��G�V��n��G�ޚ���@�9u��9�2֢��WT���^ɜ�:p�hx�����|��b_���q��#C��^'�R*�S�(��~Ő.�xV�[���EΜ��R��Gɩ��`��'/��({��<U����h�\dBHo�ٞ�~��x�J�זn�!�R����M^�e��\�!�W�(qY����k����>[��[���\��V�j@��we��U�Ⱥ������W��y��/�k9�����������]�hbԘ7��e��)�c)�1�#�S�þs4�j5��t��h����L+���a50����Ŕ��7�d�5׬$;�,Wn��q��ڛp�ta��z��:��Ƙ�#�N��^2l�7}}|���E7c�����i7ݱ�c��7�T����K�Wt���E>��u؆P�F��g�+/�i�Q��.O��������m筛�>���@�/�f�V)s]��3�޸�8=%�CIcYGu|R���_*��Uظ�ȯ��P�]��!t������.���ƤY�w�s�e�ՠ�zO[���� s�#rVD�Wo��Q��J�2���|Y��3����ψ��+�`���{x_�,凵Ҋ�t���%B�&c$�����L���/)�h��%u��琾{N�Wx���G �[9�������W�
���+ԽҎ����Ҿɻȭ��sz����0OR�|��C~R�{c�r߬�ى�t`��@�~ R�#������}A�?'�����e�Oe,Z�����F+j�㶤[�V`c���k2;�X��G���bTt��b����ݒᨡ�vi�;9�����W��`��)��2��ƒw��]{j��Z\�s�Փ]�7�/O��`���&:|�3��%���@�zq.��K�:
�Y�2WNfC��ޯ�_�L���xo���7�*���"��ro-��,wBA1+)�_d6
���{���o�gZ�}:d�;۪�JR��*�y�X��r�i�����C�i��Z��C����Uyz�?o�~���v����T����i���#�0�`�i�2�����$�oI�w'�X����nh�Y��d\�o�d��Ke?���`E9	�-�{O�հe�
��Kp,���#��b�����3LZ���+GG��E��$g��FA=;�瀔9�6y�>�Vy���͎.;��A��L�[��nx��\]'I�)˚�ʄgl�z�S�G��=~�@�s�F�y���N�x�jZG|��!��sQ9�u&Xv��H���mM��̯.���ͧu�$��a�Is�����,�lL4Mt���ƾjp������J�ų\�Uގ����s�	W�������*b�p�邡������Oq��}x�m�����S�"�O�ӽ�o��v��\Y��y0?�ƜQ���9L
4=��~Vڋ;q�'31� �"�G��>&;k�Ot���\P��˶|���C0�BP��ٯ�_����tn�V[$�mCk�E��u�8�����f��w��R>1�pl�y�ʲ�5	-�s�*���� �p���ͤ���E<��-��(^1�7[�9��5X�%c��7.�L��7�D{����&���{wO\ȋ���vk�CAlέ
�z�/%�h	�}�6�Ǐ}��N�Ү^a�P���ح}|e�c���� �m��ͧ����8�?U��ue+-�EVZ{g]�YPy�����#�/�`,�__�xJ��u�%xa<'����Av[��x�5}�Mú_N����﫰��۞�����I��g�~�x�i����h�%��2��3ܼ�:��o#�!p	�uq�����qmPq'.Ǥ�ZW=��t�Ń�S�:��yۯ���ͳ�z����������%U�����fe:�����/DOU��-=�L�N��)���z
��+ �"�X��O>�|V&��8<�D���s�N�kC�k�o���hv����x�2䠘�*��\��4��~��w�x�iy��x�S�Um�27���F��Á=���b�R�=��6���K�wwS����A_o�NN9OS#�Q}��p��@P�߮�w����G��E�r-t��o=��Z��@�O/C5#)�ck�:֞��P���t�oּ*9T�+a���4#gӅ��n۩���X��\s�
	�WƄ�����;�u�	yzq�r��*br�HE;]��\��Rn��eB��j]�n7<���>~�{@�/�����$�w4� |8�jZ�w��c{+:�k+��V�+��<kj��Bb�)e�w��\[
�7���� �㔫���m��{��;ۗq�G��A�Xs��A� �4 J������KlV�e\s7;��Hį�N�w�]�ݴ	{�u��`i��	yp�Ev�:�\��1w���)>����L&S"�!(s���W%�)�y�u�'��KQ��wYҦ��$9fz�߱�b��s�Um�>G>�!ەB�� U紶��ӎ7�wײ�I�$:�3JŚ\����Yӻ(|�t�VX6$4�,�d����g���2�I��Eܺ���ks�Ar{��Ma�g�=���g���%�\��>[�	�{�p�"�����i�+׽��zG���s�o�gZ`�9/Jd����a�^��,k�ǰ=��ɵ�r^i�z�[�x#ѧ�{��+�K��E�N��%*�>�[7�M�}u�DX�2J�=���(u��n��c��V�Hs�[\��mG�ՃV�q`��]�G�]ȯ8U���n[3i(����^[7׻\��r��8j!Q3���u�ExZ��h�-\(0B�K����yuw�N঍��s���t��
w9C��N�;WZZ�GKZj�Um���q��نR���~Wɉ���.s����_�A�s��c}���d�Iԫ7�Ȍ�̔���u�T<*pʹ�4��o��s��+nw5���ǐbq�Jѝu�*�ꛩ�r��n*q��%B���7~���[>��o���
o�`��_x��H�zN6�U�i:-E��L6\ꄹ\�c`��τ�g��P-����l��V��{���j}UL�H��]m����M^�F+ϲb�0�Y�`�ȹf����U�,x�6R�������W����i�x����Бi��xr}=|ױJ�;m��J��䱹���x5�$�6�CTI�y2��B���җ��s����\�7�ϕY�鰌O�����Bx߃��Xp�� ���Q+����X�\J��]40e� ]��}1g��`Ǐ����<z-i�dW��ˇe�,�6I].*�8����Z�@��k�~��~�n����m.W#��+"�]�^�� �!�uF�#��؈�w�3��Ὡ�9������Ǿ�.��G�n���>�R(Bߤ�`��Rk�Ih�2���\YyW)��+���f���o"E���`�nx��u�}�-%zయ�,0lIX֥'x�F�n�F�<m����M`C�]�)��+>�,�z�&{�׍|��5�%O�����	W}�a���<y;�q>���:z���uüA�NbR���(�)iD��;��)@�Ė�^gw�0q�3�Ǽϵ�$ڟ��
�C���PBĲ�a�6�	*Ȥ��J^�i�I�Xa��1�5��ۍR�7�|h��9�B@a�3zL�5d�ȫ����wG�V!&X{������T,��0 7i)��f��Y���pT�M^�m�5` ��j<Ɖ�d��3|νb���A��IǑ��V�nJc��Igp�VŘ��(����-�Z*ctYM����Ea��Ư�ΐ;�2�ٌ1���EIk�q��f�b�^T,���]ǘ���ڜ*�\�����+��Ӥ�u�a,	GA����Ѽ/ �5)��~ݮ]�g �gv��o*���˹z�AB�)L��˄�xH�ȗqa�{�t�)�<s8����Q��ї�j�%\���Չf��ݠ�&�F�j�a!�۸�f���9���ثbz�Q)�e�:<%R��|�=�����(�����A�i�{�x�4c��;-�W���N���7���/�wXj�^�o��7��i6�U�âls���W{W5��K����2�'�W�)�Ю��{7fmH�^̾lF�����#r��7�b�7i�T�`��[�dЇM�(�\�Mj����ysSk�
7����ek�-ʺ(R!��q���f��a]�~v��%h�Ys�^�
b,�H���T{y�V+��'md��Xo�#x�O gSV��SVK�"%��j�6ժ魣v�̽��~�/�b�c�b2�,0\[�)���}�����y��BPlO۾��y�D�t�����s��fgQ����*�$nX������\x�J��[��k7X�X����iR�FHB���i{�C�^��!�/d#��e��#����H�>�ۏ���P=n�[��f�ݻ6��@j`�6�L䯲w���V-+�����|�p�ʲ�`����:U��5S���">'Ytc���n�zsٴ�#�ox�����ށf�[=gϲ�I���
tA ��x�f���6)TiQj��>��:�G/u\��6ݪf��U&8�̜���/id#�en���%@�1cȗ,[���z�ie]�N�̕���᱇�hR��j��{�1=��J�M
�*T8���+��v��)���::�=��;��p�,l��2:X�"i���z�eB=t�VP�|*��K#�{��բ�5�:�X�O^�ܛ�.<�C��r�<rLT��XynG��五G�	�QY�ËNY�ʌ�Cm�[��L��c�Oq;N��XN�w*�X�b�8��P}N�d�ROĳ�S���U]r�����t*�Ib���ǗN���j����gx�͢�c��q��B'�����z'�d�-��o�akmKǏ ����/����&ۡ��n��B].�i��.+Pŭ"�6�AH�Z�[ET(�AaX,U"#[+YF6�EIX�b�"�Zѕ%F���#[	RV���!im�R�0QaP-�"Z�KlF1�j
E�E#�d�AQE��V���jA"���Y"�XU�b�+Y-E���T�"�+Y""�RV��PZ���*�[b����edD���UU�*"��E�**�h�-�,DPD�¤P+X�
�Z���V5,U�*����QT��,���X���RV���J���b1T�PX����edjڑb��jE,��*��TF1DDe�D��*�hTYY�E�ŭjQ�b�UUb¡Y��aFV�,J������q��f\�
�AX�T���T1
���*Ŭ�*��Y���*>�ϼ>�Ou�lr9��=Hs�v2ҿo_'����\_Y���q���#�ਗeFL�t�Nv��8��쥮J�6�d'_�id@
�U���؟E6��'�����mK�#xm\�jE���5�+�.�3ϝwL�X�σ�m����"��oi���d�ܵm��/W����W��(y��7�T����)�0{���0S��Hq?'5�#}����Ƽo�q�--�D�??V�!��j����ZRh�W�Q�,�C�9w��ޡ��r�#Ҕݓ���m�z��z��=9UP���__
���KecF("���\���
����B�>��1�:
�qR^K��+��ϩWR���r$s`��gݤ_z�sR�wnM��|�����:D�/3����ڨ�4�$���)���Ϯ��s�r�|��=��cts�
[��,�ׄϜ��̎��
j�)uH��K��!��3�ų�ٺn{���IJ��σ{�x��)��f�*ƑbN~�	�s�=���tL2�'��H�Dq|Q���F�wS�լ���Ѵ��Cq3�O����������L]�29��P�)&Mع߸�X�!Ui�,LΑ�aa�v��J��ӫ����3z���7vy�r�ISL����B�s�xt0.�nV��k"r��=�#Y�
+����g���D�t�*�=TX*���(��E�<�;��g��}w9^>��%��*�|�W*�MIY;Y���t�mԷ�K2��V���E��`p�r���9<ݷ*�����sӰ^�&RK�#1&��I��^�t�՗�-%`��xe�
�i��h�nϯƔ����wu����y��m�x?����������wW �{�������dRҍ�]�^%E4M���&��D��yV'e,A���>�ί'��9x�qQ�{Bq�QV�\Ǽ�_�ڼ�:T�������](��_�C��}z_�W�fU3骤���ΫW���=��ݎ�e+C����Pz�����қ�gw�<l6��G{�}��l�/����i�� �XZS%3x�2�\D�aĜ��W�o�@���p[r�G�z8L��>�{]��Q,�=IX�b倹�|*Dpy�Iͺfe9x'�rޮ"s�M���U��r���>p�U�B�ԱM#�QJ�e0h_
q#�b�K=.��{J��v<�N���������si�kY�ʇ���<��g�I��T6e��ZJ���.�I�.Vq���e��U?6��=tZ/|l����i�I�6���gX�%b�G-�s�)���|(�(r;&C�781g0�����F�u�Jb���F�H����7Z���[.?N����O72Pڂ��;Tj�TG����`�v�vSU;%�"�ޥ�M��sú3Nf�E��a/k�y�9A2���'J���>	�zS���Z�E��ӱf�TG=`z��}~j���g�س�+{�� �^}2��(�y���3��F���)�7z�AB��"���W�N���A��.{�{����{����e�����09#1N�A�`����q�eȫ�A�\zmw�wp�^���N,��1
)��xR���3�cy���~�j����@�:E�����wv�%�δv,i�ԫ�_
G+'��6�5ٙ��?j��߾�S��f�*L#�I�rV)�uP���܃>�I�G����C�x����Ə���=�*���!���҄;`J�!���{edCpts=�QG=D�Q��J%oNK�-s����Y�7�@{�3�7�m��CORΖNڳE�� ��=Zz����'l5m�K�՟Z�+M����5�u��(jPpXV̀�L���	w���^�R!UͻYf�]��ǠI��ӷ��i�����L�_�[�Z��gz����SW�Ԛ!j3��<�!�s�,a����:�м~rV''��S��-�W�ٵ鬳��7e�����g��Ӷr�I�dҔYryU���ek~Z�G��t�]�3���:ӱ�ώpp�i�V�x0�:)YZYPI#�p@�b�;.X�m�8�4����&�4�u��u�H뚲_�ǂ��՘�r��k�C���x�jǻ�u�I��Z �����r����wڦJ�Y��Z�0�/�R:)��
�����m&:�U!�8	��5�xݞ�=�{���3~7>��þ�;Pɮ���VR8Xzj�Gi �V�;up>���m��G��.�W�$�,�˧s�>���X�_���֎-�~8���}���S7��޶-S~=�ew!DJ�-NM+�ΌQ`��a�\ꄹ\�{t�g�
�\r#��#�*'nW� =1��F WjIB�]Q��+Ag"����1X�}������GAX��ח�z	�OUA�����^V�,Y\\YA3,we�;�bynmo�E�{��ʐ ���ݺ�y��:��'�4%�%}.�5�����e�L�M)��4�ugj��M΁{(5��/��"�Xx��3�̧k�8t�B�D��5�B���D����p.'��.�=�6�$�"����L\D�����%�D�g#��{�[.�~� �=S��;�K|LT�*g��͌yX�}F�͓Ü���ٌnX��>�ʺ67Z(��k�ic������ٟ\d��V̛��͚wٲ�&�9�GY�3]����k�S�;A��Ǯ;�0-��LM�1uy�։b��V��J�zx�R离�e&�#��%dA�T�w���>�!�.�8�i���[�7x�O5��|��f�p�i���Z�co����;���%Bɘ��)5�$�t�"�n�i={]1��s��`����,�l�J��=x_�֡χt���(-���+�:����Vsb7=�N��'��]VF�'Z6}5xi��R�c��r߬�ͽs���X=�2�WzX���w4��W��_C�O�t[�shI����z��f
�8�+j�㶤@QK��6q�vE���٥qv�n+��ǈ�ݱ��Zw�{���t՗�^�0T�����Z&�f�yj�� �.����A�rىԵ��z�k�F�o�ڳ^W�Ա�ѐn�7��`��M����bz_��Ŀ�R���U��P��x}NfC�[��cP��L�ݾ[���
�([����=��D=��,�����eUqy��&�¡&�u�X<��qH+Ư���X�Tf������+�O}3�j�8���Xҡ�Q6N�-LqGe9vZu"G�!1I���T���-�9�U�H�u�*�\3~��^�M�%��*��s�>����j�{4���D��+���L���,��v:�l0t�UM���W�[Pi��[�pg'V-��3ƫx��ڝ�¤�ˆj�t��1�ū�L��c��;��R(�t�o"�DL �=q�ͼ���ޢ�ʘhu�Di��&	;�U��Ӵ�r��myz_+cQ��*)8�oM������^������<.Չ������0h�|h���n����!�E�}��v�&����W�ۇ^�V4�s�����s�_�τ��0@�Ȁ8s�3��8�.��L#�B�!�1q�'�;�5��W���T/V �L]�ɐ�ɂ��i�<y.��{�'{�}��Wj6KKH�Vgk}q~�5��=�`p�R��{/C��E�l��ya��x�����vRJ�JE�`�\E$� vע��������A��׉�TY{�,�{�v���(��o�t���u��C��.֓R��q#/m��2�9?l�v���|�o�&�:h���k�h��CL�c��j��zאy·���f�i�>*Q�/-���#��&V�+q?:���Pw��8"�z�t�)[�^l[��I^��ѣ��qwh�M�{g���3�v���Lx^�ذE��S}L�t����V=:�v�l��WR�ʵ&�^�7�����m����ZÙkK�-����R����#�ą�9���_�G��,pΚ,����Bq|�5�0g����U�`�.�Y=iN�2�q�o_Q��r�:����[J�^(���I#�$�z��ޭ�<ލ�9��ft�����ݙ��q`۰��Nf��ZV'���G�v�y��})�}H-pWJ� �]���债�����E���c]|'WKw����]F��ppކ�u@:'�祍���+#�����E+����|)Ď1R%��,�Uֻj�2v�}�a�O�\gAZ�2��t�-4�:��J�̻����|:�T�k��*WϹ�v��RAZf��،�=cL8��r��*5�L�z��<mi���1=N�`����0��e���S�۱2�Ȗ�,�zY0��x,��[ޯ	2�e��ĳD�YP�.X�*a��s���+W�@!Ǐ$'���x'Z�ՠ����1w�Y룧|jc}1��)�^k�ǾV��{L] h{iD�f4�dp�4�=6�P�.��^���9'W��=gEѯ�ܪ;^�2��6��g�)�ϻ}���K\�9��5�:��Fx���wo����Y�bx�W�ys��w �� �P�a	疒��%
��7��ޚ�ܞu<Q��>�����,�gm�׃@��[���mg'z)�1�ʙ�W�T��k���P��L��ya*X�f� J��FR��*�W�\J���!��\9dÜOLؿ�e�n�W�n��d�)���׹<;LL\ٚ�ewSAXb��^�Z��nP��؍ߡ��++dJzQ�|�s�/�0�U�NHi�8%v$D>xB�:�[e��q��a��a�k}����5y��5�q����5G�VX�� �ݨ=f廿
��b9�M\�)3ݾ~|[����y�7_�Ħ.��,rX5�a[ِ �&ut�|o��~��z�X׾��n��+k��#X��|W��qpr�Oem���.��E=pX��m-B��c9�V0�̗�Z�>��x�g�k�C���R�c������%ǃ�"�<���|�Y�}Q�kZ�@�oS�N�]���O��c����Z�Ŕ�����_E���W���y%�җ���P��`�3�;P�5�}[��ܬ�p�f�,��-^+	��7[Ò�m*�k�)X ��m�9�*��̺w9C<s�N����j�'J�a�d��Y����[ٱ�յh�Ȕ�	�D�ъ.�L!Ψy9|���Cݓ1�?U�3H���={ٝ{K�_��^D-��I�k��YȦ�}��V'�d��a�|���S݂Z����r�Q�s���dac��g��]gk�ƖEf����\:��hb�%A�xsi�V�,�z4���i�B��'eP^��;f�6�m���>^/�FU斬�h�};Uu&��i���a�p:y��,���-0f�xAV�[K�_5w+�E=���j�u���xzm��i�,Y\\YA3,c�-:ߓ�sk~0����^�I�s�J�����]g�I�q{�Aڄ�=��@֮J`.�^}B���SC��4�߬�y�ہ^;ݞ3϶�����Eç�#��~z�,���A��J�s]��3Գ'�1BӺT�������).0	:顟t�5�Vg�y����ȯ�˗��d�f�!���Ӳh�n�W���ͫ�vV&���Mf}���+"�]�^�CVxg҄;s.�:��>��\���|�h�=�RT��kHpaB�ߟZ�3�`IXT!\����]�y�E-�t���'��=UѾ->�j�ц�t�o3ׅ�Jt���1�<��X��0ڻJ��шQ��7���E�ip�L=���Ɲ�c��eo��u&o�Ul���e�Ә|�X�S*^yHn����g�۱XO�@j��\�0��&YU���OQ<�>�줠οCZj��WU�����,{���N-�g�~�/�e$�%�QCN�7y��O���*�F���':���۝%ُ+���Z/��ӕ�崣��wS��=�aN�8������Oj�f>��[�f��y�Fuz��H+'-�G��[<�-�v�~o.�O���1�n��>��o�T �p�\��9�1EX�/-��dS�' �-Z�����A�0��v�v(=u�AN�-> ����z�O���W���ӘO�
��:%;y�#��Ϳ �@;@yЮ�:5*��c%��}L�r���^1�u�B�w`m<���1��#��Y��V�-5�W��@_
���Kep�3��^�ѫe�W�~���?}?�mt�(�'��Z���ҩ���s����+�SF�a�ӎ$�>��f��Pt�@5����b�,�hqDiĹ'A�9��H�>k��G.:	eS�+��P�܂����g��#�e��b�C��-#��;���0h%�JQ�V.���y)s=��Q
�f!qi�V�bN~�OK�Y��̙d�ba�Mg�?T�&eM�d�x���y~�xB��Bb�S������z�9Sg�d8]���:�������V1�;��H�:Q+��u+3�����,ŧ��U������Â����x�:�V��b}%���C-$��"��\E$����K-aϻ����g��u���s�@,b�	7O�Ξ�7��9j�+}�e��O5�<hQ��1l}����p��ڿ����7z[�#6�O�F��x��+Z[�6�*�.�����K(��u:�xu7T�v�=�8nm�׽���{j�wr��沎_N��ݳ��7mBy	q
`���"�c�\����t�C{��R#�٘���V�ϡdc�/�&�i��#��}��uc{�͋�F��c^�K��A8��Q���Qە-��Ly����(c GY�Z�l�*Cw�I�u|�*�����N)Ic{(o)q 3`�vs�Q�f`�z��<���O�	b�]y떄�2�an�l��lIV�=p�.<���sQ#��::4�(ȜkO�V/n��G�R�37��q�(�.�nom|WW2�������VC��QXe�o�71If��*s5ܓ�QX��{�j]+���-�K�G4��ܺW�q��x8QɎE�π9u�l�����O@|#�!��헠!��'/P�ɜ�Q�	����u�����R���P�%w9U��t���&b�QFi�Y�Z�mq��<k������4�J�ɮI�U:y�y�6�n4�m�.���
b3��W�{w6�P�Cvx.TB׽�we��s�|<:�[��e�� 
vە��`��Q	�����)��.qe&�v��R���-�ܝ��oܼ�E�*��(^�}�Z�RF^u(���ZI7,5g�s9�������^�t�9��WZ�^޻��R���'��r�p����ܢ(oE&�]մ��)�d�]�����؍����V��C�Ы���7�]��B���S�;�MXZ��v�k;�k��c:EO�`\�M�m�{����$%<�@`7wB9}����s��>7*nj�@��K�=�Ә��0���Y��ƥm�_֤0�k�@�z��S��)�e�Jeެ�AKzoM�K�nv�F8]ݮN�-�R	��|��h�����d����nt��pT��g>�"H{0���	��{|�JC�8�5j�c��a�Gb�XRM6�%sp±
��S��ِv��dS)��nT�`}4��mSm"����HF����:�mk��_q{���6%D|�>����PoGFK������DG�sm�}ŷe���
y[���G�<G`���:]N�X��{j�+.s*�ԩ��4t�,^�BduMUa�]O=�r\�1˿f��@���*��ɝ���q����:����jn���轧+u�\�T�ՉE��9@�W\�֬�"^f.�ɥ&K�:��a�/^p%�,����7���A|Y�S�fVR8$�A#�]����p2�n��j�
���E��h���/U�x	.�!S+	Ō���?y��{"�nȌ����W�j�~�j�T@j����s�K�3,Ԋ��1�,��~��f}�3!m,����H�
��B�*�I2�k
�Z��YDU-*bB�*6�l+s.@Z�H�m%�EP�V*�FE�*���2ER*�TT`�Ak
!mR+��hcQAK�cb�
���b� �ciDX-K�V��Z.0�VTFЪ�al�Q����EFEPm*KKX�	Qb�ܴA@Ơ��,�-J�PE���""�TQb�V,ė(�(�aj�LB�*c*��YHb�ʂ�EPƈZR���U���QJ�P�E��,���-K�UAEV�k�1��d2�EPĬ���n0��*��F"Dq�11�ZE��j�bUH�����LC�E��Ȣ�T�LJ$QV�DE1��,P�̣xF0v	_b�7��jg�-�<x�������J���ȓ��la�+ߖ�˂��/�����o�%����~T�f<;̰�,/��GD���l���lD��}e�-�M�����zR�T;(Sa����7��-`k�J��1�d)�w�O��bf�6k�m,��Oίפ��@<�=��c��X��P���n(�:Wk�
6ǈ�^/R�:Y"�~�����q�EIO��y�N���gZk6
ҷk�3���^�ذE��[K&�ݠT<x�Ӡq�.o6{{�'V��~���?fFU3�dP�>̀�r��6�8����*�rW(�}��eE#��ͭ/�}����aU�-z%c���������%���#�����=�Cau�[��iR�=��A��{&��ּ�8�j���;(����������W�q�w��Ckjn!w]Bs��p��K��)�yL����!kM~䟩P�B��,3��zX�3=ѯU�f��^a3=ӱs�4É��/kɔ�_��6���)b���������&���*�����؋���j���}�	��ೃ�fں��p����5��	�Ҝ��Dۯ|�6��v)D ���ŸU���:4�h*�J��.J�1\úS5G�tkoY�)�;���u{Y�r�X�n��.��D�Z�B���h
�],]��ѓ$�꽭��L�q���
�!Ī���v�	
�U7���7k�yx���徶����R��&����ś!�Z�A���x'Z�տ�B��<�)�v��%�7<�����P�$D�\*��`��/�k�M���C�^��k�wA��Ϳ,�c/�⡘��!�����JUϣ4o"8��xs��k�t:��"���=O�8�͗�o9����3��-p92���-%J�8-%���7�����33=[s��n�U�CŴ��n��"��[D䆟#�P�lJ�!��З»�z��	ű�g:�Ud�/��j�u���S�23t���ƨ�VX7!��t�}�z�˩9_a�����s
tÇ]�b��n�T9׿�W���E��PU�
�̀��y3��t��܃�{���T�q�;�i˾�3�a�:��gʡ���g=�p�;�ؠ>�c\<��n��q���MO�8}!�	hX�k�~�X�t�����c������٤u߼.�ȯp?/m 5�c��7���u6Ps\��FJ�Y=�Z�V�pe�r��wzvƦ"�a�گ�.�o���	>'$�/�z*�.�'ˎG�c�z��3��؃:���#Ox����˙u���FǛ�ID qp�1փ�g���I=�Ld�w*:��r7����Ú�\3ظ{=z!R���K��DP�ǧ���I�y�����ZSrٙ�9�w�;Pɮ��ܕ଴p�f�,��sݭn�6>�N-��g����B���{�2��f'SS'�8��켾/e�Ů{.�m#Vx�G��]3e�߀dh�R�����D�ъ.�L6�P�N_4=��C�����z�޼.9�.vΏR�Xtq!���bKG�"�־�`��;B��7�ܣ��9.�9��a�r))x�'>�,B.Y����k�,�.,�����v�ϓ�sj֭���c�x`�>1����}=m�b�:P�#�@ϵrPu2�P�e����J�gժ�%���l��_����0�g�z��R�x5���&g𞷋�C�@��Q+��5ڰ�ȕTG����^��u�i��顃����Vg�2��<dW��ˇe�,�6I�3����H��8�υt�ƴ�}��T7T��n/l��ds6�dA�+��B���BJ��&��{n��y��l�όƑ���Rge�L�+�����Y��J�B�3"w\��Y�45��Xr�/p��x����/�ފ����|7��+]{���pkf�<zv�0�v��}���;��1]�0sv���d�����my�.4�n
b��ǫ\+����P
�y���R\�CҼ/��k8.�����uj%eK�X�E�ޱ��cf�V�"ǫc~��>�j�_M��r[���Vڇ;��������{/Y�CPӫ�|r��ב�c7kE{�ʥʤ�N[���G��ݝg�U��yۼ�߱:e�J�I&[Ҕ�HE6�ZЄ�U�0Mg���)�`�)�蹵_�鿿f,ň2�k^ͫ0~��`N+:^�h�z���uǳ��`�i�;{��_:wM�Vl3:)�p�p5>�E��;7-���b��q=Y5�#}����xf]S�M�ww�=�{�vƓ��%�	OR�OiWQ��E���+�3!�]-�{D�-EQ�+�*�h�̭\u̘8�ϫΏi3��RKG��=�����U�5�N�7Y����6�s�v��a
a�?-����`6�i��%"�]V^R�/.]��
w"F6�29{Xm�G0&��s��v��)?N��)�	��F�K�`�[ϩWT}�����C��m�>����Xg�:�QyP��Y4�׼�����P�R�;�v�x���R�QWG^�̈́o�uJ�]�|�He*g<��=�;4X0�}�>-�B[��]d	�I��q`��,]����>�=��z�ӊ�ϯ-U�}�,p��KW��/`��;�|����=L��=��3y�N8}
Wn�>������,A���l���y&�빴��=��-C���^Snz%X�$癆d��'�-��2Ɇ�Y�1ޱ��ҷ;��U�Q3�ґ&�_ZY��+�ꎥ�8���H�^���6��oM�H�;�*}�w?=�������9�iX�du+3��l<�Z��Zx��^L坽=~�f�Q������Q���9d�ne$�����R����*�����q��ݾ}���/��{إ�Iէg�]�p(��l}%/'uU^ Ku}�U.֯z���c%�L��B��M�<k����_'��R+�����3&���$��(�;T'e,A�^�>rt�.Z��}-�S��\��ہ�r3�c�ܭ���x�������^<��˺t�mz��> L��5�/������	g�o�J)�]j��GR�v6,��a춖M�g�/q�2��w����Cz��8{�_]���[�O��ԯ�>����qf݇}Nf����ѹ���ik���xWM�[ck#z6͊��͖��g*�,rmx�1߮�͌e<�o�I6�߽9�pJ��>ڰ�6S8|��Qّl���鳧%7]*�Wܪ7�k�{��e�H�N����i-1m��l�㕶�_v�u�j�A@��Bʎ�Y�
�[�:��X�����(�+LU��tD�y�VQλ�k�弭�|���{��Wi�\��.[�qw��&��ּ��"��^�0}R��)��O>&��+Μ��Č�H+�X=.i��<�����^��3�����Mk^�ς����>="���w ��a�\ZV<�C7ӱ=CL%��W�)�}2���]�����d��o��;��g�q��m_���.v��3}��&{�2��T�q��� �1���_�k��1�<]L�R��+�6�]�"���&�T!�&��|�rsق�ч�(m6�tۼS��,���?J�2��ú@�:Q+�f4�dx_��XT>�=�#v/L�����_.�"�Y��%LB�\��XA��@�:E����U7᮷���4��VGb��V<d�>��Z��.���(K\����BXyi!Z�rW�:�,��߈��(f}b��8d���%��϶RyX7zёY��Um�|�(C�*��� ��&s����ѵ)/`�=w{��S�>��vp�������tMI�@.�p��Y`��z�t�v��uYB����Ⱥ�
��b≸ޒk���e#]�}��U����E���\�:�f5 ��r�@�ٲ�#��`����ST�37�o�Z4>�8-�=�=�H��T���I�ngb���hn!f��!�����<6���R�y�l�Z�ٗ�z�`���؇�4|%�g�T��z-�O��,rZ࠸=���k����nse�Oy/��	�csm����|�j��tg�2��}��˺7;+Ϸ��>�k�iuty�g�g��~80<��%e�F�|~�ӥ��g��æ�7�c0�:�x���>����g|�/L���h��\���ȷO��g0�/�R:)�eәl;�Y㪷[疯����<-2%�L��a��=C&���@�P�
�G�j�={��<q���[��×�+�k���G[�-=�̰)��	r�Y��o7̞Mx��� ݠ:��}o��y1q���mr(q��D�yъ,��a�\� N_4��݇�N�un�u�ᣜ��x�a�6�h��E����TG]u�V�E5lF$˶������NfG�ԵWn(aqf�Xd_���v�X]H�eqqe̼ww0�TB����ܕ�!(�y�qv{ީ�gM<��yQ����;W"W��Z�(��^
��'o�������N����t�`-����8^�KeZ��ӫ�4�4��PF�ǻׄ�1��b��B�u�7�T��.jI1�<����q�-�S6ҕά��;̯���SlK��,;�r:w�@���2����j�T%���t)>Q��k�=ǂ���v� =��t�W�}�[�8�a�r]鹕օ�9�@��D�����ڃ��ݻ��N���(V��޸�8=%�C>%�q]���5S"�G�\;�,�~�]����o<s��/;�#�+*
Q���9oo�{픚���� �+���Hj�
x</�ёn��Ň=:*c��4\����<�L�+����Qf�%bJ�/��]y|���o��~Uk�)E��G�]TU֍�J�@�pbo��}.�X��Z�]��:K\�Q�� 1m�OT����p��!��F�'Z6}>��yT�n_g�y��h�+�����^���;Ə���c\�W�BH��S+�vu#����`L�ٴ	��e:������N�fj�V;jE���]x��8����<G&��Ӽ;݃O����)C!��O����d��]�O����
_>l���l��Z���z���,݃�&e��J1�*�g��8ʣ��m<P�W�P�0|3��S!�b�̄�Sm�!f����<��D�1�G�g�u^�d�0҅7:��w�j�8P�H�NQ��(���ͺ5������t�SZ��H�<N7�ò�+sw'��j�ķ�=�U}L#l�b��@V�v���t�?�1��@c��ӏ��
�֖u�n^[緪�Ύ�����d��f���I��M$��.Y5�	63��ʲ�;�^�/��ZiMZЙ�rޮ�({�6�i��R,�����\^�eݹҶyb����y�Ui�y"�=�pJ�y���a�֨�4�7�[k�Q@A����t|s�~�������P��l�^z��~�<s�j�R;aݠA�{{���<$Ύ������3�/`(7c/�B����6���Ni^^� UoY�H+��׵g|��έ�'�L4O�"O�_rW�q����uOs�}*�P~*����u��.�א��W�{���y2d8p<���ғJ�S#�Y����R�}����3{&(f׃�y݌A|�C����#�kF,NS�@�I*)傥qb�����,��$+�E[^r�:sY�0���J��%S~r�D�x<�Z ��C�	eߺ���x�(�����~#+;��=R���W����	��6��&�Q>��L�^A��8��z�Z��j�`!\iF�Z:K�833�MK�k� �r��[��T�F���]L��b���Upfd�q3jg[1�'\�R K�-�u%c��rrFe�#�觳�El��;5+V�&эYA,�[��nu�[�35��FܫP�G�E�-㉽�;%b�ٴ���Lg��5�[�5��]�Q���9��eo�5�#3�.	y���M�X�p�T�LL]��ʩ��)�]k�rԾݱ�`����]^��]�~ھv�3�e�~[��
�����o�z���]�gRђ��}��\DnÊRZ;a��_$��}��}�2�}�{������ث
͖��g>\�9����Ft��~�(H�������:I���)��<��B]��M�;��^V�)��j`�|V����`ՁѺ5Ry�J���SR>�H�L��sp?�����S<dv�ƃ3��[ֱ�ӽ�c��AJ����ZZ��f��L�=cL8��r��X��}2��Z������i+�ǒ@�/o�eUݻ���Ձr�vW<i`Յ��f�;zeoz������ީތK}��Gip<�x�OD�<Wm8�]H;��y:�&������oeuؗ���@�ڣ!3�}־i�k�e�F�hJ��Q:;I���\7��w���B��d$�	'���$����$��!$ I?��B���$���$�	!I�IO�@�$��!$ I?؄��$��B��$�	%!$ I<�$�	'�!$ I?�	!I��IO�!$ I?�	!I��IOHIO�����)���� ��o�),����������0@o�x�T�QB��
����P$�u�PAH�󺊅)T��T�(R�mC�.�����X�v�K�)�.�v�]�������΋f���H��`�@:	Usm�(�;���U�2H���RB���vȡ�lmmm5)hUB�dvcZ����m�l��Ɖ@89�cCm)-�[T�)HdH�&�`��J��D�i!���l�T\��j�QV�YUT%�p      ����J� &�    )႔��014����0#&�h��j6�h4�244i�2���R�H` � 0  �0# #	��14�I���ІL� ��f��hڍ�6������������! D?�����Id@@! }rHI`C_��52	nH:�6��4����S������C�	 ����QЇ�@$�>L!�`#	�J�+B@�H}ߏ>�񽁠O��?��?����$���`g��X����L�u:O�g��?!�B�,/�{�s���sv��f~}n�us�뮹(����." +Tp#�ܭ�4b1�aq��Z�sk/F\�u&u`YIմ���hn��º�M�yٗK��f,A�{Z��=8ز�c�؛h�$����d�����ha�ˢ�L��.�,�%V�{R�/]��m��w:(�㤂��ح����fC�1CØ�UϤ�]�5<H�:�n_2HEP�]�ׇ;R�M��vĊ����Xjm���˥ji�LB�����9�H����|΄�/���z��]�^�U�eab�I��v�,dݨ"�(��wn���xɊ�El��bfݘ3mEX�
��Vw%,;3��C���}f��a�˂�D3��lb@@��fm�V�X&I��:��x��Jɂ=���7OV4�ݱ.G��0���ݧ�X�h�=�E6�1�=��#�fo5�)�ڽ2�e�
2���ܼ����I�6T+ni.c��k�܃z���;7yn�x%ea;��j�f�B�E�7��MXG*��D��k�em�混�c;*d�@ct�ب<5�%i�������X��+N�զ^��X:YB�R�{�����h'Vm�v�Խ��������o�j�`��>Z�5l���F�)��un}��R4o(��#
Ƕ�ٺ@�c&�Yw�YStĞ&�C���nƨM�3F��i�N�i�c�X�i�5�	)jy��`ٴ��֞5*[���e��[��㹡�t�
�E���Ècse��xF�Kj��N�f;�����^�A t��FL�n*�²&o&SwR�4#�,�����mȂ����%=�B��4�(V#N|��%D�.�R��)�Z���<��r�W���FɫD�u��a�Rc�E�V2^�G�[��]glca"K��h���5gM�%���іD8�o^�;u��Z+N�]@�2֬����
Ia�
h�ʼ���B�@�e��塵 n����;A�h�ƱW��g�t�ۺ��LA��d���;r�Zm��Gr���ӵ�dK������Hn���hpTX��+�����W�;�m-�٢4�����)���a��хe�6*G�9Af]�Ï
U���%����֨�,����7z��p���˛IYe�ѹ���5�vj�a&5mm�C���Q�*���e&�u���ya���P�2I�,8a:v�7t���ַem��$�`P����:>�)��3Tk-��;j����S���t]��3�֫����(c�4f^yMV�F�Uo`�U�w[F�j�,/��gbyk���성%���g%��A���&�)��w��M�E�EF�Ot�M�֯%]+q�FY��W�f���Zh`{YOHb�0+�E`�@�}ڊ7@��ywivE��n��{BE[���V®5��H�sVB�ށ��R�$ck(<������ڇ�l��5>o���Ju��!�>>�ϗ�!YN����}�Cs}q�OO�z�9�^w��;�n�!6Vv �"���lǝ�3$+;�bN[.J�8��O��j
F��tzݜ����	GSy�1vԴ���L�Դ���t
�XT��-EӸ� K��ө'l���=uw�ٻ���J'ٛ�島ps�|���]`!�2�\we�(\協0�}kܗ;f���\��iL���N�O����-Z�&����á��+��"M��t�7u2��YϢ�-���s�j0Ǡ�풎+����v-��5(Mr���t��[Aq������Tܲ殭1�s)X����ζ��3���<�"�v���ږ��7���勧��Z��tQ��W`�I�Cp�mP���
�٣J��Z�.�9T��D�	H�(�C�D��;o�T"!��b<@��4s7rv�c1�{)��(-��pn��c�K!:���u��\8l,[׫�f@��]���;���]"�Pnr�^�ޓ��m�r�g.�v�`�f�0�A�c2u���V��y�Wi�=�S���r�d�BN�j���=t�:���R�kY���(�CfP՚���oF]e-��th�زK���&\�x^N����'|���\�ī�-�M=ݒ��2<�ҷ�M�oy��/&\�t��v1�/"xڃ�w��)+Q�ɔu91��w9�Y��.�ut�=\�s�y� u?Y�;[5��u|���uo7R�fv���]CZ$���,,�\�n���U:�p9@����u���`*_'��庞��<T�/ z�psC�R)��o�}�q)�5�6z9[.��P��K�іa��7*��7;$�]]�)�(�'i�mdS�'3�=���.ho(�b��=� ��s:"�${��K-�������u�l�5�<s��[SU�I��S:�����(+6�)Vk!�j-��+���sz���+�XtP���FS�Ae��E�Tg/xuȓ��rO�P�,�S��}M��Ɲ8��x�9ݺ�@^c$��L=b.�򴤇�c�Ĝ�S_RX�����c5������W��+���b�K�ʾh�Z�X����ufᣝ��m�;���n�+d����΍����5��J��`/��xh��Ӣ=����J�Ysq#)M�M�
\W,g�7��4>{�W�v�.�t1 %JJ���F��8G��R�A��<�:� oT����+fr�@�-'�A�1-ӳf��D� �%��*�k8ؤj}�������A�n�(�f����-u=r����1��d�z��Ɏ_
[9;�(s�O]b{��Z�^��r�p�zb�nܹԚ�/=V'�[�M	�1�F���n��jV>ZN8U�:m>E-;q��m鷹OA�95̪�w}H�_L���o}  ��Z3ʛ���d���p��n��ھ��
L�tj
�Ԉ�	�lmH�����^R
Vn\�g+�D�&A��@0$����X.�	�T��V@R�]E��B�3�	���� HB|�I	�w�ʭg�!� ���g��������}_Kδw��z	��Y�������}����/M��������	?D�RξiR
Ѡ��:�����d^�|U�y���d�D<x�
�m�'N�O+mV���1�������[��eͤh�H�S��vB�j1ʱNR0Wa�M�ҽ�f����c[��<B�.7�|\��2H�(1���o��+��.Ė+V	XKMu�ep���K���Ү�n۳Ε��ǲ]�d��hPL)$G�Ca�ַ������σ��(��t�ͼ �q�P������$m���q��-��x�k�
*��J�]g�����*n�ێJ�:Su��^���.��c�-�R��f�Wsq�����A�WZ���ǯ�t�O���b�t��;���f�f��� D��3&���ϊ�k�K��������8�r�F�v3H�΋��̲.Ee�M#}YK��IֵX��"@�\�
'�����*���<8�b��t�|7ˬfT�Df�zk��X�2�됞��eb���Hu �{�f�Є�{�)��;�,�#>[�B��6b�4n����u��\0�����(F�it�Ӱԙ|Fu�*ni�jQ��<2S�̭�C�������e;s7t �,�Is��5f���_4gn�8]���)h��(o��
��Vw�}o^[h���W��U�Z�ѧ�#�c�fbv���K��e�|ީ�lG��r���kv"�&�Mi����QX��!�(�ŭ 3�[��{�m�!l����t4�v�.ٕ86�d�hJ�3��T�Bef.�^%��CK�q�r%{�ˈoi+�L����#V�t��%宻_=1b������F�`WI�,���r�-G�=y	F��(�]S>9�Q�9c��<�����5�#�&�u���%+��0]Q���=�ԃ0��v��J�}�z>8�L��̼ȫ^�-6u;��a�0�b]��e	�([ül��s 9Z��@�!��M����06��ȹb��1��A*���r�o3��|�}	k�p���T7���rb�Y�\:��f�����)SܥJ*N�/;�{/����|:�ȣ!���,ĥCE^#�0���L�qnGI5�]q[�4$�J��^MۼuȮ��	K*�c�5>�à���4Be���D��\k��u�B>�J^���H�\ͼ,�V/�Yj��l�DB��m�w�P�ܺV�3�b�p�b ����W�A6�	��u3#Nn.=��.�x:�:��	z:�2�fnԖ4͘C��M��+X�
j�#�T�x)e��s/����_J �D�Sk�-WVPv`T�7ݱ�hͲ����U�D�NM�LDn�9��ko8%q!|j��Hn���W��9:��vQ� a�^r>h���RҼ��V�2QR���R�}ʮ�U�t��j�a*í�%�����|���E�W��z #(m�U���WƅU!F�֖����hd�������=��7�Ԡ[2�p�e��x{�)��\���H�έi.V@NZ���0�d\�&�Vx���r63�*9{�v�Z�;�]�+��Y�!KR�Լ;"o�(Y�U�.�`X�g��)/2���ޔ^d=�t�=Չ����T���)qr��.4�(���*�M&8��nThԵ�d�.S�Lm̢
�-���ɓX��U�J���eb�֕��2����+��U-��S3��ʪ9K0����癕�dD~&Ò��lbdj�}��_������Vt���L�]�G��c�F�:T�oޜ��>��v����U��V�W�dǨ"�L��������O<Iu���h�*�^���;��.>?R�!���f�����6W��F�^�Z��q��#�;���Pg]壞���a���V�M�Z�m���߱���,w�)��&�u�� 9�ھ�Fp���+����������i-��^N8ڰ�Sצ*J���כ�4���JH�Y"M�s���.���o��^;��G[��<����J���]����X&�k���q�K2K+P�Ȯ����^���S9�~=��y�b^kY{����^�6}/�$���۞2�`�,w�p+�2Qs��l褍��#����h��~�h��(z���њ����]�I2���>Ǉ�b����s{�Aw������~6k���5P_�O�lk���{,�����?WOt�<�������t,C`f�3"�׎R���f�]e���Z�D>��j]KI��q�4������{d�:t��=t��h��:�}b��^���b���y��n��DE�_�H�޻�o��Œ�^��w��.=��.��0�*J�v��/i�/N3ۼ5�dĩ�ﾰ��M{zN!��'�l������3��O7Kk}Uՙ�
{ځx��_)�M�v�؎�������@	^�����"��qє�٭�|�~��ĝ��D�m*Vh�{��S�^�a�3
q������k���É�o��КJ���ؾo��"�4X�a���VL��\��_U��Ai��2����"�
�"�-?��ָ|n��4�:B���i���5����R�N��8Yί��&�f���~��7s��©�<�r���=��y�wl��`h��nv\v���mv�ng���3]���P�y>����*���j���
�xkEr�e|�
��c��~'�����
T�t����M�K�_)Sl���c���y�w��O�j�tuaSW2v����^y�x͸�M�"��)^v*#�G���-4Y���`����HUU�"�t�:����f��=��:��KL��)��B �Z,������4�z�&OY�)��v�W�1E=�s˳L�{�<zgٴ���v��8���a�i��b���{���\zgN��l��k<�<OQar�������]h�=��^�(�awgne���wd��3[�����;s��p�וT�>k�g�p�ht����O|�{Sg`

슘�V>��7o=FNX(��9O����O��;]�ow���G�q4�v=P��^Rw���}�bVVt��gg�kJ��\���bx�N0����{�����x��f�۶xmx궇�qW
z|)V�!� �(NBy����4�����;g7�󫳌;eJ����i��z�Z��'L^]�����b?X{G�(
���1������msO��3^�ѩ�)��ozY�1�ó^g©
C꥝gOv�7�鮬�E��}{�#�Vc�O�P�:LN�_n�}���O=��{�5�eC�L�4��ڝ3��5�:���,I��+=K�{yמx���q:|ISl������4����j�N>����v��?|X"�q��X����m>�;CĬ�����>p;J���o������~ю�3N��o�ݝ�1����q��M����g��,���j��鈣�m�0��R�@�qd��[N�ϰ��J����ۭ�8pq��*� ,&a�tS�Q�h(T�2�㝝�c�5��Kp�.#PӼ7��*�v�A��4�.�W���C��w�[?����~�M�8�v^3�'H;l��j�!��u���/˘Z��+��Lun�m��9��BNt�)��c:]����#��B�D��г7%m^��+�9yo��zl�^��s�jY ��l�D/����2�X�O�k93���fY=���ӎ�0��Bb9G#.���L��l�r「[B���Ups2�(f4U�3ĥ�Sn\\*�QK��+�D�T��n\�Q�S-��tN����yώy�@a��̛_5��]�"cއ�?;A��3��ܭ���*��}HW�}��{?g��_�U+:=�W��ߔ���գ���>�Ͱ��:��ĩ��f���I������x�f�Nn�w�έjE�Me��z�s5���x�0���i�������Γoh%N32�^�	˅�*
B���A_X��۶W�m��Ǽ�W'+v�h~��/�����"݀�I^���a�����ޛ�i�:󭳏q:`�7a|���}���)�״�M!�5�3��^���t)�<v�q�(��o|�y6���i�R��]3�<֎٦g���f;I�^�Ag|��S�׉��8ü�Ӷ��n�坾�O�޵��(e��鞻NuM&wW�S��4DW
h�V��+����6S�ra}�������I8��FK�-N����m����Y|��{jk���16�S���
4³&�|�H��s��=�=���:�T�6N����s�N��t����f��Kw�C�c�:���]X�rx�iS��x��u������ºY�3��YS��T��q�g�ޯ�]t�E=���'/����|z_@�r#��$7F����.5�q�e�� l
BN-J�;5?�
�}s�ݷV�N�l�%AN�c߷3��͝�}gi=@��f��{��:�x`���E�S�����6���|�����"1�m���(�b��-}F�X̎�K�Q0�p��V+�v��Tf
�.�o7��u�����g����S�����]f��*�#��>Zi{_�W�m�V�����WG?Zx����j��'q"�K@^O���[���7��/�n}g��v���uO��q���xy޸n��rȦ���_	���ZO9{g� ���+8מ��3u�gz�!�F�K����sXq��m�T��E��z���s�����1�w���ǈcz��f���Čj[G��UAX,Rت�SOSW�t���S��W������?_��{�S���.�l�uO2���3'�����ݔ-�'i^����sZ��G�|E>-�(��x�m���*��k���&����s�i;Cl�<O^�s���֩�4�1\O2�5�c:g����4��y�7�3����&��wֹ��M2�Ĩv�vy����hm<x�����P�O�y�h8j��)��t<ji��w�����b�\U�w�;����s�5H-4Ԯ����ϰ�*Z29坓��v�w��Cv��N�'��:�k�vΙ-,Qx�ͻNw���k�{={jaX_i^=rحT�>�#�<kz"���������6��/��a�+�S��j�g�z���q�8=!ǉ�Scκ�gL�c�z�<q63HY�w�;C��)�X��M?e�\Q�AV	
p7\�?ͼ��;9�1����ZNd����B��2�iY��]��N��a��u��{���tμ���q�t��D�_z����G�C�+���0e��$���铴��\��o7׻��T�v��wNw�o��1��6�L����i�s�c��AN��;��!^;|�i�&���έU�Ex!��CO��'\}7U%GP���f������w3�d�)����y<C�;J�q��:C�s9����q<gi�zy�9�Z�z�	8�ĩ���z�Ԍ��ol^]�[siL�q��`;�^>�[���#�.�s�@�y����V�X+rդ;�ߟ4��2zČ�S�'?���֏Z�K(6�q�:~.����o�s�6���}������n�؁1=�%a�[�
�\�U��FBX�9��N��g_��j�mk�==Q���M���EV~����+i��<�8w�;k\DԵN��K���ś�FOF�^#c����;ػ^
��T�[%+8X���2dĳvds��W�Ǟ]�R�w�:�ԍ�Oe*�o��EM8��Ys�&���^j�d`�묡.$�đh
��c�AXP��w��4�r�C�
�?����w�w����ʸ�yH+a,Sl��^<�������N��c��Nc}��ˆ�%E����:IW�6���T\���ֆyQ�������:D��gK�ػ37���	$��0)qw*�$��ċ/�:��S��^�n��awb���쏽�_��_[�(�A?��28�«r�r�㑭D��1`��3*`ժ�����ETU�ى�	[[F*4��F�#+V�[[U�E�Z�T,U-*�ZF�D`g]�����|����፬�6�9�,>�v��,V��Ɨ�1oN�}��pMt,z���_����f�HC�t�!Y��ז�Xv��	ā��߾k�$�N� ��{��g�!�Xm >s_�
�BRI4���O}���	���L$� �d�@�:@5�s�r�L!��$;��'l��+$����Wd���v�L
��� ���5;y��y�|9X(��&���&_K芧Yf�Gsf��-��U�7����$��a=`t�m �C~�B��RC��!$�d�$>4���v��$4�6Ö�y�y׺�� V����Hx��ᓌ2C����u��!�)!XI��bCI;I'�Hi���\��<�@��2C�@�`LI&0��$*ǽy}�CĐud��!������b�C�$���<��=d�!�)!|�q��	8�i!�k~y�N0�L��v�A:�����R<�=d=��ώ�I��ԐY���Oy��o���Y�����Gb����f��r��g��EJ2\'����_�x��M%{�5��,��/NCN�[��o���$W�"��T�+9�0Y)���(���􆅍2͋f�2��dZ�Y���V�7Mb�����j���w�_~��4	/��R1)
�˷�nӖ��z"�З�v��N�HF�������������
�������~-Z�6�b���V69��~�;[)yM�7���s�3�^fzWjm�ѱ�<���-��Q�l��z���̳1B#�
�|�ma�䷒��ڨ,�ٯ���V�Y}��n��Q�C��l�ѹ����9vh�����ޫ2s�R�2�U���9���ޗD��������6S�(��q�{[�D��ϓ�:��ǻ��V6�!���2���u�Q�Ǔ%oW���;�a�����d���4PS��+^�n2SyN��Χ*)�臟O\�De�WEŃ��KA��P��.N��5M����:����l�.<.�4��ȎP�Z��Ϭ��������=�=v��u'N�vH͘T6�o�3qb�4C��s��vɭc��I����Y|Flr�L��J��a�����Ɲ�_�[v��#��>YG�8�K	%����G�/f]?z?���W�ϱ:��!�%��GGv��yILo��q9z͏31�z�7�oW�'s��J��e
6W�;�w�./�dp.^JRC�.D������u��j�;�f����.�zׯe���� �����Vk��Vq���i�^�4���i�{��Bp�ݔ��.�_���(�� ���n�a&�'�M��{�[��`��$���>��H�á���\���,��Ě`��gr�'�䇽2��<𷙼��2-9�#�������㘷�@�k�F�ԛ�I_��Բ��=��@��j�SՃ�� o�S�[�F�t����㍘��k�c�#]zE���m��t�"y�i]�-Y��P��.�y�3���epT�;8Z�-*��43���'Yz�#u��Y�"@fw�m��-!]G�u	��Vډh�-l�Ȅ��#}d��YGG[&��޵7uw2tC�'�i��ҰM�����)4l�[];u(
z,y�g���[��.���MtU�%��cQy&��5�iF֌��s�@:2*�(7�Z��L��]:a��ahaoJ�;���Dۄ���oY�T�赗�
��7O+�Μ����5�vZF�ڪ�mA���R���Ԫ�аee�U�R+mkZ�Ql��j�PZ5kE��Ek�KX�R�l�m��[iKj���5���E����.a�XV�z����F��'���p�2��1�V�>T.��~��f,��u٘}��cl��Ձ%ˢ�e8���S�����Y�ç��m��������k&<�h�'��VQ�)���]yOa�꣝~Z�jK�R�OyY�S�^�6!" 3Uw�f�[����eؠO�z-�����/lI�{�t��9��ޝ�)�����e�-����������!F���Z��9���<���� �ग़���*�w�zR�n���2������/�jDc����}h#}J ��Gt�x���y�﮳�һռ��`9DnIe-��̆�b�P�( ��י�l0��v1�w��*1̹{)>Ml&�HW���G{\T;����_��?�λ��~��p�'ˏ:(���ԏ�Ok|��s���5�8vy��B��5���c>Ԩ
\]כ�gs��qg�>os��;0`�#.ܮ���M5+T���yʤ	��b�_��=H�OP�/��M�ck�:��ǀ�\�E����Y;�/Sso*����P��"޽��}'��KYwl�}�E��q6�����6���	Eŗha%��XUދ�V#�R����F�����ݾI��n��!�2�[���������P�V�O���E<��@���=g�R�;נr'�|�CzU�������|�����L-Ե]�QʐV7-�}��w2Q��J�0�?���sH�����=�m�!��^��z�q!�1\����mf�w�87	Y@X�n�:��ĳݾ��9�� �1�ex���R,zuۿv-��KԷ��?ͻ�9���r~��(�߽�W㾙F��?K�iT���` �'G�5j+T���{���{�ޮ�@؃c�ڱ.���ޯ*g+�n#��439o/R�9��B���x���u��u���*LRE6�K�e'Ql�9?U}�\.~�F��~��q{�u%�~�)jo�	[�R���\ڹ8e�2(�Q:�
`9v4�*����U�3�`���Ii���k�|,!���ɄY*�mK7ݗ��50��)Q��'���r��Q�]q�I�o���zt�'�߈�W�S
q�pC�u�}�D�:�����m��2��_es�l7uo��p�~c�����t��-��t8��`ދ�f�j8�Hu�wM:��	Y6��XfƧX&[�U.�w*S�(�3 �]��C������tɆ��0$�iY���H�{jVb�Ɩj��)��`Ϧ���*�(AR���}���\�؋2ܦ8�v��y-�o,��X��c4WҷPC�s.�D1:��ݡG(�\qix��C�\��Z��}b$���<�MX��A����޺�8��G����X�1��g�s-ZN\bV[8.=�Xsf�]��iK9أ�aD�#���3;7��8�<4w$��v��$�|�`{ze�����I"����qj�ˏt��O����b�R����k,PD=��-hZQ�H����ъ�@E�"*�у�u���~�̵�j�9�?�����<��Gs?r�\v�8|Sxr=직~��=�, ����h@�(�Y��~H��p����(��(+�Ϯ�[O��L��1z馢;w��v�B������\�6���=��m�Ҟnt���kQS���N@���24��+�q��^�z���𡿵�D`�1?B��r�����7Nԗ�1-�J�O޼�X��p��$f�����=b�r�������5eh�dg+>�8�֊B���ޙ'�c�[�V���t�1��HqS�c2T>il�n~������^*����n����)�*�TE
���ޢ��Vi�E��
�9]��7��3�� ���Vky��}�{R&���0s�Z��&��=���粍{=�|K��a�/rì[�ᅱ�����7��ٳ���T��L�'�WX�p�~�^�:A�Z�	�u�mo�q��C<�Yz;��8b}S o���{P�����rxk5�`N$x�Rh��}m��PQ�J�,�������Ռɾl�P�N��#`lҷIB����f5	�gy��}��yh
e�H���^�R�� ��@�����u�Y��ap�M8�l�~��ν6��<�"�Ȼ ��8V�N��t�-AT�__&W���b8�뇎֩�6F]X2���P,CXnnw�_}�}����~m?޻b-��"�{�>A;�ngU�f9�&<��r�]G(���G*��h����In޼�F���7��-�5͡i����4���ǜ�͋��q�{����F��x�x�oa��V�2 �d������W�Ƣ�{󡟩1���൪���wB=oŦ�\���Ӹ{;�(����2�ɓ/��>�)=�\�hyu��[�C1ȡ�0��^_�٦
&ny,���X<��V<!:�5��������w����q���8�����n��e��m]{6�����@r�)۝<�����̳�C$6u�G�Iv��/Y���sF���{�$Ӑ5��M�3V���;��]�z�)��.聻:�tW�K��c�ԍ��9un�>���$袹9�?����䴯ߡΞ�,#��D^8+NA{Ѡ�uؘ-�Ǜ�z������%qh;�}��G�����7�XO�Ŧ=Y׷���GØ�F���a���[���~����'��E7��)`�4>o3{ۻ|}�tJ�W�e,�u!I�45:�{�2��j�zjh�_��^�y^K){Y���I�j�k�P�j��,y-���l��1=�q4�}�]����_®v=���ߝb��ۙvfӾ|�v�Fd;���!	*����SX� ��b������ǝZj���s�%=����X�b�`�L�յx3`�9�+��3��AaP����r�c_S]sn�&Ȇ�k���;�Wt�2����B+�&��R�$��}��A�-��L����Z�۱�ԫ��4ch��]A%6��;6�U��G"�AwK�z#$w�R�2���h���`��h��;�%NOF�<CK�d*;�9��9#Ul�l�>��A�ˎd��Q�I�� �^����8�]�z9}:�L��}W\r��هB��R BhP�h�H�[jZTZ�Kkb�EcUUTm��F#R�0U�mm��R�YV�AKmF���#EQ���j���P�@�F�$���s���?�گ3�p$���UW�>�����u�������f���&����h߳�!�ͅz�t��.�d�F8��}�H
ۊY�����x��N�������`��֗�kmYp�n��"�~�:��K���&ʩ��J�^F��N�>�y�����s7�y���_�ZmX�����z%�t�|�YQ9��j"���'�sme���w��᫪7�����<�=0`鹖Α� �ݖ/c��h��aW��E�Uo?��Y�m���ݷa�  >�������*�j��4����i�Z�#�YZ��}�DW�]|67�e��j<;�p���q��(�����|y-��e�,�m�%qܒU�h���Z�k �c��w���8@QΤ�O��ikc� -����ꯪ���/ߡ�O�P-Y}���Q��W�<��a��r��o���׸/�fW�c!�i�لM��V41HpD��^�lp�ev�~waA�����cuڳb*M�C�έ�^����y˅�Wn����)	8	h|���[�^�ٞz�5)�)� �~�������+�������HcH��o��#&��-��S�pG2^�S��\x��zK~[�K�-�t��:}����s���J�K�x*Nn)2�/UZOP1a;��Z����{خ��1���_��Ï�3k{�]jX��[���$���-7�����Қ�3�`���.Cwcf����9�=��o���=YKK���{�n޴�˻._�p�.���Tkr�H��1��{S����JDTX
֟{��o%4��@�u�L������]�h�>F�ec�0X]�w��f<�J��xI�|҇6��禦����h�҈��Z�:�L�������j]����$Cd�+/t.Jn����C�mX�QW��[�j7$i������_S�&N���.�Ӽ��i��=������6�N��hd�6rg˼/0������^�a4]1B8�x�2��A�����áŗ����b�i�̲�Y��Q�c��܇�7
2�/mIn�n~����KW�ۂ�֫�g�o���
��QW+a0�uh�W~��C����k��|uAOu���Z(��2u��:�+"��"��YٕNݗ�����5;H�sLh��R~��~�pZ.^T�ʴ�`lbd�����o-̿���u�y�V���'��ỵ��=�^Kt������e�I�`���o��N����j�=��u�)�[Qx]nf�J���7Cҗ�%6�bd����.U�vx�g`��4�8���;�w���9�S�@+޸w�5�`�ѽ�R�AQ;�'b�&>$��/Lgr�.�R�9�{�ؾ�h!j=a���cK�z��>�s���l�+{���������a�q�A�ζ�%�v�^
���;������D�h7պxqEz`�D�2�H
�R�k��S�+���E�Yժ�(�Q�B���[�ڐ�V����s�� gK�f#�Tg��H-u�a�%�JKL�}W9Q<�/+z۹�$n�)I݉V5ə#��p9�Ad
f����|ӣ9����b�+H�WWw�e���ZR�m*	[iE���XZ-X��Z��ZR(�T���6[DT����ڵQE[KR֕U--FYi[Z(%[[D��[Ub!mX��ш�kR�*ҭkmcjѭm�F��UF���Ts0JZV��,�r�[AnZۭ��,6�T��-��y����!��%�U��Y���Uo&I3��wQWx��w�2wu9�F5�"'E����W��@��[����<��ik^�#t�'4G�c��"�U˄���	���^?��a��|/����)�#!62R�[�7t���y�M���-�'��9�V�{zr��,�\��>�6�ـ"{r���+Ea;��� �X�K�-��@�v�²���+'-)}����z��Gc��X'�1Ҙ�*o(��c�屰6i[�$� ��o1�����T���	@�ܿǚ��Ռ�mL>5��.`rp���'3h�:��+BgҎwYc*_Fuw�1����_Xt<�յ���l-:�b�w�W�eR#�w��C��'��E/�]�{�+�r�B�@�̖�*Q�������-?�ޏ��\Me�w�"��n�E��� �[�Z4s��m���g��}s��f	zqo $�Cnin$��p�� �S5_�pz�9���������G�P���R���hz��A�$���f���5��E}L�~�"��g��nE��t�GR�(n�g���w,�.�&��0�Ğ�������FlN��!v4���mߞ�[zM��x��=|�g4��f|�^��A�}8�S�[�N0ѝr8��U_SmQ�O�>�YX���)e�2���{?>=~r�t�Z:�q��9���N��	f����qL����\\�d��ފ��2�l1�D�����o����t��e��+�4l�*Qt�'���Kn�ԍ�bj��f��T������u��_��Xͽy�pK�����[���Y�v���`�)�#�ޗ�9�g�<"�}}8��wz���v,ج^���[h�潯��hX!�s���׸gG��̈́�����Ő����f��U��>������J��5���' ������[�oC��9Z�݋$	��En���0���f���1I�.���Hn��U��H�b�~��67��/Z��{�wP��y��I����øxs�.�_y�����6�ﾪ����{��t#�C\�&�3a���N�m�Z����j���w�oJ�^���%�R�v���K(�*����N������bn��| ��J�{�y��~�����wg{c��Lɏ2�� ���)!5�+4>�37�s;�}�~W�|UD<^��������w�G�?5hE��,�]�c��=F�� WC�� c��츂ޗ�_��kF�WjY�|6��=ۄ#b}�yc-֙ ^��Wu�~��=��n�v�\�[��|Z��elMXu'i��(�:��cާ�D���/koxO�{����GCqt���T��MҁgÒ�p<�rr)}�φ*U���;��(��5]�B+�N@'�"i�b=��D��Y�}EL�6��ujfwwl"7(�a�fh��НzK�f�urŎ#4,R�V�Ĭ�%�+�ކԔs+�����r��OQ�+��F][�r�	}��w�a�PrES�j�[�ɝ��p�׍�7�R�_p�nd�5���`�4M��/ml�kh��7kE���#��M϶�Z�Q�\��TB�c�֗"e�(%��F�pY���նֶ+X�Ym���FԲ�*���*��Ѷ��e�2�*R�U���hP�r�mj��m�V�E�mR҂�b9�b�mJ��RԵ�C*Ih�r�����m�Xe����u������ܒ)'�U�U6ͽ��Ncm[��[?]�ry��lz�_�3:�K�AOؘ�^k��#ޞ�w�離�lo/
���=OC�o����Pyh��ѐ����ۀ:3漮��ޕ��
�e'�$y�vT��j�d��꯳�?~��<�B�a�:�-����4x(v.����G��wʝ��6d�6�+���/q��W�����g}��&�S9m�ݭ��ʼկJ�Č�Z�#oB>����[xC�^���O\Г�nl�ʷUk_`l
BD-��Q����?rv&1^7�=ͭY���om�*�A�ў�d�U"6.d�*��Y1p�4ʮpOn���̹t�1M�ޖZ�{���>�(���V�h��[�P������G�)��NO�P�~�j
��ӵ�<0�|���|yL�7?;Z g�Ă��V�h�9�ޛ=�L~����(�Y�/iO˙4��	Ǎǝ�ʶs
��k���CT�z��\�����%�ה�a�_�8�	�R�4u�Aha�{K��	-�JR��~Hw}�u���5,�*�1��_n��ڞ�w6��C�x%���y���ރ�k˙���s4�繬Y�{�o�NrF9ؔ�"k!�ۗ'���}~�)��ěw'.VfkOV!���#fCt�R�Ac<8�Ù��a;����k�c"��{��gf)��>�Nr!�[x��R������
m�M�t����M�$!zwsi�1W��C��7�^�clgw����i�`��A/�`D��TƑ�gZ�$�R0\'O
���{�>����@�/n������57�|����w�#С�(�jf�>��Ƿ�"���p��3S���㛓Vw#�?5b�TK�y���J��ӎ�α�q��N���T�m:�h��^�6�Y�P
�eژ�W���ޠ�oV!N9�w��&���tx2��-�"W���={�n�׵}à�k��d��e� 3��}�k{��aA0���?b�M���)���#�)f�K:y��t��IBNe.��q�@\�ɿwZ��d���Sqeidf�^D%ݺ�i+�g�9a9��0)nL=�^{���V�ɪc�f ;-�!◯mp��� ��W��<Jφ�5<4���{��b�d8�JN��9���~`��:1l�������]�ڈ�`�g��]F�:]��kN�99�s����td�ڱKT~.� ������ܧ`G1+=s��#��oS��S�zQ�i�������ʖ_��o`�y)�j6ݺ�YI�؃����%u�:�=�yY�,p���l�2H�6�7�T�A�=f���6H��P$[R���ܡ:�7r�[)r��x1t}�ɖ淚eI,�ۂlM��Yd�L���sP�5X�X͠��s�}��v3=�~�>�ɝ��3�Jz��e����,㚴`B�����RN�����\��f�R�Z�k�l�悎�:zqj:LIۧz�n)yGvi3z�����$)q�g(�����r�(Нc\s!�p��J�Ú��;��2HgQ�j產�%�eC�YUU-���-��%E�\®4�Z�XѦ4C��k��G\�r�p��-�J*6�kL�ʕ�fX�l--��q�m1�����m��[\0�r���.1�pZ[+D��[��ƘJ�TQH����3&xޫ޽��\�I"ۡ���NX���w,�g�J��4�oOR��w�5ӫK�Ś���Y�"lf��^D!����v7�a���;zS���8���8���X2KB�o`�O/8��Zn���be�-@�� mBp9�We��o�.3�3j���-q\����Z0u#x��E�i�o�no�O����P`�V<G��["�݀8�c,��f��հT�),�H��3;*��[������z��e�́�&A�Zb�ک�W�gM�<L��vX";=��k�i
7�ׅ�{�lⴭ��^|ߺ��/�:%��x:ִk����ӆ;]��NS����g^���˵�x_�#ݔ��F�U=����#��1�0��N5��1h}�N���X9��������	2��Vo� �ΐ5���a�G��e���N��i��]�AY�N�-���7�o���ԑKg;�!���r]�ݞ�wH�Y���z��F��ӈ�^7�\L���"�Ջ�7w�0'bqK
��.�wj�8�L4���љ���5=��e�����~]�"$.�pO=Tt�β���Ƃѥ������Wo�������Qs��l蜍���=!w�ä��v�f��{<0��r�\@�@������ ���]�����)���w��W#ӷ:Cl�ܝ���df�SՂ���]O�����WX[j�Iij�]�^{W�y��#YR�����;�f{gV�Qe(���E��G�l�����1��Ҳrb�A^�+�o��������1-�]6>���:-]�箣��j*�9�Z��Ւp�w�L�;�JHc�"�H��|^֙�{j֒�c�wY�,�d��y�ic?L�k�x�=�VL����ًvMh-�~����=�J�ۭ�h����~� �⏸�z�gx����e��2�G�=�p�D7q�:.Ys��d�7G|ޠ���\���!�,�}��,��w�i��X��U�O9�	�q9y֧z1��ȅq'SZ&5�	��ƶOS�~���)����y�AX:v\��݆Ck��v)X]ĂyB6T��j�`�N��9���X�{{;���������$�����ds���8����VUY��+#��z�>�<�y�wy���������Hf4x���?�a'�~��V�a����z)��d�:h�zU�y�F�wn�q^ބ�&��=���;�h4x�G|�����e�lp(��4�wӬ<`Y�{��bB��IT�W�K��*IU�H5wڻ��:��P��!��z���J�:���&h!Ϻu`���48��P@E��$<��G CU�k&�qq� �n`�r�q�!ܡWXep�][b����ֈN���;�P� ��l'8�F�22�� �UىF�ʻp�ތ�e_;�;��ٽ0��L�.f)�6<}�|����ݲ�L��Z�s��k]h|�}7[����*���A��TG3�0�Z�V�Q��E���L�fQ���n\�ʭ�-�qi����6�2��hV[m�\pe�%mj�be�G2�ڹFZ73*�\r`fR(�B� �F��B�۾�S�8�_s�I�5h����&�:�x6�ߢ!u4�U��4��A��>��d�׋�Io`Ub�P�a�O��Y}��xڧ�pu�wQR�>��hｆe���/�.D�lC��o���Q�s6[�`gi���̝n$�����Q�u���߱�:�<a���#��=��2�v��N@��9���WI{h����k=3�lv��|�N�v�_Z�Z����i�j���\�eeߎ����+��U��k���1���2N�O%o)s8��Z���d�tp���$�x(�mڞ���Iw^\uiWͥ��������Yc�'!�����Z�T�wiF<���f��oyM�:*C�AW͝\�����ӻ���3#͒9#HF,��V�*b��[�ooӅ�6��+]y��b�Mp��k�����9QaԪm��uSui��Z�t�wma�P�y�xy{A8��6���w�O�e�'���wn�E|���ʄi�s�J�ڹ.���<Nߗ7�j�Ԋ�ۣ�4߸_gI�g�[��
��V#����0ҧw���yX��0(J�����y����3=�i3���Ci�6�����b�W@��"�����$��ř+���Ja�-�{|��-7�4�;��8�*m=�m����LL�w#�-G�����S3��V�k[�{l���j�/FCnn����Z����7ա߉�Qʔ�1X�,I̥��οza���������xm�19��sz/.����6+���@[���\ �W�����^=ڎ�8Q��w<����@�����6�k����|3%�u�;�/3����2��EE�l��ǹ�[|�/k�5l����^�Ћ��� m<��U��ih�[�J��<�X�ej� 8)�U������He4q˞}���2mmM��_�5�d!xK>��R�̻��p��dR4N;�Zs�����J)bTܤh\E�Ez2��^�	�y3�t�Gn�u�f�p�˗%�ʝ1V[x��}�ں��я�/z�| ��������t�}g�ײ��PH闖��	R��ۄ��]N�ک�}B������W��e���V�~���T���{��]C�eY�zC������ן=�-Qm�6��'����Wh���œ�љ]C6���~g�~A��
�m+UQTR4�r���$ �'���,< �>V�0Fp>?�0�h,�:2gw��Xi��a�?����OD�tɴ6��n�!��F�����!"��M���Y��ą�P:?�2��3\���p�,��a����` O�H�7�'��S�w�������`}���>�?�DL��f�텟hD7��f�t�w��:�dϑ�r�����oRu�#�ǰ�u����	 �'������3�~�<��$� }�@$	�������&|>���~D>E���'��'�!�w)��,����~Sa�C��H��~� H������Y��p}�b�r��$���?ZL	N��HD���Sf$����Y��!�������AY:�/���~�rS��e ����g���ˆ���@���?S�$���<�,��S�����^���C�>����~� H�'pEY)�N���s�>�0�Y����.#��vxM��ч�>����� ��|?�~���)���?v=}��������	o�%�����!�8}�?̇��@���
�>��ҘO`Y
?��_��#�w��.����}��v��g�I�N~�������? H���~��Ϸ�~� ���|�N��a�`���P>?h~��Q��k�	 D��@���O�'����C�K��^O�J-w��;7
3`̇�! N ��X ��2`�t��;�_�{�	 L�''	�	!��prM�������ÙZ����������s���LIi'@of�����A� $	�?Y�����d�� 	:���'�$�}s��@>������!�=�ȇ���d?�>�}`H~?�}�|�R?�?B!��?PO��|��a�a�HL����k�~ϔ;����"�@�q�O�����$ ��������C�?� ��? {��?�������������|��	�̇����\��Pd�~T�Ɂ1�T?� o�~�������C���ܿ/���y��鯠��? �� ���H}�7�o�}�h8;��60�O��Q>��>@�Q���Q�C����vl���$�!�~g�D#$@���?�����?�C�$?C����g�<�'��I �'�'�?Y>�I�h>A�}�}'{��w�?<��s6rC���� ��RC�|"��:����"�(H�DJ 