BZh91AY&SYŏ��<ߔpyc����������  `�~�K}�  � �P  
�(U%!��
JJ$D�(
  �@���k�<   �� �  ( P ���� y��{���4�l��t���q�|�O�0Ϧ�n�;����u�W{t{�u�S�ܵ��0_f�3�v ����z��/6��˼=����Q����|���:�k�O}�������y|�/�uk��������s-�Ols"�k�F� �=2�m;j7x]Z��ݷzә������vΥ>Z��[=���\����֖����ý�r�m&J�����@R��m�֜������m�um�o��ﹹ�|�^�=��֞�u���6k���o �� >�{�w.�wn����kK�Mwf��;�=���> ^�ܝo|w�e�����mxw:-��x    �      ��@ ���jT�&����  @ 2��JBJ@       )����� M0� 2`��@��Hh���M# �`���D�J�e0CDё1�JxF�ڏI��Ч��HJ�hL��  0�>_O����%7�Y��R���#���$H$vH�D@)���b*�'��P�����˔?y?����B�TH�'�T�1���/����ԍ��=,��m��m����2�I���?'�'�+������Y�����6kF
���1�'�T����SX���j�d!?��k����ç5���XkH�0� �&k�5�d'ң1u����,�2i�:n�2G#n!��#�}Q�8�gfIR5�0���+�������X��>�2"#:���Έᾈ��5лeZ���P��ס�w*7�`kY�b��V��Wm��oڳ�
9o.h�
S��wI���P'���;�����7�沔s�Wp�j9�4�ƃ���ߧA=�h������N���՟n��d-�x�'+��2y����
�`o��ܟJ*S��<Q�b�gn�u������;[{�ɫ�kK�LFa��|�V9;�bړ�=������7��n#�1�;N���UDj�B�*ǃ܈kQ�C{{Q��fDE�DXm�v8�	S������Ю> 4,�S���#P8DC�#`wWY	�|b�>�]�e�;!�OlݖDI��E$��0h��Ϝ�A��E�_8��|=�-�E\C�"�s�+*��60�dC.6#&b3���l a��w h���V��*�n�'M�0�<9�!�GDX�vk�l�.�C2�P|.�&���F�f�H���zCa� ÃLQ�i��rzC`ˎ��N�D�D2�*�#Ġ���k�o���q�����}����gk �3܈������65tLD���s$N�Ұk���c����C�`'��٬�s��q�ːa�18��#��89�F�88pgDF8!�΢9�C�#��*ʦ��
�����z�/,9A�Q��b�Wr�0��.Ɂ�#��啥iv]��qnHv9;�b�pR��D'�5����ۈ���giѱ�����/���D<Q��C�lu�"o&"j",���,���n����p�"44VZ�)�tC`88DE����AÞ!2��[#TffX;!��bl�dJv[9E��I��\-M����6	�"�=19@��W���
���' �����b2f#��]G0!�ddpB�=����3Þ��qGj�|�2u��M>۬=��W�Sl����OD���!�5��^i��FaOzc�"B����#b�zCa��D9�=�H�|�;��<������N"mH�U�e�!�{��;Y�a۱�#_D(9��BF�b#fb��`։��ܞ<�4��ں���o�����rts��pC�Ӄ��%���G:������7�Nq�t�Ds���䑀�
��# "��#��#�\��؍��>YwE��cM��IR�+�Qe؞SП����+U#�*��8��G���O�!p�""S
T6Z�Z����Ս"5�7���dCSf�Om����^�8�>�¤�)G�ȊzCT�"���V�V�)���k��`rz!�M^f�i���#����w�Q
�P�"r	�է�-ѭNI1?�_�8!�OJ�`Z�N=�TDMA��Dm��dCQd'�'��+T��j["4�
�P��F�!�xGXթ��6D&����G����.����])R�"^�&�\�[�#q���dE0�!�9=�N�"�i�\C�G��?��mD+�-�ai��'�.ѭs&�B͈�pC\���L5<�&���i��d.���r[DʅrZ�^�=!ى�''G*k�Չ��>����'l��DO ��J,sd|�O��h�D"�O,<�,ߜ�d5�tz�pp(�jt5�"9��dD2Ȅ�;��������%��O�ć���>1���F���ȵ���i����p|�/��/Jߑ����Ŧ�&�z<����~/�G���Z��8!r5J������g��?c�F��hk��|��J���Z�M�5t�!�ȞD<Q�N����Z�=�}H���Չ�T��a��Mr�P֡F'�@�ȇzE#F���G��?�im]�ȉxF�j�үk]Dc�9gdF'�X�,|CX�[����a�=4�����ux>Fy_6Z�u%+�U|�'�!��Nƭ:ԏ�L��_VN>���5��øg��:���5M�_29j�]-�F+�/�>3CC��Q�2Q
Xt�ٿÞ���}�É�_XCIf���<r�x�Xpv]h�ˇ��`SC�,hj5��i�U
��<r�z�r��{�f��x�&�=Iꇫ����Oݮ��ѳ�{�0�?�b��?��5��Z�B�Q�CI��d(O��V��յ����֍YʱZ�I�X�4�-i��J�n!�i�i�臓u�Ғ?P�����B?FS��}�����R�H��=��g!�_ȅ�*5^1�lh�q�ݺh��|�q۶�:{A���t�c\m�w׍U���:A@����+N�9CZ�ޙA���������8�Z��3��� ��K�(���>Xa�3�S$�Θ��;{v�n���u1*ݻ|�l|�n�<m����m�5��漬m�D�!׳�$�4��� �β(�o{\Y��OV��G�s�8�
'zWl|�N�&���e�8�<�YG����<ideK��g��,g���o��A�I
<i�
 �#�:�8��J��V�N�����
���'���7*|Qg�0��Κi��[s�3I4�8���˿ͷ��'P���$ �(��0χNd���ʢ����<�ic�&}��W#O��U���Wt��;54��ת�+��|��/W׮���<�E.�x����n:|鍱��1�ݹ�nf:qێ�;|�{�����CMVNK��=t���x�>x����=.I��m��K0���qߧ�*>�=seM��2�4�Ƀ$�ºlgN̚�j���]��FO^\�vPy��t����̫���������kѳS�`����������3��Ǐ�j�n�&v���W=x�t��v�+����t���:iMQz�}:Y��8�Q���8��j����8��جt��]��c�]�����}c�<z�Z�t鏞+����_]=z��+�&f�n�xL�ݲ
�N�g�:��\?GD*������T�9Nt�f�3N���]8ju^�I��ݱ��Z�_"�m����5{~z�=t��^<|��8��rv�/��v�ݛ��]W�6��������ݶ�]�v��m�c�;��y�}t�2>�c�y��j��N�x�K�:��F��4Q�I�4�q��+6l�N4����9�	鐁��R�t&q�r�:�^�)*pں��bj&+K��|��z�m�cǝ�{ٵ��!���'�Hu�T��6Of*�ܚ d�9�rQ'�ߝ���M\��N(��LF8�&�I~���ӊ�6k4��8�g�]B?:z��v�y�Ӝxd��}��z�m�b��ˋ2񥨎���>g�n����M(〓JwEE�]l�i���q�L���捥d�yv��]��^6�������om�����K��F%c�0ț���-tWl�20�MAצ�T�U5�p��V��Ω��_(0��7��8�U�C�囑y22���,����W�V{����V<u7|�z6�D��RVl�f#�w�A.2� �M˺i��꽎�w�=��Iu$IǊ8�J㺞l��ruK���v��4�s'I���|����ksW�������Q�ԳG�lu�S&Lt\�NY$<��)��d�ƌ�����_l��Ȓ�7�g][\�Bs?|��K ���%�lWx��]��~rL_+=vq�%�e�@�z���/B�I��Y fG�}�2��K,�r�`��:�8�����S��~�_d�I���	�id�x�Q�n��yc0�dHq%��+�`j��/�"X�>��(5E�s�$���� ����ȆY�w�_Z�Sr�]Ae�/�O����E�垎.�ve�.�t�8�v�,�Qf�}��v�Ë*�.��/��f�W3$V����ŕ�:�HǷ0USw&S�(�&`�eK��$���Ң�4{�+=���2�[ZO��:���֛l��U-C7З��������/�8���g2�>_�NY�]��,�S<2N0����Qe���#p3.g'
���;_X���#��4��w����i�6%�g�A��Xq��mݖ�ݴ�3�s�i]k��Ϙ�f�ȒJ#�.�ѓת�TQ�B���J��S1�u`�+2h��cf�A������vN�w��j}}1
9lL�b_LE�t���c	����Qq���aDI�/����\��϶g�/�0EL�ݞ��0�	��X����%��x��z�ڭy�|y��Z�K�^�cUm�6�׏����m�n��(��:�XT�q��]6�.Uos�t��^q��EG�\j�t��Z8�Ӷ�Oy�ˁVۭnèm3Qv��fr\V��Nn��� ]�o��m����Z���ݡW'x����q�#��������5�8��ͽz�F/~�ڝJƸ�w���q�g���Zw�����'��V�;9(��x�j6�yzV�����o�auY�;<���?x~O�?�������t���MR?�m�/��$�BA���~(��non��)��"~*^x�F����/.��&�Hl�3q�>����Xޅ�1&�:������C�*��İ��-X!��ayc�a��F�+v��v�%l����G����MXք���[�;#͠3*�`pҎ�EP����w(
���1���Ҽ���;@���h�e�8��)A�}g��}xP�g�>�:����x73���[��.�h�f�c҄;�{7�M�����ܐZ/V7�zN!�8$��L��� 4@�n�ԫ�����)K�]^�yA��E1
-��X�M�o6�{dAkct5��9үVޤ��v�4h��rꎻKiԥ�x�D00�,J���8kVW���A�8��4���eӧs�p���i<�ZQ��Um����h��͙�"c���ԕHfTR���Z����wY���Z�r0}��|J�;J��dƪe˥�.��A1��3�nt�"湌E�t�@%w�q
��%m�F0��O%WR��]ݖlO�yƁF�~�K��p���g�B�}�� ��>����O~�������A��`���g��?��_��?3�ߩ��_��w_ѻ����pܶ�浶�o��m�m�m�m�M�ݶ�6ۦ�v��ܶۦ�vۆ�m�nm��6�m�cn6�m����m�n[m�i������������s	|����%�V$���#�_$���Uu�>��t�n�p�m��M��o��m���m��-���ܶ޷���ܶۦ�v�r�m�nm��m�m��n�m�m�m�i���;�����oF��%���}�/���6��[�m��������m�i�m���m�����z�6�m6�m�p�m�m�m�m�M�-��4�n�m�i��6۶�n����n���;��m�m6ؾK�ė�}����(�{�wU�{��m�n[m�m�m�m�����o�m�4�m����m>m��1��o[��m�n[m�m�i�۶ۤ�m�m�M6�or�s����wsn�n�m��>K�����������m�����xۖ�t�n�p�m�m�m�����c��o�p�m�i��m�i�������ܴ�m�m�i��xۖ��m�p�r����w6ն�66��_$��ۻ�m�cm��4�m���m�m�M�-��6ۦ�v�r�m��v�r�m�cm��4�m��M��7��f��|�&��m�pۆ�m�m�wuwͷ��o��0A_ �"B2$��>?��|��UD����������`����C�}�eڿ���ONϊ��͛6۶6�N�m�m�m�ͽmⴭ��fͶ�����ڶ��ݶ���+��|��m���6mU����t�n�v�o=m�ͱ㶝6�o6���m�o�|��ޫ�ݴ�M�[6lٵv�m�x���;i��b�lٳ��V�iӐ�_i��_+A��-n�M�F	��wm]�C`j�mc�͙��.�P!���Kl�T������=<�p��e��ظ�M5u�R8˳v.�X�B�Ա@e��STX����6�]�t�M�D���J��彋��6HZ��Yb�m&ѱI����Kk�3.Ya���t��&�kQ��mm��Z`�3ü6X�j�V�-[Λ�
�)��f�lƘ�K�i���{���XMMr�n�e�N��F�h�
9�]l�[�ܟU���ޮ���t�an�ĥK�Q�ܦ]� �m�m���\���7#v��l#�SPF��˫Ha.ƒ�+���vMF�X�wUc�ғB��1ک��vf5��Qք�i�me%աol5���v �5�m#*R.�fH�u�q����Dc�I�(;�*F2�MM�m��{���_6	`�U4#n�����m�h�u6�3Y�l��Y�be1H���e�f-�e!#55lnc X��,��.�bI���ƴ���З[Lb��jm�����E���[�w:���q��+�뉱�Y����4�l�Bܠh�:��)4a�a�i���Y]���Ms���r<�
�g�(�8�XV/[��T�[Mz�/߾�_J��6�������l����-�A�nn4r�L��[u��lѸܭt��rJ,6ݒ��s+@ٖ�ِ�M�b�44�.��묥�Ҡ�����S8)P��{{�z����6�m�h�In;�D]JэU�v�6��6׌\͛F��SVkM2�麪fc�+qNշ����L]�m���0�v�����3ȇZE��d�%i�jM��~zʘ=3,+�8��bK���;.&,6e�CL;U�I��e!6#"Wcav��@[}�k�KrM�4����H@���,h^��>�������&�b�Ps�[VL�!�`�j^�?]�>N�����61�mt�F�3�q�cK��V��ô %�M�YF)A4m��1v*VC��'�[H��&v��0�!�P ��\�ڦ���@���mΉxA�!�a`�k�k1���Ҙ	R�Q���di3v�vb�JI�:6u��K�2\��=aOl�,%�5�Yt�O#[e�F���f�)@����6�Xۦ�h������ڕ�:�+WĠXwm��nb�Nf���,��ZͶ��+���ctX���`���c15�SX� ̎�hݝx�6m��l��Lh�\RJ�%��ii� �\[�`�
f�ɺ�az�΀�*�v�%�ɕ]�E"�a4.h ���U�R��0���]-í^�JCq����-���lK2v%j��Ad��LZ�c���H��K���n�+�Y�-��OR����4�c<�B�^��D�v�]��Y��0�/0�,���l�sr%���7IwMGj7u$"�Z#�f5�i�`�Զh`�F�F�u�[�G6l�I�b�J���%
�4�Bw�ꪩ�����;����1��w�_DIӽ�{�cs��[��x�9�u�]uǼ���{����n������#����UU[���E!Ça�*��q�c��>�|tg�E+Im�6��Y��,!���=�_0[
u�r��
�C��	6���S7hq.vںj���t%�����̎�e�ٻiR�JM3�E򭅭'�5E�8��`hv�h��-�06�Ń�2�dB��8�b6\m�f�q-nZ4���[Z�2���<��6"����O��D8�h�݈�C�Vb�Z(m�����1�Dy��e��1{�+���J��/n�&եN�0	e�c�6�8�&���ʚ^�_�s�t��*��� ���b�,��G4�%�)�Ac)kF�,�D�H%m��#!i�*������I��D��c$�Hu�F5���B�RK3-��HkF��E��Q=Y�0~��V�[�;��e��=���O����P�,/x�M������UW�z�(�W+$6.Ӵ�OgL��=�f��-�|m7��'J+	�y���1�q$���F�,ke˖��$Mh�S�1��nJ<I�qƣt���Ҫ�z��|���`��P�b�y��g�X��&��)�\-������]n��F[e��Ofb9v7�eM��t0o�&�S�;|S���T��C�/fk$��;Mb�27O�a�UU�B� �yz���d�[:8�zd�5(
ӫ��yiF��X�Kp߅�*��x��f7�I��b4��xz(�t�r���̣<"+cU��X��t���M�����&����ֽ��e$��9\ҫIB[���[qkj���eJ6&҆M4�#��6�guu��6�b��:���e��2�K�z�hjR�#
����Jه���.fUUL�E�q6��@ݢQ��Br���0y���-�.�eukg�˳z�����$��ȯc�$��c���tr�J�s��M�SN����8"'MB�*���� ��!4��tJ&�H�w�g&y�Y�SḝTX�*�h���u�W��W�}��~��A�k�2-���V�Y�,L��4g��� �SE[E_o�$$���sƚ�s��G��1ڑ4|YJ���I'�ʘ�P�6�%M����I���r�Rk��,0��汻�DM��KK�Z>&��������]0�����ˇ�p�f�a�5rSUFL�9r�8��	�N
R��}�<�n�	V�o0`Rь��J8]�ų��$�,�E����]���TOy\)�|b0�Q��`J��l�˽W����w��9BbI)����.]�	G���5*T�R�h�߮
�rr����{y^��~Iϳ޸���ˍU�]�h�g�f��ڃ�f�e6rd�RfU�)]������[��f��I�!�B~����\��k�?U���#R�����(�x����/3+f�J�%�g�kb��������M]���lu�Ge�h����	0�;�}�}�;��s����2���ƚiJnOJ�ef#�Yb�뎻���J��r+�"��թ�#�uj��i�G���>�l��	,.�.˻�,�T*�����Zo�����<h�d�)�q�������{�����&
'UG�'b���DC�'�^�Uū����UӌU⫌Uⸯ����{^+�YŜ_���mx�+�q�1j�j�/Lc���|0k�ń�#�dЛVqq���x�Y���\_��/��8���|��1��j�,��-\qȄPG�~���-B�ylG/(����+�"9Z�Fx!ylG/(f׊ی��{o�x�wnt�^��L������x^.<c���9����l~4!0~[!�d��?�������{�h�;3�dު4LU�Z�n��J�J�p�V���];�N��|�҉B'cj2sb��n@�����áa�k^l�|`B�������O�	�K�|��}��Z�������Ͼ��W~{�UU��{�"�Ǘ��z������������UUW���	�����UU^[�z"e��{ު��-��A"��s�뮺�y�yG4�Z���qƚi���J�jիV�JEC$�� 0�1V�9J������A�D���B1,RcڪK'f�g�T�I@H��\b��z�x X��i$n:H�EX�i<H��J��T��� ���#���>w̗s���w����0�X>��z`��2I䣪�w1:����M��z+nYe�Y�Sa�QDE�����68Ԫ�E�a`���o�'"1�Iވ�75W�P��B�v���ʟ�jQ⡵I�#&Q1`Qq�%ЯH�>��m��� {A\�4�ETn�\���'-���U)� ��:�I(}5$��12�h���Ti�,�נ�<Ye�]o�?&1eLz~٢��
��ܤ)�ٽ(��"$47���Ke���'C_����FR�dvvM�0h9��M�\��aa]�s�B�l�IJDZ�"�L�kV��2�ͭ�g��RZ�������w��[x�s��8_��@6�D"E#�����RBaC$G�B�S��hf!��PF%����Ӳ��"fzD߅��rE$$NְOu�@0�8R���9�I�Ƒ�q"9tP�:be �`���G��
�*�]�Jm�]m]�]���9�@>���#��XR��0����$�i���s�!A�N�<>)JR��<��rfpQER���J+�P���2И �W>I���P$I�>�OR�l�I-�ES96[�)
��;�t�(�(i�@6��"q��%�h����܅�.;l��$�yg���>��,�O'�@���:s��`z����+��;�qp��^��gQ�vP�YF6�4�,��,��,z���.\=�Ej�}2947>Y'c$Kl�|%��u/�M����D� �R"��1�8����C�E]e��Q�|0~B[tX��D�A�81-�56A�#�ɳe< �7r�T�m0��i�}.�H�������;]�Ҋv��C)�,���;$� zdv�Ne=y�,9�!D��ON�R��
E�xᶜF�)���c%�+�`I	���+zKL�$�G�� o�SX�1"� D�l.��P�Cy�Hhtq��<>䗍����4r��0��'W�!���6y���M%���(�Y0�����=�y�)�O����1�ϊR���ϲ�<GI����Ў�L8�'K�)�:y�[-jlfե�աf��ZЍ�ъ��]6�
�-�J,������q64r0-�2��%a�4�1�Am0�أ��:<a�O���'/�yp�ud��
F�c���t�pt�40�;���x�ߤ�p��m6JM�̳� �k\9�eU}0��
pSf�*�<u��S^e�K�f6��٦n��>��]>t�L@!(�"��ĭ�$ �Ca�JR���M��lvݕK9>�a�<�0��F�^�J�`�zi���������o�6�zp�N���(�Xm�7\�!R���\�%�|�U��z;�uo��M��o``��$%�i��+�	 Ɯ���H�s�=t�L����z�y=�q�thۊ�LV�����,����:��$hZ�jMK.CRJ�W�Z%|~�%��FPB�L�/�8���&�RˊD���=EEx49�s=��9�{eYQNlc[aD�&s���1jUT��*��/CvC)����9�]��`?ivq�47E���@�Ei��II(��tͥ9zlɜ�d�B��'��"S�������N�Nz]*�Ӣ:�ze�d,tɩ�Ʒ��z\k5we����N�vG0����{*L����<��&x�3H���C6���� ��=� �Nv�M�!Y�Q��M��q=oFR�#��h�j��VȴB���l����Ǝ�'�Dz"r(������Q裂#���b
��U�x��'�,�6����~W�����?8����_����&/��+�W�Uӌ�Y����U}Uz����:c����8�>c�q\m�WM����������]����?��;?G迍��,�DylQ��<����WA��(�o�]��>q�]��gck����g����k���4ӎ����Ux^��c����N&��D��|B%�L��x�\/��k�3Oξ�P��(V�鮃N���g�U�'�O���O&���bܕ1j ���O\� ���$F){D���t�ڍ����;J�ST�Pl*�4����ʻ�뼢o���o\tFQq�5W��\�,-i�j�.��M���
[t�����ܣj�j����<����L����ro�����Msx��̻��˗l��W���=p�N?^�ɊA(4��0�ue��%j�5��J4	X��UUyw�<z=��uU^]�x��W�캪��x��{��e�W����{ǽ�n]��y�g�{����ߗ�̻�qXi�+4�cc����޳[
�eJ;P��\j����mcmٵrQ�]l�L�j���+��b=�%k���W�sT�Tn�YaQ)(\ɣ^]�n	q^�4�n�
�h^�v,�X3SU�b�����l]n8f����]�V��f�����T���a�:̽���e˳SkE!54m�X&)�
��B,>�Om��鳄���Y�N��靆�%�uJh���LV]ɯZL��F	�"l��p�Yi� uʭ�R�G*�]vaZ��,hRRQI	j�vj�D����wE,5���o&�uK���f��W��ұ�]J`�k��c�Rh�͚�a��Պ֖%,�X�}���l�, ����I�- N����5%xj��o��$3y��4��O�92�9�
�2쫰-�ORm�� p(��%���,���F�,5���_�N��r*LkRpw��\�6`�q�����;��l�j0�j´��)�����<���EV̱dǢO�xR��s�T�B�緙�=��nI�פ��� a9��*P��)`a8a��4�=Ł�|���K���t�m�����~�h���,��z�l�l�s@C����*2�@=�+O^%�c���&I�D�.\)x7���9
t|"%d� @T�}7�1
��RM*n�O�}ې9��L7�4}�Z7�]�e�*�]�V*~7}�ɎI�q�Z{_��UVp�n]:EQz���HN��И���� B��x�Ƀm��i��uY��I�>25<��u�ڈB�D�)������ǿXGgJ�Ȟ�3��ReN>�dɨ�#G��Q<H�6Z�a#84�B��cǗ���X��m��;���`�~9N�>�4�X}N[Z����v�$��(ӷ�I��{	ħY�FOY�X�V��Ǧ��1�,��\�����?M苊m��Bٽ�����w�>��k~���M7|�ӧ��[< ��,R��Wb\�S������k�L�Sch
v�B�f1�.����f��իr��fش�R�m�3|��9ٮ0k%M%;����\]��ӗ,�.	<8�מ�&̛��	jsO���c%��#é�6�ZpT�5��R��������������hۄx��X�`d���(���W�<����|�G�L䞫M����q7���cSI�y8#�	��c� x���e��4�	��.Xq@���& }���W�)*��v�j�J�����EQN{���f�"�˴�8�ƽ��I�8�+I$���B�D�)�vRs����D�(N4�0�f��=2�9-#M��&�BC��c h��i8
?y��٥��X)k`ɒ�U$*���m���0����p��,��OM������H�8���I=杦h	D�-�8���,��NO#W����>iXV�c�>R|Y���nFr1V��|��P�%�+	P�t�2�@�˶5/�.DkI��RUT�Ü��;ɇy�h��8K�y��Cn�Qی]�|�0u��]�ru3�9��z��=܆c! [I �sI~1ܽ㍸���ɬ�}Ƹ�@�I��ӑ��o]��Yb@K,�?�:Y�kL���?�[-ٌED��R��f�N���x�̿rt�����AΗ���E��ٶmSQs^yM���)�S���oV�Gk��ɉ����Icy�1��,��V�+�(kr����O����(!��L���'�HM�:�諣*�ʠ@��O�f�cE��I���!��L��M�1�4!�:�>y&vBC��i��@������5n^سMi��[.c�/3H�<��7ӣI�+a�h�iL>t�+��Oʯ�wk���Y1;t�ʕY���8	����1�^S mcTjb�#
y�<��޳vkf���:�p�w���7�G�h���m� =L�0�-�6ÿpOϜ?E�����e&f������֭�O'ӏM���6�ںkJ|y�	 �ΔUJ(Ǟ�U�)�F����9�z�;g����b���į�ū����1W�<c�N1�W�m}Wk����8�+��⸻_���0�����Q�5��k����C����?���x�=g8�6�+kǌ�^+�2ڼZ�+ժ��ⴼW۷��=gC���v'ǌ�~=��><���9b�G�(�pj���yC^Z����:}G�68|L���,��?|(�òɱ�d6}�����.8�Wi�8ʼ+�p�q�↏��3�Z�W�).��n=?�'��Q��b� �D".`TOd�T��i�v���I7�M��=/�������im�d�:h�����ٕ:���V]Nu���z�1�\m(�6v�C�bcF��T]>����Ɯ�}�ךy~¸���.����C=����.����3�=�{r�����C=�G��ܻ�/?A{ޏ{׹w~^~�8����r����%)yy
*��N*���쌚U�d�S�].�!������\ː=H�Jє�&A餶Ҟ�;�L��q/�(Ճ��n�gX�xs@��&��
(�����o�@ӥ7� fm�bm=��a!6r#Ba�aafH±Zt�ӊ���]dn��_��	殍��k7<A�ׯ���KN$ΰ�:�n��|���ci#�.-f\g��;���u/hs��^C���)]��;�)��4 g���c�OOSN �)�x7! �=l�4(H��L�n���ɶ��I��G����:�.�֍:V�ӥV������J��ͨ��[B���bm�U�[>�~������o�
Ė3F9tX�8�Jq`2���[�"Z񮩘�k��u
-�R��d.�D��"��
��eh��4��`ɨI�1 .��	$ti穷�����N�<@��3\;X�P��0��*1`V��p���\}�y�v��)G
R3<�*2<�u�qI�5�Ky��Ox�A�ɂ�`�,�t��s�+`�tu-��P���߽���`��L�ݒ2h��USTV�'��8�S�(dΏb�Q���r�5FU�s�\��1dX�"���>��� �n����6���O`a'Y�,p��"շ}��s�txڰ�V�*�ډ�_��O�Z��-hK�^f�5`�dm�q����v\@��� e)+��Hm��aQ��ß��Vߝ��R��-�QF�ΌFF�!Ŀ4��i6�Ni�n'�OL�N�	hl1��pܲ�%�r���N	�5䜒�-CP��c����)�±ZmU��[&�w�ژ�%QF�"z�s�X�:��N���ɜ����r����Kļ�m5��ǩ`ZD��Y"h⪧}���*�����2��'�FTz̄�=��Lq�MYekh�5L �
�.���`ݪ�Ja��V��Z|��N�r[�șDC�� �����P��ɹͬ)L�<'�v�e�.騺��J�omͱ.�.�� �
���6�5сz.��YE��steHZ��v.��ˮ�֎�rW*����?e�s�|��ۓ�Ic�	�W�@�$&�kz��qI'������e�0֭����,�d��d���buɺ�S�QҘk$�Ck���}_p�;F�?~v1v����#r,b[��Q~�v�h�0�kU�'�^xxxڰ�Wn�Zx�����B�%�hEh�n젹���|7�U�e��j��u)���3�%]��0��4���'we�6�٤�À;�&�sr�|^%a{��Q,L��N��8w�Qn���X�� ��4��z݇�8���p色�Ā�O"Y�D���M��݉�XX�
6Ren�z����LV�@ӄ��L8GI�0�a�C@�Ͻ�-�֖�-'���y��C��e��4��E!\�x��l�Zk�^�b9v�mJM�`02��S�~���f���+�U�!���߅��T%Ⳅ�\���>jfHUz���� JyI�u�e����cP��j�U��&:ݶ��S��1�M
m����3g��4�����9�m;iّ4����ҝ&<�I%]h	t���&͸L�)����Y�������G���Z!?��G�~؉d�|"'�	��4����i�W�ڼ^��{��x�o/8��彫�j�j�W�����tU�Tz4����d����?�K��G�>�ǣ�	����>�#��+�G�J��/K�t�8�/�j��/3��~G�Q�pr�T�XyF.Q���O����x�������<?'�����68|LKƝ5��xW�U��z鞮���6�&�����'ֲ�'��!y#������8�
}9�VU�t<�P������W�@��*D\�J��c&/�A�J�۫�_i�qU!OE�YL�.ޘ���)`�AwIu*.�&.�r�eV��-٭����]s���է��&��y�z�V����^OLJ����}ӽݐ��V\��{vw����棷b�ul#o���Ewg�}�b޹���������>�Q�h���ɾcᷭB�a?>�Ͽ|���M5CǍ�+յ_�1���鏨�;�~�;]�]�/?A{ޏ{׹w~^��#�{��z�.����Dq�{��^�]�{ވ�=�z}�˿/{����O�w�w��z#R���A>0D����h�����J�n��7h[6ode���Z9��6%u���Ѡ�k+.��hW[�0�$��mp0�D�,n�Gke)��v,c�7U��LM�˚Xhkt��v�؁v^�4v͔�Ŗ�5��%�q���6�e�gL:0e�����I�mhh�e��v566�i��Z�v�Tm �R\�Rk������\�tf���:�����	���MiHK-ͷ*[��j�Hk����Z�Й�F;G�{��^z�i\C,x҆�j$�s�(nζm��4�׶%��j�z�cư�]��%9l+�hn(�����ёw����Cl����ɰ2�C�����8R�]���5``6ɺ��҅
b�5�O������<k�ti1�7�=Js �N�2Qd8\�[��F�(����Ě2`�/o�4b"��|kB=$m�&[8,��0	�L����˅Œ�vzw+�o�L'R<�W����aX�N�Vد�|{	�M��y�X|��,&
�l�a�ZؼK�.܁��>�J���8�C��f�@�{$��Y�������/.T9��F{�mO �F�4>�N�Lm$���R�᠂z �)Ȉ��V�S�Է�A��^���(���)����F���V<kXJSq��{��	:�%5���[�������<�]��J�)�fN4�9��^{Go�,�R�����+&�n3�G��c�Ҝ����p�S$fPUY,�؆�(�c[.�F��2w�_�Jn�-�7�<;g�=m(ˣd�.&��d��8zXm�C�qi�8Xq0�I��ç����Zz�5tVj����y'[�p�i52g�?��q�1]4�����a��Y�&�^fhM��f���Զ��{W���M����*Ĵ+6�������H�H�Kv�lP�S]n{k��7]�2�^���k������d��G(��+ta�h�+\�]7��Hj�tif�Xh0/]z}����7-����S�5G�XwHMT7O�����;�oc�}�ϫ℻XZM���m.a~��(���� \�L�2h�p�S�L1��U�M��~oN�Z���k��=�f})v�R�}L��d�/�lL�^�G���<xPq/E�����]V����`�e������+'$���L�\���w�V�#0�T�p6S��x-��ܧGa�W��t�X���zI����
I-�ՙ��N�<O�u˔�GpVp;H���L��g(4j�!�oC.�3�w��Ys3l������Av����|�=Gk�e����j1d.��)v��<O2�������������h�ou��Xt�L!�A~>�6�y�M�n��+�7�����^s/�KA�/�-�F;q�N���C�g�b'|�9�����l�S!*�A�'\�N�<KO(p�8��>6�'��9�΁����;2,�g�0�+�V6��>2�����~�]�2ԙ�i0��0\��<�L��6\8��h�F;�]6��iRf��4���r�hF��u��e�mҐċvr�[CZ��$�BH�]1��d/"��:�$WF΃D�i�R2;m�����~��&E;B����k��:�M��L��˫�q��И��K�����Ar��;�v�0�=)��s��KZV���s�q_)�c��~y����}��㇇m��+�V?;1�:ѕ��ǆ,�Ͳ��x���� �;���N�:<&��!�;�E?��%ep���y���LHCC�:����;il�&�T�c��;��Yeѳ(<B�=�+�W��~�FS�Q����[��!W�����ٶ;Ucv�\Tk��:!>��!>á�������Wn8Ӌ>]/k�1W�W��ūūŞ*���i8(�i	�/�C�O�h�C��lq\Y���^���2혮-_��KW�W�q]8Μc��b�G�(�pZ���y)r�W���^\���j<���0򆼡�˔-q�/2ޜgK�ұ�WW���������N�����;'õp�L/J�4�t�/ūÌqq��N߇��4����8��p�Y0�DO�n�&T�� (��1Tљu>q�M��#b	VVM�Q
����b���۽�M�s:�C�NEU��r��y-Բ��v��V�U2�TmݵD��svo�n�vgl�ٌT�M^��������Ϻ�r�{����O�w�w��z"4������.���DF�������_��荟{��z�s/��=������_��z1(K���*��f1�����q�Lx��Uaם��44��I�<*��~ d"��J
�(]]t?a�9	J[�"��dY8��ƃǵ\�ΌK4	m)��m80(3�!&L�n9��N+�&1�b�Uc�h!�fA-cXP;2���UG����񾪊�l��Yd�	w�˹q��Vⴥ�I��$���u,:�F>nadm����[W�N�Le������'��(�K}%H�7r2h�d:���\���s�	��N�!�'�8�_�~��t��r.�%�me�O .���D�h�ve�FU�B�mc�J�k�GF�Qafы4�$Ʈ�161�.��Lʼ�����o�V*�����!�\�3���`��l�[z�7�`8u�\�L�JL5 m*͜Ԓ[�4)ݥ�VI�%D�I$�2t}U|��S(��+%(�r�O�A>!� �3����.
]琞�Ͷ�W����������:�=��8����E&ir�I~n��h�X�p�Εww%�a��]�]��̟�TZ�\DI�shꈚ�jHBB�b�6�{6�<=4��1[Uc�Wg�:�w2V�dLcW����(�ܫ��>����r�.��9@ך���Ꮨ�K���t�$��{��ERx�����:��'��Q+����o~U٣T}���2��zCT4|S��WJ�U��]�4��?kl��������pC/��(ؕx"�~Q��"�+D�H��37<��oq��M��U}���xP�N���R`|(p���i��a��W�l����G�W�|��B&���U�vǍ��D����{I%�Ԓ˭��z�칕���+mJ�bT�)�qt�v�Ď�����A.�����Y��w:k-Ќ�318�8t���͂����VET���\"�(2�E���Ә��R��Q����=����|R�Z�o�j�F�1���!����T�\喘������DY�!�������]�V�4�)9j<O�m}��Ur��$:��zy��#���=L㤭ԗ+ioJ`pL��=�+�l�$��"XK�i���1��������~~2ZW�w$
�:�q<�iu۪(�,�ݿ����+�z�Ǌ�ͺ��Ԅj�k �Oui�f���|-2��k�&�=�T��˻���f�g����.��:���?d�2HØ<m�d��e�v��<ã�O2nP�ӓ��tX�,$���4�̚S��;k�U�2I��4��߻F��H|�i^*��Wo��|�_�+>��+@�I�0�E����܇N���Q�\ˍZ[L�J�F��Z�w�&a�(d�*Ijz��aSS���Y��]ʅ\�[t����ف鲫ڣT'�^���&
;>��F�>v'��O�Q�~Z���j��x��g��|q�]�����8�.�cn1�{0�*?
?
'¯��[^G�\$p�Y�t?��֏�~__1�qv�&���{|�9����t(�G�U�C�>4L>'ñ�5z�Tyy52�!��aK��1G��yj�����ɨ�(k�<�F��ǙoM8�/K�.+������'�d��t�>���qL>&���L�ӌ��L����qY��V�f9~o���L���1��5�\���{�E�Ր��ig�b��ݴb,D9�^�Z��Ǘ
o�$tOlN��UU�'g����ZM��J�'�u(�F]M�Nn}-�!�;�����L��TQ�Ԩ&�W��狫���}R���v[��6yD�u�Lӄ��:C��RP�݇�Yξ�ֶ�@��<yУv�G���z�}��)~��ϋwϣy_~��0�%Ad�����yo����/���b�{��z��/��=������_��z2=�{�UY~���Ed���������=��ꪬ�y{ǣP��	���D���R�]���-5���x�+�V����\͈O��G�mCm��-��m��mM��YE�KHn�#Bim1)�4�VZe��:��$ʖ��CPΫ�+)��Д6���1\�[�ic1]B[X���W8��M���OO.]e�I`�SQ)n�u�1�#6�d�Y�ڛY�[q^����Xf�뵶����.D�t�X��gp͙���l��x8���Ť+E�9�hǨ�Ͻ־&��)�e�鉤�vu���]!��ɔqEqu��-�%ִ���z۝6ec�u	vbhQ�]Zґ�Ht6�qv���W��l�ˍ3��u�!��[s�2b���CmF,%�tM#� ,)�#�f�bb0�Jt�lb�䛥�VE(�I�����,���Y(0�n�)҇�&$����e$i������zE%���G>��ry�.!�e�U��i�l4��zh�����d���C�G����q��7D�Pp���F�Һ��q�m֜�Y���!��޾}ָr��N!���͞UmQ���ʭ� ITϰ�,�}��!�64�PCb��<y�"�+�g(���iJ�_�X����z�Ld�[�H��\] r����.�p���V���U��MR���1�*��$���ǉ<t��bZi����$!	�}(�OK
=,���^'��7��Yzp5VC�@6 ��7��k��tL޷Ϡܶ���'O�����"���N&d/$Lk��9A�h8N��6�8���ѯ6�8�����޶y��2-m㧷��|5���	���B�{����5y��"w��������������酋�B����lWֺ���Tq&�V��KhKx�۸bY�c�J\�M�-\Y6��]{j�63\����ea�B�.���RXb��.0m����z~�"���A(�E���׹�Q6�r�V�a�Tp�~�WL�X�K�b�4�gP�Cz)�Ì9�1����[�bM�6�sv�%%��H}��Fڇw?3�q����!��=�
����^��9�8L�����-Y\�B�}�.[�4ȯGq��>��i���UB�w��I�ԍB?�DƑܻ�]��q)mL�0�;Ώ���I�q�YX�b�[+�??0|v�6!�!g5��3Hl<U�G��&�K�S�FL�#��1"��qH�m��$��d��W[�J��`a����֨�2�n��kTt���O�w�K����:hh�{B�dT]}�[,h�����pC�9�FW�E%���8ˇg��M�r��E}Z5Z;F�YepT���.�lwb��q��[��'�9�g=(7r=�I�I��=:�M0��l�b�F��]6��0ܶ��l�?F?n}���6�~S�>c���'�+"cr`�;"�\�]�}9W�ُ�˽nk���o/1�Udͤ��1�8yj���V�k�R�%�*"0�D��:�V6���"pJ�Yy��j���n�e�7��S���t:�W����C�h���T^W��漞��A��XuaDO}'���LK{dNIZ<nA�����ޝ٣Bh�|���+�e�K�K�}Ü!,���Y������R�Sl:QE��Ą�f.�r�.Ջ��Xi4Ĥˮ{��Z���x�t�i����pNfg�E��-��,�kD��ƥ�����7F���(�w�|�¬�U�L�Q��+_٢��Ӈ+��|�8p�q�m����6�k��mv�ⴭ�6lٷggn+�Ǌ��8�{���_����6l�j�Ͷ�6۶�6�ǯ[m_6��m:m��6��o�|���6��n�v�mb�lٳev�㧍�z۷��m�ئ�JSI�	��MB���;Y$����'Jq6�wRN�ҹ.�x*D�_D����PFv��y�֟Z�9�ӳ�w5P���GK�ܶo��]ڊ����.07#"�G��U\�M�7�S�ʇ�$�{�AN&���؋w/�r�3VM!�.AyK~��|ꪫ;���\{�����=����{��UUg����q�{ު���������UUY�/x=g��z����^�{$�/!!x�螈��Ǫ[�gy�;M::Ό�z���.��>U��yE��,����kJ�f�]���y�����09>�tp�8J�D��E�ܑY�y6@]0�h
pq=�a4��F �z@��>!���~J�V9�mk삛�4��z�<U}��N$������䇟~��� ɝ�idm$[H�Q���6�p��.ޥ�L��;��fN��3C�������*��a�q<r���׶��β<��ߞ>4�aҕ∝!�����l�fz�.w���m=��a��-�߹;O�{f�Ke��2���h��K���u"��ؗL�YT�W��v�T����S]�i��$uH��e8M�;����Ԑ�pa18v��h˭W	K�Z�,���E���	��q�AdJa���a�U$�DVFQ� ��U��\;�>�%u8���Jڪ�c�1�6���W*6�
ɜ?{�v�C��J�.����������L8M��!4��zg}"���Guũ!d�i�[��F�7���dQ����ꯞN��]�s�&Sq8�1��ydnz !����!��'��W�����W���_5���k�g�-+`��!��i��:�����z�ם�[�����n�%Qi�I�a8lɓw���@�Yۡ�~�7CF�.�Ӹ�G��W����GP��O����GKiZ�YQ��viy�;M87�*�U�uUM�2����h2���P�����p�
xMa6�si�J������Q�I�E�V�~2����B	����d%͗��;k�.�/7��"�S����D�����=��5�=o7J��L�\�����̸����6�R]Tv�v�(M��I�#.�JhԺ�h�H"I���j��d"6֓�l�-!��SҶ{����&�`d�:56�)��2�۷i��4jn�W]��ap�Op��X�;l��.�`���l�bą.i��Y_��0�a.	���{Ϝ^7um����p3���Ј�!�C؂�GW~33+c��L��Wk�*˻��Y�×����S������ӄو�2e��x	���H�].2��[*��'M��A�k����}��4ۣE�y�sq���z�ѥ+j��Ǆ!�t�}"�4֘t��������?L#�a�8�c�[e���C�_ۣ(h��HĘz�����q��y(�+-�*��8'�|��38�]ܪŜMrl;��C��+��q$��w���ޙ������&&�IV���T$�M���!N�_i1�kPb��WIF�eb+��U����.ѥ#w�:o)�au*V��s�����uu��Ǳ��y�:�aqf8O�ubWd��HL0�:L���|4V{8�OX�ӳf����n8x��:qӍ���m��oV͛6m�vvvvq��qƹo;qƞ��m�v�J��e6�m[m�ݶ������|�M<v��m�񷭶���6��;x��n�m�جlٳf�㷎�6��n�;i��b�lۥl����n��~}�[캹4�[�ob6�j �ZI�YgEཱ�Qg�8�]*ӥ�3�E�6>X+q�Q��zsװ�R;�)�h�W�c� wu}
��yD���S��*6[F�y���Np�%{Sn2cffj����]�]�s�ј�"�I$�_w+�B�{�}j�#&o�Uɽ�3�d�f�]��dL�x���e8QE�L"V�UT�%�M�fJ���lڹ^�朙�fE�]B�"�%TEnFT��rb�_��[ڪ������<����UUV{��Y�{ު���������UU^�/x=G��z����^�z�{��]u�\��r��R���1�0�ܲ}����jr�rڥ�l��t�(�PN!�m�SZ�1v�=D�lCT��'ט���i[j�-{�"u֓:���ZYn�+.�l�I5��3����4���[+WmF� 4��l党(�a`!nf���>>��z[���mJ�>2���e��-�8ⲋ�0@��4l�6��k,BZ�����-���ce���[X��B0%GL�Jٵژ�Jj�f4Ԏp٭I���s�Xk�����|w��&Y��%ױ��к�Ym>{�r#��7��/bitf&�n^��2"Ѣ�YX�i ��]a[��lc�9�o4�C!3�)e����,u$��d�����rUѵon"��n�V�d���m6/��]RV�Ѷ�R�-�ZZ%ц�$p��g~L�G�{Y���.���WN����U9a��x�J|3�$$<L'r�����c�B��^�Đ����&�.��	�wD�7G�k����T����Ҫ�ǌc�Ӭ*�S�WD%�����F;;@���)Ԍ�T���U������9�nX��f}�cn�4��[璷��FyО��\�t٪���x�3�4����KM�jW����1�m�l��]E��Q6��x����Q�a�WT��U�ɇ��u�+'^eXK�K��b���)-�%,b�e���u��u��O5��3U�X����]�M����溋cR;OUZR�U!����mɔ�,YPeǀ�y�Utv��J>Y�%_e�c����E�Ǔ��Si�$��N�Z1�v�����%�d��w�]Y��o�\M<KKL�ä��-�XA�dA4"'H|B����fU�޾6^��xE(������WP�-VJ�U
ck$��ox�,G%fv�n�
f0 Ѕ�P�ję]*�uc��u�,fj��0�j�,BRY�+h5d�����:q�\�&�މG֞oB�&'�$��IӀb5�q�]�UQR�-;�u�m���j1�,ښiZ#��$٬�m=�ǭa/KC����<�!�/N�7v��3׌�0=�4���K��B�&}4Y>�c/=$�%	>�m,��]Ylѣ&�]d��sʔ�T�ad�!�h�WP�t�A+J�ǌc�O���=y����|眎<�q�qU�舝!���_�Ԅ�U�z��F0���_V^�Qi9�����{���s�JK����-����+��@�KO��N꡺.�'�Ivܫ.���WB��O��He�7ԙ��qg�Ś�N0ҕ�ꪾa��Ϋ�P��ii��W����k��	��Y�����%���Yue�wwuw�I�2�o]�Y����=�vV�U?
sTp��OK%�th��%��5�u�\��k%��Fr�i6��ҕ�+j��1�jh�/|�6�W��Q���7M��nrЏ5�!QN2hZ�60Q:���	�.�V��c@�Ζ�S[mc�(q��Sj��2���+�iWU����/註,ҫ�Whh�U��܅��'�R�i��)ì0T���GNQ�����󇤨�E�8P�a��u����$��2IQť����hь$h��d�߼����0�g��=қUW�+�Uz��1���'�32�K�����8��F0ٞ�_XC	�vv��c�&�`�m�]$giٴÙ��<�����0�W�kp�J��]t}Yl#C��3�Ƿ\Q�v�TSϪ��k�<�O�VQ�8��ڶzl��>>+g�6�6�N�u��o[m�m�x�Jp�ÇWggggN���u���^4��6��m+g͔ٵm���m�m���z��m�m����m����|���6��o���m6�lV͝6lڼx�Ǎ�z��n�m�ح�6tٶն�v鯽w�=݃�{f��cfgg:و6�ݫ�v�".����&��GK�Շl��O�q���W0���%R+�ssg7'kTe�u[��7vI�+�U�4��:W�5�&��{JreQ:Tܵd���}�Kc����X�̸���\���4��̢*"]�8�"�>X�fydE�M�]Y�ѹY�.��O�w�UUO}��g��z������޳���UU^�A��Y�{ު��o�������UUW��yz���{�UU��^�iy^P��U�8�1��t�����Z`6�vEy��a�I�%��$su7E�]�]�v7ZQ�4��N��s����:Q�G�z��9�3\Q�Y��w����]}d�����t�;=+J����x�1��c�}�{j77���v��/Ԗ�(��/3.�&a��a/7�	%=_Uxaֿ~/�BHC	���<��lh��pўE�FӔn�H�Q�ǎWw\d�o�4t�|�������m�%L���"���Q2�cj��}z�C�Ʈ����fe4�+5��hy��1l��%��[���%�h�5�Fj��,9Vʂ�!�|�n�����Oh����
0�V�;-=3��d����|;r����>m�:4{=�GO��g^��P���B`ȑZ�)R+��p���TMQ�g|��#�!��lDM�؈�q��lɐ��@�a�d��'�5��G����m=}0f
��hh���'ke�d�H�Z��&�:д�[�BH,cч�.�/!�Ɇ����Uw�۴����GV�.�����a��c�Ux��"sd���3{Ӭy�cM�q�ÚUj�j�Q�hOҎ�ٞd��iK�VbMߘݷS|Ύp����a���ϵ�r�Z���ٮ*��գQ����G�����Q�7����Ј�!���cY���7(��u���~Ҝa�P��̞���Ѧ&-ʃB�(4�ʞ�����5_�}�Pؐ.���UaE�u]!{䓲U]�{m2�pp�It[�Ô�)�<;����wvZi����}0҂� ���'3�zU:&���f�X�x,ڒ�j��H��.}]�"ݻ���k-�/;��͹���f��@����a����bI�"��R�۽��0�����7gfֲ�IN��E�kK0�,#�%�6�M�FZ+�� ����2��#$-�ǈwܚ��\d�(�p�`t�|�e�"��$k���2B(�I�f�'G�'�ߐ��R @��"'~!g��n�ܚ�i��:��lõ��u�(����MER)���G.�y�T���х����]�:1Xŋd�(���.'���>�.=�j�7&���(�	�C�<ݞ>N�(�N���):��n�ʗuz�IL}OS��ߛ��4N�܌*�)<�q�9f쵑�VBtu��O0h�'k�v�Z�b�Y�R�,Q^[m�+瑭0��1⪺�7wR2�c1�+1W8�/��
.I �Quä.�he�<M>���2M��;:�G�`t�FXӔ[9���Mf�FȜm�&�O�rJ�^�#��yl��ۓN�F���J�x�֏����>Ԑa!O��I$�@b*�%�����?�p���$�s��[,���A]��R� �Hds?q�%�΋e�
"B��GX>��DR,����Y"�d)AH�H�Q��T�IbiQ1IARYRT�RP��BQd�EE�Ȋ)"�"�"(�
*H��(�B�(��Ib%�E�QbEBQH�Y�Qd%RJ��Ȋ*B����X�,L*\f`�F)E�(���Z(��kԢ��Z,QeQeXeHȢ�,Qh�E��QeQ�F
,��(�X��b�YF��i(�G�p`��Z*�(�EM`�3�J���5R2(��YE���,��(�E��jP���X��(��,Qe�T��,��Qe(��(�E���F�(��%��,��Qb�*FJ,�T�b��,��(��(�#��X��,Qe(��(�#%(��TQe(��(��YEYE�,Qb�(��YI,��(��QJ,����e$��(��QE�YE�(���DbQeX��,��,��RKQEX��,QEQb�)%J*QeQeQh�E(�I,��,Qb�YE��
,��$��(���E�*Qb�(����,��QE�,�b��R�D��� �bA�	$��0F�(��(��(�E�,Qe$��(���,Qb�(�EJIb�(�E�,Qb�X��,�,QR�E�X��)E�X�-Qh�QJ-
)-D�IJ���,��)(�b�KE�YD��E,��iT��D�E�U,R�R�R�,�K�X��Y(�R��K%,�)b�R�,R�b�(�JU,��K)E,�Y)b�b�JU,R�,R�E��)"�d��J��X���)TK�K%JX��U,R��J�U,R�*�)h�K�)K�X���K�KX�R�)d�ZY)b�)T�K�QE�b�)T�K%,R�,R��,�Y)b�)T���D�E��)b�JU,�X��%��%,R�,��E��*-E�	�K%)E,R�b�)d�U,���)aK)b�J,Q,�ZZYV*�X���U�J����R�H���X�U�b���R,�EUX�Ub��U��R��Ub�U��YVJ�R**��,U���U���UX�d���UU���V*�Y$�*H�T�"��b��REB�*J�*JH�T���dJEI�H�T�H��EI�H�T�H�e�0�QAH��E$R,��P��H�T%"�)FA�T�׺9������	Bh�<��ϔ� @�UBBDF0s�J�����_��Y����/��'��>���������~|�����c>������>;�e(Y?���>?byό��a��9�BC����Qg�Ο������>'��y��'O���'����y���������PP�C��EU��LB����|G����}�h��I��bP�/��?�o� ������HC�t}�"��p��*���'����BH�I{Z�T��B��p�1~J�'ޚ���))?�7��i�k�ַ�F�~A>����V|��Z�1���?��ӏ���LD 2D�IY�b!&TA�(z1ED�G0�B���+�3�N?�C���O�>$�?��,���T�)2��KEP%��!D ��2�g������0}b�������w�����D�A��xc���B��/���~��A�*���k@n����?�_�;?h����������a�;����G����h�?#��d?�L��������~���O�?_,�{?����UD������,��zW�����g��G���~� �)�}��UD�?�,W�?N���h��>���>i�	�ԚH	FP��E ˕��HBB~��IOՀ�D��U�
Jh���㦈�'c��ID?�пMhN]ꏽ����R��ƪ>�oh��l#$<�9$$�?GDg��C?ATO��̡��R~���P���C��~�������?��>��'I��O��B�����z3���D��~���G�����UTO� w�S�/�~�?0��&��2q�l����<���R|O�����'�x�~ZI � 0�㟰p`�Lb��t3u��~%�_��迏��|�2%��I��ἃ��;����i?��X���0�R}�>@���P�=�c��8���9OD�+��HV�`r)@��G����D����$�

LS��v@O�w�ht�S��A@>���Q�����������}���S�����H��߂o�����w$S�	X���