BZh91AY&SYXX�P_�`q���"� ����bG�>         �JE*������UJ�U(*T��*�J�@��RJU*$T�R�*�$�J*�%%AB�QT(���J�$��H���)
���RE	Q*�T
���ER(TQ)RB �%QA*��   �$���
�,�I!"�B!UFhIH�R�$�   ]
�R�J���UAR�$���Q@P��oy�U	A �  b��)�2h���F�m�km�Zj�5[U�����U*��ݲ(4�2���l�J�e����:P���K�T���'�  w6z�	 �x�ΪR�J���g(�AN�Ò�P%w%�-l��ڪ���t�:��[dX��U)EB�K�zE!]j��n�P��T���$�BE!*(��  ���
W�gHA;]��8�m�"��7�T��A���
z�Yӽy*�%J�z�J�[IK�+�x)=�^s�RH�����JU*��BJJ�QU	*<  �����н��K��AUE+ީyޣ��jc�8yUE)���=R���xoG�BS�W��l������%z{�/m�������B�����*�
RQ(T%H   �w�@TU�O�ʤ�A\z��R��M��E"T��yT�QE��uR�<���*���m{ޥB�ޤ���$x����*�d/:�"RR%R%@Px :  s޼�T%S���%*�R�z�v�e��zH�O{ҥ=5
oI�w��Z�V<��*�*��z�Ҵ� э8m���R�HHRP� JE%T�  ��B��J����	$��]���u��h�%�{4R�=L r��9�*�*�]�f@ju�*�7�Z	�H��(��UQUx  g.�"�hR�9&: �8t�t�tI�Vt㠡U���U��cN�*��N�P�9��٪����	%T�A�  68<E+P�u(Q[C����n�T���w  �)�T�F���L:$�7E�HV�vJPQ�h
�QQ���(-�  ����DWΨ���US��:R���� vV:�ju:��궱�������9w�����    T ���J�`�  L� )�IJ�@ h    T@��0L���I���Pi��H�"x ����0&M4�44��L�����OPh @ $����&�   �ώ��\wjy���w<�89睶������<�8�Nw1�7��ӛ� U��� �*�"�Z(��ڢ�*�������uO�Q U�~Y�1��EW��aS�Po/O��g��;��9���9��9��9�d�`�Nbc�9���Nd�N`�`�9��9��d�i��9��9��9��9���&N`�Nd�y��9��9����9��y��y����y��9��9��2faᓙ�d�`�Ng�9����9��9�`�N`�Ng�g�9��9��9��9��9��g�9��9��9��9��g�9���d�y��y��d�`�^`�d�`����9��9��9���`��`�`�d�N`�Nfn`�N`�a�N`�y��d�Na�fg�9��a�^d��y��T�9�Ne��9�dY�9���Q9�NaG��9�Nd9�fE9�`S�D�Q9�NdS��9�y���E9�NeS�D�P9�N`S��@dfP9�Ne�T�Q9�NeS��U9�beS��A9�NdS�T�9�Ne��	�NaS��E9�`S�P�Q9�aNd�Nd�P�9�Nd�D�D9�0��D�9�Nd��E9�dS� ̧2	��9�a�D�T9�NeC��E9��� y�Ne��y�Na�@�0)�D�A9�Na��9�NdS�sʆd�D�9�d��A9�d��ȦaS�D�9�NdS��y��A�9�Na�D�9�eG�S2/0��A�@y�`�Q�Dy��f�U�UG�̈s �eP9�C��
s�a@�Ey�`G�I�`�U�y�NeS��g�"�"<ȏ2#̈�<�̊�y�L�2���<�2#� ��2 s*��̠�(�(̩̠� <�/0����$�� �*��2#�(�<2̧2#0+�(�(<�2�̨�"�(L����
�(fE9�0 s!0+����(�<ȏ2��(�"��a2#� � ��/0�̠�'10s0�'2s'2s<��<�̼�̼���d�<��<��<����̜��<�̼��L�'2s0�'0�/2s<�2s2s0s/2s'0��0s/2s2s'2s$�0��̜�̜�̼�3̼�̼�̼��2s'0�'0�0�'3����<��<��<�10�'0�'0�2p��<�̼��<��L<��<�̧1�ė2�f� ̡�<ٞd���<�2s0s'0ss�0s'0s0s2s�y����̜��<�0s�`̜�̜���̜�'2s0s'2s3̜��'0s2Ā��<��|>?R��m�5�,�;|*�p����j˫�(FKR���;`5�^��h�y	Ӧ؈L���%�J�qP�&�̠U]ju�GWb����Ӱռ5n�<�Z�eh�&�ה
�r2+F{ck�;w`��(5*_ƢF����h���R��8v[�4�⽶�"�1(��Ҫ#�b��M�5�jd� �բSE�D�g08�`���EaP�j��DK��8�(���5���Wef��t�J��p�wV�d��6�]�����02���e��Ň.��S����e�W��H.c�d���^�i��7����,��D��M�0[*�c��$���Te����[���[wt���Fm��-�ȝ�	mݑ�d�U �lR�f��E<���a�Ҷ�y�6��Ne20�A� ����sc��AnR��:LE��i)�+n極�QDKаCY�����6X1��l�V��Q���(�334�Rzb�Q	m�P�h�/3u��q���.�5i�LPB�wJܛ�Ǖ��^%�hY�����(�h�P	��ذ]��7ne�Kd��˽ePz� ��x�4&J%`ZM̕�aؑ�+7c�0��#�6�`����kcHk�P��뻄��Q��,T�o�{2��,CC,�H�6����&���7@·�E�^�,�y"O6�jݗ�Hp�J��O�{"zcH��;e�p���@����X4�n�X�"��W���P�qߖ�.��t�ݡY��X�h��sg�Fv��.$ݩ�J��V(�4�پ�oR��ܩwY*�t���ork��j݋0,�f���Y��mn��iY�"��
��{FXhB�Π^�k�HZ�ǣ	���]�E�h$.:��{��R�N�P��b�th���/��H�� yj�Ԍ���cc �Yv�!Sh��IEE�.�
�r+m�N 0�/Y��!Nf0>s&��NQK���	ն����&���f�t"�����^�6�D�1��7.��,ƳIZ������3���� �VGb��J�iD%ޠ`j��`{�J�JZ#p1���8&�N���lұ{nV=+�L�L�`|+^�yWX���7R0M�ti ����͇l�3nM���FP�(�MD� ºA��V-Ru*̱����Y2�,�5TGI&  ��S%RgK�ܤ�sw*U�M��M �M���+V������И�6��o.;{-n���ҩ�0J���� b�Y��VMT���)S܎��5��֥��X���n:e�Z.�b�^�m;�l	gWȱGnQn�u%i�&���,�1c���G�%�0�Iqct�0��L՜J�zv� A����M��$�Ì��6�ⵡ�28rz�5YBn]K�R��GE=�@emkcX&�U.z)d��ɶ^)rZ���
�L� �m��1�����[��5�c;S�I�j�uf%Roce7�1��l�� ���6Sڵ*�I����)d"�L����X��YF���Up�tr��lDyI�7X�]�Ł��/ ��uliI�>�oV�)�[��2�-[�*ܹ�9�(ް)�w���3N�@¹pE�7,��$˚��l����V��`��f�F£@Q� ���[;-E�{t���&���r��4�r���/Pj��p��"�V�ͬ!��7����:)9L䡗W��k���U��x���^�5�H\��B�e�X݄�}�XkfQ��Nk���o�8	�Mm�7%=��wy!ě�� ���9H`m�̊�u��V\�z� U�B����X��3d�,�B�.�T��fJ��g��r[Y��z���
d�[*�h�xaR��+Yl�:�K@Q�Kk@��5l�����aw��I@�̴��'��a�%KX	[�#;jՒ��B�e��u�"SpIz��3d�!�8�&�Ɖ�R�r��y�wc�9��s9�)��]	H��� lk�3J�:壒�
��-��z�ٳh�&n�H����M�t�ǅ���#�ł3X�1rȆAU�	B�B!=�b�(Lg��r��#���!�+Ej����k��*1��W)��wz�`�S��-��u�"�'֞'WKF+Ci?�M��n��56���L�H%G �ض�@$oI:�[z��dP��Ƒ$�[����s	�he��$v��ԭv��o](�SMռʙu����kf���SI���n�Od��b��CV��ʱg�bRtD&�VC8����pF��L��Yh��M�EC&7KQřACu2��M�t�ͱ�mҢR�n,�H6��L��f<�be�D6� �ő���7[!�kF�1a��h�4�G��Ŵ�/RZ�V^S	�6�]�-*(G���%�	��pn0�[�Tq{u��(Zj9��M��e��Z#�������Y0\De��a]$͡B�e


h���7��E l�5. j�"�\��H�{;3-g%KilÏc=�ZZ��5,q�nLF���V��6�ڌ�+����SI���P�R�����2K�0� 9�[�1ݭdv��§��QR��Z:�	CH�����l�X˕S#M���8�P�M��v!�b���Aب�:p�O
Y�!cl��D⼺7y��B�hYTCYqV�i�<��S5P�E+��Γh%�[������۹�49n�+h��6���� �M�Y-1l��c�T@�6�����P1S2��T@��Q�I5,ͣ5B.��f��k6��r�V�vr�B��H��ʡ�JJ��t��({L��]�M!!H<,x��+3e��l��1�%M�y�bz��l!��;P�FVYKSL�7i�U܆�P�&e�e���`�Ng�w�	;��3Ul�<��ZTX�ݳ�)�d�1�����mi�"��=
��T�ô�z��ax�A֛ɾ�j=�m��@\�$=RP� �U3JG$ciZ�#U�`)��L��K�;P�L�5��Ŧ�LO���q5��P�,��e��U�ӱowi憵����?VA��Y����]���ͨ5�YP��z��
V�$��u�oT��6�č�x�^�ŒkVee\����m��Ej;��בU)-�q!w���	Y�ۣ[W�S��/!Y�XFXj����33Vh̡@,�-�w��aPt�o�h�^i�_lEKJ�I���t��k��ܥ�X���1Y�C>���F�R%�r�1ԕ�Y� A����TiS��7~O+!�mk:�S[����ފ�5��[���'skt,Y���f#!��B۸�U��wHT��EW��4�
���\��@ham& e]]h�
�H�ö��6�&6��Y�PYF�1�Xl���r�GQC
Hcsc@��e,Y��jŇhk%MМ�b;Z�R��ӊJf���1�3Rm<�+3�ᲯGv4��jSWR^f64�(ïl�3r��+�详��	&*���0�Gr�љ���E*I��Ÿ��+4��z�էq�z�M��!#h��v�6[%��̠l�'J��©G��2����+-�Um�	��iEw5խ�W����m��!ۭ�x��+p�.�6p�a��N�<Z&/.����(d�L��1�_S�F�l��v�r���Ҷ�'r�FP�4Vꙵ�R	����:B*�V�d�٘w]*x)T�Ecm�Y[ �ēt꫘�
���C)f�^�.� 	�{a��X^h�5PSl��{)i服���mVL�$�[�� U�XV�Q	���Mc�EP5����C3!��;bf4�{��V�bK؍Ի��g(G�]o�6M�aeXZ�.�wu�5�̣�(�V�o.Uز�&��#T����ۃa��ݐm�v�g���V(�r��$�c��4Pvu�[.�o2�Ie=�Z5G�[�����Ŋ'��̙&VT�,�<�+1j[���ʨ55��9 �"�ν��´�9xSe�˻��Mqc^%^a��*��]�:	�r��i�D��d41-�ͽ��K-Y�jem�f׭РH+둊��lTP����2*V�d�{y4��p�ܦ��SY��j��6�n����t�"�D��oh� i�*���*aj�5x*X#�Z�n������m�ze���zB̹�r��b	b�w�eJ�<�y�k��<�%J�zcHԵr9%�ܸ,M2�(�+]e�B[j�@��69A���X�:�$kv@�N��QQ�y���hM��M�y�+ ���-Z$])d��*ʕ�� �3SɆR�RhT��l���6�_�����@9N� C���;�%��ò���7CS�
$���&��\�bQV��41�8���CT`X��id�{{Smm9x���]j�˔�V���G��V�U��F�,ɖ5�/e��E��zliR�{�eQ�i�Tl�ɮ����q�m����O�[�v
U#ŗHEoV��H:�C���c�2�t�m���
�(��e�l׫i�l�qV��II��U��� �D����Ҫj,���
o�n�؃k�b��MTh9�q)8n��p�ׄQ�1e[YT� 걿Sݛzt�D��2+�(6��o2R��wtJAܔ߭64I���5"�1�����է*�޹3E]����*�m1b�h�%�;mHL���kJ�
d�Xv킠��r$�$�7dr�^v�^��˭�ZU�V݉"eY��B��!��Tx�)�AAV�W7@ɚV%杤ءŭA.%K�#�r����Y��t2ȫˠٮ�Jb��F*Ӷ#N�V1cR��賴��%W���Y��a��m�޺aLIޘ������&�n����
�U�)��#yzM�7�U޺zK�������IT��s[�R���Y#]��ť���ynX7xۉ){��E-J�C$�����B��k�-�u�t�+P]P��h^e ��hMTc�e�0�Y�װ�C!D��ta�zһ{�dӏij�J�r�΃�*�MB��.�\���z��O��zwm��h�ҵ,(�m\������� (B�&����<�ƚ˻�b�tm���V��Qۓ��Q���N��OoXr@`�;��vU��R5b��%���!R>{pRguxn[I�Zɫӑ,��w2Q:�Bn"�輳R����{�r�dO
� ����"�Q�x�J��!6k���@�h�b��F�VWr0T��|+>�� �jQ�d��,�	��b��\��	�w��sq�Ɯnm��ӻTM��c�-�݀X����ژCݸ�e쎀��!�VV�΄��Y�rV�k8�/h���o�JVS�#4��`���6�`U�6�<Θj�aC�����Z%:ۺ ��՗2[m<�K�iY_]�ڼ���ˤ�R;�ܘ2\���65�H×���$���e1aQW�J`D�z�Hl���kX�7��,��j�]K�	�,q�j7�yP���]Eq��6k�Ϊ�R5LS[u���T�S�W41�㕛�2NM�o�j$��h����"M=n=�㢌v�Ƒ�K�_eò�85m<��o$�̽$�oM�zs���_�hm)�:�"�P����e'�3n���*:/\��+#���U�d+��^ʚ���\D@R#�N��壇(�)
�7�-V'bŧ!�J��������iGE3{��m[���U�6(���m�ICm�F0piV�軥Y'�Xh�h����cR;Ch)�Jv�4�c���2m�.��,Ruf�miWH2#�Y(���f�.�h[n��w��/DA;�v���l�l��Tx��Ӗ�n�������yIH��⳶ݍ���R��Hn����%ͼ�t�aG�*��rRڔ���*��S7B�,�QçPUe�����������x�Zv�dމ"�T��'+r� �S�
m˛R�N���w��wps�n�ɐ�P�`�*؛��^Ze̅�4�&��s	Jv�*؍-���N,�(XORa�u�-��t-t��sP�w��X�-=�G)��%<�V��6��6ȐF4��U�o]2�P;++0�O�@�G$ͫ:��X�Y5	PV��β>�u�CnX�#>�\)AwWB� (��Y��G
/i�uϷ���	q�baT@��s|�"��N%���&��\��,Z�*�H�C�¨�ǝ�P,�Dȴ�ư�p��V�u��<�����s�a�E}g�Ӡ�̏L�p���f�D<�(Q��.Ch!��Ը��T$WGljd�46�%�nm�|��I9v��A��J1�j���t�3�Kg~�Qj��ԩ�x���v)��T\7���fPBT��ݬE�S�c��:�G)��r�m�G�T�0���a�V�u���ʛ�cb�^��j�
����㴔�Vŷ}	7��H�d�j��3p���rF�5��E���u#�[ʙ�L`��4���o5�i;(>�݋yC���n�k*�b��0Mu׶/�a�k���I��7y|m�,��mQ�V3%�K���P�zy��fq���N���(��E��;p�ٵ��⑵�L��lR�7ZʧlVGrJ��at7�Yj� �4Vc�C�Pm�˭��� K�M�e�p��[D���hj�gƓS4�BGm�����j:�lɳ�v�+/�q������G��ݪx�3��GP�(Sx�叇]QkxwG@0���F�@JƓaBT.�\��m��d{�6�
�Ln�C]̻*�7M+��F��M�Fg"@Ż�g��X�Z�u.")`�z� <�%*r���=ٞbgv|pBi3/
XT�"3f1����R6�kr�B��{�4$*�V�C1��.m�u�HoT����#��ͫ��:e��x��a��cI�M_Ɠd���[X�
öm܆2�%2��&�S?}#��~��z|���hXI/6� �s�-��� h��Т.���i��
Νs�������O�:�c� �_��]��$7w�f_��ο��g�����V�W_���7s2�ֽ电���v��rVG;��7;�`���;2��u��vTvj-���-������Oh���L�̦u3�oe��l����q��`�{t9��Y�����gi6�q=�ՇdĂ��Ek�v�v����ޙ�]�$��2ܙ}E�5�J��$��U�Sf��!aZ�Mwj��XY�+��m�P� 4��]K1��IG�����3�@#r:۫;{�5��u�
�bj�`zujt�y�s�2��N�7��E�B�A�;�X�aa��M^U�^vA.����[,��$�k���*�ʻೝCԵ.���\n�T�������!�����s�+3�@�u��W�Z�k�*ke5��]��m��p
`���Xܗ�X��g�V�p&�i��8�X���ƌf���:��՛ɚ4�>�+��Z5���xo]�Ls�}��"�3+��{��]����l�	�{mg���Ly��E�A�
<Ww�V�w]G���5��[0-��m�V�7���30d�to��wǣ�TUu�KӸݾ�;��R�2Pi�M^�lmۺ�BXZ���Wr-�S��Ӯ�v9g����3�;���N[H�d���ɭ�Co�WJ�o�l�l������ˋY�id���;�5qE�g���Wev
"�ē���.�SL�uչύl1Q;q�fR�=����?+d�t����CwwS�*4��5l^��s2�]�B���.c��9j,��;[�Y��kD�ݾ%A/x��j7J&��a�������|zt�V��7}ט	���[�h�z��n����"�i�B�n����'.JQ���cb���{�7;!�����Ǽ��]NΙ1�9��V*��\�$�!��t��u����hyo{*�=�B�;$��R���o�{^+�R����cc�53i�+�������WH�6@]� ���G`̝�ԽO�����;�Ěͥ2��m;8�&�eꝀ\��x�}d�:�];�HA�ENE3~�cil�tCw+-�y8eۙڥHRQ���V�B1.�"�OwBU�ͧ�N�u#��Uv��v��zqXx��ë�$k�$;t�։�bݺZ:UF���[�%+RS�H�����$�P1�{&)i���A��8lG�c^�֖��:��9EM�:|<s.�Tr�WR6�9��WX|U�;�Ԛ	ބ��ث��F���['�
�[�)weK����[��i�I�<��v.�ˬֺ�ꘞ��\467���V��"VEDu�S���oY��/���-P��zڵ�&�I۟��&�<��I�������6*�;�Y��-�[Go�8�2�&�.����[�v'���h@�� ���X��\c��m��l��=�+%�E�-i�;*a�a��Y8mb��}��h.�X���rҬ-�)83[x�4:�9��Kr����5�C�86��-k6�����̤�1���0r��{mw�6>�u���OJA�ڵ�r/]������KM��N�e�Ge���u�ܳ�'�Ze_�m�z޹S�����ɴ׼jR��-$F��Gf���ј메���)���]�9z(D�<O�y9_�����Qv��m�P��|���-�����J|uCn Nv A�.�]|���e����B�����wAs��-+���:^@�&��[��v��%��!)��S�"�����'��s���� ��2�vGm�X��tR�U[���oS��J�����;A�R%���HV���zpd�_|>��C����d�\�y7��nTН���Pk���P�	c9:U��0����(c��N��EA��#\b�T��3���=L���]f�ڽ�w�ri@�w8e���ikL�-�ߧ�O������f�e���X��c+�U��Bĝ�)j)�4��5D��V�R��zB����pr�9���.9P���:�ͅ���h�:�n����b}�f��cdM]4��c<���m�s�uu%�z�n��ۄ#�Ӊ��A�����yae޼1o6���K������g�����+�)�O #��߻�G���az7T�$�S4_M��F���`�\����f@X��(휂�*�@��BV�.]�7k@e]�W�������E�}/`�7퓭N�^9r����dZ�2hc���T��Jz;�KU�s\�u�ܭ�
��m�ګee�ܚ	֘t��J�	�8��4={ E��ɑvW9^c�6�b����v����&�����R����i�\i^^���j�.�Ü���@�����_Au�1��N��r�Y09LG���%b�M�T�MR�y-���6��ʌgNA�n��gn�Z��!mX�ÝX3vZ��ziO)�Ǳ$�fJŴ�m��x0�V�|��S^�M�Ɵ�Y���s�3T�w\@���
�ȫ�],��m�I, f*��W Dh�n�s�����N�;�S�׺��A�Y3 ���u�a'�sk�%0>R��cf��n���㚩=�hV��:*݌����([�繥۷Øs{�W��]qL��Q�eg�d|�Mc�6p���|*R�a�q�΅o{iK��9K\.�]A�ڰ�&�����jLm�l ��gY'DC]������Y�:U�+r�6kH�����.�O�/���w[�#��_Q;4����tP<�G��0»���{a<i[ڗ�Y4X�k ̚�"̺��v��%e�̺�����>}�r���Žw5�+E�ԏBR��v`z��̊�T�*gwl�c��X����r��$]� H�wn��"�lݝ���_E@���f�u���
���U-�X%��nL�2,�(�\���T�&7�RyB�9#*QٝF���D��]BVgf��3�X�[�c�ib�k�q�L�;4t
�8�nc�9�x�ڛN��d���JX�������7<V��oڹ�u�Tj��Y[|��J�N��ҵ��u^��A�+:��<���\�9 ��zh�>S�3�:�L�}@��O��`�ڦ�f����Xb�'!�ӪB�,>�q�qO��g Z�J���F���op��b��eu��MSt���p�Ϸ�_t�v/�hc��JG�Wю�	�H�� RC(Pۼ�#�l�VԾ����:�ɐ%��s��l�ҕbO.��j�Q�齶R[��'L��b����xn��4�[�׿-8/B�(`�	�g{M�OY�%��(����w1WY���]s��9�����4�����N��3u�5�ً�o��Ļ���{fyf	�Li��'r�;�fA���ɂ�����oX
�w��"]�evƩ�{v�ĭ%Vt�}{j���C6�'�W�\��"P�h���\ୠ�R��4�Ќ�1�[xjX���]�*���^�S�`��͑ϯn/��P�:��V�Ý��c���1�1wt=}<{ul;��V�J�Nr�I���Lv���u��#���jc$��r��,w0ӭ$����]'�7^Н�q4�"��C��v�e��G1�E�-b�
�vPx^3��Q1�U�|D.�
����EA�uƫ��6,��(�o���ǫH�^'�X�������������V]�h�A�u�+��*�!�u��uQu$�-�: =��>/����x�qcX�/��V6� t�����79�nP4#��sWM.�=�Mb�ިR��V���lڗ0F	�3�C|�f���wFr�wXC<#��A�T�u7k�w�Fq�#��uN.�쀅��d
Ńݵy󛣖b�M�J:��-���B;���x��0\�hsO,d.���ꔹPd.��@S����.���z���A�c�Mr̙[s�\��h��<�h�{\����B[��Q���j��5ґ��ՠ�JG�����홺��N;����0٤#�9܌9-���u5�s��X�$�P���_2�v����$8�A�z���ZL���um�t�4��U�0ɾ��?r �t�+3繉�QWRw��eeB�K?z��|w�G���5KS���4�Y8�S.��w�X������ڮDPwI;5oN��/6�#��z��ރ�=�cR��mA��"ioz#])G*�:s�Y�S�z�ح���
�Эa��m]�qX���w�X�d�)��1��t/���-4ۆ�,���lʊ�1ֱ�m�j7z���Y����֩��"��J�z�	�Ao���첥٩{ڰkEu`��a%��1�5���PǿFZ�9�F9�[c��t��3[g����|�u�9 ���;f���opb�M�L[$0���9�p��.��j,@�B�F�1/v�w���ʏ�{uK3;*bX�V�*A���m��l�(�M��:Tyա��}�NY]�eZ�'��y�a=��{�I�v�r��;Y���u�K���K{�,tl��XZ�:�%2]�e�G�:�݋{]]>�qb��1�g;;�	�g5�iV�)�W�z��w�h@����fc+M�.�M�F�Y��������um>��W):MH�Yb��\�U��t�=�<��FV�Ov�T��/���7 #�q� �u�U��:U%r>�~��vg"��M�+]� �mw[>x�/7Z���![ �\35R��J˷}�V-�݌��$j�H��a'u���;t�ۇ2�� ��ZM����]�٦%��*Ms�R����|J�y�Z�f�[��B��7�k0_ :�j�9��jU��X���%��(��G�;�X�;�#�������T�ʓ3=|�Kz{rM����L��й^��C˳2c+yR�{��*�)M�j��"�qDҺT՛�uC�M�����nU[�3xz��
���Ѽ�@�S�_J`M:��'q�04�yW��9�ݝR��w�g�K/еƱ�v�:��ytcv�ՂS�W�rED���݉��.��b;���p���ѿC"ۃ��,h��a����ܨ!RIR��ib�Z��d�f+K
?9p�{VfVc����+�$-�]�D���Z-��G�M�B��n{�̸�wu�4��v���@of�b�(dj��8�Y��R)�y�Ec��Pt#�T���3�.��<�@��Q��1Y�����{��(ʱN%r��ͷ�gaW�a���j���j�]!5#��F·S�5ۏ��D�k}��m�ơ�駘��꾬QZ�@��K'���yh��>
`�X��ՍR/k�3�> F^�d3 췰�]z�[�ʜ6eK��9p�u/��ih�&���Q�Au�|J�սeå>���(�Ƅ1\�"�y��^�-Wx핢�tn��r:Vs��SeA��F��H3gW`�U���ot�/"���+T�n�,v��1� e�Wv��;�cs�;[�fe�6��6Mwn����++�`瘢oM�͗=lj��վh�i�>q���j. PDt��u�}/�P��h+���i�b�������ZŔ�T����KD�i���"q�ⲵbi���]Gkj@sL�G�i�kҘf���D�Y��֩��62��wt�a���x)T�%�gHG�w�b�h�d��фջ���@m]!GK�s�.t�q�{�G��f-5�I��p�gt�;�[����5�(ևA��k~E�X���7.:|w�|������jmo[|')R�]k\z���i�2�b<|�+�����ƌ�t�8
R������L��U=�V<�î��B�<n�H*���W�[n��\
�]�����|y �RPÔJ�p���ۙ���33C��G�Ǵ��F����K�h{���5�"hv�m�[�Y���H{/V������L��о�n��OUn;��4������/1��m7y�YQ��yW\�⳪����q*T�s�j�8�p�b�+�e~�|z�R-dz��p��SC�':�nb����s�Y�V�;�)��J������!���t�t༵�=Ev��L2ٳ\���0ӛ&{���N[��Zq.[/�G�W�u־�Ƥ4�T�W]v9Y.����� ��4���o�}�o�`�X����W-� nݩ�Ѭw�M���P�Պ�Z���Ӏ��b=�{ǲ�
�B��c�;K�wC�\�u�O��k>��KZ7���鋮�;�G��oKQO�V�嘷�<Ω�)ʴ&3:�oNN�~�P��������z��^=�i������7�x"8�ueXUA���Z��H1���"<<#H�!Y6 �<a�	W� t�%S��ѐ�
G�i�*1E��f2!%F�:�j��-Ie/-��ax�������$鄛E��Z,&��S�1�X!+A����"C� �&GcB�m��@T��wL)(������d�TA�r��-��a�݂���MYE�q�ˋ��0K�[���ô*,E0hP	��,P>(Q5MM�@�Ɵ#,rV*$,��'�`J�:	4y&�AA ��`���O�J��T�`HP�j�ґ��a�a�n�:M J�H>�wXN�X�y��1���
TX$���c�PeQ.�����`��	F)#���mG=*G��.�-
(�Q/R& t�	QD����f[�L
@�L�6��j�(�!)"��.�B�b�N�I�){ʯ+Xh4]�s�받��A��%ݔ�(��j�D�*e�1Q�-5T�ʇ�0h���T(�Kŀk
��R�eQm"����I� %$�f���C�Q��(��R�0)а�RH�m8��TD|���ݨ�"�uut����&DD~��������Lu�\�juclgn6
����s���C}D���3Ty���"cX�"�v��\���ѵ/�*�s9ˁ�Q����GgPC6�l�uԋ��vUտ\*��:��@��]�U�t�V�&���=j�u�b�g��)`ͫ�D�XR�q���L����4eKW,i��.�ĸ�̴e�?g-1�A�^uH@զc��qd���X���+��.��Ai���7b����૪u`R�N #m�r���m�<_
�7XI�8�YL�lɫ
e��*ܺ��|�JT∫�ݥ�>��0^5ǌmQ�g,��4�n,wyȌ�[Y�9u�ԅ����@�}6�u.2��w���q�[�cf���FV�&j���Ur$N��bН@�0e��c,����RJ��Xe�vp�X
�MCz�C�]=~\3`�8kEz�]h.��S�b)r���	�'&no 3�)�-��*��4Fdy��[U)`�}�2�U�|�!���E��Ą"l�F���o+[�ׄ��Y�`<"�2ښKnRc���
T$��#�J��쇜�-����p(��N-�B����⮷����\:���8��5WS˽�ɭc���ھ�ĺ�m ��=f�ݵ�I	��%��"���5����s��	��u��J�.l��3U�^�O_�����:333�333��ftfffwfg,�����ᙙ�������333�3:333;33:�33�33;33:3333ÆfgFffgq�ffgfg,�Y������ffg�����///,���Ό�噙�坝���^]�fow����{=��gs��0̈́�	ZG��nҀ�H��WVo=��^l$sG�\��6�XR7���n�{p�:i# �5m�Tgu]��R�w9�R�7����ǟ�Mȅ_R�՜�Jՙ������`t:'�ю7��y��T�K.Tq6�V��t 7���{9�c��ۡ6�������%�tz24(����ٷY2f)|7#��M��UK��Q^��IΡ�)��ӭ��w{�+b�K2��k7�HoA�.�'�A\�'m� �*+9K$o]Y�,�;)j����]��w�\4
v�Y�}H�p�ٰ8I�ݏ8�4Л�^լJ�o`���7>��e��'�g�I�|{q��������
�&���n>��{�v�D�g+/�̐r�BM�-GF��4:R]���,*�8!��% X	�Ø,7*VwKCk-��l�K���j��Z�mw{�1���EÂ[���2�Ê�b�t�5ʊ��vZ�ܾ4R�6�\�ysnP9|�U�!TQf�C�ZH��:̸_uđ����{5���H�..
�P+og:��`��[���[�26|a3�#M\]\�QNn�YW��n�]ҷ��^�R�u��bVEJ�'a� �lv9�h=����F��ΐ�0ĭ�}��8vvm+�"S�LW��������}3�����Y���ݙ���ՙ�����ՙ��;0�����33333������������33;33:��������38fffffp���������Y������������3�33�ffufffvvvvvwwfg,���}�w���}��i��d�J�A�*םn�D��+V,�k�_b_q]�[K�-��B,}e�w�y�ih�r��(ju)f�ꩲ�$�&㱩�{OjΤ/A����E3���;�u5��G#O��3��E���˪̸����N���;z����s�eJeP�tK]uo�����x��)^��K]��RӼ9�r����oE�-���c7P���7nnۍ�f�y�u��銼N�!��w5W�̛NY9�M_8�#e��Q[Ozt��A�p��՝ʷm�Ӯ��	�K�=�M:��u�n�-�G:Z[� 1��s��}���4_�s�5�@[�"M⫮\�}���#���X"K��gC4+!Ĉk5Au(ѳ��xq%)���l��#��EU����[Y��g2#+Zō�
�Xu��w�պ��0�=�;��̠u'R�ģz��t��5`r�t7��t��Ee�r6�5{�f���\�?_hŕ��r���Ol+�;Aƫ���ѥv2�7�N�0m��	�����Cw6$V�wC5�[�	}�Yʹ6o5��2[��\���wnj�-.c�L�j�C�Sju,8������R�t�72�]�s�N�p�[�����<�A�g��F���U�6(� �P�2Μ�,�U�&�<r��b���%����p�j���K����y����33�3�fffg������ffffxfr��������3�33�33:�33�39fffg�fr����3333<3�:38uffffg33�333������Y��՞^^]^^^^^]Y��نfffwfvvvuyvg�wV�{����Ow����gW^��y�S@HQ*V\��O�!@��ڕ�õ��vs�4�Z�p��G%wn�w�bƵc.�g�1j�X���8^;PT�gw��:���CM^�[��R�Aqt�*�:��lK�lu�)XX�S7�+-퐦�˃Cp���ve��d�-��Ċ�]֦S]���T]�[���Y�c��*��cJ�L#t-�۸*���.�ަ�k��������g��ɠn����k��u�ŻR=����KuN�B*υ��`@0���Xy�=��y��y�]gA�+K�mi;U�5b�߰�w����e����	5UB���3�������T�GS]'ɸ��V�&�B_[+�ٻϤ���&F�7��ר��4�B�'2.\�@��HN�U��}I�ᎂд�3l(���{��L.#4z�£��� z��omRj�?+�W�JXQ@>��V�H�ڙY�����KmA�u�^_6뎾�W��b�q;M^��{*P��GUT�F.j�ܾF����i�N��|~���%�}J��7}������ ���=���&��б��.��e^d�X��Al������o��\�r�a��A�L��U�9��R����M3�<!V^�.�������)�O-W�w.+�Z���_i�������C\p�������zm.�Y��0rF@;5+9��y�X]���)Z�l��D�j�V[�Ԝ�����7����Phl�g%l�J���Z:.u��w)[��f�9�u"�]9�ۮ�UOhڥp��(�-�t)��YZ�:�a�=ɲ���q^S��5��ՠm��|��a���5T��7M��l鰽1�b{V���.�Nmz�ٷQ���h��B���f�M�)Cxn̰�w��qe��5E�L����t&��M�\;W^ݵD;�N���<J�o�9=]���G%p��wޮ+*]�}�"&#���C�s�����C�&3z�6]l����յ���Fյ�И�7��o�����
ًۼ\C��cᗆ+��=�en��҈YꡖT�y�_W��+v��ۉ]+7�Vѯ�F��,�̀?N�tNI��5���`������\.R����&�A<�i�NY�Ǹ`�c�\���w�nt7Yl�6f<~��8��9(����1i;^VF��>u݌�cq����Ȫ�X�2�v���,�/�r���Ct}J�u�+Uí�.�״�V+xJˑeS}Bnj�����@��*�+	ndd�`�Y2�U[J k_��e�G%J��k� 8J,;�刬��ݍ-K��L����������x�f�Y�"D��
���bOg�^QW ޽U9���Sv4�hR3^T��(��=ڪa�͕�6�V�9�R��`���
�R��qO�����,9F�kΨ���.��_�J���M�*��)�a�w��S�1yBI`�C��ej�a+A�;ӆ�׉(��\b�YPC!"JM�[P8��Ք.����`m,�޲������1�i��d?���GW_��U
D>�( <ݷ�i���(ߌ.b6�⮶��oZ���xK�U^8�>ǲ�����>�םC�8�f+��]˦��N�i��ҕg�p���㪱kh�`��7Ps��-L�70K�X(�AO�[���{��Ư��z�٩3�q�q���l���M���U#�_t}���wT����P#���
�8�n�2ocWǩ0

4�0Ɗ��;���Zū�q���9YO�oykX��U/m���.�T�+fɅ"���ok��b�Y�V�mɹ��7(�J1s��Q :���a\��YlKk!��!t5Ya�4-*��,���4���s��v�t	��b�R#>Bt'�Ps�+H�joh͚��E��J>�G��B���[+9	���ۦ�ߧ��*L�n���:ޢq��_1��h�w|:#%���C7��OEuŕ� ��np�|�\�UGؙ�#��h��lǲ'ꘜ��UH�s���qA��َ��V�	2p֧�S/d[�z�4k5jP�zu{*�/*�V"��r)lN�.���[�t�btx�U ���ra^�/�E�Ø�+�C�Z�th�W<�M m�(>�^
`\\d�.��u�e�ؼ�����Dm+��}�@�����}3�9.�ތ����If�k���P%��p��t]�unR�����`;��R��Ii��ݑ5u�l;o��r��s0�ZBSJ:�I����ɫM��WA���CY�d���FQ��9�8�2�K���X>��xGo�郍c���te������+s-H��kbM������p]d�E�
�F�w�t*��L���*�]h/����L=�,T��}�,��>*���ejAv����{M>д�&��]�Bq�ܮ�e�hd�s�=�6�{e�t�YX��7V�m:�o��MTw;86{
�9$o8kpn*�t⾿�憎���l��p�W'�4MЩg��b!u�o;�i�k����X������u5�΋]]{� �K<��4V5Np,�\���5:�i�;�φ��[inp�[L��m	�{VΩE�b���*����:vQ	gpL�W {��&�s1f�3rv$0[Z��we�Y΢�m�bUX(�r"�mm�,f��i��7Tw9��Ӄˈ�n�Ԭ���x� �re���>.f\�;]˘� :e!}ˣ�C�u�����ڕx�	�7�/L��E(2k���c<'1'e�ؘ�Jd������3��H%�2���  c� ��v蠺��8�v��hH�7�K��h��Wt.�y|8t�-ڃ_��% ��X16�!�^�S�}:3J��b�����:�O�!B�h�Yn�WW�l �F���0u^>@ ���ap���$����ŵ����hy�u0#�=�[��]*J�-��ɝ�#�vR��W��N��#�d�ˋ$�_A���3�C����S�/vjv�UVۖ� iGK/����#����l]��rr��l�~�譀�4Cu���n�������G�ֈ�С��N�F�N]5t\�t�p�T3��$�t��B����]7��:�m��$�7���&0g*��ԩ�ar��J�Z��r�P�z�#��	xga����
�����7x���oh2ҥE+�BFD���#���jƮ�Z.p�z�.��޳�ˠp�����ξ�jl�Е$�
�0�����!�c�����oZ1�� }��+�v?����1�^w.��h},�W4�8�j7pu�$��Ƙ"��׳j�4��k$�V��C����z���5b�z�\�O<Mk>�lo ��#�.���Σ/q�t^Q���~��e�es����AV�!����o4�����3^V'd E6}�>�wj�#�{�'�O�k@�K��RZ݁i�'h��3O 98.�a�5����d��,[9�XI	h7k�.��ˬ�#��-�s5�.�#7��@�鳩�|�ޭIT���vc�eݷJ[J�� ��B��ՠ.�Y���G$�� ae�u��B�o�c�-�;ڍda���ϳ��[חץ$��h��ϳ$�+40��V�ԭ��]���WY[�
���Z;�������u�sI�:�]h�M�p�tZfE��R��Vm8-YE��r���frh��>�uy�K���)L��^R�M[���r��+�޳mkZ5fI'D�����>ÙfK��q���d>����^$G�^����1�]�[:��e'Vz_ ��{ز+�W�qG*�cÏ�ӍI@�:��+Ց�����>��u��M*>$4�8b�F��_*陭�Ȁ�4N�EܳH��<��*#�Ջ����{:��PÕ����ٷ��k�,�3�W#�`ů*5�r��[Wu�%+���H���^p�V˗(-�^Sw����^�g)��8q��4�_S��nڜ¡k��KP����(�lU���%Bܮ���"��}åӾ�E  ����Ϊ��C�����^��`��FI�/,j��*��]�p�W�T����΋�G\˜�ʶ0;\w��&�h]���hS:R��[i3{�"���s��ݴ0��S�)����O�V��G����!�#cFd�sXu��8鼥�V�X��cjث�
��R�a�z�n匂�oeo-F=��/c��Z�R8&�q/a�0f���s�T����Ƀ��X���z��=��U�@�6�}�po](@�z�f�Q�U'e�����ᒻI��j_Bjb���w��@]�=Q�H,��)&mp��e��.��d�^*��{�#��8R�1sO��"�5��e�4U12��g�q��j�00���4��˽=B d�T8���xIw�zu<-�|�t���qhє��ï�NuF��=Ն�u����ޮ��p(�*g*�O���Ŕ8�AعDM�x������H.�s\z%��^��I-F� a��|��쫋:!�/kk�U���Ȯ�R�[�ܢ��e;2��:,�(7Қa|�칯GB	�}����������l�*���j�.z�:|/���l��5�u{�����}$��t�~}|�ĉt���ªeY�����>°��u)��/��B=,j�e�lcᗑ��	�v�Y@U
���������T@{��i�������{���o�v���w��:�<�;�<�#�v�,v�xt	�)Pe��QԎm4�
!�.��C8�)�eR��CȺy6�_R1Q�X丂��/�H؆�^&���8�`��Bf1���A}���[ŊW��Bu�ݦ0n���}imF-�4��!�rV��vo㙷J�Π���l�.�L��"���x9^�FR��h��cv�t&�w9�;��&x��
�Me\i�L5(n3�*�s˘���ɞ}a�u��Y�`g��35��qդ^�ö�C1�'Y�#��"t)R_�YV5V�9?�}�O�G�v�k�Z���.9c�R�M�/���{�{��J�4D-fuX�^E�h��,4�r!��W�k�8�!��ujj�HUm-����pѠ�1���+���+8d�+���:�5c�t�}��q�T|��+owq�`ۊ=֞ǧ���/�c��śI�l�t7�ܝ�ț��,.� �WYB�ilWPvc'l,w]H���!�l�	�A�=f�ae�sHl��a�f�9�܍={
4��s���3��WImgnL��V[u���)�&7s�i�59B���9Stmk(e��"�kkgc遬�ݝH�^�J')�L�]�jpL�����)ͱ���ιχS��n!k��=]�B��3q���Ż�SO�q�Pˢ�4^a�E��Ѥ�	�'B�m7L�m�I*B6�$ԡ�%$Q���T[4���DE@h�	��
!�["�d�YHXm2�L�(	^P�=Fhq8���)��t�ߛ�8�FÜ�����������������������o2��%����Q2�lP��GĚh5Xg<�~���_�g���`�� ���Eqh(Л�]����wb٨����c��N-���|~?���������_Y������:}�j(�軓��i�k^Y�+fhs�T���Q�1��%A�=)���q4H�v(�Z���u�5ZҚq[��wj��g̹�R��Qv�ب�mb���: j��:�1,��C�%8� �d#�&����k͗�y"�ۻ��tr���؂�d���v�ܚ��Dl�4^]��E^`�O=�SQ��8ǜ���L�7��ƂO�۾�:����m������A��K�ˢv��1k<lMATMZ|���]tn�;�U�b����S�O\) R�(��ȣ�T��B�,��v8�ui�{�.|Ǖ�EOh�lwd��Ʈ�5[������d��|��� ��Eyk�7ml�cF#Bu����<߉�}O�TSm�����m�v�����y5�m݈��UZ5[����Q|;���n�h)��~>q����;�/?w�G���Ϸq���;����foy��fcÑ��ys��ҦqGs��o'-�:-��Y{]�s�B(Z5�
�O7B�n�"�$�hB���R���t��R��N�h[�z�i�ô�|Ŏ�fZ����=�IN����]$Li��~����y�I���(��|�?`<��w��v�9��p���{�N�
�6�-��w��.2]g��iz��_�e�w�/��^S���A�����r��Hq� I5NbYmC���"���ʓ=����Z��v�����>}Ϻ2}S������)�[C�M]J�����+dK�s4�v�Ҋ�lyYl��33ѹ��6����~��W���z[��W��/e˼ﲷ�Y�n{�޾Y��Ƹo��f}`[�mQ��[W�)�H��z����i�=S=�����zx߻��=����R��+mW�w뼴�k���� ��� :�잿����ױ�U;\�{zت��zO5CݞvZ����^5����h:�B�Ӷ	�,v��5k�* )�wvg˥�=U>"�XS4��
+}��[�Su�H\=y�yr��M�NܑfV9^��yc�y�|�C%�(�C��O��e��;��[J�/����څ��%�W�7���o���$rsí�;������)��hԣ�J^iC�����T�EY��Z��-���gpFV���}P9]���x�76��3�>�c�-���V�;#��K߯C����K�����lJoL9瑱��=4������*�V:�|�.O*����F �'Y=��>�b��3�C����:*�ǧ�6��#R�	G ��&���WYn�#���"|��۟6�'�o���N����j�h���yV�5n��y�W�Z19�93���G��W�[�5:�����/�o�r�u�f�4���st��{�F�Scn�(�p�2qƟ4NQ�)��Ld��čNXyl�>�m�x���$�.
�<��='���n:[�ޟNp�s��ι��)<1���>�ؽS���6K��ͦoě�[C!�x>�7��s���M�+�>�nw��W������v'�$O���i;�ۺ}�����gx)�4gY{:�ʹƋ��>'vs_@��z�٬̑y
 ��0���T�O
���U��I���<��J	��wܲ� �%
�,�$筌����}�1blh��󾿄O��N�|J����ө}�9����&�r�31����S�{C��4�!E}�����P�-�a��s�B��e�u��LiŽ>��a��xN{�U�EУ�m���ؼ����S��݁7��)��nu�w�M�_���I���:�J�=>V��q`���7�aeM2��h�݌���2{ט����dA�u>��*�q�y��}�+���D}�#�N_{ս�xK�%NStS{���P�z���e
�w�ʫ2{�"�"O��в��R�
�:z����b��G�PB�]�~�^ݹ�"�^/%��F�`ݟ=VT���mC�l�ӧ ��P��_��t�|���sϋ�2�V��Z,i��,��8��n鼊����:^yV�5s�����_)���ݖ��ٝ����	z��~k�>��E���V�ߕ-�N��i�}g���c���y�H=��Ƈ1q�Ꮇ��U�9C�U7O�b��r�w�M�x���j��+���k�8��hj�?`?k��>�f��Ä1-��=ٶ��U��-.	�H.�������xf�n�
�w/�;޻>#3����FG�>��+���V�=�G	�����̘���`"n��s�%m3)>��B���=uw����F����'fX��"�At�R\;���w���@l�b����l�pMb~��@kG�hU@�����w�_9~��wn�!a�3�@+]N�v;\K��&ww^�{�jձ�FRP�f�^^w=�|1%;��ԯ!��,�&w�`[{�Ֆv$]����4�槒�䮲'sڊ�؝��&Oy�2��#�7˵�*y?���?/U�I;#��}ud.^���x�z���I�/, ��0d��Q�M{�1:���z�iI�Y9�t~�(����dZ�Z>��ܕlڵ��N�]f}>i)ܮn�W�K!{����T�N�w��P��.���>W�������gÜG=�Y��gӪf�����n��i�tL	;6Ⴣ������]~�Ic탵%=U���=m�G�E�$�6�`n�{h�"�g���3��p���+�>g��=O�n��o��Ζ�K�����]��Q�Iĭ�~=�Z�5 4�g-�¦��������^L���R����X��R�;�.\i!ef]��Kx��f�����,��:w���u)G],�$:��y"&�e]�9�O=���]�!��I�kXd�Auw�H-i��7R�6���_������OFr��<p˘cU|�jS�ʳF�:(S A�TMF Q׽I�51WA�1���P'����\֐�G}��}i�*�8f���g��0n��[�Z�
�i�13T���`r�����4!�K��t٨�vxI���^d�ロ6�k�}H�&m�p�9���z�u��nF�˖����������Q ��@����3�M�8�ss�X���w{io.Y�{�c�52�B�Ϗu�����J<��ߙ��S'������2>�{�{�zL�[������'�Oy��{�y�?�� �\B�x��hdڼ�F�Ȇ�L�8�8tK�R�z�^9s�����#%k�*(ζ�Oz�]�`��6�h��>�;��H=�oG;6L���q�5��`>���E5�+u��O�_WzLߊ�{A�+h{�WP<�h�Kp-[��G���z������N}�����ʸl�g� D8�M�MKXڳu��5�J�_��萦pp*2�S-��۹Z�hr��Gz��ݫS.�UE���33XZ����ۅ���
��߽+�{���>κv�#��O�j�`��_vYn�r@��N���,9JWJ��w-�_+]7+7�K�x�����o
ܱm����Z6������us^�<�]����>�J3����6�h�Ǘ���^���;��!m�!����/��Jv�&�	����<~쫻���[�P�Lm^G�ik��@`��-���ъ	ݑ����F�����z]zv��<�y���it��7t���[/�uB��sɷ(���7q��|�[W��"�5����=�hh��5���@b��^��о?Oxnm8��.#�x�X�`�#��U8����%u5<N^�b欰�
��ԗ��rh]mf\�Y���)�BQ�Zu�ﹷ�-�� wF��7�N[����6.�+�f������5_��{���2�ŋ{��P��{�2���O��������S��Nz�W�&��}�=p��x�=��}�!U�k���Xȍ�4�!�wPy�ּ��R�Ć�u�H=���&�QY���[|b�6Ob׼wb�����p^y1����c6���%�j�ƕ���q��1Hm}�k��u�`��Bj�N?fE&Y�����L��%4t�QVҷ��xY���d]5gk�W��>&tK�x}]�� eM����b���up�[������Қ�!���zв��<��BuW�yk=���z��L���+���޺���S�6�zt�L��ށ���7��t��������H��x��_�>���:9�J߫���۽]㼁���l�����=���>�{^�^�K7����q�%�C�:��]�buI$;�����&���e��nt���>i{���So�N�$��W���(z���]X����[Z��XL��y�nk����c�#{�u'>jy�~8.e[Y�_;�Jg[K��Mj3�繶��(]�]�[�S�R�A��!}����>�K����:����nc�fM�]ŋuK�dW�_��pNOy�����ƹ�{��vr|�C�� U�9�X��0j܍mb�^j�4�}�9��P!���;h_ݫ����(O{Yߕޕ7Q<����q޹F��[j�˕�:�8v��"�|�����u��Z���݋0_λ{Rs�^ c�`ﶾX����c} Of0]�#�����9y��}{���NurU���X�R��t32YC��i��%ʫ�Ë��~���yMJf�b���{�WMu�/�;{�(I`�y�lL�{ރ3;ym��PU˿+��R�6{>f����T�e�����[��fl8���rz�$l��&ĘM�Ň���O�k6��k��<U@M���5�2��d�xy�����ky��=�}s�2RZ~��XI�y�>�q�M��n�<��/T���<�����~B��eN�)���o�C�`vZV��]�k��˗��N a�v�z����*���p��%jA>ܓm���^8ϣ&�����|~����{�W�}�ŏ0�^�p�7���t���9m��w��q����bM���U��r��Uc��Йɮ!̝n>���'x����uz.�z��z����Of���W��&�������l���(Bs���>_}���Uk�S�<i��F���F��VT�u���ی07���G����P=4�^Vu�_f���ϓ�����Ε|�d�H�띹x,�t��Lpwt|�Y��|�3����\�����&nF���Zz�s���MS�Kj�����ohS\���ě�M\d�#��(�D1@Z� *UW�;,�`�o*��LZ�A	�1�qU�>�1�~�y�^��N�9��ݸ�e���:��^�O=�{���ݼ����͐r���6ـ9�YA�!�kL�_�'��s��h޻oG���`_ϟ�ۯә�p{�$G��;��(��j���c��f�^_o��'��s�V��-������g<kpn
e��'�w����ѕ;^^:��,oY
�q��m�$^S��#L��r^1+�6y��ou�*��|*��2��ܯ<4f|W��Mw��%Ei�k��m�����/`>�c�Q��{C��~�.?ӿ.��&=�y�5�CbD��a:+J�ͨ���	݀��=�2߬3V�)}���(;|��C���O�����{)+���*�;��~V�S�a�]9����,=���6��ׇ�ܙ�n̮�+�����x�??;���cB�x/�1��Jĳ��ZF��2ʒ�T�'���c"�izK�o�Ԧ2Д�z�J�RAqW(ӥ�KjS7F�BfUS�X:��A�c4���ce�YKeˋj=�ţI�@M]�w
����u.Ι���&˖9Dus����K�A/+s{�vX���.�d��cP^^���k|��j�������[�f"E��Fu$�Q��e}zpO�z���XQk�S�����;b�}����n�[�>žkL��M��� �<X�Ͻ�w��H=zk���O�����Lwz���_{��B��5��v�i�;��^f_ym�n��L���,���[W�XO� m�>�խ��˨�DYw]��}~a�S 5��	��������z!�mz(��s�+ű����{�Xi i���޸e>�q�C�F�O�m��~ϻͯl!����Q{�ǻ-W1���̿
5����|�*��z���a�G -���o�o+��mc��+=#�{|��2����Cj߻~ʍ��8�\�i�Z�:30�f��R{ta@�m@��o������[��Ü`���G���<? �Y�f�8��?����9��2�t%/�N;IՎulS�[/X?on]o-j��9�� �j�XP]� �$ep�o	u5R���M^�/(wbQ^�eF���U��e�=G�<W�yoA�|]�P�Rgk!���sx*Y;}��������Dө6��c��z�*�S
A�V�Y�e�L�C�m�����u�k�(a�f�M��c<ol�9��#�~]�]/���Ɓ���u�1�'9�s����t����t��9u���gY�Z����y�qҫ���RQc���bF� F��u�g6�떴LX�nC,��Q'4�\X�V�Pt�ڜ^K%@���lg�����R�]Ӎ.V�}] ����~��\ʝ��]�ʖi�u�K�Տ2�K���EGq��V��^q���єkV�UJj��:_�݄,r���m�]-�z1�(&N�r�����2_�K7�tM�Uo<{[t�l�7�3�Gm����;��#�\�����e�^�w%+f%	�Ҳ�9�DbV�0�wm����5�ػ�e�!ʸ�rP�B(��m��x6���z�vr9����Sop�ԩ�%�]z�bVq�ܪԨ�+0��J1õ]�ñ˒j��OH�N�h[ʉO,�-�y�6���峭�y����`�:��6�����ƒ��ML`[���ڎi��[y����/$2%�XD�f�\���N�����l]�wyf.Ӫ����~FQ��q;���y�Y90��\�?xd��� �;���E<��7�@f��;��$O��p�^F�"�z:w��ʍ\Xu_1LZ��6��ԋ�z�@h�s�g'��o����7��N�{4W����l4STFG��9�\L<̕���+�1�y[ki���S��f���)���}����ܶ�b�Ų���]QZ`^��t���\�@���;:3gg
��<��]��Y�3�nnӦ�0G؅e�C�B�MYu�A�����O}�L��}��{lZ�E�E�(f��I�Gj���."�σ��;o'I����F�
��(��uadznc�j�o�qgV�X\�ԜN�������螗A]�l�ܽ��"S��e�>1����ҝ����2���du������ (z�s�@�x�θ�v7:7���\{����^M�p���pHyK%2�}�4�P�W�X�wWob]�e�P��8��RFCjr@��E�YݜS���A�"�r\# =r��	��m8�8�ģ �:��&�ނ�5oV�fKNh��G�YV�Yk4n�e2#����ј4eZRr��ɮ��T�mu�V5��&�&-�$��u�S�˙v�Mm�,b����)�'r�7��ek&ݛb�N�����M��������޳�|�����Y�gl�i)����QN�1���F�Fs9��~ߏ�����������<���$4Dӭ�����h�H�E%��'b�5AE%:"3b	��>��G����\��?G���]+֝[cn�Jv5WE1���5���<���~>>>>����ϣ?�������uZhq��|y=h�1XԚ>l5رT?~c���)�]	��tc4X�;ƈ��Wl�\n�vz�m�[:+���*��c�����c�x�A��6��(�4y�;-k�r��Zɭ|����֜AEu���mm�V6�6�v���la�G���i>yo�4�P��'�����n�Z�#l:���]5V��"��#����[b-'��:c�k�X�(��)���b(km�5TbI��Ć@��[�F�ͭ�W�%�M�bgm�Ζ�J�y�u˂����jV�"9֩���
�N��z餫���W��~��z��0���?{�{��ߵO>o�[�0��at1c�Q�>Xը������h�6B�(֔ No5�S$�':.��uvC��>����z+��ơ�.h�&��T@��qv17����⃎���H�t�s��˪|H�lQsGC6g{�e*<�q��� w*�g"�������d@au� "�;\�5�n+f��A�Nb���=��g|_2��p�%�	���0��eg ײ.^O�8�=�y6ޡ���u�9Sk�}�kiǭwۀ{����3�}g�Y�@ܧG��C[��w9I�5�<ʩ8]��*�����h�q����]/r��]l��@x4�s ���Q��V"Iv�=@rGuF��j>b���ΐe�ˊK��B�å,f�$��A�{�}�����Y�^�+G��u�2��И�Z����J3
����g׎2\z6�1Ȥ��2��xRۼ�cY���a�/dF�χ�'�a!�#�V5��R��R+f��> a�닆����$"+���P׬=�����y��:���/��|| # e�.@�a��x����l	H�kU�7-��J�LvT�ƪ�����R��?\�0���^�RX�~���:@�c�d`Ml Ƶ?�� .d�5�uw�+/U����l���\U(*T�>��Asb3�:�i�tf6��T����Ҟ�n���W±���m8Qhu���Է�;�/��o��f?Vؕ���\�\C=����#�D�Sm��js|9�qc3k�_nq��w۝@��^<E��^���<||D^���z���i�>�����{VH�|���di+ q����P<{�5z����y��s���G&�wQ/��H4�{������C�_�On>��e�2��d�=h��@S��DK�Z�L4cq^ʐ�+�.{�Ub��a�Z��`��KMx�e��շ��\ n�)^b�&�8f�cm�7�d�g�Y�O)���м=�w��t�a���bp�şG���y�n?��}�.��^��2�j �~�مu��;�gb�٪�@Dl��;&�� ��4 �+V}���\ 2��'O��@��Tx6��fm4-�3	����ZtxM@f�Zt����?��yQqVx.9��"��G\U8�z���Lia�4P�:tK��Y���؜>&�_%����_�֟��?��HL�����$���O�<d���V2���k�Iߗ��?7��:�,��Ö���=�7��{@�}/M���S�Qf��@�&ꎮ�6�&ފ�oI���6��G.�ٹ����3��O��|���;~�|n�q�py@��Ǜ�1�Dڡ��#]È2X��i>ҟO��@������+�	���+6 g�<����^	(��L���cp.Ũ�Q�z���k-Nm˽C���r����eb��1rRy�AۨA�ʛ�v�
�"rR՗���ٽ�
"�A}v\9H�d�$�$�
�G%/6XHi��v�Wz�ku뼶/�L�ӟ^Ԗ�>�1aݚ����E��o;jP�ɷ��9[ڌCDCV3,@'yñ	�$�䢝���>#���(����܉�ȄJ�Eq[�z	>�i���\�p�@��p�F<��v��m��x�sTz�*���ks�/e۹�N�^�ۀ0�I��@b�-���c"=G_�O�bO�}���t�sL���3gd�c�Am��d���ڔ���b⩃j� �e���[�\ K�i�4�ڕmaH�v�@�p6�������Dc�����כvÑ�� ePI�:�b��A1@И���{m]Y��;�����Q�@͘�=�y�4���ɴ����"��t3w w�<�-12�ǘ�
�
y����/JƧ��[�^����"6�N�
�]R<���B�ik8@�f"�>��`�Mc�i����63}�t��;6- 3.Ŷ!�������j m�7 #ԟu��J8�,2�]�CL6B�J%�V�����O�)�8������bF�k���>�]�w!9�j�f̛�	��<�5)*��3xo T�ĤS�#H^zq��->����T�9���q�W⑜�x<@�~{.����d�,�~F�>lXb��R���([�jh�l��#C����$�ᑴ�v��;�֠#Ώ+>�/���k.tdk���{��]�&@͸&]�B���Ki-	0w�ovgPSkj��T�i�j�L��x�	k�O, �;��u�J�X�������2��V�w�;g*���#u�6]�&��k�Ĝ�Y���q���m��qC||G���������׭���=L�W���k�@X�j��J�:`SC�Q�^��=)��{hݿ�75r��5���T�ޛ�����D�q2�ݶ�Þ�p8���%A����y�����LK���v�()��'g��i��u�D�U5;uNh�Ӭ�WqW�x8������0�)���fD���[:oR k����$��Az T[D�t0��A���L�/������~(�U-�]ݑj���耰�X����᭥��vd��	Ip��.1���R�A���5>���I�Nu��l���k��ά���[��fl����4��Ģo����)8J����[���n��^n�єsc�ڒ��{`�M<���F���+��<��%sdH��p�E[���a�.*��D���# �-9�-X�{���\�~֯P}�L��r�#N��)��������|�Q���=��i�X�ⱃE�f�������v!>G KO���Vs�8G2ŉ?*;�5��J�-�#��=?@�ݚe-�\��:�L2�k��Bm5�)�����s�@���G��k�����m��QZ��%[^B-���s2T�E^f�$�XF��^���H�93*��]��=:�U��6����Z� ��h"�?^(��{'���]N��5�_X�7���YX�j�{c�=��wqsh��*P[z��6�W�V���f�u~���>>> Nw+Yk��X��FbԖ!P
�Ca�a	*�%��y�\*>�� m�N����i��5/��/z�Yz��6�a�a�Z��L,�܁���O��y�T�*�<�v&3�y8�m|�P<�
����Z[��r,���x��ײkP@C�:�4m!f��:ݪ<���6�Y��b/ێi�f�����A�*��o�Ue{��]1ָ�yo6�+��+Ā��~|(Oߕ�}���r�X�ʮ+����|yp����H.�7��I�cN����m��ʽ�D4ۺ-ۨ��vnk�eyB�T���^:ዽ�Fa�.{ q�S��aR2��q�eo	!(�#\'�kw�m�5׊$=�ɧ}\�KI3�U ���9���gi;�Q�54�hf�c���9«�b�ӅT��w5��ρ�{��D�<3%81Z��j�w|�,r�A�f��T�}��qz8��5�=�{
��P����+E ��\�Y���#�D��m�Sӻ���)�^eE��q���^��JB:��\�^�z�������Z�x��9�iTA��H��ݜ�������Y�<\�ʈ+��0��Gx�w�ꄬ��;��ރ�˨�Q�;p���(�q<�KT"�,;��2����fbj�{7]��ɏ��(Ƃ�wJ��+6-D�yÍ`���o/NN�Ki�s,I�t�b;)�U��gVg+a�(S���x� @�D�~za	8��*�dbm���$��V*�� ��(@��dW��'��i��t�v�xGP�}̵|�gxxY�\50W>2�N&�(Z}��
V5���Z�7� �ұ�[VnY�`��*2X�պ�O[��r!g��g��l�oD���K�|��+a��ן-i�Vh���[�2���z��{݌4���#+ѷ.F�	�/d<s�i��t�3�cӻcժy�)KH�/x	h�/d����v�_�n<?=#{j"�FH�vX_-ؠ9�%��{��[y�Tb~n��{�/{��0�j{���w�=�yk���A�Ƥ�`�T$�C&�jȲ:+'O��V׭;���T׬�,�g8��O��M�o�}u]c�b6|�O>�\N�c;����2vi�����
�Zc·^�
Q��^�qv��Vn8�of�@j��sS��=7[Bg.kq���3xY ��'�ԋ��� rVP��k��jN�^6��)�a�F2q�:��<e��-��U�����O"r]06�-`�54�y�ǟ���إϙ�g �qd�Bʜ7�E��ƣzy��ܩۂ�.̇��Pɺ*��3Rz�h�pL�����Pwch[�#j�`�v/ᝋ�'W٣�����X��O��z��W���WR�0ģ�ݴ�[�^s3
���2����p�k�9����R�f��Ӈw>(o� ����0��x���F����M��^�_LfRB<��W�o�V�����惜��Χx�V�e�WxxY%U�v0����F�}%)�hoD���7���E�B�p�W���c�И���9]��=�-�e8ج�/6�y�S!�V���iIvs�!��-K�+r����3+VM���]0�^~�[��C���j��S�	�EJU"{�z�H�5�폍����,r���!>�{����T�X���@��O.�,�0f���)��I��\�2E��x�y:�9L.��=��Ў۸b�L�`R}7%ćl��7
,ߓPw�o�Ҏt�2�C���7^)]�E��j�o>{J�*�D���D��ۨ�Q�T��	�^�Q�2���W��e���XIfF�#����BS�e�:�;u�m��˚
��J=���fG=S�bI�RY����F#U��/<�b3�`����H��!;l{ke���1�u�������,o	t�!��س������N�jx�੤��Mykױ�Z���D���a���WN��	���挌�)z��r�.�!wS�6V�F!Ђ������`���l����H���(����J[�տ��h�5-����j�Q\�&�����[6�%=�ݧ�	�z�8���2����s��S�]��P�<�ɛ%&�ʈ�ޠ��5���ʛY��W�o��v���K��@�G*�v��Tڴ�N[�0��p�4�����Q�SK�����nvBYgMo9{�,1\A,5�y��)��[����{�эox��1�+�Lz]�Bӻ.��k���<7r���AY������㮋����km�����S�Ҭ�n�ve���qŦ8n���������	�NL�\+@V�tyQz�C�W�r&Aͽs�\�361���<�&��cZ�q6�S-�o�\8xٞވ�0�-ʭ�
qm#H=S�qv��w�H�-x��d���nYN��-=Fi^�f�j����d"R<�Bck��D2��o�櫖�A�	s�J�S\yk�������\F�M�=5r(<�4�;��f�9!��ͼIw���S�aÇ��$���w!�4B5��ߵB���T�C]�:t��({��G7����C�i�j4�F��y4�ψpz�G��ɓɭqT�sX��271�r�oq0�mଡ��l�}����VfC2J'��'e2���d�Éa�}�~�9g#�y�RȨ��YC��:c3i����������,�ً;�-��i�̖cC�+�\O
Us/N�K�C�z�tjw�ݛ׭���u�؝���ٵ¸5:�C\�����
M�2j[�0F�`�h�'�+�� ��hJ"_<>��7�������Ͽ?�}�g�7]�E^%2W5�v�E����/��O"\���:�d{p.�z!nKc0�i|v�}��!y\.�����/�kH^�)��E[r�jx7	��{�,�4�a�bo`$�!��e�`/�+�=�tC���js+��K��f�j�l^y冇,9��*�-P�ĺ
=����t�:�6{�+V[��~��\G>h�JC�������B��ąΠ�Y�s-nZ�h83��xZ]�ƣ�9L��+mG�Ȅ�BK���D����u���Q�7����DxJ�5Y���(sá��Rǿ:z��`\�o#��c��D�O��9}dlCA��j�'�E�e���=��[c�[�4�z�����5w>��] _����
��s�ڶx�ozE(���q-Ԏj��5����=�|��ϝ����2�������y��	�0�@k���X�U4fEk�^���v��1��T����W�2<m�05��qP��#��#��3�}�'�Lջ�G\&7=�������K�Cw�)G���EG�^WH�,8ϯ;��(��D�m��� M���������]�'Y�8j��w�_F��_�}>�u���%�{����d�񭛖6��#B��u�w�	��۝����a򸫔��#v�[yW��l�;�L�)j�����Ł�����B���W����G����x�w�2O��_V[G��lS�-,�&4��S�����NuS��#�2Ȱ���F�W]	���i�s��:���rG��'��W��8�N�� \��P�	�̽o%8�w!�� ��y6�ۙzK�!]�S<��ğa��f��B!����ϊ+�ժC)^�u��0r��B�dkC�]�Z7W�������Q�<�Q��a�E�H�ON�o���3�2�H|��eKwe��pK���,��쐨�h�tu��t���u�q�r��u`�*�؈wz}��w�s���jyRy�4�*DG= r�@�s��	8�U��.����2�Sn�)#O�zu�o@^REo7����Y;3�	��i�jG6�T9Y3��D��am��ʫ��]㿍����
����c��T�$&��Lt4%1��3E�LZS�K&������޽��[>+�����H��I?�ڈr�q�=x�MСӒ�v���Z��T��T`U>�+w��A���l.�2���+�+-�n
H�"
ਂ<���fηZ����a��`�Nk�#�ӯ�4�����2���(��;p̾�4��N���໿I&�ty]��ci��EC{������P�)L��fi��9��i�|i\[a��]������C�H2�����F���>�������$<�5���WX����H�Ɯ�L-����u4�1�K@�����ɗY�X��1Ѡ�]������-�y\E6�LS.
zlN��T��}{�0t�^ƺ�jM�j�3
+@R�6y���&�m�)$'G���`�S��p�B6V��ޫi�8���6�7��Ȯ�b�����<����)�n8iK��e��󳕹�6�pm�;�B3>f�b���*�N�1eecɭx8+z��)�W}�Q��se5�
�w/=Fբ��גG.v��ts�E���+�j܉O!H�=��z2���m��gA�ڡ{}��T�M�o\�g:v��8�<�U�TaUc]����u�#o���d
s���:D4�`��ܑ���.�<�� 8h]K`��ܝ!�7���tH)���V���VZܦ^�wYy[QmܰBZV��6n'�]Fn�Xz�G ]��4f]d��|�M�V�՚�f�RE*�e[�W ���(�]���j��	��5m>���f��/'q��6y,���[�U �D���D�#m��ι�hssO@[r�Ý�D5�C_vEGR0��X�9�+_�[��yu3o�\[E^�Z�^VT&�Y�.:m�S�B�މ{��lCyi��v+�xE>�R�BXui	�jv�����-v��]�qu��RÒHvA;X�E%A ,�Q��i��ЛT<s+��	�_y� �y�d����@:��W�;����S��qLܑ�+���]��D�sN�8Va�W�͝�Y���`����u�����{S�\h.�C��:Z�r��pmA5��BbS�-z&�Q���(�bEpX��沕�����U��f��Kqĵc��)�3)d��2Y�{��R�؎��c����J��f݂Խ�'��m=B��W�Y�W�CR��6�I`*�۔U]�|��2��wGJ�qҔ���AU���O��m�ޘ8�i%2�(r��
�]�9���k��in�h��!�h�e+o���|6����hR��+�:m�ټ�S��F��̆ʸ�°qu.˦��y�S��ݣÝv��r7@Bj>%��gX.�m(D��(v�9h๡A�U�iw�˩ryTtb��,�8��A�|�J%�-�o���=�W=��9or�Y��nn�ƸS'z�e��ڭOv"�L}��hٴ��H�£�Sv��u�=�#v�t��
q�����}�Ƙ�N�&��
����f�2*'�N@����I�V최F˘�X�z����ɺ2O�eb����4��'z�d�y}ǎ�R���6�i�S��{j��w��n���l�[n�*EҶ�>ӳ"��Ҵ`H���.�o*��
h��_3��4���l����H�R��`�%R�:I��� F���* �e$���HSm�(Q�i�
�4�x�5v)5�
�E
�M�JN�a/:>`-R;$6%\��r�\*݊(j�ӉT4��>����`�7�[j�jՍ5��mlUA;��[`�A�>�	�|y�~�������������}g���U��iݷF�&��T�A���h�.�DELQтs�}}~ߧ���~>������?���ޝ�]-���1WN�ALl%k`խE���*+�m�+�j?m4��N&�y�?O���?O������3��}��c{�"����h���w��u��"�3Ӫg����cu����.gc6*���6��[l:uIG�F��n�j�4j)(LF�h��V����b�-�D���':u�M��!���+E&"��MccE��4m��憴��ں]t�蠉�A�N�
4QM5T��9��i�5��ty-WAѢ���F��M���U'�b5[�lGE�E%]��qQ]F3�6����Ph�:��1����0yU���b����%���i���6�κ}r
ާ׀�D%���\�cq9��"��G7��P��T{������K�Ѥ#I:m�,��_���d�ee R���}o�n>�WRO�j�R����W�����/��Oe�N�z/u�(�2����,�}P��}���R�5����y��V�t,f�J9;^�q`[o!R3r��Q2s�D�~�y�V�[�ڒҸZ �eL�nc�5�2�Y+ݳ�N�O3G�������Yz�jZO�3/h����G���!�a'4�m`\�ji�y��҉��<�W->k3�HG�.�[��ݮ�[�&�J3�P.����%�F'K}�,�����d;SQ�W�r�T�m(Ǟ%TQ=�\/W38��O��'F�z&Q� �xvW���:�δ��������f��ׇ9�.�]��<�8T��{����~���t|
����}0��5E;�C��p�3o۲���ӵR�O����e�ϧXH�%����j߁N�+��U;�j�"�k�"HuF��ź�����0(V�V��ˀV��g1Oɚ�@&3�&b��#�ל�JmumZꞟ{�ATWY��t�ĭػaW��E�3����}p��,�����G@2>�{�Z�L!�%������cR,�Gv�6��E;�o(i��3�M�J�h̖&�E�d{&x��6r��+wT����m�-��W\�\ͱMu�x�:���Ɏ�e�ղJS'<����HE�ν�Wڧ+.@�`�m�'cN����y�[�{���� �� 3�{�ͤgt��륳�]�+�M(�UT�t�:�*�\,+9��A�&���5146�|�Xg��6�n���d:M#y�mIz=�ꎺ��.�1	�㘆�����ŭ��0z:��嗚��A�]j=��^8Oz�|2Nj���r{�4������T�ul��`�.�z���g�����·`�Z�Vy�}�X�Z~L%u)�).�>JۣHX�p�Fɷ<4�ZZ�ѽ��'a��8l|*D;���6�?�}�ș�(�o��w������W�Yk�t���v����7��C�p��'c�>x2�����4��휀�N@�M��5��/�6M+�&i\T�|��)�nĴR��洖��7��)	���x�q7wQ%&Y�j�d�Pj�N�k��y���\��z�*8������D9ٝ!���纇6���x��&�Uu8^�z���*��aqך��H�Tm�b��K��i�kC�N-1T��\Ӛ�g�_�U�{˾��w�낱��U~؎�v`^�Y͆�b8�uפX���0+�K���n��U�
����6�3������/�*U���qx�u�.��h���4���Bܲ`����ET:t0�B�����)	%</��RЭ�u�ڍ3��f�KgҜ��]�3d�r��8gv�����7�s��o��_\�ԔU2\���߳��q� ?�
Ȥ0�H�x� O��wmxK)0��g:5��)'����� S�5��zY�����/-�I�ݶl|TF3(��v��+����dk
c@�sA���:�S�G|�k��x��k�y9��k�X\�T��7��0߫h�/_lH�0�*��x�E�1�5�%��w�{pzԵbj̫�Q:g#{
�s�Yʩ�����)&�ș��<�{3*BPd��^��ï��\�f+��8�c��
�i*����L�\d�DG7��W\�J�{�'��\Q��zzf�T���Z"�L���j�ؾ��c\��><�ŕ�g{<���SV7׎dEJ�O�|�=)d������w@n�����z�r.!�Bǹ�;Ha�X.!t1�8�p����1B���_5N�G*=�	k�g{\�&�;���W-�v�G�>����A0*$y7��FU��m0����<�M��h����b2��v쫞���	��9�A��k��k:`uy����������ٸ�L��J���mZ�~�Y�Fр�t?]��k�\kc���V�:p�o��Wi�����p9�,\xG�P]6�PK����<��ؿyhޏ����H?q�];����vÛ,S���:o��^��M/�N��f���i�p���q[���f/(9^mwNh��V�9��ʲہθ�:�=\�6����knR��v_^nb'&�4���{��x�4��Q$�<�{�<��}������(� n(��c)48�3醑��_4ˢ��;0�o)i:U𺘙�5���=t��r�Q�ǥ��T٪dx��l8|��+#�	ԙ��mGY�ao��\� �5v�#�1�S���ޞ���጗s^�R-Y��[�o��fm��V��`�Ƨ8���8ӕy�R�\�;�ݐɷ<���`C��"�Ί�.��*��\�Y��[ �xZ�a[��#d!B��hpTN��I�8��.6��s���^�ؚ���?�3͚����S=���g�ȣ�,h	m�N�4�bqj������^ёi��FH;���Μ�:|S���<P�����k�b�D8�ifg��Ju#$�0y݌x�s�Ή��:�L�����*������@�g(�J����[�T����S�2B<��/&���U]k/;vȐ���giqV��n�T׺�k4&��I��mY�==U:����f�ەeʺv+�z}��h�t��)��C�}��|�kyq̫G��o%&��ca4)]]^��qy��]�t*k��9D�\hA9(�u����|^W;\F�Q�!m���f���.�'�Ѥ)YV���X�ڔ|�f�î�b�v�;Y8����m���T�mY�������Х�yC��y�ib��8���E��h5J�h ���J���T���]�?� �2�����T�a7�����?~��ͥ�
I����2_��4�m��O�X2�Q��>��)���U�	�2�K���e��C^�"��ӲHsۜh��@%#LJ둏����ƶK�.HP��Cp:b��39\ɔ�<V�)�V�6j��1CUD���B�����֐��j7��"-)��'���1]�ܶ��D5Vox�;K=Lڽ�!4V?�M��R袹tqJ�ty՗��]xfb�P;��f�wD��e�2�͞�85��bܳU���z�;�[�Oe�D������IB�kqM�KYO���M��Q�6���� �j��Bz�_��aSM��׻`I�����üʹSm(�ϊ��s�h-kI�x$M0�d�|>Ҍ��"�UKb�կ5�|��������(�3=���y��n-�?v��])U]�������%k�kL����R�T�qP9 Rn�幤�L(!�:�R���C����,Y�6<�����I�}����6�����[�z�%�L,��w��[3��
o`�.r��h^P��[�o��+�c�ƪ��JS �<;#�N��%cg�`GW�3ם�Zk�I̙[؛�Z�]���-U��<wyݏ3Bn�ɳ&�e�O5曓�����Y�>Yt�o��:Z�n]vA�U�i^UWm��ZooDT�p��&�\���m�V�}R\I�\��ܲ��K�m�mX�tcDT��ӳ�f�� �x� x��	p� ;������?���Ӿ�q����$�S���)C�})�F�� 䁚��E��I�s�!�-��j����쟶�+Z��	X?3OK8|�aA�ʚ@���8WΎN��7S�Y�
%����S�ï��v�� �ۆv�_T1x���kr^a��r�T�=�1�_��wG���*��=�^;�Z�`9둝�2�Uq��"i#|S��
M�[�8�Kʋ<v���2��UT>�gQ�U����u���5��3KzB�D�:��@�G��I�hp������ʵUXA��c$���s�@+֜��~Ɛ��V��Zڹ�Y�"�ϯMM��&KƅȎ񶪘"(�Kl���#@�-����E z������;�(�1�tsB�ӳ�0�����I{��,�]0�����}���L+�HC�ܧ����5�:E��x�a�4���`�����?v��6xfy��"���f�5���P����"��P��v���)��|�>^[�Ő�W��H��"��Κ	�ޏ�<t�]k^�eg�iӞv���#����v�u����2��ư���G�d���oں�.����A�g{Y5oW)��3���=���[z�UϾ����~"�"�e�i�pV�a�蹢:���\��C�vgV��i:�����*�lNy���d�ݢ�[?����~"�¡*�V�g������l�uq8��4Qu����_٭�i �XL,��
�6� g��NVo�k^q���C*�3cm<�˪���Z^��| S��a���c�s����@t�t�g�T�X���]n�΍.!�)8�E��Tx�!���BI�ٍ:��)�� *[�}���F��7b�{���CЎ���I���\�M�-䪪�5Y����0Ws�cq�"��'���_�T`g���ufr�l���^2P�؆sb�^e�l <4�0[�,K�U��U��^v����f��¬֫Ι��#���yJ|[v]��vF�O�0�o�+�ȡ����b�3�FCc�<Tݛ�ne�(.��*=�1���ˊ�fe#%%ғ#��sɟ;3 '����q�fT���Òj��s�+�P�dU�%/=��Jl�#z�`ʮ��;�
D���S(J����i�5 �QJ�n��SHh�g{�����+[�i���A,�"y=�0��ѩ^ɻeч�ۗz��'4w�3�d;�-�"փ�q���@`Xϫ���a�Jh�ҋ9��D�h��O�:su�U�\��,I��,v-�:xߨqmPy��ؒKΩ���f����ъ=��et*�Λ�g*�FY��e���;7�kWo՗.���5|�S��b�F�9���p�(�f�����C�ڞNޛ*ⵝ�r.ث�E콽�Y�N����m���g�������сRO䨘dTu@�!*w߾�z�?��Ͽ���A���0�x���Ez �>M�!����N�$��aK�i	�u����Y��S������_W��]�e�<����a�]����m<�:��}��;���dS�}�f"rm��Bk�E)"H�X�Vs>���f'͔B'��օ֟�gЛv^c�uٍ�,l��>3��Bz���F�NJ�'eY���;�N�{t�=VjE��@c�X`3�V��sf�lȻ��w0�{`��R��Ӟ.�Yd-n2#�����S���2�S y�Yh�^�e��-	�΄%M�^ZgWR�J����mex���&�=O�ex��r������m��}}���&X�B=��kV�4tzy�a��(�5���_q�dҫ�:�S���G�M�6E��}W���i�Bz!����~x 9uoZ��P��7���f�xc��F�vSW
V���Zc�m:�D�<���۔�3��J4bc^~�	�zVu����vmU-I�
Yr�vk�Bo�X�w��.3��a�'��#���H��9˱���|֖f`� �w�j�Wm :�.J�o��ZF2�����d��E'V�n�Z�6�Λ�gm{k�1�����h7�.K�� �����.gw;�䏕ff���()���n�'R.W�T�M�Skη��tʗwח����;wi�;!D�*��v��ͭo��FTeT�ZT�o7߻��o�����l���SP�/�_v�7-���uo��ڍ�sP/�y�,�X�*������>�j�Oc\kEh�u�r�'�jxxL�o
W�����6e�D�q+�9��?
�Lq��6��8���ͪ.��Zʭ�%&}�Ra'q�8�u��+�,���X�SuZ�v�YMGZ2a���n��{���f=�Eq�B;^-��d�N���ȋO����
2WyW\B�Ǌ�����C+��q����;���z� V��ֱ�r	���;�`�ڥ��&\����M}G��x��RڊM��(�1�J�ez:�9��+dKE�W��x֑��w~i�Qs�|�`�Y��}J���#�o\f;v.���?��YHX�J��d�J���u8�gM|�h��؄ƶ&6O��T��y��	ƼP�B(�����Jۣ���浀�^>s�n�N�!�3�V�N1�R&y�6���۫�>.��MM㈋��"��r�;o�n�\�of����s��`Ure��qk�j%���ܸ�Z�����PJ���6�9�������f,�r3�"�W�ﻛ�H��S0��^�j�1t���!�.��K4u���_I��n���Ӭ����N���	�� 5� ��/�]f���|<�.~dt�-�Z�o����h�j�Yae�z�bGOU�1v�]_c���v�k��h4��M�9�����A��"8'���&����G��<�����S٨N��eR�	�����i ٠�4��2�|�����-H�PAK�D&˵l������uM;̈́Twu��a&���M��kj֨�q�
�3�5X8����>�M��/^ґ������P7:y0ʓ\�e�@���lhM�e��p�8�[�����j}S�ՋO�SE���;�}���N4o�V�?�W������e�f�2����9gF\fϹ�Hn�C�X�UQ(A�"�6������m@g��ᲤI�S��
g�=<��k��2+���J��f���g������T�� ǝ(VՍ��h��tT�6��fbf+b+���-Fă���'{�0�A��t�k��n��Oⳗ�-n��߀MW6�,�鵶GZ��y���̃5�_˷�W�N-���L��;�PU�}�S�P����.D�%�z[�s�_�}S����[����vr�.����VԳ2D�UFلg�@�z���F�����R�/�8`~�W.6�L�����m^gzL�<��֔{"W]~ػ]��5=�3�����d#������Zȴ��a������'H��`$�z%���ڝ�>nP�C H�h�ݜJ���̳g&+�0�VHK��K��R�C��1m��wUЍދ�v�r.(���y\�}B�������mn��E�fҽ��?L�R�AZ��2�ꭲ�Q�;�#I�V$a~��L)��Dp�kT��3�{�w�B���ֺ�|ۨ�S��!ݕ��G�u*h,�t=���t73{ZDU�n���)�%eu�(Y-�]���ڷ��k;{gs�n^֡�0b2�H��H^w����!�nvp����'s\n��M���)���Ε��H��Jh��Å<W's�][ZJ۷�lY�P��ub�9�
+zf^)�iA(I콤��m���qU�L���Tz�t&��>��[x0Q�b�, 5w���T�y�v��>�}.	��s�=݂��2��
��7���ڤdK9��C%���E�Ouf��Qr%��&�wF��r� 8�����I�M-�c��ZTy���K����y��L��G������t���|VY���.�҉��l[�L<,��S��N�I�n�a���0�4j�-����}�Y�V'}J+�t��U�ۥ�oc�Y6߅�v {ٕ�F���n���fi���g^c�ݼgpuZ�dzb��M�rs�ɜ����$��L;�x��`��t5�����x��b�V�!��Pj<�[6,���<q	F�q����L�÷�������Gk��o]Z����o]�!�}d�[���i��\�!�k,�T�ö�T�l�ʽ����Ι�rĕm'+�7s�Q��sw=��Xh*:��,;zvԿ��V��5�c8� 4q�,��RA�Z\��vl�U��B,s<^!���[���N)��5Ϯ�[��(A;y�o�lJ��#O]ҭGU����{YZ��ĸt��u�(�4u!� �^!J���h񆁰�N�Ʀ���x���\33$�J��P��7��͔I���[tތ��(�;r�cY�B^(���:�����}4�Y$ˋ�vy@;�p7��M�,�()Y�A��5|1�A���[����D0i=qft֪�U�j�M
y�9�+�{����qn�v�K���8��ǖۣW��a�eaT��5:ז�	}v��}{n�'`ޮ��U�I��k�~��(>^�QU�Ҝ�ŕ�8�x�9�ڝ��^t/:����[� ⻯��D���lwf��b19WO7X�Ŋ������'8}�%�-*2��K�v�b�ę @�{,���vj�G+�uoQ��5�%�[p^��589jړ��%s��׻J���e8-N�c鹴;���^E|����lh)u�]��X�)Ag�t鍵�k�.âg<����?O���~?c�����?��UEU����;��Mj��(�V�`�b���A9�__����?������9�g�}&�c5�m�v�n�65��	��ۨ�E���-��ϯ����~��������s�Ͼ�툏vH���:�d��#G}w!��>�QSDkj��
����CE_Q�6+U��X�kZ�-HSUڪ�h�+���W]'T�4�DDS�+m�2ɭ!��*I��1/n�Oܾq�Y��#�z�'X&���F�UA�b���N���<�έR�gч���%�q;fcmm�hnέh��GF&����U��jj����WgMۻtcU�bM?��y�mܘ���Ѭy{ϑ�W�h��Q��*�k�D��4��Ǒ�V�;�|���;���uZ�JTN�Ru�U?*ox :�k���о�uu\�S����1]-�����1{r�JR�]�����?T��0��W0� �PZ�_����Ͽ;��~��������M [#]���҈�l?�7L#sY�J`����~����kk:�w�c�����Ly�<�&l��t�r�㚨�)�q3ϚúTi��u^��N����č!���=�[j�B������fgd=��("�D3���K�/������H���ib�®���Q�{'S�.��B����2�cSy+��h��a���mUo���R�l�Y�AQ�������vS�����{��g�X|�sS��Z�7��#5�`,7`Im��Q-ej��.7���5��x�[�뼕�t,	��1��@jI��qCzC�yn�Nr�2Ł���	��{���9��Fx�$8����=HI��N(�$��},�&����;�x���+VϪ�Ɣ��ptlx<'�aOɦ��b�,��K]�뇽[N�	^�v{1;ٰ��A�ǂ��i�:Lm�����0����^�)�0�����/kN��x���6�;�NE�Ȅ�w�:�^ځ.��^	��0�[$kJc4W.�Ϧ���/'��t��
�8���G$ew��ǒK2�<����'�ѣ�_-����a���dT�)Z��-#0�(�6u�v�5�-b���t���G�����}�*Ք����k�iw2�B��ȩ�����ll�� �UUz��`A�AHe|��D���%��.#�6�qy�ޠ�ژm>�f
�vd�T%%��f�.����'.�#�iJ빛ٷ�C����77<��
i�e�� FH��R��,�D���S*z��ldb����Vsnz�9Du�h֩�gr=X�~"6�Ya)���Zy9)\��@��8�;wR0�,glBӮ�{Kf9!�`T��aXm�X��*��5<�ݰ���vO�����z�l�n��(�q�zL#��>*�y��7�8��?�^�b�_5��c�Ɖ̓��vr_��Q�ү����X`?0E��l�M�o;7+-�ڡ)�J}>��]1���H�h���!���\�,=gXQ��&�jĘ�ழ5��+��l��P��=��}�*8�(`	�v�'O�>��֞�8�!���,_�pg̲�v����(��B4�/�GM%�͈1�փ��!�^L+���/���B�|L�ta��P���'ab�yJ~������+:'g�+�U��n��֨���
�9T��������z�Fϓ���_m�ȸYt؋���C�m��W�p�Bይq�7/m�-�ř{�M#�R�%@��ikb�ׁN�������E��`y�v�U�°�`n`Q�RF��d^�x�g<]���XY�4b;���C�_n�6e�y˴(���e+�	i�h}kHxv�/b���,`��}�w6�^+YMS`6Y	�gQ���8��y����"��e��ʀhT�A��~�~���ߡ>�,����2���I; ���{�r�Rd��
� �Э�S��HR�'Ouس\l��m3P�5��D�wcL4�dI�r����U�u4
�F���Gl���Se��º�������k4g��8�l���:�{Z]�@����!,c�3����Rj�~�KS�>����Cb�M��xU������/�)�~م�	7�"Ԭ)a'g*�{��{��3mE�k/D��=;B���NST�P�Ɵ.x��R �r$U[�FE��_�����~��p"�Wp���tq����a��a�>s�)���Lx�o\�Įq�t�8�	��|�]T����˅�{X�5'e�ֺD�J��4�F8����[V�3�Qi�Rm����Q4Ҍmդ��oޮ�CN�ػj)��$7�ʌP�E�8�
m�'�-6�\�sLc��Xs �9gϨ
�C��ޥ��B�H�y���6���I[��������,|���3�"6�o��aݮ�s�l�	H�W\����b�c��@{!���ֳ�v�=��9�-K"(��uI�](e��T�e+��C��U���ܭ�X�N8��5� Dp͠77nJ!,D��nœ�����w�,�$����\;qǳ�}������q�i���Ҭ�T����٭�7�~��~�����A?��(e@�T2@��"w�������=����}�,x�5{�s|�wC�n�.x�\�m���m��;fp*{"̨i���8���6rqM!j�Y�̎����I��kHۨE���� v�
�ɽ��eE^�ٝ�:;�֐��<z����p[Wo����`����H=�傷�� ��&}��6r��:iڛ�41�aL�K��9��CqI�"��U6j��l��~v��n]��jW��5>ř��� ٠�4�^�zc�2�Y>��Jz����S�!6��m�,�2Y"�e`ՄN�>�8��G�z�L�sY���YU!(�y�L�Ǒ��Y1�L�_�Y��'�<ۏ]�Q�S�F�	9Tq�w��kEy�`}Ҵ�%4jl�{�|aO������z��P^P�B�����M�Р��Tד�=�t1�8r!�b�γ��s�;G{�[uõ�r�L4�f�i�E�-�-u���f�sU�{��3��Z$U�nGbK)Dk��=�W����W��^��]C?�uM"��<YCn8��kϒ�o%]zMp̓,\9���+9��+�Õ|/Ru���KWi�Yδ���}���7Vۜj�I�M�^����)]�C�E���ٖ;�d[(=�����k��72<�&�V���C�3e���[k����G��p��%��7$�o�W���?��H�C0���{���=��}�|J]C,����3n��W�E0��id�	���]���II�4[xmm5��غ�i\FfR�UEq�X�{��V�FO�E�
�p�e[�Z�[�4f��;{P�+jR�;�>.r{����@݈I����c����2�­�����v� J���(F���6��Y����8��tܨ+��VϮ�\��J9�}���y��5�R�d������yS5 �-�r�4���d٤����as'���+m����В$���M~e1�V����2��Z�@��}��X/>��.Z)G��M��;7�'>���z���Ou)�;ya�[\�n��Y�b�r�W�`����EOY~L/sGMZK�m	k��u
����W���yhe����R�X^����͙qI(� -5u���[0� �\٪���D�m\���^1�2�B#�:����ϹO��z��h.��5o\&X,��U����6Wx��eZ8=V,!8j)NYE���h�!x�ܑ����/>�`3\;�`JԽ������N��v5�r�f�=C/���Iڃ���ì-0�����G,����=��lGx�*먂�XMg&>��]uh.eN�I�,#�c
��y_S��(����I�`q���]q��̾U�K�h���`عT2��X��������\2 Ci[�����"Ro��P!���Ck"���UA9�$�	�k��qD���[L���"M�-T��{y�b�d1���K����6z#��Ƌ��BѤ<ˢ���ƬPJ��[�*�/�LNM��bW/H<c�nQ��ΜRr�a���F����-��8b�N��a�ț��(g�\b�@��P�X�Y�P�R�FC�[L朮�O������.Ĉ�z4-O�#F�!�����F��D��9>�b�z�˷���vd�1�&0d�#��ɇ�ɷ0͍<���!��I�J��I>�r�nz1Wnu@�g�@�>��R&G]�d�&�]���pb�?.{�s:��F�v�j�s�/K t���F�*�%2W55�'(%��S�:�Tc�O���A�s�n����l�^�c��.*qX�t���b~֐��̈�S�( ��j6_z���Wa��G#ݯL�|��P�h�kJ7����a��1�Z��
M���o:��{u�Gfj�d9�R�ܰ�{y��'��m�a{de���b6�Jc�]�v�`s���ěp�񮻼]Ī�����bL��*�"�av�x-�)�\�%}\t�_]޷������b�Ț��1t)何�9�{IIk�}&M ���s��#�4��Z���>�}"q�\��[��]��et�s���A�]��͞��s���U�)��UQ�ёaM*��<jMzY$^�bE���V�*�3�����O�t� r��ƫI��c���`��"���.bLMp�{�Z��ka��%?���`�>��uc߮�Lj@����1y�z�bWu�\eTpT�B��<Տ+��e5�S��c��xg���5�X�UA�.G-�^1t��Y���^ANM0�q4�Z����/���hT�[?vE�z$���l�E3T{����Z���/��4�k<�c� �aF�d��u�T��˓�Zs��*ށr��#��!�<��Sly� *p=/���v�E17=W}Nj�e��k[3���졶Xq��Ƈ�y�#Z]�@��Yt��3���׊�b�f��;;
��F���~�Pc��Ą�"�Y��<�W���Iq�)�p7f(�M�=��R�p]�&:��î� �����ӌ����a��z�\�g�s���u6�9��tEg4�66�����V��59ܽd�W@aeZ�!���!�&�R�HT��`������"�ࣔ��Q��#8�c�aq{E��)����m� �@�� ��Z^��e^Vkk���T�������`l��P�G��
�Q��X�u�sV-��oN�8���Pu��^��ޘ.�tC���x	�9����KD:� �������FD!�a䪴�< ��Ӊ���&񏽷�����#����Ј�c��aYĂW��΍�up��p����)�����J[wX9�܄]��l��+] 1 �i1L��P�M��z�a�^�]���um>l���u��6��c_s��BԊ��)�,�����z�'7d_����yn������hZ����k�����B�a����$�<�nXJF���#*:�ȁ��K���P������i�ko��*�8`LZ�;C�N7e�7`֨�Z��4��R 6�)|�p�+�x^0{�)��<�W�27j�Zwc���)�k[5�j�L���╷G��oB:ȱ��յl�\ѓ��� �"��5��Ę�2�e�D=0��tנ%L���mL޸���^Ƣ�D��O7��
��S޾�|/�R��)y1et�6��H�q�:;E(��\<�ڱI;�[*/�~�Y�3w Q��J:p�5���$5䉦���\�б�NJ��S�n��Y��f��M޸�\5�>��/aF�i�y�#ZC�(�J�`�u]�R鳹����QM��]��^��K��S���A�
�S~�j�ù�����@v=\�ՙ��V����!�+%�(�b��8(k
t��^���ѕ������S��	�g:`3�5���S���b�� t���9�M�����}�]��������FT!�a�� ���O� �}p��:���@j*)��	I��5�{�bj��a@������t��N�tfj�}T��~ۓt�%m�^�<D���~!�ڎښ��Ī������b5���Z���ʥR����p�7'}>��}���>�>j"�*^.H4��C�ia%�2��ӯ��b�%i�U�΁��n��|���6v�4���t���u�?�^�>��O%Z���؂$$ꚜEs��{�HSU��b-�	'�\Kf7Z�`͸��"�ü9�v8����z����t�EveA�����Y�ɑ���o_<��J�M��ӘBk��r*�=�ZO�!�՞eݻ��!�İ�>>�R��c"_�qg��u7c����Dw,�
�U;�T\5��y"v�OF�*�TF�u��
�y)����C  _�_׷��il���7�(�n�^��X3�롛��A�-��W�7)�m۽h)�`���.9j<�A�P) ���w\+��(nC��G^�ئ؝-��&&r!�̬��}��h@le�:������g!��K�㚨��=�m��i�0��K��̟�:lq0�U���8�����r�&�>��}�7�ߝ��h�-A�:X��/ =ɖ���/5����wX�x$8I�n��)��t�Y�-�v.�u��~=��B Xs�s}�6��m_ISv܍��Q5ن��\3n�v���?u����D�)�;+�7��#�}���ʨ�d��#��R���u�6j0��H�$r���ؼ[�(K��ۻ��9Ǫ�!kqN�
��4�6b=Ϥu�i�����aa���z��[z�(����T��FY�EG-0(���c!C�q�	����ַ�u�i��`����A�-�n�[��z�Ⅾ�wd��@p���D�1�Of[�a;��ƤwF�1�O8q]�<9�Ԫ�ob��[Sl�&�"h�pl���PTC�B���)�8��4���3I>��n}s�,�Muo��[d���	����oP͇���A�����e����{Vg��ů3j�Np{��<���88�$��y-�1�X	�]�W�]�{�C�N�H���b��o�'ZT�|r2�ruֳ�N J�z;z�緄
�|�C:a�qn�<V�g40[9?��vcO�V�dK��Ym�|8��	��y�O�E�������M�g�(~�#|a6b­G�~�5[q�Rٜ�5*L�),C�K\zc��6<���gD���}���M����^��=���>:�Y+�t�<��p����[7g-�Vz赜�f��`ֻG�*6oRov�!���3L٨j��p&�iX.�W��<)���Q>Gj���.��Q^Q��EGg
U�&��ǎ���J�6����w[6u)�v�us�Mz�e�Wm�+�1t��3_I�=�F����ھ�\�r���Φ/��#s�_b#5GԪ�0�����K�kq;o���{�N��C���ˀh�\���;�qSq`q1��ce��[4��_Y�qx6]ս�5E��V���c0%�wn"q���/�>n�;����8sm�(�=4���B�wrت�QcVV���]ia��X+ �N�;��6���y(��t6�Y7�P-[p;��/z���y�{A�Im�k�Sk!�ȿe^��ԁqS٠�@ʯQ�Y�+S�b�f%����q�r���b����uT���Qε�·�n�&f�Q1�|�(^;]��ӹo�iu��W�2�B�K.�K��59q�]y��G-��P~ų��j��\L�N�r3ˬ'�)Vn��%���c#]=��{�&�)v���!�5�`W�O4
�C��k���>��w�]̓'oGpQ���\���ʄ� A*�͖Yu�ձ*:�PN��h jb�a��P���n���V�u�BݹƲ���X]7P��L����c�YFڷN��px
�x=��n ���*�Nʃ6�\���J=4��nqį8+ū73��B�;2�K�6��%]�n䓑2�(I�-���t���VX5�CUF�t�W=��_�jZ���5�bv��T��T4��?a��DY�^H���A�,ƫis��u�{g������Ә�E��`�da�՝����2��,F9r�l-�DZ�dt�ڏQ���t~uZ.u�s�on:=#�&��B� �����<Z6���b7Q��5o!�Cn䤵N�&w6�l��jc1�Y6�2U�H���o�����Yȟ<ߛ��|���V+�
�+L�X��J������Z�=�jK@!.и� �~����)ջ�e5ܪn��B�Ǧ���(�`y}���wpޠ�j����U�%�
�.Q�$/��8�f[�_h�]+5:9�Vh6h`v��M8��=z-���T-�h�g,L���1ٖͮ��$B� U���oes�𻮦B���{�[`�e:#\���q9��G�r�T�YW/����
�#�I9�6:���V��
j2�j�cQ j���έ�}Fe*�/���_\'�5��&�����~�R������ѭ;�Ó��{|���:���3s��`a�x��&@�9x�G �w�]�A�6�6ƎD���n�\Dպ��m6����͢���J�L}I���8���jv�Ae��#_^np��v�[�\���݈��.��-[��vbKg8�K�$/{���� �5���&i�ر P�r����a6��TBqK����((��A�D�"�$<����\N)�L%A��� �`�hn�xPVk�[ˎ뼶���}�r}���b��wK1���(ti��mh�5xh"|��QG�x��u�����~�������������V����*i6�4SE����WZ���k��J+�Dtb��s������~�����>����g������Om���lQGn�Q���[E۵���1�3lѨӜ��������O���}}g�3��羺31�Z�D^��j�bH�����-���ض�눚�4�l��c>F�<����`"��Fu�4�v��8ѷwWw=SZ�j-�]|�yY'��v3qth�w]�v��d���l��(�n�`��d�F�U1�`���]�A�bۻP[�5��Mt]�.�-m$�Z�{j<������t�Q5֊���s�wsMf���Wcv�mA֢
J(f�*+X�"��]�����E�c���-��lf���5�l�c:��<��̓�����wSF���9�::5][j�:�J<��U�ߑ�ű��ȭl��.�v3�nڻ8��pq�� P�Y�A5�]3O[@
|.I�Gs���U����ot�̏k�w�B����`�6AS��{sS���x���iŹ���k��;��|�������k�
	�%Ƙf��PR.�)��7��	�)�#$�W��Ӳ!�e"A�� �e���Zt�чlƩ�����3�x��[��wEvy)���Zy9�+g��jf���m�R��7Z��@�e�D<�ʼX>�.*�.�B��Az��&�q@	6�0]3���B훹K�M79��^ě�׬���ظW)�)�aW�>���nP�~�X��ݍ�u�_Ym��5�4!.���6ۉ��9Y�ϧux }-
`���k��������q���tͶB̓�nBeFը����\�SK'�`*;1�'��Gk�3��^/���駪'MQ{���HN�G�bؾ��>u��|6�s����Տaӹ4���G�7R�/yI�����YU������@��I�F��~0`�U�点q��{-�O�^�^�s�Uܰ�t�b���Փ
�V1OFD.�p�a���7�ր)O%hQ�������N��q�au�ꗙ��w��Pd�޴4��y���ˎeW�D�x�i�k�Z����u�}���,Qd+zD��>����+n���<��^�jNE�;����&.�T�.N�־c�g~�\����Y�[��ʖ5�{/pp<���m��2�3���RZ�H����,�7�R��v��cN��y���]��Y�(!�5p;ܛ=�{����dbθ�s���D;��;�B�]�j��n7�{w�n8��"#�L08����	�qYɻ��	D��9O�b��xP�V0xi(>��!��P��Yt����)��z��rT.O�h|l��)����9T�\e�t �Io�Jq~�F�J���k8z�"r�j��{[\5�pz��&�"\z%����^��<�3:8�R}(F�_T"'��2�B�h�];����Z��JRY�"<�LT8�j�	2��V�5����b���ELm"���{nTCw&���vr���bfQ�aA,t"9y�:�f�ڐ�]̢mۂg;1q@	�ܗ���I��1��X�\*"�!�`�o<�2��A�[���C\�Q4DT_d�l����o0]��'��cW�:=��R+)D�f�u=:���9REo7�T���-3-)�";�Z,�m=�"b�@&�>lq����SNcx�\� 7G�vW�m���uÏu�r̓}�YX�v��!^?c9@�)���`V�o�[�g�\����s˲���喨�T_-�lhݴ)���G�ێ�M�c�6�:/���9q׋*w�Gs$^��c��Q�q�&�L;ì��r�OF���4r��V��sf�^q�t�Bg.��]fa�� �+�2����2@�h�͡D�"����]�K9u=dF������,�}�#�'����7M'W�{�uw}��j:DK��n�l`��7&j]Z�O)�+�c������W�20���!J���﫞r���~
��T���?��c�d?�Z�G�>�����ĉِg�:�nu��D�}Rkw.�����{��tiq��W�4��|�Q.�,V������&n�ѐ�o���ٹ��1�j����aH.�g�{�zO�Ն}��^���hk�\�����[R1�K�v�lri�Ƕ�fk��6E=�����a�\���W��E-h�+Z��c!���	�k!�'�Ϸ�*1�i�@Q��'l����	��^� ���Q�p�;��؟��Ί7^�g�b��"��}1��XR�8��ȎX���4��Z�
=�v�?=�<��M�ܯ[AK�}�'�i�Ca9�~���#vܪ�;��ݳ����Q��)�p�_&����^��:�jV��ͼ��l�\�r��ۘ-�b6� ��� �Ǥ�����N<�:��7�/	��1�'�=��$K���2IT{������3���v2�X�+���tq0�D���"�du=�!Hk^�'l��_�M'����]-�J�x�G
*�k�Se�@�0�l*��ʃ~5�>�*k����J���T�$��m-�9�U��*��]�h���	��}�_r*����Q&[��3�d��a��2�1O�7Ye�v�a�éwa].�{f��s����7���W���_v˕n=��{e�W���6*ݤ^Mn��g�|<@x�1a�0�P% |��}}����������[�!�0�h�1�{(��!H��M�9G�uv+�WU5Tl6�X^�Z��D��B�sp�hWg;�\68zL����Slێ������#SW��J�ԟקY>=[2��e1ډ%ﮟjF6h!�Ao�.��k�P|���a�Ϟy0��� x2�Kzs\'�~!�!��#YS�D�]���S������H�0���Zkm5�}���8Gy��i�q�:Ş�
��yvh�8.S�{[(����+Ѥ@V�l��i"$��Q�A����¾�7���y���/#�z�%"g�0��u�w���&�O�	��Q�y��-�Ki�6��1�3�,=�VզeZ�:sj�O��zI�|TӨ�6���	}S�xv�ٯ/��T��޺r8A�K��q톶ED��c|�cB":jXf���>���G8�|�h޾��"�-״+65��$g�l	�N��H.�
�j�G���Qd�1�Q��'X�YLփ�>J�v�4f_'�&4�և,��K#��������P���P#H7�
�E{կ3F���兗yJV����5�E&�\tk��֩`7-u�0JW3���[����.^uD���7�X�N��zP��/ͺ$�hY���`�xk�^�vb��n�6�@��e]�}X�g�r\���uA{C��9��<WM��c�9Bo�;�Z<���q��w���C C#�D�P�OÏϿ������,R��R&�}Rm 4�ż<lGs����Z�2V�Fh�a���Z���;9��ꆵ�v��H�Ѯ��C%H��c��>��'tO���X�Y�V��"7H�c��������B��8�EWf��cX��]̄0�9�>���Q��	�'Fk�^W�� O�Ҽ�p���fN5BRpt4+�]+UQԬ��i)�A��b��Q�.9�<�Zs͢�ଡ�l�9UH��������z]s3�ˇ��b!������2m6��@��ڼ؃���.t6�еA^��W�nQ�6D�=���U��hH^�	Hq�Rp��uϬ��R��;e�r��O��-�Z~h>vc�P�h�S�G�)-��!&���[(I�I�Shtr}No[[f��" ��Դ�<l��A��E�	mQ���6	>��W)Z�hF8b�����t�T؎9jf6�+R�'j�I$�|]iG���J�0ùN��8V��9�\���738|uカd�җ^���Ki�9k!���)�9�A����L�O�;������8��H��-�Dj#���TûK�AҞt����H^��,�.u=ߌTm��^C���՜u���o�Gʹk7���ލ�@Ѻt�|�w)�$�8��f�Ɣ�]�qk���}X��''���8�S��N%�oXR8vI_u�~�_����Xga�	Z��)����|�0�Ŀϼ�_Y��^�DF��]�#*����;\V��g�Uhۖ���.r�V�r�Y�Fz,�s
��pu��XkU�M6��5m��s�#mAvVu���t��;����/�,0�x��hr� 2�ց�}=�Y�d�N�����P��wu�'��f�<���n����'��l���c>T�"��P�v��}a�ά>��Xn�΅=��zܔ�E���끒��q��8��o:�kHܠV4$Ƌ�f��d�y��ݣ�V�Sͅ����V�?�ܞ��oe�@�\X��rCJ��N�.QM4��	��Ȼt����)��9��>�V�T��|��z�E��^�F]��S�s�6�۬���6frYuG6�Dd�fn�iI�@�J��a/, ������>���&ih:skQ�4�Х�*�f�V�����m̜]p"�ӳ�{6�C)2����lB#�qa=n1�^)�C5������wev��s��kCF'���nyE�W'��*݊�Ə?������3#���G1��@�\����Le�}\r�A��ǵ�q��o0�Pof������F�bW�^v�Sq8* Z�^S�Y�%r��t���w-���ed���n�m�%Rf�|�8%;��J�u>�&�햞�8����|��m��0�!~IIA	ڸ��jt����~�/��S$����r)M�3���v?� -@m+�S�j�;;��j��^n��M�o�I䱼O���j���2�R4ǥu�ΧSQn:�r�R]J��/x�6��i�ӔA�9Fg]��(�م��Ǜ�k�u��e���K�b�eL^�(���(�$���d�0�`�u��9�)��y�_эx��R��l�۴j���J��6���x�J`�!����i� �C�����H6�+��z�ǘ.[���嚤B�Vk����p�[��l�jx����Z������ڧm��gtQey�i[��D�@���rF
�h��!cF�;��˨Yl�(��o�e�l�=z�n]�,��h-�=��e�D��Vj�Rg�I;�[��x/��^�&�e@\�=}��W�/e@�l�!m�0��س7��Ō���ny�FFO�0Efy��zî%��[�Ww�G(�ԳPq~�ܭ��C0�Ľۑ¯���9Q�p�|�n@L,���a=�l�GiP>�&]��-�k�)k�:ι�
��S�iL�k�;��N���*Ժt�z�e�1�V�g4sq��.�뀸�䲑4�wnᓲ��Ps�c3�� �۲	�]�N�������O��fM꺙����s�2���K+`�P	�.�Inuۥ�`Nxu͕z���/f�B��2:��szl�;�翕�UB��0R&B������~y�����x,����jA���&��q=�!�[\�0p��jD�&�S��e\���Y(�<�`�\@wd[�*}������Vs�!��-�`�Y�ށ2���:�Ku��s�}fgn�Eйh*����3�%��|;H�Ў�P"�"ȨK���-�dmâ]J+9{b������N;,�v�Xg���3�	�@Ƅh�[�����m?����L'�d�=���Ӟw�A*�+m�gu�wc�;,a���Qg��c�݈R��ywP�D��=y��G9�+q�C�'f�O��rB���L
�	�����W��AoV�&��U�g,��\BΝ�[we�T-�̽���>Ww�#)ڕ3��Ғδ��u��(��m ����9��j��<���{��f'�CP�\gs�J;i��r�l%Ҋ�3,Hۆtn=3����3�-'h��*'v��L/a	5�ԧ]��r��H�Pl�+I�(�y��fol&���v3�F4��9�)5�o���Sy�&���K�6=Nܣ5����:�5m�Yl����ؚ��d���K)5T5�D!vX�c�����?�!�Jʒ���q'S��QB��'�Ϻ�n��o6�-�/.��ut����,7Di�u3���
I]�/gm!�����r�0��35u�N8-�;���̵[EQ#�j�k�:3Xz�:�f�ry�Uh�]*"H��JDP�6�*� ����цa��@�@�>Ͽ=�����y��T� 5���&y��z��=Ɵ?�w�T�*h�f������_:�c���m_?tF"ץ���8i�O�@p�kf�J0�2Σ����~2�Ѧ��N��L�p�kp4*�:����"�˴ w�;(��0��`ث��:���q<�][	4��*��!�y��#�\����4�I͇��yr��&%Sj^���^���5��~�iA/�:�������eL.�R&������C�9M�g��Y4l;[���D�|h���:o��ʫy�<�gfөe����;���X�zW:5alS�h�R����o��(��hs*���]2i��L���%��i�f��@;ȱ&��D"�7�#��)�;@�N��c(trd���)��q��O>w�M+_Z(��&���Bv
$���<�\�VRSg�87/j-;��Nκ��I#*߄�ܸfO(���|�N�.��O!Ƅu�x��_�^� ���[6��.z#�-q���sAĪ�H~Ow'�e�4��|_8
�r�+Z΃b�@��]�������G0n�b�9�q�on����b��{I ��M�z�z�F��g��)���&��"�7�`UuU&�*s��niZR��vՖ�����G����}��#W��fTN��d8	�!�[]k����������?�ԕ�����L{Úo�'ԥ�S|^1���ڔ{�D�q�>@T�=�W	��&%��?��Y�xH�M�uŗ���̅�p�u�`v��O�To73Dy=�I��'V�w��Xn0����묞�����KfX��h*5�h�s�4�O���C��S��2}+$-qv���D�:q,�vV�����FέY�����q��ï:��A�����T�BO�V=�q՗!���o��%�65X�%[�w�@e��9�f��=
1q�:se^g���Z��lY|�m7�Cι[��x��W�co����HY9��-�g>��֨����m�9�%��ʏ[��cc|*ȵ�ڽ_?Xu��r�O*�l#�WQQ#
?/��;X\�D�͉f�n;��LvG��j����wv�7z��("O+l���sH6�ꁡ�h/ ��iD���w�.���Ө��K�!�qAP���M�]��fvH�G�4w}�'����u�����r�c�L���҄�8K9^�o�xz=�.=�)��ށK��5A"K�)g	x)�#�bi��;Ѵi����ަ�+X��R�Z���/����5'�j_N�u�6mb�͔r=�1�a�H�ΡF�>Yk%��1T�)J�ӏzhP!\��أ�����tF�!f�^�oi�D�ٻY]��W&���K~s�J�6��N�,�ǁJW���ڒ�x�j1�9ˊ導���
��CP�t&�-`�dsU��b��.Az�X��c�D)�2�3��yyy ��2�h��pu�n3��ƶXLRǹ���q�.�f���u�܈xx����-`TlP��4�>�-ES�q!�M���ř���ʃq�6��k�ض"zu*�8�6'D�8����{6�*}��˭gs��c��{��⍙�@T�k�n�+L�tH��%���;2�]�����[�����Q#W��0m 	�ᛩ\�C]�ίF�=�Ct��"o�Ĳ�l�![nH�]K|����8��3�-��CBK����%�����5���P���2�>a�W�G��e�-#6�*�@�(��kmʺ�x��]7x0��.�o430���"���{���Rpe_6����Ib�%���}�ksN�c�\��&j��mf�LC�j= ���Ƴ�ٱ��z��s��l�+��=~����<��R�5����o��/e�Ђ�u�؍r��!7r$�]m�諗�c�h�:�n��k�'B���u���Am�qk|�JvH�FڗG�R�*���wf�eLe0(IOJˣ��.�bږۈН�ng`�]��K��h�;�#,�\mZ�3�t�T��4�;x��+[�D��Q�&˘/wrݧ�[�t�
����s���3��^:�aX�!���΂W�&��^d�C�a���K�Z�3d+b�Idմ�{BW��3~mB'��k m�K6����NQ��5�B,���r��@p��m-�s;,N�{��BW�a��.�n�'o%gu`Cs]��!ʗo'ղ6&��M��b�m\Z- f^Z�7���YM��YБ�_L��i�Yy|;�"��1���E�	��nX�1t{���=ö����C����뷠���oQ�T���I@��-y3[�8�;貤0��,��عy/�^k��YA�([YwB�q`��Bعyb�0A!\��(uPt��eg!�� AE�6Mv�}�;M�@��&\L�v�)�6��T��ZA�.Z��|�-$�r���0a�L��]yimk�Հ���_.bt��%t�(�&w{e��.B�<�kc!J�E	σ�X �tw�V
xz�H��	�:�CU�v߹�󨌏p:�{["��u��o��IuE]�����r�vs{�Aaĉ�Yi���ܔ��=���=�8C�6��^hD��J#mDX�6�V΢��5&������.�4]��늂s�����~?���~?������g��'�Z����8��ukg�ѭ;4D՜E�<�:q��]X��u����D�ŵ�0Ny���~?���~�G��}s?l����v��ױ�h��4m��3�l�F6ͥ���5S��Wxn4f"*�5bƚ*ڌ��?_�����~����}f}~������ڜEv?{y�
��mxTuQ��tcc[&&�>�(H:�2@��`�$䐉�H$�����b���h�lV؉�m�[i+l���v�;�٢-~:�"�8��U���6���n��X�:
���5�i�"�4��Mlkf�O!:7s�֞�]�ULQ�kU�Ռ]�j�U[a��T�QA�[�H��
:�LA=[IT�j�&ڪ��y�8�UV΢�"�#Mwh�ڪj*�c:�t]���&������m1t}�A�v4�wtv���ڣ��:�⪥�"��Gm>Z�h�]�U$DEQ1�Ttjjc�Q;��rS��Eظ�vb�j;�*������Q�%۴6aG�#�=84y�5���%�RH79�[Kg&,es��3Ή��<H��2|��m���a���=� w:���f�@կ��3�*(�K���z��螯=^�X�vz��S{sX�V��oe�";ۭ,���)䌙��q/P$�!��Oo���1��M��9V[�����z K#��rG+�2-)�h2D�12fA�p�	c��Ƭ�Oi��#m�E�~��C�-vѺ��i�6ԋR"�MgϽϘ�����ܢ�C5��R]v��t_s�V6=�!�D�)x�:(�<�M�	�K:��C����N��Z�#Nou��V���*�e�b0;�����&q�	9{t���	{���5s��=&�J������~�x�.�bE��J�U��C9���_Bu�>��t�b�N�1�Uj�/��[�7����˲��[b�b[nݬ��|2��Ban���Y8��[6x��(���\sc���?��9���͐�)M&MS�&��)��\d��~��u��S��cRY��\�C��٪!�7sT�j��I(d�g���hZ��E@�{-�'m�07_�k|�K�	��n�X1�-9QrU�[B�+����.����$W����u�&qìd��DŖ�j�-�!9�x�c4�jB��D4��.���hͤ��'�9-�x��̲u﹫�(˩��Wa�d+#���-����WV�gö��΀�����ؾ�L�u�E���[c����L<�0,<| c����uwH\����Q��U�qV��T�܁F6��Sk١��[T��e�H���{w�c�v`ض�+g�C�N-��m��vR0�l�!o0�mI?�B�0��!��p3�En�!�죊�Z�&6Dxsr�,E���X�!�Q�&�ͨ��lî���m�tuaZ6���й|Y*�-ak���S�}0�ʵ�7C��CQ�W`�x�1�Mrو;F�2��Ѹ���'��_v`�xeؼo�����p���� %��a�:m�-\;��\ʜ�My|H�2�xp��ru��hIg42�ʖ��w�Dy�vX,�Z�1�oY���Yt��!��in�N�\�䄪D�.���h���<:]�ǁj5Цq<1�\1:�2�t��p+�3��~֢c? d�[����	�m\���Q�·r�\�����]v�Nξs�Q�,�~ZK�Q�Wo�1.�W��K��
����1��� ��Z��7&�pݗ�@@�I.��
�z0˘�ާ�8&�v5�#S�w��g�d�;�d����#v��ػ��+��9;=8Q����!�v��3��nEG( �I�C��/��F�� �`Ɲ�����\��&�3X՗;�p�:Cunue]���3D�=���I���N�iu�&��]	:�e^�Hy��]@B/myo6�?��0C0/�__[�Ҷa�6`'7���o�o)�V����y�g��2a�� :�{{Ը��OY��`[Ҹsul��ZB�{[�ձ�9:������1�F�c:��q�5�9Q���%`�h�lԚ	�_l�Ul���+���S�PK�9�G�F�c�5��F���ǚ�`|��f7��1���1Ki���&�DG��H���*ړ!���av��;�i���)��7<-t5i�!=_�7�e�^4O�7�Mj����Μ���ށS�܅J"u
s\a��-g��ZכK�d�+�7����-�p#l,��e�\W)&r��jDu�|bxe�_��w1a|d�#dn�dz��֣,Q,֥w8X�U:+�Z�_�Ks�ρ�E~2W�ۊ�.K���r���c��]3G��[֔U����`k�t��h�~Jb��>���iu�n*���3��JI		d�.6�rT�e>r�A �������~S����ۃ-G<ys����ڪǱ�̩gk�"_�ޮ\(��2@ldU��tH�*<�����Ȭ>�b��3����]�TвK+���0� E(±���v��T�M�bP�AD��p�7U��;���ԟ�&�B��9��Ƶo-��jMBF�`�sY��@�	�a1�wmm**�_PiΰԖ��|1��ʹ�L�u&�mԥ��������p0�NGG��~��_��{�����0����BX#0)��U��a=��P,�U9�O�{��ڊ�CF��3�z:6y�p�	�l*�%�7��X�3<�z*=�SQ������\�Uʵ�э��Z(����j��˺Wӕ�Z����R`�o2�S�qh��@�)�]�§]EbU�v��+-�зW^��Ζ�,rz�qV̥�3� �p�>�"�A�$UJC���DSN�6B�������>mxL��r�Gu(�z)l���o^w�]�����7=���j�M�@5�0^@h:�;ϼǚYA'ӳ�P���'_��SyE��6ΣV�u�*zދG��+Tx?1�%~l>�����W6���j7���M5Sj���1M�6_�XWR\���+S��B��q�vcT)�	�Yv�'O�>�����<�]��Z�qv&<`M�y�`.ې!�����#~���<��&|-:7YA�$���sy��ѓu�Z1�Kp�� �����F�3G�W����~�>+�Mv�gU.���/�nV[�a��kn�2;�uֱ��E({yL��F�2��i���t
���oA��mӮƬ��Ai��Zţo����~��^�1��\�ȬΫ�+n��G3{*�o>3����K]�6p�-�������zֳ|�����}����ן{���<�V��X`��T�{ď}���AU!d�u0��l?����
�>Ǜ5ܲ�B4�&�61D�r$k\��w���.?#�O��ހ=?V7����28�d�jl���1��;�bّ���Ќ�G]����-�S�N���"b�����kH��7�w>|ι8�?�\���/��y�7�%4�p�A�v�[I�'�����ҕ�Q�f&.����]X���˸c}πs�T�D�蹝p؄UW���&S��f���f-�օѳ{$�&��0�ᥫ��PV��?L�>*��%p���xH�5=�?U�k�x�*�:!�ZY����Hɜb+��&���v��0�#����B
�&��M��v1�|N�<i%s'���x̵��Lp������p�c��Y�/��Āg��K��~�C��� ���պ�j�yM��A�OT��r�vV�V�/�Y��J���{:���N�T���+�j5�H�P��rt{��D��rd#>Χ�JfR��isC�U��5�؁l>9'�6�M�)����K�J0ϛl�:8�l�JF��:�lvE*��ܫl&+z��b��m��2Le+������]��dU9ɘ`B希�W����ya�@9Ź��@q�Y;�����җS��5A7{/��o��9� �\�9n�:8+]E��!+�r�}s�s��+]m�Jc��9���˟�[w�:��0�0¹H �|<O��EWC[��;:3���9�N�{!�O�kT�'�[J1=�C��vcn����?rk��sN=�����|�3hom�x�д����@t݉�ۧ�ǧ�9ו9a�7I\N+�]&Uަ/���wsd.�]�/����}=Ե��S��jH0d���G��ʱ_��Wr��G6J�t�]Lwj-�u�n��y|.Z��r��N�a;(3B���l&A�.���Y�5[+�t>u��¡�$�cZ��H�nL+{ Q��[���y�۳�C9�!�u�!�G'��3-�8N�0��F���P�t�������Nj�w���\�Q���.=�~N7��sJ�M�&���4��QNM�U)��:0��>�S�E��x������ƌ�� ��aĠ�)��g���t�|��?��4Վ�n�߈�h��so&r+f�7�n������I~�\f�2��7��"֡N�T��:�BO,m����G6q\9�^�g�v����x���OL�sK!"r2��,��
\�jCcJMOFjqы>m��9L�Ve�@_�aq�V��"�}.��n�8��ǧ����3oꏱ�Y�P�i����E��UQ`3�i(�Y�c���@ݴ���W|�Ytw5�Ԝ+�ø�k�VP�p�[+��w	D�]W�t�9ۻXL"�R�����B\w���ǟ����Ɠ���$z��K.<�\V�y`Y�Gs����h����y�E[�<�"���	T���)�$Ȯ�fO����l
J� ��:�^����}���<Bjq�ڞ��+����mekJm�W#98L%�Rӝ��Uy��n39�B��޺d{�bx�/@��h#9	V��La�`F�G&ğ�w52g��׉�:'�nxf-�P 0�@T=)������e����<�/��X�'�d�.��V�#UI��u��w8y���	����vԋmi�l"XJKt2=j7�A�S�j42[�fG9�~r�"��"���j�"3f�k�GR�㜝ct�\��ΨHc:n7bJ��݂��9��I�V[Y
́�z���Z�>�Ӆ,g�+��3�X��J&�cv�F�ba��#��l],8�;���6�{,R�8�y���:i���-'��{)\޼�c��0��9qŪ	�)H�lW�f��sf�wk�t�6G������▁:�q�ב�e�w�M�oej�r�c�|c�j �(��M���B�^h��WQ�Of߹���\�=6��R��&�`b��a�l��Ĵl�P��j����v7c��Q^����[ޕr	8�VǕ��RM�Pb��:�+�X�a�Ӗf;uT��s��"�ൻɭ.4��؎�Wb}ʸ�j]Xz��[s��ܧ����Rǡ��s����W��
�>�=���gi����5��@�;>�֧��˹����TG���B��BOkꗇv��+8Z�i�Ez�g(x��^y�q���*�q<�v�g-l�����@g~z�#Xiހt�ɚ�	Mr7���}�*�cvڙ{[y��B��$��Q_�"t�(b����n���"Y}�E�����Ĉ��o^�	�e�s�y�:���3��DS�h���f�S.��QnQZ�����Q~)�����P��jE=�j<�M��^@ހ�H�"m�Tv�R�fbvdN4����vd�%%����([�F �%��x����s����j�r2�"��k.Y�9��Q��K�Z��{>��3]p̞Q7��L�J�i��kL�oC�M�eH�e�Ҁ�w�8F�Y\B�{/�d�kM��!�'���	�[���3	Ψa�dY�5���U�ӭ[����u��zCr�dX�z}/^�dBP��%mR�9=�n�x�.�O:lE�n�I��-�j�yy�:;!Y��=v�C[-`w���9�)���N��
���7@܋>������y��nb!7r��v�E��&��*Z��0.6}��i�� �2J�[�b&�i�?؜/���y���2��K@Jm͐��[�;�7�w�V _Pq��!�)����a�ŒpV�6��ͽ�q s"���7��{�w/�xw��1�q��ʀ&��]�{�N&�7>���f3��VLS7Z���J7�E�E��x��V0~������%�|G\lkT�I�Yt�&O#D����x��F���u�����\&�b�l��Gk����:z����v�x4�t&L݉��=���s���k���1��hn�)p�����)l�	����':nV�F��F)������N�1���>�.��0~��n���]z������<.��%휳�����\qB���g`VwU�quu*8�V���h�V��םQ����̫[�n\j�dV\�F9Tz��:ዽR"Q�!s�&����fϱ0�y�����Ct�Xg��A�ؘ5sv��V�,���g-(�c#WOGUz��j�������9[�v6�tm��3��4vR$Q��p˺��bqEOH�LEk���4���U���l�6��	�7�.sK��m&��3���Dg(fk�	N�e$���L$�!z�k�r:]�7EX]���l��
�㜟Wji��%f��E�>O���@n�9�t��2����g�K��1�r�l̽n���-q\���͆pFDz�o9�𜕭��Ns8��K�M^K�"�;![w��
�ڲ�M�3�n�]�sHф�4+���G�!>B���3a�!��Ek���I��i+��6��y�L{#�k@J�?�ˊMs�+#�����n�����1�/9�;K*kݏB+Z5<���q&`rSi���b�i�mϑ����	��mg�z�5���q�(% �f8��]帵� p6�� Z{�qB�k��yn%Mg�ۣ���΢�j���mw�ښ�t}�O�r��|��79M�)���64���G���4����5�؝���긫�k��HaC/���E�F3	����رւ�ǌ	݆1����eRUFH��Q�{*'��K�{�ZCcY���ZH�y	0��l�:��!��d�֕o��%l�>�j�d,���W/�履#��E��53�GĞTB�x��.aִaM�^��f��*��B�ޛ��������<�g������(^�ҷ�M�r�c�RY�E_f�J�1|v�á������΁C1�DO��Y��goX4����B^kv򘭻}��W��bȝ`VBE��p�J�^�]�v�3뇼m���W�1�qk�3�a)��"qV(
��@�uo8�MS��n��n��}��=���� �����_u>����5x�Š`�hs��T�E��Υ��!u��q+�N&�k�=�;J�WTHVDٶFN���<�o0݇E,���'�gy8yO����JI�G�r]С{u��m�ťf���K��{z�-�]�nu[tx��v�PyZ*S�L�}�2]�m�-��N�j�gq�ڂ�8���J��HrR�Q�&[�5:vM����	�r�ff�_B��]-���[uԭ^�n���Q<m-�K7�ie��(�+����.j�����ٙ�y��i�Ş�u��X��<Ԙ�j��;3x���fP�r�l�U��b}��-D+��B��h�*f^�������4u�
���f]�	�vö��Gyc`hђN��xl��͈2�,�����ooR��
�:�w�m��kQ��zmZ�_��-���m��@ܡy��݋u���e���m/�'y�q�p�q� �_E�k�pW}u2H�.����3L����b�
��1DV	�f�����h�y�Vh�fJWB�|�-��늡B󁣙&]:��"�A��`�VE!{�)������WH����T�v⭱���&S�@�Kb�dHX����U�l5g+6�`�I���ӌu[ɽmV��tl�7�<U��=u�3{x	΃��pB��;��D�y_O�o9	ۉ�j9��Y�&Ωk��1K��}
X�13�asV��$�n`�f���W�\�,w+��!��f��8V[�1 �VvvҐ�z�Y��=�-�MZu��l;�ba��c2dR�<�1Xb���L�C�H$ճ����Q��t�JoAy�s��DI|zL�4C[�&-�6�e�b>���_�)�m�{���ۨ%��c:�k�(�u��t\6on�)};{�t��'+��H�$Rv���1�����d��_c���C%%n�F�z��z�GR#u!��:���z�*�z��#7j[�����x��{��Q�!ޮ/�]sC!V�����kGŻx,J��A<&w�i-.�J%/�������bm�8��܂7��ru� K}]:e��+O�ɻJ����]�ym�7MQV6�?L��9ӝb�;�rp�]Ά\��,\���V�!��1h�7�6٫���r�V*�q����Ww��k4N�-=�[�2h1��h;�̡�{�³w#�)QN���t3qv3��ܢ"�ʌ��&N�Ց"�]uZA�%��;&�D'{��uM���T��w��{������\RY�֩ �Szw#�m�>�aX��H�y'F� �\��P�E�)5���P`�إIQ�+e�
�.�&5mP�. �L� �QH�M�&�a�l�d�!�Hv�M*D�/8P 
�d�DG���b>[�+�]�E�A���(�v��;�MӪ��ݫQQ!�����~?���>���3��ϧ�E4{i���Y���{�Z5Gٱ]���ѭ��6�M��t�)�g<�������_G�����g������SQ{����l�u��Nت���A��[]wF���qPN|}|||||_��Y�_���M�2EE킚�h��֭�i�
.�Q$q������Vڋ�=X�=:������N�E��FƢz�A,DMTI���*�����/+i�c`�]�lbj")j��Z*���N�	�"���������*"��TRѠɳ�7QA���}ڨ���>mAEy�[�����li֝�*�b�bjo�����:o2k�LI�ؚ ���](���>v��H�����h����Zؐ�����"<����m�E�h,AWc]w}_�v�^c�l�� P����n����/���͍��t�.Ե�]�u>���^�aQST��;��hL��z���H� �ü�/:��xU�uU���5��>#���9�K��%�1��a�O"���ph��S��. t�d�O4x��fua��i�^"�D��
�oR�h�
Ψ�<�E�ivlX�O�)11d@��k�j���6��㡯��۱6�Uo��w_�Ƒ����H;�캱�o�� ���uÆ��V����]�L�(FL@j�ʍ���
�S���������}X�h)�=;� ��fmO^�p��j^�E�����Om$O����(V�x�D\���)Ĉm��)�	�4	��S������<"���dZ옆!�	Q=l}�kUˬ��k����/J�s�D�*�h(��2�־hM�-\����j��y��nr�a+�%Ȋ�c� �z��%��-�,Ƣ�:*��ճ�cs�->����j���Sϳ��^ΡV��������A��p0\{)��S�	[|2���xǧ5ݻ��f�t�%6Q�.��y��4zBQG��ҏdJ롕p�L'	I`q�P`=�/�q�:�ſ0�j�3_T�2��,��6�x�O�=ŵjv�W؛�w/�BCv�$V4�p�oOZ:������T�Jp�3ݫ{t��r��������1�4��0�a���s�n����ϰ��_wj��p*©����q�v�!����N1�n����pUn���ۂ���(]�N�ƻ�'.�8�9*jV���� �xS�	���>��W� �<��Wh���w�!�md����XOu)�).�+�c���K��q�m�b&�N��W�o��HQ(���RDA�Djn�K�\U����7�u�nM��qhB�!r\nu�x���c��M,4IͶp�'$����-	�CAP�}�B2.��>���1��׋��.�8�l��,���m�7��0��lTs3��%������u��󝗱�إln8l��|FIAg�]ށ
=Jb2na%E�\���.�gfV2z}�u�G���S�d���`{P̩ר�u9�2饴�[J�CU�z(S4�B�6�W� cǨG�R=fY^�Κh
t咟=�Õ$���W��G�W3�E
}q �`���#b�̴�:�l�i�5��ލw��ensR*��zvbgR��b�oG�o;ddj���g+쟮~e�����l���	w�1�с�&=��5�ɔ0qW���<\R���?��݅D֜|��K������q�G�з�/�
&�w(U��(���S��kk^���J�j��tx��6od��`-簔Ŧ�ȉ�,�^�"9pvvq��X.��r�8����kw
�XU�RȸM$���{�b8��3�^�Y��D�����%��YfĂ	�;5��K{��R�:���v�%�U��غ��^>)�J�(u��㺪�FD���U$ꊂ�'k_F��>F��aUJ���s��}��}�9J�\��Q�M��;�"���g�}�q$�R|�����xfJ��;�h���vbI^��~֫�5oxYG+;[��li5=��<OA��2y�:���Z���v����{)�f�X$���q�ˑ0���VƌF�ml��p�א�q�<��l�����a��л�ݩ]2iB+��6	�ː�<�z<����0��7�sS�2�qSf����xm&���1�}Vv��4�K�K$3)��8i��e��x�љ��vvO�Y�^���r<���:�����CCx��9�e�Ӽ�MM��:m�����l�pëe���9�ִ����u�-8[O!.�v��!3�h ����!��E�d����7k!�&R���u�p� �/����Xn�Yڹ�e�$���!q�T��Ô���:����t����w�X�\��m���\;�V�����N���V!P���f�>J����[{�]w���a�o'�fcaI,؟5)}�5s����ս���O���3˖:�n��ϹO�֜^w����}�U��/6����Y�~�h$>c�H4Q)fzDp�
�[�T�)��=����|mS�N8�v�o3����h�\+v��9�=>J$tǷx\o<Ū*�fv���"^���x�;�FĺG���OO/��!�{���^Ô�ꋔ�)e/Dg�)=�
���b{	xx[G^�s^<��e�]�}>�V��e�?WWr�UOc�5'齌�m��wU�c�F���)��tW�B��W���]rY��]5%��fq�מ�OE^�4�;��יf<]�HӁ�eW�N��Oj�9�:�|��M�s�E�D��6J|��[�K!�f����s�Qg�j��ke�նp��&����K����4ڕn8�n���vom�ͭD甬�ys�CkV�u�l٦�����Zf�6�M�;�[[��ʗ�h�ڂ�P�#�=�B��R��R�0Q��4���AARQ��c�黻S��<��n�g�ywgm���ϱ4����4���<�LI^�Իޓ(��4G�J�_�3gE`*J�ӧI7F�>�cwtcU����y�7�?�	�F���'F�d���m�h``�|6�N�gu����wz��
�����`UfԲ�:O�-��w�Ɋ�o���=}��j�?�is���b���-�1��`��=�/�����"v�@Ԉ�Ի�4�|�9��?�M��?\���=�}0-)-60�T���������0 ��\d�`�butX�T^��1��P�L�N	��g�k
����;���.q�֤w�T��Ä��gjCŬ��b��͖��w�r�:oN�R���#�s ʺ�+V���+�&�1�{����/��q������ �	~�����\�8O�3^�M!�����C⚇�gx����<j��(���е�f��"�a/�R��sV�hFv8��CH��x}�w���4kQ�D�;�;D�&�t��~�P_1!<�Ot>���*�[إ~(߻{
@w�neY�u�PDy�=`,�Ҟ=u˶��*���ɫOڣjgf�Q��o�,��3���2���5v�}��c�.�0̜�35����[����� =v��� ���ܪ֝L'��������|����m����喬M��A����F�k�3֫]�T#*�81}W��I=�1�ha>��j�SP�*���n�VwcƩ�h�\�xe���8w"v��%�m��|}�^���ո�VM+��Mh�o^��c��A��vk�q~yݯ�R�� c:R;a^w,�J��~�xه���9N]!N�L&�2�؛^D�_4������9�d��p���K�g�9X��*
]�%��C]>k�^j7H<�ٷ�eE�=�ѻ+]˓v�Z���ٌ���uѴ����؇�٣̴87j�ٹk�{pJ7/zjWofRY(Hl��0�5+�ߧ2j̛S�b�&3w�sM� ��J�Y���v� ���X��.J��/�D̺�R�=�|H�0�|�&q�}�B�s�7�˻F�dφe%�ޭ�i���s��Vﭳ��*�WY�S�w;���5�ۣ`\�����S�����BWqp���6�J��K�nv3��-#������˭Ǳ�?g���{ȄJ�o�����w��ֱj:+u�[U۹ՙ����K.��xƖ|��|�mB�3��5�w�w�\0ܸ�s�D�9']���].�BT;i�}]cۮ�Bz�Fh��{��M�t���4�8i�y�&J�ͼ9��V��<�+��о��c �q��!�{(�|�s:J+����T����!��i���{~R�	�����ϸ�˧7md�AZ��y��M/�ِ���������(ʗ3���UlS�E�GZkW��F류�I��iCU�=�i�od������S����vn
�٫s�"�D��r5�[j7�d�w[��Z�ٻ��{ZY�#Y�ꎦV�Z���W<\�ط}�M�L�+��~Y\�l��\wU)�mp*ʈ5�7KGn��w+J�>(��������o'���ߌ���؉n�;�Oөg$���:����e���&�`�ʔ���l���;
�y-ܖl�"^�{>�mD�]�o�Q����ulO��W��<������<@�Z��9h˥O&�6�=��xe��{�_Og��ێ�;f�wY�!�Vy�wo��%7ViЬ��3mK�3�i��v�n�AgT6\�i��s:U��f���Vl���)�~ݘ{�]J1����;{�^�G�%�s]�Yƕ���b\�yV"3%�1�&�Q�f�_p�vp�>���2�Zoen��*�SL�'U�5%�rp��.���k��X�Ԅ��a�A�#�l
�e�wĚ��7l�ݑ�����	������Ǣik�����i��g��Ylg�͢1�^x��O�fv��W-�W$�?$�mV|�sr�k��s�7�7G{=�LD4��S��3:${4��=�6�T�)*�!{Yf5�olbqR_�b��^nBQ.;�e�B�⼲1�go@�Z�e���m��wha��nUh�|�ؽƖ���P���yߕ�!�Թ��dP�*��E�#875�l���g����Vǔ6j$���n��z��Q��Q����D-|���vjԧx&\�_p0-QQ����u4�<�++�{����u�y�uJ�^�N��3HoW�ե7���u�@g�Oݘ�e��W�J��̦�Esw�q�j���f�S�����r���쯧��?)�=��r$���f��uAGfɮ�����1ޗ�@�I\�������mvoT�(;�����鏇��k����+��wA��ۭ�;�sN��u �n�Nk���S|*"�jt���&�S��d���X��G���Qnӛu��b*;[�U�`m���F<��x|<���5��D]�����G�o٨��B�ڻZѮ��KvIzr�Wg0��^�o��7iS�z˹�ޕ���n�4<h�uԪ8�X�`^���kw��vb���7l-�^��ީ��Q#6��X�gm?`0�U��4@�_n�@�w[�����xް�����IXm����c7��l{�etCU��h׎�n���~��
͍��f,�����.�i/���4qt��x�����~��fY�#XM��@�X�t��u=���Sh�j�0f�ܿU<�8���~�la�X�G�u�W�otng��iT�7:�u���i�nlV�����;�~�d�_x��5��F8��X��i��PԱR����vsYE�A"��DfuCd��p��V�[�ʽ���V(R�[�g[5H&���<�������>�T�'H��:兎w
�V"y¢��V�j%�ml�]]���0�Q�~��s{�#$ܳL�+Fl����G_���WY��^��RU�G|U,PL�dv(u��6��ܯn�z����û��C��j�Ի��j,���]m��^Ԧ��k�"��M._ �3���YA�5Y̷���<��-l�S������5�{��.�h�~�H�vT1E�����]�!�����{�ۍ����0&�Ȫ�)�\еg�KꊜVK�RŔ*6�&�_G{��]����W��j��3�������/H��y���ݩ��TH�
g�yw͢��g�<&g�^�x��I�Ͳ���ܫr],u�=�[/{{���wWU��������ӷu@\%_��"��c����M������w,�q
r�u�@�="�^+��%��`4P��>g�MyQ��H:(��9�e##��k%���r���_��=:�*����9-��~|�c����O'к=]+�ޥ n�oSs��Jj��UƮ�!ֲ���*Du�1��f�N0v��sc���.q5ۺ����J�ݵ��P+�L��ձ���sq�g�+Tly۽��_r�K���e���gw�2^JTH9Ȍ���mu;(��N$J0Ca�c�o*L͹�NC�q;�Mu�3�+c9B`��f�z��e�z�w6���ږ��U�gJԋ̬C��`;VF���ɜu���d|�;8o���Z�������7z�F�VV���_�L��vB%�]>� �	���}�Z�({�KB㮉S�s���٬��9mTu�T�"n�qn���}��B��� [�v�qֻ�t��ctxq���
ܺ0mѵ���b��K��΋T���J���Gr��}@@Ɋ�7��r�i����ߊQT��c�o��yʵ˒;6wchYܱ��>������)���:�K
�
�QȜ���3��j��ʙ��u�7�ow��F:%^4���C��1#0�i1��3��͹�i�]󫋘sP(��hk�,���>ǆVI�]�Bz(��Wh���ga�͸le�M�������G���8�>����4ݪ�6�R{g�m ���ɔz9�5���6�-N[t����[�O"n��h�0���a�N�򇨍�a��Ht�윯c�5�2�^�u�qX͉"�Qj�i@:��6����.Z�����k%6Q����O�k0�O����N��ky�PN�`{B�,J��IXnwp�����eμ���S��it�N�%���q݋�kJ�=��t��/�����]uf��a�=b�X���Z]�-�Z����4u�0�C	ʶ��]�n�a�7e��'�Pjy��t�C�㜍b���t��4{Ris�V�Po���7W�� �]@���n������Y\v[k�k�/Li��͏�n�40��w�|Fˬڔ��F�I��vA��t8�b���o\�;��)T���S1�"^�Wp:�":�r��Sv�����=Z�V��-������0�
o�^L:%⥀J����AD���4��0�����]�AVFA��,[)�:��ް�j�v��b��.�]�:�k�B�nnڎ��l��a�e�Z�B�V��kWj�x��gT��j���i����[]�2�Ex�)��39q�KV�&4�t�䵢���eӏi��
.B���7xZj1BH��)�rNuoM�`��%��Uj+:�H.�y���P���ok�%�s�[bS�φ�OSu�B�J�5�΁
�d@ǫs���5�p</���]x�ך�vd�x�`m���h.M!���t3]��8�H)Y����9���6�ƥ�1�D�[�����I��L[E�M�g3U`��x�j\�Uk`�gh׭�c���k��IoC:�b�;L-L�K��gs�;Pjy-[4�Eل֌ᒣق�LIg.xe��a��T
��kq��T1n�*�#�y�����4l�7%̺��N�yR�纺p5*ٽdֽW��ڸZ��Z�� Δ�
c�vn�^�G�Yw5r*�r�S��x��Y�-�uݬ��c�������X
)$CY���ݢb킩��8
"��������	�J"�矧�����������ϯ�OX���C{�E��CTMUQ:��A��6�֒6�9��������}}_�g��?���"��j�����5���AT��P4W��l�_�����f}~3��'�EUT[j �`5���"j��6���*���Q~�D��% �M]�u���[Zo��St�"�i�z5D@Ql�b�MV��MMT%-i�	�i
B�����B`��I��'Z(��"��cD�	uE�����U������h)bh<�Ey:+��Z���m.�h��gA�-�i	��c@CRPU�j��"�����"����Rh|�LM��f*����*�����%}��ݪZ�����6���clj��6��W�]��`�G��x������}O�t��p���*�`�}wW^Y�������/�Q-X��be����^��^��b�_/��{g
�k�C��.T�|O�L,��0z�\^!��WJ��p���̳1��ٶ�5K��k����Jelsڳ�ǣ���l^ڇ}v�#�Z�����p7rY��z������b��W'�P_Ƌ�詢3Ѣ�+/���v�����a5�X��߯�O�38P{��2�uf`�:�Z�ݷ�mq"_%��*�r���!��E�y�"}���k���2b����ByXu� x������{|�bg��⪱<�띬���[2;�^��:j`y��3��!�t�e�iq[9
���p�qc,�ז��<��Ue������LKi��TL-�ڭ�����x9�G�l��f}���\�u_��Wsj��	2" d��B;_'
U�Q��sb*6�{=o�6� k��:���]2�uw�p��㌴��v\>�ś�)�3Q���[��;,Fุ
v�<�ppĒ��y;%T`�,�������"��xB;�=d��\SX5o���>�Mk��_kVve��gvZ��|�?����r��}id3�&�-[+*V��_��4��q�;�K�E:YՖe"7)g��-�r�|�R��˶4;3����.�0��տU1�O�A��YP��K䥣�p�*Q5lF-tK:d��3�s�e�:�H%�й���Z����L�[ǩ��I�E-ج\���⊬������e�+^�������*��d���l�z��O�;,��-�	�ͼU��
[t��ۣ\/�#)s�庮�ɀ�"���C�]gowuX&e���{S�S��` :b)�ȼUVݵ�;���f�����jh�j�J�C�v<��S��w��"�]�\�Z�nnVը�wRb�@m��;��Ѱ��,��;����Ԙ.w���_`���-ִ�|��[=b�]u	�󄝐e��5\���U�ƀ�9�E���2��>�R,_:�n+�.�1��'������,�Q��3���,cK=��g�3�{P��zW���z��Z�b�I��R6�q�Ð�Ϛռ�.���s�Z�a5�6��]`x���m���=�]��N��cT��$�
%��T�rz��E�K�9�R4�W��ܳ�B 
�x��ft<�֮[�Nu�v8�cu�tU��SN�˸�o'xV�Q���z8zh�,� �4�iP�Z,R��<}�=�q���o��A�� Q���'�g<�@Jظ�-������L�^�:k�����gT��,��o:�e��ѩ�o
�O��J�ؔ�F	k�E�K�(wy���Y:.�/�Z���z��J`	�����Y)T\�ydȺ5p�uCX���;�-�7�	 �Aw���`zʯ���5�q�V��r�������m1[<�̀
Κ��^P+Cy�խ��t|��=̮�lZ�DuԼk����ٮ�J���̑S�|��@?��:"���]E���>��������3��N��jא����������3�qL�"^x�F�%�7'Z��]��7��ٸ���w ���n8��Yd,���K�V-�z.�9��j`'7�����yD	�ͧ�%[��#ܨ�h�/:���ȹ�����O��;�y*��y�T�a�����w2�v��A󙖞\8Z��Ox� ��Q�Ў�eV��1���իio6	F ��=�c,�W����>|/c��QE`�w�e��1�
��܃,�z�We��٣9�
���[�ۇ6����}��=�U��k�ѫ<�v�&@�r��z�3��D\j���M��wMɮB���琂����M�vλ�6nu��\�+P����S�|����l�Z�3��L�	�����~�ɝ���n\U>�㺿=of��{o������Z������b0�8�b^:��y��}F5I�swX�5���Y�K��5GiR�u�(��\�A(�xǋ����o#n���I�5O��L�����Co�)jj ��)�ɝoPG��1ݺgfj�Rեy�ٸ�!�ndUnǮ�Ot�O��y���Y8!����L�"rȚܗ%�����;pc�yI���0���"y[���|C�~ v��;��Bq���K�
Y��L��VeX��>��|��q��t��>�ћ�-tZ�ϫ��z��QVV��|�;�K�56B*I����
����u���^�䏷z�d�oJ�i!�$��[./}����+����wN�K��sm".�G,V�f�w.��S���ƎR�#W궫}걚��zg;)}�d����;=/���c{��'m[�;s�=��]�l~�F���u�vu��,:��哝��܍	:؋����-m}�;�ުu�%�>���ޑ[2��Ǆ��-�&b��*ww84�({}����Ht7`W7���jY��.VB�.��z"K��aO���2��]��s��XͿ8���P7eV$��B`�ne�s;}�3~����)4]��l;c�%����:ҭ��Ex���0�|�Sr��(�%U�'pTx���������e�Dّ~��o]_37',�g��f4Lӝ�;�M�Kږ\��MH��3i�{��x�7�Ӛ�.un��Ui�.�cĞ�1��\i-�'Ƕ�n׿9�L׽��
�Pcڎ(f2��p�g�uL�۹3�-��WJ�p�V���*��l���׵8]|���r�����m|�L]�u�7i����m�$MUQ�ݷ��;����q�d�^ї�{��E��-h'8�K�ݼ���B ���a�Qn/���~�F���"���\t��x֍�1�Rr�t3�������@7���X�m��2��gR��˘�kM:tE0��r9]�X���s��CA�hʋ���*�m9�}�	���q�A���W$h�{��-X��]y�������6X�͖Q}���ז|pT;JP�&#˨k�w=2b$�*g���M�Ɵb쁽Q�1Y�t��ƸS��;��T��P��#ٴ��#n_cdA��+��~m��|{'�\�R�UG�`Z�j@�	�����2�"[zw�J�=�(n�Z�+zuҹ�	J�j3�e_+�Y��	z�
Yl��g\^��蒷s/CJ��z�@�԰R�itP/z�dJ��R�v��F��(�h̞���X��m�IopW>�׭���`�ْsH��K[`׫*���l$�gι�v�CW<2����~�B͗I�r�gR�4'-��ޡq��w�Ǘ�my�1�[{�y����o����;a/˝�ݽ^�i��w5�IRܳ����&����p�#�B��6]Vm�|�v�i*Խ��}~��Ͳ�Gf���a��/�����,��Gr�\2*�-����SwQt77���+{zg5F��.��6�;ek�C�Ȫ�sPb �l
��A"Kee���O>՛�)�Z�x@��}ʄ�cZ�jp����^�=ؙ�����c���h�<��X�i�2`Y�6�75�0�3G��钕���D�D2i���%-��Il���,�[��6�Ô�c�����L+��./U�nTmcTy�ן�wW���/�Q5��p+�]��0"��}�逯���I�^�֖�ફ��c�ݣ'w6s.������.z�*���5 FO�����
LnX�6���bYv�6�u��08#�TsK(�9�g���,����|]s^zk�h�݃�2�[��}��9
��H)�P�/�YV����c�O;#�ll�.��\L������go�@S)��q7�4�\{��ԕz����5�X�'���*�Tq�^��4��-�*��`��Z���V!�k�d�Qs�W���yT*��}����{s��O�=��۪f��cۉd�]�t�ϝєdq���"�/*�^H(���Q�*�>]pu�i�8^�
׻�t���6�vls��%��mM�C��;ӊ�[^K�=�<�Hv��jk�+B�#�z���Ec�t�AY�q�,v'v�F�F�d�|^p$*�A��,���	ݚFar�zU�Vԝ9R��S�]�8NS���jG�i3ݯy۴1�Y����5J���y>��LL���r���c���x:==|�L9v_h��@ޭ��x�[�m%ãЮ�v����묝�m�,Z�/1��R��=)crx\	��2m��u�c���1�o�;������T��7ڏ��zr�'scjR���%�N���[������sM�ְ���!Fǝ�t�{f��WW($�{\�J��bUl��ۤ��P�m��R޼6#X��py(�} \'��|�ck�T�+�f��]�.k�������qo�\h�9�$��v�{RƋFJE����[�m�����:���v����58Y�����t�j�� �(*���Z� M���/z�f���7�[�[-��7��ط��+!���w��B�j�ѵ�)
�3}U٣c��|)��Y�{Z/&Lwf�x��ox&�'؛��A�L����)�u?�o�d����[I���.jne�l�`jͰ���;<҇|9�׳�_e'�V����v���lh4�g�uE�>}\��;Z����gT�24��H��0{;\��������f�5f��>X�3���;�v+���I�:�<-N(�y����:Q/v6��!w��61��V�)oG�� >��c�����Wӿ���(���O������=�}��z��%�,�|,Y�ת�b�uݝ��{o�fR��%P2+��U��S��=�ށ/i<.S���Wz�,�;~��}��� J�]&bO9��"m��޿LSs5x̚��jW�ϬΫ�y��7�vX8��ݙ+v���.�m���͖&U^N�q����������q�I���u{Z,�ef��`�v�ת�Z(��6�e�Nul�{�oh�Ǘ]����Ҷ�j��n�z��]�Vn�ʉ�݊=}X7���a<����%te�[�;�&i�湜�����j�O�S��g�c�qlB�72����̈#׊"���zZ%�P����,���bz�-��}O��A��tq$����%u͗�0���l(d��G�A�5�0Of��w�ռ��WW�z3E
�Ǜ�i%^3��hv�ՌB�]:����]��ǽV��A���T�a�BTh���R�K�<�w�o�K��8;�\�m�un��X桚��z��-W��~���]p{��y���K�}y�����۞�`�FI���{�+�{R��5=�;Ə������*^�Nުg�nP�-�`�ek��dX�{sR��n��RD?�Z聗*��\�uk��+ϵ���g��_�������J+V�m��� ,�F�7@�8�-N���ϗ,9՗�=�'5���_E��÷ˡ��C#xw�¸E��.qnkJ���������\��l�S�z6���w�m\��TZ۩�J��p�	fY̯��^��k	��hm�Y+i8�^�Z'�-oD�J��Y o+UC �k�H�P�^���d�y�.�xUS�ۥ����ח���2��k).��oo�8����1xk�ZGK�X��ݺn*�U�i�M�Lk���Ц��d��RR�j*V�xWe���4匬��] n�T��T���B��U�hKPk�7s`Ҥ6�_�a�4��nu��/��'5Pm��0h���`��C�+�T���)��+�ZڻE��O�ڄjiJ��]��m���A�+�l��!�{ӷ�-�)�@퇮%u�۴�o:5�:��ʷy�WC�!C��h`���+��ef(�(m�]fb�X�PL�i3����J���g8c���G�}��s����8\���ot�)� ���v��)%*�e���&u;�N����U���RB&i�����Q֎������m"O\7\6*�P�W)�]��AW<9K�t����B;��j�b_Q�ke]w�e����n�lQd����8@��U�vv�VkU���69jHyu�%��e�wմ�u�#�#�7ٵ��ĴҜ9��XZ-�U��Y���$)�����O�/x��y��6F�h��NV���i]ͳ�@!���٩�Z�>�λU��ۥ�3�(�jñ�{Y\z\��������8��5nm*��X|���2�#��(^ޠCs�/��m���BP�EsY��3�s��/�p��`ıQ�l
��t_���U�Z]ρd*���:;�vgwB5�kxӡ=��s���֐=8�棔��]��ު��RG���i���^i����,]s�G��^��b�{�� 9�ӛ���)ů���ҝ�^�gf<U�H��mYGJ�'�ᇂM"�)�1�;�U?J&a�f��w��e���^�qBEp��a��@���i��8+�v�T��_�WBz�Vm|�(e$H#��DH�D�c�X�[�`��˞�2��4U��4�G�����[��Q=c�;o^���4�)�{^;�M�ˤ�.�����k�&ٺ�����;(=�u�nr��v٣�wPfRA�#��C���+:hp�����%�Ql��2Pw�I��yuV�76eJ���uYt����Ԕ-h��s���iR������vx��1��ѳC���gq�PZ��,eb�\ھ}�铦{GZ��޸�e�'�F\���|%�Xn��y�SR%.$�;z�1|��j,�y�\�$6�T�twL�����-pcs�7�A8c�4��<}R�5Gp�Y'
�ܯ��`j��9-�Mf�c��E�dn���J��r^��+r���Z��F
�6�.>"9պ�	�������LZ�Hmh
n9��J|��h��·�`8ɗMv��ll���Y9^SLf��}dk���<��n����e�00:#�0�c$P�e'l�\r ����EzAݵ�v=�"��+zEF�B��a4z�W*q���v�N�޾͵���i�!Ҥ��q��f�m��^d�Б�z���oYS}*7]"N�����^�$;Օ9j�h��ؽޗ����u�/��v��X}#�JKQ�4 FeOd#f�#�?9�5i:����4<�T�j����ea�I�5LU�LQ ����;.S�*�:��[
 ^ <��ׇ�_����h�����+l�b�����H���/>�x@RQT@O?�������}}��f}~3�^�ݢ)��t�b�h�j�Ju�:�ݠ�a����������>����Ϗ���{'�D�ZMyhk�7�-P�Q@U4���t<M�ns�}}|||||~����������bb��Th��A�{�C6�UUU�n�D�KIGN��(��N���
<����hѼ���&��4y4��o2k�m�#TbhiҺ(�:���GGZ6���A�����*�����:꺠�Z�q�y�և����;����R�4M�4���|'OZv���O%.�WQ���*��4D|�M'�:ꅉ�y)��i��b
�C�����
j�ӣ�{�������|��\�q��;���[��k&d�Ax:m��dvw`Kg.7�xI1�[�v4��<��{y1���ƈɸw�O��$�ɪ*� �4Ax����1���:��]�]�|���Gәk����sg���qey�c�n��Vģ$����h�WOlGS�^�Y�>�+��۽�[�v���lڗ�2BۚV]@�Y<��wy���q����Tll�N����*//|tY�uDeRj}Y7�0��/�kS�����V;��\\�����^���i���,�$߱�2��s=��B�v9n!O��6��W�������2��z�;q6i�p�	�t�N`Ψ�6�D�ש�Mk�*����j��h�cȚ��b�'��MUz�Fap�q�"O����_�E�l��b�+�}9Γ@����^\[�ت�ʾ̻�����,�c�P�n�f��@ݽ�8�F��R�z���L<�b�v^�:�63B�	SޖQ�ӳ�-��~��`�u��2>���P�ңR�U�^�h]��6�jeIZ��wt�W��{���b��G�W>)=7ח���]"3�m���VL�ꎜ�ɖ��)w�ͷ3eF�^oT���VDK���GWÞ����ǒ��{�\J����%�=���+1�,q���76��+��O^��V%�zoiJ��\lh����śh�r�㺎�����(�����<���
~�ͽ{�h��-�ًne&XG,�1,z&~�h���S+�jIU��,b�K�{�TK�\�nf�p�S���s��ꡖ{�����
��&���ͼ�mM�vjVL{S6T����ؗT�uU�fE��?�r>��,��黝얱����y������^��t��JǤ��-��ܷRm��g��ټ0m���et�{:0r�[��^w�2h�H+n�v��WF8d�$JDB*$�gP�!@!����xg�lI�˖���xN��BX��qՑZ5H�7�;��������z����k�K� �]-g\��+�:�L��˵��iV'w)��u������1[��Q�gs&�X�E�9�X\Ô]edOV罵q�rz�O���c�w�v��̅!h�ǟh7-8�8���t���IfU����:�WϹ>*��1�4��uYwq���y�E,r�5_��J�ݗj�ᑘl/Ě��^��7��U��]}��{ke��E�8b+6:R�;Ջqڮ��]9�O^����w;�t�f�չe���fh�5n$�FP��Zͳw�-�o	�O>�Ϡk@[����i�]���F>M9ƈ�<���<��v����"rv����m��z��0�u��.���E4v��~�Sp7�\��g�~|�A�޹��7�ި��ŭ�͖y���h�n�v�z�Iڒ��;UF��\[�]�j-q���:�ޏ��sw��O��
��q�%�e�k�P���tX}��IVưq��8�4��P�o���������U b�2�>�����NF�H�D^Ev�M�9S�zw�X�2�������ܪ�Eu��U��S��5����"y�D�+�Eo,�Y��>{<�[�ye�)]��sCz�at�Dю���!��5�;[X�o`7fEh`'QZ샏����r�%u�	����:,>�e�1o���Y�ܗ��"�z���˻�7�������J�;1N�{s �b�+�ſ��.�T�xӽ�Fe
zw������c�%��<ϲv�p����"+P6=@sC���&�>��7l,��X�tzvT�h!@f>�;�v����7����V�Ժ�pq��~���~>��n�\�g�nE���.��n[��k��R��)�t�1"j��qw��Tk{�ad/l��r���l�C�-��kI<ӝ
�p�ĵY)q���%��;{:U�@��WIs�>3��8��x�+8V�Qȇwz�MB���5m�����*οf��Ԡ�/u�G����T��w<n�TAF6�UdLNokn�x�(p�b���}9�s�:7-qz�S���h��z��(�~�G)y���e\ë��֫�jʺ5��V�*'a,�G���-�Z-8U��5��v��z�����|�H�6�{�!�+/�j4T!��m�6(fl��V��L�����v Kbg?�m�z�kZ�u�NI>�U�>���o�΍�dk��q�>W��!Mu��S<�'p������̺�5�Ԡ����{�/�,�x��*I�:��u=��j����'R0�m:�q�̈ی�D�Z=H���/��|�n���v)zݘ�S�r�I�9`a�8���<�9����5G��ա6�q��	��"��Iw׀��4��um#������Q#Cwl\:�p�2�i��o.����8Ӡ�������K�c��~�x�z��>C���HE�n����n��o@p�D�#/�@�{��Ie�y]�R�g��u�l���*��9SGrR�!_@�>�륛�ȥ��*�#dz�_6S��UZC���5Y׋�0��}p5.��{��8���qg�d�V�W\�<5�6;���f�ӵ{�/Z��ũ�H:��q[�Ƹy�תF]W�NW��c�R[������^vY���[�f$C�'�ٯS�2)g?5�Wb�Y����Z�^Ҥ��J�xk��<��ε[Tž7l���'�Eܤ�+&O<+�Z�H庮��Qz��ך��Ί�N������q/�w�8㷫�I�5;�lZS`�^���֦��lõ)��ʭ���qPı��6uG��7�R.e&��>u�}b�M��!��钠�"�f5fKE޵������=H�Gw�����q3��ꦄ����u*`��{��)w+��b`ӑ�6�՜| 	���DZ���N�S"=l���f�-د��YJ٪���4ծ���;:��p��C�g�9teӫ�sv��s�[�S����UǢv5�/ee��3)�Ǆ���_Uh~�t�:��㹗�Ƹ��k��(q�%:ڹ�[��������l�0*�3�ѵ�.��a�+��S(�3خl����Ղ���k��I?�������q�
��<���l�Ӗ��ǜ��u��f�[�j=/����κ��Ґ�M�-Q>[<dZ,�I\���
2��S�����P��wVIzjC氇`�LM!�=f_]Em��rܩ���8�O�z2��!.�{�pfX�]�9�t�#׮��%�ٱgVeD�27�n�Մ�LTSVi�C������J$���ؗjq:'\�[z�WW��Z�4gML#�1fǎ�W@r���꥗�ɟ���S �{1SR�Eg�.�q\�w��רT�j��"�`���慙A+qj�ϴ�7v�P$om�cէؙ�%�f;�:��1� ��tG���vϣْ�h�%�ۀdr��/ ww�\ε<��:����B�ȷ/��[���`����#��7|���g�sbz�^S���3r0�<��S3�1d���)�ú��L5*Y�7�kZ�wo��y�ufe���͐;o�W'%�)��s��W(|dmd�G-�
peW�#�-Yx��kir����@z}�0�=��R�"ksdL�`i$��&1�Ke���3S��n7o��Y�쬧����\xF���ϖ*������i.�涃�9:FL�^{ۺ�s����@9~�><��.�r�g�lBΙ���������L�nWH;��6�k&�Nz����zݹ�E2/��7#.�\�2,304�&ㆬP*�|���%�4n�\�S{���A�/5T�Y�2s��"#�N������
�����y2�K�T��������O����_�>��;�[�Pߣ����@x�Sb�d��ݹ�� o
uCi�h|X%�v�!��ݺ��+i���f��%�����۳�V!���5�{s8օm_W���)7�]0�"H�n�]�
`5GG�븈ǇO�TI�neo>^1���~�����)�ˆ�A�����ߙ���_�bc��[X��x�%�\[�~�iSTN@w��%���p����i&��y�MOE����wE����9�ݔ��woY7�q���;jwo�ґ+Tv4���D�tF4�gݲ6;�yX�'�RR^e�c�(x�7t���ͱ>^��^�1�ݥڝɦ뉫�U2u��
���d�����g�w��S��Fځ��3+�����ȕUK��Td��х�27�����:'�P�����*q�m:f�� }S�2�y��˙|M;��f�Z�q�S�?o:����[dg��/�����SM�s��\S����^���ys�&�X�.�k�����ڹb�b�!QɡX�BJ�����aܶ{Q]XMЂ�`l>rܶ�/�]�_&��qs��-�9��J(Ob�e�{2�y.u�kע�$�l��6uƫ~�m�f,Fm�_;�3\��]��^�����o�CKl{}y�KN�\9��v2#!���T�uQ���w�׽/�����2Ն��ښ��p{֎�^�ˌWS�]Gƶ�,��U���Xޤ��|�'W�sks�]��gq�q��q��@|/���F�7��[�C�GD�C�,;�U�Uɂn��8�����n��6�Y�ƻ.Y�I����]�U�B�$���;E1x-Ü�.��;1m9�S�3k��`5sc=���� �+(1	��y9�Fu�4l�F�{|�jp���m ���&l�v��8ª� �o�!s�d1���p�����F�2�8��}��@x��!�t8J��#�4f�c�#KMv�q��ck٢��u��v�Sq�r��Ƈ��X�ú�s�S�"�{��|�W�!�yd)}��.+��������9%5�O]�نQ0.y���B�� J{��W���Q8&��s�\S8��}[5,�C�Lϊ��X��S�0*��� k�s�}M��u�z�xv�;y}��ەJg���eD�,�긇�Y�g���;f+M�CO��q��w��u�]�K����>��u����u9��L�M�m�UՄ����`IE6�Xͽ��J{� wu�����jZD5 ��y+�;�}Ց��"x[s��O��7�W��)�}ʷ;Bl���YF�B�H��Ӂ�3�����Ҙz�Vm���Ӎ�O�`U�#@��g}�Tۦ��o$a�,�-,�iW7/*�����\����cZh�2I�:���Xa|��!ԍv�̹7��bW,}��.햏f��5zG;]}]��@[;ۮ+�U��꣙�Y��e�r��ͩ}Rw�5�H�L�9n����/%�y�,l*ja�sv��yXv<}�Y#�	�w���k�����·������f�t���ٜ/���9H�ѥ�$�|WH(�]z��;�Ok��T^��x��w�P�{׎8@�\(.ֵ�����]��Aim����nۧN���j�Z��E��[�Ϋ�	�m����2g*�p��xCu�@�D�lU��]�������9���u����nĞ3[mp:v7	�!��[���x����Qa���
�Ъ J��ޖ[=*A�Y�U�110>�>9��,w���ǋ���FM��h����EvrQ����U�n(�_JI��
kǆ��L0IG�CR�f����W'U=[��bﶯ��㷮d]p91���[`Z��o�{� ��9N�7"�0��3����O֌x�V������{8Zrq���)�r�&r�%�ʴgki��������{����׸,K����o|�z�+yv�э�-�!�(�#�1]��ӎR<�Sw�lvik�n�:r۽���Q����V��k����M�KD��1����K�o�Vv���\�1jy��w�Eº�Q��Q�]��ƙ�LV�$�&��]6�`5�s_4�j�u2�%(HD��B�23�E�j��j���1�4�H��v�(b�һq��<M/��s��hRv�3�VOofs�.J�k�IZU}|��X�g2�n9۴��2�'r��}k6�J���Qn��B�Q��M��G6��7@�Aщr.�n��E�.�hծ��v�G��W���2�Kv�v0u��l���EKVܴ��X9�Β]N���"H=��k,V5�֪��v���wR�������$�V��`�nkݓ��-�.�*���5����:m���*YL���
�W�$/\ﻴ�7��.�[Wt����5�uj ��V9ɚ.Q@=��K>
ϑʴм�n�:깠�4�E�=�#��ҏ�in�j���M�e��Թ����˻��p��ڃ������,���Ҟ$�s+���!^oh�T�쳄�X�Hf:�J���V;✷4�7ʝ�-�xG+���Y=	N��y��!n�Ԅ����5�U步���h�U�G�s���A��<%�m*�1ҔJ�%���.ZP�mT�>��G7�+O�8J@|sX��)l�Wub]�[2h!��}�XE,��֚�Aqo�oje8�T�l�kj�OP:�=r�nGs�{Ak��'�w�.Ր.lT�0,)}c������n��n:�f��(�����it��͟�]��j�5�Z�7\ľ���0(p�UR��OD��Bl����+j���|���[�6�=B&=Y����X�U��%���[*���Wc��[��Sz�v'�oc����}sB�@������cFC^��/�����[.So�j�U�I�	*6��iջ�Ƥ0b;�"ӹ�O��@J+<H��g�(@MBC���{�(���,�-�j��<�HvE���JnU�Zk�C).��M�+.-�� w:]�l���mgX��s����u�d`���@[���c+e>�ޭ���hU�-a��>�[�N��H�ܦ�o�c�,9A�當m<Wx�pJ�A-�N��m9�=�z��\�Q���'Ht���d'f����(����êZ
Y�H�%v]m4����+�b��`�/���]h��v�/����@:^����7Z]SA8,�;����Z��cB
ve��ef�����Ҵ�v7 C(�2j]�}�e�}S����0�xi��U
f�hd	`�b����.��+�X�mw
�zf8x�V��B��L��	#�I��{����$�IX�PD6�:�U���Z4ih)B,�y��|||||_���}__��d
b�):�mTPh%:Evv�v+�
K�<������������}_���خ��K�(|���4��i/2i4����m�G�ג��<�?_��3�������+��h��b"����1SL�Q֝m��RPDa��͊�މ���t�"/6�w=A�ш5��Gm@P�ڪ
 �Uڝ��P��E�3Hh+�飮�a((("z�LԄ�j�>]�
*�jI����c�1{��h��P6�9[H��%=RtSX�aЛw��������.�������j��ӡ�DIv8�'I�iC�AHQ�=^��f]����仗/��,"��;��-���QȱL�ui�RokhC|�G.�fS�{�S'�Zq��Pm�ۃ�����չ=bb ��9-�j�~����y[M�y�H�u���#Ә�u��Zדϱ��{i?�;`t��[���T�T�u��s���;�UfU�~٪��#s��h��w�$]x���г)+x[W/���H+9���2��:3��ъ��Ռ�p�.UC��^���~�������z�
J5v#�#_I�(��`E����w���W��;�W�@�]���ļ���h���)Gxߝu��"/!�{a���T9ԝ��UNZؾ���-qw1��6�ӌ�[*�� �j���k��������}���~w���6�H�����;�)e�ڝ��Ҳv8���k� �*5���M�����:�Yf�Ftn�n?W>�`��і�*��J�6�d��'�f���7�RX)6b�*��>�ۣ����g.�]�Vu��v�]� �I7�ܼ�(�v�z��Kj���@Xw�9�2�,b�bi� ܕ��l�d\{yc�)�$��t�f�#'qh�[͠ �O����Ʋ���%�}�ylv�����۟����=���/���{���&D����H3ٗf��۹�ԡ.��m�[j�z�w���d����l�k�r��ڧ��`M��m=Gj$��>�j�j���RIbhn��$jy�$��,���<�<�� >�0~�)�h�ت�E?��J�N�M~J�C�z����a��˞H�J�Sv7W�y<�\��k^�=ivϫ�w����%U+֢�32�]�lba/n��2��*�L��E*�2��cZ�ދ��o2!R�v���֊�ƚ���U�U��dxW�o \\��,����}�W�,��V��	:�����]��o8Q�wc�%���>���L'x�@�t�wP8���X���/��vOv���K L��q�>3�����}��ngj~8���5t2�;��Y�Ս��.�f/,��5/t���gL"����ż���u`#ך	���;!��M����g����z�l��f���-�X�n`8�PJ�.��9�ܫ�`��e
h�P����P�r�e�����3��$k�תiԷko���;��.����qc�>����8�Ϧ\�ZW6T�vn�7J�`�tz�wt�e���S @*�(3E?��T+���[���b�%Y�^����F�b���<�Zģ82�g8j���ʗ�<E�!އu�@w�[��k����Q=�3�ٷ-���撍7UԿM,�юo�کR:xbl�ʎ�ʜ����t�C��,uՆ�-���k���8��+b.<s�\�y��Y�P��u��s]B�؄�JY��4d���@a���&�묦=��ut�2��CG2�XPg��y�E8��d������xM=�{.��oEo�i]����;�ݧ\��EW]U���Y!����Y���xު,2�kυ��p_�oH�[,s`~U6߶��t�3��#Ǹ,���8�M��;�q�S��@lǦt%^��5�.�$�2}�e�)f�kɬ�w���#5��D�%��pw�����M?��*�~=ޒ���
7�|��Â�����w57�6��M@lUM��*�6�v�Y>�(�< �&�d9h����n�{g8�OA��b6l��/��i����+l�8&�z
�e򃍤0�v	�� �\�8&�ɵs����G]ě�g:��}eS9�f)Ϸ�V�7ukꏈ��ռ׳�p����T��e���zxW��k9���3��׵��յ�uP9V�Yu`7{L�Բ�7�VI}�Mub�Q�|�n��8���q���	NJ���T�R*_�y���;��JU,��>�d>��ڏ+�~8�F���Ku%[�u��v��J#;nMH����N)��|�[#�Uosw�-Q�7�����VF��}�v��5E������l��Wx��;?�L>�ș#�9i�'.V�\�Us+c)��el���G\<�fc���k�k�Ǯ��5,�;�yV=w��c�᲻��$j�<�b�m�_�P9�bw�n�zu���m��X_X�,�����
�z�7UOa�����f�i�]�X��Q����p���!�l�˒�[���[{t�T�z�混w]\k�Š3�9����KהbϟjF�[���f;}X�̖�Wczj�m����h�%V1\`E���ia�yz�uVᦩ�E�@�4Tn�QAx)%�n�Qܥz��l�{�C���� Zl�
ٶIVBP���v��Yoc`���M�S���� �z0��`]�ڸz�7+0q3���D��6�FŌ��{�L�q�/����z�'��l�g�n��s��WaM��ܽ̕No��1��2j�Z�f��o'�2���<T���]o���ѫ���9i�����W)�9P�����n�L# ���$�,_��k���R�ص4uuk\�l��ո�U��[���{��Y>� R�g�+��8=#Y�j�j��8�"���H��[�A83<�y�T��{�{<Ͽk�Uܮ��Dw<|q�����p���MŻ�>��|+� ������,�	 7j�k�p�V�2��Y��6Ey�L�<smR�g
�E��\��������hY���-�|y��,`�{��E�S��'����<�;j}
l��N3!f��j�0/���A��������[΋�P76�ò�u� S��;�u$�[�OWNSn��cr�[����u6��&�7��=��Y����q���˾�*�`I'/�ބ��!��d���cк14{��Y]j-Gco�,�D�w4��]��j{�":Q����2�Sᜫn�m���48�1o"jI��PŖ����S�t=�6�uVn6�?xx���9���˚v�'�*W&����9�����^0w%GoǮg�E�k��u��oo�3��(7n܉�4��f��=Z�Ts�I7]Mo`�)���9�çbWtnyl�Q�ޘ�Ψ�����m�h%�k�ٱ�E9�୓*�5<�ֺ�pWm�����"�IR��2�aXիg+mt�@I�ubu8n����J���]�����0��HJ��mGu�]�;�(G���j;���F��kW��>��>|��_����=B{+��tƟ^�q�����Ʃg��5�{�(=-���׊L><T��M�6�:[}PZ	�	���̵2-[3�pfu��`9�!�\¬���ݣ&��&��yP���k���gՐ��J�9UL�W[ $ed̾ձ��/4�\<l+�YƓ�����4j��n
���t��r]�jqT�-��/���Y�Q4���m=,�`<ưl7˭PS���g	�c�l��3.Nʱ1UX�J^$���N��mwV��u�ϕ_�77y�p����;cm�����E����)��w��o��:.��`�n�xf��D+H�*������&)���>���h�$��ղ����,�hf����dW����d}P��D0��RhMC�n�C��w��Փ�[d�>�я��iod˶��]~�x��Xc.�Qj��@��ɖ�Uۢ����9�d����؛�R���-��y�t&-�Xü��&�Mp��{�g$�xoj�[��^ݕ���~vj
����DKͨ�F��۩&��B���t�[��L�71]���k0&���YSs[�7�u�����V��vý�x<� ��H�U�v�K�ؖcZ�O��f��ǵ��3㔋�-&Yu�Q�:�oWB
�F`g筚m�ix����Uk]�@��S+G�z�\�Q��+\R���zQQ�m�Nq�k�d��B._U4�k����W��T1�*T�Չ쩈�g5�ߏ
Hb3��Y>�Qs�,8�(�*n�r�)�zF����7�L�%�MmF�\'
9A�]�첦m[�z�K�n�H�Y*]huwΉ��
v��:r�R�K^$�EϠ�q$��9�n_z������
�W4�U/�[�Mк$���g�s����}��ڝ�Xu2���f;��s���͍m
뻬c̮����V��#_�q�ڟW0�,.�O+����ϯas���ڗ:[�u6�顯m:o�C�����D»��	�y^U8���S��:�|���Rg�K}No�J��4�#��hp�Lz��@�uM�&Km��8�%?f���_����[��`eQ��W��s�G*$^�~�qk6Y���ź�V�?n{1&����������y������1�������;�.!�Tҷ��]�g|�ooh֥�p%+v��[5W���S ~A�
���z*#^k]�0�4��L��(K���X^��ᷚd�W�8H:�*�|�>o:݇���6�9Lm����Uf�:�D�l
�� w-R����)����&�UUs�n��b���~�v��B���N�ܴ�iv[����;��uO<6w^�	����+���f����V;�t�'t��ڨՁP	�2^�����غʿր4���h�%���Ѡ�5��.��������X�}3(Ak�����7���	�*�
9=Ƿ��J�}��&f�����]~��Xw�g9M[�5�j�2�'�6-�Ұ�`7ie2�XzC:O�;���W��-��7y�r�I��m�9���� ����Y3��f��r1�=�6��Ie�F�5�}��w�DS Wi�a��`픱���IL:�L��M�7�c5`�P�;ր� c��.^٩uL8es�9*ܚ��Il��aq�w�v1���P�r�zS�FϜ���e:f͍6哎�)��|ɳ����z��T�k�TX����/4)u��*,ut�wk�R;�w
_�(d��:`=j������{�y�Ѥ�9�	�
������DN�i���ԓ��R�Mm)x�i���ר�05�/�5�����k�0j��a)�*�������1�z��pÏ�OL
�~W)ڙ&o���߿sn6���>��W%��򋹗��m������+�]�v������-�}�h���x�5��;~�W;�����0��b���T:��r��Z�3�Z"Ğ��+�\����{�9j����D��쒻���U9�]{G����+M��wBh"��$��^B�
�j4�0
��sh+�^�� ����k����>��6�&�����9ڄ1:�)�3Z�4�)��й����=�_dn��ݝBP�Ճ���"tr�7����fT�N�=�{o�g����{������תd� U}�SMrֻ֍�]����N��M�[�jF�a�R(Yx�ܽ��W��qg��M�چY���}�J!������ny�h��攧��\��{�'������E�^ۭ��y�'���|�:�cVe�{�W��w]ƪ޿]fg���^�y��a�$�m^6/�+��!��j+,6�k���%Yv��*���]���7��}\�+8'Z��N?mE�"a��v�b�t���9�s��L{/� ��t���*�nC�1&'oY'�Vȩ`-�Z9��9>p�P�q+�ٝy>;]�|�UuJR��:����%�t�b7����ΥӲ�: �l&N�Ԗ��I�l��ȶ���=ܩ��Z#��^.-α�5]�;@�9�6�������w��9G� U��AQ�_#�ʊ��
���}������~�7�� @aT�$�B!	T� RD��T��T�ah`BTd i�`EXBQU�$ �%Ap�����!Ȫ�(eEN���2 ?P�y����=�����
�B �`0���p� �J�*J��*J�*�Ƞ� �H�� �B��B���B �*�!" B!" B�!
�B(!�B�!(�@��H��*J���@���B��J�!�B���Ȅ!���B	J$!
�
B!	H$! ��B	J$�(HH$��B!)H�!(��(B	@$!
�(BJ+C*�
@��$4
B#C
��42)J$!�S=��pq�ɾ<��p�aTÀ���~��7_Xqӏ��>�F��������F>x�����?��������_h{_�{  T_g.\�|��c �ڞ8_�~���!�� 
���:�ϣ���3��zp/�?a9��x��vX����E@Y�D�!�I�H�I�H�H`R$RI�T��H RXT�E%�I%RXD� %d	D��I$R e%T$�HeF !XF�A��a�d�e$X	YHR��``XYFVQ��dH��YRE��adY XB�!Q��hVQ��idIFR�E��`�a��hE�Q���)
QJPB�?Ȑ(�@(@(T�B��T)h� JQB��h@�)D�D�F`RID�L8Q0ri�1��|<|����
4
�@��H����ϿǷ��1��]��09�@t��O�ոk��{vO�e�����y&�cШ�*�ڇ�=���P^�DWևk���R�
����7�
���2��&C���4�C��['H�m���4P5T@qԇ����@{C�� �ѽ��Ӵ5��:���0���=��� U߸=~�DW����t5a;�����2'�!�;�0:�Bs�a8��Q U�7�`0��ޙ@�@���~�/C�K�z� T^���d:]� Qs���ۧg��C�?��
�2�ˈ�\ 0��� ���9�>�
��ޥ(HRRU*�"�
IU$���(�*�P%P���J�R
���P�"U(�@�@�@� DB�D��J�T�P*�R�B)U! �H�U*U*�"�B�J����%TT@�� A*UTU���U#�6r���RU$���D��J��RQT�DRJ"���	R��J*%J�BP
)P�Q$���HS���*��;� ��S"��i@kM2���A�M3Vh
ҚLE�ej��[m��aMBV�V	i����[hҬթ
R���B��
�P�l�
�Cp  CB�
(P�C�;��B� aaB�
  �WrP���[ iYVѶ���1T����[leA�5�S[kMI�f1��5��� �)(5�*Zʪ�   l\���S+%6�(j��SV�e�hT�m��c��[�66�T�eL��լ�++@�h�1�V����m��
@��)$JT��  7]�m���)AT�H�m[CDA��R)U��*Q-B�Q�%!deZ�6�QUUP�Sj�TP���UH֫p  wV٬�3FE+ePDH� La�P������+F�X�)R6���	*�Hh� B���   ��	R��5PP��+$(����H��b��$���hZ�P%R�ZET*6�AEUm��U[fI%
�)
��P	R\   
��[@ �b`  6��  lL ��  X    4m  h�4 mTIAP�

�J��\  W �lM��C0� (H�@	�U�P�P �d�  ,� ��X  � jE*�RUH�"��  l�@ %`@�� (ŀ�
����j` �a� 4�  j�  �eV  U,"A*�@HRH�R�[� �p  1� 
 ̬  �`  C,  	�  �F j� (PCK  YV   E? 2��A�� Oh�JJ�L����a4��M0O��D��O)�Pi�  M$@�SS@ ��BQ����'r%ce����h0aS`
7}O|���k~玼��u�#��B�u�����!I:�$�HH~�!	'� �!$��$�!$�BC���]_�����*DV��Sܔ��)
�b̵բQ���y�Z�d���Њ��k%-�%�,��<�2�J��_��6E��Cu��ŌiY4�Ж0B ͂GG76�љ��JF��L��Z�
h�M%Y5����V�Q�S�AY[�%��l]6�xhSsf�r��y��T�&H�����(9��太Z̲�G$x.�'oL�X�-P5��)�)P�U�F� �(��1���Gn�E�ʔ,;��Qn��pS.\��4Y(c�at÷;kLw0K�h]�9�&c>t��r��pU�&�F���uG,0�Y*U���l�x2R�(����4 -T@��Q'���m	*^�Ч��.��nn�����fxN^*��+f��W�ltP�42R�����ma�i	p�ҞDį�.�b�e��Һ
+D{^X.e � �:X�AB�鱛xu6��T�)I6��R� ��&��swR��2]3r��N�N��om�"^E�����R���R���YG㨋�V���#Xڬ��1[[4�-b6f��[�W[[	r��gn�aS��n�J7+*��[D`�phО��p%/2�-��	�VE�H�T�F��D�@�Z����:��AS�H��%�����cW���ҙ&�����uyN�Q	M�z'����TZ�Z�m%�maAX��5��d������e]ƥ�-�V��)3�xX��&]��Z�ԮÐi�=OL��
2Lne3�{-^z��N=5j��V�D��$�?dU����w�c����F\*d/,;96�(;�Xk�<ҝ$��;Lڃ0�";���[	�X�X�n=.@��aB�jI��"���d�K��w&V=gH77e���X�/$�7�jJ�U���sl�6�ɘ3C�g(ǲU�4�̃�SX��"Vn�����ADLa-�VYObmmʄf�yjP� !��Cr�h�M��aR�;���nd�����d�˰,o"�%���@WSr��Fm!���!�wv�����C�-�4ē-�8�]��Qi��bf�][�ITKU�Ԡ\�6���62ʶCGB̻:/��70KQ�i!Y Ǆ�Z�� �˧)��4&�42q��p�Ŷ�*̨�h0��L�X�s�ē�+�d�sN��pZOn�6��ܲ64�t񄦩Q�ݢ�p�k��/+NX��*�	S3>��u8AhY\�4�{���f�V/\Z�%��1��F�9��8V�'1Ci���(Af֭����^U�b�<[�5�N��!L�FE����h�aSF���>ɒއ�9�0i���e�uv�bU'µQe*�74�mbwy�b�+8��۵�s[c�v�ӧa�29�7�^"o ���l�����
�3�U����m�4�n��𹕰�x�n��e�qc����G�%�e��b�:l���Б��jRɖ�¥[���H�լ��6��)E���^��H����P�Q�Cov�Iw�ckefh[l��vv�y��PԲ�`�V��8��9�^�e�
�	nD�}e�L��Cn��6�Jf���v!�OR� ��%'N����=�qހ�C1f(�M�P�iN���������Ι��яT�@��Z�L�;@T�V~��,��	,���u�0��U�/�kj�!7b���;y��!l�z�ma�J�	GC��Z�G���n)�[șn��<�nB��C2N��(��e�"��w�D;�a�q�Л!y	�s��	�+�f�u�cLk�C�۽P�8�L��l�"�1n�ob���5���`�F�r���|��^��Z7j�eL����(e%dP��f�iV*��N�N[oQ�m��b�1Cs�M���*�&���$vk2��f����Q�6��v%kA8���q��.X4�뤫�6T��T�b�l����Ceɍ�e��%%�	�%gZ����ECY���1cz_�/mk�A����E���ec ZTӚb�ũ�א��w�Am�v��P{r[ҫ ,k`V�&�D��.\zNGXgt�8�^����j��Eac� �i�(J�AMmG���:,�{!��@'��r�̭(�aݩJ�k.F�9 ����
�h�: �y6[�eQO0+�%�xP��݃�@�O6�Ijݔh �g�L�yTd6q��������.QcPI&4R��P�� �(n��Y�p��*�Sr,��[�kU�[�Q�#*1�X��YY�`�x���Yp����ܹ�X)7gi)5ą�n�`�j^U$�p����3\��=vnD4�<�<R��Q��-��m���X��C-l��-��Zə��.Z���S�ebyY�Yqۥ�%�"JQ�C��u�5���]��4sr<��n�m�1a��M��e5IMvP�,�,,��
DG�A���@Xô�{�.D�Iݗ�bh�z�)b�@~�:40۹kcw�J�ubD�n�²#y�Ԛ�kϬd&-�rm�ol%� �����/�u�����vV�2�	���SX��nY?.���*5��A2�v/h醲�f:�̽ҕAx�����7�i�2��j�����1��,F`Ƥ8 &j�6�Y�����Qh���njv�r���n�m:r�GkpY3eM/1)si��ܑ�B���wXԌ��f$��Z1bK.�1M�KjV^؆!+"%�5��v�0�Sy���<�ѭa�t����f엲�L���w��ki����bb�؋uxZ�)�]���+ z��7"sb���X.��Ɲ�c9;�ҷq��Е��	���;�3r�B��H�$��W6�Gm��@�ޣP+`�ma�)��6����e=@�دrV��Xi�ZE�:�܉r�`F�+��W��;�b���:ڒ�|�a<��DCj���ݣhm��8&�:/L[A]�Р��*#u%��ӣWt�W�x	�G);�z:�ۥ�]_]���9>�0�b�u"̽a��ה7nۛ�B�	36�K{�I��:8��d۵7#�y���Ácӗ$MS�Y�s2a[yj���t��n:�jSȍ5*s\X��T<Fޕo7l7X��Z�V���BA�Ҽ�&`W�l2%���'M�Yۙ�~bm�f�\�1���]�D���Q�7J��_Z��f��*Y.� �mnc��g7J���e:"&d
���@
�����v��3z��p�*�;Q�"u���r�b�kie���RԍI���د����ŻƘ(q.�(ښ�r�S]fU�! ���Ř�(���ঈ�Ib
�*'m\K#ܣ[,S�j�b=B�n2m=�i��͘��z3EѶ��R�M���!��";�̀* �'G"�D��qjۘkr�ʲ
YBe�w��J����r����1Ǭ]�t�+�(ԽڡGl`2@���LMMX7Q2�(eq
�8	i���D5fjʆ�L����j���E��U4XT�#z�Fr�X�BN� �Zoo�V�mW��{i��Ԭ���NŋU�.��2��s1)��r�7�%X����5�ɖ4-&�U�c4�mT!]�5��Ѻ���$5�M&�$1��q\Q��'fUǎ8$�m`AVT�"�%��mf�PV�!z�l�ϊ�t�G�H#��L��C!�7�h�ԗn䨁���)���,k��f�R��bЙ&#/+q��T��1��lV�%x�J��a ��F���&��L�����L�ܶ4�Ya��U�:͎�dâ$�^a���z���4�&�h_$������ՠ��M�1-�0�iaۍWij��6���d��v,m\%e�m���I���NU޼�X[�(��0��T��_\�t�9ݨ�n�H-���9y,,8p�3U��O����ږi������x�M�!�L$n�qЕ��cΡ�"%����Ë\�]�	�֘X)2����ُ!��L�xd�d�.$����śG���Mh�k�v �wE+z�f�u���]������Wh�[�k"���)��ն�<�x��T�W��&5�YI0�� D\���6��Wc�-Q.�PT�~6����=m�����[1��*����s%��I �e�xM����GC�w"4��f��іpe��_ŕN�JP�bї��HB��p������GxLA	b�����Ɔ�J���e�^%L�v2<v�7�o3jV��?)�:�e"Su�bX��̀��2�S��㤷\p�v�*���:�kVf\�Ai��)�2�4
���fi�RM�C�y�,����p�Y�.�$ˉ�*��f���@1�4�;�jbݲ#sYç/V��	
��*`׬$��b��aB�̔�Y�TfH�����G� Ɇ�e^0S"��h�Yx�`m`2���v@���	�f�ģ����+)JQ�&� �nڃ
!�"�f���(K���uf�|LE�ʼ�]�k&Q��r��a�HcHZ��tZ����ݤ����Q��y���w���Ǹ�V`��]���m��0:��񜅚����2���p�X������x3.Q{16⼱)�@M4��vűmYoR�&�<��u�H;�N��f'��R�B�Z��&Y���),��*�ڭ^m4�+5���l1V�l�m��IP�ce��^h��с�+s%�4�`
p���W-K,� ��i�`ZyX&b�#���.�6^���,�Z��n�E��Mݙ�����,0Ib�[z^ɴ*�*�J�&�U��Ҩ�2��uni�J܅�0�#����
���cw�ڸث�V76)�l%1�J�1$x0��&�sfS[��a8���Z,�Ժ���P�{��յ>�)��-ͭ�T^�%axð�p;8�W��Ņ �nˑ��ܚ���&�a���4Ŵ�!3HK�qX�,-7錇Q��R�VUc���u�e;ͨR�p�i�f*��&/d�飺�Ѳ�E&���/p
ƒ��^��ӑl���DQ�h��ֳ8�գ�3�7l�yN�����T�Y[� �+s0̟aq����Co3*ƫ��Z�f���b�`a۰7i*�lJەj�:ֆ�x45��+2�: ;v,X�J���w��-M"���*��]�ڕ���Z��:�ZYxD*��/.�%�G>�a�,�bO?�fø��=��T��nT��,G"�N��]�ǁD��.����Z�m�V�a+G�O
��ǲ�^Bn*ִ
x�(�i��KVJ�y��cF�wh+	fjem�_l�j5���w�k*պu�t6i����
ڽ�.L�v$����F�eѱR��j�[N�͎è�wa�mڛ7pe�S�r��1������eY7�Q7X�&sEH˼��d9.lZDS^����ug�)� �7V���	zZUb���m��W��*�UC�l6��࿑2En��j���E�P�%]M$��pM�����k)<fFE�ui�n(�[��� �x��I�nK{+����Вk��d�p�fG���	ɒ��tRxoI�I�J �{���$&��nbl��f�˭��J�l��L�6n
�ʰ3n,�.��a��fb�T��k	�X֣��ރ��Ҋ�VM�d����Tְ!f�Mڻ��V҉dXD�;�n+:ܥ����-�>����7]ފjm$�0�fnӰ��+U�<��4���境�*̅Js[8Ҩ&M�O
���S��]$���FhJQ�V�0=6��we*ǎ��vQ\�ϕ$֬,V:�k$��:7�b̔���+Z�'%yuM��;�4d�S|ҩl��.��V6֖Cq3���t�]�˨��@�d}	xR-V��6h3y@m�ݠFP�)�,�����d�A�7+^�[�!�VQ���te�dm*�Щ�hx^��j��ʌ)%"M���#b:�.�� ;�Vm^1��kV��.���E��a8���c��Z	m9��Sr�ۚ,S۠�GR2�0�B�J��#����7�5���$�B�2,��j݊y%1�6�w3~X4#��4̱,l3SV�Mu 7p!��2鶞�W`��mhHaa=��"wRT+Kݼ��*� YL^V�V�lA1�-e�݁'���xu��B��P� fk���;h���1���wN�J�v�f�WX7�y%d�j
��&\����Z��j'��i[v�
":�����F��ę�]c)25PSH(bY�,��U/s[[gV]i�E��q�7[&a����.���Qk0_�wK�3q�U1�Q���X�c�p��[m�ьb��L�1y�^��Y�X�4�U�$�d- ���+i�e�1�v�x�y+I�; ۖ��n�*2�3ZKq^:) lL�w(Q��b�K���P۷��p��j�;
�Z�	�DI
��IZ�LߤU�	�N�r����_eE���^h�S,�1�ń��6�FP�K�!��E����y(A��MR���)m֨��I���٣{Q�qThb	�����Yy��������Ӯ���5��q7N�w��-�����H��c��Q�S�At�#���f^$�Wr�Q����ML���@��R[�u�wD<16�$6ۺ����C-əx �e�3h�(�JO6�Ń�>��4L��^Q�bә+���)�y�Mm�3J�˭�X�%�l+��31�"\凗�N٠�*l.�<�.�k��'�V71�LPҿ�w㱪�c��z�F�ei�1�E0��iM������O���!H
���n,�p��/>�&n�iP�큛vf���nl����y�pѰޕ�2��y{`.�kCS��(�/A�H�5T/]�`E��e7�cq�LE�,���(���̭���v\ǣ�Z.;�5%�(o���q�S-Y��\���0�Z̼��HfCx4�T*PXTH�t��4wK�+h+5;aV�(V�;��sM��A�C�վ�V"����k@��v�R�L5��K�YݲLnl��-���qhV���;�׹����g�J�|��\�9gd�kU޼"rN����C�2֪go�=�ˢG�g�$����w�H<��A�4�����>̥��H:r*����A�vq�=�l�v��������A.�Zk02�
I:�L�F��b��u�Ι@��h=HY\P�r�^)V��:�j�ܒ0��eC�1�Le����i��3J.!��-�3@�F���].��21���:�����K��9�%�s�l�ڭ�Y�L�eݩ9*���{s����[[������Kiۤ�\M^�y|b����|�95�cA&u�A� �������D�-�ȯa����c�U����^���e������q�\�ŭzM'F��*i�d�v��F"G�*A5B�.�绺x�+LB�Fnu�b��R�
R˦"�7�}�v�r;8�0�I�pn|��ȳ�oQ�����%Cר8�v�xq-�Y@n��e�7���]'\;�چ�И��b�hX��]t�l�վ��ɪ:t����A�<����eZ�b�DOU�K<�ު-T]��7,ќrp�hYa���\�@"�WU��4���庾�m�����F
M�N2 �%^_vк��!���o`�գ�2�L�a�9���XU�b�����053q���<�Vf͞��f�]w$K��Ǖm�oX'c�52�k�mc�e�!j_;�ԉ�<�	��s�	Z�ȫ��_ 6`oVܲ��,��0S��`�2��V�h�ێ��8�7g�f���s��(����};0G��sR���_1,���wD�P
����gJ��L����a�����8N���K���6��������k� D0�c+�Zf;h��
f
�ͥҵ�F�cL��W��;{>�uw� g4!�l_�mL9e|ܚ��=�.E�`"��^|DS.m��[�\5n���.�w7�%>�p��qt2���q-����QB�a�w}Ýa�K���m�(�u3�̰�<Sv�9�������cG��n��[��[�1�Koo8�;�{�.�
# W�m�k�|�h�D��[�CM�,m�{[����q�2�^��+'�=��؍3���)G�r�=���r�X�=)[���ҝ[U���l��6�ҹӑh��쬇n)n��Jevbgo�jY�������k�WP�OG�B���t�âd՜�Y���ڗΏky  ���#6%���i����%���� ��s@|m��0��T�\]4�qټy���=ΟϷ0Pul�̔VR�j}��9$�����'I����WO�l	w�"�7�:��Ew�Qo�$�GT�mk���K��-��8���DŴ��=g�M�#�����Q���C��،�Il�xUi�KB���c7�J�k)3��^�f��l�8Gs��9���ob��wN�5('��<���M���ɾ���`Kmt�@��f=o%�:��=I��.
��VK�X}�"� ���4@����.���
jor5�N���\�K��4x��P����4���d���5�]��E�)�)��
OA�kD_r�'
늙�鷵.��.c��}�r;�2>Fф�x�gLJ�]_�K��e6GL�����V�}����P����0����M�v���C�|Ղ8K=��ڣGzCA���xښ�Fc�g�pެ[�r���:��MP8���k]J�S�k��7�w�6t��C���3��)m�.���a����q�2�՜�9��5%,�yr�6ӻ5e�W�_i�9��Ҭ��I-S�غ���d�SY
��Q�z���$`�W��xJ}��X�n<v�B��jܹ�ZOr���{o�88�[��*Qֶ�D{�?��������\��u,v�nG�j$� z.��J�`��&Om�f�����,�����uj�Y&�Nm��LD�Yw�����#��W]�j�Փ)�0a�v�fS��>�ֽW�6���P1�щ�ҐAQ5�wq���]�ѽ���k�]�e�mQ���@�[Y� �N�M�+��9]#W3o6=n㜇�Mԯ^u�6���yT�Ⱦ�S1�xm�u�����5i,+�1cn�\ �ކ���9I�)r�o��؎�G]������,��=�$�`�=��.�f[��j:����f�E�v��T�Üc��hc�l�M.�t̴�c�r�Qh�� �VNߍ�.�}M�������8uY�xE*aa�`������^�iԝ��o`r��b�MoT)��H}���r��2�1Z���`���pi�Iޱ����ٯWe ��rO��"9����xU-Z����&
޳����1m�!G�����.�h�i�Ô����ct�(r�"hn�.w
:a��v���������6M����RŞ�:�Ex�a��kw����(p]a���:˭�A��p�K�b��\�w�����\-���F�,L¢�����jN�JD蚥6р�����S�`r�<Y��`�r�M�Lk4�s8ڋHm0F�$puFY4��N�3�֝�O�:�"W�.D��o��>S�5���Χ0��C�8l4�\8Q{��oRp#��ᅀ�_�n6{���c���V��u3���\e�������p�ׂܸ���W��l>W�#O;Z��;e똀�X�^�>�򎨱w.�1�%�p�J*��՝RU�Y�Rf3�/�+f
w;%�Y{��Q1u��\�^e�4���+�X_Ru!ą=�5�� �_��uفHʢ���s���:c�w,+�c�k}�z��k�ل`��\�y^Җ	�\ٜ�bӲ�$vb�.��-��u���|��`������q�cu�<�y�v(�����:�k�1��~�k��W{���{z:ItYX�b��6��Z{P�1Xkh�I!���	� DΤZ�����Gs9[���B�i0�E�9��m�t��R*M����w��_זt7Ǜ��|�aE�VW�'\Kոb�lWu	J�hՃX�&�iّ�����G��!-�h+oICa}Γ�=s�Ё���FC�o�V0�ie�^���WF�*T�ld�4�R�9����n��Ip���?�ֶu֭r#�i�f<#Q��{�n��6�T2�|������[��f^�Hd��>����v�݅���1�p�YZ	�Ĉ�>�m+�(�#7��]L�K�܁��*�wan4�tév��-�4�qΐ[��h��9D�C��s/vF��K'U>�n�(t.�:�����R���Fł8-('�*VX�o׷���N��}�]@�j�' ����B���X�+2���N�{9�}�@�5+�O5lI����9��5j���QAg��y�1��L���38-�
�ݤ3�CAm�#�/u#QWüTy$3F��W��;��N������F��:�W�� u��f�̺U�[��fU�+3R��h�wW�E=u#� ���:��ծhG��m���C�Ol������Q��w,�feb�c8��T�LS4�BW�z��rm�e�x�j;��1���m|B�7�3�Td�7i����l�]A_.km�,���!�]���x�������7Z��{F.�o��4�H�@�3��a�4mj���}��X�.���LL��s��C!�޸��ˑ�d���P����Wg���_7Cq
ʜj|�f�J�bzjEe�n�J�@^IB�7ZЮ�`u�'�;v��,m��L�y.�jߞpɔ�
VW+��a��M�yj�E���%�5U��b��+[�G��NX;�i�j�H��xR|�� S9$.���9A����S�P�I���y��c�8N4�D�Aft�����4a���4܈��^l�|��k�l� Q�  �y2�R}wkm;Q��6�[\;0�b|ۍJM���f��k5ϦΩCG��{k6D��/i���WT����cν��*���~�sh_YJ�V	N=�{u�):�^���h[-��ʀ[V7���D9�Fp;�����n��ǅj�V�$��r�x^�[pᛡ�ZW:�C��T��:᫠lSg� �,�=�:���+����+q�s1��6����e�b�i���7
u��H<�=Qjȍ��PYo���U�4,�쩐$��l��=j#Ȟ�]��h:�¯��PNP�©\7c��.��d&���Z3�d�k^kH�\z�V��pw$��EvuE|r�[s-�C`��u�,�m���H.�)|��8�(Lr�Cי�����+�1���1N���{f��U�7�!�ۚl���.͙/!:�y�F�]��f���*�h�w-�G���lѦ���{E���aީ�ff��� gn@�#�Q�ً��Κy2��Wt�F�c�ڷ�_Kw��dsy����[�9��l��:�I
7���w)L���]��e/�c�
�*ͭ��ym�$W.
�_M�ڈ2�6|�'�Y��M�O/��>Gb��V^nM0�R��f:uwh���k��mr燛�x�J2���Q M�M�G{;4�[[����Z�\sK�q)��Y7DH�rJ�E**��S��Ŕ1�*e6.��\�Ͻ^��+��Ir���%^O���Wnу]���8��Z�%T�kDʻKk3z(�ԉ�6�X{f���۽�6(0�0rZ<tq��;��{�`c8�ɠ����@-쑍��N'��4l���+Bf�s�mD���gj�qڶ���gZΫ�\E�i��`���++2� c��wY{�F^�;�
��a�7�L�-�Q�iҷ���A�2��i�4��U��Š���[���5w��uu:�[]�hŁ� z��:;wI[�}d�N��]��� k-Sf�+f������9P��y�X03͛����:�ĳ��D�$ޭ���<v)�;`2���z�ju�]�',ˮ� ���l��W�ë���#_�-e�W��$�K1�W�չ��"���6&^���W��`vm�2Zj��cbU�g_\��>�!01>���5^κ�iP&����E�V�В�-if��V�g���_Xn��V/Qx��Mj��cÄ�ؚ'j^�L1n�(RK�s����ϲ��Wu�SU�ga؅�7�ȋ:5�6/_�ݍ6]JL�ŷօ`Y����U�&v��Qد�h�Ј׻�6$5�s�����]�3��OC]��K�r�5��˱��Z���)��A��;�d�$q5�%ss�m�;�3�;o8��*7�o�y!��Q��[��Et.⬧��֓�{hN�,>鍺�aV�WY3���^�]u��m��6��z�8���V�竴ô+1�:��w���촆�y��ܝ�$aQW]�lچ3^�����ն�����3kn�ڀ��ܻ�w-ҥJ���ֺ�x`���K��U���˵-�D�Bx����՘���Y}�XA��\&��Gt�]��h����Hfh�q�^,j�%-nѭI��}6�����j��k��ܣ|@���&�ݘ���I�*���n��OM�.[�Ƌ*G2����W�!0�=[��۴�zm�ˀ�-����N��]Y��Ds/.���}��ĸ(�J�N��:�n�*=��+T���Ĉw9'xt�4gI�N�^�5m���JÕ}�E�2'`;�gsa�Y
�5λ6�߬:t�Md�J���E�����56�dF��A�30��z(l�1�v�E��ɀa)��eO@�ªX��[��VM��QS:��V������X2u0��fWWA,�Y��c� J�����ʎ^�S�����%[��Y:��l|���`��u�#��u�ǹu^��h�w�p.��d��Ʊo��7�2�X���z�t�6��,�oDdf��Tj����uuԧS
�CN

]��8h�qΛq��W;�!�R�e����v���{�&Tt�S���Y�.�N�7`��R��(���M���r+��"n�Eř�����h��#�T$d���Ӏm�O}��&�����*R��2�Vb�����ޣ�AT�e*"Ή�n�t�s����Of7{���� )�Ji҇K�\۴l�k�m,{a�N�����E��5�'��-����8��][ug9�o:S�w��ip�O%��A�y���7�x1�n�w}��y�o�h����=�ܗDz�01��i�R�een�ٓbEP�V�s6�^&�R]��N�Q�;��w��G
	�v��q����%Q�S�9�]����n��B�zw�w:����"A��|E��on=Ίa�.ef<�1�rc{��m���wt;�T��{r �D�۴2lMcW:�JF�䋕�6�Wr����[6��v�W���CF'��vF�ei�ULu(�w�a���ي��<�m-3o$t���1G�yb�GQh�|���T2�f���]ϥ��e�ր�n}ŭ$�#���ʳ�h�W�D��\��C4��+v�=h�YR�5�.�ެ=��j����⋲����]�J��5-���*͓p=�����b��@M؈��w����.����3e�0脮X�fS #�or��c.v(��c����-Qv��c��oB����<(J{LQB�V>�k>Ǧ݋Qv{��(k��1����.��rq/0e�\�u�ʼq��iJ��Z��hc��Ea3����}����\ZC����.�[�K�*9ңU4��{ù�ԡ+�U2�+Z�嫥N�UX���;���m�x:1����Sz�1�p�{�:�K��n�w�%]g+I�ڬN})������#�nY�tOP�58��۫�BS-.Iv�=�	b3jihM>E뵺�>�!J��,}�s��٘�']& ,KPw|4,e����8�����ν�ξw����k~�W�I$$?!	%����~K�s�w��s.���;��;�ncn;�ĜYs�r���A%o�k`vۉ<�Ծw�-���u�k��A���b����ŵ���q����/�M��s�/P�ي�Uu�4VI��=��:�j� l���˶g:�0)����t�n���5�Gݩ��`f>оB�[Z>�p+��J���i%����z�@��V�h�*�����  wZE%���O(��]@����{x:�]��f�����Ad�M֠�!z�tҧ+ʎb�*�YW0NCK|�]Y�&�D҇_^*;(w"�g�5ֲZ���B�����N����
n0�\4����7���������/4���jG@��#�Z���w����ֻ�w(L��5��8��`�_r��z ���a�@������"�g�s�h�[�Ŋd	+7ה���va���ד��.B�v�\��s^��fs6�Kjf�qVTM��,dڂ�Tx4c��&����U�)~{�0�%v����r؃�t:L��o����fN'M�j�146/���Z�X�����VG%��w��ԖP��cWnsq <�U�S�˷u��Z��p��@�5g�vҬ��v8�٠Z�t�-MOlI����V�[J+��4��\��r��V�v>��n�F��l�7��vM.�K�3
��"�;؅�{�Y��I:t���EPCmj�7z�!}:i�KR��hs����Mm��Vj7�Sy�"�T�5��b��e"_%�rʴ孵��k�LYB�H�0�h���;���\5���O�1g[����R.\4:��λ�����ȩ�c�P[��ѷɰ-�i "�5�ݶ���w�'4�ٯ8D	}[�s#��g�έ�f�O�4�ڽ�o�p4�Z�^I��wE�u2@���A��1̳qљo�|V���Yz���n��ٱ�Ѧ�MG���]�$�YD�������I�K\En�o��27B-��+��UC/��[����޶A��Լ'���ݩ���"V�jb����r���a���%�l�G�����S��A��N�+ Z-�������|����Wr�@9t�c����Pݹ�Z�9�����q��>���%9ǝb̻O�5y��3n=3������uq�*���ouuX.S/u���PN��vkq\᪥�l,�Ȋ�H��خ5������[��8�bq�2���<���j��0�<���or� �e-�a� '�j��%��<aɗŉw�l
�����Zo0n:��/�Sf2n"��_<��r�%��v���B��i�qH]Ԙ�N`+�&wPb��ݫ���xRLh:�/e���K��緷\�b�0[�h���,\.!;�l=�����ݣC\VFi�qLޒ]g�2��$$��;6��l֣H���}[�Υ�.D��b�G�
Y��+N�Yz�g��}�&pM�G��Cp>d��nXqD^��_We_!�sc�Y[ϬnoEc�j
ꢮ��<D��	*������s�ΝB|W.�%�w�v��Ī�ΗCp��(���JxWjJV����DW���\UkXm��LR�ViV�Db��ŷ��έ��.y¢P��r�W�\�R�b<`P���4(�2���{�w��.�/����;�K��'sޓ�*k��SA{�,+!����sl�۬S�Ƌbn��24p{G�L��J�����ܽ`GmW`J��K��R��+�5}�]H��,�DWu�;����WN<�j
<��{LW˺�����y�|"�A���6�b�w�S	�s4M�jvL����A�T9r��;�[�j�(n8G�3��e!x�ɢ*����Ё��ȕ|�]:�Z�ÀQ�K��y�݁x�d>닙�W��wT2�[]�ߚ���V�6r�p�v>db��flw��kh��H���mv���� r���l��;i� �ge&\%�k(Ys�9=�`���u��rW�Qʀ����N	=Ai:��E	���Jޛt2�/���n��C�޳�۵6D�f7ux.Ҿ�r��h�e�JZ�֚��h�sS�� L��-v��6��jn��@ ��V:d�C0�_5n�.�|4R̽�!	n�u�Z�A�]1��H��WX^�4e�Q��
_|#k��c�Z�Jr�i^+gs��^U�|j�먚䂼B�4��V�7(���`�j�G4�s�n�)�__V�n�t�d%���	��t;G�]�u�'hj�����jp|�*�õu�m���2��t����剂��J�v��+0@VJ݂|�=/9��Gz�7�0�� �z��GsFD3U�Y;�K"C*mheh��[l4��ʐfE{�r�c���v���ѓ;$���h.�Q��nS�
Ti2��}��X+�EYb��sU��҂ݝ���o�;�x��v�pvR��`�}�^�:v�J�,gS��
�u���6�4lD�^�Ɲ�S�C!ĕ�$���	(Gn�l�Z��7"��� �as9�V2��.%��2��^�4����Yh��f���L�{�_p�޳K�6a=��6��ԫ�N�=�7�ө�\���j�c5��Hz��p�-�ܶv�ޓRN��ts3xP#�c
���-u&�%ϝ]�o�!'Xn�e�T���V��m���M̚������a�tI��9E�\K�]�9�Z����u��to���u�v�B����+�ۊ�g�f��>1k�`�%]�V�N[�ŉ�)����̮�ˢP�GY��5�����J����ΨK�Y��(�˵ێ rQWBeeJlj�H��X������E�8i�M��eY[�;jMU�8��
�k�*dB�R�wk��2c��v��1�tP��b�U��r�V�<xussb7M�^�
x�r������̂mc1��>�{�	̺V��٩�*FȏF���P��th��e�/J�;�˹�M)��\�B�b�U}*��ZBg��=w֕������ۣ3/4D>4R�0��8p^^&�/�N֠6���2����Eۘn
q�ʍn�n����,��PV3�����F;�@d�O,DsTΊ�櫰a�$�4��P��w��xT��{z�+�Вȹ)���rC��[i�,-]�9+__9��b�-�;TT��D���c�j="8�=�}�ʵ�v�d}�;�M2� 
Ŭ&rX�����*���w�S&q�m�G�c��'��L�^>tl��s���E�[@uv��fګ�Q��9��3�:���hd-hh
�U�3�;�}yf7G_"L;\ĀOqo=�e+/.����7��]g�8���6�rX|v	�p*��*�1Fe���3�|@p���ţk�S�g�e�\���h��^%x�WT����.�Uu1��H�l�k�<T�r��_$uf`�PǹqC��9�Vn�r%���;�@?��yM\b�_=U�?�2�����hT�� 5˭Sz�,��/j}r �*�X�;4�"Sj))^-xpkwds�iA|���H,���1Q�t&�%�Y��X��U�e)�F���N��j��{�^�I�٩հ�*:jذ��4jbU�}+�����o6���:������nK��2��f֕ƓW�*�9�}��aۖ�X�郐�������r�Y)�J�ʻ�Z�����dH�3y,eF��dp[��SO�y���TN�k�ڛ7���S;M6^n�B�γ֢�y��ܓ[ͬ���s��i�����^�6�B��sx�>�Rٷ����Y��PT�nVζ��u�$��*�-���a���ll���z5f�Df�{��]��"&�Y�<�:�V)Q�P��-;&�:r[[�+�VD]4݃[ٜ�:C�Z2�eވs�l+�pQ=1|�]K�b�mr�"|�wrU	u��-�
;]�!�8���f��,ڬ�ت�&���(���4����gΚ*�|�ցTl����uY�rʸtR�}\�+�mV���^U��Vr�QX�iR�\S��4.��3��-j���YTz�]]��4����pՆv̡�@:�^�s(��u#��p��X�Ч��
��L�,vn��p�ᗬJ�hY(�vZ����4aY�$2�bM�q��wǷ��Nӌ����cw(p�׳L����jL�i6����ҭu <N������A���3,�f��3Vwqu5�8&�����f�ҥ�f_7Vymܺ�b:{ςՀ�W�_�t��P;�Ru�r�k݄��n��6�5�}�L�w�QPz^4z.��̪�%Ct���g:���1>ԱV�;���i�3�0َ�'BݗZ�S�]/l.��]�Y7u�b� ����3rv���7��;�K1����H���cl�wBxDJ'4�!����A7E�������o#a��&:��0���J��o��WB=`e�(�ǻoE\����Y՜{�9���8���	˴Mޒ�o_j�����e�	�A�v%F9IA�]�n�v;F��h��i���;-P���ѡ��9�ͦŨ���f A5�����Û0 �H+aow��;6�{�|��וz�M{j:�X��Uˆ���{���sj��sܝ$6��O�F�=����b���k���c��Qt�_%�[�S
l���Պq����q���\�Z)��F&D�e��D��/�	V(�X�ɨ���H���ﯕ�d�S����e�ƎR-����Ed橘���ֺ��.qܝ��+yJ*��8�V'�ͫ)q��sU�z7E�k\'T}nt�w�+0���b���!K`5��#�YO�7�#�P��k�CXj�w>V��!�0��i���������Ә�J���b*�hԊjQ�ϰ�P�mc�����1*d0;: 6��J&ý��`S5n|(����9۬m�V��]Yc{F���z�թIE�����U���hP�Z��7O�s�j9���X�w$��s�Y����x�bwCEEj��8�+V)��dEnU��}�]+Rzؼr�4���5<�44|�5�j�nu��]��
�Ӿ5;ʦ��ޔ��{G����ۀ��V�H�&ő�>y�i��&v�N˫���s�ƌKw�:̴ѻu�[���H=��6��I�.�ͫ|
�u�KoV]���t󌚺�|��K;~��߭[��<j��՝.�Ʋ�:�����#�����NJ�`8�Ww@��5W�h��m�e�Đ)s�Z��]���8��0����fЊec��j�H����*L�<�#��V��F����Y���wAҠӊ��Ml�[�sq����b�b�j+����@��]8zpm�l��gv���ի��ђ�`W��H�`>�w5qq�������� �-�/~�fn�rЊ���c]��r2忺�����w#V@����e!7� /��iln���L�P{8�ί����G�����r.�ܚ�P �ִ��v�1�W/�u�}@�GV��s���Rm%�͏�Y-�Zt#��;P8�ۭFN�j����P�����d`�ӹ\��yv�.�t�mt�۩�7M` ���JVɧ�e�7;�EѲ�}txg�CSXҕ�r���4�S\v���{����8�Bt���Q���G' 1��M�<'nv%�i�y �u��� 0�a��k�CQ��©�����u�`��a��x�,E�L��O#�ʖPӹ�_f�Z���J�3H�Վ��$VA�2�����Bd#6ݩ���h�JÅ�Z�K��l�R�:�H�-���+���z79�a�p�u&���p<���r4x[�v�\m��W'����6��,Cϔ�u�L�4M��Gn��#��XiԱƞ�:�]����*l��cL���'�a�xgBsx���Dy��a�|e��c�ڮX#���`>�߶��:��t%rzr��L�ͽ���6���U�,ǉ�IT�D���A%I�A�m �%ݜ�*�v���-�U�%>�И�d�]}ø����'8���d��/]��3���F$Z/�(d���8�D]�g�Y��64�:Z��һ������wE�$<S"
���hu^P��0��a�2îc�����ұ5k�H;Ηu���pʎ���=��]��ܹ*u�7a�Ч/k����o>��ԫ����ÌUMVOA��4�w-��J���,mŗy�d�����6H����x�շ�'�(.�˚�������Sh�R�W_*yg+.s ސ��t�Z��hKt񴍂fX�&u�\7)0-Zݮ��d|�;�֣����.K�g[pL!X2h0/l������x-�����[ni9[�z ��TL�5̐E���5�f����M�M�i�ܬ{�;�ĕ�''ۮ\\:_�f��F&-=*�icK�,Ia�����B���[[ ��^�gY�5�J���,C>�@e�t�wQ�����)��u�����cT��zA���{Ny��R[����u,4%Mm�]^D%	п��Om�N�Iv�(g.n�=�z[ r�Ӿ�'8�pN��m�U�yV.��}8X��]ޖx+ݪޕ���݄��W�)e�"t`)��L�lz�g��2k'˻�M��E��ݕ�pEs�X�x(�*�E.�N\4g;�]�Ċ��BJҧrw'u��e��፥f��d]����8�����޺�ɻ�uh7Wp7	��R�8�jL�G�	}��lu;����\���ݻqq9�zgZ�[���xi��&�(���Z;�Hgz�#Loj>U�Y�RU��v��
�a������m��9%�d=|U[E�A�D�����-�����ۣ�qC�PwRw�)�hv��&̂��m
y���2��v����]oe_CK���
���iU��E+ڙ��7� �����-tw�N�-e��κ7OJ(�J�m��*�]�˃�u�@��wu�qR������|��T�t���ִq0�tr��T��Jo�^�_-��H�ۻ�k/��d)o����8��
�(�Jr��o��x��m���;|���3�3B����ti�:5/��2�R7[wǧ@Ԝ��sn�i�I�vb��+�2�����e�[W���	�޼�%�v����<�)loQ�pu�}'���U:��Ļ��J��Ll�;�GDh4����$�JWin`
���^l=��x����#I��me�������[1�%n<�z�cNh�f��T��,�T�BM]�����9WM0#9�N5�qKq� nDt��ϱ����H0��/Q<��Y�}g�e�W�a��B�S�kN�%�J��5u:�3��b�wP�t�ۙr^��a�ٰW$��@�Y͜\��,���>���QJ�R<wVHb�G��WR�=w��\j�NV����+n⃃4x�Oz
�W|�kXj���\�;N�J�X1r|"���:m��p���3i��}ɶIm��>��B8�Wz،��h�u6n�욪��{[t�^��t�М�<�*q|9 ]�Up�]�O��Wm�t�O��Xm����t�tg�!�iS�Yw���6�7'<�������u��)���c��ܶ潮�8�� ���)�����w7&V3��7�WW	��
�ҧ���ƗVv��:����p˛tDۃ�?bv�y_ �X��C2��2Fi�יdl�OvfD��7cU;|��=tƵp�V#� 8\��f�w#	8��}���8��3�%�W���t,U�T�R�P��}B'�%QT\a�&5*TĦZԒ�# T���@Z0�iB�VQ� T
�R��V�CcqVB�*QQq�	�Q����*�˘*�IRcr�m�J�j�jJ��.YYP��)����lc+I�YU��\��
UAf!3�Q.Z��T�$F�ʸ�X֥W2�*�,�&0.$rȤ�e���T��[d�Ҍ�b�R8��(TUr�,��e�.f`�`�X(#�U����"��E��XfRF����ʓ��LEb��m*(�@Xۖ���Xڰ��R�,��U����2T�+USH&Y-X(c*,
��*Ab��O�DW�|���ݲsޤ�e���K4����
AOC��N=�!�=p]g*���C6m�%��;gr\ł�.�ve��m(��=UC��Oo���U��=�Q u�>[�ٖk�d��E^�U�Px� ]EZ�Vm�
��R^�X �|:�3Z��pͅ}��9�Z;�ito�1�x�	��{����p-�y	M�Kzx��9��E�#�	����WQ?
�(1�n����YV�aK=��.���̬�Չ���/��`���4�D�=�f�F Xo�ъ���c0��j�#<߷pǊ(d����A,g�o]��*��v�T}3�������(�U�`�r#�I�*�b�[h*
U�ִ\ �J���`�5�@�Q������@����06�ƪ�Eb{7��0��s����p��G�ԥ���[�	ʷ~6m]ynٿ� b��E}��[9Z���-��U�1�E�;عtа�����QGq�h�ӑE�WX�gl�+��_jv��Xk��*t�N�b���ct����t�עL��3ҺU�����>s�0@������������o��2����Ɗ���2�U@G����@U�PsHC���=2����j�{��,h�t�Zɪ���ʚ{2.�_+�vjS�I�듡��.��5뛘��x�����w�:�;�n�s֟s��}4�'�(��(�0k.\��"��od݂J�z@��!�SyatW��E���ʗ"��w�:��]C��fJM�aox;��w�~�Vb�{M�r��IX���ʄ#qD�,�y+^�Y\��븵��=�,?U%L4�5�(D�9��6���n`���1��7�!�] of�wj���Qd�\��<�>�tMh��n�]GX8g7I���C�9�U�v��7��e�nS�}\d��zd3j�Ȯ�V�ÐJGv�vd�_J�l��.��6�m�{*��>Wy��u`�*E|�$s��`����%N�̀S;�"	XW]�l���+e��5�����rvn@�M��̨� ٺB+�rC�1�}��U��+������t`��a���a�r�71m�ϊ�P�9@W�eyf�U�
U��y�Na�t����=�ic�tbŸ�C��Lg�Pu�W%	sڡ&*;]}�V*=�[�C	/=\<0��1�R��ߞ�q!^?d��_k�kjs��.:g�;Q	� Eis��{|-�ʶ����|g�:o)c�Y��9j�;=� )�@n�x ��Y] $Z}��0�m���x��[ۦ�ui�rve>9���~+.�l\��z|ĎK����5�(/�-��V+=	-�2��m�u�,����K���t�-���%��C=f���;',��Ⱥ��'�L�j�T�Gf��\&��u��L.�l����I��[�������2��U���@Xu^�gJ�$D��knկq�uG���\>x*�p�Bs��7N���U��n&����(�Ӎ��A%��ҭ,򦦒�E�4y^�/ef1ʻ����*9,`����=�`�lmw��z=�����Z�E���)�b����i��v�g�����3=�	\Z��
�f�?g1/NgŇƾ��ˈonY�0�M�o��yO����K1�IlT�.*�	��D
��0�E̡�eYAGL���99znVW%X��^�U�*X����Z��t�=t]�Ù��K�@��Ӿ<����\�J��C6���Us�s��I��������1���(� ],�0��rR<���mBF���Wě�x�3�Z��X^�5����O-]��B�2F���9)���5*�p�2z�"2��=6��\\���8^��	OS���h����Y� St�TbL����H�����>�I���lߨ<�Q��s��y.���&�9�u1I�Ĭ2�z
��v\�����ӈ^l�e�4|�j���t�ϭ�]���=t��7�b�H���w^ӥ!�+u�\�IWXt{̟`�Ԧ�pzV�K�dX����BM��_k\�Ȯ9�����;�m�#�Yo3�n�a�+s�ǒ���n�F"�f��2�
�G.w���N��m��(^;\Cѱ���[��S��`���z�u쵖~��k
�i��u�B�&�� ��2�cl� �ؼ�r�c�JGq`�ap��*���xo2avm>7�4A��L�,�bh]<�/Sз,ğ-��CDhi�`��h�~nL�XnL1u��r�o�({�VC�h�IK53�{5��U�cFu)�/�9��o(Ό�&�?4[V�]�+t����U��^����K��H�u�\uJT�gT�s����	�<k'�ۂ�p�h{ ���0�4ld+�\^�r��/���q�0�c�1�ԇ��hK=1��F�B{|;>��8Pe�3*z�&g�Y'�vSܥp��xc���\�#q�,B��m�Nޖ�`�釸��݄�dt��;z�Z���tg���>R�7�O�+<�#���C��Y_V��ʢ�*e�w���ƺt���rH��$O8SH����S�TǷ�oƐ�<�����~�F��їX��mu�G9H��^r���������=&R�3V ����w:#H*k�ۧ��l#O.�X���$x��7��vXJ,|LF�ǄRE-���;���ّ�#��DS���T˄�����' �ʹ�
����^��T�*�W*���l��l�g�w�J1�ldt�VD�!
r�_<�ego]�3���b���E&�q��GF\��c#�*�r��.�W�yN����K70s��Y��t���ͤ�(S����8�e�W���K5�=��U�oƑ5[À�3S4@���4������n�t<7�+�e� ���Ͳ�]4>TX=�ހ�';�c����4�r������J�̙i�dR��7�݃Fw3L\C}V�Tf��]q�z.���]�`F8s M��,�t��1�f~C+���_k��s�~��ۏQ�Kҍ�k��X%w[�[")�f�͛��e�͈� 漎�D�+�ǅ����Q_�Ä�(�&j���Z��3.>Ӄi����]0Y��E7	�hld�� �Q��vX��*���*ܧ�t��n`���K#@��0&3{��ۈ�NQ�顭�N��{N֑��N����[��x�X�����l�c�!�@dt�"w=�S�{^_���Y�{R|n�j����Y�u�IuO���ũ���8^;M�i��W+Xѹl��:�K�h��Aٌ΢v���Ӳd|���\�ޫ�5��:��RU����0S�$d�=&��`�w�y����ة��/f���9�ٳ�b�g%�/���()�	J���{G(7�)q�Rp����6+�O<�|8|��/��Ӝu���?�(Ro@\N6�r�����x]f��N�_���U�<1���W�c��r=�!����;!�b�S33]�㭎��G8���#t��J-���o���<��u&�:�N����P�p�e���k+���@������!<9��>�u/��L`�s�� z*�����q�ڋ��~�����"�<d���_*�+�
�7	��q��~5P+��k�;C*��y�@hn�R'pŽ�٥��зT�x ��=��"����ϰn��r�3�<�.8MNN	�<h��f�p����{{��#�A����hpk|�K5��U[��Q�����r�o������T+u�q=��A�?]a@RY�:x�tw��l���l��n�-�w��\ۘ|71�6�dU�
^_����RD��]p�2�|`�L��g2L�CiM��`�5����ӌ\�$�x����t7��ϝe֞�MG�*x ��B2-��9�5]�Nq���;V�KD�v�V�5{�p�u��F`�۪���nd��@�}�)(��m��u;�n�uf��mZE��AӁ;'ۇ��`�$�b�8�k�̜{A�\�@�p�����B3�{�/d(�+/6�;ɼ:�m>Crj�yRt��c���=��'�i_A"D�E�D�����G0�������pHc:D��T���s��%u�3�B�rP�cGte��0_V�Yd��]}���e���:0�뺮J�5�@G3�� ��A�TP�ɳ�^Z=�G���.�a`�?f|�p�\~YMj�j"~`��Sd)�ȨsOY�!�MK.b�;��引w�kꄔ5��+Ӈt9~_/�U��qJǠ��0��2/.(��\�ВıF��n��6dȨn@�MH��:�}9(fN�wFK�_a��Uݘ��t��*ց�<���M_y�n蹋�Ͻ�K��f����l���`��R<-�D��x���/3�^�c^đ�N:6ey̻��C�uN]`�s��2)���my���Ԁ׵j�<z�*%vY�n�[���V�;��9���$�e��������/��sM[�lC�< uә/ީ�,:����7 Mgu9WQ.�Ζ8J՞�f���Q��zڏY��2P��y'�gw`�}AV���e��Umϗ҂�@Ks̬���Lkʅ|UG
����t��+�[�T��ƭ����8Nsw
���~�++ն��
�5�����=@�i�z��P�J�۝�t:+b ��݈.�.{O\��!�T�gtv��MB����V��u���Wyv*��rp��M�o]�u��W.(&w'#���*\����j�Uc����m>=�H	MC�@�=�A��y���	�=ǥ��I��1�{u�V�����x'B�닆��B�2F�Go��1Ce�Gh{ׯWb{r�.� ��Oq���w3���h���*���uS��jW�J�:4tuѼ�JR�-��v���-娟LU��'a��e�ڢ§1AyH�";S��Xe��R�@Y��u���v�����enp�[�]F)cw L\��~B���d5!�"��/y�H�N/X����A!L����-G]�����C¼�>n���6{+׳H/3U{˫���xŎ�P��$ƀ19b�s,v�A��ݨY��i�l�g@�]
��h�����>����T�p4p�	�`y�M�~e�z�!��M�Qs��Qu1Y;��d<|�j͵йr<$�	LD��+��β>s:z���u�[�7��&�?4[�n��́�;w[�س#�0E_���ٕ~C5M<��1��΃��$n#�+���D�ԁvF�T��{�Kr�K��R�MMdܡ��2���zԢ�ӭ�R"��e��쨫�"�ˎm�9yӏeP�,Af����0.���6m{����{0�78g%�9_t�s�ˎ�����g�Y��q��NM�p9���L݁7p�xE7�X"���sʴ;����98p�^����	=�WI��ӌK����x���6a���,Y1B4�zcd�蹜f�
���eƧoN>u5ٻݢ�CP�h�r�t[��/������2�qe}G�~u���ļ7����m]n%�c�)dL�Ē�CQ[�<c[�c��[����!]~@.����4|�M��A�� d��<�c�>���{0�H`�����P]�b�:�#Q�ז�;"xv����q��w�B��`8Ʌ�*�E�
�;H�8S��0Rr�;���y1+���Z�uIYhnng�9��#\L���V�1]�?Rߦ�%��Y�y������M��c5M#5��o[��&/�� h�uHD����+�d�uwX�K����W���q۾\�e����e@�d���%t��0�e�&��f��+�roR���W�ʓ�r(�P�P�(����\��~���n��DO29�<E����j�����{�,��5��A��MZ�H\�U�'�NP��Ja�X�ce����,�u��o2f�VX�[���G0^�];��*U�uԈ�Pm��W�:4:Pz�vkF��gȅj�k��'�i��,I
K�-����ͫ%o��o Ⱥܛ��[����Z�x�⎭��k�b��wV��%���g��ъH���՞���éb) ���ٟ\���"殾�{x���e)z�ܮ�`Oy(q�Ђ�J�����O��=�{k�ᢀ�_���{�6���w'��K9�7z��'�?�,4,p���f�);��jf#��)�ǓBi5s�
�~3}�i�n��A�#E��џE���'aBl�&:b������ɑ�S�g��XM�����g�zu�bV��>D�x��*f
����`�:چ"~�T!�7�W3S��w���}sIΈ�ǽ��3�_T%�Q܇U�ON3�[*f��C4��^M�l�r�oQ����撴.#0��Zk�����i*l {*��P� ��؜��ֿKοM#�|�wj�_&6��i�e�1��^�cS��������Y9x�6	)lT}q(q��c۽�K�R̯mb��i��
����E鯥]}Q��h�3m\�-`gr�-�}�Ye��ݑU50�ǙU��/���Ժ��Z%��`D}V�����k�.E�V1oE]gA��=PaB�t��>�3EN��x����(o�K�l)����M%�v�|:뺖 k.,b�H
!���Э����.�<):J�ݽ���0%��� s�_D���i�u{Y|[(��S�\`0\]ZpR��Tn�a�(�6��cy/7i:J��76�_M7d�Q�q
��� �jP�@�2�u�qj��we��tE����+�Au���IS�����le*�n��	��Yl�SK+����]:�����V.�8b����h���)���Mup��DM���U���b�w�3Z~F�N��-;�{{։h2���:Ƭ����.�~;�#P�x&6��`ɊrL��Kc
���2����ӉV�["�e���vm6y��������I�\��Do;�sU�m�k\*�LT9.���ҁX��o�ņ����J�� �͇��Y�sO8o�"�^,|#�QLN���R��ϥŕڟ53��Vq�\jKc+w�-*�!F��$Gr�h2V�Y[C���y'�R�佛]V��u�KՕ�{*��׍$��\-]��o7M��9�h*�&I��.�Z��D{s�[ƖAUՓw֢ǲ�A��L�[Ί���9ݘ�(��-E��pP|��I4+V^M4���d�?gp�[ڴ�+u�VqK|;�P��ܗ�V���sJɰ�f�Qں��]M�N4"(Aۥ*H+}qu>��n��l-�m�����ԧ�Eh�=ݏGC�p�غ�d��%\���٫t%Ʋesm�z`W\őܒ��b͊u�wM����+����×���bv;0#5�oE�t���޻�dYմP���p�W��3�K�����{r�yBɰf�$��3�h�'�V��/��j�(�v���gQ(9\�'�Y�79�Н�-;܍����þ�l	��LZ0F�t�˱
��q'/�
�T�6.69jv��Nu�yWAP���H�����b�����J%6�?YK�XgH��fc�)���ަ�s	��Ҷsr�k��ɍt�� -�|ƪ����Y,���CUY!�"�#JE���bC�5>��4s#�,M*\���wٓh��j��@c+v�ʊ���.�Z�*wɧ����vI�ᒸmo!�=�S�Ww�X���w}��k8�x�}���m�����3S���KG�
�;6Ѥ�&�|h/3�C�1u��zxUɣ��C�����Q�N��kWu���W!��j�����\z�� �Y�<�%��>���m��`
d�;�sR���E�t�i�] ]�K$;/)���^���ηZ(1eƶ���q����5�S.#p�VJ���I}�Z��+8V�p6�G���Z�$����L>���A���`�/�M���n�ňp�P@����f鼺��c�Q�7]]cE���{
!��L}�XGTl���y^b<<҃�/ה��t��U�t5�P�ܴ��h�;S�R��}�.m�l��wSM������巻k8�N����T@��ҋ�H�rY��E��  � �e���[l�T�`.[m��
°�2��Ԣ%J�d��m�EF���&f9IR
R�H�j��m��[`ԡX�YQ�%�+AƢ�\�f V3,mF
,�e(U��
�DQ��b�E�������b���J��1��h��n7,S0�Z*,PUZ�ҬQaU,b ���fT���[h�1�㐘Q�P�C2��Q(�F��J"���TQ
�AQ*ḙ�1�)�*��UVڥ�
�*�W�Ƞ���T\h"��,b[
���AlVլ�m��V����5���kB��DQa�2�m)Z���h�5J��m�Ŋ"�¢*,Qh�DIV�ъ�*�k�*�X�eU+R���
�0Z��^��=ٙ׻_:��4��������$˓H��y�]��Å�Bd�0�V��&��g[d�7Y/���ei|ћ9q�⼐Y��?#\ԕ�H*�["$�������hP�;N��hJ��]�S�q���UC�8��������}�ڳĕ䩹��h�N�!���������$��
�΅��G� �&*O-�N������i��ߵ���i��3!���P5h�|a�t�w�0Ӷf���l8��veg�|�C�]$O�> �t<]1}&سD����"4}��k�6��_Rc'Fs:M��
������$x�U����I�+ߵ�c��B�~�&��8����fE�Vk)�
���P��f=23Wϔ�JO�ucM,�G�E���Ou�4�$��t�'�AV�<M$���=�[���6�=�'��J�Ϟ^��H,���VbJ��ɟeB����&{N�zd��Qg|��8�Z���M�����;y_�$P�G��ދb�d��`::�q>��|N�b$�ho�d�S>a�{�哦bAz9�j$��1�O��i�jN���6�R�9�Y�q�C�
�_W{W�.��U���r��F�����m��;N�vmY�J���Z��J��d�ܴ�_�CS�I��&�׺/WLC��i�<v�Y�ϲM%d��G��j�^�b=�/Gt!5�:���¯=>���H�
��y*4��v��$����v������=M�C��H/�Gt4��yd�6yC��O���ެR0����
��T�}�M�ۮX"�תk��O���9��[� �����9=�f�*A����&3j�Y��dP�P�&=0�����x��4�Y�N�|;��H*�n�I��!RnuC�qC�Htyv��VJ>"=>��b�9{�r�бP����?vͫ=IRW��M�����:��$�Ҧ��7�+Y�%a���%d��d��a���|d�1�]�!�J���ה�Ag��wC\�m����~��w�bv�[�E�u�g��� � @��C�V? -C��y��:@�Y���C�O�ͤC�<��<Ci�5ޡU�$�����mI_�L�ވi�_-Ld�>B���|�=�������شi�%y��.���;�בa�:��Y��,b�,%�����}wx�a��׉�xA�
��nr[�`SY3����܋�ܞ�)�2���u,��{M-z�H|�v��y�D��4*g�cj�]V;i��ެ,�a�Y�bp��ݻ=���+$�-s��U�{�]�秜��t��=C�̠z�� �<�̚J�U��ɉ��w�0� t}�m��bz���ϻ֠,�Y�u�;�6�Y;��C�1������ ��䘈�ל��}⽻�w���'[}���{�H����}�O���1'^Л�W!�=C��&u�2|�l�쇨|��;gf���xɸf��t���^y������9�k~���o�5�v�2T��w�ISI<B��s�2z��SI���IY+57��?$Ă�:��4��+�]!��!_S�;��:���1I}�d�Y�%g��~��x}�#���`j���8�'�˗�)'�W�Nk��g|�*I^��5&�M�z�9AM2i�&����Ax��j��jf��z��*T7:��z�!�Y;<�I��.�Èv�����x�xW�\Y7�:�ߟ/}c�g�+��M!�J��0��p� ��K����m'���{ԛ��C�;30++�� o��L���d��H.�����cWlꆙ�1#����K'��N[���~tg����>C�bu�
��OY�=OP�N�Tx��9�St�O';�_2t�Y���d6��R|�;�4°��X��)1�1�:��i�d�������V�5^�x�f�}T~��� r�=B�d�1����!��<M$|���5'�r��Rz�OO��i�N����C�%d�u��6ϝ$ă��jE�C䕚�p�c�cK�?�bNS�]�+��ꅛ��݆���1[�E��gl��
�2m�v["��+�y�N�X�I�k���N�M$��:d�Y1��T�?}ϵ:H.�5�GFu���}������^��:M��*s^䋦q�!��;Xi ��4�\��1 ����4��J����4�W��;��I��3�/)
��+�߰�&��`c;3��M���뤙z�9����:�>��׽��^s/�����J���~�JAH.��Z����XW����!�cS���m ��<g]�ĕ ���8�!�ia��1��Ax�!�)������:q�i�����}&n�!nY��Eoi0<�5R��}�EԚ��!x�EZ�R�L^@�ۉ����|g���ߤ8)�/(�Vڌ�����Z��2ҷ����w�� �K��Y(4n60�b�E1!�4U�nq�r��9{"����i/F��@" ��ѫ�aXW�l��{�P�J�hq1�gyL��}I���1XvsXI�/�O�.��0���'���Ϟ�x�'���Y���T��7ߎ��l�'��YW�7}@>�#ܦ4h�H�a��i�g�bW�+'U�$���&��NЯ���P��$�8�TY=k6�Û�i=d�Ǡ�d'�W�nuC���C�����j�{+pe�_w��$X���P�#�Gz�~�c17<�b�=��3i�O��:C���R�9��q�4ϐ����@T��h�:�6��HbG��V��C��|�J��+�xy�د9�>�2ND�[�OG��D} D`��׶��3��K�����MZ�!״�ϙ*V>��*AT���0�8�a�
��(C�>La��w��t�Y�<βT1%H?tk���������οU������"$}�]䚴���=�P>J���14�ɉ���4�+7ݟ!��{���4�$�q�|Ο����w`g,�3�s�M$��}�}��;�K��=N�S�\��!��"8}^U�>�|��S��v����+��CJ��T�=j�$��lhx� z���a�v�&0�d�*��<LI�T�!^���d�xɌ�eﮏ��y�w������:���!SH��+;g'|��AO7���`):B��;Ԙ�|`T=��tM��SL�K���2_���Ă�M����m ���Pơ�z� u���Y�3�_y�����_�����7��4�����3T��ğ{CP��+<C\��>J��+�����H(p��46�'�I�4f2]ߐ:�Y�>IYX|��;��%B"���@� >ۅ�Nĉ���_���s�'n0�6�a�at��z����~d��'I�'p���C�g��B�8ʇ���aq�Af��jM�z�%�&>2b��c%W�
��q��+��_o9��3K��߻�~��׾�����v��T6���o�
ʓ��0�|���/�7�|����|���zI�|��{���O���
�B��Ud�+}����N���m;a�%�h��/��˥�5��Z���R��Y�ۻ����+dչ��}L�k�Y�ս@���]L�v᨝�u0�Z�����Z�hʳ��`��ov�q�Y���\�����r�s"M_:�ݥ$3�V�t���Ǟ�(�^�,3���z����%b�Au��D�]��gJD��ob����1�>��2Ɍ�2�;Mꆒi
���SO��L��i1��'ɤY8�t�wI������\)�x�~S�MÝ���@l݋��7:��<ʮ�>��vo��
d@Ж�HE�A+�e�������X��U�FvJ�أ%6�>R/2��m�.��{2�P�U�'�^$au</����tMx]�����&��������R;�Z�Tz���� `b|����>X��\3a_p�<���k�^0�Վ5�y�ó3
.�op�;e�%!0�:�:ڠ.n@��l �K�շ4�h�ZH�O9�祜�����o�7��1�	��4�֖=IY��Lb�5x�7U�n�K@
�{q7��e����n����(È*XVc0����k:ܠ3i�0ڣQ�zvnڱ&�	�զ��׫ݮ�5꾠��V�j�x8}����bp�b� �l����s�`;ϻj@cШT�uRZH��������ł{M��g�,@��j����`�����9�Sk��.���\��rw�!Z���2�g���+�o�ܴ0׷]�1}����Y�h�^x�p+��8�n� �(�qa,�1�)�j�T�݈������'h� �v�����GYKa����oh��*�Q�qS���/��ˑ���Nż��nq@���9����Y�t�)mh3�6�#�X�A�3c�=y�o`����.c�T�Ц����V�`m��]H��1�q�gNU�5��@zHE��Y��8}G�:GkY�{\��*�ܵ��V���k��g*]��9L�;���_Le�P�{@R;�kpFiKK�u�Φ��P��f���dT\�,\d��~]�S848e����7;��jt�^�L���"q��ݎ��S�qU �*�
0��̪��B&)�8���h��y��c��XJ�$>����_�F<~(}�7�%_#_6��]ω�Y��n�b�<��ޞ� f�Gu�K������H��3p��2��j�hQN�A)Ϙ�7ϙ1�aX��|e���x*:���|]�؝��)�ԀD�rYྃ���@7�a��;r\�D[��k�@�9������K\�'!�Pp�܊yUA�㹐�N��BWX�w(�en_q�H��0��X�h܀P�
�J��ų�f�M�w�+2�
�N�}�}��WC��8����J�T`VX�:��F�3�jJ�2\�Cj�1Y�c阠f��Vg��1�R܉�ӼF���(���1���c8ew
��ں������/F.���6���Z�k�lJiG�vn��8ӧ|EYs���mct�9X��g0S��OY֌��Nu�<�҈�/1��q�-�m���)wWh�.��9�Ϲ{�@���2�����[���KU�.���50�ʰ1�hjq 9�Q%&�B�����$0����Q�2x�Ʌgo��uRՇg�q)����i��=5�ݳ`2�p_Ϫ��p���7�L��]{�8i�y"6�V�\����-E�f�xFcȥw�^�g]Q��īQ�n���γ�~�p��$h����F:������k��FS��*�c���}�i�-�ߘ��Z��=�	��lmw�?z,{{�v�Mf�	���k�F���
�mE�|߆;Tǃ���V����r�Gu6~���s �/�9�1�#7����]E��|>�·_]8;۶�T�(a0��s(sȍ����c�<kk�I�V7�d�%����
�hC��{�&�*��e��UvE��Ws�<��ͪ�����ݕR�WWw=��[�T����cw]!���yp��x�H���?b��t�V�PZ�����y�(��rZ�ŲV?���W�_Trt��rj6�N
������B�� $DG�s3�赁��2�����e�#mCX��m���T[��3,���.���={;�f@�[�UH�o�HkU��
܁��F) �{;���R{���d���Z������fJd��W�\�y��u�묙>Q��)�k�-ص9pj�͔�!�r�ňБ�/�}}�
�gC�q�7P�vw
�wDLC�v������u��(ě�����ȸAѣcz|ޒ���-�R�w���z=iҷ0==�s��Y��b��/���U�Q��r�R���x�UO�������ۃC�ճ3��f�WzO �6�������u�L-f�M�a�Q�d����~V���
�c�c�	B�y����n�oalT�Hz���}���c9 �a�E�X��6��ݨW���nX�5�񇔺��Z�$1V_݋wD�W�4�+��<���'e��Ęc�a���M�\gt�q95c_���F���17��<]5́�4�x�?g��7�+��{O�rN�YSra��e�b��	�º
�!�S�<�뒩�k~�)bW��m?{�g#��
{��5
-�2L��<`�^��h��{xEQ;<-��h�iFԇ����)鎙t�-2�zu�Y�.�N�:߾�̸���jҳ�g����Ƴ�~9~@W?�!�Γ��=c�yêG�����~��/�B���ʥւ����]��?r�u���iշ��ĞO�V���0��I�ðyĖ�r��֘��n�Zuܫ{��
�8�妖J��ow�t�԰�����4T;.j�|l��!���8�7g^<l:o�]-��}S d�|��uf��N���'|;>Z��������a����O�?<�M�>yP*���\kW�xx��e�<���vu�L�dS�8}X/���J�Mp�"����q�9�K����z���{Hl�م��Rӑ��7M�r�3�~�6���k"��k��A���q��٦���h[�c�E��jY����S��8��0sSe�eN�ܵ��{���`�r��#�-$5��{F�(j���QA��C{\T��dF�"��wZ�c�JH�]d�W)D¼1-�fT�Ϡ�͒��@A�vV�������.*} m>q[mj˱��z� C�ȑQg�EBrZ�"��:2�4�zҨ|-m��T��cm��SQo*$C��4�]4�y(Ajb�I�4�܁S0�e���$8�R�T�UJ����$M�u��	��&w'��Z�l�l��K��۪b4N�����ĕ���ϩ�1�b����i�����Ѓ�J��K�0��8w�V���I0���F�,c�X�u����h�܄�L�s�+~V7=]Y*�}���-O�Ĩ]='6,`����2�&A��P���1�ҹ���A��C2�aw��[#+h>����cb�5
�5��6�Y޺�,�i7J�+�I�2�wr�4+U�[�>��}�W�~�'����ޱ��[���ڳ|��
y倧�8��^\��?����7��l���v&Q��R�w9q�I���[fU+E�n�?��XVo�����*�O�T�����5��[t����X�b��Du}�/�*�X.!��r#�9)c�R�k��χ /�ߦn�w�����Ԣ�����R�����&�θF�u�F`?rj��L���qEYY>U��7<�RhW㾣`9Xc��AIzF�!���l�{0��b3�s��ף�5��O�b�bOk�o����!ȝ��*9�Ο��gQ��	e῵:�Wf4!�b�U���k(]b�/��#cV�n���9 :T~~e% ���+�N��W�AL����'/�ּ���E2��׹n�3_wl�<5¯��?C9k�۰�W վ<��M�8���kz�ZV�#�k���d����j�Cx*�����*˪��]�B��[].��m�}�;*�ر֞2^���`������PB�쑂��dTCt���2���G,�����Nz˾��=;�J]Cr�S*��u0{����@�N�1��[�3;�3�>���״�i]�*�)�W�m���PLf���c8P#5���f胟p;v��7���Ž�+�#��,֩4���SJ�W{�M��JjJ��C.tζV�7����?���$������/05�O~�?Ww\<���A}ZbvF���R!9�Dl)�P`��Ŗ���T�5�����J���d�s ���^���p_SZ�|���ew� ��� �ˢYg<�ĺ/S���� \3�(�S��CF��◧p���
�U�sO�*���#YK�?^���ݜ��ݏ��3��h����n�s��18X�u�u��<%q��0�Qw7=0�T��ϝ��a�����T4�%�����s,0��F��d�;}���tB��]�����S�\G*�O2C��}Z�O���Ӈt9W�:��-��k�$t=�e-Gd�������b�*�`[�Bx�y�"��0T4$��̑�o��C��|�R��!��Fݞ�:��n�i��F�;U�g��}��K�����F��[#0�w�7��y#^��K���=T��v}*��U>�!��}�W��s�ygxy�EF6���,��vl�^������fxՊ���݃�M�c�Lpq+F�ɗ�q#6#U6~���|uDD�,qq�>�;�5N�j�B�Y^%�qZ^�h�7�ޱt�մI�+(�+Fq�&��ض���{q�f(�q���!p�v�N�fGwztٍK�Y�l|w�Z��B�R}rb��N%�ٴ�+��M��Hѣ�Jɮ<�s�-a<**�B�w;r��v	��uI�����xk[X<���n�:şr�zR�#������gv��� 3i�3�7p��I��j��1��lT:��Ѯ�J�g
����|��7����x6��4B�G|*qn`߭0ۙW٢�v�=/�5�[�[%���"�()A��@�p�뽴�n壤9��)0��۽�-���\ξ�N�欷�a�g��kj|�	;��+J�ѵ"�F��j�Ү�
��$k��w%�զ�<�f�x�����6�[�ի7�H:6*lwi��F�B��婸~U���Cxw3�kR�[ջ��4z̃�۴�Ǩޭ۫�"�
�v�ƻ��-,ͣ���M��V_��yVo!��ם;�A�`.��_-��tG)[�f���v-�L��2�u�B��Ɩ����[��E�t|*�lNa>�g���U%�ը	��C��a�V�����϶Ȭ\s�[����k����w��쫷�N�_3}�Z`�$�|:�aK�+P����i�Ж��+�6/��c����m�+��N݄��:�ضN�NYu����E �n\k��'� ��׺�uK�卋<��uy��<,�Ol;���jS�3��xh�tl".����'SG��v��L�.��Հ�Y%S���b�4�Å�Ylhu%S�h�᠇���_-�9Ȇ�YӰͺ���'2�sɱ���;�:�[��U�a(����	�S�W�$af�r���-.�<pNT5`ͽ��xtG�����;%R��:u�E����G]]Y�wj��fO�6�R;Sp�Сy���C�{E��gJu���g_(7�+����k��%J;�@����X�Ď��ww�0��2>�U��|�Ř���Sm��ٶP��{Q
n��SA$�R�J<��j���(�e����!���X[���ٱ}r�&ޖ�]��G��,X�ʙ�%s���׵}��ϛ[Kgq{#%��	7���eC���3���X�g������ͤf'L�vl��͒sOm�੥T���^*�1�x�T�>ڶ�T�YȌڹ��V�F�;96�!K�S㋻�Wf�Tu��H��Sf��e���ŵ�X�R�=�c�NS7�:=x�h���7J�gi��-��p�MX)�V���)Qξ��劮�&��s���YiZ��5�3�w2��^��016���7k�`�:T-��\8�:T������Ywux�;�B��m2(�8���;������FۗL��� �L�:�v�͚�:� -�kiqs���INZrV�n�u�C*�8xT�f���NS��ٝ^�F��{�\m+DUVEJҥfS2�����ج�YmĔV
�L��TH"���PF�j!Z[
��R��FڕR�Z�%�QTX
*"��%����"��h�2,J�b�j%iU��*���-*-�UU�Bŋ����[`�Dm�r�Ghъ�A��E�[Zŋ�QTR(���s0�em[`�kX��X4���R�[j�,�PFTUb)n[�[eU-�+*--�� �Z�c6��c��UE`�P1�UUb�T*"("��bW.e�V
"VUPb���Q"��"��*-k)s%AƊ(��m,UX�QQPFұEEA`�JԨւ
�1FT(��Z�-r�X9lV(�Z��cR��AU�QA[j#ic�&&(��ł[R�Uj�TQ)*e�,QV
���UV@��|><�����^��WQr��n󆛩��n�ԕt���m&�]��s�z�J�d�J�9M�x�����z������U�xQ�]��=;]�����Z?��S�)�7 _SY���f���C�ʲ�'t2]�ra�O�޴R�8m��EQ*�G�p���l�S�j��R�P+������5��=d�y7Y�R��ǻ�h}�P�4���X�}HhR�=%Ā�ә��>��ղ7z'o:]��B��-�e��4W��_WǓ���rk7�NVU��[Y|i���`s��Xy��-=s�k;�iF���/j״���X��8BI��]H;Ckzv,�N���go'�����*�����*��>U�bʞ���A�޲��s�)ȋ��
ʟZ~��=��*���?V�����z��K�T׉��>�H:�^ÖgC�y��H|.v�¡��m�E����! ����?��o�v�Q�e�'쪧9'�o:j��v�'�Ň��6�6bG>���.�l������_ı��ߠi��C�<��]H��g6b>-��Ρo�T��*]�ew�#֫�w<. #�'T�C&h���C=3�����x�����.\�˷r�u���ͥ�hr�,F��i�z�+8���v�����bW�h[��U����+>�l�T){2��@`y�n��0�Vr|�y���u�ui��"]�&c�V�})�/2�es�@���gAˍ��6�n);����ﾨ���d����R��5\+�4Ǽb�S��^U�i����x�gU}M���v�ˋ�"��u/�F��l&��B+x.}z��;8��=�ʨ���΂���=��Q�����K���Q/'���Y&�D��_�0�؈��V���n����#�b��L�^���[�a�I�ϛ�C��TQ����I��3���\�3���v`���ݳ�Kݎ\�pO�J֜|�8nE:ѷ�=��_����Ar��v'��u�Q�z�|��L��U��y�U����a������/�r���,h��8jj��� J������+NMo�\�ؽ.@���Eޕ�bB�յ
㊥�4��鸄刢��;E��0��ӳ�mW�G�yD.��Yw��eOR��taC�kv����@��ҾY�m���Z��h윻eտ|���T��:��RHk���l�QS^;���Aǆ��3<*6���U��J�lܸjHڃt�!�Ʌц%� pY�J�T�ٿ�\c/�Ps-f��S`*�Y��jމ�M�G��q��75�����hw>�ށ-��k�c�F�j��86�{_�^\�ч=W�p\G�f�Քr�5|޼}p��&l]s���S��*�����X�������eݝ=Օ1{����N���eE���������5_	�ޗ�KgDhVt�T<Y*̣̖�I�uyYU�5]i�p{{\A좞�%1�]�2��i#L\7�l�{LA��5 ތ���`JJ�nB��}UM{8��P�K}�DsOjJv�/��`�)������{͇ݬ�� + ���9��ڂ�"y`߽��$�]�4[�o�:��S��
O鋼w�_ei��TG7t�:�ᾇ�`�S/��ů���t��`��u+�\�6��aN+�<���6z����˪4&ݸ ��w׶��:s�Ş�7����q�3�h���n�:��xJ���G>�븯7���m� �����-��i���yP��mh���N��k��y�)�sB{���zӗ˺A����'�@W�X�v��\�H�Ǧ������uZ4��C!���T�D�k�|sl-NIߟ��5��r0z��\�e�w��2�
{�t�ݢ]�E���=3s3�lL _��}7���:~�0�MƩ���^��3�"��l�V=���ꗜ�Yu��y�\l۳kP�֓`���x�siP	�d5z�́n����7I.�]w���{���|4�9qG
���Q�Wm�Tc��\c�Ai9,����[d����x�^�Q2�Θ��ڿ�hݽ>����|��]�\�2|��zy�����Z�ꭣ�����}_G�|�]�un��5�8���q��e!RP�i/i�d�����J�`�C}^�>{�kZ-���tߦo�͖ǩLW���e|�S���z� �<y�}X�S���{�]{i@�Fu�v�<��1=�r�?'o!���U���A=d�d})R'pwyGv��u���V�OD,q��C��G<0E��]RD��Bρ�����<d	�r�H%V�=�&�;�w�雲�L�dm|�n�-�Pٸ.�A�N����D"T��貃��sr�JY�#�x�R��H����<�g��;�gc�W�����Fd�>�:�9ˡ�������7�s]��Ҹ 2��\�1��C��Q����2�h�Uʝ����
o��c�.ݬ�:�>kyV@���*e9(��Z/)7]v�g�����k���q�*s#��H��Н���Ç��#���.����䖎��}�r�-�ɇ��N�;P�]���4K�[R�[{Hw�c���Y��v�:��6g���/j��ӓ厺̿c�'� �<͡Xi�=�e�)2�����
��%�h���5p��̑�}Gv����镨�W	�B��z����yYY`.�s�9R�D3�3��_��-NYK�NoW-�uo"�b��d�v� ����K�]��x/��nf����71�^��F6(�Z�S�#菣��՘�c�o�z��i�vF�  �����X�=�ڠ���VI��H�8�������pW�u_V-+��ܖ�T���{2wLF3ZT���`TgӐ���]uD���y+��'%�!�V�}����H�}�+'����vz��*��0�����F+@���ȳ��]
�)���aHW|���]9��G��s!��96��V���%|eZ^��U�u����,{��֠�W��M�����2�}�ȴ�>�
�p�ǖSpMg�	V�pu᾵1����`����jlΌ�Ɵ�_��� ,����ҙ�UvE�����ϖv�#mؼ��/�Ѭ,������k��vԲ�����=|."^T1p{*Q@ ��x0a��1)�NE�W4��d�t�m�3��Aw:�܍�H�l���$s\���ƴd�@>���F%Z��GY<x�a�}�Yq��2/�`�9���ƯxT+�:ncD ��*zO'jޛ��|瘝k�b�sW����WH�2
��S�\=��G���*U���uw�>T�J�M��o]�T��m�� ]���Ę���"�I�ܝemv�c%L9$Ɋ�Θ�t�E5X)d���y��\V��;��TJ�xw�F8d�ޮ+����ͳOP��e����2����"���� 	v���Ot��������U!�v���f��LB�y��ˢk�����M'��|�3.��g5��.�f@^C�o��)��MW��=�*�u]��'��h6���-W\VO�Oذmc��*}�zƼ�P��ts6��{�%f����
�� �!MP�r���<jU4�7,�=�\���͒�'q\79�j���S��0A�	��;�qS<��()̰й�8�	�2���r{�xuxL.[�gqu-x�WƖ=xi���i�?oS�y��d��S��Ӕ~���o��e�fx9*��o�E�h�R�X1���8a�b��pV�R5��˸��7z�9@��m�X���eC����������X�)U{�]�V{.�CJ�E�D��_�0��}1����}3:�L�<��wqhW��\5S����}�q�B��*��X��%]e�5���m���sֹ��@�qj�p܍Jޜ��0�\V;c�%���o���"T��vRVwt���^��n,�ﻖ����Fq��g�#�ʫ�(<6ܦc����)u��u���+e������z�i,�:^�ŝ]��_CL��8k{Xu];�~�[IH����4yn��'3�qQ�*�����C��a��q^���o��\�<�dYy�����M��7Ӳ˻�2���TO>��n���MZ�8��Gp�^>Ȕ���>�t&]k�"ֵ����������B�(��ަ�Hg�Q�'讨����:�atGL���0��L��;B���ns:�T���e�a�ͧr"ŗ ,��Q*����\aC�sv���
��� bcuX��������R��vR��}���<��i!�-��7��^�ُ��[ɸ���.�����*��:��Z.w�xm��b'��2ad-��BS*La:�� ��{�y��2���v�!r���΃��w�+��� T\�<�:Hp?j����J���VXu������&8f^��\İ��3�V�n���(
���a�W�Ds��O��{K��c���3���{�9�@�	�Ĉ\�M�@\[��"� 7f���e��0ǹ����x�tc�W���n������k��a���}�hx�}����C�hI�Si�Ts��]o�é&�B XH|cNK�*����W��A��@N���:^J_5W.Zr!�ܱb��p)[�J���h��U�>��xO��e���}����|ݨ�}Ամ�V���"RW���|��sR���x����"X�c��u�y��NRt 9t�̾�#�u"��Nݩ��yU��#	n��ȡ;��<�4���k�꾽i>��(���o�M|PJ���<4��Ƕ�(Y�����艚5���{��&+��q����}����;��ہq��ͫ��!B{���^fW-v.���[\ �� dqC��^�)��ބ%_������V,�{��**b����0S�$�[�)��f3�ap9��C��%�3S�XBƽ�<o���T������ܕ��F�ł�U�z��Ο��>S��\K/�)��m�h�WP��sCn�9׉dƆԄy�(�ʲ��q3`Q�#._'�ih��s»���w^�;~0EzUqN�:]�EiIX����a�LS�� ;�kU��o�;�|+���c:e
�[���+�(���b�9���W��9n`a��ڸciW���	J��j����ݼX�	�{Ԧsx��F%B�{Q�Qu)�q�n%d��#!�f�ti��T�Y)�Ҩշ�c�d��O|O#��_1?Vh�Z�!��;���z4���6�^; ���[O �\�d���2�(|g�Y���9�5ɫ���,��.K��;T�Wu__^��؇����cJ�/#��h�t�Zq1�[F�rVE��va�^z��| �.�1�����l�)��W���҅7m�rQoN�Y���d<��Yi�ڼ����nB�J]�u�NV��MÏ���U��,#�7�;��U_}An�%�{�l���P@�, ���(�S�y�6���{X<-�jd�=�o*co�G���H�7	 ks,X2��>��P.��`w��<JF�^��U�����v�,`���6sEw֞'��0z��8��s5>�N6�!��[d�s�"�ÿ-��
�K+�T��kd�l��{ק�m�}�@��T`�_j�\t�29�2w�}Tf��ܒ�۪<v�j-6�o�[��w97�7��'ޥ�u��ٽ� �t�J����7�A׼����5�z֟G���gR�-���F��\~Y�xX�^T�U�GV��u�.~C���'!�vf__Q��5ku�"$>m���N1YsXU��:�5�7�?<�ň�T��9I4:rg�P��W�4҅��ۛ\.�<o�c$o�YXeS_d�*"�q%�K�F�+v\�1��� d�q�Mr�?8�ѧ�w���S�Q���~��#���n ���*�I�o���E��M+�$���_���Z����AJ�����`�n�kw�|�sU]�}(Jh��"�{9^���Y��X�@���p.K[�����1yL���2Rь�[6��@V�܁�'j�䇕�׸@�9�S��z�a�U�X�w�ܟQZp#�,^oc+G�M��.��G?����4��;>��>ø4�εЫ��/n��5���2U�'����O菾�ﾈɐ�5��7X�s���~��O�k��,���W���f���vJ)�R5�萸֊�ĕe�Y��a#���(��2�6�#W�_W'Id�S�8*Z�6�	�v�	�O��y�ڮ�D�# 4l��vIz_�s7y/�E��
�'i�nc� �ټ��������=O���Wc�rX�0a	0t%q\M#X����������:%�ؖ�%ۙ0=-��U2�Vt@ߺ��{&'�ɉ[1#qK��>�u8[Z�8�����s"����+�t��Ď���&)1\�S�7P��+I��N'�p��iU�:O�	�����u3i�Z���b9���6��̋f�;�i�F/�c��W�'\���@���%C��׵6\��4�30����C��m ����6v&s;T����ٯ�ﱿa�F�2Z��6�ea������_�<��\�9�=**9�ȓ��`b{ˡ��v͙�@�����ڷ���WmEaٗ�g��O��V�Y�&�}v���	�:�nt�h���CJu��*T�SbG��êIp��Mj�+���V�v�>P�8b�Ȳ�❵�|��=٧m;��I���k�ui=xK[ܝb����3��c](:C��@M��*;ͺ�W�&⧴l3�;lD�
y�`�:�����
���������R��Y���8@(�Ǭ��L�ڴ!ݍ�Ti�x;ybZc��WO����%eA8
�UJڌ�wMf4.��u.͆&mlE��kq�d��dv0<�8j[��m�Q��-�Kv�����έo���J���TX���VV��G��*q���`��*��.���3I���0�[SU�H|d�������y�:)b�́9(��-�j���~".{z�M�'i?be���fJ�o8��f�1��-��K ���#�{��|���]vӣ귥�^N���T�[c��jOh�N�x�z�b�c�Ș����nѽ)���h�fTj��j1�C{�^f'4V�����|�/�����t���.`=�g�F��4�f+XjV��x�d��..�1^R�2-r��ë3]o 3eV��S���i�T�����<��t��Ӧ��஡�Y���N�7x����goo�R,x�1�P/i�Ć�zө��uٔ^�+��3�E��f|:;,�ځT�Y�E��8
;99+��D��t�R�н/h��tzw���+��N�eop�X�)I\���=�O����ݟ7z�u�S��])]�� 0)-��un\}q"P|�����S*[���sF(����C;V��R�ui���<�:�F�����EX,�h5aaO�O��+I���퇀���mv7R����]�waf]��FpѤn�WS�ޅnZ�yu�K�a����Cx.����zN��;4��J"oV2���o7��̬�kL���*5���23���I&e��k�����cU�ҩu)p\o�y��Ѝ>����i�x���u���t����lK�SK�]�b���h����2�B��)�R�^��:M*.�5862�}�D�1w:�ғCzЫ�(b���4�V`��O�}r�1*�ۺR��{��nuj��wj����S�P{g�2����x�-�L q��u��c���hr���8���P���/�X�(оs�B�-��Nv�Ū��Wצ�P���.i�	�̬@�{n�&�Q�k�%N�ơBV<W��X�����bp$mݲ-ʣC��J����+
"�˓#���G��/�O�*���0p��b/�U������*�t���
h��>Du���ܦ
�/o�6/��6�ӣ{ې�$$`q���N�2R$kU�g�����	wWoL���M�aD�TW1�N,�+�3��#�Zl՞�ބ:3V���Ԍ.�u���U�c��A F�F �,1��** T�V���T�fZ
U��(
���j1da(ֵ+�" (�mEƱE�EEU��PPb5�[J+AT2ت&R-Ub�+%j�L��hfU��E��DF+i(����F6Ѵ1&!�X��(�X(��[h���DX��ZQH�ֶآ���R�SU(�j�"�VEQE"�*�r����R�J�UA��+H�V�J���aZ��"����-be*�*�"�(��nU`������*0EA��E�Ub�±��T1��c(��Qq�U�(�X�s1���T�l(��)�QU1
**��3$�QDb�"�Z���TUU�cQX��ZT**�DU���^��{�����Y"���U��Y2�#|�O�|�F�=ϐ�:�,�{��������9�������9ZѝL�i?������Ք�8�M,��7I���Ȝ���ӯr0�^@U�\"����*����R(ܕJ��F��<����O��Eܴb�C�9���{R�(��
�>�Ub�RU�_�Y���J�?c��a$�2��.��9��!���Q{j[U��l�<����./�V�W�o��[�;5`Oٌ������U����]I�9��U_Wt���k��vEJT��C#�Q��KL���ࣵ���qz︋N#���"��ꈚ+��&{�[P���i�?1�n�#��0�#h��=��j�-z�3�$���P�Ϥ����UHʕJ/���]4�m"��X�3�P:���.���������W��a�T:ßT-t�tr�8��V�UQ.*�.��{�Zy�_�F;�8ܲ�0�_r��zak�j�qU�N�����)��١R��y�cy�]�B<a0�vN�'b��v�j�j� ���2=N�n},��y��K�7
n:�ȕv���R�Z�[p
�Iݴ���o5ya"����v��bP������+�$@䥰���r�r��6lZ�e&�F�Snvμ���M�bʋd}I��c��]71Lg���9(�F�wr�-��yԲ�)r����Q��I
���Grq�n5����ǋ=%�K� ���E��UO�#�����ՠ����~��ʴ�a�x��+�ꔓ2�}җ�t`�^R��'7�i�y�y�ٵ~�8C���D������b�g�O�J��^�mp�Y�uc֒����\#�K�:���h?=)v����e.�{>�gǕg�5��vf^�����:�����v��9�q]E�U����B���O������Y<_��v뢻���|6bݳI�ʆ�n�*��ڌ8A�&n�Z�����_:�q���q���b:�=�������w�����զ����n^{�"�uc�U��jlS��r)��x����qv���;D�?N-Z��j�Ò�2�kV1lY|�����Mk=6a�ۭޝpA�����OW[�:�n'��l0�w���5[��D?m)��4�:�\u �X4�jiGn�Boh��|p-�L:��usC��?L螪Q�כ����R�I��1ss����X�5/��T�����1Z��u���zT�����J+.k�M��Ǻ;߮�f�m�8�����>��sb���,��$��uK�N:��Q�;���Ճv#�j�]oX����g���C������=��">�>�X����y��u�%���m���:n����C�0쎸�K"�E�\�N���O�[��
}��j��&Җ�*�.����pyY�#inWJ��N���ʙ�;��.���TV�q���qS�5veGV륔���U��W)��/B��ˁ��.��
������v�&�ܞr4c�5�7]��s�w�<�C�+D�Gy�Q����j�{v¹��+t ���!���܎v�̶;j3��^5f���K9����ZR�>c)r�*&�Ҡ#��K�}���R{n��M8|������P��٧����Vu��P�k��nE�N�I�OR~���\K���v�Nq�8j��NGfO]̯7�����Ҝ�|}_{�(��oڠ�巐����X�7��bi:B%fE���ۼ�|��o�BB�=�~]K۪3�GS��C}��tUoESW"b�H8�br���Ed�Юf��K��,�r�I����X���,e����z"����Q��9����wW}��ر���Q>9V��9��t���A�i;�u��S Q���mdR��w{��舏��\�qj^��>��6���ȫ��tU������י��.�%��pt�"��l���
q�s�k��{�if���/&/�W�qTY|��\J�f8�w��Z�\��m���r)���7؝�ތBUB�H��N�>��Cf��Z�OGqw�9�.1�����H��ج��7)(���P�����E�+��m�ȤM[����t�LE>O
�ת����u�΂��R��[JԚܟ����6�\����g��s�:^�{ܗI[#�=&�R�k�L���Q����Jߢ���q<�	�8�Oe]>��Л��W�k}�9����5���o>WB��C{,�*y�|�G,��V���z���z�+��8�':�)�V�-+Y�
ڄ����Ř�!wY�����9ք�@� 
�K��k�g-�s�H�O��P��u'��O/nJ/������˂��ʨ�@��`��{<��Ssh�y�FV�/}[���ۮ�6;%�X;�E�e�+m-�uV�|㫨�T��oy
�r��F���5�z�@<V�7�,4��,m���� ��;(�'���	ץ�m :�n 5[����v�[ݍ7M-�+�og�W�}�}Jg^ݝ�z��^�Zq�W�%%��E����.l��Mܕ;�����=��2�Y���3��J^ߊ����R�d����m=�;I�8��}�s��"�E=���W�e��}����;��u���/��'�����iŬ��w����s ��FA��l�6��.+]����V-�]K���֏)�n7�����}��G"�o���~~0�y`�*�e\��{R�	��v�D�o~�N���E�)[S����g�f����n�F��A���ߔ�	��q';\��Z���Jʈ��\C��[��ys4����v�cp��K���kKnE9�1]΢�*���ڥTiO.5��U�L��.[�5d��j7ϳM���'��[qp~�蘧�^Ju�UDi]�����E��ϭ�yv��O���*�T-�7%(��jo���OH�B�F1��w&�޷/�;���9��:f5��ieUf��e�d���]`!F�0�j!�m�+�Ѿ�)�蹣���I�8�{Ms.j��N����v@:ΚGh��|﫷)�e\s�G �}cPh��[�A�r�$JC���h���ݡGy۶����5)1gv��M-���DW
W[|���j�ݴ��|��U�J�Bʓ�y��\��F�T��f,���h�z��`iwt7��n�L/�aTa��j���S��ݳ��v��m���Prn��,r�����ގ��C�3�)F+�k�^02�Z�yzɚ�o��u8�}-�G+���sy�q	����5
n:����iU]t�j��b�Y��v�Z�ת��o���>R���Drf�����,��h���ݒ��J���5��{&`�W�aK������|�ؤ#���H��m�ںƠT���E�Ӻ�)�D\=]9}�^��+Ǜ�k� F�^�\w;3�s5��յ^p>�����Z�V��츴.;GϨ	��Z���/�I�t�=�Ô��V�$�q�yg[y�Q��5�v��̚���� �諊{iX�w9��v1�=q{j:��狽&��j��i��ԕ��`��7��^��^?]�^�n4s�t�.V�I�ѱ�2�eX��b���>�m�aP%o����,��	Z�];و{���bŝvԙ2�5�*��`wG�0j���Í�ׇ���'��nu�gm�cL�yC�?��[���u'E�S[��=���c������~y���:Z�n�zVO�8�,�Qʣz^��͋Mܦ�����`]wC���D�]����r���&��V�_Y�a��R�4���Lv.�2�봹�Z�o�ޅ]y�z_�ĪSi��މ|���}�n��z�W�.5N7��uc�j�W������mNĥw��jd�E�ë�Xi6�'k��u,[Wu���n����+�U{6TQ	���=g=W�|��Q�hq�e�.�հS���k����S��mE���xۓZ�=Y,E�Q���.˸��+u���ގ��������[���W�c�D6�U5eDO	Z�>�4+��{No���f�Q�^��M�m��Cb�`l-�=j-�]��������˔v/-�0zs�bOt�Pm&���V���}�ieE�+zp��0�>�oM*�J#�S�gi�CKH�-t�N�7����y.n���1'�#�岶nd�w���7Φ�}Er	�bwy��iw�s��m)�i\�(����U���9�{G��֤��RW��������9��}ϳ��̞��w�1�7)�w�8D�l��	|�U�jW�l�5!m�Kq�7v��c�T�Iq_=�	�4,��6�l��NK��'�k��Nк���-+� ��w�58��*�u���®�&j���X�(Kx�r;(㺋�����b�uj���Q?u�z��U&&fÉO��z��.�4��CX7o�"�%]�T-ڋX�-��Xѯ8��D*z�s�M�"^��(���6����^Į��>3{H]���ܵSؚ�����؟a�xwj5��S�_S{Q
o�n؁O���З��ٜmOk����J�f-��l���
��>=�w��=�(N]�d���Q*�$�х�<Ύ�pbq��氮�{8{w��-���Ol��#�u��MWf7��ۈ7Pʅ�&�­5����&���3��b��t&�jI�wi��j���[:#�`�x��i��0��o�&o�m�7Z�d�3lKU�3Z%-B�2��` ��ݝ\f���%� 7���\�	=�P�F����!V{�r]�� �=�WB\:����[ܣ�"O�2�H�n�h���(��5�vq/�}G��w�'�\�z-�8V�X��G,#��밹��>��Я3�C��Č=���o=^��k��)ݙW=*ن�G,<.%k�����N���%>ro5�Cs�����a�N�;�
�B��0�b�u�j�hR$�7�s���S��WT��{�O����]�}*��s-lfE�Y���ek���qu�;�W�hk��qc�՝�V.f���>�S6и����t���J�]f��H��Q�Exe.V3W{~p��|ꧧ��ٺ����SX����Y��;<�D����}�����K�Eb�߬b�>��i���j����a��qܜoV����G��ד��1ι8�X�&�&AvҪkj[W�|�>ڱ��ߚ����	%C�qË�m�}Y������ύ�R��k]Y�<��W�$���y+�}�\�����^��0�X�U_�|q]������i��*����Ì5/����	��Uq�K�3v�{X����p��,��+tA0���A�uF�]��u)9uX�
c<̆e⭼ǝ�sK=a�5IGj���nݡ�o7M�K�֊&�U�V��R37���舋ڬ3�O���wN��ڎ]��������ѯ���qjy��ڎ]�c[N_T�T��1|�'��<���?V�Qg�Y|�T��)���}�M��f�E�q|\Wr��W�ͥ����P��m���蘧�_�+�O�m1�<�����'�����ҁo����Z��B�OK�TIق�WsS)t���
YG�Έ���z���2&��7�oFL'M��+%áe}'���pO�<�u#�\>�s�~p���x�=9��(z1ܩ�-�+50#R,�2Q> �τo�/'`�Y���č_��Q�+[��GZy
�a�R�0���"6vYK��U�E��j�>�\���YU�7�\��-����&Q���@�Yy�-F<��Ū>�X=]�O��[�\��_�GmT�c^w����ʓv�C�8ŕ���57���x�&�Fkἴ�����Xϗ{�|��H���P�nwʭс^��b�����u�: �0�˻'[Ǡ�V������@s'��3|zs�yX��I�U���� Rݿm��b��z��N�X6�2��!��F�����$��t�A�Mɫ�|�Ҝ�h�iv*t���B�t�k~ ��0@v��Et�YՈ�����Q�:� Y|kn``m�2� �[��Z�E}`o.(%��\�n��@�t����{��MBX��Y!	�����
*�KPf%�}��0+�<G��6�qU˚.�f��Q�����*��H�bwvx!q�Ŵ���i���c~v�l�ظt�{Pwώ^�Mrө7	 �Oq%���e,�XT�)�\�z�����OH�n�u��E5T���e53N�ҐK#��[�!>������o/7֡��;nh�v���z�m�N����N�{�h�P �,��+�i��jPf�,�u�����L�Kn�j���w)u�V뚹B}�[�Z��g�ƾp=i*��-w�rC�j3/�W�1F����P�[}[�y\�iS.��	�GV�Q���p���҆&mi���×�$9�F���`vU�ml��}{[H� �����C�#�O���)ni�t9��N��r]eb���Ǵy�oY�u��{�R��R�[�#�]��V�ae�9M,����e'�9���OLg��ݗ���m�j����\����=J����l��'���,����M�^�Y^�m�(,l�;r5Wk7{��{ .Q��QS�χl����+n�H ��B��z6���Zڟf�[�9���Vm.�|�ݧ͙�%��hN�˨��!�ڻ�D�v�U����t���G���ۇI����Wdqf.vݩE1b�8s����(Ie�jfە�>�n@,�}�v��v�6B�օ��âv]�*�ή�|�ܠf���f^�w�[��Ě�θڗ�'2ˏ��Pr��-�-�s����Ħ(�U`B��p#[^�vL�^͑�l@ת�=��R���
��Wt���TD���:Imڥ������.u��Y��/��wo�2���U���� �.��n�闽*�����|��_*
�*��/:�y��54���-��l�YJ��ð�ͬ��bpQ���-v|6)J�e%K
�;��v���\�<j%�3��XJb���6��qM6��a����/�K��l��k��w<O#U���L�v�|��Jă"�zed���h&Wgs(��_+Q�l#>���u3��ʔ���v띜�ޱt��s*��GP���Ԧ�R��TJ�Q�i��Y�mҒu��k8�����vʾ��v&��R�h�b�����A� ��Tl��w)M'YId��H��u{^6x���sp(���51Ԕ�;X��0�
׮�By�N�tb���Q��* ����������η��d��F���
��ꓮ�t����W3��fM6_R���j�X
㠈���R�Jt����#��>���	�C#�8"�i-�Z(��Ԩ�VU�L�Uq,c*�jS-�Ub*�F ��b�R(�,DDE�b�F�E�ʠ�����2�bX�Ve+��(Ȣ��A��YZ��Db"�Q�"�*�((�D��V"�Z�kDe�eJ�S(1�¥UX�"�Eks(d�,bcR0D���"!���,V�"�ZQ���A�b���j�"�*�1q���*��Ҳ�����Z�"�*(%eU��X�X(�*\�X)UQQ�DEX����`�5���X8��l�X�m-�Z9��*V(���b�Fe��"�YH�-�F�\�dm
��nR�e�[&P�f\V-cjL�̡�[�bť�q�V�QEVE`��"媌F6�T�3E�L�a2�{��3����˻Y�81;��l.:�A�C��ZEÝX��|���pJ��*�׈��08m�Z���<1�	�ruӗ�W�WՠK���S|���9�/���ͺG���u�{=�'E.ߊ�mMU垺yt�K�RY�H.#r9O<]%��9�'�j9���3�2?��ؾn��4�B�K�j�.�Dߏ�j~c~}B�ړ��kӄߔ�`�yfSX7P��)��oB�N�e3���:��UF8�5��(�mM�k��qn'�8t��u�{3;9�g\~�+��zԜUq�(��F��<Ov�̦et�C=v��nl��^����Gsk�_q�J��~�k����p���Vڨ���'3	e�ө�o�[�U����1*��p�9G}9�¹��n�ȏ ��t����.�Z[�p�97��Wʯ���=ME��d�N���.T�^.��kM�.��⯺ewdr��x�k�)����������X��ʻ���5��s�ss��\��t��)�\Cqڞ�u*g�IV@�=n�˂��]��s��ϻ7�~�u&I2���EF�V�ǌ&�T�t��o�hD�z�%�>@n"�֠3�+��5�t�Kkq�Or��Yw�R��o����u%��5n��u�K�������.b/{�=م��m]ML�\W���!�ָ�9�
�0B﷯��?������Щkp��SWA_D}3 .�&��n��,ĴW�ʞ"V����ˀ�w�5d�M�u�M�|��6�J5�<2�\���f�U�bWd�F'����XJ�#�y��wn7:˾n�Gϡ�R�C�!6G �_�.J����Ѣ��kO��@J��VOuK����>�3n��%�:���N���M
H�#�;6��#�}|��mDk�q<��۵�R��4:�N�np�UNmx�b����$����꥗�	V�/'*1=5��?u�w�\\>GLܫ�us��V��FIow8���ap�W1mo�ˋB�B��>ſ.����,��L�}��Ha��g*Ya�)�\Cx�����������������_H�lV)�}�On�J�m�9%��6��'�w�f��F��{�k<��ޣ�.��g���yX���M7R�#,
��f�4i�pJ�A����U�(�L����T2�P��6P��B~7]:�����V�k:���0���chǰo�Y@���H��C�Rӛ8�E<эq=1�
kh\T�R���on;��&T;������ʺ�w��+�RWҺ����oS{_)X��K`.�O$i�[�"%�ۣ{�|r�[����t�ǵ��>s�g��|���s���)N������}�+OFc��?Jq4�,+�5ꨍ�Igۏu��O�[�*:5�on_<Z���u�:�в�$씸W֚ˌ][�c�HQ`��3FE��W}vAT�|2b�V9X!/�Z���\.uoL
�oK���HqnS��g���z����O,�+�=q�^���s�ӱ6&&%���Nj3=�`9L-���쾧�wBy
���W.c�]�ab�5$	O&A�{.1e�ŔD�l�ķn��^�}N�P���.w��_,�����r��=C1[4��=�xq㝽[_oPU�*�i��S6�հ�b�{ջ��1�"튇�u���<t���fb1`3��w]�]%�����ˬ�7 �:���Ċ��!ɣ�L	CuI�ie��"b\� �t���g�ʱ+F�u���
ݨ�#4\3��NmBefC��hf�(��K�G^�43��˷a�s)r.�D��nGS�t͓z��D�#����v����oWa}�w���%?�U�Q��E:r�{9�Y��Yq�=�;��uy9���(����PK6����9O�����T\\�p/yZڧ궶�������X��g�<ko��*�1Iܥ�~�uvV���׺M�~0/U{��~����M�'��0�7�S�mťU�1V����.^Y;ޛS���#|�L�ȫ�����|^��.��ﱬ���h��}S��O�ˇ���=ڎx�Jou�Sx��̀�yS��)8]���pkZ�<�>}�TiO���(��ۻ$�ĔƫyR�*�w����-�oJ����N�K����%�k5W<�ʾY;U��	B�M�T��m�
�!�nM�����o��8^=�CN��L�:�α�t���a4��5e<gQNv>=NWܶ��Օ�܎3d��}3S97q�S���n����7��F;�9�*��W���f7H.'g!GeL��_Mt޾�^��/0���ƴt�yX�� ~��+MX�-���=����ӈ��:�w[���v�Ty6�r����"�W�~	wۘ��R���+o�S-s�8.L �=�`�H��`��*�Ã)s��ؑ����o:�/���n���R��@�:ar�ٖ���5sp�G8j�w o=�;2]7���w�Zb�-�
�W	[��<�
��{�;+�33�M�l���}%�ʻ�U��&eh������_��g˗�¹�����J�gn��h�g�\'i,�u'�5}+�ۘ�|=���k��+���~��a�Mi!/>Ȏ5��SB|�Ve>�������;C�ߨ.��a�o�em"2�C�bޘ��c᳽Z�3�'��ĸ׬�B׶n�ޡ��{."P���]ol�^��\�J'�+���>�P�V�'���p���Cj��,�עa�%@�C�>/�K�"���
��/oǦ��^ߩ��|�umT�燼�P��������4���=ҷ�Yv��&�wg�,uD���V1�b�U^Rl ��V �٤ͷ�շz���CX����Ya.�9��&�ֵVqTY|���p��8��)L��U�.$Em�p+&�t�"�+G_��l7v��Ǌ�Z{���χA%�Gz�ZC\�a��Lb��{�{�	�#f.7R����K���#[P�΍���Ϝj�7�6sơ�� ���sr���Sq�ѯ�_Ue
����z(S��F�ق�������%R�H���w��Y����bųz�»��kns�?w�.�z��i��������0�j�s�4����R�B�܆��E7�sx�i�+�hy��e���RZ�w;��4��j�k�p�h�=�70S�Qk�\b��a>��u\=W����/���nS�}]0�ԋ�0�|#VT���>����Nb�U}�Zܹ�f(�ު�����S�!��G)J1Q�5P#�W��V���.��Ĝ�^���Y�]RT�M��3ޓ�k�k�<2�\��]�U��Į��in��`��z:��V��E�J�����j�Pب�j��q2�n,����\u9���ޜ����<s��;��㏓pz�Т.=�l���<KbWV���f���\��ƞT^gU��Z��]�ĸ�v�9�X�K�
�a�d��&�+C�ve�'Gh��DDR�/�W%�I3	̱�hZJ��ygz$5t��'�$i*6ELTO:�J��8����nn��o.�y[ƍ*�)�4��2jx��|kt+ |JÖvL�W�"�*P)�}Q�U<r��ah�7���}@�̈́�zD3�%w�{.-��w����y�}B]7q�W8���b��o�x
��#[��?$6�K9�K~�_-��SO�oأF�ͣOe�+����.KUí̎�t����5okܭ��qË��+�q3�N������']�Gkɞ���*�y)��s���w�,%NV��������k#{��e�uԸ.qesгcSxkϽ���{U�b?w��u���xnb��Qz+{7e$��P{��<�"��z�W�Ҟ������4�y���P6T�Xz��Z�u���tWYP���i�W�Λ���}!��V��i�=H_M��C�k*���)_�U�ZE\�U��U���_t��Ox�"�j��7_!�<�uc���F�ʇ)T6�d��%�I�<���j{���Z]��4މn�S���G���y�_�F*��b~V�T3��r_е@�u���3w)�NPe:��7Q��1va�4	������Z�
ׄc۸#�T��jwW0�t^I� +X�,M.>7ϯ'L�8w'܈{C�����e)mQ�y�cwC&��wAwo�N�Һ�H�(w���Y���X�[���K�L���_W�7=*3a�jf������ʾ]΢�v����w�������"����d[�;�U����k&���s�ˤ�������jw�c~	_�pv���(��j?3�����E_o�_R���|��aδ����6_uD�oMQc��|H��D��YSܰv����m����fq9�B�����v9SK��[k��8j���_���ۃ�ڋ�u�ג��߬aj�+��8LT�<S�kV��ᡝ���_7�+\�G^A�u�O)�H����۶�惘���\b�(}���<�-{��~0/W�[w��SD'�J��+�U��{e��>x�z����k�!�犷ޓ�^�.K �x��n(QROG����_�d��8��r�++�M���%�t����,���t'Q����$�e�0��Ī�7ï�1ZՎ[e��*�Ҟ@��br0E���,�yM�=8��n�4����@�.�}��ػ��z�� ���+��L�4F4ۙC"�u����3�(���^e-Ì�&��m�{�=΄�Y�Ѣ�LZ�Zⷍ���u���̺w�xhL%�V�Y};,v0��.X�\������ĊK��������o1e�	�t������on�������7B����#�7�QSN�b۸H���
j\�����Mm|zӾ8��B����~�s��N*�.x���Z��ѩ�q.�s�ݮ�:�����Z���U�J:�}��8o	���.��e�Z���b��u4��
�#�MCr�w�;Ɗ�u��d*���l�9}Ѻ�jʞ������ˀ���[�;���+��QY�,�v�Kf�m���m�a��\%n^@O2�+��e�CM\�C�̐Տc�x�:�O5�����ޔ+۾��+�������.^Uڽ��K��+�[��-3y�ut-jn���T���j�]�����C�&��ᇣ�{�\��w7T��m�F�p:��8��om�u_hׁ�����q�(��JMݭǯA��z��]%�C�;I����p6�Rྙlk��a(�nb�o�^UewKT�]6$��k��.:t���Æ�'i�̌v+|ݧ�n�:�izt��p�xO.�j����n�6�y�}.�0�i�)-c}ݕ�:�"�^����ö��[Y��0����ǘ�8e�q��w���U�Ι	���;���y��X�w�}IDz��~���^�y��1Y��N=�A��z�ACX��w��Χ��b�u�'qD�Zǲ��˞
&k�����}Q�5r}��5^Į�m����kR�����ǆ��{��u`p���ϛs��a*�+^���=�9�ݠ�8zu�r ���Jyq	��-�U�J��Ī�M�77Zߏ�3BX�;g��+�K�m'Ǵ'v��(��ڋY��hYQ	�wb�0�h�Gs���\�m��ʃ8�5=�b�*⻭h{��d�M�`�<��N^�5��󻣶��*�I���\��uwru|�jCE�#*���&�<�,��-ź�jeR�%0#����	���w��n�{�dL�o>���N�rʶ�M�\��Ҕb���G,��xZ����T�U�`}ٰU��wOoԫW�;i��{D�d�z���;1�Z�#�v�,���9�EGҔ�u0JVN��:���+���e"��iu�_Q{�3�l.n�ۗtK2�owt��p�GQ��P	,?[<���p%�9ϭ"�f�V��e�"��F�������uӊ��ל�0�#���wŵ�󄮩NEwjn�h�U��Z�.�ۻ��Μ�Q*��|�ٯ�6�s�k��ea�7W%,�%p�{��K�[��`a�k3,*�4^v���M��ؘ&�F�0Ck�&�Ω�
��ٴ�u�W�'Uǩ��N�µ�*�VSk4��Ѭ���X����J¼�t�s��x��uo2=ڠZ���j��v)m+6#�RX�r�Β�Ԃ_	�]]�w��'���v�N����zi%��k�׉��G;B�z/b�5њA4��#��7֬�n�V��5���Bc)"F�:�:o.y�>��J�=|m���8��xF��WN	�$�ih��Q�@w��FoR�-�jF,2�!k]p���M�rĕ�d�b��Q)'��|���VC3���q�U��Lu�Q������f[��R�����UXksFԽov �vl���Դd�aC%;�z�_wŌ�+�OBxi��X�qA���j�:�P*��BfX��p��J���0���FsMe��C���3�����2m��sy���Ҿ�tk�a���n�F�ڪϵ.��������]�1Zz0iX�3:�V��V��k�	��n�����QH���z(�X�-|F�dt�Z `z;U\N7���r�!�깎�|5ʜDΝ�Y��yz��w��<�]3}+�XL1XU��۶+�� ;n+f�.����Y2�/Vu]X<��;�V�3:��l�[�E��'��ۢ�E�K@�A+����z3SШ{n,���։��"��ܻƥ��Uf��۔±�خg5x9���m��z��mmaj��������6����d��r�QҼ�jk6n�r���1�Q�ނ�dM�Q=����
Wh@\��r��t�{q��{۩nr�^���";kRɮ� -ފ��yM="؃���~�ٛWD��i>A:'c-�E����yw�)Ab!�qQ���"���Q�`��x��4�;�Đ��ږ�����
J�׷��g$�Pg3���'���l�௎�y��Ya���J�@�|�)n��]��|�}gk�M3�f��	�Ve����O���Eq��]�0��e_.�Y@�q�6�4U�� ]\Q�
�)P���(b����w��B�U|�c]>��A��kR���1tUvcms���.9/�ϖ�Y��M�Oo�}���R�u�.�A�wNO�In�Xg]u�%��І
G�OF>�0	x9c��#�i�
�N�X�"6jIU����˸˰R��x��!�7t�h�x�Ƈ<[��{������x>�LT^���\KYQ�l�AR��3(��A���\n5l�AE��V�(("#����U�(�԰��C-��UQ�-**"#[-(*ň���Ķ�nZ�2ظ�P����"b,
Z�T��%J���dQ[h11������R��� Z�6�j�"(EQ(e*���j#�e�Ԩ`�UPUXcb��T��
�kiR"�c�!�ĕ��AX�J�*�c�b1"�8ш�ŭQ\j�W-��X1�
�dDdm�EIiH,��IQ���V��(��E��"��H�&YZ���E-�TDTAFDeJ�Q`��Z�b"�LJ��%aZȶ�Em���[
�ҫJ�����0UU�1��B�6�b)PU���Qb�AjETkb(��D�AT��8���T��`�D��N�޻}������9�i��m�ѽ�3հ�=��]����Ub��!�t;Gq�H�\��{�K�B�@ǘ�זo���W�T�QW��9yb�3��_�̳�ڞ���W+�Cy]�g�X9�zB5�^�|r����Nˍ�ݰ��K����j�P��n'歞��y�v�)�4u`ܓ9�$���׮֜X�~ד�U.���P�N�G��Brg�������@�jWm�YQy���ڴ��U<]%�=��W�S=�s����W.󝜽H!�N]ý���O�o�b��ci�
�}�S"�n]8��眱l4���{��y���^ˋ~���6��mR�^�bh��xe��B��%)ۅ�����h&��P��X7Y}�J���S�������ڃӶ��E�g��u�W.�k^�wٿk�ԳW����-���9�r�s��ʪ�qg6�s�+j4���{�"���p�y	5��:��ev���j��e�凘A�J"v��Ɵ�;��y�I��7���s�W�L�Y�eV�s�d���RYOjl�du֫� ���,�w�f���v��ʃG��V^e�G@��MG�I�#ݣf�KRs���B��:�'��j.t*�uݹwGE�\�X��+��(�T&�Y�NV�����ǆ��W�Tܱ��ES��u�Ī�OB�Qq)D��ΏϥS�����x��05i����8�[G����X��Gc�s.���B�T�	UG��|�3�$�_�>5�y0nW}���+�<9�wKJ~엓;FXv���,�r�wO՚B����!����ZV�3TK��wGR�g6�+�bUv�9!�Vwe��̿�s˹�}N�;�֞B���W.c0T�U��R��+}^M�f�7P�z�F�~]��+���]����mp�dbu"k"��݊�ׄ09�[x�<3��ڲ{�����_wd�3XZ��ڄu[\�d�cs7֎CTʝ�}��T^b��q`9�Ȼ��ٹ�R!i�4c�t��8w!�P:�M3sY�g<��>{pw�W��������ȩ�[:(ޭ���H/�9O5�(|��<�P���r������ܺ�x��Z�r��JVw�"�o�a�97��m�X>��N�u�n�%�"ľSV�/Ԑ���kY�Y�p���¸:�m�^Y=��d�u����kƄ.��,.�zQ�75f��v%H+��fN(|�������X��{��f��'̜�4�n�,�'C�T7��eUU!��zk,�����m/R�����S�GD��mڜ�Y�M疌r��fs(o;����j��Q�����*�/7l<���nT�l��{=<;�{��x�$����_3�J��,�7���>���s����os�Ve�e��I}\�,�׸�o5,�*aJC��5�W�yTY|�T�+eY�i��p� ��z�.�O���vS}E_e��B��%T)P�����D�>]s;_��DU�8�ɘ_���?k���q��oB��c��|]��YQ'c�j�ul�߳g���3u�.�����i(���ZrӁ��^JU��) �]j$�y��ˤ�X;>
q7��tĻ��{�����wJhnd���6V*Ƶ�T�!��YQ=2���2�'=��
��֎	-|5q�U<�X���?��r�|a��p2�2�y��#y�i��y�v>ۉ�c����ʁ�P	�Rwu�,U�擔�*i��,5�m{6ȹֻ.�/rm/�{M[\�V+:H�J�_e+'&���t��}�.��I�B�
X�co�	��w����S���1�5iڴ31z#��wi��Y��x��VB��A�Z�* �.�*��s]�c=�>i���i��n�.~h��Ij��BYM8{�nB7c�=r_f�����*��h�$Aʷ�#8��x��.1)Iu	�Q�q�8D����/�ż���J���g��a��+���u��˻�SSk��o��.��U7c�=q_�'o���"�����m.���;�'��W��i��v�uz�٫�"�^?��֕v/н�v���8��s��}X����3wT'5N=�Θ�F�C���b��zmN�W�{�r��	��9a��B�����W���Q9���_.�R���w�3^����_q��+�
�������Ү�����wvq祼���T-�����E�=Q�iTx*��ay���/jp�r��n�f����|y�x���g�����8�
����>\HѸ��9�F����Q�>���[.2L.�᭺��$��&��Ciea�Q�G�)t�kݗ��+Ք��Tw��5t�V�|6�f�:�(BE���;�M��c������{;�lY��>;�<�32�N������.�wv�D܋SS�興E����ǜ2�ǣt�\��joLu���:Wu���<g��#.f{����˃�u\�?3��ě��S�R镭������2����w������-�ҚN\��0���!>����'�ޛ�e����sd�	2s�i%��8Ja���xĦP��𿳟��eߘͭ���7�a>��3��|_S��7I��\���=��r{y����o�NjԼ���Q窗v�s�EW'N����1��0��<9��Q�j��r�Z�}ϳ-�����-韱��^wIX�K��>�S6�@q�{�X��oz8���U�CX��+���ʼ�W�k�Z���*�_.��|R*a��F�~��A�􇹀����}^nk�\V�W�˴�[K�ƾ�����n�|nSj��>�9��#��0�x2��7)���"�:��8c�*��a�Y_uT�cG�y�eG@���NS�9F)M@���!G��X��.�F�pN���u�����g:b��\���u������ݯ�&�j}�M9�	����ت�Kxa��-��k.p�ǳ}�s8�F���Mÿ���TE^��g�����9K R�yyY��>~0:�V���T9ƏV��6�R��lە�d�'�g��'���Իj���k��w������~BJ�J����dV@�w<-�{mG�Dr�#�3|ms#ӏ�V�jo9�{���T�eKpki��osF��byH��֪�*�+�ƫZ�󞑿r!e�4�/E��Ӣ���5�_;n%"�f����~��\FJ�ר�ٲ�+���*�w�oI4ΝQ��t����m	Z��*-��$��:Ie>���4����P�v.|��jC�wm/Sp�/�Ϗ�y�Y��B����A81�Ð(���l��1��.�Ġ�}m�p�b��#8�d5�^���qeהD[��3��4���	�<%�y�}�p�����ꚅ�uD'��a`T�����r���صeT����<���ɬOvgs.�>�C�i_}�xVa�%�*�1V��(�]qsî��.���q�:r�VVG��q3��fgfx�|q׶���ά��!i�φV#  /��J����`���
��{a����
�U���2��Zt1׵��������ƝIu8lE�I�/!�$V�1޶�=�#h�\��5�ͅw�g��V�w'K\�^��D��09vi��x�<���YJB8��n��(s���6���{o�]�M
���2^��uw��X���o265��M>�q�w��}���Bs��G?�+���w�W�ȉ"����}ZuL�s��}��'����.U�2,���/�f��BȬ�[U�A7��z�%��cսxo#c�P!ޭ�<�F��^>���V�����aI�=�Y�/L�qË�|�uuO1��ꉥmM��h�PU�bM呍�퇝G���ｑ\Q��D/mW*Ҳ�7����������o{nߪ������D|�H6[]��v���OEa�A&���6��}�$kR}�I��*�dB��������;"\��!Z�o'4����y��C{JwmF��q��o8�n��m�-
��k��I��m2�0��؄�������/[��Kۜ�E���ޜFE��G �#R�����Ωt���:���Ka\�B�ѩ�+}}/�j��Zx��``�5��u|!�a��W�c�t�T�՜4T�C������fr�S(���S3��Rm�b駎���8]��;�r�@�K0�P˰�eJ�K��T$����]����o��zOx���cN�=-��wճr�5B5eOL�Z����	�n���ri5��N.�7�8�3��9���S��ÿ�^T"�Ls�C�|ҵ#W�H��y+)z� &�~���7Ԥ��i�SqԞD����A�]��T[k�@�.�^/�7RK�]��#�F9��7�ݩ�u����ɞ�/�����n p�^v�'F��?h'��2�+K���UB�-56#��G�|XNqX�n.��P�2*�K�Q+���;�ux���3������qp�l���������[vK�z�l��S�r;*;����bڥ�c~}B�ޭ����'��Ϯ�kj��t����&��s%�)��E�|��i���u/?Qu���B61��3����S�YdU��.���r�&�o�-��y1�6�􁖮�\��#ꎸ�{C���ٴ�1�o��3�r��;Ev�T�p���́;�ER�[*�m���e�N�ȻW��gkj�T��\�/�t�`��79�kխ(�ot��`>���m�bWr!r���f�=�]<y��l�p�"��ܨ昧���y�����w6�+��Mǆ���(`�f�\m����r��*��i��Ӵ����Ź�__�ģO,@*�;�y���T��nꉊ|�,�w������>�MmD�|�^s0�ov�����s�b�$��S*��pbR����1t��ߠ���͙��XQ��?WZ�]�Ǣ]8�l�cUʇ�&��
��.1t�f��ioid�ڽ\�U��$���#��[�R�R�a��rʓ	�ς�xp�M��nz^��]���W���T��RB29��F��ᓰBO`����Y�1>��'��G�>�=<{=�O��2�Bz9T�����ݪ�w[��/	�ob�sQc�羥�l���4v�;��y�n3q@Ki�ѡ�()!.�
�k�����f��
��L��!J�H��\}��l��÷ �����O^2�*�+jv�te��.��O�u��4�L�����S��N��^Y4�7謃�a�zt�m!v�mu�5i��lh��;�^]��l7����������k�*�*㺨��%�ocu>\�hw�̑��ZR��b�5z���*����Zq<_Ɯg�M؄���|C���Z��E��h>�����o��K��=|�.�O���:M���B� t���妡�ӵN4,�|���\[T��v��Wy��hgT�����}6��7��yp���_b{��඙:��\v�)�p�b���-J	o��D��g��Y�+}��F��+l�,�|�	Y^W"�g�g�9<mu���K��Q;�^<O����ק�hdL���:�f��޾�Z-<���%���:�����f�o-�}�ޕD��8�b��mj�|�f���]Q�J��7����j�,򯬮w��}�<�H��j����4���rb~�>~<��w�j��[��W[YF�u*~��=���AbXR��!���9u=3ON�\b���gDm�\C���O�f�χu*���SVrH)H��ۮ�<��w-N��q�Y �Ķ�Uփjr(��`׫/(�|�]i��|���7;/�ԭ��d�7��
�e�7�xհk�m�<ƥ,��ҟj�t���ڷ��4�7[Ǩ�nmG�NOcTj�t�>%�s\/$�Y�G���Ϊ�!��t�,��kwW6���x���-��}��w�we�yEg�q�r_�Aa�l�s-�V8���z�I���e��%[O�D�/� jR��v�۹Eu�C:������z���ф����;��֒��ʆ�Zcx�)�5gsؔf���U`t��5�S�գ��4���(���C�4r�:N���ƥxh}l�w���Ѡ���G���b���|8��<賨f��|��vZU��|iΡ�n`/����qn��\M�[��sw�S{p5�5��B�U���&�\g儛���x	�Vo�EҬ4��`
����a�Xsa���hoRV�3��Rf������g�����:�b�J��w"���T�٦gM�.�q����ʖ����B�L[SH�7d��)�z6W.V��Z�6��5%��R��/zV������uut']���w��;�ʷQ�tj��&�Tڎ�+���<��.���y��U��p�Ĳ�V*	t���(2u��*I��v���x��%��'л<���GAǩ�!������S)�yW�s�5��izT�Mfp3-��܇J����7�u�[q�-����h�Wl)6ٴ��Y���
B�mwp��*Wm�$�C�|���bNZ{�f��J�E�B%�N}2q���*���@��U�XA����;)d��vj�Q�V)Aݗ�c,��j+��G,���=Md|.�NG2�c�y���; ˒��A3�6�����܆Rۢ���z�R�դr^�륰�v-h�R����:�|��/wke���i�n�m�N��ׁ����]���9��T'8���% .9n�Ԇ�a}8�{��uLP�(j8Ui[x��K4����Kj�����x@��w�]M�F���>���A�V_jH�D��g'WeYu��;_,�ھӇ�	�N����gH�ʢgp���yJV����s+ -�\�!�K r�Wu�yZS�&�^��#��^����o E��=��:�q� b�1z{S����b��j͛Sq[}z:'9���l=�\�	��c�p7�b7�:�������!Š|�e�2���M\^qT���8΅�{���N[޻�O�}�&�s̋�d�i6�L�����/giZ���������]w��#��t
�[�^+�k��f�-���hBeF�F\o��\�ܡ��"�q�<%hc|����cJ��t��%nWb��lw��6�P�e�o����p�d��r�jO�ü8�`[��} �Hl����;��O��o�
-K�Lln���z����R���Fk�[YWB����;:� t���[G�'2���d�����l����g�b�M���d6��vW|C�N��UvRV��E�Y�;����]y}٠t_*�B��UF

��U��VDX�U��̅e`)ȑc*�1�5�Ec�%kQ`"�2�*Ub�e���*UH(��1b��F�Pr���b
,cF(��@PU#"1X#�2�X�X������+%B�,Qb�H(�#�b�Ԃ�IQAb�PUFE��dQV(�V�����Sʢ�5���PDV
#V�AQ���`�T
)A�Ae�"(��"�" ���AH��*
J��VЬU�H�Db�V$R*�,+*E���@X���$��((J�"�(
��[b1���Q ��E�b�`���b��B��
��� �TKhň�E�b�*�ȡT �@WJqK\�����]�
��Ku����9XGy��ǖ>�M�9cy�u�氢[j�����C�A���1��7d��Q&r��R�d~�����ԭ��wIXs���}��5���5ue�:Nsi���O�]���+uQZ����щ�W*{�&����0��Z��������c��P1�����2����n���w�)�MB<�ɝ�3`�^"��u�a�4b\��fS�����!W}��o�ͽʎtq�}�ªzڮڊ�nCy�+f>�*��*xs9��f쉦r��������\^q�����t�D�[*n*_h�yy��/Y[�e�G;�:�D)��33}���-���ل���_=�;I�;GT?�,�O����7��F�\�=�7#���2�79X�3�8ޖ�p��;Q�����2���jDWZ�G��|_���Y�P�t����Z�K�u*��s���3�O氓,�ż���5ۺ��ѐ���철���������m1��D�Zǳ���;e��
�.m���-D��b�<����;4��:�<v3w�RF���Yo����Ƨqu��7;��צg=��E��q\;)��*�FL¸�.�.A
��8D�b���h����ܺ���g��V��ە���ꅙ�B♣R��hs�ON�xJ��Y��
6�Vt�Ri�O��F�:�%p�,3{j���u����35n�[�̮7;���kZ:�?�7۟V)�|�^녱*��=p�Z��D�]uΥʉ FCϼ��q���)��i�dS}E_e^�]����m���g�6*������Ue���Ux3�Z8:9ǫ��{��N���9E�Y�;5��׈�U���M�r[ŀ��U#+��@�r�]dm0�ӣþ^�2;�+�g������ǅ =�N��ݰ{�v�<�|�'ўfG��*۪��J�, 4}y0��{|Kґ��>��XL\��2w�N^v�������w��!�5��2<� �ߩM
����	h���~4��Wj��=G@�梕���^A�W���Q�ۑV꜑k�|X�0|2��"b�������fU �\?b��w��Ĕ�{�uTW�-�I���l���a�P��׆�U�d~���O���FsY{��Y�g��G�����J�G��MLy��Χ zᜠ*!{+�U��#�+o�R���9���j杺����+R��"���ɩG��/io��uk=�۴lt��6�)T����[՛}:�%[��(� #�����y�������Ӝ���o8������ӣק.q<�OQ��1�'N��Y;{�+�n�i�W��I����3[Lz���žW>�ϟ�@��2ϯ��۠D�q֣8A��P03��oٽ��G��I\w�OT>���L<����O;,���~�T���R�Ƿ=h>>�C�9o'`�E�𿼢O�uE���xs�0�f�i�/Ǧ��V[�+�KM��Z�X����7�_���~�%�ʑ��'G��e�83M��em¼�+����O�>F��x{�T��TB���Z�\��WX�V��o��	^�q7��|-��;�}���VU1�gK��Dz�`�9��l���^�~4�=�)sr��z�{)�����{��^����|�i�[6�ւ�Wl�F}0��{*��$V��iC�3�n2e"�B�3�|1�ב�W��K�q��u�P���R��o@��~���V�[>��q���O2E�L�d����1qʟ���ϸ���nvXb�XO;v2*������Ys1�]K��Ġ�MG@����J�u���mC�]$r&��s�ͣ�٨U�G�!���������VԲ�l����,t��FFT�h�%��ͨh���Q�α�Rj=#�th�8��R���}��]�`0{��+I�4��w��9r��RW4�D%>�on�8&(�r������'A}�S��2��3�_�5̑,Y|v���V�}�u��(
����^�f�㻭��%�d������ύ�%^��T�L�6�����B�JV�Ȅ�A��ӣ�N�k�W���2f���T������s��	����W<���O��-����ľ�x�A���?I���n\��uNH�|͘(=�/Wn�f=��0���7>�}�)��/N���և�"}J�1�}��3�S�5��y5� Uw� 3��>ݼ�Jz��DM�=��LM%[F��>�%���VK�|x�P�J�`>>nߌ\�G�l����x�+��	>z�x����M�=��0���t��/O���4RVi�������?gUv{��՝��F4���t�G��	G7�^�͏i��ڇq�^�|_5��?���ɫSS��R���&vn�.][k�<�T�/g��o�Z=���ٸ�Q��QM��q���v�E�{٫�"�G�Oqr�p�3���k#͙�=�g�{2�}���t�#�{O�0�m�b�s���U���v�����d�Zn7�5M�`mF�{�k���w���7�G\{�����]��#sᑞ+���Yx�z�o��EW�:|7&u�H�:�{n;m�)b�i�߫�[����7^�n^�[q�}hi����v�7�Be�w[�[L�eNP�K;�L�B��'˯�9�٪\޾t����M�h6�B���
}��wX��
췹X���rf�V��m�ͫ���т`���0�6^��5^w��Wl�0"�8�2�ue��Y����h�#��wIS1�6�XY3��L�'��!����IߙFsݳ�!�\b��Uϳ�g���xg���R*M�禣 ������g	ax비|��X	���vҗ��9Ke*�xpQ/��Ig{ޠ)�,�"��n�T\�9q���>�3L�2j��=7Z���G�+���i�G��q��y�o�E*�e�f�Ҩ�*�dy����� �Q/��/��'���#g�T_V�q	��1��U��G�N�e:����1-����)֋�V_f��]#��:���^��௧���kō�Ӕ�� �Q⑭�����g�/�������{T����#p`�����LM>�iωh���	c�
{����r��*G�ʎ��Tv{=z��k����nD�����Z�^G�����Ɨ�ݑaᨄ�kÔ;>@s[�p�����g,���ޟ+�>� ;�:c�원�{�f�Fm��[&��>�J����ԣ��juf<���f�ɺ�=�<�|���wμK̹�ô��/�%���׾���E�L^�FLe��o��������x�`�cR����C�Pp�7om@�a��:\�r�ni�u��OgQ�٥�����f^�F1��q�w��s��g)�X2Jji	�(�T��7�M>7%��D�o��}�r�Mƅ�vE��PiͮJ�*�V���>�a����»�v�T�b�ފ�6��|=�=]�#��^��S�Ǟb�F��5�����c�c}���������ge��}����W{ dyS����Չ�{l�r��0*����}�%Ett-�8��Y�?_Ry�?��T�]�FS b�W��N�<�4�ݜ�>��[��HO��~�i��ueT<5��==G���:�xm����D�x���je׻�����Mz��R;�Ɛ��E�ϣ�Z4���n+�w�;�>��t&����=�(��}����)���Ln�iV�G{M �H�9��U`ިw�r�m�^�5OR��yݬߥ��}�>���4�^ӑ�K�H��|�ļW�Ϭ��}DS7� �%��۽̍���9����@�s���\P��A����tf��w�'J�����=E���c��.���������g�H�����@ȋR�]f�
�=|<3�t��i�}Dm1��IʇK�C����JՊ�Ѷ}��j=i�܁�lUHB�z��Z>͘i}u�X���H���~�3�q�:.\�0UN\߄�$�א�"`֚�FxK��LM��S���LY-���区4-�c*]��<4#}'/����;%���=��KF>���p����m5..�}��+�]A<�e��|�}Z�h�H��y:�l��y\����Ot�iOi�cY˖z��.�4T<�t.=��y�G�� '�qJh��;�-�����V[�s��M�]Y�;Ѵ�Q�)�S�`��nE}꜐�'Ņ��I�a�g`-wx`���{�����>��3{2˂���NC�����C̯Q*�h�c07�|�Of�8��ҫ�fn��.��#���{c+Ð�Ϻ���OM�,y��/�+�]xK ����T��'�!��9麅�;�����k�s��m1ꄪ�5G��A��zho�\��]�YI���j�= �C�'�}%��f=�9�������3[L1���Ӫ�~�V��I��7~ݥ��G��D�xLk�8Y%�ʅ���B�ͪ�q����P�Ay��Ů����Iv�u0=z���S��nG��py�:��Df����2��_ѓ�r�OFǄ_���4:���w��@�D졺��~��u�'�3��\vB��#�<�;M�N��*�̼s��N��`��=��(�jG�%z2g�b�T���8���?g������5�y�]�g�]e{:KdB��Fm~#�{��J*��:N��nm��_�r�廒��I���Edrb#��/��۞�jg3���Mʹ݈b+:�υ.����p�Y�"��E������;v�ϲv�Ǒ@IVu_��E�Y��+��pg4!�eټN��K֦�f�څ6�s����n��9�?ZY��/#�B��3��^G��x��ز=C�!�y��@^Ⱥ�v����/}��v�I�\�Upy2/ҙ��e���xX��X3�}�m���#"�-�\���%��tz��W�ۙ`>3"��*ԯ[0�W�f{=���w�M�
��b��+�#ﹱL%�޴8_���eV]2�	ω`{��dan�;�����{�$z��JoL�,p���ͨ�ϝ�sސ�3�{-�o��.������v�dn`{3�sδZq��ez��=�3e3Q}��__�s���%��T��mN�2�K�|�g�ѱf�����ꝭ���+����D׋����ӹQ�և��W�e/L�M�\��V^�ϰa���\��ZG��z��ؖ�d�G�������>�%��J�K�^7ʇ�$�z�*���ȿ]�����ˀ+���6��K����l��k��=E�a��V���+4�b��#����Ff_L��`;���K=8}�������ȇ;@Ty�(����vA��f�C�ͯq���&wÓ�"c]˧��گ�2Amg�v���ys�F�΂�>�	�CU݋���F������ms'_)]��A��]!Ո��'::J��:&����zMm�%���;��ɘ:�t�u2.ީ��2�2��Z����An�u�:�����A{��s�k��M��f���Rg�ٗ�;�w^##ҁ��2Ǻ�V/�IG/�D-7;,fzp39/�EMz��>��go�u�k�#�֜�#����~Y~��Cs]����۷q��҇�N�=BP��Ϩ��R���&<�KIP���)�=d�V��H�O,w,�o���~��{D�{U�1]�3�w����=�}Rp�b��:2g|n5��G����*��lE��s��=�����Mό�W=��/`�r�cۂ[*=S�JȊ���U,ldγ��'�C����`��7�.k"o_>\�z�xu�:{�p�d���ʕ&�R� ���ø�)���ax��u�G/h���uy�D�:���e2�/�������1N�g��z��p��"�4��m��h�f�Y���޼r�V�����qt��r<{�D{��>�W�Y2�cd���] ��smW�W��{�'Z��|��+�.�s��^F�s��I���s�Q_20Ϯ����t|�rW�P���i�ݏ�<��ْ/�YP\����U���D��3��E�{��xj�Ú��as@3[�nf��mvj��=��!V��6��P�]d�B���4u�.��?�����C�u��U�Q
bU'ݕ�o݆6��2�u���j�\�5��KV��O:����VW�A�C(�Ǚ����%�EÏVq��@�^�ƌWE���ݚ�h�ǫ�0=��_�1>f�fQ1����	h��	c����p���:��:`N)^�3q�HC�љwy�����	�;�������T[�ș�𘘊}[F���0�����o��i�Y��ޚ����Yk 
߶����@��^�c��<�+E<��o�xܛy~�[���wOq��X��������H�5U������}%��\ׇ#�Mφ�~�޷����2�V-���{}HMl��gCԳ25U>��r��7�U����ٸ��%������o��r����nSH��Lv����=���3���W���p=+^��Ы�Z]]O�g�[펭���|s�� i�Ϥ���G�'�XY�Zu�3���Y4���~0�Eǀ����d�W��9�ߴg�,�/�zkE�z+��z��՟UCÓ��;G��J�Z��v{`Uvw�G��j{�~�_2��޴r��^�27$���CJ���_b��q�;��EC|�{���[���j��}�<5yװ��t�����/k���(���.� VEU���z����Q�8�F�S0��A}�W�e�(n�ƵU��̇6�ͶsRwuN�&'sD:c9Z��}�� E-Qv^���=u�^�
�yX�ɶ�k�	t4��]�tb�	��7�c��;r!u}�'U�Oq5j��\��n��nE�5�[�9������ʾҪ+���%���ݵRv�ɚ�c'5�L7[�k7�f+�CK`��.Q�pT��]0]��v�ciH.�a[�3\��+/1�Š��C��(M�P90���{�R��,��n���0Ǳ���aMa7"�Ii��[u�4���ډ5���Q;��6C�7J��d[���j8��CJ�� �\��;ۧGEj��0)շ�"8&��͗���c���B
o���P��}�Z�/K�ͽ���U&,-��eJ�<R%Memn��rv�����!DrYG���,���ǈ�/��aofd9��o�vݦ�c�z���K�'_p�c�k-(�d�jȩ�Ȃq�ޥ0�G6�*
32�\`L�j�Xn}+A,;�c��ڹE��=���2�v7Kx�Ŷ����Y{� �uܛ|�i�b��U3N����pws��6��*[�}.��E�[&�U�����];o���埂��kH"�Y�)O�2Pgp�ښh
H����gn����P�>G]e�ǥ其�@�b�m����;��ml��lPg"j�ҰV�n�d+��F��o�D.��J�/	���4@�!"4�=�{�^�㮗ʛ��( �\j��]�k�;���yQ��Y����6
�W)<�u�ڀB���g�e8T<������\���>�K]�o�voSY�v��w(��|]����#r��c��u٭�U�V��i��ӥ캴�YË0Y��V��d.��B�}�z���$�� �轁f�+��q�G�J�M�����Tk���G��
骺5���� 쥯*Vѱ���H�^+�MR"!��6����k8=̓ܙ���Q}�@]��Ŵ���v��2�*-�N�������VVkw�g,)PT�yf*\����6r�ɷ�W*�<Ɛn-��-�h�H�iJ�x�m՛a�-_K�+@p�C�k�]�	��j�����j�ʾ��N�+ `,���������d�%`�o��`tnX`���1��,�ʙi���WV��P�<���i��Хn둏�PS2�<���m�7���/�n�t�ٵ���Q�y���8]���}Bp
��7�IP����B��g��(F�-dR�ǡ#���V��HWk,��ʥ����ϱ�6�^�=ο�^�G=Bi��!X�����G�=���9��ǚ.<N�HTz�t�ϯ#�N�Y�'�L��X2) æ;�i�<�,P�-sH��������^'S�)B�������P�<�b����CVv�&.^�R�����jl}\v�e6{�g7_qP_p������� �X(���AE#l�"�Ԣ�QADb�T`�X()*AE$X�X"�T���Eb"��l�"**,�Td��X�"ֈF"(��b�"��AHJ�X
�Ȥ���,QA�b��bT��DH�*�AUB[EUTH�E�ID���*T�*�d*U`)
�"�X,PQVb�(�AdPR�*((���1HDAH�UT��Q �
��Y"$���Q,ETE�����X��Z`��R�FwlY"��A`)j�h�V �X+�TKdXbI�����mEY�*ʃI�AQ��Y
�¥Tr����H�`�E��������g4E'7�U�Kz ��Q9b	��|�gvoG�-@�	u�k�P���Ƣ9�����z��(5}l�����5�g*��w���0i�z_�Gm��7�U�5%��mH�4�"�4V���r���W%����^�x�����^L���Ux;�2�Ѯ=;�?O��~��Olƈ�큡�R�Y��Q��,��r�7����H��e�Z���6�V�\<����O3��f{��~�+������~^���«}Y`Al�*wR���Xr	h�3�j縱���o�ӓL06���:}mr�^�G{i��F]:��ޯ��dy� '�(�����	h��y��}����0��ٔ�=�v�\D�Y��7<
����߷n@�,��/Q�b�0|2�J��m�]��$�~��Vk�b��^�9�R;� �����G��U��u�I�u��~��y�� ���>�=P�c��w��2wu��.~�����okà1z�����jb��C�}n��@u-���-Ú�˾��g%��rz���#�7Q�ͽ�'äֹ�f���%W%�j��.��ꍆػ��"�Hwq��֤�=���R@J�n���D�G��L;�������3[L<����]�'}q���Rs(�q�\ӫ2��2��]�ɵ3����T�U�󙨷k�Mr�i��q�A:����]50� �6���rB(��<s"��٨�&��+��k�7�:�����Z/�:Q2Π���ft�;��M�o��E
�)\�dV҅��\����=~�v��e!qމ#_�Gq�yT�M�Ou�Tǿ	��@T
�a{e�{�� �5�`\yN�.=��<o���ȸ~�Z/�h���Q��b�2��|u�7�_��^=��.f�}��x(�v��X�<v���"���z7�kO�h���W�����޿Dd��֔�W�<��Ve�ɝS��B���d{n?g�ȏ*~=�bβ�j��yu�{c��zV�a�Y^����Y~�qumh>ʬ�x�Y8�dϑy2��|;��^G��^���%�A��r�_�]�c��G��ao��<�q9X�O"_�3y2��GS���=O٢v�뮊��^��ҧ��6=8wϩ���Hx\)��D?Q�͹�쉨�M���^.��h�F�Z}1���6lɮ��OL�7�ǫ���O�vG��#C�z�ɖTa)K���2������W���ӿ��9�僗��7���z���>>��Y^����z2=2�����Κ�Rg'ʽ;][]�t<rR=��4��_uC�}~�7Ģ���w�ˑne�ٕ�v^�1��.'�̙��j��ӾK�����+����y���&3G���C����h��C����b�����)�ٚ���&���do�;�0a3�e����[׿^j�y�;�%u��\t=�
�<�L�J���+����		�1L���떜�����ۊ�L�)�}+N���r����u3�ޙ��u�<緸1P;�i��۾ͩ[��W^��ڱ$
�A^;su�2�LLSU�u���%5%��O�~:٬�bW�Vu��䯲���}�\x����x�"���dM�=���0�=]&��>���Qv�y��!z����;Թq���U\[r�>�����G}3��y���^㧯�R����v�Y��DϢ6�4���_�CUS�=҄��~���2f���$������[O�F򽙱uǝn�)/B�3��X�L��|�,�d{"��2yW���ۉ�*8k��2{���f��L���7��G��`�D�C/�ү�+M��F�o�V���+���v�#q��q&�E�{:`�Y�Ndv�Ě�|f��)�y����������X����� k����Ȏ� �V���<�!	�ius佫�_�kۜ9��fn	l�z��*f=��K
2gY�ɟ�Cx#����^8�d���9��W���/����xu���ѐ���Z�˕�:��}5�z��)�<�^�{Ҫ����3�.ΝhL�VU�^2�
�+�(�m؏���r�؉��ӏ9uͅ��a[�f��pG=Җ�R�~@76n[��C:���Ic2��}cQ�z�{�^`�ݒ�<*�,�%���%�T�dT٩KSU�شs̵��Hi��/u��wc[���hø31��TK�\#�Q�J]���^=����𸗊ؼ�Uz��z���Pf�^�Oi�#4T�g��z}t�z3լ�٠Ѿ�T;��#��G�qȏt�'����+jYx6Hl���~�S{S[Wuw�����U#+���P�>_l��/�C����a�C����^�w7�f����Ln���+]u�G�����U!W�+�a�.W�fς����%�x���m"�$]�=݋&.Ϡ��EE>��һ�_{}�*S����O����R&&�W��-l�@,y�ኂ�B���d����'6�XI-���ǲ�����=�nJ����)BW6}�o��S�T���8��zg��?�v|�lwc�qZ}�
B��^6_�r3`���o�@�U�"�cn3h�x�H~n�o$����ϗt�q�*������{Z�͛���q�Vc;@W�W��e�x.3:��g�{�����J}�=��+��ft�I��X�B[���������'Q~���gjl��<�pWO�s����[�~8q�S�Ȟ�͜�'Ei�s���*�ǃS��<��O�Pm��-�ǹ��N�|<<�ҠCn�=�y��':��y#���[��+�Y\�y��mB�dp�KwNW\�U��DL�������o4�̗�"��ħW�������]p�����n^뷍>���	0�F���Y|8�N3��^�>�ݳ�<��Τ��f�FW���O5���o񩾻�l����\�!�p���mV��kk��r�;:P����vj�y������[��5k���a�@��,s�$X##cهc�����C�[�վ�������4���,�G��iS�X��w���:�kl�m��Rf�]��~4��qP72��?_�璧��E��q���߆r�����+�*�0P��Z7��-�!r^���z�U���K^��惾.��=�~)��O�������YN��5�U�u�37>�oFr��ϣ��vEV?T�����J��~s�����aP����ll�A����v_{'��5���dz%ѯ�*�o*�a-�2"ԯY�¯�գ��{����f���g�Ta��Q�zp�y�_y߲<�MCQ�Cr��~���J�,9�}�0�EvE�F~���#������iA�T��ޜ��P�_��ǥ��\a��  �NҚ_W��=y��d��ﳯ}�|���'o�a#K������ep+!�� �#۷"��9"�^����`�f���Z���1G�+"���`(+�����;U톸�a�7{6��c� �nO�DM��{n���(m����y�-����Ao�YQLɋ�������є�
�� ��D�'�N���*�!ֳ3�c=�k�����K���ޭy%j��`��Uʏ��E�w>��s�}����Q�yUx���>��VP�<�	�~�4F���"֢�n+з{��Þ��:������EG���ρxR�0����s��8�r�u�#��74��,��.�|�v�>×R�웨{q��]�O�I�t��c��,kT}q�V��8};B���Qbn}z�r���G}�7��=��k�?-lW�'����������z�=�o]�H��bU��,����j��C�Rw��������I�ꢎ��C�g���FmV�w�r*�1���cOh��θ?wn,x�Q�%����ȿ������G�}3�4�N����bdS�{��ٮ$v��t���o�W���|����Q��
X�|z��;�{:�\o��y$v�R����r�@�ޭR�k��ў����ɝS�Bsq�|v����uϏq��P���o��<vWG�L�%��W�ϽӤ�98
��&�X�ɝf�&|�Ι
�L����^G������"d{��ۦ�5��{����X�k��#��L��N2�"*�
<�~�����u<,(���HyE�O��e�C��+dW0�� �;C��mK˱��d~7#-��-
���F����!�h�ʒ�=�n^�vӦxr�+�b��Ev��ܓ�%9i��b���cN_> =m f����a�IV�X��l��䣼�F�H�o�m�s/)����;K�k�xFd��9�5���P�?���G\|�a�z����̰d�d	��
�+��]������*�&�]�>�[��R7�'ûY=��x_J�˸�!��(l�E�4z(Ŭ.����엠�g�>܈ڏ#W�P�%��>��/�p����п��Iy����!<�d���������*�5��eI#�ҙ�|�ә/Ƣ�W+��ģp�'K�����y)G��o;2�Q�w �f����4��@[� pY=Dz)�x���Zwc9z���}J�1��K�+<}���=�^Q���y��;���c܉��M* _Ң|�g�uo+���5[F�\��@b�*�,\S��T�ob��gf{l�:z����}7py獰r����y�en�w���Q���E{�f` �y���V�X�F�5�������<��P�s�y�(����p4=�~�ڇ����0�#���gz�Y�&}Ųf�j=��xl4���5,o�Uh�j���!%�U���n��=�ݼۃ�WiW{���}��+��ٽ/Ǥ���d{��3���}�q>�Q¾�ez�C�������>�[9������d��k6u��ܩ�9s\]%[�~�Wv�QZt�,�0�!i�`մtʺʟ��)Ҡ��N]�<�1��iLH�+�]�tM�N�F�5�����}3��f̂�
�կO5����c�U����M��S��G,�8d�3��k$O�� n��o=l�=�F�V�abp�k�����`m�y����X9�����@�jW��/l��cˋ�^���u�1��Oi��I���ZX���d}�#�}��
�������fǷ˖�l���p�=�;>�u�1p�E6s�:��i��]1��=�>	�B�l�X2���7�9sC��qJ֝iב틟9��w��(+�}sjr$�nnj8	�������ٔoj�2��nǟ%���w�״�W�U����2!N�g���"�����5я�?\�R�M>�n} z/޸|��}�A�w�����#p���h�w��n%����e��y{�u]�G׆MV(�v-�G�;@kȪ��*���G�XJ/�CO�ٍ�t�>�t��|���t����?�sˁ�٫?U�|���K�4pu�mt���(��V|5�,yg�L����_��K�u�7/ޒ5�w.�P���#,=��LM>�i���X�Ͳ��{�O�,��]��c��W�z����z�n�H�u�p-U��d���/��^2���E
�/������}K�6Qb�iW4;����rS|��W��\�klV�g$1�v�n��|�L�0PMݼ|z���i*�i�t�!�/3K��p���y�;�Mܐ���T�p���p�ڕ����̎��u�%�꣹�F���g�S^7��=�5�o�`U��n@G�o��Bͽ�޶{�{saǜ��8�w�+>"���i��F��4���p׮l߼�#���{����]:e��xl�{wet	��-oc=�O�n|6�ͭ
�w�ke�35_�|�e�t���
<�N��=�=��Mxb��宿M��/�T�ǏOὓ�}y:+M���m0'�W�j��j�ݺ��V7�"fn����L�ɡ)e1��	�>�Q͝�yy^���l֝d��mA�9������, {u�U�}S�!瑭x'��z���3��V�;��u�q~��R^��76�ƹR\���R�z��s�k�޴�R;��B��{�80���d�s98b�PsZ)�g�|��������/��co���s�/�v�~��%{������}@S��������[��_{~��&Ҹ���)�^L�zr9:�7������.�>�q�\k��]�xȣ�ʱg�w}�k<Q^�).@{�X�SȊ��,^L��U�tf��w.�g��Mw��`Wi%����B�ˊbۮ���Q2�mhޛ/�=d^�0�/(�PSU}�;*{���z����R���n���X�%���伫�!<���'�E%�x����M��kY|��U�R�u�ڎNۤ$� -�ad%?��+��[3��$.��-�q����/6���c��f�.�}�UHʙl�h�9�,-�W+��z�>q�w6�̪�x����V�q�@�z�p��k��di���*ۊ��Vv	h�&�z�*��Lq��[u4�����x9H����/>�Y+�e��/��z�@�t���X�yt��4�j77���a���0��]��5������y�X w�DM:�$/I���Y9�����t��n���y�$z+����� ;<�f=��w�<m�IN��V���M����4{�<�j�Ⱥ[kUrwDzz�h�D�xnzH�\�2*5���i�7U
��}�1q�~�Js�2_O���^�Η+x{`w���f-G�25�O](��>��}*�~��,k�=IU�c�9�B��ۛ�\=��{WP���9���v�Q��7�#�����0�g�z;��ϼ[�x�&��wԌ��^�PўY��S��q��U���ć`����S�r&q����xo=��`��E�8���d������&}�x��R J���%���Tģ�̩_�`x'�c:v��d^�R_j���C..�O뱿��[b��yHf'+����-)�n�\�k[�B�v- ,Otsj�`�j�	nLn��[:��0�Ԭ�E7\���hܡV9	RG�w#��e-�����y,%��Y�A�:�*���F����n�ب�>(�8*>xv���x�c���P�D��s�3�
���	��Jѭ���C�������Yb���53r�Z�J��m̲r��C��cH����bT����K�����cl1Ȏ���D�6L7��S���Ӝ]�GwwX�HA.����vnWYgj�=6�HM��V�y�*�X����j�u�#V��ɮ\�vݧwz�tFiwȊÏ�
)�q�}�'�r�a��)��.i�K���;�M:OC�v�[xٚ�i�{+�d@�z�k�����e�?����I�{
�� �pv��9�����AYt��%;�����]�k!���`c���%d���2�ֶ���';�C�_]�Dw��<)
vnՄzC�a���*�Z�]�e�m���R�v���8��у���v�^6����g��6����a˙����d�������Ա��`e� jY<�}�D�9��u�z�����t�o�<8�)�4��詼��샞J�wIFq�]B�&rT����2�X�	�a��t���u}g��P}x�Q$�nsg�h�u�����>IwV�KM����Ӓܹn=)�-�5�Ӌ�v�@��#��ڻ�H�CQW��[�RX��cn��RjU֝O����M����C������GN�Ik]�ޫ���2����]���q��6Ƣ:!hGкT��Ww(,�0�NF���+*��4�wI��eWvI��)E��������+Tw�%��4�A��l�.�R�A��K(=��f?��jYv-*�!�}]q84պ�С�ks]R�ݷP���7�F�<���@�K��U�nu�WNo5�Si	�A��\ ҹ�nh�Yo�?h7��@����(�M�~� l�;	�c��_dla��Ns�u�t9ވ0uJ��z�$�v4��,Rg����KG��#��ۭ�iV�-��v� 2*�y����.>�s6��ru�1�[��\׼ARAn4k+�������;ڵ����I���������Q:6&ej�p�HnwqڋfpJ��F��c�N[eݽ׸���/3Z+)��;vi!��)�������[}k'�mY��+bu:��ċ�-����1=b�f� �����%�
ۘ���N@]C]s*<�z�\����ba��r�Fk�ۍ��<�5{�(wom���%^t	W,�v�qZ�t�uv��u���iQŋ�4�K��r�q#�Y�s��Ï�����]�q��jڽ]Ow�-���c�h�hsg�e����'ԩ��;�:�U�;���R�uX��(�b�"�Eb����GiX�,��ƪ�Jʒ( ((AV��b�H�(*���3E )1+
�aZ"�"�&$���TQa�111 ����1L��تb�,U �+"2�1�"1I�)*
Q@U��A��!+$����DPDU��� cF)��q�AA��D"���Kb �2,�DE-�R��((�V(�VۉDq��HT��iP��EX�"1`&P�b*���,�&e���Z1d�*bV*�U-*,�*1LH,X��X#"�Y��"�-jQ�*Vb2Vb��ɉ33�S� �QU`��AH���T����� R)TU�-PQ�~u�|\�gucN����M��ض51��1�Ej��[=RH4�'i�N}��w��l#tUN67r�w{B���[oaR'7��p��k��+�V�u���s��3�G�f�.�}⫟�7�j��{n�Ü����}՛\muo%��^��Gѕՠ���cj#&��'}1��'7�G�����7��$��2ɭ˹�J���V��:�r\��Yf����s�[Z
ʬb�X�ɝg	�-GL�Q�|φ�����3�o�ޤ��a�<�����vyQ���ED�e��U�MO"��{&X^b�#}F1N�H����ޥޛ6==ף#TO��C�{������:�d?Q�͹���&� LSt�
8�$��^�kɭ��YUﶡ"��Ert�����D`���S-���ޚ�;/��&�E�zl�T�6�>�^�'��7<��چ�E�T2�Ix�:���'EG��и���%߆����,�A���{Ԗ�ȁ��dOǧ�^�ә��j���5���o�E����7qȺ8s6�sf���l�@�$|�O���۪D�S��ѐ}+N�b���d���b�Wc�Bۊ���4�&�qyNm�6gΧ w��K�>�ʉh񩇗>&:���q�û���FɟF����fQT?6	���Xb����8:�yOyu�t����v�\6�~�X�Ck��<�ϻ�B�>ŵ+P.OU�x���T5tW��xJ6�3��u˦�4�f���4nFN�d�����t��t��!���]Td�;t�%�N�l�9��Ѫ2�f�3:��T�����+zO,��!QU��!$��hz;�Z9��c�vM���W yߍ fg�uD�Cܝ��;%+^ۧ>~�=7Mvq��7�TU{գECvi�������@y32/Ŝ�y�(����p4=��$Ò�ו)U�Q�i-U����{N��Ͼڇ�P�e�53>!}�'��+�؁��o�IG�@M�y��sx��켯9^#l�螔2�ևq���zX�L�Ip'���0s�o�t�����z���W�u��>��'�n=BPӲ�ٜ+���:��OG�א)e{}<$��l?\Tǩn�������P�~g ���;���|�w֑�,nL��5�T�h��ԉ��:��<���]�o_= {9����B��;�r�=�-���VET{MF+�.2gY���/��\�0���^zsVzGfI7��w�9�^G���e��s��(+�}B�۩���MF5W���y	ʍ�ޟںL����q�F�&PL�sʇ}R��w���t�{������NQed?Q�6���R��3�s��v����8�V��T\��y47�w]$s\��{��>�W���ʿנ��)
��5'|7��-Օ ��ʁ�����<!�х�q�Q@���]ΩGp��>A��v�ٙ¸db�"��1��s9�T++����:r�7z��wVx�榞w��B6���K9tYC%"�:�Ov4����^'8Z��8��l�}w۝.�(�2Cg�z] �"�FT�`T\��}�,*�ξ��>��DG�&�޻ٮ$��=U�>8o�*�t�>`�x�a��T�_L��>.W�dl�*���s��q�@���_�'�t{������$k���D���w���n�R&'���8KGwZb�:�[�̊�Umd�{~#=����=J��������� S�
���7;s >5�1����!�Ve����}G�R=��Xj��yU���<��5�?m�Q�� \��\��\.=^B�lY��+����5�
��ɭ/O��qzj�P��9���Ùc��;`^�f!�Q}�Ω��k�[�v��Rm�����Qxd��������x�0����25U>��(�ӽ��r6��A�ُd�>���������߉e�Q������u���}q���޹��3��#�G�ֽ���NrܥW�ݤ�o�z%����dО�*8b���k��I�t�ý��qc4�� o���uh&��[ӽ]�v�U�����*���	�5����I6s�T<9;0�5��$@����u.57�ʀ���K=�n�I�p��Un���R|���y���Pngs�{C�	u��:���G]s�iH��2��}��o��J=�����ƍ�]I(�#��`�|fWy������]6����&�v�s������:jl!��:a[��u�{ւ��{q������G��Ҥ�N�w�����`�5��P)�}�w�w������7���T{���؋��q�^�|3�h��}����=痦�_l�� ��k�V�z��2����_s�㔻��\E�}��+.�b���Iu���|Տ}�O\��Jo@T���q�ҳ���q���7����T=V�v9%�>���o�y�!�Y���;7�t���FTL�@�R�]dm0��J}!ɿ2�r��%>���.J��~b�+~��5�����
�M���!���T�U!
�^��o��.8B��{�>�#���W�uU�q�^��}�R���������ơ�#�\{*#�������Ζ���������~+�a���x��W���� ��[��� ߳�>�3��Ie>�/v���tD�J{N��wO��.���gǋ�����Y@'��D �|��Jvw{{={�}���S���t����#����"����@,eD%f��u鹠����_>�O����3�Nv:��־��}�}��l�xn����a�wg^��=��C�/�O��ge��l/8�w�s�ϯR�������tR[�_���a�+y�l��G{��O8S�I��;r"ަ��կ^�1s�z��\�y�w�
V�f�$�4�����_��ޭ�륾�D�t�y�2XL�8�O�{?��9\3�G�W��9���Ϧ��V�x|:O}�t��c�;�٤V��	3/���/*:=�����<�5���Ԃ<�*�����DOT{�2�L;ͯq��eNWOTU�g�ԺO9o�����~Lψ^�Ry�d��i��I�ꢎ�ǵ������?k5��rOYjv����V�����S L-�xB�Wx���`�z��\?h�{G�O�ȍ��k6g6;�G�w��>�R�\em���S�F����������ǩ�����W/g3��,�Ǖ;�Z����ݴB����WUxn����29΂=����7�V�R:��i�>��==���s�r����خ=���^�d�q�ւ�� ���.2gY�|�Q�!w11�si	�� ���K�qc����{o��7�\nG��|ag��T��:���n�T���˼b�'Օv��߳���;1���ׂG�y��g��~�c����.��=#�5�@6f.��I�3�\f�dow3t��zu�[0�Q~ڇh�H渟q��Q����mK/#L��`��F=�f6ck:�M�",΋+� 8�$��fh=(�Ss#�f�5-7|�YTlڗ~⸫vC%{Z�u@�d{�^Su<��aޮ�����t�_p�:jt��+Ԗ�ٚ���:g�;J�u��uc�z��W)�Yrw�����"����}����w�����Σ�����=�8�8p}��0^n�wmɿ}�F���L����}���}��%���>>��Q���n�n�����=w��^4{ԏE��$���
n*�3N{�@�Xs�2�z��$���a����Bm/u��z}����� wwߦ�:gT�C���11MVѽs�ݜ�����.��Y�w���>�׊����K�`{���/	�fe��S=��a���������ݜ�r�O��Y�ƎT%�j�|n<�@yds���>9 :'O/Ux.�c5��;��O�v3E���"�zGaœ
�V�q�5��?O2�2���'K��y���������ݓ-�~]=�hx�ލ�!i���C.1֏a��ߴ��^��3;���U,�^�u.�۾�KyG����!���h��,Y��c�Z?,�8ҟ
�z�o��5k�����H��q]��0g��tgqթ���}��I�������<�{�'���2�2kKN��k�5�Ӯ�����4.��Ň�.T��ȏx�V`��xl������'��j��9Q�kw�w�L�Ƽ�7�~R3>ͭڑ�5i��oN��۟��A$�E��,9}]��F�v�S��*�9]��dj���fԬ��U��[� �Ӽ�n�'��.�g�b�މ�`���-�~J����/�<:�����F=�M��T������{��լ^Y�c����·��%��R������:�=����7H`��4���T���p7>�0�pb��/jo3���P�.�ü2Ѽ�ax�sʇq]{N{�x����!o1p����f��6omy�՜ȷ��t��p	��_\�9y�A�W{�|�o�r<{�>�qDl�є;����_�ov_=\������CgǤ��FTK�\��}��«����6aU6!�yVןP�[|����ϼ��yN��mz�`�Q��۪��^*Η+�3g�pM���G���n�on��{j�,dy�.n=�t�{�+�Nnx���0P{U"bb�W������}W���۵�R�;~�R���q/����
�����!���9�9��/n+xLӪ��;Z���;�=��ңq[=�c�w�K��2<�_�: �¤ U�Xo=r,���͔O�'�[�w���g�͆6�6��_�d�i��Q���Vj�׮l�{΀�9��zt5^�>Ϫ���`#45��e����ou��&�a;�η��s`g�9�_+����wSn�I=��*�U�'N�?�]�<{�$���������c2?	{;b���������w�N���5�]�Ѳ�F�uqb
V�)]�ث��O��'�FXZzn|6�kC��w�k�4�֖=Ifd6�Uza�y�Z�6ss����|w�pO�j���ߤ���~���ǧ����>��tV��?���eE���i�O��������h�j�Y�=;��?mΘ��	�>�QÓ�2�ŋ�6kM�y���{�1� ���UkP������@��p����Uᣡ���dC�=��Rp��P�ܼ�v4����oz�v��}��^�o�w�#�n#����������{m�4�ܒ��{bbu'zȟX��Z�>�`�s�<7Tz��6=�q2��~�a_yK�]�u�C~מ��D�v��W�w���/y+�A�3�d_z��d�s3���d=}��?K�H�r&Lu��C��Nr�Z�z}��7"��+� K*:�U`�O"+��,\d��U��c�gʨ/o�$���ﵸv��>�W�	��c�'ޗ@'2E��dEx��?�(����qBr�SsWO<�{2�1o�v�y	\{=�F���~����f�2�:���B�D�6 �3������ND��
B��Y=��s4.DWmC�V4�LQ����ǖ��F�i��;��SU�ۇ��]�M,�t{����g�ǹ�y>����r�p��.���(޽��3V�mf�%�UQw���,"��zO2���[*�nT�S���t��M'8,�H~%��3������ԑ�{���r4(�߯�G�ơ�Re�r�u����Uͭ^;� �O��4�����f_�&�o�}/��9}���~� ?nT��|�����ŕy���k�${�Gŋ0|2��&���Ȁ_��Ȃ^����<��o�Ϥ�j�0�zܟP7���yW�~���*h�@�St�^z��\�2*5���@,e%f�ͬ�D�y�\��fF��y90���S�꜁�r������G>��#�uo+t�����5�A�/}��x�k�1M�D.}��ޫ��㒹�FG���P�4�ʐF�+Ǫ|6�T{�2�L;�1���3�U����j3�e�@϶�c���3檧�_����~�/Y�6;�'�zd���l����%�ip�,>K���i������ �Yn���]��1<}w2��hDR}��������[w��L�a�Ӈ�և�En�;RϬ�/K������X����wtU�Ľ�&�̏ʼ�9[˯�>����o$������T��5��L�/\����#�|�����y�wRs¥e�Fdfm��6
~{�q���F�P���o�h'@zt��i�]��)�5��Յ9=����X��o�*U�H�B�o8��}w�o�n���m�Ϋ�����O�y����;�xP1y�'��]�^�Ӯnc�Ԣ��wg�N0+[�ʠS��6J]����|E�{�ǩ���l�*!��-�u����"�X���n>ɟ"����/E��E0�w�O�>ޮ�g���{���q���Y񅑾L�:�e�}X�� 3�9C�N��W���FL��^����^���O��}�������:�d?
���̰g���W^�[=�r���s�}��P�l��j5�뇟"鳟����t	�޿[��\��]�g����(k�]�+�|�xt��deD�Z��h�va�[��Wq�G�!g���~rW�ת��V`Ưr����P��>0y���dL>��XZs>�~7�0�5����^\�����U��U{ý��,�?��ҳ��DLW�$�����͊�L��tdJӰ�ǽJ�^F���E�;cs���������3�ԭLde/L�z� +~ۉ��^�ʉh�M�=���LM{��ו�L�����^G�҆)яm��8���VO��Mxڗ�Ҽp/�����X���t�;^s}�+�����D���<���='���^+��LϏ��w����;@W��������SW�s��V?ܓ��J�꾻�#��=�����,-�|ާa��M7'ud}SGj��Ð�f�*��zN��}ڕ����r��w&܀}{/Rc�=#M���q�x�X�cA�n��Z�֜�,�:�|X��ٽ}w��v;����S+��C���z������[��n���(nL�Η�s;�l��`Մ��7QJ��S_eH+V3�����
uma���5�/���肺#���;���jm��W� %+�u���1��&.����V��iM�n/t>�C%����g.9Y�־4�e=��;�1@s"[�N��/]ٽJ^��4t��m+�U*U��[�q��<��47wu%�"�I���f����g������aޠ��pi�(7��Rŝ�Q̑���@ �V}GdX�|jd��u.���q��vn�5̋��o,@:����\��Ht�&��[�q!� �aӾ���	�]� �We�>���9WU��2���[�jf�
-@�{2��-M�WZ֚毬���u[/�����gV$�ɻ317������1o{x�ժ�X5��q��y���Y�$���3��[/�ŷph��\��Zyr����U������EK�����\{+l��ŎQ�f8*��e�ꡆ[Rouj�("F^���v���cNՇ��
湎����A<� �+��o"�Ѻ�n�s#X�V@1,o�N���c��Wz*ĸ��{�fú�5XF^��#�)�8�&�2���^�]n�+�d�;.4��yކ�s�Y�eC��͝�r�]"��Ro_fC�:�vy.W�p�
�VM�_gpλ�u4�Ջ��=w�������:�oyH*��40���wmn���:m���G�W�`Pm20���b�u��4����'!B+����g��s���6�-��v���X��O����fs��%@g_-۽[�w:Y��m�0�>��(���u���ܳO+���
�%V>�����G����6��[�G��=ל��U����m��N �����Ԃ�wB$\���FsB�4��U��t$�g/p��gPG�sW%yS�8t������'���\�w���X��&��z�khu���4�H�\�e��L�]���*�Qt+
hǹ�ܬ�ι�	1��-��qd�v��HﯔY�0d�jl������z���us���v}�0>敦���*�j�c��������n�4���f�AB�4U�#:չ&�}A��ӎ5S3>���4�M���n�!1&���u��tAU��4�i�z:�%�;w�=����nv��k���廻'�}[��M�
�ܾ;�r�ԓ�%n��5���}մ��폹�=�E��*��9���9�HT�C��_���Z����t��.����|�-��gz�6��q7Ǩsܮ5�5i`��eO����^��]-U����v��g:AH��^�*�d%�R��r�>$������bB�(�)7[*�F��bJ�@Ĺ@cY*E�J5r��0�kb�(�Kj�*� �)jԕ����¤a1R��)Y�Qc�X(���Z ��V.e1�`�V�3*��Ŋ�QdF
�
(ĕ�"�
���X�b���ɈEYPD��"
�E�
*�ed+
1b�$F*�X�"�#JI�
�01���-�������(��!��DA
�RT�µ!m �`V)J�LHT[�X���LQq�@��+�jF-̕1�U�6�*,YE�V���(�V�bI��0��c
��k%K���aQq��T�J�m��AekP<�y���-��p)��=!&���٘V6���!�|J�g���9�xR�kg���۳Q��e�����	������_�7�ɽ��瘕��3Q�ƾX�s�a���<5���|%�bw�	n��y�{S�u���碏��L������=8\�tޖ=�7X+����N[��P>�j/��V5�ӧѝ�q-�:� ���	Cn'i���kJ��
�k����
2�LQPg-�k5{�z�w����Sf���}�F�����'
YLe}�ZX�wǦ~�͌�T�g�{�܇�]�mm��/�_��\?m����a�	l�T*��}�o!�G]�Y�������2e�쎩u�?_��{�yط�#��m������6����.*�k���'��P�Е>��?Sw��2�n2e����^ӑ��߯���������w��Ԭ�u���6|���tE&e��dXM�
��r�����*�$u�����S4���ުO������k��j�{ ���r}R2�]0*.X�>͖E�hh{����G��=1�����|�צ5�N��t�>�u���26b["&H]2�V��x�npF��)�o�P��N"��+�L�̡�e��I�B��K�Z̭ԍM�:̝�U�*���~�pI�G>SMe7���p=z3W��8�L=���0��1����M���M���֞s��];���3�ە2�u"�B�ns7V3�{u��ګ����VD]�E]�fPQ �N�H�Geh�/��E�ǶHn���0)�5
�b|͘<�R&=�����ʊ+Ƌ��{�7>� &s<%J{��ľ�g#��
����w"E����S��=�뺸���m���0c^u�o�)��0��>��_��:��� *~v �Y��qM�+�s7�V�v��N@�OR�͏���!�_�d�iz}F��5�Vj��7�<���-�G�ea��t����ލ;@W�S��.k�qɹ��ͭ�3k�j6X�3Q��%wp�,����W�m���SK�90�bN���C�9G��%�����:����;��:+N����z���X�ќ_���U-U~��՚�7�L/�V&��۝1ހ{z���;P��ō�����c�=��3נ����>L�� k����ʿ/���}Uï��_���}��_�z+��z���l��G�U�9'�������m���g������G��v��]�վ���|��q��;���G��W�}�����M��*}E��Ub2g}7�a���o����>��{\_�;�����V`�x���j�&o*��ˇT*��V��e� )��7_���fb��$W:ϧ�6���%lo	:���֐�%�i>� �U3R�Ə>'r��W�H�.�^��n(of�E���׷�\�:��x��!s#N�SA����l^�n�����ǣ����������W�@��@������C�S�Y3����4�wK�q�<�*���x�_{��]�7��&��7��)L^�w��/#�@S7�@>��3�ygȱ�2��hi���U�LM(�*\]��G�:3Tz�����/=q�Gh���)��rْ,�� ��4�<ˏ<4�œ�H*�w��>��1~�5�{_�����!���5�1-�\�CO�<�.�����ӛ\��(����e�mCU]ŋ�^��G�ԁy�#EG��и������O+҅���J3Z��[���@�l�9�O��-܁0�RJ���+�#���7���/1��7ļ�H�ܾ�s��Z�I!��é*"i�i���r	xk��G��W��P�5�8i�C�Wc<�R�n���U��{l
y��"�U ���n���3�G��21��l.��D�M��~���=\}�~V�&3��	�e��?NX�}%ѻ���7P��6�;���/=�G�|��ɚ�wm���@ϣk�5'�a�>������顾�gnA@g�}�N�{|n�#���inT���eG��Ѽ��PU��V[���=��'�JT��\: � >�.�b��l[�ҁ���9��`7���־N���k�+iVι�b�NcF��#%���Z3�'D��m-�SO#Q�]�����f�!�H4_�Z67Y�l+�GW5;=�R��oC}��f�k�	�~�����Z�%g��P�M	B��*x��g�O{^d�0/��f��8^�6vaY��
�g����`	���K��#<��G}�R2'#��F��V��^9;��ҹ�y%����7;>em���S������|�	V�<]N[������o�$�m�C���9�u�9�O�8
�c,��g}1q�Bs��e��/��=���Fm-�=�`>�:�=ƙ�=��;"<��7���[9�kAS6E�x�dγ*��/)�Nx_�ˡ�3�����~ِ������>�����/��G�c�w�S*M������S�8^�Yu[wӞ�/l��zw��2e��c��`��>����^Zb�����U{��i�&tZ?���5�ސ�j2�����+��mCF����t��\���ᢡ��~6v�.���Ùu4�=�����C2=����9FFTKv�����f*��ĿZG>��#����WD���nc�̮A��g�n��˒�F��p`�v�D�>����4��P�_���T�(S�Ec��E}s���EK�36L��b�*��n52Y��_ɜ\�����Cvӈ�x��u5�$1 M����s���W91<�<�m�S��k ��>:h:Z1q���Y�@�4��g7a�H5�b�:���ò��b��d��::�4����!W��N^(~��Y���Of�h�uNH��l�A��R&b)�x�+D�����I`>[��O���z��W����}&��ۑ1_<�I�%D�w&��ex�F���O���//��+g3y�ur�;��^�W'��O�~8|�{�N��ˀ+�<m�U^G�հ=��K��3�wq�g�w�OL,s�{K�����P�d��Ϗ�����P�r@�BA	�3{��n{lx�Y3÷�f��q�P�g�t=&TmC�N�6��~�Bx���<��W��yB����1�2f��	(������e����x��=�7Ł?-��Ǫ����ݒ��:<�-�. rRx�VTk�Që�	�>�P͝�3�]��Zn5��N|qO��q>Gޢ���~���e-��;�$o���n7�s�/���]�>�Ië*���&���\��6�}^۝�y{��ej�X�#�R�ꐶ�m�*r�q�|�V����9QF*1M�I�%	��}�gf�9O��l��˯���72�}$1��^��μ�o����u���~�H+Bٕ*�]L�˟-s*I��_U�NgY[���MY���'W	���Vd��Z����8�Q�pD��Pv��Xr�W;�ܵy�rړV!i��v�\���[�2��I��[�qI/tt]�.����-k��yû�(��� Z�gX�ޅ9fr�S莩��rj0	��p��o&X^9�'�q���r<W���_��^vM!vkl8����d��E%5Ų^�4�nr�1M�
��&^F���w����]$MN��1YU1��
j���g�^y�������#�Yk�$6n=.�}�R2���G�6XK���v�9��=�P^�y�~0�*�_���e�����r|/옖���ͪ��ex�5��㙖:�_��ճϷ�}<s�(*��.{��������$k��č�L�,��6`��'�6����u����}=����܀|<�q�/f�}/o��	��;�)���;�&���D�ޟ�<E�Zx�o�\ߦ@hձ11K�h�~;�&��k���W�|�&f�
}�nL羥<���u��'R�r�g��co6�w��8QQ���^��*�s+��^�j|��^�}�wz����\��W�#�s��mhx��6���y����~
M^\�(��W]�vnW�,�Fz9UJ��֢����gjl��,�*#�O�Ȟ�î3kG�*��}�=S���@8_�D��RŃ:Q(�ά�t#�b]��]��/m�k�mΆ����C��T~��cƃ!�dhXm�ё��v��S�4���-�����Î��R�r�]�ۣn��A�.������z�
]�����!��K0Ԙ3��W[�͞(�	e��ۉ+�u�̜;���@Ͼ���y�p=ҥʍ�Չ����L_���4��Gnv��ݧ��)��w]˾��ď�K��kN��������d�^��Uî7�~7�g�	l<�O�Q�YX�_���nor��[g�[Q׎����@��G�ok�9k���_z�u}�v�b�F\�"؞����{����{��=�T��G�qUCܙ�M�}3}2��?_��_�烶&}��Ӟب�p�U˗����W����(�P��]``���/�P��O�x�9��>���~�GI �ޅ^K������>��<o犣y�,��Pͺt��&*ygȰfb�Gg���{�#7���;�����q��+��K�T;��k�t{Ҩ��UH�X3�}�rY�*9����,����*�XJ�Z<�����ǳ�Dk�z�à���<��!��ʙq�+W�zs��w���ފ�WӪ�>��|�ZE��^��Dy�߶��O-]��k�`V�ᗝ��M�>��G����$�e�{A-�ƗuC/��(�+�U�v���M��Ǒ��S�.�_�7�����gޘ�89�v���J�8�l�'[��� ��_h'����!���]Fv9��۠��
�m�%��L����zT'v�U��,�b���K{M��V�O�E�C.����5��V�[Aĝ�8�`��Y�;2Q!�u�Z�ݫ1R^�{}�"�˒5:>,\>MQN{N�@/�t���j��{u���������!����YsL���H
��{,
�y�� ���t��z��}r�ȭs�<�H�B���+��d�yz��_��Y���71q��9�r���&�μJßE��ț�{y[��r ^�u7��Y,Ǯ�ngn��ʾ�=!I��@�F������۹�FF��Jr=顳pՐD�+�������N�.��q����==OL;��|n;���}����~UO��u)=o�@���4��Θ��s�w�Z{|���u�h��������k��Xw��g�:i�)n;ק|E�/+�r��^:l1~��'Z����ߘջZ=��o�U��,^�V�,��=��������k�*{6�E>񂶼0��o�����Q �����FD�����v;3֟�5���:#\��Wz��r��b����z8�h�������~ב�]E�{��l���*�=��߮�WP�e[���2������K>��l�鐫L����ב��{���q��s�7©��S��%�����K�ݬ���z��99��[O�e���ٝ�������Ύ�u�k5�1�}yؔ\g9*�d��C��ˑ޾ۥ%-�0xM��@_)�b��9��[ή��{���f�k�0-�Ё6�ո�޹����f^C[1q��c���;]�iѣ�cc�:�ғ3 �Z�T�{����x�������;��Ya}��z3��Ey�>��H1j}����������!BF�s2&�ң<2��3�kϦ� Rr"�]d���/�P�K�~��r*��y������.��q?i�~�Eh!��L�=Ӕdan�;����mCF����/֑^�@����#�k�����}��p�m��x�Ik�2F���TȘ.}��Ni~4g���{G+�8��ND��R�N�;�)ZDx����:_��F۪r@��Q������1N{�FĿGh��@���]�_>�W�ŭj�d���*^���N �!�r&���-Ah���>��?R��S~.g%>�c�ګ�o\�=����\��׊��C�8�p\G�\Q�6����Sw������Z��I����D�Cی����t���>���ЕcZWu�y�W�9�Ʃ9�u���vvzW��)k���g���D���A��7�0�m{����F�?�����������l���-����UhLd���IG/�D-7��\zp:����/Ǥ�G�۱(��J�?Q9��e
�Y�&�{�u������vu�:���\ä,���WmZ�T�qu���`&�v:źьݗ;�i�̃}Hr��S�,']Z�wڝfWb�T��%��bK��ir$��"Vv΍����n�q���f�T�}	�];���k�V��ӌ�t�ө�빉��8y�N��z�����d΅�>��?gw;~��n���f��tp�P����}�H�{���nx��碻�G�NS,^��1���w��o�}2P�L��H�:�{{i�:*��l_���7�;��tSe�/���ޚ�A��k/{=�M��;M}����gY�|Q��0����r5ϼw/��\*�CFye����q���YY��}V}�>�=>���nrj0
�T=��([,/w0�^��+ǻ,П^x�b�3�'i=^CG���s�Y��"[2�[.(�����'/6h4n+��wyԂìpύ�i�W����Ӻx{O�߆t�}�6Hlߥ���FTK�\��}���@ʹ�<�W	륍�ehw޶�g�w�W3��:}���W���d@��ET����w�c#f+�ٜ-��kG�G0� �~9������S����K>��r��=^�n;����yXc����8}�{;�|��b���b	h��	�=;�����t��� �y�c�@!I?����BO� �!$�BO؁BI��!I?���� B��!	'� B�r!	'� �!$��BIH�$�BO�!?  @?h!	'� �!$�H�$����� B�x@�!$��(+$�k'�b�� ��
B �������_��|P;�� [vH�����ԝB�$t��@	 $  �>���I@٪��I	�̑�I�liOF���=G�dP5O"UJh       5=4%�z��@ �� = DT�h      *CFj=�=M4P �h�A�� ��6��6��Th F���v���QAC�ı���p>�4#t E���IL�b��HXJ�S�g�O:P�����DBP~�8Dl��FA/���Up����vyc����P��b�T�(�β�xOf����L���8��dv��,�б��q�gd.Z�)x��U�̛|����X�wp��I'aJ�Z�`�~��Pi����ZFʩ5j�C×�A¢��t��1�*�Е�ui,P!P��UX[
�VT�3]�4�	�ɵ)��t�\0D��4ț����VA��V얝H�Yj,ૅh͋��&�"��b�0�RղS�����f��lM��0�|�?b�%�b�E[L������aؔ*��Vʜ�u��_ـL�[s�n�UB����i��Q,�*�ۛx�S���v�� �m��e�p��*l�9�����7w߫��^�+(�Y�as��]#!OeO;�h܍�����L�i�c������H�m�a�D�yUU9��;���������Z"w`A�%d�B����N�㭤Խ�1{�yz��l��qFcmZ%=��B6-�q��9�Dk���c��	��2bҗ�r��zr�����;x��(��D�F[�9C^�^\�#v7M�t�'2���dM:{j+n�i��$�M�e�;f�fܱp�-xvUT(�[��3^�׸#iʋP�e����Kb��m�:���ƍ�I�?�����3�rߞ	� ��!�-� �'��ɡ�ieDC�����q�j-;$%���R%�%�"�ۙ�V�ۙOi�P��2N���M�oZ��p]�VH��S���|�ԕR�cf*���M94Y-�4�,"^�)^��2�B���Z��̗���9�LL1�*�w.���؃(U65�y���ʹ��B�$i�;�@��"VR5��*��/�.�i��R�^r�����k��KY-�"d�Z�C��ڪ���W)�%9�kkܹW�L�n�:�3ʕM���Y@��(�PĨ�T�ۻ���l�wڟ�����H�z!�Y��iVK�P�A�t��2�]{r��Ù-<w�R��P�����u��ur������&@��,n��b��w�m�3�9�%
=�T`�T�p&]�jr�A2 )�R|���&(������d�� �1�B�R�N��-����mA1
K<R�ޭYl����Q7];oT��6�⹛.�^�U�z��FI�@�=B�{�!���˝>q�:J�yƵ{2�2{n7K�s�)�w���}� ��vN8�ެ�����G:f[��LzN5���8��^S�`�.t�eg��;y�v��>4�}4�:b�ʪq��#^р�u��A���G��-����E}���ͦo$Ry#!Iȹj[�q*���+8z>������f��uy��J�*j�5�Ӭܬښ�Ww���'�y����ױ?�c�ʺk�	1z,��^΋�S]��%ׅ����NF��D�
E�6������g憎H��8$T8��:f�Lsr'�[qټ�֚��,0��>q��B� �L� ��	�@�2�������Y�܆�*Lb�q=�,�l��/�>��B�ӄ��ZG<��%>qԵ���\�9�ߗb���m��]3	�HYT�"���VF��U�>sw=����I$�=8GOs%��tܥz/y������/���x���m��R��a��ˉ�=��Ӹ�v�r����n2_���>p��M������+�(�l�nJ��{�}}>�i{�K��:F$^M[�Z�n�nܬW�sRw�/{v�1ƕT�+!IBp(À����n9���5Q� *]�*���ہ�ҫM`��>4�%�V���k��Os8H��yn:��U�ǯ�O]y�D["ڱ=��k�{����� T
����* Q�6/*ׅ�{�ʬ���HBN��DRv)�aO�W���):B�&p�P��4h�����2�`�tr0�2h�ӼkG�^yܠ�Y�M��av�fv�E�s�I�R�B�kH�5����f�yYK�]��1O[xx4t+Y)��j(���w"acW�$�,\8%���2h���"����\�dLi�g��Q"�zG���a��]�ʉ^���]!�.T��I�78�j�!�A�[k�勲HRU�%1J̴�6)��   !@$	$!A]�=�N�T����u�h����2!�!��*@�$���H$����X��oo��5�$�&(@�I1B[�A$K�h$�kTTB��3jF��-D�%E�j	 �!�MH)�fI�k��� 9�b��sSj(�F�:�h��Z�!1a�!IB^q�[�7�k�IP���돾�$�u�6�q�;+2������ʆ|	��_�\<ú*Qz)]�7~�NЌC_���NuP��������¸���1�f��.&Dyk�^$g�����^���WS�Ts� �zӵ;N#3�>�=N��ʽ7�eoҏ��U��DY��	ǅ�z��K�T�p ����S�cM�,�{/f�ܭ��%�ROm-���Zq9�����1�� !@$
$�"�@BI��
�"32��¦�=��%���bg1ׯw�o�����A�=4��&js	-�w��:z=�Z��c=W��Ǵ���n!J�a8��<����q��me�
��]9,*$��cXg��j�5�5��=����~[h��+ch�����B�Ϛ�>r�ρΌ��>[JD�q�OJ�����{ﾚ��{����'4�^�K�Ox��d��<�:"�]��A�y]��ڷ6�2jek�b"����շ8w.h�J�j�a�N}��ܛ���s����bD�$I&(I�
l�*TZ�@����x�l��m�q1��c2ש�e8��} YL�E]�U�N����d�	ឿ�>�P�#P��Dm�Nle����Эg�~���*��j�Ѕ����|;n`���f3�N�ޓ�U�K� ����v��^�'��E���2r�P����F�G5܉���3�&��	�؅K�����eŕ:��V[�4��Q��+]�0nt�!�sw����,;N�J�3�v�sOՙ���M�������I���TZuPu�AG2(e�e�6��3.Tɜ�¨�鷱9�;su[T��- L$"� �bbCb�o�7�f`ܚF3bx��_ǥ�ws)�Il�uf$�l�8�ğe	�+���C�lEv.��}Z ��]�j�Nt�S��sÆ^nmԃ�'b93E-�םm&�c���Jefw:�`���
���Ĝ���ɞ�s8)�`NA����Ķ��4o�V|�=e'S�,�erMm�/��>7xn���啫_RwB+��ѳy�g/�e��a�Cr~�q�,n���
o5��˝�62��v�..��S����y�Os1%�����SoV��4$"@���Mվd��gCy�`o�D�`T��53�/\D}��FD�se�KOMVv��]:�VM�-��T6���z����r�M܋u�nz\��mʓ�5	����3"���AL�vƍ�jk6��Or�6&��}݄@M∈۲0B��Һ��q�S�U;֝�uTM�}u�f��D�%˚s�0�����f`�m+���7}z�븫 �x�ѵ���0U��U�$D��&É[ jC.2ę��^Sf扃s�n*Uo�#�U�f�]=�cݙܷ{;�p! �����������g��ed�.�V��d����9^н-�ܨΞp� 0ޅz���ys��={��A�	m�3>���i����q��N��K�륗����3Q�l�P�m�;�l�f̞2��&*(ܢΗI��P�̈�����̼C���;+U�Uͅ�n6ph�����3��o���~8d�=Į�a,�ɣ�6ID���9�vٟ�3�3�Ʒ3j�)��j�-�{�xH�li��T��D]�o;ۊ�g�7ct�.//Z��bu*�>��3-�¢�.ot*gTN)%����tH{�b�}�7��;ͻ�7\U�8�ڗ�*U�������=i�d^h�/7:�X�m�f�$؈[*;{or�t�f̬�Vcz+I�7_Vr*��8z(��4�:3{v��ٺ�7;���H��۱QMv����OJ|�(v��Tˆ���:��7ը*�bba�(qu"�W�����I��I$��DD-(��/�S�"!���$��*���kJ�E�<��󹌗���Q���X�}��LPq	�by��7�+#��K[P}�H�� �0��ʶ,l��_dq�^(�^�Z�����]�T�_AN9P���q4���Y�C�m�5C�V�*�B�A��6�8e�M�Aꂈ}�"����Ȕ�/���
N!0�_� q'��'��ig�W��Zk�� J:�"� 󯥞�dd��o���[2��3�͇�$�=
Š��/p�g|P2�%���3��`��)���.(�D&؛��֮�>V�	�DB�Y��l��"�`h�X�ZE�[��`�=F� �#P!&�XN�#�U^^Bka�87�rĈ݌����C�i=bq��Sڿ'?ڎ=�DD1�iޙe��r�T���������~�s�eY�h
t��^=�{��RL%�+2ǈ6\���G�6�Ϋ2�����z�G��g&��u�!����=�<�2ϸ�H0�_�'������M�n���8����@P�d�i$#�6lN��5SEBpP�Ђ����`o�ض��ͪT)!�a�,�sG�#h�I��0_[�.(�[d30��RL����HR��G3���"��ix{�x#ׄ��܌�0<j)e�e�L�܍�fD?��+v�(�<^�t;'b�ITR�W����!��PG:lI��9�RG�a�j1�j��\�t�B9�G��E�B�ӭxr����T�
����v��'��-
]�]P!{;����4��InU��SR�s����t:�F���V���|��xH$AD3�����T,v�)tg]�B����B�r�]\a�iu"��6|-lE�����	h�ХEZ���"�(H]��