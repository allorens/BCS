BZh91AY&SY+��ٷ߀@qc���"� ����bC�      �/�@֬խ(Q#F�R�@hHm��AU��l֙PiF�X� �l�FڪU
U���j6���U��m[[)Z�Y��ջ\�n����Dl�i��ic+Z2�-����l�mR����&��ةTR�SL��Y(�fEk@Kl�!����ceh��E)���u�eIj��^1"�Y
��N�U5Z�-���STk-m�U��Q#���kl��`
hZƄح�ւQdm�5�m�JT�fM�k.�ΦL���ZX 8   ���BG[s�:����Z����Uk��ڨ�T�UR+�ҫX�Mڷ�N�鱁ֻ��M�aԲ�1L��mL��Μ���1Z�[dk��E�   y�/@ ':PR�a�,��*�tuM
ޥ�@9ɇT ��[�ށJ��� �'� =R���p>ڔ(�;Y�%���X�Uh�C�  ;��Ω��R���� tgW�=S�a�U�R�ފsaJk���=�(7N��oG��%���@7�5��J*�tjӠ������sl�B�2f�l�1	��  ^4$(
ڮ����_}ә� �3��B��:à�R���*��w�h���m }�5����҆�^�u�AA��Tmj�hʶ͵��e����  ;�μ�(=h^��A�Ӯ9�j����R+��M8Ҁ&��P�)Eû�J�T�w= S������]� � �-DF�ۻNA��"����  	���hۭ��m�i�:�݀���N��\�����jt,�jR�<�w�@Tp��� nqnT���@U �v�)�fQlL�3l�  L��R���}k��+c� S�^��(
Fͺ��[`wG ��  �������: �NB�UBTm�UU�m�  ,x �J������k� UX r�@:�8� nsw@ ,�� 3iT MN�R5�4�fȐ�6�<  ۼ_PooC�K  6�ƀ�0th�u�ݪzG��4 =]&��mͷk@��pP�e� ��ƍ��YV�՚0�5��|  ׀ ���4 �'�Q�s��� �t8 PZ�P �  ��� ��8�Z��    P   50T�H	�& 4ɓi���ъRT� 2h    O!IR�      j��@��H      E=�5UP�Ѐ  � �ڔ�&j4�D�)���4yG�l������:o�����~���Q�m�.n	�y��[?y�:�������Þ�n�s�UE�T U�EPT��@_������:TUE�=�/�=�����EQX?�UU�t"���`�J�� �������јO���\�0���&e3	��fS2��e̦d3	�L�fW0��̦l�Le3�L��G09�̹�ds#���G2��̦c0)�L�fS2��̦e3)���fS2���&e3)�L�L�S0��̦a3)���1�	�̦e3	�L�fS29���e3)�L�fS2���d&L�fC109��&a3����0���e3)�L�fS2��2���&e3	�L�fS0e3���̆d3�L�`&C2�̆`3	��fC0��0L&d3	��f0�̆a3���f2�̆`3!�L�fC2�4�f2��&aa��f \�#�Ts(�a�9�0��E�3�aQ̀��G0"�E�#�s .`�L�#�Ts �dQ̂9�G2*�D\�#� s)0(�U���Ts"�`�*9�G0(��3�dE̢��G0 �0�@\ȣ�E3+0�A��s"�d� ��G0 �d� f2 ��@̢��W0(�Q\ʡ2�aE��� �` 3�� ʋ�FaD� �� ̀��0��L�9�0��0��P2 �W2*�0
�0��Ve� ��W0�L��09��L�as fS2���&a3`�L�f0���&a3	�L�f4�f0���&d3	��fC0��a�a3	�L�fC0���&e3ØL��S09��&e3	��f��fS0���&e3)���f09��e3)�L�fS6d&&C2���&`s	?�����w������/��Ԥ�e~�[zF��\��0���+|_5��-x��݃�عW������LK����ٻ�a�̣�	����/�Q�x�ѷL�yw	{��6�k|�2[��M���OR=��S4�M��%cpFF��ޒw)��R�Ʋ-v�JK6n�i;�هU���eA�����m��)��kV6(�.������=���A�(�sXZ�)�'~Eʼ��X,Sܧ�X��:�׷jS���N�,�H�TU�U0�r�i���ʽ{{�Ǐ"��J�����Ɛ;W3q%QZޭ��gj�#7Ullѵ7&�ݨS����5d8��r��	���n�K �p˰v<e��������Ȟ�[R�������e͔�t�5Dƌ�B05��ݣ��oS-��!���Z�7���$�&6	�f�L�u!�����\x�$�bT��`E�����jR��(��	yQSL*����34:5\"��+V��k�F�1	:0,Do(�:�ʹ�������Ep��2[N��KN,�p�ƅ���A2���R�lTN����:��]�F�g�4�6�h|���]�Om\�Q++^hqemm]��"��3r�y��Yi��f��6����ƞ��Qͬ��Vǌ�UlL���ư@��7K�9�*����d��&)з3/4TX��[�kF�f��;��ʅ�v�U�1n��8v�i{C0�:U h:�Ĕe�p�Nl�*�![�5�vrn�Z4/ZVط{ǋ��E)�=�M�&�f[�U�z�bӘ����#%-m��t<mfcyF�m��;��M�Zö��fZL$`�ݧ{	�	/mk��	l��BiK�wLLw�*��R%R<�+/\��c�AD�k5���%) �B2ɔ�Ɔ͛"��LjI��gw�(�CBJ�*�sE�Z�ZH�3��;Ie^�o6ð�uS<@Ԃ���y��h��X��-��P��L3��s�'�m��Î�Rb�0��ո1ޱ�Xۆ�R+R��������h�dҎ��[���L�5
��i�x�f�G-�1�N�i:�fj�ok�u	��iU�B]�x0�l�g�֑.�]�K�t��jdr�M�ð�7h*���"����Էǫ�F��jA�WRz�&o�Q떚8���؍d=�چ�d]���A-/q����h����L��4!��h��2(,`��-��;̖qzb����)����X�:�#i\��b��w���C5��Ԧ�A�L��Sm���-Cte&�ф��k`�[bSU.��+0�OAM$����6a�`���;�-}p��\��h��,�ꗺ�S���x2l���7L-�m8�P)f<&�$�Q�nhx����6[8#��t�h�4BC�oSu�h�maڕ"�G�ŷ��wn�l��4j����;qY�<�n��n�zi�F���ŌBab�� �gL@�C�Rw�oC�P�6�eION+z�ӷB��
������n�b�͸4�@:�2�����ܽ����سUJF���w/B^UyɁ�-�O$Ǵ�U�e;�������P��X�������J�5�ݸr��"�pP���݂%�ݧ{�ɷ�a���!�[OX�1�`����(� PҜ�=^�SU�n[���v������\�3L5����@��MԨT��"9�r�
����Ul�P]lݫt6R��J$Y͹�.+��,�O`ѨD�Kl��x2�P���r��7�� �p�R���4�X�<�!�"����ٸ�I̩�ePa����,�f��YFYZ9�`�&�V�n�h�Y%���5m�v��H=���Z�������Ѩa��N���jF��F�������+wYJ�H
�� N�4�;�#��E8�;�@Wu��6�{�V�S6�EZt�����Mx�Ј���{�0�=�s]�g��׊[�FB��h!E����*R�X�b�ɞx����I]@��W�M$��c:��i�)�;�Iźuٙ�B���p�bh*�ܦn���V�ǀ��[�^v���+9�Tv�Q.�d"�tZmN;6�ne+������/`Fdwb�C�%�X�Y�ſ^��j�t�h�B�{�cj5x�t)���tǴ�Z�Ǐf��2n<)��63z$��*b��+�3$��-)N��dr��Rḕ�A���k*����V^f&�� �Sa��,̲�&L�G@�`�@%�j��b���TRJ��Bs�(�5c�W���'1L���nf4n�n�Վ��AD��^���ٯ*�Ų�-�^�-S�9q8a�0�0�襎��X�L��뗦�K�kt���usn܆F����f��tU�4�jS�c^m�ĝ]��q�Z,j�޴M���N�;H�Q�;L��Qk!p��.G-�a]f�{����V��Jf�#I$h�.�F��H9���o�x�Q�xJ�*)��V]�$!��Tӛ0={`�`Y�@1�rXhR8&����"���n������!��~o���6��We=LO�&�P��io�+$�����]6�Ia�����Wb�AaŃ��z��6���ϋA�g�n�Z/e��
3SM�&:������,��IYP`�'w�aǦ�3[�6��8X�iW�Ue�"%%�	Q��.�� ��7�Q^n�br�[
�� cd1x�"�o6�2�Vݭ���"��m�y�tk
v��z�o%�<�.�9P�r�ǭ
á����ܗ�]ۛ�*"-82�	u�eM��2��YAU	p��������x"n�E�ِDv��������Q"�c9�;X�v��"�5�VW�)ތs�0S&�ճkCYHc"�cxf+�N��c���Z�+v�A(VfX6^M�.X�tq
�(Б���`׃f�U_�`�e܄�v�e���OTܒ�)����Zr�*f)I̙52�n�j�C��M�yn��Ԡ�V��&UH7rd�AL͠偵���qK��n;X�.6��Up�;��ѻ衶@ :I5m���zH��j7�]�fm��v��@á	ytÃOf�l;ڱ7	*ik@�Ԛ�WK�ZD��z�laF���m�68mfmj-X_
ooPx��o`���(VƗ�v�ܩM���r���6�J�����-l��l���KH�@gƩ�՛YJE�R�T�9p�b��u�dbc�$Qut�'�Аj���-6�a��[�g��`�ɶR�*"n(�`WHTB��ܱ*�V��SgCP�v���֒H�N��24��F�^�l�YHl��4����y�������U�,�����M��5����ӽ�Ћw4kE]=1T�Q�D�(`�eHs#�F�X�^����+���h�4v�r6�7x�"lt�;V/lɋe7M^�`�cv)nlse��Xӳ�ͻT��t3f�ҷ{R�LDZ�c]��ݎBA85)I�/Ye�[���yik�+����I�AX��rƬ�7��1ܧ�()jݜY�X���]�U��n������)ùl2����TF��k4�^�P�q-ݚ����ӑ�d��Y#�̡!5r�rɎiƖ"����XƩT�f����.� ���+˻ˍc�,��b�ͫ�0T;f\� ��u����1=݈^[�ٵ6��[#�i˗�2�C��V����Ap��ɰ
z�^�f �ͻ"��1ķU'�<Un��Ea���`��=�7%,CT�T슣ME�:�I*#��c�%�v�Ժ����w��r�2��kj=O+tR��EᬐS���:��W.]w[��xIL����x�&#Y|i-\F�6:���aQ�]�-�{�3��5il��۷iQX��wm�0m1G2-7u�-�D!�wP������b�cA(�3<9D-��V"���w&i�vE0��#���[z7K�v٘X���#�ZD�t�V�Qk]�:����[����ՍZh�c�
���gHW2#�ລ�$�R��+l���`����ke	Opk�f�&i���j�0�bU"��[���B�]!�cz�eC��!���cv�lZe0áT�^���RK���RL�لkx:�vY+��O.��v3ޠ�%��A(�(�*�PP�L'^�d;mT5��]!d��an9Y�*�Ry�3v򰘥6�Z��O!�2�n����%�+'65�@Qnn�N��;nT!Z�Ot�gt3`F�Sn��-��&D%�Y�X��Q�t�ư���z<��$m��îQɊf�cV�Oc�iК$R �\�r��;R��Ez,a�)���f��X�~���Y5i��LY��/K�j�B�V�j;�v�3E8\���Ԟ�P̎���*eڀ����m�e�ry�sv�k7hi�^�3(d�U�jl�?P;��i&R��x�]elf�`�	��dx�b8�D%�����	���f��<��J5*nfS�m�!��Y0�r�Ƭ�~�w�8mT%��֛�Ӌ���&�[�ma���eM�Z�3!&��)�K���������ָ���#&���Ǫ��Jކ���(eiA��4�pTn*�eRB��7�-�v���,n^�$lią*��fګ8M�ç��
�	�3B�D(Ǒ����i5����$�ӫ�����ou;��SF��γ`��h�Μ�ug�N]2��Z-j��O8��uႲ� I��/N�4]�f*V@����m������n��X�Qv���}zz��4�:0�CV(oH��70��Gm$�8�,ݗ��+xL�u���a�L1�U�u.R˰��
Q�FVa;!�s2�*n���o�^7T��{�\�Putʶl��eI����X���]��gq���v��a,H�.�VcNR�
X�,��@�Pk8,p��=d�1�t�0W|~��Ͷ�(M�:��[�v��xm[���%����0�*͵���յ�����؛��Z4�y"r�NU
��0ц���9��FP�6���8%6��)�2�6�Ō!�yf�Ub;xn�+9��������]�K�*�zN�K���v�ZE�]��Z�;Nh<��<�ņMiv�}}I`Ŵ�]��K��F�-�
X��f�(�d]Ix${��9T�M�R��6,���ܨ����(g�DI�^\��m]EY�1���b��=x��2��gĜ>u�����&6�Ŏ䱹o=-Q�siҒ��
���,gp���á�)AV��ES��&c�5��ڲB�i�z��d��+F�]@���n��A�IZ3*�I{�!�n��E�vX6���ŻZ�-��5cؤ���崚v��t�W�t�ɘ�ץ��5h[���.ɇ [X�ujG(Yb�k��j$�pZ��LS��R.�$H�Mae��6e۵��)�u��6�ѥ����7r�ʀz�Ѭ8K.#n��Q#�*�fn�6������+�.�)f��j�#Bh#6#�v[ڼڋ,\���G/40��uu[�i7v���)���W�##`&�D�CԱ�-��i��ux+#��m����Sj�L���Ɲ�����2"��7�-+J�j:ZR2�#-^��r��ٖ��pZ�������Z`�(�ڻ5�Ncݠ�D�$lƥ�=z&nC3���;��hڂ��F�N,��1��؈[լ�ͥ@���^ilsZ��{�*\��r��(�b��Ba�M���VM���XѫP'K�GD�dr�v�a��QL�x�,fV�K3H���fTcU�����d��,;P!4�Q<T���г�e�l��o�ݮE�|v�d��Ǜ8����òS�æ-仼F�S��Y���KC�������9�%Cu�
�L���^�@�˚-�WnL��b�m�y�y��le47u]ũ�N<l�d�n���y�q� MVW��$+S�sV�X�5��G�����G�]0�+�����i&mXB�2
r��Ȍ�D�2ɒ���	X�!Lt#����M����o���,6�4����<AӖ6%����0�lO +̢�����7�F�Jm�S]e�l���>�8k�=����ڮ��i�7���ǃF�e4��b���Z���bV5Me�[z4��m��V��zq:rb��ܬ{�o���, rź��(�l7���&�<,��ts� ��Ŗ���Jۢ�,���]6��$�"�����=�IK
ך��f[\
���1���R�=�3u]�*n-JݥV��Hv`5o��q�JU�݁�8��8�Ee���Z���_^��I�IH����c9��2ہCݗ�&V3D46���XY{#�KSELc;2�p�wI��A�IyotfI`9@V3wL`^+��kQ�J�����5z�׶0�76�"�SD �L� �sr�D��T�w6^ֶ�"L�/��yD�"GD�9&���62��^�$�2M����|$[�5ip8b�Kj�kT����3	�0��k9n� 2��d
�Y[#0�;9I5�w���(9��PڽcX��5��Y��rQ T>h�%E�(|���AU	������-8�*��tG���(Q7�����Cd���C	�阸2Lg�c:D@X���+$�궸oTβ��7Ghe��[�6��}_](&h0a��L�ƁX����ʚ�X��o%[,6�"I2��$�eϺ2O���(�Aa ��یq�$��)v����<�.�Z���#K.��k7&���xK=�p�4����V���������w!�S/Iq�=�B��3�i�E"0�*	g��6L�w2Ed �AX�Ι��L���2=lz���e�D����D��&�T$d�rzAeȼT���=&�S���z�\�h�u8��qDid<E�K0ipV�`읮��d��K��K_�cߞ�o��og���G�B��K0n��7�R_��]�WT=N()�&-���Agam^�q����P�oX�:눺�p�jM�L}��g64�hX�ϴ$�96N�H�s�fƭV�9ܝڸ��Q�I���,!��Ff��E���E�7�K�OaL��܊�f`YZ�h=�n�T�՟w`%�;�%y6Z��yr����v��{۴U2X`�R�E'����dm:k��h��F��3RF����U#���jCN!ϟU��f�b�{��^�x�w.�l�*-�|"��|�\���2�[ܧHl�{3QR���ݵ'�5���5#�V�eݾq�8���I�e�,��ۛ+C	㿲�3sk��Mwl�lP�6^]*�pV:��sf��K(p9���^��-�GU,���#�te!&�M��kw`p�v*���ӸeA}ǫB9ֲdq��[�-��頨�2ܸ�ǵ=U���6
��eEgG)Ֆ�ٱ][(�sqH���k(�7I��������Q�k6mx���!{_S���P~w��!e6f��%��c��y�u�4���%�a�K����|�}˛��rZ, Q����t��u��mj06W�������PJ��������Q�d�1^��M�1\:;��l��In�������d��3�Q}�M�X|A}l���!�tTY��_^����@�z��=Ot�����2W ���Z�Q>J<"�z�ܱ�������0>T�ɚE-��"��)� ��M?)�^�[��MJpɣE�-�p�t�a�+y�����:Y�6ef$��Z����W���M�����e�]E�nYv��d�#����q��
�ԝ���9��o���d�k��lk@͈Q{36ö��1�<��I˖x2��,�]q`�m�,"�u������9�yfkY)ۅYl@��\4���=�cMe�tC6����������d���F��F�}yl�]K�k�΀�y�+�"�a_ZV�����'@ª{+�д�g�OL�&�PλW�{�o�E:�a��R�s�t�v�H�1��m.-gk�H��j�B ��["����;���UoIR�I{A��+�V�n#ڃ޸��s�5��yw�eg�K]�yٷu&Ң���n^����O��*���`�,nTD��W#�FC�{��@sz$�U�|�s�������k����y|u2I
f���C�I�Q�p�����;�n�MN�X:$,@���h2�L �-��qWjoT���*�=�f�^�:��0ٶ�Iֽ�0_<�N�d��bq,*�Nȴ_c����p6_x�ޭM��5���ɔ~a]�u՜]j��:�S!�+h[��\�̵ۛ�Pg3c���_�����޽�:����u�n�(��	�{��F��qw
�A�Y�𧎄t����B�=7zm�V��qBn�˩(FƖ` ��w��[��ܕ�q�Cz�X�����to�k�/���P"�jVl��GT#��K�G�K^Cz�Ѡ�IEɻ�Z2�n���؍�ܥX��Дk���q�WWd�ެ�@�W3�� �c5��0���%���\�+���z+�f�ɖq�sJ�����s�'WSᮦtc-`���V��굘eŠ:O��2��u���p�,���_:]�Qٛ�c����B�m%g�ټ���SL'E2��YêO6Sd0P:��9�,,̭������+�(���&d��e:�5��m���X����v$�b��0���P꫄v#]���e�������
�㥖��\��e���!Ե�Q��D�n�(�2f�%W�dT���2-L�}:h��1��2-�1��,�ǝ$,�1sU+�H:@���y8�fn.�\��ٸ��sα�P�Vַx�<�7�R��u(Pz3#�meEN��ڀ�'o�7�P�Io\�q�6��v5�OdZW8B'�[B��&��b��"�k�(��u�|.��豸k/i�h�-��!3S�(�bd�����T��{�ʾ�L���\#^s���qQK�ͻ���l�����ǉ��Q��\[m����I���+
'Gv�s�Qe���w|LΥ�V�gZ� z�ta���_d���1�R�T��΁ͭN��첝3��6��x�s�t���G�������(oU��A��ymm���`JʨL�չ2W4��2	G�)@U�Ź1�|[�s�e�"�L��t�m-�3u9\p�ƆS̛;�*wX"u�V/6�{�X$ïP�ں��*[ї��(Y�!*����5d�U���S��mئpe���273�ī�Z��fP��V�]�n.ioF���0fK�v�cL~'kC*�.�����-�2\Դo��v�c�{�n�P�\{����#Y8M��I7o2�;c$�G��O������F!o���s"���M��/�D9�J��/&=�X��cr�L|O�y�f����ވ�e'M�P��N	�"�Ե�,ޮ˼�MY��`����\Tʩ�ʳg+h���en�C�*0�Aa��~geل�Y�B��8׆]Ƅ�A���@4��:qh����y�5V�銵�N��F ���3�ʡ��4m���uZ�v71�o%s�L����؁����m�N;+���)N�Q47��q
(A}W`ו:}�_}�s,kO�[M1�j}ض#����d��`��Q�|#��Y�`���.&HYI
���/t���䨅�%��ڗ�m�p�[Y�ԲV-��
�) 7Am��]>�gu�����YDT׼h�z��xh�F����t��%N�gM^j��L��Vz#9^��}p��k�4�M�R"��hpW3H���b��Gl8 �#�8�����t�K/��ۙQF����ă=LY��'1ᯭ���ݡ�E󷯥�����rv|�k�~zG�ʿ�,�^T-ޡ�����17�hf%D�r��E���p:ŀow]w���`�6ѩ����~� E�:Ώ1,���-1�w�^&wM��5١�l���r�K���X��#��3��mv���������*Z��"�.����S��U�ckPOeѬM��3'�)1�P�$�;n]�u�|t���B�66��8bs�zQXh,��O#g���*gz��0vf6w�J���@3p�o���)ݜػ%�F���blk�����Y����
�R�����D�wXt��U��[�M,-X�(�bLT�÷כ��U�	�^@�����(�t��tۃ�7�˵���V �X����<��ݱ��O����rEM�E�r)ҶK��}}��1��]*0�8���b59a�E6�f�|/j���2�wj+������<ی�nಂ�N�������,)�/����֙-��.i�T�Tn�	�M�" ��7pK�Z�bԂv�G24��G��=��]+d��:fZ���eTs6���f%&� I+���E���hm�<�'�E��un�d����O�Լ}�fT�}�j��`Е�t����Ŭe��ԗc���|d��	�wr�4pL�35d��7�JZ���+/���s�Ojw�C@�Àm���!���lΖ����5&�L��d}�sS����@V������,	�:՜�J������Bd��e��)q��7R$��M�*%��s8W�*ua�PQPf���6�b���m
�)�uw�i�F^.qdYړ��E;�H���3�;(ݭ�H�݊�RF�����Y1�o�K���������>)0N2<E��Z6�v�tMA�Wf��e֮1-�bmI�� �'^8�{�=̠;og�n�X#��O���ӒX��=n�v���]����P'�x6���Y1��7�]�p�>���`؀�#��l����͔l�/6赖�a:�{��\]�ob��|��[���Tũ�Y�m��}ϩc�Џ\}3S�	������7��U�z����xWV���׶�x�a�#,T����Z��P&@���v�l؁R�CZn�]��x�À+#:(#����,
s�n��"�빩�ć(��w���_�^k&���V�8�+Yk�[��M�\��/�e�����:���8mfn-��y�]e�����A��B�V���pIS���,1�r�n�B���ʝ2��	��mk�V��pX�_t��i�$�H�h�ۀ�khd˜:��g|���vJ���10�A��]r<�B�t���N3�9˔��Z�GC�:2f��E���u�Jx`��l��+ɏ5��OV�:�t��]>d8:}�7T�թ�n�[O8�u����
e�԰^�GJ��:�wj�rk[��={�ib� 5Y�ʴ}��]��|�SY4�4�>����\o9���T���!Q��噃:Ԥi�[�7$�{Kc�r��<Y�J�E��!fǳ����(j%�֛��)c�0��:����Y����t��4�iv[����Bh�r���IQ���<�V6믵v<�,��굺�=�U��@��V�������i���YE�V޽C&�T�
:A��]p���c��_.��ǂ�+����%t�/7�ea�4kjrd;�`�S�k5=�On�
�����Y���
B��ZHG���@�u`<砖V�Y���sJ��.=�5{�oYq'���^��p���}��WSp��鉛�Q�Q��E�h��_uh��s��NY�zWP��:��ﮮ༳@us��C��Q��9�Th>l]q�9Y1077���ap��4n�j+B��|.��keiu�Ԭ�QOz����_�I�P
�����C Z�)$viPQ�Q�2�+YY�aEi��r�p'��j��v(Z\4��`V��֍�w��G��peCD B�IQY���)�pق�ڶP-����v@-�SXo���7�Hִ'�e�s-����ÅoVkZ:R�[�<�NtV1\MN�q��_GB�ۼf�]_6A���F�6���r�����Ӕ�9�Ȑ)�}�0���ILy�f��+7��w#������ӓFkb�Su��{�-��؋�{�!-&�u�%��M��Y�\�kf�b�j��.
�4�GDl�����H�ܢ��vS����9��Gx�m����e��e^��V!J�w�wR�+�6������pW�k�Aa�j�0�$�e�� ��#)�{�lge碧E��b��CH���RZe&�D�N9��e.�tDA�sj��Y�x����
W�xBeM��+��ek�+ Rn�.����ݭyPf�^�0�v�����q����_d��%�� ��md�����	��}��N�k���.��z-�~�;���!��ou�iEN��_�6lm�\���kKk2��j k���oԕ��Ӻ�MtE�=��0_'�q�KSB��ݱǂ�M:h'��Ut�S��$�*Zu��t�f��F���e�ٕoz� �� U��d�R��&��<���Z��S�X�8�Щ��X�U�2� ���m@������0ZCyN�c�+`�=Y��ۍ;��mq�r�V��>�ܾn��+�!_�0R�8�w�V$�b��Q8��PY{�M|E�Ԣ;zS���×�q뉑�C�-���]O���k͘x�+l`�C8��n��Б�VX'p�"���: ����
C�L�uɯ�+U=De췳7Ûi�ԣ���xË���ͭ�O�*�*�^��ĿTmtx�-�'Fl�бXfj�[��ԁ��<D�=	ɌY�7s���8Tom,�G�-�X�"�P�6f�v�pR�R&pT�1'����Y(ue-Q5�e�͇��u9GE)}�rC:�Z�����{4�������i�6�݇�gzi*P�ٍ�/u�5�X1"�38���Bf�4ⷮ���t��]�!6��̽�s��W��X���fh�J!�;4���f��do)Z�5��2g�˧]��z��'�z��d�c�w6�W@���w�J�g]E���;�9C�A�
ފ�wf�3KqP.����Sn'�m��Z}{��ki��utq�~G�z�-k`j�r�]�Ɇ����w �϶����A;��O�ז���m���
���x'��Y��/�5�z�#:��(�Oe˽��]�:�����tK�N��V���c(<8VX��Q����i�4�V�l��e�-_:$M�ݮ����982�vt�z���"wF��A�]t�i-5}���#���E�)���V�Kpi�d�E֩Lx;U�ż�΄�X�`޶��%�Z���xJ;]��IÂ����
��nGI�̎T��TF��:�קV�Ǡ�'N��#��+�k�����u����V��Y*8d�QUy��F&��,��B�!S"�M���f�t�Hp3D�@$��5�[�b�f洫{'&��z�"d��Bo,�ؕ�It&�z+5�*c�Q����3e�,�k�:5blX�gk�lm8����A[���J�6�b�3�T�� r����m8�,�=G�$�݃�8�+�[Oq��|�������Cԅ'Wr��� ��߳���y)^��9�.� ��W���#���'w��o<��C�!�P{��}O]��9|��� vޤ�F��L���|���@_^d�z��������e4��磞�=B��|�Ї�0��tw�	��<�����<�[����9��Α��!�;��c��=A�� E�������PU<��_����)�/�=~_�����?��~Fw�_��4�~?����^�Suo�.��T��M�_{Է��Q�2�Y�jNV�|�멽�}�ګ�P��'`Si�A7�ڦn:�vm�Y��'��sި}��YC(o93aY&&q��D	�����eT�v���t׼�-�97sÃ���g]>:zbk�y��X�U똖�b__h�b����q2�:��q� �a̺�"sI2���׮��P2�{�ݡd�}�f�I��e���+5Ԕ�8�ҡ��eB#�φ�x3�AI�G�&��m�ѵ��a��!)�D��t���u�dǣ!]wΏd;�WX\��Pn��H�P�ɥ��K�*���o5Ϊ�[N���.i��sp���D���n�
�4�Uf�Ϲ��V��t�c�w1��3!�6���In+{~K��0��������NۇY��rEN��Q�As�.��k}�R��r��|��h��G���z���^�/��1�M���Cn�6yIm^��hC=|wit�~�2E�,�1�ۡv� ��ݨ^�.�=��.�A���㡹�]�v��A�nE�P���'��u/,��jQHt�������p�Fc;b������O7*��a��&��V����ԃu`�*��x'��:�b?^!�yڵ9Ju���k\~�`ۚ���>`=�4`9F2���}�hvr�U�*x;���7j& Ȅ��tS8�q�V�v0�͙�ȩ�eq�FWaX�ޝ�����������g��g�<x���ǃǏ<x���ǌ��Ǐ<x�x��>�<x��x��Ƿ�<x���ǏO<x���Ǐ>�<x���Ǐ������z}�x����ǌ��Ǐ<x��x��Ǐ<x����Ǐ3ǏǏ���ǏO<x���Ǐ>�<x���Ǐ<}<x���Ǐ<�����w������>�4z%9�u3Ǵ"�i�R�9cia�`�y#bJy�1��v3�kU{zx`�W�����e�����B{�;-�����K�ƹ�����>�1�v����Ñ�ᖍ���'5��X�e��6��op�)x�ڃ �v�q
k!L�&=�ں��h�(�g�M���j�L���'6�����L(m�.q�;꺳��k�74�q���+/��;����C�����Kq���	Xo3�6C.���A�nrE[ b�	��;�����aKv��������Y�2�3[� T�#
��$�ƅ��٣9��t��t����A¥�,ʸ�b��}���ܺ��wHGچ�s�)�ju�a�Xe�ڰw��H�[�*Ik�H/vv�Q]x�j]^Rړ^�j�d�]���X��I�{x�����C��^lf���ZIa������#uJN,���se)Z٢&��E	y�ۗ8a��1<z�C��30���D�E�qs�+�1̠�F(R�+�[O���@v��d��w[��8V� �p�TT*kiݛu"�{��R@=���K��uв2(����G�w=�_a4r�ZZ�J�Uh��ҬGV�q�{�Ĵ~�Tj�c�[Q���&=ۈ�뜚h�O;1��!h���)^��+�ԝ��<����Ǐ��Ǐ>�<x���Ǐ=�x����Ǐ��Ǐ<~<x�<x��Ǐ��<x��Ǐ��Ǐ<x����x��Ǐ<~>ߌ�~?�Ǐ?<sǏ<x����ǧ�<x����Ǐo<x���Ǐ>�<g�<x���ǃǏ<x��Ǐ�<x��Ǐ<x��Ǐ0����+�����r��2mq{O��R���ДZgc�)���=;Y딸�8o��+xT@�p�x����&h⥍gk�:�U��s��:���ji{5Y\�su��wRv֎�~�iN]t)l��zb��;����9���$��0��׸����p��+�[8r�E۝0��R���T��>�Ok��C_"c�3���Ļ�w��8���O�.�ϓ:[�w]�VWX梤�.6�����jE( ��+��x���`���\Y��6�^nV-�Dc=e���א�9u[�7�2��,�mڭ���Kz���Ȍ%g4��O7��Q3]�R�W��6۪��.�`����Y�ww�]���HءTd:�����H�6�p�
%e*�خj��n��f�1b�L�--�j�ٍ�]7 ��n�Z;M��M��Y�2�d�DF�ʝ�@�c��89Z�iL�@��Q��͔�j�'��!�{����C�/�ޕ�t:6��oV<(s5�ެ	l���V�|���2�X�z��<�ډ�m=�O��^s��W��'�)��*�7�\eV�)ۃ�U��;�4���������*�͋N�qU��[[�}2f��A�^�>�X#��p<�=�1�
�0Ć^��!ν�yO�`$�1T�v����{��Ly�mc�6��7=�R4�ڛ����3C�i�7"-�V�'�h΄��8��P�Vr�ʾf��"�	J8�T$Q�"�$���A0I�+um
ť�Uv"����B�W����%�������l܄�V�d��
��@P���}bn@�s+�g-�����uG��X�!fH�&�n=�7c��O��j�%�$��i��@�|@���+V$�3i��|��,�C\���:�S�r��.,tWuޅR�c�&���+��-�m�;�4DJѷ���8	��"wK[�ד_m�hi����9pX0��{*Ru��e[��)SU��ԙ3gG9�~޵��l3�7��+�x�\��ݳ�5��K:Xwd���9���0G�=w� !V̸��\K��Ŋ����P��KҤylMy+����.�8�c��gH8Qo��qL�T,�E���t��dY�)�6�x>�gn{�ܹqq��w;����t�*�O�R�@�rn�PG�dЎ�X�����5�Ze����]�.իBj�d��Vft���r������5x�5�zQ�D�M��"�u��.r[v�6��
���n����'�Y�a�)�Ֆn��+���n��,*�m�B!2g3g�K��魾�yw|6�q�p=���gP��p��㔅�9繥E��Q��wTs���L��6�m�6��!��5a�zrc�ʸk7:������{j�� P��r|:��T��7R��Ep�ՎsZ7SZ�ͬS����%�r�T3�D#[��:�M۝�."$|�v�@������c/�&��R���Ns�\*K%V��uB��{��w�Ɯ���R���ىQb�+B�[ߎIcX����ǃ�A��o��ʹEB_,�ަ8T��k��xB��NK"���g�d���<ڃ�.RVox<��y��IWZ u��oVK=�>��##�H�ЅY��Χ��-v�����D!����)�u>�N\/��Wh�j��o��:����%+�3u
a�W��O���5����V%�&t�F��gVV(�<�2�|R�c�:�����Uc)1�z�%>_t������f�4~�+�k�72�3ȷ��]�|�؃���7v6�Dp��_��cw؀�����[䷺�y����j�-t%e 7n�x��H<'�Ӱ�@
��i|{���ʈ�ku:�Z��Cw���nf�����M�.Vc�32�2}l�����#@�oygJv)��,�����Y�Sl�v>���q�����"�����[�����mv�z,���)G�#nRή6E�Lg%�����t&�m�@�<��M��v.�m���d���el1�?p���/LSe��
[0��l�k��m�/�G5�c�Wor� `!Z�7�f��K ��R{�,�|1R��jjw�p`Ll;�;	�۽+]\ė65��щ_*y�oFD��/e�ܨO$M욲��R�Qzf����&�]q"����]�#O�]��J�f�/n,�L�5����Muv�f�n�F^�Y�ӌY�y�u\���a؜���sۛ����{�
�P�zz.@V�zLCU�V����C{6�͌�Hi�EN��9T��X��S.�f'��@�**�
E������ܨ#C)#��ڙ���}���;���PĒ��"��%YV�:�H���ܢ��A;�:��ͮ;�^uI!]5��;�:���F��FtVLA�D�$z�u��J��y�QL�K
�}\`�af�m�ﮘ56���m2^�Zɯ�m�p_q�9��i�NU�/��ʋd�FS[���Q(o�=,Yɗ>��`�� 喷|%gwb��e:��)Ȳ�Y��ha�z彿)�l�>ɝn��,qҸ��3���yY5�K�8	�h�"�*P;�P�_�j2�UU9M����	/0SD�?<Ie����m�9ܯ����Ug>�1�#\��n��f�����w��}��� |��l)շ�@�X�n؍�6\��G��wLp�:�.���� ������,�q�v�����U�ٹ<�ժ��U
�X�^^Rnh�y&�s"�R��m��(�S��Ot�=&�)����꾢�ݕ�7V��;��K��K*H[5�hS��P��5�<�թ��eh8��t��C+�d�c�T�ܯy�t�C���sJ��S����
���@1�:ȼM�6m�AfV*Y��-�Ӣ�������x��ĺ���R�H�3��{�F��}�XM�un�ݻ���W�����ػs5ov�B��P)�;7f����=XvACM�doF��$c�)�z�qu�ɝ�ag�(�$�4-968pmD��k���˽�q�v�M���0���5�,�X�Dk����݄������s�-�`T{���q^�q�lĭ�È
ʛ֮V���]*�\�z��T�8 
$.8�j֝�	�ӹY����1L��E�w�-�Gv@�u�5rX�&�bq5Je*ĩ;kA�9݉�K�-��776�v1&�nʺS/	p�̛Nm8���]I�@Z3��{�'��D�x�eZ�&�W
7-�eC��`̀�y�6)Er��&1�\�H��5Ü-��E?�a�嗐�Ju;ڐ�<ݨg�ܢzC��U��ζ7�.͎��]x#l)�����-���>�_�|�t��K�/,�=K h����=��h�^��簤6��T�7	�)��ʣ��W]��2�k.ԹݚM��xʅf��ۤ���2Xն4�κ�m�i��s1_i6.i��v��8SAJ=s����0���ҧQ5��K�ězb{&L����N�t8�YBɰgP|:�u<�����_V���`��zś�gR��v��\��H�ϲ	�']���o��1���`+��ACq�&����My�gv^�p7"�2�I�Kƨ򧽀�����ǿ��IyX�T��L�}^�sr�fE$��5ZY���2���;F�L�1������2[�Ar��&�v��:�"ur�4�xq�U��[\�6��W���]��#��!��Ia��5�޳��+Ew�ph8�s�C���W����{u�P���y؈����;UU���BL�d��Dbnjf�q�B�:��mcAf��XC�:�v(�[}�Lx��n���;�����%� O#���M������F]<���7 �<�[��i"�m��r�h�T3.9ݭp0�ޚ��+�Όc]�F�=:\8�� �E6��H��c�Z�����Q(�򹲞,����u:���Wv�X:����4�os�٤̥��Xn�9�nu�����F�n��"}+J�1��ы���,E��)8!�Q�q7�zi�K7wBa$��l�2����'��wZJ�NLly���2��0��橾�4�_Hx:��҆;�p���{e-�ykq�-��@�7�]��(�'��ӏ<+�r����gS��|]c�M�����}a�y�[]b�x���[,�0>�3�Ī�僅�]�,���	�h�v���d7W����:�X���:�cL�wm��T#r �][�v����i
�b�#�s	��d;���܂� W��*�-^X��Ӱ,��M\��]�B���C���]m�х	�����*�_鷮!�����[�3�I�;zm��]��z�10]�gK��i�J��p�1e\��5F�w���]/�c߻:n���;�*Ӊ�+�.�MWҴ����̬b��aS�q`K��	�g9��p�m��B�r��čJ��\;�X�:���a��B�H����,�6y����B�ԭ�n�u��l���bb9��f 9�s5��ub(�� �$WX�2�R@洶k�wۙ�pܙ_c�= ��$6Q�W+�0�L��S�u�w�p��P ���*�yT1��Vd�X��B��[�f"��6�2f���Wj����[��qB��|��|s+0�L�?ksU:�}K�-��aˍWT����P'�	�w7��CD��CJ}o���]c��u�"j�wڙe�x^<Gv�8,��{���SJ��d�>:k!t����5�g۲u�<�ˆ���ZG�� ����eq�]t�jӊ�n���tGeu��ѧ-1�~���׫���g_
���|dne��Ag6��jj���%+(����v�;3|�9�wnffjٟk4*Y%�q��GnF	��kU�/V�e=%=0*琱��ڻ������9Ӊt�egr�X
�@%���v�JQ�w�1�!�ė9���7���u�B��'g����72a��U}a�k���Aأ�������kMU�g�՜�]�qP���Q��h��j#��P��s
�\S)��1��{/3I5�.����z����QR}»[�t���(܊��Kve�S���4��P�X����:�V�UXkWZ�<֫ S(vʱ�7>�:�IO��z ������Q_+�����������֞�e��ٍڨ��.��w�:��[�x��b���j﷠�PJ�(8��lU�Z�kKѢ��]̼���0 "��.�F����cq�	ܞ�]����Q��7���N����oe�l���h�Wb�6y�b�{Z���[*U�f����$�qD>���צ��6�k��eoPG�w_��Uu���e{�^�	���46Xه.v�R���l�����(-����(F�=,t���a[h�ݢ��o_�Ѐ�!�|�t.����ŋ��n�k��"�T���~�ETW�4W�w���������'���_�=�~Ґ Q�rc"HB`�M6
`�6$MC.`�6�ABB�䀨�0�XH�$�l�T)I#�T
���CT���4% ��"J4HB?'!q�&��CDA��0�$���0P���:�L@Y���>���E����:�C����u�dЛ��3evqZ�����q��I�cZ�i�;,ǝ('u� Z��c\��3��{�qe"�`A�oU�[oI��`��Ҏ�G�U�ԫ�c��V"T���ZW���}�J�[��Z-���ی'�I����KɁ�r�ogU���Ӽ%��!�+��D5���9ECc`�Ih Ҳ5�.Ut2������}��9�q^�7�H�h��oьj��y���q���2�&�D�s�v��k�Բ���ԋj����:��ձu<�_T�Y�r,x�	\rt��$¾X�fS᣹2���,s���b��i����x�Yy��򝰫Ъډ�R�����)���Y���w��{7{�x�W|�g;
��H�:E-#���J�O��@�N�e�)4�V����sq�Ջ�:hN���sv�.^q�:���Y�|�9��u`�L���l��TO` 漖�fe�����(���Sj��EvO�U�$yH!j��V�j\��6��@����W�m�˚��ÉX��zT�E��wwpFԹ.Ǘ��*�"=y���@�ݾ����e7��c:k�oY���I�u����f��
��=�Y���*J/mV��\V��Gy{�7Ď���k������q����2đ��L����l�PPH�E�Q���I��2%$�i��P��E�blaI�e�RT�eơE������?�4�rD�[D�X_���B�L��A҈!Q(Km�[0J��e6SP85@�dԐ� R&�q&G,�L��&4������ B�M�1UH6[�S��e��M�ڂ LP��h�4��(K ��I�Q0A!�#(�Xi6DFi�M�E�$�RB��7�abR��h���"��`�������*jb*�񢤉��c�&"h�i���}�~>?������~<xϜ" ����n�4T�STDMDUDM5Q�4�
b����g<x�������~?��ǌ�9���F��(���SQf*:j�mE�M�m:��ASMC�M-MWQ�)���j��"�	����U%����mQ1Dն$���&��b
"��`�IUݘ&b
f������S$Z4Ej��"����(�tD�1$F�QM�ƨ"b*����j*��H����������F�(�(���EMEDMTԔP�mA��AT��[�w�Eӄ�w��OQ���w�.���Em���U�FѨ�3N�F�ttΦ��n��tu�V�5�F��rE[DCFv����V���uAVgm�+b�z��:2�k��WE�U�V���-��ް���N��@�QDb�P1X��jWu�E7X��h�EX�,�?oWW]u������N$�O�!~�&�) -��6;��c��r|�9�GQ#�M�f�yW�&�f�ؼwj�z�벸�`;I���V�9%v*�4�q��]��Ő8&�m7?#G�,�Pd��,"�4��"f�	��	���_��_�fSp{.��fV^VկL��l�\i�G8ӑҤ����#�\�7���Ff���o�e̩=�r�F]�/;!�=�A�I�fMܮڼ�y���7�7��v���zK�:�ǋ��wۼ 
9�Gv��@�e�4�������.Kd<����z'���ϲ��C��9+����MD|�,{���ݵ���JA~��S������cf�g���2�vP����V��({�˽��t|�5����q�>̝�6:�6wt���1�A�؃���E�7_]�9��;�<@�֙�u�����?/z��W��5�5u�SU��w���)�Gu�>�������O�F{u�@}��ny�U�y�Ct]`D���]���z��n��½�Ja&��#?{y+��A'q�O)4����nң�`"�VI7�M;]�cX����8��Qtשo���]o;�{<�S�ƴ�:��[�=�R���a�L�	·2jk�fŹZr��,�!�s�t-���1�7�l��q5��o�s�(�:�	H����3i�jb�u?Mx+3IC���;1V�.��kTF��۽\�.d��4Nƥ�/��Ӷ_Wk�b�* �M8������=�.����k|D\X5'A��#1���W`�ʠݻ�z��X/��"�u~��;ͺ<g�T �O�K�n>��ᾆ�����C�{,z�g���h^k�Ӻ�Nk�����Y�Ǿ�ɼ��6u����� ���`�F�8��Tȱ�E{�/�Z��-�鎌�j&���$^�G��q�v��.�Uw9�5�£G�����z���G�K�C�oE��1�i �'��s��_��@��j�7@MLW?7�֝�U�í�����g����|=�r\H3-��q���^Q6�Tߏ������=��것���?y�hs��.s̛�l�97�19,zJ^2��On��U}Nu�K/y��4s����C\����swҡ�|�_	�A�Ͻ�'��y����X4���LJ]VG��0�#�}Y�+2�<{��XNx��'ULW���9L���`w���ΖR��X,9Dᝂ���O+����7m{�[�ĵ�F���ދ�Q�,��|���g��)���`��WU����(T=��$�:�!0��EdO�1�̺�8;��/���Ub����TUx
�������H|�~�1ٹ�Q�~�P@r������L�PE^�^{�=�/�6�+-����{*�{O�t6���;�����I�8�?���~�ʺ��I�}����Fg�z!<iUm��󧞧0R���]7ޫ-.5�(DU%ʧ�em�+0U�DK���~}������4��5�ش�r��}����[=�j��OM�Bi�|~�1�G]!��,R�{[]�;s��:����FĹz��ϳ^�F	��2H3�}�^h�ʌ��
)��4_t�"��|�qW=y����hw7������,wCuj�^"��n�ڮ�g�[�����,U��S���	Dn<m��e����d�kڒ�\���e3b�u��Wr�ڠ�>L�%��Lp%��l���AY8f�������a,{mh����2l��}���޺;�:�g=��!oc�"�ۍ���
U���Op���	c)u ���ѪLQ)H�n�d�d�E��YB7���u2ʙ{D30�XFz����N�#�EA�_7�׹��=6W?�J��ݒy��omܤP��u$�.���ޙj�g��G�5����&��ϋe\3����RQ�h�CA�~}Re�]2��x�nN�m�i�\�\�z�&�
�OUn����)��ݮ�g{�������h��8A����ٰI�s�Z;y�r�Z����%='��>��}oB��J���d��{���{����������G��˧o���R�����fy�2�*���k�zқ�g�JG�8S��Z�m?H_����X:;yWNe���`Gb�{e�;\/��/|�y${<�v�zOQ�1F� 5Y;L<�3`0�vw�7x������"8���A��q�A������OHg��D}h��[�����;�/p��<��@m����-��vozƪs�g��>
�W��`��i����=��w����*M�����j��+���r��!��]��k�'ǃX����p���\�A��6�g�Fy������r���ֈEI2�g�;׏{�L�r�K�����Cm�tgx7��d�4������v-��n�<x�m�7���T���u�X� ���}�bSak=���|�GU�S�;����zs�C��V��Y�-����ʝ~��J���,�ȯ������\z��#��0,�ݠ�'OtTWG���"�x�gb�*Sޮ�;�ᇋ�=q���IE���|=��9�F�h������#®@:��f�}�6���w���=P�c3�Lԟ������;�h{��&�z�8�|�Osp�k�n�r����h������������FO��/yS�)�9��]L��Q�z]��2+~�̊`�'n��ι�D��s\�Ü��N\Ȇ�l�!��o\qws�}B��,�p}r��L�<��޿��z���3O臲�܃旾�?OOE���5I�]~���Y�7�ش,��N����^�D��ͯi��lv�:�#���c��\��tO��B�z��7�����w�fx��a��[QܐI�fQнV���A
��I�"���B�;F��7���\Ľ}���6���t�QN�Ǘ[���O�Ҳ�Q}��� �7zk@��ކ�U��h�
yK���a⯲S�&M��޲kg�&��{�/�ڷ!��Opn���To�kd�l+��I�ʨ��QNݧ=�7�͚�<���5�H��$���.�������0��DY��[��oiʞ�s}�*A�;��`��^9�E{�U7ly��8o@q�<�*�g�>���U��S�Ǿ����뭾�4k�m\��-P=�'���]��/�x�����cix�3~~����a��s>��ς���<�an*����ttn��A�o3l���o-�V��nݯ�V ��Bᜎ�m5���U]�tK��@3���m�\<7�!���&�z���7^�:�Ο?�hZ�H���̷�ew�ߴLG�v5�u��υe�:H��t���=�Ɵ����n��?8���"ga��ؚZ_LD��bo���۷��	�4��)�ʎK�J )3��;w9�d����aЭ��[Am�Ӹz�4��i֎���a�QѮ��W}7�����9r�����3�d���ʎ�+��F�4�ESj�R5��$a��4�M��wfE*�nD�b��і�.����r+�۬q8�e�E��᫮�J]Vo���:=°�$��f�6<��̖�5&�A�9}|,���o�K�y�y�����>�m14�:ط�Vz	2I�0h��7S���/��f�ݙ��q7�x=C�����Z%��qW@ʇ>�F���Y3����ϼ�vV���������ި=��2��;����ڹXg�60�Iu=�JT,�0�,
͓WŠW}2t���s�F���sx]����{��E͟OW�e��Sw*u�j���?=�����.��{GK_��o���>�t)u�Oh�և��o<��ݓ�,�{�y{��_�0�W^ޝ��4fm0���� ���3�a��-��S���Iw��ݢ�/\^���V�G��f���;�^�u/�&�Ә������_}�?����]v]��?x�����&��|jLf:�jmX�/&ó^���*����;�;a�m���u+"[}3��#����N�!8�5j+���`m�Z�z+�;#֪���{0��:e<�i�y�s:Q-fvj��'{��L�S���EAF�Dyv���B8���}c6#�ys�Ӧ>3:�t�(�ͫ�_Y�-ܙ�wDyV��d�Y]�$���G��2�9s*H2*�,����[�������>=�	�r�����f���4�t}��=k��OO����Ul�b���*��w"�C?u+�0�1�UQ5;C3;	�+��o:���=/�����%���Vyj��K��Ré�}�2]����f�i�h��B�y���K�qz�=��Vc�<tM<=TX�j��6\�ӵU��I]Ӆnfd^�p7�dh�.��9W#f��o[4�;Ťh��.�Kޝi�����%P2ۄV��w�W�&��3��m[�Qܼ-˵�o%o�_���lR��	�'��5���z��ͬ,	֎$k�F�9.�{z-�亣�=-Ï�l7�1s����� �����#o�=[<b��c0�!b5����&%޴�;J2�Ƭ1�f�=^Z%6s<�c�C�Vŧ�Iyѕی6�[�
nK�d��#��]Q�Q=i����Sfᬋ9!�oS�6���	���o8[t(q\6�soY�BbYh�kNck���e���4�<��Q)P���`䡪���Y	��]����UOF+����z�&ܼ��G���.pl�xj����*`z�<.:�ą�e�˫���o���^n�u0�[;�6zB�� k�ڵ�\����󀍺���^�\m���� _Յ�N��(k V.�/��Һ/����U���|ӻnw	r�τe���-�[��r���U`���� �2wfo��cnĹ�����9�PW}䳢��IW�y���}�Cy�B.�u�g���YO(�`(`�ej��^cr�GV��Wuu�<2𵞒�{��x�ʯ���,��g�S��>�o�s}�\2�ŕ��?�C�Ngf�z㈧2A�|�gb�����D���P���7f�Z�7Q{w���^cEo�h�=�*��;�vY����y���ȯ3�ҹ��[�3~�[��������f�OG{Z�F�4���ϼ�D��|��~�Sy�yT�e�Y1����$�6d��쫒snwP��c�ɮ�V �)�{5��M'�7c3�]����\����L�K�[�p���be�Pfsz����9jr����wa��#�{u���M܃��E�e_V���o��]1z[!��N��:�k�(�wL�J��ں���y"�&��Ux�[�/�|#���u��ߠ�I0Y�8���ΝC}G�嶷l�}�U��� �.@�XO��M�y��\��{]����؅�X}����Գl�/L��k���nv�����	��VN̹;��\o1�Q�W�ޒv�g�ζ���U����xl�jf��
/=���;Ӑ�u�\Z�=}�7Q�����:_dm��!��l�W��U�h�
x=]c�r.��\��sp��f�ύÑ�^�q��>�:���뢭n�X�09,�mh��w��3�ן����r��I�9g��ٟ#�].��զ������|�E��7��0Ì���ѯ>�=N��n���?/WU�SHzf�z�M���샺�4������{/jU/{�Ɏ�2��w�B���(��m��t@��6�tl3�9�_o���<<�t��C9��Vo��7���j�\���Ա[�f�R����Aw{V��Ha��Xi]N�����q[;Q�7�>�&��ݩ��Λ!�$bA�z��oD3��rq-m꘵C���q���<t&�Jƌ�--�I"P�RS�pt�7Y�����v�e̼o+��9Vw7�s��P+&�iΗic���u����IP[DCɵ��.�+d[V�볳u�Fz��:�%ǚrCgu�W}Զ$����:�C�e��84d��=�3k���c۫=����Mn�`{$��*v�;f�R#U��n�\�5D�*�8F����.�4;�蛱���)S2�8�ʑ�5�b���y#zE�`�Tf��"��ϫ:���{Q�uB[���H�n\[ZdI���~c�5FX�3�Aj�6wg��T��&nj�t�u�]&�hޅ�V�p��(Eyf����;�Nz���a{q��M�Eow��u�u�<��;�+QΛs�ӂ��[�RXČa���ؼ3υr\���<��M�CsYKqz�[`�qwl���od�t���2�����2k�k���:3�$��6ɜ4�g7��i�w�b䧗9k\��ʦ�sP,���{[�F:spI�e���E��;[]6��M�DWG�^*k�@�Tp���s�}�SՅ�bY�guu���a���}F|�8���!�^mP��zNn?��h$���k	;^{:�+���:��u�a��ٺNlY/��U��0.[��a�w���N�:Ud
��'�:x���al�~�����_Z�^�S�Q3��s������Y���;/>�EcN'�y��P��3�xy��vHi��&��Z��j��3/����.�@�B����<9����(��7�/h���i14�]q��Z����3����w@�m$��m^��S���n*ڨe`��\U	?�����bV	�/j�\v�Hw
�]�#�e��6Y�c-Шsm赣�+��r����-���Cå�[=��<#����e�e�����Z$�J�
�o���wAԆ�ܤ X�;zk�t�+<z���Մs�˔�@N�'Y�����6��gb�2h[���ϲ�(�@�y�.�	wk�� A�x1����N�����j|[6z���7]���7�s������/}sKwG����t�x��~�t6�e��XGL�\�%���������m���+$����YN�Su��[�٢��<��.�&�F�H=d\��W.�����X��'��k�V���YjB�(oN��#m�Ey�'�v��w!�y�Y<�Nɵ�%�4iՙ�]Ğ���;'n�θ�6%�Cqc0u�R&�s��1{��x�Ft�Ǹh�h,����_5|�{%e[���� �j�p_�z���<͹5໩��\�v���R�ӝus\F�S��u�����u�����WW~�����ъ5���|��
6��޺��6�mz.�
رoQ�:lTXq���].O[=��U��Fq�س�Oo�Ǐ������||||x��~X����4}��S�GS\�t�cw�&�!��u���:뮍OU՝b��-���b��h���w�vA��{~�_������~?�������$�f�b���Ѥњ���T�Dp]��a�����Wx�=ƚ
h����������b�`�*�*��kM�h��&�����E���=U�Z��4�u�񣽊��lPQV�(���
���Q��Aը��h�f)����������
"'�b*&�������ƪj+��ULEALM2TQP]mV�S=m41LS1'ͦ&��~F�
����)�����UMD��U��5MQ�ԓL�CDLn��{�"�*`�j������5TQQ�D]mDDQժ���� ���đIQEOQ�f""�������E/wQS{�D�Tz���Q�"��UG��:���(*�"��4׫{ڊ�޽�7�ҹ����ԫ9���);/����zɖ���&Y]�vئ�+e�kK�/-R��mj�
v��u{���g�u�h�;�=��Z#��.�����=~��9��3���
���ŠOL6�o���鮡�~?�Oq�w�gOfY��y��y�sC/h�֟C�m��z/���kp��L�^�é,��0[����m>�$��"\?�� ��vԿaܥ���}�)B�����?d�^�ҧ�ʅ��W%L�`�ƖN0-����u�5�����W��ߨȞ-�����+(�����9L��ڊ�� &ً�~�gk��.�+C�S���5M�hΰ#����-��վ;ǐP2pD���ߜ��Gw3AK�)�L3;��}�Ї���C"8
�w�����+��d�����=��E=���`d���~|^7D˘��ʲ����&���x���C6�z1��ሔ弹ı+��2�u�3c�:�@�KXb�*\S&�ETosa�N9��R�h�
�����q#z�$�b)9Y�"��sc�\�J�a�������ޙ}�=��Ǡ����@w����~�{<Ԟ��j�	��z������h4�k�0��,C����!�4�
��o\?g�E�2�*`�qB7�����u�f��r�k�� ݍih.���J�EM1f�O\,���Ĺf�j�1�9&�r9��3����,��&�;��7��J��^��P�8�m*Ҙ��K��aj�A��u�S]���`{Kk&�u�z�>۝�2>�"K��v��tfv�ڜ��Mgޞ�{K�ܩ�R<�[a��rz����1.��ok����ٳ�8��Q�8�"F'�b'�
���6�nƲ��ֱ��ӭU�\��]��(*"�2
�ZC�[����j�R��Ԅ3�����!����z��<�̠�$6F�Ǿ1�oVܚ�<���Ph��AA�<s��^����=������I����h;{k�ғ��a�k�#�ɊƠ_�9`(��w���*w]K%�G!��δF0�9���MGc��>Ϋv�k�v^&h�P�Pɩ(C��z��p�-t&}6�gF���a9��)��r�A�Q ��q�10��ʜh�7�竮�	��%۳�$���LZ�ml��������<8�[���qt����I �1>�5�>F2����W_�hi��R���*�VZ8�������$;�Q�`�f�?P�,���&,y�?���5���Kr���̆v�Hθ������7557�sX;  �c�c�uk=�p1���s^��̓"ZG=�M�m�udx����v��mk��}w!�8^K��P��K	m
�ۛ����N��]w�m��,��a�:56�[�����w%k�ѓ^����V���T[�L测�н�az��1�+�e�񇺎Lri�b��Ww����?+8�'��NV�9����êމ���"ܫ�6V�����0�6-���;Q��ީ59ݎ��@����~'�ƽCo�\�d��Փ�Y��9`����{��.�0��K�	������I��N[�R-B��U���ѕqqnS;���<�0au�0B�[B� cz��i�!�e;}�=�w��T�E�&⩙D3y�hS,�����E�!���
�u�_]���$/xvτZǡ�!?C�9�C.����J[�o,�4����<rco��;6�]g��摋�|2}�:O��Z/�)�s�3B<ϺKA	��fBw��j�%����2�<��s�EoYaw�Sm�hj�r��PX�[N�SïûZ�A������`���7[���R����R�(N�6=���.��-�B�O2�S�4'�}j����6��� �\��SZ9���45���Hk���&�еnd㎿1�Z�_��^���VН.��0�UF�M�)Uo\���;���`���Ά�4�|Nk��7$����3��l2�{�ӑ}p��pz����\���&�gO�#-}��_A�"\����i���uY��%��Y��N}܁���C�-�܇n�F!��~�,�(����:����\T[#����-E�_!��ݞ��m��!�FD�+��zX��}^"�S��d?q<���Mo�b�W���W�Cj��r���%y�
�S�[���T�d�k�R6��H�km)�"�]�!x��ohJ��ȴ7�Ӑ����Q87yK9���Nf�.�R�"*u��������z�ֻwqhR����|7c5���������i[.x��:��X.#��.�n��?^-f��Dx���Ľ����qM��M`a�֫��1��jz��v#�T�׌S�5F���C�z��ڄ=����{�f��sI��Q�J��L��k�t�e
6
�������Mt ��(���[�{9���g�v&�3B���g����ڨx�?�o��|��H����S�/O%�o����}�ޙ��0�G���~W�d���!�_)殄%1|�~��C�z��1��:�ϫ�қ�5B3���6s[m�E�èa���\�o7n7�ӎ:/���t�Q��S�AY���͈�}@�K$�<SM�����g��Oß�$l3czD:`��u� ������C����D�ʳE�o��œ�R��n�c__l������K03�	r�x��#Ub�5�8u�C�)ٹ�P�ƽ1���D�i;��*��E���PX��̙��7U�N��kuz���8|L z�0~ng��ݓ Ju��>���I�V���z�R^�ǌu7�n_��ҭkyt�)Aw@F��{��T�\�9r�<zͪ�i�:N���Awږ;��O��Fa쒱��4��-u���w[��Z��]+ ���^�ʳ�Vg�����2"Ls[M�t����ݦ�W=�9Ad��V��# ��=�Ə������ ��.�=<�h�w����`d0sC�Z�Bb[l��NL�Ǥ�|���1U���v�Uv�<K�|�^7���̦n��o���à<'�����0��o#/��4�W��E���F�g������O��G���v��ы�g�3?������ w�}/��&��VX�L�ӻ5�G���]!��k�p:��=%�qh��b�'D[�Xh��?�����X>����[�Q�ι({;��;�2�/EG��<5c�w��7Nmciހ	\Zĸ�-���툦�7M�V{���k��}�R��-L�pta�9�`k�ؼ�	���7��8���3M�,:�YA
F@0���
S��
y�}��B�}��mW�I�,��?��>>K���s轌`%rTͶ�b�����)�DP[����ג��}a�[�>�l�=cռ*�S��a�E�.==^UX�Rq��Ɩ���x�e1٭]v�=Yxh�P�v�`b�b�N��o��p([�z�K�Ƿx�
N�"#�����r�{��t��= @!{')5x�!�P,�`t�K"Mn�Om����� ׅ'�o��<w�}�&�x�e�M�y��Vpʽ}��z�����.ӀX�n�M7�/n�Y(l;��{�,�2��n��6�N���z�a�����͍p��`nX�^��p�[�&k$rC��zm�m���ʑQ�>^ �8��{7����*�����!�����ټ�$�<���'�b%9]Ǌ4�����_"��B��h�V��u�8�7\9C�x8�ƕ�2{|���)�y�I���> b)9X9�Q�b�on�Ɍ��z�]-�ײ��m���?׃H@��h��o�-�#�h��r!6��m�^�5¡۬�`:�(�����^�ֹu����.���-ׯ��bX`=�E�3�
5�3�G8�xe��4��ו��L;�.v:Mld��;Hz�m�e���z �s�	��qM ~ׅ��:�]�~h���T�j��kk4�q��!���|�gu�x��F�[w�J~lF	��q�
�|3^�ٷ]��������=ӨKD����{Y����8�[yX�%�:�ƲǾ=>�� sh/���!ۧa� �U�³�ֵc<(�36���53�ynd!�bxf�3p�}��I�İ�-�LW5�1�2kC�Y���
���k�{g�`����6LLp����Kv�k�vo4� Iv�ov-o��a4���}���j��ì;�@jZ~��D����FG4� $��-���`�Fm�ޘ6~��;��ӯU\[��SgI�.;}=����F�g��j�y��_M�d0���'��o��Q^��k��o̿E�l=	m񧴥� �30��$Ҽm���d�t9�{��X��p�/��}-9�n�1uyR{�n谟X�Ûz����]���׾����� ���03�� �(v}3O�����w$�V*�i�� 3�k�� ���[a��9KOղ�j`��$��tȸ�牨��[����LbA�{��P���]���f=�1jK$��gX��6�S:~iw�7�`t�	7)�.;�xN��|����OlNH��y��!?1�A9 KO�����{l���4.0A�7����1��.��ڙ���?��5����H�#��sZ��):��_�
�=��,)�T[^Rg�z�W�ׄ���:b%� �����>)�t1��-����?�q��_O��d��c� R�@�UC�g��%�l>ݾv��G��K����a+"��o@/m� �a�!��;pl��L4�R��(���7�A��sɜ��x�yƶ�ב\�8�@�t�eٲ*%�ۄp-���'�y�%�Hn��}Oxu�U�{��Zʝ���X�!��q��F��\�%�r� ,��1�H���]����N���#���3<�8���m�¨Y��V�@E�Ғƽ�i�Jxw��+Aaߺ����KU+��ώ�L�����q�[Ő��~�R(�1&���T�l�t�*�U�%=Ӂ�\���h)=6��;�*��U�s�v��z���*�x{<�5��	��,`GW�_k�)�|)��ϝ>�'�Br�R@��-!�l�]M1ƥ�������j�{u�B	RG�J�ґ�e�̊��O\�vJ�[�.b|�&����Q��[�3�9�p��������؋���X8	�L�eB`ke�
L`ۍ!�JװT��\������cFíT�����E����dt� ��lsH���צ�N�՜�a�Mc�C��/A��ת��9�X�j[��Zr�ג�.�'Z#'��~��d�Vl�k�z�ms2�B���p�E��Z�=�cX/vD�����A3.��ƺ���W���2<�S�}[3�/c�G�b���P�k�G��@��/=���"fp�eO�nu�4`0&�2w�^��ƕWq������앯bj/��cZE�"=/B���+�5曌�M�����ٝ!�(�d���%��`�P���W��Ou���}�@�κ�Y�(�TyîO�Ǫ�?dMd�|>��z`a������!�k�9���K��[������w�&O�a8��sw�-�6$<N@�{���Nk�=[�M=��b�0�q�0��� _)�O�^.izͼ��/V^<t�ֵ�x��LB*�������xOB�}�Н �N�:���p�ό�6ʙ\�'G��\E���3�������`;���b����TɓI���`f�J�Up h!K�A��H���sQG����'Edpb��#�Tfm$�rP�^�__$��
l�[�_���r�u���۲ߚ����s�=�"�w��d�Hx�.�q��W�T�N��d�L�s�1��&���!>k�H.͂e��M:�6��孢	�=�,#].�e��'y��J��U(��7E1�����r��p��qn�o2���{Y�yss!�!���F��0u�	6_ҡ�*��Y���J]*����tn����e5$r��<��������D���xN�OIij�xj]c3WQ���;����1��-��c}����n�`&��N�ÂXw���k�	�lT'h���&�H(���~{������T!�·lq{��q�*������� �ØLx>�_�;ny=2�t���ܖ~�=�☡�����,����b���ڄ�����	p0X��9��a1q�t^��P��z��K1}[���~����l�������a��9ė��ڶ+�!�����A~C�x���L05c�f�ؗ�to��=�6+Co9!��@"|OT4��!�t ��ߟ;��y}�ن"�E`�4F�������>OA�ld�g�kw���f�9:è%������X�7�,j�Kn��v6�Ø�a5�.���&:�����\n6�K�k�N��w@���&�x��2�rt�K�[#���k��3v���e����CӹrgH���fY�q49�շ;ے�/'�Z�����}����� =��ec��o=C����zכxmhg�X���B��NlMO���c:5�i�n��P���5�Xu��ݥ��6�]ӌ5�r^]a�zs����N��-�2/qp#�=UX�.�<�Cy�	�L��g���pg��[�ǥL�D����{���j�?*��(>1�C�^xrMBUl�aw��+�D�r,,�4q��4Z�D �W�E�$��)2��#���)�"J���{�y�K�l�le������!�s�NP�;_Or�n'I��Jr���Q�~vk�<��3�\|8�n`�����~�*j�H��,�ޖm�L���K0S}%�N�I˼�+Z�1ت��0��lMɐ�p��Dq�f���]���/����c��
�i�	�����R'�)�:z޳�;_!�^u�l�^��ԁ�a'�?y큿0Q��G8�C�-}��M7H�te�s��S�ǀ1�Hdix�JF7C��"	���$yaDP� ���*��=�/��KV7^�}B�ʛ���wFi�=�%?5�FM�ڹ���f�;�nl0g?0o ��{�x��L�_���bƔ oQx��)�í��s��.���v�F� ˋ�˓������q!�.���ލ¨-9�◶���}�u!�S]H�#0�g\�����d{S�F'vjon�Awb"��8��B�:�L�x�:��ޅKI�K��M�/���-�/"帕��u���ܢ�1�r��{]3U���8��U����W^k�5wXĔV�-���e��\^�``��:Lף�U��L��j��Ż�?e��\ʽ�N���6�wVIL+}��	1�"t���h��v)l=��5��H�5���`��7%�jq�/;�Z����gZ*�8}�8Gsv�׸v��e����lu]��/�"�6����0#�VY�[v�of"9+��K��mf�h��oi�M�IM��BD�������
�	���y3l��s������Zs�a���d��Β���n+�m��,jά�4�Z��i�rԎ�V��;�ǒ������+�	�(0�dڹ����Ѳ�~��ڳ�Fj>H\Vx�}[ԩR=�Mi�-J��Y�.��Z^��(=IWc�@��qy:��`nWg4���{dl�Q����v���-����1vm��w��Ң��Y��
YډK�1��8'VX��Y���S�%�h�}X��5g^p�*As�)�1�B�ȭ�Z'���A[]�ԝEt����s�R�p!6�9T=�����>��/:�%Y�	XGobJT������n8�+���}o�=S����w�dN��E'Q
����G$�������ՒT@I����˕�J=����|������f��&��lkʇB9:0��ù�]�Y�Xto�1o�.�e]ê�pͺ&��sōy��-�ݪ�v�����.���i�0e��y9K=��_ގ꺀�c�i*pi�DhӶ>�E@i�ܖ;�g��h�.�'A)�Y�̛���2�<C/@Ӎo1��-���
��ӾW#vi�D9sE��\J���t�h���u�
��iJ36����&H�y�ͷ�/o�T�֚�)��/n*��p�:�^0V�i�P̑r�v�aF-%������;��q�W���o��PG��P�yepB�n��ɂ��p�y�V���M���t��[��kHxb�;������6`�g�8��8�wCJڌ.Ro:�>�U�*Q����\�q8b�����2e��}�(�'<�b��r���k�bjtޓ@��xa���ϳf"@�N?��B�<��4�-R$R���le]M���7�K�ɜq�Yy����t&"s�O��gq;�0VbN�#��v��S
}`3�nRW����SX�W�a�]��m��Z��{���'�Q�^>�ƌ��v��}A^�AЊ��E�ɗgikR(�DY�k��&�!�ׯ�����tͧF2O05�NgQ7�R:c-&'9�����u�o(�h*b�����J �"$�(��D5v;�����ؙ�������i��h����}�_�׏���������~�h)�(h��
(��.t�j�("�������IM-4�=N� ��s��Ǐ?_�ׇ�(��h�N�)�4b"��e�E�V��9u]f��X4D��S�th��(�"�U���N��F�$�.��ՠ��#�h(5�4UT�h��QQIN�%�n�*:ɨ�ɦ٪Jb�lu�CUԖ�4k^���}@b(�B$��(� ���*�a��"+cJPVضwv������b���$���j�j:�b��;�M�5F��U���a*�
h�N��UQIu�N�{�uw�1�Mn��zɪ(��6
E�n��Z
H�}`�GY��l��=A�())��.�����j&���=��Ш�m���!E�!8#��O����u��mX2�wC�;��a;\&e����L<��G��'�$6��ջ�k���;����}�t�p�OƐ�_��2��4����!22A�$ ��D$l�Y��:��]�� ����@�p����~u����o���k���[���*Ň�X��"Y���K�>N�P�nd��c�c����zMsO��u�� lC���*ٟG4�Z�,�����o�����㺨D~Y��^ԓ��aŜm��������=4V��o��"(~�$�W��;V�&9�Ld�n�myίa�Dėg�D��F��;�;�ϝܝ��djq���H�t�4�>}Ե�ws�e9����p�|fT�4c�RF��@�x`�̄��3��k&�D�6�῕r���`����$�?�ݟ���]��YY �ܙ�m���C:���A��A��Y$5gY�b�h�ΞG=;�����+h&��s=t�j���*�B��
��o*+��O�7�ז@�4WV���{lQp��G-���޾�]����1�l�桕�9�`�~4L.z�-{��Z�B��TX�>4tWc���<���5�A�'ұ��l�|��L@����.�|�܈��_O�I2O�1�º�[W+5c6�Ž�S�܅��N�e��� ��?5���?�r��\��Y�ٚ+����W����e}��b�7J�$���?n�
98$�1쵲m;oG�4�Q�#~�ҮeS�i�巼�-�b���p�!�S/[Z�!kb���r��%\gb�}��@�!X���X��Zcu�	�d���G/�j�;Nm)�juu���W�=������ ��v��id�G,k�^1\�$��Ɓ~�/��-��#}B~�L9��5���g �Q��n����)��P�j�����"��1sH� ��=~g��� �k������j1W�G!=ӊCF�4�'z��g4�aUjw�����	Ic�e�hO�7!��<`f~Z�a#3�-sE�hPؘ=�O� +��|�<Ө�"�x6�E�,��Ut�XHOt�͜�uë@�j��s=p��e�:�>�S��Z`Lk�[&�е~s'p=��zg֪�Q���_,L_.;�C�Yxj�`���8?���lsL��0̲F����������2[�6�>���ǀڢ�v��U-ƽ̓~^�倷c�D�y�|F��V�s�:Ɨl��U0��,�P�������,9O�K�wn�'�]��`{�[9yחx:#�@�d���z���tC0d���z*b��N�=y�k�B!�Ԕ�Q3p=2�tM�1�����T��Ȓ��{f|�o������M�8�6fƴ�ȯ"���k�W!L���]6~|e޺�W��8�)��ĳ5�Q]b�w5�i�K��T=�9MJ~�cs�"�h��x�=^3��4"���%Fv��yI;�z,(�����T��Gִ��:ƸmJr�U�W8��(zZ���F�H]e�ٽA��vkue	�,#N�_�s�߿�>|�y����~�����N\�* 6N���9N�>�D3�U۟�S<x�,,1.z�i<K�I쪖ƭ�!s��� �eH�om�(2�������5^�u�6�n:k���������~P}��_��,�%6��%L?[uffT*�oxa��z	ʇWe�w�TQqQE�v�\O>C����)�=��ιJ�e�(�j�A�G1,🴙LP�
�،��(�Oџ��ju��\kG�r���b~G�E�>_�&�௩���!�p׻� �\^%� B��eK&���!>{_g��ǙT�o�UJL��P�%��遷^����@���]���E��R��n�cX�
v�0i�gD���K�Z����q��g���	{ߔ'��|z�G�&�ƅi;��eWCը��֔*��k��&�Z�����!n%�0d0�t0t��#�kt<Y=&���9B��0�n�;a��b�����g�����WPE�di	���o�D�U�G�2��G��O�xF^ϸu�c��D�^5_����\��'\�o.�����m�tY�@A[��~��GWǳ�b�l����/s+X���H�mܻI� ��Q{���\�[�e�${א��eW��L<�7��7I��h읔ב]i�\���mW+��Ksjɚ}4_}л���m�vÍ^����ڝ�L{Z��B��ȱ�k�����8"t.��ߞ���$���"�D}����yMҝL�^w"�>�i1�Q��c��z��z��O�y�(�s�	C��Wզn���^�K�n�'�*�P�n�ߥ�_dfHfɽ�_�A}��;(��L[X�c�v��J�{P�=�2���p}aC�PO��`���WӺג��y��W�D�z����(a�ʁ���si�x�Z�/���,��!4���Z}�c��G��sT�ԳI�m�؏��)��}�����ͽ����I�o�WX(~�G�ߠ6���B�.,��|�1��^�S��W��J}�*�F>��W�9�֙��l�ʖN0,v����e���o
�H�x[@���ǧ��$�U�wg�,F���R��Kϐ)	M��Pd�)��z1�����+�J��畇x���+�/�惟ML`�_L1�u���I�j�q^�Ƚ���Z�I�����{�>3�h�R��E���v̏��y/�|Ǡ�9�#�
}���}'��DJt�����H�4Q���P��֪~���\^UJ�v�6eK'1p�y��ʆm��˽},�
}}%�N�I��NW[Pv�Jz��5��zk�y����$���:�Hv�7�V����P����}/"���0α�hu��!�fq�YS�#�g�hָ�����������3#��*â*!\��G���a�Nk���2���y���P�o>N��8��v\�1��ؼ�g�w~� g�p*�8TE��9����_F���mu9�~��w*�D�h䙭�C״�\�_C�y�CE�A��f86��4��*]������0�r`���'o����]ز뱔�^����F%�at!��|�����?j�*�d�߾�hμ�k�M1^����(�Z��k~�PK�>;���f�ڇ��N40B\w���0�u�iTm�����痦D���)�Gu[]�JO�x��y�+�@UR3^�ٷ��2�O,Az�|��4��a.�K��!�?�v���"���K�1���=>��|��z~5~3(}��~�8M��߁K��Uu:�|���`^)�֜�d��l�|��I���Fi�{�@�z��i}~�����.{r��N�Zt�HiE}��M�`���T�s�`k%^ݠ��0�3u�y��oљ�f煲�vCr]��7�����R���ұ�A����L[e9��Y���u.�{�wo����z	v��d�3"�kO\�o��)�=���B1�JuK,B��6��7��<�wR��u5s��ݭe�Pq�!�)d���{ȥ�n�@�t�9��������wp��ˬ-���G����~��c2���O�t���(f�[�Lku�T��Ä�g�}J��:��*_z�:��;����[�q��ը��"���Zn�����V�Y���e��譓V�����-2q�nW0�;���������}_W�?������V4��-�qcP���/��1��&�%yQX˜����	�,�,s���8獒�	)N�=��~�[�6�Џ|9�P5�����g�t��ǟ�ܡ�X�^K��B�s��dȧg�%�p�íw~�� i���E��t:U��=
��& E�r�`����D&I��L�m��w2�T�s�A݋���BՉTS��G<�Ƕ�c�� �3�Añ�>"�]�o%bW\ſ�5�{ײ�����+k�`/1W�"��\h��.͔��m�=�C��(�,�w���m�r9�l	l�p�4�u�O8Sm��.9�\�6��vng�`��tc#AڻHh=9�
�B�"��/<�zxУ�S	�2��֮Qy�%%�-�`���&��0�fgg0�l��O��:`3�X�@���Ѯ�	�B̓q��E�,��Ut�X'ע�ҵ�F��o>����{eOn ��}n�ks_��q��zhZ��N8�z=um�Jb�ޜ�U�(���S��A���)��%܁�l|5�,�{h���Z�];N���mq�u���p���Vw�lU��6ЎiYc����D0�o]�śiM�s�|��Z�z�vT���zVٰ�:�}��/�D����;j�d���|f �x/���"������K㴬�An�Ӆ�؟9N�r��H��Oe�}_����������������j�nV��n��l�X��h̡ިx���-�W���p�
��Y�"cq����#�ήs��c�%�SL�_PΖm�-�L+�bK׸ñ�& {ߴ;/��,�)�$��y��Jto��8��'�����^��	���6���"��q�k�A!�p�hD�4��-�'I�{DaVg�I�W��5����'���x4�
� ��o�N�Y����/ ��P��9�%r�My��N�y����8#EWN[!���x!0��)�E��x�ƞ��ke��!C�ve��(�ru���t�rx����C�5���zm���Ɗ��ئt65��,��mz-��7M��3Z����q�����!�;������ s$�P�����ߏH�C�����Ё�d��3*C3#nn2���k��/ݫ�2�)��	��)̈́�0MP��v#g1Ϭtv�'�c뼆����T��w��*�T�08cϷ/�j�H�I��d�g<S��b��=��s4n�R��uC�e���ixb���D��.�}]0�U(��%��>�����>���G�__X�aK�a����)�v4�|~����Ŵd�����	�W�ղ�l��q�Kv�K��c�n<;][� ]�/�V�8�:,�hȖQ�Cu�������sTo�s�,m'���̧5��u��P���Ȼ2�.��W��W������xx?��� z�;�o���(��fo�w��:���	��n�|k�4��W���z���]���|��&�i�cV���ݳ���"Lv���s!|t��F�C�u��X�'(Xޤ�e��W]��<Ɣ�U�;�3'��,�����P�_bw���
�c�􎀎��&��ѭ�Ҿ9���	$���=���+\�%�]S�%w,�]��zC�a?�E��Z�;��|v|Z���ٕ��{�ͱ��I�é�|��}���	�;A��r��ޟ,�����h�����^a�>'�K�>ϳ$3d��E�����-��1^�lX�M�Xr��M︪�⬠`��&,/>'I�/r����w�;�mciނC���"�m�l�X#���r��k�̥�B��g�5.ldK<X4���_�Lx�՟�L�SٛCL��L��k�X�)�k�x���0�72�)0��^M���ZfP��5���`x��#�pN��(ڠ�w��s���l�cyv�V;#�G���T3e��ZUq-��/���C���ڞ���d*���3F�4�w秪�e �\v�w��n�:���͸��ѕ��]��Q�ܾ�a���HՇ�x����j�=�V.��x�d���R�p���
ߔ鹊��B�#ޘ.��.j������ }��  ?��� xNPGSZ�.�w�Yp�qCҐnm���uR�/?}���a�{Q^������)A�R�4�®�`�_r�]T.�p�#=y�����\L����ͪK�D��d!Y*���N(1�P�Ȥ��Z�I��i���!{�}����v���*��K�1��s�6C��cH"}}'����Г�x�'ˤS���M��y:�I��jX��m�j|�������0-�Д�͵1���3����'�z�$�Vvt��������k��T<b�����\Ø��}|�>�� ����kh���gK5�T�:�s-��}�����y;e�6à9E�匤�5�����Q���~A���Ӎxr��8�T���py=�B��Q{��kXMs]���BԍcA(�zO���v�lc;l�v�,�j����f�˰�]��W�D��="���i�=�%?5��޶�W>U02��n쟕ϩݰO0�c?K��^����0:O>�m~O@K��H�4-1�ù�k,{z}[bMs���N�#�>}�#��X_��Nd��)�~�Ū[Իw�m۠��)8%��a��FQI�ZV�������叮!��%b�E�Y3��zi�h��/���ʠ�dH�.ԳS������<w�J.����UJ��}��V6$D��r��	��s�\2�/F�X#J��VJ�Z���[���b�$Ў�e�\����\�s湺��=��}��S?��9�������n�?v���܊֮~�Pw��4G3��&9�������ܰ�����٘������i0a�Ыˋ���`�0>2Ƌ|c��=N8𭦗˻e�Gi��}Ώ+� К�]��e�ډ�kljO�sͼ"���1͘���{5�2��~ృk�x��O,�֑�	㐃sPK$��(ֳ��g�p��6���K�uVfV�\m�{�@���}��¼"nA7��At��렜�d	c@��g���g��?ʥwX�y�\��T����|���6"S����i���M^Ʌ�C�e���:��3�H%ˈ�Y��bw3�%�;s��S��k
����|��|�܈���@M�3a�u6w������.�1-���<�%"���(��;"��(Ʒ�E�4äL9�:kh��u���d��k��o���&Y��c�E���y�����O,n@��lz��^�jd#�b��L1�׳�ǱL6������6Ⱥ��4���F��zw�~}��I����D��?����b:���N(NM�u���:�Rݼ���3H'�'k.�����TDG%�<���f�%�[x&q��ش��y�w�oS��|z��e�W�V�pN�k�-&���9j� ��ĺv^�6�JL�<tKVrY�8����=o�[/�[n7:gphuˆr�˵YD��^s�5���f��]��|�B�75ҡ����L�J��S� ���v:7l��R8
��̃7V�K�4���2ַY����2���n��Y�du/��K���1�tJ�ƻo�&6
TJwWn��l�כys� ��`�����S��w:
Ob���ݶ���)�G����k�eև���9	���`B���Xˇ'1\�֦5dދ뜝����.�;h���h*}s�ʧ�s�Nɪ��.�_�������=oJ��^cx�pO�Y���-l�a�Ma]\U7N7@쾓�#V ��nW>�oC�	� i�42ܰ�<P�����P��I)�u�VH4|2v�q�ys�R��UӔ.a�)-��ΣM��!+�G)wY$svX�����lq�z5����2�Y"A�BbK�j�Y]#��u��� ���J�B`bf��>�4otU{Ա_Zgtɹ+2�R�����a�uO�E2���Y�շL�%��5�oiE�����PV%�� 0eTR�5j!S+p�θ��|��z�+� D�'J�*Ц�n��"�l�ȡȝ�L׏��:wo��u%Եvd�RGȸ�Z8Gs��b���mo:yW�%��\rS�y7ϯA@�5H_c���w
D
5�Vv2�O;��)6�ɢ�^��s��}�(FZ��f_�Fj�6����;�	�!���B��h,�N���%tʂJz�[!��u�ո�zQ`m,9��c�>n���(�qnQ/���v����˦�������`|���t���{g�#����Y�3���V
쉤�d"���q�c�k+�.D�k-�Um@:�7���V��Ǩb��	[�]�h@���Ky�.��ұ"�弻�p&zpF�@���j�Qݫ7�*w�\���(X,�8��-����؟/��X��!�YB7&���dE�Mv��<�3���A9k8�ci���̰�kVo����Y��zԗu�.�남�:]O*�2��C�l�z�j��ԝc05��tn�s�4Ņ{91�@��.�JV�<��u�s���u+Z�Ω|
��)�2S{y,�[%�7r�xa����lí�a��]���Re>4k����[1�u:)����D.�yA�V���*V�5�6��ʁ��c�d�m��v�+������
-�E�o >���-f��i\�� �-�;���vt�,Ū��+jU�����V��3ۏ0l�c�o:�a��۝)��;��ƍ}h����]��;�:�eL���h�0I���hpT!��Z]�!�Z�pI� �r�y��H�����9�]��ݘ�_��c�
�j	��H��+���M��)
iis�������������������r�*�'��"�h)���U��U,Eә�O��Ǐ����������1��:���'��jt�5�("*h��CE��|�Au�t�'{-�Fئ�d�)����L�=X*
J���R�����-]mw��!T�Oyt�	�j"������SS�EbqWP�-f�N�>���B$�:�@R^�U5��KBSTC��*:��DkEM%4�]@h�H��؊��*������$��*�i���OV����)hg��*������h*���(��S���2UQT�U%U/��Gx17�b*�m�u]#j�n�U1h���{�u�]A2Q�����ՠ�J"�j�=�����y���:�%+L*�"�p�԰8@�Fr�o�?g�:��^�׻	�_�Un�7h�ɶ�T.47�focC���荒������{�{޾���*V�͡���tK�A~�2$�4�U�\��,ܢ�a),hr�v1G>�z�lJ�+��"��ć��D��������*�	���6I�c��ΞeY5�!wN�V*����c��ck�,�{p��3���5���,�:c�[&�еnd�պ�.���Y��{K���U��A���+�	�4��a.����%xk�Y��D���O�<��tk>=�Ew~]1"�^,!��P��*�U��a�v�Է5x�/E�3����h����ذYeN!�"u��zT���]V�onIa�bK����I�T5	��qL��^%�_�n+���7���>wd���E�E��z*-���f�e�;�'6�f�zdz��ә��kn۬X��L��xjB�38Ѱ&P^�w�	>�5�my��"�	 5���+��Eۡ�.��D�]�ˣ �渥��>ˍn��r^Y�>��ĸB.�����Y٘lm�G�.~X�gR1�8��o������N��W����do�m}�cC�`��4#�V�2\�1�Ī4�:��iz��'פs���3�RFwR�a�DM�B�Ŷ�ͳ+7�O�����
�����ݥ߰8gd՗F�g)��*�����:�Q�Z�MޭD�k��<�[�C��)��u��ek�/����u�
CL���=sΎ�G�.s�9�����®s� �v[5S��E�Ƈ����2*X�R{
�h]�Ӛ��z����v�[&{ѵ�'��/Y��-4y!{�{^��ނ%1�ħ6R��,��-���ey�J�1���X^7eGc.�)��ѳ&�ry��e�H>P�9�v4'݆�����x�I�s�1��&Q�c�\
2&�΍���Ң�k��>����<1�/��K�P��)>0�ʥX�ǡ��5�Kv5���m�.܅��������"p���=B1��}��i;�����7� �QX��Q�S���݄���a��w���XG�̛Z�p�n��.�OI`Y��;��ͩ�X�_gܳ͋�I�Vc���l4';Nߥ0��F6�y�;l3�������x�lդ�Mhv�+�/��
��kmtf�h�ҵ�r^�ά�iWrʹ:-��@`���h��T�SF���݅P���NZaٲ�/b�h��*Lq�u>��>�z� s�f8��}Ұn����n�ys���L'�X~�F����l̀���|_�1�Iz���D�z�q싷�J�l��$<�������,���h6�hZ���rP�PZ�'�,��S]�5�lݲ���H�'3X�������S�p�M5�[Z��+*<Δ*�V���q����U��]%oU豻+�1��[p����/C��]E������������x/��@���Du�nEk!	i�n�� }f��=a����J�X�0 [� s�~L�/�݀�f���ޠ���]����W:�˚:AaI/�k�����E��ktױ2��?^>Y��B=[ѿf�֭���=	bN4	��7<5m�u&i^ܞ`h���#&<��~����8���,���->ABi򝝷Z�i��uo/vD�kV3����.��cH)*f��;(0������z͛OX�o�K��-�hm��(�U�[7�e�Q��pγ����6�w%��oW����lb)����XQ>3��1�1զ��. �f�܇\���q��Kw�ޝ�Ed���t��Ƚ���+Ti5٢��DB&�mn˩��R������iA�e�D�_�Ȁjǩ0Y��E�})�|1��1ɝZ���=�t�]�evr�Y�����gX�W?ɏ1f?�����~��f
o������Ҹ�w�S�o���c�3r�t�Qr���(�*����e�ϑ���G���M��x7TQ��-�v�m�d�vv�iӺ����.�jt={�Z~Y�R	z���:��`y���`}��~��wM��7۪fm�k�)��Շ�F�=a�ѹ(�ʸ++�J�y8���-����WJYBu��ސ����]�#��H��q��U���/ ���]`J�9Κj,�y�cGu�0�8Y��OsȯE�� �������1�FG\M�@ ;�yǽ���Ǽ<<.�q	JqH�xeo��-�3�s]���y��G2��9O���K���wh�±3.���M
��a�{���b`�^a�>����OH���jބ�YFM���b���8��MP1��sv^�����H���d������h��ʢ:�F�jÙ,:�����m��/w0���-��qKs���#�]�8�����sX��>b�7����Ő����%j�1]u�Z�{��I�S���C��A�eh\Q�?b���J�C\�^�X��E>!53������徫.�&]�O���C�~h���dK� ��m�ݞ�q�SZ�tI����xy�[�
b�S���{)H��]����A�}�Ff-7��Z~�6
I�^�!�����d�X� ��-�=Ŷ'����eY��>9	吃sRY$5x�:�X6m�6�ɻ�e>�W��U$�k0=�Ǧ�'r⭨.��Y�A=x,�,UD�geb��Ԙ�f��t22����U�O!ua�!�#����M?k�[�2��ٰ�Ů�i|�ù�Y�wwc���4x�V� �*M�՝Y����8�]�,�mu/Z�� ����cZY.^Wf���������]G1JCp�>W7$x�^���>�1s��4���)�5k�*�on\�p�wRY��+� }����������w��Au�]��[�'��E�5�8�/P���H�ޏ(2.��nK�i�<�	�{����̜�/ѝܹ����n/f"S�	*�ҫ�!v�a�e�_�a��xc_|]Q]��5x�7/�=R�!������0�7��e�KW��V{E�ˍb:l�|���3��kTU��'�4@\�C�NhL�}YU�k邞w��"���\��m��\��gY�����%W81 ��_ �X���@ׁ�T"�.��B��¬���f�����v��Ͻ}���=��"��@+_~Aa�^=17�/:ꀞ4,��n+��akZp�8i���w1�'z9ε��d�A=����Lj7��p����c���C��ޯe+k*#Ej*�e����w�gOF����zN������%G0����W=�~������xk�ܨ@���+p�q{F������N�U�kj��m�Mc�y�3���/ʇ��_�z����U���|�Ǿ���X��)O/}�2s]n�6�nQa^� Iza���:"��g/�s#o��׊͖��}�3Nq�k��f;����l�Ҭ1=��N�{B�����8���f�Է{J��*�{�`�wMO�I���/M�Uʆ�/a5!���{oo�\K�_�J���Lr��Ln��ؖ�R�6빭ˡY�߀O�<����xx���j�ʝ��3�9<�y��ި�S�v���lap$��E@A�"f��wN�g�ڣ�u���o�5�#(}L�o�e����5�e�̝OsQx����֛�$<�_A���<9��͙���fE^���B��~���R���\v�ܡV0?Ņ��O��W��M~�]yU��)��@�~����g:�.�`�K.D�a�?_�[�ȗ5���A�2��ǃZm���X�8�VK�c�W'�[��yK[U,�

��`r��PX�Ru=�(�^?{�ᩭ��ʐ#	Sղ􃆚�۱����|^��W�5�nt!7 ^%9J���q�x����v(� �&X��_Gd��`�Cd9��pB~�pFٟ锝ax�I�3�����R��;�k�|r�fg�/_T@�7���ր�,=K��7�D��.�}]0�r�E��Vi����6FZ��Ѕ��E��eأ��׏;� ���#�&�d&5���Z�U���fV#�1�����u��t7b��X	AcK���Rq.�;X[���:W��9���>�������Ҧ<�]4���܅��5a��bF����c���۷�`~���.�����]�*%7:��Ϥi짷"��r�>s���Ā�ښɏBh.G(�oȶ%a�;6}���8�ש��3����_9��}��_�3�99ȫ�{��v�+��G>��oQeɅ�c%U9~��-���.��F�Gs��T;��@�����L�5�{���F��QA8K�Y@I���ɛa�ac����{V����'yQ�t^e��3�/V{j��gS��u�e���;3m����+�T���/{�}8�o��v���%��򝺩�Rjv:��P����x���u�3'��>��)9��=)�qh��=��F��ߧs�����`� ^�:	����;)�Dעb��>��7�~��_}���w�u��I���f�{}*W{,:}ƐEr5>/��ӱՑ,��KHC ���$�%���۬�a�SĐ��5x�ۺ��#4�e[�L�]�XrW!��O4��T9KL�P��4����"�6hV�TS<���U�K�Vz��61�o�b��o�k	A�,�`Z�Gh=fͧVtg�Uՠ�Ⴓ.?_��Kr^ņ�F6��u���U����N��lr�2���t�
 �f���QF�>ڭn;1֌�s��]��3����D?.����pk���N;K"�R�~��|<�4h�`���*�X�[C��r��/�;2�!�bX�|me�-4���Or����p�wgU>m�gĵ��82�E��"������J롒m�F�ojmn�
έmt�t����&�,1��[��MR�j�E�c� /?��8���w\�Uԥ��ҳ�|��Tm+�H���"v�xGӰ�E�}�N�� ���w�E��n����b<��[�F�[\u�5y��9.�� (���jc�)��ټֽ7W�H*��E�®rt���`�F�*��z,�c��-� �z<�Bmۭ��i�*a@���w�g;���)������M�M���-?,���Dy�tS@}l	�ѧas��zqr�����+Y��p�<6�옖��@W5�E��c�(�z��~w�(��&��t'sʦ�������}
#��d!{��.�	��N��TwU��BO�|16�=D�m�F:����]����g��"ry�P�.#��{�;k��.��>����s%�S�X��kr%t�A�k�6Wv��b��6�>��C�}���c\�9��{���,Ϸj��n4C��K��k�m7�ڻ\jl�Dw����:�_��b��a �2����9g�V}��ՅPW{J4v�6*n�1��gPmy�P����C���Lt9�g�;��Z~��D�� �X�{�L*�>�>��97Q�Y)�߳�UVR�N��#p�핳m<����V����P�u��[1�o���T3�� ��l�έ�x���0�lal�\Fmv�#���5&e&j��s2��4�卌����T���8��*ǽ��������  2��H�4�u�2�xz/zb�)��v}�hM�Eڒ�d�3>�ƴ��y�����F�޻���F;��Aa�-��MG��gc��fnCkq��Fu���&m�y׬��T�蓔��8��|;��ڃ�2��ks]��d9/6���Y�A;>��5(��u�w�^Or�[���o�C*.[�k( ����F}�OƲ?�?�u��7S��;���m����D6��ukM
V��
e>֋n��u޸�x ��(2.��N�Տ=	�K��,��ez�c�S�ד����	�{1�X)P�~�E8��&�=�������X>s(����c�胵2��3t�j�?��˗n��7�Re�/4x��,�D�&:l�6S��Mk)�پ33[f]n���1>�5́0�yYU�i��)��)�Q����Z�4Q6�N��:�_e�l�;�?��0�D?��?�W�wJ�]]F��]xi0��(�5j���ogt5��=׶>M{��չ#�h��]�!�|m���q�L��<4s�q�G�:�W�k�(m��0�i���<q��a3C�P�Vr�PHF�:�䂋 K��ݤ�˥�����СU��c���SV��m��w�.��x<'A��� S�̩ �|�L��Xz;:���r�\�������vR�ӏrh#o�7e��g��������3��͈G
��_,a���5>�U��)�Z����
�!��X=�4� �cB`kc������1,�3��ȭA�o��m�˥s�rUO��Bi���]9�8/Ŀ|~��<�\2��WD.�`�i�	�e�㔘kP�*��2�~.���KsQ��1`�sp!߫4s�erL��r��(:���չ�f��v���n�a\bK�wco�2�>:�lj�$u�%��f�#��2z�������"� �L�@��V~>;�,���{�BPh4y�\�CM�qs=gN�(m��ִD����f`P&P�.$̔��5\�=���ּrC�D뽃���,]Ȩl��*�y`�˨�.k�"�)�t=C�}6�#DS��I�T��īy۬�N`�2��Lgn���sv��^aU�K�iL�p����T9זt5��rۖ�j��U��U�ys�fh�]��{fa����M��Be@,T)=�]�,�^>�
���{gm�u�¥qu9��ׁ����*`w����S�΄&%���R�:z
��v#f�}�+��Pv�z�bZ�k��r����Z�tz����_:j#�g�tp����

��s�DէPݪPʗy:Am��G�NN�ןs�8IN���&k�Z��p��hM�4o7{�5�f�v8u��x�g���P#�^����7�{�C�ҽ�W+{7F���a6�Cy�qp�*��{Wׯ�4P���sO8K�3G�beT&md*��Y�u��Ǌ�a���Ð�F��'k�6��1�f��āBBK*P��ep�}xv�ۡa�9���޳or(2��R��et:kn�v)Rk^s�*�GOݓ�k8:"� �]�]�S���Ƭ�ј1v2M�C8U��R�(]=ԅطn��b�q�{�����8��1Lpj��3@�U�2-RdR��� ���??���{�o/����M��%n�ˈ��w��f��q�ݕoL*]nڗ��6�^t�=�5�n�oa}�,h�Τ��[���]�R�T�i�0u�v�=�[��AQ̾��'�,uc�*�8 "j�(�*��Ҡ�w�q��cmKgjV�}8�v�@�m0v�f�weꓯ�,�B�����̱�Ù����H,�X.8}����q:7������ը�ruT��l�����Y6�,��qkTB���Tw�����m�(�w3��&��L�b*@ZE���N����s2r����by��Ի��-��}=g�oV�t5����D�c[�U�dmLG����V�I�]�݈��z���u�W�o+:�>7�uS^եZ+jߖ�;�Z}�Op���]鸎��9۫^S����b+D�PT�ԫn�]5W_'X�(l��N��9��ݔ%t������K7�8szul]�[��;��[Aض��b���B�^�<:V�M��F�����gcvss�E[�:�9U���ͽ8��:X��seu�[M�k4��]Ův����-����xլ�e9uƴ���c��Y�C.�ղ���^[�ŗk3�K>}�v�a��(k5�z1�s�-��!�j��m��y\��^Xt�+o8d\e���`|�M�L|7^�:pSǰ!|��zdo��0#�P���U��8���T�M'q�=I���`����3�
�&����T�{`X�~��;��j�eiG�S"�M�����\sV��5un9>�|���WQή�b��E�K+����E+�C���,���N�;�uʒثF���LHpM���P��s�[T��k'~�D��/�j�Mؚ!�C`�1!ۭ�N�;rJWYJ­Q~1=eC�<ㆆJ47��K���@�v☹Jl��,��+��S;�]�)+nv��n�oOm���>M�;|;��	�Q燃��n��[��^s�e��^�7���[H���E��p��%RP�lQT4���%��%14%T�H�R��l�}=��oǏ���||||||~�����ד��B���,E-3Rzê
���J���s�������������������hhX�
��)=����j���&�k��X�t�SALIUCHT�T4���j�"�Z*�j*�;���jW}j�j���h�OV�V���5��E-Ru!���� �m��kBPU��MWRM!�����Ά*:��J6˧AOQ��W����:i�tD�覀���Ж�C��tm���I�:��%'P�i
(
&�v��`�M:=1ԔPU���J*�MRѢ6J�R4�5Z�S��h5��N�SI�yW}V��vh�뫹�S���3bD�L�IRaG�����X��G	��Ns�Es���;ҹ���(��e�F�v�퉰�ح����b\qS�|p����r �lg�~n%'���A��E	b8�H��$P������}WG[~a��83�--|��㮮�	w�ﷆ�E�at���T���TS�{�;Ǥ8����DE	�By�hOa�H�):�]zi�:�yc:q:>�_7ú��Pj ���_�i��9a�0\�|���\/����Ux�az��蕕0����l]з_lSu=N�^/Լi u0�����>���1�����(��5�(Dî�ו�_����.�W�6�����p9�(-��0�ԜK�v�}�?���>Oia����VnX���U����dse����Q��Q��n��X�Azp���<>��	������4.�+�/�Eʘ��OV����0�=+^ʂ^���\sHWrʹ:-���%�OYة�kN#��t�r�u�y�#O�@�n�u��yw��}<?.g;����sM�ݑ%���WO��
n\�J
>��+��	�`}�SVyX���f@͓��E����<�ϫ�	#�-s6G`��d+�P���"Y6u�vS�w�O���Cap��ڌ�K	��M��-ƞ�V�aWugZ��
���4$�P�� ƌ_��鮯ݤJ.�ta����j��,��<���{�zL�֣or�5چ�5��k�ۗT~xr����G�\C�	�����~.���������D7o[�R �CȎ[��{6w��p���[讞����A�U�#M�ɏ�vo�]�a�%�Ou:���H�v%�9r��������Q�����������('�۰����}f��nt�N��L9+���0��^M��sͼ4���Mޚ$��m�ob���LC+ٌ$�Gp�̽6�lMO����`�J���vW�'���z͛O���':���ˡ\��mfe����h�g�!��Hp[�a{q�5�j��W�H�"Sm�R�&X�S��t�1���bC}w+��Ұp��굆Rv�ۺt��%�Ȉ�հ�b7%W5tB	�q�d^�	7:��)�TN��m�w_�sj�4Z�#����^Ew�!�
�Q)ٲ�,� ��<�d�2}��#2/&�()�'/�I|�[<�t	c��I�E��?Q�}|������k�~��:|b��8d�Z�l�sӺ�;G����q<��/��Rp
�'�W0��e�>G�e��3V����|ւ�tk�S����'L���6H��j/`aR�"�&�z�(�����_y@��,=�!�s,]5����|e����1�ƾ�i�ճ�[�9W5�E�H�0��Os��plE���9�gq{�,��vB��v8K ?`�	�&��e�C������zd�/d���DUQ�(e&��u\�V����M��8��v�CZic��F��&����u�6:��z'rb�MEme@�2�y +��4�k�	z��u�E�s��!hA���E�ؕ��<ۍq6r��r^ғpѻu40d�V�%If�-2��V����|>UUS��ȳO�������;�.v�kyϡ�\^��_'pеa̖ٛ��[�`fy�oiz�\�·wO�aO6��A�#�4{O䁡�B��֜��#�ˁש����E���tvu �6p�y���+�X����ˆ/	��zh�Ӻ�1�N4��֫!�;�T�� ����gw��"w�f��v-��C�����q�W�n�����|�q�>ﹴ�ӆ32�-�Lus�N�n��3s�M���)�A�ș��o�iӭu<񞝎5z���Z�x��-�e�`L�#5��/Q����+a ��V�̖A��]xJ��}ا�53�c�G����Aʒv>c&��5���\�E,����"ؓD���3־ݦ�cy�/�:�u�f����.���u�5{*.ۆkAA�e{U8�����t�&�یi!��ӭ�w�7��u���QE��"QUE�5 ���#��p���9oj�"�t�ü$ ي�sTMw.���a�@njY'�)Ք�Z�TS�� c	�dS��ط����7�;��@�v�e�j�#����M�֯��&�+~����=goGƻ�JR������ם���>�r>�1��������u�%RT��6�WJ�S����i�`'�Nt�� ϞJ�4Ī50m��Fʴ�I��(�O�����]�򟗱~��x(���􃉇�ݷ�6{s�|7�Re�/1V9�Qz�\h�e�VԠI�w��M}�:�xa��A�"�~��G=�e]�4އ>�Si�S"�09�2U��<nD��p�b[zYW�Eٓ?>8{h �
��R�7[З��]F��I�חh��B.U��mU�7u{0�̟w���ƱD�~=a���*N��2(���WK��1���S���)�^"���y}yW����+A05
OB�01���^{�9]�w*�A��r�j�k$V?�hO�:���.|
�������'�Bi���]0B���%�P��vX���=}�w�}�K`�Y@�)�m�ܤ�Z���X!tN?0�9�b|����0��Ϡ�Y<Ԫ�q誜��0^��-�p� ����s~�:��f�;r�Gy?-�4}��m�Pk��@|�P�툈W~�i�dgםyw�	��
����E�;T)�5��`T�8�{�A!��i�!��odڌ�ѝܼ$4��6�Tw�r�>�`�1'�ߐY���s5h~�S���'��3�������=�D�\�8��ǅ��fcs�n���[��FZb�Mvٗ���U��
�n�7��v��,�o�����٦R�0�����>V��n;���K��A�A0���-�K)�Y �4>��w����S*\;`�{����S�f�z�Wݰ�!T[�a҆�h��VY����{��U�B�4�`�q��t�ê�x ���8���/Ǻ�H��F����}��m�����ɘ�=��JB/{��*Y�(�'\?�.b��ĳ�!)��ƪ�Ͷ��[��_Uw	%�8�y���{U-�΄&�P*�®�}ך]ap�u#�����|�{�'b<y�h.����&!�>!��O7:��x��(M���%P���m�$���ϻ������J$��{�/jf
V��0j����-����lA.c��[���/�O9����،��E�Y����`X|��i�Ǒ7�����E�z_'���`B�Z���jY]��5�k� 7jy�����v�e�0i�S�mxw�� ��Dp��~�TƗVKf�'_T��|���7u(v�;��J�����֔+���rq.�����0t����q��F��n��HR��zzu�jNP��F���s6)P�zdi}��v@p��T���t����J5!�\��-��4-~�LKi���DŰ�=+]{x%�^վ?]2u���?}�Vr�y�	�J<.īXD�xjZ�����z��mt���U����:v����4ev��Ÿ���'�z­qH�H��. T�?(p��M� ݕ�R�ʽ�7�A1]M̫Z��F�A���V�b׎������*���ʶ�k<�r3��A��_D���������ϩgz=�K������f�����Wj�C���uP(����P<�о�����?-����~�u���9� dRĠ�gc���^�hi+�ߩh�bՑ�k�]��9aC�p����,����/㲽����js�g�5+z�X8��Ј|,��z3�-�Mn��k�|Ş1������m��K��ʚ�Խ7�V�͡���Y�Gd�Ie�2a�ȼ�O\�o��ĵ��m���e�ulX\���##)��O�=z�1��Tͧa*��s"��z6m>b؋x6���7�ī]/�N��ŵ�����V0J���>�"Sm�R�&��i>JUs�_��>U��[��_i�x��Z|��Y��dKw���dC%W7;��t7����P�݌��y1��f��v��i��F�]�{kVW�~t�)C�d��#_�X��A����� 먡�v��_K�ooO�w@\D��|1��]"��F���9��.WG��m0��k��P{9��SfI���i��v}u5djK�p�e!�6me�̾�'D�>5��<�]��9�e��2�<&>�]]�2b��e�� V�2�2�r�
���r�����q�˔힓0�VM([%���M��]��q{���T����7�h�:��2E�.ᷤ�N]�?9�QϠGj�F��.�/3�:p5��`��D��!7W�06Ƚ�j/�C�0���='�C)��#��a�!���/ξ�ؕ}��ᨃ;�u�#���F�-z��M7X�U�xa�P1���~����r�XO�Ǻw�!�~�/�C�n~�ߏ4��w�A5|��ywJ5߆���Ǚ�r���JǾ���E��]�(uύL�I�5�x"��$N���#� ��^���6&��c6{g��q����V;_��~��=��Z����֍E������:�ۺS���
���E86��0�ŠvQ1\���&��$���pptQx�3��~Բ�{)�`�O]bT3��s-��7h6�v�ey/ʻԏ���4'�;���?HX>1��˫YP�wN�!��Bi���V&-��߆��//�H��%�%�p��C?v9�����+�7���mة��4S�/t�w�
��D����ؚ��z�Nֲ�(8�rnl�'�����!� F�71��M���M^޾�O�D����������%n����1��۳�%��*�l��1 ��M�m-��ȵ�>q�r�9�~�뻵}��<�9Ց܎�
������i�B�ѓ�f����!W��%@����im�a���W����m&z������*I��?`|��_��=�Y�{��T�"��nZ�δC{�q�Ad	cEuk=x�[�W���͸f���sb$���D-߼��
�)+}��k�}���d�'.�2��򜥭�B��,%��8�/P���hAoM�s�ٝ'u�"b9u��n��C!�ݫ`hێme�	���b)=��R��IN.����7"�R�����*��"eMf��~���8?6����?S�.�s�g�sJ��x	���"��+�
��g.%�q���ҝ��K�u<0[�!#ا��s�8�U�]�fy6��<��b��f���OM^�p���pE�v��MoW��k�p�Ѓ�����>K��4(��I�oP&�+{��&.{3�k��<2ܹ��9bF�N�Bxw�Ȉȇ5��;?��yP�y|�}�J%Ӥj�?U]��K�.� �wN㋿rTX,��TZ���+��*A1�W�ó������&��u>�٩Vaȍ8Kr�	�}e��Z��N��=+^�T��*9���:�=��CS�+�G�|)o���:[ۆ���#�s�	�v���͜o����H,�F���#u*Ôr�:]3&��ӽh:�l��I�]p�{��*N>��]OkOKJ5���WM5�
�fм��S8�uouwN��q��-+�-���n.9�Ԇ��ƀ����c����,9?V���qǫݘ�G�0�/3C�`,S�| 9/0��~��es��H%�Mc��B��Vz�Z����Y��ڣ�a�}{��g��_�
�~�	C>$}�>!���X���Pf2r~���Gy?>�c�5Z����4��R����������V�eyqiP��yXj|��t죻,�E�[E�<�r����U�1Q\�XYk߉}͟��;0N�=X�? �e�Ӥ�h�k�n`�a�r1fu=�o���8��lo��s��\�)^i�)|k���Hp�,>#�w��3��:����ѱԞ_y&�����i���&ކi���0:�R̠h'\=ٶ.b���g�ʈ���B�-o\�g�[`��v���2V6�XN��o��ʼ�P���]�(�^<ȝ�\(1��q���on�v?�w�`�����93�>{N)�|"!�>!��O5t!)��Js~JSڭ��>ߞ�F��z�%wI)Y��߃�������
V��,y}ಣ|��0�v�0�oT��P)�2�g�q��a-��������(��=��z���]�����K�dp�
��5�5\�DľYD1���#�G�����G}^��
�k+#�t�%��Ӳ�q;��{��.�q��[��7�]Po���?�, (��Ds���RW3�������+����@V��e��f#�Ӛ���w���[z�%�;K���:�����w��^�}�K���{c�"�l��ǆ.���9m��;�B
��	��͜�
ӈ��hjչ�ЇFt0nB���B��q�ʞ�������Ƃ�0���h����.�K�Ӝh¾�L��T��8B��	�L9�:�0b�3 6��ը�0T����#��8|��vu�DH�fP��~�<�>��`��>�xl,�)�Gu[
��eA/r�����|���oq�4E�f��-��:
�s�����9j��Y�w�wy�j|��:ִ�g�6�#--f�����B�5�r�]5��v3�����:.���D~Y7 '�(߄�l9�~����}ڷ�q��oŎ��u��*<p��z��!��{��^�S��Ӻ�&B鶬�/9&�����*���������MCg��fF?�TEC��g��k�X�579UY7lv��Z�B�cЗ�zW�^�yf��z��PB���q7�m���O�R�S�̺���k�3�M-7���l|�;5>����Ɛ��f���u����w��;�<42o ���
�UX���Frҹ�EL?�m037g9����I�aj���E�d}G6�/V�xֱ�v�b�D0��1ro���':�Fq �.�CQ��>̴���-�ˋ��)W'5���v�!a�{ɃT��m~�Y�������׹Fj�q�{���#���92�N��n �b��m��Д�l��r�混K~����GP�H��[��h��MV�XZ�����'�gp�*�Vͩ}E�t�a
Zb��\�q|�j���=b驤�V�_��N�7��5���eh6�*�:Ef��-��3@��� :jo����5���Y�(�vA#��U�AfA���ki�4`M�0�����rT�\ĳ�;ڗ���?n���w-��5�+�B�l�nV��&m�ym%���Fd��Kr�k>�'���J��N ����S����g_c�j)��֝A�J���ڗ{�����l�*��̙[#t��J�҅-ێ>�W0:շ���ݝ���ľ�����^��Y��*)�O���4�uOcK�rV\�o�3�Oj�[c��y{�����K�N&�٥7d`��g�jL��\���6P�$AF���t�}�/������b�Sf�k���&�w���Nδ������\F��0=[)��`3^ԧ`��3e]��%ƚ�HV�<���s�F!��h�@S�
�m�ՙnU�1���-u��r7��9@U�BO�˴��f~���������J�0U�B[S�is��}��/�=
�Oq�e�֩���㽶Й�m�Ÿ�њ_kt�IJ�2�ؚͧ�3`<�'�"#Om�s:�2�H�!�c��J�	S-2��2:�n4r&�p�39e%*�����$�/^9�ID'��Ǘ(u����άt���|�
�;m*u$��=O��X�����w;un8�-���+9�a��Օ�E-��gZ���>溘Q[���C1�y�C�ƹ�,Tn�ZZ�Zr�b�L�b����t�w=���*�yDԡ��#;]��M�c���{�8����R�n�/�z��}k���tTb���T�W��p6Y�B<x�XF��p�
�ö���ѣ�F),��&IF�jN*���L]��~��h{��Q��`(u3Ջ��7u��e9�׊�}��K�2b,�ݙE�r���y�d&h�4>�)y1ml�qPK^=[FM�+:�l��	S��u,�~z���ౘ��r��W�-�ڰ	�T8��ʶ����+�c;E�5��
O4. �\��<��]�꺖
���i��]7p��*0����2��ds�ݬ'�����[j� ��RFTi@����8Dv;/\,��6�D�Wi
�7�HKA��y��ݰd���g�:�s�k%�ů�\cBҟ�I�{�׼M���m�����>�U��z���D�5���=8�X�ƫ�)���%[i��t�I�N���i{�Hj�m�uI��g9���x��||~<|||||~��W�v��MF��
J
N���CIH��:
4�;9�ק���Ǐ��������������G�4Sܣ��)(Ѡ��m�mOZ�j���l��F�#A��6�HbKU��@յ����j����c�gl�����%��N�t�-4�t�i�b��]uQ]C��4�gAm���.`h��)M��Z֝;`)�v�IuT�[[N�[`ŵ�4Mvѣi5F�Xih���
�	�CITih"CEPn�X��ӧ�몝w	�Z��M���ӭ0��CGR��j�:u��������@��. ЕEPf�؊(GA��Z
)/\瞣�s�z�=�6�ܨ��u�3��WW��{�d��N��Ka�>������+(���\��Z�{�:���xx{���:�A�_��W��VVN��v���!��v�I�Ͱ&򢼸�M��Pd�4Tu!o}���;w�$�v�&����C��ɪXp��6=�M�`��}\s�U��Z�C��N6��쾼�#\!���Ȫ4'��[���P(lM�xw�������v�_�42��=���m�K�k B2q?;�I��JsiH�4Q���r'�.W�= ���m�[a#����z�XT&e��A���.�Y��3MI��NW4	%O0�K����y��3eK]6���^nrrv��|8`��a���'ʯ���nY'��-? �sZ�@��{�9�D7PP��;)m�p���掯0�a�i���*s��Kv��B��̮x�2rV��]�l�e��*��룛L��ݔC1��~�����H&��t�.�Ӟ�n`�������77�ꂾ�5�ۛ;?y��~~��k��K�A@pZC�[�2�x���zݏ:[�Mv�v�R���52�e�ǣ��di/�Ӵ!��(h@����Ao��9^�a}ae %�2��9��ÿ�]2�_�H�/��M@��d�t�[Ng5l?�@m�x�5�˔�ZĔ�́�����l?X�
*�\��ZsM྘7sy�����*�;d@�Xۮ�uo/i�i)gW.X��p�+.�Y8�͡Yfu�J��?ync�����0�n��'���pϱbhgJN��Švg�7M@�c����#Þ�"��;���9��*ge��C�ss�-�����B���\eۚx�C�DYzD�f��x�u^7^<��
�%�D�g�k�n?yPj�����U�A;�=$�%;r�.���r�ކS�7'�?3���+�<^��ʯ�=F+e�Q�y8�A!�[ͻ��(?C,��W5��ZYwd�j���y4ʺ��4f����Lw��]�I���\�v���Q�9㳹p�ti~k��A:��}�V��Ԇ\t׫X%��]�����;�;1��Ou�'��������1���!���ʂ�B���aLv�˚{��o���e�p�|9J���[f��吤]	��i�B�%��tBd��D�E)�RS�|�a���J�����r+W6�f�h��[�!�����rm÷���*�,/2V9�Q|Q�M�Y�dv�N�o5�~8�D�<�S�?;���Rb����p�}Y_v�}RS篞�z��4�F�}��^8�׊c�7�]�wR��Z�^��Ǚ�����rCc-ҭ���,�)�������Y���ɶM�R���okM͖s']��Ͳ�f�ϵL}[۸�N�I����ET��J������R��\����0t���Ǌ~�7� �o{�����%��lݯ�gp�g1� ���=���=�y?���0m~���@,�A�ꠂ���Ð˞��t�T�(�هv��)��XJ���<5��]'���F���P��=�>;L6�@M��Co1�*�o3���c��X�zh�հ��qS��c{ƕ�qz�s[K��p��lm�L!\�ǹ�x�������*`����E�P�nd��ҵ�$�[�~a�YBu�����W3�����Ѯ$wD��`���<̀��=��̮F]s���e��|���ƥ��ʥN[D*���!�[� ܡ2���9��gA@x�	�;�\�2O��كqQa^�\�Nu�`ʕ�AQ�{������b�l}����1e|�(���z�@���-ӶF�i�@�k�{�-��������\н[#�~Nm$�4�m:�O��́q=�\$���PZn(���Ӡ�pfgvu�吾�i����W�yҏT���.6�51p���B�sآ��
��e�s�f��Y��ױ5MږƮ�!s��A�ːt�:��6m��� ���-X!c�kB˓p�)_�fQ��_��9Q�E�@y��{��-ܻ�[vK ��r
���X����V���}�n�pG�1������z]CXPOf�vh�j"M��b��Zu�;,�+�fHѮ��S����y�>~��ՇW+g�� k@:9�C�4��|d�j���_���M�
�̖)��v�5ƥ�i��j;��5p"{W���{^���vC���CWB��1��� �f9�ЄˌJsՉ�'5�)��f�'�������u"�_�ل��"�2!��I������O���)���e9}�=��;z��-��TS)T#���)]��A�"m/��V����ݦf��O1t��������;	�B�E�X��lnWP�0m�Pw��M((f�:�gK��pѺ��:g (m@uHM�3�
�2��*z�(��֔5��a��k�����ڙ�=Z��\�s�/�����!i��-6���	���C9e���|n�U砲6��tf����ވ���xY���Vã�*~�1-���
eQ�V�eA/�}�n��I&�썾!uԳ*ض�d0b9� |y"u|Q')`����}vw�E�:`��V��WZ>9gӮy���j*��+��a1��Zsʢ?%��]���QKWX��U[��zTW�K���%*U�����Ü�u�3�Z�b����0�W��T��{;�54F_]8� g'�����%@1a\�I�v[���y�ˮ���&6&��N��k��Ԧ��+]��؛�J���s!��x7��G]k>~ ����ӟ?��p���w:��8Xh�M'���I0Xhd��uS��k��X����
�З-�����uci��$=��@3�&����ֳ�fԥ6������wsF(��͜1ae��a�jz�oF�ͯG�/��w���,��dÉ�-=U�}�#����p��꿲�?R�=L3��7����5>�z�1�rT�G!�	N0,>����9}�/f�(�Ę����2�{����ROB_�|���~��G�yQ^\D&��OMYw���Yr�ï��lo�\��s�4{��Ui�U�W��\an���V�B[E�c<U;�|k���_r:�"�[K�)M2�F�R���ח8�������y���xsDw]�Y�nz�S��r�ii,���rȺ���R)��&��������Ϯ(v�e�a��Ųu�R��Z�j���#l	vE����I��&*�9�Q��Y�_0�<�]�n6<�Oi�y��>u�	�`^����So`Bz��őu�-?!�W�\�~?|��2�����Y�O�6��k�A5�љ�﯏�b�>�����s曮i��˜d��iX��Swڌ�v��uޥ�V�UZ̔7W3n���泯^�Dqj���]gaĢ�̛�x���{�ȣ%˲,4��{��n��X]�)ʶ�"����U�@5c4N�zYY���0�a ��C�w�Z��n���B������r3����j&��zB7s��ώ"���ŀcɤ^;(��!��Q��z��j��w�����v�,G34�Uvأ�s�ڸ�Ǽ���N�K럘�����%� ����z�b�5���N>v�Y�(Ơ-�����K�1�e�~���aw=8�YA~���ܦA�AˬG����ky���w��*id=2OR��hnt:P	�e�L8��zLW1n�1���?�m�t�������w|����,k5��ny���⡅�*��|F�#G>|�r��z6��"�������A�0[���$a���6~w�� ��v��Z@wJMww���"�!]���\�r���l�	X<ă�솭����\�T/'���p���_j��#�؎o���Y$1FUĲ�#��K�X0"ä�꘹z`��驩;Q؟F�.ބ.��j�P��t�ncEuk=x�[����:��A@���sN���ye����eg'��eu<�biq�6V���Rm�T:���E&j�vb`����V_1��m[O�ȏ�W�z�r�5]=�����\Ty>�M3����*YɾЌ�ߞT�-a�*l��l�%>=�m�2�᧦.7��Gl��z��W�dɗ�j���e{�EZ)�ep��W#�za欘<��2ױ�*
VW/8��.�֣Qp����Cia+�ࣣU鬘<�>�-�{�K����G	���: �=��N��*���L����n^ù���.�)S�Qm
��oHkj�(8v!���v������׽J�nk�L����{�^o�U��ޣ�{��񊴐���>bxm�I���sϯ�K*Ɲ��;��a䖫��W�C�Wc�<��9���q�hl�T�:�
��}�~p?s�&����̟S��{�E��u�B���s
���\���45vø������M��4�ׄc�
�7Y	&�	h�R�*w�7�x���|T�
�5�I�`�{mi����������6+����.N�h0{ap��`c+�"����(q�Z�T���Q�%m	֝�|8~�������u��O�������q=ó+�e�0MC9*�K��|{`N��O�kl�+[�f���ݿa�������_A�	���4�Z댟�Y�����~����H�Z�@NE�ک��¥w1vf������:;�k�&��=���|#C�(��DoU,�w��l��N2l��� � �_D �)���DP���n|i+���7[��v�*(˄��}eܤgO�ǐ�����'�q%��r��)�1�ӻǀX�W�}_�Uc4���Ν��x.'�fD�lk�[9y�x@��h|/>�aB*-�/+6�
��_�]c��kA���݌h�vA���CI&[�}GD�9:L�`���p|����}�Z~�s�^���E�lkM�r-B�=�B5��t�:b��^Y��`l8`��z/x���Qas�����S��	W�ly@Z��Cv�EI�������\G`�e+�1�oTÔ:)�8@����!����F�W���aPP���zC2+
OOI6F4
���ni~ޭ!ؼ/иP�f6��>5b_������~����O7:c�tp��)�ݲ�׳]�@s��wJ`����]�6o��l����C�dȇ�`$����h�DJ��֫��WwW�y{6f��g�IΨ�5�&�<�=��uv����-|r[z�̻�hЦ���٢FHd���Qt��*�]ctS��:�r��^�3X�2�s5S��fJ���V�L��9m@Lm�ޡG�q�T�=r�O�~J��q����|K������Ñz���bk�7hC3Q'R�-�Ild0��� ꇅc�Z�W98�Ӵ�B���Tˇx�f��$-�f��V�sb���U�7�u����#�6-�ĺ���O�kk��D���MN�|Q�В�z������z�����fc� ���?>Li���&�#�9\��*�=j5�QT;������~ͭ,�/�����d:�<!����:��xlY;B�P���>���m�n�_]f����/��a��Ű}���Ð����_.2s
��~]-Ƽ2�.�nje�=�� �ϖ9O��w�lf~V9X(��	��/��~kNy���l2��l+�{���F��(WHfɵ=�� ���o6�����=_�F�����V�)Ĩ]��^*f�f1v����/Dܢ�%�]��������H~,��ܱm���0�]πؓ5ǲ���Tθ@��Κ�XG3��^�ǵ�oW���3Mxi�é,��y0�y�{<Z�cs�d�{w�C�g)Qt���O<���.��z��{{Nb@�G?�Ɵ�S5x� ��ͪ_[�C��[ʙ�y��-"�ٷ�k�[������ZLXB��w��0�T�o�Q^�q�˶�$�f����M�p8ܻd�MAdIz�]:��սI�Q'~1pXp���྘`[;�9��HŻiM�v~���Xc���6�:&�&a7�ov�ڻ��n��{Փƛ�Z���^�n%m3��Ȣ�/�U�N�=P�ֻJr'!�� Eʻ^_X�4��`�4J�y�9M��6���B�bYY�krao9��ޕ��$�{�P�{�	���{��s���'&���.�Ƚ���Z�B��6���=5�ߤ��~�U힓&�v7K���� g������y���'�b%9�%"��F�[X��P�ظu��IvR"���x& Xoi��l�w�}��o�!�z�)�ܻ{�7�J.�Bb���R�U�9�Wp/�í�mN�������~�<�a�"m	��� �_)v�,��zO�v�g�}Qu~}��2��j�&�Ot�a�߈?F`kÐE�^�J=y�P����v߮3*�N,�ֻ�cIGs�|wɤX�e���B��|{� ���OZ2z�61��Y��������!lP=@k]����]<�UO������n��5�3�����%;�%���T���{g4ÑXbgy�R�N*�9�é�k,{z}N[ѬZ���B�@�`�c����Uטt-��d�-0�=.��#p���I�>e�L+�@�LW5��Z�ͻ�p[:���9��7
Շp�;)�~(���o�u�����ݠuA���q�.�8˷5���0r�h�����&�ᛖw8�:(Nl�Uڰ2���iG^����Wu{�м�6uդ��<�9du���a3�0|�i�f^.d��"��������Ɣ�r�.ya��'w��]o<o&R9�.���]Y�{�����Y͵�x��K�pn��s�����0�*1��[�tL�ʮ�ݮ�X�k��0�f�� 7�oj>6h� eopӱ�'�˘���b��Z��c-��s(m���܎�dRO���g�^��)5���+����ı^5����;�k\ke��SC;�0��q���ɷ�hct�l�L���Z��؊<[�0�7p0R��pܣŔ���S0�:�^af_9�x���q)����OD�t�Z�십� htbh<���蹱��9�;�v9�w���v�j�<T�W�Eꥨ�Fi%����8;���p�NȗA-�i'l�c��*���.� ���>�4���yF�1Ic���&��c�gE��JtB����Z����t���׃�^��+�A2�e���Vec�/��Yr�d^.1Z�j�/.���ǡ�7�nl�Spj��2kF��Tu��C]�������ؔ��TM�YB�'��[	9�v�SIE:ln��Z�7��6���Q.�t��Y�84�VGt�i>YK2���
u�22�j�ss��^M�
����k�o��hm�c��5>�ur���K��D�4�/EѦ;J�T�A�<ܛ�Jx_���9]����1�]�p��u����Gʴ��)��DP�73,�`&��9��j�$��������g�Wo8@�K���'ˬ��]�n���&oU.E ��z����5�]�Ҧ�W(𿅭��帵���j�t0s����pNW+�X�ngj��vՍ�WIO�[�B$5��Ӂ�Ȟ��*6z�u87wf�:qQ6z�lq�1h��1
Q+��Pw[U��c�)ӶhuMs�w�H�k����AE�{]tD��T�"/-N��5�@��e��l�O2#�$=3g�A3��k�ǐc3��x���^^�Ҝ���`��,/�혓�G ��]�V^����[Z�P�8 �*�v*YQ�zļY��h�ͻ�.�ݝ�8��G`3.�Ё��p׉�W�Ƭ:�|�ifpf��Y�SgX��	[�f�t2��t(P�w�����1��r�83[,���׸��\S@�Gune�ם��rM��n���>�PX��V�C�����y�F��ɳ���,)kz���YT��8��H��j��~��!Z��]��uv�}���@�D�<��s�J��<'��Ba�T
i��6��.*k�3�փ��&����ĲR�Ӿ�GY)�{�1�cLpn����[���Ն+
�9qV�|
κ���ڒXfYU|��ˌ��Xb�|x�i�re�����3��{��R\,1�������A 4���Ĵ�)��C��is����~<||||'����������[���Q[`�
M�HA>l�SAI3�����Ǐ�������^�� (>$��u�
ih((5c)V�Rn�:���A��AHivlm��F�4j�h�(+cAA�@�UUE��e�m���kd�i��i�F6���(ӭ����F��BQZ�5�Ji�Ӥ���]Z��&�::t����e�յ���I���:�j�)�l�b+@hM!���)ttj��Mh(B�&����N6�F��CQhth�4��莈#�K�M:("��)��!�*��&��m�mI�E:�4ӱ���k�h�l��ߛ�L(�L��!�'�O��%a��MUh��p�����M`�:��KD�'6v�{|{�K.�5�Kƴ\�B�n�TG��w
J>P��6`-�oL068��)��H2��F�dA$6��M(R`�ȶ�mAD�`$CM�W�~?����p��뗸3�{eV�z�"ڑ���=Qo��k5W����~s��/F?����k�ֱ�^a>���>��u�j�NN@n�h�TW 3���z!�/�i���o���`0&|�[{�d^�5s�+���A���I���g9k/v��qC�njK$������e����=;���=���r����gݭ�~�Wܪ��!�3o*+�]?5���zYX׊��z1��E�T_���v4���ݏ{~�Xp���<ACƻO��2jɅ���2��P�,R%r���v�g�ow巶��׃��{_�1�H�A��1���p���Ǎo��1��*	^���$v���҆�=�����m^����m H8v!��˷�Α�
S+��u�.]�{]o3�[چ��ב\�	�q�a�/����NdW�|�- C��^�s��	e	�*���ku�^�.����4e�S����t���U�z�Õe��7;������xg|·��Y���tV��a�,s�Ŋ�
�fW<5Z�E�rč^��>�&�E���a�Ηo�x��{�6�C�I����̪R�꣪��C7d�/��coP�֟I6�b}D���ݜ� �DKgɷ�֚=�gɾjs��:���+Q(u��:�?�-#=���i�;��"��L��V���-냩lO.[Z�;��K���G_�|��������3���1�z����T��.��,(,��U~�X&���ʐIzjz�+߽u2�J�~��q$0v�q�F������д���=+^�T��%G0y�Q
S��vU3�s��Dt^S�l�����{ä0��y��0�,�>ó��E�j��e�Z�ԯ����&��ok���j������/�C��^��<<��C��o-sD��n�}kKJb*��*۰�19ص��%�r�c�D̉ �c>�t�g/�􁁡�ϢĽ'��N�y�1X��x@�-c�i�a ^E�Hݐ�9.m���;3S��b�@|<�[�I>9n�^���ž)P9b�(k��_���0�=��]�zRM����R&��gӶ�QaS��u�uG�ʜ,��me=���<��ݎ��h��@��ږƠ�H\�veK2�*8|�v�����g~n�J�|��b��88Ʊ�����v�2W�R�w��U�?h9!2��{����m4n�����s�t�]�{����0�B�Bـ��|��>y�����S���S��E[JK&����;--*�s�Q2l�:&:ɞ5�(�g)�7�3X�t�juoλ�^L-N���}�&�y�/f�%$d�G�P#��<��G�M�㾰!z�ǧ'A�Ύ��u�����|���U+oB�X7p�s�&'p"��.Jd�f���o0���Vu����q���O9HL%P���ǡ�l����Hql���'\�k�Ęrَ]`�۸�cE���{Y�2�:�Ju��)�=�cEL(>�s�{�[B}ab�k�����U3��6�o1z�K�R�6^�=}*�^ދ.�X*��X�����8��-�;��"+t<���Vbg�:���`�>1�۾���a��$YS�����rPX��0�ڋ�,p��E��Ղxp�wF2����^|ll�5�C�u^��Û9\��qTa��k���Dö��K�d����n�v���v@M �8~�^"5�Ha���u��Ϟ����Ȭ���Y�N�N��i��Ŝ���^��Z���K6VŰ}���?���GW�r�Ќ�jzsC�����}L;�KjK��l4Ƨ��)���t^��嘀^�;3��C�w���}�5v�v��n�h3��Y�2~���l��c��-���g���-�����y��k�+���;	�(aA���:����n�ws�f���w�>bI�l/�����I��(pRj�P��}����̯�` U�ď��6
-(_:�лt����h��"�+����=O���_�����;�1�o�X�5Wt�H���GJ�u,��Mv^��-v.�!�K�Yۗ��awzPRVp+H�V��˨�Sm��N��m�fP��P�TX�f��_�'��E`��斐��i�,�ץ�ލ�6�y},ӃzK��PAC���[�{r�k&��s7Fs���>�va��Zfb�X_hx|�p������3�Z|�*f���:�O���0S�C*�lj��pt6��:���
��˱Y_N���F~�1\�T���AUc
+y�����،es��=��ٖ#[���jY\��a��^=s�ș{fd���§+�L�%k��gsL�B�u�dm��j��/��bX�F�W�m�5^�h����~W���L+X���[f�Ac�vk�Lk�Ƒ�@���C�$�D�-�K	Mm~��8��M$��·�^��;��}��s`{Й���ۗf�)���ޕ)?x�&*��V��6�z�&Mb�c���ʘs /b���u�X�d1����W�����v~��yU�����E��1����~�:����V��`�3�`��J#��vC���遯4g���}luvIvN#�O��e�v�.��%n��Ũ	�?%�A�3��xwh�E���2Ϙ:�C��j�I�j�4�ˊ��n�t�.l���-CN8���Wj�Yo����6��h��˘/���N��x��	��1��0�Wuխ�N� �&r@��jU��wI�L��k�Yjh�3�^,�qvj?�^]���@?��Q��y�uǰ���o0�]���R����Q����*��zpE��Fm\�@UR3^�ٱ�1����Oo�������Z�
�ϔ�c�x^~m��B���,:�c�^�y���u�l���vӎ.�+t�K�n5�y�Ƀ,�Ad�!�3'ͳ#8gJN��8��^y��mv��u�o5���H��A!��S����V�r�"��Ԇ����8ėl���Aĭ+GW��/�XRK��ٿ߹�0��@����l'�A�0[���a�7��O�8ᮑ����F��͢%z�x��"f�5'�sͼ����E��=Ų/O͎�]��5[7Q{W��l�J�H8��!��%�CW�2o&�W����9�����Ƀ��a �Z�����+�P�^�<\iѕ=�m��jM�Ǧ�%�Վ�=�e�q�4;�2�)�?;�P�^;p=3!c�ѡ9N{���TT{�A2k�uUKZ0��*���p�Gl�i�
j������!|F
�Ӯ�V�0�<Rz�f�^y�gF㫬{E�T.WT\ȣ�~5�
�>�~�G���<��ʳ�7�)[hc�q������UVG�b���f��3U.�
���tq�1�wS{�[;s)N�{2�J��mE�rn^.����r�7a�uvqs�Gۼ{dx<<���o��{۽��8p�=�d���Tݩ��~��cH�Ir����;�q���+���2ۧ�{'�:�u�_<��$��m��5S���t�`��]����[�fٗ'F�VVn�R��L�7���3��gǧd0�mf�r�ڨ`(�c������EoI�Y*��礩�[�2���ld^�+�nMW=��a[����=L�����@,�S^��*���c63H�g�����\/��JacJ�v��R��L�&�ueq�z�1�٩�zY����=��=t'e���M�q��P�r�䍴;&��!�u�Q�K�Eu��v.F���b�F�3rf	屣�]m2n�9��n�D�U�ŷ��q�j�I�,nA1��M9��΁p4YJX��h��;�p�Ĥ"�-ѻ��}��$��%���
�5��&���=�C#$�=(kя�9↉�����-�A�s3
mڨ�p��b�$k%;�X����Ӳ�����Џ�;'7��g����|M���_tc��qF��N0 4&3c�죶�7G��`��v�r��k{(^�,Ȱ�{�.�T-�#�S_Jxp��b���W���n��_�^�U�g��C�l�SW]c6����\vQ�G�6��P�T�,YD;�t��,��N������8��I�X��^y�+Q��"7ni�.����s����n�H����g��T	���[�d> B�k���{ʶ��+�L�Է�O�&z��\�ә�g��lOy�r�{y�11�E��wSќ�{�E����3��M�IWA��e�K8���+���Ը�.��;�k�4�ֱ��ޒ�gK�)���P��t�ӭ�T"๔&纤�cu����z��7� ��t����y�7wD�E�k޸�W��1���r����#V��)���N���c&��)FKh��:�o��5Oj����h43��6ʘ����/U7D@�����.+xӼ�n/l+��4u�aB����z-��F�ch�At��9�m�hd[��e��R���u쇍U��(�i��o	����l�K�(^����	�ܑ���A��:Eot����������U>��s*����
�9���V�)�j�bk�f���ʖPU����rm�Qdl���]wSG��y��"�32c{�O�yyu�$�P
�̋���;�s��<���e���Kzr�v<��m�e9�݆�J��q�;":Cl{9��9�EBR2q��U޽7bd��d@��M�z�Pc�#y���1�롛WY��FV�_�0�~H�VHX�`�f�_%V�����Q>D�Ŏ��2�a嶛"��ot���r%,�{���tG�|IP��5z���#4�����U�w��'���ݺ����u���X��O���{�(�1�옽��껾`��3�#����+ �e��@�]�[2d����ZUc�gm�z:HٯJ����+��;��^M�9�*sJD�M�<��o�wsƹ��A��zn� V�2��(�75�U��O���k^歜�]�F���O�pd�Ԥn|�Y#��ĩ/��D�d;�j�w-G!��F~�愮���o�k�
�5�}�㰴�(���GJQ[w�X��s�573��*���7Ƃ�ޝ���&�<�"q�w��Z�-:��c�������/��;��ؚ��@�4i����gp����pE뭙��U/P��/)�z_^K��Љcq��nR��OS��d,�H1^�mR/y��$�$�M7�e�[p�V{z�qz̆�x�t��e�#��pkSsNCMB��0~0�m�N�9}kr�qAn��������(-hc�>�[}vDg*a���w6�N��n�n��:�+�0�wX�]��ǂ���������ѱٯ�Q���LA�1Q���S�N�LP�U�,(g�a[��eoQWӺ7Fuhd�Y��i�ۊ�J��ǩ���˺�������uq��h�/Q��}�Wn�D�ߛ�f��@Yg'��.�1�e\[��
��n�_�}E�n����݀�c�@h�y^�}q�*�mZ|�9B�9wtܳ�\@f�3T�烢�K�g�#�:M�l�Ξ�pT�N٧Z:sVe� x�%�"Ls��]�4[����brبD��>O좬�Պ2�f��t�S9��>�%Y� V������u�tj0K���0�e����z�Qey*��}pTx�DQ��Nb��a\;Y�WE�(��1i\On����h�oH�Η���f�ݩ��+0�{���!G���k��<���6�^�jz�=S��&W�2r�AJ�"��/%g�n�%F�_Kt�ݶ+쾍[1cO�^F��V"q*ɋ>�$�h��1�mI+����.n����c�3��썏��~(`۰�'����Zy�Y\��Dɫ�i��{&&��psԊ�����n�A���[�=�ղ)37�K���]��ڇ����;�wo;�&|�z�.T�[�́I!O���Kݍ"I!�n�{��6��Q��>���|�䒾y2$d����ϳ2<�u��h��v�j��6�t�9�v�zZ�
� -�ڌ��������֋(������_V�Z�/F�q�����U+�K�|0�R6��aj,6�uY~zs��XW�e��TBR#���^��7��Yܦ���6q�j%D,��gճq17�gG�o��ؤ^�U�&�N������<έD�J ��`���q&��Ê` ��5*�3��gE�7U㬒w��̽��(N�R�jlf���m]��Xd�9zt��>	E�1���� e��)"�<]wj��:c���ݐ9�b[���(l9X����} �UG9�*�V�ayt���#��²tb��k�ʎ�r��U9��7HмG�(���&0u^�ux�Ԯ�ǲ�Cq��j�[֏i2'19���'wb�+�.m؅óq�;����n��s$�'��2�6�	6e�"��qk���
��;T����+��u<o�ʽ�s�C�ǃok��D-}X��oi�#�l�}���0o�����W�Xδ0��'�ER��2����r��l��JS�&`��zo-��� ������O(��:"���O]n��i�ց�Y+ڣ����H\I��I�'�Hk����((�Ut�7Lڳ�ov��F��),���<�λ"V�bx5��t�ޥ�yxF�_����E�h�[\
	�й:I�@nuvI��^�꾼i� �:���CMK��t-�=W�L��'�u^�|ȲR�&�ޘ�X�w�}���|�6�]lc��t!�)�'5ܱ��YJ��1x�,n�L�FT�BgTu�~�앥�!�G.n�Gaɦ�+h"�b����ua�g4Ἥ�Η%��Ѱ�0R��:�k�p�»g���퐽�ux�榍޲u�=��AxF$��a�����\b�p)�`�lN��:�ǁn���~��<;]ƀ�f^Lx���9ueu�T��i��ǡ��<��<	R^b�اvQ��;);R��<&,�Υ�r�ⷭ��6bSVm�7�#��zӨs>�*,���D2�}}��4��v;�}(����wP�abI��OQ}�57peh6�Lm&���}�=���(f�zRF�=������Ǵ���"�:h����yVoiS�Y&�Q70����-���W�e��:g�e�t��-B�_�7������:����9�����H���H*.l`/�8)/�M���@����vv���������-b������������e��k��6�خ��xK�.�J��Z�CY����q17%�b�"�
�p���X�tP��YYq`����X)�r�A(�J�C4﫸TG�
���B�n�hn�,����kUwJ���gr)�u�J�F�t��\��st�;'�BV-��:ˬ�l*P�ajy��xr;[�Q�{�MB���**8��m/�B��a~n3��Q�q�$��Q�4�n�p�V����M��+����V[�[Ǥ���������4F�+���n��uՆ"ǲL�n;s[�����"�<�p+�����ŧn�\e�ڔx��L/����3c8�7�c������m*����@џ�I?������li���5��������j�M�k3�ߏo���������������>�GڃAA�cRN�"֖������1RSA3��׷�<||||~?_��C�e*"��b"���m�Ψ��h���%.�6��
��[V
V�k@j!��6J������Mz��w���؋S��]���(����im�@DA4�DMS;8���
it��Z%R���*�ѡ4h)��E�M&��֘��u�HPUuV��"H����E��u]41���AU]���h�$�i���"��4�h�1UA�ED�E,���iS��;�4""ӡ���bӪ����h*�i��6ƱSMD�� Q)��@${��9N�6�)r��!+��qX����♽��.[N����KiLjj�YBd�0-Ik�9�=ݰ�0aT?{���q^Kd���6�K��3��?I0�F�n��h�#z�@�.�w+�j��Lv[�s۹��{7Zb��ѽ�����<Cp,�������8�ڻ9�[l�{=E����:,�����7>&#�WN�~�,�&"�G!(b}iy�;V�x��g^��5g0b���\<;���Q�y~���,�cZ�f
5�Vwr���|�x���T=q�'�(��x����$��N�e�|wJZ��'C�}�<r)����o�x�F�m�3[>�Eu��+0����d�=ױ�����f�1�%TK���Gz�XS�9n%�& �۴%@��E��������q��{:�x�,R�u�;W"��Ϫ����Y7!���U���z�k�������e(�)��F�����ɭi�M3��gF.���-����m����j�N�y�H�;9Ғ,�w�OO)�{<�N�c�Gfm��MB>έX8E�B��)�A�'p���n�^�.��͛���+��zTOi�X�soW˕??�|��>���۶��t�i,�U�*�v�*3i:�e��9�K�HlC�IW)[8�{�H���������^�P�<�v�}����$�'s�zO�W�ժ���MQ�Eih�l�\�ԊLf���gX���"������0���#���C����@��4,��+^t��3���Q��(�Ԁ�����1O�*;lګ���ǝʑ����յ4�KȮ3s��ɍ�ӵ���N=�q�6�M0�iCz<�y�ޱ�UP���4���Q�_w3�����үEk ��*�yS��s��do��0�g��}痧�����VC�p<%\W4��Cv+��*r����X�?e"���>Pyf_�/w��ЍNl�۱��$^����6�s�{�_hfަ���p諎�L�5/!���B-)� ^�Gq#x��|i�U���w�y���S��Jv)̌�q��]�(�zw�ɪ���f*~��	�� l�����<����;�}���c�<�(v�V?��%Ys���u�����i���$o2\���U��T&�q�Ʒ<l��It�e�c�����$upTY�� �9M)	�������T y�q4���+9�~�F��u�X�Y�IYx���s;���t��T�����xxx{�V:�HƸ�}�{{I�1�ęDC%�i%����:�l��@��#6�����a�X7�ҫ�EE�GV����ԭ�ͯ��\B��R�O�^=y>��3B�ޞ��#{&'�;�Âȍ�ժ}p�u�*���F��>Tf|��a4��1=�]
��h\5K�Y�"�B*w������8�ĩ��PL�tZ:-��i�'y�C��;콙�O �$�̦�"��7�%������jǫ�4��\�קx�C6� �Ð�c��l���f5�S��m��sΎ5ټ�e��T�Xe��Z�>�>�n����Z�u���Ū��|햳�\�vr����q׮IG �t�Ƃ���kC4�q���N�z�7?f`ч�DϢ;_T�tu��R�1^4�*��6�C1mq|���#�?K�5@a��F�a����SYC�u9�����UVU�gM����+#��9�����*s[�۳�v{m)JXؗq-d13�s�|��C�5ta!	ƚ�^�M�X����(>���=���B'Y�J�X{]������`��Zi�:����Y��Q�N>C4�
	)�ٍa{c���6FQY��c-���o�w�H�5��.��2�,����"�f��|���I���v-��;�ޭv�]�7t�F�����sNc0Q�Ю�:|�������,tU��j�QQ��0��N��>�� �����΁��}xI@��l�ɍ�1�<�vn%yf;���ۮye��:(X1x{u��ö�;U1�7p���-�D������:�a|��^�+ �3e/W���Gs;wK�:qw0��+��S`���"�S��1s��m��ړEv�L�������=�����[��e�X�fS�~���]��,���b"Y�zVu��fý��cs�����O1�z ��p��Z����+r�+rF��t����G)x�R\�Px�گm[��-�B��!v����[_�ْ���B����c���W�&B\FN�j�3��@�On˝�����ٯ�Q{���p-=��N��]MT�s�/iD��+X�;#�ɻ�.'���"�$��t��}4R�OL�ۻ-Ի�(}Vs��G��*�r���zg��ָ�nS�y�b7r��MOM�k@;̛�V�Y�0�C��.,Ea���ڼ��U�u�����'�`_���I�|��
�x����OUuy�E%A�i��<�Sۧ�p�箸�����U(��t�]݄���˟D���ox�UͶ�M�l�<����{�<.��:�yr!gO�S���#�c�����m�#6�o���� �4�ҽ�5��A��Ƨ��&��3�h�#��+��[#g��̎�уy�*p����Uc��Ƽ�2Ϫ��C;Q�˦��b������pop,�.���9�S�R�hܼW��7�@�� �z�\{,��O5���`��6�z+�{7
����3cTXzE�W��<��w�3m�v�	�'�Iy4+o�%V�5�g���.k$����i�h�Bս%�������\v|�6��v;]�(�%�rz3e2�,2��-��}C8����Љ���Z��
�o���Θ�g�8J��;Xq�W�\���;��u�S��F�L��Q����㇑�_�z	�N�rN��ؐ`�y��̺���"pw}�-�K�ne���<;����oVmⒻ�&G,���*cCq36�G�R}bVW���t��A�}Y�7���M�F>����C2�F�ƛ�SsNdl��OA�GO��I�"���d�6�x՜KVXܯo$�(J6�ڹ��3�p���y{��kp>B/���7Z"k���E���!HauR�%U �W;L���5]ݾ8��gU��h�йm!�#�[|g�Ғ�Y���'7�}��.�jn�������/P��b���=��$*�*+�@͞J�%���X�&��30�]�3G�@��f�I�����[zt�p��~d��^����t^�����-�׬F[UK���j���3���2��(�km����cp�w*FOwm�s��8R�r�[��gv���y����鴼h+`�g��0�`��D�v@�L��d%���ϵ|�ݲ�����D���ә��b���o�<9Qy�y2K���k[^�x!Z�@�����M�u���r��:lܓ��|�l�D�6��m��9�䦫��6pc��A/.��G,�e�Z����a�9a�N,���zi�=�3�;�W�W
����x,)��@��Ԁ�x��v�8�w{�)+9�Jepl JO��� R8K��rh�/�$v�.������H����Ϳx��H��e�� )�M�L���iՕ?*?�� �e����1�o6�s�N˥]o���DA�!��b9V`<+.���e����$H��/�d��v|=�o=�)N�9�j!�����������uWҍ�s�t]���H'o�j��k�b�K�])�!�s�N�H�~f쇗�ɪkL�m�y^��$'��M�El�X L��-@�p~����J/�b6�Q�:|��}�{�s�;�[\�R�H㸨��.i�Ƶ��|˚��W�.���F�]�� og�VB��.�2�x�)GC38�5�1�>57�u���vfȵn�U��s�tV�y�\-#]#���;�<u��E1����2�����3�U��uә��ǝ!�,�Ղ������1�G��3�Db���A�m0a��XG�~���.��4�1O���LXژ#�~�R�܎���h�+;��wsF�&�fu�Q/��O~Ε�T��W,e﹯Hwqx�7��p�����cR�[�+y"��].���Wn.�f�5�+R﹵<v�h�۬c�;���d����Åb�߿xxW��75��O��r�֏U����4�ϳ�v}�gq�E���k���`��L��+D�9^����9=W�d
�\��K�uci�kױ4AO��U�l�{�]��4Y/��X�F����sy)��`��*��H����e��X{Y�E�W�XԆ�pQ�F�z��n���Vr�����y��_5�,ڱ���c��� '�A�o�n3� ~�\,ͳ�|��g,9k�1�ѹ""k�`�u�%��'��I�3��=�x���=N�k
C>WP�'i�ɭ��L�z�+���ḁsц6�[��<�tQ��9����h����Y�30�msC�k�z6�h[�bt��O�k>��[�#E�
UY����]X˧X��CFL=�*�M]W�3���;�J���\�T:�v��N�Q����j\��ϣ@P�U=@D���L\�K{=�jM�w;.Ot��@���n%�NމfP@�Q��v>%��=�����_{,x���y�Z�w���f=hu�۵󮗺��F,�
���Bx��2>�܉����`���0���	�%�[q�H̫�b����C�h��:�ݴE;4\���Cª^�ߙ�5��~�uO��������;���k�+�s��:�_T�Np�ϻz�7זs��U@���OL��HO�9P�G�x5�@�ͺ[��91g%�gomK,�E�)&<g�H�� Vy$.�)bKu����I�Z*�@Ӛ�#��ٱ���%|�e.2+g�T�@̼q9��6�i�vOKi�������
�&��h���T�6ڎ-�?p&L<M���Gv����Ę���������]b��Q��]P���+�h�����Wq�L���ލ�d����wr��m[�"
~$�T��\� �	���K'�zs����|�"t�򽎖�̀�\0+�Gb�/M%F�E���q�o]/c��UD���7�|L[#g��}������)��NT�m�+��ѝ�N���"���˫+�b��d���7��ۣflm�3(v����+"�Mf����XA�)�n���?kb�]g׹��=PPR�Ҧq��վxLj�,V��t�H�[��+y�[�M�a����[�3��"였��n�mw
喯�.L���� �� ���,Ф�U}��z�F���Z���R����|�hI@<RU��v/-��d�QL�C�3れ�Z`��M(�s���K��7�u�:��#~߱}���J��,�Dǉ��0�.r)�S�K��mP��l�� ��܌L�ADf�%B6��7�r���1���WDW����!�k1 �y]#���=�$�po�1�5O�D�����% $Rs���?/5(�����ƟY��ȧ]�EPF���ǓkP.���d��>	����s�$Ғ!b�J{$��U͹�U��C�{��16��'���խe��A���}|zy�S��%+RU_�/ۏ#i��?�Y�퉺~���~����V��G.�#k�l$P/	V)����vml܌jd��uM�f�7S��7�u@~I�:��E�Q\Zl�Wʗx�1P��?��u��
���}]�}��n�2m�� ��V�zMYM�G5��P�!�i�1Uo=sxrc�l�W`S����+l!���$��;�6ԑک���x����-gj���{g�w�a�ׄ<j*b�"�|.�<1���S�A^�;��Q��<�j�6�DB�y��/7��}�[���#˒,qh���{Ucٜ"�E˶�w>xtv��&v��Nc�����i�N*,a��|:Ae�+`#��K9i�b��j�c���-H��|����M\npZ%AǨ����ӭO���v$U���]����.�T��d.Sb�ٌ#wW*�YǅKc��J����ip�
)���fWn���ðL�l<-_" �"ګ��19�N�0i[G��BX��s5n��j�Ť�s�`��B_Aݵ�Q �*�u�-'3U�B��.�:Rn���@��.pȊ\g���H]�mu�ͼÌ�i���K�"�;�؇�i�ɔ+r��%e�'c�k^�����ܦe���J��ݫ�X\yY�I"Rd�����]ۈ�b̩[�+R�zu���jPI��1\�;jO"35�5K^u(j��MJ���Gd��قmn��q*4���p���^s�z3�s�n6.�cy���+����`�Fmp��ϩL"blsl�����ע�؇�q�˳��_�*{��FM5�s�!�o0I�%��8�NW�����l��V�T�4u��NT��@�&�׊V<�������p��<>�_{�<�d��ט��H0�Y^r�Pi�}����b�k�������T���'N�7����j'V]���[۬1�R�D��y35T�S�s��y^��4��b�}��N�
J�i����0��>ug}��;�v��4��L��_\�Ј��[>��0������T��]��|9����lL�*�KӄlD���q�tyu��>y�SR�F�.��t�6o��o���f�o.�A�/d�;ZR��:	������f*���t�n��ݝ;��4�˗�[�Ն��#����6Sic�a�}��XIe������륆֣L�|�y��I���BZ��VLY6�4c�P�'�:�z��n�*^V<T�6�t'��
)ƵZ!�폇8\v�<�X�h��0�л4bĚɵpsw���d�piښ:���؎�q]j˥�D�9\4l��;��Ȯ�c��������
]\X�-d���$x�}�1fe�ZDO.F�8��ʂ�L�bä�� �"�t�f�f� ���3��ْ_�''j��0��Rl*q�d�.��3���j�ƍ�h�	F^���Eeҡv��H7����(�����:��.� �b[j�W\����d+�B�fd����'�����Y�H�<2��z��"Զ7�zf�tZ���m%b'�b�zr�fpً���}6�����n��߯^�>��)�;��Z��le�;`(��z�d�ة��Π�J��9ϧ�������~?���~?����T��0AG�Zt�;��㣽cSl芼Ƣ�'�����}�~?������x�y��Z�ٝ:��f��=X٫��-F룪K�ˍ�Uv)�e(����((���5MEQQ4u[$H�T�Ur:��6Lԕ`tPb"
((���������ѥ�C�5�I��I�!�"�������X�I�+mEE4Q5Z6ɢ�F6رUFؤ������&����W��MS��;m�U�l�DHRTQUP���Q�;htf���b��������Fv���0DHE���M4�S��QQu�1,@[4�tTk��*��E��Eۏ		�d�N��D$�����3{tv�U��_=sw%���❞�[B.w<�Wf:t�=J��޼ҢbR6;H��{�6��A�:�WVpR���D�?��/�#
	8Ѝ�#Q$m��L�X?�-��Jq�#�*���@"��{��0weE�I9��s���ĶK{i�3k�ZD�\_�#=��P`��k1o s��^17ۘ��y���9���&������tڎ��QW�s*��.Lҭ�|ww�y�`��A��l�n��o%�Eq^T�O#�7���f��?���Tn�.�h��0g:��m����^ŗ��;Zz�P!��w��&�v��M�\�0l���M����P�{�SL�w[k��=3���BAa�Ѷ��9n�T=�Hv��A�k���`& xVhE�9� ^�DX�C0���6�o7�[����d��*�)��S=x��`�LG����!�ӒM�:2�z�փ9�f^D���JП"^*�N�9��B�6>]Oc�z�V\K�=���)��s;0���y�;d*(��!ܕ�(�nm7���Q��ͬ:]����y�7���ń���5�"�3p����-�rAJ��w׃uE���.�}u6�}N0d;��7s栶)p;#�iʼ�+Ώ��N+�\�>��=��\ox��������u�\W�*vl���^��;\EN=o��s�X�i�R �F�R&p��e�Gs`G3��۔�u�T5���]n�ܤ�.d�����+�̓�&��/hʊ�at��8��|���*�J4
R��^T��Q�-wo���uqurU�U��o8
:+m�u��d�?����M�g �w_7�p�4*�Ϟ��n�\�HC�Q���ۯZ����{;�Q�gsME�kv�מ㫸�3�� ��hK�J�����8�;�i{ɺ���TP�K��[��{ew7z�R�d�n��:h�!�"#vF�O_��$b�v�S�BDD����f��Y�g��2P��<�(���2�B�z�X�T������T��0em0M����&rAX��K�L�|��q�8o0H�m�X��:�l�Ш� ��	���]��T���쑒6�lo�|��؍@Y�93yP��cI�l��n�ײ�7^�c��lχPc�g��^��*�Ȯp��W]WNd�8�g�\�����m
�&�Z4�2���?P�oXt\���w�y��U���}��j��� L�����5�n�E�Ӕ�c��e�tBq���.^y��`�:vD�����1C���A�f��x��Z;wA�l�߼<=kv��7��:��6Z��:Gp�>���E�c�g���f��Z���X%�x�!�ׯ^_Gr�{����{uA56�_���"�e�]辿J#/i�߈I���z�-Y#H� �J����{�v���Pk�7Z+D�����k�� U=Wz���o�b�r[@vH��p����:���˱z�u����S��������ҲѬ�}Ե-��e&����r�LIs:��G�'���8@��BA�+�f��V��Ͳ��6޼�vw�3ᮒE�))sƫ�v�n[���׸bSC a�\�f�5��>�^��@��-�Ip/�.h:).4�]>j�7EX=p��4^���u�Èს�:DpحR��Ţ�J��W��.mi�W�/F\��|g�����vǘ,-�\�%�.�!tW��U+����mV}c��0�8�I#K3��Kc������\vb?m>o,P�1|r���k���r����%�la�m,NK�}Hڇ ����rS��c��N���C���Y�W��&Zj��E�Ez�=ů�/P����,�;�3��w��o7C<��ol��K��s�t���S�]�{���>`���W�
�L����^kˋ�̺�ㇶ�����(J�T��`�l��a��t�b�[��\JfU��������s�:r���IOj�"h���R��S�A�ܯ�ͯ�uӾ����#�C���Y��%�t�{L\�oa���c��&������O4v	cbT�f�j�������<4ɑō�%.�}P�~+n�l���?2�V?Y^�]O�c]qV����|3q�^�Im��7E���X[^�2��X��V��yY�=%"�n+�f׵��"2��y,�l��s7�}�m����]reV�빠�=ܚ��:�(K�7��!�w���71v��UW WcM�)��9����Ӟ��u���e���Ξ� ���%{{w�&#8���)*�x����ս�@~�ѽ�۠��d����Z^�!��uI)���A�	�eT�+\��h��8��.1��ή����ne�5M]�)�I� ��j¯U=�b�ln��]
��z��Yv�v�b0N&6O_5 ���eh],�p	K*ѼM�k��RKy����?�}_�L��w�o�#�?�;lP�4T�fݤ
g���s����'�˧�>��Ĕ�)08}�$�� �O�ӳ�z��vb}\�}���9JD�b6���zRV�U�x�v�{}�<�Nܻ2T�����}��b�����\+�Fl�YHQg�DK��z����>e��7۲;��mh �,�շ��2t�g�U	v�cnƬ���W�6z}��&W/('�)�kl0�� ?��fC2��B��h��\FO-��mqE�԰���6�A��Ά�M�.���Q�#���Jb7_a[��P�+k�QAQ���R}/z�ty
���o1�e�y{G8/�'�#T�q��h?-��o)��<W�m�wa�M;U����D�g�꜌�/���i��A0�f`+��dޣ�Ǧ@��ޜ�ͮ]��5���'�Zn���h�ަ����`����*-m�/�����®̶��̆*����3�Ƕ�oz�۶g�ʐ�>�z�y,'�{��z��e��EmK<�3�ȷ�[�l��&�=�Xt*�Pl_�����8B���d��,�|�/��H�#F�&�hp�˴a���Ŏ������=3n���h{�����f�׆oɎ {�`�>ا�� WH�.`���W��-���t65����;\
��Һ��/5+F�^�!V9�k��h1���}�v���΀���Z0��*����Z$D���}֨e��NЋ]nj�����h@n��s�d蹌\B��$����qJ�Qz�<��zk	Y3Dd�܊mMV��s�qp�Y�ܥp'�є�����K�wvmT\k��Վg�l�u~�t!��QZ�6�Y�h�j�����ݖ���%�z�*�$US�Ǻ���x�:A�!�8��@����s#8!�/��k"��x��j��2�}�=�Wp=fC_���A��P�ZZ�sD���������-�����r��@�Z�"3��%��U�!�/}���y�:~u��)����|����7��(�{�cB~H��C{W�Ȇ�mJ낟�ӥ��v��4/�ފ�w�z[�*1�+�NS�;v�m\.�*�� H�M�%��-d�Y�hf,U�Ao��g
�ƜI��c��ʲ��t��L�\�R�uNTa�^d`kPc^�]��^Ge�l>\m�?������<�Z�iL��w@s�b1>������Γ�ԷLOs��ùg��s���JM0p3�Flpއ	6�ҧ�=�ٔ5�P9���6�9=u����uP����P}�o�����r�T'�.�Ĭv����1z�>���/p�7��-פ�O�ٞ��=̭V��Y�4�m�>����ݺ�@����&>%o7B��/����ǟ�Fz�㷢k�m�n�T�Q��ǧ_�u����#"�ח�#���I�x喤��Տ��'�i6��t��ʥ�ѯ !w�ɨ��������}~ �Wc;,F���,߸�99����=<W���~5��G��z�l��+��a'^���w��F���r����q��➡���麉s7���,��@w�Yh����}�N�e����VwY���[��$Ʃ�^tKКg@�?X����*��ʠR�;��תc�e^�$,�t|Fk�G��>�S�_%h}��3��iϥb'҅)���\�� �L"�����y�om	n#��[����u���r��,L�.�s���K�9���\�Hi��S�����xx{Nl������1�»�^�r�1�h�0rM0K6=�
��q(����x�n汣�3�d��?#�R#G@�b m��H��%�B\d6=b���lەѷuټ�X) 딁\8e9\�l��_���[ʀ�#Q����і���mll����n7�CN�r�`�^�]���оJ��1���M)�R�5M��2�ٮ���Fe�i��T0�^|�����ޯD>�&J�k��jۯ����흼Ԃ��5+v@W�:Xm�<3Y��w�|��t�7l{<v��N��:؋���܁�Vq�|��m��??��G6ݨ�j�3���������8�����R�g$i�W���_����vY�A�Ʋ���Xn�V��s�!�P��_���`��D��&|8��]�2����Wx��ۜ,��Du��"��c�2
F�1�E���ѱ���a�<�4�J�]���Ϋ�.u�Q��\��E)�l�j#Nu<�ՎMv�z�P-�;�])�R��~�W��콺O%u���� J��Bʥ��乽�1d�){k� ���-�:.��a���13`fY�JAîev���|4q�j�<�����v���Myw���4�3_n���Ɖȼ����ؔ5����x�Z��������d0��p������u�[}�B�7���ܚE�)����P�A&��Z���[<�FՆ&۷�]�IJV�:��vJ�l��)��26Y��4/%���ƌ�җM�(�P���r��AYK=��&M쐶�EM9��)S]��3&D���m�C���h�SlP�dw���d0���fT\�U=�wO�����8L��ٛ7Lbo��X�#&���m���)+/���T<����9�ۆY��>۪��t�ә^�{�p�uN��Eqlx��M�ٌ��r��OZCv��n�Qu����X��A{���t5�8����<�F��a�7�����p�ν�������#��W[>�sY����O�M�:� :w578��d���8�G��H�8�`�)O]�!��7�:��\Ub�u�w�y���L�V��-�vs�K,n���9qT��}޴���:�=�&ׅc��аGw�����tl�[MG���ȳI�,W�Nm� �q��	u�R�]�sI���/�7���j�{�]�����[9�ܝ�N���
Q�:}�Dl��]^�KhMEFbڥ�2�#hlc5y�;m]wi�R�W�8���C�]02�/�S���v+���%��0��:�Z~ȚZۍW�F���`bm��`>٘
�{,�^��;>����}��禮.�::+���m�F.�>���c�@��F<��nq[F!��������	����	r"x���w'�+�].���|+�˪�hb�򰴺�<���;z��m��[��%']��/oB�Z���xQ�����uk�-�<k�H�j�/
nex�CEZ$������K����~4�5����m��d�����s>�\B��Ԃ�n3�р�g@s�U/�[�3k���~���z�uȃ�<�T��n�j,:�')8g�j��ʄvn��2LO�LMn��T/�ف�HP�`ڝ�����\�i\�f�`����3��,���R+xOnh`����"EU�'�sE�t!S��0ĕ�8wYV�yL� �bRӲ-NP�۷��̕�(pR���o�^����*P�Ҷ$~�b�M���y���ݽ�lSΰk���A�����	��k>w��,�W`�9'G�Op%�Ct�ڗ�,v������}s�%���PB��u�7�R��u_A����ي�����0e��!�{�\�4��z��FG�M�O`�^�����2���Q��+����u���<�P,��'˸��W,�[�u#/3N�l�4��T�����+�����rB9��U�{5A��f�z^��{Mvn�ͺ��F����.LWx�z�s��֌U�He�4���T߷hw��6�
��|� ]�Nm5���M����@;��T���4J/b�r��.��_v]lъ��M�
�k��2�լ]ũ�k��wr�i��#&Ӕ~��ː�衶���V>Q���l�k��1:����R�T�m��t�͖e�����J�Sk%�*��X/��tk��q��=����I�eY�rU根��v٘��┱w���3C�R�@P�8��k��f\s2�w5a�4���U��u�B(��&n˃���,R�+q��m��h�u��E��l��6�VC���X,T!:��Y�Q܉XN�ZRm�U:���&��������7�PuK� 9u�$	^���I���\����5V�U�'�SK1�oSdiIl�F���i#dB��4�҆�G�@<jT�ֵ���쟚�hWm7:%�W\&6GW_7.�V�.����::et����2K�k)�Qj�4��(Vj����BL�oH9��ڔz�B$l}R��|��Bn��5�|3l,���F��WjD�l�a��5����7�$.�G�[H	\����^龺N�Wv�P`ܥW�i��rH������Fq��rř����݉]�u�ן����Y�}��
ۤ	�8�nLCX��Z��]@�^M@�#�lM#P���u���7������S^�q��tEowUڃ���mT��,�JgLF��L�����}�/cN��n.�q+��`��m
ݮ,���4�]3�|@��z:ݨj�h^��|�ƚ��(�+et��}��������Ǭ��]C���*C[����"���.��䲹=�hz��3�tmu��^���*����#�Tb9rÔwo�ǵ��4o��#��rr���5m���ԏX��;k%IZ}D#�5n�ɊB���i������k3F\E�½�g6��1֕�u���m�=���ϮR�Nwm]�|v�P`e��J�*��P�w8R����C�EQE�����E%2QQ$HUEDQZh1�m�s����}�?��������>�-PG��E$MM�1MR�lUEEh1Q������x�~?������~��U�޺�6QMAAQVک���m50�Ҙ5Z��Puj�֢b�N���F��d���Ʈ��d�MTE[Q��ֶ�N�5AD:4�T�>���P�)��E�i��X�T�b���խUQk1M$E�)������kmT5MPh�N�6��3APUUA�C��XRMS�"��u�IU��b
��#պ����f*(�*hi�����[QQ5�$ѣPUMRSDSQA60T�]��u����!QTQ�QD�TA2ATK������NfdY��8z�V�8�;{���/�#:Ȃ$ov!B��\j޵R�'B�9�ռF`�ڜ�]s�!�������2NNn˘Ž����z��� J�IM�}t�}�7����M��x�K�TFT�F�_^���h� �ނ�2�#^z@㫨��������*�y�S���$�	<��#�l�jj�Th�K�S���[;aU֙�Tu�����kA�8���S���������W<��b�]�%���w��|Y�u��4�K�������θ�F'�=�u[�0
�._�Z��Wh����pv�����=�s_�u��7O����끶i[\��9�s����=�բ1xv8����$d��w�=����t�EV;��X��+f��%��ѝ�N�M�=LvUŻ	~9G�_�9�C�fO�"zi*f\*g��h�箱/��$Ѕ��;yQw��CN_OOx:�[�6���}���2�;)mF��������H��G�/���G��VW�=k=X�D,�)�����ۍ��v��c�*+�/�Oy`�5��\�6�����!�yr<��o;-,S��_+gJO�m��gU�F�)a�o�1X���uwFV�2&�E����^K<8�:�w�9j�ՙ��<�����3E� ����O��=��RVž����ٗ��#B(
��̀��� �詉��9���ٗ��{��M������R9z��lZ������k���o���<\�T�bЬ� mp^T�d���z��ө�� ÿ��W�����\�a�d�ގWW����䌊&MxΪ����Oi�ڴ�����S�L����E�0��|�ٴ5�HG�⒗$�;�������z&'��q�v�ßV��#��n��H��%�|
�/x'��kP�}m�UY��-�s�Sm��
���{��GWl,ū���+�U��aw�wf/;=��}��Wk�t���ir
�~�W��o%OYy��ee�H�.�$�=�׶�s�XOt�-��^T�kT0���սQ5C+(����nS�{x�ܺ�yIgr���={�C	�`�W�{��B�ʂ�_�g����W+��ji~�)��R����q�Ϲ�64��*2�(�<7����_/!�*`R��N;��&(���Ͼ�u�4�
nQ�P汕ӌq�V����֡'���=�i�DT�]�sn ��W\�u���@�e\x����P�S�˧��w���3���~������y����kw�|�wM�NM�ӫ8�J>
�{lm{����#ho��-5V��;öt&�<���m@�����C�+K�nwa��Lh7s9���6m���h!C��#T<d}+�YH��Z��5���������pѭ�5Z����C8 ��f¢�h��^[��S4���[K1�=�j1��&%����@�>^_���3��ں�y�	�L�8C�$�g7�� ��Q�$��yJ}ў����,u�	q�wEZ�k����y���rLLd�Ƕ��KN�HWf|Wc^J��9�Qz1��Bj�I��ͱ�z�V/=F�Ļ&#8��4��zX�(�õhM�@�}
Y���+�y��W4��������,j�$���,���Ĕ�����c��������{��M��x
������"o�Iɳ�ҧ�ONewK��7P�y�qha�'p���Ud��	s��қu��ef�N����xxgϪ�=	˃��lv�!ѤU�&�}|��o�)���a���ݤ����>rImc\x=�ݧr1NPC]���}�Ncs*�+yv�-�R�����C����f�]�1����6zx�T�]:�3=�����u��'=�H�.��Z��k�]���
�ͩ�r�i0c=>��#��X��jA	n
�T���d����A��w����hI�
+^F�:�"d./����»	�h��ې'��r�C>���8�|����jڡ���c���0:��UQ�c�}�@���(�ޘ�O��>�p������.nv�sz���N6E��i��y"�9��s���F`e���M�7�j��x�ת̘��2Hl��U�scݴ#�6��9�h� �m����i~��q�Z��I�6����ޯ��gݢ�z�8�g�сxVL�v��u�ɤ0���&����o��_�%��#����s��u������B],R��Gp^��z��woG|�M1|�����Գv�Oi=A+BQ/��;�D��Ak@߰�H����+^��{�ك컷�ط�������P/w�H�~�"�z��{���r�L�c��w(�pF��e��VFޝ�g~�<��KS�/*T��ӣ���ճ�oc����l�E�^��q�%:��g�ۊl-��h��������[+��+����Ү�Ŏp�[���/䄎�8�D�Ƶ~}�5+ղ�[g��?��ͽ���c�׻�Sdй�\B�H�f6{P�ۈj���3���ݳ9v��^H��R*��W�u� .�i�p�coC0m��湒b:�fu���R���=[�V�@��< �5B��jq�£��
]�2�g��5�z�B�T뤫�P%Q�����N�i@6�&��.u���;t��K��*.�tަ��)+�q�k�O\z��َ�6jA'��<Lv�,&�3�G�ub�4V���R�l��hp���.��U�
�-����j-��ȁ��!l����5�_ErF9h��"�����n߻n�]� s������O��q��N��v�:`�Mpf�]܇zd·��q~�������JVHL�<���7�z6�ԯ߹s��Mk�Q�C��{�+8�cTUd�%�=��&���V����B�Y�����Bo�����M�)�Ã�#����]t�`�:7%�b����Ν�W?_��Q��_H��ݛee���R�N�k�wTѱ�:��jm�s��u �.����I�~�^zN+����L�e{�u9���>���a�n��ɺ�kU捋�ݎ��lj��i��䴱�\[�I��v̎��:B]�4e�b�(����^��=W�s|�R�f���Η���x�H\-(�S�Zb�*�h���g��0�&�a��?�i��^_)%޴Eɽn�kn/2��1��ܧ�Y�C��'CXU3�,�b9蚺���;H��{"D_>��V��-��
��O��:�!?�YŃA*��D�<L��Yh��Ӭ�C�v��8�1��]�6��]� �G�D����p�;��h�4���-1���d��M/�H�jW���IZP��t��4�馔_g-C�^C����#M�,�o�Mw�E�ٍ���;�O^I)�j�-�!��uą7v"�'6H�Z ���4F`�m���(߹�J���Ҍ��-�GST�i�yҴ��uNgH ��� M5���ޚ��Y�]�����Ðƺx��Gb��E����z�r�]�[c�s��SV�-*�趞S'r�]\��bΔ�˾�.i���NS�k� -nH`��� �k��{�n��~?�걡V5�UZ}�g���9f �n��3c&��T�F�c%�mi���,WO|�i����*�J7�|�{��Y����OHa�a��~�E�?������=x��gI_���!���/5ו�4]�0���(g��g�k��d� j�Q�;[����I��vz��5�7 z�oT��M	[��_���m���׌[T����l1�Q+=ƽ(�v�&��{�Z���>���ٙ�YY�ۧOct˞�=�`����¸(�C8�@2�`s�����frv>ke醈�2��y̎&��l<e�]��e�k�d�;��+�ڸ�f�]�6r�7���2E��Q��F����R�.��^ީ��yn6sK0Q�d�u���.g�Y�8�,�JAJ���g���5���H���H�l�! �Mq�d�ژ���S��8����w�8���pjL~o㘰V¯�F!���/3i��}��Mf�θ��c�&��1���u�1R6-���Å�{�������A��[��6m.ʸ�P��6�ն��2���8iA��6^��s�h�n�r꽌伕ʠZ��<V��h%@��<=�\���;��o��xQ��{t��� �UِWc^]��T�j��]w;�9e���8��u�` $�1 g���%K�S�.�.�9�"�*ڈ�=�f�%ҫ�<!��6������9�R4��d�վ�ؽ������f�3��R9�O>ֽ��Z���y0Ʉ�؋��ȨZǮ�E���tF<oP�=<x���R�}�z���
\f\�ġPw�6T�v��Wm�8��*�Y�w��l��[�0-��kt�2������i�ޘ�gBp�K��dՔ�EkΚ:�� ./�c=����/���
�M�hX�_C��Q��=�@v��Qy���;�mv�=t���Tvp��U4WV�z�}v���q���8;��ceK��V�[EQy�1���L;�����f6_o����T*}W2�o��p�'��z�֫"�������<C
�PS�6xF�#��w��W��*M�T��,� 5��S�%�X����[�=v���ܬ�Nj�׭�
�����t�U��n�>�i��\��sL��Ԅ;5�JR�-ȦI�ޘ��Ώlъѷ0�ӑ���Ѥ����Y�������s~��O{u��wOi�:C��4���>ّ�
�=_�&�f�u�>|��t��᝟p��7�n@v�����vt;�6�����l�`w��4c���^ډ�$O0{�;y~���K�K\�����m��,9��O����W]��y+A��Q*2^+[!����n����U�8tG��j�^:;n�rB}׾�A��F'xif��=�k���^ղu�-�����w�#2�a�1��X���mh/��)q'��:�B����������9q.o�U4#��]�3Z������ȋj��w�o��k�q�h�R���Y��O�����/�1���,(���6�v�&���(iiO`�(�<�J�Y��*���ZZx��h;qu*�V�#4V��!�nS#���z[Ϟ\o�{Ɵ5q��߄��{�K���7;�M�m)�sX��u��ӟ�8<�U�u���\9��A՛�~�pz���rk��\ť�k :�d�����W:e:o4#׹NC�������1�%��/,n.`�%8f:�ʮ�4�)<O�8x%�?W�/7K�	Ӝ]x��.AَZ������9R�N�u�N���n��^������[Ւ��������o>z��OP�Gg���Ξ]����~��)��c~;��b�X�vq���(oG�g2�b#ƚ�_aˠ��<�d�z�vH�ޑGt�IT側�=f�#z<b�Euek����MKx��=χ(�m�����sˁ�{˺��t���wӠo-�w��ed��ם�:����m�ƾJx�\[�A1�u���� ��-��oQx�ob󳫡�1�����l��a����拉y����8�x���Ҹފ�'QjԼW���lDB�U5�C8!D`����<�4r����=)��M�>����]]�.����zs[m�b�v������Q-���	���I�h��.u��*=�}��Q�d�������?����~�}�Q]�Ȉ�/����Y�\�B �/��c�aE`�>�{�A̠L�@!�`@�U�!�eX` ��eXeX`@�� !�d@��a�dBVV�!�a�eX@��P!�a�a�eV � dBVV@�!�a�a�dBVU�P!�eX`@�!�a�aP!�eV�P!�a � eOL��A�E�A�A�A���a�`ea`Xdadeaa`FFaG�^ǰ{ � ���� � � �P �D � �@ �#� !� !� !� !� !� !� !� !� !�@:�z � � ��U\22��Ȁ� � Ȁdr�0��2���LL�
2�*��4L !�]� ��¢�L�!4�0!4Ȥ0�10!(l�!�dR�&�@�aB �&�@����=(�2�0� C ʰ�0� lU� !�aV �U�T!�a����������� AiTa �����}������I��B��Kg���?�f����j��q�7��u��I����o������UE��!���c��E_^0��+����� d��_�S�C�Z�(������������@o�{�����@�Q<�� ��د���,���@ �4����� @  �L $�,*���0 ,�	 @ " H���B   J��(Ȁ�  @ 2!"*�ȰB$ I� A*� L�D�R
��G�a����?j��R� �@(P����~���G���~���9���j�������N�������z�g��i�?������?���X��+�܇�O��C�ޞJ*���UE��!����E]���={	EU���&����=��`������ǣ��à;�ETV�H�����QU���(�����xp�?������?X ?PI����**��?p�_��Q_��a�������~�~�����x�ۃ�����{��y�I��~�b�����T���L����|����g����������{`��>�Qu����O޽?��!�����e5��e��>�u� ?�s2}p#��|�c@��
�R֩T�J٦��Z��V��Ҩ6�Z[3��ei���+a�P	m�F�TV`0͈�R�U$)UQ���٩M�V�-���f�36ͪ���V���h&#D�Ukm٬�Z��l�ѭk[-�i��FTͶ+lj5�M*0X�ڤ������u5���&�amiY���іi����j̪�͖����̳E�F��b������4�LcU56��M�6Y6��SZ���[j��ثkS0n��m���*�   6�^�-��.W\�N��R�Q�]:sYQ�J�N�M5�ҥ�v;f�I���ݠ��A�ft�ꊵ�Z[t�U�]�v�G�G@��Ȱ��cb�U��P����  	�<�c!E�4(P�{���
(P��{����B����СA��}�
(��l�/,��m@�p�2�(�W��b�+�P�l�5�clU���wZ�\�+�a��-e��0YU��͉/   Z�@=Y�F���P֕�wݯzwuͬVi�@L�չ8:�P�U���xP٪���2��
+om�åuU�*]Gjm� ��8e�ڴ���-�ƶ��f���5���>  7� Y5��ۦP��t֩m5�ݮ�iwp:4���vڭi5��E	\��u��@��<��� 'W8頡�:��mL�RU&Ie�m��|  Z�k@ys��SL��p�
�wKv�U��ˇ]ۭr�;�G���8P�k
%@�r�
v�:aJ���c`��[l�a�,��ݽ@��[\pt��ژR���n��eU����Ք`	U�]
�� 4h�QJr�v� ��թ6F��ٻ��mD�i> z��Z�s��4��(
�ۛ�T�i�];��]����	S�x�%�;��@H���yޕRS�{g��*^�M��Vũ0֩�J��_  9�Ϩ%�7��ުAU;���(Rί{�R�[מ�	IsǷ�B�JU{���)HUH���y�R� �y�zRIM���Q%H+{ձCm�l4hֶ���V���� |�P���}^�U^{��I ����I@%�^\��N�7��z�$V�c�Q^کCr��R"�+�{w��������=JT$��C�Y��jIL�٭���wl_   ,{�JE%+�_s�TP��y�P��J�v׼z%JT���
*Q�w�)D��]�%�9��T�K�Or]��R��z��R��P_ "��JT� S����� &�j�i�*��i�  E?��   ����Q3@`	=R�eU&� �_>���4}��OҬ\gҍ�M�l�A�K���cY���kp���ꪯ����.O�����Z����V�kk�ݪ����ժֶ���V��Vն���������^~���J�?�ͽ����cw&�Qe�E�CX��Y����  f�Z��2Pv��a+,�b��ç�[�
���EW�u���#d���u3d��Ii\������~:h%�ч�j7���RB��inF1,�y��f��`�0��ǲ�/��t��)�[oDX��#xAsc���*�,60���WYJ哣jB���]�ux�ś�N&��ɡ��p�
�ڊ��6�XN\��EX�u�"�5�SU�+����6�%`�S�~��bu�I��ؕ��0�Z��T�[j��Ōf���f<��[)�j
�wM�ӤM�M�>,d��p2�HlRC�U�>�"�cN��y,bm^,f���t�U���u�C��a]��B�ധ��q9�'8�|�繐���
K�h:׹�-��o�^�*H���Q��і�u��2A�-n�(�/E+�� 8aKji�%<�S�4�A#W{x.J���۬#�`�,|�kA�(]lP�b)%���e1vֶ�u�yP�%������K �6DB�|�ףt�1�`�Ǜl�K6�j��dA���ǩҠ.Z�1I���e��k(*͗�F�=N������"���6l8#"VU;�޸��R�.� ΊY���Z>Kv�%Q�j���U�R�Ew�I��r�Yחsq�(1�Y1�M��j���RQ81���4xYx�n*�;�pV�u"D�io-mh;B�5�l�wklhF�J�5,�\�(�u�S];�s@`�-,|�K�H�6�4aj�D�>
�!spne��
�Ϛŭ��Е���4J�r��31��z������%e��r�٦Vfb�j�H��EG`�!�f֔o^� ���xMIaۥϣ�^�/&d��p�P��o�E�@����f�9��v�[�&Y'Y�Ng��ٔ�!Dp�Wnͽe\��R(:ϯK�,�7VťK�M)a��U�"*��2�d����4R�����ۻڔ�L[6�A�f���f���u�ZjE��)\4b�����9��.����0Ru{�r�_b��d�Sd"w@�EP�`)SI;�x31]��1uW���-���cf��)n��ؚxJ�HT�v�.��T�Z;�VJ7�E�X㻩M+Ж�h��*�p}eF�sf0r���R��V(��,�$"+kB�h�$d
�<���z$ьP���(���*�U�E��*����q��o)��N!�U�Ǵd��,<`�+Y���
�p�!�yR�dy�c"�֘�h�+6�v%:w,�{�3�֊��t$�A0-^i��{�x&�2�ŀ�yyp:��oUS�����*|S�.�2
š�4�V�ݢ�i�O������Θ^1����&���{�<�� k���*��]�j��V�q�y��1p���<#
F���{��ˠ�i��++b�M�l7����FBp@7�Q�6�tr(U�JKE��9y@��zM�Є��eX1A��K
�r'H����Gh�{.�x����xE7��C�a�6��1^�I#��ƪm��a*dA�A��.ߗ��b���!D�d��/H�ׯh!�:�C�#�C!��<��0�Ӱkl`���5��Z�Uӵ��B�<0h���L���Җ���h�m�TE�(5%��B��b���(�4�S����(n�' �V,b[V�A���O`<
��C����F�d�f�ވ����׋j�Z���p����k	}��Λ�CaQytLa�0�j�L�i�M[+A��nY�x�.ЬzhX�Wu3a�:ҁC��N����i��=�Rec��Ù��(JZt��L	��
�*kE������ù�~b��ix�"���d�%�����[j\n�V`�H�yBL���(0�n73K�!������Pd���lh��iA�u�#Y7�%r{��,�`�-�FPZ�k�Yl�^�0Ջ�5�0!%���
 i;���neBMjt$�V��W��ĮӍ5𚶯ih7�m�]e�n�3��D[���S�pSj��{{�jan�-+X0p���%��4M��ʺ�.'W@V����H
<[��B�E��hƪ��tҢ,�X���l�Q����ZCj��Y�2����)�e�[���8(�I�Ż��ffD��Bqg/d\��zR=�PDm�/q#FR��3nHw,�3+҄ۻ�љ���H&�)&扻���4�[�5� ؖ�0h�	�V�PbS,�J"�Vύ�b����m],ڹO�����dA�n���=OA�VsE@Zh�f�u�VhM�4�Wَ��4���?&x�=�J��7�cK�cԴ]�5!����>Q���Ӆ6�,�ؐ�x wP��wh���Ѽ
��mݥe-�f+��ge0�cT��I�Ӗ�U�H����J`Ϧ-��ñ|��t��Y�AL���?�o������Hm���XƼ3�Z6n-�*��^�e��ܔ�.;�m����.ݙz��wj�15R6�mψ�9�&��]�GR�L�卤ݼ{�6�$�w�1�$��5��a$&$R�[b̰u��N�E�F�ٕ )��QX�[���޳��x�LJ�*��6�e��vn���B�g$�-�+-e�Ym���i�Zh	[f�Y8���Y�ZsD�ю^���w#؁�Z��q�����H�h]���Im04JӔ j��:�ԙ�U-��feU�J��Zv��Z�x��%�ش&��P��`�j�X T�<S��P%a-h-A�����4���@�J�6#6�T#�R�f	����΋2�M��I'��(s3p�h��r�
�d+2�;*�iϮ�Ӓ}�|��RX����M�o��A��f�ecIU�D�۫�wv�f��#i�rd�
��Aq�r��%ůAsj]Z��tcjc#,^ݻuk�	��_ۆ��F�e4U�
fҋ�Vy	gC70�3��JNej(�)n����0SB̆S �elo�1K�.�y��i#-��TnF��ঙ�fj���P`��CP�C��'"�l�t*C���J+^U�]���i�4ˎ�8n�MVwYd\F�<Ȱޱ�dU2�
�ڗE*���wTy3�O_pIpѫ4����}���7�'��|��Q������a���g�]�[!ݥ�tU��ʶ�[�ߓY�bQy���)�y��$��GO^#x�0�/\��w���R&ԙ2�� 	�6VJR
�,;N�-�RY�Ǖ�8lԂAg6͛o@�C[�{�	�tNR��ո�q��mǛ�kwZ/mY�`*����ˇSȭd�k�u�h�Lb�,�ϣva0n�N��F��beK�h�F��e5)bSl�(�7%��
�˕`�2�M�8�����T�@�жm�IS��
XR+5����T2lk�T��h���[�O��%Oq���%�w��n�&�8�U�W`05��v|k�/���a�)K8�jAI�fx+0���Z*�����u�N�B�<�p���Z��X�eݠ� 
�)"��^t*l��fG�;��5���8���b�j������F���5l����$�)f&���e�����H���W��dn/��[���x�Ff�,̃� �L�"����уZ@� �껚j���'�66m��Ux�̵Z�)���)�-�]h*�d;�K.���^��|���̸�A�WWW��]�n�Kb�V&�V��j��aAK�f)��Ga�b��t�����F�8`��y�`���w��Q�]$��]�tԕ��j8a�$ʙ+$�X���?n<��W�,pa��$!��y{�[2�f�QjK,�m�w0]�'J�h˩���{Cu&��T��L����#ç����Fc��6�_ ����\60c�ZR��W�*3D�HV�D�)�:��w.��0��q�1-�E���nV
�b�j^[Y��*ٶ�T�'L]��ckSBӷz�"��T�T��3Z���w[ ���e��W��J�=U�	bc�&�*���V�8M��:��iCVXݢ�'.a�R����Q���$,6��f�/8��L�#���df���e5��b�--��:Zؓ5L���h��z>)'�d��e�,R�B��ŗu�@���$0�/���T`���cr����Ժ��Ӡ1�X�� [���h�����,;:ɆWi��{�dE.�6/��*�M��&hU��03x*�,X��٤rؽ?M�I�jMXvO�U��˰�l���<���Z�"_2�Z@���A�A�#�WZ�5�����XN�;D,�Nʳ�Ԕ�M^�i�]˺�/A�R���I�����Bb������H���`qc��ȩwK/`����<�M�1��æm6E�-Ӻ�r��M�v�nQͻq�4kT�'H�hP&3���D�L&�"�R���45��Gq+.m�Q��!.�����LN�ؐw�F<�L�����Tn�=o��ا����(��ǩ˭�n�gc��!�Y�U[�b*����#�R���Z�L�s1�o0��j�b�3NГjtr�\n�,Hü{m��lU.�(V����Z]�G!J=�@��Y�1=76�4�;6m<�A�Z�@c�)ВF��:X�-f�J
M��W��=�=����?|�d8�ePI�]GDd�{zF)����1�_`�B�� ě�j't滌5K�]֪�,9����ȸhM
S�Y7[��ԓ.�2LL��6�;A��ʊ�Cm䊲��M�.��@��F����L&:<R���X�!G.�"v��F��1���2F��a�{LE�;�F��N:.��:�A�dsM�n����%��#�� '�����W��vCfa��2Rޕ��Ѽ�1�F���y�
�}Ƒ�bj��^�u�$��T����+Z�)�#6<���V�շ�2�0C�FX@��4�1 �TT!'Z�V�T�L�u� �lYV"ۚ>ej�+6��Ď6j1m�P���9�D��F�VkM�y.��'(
���5��.V�G��a�h9���;"��B�l�K4I�� �33#�Z�-Q���hQj�#��N��4�P.���%�W��[�b����.��Ej����:!1��# U�(M��鼼q�h�v�cf[��B��W1D��0�J�}�3ᜏx�]�/ �1��x�X#�<�_-H[}�͚�g�&P�1|�f�w,�h�-;A�q�92K�.�8��2V#F�Y�N�!�Z����ʯ%�(l�)�{,��f56Qxx�:�M�Gv�����GB�m8U�v��w��(ZP�lj�L(Lt����Ǳ<�mݖ�LT�4XY�nLNѫx����f����76�+%�`���@�ʆ�j�ʗ�e���V6��B��;�T��t!?`��dK�&hǓPn���ehufc�i&�=��*A�e���ǽ�fo�
-$���-S������g$���|�7�F� ӟF;xK�Hf��QX �b:�tqQ��4�k�Օ�;:�K�H�-梭�j�{�����Z��j�4��%����d=���٬�Qopܚ���E:)�*��&��ĵ����J�oRx�7q<�5(�Z�G�YX�,PST�)d,������P{l��V�-MXĆ���-��
�x�;9<���9i�q��Le���^�.b��:��b�Cǲnc0�(&�2��a�d�N�R��>Y(��ݥJ5t��:�JI�@8m,KC�J
�0Ńm���oq27�����U��w*5o�Ը���,U�l²���a]mN%fZ ��Ԕ�Bm�Q�F��H�2��:�z�zq�,��5��Ԕ2�d���/5�a(m�o
��W �y�X�p�[֦V?�����e��T۳��X��J�����֮�ʆnbYge�Y{����Js5�4V��ʏu�]�U���U�1���t �2|��3R�X
b�`�%,� #Y1Ն�;�V+��f�N*� 2�5������F��T����OvV�͎��I��Ea,�4���DJ��Cj�`��hh|�mn&�ɘ�|-�QbA+oL�cKب(�Ȏ}�k�����E�Xf�ɯ`�.�57�Ĩ!�[W��Z�@=2 x����Q�;1��M"�&�� �%��e�kol��!�aN�ʑ��nt���2R4.\�Ɯ�un1(�@h�~�AJ�v��v��g��m�o"�L��V���1�2�47�aI����mc[oQ�N��/��1�[j��unIf�1�"�b���r��Z@��� 9��~[ �RM�Y�y�`}��β�z��d[���|�yy�	���N�ǹ6��I���O$�+��B�:�܇ަ%nҧKJa�O6eA�����B�`����+0��*�#b_kV��#��Ҹe#��6���0,��{,f֚6�2R9V��V��,���Y�2�J4䍝��u.^��	��q8�k*���SSq?����5���C(�	R�����n^��(2U�zZ��W�|�6Z�i����2E(:��YV(K/��A�ee�6�
��1
�lճ��΍�����Խɍ��d���v�R
ٹ�Qq�+��\pȎ��3�J�ؙ��>Ɉ�5�.�k�2���4!�z�P���P(�i/�-�V�n��r�͝���F�Vj"Ea�%ک�V�����l�Ce*xшaf�-j\�HX-���[����wHԢƕd�ೊD6�r[YsK*l4�]LQ�kv�g�f�³U�TvS�Q=�����`���G�2�6c�P��|L�O;{�����9^k"op(���qF��XY�/}��,]7}g{�S�/����3�Q���x��Ns����ҹ�ᖸ��_;��u�X�����.}��,Pv���Uj�V�}0owp:��Ln�9��p5�[F@I��$�W��N�q��Y����v��~���MB�/qk,e�|y���^�ڼ�%v��}���@mh���G`Y�D��2�;��0v�8�D�Z��X2l>��}�zW@�`p��#��x����u�U�'s����i��賋�E-��&N#�h���s�>�BW��7�]s
��ZN씙��f戮��`����s��h��>�0���vcX���9���^՘�)v���p��"чr�ޤ涷u!�f��:���`������4�u;�u����舮$�ƍ-�D$hg#պ1q�/W���9G��I�׶p�	�1=�Q��ߍ��{֬��c�Dս�ȹ4�v&V��4_��u�=sP����ꯊo/��uf����"s�t��ld]��:��^�/�@:�>=v�2����l���VNk$7��Jkh+��#�}����Z:�/kX�����{Ӑ8�àS՜�9�9=Ε��:ҧ�FE$��kQ��N�]ۥ�=�-���N�Y�޵˰�3wMb
F��l�<Z�o��OH\gi���.0f��:�=���,�x;��:��z<��}��=����(�ӻ�|�돱偵,��iN
����*����
}�0���+�M�����"�N���	��	=�b��M�-p�l�Z'j-�˧b���d${,��K
��Z��b*<c�z���`ѱ����x�8o���������q��2ۭ�hjZ�x���h�PB��Ӻ"MAZ��h'��l��N�h��������:�bG��0'tf耹sP�87�����+䤢��i>ҏ;��$�r,�<�k�@��b�Hz�-9�z��2w�L�]cJ�Tm=K�P�Xs��ʳOo]]�Z�~�v�Ky�O������ �W�=u��pc	��Qǧ�g��8׍��(s6û=n�٧���b5�6�{@���Q��<��a������}�a��7a�W�Ve���G8�b���]�z��a:}�+=+�-����Gv�BJtt�'����%��p��>��]�����Ӻ�ͫ�흫ѻ�;��3�r�:�"ƀ��Wǌ(��P���
���=[Vb�4��i.di�<g��Y
&����kb��4�q-7�я�&^o�-N���>-���(�\:�l}���:��dx�ۜ%⡼����]���O��MX;n7��i:�yiX���Ԍ^���D.&4z^�����s��<�����A�$�­ػF���lR��"_,]v���X��w���h�o�E�\��gcmÍ�a�R�y���2Ҧqf��Oa�ފ��9v%;_y՚�`B�t��Ƴ`��kZT�Y�:��vŮ�GoP�ے����Ʉj9y��n�C3	�"U��ˋiaq�V���I����:�m�;=����W��#�As^{�{t�Y���)�a,Gm�����W��0�k���p����Gu�8oj�f���kE�-����\�^�������o2H�՞��$Nl.Ce$4H®y��W�W�#3]wBk&��]Z��:h�U��c[�J��&ռ����ޝGw�)>����=���P�t齴���ܭ�Z��v�\2L��h�Q`��c̚N�A`bchؖ��3e�!�ϻ��T{2�}îacʌ�իw��_���b����!g,�>��C���ď��']��Fe��sZ�x��o�ۡ=�T�(V�9zU�(��r�Gǋ۽�p\�Kᕚ&cͼ�d�0��=靫9��t��Dn�g�seZ��/{�"�7BA	�KD��
h�х]�����QM��ZC�,P����w���:e��V ~x����G@��$ �!)�D��h.�r�t�.�T��N�dٰ>��A�*!�X�}�+j>��B���L�j���&6����k��eH��/?ץ��dS��$��+��>G�n�L�͈J]srPCw�ӻ�c�w�C�S�ix~s'/c+��� 3a+�0�i���[�Իi�F�ox��;�)<��	׀�&�z���V�y��o��i`"��{#�����lZ4�o\��󾾺_!���ߞ�"U�ܰ*ﮌ��z)v]�*[�ֻ���.�RA��s��OV�}pǝ	��P���-��~g{��<��DCWG-C ��Ӌ:�#ۉ��J8��y�5hٶ�.���۬es�.�~C�<N����ٚ$L$��%���R�fdq�x�,�A�z��k�7=�)�wh���2˿yy�v'�FuL�+���飃�g|��Y;ԔpGM=]#�b\6_�np������ˣ1;*��S�`���ޫ;79�ȍ���4e�t"���3O�;.��@�D)�`�F�;�"��u]l�ݜ$m�3;�8��
MTH�׻�4f��ul��G8$��� \�5Σ.=�ː��h�:�_TxK,�;b5��v�p�B����T��QӾYU��OC�½">���L��ٕ�"zV��BJO"��H�]n�[��oQԦUp�N� ������G�׸�MD��DOTʂnL�i�0Y�iӻ�-�E���9����/�^����5�::���on�S��<'K��1��0��6vз�b4�	,J��.p�#]��(�	������z��%�5�%��
��dAMI�b�9/@����3��|4]
):�-�9���ǄnL��%��ge�xQi��0����oż�r��u�X���l�t̮%F#Wx~=�l�� sݏ>x|=턎'A׊F!��X(ټi�O ��5cT��W19���n,{�@�@π{��<�|�ۨ*
h՞���c���5DW�\Zjϴssb��gY1�O>[���{KtV�9����W��yk촉�I`\@�4��P�*��lʫ��pc���n���P�#�ߑ}����%�_��-�l뫾
�D۳��
�����'�A�j�����"j�	�98f��-�#�F�k^*\��w�	i��HSn�yl�j]͖ޅ�Rb��9Qm-+c�n��q���C�����66���Rf��t$˭�z�VU�HPҬ=s:��հ��=�������ɏD��Z}�j��'���N�WS��ݳ|�!i�r�a"�9�L��C�H9JD)���=�Wy�R�l-��G"ĕ������K���Bb6lb�:�9��vh�aJwA��㝧�9���V�L��$v'��Ο|߲�Ė�{��NXz=8]^Ǫ{E�w��Q�ʌ,ax�q+3.M�X�U�`��#���lXޡ#FLw܃�{��|0�]xs�**�5����{B�A�+y�@��m�;tw^ʇ�Nm}e:8{`�p��m\/n�"��=����'q��)�=�1�zňu't�h���<�	����ڰCD_:��Eέ�S�F���C�1}�*q7k4��7K0�К��ʄ�W��]�wFoAuJ��L���wiWk�1�˛Ω&��4�x��]�\}(K�Y1*��mؾ�X�?��AAU��v�۩2�b'v�w��5���C�m���sU��*Ez�tk��E��
�����"�ݲ�iݺ����ד�'���W��ohao�Wq�-M}��:b� sNM;����>=JOm��2^�7���gwדi��p��X�{�:@��FJ����lE��}�N퉸���Z��-���Ӧ���Fo`�f�v���N�-�,��g����ȍ��7X��;+=���Y�y�Y��N�y�����<ҟ'��<qםlO+�;Vb��u���]veP��[�ܯE�T.�-�s�#�Ǚ�˒t[��u��v��]�@<nk�KR�_	Rˎ_D5����b"-JJy���f���ťWv�v�ɪ�Z��gv�䜦UۇY��t>�C�1
ݭm<T���Gڄ�v��d7�7�Tӧ%���"jb�r�Lqb�~zé�u�t�l��f���ln��5��ݕ>]F#�W�_z��O�o'S7dr���+,՜.���.J�%n��c��s�j�� =݊�0�ݣ�Y�R����Xz�6hF	t���2A�[R�mc��r�M�����u�{r�&�#�L@`B�7�on&���{�W6���z���[����ğu�f#����2�Lv����̱h��a�ߡfv��a�v�gN���|B��E�}]*t�wpz8j���x�4� �/�%� �d)��M�Wgu� �U)g�j��:���u�D7:�_�)`��e�����qe]�PLC.��j_:��ot{��wy�s�=�ޣ�-�l���l����^����"�3��g��|x���'�0Vࢱ��W��P�hn�Vh������⽤ٶ<��o��:w6uf̌�k��/8V��j�m������CP[�7T�j�<��XNs;:ֻk3Z#1�ݲG�<e�p3�L���������!�`�^q�B`Y|+�`"�8��9M��O�Ue�ǘZ�H5P':�D_fZu;A ��`g7���^����~<#�t��&��3��S��0>j:���B'Q���W%����`iP�؃�2j�S.%��9����.S�l���q{O\��a�z��p;�4 :�;k���������z�̲��Ph��Qѳ�F��kV���1��;zU�0TEl��Z�E3*�EcHM����m��ˏ�kt&�)�P�f�%��k]=�:q��F�kz9}����p4�v�u=� ���a��τ�<v�˥�bh��M�^��z���:uvyݺ/T��y�[:����W��с'O\��]�e�lz�j�{_Yּ@�Y\��p4o�W �y~~ޝ��<ȱ3M�dc�	���U�����F`�i�@^�!h8��:��0&���a��*1����:R��O���{�hv[�a��
�ǎ�/����E��ΰ{����at�4s���4DB���x�Ӿ�|����"A���e�댡V�˭��Ũ[�F����]M���B���j��ː�U{�9�ܜ��E�gD��F_{l]ŧ:�+���OM�1`��$��zXɵ,3������{�Y,!�5X(��� �n���F�i~�D�����':���ܙi�c��Y���o�n�V\��Ӗaa�tH��R���ᣇ��F�Rc^���<�q3vt�KJ�if��«5`/{�.`� �0�$����5�$������y�2�s��0^��K��r��j�E��rN���v�,@���4�c���#�a2�v��1e��'Q��tY�<��r�2�S��2(����h��R@ؼ�/���xaS�Ў��f�)��$�F��[p�"��V7)���t�a'�M�jƈ�専�\Y���ۥ	��P��ʎ�,�`Fw��Iea��KEɅGp6�r�����y1�u��kE����4��[�MPL��Y�'9LpG�,��]�U��Yɤ�y��&'��ɗ�e���K���L���s��}P9�d��YJ��&��V�.�k%��bN݀�j�C�Y4��'Dt׽��k��RN�s���8�($��Z�)�wWo		��7�9�|�Ψt<���sk	`����]��mm�1+����Ժ�\�ε�s�)!O0��:�Q�]=�ԑ��^�	�i#����ڂ��s����Mgݮɒ��ۢ#3	��q�v�z�����9��QJ���Y6w�/��yV-�Ƌ��Ii��a[E�U��7��}��z������y�	�G ߎ�/k)Y)���3J�̬�W��g�����ԋ]��L�c��Eˉ%�z��j��S�{\ϻ�Z�.m�ۓ}�iR���0˻"k�fC��Eb�gh���sK��V����YG�K��<°��+_s���`��-��?�t n�^��nxZ8�̺�2m��-~/o��O;�uWm{"���+=�3Ho1��Yo�9Jp��Ycg� 0��\��{e�e�4Dt~ʳ#��d�
�Z�n��,���{*���������L�3���W�ZDՔ��9vW��W n�n4�M��Dxy�k�R���7��`�Qn=)������Tzݤ�]nL��)j�r�gDMX�\Cf�����7-]<�9�Q�o2?#[��y�*H�Y�e
s�6��μ�ش[����}�yv����6o���vNn��{"cyn�=f觕�RoU�w�;3����Fz��R��]v�}Ao-��̐�3�QW��y�x�jٚrB+�8U^���-�˅��>�P�H9L:ǝ�	�R�Y�Q��'%��CL�;,c�q�C�enaͷqT�SC��Zؼ�]�Ճ=�����ɓ���)�9{4��QC�����"k�aգڞ꼌X��3��|AYSt��s��-�p��}��V���I�����M{w0n� ;�b�	�Ų�sy�I�Ó^`�}Hdƅ���P��\v��Ï��fbC<2�)�[�C
��}�]kb�;3U -a�6[��3�:sr���Dsd��q��eu��$�`��D���œN��E\��"0=��g�vb�3{��m��z��z�3}wD����_���L�[�Yc)�)��7�p�v�Qܯ�\I:��-��{��zv]\�0n)�T��>(p��Ƶq����tK�B��K��{@=�G��D����}�O_ذ]F�r.�A������G�����i��+�6�]��{[�o`sz�.��'�Q߼��4����������߿�������m����Z�km����l�xx3��(����Np�V{����9�uvoپǄ�D[�g�}(f�'�L)�b��r�aۙ����Z��*-�TS��mT��4��Ws��&q��3Up��츢/5if�>�H�*�SWQ_=��.�a��z�:�󎥛V*v��$�=0��M�i54T`��tl�Z�0�׈�w�ڦ�<3#OOv��lRjd���s;PfJ�X��w��)�%G�I��&in�LWER�r�09�.&>�@�4耷U�^D6ٙ�(�@�RM�Ek{Kc�lN�;ST}тO��A��k�m>*���
�X	�N{uG����#�~�%���A��+G���X�=�y:�@�)����T���Pݢ��)��V�|����p�ѱƦ�fbү`��yV/`rGI�֫Z���U	�8B��=�&��F�_��gp�*1�E��@tk�'f#t�R�~�"�}8;$ˁ7�
�X�d�D��]���O���n#8��f4�{&{���QV�'{�T~�)y��fi�w�ٖW<��n���k�fk#�����U@8ľ����;���%������ʗ�O|�܋EM�}�s��^VV0v�Ʀ�W��^O1���۹���=���1�ֱ�]>.�*%���j�t�p��Y��(��˄h®�i��3�kH
��kWѾ���EE�)�U���;�,���Ћb�s_�Uk��6?m��涆9[$����	��k��z���7A+�ٛ6�Tm�F��_C��,g��顛z�0��E� �-�ɦ�`�S{1@(�7Q�He�6+gLɜ6�~C�.j�(�WMP��\�RGUEȞ���:TrU:�*���;��9�#B����C��n>��j�u
,����6[{9>@��p=cg�>���j�]<+'���YB����	����b�k�u+�-�G�o�Fs e��Y���O�ta����-r"b�;>�,{ނ�q�M�ݐٛ���v\s�����ZZ�`;��j�w򍇌Zs�CN��K[��󬪽CA�L�O2�	�S�+=�A9[&;�47�iJK�ٙ��`��C�i���Yl�OX؜}�T(��j� ӯ��H%K֏jF��s�d		\y��+��<(`���[�q��&y;j��Qa@�����-+�۹�>PV[���c\�ø�����h�β��Tm���fn�
��/��)(1�s��Բ�H�)P�Yf�3��k�
v1�.�Q͐A6j��L����RvDax�*W=��8K��9�U�Z�R���u���1]�"�[��Z�R�"��Ѯ���M|����J��t��`\��h��L�m��dk�^��wy�6����]GV�k�WdKCD��4B4���p��6�c���8.[E�QB�l+7����k}�ڄT卞���;ss-��r��O��YY�;����������u��7�1�ԇ	�wa���!1��z��TF�1(�iQ�M�\W+V/��B�[<��W�7>��9#>�X�l����+��Rn�Ǩ��iUtlNWZ��fC+���p�З��TUrǖf�a�tAu�$�t4ڄk���tm����w�f�8'��4vT}N����AL� O��wS����+:�a�`[�s2�b2�+*Yk\p����ݸq;�������z�qH���qwWgLr�6o�I��P��Fp�\�Ѿ���r�<ksgm���ƖTXeB�<߭��	�m�t��Ԯ {�=����HF�I�Z��鈑��zVr��`1S�z&}%9dvEڵ�Ɗ]��r�Q/:V �\X�>�K�$��3��o��A�Z=5���CI�9YF�0�cqv�̠'n�`)W&+[�_v,�:ª�g>$
�l9�����R��L[�c�y|7�=,�1�	s�?,�B���)0�s���T�+�z5+dBIΥ����ދ���VrT���3�k3<�v3p8�����f7�C�n������1)�Ep�2s/z�E/V[��ӲeY1 �������'�2�!9]у��.܊}���=ά��r�u�ݯ#�:���6�y�k���Y�N%�;�:��	�f\�#�)���3�Eq�VI]C��Ρ$���!�@E*�$Rb��t_l�R�gS��P�\�_Ӻ�K����l�n��1Μx�5xEKG�(mL���8���vm�ps)�ntn��#q �䛧�_}����ς��pC��TY�<)��LB� ��ܻݎ��n�}����m�����̯l�=;�3	�j�=�h���u�i�-/37�ά��wY�Ȗ�51Q92�at3fۜmk}R�U�$��lX����ww5-��r$x���
���K.sݽn�G��D	1�D����'�c�8P����VIb�=��4��I2�m�����f��ں-k	i� �^�,q�8/�t@	6�	\a���e�ާt��2h����r� ]��1��;�+:�m78ٮ��AX+�C�X��6濲&^^��](�n�N	y�v ���p��pe�L����E<����Əy��:YVIS^̻N��2���ې
q7��j��6Y�U���)�X�0�\�ڽJc�U��bEA�Ѯ�Aq���]�x|��-����4�'�f���1�i��p�a�y�)�tGI��C�����l��v>�; ��C[QT��S���a���U�͘H����mZ�6+̸�e+�V[���n�ۘ� ��w�����u,��V�\�d$(���ah�9$��C�Zr���� i��r���gHV���<%9٨ݤ���,Y�����1]ܛL,�����) ��p�k�Ϋh�7��*���h���m˵r"����u���m=��Ѹ�3��p�MIn���],�J?]�JԵ&�jȹ��5�F���鷵�#���لp,߷����y���ؽ���5���Y��FI���0i��ڙǹ�fH���V��u��w8C8c�΁wh3�e42�:�7��4k����ؐ��c�_�zy{�#�A|�B��e"���~�fyu��HO��A�+�`Z��]���?��c�O��e�s7�c��Re���W����&�Q��6;���d�lugz�9`�Z0o��)|4c�WM���ýչ�냭�	^�;N�:Gh�k���b.���Gr�w��6#�7������n�^_qЎ�:�^Zm���0c�����<�:}���0{G-94).]�a'X���f�m�#��Gj�m�#�t�	/�ٕ�գ1lK��6�[�^Qz=���(��zw}������l4���\�_VЃJ�^*�Gb`hʹ�K�S �[MHdʡ���T �f�c�a�&��%���f�]���0�)s f�z���Έ��._#��2�u�W;5��'�F��+VI�>�>��L�vAO��訡��������n��7Ko�&$�#��p�i;�V�xep�ivv���A�&�/lB��d� �%oš���
��(�켹�SWb�]t�f�{��p�%Ȼ�C4�jyI�j�}�=CU��I����xzHV�$����qb�j���M]h�O{��p��ޠ x�p�i�5!��n#�Ǉ����/Y��x���ȼ�&�*�oM�㙉�P=��i��5!��J��/�(�.]����F�q�YFfwTM@��6e[�4�����έ�
LR�o�?jٶe����sV{$F.۫������!z���`N
�%���l��ø l��@#I��G��LnT[��N��{3&uY8i]�(}���q�ˠ�0�o�X/��۷��|0�͎�C�Y�$�jθ%�rj�
qWo���7\Ni>���{W�-ڧ�JC�Җ �6ө��{�TVlu�O+/��ayԏ��{+W	��5��ӮL75כ�b/�dS�`��q�Im!���nA�d4$6^��s3B�v��ӌ�I�QJ�����F��w]���;aƑ�}�ΞƷ@η(��F�nP�'��K�a.�m�EYd��^��w9ʭ����ُ2;r��Fo`�2�G�Q� ��:
���F+Hc4�mϘWX]�u��^n���^�;��o��ye�;w�Av��3/+�n��ܻ��*t�n�S����EmʄkI�
�a����y� q����v��̲�,�,�"�+�c����X��j�:�V�5��dl��{��U��J_lyjF���Ъ'^P��Mb�v��Ef���{ǝO�A�A8�mpf_<��P!�{�Q���PBRfn��F��C��zp�>ji���n��=�𚑫f���gA��).�Cqne2�ޙMW:K���q�V����]{.U���n�w%o�2�v��v�R�z���M�>�.�;����Ǜ+C��)��#��˺=��PR�Z��a��7�P���q��4��9��dh=�9oeS������cX���U/(�K�Qʘ+�ց���vΝ}G"˹�0�9�:um!!�7�!�[У�;2�gaXuDD��j�m�c:�lP�qA���g[��`�� e�bd+g*���ٗ���������1y#:B�����N\��{ZrQ΋�;j����b�n������G�C��s�ڂ�nU��].J�6������>\��0�{7���T�܌�9�/H�ۼ��o�"���t@C&��:��A�볇Kn
dp�'O��%1(*��:�0v�(iCD�� ��Y�N� �V,K: Pv�����#Uoo먣����9��e�҆<������i�]ǚ���.����eqdk�nv�SF�ي�{`��oq
;7C�_f&��O�,�e���ۨN�,�wXUF��%�C�tвR0���Y�RlN�0���>L]��ǕW˄MEm�M7��jC{L�M�fm/���B�N���t�V����M}��l����ǀ��K�e��,R���guV�LeUh*�!CQC��0M�i�f�Ǆ+�5wۺz �a�J�gD΢�]�h��9=�F�e�}K��f@���ů�!9:eӽ�V�-��O&�z�2z^m�;�c�ߋKE� R�(t�%�
 @��뢨c�λdU��r��%�3�
9w�Ԭ@ǋ)7i�Yz��V������N�ܪ����D��i.EqQ�״�MY���6L�(�3|��9�7�R�dT���k��/^�%�?��?T�{͍�H�F�:fo��M��	n�=�/3 ����8땍�6�ܡl"�鰍�������is,\w� �E*ݸ�Aw�,b(��V��s/Qe��%r_?�8�P|�kKD���x1KoJX٤��ů7��h�,���b*�l|�`z����d�k0gM�L����õR�tH宥=��6�q:��h*�C-�#JUh�߃�{��a�w���������!{��sN)ɾܮ���p�d�\��|-��E�Os��du]:�����Y����C�n����t:<��A��Ǵb���t�l��7�(�p���;F�a��$��s/�3���'os*\y��Û3�ӲGR���K��!6z���!M�W�^�ɲ>�8�p=��.��l��m�r�7�N �_jř���w-}�(���x��Yb�o�فѮU�n�h��đ[��F��͒���܅j
����$�i�ګ"�����ZŪ�����ؤ����\0|G6]p')��TQ��J4���4�r��?��b7�]n���1�s�v���A���]7�-�{�4����a���M�㍟0o%To�{7��[�����|b�1�;�(ȕ+y�Gtj��-a�'�KVzkc�[4A<[�m�}A�4cgf�n�怸7�n^P�:�Qg�e����&0L~3�������H���*��̄BQ�1=1q�<.��Z���f��w�fMq7�7H���<y�+~�O�,Z-��{�ʈ^��������L���x�|\�YH��/z萸^;��楦k3��������O��AEJ�1�ބ�t֦��0�nk���vp	P�m�]K<�6]��g�B��P�ZP�nM��s���GVst��t� �Vl�6�^��K�i�{�I��3���5x�C��x���ʗx�i�=��tZO���f�H-g� vC���c��;i3:y-�UJ���ћv�G��Ks�ɽ���m��7��M�� 7XōRN�x��M��Z\u]��"g,�8n�(N5\�:���x��r�LD<�&�vrN���r���Lf�	(Wtqc�̣IU�"�2n��>Jqw,�o4[42&C0O�As4�9�z<�y�#�>ٝ�m��	�$v��P�QB�C�Ui������D��
簎�R��WsF���=gj��z�Q�p=»�x� �L##�+����6/1�Ǹ�PBZ��k;Ԡ��wg@AAUb�k�\��r�N�K�zyύ7�nw�N76:�}Ř{u1+�Ҍx�b�y�;��Y�5�#����g�H5��#O뫆Ci�5�6�Zc_�ޜ�x����Fl����w�#AQ���Y��]�Pfኖ�(*�L��ͱ�Y*9}��}Ը�]���L*�ZΈ�z��WW]V��
d��fmar]f��t�� o�[S3�j���c�RW8��V03g�������7.���:�����!	1���W���!�oA0�����N�L�:	���E�e;L[]N�;M��J�mϲ9n-<5��"��>����tQ슥��w6��]���q�$��m�%`��2�Ag�p[xqE�/������^��~���/����ޗ]�}j���[�w�_����R��V(�u��`-><;q*FW�kL�+�L��{Ѿ��MH��͛ @�=�"�9��s;I�WxS�ns$����8�	�<{Y"��W�0��fdǧ��t���+ix�R���^u�W�:z�S�F8�TzrP�]ʹfҮ�yq�9csJZ�_L�P7(�v�jz֡����C'��._#�S�O�4�Q�b���y�y3�b�؎��]2��۹��^L�h�|fon�Bsgz�~a7ӯ=��N�ac �s�������C5����\-�tol���7�[4�������}\>Ĭ��^���ۑ�	1{�$��Wu�Q���x��3w:��Л2C�_��-+ў}�-��>�w��dVviʷ��M������k��Z�ڔ���ǥxװ��뜍�O{���
	�z��c�G:�\���m�P.�S.�ڞ���\�[3A�״�6k�{
�*�q���d�Y�Z��n�nm8n����Sە)���7:E��l����3�V���v���{E�	����*_
�RC�Fu��m�!<����3�/��<P�}����ս�4_S-��!����l��7p�^o�׊g�����َ�'�u�����d�d����d��k�Ql�^K�L1ډn���W9����v�=�<���L��E��8��.���]���L�(���H��9b��(e6Swu1���2��2�P$THX��2QL�LAE$Q�$�I,!�)�!�̲�s3ɣ	�&�I0��.�XH�����VL)&"��JGw:�d�E]���%	F ň���6D���		�1	����"&T��w`"L�Q�3L�$��$$B,c�"�Ĕ�H)1��4Bs��1��D�a�I 3�$��ƃY$LT�Wun�*
��E@�9�616�h6�R&f�� ��b��Piݮ~X���������[-��	M�B�V��e���m}�6�߶���:g]3�;�Z��6Md5^����g!��Eڽ�opP��2G�:��f���%P"�T�c�7L�N\��7�T��Z8���H})�th�u�gvu��a��G�u/��>�n��:?<�.��9\j�v�������s��u*i����m�� *.0�B6���A+O�+��+B���������������9��c^t�;���{~�s0���N+�d.w�'Fi�b���!�2p)u�(t�gD*k;q�8{ViG�P�r���W=Q ��-T����|kk�[;ƀIL�����gv%��~�P��Y��Ӊٍy��������E�4��\�uC��4�y\��YiEӭ��9�*t��q8�?X�'D ��Z��uPb.7$c<ݾ�,�>=��n���D*r���^����hc8IÈ�Es��^��:��S��_�ՙ�;��z����U�8_!�L�z����<��M_	,��.�V]��٣.WԐ�B�uI݀�,K��o�"zX�mCθB��2� P@��OT��?;��:7V:y��We�jb���#[����S��;�t�c'Sǩ�gФ���γc-q����QnCr�|���gkg�<�d�W�2�Z;��g(8l͓���U]w�n
h�J{�n��7F��5F�EG:[͠��NVp%�Кi=�/��<��(�Τk���*�g>���E���=v���#Og��uB��RQ���2��TS3��*R� ����KnsJK]pё-�����7��m븞7i�������ت0�c��*��� fW�t�)�QȊ1���ꄭu�j�Q�D��1a���tj�W/�*QW�4��q.�4�O߸�8�T����i�7g��\�F�r�d��&{�P��t��Ry@W���r����s|�S���#�Y����;5�8��]�p��EG�W$�N��x%��w�����&�Cn��������J�\u?���y�[g쮸���j��o\>՜�+ܮK��������Z����k��5�@;m�ٸ���(�m�F��뾏���b�ú��`�M�\�I�͔��6��O�2<kk��+�h���e�'n�7�L4���w��$NO|o���f�������C����*|�3���8�+�g�[��:�2���<��r4$���B�l���t����;F��m�B%k�x��+�k���H7������@�S�w��qo'%G��)	ǉ�9�^�{̫N��t��5�Է[�L����u78u�[fR��K
��ەk�L��j�e����ρ�Ù[�a,[�<R���joX��%��*<3z)#��
�|�Nb�v�6c;]�]��s�S�v=�Z4��:.|�Yec�^K�|�U{�8�C�ַM�t=�3aj�e�Σ��͝ev����g�fo���5'Ea$�:�S/���6vl����S�o��	�g�at��(V�g�Sw��C8�< �U�A�Epw�F��'������!\<���t��,��5��>P�X�Cj��|�������]4�d��r��I�P�$a񞩂�+Y©�Cjy�����/k�PtkU2��oΈ��a��O2�����ѪLÀ�'	�V`U�O�'���8\AwO�����;��\ﻈ/m�K�\�Q��5�*k���h0�}$B�P��Dc1U���oM��L�]�Ù�	����mށq.�AD��I+g����+Nꅥ`�a��r��Y=�_�P1�u�)��(���/���$>��E*�O��L^�M�ƞ��oݎ��������7Έl�1�ӳE3��F�"�^&��'��J�u��ۙq�:!r��S��θ�dgۨ���o;��W��"���h���BI���Y^��q�]���S�ZLX�g��p֚�y�Kmr���Ru֔(���ׂ�s�A�/*����ޘU���\�5��g����y,M��n�fv�}Ȟ��/P>���y���Vaﻮ�B�'wB�`9���5�b/�]�%�l"j9���⯧$|K�
�J-����;U��W����|�"��:�"�Z�3J�
�� @�<���۵�v���S\hU�&]xϨ�:��;~�Ub�O�x�=~2��6�u�+k1�5��UF���H�S����W�Q֯�٧��#��N��[�QԲ0$�7��p��=����Ms,�5��W�[U�n Eٌ�N��C(L�ʵs�}��%�a :Ѣ��Ƀ���߀�*���ǁU���j7z�_�l5��#���;(��UC�n��-�(𸩖 ���A��K���X�N[=���E�ј�a����'�{���>���G�Ҋ��[��E�W
�؅����\L1���ZMV�=�	Z>h����
2���e!�������'�_Q��\�]�^�G�C�_��ڍRA���28q�����Y�ݚ��ޓ�J�a<� 3SG�C�R!y^����-��\�}]r�Ps
���aq��r�s��'���*y{8L�.s��(q�0���4��35h��Y,Vjǀk�5^έe�n�0�NJ����ve�f[�P��Uw@�\�k��F`E���v��g��ݷ����Ü:ՙ�����ǵЗ� ��ʨ�tr,��;NBrmC�r2S�T����ä���_\�|�F<ͷ�Uj�c�kM��5��<7�S��a9���f0ECn�v�ݳ"�L�k�Ȩ�K�ǞG�^�,�\�A�4l�p:XW
x}��]l �TYp�J�k�J�_d�;�t�7����Y3���%[�-�N���_���N����޲c���sT�y�r�׮v��D�ԏ{P��yK�lDt�ee��̈b�b����yl6���D�:����h��f�����<�����:Y=_@?-5&;�b�W��S�`Ս�������AS�b9��]��΀to�4��on�����Y�#���lZ���?��򇟭��x�9���<���W�&�i��<᫸�N��P�X6j4�c* ���L���&�r=���>REb#���xx���L
�q��ʨ�������|��1u�ma�'�|��)I�q�W��m�=EW���8���0<'�� ��p"}M<�d�L�C��4��ǚP�4F���K�.G���r��T��&l܍��s�d�a�%��Q�����x����b�D�_{H�U!��a���Wq�.��î�K'ُ�/2utb�&���{��M��6��oi�&F�}�IM%���
�^-x���n��:���Rk/�t�R�3������<j�P	gê�crFߖ��o��Yr8{ge>C�r-/W����M�$������+п�@��ٕ�fvi��B������k�G�+�P��-S���,ɉ��'����U�|~$JGv�<�d�ȹ>�h����b��N�d2������s8���F�8OĠ1R�s�8�Mօ]s��Z:��t�^9����l�7_��პ:\W9xc?YsG/�IF�b��5:�����vx�� M������r�\4g�ڿ�;�cs��Bw��Wl�y�Nh�O=C�8�<~�#A�dP��hι��1�	�ݴ���V�����gf�۪�/�n��Q"1�~H�$\J�tg���sv}���U��e����>�������d�S�B@d*�G)�|������a�k�q��(�;�.�}�u����R���Ud��o���B�UY%j�:�����T����Vө���	���ŚBb�%Y\�<���Ń5����f��\��R�� �19�ս�e��%����1�*}�x{��NgvE�~�����ok��z=�~��՜�EP��s�ƫT˖]����Ur
j6����R$.^�4C�oz�O��m�AvF���I��xt=5�.BN�g���MD[� ��{^��3h�4��QT��6��B��T�A��}δ���e6M7�t�#!s��_�g�*�J	�����f���}#� vx���ݸ3�a�T��@����� Wێ���gA��O��X�k/X��rts��� �w
��k��r4$��s��Ϲ��EVK�N��@Ĩ�+���/�d��|�{�D��J9/{ݐV��A�Z�Y�ߒ�,�u���3窫�M�jmCVv�R���&��1�OKg�z�_�u��7��\9e�Z�@A�v�Y�^�����Zv�%t�a�����*�7 ��m�edSw��C8�#�
5[$q�vz0�P�}����DH #�.Pͻ�Js�&�;c�������6�d)�g���}6�l}i����C	8���H5�s����ס��R�y-zM��j�Y����LT��ܦn_���`��zlڊ����r��(*�l�ef_p���z%��.S��L2��hFv�������v!�5���̥�w�kڂ�apɻ�:}����C.��2����!�/x>̼�9��w�m�nu3��N����^��o�9�Ԃn��d�x_�%B�B���f/�\�z+u��%��jʼ��I��'4��Y=V�({��g%�/`�(M|�J�� c�iV�`�>JȮ�����M�z��%SԺ��7뽔�'$\���n��u�
$���(� ���V����K�����ۃQ�9L��1{˭ѿ���_�� ����tTp���[�tMڔ�j��'_E:���!�W����w:!��d��N�Nb5�1q�/�aC�����s,�U�&۾D�Y��;fR�ubR���-W{�}�Ww�bW �j�9�m����7��(Q=��USZ@��x�b�{g�f��3�z�W�T�����#�ٞ*��y�%z,bܼ��g��XЅ�^�*aָЫL�A3�wj�YM�51�0v����S��������V��hp&J�n9��Ʈ�z��s���`����8b�;2}8��1�-�[���﹉k:�_>'�������U5̲vG�W�[U�tV�'�ӪЄQ�������,��=Ik6�=�N.�uK5ggd��!����Ƙ�Y߭ͼ޽r���ez�'��`����ǖyl�<{���k^��Ծ�cB�ٽU�nG^��FTlԍL���ع���w�<+Jr���\9�1uM���ǭ�0����OT�>�|����c�0���e�Ga�g1���<�v�@��:�6u������f��
p���Jip�������Ǻ����c�LBe���B�aIX�fn4̞����Y�T�k���T~�V���6*���j�B����ȍq0�WTpJw;l�3[`,z���n��,�rQ�G�*�3>0�(�G���%��Kf!�%��Rʿ*��{'��\>��gƞ�� ��=ꑶ�����R ��(F>�����m�u�����H�Ö3O��i\U̱�l��;N' F�<w#.�Z39 Em�n��ev_�<���]��@�����8x��A�\;;l�|Nih�9�����uL��O�3@�٬�d�E��(ѤD�}'�Na���K
�?e%���,�1���� C7��&]��v
�I�f��c$�rk�+�MFu �r��z���S%��fU�H8��;,v⫭I�`O��"c�'j���yPWN�أd�^\!��ج�RzMYdl��h����2	�K�Fhm���1���݅�Pt��eS��}�|���l#Gs RD����T9�;3$�ue����P��4�v
k�΋�o���&0�}���w�Oi����=}����מ�������V�G��dH�Jv��г�&��mu��sj�δibʜ��{J��䡠{�[ѶGaݷ+�X����z��ݪ��TV�kN�.t�xh!�U�/fr�1Z�6_tV���������6�]���W]������Z��L��8��ν۵}�l&s�h:r��i%*m	�{{gLrAGsb�0�����I����<�1�r�^���=j�vhq}ݯ��Z��z��U���n���.0��f8L\P���2T��X@w�ح:Zw�_K��f�a�Հ(��f1:���;c�Bn�)�הc�@n���n�Y�y�QZ���C�1�"k��@	j���Y�B�Vz�o�l�y���V�����Rt���d?lI�Ɔ� ���"/f:x�"ت쳍ܕ+z�pt�/�?0���f.Z�5NW�&'�tt�>�X�Ӌ�]a����_\8~�h��>%�OOG9�1����\!p�q���(� p�W9a*�7U�;�+ڐ@s`�@:��u�I��n�5����i�#OY�~��]B�Vm��"��u�|Ҋ/`��F@R=$Ϧ��҄T-u�FKj���e��n��}Ʈ]ܐ!RnV30�`Tñ*5i��]��櫂p�Ӆi��]��93�u�;au��7��ڊ�X�c��n8�5\�Vs'���v���)k5��x#����1�N�3��m�zn��=:��.�
!;�Z�N"��y����'��"�;�"N��rp������o���QS,�v����퇁)��Ef.�Z.�ѹ�!A�x�5k(v�7�c{I�`�;�����];�9�`Nw[�
�W �2�&P�{)�_LLnay]���W[���ef�yk�f�r���l*$w^6�V�V�T�q��|�\�É�VZĦ��G�x���o�������s�~-ot�\���=y���'op����èK��'C��ؽ���n������♋+/�Wn���$F8|u/AP�`�/��mw�w��V�L��[�ə����bwJx��CE�}p����y+uV�u׈�I��ѹg:��A3��)�����uAh��U��+/o;��W���ū��6�t�/o�]}����8��,�Mr�p�_,�e����CR�J���v�
<uѰ���WXPCg�>B��%lD��hc�8�g��SWp�{%�۔��ܣ;��~N[���]*����m��yb�]�n޺��ǯ�&��s����x�Q�f1;tp�U���cQę4�����e����vc��L3������ޣVM��#(��h|�吣nqfN�;�uz[��Չ�:�`}����G���9�C��ב�O]_L���4WV����[��7_��g�}�e��݋f�6|\�lXgV/���;<���6����:T�pN���7O:�-��tY�]�����^%z�$*��;��}0h6��#��v��M2�����说صЙ8a5�/���ěn������A�e���X�Ϙ�հ��;����m+�&>�p�JQ���;3�	=�n��:76����l�0h�}Z�k)Q���:��,��8���*�mh�@����`iݐ\���!;E�d��F����
՜���Vk[5ئ�d璲��On[]�	$�q����ù.Ҧk%�}2�����'me���M���V�sG�`9=o�g�7N�ܩK�u:�r�h�9��7�R�Qe*ݘL�3vy�:�n�+�%��əF���Ot��S/,����KFҖ�{O�I�x��]2k�E,���L�q���a�H��뀧��0�������p���!���W�'����O�{����<��S��E��\F<���O�����u�o�\'�yl�PY٩��~6���N�4Q���������=�+n��e)����l�C ̕�d�r��r��ˇp�Q��~��z���(���dgh���Q��gy�#��@WqʾJ��(:N��t0/b�KkK+/5`�-�O|v�(9���޳3�
��d��-NäQ�\+N>��)o���N�����M�WJ�QPZ1I�I����@X��f�j��M$m�!�m�Q�J$���ܮUB���h�%L�lNu&�"$ذ��Z��F��QZJ˻W���#HQ�+��IXH5��i$�F(�4&�k%���h��b�FK0�Z(6��S1��Dm$h��l6 ��MI5E���#`���1�
dF�&�1������͈�1$��D�-�)4�1��eFR�Q�3��6���Ŋ#cDF�d�F���E$���I�DcY60[
Z		z���������hj�U���攥�.�N��q���X�[�1�.�Pc�g>V{��S����7F�v��f7�bu����v�u`\�D��1_P`����V���xUX������+��x���;�77�����������z���m����^+��[��w޷���W��ξ6��~z76�����W�1��>�����ޮbܑ����)297���}"$"~>�?[x����}�����ݿ>�~��ţz^�;O:�^1W���|�����_�޼�\ޯ_<��{_V��[��W���Dp���r�� ���:o=k�2�|�~M����B��W��X��}��W��m�v���z[⹹�~�>��T[�\��o�^��u�o��/k|zzh��;xۖ���ߝ5�h�>����p�#�f":o���=�|�ʵ��r���P��CH��b$z��7�7��|��+�h5���+�ޕ�_���=u�����o�~����k�����[�����7��oG�m��o��zZ|�/K���U�t����_~�?�?߾�D?S���8uK�C�>���G�z,�^?o�����~�����}W~v�������<k���7���o��|���k�������^�"���{�>���������߾Q���`�Db2>���1����yK�G���1��nV�����������zZ}���˺�7�nU�^�.�6�x߭�{�������6�x+���y�K|W>����{�y�ֹ������{}/գ~��}m��1o�����5���w����-B�j-��e�&�S���87�:����^ץ�W����x׋����y�zZ����~�ŧο}��c��6�^��+��[w��U����~-�\�ۿ߿}zj-�\���z��ן�����z���ޓo}BW����W��,F�>�>���zom�o������k��cQ����_�ڽ-ߝo����}W����~^yzZ7�~��_[�-�޺�W��U�{������^/�~��
�.k��wZ��@�/r}�^E���Q*�ޏ��J�_o�ޭ���|^-����}m�^����[�oj��K����zo�����+��m�z\����������v�M�o׍���/KF�o�����o��w�^?M\����ƻ���9T� >�#���w��j��77���Ͼ���o����|ޛ��m�޷�}��kA}m�����W-?z�o��|���6�߯�������6����+���/���ſ�Ϫ��f�xg	��QY&��n��r�\����gJ�⾝"�>�lY!jm�V�b����io#V-251��^���͍��jnﮧG�#9{����+ʝ��C�p��U�pz1�p��.w[�J�y�"O�N�A���%�7vx�!�ym�(d�ս��k��W���o�_o}z��>/KG�����o}�������ޖ�{�{���w�����7/�x�-��}�ڼo��^/��������7��盟�+Ưw�����<��H��˞���j�jO�b�P�9�7��yڿ�����W�z�|�߾�y��ޟ����*���zߟ�=m�U�|�y�_�[�>u���~��:�m����@�d�s���Yt�k3�>����}����[�\�[������^/�⯫�������x�_�ξ�����������������=_��ە{]��y����m������������D|��ъh�k��������!H��ſW���'�Z��o׏u����W�Ѿ�wu~/Mx����EDW�7�����������������~^u�oｷ�:߯۾y����{�~}�o�~-�+�i=Т��[���}� >�����>y����Ǎ�k�}���o�s�������կKx�~�{Ͼk���Z����ί^�o�_˛�wu�<c��Qh���|���ͻα\���տMc2�_�oW{��&���G��#�"<���r������ս�5�^6��o?z�c���Ϟ}�W�{o���_�~������sr��}�^�z�-��|����ǟ:�=�u����M˚76忾���߿�?�=�e1�q3*�zts㾊#����G��x���^+�n�����j�����+�������ѿU�������[ڼj����K+���_�}�_�o��x��wkү��r�_;z_���[�wίkx��x�s]�̺5{^��y2�
��"0G������߭�W�_�^��[��n{���w�m��7��m����������{�s}[��s^���h�W��/�}_�x���������/�Ϟy��?{b����~����ӌ�Z�Ox����X��P��"0DG7�;o?{_{�U�h��{���zߊ�i��/�ކ�m��z�|^��߯���[�������=_�E�+��>}��������n�}����o3��6���jE�߾�}�������wu�x���瞖�G�������6�:����7��^/�^��W��/�7z��+����믫z~�������|�叫�����/�_W>�w>c�W߅QB�XT^h���i�w�����`�L���S.q:���܏rT�C���d��t]�x�bW��]`��6;�$��)g2'��=#�'�KT��aXG_L�!1�Ą��7�9H����T��Z �FA�}��U%�º��bǗg��K�;#���}ݕ��������G� Gބ�Q ��bo�������/�z���~�^�7�ܯ{��k�{k�\5��[��x�ƿu���Z����������Ѿ?7�߭��x�����5��[�]���u�����89��d��Z�Ξ�w��.1�#߿?=|m����{ׯZ�}�x���|���_V��m�y���~+���/Ͻ�����ܷ��_������k�����U�v߭����^-�+��_U���s|o>�i�@��U^��=���;U��8}|�x��{������U�����^��W��ﾯ��Z}�o��z����o[x��g�-s�v�u����_�A/���5����W��.����o�m���*��/�h���v55���f]􄣣�~�����s�_u�z^���Ǐ��/?z�?w�����ݷ�����u�o����;���-_���o�ί�n����*����^/���{�/�������7��+�C����fI�nqy8��ƨ�_����5���v��W,~����W���˺��o�o��~^������{����so�>u���n_V������F�����/��_Z�}�x���D��9��mɬ���#��z2���k��_�����W꿗�E��W�zoM�^5���x5���W��O�o���痧�oj�.oKƼ_���5����j�_V��m�|����[�\�������W�����D�%�%�j̉�nc�ɢ���f����u���nWv���|����[��?+�5���k�������^7��o;x��x�k����zZ������^->v����7�ż6��ە#�����l��MP�� �a���~O��ߟm�^���y���o:ߪ�o��W�:�����~~�����/��������okzW?��|��~/�����W���/>v�w���ۻ��?���^���n&"��(|} Np�l]1����������[��W��������\�����|���h���ׯ����_��W�|��n5�W��>��뺹c���~���W���ߗ��W���x����M�y�� R?@ ���(��c�O۲���������_ߟm��ۗ�/���F��}��-�_�|k����U�|_��{����V��ֹ����{��~+꾯��w��_���x���x5��k�}���{Zz�������~>��W�ޟ�>߾w���Б�X �s�\�˔����Нx��O>�JW-Nf�y�C�Z�U�)r8��ƨ�]��8A�%���tK���)�nh��:1�i�aͧ�h�$�}Nܷ��=6�//�zs'P�M�-��#�v�K9�Q�ޏ��#Z������u&�L���(}"C}�����zW�q�������W*�w����zom����������?��-�]��������[��|����U�:�/�wſ���/�w�k����Ƽ|z���l�{�^��ѭ狼��#� ��<�k⽭=v��ޯ�����W�v��-���y���W�G�����}�zW��{����o�߿�^�|\�������xۖ��}����������o{��s�3�ټ��g���Vz����D���w�7��m���_��<�~6���ί�lZ
�k���W��W�v��Z���Z���/�~�kF��|��k��+���������k��~~�~->ur����Y[-�z�ޭ2��s�c� ���ﭽ�v��ſ;���}�U���=-�\������ݫ��ۗ��y����F�z��z[��x���x5����&4GՆ>�>y��"�2|�����/s��u�X��>NcE}{�rwzW9�xh!7�b�ٜ��1&��V����-��=+�Meo����������Z��0���N+�Z��J��њj�;Y��Ӟi#*�QOeГ=��Ms�l��NI�$����@v�Yc�[U��B�^��������2��cZ�z�����tUpUB���q;3湀Ō	�V�-;�= ��+%gL����r��t^J8��}�o沸^�T����
�*���ZVr�hkc²��9�y���1�3:��dj+��S�b8���)��.����ΒtԞd?\�|L5i4�\l��͜�fD������n<�3&�#B����xc{UkQa	G�wC� �X��_;�$�J�q�Hq�r�Qv���v�����L���s��l�H[��fg#k\�{޴i��Cm�έ󘴬y�dqJ�p�>���gpn�.]p
+:�;�GON}��^;��\D�LnB��
�$㤸����|Ȥs=�gVN�V�:���mLxp�)*z\s���!�y�\C��^D`�&����y}w��� �A��OϮ�3�M��6xhs���������I�t�i�5x��X�	fW��p�� j�����ai"��ә��B)k�2[W��{,j���	/bhm��(%gI�K��'��F���F��E��M�Vcʥ�w<�4|�z�ws&��#fm�ޢ�f`�ǹ���b�&�u�;u 3���&V�fS=����:�\9�^w�r9�-g�5�Te��C���Ô �ыaU xҙ�3����pcu�\�Y��c�d�F�8S���ѽR��'��jdt,�dѸm���q�I����D���/d:��*]$�҄8XuR��S�m�ái]WP�'w�3�s�&��*�n��u�}�=4�S��u�s��۩.�!᱑\�I��3egh�c������`&"��ț@�򵰰�g�s4�]E��,0y9wս��L>
Qv���0�q�2��d��h	�Ք��jK6���&��zmN<Dk�x�]߯�Z�6�OY]��|�����9(u�=��j<ͧ�fD��ӌk4;�&\nÇ;{)������>��ەљ����������0����A#\�˯3��@��x�{+�������R�eE&�����&����yV���w�n������Nd*�ˣ�?�V2��L����Wl���g���6����t�'���U�.��q�Ѧω�r��.��[����X�S{�cX�jE���Y�p�v9�2��|Ƨ<#v��p�G��rt]�c&��'	��l��̜p��(S�2�I-LlW:�-���©+�ܶV}M��e���n���E�$�	h�� ��X���-z%d�ϕ��a:�����Hf:�rx�}Q���Ûp��{1w�sLD�:I�Pq 3��G��hck��v�ĥ���3�P���Ӻ�4���c���۸x.K4>��0��I�V�*��5��Y=�c&6�-f�tK��p��wO����&�{0F%	D�=@��� 4�A��\�7W[Uy[��.�Ec�"5��'�I�GΈl�{X��@.lA�D�_o�NXm��e�XN��W��C"����
�x;�X��굒�AiKn\<�y�B�K~�ͩ֙��pl[0]l��[�ӌU��5��U�Om.��(֋�8�FǛ�à��%��]�u��)/�Ҵ�2�m����u�ݏF���8��B6��\Õ:>����_}��0�w�ؖ��|tG��83 l�lo_r�tS1��Ͳ^B5�W�m�d!��֯��\�T,��e���1#�*3�i��D;s¤�DsN��Nb5�ۋ���V�w]�EC���l���L�~t=����Cj���o�������	�[@E��ߥ�ǈ9oN��|�pr����.�GħA]I��?e_�#�/�z)7���C6+I��w�h�C�Z+n�8.v�ཙ��i��{ʘk�
vx�t�c�����z;�ޫ�ad���K~еP!�Jgv��_@�/I�J���U1;�<��`����%YO�.E���L:Kk7�7wx1Ҫ�u2�(����|�k�d��ͪ�{�x��1����Tv�^E+�;�n���[	}�Iy�����.��uN�r�,[5���4��={i����U�q��F�!�e����(]L���*4�j1��?�æ#xR��jq�<�<�q*C��G���aCY�e��@4~����L��BT��.��o;ؚ�����_)	��,��u���ӱ�^(����5J��x�FČ2���X7�'(�|Gv�{^�DJ0�	������[\���1��ұʷ���E�udC'S�+N�.�!�)��G��d�)���+��7F�v�$�5�X��}���۾.��,�V�=�&�r�n�zn!VW�.J(q%i����EH��OW:mʼ���Ǧ�D�p))�'.��RY�� ,=�ީp����%" ޝ�(aL��0�E蹌���
�fWvh�=MTR�c��0�i�N@����eӫFmL�>�
f]�>=RJQ�ǥ�Ɗ:�d?��T�����ޮ���`��P\�
��Q9���(+0�:��a��v���Ď��Z�"�����2�K.?^�]l!�Z���]���.!Xi��^���_��y2�>�r9(%[���i��"�i�w���v�!��zw����M{�?gd�S�9`k�",	N�'�'j�����*�ׂ�U3���joV'�_/����e��ګ�q��健�#46�/�zY=@������/&{u5�`�׶qa�+��Ҙ�Q{�q����΀tpHB1���/fr���J��CVE��u�;+��Q��5([��|O�y֯�3\4⹕�]ī�tf�<�1^W��䢨�N�Z��T�eV���= �[7Ә8X����]�km�{��@�O	��Sr��,/vv(����4������W����e��DƳ+������v��/I��3�H�����t��j��6\���d�]��I�����()Cq-�����8�%��41�1чȩ�?W�x2r�iQ�d1���_�Nq��EhIK�������V�j����2�J�EW+�x:q;2���8�|�ƽ�����ߓ�k���%>���w_f��xv�T��K��bN�*,O�T]���^f|+Z��CD8��Q盞؇��uĺ���D���eX{��,�<U��=���oU5�r�:�\:f���Y��ӑ��c�~4}/�����t����%�,�3��6�����0<=t���������|��9�2�����9��.�m���ln@�C���=mp���%�\x��?\u�&e�����]�vz�39�
�g���7�� ���U�K�2�2�:6X5̑�D�KU
�R�\4dKj�kN�����2q�I.&�O�wIk]��4���Fx���4���2����5�p�}+-t����+68�K��C��v�}]"bٌ����%z�):4|ii���8�K���b��{������b�-����2�Lno\Щ�G�~v������t�z�{�O�4�A>�ّs�N}蚖eٯS��g�X��k�z�L�]^�×�=\���廐�ż%Yb���9f˩������ٸ�9����W9Ҭ�-l�[ޣ�O��}� }ӕ��9�}�X�׹��.Bb�*�&�M��:`�X
eq�jf ɾ{Y������%�
��k�S�~puR'��;���{_t6�E,�dѸm��̌��$�G!�ɘNM�bݩx�G�nX��p��"���_N=�,hXz^\,I��s�&�P2]ʜՔ���q=��u#�a�.#��.a���
�<8*+�i1q�(1�h1�Οd	�=�]6S����/�ok�w�YU�hؖZ,BRto�]���^e�������֩�����0�:�΍�m^F�e�{��ʮ�ɍ�~�?�F���Nd��������V=I��[=����}�+�v� Z�#eL$K,F����p����g�E��.&Vk"�L�U��y�\��z1����������\A,�j9�2��|Ƨ<#w�B�7'D�C92|9����ؖ�dL�^&�:	`��s+�.�P&��p�@�*�e#�"���NQ�� ���[ת�Dΰ��vpQ°�r���p�kэ�>[֩�i�=xZ��R%Z�3�Gn2(��5q'S��g{<�꩟u^��DF��P-�7��P,ü����� ��,��-����B�\��d;���k��]��!(��zUݲt:d���0�}��C�/������(���Y�����7y/^>�AE�M�v�%�or<���0��$�"���#�w�@�-Y�̒�.(�oG,i\#DފV��Z��={�s���M�ǵ���؜�e��]̈́Y�dh�u���:˂��^шQ<�9��l�|B9i��	���/�|n��ki����A��J���YW�M[�)J-���Z�n]��2�%6�(��烂�]��\�Y'pȷ�o�eR-\a�g.^�p�m=����n�!�����I��n����&Y�`�zA�Y�a�3���ҷ�]$���B�nF.>�a�I#�l��0J]3��f��N�u�Y�{�{*�s�l1�\����n�`[��rx��0Zy��\��9:����:�wB���O��3=���oAS|髢��y˅�Y5v Ydⶫ�v+�=�1u<w:� �������ö%�_<�!t�.��q��B�6�j������A����{��s���"ſ./����7;7̑�����ذf��^�F�TFr@��V>��u'��U�gms8�F�7uCwH�IƘ�l=F1/�b�5y9�z�W��#���wx�v�Ë�;�g�q��A����[8۽���Y�W��n�ݞ���Հ�FP̈ۊ����t+U#N�Tf7FwW�n>W�C5T����|��;������ef��2����"��.l0�3%�o���
٦"Ͱl��;��_	��ek[�C8(զ�E���:��5���)ї7e�j�ޠp���֒�
����p���#�`֩;�{1Z�����ȝ�h�,�f\���&}n,j;}�*Z�U���2��L���0��S�%�	л��m�f1z��St�"�U��p�w�bv�e�eJ~���Q7���*SW��RP�� �X٣6f奏.A�PX�/�{���ݝ��D�t���(��Tfqx�nw���g>v��v��Jξ]�l\���X1���o\��J[��E�֨�@�B���1ꇰ�=ʋ�^و�x7�U�a;u�H���0�
	GB&�Q-��$��Z�
�D줮���r�s�E$U4wݭ��(���c|('�! :�;�t��o(޻H���5�����Sm��ݲ��q��gK߇\�9�g-�̘������{��\�{����b���#yS<��%�Q��C��%��>v��XC�>Ϋ���QB�7:i�#���pJa{g����8�h�Q*̘��`�ѹf�#�S�a�2�K���5U�q�^���D�eլy��)�*bӈ⩤�W��͊l2�[r��9u׳��K��]�:���\�A�^�^Y2�w�6\�K���{� ylEI`�TIFCF�2cI�0�i-����(��F)6IRm&�����32`�K,��1���h��Q��4R`MQBF�AlQ�!6� ��TQ�H��hɠ�6dP`1�6,�Q&#l��F��lE�4���d͋�#�h�cQ���	��*1lE��Q�E��b�F��b�F�����6a`�1�3QDPZIc���b6,Ze2��McFI5	XCQ�6�F��5I��1EHDEE�ca���A'y������z~{?�|�H7׌#X���^�eS1��N��٦t��iEc@���o^�R��*�Iw��O����g����}� 
�t�Z�S���я�;�ֳ���J,�3�|�! x�B�ɹG�]�����M~]IöH�'7=rk(��׾���m�p8i�w�f�ѽ&a@	N���+��_5��9��B�Q��?�R���G�.���N�q6�`���4�J�� F&A��4c�hS�7aG,=5��w�̒!��'I��D6C��u�z�.�A�S$�2h���!5]5�m�cG� c��^��e3cx�]N�|��`3L���v/m)�G��0���|���&������$W���Ҵ�9!��d�v�,�/n!Z�x#9�%�����U��)V;�l�<Lt���}��K�
���o���7~�B_+}=��faU�����͠�8��e�N�s���u �d��+�(�~uW�H��/�zt񢅯ghEX�
�j:���k
̱�_�>r�+�T��\hS�<M���	�z����Y�L��/Ev���1�,>�L�����zM|�1���������`�����0|��f���Ơ��5��M�S۠-xA�Q]��P���F��(�"�m����|�O|]ř�8���y/�SkPIe[{��5�=E���ړ�Q����D�`�t���\..u�t>����t	T�8��U}�}��Pάj7�>.p9ɝ;3̔p��L_5p��S\�'EG�����Nq����W��9t�/����&�z��f�\-�K�OYA���.��*�/�+;'�&�u�0�R�r��bi������B�V�+���4�(�!Ǵbc�Y����q.�=��Sf���\f!)H�E:��&Fq��2�ـ#g��x�+_	M-҂�rz��Ǐ��v�[��m��q�;Ѯ1k�t��燕epY�(�<IU��|a$���7סo�t#����O���l�PR��>jK1��:i���T��N���H��;��NE���l=dt~|@�wU
l���aq�m\U̱�n ��;N' F���!q��+�{�\B��#�Ӛ7Q��C�"Β_���@L����q[��T�H��q1�+Yyh����y)yԧ��(MH����+X�B�w�4.)L1�:XW�\~�K���q�cVTt9e�r�pg�����s��쫀�;�f9��1�t95Eq��ΤG��M?0�$������L|�ʳ�*��S�Sq�Xa���\[=I������\��\&uz5��o�Ծ���)�|�t��q���5y{7�fY����/oZZ�/M�r�������)K��i�?7��bH�:��u�|���{)�f�g�\���u�w:����ﾮ�Ѱ�hay�$!�?~��2^|�5�"�
�Ωi�q�(u���k��E�f�:�WK��6��p�ƈ���Cj���1��健�#44;?�d�@?^�>b���J�T=ߐ�oJ&l8}A���u����X2�N�nv`u`�h!���!��C���Т�z�ϛN��x�u��V<r�[�<���S/�,�%3y֯�S0���8�ekWq)t�H�ڼK��q�;�8\a��DaD��;�~h��7>�|��uׅכ�U�`B(��3�N�d,���,�z�3Fo���˷�q�$eWB�����"*U �������:�S��%&�îۼ?��<�g��3���7�y\.7���ŖJW�I:!T'�	K�׮^�y�V��*����!����<��ۦ#��oJ�����R6��I:j$�7�7mÙ�g�k�ŵFw�&;��gb��Y]=9��\c�l��T��*���'�!S��5��Z][�L`�	�U���~�0x�q�Bk敾<�g���֊> ���m�RRwf�O��p+�pW!�26dj�T�j���pͯ֦�V�Ю p��&���/ c�c�8�z01\�q�"��pϪ��M"�1�����R�����oۑ�����:�Zve	$j3���`R�X
ְ��'��0��V���N�c�_}EZ�W.���6ѿ���t8LA,	���������L�s��-�/��H���49�H�淈U��#o���L1EIF�� oW�@r-$Tϧ3�҄-s�a'����y�|0�����ϜnP܄븛���x�g�(q_B(t�ɭ��w1啹D���f�JW��\��fnTa�&��.�?1a����-㸚0Y��?$k�@�L����
��ɛ�#t�?���*!Q��C�����E��X
�]6�~���ɬJ3�
�RG�lا�O3�ozW�O��mTH�Y<ɢې5���ƨq��>�3*��ư�݉$���W�[�<4u����=��TX�r�j���w�a��x�L����T�rW+y˩d{@�UgL�V�¬�4�v�
�s5�6�y�5/O�3�m*~1�Gĝx�-^n;wMp95up��F7��++���bYh�3	l���yu�jG�˂��M٪u[����N� �5�	�p����ct�{u��F��,�ۃ0��j�ؗcjw��^��|e��5�r�p�t��oeBiK/��,�2�62��\�=��a���բn������x,Gے��o(�S:9����u=ǔO0���y����v�ogp�8�̤�D4�Tj�6M��%d+��^��@GAF��Lz�`
�G�D}����&5p�v!�2�+ L0���#��6J��j��p��������O��ʡ�V�s����M��̺�qN���h��p�w��<�퇗�9���iu�i��Y�,�I\��異MàK�KڪU=�	��?v(��Ea�岉����[���
�R־���x�����
��-z&H��_Z������ ���dؽ�p�5
2�j88�W�ֳ�W�	:��Ht|���{lw�����+'x��hP6xXp�SFg9�p8i�w>%�F�0�T�I�!�&�k��|����_1X�\Mķq�˺|u9Ѥ���eE	�����B �J�n(u{Q̐t��W�r�ps���QY�D.5xWԓ��:!������ .lA�k�ܧ��*�aԻ=���m�����S�h���Ӄ0l�cx����c�0�J�ќ�ʱ�t��'W��${"���J��Հ�H��a���Zo����4񃯵��=tB�Y����)��-�o��#�g���;�8�oj���|�k"�ٚMG}\6��ѳ6bԽ�JW�߳N?9|���os�;]S����Y'472��鹏{���Mum7d�Ak"_�tF��x�;����y$��?i�ޢY�~�|�s��0��Yd�����Ajcq� Zx�t-}���4�k����\�\3k)­Q8�a��uq���{�����nX�9��wRd�v�Lw\@���}.s��t���(�ټ�aS��HGf�C�XX�uLB�!�_()ٶ�z�B�Y�n����{�1��+�\i|sk�eM]��8�I51�0\v�f�v�؀�%LCE�������[(ty�^�������ǧ�ʭ72�(�و�j��3��\
�Kwl�*j���M��h�Dд���gix:�F͓�K�����6%�{U���t�j�<�ּ'����{�/_�t_J8'�^8j���`騁GuA\#�V��Mg1ǬbcݿZ~���$"SGuo�8͇HE�r�������v�\eC@V/�����S��-�ڞnh�ũ������R�"�sv��,�-ތ�\L1��:m�=7�8�u��\t��⾣�n��ֵrf�2Nj�}6��"�o��<wct��}����OD�� ��=ꑭ�|�I(Rm�AB��bؒ���]]j薚+�=��j���ib���=ý���~Sbh����b�Hx\��!�у�'4UUd��W����JRqv��i�|�>��N䮹��8/$���;��@roϢ����^�P¥�Z�������<5i�Zݮy�=�?�U}��US<�w����\�$�&�D��G_MǕ�qW���ๆ;NBrmG���)�ھ�MX�U��z��܆� ��:!�$a*�P)�p\z�p�N�1��}��.�-�Qx��� �#2�W����S�8�>�\������S�*c.K.?Z|7"�'"�)dO�_Q��Hۭ8ꢋ���3_D�UQ�r9(%[�;Z8<��g�ҁ��;}u�փ���T���V�!T�\�2^@r�בDE�)�D�N�2��uv%z�Ew7��9����1�&��������mUѿ�2�Ќ�ۂ��&:Y=����H]��J��
��U��K��ø�[��W��1��gt��I�����ʲ�
�z��2���� �x:����pa�,��'�St�_].'�wJf�_Șvca�̪���p���ԅۉI�L�;�Nxc5��0��j_ƸyUV:SV�Α��n}�H
��k!�w����VV@5]�im����W�=i����.�|i�ݲ��	aU�
���N�k���
���,�H'슼L��x���;�KᷥvT����v9�;�eb׽�e��<���)��՗�Nބ6�,�1^2�x{����b�oY�(}e>��Zf)�
���h�0� EVcd�.��:Ty7�0��o3���
(=�EO�&{ι@�D}}��7ʵS��x`���E�i��%�g��٥;���T�,�����N�MF1}fW]���{w�q� l���]2�ܑQ�y��LG\�����>�hd�,$�F�^c�-��+��e������_
F�j�����ӑ��c�l�}(c�[|�]Y\���N��6�5�	<���u�����0x�%�OOG9�9��k�'����}3���U��<����C��,��&	@G��?_�uI��n�9���9�1{wh�!ε�%z���nF�������p*J= � 9�k�#(��iU	|)�1d��r��T�lkv��u;�ý�5��'�븞1���48�"�m&��=fc����a,��`9�����X���k� �P�V�|��'�,2u�Zv�'Lc�ݦM~J`tS}�Y�M�+�3Խ�p�:�Q�����{����˄��M��� ЄP�@�Ӝ׫�aFd���_��}�G���Ḭ;k�8�͕��>���Q"�Y<ɣm��g��&m�B��:
��S罖�W��2=9u��iHE���,�i0<F����C��)�ܼ�\Y�\�={C���H��g�,�-���-�6ٱ��X����L*�0��?��N �R�Ǹo.[j�ڌ4�.=l��3pK�vrEǏ�����ﾈ���b�	�^��ѳI�وe�|>���U���yᰱ��M[\�I���ܳ�&�ZZ7kY�ws��"|���{^����0P���F��^Ӣ}Y;4���fJۿ4�$:���GU)�/�=��y����hߪ%����I̅}��]�a�B���}�t����������@���ܩ��]o�����w#BJ�^'2|Uu�=}�0Su��Lܵ����ѯ�D��
3-��a &"�u�GS�l����o��A[�y���4�ր0��Ҹx�	K��,�u���|e=U^�*�/P�K,���<��y1�xF�a��D����X��o�zx;G�U���	1i���ҩ��U���_k��>Q@"���٩�R�Hv�8�!�̣n>~��O��^��E/爃��
��עd�ϕ�Z�̮�3�m\���ש�ޞ�����,v�W��5��b�!1�'��q"�.aq\v��L�ɼ����v>��RTn�1@�ō�ь��p�1���N���%��{ �(8n�	��;[Yq�Z��Ц�⾯W�GW'ov�(!�r������ޡY�����i���*�����c��2�ҹ��j�2c@�//#��5j��s3��S�mnb'�I��A��x��*�'�!���|�L��,3��4i?L���-1o��i�π�����Q|��O��^d@u�
����Ku�zs���_�fʂ�5�*qGw ��o�R��� <�`��� B�з�}P���g6QyX���d�k(9���c��I�X��vKO,�{D��0V��PK���C�Ҩ������p�,�bco�i���i�>�I�����K��ć�Q�	���5�.U����iޮ�7|��J���J���0�gEm�r/FI��]�7�s��WO��]i�u�-}�<�J]��O�/Y�N���]ܞ�j���y|��癹Z�]���i��A��z�5�9��S ��~%��Ԛ-��̵-�{O#�ގN[w��J�<P���u���ac��е�e�9Z��!��B��x�WW����y�&T%]`�.
�qYM&0E�����[�R�!qm]D��ۜ=?V���G�p���#}�f��G��Vq��%;1��WMs,���LlJ��/��m�U;R�.�Г�3�8[[�>!��y7�n�_k���6�=.|o��Q��S�׹ʛ�P֦�/c�6s�6���d仧�T�:�Ӟ4��/`o�T�]�tf�28�K�u{1)C�ݸ�x����0t籪7�qRա�x��ž�f�L��ˣ����ո�v%�d�+En��y���L��u�HLG)!i�P�#]q���s�&�_j3;�
;.U�m�PR�ewun輮�!�:�'K�L]Ij
�NcKǫBqK���][P�zU�+'[6��pFFh����0N��5�l�*�07l��<���%$�s;�:v���@c���O:�Ω!���[��;�;����8[����+{��rۧ6���r�N{V�9����}>Q�w���uy��v�j�0�c�^8��Xi���6�C��Y+�M�7�m�K���	�,��o0�Ssu�Nң`^�X]���%^��,�f�f�1;��M�DX6���y:�ٖ��x�Z���&+T��a�Y���h��KlV�n��#*I9��N�8�W�%�H�(�%�PMa��=�0.x��
85���h�"6>��O��q�t���1 �K4��G-P����i���I�\��{�םW��Ѭ��������S<~��M�Fiۻȷݩ��P�;��Ј�q���ݼ��Z{�s�ђ%=]Ǚ᧧M5	k�]��gP�{0��7�kF�4��*�:cӏ:D*�2��j�����(!�u��a�N�{y:�yٻ*TQ���%�0�����˜�M�+�Uk FC|V���P)�&�9����r+�r>����i����Ff�#7��\O�=�||Mꐌ�n�T	^WA/;YI�p]N�;� �#�㉯6�ݝ�*��=R�sI84�J۸���w�y��JǵK�&�S�u�:]�r^(w��{��� �X��5{�z��CE�p�3ʅwD��ge�|��gz��+����[���]`��"2�:�:���J�l���9�+0��Ga��z��*daQ�+�}��Ω]qls��{6/v��вn�klk�����C��pc#������K/��K�l��7��^�:2�qXٸwD� >:�Ĥ-3}4��W��x��Ys�i9�v��۫�j����e[
��\B!5�m��^���x��")P�x���8�1�}��!Z�g)��o^o �����CL,K�|2���W j�"Ճ�`�����;y�K���)�h���Y�M��L�bD��z�2vs҃v2h�7�(�+umH_1uˤB��ީĎ�T�{��$9���#Wu�k��o���yLܹ!��_�ڏ�56`�HI����x^�x��{�G�=3�9��dѺr��"�+|��]#�8S6�[�9;����Ժn�G�5��H��o.7��L:S��k�u��Z�L��K3�س�&KjR�����f���o�k��֧d��m8�◇�BG��[�PV60Qhчu��!$X��v�E!E�a6+DfljE&��")��l]�FŌ`-$lc�60�"h؊Ơ'w66�hh�71h�wvUr�nlAgv��\�DI�.��\��Pn�Ƌ&ب���sk��+&9��$`�;��IQr����9�Ph��s�nv\����H��&���wv�r-��R�6M��đ��$�6�(�ܹwrW,A�.\�fZ��7k�;��A��;�H�Q�v�	 �9��2PX�u5�\�K!+��:.W?߽���������=&�^;�pgrLo!'���sŕ�Cz��VF3�5���c�zȸ�z2��G���
��8��N���W�}UIn��6�{�x�N�=�k�f�X�oՆ����Ep��XxJixS���*�+}t⡅�$�!K�c���_ �����gTS��dg��R��f ���ə3ԃHR�[�:�8�5��y��S��fD���P���`q�&�r΄���]pQD���VV��s�֮精�O�£Te2���%���J]�Ԗcq�|��F�U�8i�sv��9ñm�+vI� �<#P#��C갸ⶮ(�;�|\��2b�Q��c�g��^�����OU=sJ��WR�fe]��;���0}C9̂*���Ưާ��o�{B|��+c��Cgt��*�[�*S)�O'ܑ��戭co�0�ׄѫæ	{IG����@p�5{�ga�\vu��C�����OJ�R��:N��G J����:G��$$�G,�+'m��Z��b^�A��d1a�O��5L��1�",�"��vM�Ľᗔ4��MC�隇:�iȣd�T1���mMQ�d()�3CC��|NlY�C���v��Ьv���t
{�86r���7��D�'z�8rlX.�C��r��w����y�̻����RuE,u�F�%{����<�oq��e�ּ�G�s�D[��^nԹ��xm��/���ې�n���EdƘ�^n�=w����7�n����H38�P,*%�X�n���ţ�	Lh���rwzr:іX�X���������-.�G��ڣ^�v�M
���&t&"�{=>�k���F�WW���2j�ZW\���=E���P^&�RNT���ɾ�@L=�+uFuI�n�K�Q���u�Ys�w9U��]3�d�a�4�*�/�{ON'e�{�)�jo[}�yT�������"��y�.S:��}�m<��3Ǣ�% ~�]r����t.�t���}e�"�Ǆ��@5���c�1�nuE�b8����J���vT��������z�'��TI���\�ra��B�w8�zr4���u�Q-S��/���5���;�����=@�iV�t�����J��G�ژ<k�
M+|y���hB�X��ݲ�w�佑[��.�2�P@�0J8�0S�u�&e����;$�F�bbs^�(�Y��ƭv�߹����+�uB�%����ZH�N�U�Α�=X]'��/�f돈�8�c����jvI[#��!�x�"����4i�]ˊHK����J୚�f�mX��r^-��fz�3�kd��w���ܭ��:C$r�mE��˼B/��2��*�˅�^:�6%1ϝ�໡�'K`MܧO��y}o8���DG�}�y�-�ƨe����Hh)��@w���u�M��q<n(�?T#������kH��%��s��;[�:��tc��Swˮ �I5h2�1��_6�@.�ĈÉ����Y�j&�q����;"=�ɞø}�3�	]8e-����u���E�1`�+�E�����	�}QO%�f����>�aʩL��zW��_����S&�����`K���XgM�����M���J�P�=0�M�>b���~6������]yp��[��_J��.'gVه�~Dչ�%{�!�}�Y�i�5P��`Uc��YC>��ɭ�>�����vf���J�Z�J���[t�!s�����,�6�Yh�3	oM��5�o�K��3�N�j��>����t>
�< �ײ�%q^8�~�*��ct߷_�둡'ڼKt�[^�=S�g"��WS��ޥ��}��M�`�Oo�a &>�]d\u:��F-���p�����P�+��g9�4�d�F����6.R^���[*�7�|�U{�;.�O3��<��숋"�[;���-B↖Wl>�J�3�[l����\-���\���S��7j3��"��n���G:k1����5
"5���&&�7�I�u��B��ۃ���q3Q��--�.���mQ{�K��ͨ���m�+��z)��A�˻;O���4n���[��� �b���v�'��J��TG��4���+c�����k'`&���G��My��ȍ��|s.�D� ' ´��"����!zx`�ǩ� ���P>��Z�J��K7�S�)>���R�)�Kc����[_˃�3"mT=�5��b�!(�'_�p�@��q��Ԕ5�~�y]a�`�lZ2���� po���0/�9�p0p����ʨ+"�Ԟ<�P`���zÇش���:���p���\Mķq�˺|u9Ѥ��eDE	h���`�ցݞ�ET��x@b`D��A�ix@�Ǘu}I:H�pCe|^Vr.�9����ۚY�>>�ް�`�Q2JR}� �g�W�V����oS>���op�B�~i�r��`�Ma)��`��!Q���V
�0Ĉc��gJ�c2���u\���-хf搞O
��vh�b1���div@P�3���5�}1i�s
�e�������:��[+�8]V�s=��i�y�tGc0/��1#�5+*�5�����֟H%��C}��#9�c��Oey��>/sqDff�b���c=i���w���*�Ƴ�u�i0U��S�q�=�{γ��h�dS�@S�^�G���e^,X��7S��'j�<�@� H�=�]d�������P}��q�8��;ط�w=���̼�պGm�z�c��oj{�noq�/���:S�{�v�W���S/�O�Ϛ�ӫv:j{�h��%��:��w_�.�׾�3(��DM�T��끊&/�w���%��"�ھ�s/���[�`�o����ܢ�)O�Tz s]/+tW�P���L'2V{tb�k�(�\8������Uٷ�,�[�	0����Ϫϧԛ��>�\9��t�*����J�cc7}	���΅jt�α��{ފ<���y����cTg��{���e�R�4��ỷ��M<�\���1�Cz]eܷ�o������W��������-���h5�c���*�z2F;{�{���:�%�<0Kj*_wn|��_ʟM������2�����2<
�18�8:ZF����"�>r�5�;����'Nr-�ŸH��:i�����V��'�a��3��Ɓ�����,Q`���-,ѣ��YC��B�i5�<��*j;�f�c�����4�U�~���Ѷ�iP��ɑ�ܳI�3D�A\��9[��v�=�;G��+���X��G��tHG��|oo��?}G�5�����g�3�cO <��7�.��B�d �騉Z�U웜u���k�=֮z�ZG�2�;LTb�f8��:���������{V�������q^)=Ӈ��i���4*2��CA�L)�R�{�'V�PQ�eK��^D�ɫŵ��yc�4ۍw�K�"qƚ�9��S����oo*�ٗ���$盕��άp�6v��L���(����ˉ�Hӎ{U����E�����y_O-{���'cY��f�:�L
�{�9,��z������Dj�S�œs�'��V���3-�����7=mU���sտQ��Ok����+*pK(���ӯi~�e����Yv�Ԅ���� c��ƅt�ld����f�y��gj)�驭݂��g�U�V5Y�]И�T��T�D놣K\1�����4�������R��ي�}ɓ�z [�]5�ic����=�l�9|����K{�kb˾�<V�%�{��J&�'�zvf�{�cv���sG����6�׭�	u�	m;7��7��:е�X&v����R����O�����a�/�c	�ݦ
�YÒD#菾���Kb˄��&�`))L΢K�PD-T�7}��m�E�����z�������h`�����	l����4�{�][��Qh��y!(Q[���9k6�@��}�?�p������A�
mi���ʂ��Q��Z�\f��r��IX����z~0�-L�gfR9�8�s�YN�_b}�[JýZ�`v�?��4�S�.?8���p^����8z��K#�Y��M+e�p�����m�ˣ(���8��|}ZZσ�~��o\�|-|�9�M�v�sX^9���+�=+�GWKU�ྷ����T{-��������LА��zp^��o	}Nf�b�:]P��%�7�{<��Y��~r�󲠼"���i�I���s�{��{��*-�_7���dF��k�f*���Y�b�e=�g,C�r7�V���gq�z�J��ykʨ�r�/8k�X���n�'$�b��C�[�+�7R�ws.X�J�G�:�E��h���'�ç�RzIۦ�p�{%e���w��v{Q1�>����:��W�B��c�8菾��Q��9ܬB����{�^��~�'}�fT�;��K�F�k�K�[�=��)Sw{�%�W�^��q1�ӸS/E���Y����eٸݺy���Q8�� -�F�N�*��Q79B[p1D�./�/W[kzX�u��$P��vv�AVNU���!�@��s�����=k+��+sS*iй����[�[0u�����v|���X�wTg��g�-��w
,��&��+��v�U���Zl5��}r��+:�]�W�Z�_<ف�6'"�cC�}�1?-bG���%(�}�����1����m�(%�v\H�uum\�}n:��!�V��*�T�BN��5��mC�9_Bt݋<�n��ۗ�L�C>�p_٬G>��˖����u�v�r���q@R��7�)¼�/��6b7��!����w��xjM%淬&�v�Ӻܹ��ҫ;ݕ��]zv�;B�~زԷi���H�����q\�R{�`C(�[�t�k�C�C=_����ڕ��->��rк���P�Q'Z�Q���=f��P�=_���i}�6_d��1P�,!�6���T�1�G�A��jLHZ�J�c���De1�w9�.�cyzѤB�����O��ne�Mo���J
�XWr��K���ZÇL=��)s�_�t6*����^�W�B�����=^�&W(�˞�m��{�/"9�&�q����D\G!�-l:Xź���}���+&�lܬq/�j��t�ԝM,p�p6����ȟ��ޘ ���=�2�!C�R��Q�*yk��{X��r��k�5�o$u��;�X�Û��)v��-����X2�S���v�^I�ZRY�]n����6A��-��Tu�u��]Ǳ6GxoQ7�<���+pE���,�j�+7\6����9�]��\�9BT>Z����hW�λ��G�1�/��Ht�[p��[��gYڦ;���ZF�ol;��9�����C(���e��cb���\&�\�{q
s�M% ��X=�Z	�0q9Z����j�^ԃ�ŬQvY�z�p���)�:����؞�G98�Nޅ�0׶@�_	�w'{��L�Žu�5D:u������r���}�gS���)K-
�Ǉ���j�U��B�E�Im֠���v>�MW���ꧫ7�BO�*��5�Z��ATB�J�Ky���m&��)�]Xb`ø5[�:�oBS�UPgݮ��.�/~T�Ƥ��'�<��=��W(���ۡ�nu���IRB�z`��&�T=�j_O�W5�a���GB�É%�c9Q��T�)����5�C������n>�0�>ոԞ9�l�v�q<�j�����v�`m��t�B!O��᠞{5ٔ�ڹ�K�Cn8�ֱv��skM��i��þ	T?�#1����Ӂ�Vx���YY��D���/�ǓY���%-s�0���q0�
��zP���:��N��1�U�;��ŵ��ycsPۍ}Y(ڻ5=6�)�Q9��x���li�K!�ȗ�Q�^꾌U����赥�q&����T�w!K�Z6�9�Tk�u�t��|[�9�y��qR�B�m�Zy��N��R��햍�x��X2�"�AD�T�JvG!}8��=�ɫlQ��_C(,���v5Q�u�z7�����zC����*Z��-i��"= �������bR�(����#P+�9|�_x������n�5��p,홍�XϝK����f>�+��k]��S�Gn���g�=+{�Wy=����0,fu&;��%�m��]u��f���ƭ(���e4�݇v������s�oVxch5QF�!�H�wT��@��������H�I�v|���@ꮘXgݍ�b���dЫ�]�8���"GN@�B�rX�N��Y��$�R;=�د<z�{mU��V���Q���=&�`�f]����~�nv^�S�ж�}:)���Z]��}�	�x���I��&�
Π:���]#�U���q�����5��&}��v���.�]�|4�%�;s��X��C���@$�ˊ�+pV�Au+��2��ڥۢ�b��,�����Y�_W����t�+����S�;^J(wt=��o��Qۣ�{�/�b�/r9�*A��w����ā���\��gZ77Z����J�a�Wi��.l���QΘ6v�o�A����Mq�]Bۼ���)v��G}Z���y�����}z ѵ���/5�����G��W����#�򜐕�m������wܽ����r9�8m��,t!J'։�x��^2�j8�[�$�Bl/�弅���yu3�坮r幉m�tVp����v$�re�8��[�Y-�h��Y�v�wqm'�;���6޸۩O��j���R���H5�Y��k% G��l	h���0ot �|����cI��4v_f�w��5�1�kds�^�w�%��>D����ە����i�V�C���2�y���<��=�V�}u�J����h�/y���-:��H�"p�!�PLdί��GS�.�#�8����C�/f����"��MA�;���=���gW8���08e����ъ
ojX�5c1�R�}���9sq��z��RO�����Â�*���w�Q�î�����MZQ�|��S���C�{\C�.1��YI�8�'W�xwt5N<������zu!�8�!K��pD��r��N>���"���
ٓ8p�u��Gt�]{�/�r�/���2��ǚl�̼�^ؽ��-�zIȾ�e� ��$�gb������\$������Y��R���n�f�dػM��mB2�\���O4BL������n�����V�x_�c��ܷkFm���5�ED�⫣Z�UD��c�L�*�P"+5�Vk[�FqxFm�E5h�>"���z��/B6V���ֻ���y�`��������{v]f�s\�F*��.�	j��<�u�me���g{u��ͶXB8Mz��ײē��\:��Z(
�
�������͋!Δns�(�LAQAY˰bƲV�ƣst�N�����Wd��\���官��b1wu4ˑ���˚�[����s5$D�����s[��Q+sX����A�\5rۛ\����nQ�&PQQ���,lE3b�w`ӎ�\�V�L�np�(ӜQ���sccQZ6L��6�E�Tm��-��4[�p�k�*Qc`�nRh��#cr�1�mr�ѱ��t�ܹ��ͮS51TTܮmE�_�v��%N_m���Z�m�4~}|7djG#ٲ�Yl	���v��Nl��d���H�pnc�9i��1��~�>�N���j�s����e�n9�}Fy��9��%�z�%g<�pvk���r��}h���s���)�	_f�*Ϳ�f��B����ұQ�
%G�;��O����7ri���}%>��'�!]/�-�}y��1M.��x��J:i�g��J�*��:w�.�}��\���m�}���DnnƬv��\����
��d�?���9�:�]-�E�n�...`\�GL�{AV�en�s��,Z��|��$����"�!vکe ^<���;ٰ�xW���s��

ToIPbp�.W�c��s�n�3���h����X�dk������J�PS�oЫ�%�����c��_+��>���}��[��ĺ�t���N�\�[��Q�l���+]�.�2�I�l�v1P�ϯ\�[�ؐ+[��P��Ƌ�}ҹV��Vt%&�5d�n��a����X�y5p���x����G���'����a+�iB��a��T_L��{�`C!#�����e���a�s����hv���r}��l�yA��B��pk�����Uv�SŐ�y��������ԭ���Kxer�4����M���r���s�U�|�W�y��.��<�1z�{mR��F��Mu�]s|�R�M@�엫X��7�ï<���'c���9#S}眓�{'5�w��hf�]�㺯m�V�3�ڠ��Y�������(%2�ţR��w,u=����n^s��[���ۈZ��<��<�*n��P&bsxj8g�#/�J�_�⨛{RV��S�Ӹ�2�\G'�ds���泼,;�X�{�}�qZ�<�I:���G���_������S}��>�1�/WX�ٲ�9W�֓�ǡH����]}�2c�좮�Ĺ��X��1�kq�C�q��^snb7��f��H����{zR�]�j���z;}\�p���`n�#��x��,qe1WЖ[m���Ϩ�y_F��T|G�*o���g�h^}N������BS�J�oI���o�uw��z�����o���w��H���a�PN��|/��F��#�)[@z�SEx]��:C�&ÀI����wȫ�ҢAf�sW� 0D�Qх�����=�����[�=�(+I���cXSk�L�O��v�+uQ���z��-m<�8��#���cn$hy���k�#9s��	J��)<����ж���鷷\�,5
�P�����Y?�&#�m��Z�h�ݴ=��w�$k)���-��X��s�[�q�.|��(zD3�=��zes�;��)����NB}v�E�)D��L,��ޗl�ЈS�H].�1=�/ᩀ�t�3�;�T�+(�����o���W�7�LGR;_Πm�AZ�־�����:��,.1��a��:���w�9	��l�[9&Ĉ8��"��
��_�u,<�v/2b3U��u5)�o��z��Hs)�\�Z/�9��E�FVu��U�N�}ܲ�mF��ָsQn��[��e�&�/��Q[[��х8_��1����X2��N�k���^%7�����C+�l�bt��CXo����{ɑ���aj[�V�~u�[z���;��W��"����D���癟oO��p�L�c��v�s���NE4r�ytә�p.�()��<j*_,���2�zy�̠z��]��c�7	���*%�C2>cg1QM�n���-�����2��<��VԈ��T?_5�w���Z��,NB�y��We漙ֆD�]'�O��-ұ�K(�s/֖Rߦ�]�3�{�N����Z�����e�.��y_���m�f�zԼ4v*�e��Y{D�=�S�������coOK|����� HӜ��=�K'��X/�)�I}S�*Z�^����y�c|���_W�YrU���U��J�x`m�p;�q{���t�Ԟ4õ�;ٹ�b�EiW�������Mcv()_o���ǳϡS��[�L���WѮ�q���n3i�9Q.�B��#�ޓ���M�R�wU��}�m*�;9m�SJýiݍ��ʗL�!O����ܞ�Aw�`4�3�-��V���_�t�����M_̾�gn�>T��<Z��&��@:�L�38^*zn���5�GÌQ�pL���{m׽�Җ�1u]�u6�締�#�,`��\b��cN7pT��E��8t�{w��f{����:�x�����i�HWReYl��p"��f���\6]S'��jAvCE����n�qf�3��X�[���Mf�\��Z棚a�n1�#p�V��U��](��t��Ͱ�=�Χ��w<wک��71�a*U�b��.��H����ՄOi��
�w{8��un����Oxͮf����޶{8����hkw:��}�t����ϥ�����g͵����y���<]Iggu�K��k:�-}͗|$��U���c��z�%!��`\�Jї�&2�h�	gm���)XD�I	n��眳�ď��ʉ-�b��HWK��Kz�^o��LSj��߼z�s�M��<�^ϗ,���j�kU[�>oe��<�tt�N�^#�J�[��_�E�0�g]�D��Z�$�揸g�( ��C���R��j�4��%���:�T���*��<��9΅��ح�\��C"�mq�8B�G��:��!�e�G���}A�6�kSh)&��ά5Ne碞���׻s̻̭����c�UN�v��W]ݸ{��R@R�q�8:��uZ6��ڋ��$�M�C�>�"�;�(^��/82�0{����\O3l2��[G���Q΀�,�w��ꆩ�YP�-f���qQ�?	JG���t�G���Tav��+�P���I�+kq��M�J��>s�Og���꒣��p�I���/A�w@�؟C{������񝨗B8�[[�y�������'�fF����k��˪!o��Lkh<b�����~�'!5e��N�w�k
ڞXf���U�2�\��GH��?�����JR�9�vZ#q0�	�Gk�\����"%<�唩���&
�3eFK��v���LM6�\+��Dr���s�ۺ̱�'�&��y�9
w�\��,[5�uQ�3_6�m7�Q���)l��׹J\+�ʃH|�s���r�*'��jk�ڷ|����^~�c�[u����nc{B�]�R{��p;&ޛ{�IX2�\�[N���q�����9xm.���n����.fi{�j�K��o��T���mT�K��:��Us�T/\��dB�B�UBBW`�;ʣک�AW�����|�.�M9�K��ч�,yf��ܙ!�9��t��nt�U��d��}yE����
M[�2��Į��x�T�N�!�a)���|'�ہ�ϸ=h"�r˩�9ZJ�!e]>�sEfJ���Yݔ2~�;(��w�"\�P�F(�wu<Ν��<�Q�zgkV齸U���*γ�M�3�����K�\ə�䤃gT�&�z��B�BX�z���^����3K��l�a���ң(����.ժ�ݼ[�i���N*9q&h��3�K�V.@�\�%������T�j
O.9���-�y��4��H���a��J��3�R\܅|9�_.�Z�h���g\�b`=3\;U�t���H۫��qs��H�	�nН3�J�����EX�T���Jv/�z��<��D6�i��.��=5=� no�lƚ��S����=�sb�z>�w��;A1P�tu#�:��-	��<8�K�C�펝�yoU�7���j�r�����;{Y�X����Y5.��_bg!�\7;F�i`ٔ�H�S�rяn���]��L[XwE@�X�Й4�T�;ĕ�cy9?v`�ǌٜ�h�p�n������V.�ȗp���ۙJo��5='���u�w 龩�昨M�4.�;��\QT�y���M%�<�!�,:�;ٗ�&�2s]��I���
i�\�5Q�{��+�#T2龜�L�J/��r���U'<׊N�����-8�؛!�F�=��9��:`[��[����Z75:��7�M�l*WV��������$�N�^7h�s�_�f*��DO�n|�,��4La��4\�~��ՎN߽w=���mW{�E1n��8%�r+�B��f�,�^�GXh��L��T������6�s��ＦR�]S֪T[W'1�ڛ����l�+'\5p6Z��61�x�v��:�q���n 	���Y��9$�IJ`u_TDꀩj�z[����6���ud�\���/n�)��(9�h?��TII�I[�S_jOu�`�4��qz�f�����WN-V�o�Ѣ�L5Ma��7�)g����7C���~�U����.b�]{9����jV�l�+nW��E�X���k���\�S���ʏݗ<<pR�蛇�{�Mp����=7oxM��Y��7P�QC�ރr�v�܌>����_J�xOOڅ����7

W��E@�;���&t�"�;{���RY�R��,�o�q�P񜨗IX��;��� f�cCܾ��0��-���ֵ�tAm+���'�3e�</����"UͳLю3�:�r��x7�5��Y�}��ri[/��q
���N�����ݺ.���9��2�J4��	�sQ�&���P�����Bo���c��f�c\>���W^��t�v�y�Q�.y^G�$�;��S��7)s�C�X��n���cFs]���E���OfZ�1`�"��n1�~��x����ٺ��{=^N���ϫ�Y���?	[�PK���/k�q���yS�Au�p����{�^�bq�d>���ܪ�vo��<��I����ꮳؖs�7w���}�^��q���2�\%��M���ꌻ7�f�"�v6:K��vv�S���٘�*Y��@�V�B����Ǟh��;ʛW2��G��J��q��U`h:�#���G㖉J=�|��Þ���,�ZA��xr�\d��J0$����h�1r��1=�R�_3}PnM7�?����j,��K����	�\�Z����Kc�b��HWK��D�|��y��m�TU���s���ʯ��.���\��w�\*�0�*#�7�k�gc�T�n�ٽǵ:ޱ燴��履b��`1=(�e�N�	k��<�NoM���3&a�x�Gz�<�k.o�O:�Wˬ��+@����;l�a���O
�ӡZ�#�&_q�8�L�I���cг�OmN7p(%�r��.�TU&�dח�����b�s�K��R�	;�o���3i�����{��Uʓ{bֹ�e��ۂ���b�>����'Ơ��p�����O٘���)��#bK4��9�xt�#f#~�+█Z�G.���ʄ�W��ˀ9=|�P噉ͩ��A�yzѯ�
b:WT@�J}%m�o>��	��/a���j�i�����V����q0�	��v8�ҵ�D��q����[p3��TKDdn؅/^����5LH����ޗy�E��.����9�ۭ���X�X�DW8,,I�Ց|�9H�oc�Fn�P�7�R'�k��t]O�nmG��9Owj]�,���C��y�5,A��r�ðUi�Q��]�$�[���5�k2���!Z� `㆛�m���<}����(�d�gq�x-#�<ݻ8��v�Z5��l5�Ȃfa����u>T���,e���)v��7���yol/3��m��'D�Uz�PT7�G!ԛE쨥Y5q���g2Ligi1C����y0+�~�}��f��:^��T;����2��{���=����
�P��A��[���oh�椷��y�B�}���/�����}���\�[����=�Fm4z�Gd��8��K��ٮ8<f���MK|�H��^��+�M�ԭ���恻 �7x���ub.��+���yI��'�_�Y��8qH�{��P�Q���_�8�����9-���f��l�E����r��n��������̬B��+�<9c��S���XN��_ M��ёz�wsG�}�T%�Q�v�\��m�۶�
�#�q�j�F2�r,/�V�I1��.�w����dP�ј�h%a��Zw�2d��ȝ � ȪY}��;�U��;�I/�qڨ�;�5t
'H��5ȭ�:��O��,.�Z
<�5V6����rXov�,[�5龧}\�Vf���k��E�ي�]��Nɠ�xs[�˓QX>vC�$F���k�#�rf��+9:ޤ��3��L�[��˥���X)�q��8��:+v��^�z��R`��_��«�@�Z�������sWLKa�kEuăp���)��ʽǻ�����v��*�x;׳ݳ��q��Av��x��X&�ӌ��o'A�Wݸ����Z�ͻ�[Πu��v�'%�
���uL�z%	v���;ԈCes�X4Zx�3�]u ���//g��l:F]����^5:�Ѣb��,��Z��-`Or>��ƕ�7�ӧ:�M��w�+(��-��Zh5�DY�:դݦ�l�·u�O�>{I��yx�x��4�`j��!�/�d���_^Y��4�8�}��=�`�j���[;��fE�I��/ =�.�-�Z�<��kf�cyRKX+4��)CEp��Z�����b;A���*�(^�xi�ޏVą{e�w�=�#��iִn{|��o֣eD�:��ކKv���k��~�KɫH��k��F�F��Z=K�uC֨������b�ݔŇJݸ��uY��]�Er��	�|pe����n�R�,.l����N,���K�_r��&��G;(Gŭ��7`tLc=}�Lxy�{F_}��Pd��@<���w;�v�����^AAۻ�r�ݽ&`r� ܬPX��!V�W0_K�:L*PW�Ej�I�#[���I�6��F�5b�\�5ۙ��\�Rb,�cN�cr�\�cj5��sU��*5�"�nkr�,\��c\���.wv*5r�IsX�-���m͝ۦ��5r�lU��9��`ۛ��F�Mwv�j-�IX�N�R[F��'-r-�\��\5���"�h���r�l�������EF�Q }� W�EW�;Ǽ7�Rr鑉����[kU�3��V����κ�`�Ddx«�����9�3-���td˻��A� gqU�9܌��2?�T��L�sLM&�]��:�Cr��Qڽ����-�޸��6��FtY�Z�t��I�է��g;����9Y�����*^Ի<�$�R6:�:���Q<����ɦ��ۅ���9\�m�tn;늇Y}�t�	����m`�u��꒰e��Q�Iڙz.|���ͮ��.���� �h��>�]vn�X̢�C�j+t�l�Ծ�����`���yge��U���{�p�޶���9\�`U{~�8B��|f�:��YՂ�����#�Cx8o����Wn�7����}LwWǶ��_bq��Y5q=]~�Й���)u�����P�_ͷ��΂��v_V���Q��{�WR縀i�G��5�5���)W�KCv�5n1��m=��9���+^	q92��z���DI�;�zC_B��E'��x;*�l��&�eW����A0x����V�s�zd9�w�[�W�zC���h��Q��]-R�;�>��I�o�.��xaD�O�c/��>�U����Q1�|ۊPL*�,�=���L��o*ş^':v}�m�2�+i���[Ƣv�d�)@��.5�u�W��A�$�%�}K�>��u�MeC�|M9+��N�ی�X�T�F�
{��Z+��]�\���]��B�c��	��k����<ְ<�M���8�St��&z[B�d�]E19�\3�ȼ�N�a�OxeG.j�7��v��n&#1��y�|{# 4����|e�]5:�s�� 龩��w�.1�#�1	�
���Г�=�O'Ms�%�.�m��̸��on��ڙ��͸�Pv65��ȝA�x�+"q��{�2��^eN-}ܫZl�K6o#,�^A=�W�"z���6.�K�Zv��Ts�u�L}C1T�Ε�j�o��P�p<�{m�;�=oS��q�7�>��׻Ѻ��̨/�3�������*��i+w�d�p��[O�S<�ȗ���ۇ���g*9���W��g?07�eJ5�Y�}=������4�3�`-\�蔇g�r�ki���I�r&1�䙛�]�ɘ M�2�x�Hh䏺�;�f=>_{W9������cY�i��Z�Z�\�W}7D��Y�5��=vzw'1^�wΆZ�WSn�(��87���5&��r�u�����M����!]}k��*�����γ���&6�mM�I����V2�f��OWӪ�-tlTF>oq�}r��s�^r�����Ś���]u�l�n`U_P�T�Kyq���9�-<]eezھQ�;���G9�Q!,��II�]_*U/*�2��ީ�nݧgzw�.�г�r�s�Վ��$#��M��1�}����TLۅIM�/�x�f�ͨx�TK��PS�oI�b�>Q7�D��P�ws�t9a�����>�Z�niC�yО诞3�.�@(�nX
љ���;���z�rU��W&������q
m�uU��Gi�ʌ�D�.
�.�9@򡠗�Jۜ���u��6�.sP���W׳����缫g&��3'U�^y��P=������W�<�#�y{��kn^tH���N��[���e�^���4qh)d#Y��W'{}����>�մ�Y���-��VZ����aѽZ&��Ɔ�;�N������c�xnl;�"7�!FZ9�B�e˼��9g�*!�q���+�1A1Zi��e�G����椄v�td��JOd���bi7��y�!}[�W�v?���۶��͘[b�V0���tz���j�םY�:��k�5m@�o*���:~�3���Ѧ�w�*���V�w��N�i�9{x�sY�̪�Y�ۧqpK�^V�,̓��.�B;r��Q6��;TN[N��Ж-�1=����x#؞�&�&����I�v:�@|�nr�����k�����|2�D�D�`9���0�ˈ+��f��f"�;(��w��gӪ�p�b��!���:�ע[�W}��(�~��Oܺ|�/1������B��G��zm�lc�e>6Y[�c�v����떞�)�]E<`1�zt��U���_%?D�M��ė����R�yѮ�z��w�q���s]'h/ZY�gl�kۗ�f�T=�5��tU*[(�{�����T7M�:2���%ύ��J�y�Ұ�T�#T&P�1�ђ'�ZX˕�^�c�`J7p���R�Y��*�����v�W%\^㑌]N�7��
��rNk��]?kg�٭�]��݃�$0�T�:C�4/G���0I���i�.Y���@�#��^����i|9ub|C}���?��=H�U��.n�D����[�r��}�c���0s���9���Hjְ_fʛ?7T�[�����o :g�쁠��Jۼ�o6��l�;g%��v���\_s�m�p醅BT��Ԏ��:�sQ������Ge6�/z9��j�չ��p�T�LJj1p�q�ȞCdZ���q�bu�AWK�T�Y��s��歨]V�u5i�5�n������[��S:���k�$3�3�]Q+2����x����9{B�^I���\;�E�q��½��2��1x/��w�՞Al}毽+������W�b���D�K����t�ƺ��a]���3(�T=|�V�|6P���I��]��S�
%�^k�ɝhg�/W_ͭ�kz�.�w��Tz/��k��Vo�թg��.��le�� РӨ�:�A�����޳�Q}=�D+�F1��g��%���`�3iR�K9+,�z,�L�l�����H��g{�n8qBkL!����@"Ǽ�C��gv=��.Mv3�M�ʏ��3��A��Ի9��#g��C�t��� .��Y�wVr��I�P�0�*9�b�7�
�v�ŝGv��
�bo�����k�z��'�q:���=VR��K-���_=
�baY1�"l|9:�7�c+:��h��T�B�� �_I}[T�Z�J����7���6��<�w:Ѻ,��N��\d�?�P��7@�+�����OHjVJ)<��jy(��b�j\��
�c�Λ�aO���*I�	uE�.�O��Onq�r�2VV�y�xM�k�U���e_d9B?��C�c(N�ۂu�_3M�_r����U��嶥�a流�
��V_��+��:`c��;���娃s��rwz��-���o�P������p�as�p�Ń��ڿ�ii�4�GK
��9���5���7�5�0���0S�֩ܧb���!�?�Aܗ��<�j/�o<vک�X�L�s���Ed:u��jGy�!��'{]�z�3��X���_=��:�.m/F�/ج�g0n�lz�O0����7�X4�W<D�	��;�=v�X�G{Tt�޻rJ`ȡ�	�,���J�<�v�=�Awe1�/�w8%��M�N΢�U���E���lx̫�Es�'<׊s�/چ����΀�K=U'��+}�_����;�?	[�[�s�&s�	�	�E��R=���ܮwe��$��}G����v��O�����8��O���hD#�=%hˎ��e���63�z�Ӭ���p��x]�����$���f�)^q�d([���HqԇJ�z�a���W��7l�ĭ����9�''�.�E���	_�e�ب���|�>������Oy�x����\�{���q��@�!��%���o v]뮧Z'�(���r1kI.���ڜ�
	hh|�$�ﮊ������ع�tJP��]�{k�Z�,w���O�AJ�z`�#�'4���˅uo��g�c�ZԾ���e�<k��q���t�HY�}�XZ(3˵U	�`Q%.��53y��R��=�Q��ju��4U��Xx�#nL�Ⳳ��ajW��]=��
,��;]�N��^}% �MfД8숾�؍�7���i��Kb�nŕ�9L:h7h�7�Y�K,�F4j98�� 4���p�]K 8�W��w�-}�[Jýz�`�x�,���N�q��z.U,!;�24�vV���b�{ɥq��CL�V���J�]��]qi��T4+\�Jܚ��P�����cݼƋ�XU��Ç�(��0�1�Q�*Bc��	����&��Ojē�E}���yMd�b�g��r���T�<LM6�]�3���; Z��D�a�0�hvu\���
u�I�{�ok]b��u�p�ځ���?#�O�]�;��u�ĳ6v�|;����K쯧���������/;�N9�}G��U+�{
��֍��8�R�w��X��3:�&���^�����ڙz/䷶Ug;��!��^AxK7Y]�F˽o��!r���!1�1GbCb:_6;o�7��:�;O)m�aeʶ�o\5�Q�gj)�ʂ��g�'T5c\%���3�G���:�:XJh����a�##P��
�㉠�9�Lh�u��Vo�4�z�w�[��@�0���vU����ֶq/.��<*o�߬��/�u���v��B�0Yu�]]"�iX9ڲž[��@�d��i�T���Cmq<t�����na�]�8�]�Vp����ա���l��K��x�3��V��y�:�K�n�sWf9�<�+X���F�'��KCc��yi��-=�S�_.����R��]s�}Yp�����7މ-�uQ]=2�x��Y=jOn�v(*Jtj�-��^_K�e,���DϮ:��R٨R�_����q��ؙ���k����y�Z:ïy,���?�Y%���Ϯ9wb|C}����VP���,�YyȂ�q����f��;�����2�?mN���h9����ۇ�r�[{��q�,l6�(�f���φ��O��V�;�C��m�f�	F󬝷��2�9�)�@vôn&!Ҏ��󎯘�7u=���8�.�4jz\}-d�vlw0�Ꚏi��MƻG#]q�n��/�9�=p^o$�W)%^�a���q��^j��I'2�ӆjp6��n�'��A�s������c�����}�`9<$�eN�t)%~Oxi�0�f�ı�5p���sh0z;jsbpѢV�v���Q�x\і[�/�7�']�nb�*�ʅ>�����w�ǝ�;��ﬥ���Ka�q��V���-��/Hn��uq�G��
�kyA)�_�Ϯs�Ny�k���s���Õڪ�3*cF���)(pv�/}�m����Sz��S���ss��):}0��1t�N�]���Y�:��U��3(���W�s�y��T��D��M;��T���V�&O6D�\���ޯ���G1�E\��uܖ�)��"f�8�8ڐ��zF8�-���6-�{q
�u�W�s���ھ;�^m�q��9j�����-WӮ�=VR��KoTK�Vu깻�
�B�';4��	3�M8��]Τ�TmS��J�ݷ���/�Xm�4���	02��]b���t�>D%��Od��w%�A�sWB�c�����G1�P��Rt��,%��Q�&(%���.���}s$;ņ�qv(iH<�r�V�p�܄�6��9R�������>���8]VV,Y��o���{3��t×�D��2������'*��%< �S+�E8����j�{��}/����Kȅ��`�j�Ӈ�aH�� ��^5�ַ
S/����6B�v�o�H28Nw�E�3731_��u9A��J=5a��1Æl�V1?O���"��r�`���z��rK�+6��u�ʴ3b"7�sM����O׸wD�Ճ�-Fb�4@j�Jf��q�[�b�Y�y-&�&����P��7xh��|�ZLxs�͈�Y�h��f�:��bʙS"bc.�AL&������;a�{ٺg.���<�\�h�Y�TjNނx���6���^�9#�B��{�%|���Xq��^݂ۺ��<�qj�6(Z�E�qw�kX"TB/G�o��	�@�o�(��w�P6�6��9Ҳ^��m����r�{��A�;�ye����U��O��5},|]j���;Nܙo�ج�4��'8�V�:�g$���{w��o�SU�����l�m�g\�/�M
	�c�#�}�jYS��tI�v�^u =�����kq��+P[rt����S��˙B)�(����t�N�̫Ն������B���ڮ�ݚxʽ�_������n�ͷ����Lf����aŽ�F��<�hj�mj�Ͼ��F��uv!xw�8ll ��OE�͵je뽫v%.��Zvb�����X�syS�i� g�	�ni��Y5p8�������C.SF�/�31�t���#%u��$��=&D��t�O���`!�0��-dS�j�r�f�i�G/g"�pP��\|t����J>�7��܎����n5��|1�ה�O	��O��
k��ܙʺ�'jX�����Tl��Q=��ЪN�9���@���ws}Q�:�ۛ��z�OE `
k��ס�+kr�ǁ��rS�����#n�=���P=�e��R��,d�7����m�C��;������F��{,�C�-.���p>#Wb�nm���E�=��6�؜@��-����Qa}8ىq�C!]8�3�d�����#�p��� ��uEZ��38ܵ�x�ڜ�p�(Ӽ%�Xb��MF��B��/�zՒ'r��pk��4޲���t�7.em�0]��/9�
�`2%��2Q�@6���@b�B�/)!o��S�"�^�r�*+6�췁�Jn�V�CoE��굹[;�_�gn�n�o��=���yV�+[;}��l�+7��Y�{���ӻT��yL�6Ӂuᚹ�`���b� �Ct��Lv-�]��ab��-��k��1��%���:�1;�_8_)R�j��Gaƻ ���,�۵�:��յ�3׉��}��<'%�C���Ã��]�KQ+�RN]��/i�+���q����6�fd��ޗUh�G�U �%d��Ŏcnj���N���)ܖJ���k�"�np��wv�Uʹ��Qr�wcr������N[�h�;�b5t��*+��˻����71��]ݮ�k�4X�7*6湪7]�kE��W�r�X�ۖ����\��®U'9����9[���\�wrᨂ�W6�G9�[�(��p�mͮj����+�Es\�.b��W6�-�����F�k���n[�w;����X�U˗���\�b>��������c�ȳ�)�OX��i0��FK�l�M�Ɲ���+��v�ư9Y�{����,������YPyPs����Jޥغ�|����ZW浟�f˖R!O�!t۶}l��.�\z��{��Q��ҿu��T-�˚��v�����"�͛|7�0ě�o'm��P1`{f?Y鶔���T�L5�.1�0R`\�GWTgmx�ǵ�z�i�a�m����+ȼ[���=<;u
���[��;4w#W���Y����Bxb�7��z��,Z�#�m\���Y1WF�˛V�ܾ��ŊҞ8Ὢ��5�����ۻ</���j�5gX��3�5��׵��S/-'�C�=P����c2��r�E�VN��v����ҧk�-���q���3͌�z�Ӭ�}��G��ʡ����5=t:Xr�s�*�k4o$�p:"��C��/S?E�"e��ߣ��5�9�ʺ<���~Qg�uBWe���}���&jy�܌\x1�y 	r�z�3�e5�����^�V��˦'�+m�Ϊ̍!x��Jʕ�렱�{r����5����*����fLG������=����G����{hypi�J����Om�L��cה�QugTÎ���rVs�<��P\w�R�5`�}N�o�k���Wк��V����"dꀫ媕X��ډtb���c����{��\co�Z{p�9D��@Т�>URr��ll�!�篳V<�|jN?�*������kn���gD9��B_gqQ"3&d����]Nr�Z+�&C�_>�ܾ�����5��5�7��+�AK�2��0P���4�Q�N8�3X��>�����-�p��OtS�pGbQc��v!v�_�ΰ�G�����_��g;<��D�q��Ҹe�v3>0ν�1�ħ�QA�{H�Ћ=_�|4��Jܝ�k`G���gmc_Qz�}㒖��	�j$%�T?�!1��N6��ɯ��L��(#dPيǸw��ֵb��M,LKn1�3����:-n|��hy��1�N,�]:�ʷ��ʷ^v��$�18fځ�ܭxn���ޓs������OZ\�m��ye��(�j3�`�
K��6u*�$����iΦVZ����rTp�Җ���+�uh��F�e�:���+J�����<�i�̙� 5����*�u���82��;�7*�N��v����[�:\��N�yf����n��k���������v瞍�N�i��/o�i��yr���'�wC�<A-C8OJ�O?������Ǔoj�qڢr�4K��j�\�������ŭa)'kf��uvn�9����>U6��=�}[;F�6��^�h�K���,�j�88�{�m��k:���S�U��Y���ٱ|*��*���쌡���{�M��uٷ�TgY��7"9Um�	]�S����b�=J�Ӊ}��]+�ثp�Zm�i�|�:�u�:�˺�F�Z�d�9B��uD���=Q��4�{���-��OmN7j�p�^�x�i=]�����`/H#�Gp�.��ԭ�R�_��Z���f��V>T��_��jޡs
����}���%��s뿇.��������λ0��R�����.&�r'�*3���D)��]0%-����+�_�\rs�Np�F�`j**Ob7̸=��<[㏏��@Z��r��t�+.��_RF���/Ǽ�<��˻���b_����O�5?6�v��|����A���
8����g:���ⅽ�R�!h��=��L ���דIu�wJ��lwF씻lk��n������.٨�B��WP�`��Nj9c����Ef4�wej܅���Is4��������j별�.�𰎹:2�z5�Y�J-��/�瓜��Ꚏi��Mƻ�r']�f�1?V�9;N�"��K��^\3���n�Ȗ���m'�:U���E��6�j�ǌִ�2%�a�_yr"�~���Q�~K.s�T�V��l���̱�W1��:2�{MsܾY���9�{�����������H���GjgFr6;����a�m^m��s|�G:��~Wf�X̢�C�Ss�g����c0MSu��.7�:1C����)�l*�>�^�95����Q�׌��[Mc�qv9ۓn'�*$�}p1GV�>l'M��ۆ�W��uE�ܩ��u���o��~���4{Zή�1k�{��J�����yd�\��ɷF7�v^\�7ї۠oa�*���̒28�3k�VZ��i?�f�`�*�q�&�22��y�=8ʛn=�8��<K9��ܞ������灠��[Ξ1��U���v# ������W�u`��NtK�:��1��۽O�A��L�k�s�~�g�1Q� w�;���]9��=�s�TÔ�;vʦka[�v�9�W��t����muP�lÎ,���D�q�3�[;ս�	c��[_<㔝7p,)_oL��.�ˬE����ӽ�r�j��IM|S�ڜ^tC�r��4�S�o�����i���}a�;=<�y]�>�[ݶ��a浐`m�ؗL�ȅDz�V��\���	F���8�Խyp9��o�� �a�
ٸQ��9R�us�,�6]�r��P6��/\�һ'9>\������t���CT�ġ;���C�E'i��G����

�Ga��53W-�'٪�>^oE`�mڛ�u^���t}�����|��㽕 �t������$\S�F�K���>���bK�*��'u�f��ʼnn[)r��]���&����vXC�3||r|��Vܶ`���lW�sZ��޵P�՛C
�`�x-%.�ߙ�կV�+wP�:�H,�(g:P̊�vf5��×�=�B��<)'xf,��9�F��,ʹ!+�K�&M^pe���v�`Rw�\3��O�R^��q�6%��<��#��嫥R�����W�;��T���id첮0U��Ɏ���-+����$\#㳳�,@���(~�-�G���t#��I�E��1D[�Ҁ����{����#��ἠ�Z�X�W�;NK
�U��4�	�Xr!���h�PlI�.�pm0*�`��W;`���3����V��oD�_Aq8�U�C�W3Ƈ��_����C���H��΀oU�����#����y��I�����z#�L5��Cñ��\�$�+�0�(ϑ����,���.��ǲ�c�b�e���x�X�S_C���K%��=����l�$��L�$yT<�N+0����-������iN��.���_��o7~��O����Y��}���`65�*�륜E�wjs�m�g=��=6x���'��R���BS�o^�j{F �/U�h�*g�ue�MT��L��2�������2�}�/�W��,+�޴8d�t��U��-��� ��0"3z�L6Už��nf�}gն�'�,�ȈT'���W����_nPݾXF�o��?|��VU/;q?�6Z��3���ET*iG�7?M�;�~���
�|пeV@Ӫ�\�7R�^�[ͦx�W;�Kn��x67��-ԅ����vN�3L	e��m�!BeB���pv<�P��֥H��c��ǎT�h�L��c���%�li>��W~�\MD9�L���Ă�}EDQ|v�;��`Czj�e��+��ȅm�M]��Wn��V�%�E����P�`�4��¢��M9h�6�V���䲘��y��n��B]�}��.�$�m�HP�kx�q��4�SG%��so�^�X�����ҟP~��΋��]~��O��x�ܦt5�hP:�s��JnD�b(3)�7��U�5�4���\��|�b�|S�'���?���x/O��C�P^��Ubz�j�ک�U[ȋl��_��b$+�ڋ<]���H<m��nO;��[)�S���vct�Wa���<ʌ�^�Z-���&]e�k���(��(�Ƕ�9g��w�6V��B���Q�}�E�lW.8�^]s�-{%��1@�F�b��&V��$��MѪ���5�ak?p^�>��uF��٥K$6����j���81�r }������ڶ��36�4�x�f�K��D�b2�XN&�t�nP��b�Yf|��g�|#+#�7�,?�X�;:v�\aVv�]�Me��k�qԼ���~zݦ<�]]�,��Ԯ<��{� V���'1�|�̛����#UΉ/w�e�Ы�s��yL�]��]�]�fJ|�%
۵+�"8��Z�<o�͊e�qy���iܵyo�e� �>>�:�eV��\y����ؙ{�XG�K��j��3���#�+2�y���f/�.J<8���	��}-��Yu�N�P�Oף>^��+W�9�>�ͿX����Ŝ�o�	�~w�d��PȁʌÁ0[�$������q'(7-��^���p��(�L��h
壾���q7��H�]�7�.j 55�D�u����>�<�ު1��6�n�*��gu�5P[z�|��{�yD^���q�)�y�i����F���V<�YV4����lN����^��#�p)L��*5�^���ȟ����&�f�#���췝�'n�z꼲K@9	���N}�ycѶ�����u>d�d��j� ��	�<54h4zszlM(���6Ց /P@Yz��`�54-����u�7��Lu�w���UAc�L�ލrD�u�{"��R�v� ׹��=�����d���a]z�Mҗ��a+��y�r��xN����6��&6qc��U!f��m~��~y�j%���t�[���-b:���Ύ�檈gڦ�7l���G���YB�5ts����1�5��WF�p��S�7�X`;BIخ�e�J1�x��]+�%��O��u�����v�@\��IP�=�6��9t�
>�E����S����Ó���׬����C���5��r��� ��
|�9���NY�t�z�<��ܼ7�3�0�̲�[�*O��1@���D.��xnMO{�5G^�l�+���9�V��T������R�כ����"�u@�v��Wuq`F+����bV��PRT�\����W�߁���x�a!z�;-�^Jo�a��ִ�S����rO�'��d��*g��9��頯��p�ϣޯx�c/��"f,�����25��3�]j1p�����Ol��FU1u2����<ybq��B�/�"�W��`�����Ed=g�� �߭�q�u��ȁrY�x��Á?*�te����px�#۞�{��r@�w[;P�����IC��Y�ƫڑ��~�p�P��jK����s
;%��<gu�/%-5q��)�V���tS��P�2U���b����҂8�q�D���\�������H�y�3>
Z/���z�0=�^e�N������P�	תr��k�,�R�y�O'ś�Fg�Q?)���w )�w���	��c ��ώDN2_,�r�{��{�f��͒���)��(���n�A���A�`�-ᅯ|{I":�w5��$}���mYt�@T��#�����ٕ8I�/�We��/�%�Y�˷$�0�x���s"�	��]3��d#����q�b�+�P���14S�i�j#���̦�O����~�O�F@���2L2CTvD���9�����q�|�uAU����Ŕΐ�@��q/��1������R��d>6�Qb���Q���U�v�g��9�t�G^�uEk�k�2D�Eߌ�)ߏ���ʐk�����auz�J�[���<	��kt9Eo��B�-Y7-���pSv"�'�1+���'�!8�XT'��oyT%'i��_>�+W���s�V�����d첦n0U��\��~[2Ѳ���,�p����6M�+1�~R�*��Mϥ���@��a��`W۞y����z����cx	8ሪy_�Ztz?:�צ.�g�B'3�yB"��Mi��.������"�s�xi�]���Oe8�/��:�3O���B�Օ<nωJ��<5�w�n���Ét�
@�`��[��o�ن�:��N{c�LydW�s��|�T���$�)�4�C��s������OS<�N���pL�:e���b��:
�֥�د:��u��ρ�[<	=�2�Q71�_�('����ܤ�>��L�mG�51�];􃶵�3#ܖ�w�kI��̧��4N,*���Mkt49����<�WK)c��m^���=,i����\�ͬꍼ�+����J�p�.��r�d;�E�Q�˄]b�љid�9�ͫ����r>t4�m�r3�ȕBj2����ۨI��/o��Jn.���i
c3��	=7P�ק���G:���&�g"�7|�UՓ
}f�4�铆na�A9#%�S�$@�"��{�m���������yؠY94w�a��L�%<0c�8HFx�/4�����+�6F��k��
{,ު��Y1��e^���#�����ÔUL�,�g-���T�T�-�V�`�5"��W���6nA�擗�_���r����Z�jަGĠb������Vg[����JІ(��i|l�靺�����sl��������G7+�T�#}H��'.шA5it����-ͻ2����R5ma�[�9vE�(�n��㷻�Jd�Ox9S��=�x��E���]�*!n��Ys�թi+�n5>�f%����{��e��ؚ��|��fʏ�������������N�H4m��g9´���n�^沐�f����-��^��I�V�%c::�Я��D\A��m�W�;];�"��)����^���V�w�*�
��wV����}��/�܄�(���g��0��Qښ'fG�:�ag^>����>�l�w+o@,�����v{A!�g���w�
<Z�87L�V��
a�y�Y��и�_7��1zwQ���Rfe�P�z�{�b�s�+2L��^�M%����z��ψ��ŉa��+�;]���k��[�α�wI�8�U�y�F%���v�y���Gd�5:�|�p^Y�M)\N���/u�f��t�f�:�;Oc�Ń�G�d�K2t��qs�y2;��熹��w�v�>TR<B����	��=@˳���`����\���i]Cz�i�솂�jvd�`�C��n�#Y+��q����=4����%|��&�qTڰ�'��ukD��6�9�&�����?���ya@��e��);=�ʯ&��G��f�O�b^Sr��jK�R�3N*`c�a1tu���u�6vX=*��Oo	����N㹆�]��\�0V�C�m}��=}�����Ղ�����Zk]sC����4+&�C��;;+~+~A;ےh�{|�i�k�岗�f�Tr��Ǿb��X2�U��k�0����Ḥ\2-Q�E�=��l��q3�hM2�Ύn����ogK�-�9bNz�f�j(�Uh�S1��R�xw�`����-�������y��A�s=e��g��>�̲�9��)}��r��*����$��E�F����+�b�W9���h��6#$l�U��]7)-�ݍ\�N�;��ܰX��k����+���E�r��ܹ��[�ͮWwP�:h���+�gv�W74k�Yݮ�sj"�ЮX�\���
������)��QsT����� �!#RY�\)+�9k��(�K��l�,h���n�4nn�s��4����K�7+�sd���k�swZKt�9\�v�gw+�4���s%n�ܱp���Ӏ����_t�6��3Dn�[cq�̮��f-���NWRv��Y��M�Q޷���P�f�y+=�}�_�=�ژU7p��X��_��3�G����\ϳ�V�!�9d-Ke�)�AS8��1���o#��ʌӰ�����|�����~9�z�HUϽhk֫S�/=��V������ɚ�.��%��Ȣt����=`��E��)̀��o�hp�����}�~��
��g_���x��������N�U�d�H�P�&&%z���Q|}��U��h���gt	��ѯ �@�����Y/�x���;ϕ)h-�
#e�C�	�����mMmot�VZ��y��q�"�e����^U�+��R���<���*��c��"#���Nb��ި/��b��ښ��\�E�>܍����Ժd���5$]�Sp%�[!\@>�nS�ҹ��Y���,����9L�)Ա�b�|o�S�f�-�7-���3���1P%�G3�H��m�9a\�����
���p(+��vǥe�e���d&*s<?m)��}P�[[���P�b+�d���d��iu`��̩á�&�N�u��7�h;�.� ���W�<��F1��/2�P�c�[���/_q I���"B��zg���=E�0@ԈZ��zGM����
�]vL��xS�b)e��r9X�]lʙ�n�V��"GVUh��m�+�E��D8�s�
 �m��l�.�]�l$�P�d�};��y�z��o�?��q��������e�B�ܼN`5�n��u��2�Oġ�!����m�u뮝�y��v%e�GR�eűLܸ���:�{%�(m�/=0���S��^}�c����g�ᐙ�Z�(	���\�d��*���{q��9'���I�z���*֟g ����Q����ϲbCI�\(��e��)ĵ"�+�C!in�X.���x`go�CL�L��גAug���h�IR���J7
�X����p�G����Gr�Y�/#2.o�Ʋ�@q<�[��Fs�w�'ƙ�J���&H�G�ڜ��Q>�o8Pr�X.T=��6�.Y��[�5���|5r"�OY׋	Yk<��`@�� 7<NA+�f@U�yZs:Bmm�ƈ]W%4(��OAQZ2����7�T����nd��D ����D�u�Ip��l��їL�e�lW6���H�'ݚ�{��
Q�!aa��ۼ�4�OD�}�;EdN�<�vKe�6�;( ��|u̱�B��!!=��[�e@����T��ӹ��*�L*����H���f����ńQ!�$I[uty}�X@�������u�F��J�9�{)}�\�ɧ�7ך�9�����}�q�E��x�� P���w��5�n�٭u�33]>\�z�^_6��ް(q�ZÚ;�����moX/�/�Q~��vJ�5ш�6���=�[u�Y-�!�ڹH"Y�Bg���e5�xj�gX�:o��f��l��a3(+��/�5��z�����s놮�1�߮�Ll��x)3G�x9n�l烙���P��E���ԃ�ĭ0��m�b�ؓ�����t�w!�P�p�ʢ�0蹕oY�ZEЊP\P��ٕ#/�N�@86wj�ey�6*��]6v�h�2n<�W�XM��Yҟx��
�)�t^�,5eN?H����X����֥1��4���V��L�oI��|$��L��K ���8�.It�m3.��>kQ�&�2/f��o�s�J4y`-�1�E���[.9�e�t�ͨ�	�2�����l�~�`Y�V���>��A�]�>��nȄ�@�.�|��s���4<�O����G�=���/��c0Ժ��c��-G
L�}���a��g��Ğ��0�k�*���H�0��7WT�u��֎n�Y�S�p	j����/"ֺ�hH]z�w�H��6t<�\�i�$��0�)��e���V�����Q��}F,t.��2�=Ɂ4���QvI���¨�t���G�����)*+�/�Y�<�f�u��W�!R�e�0[�a�ɓ^��t��Ǚ�3B[{ʤ��"Ů��rw��{�i<����ɘ��7{��[�=��l�ͪ۬ɭ��XӺX��*�6�G��{����ڪF�?]�{ %�C�)!�o$�T�[������� }�9å��˭�+e��BS�((�7 �-R0�3�%�!�	I �X,����#=ǥ�Ct���0l�d-�5��ɂ����(�$Z*�޽qc�j<���[#��,��̞5RBW���)��qN{�s���TFt&���>��B)��<����iqb�+2ʂqGɰ��g:N��#��%]�P[f��~g)��j��Ly�DxO�y���^�oES��WH�l�(L�'{U���[�L8;q�$*,Z;ئ#P�|Thֽ~c'e�lྭ��En��L�"z�w�>��>ϡ����ېk�>%@����g-ڵ�r��1���D]iu�#G`�	�v	jɹm�o)���JO<bW%���T�Bq�f�(ҏm��[&M�Jܦ~�~�E=϶J�0SfG!5��ʸ�V�&:�-%��V5�Qև�R��5���#Bj\\�B}/qo��b���1�(],���.����z��{��m:.D
�Z�E�4���ޞ�$�.퉼�\2��\fذfd���F���Q�Զ`�~�|��<����-�Q��86l��M�oރ=���<��ӓ��yYI>dg���M�,�5��o7�-�D��a�/�oGg��X�Z�u��mX6�=p��X��S�d^]��Z6�<�c���i3-�A��X�>'v����O�b�kM�K�<�m0*6�y��o)Φ��{I#�e�-g�f�\�{޺Cx���H^���q|JWaᯌ�C��U#u΀o�\�܏f�A;����9�ã�=���Ol{)�,������m�du$�!x�����DO]Ukw!��u�a��$F�g��v:�CmC���֥�آ���n7:��Az�'��}�ԖLM՜����z��S詗�c!eԳn�X����s�O���%�Y�p��o�ڮ��Hۊ�^U���N��F�{�<"����j����(R�}�CFB���=�0�uK�B��q3��i�߫���`�(҂*2�[�"�^S��R·޴8g��;b�%L��;���܇�"��$�`֥�ĕ>��fK(h�&
����@U�xT��h5�k��5B;��s�p�ݫ��=��2N����u(�_D(�g� q��˺|�='P�̞��;�U�¼�[�o昨���M���@�=> g�3X|��.�O%��������Mb��c�^�V�����4�boW$�h��N����Q��l�.�7�{��zs}*.�{%�M\;�5��sE�L�h�r�@�C�#Ǳr�Zs�_f���=�Ӵ_s�z��oӳO5C��`��̝Ge����c�BGF��-�@9��v0"�8�1�Y{�j�d�F�\j �d�w�\	{�� o2��%��aQ{�wu
�&�0��B{����*V�[�����ۇ�߮��o&*Ҏg�+Kƭ�b��w�kO�H��!`@i��2ָ���b�7� ��<같t��\���q�3�ѣ�toDq�箋L���Jɷ��uQ��8�a���w��7�h;��� s�z�]�龘*hF�>cGY�X���&�V��P^�k-ïs1:N�hZ[��,&�z�6Nz��ef�:���J�������:�Pֲ5�q��e�:�ױP2|�6��xm�qAz�%�F�B�|�{���R��tK�g\(d&~��'Tj-�K$6���j��ب�=�qoԩ�����ڒ�ۖI�DΎ�x{*e���t����Bp��t��(Hm���2X�Lu�	Ri�/�T�aP��g 8�ȱT�C�����q����;Џ=�򦎝c��<�F��x�C�+[,�=5�1�%���$���`�Ž����O�z���%����ڭ��j/oF���qZ��e��:�sw��@����`���/^��I3�����]�iy�#8x�<��v�(�d�s�;��#+�3Y3p���"_דy������[�u�sr�����juB�7]q�57NC'�o��S=j��}͕;��ɾ�Y�RkH���μXH�B��� r�0�LAn��%x��k=ώ_�=[�Y�ʏ���wr������g(��5�Z0�%L���� t���MI޲��_S��2��=ٔ�������<��&<�|�G_���9��>����K$���B8 9ލs=8OP���ϰu�r�$L�^'�pdq~-�گI_?O�>#��O�3X��\]d�VN�	���*4^��w_�M9��y*6����'u�-$��\�� �9����W��W3ίh-lr:� t 0��7d��Pb��soF�����5Ua���Df�鱦�}]�"w�����]{ۨ�DO(N�'U[��+0�BT�}	�0���n����>B��[&HG�>�v��|��V���瞙"V
k�G��g�Þ�~�p�*F\l�v���l��3�2���CU�Zj��>�&3 �^܎C,�O�IXw��/ڤ��e�X�"`N�\��Н�4W1�jmM����u,h�jE0��rիe��Y*)ϙY���|����E������f�M������F[��<�A�E��J��Į��+)a��{�yf�ZU��[5(կ_�i[�}���V�V�Է��Xn���q}�4ئ��EӺp.RU��#�sj{��A[4,=Re�8]b�gw�ɝ��S������8O�,%��5�pJ���د�w�����[Q��RRo��BM2Q�M�l��xش�S^���{�<n"�%+�,e<X���3�C-�y���DȚSU�^�/�:I�9�9)H��ԇ� ��b᭩f��Fa��T��T�F���������<�����S�����So^�hH]y�w��[��i�.K5�%Q�p$�Ts�ܕB�L��M���U�eX�.��S�,�t��2��*�j�]K~��b������ r��Ϟ�\V�՝�2��;�tc�� �զ_�S���S�	Clk{�=��ja�w��߯��g�Wӝ�]J�H,��0� +�p7 �3 )h�R��^��g����w���6>�����_�޻#?�N_��<���R!V�G�DZ;�\��i���f�2V�l1�������F��(�H���,���'��F@�v�%����^��b��z���kuS���K��z��7�2Q�f�c����u�}�|y����� �B�OT!�쨩}[�HqO�2�ns�em�;[����{��
���h�1'��f95B_1�����,D:���KM�6�X�]�G�!���f�M�Ne'��{(�9����4�F��Ļ
V�zWr�g#��>��>Y�e���y���/�Jj��x!�u�q����Aٯ}<f~����;SU�t�	�]��R��*��q{%@���'8t��=��皃6���(���E��v	����oo)�؋�"iI猤���B����"�v�NM�;X�U8!�ǥ縷���d��0r�Y;,��a�˓C�l�F��Q3K[
(
2�o��L+�����4�3���㳷2Ǫ·u9GD�?��]L
��:d�uRq;1+�ۤa1�����}�GEu�z��zZ�X�ۆ駅�����qR�,�����yk����Hu_3�fJ����qeCi�I׼ܬ���F�찆�F�(����T���K7��t�*�`7��@�zȿ�ҽ��e1�W�s��5�#�"� B�Y�2,WbE圾i�"9�f�a3�'��[��"�SZ�A]Z�INEyׇc��d��������ʞ�z���&�2���*�\T���d,��]9.s���`!�)�@�Ke�7��+�ճ�n�Y�9f;f�P<}�@�Pg�HR����r�Z�~9�z�HUϽhh^�S�?^{�W��t��/�~kh�W7�E�^,�xGN||�T�>^��S��풥�>���m�tULvH�aҺ�kov�n��i��Kѭ[�����Q�,�\~���6�.�X"^��Ŗ�7�/8��]h�.,�5��˽�^�(���/R��s��;�{��#���x�}����ߌ<%�P@��[�"���9�K
�}�C�t����b�C�ӽ�0�+téO>%`j�-!Z-�,�" 5P'���=G>�/��<8ķ���d��	�%L&�M���[yt������@K$�;ʥ-��5�?p|�K����<�f6v���1���⡦*:�5~�oޤ���y���`қs<*�;�.���q��{"�=�� ���f�s,cP�'ױ�%�VK*K�H����w�M����{ʢ�=B�u&%do+=�2l�9>��O�����)��Jy���'�n[�����k��A;�d_��!�Ed��q;~P{�������U�Ɇ�mhwS�:."��'��:����O1υ�6qF:�u��̦��|�Դ�Ƭ4��f"FX�.�6��v���Y��n-�v�VC�p�7�q�2�ջ�i���D����G[6�/�)nyk�0�>�@]�n�B��=h��7����9��m����>��l��{)������R���űIq������ْ����UJ�?Wᐇ���Ľ?h�7�"�VulWR��M�U� ���=X�k-�J�c9?r�9&hS{��{�.ާH�[k��1a���a�0�ְ�u��ڮ��oYu/W:%�)�B�ݔ�r�r�B���
���V!�q�Ȁ,nz��f"y��6�Bؕ�7zw�Y�Ӯ{�[��`�V���Y�]p�4jb,��N�����D�<@���C����砭�m�Mn1�ժ�z����	ՠ�f'`iI�l� K�Q�N�s����|gj�eX3p�7�PS|��e�lm9!���+��\~����H��
\�>;ǘ��f`M���m��C��H��b^��Y��R5m�l6d�Y̽����1͸���f�C�s���+�%}�Kw�>��/{�z5��Iv��]��5�ٙfAW`35뮁�}O�zu����g.�)��D0�3��k,�1j��D�LW���=z>��x��,|+K-�r|s`�֓77�n:��W*Od8�X���\�k@������x�u����=��+L�`c;�������&���-�����Վz�Z3d��B��
��H�n<��s	�+%	�X֎��Wf���WH��pg�*��gb�{����Jy�IF��t�Y ݇Z]���%����i�Ѻh��r�Ϗ7�L|��r'g�¯vb^��ww�+3�[�þ�.fU�39F��gQ�6ݨP�_����,�f��yDB"Σ����B���I��c{+�+���Ѷ��/*��3I�-���A�kROZ7�bsg\�����PK��^�gw���[�y0ǀ+W��@�\�Zs�q(���)Iv;��	����۹ㆣ�7��vPp�䁋8s���b����j�f�O�AA?�SԜ��ѓSx���h����4[=,�#K����<���Fx.��6�}���\�nu�(d�Ͳ/�#j���.Z\�Y幮>�[)����.g�b&��nn%{[��J���Y����g^��>R.["Q��*�ٝ˛�';��v"Hս��sq\�L��gM�>���w����0��7�lq�η�j�e�A�oi�Z��{�s}:9U�L�/zPG[��fM#x=b�Kܤ��߲����#�b���^��Ġk��&����oT��77�]�^��|��`�<�L��8�{9��-�q��t��Y�άok�-����=�W��~x��+�N�n�����f��"�T��.d�KRNЕ��C��X���mqk�]r	�[�IyI�%��s�x�J�O��8�=���*���-Ӫ��H�&�I�NވZG���Ւ�VfE�]��υ5)�O����=�.u.N��X��LH��,��]���]���F�O-�w�����ܼ�I M������俬v��]v�I�1(t�qg��:k�fU�K���o#�*���q���0�g<�&��9B�T&w�}�r��^�EkY�{��j4�_Q'�$}@}@
=W�͗w-����˭I4��Bd�b���;\��把)6�c H�ݱEr�g;��ƹp�&�@�g;��
19vɡ��g]nI�b�rwpػ�5����(�#BIQ.t��F��E���L�$w)%�u��Ewq��븇we�,фw[�HQˮ�&M�;��.n4�wZ�n"�-��k��3��g8M;��]�d��(s�!B#���sq��vLA��l�� P �u��Eר"���K�U%�vi	��ԯ�[��4�J��V�I�:gnڢ�EΦp��#7��"�k.�j�����L���d0�S�Fx��p����a��+�U,���̦�uϚ��5����i4�n�
 S�i�$��	����)��+��������N5��t�nP�ޞz��țiڙdXp�/}����o�V�񸾒W�X�>E�*P���9Ϟ:�W����������Kqu��m�s�mDh��r�e��w�=��L�%TA��)* �[S�^�`������-$D)�3��M�.]QޛzK
ᶴ�*μX��K*�<�@�v|������p
���:@ajn��\���؉ͥ<.S?�&�l�Kz�צ
������W��#n�v�ۙ.iSw�.�=��i�T)��zuR�e��
�o���9������z�O������tiE��݈��q��G�����F}+ԅ\EK�rK�|�E�vʁ-���3�U�N�-���f�4l�.���E��a�K�1ш�*6���=�[u�|�̐�xKD\F�c+C��x��@���ϊ��>�T ~-���)L��soLo��5xX�f�`͕�4.��2�#����eܷ[^�V��Άc\��\�/�Fg�v��1�^u����n��Aׁ;c.뛜9�1u�_fZ���ǮM�_/k�i�pH���Lf�����J�n��z��p���j����0e<_����wx���C�o)om���n���k�/,�F%���2uU����pr^��%�.�l�F�e��u�u=�tvT徝7Eo��S��)��U�.�M#/ё^nXe嶨���e���Ӑ�ԣ�.�iY�w�ʛ��ڊ;�A�`X��e��z�V�	�lv�,6Ye�<��*�+/�^��7��7���pF(��|6-���6�F
�g,ի��7:��Lg�%�ۨU��#h������ay�UDsϳ�Xۙ��<����.G�������/R��4=��_,����<�NgX�
�G
㥮�2�{11� 7dG=�����7΃/>4<�]J��J�hg>kF'�{±æ�dy�)�(묮��a��g��'��?T��2��f���Lr�I~�����)����,C���ף7�>�܈�P�#޶=��J@�,�ĝ���h�Q`��M��l͘�W:�w`G6�"��iٖ8�9ҬV�uѕ�?`�za�}�e:�q@v���d����N�޹�*�s�>7���+�^*��V�;	N�t%���c%����}=����yy�S�W�G��.���f[�*��0s���9X��չ��ְ~�!U`�X��m��=��d�ѡ��\I<ѹw)����|}щ�(����J��La̋[�Uh�b������i���G^���.�7����s�Kbf͘z���~�7�w`Õ(�}� zCu����2h�|��^��a���a�+A�+�&�^��<kJZv��2-̖jIX� ��42����S��+#w��cj{��A�*���\�W+��!
�Q\Sy��[��Am�2|��^2��D_��+$\BB�C}�u<��;ϝ����+��������n4
��.A��,��C�=rݱn���u�S�b��*37bam��-f�[pNj�N�A#[�~3�;�U�^��8-����X����_�d�z(h~���&
)�(��q��m��Y7-���g7b.�jRy�)�ʗ��r�&e��d��sό�b��5ń*���-Ԛ)�vO`+ّ�Md첦�XjeɎ�ټ���|����A�]���<B9�8P��͉������(躕_��]L
��<�uݜ�=���S�[����z5(/V�������ݿ��ʁ>E��:v*]�=y��1�M�N���^�xb�{�8��+U'Q�6��{�\���^ь!��E7�anQ��Jg�P�'[9:�]�*��[��1'r�J�	9HҼꄼ\�t����S%���N�6�yg�$o�2����kن��e�^��%k�am~�=�f�o(���s�<��13�/��'&n<����"����!��6r��umw�@d-O�e�㒨~�?��.����]?5�C��jQ�c�gx�������eH��O�(.��zcp�^�O>�d��Q�#u��m󻇟`EX�\֥�د�>W�~8a�&��}-=Qyr��QH+�QN ��$5Q눩���>Yu,�;ub�#��q��H�|}ĳ���"����zD�������b+ ơ��}X�`y���N��Q�u�)׷ZVܾ0��*�/Te׶[�(R���Z�Z���*g�v��( r� z`�HyM����n]fxg�꜅��e-�v0�Lz�%>[r9�K+R�b|T�h�8k�?m�`��^V�}��7�3�j�׸��Zt[�m��\y�t`��tJ-�R���
#e�C�x��ӫM�;��t�|t�"г,ْ�	�o9l�m���p�G;�rf�iܷI�fS&M$���a�Ot���B�#"���3�	"oc�Nj�d�F�Ơ�I�	��N�^fb�3�<W�b���d�L"�ac����i�u����7��٩n��S87f]%
K��8�
�0X��bV�0�H���p�}p�;&:�ŧ+bXF_ʏn#�9�Zo o�}�&���s2T�D%fXJ���ty��T9�"/8�&��l䡾x�j��*c}�,�^)Nq�����}��'oe=|��7�f�JD]u�i����"+�U���7g.�aً4ˠ,��q�ͪnD�b(K`@iz�헳o�aX��;� ����J/�Y�cwP���=�56;e���S㦽=��>(Ր^/�ӗ٘�	��w"Qx��h� 6T>=�gP�呆j.�z�W\w<����o��D:�_8�n�Gj���e�?]Q��
������/!�J/���bd�Ҙ�6 �]��`
�Zݐ�ҽ�/��GyN{θ/=��՘s����G\i��a0���/�#hYK1D�θkxd&~��5AZ�������\�+q�C����s���m~�,�x~�j$��/�����h��݈��{)��.���2;�iy���|�V_�*;e�V�l�2��I��`"ĕ(o��t�GOAs��dP)MEE��K������5�Ov��^�],������`p,�%T`@H�<[S��7��.4���*�&�Lazvu˦���6�+�ߖ�c%��x�>JT��y��nϚXCs;��G8�y�3wu]/����\:����|��o�-�wSE�|U�r�L�S�$|����r<�9h]y~�9�;�}�b���'�jt�=^b�Ƀ���6�C���X�2t�P�GQ�޾��f]پ��Z�TT�������>��i�E����\���\"��?nJ� ���͠�8Y[��x}�cT���XJ��Zr�I�Ω���TY:���|}|�CF�!Q��~��zgx�-��nF��r����c��ȑ��x�zY�$��꒔��"e������F�>G!=��[�e@���SY�I�Փ5 L��ǎ���K%��`i1\��3�V
�=�B�Ҵ�����/Qb.^��i[&׎rg�Y�mY���H"yBg�M���l�B ��2�����ö�<WB�,6�6>��YY9u.�U��o��fi��r�/=h�1)Bw>�V��ض�>%l@ɇ�wL"�u~$���k�?���L�:���9��[�BW���:���V:�?�~����lч���-4=I��յ�V�vئ�g�V�Ba�[��h�aX)�#����O���)�t[j��g�.��2���)�ʊ��ͨ����X�:E�,h��jD���sZ�YW����3����45w)���Wc���	���BZ�TE��@�s�PO�>��K��#�x��D���Vcf�{��UX�	�I�Jv[2���1z���ş���2��,]L���C�o:�{S;�'1��]F�
�6�����w9u�d-;����tfmTy��Ϋߓm�[���)	�;]h�f�����}ˌR�ju6�iۭnS��rN��f�\�p���0�PHc��X�'����H Y���v]����[�]�o�_v _u
�e�:�|\���Jp�|ȧ�P��(묮�zb�ʖn�z���K��=�=e���*3!C����N�]*K�k`Jm�0HWo���[㎶�qD���%0.Le�8e���� j��LY���9�iٖ8�8�Ҭ.t_2��O�^�{��2�e	�ʢ"�y��u� UC�Κ�O?���-��h4S�+����!L�E!�9�y����6��nji�M�bxW�H.���� <�{�A�����m�;!׭�l�b��0E`�X�س!ƴH����`N�-׌�Ie|�Hj�u2W�и�=㰏�Tm���ַ�Yt���V�OA-��N2^x�dNbP.N�0������DmK8������M���;tU�AM���v�O,�l�y�� ����j�����~ːj�z����-�2`�A�|��@�����9�4g��Qʹe�Y�U�zfK��=h��;�T� ��+�p{yL٨�۾��W��	L�X�qO�x݉cp�-����m�D�^�E�-��[�z�UA��{G���KV�;R+��d����N�[�����w-�=ø��@��8\�:RV*ȧ^"Ί͇'V�^�[��H,�y�v:����6U�_xosiy���
%Œ˴̛�Wr,�y �Á�u+�����tf�oY�j^Sv�>�i���r��%�9L����(��%�t>����WO��wKBY�'e�{�a�Yb����S⌈�e</���L�M��!\"��m���l�rrN���U���]L�@:�і�t�6h��bj�T�6:�8��B�������b0�2�J��3 �6+ �|js� �B���\�^q�N���e;��S�[J�IűG��e'^�W+:�ڲ����)_�a��5��K����ή;�����%�z)U#<�5�������{�^���)�,��hxv:�Bᬩ�
�^2U� oP(�$/@�:C���&q�{:e�B��jujY-�b���t%�S+�5�=��P��yā�����2��)��T�s�.��NhV��ҰS6(t;��V�E�����qÅvuGo��Y���f�9T`HR��Wtk��B�R:���gT��{J�t�ϣ2V�:�gZ��z�Դ\���y�_B�*�2�7�F��-�A�x��v{QĨz��j�8g�˧�����l��YZ��T�h���"Ux�Ͼ���Y��L�vb�V8z�X���Bl���[��3V�E\���y�qtSZ�\B�������qb��l��b��s\g�����m���y����ƣ�SK��M
�1C�!��;���_���P����
o��$��;������s9��9�?���)��y��h���>�"}�1N��Iw�T���B��trཻN$��\��m����t��҈������M	�p��I��R�=^ o���%w��7��E�BAYhFM�gE��D!/M��1�Yױ�'5d���%	��h����w�b3�nM���Dew��~5Cx��;
c�H��h����JӢu�x^l�.��{v?ps��k�>ɾ�����C/f�=}J9�d�7"[�%� 4�=Cv�ſa�b�N��3"y���
�3-�=��o���i��$VSU�/�:�ʬJ�u�p�*p�icv�3�sL?<%̹`f\�׼{��~�戞�<���]-���J�q]�j���ˌ~��z��@]���v���#c�u�Jj!0J�ӓ:w詗�VD� Z��*�/zM�[�3%�k̻']{�{�"�AT�k���� ,[K�U���zc��<48
ÖN��⩄���)�9�V;q�{���U�n!q�$𿯤��2���3��>S�Ar��������1���O��/ҟ�H%����z;z[&U쏺C��͗��Xq,��/t��%[{�Y��F����ޥP���g����7ʫ�(�s�zSc���wWO /s ��\�B��D�|�ެ?���\Æ�t��ku�W6�u����Xp�A���qދ���9���r�Y�q�ϋ�E��Y�� �A��>E���H\u�z����Q��䨞��vֹMWҟ9�s�(}��ovC���|.K,q%l`@H���ʗ�x�<&,��n0�y�����;OM�u�<�ޛV�mi2YY׋�J�T��'Ł�A���E�;�;=���w��x��}-�&�l�KB[Z��/���'�ч�*g��&F�6�,��ZUR�%Ͼ� ݐ ��W`�>�F���׆��wB�	�Xm�ލ�as�����Ҧ}<]������c3q2K�?���"~��B��83GK�|��sj�$�{�m�-�M��jG(��%�9��>f�
�6��\�a{B�.{Ƅ��5���zɂ5�)�Ƚ�<��Bj����v̐�˹H"[�&|U���l�B ,�=Q&X�a����_�=�'P
7{tog�W�<���xu��w����wB���1,�'q�ک��b�\ 0�CnL��b�j[z4�|W{�6�a�1G�F���0���ɹOZ�X;:�H��dS/uX�W�#7�� ǅ�SW�Zo��c؇��n�d.Z�d�#��"F�ױ��|�� ��E��"�v�B�Y��Q�6.�r�$ЈN�np���PY�Vn�QB � ˍ>B���W(�ì �8/!�U�������:�I�)Z�+"�TC�NV%D':��P6�2KN�iqԬ�z�6�����.�v-[.��[��q�r]�N�WO[�a���e�(ֲQ:����]�E�S.����z�E�=��_�bm�A�G�哻]�ol�<&�|�#Y̌j��-#<RR�O}�6പ0�hLٿymr=�S�I��h,N�Z�`�^���f�ʶ��uױ�9N��X;�*zzS��KC��ڕ���o�p��sts�E+���Z�<�7�(�`YwV�Is�WU�`�y�U,�[s+�5�V�m�5mӥ�4y��c�^�{�����.�7Ն��(�eёxTs��;�"?�CPZ�g@�VhΫ�#'�ImR\����=�K�gQ�z��5����U	�]{��;�(f�y�z��K��*����F8�^�YC1օ��r��y�f_ sc��.7ײ#{8_nh)�q�I�Fe۴RZ�8��K�}����TH����T�Zސ�U�8��+X��}
�Y��b1�u����O�f���L�s��b�V�s1�fx^�Ψ(r�C�R
���iI,}}$`��X���a���P+n�{{�\Y{;�u�g��B�b�E�1U�:+���f#sA�ns��Ӄ��ҢM�Α+.�&�yy��Ή�9Ǭ,�$����)�V�t �9[�i<=��#%}���xUܙ����\�362-�{�?bȌ���|���"j�3�o��@����/%w��W�Mf��^�>,ww<��$EVg�sx>s�XOc�4S�X{Ȭꨡ=��U���:�Z�9��v�w1���3Y��"�rG%��I�@�fQ�z֭x	����'x�)���ev�z���B�/J.B�{����Ns���z	�1'��:����XC�}!}7�����d�c��4��-yӃ��sW��\}����v�ᅯ�(du.��3wb�[����E,�̙�8y`�oM���wQ^U�Ӷ;,lH��b$,gVX�hY%FL+S
�]�&�����T�Ko2'��)'z������������*��ُ�y؂���gn�
���}ev^�۫��B�@�}#��2�}j��gjs����Nu<��h�y^ݬR��c��Os�Q�{8n�K���t9cz��VX���D�ۤ0@�1��v���e������Vh������m��r$	�o����֖�14�r���l��z{,�͙�������j�S��h�h��U�Si�q�t`,3�6]KI�����I�}�rP�c;�[|s-�f(:�)��=�C$�o_p'�e�Y��|�:�N���<���9#	�m��o���Au����e�eX���sȪw�b�3�{����b>]��^ǎ�P���$�+��$W]�H��Y�����)2)�L�ˎn\�ķv䈡�0�9r;������+�uĉ��n��(�"+�% jE+�M��
hء.����'u�$�$P��r��D���� � %�Nn��rd

]�f\��$R$�.g]L�`I���0I˻� �s�3e!@�������g:QH�n�Nqr�)�sH�]�n]wp��wD�0�N���sm�BdwvRQ�Q�Ih��@#*D��uq"�]$�����LC1�t�T,�Nt75уL���R�S�����K�w\1Hb�F���DĒ

�h  �	��G�gt�l����~�F��y/?l��[��Ws��{jcs5��&ӥo��thVmQ�p�4)Žكz���էV����R��~�j����t��%�8T.��}������
�qO���t�����=�5�m���Gx�eCaVϸ{���9��4����4N	`cP)��3�ղʽ����-��� Kq���b���#f�G=�o��Y�|�����'N��Bg���:$��Ge���լ��/��f��W�;�2S:�6���Rw�St�e%6�^���CĤ��,I>D/�G(�Ɵ�{�9T�.0�k���Ot܊CaF���t���F8KH�0��:vSa�w�PnU8�K��� �	�d�+���v�`Jm�4$.��w��c�s�[H8�Y��4>Z���z����yD \73��������'��X�wJ�^]te,!���zl��'��S�뱴6;ו�3���9�ğ!��@�z���G!ߕ�\�֑Ϗ�<W�0b.=�<]N_0C�iL=�U~2��PGQ z~���}KF��8�swR����nJR�ט3֮�!֧��Q`JJZ2|T�����!���D�^SBY�݌���q��f�A�5�����	����D॑��;}�3�����T7N���}_�h��4/$Y��G7s�����"���-9k�9Y�V��f����vc����z{��4/AۓD�q��t�#P�L��9P��[ۂ9j��$r��Մ�L�ԣiF�+��,TF{�_�}�g�#�8�~aۨ��rz��j�<e�B+��]���N�v�
�Df��:�}��<�[2^[Wd��`���K'����W��>m�~��&
��7b���,�U�v	�W)�.2GZ�~;�;�\����u�ys�����ϤFK'k�pw;8�7bM�`Z/v;�dܶ�"lkv"�4ǵ�=��RQ蝾�~^찇�f����_�p6t;���ۈWO���/��\z9��=�-}��Y�����f�6jc�9i-����B[B��:���b�W�vga1��4�r׫��c��Jw����c>�R�@.m��5z�^�T�Y;�fW�|�Y��-���6�����]��G�>��P��k��m��>ҵRqeCi��{�\����F��l써�W���Y�)��aYI�tF(w]���~kH�ֵ�e�<�h��O���^�X�(�i��Sw�"F��CҘ��YI�K1��qó�n����Mju�R�lr����� *��)�Aӳ$�un�S�~�:r9���*�C|nV\7|�و o��DbY�N�Ї|�u&+��;<�IN��׵a܏�:�S|+.�N��O{i����>���u�a���T�:&��Ӱ�y���μ�m=�p\��ѭ�[;w��C2���{=��Y��<	=_L�#�a�EL�1}uR���U��7~�wR�8��Q)��1�E���j��&�e�)�A�8�Y��UXJ��r�E��⢳;��p��i�p������7Ԇ��X��d�+R�r�T��y����wͣ z`�H��ϸ�ϽH)�9z�#9�Jz�[��&�S�����l��H� ���KD��@�[C��ċ�9�)�X#q�� 	��î��[�[�h=�r���#�*B)�̒8�*��0��@y׶����DϞz�ϣ�����?N�DI�̶d��=��{J���p��^ o�T^��~��Yw��'�^:��V)�h�R�G��K��8׿ff�`�VYo��.%�Q�ZW6�9�vȁkp-.����-�� l7���l|=8=qR��}^�/Hۇ�b�'�:���گ�gW�&*Ҏg)M��T"E�@kPn��ٷ�c
Žu�#=B�z�;�V�cD=y�x<3��jn�_TS,��s�6��F(KX�.��E��`���&�I�^~M�fY��;�H�ՍӖ3�KrmY�M�,B�v���������L-�M8˶8�\+F^�ڳq�G[O!�w{˷����Qu��=R.�μ�ew�Y���܊�7ד&iA&�{��v.��(lp�Rmu�Z����|��zkc�0&0���ܔ�宗Jzn%N8��G[j2����זk�0��XH8��y/��qxCu��YI�lI�H�� ��
}+ޒ���9�	�yq�{�iT�/��j�����p���0��l�#�����l"��5g/�a��7!0)����r��a�-4p���wg�������Iꉔ=�y�L�L\Es�\�頽�q��ٌ<�18�Gz���t:�2P��\Y^��z'�6�p8<�ȱu*��
��Rf��MUeC�%E�7ݑ�\£q��\�k�)��2<�j���e�"�e�y��� ia,��M�e:��s�Ԕ��G��űS�Xw�r��yM����9i2|��ŉ�R��3<�@��{&��t�đR��Vn̯P���3�0w�Ā�U�@U�}|�Z%�-�zf
�ќ����h�޸h!��پ�]#��'�2zk� ������>�F���	���m��L�x�z�g��h���i�B�������z��U��Ù%�U%���I�P����F�����|����15
ԕ_�_�3>�bWQ>�� ��V��&�&p��Ցz%�ټ�Α��K�ٮ�[ܺ��hҚ�kx2����z�l]:+�w;�3.NL0�fF<�z�L�nyx!(T������ݕs٣�p��R������>���^jHEbJjV�����x���s�����$T+�= �^߂������2GNCb_���1�wkLf����8�䴒5r�D�ϊ��Z�" ���az��xT�D�Z�ʣ���Ô��7��׊��f����2��L���Eф�w�Z���8��ƹuȝe���8�t>6ͦ��2��؟1��ovS��)�Q+7b.��F_�"��w���=oD��zbU\?&���C�@YqN��e�T-��X+r9	�m��s3�%���:Ì�-�A����|� E�h)m�ym��9	ŋ~�AE�ED`�����j�dX�A�:��]�ٗ����<�	Wc�Jc4mr�m�d��w3�W���X�'�芟Q�f�(M�]m�T�w����Q%V�i�e��8��g����z���Օ<nωJ̱� �dQ�ɜڂc��J�>�|O2��Ei~O�]uXR�<�dS�(HgR���j1p�T�qx�ܻ�����]+5*o��G��S��S>f��<ybq��F��s= -n�z|�k��8{�T�p�P��]_䂗S*o �����ܲ�T�JR�&3����ky�{7�����jr����|u��/h��@O��VtW���en&V�W:
���5)�)>�zXS�;i�4m�,�Kg�v*%b8��l�ٹW.>�A�l읤�\����)���)��fŒw�f:��=qF[*�,�t�K�U]teya�&v<�:^&�:ì���ڇ+ئu��P������
�#�Ua����*��)��TF�0F�]0�*�0���ht��^�)��þ���q^�fo�2* �dL끀�P�
Z+*��F��'B�~h[vT�����j
�WQ`$�E����K5
�����A�h^bXM+����S��]�h�_�Yگ�B	@v����O��:0����l�0ј��+t�h��2��K����u��!ӥ��հ��Ρ;ڦfn0
~ˁ�N	��ų{^v�5�P��XnEп1	2�r݂[5\�����]��%)�:x[�`D+khX�l�sʾ��~qN�K0���(݉7��ԥ��ۅ��y�m�gx6�D���rGQS��}������l�_O�F�9>
�l�s�ᚮ��!�#�ҕ���-��sv*tnS�����fXj�$�P头f��7�P�B[BO�큳��T����kG�߭��vm�._T	���c[�xO$/'ϖ��ݸh�R-�u�����S��"�S.� O��7�<A�����W��&��5��֧˹�n��ۯ%L�Qꪮg`��}����ԣr/#�����1�s��;n*��g�L��J^>��[��]�;��]L��uS8��Ս솯Q��ʝ6�'tw�jC�z�'��x��7~�6=JkMԺ�"��o��<�Z�8��#�cz�z��`�eʝ�5L������4תV��@��qN�� 6���C���zȸ�J���rǹ�W���
N2
u�<��m�Ra[��0�3 �Y�$�-��!h�������[��"�Z��m��itck�����o�^O�ʐ�NR|���<	:��
��u�O��+ck�������&Uh�"�n�d^Gf����L����g������C�*�,	��_����%���.�۬�S��4���ק�j�=��C��V������`p;Tdo��w���H�W���t9a}JH���`S���>�2 �:�;}��|�KF	*T�O�@��{Ł�=.�/�N>7Zӳ�L��h�∟�י��w���;c>>�"}�lx����\Ք�!����O1Qa��>��К�A�!28��>���WmB�\�ƴ��M�����]��bN�tp�z8�!;-����m���)c9�gI�<fR+Z�����*p+�v"��V;]c�}�ۋ�(;��I箅{ŕğL�S��Y,���j�0�v2#���MW��v*��>��y�������XġB�H��.���X���� S���Q�HSng�%��S���h��~;GQzz5d���n���ޭ4]��{9�B͌@-�|T�	{��q �l7�£�%������k��^+n�y�=�y�Fnk�޼	�f��r&�k_&*��s8�oz�����g�L5p6�<~�*p�j��y5=��g��'se���K)���<Vuͼ���H��gF�t5��]p�9�c��Zj)�Xn�Eq��Z�.� ��<��W���N��/~^�	-�;��
��z���Ij��H^��'v���<��Ui�_�]��`
Z܇�Ҏ��-�bVPz�&m�<��B;ߔ9����.���NI눹�Jq2�ў�W_����p<�D�@z=>&���c�Ey���^k��67�Kw�)�l�՗�>�V��5u�����M/ܪS�0:�i���x�ܕ#q�}\�����}��/NG�>�Y�y�{��G�Ze���W�X ��j���@(׌L��R9q����t�Ң���7ȧ��bdy��qe{�mT��f���z�j���q���f�Z}},�������R��JN�q�����v�c/6��pTb��KX�A7�Ǽ��aǀ�ݕ�B���B��WB����S�x�iuZ�o+w�f켺w��|�i����꾼T�cX,P�:,�`16r�uR�R�H�Y q���Z���9�/�ǔ�֬+�ߖ�c%Y׋�K(~����yB�)��e�a�����P$����+�d)���_�ğyZ
��m���{��'r�����4��.o�'�hR�#�� ~�� ����"|}�L4T>B���[f�J�k:um�i�Z��9����n)�fԦ������,T*����&_�
��|tn@��1Id	a0�^�U��N���T	J���(��;�n���f:2%��/\X=�C<��}9�ت�����:�ͮ�V��'ۨ�R�̐ӫ��9@�&j6+��d��Y=P2a�Y������7�[��Ha{��1�V�Y��J��~����=R�=���!{"�w��9�PwI�˱&��o��L���L�B*W,�ve��'a`[�S�͚)֢V
f�E�3H��d���K
�S9�-Bo?]B�^��Vn)�	e�*��1��܎C,�O�IXz5Rl���
��sX܁�*�z�-�ѫ*q�*`N(U��E�K'�����~f6��I{h��N�9���ޑ�4澎)�<e�[s��z]�F�������֖m��y��N5��躽�[5-�q�	X�Et.N@�߲T�8P��D�W��B(A���:��7�V�\�oN<�Yt/mK���VaW#YD�]hK��|�n^涴nT�l^�P�S�R�ٚ�sD��ɝ���;q2�P�஧�t3t�7kk{TҌ�v�a��q?t!q��֋>l[(�3��q����1z�����)Y�23�!z=���s���KY[Nd���1�%�qt:������8y��E=�r)�^�=��#eK4xny�x`��w,I3���.x�%k�DqO,�!h�a9���n����׭4$.�~�d��`&�M��äZU\��W�7��lßC	=Pf	��C�X��P|[��q��Ny��5����nnw���rD�I��7l�xm���uL?��@�bK�=�Ua����*r �Ǧ��ާ�m�H^��n�{>V��3�m̂�(#������`?.ڳ �s�B����S���oO>W=��+�\-�E�	"�x�L�=8m0�[τ<d���_W�\,l�MAx��)�k������]yB�R��W���[��A�����je�,@7SBSd�d��1_Ou:7Z٫�U�\�����������?3��{������Um��[m�m���V����V���ֵZ�۫U�m��Z�����ֶ��֫Z��j����ժֶ��V�Z��Z�km�Z�k[o��ֶ�Z�km�V�Z�ҵZ���+U�m��Z�km�Z�k[o��V����j����j�����(+$�k/J2� u��B �������-g��)��$ 	P��
 �TH���ER� 
U�>  qTB�������%�ITJ�UI
��*�!�R�EEPT�#��D��ITI BP�*I(R*!((��B�D�R�("
�g7 ��*5�R�j����1��Тle-�
R-2$�U[i�J��U(p   �ʑV���,p s   u` h�k�  3   �pC.7t�hIT�X��� ��3��F)U�Y&����d�!h����h�i$��iAU� nᦫ�͆�*���U���[kJ�5hV$ �I4�-3H٭�5"
�����-��5��5R56ִԩ�jZ�J�a��R֕*EE��k[X�SF�mXT�T��R��d�pj���LK6��V,k-YcM[m�µ�-4eR�Th�«-m�Q���X�*UI�TVMT���:��Uj[kV�ce+V�CXP��Q��Ҩ�Z���ST�[jl��+V���J�1 �+!TSp�rj�����laB�,��5Y5�m�"-���
�hҰ�T%�"0F֪�A,�	U���0[�SQLlQPֈU�Xe�f���ѭ�*�U��f�ITV,UI��9��Ђ$�X�l0h6YU&e�*kAJ�Z5K�z@� D�����R�T�h�2�L ɡ����R110 �&   �"@L��O(��D5(���ƆԄS�A)R��0&d L!�01���$jz�i� � ��$"
=F4�@F�  �����
�g0!bX�� �bPH�/�;�D�$4�kŜ�¤I$Ht�q �QAxT4	��G���t@��V�}*}%}��������	�ETP��oP�M$������*�ʑ�їk��O�_k���g"I"C?�.�4�h5���`��8/pt�s���~��m9�`a�n��_�����]�?�^W�UYĕ�Z����=�07+I_h�A�"���W�6�hU���h#�l�jf-�B���뫶rY���l�X�M
�O!�!�,ndn��*�RW����Z��㨱�h����x�Lb�C0w��Uy����㑰�owi�/���m�U�o,b�)��岦�I�ʂL�� �ċE��̛�^�2�c%��.J�2��ѲM�Y��M p-�n��ժ�ڻۦ���th�8����J����kl������7f�=ҳ�-wVA�Fe;Ki��kh+J*�ѷs>P�;A��O�n�ø�U�[t��V�J|,����ʆ}t�j��koC�l�ne�*�����\Xɠ�kw�R���H���yj���?e&TJ��WE�����/ᖒ��7�&�'[$7wZu��¥�Ю���JEc�[�:�T�|)��
�%ܴi��P�vu����V�oH�E��'�)�e�M��v���Z�A����p��t��l��(!-�ob�z1��%�7���7I<��/&ѨoFkXX0�.�P.�Ylm��Y��MUقVU�YAf�G+�4(d�En�=C�J�W[���[�n(�U�ͺ�:�����1Yu��Ԑ�v�g��6[\i ��5�4��f�x���6o8Dx&+W��X�n�H�n�V�wm��D:;Y�MڈT�k���
8���P=�+�`���\�ǃFĳ��O-^�VV�'� �I�wIA��͘�AmM��f��Ě�K'f��3�u��VK��i�F
En<ͱ.�4�r�ߢ�A�M4*��͡��	u3�t�6p�;9\\�c����V����4*��ַ)��v,��V &�3,w��j.[�+3%0� 0jS/���/Ne��T��0��Z-�Z�D�N;��@%-�%hNެ���%��U��k��E(d�B��pL�6<xiAZZ�6r����Ge�ޓ�a��ʸ�˘����qŖ�(Jlje�-C�E#Y[li'�r�0��d���oCk5v,t����f���v�r8s�3#d�����0�E+f2J�:Y|R�zfU��ֆ^,�f�Ɗ��)d���lJ	j�9��VM���LYx�]��cͻ��ytX:�vun�x]ֹE�ˤo"���nYu+MʱP�,(�5ٚ�����gY��X35	�ب'��tk%ڗ��Z�x�Q��c�h�@mT�H'�ʸ�Յi��f�L)n�A����v�\T�f�W����	[V�Ws6�_5�n�Y�b���v�����YR��& ��3�����E/ �
@��V�o2�р�:�ܣ5�)�R��m�XΡ����׻N��S( ���up�w�R�F�zMN�Qj�n��!��vk��7��#2�C0�ÛF���nM%P�X�ɹ6�M�cy�^��-JZ�f� ƌFY��QZ����;
�%օwO,�n�Ob����-Z�3��L�X��qV`�7Z�9�Y�r�0��z�YH:�_e�{O����k)f�[͵�ٷ��S��Ak�'j�qԭ���rF8S"���A�h�M�۩.e)L���J�4��%+�-π��+F�b�ה�xc���٤,F����t(�9Rej���wOE�n���	-ۓ젳5^;���2���RUo[0�$PĳJBҴ��ȷ��s� �������`���He욯�^iͭyg/uQ���*$63!��zə���x[ڐ��N��kR
,ж�����ȥ��+�rZ m��F�76ڋ�#I����ܫN5P�7,���܎вS�k6��؏�d-�oT`Uު�U�A�X�<�v��Tȕl(鷺S�lb���w ��$qNӭ��`Km�@B����fm]ؗr��W�Ҿ/�b�"��7�qu2{���i�`��N�]��h
XHXN�6�`;�d��O	9�`s(R�Q�v�+���%��Ҏ,�n�h������I��y��u�I��-�Y�E?�5Z/(���!�0�{��a9u���&P?f�h<�*��>�3`�!ߠ*�n�i֩�ݫD��k�+5.�b�vr	��~�!T��lPG�b���ۡ6���R�������Fа4jJ�\";}r�\��]SR�ٷ��c��3�b��Z�AB��� �B6�
��lӖ��(-��,g��cz�]޵�ni������h5B��&�]@��Z�!�ǗY�d'tv�G?�_qLQ�b�`6ç�:5�;�A�<��ZYV�ws&�3u��i�6��&�# \B��&�$���dY��R�e�0�l��v'q�� ��n�� Gd*�V�/p�<S �ZA^��
hi�*��;)���5��h�5��
S��%Gk#�R'��R�>�b���4�$id��H��`��� �u��k�c,��2ӱ7�t��7���Ԓ��[%G�����bc@�f����h&[Oڭ�p�������.����z�*¼��/0�{.pK�1�!�$����6�1V�t,'z�5A	iR��9���i�9�I�f�)@-6j�T�����k.C��J�Xӊ:�Ss0/C��E{*T�$�p���z�¾�u�7h�ے��,2��(J�֒�-e�vU8�LI�En�l�V���0m��ܲ�i7�uth:A=��ID@��^֛4/$

�ߍ�c��i䌬͕��Se�W��-�iT����(�҂FQ�%	ӏM�݁.��5Y4����y�d3�n�H|r�*�Ծ��f&��wt[n�-)���j��$�4Ū�V㰕� ��Z5����mӬ��d��'�%M5%��Y�Zy��B��0�w���تm�������ycI` m���T�պ�b���'Z͞��׽���e�$�����.��ӛa���y�!a
YG�P����uS�R:�A�t��طC�{��Ƴ8�J�m�R1��0��������2[于⣠R��+X��̦w��庵�m�:l.Tl!5m�{��O�/�5k��ָ���-��}��Vd�ɼ``����w:3w4�)�5����y�Ka�Z���,.�Q7w���yBMƴ�4��v�`kY��Xa�7�`�k9Ş�V yuPO�7KuQGq[�e���"V�I%�t+i�F�2ɺ:�+LSJ�]�2�bTbQ��R�
�#�1f|�[�|Fgǆ�`���{���5�����J�Ѐ��uike�/(��O �pfk���&Q���&U�5.U��K���j�B �:0;������6�Mըv��x�6<�x�,�>XiI"_70kX^l�t�!x
�Ù�&XG0Rc�X�b�8�m���[C6�^Y{���>��� 2+�z�V�f�`�\��o�=�cK����A
}�
]�ƺR�e*.ݬ�$��0�D�x��1b8�In="��Z/�0��Yd8e�˅2*R���@�4�U��ұ)J�ӭ���Q���VnS��m��/q��T��Jl�{�E$��&��ѯ�4�onf]�
�,ЫT�!ZB�9I��],��S&��D�R�M�m�՛�o��KL�B;�9�(V�Oo�f�`aLͶ�E��B�i�q�7r�o��k[x+[8�j��a��Ǭ��9��1Vkr� q�̻w��r֌$i9mM�I5B��n�k|�}�u-��ڼ.��˾��g��x$Y�;�������n4�.�Fja���`�1���p�Fe;O+C�]&�j&�櫐WQڴ�鈜4v���b.��k#-F{��F������RڼK�Ev���kOڔ���,E�UZ�X� ���nJ9X(fǩ��ŰJ�P.�"�^m�^��q���sFy�ޝ�VM
�+EU��{U��Q�tsi��Dn��F�dwou���4�5�j���{`�J��,�ܼN��xP��4^�4j��V �d�;��`��櫠Q����3�m:8I�':��oI�/��3/�*�|�י���uֺ��;OAA_�?�~��#'���?;�k�8v�Ο��?O�ֿ��'�\\��g���G������x9"+��         �����&�Z���^&�ج��{�@                                                                          �� �                                                                                                                                                                ���*2J���W�[���2-�e:��͝�ʐ�Ի�z<�zkq�Ǡv�g:Z�纞���P��<�غ>���Q�6�f=n�a�v)S�{w.2��ً��X���5x5h&j��d: N�&�`˭����V����,֓�וӰ�~���vݫ:�'gf[(̜���-�j'�3 ��1�pt��%��uZ���C���Y]�j�Bh�6�Ķ�]��.�ښe�S(�2\7q�3��R+����=1o�8E���� ��gƀB͛��vuW1����co	��l�p��v���N6ք9,���SD�l�ꆍ9��Q���.��n.2�D*K�\�,ט)S�%��v�K7��q;.\Y���ocKq*���g&\������N�A��Q��]m�U.�������'�fh2�\-헜��s��KWBb���ɟ&87LX�W���O�D#�3n�fL�S �Y�[�iE>�1���:���]0��/9R֒�����^'�^�"Z�������]��t�=K�r������᷂�/�m��XPպ�hv�6�v�&�x�4S���#!�'U�i:)WU�#�+/*��v�xgQ݂U���E�S�wKv9X�S���^�E��h�)��r�nSv"S�Aձ�E��eY����VX3ː����7r�QWn��s4Ύ�c$�{���f��(�n�`b�P�T5Ǜ�s�<���[Q�$�V��ܗ�r�+�urK�6�iJ�|��ƌ}[�F�|��G�7y�7)��@�[Ճ��I�k7ƘW�&�:3�Z�O.��^��bR�jٕ��^%��T��:1!*W����K��n��F; :�����bZ;���h����!�X�S��U�!���y��OQ}��݊pkR�{[؜�^��d+���HN+C�k���i�R�=��������Vj�u�],�Mm���ι3n`��V�w(B�ѬRdQ��glG����K�&.Ojyk��̏����
#8*�/5�g�eF���j�|*1�0�7QW��;8��n���u)�3&N�qq$���T�D���Z�N�5��)�ڸ�1�a��`َʱ�����CH�;V�����x'm�Eֺ���	)7�E��)H�W�_H߫�μ[�/���xm@��Os�.p� ���i��]���6�B�d�K��)Iy��"Lض��;+4��f'������-̧L.��Vd��BW�*�����CW�g�*gv��%�N�
=7�+7~��B��o)�ԥ�B����s��S�zk�� Jc�}B��J��5e�']��l��X��&���y��3�d���v[I'|�jW|,��K�.��XΎ�kE�n׏���(�+��C��fOt"�5*�3�L���u�/+��}X%*����	�ӪU�hʼәEV�ekޓV1/Z��dXm�V�h�u
A`��:����;;�Y]]|�L���a�kb��s�\���@eٙARN�7&�J����*��5�U!U��݊�{�����5��Q���Ma*(E��i�V�Wbu�n@��E�ױe��&�/���������h��s��"�x�\�ҖNï���]���5}.kx/*�*\i���QQr�5�^�	K�\=|�ћi�Bt��T2�g�G+k0�kp���Vޢ11�]Ss�#K6]\�
(ş���c��s%��e�d�r3��+�T\�d���'�t-тu����p:]{t0��N;a����V�NՍi��E���� ��̋[L�S�g*+�p�����b`�W^�3����ME�sy�GoD�";�\�&�N]�
�F�3�<u�7���	�a��ρ� �-�5�EDsj7���2���)ҳ����n;ް)��H�����a
�t/%���S��C�)
Y$��.n���8wM���k�ͬ�W���R�^�Q�{g��ە�p��ǶbiWJR���|���P�/�wt��v�����;[^�����+Nݠä높.�t-YKs��6��A�ؠ��ڳB�#N5ˈ�ҭF�4l;�i���L`�)��1���S�t�w2����n�΋��KNI0w]seٜ����s�݈֜n�&�y�',��Q]D�H#����l��N�`�w_m�d���܌�}w��27۵�%i���ᦝM��p����)�{E�N��˭��a�������e�(��U%Hs.U�wf��,d��xa����w�"~�{JL��|�q�Vi�:9�(��/����pv�@ ڬm���x�%d�u�6�s!���ݲ���r��-���R6���i��Z�϶����.Qa��8=�d�tW[��լu��i[�g7�~t#ܮ��U�0w-Æ���l7T��R���z��d�j-G5�k���ȇ2��:�[��ȩ�e#�WK�Ȳz�
��+-�Y�]lx&j��e�ÏV��EOo
���k]A�ww9�N�6�ʎ�v�٭wq��s�<[���LA�Z�(ZsH�t9��^��g'�J� ��*n��S�m[=Ev3���k!�b��p,���-��9ү7:Š��Ϙ��T��\�3X�j��ت\(�z����S���l|/�\	w3��D{�C�$
iy�F5ns��0@²�� �[��	MgW,��K���v뮱�`��H�f��;���cn��*18TBR箶Vi��7�n�[���
�P�|�<��6
6m����1��r��ǓT���r��*-3R�R���q�oi�Na�Wb뭾uf��R��Z��-���oR=(.]wx�H@A��+ �sh����
��`_rG]W���ɕ6��U����T����L�|�/VUn+K˟)�W߱f��X�{3|ov�<����!��ͤ��S7E�zI�FwM�w���KOn� ^�eF�g$)'$pE�t;���#{Ρ��o�k펯��n<83��������]����t^��/��
ۊ��Ʊ�Ә��$�]�rP�z��J�f�C��hd��OqT��3(N�e�2��7&�"f%�
����e�؆4�Mѐn_�n�Q�>7hɼ����!�wS���vC�d��59�oK����2�'�KM�m�E�}������H]W7�e|D�+���F�1gZ�6 y�G��T��g9N��u&���!��Q��Y��a�/�	�5Zv��R�7:�5��5�r�ڻ�0֟����;j$Z�m�	{v��4ҷ+z�����Z�K�U� �f]��U�U�Hw�\'�T
�7:�vosf�6�K�At����Eg��H(���)��&b+��R�w]-��5u�*p,���S�F+GR��Cn�>ź��\Z����[r.B	S`�z��ܝ��uan��8�bЯ)M���:~�ܬ�q��f�=֯%�7���_a�8'���\�Fbc�Xa���N�m�Oe�L�}�|��jI;F��#��Lw��=�2���ҭLn##���Ry�[��t�ww`#k]�{S,⎍V �v��Կ�&GK;6)����2*j k�nZH�a:+MsU�=�Ë�zo,+2���Y�\ƺ�v��y��T�)� �	`ƚۭ�#���2Wӎ�t��i�nƓd�e��q�)����^�{i6��J^��1s���i���^*��}.[w0A4=��"�8��R�u�u��tk0uqt:�+i7����e�F����7[R��v"H�*�|���կE���\�n]�x��\��������s��J��su��o40мf��5��t�r�*��U���/~5lںY_b��N����)�Yܖ
�ƈ             �3A�3�MxJ����qR *�V�u����w�q�$j��٨��FM�ܕ�ʘy�QN���A%�;������o   �@�@            ����d�|8���?�o����_�D �k�y��EAT?.��Q��{��Y?�' 
��O�N���o��ƽ�����4��O���@�*:�Q�N�,J��x�[x7�4�[ܔhW&���I�V��d����;�sn	
��J�r��r���ؘ���4v�|����S��-2� Y#�۾\�q��N�L�o_CV1���f�
Ѥ�#�;�tSo���:�سze'Y]6���"[�8��Ŵj����j�3CTp,'�zYnl��aψ=�e%,�	�
Ui�X1�!ʏKѫqr��	�N9kh��6�Ճ��b
˭�`��~�Y�V� up2\s�v�߳k����^ӡ���A6Y��aNpKW&������D%ӋFd��g-�̌� �|�/*����)�yP���c�7�`Н5��7�!7c2gAˎ`�h�WjoY�b� ^޸ku��A��}�u.�S���&:�0ޛ����J�E4*��bڜ�
�cI�l^��]ڷ����k7Q̂��I��v���VR2��(e����X���7R��5�ӫ�@�^��f*v�e�-g2WP���a�R���{�yñT������RX�.� �[jV��e�%�W�a�T�>�N��Q���ֵev�qn�i���e++�6����	��ٽ�����KS
f�j�6N�ن9y�lѾ�5�]\�N�"�X����O��r��u֦�"��]��wr�J��yH��f&�N��)�-Өyض�͵�M���:ܧYD�z���&�;��,�A��7}\��$����s[t�`��b��dh�;V�}��m���N��M��2�`��V�M�����Ya0��b]d��=�Q�]�ɖ.ž������9(��oc�j���^e����zN	��q��r��%T,�5f-13q����0
��Ƿ]���ӷy{��� �j��u��|i$,�ٶյ�;*q]��de�U�)`ulB�WmW
X����F��ժ�a��\|Vfhj�rM���d�����8�*�aB�����qYA��
��ce�=�"��ˬRI#��dJ�e�yҦ�j���n^5׊ct~HX�R��P��iLb�dA�=Q����^p���n�7��
D����J����5b}�/3n�(�o)�Q�/	��/C��Ekj��W`{��� 2n_a�Mv-[�*�;L�
wV�[�X,7�hi2�ϝd����9�e����T�=P�_w[-�u���Zޚ�8#�|�v��.uu z�Wk ˱�VK<zö����.h|;.�d� ti6�W�o0�9)����9�eJv�ot��z�^էe��ޭ�>��	�SE��$�t��n����F�;�[�M���Id�І@.�1}��y��f��+C�f
%�����a䙽յ׮���������oQJ��m��ZFh�Ĕ��lP��8�if=αB�e��[Tˑ��L������zi�#[�Fˮ4�.4�:[��oU�m���`y��{
�w�)5�P'%]f}�������b�b���SuvA�����4�Fe�=�ʵq�[\36���+���֋�"�S�Rœl�p���M�WuQ��M�Q��ə��[U�*�k,��)s���s�s6�y{ʢ�Q#yWQ�uԭ#�L�ut�'m�tu2����S��(���Ls�D��b[��JV�uw�CM�|���#�1՝�9b�U��1;fgD��IkX!���\��YPr8r�h�5Fe=��2����KwZ�d_nf�c�f%2��x~�;i,-b��w4�U�y�I29�ge,�v�nTg�]�L3umY�A^]>1CӶ�����q�!N��e����/z�.���{j���(��hl��#HiAZ���P��,5��5�+w9ӱ$_)�*0H,���^�ژ�I᠄��]1�h6Z�8��M��z'�j_P�ق��v;G\��f؆��j2������Q��d���n������3�!]�6�P�L�����%g>9M��֭��F�m�\C��A�$��x�LR�VvKB�ܨ����}�r�����p�w��)�#�[)�|���&V�2�Ng!t�i}//>�)��a�y���Nu�YwA�.�9�p��]�[�8�1�-{5Wk���E��^Sf��]&�ٷ��YQጲ9���2[���jN �[�:o(0�GYC	����nZ��K.C�i&S؍�)q�9�83rcĆP����ʱ�Ev�
���:'���'��&ꚺ�	���E�:/�Xshn?���5�����nR86�*�NP��qa�yx^�5j�՝{i�76�{D�c.���2��7����lSnZ��E��ܪ3^�Hw�1TQ%ң�y���݉���]Nwn�]��s��M<[�%���*Yv�e�B- 	�=K��z�j�Zr�����%�< X⬹;+/.�݈u0Ժ�S���"ע�
�^ۦ��J��P�K��X`7�q㙻ee�����F��A3��f���B�L^�+S���
8h����WlA�Kծ�D2q͖�Z�|�d�V��f����vUSf�e�����-n�u vI`<"�B�-: ��r��l��3���9p��	b7w���x
�h��z ����"��Ӗ�u�M(3b�5n쉅�T�S��(�(�nY����/��t3��J��HR�u �M��3$���RL�8F�����pVP��CD&�l����
\y�qޕ�M^�|�J�Nd"�l)����Ӗ�AwH`�Uk5�LTs3��^�:�T�Y%K��y $	)�8�<�o+)9}܃�fT �Ɵ6%�L����[k�޶�v��\\�hH�			\�'Aѕ��f�v���SD����$k��<'jV
��,�r��1�W���pƬIl`wLj�Jb�7&���I�U
��HB��O����֨���U;��˹F:�Y(U�ռ^�nQ�щڗo���)���F�2=��Soo7�t��O
=�!�X8�n`Z��+,�f�r��<�]�w�:�t��8]]ᨱ�.��:ʻ����e"���2�d'�"�o�e�x�K�/3��D
;pl��z�R�d�.i��r��1�[�4�mU�BCC-l.�=�h2��Y��WJ�W>��F�(d3���{t��Q�X���&�	���nF�9�:��
�"gb9Fw��.��G��w@C��;P/S2�����+��^�kj__*���(�BXFD�U���l��V١|�H�A@:�*.*����8XϺ��w]��+GJ"g5xR$Hx`�(T�.4n�������)�e�����bK�e?��K��$ݫ�P.�hR�Dh�u^q��jts0�n����m��8<��43�ռ�N?F�L촫	���n�c�M�8l(��/�]RXi�B;����k�����-�z�]��ۛJ��.r�&�[�B�V�r/�ՠ�t��:c�z�f�5V�L����2����ĦX��ۮ��<�6 �Ω}Z����%]�:`1��g����}��v�)3l����B�)�s�]�x��$�Tn�`Y�3z�I9[ٵ�V��VȮ�I��`#ӳ[�U^�y,"8(5�F�H�u���%$/����X�b��듔	gڥƮ��,W�ī�5�o�ۦ�WR�6j=[�]�b%Vh޵Zf��9��KAǘ�`h���ͧ�l��Y�㏅�Y�)��H45e�f(���M[X0^XJ���R�X�}c�Аj����"���{�1.а��*����=Q�����*f�)����:F��~45��l�qQ ��qAw���;r��&n�S���G.7�QF�e�ש*��W:K�lӤ�A�sRJ����<ayZU�C���N��.B���������6]s�cH3^����œ@	� Qt|���-;Q�i�^�?`W�N���ᕎriK��aX�Wq���V����,C��]����$,��D��WHU��Z�m��5�?���E#_ևjhB$��!�PW��hp��Ѯ�樯�/�                     !-��w]d�Hz�q���G�k[�\Pj=p��B���:m�V��13�h�v�f��V$�5>�b�ͩ��͆i��1�g ���[#�F�}E�j��c�۷���d����JD��R>`����$��٘��<������8i]�+�#tz����z����'���P�We��b�f��3V�����N��^�dV���gi��F2MWP*\��W+鰂�MLJIh�W_��ss�[�vK'Ψ�~|6;���\�ώ�����l�N�ض�tJ�%��N��ͮa�F~QՖ8�D�G,�b�;�;�g=�؍ZN�U��Br}�"�����1���nv��Sy��)����7;��5�B#d�5�+x��d���ե)%���}��h�@�\��qs?}3���1;����S�ƌZZZb��JhZm�T���ʊ)�r
Oa�(�h��(�V��##"���(������!����1Z
"%�i+Y��"�
���1T�d4dK#J��-<w�q'��E)Jд1wd5HPP�JPDR��O\�� �i�A�
]�$�5%!��?isѾx��K#Y���ӆu7�$���Wɻ�C1Tw���Թk��+�]r(������H�Azn����F���{c66ڟ�ڊtνi��M>X
�o]?;r���@���\aW�g��4Ð��_[UUu��ᇡ�*�Z��7^�lz
a�u}[\���C��}37ާa4/�\����b�J�%{8�/D�GAT	�9x�*�/��v���-�g&�K�o/C����MY=^��m_I��4ʹc��{�SyORd�[��8�"�ļ�f�}�{3�j����AޟlX9)rI�ϵ9p��ZaFLu�������?_���o�����������=V�m�cT���V{��ζg�%�4�ނ����Q�ų�vq�
�XØAh�$���q<)���|m1�d]����(�����������՛ɫk�-�[���=����E�}�����	�Mj�w
-}�i���S�������?r��3�]1����w�V�gX'd��l������������P�e���r={�4ӘG���;�/��o'�.}wH�nv�ҹ)��]/+}��YZ5L�p��Vњ�Y���LG�`��Ν�e��{;���C��͛ɰ�J3�.��C��h1����l轸ϔ����U֯g��SL�a�׬����zACVtW72�=������[���q�:�g:@�=E�Ӡ�����p�%R�n�C��Tl�YZ�Y�w���_Zc>1��+ލα5�bfbh����ù������1Z���S�5zǷޏ�3�r=���c���]����T��7�zkbg��5�/�0{cԫ�3��z��
�K����/2l����+f�S�S�Q����D��K�ق�nB�r��c�3��t�ֹ�[���-�������5O>=k(�i>;tb�²�Z�����ȳ�g�r��+Ӣ:sTʽʖ��39�)�=�vbW�ZʹW�_/]J����'�9��Nb�ć���:�nc[���7��3�Bg���~����i���	���׬z��G6dGy��\C��������O�/��W���'�"��g��C}ؚ��X
�x뢅�W=t��KH��n��d�����+rMS.��ר���M�G}�v}H���qFV�ě'G[s��r�ޞ�N�-n��w����i�4���.&����S9�{�n����4��3I�����:Ip������� �׽����Fj��S�7�}�'��O}>�̗o�OՏ��t��7-���i1A[��1c^�/eļ�_���b;���O�y���bot}5V��*�V�,<��=)9۱��0��F��d*s��jǂW�N�~W��Q��w�*��1�u�'(��|�Oc���ۊh�>��z�x���������_�B�:�X���ok.�����^nOJ\D[�K��/��$��3x�ȡ��|Ԯ^��j+5�Z�4���l�I����y>�Xb�����0��NF��ϣ�em_l��q+�TҊ����mM��#�vթ�|�����Ȱ���p�'��ؼ��X.�!t_�&k�i�)c�����u�S�fj�El��ʍ|�S�U����8ս��W�����R�g�o1���e;��W�4Ñ;|{ֻ=�0��FT�몛����x4���V#=>
yr�ƞ�օ<<�<����_��Th���Ȫԡ�B�uh,���O���\��W[���ҭz����Rt�h99�n@�ځ&��q����#%gFdp�H�s���hc&�yAgj܊We\zVV
��v����{�<����[ؐ,T��~E}��Y=^��>ӎ�j��� �+1ݣ?A7�Rgvܻn�����������=���� Fk>2l��9xc~�|��Te��=�Zf|P2nJ������ޒ�&s�8�ӹ]#Y�������#-��O��^�+c'��*ܬT��>�J)����*����Z���ϭT=C<���4ߦ+�%7�0���s|��J{��m��z�>��q�+�o���i�f]���s���1�ܫ�����bO����~}�{M�˻G�[w���Yg�����/c�
)֮G;��R���6\����X�{�7҂��q.�V/%!�r]��!��óۙ�9��o��З��3�����'޾�-��@�`.�ck��ӹ<��糯��{+�W�ra:~M ���T��&|x ^��&�R������
�^��dl7H�'uٜ�:�A�m�ǯƩ�)ڎY�^;u��ؐ�_{�e�c�m-ٕ�*�,kg�����}Ԥ��c��	�W��Dןk��^��_X����=�6��Og�/Շ{�M⛨��5�$٩�.�Y��Pg�c�� Q5���w��=~����{���V�Z�7��Q� ��bU2�j�������ɛ�Z���O~g<��LSlu#:4ܟy9u�S�NWf�n����D��H�s)�.�¢ێ�A�f�ң�N�B�b��2x�����!F2=��t��*�y}� ��>C�%lm����~	i/f��A�n���_���5�W=�׹�y+(y����OTxt�_�]?'�گ;����s��gk�~�$�K⣾���9]�N���T�ހ��::���j�QV�߀!x,g�ȶ�,n����{���S|���f|b�j�Ȭu��UM�3�eغ!AТQW���L4����]_�����V��3�����2*���>5�V��y+�)�3��t:��:�Z���.Yæ��#5p_*3k��wG���nK$���{G�u���vrKY�h�NT�u��+0`L\�ڬ�ښ�bH�j��a����{.^w�����v��Xຌ}7��1Z���{ywƴg�3E�I�0��t*s��⥶4`B�}��y�2z�AAXV}��gz$T��{R��"��m'�c�9eF�t��N��r��#%���9�-7<�2}��9ݾٶ<�b^�c��=���3Wy`U­<�R��mv�,�ߦ��A�����ѫ�.�r�����si���y��·��T��S�^��n�;���O�~���v}��a#��������6�i��Owk�Sm|U�Z]��mڮݾ�M�c/���8�r)em�C�2Z[�4��d/�.,^EG&-I���S�j���cf�F@_�=.+]Q�6��|3v&�z$�_g'^oަ|�Q��"��~�PW��������E��W��������E۳Όn���6��RL!��m���̋ѩLn�58]�e�z	�nf�^1K�p�zz��DLN�>�I5���<�ٓJ�ڧ�:,�P��ߺm�V����\^uF��n�>��2o=�4pF_/d?!��;o�E�^'+<����}ŗ�}&�4���F2)\����}�͘�3A�����Nb��[�������п�����;��_��V�W�̞�99qՔ�p#�]�Ά�,�S2����wI�X��N^�}�&I�v�Y�(vF���iJt-�V.l�gD
�
%�һ�g�a�6W+�*VC�i����6��*985u"�(U��5�X�5���;+f�Aeg-5zjڂ+ӵ��Fu�%nb��o:���еՈ1�u�pd<��F��1&Z�����8Gt�-M]�r��J��xo��B[��X̚���������U{��`�K���I1
���,���Vݚь����e�RI�	���D�A3�������]��]na��ԧ��R����2W�	��t��xo@٧|Hfj��wf�8\[Wl'���P���\4ŝ�[�c�NLgk�L3��q_c�X˾8iLDCd�gA���9�wg�����V�(�q�'﷠��Qu�/����                     ��Z�wb��>�}���ט3�9��9:+�dWc�$uKl��:�-�i%��5Ӭ��+X+PC�̂�,Y{D�OE�:*ն�U�'%l);Gq0\�P���Mt��*V�\�6v-osw�5N�[��šg�k(,ҾP��n�`BcK4�ٔJ�wj:4��P�2��뵘^�̝�֒PV�֜;�δɗ9�ε�L68����T�)`7}��&�6���Ѣ������رkɗ��d�P�<�v:�)h�--޺{b��gw���z�
܀<9� ��ȱ�ӈ)����j�nC��v[N���w��q�͠��X�X����6�E�u��K_	
l�w�Q��������x�����P<|[:�gd���გD#��|5�q7#�;������ߛ��>y�ӸJ
���"B��
�=�M�@4P�R4P�Q#M4U%%�4��ɢ����eʅ�����+!i�))5挦����EE44�KM%VA�'2e@D�$HT�SCN�uR�ѐ��CIT�F�)��r%IK��w�%'q��C��%!ݒ�4�UAZ�pwAKBQIIUEP�,EI�D\`亅�X�DJW���I�k-e9�"�M����h�a�9�윙��������Wz476��m9�ߦW{��{����5<��Zˮi�(OUd:�)z~�~ ��?~���/�]��Ex@�^�cK߿�����<k�n��M\�|�ߚ}�/>v_?"S��)n����Y��i��;>�k�=<�:1'����,��q`g7ו�Z���w��M?~�Vi��?;B�+4����Y��v�u%�J=Y���Jo%��������2�N~��{$+�U{�詖��<̞s��X9��[����);z:0�l+���~���;��?o�|ͣ[�}���W�\|G��V�sr
�#Y�Eq��.c����G����W|
��
�{�5Ȥ���7>[��a�X���z+��`S�S�
a�$QI��v��/��ܴm���c��n\�g}8�z�Ʂ�'Ѝyuo[?涹���^���g�Y��t9��6����qoy���_�-�h��&�2�;o�
nv�}^�n�aL�jTvy.�*v�KT��^��jv�y�?zV��차xż�~�L������������7��]�U�_���q+�h��[�.����+�k���S�p���y+�Ú�tW]��rG�v��G�ا�7���?�o�en5	o߾�_���1~�#��;��Dn������u-?ы߽]_���SY@�Z�7�w��\<7rZ�w0z��Zչ�zW4�i���S�a��5F����a~���(��ة��w�n�;_����9��МL��el͛PR<��������}_W�}�q���x?�,�ex����J�wZ[;&3��闐�qK_�j���v.POe{����LC%r�S̋O/*}F�@������_Y��m���]O�9y�]HM���%{q{�t�Vc8
��\EC���0^�B�\��u��n%е�M�Ͷs�6�]7�����ޓZ�%W��HW/f)��x�|ү;���ԏ\�~<�~��3*�En����II��<-��i�R>]/�gK
�QW�{
o��y��%�����q&t�o9c��ie;�5��ӛW@��:ч$v7�p��yW������[җ�<0�;T���ws�����^,|rY[�Y��EV�Xŋ���Kucrgp��/�������X�==}�7���2V
U�Ӯ^�e�M�������d���5�욻p�*aW<���b�2=o�~k==��7�.��H��]Z��[Vkm�?��KȾ�����[��#�Q)�&>������V�w�GO��q�Mo<�!�r^5��.�Z��q�J�W2��%}��a{��7��{��\qם���5)��o�e܁�o�!B�Z^�5�>Kܿ\\�q������S�Ms�{'s�q﹬�}�o�2WQ���ܔ��� ܺ�J�'|�r �Z_��:�#ܽG�|��_B��%�^a�o���~}ߛ��8��;��(:�(��%>��rBP�_<ޅ5�\���-/��M��s>}��=s��w����bu�<b�<���������_c�>ù�9� {.��]�������^{s�~}�k{�{��G����_g�O uΡe7)�������s:�$(y�n]���C�|��9<}N%�ƷtX��n������N/Y��@Jڅ���O���E�����W�>�`����^����1x����a
��a*��#�h�|	䢺����7���aOa����|��#s�z�<��L��^~��`x:� �x���x���/��}�\��������}>9��{��� �]{��Cp�d��x�d;�|�(�ة��=�ܽ}��B�s���l�|���g�^�㾺�߷��p�_ndy���_e�_ax�5֕4w�@�r�Ƥ93:�q���]q��!����������������n�N�wP�I����z��Խ��V�#�'&`u9 h�܆���_ �k>����ϳ�}�{������
C�����<��8�n�$:����� n^:�N���>BRҜɣ�}������{��u�f"n;�%~�5�������_���ܚ��w/�^�����^��!��+��Ͻ�����oυ>���M��`��D/P���!�>��M���|��9��G^gWr&H{���8��3�����g��s/��C�4y��y�@�ܾC��=�q�퐻�q;���]A��H�������y��=���w:��� n]A�����)��<�$)u��G�w/q��'�HJW2�_q����6y�u�u��� d����|���CR������]ʞf!B���I��!�b�>���~f�3U�`��������zH�
f�_���y�S<�������/��4��*MǺ�;��l;����(�<��C�u�W���P��w�Qт��u�+�u�Q�W��D\�G��Mv�&�9��]A����5� Q��K��=c��(7)�� �>c�_!��.@��ۈ����;���^}�����y��`=Jk�x��8�ܦ����d�H����Od=����vy�<@�s����9�����_.\��u-�	���e>��$��C��S���Mw��\�����$܅'=u׼��k�����{����i_e��.\��#�ԇY���p{���c��ܦJy��ɿ�S��������z����M�R�}�ě�r�!̾�����S����.��G��
�>���O$tq��C_b����Sodc��)�v�w����W�?R��U`��{��x���s;�:�r�t/P`�d�/��+�d}*k���7���_y���Bw��)���{��;�'P�q��\��w�?K��)ůzм�pw�H�:��x��}��׽{���{ߠ�����u�n�9��Od)��g�^��;�ۙ��l�|���U[}�Z�~�M�Mi?OUq#���Ԇ�è_`�u
rk�
C[��Oe�N�<��<���N<�r��;Ҽ���\��~��^���������JZW�O��C�0ܡ��r�$�^�;>�=��9:�7.����}���������_v��	���st��V=3�o�|�9u���D��˕���7�?�;7�z�������[�G�6�gU$�;&5z9f��m\^bD�x�~�����"""�,��j���^d�W��X���?A����b?HR�C�}�����_�a93pC��u�����k�8߾}���O-�B��:�ݹ�R�}�����@�w@z�;���7����^�s�n�~g�������'�`�Pd��y:��Gؽǲ;�� 5.��=��=�O%�){� �Oe�=�������~��g]���o��:�y���y���}���Mb�Z��rb������7(y�B��y����uַ�y���}�%�C��{��Q����by�8���u�}���Ն�My�A�Mϐ�םo�5q���~ߨ��rrG����s���>NB�Z��qO�t���5�*s�n�����l�^�ߚ��~�g�A��┟K��ԉ�����u�����X	��{)䦤����>���=�(=�u��㯻�{�}����9�=��B��JM��~hr��:\� 8���
O%u}����:��|���M����ՙ����U񿾥u��u[W��]�
S��>˹w+�u�^w֗!}�7��u!�b'�|vu��~���ƾ���{ߢw#�u�:���;��<��qC���;���O$=�ۘ{� �p��T�,��5����m����(�T־w��ؤ�v^���Q#�j�
�qؖT�9�e�)D�'��y*N<��E�h��!Q��(��ē�,g��	g{��_���� 8�=���w�GR��9�ة�;��^CxP{)ԏry'~`j�w/�=aܾK��;�8�8��{��>��]����#��b�k�:��1�@������qO$(�G�7'_a��y����#�<�ی�Y�<����=C�|�r�+ŝ��N� q��
 ���a{8�܅!��N��_ ��=��{�~q�t]�~>�|�����=���N�}�����~�0���%'Q�=`�A���=�`�v����$=��>�q��oϷ�����S����=�<���G���Wr��{�5��`ҝI��<�rf+ԞO]�Ѩ�|}�}�����<����Jq���/�Pu�
f���G�y��.��z����;�5洦@�7@�z��<���߷���C�1]������7/���)����!����b���98�C��P�{�Z>��]�s�|���޽S ~:Ť(|��=��tk7:��%ws�ܿJq�>��w':�L�`w������w���]���j:����'Wko}q��^v�CI����i�;������ysu��߯Z<���I���~�dh�lE� k�:�9��Z��Υ[sV���M\���[-��VV⛪��ܾ���͍̆�N�5���R���W�������������Ĝ������u&G-�}�l���53_�4y�}N�8�i�auz�,h ����{�ON[��ӹ�:1Fdvᮆvm�����]��+ч_�;��Wܒ=����3ޝ|G������~1��A��M_��E:�cP�w��a��6j��^54�����F-��4�O_��A�^����9}c���gt�rOM:8*���K*x�8��#[��������m%S��s�Ŋ��t�d�7:H��c�*�"Qn�|�}�5���_���j��m$�õ����'�^y����.��&����;������2�*�a�pa]{���xI�o�Ԝ�#J!B@@� �P	@�%"P�%IIKAILEE���:߾�o��^���
��yA��|k%�d͢��&�	�1]ƾ'��9�ފ�V�{^W�,2�#]���t+��y�%�����e]mx륾�5�do�_G4�Ԃ5��\nBNM�E�.�Ν�����g|<�����+}������M�Y�� �]����K���^oxL����U�^���t����ċ���ګ:����|E+����Qo�|�]����>��ds�&+�l����z�x�K��ܡG"ڜ�&�m��o�B�k��fE���jz�fw�R�u��r@��c����7���+���.4+;�Z[�Pt�<��@���e��/��nZ�]-��k���j�6N�zb����;l���t@�r�e�.�T.���W�"��
���O�J�Bz�e����� `*U@�f� �HL6���<7� �:HM��7rp��W.�v�0�U�y�H���lz�a�䇌�u�<��k!���[�w���%^tټ�n�|�`k�G�ܖ�\5��ۙ��"Ͳ�/��U'P�wkzJ:��5�i�È��\N�cK�(m���kP�����8)�7�M�e���M4�8;��o�8n��b[���A�!�°�V��^h��r���V�x��[][
<^��Iuw�������9ەv���
!o�Av��3�q����%{O<��w.��*�7%Kx��3S�{��K�K�Ŭ���1>�n�L�6�Y=���ѡ	����O�]O��p                     
gp�|����:��������Ł���ܢ�����Q��s��Z0d�/����
��̽�C��F�����@��[��.�@\�@��Ң3Mȯ4�K'8��Ɇ[U�porj3Op�z�6d���im���gf���+����l�eg�z={�����)�j�7M�w�g&r�i��e��Ȓ�a����m�̛�J�-�u�b�%:��t�m�9O�\���+N�D��b;T)n"sK	_�����7��nh�C����ڲ[U���䒨~�0EL��l�.Sj�]�S-�1�X�Ń��+���R��BeJ;|�wJ��E�)'v�j�R�Ӛ/�Դ+@�����K�3��B�'L�ntU�9��^c���^�����4�v�ߛ���7���ï���}'��?�h{�!H��@�j����j���/�)J30u.Z�r�(�*���A��,���%8���$hiˈy��hx�r%Խ�aHw+�j (L���Y-9B�Ak�V*H��2)��NI@q&C�0kX��Y(D�Д������(]J�oԔ�!%u#��0��`q��dQ@[��j��R$K��"\��o�}����ծMJ�Mpᣳpa�(ڥ��hV',�Y�z	����#�F%;E_}��GֳƠ�M�0����c<��~�o/�
~^�{����,���^��z/���<��u�;�>�T���O�Pr��xo�foiɺ�����i����Bj�bq��o�5���ms}F]� ���זmz
��l_/!�sڨ� ��5��,�K[�k<��︯�/�j�>:�~���qy&h�|����������^�'%��++e���l�Q�x�z��_v��y��]e������dOBX�'l����T���\�^�ew���Py�5���ɂ�g������V��ĩm{��4�r][C�7K+���׉�C<�~_�H�7����X��'Z�Wl$'}`�{�s��GB��}��ċ�}����}j�M����7s��z�˩���}��{��0�&�[q�Q���>�������H�j����&�8��z
;�W����n1	���p`z0*�t�Z��-�n��e�?*���y4��3{c�c�3��$+��\�-�U�#W�Ǻ*�\>��1U�[Mnk���������2t+W��V�m�~3g�L1(��yJs��%=�J^��~��^́obO�A*�i���o�sO�oދ=��r��������j�|o[�(��b~����Oapu���	��� ��L�I���:2w6������s!&��+oi=��t��wz�:�%J��Q���h��8����UUU�T���WtR^��v�W1G����j+��%�'�S����q�����O����g�/5�h$Q�����'nT�M���"�L�L����L�CM�F�.��H�w�se�ִ�o�����ϽPRj��D׷�!�@���*̼���1����sH͋��2)Ļ^�����~��)إ�̮�/q��Y�q��i��v~���oFò���)�_�@��L�w\��^���G�����{����㼲r���{>�Ϫ��~���뫕�X�+6X�)e�b�v�KgN�܍���67/v�r�UӓcR�P���e�w]��z����!� {�Wq1ۗ8�e�,jz{����꯰8�s�����HQswژ^�Y[��N(�+)�хx�͗�D7�ܝ�孅��rv��S�=������n�<θ�s{���+̉%L;ß�F���HZ4��9C�<縱��4y��Ӛ��)V��퉌,��ҹ�����L�ߘ�l��oAܦ�3{�*[��w�-��g�rN~	9�Y����X*�H�kٽ�sǼ����L� ��!�r�B�+>�w�d�Q�'��[�*ڀ2z峥R��᩶zn2�v�S�����ʫֳӝ�c�ns�53�+R�z�;C�1o-Y�r�N��lݲ���ک]Z���A�ޫ#/\Z�R���;�#��g�ۺ��)�[7��U vY9���n��Ou�꯾�缾���{�?�䭇��Ɓ[��b�4��7�5t��9&��
�s{~ϧ��k�{k�y��+�iɕ��7o��z�.�y����2�our9,3��O�ï�z%[�H
�櫪�-U{��{�__o������C<�2��?^dV�y�g0!2�*�
^iU��%�N�������F��~����T1.S+�/{+���E&��л��k���"���r�P�Zl��֮I{���u��^���},U��]�'=�:4��iC�'yvG��eB�(���=���uW�Z��U���_C-��K39�Ō����ޭ��Qrkn�٦��q�>�*�WU� ���Da;x���N�t��b��q��-;�J�:(����}�׵k@-d;���{�W��Q�R)�y���=�O~���^~���To%�͉���J�	N���lcW�ʏ̸�����2��>q�.����@ų��fObW]���©8 �^�ʝ�C��_�e��l hT��f�����5�U����m鮤=BJ/9=�{H���tw#�͎suD�>�2�ĕ�_��]���]7y\�v��h ���MS��^�x�|�u]$��v�Z���}��Lꭡ�*�P�}�j���as�]"���2cP��jJ��Ҝ13}�R���5w��6��k�~�O,��gu�%_�Իn>�WN+F�s���+`�����r?������a�9���3П5rfOwTj������;�=�������A�FN}�\J<�4��ډH�I~����ط�n��5W-��z���[��\M��F�q����8�o}�6n�����i���z'�n���w~R����q���9��e����4��+����� �ir���R�EZ�pƻ�Z��^�,���sԟD�E�"ҥq[_Ok���ey�|6�궟��<��r������?8�N�:+w�i�\�Q��<�������'nd<T�O���B.�*MN}��Q,��@d���:�ɬ��	��
:��iȪA
:�OV�Y֑�r�f1��!v�*�뱡�:�9��A��������X�l�����W�
b�^��k>j��b����Ҝ��S��;X��{��iQ/�e�ſ=��ۼ�%I�>L?����\rی�W΢|�:�����<����U��\�_�Y7�=�*۴a�����L�(Q�����&�F��TR��8g^�}zt�
���ryX�bV��r`�38�ܛz}}=�F*-H���v߹Oo�d;�g4�Ǐ��og�Vɹ�4<��_^��v֦�&��;:�5�Gzc��5���}N�]m�A�����iڮ)*���.��"��w���T��7OA�k)�
��Ȥ�dfZJ�*w�T�bm�Sr#Bֹg�%�CB"��V��z�BKY��4��9{�N�����c����}���=ῃ]}��������xG�.7�cծ�eh�Z����	�Ǵ����l�rK�^�����}�����
�O�eMCü��&�������w�±ݏ�_�ׂ��S.aW#�"��˛©������Nѝ���D0��[�_-���F�W�é�<��a���ZF���bջ�]dy׺i%�r�n�=��D��}���3:��;=��3�%��5���v��y�a|(�������*�w:>�VeiU���,�w�~�����!�ÝL���Oe{VH|�9�(2�]n���v���$I8k�G��c���)_V���!�3�SrE�}��@��g;#�H�����}_u�{ެ_���Xj����1]�������rf��5��}�wW\�Uǀ��u�gԚ^i�s}<�y�'5�Yʶ*�OKHe_������~���V�<w�l��e~.˳��{�J�ur��O8��}�ՑY=��h�X�׍-�2�}<��ly�^��/?V@���U�s�g6B�5Qz�S��[�\{|T3%N�]�g0J뎹��~��~�����w�:��z�-k�8*2��\�P�������؊���p�ܼ�}Az�WA*{E<[{�F��_��^�bky�Mܧ12�S��O�#Q�T�J�suݐޓx����a�����FL�5��Ʊgh�
�Df�wh�.�=�Wn��*;+.���o%L��v2��;I�f\d������RR���k6�p�17L�4��H�IDZ�YS�y��i�ThγM1�9�Yun_f�γ��tNn����K@��ӗ*)�
5:�+\a+;t.�t�t9M���T��Kw�^��Ǻ�ám<�@Ψ�W��ź��äM������u`������V�J�{����W�IcG���� �sa*�x��S�ٹ/�5�0Z�����A��M�L�S��ɚ��P�%��#�aV��S���W��5��N�r2�DW�Jݶ曝��N��8��`�^v������)�J�0�,���F���pg�{��u��J���1�`|�}���ȯ��n�����l���厽����                    I\V�]���5>ܒ^V<��Uď|�*w�w@t�@R�Xre�b��%G�{wכ�+��<яJWK����\�������B��s.i��nmÐ���2�Fk1�;���Ӯ�Nw��-w(=˝�Z�����IAk����vs8V�RA$�>�s{�u�[l�F�+	�7�fIٹ�k��Mn2���8;G+�J���X]���Jxά�9u2b2ͱS�V����f��ƻ�Z�շAkW�\�t4qs4��o0t<��cڛ�W:�X�ѡL�a��2�J�����Ȗ	[��Nm��0v�F&�CyQ���<����a���1�bH�zA�S�S��o6���P��,Ktx)������c*�+:�	٩��n�<���S�k]uE��ґ��՜.HC��3gb`���!2Q�'�� �9Sj�
("��-:�R}��5.�8�Z�tFJe��V	�k*��Z�
dgPjiu!I�ԙd�b�<E��Z�u��7����L��:�G%�rG,��M\K��d�	��@d�^#�P�q-<w�%4�8� ְN��52��qujթ����Ĭ�#�$�KU��2GD���kF���9�d�YfU���`dg�5h��i���P�wv+f�$��-'��UԖ��u=�j�/1g�Xu�ފ�=�{ڣ�Q�}D٫��g{�'���r.���t$vy��w��W}�SW}��<k¾w��83kޅꇞ��'��u����>�z��h��&�A�snB_7����w)U�3Ԫ3Xfj�}�p���M��&3��qEF��O�U�8�[3��eC�{����rw��A1�*����!-��w5�0�X���W��_rŽKyf
��C� �Gs��}F�Z��I`��q�a�m����sh�:�cE�c��D��*�p�9:<���i�`�w����+c�֟��a^;���ż��dj�J�����������nQ:&�n���sy�JiSڻ�V�ޮ�ϟ4չ�
Of�O]v*bK�Ɣm�G�UW�Vb�z~��0_��40���uK61�\W����r�m�T9��(Q�H�����nz��#�+���:�5h壏�|�K�~�:�����~/�(�$�t*��˭FkP�ݾ� �ʳCS�G�[J��l��Cq,��2�&^�ޤ�o<�ꭀ�&��{J�t[��n}{5��v��ʚ�=̕�O��T]vbX�ө�Ԓl\�Y�W6�`Q޵�Q~q��=9	�淆.�q�w��o���e<���^�g��.8�U����ޭ��e�W���/f��֤�Ǳ)���MWn��r��	����[{�����L�I"�%yw�(�����ɶP�����>z���G�<�9����}������K�����*�5,��|����\�[� *!>�#��+o�5���VAQ���Ú_��^,��T�w�]����VF�nww�9kk{����ӽ�\R�}G��|Nm��2g�],:�%�QWX-=�}��~�/��^V�o��93�j�'��=2UĮw���uǠ�ALɸ�J&�g-����#W����Wj�*��X���t>�o�����jy�v�i�,fTc<�ۖf?o7�$�/��V&5<[zs���j�+>�#�W�r�W��m�������0�W7��ˎ�76��_�]�ȵ!���)���������+��_k/�ݧzt�!��ю�u:��_}_V�䞛��x�ٔZ�{-��ѡd����l�iܻG������Պљ�k�y2�ӗ��Â�f�����TQ+A���r���f�]�+�q��B$��t��j�>)�3��}�жZ�"�c��f���' z�?K�T&yz��Q���]V�����z4x�q����Sd{ʜ��p�=Vߴ��1�[��ͷ�����~�iZ۷:���fx�Ժz�~D�i�m�`C��b{�얤{��S�^�:\@ ���6%���V��E:�ZW�4���E/M%Zt�P�[Bk��a��S�%]^������v�ǋ��b)�;m`��Ɉl��T�ݫ^�1I�Y�e��.;;�����}�D]ع6���ɋ���X<<�7���E�{V�z��-�w���(VP�4���5(y�Gp���KG;��%��M����%��:�� g�F*�j#Nҳ�n6O{ЫdQ�#��*�){(a��];�@���ha�al����vw{���>3�㮚����ʯ���\$G�����Ǚ��y�H��*���e8l5�4�k�8է;s��&a��o��*P�|a��
���<0?Z��+m�^·��Z�h�t���wZ�V�t"���UD�T)����־HV����ŀ{��z�hu����F����
��AX*�Y�8��;7t� 4���j�/z����S<����,�4R�b���WV���4f[���J<b�n+4z��P�f��u��۔���#���)zD�CRV\���9��x+#&̵ħs:�;��=�a̖���ga�CJ�շT;��]������)���W1F���WJ4��|Eڡ�&�� 
�^�~��b:)7�轘�L�*==� �@+wuj���h���Y��`Lɫz?y�&A��-�� ��,T��-*�|O��;uZ�0�-�\�=��z������`B�^#��GG�U�y��5w{�ᕠqV~�§�%\8p���F�X�X��N^��빋�\���ĺn�*�&]t�Թ�MaKO��{*Gs4��!>	r��<i�5 ��5h^: ̤�h/e�n��g�~Uh�vb��ݟ]�Vte��saљ��=1�z��xW��ӭ�KK������*!]r׷Ć�Q�����b��J�8h����4]iӕ%�
�
|1w[�M��f����I#�v��e��Q�I�3�/g*���:&[�^ܵI�Z��K�a1�?z,���ׅ߮��6֦��lSc�(
�mwCލ��	��C[d�NXݫ�N5ì��A���|mԹ3پ�r {��:������̧�K���#��9�u���ZtO=\����ǅz���(\�(;d��꾯X6MA�a��MV&� ��X83��[\M3�Z���v�"k!�OQ @�� Vq#����2�_e>�4l�zzVuØ�P��j�S `�F��`�~�9m�]��A���<��Y�em��:��vPлF�7��^g�(��*�N�=���gxc�7N��pS�a�Ry\zq����d~��XU�dB���׍Z�?=���C};��]d�D+��e���(��p�y�>�K�����F�8�8'p���f��p;�%�&}���ֻ�ь�gM��ɨKŷ؛�!Yy�-�����&sS���ٗif�ǅ-J����q��	�\І�'�y{��*Ǵ�R�ƈ�tu��`�K��\4�xZ�9ڒ�K��t��=ǆ�:o'O"0�̥��­����s\T����Eg��m`"i�G@�_<5��.��7�]��U�Yh�H��y-6�\�O����cZ2b���h��;9��������>&�K���M:�k��x�N�
���em���식���rz��)��0�xч�wʼ �٥U���փ��w|������V0��\�*x�S����Tsg���o�^Xaʗ�+�`<���]�)>�߱��ש�-�zaVX��2��a^��AW�θ
����h�b�0��6�&�.zkn�<��T�`�{y��|��Ws�t��x��9G;.Zx����Y�1�ma��/`عTG�1Rα9I�zj��������C/#�����$�w��
��%���X�\����wN�����b���0VPX�p	}HP��]ϙ�Uj�e���V1�罻�����@���֊�h
L���_^�^9ǀ��Le�2+'����fe�V]���76 �4?�G���,^^�����bB��|)Vj�X�x�'G$�eկ��ڨY�8T)s=��ٰ:�=sW0�]²������[C�}|�n#7��Ϲ3�zT����\C�:����S1yS1��//gWk�����pV���qe?�@^r���:�&��_o{��}@�~3M����"�B�ܪл����/�G�s��o��e�8-��|��ևe	Vlp�V�w�=�
�6<q��#7�Jܼ��M��u��.�3.�k#vk��gF��Y|��]�����l��8`o�1{q[Uݯu%��A��DՔ�u�T�g	��si%��W��l��Q��kk�|5����9�i��Pł�0:����l��~��Ѿ��X+��E��n:��I���<�]K��#�h]�7�����������P{㡘����]j�|���9�M�1�C�s3WZWVo��x��/�X+O��^�-{��}�0`���Ѫ��h.�xl.�꧱��x_�UT��2�s=�ʯ��  �M�|��IV
��X>\u�ͮ��g��3�h�N���� �C�߀w���ғ��s>�-Or��WMs5�˒��u��>�Z�
� Axpѭ�kē����X�&�\gM���lԗJy�������G�/`����z�}Ί/�S"����WD��#�֎�Z5}_F��ˈ��#�nV��俬i=X�଑jN��nd����'���I� �UͻU��Wd�i��mq��9��?wr\��N��U��W*.���j���[a9��32�ۥv����$y�I�
��R���+���ܸ�T�-�3�W-V=\9�y7E��WU�9uwLJqw�B\>�T�dy�m��u"%�%�]��q�6���(����\3��\�o�I�D	cyY}�ݟ�8U����6K��]��6q=C���(�]�6����r�<b����M���T��Kx�e܍���+��R���X���jmvUь�����M�>FAaS��(n�>�f�|�X�j�dg]��л�ɶ;wR��ߗ���Q8���w�{0V���75�Î]Kޤ�:�ۋOA�@��eVj�if��hs��e��t�7V��)LB�f��NǙG7w'=�ȧokGk���z�S�r����@           �  `     I$�5	�ń>23��b�P���J�g%};&Tz�6⾔6t}��Y��kP�:�7e���E�!m��WY�"]���8R��bQ/�]OVSY�l�Eu�����uR6�H��e%��g��k�g*�Q�*��J�C6��fޘڼ�*��v��ܸ�V�Z�8�ke���Rܢ+&���uX"�)~�j_�
 �K�T�{�1�b�1�a����e�=[�e:$�w���	���u�v!����%xmNӲ� ,�tWc���Tꄡ+:��-��.������ѩ���\�
�s���t�{�w�Jh�p�ɽ�pX�8�!����"0t��כ�O"�dw�.��wS�mud�v�t�W'�|�h8eZ�0��� �e��:ἴ���n�Ε�����\����&�e?DAI\E&�Q4��Y�.fa9.C@e�PqkYKVa[�B�p��Y���d�e�YYK0ᘕ��VY�:����fa�4�K�!�5�VbP�&k2�n��5<YQUMQ��SŖC�ݩՓIE�:�Ð��ITٙFFe�Tك��XA�dVC�NNG�PPPDS�A��gRs&���
b������*&���uQܙ/�NT�5@Q2u95T�����qu��RH���ґ�X�%�cq���v��:.7��W	T��5_ K6�6Ĳx��*���}��H ��&i����,T�M�mQ$˦��8n�s{{�6z�_�"�HA���hM�\�\�IZh�@��>*;��uD �8�5�u�}�yS��p(�h�P�+A���@Mz�0��4�ӝ:�u�	Vmz���q1�JaX�wdm�el���*�g 5ѡ�ʽ�󫰫]j�.���pX��ߠ7^�fK��|*/-ј�L{��'�+�ݚ����g'[��i��]ˀK�b�w�K���Ve#2�^y/�����{�隣/И��U����n@�2�pz|����{���;^}������+dU�u�^�v��w)f㻸�;5�ۊk��	�RHz��^z��f ��5ܒ����?V�`P�t����r{}�:�Uh�}�7���ͨ�ͭ6D�e���{V4�fI��ɽo����Ԑ���N;{[�����,�xt�[4���ͱ6��ٌ�[�������1�\e)�-߲���wuu�;��78��n'$�44�#�V/
U���g��8���6��~j��&?I*�eУ~���.X��&���U����h�	�y{J�y������d��\+��o��4g��1�Q.j_{"���z�z�y�J�>^��jƪhCJ�x�[{��v�{�
���bU�#$���2���p��{(�����cO7�eM*�}nz|��- r�N�dFٔ�e�4�>����fff��p��f�(L^)ʗ4����j�_mm�KO�|i�[�������_���<�?��@j<6�X��@ܶ[��{�I�G�����mӯ�֋�%M�J�<:ϖW�;��Jϡ�z��[GE���6��De��ޛ�3f����ͩ2�Tr�����>�$�M,���r�8��t�4�ju�>�Cp<�,h�/�?�Gu�w{Ԝ����r�<`9j��n�\�9��E>�n�^`�qNc�;<)��>�$E�ps�¦��e9׉3�0�뀦e�:ίD�Iv{��S銙U]�P��z���$�/zݢ�
�v�W(��:
X�Խ��)\�Lg���w1Hi�P�Wr�}�ܓ�\�nzU�E�]'�|��C��<`�uq�N���\Z7G͊8��(cG���k�0^S�/>!�F���5³�I��t+�u���3��1w0��&��\4�UL��*���P��b�+/�Rt]y�/ۛ��t��g���|)Vj�D
�	#G�|�g=r֓�r"I�G�����Y�<;��U�sR�9�w���\� �:�t�Ǜ����O{Y�.��Ӫ�{�	�Q�ٹC�XE���ۅ�\�Ge�S>
���IJVf��+qD[��N+[6&~��1�K��(�X��*%y�����F��`
�#��y�;}��R4�<�S�㎢gQqW��}0Lҹ�Fu_Wf�Oy��C��b:����q���n��]C{�^���cڅs��ޭl�>�^m�m���G�yխ� ���Y}fDc��$1E���Q�,��J�ףgj���&=F{��W=>��۩�^���n͔�R��,p��r�ۗ��1ר������6�0���g�{/��K�pV���n	z����c�^�~{|�����.�]>Ww��P@�z׼��S���;��*�2��.c�qGȅ��C>\=�g����_�V��z��n�=��m�D@�{��U3�����)]*���W_J-Zv%�Ϙ�LM�*ih�rK�Җ�{t�ʁU�䋱�9\��P�+O�5ђ�<hX3u(� �^��ɤ�C;e���2Bf2_�����S�瘭�^
`7 �`;��qvxT�ӓ��7��g��߽o�~��g��@��ӺWN����9YMlZX��_�$�{�x��|,xxx`@����;����:�p���o��z�h��^Vh����u���4S��;���g�B��L��lU`�$Q)Uݡ�
g�j[��.	�荿��������]h��Y��'�Щ����Nj$�4�Ot�i���n����#����,��pVp�g�������"R�'�1{R	��W֦-�Ӭ�)Νp̺ʅ
�k�E�p蚻�ƋL��&&|�nM4��@*֫C�0c�����*�;�6�+�o.^{�i�}�8%
�yժՉ���W
��X��`P��^�,>G3����j?J����[�e�k�@(��
��7n�� ���u��6���K�%��u&�^�/��벯p.*�	����<f�b%[�u�3?�C��I�K�UC�]�d�4ib�����/�3!b_�i�E!���~����=�<�c�˂z�:;��Y�Cl�ݝz��)��������V|�8����Z ^�Z)�"n=��]���E�s%T�V�{�}��Q� %ݸ	��3-\��/��̎<�u�po���������V �m�g���$ߤ���Z�V�c��C���z�2�^_��دv���Ƞq�{�ɿJ����4�C�k�/Y�iۢ�R�Z:�R���{������\��\
�f��Z>��R��Fx�j�\=���0R��=&�b�I�0]��T&z� Ⴀ�hCP!v���'w{����
���X�f4I�t}����t˂Yg����]��qID��L���5�w�0����X��S)U�)r9&�]|�{j�f�I��9�4���t�0�Iξ�V��'ƦsWX\V��v�F(��|�~������mX�H,��P���(2�.�*������༔�7��
�Lz�e�,��r�#�M@Qx�F0�,�z3^/9���l����_ȼ�X˜+|+�I<�x%��ܶ���B�}�]��ߞqtX(;ә]�n��S�Yn��D�8�^�fY!�N��C	��`٨�p�gGZ���ӑi�6k�D�#�����+�Ϳ��E�0Е�Bx�TԔ�Ú�ɾ��lV��5V�Žj����V<�u�����W�2���^����D+��O1[�8�o���p;�4�te9�/h+����z�Zh;g�Lt�����mW��l�V;sⷫ�p��秽��|3@t:�Dk���s:�*>Y'p��
.-}��~re�@��Ph��C�c��4T��@(�kjW>z�ڻ �7�,�]����N�雷ǔDWuc��,�I���s!=�=}�tji�^VNWfq<��A�R{ޣ@��e@�xB����K�W:5��
Pϑ�/%Q܍u�`��ݻ�3�t;�Q758ˏo�� j�ؗ8�g�6��΁�$��v`�
5>�-���byK�;�����$�dz=�9�v�绺��Sθswb�aD�gZ��$�������-����9Aۙ���;e��UW��b&T�!E�2�&zx�Ӥ����\�ֈ��=M���sʀU��ߗ���1��ݯzf�� �㢐�6�����Z�:٪٧�ʂ��'^:!Ny��߼5UԾg=e�/��E��S����kd��d�yd��uϞ*��{A���>�w�ӫ6O���
�6nS�s��s�����vpsԄv�.Žj��[����~%��AjI4�njr]$n��H#qM7�g��갹SpB������.��#S�P=�����喤��ِY7��˾ZM�R�]�ٺ�NA�*����74���6�W
�)o�	g��^-�=�����_^,M�^�i[굌�\*}�T� Cz��}�}�q���3�?YFg<�Uد,�"Ǉ����Қ�T�h,W���~�S��#���oo$v�W�*���tHCM�|��k{��-���j�y�|�e/ny
���X��! !�N�񣃼tw�\\�:�o��
`a�p��~T��j6����)�Q �6��[��>mD�++`+��+O�A����:9�.)
�w%D�{�`�l�e"9X�Uh���^��
q���'|Gx�����-���]L�
���f��F������hq^�'��N)��jdL�oT��+�R��b�4X���n:��j�M]�G�G>pj����G��z�
:��Νf <g�J��X����R�8�M7%�O���
��$Ȍ��0J��t͔�a���E����/O����4�a�+5��K;�<�ȫ��[�^�^��H�r?A���;K�Y.��k���^�l٧�Y~N��&	�������h����Po�1�@�j�m1ֶ�]��M�2�`�E��;E�N�y�O��Sǝ�Չ���up�\��x��Lrl6����C@v@��b�w���,u�ZfB=w��|Ofoucx��n j, ���;Vݏ�=���ht-�8S�#�A]j=�������@ÃQ�ִj9~g��ޚ��\��ڭ�XB`�P����h���>�I��S���{={U9p�g�lX8:��uW���o�c�6<�]�f�m������~��G�JR��szɹr�}>���1��>��U������1��n��%���b��t��.��3���l��"*E�m73R�]�X7�__'�@�D��W1���wI��W6tѳѴJ�w�4ʻ�Xy�m֋���X��e���+p;N&�i@�N���^�ש�Z�k����,�&��V\m ��� ��tK��M��Y�h��3n۝��Ü�=��Ք!7�F. m��}����f����4��&ܫ�1�:������"u����Z�:�E�j]��6�]�ݧ8��'ZBK��ssU�V�i��G1��Qv"����8�D�"�1���P$�)��Eغ˵NK�K+��u��x;�,MÈ>ʜ�C4t��\+�
f�g�������a�7�j�Uj��%��#��L�/,㚺b밖L|u+y�w���Sfw0�LրP�Wu�����d]���s�קk[ӝvZ��Hk��Ў���4                      �޳�22�Fq�k���"f�\֯۾�M�,�uNڔz*ќ���(.��CwW�@j�'i�k)rƎ�F�YW4L=t+�R�)]~���r�k�|�:�2�\~���31T�Q#2䌻�-fm�b��\��lt���p�`�H�5WM�E�`6˭,}�\}J�h���c���˲	utC2���gG0c��DM>��	�|1�;�4�����fـ�2�؝׷%��'Y�0���Ƙ݂`�[�ɣ��*_q3&��U���:��Y.��$�`���[]Z`�ð1�F%�[{�8�,�R`�2+E؆����í0i�;f��ӛ��k �vVی�n���:��!���@�zj�A)��p�{�`����7��4����C��4�9K坮�;i�� 	  �Q1111?D���R�IHEAUIDE��wIBya%-I�pmg�dQ�5KGGP�KG��E$���cΌ
i��N�2H��gbT�DLEUD��d�TID�.YEV�
�"*�%�f*����2(s���c	s ��&����2�j"j��`�d:���XSLETE9DQU�5SF$DI�<�S133�g��@g�ӗS:�ی5)�l��L�&��,uBU;7t�*�������g�m�ڜ*����y�VT��W������a�")߭`d)�}��_�_Ld����UT�vL)���9J�_��x���Y��3�OI��L`�5����Vr#C<�)?�Ⴌj7����6+w�I�Apy�Z�+|.�^R��v�(���~y���W�������g{�"ǨW�� �"�Ѵ8^�9"��ʅ�t[��(s3=(}��� �~�I��Uų\(J���9R��h@���3�8(�
k�ݽ�]@�����˅�C�U<]
9��p���ى�d��W1c�phuq�T�_5�u�b�>��/%Mn����y��,�x��3-pt8A'������Z�g��z�\�y?-�>p��"��Y���5�����D[.�*����ɽ��@�jy )on��p��Pt�@��k��[M}Ѧs
��TNk-abv3N!��0�v����7&3æ%�g�:��]��Sn��`0�'����%��`�^�Z�o�T�����s�e���"n��Jjcos3;���%¼��_<^�~u�r���g!�AI̩u�����;=?d�.��k�j�Q/v�%c�$�Wþ��c�vŢq$����+��=`�gQ�|�N���������OL��J�@P�V��(;��&9��*��K�=� 헆�=G=�^o�H f�'��*�]��^��g�z\OO��c2U��;�Tnu��,u�U�p;�x������7���e?��&�ML(�B#�HT��x֣�y����qϛ���x|��9��
@�C� 5��#����s���T8S�Z�D�F�.��k�J�<]O*V�����wv[����f,Ůce��OvV�?\�wO-�v�\��D7�}$�Nr��'&�����ھ�!L�c����V��sƃ2� �c�`�LC��8�O��P�T���l]���Y��)�:��С�Ɗ�:�1a��k�Z��\Q�n��S� �Y�v_U3u$�yRT<�7�r�xu:�O���S�8/g��q�L����s��ףѵ�N|� ����ؔ\e�M�jI�R��vzby��r��E��Z����r�kPV��{��w7��ʂ5R�z%�}aѣ7�@����\"U<�C�m[���E���U�V�&�R��T� �8b���'ȷ:�56ִӃc�����jgj�Y��q��kv�����\;��s�^{L���)^�=��U�v����n�����J��sđ�s��OMoNx|(��c[�Z3�_*Z�a��=#�ة�޼0H�*�K�j{6����U��|+w��@Q����η�5+.�8�f�|z`٨�ML?Qo���mw�� R{�V�]��L�	.8�H�E%�0�`�ˣ�J��Z3������]�O��X�dWM��q����"������p��*����1p�y�p���X�GG:�Æ����'��{�
l����m�a����WʼxU�	h~(u�������>vP���w�J�v��3E��&!⡡�W��L��|�.���l{�����p{�LV�N���+F{D�7J���UQ1/n6mә�L��n������T�\��:nN��93.I<�O���9����;�M��r��
W�Q��Ƥ}�z����A`�e��LvjV�Z�2�ݾ�o�}'�/��s�n2�S1���]Q?y�pr�,��0;M��N�t({��J���]�LN xBr���Z'� >�7�FC�ˣ����ؓY��]J[�nc+oӀƠa�c�ypz|��f�,�u��eq��
��b��"��ճI~@J\���TX[$�w�"Y�yO���O#�S���2�~��^b�OE�п���fffΝ֞j|�Կ}��z{ѫ�i
�=�B��]�Y�W�e��g-8�&�\�����ת�A�/yuWX��R�[��.���VRs�ٶ�c=��w;>�}>���$Y}2��[[WF�d���:�Zg�lfO@)�`P��X�a����G��VV�>�N_���iw_K�w��DL�.��u71���үO�s��&�������R3RfvP�qsq�����U3�Y0��0Oy�����*y����u}�m1E���x�yW"�Dh|)��XxޮV�"��y7�Ez��D;4> V�0���#$���bՃ��zf�$�M����]�`�����<4m���ݗYP�}6�m�MeT��Z�B�z�[,p�gAr�#�M@R��ՙ)�5��N5&/vZ�;`�!�Ǚc[V.�����+�3�$���`[��"�
�)=2��L�K�ݵ�\܌�n8z@��YRԏY�wꯄ���{�6���#��d�_b�>Jo��]
O.��ϣeOVn���~�@���Ä���С�+v�V��zrj�\���k|:����;W/����+փ�c~9CKk�3N�j�������~�N�yu��O��5;�V�H�XYW�rh'�����ZB]z��ஏ��[�z*����ʹ}������騾s�7J��p���W�Wsf|�0�U{kʣTT��gcG6
�%Ӹ���LK R8����Tv\����
7�f{B�dD����������%�j:OR�W�u ��
��w�������^�Q��) -'�ͫvEu�ySE/v-�i&�EOAK��~�&е�-h��{+��F� �����;�z�˹g���Bhs��hΐE�����{(a7xgw����Y��KpՌ���Mf�Dc�"�m�W\�kr}I3�3p��U<y/���@g�.����_*�S���1\�.�(���Mbϭ/4����׶I1�^ua�W0�I:��pL���Y�q�m���{��WS�|�ƚ�D�?=4K��H�hp�*��s���A@!�@��9��8_�p5��?�yPyQ9����}���<+@5�5p)�x����E_�n��fGy#��͊�T>.f�yҪ��d���g��^�ZЕ��lw��u��:�����q�a5��u�z k����|i��,��{7�E#�~	�,?Z��V��_J��d�+����p �<}��m�.
��u��6_��+�;V����,���;\G_�X��=�7b�kU�`�ܾ��on�/{��7F� #��S\��ܚ�ύ)��̤�Q{'u�?%K���Ʋ�y	N]�-��b��OSW�����.�-������r�$T��Ug=q�3�n~Ղ��?Y���.�V���0�ez�NR�����w�η�ؕR���7�� ] ��䆬��܏�6���׹��X��X$����wS}EV�ʗ;��Mĵ6�2'&�X5��P:>Z2���_:�m
��@V�xv���/��fz�R�Mi<����3��ާ.c��.��kw�pM0�c������ĕn�i �M_/l%�`P /�3v��X�
c}��-hT4VN��HTj:�#�>���4g{1�6E��J��wJ�W�������7Y��u]D�3}�ݚ�I>�@�U��@
��*�[�Y�f <R�]�,���w�����u��Y.�����הb���+׹A�EV�Q*ǟ��k�fO�.{,��Gm][(c�J�W*��%S�9)"<io%Iٰ����|l�Q�D���\�vo v�U�re-��UP]�/{�n��gʫ��:%YC�A�ʠU��Z�h{Y=/����;�</�&����U��R'�P����jă�A��b������lU�����ճ8����X�K�gk�U�9�kI���IS��~V�x@�`@���S��{j¯of��IY�=P+ϮM<�
��A�D
7w�+�2�n��u��L@�2��t�K��)�ڵ!���Z��!K�`mg������0���֒N�rs�I��$[ވҷ�;��Ol����	���V���q}uN�T����0����9q6��}|��u��qu<��&�n�J�<�����iۢ�W|����0�{G�g�.zT��U2��
}1?LA��Ҿ5�|��e��]3��6���s��r��ʐ�!�7o+{����vr�Ie�el�Xxˢ���n�w����{P��m'�n�x�%���U��-�N`G��w���Uw����s@/��
V�ת�����PH�L:8O�i�`�+�u��j�s:}�R�
���n��p���gG����B%m
��ʷ���]H�N��r�w�)u��8���I����c�kA�O�ց*{z]�ݳ��k���0+�~U�j�8@�~��~'>Ur{��P��mƞ�[�s"63جp�c�."9��YuD���:�raGxh�}~�&\z\u�z\�R�L��P��a<����]�t�fw��`���6�\�iI�_��]1ʞ�0���բR-� ��={���*���OW�9���_j�x��W�Ô+*\�,z�2�hp���\�L�Bwjb�L���YjGQ�OB-O����c�(�z�P�D��5���gw=|��G(U졷��JU�:�v��^)�(CKQ[�(%����4y���� u;:�5��;��
��r8v=W+n��崖���o2���9י-4;��c�>���,�Y�V͒}���v+F����k53�����즨�(vP�-("%b�)��iC{��Y�i��NB]N����ۂ���tu3h=)̢oe:��Gqڰ�/��ҳ�5�j���VsD�9������ΘjP�&��"oz�̷���k�D�X�
Sr?0C�{�B���2�<���x�����y��Z6e���F�U����/Zz�dM%4�L��X���R��!M⇻kP�8;�#ޔ�R���W����3I���Ж�]�A�{�@'w�u�Y�nZOFa���\eᒓ�8�ue��Ŋ�<h                   I$�D�ڪ'c��'t�ӸY�����'7����R��-����՜!j$Q ,�l��t�J�%*�5�kA�	s�Ly���	N!��E��+S��=��-f۾���f_l0�m�;�e%�B��Zs(��*��v��S��Pn�X�sov�N��]�������;����4R��X]N�*Qܷo_�d�&U�MpuԊ��s;�Xר���a��M���y�楊;��L�N�j���s.+�[�o�.�V>"eC��zԼx�u%鵔wu5�0ø%����tv2Z�_p��r^bߥ�}����D-2��
<�^�3�C;������{e�G+fp\BK!�x�T�%7�^Z�qn�n��u�$ݡ��6�����*��K��@ H  
����g��(���ŔqeMQMwaN0DFYP���E5�*&i̱ɤ�Zx�h�����0y�8L�0��� ��)���j(�+#<���ʊ"I
I��*"�����()�$���TU4��9c]FM%4q�Ƥ�̊b'�"*����U
 �@|�777�1*r��{�v��v�%���*�����IA^&b�E<�d]�UCV�=�R��}��݊�C�X8W��8���o�<�$h�y%�y��`�ex�j�
o�-mX���mPx*��� ����^��S�W���}Z>�Q��yHi�d�n�Pw^b���L�����;��p��U�Έ�<�n��u-T��G+r�^k3}Uʻ�6�!a�1xpvZ5�~X���MZ TW�T
^^��á>2%�!��a�����*����(�M��Ix���?q}����5�p�}�\����G��On*��R�7��x7��ZȺ�ꊔ+��ȝ#NVp5�\�T��c#���x`N3<O���3Q�I�V�5� .��
�~u���G��wt�K+ԇ]$(�v��``},�;/��#��yW�i�g��q��x�}9X�P��o��s��/��J�D[�S��,\��nĪd�7�V�N��XY�X*N]�QR5)��ͱ5;"�}�i.OF��o�������K�=�i��5����9�����* ��/%8d:=g�!�U���oZ�5%�/xw�3���(S�j.}��\M�z�Nۻ�n:X�޹��6�8h�����L����
�i�l��^�R� �8n�t��]����FɆi-u������E5��D*����\<�m�]���.�z��W��{��y��i�Asʬ�yGin� �����=�L�{���%^����ῆ�R��L��y��l�C��Fw��gL����r{�c&C�2�pT%���u���|+}��d�o^_w�P�D���V���<L^=q�4OK�$OM��["�9��\��:�#����u�o�ղ!�~�<*֐=��.����U��f�$�l3�9�1��B+�#��ۢ.%}Ȩѻ/�o)'R�5��6�Lvt>0�����+�;#"ǠVwi�x�$�1"�����Bl8��\��/b^���1҉ўj3L�Y1�����{�P���'���5���lDs�1Z0]�Jo�awש�S�z�z�*�Q�wUW�T�V�\t �Ӛ�c%��@x��Q����{�鵰��|<Dè`�A��b߭�XS�:��ޯof�U�5�6j�a��8=eqA�ʠ� O��;ޣ�UOq��Q�&���S׎��
M.O��kW�W���{�{��C��:��<7��V�x�=u�E�:&z=�l��>�M�z!;Zgj����P�baY� ,w�3EK��'�5����ǈ��"����r�6(
�Ʉ�vP�[�z엞�r��U����ֆ4n��UK5t�o��pЇ���[��[�I�|H�X%���N�;г;:�XMY���Wނ�=�Ua>)�J\A��K�'ݤP���*Yk18��K��5V���,ו�`��}C�Jb���T;P��禝t�9�e)F_\�emm]��²w���e�����X��53V#Vyzyh�
�k��*S���wpC��C��Dg�V�iW�*ً�@�0�QA]��{7� �*a�v5H-:j��@�\+C�WO�֒_/x�O�;CԂ��`��2^�e�uWx��]s@*�Dhg��*`r�SMy?]���Ơ�TІ�B0�a*Z@�4LJ��FI����s}����f'�����_"�.mH��Z���l��4Q��dn
��l��Ыų\(KZ�k>�33}K�����2��fYd���s������:9�es�Bc	�뙾��N�xea���Ds�R�~84k��xCY]�4ʻ@���F�Cݍ+B�������lxhg�`�~��T����I�]פ�K�Fz��:��ˇv���ζ�mTT�[*oi��NC/����_`z�sл��u�+?|=hr��;߮_'����eÂ�9���s�{����+w�C�82���.�#�
�o�Ꝥo5�����+�=���Vǯ�Վ�~��Rt�Õ���|�<|�y��۫[ ������ME;�Wnb�L���[JE�d�R��$ˊ�L���Su{*]������ �k�=r���gM������.2�^���sҮ�o"1���+Y�i,�T�P����}�4�<+�[�)��j�e��U���u;=*f%Luq^+_���H�Q�.f1
��4s���{<�� ��]��n�p����k��VH�\kw�b�[��byZ��O5=1�׉��m��m�c���f�*�5�h)V����oգ��qG���\��`�,�U1.��,�D���rHi�yS7��m���]F����쾬rV˅�J]��u9V�mY�[=�����Ow�|E���]�4��5��(�-��7�j=-4Ny�Bq�J};=݁��@�D`�d�:&�8l`Kʲ����ǳ��ԘtL��|���2�d��VKS�h�vvC�r���]w���p�J�ʕ�q|t�+��o��Ds��w�AԦ]�o�����/�0�͇/k%�ˈ�	���Ӝ(}qյ�3s}��C��hxT*=�}ָX���Ӕ���8b��ǲ{�9B���]{Iڦ'���+�5~|,h��80p��:]�5�l�q�z;>&�$;�
W_3S�[O���73L��l�d��S�xz�ʦO��R>Z�E�yp�j�7W���4:_���kA���x������檩����-P84*����`�07�L�oض%*�utٜ�v{d=�P#�-)eƷr����������@�
⺖Xrq7u4d��gYi;�|��k�e�Fb�Q�NT&~���=#� Y��J�x?vU^
*��×ʖ�G���K~��v�`�8��t��T^<�e����U�ղ͏kf���}��t=S*v8(T:�O���4�X|<Ws���n�������1�X��b�j:G�{M>���������6�Z���������(yѯU��/��P�X:3�Fh��6Ե��՗}��Af�}W���	^#��k��.b#� )�4`���?
[�D�R��8�� 뭺����Yp�v���)]g�3�g��rQ򧆼-"a�0sŠ�Y0�4K����^���:4y6?z����l��,��BtJ��B�_�A�fg����z`sqw.
�~�]�n�
��Q5��­��Щ��ky�wH�|�{���CIk�i7�ej��R����vھŤ9�XR����m�[r�(�֌;��-[����wm�E�Xm��T�݆�T¨LAљ����fg��LHp~�^'+j�v �r��`o�b�uM/	U;�.Q�����bMӫ��e{WO/
�[� �Y69��-��h��n}JQ5��mB�l�u�4)�F���w��~�O�E�3c=MW���ֆ0g�n��J�i�!I)���^�so��_��wh���`>83ܼ*J�ÜX8?����v�K���7�k!¬"t#F�?��4�/eIJZ��0��v{-C
8��R:�C�X�L���[wB���^S�[�1O6�$�+�1�;�~������a�b�UL�œ
~'�g��Z�{�$�g��K�0w�R5j��⇞���h���X���U❙��Ţ�80T�4��q�n�T��ZMbhyu*����e 39��Mv�Ֆ�՜ZSwm�^.wz5�y��X�iVjc9H�U*�\d<��V�(4�1���*R���f�M���6������D��(�.���%����|H:hH�hu�xnP��|�=��R���:Ȍ5�)z��s�
�kG�E�,�#���N�wn�z��p^*����Dqj��a�K4�\�A��j=��zV|,Q�@/5ᲵX�����"9֩u認u��SUr@��N���Jc�p_rTƌ'��mh�J��������Cew��\Z�+]���ғ�ͥ�8+�ǈ�+�;�ziyy�D��{��Ah��PV�*x�Tà3b��V��#n��ۢ=�q��>��/�mϦ*I�YѾ�z�T�p�kG:��8����b�'-!���ͩ{�W��K��u/32��- o���j���_���ݾ
���2����x)�,���]v��2�u�:�����@��%k�pR���`m����NChV:!����8S���8a�s�
�XnuM�fٻ�Z�7A��(��'^j�/F�����g5'�����?AB��;���yGDb���ͫ��x^>�'��zkv5�i�F�{�DgL��{	���-_��^�c*fe㽝�R�1Pg��"�q����i����9�4�پ��fS}U�$˲{cm�>���¡��v&��a�M`�$���j�EP@��gϪ�������D��Ū[Βz�UL8��l�&��S=>�H�G��ӆ��������=��ׇ!�/MU_?+����0�1���SyG��E����l8}ލ�˪�`��T��P
�_&P�u�	M�b�1`�MI>��L��1^��o����q��Q����ZUw����xU�	��?¡U��xAcp��}��W��+G��S�,e%Z���a0���I�-��,�GgN�c��G3o���|��!Q{b$��S-�c�FTiC�|r�!���cv��b���܆=���gU�q�*YGX��7b���N��T[�s�VTy�wU���y/%�5F�]��7�o^9�i��W,[�@�:�_Y��S��jI�~�'A��L�f��Ƶ��n�-�ϰ䓤X��$XЁh3a[�-�!7�]L�t�No
5�m���:�^��������G���i����˷�L+%�\�����҇hM!�u�.1�Z�o,�]�K�Ѣu6�=������1V�U�U�g	qc#9�3�F�1�([���yL���r`n
l4w�w�9hz����ס�.q3~���s�yf��[jROD�6vMq�1�0nZ�e�ь:���%�D�bf4kh[��4��c�d .x��L�����v803�]#ƀ     �I$�             �Rۯ�o`��W(�ݨn��y-�Ñ(l�fc�cP9ֺ8��N;&���4西��e�J�-D��|�.�;���J��Y��i�gmx�5�_]m�1Δ��B�b�MW��;;le�U��>zg����Tɿ8���֦�dO���9�]O/��[���eQ��߀���ʻM]��E&J2��	���iq/�S6U���Q�9�_а"!jj��1[AX2�9̆���"�&GW%�\��Au��,�0v=����s;�]1�@u;T��Տ�]�Y#���*B՝ѩj9���+� ���ҋ(��T�ś�'Z�|�h�`��NS�䆎�_=S�p��]uYr�.�����`�{{ȑA�#n��u_z�PRꤐ� �����������AT�F�*�����I�%5Tk���V�*��ʩ��-Y]�\w�xʟs*���Z�DI�QQSDD�QEI�����`�8���SUPADPV���jfbj"��""(��	����#x�F� �0�Ս4F`aݕ[�ț�232Z������&`�*
&�(J�����(��{�}�!��b�e���^ ��uu��A}�ݤh4].�Z��/��	.���<y�E=�L�
�3<G�Q�\6΀��φ)����{�4`�i�n/���5o�k�l�kw�8�ɠ�/�]L�t�#�N"��]�v?)��������R�J%���Wl�i��Ts�nK�X=�*v:�x^�����7� /��B��d��V�/��1�3ՉX+�?vJ��om.��k
3*�j�Ϣ���A����P���-���%��_�3)�-`'���=%1��RU�����1R�g��s�����s�A�7����#���Z8:Q�GAh��ۭ���0!��NpiWr�}þ�¯�,�f�r�Z�h� h�5��y@i�@�n����xG(q�yU�À���*�\�d��@S�`ƪ`�W��F���$�77�QV{�B�T�NM���<pQ�3�WS)�P�:�r�*��DT���t�0�B��3�]_N�,�WL�ne[��SW�G�n{���p���U���N��N���r����'�@iD)!��$�=�@x*:��J�#��D�vh�wB����%�p�nK�k�a��4�L�<~���|*#�Ք2;Ƙ�;�t����5w0Q����]��yO^?M_�>��(T��![ag{�f{���ؐb�pf��Rr�ô� 4��D%C����W���ju�K�s3����u~>�>����bb����ځ,�=7�K���JY5����������S��K�j������V#�ݾ�	�`�|mp�j�� v�Ѱ���d�*Y��o�Eߵ�ν��*�> O�F��H�x���
~�ÜX8^��]�֣���p9^�+�p[��C¬�P���ӣ����G���Z��Hw��'uZ�K�-��,eHy�WX[�!�)ٮ�������������i���R�Of������%�7�QT�z�r�ea֯ڵQ���^��L~��G�Ka^�� � �t���VT�V)���{�Ĵ=q�dx
Ӵ2]�}�</�a�'�����K�o��P���_�%]��R�0v�R5u��x��5�=�]�4���ײ������C�)b�TjƲ!�������h�ã�l�2V��}��n����4��Bז'�	�xo�0X�yW�[��Qb�6ў��1w�Z�<��^�=R4�
B�ex�_Åԏf��ח��ܸ�.k�>@S�Z'�uaٲpOr��.Lh�̗��w�T��h���U�p٪�8e�Gk�#h
>������$�~����:��GHh�pp�r���a=�k�~v�[k�t\�v���/k�뾗>�W6�ͥ�8+�ǈ�[�1�Ɗ(���t�M*WI�7����*p�Sj*/�{�N}�E�/�.�9�7����Ԓ*�+�\"��ի{�"�Ic/.������nN8زGr�B �M�}�{�򿩂?�ڠ����®b�X+�kp�vVV�b)��%>c�h,���~��S2]yw�K|ū԰H��n_�ׅ�xsƱ}��8`�R�
�%W]{T�9�i�6��8<�N��Qp���]FB.��Iq1��=J�7�߹x���~���ح�-���U[?�QY��<���${��M���>U����$h��t���|�
��^���ڽ�~42�NL��E���/�9h��j*�|q�Ky����4W
�yW�p�4ym7��/�ÜU��Y� �E9^-�*	����r���K��z<>Fӱ]چ�~��ws�qp�,z� h�,e�+,��.�A�~�f�������X�Qܓ;[���M;ȴe�ِ�5/Z�V5F���1ҙ���fV�!ޕ�E�;��ge���@ʽ�HX�@z�:|W���*)�󟉕S$�G+'��J��FԷ�������pTU��9��f�b��M mx�:L�η�x�T �f=��v���H�^�����͎�G\�,��Opj�-�e�)���z�z��:i���Tx2��\,`�Ws�32��I����̍�YIe�Q����*���8Дk�W��ƀn���o��d�
�'ø���%ad�w�\���F�N�AO��_�4��\���2�p�b�|'w�=�>Z۩�R�����l�ā��}������o�����b��<��ԓ^f�<� h��7i*�K�o�U^nRU[�
v��i�;�IM�z��U�F&�h�����qxT����8j�|�^9t��9Vnl�5b`�s��z'�R��E�l/�DnD�v���fУ��3m��[|��7���V-�qU�󐪝*fd-�ޘ�w�kYxk�UG(�a�8h��^'���~4�WJ��s�������xp�+~�GAh�ĕn�i�n�]A6���dx��ۺ&����B��P�]L�Ҧ:n�O?[�Ys�P��gF��X�(i��e���>�^\���Gve���fc��� TAm.	����54�tPʊ�/ ,#LcNȔ�fw{�v�����*r*�Q�ь���,v1d����s*z�j��=j�wDa��2�<�^<
��F\P�,�pi�c4��>�L���I>��]�b��G�%���wol����SG�ʭV�w�t����݅I�����ŋ��޴�$��K6n�G��Ux�;��}����¡����[^~���e�׭V{qɱ2ѧ�v|j�#��zi���c�g�>ׯ�r.If���3��ݺZ�r�ջ�K��Nڧ�q�4Ù,GM������� ,o�\��ã�6�k�~®��i���)zH�ߨװe�
�j�� Oj���F���UK5u�G�ߐY������»��B$�Y�ZI(�����36�39E
s3{L�z\`:b��u��h� h�F�yb48��?�[zFF�no�,ܸR��|#>�W������V��-��=��vg{�U=^��0�v��V+D��4F���4��ᾈT��o����>�օ^dB���8�Wc�^({Mw�w�]{�{����3��ݺ�d�1{vOz*6W���oǅ��*�h����7���Ӎk�G�:pq<5�	B�U4�&ns���˚f����S��*e�X�f���)=�>��ЫŲ*�Ek]U.���\�f��=���YWW�ϊX㷅uLf#�]*�%�9n�{$���[�/g4��
��'D��M�2�(�E�(h�O�)3�R�R�H��w�tP��?q���)a��GZG�+�3�&���I{�se��2��*�k§٨�p�0p�����Q,��trM���ק2�u7���̭߃��s�����b�y�o�*z=z�����F�,ΎzU_���ǈĽ�{�MI++�Ϳ�_���*֭	��Nb�!�W�U�Q����v�j����_˟�`������|)=@'���|�g	����"&����C�S�5���puG�>�\	5�_1�)iY�k�۾�Q�r��ecCb�	f��r�ݚ�r*���okX�����V�H��|@�Cb�Kz#?j�Vϴ��U)�cd:�~�M�/�]�,I���o.)UM�o���R�ۇD�d>{��m�Q�/�~�B�əR�!^Fa��n&,�f�r"M�q���m��B�L���S�頺/���[��ۀǄ�����R�������O�/��;�Z�Q�o�>u�/Mؔr-��a��j�z�-n5���"���b�&��U֘�}]�#�ܼ�����׉S��]�۞�EOirѯb���yY�k�s[s�zaç5���)����Ʒu��֔&E9vnEf���x�j�C�J2�eum����ta�Һ�j���;�0w�J{H�ת�[������;�u�K�L��Ձ{��)�~�B�>/�-�s�KӺh�w)K��^��=��j�i�CKt�S�Zo<8kez�J���͞p��]o,ΘDc��[='�iR���e�Gj�(�w��`ǜO��9�zOV�">WF�7"x1������K�K�`��ؤ���A��sbrzվ��ޞ�f��vs=l�_[�ޝ���hÜ��<��m�~K������̣����y�/9����9�����gj-������N�S�}��a�w�+���.=�h��^��j:3{��nV{]M��й�{���y:�}wKR���qw����ۥZLƧ�۩�>���򠘜z�r�E�<f������{�bT����
T�|�G"<���V�}=4z�ZTr�=j��@yOs��{ �2��?�����Ѱ�m*;���<V�>n=���2�ǽB�`|��j=�7&�!c/���Ѭm�[ci����j֓'�*��}w&8�$/T�V�7زd�\��ĻDcF\��������@ÚF�W}�C++]���}�۱V���ݣU���%�:������$�k��:�A�eq(>DZ����ʱ,�e2�r�m��,�j�㪻��ŋ%S�b�N�A�e�r��
r��n�cG��ˆW��
��)�4�$�滫�:�FV�v�4	�R��������t\�}ΰ�@Vdn^f��1	���SM��^�18���A��c2S:���ט�:L��+�Y�
�|*&�[�v�K�IR��vm��h�Зj���]*���҃)���,\ږ&�I��Q���rRJŧ뀛�ۻ]pĬ���g6�r<��:��r@��B<�LY�                      ����ݜ�7/{�+���_'&N%w�7��QNR-"�;�e��u��Z�(�8FxL�J�c@Q`���iD��:�V�/��bE�+Z��VO���,PN��MtX�9�'��aז�g+b��4B���n�O��ܠ�6T��i!{[�Mv*L�5�L�8;�= w����ډL�Q��r��� +o�-U�Y��)�|��u�r��\�����һ8w�u��V����(Q"C�[jٷwAV�%��H�8,,��xkO˹�m ����N>��,�JPh:�u�+���7�(#2!׷|����lPI�f�Q�c8����*+m��]�������Zpf��-
2!��l�T�NԺ�Y�;�IM2&��@ݕ;!�D���5����Hh��T^�O�1?D��1���H��(���ĊJ`�,�&*�Y�MMM9d�Q6��Z�j�n�p�8���)22�
'����hJ�Y�Q^XF�&w��U6�&��G!*����h��2hh����j����j(*B(�)Z��y�j�i��1é0��:����*���2�����0���ˉȊj�h������߷�mC䫞##1��»l�%�Z�NYZf��yt��z����Wԯ�����m"���]}����o2'��k'���.2�g6U���z#�j�B�jq�o�9'���.��!��{�aR��ܻ횫z*�^z��iы��g6U�:�̼Y���2�<�t�{-Hi�d'�������}4�5</Ooz0�eRO_l;d���{�OA��F���ߚw��jO����K&'�ݣn�ed�8�1aI{���u嗷[�r����2���q�@��>�'yvG��K.˾+ܗL�)�P�|���Z�N�Z\���>X�߻�Ȓ�ԩ��̉r���('L#w]��gjb#@�r�H�%.'22�A:�Vݗ�l2�%�u�-�c �\p�m
i���'����ޟ����t?eV��ׯj7�
|���C喳D��BS�*�[q�z3<zwXw�m�Z���ɿ�����q��{h�fk�yLʧkڥݽ���= waGCL�M{r�nTC<gTZÇk|������z&��?em��a��F/zp�TCӆ��qw�	�C� �0^����^p\��2�9���{
�x�s�<b����am).TJɼ�}o��Pq�,�*;^��q��׆:P-����\�OLлRa�7_�>�S�F� *���;�!{e�NY�
�lb]I�:�����]!ɾa��pm-��b�����Gtsb����v�2vu��'wݡ�ap�2��O+��v��c0�����X���ğ~S��o�Nv�gb�[�7Vj�k���g���o<��L�8�*��&I%zMU��e5�M�7�������
M�x�o�އ���g+�,FV�=.����>��]�,��)m2[ϴ�(�3���_���z\�9u^���*�y�X��K���$�b[E�-*W3Q��=��.�څ�2�����U�pp�<�PRar���u�ً�S�znj���B��U�MG�s��2|=�
��)��]�j��b�q*�}�8׫c����y3/Ȭ�sH���ޫ1XӅ(0^���Q�=3{�0��L��i>�n8C�F[vS�j���q����us�n���}�	��{ս[�z�j�_�[�N,�O`-�s�����WΧ�;.��*��w��c껎z�=ĭ��o�'��\�gV�|�V�̵�:�
>�:�~ک7(q���)�t0��˒a���[�ӧ�V�yY���n˹�Z�޴/:�p~���#Wݯ7�{��6BiOb�X�g�sR8�;&sCͽ@���m�X�^�B�>��.��u�й�f��Qz�\�㌝�Yv�}Iإ\R����bJ48��K}ѩ=���G�Y���iW븝��޳{�g�x�k�g�nb����в&*x�(�M�m���[d�+]부��9�W�2 :��s�Ð����ssN*WYˡ\�َ.���͉����5M_O�W�<�j����l���NI/=zN�ה��{����O)[�����}^�����A����V�;]�e�����x�9y�MX��<�޿��g�f�`�vඤ<��>��G<u�ڬ��0/b��Ի;���U�is�b���R�C�j���I��^*���:�=�X�y�?;�=����Y7^�V�+K(q����f�Ȁ:t|�{���w;B�w�JW��$���眔~�^��Z=k���
��W)�]9׸&|5,����cRt�}&���[���U��{�.�;�ͧa-� ���{YQBt�>��g`�y��)FO�ˎ�Y���ژ1!t0NK��`�$�?�ļ|G�<���6��|�9]����C��������Y���l�탁eOz��n�Oh��[��g�B�уջ����b�+؝�aA�|h�|�M_z^U3�~��[�>�5�o�߽��Օ"sN_���{�\�-C����=	�E�Ʈ=c=�V:����3�-�k����gH�� �p��5OSÖ�LT3r*a���2r��L�o�z��S)���G�ݣB+8���|���c}5@-�b�+��и���͊���u���̲9�@����6U�m�f��'w���ϔ�_��%���5�z�B�r��RZ�5�(i��|�B\[8+>�3��Ϳ?z;��=<�^�̜|����z�Gg����,���פ<�d����+���vy�c7V%��o�i�AՁ��l�`\ON�-L�@M�B��I� �[ގ0��1��-��o�8�NMg�FW{q��Yogf%oo˹\bێ�s��UV`�G�JQ�}��.y��^��Z���.,O����A�8�㩍k���s�؎�5>��;����zO�~�ӽ���>�4��?�L�m�OVfᙔ<��X
�UKmOM�0P>�J���p۸�x4�b(��ֵ�2��f��{�^���d�C�-HH-i�NȮ+�nf�]�[���n��i��k����2pc�V	��=(���,��>���a��1�=��u��usc6}�v����)Z��LR>;h����6�%� �����z<�Q�
=�����6���tn�~2(����5�GKJ�OړD]�ͽ�&'[��*%��T�R:��y{\��w��-#=�J9���u�E�M��t=�L]�٫Xj^d���&��z=a:�d^sM6������{B�sp���痥kUx�����j)��g�=��?p��]-�}n��k�sPl�����m\{ug�VK���3�ʕ �S��I�߂������r1Wk8���}���2C]�>a��mq��r�Q\z�.�I�[�Wx�Dr����Lq<������̤����q<Nɭ��gV�y��~a��={�n5N\�؟lX���O�ُy�9���_e�����7�an�z���kH&u�{Y�T`���x����dG�2��LI�G���̉z�r-/eϞO��0�8̕r����jϕA�=7�T�����Sޕ�o�>�N�T���ڙ�A�7�;|�J��Q1�oV���F<��}~t4���ooԮ	-=M����)��H vE����K���(�����#w�J��^��Vk'�h7J�Z6��
�|lb�c۴)q�N��D�4d���r�9h���X��c��rݢ.�A���lA�2�;
�n-"��ּ��������K����*�����$y�S��ɴ��n6��t{V�g��:ٹ�'�����;�{��/8��4��5����&t�������I�XU�QV�#یl'�p>�gG
�'���$����x�v{�S6G�����iVr����7��/Hp�P���x�-��?n���}i���*|n?�_��ˊ���g�p �
�Т��_��w�+g=�� ]4�f�/4�[������:��=�������φ��~�Wj��=��I�,�@hE�]����[� ��l�ʛ <N��+ۧ����B�O:�a��z�Pe�͡�2:G[��P����ۨ*`��������J����G))Jڱ�P�S�ޡ+朽[i��F�u{7l�5��q ,��ŝ��8.�5��O)��C��n��Q+��S1�����%�r��.�ز��_Мwl��SlGe���>]�s�q�A%�n���3)S��@R�|V�û���ô���f},�bQٝ���t��� W��h>z��r��`��i��ѨT�SI8������J�;�Ѭ
}�F��;��N��F�

YN,�'p����ӚvMt��SZx�A)1+ŶƘYۻ�m���$�b��5{p�ϕ����<�ї��Ή��f�]�V3X�z�7+r=ȵ�W�D�,辠�                     �d��N�*o����X!���S���j$G�>���螧rA�#m3�� ـ��f:���"yR'E�z��y�f�ǈ	����d��3,����k�he${�*f�!�܌gVtOh��|)�h7\����U�6zZ8����`���M�媶�޻�EV��.7���l�w�M����:y���E��8ݖ��8V�AWTF��42<z���6n��>�D�Yj�z��,q�4WV�"����V���$UVwRX��ĩ���%8Ϋ̫��p�t��S'X�5Vgښ�r&�+F`h�&��V9��Z�U�sKp�2J�
����/h�R�NL]�p�nk��`�%��nAX(j�������{ʧt^�`Dʬ�Y���7�������(��
H����:���i��bh������"�����¼�"�(i(�ʌ�����Ȥhb�(�*���+�
)(�j�s"�i=̦�J
wcLEKU-WY氪�(Jj�;�!*���
��"�))��)��ZZ
�h���.'R4T�@DQM%4�WvIE�2
(:����QT�)C@�KIHR�P�y���ﮎ��1Sϗ_.3���"뤳�l��E�N� "�@01�sQ�`�ds��Y�?ᴵe�W���`b�k/�:yH�>;v+�{�3z/�u{pf�1j�5���LՏoo�(�>�)�������%�w	׮�r����:j�eoEC�z�0����f��o$W�+;�~�xv��L)���:���8��c�{�����E��v�MF�Bc~��g�ym�e[����^����ط 6;t���mz,�p@M�t\�Ϡ�y�{�>l����
o���0���:�$��ȟb�~���8��t��e�ۉ_�w��fߡ�^�cb��3Ǟt~��]?mU��Pύז�
F�[�Q��l3�>����G"�R��Y��ȕgqG:ێ�7���CeÜ�9[���}U��6��##k���S�z�?dߊ�C
Z�w�	?/z�����*���3'+��;wt*�C�;��e�oT�
�SQ�Nj�R�+=�n�����l|�8K�5W�#��4�#�������ΛI#�,6$���w� {sT�U��M�l���Os�x6m86����)5h:�+�o���<���e:�e��%��l��=�'�0A�������!׽S�Z��_���v���V�q��,����v�^^�s]
�n�
��u�4�bg;��/�rN{3-1ȿfO��6E�ڒ�Y�����Avd�k��v��vk}�Ҳ �x��������|9�z�Qf��+}s�a�y��]�b�.�i�����l�$���eb٫����}�xo��ڱ 
��\k#}���Z����ۂ۬�ى�	����w�U�t�ޯrw���q1�)��N���U���8�dZ���U�^�l�s����}W]Jm�P�C�?f��m`$��yڵ�*��9�OT�'�/�T� �K�S�k��6��Z˺�N�U�Kʙ4�%��C�[��,9ֻ�E����R�\���EO{QRGuݓ�{.������Ⱥ�Rt��=K[�@L>���X��{��ps+)Ԫ�ץ��՚ֲ��e�"z�����V~��=�Fݐ皋q�.��NcēܿUb� �霶�c�=�E����]�5�/����ˎ4��@B����?��e�0B>��f�w%h�����'% � T�v�m���eF3���kfz�r��;Ը���*c��=O�����^=���3��ޓ{�q�z��X�n�~ʞ�h��6]��V��X�9�;/;�ٱ V�nww����dc��zg7Ea�mM�Zrٍ6�C]�i�˂<3
�t��i|}79y�H�f�銙�֍�U���
�= �^�o`kF�ܻ��;���.E�X����I�Λ\�q/��EG�_�u���!�p绢��[F<�iF�}�ټ�%�F	$�AĮ�μ2�-ӷO�\���8ےD�@���1���vm�+3en��i���o!8fe�UԞ\�1:O?�;'�s�~�L�+j;�6i��^��٤����K��;������yuՉ��S��9"1�:���]�I��sW�x���c��Y����,����.��ޞ�VZ�j�Ѿ�kq�&�#�Guu��d��s���n�N	� �[��y��h��[]��	�Z��Pm�y�s�o��yۥe���5�Qзy;�����C����1�'FAS��
b��N]�eoC�z~�t�o�����JW�nuD_���vG��⩋��b�v�zMy�s�u�oծ7Ƿz�*�W˂=;HX�|)t�0N�>��[�gŷG�+�;1ɞ�o[�U����MV�]lX�Ի2>e��	̎mj�^��3T���K�a��?{�%j̩�:�Fz�l_<�۵��=~"��u�y�u��{v{��73wZ\�6޺�zv�o?+�)D��yL!繯=��e�d#o����G�{3�TI7��h��5��F@�s�TC潬��Y�����9�~�38�Nw���V�_��ی�\N��������̻?ie+=m.���S��~����y^9�4��f��M�>$����T\z�c{MSB]QfVC͌u*� dTW�uS|��fJPoܻ�I�(�5�<�L�tБ�g���콴�}��.�|E�;��|�p#us�0��}�!hO�m䒷kiF�0^��6��h���y�ޜ{l㥸.#�.\�����\�/\��Q�ux�����P��	�׾�Z̕P�!�vյ!�a���u��;j�=*e�C�٩�g���2�m�O�m�/}<�q�4E 1?�����_�� �,��F�����gb ��\Tuf�Qx�V���0���Ԏ�.�kCC5�G���Ц�{�k��YO��z����^�����ʒ:/j����JZ��@n$���+W}ԙ�C�v<�^e��ޒMYި��ϣ�) ]�Z���V��ޝJļjÇ1՛]��p%_=�܄�&��]y�#��h��%�3I)(�V\LX�������m���]�aoVҳ�S��g93�3p~��L�=/(����q���N�a(�/$g�$���g�f�GZ��TY����`n�>�E�[�Ʌ�)m��n=�ż�����I7y��V�)[�οC�ALp�S��H!��{�Ӑ��Wk�*���-M^�y�3W &T8ǭ�B�W�7�Mp�|b����M��M�OΣ����Ɋ��m�Ζ�y�������ϳ��o��7$?B�5�.xY�=}[�8�=��[<f_���!��tEI���TGՀd���'9����y��vJ�w��]���w�W��Q;]wg�7�#}Y�H���F�=5�"�c��r�������r!zq[�.�[kn���3͵�o�	:\�B�'Fi�mH&4��������E?A�;M!�����R��oϱ��6܋�I�i�h[=k��i=��-��c�n8��b���r���5��Bk���6v���s����[��z"�b^p���='%etg��砽�Ye�Y�nn�^�gyn7�勯y��y��~�"k��=����f�{�b����^�`�ql�`���Ȩ�9������~�TNE� **�x�˪7��S��[xՊ��-Cל|T���s�=M�Ԓy�6��mj�.ǔ�Rzy�:H�w팺��������]Y����d�.G�%{�#-�<�0�Z�K�ٮ�׺3z�6 |��oQ�IH�\bey��R��8Tr��O<A�8����2������6Ed�~ү���+T�GB���Mq����Y�y���q�\����ދez���r"�_ȬX���^ˉy�u�{Li�߷4C)ǽ�z�xċ�1���ɣ�q���R���g0b��}C��SU=��*�U����|5=���f�:��=�=/g*W��b���ah�xW��~O��N�+=�OP)��l�\HN��e�ۉy�w��U��F��n�����#;J�}s���3�����?�.I/y�����,+�?r�wǛ����~���W��������KUEX�(������ڊ���q���H���SA��i�y�8C��������y���=#|�AH�Q@��P2E�UF�Z�u٧��911.p1��P���?�<L�<t��b�)�b�����L����C_�����W��|��'�~��Q��YJ^e&,N�^t������N��g���}�|h�0���՝��0F��S����UUE����l_��M6�RM�$?2��"��a�U��1��khر��~Yҏ,V~{.g����9�N�iȒ���H�H���H�[�s�⤥(k�E���]$b�y邑�\�e���Q���ڳ�"��"��_)%�ps���A���_��A9�����ܘ��(G��ɏ�<�Y�����tDp �DyO�*�.*�7����wP�˘�yg��7���i��lz$I$Hm�)*UUIgG(o&<�l&�s�#��R���M)����p�dc�:'�~ƶ/a��=�u�G���f�)R�I$�y%���xp<dmd��y�w��~�e�˦�ZE�{x����˫��X��1'��n�zͥ�I9̻�>����r�$�!�u�J+>�_�(��z�1L٘��R��a��u�*Z�0�I���<�$�$>G�=�SIX��NUiUdp\a��K0I��L�ŉX��2m��C#!�zQURjt_���O�k�TC^L^G�!O�~��y�����Iֲ�p�b>�&��܄:�0M���,˕_l�>�I$Hj�<�'sZGL��I�^.ԟ�I%�-�攞O�����#暇���ދ�9��lad���J.���y��f�u��~�葇φ��0�|V�$�!��7���[�Uz�k,��w���$�$-'�&]�g.��(y&�Y��5&�l�Ļj=?�ߢw�v�:H�oۇ�W��rmPǿ����Q���F��UV�����Bij7�ۇi�)I��GJ2�8Ǝ����mٖ*����,��I�y7k����(سG^V�a��#�\tQ(H�'������U�;�[�3��	!�N�jo�L�a�vvY:yn���~�!�z�'J~ILA�����[b&��D���H�
	��`