BZh91AY&SY��֓�_�py����߰����  aM^�      � �@ ( �@P  ���	@�PDHJ�Ѥ�
�P�P

JU(�D��QT���T��6��IJ�mǁ>�� |@  	    ��� ����v�7ov�ǣ������ztvݻ�˧;��^^��t� 

�v�+�y���wVi�;:C{���:��7סU���i]k��������/�>G�_m�u���^���������؀ |�<��Ts�� �u}h����B�������!��_x��4�}�^��i�H�@g:9N�)֪  C��餫A�o `'j�k)M���7 pnw���d6�L�K��ΟZ�,��0 ��.��#v�8�ٕ,�T�i�3�%��n�:� LON�W�d�Iy�����riZ��Πp�Y)��F��7���2�E4=�� �a�>�y�+{MhN�	r7�:�L�3�uZʍ7����3�Ϸ���� ��dSFCMv�SN��΍=F���Ǡ` �ޏiY�Ҁ�  ���h�gaѠ���y������=�_`��@x�m��7���rs���nz���z:u��!݀m�	n��]�^��3�                       (  F�hUSу�R�T�SF��i��A�2��!%*��2d�@CA�0L4�D��U7�A�F � d���@��)�L��F�� �i�MRA#S1��jd��O§�g��=S'��BfT�J220# i���7��}
��\����[�T�ql��w�VϷy�jzO/��'o�}��͌37ь6��������3a�;�v�����~o���~��O�ϫ����u���0�F��q�6۴z��mۜq��r�o��6f��Y�f|�6�-�ʪ������zX�����������1����~�Ʊ����'�0����4�k��4��ϩ��\��Z���$�l�N��q�����u��ěa.�z�z�X�ǭ��x�MN�q�Y�&R�L��%�$�^�R��M-T���k[��uzmN�ɧ���'�,a�la$�S�m8��&�I��~�I7"z��bI$��$�)�$��v=x�)1�I$���u$�z�w�N�N%��y�$��I4�k�a$�mX���{${���x�Kx�M0���'�%�I2�Zǉ&�nX�i����I7�$�]��SOR�q%�u���&�4�I6����8�Z�^��x���Ē�$�2�^bMe$�q8�)gI��=I,�I:�����$�%��I:�_�SΧ�$�\a$����z�7�I:���&Q-4���q�MG&���-�a=a�z����OeɄ�e~�i4�_��i'���q&c>:��I�rORO8I'$�ԙ�I�M��q:�i�<D�i�2�q�'�G��O0�a$��:�I�獼r&�e��M���֞"z��I4�w���I��SI��lI:�iq��z�os�'���x�I�<u1=I4�Jc�m=a�2OI����Iل�{$��<e$��'L"�	'���z���qĒn�4�K�M$�$�RI�$����a"_�RL�$�v0���x��a��y$�y�G^��'^���'�$��ba8���z�oiٗ���I'x�~�e$��z�O}�I8���^$�L$�n��	�Oy����I9��2��m��L��I&d�i׿��$�XI'�L$�x�I$�z�I$��$ƒjM$Ӿ��$����$ēԓ����$�X�$�_�I$α$�ig�RIw��0���$�Li�I��.��D�va$�2I6�V0�IͲ��x�θ�$��x�ML���I"wX�I4�2I4�y:�S��,���6�I't�Ԟ��:�x�7�u$̒F�X�I'$��M&s�I���^&jI2�u&�gX�&�m��I;:�$�����8�I��)4�5�I�RrL�ћtM�f�����thl��t'�V�w��z�������.�m�c׏m�=X�t�L��`�OV1$�9�<I&Y]�����s�a�I>�8�Zē����e.�x�^�I��ʱ���[�a��y�$��ԙK8�M$��I,�I&��i'���q'����RI6����-bI=i~�F˸�$������u����ic���1<I%�I�H��$����i�ZěI�=ęIwz�I{��bx��q��j�*�=Oc�=��q񇺦����u)����/�	=[��N7c�f�$��'�&�/^�4���4��:q�/��6�T�峬M��k|y;�y�rN=�4��$�q8�{�%�I�lz�%�I;s�Z\ik�����z��>LZ�5��������i�I��-KO[�I���'��?M:�{�&x���<�<IX�im�����0�N�q��k8�m7�~�e<�<N3�$�[�m��$�Ɯq~�$߉<��M4�q���R\ĝg�I2��&�m�	��$�q�ӭ/�h�x�z͌$�Ĝa~�'��bI��I����q0�����ē^c)-�IX�oR�&��4�ӎ�댽w�<���S��q<m��4�LkI6�N��1'^2�w�I�ĿN$����L��ĒIq�<ORg8�I��~�I7$�/�ęI5�I��I�$�n�z�{�$��$�i<��ǩ'}�J�Z�1�c��1��3�q��I�ұ׉����IcIoL��I5���4�K8�I�I%�I�N�q�I��q'�-bI4�2ĒNkI4�ĒI�<�2�~�I%�q$��$�XĒJ�IgI7c	$��=Iy�$���0�'�8�M:�u�I��$�K�N��x�u�I՜N��K�Iש1�N�I9�$���y�$�|ē�I瘒I9c�I<�$�v�^:�$�ԘN��׉'���ԗw瓯I�1$�No��1�|p�1&��0�q&�1u����-�k����/|�KX���i=m6u�X�L�'��?m8�7;T���>�ZV��x�����i8��׬�����:͍<M��u�+g8�zî�c��L��I$���z�?��i~�f&��'k�~�I5�I�e~�I&��ԙ_��$Ӊ�cm��g��0����m�s����M��6�a���2�k^�ǿ�i<�	���S�p�M~��=G�,�6ѩɳ�'�闛Ǽ�=I����O��$��'��I{��N�&��<I{�4��K�X�M<�s8���bi������w��q�m4�70����N�c]0�{4�z�c/~t�<�&}z�I�U�$�k8�8��S�ㆢ�U̝.&l����<eⱶ^=a~�.�x�y��O}��=z��'���m��i��kYIg�W�$��$��c	;�#)4���o^�R{�L�^��N����qs	�^��c���sO���ާ�X�[�\L2����'k�a%�'�.�xI�1�mM+siU�k}��Ki~�U���bOYL����N�]u�z�9Ēu��$��OY/�1�I���8��Y{$���x�e~�Ēu<�ԒO;�8�O]��M18�L�<I�la$��?mX���Ogx���x�&���?_��$��8�a䓩�S�<�xi<�M%�u{��O��e~넒z��z�Mi�I2��I6���z�&$�N'r�&^$��'W��o?D�Zđ&��$��:�d��q$�e,c-$�\ƛI����m%�IԝLs=Ncx�I$�{$I6_�I$�rORfN��n��e�I���ƞ�$��Ҝi�N��mo{0ˍ��I���I�&�=�i&֝e�^L�Z�8ĘM�&S2�6�H�vx�q��I:�m�u�Yi�1�I���q�x����Rfm�M$��0���Me9��-{K���Nt�ou��cMZV��-7������4˩�6띌��SL��	��fa��M���/=����}�7ĥ�J�j[�枷38��q��z��8���N=�	�~�rm9����=Z�î�6������sz�e$��&�va��$��%�a~m�ן��4�y�=c)��ck��N��m��M�0�w�u;�u8���ӌ�e�e��M�=��3I�ʱ��y�3�5�N�����,c������<V6�L��u0����:��m4��Ox��$��i���ؐ�6�5�՟Yv�o�@L�lO��?o�q����ϼ3s�9��T�Ck���>o�wͼ�Ϊ����R�q|���?zY}�_�i�y�n�-�=S�t�~ǣvN�翻����җ��?,���.��q�ܓ��u���{�\�u�u��o�ۭ��9�s��͵�K�Z޹��|�\��s{ׯ{�9����g<��u~v�;�Oh�<ٜ�w}ޗW~s��wxo4�s2�Ξ�T��}�7����67�4�z�"O9}O<�η���<�߮��������?�~|�ݾ���������]��w6����~Mk]�蛚�pgǯ�O�T�o��vO��OO��y�t������^����v^ض���:��x����|/ީ�����|{��ߝ�<'���ש�n���x�l�y���~r_��׳�C���1���oo��?����쿷��3�����O���{�}��������6rݶ�W�Zy�;!{�kd�Y���&;��S���;�O5V�u��|~����#sv��*F���n���[�|�zo}�ͼ�u�����{���~�_z��ϛ}�oe�νN������n_���}��>=߯�7��\R���ϯ����ֲ�k����3��zy<7�oz��o�%��Zu�J�{sJnn�w�[�������]��w������c�ɋ�=1����W�n�ϯ��咜��l�_ߞ��N�R~����(x���3/�m}Ҙ�KYo�}�{������/��z~�{�zt��󫟎�;>G/_;羾��~��F��N�>���}�*��x�y����)�\SY���B�ü�V�u{�����<w��rky��\��f�݆��3+Z��/��3Ww{��O��y�>�}���u���պ9�q<���Ӿ�T�}�}���=?��K��wx�>{=�՟��z6�'�;Լﻻ���|�h�6�.oW�����Y��wz:�s/�t����q�{��5}��7��wk����W/y||�����f�W�����J&�W�Ɲ;5�	z��g�_Ǜ��9��W����{���G�LoLWyޞ����ӧD�cæ��y��c���Ӷ3>��5�J���/��[���ò;a�o	:�;��������zzQ🗠{�~<~�������>��;䩊}�ǅ��Z��#5���Ǜw:w����@�g%�y��y~_=����@N�:6x<��v�d�;q�9�˷�f���+���/"m�yw}z��<��8�}�q��P:x~��ߜ�e�Rӡ��|�۷���o�vi�j[�<C�w�d���<D�������������mD[�P>��uP�M��t�[�N���A�|����:z~�ϠS[���c�寘��|��L�ۥxۏ����]�m�N�kק�˝��j⚑��m�=�v���[zϻ�k��?vߵ7��M4҈ ?_���M�o��{�����׌�oN���uۛ�_\}��4c�=b�m�n���n�N6��}y���:]sܽ}}��c�ju㷿^Jq)���L'wZ~ޟn�?���	�=�l��^+�ˬ��~��V�^8�1Ǉ������m��n�˳�(t���7�����m��������T}3��ӣ5�W�8��;�_�|��\ϯ��\}��;t�7/O?1���_^�m�o�{u2�]��ׯ����ݼc�Ռ��6g�t���k�������im�]���_\v�~eX���O\�y�~$���ˏC�ߺ��]�vc��z֕���r��<ܜޱ{��n���޽�_7<λV��>e��q1޹xܞwx�\���5n�����i����!�7�7�}��ߥ���ߦ��4�Ϻx��zy}:n���P�c�t��S;�N��{Șq㬷W�[��ks����|�/��Y�u�k왞���oo����<�e��ow�������^,���Z�^�q�w��ӽ��]��zpg\�w�t��y����S�4��:��Cy@��s�����鏼�~����Ӿ#%�����w�n���z��Hy�~������s�����_sN�p�;����ҟ�im����-����t�[�z�^���OO<�~���߼~߿>9O��s������.���:����/�gN�L[�����u{���߿=��ڻ���}̼�z���z���39~x���O�ܾ�W��y�k�����~�׽���h��|�~���Ϻ^�������������w�޷�m�\�Λ�m��u�p��|�;�e�㗽9�7{��֦��k���y�k_g{�{�ߋ7}�nv�{z�O>���h���־x����_5�on����{oٞ�-��P�{-=����䩤��C���}�u>�;���6>��߯<�/�����ֶLmκ�ߟgkھ��}�{��\��;�}�����7/�^���ԯ��l%/�>J��!��|.��'��;6,k��ͺyW���M5�?��\o���\]h�I��S}Ӓ���z�_y�����o����;���;�/�y�t�������?����~�~���m����=�����͘���ߴ�-�|wϟ�����xv�����i�w?��u9��b�~����������|�~�U�{ݟh�������g��o�~�������/���}��
���{����CzQ��>�{��'yV{�����������v����xo������m���N���y������&h2w�浭�u۳���}i������=��@;�|\o7�{P|����C�N�����z_f�z^���W�=ǚ�iw�W�<��\n�v����Yb�������wn����>xE�/|^��Gߋ����37�h�5�A���,ތn��f��w����ѯb��۳��Ǜ�z�����OK�r�����ۻ�}�z�y��������M\1�����=���7K��_a�z�ҹzWc~;�]<��o݆N��;��_��_7��z�y)��O����}���=Z=����l��/J�mܿx�e|(��==��z�oOGϟ篿|��Rzo�\��Bi��y̺�:�i{��Ƚ\����S��P��<����}�A(����g��l��g�M���7�>:#ٷfNo��ۗz�{�ޖ��J��5<�ٶe��>Ǟsy~�w��|������W�����n��޿z�{�e�Y������wd,�7�*}�we3�H���ϼ�o.7_�h�<�gM<���Zk={��څ콷Nf�~t�Y�y�~�n���������O�o;����������ݞ�_߻7��6��J�/��1��H~|� �b��v�{��{�����oL�;���'�wz����z���}��w/���N��Ӧ����l���}��׳���o�察kv�4���<��'�z����>/����z
����Ǜ��k�����⯏�K���>x�5����o�3~�w}��r�o����9��_�~�o����z�xt������'�����z�������w��~�=�z�c���}�>���å)�S�\vL���ќv���l�ӥz�}��_�ӧ��?=�G���W�K�7e'ցҺ��'����~��G��N���K}�=ˊY{�S����co���=_�u�o^�^��1{��f�������ɧJ\�ٷn�{�]u�]ƾ~}��Sǭ�Zzyr�����V����>��^��{��>��t�ly�U_��u��U�קN���񫽇��篝s��s�����\�ӝի�}~��o�j��������fv������g0潟�ߖv���{�M5�jw����3<�ϟ}/���߲�1߼P��u�|�_{��|��}o�����n����6{�5��ս_<��侾z_g�7�|�o:�[�^�w}�쓖O,��9��u.{���~�MwN7��î��vs6zG�߻�>��1��;�{���}'�ǳO?w=�s[����}�׮k}�~��{��[�j0�3w��k/�^�2o���}���7߽�wY�ݾ��ձ9��/Y�������׫�Ӗo]�9��:��;�_����o�[���w�����w맃{�w�:;�|���w������%���Z̼�o�{��<㝻��~�^]��s5�gw>�������g/7�o�7��:o����Z�i湓9zy�NaV��V�=���/M���i�������w_,�fwv����׵���w9�����9�g�=O��<��~)����}�,��{�~�����kW}i�g5z��4}{�w��i�ׯ/p���������v��{�n�n��]���9�l�}�}��{:y�7�%7�|0n|��|�M�λ��῭�{�z���y���:�o���=ޜ�:��ns���(���mW�s���ZKu���^���VO��>\��u�|s�Ȧ�=�ҟ�7?�6k?��)	����l-l��m�ێG84�C]9��\�ך��Z]5%6@�fI5t��ܵ���x��݂�67��d�3,�4�M���3k&�X�fK�k�it�n% �֚ҸSuZջ��&���XK[��7ZB��"����L�t�4���P�Im
�bF�2���
(�j�����l�v�29.��H�A��Nи��jͮ��],:u���̚W����IL�fd��������53W �sJF鲪K1��Ԏ�?�4�:�[G�ǰc-V�+q͚��jkDz��m
u+�҅ZB���Q��+z�h�D�^M0��KX�33136j�m�%Bi[>2S^��xb�R4���t���&�<�b�L�
۵I�W��(�m�GNs�|NI�n��)�$�ge ��d=�;����e��N;[��pḀ�B�ZV1xnc���|��{��%�iKT8�Qƨ>��ף�����`ƘH!��eШ�[f��1�a��n����n�p�9��s���4�/�����Ī�٦�������~�&Ű�{��r��6(Y�y)m�'9���S��%Ф����Km4A��%u5$e��ь�C�U����6j�iq>�I���W߷C��6�Mu�[�����6��p�*RJʰxk�v��c�d��9)�d�<�N��4��L�۰m��Y MY9XN�7�+�X�Q��66Ie�6&�ڸΌ�:��1����b�a�l�zS�q2���JoRWr�ɫ�1������ꌕf�o�f����l��&�>��&ë$�b�,�qt,���9)���������f���$���l�u4� `2�&n�g���q�e��]��9�,�K0+�$���8������B�y@��'"ͱ�ٔmˤVH;Rn��9����I��23FhSl�2��VV�I�]t�&����y<�|��I�SZ]��z�hq,ۜ-�|�N�{�4���ۗPjl��q#�Iw�B��Ma��I�- i˕�:ɡ1�
���2�kS���1�,���������5��!�%;l	�B}� �3곕��(d��Dͮ�^ff�8Os�8����������?�!�4��g����W9���lo]��yyO�����G��������z�o������$�s���ۓ�m[m[	a�a��r߿~~c�߿c�����������T���yUf��b����Z�튪�Vj����*��X��쪪��UWkU]�UX�Uv�^�1U^UU��UW����Vs�Z�Vj�UY��X��쪪����c����c����r�
Ęr�Q�k��j6�M�rf�a�M��-�ܶ3�;s1�͒�F��im��s���������U�U\�U\�*�UY�ʪ�*��ت�W+˵Z��U��U^�V�UY��Uj��U�������+ګ5V���Z��Ug9�m⪫��U[��ث5w|������DGҙ2��ELDJD;[=;q��j�rq`���0~~ǖj�j��V���������Uj�5yUW%UUJ���*��^UU��=���b����UW+ʫ5V���.ت��b��튪����gU���ʪ��U\�*��y�~���`?V�c�m��͹��[9s�6S�=f�̈v�ɜ��ڥrp�%j4����Vẍ�um���ԭ����ͷ!SE)rPZ��a%]�@�E�]��ܚ����㓟G��}M�����JU����������������M�G�?�z���	$�$�L$�I��I$e֒OM<D��RIěq�L��I8�<m��$�e$�I'��I��I6�I��֒I�ZI�Yu�[I��I$�L$�L��N��q���&I'ORI&��<e$��z�$�I��e��$�L��x��<DI���OXI'��i��G�&u��L��&�z��D�I�Çq�qē�ORI$�	��&�4�q��u��z��a��I�i4�ߏ�����y$g��/��w�]�v�Y���-e�����,�
Sm.#^CmRZ��[�r7f0�)`�5�m�mc��s[1-�6�M
�m�rRjsJ�:�jly2���;B�l���E���P�Xh�Y���b�J��V�8m����]	��ꑆF74��6m���Tv��ژik�q������4hK�5��6c��`��^&r�;Wg]uk]�N�j��4!Il��r�n����@�[ݘL�	29�;���F�v��a�Ɔ��[ô�K5�%r��4'N���9���͖��*jd�	�Ť#���3t�ĩt`�\]�fѶ5f���ѻ�cB��~�핇x$���a�Q �;�����~�.��R�pY�c�Z�0���\9K4�v�-�m�
۪����Ll���G������8Ղk�1��ne�Ͷ�v����Σ�U%�)�M�h�2��K���gl ���`mM)o1�I���ke���1.&���J٥*9ɐt]�j��Q�!iq2�Y�	ae#h�[v%�h��Y�3<Lm�nexm��[`��7%J18eK�Y��`ޡe]��]	�m��R�R<-f����h�-�n��J�ݓX��
���G5�8�Qd��A��:�]kE�Cv�k]*p��1x�iy�Лsi�5�e��Q��й�1ii�6yk5�$cim�ZGYc�%-�&�ŹT�irBAx��V[3eK�]���a�+�#�������]�(8`\�5���e�.�%���	0`L�<��[��\FR).sZrdJG'	f�&X�}�Y�[���Yq�ՀY���Z̒�R�Ml,P.��0m�	���ö��β�ݣefJ��	b	0��K�Q�,��M��nYuJ�n\Z���TJJ39��"��Y�-�rM�x�)�Rl�JHA���HM!u�Q�f ����y�v-����Vӎ���KWR���-hF�v[��uֈ]��ƃJM���˜]��M�0��f!��,���hiI���ؖYfv���ZMM��,��nΈ [�ګ6���\W���R]͊�5ZE�������֤�v�M�2��\��C�e�h�ڬ��c�5p/%n6���\ŭ���lƥ�d��B6�b [CFi[�ٳ�)e��7MB��j��pF\!L3�4�t���<e4��u��[LsB�3�6��E�6iu�mb����:Սe.Uͼ�&��W6%���P"b�6kW@�Ղ[ʹ�X�	��XÕ�-�8���	���������6�+6�>a�X)|�S�ޫevlbGU����n
Ȓ�ֻg�����'(~�gH�����]lEF�F��5D��6i@�K�SRR�!�Ts�����l�n�Ef�L���KB&i+�mm6y� � ��M���K�f��\<.����.��c�1i��)�Ň��6[��K����FcR�s^[aͮs�:д㦴�R)1 �!^m3.83kie[fd0k�5���j+�1�%ቱy�2�X�\P�����g�eػ`#��c��ܓ��>����2�����{w��B�}���f]��߽�n�\�@��ff{�www�{۾W0ADu�y�uo:��X���Si:�N&a��z���p��6�V5���ѯf����)f��%��������ଭ�iTB�)1�&�#� ��j	���;4�,�U�b��h�ڻ�f����oQ#sJ�Uvv�P�v��GE���i-�m���^1��ikr�����5ٮ��ۖ�u���o',����X�u^R��n��Mu6�������t�k��\۵LJa.�2sLc0���k �5�hZMb5��xau�F�d#nj��q��R�<��)u�R��3k�r�f5�����r��(��&Ml�훡m�@X1��N��c&�̈́E�ҕ����K��j�H-m�b#`4�"%�$�0�cV[i*	��?�:{>�vt�6I���ՖmF����=M^�W��'�����tN��˻�^,2�.�0�RvX���<��2�|9⣝M�C�bk�c8Dxhh�|�,��gG!�d���vm�����UTN�3��Z�c�n<��p�r)T�My.���q����u�ο-Ku��N�����a�^�s]c���ڪ!�z��Z򵫖�Y��y�R���e�"���	�T�j%r��Uw��[H'�X��\���q�&�e5T��*�������~��2�yt������lk��p4H���Ē�5Ֆ�:J�W� ��:w��QOh�%�G��++I���Q���Qn>mN%m<��q'\q��a:�m'RIǍ�FX�y��m���R��� =�Y�'1;�?B�x4kZUj5|�Ç_�dm�55�*��eh���v���Փ�}��<��A��[岛\��48���WtW3��=	����NVW���}=|6e�.��>��!�S���B��(������%��W�WT6j�(�xN0ӭ���\q��a:�m'Rx����	�,޻ۅ�kJ�x6B�xa�şZ0�������}D��Q��>8��ҒU�	cN��Y����b4έy�s��z�ځ�V���鳢eV\Y��Fנ��h������x;��l���X@�LM�/�4�_�0ne�f��nb���F�i4}|L�\Q0|�J��b�����n?�Ϛc�u�8��S	�Si:�G &�,����e�ێ�rū�qv|��^vi��P�Gl#��L:f�`�isG�����,iLԎ��Q�!HG@�[�5��\F�K0`@�-����B�j������A�1�k���]05��A5�Y�;�-��[���<��3D٦�y��)f͗Cq�f�3m{�gh$�m�����<L�qf�bYZ恬��sv�!���j����l����a�ѓȖ0�l��VUpΚ=[6��e�Z�T�T�xh�΍�\��!W��A�5Y���]�l�S�M��4u*��Ct��χ�mOE�΄F���]U$4n����HIv>�r�Ű%����[�7h`Nh��6��HA:t}��9U\2�˭�ۉ:㍧S	�Si:��ǎ6@MYgh��)i�|���U�U
P�A�&���E*.���~G#I��[ji(���ƍeW�k��V��ҬMMr�������h��lD!��U��ej�SZ��]K��L���S1��yz�CZ�2�q;kk�%�_�/���4mW���=1��q�(����(�x��R�WtұA�H]�kz˭�u�κ㍤��Sio-k[�|�\m���n[JI����PK���s��_�Զ�}��XzҴj��¨�eQUmU�J`��0����wolW$VM�v��&�*������oK����̕%u�p�Gpf���5&��Y�s$n�W�d$����a���5�꫚OŶ��u���ng�D%�5GҟRy��(����>�[=p�%��/U�������n��K<m����\q��:�m'RI���	�,Ms�Z[1UU�S��
�wGW�4'�F��ˣF��{rl��!]3�0r�k*�Xk�͡t�l�t�[�n�����yٹ<��1����K��F��R�ӕ"f{TQd����^��f�v����r��%PacE��!��uU����ʭѪ0��Y����Ά�0�P�ؕ��PY�/>�̳3/9j+ ����>Sj�q�O��^u�ɛu�qƜq�ϝq��$N��Iԝ�O�e��h�~�~����՟9�j�O�4!䕳��˳�q��oFTx�B�荷x�I�j�[_����ص�Mn\lJ,p	-�s�� I^�ʡ�D�,Ĥ��Ks�%m�sr��x"�9�v֍F��!��ev��j�Ҫ������@ږ��.+Z>,���*��k%}�$у\��`] j������gU	�nI�*sf��6B�o�+�M������UX}C{�C�aq|yy\4Y�at�ּ�rD�7%��x��:�@�j�����Nϗ��!8�V��m�ٕ���72�]H�&e�sl`,���3�B�+��酎ZXY��n�0�gu��[�ou:���/�:T4ӏ-�1�8�o�L:�m'S���O2�e�c�4Mi�U���=],�E/��&�3Z8e��b|�-PP���.��X�#�Z��ՠLJ�#���մ��d�#q���bcW/65����Y�����W?�'�=���.�KH�-.�6�d�be��1�W&4eh�Yσ	UW�F!tu5W)2���x���PQ_*%�r"K�E����&d�^�B�}���Y*�W�͎��ڟ���]m[N&S�8�5�S�T��bm�c�V2��1�N'�eO����1V�]olT�R�1]c�bq�����V%�+�X�c��|�ۭu�S8�N'�V1Xŵ�V'��Ʊ���z�b���+�Z�֚��q�c�)��V��X�m^�긵Zե��y��V��M�X�bv�52���b|�GX�'i�p�L�1R�Jq2�bi�ɜW�N'VL⼝�ⱊ�����a[b��iZb��b���+�1�N8�N)X�cj�����c�)M*���,��S��t�4���|O�?N��j	�á�%i�ߚ��N&���یk��~b��8�1_:���))��k��V1X�c�T����jZmj���LjX�eN1�u�c�)LU1X�O�b~N1^M's3�<~S�x�J�<,�G����k��	��4�bv�cϚ�Џ��.��d���Vwz��#�М3ގ�=�˻����D���ic��>o�}�GK1���y���:���!�Y�M��Y-X��M���02?����Ħ��B�o׬$��wzl��na���e�_.*�fHċr��GЅr��^�V�0�r��o���νM_}��?1�0J2�J$��"@�r�aa.�R�S��w��R�v�,H��{iC�e��^{�D&��s���[R��9ň�d���$�{�e��p�枓�7�ܵ�rcޞ2�����B#��;����www��=9�}��!�ٙ�̜����{�̯�ޠ}�ffw2s2����s3ﵸ�8�����:㍾H�u6��:�����4h���$����� «u����85Ub�W�n����dQ"&<�#�!Ɣ9*UB�m����hw�S�UJStVJ%V��u���[8C6<����۸܍�����[���sv��Y�u6힎lw�R�u�韱��k�V8�f�2�{�8��΅�sZ2�ٴ�T#���Ԙ������ɂ�"P֝km&D���X�N6��w���.Ǎ� j���W
�(�j�o�W�ou�SyM'�e���v�W��(8a������Z��_RG�A��<mCR�`m1K�3C�DnbZ���U)2��MW�zm�,vN�p�wM蝞71��T#��GLLB���"���~c�u��<y�^y�^yռ��i"B4a���
�[B���U
Y��o��m���q����1"V�~Z���ỤT ��ͳ����v=�gd=��,VoV��Ŏ�<�{�=�R��4kQ��̽��j���0V��r\�ٳ�>��Һ{���J'WD��zy��eQ���Wj�<h~���Б�L�KH���~�=���d4Upj����pDBv����Ɗ4n���G
K�?R�(�`��V�E�c��쳒84d����A)�Ã�ۭ<M3m�v�4����aZ8%lk�e~5�I!��Z�SyxN;-��;n��v���n&v�+��/��;w�sl�ĳx��e��xs	�ky��c�n���͎�w��s�N&Ը�(�^�)i�[��\q��$î��u:�n�m����vi��ǭ��9��^�w^D�j�Mv�˽��0��|d�3L�.^�u냶5�I�5��L�|�/�ܻ�$�� R_9��8V��Mv�6I�rsL��:d��mR�Y��t��4Z܉a��V�L�X�une��7؁ ��W�ZF׻��kKAc	�)����4iBU���5Kf�����3Mf���Ԭ��RV:l���̣�L�����l�Mc]Lˆ�fΖ�󓼜f�D���B'�@.]@�K,��~_gњj�:xT��F��I?B}-�����tM
����u$v"m?)�"҄RSlp�������toe��bf��~\y�뗲x{�=gI���c����v:`������'K%'�+�UZ'B冄���˞ʻ�/����Xqe�dV�5E~>���ѱ
���TA�p����˥����%�S��uF���UU����K�z,{&�ގ<�j�=&�	�
�B�xf��V�e�`Sk4#�w�,����Ҭwl���iȄc\��J�����	�+~�SUQ�GɈj$�b�4�.hk�+�E�'M�O����q�I0면�N�ۦ���Hh�FJ���QPh)=���n,z�q�n1�ò�p
D�}�J�j�V!�5U!
��A��B f��ʤ��*�O�� ��C��r��2e����UP�9�I,�+��៥8�h�:M������^��{S(��[�*�i�X�[��� w����q<�<�n����:�]h�C,�(4"�g�C�hI��i%��,�ڗ�5�fil6^F�gg����8�I���{km�ָ<'w76�4Cwm�8�n�Xrn��L�7۶�Y��Jj���K�4j�����W��[��ph.� �h*�5ӚYh����?F��¨�@߬e����&#i)Ծ[���u�-kyO-����y��0�R�q���><�xj�{E�8|J:%pF��<	U�6T_�f:J$���ӢMz h��3�ӏ}�x���7��&v����!�N��O��"�����Ef�ò������	�,��G���7mg�j{'��n�F	���/�T��VLE%�˘l36f��y;��ez6fY���_�x��65V��hA,t���q�Dމ���:j�~�.��rۿb!]��)�H���Q��r�a�Im�#Qs4q&�G%���㌉<I�;[�5��#����"�ܱ���Z�m���W(�g��[EbpH	Ai`B�A~Wh�I�oj�n[L?���l����u��$��Si:�u�ZXa�Ma�t��&ྵ��cB2H�)UkM)V�3e�E�h�USEs��'�Um8'���dsfY��߻�}��x�I�l�Qd2����a���Α���)K
�!�<��=̫����1��.P[����Cͩd"Oɇ�(z-���Mp�ݜp�F��սӣƱ�˿�$��z��͞�2��*�𘛄)�%��3��O$Ĵ��(_��>j�����*��85WI[:w���$ޞwMk�<i�-�xqsndގ���&�=3N�g��l�W�>~iȇRI07�Ƒ��8�v����1�:��h���Wgf�=5����L�vY�n��M�xӽY��:o6ΜJLCID�ĥjSo��~~~[�8�$��Si:�u�Z|��㳳O����bM����.�ݝz�hΚ�fr���D� Hk��������\�2�K�:Ӭ&
�7V8-��%�5�vci�qӯ;k����7g� a!3���=�+
B�ٳQՋ�%E�֡,�.�i���K��4B'k�-�V�V E�.� ��G\Qkw��7WB�2���3*�1fqw@r���T�A�X�;=}k��5�{M�S6�TT(�t�D�Jݬ��BĺCz��^�t�#�ڢ&!ԊI.���q:��am�6����o[8�V!��0��eݚ?W(.�Ȱ8!v��"�iFG"�B��������h�N	
��m�nN�_wGD�����mn� ��׏���1#U�:Y*��?V����~Iqxj�YSA����(�X5F�c�At��E�]Cc*��7�b���֌̐��%]�u�nlç��;:�A�mj�ՖI��.�эQ��<�JΗEkX�t�p�7�g���'I���;&�ʪ��!����R_�u�����q��$��Si:�t��GłA4h�̽��_n7F���(��T4�>�{�e�R���Q�@���h���Twb����?6	��(3凓�;]=u�חL���yM{Y��J�,�~	ThCCA�G����N�j����!�4�]�����뭳�l��q7|���g��~����m�UƪP	�g����g��m'tXz��Jj� tMVB�V�k���dU�baԄuͺ�8���'!��.V72�p�$����,����Ј��MŗU�h��U�Wk�
<��a$��c���m���%��o��wu���H����t��s�nK|h���[��RY�U1m����~~~[���ŭ�[��y��1�T�l��&*~֦Z�;ywJ(��@xh6a���v�����Ղo*����J�B	��~�G���[���j������{%V��s��,G����w-������yN��8B��������խ�3	�LKY�^�X��;!�l��.�8&Ɗ�AU���|YH�%$�6�C�,����{���"��$K��EU��eѰJ�ETYd���%7A�~��pJN�B�T~�[×ws���64m/k~l���Ѣ�!�Uh�M�*4MSV ~��#$�U�8&��?J�!�WA/���6%?��^�ѶS�����q�ϒu��io-ǟ<�%N)��}:�L��o{��:>k��EPA��2�H�5GԝdI��Q�<��[�N����z�y����n`F�EY����Tp�Ǘ���[��K,v��:t޷�`EEYs,�V�&Ć��F� ���~�~]���J�2�J�$�2�բ�q#��w��@�C�`wd��������*s8M��swV��L�6~7T]Y�(?	���"g�m��-�n7��|�u�����D����~N��Yl��)�d�A�F���	�d��z�54����,���(X�h�%`�)�� }��u�2�6KI�6�bb*�x�_�~k��>b�'m?4��b��k�+Ʊja���lV1X�q��+��WX�|���m�c����c��1�N�cX���+1�KW�W�WS��k�mƱ�ı���V1\1X��+�V'���'�1汊�q�c�O䭊Ŀ??���|���iX�c�V<�'�K�q���=V'�+�*-8�OS��Ғ�K)be�������bq����w3���q��+�cX�������մ�q�ū�V1X�S��c�q�q8�T�Z�+i�J��<L�LR�8���'V1X��
J�V'�[O�>W�+L��Կ+�T��N�Ƽ�'cX�M�_:�1]M1X�|ƒ�X�c�W���מW�W���j�3J�b���1��8�m�bi�ı<b����u8��ɌqQ��<N'I�^O���e,L�R�b��N'g���|���c��jY ��ٿ߶gMq�~Q���}����X��Ӿ����q�����]w��w�����w��{�潽u��湕3c&�w���P�{�����lo�x�����O7{�@:Bj�&�O|�{���w˽#�_sZ۬�fv��g�k�9�H:�3z�\d���7to
��wû�~�oI������ϟ6��΁�&X��N\���yk��ٶ�@�(h�1�'s�j���|�Op���v֐Nw��5�������0�8��x��h�)ř|���3�c[3f�Yn�[b5�I���i׮o1�%�?Y����l�x��"Z�f1T٣.�B��w�q:�:���s~�3��ϷS�4:�^���j�5����l�����=��?#a�m|�| >E�-���,Ѩ,c}i�:OK"J��J݂{kN�m���II�,�N�6�n��0/jĔ����]V1����ңv͐�ºˋf]����/u-�m
������k�3��M��V}Vb[{[`�����yk��]�K2����p��7�'M�u�W�&rK�.͖��6P6��V��f&��]���Z��AqJn���Ե �u뻪��r#3Œe��5d��/C� J5�o�����ՙ���w����s���g�5����w����>�ٙ��ʼ��˿wٟ}����2��ϒu�>I�Si8�x�gM	ф>���'0�/��v���ح�5���u�s�͌�,�I�q�4lUK�v�����!4v&wj�6�t���q�ʋi%�a,�).sYn��7kq�.KP+�ٷ�6�&� ��ivXѴ�Pc*�(�CFjCnFi�Yv��`��m��+���U�����%x;5����6,ay�F�]��c-fЅ�򚌬���ҁ�e���C��G�u�Zb���,���]Jm0gm�Z��J6͡E����3S+j�!R�	m��ih��%��Gs)M�3a1w,��1�.�6�aZ�M2�-̹�;�$$'.��{X�6d�lS6y�5]b�M��I��3YA�`,�e��qs)ql�چ�-�Yf�av��y�/�6ShD�Є5�w��oj�[��ǅ�8A�����+Z$C��.�G�d9E ��Kn�:��ӳ��m��� �E#U����F:/��,�q��
j(��M�
%	�D�7��0���~, }HW�,��E�[9����Nl�s'Q�7���t���45`��WL�Sw.����;:e$�����;�d���A�(4	V|?W�����X��iu��J��,ZRXӳ�]5Q,N�PH'+U	��F��
!*됣��~���D(/���-ڳ���f�8�~�v7��9=�I�_'����u���N��I�R^|�h�8�b�\�#��L�"�8���o�7S����&�@��cT�i��rT��Zkn��<��ۺȓ�wݽ̺ �T��Ж&Y�i�.7r�U �v�YgaڅbQ���+��}�,�h��T=I�,j�<>���q�0��؟�9B4`�=4�,�Og���+p�[<hRO�ʑ� ��R�V-�avX�V(�7\MTM7#+.86��,h����T��LC%qH�MG���5H�0�~�O��]"]�4A��HtB='e�M�<-��q�$ދt}I*�����Zї%��E`�HA�FJ@���,���N6���u�ϟ']M��N�:h��Hh��$��#[Vڹ�E),M��*�%`4JC�Y+�\ �b4�����Tڎ&mH��3p(�1%A:'j�	A����<HCd�Z�=IE�)h�L1��5G�П�I������Mz�D|ӗM)y��f)��nLF2�㴬k�.��h������$�,��G�O�
x2�t�J�J�Q�,D�*��	�F	T�% {�.��%n�IFƃ��@A��!��t:Œ�	[�C�Ubn���,?RU�����V z���cT�������,@Aj<��4yQL�8�rm*��h�[~~[�<�1�<��[�X鳦����h�a��|˦n�H���V���"te+��5(�I+�Ҕ@B���e4���Gl&ţ���!���/�����a���ؤ����X��䞡�PY�E�e�?��[5Y[$:�8�Wa�I��~_"�yQ
$�����=�b;h�G�{�Nyl�v�MQ�?���!�㧇��D���ҕ	���i��3n���X��1xl�$h,�5F�hHAP�T�.����,(�Е:����N~_�VU~<~��W��
���v��5+ּ:"�[��b�y�1�[�|����M�4|X$4CFe��L��B�cҥ��\�e���9OZ2h�&�"���_+��a�;X��|��״�%�lhM- Pu���G Y�&EXdrY�`�Z�uq�آ��fٶ�Fnv�Ec�iuE�vC6����]Fۑ��e@Y��<�8�6l��!��d�:Mt)nV��4�QQ5˓k���x�@�%�#@~�!�i?�?1�D��D�ᆎJ�5�K+��I[��-Ah�~K=P�>i�$��C�\~��u-/2��K�h�d&��EX����T` "4%��ܨi+��NC�Uu��BtK;���lh��6��W�v�vk�>��MVإ����47�o���ސ�2f�VY�W1ђ̼����"�]v��k����!G��ş�zm^UY�W��d??���U)��������X�???<������>|�:���H�n���8���ok�Q�oi��<�JQ$�qP����-���h�K��H[z���0�>�vl�7e!`��I�W�g=�����j�Ut��\�f�������0��y�΂}@j}I���g�~�_��h�R�$�u��qm>$���
�S/����Дѭ�֦�#S\ɒd�e�����>4t釰�X �~%�j�?l���b�\�K��k��z�yMG��[nm�N"_i�L�O֒گ�u��έF�M���N���ϟ$���H�gM	0��z��c��)H!�K7R��`�u̺���+��\TC��q��nx�$�3?�'!�Y�K�}Vi;Ml�@C])(�J��r��6k\��,lK��b[uiLL�l;3a�4F�&����y�9�K~��9A[Eh�V��?N~d̹�Q��,�ɛp�K>�_���ƜZ|pC�;_�G�K������>?T�U����<Y+��+��1�4Ja�J��q�8�L��B�><�1��-מy�c�>b�Z�>y�4R�q�\�1ڝjm(�M�)H �9G�יּ-�����]���ƈ! ���A���hH"l		;�~`$���˖�8��D�Zd�c6��!2Fj�s��gL����A|$-^&�ԧ�ĒA��C(���;W�=��@�SY�C�:8~=��YZ0�@CF)������{Y$����k�A���
- �d=Fp�*�>!Ī� �?X�v�Hl !��Ρ�-��fꪩ�:��[�?-�n���c������8Ƌ,�����?�ͪ��A�1�{��ql�8�#ֳ��jҀk\�Y��f��ھ�,��GK�5m55�Zm]��k��\9�sf�G2��V&,�,v>�p��pvF=�R�-�m���#i.f��f`��1;hkb����KYNS-4�[ڇzV	���33'4�ɮ�Z�mJZ��~��Kq���l����7���~O���U�����uN�M��(�o���jX��5(�lDά���V��~$'
���'�|8l���;F�:uƛ��V
K3)�zj8s���@�K��0�㕤kg��X	�T���p�ivi�c��p�ͳt��n�~���S��P�JN���?���Q��S͸��?-�]y�c�1�<Şq��Jq�ݨ�^�f2��[{R�L86~{P���%֨�X ��Ϳ��.�a�VIe���)�ý�ܻ���?�]W��-)2������}jY��ĭ�Pp��X��g꺕|��N��À����d��x}H���j�[i�X�����k7)�����1�~5Va��)��gsU[h�^�����ƖK�Tw�g���Ϗ�>��`�<���x��_��gŞ%�����C�?8򞍥v�NmѲ�?c�����O��ckV1LiX��c��q�8�b���+�:�1Kb�ҾaX�b�kcX�uX�O[V-�i�c�u�bU���>O]V:Ʊ���+�uX�bX�c�5�8��bq���S�N158�7LV1OL����1���ʧ�jx��+���Ռ��c�a��)��q�3�a>b�8����2��4b�8�N��+�N>f��ū��u8�b��bq�k�b��������+��+�V4Ʊ������+Ii:1R�&X�R�8��V��c�)���iu��1X�q��ɔ���U��~N���gj���*��+�[ji]b�,b���1�1�bq>O�U�y�<�'�������R�jq�1�ǘ�4�'�+���T�X�S��|�'�1�1j���|���XO��+lVL�Ӊ�����t���GӦ^VlI�녳MJ~b�c]���K.��O&���+_-�����a�9��g^
$䣽���з;�=��k����k0$�ָ$yp	����'ngMm֢�L6Ɲ9n������7����ZsX�e�T���o3s��{��/j��U�}����}����j���~�{����}��j���~�{���d��Ϝ|�'�u�1�Z��X�yǜcEѣ��E)�xl��+[]�ɱ���Ґ�O��cVy���즥���x�_�1N8�e6}R����L��ܫܱ.9P�-�q�	ZY�+�5�A�ݷ6���%扏�f^v��Z\�Ё���Ul/�\����ˍۦh�)K��j ��D&Q�u�Slk�Ј���� ���ʂx��R�t���r�\,F��d%)^|��ǦG�8��矟�[�ο-�c�<ǘ��<�)N0�U��HH�1�f�.!��}�i�R��!zu
m��j�e'㕼�߿N[-�.H�̌��M��b[��]5.������F+9Eh�6Cz�bt�}\8"&��Ã�Q�?BFui��W�DDL6v|t�|���DN�T���K��!xv���n�W������F�aÛ��B��.����������[�)�����V��/ъ�2�47�-Iw��cl�����tl4""dK��B���:�mlbߖ�α�c�1�[y��cE)�0�w|���ý,�J���:���x9���]�=�g�#p瓥9�fM2RbI��l��뿛s|�6;�O$g���G	��׳V��
�	��l�*r��T�-6Υq�܏��@��!;�'|sUbA��QĴ�m�1m� Ź�$�]X��M4�+̍YiJdл:���»06a�*J
d�1��k��ٔl$�U�4r�"0؈���:��WvO�$��+b"$?*T��]_p�'+d ��r�#$��]�=�U���؈�C�V]�T�A;U��,������b"'����AS�����)���Tzh��c��	�q6�!��ܟ�&�5֭Țܫcbl8��X9֛/R[/M��a~S�y�r3�4�O)�&���n�Y�]II�䍎����	�����gż��b��-�b��m�A!�E��̻��lQA:'��m��u��3�:�&��A0�;��~���z�B ��+�d>�+d8|��ٙpƱ�c��8(�p�$:�A����+��?'ڙž$����D2PK��R�]���_�J$�o%3SyJ�U��k���ZMYn��k�f�|��뾪���r1�N�L.U�,���a��	�A���.����C?
<[05O��8|�ϟ�����1�c�1�[tæ�� �Ѣ�J���Sآ�WǬ�k�ѤW�AٳB!/Ȏ�ё��j��9���;�e�� ����3��u�?Ra��.8~9Y^�s����O��>%-l&�m�n%��!�,͛9+iN��ѳ+�l�
�_G�%�6�_�n�)�ճ��~�.��S��蕲��F�C�C���dk��L��Qǖ�5ٛ�ۇ�IM�&vg�Z
?��tD2¬��F5ey~��q���y1�1G�1��-�c�1lc�0�o6Ɣ�8�fr��]i@�TJl�
("\5N�Y%���r�?p�a���h���O@8�)Ԥ��T�53�%���̴��51�ܗ'6rb"diI�F��	u����d�tA�c����Ⓧܸ^4z�����,�Wd�{���h�K�֑*�R��B;1�:��w��0�,���|xy�����՛/���7vl�f��{�䶤/�p�,��C���B�	]�&V�J�3�ƍ�տ-��y矘�-�c�1���kiIS�5���\%��ۣYuk��Q�g���C�+���m`���hwl�	~�|׽wy�'v�yjT+5֓L���� V��5ȄѫayZFY��$!&Ä{�����F1�%kĪ���xC7i1c�KH]s3��
���s�]�f�VR�;:Y��˝��%�$��K($�T����l�V|x�G�o�ފ-˻��l���X���|j����W>�*�#5R��+�Æ ��X]h����������S\6!g�|�wG<~��� ��4��xԐ�h�z��th;�@Z�ZP"���gF����Ọ�Wq* n���YR�-pŉ%�xЙ��i�=��O{Ka�S�u�W㥈J�\\�Ͼ�Z4�}�O?8��~~[�<��1o1�b����[JJ�q�c'�37iH��,H�Z�HV)%1ߐH����{�d�w���b��$�ғc��U^�����,C��`�K,!���Pj2x~��	=j����m�8ڒpT5��S�g�T��j��a����Ǉ��\?W�t�b ��A:Ĺ�[��%��*#,��[pYh�S^X7h�Mb������a�(��֪HlЕ*,,���7$`��قAݜ��	��TQ���Dya	ڟ��M�/)�I�����n6q�1�����cc�c�1�6��Ғ�i3��$�
("��,�醹#:]t����
���F�N�w���v�"W�����e���`�BB'+{f���s�����K����"]�GZ)	l�m(�>�;�_.#M>�Ii%��O6��})���*������~�p�����X�j'�P�R\$���z:'��.�J�{�j�N� ���9]>��;��$׍�6/����y�1o<�1lZ��-�a����RT�-���2֯�6o9�EA�;�djl��ͪr�t�AN,�[�;-G�$K6��ʎT�X֔fh�α��i��%l����}�KQ��R[O��"m4�?~�;���k�p�lن"pN�i��P��~�<"���P��(������.�����4�&"����2φ?��l�u�^cm������%���f����1t6j�yM%&"?20��)O�Q�o�ϛe���]$���I6�I�M$��6�z�I&XM��e=e$�M�I<a$�I�q��L'x�I&�I$�M&I&�I$�z�'���I=u��I�I�I'�4��$�q�S�#6�I4�I��z�I$�	'��׍$�)$�OM4�,�I�ǈ�$�L���L'S/��1�1�i��K1LS�0�����h���'�$��K�u�]u�c�1,Zֵ�I�$�$�m=m2�e=mi�����0��S)57���~��xvt.l�p&�oz��wg������O�o{�˥�ݏۻK���٭>�F�i9��]�Tw����p|,���fS��õl��0�]�pu�^��9�<�i;���/���G�{t観k�sBI-{����O�N�^��6�<���=���������]�2�T��^�n/�|�e���F��m�3���s9��Ӹn�S��Mo�ךע_
t�~�<|O�sygl�������Ǽu�[h����;��{�����e&��{�hv����d���g��4��MI˼���dm�;��W�w�����/ζq~/�ė������@u�=�(�����Cw�`}��ԕ��n�.�5�Q��;0����!��� ޲�M��'��ܻ���e��7��b'<��{��$��{�����]1Au���77:�n���5L4i(�1�aU&\g[����]���uDN�m6Z�������m��T�&���@僚��� Xa�sJ�-�Q����aIsM�I������X]�[�=*Z��03}����ճ"�b��3�$��{ۄ�λ�Y�G�M�߷߼���Vj��^�������5Vj��^��������fe�����w�Ͼ�|�䱎��b�y�bص��[�[n���;;,?z_ŦX�])���uC$�f���Tən��)R���m�y\�xꘫ���K��JK�mmN]�ac^gC�!R�[b��.�Sm��j� �%�m�d.+K+]-��і�h����X����"K�j�2�*�jmYf*klh6m@%"YMG
�5P�5�M����E�؆��yl�q�&vαA�خ9�s�r[�gKX�4���1�qR�:�Ie��Yq�͵�Ի��$�G�-e�u-�t�Mj�Yb���j�bk�-����f�.�C0v5L���jf')V�vH�E�6�ӎ�b�����5�5�Y���	I}��-O9��n���XV����5�`w:ٙ���A���v���1�$[[L��q�=��䉎V��֮4Ac�"J8�Qe[�HY��y���-�i�T6��:����[�S�iI7�}�mߛ|�I2%�ڥ����r#H��MA��TCV&���d��!�YH� ���Xp�IM��,$���{ͥ'ѵC���2f[i�ZI�S�(�oE�99�V�,��[JR����$�7h���I'������l��x�lCBB�49Y�.7���6��c����c�-k[�1����)JqĲ3�.���rpQA�P�[��=�Á�K��y �ώ��/�X�"4}�ч��{��b��6!�Vr�2�~^��� �kg(��ܱ�.�~n˗g�6}�< p��t�n�n��<y��ۼK�VйH��y�B��[�km�.�	g�㥟6|oGx�І�YVYxh4q���~<0h(h��p���dUj��r��V;|u������u�[�1�[���1�c�m�JR�q�������7�,힭�jֵ_��[0A,6Y�8a�zH�І�!�Ѫ�N�y]��.jL�kW�k����l��r���?kc�a�D,��pъX�B٩%��%8�6��3.K�'N�%{�����Gj��Âp�SZ9̕���1˓�]��>N�Y(�v�|95G3�}��pޫ��7���B�K���~L��g����+@�}��|�T ����B�Oʐ],���N�kt���Y��g��K���c��b��1ky�c��|Ҕ�U��L������JK��آ�!�{�ի�U�FW6l�WkAb�j�|�?:]p_óE��`�?s�\�ZE9f�-$,���-1��H�;u��a���C>O���v5���F���qp؇�¨+d��Hgdg(���˻��"h�X��Ύ�R�tjVƑ��r)��~��tk�Qb	���P6�툵�F����f���т"�s_�	��Ąr�����|tIJ�lD9��6s9E-h�UY֛K�1�:�-�ŭ�b����1Ÿ�JR�q��;��o��rJZ��zJP�h���f�H3Y��^Gnq�����d;{��l�&��%��Xp0\|�#�s�L��D�<^q'��gCU��v��jͩ]�GCm�$H�����1�>�Bޠv�j��5�X:]b�!m�tfx��Z�)c][4�-��X���m�Me6����V��b\���r�t͠@���Å���!��Y����w7��w�y))i���kLu�>�<�K���%����etk�0����ц�ֺ:8h�)e���n�Vn�_�����ΏH�����|�-��IJa�T�)9���{���s��33P����q`��6C),yYZ0��Cf�hiQ(���BV��$�]<�>|�ļǖ�X�y�Z��1o-lc[�4�)��U3��5�k���p���F�	�u1��L�91ľe����AZ����K��c�؈M�æ&�b]�Ca(��#_�0��I���%'��������CN�I��^��⍖�˳��t��A4k����J���s�9V]Ye� ��E;2�}��1�������ƒ��O[m%�j6����M5�Mj4��Ҫ�L˱ݱ.��1�T�[c�c�y�<�-lc���1�-�R���FK�{T��(��l�pC���L���b#��tv6�S��C�&F&)�},i���F�!�D5����ʳG�.�B��͍����v��75�hh�����<�9��(���Z�>4�5H�!!�nF6~=�����ɣ>h�?`X����K ��+Afj���i�,���\��>�Y��V���=G����%J⥈��+��NY	��[α�<����b�Z��8xѢ�B4dӗu4(��t�0�V�h��U���uճ���'������sw0�ޝ��ַ9��a%�T�Ck�6&���|�V��3C��~:Y������&�ӊ���g���	��s�l�wr��:k�`X��T,ÿ.��D�C[0�/�r7{��"Z/�,����]�fޒ��j�s?=4��Y�h�:���ڟ��󮱋bص��bֵ��qn8Ҕ�w�MO�.�ت���e0��t!�c�9u���Ft�s<��+7������y�8H B0�7����i�7�Ԃ���)u@�RVjJ5�p�@��i۵��n�u��n���X�<��ڍ��4F9��tBlM��'G��o��n��D�f�IWc�v.ԷSY����1+Ķ�Km�c��M��J�]^.��G.t���i^5%,Q��;ff�C�����.�á A2�>�i��zi�y2�Ĳ���-��p���tR��~�,O��(�0 ���Ώ̌n��'zW����_�C��EN2B/�a�t���_BeCb~�'�lB� �l�[R��s@���,�hf��3!�1-]nu�K�q7�K|�6i'ʔ�]�}�E*��L��U��U->|�[�y�[�1lbֶ1�-�R�ѣ�+q@�QU��k+���ș%�j�[�&�d�̖��$A�ALmй��)H��FV?�"���$%quq�ex�0�'�f�%�,٪7Ӌǜj�Y_UU�y)�y���_��8A��~?V������F�$��'�>������&g��J�fC�cK�K͕�����9$����������ψG���Ԗ��~q1��%�Û[��&��#F��91ϙ�QS3�Oɧ�:�y~��:�N<p��z��I��I��ORi$�I8���I2�L'S	��u6��M��8�m��L&�H�I$�I6�O)$�I$�x���[u:뉖�$�M$�(�ORi'I8�m�O�"L$�N0�L��I$���x��x��<I$�ORi��eO<DOSĞ�x�x��q�i�%�iK<c�kmo�M�>|�>u��q����M�k|ǞyN��]u�c��-$�p�	��I��8ˉ�z�6�/S�I��2�i?�&ΐ���}���.c���h9/U���q�M�I6&��p׵�w��D������#4Oe�����f���$�]bs<dyN�Ǚ��m�J�/R9ķz������{�w�Z�y��ӽx�˜޵�=��j�wm��r�|�`rON<LrK�/y{��Ms=�z�j�5e��$�#S.���C�]!�ʻ��SN���?~�{-����!)�r��m:k#2m$����[pOn���b�W��oIw�.<{_7���X�Jr޺q���7��������f�w�y�ߥs[���0���8oX�}����r��{�׽����>�������ڪ�]����������ڪ�]���_�m��>b�ŭ�X��-lb�ŭlc[�4�)��y�'�(�"?�GǍş������W6�4�d�1�ۙ�*8�N����g�?��6J%��)~|�2Q"u��e�i�:����e��`²�-�%�8ⱇ�~��b�9F��`A�x�r��/'�3[4v�H��Qf�߮I��6B�v���'4l�(���z�ܫ����E���]�r���DʕE�hj�R~>8~S���u�矘�-lb�ŭlc[�4�)�DEJO9)��$���k�h�"�
C���hڵ(���0�&����Ϸ�-��%�L/5R2�h���V��b�\<�]���mI�5\*>�*��A�"%�,�~��)U	P�g�9ƣF��DD~�LO�)��a��4�SF	�>��IVe܌N�����]�������a��"�O��6�!D�'�W�Q�Ԕ�矔ŭn��űkcc���Ə4YCF��ad���-��-6�V5�g��n�_A�d��@�S)���л��&�|�;AyŅ�ƅٖ'f��B��J:�O6-���� r����5�ns�9p�n�� �if �-5�͚�(ݝ(mMk�nq���]�[��MnƳKq���嚸���5�7F>�)�0�~"&�W�w��r����U�,,M����ѣ�5ыk���]�y�Z�t�,�E1p��9Z����~����MR�:�˦�i8�=���L��fTm�S2_��YPHh����5�¬K:Ο�>��]�[���Ҙ%\n`����C�fU4ߋY���֗�jωWF��X"pN� �.���y3���M����뮿1�b��<�-kc��q�)N8�ײ;�QhD!��Ѣ�t� "Xu*�*B�4~��>^a�'>�~d�
�:�$x:4#�dcP�i0 �7VX�i!f��>4�"<�v,�vI>;E�p,0.0�<Y`B}��#<�{n��[Lt�5�+ 
�lFj�X�ka��_���,��L�<Y ���hC���7F�'	*W[kr[��*��0O��0iNW+�d -o��񣇪��m"7�ܙ��:��Kc��κ��-�[����b�8┥4h�dh<d�Z���Љ�k+fT.��eJX��&T>�ŝ;X]yB��:M^��$4l�z,��5d9V\V�%�3���<���k�E���jY�m&fS��.�t��x�t�����hA:����.�U6l�%�P�A8iQ�"��Ͼ���j:�iJD��KT5Y����B�wDAEL�.�l�C�0�������ŭ�]c�-lc�bֶ1�|h�B4}G}
R$��E�|�����,�4�b-�K�6R'��5X�ĢA:`��k�,BJ�1|���:f��E��]��U���u����hd,5�Va���0����`��v�th�Y�&��Y�N�ĳ�~��R`X�!���_����X��S����Q)f�&���|��%.���٢�&T<YʳE�8'����-o�:��1kcc���[�R��_&�5�^�ާ�VMw�写��"d����,c�z�h�H�I�L�;�g�78�gw�p$��M�����e#A��1����q9����_H�v�7\[�,�6u��2��&�Pf�����EuF+Ojϱ!	�5�`7Tb,ؚ�6������&�Mvdغ�\M\3dk\�l\1�sR�p��Ի0���]��f[�m�.r��bp��i�..���B�,�_z-������>��}Ek�2'+�bo�z%����$���;�Fܩ'�l�RJaK�O}3�h��cx�2-�����,D�U4B˫�����H3�5�\�n&����6��ۚ����ʇM'1t�~��'%��LUT��i���Zc�lc�1�1�[žq�!hѿ��N����E�K�ptz�a�
�6p��hپyI"IuS^�d��>Z�btm/9M%��M�{�cs�ÅX�!5��ń(�ߕ��V�[.	���Y����N�����<t$"D��#	D�\D@I��a�w[c�yY+慶�5���W7�\�	�e����x��_WƎ���r.��a�ń������������֜g;�۩y��1�^~cO�y�]Z��-lc�c�1�|Ѣ�4h�Zm��{E�H'D�������&���%]���/2���v}u��>�C�G�dٲ�V�0�8Y��v�F��U,��Z䷝�0W��]B�١���ƣ0�r9�n����>�ǎ�����-Ֆp�_꾲:[0��	��t��镆�UU���.�v71Z~��-UM<�'�ۭ����*�4z񓶳
�h�Y�W�:p��u֘��u�-lb��<�1�c��8�)N8�L��5ߦ����]ohNv�E�;]!�+7w%������x�͐|:0O�,�ݛ������3�FJs���]3�٥��nGMy��GR�9��7?���FK_�	_�M��I�2��m���p��#�~O��?l�%�] ����\�yr��[6}V|a���0������F`�'�k�g�07�%Nb�k����컗�˼�W��,�z�y�[8��#R�%�����,>z���I6�I2�i'�8�Ēu0��'�$�ԘM���<N�ORI����N8�ԒD�I=I$�I㩄�OI$�I$�6�N�۩:��I$�I=I��)4�N=I8�m�DL�����&�$�$�$�N"I�ǈ�I0�I$���M2�$�<x��	=x�ǩ����6��1�|�6��qe�屏6�K������<�:���cZֵ��&	&�oq�����2�?D�OS)4o������f�M.�3Q�V7�i��{�I�j�<�������"�6=�ڝ��ӵ����u{�*����������X���Z�}n���y��g~��w)g��w��õ��-An�ͻOc��Χ�}�o2�9�~��ަ�=�k�r�����o7�����x4�[O�D���Y6n���~�ԏ�>����޳����zO;������[�C�h�V�ݩ/ox���=z��wg�z�߽}�,�_���F~�cm��o�/��>>�����ǿK4���f�w�z�2sD����M�"�ٯ/m�Ĭp]e -�M?
w���;eë�b^#eK ��r����w�{��Ѵ�M۽�n3�2u��6�`��!}�KC��s�}��|s������>[7���R�W�aQ�)(�;���>��t��N��P	��[��l����*t4~�M�|��=}�{�+���;T'�Q]l�;6�nM��1�8Z�hshK���Me�t�����o�z����iiU4��a�2Aik��a0�]2\5��u���ۃ�&eu!�e֚�X��J]u�֭�l9�,�vm����i�0�Ƚ~1�/V�\r��F�Jm��iL�����H]�W!�~�ͷUU�j���;^����w�{�;�s3;�Wwun�����־��}��Un�����֙e��y�]bֶ-lc�c�>><lѢ�4h���f�ZɍL�&�P�Fj�R5E���p����-k����
�[�����m6� E���YtVd�6\�j�+n������V�XU�s,Qk�+u��L�k�j�����Ѷ��杤\j���j��9�\6���,e.v�0@Ў)/6C0R�5D�V͉��&�ظ��jr�r�L�L�5u�ػ��\K�����t���5��%�!v���1]�Κ��Y���m���K,��#`[1T�n=�Knj���cl1�ͳ�EZPa.lv�Gh��*�ҡt���S�j�㆚f3b�j��!,�9Ѷ�R�-�`�cr��7[�lq�K�B7klFX�i��"�4�6�Ky�il�0UÖ-J�ݍ�	TY���irBH;\,�5���(h�el��,��bl�K��	Z!/j�W��2/�w/�|}F�VV���x�~T4gk9rHl�l�C)M�h�Jq.+���GD�(TY�°�ިC���7s/$���K��`�N�������G��l|Y�����EQЛ0�|�4�y�X���[��1lb�8ڔ�8⑺���a3V��v�����jl��[q(�墋Bz�~�.�5�.T��7�yUd�m~T��6z�C��ˬ!P���L�|v����o�܅��:˲p�F��v���n�L�~p��~;�D��h��1�i$�?���h1��u���p޵��#�vb�X!Ԏ�.x[���g��O'O��h��v~9�?��w�7���x�@�)+e'~,�-j�?Sp���fvۊO#�jK丷���κ����kcc�-�[�R��F�Up�#QH���(�$���&6l����yl�K~�[6tXY���KZ�.(��?[�?s{��s���4(&f���4Y����YP�W{|3a���K��&��ٮ-n&�DeRR%��p���ϓ�҇KҦ�?X�U�>�j��i��Y�r�J��/��١���~�0��v=,�4$�c�F�p�`�C�}�`��^��[n�������q�$�gNRg��K��cO�~y�X������1�[�-�J!�G�̒�
4��QhCWk�{���YJhф:!b"~�]@g��?6�%���05�:�U�x��CU��!�b�5�.����3�q�(��~i�#�4�h�Я�:Xh�9G����������V��>p��R[���]�Vj�,7��2w�Ҷt
�&W�X"a���X~���X�+���JNWz�Y�?C'nܧ>��m$�-/����^[κ�����<�1lc��6��Y�ٿ~�BV<
��]^Z�����������|㧞H��e�R�i+�&��e�cK�iw5JSGcj���ؑ����3'���gO;8@���f�LA�u��y`aP�1����ܥ�U˚�l�s�NmX�m+J�嘶Z&&�i���f�J<w���C��1*��9캀X�6Y���G�ǆ�!�x���Ə�^5U�ԗN�v�+�$I^E��蝤�j��Õʅ�?T���kI$�$�ȐÕ����~5Rϭ�Hd�h �	���τ;?	�沴���ɋ���K
fh��� �+xJ�T(�o�i��F~��D�B�4m��+���f~l�����mlmly�X�V��cc�1l[�R��nQ�(�`����E� ��|B� J���gH~�%IX*�[%CT�0�D!��v��T��h���?J�УTl�W�~2�h�����[ȴa�����h1��\,龘V��_����e̓��2F�"Y3-��j4�%��\U'h��T{ʫ�`�a��ς��a
Ø�L�O�;��ս������02+��c�e��u��q������X�-�y�|�jR���T��m{Y��	�������h���L:	����`p�T��]��B�8k���ep��zG��%��fBbI��G`AF��x@;?{��NW)0D!��N��DDD�]��?IOߦx�&)�Ξb!Os��n�G�!��ʫةZ.���?J���V]�~�]�k��E?SM%�X�Z�u�-ռ��ǘ�-�y�|�jR��Dwڞj�f��Tꇍw��K����{�Gmb;*�~)9��U�tg�Z��]7m��c��l�4�&��.ګ���R#�gy���,y��(������6^5m���m�D�g��X'O�Րk�??WžӝO%�u��mv2�bv�ύ����N�����P��N��v7��5���g3�E�*h��*|����|��y����ǝu�uo<���1�cb�8ڔ�8�r1��wfX~ݦ�ӝ{�g�����:c�����'I�l��c��6�X�^�w*J�&�v� &����{��[_x��<�s�\hO.��'z�e��ءY�.��A��Eѡaf�Kn4�I�Zq�;� ��u�k�k H��t�ݨ�gS.Lݮ�+-��(f�� ���n��x�59V°�Eֱ�"�XY��.V36	?G���ŕd�t���i�EaӦ�B����U�|x��*��f��ۯ�˻5D��4�_��ң�T�(
F����T~��l�z�#Æ��l\\]�ǝ�%.G��K>�V����F�Z5����ÇC�����[���])��,�QVѵj�
E!ww,�ܨ��/h�$��j�ڡ����]��Lhӏ8�θ�뮿-��ykc�c�:��m�4h��ʐ�H�u�L�Z��u8��>Z�n?C~�o��%�&4J�+�������i��i���x"y�Yy������=襛0J��8U���,�~��r��Fm�+S6:ؓ0��.�6k1-��K���p0��KJ,*���=�������:]h��<F�V�������Sp���m�J��9��浶�<'�:���>2�I=i6�)��N0��<I$�8��I'�&ޤ�M��OI6����^6�I��I�IԒN�u6�'I�I$���]u�]u:�I=I&Rx�x�)6�n0�q����$�-�I�I=I$�I���x�$�I$�e4�M2�&��z���ׯI�e�z�q���z���>|��Yi�a:��QI��1�u�|��y�y�_:�1�0���I#$���M&�$�.'�뉶e�~�0�٧��vy>�-��f2t�[����_�t�M�|/����e}w��-��g��1g���^�Qf{��jj�/P��57�s5���ײ�̂��7�٤SہĒ����u��5=���mm<�$���[|҅�[m��WMI���+�2�w���s�}s���K��{g|�U��{��k[�fe��e�����c>�9��웻���߽�g��m�cq�]u�|��Z��ű��Ÿ�JR�q���32J��ө�u:z!옞>p�r%�s��8p6B��2���Nܗ2�������ѳ���r����\�oP¢���=J͊�2n��.��G�x!g�l�g��w豣�E���!G�Q�X4�[?%|�,�2��՝���=Xe~�+:h���HY��g����Cy#fV1X��f��K!��G���<��[��ž[�-ly�b��X��m�)N8�jO�2�em�mMɚ�)��z��#�(�}>�gи�����'�$�\����gN���e���Zb���
�6��MS!Z(caln�!3$̅Ŷ�{V�Q���fN�q��R:�U��aߪ���J���%�j�0l�������Xn�(��ԯ2�/�gJ�Q+�,�A.�Yf�[>W�3H�>%�*�F�K!��lU�)��4m��|�O�8�&Ӯ�����[��-��R�㏗/�W��Z�^Zmcm� �ca*�	�.�췀i�M��kHaf�>gh��9��ʑ��E��:�4e��]���[(V0����6������ͽ� ��t�kZy�i)�.�r�[t��V]����-�W��k���f��ZBQ��g6��n\0��iv�.f��u�3+����������iߥ���}�FmN��G�r�X%�%���ٯ��dEDT>�^y��\S[vS�nľ,6x+�߆�	��6BW�T��H�=v�,��6}�I>0�&b��=]�8wEJ��ܑ���E���]��ь���x:�m��]�ї�Qm�Bv���bl�&�z��k{�Z�s�_h�:��:�[�����-�|��m)Jq�C�T��(yO�k)CTU���$��p������tG�$C��N���]/�-g����e��G��F�Kf�(��ߓ-�nI�%J�>��G*��|R�p5V�����YʽS?���ˊ.S�ŻM�+m��D��F��o.F��Y�z��T�|��(HJFU�l�Y>п��N�Ɔ�W�0Ox����|~��-�֓3)���)�L)�M���u�V��y��1�[��-��R�ѣ*M�@E��*��I�yճ�Ԍ����G�J�V4����_\�pK�V5^6=d'�z�Y�B��u���Nj��ń%���֮eά+Zi�9��[�����0�����mx7S�(�p%PyZTOv�������fC�K��uq�c�	ar��߹[}{Ց���I8@OT!ӈ�0����q�S�q�&Ӯ���ϟ&1�[���)��욈�\�Ojg���@		��K'a�g���qY��.�.V��j�Vh;Ug0��'jz���F�>�S��ˍ�.�̕�e�8ÛN4G;N�%�M4����,0���h�ރV%���&��5�>!���iJZ�ts��҆�d���M|��x�o��%�g��b,�Lp�P�J�XX&	�G�GA�N�t����~����q>|�n8���uԷV�1lc�qn6Ҕ�#���QU[gf�����+���ߛ;�v��<AKO����ēi�[BMj���3��l�[g-��m���t��M�Q�M�ՠYf1V��B��;%���Gh�k/�!:޲�K�mVXV.�)�st��]Y�affj2�V�4��gj��f��R�]�/H�x虥%�M+1\k1����K�K��õ�c�,�'N�a�=S���0�}�[y�5�~>��Aq�ҵ��tm¡��(��6Љ���C�|��.����V��'�\.�Nl�v�}�0���8U���6~��*�	��g;�U7��������j�qZZ�ʥ�:'S5_Q����S޺��̲߱��%�P�ܺ�YN��Ə�N�6�$�uԜI?��篚M2YCE��&���t��k��}%��Ct�,�EhB��Y��~a$n�r��l�ڇM��C��^1�b�����e�����<�"�E���म��~WM�@h�oJ�3>n)1$0�2�$�5y4��r�"4�`�D5�����Y�/8�t�A����B5��|I��d�.͟�8t�������,NY��,�O�.Q�E�t?�g�:y��q�ɤ�8�u���4�YCF��|�:�;������ �o��[�֟FC�4�HY�l�a�l��Z�ˏ�����J��]G)\ԓ������W��o���cP��L&��ܦXEz0�G7Bp�X~;R�|\�8��ffbC�F��W��X�� F�����b�h��[ �;�K��h����xzl��ˣ)+��:/.4�ޚ��S򺜕%��y�cϝu��4�u'N�Ϙ|�i��CG�hQQcC�0���Tz>�z�w~���o���ǂ�kg���O+\֐*�S��Y��sAXYW,,Ia�����4ɗ����[w���?W�Չ��cBm�{����~�9�[��eB��M�V�FΖ@,�M��um���h���NϛLcx�[w,t��$�B��G�%����mik�K<h!�auzV����MӬ�a�^��i$�M�Rm���"I"I$IĞ"I=I6�I��	��$��m�Ӊ�	$�Ē$�I$�a$�ĜL'�8�m�\N�ˮ��$�I��OOe&�q�IƓl""L$�m$�M�I4�i�I��z��ԒL��i$�,��i�L$���D��׏I�x�0�$��I��ξi�i�ϟ<I8���Ēm&�,y/<�θ�cc�1kuiפ���m6�OZu�����Oa?D�I�)4��;�>���f�0N˼f���M;<���Git�D�:9�O��r�׽�6{��k�_/&���y��v������=<����=#�ܠ�UI�i�#獽u�Y�wv��3�p|g���wu�s0�Y"�ol��Me�܂���=��F�9�������w�GfG9����kLt��%�����5f��5�oo.q�욕�&)�� lD��m���
/����͛k�c^�߯r����^��O;��=�������Iэ�^�f�c[��\7�����y{�Q�[u.�Y��'K�{��g.���!3h�Ϧo�'#���a��oTH��w�U�;���OV�h����:�)�=��?}���;ݳ��|�g{�/+{t{���Y��H9��o:��ݯn؅�ia0ܴP������)�;�|�����{��{�6�g�<_u'>)��ѱ���鹝���G���y7��C�Ĵ.�y���ϓ��,3�j�ce��%
�&�eCD[J��m�^<U�Ԙ�����i�ĳ5�Pf�X2�mP��Ƅ`
G��/a{K5a���jB�QЄu�k��^˛�Z{Ǖ���'-�XYN$��v��$!e��{.4i��:L4m��Hv�Ka�s�=X��yv;ۨK��Lm����G0�����{�<����{���c>�9�����������}�o����̻�������9���q�c��]u�qo<����屉c�q���8�����[v�T�CWG-ط3lGkG:7A[@,q[��p��C^[B�.k���Ա-��^,��CCdw-m�3��]�5�ۄ��T�&�����9�h"XL�9��ecJ�g�Kfx�Yf��P4Ұ�6�R7Yn�h���Gg]l	[[1��4M��.)�v�	�B4���ҀiFct6��5�J�Z*]U������H�7fT�L�c�t`�R��V��e����:X�F���̖g����id4e\�͚h	i�Ķ�s�]��\ض'1�h�4���3�e:4���4���9���| HJ�{BKX���:cR�`h�%ֹ=Rt;/^hjk���y[��R�1%�^ՙ��cL�LV훹���Ze�XV�d�VoJK�񎻼���>x���ٟ��k\��5m�_���Ѳ4Ctg�Çܔ���_*6���1ȷn����ʦ�ʊ��6~�j����黻��tk><���َbi[*?8���*;�R�2��T� d�)WQXXM�1�[�
�xq���d�6�o�2�SU1�r8��6�1�-��q�ɔ�8�u>|�摣!h�Ƞ�*�6֛j@��4�(�kPL��8j�ՒjƷ^Q���NC�������<z��*�]ivyQ����K�LE5���4��g���뢰﩯��J�$�LF�d�1E�Ϋ�6=�������a�V���r�wk�:q�6q�S����DL�)��eW�3I�m[j��v)���q�:��q���uԜI:���>i��7�(y������ﺋ4F*��z<Rخ�>��_#N���������)q�b^i<\_9�ߵ�����a��(0�j��ZK�L6}�p���Y���E���᪳aad�P��G�]��|ҲR�_��l���>�.��WM~NHH�HǛS��j��п��̌���Rx���n�\q�&S���I����|h�aa�Oai5�T�2��r�]��d��8��aQ>�õY�lͧ��~VA���R�K��lanyt���69�ٲ㋇�V��BNCe�~6 {�jCC_[Tm*�#ѳ��=_vq-���˻���ú��p�'����}�'+�gN�j�Q9�4����L^E��]h��X���Zԑ�8/�z{O7�Zo�\S�-���L�]Iē���4�^<���D���`E��ݨ����\T���{^�k��.��䕑�b����zޯc�X�F겶�M	�F�e���MA[��Ѱ��	���� HM۬��)kQv1����n�����^f���K��f���S%Ҵ5�9��6�b��5��35�v3l��F&[˦�
�Q����^����t�ߏ�2H�d�v�h�tn��c_�ׅ����G�s3�N�Nt�K�;q4'�e�%�	��I�L�q��m��S[�d��!�����th�a�V��ѧ�(U�E�e�y�1�pfj�2k�C:VM�m���I�K�a��gM�p�o�Ga�z�L�8��U[����6�n?:�8�2�u'N�ϟ<4"a`x�䥽iUN֍�G��%�+��h��F����2[P�h���tY�,�������ϋ����<�4(��:pڧ�)6,�'�����e��]4B�,�Fn���7Jm2W͙0��,�̅���2��#V�yvp�#��Y�O�L���]G5�Ij�$*��r�Z����%)�q)����u��&&m�柜�K�1��<����u��I:�>|�e�Λ��J^������#Z��&�\���}�;<(x�IXYؿ!L=رd��\�-}D2�0��F��Ag�������$��a��#H��p�2�G	+�ƃg��NyK]�����
�˒BO�G�{%W5�kCE��D���-��׋�t���&�
�UAg>*��P�@��^�ss��V�*<��4�Ⱦ6�ߞZߞu�I�면�u>|��L0ʔ�Ѓ�=(z����J�SUY�*���k��#(��z����	Ap�W�m���=l�[;:�\�4��'N��mkŮ�
��l��S��o��uu��:!g"�|~uϾ�RK��/��/���_�/��&�e4�F�7>4,M�+��aۻ�?�&ɳu�xt�j���V�����Im˶��F���j[d#P�b�������qĞ�]M�������&�Y���=���7wsC�c:l^U�|��Է�e�4t�Φ;;�M�i���źQ��.!B���k);Gۙ����h�f#��&��o5�7� s����+SŹ֠C(@����1�٦��M�mK5�i��H�Y��Kev�њcDM�x�js]�u�m��JQ��2˨�����2��$�f��)k��8vFN�*�_��=k�U��Y��<$.~��Iw{4Hr�G�C�1�Z���	zӷ���ĿsR��]��h�v�@h���æ��9Aፒ��4�K���p�.�]�V���ɇ�\���7fQ�},�O����1��������p�o�yw��cjS�X��u�io<��Z����)ĥ�)�vg��UEZK�w�T�h�f��cw�%�^�s]�ç�jr����j����O���i-=rI���$6]f��h=��}X|�~������+�}6�u3�&��~���	f�7S7}�'W��7�3X�m�6-V3B�hdF6%}�M�=�r�^�f|�v�-�=�TZ���j�����Ag����N�;::�כ�d��確Ɲ[��~i�q$�$�a$�x�L��&�I�<D��RM�Rq6�m$�I�8�i�OI$�'S	$�I&RL��a&�I�i:��]q��I$����I�L��N8I8�m�DI��M��)$�i$�i'\Oe���I��M$�e��M=I��<aa'��׉$�6�=a�M�x�a>u�O�m>|��Ԝx���$�N�>u�]u��c�b���m�c�:��k[d�M��#.&S��m<e�B'�	�Ş4xѓTs�[K﵊�p�߰����6����e�q��js�u�姧=/����N>�<gt��v^�2�]G"f��W�y�rv�}պyd�<��ą��s-'*��^泼��s�/����6�ަ��3=�gZ軇[��pԜ7�&�k7����}�m'��nr���[h�@�ZW�6��[�C��Q��3��M�njq��a��ă��S<���s{�+[�z�ywww�{ٓ�s�����{߾Ƶ�}��}��{߾Ƶ��i�O�>u�q���u��I:x���0L.��P���<i{���MW����͂j������UHl��|o����_�f��S���v�Pn6vZ�l�6[�ZC]�Ś�O��K�;�y���W���'�hr
&	m6XY��ph��\>�,����*%˸��jk��ž�?S���3�L�v'M2y���k��{��[un�Ǟy�]q'��Si$�O�0�2�%���rLګA}��Fa���6p���������L���jڼ�a
cl'�t��h٭-�U4����y�w���R�)2���UV-�ޘ�Џ�GR�n�~��{���X�B$�_Up7��ʔ'qvg�~e˹DH�{G���~7_��\���S���8Rb־'M4����|�8�OS���I$��M�0��ϙ�D�rE��jKN��^h^���V����9�~n�Q�y��^�Y�g\�n��I�۽6�n�qNRr��]��7�a�#���x�,���h�[� $:pΕ`ʔ�㬭�@���yj�ib��ј�cn/+�at�`Lڹ΋v��j��(1�u�Wiv�1���U�a���,���g��U��06���LA��Q��NWj��ř�_��	b��L{$�X�l�B?{���C�F6�F<���C�5�T��.���.T�g7,cw}'6ƹ2�F=��k�Zҕ�-w]Ni`�YS1�9�L��Y����v�A�B��(Pf��~,�C�Y\y�2e�k��U�4|a��'\q�'��Si$�|���MB�}����AE�7�V�,Yq�D*	��7j�}P��pt����8kỲƴ8}O�%eh��+(�yh�ri�Sz��5N=(�MU��+z9��G\]�p��O�2C�����|�9�a��+�~�d\��&�:Á��1c4�B���d�p�uQ����k��93Se���'ї�U|��sc���f���S2�)���-�<��q��면�I?��i�h�p���zz�P��?~!_������w��v!����~<%�J��5qn[:�4wG��[��=��g*����P��ٮ-����!�|�<�̘����ZkShQ͡(v(f�����J�=��}�R\�,�Ŗr�~8��%�65���+��7P��|�2��l�ץ��F坑�6#��8��]�l6J��a�}$�/1L˼����,���4���㭥�[ǝu�Z�󩴒I>|�L0�/��;� �e�,+�(�#D�U9j�eB	���Ɛ��~��(��Ĳ�y�Y+�:Iv���Rj�ix��Z�Ԕ�l.��Gګ;H����F����7Ł:�[5����W�a����&��'�g�l0�l�6���D>�i�m�y����W!~��~06a	ʮk���7s.���g�D|�h�$n��뇒��q��8ۏ��면�I'ω�F���0���wv[�ո��%��_��u��{��yc��⎥�t�w����'kSZMk�a�3Z͝�ff�ͮ	r��mM5�2\f���[��J����D�*�B&��TyHjkv��\LJ1��pf&����ml�ΰy�.J ��@iu�����,4ךl�6�BE�:O9g��y7�U hHa|V���|v�h�N�Y]'�|h7�++����S����WQ����,�Wu�Tk<;	U��������qw��j��Ca�a��fRo�؛��`��(��F�,,�ٵ�T��K"W�u�8�%�\f2�i;.��S�P�������cFЍ�`h����8�e����:㍸�<N��Iխkc�)q�4�/z�sF�Q)�ET�Wu�>4kB���ے]�Z2�d������~���j]��O��5���Il�8���ߧ�U\�~%�(�bH}���ZFvG�C�C�ZCD�]�V��`�u��n$��G"rf�G��k�t�����F���Õ�`j��������o��9�}�E��>mo�:�6���:�m'RI�|�b&�,�a�;d���,����#G��Z�@~�e��I�V"%�Do�UCgŖ4|A�Y��.]�s;�y�l��:_��i7T�`k��x��Jdp�Ǵsu�ܓ����-��2�������h�J�ȴ�m��/5#��]ޏ,z�;.� $�`��i�-%p�H�~�����O��8b]VO�lg5i$v1&~�S�K�Lˁل�0C��8tL �ϗgk^h�J=ԓC����C��\>6����~u�<��u�j[�-���ֵ�1/��i��ɘ��sUM���j� �lV�V�/p a�c6�<j��v��Wke!0��������po#���iy��[�^@f�W(�*���]�T�?p����#�H{2�:W/F��6~��lA,F�D�n�k/t~�����a��$�*�O��V��p��s&M���A.I���Q󝸭��N���m�Ÿi+�|��oE���3�}a���w�iK+�*���lٛ8��?����ގ����ݷN��qm���F�o;'v�On�{gZw��]w�l�وzx�gZ",���DE��ȑ4M�#Ӈh�m"Ȉ�D�h��"�DY�"E�DM[h�h�"-",�m�D�"E�H��ؑh����d[[iDD�"E��Ȉ�,DDE�M[i�"Ȉ�,��"ȋ6��mD�mm�"-�h�,�h��"�B-�""�"",���m"Ȉ��"&�5��""-�"h����kmh���,DE��"Ț-�h�dDMm���h�!DDE��h�D�h��D[i�Ț$YDE�4K6�"",����B-��Y�m""�[DDE���",����Ј��"h�"�[D���"h���m��h�4[DD�b""�DY�h����h��mmDE�""ȑ5��mDE�DD[D���""�D[DD�m"ͦ�E&�-���B"ȄM��E�Y"&�"D"Ŷ��m!-�h��ȚM-"D�BD�f�4�M&��$�K,�"Y"IbD�[I��K$I��D�D�B�d�$��4�e�H��$��%�!���,�D�2D��h��$H�H�,�f�D�D�%��[K,�D�D��H�,��I-��H��$�Y&�$��D�&�f�D�%�%���E�%�$KH�,H�f�D�m"D��D�5�$K$H�H���qlq"Im&�-�H��D�-�H��$Kih��$Ki$I�,��H�,H�-&�f��"Y"D�D�k$H�Ki�4�e�I��$K$H�K,�$��$H�-f��Ki$K$�%��$K$%��Ki���-�H�I�I�$Y��D�"D��	b�$��$Ki$H�,�D�D�4�M"Z�$�I-Ym���i$����idIi-��I,�-$�k$�-$�$����D�M�I���bu͎�ĚD�"D�"��4�D�[HH��h�Y-�I,�,H�M-�H��$K$Ke�$K$H��HKik$�%���D�k$HK$��$�$,�-�$I-��Kik$K$$��ċ4K$�id��9fp��K"%�D�E��Y�Y$Y$ZZ��M"Y5�ie�i%�%�i�M,���Y"M!$����%$�h�ki�Z$���"i�,�-"Ii$KI"[�h���K��m��Xse��X�e�-�}39��m�ɱs�^��g� �n�æ�l���l���l�ɶ�Y��l�d6��c�kf���Y�l���LhA�a�m����l�X�F�Y�̅���!f�[l����8mbЍ�fж�����m�B�B�B���F��i8m�Bs��� �lZ	
�� �"Am6�F�Q�����F��ɤk,r9�4MM&�h�ɱd�5�i�M4і�4�MI�4�Y4���4�i�4MY4�FY4F��h�i�kFH���Mi��f�4�Ѥ�kM4e�I��ɦ�ɤКi���Zi��[M4֚&�kFD�kM	�k&��k&)x�d��I�ki��ɬ�&���M5�D�k&�i5��d�4Mm4��h�&��[MY4Md�MZh��hMY4Mm4�&�Ќ���Mbh�&��M4�FI�����M	��i�k#"i5��k&�D��D�FI�k&���MZi��2&���F��i4&�����M4��I���M5�,�D�MM5��4і�D�5�L�D�5��FD�MD�&��kd�4іMD��M4�[M[M�5�Bh�ɢh�d�4FI��i��M&����h��k&��MD�5�M4#-��$[DD�d[D"ɉE�DMD�m"�"&�h��,����&���",E�h��b"h��4MDLM�4M�h�Bb�&���h�"-�"�&��dDB,[h��""h�DL�h�m4Z,��DDE�DYm�",���"""�%���Mh�m"-�VŐ�H��m-��D�hֈDE�E���H�$M�e�MD�h����-DB�"��8E��"-$[D���B��$H��"�$-$Y�Z$Y#V�dDZ$H�npv�'nm����$-l�E�E�"�ą��h�[5�H�h�ZشYѭlH[D�B"Ж�E�h��d,�[,��$H�kmۙ�D�h�$Z&�-���D�"Ȉ�h����8�D����"[k"B��-m�Z$HY��[�"h�B,���[hE�"h�B$YE��"h�"$YM[h��BE�DE��h�$D[DE�H���M,���D�h�5���,��Ȉ���"Pd������_�&#��Q
C�3�������`Zf`$3l���{�9����?����zy�{~���������7���ۏ��������.���>�z�o=~f�����||�;�y����>������v�ؿs�ݾ�{������_�?��O��|\�O���z��8�����m�����?[�C��c�m�?��^Cfl?�����~�|[�>\����9�}�L���g>=m�&6���=ϛ��������'߃�y�6�g��W���G���v����x�g���ݏ���d�:�}��o���s9��<�ѷ7ϳǏ>���}l�s��[�_.������:Օ�_����n�9�c6����fl��l�Ϧ0͝�f�6���i�g�[m���l
m��a�yvs��p�s^~��ι���;���w>�������෰��ljc6�09	���$�j0_7�����>�7�<��z<|���}}�ϗ�o���\>/!�����w�w�~����^7��h��6ϳpy��o��6�<��ޏ�o_�?.�G��]��������Fo����o��>��ɝ����|	��o�~��>[�~��~>_��o�6f�����5�_n���~?c����yz����G���o��l�w]�pٛ��oݶ��U�������?���c��������?=	v�S�?[|��`�}��=ۭ:�K�ovt{L�fØF������fw7qƏ�f�g����}^38�m+�[���MX�������u��O�ލ�fÛn���$����7��_o}�}Cfl?��;�l~�k�Ϟ������1�����?������|�_�u��6{������y�9�6��/��k�����8���M�7��|�흶l͇˙��~��[o����F��y7��}�O/����z�L��,����F���zo�~��}3ze4�RO���n��'jZ���ݚ�7��s����d�w��g����n�!����#q��j��τB?��[���֗,����#|��8�ov[��}-�o���=7�{����g���}������Ӟ���}3� ��~=~�����l������>���z��s;g=�o��������3�>���w�����OӜ�di�������rE8P���֓