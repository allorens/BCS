BZh91AY&SYt��>�-_�@q���#� ����bG�|>��� �*�@�%  
	���U*��֬ڪ�6�lQ��������B��f�iQi��f5h�R�
�mf�Rյ
���[@�k&���QV��hm�4�CISl����bյF��i��4֊B6,֍�X�6��IU�f�ƀ�تBն��RZ�KJ��ZU4� � ��V ��k� ܺ�V�Y�&p ��TŶ�ef��j��4T��[m��ԳKV�dl[m���i��-�Y���lIi,�$[5�X՚�+� �ڱ�li��  ��   0���Zѭ4R��vƆun�
�Z�%V����e�l�u'U�nں�G\-��Һ�[m�ֻ�k[wg&ӧ]��j�Jh��1-Z|B@  ��� 
_p�0
P�r� ��9�pP �2����zMv�P���� ���

�@�� �^�4�;�:PP����6���̫k+cY�B�����  A��|�);����G�;%�iT�c���=�����{TR�@�9� 
��=��ҁ�4���h
PQ��7��N�4��	�IT�+MZ�V�_|�  {�|J��U����=�����(���;ڔ� ^p�@{^o^= �H����[+��׵�q���:
�q=�{k{�յVm��6e[d��>R  <r��Р
������mN� 9�pR�t2N���� Ӛ���:��G�z��Fv�����X n��"���2�l&l��|� r���W|�{�Ҩ��:��tw��PE�۩� ��;v�Tmf�v���/`�=���M�ˎ��\���A�Zv�%�J���M�����  8�
}� w3�  ׽s� W{k�4T�����	��� �K +���j��;K�= ��F�-�-�m���f԰kk���� ��B�� 25�x (�s@(7p �7 V�9���sn ��;P T¨�d�Va��L�3f�Zf3�@�� o�q� �K ��a@�i0t���@�79ʦ��8  �r� ��� n�͋RV��5j6ʩ�->|R �z� 6�1m�ј� {� �5P 7W#� MӀ��{�� �p 6�>  � $ * �H� �*R�0#  CLL S�4�)RH     �i���	J�����    5< T�%Q�ڌ&�41!�IꒈU       "H��I$�M)�jz�Q��S&��bOMO��ʿ�/�_�g�l$J�I����)�0z
לޫQ��)O�[u��T�>����W�@b ��eDW�< � ����g���?��g����}*�� ��9$�O~�� 
�s�B'!���AE��}�������e��]��6�-vV�`��1�c�)�S�0Lbݕ�6���쫲�enͮ�q�c�+�#�)�S1L`8�q�c�,`c���1b��1�c��-�k�We��]��*�٫��f��]�۲�f��]�vU٫�Wf��]��)��ьC&0Lb��q�c�!�n�2��]��-vj��c�1b���1Lb��q�c�)���	�G�0\`8�q����c�#���U�m٪�V��m�m�[�vjf�en�ݕ2��q����S1L`8�1��#��1`��b��1�c�)�`�)��1Lb��q���)��1Lb��1��X�1���)�1L`8�1���0`8�q�c��B1�)�1Lb�1�vj����]��-vZ���&1L`���`��1�b�ٵ�k�k�We�)��5�-�6�-vmvZ��k��1�c�!�&0Lb��q��0Lb��1�c�)�mٮ͙k��e��2�+vI��11�&0`��1mvZ���ٵٙWf����1�c�	�S&1La�1L`��q���)�S�a��0`8�q���)�c�
c�#�S�0�ݗe�V���٭�m٧�0a�R0L`8�1�c+vmvmvZ쫲e��]��-vV�٭�m�k�L�f��]��-vj��k�We��]��-vL���f��ݕ�5vZ����k��dͻ5vZ�ٛ��e��ݖݚ݃�1�c�)��1LͮʙvV�٭٭�m�[��e��]�f���k�We��]��*�٫�We��f�*��٫�We]��6�5vj��j쫲�f�eWen�]�]�vi����k��e��]�]��5vZ쫱�����)�S&0L`��1�b�1�c�)��1L�ݙ�vV��������#�����#�G0\`��q�c#�)�G�0b��q������:��2�f�f�f��k��0`8�q���)�S�0b��1��c�#�W0b��1�c1q�c��G�0\b8�q�b�q���)��0b��1�0H�1���#��1`���+�G�1��P\b����1Tq��T\`� �
�1Q`��8��"��0q��Tb��8�D�11���ULb*c�b
c����1U1���Lb�c���T��1 1�	���A�"�0E1���QL`�� G�����1Pq��Lf0@c@�".0Aq�#�Ub��G"�1�c�F)�0b8�1�c��8�#�+�W0�enͮ�ݕ�*evmvks�)�S�0b��q�c���q���#�G���W1`��1b8�q��q���#�@�1���)�G0`8�{+vZ�+��e��]��5�+vUvZ�6�+��Z���@���]��������n���B	���#K,~:�U�6�O�{�Hq��7`�GN�1��)��])�;F���Qӡ�vV�Ȏj���Bi���7w�M��ˬ�5Rɦ��+�6��h
�N�X�m�a��s��PY��ů�u�Z;պ��	���Ï�hXO�'��q�,Z�n�*�"�"�����+*��1ɲL�YUm����m�Y��D�L0iDu�����r����U�maz��3}�2x�Ş7�ש�.�����[���(�+�%-R��D��ٴ�57��U#(��71�`�CO�2n��WSi]�G��!�ص��M�����;��-U�S'p5R槍^m��jnٖu�Z�I�Ebu[5�E�1��[���f)��gX��x.�u�(�2�r�5kYZ�NIE�:�7�R�ٻ,G`�%��3f=!K��8�c��d�`��d�.],�-ُv�܃#ڶH�1"����i&�;���
�*J��M-�N�U��Q-��-W�V�L7o\��eT�FC��[�E�Y��1!�!ջ�U��-,�@��Qo(��U)Z�M�`�b&�����Zj,��ZŰZYg��HM�i�0�ݽ­���Z���;c��X�5��%"^��ݳJ�d�ݩ�^�S�uU��(Gm�a�4�,�6��J�2�fijL�Zl�d1�V�qL�I�Y�ctq\&�ʃUM8t+�����餱��ѻ�8�N��^��%�x���n�X�0����x`z���vb��k�BӞ�ri��;QE��2k!��F���6�?Q:ө��$A;O1\��)����1nuA�h�S�e��Y�i
uYd����sf۷Epk���P����{P15�e�I��2e��Z����7VФ�B��,����br���5�;��=Ut�.��{���=�y�ӡ\m�qwc`�Iv6�Յ�6��z���kr1uqma�IfmǸ����$hͧW2�\T��+4R%E�6�{iV����{���ɛ]�·1�M��[�d�
�, �RɌV��ը�f��1Û����u����w��o-Y�2��'"5,��bX�	T�����\9��6�U�FTm��ӁӺl��WRb�Vlǳ$�"x(#�]a�����
����r�E�՘�M̡wKJe��S�Pfaɯ�iX7�;n��o.�fn)�+N�� i;�Q�A�iM��t49���^�m��MU�H��h�Gv��#݆X�bS{R�D�6VU��vFw]8�cx��6�{���
M2�ի�PB&h͙"�*$+q�imA��o�d>�V�y֓ǙȂl�|ݗ��m�6��6�n��KřX�dR򨵭�}.T���w[�#�z��{�wZ���-2�Q���+*���7IH%����IgD��٘���`�̵��vP�v���*�ggq��U���r��sl��z��M��X"B��,�o�R{��L�᡾��p1��dws7����T�Q��&[��9T�p�m���5P',K�����Bn�[Q�{��a�	�D�ӱe;��Oncln�	*cwr)j�UGd#�#��R����7CZꩦ2+��۳Cq�"�w7a�2�f�oD������[�N���W[X�օM�l`IЋb[�3w2b�Eb ���C{��L�����:(�0դƻ����S��[��ܩ���!S�V=�Z�)����zR������5�ݧ{������R���A �����-٫�5��O�Җ�5%�x4�)L�M����l���d��6�3�{vFi�'�we�(�xŽ���bhZ���a�ZG�q<Ip��'�<���'�6�˘6�\+L%b�e�f��#�讴�y�!Z[5+(=:d�*�&(�oE�^]�MC�����Bv��l��2<�#ӕ�U�w���\ʣ��P87&�B�)T�d�.]l�;�Fa�.n��V��-���f�[�\�5Tώ^F�Фܼ�~A�wʋ6f���Z5��x)�T�;��e���.l�NT�觨4��R66,�����7�A[�ɓ.�
�x���k7s*��#�qb���r���ٚm���d�-:�KF�SPV��KIը.�Y�jE*�ϝ�%}t�w7���x�\�궶�/k70E�d���AORUr��y {iHd�:k��D�kV��;�om�ۓ6�b���`������^Z�kl��=ט�~�yToo-�O!{����j�����N��f��N�Ϧ����r=�v��V31�5X�ݬ
i:��,�Xt�:b��Ğ���h3�r��+a�F�A��!�$²��5I�V-���6K�z�Q@6Y��=�k�̦K*��+͆��b��4���0�^��,�S5����7R�4���Sf��jn��ZSD�[X)M̬Tছ�H,��U��[v[b�M�D������T���Yǒ��[q��*�d��\lb����1�Ɓݕ(5���d��n;�n����J�^�N��)""M��q�j���&
�+Q���'��ܢ���Ģ.�a��ZF5��uQa�p,i�U���Z�(l�.Y��j5W	Af0���6Ї%�J�P�s*m��A��y����z��J���Y�, ��f�MĶ]�x�pl�V�=��n�0�ve	1�^�5v�+scU�[Q�`�E�Zt^�K~w�]�8���8��ؙ�K�87�:�ZѴ{$��
�K���_ׇYu��^�]���V˥�:(�X���j�+rV�!����՛Q�#[M�I�t��cB���$2�f]�RF�Ԋ�h'٭ALY���D��w��B�%�<��M�U1��{J���Urfl�Q�!z�n�Â�̶��$ٳo\�4*�\:F
�����1�%.^��:N�ȑ;[IKB1��m�+U$ӘD�&c�I��m#i�!� Tq�ͨI([�)�����b6��4K��
����M�������[jP�$մ�PK�C4B��5�B��vx(ok�ө�eeHH����AHr�1�XB��+i��7P�Ne\�y�@��i9Or�!�,�HȘ�̥I0�V#t�%����J�S���1�hdx#�Fn�-��0��r6j�"�b���R�J�،�V\ˏ��U�#s,�2�Ѭx�2�����*�@6�!N�CtFުT�ǒ�fb;�«-��p�")ζ`���0��o���;��&�&5O�����V�Έf�ɛW��f�O&q�cd���[a�N�ŋ]�4 ǔk4f;�2�)��gPz��Yd�2�����U)0�GU�^Q��1���0����#�H衯��Ξ�NU��%�/�A�Ei�!�hcF;��-����M�F��$2��]i����:wx�ܗ���Ŝ���[��������mm�c:��!��)i
7��{n�n�SVZ:�]F�ndۗ�f�����]aD�����Z�ak[D��d��g��#~�]��r�C��J;�	rn!w�`�Y!u��$7�ɗT5r�C�l��@������2��ҁ>z�1�D@uC����JܶѪ��85<5������X�H5Ԯ���f7h䆈�OL�ɱ��oL�����U�ZKC+���N��D�i��Y8tkw�aޙ�@��GR,���h���/`�Z�_�w��M�H��U�EKu�n�c����/)k�X��[����\ez=��I-u�0�%��S���j����g*�n(!3#!-w���-��=1���"&�
�
�ؕ�r��64i{l�5�[2]Q�m�C)�v�l�t�\����Z��RX��!(�5�����M!.ܠ�\���[.�K]m�e͡R6�u��2�u
�o9��D��骄�km���2��B�z�*��rk�m�L��p����(V�����Bl\X���,�[��v;ɛzbY�d�V��;�`V�<aץ]��1�i;�^i2궃��71fC���Yf�#w��QPQ2il[�Voqu����m{�noU�@��4By�ֆ��U��&��m����LV�0�A�ݵ6�C3�ì�eƲ9�`�j����$"pD�I7Kz���E9�wD�M�v���[��aͽi`�y��7�����\�W�^�IHq��K�qË4�b`�6�7-��n$�/^�Ymcͻsnl#)R(Y�Y��Ӛ҄^��Dk�%�ǘ�l�bN�[uW��L�t�L��H�7p3�7�q�a!caYaD��-��5-�iZ��f��2�Ö.�i-�F��d�FҲ6@�*"�9�]e;���;�ݻٷA�V�,e@�a�P�t���8�l��7���N����6�֑I<��-�e���2��*���n�5e\�X�kgn�H�^�q�iZ�EUenQ76 4�[nf�F�#
Z&b�*�_1���n�o4M�g�D]�\���Ҫ�ؚ6�����A$-�fm 01Hhc����l��媆������H���R���/����Y>gm����m!P���*Be&c����Fãʹ�)!~ ݭLM��L�V�ņ���w���uG�Y���GK{5��!:/,�'�\nV8w��<tI:�{���*ʚ���0mmR�c�O#]L�YaaJ4���
�����9�sfK��jfm��aه73b��Ɂ��g񪡛4�Z��p�%دsf�v��IBa5����k9���N��J�X�D����+�bθԕ��)����W���
v�Yy��we��Jݺ��)[i$un�9�g[`�Fq�	�hd�T�͋d���ʔ��u�i�A��KVWVZ[c5���E�:P�fndFķ
y����a��m��q�ڷz��Q[��n�����*ѭ��J�K�J��PَH�������ѥ�������+!-^ex�'���W��Лl�Om,^u*�<cyN�P��#[xX��CD��bB�ámF��c��/eb˦P�3އ�����R�aCAQݧ`�9���Ik��'a.���Jx�9�Q�8���p�Z�a�Ӎe�Y$ז��1�2�f�g�H��1�{���]Ky�NHsi�Ҧ�J�Ҝ�S	�z��*�.�����F+p캄S�Ǔua�KI���:�E:�H>�+o
֖R��wO0����{
Z)=�ͤ7^gt�T��^��[v�#Xi�IH���7jƵ2&��ni�gi}5�&����gS|5���64��V�`��C��^�w�*]g�)D�Z�5b,�c����L�8E^U�+"o���qؗZ!�a8j�{O�0�Z0`�y5t�Lz����&�T��y3t��ID��0;���6��[��ᚶ!�,�5�&f� ێ4��bdf�z���Ak�S��)��r��;)����m�4��Q:��b�]�*�ɑ�d�#�77):Oq��CŹ�mn���8MZ[[�HtJ������7����a�̀��̡����ݻ��x�Kt<�`;���X�sE��KI���mBa%ܼ9:��̘�cj{���\�32�k%X;���/p-i�`��X�x�� ���o�e�|�Z̼��i��DЦ�7��eM�wi��^՚�qB����nَ���Ж4"�1Ӱ�٣5Q��Œᚁ���,e����R��˽Ua�1m^��J*kkj�a�X�7FճG-�9qM
ز�b�Jj��-��Gf<ʺ��۽.��C�e������4aT,���b����lC��"�Q�����)���2Mɪ]�,i�^3zf�H��W2�m����D�/����`���f�OV�oL��]�$-��I�<�i5�6�%	��YP�fn�^Q����.fV���L���\�x�#-A�ihv]�n�k2���UH+}o�2i�T��p�4�[x�g5e�7wj5�	��In����M(�6�V�mE�:��w����9{���+4;B��bh���3%^Ɏ���Ƣ
!���SZ���D�׹�C�T���4h��,��c!e���H '�ƋŹ��<�u}V����wb���� �4�쵯��E%���#i5 ���┧�u��T���wH�@�[I%�E�U�ةY	lyTV��*YŉA;-Lu�ˠ�:����7W:��k��!p*PgA z5�W�g �r���P��X�F'�r��Toqբ	�iN$R�U���;<�^LJ�ݺ�[V֤�H��5v��j���jbMU�K�LE��}&�Ɲ(
�匾�xn��Y�� �@-��d"���MYK)H�$A��0�ԷU�l68�F� ��J#`�nբ5�o���.���\
 z1���8��H�0ը#��W� � &3Y�\�%M�$�*5�v���dVR�vZ�@�՞U����UJ�^<5m(�-)bX�,�Zط/.�f��Wp:�"U��¸LЈdki�Mb\��z�b�^�1U��E�-x,��p�0l�^�vѵQg*�5S��n+֨���8���Y�ͩ%Lrצ��-&GQ��W�J��z��E�J�Ҭ�)4�
i�穈Ͻ�f◭�� \��z;��qd[��9E�R؍�H�o���y
�l�r�;s���<��t]^m�+--Y�4��F+�qF�.�1d�A�
<F`5o 2��g3�	�R�.�xKڲ�RZ��r��T	k�8��i��h��F,K"c6���" � @A�����YkJ���� ��&�4�n tc	޾����+������=���-jS�{��Et)��� �VR$bM$�`��x,�����lX��@;J�\��J4�{��<�U�b��F��Ph�h�8��p� � v��lf��� ��~���{E�`v�m�)��`o�@�d�(Z����لz���-�"b�N.�i](T��R�J�4A�U��I[Y��|��J��r?4��~���/m���?=��w������?B���|�7��Ķ���I$�I$�I$�fi<��,�ANb�T}Xo�6κS����vO�o��UhZ�w�Ѽ7�D�3�7+.�M��O#-��nNC�WxE����жJ�<��ǨǴ!Ʈ�]��d,��\,�F�C����#b�v�����6���+o:�Z0"�KW�3��B^FRO��ʼ�A� �%�Ӡ��glR��ץr6)�5����o�a4nMԕr�L���T�{,<
�׭U��A�iC��&�2fށ�!�|���&���YӴ���:��m_aFIcu�Q���:d�����{oj�m�vt�R�q�;#[§9�H�O����NcE����5t�]j_j�=26t۲J��OD����C��om3b!��}2⧹oqt��.
���fwqj�AS�3��Z*G������h6��"�-SzE+�.��������ީ(�3u�ԋ:�^'�L/&���S�Mݩz��ǳaQP��N�kZ�M����rs$뙘�#g&���$�q�y�ۭ������+y-mqV��\�}),�}����M�.6����79��.����eN��d��ݗ�g"�[�N���n��y�ZWf�$g\<�".ft:,K�72&���R[ܻ����PY�D�����Ju��b'�"�|sl��	)��v�]��I,�3XLɧ���K�A��on�|���fi�.����|����x�#a^�:�I�N'[ی�디0�P�𛳃6����B���\�.,u�M&���
j�%�vb�\�9���*uޒt6*�7�}Np���'��Ý��V�M��\�Ep/9�;:aӦ��-n��m�9ݮ�S�9&Bq��&X�q�r�9N���%,���E��t��mnG#d���K}]��n�L&	*��̳)��,a�t��\(�M��ۖ�R*
��d����{i�c4�5��G�������	�h1��2���$Wӗc�txSqK�q��e�Q�a���"@Ν���H$w.)3���0!�B�ftt�q����OT<'�F�"�U���:/0��K�f
�v.U��݇G��/ޓn�VCGL�tk�2���IB��WZ.�Ў��;��<��vu��v�*`��+f�A�(�tj��r���'�#,��Ujۦ�x�ak^X�p`�/��p%��;�u���5b\��.a�d�o8.yB����^J������<os]�͖�3���}�y\��y���՘B�u�suT=���Z�ތ��6Sh�we]�^���p�i\��gw���8�.uP-�+3U��9�/�ȱU�ՕJ�6�v�[�[�Sj��v�+�Imgʱ������~��~@���[s�޸��7 �vpm�E��JN��v�m�����.�V�ʨ��ۮ��̜�0���m��	�Xƽ��թg�Lt��̨�k�]M%�y�W]�SC7���{Z�0�|��ݗ#�2�n���9�C�k��C�3����G}�:���38rm�5��M��3wM��w���Y��e*7{�FK����n�J7�2.%l ��[e�}�v�B7�}�N�7is(ůn���1���7�v�G���w�y+4�]7�̒�7Q���.T��MY}�㋒h�s&v�ږޔ{��bѯ�3�$�43�U�W���$&�����`�ݓPn��WP˓�b��� ���~U���a]-馠O	�IL�a�kYc��IN\y�)��;�A��m�$o����x�5PR/��f������>g�$u���-U��隓�>��xپ9�m����X����gHn�K�p5�&2Mf؊5y��d�N�f-%��������\��&E��=��ʅ5v���2���V����"[��z��M�Ӵ�P>�N����ox�;/1a�Sb؈+kѩ��x^��&Ƅ���7j�7��Gut�{ǯ�U��.�;^�哙 M"���r���T�^MK�Vlo�R�%�f�ljZ˾nR�X��,�����^�v���Ed���:��=�n*�W�@c+BN�݌ev�mͮg���p�'T�;c����4�{��`[�Gc~��ˮ���3ٍf3H��mw�j_[��ϳ������f��	6ٞO�������7_�]̛PV]��GB&���#�!��(��i��NK)wL���+�Kv��u�9h������E�s�f�|L�Ȫ�o�ۧ�����$p��5u3�,p�u	�l-.�&���ө��u�P�y�}F���p]L*���C!�a���
M�Y+�m���� ��9v�����͋|%���Ȕ�lN�M���|f�΃+��/���Q���΄�z.�VnK��6u*J����8�p{��{~�2+�Y��v�����RՇ�:pjUvU�N�v��<K���\+���)�HK/y��Yn�+��7y��5����gܼ�{Kl10�
����f@�4?�LPfCK]���%�z^�ǧk��9;M%q#+"7YBS�лn�'�2�g8�7wݩ�ͻW���5��]�7�V;7�3x�Wg�T{b�E��� 1�1q=5e5;�����n��!N�^����C(�w���sR�绰�3>d�bgz��������Ab��5Ǎ'*Ps�1A�nmmjKa�uI-�;�=C�]�̝�=V�q_`Oh�2�,��y�+#5H�$[���{0�-\�.�B�*b���8k��d�U�q���wnCN+�����9�_'J�=���ol��P[�;;�����-�΢1�v���	��J˼�B�D�x�h˖nbjYmY���!�z�J�'&0Bd�o{�����G����ڀ<c-�k�����'Y|�ë���(�$����[+R��`>��\uf�C��	pYkdӘh���x0N�g6�(F�v=+��e�؜t�Tc����T���&A�Huu�v�"ИL&��7��}(���[n�ek(���wc��y�!�4
��L+�0�o�LF��@e����駮#ӝ��\��S=ťZ/U�q���
-�$����e��/q���|1��c�иv%�M$�=j�f\�M2}hUv���ϔ�I��ξ�IBK�\���A�{�j��A��V�r��k����z�u��5�S�2��xt�j�K7�ټS�&�i�互�,��t�ml¶�Xzi����G�]����gVW����9���&�)sDoU���tX��/ap�����Wb�$0^!�w�f���Ձ(�������v8�+�}5;�-7���b��T�FD�*;Cs��՘$o-���0iO����L�,�oF�,��\lP��'b��vۮO�b�N���\��jiYM�iD9yJYצ�*���p�]kv��s��Z���N^@��t4�Lw;}�Էh��f��C�fF�)��M�w�7�aN��N�)Q8n�g(S:�+��yC�f�aΘC�
��,Ím���� Oq����j>j�2A���2m[�)���fgA.u�0��uQ�Q���w���Ы��I��b���76˥��(�R`�	'���nv�p������;J!��	\�aɉ[<����K�b���]X�1-7�_.�}Kuƞ��O\+�eC��0��Jń�����מ�ڣ,�����ٹ�-���..�!c��Dx�,���,jYfg��9rv�t�q��o5��\��H�F���S���l�)�]{����&���U����$�[{[C��cG5{t)Y�k��5�ؖ�L�ܨ�zڌ`�+lκ�#6�vR8���,2 M�V41���ci����{ZV�z�i�v���T��;G5���@��ϛ?��^+f��[�y�:��>Q����c���N���s[i����Q��j]���ݴ���K�e��i*zȾAN���t�M�\�]g�Ɛn�oh{����ʲ��]j���4���Nm_��g^c:c�i����	�ե���5���Ȃ�=ҵdM�c.�����Ofg���׵�V�(k��Z�M���z��ok8�jh��n�h���r��-&н�r�)6յ��f��8c�4���
Yc��a�����A鯑Ż�!�F�����\zrX9/33���ՠ"|�`q%f��6n�0�r�1O�u�>�W6��0K�Nۖ�˦�;�E��/t-%	�f\'M\��8� ���[�A�o:��8l.�L�rh��e�A���zȐ��6���,䔁��V�T{4��f^���m��k�Ǜ�
2�%<���nY�b�&Xc�d������u�tl�SF��Z��fLޡU�#�ơ�Y<�wʱ���Q�r�b���l�[B�7��ԷbӨ��n+6;2��Ȃ�iJ�{�:^�O���Rk��1�iM�dwR}G=Z+�~��LKb=q���s���]��)]����x�RX(d|�^�bo���d�%N*	j�j���٭��C���Z�4���9�o��Eҥ�v����C,N`55�#T֞�d�����\Φ�mJ]�����Ԣk�	m��*���%z���l8��wV�!ጢә��C*_I��sCc�0�ëe!�Zo�Zg�;����!M���9g��G��;�愠��Kv�F�Z��4�=pv�;p*G��	O^�:�ř�-x��z)<�8�U���m����8��ӧD7�ʧBc�{^�m���/H��}|UL�͢��0T�w2�dA_DU�v���:��xor��i���Q+�z�''u�e�R�{jQ:�������mAӀ�̂��r�Đ/"n;�ѿ];�]�7cz�>kn����C�[G1d���v�)a�%�k��`�b�鈩T�%3��xq��]�$x/LiɇR%��S�K���M+�����^��Z�ІVS���'(Y�V#o!nN��� �_+ڥH����Ϻ�����W��}�d�g<�v��+fK)�Ɵi�&��H9}��׈f."�XoXxB�h�w<�ǹy�Gv�OH��Z�&�/�6���	������Dc�3~�-�XuO�MO=���W�1�uuwJʽ����Q�Ʌ��6�z�4oz
����)��WNv��
��</�}�A��&k�ي��.�]�#i����p�x(>��$V~CoVv�Z�c+��de�`uXT˧�b����n�%.죋I�uE��ٲ�pD��7g
�����#QE���a�L�v�w�9%��H\��*��n��V�͂H���"��J8e1�/�Vy��qαu�2�S�4�ݓj������wVwa�esa�ө�,鉛��vJut���M\�[ڍ�shd�s)5W�8�,��)�a�&mC������oޔz�X1I[����Nsv���r-k4�(-�Wt�a|��޹��W�䫏^����Â*:b�S��f�Ƕ�����6��r�!��y��tm��;/vJy:��w)������YW�|��g��44Ļ%痬�[��}�Yz���꼾N��������Iרu8��82����i���9t�'k�K��cƵ��[���!3'�u��5D\�{�j��˗����U��»;$6�.j��+:��x^%��h�]<���bp��/�W9�Zùs���,L�hM��&I�(v��z�v�S���0c��	��q���un\(m�4���r{I�e�0���9|�N�2wa^7�W%�V8���6~ۉK�H<�p_'zmV��5��'U���;:*W9Σ>�0E��Ǧ���p�GZ;^.��7,������Ĵ��ݜ�*2�6��8b�q\����̂Y|L���`(.]���x�_K����Svt��[�Ǿ���[�v=����/��3��N�J:�F��._�Cz:����4vQsk,���=�qKW�;�4婳uG}(�XyC4���̰I�$KK��r��i<�T�4�(vJ�n]����Uc7��U�Q���2�T��S�I6rRI)�$�I$�I$�I$�I$�I$�I$�I$�I$�I$��}����\��Ŗ8���6����rI$�I}�v
�u[�]jby��]h���K� ��o`� j��̦ u�u�SDS5��<��;�����{�C��9��X�l�9�5�y��x��]\�x�B��ޱK�"���\�<���	�C��Sȧp��jru�HI�Gq��\��` �S���1_f{�}���/~`�u�#�!���IE|�yEz��%���̐���'��]y��9�����`�;������(d����G!�'|����L��z�]�y�'�`�P�E�C9���?��������~�AC�r����'����J���AG�?����}���?t����ο�?#�k��o3u��ov��7�J4�y��񋿾���sI���Q�;��W�3MV�;����y�.bŻ
��u[�l�݆;0S�6Cx��m��4�"˸0-�2	��gw[���.�j�����[r�����FDj��sI2w{2���W3rѱ�W��5��J��V��~܎���r��[}��MVk�&�ۮ�<&����1l{3�$�}J��7�P�*H{-�DL�ݍ�2WZ�� �>�c[�f����Xx�Z/Od5�<fb������a���qew��_S	�B��4��E�<^Z�1ܜ݂_l�(�r�J�Ǖ���OM�g6Xq]�����l���6���u�F��k����4�|e2�Z��o�=+s|n�,J	��ޫ���d~�p�K�������my������8R�aiv�53z�&�#\0*@����'H )!�3Dꖕ1�c<�#_s-	"��R�*;׷��43�j@l9n,�����l\����r�rG3;e�.�ANS�Wb��̋N�Φ�6+��d��Y9�L'-,�������L.����������u.SR��OyQB��Ǜ!���:|���Q�L�mF`�`���'���~�|u��F�aǳo��g'2�V�r{]V�������5�毟��n��Z��׍cZֵ�k�Z�Zֵ�k�Z�Zֵ�{kZ�kZצ��vֵƵ�Xֵ�Zֵ�kZֵ��ֵ�{kZ�Zֵ�|hֵ�kZ׍cZֵ�{kZ�kZצ��vֵ��ֵ�{hֵ�kZ׍cZֵ�kZѭkZѭkƱ�kZֽ��tֵ�kZ�ֵָ�k�ZֻkZֻkZֽ5�kZֵ�xѭkZֵ�hֵ�kZ׍cZֵ۷ǧ����kZֽ��tֵ�kZִkZֵ�kZ5�kZֵ�ֵ�kZ֍kZֵ�x׎(s�����<cJ�s{Zr�ȭ|a�	qDs�P�u/�5��KCj����Bc#fA{gv���k�j�Վ��k���Ɠ��J�rE�g����f��U�Ëpu��Q�(.�$�r���d����8x�;S}�J�*7�����MK�2��:���љz�L�كe���x���M���pF���1�.`J��1��V�u�I}���5��t7m�V���x��o2*.�ĵ�4 �;Q�=�]� 6n���Ԝ8�;iZ��U*� �:��G��'4���%&���mB\�U�� ⇺u,ŧ\�e����BǝZ�5y`F����6Ɯ�����(�;k7s�g"��*Q¦��ݜ�l˭}�[�ћ2��	�ʅ�}V���C�ȸʍ+*��KbW�f5����>��aە�6K�,k�y�%�)R��e���U`�Y��GT����Q`�m�ǅ��\op���2N�5�owC�E}%d���+�s*7���O,j����teVV�`ܶNq��S�u���݋�Q_�����L�7�S�h]T�sg��G_��(Z:I��m��>�h{]RR���\��ǯ4L� K�rV�oV��r�Wm6�e(TŪ�F��8��T'���6�������kM�p�y�����s0�-��]s��==�{x׍zkZ�MkZֽ��kZֵ�xֵƵ�kZ�ֱ�kZֵ�F��kZ�ֵ�Zֵ�{kZ�kZֵ�Ƶ�kZ�ֵ�Zֵ�Zֵ�k]5�kZ��kZֵ�kF��kZ�ƵƵ�k���k�ZֺkZֵ�kZ�kZ�ֵƵ�kZ�ֵƵ�kZ�ֱ�kZֵ�F��kZ�ƵƵ�k^�ֺkֵ�k�Z�MkZ�mkZצ��5�zzv��ZѭkZֵ�kZ�Zֵ�|kZֻkZֽ5�k]��k^�ֵ�zkZ�mkZ�mk}��W�m��f��Q��F�x����k!�
�9�����"�xї�R�R��E�ETw�7'+��JTх�����Q]�PBaQ�t�Ѽ�w͘��WA������#�����$&�M��gC)b�(�{;���F�R\:�_fD
�񜱤^�.��ӓ_Z#o�͸j�OX��EӒ�+���R9��ܧBQRG7��0Ҹ����THݙ�����d��>�CG`��8E[%��L���,&[Ѫ���=���_f)���e<̚x����L_t�@ڜ���4ec�����>�i�������12j[����.T&�����nWS�Ç8��b�]Y#��O��WA,3ݵp��Z)n,�}��9�%�p��1O�0��h�s{�
�����|��y/q�-�HU�u��X�)��',0�z9�]�I��w�Ҍ���C�|��Z�=��K�s��D���;�"�Fں�����u��B�����V+Z�=4Vu>����ϛ!�ђ�[��AT�9.�S������Τ�}���&�7/5�zݮtzd��#��:��n;K���-���3J��S��6���C���M1�|�ޥ��QM[�����+U|K膐TQ<}�Uy5�m�&�)Vi7k�b����f�t�ӽՑb��d]ɋ���Um����JVa�G꒞-��0֖��e�/���=Y}���yGJo�]e����H4Y�#$"�L4Aj�T��f���n�E.ؠN=Wqa��-jd�r�.��QT!My4g$��#X�L������^S��w��v3���m+�V����St����ܛ[���:����-9������=�r�s���k��C]ԙ��j��e��ݔ�ǡ]�3�wY�7Ty�e7b@u�lQɩ��*�
"P���M����/���,4k��`<����'d�iȨҘ�]���}Gh�u\��=�/L���]����ɽ�(h�tgV����'��.�lw6��ߘ���6�Th��q�â!��u������鎌�mt�����(m���J��۩"\M�4S�4+���Ѱ��^Cw"Ӥ����ht1�]IW	�-��by3�}Lw+�o������F����م��7�Ě�X�V&�?G�<���am�_��wa��m��7�c1Q��.Ɩ>�}��f�9b��`��Z�i�+(�v<��l���MߔzH�,��Lmmh�����9,�����K��ۧy���|�f^��'I:�,�ˬw���8e;�Z�͛I�A�J��؛n�YN�QoFqY�W���vn:��
��L{���f5��T���SG8�r!�hز�kC7)]�'���N`����'��fH��E����Is{F;�Ƶ��]Y����0����t/�&��&�Wp�MȾWB�:ƃ�88K��M�����ntaN9��r������}���3*\�L�A�H����^V�f�o\�:�(�-ݩ[��|V�Zp���C�SC��&-y.e��m�F8�q�b��7������j�7�#�E��Eq�d�-�to^�ռ)��+'g#ln�����5N��Q(�k��ܲ[96ę�������nB�9м�s�]xUHu��ӭyTj�^�r��
�ה
�ϢǡyjN��������N,����
�Iݐ�q��,�s��Gp�β$��9K�Z�է�,�ۗ���q��nW.G:��蔳��u�z���w�����7��/t8��[Y7GCIu�@�ē�Zܝz��7Rs�{������y�����l�kKQ���˘��T4(i7�m4"w��[��t7�������A$�X.�y�um����p�����4:4*Th�ͧЈ�/ztV "un���Z�P�6�O\u�J��ǪCo���rS��k�ruw%s1$p>�郑�st����	*���	�4��F�����8�й$�X�;�[0��J���1es��4W+�p��l��5�E���O�������Q��]c�;�ښ����r����iJ�n��>�88����7��Dt����������9�!�1m�a�1���*�XYY�mE7�Q�.\��������/cQ;n�%��|!�z��h62!���],]u��\<�����l���Nž}��w�Q�g[�{֯\�&�9�oy�n����V��V���5����T��z/q2m�3A���<���,f��y\��.�3F]��Ů��N&�V ��d˾��1�$�s��ڲu�*R\����R��y���7��}`^�K#�T��i��@�B}JSc�y�dOD�<�_R0�b5nR3S�������	Ȱ97خv�9���Q�]�\�0q�˹@�+n�ܘ&v噞�y3rT��T��S6f;�M�=�5J8C���D��N���f;\�Q�.�6L�å3�հZ�}S���m��9�eLe�XX0ٰC[%H�Ϸ;sJ}�!�<��7k�4hEb,I��\�F�U*�9ّ�*S˶�;
&�w�3�M��M��ƥ�����/)PG
���lpA�Av���Q��l��T���K�ܱR��c�Mn.��yhS9��6�[z�Ya���68�b���M�.�͔r;tlix��wg�{�dE�0i�#��[ͣ�y��m��d+G��sܸ�}X�����ρ��e��� �z�=��r:��Z�ˮ��r��G6tv��uv�N�a���n�,+��2��c��sV�O&��t���q�nʌQ�����JҹjN����1���Onu�Y�}{1t$@��o*���gS0������9v��7�U�0h�%A�D�$�{�3E!����3�LV�[b�=	m7QR��4SN�Ժ����'T(��->��w5$3:��dy,|�B��!�Gp�7c��|�-�v�KX�/��bq����X�WF�R+-["��.�?��*�M40CB��WL��$� ͖N�w��������y�eRUd'���1�^�dޟUU���P��7��*�-�=���ѷ���l�ݕQ�3����xFb����Y�U�3Y:\�ن)�hW�r롺�w;9uq�,�sܻoJ$T(�O9jD�ηC{m�N�b��9�nL�Gc���WIY>�j�ʔ�C�Nm�k��;v�3%�*�Ѧ��[ewj�� h��j�^nl�	T�(��l�7S�ޚ�d[��^�
���%���a�yG��J� �X(3����7\j}w7yZ������ʀ���(�
��fհt�Y�٦��|Y����"!��Uo�,�*�=M�x>T*���:K
��72d����.����R�t�3S(�Vc�{�ۣ��^��4�IWݐ�����Kη�w}[/�l=$�����i�Xoo�d4�ݪShn!�r��'��ųSYZj�T�{8miP��\[{���):1��2�i�^Z�+7oL%���&�*�0���1T�`ئ��r�;��! e��k	�U���"��M��D}��a�M�a��U8v]��G-�ዴ�M*����[WiŀxֽwD��y�MX"7{�	s���<��G�/L��N��%L}V�|V'����-\��W�I�3��{R}�9��h��*L�h��]qj����Μs$���n�.V�8��x���`���;�!S�ڬ��e��݇�%;�SB���gh���;V�Г�uB�N��Υ*k��CR�n�)�UW|���,���C�'.�X��Ў;��<A �� F�f��:�^n��yY�y�ʢ�B٠gaB�Ei�:�\�ei5�0P��͎N��K2m������W][W���]�n��	n�33�c~C��-���!��x���m����Ѧ����]컾)��p�k�@��Yf������1plx�g��9��tiS�C���qᇂ�R�x
�4��$�)ͱXM�����E7�wK@����TI�A]�f �i�!���gwퟧM�D�s/��"E�V���;�s2�_C8��0Xx#��vHP��<���s2C+ଔ�k�rM#�@`���$ՇZ}C#pi��5}r���FD��ڬǝg�M��{� ���nDۑ�&C� �}��c�-X�(2�U�ж+��8UgPXrKĤ���e߃�5͒�TH�C*m@Ľ.����k
�շ�Ɠrﳉ��=�ϝ+j�֎ޫ ;}.'/u�Ι��ֺ9�(��f���ó]��B�*Vrʤ�m���㷆�K���ut�RR���l���'Lbֆ��1L����fB���z�b�.Mx���p�%u����l���$ک2Gyo)��C"�캫MV���sQ&e�\������J�����[|)��ɼ}��O��r1�<�h�m����љ�Z��!u�S���eC�;Y&s�G����ܰ<��\���|��uD�:�]G�c��9�0�8�VHӚ_U�P#��F겶�, 9�ʠ�G*�'2r��'�S�չN�Q��<�M�0Ҹ�l!�6sj��M}���U��-��E��E����}�c2��μ����iz�A\i�$/�|re�5�zw\P�;��_U�t�:��z��|��#��W7�ij��{z�gb����j)ñ��7l��9�kM�mu!5�v��%Gf����q��ʳ��
�Mg��we�0�P{�mЂ�wQ��5�tF3�n��Ǻ0��]S��,�\���hk��*:�uDg[�vJ���ʈ�bYCj]4����A���KpM��u��}4�ʚ�`�:�v[s`9G�H4�^�e۾Ģ���e�rg�7Իa0�L�n��������b4�S��35MX��%���٘��n��g���8UL�|��@�m�����]�}����Mn%,ZeJXUf5�݌Gk,�v*���6A�	��Q�����1NsH)-���עX���B�?�罒ښ���"]�s�C�'3�{�+����t��-'l�Э�r�.v�KK��`��K�����a�r��ݺ�&�ְ��Z�/[�v;t���8v�[��ޭ}��C���,5{�#-c"G�z�Xh�n�k�5�._��B��`���M�L���O�V2���CS;_���  
�{!�?���?���������Bh����Z�0K1Ą�D�P�l��N!#3�$!�h*2	i�d�&���D�
 RqH�R��i8����n���Kl�=��TM�2F!��)$,��AHe&YD��FҪ��Ā�p����O
Ӓ&�E�#BP-[�D����--�U��l�қ%B�(d`�"(8hA0�HL��N@����b��q�lG�I����pF)
$���JOE	�⊝R��h��my�	$4�.)Q5-0���b-����\�?�J�/zv�e#5cy�M��+0$�`{�L��|DZ���U�YVB�]�es1�3Y�jw|���8J�_t��*N��3��4���<r���2]��8uv�o%�.�b�l�R*=!j\�����,<r54ò$3�d����`(�����ι��v����
\��:�W�Y�p|��v\ښ��gVeʁ�2@��jfnXc\�W9Xl���mZY�����5#�I�0H���L�`���2��jai�7�����H5q`7�[�y����iI�3d6;�;\UM�RƖ)�Ĉd���:��Ҫp�̜$Zvcv.����m�]��y�*kx�"�n%BI�L�+���뉎�ƴ��2M�oK�Qu)��2���㴄Ng	s�a�S� �����T��D��/�F�ˍ��;���T�yE�����oN�x8�ݚ�Gh�U��;i-�^�˪�7@��Qe�(\�F�V�qѮ�t�ΛpqvS%)��H�N�h�u�r���W�C:qurT��`�,�`��Ba<��	�rod�27z�V�u�ѥf��N-䜧���.�Թ��M�E�?2j�����Z�ͳ�m�Xų�t�a^.�^c��G�	�e����Q��*I#NI�W (h�fh���26���"P�lqBP*#o�1P2�A���d8�BH�P`�\!��(�p�H(m0�l��d�'�n6�)��
I(�@��d�$�P%8�)1���p�T��ؑ��K�"���# ��U3@�P@�����Q�	��a��L�"k�1l@ى�D�CA(�0�T��Ə��eB�i6�O"c00D�)��D(� ���	�$�É�$k�C�?b/�	P�Hi�^jQpD��F�$�	n �H�LH�AS
�Q��`I0�F$byƉ$�m��9`Ȕ("�J4�p�#l
��
%H�?(�e�Pp6"k�"�)��m�܁5'�%c&ڂ&�$�b���6�a�聁%�rG�����!#�����H��dH$A$�p� ,RUJ�
"d�dF�n �A�Pq4�N�A�Ą#<�! �A�������2Xn(�>fH
d�S��P�Sf�Pę%�cL�$P���L:,� @e�I��o���]��]ݾ����[]��;]��;��o>��y]�1�==���xѭkZֵ�hֵ�v�۷mx󄄏3$$Y/����\�o7�^~+y�9�W�矪�yp����1��Տ�ݽ>><k�ZƵ�kZ׍ֵ�ݻv�rD��0��E��u�ۈ��ߵ��=ۃ����wޯ,���f���;��W��ߝ���cDϕ۽�����S����ޖy���VG�����r_��j/�����.y�H!<+�����Q�-��_&�)��L79�J�3I��nH^�ҿ?=��ӧ.�J���ǽ���{���wt��^����s]���[��ݱ{�틎��5λ������ߝy7�ocҺ;�����o�뱗wSs��价>u��~���q>�Ϛ��u�i���~�D�ZS���[�u�{�W��9w�{S~{�qwr�u];�����w�M��q��w-��Me'�t��o�a�;���U˻��;��������+/�v���w���z� �{ں<���cݭwQ=��6��w.�і�quv����72�	J? J�3'��x�Bx��D6�E G� �(�����e	m��dbD8גQ��I�	8�l�#���%4H($TRw��~��8)y/i���if�̕
z��rIc�iu-�}՘f��`ɵ�e��݋��R��s\��k�cZ��)#��R�Q�q��$�0���9$��(S"D*\���`�$��B�!"M�Z���1�Q*&�8B�n��BQ�3Ȱʅ(�R
&�r@b�G&g���� g>ޭ�2
���-����͊n���]A�a��Q1b���r2�5B�����+����:�g�Ρ��>т:��>vX~�(�ٻݧ3�O@�!ޠmY���m>��G��ڙQ���a����TX�o�+y���4v���>� �{�zMǚ�n�m>�4O$�˾Ge����M�ӝ6|+�����q��܈p3��[�;`�9��|��F����%�ϣ��tՌ������Ϭ׳%������0�����=�[ w\;w_Or1�)�|���3������f����SK�nA�v�И$���QNzZY%��šP��y;>�?x�y�=�e�����غ�9��R��H��*?;�eVD�ߌ��+���^=�~Q���E��C�٪Mm�I�i�~~"7����s�6G�}���
{��jm%�=W9�b�#�7�9|�m�ȯog�q�*��"4/y��W}�B�.�z=��^SC��㼨�3Ǐ��뢿`��j�t�Jk�`�;���UTB2�`�T86���˜DU���"N��J�؟ݦ��c�:����+mŜv�5Ǻ��H˔�`�!�Eٗ&,�3�"�IEKMl�&�����07l�{�z���>?�ĺ<�q���l5mֺ�>U�1t?eya����B��.ھ�{�Bt���nX�|#��7�=Xi!�=Z3�0�~���~�;+�x<�~z<��U��?4{s�xw/>�_`�-m[?�)�t��;x�t1н�����}�8���vOU������{�&����g�C,���k�Gl ,�����+.����VU���
]B�	��sxz����2\#�2��ᖁ9��܅�ae��D�g�_����Mf��oT��Q�rs�6f�t��i�w#c��d����Վ�`��/�;�E�]DyuZ�.��.>Mlܹ���΅�1$�P}���4�m�N�w�ff{�Fz�9����ם��{V���oQ�<o��x�v�M6֊�9�:��ǽ~��8���}s�R�^��7��og�U�W7��o}�������U�+��#���_0k�-��Z�X7a�A1�@T�V(�!�Q��Em5�Ԗ����Y]��xi��:��<��Ÿ @���#0�I�xȶ�3���X��9����J�$��j�[ևe96i�k/'VQ=����I�����.Vzu܀ϟ���YD��w\L�
z4v*}<!,���$�����y��('��y���v��2{��Nk0�>r:<�Y"62}X�3�^C鞯���T�b�g�"�ݶ����V+��*鼡�7=����������ř�u{wV�\d��;��o���S6g�����7����ˊ��� FPqoj%dߣ���{�玦,��>[V����땯�y}������מB���T7��r�))���ϙ�_p�J���;~U~�(b�[�^�S����;>O�:����*g�K��*1��j���c��[���z!��L��A�y�Q��gX֤��'��gR��~�C]"<i�cA{>������h_���!�VN����=��W/_��������l���,u��PMݧ��z��Z��W�t���L����~�~�5W��)P!&�;R����=Q�����7h�5�.cGdz��TrZ�1g]b�wt��\殓GĜ9'N�MbI�l�E..�]��-��V�P��#�a2�ࠫ�ܯۛ)���{�;�B�}_֖8�|����8��.I�n�x~�``A���F1&e��Lo���PHz0��Z�8��[�_�{��_��=�+���A޳^���"S��&䜇X�V�Wz��>.�}�-�$7=��5�Om{ąظ����!zt�Nf�I���&�������%�4��q;M�g��T<I����Fu�v�o���׼3�z�g�y�d��{)1v�I����Y_��Ϣ��.|�|��M�c�.7���A���NȽ2���iț�j�zai��.j�O�z�d�{�j��������=��6�Gs�38�.�&�=>��nx����ssO��s��B+(|FO��]x�k�]����ެ}�k߃u^�;��=�j�ꈦl���6&m˶�!���f<�<&�y��v^��]�3�4��hǑ�gw`�ۺW^p����~��Vo�����#����r�<�S�M���'i�W���x�@��g��K��Rp�2b1�Qz��֯�z�$������'9��1gkց6�.Y�rw���{�3O+��KF�2��ξhĚ������d���t��Q���;��A�EY�o�tͫ�i�",�T��ePKE��0x���,W������?����S^Y�Z���[ZFE�z)��������5w�s�z��;�+u�_An��C4�����o=l{�&�)�y�����Tʬ����mf�L	����Q�Gp�{6U�o!�~7�_��j����A%�5�����NY�ͳ�m�>���b@��7^��h�'j���ˏTK����ȋ8j��Z񬛭{=g����tu����z�����U�����D/��K
�Ɇ���d���-�*l������)��z������8��|J�~�f����%�~��
o?�{~�����\9荖Γ���3�� �3�t��l�V�m�d k��.���F�������M\�+͐�����{�{���<��n��|,��<�kG�m�,���T	��1&=/���¢/�o�6}�}�rf_r�)@�
^�()���Z��R���v�����ޖ���B*�b��7�*�Vּ��5�|��-���\������׳�_%����Y�Ol�y����Wm���$��x��L��I���>��{&�����G�Uo���6���V�ײ:�M^-�ؽ��_A�{2#� ���=���~�Ll���߫��e���4��*t��,=��Y�&�}a���Z}Bf̼7��n��>~����h�tykij$����q#��Cg��#�@��hg��9#�{/�Y�����6���ޝ���K��ں��'����'ACчukW�˙�����3��R��mW?1��.���V��j��^�#p�<'�uQ��M����X��/���9xu�z=�ߪ�Ø���`��P>}B��p�K|y�g�Q��Lz��nmI��K�]�i�<�(c
26%�M�̧��~�|`��`��T���������eœ��;�4d�͖��Mw^a�7����/|g(Ϛ?TA�A:��v��7]���M;�4��]sF���<�]�U��A�O}�����	lg^��'{�qc�9ٹ��j�
'C�^蛴�m�c8M@���D�Ȁ~N�m.SWaQw}QN`ރL7j^	�1c�J[h�TH�[;"��݆��%��Y���I�%ة��_��B�*��ܐn݋�5�wmmzï����LS=�͒����*W��X[^=�}z㉼Y,�ܔ�S��V_����Ǽ��^I�n�m1�j�źi���3�3��bn������Gi��$�s�L���I�}��s`��	&��%�@��=�ќ|�;�5�-{�`n�&۽<m��{^�{'M��@�����&�/�"���cϗ�O�ޫ�?o��������ʏg�d�3����~ʲ+�P����x��n��͝�e��{%L{�}:D�H�|{ܯ~w���C���^����2�F������9ƥ�j���:#=�]$�����oM�ߑ��R����+�n.ī_t�[y~��Qp�ˣ;��̓i8���/��>�[V�ګ�^{�^��5UW�����2,�/���"�UUN��RSR5�j��C㧍f����2�ӫn���>�9�K�C��I�x}�&�]g1��ρͫU��X�?�ݫ;�w�<�0�s��ú,����G_.�Y'6�tf�s��B:�n�Ȩ��v���C��+��}���V�]\�,u_I�*}�_����mI�}F�^�W�Ng�~�ƺUjy6J�$��*1z�:h��-��h��<�����V<oO=Y7~��y�&x���ӽq휇�S��8䛺,=�������gޢ�ŉ{�no�t�,a��YѦ��w�^�` q"<+(챿l�F��x�w~=0zm��2�9�L�[���:��zǽ����W1�đ�a��b��<��a0�q>���y��U�W�����:�^>_I`m�B�z[������s]��q�eX��v�I�CW���n��O�x��ܸzu��=�z,z^�"?�x%w��8>��WE<��m��6��sq�c/�g19�����k�.�2꽫�ƽ_cUd���{�;<6�N�����_�c_L	�_]`� �>��`WF���r�.}8M���	�Z�j����X��9n�#.7N�}���� �>��C��Օu�j[-VE�ڰ޵� �8����:�Fc.�X�k��G���f�.�]
9���됽���+7��;�}Y�+��,��������ڙ|Õ�A�];;2f���s�!b��ľ�xk3IB�d��Y�����U@��n'��oQ=�0��g3��!��?�����v'���B�#�}!~�=��;����ǞP���=�-��ψb`_mq��x<�x6wN�H�������J���T��^DV�6��D��&$޾�o���v����tǫ{�[¾����u���"o��u��Ec�{A��C��G���L4+W���Yt��k]���Od�>����$�����G���r9ŋ�<4�� 4�+����c�ryOv��`/��c{���[C?�I�\aW��#N{5���W5�HA��i�I������}O�}�����,N�g=�ׇ�����Jv�{7܆�HP(Կ.���_N���x2I�n���f��H{g���vtKh�,�s4L�X��|Z�I���_�yt�R��n���c����ճ�	9Rњc�5z�t�W��ގW�@�!���M{�:�k:��:��_N�s��p�k���a�.�i�c\���a>�xW���z���<��L�j��j�K�7z��rf�;�X�u��Wy����� �f�ٮ�G�C�R���r�M�W�k��N�ɞ���6�mTy�.�*z��LG�*����U��gӽR
_{��{�o�9뜲��H�N����f�,b}Vs�4��}��ml�S��T�rY����7%�ɣ=ǚ��d�������g�����?7";t�^���^��츯��Dx�|׽&/�4��M2_}��� ������������;G�]DQ��;�c�0���T�s�<)��\��U�S7�o��ݵɗ�yS�jy#�]��ޖ=^Yu(�q>�1{s=�,Q�����ʺ���ױ6W��)T3'����S�NJ��e#�=�y�Uޫ��<�7��#^�{��]��RT�J���o�^�j�>�s�T7q�}ъ	�6�=j���e�eϷ_pK�g@�gy0=9�g����E>�����ֳ�����k���~��h�]eN�k#&uܫG���=�R�ٱخ�����MOM��=-ҷ'0V��s ޳���*1�$��>�,���_m�u�S5>([{w+!�Sx����(^̥dX���m��3��U��vͬ钃��i��`��WQp���7��^�����홝uʻf�	)
Փc�|&cة�NcXE��:��u�fܺ�9S��6n�SkS�˘�>2���D�ب��H�W;.�4e:�R6w���Ջ7��w�-Z`�E���㣇�f���[��И���n���Nd�,h�Xd�*�J '{ikkw!��ga3[;�
Dr4��ѣEΆeq��?lX�5���;����)�NY��k�i�����Q�k��:���u��j�9���K�*�=�x.���4�;�ޚɖ�Ɗtq��16�oLw2=iB-GyG�Y�b�i��E�dqV�����O�U�8�Wc]�ѵo.��a;���i�^Gٌ����v��.#�b�ok.�5��A6����Vfm�'}d�ݴ0���#	������b�]=7�����lSy��GR��,Z ߭�eqO�ܺ�DH�3���Kgj���G��}��ԥsݙ(�Ee	dVG]ia����e&؍h��LNw�vƗf�5 =3U�*k8KA-<%.���!��2�2��W��~�ZB�F$-1��N��-����o1Ph K���;�[� �h��}ؙ"�=��>���zy���7е�S���
�����K9�7Dz�eU�xz�=NVK^��hf�N��}q;��&A��]�)���<¬ve��޶{�}��Pd�	z��Ug��7�C28@9V�,�!�- /3X�1��qow�'6�vos�V��KC�Y�4�d�է0e��v���p;9;s{�	�ZՔ��£���+U���,���t��0+�n��2d��"�����f����Z�ErP�^-��%��`���~�bA��O���]͗�lLދ��SD==pe��8`���]󝷸GD�{K)b�q@��Y��Xliܝm��r�|�e&~��q*�J�(b�%�.��ݽ9���%�Pa攂LO�̩ٹ�ӃVئ��D�TlC�������K�����:sW��%�w>zVDc�^���D��,�n�yg��4�S�4��ޡ�k�@�ܖξ�����%֙��w�v���-!ٛ�8ݳo+QP:�2����;��{5[eᚯ�
�ǲb�ή�T�W��J��1�!����fT�^�+Y}�MrMrR��o���z"���;��;��Bm�Pq���Y�xZ��U�Z�#)��o�&��8��*I
�H4���s�V�7��[}�F�{����r�>��ݵ�����l��:�{�<��v��k7��wW�wO;���\˻.9���o�{�;h|����3�]��O;�Z�7>{������q�h�����OOo��_^>�������k^4kZ�N�:k��ؙ�B?����:;�#��n��u�^�v��Wn�ӝ]���s���{��G���'%u��|�g����
C6��=�x���־��}}}}}}}|}ֵӧN��� �q��A�b`����NۺG�����|y>n�����5�����3����?ٯbI����]u�'��g��o(��u��#�}�ߎɟ.���/K� �]4v]�i�=ېI ]wf�}��_z�F}b�s}|h��dr�wt3�JO���/��3��?����������iݹ��u�_2r>=����.���)��EO�\��H}�~��n�I	��=ݣ%�\3b��a����
c"�{�E~��$!!4Lə$��u5��~+���߶Wz��,�v���i�+�}^	 ��H�`SΎp3� ��ݻ��d�4/}��H��XI�w`�?z��B��w�pB&�t�v;���Sc�m�����L �X�ɻ��R�~��o�4enHal�t��a��,�PR�	��=�t2�����������c�����Ѵ�K�i��� vUן�u�s�8�4�%�7��;P�^Ȗ|���q����S��v��-�[0點��[���
�����-�c���cTqX�Rt�`��&��y�337���>$V������*򿇃p�YS���<�����ǣ�G��bJ�/��EE0-;۹Ԣ�DR���Ns����d?�Ӊ��{g3�)�,8��`��p0FG���[td�Ƥ%5�[�[ji̽#R5/���3�e�'��Jq��|�n�f��,.b���	ы-�O-Nz�L��i��[�>��N��qA�E�# S+��Ux(�|j�>xOB\w�+�)���r2[�I��v���<�����A�R箈M�{sޚO�SIR`-�;$v=C����5���dK��[_�����#��8�BC�^�;�gu*Y��0����"�RXsw��0�Q�ègUs��:�n�C�L:=���z/��5��[�o�7>�}ߏ;0i��k\�i�Bu6P"�]��1�o/|�(�?�|3���|���!��@�}���}�F��U	��߫�m/� ����B�� ��xg��,�k(M�]�\�_b*S��ӭt~�c��P�p�J�r�m��-�֪�ac��Rt��o#�gL
>Y���䙍��ܙ]�v�M�c��p��9�Mۍ��zge)��� �}~q�����}x�����/׾wk��ު���?&��C�cu�웎2��q��P����JM�6$=�;4��K��7�M@�L�������ʔ�[���WU��w�����%��E�� ��.���=?e����_���){`H�� ����w��F@��y+���|��b����\��K���|2E����4-��D�0��j/a�i����O�����{��)�=��gh!����z~ǋ�7� W�#;k�o���K�f-$�w�>݆8g+H��=������Ǹp#`�.�0v��%�D���!逴��<�]�P��@7�HV��S�Nff��!�s3����خ]�>���O�`����I��vA�g��%�H)�L���^%�V��vnk����9?���A�R���2�)�����Ӑc�P�a�_|����).�E�K�=u�>���>����?6�;�'Ƽ��O���z0
�5��q���z����Q�aс�U�[iS�r��o�i������O�|^���<�A��c��#k<l_��DC���3y�@T}���B�	)�/�sॼ�Ntw�~��/Z�q̄~d(v�D�������Ï.�񻘉p����o�f9U���,�$��|�]�WR�KL��� �PU��v��Zb���\�M	�j�;�3~��R�J½#�Y��W��e�#
������<�����U3�m�����.��M�TUnJz�Ӳ�9��n˷��k���,ڽx�M��}VXd���+��@�����y�����P}�Ľ��NR�	����h��0��*n�1vr�zo	禂�g�!�)�$C��j5�i�>�*� ���[8�Ri�ک[�J��f�����ᐝx���A���
���ag��{���d���VT1[��&�3�������=� ���r��&����H�A��Ϯ�mH8Z����)z鸮�h}Ķ�j���&˂�����ܮa+ג[���˔]',N�N�	��P=����G�:no@��q6����;������t%��@����y0��,(,��5j�[�����N���C�,�-��xɣx�oG�;�Y��ֆ�� �ӧ�0��Z�9.�p�9��iNCq����1m��<�n�7��38Cc��RS�0��Ia� ^�C�����/�¥"+���e�ox|��P��c��f�_�]�^�$~��(h`|C	�[��3�-�f��QaY5(�E���G���v�n����:/�lptg/<���CawhOL�-L���u�#�R�����<CJ�*l!ߛ�Q��6��	h�)o1{��d>&^�Q��.2���Cr��)?ߖU����O���bK���9�h�8���]�g��`|���9�;oxi8�0v�T����v�r�g
�x֫&{�O!���錬=���H�f`��h܁�������i:"�Y���������2�Yq�%��UDe��H���k�R��MW^�i���	k�)���PC�ϛn6��}�<������mS�\���(z�z��%�H��	w�� ���2g�#Egߤ,{΂W�]ޤ�㇯f�8�	�do�<��F��C�>�(�x �����L�2: ���#ϻ�SY�	�.�%��V�Yz������;�x����z��xi�=���[O�q,�@&@
G�h�u��,lF�Y�,�m�-��{����,9�$�[�]�{go&��{[&E�&o&�} ��X]e:*b��f����b�,�;5~`�*��C^\��eI*L)�/�P{�[Bz� ��	��g�7�ߕ�������^��Cj&A�Y�Q��b��S "��KzG�~�9��?D���q�.���Ԗk���<࿗��	��q��Z�ԯ�[�p㳼dO�b��XJ ,ip��0��׽�ؤ�f7ۼ�g{���!��0~ni�"��B^�{`-����+�ɗV��$��p6�z�E2Y����0k�d�lj��6S:���5Ko����n��U�9��+����lb r�� ������
w]]2�{�&�G(�{�e<y��,���Ǉ���E��v���]� �P�Į�0�з)������T����y�///.��������{t�B�ݥ�_������k��um��Ȗ���,(wG�.{Lzr��Nb�ެ�=��^���.����,����sߕ���>3����(.�"]�7�ݽ-ݬ����k�K�߫��K�q��K��(
<���8]��_=�l�5(wI��{��r�ۡW�vk�^ut�q/�������t������n�9P���g��=y�k˽�A����sk�qFj�:��
��˟j�E�{x��B ^9/�v�K��}�����7%o��"(�L���=�zZY�!�
O��rz����zi�0a�#F������v�7~��	w����?��(?WO��-T��!7�- ���9�����U�|��pĳ�S��ֆ����v�<�F��~�
��3��1עUuEO`C0:/1q�oO���s�xy�.�vv95f��,���B���
%=y(�l`��}׺�'���D���o�1�Ip�گ
נ����mSTm^���W���7/]UkS�\PĲ/i�M�������(W��JX�;���J���?�]߸���T�X��*�{���:���E���]�5؊��6�K�e[=u6��p���B�p� �;s6X�Qn��Y���Č���Jk&��A�;�|��tOV,m�J��	`���ދn��h�����?���}�s�N�#��\\?7�/Z���{�z!2O~bS�JE1IJjgom��ȸtul	v\
���܇�y��.��x�`47`��)}F};�J�b鸍�%�K�h�U�����[�a��h<4�q�C��O�����d1��ǘ\�j>`��=Z��q����'�Y���⨝���`�������y^9��^0��r�l#�(�v#�;;-}�����k46��]H�^�n-ݵ��{[��2~,�����x}�	�Z����l!}�>=��륵߬N�<�[��ݽz�2
,1�*4�k�q��qK:@���<f`^����fCSxX!���C�vbq4E+�F;s��[~x�R��f�?O/ᨻ���(|E�XS<Ų�{d;����i�6�
���¯���Mm>����.��jo������`k׺���f�W4��rȵ�:�v�/l�y�5����6���;����H9gh�:C;ſX����l|���œO@�f-�t�%	�m��<K뿄�z�d/超^�� �-�x9Ă'�+Y�_��돶�;���.E�D+��W��)�fs��NCV�U�����d+^~��>��?�؈���N
����f��	$�O������f�j�s��޸��E�rἹ U7U ����ufN�wkځ��1N��e3$Ԏ�r���X�o����ǟ������p$ڒ;��lO�i�S��ͩVwN�V$d���8�H��V�v-�I��x=��q���B-�9��oY'��擊����v���D�u�=�L�<����Ũr�W�2of�P��:y^�w�`��a�u؉-EI� v�;���k=������3Uʹ{�|l���	eA#X�=�q71P�6
	l"�r�X�����<�c���@�&v���[���82�BehȕҨ��5�Ƨ�`�tKJ0�q,C�0�',�����S	<�Ϗ������Ϭ/�O����h*���!����Ŏ���/^m��ow�q��czS`aC�`eu�w7�"{�Rdu��Lʲ/A���C�_�ٽ::D�DР� _*+�ȃ����<��.����z��>�Y��X����֝�CǺ!��R��QL��n�� �֗��������!�Z�^�!�k�Q8�]��TVb;��{9��:�R%W��f��� 5�e"�P�o)v�L��!���l�m��8n�'b�mFn�{s[��6�CF9���2��.,�%�Y�1�
�XI{mi�@�/|Ǜͯ���2S�Gw�lYO��:�\��SE��Ǳ㡙���u �B�<U[�W`8.}c�[��N(*I�0�K��f�{�j���]�(��+���ʴ�51���xs�Hs;^��C.�^A���pܼ4E|�]W-�/������6�z�~;y��}�oI��\�Z�����H`�
6��.1��
T�G�
��{J{kU sr�v���\r�����n)����0:<��lsH���ٙ]���&�{I�X/�X�̵sv�O��k���C�M�h�C)��!tx_=i�恐�F8}�[��t�I���_~3Q;�����Y�v��[�]��1�8�16�qvn��`@:"��o�c9p'�����yY���y'*��<�槒w�񷆼!Ͼw/"�'vB�Pi�e�A� [N�Sץ��_�;@@��.��(���i���ۋP��|��_ך�`',M����+��^���*�!\�y��n��b���-���;$':�߯}���D��E����:�]�s�~��k�"�q@V�3��T-7�����Nć*#�r���?�����GMek�����͎_�!r��K o�xH	���&F)K�vҹ�t��s�,���B�=�Bޭ����C3�[Jq=��*`���<CMj�j��0�ާn�����n�W!�:#�8ė��o�	*����{gR!���Cx[G�ޔ�P�'��T�=0��j�QQ=]g��W+�ߝp�#��1�bª����<�3._e�#E��B�V��B��@�
��\��wu���� �A"���|C@/ʏj��tv���WR�������ƺE���v�lll>ݭ�Q���y^�T���vG,m��O��n?cX�N:u$T��_����{%i``�7^��d�`cȺ�I,^��%���q ���S��)l����ջ�G���c�K�y�m@�ҟ�.�X�R���2��C����-���}�Tr�vKe�f��V]n�]�zc�m��@�����-�@��'��%���Y��Y�A��.ޓi��#;/�C��8u>j��y���C��k;:�B�Q-�k8��7�o%�wغ�2�F���u#7���b��웞�#�[�"IT_g1f�In ���s�<æ�{���&a�P��vv��Jdu��D\�j��=���j����8�U#5��s�{���~@@�>߼�D�����" ��Ise�C�ܱQƁ�^5�[��Y$����c�,_ (��K�ď]���e�Nb�����b�=Ln�B^�[�W|Vz���ojJ�h�~���<������mmJ�u�<��50A�q11��^�����e[i݀	rE��w�F��E�^���\�+�������ԕ�i�B>�=5y�i�E�^����#�w]Bw`��WA��h��B��Fm���vm2�2a`�/�+��˵��CY�S�s���_kc�;��z�Mp��MEޕ���,��D��<�YGu�jR_����υ�g�a��������(���-�Wϒ�T�V��J������y�yof���[EQZ+6lH� HHI$��$y��uoW��g!�_��ެ�O\�n643� ���HR$���c�a����K�"סw>�=.��F�=f}�fŰ����6q;⢏��s�'�� ����x� ������nD⽸|L�y^�<�����֥�<�j%=$gP=�m4�_-�'�P?@�@�/�5m�uOտI3/>��{M8�`l����>���d\�Fi��@*AGc�y���ȷ���#x��$_ZP�s0�C�pjcXt��O��s���~s��R�~��	*Ml��1D�֬����R�fC�qI�h�����?!f���#\�i>?e����+I�<z���>��=ߜ�1�-�;�{'��iv�^��|�<�-�y�"l?��Ǆ�P훑̥�i�K��Z�[�k5?0C�\��{S(������7W��,#���m~��L��
�-�-8��
����g�Dx��@�����܂�\
�s�,g��q흼 ,��:�t�u��Y;�]���<Xp9L	b��Z��Jq@,�$/VϠ���:y��#�7�&zgf� rL�����E�%����8�B�I{��Wf���hA�=�"�m�/�"�B�K�@���w%_<��,T���p�{y��
���ā��΅l���v+��f�9��]Ҙ0]�� q4��@�K�jaB|Uǐw_�Xg�=�c�l�i˸�d�w�V���VF�7YJ
�'A��x*<�VE�݂��j5�C;�\�n��K��e�ld�ъu1:J�s��zZ�ӑ��Z.�҇O�U	Ze8�Li�m�s��<N^t��uǺ��T���w��Z���2�o�����5���ы��]lBힼ�8��ڪ�y�o��Ln���[�L�c���5r��#��U{���@[p���䊦�*�Xh�^�3�W�UMmѳBKd�3�]t�sm�@UR��]x�-q�M5;u��;09ܵ�Xr��o15�2���}]o�bZ$Aq%��y2J^\���pu4����_rm�u�ۊ��KV���e�sU���Z���x�׉&q��2(X���5��o�7����}-3�.�[;%ֆ�E)5ي���o��\f'��3�ـR��Hz�}�N.un 0Y��v���y�zͪ8sL+P���!��ė3kNi�T�4����oo�*���oo<WL�F)���ǋ�>�9��O
ܗ���ͳ�G|U�1H::ъ�n��7�n�=8u�Je:y �=R�e�K�(�]�;A��%��yE'm���'O0�y h���I�Y�JP�n�/�i���lՙL�T���Czщ7u��ėyB����MÉ�V���e��Jq+Vek���`/�ۦI�J�f�|�>��B)��Y3�W�����L;���<��;R�u1����7[�b\�Ұ�n�5�_5ͅմ�7�������o`uT*m��s�pҹ�{-��DfBU�Α#fB�\�V�霪��о�t��͍��J��޻ܪ��U�'���6��+#ΡB�+���Q�a74�,;��(/]�}Y��4nh��3�݇�0n�-y���upP��-�r.���<����j��ұ�V+�[��e���l�����ĈN�Y֞>uFw��N����S[ٹC�:$��B��v�QW2���Ǯe�8b蛳�F�������-�5xg�O#���DZ�,.���t|)�dUD8�9���7��z���Ao.�e*϶��Juv��lk�2��=���l-:
��>R��W5$�zy�c[�뛀�JkEQO7��T�����)��4;�_�q��p��R��8r��ðr���!{Nd��\�!�l`�<���e�*����W�./;��7��j[�_)����U�Fʳ0�+`|�q�DYe�%�����l�W\l�;A��֯\��X�]R�]ɺ�튘�T�u��&�YVJܒe_��`��w>y�&iRH[rI���(�4囩��~~$�Q�AK�Ő�
D��|n��W��`d�O02�$$�D�O��^>���q�kZ�����������:t�׏��!����3����D�1��7.���>��$�v������צ��5�kZ�Ƶ�����N�:}zx��䄒L����t�Q?��|��盒���.pK��r�JH2^� 4h�����SM�Q! ��B �	#t���L����C`�wW>u��L�i�F��/.�s_k�_��!�������J1&r����f�\o��z$00��B&���C��Wa	3�\Qi^�$Qˈ��2��"|�I�E��ؔ���i�Ra���}��YR9�!	��h>���re)��H���>��y�3d�FBFB	� �� �@)�2y�K(|�4J0�[A1�|�D�'�0cL2J��$�-�'� A�E Hđ�J���.�{5P�V�tw-�^��Y}���U��Ҕ�����ɭt7�EoN˚��6��Nd��9$L^VS@���h�D�n>L6S��!#$&c%�#k� �1�h@YEH�-��A	4�~m�A@L$���A	�$�G<�iƒ@��		���0���!3�����.:c�J ��k���Ws!����[䜧���+����b�ZH*K�L݁�]z��~d!�)��zuNҮ�GƄ}K�Ǥ��g���){`H�=�	va(��?5�w��q�=��`�D ��D:m.z]��ّ�/e'`�M7�, v�<עl?B"��V�ռ�����[�w��vy";���*<B���\���f�{�$�^�tVB�.�Vh�6G�8���a��yOz������B3�1���^j���~��s��ƨ�x�כ[	w��>סHg��0 �%�8��o#.��5�=yi�������|������	����)�<�ө�o���u�K�7�Oz</b41j*�����^�9�3��zw�`�y�Q>wgt��Q����{�Yp�<����-�Ͷ��klЂ{O���rc��.a̖�������uf��=,�!@�"q�Á	佲i�Ə>F�6��bE�B�z���%ֳ�6���]��,�M���?�A��}煰�ޡФ\8	>Gd���M���f%ؼ'�y�K���0�d��Zx�oD�)��]���"n; ?�:a��}�|�y�OS���{�u�k�!��߂�\�Ƅ?�����k�(<̪P���G���`;�~���t�NkP9);��wjf����+�u�Y���hvDG���Cd�Ym�5��{/�:H�b��'z\3Wq��A�Y�_J׆wW�x} Ӧ;t鎝**�������;<���(	�*ۤRz	B���*�dL��������/��4��k_3��{G�xK�j{*I{�2.�?�e��0��\���^�A���ə_�M��3��I����@f`�v��ݎ���o��o۝E���yj9r���R��'���F�>=JG]t�uw�w�;����0����	y�5&G_@\V�TX)��4B���-��I���m�X-�#��3{�;��0g?2����s���uC�T�o&��F>���%�_v�ek��c�b̛��#�_�M� [�'�s=���g��8lN�̫=S�^璡�ֱKLwf��T{{��g`��Q������5P�<��W� (�Y$���о3�o���3� b�!=ai!�y,1�|��3rZkW��S߬,��@�x,y�3�Ƈt�7�#�H�h��ε�[��r����SZw�e��_9O~V��?X�O�C��{�<��fN�=X������c�����o��6��������S�_����~����oKW�`���B8��H��t�o�E
9�6����ۇ�����ߗ��'��z.n�2���Vν8UJ��1�C�:sZU��{�t&4c��:h��e�^�Mi��$\�d^���]%+��t��}6����L�xf�����X�YPL��>��@�+��@�:�7+���矏�y��t�N�T7�_|ݿ>u��w�f��u����΃�
�=r�z�OW�ȶ�JE�{��[�5 擜��;&�vY�~��P]{0����_: '��6��q��*�H���� ut�7�Ҳ��H�������R{(sT�U�b��TQc��f~B.69�y�8ݻ�Q�3�-#�w�u��	��弋���~��zun�����&��a�����'fk;dTo�N����\���N�CH`�B��8�,�zOG��t�#���{�ec�aO�m�aA��OC\gfkD[VmYI���Jq�)��D_�<�ǂ����]0\�Qu��L�-�\ۖ���ڍ�f�ݲ��CӾp�٭�̃�m� @���*�S��1�^�iN��X��ğ�ő�ܷ����r�Ѕ������g�����>�a���4���,2���H�EQ������^�̜��:z��b�ڱ��\v����;�^���=#���|Oں�ԣ�6�����P�!�qYp�f�i҇�؝�Ms�a.��{oSZ�T�צ��`1�~/0�����>�M[cg0e��3YsB�Lo�g�/���f�sځ�)����z�j����k7r�n0B���B�@>㗦U�e��s��#�'�V�!�1=v�Iu��[7]\����@�;$���xXR��� o��<.���} �X��1�:&Q��6���I�@�����<j|�L�u�ގi=S�#��;t�g����j6/"�&-ʣ݉�.�� ��	vՑd/�[*��p_���v�g�0�����f��駻s����D`�᠞p�b�Ծ2U�#�������/`� ��m�mW���kU�]����S�� ,	�����KA��D\vL�����kc�Å�zˉ= &��b6�6U]��|���o���%�M�_g��[��yg^P��?���Ǉ�2�$�)g����\�^����j�Ś�����/7QSm���9A��kS�S:�>�[@��<�ǥ���ThQ��h���f`��Ἄ���Z���ɪ�Jp1l4�f=[ռ�n��Z`=��m��y�yHjaJ ,y9d\���a≉d]#��U�T�����9�=����I���D�G�u�=.½{��>ܞ!l�qX��E^ε~>�0�#��ؤ��-�ci]&�j&�Nq��]�m�og�ʀ���Vc� �r�X���}WA�Vߜ,�\󿄎�T��t�5OD�9�۸�7A�ǁ���L2���"��|w{>/�DF�B��ܻ����H�"���_@���S�C.�h�1�7�WǮg:k[k��`�@�]"��7��9:�=@�#W}�q:)܂��A��]#��xOl��J�.�)���;�fj�Fw�<�vJz(O�t������ ��k���}�,��J�:۽[���'n�lg!�4��$:��sb�t��mR`Z\}�=���!��_����E����_���F�f~.�'���z���n�\�ӥ��ÚV���?t�'s�vC����9
�^�,���YZ�q�x���k¨vI�9!1��~JI�E�C8��GC�}g`��l.F�$7�MvϘ\���=o�τ�rڌC��m�@�����W>���q���1�7NϗN�O*��զyg����!�^a�9/@K�dق����#hOOد�t�W� � �Cy�:��6t�NԦ%�nٰm֬�Hy�;�%�A���C�"�.��lφ^�O~n��4�"k�9�.�L�����W���~u�|�Ʈ{�Y�����a��hP!�.߬L�%C$6<�4!~��_
�U9�Nt!�/��gC70˿B|;���]�#�`�|�3E�2"`��zkN|{��N�&92�v1�C�T^ 3�����_���<��֩��� 3^!��\l�]���2���WC�n[-צ��>����
ʂ�_9��W~��nff5~`ƙ�TgN�]�/�P����+sE�j��Z���������M��Tt�bTO'� ���+G��wϑF��!�t~�L��<.�V���JCz�h��z��fN2v���d��0�R�V��.���?Yk{��E�9���M'3u2���� =�{|}�������7�� ���W����0���A��ݽ0�E�J�z|k:OV�K*	�v��p��"DB�����p�CT��@���A�ՁO��4�M���hb�c�+p,v�cBѡKv�MɃ��%�rou����/-!�x�&i��C���"@Pd]	��}n+�&��Mm^}�ļ�tlrی��Ȏv�5!��{o.&Au	��|ճ��7#t�z=!퀄�v!��kpi���j'2�f���ջ����q��2X���$�	B���f�xay�#��vI�D�`b6��L����G���t_���}P�7*y=�b�C�&��6�MsӸmp!ޙE�A����OS5֢P��wwfv�
e�NC.y��V�Gp�>��ُ���R˞'сD5�S����L_�-b履�bm������	/ȅ�O�C㼪)���רu�������b�gG1���~\q9ጛ*{of1�=��,���� �ƙ3�� �7���H�"���qqrzW?	!�t����Vq�r�֦谏��i��������į��(�"2���0L��[�``>q���8㡻H��K�e�?X<��fY���{�Q���1RuacW�3�ؕ.v�K��af[��B*[� V.\$�{����l����L�l=��	ʮ"��WGu�r��m�NwR��)��ƺDLt�N�N��:��{�!��,᳨�_&��qL�`	����[�`?������&��Hy#��%[�ɝ��x�3Ӯ ��+�ƓxX�O@�3v�<tE1��-��ZF��ǐ0#lX����j�z������GX�;9���$4^;/u�ܴw��~&�â-��^�ZŗQ�.��%܇��2@����c0�qQ���	z���omV�"����Iʨr�k�ûi�	Z3�5.?.��������F� <n�V�ߔ)�a�yx~�� Z��ݕ���;��m��0ޭ�s�b���@r�]���#ǲ�Z������󳌁�uOwqL��k�NZ��s��I�������h7�U�v_8�Y>[���дk�7 �ݾ[�yn�c;B-�'�"#�����r�Tl].�4�r-���gY��-��)��PX&>���s֡Yh��J
�Rp)�eMw<����xkp��]��C�mݘ�p1z`V�ځ�}|k���t�"�-yb�T�Pw�5�{���ghyh$��q�U܇���q�s�^��3�X�>��_Aw�Ȣ�)�]clLN���n���̎#NowRC���F,�LVr��9�B�^��N�:�8��-h�^���&�����B�5�O�{E5��b���Ϫ�M�T��N�v �y2��]�%�t�>S�فS��y#R�Ielۅc{B^E�I(o1Ħ���>�S��N�G1ӠTL�#�\.�J���==��zh������K!���Bm�Lx&پ�&��;��/����l���FN\�j���yq{lVg��ܿ+o�=��=�_6��8�T�0֚�F�?8�vkLb�ǽr�t��쀇�7���\��P�z s{�^�{�x���;܇����.��ϸ�5�N㱿[wUK��9Cņ�Cd�	�q�*\���t��#Y��φ�W��/�`C  ���
�Թ�S�����z�f��vf�t��6Ѝ46��>�/�	������=P9�3�nߤ;(���,���=\��[y��"6�.��n���(�����ԕ�ѐ���GXn^�j�Ku���|l7v��L0��'�pb¼��	��U��4S����Clx�[m��$�$��;a8��l��VU�fNr'a�z�����u�3�$KA�ɒxi�MǴ]�P��ٮ����:���p�=�=��c�}��=���&`��	��|�	�����1��(��V���9�=�,�{�P��h��	�H܇�����超]>����~�����#��9�n���`q�?����=��]����Uc,D�ą��yo�G��G.��挮���Z�a.���G�m��A��W�F��E�����\'�u<���#xw7{�yԼ�^�����?N��t�8Ǜ�����=ᣋ�9�A�e�xg�ՙ���2K/E�>qrB�%���B���|=F�;����P`v�`O�r"SY�L'���[�z3���ո�?WE;7ms�V�}ZW�cǚא�aR"k�p��P��	��u.��e�R�
����,�k��=t�vC0`�Y��r�ޑ��E�\:au�^m{&ރ�LOnbS�	H���������WY�����t��������?1�5���#���M��� $��t��=G&��ww7sU�x3�k��&�ΰ�cג�'�vk������?����fn\S�+\Ӳ�t�_8��y(��R9�iyz ���f�lOm��7��Κ5�����{�w:�wj4�j�BLK��Ad�yop���J;��c8�^��adR�X�G{(�qń��w`�}�{_�~�,�C�?4�I���]�It�Ύ/D+����H�zw�\�%=^?O\�ʷ���y���2�����8���z]�0��Xǟ��RA�#_*��S���~�ӵG���&��1 ��T�4�Y�q�*�; �A�@Bs"�vO�,����㬿M0~�^?�]+�b���32ؑ�U,��k�Ώ��e�>&�����T��ه���4�eD�4�(p�G*y��gQ�۽�t3k���@��Qd+��9Ȯ�@���͡N��DM1�s�]_eg�� �N�����n���g%tv֙;g]\9�uէ$��(����n�G1ӥD��_=���y��/4ω�}�|�T��/��XHk��\2���ƍu���T��ƿ'J�Cs��m��	]D�5v'����\s��j�0�tE�k�9��.���` `������7"��O,G�xk�M���.����+H>��a�� E��@A�Ñ�b���M���Ǖ`t�����G��:�Z��>Z囹����6�l���[��^�-^*�H�/)�ڃ(���������a�L��+���� ���ֻ����\x��h�	>6s��ځ,���}�z�O��*ܮ�����5���az�_�� �O��i���hc`?k�`�'��&_�e:���9�ݮ'ӾC�f-��L�;:�;jP
�c�|�������"{�F �
�M�U���[����eu���t�%8e
�)IžŰ�ȶ��1�C�@	�q"�y�.�{Z���/��ϐ�����7S�����L����)�$MxP]S�)y�?,.w�D����W�OB����B�pכq�6��1����X�&���i�}w�����B�p6ض�b�CS/�f�i���
:�f�$I���N*�0��"�GE�N�,�Q��q�֎#�.��wE���,��e�<͇b�#ai"�Ɔ*sU�oN˨�1M���8åǴ�C�#�lcxB�o��V��cFh��&�����Tؤ�>�	ZGQ���&y��7��R�yuE�f��A�IW&G���U��1�����6يڇf
��/v띫!$�/q\�o]=��o�����hA�'��&������F)��0����(��!t�P�:%��u��k`���%�b\�u�9��O��)��V[累�4����M�u�77Z��{�H��fZ�ud��e�B�!ӊWn�����S��Ev+��p�gE�x��n�](3N�f��v�i�;��Ď�V̮`ۛױ��EB��7D;L���r��W��Q
3�+��I��h$Iqٌ��׳cѺ�;e�\+aVqj7"��1�{՜%�Mˌ�x�*]�(�Id��������U��(cAiZ:.9�c���wt����Ӯ��E/'v�3L{��h������	Jt�)��:��I:�ln9XU�W�[{oE���-ؼoFjQ8sl�UbU�5&��y5�o
'p��:>ï(!7�wX.�푏b�ȝFp�%������
OfH�:�X��1�P0��ΗT�#O=��� �P�)�=+��Ta�Y/~L��<Ǧ6����#�҂ea����Ǆ�FY�ְ6k>c)��K�-����Й���D"��eo=X+s8�ڱ�lf��VM�i���n�Z���,��JS-�w;�L�J��+�YN�%-e$���Gs�ڕʗ@���}v��d�J�z{c�h:u��B6�7���޿�κ��Q)"�k��;"%�����������ڤY<��������4�״2\��.�+�S�ȅp�T�bX�eg�t�n��.�rp���u�wF�5��u�M���N��9r����:K�D,��t�2_���+����n9nJ5U�\=��U���N�u�gw�w*���Wy)TüDPR�첎bVu��][y��\���·~�(RX�ӵ���������8�*�]aJU6���Z��'t�2���[VӦwmi'��j��Ӵ`U]4�4��;n��ⅎ���\{Q��uL�^X�C��A�W��Q���vMH���.q����
��=�m�J�6DB��[w��e����0�(���-R�zb�e�T7qr���]�AM�#������p阊���ٵc�#ر`�ڐM,��e��w�D�[,�$I:�79"�ÜԐiRHZrL��m9W��<I �A �A �@!�⹅��$�43 ���#I��׍}k�ZֺkZֵ�k�k��ӷo�O�0�!!$���v�{���?}�BC1|�x�������k]5�kZ�ֵƵ��ӷo��<HG�2H��I��31��v"��d���Q`�Eb�ݮ��_�?���c���V��W�$�f%/:I����iDi%DD&I��� ^[���h	w^��_5wO;o����AD���0��H>�A�BPؾ9��	$Lh�I�2�{�k�˚R��a�F�:,n�P�{�I1&�F�$#D�7��a}���5��z�����2�"�$�fNw�� �Ѿjr1E�I��%"0f�A$QM�A	�g�0v���Q)�婄*Tk��(Y���w�fg3x�����%c����Nj^6�+sL�3Re���۽'�~���H��8�D��^{o�7m�B�O��SO3�
z�-�f|'��0���,r���Ɔ�N�u�2�wj/3��]��yջ�'��˟@S���t��[�y�i�K�����x���*�
#��ƻ[�'�n��Z����l%��/sӼc���#[��3�*t8�X,υ*|Y�L��8��љYݽ�W�N��	_��K�xo�^��%��\+�W��� 0(-?&v�;����۹�n��Se��l9���l�Mc�~&�~��^= ��ރ/^���Ah_��[]��G;��%�.ob�y��w� p��a��_A0ǵ?z�{E3�:� /-4��&���u�SWv�0�3!@C ���!��Pk�l�c$`�t\̀g�r�?1���G�j�c=dڜ�k)��`�S���:�xkR�Hv�!��<��I�Kս5\z-��s�-��K�U�kpƮ_sVw̥H�΋��;/2��|j���6��
w������r�&|`�(�P)�4�gT��Gs�ooޮV��u~;}�����o:#�MutW�5a{�ZD8�y=�I��D�]��q6)�iᵴ�*���x��l�T�����*!*���d�/4m�Y�qwOM,�L��M����_Gį�I}���d��Nr�Ys�S�N5�eR��N髌�ʂ�<�E[]���988Ϋ^oY��}���wצ��ys�0��D~�<qҀ�N�t�"y��;���9�9~=y���_��U|hRxF�{����i흡��k7t�3:������1��vu�H��LJp���L��IP����ƨW�4K`p{y�xu���|��h��Y�)�����<���\����<�z}>a�&��fu:�1,���TT���.aq�SP������+�����8p �vL1�C=!H�]�(�c�*�.����`i�{��Mr0x�ooj�-��w� ;� �P~�k�6Ⱦ�&����<(u�~{��(�}1���o�:�ze�*�]��/I�%�v�}�������Q4��:�,5���F4B�TsY��k;�d;����җ�#X�{�w*�x���~�~	���sh%����}�E���ևcw9�wv3���)�,v:K�q��iA/t�Ǆ h
����s`0b9����ad�[V+�kξ�{]C���=	vmǟY^�epj�7�����rLs��nKu��0d�7����A�&�N�ɬ��]�䋏k�VJ/��Ki"eC�3)Q��(����:��x�3{y�ib�uܶ!ɢ�t��tJ��GWm��֩J^�v����yγP����y������S*�����Мȼ�K)[���kR���ۙ5���EYKc㧡t�e7�8�<���H[ړy�V�4���Щ��k��X�ӎ�|�������]�k�G{e�j���5f}��ִH5�Z	G�i�%`%����b��ca�B��,�3E�M&?��F��ǚ�Ϧ|���S%p�Ϫ�C�]��%�%�t�v��}ao+;.�z47���7m~�p��@�Q"�w�?�fŚ�5����;,��k	}G����9���8�0�08-3�����0��m j�;�0ջ��Nϰ��s�f>���^�u�M�С}�Z��&�$r��ŧ�{gS�)��Ëc:'Xcf󆪽9������:�w�� b�Q�^�q�)��5�U�����xW�Fcս[�{"Z�Q<Um���f��L��Y��@�B Js��Z��7�xQ1,��	�V%*9{��߬ӫ�V`�t,����'�}�V��r,����A ���y�(���W;���Q��&I�΢q�{�b�d�����I"{�9xkki5�����^��:<��c��D%"@���EOG�*�]�(��\Zc�+�ˬ��q j9ӨLU�H�IQa�K�}|�灱lO��"Su�L�:��Dӷ"�O[K{Z�;����;.�,e蘴�����iK�����5w�S��l��[������aG��?>��)ebס��YW���	<��7�$_D�2��z����NV��RW�}��A��@��3��C ��zφÝC�^�[�I���l�3S�u�]زr]
Iu�7[/�G�`�}b��yv6f��"��mMy�ݻ��J�۷1ӧ"�I�� ��qK�q����z���~��U�'�h��^�q�e��ן�b��r�v�cV<wB9��;.扺�7�Y�O:�A�w ��P�Bǻ\n�t��Y�����} �H�U�5��Ïʾ%O���w��;�t�d�'��qxQ!��|a  �;��Ӣ�/����xZ��4�k�}:�8�����E����Z��77�?�,���,{O�ߐOBA�6cp�-p+�\�I.8�������c�w-`��k�sI~�-E�;�� P0��b��?*��5�#���mN����������{Q��	�vnb	�a��/ܡ^ޱiTQ��.��o_3�*�fww6T��UM[�DUL{S���-<�y�e)���T�
�d�9v��֜�S�͐�j�^UC��L�(+b�Dc�\[j}����'�s���Z��A�$e��^Ͳ�ʲY���pFФ���t)�;Гۼ�qV�ϡ�ޘW��.��o@�	>X|�A=P%�܌k���YU��J�ݝݫX^��q"�*7�������X�.$xFz'���5��<{6H>j���e��;�|�-x"^���[qU��N�Su��ne]�jS��+5��nȝ�=��rj�}�����#MBb��E� �Ò�Lywf(�'6��.����������Wr��;��g�u��,�Yo�$��>����D��8�	@3\�������<�|���ƍ�9)zم5�8�:��柽�DSzS~���8�7�}��Uku��j-l��L�ߜħ6���BN+}8�w"��oD����8�=dٖ'/c�^�8�6���d���4�`c1Vt�O^H����=��O� Tu8�6�Fa�淼�L5S(r�j`h/ \��,�N�;?�r'�߉�M�oZ�M;��m�\�aCU�Lm���=����D�f�^��Z=΃w<2n�;��0���-@�E�(,H�{�ۍap�Q�_n�h�;�v����ލ��,V�������yP��6x�yg�$d�%Ia�&�tƝ�]qH��V�H�L'������C0i�'��k�- ���0��Ex��5�[U�lv����U�ce����
ʕ�eA =���j1������p�1���<�|ų&�f坹�@Wwo3P�Ùz�����^�'}\���y�l�3�!�������8A8��r��x�O��ٯ���{�[�XWtIz&�^�L:"��@�r��8��P��r_��H1�T1n[�uu�g��2B��] l��죝ΐ�|I��7} �H�F]��u���UD3�8�t��\�.��VzاO��gs,`�ٛ��r/��]�F_n	�ܗJ*¾����;�K;�ռP�{�����w��#:q�*�����N_��]c�zϱ��F���R{�k�_�z埿f�	
�E��#��ÔG.�Ꝥ���� �mބ��¦T�Ou��N"H�.&.z�oMl�oV輷_BOSPc*!nm��gs�B�4~��6%l\X��]>M�0E�A�qqw4^ĸ:jw�l�X�\���sc���d8��5 �2q��l�	1P�)���v�f���Vg���1�|�d�W^v�m���Z�@L��g��O�U�
���z���T�-����u���/�Ygut!�K� ,�>��j�j�Ijħ6��	�T-�.����~�0��-p��mV��|��-��u:!�4t�ѷP����b�׻�u�bY��)��&ٴݕX�Qcd��R�p�Q�O���`[�a�p��]!M��y�tQt���.�]u���w3'7�8��khu(8�;�ׄ��������vz1��΂~���!�4���Ow�n_^�r�u�-:k(,h.���^�X�al��!}��MO��c�k�0�;�����9�I��m�\�*s��0:�\�ͷë��	�
�!�r�+KY��3E,΅�H&��p����Q&�f���Q5��E.�]L���梕����b��b<�W]E���`k�Y{(�O{��zn�_B�՝��"|z}q�t��J �������uͬ|9\�'@NnN0�������Ȉe�<}�p�wUl3異��W*ܤː�5�ׂ[��3;��8�~U��q�[C�v���O~)]<�]g*�v����q	�-����P�W=����W<j��(l[��5�`{�wi筼GT����A�^Dg�����-�Q�d���Cy�S�1���}nځ>�z�3�����gu1��м�3?�1���y�9�W�?,��	�Y>���?Cp��n,���0
�h���3�ۍ����E��Y�c�4_&������;�����Oech5����.�6���f:y�:��i�[S\{:"��{bY�k�Ѕ�4��'�Kսc~�s+�M�`~̬GK�r�NP�ݞa>�S�b/�y����/<��v���r�ԇ@�L7Q��+ޜͪ���ۢq��n�=4`����T/��C%1L$�Pz�l�z�Χ�S��͵�J�fB��B� ��<����Ql�s�$Bj��5���3�(�f<�7��l�ws=���)�]y;2ߒD�2�8FF�ߔ�}�r��Ԏ��ApK�$�3L�j��D��,,F;k�Py|�x�o�H���q(����v]iq����s��J�O'��?�v���'ă�DY��w3o���Y���K��L$e�@t�P��JY�q�yc;Oc�)[��i�����o���^��V�[>��k� @ӧ
oxx
¯'�e��^�/~=���L�����"�@,���p�z���u�d�}&��j�im$et�k�^�ǵ�2)���+M��+$Od\:��?�Δ���j5�"�چ�ֻ/N>���v~O�6�s�:b�n�J�^�f�XCQ1���<�lO�D&�"��d����k���PmA@�y�.ӹ�^��O�({���cX�[/���.�XEl���KM�CM��2�q0�؞�ǌ�m�;�+�h��^���2�pY��ή�x�h��j8��wk�g`y���]C��^����6�n�5�t��t�z��|�ۯ�Sc$�����7~�͆�M�Z{?>Î�`�6��}���xml�fE*�]~��y/x,��<�[*�ӄ�'=��?I���-{h$w�
пx�>1���͟��i&�x߫<�yӡl����W�|ҁy�aE��6��u�k����g�DQ�>a���ο'�0��kZ�\%����wL���CF.����B��>�NK��a�7�W=�l�;"]� ��p��l݄���|��v$��
#ml>5�>�y뗕�n���@ܢ�ꗀn�Ɏ�${3�vñU��&f�fQU"��|2�'��_���\Fn]�)�oM]��}�S�V��A��a�˝ǋ�4e٘Sږ�/�T������|��sg�?Mt��ӎ��=�<�$���V��=�5[w���OB���y��Ѝ�%��4�F]��kZ{�<	�><m�n-qܵ��t&�3 �0&xBa�-���n=2*)�7�/c���Hj	^g,�؊��H�l��׷<�~�P�j�M*��
�{�JD�=�=����I�|��'��e�PY\b�Dq��Bە��g� G[������P.E���}��w�Mm���M��4��;g_R;��z"�:!�:**M
P��5z�Ol�W�T\<��э�oG��r�C�󵜥�ؚ�������=܆�;d�o�� �/nbVz%~�	�$�s^�P�x_��x�Aa��d����Ԏ�����%˅�Cd��6���"{�Re���[t�OIB�Ǻo�"/d��jZ�=#]Vfr����ˆĴÛs��q�սN�7*y=��|���s�`D���`�d��9�]���YP��)}m|�	Q�g��.���"z�:���y��nRv<���u�Ǆ]��Z�"�~��)���̛j &�s,3�P�dȻ����>��0�/�,�_����<�5N�;vX,҂^R=H�k'�+g�kuPHU����2�I�[��c�Q.�S�����}�!�Qq�{^n�n?v�j7M�E��}��ՙ�+b�3nt�l�_"��7����3NWj��Q��$t���ǒs�}�~�:v�c�N:E[�����Yٝ˘|5t��+��턂�����1m��� +��\K#AV:U��n�:%iq�R�1<�%� ���a(%��"Ǻ^��%܁�|J�������}�8�!_�3m�ow�(�k��YPXk`�&�_���=�v�49�8,g��y����9�^5�2'�;4�8�>hDD���V���f��D�vk��Eyœz(f:�8��)�g6����vAm�D�!l��TS��}.���E�9�*�'2Gs��(6�<�3OɆ%]y{+;�؝��-��6&����_��$������];j�V][��˼�t�{}@	��S���Ცg*��d��L�0}�}^2������,��]�yI����{m�4�&�-�бD�n��;:�܄��2-��41�R��8��c�gU�\9����B�z�f�"�#d��Bi�kf/d�u�����=zѡI�	G*���Ѻ��Wމklgcޔ�>ݚ�Ô{�i�q-s�ڣ���:���,A1)��%%�j�����wK� ��}�ś+���������6nnE�2�y�EX�	�J�#�];˓��xJ�+�G��=ƃȣ샶iOU��p�82���Q}X2�V�]֦�I1&��\����fY|x�{���u/vy���W\:�w���R�r����V��/�{��K4ֆ���ײ���Ƅr^��wt�FB�|��F-����L"`Cu�Mp,Z�����u��5��pܪq�"�P��s+��8sU;n�m�۬��n]������%�d�=�kNQ(�38X'. �b%����Z��\>��%��[Τ�K�uoz�\|�,ɍ�]�/E��Y&��L-�7{�"�U1�0�#�j%�^s�!���;u�� ���^f���սid��6��	V'����+P�I4��m
;D:T�3�Z�d_�;U�O,��WYzbط���l�W�39�2 /T|49kB���k�JZ�*X�7�]2�v��#2���ِ�#�ѡY���tB�%S����������2���V&��Gx����}����n��U-�Lb��j�lN�;�1cg���](���]9�6ܐ.��f4֙]��<�Ө���-�X��y};�A,�7}OI�j�.pL�FVg`=%ś��.����"�R��ݗ��v���o�+Ak�Pf��`��{�`N���)�髯M>zc����sԚ�O,sj'��3�o�y�����zιW����B�>�]	&'/���JoMܬj���dڨy�2hE�+Q��z�̩Xl������{��ݒ���BWg� �(݈i\c��Jܗt��^:;P�)л6A�:�f���륅��<H̐�����G��=c����N�.����=��l}Ԁ�����Ħ���9�..��Mn����\�h�	��YYA6�Fx��|��\f�,�������j«�hwU+�p�U34��Xۈ>'���akl>We=X�`�4����:z�v3���2����c���ve])�#y{ra��.uB�+o.���4����k������Jf���۵���ۛr]�ڸ�%�L����`�����W�pu(����R����Nn��2Fr���x��I��L��ஊ�i�2dm՝�.&M<J��:m��o�v���fu�RA�M�v���e�;�nu��|��d���ɰs]�7�&���GmI�
��kl�;2�>�bjJf���؜ÂG����G0u�����zq��[�y1��84�P�wp��Jȳc�mu\ø��m���nw;fp������N��[{\�r�2Iv���>V�������rNޭ����߿?/�}��<����(�"��g	M � @d�F:t�׷Ǎvֵ�vֵ�zkZ�Mv�zzv����$� F@�_�蘦������&�$d$;t�����붵�k���k�Zֺk�o�N�]o�����������˫�&o�����&��DRc]ۄ��&TBZJf�+��J0flI�����6�JC�G�Zy�ϭҠ7����فC�u3BfE�=ܥ(̢H��$�h����"RE���Q������b�$��D�*s�^�>8�������H� �E��ܦM�$XMs�ݹ w^�d����PתnQ2��c4���>5�<מe�Gu�B)�$DD�K	e"S��(���n�p�anK�A&�,4�څ�T(�!�B�!$}a�*P�٘�E�p��fN�IWs�����橉̗�1����wUrmtOK7�k����Ҋ�q�z��Y�y�\5���4�#e)	HDQi��E�Pe&CQ����H$I%��$�E�@�#���AL6�4���(�Z�M��%�d`-6L-�W�I�	S&���|{q�GN�t��H"燿�<�X艝7����}�"���!����]U&����ծ�F����_�"R�!űd�0L�o� __����R|�1,��yd�wiINFѦ;��z:ηgowЏ��������\� 1��K�0���]!H�]�(�ay�=�3����u1���]�)�)���C��9jw��w���������`&�0#�v��wT�k��^r��N�n�w���Qi���Ao�s��?�����/O�����y^1�"�]���ڍ\��zy]&	�i*�.�*����3�*�K sH/Nb{c<Ѓ��o���_e̫j�l�����?T�MW�f�D����a^�R��(%�S��FP=8×Lc�qԉ>��ܸU���A� ��c"Ht�a��@�f�y�tS*�T7��=N���Ls*�u���::��SvooVJ�ې @f@�y���>���C���@f��l��c�=-�{�@ Uɗx3{)gl����x7�}A \p�y�u�v�xw���0:.'�*l��_*�ڵ#3'��o�k%,���dS�����<�t@<L��S�����~��gAô�q�0��B�
��{�N��P���[G+�s�������p]ةXG>��-f��qBGI&��*� i�Ww�M���
����O�װ�T��+E*��8���J�븘��5�^gMgp�:�[2��V7Q��*�s]gv>O4�_��}���>~~^~��7�7���a/%w?�+�����u�"�o�;��1�7�&��|�*7�ʨ+�Y^R�QJ�v�o!9�O��By���JF_A���	�#���8���n��*%�H���׽݌��pڷ��r=R:1�����!5Y�A�U�����x'hkծ���ձf�ս[ƽ�C���X�as<��Ū֠�LK$�v��)��*�eg�{б�	[B���a`r�yXj%_X��y	K���tu���r��8��Iߊ>��\��0��"�$�57�$vEê���ڡ)�~�1�vN��*XM��{%�D�L4�q��vS�ޞ����b���%E�1/e��ϻ�Q��t�[�wU�˙[�$�:�-~ܕsR��9/�/}���O���Ac�Ҩu�f�����ű���Y�x#5�Ԟ���l�d&�tך��^��Ke�B�!s��t����3���g�/�6�w٧y����S�������y�:nT&D몗�	m�<㬶��:@��Gr$)��>ِ���o��*��-���JO�+sM\�<��Q�*�X=X�K�eì;Qp��y�NŢ��J��}q }���{ʥ�CŴ�'f]�,��.�.g�����{�/.qf��dp\����VJܾ��·/zq>�������???�����W��7TW3g<^��w!W;H05~�G�8���ʃG�*i��RZ޺'�mó��FK��7F�9՜�~�����W�4�Yk����5�t���)���/~u{��{
bnˎ����tQ��_��Q"i3�[i�^�� L<3���с@���u)c����}�z�z^��k$6<vY���_A0�ZA+��$�/]�h �Ȑ��[P�[���9��Gsc3d5�HdcH��^�鬺���ýzFfu�vI/E@A� aض5'�/1���@��=�ln�(�fHl	A텽Ų/����(%�^�,UB<�o+�����9��w���z���`[9y[�灁ޟh��Do�u텈�>n6'@9	>4IU�H�3�:��o�o_�L	m�r5��v?����s[��
�x.��<��5樦�Bo"�+�f�ܮg��^CM>��s2�
W*�
c����{�.}Ol���H�U؏�D���/7����ӺOq���z���Nζ�k�"�ħ7��z�3�[���ݾ�oa�Riط#/�M��9R�ւ:���o�,Y�OMIں;e�ͯ۶�Ǿ+=�!��&��6^�)^�.�5�&���"$8���� ��)�����o\�>�T�8U1S(Z�ͮI�|M�{p[�&u��fX��Z:�nJ�&u�?����������y� �c�)ݜ1M����@���EGx����;��Zg��b��^QiB����'7�� �d���  �`gd_�`�"�C)��)�}�S��Ⱥ�7@La��v�B���c8�ބo&I>����IɥE��1�z?\�ɻ��ҘN��O<�\o'�ҥ5��ݽ��WN��zݞ��*�	�>B��oHo��+͏�����?A�E�YK���dNb�]ܺ\U�`�t����H߼��|�@V A�8u�������P�Ъ��vliqʼ��r�n�yœҋ�F	{k��z�m�ߧ�u(}w�x7��"�����Mf�8gmR�˻3e!RX�/R��_��}�`V�&�n���E��E��[�nr�|�y��;��D&���'�vk��E�{��b�0���L�O{[M1�>Y����ݼ���h2������Y"���'�a�C��e��~`��pn��_;9�;�5�U���B��hd,�H��E��^)�8f �y����b�'�����| ����O��e�ۣc՚+$ə����!�Q'kMf#�;'��\�E^JK�Os�u&����[x��fʮ��=:W���u���9�K����9@��"1�+��@��;w�^��з3�;�m��^:oͳóz�a ������:t�j�@����ϛ޺�o���{�LD��}�,�����k���_k�n��{o��I�7!
�#^k}�M���,����>����͙��8���Sj�e_oj�����;�j���޺�2u�׳gO�b�׶ �xB4,{�٩�����]n)����;�Z�بd�u-VzBeV�
Or�P<�o�"�ᢏ4:M��?������;y �&�_�q-oހ��g�7_8Sͯ�$�/	���MP��k��lûKA�]JsstLQ*%٫ڴ�B�K�o�.򔇼�4=���ۿy����ƼHť:!C�Gb�`�;}~:��ͰO��{����q ��	�3��6�B��.񩐱��R��Q$���̥��9��*�2�ؖ5�Aۙ���e�����  ���Bm�0lŷM����Y�אy���mq=�z\�����ƗJ��L!��솁���c7�
�fdE�	�����FXD��Lki��^lJd�.VF����;��@�^��n@z���V�^kX1K�	�rw}�Ϯ~��-����~��l4&D����0�;��{�%������$ �bÙ�E���I�خ�n£[�NW1���{Od�n�q��}�7���%��o��v�Z�:��UKr�R]�U1��$.�Ւ]�
��6��GBn`Ä�ěZ�CV����;'�vi�AK��.��GZ۽��Ѽ�ٛ�������ϟ�������a�lI8U����8hC�D���]3�6�Ek��#9��&}:��i�CSf��;��z���W�#w=�oP%A�
��_��RӞLZ?�D	���-��1u3WǱ��9��Y>QQ���m�C�C�xw��``p��2K*czVe��%57ۻ/��Y�{U�3`NHptq4�[E?�۞��~�lK<3�%��-;�4 �z�d�깹gwp���K�=ُ0љ*�W�������`o��6���*8h��R�~�_�M�����,����nc�^E=4{
T*�eEM�MA#��l�{�Z���Mc���#1Ov�h����F=B�C�-�Xs� EǦGDz�#~���"S]���A�\���"��(�w/�7Җ��c�iT��N*��D����� �"L@<�@Oju�ϧ��������-*��@���[��͹������f��i$>dМfzb�Ed\/0wxz,�o-}��F�0�N��s��R)��&�����*]gG��m"'�P� ����nh�@~��뷧3�h=X�2�8�/�n�x�C�Bm��6ݫޜԜK��_+�@�ed�<W�f1��nֽ���so�'�q[L��U��TKx±��r���b�hq���l��|��9Ύ�|.�w>��t���A�`�ힲFj�� <xe���&>�)�M�Z������5�y*,9�{/��獋`�4#b�L�;�j}�E��'"e	�K3�	�V�v�~e.K�} ��Y�F��w�D*�㚢"g�4�v(4[���>�C�;;-{�^�n��U�+�Nw�&yt�[��];�J��#��[��	xw�~gaw�A�K�:b�L���}�7��q�\�c�Rp�c.�u�b��̥x�0�~�ɨ��,�^�7>��V3ɤ&"
�ZE�o+���*��`��|�R)d��Y-�������ƹ�j�����]*�O��K|��!�dl0m=�s;c"���Z�U9qP�98�ӵ?�}� �ʅ��-��IC�jMv���j/a�F�3ƈ�v�S�j�:Չ[��dp��Z~�05��$6<vY���_A0�ZA0� u��<�3�ՌcpdC-���H��ig�ˠ��h�Z=���9����CvIzW� ��˵�HT�'��FP3�e��\���6�s^(�������i�t�= �MI���/c���nc�
._k|�pv7�f����g�`�T���|��b�����u����y�p��t
ó��bO!�뻟=�-0����O�&C ���漊�X{�!�]3`݅�:����#i�8�k�D;�H����÷ �9��������������yx�����`�kV�Y�Դ7�ɐ�/f۫�[:y�^��
 �����<��0�E�F�sl��v�{%𥽻��ˋ�"����E4�H�3ю�.b�θf���sb���ʾe	�緕��k꾭#�:~�ր�m�v�c^�hRo\�,-�]�Y���y�=��g����m*ƪa��i[���Z�Z���[C�%�9�No�=~U$�,C��WdcB]�d�0�s{����Q��>��.�e��|���Х7/1����m�=�#�;b�B�/v��ns]�����t����H9Q�#��=����#7�%�]v�ʞNK�"�o,Y��ҭY8��s�!����y�����^<�M ����s��lȞ��M�Y�ܘoW9w��������<��r�I��AcCR�a)��F�>;0��M��o=z^K���N��7bmت�ջ����;���?��+:q�_T�7>xY��%�`�,;ZF��S��^�5W���푫���dWP�N(ҹ�rs�l|�=6�j�=���;b6� �X��)���S`͉hh��mY
�O,��o{���	��:ַy��P�b��S���T�v?����A�rWj�t7E�ˇk4l�d�X�T�{���rR�6m���.�zrwz�����'���������y����Ek��X3	׹��������K�2�Z�Y0
��8�(ŉ	n�����P+���1�=��_~Q�\���/R���X�LW����n�09���4ft�֦�yJ���u��R�q?���
��&��X��|���e�����^��n�2�R�+���S���)��^��O#^]�N(h|.�	텈��F��0�{h��Klc
rr�����۝�e�y��G�5^:#Z��`	_~�G�L���^���bv+���n�����͜�ffm��+�	ye}����U�!@�h��ۦ���yזx��<���sB	��9�w3o��۩q"�S@�R-��81�f�O�����5���J�w�Ws�}��o�$̼��6z�˦�KFX�z7xJl��!2�hФ�(�
���~����gGTꝭ厢^'�v����K�k��HF�*󆮟)�m��bS��RX&ƃ"��7�q|���0 ���{�abC�c�On�[P.��6�@I�т�׻�t��hŉ�xm�[Ͻ|���7�� �I�1e�]D�p���ce�y�x2�
i�hkc��L=/�U3x٭�9n����1
���E6�+]_]�u��۽�e��n<��:�xL�Xf���`����_ލM6fI����Ʊ��\�λ�lef��ݢ�d���r�e�u�`��a�F�{�W4T����ͣ���?���80�Nl���d]���%�f9���!�\�f�C�4 ���&�i)��9O�"^f������
mA)�52]�Y���zo&�^J�C�&���Z=�O<!�=7B��i�Ze�X8`赲��}���b`��|���g�l�/K#X� ���ٿ45�s�΃@��7��'���d!�H`c�����XD�Ri�,�ry��+]'%ꜫ��YdN�l뺔N�e!J��03��n/p�ٛ-�WE1}Sm�|O�r9�`,�W;϶���~�-/}�N3:��v{X%h��_���<����ĠL��w���?xQT�r��.�>(HJ�r�Ey��|�(w?W�hvx��<��Ġ�Qx!�9�׷\W4�Um��kn۶���;^�َK���iض�^�T?VD��!�k�4k���=�}�L2��X�/V��d��}}Bs�S	*�!CL�{_�)��O��V�t(g@�--<qz��ϔ�щ*�C.*m�j	����f�Y�^��<L�;��ܲ��[r�Qk^���f�ʇ�b\�ˇiie�}{�c9B�R�B�i���B�W!�u���2�*W�)(�3�g�����u�h�r�������r�/�+�g�8�<k@��U�%+u�1�8���HK�˕=۝VΩ�+��[���cv��%�o��cY�gr���Ӭ�5�	6F �Bq19�&sRv:*�#��ҹ(X@�A���{7{KU�c��;�4�<�l�r^%�+�ms;���U��<ү	&=6l��	HU3�=��j�fi�=n ����0-�sL#0�q�;Co��צU�����x`���L��C�Ag)bv���R���f�Z�sgekۍ�$H+��[�s�B���w�Y�l�C+en!@Ө��bD<iy���&;�F�bV����kJb�Z�N�ڸM��K���ڸs7ZT��oj-&e��4��vo֦�=7��L�؄c;�
���ж�X�/�N�8��ye��к�V�{#9�h�kn�ǼRu���].r��6�૎u���9n�ѓ��-�Ԛj�Fwc��k��
������ӭ۩Ʒ �[szRZ�ur�Sw�;�&�Mb+3.�:ް\p�ZK��oub;�}�.p�sPHA�1﹡
��k�kUu�@�J�e,R���2�i\�t�q5��)����1a�U4ɀ��: �L��1�?u�q*T�Vz��[}$/V�)k?#_�x!��k	6�̾�u'}pW��A�:�	�"أ��Fo�����˦��t��C���4�hS�����[y{2�n@r����W8zƯ�3�Շ�m�ٙTJr٥���To6k��)��P�4̘��jYq�U�"9��̚����E�K�o	�����"����v��kSp��L��rv	{8��ë�ßL��M�;8�-��^��/7�rKъ���)��.e�I|�쮶6�L�qrϟ��u�~�Y��z���xᅕ��ޭ�9�g4�r瓨f}���YE���707�"*;��кl�V���pZ�55�TR�	K�F=Q�%a�����tm
0!}]O\s�S���eݮA[�5զU�`<����k)��}�n=�²�7��94&gݩ���7a��*�v�۪][Ǵ:���(m�P��jI�F����Jѷ����qھN_�qf���D�굖(E�tTZj��ꩺ�}�D+e����
g{x5�R�6A�w���=���Ֆw-���n��G*#�V�%m2�J0���I#��J����5����r�����ː��pf����3�^T�N�i��/��:����f�Y�������$U��$���ٯ���B�m�#��́9bX8�I�y�gwv�f�Lm���3)�ISq���IŌO��:�/<��^��G㦉><��9]II3	 �I�mx����kZ�kZ�ֵ�����ӷ�O���}_�,VE޻�n�/���B���<�%HX��A��o��~�����w�kZֽ5�k���k�nݾ�>��o�b�̓�������+%OZ�15���7��I�4r� Ɗ����.��(�1cF���(�$� ���h�a)��_=��ۙ��ܲl�h�I����I3I��c"�I�k��c$��o���{�l�߆�W	"�5��"�̢4h�+��[�Q�����1 m��
0hۺ�Ȉ&i�˝+�U�ss$�"2 H��yw՗�k���漝�l� L���/�HBo���;NZ9G�l�����dݙPң6��gE�w�����s~c��㎣�N�E��ʻ3ɸ��苙�wx�jr���ߞR)�=aŴXr]����p^����Q����ɪm�6I�7l)�[K��j�z;���}�u^*��T-���a��.��y (�p�[��Z�f�&fj�7�a��*%�=�f�X��U��\�ΞE=�ă�Jq�&)�ۭLonά��{\㸎ҋ�V3�$�=Į�,�"��%I���ff�>�`�d:�x�s�Q�bNu��u4K�3<�9n*�0�1��;�RN�=	�I2Xk �gx��>ǟ��Lz�m伈�+WuwO���c�]��~.�|�a��o��\QzL�~�-�x�/#��[lmrrҳ�V_^#����yz�C�h�����q"k�<6�U
��\�G$&2�ǹ��n�Q]���g�xwƶr?b���(�ǿ6��1ǻ\o�N���6*]�յ�Y�;;"��{|��@џj���?UA���؈(~H~����/~��oeds�cl%2/n���n{ԇ��UK�,+�~�zo��u����h}Ch�� W
~\u?�Y��o��n	K�2"�����+x\����V��LƎ�	8|�{E'�+/,X֨������sC\uW��OI��9#�A]���a�N����5-^��#�­�V\Sqo	�t�wWs'h�9d��J >���u{����}Gǎ8�0 ���G35��](���%۟&�	��j���6���|H��D�4��n�.Z���k�:]=$��]��n�3�p����չ�05�����fFwD��L3o��3�q�D�W_6����w����N"S_CU���$��X�o����Zӝ����P���b�
��A�na�̇+o6���ݩ�S�Y��o�!��(|�·g���^��)�b�� ���w���,4�w�7����ͨ���L��{,�����[�RO0�/�HݨE�;`��Ȫ=U)?>@��Zv���r�^���ư3O��z��W䮱��1��@���:��
ϬD�s�㫥��f�m���:I��sksk� ���4�D�%Qk�[X=��^ꋇ��m�-����Ki�z��q���#hK�;��`�V�nj}�^r_���kL�P�+��8�q�bÜ�E�¬�Ĳ3ڭ�syH^�i���c}2��bo��Х2�n(7M����$9�b"��+������?U�(Y�L��a�����.h~��~��ܩ����!�oS�cs�Q,"hH�����F]����\h1�V�YzM��#���u����$�Ҷ5�MC.�زK�h���|�!Zɰ�ۼp��Jm�7�1���U�`oq�]�1����x�6s'sh�dmeh��Y!���'���ӂc�:� 9������]��̖r���}���0Z���-m�gv�(p�!�K�K�4{gls[)���07��PΕʓ�TU�K�!e���P���b<��k��Ŵ�w��v{��
Xe'�Y>�E�%��b޾J]��xw7��䎿�=c㿓���T���W��ͽ;q����=�R�Œ��>Y���7��|E��7�Ҭ@���ê����ߟ%��Q�·���qP��`c)�"�{�x��|�I�^�BOmaTs9�s��#�+��::��g�s}�k�y� ����y����]ٙ]��`�}z�-�6丌 C����}'c�;\+���-��u �fp����L!�2߬L3���u��
�^�[�7LR"�r����ؙ��{T���gO#^]�4,�W�B�zQ"Az8����TT����9�+gZdv�{�x�v:�Y�����.!�p��'��=�2W<���<�^��F4���yj���W!
�#^in��H�ίE4`r���N{a#]ݚ{�����۩�@�p)�g)�{гtd�͋a��*�;��?+�S��}���8D��ǰ�b?Ѝm���N�ۢݛZ�a��Ҋra�N]n�d�k��8w����e�����c?����R�K��,7ÞV�i����6ǁ�Ӯ��q"�N��L���I�F�jv�#����I�֯W�o�>wu��3��@Ɓ�F��q�=�U�9�Y�x7�0)6b29�z�hfcb��[#(�s�����/��7Ϫ~x����B��j�G8���ʟ���:ͤAb^�B鋮�t�0m���̥��Y	�5>k�'&��\g�*=3r�(8�L�����A'���x꽓�dF�el�4���������Cz]����ßb�י��f�C�D��)h>Y=������3mw{`��1I�F�?�!�L�t� ��4��ký4y�[َʤgH����6C�m��<��I�O�)�zŧ洠���T?5�Zl�e����c���]=�wP�׵ ��H2�<�cT<���a�7�л�2��+��%C9�dg�}���E���eN�ˠ<,fk���<.>�TĶ���P�U�XW�Ru�%����s(3�{0���#���� ���dl��AC����x~�(:�H��o5�Lj5Pي�5�^E��8���Vr%�.�N�r�inD��gn���h�B.��uC'����BXė��"{�%owк�V�ZJ����9b�F�v<o�hz�l��7G��{�yf�ŏh&Lܢ{�^]�/�,��wjgM����w�s��]��]IJ�a����jӆ�ZWiT��V�[��3y�Y¸_5�ɡ�������?��0s/����3��8�q^g;��ܯ����Y�C��#3�4�~a���mq����M����*�m����C$6Ge[m�%�� �;O�Z"��ڧK�VT��!����'s���A�g�:n��/x�o'�.�hEn�a>�R�3������)@'r���Sd�2�xd�Y��c�J�ӛ��sȬ�[:JF_A��`�.N��j�V+�.��_s�{ض�2��GH�x��FI�z.=3�l	��j"Tx��B+�4�;�z�Xjd8���1l7ǣ1�����3X(>��� y #o�H�_��+qn���X�9���1,��bY)PoUT���=������@���^�v��m/Lhdd�;{�W��]��N�r�;�����eI*Mf�dv;k�C��hk�����Q���9���A��_��� �p?���K���R��s>���jE4��(���(�s�F��΂�a�BuL�75�K��2.K�} ��o5Uq�l%��M0�.�Y�B"S��"�m�ܾ����!�anuض�Z0���@�CE{#9�ͽ܆o#;7��kH�>95=�y���[%�U����yR����c��(2oI3WNg�X���,5��wc|�/��>�������{��x	9� �K{z��A�p��Ϙ\��m��(%��O�;��P�]��\��S�^�bh��z����jg�@j�@pq�`/�1흂>��v��+EH�{�0%���Pl\m����]��9���=�2�ɂΎOI�߽�H��Q!C}ഏ��#��˞�7��ȧ�U�������Eؒ�X�O�S��~!��w��d_^�H�1�['�ɗ+r�ogo����v�:���ϓjFH��8��i� v׉�b�N[�`�%d�-;fs��A���H�k�.�������Zz	��&u����n[�on~��~�@ۑ������^���>����|?c�1�I��ӛqw]B7`���mM�ۚkmm�=]�F�@Q�v+��e��x] ����E|�C��\���2r�>�y�OKR������⠆梮PjH�i��g�����~4���,�U��n����ɵ�[^Ge��ݭ���7�M�{v	|kЃH�2�$k�ק��d�Üp�a����j�/1��7FԴ�uk�q9uP���Z�/����k���p�%ӂf��Y�"ܦy�5�C2����aۻ��*u0ȱ���S=k؍��P���:�
#�m ��vv0v��Ebƶ9ڎ
ڃ��jM�f�6^����B��O��Ӄ�,����v�d������yrv=�6�i�˳"Q+vZ�mu:¤	����_��3�_�^�ZE�4y�n���	�zѡJ�QaL_�so����ˢ*�.V%���5�|��l.g@�M��2.����n8@���ͮ��b��B��]�!���n;νf�S�سL%=4g<�E����ޒ�y�	rm��l��"I4��``&+In1��K1Ge��-�CK�Z�W���M�L����tQ���#�����a�4w����2�zV�훳?M&���/�]υ嬿&�1e��n��\��]��Pqm	�2�tX�MC�rdb]�=�����l��b$��E�Vv���-G.Qt��:�;		��F�>;0�6��X�>	�1�n�=kv<4s➑�}<�]��¼�����+�a>/m�<Ӽ�4�Y��r0���Q��&L 8Qʹ&��z̊U�<\P'��a(%�Ts	={�fy�g��C8UXp�`n�!fp��4��F'�!ٖH��	�R�ŧ�5n@&�: �W+fE�oo!̽Y���@k��&|<�пVE��}��[�\V�,#:u�*H�ζ�|�W\y�ZJ�q?�Ow���5��/jޡ���h�X=t����^�����s�J�L��-��P������˭�v�c���Rc��qau�f;�%mι��Yے>σ�����6ܚ�đ�Ԛ:�oS�~�vy&a>&ޜ~�iӎ��H�F��^�:x�~�9oZ�ۏ�����)��l�����4>�yOl^��=���wsG�Rμ;�������>��Pb�ʇ������?�ӅC}�긬�@�B'�E�K�E�93+mLgtvwocx�:��MmL���U<���T7�25^`�V��X�J�+)ȟ����u2�l�r{;ǚ|� �g8�̚Ob\A��MT��g�~�W����&����HM��O�����C�QL�x"E��t_:�Qz��[���%5��	�F�'�~T�foT͸RUl�����f=ϝ��S�;��ˉkwڟ�Z�Z��D��cL_�GZ������a���P�����Ο=��[@N��m��OCwj
2�&C�q���3������W�{M��Y�ؖE�tS*IR`������x\�&�1��^�q��|���!��6d���.�_��E��K}c�z��ŀ�:�fgp����Uuě�E���!6W��H�y�"U_Rw��=.J�[�7%�.��A8�m6�\���mX����_fmI��٥Eb,�b�hk-ލջνQ��;ᧅl<�����Xѩ́NEn1\!��+��]w��ZpJ(����4oGs��8G5�լ�Yb��i�o��Ƙ��ڂ�	��Ι�����>_/�0�fa�3l���؆�"Ho�`��΃�\<'5�a�7�л�*����e)�r+�#�+n�*�%�wvb�R���a?��?{��������ϫ�~��]�qܡk������fZF�e��8�N��ژ�6�@ç�0l� �<��++�$��OΏ�5k>��|�oO��vu��^ÉI��O:OͫnG4�v�p͚:��ϡ���m�0�Ŋ�oiNo5��J���@����π��pCo�{�h��?5�v�wy!���Rov�L^5�L�'�;��p�nV���od��l��%ɿ4��Ӵ���H؊�Lt3n�d.z"m��ރ,����C����\�s]{[�z�rO�I�L
��CTl� TԻteH��Z�5���a��ױ�A�,Bii�
7�1��͉�Azij�ʅ_A�Y틭�~����,�s���$i�?{Y�9h�
�c�4�����EǦ|�ӌ	��kgDl�t:ūN�ɮЋ_!���A#8Fc�M<�n��~�,AVD���x��w��t��O�����.������Ef���G.�f웘���D�Ok R��]�]u�㰊���I(�����|]ǻtʢ�|����[m�1�9|���y�_
��*�NfW�s7��<���5���]��sz�䏩��8�QB7__,U_k��{dֵ>��.(bY��xղ��O�{gO"���A<;�(�"��ά]��t��&;�9�½}+���$��%9���g�$�5��@2$��w��,v�k���"��>�)D���	����>�=���(a��������<��c���T��LU���V��0��+���������z)T���y��/3��"mLpm�^�j�i�ȹ/I�Nhs3��Q�{�9���my׬���=4�{�?O�-�x��|9ó��;�U����ؓ��6���E�:.�/��9HM���z;�,g��������6��=�u�~7R'�p��a�&g��'����̫����%�Pv� ���.�N(�<^�+^�+��N��hA�����-C���c�&��xmk��:�'�~�/O�Z~��~�L�נ���4��xz��W8A�=z��z7�.��"Ԍ��I�I~�a� n׉�i/����;
�mv��2�ml�;��?y��,�2��#���b`J���}fFwD�����`�&N�z1V&�2��6�G,݇9Ը��[D7o2���ged����y�g��.�����F]'Y�\��kEEЌ/`Ե��\�2+64�X��t������l�'�5�����ή"[��j�w�e�
�I>�`+�Y|F#��h\��2�U�nc��S�˦����=���`U���Yr��m��"���+�>ܷ�d��Hp���["E����v�'/9v�[���l2��_5Z2�sB,����n�W!˩�c`�������g���UY��z�W�wg�:΃<.�~���7���Z�wzp9&�ZҬ,�R˗��\�Y!<gA��n���7EX(E�N�[�.�+�V͗:5Pۗy�Fs*bN���[�9W��|�	��l#4v,�j���\J��]���R��/�[���/gV��)JT^>K�1����G�0�	>{��-��$F:a����:��ѧc���0)m�ۼ����h�/,�1���N��J��S��Ů#�n����d
KdY��[�՝�_H�v1GP�Ul����y��5ЕDD�mh��7x�;f�SĹj#d��c�	-L+ ��I��]�]��z���jk�9�V�nK�:7���+v�u>��4a���6F�9�3o����1qu]�Z�kt�'`�Uv�Gm�*��yܹ#]%���#v�':>+�.��-�T!U�7Si�N\ ��0D��mEU*?Ed����ܯ�Qo��5p+��Fbƭ]�5e�����:�{�s#�SV8��+�(X�8�W_s�bV	���U��k�%�h.�� B�`X��r{���wr�an���=��Dm	�ob/v����2�ٺFN�����%c	��+ee�)�K�#7B�Зv��"� �ޏT��8�QN@��,��IfM�D֌k#��en�؋�L��sbT/[� toC��:�\ی�3om+���v�'%v��Ew�����ӫdޅ��ح�G�y�8��2O���a 0�ޖ�'�9�6��Y�Gf�i��A��O��Y,���L��#��3Tp�3)��\(awm���rc�i
���qq�����u4���5�n��l�Ȁ̙���!1���V�[Y�#��:�)��K���C8���%�ĉ�9.�o=u{�cg���+&7�K�_L���k ��ȱl������Ы��@m���2��Q��%��^�F�'����B��7	�o�x��(���R���0�U��!�[�6�ҽ�l�}�F����wT�a�j��w	���{���j�<�f�,���v�6�@��-��n:jrx���;&:gKEL���}8�f���ۛ���� �x%��@Y�6.�<�Gm<�Nl�o[�	���$�2!%��1���W� j�������ƵƵ�k^�ֵ�Zֵ۷nߧ��<� r!�ar��ذ3��!�۷�_\kZֵ�mk]5�k]�v����<8I�7n��W�0W���]3,#i ��
�V�`�SO�r6#!D>7ǢlO���L����"K��9��pDP)HRW��x�㖀#owH3y��6����縬����|q�\�}\��A�%H�3)66!5؋&�{�M$c��/��>��K��Fũ(/����u�]$S��j�,%�D��wlh�-�|k�����ME���o��1Gw���6&Z���q��B�e�E������~M�ѤMB��"�M�Hr�+6�����sw�)|h�I
��Վ[N��=.�Z����B�z�f5���3p>����r�)̈́�"�,N2J$��b2b-�Ya0Ak��+�@]��
��iS �L�h�,�SA� N�q�d��Rd6�D&ZF�A��F�"q�����?{�����|����<I!�}�~E=(�W��GB�2�~��%ch�j��^��Żz�٥*e���^�	O߉>7A]/��?;/�a����8���~P����~[�}b&K���eL�^�n��=���e�ށ��{֍�-3�c��^���T��-#@|�d^��LCVZ=7��Wn�uv�݊��>*�K�VR�V롬a(O5�Nƻ�$��}�]IG��g��B�ޚJ�y#�z���-]z�ʐ��q=�wM��g���yN� �R����z���et�J�]�T9ۛ��c�����8�� �h�^0nFJW"�Hl�M��i"��U�_�>V���n�����j{-�fg���WbPo��t��W��By�ĶE�=\�uy����2��s����з��u�BKn{if�Js3�vx]��s�%�����&���q�R]��|�zX`�L��\49��D<&�� C�fY�M�n�a&&Eq�WgQ�
�C���)�����td?�ώ�Xh4������D�;�4�~��U~�E��'gK9���II�M*�;4��9�G�H�*ot��:O����k}���;��GQ�n�;�~�����{Ư�0).+ʕ���$۹�x�v�e{V׏:{���܀.�����}��?uN�@$d�3�qV:��[Q�Wi�˕ ���yV�����d�ѷr:Y]*:�G�����c0>o.�Dv-�(�=�k��R�Q�֭�Y'
b��)��eI����|w"7,�Ƹ�g�M!0�T � ��r�^�Ż&�8��ք���V�5�_v��a��jRh1����Y�.���� m�]b�A���F�5��&�����M��vG�$���i��q��475ƪ$.M]�ӽ����
w�|��ȑ<KA�Q�/���p��NU5�F<H�Y}�s���l���R���D��Ǒ�U�8ykײ-s�ėx��\Wh�7�_��b8r��m�}g��!�&^�7W��hِN�l_>Ek5�gb��<�T����S5Ce�
jh9�����n���R=�4_i��w�Y񊧜ړ9�ϩϢG����ԫݕ�M�rU�:�B
�Ajgm����dN���?��'�<���>�mA[�]|���u]�����ɹf���uɊ�91��S���y�5�_~���
c��M̺��G�NR�Q-g�)�	�4�y�,l����{ǲ��J�fː���u�yw�ﳒk��}�>88�jF�\nv"v2U���i�~��=�IU>�첹�q�<���I(|n�Q�X=�)��V^h���A�iRJJ�F�ɒIT�}!�z��k85T�9��71�q�ƻ�s�+ֱD��W@�M n�$���t�`��yx�M�/A:ۚg*bQ����CFi�+����?��mY�;��$@2�?E�`�)�zм�C����xwf.�_1A��09�`t��p^�T	�#4�/�p��;�o ��	�����sh�g�����0ހ�o;ױC���:��-�8���役}ݤ<jL�L�J�����9�����@�׷ii�|�6��\.��{���7��x�;4:CnsP����yG_�4��ý���\��e5����3�)�}�X�lÙ�[.���ݥ���RB�<�B��<h����������"���/��/��B�B�:W+�(Wr�ZU��3[ww���1�ʮu�1y˾����%t;��-i���p��Ëb�͓ͩ�v���ѳc����	��idZ�?0Ļ�P�יE�/	f�KN����o�s�ߞsξ�^�~�ӧD$o�DU.K���߫�C���@**�ж��}�n��T|Pr�i�������';�Z*{]!���	ک��+=p�*��zB���\������?T�&�݌�����8�R���Ɯ�R.�F�=�ɟ�ǝ�+���(�B`�	`n�f�k�rB��]�|CO�A�OZ�̟�U���G�A�b�m�Y*w2�뜉�9��m�s�Ƕ.3e��TH�y#*�;UcU���0��e�0�ng�ǅ��%�Lbb�ղ�#@7_���Ue$�7T<[U9ɧ|�]���po=L@*���@����;�%~n\i���_GC�V��\G~q��߹��i.����>���f���s�M��Rݶ���m�E~�t����g�@�2.eU���Cy����h�ٗ�vAwT�n�N��٭zR]��X�]�-�=!l@`�= W��/��3C�`�$r�+�>���L��q���n���Nj��Ë�G�iˢkӨf��y�	LG��ḰV·%�c���u��(���ɠl	Bg%�s�+l_s�z��m^͒?���ܝ�Z��9Ө�3u=�*���y//!����"\°}��e��"r�T�\�6��gZ�A3�w0�=�*r�80Vѳ���k;v�"n�,�z�|;~�<T�}�iRR���g�7�Ϊ�X��=Dc�!��gF�k��^��g�cV�1ˬ��7aO7��k'�A��"6��U9o�U���Xx�}��KK���3��-�}�@��v�'��v��ٕ�]�YOz�z�k|n�(3�x�[�u[B9*�邐���v��EGm���U��v�P��|8%I��O0�TH(��^�ɢɥ�3|ь�%5
���ήr8��/�4�N�[ix�>N��bZ�|]�n��9>��hm=_v��AT�\&�n�u��`�n�哏���������\ې�O�eߠ�^Yq��R�~��~��h�wVw��gE��I���WOR����d_�!A"2�@ Q3W����~5h`Ƣ��T���ꖶ��w��]4�M<	>^ȟHڎ�s�J=�>"�ny�� �.F�YM�9v>��m���N�=�w�z��cE�k�e�=����ݽ� ���޻�����.�`��;o�� q��|��{{kK���hae�|�p,F뜮�x�U1v����*��E�ZW:R9�i�5��Ss�g�s����tO��G��.8�j��Wo
K�_�o��-N幑ِ$[���x~��q���wwYig���@�;u�E���.5�i�Bm��Pk�3��,��˨A���g�lk%���Z�K���fuEu���^=+���)K����/K�bE�z�n�{ݝ"����c �E3s�?]w ��D��h%݄�|��+�'��{�[�;��WC�z�8���U��ʼ���Zy�|U�p�^>9|vh
oNi�X��8C��C]"8�SS��Oj��=��[w�M�eهvo{;-��7{�������7�Y�r7�8�D�W�sGnk�
�f�9ݘ}� d���ɠ�47���E�l��kz����+�c^�>9֫���U�Gl��8'�M�����\1?�;^���ҙ��HL_��:��q��'�)�~���_�x�������btV���Yv�F�Z�rvb��/�n�l�&��S|�V���5�$�h�@7#�7�4E��x=�%Gwbo-Mw(u=(��j�1e74�z�gZy��]�E�v����E�ޏ`u���]�]-fUeoI����w�yy <� ���M)Wk��x���]�S����Y�'}ʳ�S�M>����-�cy����x�9vajP*�ɨ~����н�f�^i0P�X����~RG�w��mUv�7ݾ������Ø1�z�g�Tϙ��^���<�o�[��*�in�T��^2t�n\�do[T<btj��;w]o`wv`���i����x
�T!%@P}��ebi�uהy�����o��ok��@��	�>�^&U�]��I%W�����N缪CQ�	�L�����d��Ɍ�:`W[c�8z��t����Z7k�z����	�;	����1��s�Ц�4u��ԵXH�=<'�2m��[v�ވ��RSj����~�?k/��$�2��\E��%���8�I���=���5��w����f�Db��$cժ�A�D��h�=�Ó]��3F���0�"֪��S�|�i�۾pk\�9ZK{0�9w�"-��<Y�Oe��R��Q�g2=��ӹ:����ad*��qdD�H�k�F��~�� HF���t}�c�u҈�2E���w���o'R�l�OO�8�}���o׿>js���k��iU�&������[;�#��N1r�����é/'���B~�١Ŭ/s��:��C�6�sh��bM(�[OG�f���@�me.����y�y*JjGl���르;���|��׫C��J��°�K'<�7D�ܿ$��t�<sM������ώO��ż��N��!��/�>��E\�oX��y��(T+�&x��]}�x'q���}�N�d��,tB	�U#U�!������׌[�}���bWU� ���e-	l�U�L�h�a��k9��\:x�?/C9��O�t�t ����'��˚�A�, �gy�U�om9�s]%�t�	�z����f����L#�HʯB3 �܍V�u�7/j�j��wfƲ�^�h	�=6� V����H%R��Uq5�.�F\0��r�ɓ�Ҿ�F��_�Λ-ڹ�:�x������K�7*u�́}� �v���#���E�lٓ�!׆�����Go�ɷ6+��q����v昻p͗W��y�l�̗���ә�����<�7��8��?QBF^����˼ߛ�f��I�6�=H��ܬ���yYP��{~�������^�V��n��S䱭qz���`�1��Z�T^���m�����4quy2ُh+b�p� ��^~&�
�c����%���:i���$���|��O����K�`ˤ#��+�r��Ʌ�����ݭ��}��#o�:�3�wj��\�k��|�yۄd�ȥ:���̻{Ol���=���i��;H|�Ty)
�zhҏU�6�����Xȷ{�T,�Oq:c�2DV@p��6�½�;@s�u��>��z���d�l�&"��k�h'��c5�#�ȣu�o6A$��n���m������M���e�Ag��W���`ǣI�YZN4FGELm�9ё���'�+��^ݷ�����:���<�'���7��u����֞�V{��ADi��mP��s@�H�ހ��v:��ow >^�s��0��[�׺Ἴ���K#Y���&(3��u�Jz��)�T{�R/Y�wW���%�>č>B�$�����`�`A�U��V��m&�C�쾜���Z{}�.$��9N;�Q��ز@-::'#��U��n+�����z<����7���J�{(��믄R��zҶ�x"�K��E�~̅����n�/Xu>�}�'��`t>��b2�z��o%u�����1�VRZݮd0���w�.�7�(] R���t�=����,B���cH����A����=�I�su�}�w��me�ĺL�.�����h��Œ�y��o0o�a����ʩ�7ۖ�,(]�������]�~k�W��%�<�\�x�����m>�wY�0�n�7�M���Ԭ7MyRD�ut��}����:\�4�vz3nѶ��í�5�%E�ι&���ח
����!t���7q�,��U�Fu�5_b�
��_ue���U��M�5仧��u>P���c�F_:X��ݮ��;�d��/ҕA��3��r���h*��Y�dT������3,��:}������,��{VO��NUv��wL�9\�O@Ƅr�YИ ����ɝ>�=>�������R��p�=�m��[��B��#���"��2r�`L]�����V��J��t�p�9גo!���jh8�X��%�$/�ݤ�ٕ�G0�
���ص���&���'�s]�����`[���؉
o�rVoX;�*�i�w�a�G6E�sC83�RK�f�A��:A2Jԭ���8�nG�J ���<Bv���b��ҼR�״�	�b�N�"�T-Bc��
��d�ϥ��Z2,˫�E�N�{��ڊ:�(�$�l�O����bL�����t�8�Tר��32l�>���������s��17oa�f�!E����ԡ��:Lr=KM5���]��E��s�²\1��1�Z�ݺ}��KA�[�bl%��ԙ����۸Z=�R���Mܔc���Jb��8Kz3����v\�^
��Ʌ�*+���΀VQ��&�ժ��7���dJ��k!��S�q�^��bǻ�'���T�=�;4�V7�\
KX�2�Y\rPoQ�4s�\ͣ'�\����	B�ͣ]äQ�v�[�&��hЮ�3^�X�]#:�TV�aLa�ٽ;_cR�>��z��&N��q�q��.� ��t\�&)�&9rP�d��QY��]孇��O��2��
��n����{0ѱ+Jdį��$ŞU�V��g���H����;�3��7t�E�����O ������3�h�^/�̘�R�r��mܶS�EM�+��9�e���n�NwuI[���5i"�^���9��t��|.�i�7��S�4Ѹ{�K�r��P�s%%a���uN�mAq�i��]U�.]b���xb���{L�3�=ي�jw�mo	���$O������M�;�7i�oI���㫆�r��w��R
z��'��h<x�N�S�ܝ�J��y�Ɍ�;t��R�(s�twC��8�nc)�wծ6����$Ĥ����Y�\����ƞ`ܲ��b��UW(�kw
�̓���VѧWis#u	�Z�j�je���m^`ȹiP:u�\��W��:/���t!�xQ�c���:��NNe���2���e�[�E������%���!K�Y*rS�]���7���������t�e�9���o�KJ�qخ)=dU������T�fu�*�S4��;sGK�$R���޶�R���%#ꜗf�^B�o(Ռ6�k.���"�f[::
{�tT��`��l�N�GT���gj��l��E<���X;��\�h�3I���{eYZ���֜ޝ/����ESi��sVmZ9"[�aRC��IrHk��~���|��G�կ ��9$YD�$����k��ֵ�k�Z�MkZ�nݻv��Ǐ/��"�XK0������H����$�����׏�kZֵ�|k\kZֻv�۶��rZ�m�i�s\�a#FأV-�����u��RTm~����^V-�sNE�{�|��_X{�tJ�6M��RܵsQ�ͷǆ`�\�����F���봔mym��[�o~k��b����M����+���#�sW9o�����YW��Ou����*�q22�Gy���"ȜNu���@�mrx��Z�hë�VEԛ ��m'|pݫ6��z�+;�c�bP=�ٱ����v�'��g�������������Y����g���_A�mm�a>1��g��ʮ�<�����{�5�#�<��w)��T�-����SÂh���|�z��0��y���S��7z��\WU�*A#���zt۝v�/�WS�-�\'���5�1���˛���6�e��xL�%�D�%�^^,��]J�8�Q�B�~rJ_���&fG�=b}S�뺳�u�ϹR���Eu���0Wek�3�s����w�_���~U�U�Oi��q�x{�J�6��4�v��O�z�}yj=7P�vYȧ��*ҷ�OA��<1��wv_z��Y�⑫W�J��ۺ�sb��k"ؒf�ܴ�['���p���F��i��y*��}���[��[<��n�\Z�"j��WFu�vYH��S})z���4�JD�����ӦBl��u�*���?%S���P�,e�t��F���7���v[�ɄLF{�zGK.���gPn����O;�T��B��'�N�a�������ݛ��Ѻ�P �$`*TI��³��c����0)�2�X4�/�ę����0˝�_h$�Y���h?�~�8������o{8�]���U��������E[t���m\�n� �_S�ӽ0rO�8p8��EߺM�����R�ۂ����?�M��3OF>�Ćq��?u�WG����Tp�����5w�&�v�vgv��c���mt�g�gT�7����.���ޛ���oz4�r�糋�C�Z�x����5J��f�mn����IV�|�UJ's:;{�m���Fv|�ru֬�*z��[PHm��p�ݶ�DD)�;�����2G�( =:�i1�2<���뿻��M���/V�>�ċ�6�C%ޓ;�`�g<��0�l�q)���Z�I ��[�w\{���Nwv1c=i�^���r+��O5�c��K�Wf�7Qx��7X�ZCz=X(i歕�/�얱� ��T� �^�س'�+�}�T=�%��׽�CY�\�.�;�������bH��G�kolv�p�D}H��]1o���c0���'��KOh��m�ڙ������s��-�8�*���u���0fD�*Ϸ��N�'W3�ӹ%)��Y��3�ܝ�_@�t��:�5�2{u�d��w�����u�z�/M���Q
X�F����f�k@ ϸ��#m���Y_�Y�@�XF-�AԌQ�͵�J��٫}����Pd��G�.%�н��{D���e�r����c�`
�B��q&�P��5G�;K;����"�n窋�'��d s��S�b�DV��2H�Xs)�Rگ.qU=�^��Ŵ��8����q�Oө�p�7S���[��/�%w\��fz[#�󞮨������]@�2ُm�L��d�]1!��.��e���d�^��i���z�L��r��@�k�ͱ�+���[�Ñ�n���W�9���{��0�����bGZFk�wN�i���k}�r��"d_�|�md��iB�s����m��U�^�I����h=4�m|�|囗��ս�x�G(T��`��p+%Nƭ�};C�uQ��&�ʟ�+����Nx�Q[-Қ펤��k�4���r�@=�ܗy5_��?x���Y҂�̹&��\C � 2(��C�����]>2
w�Z��0�������bieZ�k���\�!׏�8�b;8���>9�S��=��������y�=cƙRJާyj�7}����!=؍ Q� V���/ҸnLf��/��yU_��1W)tw��/�����)��}�8��*�I`���y`9�7�[��V�<�g�#�\��H���M��!�/�஋ù�"�i8͞Gq�{{������1=��yI��=�����*zs��`��;�U^&��[���xbn�hE\�O[>'k5���G����H�ټ�n�ɸ� G�x��{�D1sy���R�,��<�p�d�d�($q��V{|���F�4�|�� U��F�̇����*F@�v�l����]�b+���[�ݰ���wv�q���vN�z�g����`L%�8����B����uٛ�����Ġ��)x�J�k3ۖ�}ّ"��%r �xA7Q1��w7�{=�B�17��L�qA�T�N��ߚ��9��Wrvz7O�H�h̖��ؼ�w�������/MP�:�g^5#';6�3.�<�A��U�Nx�~!���7��F�Xާ}\��"��E���"��JB�Ƿ�[�O7ڭ��&��mj{_l1�=����?�z�i��WU�<@wmτHȯ�$V�ێ'���|RZ_t������.´S�ɋU���E	jd�F/�B�����i�H�K��:�X��,�
pb�=�b)��a���D�o��%U��Y�fY��i}�\���oO�+��g�`�f�vt��S�q�OG�Ǫ�6ea=۵}^���6iZ��z����~�h�7�>y�@p��$%�Q�1۹|[.R�:㳑z��Fwn�gƃ\���`Et�k�.�;�l⳺���_u��S��V�I�My�+Ľ���6�|6�JͶ�m�q*����%y!vή�kyc������5�Ķ��A�v�*�8hw9�f<���=��3�Fp�j1K�A��h�ok0d�
��f�ӛ-;q�wf����վt/qH1O����BP�rj�-#@�mu3�m�9yT�7�қ�hf���և�g��lZy����t�f��K���-ׄtU�Jon�/�X�?H�z�����-���
���f.4�����452���d�gX�<�0�:�b�ڣ�vF��8sK�v�wݧ6IBoc{�i>���yx|ޏG����z�n�#Up&�l����=k}��g3���B}qa\ ���
�R}������g��ƗAB�;wQ.o�q瀁��EF��U`8�[��։{�z���zF-�:gͼ�к��UO�{,�i�oR�4:����b�3w����a�6P�(钕��il�IT�|�HzS<^m����F�\7���E�:����lUś����Z4��� #���U�u<(�d0�A �y5�����〰m�6&0��bH�dt�m��w�N�q���qC?xN���H 9-��>��D��m���0Y�aܭ�f��px��?S�J^v��z|���6�I�6�|3���z�0ހ�o�"�k�4;z������"9�y`�+R$	�
�t����b9w��h��i���Y���8���@ˊ3���[_��ƶ�H=Pd6�D���i��S;��L͉�f�9�m�[�8�#x7Q5����b��q��c�y�[��	��w�+�Ff�c�h�1�ޫ�&e띹e��c����{�+
�xLZ�Y��Û�Ɲ��2�¢���3a�[����u&��ۚ�~�8������3+.��?9�=����ra��F�3׬����_w7{3�so~N~5�D�:���\{Ո�~������v���i�uwk��К����r����a�ڲ�q�E�|��mWY��T�5VA=}c�Ǝ�Jv)̌�rЮnI`��4-A�i1U���m�������>�ȩ#N���oF��L�z�6?��]�נO�`Z���d�^Q~���w���܇k��dV����y'�m�6��޺e��������p\�������݂����ۏa�� �iK�'�G�$\Ӟ���<�z����ݝGUT��G����G&Q���P��
2:��L�'���w�x���sDR�Ul�s�T������;,�4���z�k�;,C3��Ot�l@n�`�]	]�A�פ�� �3�JC��)�}W��ԗ؄�C���2���7K�l'�P';Ƽۯ�`f[9_��v,���ϻ�	��j"H��C,#�w6^v��fI�F|�ᠶ�\�>����Q˭����"Y;a�1K��ni�d췲通�n[��{Y8�p�4��8j87��Ӓogi��3�Ic,����Z�j��H�����7DdAE �}w���|����?�ݝ��B�I�g��gA���9��Q�]M���-蝜g���8�>�
�wv,b1�#ckTf���(���ڱ�g�[^u[۵��N�UFQD��&;�X;º����3�Ч[w�;�yHW��F�ˮ�ۚ^�.b��f-�]��=�-� ��������S��hs��=��nq����T��ˊ�zF���F���\�v#�Q������-�-���y�'�E��ʉ�|�W�{j�XX<w�gl���+dc�G�>�z5������~��'�b�L���WN�t�p����eL���c�+��=;��¤��q��=���Y�AUg��=	ө�2���P[�?o���������j*��"�y���^���5	�1�ͭb��	�uO��T95Tuź������y^��76d�j�.X=�'|�L��h��e���ж�9�7�
��o<�T���gr�Y�tzu-5}�vVboNR�n�2��-m�d$�$>�c�y����y�:ҊU��nW]��9�i_tX9�/w5jPA�����N�w���F��P�5��?�`#���aR��������<30l��������eW��+^����;I~{�U�^56��f ����}�wd�ol�<���D�Kw��A�hJ+��lk6����}[����$��.���9�fY�)f废̑u��1{Κ)]W|[;�{�v��q#�)y��J�6���[>k�3�~g���޼X�P]����6�8�����R�5��6�x��7�ԥi}���_v��Z��2ߢ���`qj|c܇G4.�(�5��n��{��#�!��N�Kve��53��v��d	l�1�dy�olAR#zt�M�rť_E�݅ӹ�����V�]{�,�l��b�:<��H��>�*�s����Ҝ�Ъ-0�/Lt��Q=�5N��8ω���J����l�����G47��)�\��m���=s��R3|WW�����woi8h_�ϝ]m�? ����$;RO7��7��0��ݘG��;�6��6z���Cm.7K����	wJʲ��ׯ�,�"�������/����r�훻q(7%���V@ź���^�ˆa�VQ�V7Ldю�֞��3�h��I����W��7���� ��Yը��\@͏P���h��G��K��=:m˫�uR�D�w�ִ�D7#A�x4��Jƍ�S���c��l������8-�߹S�M]�]�Gy��ÞAY�'���UEw����0��=�u�p�~�^�GʽFO����T�1嚐��%w&�b@����
./��v��Wj�8��FI�i�2�Ĺ��t)�"��.����掝�]F��l�h�ԕZ2��3�SNdU�xsm�P��ޅƄ�n�x��t����J���d6�d��O$�*�o�s'i��'��:���^�i���#����"ܦ��Eo�)+a�������QjY��;��U�^]7�3��xy��WB���|�J��W�n�%h�"��D�as��u^<ɼɳ۝�E���m���A;pY1�d_A�\�c�?HgؕL�c��eÞ�-7����Ȉ,��S*Vq�ˎ�ln�BW�q�ɠ������B��E]��t�O�J��1S��'*aV����v�F�Vx���UL��ۄ�(���Fp`���h�Y.X�|uJq�YN<��֎��[�BY��^���Ozz�k������;��E�+.V�d��L�7��s�"_l�J�=�osI$���;(���H�)WgCUmshc�ޘ���
�m��������<7h��|��,U�k>�sY�}ݚ���H��{m�%g	�z�ܹ[1�:Rvb|����dS����������U�ӎdtU�2`�]��xD��AN������*�(Ďbq��Ev�n#�Δ7-�r�1���֫a[���[��;��u�Z��3�Qf�U�2�8��#����oL�C��y�{������E�.EcT�X�FgZ�drs�%�ߓ�۸&M�ݚ��F���F h�<F)���hkuY%3��n�}�'cC�v���&����V�mf4����ܨ����7F� �C�N�Z���>��j5v'k�y3�,��NLw�� ���a�n��gj��޼��1u@/uKN���k�Z�V��:�y�� H�����X����:�4�U!U�N���K�b�J�%�h����L��Z�y=��m�UsY�]���ow��4C7H����V!+���V;XEH�Z����MI��y���L�A���â�'�ຩ��k˵ڙt����Ao7;<��캝}�ul��d��/�m�:$���t��xw�mۓ0���۪9c�+#4�k�s_&�x^J���Sꐬ���Y!�`�rfVk��J�Ֆp�y�f&���6-��m�����6�T�)�6+����-�m��]y%A���p��X�M1�w��-�V��Jhe^��w����L��e ��uk.�l/��v1���b��s*]a�;.�=Ⱥ�Ɂ��|��kԶ��㹵�q2��txY.-m�Ytc��ec��@�TPN)t3�'N�5�L��dXZ閶�����%��k�ns��7�ieξ�c{tXӝ�AӮ̒eV�sj���&VkG��z��`�E���Z�G�#1b��)Х�˚/���֚��*�(M��pL��r�T#2�f�.ۈ��Ȯsi��Q�u'k_t���Dë$&�E�:��枓�h!ܔb���ܼ�����e-	}�;�E��Y����h����2jd=ᢸ���{.����l�j�HDHr���Q$�U�Ȋ����ʒi�Y[c�C*ޜ�Q����ט�7��_8���*\L�p�9j����K�vo)$�I&��������}Z�}mr?��Uy_5+�$@��DcӧoO�}}ֵ�k_�ֵ�ݻv��x��$��
�~.����]1��ut�2&� �q�����֍kZֵ�x�5�k]�v��_G��3�25�忛��nsnk���������}��ٌ��ڹ�щݯ/�Ƽ�6�Z�r��p��U���y|��y|[�ݨ�r*(����}k��5r��k�_&**_6�y����ط�5|��Ɗyڹp(��:�+O��w��\�{��᫗������QN�v܊��\�髗9�r���nV���F	��.L�� �fc��by�o^�I�MQ((NU����`R6�~e���E4�h�Be���Q���0g�g:��*�a�/{s�*j�.��T�7��el-\��c�Q�X����Ƀ��Ә�X���_����s�����A���I�JC���JKʍy����N瘅�K%KM��i�a�2ADIe��D6c`�C	
��I��H2�.%!�2�eG%PL��-4a�~?8�#�N:_5�e�o'���<����/r�t�|��9��ZznV�5�ث�ژ������'(��$J���w�nƣ@w�.覦r���;u��[2;�7��WЪ�'v�E�H=�x�gq�Ï	�=3d]�42w��wG�af����{iפ�s�t;���D箕gL����H�\��w�]ݻ��p��T�ˊ2�ϫ'_׷�����v���Z�iÜi�3������q��fDtZ�����ل�R�]�4�\n���{{y!6*�(3㳐z ��zbV:��t�Z9�8Wt��Nt_X�z+g����z.������8���`�U�>��].�*����-��|s������3'ڨ"�D�%�����^K=��!�E�/�b7i���(��ucD�4D��l�N#j�J���
��4�$r�����L�t�M$���^ndv%lΏ;����ґV�Mx���GհI�Z�̗���_A�`]o�u�W�u�7�����5x��o�x�����=F�&<����-е�N?y5�{�~x��*�-2�]���y�ޟB:~�����"�w�C{e�ʟLp�G+Z�'k|�GjC��.o*
,bm�汐�bo(�uTz�0�;37+Y?{<}������I���&I+����6��#����R�{R�S���r��dc�{v�o	��%�{�rn�?M2�9oT�5�/�ZY�����έR����ݦ�-��PV��*�.J�����O���t����Y�	ֵ��qdn��b/��lO�dˉ��l �tǜ��[/�ܳz������#/�����\��XAĳ�$v��ncۻ���V1t�u|���
��R2X)z�K#h����N�h��|�Mӓ~�g&�mohve�H�0=�1��T�Dg��/�R���w$�@ޞ��֩)m����wfT�U3��ޏ8Hϡ{��M�i��:��Ϭ��( &�������7�J3����Y�oD��Fy�܂�s��e�;�wzZ�n"���p;՛�БC�I�5�C�1�̯p��/��_u�|H�W��2�Ń�w������u�i��U��]p#�v�󂤠^�F�f<��Cc�[®9��՗D�v'�dm��y{�~o��Ⱦ��lFl���5I�k��b9[IE����/0���8���u:�ir%�W�U�kUv�o!����x���C�]��N.�������s�qJ����@�!��'�[�!9�T򼨋�e��j;Gz��k��F|�W�i�].���U%y�mO�t�z
E�ín���p���-��z�=5=w\����+=�RT7�{Y�rg-�zvnvU>!��z���z��g��O�+�z��1�9[���4�����+��V*%Ԍ,��
���B�f��gG��\N�=��k�u�8��=&��Pcٕ�O=�E�]
���ג&oVn��.�f������la�D.I���)�vdzE�v�*��E?e,{����3g$ ��e�L"�ߧvR����ԩ"d7WKU?B���T�rw�>�@��D�]��lk��ky�m�*��Q�#_�r�{~u�J�d��I�:w���5�,��tn�W��z�����b2�����w��z��Ŵ<Ϯ��þ��R����*�ݤ躃&buXC-�h4���}�i��]�=ۂ�`���}�hv1Hvw3����sm�N'C�م�w�p�����K�Py�0�a
�<�w�;%�;��<̼�o|�7��f%іWoU�+�����^mv%�o;�@��� M�U]��p��;�4���ݫ+�U�v�΋�|��3`0��]1ت����R{ݧ�8�u��3�PfP]��>8{jy�I�Utճ�������,�F�)X�A�Lr�ڷ;��P�!�d{�W^�Ŷ+�Fww�y�)
���W&ٚ�+3Vj�q޷�I����oE
q8I��&A#����/��t�v�DOu�!g�%(g�1��* xTW�M��]�fwg"A�<� �Z?ZOQK��lR+�U��}�:]xZg�f
u{N���z4TI��F!�b9܏��!{�n��˅&U9?[�}�jaN�^��k�3bc��mʊ���<�f��ι�^�/z���J@9�z�����ә�gB��3���.[�mw���4��v}`0�^
�JDZ2�З�_�v싚����	���(U����QH[�11}WӲ��*-庼��W���¸>��0��o���Xq/P>@�j�KeJ,K;���+hݬ�J)8ݍ�G@��2�܌��Nr��ɝ��VU�&n�Uå[��}'�yx�?s�{=�������lj\h����ܵ������� ��`j�v�dߩw��9!���Ѐ+VϛH2zP'�t�N���>~�O�ND4�y�0X���+��ְ��Ў����$�&=ې�X��vK�VM�c��>�^L���Z��{�5�=�tvc�@\������yN�a�����+}ߏ��K�՛3O�t�6��g�v`�7��E������U-%�g�5�{�:z;��$�\�����Ό7_�P����շ���ӕsV��g5wV�#]�W�F$+|�	ݐc��\m�V?S��ӭ�K�ֿe'�e�?~�P���9w����K�MM*q�6��2���<c�0b/��e�㭞`Hn`8WC��}.+�6ϖ`�Օ��gh��|fm�L������=��ý�E���J�p�0�
�\V#�9�dzE���<���6j���p�E)A����Y�S癳QiM��/o��^_�i���4��ظ�V�;�,˩a����G9L��y����c��������f�(R�k�:�5�U�S�e���U*�Ϭ6�����8�c*9���]�jG�K6e*���ν�#��p���>�"���������x��"o������z=��eR~~ߢ���/�2�;�
�~Ic��U�U�t�y'����dkz�u���W)#<�\s�W��"��bn�o/^����棕�w,ۧY��JkHO����4�ڟ]2�Q�}�e��*s6;����W�mטEī&@�����7�֢��P.�7̩̳	VŁ51/f���mD�W0z*u�7�1�ewWP��e�}��ݝۯ\�oOmM�3@5�!9�� 
�Zt5���l��`z�,d���ױF�����JT�V]:�0�X�ʣ��3|���7b6�x^�w.L<&�{���+�p#����N����vXY�35�2�q�
�Ww47�m�63Ƕ69��ˍo��x)���^�z���2;.�}��W��{���h�G)�Fl������P�>Fk1a�	wO��m}��p��<�3�z��Oܖ!uu����e^�27�ҟT*�v��E�y=Z8���T-��2�-�}3z0 "H�V,mA�{^t�^tS핡�ݢ	-�#�O��t��k�0��H�o앺�j��ܒ�9��srnW�y����g��?ot`����ߐ,����Su�zs�)���=�+TH�}��ٲk~�E?a�~��/!�>#z�����5)�eƝ9��{e�{S���7*H��������iWLռ��{��؍@X�M���1u4V�\.���������/d�;&�Ǭ;x��&9,���0T���6�?g�"I$v��m{8��>�=��`v	����uD4΍���U���֌`�y�܀�C�s��&�W]�IDi��p�ب�s�X�58�9:x�U<�$d�Hua�Ѩ���D����QV�niZ�G�o��;;G67Fu[����;����B/:n�ڒ��̇�O��L6��#M�?<C3ض��ʮ�5v4���D��v���.0=ϨEOO�"�s�҇�7���5�zEΰl����uY3t ��|�5*����Q9��J�5�����¸(���;Ӱ��y2�e�]���vT������r;���[.�Q�Bmm �)����λoNJa+#v��e�S�ڙ�Y
�Yu,R��R˰e=�ۨBչ.ݳ���uh��^�0�y��ܴ�xl���X�����7���RW��5A��t�r"Gf6n(i|��c+P�Xp��qN��n5��Q���#�RI�|���s\����n=�QP����րt�ȭj1>Ty�nyP=+��ԯ�t	���j��[�7����t?��
��B�>�F�Bl�Oxbܶb�������:�=�ޣ����xJq��O��(>�ʈ/�"O-����z�e�:�$��]ݱ5��yb�*��U�_ٳ��-��5�k�u���m�e���͍�����r�&@=�h��^J�݆+g�M�7ͣ��ZZ���Q��k�Ńq�O���"�t��.���B[�=[`΍�L�=�<Ap��yk3�-�َo��<��Kh*�2��(�
q8�;	Ƕ�vS笜�.{z�MJ�$l3�\h�Ψ؊�k�1���3;�!L�KV�m)����|�n��n���`�~�]eG�-�g�%-ۦoհ֑�4N;կ^�_<6���b�3��a�:�I��d}��Id� �v[�_lᆵmМ4�}[��wJ��5X��D��×
Ɣ��������WKl�&�
|ɐq,}��>>�wv�4��'��g~���{�˺Vㆎ'l<v���2�L1"e��!���������c���Y:�SS�.�l���%,������^�v�/O� IW��\����!��0�k�"Jw�M����W�ַ��8�q��}��8	�i�g�l*��XC=]A�m����95s�{�OQr6�O���qJh��=X��z����t����3�hv���6ڐ�'#�=
��L�P����K�\��l�ܽ��蹢S�g���ܳ!(�G�x��������g�W]�#��Wv�g8Uy��/eDX�pk�>�1���\Z�%h1QݓGw2��FjER*ۤ+;g����S����n�'��1)�E�ؽ���jȋ(
�R��y�T�~�����7���m���=��Ad�5	�[�уO��&1m�;�D����6�G�i�bT�5�d�{��Z{^���ݻ�]%�^�l{ދW��Mֺ��,r�Y��T[�LE�q�Vc�B��]����emБ������n�vQ���s��z�U&
�I�.����ʼlS��v����:��W��<�o}=���WG@l��'����p(��^�Kh$MM]1a��C�T��z�M�Ja)y�,ހ ���@ˏWImY�k��o[b�`�)��G\_vE�ooj��"<���X1m!Sm����=E�b;�By��R�������}�\k�O_Pg�u`#!�Y���T`�F����\N˜�ڝ�Ȑpi�H�f���!�˙�W��{Qr,7]]t�]g[vg�v�n9oUJy�<�U!����#b���k��7��Q�7�$�30�$[���9ә������>�IPH���\���Y�5��&hVt�wV6�k�!d��]�z��Fob!Y�Rp=�����/�E��f��o_wn%{�74�43w���/�RaP�[�ݒ��C���F��_VV���2v�U7�g�����sS�]Y�p��oD�]��a��s��}���v���-�&�\�q�Dy�M���M���k1fu"���W}�yMyR����$��s�^��sX�tQsXj���k��J�,uF�C|�;��q��g0����8غY ���n�S"Dnލ���F%�kw�M� �l��� ���	��=w�aF��L:���n�:hc�82Ћ��_U�r���H���!Ro�f_j�{����ɪ�*F泬��>go�����u�,ޫ.0S\���ORw
u�M���d;F/lӍ4d�So�r���P�w�g�a�erv[Z��*__��ή׆sN��Y��s�Tg��Z�6���:��S���.������uA�RQ��{r��91
�L�v�UƷ�G��X=�'�Vd}3���
3ܸ~Wǳ�H%�-�a;���<�&/�ј�w9J�v��7ҟ;���N�|�F�m�W�Ls:*�*�|�	w�h9�)�f��ԓ�VF(�Q�r<�eΤ{.�<�k�����31��(?+�R�7���l�5�"Ӵ;�R���r��ۓ�GΗ�	��h������ʂe�����H�p�P*�����v���!�wb׊�/��2^̍��[
�Tv�s*k��A�yp*�e�5Y�K&�%,x��yǯ�
%� �v5*���	��w���n2c7h4pf�l,�ҭ_[)�M�sb��"
���� �ъ*Pm�n�$� Ϫ��Ge
��Đ���"�(�`�7�t�2��
͓x.��eA��P��z#���Ij�x�	=�ۮ�za[��n�T�g5����,3:�F��c�<���f�Ov�Ω8:�<�|l2�����dӣ:�*7}gD:�:����ob[�G
ۚY�vUUN+*B]���We�v�euH����*5N�WzHۼE�M62Is��y��ݝ1^h����m�&�w:rh`ԡS�X1�۾��ZJ��ь����&85����e�L�ɻ�2N���X�Gp����;��\�y��0���N��H����]M�v�`nƔ:��H0�qݜ�)����z��!i�8��˘2���ͱMf�cx^G�cظ�s4H�i�ˡ�*r�rѸS�c�.�z�f��՝�lk!��OW,�$9v�%$����{y�a�Hf��΍���1��y����S8����nN4]Y��h<i��T�P��[Y���ۮ��X%�%�]�:���:R.�y,d�y�%��c5`VH m�Jl�ӤXYJ�uL���k)t��1F,�G�Ϛh��'���:b��꺊�G�;R��Y�JŅ�W,���\�̡�*�-}s�k�э��,V�v�����I�9�5g��-���Sw�^��Ҥ�9$�S{N.D$�������W�w_��ɷ��˕��B8Qߎ�ݮk�zC""�ێ:v���hֵ�kZ׍cZֵ۷nݵ�>"rLø���I�#|�rC���zN�s=ث���~���u{|k���ֵ�kZִkZֻv�۶��(y�b���L�b���nnK��7�sc�w=k�+�X�W�7����/��{�w���ݷ�����N�E�Źh�d�\��/�|cQ�uw~/5^�س�s���"wQ�����s��]r��:�jez���Q`�W�sD�b׽ץ��{�ߞ�������o1����{n�*��G�v��9��G�y~�|U�ۥ|Y�m��/6-��}��u˜خb��ך(���|o�"��ǘ�������۾�<Hc�r�1��A
�n������%������s���n����������&�w�.w��g��{n�fAM�������b)�'�כN�=������rg��	���h͘�t-�0�������^�w�����k�nϘ���%R����t�t�y鄷>�D�dMu���l��A��5����7:������N$6c���A�SN�m}�$jn��Ly�,��"�]14��2�9�{eT�i��x�N�&���f�+�7a��1dGFϫT��*M?��y��j���ƙ�����	��]U���}���ն�+`y����3��Ӄ�%Vj���Mq1�q[���>�nI���e�[7�o0(�m��n�)y���s���}3����k� �wI��.�����}�q�X�d]�6���k�=�37��9���I��s�Y�<�$H����g�1�l3��i��*�s>���i��>��*����C�r*B��w�緰i�C�	�M�|���ʕ��I��v$?�pF��Cߪ���WY�ID`ҼW�v����+���/7�ӹ	:\C{w�5��������}6�#�R���Uq'���*��̬ש3��}tٕ%k^���h�<���jV+��:���_@sr�:�4޹v�Zf�Cvb���H+�esj��*��Sړ�vuN���fl�w���ޣ|8�[��r����`��C�s"�ԝ�N��C��+{�tw�����m�Z��!�f���>	C�OM6zr�	X�C�z�kw��d^7Ḋx�C���E�EI��4��Oh,�+�`;�ɶ�z5�@�jkp���Ćc��Uڌ��.yN�ٓ�x/N��DkI��f�*s1j�1rr�=�����b;�q��$Sc�Y;���F	~��-۴���N��ө����1�V���Ҝ�nH�з�{��Y[�ʇ,w��C'���4�/>u��t�c����#tQ�"��6���>�?��b�'4����Z�}�|h�W���adz�.���cdV�~�7s;�sn>̏ з.������h�o��S�
�y�y��kT5{��/�s�bd�u�M3�Z��Q��<�wx�6��^X��1AV齏t���Fl�ԥ32p�48��)�V�����eV��OQ{�2=�{�RY{GrK>?|1�uz[�1̎Y��C���)?p�D*���I��B E�����y.�iʕJ����bT���M�s��R=g`}��fi(Uؓ8l��%Y���^�6wu5Ͻ^o7�:̤b5�E��R͊���,�fU�"y=���v���mf����c��ok���� ���	�*�A�����1���r�y\�zy�dEd�8ځ+���.��<�#�`v�0�n�1d5t��n�����3��5@qA��$xO8�TP7�J`L��s�+5Q���֜�=�cx�lM��n�m�^=�?�OR���S���b�F}9��r/a[���.ޭn�E�؎��ϖw��Ě�!h{a�.N�b�ŋ0�����<Tl����v�Y�u<�A�����x�#O&�{jz)�a��t%�v������j3./
����lω�i���*ʷS�KJ�������Q�g7r�0�Xa<3�E�l�u�m��Uv��֌���۱��a�����?E|�7xsw�t'��߾^�!�n}�5 8�`����գH9�к��g���ռ7�fQ�����^�O��,l	���Q�f�)E���2��������;C�����>U�:�o{ՙ���m��ӅUI���*�kޕ�3�-�����vj���&cʏY�F�q��G��S%7}3���*K����\8̵̕1�Θ���Owk��>��DY'G3}���yN����}7�u�ޝ��$�~�oK�:����#�<t(V����Cv[Se>,�8����o��i7�a�R�������Zނp�9��7�x�n�[o�h��A�ZZ��#���H���f;���]L[gh�n�v�����iӇ�t��8fDrٽ&��bU��	ݟ\e�͹��Ty�ݬ~�ۂ��r�y��(|���Ĺ���K��tl'�޽��Rw��*fW/!���@�g�|ݒԦ������L�h�w����ts��^�b��T���q̀�`>ّ\
-r��E�#�9<��8\�7�4멑�vwnv�����c������V��r�m�ώ��Tma\�hh�u���R	4�C�u���8�:Yz��cX2�j|���S�M]�U��έe��V��t���O?K+j����;���Y\A���#�>�}�[(�jn�CsF��pCO��,8�,^%���{�S��t�2��j\��Ǖ}ڙ���MDDr�V�M>��mn�X�w�����W���v簢m��t�^\ˏ���w3n����=]��Ot[�;<3�L|1k�V�O�)�i���q�ޓ)s�޲+��8�L����Y�j
�qj��+&E5���Ad5_�dmkVpk����ݦ����{2ni���� �,A�3�+�Yqx�u�xgn��Wp䊕�2���W��s)��<�9�I\NK�kp��g���j�pݠ�:zCa&�t�OX$IrS�~����S��»��*�ꯈ����ќ@~V�맯G��$
(��&A<���!��2�=�Mjޮ��[
(9�2��w���6���(������B�biScem��sԥ\��������kT`�[:�^T7��W,�����ۭ��
�h�v~��Y���TY���Nc[w��g�w��v���>äɘ����j�0#6�
7l`\��1�'�34L4���bM�S��e:.L�/;G����z��yyۿR7x��L���f�kQO�->���x67r��F�b�R\b����:��z��xW��
�}y_�˫�����ii{�HNZ�Һ`����}������w�h�]~���{���_N����Ӈ6��>��ܺ�т��ja��uG�rc�Gd^ylܓ�ϲh;w��װ�j?����5yH��K4����OL0waNGo?����I������2;��E�	�wR�O4�zZ�Z���jh&�0Q�ۀ��|�IU��\��|Q��4ם�n6��m���hWY�-�谞��ѡ諚�ff���{�l꽃��޲����s_���8�!#:�{��g��XJ&SI�܍�s�4Eer��&��W0�q�uy���Z�x�Q슉�A�؅��,IQ϶��D�^\���fb�܉ Ƿ	��*���.�PyU̞�xM��kb�ޣU�-��ϭ8���A��ye�F|l1�k�.bL�ҭ�K"��e��\vc4�l��$���ld ��^`�@i+z��b��в&�7��(��V�h�-�� �j�2���yTy~q:A�/W�˚Cʒ	��%L�4�6Z����u�>DS@�*� ��D�I�5�}3{��!��عm�:���u���!j[��t2���p���ʐKh
f �p�2����x���+����
�%(I�j����=�a�i�3M��M*�.JB*��U�Sym�
Lg��uz���V���u�#hǡ_�y�nyPN��&���_kwWuΖ+������������uǗ�!t
1��I�5�;j�{o5�ev�\%4R+��s�3�6G�|�|����S���=F�>�_wmƮ�u��������<�����HU�&�=��l'�f����F�NL�����fz�Y�C<O�o'лg��g�wŵf��J�t���M�neAظl3ݛ�h�opo'CB�Ä�=��<���~�:�����떙���=�^�j�1�B�L������P��N�mN�nKL۴�A��w�	�5�q�uS��d7ƻ�y�R�xh`����2jK«s������;rw�8��I�h�ק���yY����.6No<�w8QI����tr�'O&��S�t���d��|�&��	_����Y�ޠA�Պc.,�}��M{�ꚻ��h��uf��f4x׎Lo����8�v����.ƌ�y�oV���ү ��v�I�ec[u�kO,,y`�V*8������z�L�7:9=����fl��2���ޜ��$��\��f��e�u{�ȣFI�i�^�[ߗb5CS�R�=���X�9�n�qm���
�k�)Z0��s��𜣝��ƺ.nb]M2Cn;&��LyY�m��Et.�f#ki����裘�n�+а�>���������@̆��JqFO*5KC�Ny>�Q�o7����ޜ����N�_����"���je�A��wn������/g����1��oI*�4���K;{ky���S9&E�Xp�@+���8;"t�GMq>y+�~ھ�E_g�˓�1}��[Jj{M2���ݲOOt-�b4�vc�h�c��D�wM��X��vgU�,Φ�����LDk8!����zDF'uO��^�>M��5 c@�k���kIܺ���>��#h���z_~���&L�2C�vh�W��^}[P��d�u1���P�{�箛�P�y�0��YZ�5Mk����/��ˁGVX3�v+9z9�tǣ�y}�t�և-�^JD�tZ�	��&�\�@��Y���e%*����̎7��fMŹ�v�y�;��c	�������}��j՝B�s�n�Q�j~c�!�s?�s���v��Lc�\8�l��ތ��~h�}����>��������!�����46Tj��)��ɮc۝�]�}�b�n��H04�G`��.X�e���'%Z��]]�,�Up�wU<�a�����h�b0=[c��r�5����.��:����X��>�|Ԧ�y�Ʒ�o���������;�;�{�n����+�	���.��Z@�q��}ܪo,����o�޾�$���֏]��9�PdF[��n�!g�5p��W����۽��[�C8j@���U�Fd�܍V�E[�(q!<��i����u�1������yv�t����I$��:�ݔ��<�K��SS�X��׼_D�%����)hn�"�l�ywp�������}|�R�yN��u�6��ժ�`�,n#�����N\�5���Xe�t�#�N�ٶڄY�?Է|�݇V<��N��(b�7v�j��	���YÓ�'gs��:���}u/lT�6����t͗�������[����Kq��vDO�lŰ�")8�ݞUd�;a��kg�����e�;#��ook��%ɺ<ք-�@���@g�Ѳ+T��[ꌧ��2�""�|g�mº�"gN4�C�S���6X.��硕�N��M�����~������Mx҃U�6�= ��#y��G��1���Cv]^�������K�-��|t��#��{SA�}�<.�.��1oL�ᾞ��ʎ!r�[Vߒ�Es����<vI,�>��Eik�Nr�ڙ���ݹ�>��L}��>�:H�1���g���&�tɡ�f]f���4ES\d3�pQ�}�&��#}�VWo��ʐҤ�W��6�<gJ����*~}U #ɏ�* ~Ԥ��)�q�����S�����[����dqz��C�ɟ6�Ezz�f����9�u�?���_����� \�b�����(舀��"����0�0:�Gy�0b*,���-��T��Y��5�f�,�e��f�,�KSU,�e��eT�m�[e�R�jYm�m�ԭ�[RͶYj�j���f�,�K6�e�Z�T�U,��Z���e�YU,�K6�e�Z�l�m�Z��T�m�m��T�U,�e�YjZ��RͶYj�UK-Rʩf�,�e�l�6�e�YU,�e��eT�ږm��l��Z�T��,�K*��l��,�e��eT�m���Y�K-RͶYU,֥��f�,��V����6�f�,֥��b b!*��}t:ݟ�V�f�Y��6�e�Y��5�eT��,����,�K-RͪY��-R�T��,�K-R���5RͶY��[e��el�m�UK6�e�Z�l��Ym�mRͶY��-Rʩf�,��R�YU,֥�l��,�K6�e�Yj�UKR�,�K6�f�,��-RͪY��6�e�-Kl�m�UK-R�T��,�K*��ԳU+mRʩejYj�ke�T��,�e�T��-Kje�jVdT:�P��@H ��Q�(`1@
�����+UJͪ�Yj���j��Z�Y�U+6�R�mU+5Z�fժVUj�K6�R�ժVUj���YV�+5�R�Y��JʫR�V�,�UZ�j�mkR�f�j���R�Z�{ޭ�VV��f��%��+5�V[l�f�K%�j���X���%��ݭ�X��+5��֥f�,YmK%��YZ��jX�Z��Z�����\+���YU++ef�+6�5�8� b��b�;b��`�C�'p��;����h*"�
�� F'��g��~?<�_p}�>��h�S������������?�0��?�����������  U���������(���@_��#� �@bG�O�/�������?� *��������Ӥ�����������~a��I�X
(�
�D@PaU@�-�E��F��*�Y6��UTZ��V�f�T�h � �REqm���USl֪���R�mU5MUR�kUMSUT���R�Z��VU��� ��@"��1@�U��U�@���m�j�R�j�T�6�ZZ���[*���4�f��)U3j�m�6�%fD Cz? �և�������""2 �$�  �H(�?�� �������@��~��4�y�>� \ف��.����y��;H~ o�����I���@ U��P���|u��( *�@ r������4*�����:� Z�����-�C������Ϯ�g�������� g���>�����[  �OS�5�s�������'���?�A��?�}� i������ 
�p�6y��!�H���S�	����?����s�ϻ� W��H�>>�b���<�����}_�*���O[@Qrg������b��b��L��L��^�^� � ���fO� Ć��=��6m��[VM�֙Vա�XLf���m5�J5K4Vն�6�ڴ�X��l�&mC4�B�kV�-P3kM�V��Vz�6�Z�5��6̂�k�Z-���kJ�U�:wkm�����UFb����2��(m��՘I�m�F�Y���(�ɵ��֛5��VUm��V�T�j�MZ�b��	Y���ԣ�6ll�MgwS��M-e�[V�M�ڬ���ɴ�em`JͅcI��Z�[#h����6�R��� ��k0���m��b�R�i�Շp�\� z��)���W 
�a�8��+��wt�n�:��-�wz�u�{�kL�޺���5����.�U[��{��ON�v��S�J�.v�KB�Pˈ�Ҫ���jm!b5jگ�  l��(P�B�St����Ht4(R�Q3ׯB�R�	$R�{�b��6�_{{�[��ӭ�\iMzGj<�N�iWww[��aCOOM���*��Mmָ����Yc����F�lʶɪJͭM�  <��C�����빮�]wd�n�k���m�+�5z�+D�Ү�Bweu;a�l����Ѷtm�ݔkbT k��v���׹ҽ9�ӆ��U�R�ڃcY���N͚͘�T��   1�� ����Q}ht5�`�i��}��V��ӧS�8t�@cU������]���uN�7j\���]V�ZE]iݳH��Ͷ��b�j�U���   �@+�hUW�jr�V�e1� зj�n��W6�v�]kwSvT �q��غ�p�l�9��� 6K��AhkE,Lf֪m�%x   w^մYͼaE]���@���ή��'Z��w]�ô�h�]�u��Xh���4�US��+@��kV�*��ZֳV���ż   ��  u�\  �������
����  ���  v�� ��  �yv�  {v\  �kSjզͥ���-Id���   �� ��OnӠ
 �wwp�h���� �Q`  6�p
��vp  6�p ��P �;��  ��J�meLZ�RF�j�{�  ��  ����۶�  ��  �ٸ ���h h��� ��� w[8 �ݔ 
�ݴ��f�4�-��}����)�  w�}� ;�0  s\ z y���  m�� �c�:P ��� n�4�wN  =׳�@  E? 2��@ h �{M1%)P  �JR�  )�CIJ�� �D��
UA�  z�"&ʪj  �����~?E�_����_��m�D�dU�a�)%6&�Ƴa���[`�4������������u�k[o�m��kk��ֵ����ֵ����ZֶͶ�m������>��������M�or�����&@
�Se�)�F�6N�a��>�õG� =�^6�Oh��ǤfE�u2�U�vb�PZ�[oo y�pٰ��i��Q&f�)�����C��8���ËV���V�h8�Z�XfY��T�Y	^ ~�0] �w��.��I�.R�"�jԢ�/��F�HCʗ��сGN��j�r�PK!�W.|q��a��'���
�h6n��ۦF�x����4��:���`H ����k@Z��
EbUw:toJZ`�����µ2�:�H�n�uw�ʨ�B�ͽ(8Eзl�O�����.�ҕtBEk�Th޽�qFj6,AVգwe�M;Z��& 5�)[1�����)��)*%x��M���B�2�$����W4����tݤ@Z�J��n=�a���8��%]�a:�T�W���񳒷J���;����N���Zۺ"<y���-+K�b B�ܻ?Ma��0��y�+�)
��!�Oib�[[��Q$Qs(���»,�Z�-V���u4����@n�؂�@�h��@6^#N����̎GF(�3u�,#��+d@����<.*x��\i��S����n�.���ۼgZOn\ܠn����Y��,��Tŭ�v4U�/6=����7nm�t 9VY�0�]�b,�0�H�QjM
��R��e��� +oc�YIF���C#�4�v���*�r��ʻ'-��ݳ�h�t��d�&èN�.���	;� 4�:r{a�Ml� ���#����J��P2�mv��GEt�"�E�v�I�y�-���%4F�#o^C"Vr�,�����wG
Pަ�u�0������Ei$;��*���a]�	��WL�*ûkC9f`���v��BP3ZZ�V��D��t��w�[ɚ���c��pQ�J�;n��f���5��\�*�(T`�ґ�Q�/+U�?i?m��[�,F6�+7�6X)��4�a�K-T;Ep�[���U�SF]�QX�N����6��Ÿ��,fD�E˭aV�St$�{.�lq��?���h@eM�	��<���Z�'E�J�Z�dcY r��e�ÎKp��OE��e��ã�EU�o@�gF�`�͢U�sb؍����2��t�	3V�̨�F�*�֜I���9��[;b[���&��s�\�N
�X�MZ�(��)]$�]�hr峍�`;ݭ�f��.cEcӓD�qc �C2����h�[�g��9� �
�9Y;f!Z�������J���]r�.��C��XΝW�GM�Zk
4Y�1�חWF��Z��0���&���˽�`�VK�e=����]-�kn|��,y��Hf���d �R��˙5��-��X6$�l	M�f'�ZoN���,J�<��;��`�Z�N����Q���2)J�=yj�*��AQ���%�ӡ��-ouB�v�XT@=��sA�.�
��ӄ����0I!+I ,�na�kü�y���s(�A8�;J���w�5޽�i`�X��)Cvco-��Mi[b@&m����qY�B�X2�))�t�G��Z������w%#����FE������D��QЭ�*-�
�PF,�.�M9Uk�ʥ��=L]X�m룩v<��T,�EC�SkF�����k�c �홋q�,��Eh���x��l���j\w%�0�x�ze:{y�sn�B��X��jj����W[� 4�I��ki5����D�*�2�p^����L�S�hE1�4)�%�l;�j�9"<��h77#�ĥ��[`}(V� 6�s^���j�m��V����6��b��n�NX�F΅�U�T�q�zv���O�4^���R���#���n@u��kv[,h*�S��uI���)K�+c�[�B�����*ɡm�X8P�\4��:I,�o%X�w���>K�����k�=Rkձ(�^�YX���W��KRWM�o7.1B�=WFc����y"��1P���Hgf&hA�b�v�̂+U�8M'�YG����m�үdm�{d�ڀL��Y�V+[z�COM�܋!�Ǆ��M���[�o��r��,�Ql�aD��7�ݔ�laa��vj�r(���5�`ЙH6�j.��:9@���5�ѣ�V,mE��c�`֥���ƴ-��Tݲ6�6�ض+q<��zY�ɑ�[n�cx,&����]�&*r�EU��;{]$�|�[D�"��l�DBޫ�;F�`�0]�X�%�GiՇ�So"����;J�	����	
�޶�u�m��c�S�oB6`���� ��ƅV�1��@+"�� �),%����!F�� 1��؎Qw� ш^�$W�,Zf�]�Ӂ�/ee�BioR�(��4͸�k�ǻm�����hXsv�[nm��g9��"��T�`��;X�[9���,֭{`@۳Z"��qf����J �A,��e-ƙh0�f92���A���l�)0ʱe�)4��u�4<p;D������Z����b��E��M�V���Y��[�Ģ��e7�4=h:٪�I����,���U1��]Kr��#�Z�Uiaۍ��!ܚ��w6�#N�0��v��T��k�����*�2/��2��d�E�F�,��m;Ri�r��`&*ݖ���$u�^�`�Uܙ��J�0:QHe�*xm�*�[�Y��ѩ �rE���P�p]`M��+41��D��ƍ]&�fj)*T*0�֍;N��NV��Qz�V�m�n\ś������qŊ�IAv�P�Z�;����>�(7����Bv�MRl����*��u^@����vh�Z[�M�tt;�[�1w��J)b	�� �d��"�����N5��a�#0T�-����
x��ғ*��6�J��ޠr�
UJ�`4e�fn�*�`V5�p�J֧w{w�`���ȍ�363Zb�j�
���aV4�
�bCt�4YՍM��Mu��ǆ]c�iʖ�mDܠQ�3U1��(J�����s[�Y�+>N�l^���fI�2 ѹN�	����tM6�0T��L��ik�WEZ��T�;83�)K���*A�%�5�N��B�6�S癉l�$-��mcA��V�E���(���B��-;{Bm�Ug�F�ix�Z1G{k3B��BT�� U�+'י-+B�[l*Vř�8t0�Y���BL36�`�����ӻ�b�ȕ�XK�������&��/E�3I"���{�B��1�e�ᡭ0�,���$2��U��uhY=����W2�QSK�����Z�4�D�B���pP�X�W����7H۽�k�[`�M��p�IK
��V��b���kq�t���C�5{Y���0��#�7N�]K��VQ��,-P�`qlY1�A�,+Ɛ�Q��j�gq�Z&�rn�����{Ywy
�p�Sn�����"V\P� �d�N6��!X�^[/Zbo�9q�S"��@��2.���	wf��[����,�"JMOA�f��m̫��]K�4r��tZ� �0��Y��`��f�:�
�CH+���]��ڼ�N�p%E��n�m-�T.�����Q�h���ª,9��`Til������H��^j��%,�E�(V0*ښ����̆`7ۚ�!v�5�ƭmFk n�Ïl:"a�b�t*�&�S/4�Q,���/	�B�ofZ�%DJr�Fm'�+��l�pmL�"�[zΜn�0�]��%��!�%\�vrn��ς-�V�&�T�oZ9�I����w�����wv�	�^�b���8e���sU	�cIG!ٙ�ޫ����wYi���).H�_M1�
�U�芒��������8d�u�[����Iw�����7&X�n6[b6�=�VͰ��(�΂܅�N�:1�ZJ��Y�gǵ7T	�Wt��&Ȋ�df�+���a����AYx��%H��&�/�ea��6�����X&&2��3ӵiPGC�SX����� y��b�������[y�',ϯiT�NI٫@(���U�����m�t�Vj��0E��e]�Ѻ���n匌K�L�L*�76\Wb (�O���#G(�VT�)�����
��4FFM���*x�:d�*M+`PM�騥��\/]������f�D3d�N
n@��##�N��!�F�m�ǂe����$�GkB��35�6��
4��k\���[(ˎ��M١��VV�v�-Ԙ5�	���M�@�iU��|%&|U��u+LX5eY���;��Z:�Ÿ�"�PF�E�$�ˋ/p�r�-�Z��f��v"Ki��eS�n��@�umf� �fV��5v�p�$ͨ��ܡ��&�V^ݷ{��v/Y;����e�����΄�sBY���Y�=J%m=q��7��.�i+��R|��	7JR�`��Cq�[�K r�cu�=�VG��y�0�v���b�"Ie8�$ƙ��۰��$����lI{)MǶ��ܥ���F��%�����V-��3��bD�^ʍ��,
�����Cm�n�ƉOǹ����I�˔rf�n�ZQ�3n���X;MM�1��@^���Ś�5#�ʖ�R�{A(Iv�2���Б�W��#(��h���k]���d� �7[�[F|��m$@ �w ��/cu�%Ʊ��{��Ъ���h�L�~������[���H�T� )hFe��N(�8�
���{&�ֆ8�hWE$++nR�Gq=��fi×��Y%waչf�5�|�J��]�~X��ք�c�h� ���� E�6��_Y�x�D�г7*�M$�n����{3*����͟���RN��}���wj-��r
�۫�V�j�u��5�)�w��{y���Ś.�K6Wٮ	��ސ�j��:���n�-�)�Y�^��3aDV^�0^I{�4B��(�v�L�iAoduw��qX�liە&6��&F��tBX�D���x.���z�n�.;�\ɵ/P0D:�6:���SSJL
�j;r��JNۼ�mۨ6�ӳ&���u����#���☓��yxqVcNm�%0�v��ǈ�^a�]�9h�b���V��Mm�[d���Q�[OR�r��	�3h؇[��@��n�F����f��2��f�V�j:�/)���e'�FJyQ��;,��2�T��r,�P\�o0�� A�.heU��@X&(l����Ȱ��޺pH��'K2�4�Ҩ�H�p]
�Q@޳�Y�T\Ȁ�̖ˈ�Ӳ%�S���ÖI9a�܇~c.�B�2�!^C�u��&
��x�:&��&�b���U7Pڱ(_����+!7+ّ��I�q^��{�D&�_L[�{��J�h3[��r`x!;q�9�`�5+oJ�>gU�i��m�0j:	%aQ����l'Ws�)]bގV'�HlR-7u�I%)�����6YiuqT�)M0�[`��{QR��]�J�^���e�o`����}�)��NMHH�'�JC�XRZ��"�\��7u��Y�N�R�6�m�i�o4�R�)nT�^bW�-&��5�i�+]l�FV��x�el��[���S	�f��>yZ͋��*���J6R�c2�'O^���u�Qc�f�d"����`���J�f��w45��t�a��֪[,Zc[f�Q�A\ʹF]� {z%^��5mZ����Z�m���6��,����.:�!;{im��.9���U,k��-*���r�Z�Q�nk��3�%�ōx4���K����AL�F�������MA�li{S��������Zi���C-�y�\)��Ʋ�MAX�7Piu�� o>4-�XpE���0�'R�$V�-���7o^;J��^P�&c�
4YE5�Bʽ�3-�]��s�Q�wv� �l�Ӕ)�L�Ө#�F;_`$),��h�-�6n�u��6/m�ȫi�4� ��&2�Pݹ��ɢ�),� Ӹ�R��	���Ff��h��h��2)ӛ����B�D޳����� دtң�Đv�c�{Y��`B�ٸ��� V[I�rK��0)���f��[����0B*j܍L��
R�e=F[d;�R��n�2��i�j+2Z.��0�O��{�K�������a��:�bQ@Z�5�M�f����O&n�a)ki���Y��q��RƵ+RbI%!��YX�JjF��Yn:8�e<D"�L�mf+���r��B�%%.��m`%���	���V�+R�m�$ 1�q�&jm&�f���:t�j�FQn����8��6�7������ƆN�b�oA�p%�[Q G2°\T���
�m�2�%9C5�{D$0em�\x�՗a�T�G����Q���*�j�R��&�%7F�$��M�I��޼�\[R%i�O6H)=R�A��VSyV����me	�kͻx��q2[T�"�e�+啪Z*��.�r�AKkCG4k�W�V���3u�Hب�e��t��Zxb��%q�I���ѻt�X�[`���APx���+.m��An�q�Ƭ��&EZXF���v�]�c.�aƭ�#�5�:�2nTz,���H�b�^J
��z��X˕O��XЃ��q�0��2�J+�x�d۲bLp���2�,�.�+� �ҫV�wP��N�SK%�Y�ܷ�,ܼ��^�HPZl���{f���Y��෈�&�"\�J���I�pI�\���oi��0ͳ-#j���E7c3�-/��Va�823%F�n�?����t]��3e�ys���]�C�[ީ��rCm�g���3F�(�����#�9v�;����[^��<��qRT���Dk����;D���܌\Ev�j� ��|T7�s�����5q�1ΖY��[X����CȠ�2��vunPg@R�6�60� )��2�Cx��N���<D= 3��5i��9o��\d�*�۱u�1����3%
���k����Jc;�+`�G��/%�F�M�Sb��q<v������E�Cm�[wn�b��+��Z�9huc���_.�]��9����]#t�G����u� ���8��ƭ���Yӊ��j��Z����P�6���j�)#�v����DxQ�����q	:p�T��Sj�*�w2�ȩ�]������[��++K�N|�pt�]�+�ˉ#r�9�=9!��)>�l��]���*�+���w�Z�ySx�({�|fj0Ѿ�U����9��EE�-��A�K�v}�=�o5F� 7��
q\���;�����yRmB]l�wIw0[�`����蒄���d0v���h�n�y�Os���2��(嫮Ǌ+Ү��ŏY�c_��7�a�JÌӾ��ժc�H�Wkza�����K6�Z�Ssw\Ǩ7ȃa	��͇��7��W�x���KR�R�Zd�(r��}�w8ؾ�4	����:�.�e$P�,�e�v�Ho;;Ԧ��L��ރ�����Ǥ$	���sة��Z�')����v�
R��^R�(e.���D�w&J��E���p��לee�4˳���iP�Fd΀8(od�.�J�|��Ms�W&�%�.�.�kc��|��M��r��. ��Uv8l�-�`Ei����o^�����u�Z��n]1��a��D����(��Z���-�+c��;@lY��(f�V���u�
��X^x�Se�$�����H�F'��Iar�I�� ���ۓ�yQ�w����(u�U��myZgpr5ڥ�Dwd�b���$`�ZO�	y��78���s�ڌ�p ';�����{�O��x����r�x1b�s�늟h���B�-Y�Wy�&	�8>x�'3�8���nc��"6��aHh36B�-p�� ���0 �J=�$�ԯ��oV1E�]�I���v^�tu5��B��̐<jS��ν�Z �ކw֦�,���5��O<�@�)Y{tBR�Z#&n�O���f{+j������y6D��{u��~�xSO����5�;mj7�J��A&�LEWn\��g��u��&J0�Zo����˼�`-�0��\ݼ�W<q븏�1[���^o��N�hw-�*ژ���@ �B$G�ʬT��a�2{`����u2�WkӘ&��k3{+,j`x�s��*��V�;;�f�|>����N�" n�t��Cڠ��ט��	)���wK�+�����z8uKA�X�rk��֨�y*΋Ѫ�˂�'�Ժ��ݻ��0���Na�`G����9�3����p6�
�sy�S-e�'Z�3Z��f�#��������heg���輻�y���i޲ehR��bT9t��m>����[����Ш4U���2X�0Q�Z��ƍ��{֞�q��9ܖU�jfά�T�s.#]"�zUM	J��}yΜ���R�n�Z�4]@Q�K�5�
g�i�e.`��zM ��[	$�b����Ny�wZ˜)egZ���eƭ�1��vofNU(<�]�{	�]3׃s��6o�vC�n�r��{=���Ij[!,an�����(xa�`@^֚+�Vu�������+q�@�J�o�[Q���ė�۽��9�s*��i�3�&��3}��n�=�s�Im��jMD��>[f��
U����M����=���3���]�������jp9}������J�k�W[��Z��G���n'��v5[Eݭ'�Їii��V7����x_k��|�G�dIR�ٔCH�ìB���C�oggbz�����+��u���]�TX9��<��:��=3{c����ڧIUocl�Rj�e�7{��p;�њә�;�7i�ˢx��Y�

g+(X�!����Щ��hT�]ފ����n�� :wXR��w[+L��v��B,j���w%s�|��}�{�v�*-	;w���$
1�v����_oxb��a�Sku�XB�E/+z�eø[g���h����T�	���X0�������NP9r��pՕ�9mn��3q.�1��6�16:��z�C�|����9p�p�(�ݐ�s6�i����\��s�a�2�R�v��(5�g�ʊk�}��}��Xn�y;O�����:��$��}t�gp�[U�.t\�j�-���Vٿ���Or�ӷ��
�48-����=t'�a��%��¦
��9 n�p��Y�æ��j���˖J���1�}��upe\�[�t8uV�%5���>O�+�d�'u��O �]�w���.��]±��4H�QN;����()3�.RZ(���h��%X�`�u��q��e��s�a���Jծ�(��n�'wZ/v������'�(�e���u�.p,ڗ�X�0Q�®쵃�t٣D�4��lM:(���Vu��1/o�uC&�4c�=;i��DPͶ-Ҿ����R���T��Q�g\An5\U��i�Uڣ�\�Ъ4v���wV�����[I���z&�3�g3�r����Z��k�Z�3\�6ͳw�:� wC*�c���t>'"Bi]�l��}��K�8�O������o���>�R�i0�
�jL6�<�Sfs;z7��t���.tI|�� >ܡ�R�=Ơc��ѫpِcm�h�f%q=Q��P�ütU�3��������9k.�'����z�-z[���vpH4�&=�6�\��
Uͺ9���2�}#Ϻ"�5q�5.��0<vS'_"^c�4�RY�+�����:�����Nc��/�U���6[�2�C�)�h�=k�o�uk� �1B�R:�U؈��,gn�
�>Z@_tY�!V&@��g>/jr�]m�J�󾌥f�ʵ�˹&��xv�!��R ���]mlG$m��`�n��{T6s���v3�j�D���b�N�z��6�U�e�WA��r��@dO�����r�{��&>�)v[QVv�04 (3���Ԟ2';ݾ�kz�Xm�]e�2���+>i&�+�L�J���驅��P�+;AT���e��!�K�)��N�u�e|�B�S����Q�d�9�.S1�#�������D�Z�ww��I��`J�0��ޫ�.4�T Z��&�x�K�'@�y���J�@�j�r�F��Y�u�=R����0ܕ}��ě�w$Vw ���*c��j�ήY�6ܼ�� ]��{ѫN���(�q33�J��t�q�LZ�O����Q8ѩ�Yy����[sʱ�1$���ҠCY?�����\���]c��Y�� gY��Y�Z:l+��;�b+ ��,�NՍ>��릵)-�؃�K����35�[\�1�#H��
^``�Z�I4�m�$�"����y��0:i� vi�k���3����ˡ��r�b�Oh
����ܝ-4'|q]��ݻw�g�+EZ_3��A��-��r�ۉ��t�\x3�@�����o�,��
�Q[hur1WV��X�Tx�k�K�ݗ[�3V�8�.�e�u�5769{k�����@�w6���L�G]��6���ѫY��$���p:�ܠ���M�]dJ�SZ�u�.�㓭[�X|_![I0u�+n��:�Qnl�c;4j�-��I��3y���+ed߹�v�����I��Wr�V�%�v�Nڲ����GbN���+sH��8v��@�*]�Z*R�H��EnV�
v��u���IK��B�:M����ks��u�����"�u3k1��Ofk��+'U�My���N��1��0��ۛ\.G�#�q]4�h2�"��܎�u���O�(�l�Ŕ,u�J�P*�.�X���d��VH���Hǌ�AŮ�̿�!0fk�!�)�Pj�����T4�6r˼���:��j�����\ko�ܮ4�f��34`y*xb3�ک]���fh�i;념�ủ�&3o/���d���V)k*�;L��ɬ�l}��be0�e�x*jSa����Th��x�Y^񱎆Pt_�e��J�%\��o�j��ʱьǱ���Q�>�Cb�#�i
= ���nݪփָ6~}�[�]ڎ�A�_d��Am��s�I�[���Җ��)J��n��La��VY\y�X�����.V�R�v��*fӏ&�w7d{�u�讞�Cz�5>� �]) �+���/w��]� �v^f,U��0f$Ƥ���DQ�J�}��e�F�
O+nc���Ńb�
m�uʝ*ޓxq��C�u^_9��rD#��Ѿx.�+�B\�� G>W�b���q�ѤA%<���vS4a���<���4��ҫ^º*�-/�����VnŊ�U'{ �<b�.�1K*-�,�����9Y�f2�cc%���"��2ev�S|�H�� :�������GN�Y�����R3��Ɛ	�_1�����f�Iw���Re�\N�ubn3vj=�AM��h��O2�j�I�L�S��I�%�h���*^}ܺ��v%��jtZz��LHRGs/4e�;}��"7JwoM��q����
ݫ��|nlr�N��}b��� Nev!w�%J���!�`�m*�r�%�[�I��������J�@�}�LP�f�|26��A�{��ɵ۵r���ـYM,u �i+��s+8����L�Z�<�j��l16���c�ULR_˙�F��MS����:�W�Kh-+8��8Y��gp�#���p�O�Tz{�<�%�h���v�b�uu����WcZ�oq#t�c��T�P���5Ϡ]�h{�LLL]?���+۞�x dg@�A/�]yG������<�Q7���-��g���7����rtq|Ž��ԍ;�����]�|�a��7*�o���/%4�oML�b�ڙ�]C���.���:�������ذ_*]BI��`�6���[
D��6։�Հ�՝���ȝ	אQ�RY����p�QL?fA��biuk}s�n�S\$S�l�7��V�S𺍻T�q�yRQ�':���UL%�9���`�	r�ێSv�z()�������]w	`�q�����9�4J�T��U��w�44�kU�Z���\RV,`i�j������ޱ����Y,���T>:�Q땄u�k;,�%%>x����Vdu�K��N�	�������n��/�Ѫ�;r��~U6�z��y��E-�[רgi�՘Q�_eJDPf��i�OZ��5��G,A��Vi��m]_Pʁd�]����R�7��'u0�usE48�P\Sa�x!�EgE���,u��]��-�U5���5p�Ĩ�����P�����z
��ñ�v�/��7wg:��3��j�ۇ9gs��"&��������I�[�)wn�2�n�ɸ��:y��hC�}����x*J�S�әQ�/&M,��Ŏ�4������]q�)��}+��}�q�ǯ�R������Y�FN�F��C�յ��)Y�K0Uέ�V���ϠB��}96�O���}N��3:<�:p��4�����	�vs��y�u�B1ʻ�A0X��!�c&�Xute�mt���m�{w�tY��%\�-�h\OE#��X�.�����M�|�-��%4�K5z�K��1nC�fb��S�O�.Ĩ�_e���S�җ\i��;$u�s@A��0�lVJ��I��=s�2��ظc�ѡ�(o�o'y{هP��T��S����IK���+����&B�pg�x��.���r罁�5č���}�j�;��F���G4�ȴ�����h�;����.�q�:@i��=��n7n�r����dޛ�]�Eq�哦�XG���iV�z��kB�kvMc�GG�3���!�|6��gK.���&��yĶ��/��t[N<��=ki���x���ƪT��<c��{��)�);�T�2^���:tQZqp�uja��i�u�0i�Q�o7��{|��.hr�]�O':��Α
`��Ń)DOf��8)�V�5�՗�euty��"Ko�d��\'ut��Sմ3�;gyv��Я.֡��'c ��v�B1$�Y�e>�f�+��ݵ��Wn�����0���
͗�-��8�MiA-�u��N�6�]IOx��,���t3��sͺiM��|�!/T�����A�����!���j�G�1.��9�g3��L+	=v��mԸ�3�M������`�~�;�iUσ�
�󼨄����]�ER\�ܱq�:>�
Ȓ.�n�����#��j�w��q0k��93k)qՁ�&�[�w��������wO��7�v	U�N5}���a��G�Z�[�G�b�qj�ù0�2��k'$����vBK�Q�f��V�+�BX�"�''n�}�G;bW�U�����ơ9�[Y�lrK����U:�/�*����rܽ�it�B�����.hGn��px8��wkp`Ҿ��vu^kt�ø���E�sz��&G
/%���rr�i��h��%c���6̵X���m�B���r���_I���h��.e9�ɐ�w����@!l]��K��y��%˕�h/ 6�z:���׎�u��,낸�*�kd��fͻ�������W�Ӭ�V O�$�E�Tྛ�u83���G����&���kI����~i4%)�r�d�c���`�m%V��t��
<�; Jfs��s:T����8�q��p��qa=Ϸ��'�׫y�k�t�;{�w`����ľ+h��z�r��}ө]�Ν�_W�}�}U�}U����}�D_��}G���w{�R�'���þ���Yܮ9*�^@���xڠs^r��a%r�0>�upwr[�2�㲢[�;EP������Tl1`ݮ��+w[�\kw3��l�m��l�M>W�D�O��`��1��<z�l��x���%J8CYt���(�
gs+r�J�3�M8�-�k��ȸ����c��+���q�����^���:#/�h�[�si���X��n�^�J�y�6=���t^*�&���w,���3��}�V�$JR}v���­U������
���o�$f˨Ը��ݣʆ�1��C4��[���:\Ev�m����}ή�t2��+lw4�]��I��)u�����׃���^}>�� �*p��7j>�-5�ے�<�ʺ�&���$�
Ք�Hv�N�ق|��=G��2�\U0��$�6��g,�ջ^B�=wAu�-�޶��k$v��J/�+
�m��wy��HA�c��|�VH�Ճ>AmJ�	�C�V3$fU��'�G_�R/u�k�E=q�Hqmj.7Ʊ��!GX����H���بۨ!9Fr=�*ێvW<�7�oxɕ����HIڋ��0!,!���ҬX���t�͟wL]��mŴD�Z+��NHp�d�XF�]]p{lVζ��9�u2s{�E�,v]p�o[�E޸�g���7�u�z8TDs4�y�>�����\M�6�@,f��/1���R?=�=��d�l�ѵ9��A�j�vϙ���{e���������i�Ո�b����m��|YVnf�����:���Ҵc�PV�K���5Иv�j�7Rff[�I!��L�U�ʂj��1;o�	�e����K�m��Ih�#�ܜk N�L�:U��X6\n��R��M�\|��t�۬J��Қ�m�		�����ۥ\3��s�y�G�+
�暝���Ls}�+�!��u��!P�5����$阻��d�0�e�q�����u�;�c�W][��ibuC�+:w��&���f;�w�Z��DR��oCC0�]V�:T�f��R���;6�`�\� BbaU�Z�ˀ m�"��V�<�z6�>�G7iJ�,K�_I,,Z����6z���>I_:r/��5�PPH�N���"U��Z�U��h�T���Ɠw��H�8��D�"9�m�<"����ܚYǵڢ����#��Z�T�oD�9�Smr�7�9��Y�pV�(���u�����G���9�Wc�}6���cxY]Z9�nD���ۛO^T���e	��q�%7U�~S���$���X��=[��©6�C]���M:��6��F����:��7#�����5ϫ�Р��O~�7N���n�̉������5��''��/���3����V�Kq�D�_ �q���xE^c�ú2�қ�WۗEwB��A��][qD�U�Nܽ�X;WQ9%�VʅYm���.,մ�iNU}X�M�B���HV�g"�pK���n�c��[�oh���S�ӧ�����Jڛz�t�eN�`�d�R^��-ncO�_�ϻ����q!�E^=�-�7z�t��(rv����1R�����w,6�Vݛ�Ĳ��V��+y�-�9��p'�^�pq�f���C)�J;}�U�g/2�����##���]o[�62��v�ӎ�07�s��b�']�gd�8�H]r��=Â7�>m�Mڍ�K��˘�z�̦��2�8rk��a[�aK�#���=OD!����H�S���+8��f��	�Vlvᆸ���]J����8�<�D��	�\q���]���hwD>��1��}�]r�3 }�)m�yGj��-�u{�����PKӻBoLyt�@f�[�Z&�xR��0�G�F��]4B`J�M��I��,��Y\����y��ām�8����k�'�u#RX����M��^Lb�S7�H�:ڙ�+l�U�-�S���^ިjbJ�9k���������߸��)֐s��� �jʡ�+T��H���{�����v3헍���m��8��͌ޗ�L[J�՜�s�E��e_�ή!�o�h
<�(��3�Dȥ�M�"�����à����#ڄT`�8��*'�l�j��Z{� �uy�����C��7��cB�*uб��nl)�1V^�PNr��h,����ݦ���6c���1�f��j��9�:��r8$
����D�E}��$�-Q����"��e�; DSq���E������X0ٛP��h�4U��`��1�O��"��x��v!+�,m@ش�c��B�d���5j����:$�����jSD��)f"�k�k�Z�^G�ow�9L]��_S�*=���9+� �JLw)�O���)�T7"�Y.J����o\<��S	�۠iXzb;���J{Sp7�/����-Z�VPp��X:����(S{cXI��v�W���V���I�z�K戆����#��&�_98WU�]������<�-�����[��J�WsK�U��xk�xa˺�,Zv�`T���Ȱ ��~;��Z]3�j�����c�p��6��]D(���ttt��o�Y�6n$6��V:L�W�R��9��i�PAN���B�ᘆ;�Ɯw�gϜ8ɣ�et<�v����Sޝmu�#�h6�:m��7��{�Ѿ�'!g�0Ky�W�iMns{���>�ra�u_-�M�	�n��Z/�2�U��r���N��o����kFՃ��7RF��r�;�8f>ާ{�K��mJ7�)�^�P�\���F�!	1Ө�I)���uX��:��b�ʢ]v�μ�����SMc�4,: dm��|#��ڔZ��`���Z�ٱ��M,��d]]�bwo�oH��r��!�h�p��{
��"_�N�}�n#u�[
j��y#Q���Z�7���:@.}�k�9��7�gV۸!��)i�Ϊ����jj�v�4 ��l��n=��˹L}a��*#Skft�mƍ�`Z�2au�u�x��f\=X�l+�WQaẝ�%�pI�TU7lo%��x�3�ʰ�X]Z$�h��S� ^��`	jx� UV�����w-=��mgw#W���n�6*j��Z�n��ȍ� �� ��T�y�e�m�;1޵P�j
w>A8���oF�)H<�C�mu�\UD����Wni�1�;�^	-U�մ7���7O�e�ix��Ґ5�0:�	ʳ���A?.B��Plr��C��Κ'%GӍ�{ugJ�b;������o\��<�Mj��J� ,�]�`�IZ�D��z�=�̨���x���������	��˃a4��:�i�E�7�zf&�{;�B��.[��{W�]�t�25�	���р��Jt���䗌L��3�Um2�G��2+H��b�f�[yxil�ι��6���H�@6�1���޴�"�n��%�����)�W�e�7t˷W`؃�3v.�7[��;R�*�	�D�M-������1��y��2�־ɺa��e;
���_#�(������ݡ�k����acs��O]�bj��f�+^M!Z�����h�JKB� 
<��X��Z���r�E�=����5s1f����ud'xL��t�7%�+��f�=t�Տ��2�3��kI^��U)"2�T���ܝ����w�Й��,�r�9=ᳩ��ڎ�\���&'�a��� *fR�@��v����Rq�6�V�+�h�����mŖ%��(��R�.A�0z��"�栀���6���Nˮ�1c�wt�ܝ���&Aj��4K7� 㧺���mN1L������f+7%��ӗv��0W�{�km�����7S�+[:��;� j�ql�U�6�X:���Os�-u�8˥1�6�Rp�tn�a�y]�6cn_gq�Z�^1��\�]F"yzNc���ýY��NTFLe�ƺ��[-w�k�9`�2��:(��Cz�)�n�cg9��Ձ(N�v�n�+�̮�2�>T^]G��c;6���i�l���_- *��Ǳ����o���ڋ�ˋ��E��p�"�g�fb�d�`,Wj�����v����Ò+� $"�b�fa��̫�V��(<T��xf�Ӆ�n�jWwdT� ���P�`۩/k0Wu��5��;�G-�BÒ��])�ോv�;�M�!#��D��f�R"&ٷ����eT�
K�g9m�N���ֺwlO�D����+���ܓ�jL'5!,X���7O:�V��p���VE��_nlh5�I�o)��ܾ�*-y��üf�;�󝒎u)/��;{.S� �$������7�l]����2[w��ȗr��j������q��0�,DZ��P���Ρ����S�"���\c�w���i��#Wb��A�ZŘ����Vab �e:y��}�|cXԬ�)�p�;����EfX��d[��$�W��Je��v����2��j�4�EhƏ�X6��1ӻ�Ip�Á�]�\���-E;^_:��1}uǉ	=a&�Y\n�ʈnP��Y�GtW���"wu�ja4Ř��R������u�\�_oW<4L�:�ll��s�"�X�\�«n�v��;*s�l�����F$�v��3G���R�m�A����E^	�dLz7v���w��t����q8��j�䯛����=���6i������n���sDm�9de�ӏ8٢��0!�����WV�5Ԇ��niu1�9��]�8d�H�=y���u�[������$�������gt��j�F�8������Tm�6��.��f�l�GoE�A����<J�ރ��oGR�s�%;z�=b�`�*�CS�YZ�Gh��W`�iV7J����c���� �n��vQC=F�K�����v�6��_6cL�h:�ڕ���J�{N��|Dɮ���j����g��N[V�ڲ�ӣ�u����tK9R���k)��xy����᝗����]�6��W:�M��NK���Z�i��a0Ł����SY� {��A�R"��X|�!�����8C�a�e72�a�Y�ɗ�;�c�=�кͳ�ki���؉� �E����42�h&�gF����,��
�w`�&�$r�H�4�+���9�wy�eս�ͺ"���Yu���J=h�0� �{3��>}�lʛ�H{0�/S���b�ȝ����|$u{Z�X��ǆE�|��7V+1�%)Z��;R��tS"�
K���u��P�c�rS�|І�u�Ї����椸���0�E,�X��e$���<oWi�C
�:�	R�$�L�v2�nVb���W�u��B8/(�b��Fw����xtKm�J_fV�p"]d�Va�����S�h�P�A���#nb�ci*ۓ*�Z��;1�1e�ݐe��R��y���x��;t9#u��k����Ϲ4�f��59\�]B$97�n�٢oc�^�ύj4����
����lU@�Ի���3��
46$�ܸ��	��d�7�d��:֒ ����ye�"`Ό��5���b�cpɌ�Up!CJ1`��"���	�ָ%�Fm\c8d`	�s�-9)�9ɭ6{�������v]��g�̌��D�y�[.�Xqmܦ�y���ɶ\<HR��7�>/E��0��}5M�b������"�Y��r�*V��}�vQg�pp8�:����5N4�j���R��ޭZn�,�uF7��+�>�u�2u�M�Z�����l�N��݆��Q��}Q\w����a�H�w.���]MЛ�g沺��v���E'˱��@e�]w�o�٤WM��=�}�<�cqF��16@¥J��V�Z�N�����������os���s�7��o��R�-Q0KT
k6�Gq���Ͳ�%�;V�]��;���s�8켠@ܣ����wI�r��qCӐ�CZ#;ka�hK�ݫ�DPB�;����f��9����oe,�a��/'\�h�]r�mM6�:�B�0�f�;�>��s�[`ukyh�gnM?w]�a�M,��Ҁsp�-9)`�J��!&�|�2eͮ�Sd:$���7[;��r�+�92�uu�c-M���5X��sUj;w٭5O:��Y�����kBSn��7�ll4C.ʄI��g1x��ͻ]�O�o&�Z�aST����u6P�7w\�R��>�XӲ\��i�oq�p�o�7*�X���m.�!����̊-w!��l�L��Ҙv踫#u-�\�"��J+��3@�ٷ�d&�Wk�����Ի�w6�a��o5f��t�'ú����onoE��\�K(dI��@!,%����h�V�F�
�_*J^0��۶c���y"��l����z�f�6��	it�s�CKx��{pZ:n����\���GG��Uպ�mK�7.iR{H��5S(��7b{j9�;��bݭ@K 0:��-�2>qq�7��m;�@�6d���<��R�CF�(�3��� 54��mZ7�7�Θ�+W�0G��>�-��-��O��	hH���ۇ��x�l��Ln�ܭ�P�G��:8���:���q+�'��]w����5�۴1'}�5��;��;"�%e�;Y.:	7��N(�9����^�m�!dda�ClڇF��c�5��)�+uTq�)�3$Hta'�J�XFR�*ze��&� �r�,�^P�gv+"�"��2�0SUٹt�/u���s]W[Ѭ�2�=ݔ�l=Q>�j��?;�K�n�k]n�%/�}��î�Ԇ��s�򚮊,m��De�恰!�����R1����O(P�j�%-��:�1�Xb�5>���W����T��o�P�ܗ��6�uq�<�e@"��o/�����-�;�#g�pX��ab��y�G�Fk;­��8fr�
�-l���晽�0��6����ѷ��U�Pp�̊v]o�敕 ��nN�1}�z�¯��V�y��=w���������+��5+x�y]D˩�Y�W�Ի����_�.�C@Z�_k�U�S9<�����z�^�P�.�a�b�ʛ�����)��@�$_vv]d�S2�}M�v	6zP��F���$��sWb"�]��:��U����R��V���WֲS�Vi�lށ@:�[.m��X��ps��pC\�U��T���;���mVb�3:u�%����%miwr�b�]���?�>��-�;z�`5�)X�����1WD�1�3�-���k�Tf�/a')PQ��T'y�d��6禋;�Rñ3MU�Z�b:ykZ���j�@�N�o���Ղ��N�(]Ej=seh8���u_u]��L�Xъڈ	G~v���N.^�yXw�&2{{����ue�1�(��eF�t"���!ԡ�y��p�΍�Mc�5����̬y$E8,�KfK��yV���"+N�G��U�=Ig{�� �6��`�_49�j��֩չmAkd�Z��tK��u�2�ދ�Um���u���:�*�k��=Sr�c�\����xME���z\�Y9P:=��'H�$�x��u�%íZ��&�2�b�&��գ�����\|���K����ok7�g��� �d�]���%����N�޾�2[�#��� ��hC�]qj�s7��Yi8����j�a��U�7��tM*����ʺ�܍>��TTDQ��U�t��32��]�a�b���S��/:���\ܶ7wr�7f�'��EF�;1�:�1nr��3��wtn��k�����W53I�+�����˖����6ǌ��EW.W5��Nb�ww.hs��F�5r�Θ�ɭ�wut���r$�ί&��F��îӸᱱ��W9n��E�E���:��^K����5E���.�ʻ��m���^y�(��G�v����ɢ�ws���p�]׊��!��˥��/^*Lrط.���#s\�A@|�}@Uu�]^�ct��w���N^�6XK�w�"��ٓx��i�Wt��;qU�n�}�h==M���9��}�:v*�;N��mW��7��-�C�ʡV.���t���m90Y��Kѭ�����gT�_��&���R�y�xW,sP��6Y�m��Z��cH�={T�m��[���gL>1�J�mNe����t�q���n�e롲[뭻b��?j��z���0k2�o��Y4�d���D�/��}Z���V���%g�Q�3&��d�c�d�����u�x�#�%���ꜭD>�VL�-ݦE�Y3���g>nhof��b�8��v�K���s��{���{Ք�ۧC���tP�P00&;�"��i��ކ���p��	�'�6F��X����t�k��b���@K�C�p*����چ>�@�S�M8�LB.�U��|���\d0D�2�^w!��P�p���	��&}ja#��K��5�.�J�~�珯;Ʋ��C��B����N��CG���WE��	1�Z�����i���l5+�n
��L�=��K��]��5%�. `�2���@2x梓�%��-&�ym5�ܼ}a��:����E��̌�)��\�9̖:�uܷ��GΖ�j
U&i�#�Y�|�x����'���-&�
�����_mΧ� �8[ѨoQ��Y��9�&��v���L���J���|�C��O.I���vl��*�{���2�5�D׭V._���X�qPԝ=pp}r�B�ʖmA�el-P:���Is	#�F0b��|�"{h�R��B�c:��o�<nQ��r_H"�2��cNzT���DU@��&4;�j;n B�I�A���f02N�sU3�Għ&U�r�����<�6�)�#D�8H�}G(�;��6;4T+J���2�|���Tj���7�f`���46c ����7
�O�F������b��3�oJӻ,�+��9ʕ��7������*�*9�dɶ�͉������ua�N>�W�����/h���p��}�"ְS�Z{���'v"��̖ˀsa���S�iA�j�y�t7ݹd��ޝZ�<��Z�
�+?�(���A��:^�br?��0v۸�I�]#8*�U�޹oY�v��-NWPJ��u���vcn������T11X��*lJ�9��4#�vʼ׀��)�����|ڼ�39i;�EWag��TZ��g���*�U3��3��׀1thm:y���-�[�	{���yz���^�E��I�w��,վ�(�T�)=ȕ����j_|*�q%Ι��-r\6���W!�:�0C�Ċ)��{�{7^�z��%�RO+:d҃��C�Q�BQ2��J��y�C_S\��]W��ĺ>�����Ws2�jy�{T��"�� %�TO@�k^K�*��P����e򷊩*�K�^�� 8Z�qGi��!��{κ��,Cn8F�@u�d��D��ۻ#�7��e��k�.�r@��L!ю`oLS7�eg�����I��m�A��	�M�}�{#���s��F�nt8���*̈]5�_�C�3>s���W���~���%�Lss�:�3�
����_�I~* ���`�iW��fxsϖ,�B�K9�h�YۈsiK� ��@s�l��3��ʧ��g<n��9[@w ,�wi}�/c����n_N�)M;��7Y��\R�	��D]�� eE����  �F)T
�S:�L.+{��z��N����ں�f������㝬�w#��X��R'���讉��0S�G��b�	m���_�������=V�����h�9��2m����):�h\��#�#�bbp�n�ᴛ���ޛ���$h��`�1�����!�Ƥ�}�I�g!��k�j2):@���:(*-R�x��T��cX<�3|8����t�x��~K�,c���җ�&��_W��j���:.�r�N�w��7�:BS���=��6r��_p�&����Mt�/�9-�}�h�3��T���A��f�.���lK�%
��8w��B<�4B�O���c���9���ͨ�q.^�0�Oݮ�c����2�7, �?X�"(GRѐ���WűG����LT���bC~#�����՗g��'�����(�9�G�����b�DX.nZsB)8ʑ��� �|�1W?�^��
�R��Ǐ��O);�8ZU���s0����T!xꘞ���4_��Q#�6c~��3rp+���M��;��%]DNx�/���s;U�vu�ȗ5̀C��Cwv��=�b����D����դ]����֓�ر��H{�py�+�:����yO����㞺Ok��?y�۩3[p��^��{#��;pV;�
��א�цC�� ��̱NS+)�� �g��ej�{{�qj�Sjv��0)����K���s�lp졾���K����3��;�9�8��Ԏ'vA.|���]^E#�f� ���6��O��F)L��-T�֮�����pVvn�W�$酪@�-�R^WϠl�p��:�` ���(�7���:�9�IΒ΂���7��:�v�>�%�z�����j�ҤM.��!K��e^/4zょY��3n��u[��>;�]t��Q����}ǅp��h�ܜ�;�]$�+)�.Y��\�i;\B�ͮS�J3&EOLg��)��0��nK�7GH��*_H�dQ�Z�����+I��p���
 ҉P�tx�ٿf{2J��3b���f;hx��f2	�/N71�+玢v�����|�\z�*�� ���м��ͶR�60k2h\R�C,:�t|�t�	�VY�c&��C4�)L\MIݼZ�w�K�Z0�2z���GG�Ai���A�oY\#��M��[���j�˯+�U��t�����f�~���H��A�^�a�������2)ij��,v��nI��{��h"C�a�{��r�5����͟#݄1o+�2.ɪ#��LR�"��Bׂ�,�y�!:����3B+����R��mCuC/Z�%�뭳�g�j�x�g��g�����#d�Z�o�&W1K�N3�e	�F�Nc��Ɍ�um^9=��Ǳ��yD��Gp|��}���ֲ�uX>�Iֳ����W����P����śgi�x��d��T�f0}�Xʹ�7NX"���y�pK��{!��x��:�''��߈OҶ�`��Z2Ըs�Pm���,zE��v�����]�ep9MK�%�v���fC�޾����Ͳ��]w�3�� H�1#M6�^�g��,�/��W���y��g���S:�fwI�]����+���r]Qǋ�V�9K���cJ��r?�;��9>��J��m��9�y;�C���Q�G�6}斗u��g֭��M����،�L2�G��*?�5�X��8��o��Ƽ.g��&�~s|�'R�\�Wz�j�{���]������	1��W���i+=^��X{��޼̓Ӹ�E��V�Ȇ���ƈc�Y���jи�r �D�&�9�c�b�����[s@��L]L�3q
�}5�)A��]�u�:z�q��b|7*Y��-�	V'�;�8���e0@�1OD�3�Cϥ�|s��y����Y��[
�5m���n{C�����H�AE�J���cC�{j A'���F3���a�9�8���S<"E��u�9�qZdHB��� :���3�����^]�`������{�ݖ�EB%��W����`۾��J�Ϯ렴>t9�Y���p�/�C�Q[��$�Y��ΧGDwd��M�؜z~�'�ua�NA�b+��nm��ƙ�n��w|4���!��݁f[��;C	ٺ��l�P ��J;���k��n{�˹ϫ�f<jnދ��\��4um�1�s��=K��w�ː붰��ާy��L��k{�&�'Z�����檼�c�on�:�\���')ʷ��R�_�m�^�Z��Q��i��[�:���dS�?2[.͏���t4�< uv�|��9�;��R��jX�fģh�҆W�(�B���F� ����m�����"s�����Zw���`�(��?t�~��ƂTe �^�B:T�6�>s��fm�f3�����ĵ,��c�����\�p�Tt{�Z�O4*��G�+1�;����`�B�y�˩n�;���Ok�s����b��v�=�qV��)
�h�=z�=��t�&<y�۝#�}�.����2̺��P_�n��j����� B�L�Nz�
-�m���9�OW�ۻ0�dra����WLS-��*j�낆q����g���rE8�m$�ֻ�X��+J8-�Ӗv&+�o�������0��C�*������h�����E�h��ĞtV�����"a�fxsŋ4PRX���Z1=�Γ�<+������ON��P}={u3�5�n���R�)�]W�*:��R�U�>�p!��=���Y7��{��r�\]p]u''��U�hI�̳��=}o"�ϳ�AG�h�ޥA�r�p�I���]��ﷺ1w���aQ�]q�p%]F}'��]F[�j_vj"�4iξVe�&���Ha�j1O�u�ҫ���$F��Q;��e��\mp�95Rwyvr��ol��������'!:�sp� !#�)�@�ud	��fw"ci����Ogrܼ��)U��9���;���u�������7�c�8��!4��z{�"��Z!Z�P{�Lu	u�r�p�-��%dC5�'6�Y�hY���2x�y��Qj=Q%s�+0z�U�
��jǼeM���дi�'e��3���Ȥ�a���]̝���a�ٞ	}΁�4�{]`��y{������.9+�!̶X��f��xi֋����蟨-���z�0���>G�@�C���\��	�����$�����KrYy�xq�P���i��2##K'�X|t��+����+�j�`�P`7 ��r�5=ٍKrdn܁,uLOg�١��$Z>�/������b�FƋ���m�t]�n�e����T�2[;����z�x���ଷЈ#'�LyO��=��&ݽ�{q�/R\���=�\����A�\��Ur+>�b3n���tOUL���������kd}I�)qζ.���KȖ�*c��2��mˠ���v��(��G �bM�xEyӹ�9fk�vо�˟7x�r��R>�G�^�)�z��p��͵8U���܇��w;}�Z���k��n,Wj��c�{�ܸ��EZ�Þ�->4/������J륝��>�b�.C��(zJ�@?�Te��r�YN�5l�cY+�Lӧ���l׾��M?z�Q�iz|��P�� �kw�	�2�]<.�6���!.v5���8.�V�����pX�I�E}F���t��6��p_5��W�W���a�[�^p�Z_��F6� ��ޤ8���|6rJD�H�:����� u/̇�,�G���8n1�9U�l���aq��Ds�R-��<�9�"*�W� j�opT���'�ib/�����b��:�I�)��g�-�oō����%S��:��͖c@������0�@C����򤝠�D9j�0�u�F�@Z8:���e�wљ����gJ�}�$G��&3�:�LN}����!G���<KKiL׶5:twһ����y�X���Uů ��o�ةUՈ4+�
����fz>�W� 9�!��l��i��%�<8I�KȄf��`g:�%@��ߎ͇uպd-.��W8�R=n��~���3,��t���o�j̖�N;�KnA]c�uڤ���vk������2W�sP���-�aԚ���b;
/�I�j̴�7��/�ZbY�NВ]	3�;5��]����l�qq..Z�.�Y�h0��Vu��W2�>կf�NWF�t܄��ޠ��,P�Pˈ�Cfn���YC�G�C߅���Y�o�NW�+���� cX�Ο��ey�]�����O�93L�T��	�q��P!�  W1��Mn�O��'�`릲�Ԣ�r�����å�`��u�������`��v�"b�3�9[N��kb���q���!qBl��,C�W>w˨�{.���^�ʞ�������k[T��8Oh?1uD���
O��C_����]�8�DS�zx��ͧy�L>���WZ��_�=�lL�	0��s�����_P9�B�29c'�&�i{��6�&S&�h�[w	����c����Ӝf���5-P�u���:�S�S槲r�q'Bf�H3ح3�Ie�����C�S��ӂQ䤂-*�wPU��Z��]j�.-�pg�`�sS1��B�_M)A��]�u�:z�q�):�!سo�܉�&�%;��R���[�tg��a �}5��Z(\*]Z8�nwID}:bru���o�f��C�iSz�Z�૖I���w���(�*ևi/1��s��m��׳���ӄ ��w���\�=]Q�W�g�;�U ��i�xh8mGEf�Rf1�gkr�c"���[VEE��뫥�wM�uӧS)!.��,�s��X�A�6�i�5�:��![Mh�����ĭ���rJ@�I@(/(d\�H���N�����7q,�Y͹{m�� O�]09�ǅҺN+3��f�-�荮,tj�����,iR�K�[��'\��6�M)sΊ`EVI��]����TWG54��2��rL�����+kZU�����[Aa����:��v%�(�F�����P��+Y��y��Yy��쫡j\%�hMD�T��&=[�C\Xj �H�
s2^G�z�m�(1�4o���]+�g�
��O,�!Vp�1�\ o�{on��&��YZ�\�j�l��衲�͕�AVF.<�Z�E�q��7F�U�pH;vT�Y�W����X>s ��P�2�����l塔��v�r�z�g%�X7������������ml� �a��5�ԠZ+8�NL82��T�8��3`R�k���O�|�_n���n�h'e�Em<?a��28-;H;Y)3,��cBa���N�a����lͳn9ewa�u(#}�eu�PY<��RgY4���b�.���gk��!n-"�m��,%��u�\�k�Žxճ�]K8w��f�ww��,�@� ���
 0��]D3��4��;������	;-�.�V�EK�m[�t39,b%񱙆�%�X0��*��c�0�'w'�f��Wu�8k�r���t��>�n�5v�F��k�ڄ��Wp�\EWi����ۼ��{�+�tb[:�w�X�ёnU�۩�?�*.�OݎU��-��u@�s�*��k�۲Ҽޘ��oyNv(f�5n����Q��ژ��խ�?✗˓��WQ��V����х�Uͻ�=L�A'zs���x�:�-�D,�l��|��!����q+�d����+�#���Q�B���գLIr�*K�l�,op�]�V�3��P�t�
�ꔥ�/�԰n��y�s�|�Ï��\"���u�P�\h���)vJ���W�Cy)T�'k�P�@�Dw6bbc�Uwe<��)˝�6�Iէ,��L)��� Қ�H��urCm�W����fV�ųe��:��'\LU�l�f��0Xz�wW�^�92��dw2_<.nl���{�n��Y�:������$jZ{�*K%�s�f
����nCy�6�Z�;�\l�5ƴ��7o� Q��6�c�nQa�fjp���p�K�2It�sn�^��v�̆Hh>3I���wҐwY|53H;əJ�8�����
3x�tr�<��GSN���)s����Pިە�S��t�� ;����|��滦<����P{������~��w.�k��ݢ.F�Bp�qH�GwZ��^H���X���\��ۓ�����j�-����J����ܴk��W-�滝;�&�F��P]�m�x���nY6���;r��8�wNN\�8���˺�twr���]�vwI���#���vN�/���#r�\���[�r4�p����7
+����Nk����.�˥ʈ]�*+��#��r�I����;�����7�vk���'�4;�h�s�E���!ݻ��6�W��nss�:�rcL�.r9���N�A`�q�W6�9�A�ΘwnM�w���9�;��;�M&LW;��r�k�θ�r��ҹ��Mx㮮����4��n��P
�j��
��]�����>���2���ԋB�������#��B��0rg2��W��{��Ε'�s�|���%�5M�ա�i��;�{�����-ƿW��5�W�������H��x���^wlno��/r����/�;o_�W��^u���}�~~N�KO��{��~z76�_/w����0|��)�a��n��vDz_��o��ߞy�����/=�>��k��wv����_W�ѽ���v���W�u૜����;W�ֹ���<���-�x����������?{�#� �#�&f�һ[���v��g�ߵ��-?:����Տ��o{��ϫ�6�;}[�w�_���n����*-��\�>�{{�ֹ�W�]�/ž��-?����m������^��^�����}���+�	d�2�����vO���_��_���}�ڼo�������ֹ{Z{����U�o�^�<���^/�x��>����k�����[گ��s{��������}�ڿ�����i8>��DxA����4�Jɭ9w��5iw���ۛx�^�o��j}޼������W{����zo��5������_�F����������z^-��}z؊��W��}��޾�����_��|��^�6�/����m����F"$D����r��ׯg_;褭��B����/J�i�����ס�[r���yu����~�������?[}^
��ݯ��~��y�����Z��ۿ/��~���_�F�|��޻�狖��>�^��D}<b̜C-W����nڇ�>��=u�|�u�~5�{[�x�����}^5��+��~�KA��������x��ץ�����������m�v�W����"�>���y�v>�>b �Ȃ�����AH�U�<��Uo���Ko�}�H��~�*��׍���u������5������W⽭߽o��M�W����~y��h���=�u���������-��[�����x�,�
#�#�"��^����u��k�s�^���*��_}|�������s�ϾnWջ����^���~�����_���5�om�ۚ�����^�ݷ��m��u�߭�ſU߽�W��oǍ�yצ�/kF�oK��צ�"G��xOla53]��֯R.�|�~+��Ϟj��77��|�*�Ϳ���|�~�|b"G_�} |Y��LB�����}���o������ϋ��6��w�~yW�����^��[����U�����+�G�iK�t'���u�4n�9��� �!}c`�9�����V�i��+�Һb��ӕn�a�J��ԟ
T:��l�����\��buAԩT�ɽ�o�	�ή}ʫ5A�K�m�cys�"PW� �А�m%�4����i�l�]L��z{�*�P��}|��B&O�hb(G���|m�n.o~~�����[��~��^֝ڽ�z�ܾ����������^���׋�����/Ţ����盟�+Ưw�M3D|���>��t^t�l��;~�������}��\ۛ������o��x����H}��W����¾��}�ت������~z�����5����oϝh���Sf������u��͉'��
���}�oֿ�E���+�^-�\�wη��o���^��ޕ�5�z��/���*��~k�^�����{�ޕ�_�|>�a����"",A�w5�����#��z~�"�~���Gƣk}���Q�N�����żoo�_u����u�o�x�����o��h�_������צ��[󺊈���^w����7/W���oj�r������m������k�ѿͻ���V�]V�}W��ǥ[��A������H����ۚ��כ�{_�����ϽzU���o������k��+�����5�y�szo�z�z�>�J��μnm��s����r���ϝ^֝��wW��}jDp��+��W/�D�{�Ufn�~B4o��׋�����}_�E~o�����ƾ+��|���W,}_y��*�^��y�߿|���W����7��5��rޗ���>u�~��{m�x����~y�x�ۇм���g�ѫM�Nb[��Ѽ���>�k�����_�⿖����ڼo��o��y\�Z7��|����_�_��^z[�\��r��U��[�^>/�y�j�˚��}�{_���U�w������#�>��*���8�߶ŕ}��̏-/���~+Ż��+�ݾ/m�ە{����m��ޛs�ݷ��ݷ�x����ž7׋�ʢ.L}|�}��H�,}B$G��0�����η�������y����i��"�߼�=;�+�L����[�\��;_�鿽��v����zZ7�����[�^-=����6�7�no��k�����x��4U�s����/kE������6����\�.����wm��z[��(���gm,�{�,z"��>����1��祣W���i���i�^��yom�Ƽ_�{����h��O:�-��Z/�믫z~��������W,}_�8ň�b�G���u���A{���\<x�^͒ўJ�U��p�<�s�;�H�^���������j�zN�{]�[��jsYbE��W��yA�I�U�-�����V\f�q9P�޼y����IL��J-�+�Ss�a\-����B�͡(�=ݛom9�Qch�]�;�=�a\���|�w5��������Ǟ�����.om�}[�����~���{m�{���?z�צ�k���ž���k�wy�ֹ����_�ο��/kF�������ֿ��ߛ�o }"��D�=�ET�f.�y������oj�}�����m���s_��=z�/���*��|����[����?~���{Wջ�/�~�m�ۖ�|����ͽ77�_���J����ou皼[�<W��_���c�#�>�N곳=x��}��9` �ѭ��j���k�x׍��_o��*�6"�{����W���m�z�����ϫx��~޻;�7�����o�|���Z����~�����w�.������w��*�^�H��>�T/a��`)��{ޫ���^�?�}����x�������p�1���O� �P��鏨}��ğ����H\�{�������z�Zw_���*����^/��^�y��Z7��/���7��-������Ȟ^^Ҝ����6�����nzk�o�v�ήX��/w��J�.oƽ�^z��m⯋����z�j7���so�?�ߝ��zom�}[��w��ţsn{���^���׍}k�����zG�G�H�c�{��]��]Q��~���|�ֹ���]����Ţ���|���~7����~ߝ��\����b��[�^z����m�W���x׋��������\�;o?�^���W��g~=�������#��{�#^s1'o}�vg}B���>#�y���Ag}���j-���?=|�_���ֹ���s^7��o���k��^7��yޖ�b"������k���>-�^����3��Ww�Mn����..�Z겱%۹�B(G� ڟ��c�#�Ƽ󯍼����|�����o��������گ�������_�Qo����z~����ھ<nm��>/K�^����wP�!G� ��3�ux��Y��V��X">�1#�3Ah�>���T|�bѽ�����Z�-��U��|��7չ��y���կ^ur�����ͽ������������o|�}�����빨�|�D�#b/:��3젺vt�zV��������/�}֍�{��m�������|_��~��o������� ^�a�zcEC�Q;n�١1�E
H{�[�k-w>.����=(=��ʹ�4�p7��>���	^{��غm�z���}s/���s�TT�2v	�^H�=�m�Y�����z��LRJ�]rtpZ-+%_Ui�*�s^�,��j�D�R�����۔�<8�jP�$=]W�+7y����wF��I
�� ��BQ�/AC��Gʢv�󖬳�1��$�Pz��ECeGU���C�6�*�T�I�HK�O
���_���N�M��7�����;�3������[�*��h��Q�*�?�ܭ���0�t�G���ׂu���V�+�!اG�'�������aA�*����,�ȎuJ��}��~�b�;Yʻ��s��,�W��q����+��w�W�%� ��n�e롳7f��P��ȿ�^�&'����o�^�������GO�Rey��ޢ��>���4�5��W�fO3ڢS����q�3���5�����,g�s��l�+\0��`��u�湡���zeB�1iը��c���u�0P~*�*�x7i῟/��L���ϝ��Z��K,�=��1�j��nﻏ�	��?t��V�=��m�41<el� ��FB��kzsw;/_L��K��ۦ!\��s���ƶ�r�� }�P�~8+�T�޲�%@��i�m��6�v���VN;�Ɇ�Q&V�l�� �Z�uctY�34�:�����uג۱E<��{���6orÊIB�bԳ�ccs%g��O��h��-�^�f�X�����+	���F�B�Ģ��jR����niyd�6']PR�6�6�/f�O�i�Ү��W�w{�������/���@�L��;L��T�F\���Yr�����^��q�^�ݹ�w~�<�+u��������W��s椲�ƈc9�p�F�|6tJ5���B0�~e�,euU�*� ����sS1̪S�����]�u�:z�b��Tdp4�S����[�s��56xv5�Qs* �� #�z'��Z(\*]\B8��y��c���c(mW_U����*����΢ 5R�&�&4;�0��n C1v�A��12$܄�vzK�{�)W�;@{��w�y����d���C��K���d���][YKZ���f
�p�C&��\�kC!'v���V:��B�Gg��[h��p'��ok��/�
u-�q���b~�]DT%)�&�7@s�f�?Pά:���b�-F�5}�㮋Uu꽷g�`�{��ʇ�/�u�]>��d�㟙5ˀv��t4V ��[�3j�nR�6/L�2K� tY�܁1���d�/
�c�Z�o�T��R��7b�46\hq(I��W���n�*�����,�*��r�
���'��U�"*0_'ۆW�J��:�{R���t�L!��
���ةg)*AރS�M~�@ܭ}]DqWo.�6�o�x.*`��9�����F�j�ξjXĶU��_N]M?"/�����a�I�y�oH��`ۄ�(T'yt�}œ���ρ�0��`9YH1Q{u\�6H��N�Ŧ��f�p�w)��4 �Ƴ��զҩ���\�g�Z�<tʠ�4��{yW���ڌ -ͮ]T0.
c����G<��+h����.&R��ړ�+EE�h��OH9\�Aш�#����s,�S��W�|c5��;���"�ON)���c+S��'���m)[�TqW����:����ܦVSW�_��uaZ�>���T�u�t<���{Z-_27 ��2_)K&�+鏭�t�3���K&xL�s4�-�玎��eֳ����#Ĕ�pℓdL�yh�j����ml�h�W�uڼ���a�Ԟ;p�8)Ө|;jQ��r������_)R~�,z����SM���N7;#�����s���rFqOf�sA	Nf\�  �F�)T��)⛽�{};׍Kl�ú��f��_֥�G"Έh㝬��ք�[�I�O�h�Y&��1�4��AQU�M���fX?\��i�p`I�Z����b�c�ׂ3��tY����meͲ��K�NH��EhR*����6�c���>���ћ!6�:��f�[�
w��{��݁�\z�_l��J�Y��}���uus�b��e�oWN��a]�4v��|hf�
���8�c��q����*!:�hK"� ǭ�h.��z_ ]�/�å�^1�a��z�Aq�1��vY�s1�+3']�V����m������	P�w*��3�T�R=�����'B���?�o{�6�g���@Z��rU���d�q�3?e����<lm�t��|�=����3֯�zn"�m��В�q��a�ώ�\ct�ć9;�Ўqs"42w���1���>����#>ng���ǽ�l�P���W���>�!a���\}����{x+��F\t�p���w'�߂��^����G-{�`hw����U��J��@�,c<�W�Ѯ���b��޵IC���l�.�И�9'� 3�Vt"�Β�p]|�EgW �\	�<*�q�9��l���L��<d�e��N�5:'����`Δ.)�(�{~4dW TB��X���s!�)�f�cݮ]�}�q�WS�7��n����_QQ�iz�
�ŗ�x�C�������|�::�QhSFa{w5�g=ΰ��e����qN27������$�:3���p���ŵ.E�
�*��$�D�ٶ���|�aκ����HA!k�[�q���Һ��̱���9�*{�����g;��\*���uܖ��2=�{�xk4��@���z�v�U��6&ˇ��ʎ�v�}�Ŵ�F��`���]�s�Wq����ӟ��dޝ��Ͼ�~�z���}%��� ��Cޤ8������� S_I�*�uȠ�-4�t�]t>c��QFBf���q@��u)�}$GT<w#.բ��>��"S}�o���I�ǯO�$�GA�1�����c�>t�Niz[1��:�ؕS�zv�9�����G^�UT�P �߁d{4.�����򤝠�|�,�>5
�M��\�*xD�ly��vZ����gg-s���z��oQ	`����.z2.i�}}�o4R?.��R��Q�',}�n��o���Ո?�
�Ï�Y�7��[�Z�f��C�̽�UɸW��Kϑ�p\a�1Ρ�P>|t��{b��Sr>M�������!�+ʏL=�U��S���,_7T2�5�ٛ��1+��;�{Mn����A?�Oܨ�#�X7�|����5��z��O�����!� W��M9�p�1��:�{wN���	������{�؋�� V������x�����[6��l�:|�õ��aG�U��X���n�J4����V�i@���z$�C0as�m���Sv�:���b��c��:�{g\�z�k�YĎ�5Z��*����ﾏ�K��m��Bp��!�6�N3�J�'.;iW�d1�.����f���xY+s��j�3�8n���xg
��&>(TU�a�X", 6�h#YѴޠ�S����k3�;��ud�J��=��}�n9�p����F���b�`i�;J@|dD�tm����O�w�g8�.Ww^����N����t�+�]p���_���˘ ���~ҷ���N�uyK;�=��+ɸ�/����agÝ2lh�[w	�-K�+o���]F.�OV�r�qk�=��o��~�p�ߎeˣ��9 ���2�椲����Cjዣ�<}�d~����5���T|oV}܈!�/�P��]4�x�u��?�Pc<t��'�
V!5u�b�T�fv��������R����� N �\ g�t8WL���.���DZv���[�v��Mۮ�n1����R��9��[$�J��#C�0��*�O|W��y^��c����ٸ�=|4a�0���h��U��!
�0�D�����Uc�̬�g�­@٥ڝ
{ڮ�����O�ne܊�5�E��~5��JA ��ަ+�{�Kѯvyɧ���������Qo����@�3Wvk��UsR�4�nҸ܍��Y�	�BgZ#$�1n<8"���Fj�Pr=BʼOu��NQ���~Bc�EC��-��Zf�0E��`���UX�b����5ϊ]jᷘ\���	����<���~3�{��2Sr�ց��$�������f�r�,wXx�z�F�
t4XT���{�aXv;�.'U&c��5ˀv�b�dʷ+��+��op{��-�T4�(@���	�
�<8*��1q�&�wEL�p��}�i��HR���~�q�%1���'qB����9Y;~�A\ѯhW�,Hz�}r�V�� �����s���A�����S��W��7�˼�W%i�3]��_"̻��W���	�F��]��z�+�w�E�hd��`YA�}9�{\"��p�y[F�l^}2��O��q�����T����9��O��t�W�z���	��s��~�0����!X�m
T!���@D62E�sR|��¼�UVL�"}��ra���}ҁeѶ�2��_���!����utŹ�|tg���2�#�+��J8>��dЅt���:cDtR���bhr����F������l������K�}�G/�܅�g��> J[Z����].fgwS�!�x�u��<����.��v-�V}x,���ĉ��#�St�����gAԕ�ʞ��
�Z���C��NY�'�_>$�Kr�M7�9��JM`z�6��1�ޕ;���
�5؀4�}�˳/D�J�I*�%j�k���YV@����w��c�����[�+E.f_���%�Z�������-9�T�t�t��z���W1aC]|�B�ߢ����yG)�<�M��ɯ��b-=T\��4�k��>#T���|I�ڼ��6�[�n� �}v�F7&r���H���4�/5��V���ٰ:�����g;�c:�Z�������ݾֳ�"��n���fmϮ<,�"�����N�,U;=*�'�w֠��+Aͮ�j3�c첺�i�K�۴�@0e�k2L�.q�݉��q5�ӥ6�n�ާJ���Aݦ�!��Fwc��]�K9�l����q1�զ�Y�k�:�V�3�FA�ۄ䣱r��Sv*aņ��;Gl5�t*�c!4\t�L^�V!P���%���ͺ����v'Ԣ��x@5b�ЄMzތv��S.���z<)=�Y���G�j��OK� 啳�Wu���b�^�h��	�o����ܢ�.�n��h��S���Z��m�4�u}���`����X�@]���G,R.bj�ތ;Å��\�C[@яz*S�N�O*G���k��uY'!�V	E��a��MWx�XH4�2R �R��\z6��~�Y�+άp��@s��ͨҐ�U�b=��	]2|��7��. ���	����N��M��$������� ��;��U^*��o��GaN�]���*%<kN�]�.�԰@*����d���$~�nV��C�ҌXˬBP�y�9�D-AլǷ�f�n���q+��-��E�%�Һ��|Մ����Plu�m�-�,� I��(lHaV�f�*�C�g	{�*��F3hʽ�8�f��;�����*{�b�l��5�wav9�z+�0c{��Q�䫫XY�xB���j]�m�pL�x�Պ�K�Ĳ��Q�X9GD����y��6��E�o�n�
�� On��}�,��[����1e>��]�d0a��mc�����匭���9c����씛�w���ϭU�ّ����9�{���0X@����*u�Cdb��c��*uwE�Z��>� �ӋQ�Ǿ��ia���Dv5���D������٦��MAE�L�{b	#ʖ�X8p�c�*pS�p��.޳Dڗ�gP،,�h'n]YHd�{3-���uk���+�^Xp!�Q��{A���ܘb�41���y�K�N���ǳ�g�InQ�u�֜�+�����o��&I����
��\+��2�M�s{��,`	�!J�Z.�nS�H�(�|����Z��!ޗՍ�������;G�zT��v�P�pwDȈ�.y�r����WX�Ns���ɣ$E.�x�9p����R�du�5��p5��ݸf[����8�;��·;�+�+�ع�gx�<A�.p�wtk���(��qݸs�9s�.]%�ƍb�n��Y'wJ��'7H�1r����Ӌ�ۺw���ph�7�fW�r�`��F)����d��I���;#���9E�u݃x�QF������wlF�]4�+�t�wc\���������!��(��l�;��y���-ʍ�n��n:�wqy�Sλ��+������ww8i�۝cb9�tD�˔Z]�2�.ng]���\Ѵ\�s\���u���������9]
I����.��i0��vv�T*�
*�gp.�t�yӍ�����K_R��Yp3��L}8��Mgu�`j�ө�K��݇)�wN�V�i�ڄ���h�_�">�17��s�����_��ݸ�q��(G�*�3�O��x"k�$��ϻ;400?{U��,т�l���ռ%8�f-�u��l�v�@�F>�f6�R�)J�e�Q��&��&��;�9R�r�[o�v!�#Q��eC�Js2�Q y;r*�����ߵtcӌYW�9ǫ>�-r�d���Ý��r:��X�F	(��q��)9V�q�5QuK$�<"�K��`/��aW�u�r�p�.�2V|�hJ�����ļ�O�f��,z�7D>H�K�����A��3]�D+��Ԙ����^�R�
�"uP�S+��e����q��u9� N��zPK���Mv��x�Ab��~?z���@[���V]Dt�S�ͭ2��i3I� ;��k���,��s���%�a�(C�߫S�m��H�R<%9��"��2���'t�y[3(9ٶ�Ts��QY=P����B�X��7,���ԇ+yFD`�0�5����'@C�X�����p��2��1{�rwq`���v�#��
�9�Ƕ�-���Q)}Fk�Q�ӳ��6B��֮�])��r��T�6���h�8��U�%�g�_6@����4��K����W,mi��i�B��:�QB�������]*�+���`���1�""#蕏�t�(V�����YU�G2p�鈬}P�T�2Ic��r�����,t�pX��r��]^�!h�0�y'\����62)H}7e�v���c��Ý
�fe�0�y;��U��4׫yhP�
�R2�]��|�����8����t ��McH�2	�]I>{��w�qґYN�5�VCO��n�@TT~�QQ𶗡��
��I0�7\eLs�hv��}=��C�0�_�i�N�|o�Y\�$�A����yp��u��_�K��sFp�詜����Z����Y����M�ޤ;"%����IW
@�#5�v�pB�i��"��H���Q�[9�U��{�S.9�>�#���c��P�s�e��sIRY��V$CpB.�d��U��g�Bӱ��Cr� ^��s#z�I��
gp���	��]pW=���/�kǨSAU=��|��.C���jN�C��&�p��7s��/u����f�I��+�6�*�Tב��DwQ��}H��-��I��몥��d�w�K6�M�uz9�%��Fw�U�
�_�#�I��d4n�7x檷-�}w����T7�n�
4�w�`M( ,�f\��+�n�j�s����UU�ܔ��v�	��[����aT�jj�iN��¾�PW�w;��J�#ƅ�}��}��딞��Ǉ0�;O߾M���<�"0	�鏪�:7d���[��!�t$Ցw_t�c��`�;���%5%}���������	�uJ����q���$n����;�:r�h��g��3���M�#c����9I�������J��x�v��~�s�RG�B�`�LFoj���zb�8�g#]S�ٍ6�M�Ǐ��t<SE�>��8x2b�!�2e�Fx|��G[����t�\���,�ݙ�q�
����9�f�)W�	��WV�\*�u�������R��C����sޔ���Nc�k��p!δ�K��{>n��7�=��u�9p���I:#����<�r���Wg!t[�u P�@���\��źb8�Ac7�/��&Z��]R=Ɩ�O��f��5]�^�{�O�_#Y�R��u�T���cD0�Ễ�\�Lv}+o��;&V�脓������G�$�P'P��G�,r7ģ4����,�Qr�.�u�	����B�"�o4'��B, �]e:����;}�|i7�:j���I�u����]ޤ納7��v;�1S��Si����ӕE�k�T�:ˀ�G"yt�b����7Y�mS��a��}r&`;:�wIV���n\h[G���:X���}_U}�D��o���pG�@S�Y���&	�$t�5 ��.�c�����j!J`��z�#w�m%@麲Э����uxh�;�쯹�1��K6��ʢ� ���0�u���h^�.��;��}����<7"��o�n��?bs�D@i��-���Z�����CSM�]���e�f.�* ��6�ry�Qƌ&��Z���vPC��h��#M�%��jˬgb����}Nu�L��n�޷�N�+��-��[�#�wlUX�b�$.ȫ���Bam�r����E���;�mzf���'���::#�����&�y�h�]�bm^��9������|�0V��0�k��;��뎺V��"����U�(1Ȗ=۩��l�"���������iD���"��٩|��z	j��N�u�"����U�����q�<�KrJ�"���n=����zPPxj�gҭ!\�W�7֬!�w���W��ɻk�q���~�;����u*|�#�Ѓ���ԝ���(��@�3����9����W��x�mvԝ��uѻlHG;��y��O�
�ד���͕^�p����<٭']3}9�Q[.^�xMF�n�yW�N��{��6�M'��m�m>1�n�=:ۭ9B�������*+����
ju�D��3���<O�U�������]��>q�\h�D��v0Dv.�2UT0,��>����G<��+hţ����B�Tһ�9���7�q�9�*�2";����@	�u̳��;��p_Ͷ�u��עȹ'f2�͡��˾��Ɇ���%����T���U��@��.�e3�щPn\&4���o1����ై�r�K7]$�,uP(W�p[kӗYB������ځ߈��v�[���508�Bj��Z��7pu�y��P�<1�\J	᝚{չY��9\��P��ѽN��	{~�h���,�Bv�|;jQ��r���l	)P�"��t�;R�1v����a�U�/j+U+�ܾ9����=�#*�Bi:�s" 
���? ��Y<=�a���tRtk���_�
]$s�3�9v��m܎�wV"E��9UX�>ZiD�'C�RqM�H`$xED����_�¨K���f8C�d����KM����
�w<z�Ny������H�����r�Ä�X;�~�tz�`�� �M��b}nc �>ʛ�̧����&�R�ƌ��	�=f4]�����V��E�8��|�JK�5;n��B��\Bop<��FSF�r�+�jd	v��5Æ�j�U�Np�e�q�;R|nt$&ɘ�k=i�A���C��>�>�蹰����_a����UV��]e?��a�c�=�����4�%mF��B��C����Q{ T�[��v=3_P��6C�����?`�S5s}#][5���*>2	��:U���$�{�9k�n
��p`uV]�ܪ�_؝f��dF��2�Eid�����Z;Z7[.&2��e�nC�+�]*�2#XϣF��C�!���T��}�ݚ.��F<��0ǰB�4+iye�8G��<p�#klA^���_�+*��l�:�b'���%Ms ų��wvL[��Le'��ݫ��y��/h�y'\D�?"jM�D=����[2�t'��VՌ��nnů{�V�?|Պ��<���hPث#��[����9�����ɠ����>cG�`���Ǘ��T ���(D����Xf3�W���p��?t ���f7���J�ٷ�3{��#�S�,���|&��� �")�ωW<@8
5�'���&��Mԏdu����<Ί~"V����@�S�B�OND>��m�����W^��y��w���,�,K�fV1Zs��Ӗix����!�w:��`~t���9P�!ܔ��깡vWeN�	W)�|��k��a&�2WS��g۬�x@�gl�IѪ�G$�b\f�jb��l�`Ũk��C�>�c�f�w���lʺ���rƩ��̓�Rk��1���#�\�r-�~e�:��FB��qtʇ�r�;n���=��)�Ĉ�n�\����=���9L�<�
tH��qU2��|s<"���v:��Ӷ�z^%��x�:]'_q�(�{��k�wx�%�z�(��L.5�{��8�|�F���"1��%[����맚*��ܥe�c&�w�W�m�U��to�HJ��(�~!!�(�>���]��K8�y�"�ݲ�y���\Kϙ�<�"0	N����:7�I|n]GH����b����i���_wQ�.^T!�-��J�M�A�)�`ix���.0����C������ڮC��,JZ��"�=6�-��1�%1J�<ۮsġ>}�w�U��#i���Q�s�P.zD�3ed���-�=��4�������#�bxz��2��o˽E�k��%�۱�{2�{\�V'��)��6sK&2��n|ў*<`p����t�]�Ǣ0n�}�@r��x���	Ϊ{y��5w�a	��QW5��KZR���:�� �OV��E��(�XdՎ��r��V���]®��1r9)��Ͷ>�(3٘fӠ�B�[\&�PV�-
|����u�$'g
λ��9��{OP�81X������nP�a��g��=X德�W��3cޮ@�́,�ﾯ������{g�(`���.%��K��{�������s'��.�� �.Լ��*��}�ނv�.=@M���
P� *�W75�[�!_�.�`�k��k*�w�<I��Wl�ʙ�{1=X�ZY)H���Ƅ8�D-�a`�L���ym�&b�{����pl=t��]�rqRoW����z���RZ�H���S�G�q�1(��OD5%�� h�4}�ڃ����O_���<��h���4����	JH �O�1�T�s6�WҊX���zd�'p��Ų���;V���:z�q�):�!�ܩf�A��$@	��Ϧ�B8mnF��N:wx���}��t���q���m�,U)���,�"U@��%��@��n���oKp�X�bc�Gm�$� ���3�h�i�Z�ǑVdHB����Վ�uSj)EM}�rK�J:P�஭�t[;�~Cc�EBJa�ͺ�^C5��.�a;��1[�ɱ]�)r�J'f�a� ](-������9��'��~��S&OD&�o^Ue�P�츷sh�yЁ[S.��$�Yl�%-9[f��f��8u
���ܡ]�i�������&
�s�t]٩.�\�N��*�sE;����{�c���
���W(�2l��X[t�}�F�8����(�D*\Q��Im���#x�I�y</�}}�DD��'5��{<2��
~�&;�ޭ3�ϯ�o��`���=�}��US�����كց��_y�=#��s������;u޶6�y�(�P�P��L`Ta��Q�)�b�������v��׽�IQ���������7b�o;r.{����u\��p[Q�e26��e �I�; ��j޽��tРi�V�*��8_åNiS�<̈:{��	�Y��0ѕ�X�m{&9�w<}˻śx��(�CG��tp}3��1su�.�_�zb�y�u�<̽��Y��3��!��䟘0��� qW�˒�Ъ|k㒠u��ι�v)��+���n���
⸫̷�2ҹ�a鸠�[G�^#:�|-�����Ut����%�1T
�@�����oK���HYI7�\�.�p�꯴!zZr�K7�A��� ��LPkkӖv&+��=�Eec���n��8��Lc0�m\>ϊ�F#lƫ� �a�'Ga�aݵA��
��qΚ�WُUIC�_^
�R��ы��v����N�Îɔz��L��037� �X�/{��{�dv-���1�S-|˝�g_b|����p۽-��ޣ76͊��x���g��8�����t�9�жG�����q:S��[9�`��L��Y)���u�u���ܛqp��}HV��ζkf�%�����[���r�}_UU}����/���<T�^E�}���{qW�q��NS��tF�p�`��4�N�\�
����XQ9o��o4�����Z���L�A�ǖ�_�
]$r!�膎C���voo�{�cu�=�{�ˎ��M%�D.��@�9�RV�3|k�$��*�p��Wӗ�;�$+�l��<6l�p�h	ͳC~�Uq$.�V*T�!�S5�D$�R���si���o4IRav�\9��w�dT'��U������C��p_���±>�W^^V$�S�����Zp�6�]�9Q�2&{lCg������d{�I�9^��,�K���{&���s��N�t��7;�,�F�Ҧ�uF���稵j.��v*�meD�Q��++U��	8�x垸��܏:޿S]������z\��Q���#�}iq����y����c�<�'oJ�0��mG�
�����q/Wy�^Տ��Uf��ȳ�j��Ggm���ϊ�<oG?c�IT0�O��yo��VV;8��cʺט�e��� F�^�����o>��v��5��;kZ���9պ��4����9ʭ}��.��.E��i����kf�h\�ܨ��ϭ[��LT���;mu�1u��[u��i�O�u�;�z���Ѡ���)ͣՑQ�^iܽ}׎)����:]b
չ{�BkBk��4�15������2���XtA��&��Z5�ofZ�#���7)9�l]����)����Hv}�Ƣwq�)��&��޾H�y�V�!8֚Q.���� @8r������@m�4f��%���U��D�]蹼�N�=W]W�ݶ&DyB����i5dV�H�5:�M��1���`�2�l�U���}�P��0��6��w	Ifeu��>m�XN:%��ݪ�y��L�7�Y{�f���o�o.�Q��ˇq}}v�sy��5q��3� �0T�O2Vn��GabU�zo�}Ǐw;���E^�V�D-�#x6����]�Lc0(x.9���ՁsD6��{��;|�]^7΋ZH}mT�ʷ:l�r���Z��ibvtf��Nibjn�7@�]WKoqw0�v;A�_n�Z5�=��񙏹r5p`�˃{���G7̚�=�;�@J�8g_.��.S뾮֬�t�2^�nN談����7P}Ҙ�W')���Cm���ws҉��Vݭ�V8zR�<�98��,���
�"S�{*�h��.�����R�{԰�Q<��
�	#%��E���WC�B<��H��uu4�P��3�W�wδ.6���j�w]�r֠\�����wu�r�,�i8���ހ��*�Sy��í�6"d��5ngm`G�
��0r�i;{e���� �Kt��twP�D9��Q3�5+x^.ʙ�;��K(�����s��%�y�,�xk�M[,K�j��[�=�@俺����@S��^8�^0]&ł����۬�u�ӻX��\2�2Ika��t��ݹ<cvMͳ�"{a��1S&+ﳨ(,�_��G��o��g�V���rY�c�U�D� d��c�WR�.��o*Gʄh9B�k�.��mç�}�ݑ�y2�"����Yok]%���Σ���d@$xmpwyY�Xs]F{��U(<�{hw�!:���50�اM�{�00�����3m�-��v]XI�k���Lwm�>&n�6�+Sg{^Cؕ�p��J���A�l�Ws��9�eŃ-E�pm�B�cMf���-�D�9�[�Mg�Ԧ�B�M]�̲ز����p�ϫh���#��0N=&�	c��[��B�I*�F���͹+/Y�ܾJ��S1��BH��%R��;Hjz�ue�4�Ȼ{r�#"��p��Aǫz�YPI��sQP�q�r��
(T�e�+���+f�vf��-iς|��l{x<���{r��q��%\!��,���\xÐ`���xJ�UzY{�;,&I/)<$��fHn��BIr�t�)��v�0�SNtd�r�QﮏC����2'�љ<��0���!;qs���眙�I�<p�wX�:�f̒y�o4L�த���\��1�u����y����y���A0�Q&��7M�B��<yKƸ�7c�̔`�	�4\����a$���rR)�DFf%�أ#ι���;θ�Qn�a�.��ݼO9��v�2PL��;�1��Sx�Fh�e.���"\��6���ݻ����QD@A�EJHjLD&;�H���tܐ�Idn���Fh��a%��M�&D7d�<�;���y�,Ax�2�u��C3��I���ff�H,i$�'wII�����+��7:Դ
����L�o�����������bau6�V�)�8o9�3]�4:p�}���Cz�7\G�~�>�">���Ic|�wA����D�ͺ��:�v�nĎ�Zx�̥��H:��L̸#~}�9��ꊽ\�=�UE���|�+�Ml��W��]0#&�j/E��+J�֝4����s��Gl�c[�����z�\KO�
�Wp��\=���}n���]�T$7��rZ!��j��j{p�5�Cڇ����U�4����mGS7&�/�����(4�O'+Y4�v\%�s�ze��q6��Wn�kMuOi�Uf�|_/�O�6�y��[=�]�iUĖ�o9�.c��˵ϱoG����T�L�Q�.���d�w�w+�U�}��oW;sS~sg,�>�������*{���)�<���k�r�U-2����{#�i��}����¾m�l8ƅ�NبSnx��i�i�|�<����WG|�m����¼��.ډQ��I�Pۍv��Dk���2u���y��՝��u����<�]�伯���\�;�zE��:F���F�D�ʀ��WuBm#fqᦠ@O�K*>U+����ܞS����N�b��y\��__[j��ᲜY�A��x*��*͑�}n�Rn��z�P#ypQ�c5O���>���--;P���Y�?[�r$9{R�Nx�ޯ�n�mhit�ř�1':;su�{�4�F~��[���H����=�Qސyo��/���U���qԱ֮����Mw�bߟ�#����}��s����s�*l�,ǆ�3�m�S:�ǧpZo]ƹ{ٯ����\��s5~�TY�x^����Y�*�{{��H�p��|*.qpS���ryIK��m���YS�+�����޳t駏/'��*UJ����P1D�ܹ��i���a�U��V����q=o9.�w��5j���T��Q�����|�Z�lt=���}q����5b�)r�p��y��_��rn)� �i�Nt���KӮʚZ�\>gF��]F�l7}��}ub������w�©p
`��c��#��Эd�G���fp��gc�����"�y�):n6��_r����Q6�0}5{��G��W�>틭���c��jѭ�ԅ0�X����s�C�4
Qa���IK�c�Zjë�B�ER��Mb��*�{]8L��8u�b���\���)���icY���W�2��f]�}��3�5W���u������}_UUU�{{�$���q�+���ۍ�����ΩM'%����n�D�V��$n����G�vpp3z���{4*��W�9��C;��{�r�)���O
���m�<�DLB#WMD�̄���	.g�|��4.�C\b.�2��xf�cK� �C���%�MF,�ar�+��y��8�Anc���n�u���:5��v��*�� �n?�rϪ3�'��H��19|��i�_������s����5��Y�1TH���]�?��V{ȗ7�l}Nou�o*��J�����3���;ɻ�Xȷ�v��n\��H\��Z��c�\���좋����~�����qy�]�X�+H�M�G��Ð���.kU:J+\@���&�*'P�����T󋂞>��z������o����ws�w��r*͌�\�D�}Ctb��|��i���DH������^�jX�v�G{��n� �6s�#�pw0��������yF�e�֣��D����B��2i��uB�u&�}�.�|1�B���ϰ�uE�;Ǩr�w-/��и����E�2�9�l>�_k�{�]�}%�����>���>����m��u�^�Q�l�Ս���g���ڪ�����%�4�˹�U�wk]��Od��u����Y�	�^� ����g4dizu_x��6ǽ]�n�+�7Y��������.woCyoC�m=�����*� � ����byV���i�4Ys�������������U����ﷴa('�5Hߐ<���(�17-�c����)]����lg<f��)6"t�j�{d�E/�3CQ#S鰶{qW�_u�楟3�.&�$^U�[����y��=|�O��aut�u�9�ԭya��hIsP0Y�!L�ֺ1iwn����p�pw�'Me^.��Z=�G���5l�#�z^:�[k{�r�\��q�����۞�_T��,��#����.=���dZ���5���� ���q�ќ�Y=_
[y\�Ofe��t�G%#N�6���t��yI��冰mX{s؈f�im�t{�1�˨'��_4�[�v��k	rN�Fw#{cj��H���V�I��J�TJ}&��{Z����51v'Ɲ%;3q�9���qi��U}�W�6^��쳿�4k�j�,����ż���gn��q���j�N//�1��X��^�f��k�y��++P��Rq����1�S�Kin�F/�[�+s��0{�����*'�3�F�c��yw�m���yN����d~�ܳ^{5T�аfW�¡��P\i�$(�����]�}���x8��tYm5�.�o�����j��H�Zy���J��q�uWo_sY�dM��J��{79M5r��|�*�݇N��Չ�����>-��U�9��9��ξ[)\n��zˇ���KO��]��(.�S�r-�t�C���E̨09q�"K�p�T����k���y�f;F�g�����VΊ\�����lT�"95
�M|�vZZ�hO��iNQz�_<�O��r�SW�t��&4��F�鰶~�zک��I� �X0!X��������:+����)߼q��f��
�e0ߎn�#{p�`��R0,�|F|��bKfPqu��Tu:��t{Jh������2�\�-�-H"�<k������6��k;�&�J�V�Z��̆�P �>������������|io�����E[ci�9�2Uw˾���9�M�]dr8ۼ��+���>�گ�i[/��gm�l9�4�\�q�m�Uw�jZO6��ε�=��*vG-Tr�j|�ˍw�9��_)�;���z$����j�w���2GޅN�u�J�E��m�>�g"�P�!6� ��1P���R�wF�ȉ�±����w�������3�.�J��ޚ������S�u[�/�_G��/f?�K��o�����jѥ.��y����ڜ�%k�Q�����w��'/X̢�j���s��VKr�{\��{�G�\?�g+��x-'��\��{}�'-`��zr�~|�͛���\�N��KӸ1�q=��A��.
x����{Սl��V"���wi;�p��_5:{6ul��c��uQ=˛�����}�p֭�P�w���{��v�^f�:�v����K=�/��G52��N��+7�wRj�`�] {����q��^��{�Z� �fz�e�0B���\�b�oG/��9ݛ|�[t��N�p��Kf�ͦ��mF+;�-@:N<�D334]u*��ګ������R;u5jg�H%t������Tr���kc����O�L�W�!R`b�.ych���AZY�)��~|��=�2�Z�SK[®yF�n-�B�ĵ���;/�nr匬n���R�;h��H�sFO/�y=t�>�%����{^��+r�ֻ!�ͨy�):n��u��?Aߒ�<�]�ɴ�ns�k,���bq�f�J�B�g|�h������rZ��Q�9�=���es#�1���C�]�[1١W�4�!�������sn]�T��b妔I:ԌU6鸕��9�Щ.f����8���߯�p�mZK��p�|��k�8��j~���=7|�c~�5:d{���E2�M���dނ�����F����۞�O�����w�\��]�q��"��G7����Q�n���s���; Z��E�ډ�vs0�=:�TQ΍ C�<�G1��x�:���ta����"�}RY�~��z �v[e+�@ȫ{�hn�,�v��{�.�WH��Q/ �]�zFN�{"�y��	������>�8o+]>�u���)��p�����yʥ��[��Yݰ��U��UU���.<�Ow���?�XQٵRg=�ޯZ�l�󼛿���o��PI��7�S����Xw4����Օ�����$���垼{���ї,�l�z�x.��;�V��Z�\��Ss���:�(��0�8	����߯bn̺]{<-7k���ep7�"\�P�`b���'��a�p�9��T����;��xߎzgzv�{�Kv$tz���:GѮ���/D~t���6�m�Z�+_L�\���&�\K��G�?�ݫ��E�D��2U�Y�K���=.�����FU߾�r��\�7�CΆ�����p7
�\����"{c��k��M�c���\I]_I�v�dҔ���[oC�y�):n�n�#�gGl�t��#�?|e��*�'��]�?j�R������ί�3�-��yT�4Z�b������'�ܶl%�O��ݛ�Դ��jQh�������3^�=���&��{يGA�9z���t�fëy�$t�(���lgM�[FoU�Wj�ɍΊ����w[Y��Qh�/yQS� \�Z�ER��/�����N�l6��y' ��K��n���e8�J�yy6S�U��UTSjN�x�1�w�|�,�:�.��Ϧ���.��Г���#����릖>�y����{�b�]�R�����/M�k_�'K�!��EԎe�J��j7ڋ~��D������a�2�]�9	���=�6���=1eHc���>��Ͼ΋.YQ����k�N�mƴ�F�ȟ��{GY����:�oRѷûz������9!���"��w:یN��L�:���b]�}8��
!��/M[�Ury�K���JV����N5�1��[�D�;yx���F�߽��zmx]��nr�{�*;TOՏ�ŗ���K3lݧ����:��nH��ͧ�
��{�+H�ܫ��Y��uzk�
)���>D��W��r�ޞ��N��]��7�Q�l��X�Rz�1��6 �N�9Z��u��zm����s->R����_&�z�+�뒱��.���7�w�׾m@�JR��޳�iM�t��[�1^s���W󶋒��:�?1�p���J��{�j{�v�{L^�����N}�;"�e`�BnJ��^fTˋ
���C����L:q�Y��J��X�V����B�Ҧ����$��_}�U|�\��{�w߾cFC��al�p5��z�z�_��ௐ�'AY�`ד�^V����;���G����p�T����|���{J��%ۆ��/4�3�k�=��y9���U�N���0Drj��R��agt��I+�m6�uB�r��%pP��&6�Ϧ��u���b����H,�{���r��y�r�m��uNiL�Q�.�b�NRE��7�[7��h-J��D��&��L���snj˚�Js&���|cvT]<x1��"Ý�/tr���[|�\k�r�;��s����J�&��	Pژ/rKw6�cu⿹*5����!��V�7��=\��<�c���d�Y��|��������_8�G^�}�wm�M��%��v0�K`mBx��F?[��֗�$~�V��{�|�'u��/8M�
�sȰ�+Ajw�$��Js��[��F��f��jǗ�N �1�;��l�;��l��}֯Y�rJL�����N�9�m9����2d�A�	Z�T���k!�N�~	��;6	a�MU�(�u�Qb��o�����fG��ʛ��#�-�����V+�Uq}�`F�.�>7��<�1�;���n�*;:<t�����sk�]�罍��`qw�˜$���d��}]�N���
3�t��
��Z�2�t�][
��i�bAP��tN�-y��<�o�9v6�v�e2�/(�Y�UoW7�r�؜��(��y�s3nٍ]�=��J��|uE�R��-��(�sui�XE��C�����nԈ�%#M�bZ{�ʻ�8M��}���;��kQ��&,"6��wj��2�O|�\�0^|��;#Qj�;����)��M�m�k�/�۝���я����.%wON��%b�4����U�NTGໍ��8h|���:�E��	n���a=�X��y��9��K�*J����bΛ�v��.��ЧÄ2̣z�-s�`SJk�,N�v+�l�E�һU�/����5�Ha�!�b��&�^]l�1��4uی�W:ʅԺ�Z�i���۱���
rN�ea�ZLgwR�O�'덬�a���7}�j�=v��tb�SQ��0����G_>y` ����ܠx ��Y��"�Q��M�Dp��2�&�%��7M�gh:A�)Ϸ��y�Ŭ�]�8��6��1���zn�u���CU��̬�"]�6�(�(Ŧ�]HA�q���T5�������dN�����A��rka�dRȳ,��LMR�ʼ������9v(�AYj�V�'�������]7Y��6��ht�&�c�@�-�B��n��Y�O�$�GR��OgP����ɼ7�lc�KM�0�����W+8�LlB�S]Y���5 �����.��N|�vMc��S7e�N�C����[�("��t�ט�<�{Œ� �}9d2����A�
}f�[:��e��R�|��,��(��ŕ�ʗ��i�ɹ))��J[�� 3�6��r��6Ru�A㻶K�[n�Q�$�+�0�Ck��غ�>x�֔%�5���2f��@0���?�JT�ct��gqx�.��qʗ@a�v�;�#��	�Q�z��+=
IZ�E��r�:����t��`�;}�q�/^Ջ˺ސ����(*YAp0A�1Y �l?���n��ީ��Ӹ�۫y9ۚ�:i�ú�gǕ�P�7x{b��1��@�I��R���T�u���)(�� Y�	�߸t�lQu�x�%\]{��w499mJz�ܼ
�xn}�'`�WL:�wm����$%(;����p�����[�rѺ�.Q4)vffjƊh��LӾ\jq��-���+>�f.�3{��`��0���L���Y�딙B�Sre��.u`Rh��77)>>�`�*���������GwQ����C��"H�]\�wN��-�q%9v��c��2�x�$b2L�rݒfD$��D��� f<\I�"I��,ĉ�\�4��"����
�wq& �i��!db�`��'��.�LLRd�e F��S�p,��D0�B$��0�%&'���$�OB��ĀiC&d��ݹ2&�	2h3.uwtGw	IH	@)�FE"#%	�� ��7&�FY#FL9F��HB!6#�s��)���q$�"A/;��M����� ��ιd��3D���idJ&D�2#B�(hWv���F)!2PI� �� v�9��xJ<���GZˮ��Y���͚�̝Ȧw��kb����_'��j�J͂Ve�˸Y�W"a|#}�G����k�W�����S�q�ƻ�r�_���;��b�~��Fb6����t����n�nխ5B�k�7��zV�I�r������'.!`̢�z&n%ƛ�Q�,mV��K�:Z�Ob�_|��)��o7��v5��Q���VA��j͵)�[��k����OOTD�}Ctb�����SM\K��C�WY�=��Յ��od����U%�Q�al�c[�7��g%�,�r�k��^]����6�f�P	�h�=8�2����\�i� Nښ��c��ל%k��<���}������*� ����CK�� [br+@�Uf^�c��eu�k&����Z���ޛ�)8���l�#tX�l�ؽ�sz�|��M)�g�ǳP�w\#��>o�[c5�)�����c/:��v���ٲ�ڜD7��]�[١jM+g5����_6�*3��j���4�i���xݫ�"��jfq<�,��l-7q��CK��]��Q�{dJ���5/ū5�W�	E��hyS�ݽ�CF�r�����w���T�P��u��y+���]�6�����9mEA<S�&�ꥲN�:W)��D}	c�{�'�ެ`b��WLU���iWy�N��tf�|&n��'*(�	��l�G"y�Ӝ�!u|6���D���y��
������ebt�k귚%wP��w�LF����۞�O�m�ٗ���W�'I�ȫ�*{�/p�N���n�s��q�N��-m}1G�������\��NWz��=�şu_t���8f��L�g7���Ʊ��r�0�3����i�=�ջޫ��oC��.�*�_ǥ`����r�\c�S����`�����m�[�#=��T9��ʨ�c�b��|�⧜YO���3=q�98�No۹⥆��zs�K�P�W���r�T>��(ꁊ]�wu�mLO.��n����W�K�ۆ�W���_�c�*��zή��Q*�V��v��?$�z�������m>��������˿����V'g��6�,IP�OvV�y�O�Iz��8C�7�uLJ�Uc�/�R��Օ�W.֬
�6�i��'Oh�r�/�vTgGo*����]M��Pӹ��-1(ǖ�Q�wYmӤT�+����i<R�!6���\�ŝ��V�O��ZY�S#�����d=���$#7���}}��j��Jɬ�DL�w�\�c[�������Ci����nP�&(�Ur�.}:�!��_eIh��U���Jy|᭸z��8�Bt�Ђ�賏.w��O!rk��Q0]'�c���.���d��I=���UK���֚�ӎ�ɭr]|��1�!(�����ٺ�������اo�,�k8e��:�\�+�]�#L}5+^\@}����=,eܾ{�ݫ�k�;����8¸g!:rg�����\��y�<0w9�y{c�آw�����'bL;����N.9Ӟ��T��a��|��u���;�}�q��qb����㿹*5i�4ۍw�V��p���߻ȷ'K���N����e�Jf8��u\����u��3_E�gj7�n�XV�F8����Y��h�T��ފ�.16���~��W�� �I�u!i�ǩ���6���ff���F'}֫qVV#���
�t��cX��CB��zN�܃��^�d���:�CHɏ��{w�@�4��@8_]���[\�k:��.k`e�#�ؽh��pˡ}��N�3�KB���j��;ht��4x�#��G�u�ͭj�.v/;��+�~�9k�2��Fb6p���j�M���ݪ=il��jg��������{�yÎ�\�s?_��fI\s7q9:w{��jF���j&;˜t�Y�6���5}=�u�{�s{���?l
m��^r���J�_D�>����(�\ܨ�i��|��+:�[<	r.�չ'm����E�9������qʾ[)X��ކ�ާ�->Yy��U8������gE�8�T.���lIJ��W
�M-On��]�gMj��=Y����Vfn8/��T/�L��PiW�y;�k&�;��**r�}�x����{˟�x�9]�T=�λ���Zj�u/��DW��2�N����;�q�n7qZP�^w��lf�:�4�J�h���#ue�'�6]�Z�;�Y�o6����hU	4�|g���C�sJe���47=���C�`h7ԅ^�E�R�Y0ٽ�6v������j��mOf��9��r��i������Y�D뗐;������qv�����D��:ݗ�K$�L��+C����X���
5�Ѐ5�yop�b�J`Vh�}GouL~���Vc�=�d�^�@�Z�j%nN'��}˙�m�wˍv�D����u�ºquh���_��{����w�������� ��&$�tc�G6�)gg.&��$��u(����kگ��vE���C[����b\u�{w��noZ��Fہ��s��Tk0-tf-�y�+/���&��?s33Y�L�k݉ǚb{�9�<5�\Q��3�w{�u�ݪ o�.zN��u눞��>����=+��޹{��+ڱmr������<J�Og��S�>ꉹèt[��\*>qpS���os��N�ieQ��b[[V���v�S�*\��\�J�ю;~�{�79�S�*v߼�:9���k:w���[w�����U�I}Q*9 ����CS��ù:�f'�v���;��{�/�>q�i�Dv�Nh��/N�w�]Ԟ#��u�f����9;�⥲�zb�p��@�e=�z�Y \+Z�����a���U����^vݠ���V���˅�FU܂�|8�����=��Y�̻5; �fSݤ޼�v����MJ5݄9{WWɫ^�0�K�Su�`��B'������Z��]��>�����k-�{Q��V7©p
`���䮏\V4Ӟ����!E���u�Ю=������k�~�������N>��@Ⱥ�;\E�&�E�saoc�En�������?�]#��7%	Κ��sv.��|�\��)�����K�Bͼ��!x�a�������w\�Ƴ��J!�'\������މ��̿�yL�Ϻx���!���K���tQ?qIYv��9��3��1�m�q�f�
�5�'��/cSލ�k:���ǆĸ\��L�bp�DƸ��N{E>�s�]�[.J�
P�7�0��{��Fn�Ŕ���|��Zp�6�mDs���Hŷ��5d,�Dzn�����rv<�4��q���T[�v�nv�������7�H{pɯ7�6m�κI�ރ��{Т�����O]��Y�q�fDl�a�p2¨{��Y�i¡ޔ3�i��7�^4+c�݌�v����u�y�w0�0Z��Զ��:���i<�z��7���n�r�k����h�vFr���U6�s5�m�U]�{�[5݀��Ư�=K����>����q�Q9ʆj;��{�꯼��3������p�].EC����̉�:�b��;;�*yľ9���=.�S�5��%�ӱg4����󆗵c��i�a���gW��]Q�Ǻ.�%oz�m�^�������oD��m�Ƴ$���hv�X|/Ѯ9˞M`��=:j9�J��{nn!���{����}\I|��P�����]�N]�IV��9���=��\�c[����zt6���g+�:�L-$3 D���Sn��ﷺ�O2;��Y5
S���5�Cלl��NT�p-�m`s9�XTΊ\���ܤ��L�IYQ�ܢ����q���l_Wb<ّ��i�ʲ��b6�S��{����6��M����9��N�j꥚)kg7�3�*!�v�S�IY�GB�О����	��.�Ag_�����.#�����_Ű�����AR̻��x􅾷�HgUiۃ��pP�Xo/�_P�z������6t��)v�3��</�"0�Vr:坜�Yu�柮r���N�{�>җ��Y/N0�g
V��阐�+1��ۻXp��F��\N��'�rɂg;��!l9�����¥���|�rz?S�k�~��5�s�_�N�ww�����qq?s�=b֖s�N4*���|���0�~���\Ky5���߹*5�3M��#9N{9�;���Z��evG~��kճ@��g�[��y!�ɾYG*�s��N�Ō����g-dX�6�����0fz���U�ȿE��&��9�l�3v�]��Ԟ�{���q(�c�z���)�����79S���+P�TX8�U_:��p��r���o-u�;��X3(���J���ܩ<�c�ij�u㈜���ظ|�i����^�NܗBN�}�>|����<�u_z��������/KԾ���Y�4����_ ���Y�}�F�0��L��7`j!k�Tr����5���������c�'��M�kS�<;i����.��Q�?Nt�q��]h����j�VQ��[�.�6��rF3���:L"�9N�������GYC5�Luoe���L�����N�9�z��Gu�O<t����u��9{�v��s�=��X�����K+�a��<���ua���%j��[Pg��PFp���>�*�rOS��my���qx�m����?A�#�L�D�M�slfuGT�V��ه^����9[������_<g�P��xF(��T��4����խ��Բ��\��{�rҶs^�|�h����:�(���\q-�}"�г���Jx�?���\�`.�з�L>�A�ob�ۛ8�vŞBhsoq�wl���J$Կ���^�+nr#��
�s-�C.5֮S���٩m�j6�5���T8�V�b�/�ճ�C�Ý�r���~��/��Q'+�]eyE=ť��z��?o�eDk���v�\
}O>�̯�c��X�s"k�yuO;{z��kUm���6�u�����H������%γ�
+s�zT�����DU�LҢz�Oc���:�>����ʽc0>��`���H�ɛ�V�[�˥�{x��b�oU�zV�'��\�6V{b�pż����椵���pk����G'�讣GpI`R��B�Ly��/<����W����9V���ߜ�&���;����79����Fm���n�}��f���og��1����{�.n���U����yQ!ǈ����չȳr���s.#�5��_>|^�^����.�Un����0;Y����:�(��\>q�<}���_7j��X�i�;�����u���_:��|a��ў��u):{�.��H�)�H,z"\�=施�c������Y!�s>2���C�S���܅�{޴ͱ3��e����g;�4�����ꅽ����;���%9����C��_�ot�+��;�5�����k/��|�{ecv7
��)�;���HV)MGN���]��݈��'����MD)O9�Z�|3i��黁�_2����s�6�^C*���S=��&s鿂��{5�)]���ϛ���ݞ�q����R�H���/��`%�ƴ-���	&�g5�3"���a� ���ڙ�4ݯa�S��J�����'�_J��	�hJ��19{��$gR�͵�K4R-�������1�m�q���G?`���W��.���S<��kk���|"#7* �k`���:$�a���v"-�k8��g��ӥZe���tLɦ�g8�k��c��.�mLё������
��;Sz`B���B濫�4\�Ȩ��M*GKݥ�%w*�,`%�xw��gU.��*�Z5�;���o��kd\�����\]F�2w 4����cS�j���Z�1��*�zHO�}2<
��Wb|"��wl-Sx�̔e���e!қ�����+���sF� ���Xv�KZ䔫�Iι��y	��ܫ���$��q����<��Ym�(��a��6�]��2��wo9FL6�a�6�~���r����
���kü�����%�K^��8ꯐ�-^Q��7�^e�Y�z��v�hU�<�/������c�a���TE�wwM�(6�]�۸ڬ�ц�q�1Z��-]w ��]+�
Sx�}O�9��^$�%�!�]n�W�fm3'M�8.kQۑ���9ʎ��hbü��=���Z�E�̼�-)�Ѣ�p<�ŭ��0Pw�^"�t޾��ץk�g��5M���dΗɖ�����q�CT��.=�ť�����;�5S�u�ysy)��Ns'4q}_T woI�e���S��Z�@��Ԍ�ۂ>���A��.��E6��T�,-�C��u)�Kx:^�#91�7�}t�F����۰�Ã:�
h�7W�1���jܓ^���eK�-���Y���nQ��^�M��j�c7Lɉ[�f ���˹��[i��	�I�QZ�9�J�b�sP̥�2��|��du4A���͔e�A�u�;�4S�2�a�tF,���LwFB�IV�U���J&�91*u�X\c����X�L!ot�F�ɂń�:��9B��a��Jk{^dv��I �'��V�h��8X�pU�Z��60�^�7-��e�s7~wy�Ζ��}�V&0x�\��0-df�d�Gn}�@��˩�:�+j�A\h�Q�n���[!���-��zꊭ��^��ۃ,p ��=��x�}��S7*�|)`̺������y�ćF�
��)gVq<�B�=$ô���7���7�O�,�t`64�LG���B�-�I����u���z�P���]A)\�jR�nc�rĻiVv� I@��ܩHjiꇱK���{8��#�G��2z�ŅI��E�j��X�ԉ75��oe'���xw��7Ul��Ig��#fUֺ�l0JV��<��/,Z��Jݕ/nҺ��xM�u�=� �2>�0��'n9�[<2�1��{S�̀�l��	І��\t�XGm����=av�:#�]�@c�݌�ꇌ�Nd4GJZi�TMBE���q=��c.�N��A�YE�Gd��^rt��Czr�fu�0���j�]�𤐼��V��I��KėJ�.�f����K����L}R�m�1��
�]-�ۨU�B��4���%�Y� ������^�p��Ju�&$!�6Rd��""CB�d��]u»�P�1H��a��RLT�	L��Ӝ�H�\��.W3I�7F)�dR��I�0�3	0]���l.]��C��� �)�"�2�f���H���
(D�$�Q�30h  @"D"H.��2Jfƀ�"% ��d���``�(�,� J(� �#aH$�fD�@��Da(4 �aF	��B��	$FHQ%�L�AiL23#r�nn�1%3��&�3(a �Hd�4C$�(i��P@Y��P3H� ���2dɠ(�JI�Ļמy������������fv�έc���٫���vഞՐ�v��.	d��S�&�(�]�Itl�o_c�������S~��+[�;v3�s�4�`�ɸ�p�Dƺ����M�ϡ�z��^2�u�Ĕ۝��[Em��j��o:5i�5�n�9�~�YO�<��/���H�^C0�=;χs�k�W��ǤT}=���TO�٧��z�*"�#��蝎��2��${M���z"3۷�ړ�_�Q�qT�s�������Osʞ^J�|J�����/P~�d�&\��"�s5~����G}z�u�>u��ɚ�sKrJK5u��'T��i�<��X��V��߬8s؎uz\�	��c��y�o�Ջ��J��Ӝ��:.��O6�U��\U��*�_2����H�	�w[i�J�r��Bځ���(��E�����|���Md������09�λ�}�����&eD��W%EtcTކ���z�x�L�U�9��`��
���F�ӆ�Rv�RR#��+Y(����_.�[l���֧;y�c4%[�!&KKj�׏Y�wYw�Q� ;{]�_giۦ�%��L��ګ����p�����&��q$	���+�kr�m{9w'�to���Ʀ_
W��Ց�VE�>�������j���Cg˹���q����(�3,�%΋��|��jt�����Yf~��r��BQ0UVTm7(��P�CYב3\���g��c:�3�eN'%������J$j}0��
�4k痵:��և��r��9\��k>gpSl�:�5�<��tt+H��w�3�O@��t�ٝ���9Y�������|��a[9�v�"� ��!�Ր�����Z�y��4��lԥ���hK�Q��L;eƻG"a:�_ <s%����q��zǺ�)z�Cn`�̸�o&�v�{�Q��N�mƶ�rl����/Z�k��ӱhO�t��reZ�*��|}"����Q>{�X]ɲw�I�`�a5���{��1& �G8�Z�l}�f���3�9
�/5v�ͧ���g�r�q���,��e�����~��j��E�3��u�w�.�N��.5B�rq5���S�.
x���Ů��y;kenE��z�������+�� �T�OW=��ީ��>��XnrUJ�3P���E��e�ܣ����H9�f�nr��Ψ�VA@�����K
��$��e�w��#�,{Y�u�Kz�ZyȞ��,������W���Zw���O�%N���1D�v.�8	����͸o{���損 f�y-�Z��pځi�O��ށ�'���̴��Z�gQ��T�r�f�6��a�o��O��JK�Qʖ�V5�������nT9��t��M:�}�ɣ�vմ8�����X;��s��	3N��1�I=]=<$�^��+_͎{p�=����n6���!�P;���pzQ����9yڕ���w�(���-k��|3���C�J���)1��%�R�˳u��*���!�қf;�ZK�s^�7�*�P�ҙ*U;�,ek��ϭp�e��8�od�w�t�hU	4��_l���v�\PSUJ�N�b��N���P��\ԭɯ�9��s=�zH��]S)M�[�j�q:�ȞV�4�#�}Cj~+rh��U:���YЉ���U�3��\R����~����{�ٞ���rD���&��J�6�u�;�+{���K!��hJ\�^}~u3&^"ٲö��HjZ-��gtT��쮛)TV�u*U����{W�W$[Ks�p�(�cs���h/���N��le�0u(�5:n���G�\�t�շo4J>k���k�g*5�G:r��O���'�*%c��^N�����Sx���vU��U��2�ہ��V��U�O��Fbq�]�u4��4����qg����p��<��ެ��x�k�'��g�������m�ZB��J�]�.�����F�OX��oP�(I��/{5�i�;X�}9][�1yX�z`�g��լt��?�u*��:3��e<}2���;�����7^~ެkg��L����F���GT3�������y����3����O}ύR�<��p]`�!�D��#�Xh��r�V��י���lO�N�m>����Vu-ힷ ����,IVI[����ܻ��%��\������5��=m<ⱻ�R�qƔ�ɬ���u���	��8���r�Jy���mC�9I�z�)���<b���Oz�p���8A����9�Ţ��u.Z"륪��#�CI��m���x��J	fB4WZ/[v*�ۇ�Gq��w�#s�Qha��1P�ڛ��S��A�h�ֺkӯF�f:�p�b�)�z�3�<���ʹ�m�|v�n3�W舉�s��O1rW�'0vj'��l-��ǳ_B��h���o�k��ǝ�>�ԓM�ݞ�j������j~�Q?�B޼	BM(��7�bR>�e�ZA~�S�~^ج2���Wy�W���ҙ*��.�B}5�2�	��oʺ����>r?!�c�N�}��G"S�*ۚ�!tl��H�βgSZ%��7����n�s�Q��Sr��r�5	&
n1�#�1��c���O�J�#X1__��07����*mZ��tjӆi�k��k����38�R�*'���2_S�>��djf5���d�eZ��{x�3nQ�U�/��lb�ɏ���!+�{\/}o*�mI�{6�KEw����D�Wb�}��2S���f�s�{��u=�w�1�f�ӑf#���gVYN��Ȳ|�o{_m�D�z�]+h{�������^Տk��GnUXp�{���מJ�3�C�kR�G^5H"&��J��L��ճ@uw��ũ��Y)w�������x�<������(�-�װ>��8S�[.�Z6�B�
�g}��!K�G��wI��E�g��b�Q�=��S�R�H���j��e�
�5�u��M7�U�m*���N�ש���qLw.qer��m�U�a�I���s�`�'1c���u�d��r{��qTOC��d���&;nnO�%�낳�5���e��NU쮫RP�t��R_TL�J�Q��z���z�xB�%JOt��N�xR���#���)p~;>D%�'��W(�o�p֩�>���dDG^u���v��Sl#S�ޱ�U/�I�?�CJ������_T��/u��综��^���_oU��<;*}�Q�"O�t^��?^\�^w���t�q�rҶsZ�gpTCl�:�(���}]?/y�������/>m{��_N�9���{4*����_p�0��N����bL�nA�赖�z_A�U'WMD�ɯ�9��
���jL;�eƻ�r�����؞rf��LVת-�5\$�w�2��O&�v�{��N��=�j���GVə��J��=��+lc
k�36M2��-�O�{:�p�|k��$jȒ�%I��"�5��5ĹƢn���1�+��!.��=�L��D�B����n�I�YX:5
x�.[c���џ�N*ޓo������]���
7:�[�y��4��Q𽽣߫��:��V�\|���OL��~Q>ޅ��b�݋�,t��o�५�8Ҕg�㊾�T	g�M�j���~��=.&f�{3�U'�r�7��K'1�+-'�w��ܨ~�9k�0{�b�����=����,zwE��\V.|T�)�l�Zƾǫ�V{�-/q����}��Վ��Fܨ��{
<���SMg�.�m����+q$���S�O՛�7���;Qg�����}cv.nU4Ҍ�U�r[.��<'i�x�Y=:�] �/�"Tr���W[���
E��F����ٚe��u�O�
�Wp���pب�IJ��Ih�p��cH��؝[�ֻo�o�|��=����n6�؅�)��Gp�p�Z�����z��56����_)]�cZ�^��3�꒸��*צ�х���;��7BQ�}7jZ�ʓ��d��Gq���i�*�]D��3981�bօg�����
�4��=OџWZ&>sx��*3Ϗ_%���MFE��+]�(��h�z��ĝ9b7R���Q�;M@O�h]�j���\�m3ݖ�6�e��K��/כYz�����v=v�p�k܈o�TE�6�S�F&^�h���
9�u����2S��)�[5+^\��f�P�J���lf��h�F��O�o<:;!��(���:|���'K���*��s��OT�Ci���ݏ�n`���z5�C9��_)�5��6n
ܚ�O&�at�QR��F�m5�����p�Q��<ۍw�V�Ș�nTK큶�{3�5*��}�YoS���ws�~�ڵq��o��nl79�,�k0-w��KَPW&�E;I�T8�ܯ�`�Ʀ��\wK���w�Y��)�J室�x�y�l�����z�fuM�/�b���qV$��/5s���t�ܗ�mXzkW����p�7�Oz��Kbzz����T�>ؔ��(�JMO���y7��V5��~ίCk�:����"���]|b�$��2�}jV�C͙ �k�k��=V������ۼ����j�B�rw�$��j��;�іZ����N�Rj�N��r�t�k���}\ٙ|)H1�i�}�.A>�og�3�-E�A�t5ju@x��6-�Q�䱗l*� ��}���2���gN���O~�>+��mw2�L����}�u�Ш[��N���/�R�����'6�\���Υ����.�Z��Sή��*��/\�s�r�kw�>c����
��l��*�ϯ˿����2��*Ob2z�V�j������6�q̋��V���Q��utݺ�R�\�,=_/�O�`��C���_<�/<=�&���>���q#�5��v�NC톕m��1Īf�9.�|��#L�X��[=�`#��[u8��U,�KP���gpTCob�ۚS%q
;�/�0���v<_a�I�>(��h��|�6�;�q�h�'Ld)�5�t?U��K�TL��}[�͂ϻϟ�ν��r�d����Q��7������RԶ�f��y���Ϩ8�ķ�X�b;j��o:5�3Pہ��p�rq��7r�#-T�m:�!�lڞc�Nd�i�x�hѥ�*��v;sJ�����;���3�o)U����eu�ؤِ[4��
�r.։�9tй)�J�-�ob4s0��t�
}к����P�w;��3�	܉k=]��]4W�4oP��V�R�J�f�u�銇�s*�g�K��Vr��|��;�)T���F���B����Rogw�=�=�p�Q�d��ј�&�TJ����V����x�׽���a+�%��\���+���ەC�zt��1Q�^���vY�^�_sڸC��<�৏���z��Kڱ����Xrߧa�A���d�����׎'#���c���;�8{T��m�ƶz�*�v#����UMv��甐���=���/��&;n[OTK��Vuѽ��{wO2JZ�Tڙ�\��I�%��r��n�硼����b�t\iV�zo<z����L�n��u���vʢJU���\��֊ɛ�(��E�*�v�W�Ѵ�4;k�r����U�Rw䢃J���s�9��F��{Hu\��Η��r�Q�HZ�m��޺�4��P��#h%��R��ߧ#�5:zA����k6�!Tk5�9d�*��g�I�V�E�³Gڲ�gb�oj��fBӠK`�pu���� #�M���]eG�(]C�%�=��A/&5E��3fT�m��^)d��=g-Ёu��B��W][O��%���QL��5�lZ�M
��:���T�g��I�6��Avv�:��Ej�����}�)�ݗ�y��{;l�6(<lk��1��
�(T�bd�`�k�gSG4�+�A�Mu��ᖰ�86M��-�Jq�n��A�^���TO,�S��)Un���n�̣D
�.P$Et�1�����Xh���q�͉�9n��d���l�(*����ih#o���G��8��걹/ �ۻk�,��᷃6p{��tW�)��I�*�t�x����ޢk1�D�J�;,�@�N�$=�A넢f��:W%��i
�kp⇊%e�۱��h�څ��+���v���i}���J��wG��m�M�7.ɼ�8��R��DZ�9wZ��%g�G� [m\|Խ���Al�#��b;ӻl��b�ˊ����|O֋��3�f�/SqJ;J�L���Xl�S�flE�ݺ�h�cǔ�X�n۫�a�%W�$D&�L8>���86����5&8���ٵsL�P��XR�Qm�t��t��t����$"ޭ]�0H��Wt]��3pVN<��c��՛�n�-�9��lpE[XF�o$萳�.ݓ{����	�X���u���v{�KXf�(֫�e��TR�� �e^�d�g4�^��Bȫ��Ci0���a>���S)ec�.�Q����)@X9n+h�&.ŏ4Jt{&�.�Yhm��[�\�)��`-'�Q��]���hd�б�������f��e����ЯR�o��cX������24�m^�u�������c^�q-�,���5�#��3u[N�Qmh�25��)��̳\%��N����15�"�-/�M�g�뤸U���Ve��ኞ�MµK2�eE��a�jw�V��t�t/w��{�Sf��8T�*/��7��Z�s{������1��`���园t������k����&!�a�@�[�;'
�J�.�l^<��a�����X�N%���u�����\�OuE)W+�	t1k�����w|tt�:6�!l����4X7x����(��.�|%^z��W�
�@�vpn'��+;��ؕ�̡��#7t�ћW�Co	�W���2��x�S�6��=���곴��	o-����i��&���[+衭������t��ؾ#��}z
=
TvE�Ư�GG�<'��{�|�6��Pu�����6^�h��٦��On����P%�[�Y��8HTι��p�7�u�31��VV\�\&w)��{}.V�� P}(��z7�����=�ZJ�E��Ռ7*�j�7�s��ո�l	ؤ���C�Ѽ�����|b˺u*ٽvQ�@�4����Bo���%Z<�9?���h=��X" -$��� !�$a��Q#�&�"�9�(@iI�06%#(F���\�"�DѲ"F�	A��3;���wv≑!��\���rsq���E�;�M"��@fLb&�2L�i�d�0 'tv	�fB .�5%1��M��I�
E��2I��2#$�3	�D�)��$�.q&II��Iˑ2E,���H0�]�h�$J@(�%�10���	$SI�"�ݒ"$D�0�12B6d"R�\�"��$�I3
6Kׯo����{�=~�|o�q�N�p����M���Q�#b�n-ÓOot@���\ߘ��wPol��k�"��}�6�3b�:��9y?�r���jZW��XߛgjS��9V��p23p���<lw���Ec�7sR�e���hT�5p���a\C9���ţ�0v)�~H���S$j�=f*}��7E����c��.VC���m��>�����������ت��ܺ�8�����E<�ʊ�պr��ڽ�ziw��2ur^s���pşp��x��̝�)V���dg��p*<�&e@������Ӹd<>Ҿ�����_���ou����[��\f��|�����P�y�	����\/Pٛ���A��Q�C�+�Jy>�;]15�u�/#=�>�&���5��"T��ߢ��>�UxJ����MǿNx֜���������5K��^�~U�u�+�*��r������\x9t��2%����23{�w�1o�n��=�~��z���G�K��ʁ+���Mi�r�l�:�B��쁟K�?K�M��=)Q���V9�v��G��r,�)_�c�j�C��R7N@j���tB�Kޚ�d�+жx7f��R��B&�p~���AdR���=�i2CF�ͨ�/2oyou9�F�H���JG��g��y6�6�_�s�W�`;�a� S=e�
�o${�������hٸp�P7ky�]�A�H�Tfu�Z[ �W3{����RꊹT)��{}`�zsftKKK�����m�qϮ�ȹD�jKD0�#�E�L�>�a�ո
~��x���Zg�����{�����^"%���;%�9@����$yT;���98i�7�|��3��*����M	��~+�O��{���ǵ\>���ӢY�� ��>u/ĩ���5��9���@)����S��s������z�;�'J��o�'n=wl������^7����q�{yj�=z�ǀw�2�Ȁ^S] ����_O�0���_�l{Ը��3޸<o�̮�ɚʌ(_��;:+=�U5:n�� p�+��n����0�-�!�����"}��c���ǥ]-�}×&T��'Ͻ\���Uê�T�2KF��>�Q�/���?�r+���ew�r�z��ݖ�Ey���j�>�� ;��5�?]x�U����2|�q��/�E\T��зd>��_U�>��ig��B�ێ�M���_�����@w�����B���9�7>
�N{�ju9����׺��\hK��^�ei]WQ������F�EzM���@=�T���P�6o�>%[<�M��������Ҧ�
�a1��P��f����u(���تvc��P�]*)�unT�ȁ��J�C����8�.�Q��f讷O���>yN����r���3b���sڔr�Î�ѥ'X�"�/YJ����/��|�֭�/_ Џ�Mk�vp�}O��]8�^��Iۍ�=W�x�J����;ӟo��ef���۳Rׂ����i���{�0�@������s���0�{���T�A�n�ޞ���,�}x�}3��^���h�^U؇:N�0���wYU�C�*2X-j����[+��v;�<�^��d{�t��;�\B�Z�;E&`x�������W�C������}�󼗽�3��d��OԼ}[���ʣ7���b��:�(e�$�XX&x:���#=�k֒W��ݘ�ղ��]5��z�S�,��z_��:�r���m��4�E� �zw���eG��Z�5e!���t\T�B�*��.̇]��g���!�cr=�|z��w��|c�4�����&'
�W����<�7C�;#tA��n"�P^�x�E�t�z3��2�<���z���z��W�&��U��'Ϩ��g���mO�� 'Fc��=+�V@�|io��5�jw�����:�{9f�>�/�{ԇq��G\W�؛~��K 9 i��/O�|D{��e�9F�c_f0*~���M���u�x���]����d�
�/w8�ê��i�����NշK���t�� V�1�y㳟
��:� ��fnβ;�ы��\��o0�逰����t��K;xV�=݈s�|�n��w>Bf.�u@��S��b=��rǢ�;^9�����h>��@�Ug�[��,\B�-M�H~�+�[�/2N~�����}�<�D-�Q�m_��{��O�zg|O����<Hss�;
d��늮�Le8�tw{Mn�s�3��gg@o~39���I���5w&/�߬ɷ���|�F�zE�����-g3u�szǕ�>�=a/@��巢|}��e�]Ua�����^?P�����;�@�c��탆����#�}g�Q��O�T6c�p'tø�V���{��cE^�[ʫ�m��j5�g���Yyg|8�SCgg�?M��ܡ���v#�v��eyIú_��hŏ8�Ǯ���9)���U]��O����UxJ��f���B}��hC�;��Q,;3��^�?+|��k����p=|�K�^ d�V���{n9b��X��S�!�;L�����ɛ��n����/+�W��ttJ#�F/�k���x�ȗI��O����1q��H�]y,��s��u�[��%�C*�<.�|��9��#�1� �k>�
������RQ���J��Ld �K�m����%R��;r���s�ln��0
�!,�a��[�ĝ\.�9u"��k:v��@�|h���;�<x�
~=�uc�@�/9��su�G����O*t)��|־����f���|�����h���g�ܹ��JD�L�e�V�e�imR>��(� �c�e#uS��<�8�z�/p�x����ǵh�K���w�����i�ږXD��f:�ʡ�-���P^.�TW�����U3�ϣ�B�����ռ'Ϗ��/Og����j��U��:vK� 澓�L�x�W�6�^�/Ԯ�r�9����}늷N�8�w�q����W�{}r6�ul���T'���������׻W9j��ҹR�@��� ==�:�z�1����;��{I��Q;�G��ƃ��d�z��Mu���tG�����)�����|B޲j�q�+>9���<j6E������D�v�Hf��Ez%MzMÙ#������}��2ɭ�c���d1i����>y{Z�\n���Ԗ���)z<n4
�8ˁI����#��쨯��n��/�j������w^�Y����u����|��>��M�_���f��w�nG�d̫��4�{��2�iPӼ�n���m��U���>���>�7w�5�����]xOg�t:�z�����hC���e��LA�y��^:��m9�^<op5[��+�m���Ƣ4~�E��G{��U��/a�Νj/�ZY{|�w(��Z�W1p���04�n	�����w����F�Tx��.���`K�s1����K�g\ �*�S�q>�-J�c�c�J�V�Y�٫�'[��\�s�^��'M����뇒����N���W��߫p�{��ic������*����u�7Uz��X^
tt���b�Y;p���ǂ�t��2_�|r=顽���<��8�95��s���g�:N홏e@��Y5�✁�p6�]�E�J��@�u��k�{��/�w�5�3���)���k}t�%.��<4g��e� 5cj�������g}��n=�\�{w4O�)�Z�Ϣ�hx,�{h_�Ϯ���(�}%�PeT9��p9?*)�,�]�O�V)��e�?@}^Ñ�����\?)��^R}�d��(Q<�*�Y~\:}��f,��ír�WsSޟ�[1�*v����&��T��'��Ͻ�|{ڪ�Nx��ˀkTJ���uZ�verc�����}�Kx�E[�hh�o�m�):UǷ����a����KI>�]{��%^�}���� Q�^SY����z�팏N��v�{Ը���?j��}#/���ki�^���+�\U����D( p��]F���r�������ݺn=B>��}p4�0�#�y���4+,4J��J2d:���x�sh�yЫ�W��a�8VWH�nF¯[-�9c�2p�������ʕۮnGdR�|��x�z��OF��d8�q�D��9̰�r�q����}�))������ftq6���.=Y�s3Ꝅd�����W���j�ڇ㑋z��s[Gǵ���xpz/�;Rn!�ԁ�}�^ w���~��6��1q
d�H�C%�h��lcA�E��_]�Z��%�9G�����w�]��_�������j��z��_/VS��7>
-��3Vn��to���$����*��ziu���^����^�g�����Co�CL��o7{Ǎmyo+��z���j�mhW+N��N�����/n�1�W�##_�w�"7�^2�+"��/Y>�Wv�CݟEG����|N홆�N�VW��9�v��~��u���ނ~�o����?LQ>{7?sy�q�Oج�j�}z�0��}P��ʭ7�:�J ?m�j,z&nm�����ie��g�G��M�>��{'G(^�B�|먬���P��e�=P��(�r ��+*��s�wkV�p/�⥅p7�BN����P�S�+����b��QC"ԒUL��'6��1oN]{�η'�/Tι��!znMx��L{E�����^wX]j7�q�D(p�[?#6�Y~7�L�"-�GX-�cTo�cj�;\�8���s��8����m���朙	�,N�%=�=��,Z�͉�D�����s�{�r��2�aۥ-	��]�e �{��Wj����[�0ľ
����m�����m���v���X��7��P(�T�����s�&��}����=,c�Q����w�y��[�������
v�c0���ߊ$�3�L@)(�[72��Cǚ(_Ο�FB�W�Q�׍hm��Cr7���u~4o���t�W�<��>,	����J�U�&���ݒ{�V�{����Ɨ�3��w�ԇy�Qu�&���}6��j	d�P(��,��J��4�u�κ�9�y_�,�w
�p��l�zgx��c�ՠ��������ֺ��Ū�����MC�^��t%wz���F��¤��W�B��W�>��'��g|O���)��ċ��W���L��KY�;�Ϻ#_����OKF���5�F��]ޢ�������6�>���f�b�5&����ړ�.7�f� v\�+���=�[X7�s�5����x����#�#�������vn��,< ߡ�"���m@��d���N�q^�Ƒ�?E���^����=���Oٸ���׋#)�>��Pfn3�a�O�dj��з�?�l�}��p���i�u��6�.�g�iv3����܊��q���}���a�M�#�ܺ��R-�U�T%֎�����(��WA�	n�Ή೴�w�RS82҄�f����c��!8�n!�@��}hV���1���ܣc���R��S_f
�K�uof]Ӕ"���K�o{7�>�^�>�zN7^��	Y�����w!N��ne�:�l�P}�?Ofz�w8僽�}���pv}��q�sK��~��^�To(U�k�jx<'n���G�Ù�~z�_(����eqR�迫��;>X�p*����L�����=��b��#A3>�˜���޳V��>��ݙc >S>F��rW�١�w W�Y��V{��T�x�;��:Y�cOP�q�MmS>��*�3F�ʦ.*e#qS�����_@�z�;=~��{e�*�u.��Ӟ�����l{�DK�A�d�=�$�3 yL<�-���Ax�.�c��;�VVy.���S�K�ޑ�=�=�{UH��/�N�w�sRxn`Ws��蕙�ɼFk�5"��:� �g���qV��G!���{�t�o�Fz����T'����U��{�ǜ3�t���<|��YP(JX��͝���c#ӽ~gc�=�����'�=w~4*b���Os�r����]��$�Q'ҏ�I���jh]9��|-�!�6����O���L�w!ҩ��ƫ�:����Tz�|2�N�.���2/+�`����U�j��yա��9��U�3����On9\����#8�%�ã/�s�E���"�7�X�R��]::G�Xޤg}|���A��9���Y!Y#�Y,�&��哣�p<�z��sJM!��OY��}FCY5��z!r��M]�wc�:1��>���E���r���'����x�hї�{/�P#��ʊ�_V��/�kfI{�j`��Y4��b��Ŧ���4���{������q�C3Co��m��:əV�����w^���|'��1r�k:s7��nSXrϸ�5����I�i����z��{#޺�#&kz|
5���W��L쮺+����H�c�l���}R��7|�E���ȕ5�0ߢw����	Y��}���sƴ��m�ޅ��0�������:���tmz|N��`U�G�r�p�^���Fl�N	'h��_����i��~�m��'v��{*�E���kM�N@��v���/d	��7~v����z�/�%Y^kg}J�o~�B�|���8JVf�=P���R7N@j��"��;M���^���tπ��SNko�ǞW��/m~}tE�$�CD0�q������|�5w�r>P.ϡuSz��"=�|}���9^u�^� t�p�O ��ڷ}�y�d�N���Kw��/9#���u��,��ⱔ>w�h|A�u`X0���t��	�{���[M���T]/+���'6�w(��k�ʶ`36N{'`
��Yٔ.N��Y�ub����Wiԡ�W]�n�@V�i6%�֨k�d���:��6t�qe��nII13�@��wu�j�����j����|�0y�;�Q�� �rEt���kj�4m��F�2��G
v��a���,)� v��y8�h�����t ,��{��A�*��5�%k�\;4�6�.���Q�ճy�ŧ�^�#]��х�<�}A�e�B���|힧���7d�kNՁ��a���]�"�䄪�H͙X�ڞ�w����k{�&z��a���!ga���fe��K0.��n���"�Kvo�J`����0�HR덵�!b��\�L�b�e��;D;zc�VU���쥔�3�ƥ6-��wa�{�����FK"��ƫ�WV�P	��[j�ڧ�ܨ���C߷6vu���Z+�x���Z��ёJ���o���h81��$�G��{�'��%��<t�-"_B�K�79fi�O��6��	�6��BRl�ʙO��3�		������[]��![0��W(.J-�-���Z�P��*gQ�����-�u7.�jݷ���}2��V�S�8�:e"���1VMڃf����Lv�
�!���}���	����Nڏol���N�\�va��"��Z��t�i��v� �a=.�Y�嫧���B�|x�վ��S�t��]cK(�L���`㸆#xhp������ ����9dNH���v���iUŜ1��:��Ʊ7xm�١�/$��z�@<#{���Zo�	�s�F�ڼj�_�w'\�v�X��q��:��ܼ|�g'|)�b� .T^�����j/):W�I�Iܜ�f���5˸�b�q�^��pZ�����ud #gz�U��-&�;Џ�.X��w�����]l�3W"맟)���;=v���B^���t�o��5���(9 �K��f7������웰5�\Ѽ�d*�ִq�wx��������q,�S���P�>o3a�Ff���'y"�Ö��C)��o�r8Wh#���/tG��5��PX�q�C*�H�?X���_fS˻��{�ry�~۔�<Lq\�� ��)l�ISܺ��>s*�i�r��Ӯ5�ڟV�}+�n�|�h=�Q���d饻�}Es�A.�����Z�V��i�Ϯ��rM<�r�9N`�[� �c�mw>�����#�.�s���,�xVizݑ:��c����$|�r�B��/�d9e��}��5e������v�s�3A��YcT����Ԧ?�T���nĳ�u�\TεWu�ylk��|*v��Բ�F8������d��FVj.�u��1�.7ïo�^T���(I�A��zo냩.t�"���V��uz�8�ɼWBv�Ot�n�~����fc(�M5��5�$�&��a"�1&$��Pl�d24˺��w\#3&c!�(!D CRd6LN\�fF2DcD�1��)P���&	�F���b!�hEm(��A(�a��lc0��NnA�#�@
i$ 	 ��D�L(�)��X�� �2i��2��"bQ���B �)��T�D�S9]C��4�A��(�4����&)2D�\�AH��ى�LID��Tb7wb0d��4&��a %����!fh�A%bf@ �P�P |Q�Z�MN�6N�8P�]�e9���R��]�
��U����(^�8v0l����W1���.=��䢐�2��_<,�ɉWd���%l��T�]��U��"<���9����W����d���f}F��}7w��>UV�ǀw�(	�(�����~���n�����>.<��W����p��s�n�>�ҡHz}l���(ۂ`�� �@�=+�j�-�����y�9��]])�B��}��+���uz��oz���S��&e����8\��2g@�ioY��y���������\����h���J�O��tx��{��_�=�W��Sh�-�	 ����/��F,2L��M���yOy[�G�B��W���xİ�C5�S�_��uY꘵2|�����=ɟE���z�j��_{�{ꖎѸ�/Mw=��|���F9~&Mǽ����͎�"���ȯ��ޑT������nÎ6������W/M|����G/]���I��O�������g�Y��vϔYE�/w�I���GͦǕL%ckG���t]9�v�6P�^��c�vFk������A�������}�f�Vg=�?\P���˦xx��c܄�wY^�t�A��`	��u��c�W��7�}o�1^��^?l1mx\մ���̌E�b���5��=�;��N�W�m������J9@ǎ��sy�k,�ʝ��9v�Y�Dk������*�!X�F\r�Jט��S��/8�]'Z�)��D��xw<�,VVʃ�P����H����[�J����s���4=�v��.���=6�W��������5���Y��Jk���[�_���IV�z�,�h����>���׆�N��\��
7κ��3 ���>�P:��W�\���O��|9h�b26���
5�����߯���y\og�c�u�PϭI%Mz���z!叕����JC���EL�1u�	��>-D�@��Y~9��/�ey�yau�ߔz�e���Į�s�%n�:��X}����
G��U!qU>Nq��uo��3�z��t�i�.n���9�gos�:;����ږnD�_� $H��l�T�������ry�<k�{d�u�cW�����>�r�~�_������!:m��q��>6Ȁ���?��x��0��\g�o��3�w����gw�/=�O��=;^G�=�C������U1;?UO�� y�8����f��S7��\5-��û�0��[£���9��w��w�ՠ�{޾�=U�5n���p�KSկd���� x<�攩���@]Z*�[:6��o
�pڿI����'�#�;�}�ցP�Y�G�o��
53I-���ą�j�t�IzGKs:4
��|Z������΃Ts�h9�Rx�0B�-��O��v��n����}�ck�J��&���%&:W�	Q��u�3�;�-u��;R1њ�>�v�Hls.�v���nC�}J*��:��W���ǋ{�K��G�rDoTLeO��h]zV���z{�$>M]ɋ�߬ɷ���p<���O�竖�EǢ��
^�TTQ�.�=�*%��N}����j�0�9z�A͌�e���+^ԕnd�����\?dV���m@���l���a�z�M��ݑ�Ɗ��q�.<�=��Y��.Z����s�\wޑ�.3�a�NG�4:�{7(ft������ݨs��\��Y[�[E�f{�����C�`��ǯ�"US�[��q�	Y����V��r�h�!ʜ���[�:ʛ�⎟�T�ΟQl�l��-��DI������+}�����o�6���_
��l߄�|���$�	�῾'�P�R<�]�NG�����D%�^02]&VS���{D���e74�N�����}t�%.�3��<X���7NC*4����~��?��jC��y��~h΋w�z+������a��W���*�Ǒ��*����H�UO�y.��/�>~ǻI�\5wt��)��{�W����j�z�����χmK,"K�1�$�T;���uG�e_��n���yG�-��*�o �M+]��f,�@�*���*=���(o9ղ>���V|��!a�Y賃r��ʛ۳8���нqwe.9������Ŕ��̖�q�T�4.��g8evi9�5��{ҝ��]N�Y՜���IT��}�{qW�w�8�#�{7���{UHۇ�`��-�s�xA�E�ub��r�׳�8�,p=ϙ��������*�t�#�g|W�zN�~�\���ճV�T'�g�#��{cnn={�ٞ�*��ǃ6H��P*��B�|ioW���ٌ��_��L��~��'���Y�<@a�ᗚ�[ãצ��UT鿕IX�:�N{�r�Kz�}��c�ʏ�M�\E���X:�ϓ���;�j6/c���s^��!��b��z��kf�e�R�d0"d�@�WP�{���ynߕ��Y���z<�"}�|�C7�]@�^���p7��#�Y�߿�=�z��/C���<�>[�|17W&��~�=7��~���}�ہ^u�2�P|t��zv�n����l��󷻚�僽�}G�W����{~K�|s_�I���^�����z������Q^��WMuzpN<�=�E+Q~���w�VSqR��:�emCQ*k�c�Wx�o��%~�[�:�<^��_�UϚ/'�f��!vv�e�P6t;��������]L�+��{ g��{�o׏�:�{�Adٽ�n�Qm���1�)�c�7uP[�-,�q����c�@̾L�߷ ����~�f�p�.YV��7]�S�y|�V���#�+.Sk��
샓�u�R�rwOL��`�׷\�Н<%�88t-��[*�󩳻Xާths����v���*k{ۜ���7S�F=�ͺ�C:N���yP'ȱqY5�Yˠm0)k���t3�zzrмy���t^��]&��W���{��>�G,�)Y�xj�C��R2�0�N�U�������{^g�h~����MW��^�<}/m����Y��$�RZ5UCR{�絛׵aƟ�'qm$���{��z��^ w��}���{���W�x"�jN�w�	*o�~�[������BC�|5Tm�Ϝ��O�3�<��W�TyI�|r=�|{ڪ���||�\���\bW�=��LߨM�8 7FxEp���S���Z*�Ӵ4d7޶���'J���:���v@~���M���~�Ww�:=�>. ِ:~�[ TA�^SY ��}\<z�팃���{�[�c.����w����.&��z���W�)əe" 5_	����7E�����a��O�δ��y]�*�E�CM_�z}H�g���7�z��g�*��W�n�Z qϫ�q�Ӓ��귅�߼�5���>�9[1��rMW����� }��^ w������:��LZ�>R�{��I^���y�[�L�m���7Hx�FOk*����B��^�~���qz�㭗)����V]>+�O��xm�WxY,��Έ\���R�h]yhU���.b�D48��^�s�p�䥲�j$D/J��Vu���o��m���Ar���;�b}��)W
���v�������p�wro�&�=�P�f�m�w�iG��iWc<Տ*�]>�7,;�Ӂ\T�:%��WF�Һ���r���~����=>�z�o/[�&�/3�p{���*f��>%T��Z�O�迩Γ�(z�n�0��n/�� �Y�P��ĕ^d��ў3ލ��
��˦r8���c�D�s��!�;���߹�k��滔<�~���N�������)��*�{�ۡ�دhC���K�uc�l�߼�s]iU�����o���/�.�7�w������[�]EQ�P͙xm���]a�Z��=S��[w��+�ꙺ.��;>��k�r�}N�p�^Ey\oy��:�(	Z��Dzt{��������J��BgGI>SNBsp�k���@�{E�����+��ˍ�N�O���Z���h��Y���4�}jH*�3�L�X��T��T�9ǓAվ�xh�!�ck�C����Ld�Ǯ�3�q���7��]�վ1��g�D�_�&H�G�ٿ�e쇏6��]��Y��������Iwt���T՞ͷ5��)�:�^�7����@OOI�
<�eY-��徕ŖkE�����vL��ؖ�
/+Ӯ*���޽�.Hn�Wk��`�mp�x�0����+�*.��q�*��c:�I��q�7���vrW.�ﻖj�e�R�.�:L���p���K�yIë�HN����ǰv��� &l-���^*�ʨ�j�]��g��_�N^f�~�·Ey�X�C��#��!��g�Dt���~��K����8�'��'��y���U��/N�0��o
�ߩ��sKgޞ���_~���uU%��B��r<�F�k��>����HT��h/�o	��Cj�&���'�=3�'�ցhF"��P���G�f�^=��&�̑�c�����zV���z{�$>��ܘm�����W�ɕ�V�_��h{ S�x�lT'C�W���sPz�dK[z2��M_�,m.���n3')G?L�����~�՗X���GL���^��;ލ�|Jѳ��;�׫t�z}���̟+ro3�����j�E�=���UO��H񗞫zsޚ�yt/~��;_���ݨoݵ�x�Wz`y��e�=Hr���}R'M��x����dJ�zKs�.;�^���f��쭣��N�Qjdy��n�t�z�����YU��(�%;>�Q|�<A�:S�x�{*7�B��5zb͏{�I�G�r����,M<�tEs�[�Iօ`����5��xe�1�	\(^���'{���E�:�ܧ���j�j�ML��΋��4-8�t�V�Q�ˋ������x��[wG*H�u6X֥�ڙX�ݵ0M/��,�mr
�Sv��W3�g���w0߱#��U����Bg����NG������R^�� �L��v}��{�=޼���������1{��H��p���,e@3ŋ��#qNC*��,�� �G�н���+�=WZ�.��'���JG�^�<���b���׎E��1�hʦ/�H�UO�j<g�+�^�X�ם;˲��C��x3�'�;�D{��u��[�K�A��f�D�Pf:�*�x�7u?4�nϱ^mw5;�^�>���!g��;���<�_���o�j�o�~�9%��@	�V��HF�����i}�D�����2Zv)��ۧiNx�*=�:UǷ�#o�][5b��U2�w��/v�j+�%�}�!�X�?J��Qz�7>��8��_��:Gۺj6k��{!�h=�3��^�(��߂���F֒G�ā�9��Y�wf�RV��fH���9�-�7��w�J'8������z�3�;
d��OY��_W��Qkf�e�VђIZ櫽�ջ~�Ň<E|ӻ�����ǌ��|�ƀ�P��E|��#ʂ�w~;Ɵ/Md�@t`��뜿Ф��d���%��PS�0��[�=����շ�u���
��ڼ+;���:�����M�
�c#%y}+�\9�>�!�4t���MwN�i)yY�.�67f���\�����]����7Q�;�JB���E�-}�k?r���;MGr�curq�@��z�d346�p*<�&eX6���{��f�q��ʟ�����~��1��%A�5�5��Ĳ������=u�=��]��3w�BNk[�y_PJǬ>78:�Ύ��cn"��N��+Ưo�J������9�	\^����ڱ�;��W��C�������sƴ�㳷3�l�w�NQ�t��;.�E�G�K��r3�ѫ۴�w�z罺}�47�լ�m�gI��@�"��;N@����ߌ<�5�^�e�� Aֺ�z}^~�����s��B�7Ϯ�ȋ8JVfza�z�msI��p���9���Y�_����w�o�
�Z�{�[����R��oϮ�ϮQ%�-|�������y4�zk��X�T�TF>E@^7�������>>�uC�K�����x:vK�=��J	�؜��a�U6���J�L�$'P��^���Rg!�К����R|_�I�������;��U�un��f�vΏ[+�Ή�� �<�(��]L��v�s�hh�����B�O��+c��H	��9��Ìl>�x+��`*��^ �j�"�fݠ�ў>*����qo�����XU��W�T�d#n#3�k��V�j��'0u�\��ۏ)I�J�C�tWs���*ڼ&r*\W�늰��ցx�9�d	��BXݮ��'e����������mO�Âtd���J����[���6v^��׼�^��Ts�����^��N���Ը��z��]�✙�P/���J�u���f��T�ֺ�n��v��ї�]�C�tÏO�������z���g�*�Uz�ђZ7����Nq�Vz9�$��To!��Q�;WP�W!0����G��@�#Ƽ �d3Z|���nVz������뜫{�ete�F��'z�U�S��q���m���ܛ��'��bdefĖ�g�ѣ[H�>������-���A�A\����E���/��ˇ���|c#_��&�/�� �}���ڵa�~�롷	��6n>��Q�ѵ��T�N��:N�CՕVɝQ�!�L&�s}/k^㗹���=��s��Mx��TH��˦r#��ݳ1�_	�0�'�z>�:ؼ�U�5Q�A��U�Wv�� =������A�n�ޜ��4=�w���ͺ��Iݸ3A�}�����Q�f流����w����w�6� ��kVEįR���|�c���{��:�*���W���,~g�<K
�LSO�Mte��G��Ѩ�q��L��U����U AW��fj�o4\�ZVU"�	Sh�]��"u�2+8\ᓷ�{C�õ4�LN�6X���:�fL	S�y���q���lأ�Ak�!>;;�0�֜x���Άqd�:m_:�t�����������w��fݜw�L;�:@rg�YF�L}��Ju��w��9���7���h����o��b�M$s��jC����+X��F��5��d�̖9�c UC�j=��Vu��\�N�і�3�m�\�9�%��������z��ǈ��N��S��>��B���b�tH�Km��a����I� 4����w��h�\���C\�����c�������y��]�����u����P��m|@�|����{��
R��}�n�m���e���u`��h˄�/�.)N@�Պ���,����i�x�wLkK]��y���us����*�3@�bt��Ԇ��/����j��Y�8;Q1S)w��P6륚�Y61.ODG+rX����7����j�S:(
�Y�g!lK�d��*W�o�㛦\q⥰�Fi@@���`	�9&V y9�W@i�'��E�fth]vp��dm��1(�+sv���1:M�}�:ݤ�+�I*ԩ�['V�v�i�mwpn�@a���f��	V��9Y
�Ed�ζ�Y���ɕLT۸i�(�#:�n�ܫt��г ����Ѵ4u��pMupܽN���o]t�uݗv��_Q�OI��j	����!�Bi�|�Ib�cN��կ#�qy�";���Q*٧pVM�x�	]íp��՘!|)���㏭+&��p;�s��Ru��z�IzM^g5�W�`���� �X��1�5���r#�>�G� ����:Xb�;^��mp�|�5*Cs�Y]D:��뗛�A��5/�t�]�L9z�P�L�ٛr������t�#hDӬ�k���㷣E:��q@���؋t��d-�#�S���a�}7i���k��f&'WK��G.�6z��ύ��x_R]�e�O�ޜe@��/;�)���=���0�v�wuיr��y;d��� �+�����U]>���
黢S��BS���]S��ŕ�:��p�|i�Ky3ǻ�
@�7]m�����3��'��\�	����eS�5du*��j���f"�cx�MƺԹ��2��y7�˹t�.�9�u��Vw-4:+�Ĺ��J�/�-eZ�Ά�8Đ��w� �#>铸)&�§T�#S;�'{�JG���yb*�l�Q�Z{�4^�m�,ֺ���`u�cN2hP�����<)S��G`7�5��]7�s�,eŶjX�U�ϫ�����\\s*���z.��].Q�oP��|)We�e��1QK� �8ҧ�>*pwsrNWaW�2p"����fn�]������`~B���,E�Ɣ���Szd���(�wtd�����ab�
MY� Ғ($QbđH�9�����llBY'�WPI�q�&)EDTXf�jB2i!6&TQAIL3 &cƈ�`@m�wtD����N�!�B6I-%�$^u���&�Q���\Cn�u3!�n��s2(64Y����T0�8�x홌�cE����r(�F�QF7+��� 
����E�ӝ%�N��"1"yۤ���#i�PE
c��P�&��1�!"�o�B-�0Ƽ�,A@Z#H����:�x�J�[&1�l,��v^;1�ы3�J�� ĤB4Q���������wh����k\����]ѷ&�5A$�=G��l�`]��DFb +br��2��c�qJU����v%�o�~�?�ʨWJ����4nϠ+�����/V����������>����)غ=^�qy\կU=nI,�|&xz���)��!9��^/ w�C�,������xf�F!6\�g�:xw���վ>�׊�$_�&�,_�*�����s�&��}���goLx��e�I��o.��9��|�z���{���gö����Iux	"EKf�P^�D�qG;g���;�˷m��SW�#���+�N�O	½N��v��� &l�����{��a�y���q�e��Y��	��[t� �O���!����Qq^�bo���� �\�̽���'nk%���Ɵʁ_@)�L>+xL>��m��L�x���=�z�LߍC�Jٍ�U>|Q�˥�ziD�d��Τ�$���!WR���ǖ�vڿI�z|�������E[�k��Ω��彳Kw���X��#�K�Rn�GM�=�B��J�W/Mwz�w�&����ߴ���^�C;��ݞ�w�5�2R=_�ƣb��� /\����y\	�1R�ތ���Mic=�<�v�p�Dхg@�6,i�)�(	��(�����e�杫 ^��
��|�;7��gwB$�+�b�߇v'�\�}�F/�ҡ�3�޷�کG�)�v�vN��jԗį<6V�m�;���K����S�K}I��vnowh��p4fZ��]�شϬX�N�F{�=3��/dV���m@������}�z�O����~��c��ԙ{���Ƚ�G��4T^�Zʩ��~��7�z�9�����:��"�4���`��1�B/Y���Q۔�g�x�(�'N�x�E���T��z����UxJϷݚ�r�t�%�[��c�����`,��w:=93�`{ģG%��[�q�̯�V��{*7�Y�Y���s!���\�ۺ]a��a�����xNٟ�x,���򑅁ю���g�_�J�ڕC浙�V� ��i��k0�Ϯ��d���,I>Gi�eX١�k!P{{��7s���2�>��B���~++ԇ�Au���Ϯ�r�$��3F��b�*e#]�FןZ�����/~�w#?��WR��߽x3�'�;��#�~���9/i����%��tc�*<N����6��RڿGz��n�P^9�Ƿp�ߴ�y����P�{UHۇ�d��ϔh⑻��f��]b����I@G����x�!����)çi�������{}r7����Mk��݊s0OG^��ј��s0"��X�n"�*@=<:�;�WQͣu�śS+�ov����7ť|�6����3�$�S�V8�̡�:�ImV��� ����7i�N]c	�+}
]��ϐ42l!gd���*U��c�o_v�vt��+oN�HZ}lס��(��E�L�������
���py�m����_��~��٧��@�v��j��VO�����f��Ϊ���RCW@�yM�=�<-�!�,��Q�gXp�8��k],�^c��ҕ�������5��������~�gX�Gڿ ��aJ�5>���r���W��W�n��T�m׉�G���D3q�T?F\�Q�dy��TO�M��:�w�ܣy��}E���
ו��M�ɸ���~��>`����p<��e{������e��ݻҕ�x-�8�:�7}��r#��{WP�/]�����o=u�=��]�̩�<E�~'��yB7����B��9,+����Y^u/I�q�x�^�\<�S^�ߢ��mf�F���e�yx��gz��~��C���ZX�rs�P6t99'D���Q��W�Y.���0}]Rs7��ŷ�S����9�C{]o�(�f�q�gIݸ3 �&��ا y+{ ��"�Ϋ����^�}���]hs�/d�]y�^׫���PQ�}t�E�%+�0���z���5Y+Χn���Cjn�f��X�ϭ��3�¦[��F�O��u�N��w�ȕ�ɭ��8��Ր�~*��|9T�w2�[\{�E�5f\)���?��W_�՘���ܹ��m��Wy�v�J���H�ԻoE�Qn���X���kޱL��[.}�����{�A��%�ӥΗ?&1�;|6�x,����Z�{�U�c���C�dK�Bߟ]�r�(�ZoΧL�;7����y�,����Ute#Qp6����;��9�����\?)�9���,J_�uoW`�{�=S~�7�K�S<�������O�2�ȝZ��9R|_q>.��5<����Ӳ	s�M�C�pr�ӢY����P; ���%?O}h��N��}�nX�p���W��g��'J{��US0������	�\��J��X���yto���V��	5����grܿh���5~9��=�\N{�ODz��:��n� p��J�[qsh��ͮ����[�ۇw�	������ߝ����"}�xΏq�z��V{"����Q�Z=鎵qus
�<g2X�y.t���][F�v���5��*���o�� }�5�{"����xܼC�,���eh:��OM(�M�Ǿ�܎4�pWT��hޗ����wrq��d���@w�@{`ϖz;�M���ur����F�����A��V:pzJӃi�xU���P����/]���A���T|qc�5R��\�}��9t��]-��	��m��qh�QW{W����r�i��=�j�%ի�o7H�%tW&���s�}���Ov��! �+�gJ�T�V�)���W�^!����.���.�S����d&��:�]փw�XUs�)��K��[y�c�'�����Cn;�4͞%pɆ�ևT�N��s�����{��-פ�Qu���bF^n�ddo�C�9��񕑾��P�yt�G�pf<��wY^��cW���z���˽�R��^�o% =X��*]`-ϵϣ�4=�v��.��OM��`7�2��R`�Q�߂�̛9Z�y���z+���2U��`
ZՑq+ԼAs����tw=���:�+(��;Ռ;�ڽS�U~��%����Pgj=*e����n>;>��k�*t�}[��������f�~���ҝ�M�Ǽ�u2ԒUDL�('��|�:)�N_�k�ި��/Ǻxv���b��n�$��D�&�r�����U����	�ȱu*��>Ny��u��yo{�D�$���V���86:X�{������ݑ��ǰvԲ�$�3�H)�d�Wtwk�o�֯1os��=�y��ǩ��d/uy���GO\{i	�o��`��D��@����n��$tǮ�T�r>�<���.�Ǹ�-�\S���k����RN{�FϪ���S��O��{nẗ́kB�%�� �G�
��e��Gw!Bk	���f�NA���evu���]��q���^�v_~y�)]��G���[���Ni]��u�H�81�K�Z3�ܕޕnQ����O�	
6�8#������8]���m��6���S�Wl�J> s���T
�|��ⷄ�[g#�;��;����h��.��^�z�^ͩ�ãצ�
����T�� ;�!R_� ��[¡�6��}��O�gV��>V_;�w�GC�'P��/V2E�/+�n�\v�g�~�������?~Um6���X���Z���y�|�Ǿ�J̛����|�F�zE��}G���+�b���ϰ׫�zM�*|�++,r/ж��7w"����n=����'�z6�WO�UfX��8(a1�l���#ݹ�������>��Wt���o-�J��u�G���X��������ܡ���w�/�)�	��]�=�˵��V��1��0�YMIú_��u1Ҫ����xw�zg�yo�4c�Y$�g7]Z��^Vz���:t�g ��M�^%9.-��}.ix��/վ+,P�7ab����ϵ�`>��C��7�5�2���ۤ�1��믚�΅�?r�Ge��]@��ղ]^��)L���w�f��F�z�*}�ޏz���=�EY�R�,e@3ŉ'��S��{w������
����f�)n"�� 
�Ň�l��V���,���Sۏ���S9eqq]�ط��>!�x�]ȯ���,�t�a߆o;)m�9�����k���5ەz��'���}��u!w��r_f<�������;:�)���:���4G
��]ݷ��ڳ=�_�����)}�S�Y�W� ���^>��*��yT�����X����{���Ot�*���|��x8�z�(�	�����j�z������ɖX�Kn,���s���zuBC��<qTmџ3qS>	�o*+�t��s�O��}��=��ڪF�?]�z���Ur*s#�wP�q]{�b�Ro�� ܑ�Cs`z[2zz��n��q�����+P�
���^yA�IuO�_T��z�O��8!Ha��_�҅@|yoW���ق��Y�����ѵ��}�;A�_C��&�~������h_Ϊ��$�����+�1?)��P?�'��c���v^��M�;}��E��hxgޟ+>9���ƣ`S�z�\פ�Hjю���3�^@��S�X�}00s��I���>�ɯt�t�Y&��sn�O���/���*�./e�����#�s}�F-�OfG��7�ɿAޝ��<����{M.�߆Bn�M�?P��޿������m��Oǅ���2�˥z)*�陞�@6#M�*s}E��^�\4�U��'ў����S~�׃�eT��|V��V�.Y�����[Wu�ڄ%�����]�<�8 RdΑ�7}�S�b��Y��iQ��A|�_���p׫�s+J�xvm��s��t::��W�鵔�tey��L�F�M��ɮ����s!�O���N��s���eס�y����v�`qF�&�_5��{���l��B��|rXWgC��ةzN��߂x�ץ+�
�o!$�F�+�������*����i��R�~����9�Zr�vv�����r���S��],c	�dz<N�U���]��L���J��O�{��M��}��o�n���Γ�pfP�"��VMi�Xa����e综�5�/==^�o�.S^�.��.}63O{�H^���9g	HvM¸�0x�-l_���W/j���Ez�S7�+����]K]/zko�ǜ�����8~}t��mؒL����ޚ�Q�$�F��.�_�F|���;�a��W��O��#�p��>�:�^�=�O��yO��7�΋����d����S<yL<��[���Rg!�КZ��>D��)v�O71��	#�}u~6owj;|}[��:%���:�<�(��I)�y�~��%v�{˳��	�=�r�#�Rt��o�'}ULÏdϋ��� t���=+�jg���g�(m�o�&�1r��=���W���zw�ö=�\M������TVé�f�����>���r~�J,]_`���V"���uHGZQ��c"��� �z�{�-=�jk
5�1�1X ,Yz�盦���%k���=����d3�G���#���C��=��. @}�i
|�-�����݀0��p(�ӈN¤1k|nP�.^U�-�\�n�x��k����oa\7�lg�ԉ�G���7�����g�*�Uz�p4r@l�����j͟I:Ϣ	 ��J��2j2���Ba�&��n=�R���x��k@��U��2�$���7�ʫ=Sd�6zlT��u/�hޗ����p��f��%,>�[S~�"��U^[ZM�`Z�x���i	�S�7>
�N\EJӢ����W���_.��x�s���{���ϳ3���=3��'�����H��P�6o��U&�����>ӢY�rs��	B�V�M���_��G����O�3_�w�|g�yo�(S���<<3:Ǖ@��
P^�նw**�����9X�oE)@�π���>�N�����ϻ�Cܧc��F��fÝ'vs��
�6J���WiC���)T+�ʭ29��'���C��^#%׆�N��mpX�և������S�������z�w�Jw !��gUF��(u������x��u	�5�'�rU����/н��q�u�P�I(�9@�����r�}5��w��*�Sꪜ�s/fwq>�[��_f\
0�����ݧ.*к�3!�����f�A��cQ<��P�e����#��V2�Xɭ�+S��pB;�[{`����@�E�Sݴ��� q�-�7ɽߍ&�z{z{)�Ǔk��fa%Aa�pDwp�B� US��j]���Gp�������<���Q�}+�3����� �.�RS��cl)�3���g�}x�R�p�i[(c�,��q�Ȃ�|c�;jY�e]}�`�
�Р�0@�ާ�ƧrkՇ�S:�g�Et�z�|�8򣧽������ǣ�gǡ�=�%��Q�K��H��{�5�|r|����K}�n����:�=�C���z���S{[lǍP.�J�ݲ�Ez�ϣ��@nu���><��C�o���9��.==Z��~��;��>}��d��h�Ug�\:���*��M�C��Y�K�`?[¡����|.�3����%��_73%� Ͼs:��G�h�?Vx�K����L��rc>^S�b��]��ڽ���`��7'�ۼ��ob�l��4�����)�}���F�}ޡ��QQF=�Oa�������M���q�ڽ��kr�ن��6���1��HX�C�7�O�<�q8w�P+��l���.�9קj��t祖c}�:�2;Kގ�{yl%3�+_�x������x͹]�4mJ����iq�β���ԣ� �nV`�;E��ﱢ��>���z��=|�8�}���
��(!fg�Jh����Į�ҁ�EJ��8A0�	䍾��K��,�q�Yp
	�<�o�6����F*j�īn�(�_v]��Bd�T��Ϋ���ZPoT�+Ǧ�RmG7�e�Ǡ9֮�ʚzr5(#���Eg%4$rq�
N�����)'�[�wLbڣGEsN	�k�&�f�f�+q�[*죌��L<�/�&^{\�rQ�	|�W�LFmԍr�-N�Ҵz�u�V��
��-:��]�F��:%|,�6��Sa�ݗnC}���V��iHxb�����@y��}f���+֍�sȃ �!�w�w�I*�F����cX*ɽ۪1%o.��"�h�s��#@� �����ق��Jtl�LU��#j���H�X�g*���9�wX� 
ν��Ss��a{9v����B��2�?�౽:,ߛnj������6��-�eU*7�G�6���QD�ϕ�e#;Ӧ�Nppv\ݩ}��M�9W�q���֌�i��C:
�*A�d<EeZ�r��g/��1����̳b\��D/[<S�<��xt6��N���.�s8(�0>�Q��\�`�V>o�M�FZ���b���b�\��&eZ��'�.T�D�����Y��}��-Ur���x�v
7ʗ ��/�nm⮻����X�C�(�*��Ϣp���c��z��k��
&r��;�D�7Ѽl�@��H�).��F)�c�u���[��
v�GM0kE![5�U�ǷpZ�_:��;o�� �.(��ô��n��_q�G8����-툻;{i!֪��t�4���:�b���
v�"f���sqMӊ��f�qТ��^&�oyi�����O5u̵�
Eʔ�v�q-b�kS��E�r���D�(>R���]`}G���O�T�h=��ڳ��\�b֪x 7P=!�Y	��Z���ω���O�Gx�_vb�*�9��jcdۺ��$T�C �������\s��n�SO-�\��� �64{��|�BWNt��r�w��a==�SQ�[Ȝ����.Y�Tr��!��l`u� ��")*]��z�*�+Ȧq����r�)���&mh����k%�!w�|�PV��	��򎯅AՈۼ+�}QH���1O^�[�5���B���\!���!��tXHqv-�'��{t�MbA5�Y�L����U�lĜ�Cs �f�K=n*j�R�\��8���Ad9x�[Q9y�v���Q �����5��d�T7�;V^�NR[|/�������qw6��U�7�OXp�Th��C��k��r����:.t<={O9�uv4e��d�g:�:�	�,e�u��Mvi�0Z� �J�T�g^J��[mX�=�{(���S�Z�E+���X��m�{OjȺ�-�+��s;�L��}������|�����������%PElQ��r��w W+�"�CRy�DPD�X
4�s]�*R���"�]%)%#��] ���R�� �)���q�$	WwQ�����ni2$Tr�DRb�B���^wF�J5�u��$�L���Ib4X�wv�)"�Q�J(�.���7<��V�.WH�b��Q�1�`@k1hI# ��/ MbΝ؈K�fC��^w&�r��PQ�f��u�IΗu�DdM\�0�X��.4E<�@U@}H}T|@6�K�zn�-hZ�!9�6��Ga@��ID��	!Q�sqw���*��CS$J�S;��Ut�e�5%�z���(���T���?S"Ua%�6=?i�}ad��79<��US�s��ür;�^�����_/o�-V�o��{G��+h�D9�t헄x�y�eW��J7��p)o�ǲ%�/=v��w�����ks�.+%=Ӟon9dB��7�f�}�GN�%Ꭸ%[_��o�~�4�������;|�k�߲��Ϡ-t�����*_�3z=��b��>�G>�����.�|���r���ɣ�y��$�Q�
;ঃY����}~��S�Y^�<��.��~}u�eUA��=B{���{�;S�y�η'	'8�*��yty��z�g�O�w#�D{�޶=�>�{H<��Rͱx|v��^9��ѫ�o�|�7�3
�U
���P^<���\:w�9r|���������mk�u!����gEy��vO�� NjO!��C�ٺ2����*�;H��g|W�BY eU�=���W��w�/ƍ�#��#]Mx���P�pB.�d��@����B��_��\>�nJ{EϦ����ޚ����Z��;��������п�UK7�!�L���Ӟ��L��j���sS6;���>���9Р6�7\|�����(m�r��Ec�;�ن�e�����9ҳ�� *���TƯh:\�عZ��=�*���q�i]��j��*vla��!U�o��c|o{W �n���f�M���������J����/�+�ٔB��3�O�������5���Y�I�2CPz�i���ߙS���ڣyO�����iA��dx\&��[n�O��|y��_�.B�_��������z�q�]�d+�9��d6r��MB�m�d&���c��z�g����=r:{2Mԏ/���+�=kʿ���l����z�M�E���/M}{yp��V�����s�%5�;�9Z�y��"�{���_��6f�:|
5'�\|6t;���ۊ���мk+jŎ
s��ģ/k��{s0�>1��W3��������sƴ�?�Γ�-����NQ�t��;5R�՗*2zo:����l� �yj�c'Խ�2_�|}�#7��x��o�n��C:N���yP'Ȱ+ܟ�}qF��m��pX;٧�[ .���*!k�����\��T�lf�G�Ԇ��R*�����q��u�Cz:OJ���s|�ь���UH�W��mP�X5��������1��C���<���o����!=r��O�/\�K5���A�Q�3�n(�	�}T��ޯa�t�nD{���u7�U�۸}�~��}&B��E)���[�lf�v�\li?j�����Cw*u��*^k4���k��\�|���n�i��z����O��d�t�K���ڃ��W+��}Y�L6�T���X\k:<���Ζ'j92M=��o�u
�|�'�f�{��Z�-l�8�~��U/���j?�xWL�<���s>��D<��W�Z�o�R����y�%��Գ7��g�y�G�=���V��N�e�>���n�sJ~��^�<Eue��>��[���S�2����):W������y�S�n	�� ��r�;=�>��"sԯs�5,�.�&��<=K]�����=;������~�A��]��MK7�g��*��S�<sw�R�,5��n"�E�D	��oa_����R'�3���ޝ�Y슊�p�-�7�y~��Zi3��?��8^�	��G�Kz��n�!0�5~�q�z�>�� ;�ҳU�˳8�(팤��]\=`r�`����)��7��K��R_�Qߴ�5��x���������ص�nsW}���d��@w�<j���a�cԤQ���a��8=�=�
��zk�4��=7�-z�j��v��3^��CN�g��EzM���������CLٸ��U@Ɇ�և'�p9�=/�`��or��ڗd�׷xϒ���#}/}5�+>�\P��˦xx�΃1�:՘a+���%v�b��>���[��V��ٷ�eC�R%s��P֏#����^����:O�mK�pj��7s$YX�'by;z��Ώv��ʘ��ΣVI����L�ͦ��p$Ow<G�ub[m����5������|��;�cҫ���������Y�r�x�u��	��u�T��z!��zr;�Cܧ{ʴ\F�6�mFч^�z��!M.�*�t}��2��~���qG�%\@�`
��Y+ԼAs��^��{^��õ�t{�7�\�=7��7]EQ�P�}g��B�L��Qp<���@W]I:^>��l����*���^]�~�Þ�w���c�u�PȋRIU�L���I��r���׋���H����d�^���\CTt���~+"��<��G�J�L�֤���/�ȱu*�ԟFm�9��k�S�F|�'�{&�����C��纏�_���9�C���%�g�����@޼���,��ل�-������V��2�ʎ��������ǣ�g��H�&k��>z��b��~>T Ex��0���u�9j�_9��=��RM��{�G]�u��\��H˾;�ck�JS3��@sD�3��@�>ya�*��l�ޙ�>���'W�V��� ���IT�`��޾�=U�ә�,)%��@�~�+*_���QJ����3�,���<?o�8��3ӭ�,,w)qSk����5[����n��f�H��Vٙn{56,[[��i$�We���_߬�9HF*gp;��o
�mG��-��&7+����}��.PX�����16��k=�R�����>�}�K4W��y�D����>P�h�~$s�<I�ê�g�hmzV�^�t䙛��ʼ�j��>ֳƏ������o�d���{!����� T/ez��1�l�U'0���^z3��X����n{w�F�-o�{�r�֔3~]w��9z�E��L���+M��z6�TGO�R�k��w�^vͷ��R���+L9s�w�>��Φ4T^�[	L�J��3�����zhq�Y�\�7W�ܯ'�Ϥg��*�3~j/֨�@ pw����%����x�o�rc=��ͥ�x��gz�矻4_��[Gs�00�|s����+*���E-��o�ǍyB�L��;�%��=�����/�QZ�Q��׼o�����Ųt���\�O'�tK#�7�hG����n�6���_+ɵϳ=�{���I�׌�t�����W��.���L
� $ѝj�ASަ�%u������=�}]!��2<���
�Z�~��S�y�C�>.�~{T:(�'�ؼ���+�s{���Hz-�zpz�R7E����A��;޼���uG���c��K�A��4�U�j�*���);�Z2��z�\3>G���t�Fn��x&�n�l�`��?y��I�Q���6����=��ViW�:%����P�S�L�5'�$��g'��ͫ.w-Y{��������f����+_�S���i��S��T�;WAV��T��l�Œg�c`OǺ��FR7�L�/�㨚����#�O��F���lg�݃��Fu綧�w.�ý��;>j>�� w��`r����m�;ǫި�t����k�ս��SJ󇧎3��\=�����VͿN��"� %{ʅ	���=�G���� ���M��_�c�\��L6s	m�N��f���T�p�P�:~{����R�K(m�_����s٧} Ø��#�:�a������{��~�\UĹ�ID��X���lEs|+;9ϐ��肕m���_ѳ��+"*#�z�6�����5������<�W5s����b*�]B26{**"}ՠ�x�o�P��w����\��s�鸏z�ߟ9��q��n�Y:=B��m����*��4�{��7^����-��y	z{y,�NB�gcKo0��>nx~��w�l��O�F�91�����+��/Iӡx��wt��FώןS�Č�;���i���Ew�F���VG��£ߦ�k#����?��������y0�D��l�J�}�.*�qQ�L�)j��,y��Mؚ��ܫ(��1�3R0O3��94�!�I���QR^�u��%��9��ek�9�W}�R;}8�P"�\�:��[��T�ST�����8-K���I�л:�mX�4����l��v��Βs�Kv�d߾n�^���}.�p-�^��������}��ʡ��9��xǥ��]��5H�v^�v�E9�7P��Z�
�z�z%׼VD{Ճx�ԅ�]!��۟�䄉�d��<��=�z���Tz⺫�Ґ<��x+�k�*t�魿Ss�B6~�A�����*�&���k�-4�{���Y��$�Q'Ȃaܙ��*#.��qޟi>.�B�;oz@��2�wf��ո�ɝ��ޟm�p�vK�(Q<�*�$�3��qdИ�J�w�_�͖�^���Ųx��l��������/�N�f��3�B(�|��a�D= �����r�w�g�ϣ�Ղ��J�џ'޶��8uG����S0����p O��{nd�6�5̪�]=E��- z�75��u-���rա�w����R�sި:z#�uK�R��
}�s�����E��@bO�\�\z�oa\7�lg�{���:<M��z�is��v�l_u�P���y�Y�*��_B2K�d�u��FC�a��h�o�m_�߽�@�E��f�Nn�)U�^m��s/���S������~
��֋�&���!�_�/��;R��֣ͫ|u�cy���͝���3E��,�'P@�2���*��n�؉��ty���+�}9�L�T��)Ia���K�<#��>�F��N�1­��kot%��`��xցK�l3~��I�0��[^qR�v������C��Ʌ�����Iou���'��)&߽@w��ֹ��!�w���F���B,�^�
��gJ�/�Mzk��\��Ϣ�\rn�E�D�>���\{�Co�CL�%l�}ckC�o���X���f�\>X<����<=Q{w���J���k��Mx�dG�qB��.���royL���ٻ���j=�%a�9+�E)�v�j<+=��D�w���׻ӑޚG"7�X/Z>���
��5T���������u�M�a���OX�@
�o���W�x��^�>�����ׯn�w=������7�$�9�PۙxA酕��W�\q����u�T͵],���]�Qx�ܷsD��^�U�������Q�]E
K�<�L�L\E9��F��z�=����f>���@{%����{��G��*���Zi�����1��>E���6�ǇK���y��)Y5��語~�Y4=p����=>����y�{����J7�%y�}�ٯ�"�}[U���א�8F �!��^������+��ා�ͣ�����:�-w�yq��ݽb'}�gpu��Mv���w+�j���/�ND���j2�����V%9���W-�́"�Z���5���T�,�k��f�ß4�w!��ٽ�13�W���H{����};>f����O<�A��`���=���m!:m��q��g�.:7���(�B��@@H���GҼV\��K}�n��1�ב�zc8��$��1�L{ǥ�z�cO�Lr��Wz&��UO��:H��
���Bިv߭�]zr���a��~��ۋ;V,��7��7Q�f٥32P�*�Ԁg�=<&�V�Ȁ_��oyJ��w��E��{u�v�6=条?O�>9���ƴ
~���&��X�R�hz��t�����]+O�Nve��N�]ʈi��1����o���f�a�E��}G�G�j���P��.�Z˜1��עx�5�1���1��w"������z|Z��i��m@�y�"��O�����O�=aw�N�U*���۲������~��/��X����uX����W��-�t/�[r-��F��C���/	Áx�^�ZL�
��s�L��+u=J�._��ꐕ����s�s�3�`�|�����~�s,�4>iS�"RN��KM5
��֥xJW��Z�6.��9�^\�|3F<d�^,�8p�\��%77��YZ�$��^�mf�-��^÷��Z76��k �qGS_WY)�ka��ސgVd���}6�\�U����w>�ø#��Lޣi;aWP�7���6�D������p���|VǽQ��׼w��-��nf.<x,���tT{���}���+ԍ1y>�倷�Rv�`dK��Ȋ~��ȏz�ED��ֈ�u��+�3�3�W`�-��<�sԌz"\�2��]f��k���_��{��^W�,��Q��AS�LT2]+��uκ�T|�(�|e�O�أ����<��^��'�;���\{�Ǒ_4.��O�]<f�#�݅�jY��Q&A��=�"��R��x�C�Q5��O�>s������̶+�;� ��U߀�>�ꍵ�`��-�s�xFDJFA�c�޸���^Gx�u��]���1���G�9�q~'(���mǮ���|\Ÿ��7P*��s��R����I]v}W��_��nKˤ�x�z�3ޝ�n=�\Oz��h9��T"U@�nz*5zh�b9��<lo!��hz+g�܈:{6�W	;�c=>V||Nx��z�`?_�+b\ׄ�E�C�STC�lxPxC:����5q�{zȊ���Q	*d�zF�*ֵ���Zֵ�����km��kZ�۵�k[o��Zֶ���kZ��kZ��Zֵ�����km�浭km��kZ�����k[o�ֵ��kZֶߚ��km�:ֵ���kZֶ��kZ�ҵ�km�Zֵ����ֵ��km���
�2��j��.� ���9�>�N�� EH
�PUA*�*�BT(*$QU("$�$A% ��
T�H��JQU$(���(�RTTRt�*+cI"�U֔���v5P�UR�PYb%R�h}j�P	D�QD���={����UB@
��
��OZ�9��PS�
��T�AJ�J�H�J�(%T�RD(
J��@�4ҩAEQUT�2D�TEEE"��D�	UBm��J�ER}e\   c����vm&v���j�"�r�
�A�0��(�T:��q�U��%�u�j& U����9�G���H)))B%�   X�/�A�*���u[�����=⻀
  QE�GQ@P�(î��(�(��F�(��q�QEQEE���@P g5qEQEn�RG�!(�R$��   j��k��P�S�� 8f��USuLQE3�W]U9s�:�ZӦ �����T�.�v�1R�j��T�DRREEG�O�  o��ӶT�����]�ܤ��U�U��q�۪�vն�sk�wv���U*U[���g3eR�ctv��6�ݭ;K�<*^����t;m�
V�wT*��AB'�d�=�   >�.��u���+�j��7[���kiZʷI��K�mSu&t�.R��cu�L�ݻ��͎��wr���tn]mw��X��GN��nlk��3.�j��lĩR/�!J���^�   1�7��ӆ�[F����-;�ɶ�*�J��N�k���sv��.��ݸ�t���iV�s��횝ʭ�)��:�հ�٭��V��t�p��5�D�H���J�$�>�7o� ���N9����v뮴���*�r��t�.7SU�Km��i�E�U�V�m�����ˎ��i��*�Zʻn�w�z�{wP�ɝ���۶�ݹ�$j��5�JV�  ��tr����m���ke��핻vӭ��ejѨ\pۺwf���ݻww]�Vֺ��eV�UKW;�����T�#���lm�vuVu �kt�u�*�)J%vj���x  =ǽt���Ԝ9�峭����wl�ڴwj��ڲ�u����wt;m��FW[]cm�\�[l�V�6��nݷv�\���[�V[Z�:i*�:R�٠UN��U*Ex  ��T�������R�۱r��
��v[���v��wl�m���w����u�U�5Ϊ�˷SS���Z��n�ܴ8V�SA�
�OF�*J�L���$�*4  T�T��O�CF�E?�S��  5O�LʩP   �JMOTHA���ʯWu����t�k�[�oF���;7t�\#�7q��~��o_8���Y�`IN����$��HHHB�� �$����$HB!!��N������c������M�;����w��gH�zVC�����U�6�ʷ�F\�*�q=Tp��^��C&�Fɭ5s5i�Ԣ�+s�h�#Ӥ7��	r]�m��'Ζ��岪RP'�Q9�[�ۢ���It�a:�@�/)$ɹY2����e$�{cͬ�R�Ǘi�{N��^�q$*�B�E-��k{N�j��$N�Ui��6�ܚ�k�@AZL'D�z�؛i�ٸ���:�Uǲ�b�`4'�f���7+-����X��2fǫ����L�������D޽Q�nH�#7J�%n��؁�.�Y�1�Y�eh"�E4�m;-8�������;%d�	J��S+V��Ţn�	?��2��q �^
�eb��Y�̰�����n�C����vѸ�:�'&3�U����n`QX�Z�ʡ��6�D�b�^h�B��j��IJ ��6E���36�u���e)��j�C��p�;7Ou<��	;�ՁZq,6��W�iÊ��0_�Mh9R�SZ~WKS۩gmTJ��鐩�Ù�-�{�d@,��Y���t�P������5�/0����1+6&�v�9w0;���w��Xe���HP״�4D�4�#���m�4l\�5
�����J�1">3�CX�fM�U�0����!7wz�o6*	5+"[�٦n .��I�^K�p�J\B1P�Z%�E�)n�MQIwSmK�X�l�QG2��j��W�bx��j�г�]�ȫ�e�(Rp`��wv�h��(�ĕz�ML��5�#����Fm�(æJ�BAF2�A����mЌ+{<m�X����(��aR�r���Y����8�K�+N+���wL�V�A�`����6�)��
��4�hM�ST;�;�.Ö]����Ya�x26�f�Y�kGt��)�M�ĲȠ���h��v����/ 4k!B�0�*;�BT��������wB��f�M�8Q�棵 ��m8��kKcqc�)�
M`���a2!���$Ǜ��m=�U�x����.d��PU73^��%�8�+Tkq�L�� H 4�'4NGff푆���Wrb������E�u�3�o4ڀ�iV���i%
��`���.U��3��	L�Kq���2�u���"��4H�iV�j`�z��Ú	��b�����B[or!�M�a�sX���]%�D&���7��VҫR�<ʂ|]��ue̤�A���ҕv��$��o"6���㐷���)jr�x	u��M:M�#t1���:{P�cP_&�0<�
��uv̕��eFuT5����V#0��n�BSWMf٠#{Ij���n��AjM�^m+$@B�ݒ�ǵ�l�hfS J��{��36���lFBW��N��sJ�u�*5z��u��H����b���#[Q�YG1P�N�ɳ.Π2���!�h�4L��R�S�F`�V�RV]��R�+˶*�[�n�$V\7�2�a,���Sp�F�T����:�6m�IѢ��v �+����p-{Q�Rag��Ř蜶��Q���r����Ո�G�;6�w�e�M9�5�+2��)]CXp�)���V��Ѩ��J9�g��M��5o�ُ��aְ��y�D�L�3P ���N�M�TT��֔������=9��L���Ӵ1�)ͭ˦�W����O~ܘi&�F7h��҄7��-AaD���m�&�D<X� PA�F8^e��:;��yW�m�N�䶨�2ŗT����iWoh�3>�%��N�L�(8N!��]�D5��h]q]���0ܗ
w��Zl�	�]A��o��^4kC��^���g�7en�_8�ĴR�&��"�N���T-��j�܅L'ZU4;�CP�`�f�iKD�E�hdY�����a���醵�%V� BNc�� �a:�/.n4�8�$!or�mX�CrlX�e���˃Akj10V���ٷ��
"C�`$V�ÉH6���;3`Dj�.��DP�أ��-�ܻR���L=u��w���2�l�,���
�Y"NP��$Z��iV,�3�Vs&��{����t'��ک/��h�(�Ҵ�c^��m [̗��BK�,��մ0SM��HZ�݌A�I�ihM'`	��$���eoE�Zh
'K�;���G��j�X�m��v���ķ0�3[VԢŬ �W��J�Hk.cv�i�*���TT�r�(W�t�MK�����+ՙj�M��1--+n�H\x��I���w*-�͈�oB���v3��v��u�+,a�hu6��s]Z��jT�4��8R� A���Sz�-Va�u6�cUmi��!6��4NV�[Hk6�¯˼ɴ��&f��D�R�o.�5B)1����-���N��:0J�$��䣰k����^�-���6.�ʉ�"�p</.��$6rf���\�׺��BTԶ�%�G�GV�L��Y�1�#w3cq���%��������A�r�n�m�CO2��fn�9inE��)=���*�K��Ku�:2�*��PC��l�-��I��!4��Fn��i�P�HX�/��+1�!K0�L�����ӛ��Vh@և��q$خ�*�}u6�[;p։�ҳ. +	l��'�[E�R F�C�mM%�S5��0���>g,�Y1���5+�C�Ut�In*6���6��轍�>Cm�eF��[B��y)SW/0���՘L�/H!!�ԗ��5m��G]ܭ�Mt4:�%47wT�)��+�TWY@Dĵ5�Fjo-�̳NK��,�!@j������qI%9ј��� ��z�!ݶ�Ur�V=	��@nZ%dwz�c4|-]��vн֒��;%E�[i���^�tf�����*�'l�h�DAN����%�pm��ۂ5gTc1�v�ͣ���)�Y�)��d��E��[�0��}����`�Z�tuZj�٤�Uԡ�!8�kud�4�"xV=؉V�B�U �j��܃THݩ�/]&���L�&D�?<ܷ�f	�m�V��{&i �b���Kn�;�A�<��R���k��)fY��*���u�2�B���^��m-N�n��ɻ[%ِQ"9W��j�ܦ�8�"p��`��C ��)�N�Y��X���dl*5@���'.u5�,�U�]�n@�h$͆�HB;
/hV��u�˘[�x�D�)�$��O����&4v���3E*,���,:"V�6A��
�@�#��DV�*!� ��.]H+ZҦa�`��V^�M1[eݲ�޵t����ٲ��2�b�d��V���ڻ�[���͕����F�������Ɯֲ�z{XlfJaj�Zm�th�Qb�v���P�M�7T���oH1����v 8$�YS��Ʋ�#$J�;���K(Pt���kq 6�6X��/B�Keއw�gm��F+ l�oNڛ�Ɍ�{S9!��b�OWV%��2`T�����(e��t�V�QY��\z�!j��1��ڕ���:4@;����L����7@����²�5[1�j�e�U%�ڕ�)Rͤ�a'7%��0�7���˼q֑�yd�Zцn�z圍���X�Q��1��,9i`�@���i�f�k�iK�TSXۖ���3^�t�ٵ�v�7�F 5�j�;ToB�i$���ĝ�����r�l�DP_C���w�6�ÂJ9{�[�D�v�%`��ORš!���՝
P��t���其Ԋ���n<�6�|NU���5��d�h]*�tMV\���E@���e
;o] ��L-D���R����ύ'�j�v#�����p�Ӆ���Q�dKЮ��ۧKqD1�v�j��ն���٭��x�Gt a��a�̹�7/&U�cxӨ�%��#�*�j����!�e��%7��`eeR���@�W!�QV�`ˆ,F���9r�������Atf��F<�gfke��O#l��#n�f:�y1�z�m�2��U�t�c���#�eb�h�0]�C!��Gm3�IB]ĵ�j����彶��5rb�]+#���%^���;Z���r���ۑޯ���tw��U� ��a9kT�&$O�b!�����	
�u�[���k5mm�V-R��F�K�`�6/I���tQ�DaT�off���,�b}Bd�&Û[�݇�KIUԦ	":wh�3j�^��o.?��[KAq�V�n���ᨥ������nn4@%7��(O����I����2�Ԭiᩢ�� U��ѣC@����D��u�i�WxH�y{�^�ɋh��Sٮ^'DLgwIJc.�B�L�5
y4��[��t�CYI �\�VS��{�)5�y�K�3H��^Z�e5xƮ���x�փv����YrbBI+.�H.
��6	S~��gڋj-�+I�c�1�ԫ��)Spi�x��2��P�+��� l���1%<"Ce���_]l�oN��q�����\�&��S�t1�	��K.�<L�]�L^c��0�(�V@ f�R��u��8��iP,�(C�qՄ-��pVt�c*=X�I`(�ުV%���i��"�-�EI[4�c����)��F:�6��3F��Ȗiq	�I�B�N:�QP���!�8�2��;�WX�ym�vcT�th���l�״�V-��d/kt�÷M�iIWB��}t�Ymͺ��>f�ǒ��-�Ȗ�����U�%J��b.;�W�:� CK\x�P�4 P�0V*��l{+>�ڬ����3U���pޤ�s`�ԍ���9X.h��6�E����㷙+r�G�
��Y.G���r�C)ئ7l�e�!�pV����F�6˸+-nh�������� �/6�,-0�������LZ��2儌ЅH�+&nEz{I�d�MC�qT�)��̱oBWx�v�9O�4��bZ��/�5"�$��bҬ��Z��"@��1
˕��J��@3n]n�S
�J���e����i��� �Zڭ�(�DP��LR2�Uۻ�b@�O+PB8-btӈ�o\�u�3����6ൄA.�:A�Q�tH|��PM��t����Lܝ����ՉX��ج�<��K��!�M@n��B�VX��f|��j
٠�o��3	h�x��Yr�6F0F�@�-ʈ�x"�v�[݃olP�.X�sŻ��8z��APN��ɷ��J��Zi�Қ]�IGQ�d�$]�7*n)�wY�5���P{`�Z
){N�cH�e�&�����&M3�(�BŦ��+���b���T�AR���h��h�h���m�S]J�eV~uo뱫I���ֵ�-ST�!,�L�_BYʹV�6�Ff�D -�"��7
�
�����h��K2d�6`wrea��i���G)ɢ�<�M�n��]��ϰkZ�|1��׏���"�j)�Kt�I�qnXhM�::0��dbV�u{��[��l=U�`T�H�K�CRq,�vv�� #�6��q��8d��O���^��V]��K���h�:qb�Y�-�D;�ϭ;:赟<]���P<���g�(:� `�o1;�JB�⽫;��b����� L��AG�Ci�P�FL�D�%�(j�z�V��%s*T��LF��x��Xr )�oS�!�.RNԨ('G�����-��i�B��`n��kA���h�)-V��+-cG�6
ڛK�(��D8��VsX7�ӿ;�~�@���nϡ��5�ni�;���M�����(�{���D�����+v)2�5��3�7����YA-Ů��u�4]�	q�f��:r��V��`1U���	�$�ko�{�n+�4ͩ5�&���]c�6�r�%��5F�MFɿD$j��Y���	m���?�Cn���X@��%�3m^^�9�$1��2���k`�]��&��L����FP���ȹ�I`Q�W��Vۘ������t[c)����F��f_e�1�ŕ%�4�@F+�3A���r���S���Rj�ba���R!��F��r�0�lP�OQ�q	b`��U���D�[����%�X���4��ڝ=���*�J��l嚄2h4[���^ˣ�JH����v�vQ��al�Z���ւR����/F�)=�j�	�30X�SU�x�Џp(zu�,��]�X�jV�KnVJ[R�V*\"������yCU�]k�6Z#��t�˔rmIV�+Y2G�*�m�� KÈB͹WB�.U�4C��]
 mˑڵ[Z�����_Y$�r;̠2g��M�6VFe�/�e������U�2�*��a	hq��̠�oSm_7W�����\��!�)IgZn[�Z3rڣ�P�Xڥ7\n�l��i#knѸV��&��A�y�͢��m����1��gFDԼ��#�<@�Gw(ҨUn�
]�q�9g)VĄ�������a��M;��V�3�HªU��ܩY�9�����:��F��5gm�%�,+\f���=ڽu�W�LWl+e]m�ȧ�@m:��A���H�S��t�++5�,f���-�e�r�H�yG㥴kMfj9f*���,<�큧�+21J���iY�emi'ljuo���qf��l֍F����f,�y�[gs�z��m&�e���r=����x��K�V�����@%�i��i���r��v�������THV(ZѼrmI�";[x���b-a`	(kM����7B��W����]G����Ѹ��a��E�k�<;Lm��kUb
ʨն�l��p�]8Ș������
�˫+��-c�h+KN%�b�m�A�*���w�8���rw>�>�V8�ǛYHR���Iδ掬�r�!�
����ĳN4��K肖ˉ%�t١��������qQ�pV�>��6���+f�⯅�V�,�ꕳ�$"0w�&�쾲��ѫ���[�����WMpĶk~�
�N��2�9;+3i�t�Mn���uRv����LN�o��kn��t�Iʛ*��0U�ohZ�KiE,uc�'�1X(nl�����g=�@�Q�t�V���hUf�h=���3G�Xz�8��P�ޠ�L��v�=y��é�}���GN�q��"�=M�!}�U#���w"6�ó�Jd��P�����`�idQ!�Py`�l�v!Ή8E%;�s����g�Q%�2�V��hT��.����&#�	��Վ��{o3�v�]���Y�VčY ˦v�uLL�*�2�/p��qe��w�%�O��y��>7����%��� &#{�[��I���C��r*��P F�a�v��Y�wQM��8����i=t�tgq�iVgP���L��D���!�3���"�"��Ր�	V*q��o��r��=���F���=��J�ޞ՝�JY�ݮ&�ӻ|�R-�̒���C�U���
¦�q�V����n(�B�s����*U�ZӦ䙚V9��p�u�a,/��3�y�dn�kߘ1�֚��6��wKY�аK����Yzj�E$ȏG@��v#�g[ޫw���݉
�u�a�0p[���&M1K>�C"�=>��ַ��Y{5W��#�����մK�uɹt��)Jvi�����
@���&���5>P?h�����K7�P�R�b��t"���ʕD����s�����jܧD������Ji�|��xC����T�DD��� ��K�B7�h*��s&>�K���4�-6jZ�EJ}/m���V��b���59LK��E����1o=�V�Π \3�T��%�f��M!7EN�Z��7�V�"=!@tf�WM�\�D時�5p;h�+z����ǜy|eX���bndg�^Y��S��z���7y��X�|&�����ljͷ�6�(�؅4�N3h�wy%$wt�;�>+��1��6��x�X����Z^pC���s���q��ݾ�qV�����Gx��hSձ�`v9+Un��,�,aX�ۀqΈՠ
�5N�2�&4V77v>-��Fz��N��޽JWY��$M��<,aOU����ZUl3]Y\���9Z�����V�foege'Sw�5u�Cnl��ݻtf^�WZn���TY/r^��e)�"�X	6�Ho�GC}�.mtT9]A���B�;� i;y�փ���{Ҏ҉�;�e���rp	�����A�����Va�R�T����m1�w]��k��s�)�
�G����!��
���"z���	=\:q%]L�g����u�X؅:A�!37�h1��P[]jYa�����z]oc��+.�N������Nv:�!3�W+�N싔����3O�r���Zy�̶�b�u�e�Rm��bd�6��gV+�k�)��[�*һ������B�ö�㗳/d�����S�S�������$���P����^�w�Ͼ�f�%�K����-��nOf���9h<A�E`�\�8���gfuн�㳘l���/F�ԏ�I8gٛ�F[�:UX��w�ݔ(�aeI�O�]g�Z�j�=������6)��%|�M�A��J�{bK�I��B�������ں+�n����U� jыh�Q۽���A�d����w����CUf�=�e�v	#��OkVe�:�P��R�;]�e��V�#�b'��8`8&�n��[��ɂKĥ�֓�Re0>�
g�L��+V�HIu�;�tT�Y�"����g�W�;sa�Mv7��U�N�q�֝@�[�Uh��q9.����}[C�H+����Q�'cQW\;2�@Њ�De]m���yzF:�������-�a|��+;�h��}ηl�3,��ύ�7\�Ԯ%i������P�����9nGmK�w'��2&vDY;m���o�y:��	`�;���/;�����ׂ�FB�+�
}��S/�齺�Y;(+ug/~�7���v����]N�ouu�w9N�����㢗�7W���wY�cqJN�"l�G���΢,o��E��cig��C�Ԙq+�w�$�����řʮ���op���*�x�}�8iu�����5��:6.X��N<d�s��0�û��  �S���W�	���q���gk2+PW/�so�>2kKG*��r�N�_^hJo(�`�z�ZB�Y�k���)��P]�47S�U���B_ne�B�h��󒶘��w^"n˵����C�
C����;�e+����T*r6��f���(Tv���Z󻧖��[<kqiU��N�Ռ�[G����$�2��nR��{��N���r�����K�>*�u���mc�_��8�xO"�K]_�X���S>�n
Mu�(V�E��!���ݧ3w�u�s5���yջ��}Bt�h��R�]�1T2�Č��.P��kSJ�*$ەd�
�.��$��*��Z;wI-�ȩ�g�ʝYV�gt�hr�/�`�3����a�P�a�е�뵥�;4�\��5]vm>�M"�À���AyP=����^�K�����d�0D�]��2 Eff�ozC,���n��0�V�]׽t܏h�w�D�-wF~�Jk`ȍ�A�&��Ⱥ��T�t�t�=���g
{(ip�4�]|�q���U��v�Λf7E�ZUݼibkt�
*.k�s���գ\�f����s�<��R�N�����G:��V1|䐵�@4Sv�]<�;"3;�e�[Ym�R��*4�R���6��F@��e��1�8�f���;�lE��1�C�#h�Q(Z�z�@3�X坚lY�J���/�\a�ˏT[t셷��4E5	vW:��+��������ɥ��m���.��Z�K����J�ȱc��*^��#��bZ���ڼEZ;j[�����������eNQ��#c��|����}��$"�9+t�v����0����Nퟮ�I:vqz�����=g��]���<3
�lm`viΰ���7lL�=2�GrM�Gܝ�'�Qal��.��L�.�����[�Cɞy�h�㓨_$�z`�ZT��Ƣ$���n�E�%���o#�iP[P݊(uy��[y4�rvX��CWo��0���%+�hÀ�0�ݗYu���0d���L�13�NVһO7�9@�[��w0��6b��C�h|`��0��F�.8;틥v9w�����ow�ڎ�����Of�^Ǻ{� vX��p/�&��*��[�e�R��D��� �K,���\��b�ꥳE�;7���c�d1ݵ.-j^ۮ�
��33349���
W�rX�s��r5�r������w�����.��j�dK�	��r��у�d�R�\�9��1�^�+l�f�-�WNq	S���H��[(6����	Q�h,aO��Yؕp^�*�!XP>R,�/W,��!<�ot�OA0���h	|�3��v�wŇ�:'�o#�ɼl�n�f�cj�vW\+���kB�1�*�fNcx�Mìh Y*�Aʗ:��{��7@'�S�|��ۡ��P)�0u=b)J����q��+w�R�׎���N{�[Ė洭 3��",u�\�0����OAN��	��e,Ll56K7�V�;C�eo(�Q�^�B�F�e
�c�W,�7�����J�4�<8�\7�6(^wA�C�]�W�1)s�(�d�ϕq�~���9�b&����0�F����uwڒZe���wJ�i*u��dP�v�sN]pP�4��NYw�n^��Պ��ӎ�K��HQ�i0���ǯ�k���<���q]Մ�R�kvvR����?I�U�
�d x�E��ծ���<�RZލ��[������*o<D��������f�5Jۛ^��m�O�$󣙕�$�-D_rN���OU��u��	]I�x˻h}���V�ʴo�cë]ݑ9K�v�i���Q���N�n>��P;!�A��V���x]�ێf�o����7����(��hfF,�]1��,2[B���6��wׯ�=E ���XgQ����L�����:��:��*p�ՊŦ9�fo8���΁�2F��=\���͝zP�qJ�{G��fsu�OP�v�-F����b]z'v2w\�*V��V��Ǟw0.%�)[\�aзh%t;_i�[�`F)w�Oqa=�r
���^���NR:���'Q�%^�5دH�Yf�9-���/P��k��Q<�W6�����[+�wP�{ҢV�j`)����o�'ݑU�atf1��|���6�閟6
�u��KEA��Y`6�z4-�/���l<�H]Y;��}ǦhF�S�[ׄ�ZO0>���B�b	KH�Ϟo*R\��,o�{r�^��Z�ڶd�	ջl����%��P�����k$�^S��	(b/�=jo��db�s^����o%�ة��J�M�f������L��,R��C2�w%��O}դe2�O�c��2:l��W;�3���r�/�3�B�1�c�
=h��s7.������ѳ�ڰ���ֺ�
f�T�z7�ٙu���M��
h�SU���;{�z�3�ӫ�j������'��]s �C����͊��5q7����Pݰ�Kh��.:�J��s2��n���Z+%N*�Sq؀�J���"��˾Qmi�S���RЃt*���v����RFWwc�I�z��e�{3t5ET�{Or�$�Đ�\:A����U�! ��/N3������2�f��������Jh|�����ʇ[�EL���c���ֺJ�[ݎ8�_k��R@J�k���_-׵�N���<��h�N�cr�1�;�U��WJ:��'F�z��3�&����*�X�~ՙ�v��{�9܋\�c�x�>�V;N>�;$��͸yQ�2�HX��S��zLY�f8N\6�Y�Nt6*��W�ԯ�M�`M��}�:��^�eǾ��&d�({���[�.��[�ȵC���R��ƹ�G�Ι�y�q�h9f޴��lk��8)x*�S��:�{�۷N��;#<�5���ʳA"+3aci��$㽪h?/)��ݯR�`���B��k�K�����]�:�.묛���c�t�Ӵ��G$���LQ%��]��۵���i���fQ�J��/���Q�3l,��1^F���+�ɜm!��첢ۃ*I�{ّ�m:\��k-)�� �[���������x��@�uCl!�:ηY��vs�}r��Ҩ��ƥt�ݕhʸ�d�������D��+<В��`M��p������ەy4dި8��"��"T�u�m6��Y�/�ܔrѫ;[�;%Ւ>�κAmGKlD��̽4�Ye�H
t��g<<�J(�
z(���b� W4�iX�T��2���Ӣ��i���&��32�c��}#t�%**��4E�ܤ9O��I�:����h���V)Lf���w�Bi}�w	a���Ka��mN�Ǭ	��*	`5��,�� ������Ut����,^.����w`�|s�";�01K��w���c���wU�m�c�K�����PY��i�Mr�S���T޼�"�벺��;�3�[��h�:ȧ�[�Γ/�<�j��A��g��U�8tͷK���k�oZI�5�h�՗v�B�R�}�'� v̩g�E�bh�Y[��Z����E�t�X�&=��;.��
��;>yf��S6��b��/%��H��M1��u�h�L&�n���䂮{ؤ#�qon���[��X(c9Cf":�w�l����ubF%�vb;�a�����I3��fu)qZ&k"�=��bnvTmGm�<�r��"6���b�ַ�F@Pv�-�x1� vi����|Y��%�{MUܨ�g5u5��з�����e������%�������6`�RN�|�����}�\K/)<�Bdo���Pr ��.����f:��^������)�5�]4��b�`N�v��)9b������5�g$�H����N���2^�B΀[����)p�Ux"U�cf���qE���ۧQ�,ћ-�e�{u�c�LΠ�|Otm}2�� �Ŭk�5G��5�OJ�z�x�1L杽8�@��3+�vы[�'{ �T�8��F,�ȑ����Z�p������o�ձKڻ	&K^V��^����޸5g����*�������]5j�j�]�
l�@ϛFk��枬oX�S��	u����ݵֲDh���A1�8�;֦Ge{2M�h,"X����A��Bӭ2��[��9�Quc��n����̦rUϕ�mc�,uI��.ga��(�N���!����U���Fn�r�q�)h=�u�ٽ�=|x�W7�lL\���l��x�ۡk7q��p����ɌS=ݖ�Ӽۣf(����ېΜ�+�����K�i��.�ws�R��&5^Z]ݔA]X8>�2���k�V��z�ګw����G�'�p<�0��OYu�#�Bbaѧ����n��v�QYv&��%������Q��W�����aKz��u�E�G~���9�wX���]d0o:�=*�o��O�J-6��B�N,��暡���v]�]��K��t��0:��@�&*Ό
�ޜfƕ�6���wic�%&aS��J�īy�X��$=o4�}�EH]_-�ǜ�D��T�S��5.�\1G�Ƿ�(=��ɐ-	��s���!�l4C�B��4�5H��Ȣq�ѫ�U�N������y[�ʼk�<�����o{���3�?�B		���$������5��������T�AS��8�6�!OE��X�F�j���=��Pj;���P��?,�o�cy"�h(W]��S�:��%k!9R�;�W�w����K�r�Y(�Yb��)�,��̙S]̷mbw����M��6�nN��m���hK\Q��.X���j⡧ A��.>4f�
N;2�^�Z��$@D��e�dPˣ/;s�q�R�쫳ZC;9:U"�Ĕ5�c&�M���稂���̦%3�ϫ4t��LЬs1s$7Vr����(4NT��Ǉ��1���m���t`��Є��:貖ӳ�D��]lZ��if%W�����Z���<7c��â ;�z��H1}���a+��\KU�#M���3��!���"l�]ɝ{r��b�l�۵�d�U�Ԗ�;hңë>I!���Ŵ�6*�`�]*�9"��Q<-����@Cp���rIl�4�
���1������H\��/��i��[J,c̛OG]�)ˑKmlU�r�
wA�Xu��*U��ì()�b�j��uC1�j�{O�����K5�-Ϙ�+(T=��J�ړgw-o�d��\Pd�e�Ց�n�Υ���]���c�t�@��;����wN�a�>O�,ʻ'�ZI\,�ҮZ��Sɼ΅�C���W��;�bM��gA�q�ë##�`U���˦��n��ȶ�9��u;�����&A�6iP2��;m�a���-�SP�%����_qZ4�'yl#p�E�ʾ\5eʾY�	�a�#V�hWM��+q����;��]��qJ�	��ge�;fā��:�V�_QW�ʹ�Eᵩ�*Vo�j��2��_[��G�[*bANe�&�G}sX�͟�ڽ�s3/$���\v�bK���h
����V�C)���'e�޽ֲ_�4]����b�ZQ&��Q�SO�C�ﻄ/sS WɃ��[q�'_C�8:�K�*&U�7X�Yԓ�m[��� #kF��cV�ۈ����	�$Sj�Pg_e�v5/�l{N}ù�d��nQv���M�6�c[�3]K�LQ"���y��u���@e��K'#�6�NڙT���F�帳^��jcb�t��n��W|:Uq:��7�o���Yv*Gif�l#�����L��fWp��B�:ghB��$���\��P��6]��`�9�p�-N+�`�91|m��i��^�C��Z�"����+gE׭T]O#��g_օK7}�+!{]�U�=M)o�uF���ᰋ���m����O� �R�V�]��6n�j�\�6�ޥ�5S��-����"��m���:�����Ց���i�����mUy�_����Y�y�S�!Z��ڙ�Y�+i���u㩘i�1���n1x7�L��K�L髐�ogR�����Ȟ��(�����v��65�2���Iz頄Sm�Nt��뮹GN@Ƭڽ�B��67��wWr��X��1b�6j�
�E��u�:�Ŏ�\P�Z��WN4��#-SMם[%����
Z$/a�ƪt���Û����v��M�z�9�'�Ӝ�7�خ�Q��ڝ���-��X�YsV"Ӿo�=v+�7+$��6�t-wc�|3bmu�V�_���_vm�i/[����c�p�l�-(T�K���P���:L�g�S[w�K-]Lgn�_		��������V��)��@+ǏG�˴�]1Vj�>��;I����Dwav�Y����bm���pÕ
�w����ٔ�T}Zqom������A@���S�&�ѡ[er��|x�kG>�Tzd:e�X��G���嵪V�M���%X`�(#9����YY%N$wd�;x��Ί3{�(�li�qq�l]������rd�I �$f��}bˎ��SMha�k'�%��i����� �zxѷ�N�N��s`NZ���T�BWf���c�ݢ�ݚwS�X���r*e�좵���ӱㅩ/Rp��uԏr�l����͝W��Uhi�	����=�k�;���]
�6��ir�q`:,�	aEGt�l��f�|6�Y�^���f:F^���-�S �G6v�뾱ʴc:�h|�����E��W@j�I`��W֝9ZyEGj5b%]�S��ǭq�j��[��Ƥo�d�X�ٳ����}x�_6hgu#]�t�G��m�0-��5f �¶��mq��is!�w����7�sk�P�/!�k��q�Ѫ�����͝�9,O"V��M��mP�wE��h��+^\�:��c)l��-�`|;�(��y��rV�Ih�,�O6>ݶ)ĥq�s'w]]�K�z�R�I��*��+:�;��`��s{L��d:n���,���L�R��� �C�U,�V0�ǜ����ݷi>ʽ�i���@Zɘ�dٝ��s��xE:�K��b �:��:�%*��(o0-�4� u�����f��/n��'��n��\B9Gl� �e�x��@���]]÷	]5��R<�yێ������2�7׀��k�VZ��[m�T����v�1���Y���Ul��)n�����S?4��&�ӫ/�b���Ts�d���gɳg�=��N����\�-��J�*hwr�,5�U� 4�9��Z2jR5y���9��@R�e蝯�>`Z�LY�7/e��r�ᆠ6��Ў�.<H�����!Մ�"���E��V+�[���.4n������:���V����N�Σg��i�Ej��+���qR���k6�6�[��s;��uLH�^�`�DGq���f�{�T"�Y��lP�N$��j��t 뻧V/�}���'��a��r��V4���],HUv��*�[��Mg+Lֵ��򋮽�����\zfo��{Q������5�z���|�w$8���5}���Z��O0P��5y��v`-z� `V�p
�W(���%I�i4�c�*]nYk;���4��ۏh�s�zWuZ}>ֲ\Xu��U�j��bj@�$�J�U�� �	��ؖm��U����b�so��R�eF�����}(�k�v��d���.�89�z�kƝ\ ���!�N��&�֩������;\�n{'-�����+e#���Z2���h���˶�mm,;d���qZ;V�2�(��:�Z�w-N�ܤ���b�q��Z "�Z��ٕ̝B\�q�4�s����S/(b�1���N�M0C�\�u�0̤z�ww]��N<���je�{��T㕯�肭������YFX'�	��}�g�1�$`aQU�m�Թ���,��2�3Fh5�M �p�at��6t�ioQ�6�� �M^����M�{�����ϸ5�����_>��D�li,����:�j\	��"�p��m�"�W[��+n�;�ǩE��^_K-VvN��	̴��˲B*��Ygu�&��kCc�[�iN���4jr�0dʕ����{��ڢ��My
׎U�j=�Q󖫪eG���i�q�p	�u�*}g5��C��n� �wkZ�v�L�*��(`�b�lj�Z�w ����:3�����>�g�`����(0��)G�c�.U��G���q�-��y�F�u��O���&���nqNwHR�Э%�9ɨ5�:X��b���Fsq�9�ф)�c�*��G���Z�i:��D�Wl�ϵ��j�����oAҦ}
��}��i��4�*U�0I��T�9h�,����b��wг�Q��n[�
H�Qغ�3�I`��u�� q:8���j��\�\�B�wLR�$��:TQ"%cKXl%G3��V�ެ�j�'X�;
�ӚT���07yN������ؒ[v���������[�:6(H����K�2cZ鯶�A,j��!@4�}���j�u�MM\�䗃�W��<J�T/)MjϹ�'��d�l�������c�B�e�M)9I�T��,��{���5�]��韰�FÙ ���[�Y��sδN)�+�ȣ�ʺ�m����\�6�`��v.�r���9E'ָ��4tS�ⰱ}wU75���K�i�=V�l�ޒa��vWH�Ը��E���o.�3����.�K�}}[r�`<["�-�k��_;=]��]J:�|�]p��_�ګ�4	�u�8�Z�|CK���M��2�:�.��k�F*�Nu���5�rb^#@�u���лx0�0�ד����_u[xB� v���݅�7d�&��8:�T8�#��<i�T��e�%v.���w��۠���.�����rY9v�9DJ�r^�ΰ/��):	s�����3"\��z�q�GF\�ڄ�2[:��ྔ762n���6w�J��n���Y삘���J�r<����L|�H+�
&R�W�}ײ�Дj�K���{wk\�U7a�_:-�Z���k���Õc��ky�ۣ�+%jq�v��Ԉ9OWu�u)eD��m����U�/��ә��b�b�E���f"]�_"�[��4�b��vV쵍Ó��pE���'#Y��ξ�ib�ʖV�בn^�F�v�}��Ci-�d�|���ҭ,K3W`�9Bt2�=���������U�r�EӅ9�W��Y2�U|�oS�U�|�ՙ�����*3M˥��hL[ .�lg��Vm~Oow�q-V��b�tv�;4��t}l���y³Nv�hb��ގ�n�¹I�~&*Ֆ�>/�� إ#t��:�;h��\�-���:Gٻ���9�#��w�ݱ}#�Ck��m�A[r�d��w�����c5�ĩ�ʵ��{��-�������<4ha��aP+v��y�Gq}�!��ȽA�(̭B�f@��y����Z��)�aֽ�}�3��\�.f#.�;J���ke�h�:�\n����ݕ�/�D���1[V���t�E��ƒ"�UY�;t��[�,˭,�\�U3N�;i�aX|@�U��!��Nπ��颱K�a'x[Ϯ�p[wP7]���o��͓}��u;Y9ʝ�}Q�cXr���� �7��������8m$��0��Ys���Y���aY�
=�Q�e]_q1�
i�.��WM�ya}��s�J��v,�f��\+Ⴎ�u��7j�Zyhjf�i�F�Kz�Cnκ:�/Yu��� U���I��4s�l��-�c�#w��J�T�ˍ��l9ٝ1Α�wG; �"Wϵ(iG�c�v=��i�Ckh����ͼ���#���NY��A����W-�k�ý��Z��*���[Z;7x3��ݹ���d!���&�YKqV�q����B7M�*�^�s$����r���¶�L�o���̛h0f��78CD:���W��_J'p� }�������ب�)��i�̅`�v=l]��ϳ3��V�*����zα�C�.�1�Jعӎh'/,.�It��-S�8j��8����H(2^���M�������\��P�k,U�*1j��ɻ�f=QQn�2#"��[U�{$V��k-cj[��c�ܯ�릚N=K��J�,>VX�z��]ி�(�Q�eִ���Ճײ�^N�|�pw;��>��>�����P9�L�v���4r�hYס��b�^-(���[lQ�/�<t��*đD`�y2vj(�{N	Om���n^
eނ^5i�2���]�yZ��/ �Xb��Ĩ���D�nLe[Uz;�)�q�3.�nY�+"�N���g��OΑ7{@ɺ:�:q��eoc��-6̔��em���C��Ŝ���]�_S\.��O;+;9tV�>AE+!�'��wy��ǝʆΥ��}�v��M�xű��t�(Tn\���ʕ%]�WGR��Wo+6׎��c��^A��x��E�z2�x�)0��B�(W�v��{D�C��zoT�:�u�Q����V:��N����XFmĊ�N���)FJ���|H�=A�׋a�SFn��t�9�^�:��͢e9]C4qo�-T;����%١qR6#u� ��\y���ݣ�W��0���s�:մ�噒!Ϻ��|��Xr�2����
źƢc����]�[�k���&A�SY�8����zf� �;�#u�K�69�z��E��ubM̵���n�X�Dz ��\a��M�ݾ�®���;k��ь� ��UR��x-��ed��0lվ�T���;X��tNY�\6LT�:�9v���Am��RaCҴ+�ۣ��f��]�����&X!��p�N��S�wV9tĊ�Ta��XX��uf��L"��]�s[����V��u`M�=Oy&kke�߁j�}%�+�B��0Xӗ#�휊gt��F9��0;Ū�9|��D�X6ŧ�m���}��b���o���㫥"^�_u1�',��H%t�f)X���"7'l���gU���2WP>�\��!�S�Tס�LU�^t\ ��n�KF^��d� #r�p�`�(�?d�ञu���Y';�ev�4�r�7��(�Lx�寻^Nݒ�|��+�;�	Ό�vS��KDJ?�	�����דH�Ԓ��]I��l��Q���
X���XoN����t�Y,�������@��vs���i�h)�3O")hR@�ۊ0��8�eː�t�7h ބg8,;���f��/��tR��@K�+*�Rk�z�TǮ�Zn�V��G*�f�u�����LM�כE�y]7Z�fglp�2���p�=T)���Vtz0���ژ6�,�=E*���,�]I�`S�����71Z�B.��JI侾�4����Ve�_HzЖc�]t��%>MI�<�$(�3`�VMX|1�6u����ʭ�,��|9�`�U���˩muL�N���_�r����3Ky(���k�U��4V�p� ���)���\ߵ���|����@IJM�WbX�`Є_��"֍�N����ky�ZN�ؚ7�2f�|�..|�J���z	��M��#M�μ}h'Lvp�����,�%�2�v}|��z-�4h���<4N|�Y���1�G{,�V:\�(q�e%�wԍؠb�+�z�Yƌg�eu��ٝ�74:)I+k��"�j؎KV���^�K�;Q���2Aج_]�we�j`�]V��z���s�ū��j^,��;��<�e+��S��z�u�˱K�,@�9�V�B�����J���.j�O��rQ����ٵ��7��/hS�N����o�!L�:�Zż� ��r��LO��郖��v±���4µ[�Q�xk�^��n��q�G*s�Se���`(Z'aE����XK&,�tV�=�[{Y&��L�^�g����nx6���eE����_5+r����ڜw��1�{��iG��pV�̝�vA��3kC��UpT���7q�
��gl`=!��3���6:�å�`�T1.N��,�,,�T�p%�8�⩂����qܷ����x��ѩZ����k��V3\q-�2�1&�o��y�z#˧��uv�|mg�q-|=X��^P���h82]r�2
�/�u7���ii�e�"i���NѭQ��\������̰snȔ�Y�@�(P��)J[R+j�TkBڶ���[]&0Z��E����1E0�*��h5ih�m�ѣ[����*4���X֩Z�B�%���*Ҷ�B�RڪU�-F#R���mmiYF����J�R�j����E�)(�����FԶ�ѕ4El,��0ي�[klK`Ѵ��kU��0[FX�5Kij�)V��m�F��J���Fа�J-)EYQ-#mҶ)A#1��[e�U��Z����Q�R�VRҵm�#mj�X"*�����
�����ep�qj�R���5F�����E�)j�[j�-�X�k(���.+U
�ҥ�",m���Z�QkmԱ�YKE�b�X�(�Vؖ�-�TD��7(▨ִ�������*��UZ�)FUHղ�*�iJԪ�mj�Q�"���V���֊�-�*1lP�֪[eƠ����(PZ�b��h����l���%�����nI���k�������҇eu)�U�Lj�+hp;%�|�z�؏��*<�㙀p�J]�n�6�H��N����t��s��X�&A��\����`s��W�2aCAyҨTO*�D���4i�i1�eN⯽�l����j^��`&�R�tNgKU�q5�C{��f0s_��<k=Y;(��c27Pf[�%f��[zbY,oz̛ �[g0t���}˲���;��ٹ:�_���_f2kzE%0���R<<Te��$��ԧF,5�A���R�n�\>�� ���,Ν�1ZH�}�^(�3^~>w:ӥ�a��N�˞(g-�U�e(�ҤR��`���q�Ԗ	篠T_4�;Z.�/���X�z/(-{J���i���Jv8�������]+-.u{�-���ͥ϶�oe�]�2�e�Ӗ�8V�t�ʌ��-7�k�E{�>��g��I�Ɵb�y�~�=#S8�dO�+{;J��9�FV
*&��=�0V�e2�5������ӻ9b����VT-�LD]^�]��ws4"�a��L�Q���VN>�Z� �c;�׮����.�Ys(�C�FS�	}o�y�Z��e�
	K��3r렬�,��X�7����y\y�v뙭��)�_L�h�ı��
����a��"�$�7Ӧ��%ۺ�o˅a��Fg\��Lw`H�������ʙ1F7Kѕe4op���`�H���١Jv�b�u�Ǽc3t��,��4��O���<�z������v4�B�:2k13��ur����LK
��JU��m*s�����3z�B/{/Dƻq��C����h8���&�Ω/�R�V����t����Zϛ���f�_��1�BX����]ٷ\��IX���3	� �a���V�R�4�O�ΘRV,�u5���\�*��	X���R�-�PxeF�^ធ�g:g���ί^l �ߧ�Vt5�B�Y���Cl-u+z,�6�1�*�w���
���崭?tӃ�P���p�}��Q+o'�U�UXj^�����Н���B� �(	5�-l�wX�cc,s9
��fb��c��Z����^��kO0�Y��:�I�蝥�r{0�wf��a+r��,�2�0����us4n�qD�>4x7����n�ή#�;�jL��Ed�ě�{��7Rl�<.G�Vd�1t ӎ��,s$cPVD��Vs��:A:�n��������zo8i�|�����y���6{C�u5s����~�D�ֽ<r[��Pk-�.q�14����������\<�/_lm:u;<��3�a,Z����5��y��$�T�9+k*έǪ7=�J~�ٞO^��4��z�c�Q]똧yu��^�ْV��q��Xi�i�2�:���a��3�TAQ5��*����=�������h�1f�o��M��г�xUXDh�
Vzg_t0�a�j�1s�ϻ�����+��T+z��>W�p�5���8tl�*uA�E[�}Y�Z��s-��\}+�{�'��w�J�m�n�GF��RIT��-���C�T@�Fc��e��K�n��C-ٜ8��k:8�vx�����XF^Ї�c�zV��x*�}��Qv4{�{�S4OH3 t�i�r��j�.�b�Q5��<�^r�w������Z�EOU��:��C��S��}ι<J�y��79�^�{���]�iq]�=��0�J�Kj���=(�]]���[�)!}NV4�A0+N��'�k���n��67
�XwyM���_6S!�,��G1�"V�����<2��vX���FaĻ�e^����zۭ��7�Y�`"{P�Q+]J�-�t��=ۖw4Uv�H�ۍ���b"�y�(0�-��އT���9N�}�v��}��,k=X�(����I��������A�C*��'�bZ:�t����s�ʙ��C�3گr��נ��V����0�uc�jkn�<5㾝 ��z����SW�Jn3���J��N��	�XD�U�C�;z9^lC��9y(�E�1+��G)V�^�-Kڑd�B�˝�����x��X����\FsB�{��4�}�v_^�ֵ2�]�a��t�}�vt?y��k9�F�5�9v8v�m�Ea��;*��;^Wl�z�y]�҉�ģ�4:���yoyje�*#�K3�F�ޮ,�C���B��&�c���G��`����K�F�}J���2��_V���T����`�/"\�-������V�M��/n^��Č�3��|�u�n��Yj9�X]e���i�.��.o`����Hwb.w3��Y�s��sZ=����Z˝�-m�~�'mgT��G`H,
�|��>W�p�#�Y:2�9e6���7���ɪ����^��Σ�u�p��M�C����f��8'�ᘾy}m������>�G�{���#�/�eA��Z7ػG�>Tr��|aQ?r��㞪0�+7���8Ȋ�!�A9u<��_i����# �roݻ��@�,�U���Y��v�}[�3�v"����Ü!l~��1���n'��k�����n��Rs�����qM���	��9��Zn*V��W2��ˬ`q;}GԶ�Qc*7Pk��4�ӊ�m�Ma�p{�KSj��8��C�=u�K�,�7��Q�ܷJmg;�+}�/3�KW<ȥp��+)^����Һ��:�'-^e3��`k�ˉ$��,]#�7�R���A�kE�6��=bяl^U��I�w�ک{��C(��P�pf���啼��+W�u�S.z�d�����Vj-�p��FU�����c�~�[=��4����CX�p�r��{�fѹ�%.�V�O�h
�y�
�j��w)1d��TC.��E-e���wVq�|��f]�]�q�(½T�@�M��h��K��1�-��Z���ӿ{19&�.-��ri��#��<�[���s9~��1n��G=�f��`5J/5�y�.�=7(��⏨y^l��|Sp}Y��#w	5���P�7S緕ӷs{��cU�8��;�����DW�G���+S2�q�\v���}v�[d��Ի.����F�°�R>��b�V�:�AB��*��.�/<�L��9^�7Ր�]�u��6�tC#F�HYN���b~#v{x��:�gG�;O�Aкy6�O���dn�B>tP�`r���X����W���r%���v���/�^.Q�^�^6��:��C�V�J�Y�Oo��n�R1:��JYثYo�vݛ/��wt�ª�RFv���SG�C�C�z�a:<x�a���V��%/�#w��B�,���m����e� ���zZ��Ş��x��r��	ب7�X����X��0���&����-v{R��G(c��,�����gz��K�!�i���q��wBJ5�m3���P��S��5uA3 N����&�@�ԅ�Y������/�k3��5BK
�Tuw!��O��r+ҷ��ڏ[
��n�w�E���i�="�Wb�N
(���N����v]���s���X�H骷UWJkp��o{�� ��Z�SJBp�c)�.���T9C�G'�n��a��I��i���߷>�`g8	>��-!���� ���*�W_��׵Ô)���M~�x�r�c��1��TZhNֆ�<9M�G�ӥ��|e�oZDN�cOªSW��Pb�و\�14:-�݌���1�MY�sY��W�{NS���������1Y��3sJ���.�M�v��C�Ϸ��t�q9��J�EEkQ�Ew�'���{��o���xt�n5�����p��HV�g��Tng�@ƨ-�T�+o}��L�d6��s�@M��г�w�Ua�pʤ�[n���wq��Ӧ.��n����2R�����je\)֚���f>�e��:ϩ�z�
6O�i<���jͺ�2��A�&۴���f�gV�j�]u'[�"�z�W5u�V2���*/ F�][�E�e�po�h���l��Xb&���D�*��J�
� �ܘmuu>9H�o%��uc�Q�R��X���^8y��q��lq��[wb��ɣ��Ho��N�p\:�x�$si������Y�����g5}Aj�	�;Y��Tz��K���Z�m�*T�d�ݧ�*/���;�x�+�D=�2"��[�&9�=��`�)�5�y��/a�`M�9	�}����w�NV�aܘEt<i=�)���f_?Ӈ�$v?7'nY��ϕv[V架�c���,�>��h�Z�+rl���q�r��|�o+5š��3�>o#�"�,8�'��.� ^=z`�߽Th��9�H��36�݇Wm�߳�ܟ6T�h-N`��|vuc������L����r��У�>���j��נ�(��wIy���s�i楙���Cj1^���d@N�⊣���ٔ��n>�,q�:ވ�a(K�ӑ�k�p/���w� uقpCvk�A�j�U��}L]Zdr�#�J�"f\?#٢���d��o�-"���YȵK�.�r�Y#3o������4�bj����]쥋8��\�q�W]J�S׊,O
��u��5�Fj��2�2�N���J�q�X6�h��O�_Q�e��xB�iq�Q�LvW6s0u�rɮ�J�R����q��0���{oe��'ҰD�-�x�:.��T��Z���pb�1Y��y��m��kYy����6�ɹ�eR�д�������n8��zD֧݁ V���	�{�9;}�7R���u�#�U�|�T1�a`�y3�\v�v�XO�x'�J�H�B0�8wsS������;Q��.{=+�UE����\F|�W��46[}�fg���\.8�i�DqtP�fc���J�r�f;�s����9���g�v���j��ЎCc�o�y�`ٻ��oZ[c��^��Y�q�|��!�<n�[�f#���8B�{YP��(Ҧ�zvo�s�]i��s{�:��K�%h�M�,>�)�b�-[��n�h�xll�6����Z��׊��ƒ�I).�T]C{Y�D�/�FoFs�K:�m���qA#�I�=rp@Wk%�\M8}P٢f�p��{ga�PlW�N�)1��%s/y5�����p�Vqnm�s7�.WPN���9��駱�
k�cz�%��q�4T�Tim^�,en���}�S���Z��S`�����I������v4���Xz�V���1p����}�5�ONn_�k|]�ݎ�� �&�g1�.Ջ}rW^]'Q�̦5�
�9mc[��Z&�w=\L4�z1a�zZ�l���l^P�y4�Z�][��R���<o52p���?v�;�E��N֋�r{^�f�g���ǐ��zp�k͵}8�8��W�N'
\��&��v�s���1�dC{gtwK�Hp痣��Gi�J�PS=*2�1Y���7p�[~ƚ���5|�g1�"��%�u6�Li�9~��b^
*&��=�0V���׶7z����wt�n�s�|���_4�d;}���\&�')�)Ejc#�$���$�-=�f�����Bj��^�6وtC>7��3:���?C���n��=$�֚}b�yt��o��z�v-X�W5�dW�յ��'u���-Z��`|��|���>v�A\6��)�F�?X��1o]*<U�Z+evt�5�p�#��h�0r8�l�᧡�Ǖil�D@���WT�X���<���v $�r�C�����3khQã 쮼<��9ֶM;q�K����]�N*��/c�]�ÂN�W0�8�}�7�����+�ؖ����q5�P�P<�������m��^KiG�"ϊM�/*��蹑۲��%;T
��RZ���kJ���j�.�U�	�̹�)���C�cL�r^�e��d�N�'�gR��R��F-�t�WYm�@+��G�"��a�(_u��__ڝ�7gV$����z�]sZ+�t�b�J�IHe,�p*��rOHA.��\q�)�P���Q��~׊*����o�;*����r^�����DN=�嗶r�b��'�bʜXk�b�co��Zrk��b��B��u��B��9�����;(���ǑL�YkY���ā�d�1n뮱�6T,�Y��gާ��<��c]f��7+8�S-���GB���� tm=�[WZՅ��T9��`&iUz7�U<��t7RP��̀�� �it��R�8Fp]s�� XC��B��2�M&��7�>۬J��y�h�n����ǲ�$���[�p�|��.<-o1B����	��Kz��۾-�ǼhT��ݮ�ӥ́M^=J�f�Q��R�l�]��ϫWLB��z�E�Ԇ�����^Tz��&f�-Z�͡��'}�4	���|�)j��[��:���w7C+�b\p����K.�9�j�ݫ�X�C�G8�n�4���*�D���Gt�K_dV����p�������:�k�k#V�	���bg4��њ�!lֺ�����G:Y}�oK-�3��#]�؍�k5-���{�oBWh���"��{`L����s AЬ���@�/x;�g֓��X�S]�)��0���N�Y �]6з��W�Nf�P�������q��\;j��Eb��W�vJ��k���F�4��z��QJ�M�*t�r�.}7a����Oq9��]bG�k-P���.�ev��֒4K�W�k��/�:� s1�ճr�qk�����K��W K�����J2��y4Ty�2཰��O0�z��9�	��6o�}W0��:����'��U�&[Щ�B�*��UŮ�Σ�$s�������m,᥿������ʫ�y��t�U+�	�T��$�^��{9�B�J�f�W�m�V��(ভ��\\ ӝ��������]�n
��M�[ì�������C��9�����P̅In��Zq���!a�W[Z#s
�W�G+��y+�z�T�������-��B���ݣ�F�9U�.��zy�t�`��r!�j����SK��Zp�:^u坘V�7R�P��&; |�������-hV�[*UF�Z!�*1c���ЩYU��%j��[DQm���F*�T�,�kh�J%k-��
�h�R�E��V�P`��j*�i[j��+Z�B�qj#V�m���1�4F�"ZR��ږՂ��V��Z�0%q�0b��T���cF�ڔbȉ[bV��j��RՖ�5)KX�ZX�-�P��mTQ���1���-R�m�[JT��Z����eJ�.-0-����A�Q�-�T�����j�EPEUKVʑ��T[j[mZ6�!mR�Ke���h�VѴ����*V�,�kR��X��V�6��UbQ�-����Q\[ ��0U�����mV�jȍT�-ZUU��E+,Dm�$��+m��`������-P�-U�UF�X�
ƭiib��$�X��c��Z(��U*�j�5���Klce�(T�[U$�EQ���UXV�*��U0��QQ�X�*�"�ZYV�ږє�[eT+
Zڈ�ʣTEX�J���� EF��T�Z�����������Oq���������<�<r�ܖ�`l�:�s��]96fA��S3��c�t�:�����hU���-psc�j��:(v��p647�pQ+0*/����N�?JVb:Ry��w�Z�����>�c�c"�ֶ��������tz��s�,�8����7�=F�r�J�k��MW.9X���
��}0���f��v9�=�'��E7m�>� �6�����-�.����t���'��|}@n�K��
US�w�n��x��n6+E��f�^�6̭tiuY�n����V�����\���|{�5niAN�T�s�e�����47���Sa]�n��*��"}����&�S���C)�4zŮp �ƴ]ը��;�EX$�sX�뗱��o8i�S�����v�f�+�4����8��U���-����rZ�f҉��8�M��~�y�۶�>��2�-�"�r�l��W�|���ْ���k�5�2���9������ܑ=z��w��/8I`e�{a���V����R|�U�A��y��� ��e�i$�y��Vq}����R���,�[O��FӚ���q��WcR�S���9���frm������xL�������Vr�C��g�{0x$ej)ñ�N�ޜ��S}�|��m�hE{(��1�9�N>wzq���HO^8����e���㷻p���[@����W6Y%��|��J���psba>|yoBθM�Vջk����E)�=�S���'�T�+�`j���w>W��^���[���y�j2�_7��2���e���:��v$�N���"��EE�3;Zz��o1�:���8Ȋ�:* v���u�j�;�]'��v�O��{�Wy̦�ͥO�;7{KD=�dEr+ҷ��;�[/���p��>O��k�y,/����!�<l�LK0�7b9����R��YuV�b�Ӹ�8���#����j��=���oO��g�*5u�Q���kz�:�|{�ڻ�>��b�����|_�]>ǚ(9�z�;'v#Ӑ�Ѯ� �]R�2L�R�T��ps5���7|U�W;�7���
�&���ܜpN�!}���Vs��ɓ�.���ٲ�������[�kr�W*���s}	[V�18��I6p�!������jX����ܣM׬��3�ܘl�N	�ؚ@mخ3v���Ym9ѯ��4͞ڕU�����G�����N��o��;��f�j+�r^�0������r����k��+�Ʊ�z��T��8{��cӂOi���1���t^�핂�(7
.�n
l�.tr�v&�5���hi���퉲ǋ�DnQ��RsԱ�>�H���=]Gk���0}Y��y�\����睽�F�v�7����}�[M$2��r٫a}[ ��-�z�s�|���z�z���Ί,�Y;����ٰ���g)��gޥE1]� �$��J��:8ȵh_Y�f��t+��x�����z�`�8��u���$�L�a���qɋ��+�k�O2y��=����#*��t�N�^�JZ���Ū��s��I݆��7�>U���Ц{UYG��wk<}P���jo39��uր�C��u��}�Ӭ��Lv�V���F�¢@]����=y�w�KThT��qV	(�����霣���%]�G7*wo%��z$DC�8!�|���py'����,'S���pJ�m��s����y
����d�Q�q�Y���|�8�s�q�wϳw������㟿o�ǡ�'ݲ�0d�']!�X`y��=a>d��=d���{�L�d�|J�y{�IPP��:�d��6���=���~riϵ���6��sz�0zI���8�I��6d���y��:�Ow�C����Ri'=�'��M��pϱ	�e&O{���O!�^���	��|��y\�.��ջ*���w�#�#�="=""�����̛g١�O'�6I]2�'P<�ok�`�ɶ��n'�2�h���<�d�?}��I��y��]����{c���s����Y&P�3�*T��/�T�ed��d�'�Ϭ'P6��i�'}�I]2ݝa*y����y$�����'Xm�Ï����c��~�w�����(|��{��N��L���$�׿���I>7z��s��Ru�l�~v}Bu����C.�N���A|���c���a�cXޱ�߲��s��b�k\�ө?0�Oo�2��NwP�&�Y��'�M{߾2�<��bJ�d��1"���ؤ�'~t�Bu�����2��9����[�sn7�gN/7�^�1�?2mr�VT=���$���̝A`w�2��4ʇOw*M�{y��	�'㟱%2N��$R~tȃ�B��`����q�G���V�О��u��ֹ��̝d<r�gY2É?�4�2y�7�M!�3�`�$�����'R�;�2��4ʇ�`~d�'g�#�""6�="ǣ�FN埙�����+?g����E'�LKa��q����)�a��<��&��'P^k�����'�,�L�k�<�ԨL����'���1������C�Uk:��}W�+�u�5Cگ���앎�e -�)��x���-zB�6� ���cP�c�D��N5�fh)�$2�G@B�po3h��C�MN��Ը�ĺ�qv��f�rQܖ�|�]i�Ԩe1ݻǕ�}Z�<�9\�܋�_T �29�`�s��s��/1`zs�	�'S�	���&�,�$�V|f��u	�o���,��4��<���	��C��'S/����>�=���Տ%��G��Z�9��2���[��l̚I��=��6���pM�I��eBi0���ŝd�eO�C�,���<��L��	Ru�|="LG��|=8��_/���9�y��|u6�m��}���t�{��'�i�'O~Ğ@�M��s��+&��2�|�HdŐ�|��Ɋa�m&�=��ǽ����D��r�,t.����~%I��eO�$+'s��ē���0��XI��'{d�	�����'�-��m���Ł�>d�g=�p�b;�MbB�pU;�����x��?��}�k|��CI�I�ء�N�`sT�'Y=����HVN����v�|�>�'�q�	�I�L����Y&�>�~���C2��+'Xh�7y���Ӽc���߿~﹟@�d�{�	�L�a���q�(u���C3��u�����$+'�|{�6�$��=�$�ĚI�׽�N�c޿w�}=�!啺�P��ﾹ���"��>�9��Ĩ(OMY�+'PX|Z�m'��$�O'ٰ�|�u�1Cl�2����I��h��!�0Ͻ�=d�&Y=�O3̙a��{��w�����Oٔj�x��{�#G��� {�">�XbT'��B�q+'ؠu&�q��,'Y<���RN�,6�O�CF�$��5;�m��3���n=�v�7���yx�'�@��`�fY8�/��<�Y/��,��k����+	��y�d�VO���'>�O�'Y6�~��XN��3aĕ�!�w;��c�}�w��ݽ��s��y�A��1�ژ#�ǽ��9����6����>d�3�bC�m�8�~��L���*T��w�+&��1d�&�=�3>��d�9�^��m��������vI���VMiNּ]�z��0r�,r��x��p����U�e0	Cu")v^qp[9��$�N Y���^sY�1��,��8�����a!譡�)�n�ЮښtV&���;(�y
�i\7N�b˹�T7�q�ͺ< '8�W��Ew	���G������>��I�ֱ�IR��)�d�����'PR��m���B��O�{��)'�~/}%J�y�)N?�?w_��R�g3�O�z�R���p�X�"=� �=�2��'��5`i�d���<�*V�:��+����N��2w؂�Y6��}��4��{��,'̗|���kf��Y�<3U�ټ���H�����)6�@�6��L�M}By����y�):��偦|��39�y���C|��IS�i�N�d6w��:ɴ�?�����W���[����}��6��}���0ə�ؒ��N&ydR~t��Zd�|�5a�a>�I�'�u'�VM��'Ps��$���g���Hs�ڌK��P�����V�ϣ��b${��/��<ɷi9�L�d����d�2d��NO'�t��ku�i*|f��:�}�i�$�
O�M!�N�߷�⾏��j����T������b#�W�q�I?!�|��N�d?z�d�&�$�l̚I����ě@��m�&Y<���!�m�)�Y�I���AI/SK��W��zG�|�B#Dy�"!�{GY8��>�q'P��0u�a:��<���	��c�I�i=�'�I������L��R�|�Lɋ!��2y}�S��3ע��]a߻����=b"G�t:��`���u+3��+2u+;��<�1�Or�<�����O:a=���O��s�Ğd�rw��IXu���o�.����1�s:���i&Y�C�|����0�u3y���u��XsX%a�N�C����p��On�<���$�ԓ��b�i�O����~�y���i��"���X��=�1߳���Y2���8��:�+	ĝMO�y�$�s��q+��u���v��d+'�w߱��'�y���3~fj+�v�]1�A�����/������C�ٺqvIK�{˳��K�J!�6��N���A����r�t*B��e `�/��G���{�n 3 ��b�w���Wռ+ŵ�N��E�L���!�i��F�G�*�yoJ��=9��{j�7�I������a:�2&���VI�׾ĕ	��B��
E��6����d�I��f��	�d1C̜$3TC�yޝ��g, �}w��޵����0:���6�$�&{�I��'�C>�&ٖL���XO!�{?IPP�rΡY8���P:�l�L�D#�>��)�{�x����h[{bNUdk������,�x���18��M=C��4�w�O�2�H=�u2�ęg�	�2ə�g�RN��{��T'ӗ�+'�T��'��s�5���^}�������O���I�|f��WL���'I��w�O2N��̞a��{�2��,����m����y#߲����fW�߈�c���^���u+&��zb�l��8��a:ɴ��t�q��y%vɖְu����q?0�$���̝AHd�����LG�=�]V
aY_\_.�u||�:��߾%ea7���d���Ryi4����q����ΒN������d��X�IYP�,�0�M��2��@�߳�O�W�y��Y��G̝J���HVd�s��IԚ��IY'��H�q���bì$��?}d:�c�>d����I�'�g{ǘM�"#�?Ni��hf�6�t������=��o�8���g;��'Y6�����
�l����0ə�ؒ��N��"���l:��OΓ|��&��I�'�1{|3��_ەA��FEu��r��#�G��甓�a���	�d�q<����O������J�����6ɟs��d�2d��NN�yH���)�}����|Uw��R��J��h�p�{�t�|��L��C�<��T�(y���L�M3]��:��w��u�̜v�G` m'��q��{��m�I��fϸÕ��wEƓ���cR�u�kH�(�4J����!��V�N��E��a�a�ѝ�l�Ch]Iw��)E���.4J�̵݁s�{�}���w�� =R�U��l!�Z��2wBv�X��Rk����s�i
�5<�K:s�eU���S}L�Z|���B�M%C�'�T�L�m�O���'�Y3���:�䩓�b�:�8��Y'�~��'�;�	����O2u�M��<�#�{��|S��l}7�Z�U���Wޏk�t�k'�4�LY��'�q��2è)'���d�
y�B��'R�{�Bu��d1�x�<���{�G���t²��,���뿷��O���bO��9�'XI��?����'R�ÉY8�HdŐ�>I�g�h	�Aa8�͇Ry����b'Y:�3kމ��u}���9��{s��I?i�k�����I�/�q'_0��P<��N����'Y��~�J���aĬ�Aa��8��u�1p�6�S?Xy������!���������T}�.��9�9��z�i�L�x�v�T����v�|����8���aa:�dɯ~��$�5߱%a�Ce����Aa���"8{�����1��{prqH�d�7{�s����$��Xm�߬�C��q���t��`m��=��x�|�ߨ�2e�S���O�=������׳��	�DH�������e��~y}r~�en�����q�)FI�g���Y'S�6d���g1��'Ri�C�b�C3��ǩ4����I��'e>����t}��=�|"7Wˬ|�	�ny�⸵��3�zJ�����J�l�*�m�����g��5�u2�i+�C[�'P<�oh��?2m���ۉ�L���{y2��v�>+���o�'�ױ��s�s���~Iu�d�C��朗RN=IRq��X��&�8����_�i�'}�I]2M��%O0�5Q�=��y	�����u��e|�_N��s��'�@�=�(|ɴs�'��&���e�y�����T�&ޤ��́��N�m���C��'�>t�u�R�{�"'p�}����8��N�ʋ
ch��S���f�I����ÐC�l�l��J���t{��i�t_^,����ѣuj]�z�p����2>y�`����m�u)������c��ѦJ�cv�����9ؤ�Qe�;\N�J�2VG��e��6��"��ٿ��UU}�k�]�u��X�x�*V�k�6��&3���N��3;�AC��Ag�HT��=����y�N�ĕ��=�bE���
���I�I��N�<���nY��~��n�ε�}�ä�$�O�4�2q�x�$��}5�Ad�;�y��,���N��*�!Ri�s����L�~ĕ��;��H��遮w�����1��������k���q�2���Y6�|f�g2é?j��|��3��&���<��*l��d�T'}fRu&�P�l���h����Z����
ǧ+��{��ĮM��dR~v���a6�fwC)<��i�d�$�Փh|��'��'�:�{�O&Y&���py��P���b~I�M�^ީu���x�΍_����s��,�d�3�0�`zo�	�'3����)�Y�I����$��7�|��L���C̞As>�q'X��^b,{���>���C�x~ɛ=��ύ�e�	��u�̝�&�~�2m&��=��6��o8&�$�M3�I�'�3u�i�2�PY'���d�'5IRu'�S=��cʴ�������ַ�~|�N�����L<^`�']0���d�M�d��ؓ�I��w?���i���8���!�CI�'S8�&��d��PY&3��������u�ٷ�sZ�q��M�`x9���O2�{�HVO0��py�I��q<���OƼbRi�'��bO0�L���%I�e��VM����0��q��{����g�q��u��߯��N����É�$ۓ:�Ԭ����'uC�wx���a�`��=�O$��~,�.�6k߾�d�L���J��N�8��K����7q���s�����Aa��CL�L��M��f}a���q�(y���C'1��'Y=�s��=���I�&���=������y���3�a��E��5"�Q�x'怓�;��"�Xr�;�S����n�M�˯�w�hw�V��6R��N�7
���[��[�k��D�}Y�7U$:S��0�p���MqT�� ��sz�aJ�nP���B���s5�do/!�Ċ<I�vR'�r�߻��ܮ��Q��z#���U�&�W�D�{͟�=��PP���VN ��-�6�̢IĝM��|�u����O?�����I��w��<Þ�8����X�����;գg�2>�Y��ۏ1�q�_{�N&Y;��I�7�~��	��:�d�VJ�ԛI�k��'���q�'Y�I��!��XI��E�)߇XF�۩�R��Ϸ_,��Є'<r��&Ri�9�u�d�����d�ǳ�,��f{߾��a8�aY8��X�u&�9�3>��d�|~��_G��lci��®�q�࿎D�c�\�ޏ�WL��Sl���>a�I��>d�M�w�
d�6{ؐ�dɏg�XO${�$�RM�aY4�x�u��{����d웿�~6w��>�z�����v�u���J�&Xdֱ�IR��s�:�̓��\O�u!��P�&�Y���
�I=��|�y&���IR��|'�������D���Ϝx{���ӌ��~x���O u�f̺d���?MXg�2��|�*V�N��J�y'R��m+��T�I���4�0&�o�OW�#��=���X�OϷdRi���0<����	�C��y�):��,3�O!����&Ь37�Ad�>��d�VC�]�z>Z3��7��>�_^}�у�b$z>n��)6����y�a�3��%0�N2)2遫C��/�!���	�i>d�N��jɴ>d�O��'�<���{K�_�v�/�u�����.���{�{�cE:ږ��
������,X��G�U�:M�[�	珖M(��~��ߒhi��qM��,C=ed�����aޅr�^�l��v}o=�|v;ɉ��Tpռ�݀*����.���D퉽҆0��h�A���h]�����Ǐr�r�I#��n���ҽB��9��X�}H��/����ov�##���J���6�+) �R�*�G@vR�w8jS�����5�q7��t��Z8Wum�_��o��w���"k��.�h�P-b�:��f���JεS�o�h��9u��V�5���S���y��tN|��Y�i��C;HI��;�yNqCa�&Q���NprM{Bc˽��z������#��Vu\�Yb��jf�u���Y��W�;;��MGs�<�'"�5#��]��8b���\Ƴ��?-�𵐕��YU�����ӽWpv�1��:u��
✩��,�tP��Ů��OU݇�`u�2� ͧ��-=d�7���@�l��NXne���]Yd�Z �P�Ql4��� t��F�~90�q]-�ښ���j�;�Â�*��rt�B�m5�
}y,W�tf��y��67d�����zL��tz�-��U�.�2ADő���AQH3<��1���תU�OK��	9���i��-�XG�.�=�M#�)GK�o]���n��̲��x�t鲍v��h�v�O"�� �C�8&�afN��(�0a��)wa�Vbŷ��.���\�.��v���b��y����H�aݡ(�9֨�y� 6j:w�`�=�8^�bضSoi��]�fj&�[l\�Q$k��	q�P��-յ��*]��D�5@u��>�x���X�2�)�0�so���זq-r�,X�}���ƕ;��Ь5�o_�m�ޖ~�j�.�����X;#wu��B���\c8h�e��6�.�L	mc;w�dQ:���SZ���m=�J�o]�-j�P�踩Y�oeMVx;U�x�ou���S�ctwg�'j^G�{�u��f]�b��h������nM��I{HSyMjgh%y66r�!��q�n�s�]u�
ol`푪�tU��t�޶W(����**ӏkOYʛ+�	�Y#�t���oN�v�U3x�36Hu�yV��M;+����92��/�E�ÀD���,Q]Dt��+E��Sx;�㯯�0�Z�\�.�PV�C���qJﲙc]_^о��vE�k��D����H}��k��|��[e p �5n��ל��\�(�Ԫ�	a�cyӝ��W�&^�l������j����i��j]�m���ѵs��J��KQͥV��ڷWZ�Z��q�a�7�Փ�/l�J3�t�>T/0J��s��*e�M��:�g5�w1�˖5�0q�6� �0�K��������+%�w'S@e馱i"�AawWwm%7Ku�ymɎ�a|i�[a�u]#�A���=��j�ְ�+l�M=���X�NfH� �o)�����wՑ�(���7(�:8,a��IJw���xx;:�4��H���~F����9q���*�E*�AĢV����LZ���DU��RڌFբ ��-)R�T�,V��)j�*��DZؠ�U�E�UJ6��Z���e�6�ҢUeb1���"	Z�V�P��p��"��F,F�RUle��QQeE��jV��-��KV��*�	Ub(���KeeD`���2*�Ԩ�"���-m�A��4R�����k-�-�DER��--j�QPm*S�Pb��[E�J���-emR��-��ËL-�QETB�Z2�YU[cKk+QDm�-����UUjV+m�#[d���AV�,b��(�1cR�--)m(�*�Q��
��ETEE���TDUEBإ�Ub��Ԣ�j֪,QX�
�
����m
�U�Xұ(��V�"+[m��JʊE�"(�����f-ECj��b6�")R�b�DDTIDmm�"��Um�
�#"#��YiUX�E�T�Q[J*��QE�E�"E3]!%V�qT�cX�N���	Z��[�7�ƪ��v�s3�S��@S�1;�[k;���io,��������#ވ�xy%�ֲ��~���9��E_�5�����q�HVIY�َL�e�r睘�G�kS#�$
��J|�7|�,�ݘx��}���.&���
�{'�j��TB���=-��������h�evUxqf���`F!������4댮�=���_1�f�s]�3��u#iS���y8H��1��tT�}1ʼz������{☌"�J�:/���ٸ��|��Ta�����V�DTr�ώ�Ż"�o�Z'M�9μmf{��[�S�	k��v�^r�)aؓ�:+z���˂���7�5k���<��l��Ͼo����ǑT�K�&��X�ǣ�o�P�h:��8_w.˿RW/(s���P��:I�7���z�pV��թ����ƘՎ'I�������F��Y�}l���/}�vC��m�}W�A1��(�[G�� ,پ�×q/h�ڰ��&f��8�^��,�/�� =�B�5���b�VNoWZ��J��3�J��oFd�]��Wv�rɲ�Ʊ��Mk�{�	-j�W�9}r�� ��<�9���x���S��<�Y�}'��Vm��k���M�h��4�D��9«3�Ŭ�n��Lyj\N̿y�<����`_5��hhf�;�=bю�ʀ��Y��"z	*���w�pz���Z�Qd�ۈ�8É�bݭ�i���c/%��˹dQf���96����6ej�[G�Yh�g/@�O����l	�#u�:кX�RW��ۜL�:=J/��*8���=Miܡ@L��o�����;�vf����6����k[��/\���	[FOiΕ%��Z�^�o�ޒ�z���j��p�+"gY�E1]�!�5��u�d��k���G�.�5�k�'���u�ĭՆ|8tT�fuu�]b��sv�	,�4�w1V���B����h��\F�\q�ӈ�!�����$b��sr����1�㺴�Vc�'���yʋ8��7��ϱ��r���)�W��4�Y�k$����01[��Hڝv�+��g�Oy>����;:V��Ba��+����%���Fwn�a� �Y
�!�Q%�y�պl�ܮsg�rU�������`_���ǁZ;3)=A��9ŉ�G��;��Ӌ�n�q�z#�
�,\����3��^�K;!V��,�v�}KW=�o���e{:7]b��S��|��r ������n:�6㥝~�\��NjCvB���\���7o�Z�ns®mIK�{�z��qJ�E�����-�i�M=���oL�\"���+]R곊��!X��7�os��z�
Ԝ�ʂ�-���7e�ގ��ׂ;��N)P��K�Aݵ��,p����f7X��T$��hhf��G�Z��褢ͳ�gEf��]��w{~���.��Jn3��W��@�v�[Y��y��'�&Ԫ�q�-�Qy^���,����҉²3��x^\*�#��Ӧ����]�����w^K1v�����Ԡ��pb��c�w�����j�(:�s[���r��5��y�|�N�����J�ED�?u�}P�������]bu�n�	i��OJx���{��>B�^�bXx���9~x^&��ED��]�fdHZ�n�ؠa��U���<� �[{Sض�P��C�\+4�5���bc�ο�QwP�k!�`���[ے'bG����L�=Y%QG����{ތë@���}���7�˸�[i��v�n��к�m|v��X@a�!����W��70|�:�i�	��p��!�ˢ70d�L7�/�,rZt�n����3�Ү�{�5�B�oh��^��1���,n���r��}���8��><'��13��up|r:Ry�|y��E�e�ZFAEd��0$�J�[8�XG�td��c�D�g]�t����]��\:@��5�����ͥ�N"_��$I�zY�Oz�r��u�＞n��5J4�̌��}�2�S�uj0������[�jXv$�k��A=�)�s/Ve��v�K�K��n���~����Վ�Q}�S�pV�M�,@��w2]��YÖ�l�V��=��q\��q�cI��so�Tŀ�z$9%�,U�>��&��un���@��R���M���1����P1&��p���4�|x��<�xf(|��2�9o�tW�����+�I�0�ï'*=�=���7����״`��$��e�uj���/jh���ee]c�$v�|��ť�
��N����!\��[; �x��1q�M,aS��W)�]h�HVq�ñ��~�����2�U>������af�]KW����q�O����p/�-���Nm����J�l8�oE��ڌw�zţ�yA}�����ǔo!Ew�G�qnz�~�����^oy�ձ���VJ�E����/	�ⲭ��ۇA��g��I�}m>�W���i����mW��T�N=���{�6_��O��(b����^��v�y~��e���^gB7�7&��7F���\���&��t��)
*&+S݁ V&e>w7��,�ig��� �}d�2{����7)�7ç�?mg�g�p��e�Ы�޻�&�d��[�0w8<�����<�Ճ��!�â�j3<��d�ؓ�c�n�����Ub�����V:��� n��=c�ȡ��l�9��.��}8S���;�uT�%��s>yʝ6N��'�Xx�G!��o\N5���A S�f��l���+��/��!��ἙECZ����;ؽ�秱��O=�OT��o3j�*��\��L�������۝��n����t���W.�Y��~�6њ�]$*$T���;A��R����4sA;����c�`�F��b#�Wޏ{���g�������������K;<�i-w��7�2�"݈�`T�)Uv����ļti��n���<����`�7̞�U)�o>݀t�ڮ�O��+��Q/]{C/ݐ�h�����*`����{'��+�Oc�:��̊P�-2�P�b:6*=���*������h
��{UG����u��r�YQ��C)�.�X>ߥC}5*�����JF���ѹ<E�v`q�@���&V���c��bѩEW{U튺���^�m�$���81ی��8�-��p�i}}F#/%U�3*�^��(1���J(�/�fj�A�^5��\�bh(��n+͊v\����]i�T����B�M��R����z�y��{�;J��l�����c����ɻ����׎)��@[�[$��>Z���!/NY�X"�h�y/Ɵ-��q�����F;n�횔�8�/�x'�\�p;~ő�,m{2�+�B����青'v�
$G ��:�0�Hc"��ۢ�md�A�� u"�Fd����}����Y���[��u�ȪѻzE�TlX<�+��������s`���N�����ż����ۄl#�a��}:�R��)���u�*�.ms��Ӵ�0l=@t�0��>p�5�W�8�ѐ;Q�դ���f�N^>Y�����fk��*;9=�|y�m�+��;}��1��F����o��=�n_+#s/w��0������)<}�C�T|�+-�b!�}R�M��8\Viq�9�o4z�_��Y��x,:��JY�
�������yE�z�ɩ�F���gW��m������~ۅ���}�8j�7빃����J��
��ä�:�������GԶ�x:�X�KsB��^8YpG^wM�z��]��ۿ)����oL�\"DjfV�4����=�z��c"rv�*���O��ޑ\�Ň�b3�.���8v+ts��ۘ��/��Z�3�%���v�P�$��h�hmC�5���OA�x�̶�4���m2�ޖ�\�I�J��멲�p�L��5V\�D�[�i���~�'J�9�Yg�&�v������Z��K� wj�Z�{(�t��ǡ���uv��\��|�K��Jb����G7i�G�z#ވ�xѝ�kZDN}�ځ�yqE��U�e(1ۏy�)�I����A�PCt��\�5#ӯк��X�=���*��7y��p�ά%�K�G�I�ÑM�2^�U�F��-�����}w��V�t��^7�����]$}!���{�'=���=4��=��i�f�69�;'K�J�PT,.������!��|�_C��S	���[i��ovѱ���NRu'.5ꇅ��̦yoo:ծ)D�� {@��|�&��1�ο6هD>�S�t�m�*1�F;�$��.��L�:�u��yhU�oh����\^�.�1p�����;kY��B�:0v�<�uq�}g�)<�|;s=��2�?>�/F`w=䆆�%?����ZJ��q��E��r�=H���T�Cg�1r��Y^��,�ߧ!��-[vi�l7p������0�ৰ:��]�!  .��t��;뿃���"���<��m��3648La;�2��"z���p`61[���"�(J��I� ^�m�"e^�wY��0޸-K�4�
�{ј����hm�%��{uL�s�F�F�[E^EޙDܬ��{���iGo���l�Ŋ��)g-�x�L�P����+5=�Y�p�T�>j���e��?U[����Ʃ�xhM���,�%�P><JQA��M�m�Θuv�}l� 7��Ĩ�'a�wUPuk�{6���$�3�~7oeC�C̣Y=���I���(	5�-V�ΗR�\�M�
+��#Y��N;�P��ӤpOs�b���{�D�D�����:�X�W;�KJ��_ yZ�m�w�zţ�yAc
�՞�#���Ԉ{�Vo5'!���YԣF&����M_Q��f:/	�X7���E�|yS|o�#��)���85���7i4��ې�7n�>Ӳ[[ƶ��[����K�v�x+�v+y�E�`����E\kO�y��+>�X:�ČKKȪ��ҕX��V����}Z�1�&e>w7�kq&�fN^[�\$���;�^���&*%d0�D�����_UݑZ�=��f��y�y)�\,#t�>�8��M=��������w����Ԣ�Gϥ-���/�4v���f%����:6^v!C�\X��E�K@��hI�W@]vU��s�����DBe���n���ѩ�z��*���f�uD¢;Y~Z�a�L�����ux=�<�<;$�,<(�O1� �~k���� �i�Ή.������"��!�Hƻq��Fxv���Zsgʗ��r�vn���[_D��zy�b����Ta��ߋ�R��c"*'\�x>�ˎ=rc/ty8硋½�(*��M���a�`-u{8��eS���pa!�b1bTt�9�Zڵ\��n�<��������	u��%㥙�YP��0�Z��� ����Z��s�q�>lX���ZHk+�Qi����{(`��[���~Ua��`�N%�OV�w;n��u���D͂�#�:�F�P�'nd-�+Ġ�����N95X�%mu�Xe�����/��п)!�a�OR���Vh���u�"�f�֎��P_<Jg��v��-�=U�7e%��X^r�=�XYՑ�:ll�e
b���!��Լ���*���8�0�+C�`7���k���C�lٱ]��ϡ��M��;�i�ł��N�1���#��p��b�yI�ua{��z� ��)c%�qQ���t}L����h��ws��j�k���%��o�y�`��s:�\�՘! ��U`X�[�k,.��)�^r�\�/�"F,�p+�A;�}�"�����i0_	�x)�{�rn�\!|�ꬖ�b5��tL\u*b�r��5)����%9��X��h��[��D���N�t�2��bٔ���W2��v����ݙK�պQ=E����srm=\�ѡ�4D��-MѤn���[�
���hpVb����������FnI�&�ꆰe��,�}M.���L��e�����eVU�G�(=�u���v�<�w2^�P�M�t�S1��箛8��j�jzw`����k(�]2�mtYx�l���tw�����+L����S�Xy7����ol�.V+{	_N�o�m��,�xr��L��!p-Tt5��4���#�N���]oV\]2����P��F����:����g@������iW#˸��N>�3�fc��|˔̡w+N^qƻoV��m8���)�O
R�����}�ҖT��%���[�8�uk]�ݭOW��]�i�/ lҗ��dT_Ϸe�WK��Gz��ڰ5�K�|�KN/j�mY�|jqI,J+�6�F٦�Y��^�|r���7o������ȥ
u�7�[5y}2]����*�R�"`2����+;'Z��2�_gF��W�	ك��/�k(?�N���[��He@6K�e��MĞY�����GMnm�A�gk��A�!��b�(��Y��XJ��5w_oʛ�U��n]ΰ5�k��>^u�enl�K9�u^3ɰ-�0"7%�7knWe)���qQ�&��+��5򧗁
*�:B�j���|��KFg6�L�PV�qdij��R:�/������A�cU�rHmt��!��g�a���PB[���M[Z�m����KJ���t9ѭ*N�yr1wg1wX�=i�jp��%=4ۭ�y+!/���`jb�j�5{��l���k�+B���rH�uu��	�ܮ�!R�m�2����ZFﳏ-*��5TS4�u�[�%
F�
2/�=J����;E�>u7N;an�RS8�vJ&=�pXvþ��{�U���&0�o�s���i�[�����D��)�ˆ�SX��*ٙD��H�N��ᮂ�@[��ӽrZ��JG$<e����>�+eܹR�a��z���ʖ	���QںI�6N�D價Hǐeɣ�f�V�<XR��u�Vؼӵͽ�tD�{�j#)v���xr�F;{h�}E�]�w]f�Ň�C8�ᗶ1*e<�B�ǩn)�WN�&c��6���\�ޱyf��S�a��)��*��1J#Ke+A��eX��UkLc	R����R�H�""�TY�,Tb	�T)ZEb��[��dDX�J�UF&\%VZV#"��*�����UJՈ��
��QTQT�H1p�����T���T`1TV*b�ڴ-�0`�Z�b�ڢa**��\%b�Vč�V�JYQb0b(���DVڂ"(��V"1�Kk�kT�TF6�0�)�T�PTT�mf+j*�E��U�cF �F"F��Qb�[ek)KF�ʴXV��TE�( �Q����Z�F*���m��*��[R��,QV
"���*"��-J�PTQ��V5+iqj���)�����Ţ(*�
"(��JZQ�e2�Tؕ�h+b�b0E�bZD�*&,�*�F(ҶU���,EA�U0�0� �DDm��*��1lX���
�������*�+Eb"�mDV* ֌QE^&�����e�]*�&"�%�>�O�Y8������b��wA�>�f�O���P@����0��U��r�]�.�R�U}��URXڗ�>V8u�Q�*�w�2�.�����beL�u�zg��_gYu�L�^�Dfɥ���ׂz�U��VLW��K���~��܋�Ӂ�4H��E�1q�;]6�[�;xRKw���{Z&Z�tK:)�<*ʦ��4��%��<��);��0d�fV���<�ث�]��j}=P�K�:'�H���t9_���e���H)��IyQ�oټ� Bt�)ᒙ����N���$1sםl���K��)��Q���1Lh⩻�U�J��k>��Y��T%��Ѯ+���y�!���Ī� �J�j�9�gT�ޝ�RKW�;��!���T�W�8��	Ԣ���gqsY�Pd_�x���x��ti���\)��M/4tB�֐<e���P�B�S�6�D8˞��y2��b�C�n�qua�G�?L�?I��Z���ΐ�|x���<�tT���Ҙ��<�<Z�w|d\�=m�{GH`����vIx����}��D��`�(t5�X��r	�ѕ��j�;��秇���(Z��*J*��ۏ�Ɋ�Ŗ	�j�sA��.����7�P���rv^b���_�	8��G"nF���VyG0km�#W��d��ˮ��7��������f�qh9��� Y��:K+�Zc��W�P��I��̀p�U��v����������&�_N=��%R����J��D���E���.+Ԧ����h��e�X�rc�UT��љ���z넃�V�s5OW|g�(a۩��'�h�ő�&�f�(��T��S��w�r��q�z�+����5M��09E�%��ώ�����-ڮ�^W��x��v�*�xtx��V,g�n��]gAa\�.+k�lt�vM��i���%e�������C�ʜ���3d�]z��(�K2��v��q:03��	8� A��\��kF��H��-�Y��	m���ߞ���(X9�T����m}�[�y��j��o����
m�r�l��:�A9��xcvy��kG��0��񒗝aup����&��z"��2��� �Ś�ET�pY���E\��	��?/v��V�U<�Y�`�m}��x[K=�ѷL�Pe���;��l�o�r�|�(���+�d'�?&Lîe��N�eY��C��^o��U�Ս�r�;�US3 �d���	=�ew�iE�' \��qL���=�.���k�d]؝����j�D\�RtwA�cJ�톓zj'��K\��m�nf̂����[C5%wꝲ:��TݴwN�l�z��q���u8C�+��fb�Ov�R��TѮ�v��[BN��}�7��!��k��]��������7�DG�#��d�Ji��'�2�n���)W���iF�����.��ӕi�ezvP�Ttf/M��"T�9�'�ڤ��!�	D�	v��R�/>�v��R��R��u�1�,b杷������F� C���Fl���k�#��@���8�'�e
�e��pWT�橋Ǳ�y}�˳N]5���c!�/�.S7�b&�6O4�>!��B����)z� ��g�K��Wy��{=i�*���EB��GOg�<�
�..��S� zo��s:�_��l�,P��3bX��gK>����]�8�kD�&����폦�<=8g�M�^k�˰�=M฀�.��u��W�烬87]����+�(����m��_-����C�W�&����Y��=d�虍�˸�X��^g����6��v�=6��:MI���X6��)�*���pn;�¾�ܓ�T�n�ו�G�J��q^P�^}'1/
���G�ᘞ���"��n
=�(s���hg�����k�m<��/ ���2�V4[�6t�t �{zq�M<ۭ=�� 
�Jn��Rdcx�{Od�s{ ���ǥ�+9A�G�J�t�szJ��A32#��4YU�,%�.V>]���\7oH���t��nH.��짛&���@.YI��������1Ҏf�Ghѕ;1�n�beL�cv���7ї�����W|�xt�mc�H�Y�����o�%:`ޒ�_�tC����y��T1m;�^V��u�F�m�+��^1X����q�I��.X����*� �/Es��˚�..�?|3��ݒ�kY�/=Çd��*�W]����!�V��V����o���{_o�����Kay��oְ띧Z9O�=º�ٺ8R������;���.�<q���3��Rst��g��-���Y=O�]r��c;��}6�y򖑆��m.!�	�T�vQ�sk;�ݛ���*��{�\典��0�#��{+!���<�p�����*�������3����ݭ����R��s�:�4�oǺXyṞ̏�1�\%�����/'U�n�K�U���[T��7�^JU���+ǅB11�(�S��ƴ�^�y��i����{Z�F-�/3����媠��R-%{wX�]]r^7��ެ�p���ct�ou�3��z�B�]�lu�+o���s&,<���do�{p���8A�
����#Ҧ�ヤu����1���w���+9�(��ӯ�z��[!R+'|���o4	]*�+ܸ�N��.m���K阗�;��_W�}�&lY���U�����[�E���;���՜�x����5�֦�i��2=t�g�����n��gҩ�`�)�9*��0bU�aߺ+�d.�:Ja�b����e7�������Ȏ����������,���V0��g�vQ��C�h��"�S��n����2�>�7��cR��,+��"�ά��E��~P�7F�/\�Z�>�!�L�}3wڄ3���V���7��Ō���˫D�pc12�W��9�'@�q��/� �/ۖJ���ó�ߢǃ�D^>�X��"�+Cr/�Np�"2�hL6k!�r�.���ɘ:����tӫ�����o�c�C�딄�ݩB2h�����\f�s6t��7�����n��Pq�Nʽ㙇�Qk�b�u�3�g^[Kօ��r��e�t���Xywr�Ǝ1L��2S1���[+^c��_�P�7Vژ>�C��7q��:ٹs��U���0`�Zy*�R�'��<s�	���ol��fV���W��,[���L-��霮��G��R��p��1�tl��"�6���vw]O��Mpy�Ed���9��|�.�W^b����k�F���Ҫ_Q�@��Ry}��nآz#{�.�ޅ�;�3��*
�v����Y���Q�3��뾕:>��2~��z#ޗ��,8����3:;�T#�_�A�5x	Ԣ�'�e����(2=,��ͥ~�"�t}~���S^P.�`�W�(&f:���v!�Ӟ�F��{~vuN\ޣ��Tu��Q�fJ孎��'�������:��P�f&�ܮ����ʫC�_t�*�1����y�mx��fq�c��X��`�+��J�=]�P�z�TJΥ��ւ��dp��.�W�O��BBY�X="�1�S0�r,$�)qV)M]yv/d:�t㋃u�q1U۩#a`q�R���bA]V�9
���N(���a�>�wa����`Gbb���+B���=��6?*;�����ÿe$�f;��1ʘ�-ݰ\E�R>0�P�7׫�x��I'��̠�n$�rjm�*  �r�i�b�s��kmC�)%�బ	,0o�+Ի޹�Y9ķJ�bR=�&=^w#�l����g��s���z�<�C�~�<n�my4l�����'�#|�դ�:e�+������R����8���z��>�Ֆ6�W=�)p��=�[3}�̤�I����+��������C���hQ��2�.�:��Gs�����gի�u��Bd�3K� g��|4�
���W<A"�rk%��w�B�\����>|V�}{��ܘTW-�}����L����G���)o}�z"=�=��U��[V.��_I3�2-�Fd��Z:�ő�=���Ͻ^k2��W�.Q�l;(��܂���̽z��E½\^�[�����+ݾ�k�U�'�;�m��z<���N1����/�N:o@N�b���ʕ.m'&��c'�[8�5d<�=��獿z
�:���ج��|֯%���T̩D���&�ԋec�Q_�NBal��|)SVU��u��ӷy/���#����-�MQz)W�.�J4��&�Ԅac�v�Gy�K�w�?gdwᵔ$b������VC6�K���j��/n��r�?,��=�q>�ʥ�,��j��y,!=[h~V�f�مڰ6z���fbYdp4z�P���}i�n=�����)���-�T�u��žY�1�/&�-�.�.���`:�D ��5淒��[�o��ݹ*� v�x�uru�U�>P�(ӵ��C�L�#ʽҧP�����*�>�^J
�D���	�c�];DhC�6�9
���N������b�z��Iy�}$�'rU�1��H�Y�����Y���)j��7�`s�h��	7:E�4�H��b 뱊�*�O�����T�gK�뼮F��wQ�_�P���U�:����gh���.�@G#Եk���p��@1�)A
��uoQ��u)��գ�G���E���g8�[?�L���Α�%Z*���#1t�j��3&9a_���.7�*���R�n,���w��P�}��9%,�����(
�b�p���Q��H*�~ѿ7�'F�I�ܴ�ۿA���3��R�%�X� ���[�pME�
�A��;=i�z����T��sk��(�K�x�>�,!=1۱��z�^��ȿr�f�2#�3�a�~��}#��G��p�/pwj�Ϳr�E�Z�tˋ8c��X��ʙ�t��38��xh>�]�+�����mhͯATΥ`c�o6���Hb�z�5�КK�=|�v����r�Q6-'1�������{�5e��X�bՀ���܍�V� 5��]r7e��Ǫ�x �}�qD�Ǭ���/l��⋿��bF�M/�����N$_��'�d,�]��k*K�!��ktz�5�I�Fz
z��D!���MM!�v)P�U�t{8,`�6�W�;��������1s�4�\�e�5�OR-�il.5��K�v#���z�'�?e�.�}\C�:5x�ȕN��;H����vq�r���d�	o�om�J�'�R����;I�Y��.�+6ڭ�HA��3����P�ua�,��4�f�7q��J�5]��`{iu�v�C�V�&X�����f�z��˞x�M�&�1�DV�2Ft��!��`��VE�����n)~�!dP�J�7��)n�Xt��K�Y�Z嗾��1x� �YԃN��ܻ�|{�6'�圙P��0n,��>D��7i{��gdގ���&���z,"��4�הz���[�k��ǔ�`��kW9)�N��8w�()��s� 
u!L˞�c��* Tk�p�A�VD#���^�@I]��R��U���fj���P�(P��������%b�q�S~����}f�4�7`o�ރ&��{+�sk3�h�
|�	B�D0��tWd��Ӧ�A�\Bn�MaC,c/�n��P+��Kƀߔ>��Ϣ���৩`��ە��,�BoQ�U�zd�T_^�b����X�W���
�Qȼ-�7e%��XW�2�,,�ϣ�5��\t�,ͳ��]�kH���2�Α:md����{kL��H���`���J�\��x��_����ޔ�����\e��!`~En~-pى��x�O�Osb�r���[�`� y��[ۉ<h,���m�$�Z2WU�s�ʷ�	�6%��PZ�>"������2�QXY|����u@��y~�����U���m�Dufi���rʕm���ͱi��u�5+�ݘ�`7���J�sW�؃j~�������77˟�lW����c�ߌ�e���9��]�G�w"������I�w�יs�D��N�����j�fr1�W�g����\��*w�cx���Pm��*;�i�>A���a���mvV��J
\V��E���T�`�{�l���av;̐�BP��V�s�@�4r^Jw&����dJb��L��w�D���}L\Jg��k��uƼ��p6�SӏxKՃ*�_6�-F|T:�}UL��]Q���8���D��}�C��c`�Ȭ�O+�8�5������>٘��)�g�@�;��hxu;si����Y�Q��V5�`��k7�^{ط#�A��Ǧb����l'\^}B���SJX��<y:x��-�lڽ8�W<��s�Ɔ����`��>��AC\��z�
g�eD��[4QF"0�)�v�y�oϗa.�X��0�Z��p�d��E��_t��X�5q�[���6�;�}y(��fEd���D�os���Ց�]�^
�����Id�F�@��j�a%�Pr�j].ܽ��q��4(��M��зC�<��Q�����賂���D�3j��Wά��ӷ�s�9d[\��;��Ĥ+��(���Ems�w�|����9c�]��X�^�N��]��
�4�w�qT��\��x-Z�9[����֥�ihu�m��A`��p[xf$�[*E���))����0���N��r]nf�H�щ��EM��,ni�!�$IDn	Hm7��#�b^�i�yC�|o:pLn�E\��ʘu�V��4�0l��X*��q��O�b���	�y�l���S�6d�!5�q�E��Mr��m%¢�`��/2�U���YR�މ]�c�$5���Ȫ5�H��֊Ug� ���@��P��Ry4�ܺ-�|ܝRK���vPLGY/�7}��!�����yS@Y�6�Hx ���n��z��n�>��aّ+����g�{f�D�������R��pq_wZ����T:�]��Rw�4cg����Jܨ�;�B��9\�t�YA��f��Xkcq[��mH'@+Ce��%�Y��A��ɖ��Z//&Z��a4a]�7���3��ɠ�j��X��wzR�L��,Z�n��;��T�v@���J0z��}Ӷ��{�z�������mL|q�lӫ�}K�r��b�,�_F�퍫{�Ί�	zI7�&o�54TX\s�f��ɼ��oHW�P=S78#o7f�KH��܈�C��b�"�\��}-P1��֦��*ov��-Jn��m;�����M��kN��wz*�i��N�;@ח{R��[�y,\,w�$�$����;�7��6�:պJb ��V�ÛV��f���@:�,�w�r�O;8v�ް�N����[�L�c�劶n��WQ���t� �
H���5���E�$��GY<���p��7��S�΅_�:XQ��tL�L�6_6�̨ͭ:1aÙ4��a"J�B�n��H��duAR�5��r\9��x��wM�RR�d�þ"	��[4-�|+
YE�NP����wU�����I;pT�)�Li�z�����+�gD�⨍��&�9�S�k\���S�]�oze�iv�q�bae�W`�Û:~*��
�vlՈ�nI�v��o!ui[�ڏ ��&M�ti���'&l����Y�W��8ձ�e�)�����W,�d�얈�QT�r��yԤ�^<y7[��S(b��xFk�֝j&�dM���G���cv �ѷ�CZӜx��`��w�Y6���j:�C�fZH�N�'m�_ss�iͲ��٘�K�r/��7B�jys�5�1�#{�i��VV/{0K�L�����-ռ�?N㓕ug��f�[�idyJ\��R�Y]�[��/��V��p���;]�_d��Wڂ�.�;Q��f��2f3Z/5��Ц�r�ը1.Z�9[2�%Yg��+��D�<d��?f^��a�Ep�	?8�J�*�E+b*��H��*(�����T��8e�*ԴB�.�Z-�ň��qlEEQb4�+�PD1h�"++Q�Qj���"""�Q����J�eZ�H���8�b�
�h�ڢ�b(�Ŕb[
��֠����`�(�m�1-���+�F 1PUX1qJ���E��-PQ�jU\5U�TUڈ�ت*�(�("��PV�`�1E��(ł*���X�X�mc[J*b�U��UETA�&
#m�(�a-�V#Zp����+U�a��*1DX�ŘC1���*����QҠ�-lU\5m�"���E�AX�����B�Ec�,X[V,V+-�QFڨ���UDF҈Ÿ�b�lUU[`���05EQb�b �C	(��ETTX���E"���d�+
�E����U���V�"�4�J�E"� �"�Ū8j���l�+"*"�X��lh;6��-w�7v���p���{ܷ�T�T���[��s w]`|x��T��z�����X��WD�Tn.����G�ݽ�V�s�#.T��5A����=F+��L	+��Bɘ��(���F���w��O)\�GzA~���.���g4�Le��\<�L�:�3���Z࠷�,0H�=�t/���8봍^ry�p��C����<je�ch��\�1���<.��4��#;0)f�MޮZW.9� A�eh��6y�W��g%��Q9�}.����RDeK`ԛ�S=�H���)��I��Y0���j�R�q~�ym6'���a�}^@���{i���Ϛ9�i��#�ZDr���r����̮�������N^~j��k<)��C=�ﴔ{����:mv�AU�y�w�53��S%�λ%C�Տ-�i���.p��:��#.�i�)Zܪ�q$����@_T$��-���(�E9���$�v���TX��ɻ�j5�uF�U�KR�,�VZ+��T[��4�҃!������^g�j([m���3:����M�������m(�a.�1���s<�BG�xժ~κ�]�t�u p��w: n=Wty�{)�ێu�����O+p\,o��ô&�[����Eه���v��T]�Z��������w.U��N��]�۫(hUPVI��C���TV�q�#w:;�!�v�tv�
QV��%h�ҕ!�~����It�Z���f-�BfCy��
�?i��]��H����c���i'�e
�\��
�f��k[[����u<��H��]-�̱�y7�l�w.�<S N����@�&u���,��B�5c4�^�Χp��%_��&���5J�"ձb��7���x�)ss}��$&��%�\��\1O\�Ӊ����g9�[qn�w�F�O`"�����ㅭ���g������"Fß/-�%�Yb�8�qA�ȓ�|X[\,����.z���&�;�Ԫ����D���K�L�A~��8�~J.9�JEa�2<039w�=J��ھzf�=�<��Sf�*��6�I��I�u��Ѕq����[��]{ڬ�UϞ�ۺ��ԉ�;/�8g���cx�1>dh�=���2){&Jbm�u�P�WS�&d4fu#Xj4�ӈ���L���6��A��Ը1:S=�
��h�b�%�,�d�v��q-i���'�p�\���c~�cuj�[�R�f5I���=ʅ� ���pw�Y���5�u�xr��qͽ����KE��á�6I�T��*a�c�LB��������D�9�V�@εX�>�I��	�73�a�)�����.��\��ͦn�ά�n�-�sV$`��kuy�:u�}U��;�;g�[�4%60}�&�����:�&�S��-`� ���Ky�曥x��]ŷ9GZ�z��'+g3Ñ��~!�^V,�2��VS��8�zT�_r;�t��U��.��[~/�����=A�8��^|��4=��C���Ug�7�"⯊��������O��Squ�g�hb�%>�25�=U������<ж�'Er�J�噪�˃�9�贎���n
vҰ|�3|�F�p�{+�A_<�^�wooޯnZê��oؼ�:|g�4���v.I��Lܡ��yg&T#/>��nGCF�㲰Ҏ�˽䫈V;3ĚZ*�沂d_����P��߃kEvy;79=o�Ev���~��i��֥<&I�@��imJ�� ���z�Pk�p����:�ݑ����J6�I,vzPfz�LA�`ø
����\�k���w��53��AyLQ�r�*
6�{�03i�FB�Ua�n���
z�	B��dC�<&��»��[�Fpbצ���\r�ϔ��+l�8痫�˯�e�;NE�wƲ�#u�ŴU��L
o!�^J.��=D��7�M��^��_:�����m[m���+9s�6,ѽPIܬDl��w�޷��+�viD�{�R�C)m����)�*��|�P��,^N$z`J��c��}��)�Q�>�Xl�jE�4���{��v��r+�������f�b�J6�=:f�1�7����e��C�l�W#F�@�r����(��uV�"��.p�A���/j�}�2�.���pc12�M��W����Q��W7�4�U_ �jE٦���T�+��ǥU������k�B���k�Xqڋ巛����)���4�q�Z�2�f�-b>����)�x��B�J��5�Pv/(�d�f��ҦYgG_����х�����1���`�=	�#l���5~�U�D��s[����1�,���2�\�t����,
E�����z�N�xX]��2C	C
��� ��kEy�˹��]u��YR�f%_w�4��E�.uB\�i����k�A��]9�e�=#	�I�x�Qx�Z*���uDrO�� ⚽:���u�	�)-�tLv��v�,�cb����1r-"ƀS=����Hu��nmh�q� �PK;�^җ��ξ�q_G�N@P�6����1;Ycr4f,��DQ��˅���� �U�E���uʕ�� ����ޠr
�8e��@��.�V���[ի�G,����s�)�;Yq�`�i�롸�vUΦU�m�6�*�pm��T��1j�:W7D�u����ﾆkdO�xcx/�v_9[� �_�(��zf lrip7�u��
f^SJb�0�|D�SNMC,���+Ky�n�Jp����)��L�9��dX��]rW�'���3�Kvʛ)ĖҎ
~�����3��V3��Wz;ӹ���.,m�;�8O ���j<��/vor�����ӹ���tޚ�W�]�k�T;�����6VD;�5v�80튙�a��|��$ty��=.�����B��)�6����J5c�e7ƀ]���d�S��u#�Oh�b���4�zE���=T25��l�֠*C�a��8YW�,�R{@�մ#e3\�u�=Qf�i��oc~�'F�p�N�ע1��Z6}>��~wt����</1>Gn��L�b����-����A����I]g&#��;�}k�jХ)N�n�����σ�w5:��v]!��ul�4'�ڲ��E�^[M�U=��r�R�+ܲ�a�w��T�k�Jt/�XK�_cY}/�p������R���৩�	�d�Ƌ�Ռ��s���|}�߬,HV	|eq�h<p�X�-��'�Q�~Gee�U�ի]/!6L��k���x�9����(��܂���!T!2J|j�_j�Q}���Y -��흅�VuprZ|.���v�X]xs;j*?X��|jΫ�cGH]V�u�5���ZwяWa�U�������jV��ʕ�S2b�TW�T {�58�S����ޯ��ZUӱg#�5Uӕ�����sG��l^��Y�p.9I-��T�x �m��������8�ܦ�GT6z��������6����ֽ"J�b�Z��`�&:"�t���D�ć�`U�WQ^��s�f⓫�.����R=�?hNt�]�^���*Ȅ����S)WpiC���y}�û"��&k^�)�*\GS,F.�C;\y[�3e�d�^Z=���#A䞨5�������|�+��N��
�<�:���O�'<�y7��P��r��>�H�_��nK2��� 
�f�w���3�ugé�:�!b�:x�=�%�H�s��W;��E uO{�eC~��`��%�µB�d�U�Qi���X�;��I��V�q�l��[�7���׸�bGbrυL)�����y`�\i:K���9��(&g2Oym�83Ers���雮m5�Ϲ]�y�G��)y[yw"�3,_�J�4�n�T9t���g��p��Х��>���4�H�}e͇w�UyŮ��*��qBa�����o������:Cv�Z4i�>fֶ�W��=�׉�z���XPC����بܞ�&�Fj��b�ņ�,n��t��7\j�-�%n���c�N��4���'k��.@�8�S��@��,w���]�?S��a�d�LƉp&I��X�ׂ���� �V46�;=iӻ/�m<�Gp��l�o����^���Z���^ꀢ���D��r"��d�LO�ź��Wj��(��2����fS�΍őF����&��2���(87ؙS8���cG�v�p�ؙGSjU!A��j�mbL�[��ͪ�������kt��_���֮�{����[���F�+a�-z|�����r�s|�7"�2�0�epL�\Wh��-�3��m�J��E��	�d����W���p�e����r.����	�+5H�8�`Y�}ϴV)��1-���M�}8��^�!�<��C6�N�P�F�;g��n�};=���-I`�m4�Jfzm�$��0�s��l5�OR-K3!�º��Q��Y�EevVc���G�DH�wc���V|�3gZ0��VC3�]��W�.Bz��jU�y�G]G��7�4lǉq~]H;�}��m=Zr����reB2��Ŀ_)�hU ���Z	�R��:���VemNɜ��-��)n�.v��U,b�T��]{)�
d���(Ճ��b:�i�7��p�@���`��|u���(_3Vu�H�_�����sq�z�v=͏pus�Z���.�$�#+x��K��j�T�(�t��D'�ɪֵ1��� ��|pk�@۔�V*��,��A�=\�/�\��+#�(�ӧ[���siV)~Y]sYT�n���ݙ���8�K�G8߆�T*kI�_��]���5��(^�ںA7$���a��eB,,X�yi!k5�]:�/>����UMM
����3�̨`�a��{Α�a���ma�OQ�BR��o��+�VD%�=���1�r}�k�/��@�^�/'��&Nu�4.!�
�qKfm�#K�1ގȒ�Vp�t���H��r2�F��e�1v�歴,n��o1a_��6Y��n:\���J�y�u�0z{��#��qzʆ{k��3n���P�Hނ�yI;B8��Y����<�==�� ��w�{oc-b=>5R�t�X���&'�O�`n@�8q�q:�w��\��Y"3:�(?G1����Y�Y�N��P���.��D�7���
;�t4�>�:�ti��i���a������>���3�r�4���G�a�٫����%K�"-��,�Y�s�ܴv��kw��
(jq��\��kT�ǐ��a��k9�:��VhΦN�l�*�{W�:`6���h��~��O]����7�WUݨ�9_꬞P�g�Sݡ��pB��Ӓ����9�������^�sȺ�*@�����%�աi��*f0\=�{|��Ha����m�����QR�wi��^�ȡ�(�	��w�4�=�YuC�9|׾�+�tq9���J�չ����GP.I�(h�>��Z&}uDrO��܃�j�J+�}�M��gv�gr�ɑߵV)�b�#���<�#,h)��(&f:��U�,u;spt��ם�O%�ϊi��*_zy�w]ν��Ս�Hv�b�4�:��P�e����ͷG�#���)��I�u2�R��םr�1��-�Ȱ/�KC��J�=\e��ջ������t�]�Tq�
�er�v���ì�=�b��7�Ԩ}��`_�̀#.3�-7�F�V��}��'��٧�:
��D�n�A���Y�:��H0���vyI+�!8�:aX�c�6%V�V@5��U�d ��2#�n�;.�����>�j���0$���+��^��'/�tma7<�s#5��g�ݬ��F�C�͟i��6�5�Τ�c��c>�|�<Ԣ���V�"�v���y����'���a�`�Q7��
͏cٺu6�ƫ�|Ȯ=�ҷ�{P��m]�%�oR�غЦ8X���0%}�`� ��ə�4V9�������a()4�n�
�<�:쩊���R�B&�Wʬ�DT=Ɋ�܋Wpʾ����6�G5���5�Pr�S�8�OK�$�YS��/<���ס��P��sMpjY`Vc��`�H,fw&��'ei^�����^�,P�/j��*W��ڙqr#����?r)�}t�zI���ǆ����V~]�"���l)�wW�r�k����Ч����{��X�/�2���E�c�F6M�������ep[��p`NV��,F㳃v_#��'L�sλ#�ܑ���<�xw«m<�gR�������Rj,w����|Kz��>���%�q�a�٩ڱb���a��Qg	���t{����������y��~�����m�7�~��8gR�ι��L��B%˰b��Է�>�VZ+��r���4�S�R���n�̏��i�|��H�Ӽ/�9�͂�z�:i��	VD$ĸ{�u*������8%w��(K�L������T��e��-[�3},#&5�������2�������٫�D�5��f&~��P�WSɿ*e�Z���o�e������e�K����9JXǳS�tm3�A�
ӣw ��ŅV�&^����g1��8�6C��ܥ�_��<:�ͧ.���L�s;��e��A(2˄E�n����N$єk�F59��y�	��r��Fʺ4���]�[Ud'e=�1�@�� j�(Y�@4^��W��vn��b�`�C'IR���8���,C�'_V�
��CQ|�!;~�w��-��t�W-����"o4�q������ř9=NW^l'����wZ�Y�-oA���V!�M���tMe�ٚ���w�5ά���^��g�D��%�JI�b�H�[�rKU��g�/cR���;ԍ��eh��ʲ�����2m���X5ѾZY����s�T�T�Kb��T�gjܳ@XG�w�r����FR�b�nhDj����Ƿ�Q�ί8E�&w���y}���r��b�b���<^�S�M,xy�ɗ[�59N{x6�"���6UB�k�y���Q,��N���b�i��ˤ�E�}�y9�Wκ�ep��<��t�{�x�5v��̗]\����Duh�k������2�ɩ�t6ɷ238��e�pn�!VmY/	�\@rm�R�X��ٰ�RR�KQ�i�w���Y�]�){k%6,��dzӗ��H�M�^�yguw#CQ��H��Q)��c2�G�R��v�5�F(�"�U�rU�&3׷�cn@���d�K묮��5��M�wL��Kո�������
�^�)&nV�jb.�S��=Dͽ��qfNr1��N�lr�<�ژ��Gw���{�jͦ�b��o0����n�2Lk]�������*��&Z՝a��H�q�Z�Q��wgX!���W;�V��Vt]&���9V�e^�ҟo&��j�Gm��yX�A��[3B�k��qd�%������Q�j5yf�.(��;���_n��5Ä�S�.~Vi&C�n����u�u�A
���l[��ݾ��������塨��RJ����j{0�-��_kD^2vY�ŵ�`����d7�/�r���6"����ՖcZSv�k�ͥYl�˶K3,�CD�M��	��i���ި�5$��N���vP���W@�H	��3$svh���w��%b��rOXRb�Ҕz�k���N�,.��88%(�3���՗����!v��2u�D�dLv�W��9m�拭γ�\@oZ��e����I(\a���/e�Y;vdz��e�D!�Z�g[�{��>��^`D�����=	M�Һ3����f�V�'VD�qp�F��7��[��#v[�N�^IV�$��9�r��Cnh����;�~|0�Z� 1�n��|����d=f�d�b��K���.���C�;����\9�t%M�)`|�3���hq���lLUˁS��J�4:Vso'l��$xʾ㹻�}LօF����w"�m�e�3��K���f�����	~��^`*�j��)AQDUQ+d`a��"a�UYiU�)DDQ��2)mEU���b�Q�QQAX����EF*���0����X8��Q���A`�1j1��*��"�UDETe�[J�U��������"�+��AF"�**�QE�Tb,V**���EF,UA\Z���(�DDEPAU���cEQEU"�UUT`��"ň�(�AA���b��T� 1DQVEATn1�T����,U*��DF"*(���E"�TTQAQA�(�"�#EQ�XVU"�(�
�b���E�EEQV ��Q����#Z�1DV*�������UQF*"*E�1UH�֊��AUE���b�"�Q#AQF1E���("""��Q"����1DX(�$EDQ5��_c_����7>���V:ý���eg��[�:���k�ΕG9��b�[;�ޢ�1���>熟d\V�U9�����Ǩ`�UH�!�fb�9>�
��'}N�עU�T/�t�v{3(?I^����S8ev���}Η%uL����4�W-�:Yݕ���:�Cǥ:<���!�pQT�T�^�S����~���.�ȍ�)yh��ᮋ9�*-�2b��XOI׺����;���$�j�`j탎Q#A�$��&]���ZG�}�z���3>o�;�A��bՆ �s:w5:��X���2$�y�m��L�b:G�'��zאx8V�t�?L�[��x�K�~���׾�y[�/Z���Z7���ǈ��bz�}�(M��f�M��MT��Y����;Ո^�4\��9�S���g�;u~3��X���g�ј���?Rŕ(�j]�7�6���Ձr�*��"\0����T��BU���V�xž��p�j.ʞE�v��噧��S���}r��yX����*����\�9����nV� Z�V��X�S��SX3t���	�����l��xvB��B&�"�������PԥU�aX�����w����[�:� ���܉�9�2.���Nf��T�$�a+�Y[��'��s�Hܠ�A"�-"�gaZH=�5�h%pGa��t�`��<Ҏ�5su��L�<�oR���Ze)T�&_\�ږ:u�y�w�z���|BO�}Fi�6=�u�꽙{���o�Ke>�yS{Q�q���"��y�&��Ԟ>m�׸u�f�Ób�����ޫw�{8MC6u���0�Nv3킦��鶋���a��y��%$�t�puU�m�kA�%w�DlU*�xS�J�>i����0�!��ۥ�n)9F�.*u;-ߛy�h��6M�I��� �	�F)��锥d��`��d%`���ot�ٱpn��n��,���J�1�Ԃ��Ri]T<�
	�Wƃ���U�T-��rW�{�)�='�6�r_z��b��?T�,�ʘ�T�a���)��u��X� $u��7tQ��r9��:�3��Χ�ad9%��a��]2/�,X�^ZHk+��u�Y�ac�I�q��e�劆5W���Fi���2«0�U�N8)�9(C�U�xM�#�s4=�|�t������uS3��_��%�r*0Ee��O�lv����5�
w=�f��kq��E�9Cx\8�\Oh�G}����V���:I�'nGEъ�J�j;�
�^�ĝ�б],<�Pq�#W`�ۺcc1���KI;F��]4�3+l�tQl�z�㳰j��O�Z����g��F�<��w�L���֖z��k��^c�NՋ2d�}Oj>�&����X+8(�� ����m�Ej��M
��������&����y�,)�20g^�a�9�Py�FP�^�����.,��t/Z�o� �@jWW�n�_O=�u���|^�� W���m�x8��m:\�zU���S��wd����y�����8:�"2����4�t�,p�C��6�P�2n��n9��S�k&�^��\f�9�:Pw�N�fy�f.��V��1ݐ�24[��{;��tO��}/*��;��j��|(p!V��_�E ���i��yS1���[=��\�UD��#:o�oEW�Td��WJ��C���,Ļi�ې�	�1r��>��glwv#K�51�>݁��>�_�Á:M3�$���u �aA]��z`𤗄*�%OY�_�7w��^�����Pd_���1r�),�z,2��v^
�؆P§:��=,���۽�S�9���y2��o��"��C�L��ɥ��N��)�|��՝L��k%���&��d�}\#��+'���:�88d<w|s�-��%�K]rLwM�����ta�+ioQw����+j�&�e�x����k�-�`}3����*�]C뤻�0�Jk��ޕ��Y��R�^����:��G-��kt�Ĳ�\F�q{�gOX�Pu�Eg-���鏺�u'v�C�(_ ᝱�u�QM�!_o�n'qܟ�菫�/���;��K��^'��G���6딘6��:.�zE�e��w` �R��:��⷏jk !�eN�1R�Q�&I���JZ�wK�}Y�5v�{�Y�GU�v�1M���;�І:ۻ2'pp����X�w2WJ���O�=(�������ZTJ���=o�j��Oe�J)�f��Xg%�u(!�9f�f	e_*x�z�>�r��{=7mԎI�'$��8XW���my-��`N�e�yS���@f�S������'Չ���/��y�8gC���w��'`0���s�V��X��᜖-D��+<jVx/1�j7�b��T���8�C��ӁsB��&�F;�̞s�SX�K�ՉV��OP�ؗG����Z�"�Xb�
���	B���ݽ>Z�
�Ø^�����Wa.p�Cz����|��m���V}�[i��P�V2
�y&�u�E9�����=�G �d�嚵ݻ�PcVD<�=��l^]Rgn�ASuU��@=,��ʐ��+������{+#���PVVGz��fa�6��5㓫���MfN+wd��y�i�
�����M[�q����wZ�.rW[�+����ـ��2��ft��ݶ�pT��D|*#x �G�8E��q����/K�3��s�UW�n�\���y5㼆��S�gܜP�b7C�'!���)���c��=Vn�y����o�u�@_��* j<����Ntv�xG���VD6�K���e��T)�LmZy��R�i�t��ڦX���C0�o��W����xE���"���Eu���;<���yN��Jyv
6^_Zg>���Ըu�xx�|�,d<e��[(\�T��*&��/��i�\d,	T�<��zb��yƃ���uru�U�t���{Kэy�̎��y�ܡ�zz�NO�J~z���$�K�3���w�W-�:YݙV`�o<�0�P���.)�,�+�\6Ɯ�7F֌X���P�i+�#�Qyh��.�8l�.�ڲ/vA2�d�ҍ�W{I(y�^��8�4J^Reؚ_�%�Qi�e_��]X���y�������hݖ���I�A� �qH a�����7�3�e.��Uݴ�G����G=)�=X�Z�]�+��r���P�V7���v��{	�{����ɞ(�L��>�[�e�/���v�nq���@�n�)�\�9�su:��sp픣���[��w�j�ãv��`�s)���<�N����f��K�dɹ�2J>9�f�R�'PK-o�u7�a�1�| sY1,��zr#c�����[��&�V�#�����fX�yF����a��L`��>@|o�[Hj�ٸ%U$�՜���e��ٍ�7/�&'��&x�;>��Y�]Mk���·-A�V�����VV���H9��c�r����,ea�-z%c!���0�܅ܓ�� %�*�V�J{�b�@�`�J�.��{9��r�q�<;!^^���C~�tx{%�%�`C�yn}=�t�����'�d@���ԛBqS�;�
��y�^R�U��)+)��� ,G|�H.�]���ޙ���:�ǖ��a�ym�P�tF�29-(�g���U�9v�mu$|`R�6�%�#��L)U�:1Jr\��r�/���\4�*.=9�1����y����hd��E�نɰ�&���A.��Aߩ�ɸꤥl��`in��{+K޼�Mcn���ix/�n,���͙hRd��r��zs�Y�W0n��!,}�;���He���;Wac�Y�+oʘ�����)���������<���'/qT�ۈGCM%�u(>�X�+	�����P��Kb7���ڳ�9�ug%�A�
����;�뺍�J�2��W��wټ�M�wj�j�����\�&<7S���I�goK�q����4���ڏS�2����\St�Mk��U�zc׵��b��p�Ewx(e�>�P�Rŉ����������'�{�y�[��}~��=�W�;Fc�0�U�K�=E�1��"�u{�q&�&by��j�P\lWd��Ӧ��>������}��	w��(J�:��R�%�s��멜�k��㌌��`�a�:�6Ӭq<Z:֓����� ӝ[A�e�0��(t�#V��[��5d�a�;̋���O�=Bu@������6�ˁ����[��{�+��^~����<��^
�
ߢ�l�U�(D��R���7u�iS4]�:w;��!­	H�������&,z9����Pޯ7մ����^C�5�p�׹Wy6�/Dn��=�4�ەf���o�J⓻���-��z�][)��y��eA�Z�f
ܽI"��fFR'C��A�ղ�9�i��V�e�)��c!S1��������Fdu�eEP�.���6�}�[��Y�3L�[Jh�C����i��}ޤ�Omx�T%�--42��&�������Q��ZN�u1.V���go$ �v�Q�E�]D�k�C�r\3s��:$�t[���l��v�DZ�땾��I�K~TtsK�F��Tu�W���H���9���K�/m�mf�]f��η�Պ��hO҉wP���`�&]���&"]���e|�7�Sa}��y�}/��-&���E�%�ҚB��%��5�>�3�m��s��xҞ~��&���p5� ��f����\�)H�`�z,2�;�팪'(:�̶�Ю���b��ʥ�N�|�A�v{�nN��d�!c&`g&�a:��u��1h��]��+}��E!n:�e�]1:]+��"x;�S���N��e\�`C�fRC�9��7[6o/����Y�T�5���u5V;�����3Oy����j5*=V#�4��?�sdt�I�XIҗb��ׂ�>V=����R�wK��ȇ3��t+ƅ�щ��������W����.�z�!���G�y��uUs ~Z�_}�0$�	���z&R��y�<!M�����d���3.����yNDA뜳H3w��f5��^�t�k��7�9�^\u�$��,+X`��V5�߹>��]h���@^��|yj6�{=K��a2�~�o��4;Hg�x�v�E� �vV��5[�p�+�~ա_�z���Ƴ�U��" >s��gPٶU�Q~��^��y&32�S��G��ԏ.���m��}�rv#�� �)��LX#���|��;c�vX��	R����7������f+�l�����E	�/�:N�2'�vrJ�#ϺSLZo����K�qӁsB��W"�ݜ��Z8��Ech�e-��YW�q�M�1����B�C�Xr:�J��� ���+Z;���x'+d�����I��i���l��Ԗ����ݞyZ;���lnz�L��cR�����ME�;��|�O1�[���+o@]K%��jǖǶ��i(�}I`|gԒ����OW�+5I^;F���t���}c�=����`.[��8�:ע�K]�:��QP]詮	��O�j3�R2Ϊ���,�ó�izhO'��n���C�]�^�=VTD$Ĵ�
��eoz��{Ϟf���C0]KL�J~X�\#�q��;\+|�Fo��dƼ2;�
2�w{�1����#uՈd0i)� ��Ş2��WS�R�NkG���c"{|��\_³}��#��b��}��A�{a��Ȁ>�(�x�M
��y�jE�Z�����?j7�mm,�Xw[�辜�����^�� ���GIip�E�¸d�U��������$�<ƆC�˙��w2p���[9>�>꼼�8�Pu6��vehn�7u�cU]����h%��z��w�St0jC&ol����l�ݡ�^h����}����=n �Y�r7��iU�z�����*�>����7���8F�֩�rWG5����<"�pIF֌��傦�|}%��Dm�㢖%�{,s���匴3{!�������,[Vg۲�C���Wl#���R�$�`���P�.B�q�~���'ܲK/۲�*�j9��>2��V�焫	��6�I�����Rsg]�`S�N��^�]=51�)m���ļ+^*|g�m�M^j�2��Ј=a$	R=3� D�%����Ev<t��g�����kjcu�U�g�Z����,)Ș���o�X9�m�q�&H��[듲���=���)��Z���a/���1/P�8+�}�ٛ�
��s3Rמ���;0{�OOs��9׏F��V0<5��D�d1uh��e���X�Od�N��Y;���"׋$�Zz\��r�|aps��..(�����������oj\���2�S��W��G zjD�m�-9� jOPs�Mu���y�%1� ֶ%i�[*��]��&��<�r(s����:i[�P��ӱs�4�?�=o�<�o�Xd~˳�a{�h�M��'r������j�)���(�OID�e�:]���\�]�B2��Pdzp^��^�yi��*�2y�Z�[��"�����=�8(�&��sM�6��[�Z��i�ؠ����e�"#�f�"��j�n���ʉ���c�+ �6�)*�y���1r�]�1k('��^j� ��rQ�;��!yܬ��y�Q�y���tA��(��Y�r*�/MLB����aMʾ�Wԓ��j��M̴�$�v���b��d�-�VJ�F��:_T��][6�j�C{�p엵k��zX2Q�S�;����[7/�q�F�� ��¢���)�u%�j�0ݲ��uiZkk��;�!:�T�E��v�oj���*Æ�0�Lα��3��:��,�]!��d.�\Rܷۡ����yَ� X:���ӊ�G�*V��-,���V�V��W4�h�lfAEc\�Q�å�'�:r��7��S��rk�fv����+��}͛��d˛W��ٖww!��Y�XB�C����;Z���uj���*X��١|�Y��=�nъ]�-��v���Ħ�k* >X�=ZՊ�[e�FEih�sU��oSi^�}]v �M��Pe�.�����w[M�j��ج1�F�����.U�X�	���-̼6�t�m�9H����[�)rl����W����Y��Lq4��:`0�4�_t�,d�Z�{�n��SB!5w#֮�35,�μ��3��ڙ�'=n	[������ՙ��υqwH�uӮj��1�܂Q52i�V�Ci�YD�5Œm���6�Qj*��L���[b�y%�ż�h�c,B��.�����ܕq�4֥��f+Ok�w],{L���N�BZ�z���Q�����;���
7�R���o��J����EhH�w�aoL��Sm��s�X)��b��qv�MYOp�d�R׍w
v���ԕuq<r[��d�!Un�J@�x�#�4w;x;�ɝ*,��v �/+vr�U|yfrs8Gd�FB�4x�`�e�0gn]ڠ.p�/�U���e12���#��4U�	*5����^��/�ӝ�2�]Í�,��R�o�e�>{���W�e�S4�F��0>�gF�B��x\�k]�k�Tm/�4R���䄚ɺ]���PD$;�J�������M���]!��3��f!���)������{Z:�;�%/8��u��m݃��:���۴��C�, �Xk�f�B�!r{���Z���f�o(�/�^a���F(�1�ג�3w(�G�Vh�,��?�nY��}���R�loK8ݤ;N���}�,�3�)�V���BIe�u�9k�:z���p�m� \w4�QNkm���7i[����O][��ᕥ�P���H�¸c�������:Qݵ���Jn}�.h�<kõ릋���K�ɿb��`���:���7b�s,oe�� mcֺ�}�������v\~2�Ub��E*,Pb�BX�UE�,b�DdF"�b
�+1Ab,UQU����V�b(�����)DAT�#Q�mcTH�Ȩ����`�#Q(֪�EDDDT�QDQm��U�TTb֌\R�
�Ŋ+��%h��TX�EQUUF҃(*����p�Tp�hQAb*"��b"�X��R#1j�TŨ��*(���Pb�Ub���VA��Ec�TA�0L"1QX�b�H��a
ň����1UADA��b�EEEE���U0TD`V�V
�Q�aETH��`�Q�>���1e�u[1�ܹ�YWIV��v�]�݆خ䊮���,��\#��µ.����_J�:�躸�u|�3(�$��H_K3!<+��L��&&:���R��}r/9Y��<�*�z��L�y³�����؋;,�.%ȿ�g����$��}��6��l*2�>�=��~�B�O>;g�B2�\�����6e�o�)4��y�"���z�H+o:U�AO�9ػ�U����O�{���LB�E-mL	=���E�u+��%��9[7�y��w:kkVH�PQ�3���{Ո��᪇x���P�(P��$�p#laJ�5L��w>!lˎ�/ı�*�P�d��F3�Ԑ��4T�i�.�~�Vk�Jͳ��=F''�5��w-HW@d���Z>ӎ7���s��b����K��{�:��"Dx���s�o5�'%Kx	0Z�o._�Y�m`��kh���z)�e 3=�n減	|�D�����YJK�}hk:�<GM��edY~�������FPؽ%��j+MN�j�es���9�\�y֑zر�����^�����{�k�F�[N�+��o��X�t�\ޅئe�����j��`��.���8�8pl�-�	���'c|{2A�����XG��I��,�륄�sn�]N=�A:��A|:�kֳ�x���r�gB:�9]��.WR�$��r�\}W4�ܮ;�݉�Eg��&J �9��d�E�⃿SY��=�Vwd{Σ(9�c�1n�/kǪ�ǃ�YY6mpu���ǭ�r�K��2j	���nm'3~:PwI݌�h��3��꘡������W{-�o3[g��vS��q�tuV���QY����L���8S��:�<mj�`�u�G�D���'?BZA��o����R�#�:�[J"�����J��Ri���"�,�q����쒮�a��7�XD�*/l��fc,�%��8t�6L�I	~{�u �`\yu�5��cB�J󞎽��G)Esϲ�|\\���#�0��y��)�g�ߨ&c�n,~&����K��֖Y��*����W���<�y2��o������zf o�K�~��voi����p�QL3t�Y���������r��t_z�W,��q��f�Q�统*+�v���
g�eD��KWl���:���T���+d7��V�%gj�5J�6P�Y %i�
_o#���:��.�.%-]҂:VD8򫱕�Լ3k5�y�֎��ұ{����
��-�+sIV�`A��sjQ�Ĭ��)J�5������u�+�sg$��������&N�'Q�ݕ՝ebcNwø̢���:PY��e.�d�C��.�z�խk�ܩ1�NA���6r�(���*(caa	�Ƨ0���͹Y�f�S3>	��7�dv$Y�u��3Qf�=��"�z�/�R�ŢTq�M����ҡ
��0q�-p�%���Ƽ!�fϯ��@�p�n5�ֶs{{N��(�in{Bݹ��K5'��k��\�kR�-Sr�������E�'��X1l��LX�x���K5,����#E��C#v��q�>�v�FE��[ҽo,�೹�9��t�F�գ�\~��0;��*[�ྺX�͢YӁ\�0^&�E�ݓ�)3T�p��4�����^�h~�Γ
��1U�S1�l�z�@�������Z�{Ճ��F��o3	��9�gխ#r!���9�O�u���Ze�S%��*OUu����|��w�3N���,�.�]���V�y�jǖǶ�Į�Y�I`|e$�z?0����z	����1.���]�$�H�TiEb)�L��oW��L�^ Ȅ�vV�sٷޒ�2�u�S���g)88��U�R$l������v�x^J��+�����!�嗷�Y+��3u�;�#D�����:�".[�8�s�l�UX�诡���o<��!�s��݌�x�c%��+��R����7��q�s��uw��:�(��gw=5�[�읕��kt��.�U4"޽�p��-��_f�i�w��&�x�ó�V��s<"��3�����C16�p�����2�ESy��c{3����U�$�V�O���1"el����G�x�]O&�S,j�G��{Ӓ7I��Gk`���K�O#��l���'�D�!��Pq_�/+��l���ջ0iW�,�Q����>�B����.�y,T:f�t��$��_3��l7��7��p�u�g*8h��q�X��܊���fM�SÊe���#�YR���������6[|�hc�4#Nv�^�32G)aX�탎Q#A����c�=� yI(v7��ۋ����&o��XH��1Z�w�Td��03'u�}��	2�RN) {��y��G$�;������#^��ˊT�nA,E�*o���cD���H1����"U���`�����M��䌊]�%1+l[����d��OƲ�7\�SV��܉���d��������@��)L�Ņ�cGθH9xh;�!x��.K�^c~�\�z��M���(XZ�I��E,;Qj�[���`᮲�L����h|"��w�j���x3�%p̙Yo�/GڒukVX�$��"Q@�1��ֹ�c]��+��u�r�	fm=!��bu�p58���S������� Ѹɜ������� �wlX�7���׮+�A����HWW�s���;���=|�v��V;sحޱLnxoC��b�%���i�kO�}#��q3r�#��,�u��0
�xr�����Kx��W���!���!
��W^��|�{���>��h_S�zjD�m�-9� jOPbq���"�|���nE�Uu�.�jCC���R�*��L�Z)����2�Ɔ|P�`�#k�G�v˞>�i�Z�[�W���
ZFq��\C���������fo������8f1��v����K}u	�bqH+�yr��v:M)�6�Y��K�&Ϧsu�>yꩄj6�h���o.ӹ+���9Y�x.`�X�pl�@۔�V*��P�3׶��n���Mao��٩t���f�k�㸟J�/OT�,�S
�,92�:�"�������K˭׽6Ό/��Y0�]3�B:�,,�$�����p]1Y�s4@fԉ۸+���~t�Bn����UC��53y04��b2«+�*@�N)t��׃�P�t�mX�ٽSh<y�5�N�u�LV����7w��<�I��0���������т���e�!�7��EJF#43�ZOp_m>�a]l��bʸu�2�eu� �)���ʐ�������i+�+4s7#�k��Wh���Q˗M�ub�6�ZH��@l��[d�iƗ������(}�s�"Hg�c�<���7ݞӀ��TԳ�v�ܬ6a���%��^��*�ִ���z(�on���7�ۣݯ�j���s�6x�A#��b�:�!�@���qpn���;<�%L{Rs�T7=]�GU����(f9|���!1x��vY�����!Enz3�1&�h����q������V��\8�D�ˌE�1oS�Ӱ�����R��kg����z���:tA>�#&�NM��^m'3[H9L�n0�bޢ�V�Ӛ�N��]��^m���[����W��)m�aJ��/�e�{Je���.�����;�F�{g&��]�4^�k���w�!��)�U��(q���Ř��ԚhU�-�B�r��Ko}��G� �u���l��L�<\��>N�F�g�Iq���u@�3̹~�s�̻�Pr'�ϩE<������f�A�c���瘹b���(s��p���L�]P1ޮ��˰P7���7�*qOoM�� ł���{��w��\F���ɜ�
.CY�R�B;*D�qN;w;�}kS�à�V����]���0�c�+�s-���37�yV2�v���j�Εv�t
1���|r�}.n�)��������ͭ2�J�ޯysBZ�����+Zf��8�MW���K�ς����+����R�Uu�磉A�C�S���N��e\�qߵ��ʘ�u��9� ��T�����8��̰o�vO����pr���,����2ge�)�q���t�Ña$tK��5u���M3�-[R{h^�K�8��5~�=�
X��o�Vw���� Tta����'�h�f���Hp��q���Ozn�;GɅ3����:<	+�!\��Qk�	-6˨q?Z�D�4Y�K��λ���d=��]��M����S9��%k(7C�毗��:�=���d'�!՛@l�XV�o��� �pb�aC��]��b|D��Ǟo��?  �;+D�5[�c�2��:��v��O�m-�Pl���^�aJlj���R�{U:��^�Y��8����H{��L�n��25JS�\BX�8ggw�q�`,r���"����
�ql������}X#�L]Q!-+�^ߍ)�ƺ��;�1_S�ua�Ww)P��C���B&�I?;3I�Ω�Qׂ��$���Km�+ ��kX�؝:яy]�C�=iQ������eG]nޤ��ʘ����A뼹-,��׏��\xR,��*�cgUk�Ӝt�
�����+ݾ�k���m�<�Y�`�mf=5��	sԩ鮡N�m�p���x�¯@���ӷ�&�_���I���oW�Lî��<>�\��;IF���ʤ��V���m����Z��fp�� cr�skiEqNB)�M+��?��K]�:�������;s]	u�s���ᮦ�u*�ڨ�6���.ߧx^J��[���UrzD�^Z,����q�+ğ%����x)W�N�8J~XK�3"�;"�^S��罷y|K�ow��;/�0�W��`y��镳0P�����+��Ԩ}�V�5��zu�� ^�y�8�7yͥ�a��/&���9�LD�O&�:D�3�c�(8�X�tf�1���MC�`:�:I�w�<�ռ�+�rj�wjKR����bŁSÀ�))rW�S#�X!���4�.��)�W�f���S�X��3eyߦpIF։(M\*`�p)%���K��-�M_yќ�pr��y�f�PUqw��/*-�9�-$:(_C�TN���[��-��=�W|�* ذaK�v�&|ld�S.��u�"Ʃ��Z{E���	����!���j�.��`�$��M]��s�ٍV��c�cmc�=�%��=`^16e�v�Q�W0mu�^�a)/��;p�v�K�w���ݬ}I.�;1gj��I��	�q���Ϲv�V��gd��n��5_��e-ݖ����a3&Â�%����Ľf��ھj{�s}���� ��·��J���E^ж��)��#i��X�E�V�.�B��;��46�׷5�����SspY�;��#�֗�i��+��GSQ�X��Wc�g�WLݑ��Mi�p�䧧���B��-;����/'��O/YGϳr�"^�y�᭪�j�ת�mN#���T>��Ӱ�O�:����ɨ���)���nu�C��!������N����^V� 5��_���Y2�s�aq=^��ǽ��f����\aD�����ѱ�{���t�ܦ�q"�T�?S"�`��=BiO�H�������Z��yL�{�|��=���Ƈ��:�1SQ��p8Z�2V�a�C�����CsI:���q+H����C��ޤz-#�ƸK�v�Ջ�c��������#X��h���f^,����תȿ+�����W�.B�v,�r�F�L�C����u������{D�@�֌甙��x������ten$�v�ۙ�J�콭=˭VJ�5�̓U��X����L��t��ŵ�������Ƙ{:�jx	������{�lZ�֬�x��O6D��N�϶}$3e���fMw�&�J�^4�v`����={�8�2�u,m���;.�:�&��C�C���č�����-n��Gp�B���^�k�������15���<�W%�s{\���o"	��-��;f���e@�k�pl���!,,rK�2���B/��V�{�̽�u
u�HA��%�.���՚��j�و�jHas�*@W���y�m[���+�v���с�gn���O	�3�vI�J��pJa�cc'��q3c[r���V��J�`O[�<��[��V��}U�dc�	�C^z��t��V��͹�p[Lnv6I/N��εy���g�[��2�agTv��Vz�!:�!�=15�S�޷յ��{nZ���f^��K#kL���Asմ�.����`K��ݷ�X�w*w��h���O^DS��Enz�+���^�r2t7!8�H���E�0�3ڜ�w/9磼�k�ޅL*�q�N�}��4RϏ
��o�.jc�J���&z��'v3!�f��mMc$q���zנ�S�l�'>�7��՝4��@�������0�$�2؇�*S� +�2S��gv��}n�Q�K�c�"�:^�+y�
ne%�}ϱ>�����`Ӓ�"t����Wk���9�'OX�nc�f�����Ţ�H��ZQ�Q��ۚ�(fh���xn�T�A�LHȻ�X%�s�d��/����4�%��Mv��ý��מ����{
�����)(G�i����x�f>t-�( _��E �S�N��E.�݊_.����:� ��&��I��ܼ5���b��<�ŵoGd��e^ԲX�oB@�6M�ۏ6�p�����y�r0w��n�TcT���}Y�-�]�!�9�x�]L����B����3�/&[TU�����@�x�\t5,n�3͘8��T�ۘ�6�?MS��`=[%
��s�.We�v�v�n�r��9C������~��׊g����C���F�	2ô{*�ҋ\�m�����t&�#�c�GN��L�(����&9豸�	�*i�u��F�b�I,1X��B�l$�j�8l�1��l�awN#D8zeU��tek�5V�1�{I�{�LdWw�/���U�<�'Q��F��`J]��M}��/@���̬��W}�8gAwN7,D�Օ��c�"�>({���Ùz�c	ê��6VWv��\*��ag*8�4�?e�`�p% A��^�gv
���+��sF5���௮���)ܘ�\{`�cY�����c'V��\L�h\�|�QgF�fGv�$���2@���s��1ծ�]Z�M��ù�,]��������m�+�e&w�H���{-�n��L�h��ܭ����J/�.}��W]�*���±zNq @�ڀص+WG�u��:�y����2p�{V�-��#y�V��z��)}�m7�dd��@m�����R[����@��'ž��^���9$�1��A-)�u��u�%=�����|�]��AY�[m�%�œ�fn�i[�ͥ�j��5;B�R�~�m!ܾ6�Y��I�xv��m2��qr�'���8K��;�%��U�[��n����|cnY�io[`T��7!��@����iƅm=�Yj<�w!�]�X��gS��c��6t?�ʅ�+w+��{����=5���3����Ը�L1�Ep�%	SBH�C�T��ꚝ��}7�ε��r��v��BxzKU9�k ������D���o�f�}+c�5��3��a�}�Z`?_I�� �]�6&t3z ��dvs��]g���S��V��	�7�/2��/����G�Qȍ^��*d��Ώ{�O�WM�@��*��xVn�;5��M��:����t����W5ʐñ�4��6�#܆ʡyv�Zkq�����,���:�ᢹ���ٹ�[`<��|/SR��#;Uk�DPd�G:xփ�W�a��]h�G�?�x\s��* �(�ykb��QUH��EFҪ*�F ���#lVڕ�U�Fڪ�1�Xւ�U��4�X���0�������p�,X("(�j�R�ZQU�1c��%F""(�X���-�QUU�ֈ�e"��R%j*��UVPTU��Q�ZETih���L*UkPj��V�L8�e�m�(�"�ֈ�ō��mA�J��E#�ڌTU�X��U�D6�-�1��,E���X��*(ԭj��TAH�,V
+m�QE��D�Q-�m�[J,"����Ub"Ɣ��PX5���+JYF[�Pb�T`�"&-chР�"+iKeEjX�UKj*6�[J�b"(��b�4@(
^ڊ�-�9-���{/�Yf�^.�:��Ե�>#��͝-_+�;t�nB�xqҬ�Wj���g;��(v�s����urs�)��Y�|&{�N|&r���[h�/}A�l�iL��ifU$�^��U�3��\��lvu��#.�[=���Hb�(R�}>EV�.�Z�<<J����r^z����9�o�������G���	��s\W��^bg��X�U*A�9��d�Z����{�R=~|��67���qPr���Ԣ���d8����A�c�Y/�:G�H��}�L�z��b�rl�z{3QzP�C��=\"e��~�/���h�;[!��{X��e��y�u�H��`��W�P�e��2�xE��R+'�<��88c�w��dW�N�F�7!��\9���� "��䮓��B��Q(s�գ�_�ޅWz8ͪ�l�ta��n�K%kQ��}L�Y��#�ZWR�����;ν���&��VR�1M�3T��ަ�Ҳ!<�|�g�|��n�e�2%`2B:�B�i�;Ɣ���ݷ������)z�1�M7�@���L�(�����3.���k�r$Y�;/Ǐ
�0U�|����ΦM������=��T˭�V2��� ���C{4�V�u��DD�HL����T�Y�Yx�mk�ۢ8�.��/iN�D}��#a�M.�r��d��sRWA�7M����S7:���ۘZ�����9��{��[oB�]iw���������i-pPZ$��q[6N{����m��fOd7Qm�h�q59��X�л,xL����_j�֛���w��&1 ����Vͣ���Z���i��,bC6�K��A1~-2��V��e^&:�<v:�b�������ߣOo9��'�_��i��v;��u�֍�Uz5>^u��p������W�6��v�R��l��Yi����+g�#C��vs��zh�ڭ2�*�ٓn*�ѹ��V�[���|�dtΥ˛�|��Rwld�+g<�5g�x}���,N�YȖ�J튯=�q�+N���ZP�(� d�hOy�(��!0-���L�^D$�'��6�m���l�[j}R�������x*�H��A�=H�~��y��9��~��c��y����g��l(�.�����Q.��S*����g>�O�!S,Fc�!��������N�ۥ�Z�ю�����i~�a��u#�������=S(P�ԙ߫�y`u.x��Oh���k�3�!�wDҾ'+\%�q>0������|��I��]���t;����>/Lɤ@٠�+��5� myXr�{'Y{m�c+O�}LsʹMuf�ȑHv�Ӎ�|��c���[PU:8�����ti�]t�Q�lB�wc���Y\ܜ�u��|����<��%��򘉇��"O���A�yƃ�"����U�G���Z���~txB�sPrm�W=e�S�,_��"瀀,κ�/�v�ԯH�8uH&�c�G �6�E�<we:�a��ӒQ��$�9g¦��I{0�95�F���!kӦ�mVLwY��sFߋ�����Vz(^��."G���NM��;V�}Yz�O����O��N��Q�'�D̪o�/�w
���g�o<%Zf4N'�����
���k��v��`Y�NZkMTZ�X����]��J�*|tD}�j��N�U�Q�t�ӍSy���`��x��=K>�Х�{&Jbm�uҵ��~���4�7\!��${]rv{j�t�����׾(�tߺT12�o;��:�!�r���^)).I�|�r*E�37[�^�z����1 �X�WL��`o�u�!X��6���1����TE�%>��h�;��ǳ���kfw����� 1Y\�r7 &^�����"�c�p+Vg�l3C5��/m<��+���)�3h�z!�w{����'ق07Yb�X���կ/����]!����M�;څ�4��b����&[�:r�/�T�K�9����*�8�q5l/U��'�]��y;Y�y�wh�wwS��s��}W,s��]6�m�m�Y��W�9I�S�+�_S��H�ni��<]I�;����gʲ|�Y>s���g�
��x�8Q�q��du't�l����tҿ��P��͢K�W}I��;ٻ���G�|�<�`S�O��,�Hë�p6\C$�k�\ݨk;`�V�S�%�lw�:'�s�S�s��C9:�oecqH.vd!���6�Ѱ
g�qgf����_P��㜛���e���V��zg���;��b'��eB2�\���7�p�ٖ����h�=Y��<vd��/'�\ QdK�A�Cg���������J�/OT�,�ST�aڠ�d�lS�*^���� `ݤy++���{%��\���fur8XYIc���3�5l��V*uj����D
�X>�Ier[R���K}W��U���v��t�����C�-g���ԧ+n@~�qO�\*�4�$C*D��T��6J����N&9E�1�zt���.{���"e�]�Tq�,�ORϣ�v����8��'�Z<6�]3���Kr���luv�f��51�GVc�"�*�|�1���P��v�&���ײ�j�!w:
��W'�^��q"�Ǉy�x����bgh��|�:{J*��k�rQ��)����C(ڊ�_=��V�c�j'eo��^G�Ro3z;Js�z�T�r�CvP�Z7���9�ac��B0:���BP�����ߥXB�;4T�X�Z�Î�7\�<mi� ��ֹ��Ew� i{�}W��z)dBn��;=��Xz�$y�]�"v��D�_5Ձa�M)8�����$G��;��5��X7E��h��w�߷��P����豢�e7���2S�GJS$]Nʼ�I����w�觨�����-ul<�;��F��}&�s�;hZt9 �[.���h�Zo�邺ZO.CI��K ���zt?*f0\=�z�g�����f��[je*E�;�>�R�[u�)m��J���M5��� B}L\Jg�港gk�A�,\�� �C��ɟ5j�!�E2En£ϻ��3��#Rl�}�8��N��>�8{�p~�]u��2�� �����̌����so: )�k(.2�;��U�/�H����83眲���U�:��ִr�y�[��G}D��k�@���t	U�]E Ϯ��1u�0�Ed��x7=�޺g6�
�<�)>!�qN�YOd�v�y�c�W�݈��˥�s)V�Tv
*��y��L��'���ή��ˬYlH�rh�5m�ym u5ڑ K�@	c��%-��g&��n��e�yKk:rWi��Խ���(�<�5���%b��Ug�v�b��<�91�b��%�X ��r^��r	�Q���01'��,�C���g�x����~N�p��������T�'�� ��:�>î|�v�W�pQ�N�Q��:�����N9�R�/~�2!��=NGAe�J��a����6Yr}R��U�ʰҗX��jp���`C<� �j���v`IXn�
��`��[�vi���r\Ur\Un��#�$���z�7��!��_mʿ*y����i+�\�,0\Vג�-M�]ˀ�7���-���3;o�`A��i�S�A
�fP̚�
t`gy�q ����?jv��F�������kܺSȌ>�o>U��|X�G�3���V<7�-ڞ�5~��7��uF$����y�:q�܌wQ�;δu��#�{��Ö��ʰ�G\)S������ݣװd�浑U*pm��W80'+f�>�j�u[a}<�\�3m �zfz���lU�y�<T�>ֳ#!�n��ܙ�sЏ����<���r�������#b�]v��k=5�����H��r:j͝��$��n�b��ޔ�0>$em
C8/c��ޣ�r7]�,�}k(%;V�$��&^���N\
�͚�Pcz�QPwT��L�h�6mݎ6�&�@oB�o�e��%���ğ��o"32���,J����O�6�.숩ӓ�?DUR� W�S �		[2��r��{�ƙք�K�����Ŋ���y4��.e̬�����Œ����҃���o����J��]eΗ�C Ý�F�r�o!���O�ɇn��o�\	=�"��.��TO����|d8O��9�����Ǧ^��mR?�9�i��]���G�fbYdp4z�s��L���y�5Cw[����;���٧'
��fX�x�ɼ�P�
b&�zx�<�$��w�A�׬_f��2�=)
ǘ��	�t���e�{*��
�������8T�P��aH�:�������hZt��8JOy�،�b8+B����ѡ�Y�q�&*��(��%	�K�O�bz�$w�Н��r�@��G��]f�fu͠���ʋk}��%`�S\�FՑ9�l�>�D���=��C�ݧL�'F��O��
U�.��uBǙfy�^o@��Y~���x�Nx�Y���B���H���q�g&���$Ҧ}�p��-��j/��E�&`ik�iߡ��'�����!`o�;����V
�Ԩ_:�@�I�|����H����T�;��],�*�Ǚ�v�s�N;Ra=9ꮕ�X�oP�?:�N�]����Y���A���۸�)w���e��Ö��7eu�8�2�͸���f*�~�{�E�����dCӦ�����fщ�3Es�ČL��;�C�)�jN{5m;v�:Ô`�R��&T��<(w:�5Ή�xh;��i�tz�B�=�
��7�{�W�z�R�zJ�~���r��s���*aL�[E���,�ò`�gQ5�r�Ӿr7��W%�mAN���dо���	=�z��ʇi�n/|aq=\Gl���ڲ�yj�;{�.`�z\�(V�VZ1���B��_S���P�	��2�ۣ����Y�vd���ʴ�;wP��S�X�w{ɡ�q��`���Cg��<lt�O��a��7���lV���Vo'���:`	��}�T�^���/��6��%�;H�j�P���|��`(z�v큉�z����\jB/����r�ǳ�~�x�D�G����emL��:h�S�Wgr���N�Nn:�)[:;��9Y7�m��,��v��ԬDη&9�{��/%*�ֲ��/����Uޭw\w>O�{���LB��1M���Mь���g�u�
�+ 7W�sBs����$�f����e���~Ɗ70��>"8Q��2zX�p���0�V8��*�/�|5g
@scbz��d]Ew�hv�i���r"��r�c�.�t7�a�[��,8�n�9E���v�٦QW13����~�����P��7�@��R-#N�#~%�ɀ�e�J��LU#��!�a\T���k3�}Y�L-�4ʥZ�o2M:�Ik��8߆�S	�M�FC�3�`f���t{�T����gҩ�`lS�b�J�!i�6&p��E�۪f=�pފ.��{쥾\�n�^Dtg`K��Tx��l9K���dc��	�y֡��<6�A�7h����޽ַ���n�NF��7e%�b�~s 9�XY���=�B�,E��.���v=ȭO;�X��aZS��^g������Ӟ���x���0%�|5oj��aj���m�<*�K��ǥ\|���k�D��Ǥ4H��E�0d�����j�`ΓH��ޣgT�<��z�n�mK< �L�+��uY`��Ӊ`��`E[x�%n�㹩YW�3f.1��V��_{��ӂg+�^�����r�A�հ�3�D�|���g��}��S(`���g���7��ힸ_zg��8f�dK�EV�'7j���Lw�|��x
ui��o5[V��¦�9]̤�%�}4�{�)9nr��͎��i�Y��˙�h��ű^0u�"���/=�i��!?-7loڱ��FT1mCLM��F���Vv��&�Gո���Y�崸���;m�}����b�ү�Ԛ��E�Ψs�����/�fz�(��G���d+�l�,�w�,�%��HV���Azk���:�V'�e������(2,L67��y�V��rH�SZ�]H�eq貂f^;��U�/�ۛ[�'�ྙ}η˥k))��;Jgn�x,O#��1|�\	k����қ�W�}Nߗ*�z��0��e+���R�Jp �������Y%�KЮKԞ��B��*%��Z���Եaߩ��7��}�2�ڶI��Ц���,�e�6�� ��#��}�\n�NC���n��{vz�p���Ѱ�>�&!s1 �u\C��|�
��Pö*fa��4���B#
��<�m<�ܺ���s�����Z���f����+3�ف%7P�rf0p9E�$�t�3.�o���!}���%�7=׫3�j�UC��q�:�3��kmC�)%�$����kR��;��D�,ɘ�.p��y�v�SX�4lK��!
9N�F�7��dX��,O��ɺʌ�t^P>�U��ݵϕXQ%Mv�ԛ�`�G���4h��;���V�mn<<j�O���,Rn��V�Ϝ��;D��s{G!��F*��Q�
���E3�Z��AT���&k�g2��f>��:�e˰ X=�Gn�M����m����ܺ6�#�y��0d6��QW/X �/���{�9R5G�{s,{��iP��l�����!xe�yS���k�o���ܳv�BF,�;���n�e�x��VI�r���u{WR����;%S�_1A���L�c�_t�ۡ�.�B�7d� @�'Ec�
33$JY��Oo��Z=��2��
,�ϛ7Y�Z�ArԶj��xoK��R���vRv��;6G�"'AI�0�e��Tq�T��q����gI����*Y�b��]��j����V�� �bo�f��'��yQψ��W��nU������K�\6���w�Ю��_b��yY�u(�ev�>�nYTt�Ysc��_b�t�u��Kۛ�f$"��[�����{�>�_ƨ�3�W1��\U��ޱ�\п^:+iZu�>p�พ�n��=f �۽�U��ȃg�>��1p�ox��.�v�9Y�#��J�w)k�;*���)6�2�t�p`���f���hjTf�Bs9Zf:,�ú�cZ���������,�I��\��e-�}�wJS�,��4P]u˩Mq���:`�Vtڝ�Q�ki�,BH��t��q�����J����W��B�۫��!K�Cwyp'\8V��/�&���p��*��DK��j��n�{����;6�*���U��x�ˎ���R|f�<AW��ƱZ{E���DsJ� �X7'�h� �����]Z��=�nЂ�ϫ�����h3b��s9]@���j}BO��M")Ӱ��y��);�C�T;��G[jl�s�u���� s���2.;�*�\���H���і*<�].��Y8,�:�gWc,��sᩚʈ���O [�}��� O�<�����eV6�Qp�u;���^�X��iƖͤ��V�V��1�[ڮN�``ہf�lF��d�Ltm7FT-�Q��d�g"�xGXU�T��8�skfڂp6��z
��T���=۶�ٗu��T[Bյ:J�;�&u�J�W�̝�[�Lf%Q�,fmf9nҙ�-�A]n��2H��λkhk������cS�Fpȵqc�턯�� ��o۠��J��a�H��]�,�J�gGP�uX���UHGn��Gc��Kw�k�չN�4"�1W��{���1��m,�g}�ž��͂��Ђշ�ek����!�`�ʰ8�W�RVR�$եK+&��Ss�|�\\��T���HjV3.�X���z6*�����2b��^��k>��v2����:�����vrE* 
�B�G�YQdTAL[*��cR����1QD�+m�eE�Kh,1-�T�V�DE"��EV��F�Q+[j�"յ-�J�q�e���m-*�mF�
�1l�UKiZ��(ضV�*�YiD��1)m�+Q���mB��V��Z��j�V��TkAlJ֊%���j6�T��[�T���Ab�R��h�Z-KF��e*Q��U+\%Imm��-j��Q�����K[**�m*-)Eh��Z1�)m��[V�Z6	�`[J��[K0�[iX�Up�10�R���-��Z�����J��Օ(�V�b�U�m��R�YA�U����2��Ja�0�m�-j�jV��Ģ��b%�*V��$+�
)*�F�AO��oº�f����� ���#�=��bVj�[n�zt�V�ek�u���\�T�%-���8M�0Ӿ�Bf<o5���NŎ����e��\>��7Xg%�Q9�b]z����TG�e�ck����d���[�7M^�>�t���������u������nj�8����YA��ċo��q��)���Cz�x��88tu�s�r������ݜoO=4F���&��y+�����S���=󕕚�^�H9�|������O2�r!�&i�_Q�6:G�m\U��cD��t���f+ز�2�Y4/�{����9	��sW�gZ�8(�ڦ���ͼ��CթP��&ɻ3婍��)��8�ć\�+����^��G
";ν��"�;���1Sz�ޫ�"�"tw���i�R�*&t���2���ʫ:�gf��d��5m�E·�4ha)�t�n���Y%�.�쭥�=$�-�P����n�ʗ������fXǌ���z�B�]�0q� r� y�j���i���˜n���A3����oVu;�\U�t�/�t�v{C�L�=��̋���_�GC���Bo��Ebs}�/�U�-: X��۱v%������r��&G�;+q����9E�,��p'����̥���ح�"gWo^���LΦ\���zˢK�HH�_q�*�r6;��d卝��}�Q� j�L�+R��m녺��OϬ�w�b6O�^�_¼1OK�p����Y�Y�$Ƌ�tFŶa��u��*�]K���n�oG]BفL���x��J�*�S:h����Vtnъ�E
�9%@{wm۪�s_7�w�(p>�>�ͺ�l��'�G���p�ˑp�e-�v�tU�s�}^�{�z���(y�ls�7�t��ʱ��X�ϸT@p������h�������2���^���9yt�ӥk�
;�bz��^ɒ��b�`�������o4s�\C���
�=ږj���mE���L���xP�Q�A��� �eᠭ�U�=��$e<�M.���1M�@�S�ѓ�V@�wq�
�S&-��r����Y#�d!6��+.�si��>�VZ�lc9T�`3�]=^��X< 6t-�F���/ep�\�a��nl�d���$7��u��ۮ�0ATa!��K�����H���K�Bsۺ����l>��#!��I�f�t���3ϱQ��y�&�Ƈ��B.�*�L;�uD�[J֗��~�N���D��\319+��W���kk������em�mlY�f���b�:N\�]��9�SF��vUJG�y���ى`�Y��$d������ewaD�����m?�d��oP���:3U� mw\aaw��YS�/F�76��q�������K�v�еT��3�����󩎛a��LH�aq����C>{`���cQ5��N�/V-�R���^���T5���n)q�.BȨ�'R�j.��it��&-n1��s��������q`ڮ�5h��(lOs�92���0n,��)h��WX�z�9�=�۾�@�:M_�C�eȾ(?!��`veD�T�w�C��@���V����X.����36Gl�n�W_rc{C�W+3C��J��\^
�z�@�B�R�L���#�:��}����e+u��v`��T�0[�E�,X��$=��%t댼�����􊵹�u/9_�]'
g>��ȋ�Xa��hhpS�rP�n���d�����R�R�]�f@�Q]{�[�}.�|g/��&��EF<pSՂ:Gy@Ǆ�!�:�6���{��ԍ��g358�P��]��9��`� �B°�����x���g���E�)�U�ך�$DHːg��Y�u�ᚽJ��i7��x崜Y�+�O�;��2*~g��^���c#��'���<�,9������;�k$b�L�p�4��a[+ºfU���-�킀E�ɩ�ܷC@t����LԹ@ Tjh�w�C�'cb�gt���{��L�ҝ��[z���w_'�i����c��1���zgK��;`�U�C�Z�z*�H���֍����8=�(=���]�[�#p�̸0]�K8�Z��^ؘ~i�jqn�3:���V҇��A21Pq����м>�h?-��:�w�{yܰm�⚻ʡd�Ƌ]Z�;����0�#���B��:޸g����d��ow�����0�t �"�a��v0�oWl����g���#4Υ���8*�U?fW\{�η���!>,�����m�`�'��ĦP���ۆ�C�p�뱥��"=E�\�U\�x�@�9�$�z4�kK���:���/����p5�`�-��>���x����y����h86f&�H��3�e&e�we��rt竄_I��,Pk���~W�,׉JE�*%�W�{F�e�g�}����h:�����3/)�y\F��������E[8���N�MV����rg��oE��~�"�-J�w��\�]9�#t�M��E'M�ɫ��K�����b�Uw��M;���NX͊w ���o��]#c�����n'PT��傡w��ȸw,��vE��c�t����\e��sz�>�g:̒"���٨ϐx�۲1;�H۫I��mlC�FK7�J}:�N��wEg��v#f�HUo$��C�L��Gw�Y<x���K��9m�	��t���^u��6N߶�U�;�]�^pU�}�T��xm^�gK�: ���6����5Z+he�yE*�n�	+�"�`�r�\2KGM�=���ѕR�����]UL�����@Aƙ̃\�����X��RW�
JQ\�W��}⯷_?b����Q��z�b}֍�i|y|䯓z��Kt�o��v��A;�ȶS��*�{{��\� C�eh��5\��k
�>a{U�+�ʚ���̚-�3݃P��d�.y3C����n%)������u����G_�Ş���H�G}L����B2�:6R��U���J�4C��8_K��u�\���j���(�f���ץ0�l���C#;1�S����>���U�c8P���f,�ߓ���<���r�
��c�;w���l�t�����<���ȳ�,�#���,��	=�ep{P�S���4I��X�;է��;n-kuy7����b�TW�^K�YN��
U�g�,<Q�:�����Ӥ"����Ŕ��P}!EEyJ�,��9-�/gU�{�M�*����R!�e�sU� s�h3q�ʲ2WW{KS:���3�ܺʞ�G�N8�\���3f�7�ŕ��|���|���^TI��`T�.�nJlB�O���}�͚�j��cu���7w�Φ4��CO�S�� �dCa"tK|�+OR��u)���4SIyy*����
�R9�;��������.�<�fՍ��{e�idp4�f��zl,�f�[�Ƙ˫[�n�O]O&�R,,h��o�e�x�ɼ�P��sx9T�;��ղ�{R$�g=�ч�B`Ƈ^m�\�C���|E�%ɶ�\��X#�����Rxu�i���:(Oz��b��_��w!��֯U�`��ҫf�$Ƌ�荌��JIY�ٿ��=�ڮc��l���@U;˰�q`U3����������������:}�q�p.*���_�b��%z�l��:�Y/-).�r.�������7�\y2aOA���JEM��1�w�2M�H������K|b�N���B=*������ע�G�������-n�t�޸
6�y���NW��K�d�LJ��n�a��Ջ�����%:q�C5�����Y�2�[�Z=5��-����<t��ZQ�1�1��!�����`Z_E�2�MC�l������4,h������T]G�;�2	u�|m��}�]a8�dY�SE�(ؽ�h7�yeu�f���7	���U�������YW׈>�z����f�ۣ�»����Y�	;�j'���ݮ������!z�J������m��d�"��˝�fB�ɶ�ӄw��}Ŭ��c�eS�w��9��Ly]vU㸓ZU��H���IX���ߖ_J�V�(Y8�(�|oQ�~'=��~z6�\��HH��s�\[A=���nea\4�c��X�;B%椰+"|�<������k���ߗ��ʑU~���0c�ɺ�f�覹�s��3�J���e��J}hg�
�����30��\���zWox���W�2�w���0�[v=���rfgC����h�7�����<�k"��	{�1�|��FU+Ԓ˜��'�� ig��śUܦ� �(g�ݞ�_]6cL�Q�صw��v���
��s�@ܔ���<��\P|��U���G��"W:Η4����z�ٹ�㶎k�`�͆�X�e�t9H�����K�\T3�غ��٪�
256Ǐ��ݑ��W<�a1����f\.��,��yi!��I5�]T;=ZY�Y�~�s�ec���}�M��i���wjܢ�6���� u�	�nS��u�ۧf�0�mq+3�x�W�׼6�����Sz�����_\����4���qɖyi��� ,���%���o��z;�	h�+C,�x�vҝ,ַ�w�%2i��u���9K�ȹ\T�ەi����:�Ϣ�hg�
|�J�DCtz �(c7H�2Ai_z�r�Wqy����%v�y>��۸�;֜п9���=X#�v�a�4q	��ol�5�x��OAzs�X(��G�m�x/�m��(��,+̀�XYՑ�:s�҂�Tu���zQ�MuVH~A��@�md��8�6�ˁ~]Z ��[G����%o,a��ny&؀z���{�e�9Ѫq�K��K�C������܋:p0l=btb��'�Ko7�[�/]s(?:�(���Zw҇j��|xT-{��Lm
 g \�#ސ9;��eiR˭t����f�cT�iCYQ��T��������u�X�v&᭷�ŝ;���"z��87Mq�if'L ���X�����wLv�w�"B��j�~��A�|�Ϲw0Ŋ�^�
 ��K�.�����9l���o1;ra�C��c9K֐��)DO�EUq�.�����c���v�z���;�x������3D\J�ޙ�+�.���~���k\�f-X�й/���<|o�	����w^��?g����r�B�Ǳ�-Ԣ��Q�甲.+�V�r�LO)̝:�{��n_S3�$IW�ZKw4rW����!�VvV� �}8�jƹ9���yݭQ:E���z,���TZC�N�z���Ҽj�uw�Y܎K[�����p��+|� �^�$P.�:y-B��2�3,e3/��a����<+q�=K{D3���n�'�2�ҹ���9r��a���A���yj������2+��KL��;����v*���K3���zl�co���B���o��V6άoܓ��(�c��ۛ�L��&3�1ngg{���\�b�W/Y�(a���`��
v�o�J�y���q�ܻ-��������O�P��Vf�����B.K����
>�>K��#gfOo�,z�F�C���
a��Z<��%�f�|'۾d�Y�tx����S������[�h�g�*K�8]{�#	�٨
�/������A-7��>�̀޳�"7ڷ\�Wbߩ�7cTڬ�۱X]2^�CoR�BYty|� K����v����^x��^^j��{~/D<lyǈ秬n���a��ck�,�m�%���͖�}[�tH�|��+�i문;*��o݆�bb�te��#�p�R��wY:���¥��S����I��yj�r�}A�2ki�j��s��m�יv�[�Yɂx��Ņ(�>��KM
�=R�N���36����&|�����n�mY�Y�w4e�W$o��&VUM�"����Ơ�V��똼|\L���K��l*�����2�K�x�8��wcOI9��ϒ�
�7ަbu�;�:Y*������ݓ�;�S�;�.������T�ۊ�L�m�+Ǫlw��ǵ��!'����\1���e�w�~�>�jk�i������ɍ������^�C�
���c����I���~)���0��C�)�4�y*Ȅ�tK|�R�=JRd���b��SJ�󐙭[��h�J��~\d3���6p<���L-��H���p,��^2���v^�Y�7��펁�u�/���ڦXMV�7�wa��/&��B�3[�@t�U�U\.����MOUcƛ�D���B֔��՝N�עU����KR��X!7�w���s]u�W���m�P�0�(tK��du+!��`���00pz�<�;��T`ł�������r����',0\8�ZJ�JG��\E$Κ8{FT[XwQ��*y��=[�x�ڝݲW��8e��ٜ����i��p^])6���� AoPa�pZ�غ����=��V��|VD�v����N�>&;�d�iK�q�"�U)ie{5Q��+���i+Z��o.���zK[P�hp�[��kr��.�"���1�-������9\��n���p��T8��8p���/����S��v�KMNڕu[�놖�d�A���6�#�+�.n��������k���V��a>oj;B��w���+.�w�����vU�N�*e���I�嵌�6Y�Gn6��߈�R����us졷��el���u��AN��u�œ��}9��xc�����Xz;Hp	q�珫�;8���̷P\��
�&V��sv��w<|����=:�B�):�_V=��`�]5\�n�J�z`����a�����Ǔ�����dN�
Rk�X7sf���ˆ��<��鳢�
���&�zyD����%;f+��h���ː����0<�:���D��3I���z@鎧���Ηy�!սAS�t��jwn�O�㮎h�X��a#�;�����㲅�������������M�E��a�P�[۰�!�h,[��cO�<�@���Igp����w��n-u� ��Ur:*K�3��Q�B/ =)Od
q�E4���ֹ�c?���J�
ݙ��Ļ����w}�S` WB][]z7�z�	}E�o#�L�vup�{�yZCO��$��B�n���%�����.Eћ��X�����kE�bu���+�|�z���z�*�Yc���KJOzK���^ѫǫ>�����Qt.�˽�Hi�;�%C:�m؉�0V��r'Qdu�w�ù�M[���8 ݦ���Hi�t�Vg9�rZu�naA ����Ȑ��y�.��x�q���ޮ���Yʬ�n���R��Z'lB>ŧ�J�y���m��SWJ�Ժ`b|�{t�m��Y;g���.�m7cl8�%��Y�w:v�ܚ�C(�U��B���f��%e�� �Ɍ�dC2�k���^��1�v��]v8(��1�7�͜*�G���(��;�sM�*ii�q	�w�Rr㋭�4�%f �^���jP�;��C�:8]���J���q��&�۬�=CW�SƉ�k�0�s�I�<���yś�9�S��9�����Sܡ]z�pQ���Jav���ו�h���"�8�����V��u�f�5Pܜn�8-,�H!�#�:�gV����.�,���5tc(�୼-;��}nk�6N�+�J�u���1ϥ�zi��滷���@f�9b&����Ɲ\��KL#�f�V��#D����z��)\��g:�IJ<�Cg�eZ�'t9p˼�#�j^��t��Wt,�:�4��(�* p�ۛE�Ofv.��=V�v`����ȼܡ)���߮76�q���Xҵ7�E�V�ňŶ�m��("�������im*�6�L&(-j*�Q�+V*����-e*��R�kF0Z���%����j���5Z1��Z�U��Vڊ�ҍm+�����m�Q�h�DF�-��U1�p��j�ұ-�ѫj�E-�F�V�Z����(�F��+e)B�l��R�`,�h�n�[KYAm�jPJ���B��X-���E�P�Jմ���m�F�ե,�0bPj"b���m��բYlҴ���+E[@�P����kmŘ�m*�+ZZ���գX"��-*KmR�m��U`ʍmKh��Q�F�TT�m��-�F�(��V�4�����Y�pʌ��D��-,���V�҃m)K�����KYT��������1��,�m毜�{�D�[�'��fU�� qrt벜��ګWL��',��%
�b�ل�q1[I�W��қ��%���@F�>n���|_�%0�����r��f�霉G���on�z{(���Ή�P�h��Y��
d��9�����Ky»��������U��iZ��7�R�!��mLP�[��G|����1=K#�D�ۭ��V�����$x5��ې�be�{���%��j����bʋ�0,9m,���zP����%��:w�J�	#�j�m]��1I�L�n�9����׬3`>���B��W*���
���m��[��'��j��*�^�X�e-X�t��x�k�Z��\ޔ9,�	Y�+���Îh��������<�/�H
Wj'ZV�p5�=M�vQ��qpvS���h{�r��eƳ����yS{Q�}OU`a��y�&��t)P���mVy)R�$U�����:wW%;M32m�.Ka��c>Mu�6��0�+�j����j��o�sZ��$��̛��}�\��Ζ�����h�7���C�<�,�>5#��}K���h���&@�0�x���v�z�	��c8��"��Ok�ri�����|��	��ܖ,�d^�Q��z2�Eo�#��;s'h���tc��en�l,鉑ݍ�Uy�ڳr�W4�{�*�W��A��"�㳯�5Й��2�&���Z9�F���eb[��kp�uz���|�׈PNY��&�V�;b�\=�xj507�)5a(y���d_�Cg���]K�:(R�)��/�{�7^j��B�ufK��@��R-+�\^UC؁.�fl9`
)�;i�75��(f�q�lʇL2��.T"Աb;����k��U���;s7
�yKV�b�n�F�XcP=uw���������!����xM��3�ifM[�o��a���O^�0zr�\L��nh[�6�dt�ؕ��7ܝ]G���P�Sv���8���=G}V)�VP��y��m��6=�XW�nd,��� �-^� ���E�]e�x.p��ma��8�6�ˁ~�բ���S&�wm��+�V���jC��������Ds5N4���ǥǡ�O�Ɔ�QuIu�չ�[j�:�{���N5�#/8�&/���N��þ�s�,X�����A-L#�<�"��󻹮;�� �h���2f�MZ�
%86S�,'���v�տk�*Q��B��`R��߇��߷���,�P�i�.��:��uj8���o k�+	Ћ�ÝMM�J�e&�x�?t��6's�y��I`�U]�^f�}B��܇^���S[(>�N�f6al��E�������S�����g�]�?�������y�C��ξt�bu��t�s�b�}K'Ty�av;̑�s���&+w26��䲗JT�1_3��\�`��auC�'-�������A���\sk��^8��|Yu���:MX	3�eUq���ⴈ{{I�Ӳ��غ�l�nA�s�n�9�W-�����1��˔�X���RfX�v^U�/�S�+FS�V���l$o3/+����{�/;.s���v��H�T��\��`L��C���_���|g�d2¬i?#4!���[�On�Ne���"�V�,K�"�-J�w��W�9����gk�j�����P>�Zw#���=�b��"��g�*�*f�E��:u� gFs�<���lf�"IV�B��3���g�Qs�I]9��踖��3�%k_a̧K`�֕u\ ��Ep�f�G�<�f�UGr�U�)(n�	+n���l.�3�`s�j�z?J̦Mr%���c���n��
�h�|�af��_�g���F:x"�t��T/Fmu������{>!U����BS��u(b��ƅܱ١u�uͰW���(��v�,˾cV���3�\zmE�⎵WLr��`�[����0>�,���U�t��]�2��ˌ��R]H}Z���ܦ�yɒĳ~>�|�:���w�9螭��k��0(6X`�:gR�r8_�r1>�FϦ�0#��%&8*v�D�F��w��t��Q�q�0{��V�kxJ��p�-̷�xG\lN��o)bcbNl�u�0���F���Բ�e�ʗ�y�G�[V���q5r.1�����>���T�^��$��w[m�A�T��s՝Ug�h���*x�:�o�Ws�r������ݜ�i�2s|
o��R��w�����\���.��+��,ţ��j�s�g˥�\߷y�Y����D�6��_��6	bV�,�8GG�O0� 6;�a�B��A���i���Ϸ7�%gR�u�^�3�x" Z�����
ug�����驑ԝ��")�X��ozv��t�[���Bs���Tޯ�]t�b� (Br�J�VWљ�yy�ʛ��K���j,Fc�!�y�������:��l���.�#Adp7��YK�{8��_�����:9�f.��q7�쾪�Y {�PyM�\�(ƫ'�CMM~Zu�׬�I��K�p�5����뙸ȤU�cu�lT��,h���t�5�y�Y�j�����u���̸VʱԂ����r�c��@d.պ���*Vi|�R�EECg�t��O&�S,,h��o�e�x�ɻ�|$��k�h��3�D�nB�Fd��q�t��bsW���1z^��R,k�W�X���`���Z��o%���Y�4����<�S�(l��:I<*`W]o(���C6����*�^5ȸ*"yu���.�q_i�S������~�a��S�e�K�t�x�
WI3�
Ϗb�jϞ���H�Y�x'ww=���b�cWlr��yo�30O|_�%ɗ<4�B3c�t��K��;�t��F�`p0q��ȝ�X��`�8� �5R0��p�a��v��M��OE^t�4�2^c{�g_�O��j
�R�X�>�`����p��X#�EM��g���;`�ަ����V�RDJ�~��{5qͻ����;hz.�����O[<�g�m�Y�T�1��t���Ѻ�m�&'�xg�����o�'�pWS�[��}��+ K��;~��j��vsN�T��\��{,��`vi�cs�1�+)֕d�q����i���k�y�Y&�d׻�l�*�ι��.�7h�.�w�w�<��s�
���[g�R���V
�"�`��.�Jd��"�fny]&0	E"�p�F�-�{%,޾����컾	�u��y;4�\�SQ������i�-�Е&fM9��V-7����p2ZǛ��r�o���};��*K���Ǽ�f���"���Z�)ނ����e�&����8�3�uL$�:�)��x�M��9��[��n��h(a������k!Z��T�����v��c4��\&�2���K�l�����ˁW�0���J����g	U~����0$��Hֽn�u�=2F)a�C��x�ȶ�9edk�Af�i<�����注�Aƻ��I�<H#�:��/���mM[��L���g��ﳖ3ub4�1�}�i�;���MC�eȠ/�j��@:�L���Y^~|f&ܞ@��k�r��LB�}r�|$�6e�u�E�u+��^P%��`5��{9�
bd�κ��5qz��W�sR����Z�r�B-K	=�!}4�T�.�Ӓ�l7]|������\�61�ޤgXax"�kK�V�҄;u.Ȅ�&��>�{�i�霽�ψ�ɑ�<Y, b2���ȑU�c���Ȩ��Y`ۂ��#�n�W˖7��u�r�r�p���)�fђ�3V�y8�٨+)^s1�WV��â��N�,�Y�)�K���:��|^>+��|���ťIV�Y�JFW\�na��V��� ع����{['(7��HΝM+�e�����(<�Y�},7��,(wR&>v_M ����!�դCX������l��{y��B�e���s�24�2Z�h@
�n�o]؃���3�hSǳ���׊�\L��mP�Ղ�.A�vJ+��2���rB��N��z {ؼ 
�{U��?SX�՘��,�\|��|�ך��c�ؑ[`6�>YtHpQ������&/;�����v�V�ǃ�~A]n�:�	�0���u��j�v��S}V`>��/m���������(�v��x�m��5R�C�2���3���9:��Μ��P�JHh!oT|S1AZY�N�(|K8㹩�<,.�z��Op_jQU�_4 �jΥ��ҡ�X�(P:�K��Mp{r0�b�S+fAs�I��gz�c�����u��a�g`)�92�9QU\���u�]���4<z���95ꔕ�}
�0_L��:���s^a"}���v�X���US3���
�؇A��T+i�ts�,ft������D	u��
4�Vd�9�d�]q��ҤJ��/����_ �Q��	���	cI�g�;�:8�sz�m�����Lp�����'N��#/�b�9CI�n6ZRWb�v����j�H��.�M�+l��Gy���ط%�,G��b6s�Mz1ü��wQQi���R��M����F�pV�{kc���kޗ���C��.��L��{Q<�:�8vٱe�`��������ܻFP��9�잎zr�����7�[�T���u����U1q��z-�.�݀���VT`����y,TI�x�)MN�吨X�KWt���\C�����Tt����i+ӵ�������t��na:p-�h����
R߷����5ƖxL%� o���R=�|K
?_��W������G-6�^��O��j�C�Cr��u&K�x���[0���3�3ٮ�s 5蠧��0o�(��g���r{2�?R���Pe��}.Rc�e���^鍴��ģy���3�rke�k�w��'؋ �e�+���N�`�~���
!�:�L��ɏsQ�q���PlWK�͢YӁ�O9�M\��xcvr�~kA�H[|���qv��ɎuX��s�/��;o�AW��ݽ>ɾ!]w����KF������c������:ԓo�vr�/�Uo,�*�ԯ삅}}A���E���is��g"��`����s�*:@����m�@�#��*g�S��woT�T0!"��V�j�HN�����ao���W�&u�f̽�rkb�o�rt5�[���/_U�*�8�m�.�7N�8��27kZ�HQPVӛj8�t�dwd��fr����{9W��ޒ��ks����60�B��S>�|(�����`H]u��"�L5u;�9��[X
q/�XM��г�7�U�F��*���b�w���V.�����&��e��*�V�߂|�<�x9�`p�ڊ��6�eBb�q>���A���yQwy�K�Ux�����n:�v:�3�psz2�[i,g�U�}g�)vg�s0��mٸ/� ҵ�����*��DRB^|9�=��V�-�ܢ��}�ڇf
����ƪ��e"bQ�a�\�
=���U<9=�;ٯX�OoԶ'�n+�k)Zq�Om&z.)�>�a 7������b�;�t8K����<��c|���sJڸsJ
p�6��%�F��R��k
�^�p�aെO��X��*��g���Nu��8X5�����g������kAAZ���׸>�r�{͋�IX��\8�b��+;evoF]]m���qq6�d�+��GTj4�r75 ������b�1��8_fL��;:Z t:3»��')J���wr�����gb�pG�7�������ݕ��u�ipޜ���G:V�KU����5��o���꼨��Nֆ�]�T#��;�:H
�w%�[:A��ʀ���G)��e(=��o8É�s�X��W��Gwu>���fɳ(t�X�r����՝E{��k�,E���g�Nq�z�u���Ѫ���m�oe���bV
�n�R�ٜ]}�5f
�y�H[�K*�qK4�F�5��5����7���r�W z:v�K��c���1�	�R�um5s���'�T�3缵2��p쫕J���v6+ܺ���坘��Q�1�� a`T��	�X��^�K��y����퐉�mOP�A{18��F�q�»{��:�w�E'˥WH��U�k-��ՙ�����Ɯdq��E�f9T�>��zRy�����x����76�秉
n^ɝOg?G��]�>�bcUGV}�{��{����$�b��$�8B���$����$��$�	'���$����$��B���IO�$ I?�	!I�B���$��B����$����$��$�	'��$ I?�	!I� IM@�$��b��L��Ye��
Y� � ���fO� ĉ;�>�թ�ڶƨ+j�h$Ua��A��2-�Ud��Z�mUm�)�ؖ�V	�մ�-�lE-6����im�lı�	�[f���FC4"��H�S[o�.�݄R(	P�I��T�RGV:�$M�2U�M
�(���kQ%T"D�I(5��٨%	:
$��ְ#B�R2kc+lR�^�֚��ڕD��P�kfƂ��J��	%M2�**�R֪�0��j�H�6f�5"�VM%�m�kT�>���(� O���t����f��u�unwv��Z��,)B���ݝJ�Õhn*ƫm�;������T�Ue6;k�!OK^�w��t:tX�`�iة7����D^�A R���  o�|�*�Q�����˖ձ�Kmݥv��ؚ-ZP���+���*��A4�;hP�ձmJ��GB�ʔ�F�Z�һ>�XYj�)�UP��D\   1B� P�
�� �
(t7�    P�` :44(w	� 
 @�w P�
; Р
]]�i��YP���}���#Z�ii���*z�R!B����N�   �a��ڃg��W��[mMowG+{j���U��ʦ�.��֜P�����]�N��+hjae�k]�͛-��R���6���"�K�
UP�Ck|  <�*T0�Q�_c*N�e�@�;H��B͙��Ҧ�0mv�髲�r6�UlѶZv�T.�jj��ww]����`3[��R�T��jQ-b�>  ����GZ�j����6���v۸:j�1�WmA�[8v�B�T�,�h�T�c-�S����U�Vڕ{[��aID�)�2���dh���| ����l��v[z�N�5;�sYRB����)T�SD2��4�f�u#@΢��Z�
S�om�7s\�h=�I���D�`2Z�  -�P����*�X ��T��Z�,F)N���  O^��]��A��u�S@4�Y		졒��lĵ�  �� t@� *����pt�(�_Z j7@��F� �0����X �0�B��u�hJ�a�d�-���G� �8 �CX �+  3&�>�浇@5]� �P�f�e�:�09i�C���[(O�Lh2�����{FR��  ��J @ j��	RH5 4р��J�4 @��L*R 0x������'��C�J�G�����_^�M&��!v�+��[�-l�sPh���������$��HH$�	'�$ I?P$�	"H		�|+�>'��#����jW�/��f�YR�C�ZT�&j#E&dҘ�|�"�dİ�Y��������hKU6�i�fX��@U��-<�O�j2��r����b�B�Q�kK5�!Z^�!sr��.�#[�*�<�P���;fА�CX�3�ؖVު;`�y���2L�qk���ۢ���=��=�H�0�ćhɰ)գ��./:˺Y�;�Y8��t�otU�[cY����5�Ϯnǚ0׳��w:OvV!�w`a��Bk��2�����U��<j\gJ��
K)CI�d"�}i�/B��6�ӵ��x��6^�lR$�M}L単Q�)�-�w��Q�n]���Eۢ^Ɏt��Vu.n�ҭk��2C6���A��w}c�:x�i�a��	�N!wi��Ap^m�3�i6�jn�v���,˺s~z%�I�oB�x���A;��bӮe����2)�$,wud��64���PtѥI���)��*����8�5��4/��,b˒�9I��)5c�yHY���&�
֪�`�=��WK$�fmv������#u2���^Ћo%ԧ���?b̡1�ѵD��2�M�Աݼy��OxS���d�七 ї��{�='.Hܦ�wos��^��3�+{�$�wQ�;�|(r>Z�j-s,�C$.=�)�d�J7�e"�Hi�q�f�+e;&=�[qoU`.0@��{�)�8�d�n1U��mל����%��+K�3d9���%���L%6��.�w�TBF6>܏u5�n�LkP����b`�mQ����&��e����-}�c&:D�%�Y��{r�nމaZ��KŔ����r��]�ҟ^�\���5��7	{#���Q�C�Xz��hX��i��XN���CH�V��1��/*�J0^d�eB�X!LV��V.�cV���m�T��B0���)-�Xi3f�����`;RԵ�Mg���Mǹ�5���ڰ�Ԍ��&�b5-@�*e��1���d�q[�ͬ��Q]���w1����z@�A�h��2&-�)���\��]͚
tR���m3U�j�2���Y���bL��X��z*c�b[�qcw��o �U��O+S�6�ۗN@��ͼ�GbÚav�Ob��p]�c��&�� ���_�+{A�R1�y�J��|�j0wcv�&㭮k�#�{��x�ڵwi�)�.+26�A�/F�6b�ך7R�C�2�Ve,�u���zIx�v���&Y�7���\�pJ\'�l�7-c_C����H����mba��C��[� s��L�pО�v/���it������j\i�(��-��o"�Z�p���\�n|qS�^i���T���w�uZ����7(�t��v��kUQ�ݷ�b������=��k��2���۹*��7UIOd����ͬ����4���2VW�/dvp�lPX�4����&����(�J5���,Y[s�V��-�4�BD% vMyS���J˳�5���ةz����rn;�ưJW��ܲ�q��Pb���@(wRL�r& dsGgv���#�m��ψ`�-tX!��􋜒�G�	��{�1��H�;��)��LV�v�0�/5=�Ѻ��F`�����f���/�;�DP���p�GXE��Cⶳf�YHNH���Aټ4A�f�C��gv�d�{.��
d�-�R�,�K�]˦�����Y�f���wtۊ�wv��)�uJO�̂9��;%ZCj2��yv�v7 `�9��ʊk�u
�������l��n�i]Z�������[�a*$z������)�rc������>����JcX&�.c_%f�I�۴Ubb/�--PN��Hi�ne�e�2JћR��F�*�-�:�L
@�N�m\a���T�y�X���X��.�\G6��ٻ�v�2^��F;��\vN�QǑ
��u��4ܖsT�	N���di�l��j�7�3sm��'�h�����o�Jˠ��j�7 hJ�2�
cr��e�1�X�S��j�n�[٬&��w�
�M�$� �x�)��2�h˳�����]�!�d��-�P���.D)�8�vd9^��;*��� l�ɰ��R���T7��P���!TۡE����M��tU�F�i�S%��tR�)-ݩ����d�!dsu,�ʅ9�Ah���w	e�*�7H�̉�Zn�;k�s��gv��vD'ѣ۫�?0FPZ�*ՔNE�d��\�]i��^R�.�Si^B"�[�F����1����$	��NSU��fk�w����#T�67B�ː��7��q�9�n5��NqF��Mn*kD��d�9���;�B�Ex ������m��~2:ʳe]EP��hj���]8�ʌa�De�(�`�Z�՘�$ت��c���6�+b��0�b��a�kZ�A�f^�������V��[[�ZҢ�b���$\٫]ʄM�F��F���:��:��-�S7&�9� 8`7��>��EcG�yti:�q�fL���(�ԐX1�gG��)
(���Pܙ�{p=ۭK�!nڋ�w��y�Y����Emg�{L Bɢ>*�\�VV��Q��F����w:��b=r<X��<@�7D�����B,bM������5a���r���J0��t]��5���k{VƤ�5��6o-R�#�i�%���(n��u;�#�.��)�G.��6�� ����i�Ô�mPɺ�\�x���:ʂ�-Ɣ6�3vi�t�8d�6k
��"ʎ���`fN��-,ד�Q(�c,\kwc��;�U��Ya�ó�Gj�6���0�'[U�V�6��]���HdMX��X�뱚�a;��y+�x��tdCF�lG�͇VEs`���ʱ��D� 1��@�
��²:'���ޒr4bS�I���U���}�]�.q�ǃ,ķ�He�L�l2n6FY�����@f(*)�xRC���̻�ZL�c&ǻwd���Ҩ��.�k�d�J��v��Q�Ȩ�SKo��4.�⺅�j��L$6	q�����m��Hw����[t��5n�64�Hۯ�#p���h�P����q�oZ���ͯ9K,�v-Y�u��c�-�BY�҆}2�ٌݤ%�`��:�t��Z���H�F�1*������ 	5[gr]F�:����B�_J�{5����ܷj���hNe�p��85(� �>�d1�7v�5��2R�3vu�xg-�M0Ž�.+�Y/!WzӤ���s-����� ̬ʻ�v~r]I��M;Q�0��3:p��D�p;�a�(q�2���л�+��8I�-�yŕ��XLŠ�0�S۶M�Ӗ�l�Y1(U�Sjj�DCVY�O���[o��w���v�@������82n�{��6�m�a(�QCp�D\D���6 FRd�E/���K�q�U�K��S�W�$�B�3��m=�Y�D͔�+"�d��G/ᮀC	�ͷ#ܓR!�3#9*�H��b���۽�b�l}��1tDkwr`:��oϑ�I� �bڇb8+�R0�\ŸP݀�)�2l������S&��ȫ3�e:,{Q��Ȫ"��`82�wY!���vQ��)겠�S�5��nG�`*ΑU�Gl�8��)��]4��uj�\��jŰ���}�(@���	�ݰ�	zZ�B�݌�u+��we�S�ևs�mQrG���/q'�����0 ��h7n�=�訣��-{�Q��7w/HOWE���G�T���d�/��ww^�U;w$\q�{v��ݐ�z��a���2��Q�Pw���.�e.��8��h�,��J�J���@&]D��RF[���5�jS�-�A�W�`d��-҆m��S�b��u�DK����zzL�q�>���h�r]�m�U�/kɏ��:+�7̹�J���h��y7�������n5�f�����ɴ��X[BI�RT�!�R�t�ޛrȭN^�P����+�l���d)�XPτ��(���Lf�Jo�歂��\/a�ԅ��ۮ,,'�zj�6"�zCT73T[��c7�7p�3Gli��m�!Vu})����Qɦ��㇥&ٴZ-ӳ����I��y�H=M��^������k��9{�[�����&��ڴa����Hn�(�C2u#8^��f���N�18e_:�Z�O���',�e���fS-����z���&�H+����,���ț4j��f�ܧ�W���
C��@��FU�� O�>�D�	�D`ҖϩZiңyn�f�F͚lI�N$�o5��ލ��t��*��K29���!�e1B&r���74d&f����ux�1�8T�>�guv��:�m#�4`'h[�11�����;t�����H)6�I�tr��2j��,82J���V^�t���g.
A��B���{�o�y'TR��L�%�nB �n����(�<}�q&	�C�X� �<k���+4u��Ze�Pc5%�U7x7pd&�e�e�(���
k�C��,:0�vm��䛃�d`ʲ����8�~���	o)�^C@�OM�˦�31X�N��;���7������AZB��BdD�0<�`��c�MX�2�Ó#�R���u�G҂x�Dk=�$Kt��	�R+N F֚����ʑ��;]�Ɗ�\���hh��(�r=+�w���,�U��K61��^)ET[O�pJ̸�E6K�G]���Rj��B2�p����9Xr���Ϳ�Q:/PkVfF6�I��1��wn��B�@�n� ����p�udm]ȥ�af�A�A	E(^lyR�)��jiMX&���q�R,����o�o.d d�˰һ��훉ff�,���e۔R�t`%qcl�l�o��c�|-&�}�M�,�����JUHV��^i�'�a0^bd���8�#gf�ܔ���7�5� "��2�e�j�匄�����0e�qզ�1���_]\�> 6���˂e1��,�l.��l���`=ػ����n>��u�+��j��ֹ��1;��棲]��E���0RL�Kp��4F��;{$7(��zr��˙��'�$$�Gb^yв@�)(8�nI��\�'f��Q�ih�*<�)�07Zi�dX���c۶�����6	n�����P��Y �Tzկi���3����G$�w9^��:`FgG�>�!��V�ra����8�G�wVKHv��-4$���	�j�{t��/���V�̬�$�Gr����n_��n����6F��6 �dŘ�U�l	7l8�n���&���ҭ�V�l�RV�
=���V�OM5	*�ǻ�sYua7e4�W ��Ց^ؤ�XEu�8-7s3j��z�T9��y���Q;�̼Xn��'q�"��)0`)�ѱ�ì�T ��wZm���֡��r9@�.���Pok�]�И���1�7mnZE�r�p�e���1/陏�PHe���b�2�3�m�TT,�;h�,7��^R������"��4�(���tj����z��\׏3V�t��"�F�lqD30��]���㲵�lwW�+{-\�K7)���2�U����P��q�/4v��9�������흚��8�u	��2Kh�FM�t�G]()̫��m�:���u-l�b�nb"�5��ܤ��۲	y1⡖1)W�]b�-3�ۋ-Ñ04���P����Ǚi��ULF�^$�䯭��q���<�=������U.�b6�"0\q;i�Iq��(���ZMUSqw��V%�DS��N��h#@�0A�&�ù/u���XM���N�
s�F�Vv��Ј�a��eT̐�UdG@�ѦQ�&f�ܩ�jL�.i�4Ҝ	m8:�rdȎ�63,t�r�����aYTӖ�FAc���H� V�3�[x%�r�f���pǴƮt���M�*�ik��[[wbĊGV�:`�0[]��Y��w�۱mcY��%h�;��u�G�vt�VK�T,��i�!��C����8%�S�)Ҍ��� �;i���9mcߡOr�;�I�'.3�o�������J<YYoTn��f�*7�h���4KŅkn���9�YV�}S�G(d[!غFt�w[V�:�qatٯ�w��U�Y���vM�����|s{�*ul�o��*Aq�yJ���f�I@`�xޝi
,�aPy/1�u7��Mm�5i�|ә�t�/�QQa8R��g5��φ=k/D�"7s����8g	1^�@�z��DG�&�e��k.��P�(r���^#I��p�׶����P����$n�#,���nD�[g>����'Mvd��*R����u�(�0�Ҹ��hZv&fD\�˰����������m��AW�Ky�PM���s,;���$]Y�л)�&7�r�s-#6˲��S9�*��{c<\ʉ���zI��I��86�]�Hk^��m#r�)�
�Ae��� ��2^��WI��9[�e�u� pdRD>B�ruK�5p�AX�vh���s����r��2�QA�֦�C�F�63bw ��K���DC�Do������:�w缕�^K�)�ɩG]kM#b+ܒ�,CKB�T���4��2jy0mɆ���*^�]���y���y�^d8(������蔏��]��k�r�ac�x�Z�{�1޵W�a���8S"q�Q�\!#�qT�5�4o�c�^&L���x�.*�L�#��#Uw�q�*c5��FQ��w�B�/{0sԉ����\�6�MZ�x�v(��E�x��] VF]^ǔ�*4��mD�޵���\��Vv���}&qg9�6�����?���xG;C��%^�=�.�WXq�#pK�!M���yꞘ@���x4ٲr���J�.#E������y�����=�d/5]Xd+m�ݕ���X7�2�|�\/��iLn�uhͮ�wo2�S��X�n^�s��<��/	q>�]O��Yg�c��۠�ʙd���GqZ�v�+��51�},��J;ۘ�|���u�Dg��r���lU�WK��@���V�҃29������9������ǅe������޾�/��l���q����o����_ �$�|��jٝ����o�:�:��EK��h�)c�p��m'bO*WDzn�hv5M�X���B��8��uP�h�ef> �ɦ�r�b���M�c����D�*e�\��D2������AM�y�=�/��#����l0�uy�}�G~n͎�vse윯�R��yF_E;��r�E̱xw.͘�8�_Gr�Yc��®�r����թV��j)F`��M$e ����^{��h��Z��>�L��y�8.t67r]�:P{�ov�t�kp�O�uj
�
�pc��^u
�t���[yR�&�Xj�T����;����;���=޴u�'��P޹���]�:����v��������:i�"¶���A�K�Jb��Y[;���"D�mv[Z���?e�ˠ��]`���OK�ӭ]�/ �L��7ۀ(�ReUK~��H�`���IR�Ԏ.��-+݆��<�a$�1Q�J�B��N^.[`�wG�c�;��J�H{q�f�S� ��s�&r�MK��'V�c���t2�Һ�ͮLe쬽:�>RS�bF�.�v[2m'�}���V7
����^-��z>7�k�#���W7��۷cy����hے��K3P���sN��a�����?���*�]p�(��fY�9Z@_A3���}s�p^�R��*v�.O�j��(!�t�Yf�C4�.%�y��\��.�A��,��M���K�C��b��S�i�Y���
W;�SZlkn$F�'���ۊ�
;s�R�޼�Un�̥"fP���1^��B	]rk��!���n8�M��u;�����i�ٷ�x%޵�f'ZpՉ:�k��D ��=\�2���<�������7#�X\�����rY�srv�]kK�9����
ƈ�D�;�Ap���9�Lw\5��R�nH&�F���m)l��K���҃&��K�v�if�Ul�e*�b|)���;�%�-.��J]��&����74��Np�|��� ��4ê�$[���N�n:��c��Wx	�E�I��ˠZ����c4��9�s�g��P����z�/3nS�L辑1�`�
�`�6��	o�-,<�G���|9�9Y�}�_���5ۻ��dkxS���Le��*�yt�z�ܕ:�����zʍ�Z�c�6�JK��Ȧ�eټ�[����!��5��t����y�Ixsި�隽��û���U��.�<��M��[�8��"���x�c��xw8"J��UwyR�vF���y0��u��i��ڕ-�:'���kA�h�	)�}��ed1v�ę���
	T�C����wFq�&�����
ΕF�7I�++X'>�Vv�.fᦺ�˦���&l���Ƿ��=�;,d�-���8�c3"�Nu�no
6��-a�|���f��Y���<����0ɛ��n��v�I��m�^��yX4��E�ٟuZk���uA�4�Σ��_A���,���H�td��z�BEc�9u�ن�a�����
�_|3Y]�������N�f������![[u�%F�z�TV�4]�\����"�`z�p^���^ �dk1[x�s�դ�z��mpA��j3+�\�:oL�^VwT|n6�`���N�5���m7��Ţ����yC�rXx1��Yv�^��̑�Ց]+X:���S�K��I#"�v�q��ܪ�n��R�ԟ_^�OO���W��W�Ξ������Ъ{�E�4C�S�z���uă�I��ox�O,��K����:uк��b��P5!���zee^æ�r�x�"<H-�az�L+bY�q>$t�
�����*�]U�
|�~Ն�靿3;�.;�d�^�v�A�U��>�Z��9V`TgG������f˼Wl�Zvwl��M�Y@`#�B��`��|=���8�r��;t����T{fbEnY��'���)�M���@�p�nݒ΂ܕ��!v[�b��k���VsU
|�\�n��G�S�����Im�n�ޢV�ׯNV��N[=�a4I�bF�!��E���f
�z�­Y�c��^	[C�2�p	)��HF�#Φ�ʽ��I� ���}W��_h<��>�wYϴ���BZP���T/;e��	�c�a����3�i����:�(UUAk߻Y������R6����p�:�L�}��F�[z��ŏ�$\�`l��N�Z��Xz�.�'��c���.��zAk:ɝ:(��v�3.��O(E��T�wuK��f�X�4W;�*qޗ�͒wQ�lC9F=��ո7z���Hq)
���ym.���Է%�_��u��-���2��$�x6���q��gT�k_5�	N�����؇u�-���@�8�ثf^D��C�ݩ��(Mf-�GD�r�ؘ��5rj	W��X��::#>k4P��ƾAU�o��Wm�яc";N�pZ�b���T��u����u����=�'��T�%oВ�0k1g<�{"�c[<��{�sE�p��uշ%3�<�SC�.�ݕF�Tx�Z��.dK�,���ŷy�˼��e�Y�}���ܮ�j&���x��r�+F���Ջ�ٳi�B]��@�����7r�qj��b(<�,��l�2��	2想�	�x��thᩭX�\1���[����ٮ��0�|�d�����cA5�6w����J�*�_u����/��t�g03�n3�i���9�i��N�Vd�`��گ�Չݶ���VN���B�;��2f5�R�ó��X�rSu���۠�wN���|֒��Q��w�u��
�:�ίce�G3cŹ��o��XRG&D�^P�D�+7���Dԉ�r�Z֪J�̥S�4�ڂ�86������Lf༤7�돂ڳ�nd�O�һҳ�b�h�w�A���nYf�T;�3��ç����im�Ф�K��o��wufb�HmdL>Xl��Ւ��z����6UNvQZE"�"�<����_7�9_�/���F�t�C1�xgIQ��h��X]��d&����^�Y��w�s �J43z���w-#���������y�.�B~��-箞hq��=U�����:ܪ+gG�Þ�[9sr3���KK�v9��j��î.� x�kn�U�\1kq�*����v<��:�*�"@ݐ��Y��+1ڭ���.��t3���vaԷ�T�J�j�7u��1tuVQ��ͮ�_-�<ӗ��RM�^ÎTc/&�h�w��e:Gn��w�7�J7ZVH0�����\ҵ�v�������p�FU�Z3^��㤂�)��S5��F����̌�U\UNq�)���t��b�QW>�Z��
�`�	�������|�iqK K�j3��Ko$������CjB��YڤCy¸+\�et��n�^Q �����A�À�p|��Meꛝ]��J�s���p�[h���=�o�,;'�]���ka�+r���J�bWK0nm[_9��^[y%􋚳Ƣ87':Y.ZL�3cŊgw���y-��[�堁[����1���F�rj�cL;������J|ڻk|���ƻ���]�;�!���Ϝ�c��N��Ny���}��,�e�:�f�+�b�OKNcf>�q����nr�7O�ΡǘU!�']]����&��ϯ�AAl���{���jù,�q9�+o�n�WV���d�8���A�|�ҧ��[*�)̫��e�.�NP>zG}3�4l�m���j�XZ8�;M����]hJH�D��`=(0�wAr�2���U�B���}���75���tB�����yƢ��	]Y6ݚ��	�����
5+2������i3��d�b�40͛}sO3�zT�Nv�c�x��&|�%�)�Tǵ�"vq;���p�.�������k�WY{��{I�/v��8�u�B��sۤ����y��*����YXW&H���npF�b+w;x�)3Bgl�u�B5]ʁ��/Hq9�s���J(R܂��Ϊ�*��F�z� xn-��C	��o�+a|&��\!�BX,���:gY,���mƦ_�eP�0���|����a�[T�ӯ4Ӡ��Ɛ�*V�;؜�u�����o�N�������5�N�+�Gכ#v��Y8��z��8�%������9���`�T���7�B�JX3����s�ͨ0�v�v�t�8]sT甧F�ڸ Κ.�"�ݝ�qy{!x�uJjN���Z�X�޻��6�ʝ����1��Sghǔ�xrq+��,A��m���`�xz_\��n�2pdM��s���y����9^�A���cr^t.䚮]�j�Hp�9-�˘]H�۾#/ze����s'�r�}�j��_=��nd��1i�x�9,V�<��/0^�/s���i�E{:>���5��x����8P� �!hۗ�|kv��v��ʳ) z;��%��[����S��4��J�$x�TTs���<��|j�����t������/�<��u]�U����p�����VL�%��,����/���Y��tu\����Bv�3o)����ƑB�w�ٽ���'o��S]pH��r	Z�y1Ìe�dǛ�Œ���B�r�qOY��n�`��q�j��K��Ī.��˳��8f�0���L+����o��oox,�RR�4�]ӈN�I|�0-��|Ttj��w��ۨ
'i9a� ھ#�]�-�j�c|���r=\�!{�gjm�{��cfHX�"f�z�s�oEvP�}^%Ը����݄�.��Mt6�6�w�p�C;���F�ޕ�9ZOg�fަ��f�h���"��9Ƕ�'t�灦�92��;.�\�M��7�r�󴜩6�:���q��l.�r��Ӈ�M�$�	���P�����f`�5Y�U�ɽ���\o%�1-��Ҳ��gL�|JA�%\`V������amsʌ�x�PC���v�����] l�xY>?kC�$qC�u�@��,����Uҝ��k�J9�_��Y�y��ھK�V���2ob�Xl(��Ӝ �lu�)��
X�(���
��;���"*�t�N��3kv.��#u�g�*x�J�a����e�nq-�gVA�K���%]�^�5<�+��]��l�|8�:E�	�nq�PC w���$�&�t�����v��m��4*)�](p��7�pp9��L|;o�C�yJ�Q,:�ׇfŠg�qBh�+����c�	��{�7H^E��'����8S�cU�j�b��Ͼ�|��af׏D��+vE�tֹ�}�\<�feg(�YɌ���5�a�Nq��H]l�v_r2�`.�unFي,}ws2��+brd��]��@�ڼ���`�g�X�������V�3*���p8.eeS�S�m
J�vY�� ��©��vokn���&N�"��] ���8�G��L5��d�U��l-��ۉ�����跱��y�;U�]���<����>��x"̜wvo�.#��s͢z�����sm�&4�N���m�[��j�E׊�̃�сxV�4��S,V6Q��K����Fl1vj��՛F�w_#bTeBU�e�z��&ݖM�f�p��9�-\����R�s�Vvl!�V�[��9P7o!C�g��Jn��ʝ$}n�/��w���<���$u��+�8+�����t��G�y���g{�!��Ͷ�
�۰>��u�u�Ta\:we^�D�}E�o7y=�����c\kܔ+J�έ<j�\�w�&EM�ݖ��L��E;�r$��$�[h:��b=(O���6�9N"ƚ˴�\]��5�Q��w�T��ʖ�������s�-�:�7������H;7t�D�x�z��Ѥ"�,A_ ��.ə:�	��՗7�~Eni��¤�&u8rp^����f���x�Ds�lx����n*5�[��҃r�~����\���O�v;d���W��GJU�s&R]$��ق��\�s:�ej�ɓs],\v�������[A	d}��3#l�QN{���4�yH{Ϳw}
@j�y�3�<ée*1��Q��S+�x�>o!�%5��;h^�}�5i{Kc��S �3���mKy����Rű?�[[q��.�n�)_WX���]K{�竖v�
n�m;���l˭!����":ӡJN��T�}2�@�a�0\�t�;r�Y��R`5�ˆ��\7�(��&��	�v9[ݙ�{���VIS�g�]Й�~�Vv�&aw6�}�,��m�	��7�>�4���|sqɺ-:|�Lm�݇Q�C%Z��k��jd댍�5���ue^p�w^
��C^^�6�E���,驚�v��W����#��9�'J�\Yc\O��	�)�S���롗f�
������M��w��e�0u>ڹ�ks��&̪7���W�5.���M��~�������x{��{�ݼ��,�L�}ș��z���`��ƅΡ4��Y��5��9)t���e�<0�VWR�&h+v�[MW�c-�y���#+ph��r�^1���R�+}FeY<+ks7K�����Fuc������Ĭ�m������u-�F�t���S3��9�+Bf��VQ���q��� ���!]gp�ܒ�[r�N�a<��F`�}]�2���������'�f�NO�O ʛ3�{��:c�����H��Y�9t��<�ޥ��y���M��F�D�s�[&Y쮦J`�� ��cC봲kH?H��[қ��ϼ��i�8p�jg;�D�u`l�ESܧ�HU�xs�6��r魂vt�v
��D�[}4����YM��tc�!p���X������Ӎ^N0�p����ִ����Y��Um�X����<1Mcv
�{wf}�Ꝓ*F���-T�|�`�W}F���L�)cp���B��;���Y��:L,x�
�np<4��+�_g'�%�2*=b�'����*v��r�`O3+;M�X��g!9Y�\��l%�R��և�ӒC�L�[���s�n=U�W
��j:[�;�ɊA/�k��]�i���Z�[2��m�]�c�{0�X�8z�%�Ҥ�!HS��u�+OQ�.��s;��� �6����#��w!˳vO=�������Hu��ر�K5.�h-��Q�E��]J��*�0h�����wp9��M�J��d������cYB�&�*����|�ͅ:����nL�M.zceh\Ix�N�X�Qaȇq՚Af�]���s6��jgFS8�CU��ht*�kŝ�f�u�t+�r#B��쳤�Be1m��N^�:��K������։C���ŷ�ԣ�������H�+p���Z����	��Ѓ��'G5��_/v-Ã��ɏr��ܢ]�qU�А ��Fu�yb���O%6L�y�6�z�7�������܎�\�����U���4s�_ZO^ǥ���,1�+�8�������r0Faz:�aPu+*����fÝpt@&sS�o�Vv)��6���ˣPcD�5˻�`��?)uW�J�w4.A�u�&��Un7Ԫ#6Z��N�Er-Lam�;�F��e��B�c�ے,��O��X�]�'8���2��G�s 4��zr�w!�o���r����'}���RD��[�6�M�)�� tچ��g0Ne�2'��4��EY�d���d���rm���n�wRU4��d��ê��Gcܒ! �$_�oa��9�S�����z��Q�6����uce���/2>�a^s(t�)*�7nB`[�%`ݠ�F-Ͳ��^AP:����E���Ԣ��o��r�*�c�#|U�ܭ��B���V��ᒍ�c��:��o��N�X�����c�t�N�>��ս��b��Ȳ�hV������g��1j��V��y�tɖ@{u"H���&]����뺦�
����3��<S��[���)�ޝ�j]�Gy�ޓ['Ў=���ƽ���fM2�7�ho7k&3�:F���^XՐ�Z��ʽ�Bi�uWN�
��dm����r��w�֖3�|�%����l�s��<��L�dV�"��l|s���777	7�>N�lۣʅ���/CۡHe��2U�C��i!���w´��v$�wU�Y�*V"sJ:�Z�Ll]��6#��lڙǫ3���˹�ĵ/�
ҙcSu�h��s���Mˆ}�%ٌSͣ#��`�W��l���a�8�-��{E:���.�ջKZ���r[�a��Mb�Pk�#)��<O|w�P��ݑ�Q���=&-�vdÕ��8Om����8^���(W�Ў�����y�s
����a�݅Сn^�ܢ�iٷB���w�wH�a��E7$;�z�`���o�t�#��k��gW�R���2K|�Ҝ3aEW�"3�te�]W��p��wɎUٰ��+�֞��ގ�u�����H5V�qyI`�[}�7�4.�>�����<��L��:.��M];�/ ��ε�ѫ.�v��f�}VY�VS]��yr�Ԁ��{Y<u�aų�k.I�ən�i�|_c�2�;P��c
�w:.�r�R������pG҂���]��p�&�b}}����*��A�펧ث�pq��Y\�8�J3�̷���i� kO�������\�Ժ��<�6�RL
��s���I=t������6$׽e6r�+��.�.�UC]�7����5���۬"�����yl�t�짻 ��.�ea��n���EKGfhH_o
��F�kn��S+��y�ع,:X#z�Sw��{s�)�Q �L]l�ǱE�L�tM���t:T�X����,�VG�D7I�O�M���9��:�D��G�v�v���\3���8����(+�9��C��0���|���g��;:�8��c++د#��R�Π3&.�"��vG\�k�h:霼;F��ke:��s����:�p�m��׺�q=G�a\ޤF��H��I���+����<z��6��+�@U¸�[��/�gt���΄�z($�7�=�hv,��]�KB�ư]���<�!EL�3C��-,6'g�*�w���>�\���X����4��ES��P�1��H2�Y�<x��Զ�E��
\tQ�+��:D�t�7�`��7,7�oyb:+s��*S51�璬W7�孡����c�s,\��UAY7q� �:o�R���@�D��C�5W5��*E�V�VoD+�4�6>�ڬ��Xŏ�\SOk������Ȇ�8�0��x{'���!�^�P��,Q�Q�.<v�ܴ;׹��PNkr]a{0�"Ӓ��.Wl�O�.�Y�L�B�����R�2$��͂���J��+N�W�I�D2��V:��B�5�7d�Zr�wT��*�u��j��G&��\i��v��l��w��oN�Q�0u�6S��n�uT$��M���SSVsj9}]�I��NCaHy�8x�qJ�w����v�P���7EH�Xz��74̻,0�w-Zq���w��<�݊�Un����,�� �ܩy��(�ѐjf��}0݅O���7!K��[�U� �wA溸IH��YH,�n�y�˟p�C��t�\r̽r�<���Křp����L�x%bo�<��j�	�l�Ů�l>f��%*�:�7.���4Ywժ�A/�����*ɤ,���^�&.����2G2Q\e�ͬhY���9�:;O2����>Y���LSיR`�|A�� �M�������Ya��E�;3����v��9d�h��7��m<<��/6ݭ�y�m�1S�:�8�ȃ{ݸ-�aL.��a���8�|6��p��!�!�kG>�عo:��Բ�w#�;8�bs	v�t��r���v�+��(-�q���TA[L�'���7$n<%ݜ~j���u�)��j+�.N9�-��zt4a��8�	N�{�6LF���Fܫ�ΐ�e>�sw�H�+����c@����-��£x��чyv���=YVU7p�Ɔ�	�Y0�#�ϸV \�]�ane՛�v"~�h�4�u�"]!������{QoqG��6�?iyZ�c�I#�f��n����4F�K{-v��Vv��7"5�������:�����ޮ��-v7�3��V�riJf����Ņ1��m(BB��
�:�Q�u��^�-��ms���Ʃ$2�����k.�t:����m�W�κ�������K'	a\wWյik� �^\�S�	{kX�h`q^���HҖ(�'i���z��D���8)=!�����Ж�m���WAV�7�KW�g+�pVv=<6>�la����6��ΔNp9���2s�u�{l�ꪎ��v��d.��6�k+]�����Z������˔�IG�@K3�k�e;5��de?�qd�v�8�)�K`��}g��̨����3w»po��I@]�.�Ʃ�h#@�IfG�P��1F�8N�p���b�46��B�̬��)k׆}.s"��[��8���{�E��=��c�3�2�!�m㎥��,�̮�ю:h�vX������<��:�z�V���4o��3]f	bŅ<ݪȳ`[L[N^�Q�
��Ï��!��;4}���-�C(�v�	�g4,�f��R|���g:��� ����\bR�1X\h>.�Y�ȸ���cB�Ew��y�:[E��K3`�u�q�����6�6:}^�UHj���R���a�F+*�B�a-�<urɶt���̘j%PWF�k�S����]����f-J�t^lј�ۜp(qu�-G3-�VX���2�Y�ː:	R���<u���o����"��v.���������kCn��n�'�khmbl��9'e���M�%[�/)a�`��{S�[�3�i�U8WE��b�S\���s��ݔ��k]�Ɇ�=dͯ�EV�0�f��1��L"��md��4d��WR.<���^Fq6N���q��f��b�͂�,A4�]IdnV�#K`Ӡ�W&ug�o`y��)v��%Eq���(�{��]6�1v^���,%�hg,X�N�|B���`�P�ʾ{]�(���hv��zඍ����� 
�EG���]�5��"��N�Cx_X���P��X.�a�t��:`��7K���M�o���ł=��oa��	�FL��_gU�y� ��2������J��3fA����3�Г�Ż��&YM9��
��L�էlQ��dDKn�iS�����1ü�d�X�ga����n#���'�:[�]��;OH슃=ӳ�_\�=Ց΂R�:�Waa]:͎ ^�8�|����}�0��Z�����ߔ����ہ��n�v(D���l�V�m�pW#5�g��KqR:�]ء�6������5��${�ä˜�M2�l�N��Ӄm�\����գ����r�#׏fŦ�f!�y&��t*��a�Y\FR�Pۣx(��Y����I{ɞ�;l����Qc�� �V.�lߦm���zf�1�?m�- (��C!� B�!]p
C�v�(1�]�7T�3ݓ�� �
+Ǆ��׌`�b��`�ʙA[�c{����Ϗםŭ�A���
㎝��:G=��C����E�%a�E��p:��)}y2�B�V[I�4�9����N�/l�����F�(�e�cN��4�e���[P-��6���:n+b�n�Mݹ����"K�ī)GW.e֥��>��t�
�!wq�M�e^�6�56�ϕ��-�6�1��l�mf��#!��s�q��t,���~�Nsok��ѳU��>�9��gT��W�Y̦�]�Π������)n���b��S��N���jJ���:z�J.5fN�q���ܹ�����E:�*֎�HI0c4U5�Q��ҳ��f��g���UԜ��ɫ�ۮwE�Fn� ��l���C�B0�Vɴ�me(��/��)�:������א�-�$�rZs��u�Z�,h���֦kQ�w�=l>w0���J�j����L���Ybܽ�!iI��}����9F�������M�;�n�*�ZW�xxN�ݹV�R�-#Φ�X�ZlZ�X��B�6����ĥ�/v���S��s�r�a���N������Ѥj[��+�@·q,3s2Z�
oI�գ�n*W�eN�'��t��U�W1#�y˝f5X!,U�+j<����_m��LRb#6��3Հ�i�!��'-Wna,k�w�괄�2�Si�c�)|z���J�ee�;;��lX��:�Y7Wt��B蚜��n�`Ԧ��)>���v�-��+��ΉZ-�W@�J��ٵ:���SѮ��l�c˳�o�a��g�c��Uv�{����� r-:�t��s��ՙ��X��He�rMfS5��fZڰFKظTcs�0�$�c�{9w�s*؆S<�7%�������-	A�����&:ygs:�΅������Z6.�qٛ\U��+z�5wD�B���gnY���;�I��4�3C����5ۚ��꺶0(�,<{[VY���K��JkW��9��}E�1Lf��L~�d��N/�s�.m��3ws��eg��uɗ�&xs�2��ixv�jE7|*��Dd���Dqu�G�d��E�Ӫ��h)',�"�7$Ӛn��ckM5�֭�tnn���{�6;Z_j�/m��R0<�'x���oRV]V%yq6WZ�t�9/�:1vm�f��U�6��`�:��엑�W�����p�̖4mEQYj;ҕ�/����a��wL�;�,����0WσvI�J9��Jv��6%s��Y�ve7R�V�b���u̲��a�*oE�s��{5����m0�M�W��<��vqn�/nzE�/N�g@�9B�x��L�x��cC@![%˫,�eKAB�W^�u�^�)`,�ڲJ� ���ݱŭ��s�En�Or�\�������.b���.�R��et%.b�
�m��XHߴv���C��A=\W9S��88]9f"��p�����cfP{r�9VO/��m�am�T���7}����u���	��q�ʝ����XN��^����YwAp����!���1�w���{��!��Ȭ+,K�M:�PvW`��2�=������`�ZB�+/�|-��Yy�7�9�[�<�V��k9����}&�
��0����D��o��8kU}��U��R��Ε���Ў˷sq�£í�{�xv���g���seb���1|T�U����v����K�m���VBb�8u�
gJ���D=�Qą^����x����|�Ѡԏzao�e	L���&q�Tԑ����Y�O6�$�	&I���q��F�1E�N�xl��8�ͩF�M�4��e�w�aɵP?�N�}oO����GV���n�E��x��ݠ�ǩ��يh�Zo���ǲ�u�qS�jY�h]je�발]{մV�7Ny���)��ޓ�g���r���%7c�/�d��0���w���6��r�c�!�g�Y�~�_�7�>63�����E�m�T�D�=���?���z��+_�B��}S�L�%��t��|�h�F��M���E����}��#����
�֜'\��Ye��lҘόSK:[˞�y׫�;��ͮ�]Ys[���[�J���5t%�y�Z=���z�����q ��'rY�C����gv�yO�K�X+��Z���6J����L�8H}�Rh�˲�WTѳL�7��@@��v�pf������O�)���j�f;��b'�*�����������&A:;˸34Z7��f�S. ����>��a�U�2B�t�gj���6�]����z\�c0�KP�K����\.G;ͥ\k���n�}4̨�.�,-��gq�>�F�Nu��v�껺�I�˵��ܻ���s1>�T`��t��9I�����|E�2��`��ǀ�<8fYp�{#C/f�ݎ��D���}w����V��o��������+���2P��&b1�5M[�%�v�:�9�H�$����E��!!H
ST"�ȭT�UR��E�TYBJB��
,��PXE��$@YR*�$Y)�AE
SP
H*0���P))���j�	LYC)�����B�,��HSYI�H"��)V�S)�EI�@�PE����j���Y���R��)X)
E)��H�!*�)�E"��e$�Jd����)L)�L
��YU@����R�S)�����-0YhR
Je!H�2�RE�))�IH,��R��IHA ~���e�<m&zoj�����<��Q���wC�q���*H����J2�*F������2]��L��㽗]�����{����?��˧�3j�G�� �o֯��Z8�&BSc�o�����?�Iu�`\�,��^�X��}���W�	�ό7�Xx��I�Q��M�������̽��X���yU�b��CX�$<��kt�H��Q���h=S��q��������dbz0a8�]���B��P�9y��ք(Z�Ʉʿ#H��Y(�����^,-9Q�H[�N.�K}S ����y;�2�\�s6*psf�����tƎ���yl��Eه՞�+YH��Aݳ,&��Tcٺ
/UI�͘���� ���4C�j.!�V�l\؃W�T^�S���+��Ws�����v�6�r���t!K�v�Ó��m��G�_$�4���`k���((i>ȻUqlӃ�f�Bl%Y=i�1��]�X+�zg��MFx�0���cw��K�:��w�VD���>,Ut�}M��,-���n�]��q(ɋZ��ڕM�;|ś�6���^(e����c&%\�5�W*|{��k-S�3���7��j���Y�]́�%i�[3>k���y�J��Z�b��nfꝨ%��_Au0�\��Ta�0�3`���vJ�r�yt��+��9�:ƴwwF:Uǰ&�eNO']�1�J�H�N���\̷�����;��-��k�b����gG����:C�N��,�^�0���ӀW��C�1��G�y`��C����^���o��u:�	}P�߶��y����	�2�lg�EAO����3�>�!+Odr����VΧ�g<s�����*zq�	����|�0��[n�Yu�w�����P������sL�`}4� ��̊A�u�)�h��@ȣ][l�˦ R����r�8w��cR�5���BM"$��j���>��Q�mSr�\:�f������(��q���ř�t
^��
�	Y �"�z(;�x�ĭ��<���E)S�A[x�t"�n���̮�\�,FțӉ"@��6�w�1:�2)lk�����;-���^`�!S�}�W�ܗ*�����wg֙:fԸ1@�
�*�����)��]�u�^�6�GM�軇\�X��k����,�s~���d�pBs�Rm��siqIwR�D���8[Q"Xa��� v��A���#�qUcUL6��H�QR���T�m��wW[���-@�j�D�>���wu{b�D1U�m1�!$e�ū$�Y�h#E�2%�h�w����f��Y�ӱ"�Վgpf�6�5�#��p��eN �e0l���57��\:��D%^����\"p�w;pγ�.�fm���GpBQ|�e�� Դ'Ђ�[
m��7�{��ӑ-MnOZ�1�$�a�������N[�Q��Q-J�Lj{�bNa'K�V"�Wj�����x�S�,
M����r�=�Ɖ��vQ���b��g�U�}�$st��њy`k1Q�,�r|)f,�u��}����&eR��{&����Y5�<fㆅ��˟o���DG'��/=����͍.�u�j?o�K�g�;�3~�t��^;BN�ۻq�*�ga��
���a�'�q�W?5�z�^{��*|�]'²��`5�U��E��Fܾ�P\�e9Kν�S۸�!ei�r���Z�b�����@�A��=�K��0�ɦ�k��k�v�����q�"邺�0�����m����NX���(��W��ԧ�i�aߖ�p�3��3]�a�N�˾s��]�\8�Zj8R���us�>Q^e� �WKȑѴ�ª�'۞�`��)�"R�&�5ܶ���c�E{�{�#txc�U>��Fz����e��i��]Ӳ��:S���{eIނ��_M�� �%Ӹ�=��O,�L�Aƭ�Ŝ��C���сL�1N�r�:�+������*[(������)����Y�Ջx��H�s�BҺ;�4��c��;�w��]e�kfe�R�59�r��i4�t4z;/8rv��ɽ��h�^??D�h��q���#'e�dt1ζeE��l�R�%��@�VKW4ۜ��e�񌀧!���3�
+Dul(�ݎӝ�	MŻ��l7[[�32�*G�%ַ�W�{Ҝ����嚑7Ϛ$:� <���8�?&\<t(�MY�2��w�VK�jX���˿bT0C��Ћ��PpzCHھ��b�_�߼�W�
VX1�MK���OV7z�N�R�zʋ�U!��=Q��3HK��:劓��,T�MȢn���i��o7�PY4�3юC�0�����!��f*2�/p~2��� ���H��B�0V�f��8&��e)���8@�ns���,y�\���Y��;BDL�i��
VJZ&4>>�|�y�U���$�l^}W����[�0&Z��Jr�y�n�;�q�g�������d�R��'��>����ꑐU�NC>�.6/
m����:��m����0����u�����w�����nE��T.��t0��%k�s"��E�Ö�����Y^������ݍ�ޫz�|�S{x�F�(��Ȕ.��b1n	�Sܼ3u�Q��('M�YC��Kd���)��tp�O6t���X�=z�X33f��a��j�:n��kg;s�\t�+��)�h��L����b
�rh�ƒQU��B#	�#7���&)��s�z9��S��CRb�=qd[^�z��5�7c��kM���ɺ�HJE� ���,SEŉt;gc<�(�}J%XDt�_0��i�����"�<������ZZ7�TOl�����F�)���7u��޷��w��=`З,ÞX�x��Y
�Y�i��ċI�pYT��j7=α��@/o�GZd[���,�Eu��or����G��F��'�SP�U�̨ﭕ���Q�?�7*6=���h�L����r�q��Nx�(��/���{�A4���K�ǵJ\t�q��c�&��L��p�.����rAYJ 7Ne�9���ʂ�z������ye_��ƺ�/��2/ ��8��q��9y�L�	�9���e?1ZGr�E�ZÛj�1�s�w;!w!y�)K�mD�p�x'~$K�r�âp����k�1���B�����5o��|z�*�R�{F=�t2^��/�7q�X�9"kX �o{�w�6eVi;��6��2��B�Gy�[��<��h��oJeO����wg���v��������/��ޜ7��r��L�S�D�P�.0_#/w��c��S(�w�4N��v��lw6��x�[��{ҖMi�AG��R>}گ�<�̭��u|G,T��vj��\T_A��܋�`0S"��jW�4�,�Op[��R�15�%��4<���'��>ȻUv��㾽)�����m=xV�Mդ�^����0�ڽ����I)�u#�zn�������+��'���~�0�&LEL]�o_<1QAK��p�26�f�������)���J��j�R��{�E�'9r�Nq���֍�T��whp�bw�~)fŧ�ttf�SG��ϸ:939����5_`�%��syʳit�꜀��>�BS{T\�u�r㔆��	��<���՗G��C��k���]f��k��x���9Hq�=e�&b��b�|���U�{0���N�8���-����z��`�^��z�,C�(� ̐�k�ִ	�I��3�����K|����tk���+�&5)�|P8���_��PV���S�Iު7s��h�[��z��Ю�~t�c�z{XN�Y�~R:�a
�	U�|B%�&R��_��j�����С8��o��i#��
{�vOVa������:>�5V?|}c�Z����Aآڷay��<ut3x�z�I,�G���8��:��w{`BqJ�*�D��dܳ���IlZ2r<�;2�4!1��s�3�=<����*�<�1��Nv��|����o���S;2��뚂#dKr�`��Td�R#aX��Y��;N��~�(t���nt[������wg�'Lߔ�1@�
�;������7��S
������b����C�k�ok� ��̵e�zY8 I�T�bb�a������x�@�:��NϜb�P@tƢ��#�qUz�`���(ш9/�M�	c)�Σ��m`��:tA�� Ҟ�8<�KC��6`>���s����[C����s��[m�5��0DJ��;=��>�'-M�%���|8< �K�L�U�ϊ^��n�˓����!Jj5K�጖�b���@�L�jH�*�`����y#���}�R)�s���yǥ�9.���h�0�^א!"�G�ᮦ{��/hh�W/A�v+�A����/6_�L��c�Xes��
c�E�!d�]���x�ʼ��!����R���T+3Ez��|�_xpO�v�Iᭂ�$��n��uQr�qQnj�m���R�s��4��j�.�\7sl�ݖ�R
���{�-]-�ku��7MPc0)m�*�jf������*A�����1�����\M9�#�X�j����.��
��up]'w��0N"�f�t�SQ�̠�kd�RvtǷ��:oP�6i,�F���_I�g�� ���Gް$�U��k��uw��yW�,���
�n���o{�\9�ޮ�$ު�yf(G�b^i�w��c���]���nIO��Iv9��ֱ��]�C�j
et�$i�ι�*pc_X#��k)���o��=��ҢH� ��.z�Tې��P�v˄;�h�FJd�+��=S6�0��[��j�W^�d��!b�E�5�����X򺽗x����fT[�8fֱ�g�������-Zz����{E{̎Z`aai���xx�۶�9ې��[����l]���WU=�g7����e���e(/N�51����r�x��P{Ek��8v���]ي���ՌQ�-�]&�~E_��F�>�~��|<�఍Hھ��Ɋ\QKm�wu��n8�z�T�u[���d����w�{e��Rs[���҅8��Y<7���;��C�׻Շ�O>0����V+�V�=������f"�͔6^L�F@#��M �..��l8�i
9���}۶֝�ڥpU?�u�X�4cN�]��k����:��,cr���B�afa�B��ڷ�V���&N��1D�R�G("��ܩ�pN�����n%�����e���М������ʎI)�0������^w��ȱ���|:�ka���U��=���2}8Yv���-7`t�U�.��*�4����.��ǒ��	�**�Z�Gg ��5s�� �������X}<ЭR��:�wR���B.M���`�ܒ�V2�>�ح�H�X'!�S��P#o4��Ϋ��5��%���N�5:i{ԡ7���@�^��U5
b�_>M��>e�zi���-~�t��2������m0;6��q�Kzt�鶥����B���Z'bK���13#=|���Q��҄v�I:��9Z�����Ie>�GP�U>t�,s�r�h�z�'���E�!��<ni����@���
����X��o�e;�g����6*v6�W��I���lH"Bb�ǫ��a�(�9α��@zz�rt
��m�r�r�L���_g�W;3l���ίV9mG����P<ʋ��j/=l�Ҏy�a�F����T:Y;�{/��ˏV*���Kȧ��!.$>�T\\�����)���U�]��+�C����o�j�hݺ�c�d��u�`V@�����\�#��^W�v��V�W��5EL��B�b��c��1:O_n6Al��}�� �%e�z^6Ei���ߋ<E�I!�}/%N ;)��SOL5��2�q�������ǫ���.E)?ð�7݁�E\�YJ-ә/�<�b�@�vѮ�K>��rΥ/�ü��l?s����AEՊq�σ9xv�MhB�o�&*��ar".����\��)t���Y�����<�����N/�'~$K�r�âp����k��"z���b��^�Ȧ�0�!���GM�E�q���(�3R��7q�X�8D�g.v�%f	�n�{�lj�84e=b�\X���F��0�.*���\m��3�	�v�޻S[w=�W����#.�����j��|bdW	
4FFCvO�*���e���hOb��D���c�����J�1��ڽ�N�ɚ�BҀ��;�"u1g��t�
�T�TGL�ǰ��<lL]+�̞���n��:�-��g6L�r��CN�0"-�Q�o�*�윆ΗZ���b���'`��! ��A�W�ސU��b��4��ӕ�ϸ:9�<��>�[]{8��J��G$_�r744�P�%7�E��g��8NA��ccEAZ �k���R�]6�e�`�wǝ�}�ZY������)7*m[�m�3m�A♂��c^[hb�S$pf	���vʴ���6F�C2b�G7[��&*�2�j�~���c��Ҟ�o�*c�٤���y�e��8Kk��v��þ�V���¬s[>�:������Sc`�c��Y�/��eC
��'�uΕ4��[p�D�d��)�w�n�y�\��'��r�:AOh-�����,ׁ�[�}4p�]�_I�D���^����v4�w��E�}��Ob�e���p����h��:|�nO����� ���7z���LܫD�k=;7P�˶2�.�]˲ovM�ncϦ�`�;̕�rszga��4�4HBU�,eC�Az���j(��6�S*��S�V��+Ѫ���m:L�I�&'z܆��]�}w1�� ��m�����%�.�4kY̤$1Ӳ`i�8c��}]�j�7e`���n����m9��c�J!O*+d"ٳzřX�c��1[w(�w���89_V�9^��v��;x��M�k6��6��0.K���+��9��u:�`�u�Z6����Y{�z��Yh�b���E��˖�V�"C�={�	�z��Q���w-rZ��IEG3��f�#J�:Z�8e�
h����	��j�W�����'@L�9���h[�]���=C�EN�N��\Ľ�'���=�[,wV�����#����
�����p�N��]qn����>5�IG��C.R+�ޅ�$]���{zl7�{�˩���<8d$&.J@f-�f����m��*�ܾ�C7���Y��Z��
Ѧ ���j���NN�d6��f�Ư�wj��� ���5�+0��$󭧚�ҧ6�G�C�k����J�Ώ��㮵�;M�[ <�����upԗ3�K] �v�����4�h���{g(Z�ؽM�[W���M�z-Ǣ��p{���#�˞�g�g-n��u*����s�q1V���U�Jӂ�L�-4��«vu6fA��+Eu�Jݺʎۧw��b2N���.
�� �;s�R̗�X��)��Z8�fG�պb���]�#ɳ#!N�3�6G� �څoa��fִ�I�Ldѽ�2�]���CO�ݫٮE˥^"s+��K�Q�آz��
#h���%��K�5�װ�ݓ��lؿ���m�J�/T�.㽕�[t�S dx�h��:�W�p����@�Y���¶��_��v���f�Nʽ������y��E4ݳ)���/$\,�wTe�:��6Ü���И���ɮ�s�*ՠ;e4�>Suu����9�{gj�z��eQ�	�O��l*�;r��W��t�F�F���J�:nh��יԾ�ur다Y�����>��%Q�7J�-�ĸ��>�K�w�V����ks�Ҹ�W>�s#����z��ٹ}�CG{��Uu���g��,)��)�
���%	���`(R�LYJ�M2�U% ��aHUP�"����-@PX,��Qb�*�����,�E�4�@U�HS!HJE�E�X�ȱ*�ZBR��B�DH�AE
B�JIIJ��,��"�JA*��4Ƞ��X�M$X,E@�V,4�*�������Y�)�cU)Eb���
�0�X��J@Pi�Y%2�(#��TR�,"�B"(��RUP$��T)UJ,U������H�(� �)�����"�
, ��
d�X�I)D�d�
(,`())(a*�,P�B(E��)��'*�3��������'3-_����*������qO=���+��Ʀ���0ӄ�̭ybR��m�t��d��:S�WN�v��|_y�����O�[Zx�C��~}�b����~N�{)@X'�t�٪,D�v���.���=Ju�j&����y�xc�^c��;˨N�j}+����gD�����@�ޝ]45��y��l�\�Ԡᯌ,0�t

�W���&�L(SҸE��Ρ `��'6�_�(���kS�dZ��(/HU�����5��l�̪�K��w�Sg���jlv�9,�=���̫t:栬Fț�t�O��!�yl�S�Mp�Epu�nlvV��K����ǽ;n��w}�nO�&N�����w��g�k;�X��/Q�2�Xu�{<GMz�]�u�B��`w���!g�!\��./�E�
��v���}��?�<O ���0��S'e_���:�v��.i�̸/e���)
Р>�V����IlW�	�9Rq�������9Ou�����������]i2�t")�)�C-�d7W'=���X�i:^򸬎 7��<���$�?$�ANq����W�ֺ��d���O��.$i�Kr��Xcoa�pڽ�hfYuݝ�.�ɂv�:Q��n/��gV1��
�Z9Qf^�6�@�g��$���qw�Y���p�$�����'5Ɯ���{t�8W�o���H{�]�=!���57��^Бw�� 2���L�����~̛��V�5\�Ը��T�lд4-��ٶ�[��e���j�]$�e���T+��J5P���2\[[n���"����>�v�,�Rd���U��4I:�')nq���������.f������^��Ρj�-הm�6��R��UqVԞ��E��W|Pr!����+�/u�Ʊ�dp����Pݓ�aX(�^p�]3���zyE�s잨̵���5�V5i��;���"�U��$�dT�V���q�����ܹNq�a�n���DizW�{2�:^��PӐᥥ`�����>&�r�]J�LY�8V��s+4�SDI���4�{ګ���]v˄;��.s����i��<�S��0�q����dWMz�(��nG�U����2::ٕ��"nR&��iX�7���Y}�iPy���D�4����3㱅���|��mQ���������vsAg��zy�b��)FV.��/Y>�X��ľ�+q��Te뇐[���R��������Â�����K6���RoS�҆�\�A�;;�y��u��6�m;-�T;{��]��m���9qvX�n�P/�"y����Ar�y�T��b�́����z��Q��:���:T#$!-���\`�<��t6�^7ڳ0*�O�՞���\8$3��N��\���Bp�
pzC#j���*<Q�6Nbd.'��:,�z˜<��{t��s�..ꐀ˚��A�͙��8�'��I���m6�`��!����1���"����7J�S�
����[(j���6D��~�<kյK�Ѣ�ɾ�&�^�s����ezh�p(�۶�Znr�U�.��ʯM4%v^�V�OR�WU�����x4C����ݹXk#Nb��c>�����V�	��X���M�V�׶��T�Q���)(���'�Y�gP�Ϯߍ��Y@���������TD�&�Z�Fe��;���:��g·��}����]bO�����v�Eg���̃q6��8�N�Ѹp/ݨ��G#[�j:�S���!z� �p��W.�-E�!�Y�'�&G�~�ѱ.~�ϳG���6�*���M.�l�$�������t\>��<:�:��͕���N�w�7�D\�:C��ᓷi��:��{�pՐ���̱��Θ���)����1���r��3��3���H����Zw�l�]۩�\�H����c��������^�����,V��ZOGu7) F+U�gB�1&�"���jw$�P/ѱJz�-�C����%�حYՃD��>��wnOn��P����("*�z���p�F��-�u�^* �o�G�����@�t�k�0U˝GL���|Xή0�Z�>��~M��3���+��_�n+e~�*����{|�x�P���\歊w�)���/��`�W�	�zq�N6{/�«�7�9�����8�bv:�a���O��OA����?%�[�8�ƃԥ��dWdʭ��)宎J/��t�[�t]_��C,��v��`F9��)D��l,Iճz�V���u��R��s^����tv�@*mp�ɟWK�r��0օ=�7���:;��]$���õ��{����,��:�o@�d����(�j�2��\,G�|��ms�s�wb�~x4_踱a��ܕ��0�e�A�`�\mȾU0��m��3"Up�+ޜ�����	�W��X�s����BMqf͟z��˪�f���s���CB�����o������,�v��z3z�ˆ��0w����e
�If��ߤ��w��Aۊ��Z���9�A�j��f�{��x�n{Ux�o(WZ�U�R^vd<Wu����Zɯ:;)��Գ�Y�pČ-�۩;�p��C6���8��ئ����P�=�k'.��*�����]i"~�Y=a6f���Wޕ�J�J���+򶬉��q�v��}���mf�z{y�5��jw'`�lgi�y���#]�V3����M`�Ld"o[��C6u�R�-w���(b��sѾ�H@=��s� �)fń�����uMl�V��Y�b0.��u$�NH��j��V�R,T�q#r\!	M��E������9|��c��>����P5��X{�p����~3�4G�>
�kO��L~|t�{��[G�=h�N@�Oi����z�<�<��8%�@���D�:�R'��0��z&�AA�	��˥Iu����w������ج�MP�.O����w�,㸇W&5(8k�>a`!��ǻ���u�\�ab���+�I؎+\r��uyl�&)Br�c���5~N�Y�jG@�/HT�`�����]-�,�av��~�^�,���RY\z�n���̫�\���ܸ��S���3{�ׂ�uQs��;&�"�t�;-ʷJ�׉��f4>�f-O�\�Į���*��A��P��J�W{�!���*�}��ON[���z�z|�Ny�yu�?�]w��au��ިZXf7����ͮ���;F���e\�\Oa9��T
���n<�p�ra����X,T���{u4r���oh6�6z�]����;�3E�<&�H�r��Uk��:�"����^��!`,�s�vwoR��VU�k�Q���w���~n�"��>A1���Y�@y	��2��Ǝ��Po��ʈ�T��ւ�yβ�)M�O
	�玈7�jO�蠅k�*e���0����GkC}Qsw�����tV-���VK�*Ĕ�!���C�4qJ�Ljp,I��'K�W7��_�//�S˞��vm���NA��nW-7d�31��~L�jO1WR|�T���ڰMm�/��(��n9�t,j�FuI�+*N��c<�p�}K�74-aY�#�i+�]1c����f�/�1�ce�����g��-�a�!�v�,�R���z��7�X�J�ȇ���j��x5�:��1}�� v�Iᭂ�(tm��Fܶ�#�����m*E���
��=���`bu}'����W�5�}�J�R*�z,�]���@�m�5u���q��������]��9��q�8��Wt��t�����mG�`��c�#�cӻx�3*;���^+vo�Fٞ��h���żim*��"mF�Rf.�"ыw788�k�\��n���mݑ}o�m��p`c���mu&�6p�|��솺饋q��g$�u9˺f^*}/��+�t��;�&u
/"Z�>]�����Kt�:�E��^g�U�X)����Ѵ�ª�'ګ�%.b��\�ٮ�K|�tΈ>��&�8�EO\�r1J��U!��<%��X��7�,�]���V���j2%��]QpȑNhR�E�nE��U�,u{.�;
���g��22���{��ʋ�v���*y���aa�Z���<pn߫�`�Tu,��wLN�xL�l*���ߟ]�Z��
 /F�ʘ�J��������q��.S�A��Kr�ww�}r+�
+�=~��`���{4"�A�%
���<H�)s����7����}�^D��T��{����{e��R���F{�6f��J�K�5��$�U�n랽���4|�k��D�������q�P�y阨�b�/eEa�A��e�chm�a
�� Q�j/gs+�^,���nq-7c�'֫�]Mپ�����"7��K]���ax4C�mxϝ����g �V6/�Y�xB�%���n1U�7 G��g��l8Jw�,4L�U��	8�&s>�5:�y�隄;+�������8��gf��n���:�r�B�o\��/y�\����8uB�1���Cz�h�	.��K�0p�s�f��������P��� f�a���Y9�r�絛����N-u������TvI�s��Y�F<��fu}%�O��|�콦V�i�dM�Z����f��R��=;wڴ����1MNş�*v�k���q�
~Zѓ�.wZ�7���W�i�]�Q�)�ذ�+P�s8����:d���

'vL���Sc���t�ӪX;F���#�@� ��\M����wv��^���#3N��'���3�g+ü٥��[#5t�r�jyqE)���a��Q�j۩����\&X�dӮoϻ�1EﳫJ�����6
��=b\(PE�[��X����[�{T.)�[��kμ��l�sr�0�_)�|ή1�c�ЎF�����߭�vz���@[��[�k�x�,5a9�FG��Q��+��%��~�J���H<e��ݫ��y��'7������C��q��J���֟v�zH+)@�7Nd�O9����b�<�Xŭ��t�⺇\�)�q�:����:
.�S��@g/#�3|$\c��H>+"�;^T�r��R`�_ctF�9H:�j�hn@��b����V�D��Sp�ԨƩ��F�4�k�5�̮�Α��{��@������q^p��V�&�)�l�Hf�C+.���Բ��Ǎ��2r��͊�vSi��_e�B�WԸ�� e�۾��Oڣ�c�:j#g�^׈�nwݵ
�\)����#.4:'���|����F�\*{�'��}�{���<N-7�,��ϓ���8}�����T�}�n�}-�]��7��h�?9"k�>���
6�nJ�j����Ղ���]��U�&n�tf����3-�
Kh��'U�P�O�E!&�8�fϽBO����@�i���B8����_a-��{�m�	VC�Zl���bӣ�O�d��=X'�\
B�T��;�3xYM��X&6x|}u\�pN���v�����u�؝��P��}-����~��V[�R�e��5>���զ
����B�;�
��b��::0t:�����-���Y����Q��Gg3<���"�r"憙p�%7�.^{��w�N�E�uQ�;uۆ�tս���ݱg�wt�;�>;��#����㔂���Jzf)K.z���X�y�ٌM	9?>� <�=*�seD�X��	
���p����`�1Ƴ^�-+��=v�f\�WG���NQ��f�����3;it�\�3�ORm�Z�V�ٻj̮a�*�2�s.��$�)jK�c���UFu�ܙ(8��-���52�t�WM��"s����ܺ޶PU���3H蹒��6�w�L[QY�83.��<瀠w��_}��bQ'����߼�K��䇽$u�� _��b_LjS��0C�:u���L����if��R�tKiڋ[�t(���b�+t�c���i9pL�`//H@�"��۷�ߡ�t:������7��^�,�ٷ �-��X�~��fW:sQ:�T��yL��z/}��� a��ˎ�h��tS�8v��%ʀi���E�� �s{v�����-g|M�J�\d�>�'��s$q`�~\��-q�|��Wp�p,U�B��w���3��{�ק���n���rX5� x� �SӁ�,��2qf���^�T��geuy�����Uu0�L6t�H�u`3�A����.�䡣���'ѱK�Rbruo������yWe\SBu�g���I����Њ�+`��g�M�<���(ķ�w��P*<8�C���Z�)�<kVm�P>JI��XS3��&��0�
Oz�����6�Xi�z�>�\<�aL��z��x�H�	4wהl�KL�� d j|;zE�/�!K���*��aW��]�ON�qD�8���.��m��JE��Ii�N6�&���$��f̰�������ɔ�uRS2kw"�S��g{a��>B��۬��&�P�
P�g~�=�cۖg[�7�3]3���\ov�c��<�&��pGs}�I���N�;�ޗL�A3b��o��dl�ؗB�ͪ�h��|_P���=�'�Y]�#ܶ���k�:p�l%ݎڪ��ǥ̂`�_F �e��t�9���� ���B�+tU��K���q6q��L�	�kz);7�e�t*^QHV��c/��,�Y�餼[ը�8�[��������<��YW}�׮#Mfb�lod��d'WD�cx3���d)���{�� �n��K����Y]�<�i1�JaSx��!�Yӵ�%*獚M�u��(�u�ma�,:�S�.��s-�!54>�{�m��2����|+zA�˝�9���}m�FV�P���B�	�s<=��E͚���gpz�?Ogl�B^򏖮ܱ	��%tve*K^������y�\u�\�i��$t��`4��U���,mB���NڹJ]hu��`Vo�>:�$p���݁U.�2���wv�%��E��
*�λ,3�f6�q^ܠ�F6��G	�x�L[:���d�X|�Y4RҘ�3>�T��*�q�-W��.d��(�.[x/'<�|-��hB�r�<}ٵ�D���;��^v�Ә�Vf'��N��BA|��۔��{`�:��頉6�wQs�%�z���㉚u�yn�X%U�=��H�eb@e�;�P�G219'/N�v!/�}ّ�����d�;�Ƌ�;�"�݃$w,i���c9`8%]�9�_X���xJ�|�G�s��[˜Ybd�&�\�8nn�������B	��I�)�M�8�����l�u%F4��ۚ�]��񆌬K$�����0a�i
��O�x���r�ܜ�2	X*�5��TN�����J܎�%\4#|�ۼ`�	r7QS#'��Qx�-�O�W�y��-#��5��1GLi��#�F���9R�;&�|�j�hE.��!�.�^=��Ez^�K�+�B�-���=v1=�����8�Gwn�5�H�N} ;����K�;2�^�-�sc׌V�ⓈުY����E�tyw	�w�f�S�o�FҢ;=���'u�WR�|��b��Le����*���\)m� �ݱiܲ1�l�n�H�"+��)���"�ʧ��p�@���4(Y�/0�,�8��l�|nj�;�{��ͦ���_;1�n��벴)j^�%@l���yc��Ȗ��a5ܛr;��%�-��%m�:����-�� b��L�$����4��	�me4�s�z}v+7}��պg�0EU6Y��c���;��%+�g�Cn]���Yב�����D�$eQ�z���N�j���;5�d���UrJ�ɻu/WE����k��eY�Ĥ��2N'mX�lA+����*���m��щ�%T�Ie��mU�GDX���'�V�rAݨoDp��gz�kGα�Rގ��zr����wݔ]Y����(r��2u��:m�ͦ�iJH�o{ol�i���,e�w�z!7�)�7��?��E���YF( ��5T+A(RR�`�����Ҵ��Q%%" �`��0QdA"�E#UQ����dYR**EQE��
(�X�Tb�AU��AV
��,cV,X,QDUET`���b"E ��(,PQT(��H(
))�((��
,��E�F
,i�("E�X��EX�*�D�
EU"ŀ�
J`���E�FEQA �,FH�QR��,D+"�UX�FE�"���TD��,,��U��QdX���J�)F��dR((
�,QH���
�# �$QV*1Q��TB,""���0QV
�*�DU�EUPQE�A`�,PJ�$TQQ
����`��P��#A`�0dU"1E,D�
))��TE"��ŌF��QH1��AU�Ȫ(�ٺ�9*�_s�}��A�=V��m�˪Q���Z�)-i+�����J:54�b�`Y�&��0�o{�+ɱ[Js��������=��<��KL$1U0���(
)l0{�.R�)&���e2m��
Kf�[�L��0�jͲS�L�����:�d겒�3}r{U�γ�{������9j��@���>���Etm�����
E �7��:�I�B��]�V�ah�Mz�(JC3��I�K@QO�IM�@�->B��L߮L2�|�N�^pAg)5�TDD8`lz�l}��Ʋ �w؍�$�2��Ӽ�=��L�_�5p�<��Y�~��i�H���0�a�ZN'�͊A�IL\��ah%!��-��Ii3�-aI�W�`��&<xK��}�M!-�F���������+�ɇL2�h2�z�H��h+w0����ɠߵ����=t}3뇙�Q
aU�×D�:����fĜm&R�׽�N2[l�T/���&1B�a��������W����Uw\;ͼש�Lʤ�ة-��&!��a��l��K�N�{��r�����*�o��aE<��vt�@��~&=s)�N7� �P�
~g��cɚ��yG�1P��@���׽��}���� ��R"L+) ��b�{5*̘�é���fu���)g>�&Y��CH[���C�-�=k u)�^�̽L2Z���q%:z�i\៰^:�}�/�;}ʽ��˟}ε��g̙��<]�)��S-OR�(��2bwRJUI�)8云I�y��n����e��䴂�Q�L!�)s��0�a�ZM}�`4�{RR_���U������l�>�F���@�� d	�����e�f��4{vE�XRc���I�)���V*�����
L∥�d�YԶ���R�e'P)&P�s�l��
f������䴙��CT'�~����z{]��Dy@�:���i>d�o���ô) ��G�a���i5�������a��R
|t�In�uC&(�U>d�*MC50�II����% (��~�\������i��m���� ��mC	�O7���̰�
|�����!L�%8N{7j� ��0$�YH�����0�S��ذ�e �ܝ�C�
E&.�ҙ�O����駣�b}���q�v,%l��2����Y&*�mm��볺�ÛH]K(���MG�HqI�b��+�{6q[�R��n,^��#�SG���!7�GbƑ��y���s#}j.P�[|�ߗ��N�B��[�g=3�Cq7�ɥ�&�@�,ZKe,a������+k������~u �Cl-;U4-)�=�a�u��9T��S���X%!L�&��};�,<��c:�Q�a��i)U&��{�2�L�l��lXc�B�[�k���=�֫5�W�s����xS,:�%�zb�fXu-��]����Z�,�H8�2�řN��9��)<�3�Ԗ��%"�)=ʚ;높R�)�޹�вm�a�.�	O̔�7�{�6�g��~ί��N�u��h�@Qmz�O RM&��qRm��!M���iԶl�Il�&�I���)-�}y`�B�+��2�a�T-w�L�i)�V|{����E�����:��@����0A����2gJ�p��2b{�T�J@S�)��Ө̆*|��O7�٨a��)�&~��4�Y�Ju>���Фï�L	:�������3���}�L}���?}�]x7�!��uY�~���8��]r��:��l)5>��	�m��Pˣ�����C{��aHJO�B�ݧ�-�a���$�/Xa�I��2o�쐦aL�νQeF�v~�1��	ǩ�����#�#���a��JUI��>�O�)&���z��1�!HoՖu2�l�ZON]��0�ZB��ׄ��a�Zu��~���,Y��d�b�L$����6��oȊ�����o���!��Rw��0��)����1�N�Ì��l���2R:��:ɔɬz���m�k����:����Y�0��2�K~���Im��Х�� d �s�_|3�c쿮ԣ�������S�O(%�ת�����3��D�O�RӨ���8�Ջ �;�8{�<�(%0�=p�jy��5/���6�m�����޸�>U������q�7��6��0�
m��P���m�qFd�Ф��,I�e!�TGtC�P몠�u�R�i�g��u�"�+v&��f��P�A�C��T�,�@#o�w|�G�(�
�~�~*n� �%9M�[=/�"��S�l�{p�N�L�5C�Y
a����� ��1ra<��Rb�a��$�f�tì+�B��Pe�L��<��=D�j<>�P��  ��=�un��G*6:�\MU(�N��h�|�D�M�$`��cn�3&�Wy��޷�����hL�R�[�Β~tW��G�Eб\d5��E
9��C�+j�OG�֛Ig)u�Qk+�IJ�ܹӎ�:��ۨ�͓���3���l�9t�.u��z���I�֊�^�Ϲ���AM��~sפ:�B�h׽p�i<��j�sɔ�B��Pv�a ���ŕ��u
e�¾�d�l9���2���3�gY) ��.O&S�����׾�&*��s�t�/��w5&YY�x��2���'�/�YH,�O6��p��S��۸q��ɓ���PKa�P}ۼ�y)ғʩ) ��j�"������A�N2X[�9w�{���y���~��za8åT�g��p�&ل��M�uÞ��6�l��l7��u��C�d1�\�Ijý�:��>;J�m�X�ǯ{W��qڿV���>��L2��-�d�Y0Ͱ����8�R���<79��!���<�s�!�:��8u�\���S<̞͇���S3��̳L8��~�̖�2R���nw��kG���W7�߷[����$�z��Wj���g��d�l�KC��0�S,2W�0���ZCA��ĔřN����Y�O!L�(�H,0�_���I�+2癞�>��rs_s�������i��Bɖ���Y�@�S��Ŋ,�% `;E�ɴ��9�C(}���Wh>�)����r�&R0�:��&����7����)o�L]����2�1O���v�n�=�p � ��}g�T��Y��Ȧ�IM����2�sS2厪aHJuUuS���d��'ͧP�4I�)>d�}�Ϩ�0�
s�\��H,���s&�cG;��[���3~'\�e-���\�Z	<����j�z�̞�Ϊf�a-��}p�4͡l���AL2�{����- ⦧(Xau�0�T�)�S��&
$����ǜ5�o�ٙ����-��z�	�vϽe����۰�4è�@�{xg̔�d�tw�!��
C'�f��L6µR}�\�3�l2̺��I�0���r�%$�1�0���-��s�{�>k?cY���o<�^��ILY��(��y
fk��)���i�P�����a��N���Xm�P4��>=�Qf�)&w�=d�Za�_z��7u&YT���`
??�Y�\ਫ਼�c���Tx��L��+w��Jn�����v�x�Y]�r���늽�������{m�:{���t7�J��:��rKs	7@lE=�7��aw/��[��P� ��{�oV����@�A����Z�/3.љù���U������\��&�8�m&�H~B��2y��)5���2��5�b�Ĥ�6a�T���7vAN����/w8����4g��������2��T�%7�����{0|v��o�>ߵz��KE2Ɇ�	��0�hRav��TB�m��4ɟQ�����2z�P����
uή��e��uP�u�R�w@[0�!l�s���R
e�f��f���ժ�u^��]�����'��}/�fa�Y�ϧ}p�e��)�}�XiE
Ch�NP-'�S��,�Ǭ�!���3,:��4b���JO$�:�Ru
N Rd�Y�,:»@���Ƣ�:k쉫ϻz����<`Tx(�	���0�h�����AL��3|�B�Wjʒ��	�{�e�I-
}5Cʓ
,�t,->�i9��a�XWhY3��Xq� ZSۺ��|�<��3d*�7ӧ�۫����<z��x�Դ�n�a&��ԜO��j�S�����q-0�Y���Xy�O��d�z�'6��;x������hJa��mRR
w[�Wπ��k�r�v���
��e���C)�k�'�P�
Iߨ�a!�����aE<ɶ�}ju
N����Z�!L8��L<d�h�}��d�L���۰�>��Oi]h��u���[�yDDz�xEϽ��8�iP�y��Fsde�Bٙ��0�AJf3ˆShu@�svcꇘZ,�
tg�'(q%>L��bM (���}a�m�ZN��K8ɛŐ��|�����r�S'���J�����E��߬�gY)-�eҪ��RyŒ��l:»F��a�q-�f=sɔ��0�v�!�)�g7�a�ZO!lϪK�ILY���j�HD���0w`���scaV_�ǹ����Z���a�������!L2±B�sۋ�aH��a�JE�d��TE�O%�S&h�IHr�M}R�D)�X|J�0N'��
h;�Rq��#�w���や�}?Mj�9����L��x��,�A����!Ϫ@�S>�.L��II5�Y�R
Z(b�e4��ZA��,�b���ؠ�a!�T�5.�@QO2gu��#�@Df��}���-���f�0�c6����w���Z��ȯ!��YYwS�kgǖ:z�n��A��l���n�7���z�p���ؠ\�0�Z��40ë��#�#q���)�Qp�)����(-V�t��[Uj1�����U�u6C����G�U�@}�}Ԍ�HU�n�yE� C��	��x�d�߮a��NY=tk��)�
�A�f���9���
fXk�,�AfY�/3��Xa���v��hyI�P^j0�Y�>�ճ�z�>�}��}����+���@�RIO��y��P�Ϭ�r��e�7s,�'����ZS0����l�JO3~�̪��
O0׮�e�6�,5�e�
a�a-�vŔ�H,�f�����w�z�ؼx�c��襡�)E�u����-�5��)�1�Y�@�)&������ξ�0�
Oz�����6�Xi�z�>�\<�aL�z��x�H�	>���	it�����>�w[��4�� �0���zŘ�!L2�ctM������M��IH�X�-4���fj�RA���(�z�h%;�ܙJgU%3;��R
u�{a��6��5_w���vS�(���XN�".���Z>�P��ݹ>L�1U0睲eE-�=�)h�hfoS&��!Il�vɞцaL���2gرH)��d겒�3��Oj��B��{_o����=�6}���V/z}��	i�g�՚f�R)��,�'�mCa^�V�ah�Mz�(JC2v��i��S������|��M_�L2�m�3:���8�H�{�i��������h�zb�Ϲ�'URi
O���\2�L�l<Ϲ�3�!L4�%�u�KH,�}�q4�ФR|w�M0�-��f� �.&hS,0��R��BٞԖ�3Z,xL��{V\���A��;���]��)�V��T�p�l)�L>d�Y�5[����Mo���
I��>3뇙�Q
a�]��r�N��|_l�8����R:��C	�Km��B�
H;�=�����x~�ux6g��{�ׅ2ý�ZϳX@�S6�)Ɋ��H)��Q-�!l��y��Ob��>�^4���Q�}��
)�f{vt�@��~��̧Y8ߨ��e×�����[!��_�xt��(��3}����3�JmOTqB�S�.�I�+*�P�LɎ�:�H,�d׬2ΰ�X�ׄ�:�ӈi~�n>�y���9�Xa�Hu�r�^�-u�h�}�׻z���^�<!ڏ��Y<��m���ں��s���+����E�<hP޸�8��c���ܕ�k��%9�@]/��mNLu;���r:�ŕ}$�]u���]�-��M�d"׬�Y ��ޫUy�B��,!����-m�4�ҵ�Ӌ�!g����F���{�{�����q��:�����Xy�����>.�Ì)��;J8�:Ɏ��IJ�:�'�H��<�c�v�SfC\�,<�%�E}f�u0��Y���0�a�ZM{�w�{�x�
���8u�^��ă�����f��ZR��p�g٩-��a���C����O!L-��T,�m�XRd��)n�)u2b�������@�z����=.G�Ƕ�x���[X��/z�gz>/����������ZL��$�i2��`�AM�y�A�Xa�
H=���Xi4�y�ZMwvy2���eXc����t�In�uC3K��2{��ja��ލp�����m�[�(�{ڭk;9�q�ޛd�yRu��0�7jM�y�P�a���]�h�3���<{7j� ��0$�YH�lǨ�B�L�Ň�)���
gR)+;�Ѽ��-��_R��w�L	�txT 8�3YH5P�L��aH��&~�a�u��5˵8���@�3d�)�d������aL�]��5Dy���&�R�L!Y�y)4̶�mO��b��̬�p�m1�G�ǅG�P�y�K@��a������iL>e��Q�0�qR|ke:��0�u��B��Ԗ���)aI�T�}p�JB�e3=��&�a��X~��͟�)M���������t-_�R,��&[C�qL�P)&�GhqRm��!Nf(2Ù�m<��2S4�m�֨�R
[&=X`�B�+��ɤ�z�h};��P4��,z8��N�鼹��L���?8�S_z E��z�E%:a�-5�X�M�g�B�0���yq�Kd�1˲�>m:�L�*|��O7�[0�l��}�H,�%:>���Ф��7�;�7(��~'�z���ܮ������I����������aĴ���:����>��	�m��Pˣ�����CgٵS
@�Rct)-�y��fb����)���L����������,~���?�OG��Y�|B�e�3��p�9�6�}��RR�O&��O�)&��߽�0�(�!�VY���ii9˰Y�KCS�z�SL0�L��4��.�ŘN��M�~���1����ضݙӞ'�*&9���}RFp�v����R�/���8I�X֌�^��j���L�xj��h��b��dI{z�ʂ��p��J��&L�ap���u��K�B�yS��6���j�r*�uv)�=�3�n�43��Z��q=� |�[�5����o�c�Ii:�3��?��Qa��3�`���_f�P�u�g�;fP4������u�
/���é��$��a�Ԝer��s�e��;tL�R��@YĖ��y|�.�f�k��=�w|�W�)��Cݨ�`�B��~�0�ü�Zjf���R��A��0��Ƀ5-:�JxÈ}X�*q������0��L5�\;��d�_��N2m��Y�v��k��7�]h�Sgy��8�0�SL�o�<w�&Xy�6�3T=�)�a�a�M�
Ap]|��'U��J�;���]U��:����[2�!l�
E��ΰ��97�P�A�Cɳ�����3]1�����W���Wη�t�8� dǳ��Jv�d�W��$����nI�)��:��,�0�
mF��}1ra<��R`��a8�I-���a]���Y��3�h,C�ꭘ���0M>��w�?dyG�R��=�Z�AL��d��Hq0��Q���,�y�����)6�3>������
a��Y\�-'P�d�������*���̟c,�% (���^7}�{}��߲�{���:��N��)�7SHo5'�Y�g�a��'/;��Ag�y�GnᴤR
q3��8��
d�_���Ϩ;U�% ZRx�*��Xu�'ȣ�<}�u�-二?uھ�f}���̞/��<4��R{8�L2sw0�u���Rj�e$��d�y����,��,d��C�P(A�ә�,��@�z������
�����dXrv	�nX�AE�ӎ�C9y�{L�K��|,WjOArE�{ذ���<*x<;8�ʄG�b��^��D�R�\)��g�'v�1(�k���:뢩i�����<x��܎.)۳�O_2(�zn<|7C!FrM�ed��a��}�&+R�=hZLёY����e�m;��t��u��H�\z�8�E&`�Cj��*c�w7i��-�W��T~U'':Jݍ�w;$�#�E��<�@h�*�u�nU��c�f��};�Z�Ɠ�+8W�^Ӿ��n8J�ϛ�Ã������W��dԭ�k���x��!@��a���+�8x���\�7n�T8W�wL1��x&���[�SF�R��zͩ�`0�R�@�M�W�T�3�}q2	((���n�r�Aۆ�D��k��s��Y��a�9�e���lM�Y<���{j�/<���["�v8G�ft_�ܥ�%�����3�J���6�j�`PW[Ʋ���f�@������G�����#]�W��ɂpI-�TfM�=�ts���º�Ƽ4S�2(%^Cƚ�����Q�"n1���A����v������\�DJ�]i�����Y�mM1^�_X�g19�(����ȼxBS{T\�ه����Xu���ש:q� �α��4T���f*r/�8"��~��pE�Q��6�:�I�+�8Yᜐ�F1���.ưE��v��CΫ�as�����3�� ��k���[z��{�5���Wk��X���a��!�V6j��B �/zH�	��;d+
ht�C�Bi����o��Ӥ֋B@�=�$�[v����7⏟M�)B�(����Vt�̇҄��ݐ��b��\�;��-fq�Ʉo&=���3��?�����ex؏L������/w.DxZB�)sL���Y�{޿rΓ_�uc���=r��9�N���5���w"�嶘s2�Ɍ_,�o6!������Rl�{�
�˄�Z�� {�oqv�ݡ�>~��°C�$2��g����� ŕǡ���BgfVd�v�=mW�۷��O��>�*@{���<�l�����Q�A����
�dTQ�;�W�>��K\�Y�-e6K��uXgT�1@��Q%T@P9X7.+:ɫ�O
��_�4��t)]'���H:`6�9!\��-�D�4;���|�cE�08�� =w9J�����)z"�z�w���oY�W7�Z����t%�C����0A�-��c��'�2��k)�:�Y}{ڧ������pDoO����iy/�LJs�͟d;�sG$��bL���S|�oxj����$�f���u],��rהa��Zn�nf(c��+��[����q�w�mwc�ږЫ�!�S��$n�#�()q*Oya�P�9k�[{<�J���]���U��Y,��_��y�j��.��{CG1^;�Ǖ���'½>Zr���gR����Aos�[�j彑I�n<Ce^��8��D[;���	�&����k`���n�IѦ����o����1
!�&��jnd��hJ�q���W_l���h3f��xg���.A��5��z<�ҽ�I�8�2_E� ����[�\16�T[��������2�w6��pa��8FI=فOJ�wd�ԥ�"�x{� xp��N�_���n!�l��7��/�'"q����O`g��5�xIS�ɥc*�-$��:ԵF����y,�^p�6����e���N��U�&��a�9]���Ӿ9�3�Һ�
\��A��5�6��g����
�z���2�Z2��u�F>�����k���A�x�1�*�/�����I$[*좧�s�Uc��J�O;Gd�8������6��?7J-�	nl^��ҟ|�1̟��A�?���A[=�F��J'��w
U�*o��
z8΃O���^Η�!}��Vy���aakǌ�$>�OW��uu\r�*��s26�[s��	Mŀ]s~n��>��6���,��T���Kt�[��lok���i�i�G�����'T��p���.��X	���Of�XD�ӄT5b����u:߱@s1�}d�ٯ\������O�
���{<�qw� 2�Ǫ$`�{ъv\u;0�X���<<�F�,"�hڞ�鈦���)�P*XN��
t��Lݻ�B�q���wK_Q����DUꋮ�t.��$C��;���K[X����L���kt7�FUu������8�6����� {�#00;��W3+FZ7Y�՘���GyPʈ�8�l�� ��C�ȟW}��s��Sm��U�Y�
(�3f�\�7%76b"Uڽu/Y�&�ƪ���bӋR��_�c;uϊ���#6n�Eh���ƛ:�x��Q��%�c��l<4�����K�q��]=!��ޠ�[atsl`]�o[x��l�Fq�Pкc�^|��ٲQqh�+�r~r��&,���������z�v�>��֧��������oY�Nhw���s�l��K�#W�F��F��*
z^	T�8�Ǵ웭z��%N>^siw9�f���;w��z.J���V���]�o0Q���<v41t�`��E3|q\�p�[.�:6v6V�F�M�ZM���Ng|ԩ[�si�d疺�Z]���N7�0����i��0$ʲ��vp�'d�,��U���xu��(���q�ꛚ�ow�ӷQ"1ܴo3X(�z��j��S�@��j*xT�7��}O��Lu�-5Z�/P�iՏ,�5s[���]�.�'յ��V��ʹ�:�H94��TV��v��������l���m�F�vr�������Q�U�םw��f�1�R��ŝ��T2�lO�����M@T��-�x�m`�Ҩ�
��7�e��i���I�B�t뫤�%� I��gN4�ʵP1&�u��} ��a��8,ǥ��F��3�ke;�]�3.�l*&�S����yܻ�e��$[˧����D^ohO^��f��c�8s2:���s�Ԟ5�7�0��n�*�ˢ��ϲ���K�5�fJ1�h#r��uv&���6�0#�er�73��V�K�w�NݦOqH_���ff�&���:�	-�=׿d�wK���J׺zM�uP�]b�kW�S�c)�2h�]��8n$d�K�o���������tKE�1�u��8�k�3;p����_	Bu��+sr�
�����\C��ljв`��M�ñkNٗ`�n��VCV����P�u'�`�:;�\��u��쇷R�s�Y��vPYrť�֗}Ѡ��8�&�Ru�u��*�ԣ�{;��9u�S3���ӏSnp'BгnR���ڤ�S���-�"�u-L��q��+��>�����zJg�o@`&<��}��l�u+qrϖ��'j�~�5|դ]�=���cu[��*s��UB��4�w�Be�^�����mSE��g&9&^��-������d08t3L�2M;��D�����r%��ggxu�U���y×�'$�Z���U�7e�U=l@w��m�Hl9}��/7�)��g)Q�4]���Rg��.�"��*�AEEAAb�AUY���PR*��X�cQ�" +TV(
�`�(�F*DQ ]!H#X�X�E��VEE�EPX�#�T
0A��(1dQII)"�U"�"�UQE���`�E��F(�2
*�@Yb"$TdF

��1EX

�(DQ��VE��F**�UE��"�Ub���Ŋ%4�DQB"
#$D"E�Tb ���"�*������DF�UB
�dEUb�����R*ŊH�Db(��(�,X�b*,E(�EE�III �
*��@DUPXE"1Ab��(�*�E��*�����AAUAB,TdF*�� �U�����Ti�IL�(�EAPEb�ȱV
A`(�E���"�����U`���U�Tb���Abȳ����5XwϾ�3O0k��հb��|���+������:�+6���ʸa��!��䪬Q3x�!U�vtL�����Ѷ�]�Ǵ�\�ޙ���CB�4������s�3�'2�4d(Gm�r�O��X>���Qx�����ʡ��J�������0�Б5\`v���#�����1}5�4+�@��e7s�֤
�S�G>]V���`_���&�;N����:�Ԍ���O'7f��Y[ï�eF���ؼ(��\y^qȷ8g���(���eU�r��X\	��uok�t��Ŭ�>��_��H)��Áګ�SW�m�y�RT�uA��)us��V�V]��bZ]��=F��^�(Gu��A�Xg _���#��Q(���Ν8��P�rL�'�7�O�tg�[#<���Yjyq�
S֩e��C8n����&�
��aB����0����Ӧ �6�z�*�&(P�*S����2�šw]Ð�&�t�JaP�{}R:�"�ܶvQ^���PE	���j����������TA�0���������s�G��saNǸ��'N��c��ع�WyK!�43�q���84�	c�o8��� ��<��G;�p;�]�5��2f��W��J�;=���ժ��C9�2M�(��o�i�(���6�gNid�s ����nflO�J�٩��
��kz��/��9��w��K�Gb���^�,�ބ3�{������+淄,��N�&�4�7��K����v��`q�W#VR�B3��f��*�Ej�i��|sW�G�!j�~����8�����΂������ЧX���o`�/��>%�8���h\S
�؃��T�ʱ|�����H�����kF�6�c��]��:��~�
�E�'M�f�߄x�'����3��}�p��e�����0Fr�FU�v�s�C���I�؝��b<\�45���\X����
hq��i��8�EfkII��sկ�����\mȱʦ	Ї:@�M��X�`4Ƕ�BMq��r�X�!"NI�-�|���޼�f�+����zz��Y=a6f�W�x���m�3�xL��eSܒ���+z�0~^��TY(1g������7;)Y�n6F��Alֿ��ܣ�щ:���	PηMh�_���%^C�6՟yi��{�p<C���S¯�����d8g��:�f�=�i��5�^x^ptr}��ab~B������p�%&X�vf�=�;�3�I������� �}��"����&"�0J.Z��lcr�R�K傝�]��κ.�>ij_$:k'$��'M"6��M툉\���S;jof�b(E��X��f�$�u�J��Y�1u,%̢�N���"��#�r-�5c�{������|ﱛ�e|~�	�"^u��	�������9����z���Xy��<�§��QߗNU�b��ǣ�f)K�`�i� ;ھ�*����Weo�p!���P6���z�<-�w��N(�ޭ��i�����B �!�Ii��!�l�aM�pk��/�"�+�����"���aP!̎^i'���-��y��(V�B;=�n=�&C9;��UM����p��������S�:��<^�x͗�>?Dz�Z�.e^������œ8�t�A��Л�t�L�Ш6mq��9��AT�O�b���� �*�;˖���]vz�>���k��2*�r���W̑Ń��sGU�R��Uc&����k��1om(��!�a�~������lS�j�F�^A��� ���c�Y��X���w�����a3�Pm"��p�*�ڪ`��7A@���x��|���+�;z,�
\tn_�n����{��x�!��tl�G)��T��/%�LIN�l�!��r���w�k�$u@N�{0�:���ŭ]jdY�o�f�Ŋ���N�q����L����Nc�ހ륓U��
Osb�ͬ���֪���7�İrr煄Mo7�r�D�`��� �]YE���:�hҎ;K-�.�$����
9ɕA5%�;���W�}���o0.�����4��(?���'KܬEd1v�E�pT�yF�YF��c�⯹�;��/s~}U���mI�*�K�S���f*"�U�."��'���(x@Y|M�}���e���⏐~�V�����˟o�ɏh���/�'<v	��� ����f��tU�kX��iB	��*�x�Nd�F���G"��#�C ߱g+3|�x<ə��we�w(����c�/��,NA��{9;']{` A���y5xcY��u��J�%3`�	�0�c=�i�C���N����<h%z��N7T����P���.����S���E�����<
>w�5�7�%:Y��5
�/U�Ws/_��U'�e�{O�S"�4��\ޕ�`����I$[*좧�sګ�h��_ee���Cj;R*���T�;��a{�b�����|�09���H�2�D�Ź�L=���XP�1���є��{uj]�N9�̨��3}�B����Py�\g�,#�i��5S������Ü�W���'{n�N`N�E�g=��d���ƛ����6\�f�L	�9����έ��tu�۲����q�C1u^�&+�&u���έ��(>�o.CܩSM�W:R�De�{l��%N֋w�yQc}fy
���<<Mr�M�j2/�S���v��	Mł�k�n�|Nе��,���4dB��%6���5�$cUc5$���!�=����.:W3����Z��B;S���r����Z�y�7��4���������77��gx&\\���:5oF�	�A��LEdz��f��B�I���)�S��b{�:A�v3'���*Z���pP&&(]�ۊa���*�5�e������G1^��\]�+a��s�3�'2�5��P*�\S�f8Q<!��v��mv���������j�E���u��<!���j6��n��q���ޝY��\NMWb�u���:>,���!=�nX��}"��T�sY$�;D}��5��b��Cj�u������r����
m�Y�p\�m��<|d�Xˇ�G}F���e%���5�8�Ѿ�����\�2�zi��r��Ác�9h�o��j�S��m=CC�Qm���8��i@��Z��K�l�Iv2k����*�6�G�v��=J�޵ͳ-:GRN����*����W�N)	��4�^¬8�Z�t�jVU&�B��3)�pISz�\����Wgu.�<�=g��y��C]ˈ��x{wY\�>W#�$��쪃��=�a���y�K���6�+<ɰWkg5d�R����l�-�¹��t|%��X{��-�=����n6q|ձ��Fyuܨ�."��qG({rݔ�wwk�־�E�NÅb�Q�p	t6+lr�lW(`Cm���q$��V��_���5�ܹNEFC�Js�c���<��H��K\t�f<Z8�p��1MivwMt:b�4�L$��Fǘ<����Qyl�ҋ����NǸ��b���ܗ�R\Lg>�9�]�X�-�l��	� �T\X;
m�aGG9+�GZ}�x-2Џ{��nԄ��n�R7�]��J�>�{㼳�.04�>w�P�pv��ns�R��Gu�Q�lDJ��;8�����7�}�r=(J�HV�>Q���#��?������H��W�ǎ��\�e�^��P����D�W./���S|ܣ+���N.6��<����kor����+��S���6���u&_cwKe��DM�`�E�aEz�nJ�eY��Sj'h�W{��s��/Ǐ�+��9T�a:�[@�M�:��j����R1�����\�%��Ώ�J����f��7� ��1:w2�5n�vΨ�1����P0fKT�1���y;D�}DQ��އ���޾�c0nq��{�7�:�Rٜ�Y�kwh���9�y�wu(��w�Oa#3k�R����yW�&�p��F��>ȫ�r1pxf�BR��MTǫ��vW{L��@e���&����GUރ2�G���rjr�2P�G�S~��Xa�ʅ�J>���0��u5D�XY�s�Ћ�H�W��6�v���V&��\S��-0T|�C��۫6��ڇ�ҝ�&�|�A羞��C}�i�y�5�+���b/�X��֬�����W��<��A�tKy�����uEK�����	�2�lbh�+_� Fb���x���ӖrP����v���ev��Crl,�Y�J]�[�������]��v�`����T�wZ��9��k�<��}H��"��'*�mZ�R")�Κ�n�(����&�w4똻Y�bS�xrsy�IpŇ������W[���Li�">}6��
�(�ꣳ�/X��שD*��i�6�Y��t�	y
�	_�̩�X<uM����0�WC����ݥA��g%^����r8�F�F�M����
�6����~�@��:Z�RЦj9�=J���<`�m��ꮴt�D�u9,�N�8�Cո~}z�U.�KۊF�.B�l�Noj5�F�܋�`4�b*���.�ns��Wi.�v��R-[:�m���(�2C��3�xļ9o2�oM��J��Y.��c2����xs�ႎ�����?T�]_��C�N���'L�R��P*%L@P�]�Q�+��A^te^���������
���u���T�#=O��g��/�פP��Mz6 �7�}1�q�e[jx�<' 9:\T^*p4Fҥ����(�Pj6�A|��Q��������A5B��[$
��Ɍ�����R{iܴ�DSS��[>�o)nr&�f`4�6��19�%�1��+<�a�^���Y/������|+.U����>ʔ��q[3�t
c����
5~�њycY�����)K���B��ED�V%�.�e�=�1n�K�uQBuy9�We�1aν9���n�c�[ٖ�-I!�o���\Pk�ny��j,��B-�+Bj�M�Ǜ�s||kPpW�9�_?�'�G�5ⷩ��5YZ��7}��5�U��n|�7ڍ��7e��~�!+�k|��G���7��».R����o��V��)��[�[��E�8
�my=eE�E��#:s��a3^�W�Q�ץ^`kVq���B��4�Ck.�h�]o*�E��dtfJfZeq�ͮ�Z�9�q�=�VH��\)r��RN+��j���n�te���Vdٗ�hK��b��}�}�gOii�pJ�Z�G����:��3���0@ݾ�ٕ{���W)p�oKJr���0!�]9��W��j�3B��_�BO���rS������z�y�v,�nW�����7ۈ���Okk�z�ӵz�q�oJ����������e@"��{Xj��6�l�e.{uYH�m
�vR��E��%��^	���h�3��QW��7[UU�:�:����8�u{.�
��̨�=G�[@�+�q$P:T��/�]Wgs,-�Z�����K��t㣺�NL�0ˡ�[���Ϯ���F�@p��0jj �=�n��`B�u1�N�D	9N<a�=�����p�ց
�>�L����'��ż�U}Ny�N���`S���W�&)qE�~����AK�C3�҂�\��X�1BN���sپ�U� s���AM�3e
q(N�`jb�(4m9�@�199�d�_irZ��U��&�N	��ac� ��C�(�7�����'�P�����<�E{'2�=%��a�`�a�T��qK�7��Z�����=79E��S�N�xC��\c�~^��L��¨{&����v�m���A2T ZqI�Ú���V�9����6e���>�WݝY*>���a=��"�c�Z,��QҾ��8;�Gxzi7�nX�y��Wݘ��q���0�Tvx��ɷ�қ���<)��J�T$���������_(<�]��}cb�����;�ܱ�2�GE)����69��!�Dlwf���O�)���8�WT�����9sF��@���\yX�9�[�;��LL�gd|vU����Uco8WT��B�"'Ԧ�e8�����l�_��
{=��8ڏ��W����j�ͭ(I+Y�*r���jZ�b�H^������+����qp;�X{΁����;bx<��AV��!4��Q~�C�v1$Q]~��AC��8�6��yv�I�'��:5�Q��X���8�ǔOJz����p��Q�r]���+Q6'��E8�T�ǅ`��1�vV5}���Lt(�b�-�u�^ ��OT��ȷ6%��^)>�U*1��u����+OIh����mU�Ql���v��[9���!�~
v=��X�)ӹ/l�u(�F%GOv5���8��Q���>����W`�T\Dl(�v�}&�GG96�O�Ýuq�;b�����\p���@<�%����\`h=Q�AT|�7��+�1ƪ<��~�R�#_E��u.��
C�!��K�ֺ�#@���=r���V����ĎP�e1a�z|���iT:���5d���@����.�� ��T�ҽ�՚5�����\��� ��b�F���s����:]��.����_r�k��n
�>W�c�{X��!'��*]�{��嚍-��K°�.��b��s���Qvm����R��Wi�;��P�;�Q��kwz���:B�p�r��
��S��R��Ÿ���fY|���pY�B�-���C�tu�\0MĜ�|x(�i%:}�������c��\�Ӗ1���nj�=�@sS�et��C.�{Y.$2�1���������oM�>��=�E�KH@����\༗��3Z��P���*][�>�z��{���kqqh}��E;j�23AVV(.�5C9�;�3��r�֑p�vuU�+22I�xfַ{�V��3��E:1�;�y\&��o���(���.۩{��n��j�."u�KЇ��W�����b�+�>}ҠY�bK;u��s!Տ�B(�џg'��h��n�g
P������:mJk
��B�(���,S$�]����t�r�& ��)Gk�8���#���gm�=pM2I�P��+�-�i�<�4)��U-r�+���#%f�	�?[�]0*�ޘ8�ҙ�W!��U��%Gk8]��q�ʻ�n��ե}j<KGS5q��r�r����U�g������x��ƃ>hw;��W*������n_mI[� �$t��W/�m[6�U��+X�b<ݮ��L���DQn9�i�Z+3���qv<�����]iVj����'^�ko'��{�S���E��B�&}A߹�2�L��2�G(�ƃ�d͔m�{Y��ܬ'�(���!;,�v���C.S;/�M]n�k$_*Z��u�޻�'��7LΩ�0�QG5�����m�&Vd-�:�̱�u�{����i�|�xw��F��9�>G�^�P�����7��Y�:����jŗ��\�j.��tY۪�nC��E
[�7���I^-�LJ��i��Ռ�9%[��RM��73$��.�WVv�3nv���C�2�f>t:𑷒���f�ǐ.ע�ݩ�k٨�Bt��ً��=�R��g�jb�6�}���)����޺O�Чo��Z����n��,=]l�m�\*�ڮ��3���ьs�.�2:7�J�z�+L&�B�V������E���l���4K�Zy�j�:�gGl��3��c!���0I��ۛ��'��KMow|Kֱ��Y�����U8�W���a;yIa�E#��:z&wh)S�}fȪ4����U8\�fC�v�H78�-����;�fm��u X����a�;=2B-�w�K�ܾWƞ^�٬<�j�܄��Y]�޾�u��'XrH��:���=)܃WPD��t4�Rܸ{�[:��g;Gf0g��5����w�ssLFH���VDF$X(��E��
��E"�`��0QUb�DAUATR���*�H�)XU�*�"���
(,UX�R�+,H���FT��AUSLX��F
�DH���AT����VS%*��(#
#�*,P�0X#Dł��,Q��)JJPQF
 �ł��QQDb��Q�Pc"�((�"",�V0Y*��X)U(T�(EX�PX�PT�
1U��#ERS
��,X%T��"""���)X",PPQIQ`�F�",UPPU���ŊE��d�(S!LJHRH��Qb�"�������F�ADX�TX�,U�1�(,Q7x�3���~>\�֝�]k+L�%����>@ٰ���c4��;mv���N�k�>�зM�uLlg%RgUپ���< %c���nbw�*�&o���s��BTN+aUF�sQ
r��H��滔�7Ț�6�ڬ����j V��1N/�7~'��\��K'M��7�y���1�������9D��';OvJ�E[ܴ���1J�vя07C!ōU&_6b+�,G���45�#��\h�x�8�t@�b�)��v��c��j�f�����v�6�_*����;Sa:��j��/�BS�W]��+ó|9QH?pb� ٳ�R}e��9�v\�Л	VC�Zl�=(�]�[ײ&��J+���+�$�v2dǁ���@Ց:����]>�߼��g��ܣ*����q�w=����{��^�o��O��^(f��X4S>��%^C�6՟yi���C��{�B+�m]�G���b�&'�Aw��l'�668k��9�zapptrfs�A#���Ǫ*;,]�%rU�-�B�7�*^s>.\'#�%�X���PV��Pg ��Ӄ!�9�J��o`R���U����
�C��,��`�����ǈ�b�|%�9��~s0o_�kդ�+|��qy1��U>��_��L�y~���eח�>ُ0F���/�nY��=Ww�~:(�8|	��ҷ�~��WMU��bod��3�r_�Xoz���׸3����{���D݉MH����[���fB���WTop��8Ψ7��@�`��]��o�zD�.���u�1��(7!9V#j��*�T�֛��o;����39����2����J��p@L�"�DI�v�m��<Q��&)B��ڑu;��T��;}�6�`���Vt�̋
G@^���VJ����^<uI���m��qG?:s^*oc�f�+~��"�ٔ�q����t�L�Ш6mq��K�bQ��K���,�U�8��k��jtt�]Xw}�'v}C�&EC��,>��d� _�Vm�Q�Z�5b���m<�kZ�<z!A��p/Us���ͳ�n0:'D_��H�QD��#���N��,�Myn�h\u�v�Tt㣄qU~�`�nB�����C),��^�}d��y`�mxg���,�Դ=Mѳ��s�+p����E1%:�bO:v�z��W��_��ϡ�'-J�Ơ�ă��SW-�E�%U�Â��0�ܪ�I��C�ww�}q/5(8L 婘�vz'^ư�t���3B�,f*!�
\E�GeJ��l��2P��k��
���ʒ�Ixs�R�֯ew����r�w.͉�����m�iu����qNt��a}|X���[r�SM@�cTk�k^�l�&®5�=��_3���_�\%/�`�e��A,�9kv����sG��:����ʲ.�xr%t£kSVOG��a;���+f�(=�b�}p2��O��4s��\笣�2���tZ��z�_<��a3�7C�7�؅�uH.�q��e^���(��أ�Qs�wWIs��Uen:x��R�:w/<k`��#�گ(�T\������C�9W���Y��/�;|��s&.K�u�V��O)�A�����-t�B��@���z�F9���T�Mr����&o5&��.SW������@F��0��Zg���ʁ��Jt�GU��kw*�N���s�Q�1|���p���k�$tm*�*��(W��>�kB���-��97��U�-6��7zNKV9�b�+|UH/k���u�Z1�4�*
	�;>B9vM𥥕7[�=z�j����-H�n����e�x7aA�fT_���o�h�a�q$:�ң6�g��:����V��[��S��H�[/��&Rb��R۬��Ϯ�ͅ��9�B)�Fw|n+�c[t@~~�Rjcu��@����ʃ��Z�N�:)������L�����SJi� 3ԑr^;���{���.T��'��S�^�B�P;�-ԂO�]��s�������H�uӇ"���R��9���fNW�)L�O��9>�������0\q$iU܄�x��]+g���Ap��WB�%��)c�n_9z�L�ޫ4j����LØY���W���:\Qr߼���Z�w<�
��}�L�}z[��:��7J��>}�QT��T���(�ńSF���v)���Wo;�ٵ��V�)r��K�T>�� ��/&b� s馁qv���sQ{+�;��\�GQG]qmgu^� W���
=�i�{�J>�r�cT7�dtxC�ƣ��GɑyF�K�Z�y^����d3��cb�� ^��V��e��*v㣲M󱔪$k��w�Jm�Ƭ���:j��3jK=.����~�$3�E��6�G2��*uT��9
���t��U� M3؄k�)��������}QE�ѕ()�Ta�����j	��7y)�Ɯn7��|�B�g�85I���q�����S\=_Z?��wn�SM�Uޤ�1@��ﱛ�J�����qr�v��$�2�>*$�Dq�6}Br�Dr�q��,�YS[ڶ.�[5�ܕ*=�.{���`7a±L��+�ay�8��001�|-"�����Հ���H\�!C3�ثKЙ��m����?J����n6�Qj��u�w!�^0��ll`�v0mF���"��I��W�Y�	c����3B��y1Y��7�޹�i�5�"W��c��/���t��j2����63,��e�(!���>������y�{&r��	uq$OC��,���:�/ T����u�E��-���}[)��;��\���2���ٸ�t�h�>�
=@�*/�����s�G Xnl)���b�+��i]?S�+�*��^f)�^�{���,��A�%�3����}&ts��͗.�{{�NZP�L&.m.�}xE{��������|�4qq�4�|İ|�+a���R�S�T}�d`���W�g�O�]Y�ޕ�
� �-)����=��Z�԰��ኇ���bc�[�z��uM�_bw�@�
��6�5c}�FTx���qqNݞ�W:�rY�8P�S��Il�K>"�Q�`��������-��E����|/��Z�AUq�m�a�e�Ν�X�`�3�\fu(��,�]E��ʦ&D9#��1��:�m��W��=i%�`�j}}E!'����g���l
�F�)�ќm	Jny5S\᪥g����{n��\[�f�IL��#��c���K=C!�z��nw'`�
qYUd(��zuk���Y46��ܯZ�G&lK�lBk��1�:ӳ�7�Z�\A�˗@սX�P�hT�b�2yq��t]~F����y֣�t�4���ݑꋢ��U���M&1�������Yy�%.�Zw�]�hJ�8g��;�qJ��Bko��7W�k\t�fn�w��F��v'__��V�[S��A��J���r��--%�3��W��³7��:C�ސU��lZ|GGFt:����ϸ:9��b�9���k�`==<m*�������ި�sC��!)��E��^��)�r���*
���Pg#d���r�Ӄ;G5{gyXZ����	�S���8��,�XH�.��-ߓ� <�7��c��y>U;�L�X��r�2A��¯@�r�ц#�0}n��.Br��S�DE9~T�Ќm.N������d#���CkɍJp��0��C�`4����GA�Q���wsY�H��^qR	P�;��G3����vM���ƥ
�CH��
�n G$׋��h�p�UR]'1�l��� ��] �|T;�[�q�gfU�C�j-*4'Ct�O�.A�˅���+Q��kLv��S���b8�v[�n��w}]nO�ɓ�o�\�HR��*�
2�7Gf-b���|׵M�Q�y=!�)�q����T�#<����G;�'�"%�zF�F!.���c^�lk
�krKټf����.
�۱B?d �vb=�}�{�扏�zWh���jd��՚
�6��1]_���m[淔�9x�f�Q�Èq�f��b�b����A����Ium�4?$�>���]8�F�⢧���Jm~�;ݹS�5��'��ϜbϨ 5}2x�W��A�ΆsFzo��P�t�3WlPe0w�C贠ۀ���k����y䋴9(h������&�K�x�DSVb�J{��zi��Wn��Ƴ�~�9&�3jO����{����f��ۣ��p��+#�ť�&
�֛�3�_�7��}��5�:j{CFM<��R�r��Vi�=&-�Y۩k���	�^�$�,8Y�te��w>����p�������zVj�[��נN��\�;n��b�L�&���B^;B� �.�y�G2C��+�l�V-�E��]~}y�6����'�;~��#�:�pW��6�r���E���)�"^u�YI�tu��a��n1VI�tA���K�R*��W
�84�!���]��=1^���ӂ/"Fe³ӂ�����=���=J4�A_��p�1���]�a�N��E���Y�Mrz��\����7��J�]/H��T�z'@B��'�b��Ws
-���a�T?dݬUw��p)��e.�z{Z3}(맻�W+uE�i��:�vF��^�<�u���qח�h�4vy����s�.�Ͳw>��wS���NQ���]����g����o�7����Y�%�W�g]m���;��.�I�WV�;�8�>�D����U�oE�.�0���k�)�U�E��_�R{]��x�ɘ�^��*��#`<���hD��Kz����]�sڅx�C�8�����X�;��⯇c�����D�1�r{�K�~/s-��l9��3�
+Dul(�S�r��r5�7Y[�3���(��Znc4i;�70Y�7�Lb�`�@����ʎ�:�ˇ��E��e�N3E���c�w�J�v��Ћ<=��I�|�>YK�.[��|5}�v��tq��瓱�X|\]�!�+���zTO��X�H�XE�m0dU�E%Q�D)<cYy���V�bԱC�N�	�6^	�����M �.-	�qr��UVb�7*˞ջsn�im��n�4x���nsܴ�xy�W<���Y�CDU{by�5�;����/��c���fҿag�oBu[���6+� !���7x�޾��:��qe]�5�荆�s02)`'!�f0�F�iq�c8�[�o�/���s�f\��\1�
�nFu�|�#���(�� �ʙӦb58j���E��J�݄.kl;����*��q)W�_��ݎ��(��YB�u,X]_��ֺ2(\��"n�7��s�Zf�Q�YH�'U��y�Y6�u>���^�vU��s����^��)�8Sϓv�k�O�sޚk돇-��G�p���{���V��M�o;�Uy?S�����r�)*sdt��8P��׼�	��-?�e�Io�����dv(ˬMB(�$t۫��M.�l�`Iec�H}U>���dO��+>����t~=8��3�(k����P"�����Q�a�Ȭ�Ǭm�r���;��c�(�G�{�@��Q����*("�-�9�-�@���CkϤW#�g�����T�][[�+{2}9V|±��>���ǝ(�;�;Qe��(������{�Xs}��R��#;�����c�So�)��|�%��x�eE���(>��Mʉs�v��n�>3�XU�e�P[s�d>L��"������G3�B5G}Q�E��4*�H�D��K��w���=-�.�S��@g/#�&o���a�|�NF�/yW�G>��ߴ�<�W�:�������˺��g��N�a�2�D�pT�6n��JceD�B9TU�le.+ra��f�[�t��s����`�����p��@�s�^`'v��z�-��ZY�D|�|X��oFuk����+a�"Q#��U;�&�f��G�
����`�O�m7jۗG1���S]B���{̍O�BV�U}�<W�
��|��zn<F�d(�j�2��\,G���:�
��ڨ��<q��N���mpc�¤nK�1��E�A��`ߗr,r���	�Hm�'B4ggF �ʗ��Vܖ����BMx�fϽR}f���S�P�6��7=�q��=��)EmL0�V��Z��AM`:͋��VD�]���{~�9��wo��X�xY.>3�X�n���4��O/��C7Κ�)�۬��u�B��ك���9��(�&B��N�+�П�ў�C�h��آ��#j
�ţhvwZ\/��pӥr���]!�� \��.���ڢ�繟~�	�>��ca5]��@ӱ�\��%z��d��` i��P���P|.B��,��dH�.ưE�	ۏ:�L��21��8���wKv{��!�έ(��h+�ڎ�Ҍ�8����嚁/ɘC=6v�2��la��n�~��q��P��0��C�~�A[��]����#�q�^��������՜!o���q��*�e����ɇ)�(� ߅6r^�����[At�<�J�s9+w�w/��ח;x�������f�|v�9�(��QoH�m�냈���r�k�yVnf5��,DоE�xW1Ϟh���x��m���;5WE���T�␒{�r��5�d�k�(P<XBwS���ޫiS��-��j�lwi�LK��X���	���Y�h"�36�2Lm\_l܃cu9�ښ�%���_FX�o(0'R�7R��^rf��Z�Bc�A4�M�q�W��+%2���8�X��6�����/���LTw�p�oR�L��>�l`��Nx��r�CD�s��]-�4l郃��j�p����3�]aD]��D��sq��S�q'J�A61�k�*�O�C%gsDU�G���A�ֵ���Dņ��
��^���M�d�J�wF��i��u���hP�����͆�m�Ρ�+iS���*$�	;*�(��GN�Є��鲊��Uqv4�Bv�l������ȫ��Aø���tFd�)-�Zna�:����y�oe����-�Wk�`(e1d>��G:fm�`U�w\g�:�bmp�|;7�VN%rYx%�?]�X�.�V3N+�K�op���s*���'6Y���,��x+�hB�6GMK���S�:�ٯ�,0�+�JW�1����l�������,;���ΪX�]�M.�F��x����^=��� �#�a��;f�+y�q�C�9�Ո��W"�*�GEG��rʱV�N�W���8
���.n�f�(Mx���K�ͬk.hֺ��n=�:��}���q��P��˖�ҘEX�pD9�)�u���U�U�瀙�O�2:߄�O6�\;|�Ѫ����-P�pb|��.��T���m:d(�UN�TO�"l�%���Z�_K�*�Ob��M�㈕	�h�f�!c�t�&��%�[�ʻY�t��g�[�Y�%s%"��{1��w]�O;u���U�>��͔V"��\�V�4��9�_V���a�cm��=�#�9���y��&1�<cEi=L�޽�3��tk�Z_r�2Hs��t�>,fQ2�ဃ���Is�֟Q�x�K{3��ќ{3�򩳠�c�VYNIW��1���x���\��u}�=�[i�[p�����l+m�	&���dS���]�<�] y��n�%=�\-������.3��9T���=�M�a��7N��A�eC&���������w�#7EC��c�o�c1�o�3ʞN����u<q��ټ��������Nb�k��b�򛺯3lZTm"��īt�Ŭ����nv �n%�㍪�F��XN�;;�Ns��<��f5Q����=��tp`")F�ݲ��wJ��(��
��T��V�9��`��F�j�v��Q���x�5���*�pMmU�J	�GpU��*�(�J�!�}�ڤu�i���M�����M*RP���A�EX�2*"ň��e4*�U���U��UPb�EUY
JD`���U
��
`�"��H���R�SET���dQb*�*�bŊ�"��$�D
)#��*Ȫ(���Ȋ���E"�X�X�((�,EV�b�@J�B,QEV �QU���X*0TAE"(��b��)QH�
��c`�QUQR)b��� �*������`�X�(�b��1DF*�(� �`�TUTPU���X"�UP� �"1�����QR"�Dc`?I$ A�t^oN�}y�x��svg�N�9�rz�c�>�$jo�=��?t����_9��pk��_%�辸7$�]9j�wL�{���o�ϳ�p���^��V�8�"�(/HHM�݂A<����+O΁{��+j�����y���:ΐb���w����gfU�sPm#t&�t�H�:z�2T$�1,;���ܒ\x���b�w
�l���[����C�gv}a2p��)pb� �TN��N�]�y�Ҵ�{��u/�_�`�7��qw��\:�S�G0Y
���j�Gu�ǻ}v�u�N9�z��^�
���sq�>�)��2��Ǝ��������6uI���Ȳ�
K�sʿ[��C�=8"�65%�^�B���d��WCs�JOe;����~��y�tv^5��`��%�[��!��`9��k}	�A���a���Ed:��Wk퉷=�Qm���&��l\+�Ǳюs���1�[��l�~L�jH�*�_	F/�#9H����մ�-����y<���z[���U�r7d�w+��ٱ��끗�|����tf�uCkf�N���w�GS>���qa�WO�S�/�6����W�;/�Ub�˻�4G���2M����	}�ؼv�:�]:u`�^y!;��{y��tns�<C�:an�&*��(�����ⱂ���o�*�4��u��mC��u����f6����z���ԑ���-��՚9n�4�C�s��x�yNoj�؎�s�u|3�^p��l�3K��>P;n���R������7U-w���"�7��rB".O�}���d�<;�j�~�i��
r�}�i���M4.?������k�s���̆�U�y��ƸO9�A+Ս_���$Wtj^�1^Z�<��"{�wk���n���h���5�up^�^e�)���$tk��iY��?������A�<.�)F1��Z�S��iQ$K��}sJuNq|�{xC.�e�;#M5k�vWZGJ^�����9��Iݸh�Y�TG�s+��Y[}l�"�-W@�+��w��PG:ٕ�3kh�"�jqe�ʮ��u�29i���j_m/2����I���@��۬��.�e��*^��ː�n���H���F
��Y�~kA�� �(��T�Z��L�x���d�f��oj.�BaG4U��dh�j��}8z8=!�m_P�&>���nL����+��[���}QZ����ce�̡���G7D�!.%+���ńSF�����uU�����*\_5uIFރF�+{n�0�@�l��|i��R�rj�Ru�[Z����d�5��}~�����LȢB��y�:�ް�B�ʸc4w�	Ʀ�������;ș�x��=�p.n�N{sv�;�y��c�)�M�ѥ���ӻ܅+��Gt��9�P*_���[(l�f*2�1^�h��8��(�S�Z�e�m+�g����,���nyea@O�V����*�5cЄӃѐ�d��ʖ�¡3���A����5��1�ر��U�#}�V�L��?A��=
�}�x���X}Il�ޭ-Xj�Qg��uɩX'!��\l^�4���nr�"��l��'XiwR�߾~<d
0e���G���>�4+)Ŭ'�g�*PS�5���Yvb*fݥ���0�>wM�ņ�Z�����r��jL@����8�-�yW�\�d<��d<�s�'��|�U��6�:m��^����C�v1$Q���ICUTl��fx�^���\�$���s�\�S~�.T���P"ݷaºeF��K��[|�D�f�P�#0���|��������(3��.�&(Q��-�9�]����rA��5/-��%T^{��vf�3��c���$8��Ҏ�;Qyl�Ҏy�a�P��$��ݺ��[�6soK���Bn�]r-�Y���=Hԫ�V��a�2�s�d&ihZr`ye�GwΜ�������Rݷ^�TZc�4��lLήt�9�u��Lk+�0gv3j�5��=N2�
n��~B�WV*�v�r)��}�JT.Ia�J��>ݸ��ɫ���%����4�H&��ƍ%�����XS<:nIA<ג�\���\�h�[1Hw��"��䧼��'7�B5O����r.h�xօ�3�zA�<�^�9��jy�Pi��L3�����#�c��J�s�V�"�6[����ѽ�K�v�b�^$B���j 6�S��	߉�
���'M�f�ߍy��k&��]+)o��g�l÷��zd���0z7�����An��8D�/3i�8�ٮ��D7S�2���6P��������"�Ճk���`1�2!��GE�jz7q�±c4F]K���c�E! ���gޡ'�]WK5����S����_�p���y{��ϟ{%l�������ZtvI����>���+�Vu�r�����*N
>�[��;dg�w�I�ց����.1s����C�:�x������E1��0�y?�p�
���M��].N��! �1�x��gu��kp�y�i�^�_!U�+����;�k�ڲ��QN��1;,ғ�p-\k2ٓ_;ժh��WY�a�ډ��DV���7�Yf����B��k��/^�V�v�dh�JVmtD�]��Sw�n��ph�Q_*�p!:|Lr�l,[�Y͞@Q���E!��Ț��8��]Aӣ�.� 3�@�BS{T\��|]ӄ�y�614T9v���q��F��=%���7F*<�x$t��C��~|x�{��E�N�{����^H�1"&���\��=>_����5��W�<����("�'*���S���N�ոuz��U�F�� ����H��V}�m�����lH�w��)[���=LޓF�����7��H5��R��Xt�c�=��w��D(rC��`�6�P�3�zU�:��2�x�%6}����rZ�=�[�ru�+���5ZF�M�N$���YW��Z�.	�J�쎕�����w���nv�(V���gv}i��mK�:��	�7U�2�9�W���E�]�C0<}|��Ut��C�r-p�p,j�r�W6�e�E�:�]��8��޾
����>�|�!�'�OE�1�,�|��'g�~�4�vs��ўF�{�x�^��n�=����*�lV�7��b)���Ag+�6�JM���^�P��Β��	��#��)em�+Y��MK�P�d]a�ū��ĂZ�`��O��9T9��m����3�)罚�4��k�Ym�S�qB-�c�D5j���QwvU�i���4�JX��0u�z-�[AY����y&�R�J��.�y�OrH��r�X{�v���&R�(O)�M��a˖�}��Ƨ��X�pxC	:^��}����d���ԙ#�w=�W�+�VNs���!�F�g�L�jO1WRC�Hɡ�X�ǋ�u�y�޽�|��g(v�d�;�a;��H����(��I�}1/�i��ʨ�����t�a�d�>���X�l���0�;B� �eǴ6U��,������qיy�
h>Ǉ�s4�v�z/`����"�yFߵr󸨷<=��^���s����9���t�3��0a�8�A��sa�);2�������=�������϶�1��q�8��(G�b^#H�����x~��/�qi��z�Wj�9��E%\����5{4����^i�ϒ¸pc_X#+З�UF0���C�K��-��m ��s�uM�b�+��A{]�%�f� .X%�|8�m�#��^�^����~"j'�;�����V�y7\�N�]�B�ζeE��8dT�.�]("5en��\�T��ݮ��W�y��Bb��ʡ����8���K��F��F�=���y�*�\�˙�=s�����`XْM�K2o3���"�ݼ&���38q;.'t�&엨j4r��2���F�.�$�v����7�ӻ0�޷�R7�2mb\0U�rpY}�SJ�y�|x!`��T�PO��aE�c��|.BSq`��=8�K#,�yO،\�WK��/C�F�Q��T�S�_�D	��P�Q���\iBxWq�8�z�����A]O�p���_��#D-S١�"H�􆑵}R��qDk���.������笹��}װ�7~"*�o�����5��9�fl�N$�\䊓��:ۘ	�ZK�7��R�/ɢ*�WM`�F)�B�P�3Z�B��F@>�+�M����Om��C�`vѪ�Y5ܽ�*qN9��>�T
��v���0��W<���Y���ζ��E{/��}(G���c�������WAg~�Ϫ���r�&_H]	�C#*�m^���J��s����Bߟ�᱁g�hdU��م�Ō(�3K�.u$a�v�nMn�z�Fd�5��̳�<:E��[B5�!X��a��o�n{�O�v��d"�o�w"-�`�׬�p/ݨ��g!����s8��͑�4D��ɖ�>�r7����ݨ�'�sZ~ǘP���ŗRѷ�g�_�DY������9R��|�)�Ww2����훜��쫚��b��0�V��qc��{]���wx�-6:���B_j��yk�[����p)H%�Jk������Ɖ�u(���z��}�=�s^�,B��I�cl��4\_��흌	"���z��ʇBum�y2')ˇ���/���*b�����R~�e�q��-���m�p�Ҍs��lV�=�I{��;�ˉlR��=CEES�B���p�AQns�c�
=]�u��**#���%׻�.g�o]���|X�uq��`�J�Q��J;��j/=l�҉��wq�4�o�"�t��{�ޱPBt�K����=��Vsa��ƍ��C�����9�;�%Y��(q�ǧc�97l�u�ہ���VR�B�3��y��Lje�vjܔ��Rc��ӛ�gy��tv��nW��Qt�t>��v��F����N`���}D��O�_�������G�b�Q�ַ"�=Ƶ���\+��Fl��.F*\ή&o6�1�W�aʂ(��xj:j�F��x�n�B�S5/x� ����ĵH�v3o	�=~0W���#������hnJ�1�1��uq�#���d���a�}�+�DQ�v.��w�mBøs6<����h67�};�N�esT�-�l�i|�enj�J��R����1��W��(6��VBoY�ے�ڪu��Ɠ'kȣ����c���H][-q�����`�ؾ\nv�?Hh�ЬJ=f���V*PP�k���,k`�*�X� �m��CY�gީ>���G"��pn5u�9պ�(h<ݥ��I�7
<�f`��{���%2.�p�N�w�VD�,�� ��h�Vsͼ,z�-Z{y5�MN���A����l�3������/3|��Ld�f:��y��aAD����WX���o�Y��E�1�� �P����w�:o��ӟW����Q���+�%�x�������*E�S�46!	O{j���ϋ�S��/:���͒D�t]����UQ��>>����?��
�kO���,��g�E)v5�-��.��ZNo]���	d����)���u�׼z����+�ڎ�<k�q�C��>��$��8�(b�-]n�4�����6�ޫ"�>;�w5,ᯌa`!��A�D�]Dr�X�\/7���7���
�|�l&)B��D���Մ�ř�!��s��{���2T�9ó��=!v��t��@��{fԃ��C��~���%�<��f��a{��5�̧��{s�N;���ύ#H�/rU<�z��+��TZ��A�7�d��%Q��kW���OE�^�z_�r���k�?�ym�)u�z)���G��١�#/iib���s�p�¶�������l�@Y� ua��M�kP�5,Öv�ƚL�F1We�L�OvM3Jj�﫬�z��ɦȻ���W�ܗ*�NY�����%�U���5u}'�)�,>vW"F���>��b���|�v��Fp�;�k��I��Ƴ�lO%���j�O��������zl8ŝ��**�.,G⨜��Wm�w�xݮs�1JmH�K@�~��W1B�w͊�!:�*NHV*�2s�R��9"�lfE^��Ų^��Z�,Ox'Q���g���o�1�p(;���N�������4wOKw/a5��Up�ȼ����M�."%c= �L�jH�]I|*L���ه���6���^g*"�U�R�.��+81C�����t�Tx��"�,"����s���]ຣz���ץ����qx�<�;a��>�Lp"��8��?zz�@bi9o����I�tw�ɪ��t֠�t���i|�'�|���ᭂ�$��-הm�Fܹ(���6�&sX�6�clO*Y��Jν�����������Ч(��$�U����8)s�`��k�o����+��M�e�}ٛ��Zw���3ѡ����"��V�"/sqj��� ����DD^B9Vp�12������e*��¹e�T�|a�]۵��rN����ν��;�8�;T����$�b��ӳ%[X��e�i|d;8���_ܬ6��=y|iR��lN�;����ٲW�h�<V�6��7�KQ�&���m%�3���]��A�-�ϖ�мe�M�0z]�ܹ|+���4c�#=�-�g-�nݜ�������C"�;x�|$���/�W❂�QW�,m��n]la&��46m=�������f�L��\��H�,�39��]��f|��@v�ᛆ05U�D��x�$�	J�t��)�<W��ee�gJ�h\��j�F���gm��lи4�Kz�u��O���S�,�w��q���r�%s�-b��%�:q���J}� h�&��u��y{�7]JY�$@���(^�ֹZ�3_u��	�>ѡ�ٿF9��ρ�M�1�R\خxna=���P�� V����(3yg�N���-eq��D�Hu<��3O�-	�)rdf�!^�Rl���ۋ�q�͙@�P�A!�^�RdG빽I��.:�#ئȚ��]C�$��{�zf�Q�$���bp_b[��+ǹc��N!P:7U`�����4�Î�ˣd�8��dYٮ�Ss�=��ۚ�d1$fż�����,΂��|v��˯^عc,�Y������:�}ot�q#a�̋�]�ʁ�J�=�ĳ @�:�j=}�mL�Ks���G�K�ײy{f,e�T㨉ܠu/V�Q�w��y#���1��ٮ�Vi��	�A��?@B'R�G�W�J5�s�H�h0pXݾ�w!��~}��H�LN�G��:�;������0F��vF�М.���uԈ��.��,�!���}v]���f;����pV41�p�i���WYYƘ����dH��m��sZѯB
�k��Q�)�Wkn��3�G�75��e1ص�8���=�ˏ[���a6��5�H�5�Y��F\2�F���f���y��j�a">�̂ �Naf��F�{2���{��%Ն���'<��/Y����XZ[g�lɠʇn�����</o]-��s@'�u�^p�m�8�ɗ�X�t�U1��E����$ٔ�G�brK A踊��)�i�%ν\���q���n����K��T#R�U��}����cڥ�J%d;�C�S�b���C���nf��k ik4�fS6)ýgN����Lں�zspM<�o�ڕ��D�4k��������̍���a�AG� J�t!��]�{}�d�n)�e�w�T��^��0�2�A���N��ř��v���r�N�3G�c���ٸws�6̮�Ve�r���O��&[w�D�`���OvG9���3
��MJͪ|��}�݃�'�O��A$�LV1Qb1H��UAPAY���Tb(�b��AQDUX�F
�����"�`�
�f�A��b�(�DU�*�(���1ETQ�1H�H�DbEQU����Q0UX�������TE�X�UDPTA�Db�Ҫ(�Q�*�Qi��(�(���#,UQTQX�EX��YDc0QEX��
1DU�FQA`�X"Db+QE�
b�PQX����0V(�E�C�q�����3[�}U�<Q8��ݵEA�K.dn�����Ԧf^�A�ͨkz�k�Nϸ�����9��r�a�^��;;�1[7�:��/�漝�v��h��ΜSޕ]�`_���Ժy�����궄nF����ǟkĳ}��v͇%�C����'̀�Z���]/ �J��D�W������S�����;A�����!�tA�D�E�"������
����|��-NKg���uF�5Kq7�v�ķ�����T�H�-ȱj��ux����27�g�����z��xi5y���ʋõ�^��*y�x����|x�:��~���Hw*:�V���枉�m� �⛀�}w�V�0Es�圑7��#$!-�ظ������ʥ�	���FEa�[]
����/1`���ؘ58z�06���u�.J��n����xU�sSk�{L��a��	�`U!�5��6l���N$�+��!���ݍ��s��#Y���=�5q�N��)�����|���@N�	l��c� �W��ys�_�&R�6���(�>��T���̯It
�%�\��0�������λS3>���ԍ���އ����% �G���'E"�ur�t��'}vT�������[��x�0��1G�/�2��+ٽ��1ͻ옅��Vv.)��;�	S���
�]�ӒTt��}����j�tJ���
�w&М�;��M�F�Z�x:.��nR�˯{��j6�c�~^����,��=>ulp;�y1�,Ì��V��яPW\�`^'1I�����8^�Q�fsv}�s�	�oV��fz�dh~H[�ߌ�/���ȷ8�=�;����Pmк�C�J�{3�=�PY��k5g[{��9�q�(F1�T8ڏ������F�_)���5'���ۗf�/��f�H+Vr��U��ݫPM�m��-S��v��$�2�R��ͫ�h�8�ӽ[��������9A"���Jo$�P/dR��@�m��!L�֮rφ����o�w��έ*
N��67���.zT^<xϪt����y|:��~�fևuwY�;��8t��j�
n�˺p�[S��P6$˙
<�y�}��_�u h}�~��6l��uY<eV�
v=�=��ܗ�).&��T���A�,�������f�b�] [�b6�p��|=}�ݳ����p8諑�YJn\���O�����ރ�l�^�䊥��9p�+.m���@��I�+�9ا���w}�natz�5���.4z�7�g-���;ۜ�Io���\���^կ��W���t���z� `$�1��8WQ�����_Q�W^�zZ�ǫOt�Z5��e�i���YY��b�U�WP�OH��th����AEղ:��v&o��1�ǥ	Q=����fWG$�7�{��=�e�|��׈�ntڈM���w��%�`���Lrpb��{;Yܱ���C�8��nϰF|�վ��Y(��<���/�7qh�.�}{��mǝ�p����W�n��W5�x���J���8ˊ�/�X7��܆_J1WUx�����q�k58ɘ?[":KHj�αJ�i�h�&�8�4}�������7r��kS>�m�{7��FV��_���M��c�{:;$����#�zl�O�rW&�3g1�l�)!����o�����N��#r�C���,��g6L�r����(c�'��E\�7�_P:G�	W!��W���0
��;h!
��H*�Y�a>#���SO�[R��j���+�QL*��:[EȰ*r>���K�!)��.^g��;�
N.>Í�ը�+�snv����f����ň�Vg�#������?=;���<&�8�8�m�>�f����j�]��eeXIt{}yW�m�"�(8���s�m(�ެ�Y�b��GՕ]��&q����L������LWO5�*g��oC��W]%I��:�w�b���fJ�G���}"��jA���e���˜�Vy��BE�L>�>��X������D����W�<#xx��X����S׹�턆S���Լ
�Ar^�#h��ȣ㸇qCRዏ0��C�v��
F^=��v+z�TN�~iڅ�C��>�	�P�҉�/Oa��t�̋
G@�/HKY��0�6Va�3��+�P�l�zO�k�]k�ɷ �Wǡ�g�ɝ�V�u�AX��%��8}<���[���O�� 4�l����Q��UzA��e��t�][��v�ݟVTl`��W���o�JN�˳,9pb���!Q#���~]gUZ�,=��\"�g��|t�0����!RK���90����.i�1gh <�Ң��xˊ2�� ��j;�i��U���L)�P:Z;����`�R}����Hv��X��k�K5�Rk�ƫ7���m�{��""X��u�l�!ۚ9&���RZ@�;b�]եG������r*9V�u�K�f�e�7�a��Zn�."'��:�T�1�R��fg�H�u������ՙl�� �˶s��u���T��]T�*��0��Y:�k�'� �]_f��[��T�uq��m��łt\��;�$����w$��s������)H�xj��㭋�[F�fI/S"�q�j�1�]\c{϶_2�j׹Ӈ1h�}�ި�TB3U�^"�I�,61C�ϲ��'t�U��7*�P///�[xw��L��0���|���A���t��;�g�E�Bx�Y� �̀�ʨ�s$������*�,B��o���/�����^��ΫPi�/�܍3{����3�q��=��+��
�e9��``	����3�^ �A��$T����afvA�ˡ��AP���:�N]CYJ^�y=eE�@�\_�sV5a8�RE����b
�o<��|�P��Q;���T�(�-�Jt��b�ӌ/v��L���s�CNC�qV���~{��8���p3���@uL��"O���T�SnC�)B�>*�=��Sº�����c���/u��\[�Ǿc�s'�:B�ϊ��yȰ#-W@���e�7aE�r��+c^<��J������	��l=�b��.$��(�!;U{�\('�հ��ݎӛ	���چ�sô����*�P�6����V:0B�D
�����J�5���"�|��ğ���`���D��h�`�������_2��]Æ֊Bʷ��#�xwDB��xE�����,�[�{�8�Zw��g���0vK�t�n�-�uyۄ��܉K�Y�?�Xܮ���#?��0,wK]u�X��6�j��
΋/��Ю����S:hoq���v3��a2�㭋����u�� �j����"O���8���n9y�W/×��|�V�Y�y��tk�!��t����ߜ�Ǫ6l���TM楠�+,�eg?C�ЧU�P��DQ�4}�\b�����q�P� ��u�G�����\��}/�5_x<>)��Lլo���qʦ� �F�@30L��V�Å��M؋���:���������j4���ߗ�Gg.أ
��έ�����1,{Ni����J�t�k.f��N��7��Q� N	�&�\`��@�*6+ԕiw��q�]d�����k�����qȷ8�=����c�Pw��LJ���<a��`qyg�鶲=��xv,a�#o��s�˅%{��Z����&/$l�!>�40]mWB��X�(b��7�5���x�ݼ�U�m�CT�e�ݝ�j��M�r�ThL�W�,L�F��P�l:��FHb=�Q�Pb\��].�5-�nÅ���:}df��NQM�����o��`N�ߥ{��O)t֠�DV�:��V�q�=4K�;K��z5;%9���|^ߧf䣸ᰟY�M��%Ib�c2t.<Ls��F�R�2�^��͓uc���TZz�ە�PrЂ_G3VL�\��W
.��9�ޱ�2��5�=`ЇN|�1�7��\���ǎ}S��g:��AKGU>�u�x�_GL-��|�T��1<���5O��YŦ��69���Q�T탎����!k�:���_޾8�ﾠܾ����T�r^$DW�����������1�|�I�}��.��������GXO�;�a�Bu�!�>����{�Y�^ĔW�NT��^�gW|�x�kϘ�q�nps�������ؙ��c��$0�4⛺�G	�{�N���d����Ɏ8h6��iK�o�2շ��>̶@���C�V�w��`�/%)a(�+��1%]��yҭwT7�.�o1*ׇ��cZ��4��>
�U鬵'0ns^�%M���>��6R��ǜ�s3��pa0�6��(�5�U�ۚ �;��KJ7Z^���`�}�����ME������ן��w�,�@�'k���ԁ���2�x���V9��K�]�<�{'���3�^�pf�C�rg4��q(�%�E���:�����.I[��`�l0�%x ��C�p=�Y���L�!
r烧j/v�J�'*G#�R���}@%�6���b�{�wU�ȋY�C�.���[�t�y�O` nZ)-8�m^+ڮfm�:T���{�F��=^�eNN� os��*������Co72�pf��J.MS���&-�~��@���[���h��@�[+�{�bs���.mw����6�c�ꜧх��t��AGSQzk�j��F���Cm��k����؟PܯH��fJ�������c�W��=8,~�gt����Ag�W��bm%�L�9E\L��i.�ZC	�)��}Z��|�v��ٴ��;|֙�UnIfi��Vp�<[8�3��{-�z�9'y�myÖzR��՗�k :�AΓyLc�?s��]R�nv�m�H�vٱ�n�M�n4���P�Ź��͝�3@�IPCTk ���75J�[�yK�8���Ƨ��oY@����3�8N�Gס�x�Qwf�+���H�T�"�����=ʺmk4!B����'H��-cǼw;�{7�YI�d�AfXe�6Mf��]F��]���N:G4n���w`���k�̉zr�j�S(|-����\��sמ	�ӁR��������!�
rcvJ�����j��_&=�"@��������$���C]	����k}6�w���=�-n0SE���_(�|�tC�沏���
��Y�����A���14�n�+�j�T���r�ńĀ�n�#����I̼���I:���Rǵ���1v��Z����� Fu�BKP��"5��gz�⛛�a���r���F�5М����\~��[+�)W�Q�پeo�=��en��}TE��!WbU��U�U�vf�	��ʹ�tؾ�1�����|[�v����y���	�W[ފ �����Z�m�!Z���Ѹ�^+}�P���ջ���<�%�]~o��Gm���Y*�V���'�:�����Ʈ�)�m%c���+�{1Ȟx�UeB���/d�WU^{dG��W{ӄR�H����g��w5�7��'�^c3��]*_~�����è< ��Ԡ؃����I$(ּ���#�M�G�L�ov�_>�`���i�����x���(:�Z���{
+��sY���P�R��*P�}�]sV5[V9����jK�مΐ�uo�2��յ���poǸ��1�7%mW�>�3�J��ǴvF��LEs�E�h��W�.+��,]a�a{���v{&�²a˿f���\]o'V^�{����,�Ҡ��{�c�� ��~��Ig��hιrLѭ�4���2vu�tOdK���&�U���4��>���:�]�4�\�	�}-7Eg��Z��U_T�)�:���0�&�ߨl���+TK���A�7ԷFUM<��u4[����ݣgFqWY�5�jzX�-�*a�����t�̭ۉ�ͮ.h���9GX���\-W�1������G�d��E��/qmw;�����,&�ʺN�����|"pc��*��؎�g�A�����Ջ����N�m����/(��U��0pw�Y)����C�]U����Μ%m�ZF�;8y�MnVԘ�Ę�r��/��$��SEvf@\޶tK꾙��\�י�D�L�<̭J�]H2�`�z��Óƞ���(���7����0�����l;�ҍd��V��%�D-���.^t7M�'a��d�b��3,ѧ���j�h��m*��!Uڻ�պjp�T]���7>��(��$��چJ�8�+���-ٸ��n�}݁�Wn�vӼ��[����B�Ŭ�9��RQ6|��wv����5º[)���BdF�7=!��H"�^�2��i�ɜ*����m�(mysVb�:B��V�0,c�9�1Y
�YF������#x���	Ha_���YC��e��t�Q/
]��p�3s��'r(���5�^˻�{���
�0g[�ȡ�6ͷ�vm>+(�K�e�֮��F3����j�w��,��o���~�����e��J����~y&�������^x���k�5�E�z��lfY�Q��*!{D�e��V��S�؇s�W�
χT�j�`�¶�i��,��,2𚡯w�����p�ؖXV�禑�gpe�WF���wX�xzi�3��������\��|�f��yK�Ę(�'��,>�{
��I�nb�����fE�˄�KvIN�ܦֻ�9d���ss�[(� \qiBS�ݡ^�/r�n����3&�
�\.��x9���P�����{��dE���_o�����z�&�,Y.qW���
����<]��ݱ]V��c�q��b:&<�uy7����"����k��b;栽�p[9��5��}Z�9�Z�����(��]\WX�'95s}�>���V�{XD�8 �gD;��L]��Es�����yţ{�k���v��'qWu�DF�df�YO���vmhd�ڮ�ɍi1v䂄Ի3�����WϞ۠+��ε:� w%7��m�Hg>]�;�W��śF��y��"��fĽ��2r
�s���f9��Z����c����i՚�P�Y�q:U�J*ӌ�/It����j��еθe��l��ެs�1v��{��8�6�Sۀ#n�f�Um��{';V�ǂ�ܣ�;31)T����jE�&�u�:�N�1ΏX:ѫ��	�{Ah��yd5c��E���^�/�&f���va]�P���*�¢��s�3;%V.х��W�Ա�ԩ`�)$�P+���"�%�����_k�����!=�Ev�dV�{�q���e��#GfS�+�9(����>e.E.� ��|S?��pM�5s�R�z^���G��-��1�v����?{SZ���j��.�'�n:H��x�"�[�G0\1)���g�pɏv�c�5��-���B{�*BL���p�����ƹ�oP#���`����X+�z]����(��\�h�V���>	�V���$�C�Vh�QAQD(*�*���((�Tb ������"�)�Ub��X����(��EU�B"�0U�b0���"��b�QEX�TU�QP����*�X�AQ*�UPb��"�0�4�$D�Ab�ER)�`��F"%4�������#�������T��,V$V�RER"
1EX�R�RE�����S
AdPP��b�P�$R1��bȪE���*��	UQV@K�)��P�
E �
[�H���c�^�鱽��cY��c9�p�����6��2�d+ͤa����=ρ��G&��H�ℜ��<����fj'� won�i��,���x@�H<�ͽ#Y[x��w49X)m0���u��8�R���+���=�u��H��*�IaOWvk��-����emn�Ď.S�"��Ӕ���T��&��L�-3M��2�TX.a��]�e"cX}�9�t22}�xNRu��a�h5�Ơ|B��7�֦8rw�+�v7ޫ�^5~o6�Q^vБ�BZ+��it�[ȮN�j��j'tr����&9Ag�zx��ߡ�7�F�)�	"%��}n��W�{��^?gר�*�&�~Q�=�f����wNp�+��D��Y����l���k�.�K��'���#@��p�|�C��ꨕ=����+l�l��*[&��msJ�þe�gZgM93`��WLfZd�n���6)�ꑊ�#dU�"g�iV��MSpg���o9��#�����Q�`�����7���;�*�ͩg"e:��l���:��,�6sd=��=���=�d�cm��U��V�G�u3"1@��
�Uс;5������F�)�:�ܶNY9���ܱ\�9��RE�e���ՉMj���=w�C��5(8��u	�αA��궎�e>���F��M���u�T�J�R�H2ؚ�*k�8ь��qW]����UJ+��\����T�oy߹�0S�C����b�� �wyJ(�Ȅ�nF�-���w, _Gׅ��l_�qX��N��fh>Jr��e�T�o#l�,M���A=f���Q��ܚ�j�ϯ^p���ڵ<8VfZ���5,p�b�t�VUx�^#��R��7�o-��{�:Ů+*�S��]��j���³�[nrV���X���r\�6{u���lMRb�pYٚ�O�b�+�E*��}:�+�M�L�|Fu�XbΌI��!�z��	�D<�Y�]�������H���\a��:B���x�<��tk�t���yޯ>�5�����蠇_)�f�B�B�!ѩn��h�坨)q�b�܅��2���c�:��dt����n�zW�rz:�\V;��.D^���gn�}�N�V�c����ƅ�}cH���Va���ө������xNO��7�v�ن�$�Cu�R�Q��B�ڃ�o"�\k��ІE��Qmv.��o�0��=�{�S{N;�+�x���l���	��k!z߇�U	�R=���W��}�'��s��[��ާO5�3T���P~�^��*����7-�M#Av퉛�J�l�`�k��`cX۬�X��J���F5#kl=�K뎒�ioD����H5��'k v�����y���W���t�����s	R�8�r��M�������h�KA�}bH�R�q�ykj�&�z;��_'�VV��N|w��¨�uڱ�)�æ��nk+��=C5-o�9����-ʚ��8J��Q�-�克LH6�P���ܦ2�c�v!;��T��Up�v�
�Wk�l��@��BvJY�C��VW��[�}������-��w�4��Ѯ�9�-�V��h�R�ţ��<iO�Ea뽽u/3�1i'@�xȍ�}2,H�\F�C1�Mrݧ6�`�l����L
��^MI���Xo(�4 �ؔTV��q��{��z�k�*<s&�PFkG���m�ݙ�i�l̛�]�b�D[��Nȧë^}�4�����5ݹ(MQ񜶨w�z�	�!��pw�F�HB��R�N2����_����Ʀ6���t�IN؇n�&�Qv5A���N������xJ"��͍�km˩�^闼�Q��9<�v�+���+�j��L��Իkx7Ѽ-��k��읛������.+��[�Sj�W��IKZ�
Z�]2/h�����S��p��p�@/papA��u�^�k���ڇZꋖ�ëMu��Y�%�ջ�����OE���.�<��l���̡���䄻�ך���~�̎{�sF��.(?)X�]R�����Ѳ��t\�$�/^��~��Ꞷ���;D,�ҥ�P1���ą1���m���k�	�";��jk�V뛝��X��/S1��A��i]w�g���#�������hү˃=~M%�\�J����t��̶)�Z��8j�e�zg9��nb��E,�>�R
�A��B#�!õ����&�
7Y��Ï�o�LnG��VM7�5ٴwF��R�!0����4�7��b��kC̺��&t\+��JR�aE�J��p��#���������Y���S��V(9���n��TS���Ї������{ՎPe�*_XT&���Z�,�=����%�F]J��k�f�(;bCz.O#�u\"H�j�1��̢M�LهB}��g�O?uo��ж8�t��3�Ds���D��	�<|�5����f`�:��A���i����Y�]���Y[~�v�󹠁�P;uٶ���Wskݲ�^���;2�0��}{�X��=[�����<����f���V9C�T{�eh[)�����pӻ��1���n���f&���IR���2xc��.u���2��'�ڋ�q����F3y	����b�Bݭ�4��큛rР%tQis�Q�
�����g\63��S��{���ջ���N�pޡ#���s��јZ%u_5o��>�A3Y[j��ԱwLܮT�V���0m���n]�J0L.����*feL��z=�-��y�7df��K<z�\l��v[���%�Ѽ�Q��z�s�qY��A,w\���6s���_��1p�T7���$'��睭��b۫���(��-q�wf���������G~Q�=�f����]���1=��e�#�pV�*��4�{��|l��X/����]o�#A[O�)A�<T���;�����cσd��{u�igR���53u��ٳ�\+�F��h+��j���l��"g�=��w�o�h���-�Y�=���9Z�U`���J+�gW��:�3�jڌUT�#U�Q����Ъ�梟_���h2���C�oT]:W��B̞]��{���w�*w*r�&9E0Ba�m!:�#��hD���X��wlE�Cr����g+t]]�e��=�ŀ���ʴ���35��Ԯj�t��n�EB'��'0���Y2�ni�R]�؏m\�O.e++��/h��Q�U�J����h�0gT�*�YT[�(Y���s����a�=l���lLR�t�Xŭ�2�+)>�qG�3o],��m"�r�y���J(l��5�������kEoF� �E]~i���qvz��v�k�'�Z��ړ9�%�)�������u��J��4#6�f��]'g<&�+�阙�ռe�{7��]�殅yqy�������-�u����-�2�5�P�j �m_c7T��.�D<���w�͊���zr�kOvn�mB���klu��[Uӻ��N���l<�Anִ��R-�̗&����Qϥb!ɐ+�I��+�ˠ��Mc������L��}�)�n�zB���4Gb�#U�L$��<��4[��.�[�P���ܤ�v+��BL��Z�/Ot��q�%�E����$��:7��n-����h���ʽ#5]B]Tnq�ۤкP3����cC���u*c�Ry�i��3@�T���㈋�s��8����{i���>�\�c�Hu؜�i�@J8gd�u��&��
g�v˾�kF4�JKGp�GhO��>��0�đΦ���UKDogVH�fi�OAjE�Th�Y޵}ʛ�������7��h��[v��(�xMm� ��ч���l�G��r�C��zd���M�O+n�785M�����/����t�43���RK�.-�r�#n�H�,�I�5��:�I����Z'v�f�5�ez.u��qw�߹E4�����e"�f��;eL����e�AQ8�U���]*#����	���#6�Ee���;�g�d���r���|"��2b�/���t����U�Bi-��uE�jqX����q�ڿcٞfl=��]	�$M�-���ۣf]�+A��hkPW��m���s]�Q��Bl��N2��	{*MVz/O*=ϥj���PP[cQo�S�ͼ��	�W_��W�/
P�^��t�"�Bv���i�����]�&�Xm[�i�yڔx�VE�ț K%x��3E�g�V(�#;���K�v��(�5�%�7�Y�{ǩ�y�sq�ݥ��hX��u��r{���a�tk��۔�oR9��丮�����)`\@�u=��������U��#K^
n�����ƻ�.����$Aj蒘x�x�����X����v�;�b�v�mɎ���)oYj�G��/r�d�U�Ƶ�ʇ9 R0�ΙՇ�2��5�dGX�Ȳ�-�k��
ܹ�ۇ�#��g���āށ[7e)]�)�ݦSIsد<�G�4�9qA�,K��^��r��L�ZɽQ�F�&��m���T�0������W�Kڕ��A2�aB̿-��wT��c\ݿ?o�ַ|ҷ\��gXL�>��@��˷j���ms����	P�mC��l�ѥZ��XM��kqB3�s\4�p�/��"��� ��ى�����8Q�e^���cgPQ\\Joi�C^�M�3��h�z3�O,����9��9��r����V�J�z����1!-'��#P��'�Y9��^3T&���5�k��{y/ۍ��!�������U���w/�^r0T��w_��k���ַ1u�X��k���Ƃ���߃oH�V�^י�S�Zܾ��de�����Zq�]R�*�OM�9�{�J���t�k.�C�!���
�|cb�,h"�8��#`�Zz��ƻ�$�cwP��dmo^h��"b��@��Fv'e��6Zٕ�No�wGu�j��oQ#�>����XV(n��.����\�mO��㐤�C�h%ǚsN��Lwiu�;Js��.�#s�W��*�p�^��� g(���Ӎ�G^��p�$'�\�rz��}�l0FO�c��@�֍ʠ��[�Ҧ=�4��u���}��L�}��-�����������Q�G�m�nf���r��a�"3���O�{��5l;��;�z��P���ZqCѝXֺ�����o�?#L��&�����޺>M�v�p��nvV�yc7m��v�/̄Ȫ�J�j#��]Α}�'���4��펗S�T�拘A_u4M��������)�h�n�|Һg�7)vҙ�ٓpw������J����Ԃ����1ԍ��!���Jh�����Бչ��[�����O��a�9��A�y�������o�;{.*�/58��1�޸����!��z�M>
+����UV*��co~
b��j��mN1uK�W�Tm�m��S�U��`cj��p0nS;@�`60��e'����7HL��jm��c�Ø�.ڝ����5�:ُ�f �,z����:�'���]M�͖�s��y$:'�X��%�wǭ��Dk-i�tFa�k�
:٩���I��ݨ�����:�d'V�E���U�bt���S�mDё��mb�ܺ���י�Vp���oiVme���2ge���M�y�����b�]�.��ۇx�[]�9@4�T텛�yf�A@ &�ڷ@����t{���`�=��n���m�E�2��� ��u��'��-��I��2�=z�eM=b��i��ˮ�ӝ�ݥ5��<,I� ʽM����C�.�[kUc��F����:Wq�fm�Q2R����0u5��3:ȝ�-w���9-������͇w�G�ɲV�:������&��>[���IV�ood�X�-�qF���Ѿlns�󃙗i}t���{F�}g:��"��_LW:��Ǯڳv�uƁ��K�Aˎ�źd�1L�̷�Ľ�,��q��k�ý#k/��S������6�H��<@��s+o�4z��7G#�[}v\RQ-:��f}w�E���|+���v�_܉F:6���k\�1�V�[���0�i:�N�~���� �t��T�k��ܐ]`7��	q�ۚ�s	:˦k����vaBL�f;�����*�Z�c��М�'*s2�-5}�ܧ	= =v)�^�W]��.iL�y/��ssk�$i�c/��l.���\{D�5mmu��{�����{�� w�3,�m6+�yp���kx-Oou��w�p3{Ċ�i�;-�N��qj��Cܡ]��Ouwaf�,˧%�����-a�Np����je<��θ���Se��*[�vo�ת�ԙl�>�⬼��"VFx���U�$\�G7�����ő��,L�dC�����IW��'�C`�н��q��vh���c3/VP��p�s�U�3p�t�@��e�}����#�C��'o�2[-D.�<�)�	�9p�S���sxR������t��!��)�X���;U)��s�=�'KYV��+jf��M�}�P�mҩ�y�Fn�.��X8�:���I!_lT�B���CX�;0����.s*�:��2�en71�ř���;-r:
�l;�*���v!9�֝��v㣹ڊ����7iB�;��1i�J�j�YM�y/F*QӲ�m3Y@�3M�T����pf�w�`;��5`���iR�0JZY��/;�5�,�v��NR���o'\qfMh���T֩���V��h:`�z�HQU��."�q�z�*+�n#�w�1���ӥ���A��"��*���x���Vu_)�o��.V�u!1E�ġ�-<͕sQ^mn�,0־�^R�g�m�����:k^�����޹[�q{λ۸�A4ҤY*�PE�Q@�H�(�UE��
5AUT�H�QUDA1
i�$QE�ō% �AAJ@�
aB(�@YL��DZe	AR���Db
,���b�(1�T$U��M$��(�cIH��!)�1U`�"��Y��� RJ��AH��RSS� �,��R��AAb�`�B-$"0)(EDDX���R
��X�VSHE�E �EHRȢ���R��XJ���,
D`")H*���PEQb�)��)	L��XRRUF��JH�U`,P�P2,
eF1� )�`�e2�R�H�|n��_A~2��#��Ӯ�}*��fܕ�__R���c����M���3�t�t�kG�v���*S;u#hť��-���Uv�w�)��æ���n���hD�f�Lev
ks"KjS�W�*��^E��7�ab�qX�ʰ���с���]m�@�lT�/�c�9����XE�{y�/m��%T��]��Wd�SswM�ڢ9\״=��]	�*rp�t�^p������̳5�!jb��Vc���������y���c����Έ�����E�Ɓ�Zд/❎�]�M2!�n瓾�{���d���V&g6�٥���ev�k�r��6��}�[t�;B��\��{B\�Q�K�,o_KkV�T�0��|�i]k���%bZ�byݼ��)l��S�o��Qe
��(HiE��+����E�t��;W�b2�X5����*؍[]nz)yO����:�Q�ϻ-qD�&)A�o2Sk�pRe:��]�'��ֺ	��r�ի�T������uTaQ�vo:j�"�� �������ڴn9}/� �Yz��Dk��)�t��i�Y�<)*2M�qm��cc��M�н�[�"B���Q��]�N�t��؝J�Ww�re�8��+��t2���X�+\W��P��U�-#���̞��5C+X�E��3+J`�wV�YouX|v��3@�J��@Ʋ��0�	�j+IXT������pbLsJ�*�:��L�>��P�P�69ݮV2�a�s�'<_JB`㓜��qV�3ͪ�h2!��>��l֨ZSt]��C�[Bᰲ��c�%���Qu����b�B��ۜ�v5(�P�1;tފ���C]Mn;y@]��ʣ��ݎXX�W����A73�5nh?[�rF��:��\"�p�S�݊����麃��3�LG]]1To�3��\���ց����b;TG;�����NaV+��c\>�{�Զ�r�=�E�}La�H;���6�en��Uw4+(��/��T�9����A���ެY�ќ�s-�õb��ޮ�gkx=��#S�DmM6C����M؅U����h�f�W��n^9��>$�4Z˴�9�LV4��������י�/x�|]�����Dw�m�z=��Ξ�~��9�ùn�9�=^ �L�.����P�^��c´�|���Tɗ)�ޘ�5:��v�g_sg�vlp�8!V}*�NR뮤nv�C���\�6��O�<��4_�z��5C���mQ��s�%�#9H;�g��M!���������O9f5;[����o��5S���vԌ^С+����7[SOU^�WVtn��ԛ@��=�5nὧaOE!ʤ`\j�%=�P����*8������c�YD�<�Ds���]�4�K��V���ͼ�@���n�Y�۪����l�B}�W[��n�7��>;E.ܯ{���!��Ke�<o_z���<?N2a�#�kv9�u`�e�_ZgD%�}	�W5�]j;�o_��<�0�����O�"1��J��3֚>37��37f�m����GͳF�qHj��R��h�Dn�W>
b�;�+���oS��X�A�6&�������	��:�^���G3�J7gb�}N�j�P/��(���M��;m=�ݿy�8�/�μٖ������b��MFa���v��8pG��mv�4�S.�슕_m[urNc{�Y���vܖIWE��J�{k\<��h�<�S�Q�zz�U��[G� �4�:��Z���0Ba.yU��5��*�ኽ9���!�5];*���6�N��e��|]^S�m��p�VU���9�ן������t2[��+�U�.mc՝w�e<�҂��.�{��V��y�P���v�c|{����z�^&�]bm�98}r�� ��b�`�nQ��o��բl��T��f6������+���������Wr���ę��X��շ�s�T���vf�4�[ފ �oC�V�E��)v�%���g��SvtTc1�VÚOX���ȇ��!wW6���#T�[s����M�}���X����tڰ6J�������V���P���wrS�{c+�3��:�d~kB݊-�;�h�?w& o�8��tBlӓq�²��:���8��l7쐰>>�U�J(���o����T��=��b�9ś�R�M����u˯/Ip�4OW�����R�Qp$�AԚ�Y��<��
����-^%Sj���}X&�测�v�����}^[�`���5&q�X5[y4qr7�m�4M	;����e^����;�*H:!K2������T�6�d������ztI:�2��j�i�y��	��X�Ɏ�{o[���;��9�-H4���K��Y��[I���X�H(�����
'"��k�%��Α���%�ǹ
�~���Z��2ջ�:�G7"p����οPo%H��,�m����@찓Dw.ƨ�ͪ�H2ؚ�*h>
+��$��z&�K���.���'�{Ӏ�U����	�@6�;k(�<�dA��\NԇH�hnW��z�^W��eQ��克M�:룮�fD0�1a��-��L4�b*�U9�][���齿f�/J�2��pG]�G6N����������{Ty������q�K=YT[˔-mL\AstU��=˯����������v�����e��q�9)v�LUݪ)��u�8_b�Ԛ����������xXu�iHA٫ǬZC}gk�"-Y�ȯizj��,��A�̢E�`Ӹ�wR�[�E�Ә(��xh)֘!Anrw�6��fY#��:��šxҺ*�}-���]���nU�;���Bzb��u8v��V�� Q��ج�M��mI2��Hh���v�-�/�^����;���ː���Z�~e�!�b����I*�}J�lҶ��â/��c�� �.�Ciwyt^��Z��G<�U��P�;ӆ#Zښ{�$�k;�m	6������v�ƫj�0��℞�}Qo�J��m�~m[�C{N��h`]2�(�6{-q��I��y��{Lv�k��E���{��#J����P1,���.2wm�&�i]TutoE��n2��]�XZWL�����ic��J���1�3����583�+_Z�o��"q�S�iZ��h�볬Έ+�Cp�z�9�6�����[y��4�g�o}�8�\��h�%����F�}k�b��x�XN��J~~
(1�'1Ⱥnx*��]����LS�wv:�1���-��tA�沈HT�A��S[�����eQ��AӲiݑf�n��ۃ)�'dĎ�մ�c*�s9�uiT��B���36媀��y/��Eі����2�[��c,�*�8���;Y{ۺ$���de󡸛�q�.y��ѥWI����hW�D�k�g��rN�� ����%-;�un2�v�f�O��R�����\����\1T�7uyD��Go6eAgыY��uo�핿>���G��VUs2��CF��U3y���/�O;�C9��%�%-+�W���m�������ٜ@��+���I54�<��Dt�-�98�"���E����5�����v�Ls�Lj=7��d�`��r��
�F�k���FMr�6�ئ��
�&Gj�Wٷ%����$o�����큎�);�;�:i\m.]bH��<7�����֦ jc_5cr�J��$`�Щ]J�����(:q�]�c�ΫmZv9��=���|7��)蠇*0.>�a��f+��X�˪�����JI������*�U����=��S�������RC�[��u�\�UћV=dv��ew:���oq[㴱U^=`�F�����%9eN/Q��H�$��V�\�8ۢ1�$ם�щ������u*��%����U�6�
&wؖk�N�z�*�٨�^�qi�ŝZ؍��f/�,�A��oн�#�bh�l�7:4�V�<����,�lǪ�Wd#�u�[��R�g7��`���8�z��kw�i]X/���7�Ĉ��9;�.���k{ �j���Uq��ѥX�=�o"�G3n�T�1�*��P��+VՊ<٢)�5T�g�~�{������������ʪ��S�LSh=sbkX���8j�5����f6�9St[���@�c��>�)���	���W[�B�p��i�.7kX������r�:�@]�Z�[xP=�ش�V2��&v�����3�8�5�o��:��Z��Ӟ�4�A^v~m���}�쨅=,����e+�@�U0��9CuM��'o�Ha�r��F�\�0Rnr�q��8�s<3�[��O��,>a[����Kѻ
��޸dsV�J����x����������P�p�Br�"u� @k<�jt{1i��i^癸o]��͵˩�w�І��_D��nZu�����x	�%�F���dHd���ĸ{<<�RF�Q�#ܞ��"�@��J��뱕��4��[�k�:��vD���%�Ru�3��]�3tC%ԌHkz�p't�;p8��#���qwwc�]�cf��`���yڰB�P#��c�rֻs��\*s9��u,DB0����I�)jئ�gx6�ߡ�Ұ����@�pٛ�pa��vRp0�H!P���<���l���0�ߔq{�N���Lj��.��)$��)=���`K*�	J(��;-�Ws�}��l��a_I��Uwַr-���*�����ʽ#5]^���Z;o[���n�����ŉx�5ԩ��ˬδ����h)j�$cF�O��cF'�w�񮋓���1�:�ţ���ZZ�s���D�n�:�}�Ȅ_�Ω��Z�3���7��u�����g,�RG�qZ�^�h�:A���	W�4����:s�e�É��~��W��)	���5�}:��M��t�ǆ,�S���z�N�0\�F�og._��AQ6�W�.�eQ��兄�e��fŵ��or�YQU��t�V)��͌��7�}��Ɇ��sX�o���2@}���g�"osO�}Nf
Q@Q:�v[��K
�o�Ǌt�h�ْ�k�o)[t"���)wl�S�݃�c��`�(L׼Uj��4�J��C;C�|㗂r���E�j�l�h�@��*�c��*�[���]7��҄�cN�n�y��'FW2�*�A��#��{Ty�և��]9�]eQo:���{y��zlV�H���R�#ڝ+�gj���hV
Q���[�1;���}�����������v����0�q;��*���Z���w����*��S>�}r���N��vl<�An��\��޷���Skn� cX*���c��|2�P���*�x�Y���X�t=N����y����#�Ҋ-";
�cU�K*���㬗n�*c*7yD	篧�޵b�v������t˹J(�f��]c��FR%��f�i{	��,F��.(?r���c�邜Gb���n�G%S����i][�d�S��Ռ� RT;��>�O��\��E�F&���Y:F�"J�W�W��D)'�)x+�<��rƢ����S%Ö\WDǆ��y����Q�plot^�k��5�r�Û},��ul
��0�q^�*�#84�80ֵQ�|_�m��S�𣺹���1R��3C�ɳ�6	ͷ�:�-Z��ɂm�s�3cG��'�L��۹Pm��Rz���9\8�vtN3}K��o�bcvĖf���j���^����)�m�:e��eus�+b�6�0[�`���ĸ:�;dr�GJZ��N�i�󛢛��c@��)9�������v�Z���7�ɢ���)��`�h���ރ#v��k#�{7.v@jkj�YdN�mf�iU��ݹ8󗵂W0L�YL&:X[c/4ӓS�V�<�F��P>夾�J�I\��,��c������t&�>.��6�w��o��7�m�H��U�YN�����c*m�ir�eZ<(�e���w[{�K}W�NJ�*cX�$�[g��ҿA��@�*��Af�Go�:��-D�@�+AKs\:��Φ#-�X��
࿴Z	%*wh��_��I��p��
��.�*�k1k*34>��WcP�&x�a:���Z�l����p����:��^p�f�aC$���f*M�t�A��/�:��^�YMR�˪%�S���� 0&ɸ;}d�̖-�a�9�zY�7N��ݤ#:�ͼB�ԣ��	����A��L��f�;��1�4Y����t�9q�Qfup�҆�j��r�G���йE#��p�.���!*�+a�}]�wٸ9�|��/-��ܲs</��lB=G����tұ�DV]Tq���己��{]/��*߻H����� \���bc[�x'C7s%�[K�ա`/��d�O^o�}�YRg2!�۾��z�l�_j1Sa�WdV����ܒe�$�Ԡ���`���@u
��8�}��o�}��k�]�z庵-��#7�;8�@��-�7zt��)-�����'IA�V�9gK%����4����FvvR�%�=�Cګ�ߥ�MrT�Vl��j۔���M|/�[�;��Y�̬}�oJ�l�K��{�>���̳-�r�ëw�;!��@&�G@�>wt蹶��޳�X�jmWt�>&i��WҺ7�������#nV�g�L�5.�9�d�PUe4���	����!�L�V|s&�q�)��;[X��r��y�V����mMWL��h,�Wq��.�K�մ1����o�=+��;����jU�o�}������͒�±_5g%c{k�nZz�c�}��5�vv���,�k71���-�j�ð�gb�}6ob7,얆<[r�d�q+:��I���N�52��d|�[����A#FJ���[�#u�����'�9= �`��oT��Y�R0���ݤ�E��4�e"�,�P�PƘR*�A`�E��R�����PE��`�U�����FT
)DE�
�0��M2��)�@X@Y$R��)�H�(� ���Qi
dR!*� UQI

H�,���B�SB���4ԕTE�1B�b�TZHR
E��H"Dd�R(����P���`���B�"���RS!M*E�����#)�b��S	LXU!L%$)��Œ�HR*Ņ0�R�S�
I)��)
d�"�!BBE�HT�4�_A��7ғ����K�r�`G�$��b���'���˶٥�5F��&�����/)�Ck�XW)+���ip�Hj��l��|!�>���J�*��g'X7֜	]���5S�f;U�ԭ�ЂO�3:N9�q����_�z�h�-���۟V`�L5�)�b0�X�� ���SY��anl�Tw]����n�K�ѷY���m�B��hb�������h2P���+�jkŕ]�O�whNs��;%�Z���WH0��kE�*��@�yp���1�yڸ�y��8h��׽[��O�MQ�(�hKH�{j�#�G��>��[:a(	�o/�J.�(��+��x��KJ�W(i���Y[����w*��l0�&���{�FH��:�WYTO�H-�j-�j.�oV�w�ُn�$n���j��qsu�sPE]�Br����;E�\��m�3)wFVɥJx�n�����1;w<�T�=��R1�� D�Q��-#���Q�^��1,~����V���լ�Z�{���VK�ptw�I/��� Wc[8З��\c2������L��I[�L���
�܎u�8v^�~ ����*a�{���(L���l�ա�s�PK�L��Z�9��6{Y��K/6I���5|��Ѻ�~���H	k]�}��9(�;k�0mKB�tD����2^��k�(��rW�ڱ�>{��5l7��l$9@��N��3P+<���aw[���v[�`�}I���q�޺)�L8���|��;k�/��T9:��H����<
�u`���� ��Vu�Dn���j%)�w)Svs(<}@?r�HčVׄ�$z��[摤_1Y�2��N�&�����:�2�΂-��((CH��:|q# gF�F���nB�UdWZNj�y�XޢD�nÚ�G�5(8CMf)�4�Yֻw`ԧ��r��kQK����>�6*�A�6&��SO�'��[�/��L�Q��8�5��&������D��ip�<�V�3�\"�/�س/e�ۘ.�pi�#�ά�yB�a�]qlw�qC�:�y�pR�w�)kʘq�Gj����1h����|=�7�K����+P�f1�f����lrp���q5¯�����+��f�^��]s�n�Iy��D宖a���G���V�3�A�)�]\�����D�#̢���{���˪�c�L���םI�q���X�"�Ǟ���X���oo٥y�]���
	��(캎����},�3wKNU>W44���zm�b��ž>�C�A)4�b�W���%(5n#7��WJ�|�wk;U���y�0R�	�n�)\n�Q�|��*��51�X�Qnk�j����q4�[ފ��r��S�9=`���.�k�{Tv;����w�`���"v,����Q���5�W{��a͆�o���-����E�"�5cd�]��<Bj�}��Y�6:��`����h�vԌBP�4��揻�hߋ���	o�;F7�Q�����E�����4��F�Þ��V���	J(�Ge�6
�t䞅��s�a���s}��{�G��Cn)��zF$EWCt;WV#+F�ѭ]Ev�fV�������Y�a3�V3@��QHj�#4:��ϋz��Wyo��}u�MMQ/�cDfY�BV�gTN����t�\m���E]n�v[��iyy
�D�#�[X�����C�}w� ��;�b�K���+��z=rnh�tS�t��[�c89�>�sj��t��WL������wOe���/5�M���˹ڦ���a��ȄZ��S���;u�9�{��q� 듉�p�D���.�d9�:���3(�l��-NL&�m0��5��U�[s@�T@�v�S	�����5�mЫ�����ԥ�N�7������[v*�v��*��v9a`��h@k���-���D�����=��v����'�8c�9�X�t��.���̜� �z�.�u_;5A��ܖb�ʴVd��2�*ۧ�'8}M��9�)�7�R�5����Os��{HL���}T|-�Yx)K��G/U8Y�H,�ۖ��j��1���cQn�QwM2!�n�w��;4�օ7)�)N3/+��V��	�}uԍ��.�V#i=h��dy؛軅X���x�{�qﳸ� �a������n�>�P'm�<�ԃ���<�o�m��V�*����7���_���hyP�&R���2*�3r�e�á1]�㾪�VI����v����&�6��d�i����o����*�3�E�z�@�v�L9����:mX9'L�MF��.��G�x�p�[Z��դtQ^˯��8ljv������_��<%�۞��hO	iE�#��,�\w@˘�[���Vz��oN���\7��)����R�u�P��z.�&���w׋����zͻ�f�H���!�]�Ӯ\`w��ڹYn'uKT8�|��ݬKd�o��� -+�޲�O�+V3@���4)]Q4��2�s7����z�����V���!�g'X5��0�N��Ei����,(�3jFc4��k��d��X\��Ovi�w{/V���V˝#Ta�&h�ׂk1X��[�
���/g̔�\fþ�/T�N6%c�)�-����M4C|�5�XV�{���	j��x1�[�����|�a1"֋����\"x��>[�uT�\��kY5����̹�[xX�(r�^�{j��>�r�F�a�9E�+f���vNIz:?zMJeXa<�.��4�Pe�L���-�|� r˺���X�9cog-����Z�b
짽�	nZ7�G�pK���nh����k-5�_V��ѱ�p7��G��J_u�����²gW*�c�W1X�ﰋ�0�4��.�zF��s�襁�مv�\F�g�Ż5<+XR�t�VQo���5�v��SZ���ˎ�&�]-;�m����i�օح������8nϭ=�t��8z6��N.bkS�4�<��I*V����1�� D��{4�S��8�/#y�U�C��k��W�k]�mm�����$`����uJ6wu�j���.Ze$��ms����M[�oi�S�@!��ӧw`��Kƴ ��uN�P-#�k����_�K��p{�G�6i���Tc0�w�H�'�P��z�����}�o�.�I�qOuA�}���*�Fm���0�2���h4�?s���؜D�C��5�}ơ^���7��uutڨ�m�.��gA��A��5`���qU���)Z���i�ɹY*�
���v]�4�Fmo2	��!�D롚��D�%��Xi��7�\syP�]���mȭ��v�.���xǘ�tHg���s/��d�z����vهM���e���!�ZF���`9*u�t~�S�â�����k�Q���^V�a���&Z�`9�G6jPp�.���+�ou����V+��1�OVp���eި��ئ�n��My�G��j����W�����7����έн�;N�ݥ��(�
bB\.O#�}�TܛQ�pY�j��o��P�H)<2��oX�ʻXm�F�}�m��n+�J������b��(Y��]Z`��0��6"�:�U���k�olf��a{j-@��d(�Hc<5�iN�5vE�\^d����`�Bm�~���B�l�n�U�ŕ���܄����5�'��Yڮ�i	v^��o��Vo��y;iZ�ܧuc]'y(��!�ri;m->����M*W��A�)�L�������፨��	����i^�'`k��a�Z�]��ڎ�Vf���mc]��k�S>�b���-#t�إܺ{���WvN�:��5�����*�����@�ۄV^$�;RP|F�i�t3����>E�͸J�5�Cx솠����^�!�����'+O^��sT�ND(��w�&���SJ�)`߮��,��sI�E����Έ	��� �/[�����!�&v^s�w�9}B�<���k}�[F�.���a(��D�Yq�U����ϳnO�5t��MF��B�ݹ���{8���lF����z��ˣ�u���w]J�=����{�Eb4q�~�BF$EWP���e�����c��o%���5��������3�&v�X�H(CThVq�ۉپ"�ٺ.�e�Z/���=�K]��>��j�ë�܊�[���n�J�����̩�^Y��1�s^8�Ê�QO�͢] �T��-=�Y�F"�gv�K�|��Nc�W�-��t�#�۱�)����3�p�]ћ�o��v<f�<��Q	
���	�n��ʻXm�W�ܼW�����G��kPr����3�I�V�_�1��~�t.�GE����q҆�{��~�P"��I^�G��{�Wz+���`�ܜ�Jm�0i?f��	��5�!+��E��k�A��Y������G9�}an��Y&ۛ��{.bI��Eɲ����q�ݽ�(%
l�{�J����7]yi��|��9:F��-�++��\rU�5q�rv��A��	�����s��^gԸf��b�C�v��f�D���wt_,��J�o�A}�X����;^L�͐���gb�
���'h���[�Xqf��E*�R����Ld��E��Fܼ�*-�)�2�`bu}'�m��u�A�2��\N<�L���"��	����
�J=�4�+����˥�&����5Qs�ל�(z�Wyl=RGrԽ�^��尠�Q��%F�qI�&�}D��:,چxW;1��Iϻ;g\�0���oJ��_X#*��4�It��@��F�
+,�`���Σw��Xj�Ⱦb�'ԪG��jpKg�u����h�3�.N�s�ޙ�W>�kQ��))�1,�R,F[�����i����̨{�fx-�b��9.$�����&��RVxוɣsǺWu�������8�ݎӝ!)��t5�s��zek���a�n��ۑ�¥����z7��S��r�x�ʃ��Z��L�x�D\(.����uG!6*�&��U�����@�àPhxCHڽ��b�_�߼������'Ե�)��]�+���X"�~D^�;U�����xO�uf�Z^xi�~��s9�gv%�C�EXyb�v��n��6�׽�#V��W9W+��6}������W�pQ.�,�/�@�n�2�(��7s��:�i&���o`��9��6��_�Z�b�	D�z�6l͂�8���O����L	�@�''�x{�{����ɾ���W\`�~���f#[�-z�	l�3����	�T��=y���N'erq�s�9Vwrz_i�U�[����¹�4����0Zk���u����=��O��:�5��0��"��#zK�92ԋ�*v�c��M�v2���l���	�p�7q�����6���d�r�.6/
m��W���mV���t��F��_���o.���>�)�����ӋU^���豒���F�������)�ײl�x�4�Q��s�j�8���l�I��������S\=V���;�#�wp��,����F�%S��)���.�l�`Ieg�E�G���NPB��V�W9�2�����W�F�z��Z���X��sרn۰�]2�\��^W���O�=:g�`cl}R�`��-�3=����|���8eM�������}g5�����`�+5��|�q�B���HH@�i$$ I?�B����	'�$$ I?`$�	'��$�����$��$�	'��$��	!I�$ I;$$ I*HH@�jI	O�	!I��$ I?P$�	'���$���$��HH@�}$$ I?��d�Mf�T�f�A@��̟\�+�<*E��
U@(��PPE � �
	  J�JE@P� �R!TP�RI %D�Q!*EU��*��U-�@	
��(%�2���	
�"����@P�UH�P}{��J��$J�*��*�*�UDB)A$�RDU	
��J��@���U	UUD���
HB ��(���(��  n�+[Y۹[�[k-u�`:�;[��)&�QU��qNs�wf�]��J�ڤ���㶣]ڲ�:�ښ��;'rֵ��k����[kUm��wcYUR �ҔQ"T�  s��[m����v��N��[[P�j����f�)���wjڄ1�62�.�º����ۥ,ܡ�w*��v�:۱��;�B�U�1�V�u�7 P�AD�J�A#�  ���ض�8v����mv�U�v���ʗ�[n�v�c�v�]�v��ulcYV�Q՗u��.��-��(t С�СBí(P�
(w�P�Р P�!�EU%(�!QQIQ�  ��(hhP�
 s��P�B� Pr;�
(t4(h8w
 v�a�.�[vft۷u.P݌lS��6�ݣ����\���:�2��	U!(ERU@�ڄ��  \{�(*�0l0�w)UB�a�4W*ju�A�0UM�ʠU�û*�.��EB�,��6�U9UUR���I*�R��  k��Ɓ[(ƃT�Ѯ�%�1T�	]jk0�*���`�wcZ��� �Ê�`��v�(��V����*"��Q�  =���UOUʜ
 �r�4Vh�Z�N�����\�e�+��c��ݺ���U�w4ʷTV۶�Ҹs\m��C9��U(J�(
HQ�  3q����S�V*�X]�wl�MWv�CNv��ͥ����5��n�Mb7wn�m�s[�ci�΍;��wun���mv�܌�N�4UU(���(��G�  �x����ݳ��r��N���ݬ�ܢ�J�n��Z��M�J��wb�Z�s�T��;���#��]�Z�hwwKZ�*��6���]6��7gZ�V��
��P���Q� S��[]�U���T9q.ݚ�4�c��:��55�tu���T��7v�7h�ڻ]ֶ�r�sZ�n�����77q]v0�S�Tm�n����RR� 4 E=��)ICH ���A��  E?�   j��L�U&� �I6U*h �C�R0�Ь�nG%�2���ō�RCUk�����_��~޿;g���o����$��%�XB�r�HH|	!I�$�	'��$ I@$$?��t���iT@G�C��`{��.[
��j��o	���u�.�Ք~Gfp�w��DjUj�N��i���iR�g�vg)��yX���헭iov��z.�0~�m��Um�k{Ub�ݭ�]ؒ�(qX�� .�-IE �W��&[�����˺����_[D�K%�vӣd�N����5e-�j���jɐ�=6��oF"md�+,�Z�9$�f���Ħ�����G4�6	)�Y$ �u���٫c��1�R�z����7@ ��`�u��GIA欬�`�/*���!7v����W�T�؅����Ӡ�!����o�Dʽ�Y�hk���V�i�O����`7�iEgA;�aWc������7y�4 Wse#�^���[t�-i����ۭ��fS���͊�3o�Cv�<�� ��`J�,:�׺��e���[��T����SŘ(c��Ki;H��H�bIW�u�u2�4���ە�Uk�	(�ՙ��E��i{�ZXiR&�4���.�U�<����;7cJE�{x~#Vf^]�2bm�υ�6���Z�o��T0kTL��֊�u�� �#EQx�{N9�mf�<+2S�/,8��v��t٢�/��ޒ�A�X��VPC/8��!��K.�)lȮ��5�L81������@M��	�kuNa��c��%��D�RŬ��Ȭ�-2��0CGf)/VU��VM�be��fEZ�j�n�j��5�A�� 2��N��]��s걎ֱ�Y�a+��E�����%?����U�U*�o�������N���E"r��Ԏe'�
�v�Eb[wX�r��ò�E��tP�M��I�&&(d�8��v��#��/� V�i��5D)( �:&���ս��R�6�o�G�w6���2�@t`�R�l#Z�1;'ri�EQ����+e��b[�ȫ�7K&�uwE��OZw�l�R+���l����*��:�c �6qr��6E-ɓ�H��R��K2�7[yL��<6j�iܶ��*��Y�f]mbO����l�y��0i�a��V϶�+0aV��cs+r�T���:�8,H��xl����Mj��N��Y)m��	���H���5�J��W@<M7K��܍�1�i��U�U6�U�`�(�T�����bխ	� �3n-��N�W{Z�$�`R�a�͞�T���n�Y�T�4-<��;֑�h������F�n���g2/�u�W�:�����4��ԹH"l%/��)��8l�w-���Lu��k���{�k�K�&��༻�n�̙�ܡ
���A^"lR��J�͆J��e�K)�L�p80Y*�̓BԘ�P��2��k66���E�c+�6��F�e=���һҙODm�M��+��ۧ#�{)�
B��]f�m
D��RM���H�M9FR��BV�h�n*I�)�-��w0�2��+M��B3��������6���!���%���Z�d��%��wTອ���.�"��S�jH@ȕʐ��wR`Z��n�U����
[�T�uu!��x���3&�0v���?]���F�.�Q�A��0e	����ۥ�K�ӟL��B��哵W�� �*�u�)�Mqm-��Ú�u*"�co���5T;u��^�Y�tu�?���u�jB�
w��^�bʅڽt�mb�9e	7�M��&��"�U��`r��%\�R�z0��{%���d� ��6`t��N�Z,��++�%B,9(�n���­Å�^�Y���8�H�7[2�(��ⴖL(���2�Y�s	���4�q	J�B�'R}rk´���kY2�*xh�@�C!�.G�*��c��eSEM�{P��#���K�a(�\c]%m�hY��ڰ���q�v@z��1{�(�z/���xl�(�b���m�t����ӫ�唆Y�t����b�<.�.#p�Wn�Bդ'����W�Kt EX!�m]'��NX�1Q�%©f��p�onԶWGL������2�4��H��0�]����6�]�0^sj,x
��k���]`�MX��a�H���]]%��U�|	������;��,0+T�{���3i��6�$��u�+��S��7���xXD�%�b�ۚ����	�n�ouz0&�CuS\IѠ���y���%U3i�m�3�"�eH%1)�짖h�k^�1I�'���3���n��|�K�2c�qV\��R����)U���%ֵ׭�B���9�.<bԬ���*���n�9IWPn�N]-:��5h�4�I�a�*��"�^��(,/rH��(,���VLx�|N���&m�ZH��$�CK#m��镦o)3����F���"��-���İ|y�b;B§�,�ŗO�qkn�ܟj�B�� &��UX`۵H�Jkŗ���X�f�T�Up�VLܑ�3*��re�-ꡮ�Mf���X*����o��WNj6�:y�M�;�d���t��+ko�r]�X&a�Q�Q,%wkFƌ��˺�}0ʔ[��(�+�[�e��O�i���x��]Z��V��i��,Mӻ�ƒ(� �#6N*EBn��c/\ZP�K�z���厛w����t.�Z�$^��W%`���Y"-*�I(ҷlXN�3H�zͺ0ښ�(�� ;,�����C&l)B��)�a>x�Kl {�0����ނ��wan6�e�r��Mk�XrV;B��K]o�V<���\���k��n$��:5�<�.��U�utN=(*bT`&��+ܷCU��Pn���NJ�e��(%�[j�ˡ�Q��:�\��j@f����K�YubL$���EF�Q��Y#�Ԫ��)P�ib"�ZvN��.�����t��@�E�3��T�`��͍W�43���s'�IB�:XZ}�c7t{5��Z���905�l��r����!��������8�eǪjҶ��X7z���c �ĵ�EAVV��Orm�����C0己��]5�6�^+(+ӆ<q��P�FR���ˣ(̏Mm��ZRR��0�+F]a��,H���j�ϵ^�ަ�;����V�U����bUkR�˺�L'ofLb����v2l�#f�����7[K\����q5.YV0�T��,�Q�nS�H�(T	�d'����⧲�ԉۤ%EɆ0��6R�HnFL��(n
`��0�v֗��|����[�L��!xb	^�de}1�ac�x���7�Լ�����f6�^��.����ܻF�?b�-�c+f��b����Xn��e(I�L��8��8�z8#n��!��;\���&����yZ��C[��Xr=T�k6�j�U����L���;�i�.g��v�":��e�X�E������P�����O�e�����́JQ�DǼM�#i'�u�-��B+Y�՘D�kPF�&%k̊蘴�B�Ӡ۬)Uֲ�=��W����Z���bY�Op��ƽ��I:[���vfTn�SeebE^��Rue���ԛ�4@��2A7zB#-+KVV���g"�N�y����n�|�o0 靲�щ��V�ZЅ���Q����G��@��"�X��M`c�rY�ټ���V��Lcv�æTt��%�V���F��;��b�v�/4�Eyd��]nd�zi��j�Tim�#ܚ�`�v� i��TE��ZҤ�ϲo\�Ɩ�gk ��
;���U��1@ڙ��i֤�Pޗ��TFmڛuq$�6�Y�d��G^�aʳL:�3F,&ʬTL%���WtKY*|7-�ɛ�m�R��BCH48fd5݋��z�*ZPH���]�V�Uhm�B����dq� n�Y�[B502j���h�fhp�@�B��7��N���Z�4ѡSr�t!Wc'�m��p	n��p�#(*xԗ�}"�{����x̼��Y�Zۼ�j[�c��rA�Ӳ5�^�	�Ʃ$2eͽd +h����d��-n_��/4���h͒�����J�b�w��]B2����Nj&غݬy.�8��v�2\8�L�T	m�dWYzC.���b򐰮n֌�{�+�'M*:���3LW��k7X�׭�f��v�f�+6+oXJ��V��kQ%ӳce�`�V��7
�VҠ7�x]�.�L��#JseC#��[���aԫ ๵�Z����m��4�Y�Ӵ�����W ]�Kwp�+p�v30c�J��1/�8��a�6�Ђڕ`�$ 7h���y�S�I�/n�f��ж��D4� `��邳)�YJ\��6m�A�&���l3Zه5n��L�*2A[՛d�9�<��5W���V�c�O]�VS���f	S*S������ )���1Ň^�o��c,?�w��;l�C�|����[����b�=��m8��dh�D��e:�	��6�be�N�Ԧ�+��Z�2����g)�Иw�N5o(-�՗��K��-�e퍈�n"�UbZ6]�N��MC(!�������E�mK�ԋ˦k�ytJ�;SY��ѱ[F��v܆�Į��R�l��������HE�6(�Uh*Q���2�#Ud����G,�;�˓�k
�.����Ѿ|z�
Գ�yl�Av�Ww���Vmq.�Qm�=zR r)S�P����kF��On������XC�1������!���օ{�,p���v���
�ER�F?��{#̙{k]є�9Z�ʚW>x�
���*Xz�H,e0�4��D6�7a�W�I������]Z����t��xvS@޷waV�4�|��;4��]�i$��5k���uAS*�L�gj^M��������Xt,.[t7U��J7ir�Y��pc.�7Hr8�,��ִS�����A�#.��P����eE�w��'&��%c�Y++�D�vF<�k.^c5ޢF`̮A[i��ۼ|f�$��/��v/(e��<��]�Kx���ùGK�{U���E�ae�KW.#�o[9�q�x����;r��X�,d�
G��Ot�vzvݵ�]�WI4�޼�a���˦�j�!A��WUt�]Z!�Yh�mZhbǢ�9tqm�z58k^��K�{�,; ����-Ȩ��*;���-�̻�d&����jR�ۧPX�
EFC���6
4�<=ɰV�2�.G*�vo|�s`]eҢ5�=�@��d�זҠ�Y����eM7���0��W��^Çb�IJ�� ��2�+v�-\̹yr�H�on��)���/C�6� 5��6�DKF�f�\ɱR���S���/K��,h����{1i{�5�
��.ցE�����m�!�U����#e�;�n�Ӂ��G(�mdʌ�"ɺe�wʚ2�ּ�7FG3MZ	�H/�=�ˏ�{��m��S&]�4�r�-��[N*�]��q�`�H2�!��cJ�J�Xm�]�O5f��3�R�8ލ�N�e� N��7gV�l*�L�g2�hS�A$��k���s��n�@Ɲ��31w��
�)YW-�*�����3C��0 �rG���F[ԍ��h�����^̏HV0K���WwI:�H4�jbhnT���a�NP]A�n�Ot��GE�v���0�0�e�U����#�Q;��[��Eۤ3�Ю��L�p��F�fV�䰪��X��o��-�',�$Q���`J�2�lM=�@�-PO5m,K3#�d�a+mML�,� c���]�[[I�c�:�z��L��˶N�[�dm��k����5)��,ȑm��S4,��wvt8�Շ��D^�Zs�6��K;����^롩�͛j�u)�[5`WZ`՛b���7�6�y��iỒ�Tm`��<�)��MCF|]�[f[�Ǹ�+	fB���h�u�`�
�d0�S.��{��Z��*���K�n�+ *��p�Y@��̈R�� 
�.b��Z03*��5 Y �M�R�
e��
C4]'�biF�m1�l$x��ᥫ�X�x��:���;E%yv0��1�cIS�d�7��mP�yr,�2����W�)��]ς#paL}a�1���E��]���u
Ɲ��;G�P��)�gxuj�\И�B��v]�Mf�=t���Kv�1��E�e��C��ٍ�C�ׄ$��v�F�h��a��Lc���Q�U�F�j���v�\)L5Y[�Ӥ��jЮY�̾�B�e�Q	��^ֻ�!U�Yg^���z�ڱw���&I�3:�Z� ڛcE�2��k)�(��p��R�$�z]�$-ӑ-ܱ��n��=�O�Vr�ێf�kZUuk��o�u4�2�Y֐��x�����Fll/o ɋ-��{��["�ݓ+v2�GJ�k*�m��XqZ�2�g�^ ��4�'�"��Ӝ� ���ID:��e�h�L�q=HR�U`�oV}z�E[�7��l�=�����b�p�-��;����F�}H:]�9�h�%
��ε���QݣO�+��
�N�J���]g
`�i:�I<�B�}��k��Z�WKq�[�P[�oS��� ��R�hC��n�±
n����5Q�J��M\@�Q����>�˛R�+6m�[���X��N�=�]Jn��fLi�X�X�+3�D��@�M!htfd=��2��-4˧E^�`aq*tJN�j�,Y�{���f�Z�8��4h j�Wl��Md�V6�v����K�B�wvkbU��F�Sţpc�)z�j���qok��|�ֆ�[Y�&,�H��kvX������V�b��EQu�n�
�cg���`�`�+&\�Ĭ�v�ۻw+q��^툱ūvɇ �"����0����>vZ��Zwwb���`koF"�L�e�Q�{�k0�{�&��$m*� �O.����IoR��V�FQ����k�{8��GG;{H���b���<Hc/�䭰�/�ӝnR� ����so���N2�Бɑ��vz�y=��=��;�"|�U��ܥ]Ъ��*���a�ڝGFi�r�%(&��9�|��핅+��˝[�����ln�������k��nK����(������qs��U�>���&���F���9G8u?�տl?!�[�V�9��;D���e��f��"g �L��h��U���;󔳷ڕg�M���c*���uD�7��9��ʴ�Y�9�F�ĩv�����u��t���n7&���;L#
ܱQ>Q�'o���y1����Aq�V�����"�թ9��Zzb8�rge�s�R ��X�/�LRf�^ъ�7��X.;�;�n�CT[��
暺	���s���k��r��*>yF�����+p���maN>Yka����;@[�Fٓ��u�"���ͅ���4k-��'�սrԚ�
����w��G��g.��a���j+��@�TsC�2E� yܻ�ZxH����3�(Q�X��,�'E�4��.�M��7E���p�o �Ø���f�� 
�G�����ģ�;���y��CNdޜ�mn�$���.�.�/�@�śs�HO:N��F�	�NW^�J1�35�Cm+��7�����i��ьս�{Wk��;(�O*�l��βR��~�<��\|����zi�{6�Ы�JmD�ۦ�o�eMr��V]������M�)R���e��s���͗&��Ry�I�z��fvL�w�iB]CI��}�WFƛ�umrc.�+ڊ��� �xLnŕj����U֮Ox2��2���eR����y�ٺ�/9+i��c��	6"5��y£/��_-v�m��)J�"D~�+]�!�����ˑX.�ԏ����4jR�^�Ҷ�,����<�E  ����h�g(�V���;��;�����#l�{�9�r�p
U�a�ɽ�)[ΈCef]�i�c��m�a�u̢�A�<��ft���^��<�
]bVL@ȹF�7]���k7��Y,QRt8��;Vtuq/d&T�\�q�NN��J]YPp����V�B./.h-��34GWy�$��W�vn�>	⧵3mr��T���je5���έ��m���!���wD��z	���}!��`r;�e
�(��9�U�6�d|���tj��("�6�<�h��n�*�#����.���.w��&k�)��6�dut���%���XY�eX����6�B2^jd1W��2䐫�t�M
m�,��ژSOhE�^m�YS�,�@�+���i��&�z8l��2'����V����́��m��''���-�_:�M�}����m(9� ��;�hu����Z9���!���a]�oi�m�.�񗘓eh�3�Bŷ���<�/+eo"1�^��ۍƅ@�U����su}+E�9��U�V0k&��� ��6��1��ʂ��Sd���#�6��������_S���uK����}n��HMfQ�"}��S-Mg^gm�G�i,�R
�E�42����[P�	������<Ot�6�]'t�Y��kv�j�'�Bh�����^��m>�zQV��Wq��1M���.�i$J빹|n�k4�v�Q�F��]9�&J�I���5ԃ���=1�cqMnp,�u੝���%�n��{[�9(��fVU�����aήHWRw�h��h�)Rܡ�"�����N�;�g[�wy:RT�>���%�,��P�u��,����E����%V-u���R_Z�����b�o+����!�	��̶r�b�
�1����,�fk��pa*���jۺ`�� X��9ٯ�q}WwYE0&n}�f3X:�X��*u1�M:�EX.��دJԚ��s%h�T��Bc��;f�R����|.˶p7��r����]2,.��Z]�k]�$���2:��:��=�I�X[j:�����Nt�%3��-��y�`WyP^�9���>�z`�h���ǌC\։ZN�λ���(N#���-����E��je��Vj��u�4_�N�Y.Z�]������Q!�wRL�F�ݗж/V��$wr��$ɐ�mn+t{"��OX1�1��-�{�Q|Gl�+�7�:�n����`���ʲ�W
u��s2�1��V{%��B�oD�˱q�)����C6��uf+�},��JS����WA�R���z��׹�!d-\��w�GA:�Ԫcǵà��]YI����Af�W��8s{��Y$�n�:�4sBCt�lxf�ӵ9���퉰m%��@)8�eS�n����n������ˇ�>g\ں
������ٵ.���;���)�+$y�x�)`�V�ˏ��-�b��w�-�Ͱ�5�T�z+���ס!Yۣ��Q�.s$��
a��p��}F9A3G\N�n��f�Z�֕���L�d� djo�u�&ek�(H���`�3��we���֮F�qW-u���0m�pխ[�)���`Q����/���]��AJǸM��P+��VQ���{�`���� 5C�V�fm4�qg�Jkrv!t�����m#��j�+�0q��k���7>�(kgL2ʥ\)�n�\��S
puf	�zj<y%YYJYѢ�T0o.H�e$�S����wg,Jŝ��7ŽVt�7�ݢ��+����:�ݨ�3tƮËFB�;��9�m3jn�)1>�\3�JN!�Nph�%M�ܥ��S`�9���N��-g]9x19|2��VOL��v��Ž�*=c4魛*U<ʽ��AN�R�JWY�i<d��)[�cy�ؙ5�t�6.�tU��#{�܌fN�c��^ЙAlγV��������RPT�=�p��1f�򔮜A�z��/�Zvд�ǧu:�îb�]�u�*��GX��,,����ʄ�h�U�g�_�A�v�nb�hM?�S.��#�;*���'�Yb�Iv��
�e��f���Ik��{M�e�4#b���Zwr�˼ݹPV�mC T�nk+ww���UN�QCfd��n	��n��@���������u���mr��$�8���#f���0�m�ZGs�3�;D�]X=�(������J��ft���:ZU���k�H,���Y������	�Yz�H�m9h��ehL���|�q�t27��qqoi��\y묕��V�ƅ�#O�7m����!�m�=u����Ld�F�m3"�7���l�l�L=ghouL����m^��R���2ԩ(L��ổ�h`���v�)F)�Ő���O�$�c3V�qr��=��aX��]��2�f�|�7[��3���C;����E�B����x.��y�t��ͳM��u��u��Xh�:�����~�Aq�o-R5	2^.�oWT�'q��TcۂVnQjS޵7��4��5w|��-��z&�3�w\؆`3��{[��"�r�ז��Yu���QN��[Q�O2Y0m[Í�9�ސafɴ��ܶ�L�+DR�F�1������|�+/�Y������p\:Z�u(v�s6�-q}��YK';[�6.J�q<���۝ n��7#c�vB����l�Ҵ��T�>v(.����Ȝ��Lu�*U��bq\�R`}ʱgE4V�έ8y�2
{��/(;4��4�+"l�S���W(s]�9!�����4���p�ҷ&`˓��o9�֚G�����@Xȸ�4k8�9tVj���$γÌ�&��d�2�L߮j��M�+�U�	3��.QJ�܇j��Ȭd���:s�����x%q����m�rUb���=��?|B��f�|�Q�u��nX��sٌ�l�Pb��]��tD\�k����/WM�"�n֤�=�u<q;t�sGCov��v9V�c���B�U�:�0mk��xu�.h��� mk�μ�' 8�E��	�ӝ[�ṃڨ�z�)�I� {��+B��z̕/(�:�r�®����������}�1t�;A
��H�@ioD�w�@�T��
م�D����V����
gnѣ.��3�o%��$�M�7�|o�sw��zi��j��ٴ�έ�FW�Koc'�w�k�'c���t<F�
壭6��ኳ���3��d�����(x9V��̭�n���r#U�Vv��l}a���S�H��������"�l�V��	\���#v�M���ֈ��n�|����}�3Aj'{"o7�16á}�ԋ�	�OVS�.��!��ͱYA:�T�ġ�*���wi�?Y�ȝ۾u��;,a�+;��-Z�fTR����Z�;����w堕�7w'r�H��o:�ۮ� ��ZD�T�f^��z�Ń*WV���5W����uu1��R����MK��7�a�.��7�n(pX�Sw�$�+n��+:�B;Dni�gK9\Zi��T�0�a�3Fmp\2�A*���8*-��㵸S�:h�X�Sp�ۡK6V��[AhUo��q^��R�w�/٫��]��/=���[�Ζ�g]*��&�2x]h2���m��������{�2����W�˻n��/N$To\��J��EX�f(�S���«�c&4a��m��ˉeD)2���6䮧����e�RwK׌��iV]ɹJ�pu���y�,@�=�d�:��P���e�}�u)���;�]t��Zѹ�J�]�z�jRƃr*X�}kZ��5��5\�+5��b�N�@�7��Hsĸ�5�
�5{Ў���ۮ�ViW1f�wԹ��؟v���-��e�g*����f�d�ƹG�K���ri_����hh����p�Q�)�>�Wv,��������R��Rv2n�%�굦���ܰ�P�8��U)*wwn�u,�w��(��#jܜ�S��Z���d����r����	���aK�,G]M��:|ɜ,�]�V�j�K쳒d�U,����}��W����1J�B9��Kr�09X�E��SUd�v�Y��@�̉Zx�COz��7b�
�Q� (v
l�ѡ�GF�S��Օ�ZG(+����v-�wBs�i�R���69Sz�҂��m�ˏ���ѫ���ٶ���]�Q�x�[�W܇]���]�7���c�n�D�B�&���}��^�0�p$M���,����W�
Ή�$���gZX�mN�gY�y̜&̊�^��.7��d���q��VcҴ=�3���ʽ��7����S�ԗ)�ˣ����{�N'�]lڌ�J���묥�Z�iT=�����+q=MMKv��H��ʹu��D�i��=�v:ͻ�y����o��xZa���ZHo�{yo3����Jt�B�Z	�=��4��;vgW|:!�]��]ۏ0R�6�aL�=ݹ�\�X4;@V2��jީWˈ�j���|����*Q,��)}s�� �3J��Z]ٳ3��t��N5m>Ju�ea���l��+�nu�f-�k3�=W� wJ$k{p�-uXj�v�֨X�P�tfs��W�Q�� olER��*�(ѰP(��:�e�A@�u��6��qˉMn^�C9�{��s�Օ�qԬA��w�X3th�y�u5uh�j�k���|0n��Q��Uv����mK��l]ؘ�Z���G��C݋�[Qd,�)���[�u���-��]�gs,C9�a�:�n ��Ҵ�n���{�n����PQ���n((l�B��0����U|�fM��9`��"����k;�� T���LՔr��0�u:��ecr�W֎�@�p;���w�.�=6����rmіO\�8y�!��je⭳fee��EF��r4�}X���!�<z�1d�(۬h4�y�7�]q��ܫS1�^�d��-��2Zu�e�&�q�%�~goX�K`�;���p���α&��uR�(hw��_d��Ս�#�x���9�jrՒ�lõ��P���4Ib�^�}ݮJ?z2�P9|��5��v�)���n�Z�s��>ה8�4mw<�$����ݺڵe��I�,*��:��7K�V�S3F�I�o{$�$�䳐��k�8_9�Jg&����۲��}�]ApK���ˇ�	�0h;I^9sR:NU��k�s��mN@��!�Vb�4l;`�t-ЫN�D���q���n�{��r�.9DL�76�S��rau�L7f"�і���i�י����u�'"M��t]�����ɿbM�U��#�ڱ�ԉj���wm��ŝj���W�1��e�=o]�A�; i��Da Q�wJ�0Ԝ�V)����w(b#�q}iq�o�]c�=œ4J.�4�L�Pfj�9;��UN��4�`�I⨘��0��31c���8(���L}�}j>��V��7�D�"9����B�ɇZ�y-�4io��o�����7�u�n��.����Ov�t���h9�v�:��tg^�O�r�`P�u��5.���nμzΊ�Ӻ-���s_R�+z�}gc\,�
d�;�f�|@rb]scwA��N�dp���������Q�;d^s�oL_�KT֣�3Gr[^�x�%K��%��cԳ��b;�I/�<��bm4+���r���H/�w@�.��{8�ѢJ�Y���fv&��ǲ���=+n��3(&����-hM�$�F򌆲� 7/3�D�ճ�:�m����%D2Z�b����%��je�-����p���a6U<�˷p:yN�n�Z{R7��S���&���+�L$�d�<Iٓo�����i	��^DwG0��k[���{�؛91Xl��"̂��J�t��ǌ�2���(�X.��X��[ףz����̆�͢�\�ܷ�j\m��4����2�N�]�Օ��X�m8gV�EF`2����nϵ\9�`���"�i�]�F�cN��MDիIf����
1H��a$2���r;�XΓ���@$$?�	!I���u�;�u��벘��$Q�՜�p�:/5�ӹp�'�u�o��6 ��z�T(N,G�']c�{��t��,��el%�T����<��Y���Y!��
��L��0a5,�1� ^�g W<Q���q�K��[��ș���hT���
3X���\zv�ɺV�-龦͒��r�t��S���iHkJUNo+�#���U����5°�<�7Yc�k�̍;n`�/�m�}%"�a�\��w��8��8�]���q������`�ݡr���-�A4�4AWf�RJA͹�F;R�����"o 7�.h�K+���H]n�3$6c��i����˦��4M�Q6z�>������v����z�w0*��S5t�z�{�'8m*ul�	2��;	�h�1�3z��Y�v�T.C�\�F#��]�z6��ݒ
G6���WF����k�;y"�X���S%e��f��q�\9�>�\���c��1�3Ҭf�ud��V(�ht�M&�c�rn�\�{�˭���%�3�u.�G�c���n��ҭS�jώҵ��:��AH��8W+/����N �ە6�^}��V������˱5+U�`�z���)
bD.�p�6p�Ԭ�t�>I�{���yT��iXkw���'0�-&�]�x���4unb�$�8np{twr��,#�U�Li�=	\�wy������2s!��N��rb��g;��.y�e��YK���M�)��B��`f�TlÔ�e&��1b��V��c0����뱠%Y��(�3�e{k�7)�4��������s[oR���Yʾ͠i��'X4�4�ou�0���0t��&��42��U�MƙB�X�ur�=@�7���0�f9o]�5e.��那+����[�]O�Wu[u�����EF`?e;#:�2��E\�[)M��/����Ċ5fao&&�fڅ ���=�]P�B�h� �a3fJ?A!"���Ӥ�5�\>=�b��m����ok�[�1!N��k��(�#]�5�������)Nv�c���B�����溭���E8G �]���V�.�Y���Vْ�O&��X�j�ى^+2��A�W^E�랫4z)V@8U���7X��Y6M+�m�� _\�r�n���g�{id�E>`T��e/�n@�hm�J�9mkwGxU,�cYl�bn���U��E�� ��VY�-¨��-���K�,�*:r���W�v[25�k�D��9�S
�K�%F�l�R+��������٣p�5!�x�i�J�Ɨ:��[��(#n;���-Ζ ��`}���weO0�;2���}�J���� ���A����p���;z��N�U��4.I�d��NS����+��;̴�l)�*���|����K��A5D��j�tfM��9B��w'1�;\��u�&�W��b]��p^b�:��nJ�++&�sZ)N$4��5��;����[f�]�����#n��F��j3M��I��f�Ə*V� Sz�pWS�v{��Vm�TquLu���B���3!;6�[�ww�D�kvƲ�]��ە�Fb�^�;2̵%D�d�;�E��G%B7-RؤэNӨ���̋4�9Ymm�h��[��ڎ]�j�-ܭ/��X�;,��N�z6�<���0�uڶQ55�бi��1�R��0�ers�4o�+����t�}
�TZgV���:[��7������������%���t�$�u�v��mS�Ou^��th����k2Q_u^]�%@ꝥ%Q]d�{h3t�d�o�uyB��
֍n<���Μ9�.��P�4��֧X����v"n��V��Q�f�3d�����r����	�r�ɽn�r�t���
�-%�vKɶ�ӓ�A�
�����Y���cz�s��0���Ñ͛��|���7��Z:���$��ɵ(�Es��DK��t��;֭F$ p�A4]�el*�j�x@w�t�9q^F�0�p��	W	��x��v���\�jLI���n��y�o��I�a�h�Z�0:ɧ�%B�"�9L2�̓M��/:"�,��5� �O1wNY-� H����d�le��
�gt���kĝͺ��w*6��=oi�:j�OrZ.��Z;�sfK}DU��03�'o���am�jSy��P��[�v���&2�:�}��4�u;�6�V�����V��<u��<N=�:��PWo.��v�Dl����^����-�|%�\ƅ�*�h:���jt֜�sr�T^jk6XWE�*bm^��L�9�q�N�R�r���	9VU�]� �0�w���g!p��tw���Cn�i�I��e w-��Y9;�U�i�H}b (�uϫ�ܤ`�չԶ�N��R�ᔫB���Z²v�:/78^n�R�;V�H���.�A�j���q��A+{�:u�3w%L&�WHHJ�F`�DC-����̬�&�=��·N5�B�'R��Ne�@&�e
:[TOdz�t�*Ż�9uڵ>�K���M�4����oP�1�0�C���1��'}�⭔l]��Djۧ�b��p�y�����G���s ���b;S�&zr��<��+�h��;nuAh(^5/o���m<�-�5�+c��3�,�啘PB%Z�s�-�W)�C��Lсm�/�6Ϊ|&��Vڊ�e���c7;�=@���[7h��5j��	���,f�N6�5s��pHN�jS��H�e�ŭ��r�*���nîPշZ��`��V�)B��R[��]�%p��[��������,�a@�r-��V+EB�Rf��owur/��G����;�r��u>��#fSD���Ye�ev��F��\����5���|[ܺ-�V�n�z���*��Z�
^i"k���V#J��
��,��%K��!K/.d����o>m]Y���uj�4x8��$��9ec���>\�%���dւ�W��Y�,��L'��{��/���yG`�����nt�;*�*�J7���Jp�=���Y��'�EK4Q�7�!{��V��_w}��N�>B�P�{{��;\�JC�I�w�{�������ye���5e�H���j��oʧC����j�)yr�n�\t��j�Vi��@�&-�¦��\�&.�q��D�0E/#�x{iŧ-2'r��-w��Dڿ��ps�r���;j7]����j�/xˀS�״�O.�V��ud;H��㥺�7� #��wX7����Mn$��V ��u�i�z�앴fI��L��fPAj�������δ��ue���}xM��U& ���R�KVgp�T�`�9��\��VGvN��N�N��h�s6���վ�t��3�$RVe^��;�Bc�]������V�����^l	Y��l�g	�Α�e8j�;��E#۶9�Wxl챙˷h�R��&΃�e�9-Ѭ�����K����ɹ�|Itn�t�bR nv�br���r�z��2�y��\Ȧ$��Fp�sF㵃Sg
��٭�Qs�kx����䗚�U]=�Z��������u�7B���}�����x����^l�J���Z�r��9�^�)C�Aw;�wֲ����L!�p�9�k�E��ׇ*��d\�<����hK����>2��tiQ�ڻ;u'+kʃ�W7+����mϙ�OU�$�*��4r�nGc��n���H�E����g)Q�yR*��z��3s�z1����h�L�:ȅq�@���&���hRZ4��΋�x$�>�y�ۺ*��&Y��Q��:�At�����w��m�ט�����)�$ϰ^������>��iTVMCh�`��.}�|�
�j��ܻ
�9VT����p֚����rj�'k�͐��(�׫1�"���ƒ��N�,���a4՞��6��B�k�N��>�h��=�	sf�};6�4��_p�[�j��4_ӝ��[�K�����D���GZ�,q̝�r2mvH )����y5����fi�r�t,��q������k���e�xV*��B��G^�U�����q��&2ʢi�Kx����[�=���F �dN�e�Ƶ����G�ҩNMr*����)^ɕ��'��{[��آ����^t�,�#!ZC�G����V:����:�JqL:i5V5�����A���;�,��EN7W�|a�E`�U��]g�Pv;�0nK8k�kA6)��4poq�Y���29u��[���(g=܂��g,-C���6ֹ���w�XF�=��[���懡���\��ܥ�H4���>*�:��|��p;��b���i�]H%^`�����6�W�7.��ɮ�����ٻ�E_.�y�H��cY��
�QAf��9�y�8u۴w�skn�S!��v����o��`�:�)��hP:�s��B\�\.��gs�Tgm	��o��Rb(�2Kc5��x=��\�eҦ1���V��]e�$'I	qn�S�ڡ��� gP��e�ԭo9��T��P[��&������Ն�Z��bv�H�GP����N��磜��g�霦U���X�3ʥ���h�m뤛78��V�Lĭ��>� �y��n�*QZ8�={rT���y3Wp���ӊ�C/������t�ʘy�ޒ��,w
�a��K��J���ڹf
��\Ӗ�Y�z�qAF���y���G�
��sӺ�ܑ�U�[�d����E7ͺ��Z�a���u�q���ʅ_g gJ�X'���1�-��0���{���V7o&W.���-.�ʀ���0�5���ݣ�i m��r#�Nnކ=�V���<���o�hg�t��1b�M�\�b�]sL�+�%�zi���7{���y�b�km	��V=,�5��Ŋ8�3�d�K1���m�Y7��u�AM8Q���1�shi�9I�g=%֊3�B��W[�mJ���'[��[�Y9 q]ּ˨�Q[r�ej�L!f���3�Dm�O/�m�2GK7�wF���V�ٴ�4/@��]����fhp��1e��V�N�-��Cf�es&��� �L�@[Q��#J��:^7r��la�b�v��y �����8���j[��FoR�e�`*�RڼK9�&k"���\9�7�]uj��M�+0��ޣB=��L��E�5��O_5U�]+)��:qε3�����ˊ���aݒ��
�mᏴ["����c%��VOv`�K#5�Fu�r��0d���AJ��¥݋RZ2�g'I=�]���gtY�v�{��i ��ƺ�KB]룚�(�ǝ����=�-�0��/e��A-��9P�!��0�-���qއW�X���b���Z�j�k�m��V[��ڙW��m���qK�66�2�[�D�/U�{�-�W�IZ�D�ڊ�f�v�JA�Vh=�ѻil�=Ұ3�,K��U[�Uú��"W�lE5�%�f�>޷�pw���ԽS;�)�P~5j��M��t��P(w;E�VT�
����cxS��-;�2���6p�䕚��	't존�ڋA�U�.��L;&��^�͋��Q�ƅ���VCV�>����cUt3p��z��U�($�7�5G4*����u��GV;ÃIې�u�S$�)�ݔP��QQ��KYΔ�7���5`b�eN�F5����ZS�Xyi>�k�pK��ݘo�b1-,�)k2�����u����#q�h�+3�b�r�Vr�}ؐ5��]�V[�RM�=KF,܆�^�o/6i;��w��L��h�He��#�\릎*dl�����Y���vg8����>�jk�foU��Rp�od;�$���x�y
OZw�V=��{ƖQ3K���-�ݥ]���b]��2E����fV>���ڜ0�E�5��6*É�,,l"�IV��ymګ�gI&����iD�l;J�m79�״��� r��q|�]nuAck�e�)K�-t�V2�OY\+
��ajN�z����I#��f6��[95Ӕ�^$3 ��Tf�ѻ�P�#@.��`����]��D��Ao41۟7u4M�.��o3i�XXܣ�;�����Y6-1�[̵��է»Eʀ�R����\�=	����ZWr�*�Q`u��'��t���,��40�4#�{�-m��pѻ+,ӻ{h1��q�!� �	�1%�{�	�T�7� 8����v����5��nܻ�rq�W(�]�+�u����!����4hM����,�/Cݔp�jR�ݩ��pwi�_;�L������]sڡV�U�n��Z�&�ʷX[Mp����	|-���[i�Φ�̅a���̹�#9�x����p���]�u�JP�����v�	RfZ6���w�E����P���tGu'q�J�.b��.z��f���\bj9��9�u�Ei�@5�l#�8K|-p�xM�!m�ȝh��5�Kz� ��B\��U�)#F�<��`O���kR��bk׊N�7/�N	B�:�`ff7K��\�x���|F��,M� e��1����;c����A]�k��UJ��Kvmdr�p��*Y��s�<��ovʌkH[ޝ
4>�.���ڎAۧz3��l��0�#wx�(��.�sgC�F^�(_�g\�%c�����5+*E�(�wړ/C�F�R�d�����;=�GWl�vu�'�4�Nm��9�u(\X.1"β���&�������y1�рq�5��70�n��sC,-�C��V���� �Ru+N<'f��DQ0��z%у'K�t�){��a�Cs����u�]�us�ܡp��3�+�Q_���W�}_U}����]������V{u�r���}yP���ܮ���ة=�jS�~��i�8Ch�Mp�ӛ�ǽ����ziʃ��ս�9s�v��<�T�#��Ɗ�Cb�b�O�G0EY�X���25���Od�#�O��,����z�J�v��wP^(�� ��QK+�'X��q��V��;�-�J�(악>2���[�c�����g-A���3�ay�GR����o-�D����Ʈ�`�铣�̞j��ʹ�{J���ee6���D������cf�&������]uֺ؎B���k\����G�캱��pPpr�a�B�N%e�5}�j!K��@<�Wm��\��Pvܓx�6�^�FX݀я/��=�YS5o;Vy���I�@U��,B���ľ�Ν0�Q��	��D�v�[Dt��g:�Y;]�w�*��5�.IWک�T��U�S'$k�<�WF�w����}X��6�)G(^��dr}���w�{f�6�`t���O�hJ�����u<�e��b��E�UbŤ=O�;��nm)[5��K���gެ��g@�M��Jo�=`�6��t�7�ݑ7S}�9ŜhJk�GT��������U��	S+�wy��t�zi��nF�&�3j]���޸ts�#rcy�1�ARz�ۓ,Ӧ���fq����Ԙ�qY>۰����[j�%\�!�)�Ţȥh��*��pTR�ڢT�H��YXVڢ��(�%b�AP��AE�"0����VTUU�(�.2��U���K[X����L��̨��YZ���eb�F�mq�mh�V�+X��Q�e���m�e�VZJ4[H�-i*�+ZQ*�����kliQԪ�U-Z�b��2��Х+R�ie�e�Rŭh��,U��V�Ĥ����[km�q�Jֶ�Z��*��*��cR	�R"[*U-m�$�kQZ4�VՖԴ��Q�[k
°��j�Z(�-�f9�ƉQm�mh�F�b�"��R��ib�����
�մ� �V�E�h�*[J��J�lb%h�*��EJ�J�Db�ŊVѩT��"�QEKmK
�X�cR�+,�Эk"��*�V�Z�%��\����*��ł*�mm*V���}��s�;��%yj�S2w#,�)�˕yövS�R��u;a����(pw1�_Mf�a	a�Su�L��2v��tum�����J2~�i�G.��t�4�`��]��`\b
`����2�t��h�.v���ËS5_ڽYH�e(Q^���ޞ�l�4�����uY~����S+7::!޹��m+�,�qOg�$&���������nY&+��A*�m��E���Ou��O�&�u3�wU�Ts7�AWG`�F*֝"��B�[Z��D7=�O޳g+��5��m�!zDEx�d��(�K�s�3Oa�y{��O�:j�������z�-�G!���q�[��pޠF�
OR�Y+5W��wz�҅�
/��y�~����Ǎix�
��W�G`$N���{��[$iw���6��F�h�RS�ù¨�vR%��C�C�.��w�eD97&c���S��nF�|�_)��̅�S����OPF���J,
8���N���#�G��H��ӕ�=��nv$��Ϙ�����=~�[)Tj9l��L�q�W��",� �9�¯������v�
��s��F��M�j�-]��uscѳ+^i�Sv��;]rWhTm���L�cWr7��0)m�R��`���'��Tc˃f@�wu,ya��e
��8��w�KG ���y��ս���{�)k`�~���ʿa�1�Y�0�i��f�M�o������X"��'q�=:���Z�иKݯ6��Dn�����J�(lT=Lq��U}����t����74:�s&�K�kK�5�z��9-��X�Nי��F�;;t8R��� v��V>�=�l��c-�h�չV��C!�3��,��1�6,H�W�-l߁���<��L	��e�� �[S��Ԭ�W�����SH��B�������3�Y�yX����D�8_�vWl�ǁ����m�/�#־������0����%J�,rӚ�H����$�4���:T���=�6~N@h�2�� Ldr0*5�1|��5��f�*P�Ȫ�Q84>x9�qn�a���c�toP@[�t�u��i/�Ɛ��m���	;5u���,Y��g7��w�z�%,���G�o��9H�C�������X.���/1у%����gw���i�j���=4����.�:��
�G[�����ګ7����Z�����VVQ�I�g��n����=-������:��P�r�N]\g1��{k�G�Տ�n�ZZ�}�:���hs��# ���s7�����RՄ��(lg2|���
�#�D�����Q�zt��9{;�jg,��30d��:<JkK��Y�.�v6?a����!��,;m���D�U d�e��v�9m�a�q�!��,����`P{�64��V��=�1�CaG|�T��u��kk/j�rB��qx�a��"�ˀ��mU�Ѭ�P�'\K�r�ƅ�sZ�=P��)-N������KV�R\��#������	-��+�^�~������O��l�w!q v�9=h����y�B��/�}򚼑���R������^������f;��&�f:���Ş+V�2r�2�P�Jou�SXV�	�{�9jץ5;�"�dds$�"�4w���BW���{��G=UX�I2s�6�V��GF,+��칝"�J`����ה�XJ�%1����i��Ny��Y��-���&-��v�=Br���=��:���<5M-���'blΝ'_��,c!���c>ڪ�CFoM���i�l���������������R���C�V�A�&m�q8��;�z!�n{���8ۗg2�z��if�M�y3�{��7�aU��a�M�MU6@��k���]n"�ո^��;��w�B��pXLޞʙ�s+��H��uʭcwR1:����,㭼#z�`kS��:�TOHxk������� K�S�n_�C��cۧvC�O��wW�r�-RJ۾,\Lk���������-��ڻ�C�=,�uҙ^��������_��?�D����޻]R�V�}�=��;�5���|@�9���R�{��
�	Sx1�IC���{�˛�8K���<���u�<#~����hoI4��"w?�fdcq�4�mm�U���.�¯O+q��8�(k��O���۸�џ$E���О����ׇ7):���R͓A�2��-�E�Z�N3����^�.�/n���ΛUs��Z�"�g]9Y;m�k:� �)����/8E0��|���ښ��쭊./Bwn=�p���VZr���-�VCv)�X��)��^(����`��쐻Ǵ����Co�tn:3� ��ٲ���w4HP!�ԫ�{��y)KS���Q�=�]1�+.�C!c�O<E�[��womf��"F�8I�;�`�(!���,��x쯆(�x2����]
ډ���]/����QPz�������wQ5�ݧ��c
"u14Z���x��Vd	y���S�1�,]_V#Xs3l���I��F�s�x5H��K��9يKeJ��-�m$���}���훥\�f�E��tM�u�9��To���nh�|퉘���o�&s�V��4`q�@,+n��BH���Ч!gx+���ؖ_�Up(�H��)Ѱ�m���+/��T�j�p���R��LԺ��N����U|���X|쬼�3���ͱg}�M�jfTͱdFׂ�A�xm�W��9|��|�~�1��U!�4��Q�LP¢,�.4��G��k�P6��s;����a�p���ϱ���ϛ}�p.>KЭ"�:G+��f����\ �B@�-��&;�fL���J�}��r�{3n�S�G�ê�_�w[���ҭ���h�������&ec�%�h��U�E�&���Y#��[�p`�j;L�'f[7�o{�W�9ܮ_lzHo���c�z�X��ΤT�����	�a�FFq�b����$�!9��a�u��ׯV�Zb��TX����7��n ��Vo�:�﹘�ZӤI�Hi�;�Fi�6�+U�狂���:`Gp5�tX.�Z8FX�Gr��f�A���J8���γ�H���o�iݼ�|֙���1W���`�aw��C�VPw�����إ�����m\u3�.&��Yu�=6�F�s6�����Kq�7�(
so+<�ҽ{f��P<' :�]<��k	-Kǝ�W5>�k��q_[;�nF�T�RAp�����(_8��Sf��q�|]�TSfQL��ݭK�(d��곲S��L��f[�T`|� .���w�Vl��'{�Ƕ�J�#�	+�#���{�|������ݡJ�Y��s�o��-YM�� :C9Y���UdG��E�B�8��j%���%�0C2�:��MFeqP��~ֈy���k�Y�Rr���&���Z�0�(���u�W�����^���\�̗c]l;J�����O刦��h5�:D:T���<�o���j�/�w�܂0V�#7b���7EaqzTe�VTX������@���=�����\�|��1�uw�g��x��H�@��+��LVif1�-�ۿ��B��;]�<��q/�����7���^Y���VQ��TI�fz%y����ı}������J��-�ǏX��[SCaA��'T�`}B�|&<����W���i�Z{i�-j�Bʃ[7մ�g5� ,5!�iFҽGT�!�3P��&�d[�ZgN,�%_��7�ˤ4��W>{w7�gZ��S�P�D�������Z{c��H�T�"�-��}�g���{�8��Do��5#��9�|�y"v�-�4lZ�u�|�z6h����Y��Ǎl��:�(��^�[oF]��⽴ssL[�n��Y) �|kYŝ�e��Pc��s�r�P��i�Wvn'����^bw(�����8vq��I$�;S�)���|9T�A!X�.� ;�WP��E&kp٠�R���9-ۧ3�5;��Q���2�	�$�G��
�*�4��sDhʾTÚ�ک2�2�'��R�8V,�v��[��\8G��c	����Z������|�-� vz���Y����x�+����`��[��e��@\�ўU�ā�)��H�*�ڽ����\�Up^=.tڇ4��DRR�)�u�p��N ���n�Sj��H�˄��%�Y"�;j�C�9��_NEW,k9!ĆN�|pX/�y#=�/�`1�"r�K�=�:ȆG��9Θ�M	ʯ��w�z�r�;вcx�~��q���z��D��Z��c���ck�q��W�x�|�9����(���[��`�|Oy�p5�e�du�~���̭<<J_���#�]�j�k�{}Q״{����k��J��� kM�����.��AR�G�d�̭2�w>������VSW@MaZ&�i툫�^�ux��DX��\H4hx���4r:�q�W�x�L���C�y~�-���E��C���ɳl�u�ճ�{���P�����
d�E�6v8�n��ߺ'+3�{�T�s��Nb�Iޅ!%H�#��slEHL]ۅK��v6^����KOA�y��1�c�ُ$�ɍ��V��~����P�ZI�V&�J�F�;@���ev ���|~�u[���;6�ʓ�d�� �[A_T���:���E��Vn->�ȱ,0e�֕]�~f��
h�������u ��կ<B]�F̽R0uU.s�C���Ϟtl?wPL�;�3��x��3��"���Y]�~C�6B�L��'�=�M}���,uKe������T����s*:9����;���!�"�PO�:�'5X����d�8�/�DR�� ���T�o+�V`yA�z�����	��˂AP}|�Mэ���R��I�JW�z>���@����TU�E�8�C)�PL2�`_��t��I�p�R{��V~�_:�{���!��}8,�"�8��:;��H�SvÓj��F|������J�5ƛ�S�U�SX�[H�8=fyi�l�[��<��Q��gcp'Cb�ˀj^ݢ;�+�sIR7r�:�[\�jQc:`���
�D�.#CqY�pM��N.�~Ub��o�������Ek�,�{[̝�m��y��G�^��\m��6A��y��Xi������
+���[kӚ���=: �τ�}y�����=���03��[�t���0zm	(�w�g�ǔ���:�+��l(��S�R*���2CWc���;�&4�p��%��Q�ٽ"���J6sd��$B2N�����"D��	
��.m�^�����M{��*�w[xU�vvtQ�#c�����j�[���S
�N���Lr���s�Z%_�o$FP��F��hN�Xn&V#S��m|b��q^�����e�����7�u;u�4rߗ���du{���Va��;�ۭY�*�E/tu�E}30��N������} V��y�1�#��="�X�F�{6�X-*+�t�g���7���'֬���T�>>\�7*�<oG	ͺ�3U{|���o�-v7$���~Jx�YF��wo}O���u�Uٮt�xg�����/K��UW"�mε2��H�S�j��ys޿4oϞ����1��I�fzE�tW3�aC�{mWP7S�C=M�C����He(�t��US�����/��Va�b�L6htky��>�6e�ñ��ʝ���T]��@bT"�1�!T7�JvD��l�jf�Qs:��$;�|z&K��5��у�o1qx�o�uKc�u]Vh�j���ZE=��w3�+����N����q���v�;�J�lu,@�{�1��L��xeJ�9�����%qZA�н���8������v��I.e��&5�2H�Ѻ�Q�r^�00$��7 �_:�ΤT���ϔ/I��Pe;�3,���a N�ن��5�2I���$g�i,z�ZS�K�[�����OU����ۺW˩W�[U����רd��Q��`BVd!%$���WM���"��e��]�1�e���i>���%��J�>�9�_VK���+��ݩ���ޠk�C_0�߲��Q��\va����9�۞�yf�9C�Ç}��9�p�VIRW����l��L��l]�p6�+���o���^d�/
��Q�5(#�)"���V3����&�&c��TX�56�j�&T����3�Ó�u�Z����(�G�'*bB��'Vћa`H���r�=/��]���>#�x�Z����%F޺�w�Y��-�94�!�2���&�0�i�`ˏ�����Q�{E��H��b���-gԻ7��(��?w;1�n�,kj�/ �n1���]����(}���)^�.��+h]��R*&�ef��(�x\����ct�k"W�h:�m�w&<mn<E�L#�C��ĵ��]uZ۬*��"7�Z����h�T*�ZV���{�h{���e�E�&*�Z�t+�F����P��Ȩgͼ�'�3g��ީS�����v�X��r�\r�l��!]�_,6�!��>+��٭P˧��g�U*�R�*�kmꜻs7�X��ҽ��{2��8/�lTW��t^]N1��H����%Z��|��z��@�"��6�b��q|���|�*U2��t`Zi�\GZ�^K��m��K���F��>Flkr,��Kǥq��
d����%sS�gU���].��U�^5h�Rq�����ݶ%iS�kMm��e��{��f�jnM�0���ފ�8�;Q ������5��=m�oJÊt�"��s���G�����y��\]�m�50��	D�ݫ�9�姷Wv�%L�^�,˹S�ǹ��c�};��t��uz�:�q ×}�*Fk��.�KL���N���FAJnA���7Q�s7��z����*�I�޼�^:b7�>��GC���e�݌��W�S�o�vզ�#}RP]�:�\�GfgF&.�x��f=Ѽ��$��v���άk4ޜ2��̥#?X���--	�l��\�Β�ӱ���v���̕bl�N�4��G+�3F��Ұ����q�P(���� v����YVe��{��*�B�Nܩ�^9�vV>��@�R���)�r����]�Ԁ"�{�o���oqD�[׽}��jE=�.���6�5K�������PC{)�ko�i�[Y5�&g慴g��3U�z�V�a��Xu���o4'���O_f�z�V�����^PǋCF��{Yٌ��@|�h��t]�W2h��Y�' T� U����H��;��3X�������v%�l�/��Nj���������25�2�E��{>B���Eχ\V�m\t� �㽎�̗3w�ѝ���`i����^z̛a�&Ձ�iU�K��8�!ӥ��~ ف�w����@LҟQ��'�]��i]�n�mMT��Y�j(W�cu�s�P�Ƀo2�M�"��O�E���_>��:�_ui���t�V�����.���>
��fo!Y����2j-��f�$v�X]��e=�m�*ńۖ�+���9����pmr�s��IsS�ܾ���՗5#.�F��AwY��'/~n�ì�}hP�^�wJF�hT:@�fTW�ֽ ������9���o��P�E�j��8	�AY0�7M��׫��%�i���1R�u���ӭ�����������r=I��L<�ۖk g�0{�v��v��;lt��3XtU�uxo�R� *G�$N��l����}p⮍vThQk@�#�d�(st^'^0n��J��&Lcp�������-�T��vu7Yέ�N�q��Hҭ��9_rZ�H�b'�z�_9e�"���\�Ea�N^�YZ����8q��5��@� P4jڢeJR�b�Qh�[K3GU�[J�U�Ե�R�Pm�32T������5e���[kJ�-�%�F����mUF��Z�(�F���R�m�E�m��jҶ�"[+-�KB����Z�R�����*�e�-�mib(5��-Q�mmkm�kq�֋
��։Z6��*,D�Z�X0��Z��(e�-cK[kk)Z�m���ˌŶңkeiF�2`�8Q�j[V�[,A����UJ*��(Q-�m
�XUs&a�Fն�4�lʃQ�\�2�Q��j����m+[EU�[j��R��ԩZV��h+�1pKKRe�̶��c)F�PQ��b�ơm*��DRؘ�e�m�̠�[iZ�����W)qXZ1�UKJ	B�լ�JZ�&R�-�	kKmc-�mKlmke��UJ�ִR�h�R����4Q[ke�%�Z%ee��t.���<�e���I2v����Ϻ%pJ}`V�͹OR��u�8a
ǅ�+%d���[z�� �bɔE�)�1�G�L�y�c��y���~����Kίkkobp5D��;g`P���Ry����͡��\���؆{�1:�u��B(�ȷ�T=�hY��1�r?�u�Z>�q��=�?t�ɾ�(���<"a�G���8T�!�y��a7c!�Xg
�����a�IsTե���.�eӔ������z����0�]6�:��Fq�	t��U<ܜ.�-��u��@2ߒT�{e�!�ۚ�W ;�WP�Φ�|��_IIn��	�Ju�W˹�U��=*�f��:,��y��Y�9�8�͸{�]3����v��Z���}{ټ��-W��i��9��:J����"@7�z�e2�׆�k�YJ�|+c�ݛ�Dd�yB���g��­�(C�H�lN��ux��B��⬴�[6�ŵ2���pR&H�dxE�[��&-���y.Xv�ݑ�J�_H2n�'���nG/o;�U��fǝ��ZGk����Ƒ��J�3\u�	��W@�X��cm�Mᙐc�r���vT7�ӏ��ɛ��&�R��c��q�ү����9��w�i%�K v���@d���]����d�8�O+7����h���EC�^
��#4�@�2�`,}��9�Rc��RcS��Gȩ�����'Ӝq����&7��܂��eM�:�mT�D�oJԦ���noo�:n�Q�|�wS�ViB��郪�e�ڱF�ۤ#�nQ�����|�3�߽����F�z������]Έ�{pܣ9�o_;*pzh���t��_��ֹДm]K��ǘ�v��[wֺ&U�C�)��&�������9`Z�:^�.b�}l�����M}����A>��1�1n��~��%CW�\�XB���Q����G�
)���zZ���8�(�s�@\��WymG�!��{}5�Bz:;�yr;�
Ϝ�a�k��k�+%00��N�t&n+M��%������s�ƶ�����\3+��r{��sW�Ocԥ�Hz�\�b�'�,5���N� =��|��]�9��)9{2�Ʉ���9zC�{����2Q��=��ߺ�J�
zA�]�RsU��C����^x����r����&����Cdړ�>�_}�}W x:�T)Q|@f��)=�SдZ��z��{P�[���w��J��+��@�/m�̼��n�^<�r�|;�8q��=h�VY���h]��ĭ�����-e�M��S-^˵�P��8;���4W*����"l�����-q��(�լiƍ̓v���U�!�eժR�4R���wbfL `(m�<C���tQ~�B�Ұ�2�`^19�	P�71���Ga��޳�Ll��ԗZD#�i{c�gk��p�}��;�>�d�*n�w��wz3�k��ǫ}�]�C�ns���ʟ'���ȃ�Ň�߻:�&�۵@��m+��g����<\\�Nw\�J�����h��3�։����T~�}6��8elO0jr�o_Lk��X��tUmVǘ*n!`s�O���)�8Q�z��XN�����-���9rq�-�c��n��T+�vf�lВ�B*��L���Ʊ�����}���Q�m���-�Y����dK�bW�=v՝=5#���ʰ��2�����Ŷ
��3B�OI�8��~21��E�Iam�n~��#�b���{u�ѿv��@�Ҩ��5dJ�T�{Ѱϗd�ǻ������E��>��"��O!c��t^�F��Dm�m	��\+���4ʎ�Nǽ{��wi#^��u�v]#�P�ʊ�|f�Ui�ͱg���ÂY\6�}h^y�_]�6�ޒV�ц��ln5�:�r�nolS�
xN�Q�aZ�u�B^.�.Q��Y:��Z�����z�wNe���1N�4S�J��f�ް-l���&;^��#��,���C��(�B�_=���Є��ΧQ̜�n�Mlg��x���}r$�r�΀�T���5����U�E�>��Y���*��5����Ie�j�ړ�>(>u�`=ݹ��Ti;^fxU�N��p,-���QD�Z�6y�w�6<��/�ձ`ꪆ�����~�j��a���<v��o��UXs�s:��m* �~��g��\hg*����z��d�dK��V	�̢���H�98��s8D����w��њ��X:SHV��wr�����J�����}-�I��b���L^��X:ï�����yA��$k���ʽP����7��}M����ë�׃.�X��H�T/����W�ݛ����hB2kV��A�*���� /��q�4�p�2��uZ��&��-��i� A�a{���oI޼��
��G񊾸�=�S]���!���WةvXQ�q%{��G՝B�{��(�T9��rٷ6�+$��+�#$��{������_����r~�ݗ��/U����F�xX��&�\�b�h2��RUdG��֙���U������]�.�o��:Kvh��;���/x��:m��@N�2�u�6ØƊD䗎�)�+���I�v��ʦk���9w_BY�P�S�5�I���N뭆��X������*�1C�/��tv��Y1��uR�]5J��s�k�Q�V=Q���I,����a�'t�;)��`,�b��)��,ChȽ.Hȋ�AꞚB�Kp��>��kV�j=�F���=��9��X������?�]e=(d���)�n��&oo�0��o�ւ9:��X��7e��+u��	��4}u�������n��從���$:�����	��rñ:����#dm��|���Pت�]��#��wv���b�����O�_}�1�w��[{Ԓo������EX'Y6bl���[�wa��|��W�=BX�t!�L�賥T=�m3�c��y_=�s[�9^�ɗV�zl�TvS�^�L�C��A1ꗨ�SH��Q֛��a�3�V�L��������-�'��..�YWꝥ��s$mKޠp-=���䏄�Y|��m����l���wհ�c6TQ�:.$�{�pt���T��+������[�)0���s���ߦ��j��j��W���adQ%�y��m�Lq��n�h��*�r�re^�O]l�/	�Aۛ�W��g \��#��u���{gj.�N�1�%a�`9�݂)t�
���,�˽������lfswmK�f6�I�Iy�֕�+N9a.;9��x��}�S1�[¬�M��C���v/s�2��.o��Z��;%�U�xd\���K�#nC�!�+�B�{)��N��d�%@��o��9H�h�`���#%u���b4B�U='z���l�s�jڠb�=4���:K���"�@�J��_����K��D:��a�f]ۏ���k�N@zq9�7�v�M�_]Ǖ���x�-ȫ�i��o���N�,��is;@������	r:�.m�м%,�����c����2��x�Ӣ�Hβ��q�F�2�ԏPZ}�籁��K6~Sl����NP~�F��)�d�ܛ���B�3
�H4{��+���/���K7����E�pɚ�t�)�=/�刿5Z�\���kM�k�1]."t#�;�g��Y�x���/b�>.Д'���Dʌq%xt�&j
�ɯu:��GV�2� �9�6M������#LT���_��u)��o�C`OUCVzIrua
���tS�����l����H�>�=�G���s
��V:������ɮ�=*ȞJ1S�Yuޝ�Mj���C�]������*�x�"H�K8)@��I�r������N����RN���	�Օvձ6�/�,�A��艙l���v�WL�b8��	{��Y��x�q��{�_e9�3Y��.fٜ���]�u�v�8*b�n(^��V�˽���Ibsk}x���d|�N�\�U���g*�m��l��T �Ў]cm��^zz�a���3O�M~+���0�B��-�q�1�&m�˼8�<�굛�t��0w�%�)�1
�T�)��f��#�jژ�r"�(��S��
(@Q��1զ��N����b�W�On��h��Ԑ=�[���P��*��pH*<+�[U}��Ԣ3x��7+�ؙ��e�PQ�.**�QDM�T!�	�a���1��=bT($�LδF�R��չ�Ԙ�\ ���*\�x-Y���\9�(C��#EM�ď��C�A��ua��<9q�Q��]k�w���C��c�����F�'���t6'p��|Ʒ6���2�~k�z���{w�t��Wt(�ev"h/>"�Cr�����5iYB�,�O%�OV�i=Y��22��ۏXͲ/Ý�|�H�)0"|Q�����tUF��u'qս}��c	g�4�t#�6:(١%P�X\�6�2���Gk�����z��g^O^�ޠ�h�:ɺ_v�\��l�����Z��Ȣ++owPX��ܝo��xn��v�U��ox������Í��%K�(��[�)gQޖ�u�;�r�A�3�n*{۸Wf���y�K�;	��ZL�]�B�d����{Û�N���G�߅�Ef�%�]�c㧢FE	3�>�X���Ϡ�{��9D�n�cl{���ژc���nz�#��E�{�T7]����Va��'uSv�"�Vcf��͊��{�=Z��{���I��9Jq��t��Up7�xF��N��H�K�+����������彖De*3�fH~0Q�7f�G��Q�����u���9�2!�]=�7U��Է���j�`oMC����}�U�T"6��0�^���~�̘��DR�ͬ�ْ�|���l^�rUS�:����w捇β�T�B� ��1���߂�C�<�ZIn;��uu�svc�d��\I�Ǳsn3P6���Z�['p,�����#��<�1��]��;7{��^�k�X���hb��f�C
��PȲS�%���Y#���c.��f���x}R���;j�*vv�|v�6F��vG_ײ��Ԋ���94�4�֍3"�.���5]���L�q.W�GF��X^�-.�|�7~x%��ߋ��ҷD�s�}�u�]\��"ͫ�:{�(�̙-�{P�� �u���J���M4���W����ĸ�e�zuL��JC���,8b����qՆ�"������0��+�+�̊�1���u
솄�;Y�l	��\�Td����:��{��^��a�ʇ�Ϩ8����9�{���
Ij>���ŖG��b�#���Apڝ�׈�+�8l�;��W�:�f�^�����b�q�{�0u0�ڽ�y^�wB{���m��c��1U��B��%n��j�8p��rٿ�۸q+$�������'lQ9�)�v̮�I�;ɇ>o6=�d�,^:��&��s���e�#B���ȏ[&5����O�lz�!t�{#g�̐�����dl�M	��"��L�Fv�1@oJd���b)�hf'=Q[��P���IV򥳍h�������k�T�z�������2��/���s�(&O%���U��C��4�\�ea'�]}�LR�vg��Y�x[�N��a�W@�T��^��ة(c[��4W���	��e�s�;���6��Ar�Y9qw0��/�pnh���7�b�GB�3��/�!}�����O:�M���ƨ��x�^�y���0�37�����&]���,i�\K-��o|�fӡ�Ʀa�Y�J�{>�B�	�1�H�W�����N��JV�w�֖J�����:��V�P��`�3`������.��j�"����)�s[�����<���N��w=ceR��Am%1b�����*u ���s���q��GJi!7�dYeQ�v..��#��O,���h�O��{��7'sm�i-��B��S�zH��д�;N��D8�jrn����Z��X��[.޵��h�/ma;>���XzS^gD������oAB�"m]6���{��,Z��[�"b�5_G^W��%@��dq�ۚ����z�Zؾn����:��u��;Y7}�t��.�E@J���˫ǎ�0�4$q%G��if��P㍸{�o7��̞ɝ6�\���KTé�8�.��r��[���#ꑌ�W��К���3ޘ��ҹ�Jw͏}�<+Dmpk����s;}(as��C�_�lN��DDD𵜂�tifno$��@�S��R&Mw��un�\����=�݉�/��՛C:���{��,Y���2��@�+��'8����H�;P�C��X�sh�<˽F�<�n�_{�;׏�Ǯ�P2��i���W�n[��Y�G�->��)���v�'�,y^��-n�+��ݪ�܎�XeƗ&����=���E������"����u.��3V��.Uⶴ,��c@���+�@���A%�ڞ�X��ځ0��B�r�o)�z��n�2v7}EU3c���w���G���B��}P��_1;Gwg�t�sh4�g!lu���3P֥Y�{���U��P��:������ҭ���r��� ݵ(Ŋ�ݺQ�M���ń�bY���M���*���w�[X�pU  %
�����f�=Ed�9l�H`o��.�QF����^$j�Q�ק�:�j��;�l}��a&�w��Lk�(�Q���Z�ȝϖ%���Մ>�˴��%i��L)2�c׎�Jŷ�f���}�{�f�QQr�n�| �x�u�&��sj#�c��[-�E*�M [�Ýя���t���m.'x�b� ~-Tҳ��&�o0���GJ�EX>�ei�M-�A}���3�t�]r���Pa6;���G�[B��L��K��̙�F)����r�S9j�\�I՘OۋF<]A �sb[F���ܢ������Z����r|�˰�E&Gܛ���'����Ht+6Pb=�V8�H*�^�`���1ƺV0;k����R"�ŹWR[ޕ�4�*�����[����vU� �G�C�R&�\�G۵����ڧ�:1.ZY���=i<XwHՈqڔѴ�|��,j8o{-'Go[rrY���!��˨�,�*eV��ʄRk3�.�kR�IVW	�S��ҍ[Ƀi�L�.{�&�[��⭠+���z�mcpu�dԚ��xq9���(-8�o��+�,�]\��ަa���i�tn�RXP��u��M��]k�1O��@u���LOK�n���2n�;wc�v�𲸆�5{O���5�����	B'6�����K7Mi�JoU՗yl��KQwR�g�˙R*��9i�rb���c.	���d�`F��a�0 ��]�B�3�`�s��V�y#u����[}��ݱj�,o<�/��lL����[/1��W�&���jȜv���
�	�|�ٜ�W�ma|�C�:�>�U+|gP���o;� 0%v���k�p�i�B�郲𒾂�RǛ�D'n�\�rň�Y	zX�����SZ(+��u���7:co�b�zl�}��R_���YPᙪ��9*<�Ş_��P�3��C���
��&��ͬ�u-z�u5;C��L�<���ՊۅՍU;�Z�WҬ�!]Y�r3�X�:��܈֣ۭvT�2�&��Y�zxdU�v:-�G��8�w[����Ų�㣋�x��� �<���I��:x�1��2m���+Rxs����nʠ՘V.�QNWo��ڞCo�SYiV�M�:���Y=�+�̉ڧ6��ye�ՙ�<�]�U�b�8���|�Ǥů��y�:)oi�j�ZO�A���@���uR��
Xe����EDm,X�c\l��m�VT�-mj5lU�Qeb+b�*�ƴ�V*1k+XZ�E�-�Rլm�\�"�(��fahֱk����R�E�Q��h�6����j���A��6�3+��-
ĭF(ңQ�UkQ-��Z�V�Ym����¸��T�e�iX��-�l�+cT�[e�QAjR�,������jR��QJ�e����"��K��Ĩ��3Z�+h�V�+J���iB����Y�Yk)kKl.[���0T�����2�50�+�b�s"�LCe���"�X��LAűR��UJ�mr�D\k
�F�KmkVز�-EG0̃V��[m�ѩb�QQ���V�bE2ʨ��J"�V���X�-��Tb"�+m�DF"��0̠�b��PdErƅbcD}ޒ��K߂1�x�5h�%:U�ҟ]=�b�~�hL�"6m���&#ک�f໵�c�I5�V�ȯpwTNg���W����j�7�븤�l~������4�BhN���o�X3�F��`�٦�s{6q�*�=Γ�[#���Phu}�K�/���eX�S��MMaZ5�Y��o�e����W����p�W�õ�E��,t�b֧���g������=������B�ā�K����c�2hÐt�;�*0�������4������L�QQsR�'f�������~�=i
�������W�뒲��W8����X�<C���s��8��������+�5��٩H�}���O�5��."���.������>N�˷q�R��R\^?{��a�v�wj���:����#�jژ���P'����S�8��E���N��u��;��?�����Q�L�Gw�;��g�,�w��K�X~���C�&M���*�����d���2��-�(�8���E8�C<�Vy�[�¶�f������;{�@���!�G���M�ǟVuwT7�!�^����e&oi@����b�e�z{n���ݎ�� �ɸ���eP���$R}D�x,���Q�ު����Cp�֡Ռ2nEb3���U����;�J��D7h�nK;���2��jK�7Y���J{�#�Zޞ�Q,]���sRhk{nmM��,ʄ�ݺ,��������S��u�?oLi0(bb;�Z�{`��,}�q�P/�n� �$�˧�����	Qy�߫�">��!�xR����"P(��ay�������̗p_!0=fO_s�R�p����AIݸ�3L�hL���JL�ȟh=}�<��q�o���V���b��֒:�Z\
�렼�Y㢍��J����n��Ew2Y���^k���j�c+b��kĔ��*C�ʑ�/�s}vՃ��F��jw*�D���3�&����5�ٲ���e-�s�����b=�ck-U�V`�y������2��9�D�X)�����x$�93���6.����gʇ��l�S��{�F��\���S����s�B�r	�E�y�n��0U��N�b����B!n��5ء�y��y�=K`0s"2�
����'ݸ�t1�#�<k�*{�Y�g{�F���	���5�
�5�%��� �����	�}糭=cD:�G��Us8U{Zu��>u��N�%��c�7�����_!h1f)���e�D�Uy`lW��.��8�X�ͬ�ω�,��xӾ���x��-�!�e�<�b����8���/9qIײ�ۀ�l`p��ŉf�1�5��6�*ps6�n�1��h��z�6j��uh�F�
�	|<=�$��;��o?Qb1��"}"s��4�v_���ͺO���覬ê� �Y��� ���۞�����%�O�k5P"��E_f�_c�!U�PȣTG�@���|�)4�K��,�OŲl^�A��*�T����v�(���u��y/M�����h_�N���'�P�(_����r8�4ZK_��q�TϹ�����i݈&�m,�ٹ)䵶�ә�Zͯ|��n����׮���4�^s �XLp`0��X�������[�4t�o��Fʕ�.��ޝ�\�<��Q>��:שq��*��=֝(�:k�)m�(�&r�<��� U�;���GS�{�<��͟t�l�sn�I勞��F��`���
�Ջܻy�&�z���G�u�wN��%���5_˜�0�r��,ԕY�O,�bU�7�"y9P��}�/���>������sE~ֈy���k�FU��~OX�=�;�|Tq�6���F�k9��1kdxO� p�Z�.^�*�pɞx=+��,֭�;��L�Ӻ�t�@�z��D�VN'��Rf�o�fY��� :��@�C3�fj��Sy*T���nmAw�[��v�gZr�������A�H2�V�yЋ�qY��H���ܡFڷ���dk���Z,�YC�L���n,oaW�	������q�j��L�����P���i���"�c<�ч��Q�,�V�*1���ء\n����b�i�c]�.s% 򼦇N�MN�����h��|�ŵZ�q2`Nļ��U���
��.��^ڐ㿓?a�_TB�>�������� �W�gÕm��f�p�y�v�Hȩ)��F[�
��4_��8�r{w��{]{��}p�kL>z.�+�=��͝��Ej������2��-h	���ZA�m;�s�SH�&j|M�d��Po����ꔬ���=U 'Y�#a�יи�[�Z���(3��ʰVB|��Y�[�w��S��k�{�M�:oT��X��|��y��-�ƛsU� ;�Xq����������o�,���Zخ��T$h]]U��4���ډ/cA��C�C�[�E
���o����b�0{��L:��کW�ӧ��#�\8=�]��ݩ���W�Y�sT��ԣ��~�<C������./�ҙ��s�h[TP��-���J��D'X(��un��2�w#��� |�n_K�]��wuƏ%na]+��U���2�ӊ"֡�#yw�M6����v)��]��-/n��1�S!�w�%��L��y�j3t=�)*���}:�]щG�[e�f+���^�QW���57u�/�  �s}Ա5��" W� q��"��9�F#{]��=�uj�O.�1nK�i���u�Ng�4��zf��L|+�! �{&K��B#�}���U��Gk�ӥ�~�w^�������R�yvp��׏em�3ol{:Ȇ)��44�u�O�+�E�7-�C����x���v�_u�M��My��3/eD���T.D� ��\j�:Hu���ޠ�=��,jVS����3��>Gvs���q@>�W��I��P��#�|���:�H��Et\8F(i\ó;�J����j����
�q׬���Ϋ3�
����uĔ���L�!�^4��y�WV,��r_�N��+5�|��Aί4(�6v+t�r֧��Cs�P�Ǥ��A���f7���7����R�5е�Y�{�Ta;{ [�:���t��f�CA�����d��"�Ery��Y"��6M��JQ�[�xc��v}���X==jgІ��C'�)��>��{!����Y����>���`���� �����,5��
��o"�>�A��,ah(��=Q?b���+�&J��G|d�w�#���o�k|���B�8�A7�gJ��)��n������-�Ulu�H������ɛ���-73N�|��󣇷*Q��{�64��aP����v0�	)�f<}�ŧ��=X7D��l������{��w8Ž��k��Nq��LlB���gҪϯ�5a�}��gs��!�
�@����s|��Hy�L�kz�=rb��(�cgM{�Mf�"�uL}����;7 X'�=`�ua���ʷ\����
�:`��4�F������%<1P�SJ�qӐ�<�duUn.��[X�<\
��OGA%��l4�D�b���c�VuwT7��}圉��$����n�����ŀz3䈯�Ou������_lU��y{��W�7�����Ұy3�@C��z��C��B���!�xR��FA�D�V� �@�z(GV�]w9�֞�wv���~��EF�̽����q� �q�R�bGiI��ɥ�eM����v7�j]���d*�$@YSd��ip7�ҧXe�l��UE���w��V$˩x�O[/Ky��\嗞���^�ۃNV]Ed,uf��:z$jG	5;�dXf`���:b2�an�֭^��:�;({�k�8'�j�:�0W=�wF�etn1�9�SQJp���_�Ӊ�'�o-d���-Rx�t���+b��j�w����AV���J|�>�#ڷ�ݚ�;��26�-s8���&�r�]}�LfO7�u˽lĜ��>��iݭ՘*h�����r����շ��f7�_ `s�G�磌��(ww��]���f�q����mz�7����Cj��H�o`;h�Vf����\tx��7����mYG�ShW�YB�X�b�X|쬼�N��
�����&nvgS��[n�^�c�&�2��ŝ3��V'P'��f�S;1i�'��d��a���������r����x*����N�ѷΰJ�fD2���q��bi{���.�{�{M���U/�� >�������37���j������z��p��M�Zn�T�`%��!q� p;��TU��."��C"�NȘȗ�(Úp$6{�s�� (D2���=b��m��3������W�v�)Ԝx�["�d��<O�M�h��m�N&��J��85�+��ʾ���{�g�g�k����g`(,�*��i�C�3Z�=a�c�y�kP�c>C��c��&%~�a�%aSV�O�1�|7���y��ݚCH)���vAH���kܼŷ�'�;���y�|���,�q��}耨��+�{��I+8�N�g�
���,7;ߵ�:� �����ϓ���M5�J����i �H���A���T����L�,��&��s[ַ뷹�7}���^vT�&Я��ى6�H6��d��
E���C���O�3�{��6�R��<�0��I�+�����c�g{q"2W��>;��VF�8��ˤ���|�������_,�.�D��E(4�}��3H�`����xh�uג�ŲLd��©�Rw��F�|�����U�L�l�>�5�N�jq*j0J�3���9r^����b��`�xO \ky����N����3Q$@���7wXsz�����{����+/�����I@����l>t��B�n�b��~a��I�T��޾é<~a����CO��&=eC��*�Y�%�w��M�i+?�ړ�/X'�3�J�Uq�L�Y �5�녝�DY[�{��o��R)R|��ٖ2�W�Դ;��H.�b�S��a���
�ϙS��
��Y����6ŝa�c'�9�OX|�3��/�8�'��������G��)����/������7�a�q��/�0�%~Ձ���i
��{�x[&�R,��Zq5����L@�?e��W�X���r~��i�AM���1+a���8é�1�LN���}~����}��;�zϵ�s�~���΁�E*�~�Ci�'�9�LA���T��oRz���ɉ��m6��R��I�T?S?�=t���k �i:���{�I�%0��N���
����f|~7�o���KꉼW��q�����~�q�d	�� c�ɤ���I�s��β6��w��&���>׉5��$��OALB��,�i���b)4� �Y�L|a���ɏ�Lz���y�5���}]2~ߊl�� �c�<>En�1�_w2y���Y�>��6����;��R)Ěy�g�����y�I��Ă��&�Xi4�C��3%|`T|�qP�1 ���K3�����Y�Nd��;���������1�m����1��_Y����g��bE�Y���a�O���}�?��*J���t�}��6�AH���ځ��5���z�r���=;��bf_{`'?�󜗿V�M��ԥ�Tlx����1���=��x���Y1��0�cg��UH/����~Ci�j�� �~�5��u���d�y���N�^'���ԊO���cIn`\���6�We^m%���q�i�
�L@�*c'�=�X|ɴ%}b����Iύ�i��i���AH��~LOP+8���8�LH.$��u�Oܡ��oZ�AN�0/����#�rޟ�^=���P4��'}�uI�T��O�&:a���膟�Ę�<-Ċ�Y�7-՟�1�M�u�y~`W��q%d���Rb
E:��S珉G�}b��xy��)_e%p6yL�ހ��8�+(�
[R�<������r�M�ly�y��YL,=���Kw8ѻ�.P'A��$�����rYRF�`����5{@�����R��9�iA�����,���0��J���o,#����ǟ����}TZ���w<��Ïz����Q�ے ����q4���tM��*<9�jT=C�ć�{�N�X�~LOy�i�C���!�����S�P8��Y0�u����8�B��9au����n����yo{���@ ��dL{������0�
��!Y����q9�Nk�~`T�g��ki?!^0*z~���ϒ��l1�a��1?�4�_���S�6�^'������n�}ݽ�w�w|���B���+f&2q���a��@�T�B���i�I�+6}�i�̞�AO~��J�d�g>�3�J�įs����C���CO�LLx�ܱAH��x��^7��f�p��?\��no�}�<"=1�A ���i ��B�뤝��2y�1�\AN�|����Y��a���Ĭ<��COԘ������Ak=I�<�56�@Ĭܽ��3vq�g��ɒ;Pq��wj�~Z��.<�ޙ. �A*+%W�̀��S��C���*+����L۸�~a��4��Rc�����4��?&2p�d�=B�gX~L�9�����1����is?M���r�-��9�� �V�ĩ/|ь+
���Ȧ!RW���I��
��-� ��g�L�HT�n����~��Y�4����y�_q
����������V�]������Xz�6�;��g�8��Ü�S��A2gs!�uH?gu�E�A�Jǖ�Ɍ��,P�
�'���%dRbԶ����7�@�T��ww������.�Q?{cc����$�Ǽ�K�M��P��&&=g��H)���14�Y�ON�[ܟ��$��i;���d4�AN'�������̜O�6�M%c~�e�>�˙������G>��Ly@�Ï�9 �z����2�P:����|ɿ,�&!�فĬ�&e�M�w&�u
��gy�.0*
E4�������<�y�������<5̚|`Wu8�s����bp��i��q���*<�}G�*C��n���:�~�����������^&�߲uĩ�}�&�V:�'�w��RW4s��T*�0���1}�"5�G��󦖛��B��G��x_)�a�'���{N��=�����5q�ڗ��L�R���VE&�m��q���]Q�)�V��8娘vz}y���'+�;A�H,���ya�و�j\rc�]ݴ�B���#B�H�Lv�`���W�~���m�oq���{c�a��X��3l���u>�{�3O�
�3��~B����4��ưY�]��g�:�͞�l�6�^!�}�I�u?!�O�a��T�W����Q�}1�߯���Z�u}x��o^}� T�;���m�+"���f��2x��Y�J�"���%d�W���N�? {���B��bc����)�����6�Y�<>�Mn���bA���������%���g~���UZ���1���I�hq<���6��T��+?'��M%|;܁��1&?��O��At���4�eH�q�5t�.��ɉ��8�gY3/���q
��]��qs1�ߞƕ��vg!l8�L
���������AOy��&޲}�i��/r�^��y����J�`_N���?2��~Lg���,�
Ŝf���A|a�xZi�g�1 �`��� � ��@i�Ն؄���s�z������gC�
§Y�hm�T+On���ĕ
��s$_�`b�7�i�a���=;��g���y���OY_�<����|��HW�=��!��<�H,��<�{z���y��u�o~w�~��aY��A}N��bi'PĞM���*(n{M i+'Y]�O�d�J��~ÈmĬ�L���m �x���6��@�T�s_jO_�%`��&>�i1�N_��}��<׏�޼�sϿv~I��LN�Y�AH�P��bAg���O��>�1�I�P�l
�g�n'P�J�g�a��18�I��]$��1���^ �G�~�O��~����׽'�R,���)�z�r�$�k�P8��əx�j���!R�V�+���RاRq㤃���&��>�4�O,�����nj�8�!ԕ�����m#�G� �c8*K����\�������}�`xʅb������ �a���h<g����~�i�?!��R.�;�)��N<|�I���Y�ُ?X��e���~큈��g�	���|*=�������'�Jh�׿Oz�'��9��@l��1���L�l{������&�X~k;�:� �~�h��bA{�rE4�'P�9�p�jE��ݡ�+'ɫq��Ɉ*o(~CO�(0�?o��_��^_�G�OQ5��.׫F��V�J��h'���� ��`ü�$:BCe��ٚ��J����Vl����w�8s�|�!#u8�U��=�9I��uN�ޝ�)���谱,q�ֆ��g&�T��+t�c���or�����X䷲�-׶��n͎nZ-\zhӡL��V�u-A𳣫�낇*۬oi�q����vJ}��ˢ��'D�r�2� t�r��5��p��3褚��IDi6�6\�����5��TN>�)�|�S�Pl�>���i�sY�,,Z���X;�����NlՋ66�7��$0�>��7���)c��v]�e�+�y�	�e<�3hM2�/Vڕnh��	�<^�f6���e\��&�!���Y�B����s���Y?*4��̬��yWwPRU���@�;w�+�{��ʒ�&�2b8���y�rHM���]4�|�pe�/�
>ۛ���y��A܇�z��s�a!������zc����a�Ԃw�$�,�R�mr��TNwK����ͼ�gmlU�{CC
e�=b�&75H�&뻹�d^��];3n�3�V�ָ'7��!�b��쏡ݾ����z��uNz��)]�+]&�zr�R����-]ϐ�;����铬����>�\D��F��zJ$r�/)��L�٩����t�f�j�&V�-��wk�T�^�(JI�����-�}�0*R���u��u	Ev�V]����ùc~ݾ)�����d|�Y��2r�٨3@�:��]/0Y���H�J�ܧ1pB��K��!Y�7yK\��{[�)G�^��3��u� J�v�]�}&����M�o�Wx��K356�9�XjQ)Ki;m_l� s{'#iSx��h����V��@�ɝS�{C�	,a�uJ痺�,��Ŷ��(]�5,�g�bR=��)����y���vV�\�
�]1�/�����t5�ކ�sv�v�j���C���=CFQw0��&m�2��cx��� ���g�$�D@��[�R�8(v|���ނU�õv�<M�jL�ھ)����lݺv��2ݓ��3"E[�R�U�<����V�CQH>��>����s�S�k�:ʼf ��z�Sʁ�]���܄]B�L�zƳ��s�il�x���{}����2(��^�P{nm�oJT��j�˨�ήY�C	G�z�6,�ν�z^)���<��v��6��ť�&��k�u�\8�z������a�w�f��]��BN"�1A�nJY��*�X��h�J�=+c�$V��5�W&�M]#��;�i��m�̐�gZK�sxw_�9���N�m�q�Y78���(����:	/a;�v��d�{-T��.�(׷���_fp���\˅�Z�w�>����ޚV�=6c�闚&'LSyR���؄tM��!_|nv��q�~h��3��8"��DP丮�c��N6����$����2=Ô/iv���x�D"K(�I���d$��KF��E���UA�Z
%,U�J�e�PkJ�F�����W�TTX���[k
�f5�љB�YV��ʅF�%B�jѪ�h�(bUCb`�\J"�*��"V�DVT* ����e��m�Z�Z�%J�Jʒ�1�Qh�B��FV�hU�(�*ʗbTQU�VKj�Z��ʅj4�H����B�k�J��0E�[�b���"�j*
�J��֢�*Q��EV�T`���eX�T��[Em��*���*JȢ����U�dTAbZV
+l�Uem�j-��R*�[Y((�`�J��P,����U,\b�mAE)
�T��ij�Z�IJ�KB���Z�meQm�Ub���VZ�X6�O�&��c��a�
��M<��/��4�s���ݻ�^�΀F^q����_.:��y��)�uj��o
QO�xx{�jw2덤���D `xD(q����AH�q5>��u���%Ofs	�m����P�s ��
�ɳ��G�X#�gsRx�1 ��皑ݓ&$�;�> c�;�zZi ��GWV���ٿf��P& 0 � ���q�$��Ă�gl����!��>��LzʑCs��|�rΡ�ɴR����9�
�hT��ޤڽ`T��CI�N�t��6y���Y��7�����nRφǲ=��dWsc�z��|�&��J퇆�i�2������8�b��u�M$�߿a��4�$~�^0����{q�XV;�sXɴR�nV4����C�<���5m��c���s�W�l�
E��C;��ea�Ϭ��1�d�?3��VO̯����I8θ���偈,<k<JͥH,�=��M��6���}�4�J�� LI��}:�����ߵ��� ƒ,�:��H+'yϵ6�{d�
��)=B���MI�`x����{h~v��dї������%�����'S��LI�+�~�i���" ��~0��s�B��3�s���1m�1 �=�2;�u�c<��O�q&���l1 �_w��=B�bW���'��4�a�o���T��>f�f�Xz�07���LzʑOR8����l��������;�s�o�ϼ�>J�!�kW�
��/C�ѶM������i"�I��L=;�CL�%zɿ'sg���_������Ci+���2M�����7����Af���=a�bAx��S��s�y����ߟ���p*��|�!�t��èbbVn{f |��a�S��L@�T�}�6�oܰ1��7�Ch)�l��� �Y�L���3�Jώ��~O�Y4��G�ːtzb`{�m��T���I�����o������2�3�R>vC�Vg�ě�zȥC��<�v�^$YSԼ��*���m�vɌ���i'P�R�w3	�*A}zw����
E�?k��xs�{ϳ5�w5��y�����z�dӌ�|��=J�'���u����_S��M?0*
l�:�����gd��1��] u�=��r��X{�q�)�*?��m�Y��M����k�uö��C�;�k�dŃ��6��A��i�!#�0e��r�zu���w��
o*3�n`�wާհRa�V��X�ܔ�)@F�{��'2�vq0������2��+.�ە��G	|Ӂ���S4NтܧӰ�to�1�ێ����j�T�Ǣ)_� �ͪ�x�s̯���������wD����Oyܚzϒc�T�w�h�f2\��d��Y�yl5����i11����ʑN���L�,�J��^S��Ă��������:~�O^)�����Us�C�	��* �%w����eC��i�C�f�z������!��|�'���z��ĭaP>J§��O�1�uCc�X�3���Hf�ND�����]'��}ځ~ ��i�L��B�l�߽��쟙_���&�VqĜ�>�W�Aa���`��R��pXz�a��1y��Y�q8�e�H/)��}����Vuf�F���m]�]�|7�����c3q
����m
�u�������<��&'Y?8����r@�_̛�w�<z��4�|�~ԛLx����i"2W��6wL����}��{Y��jetO_U�u}����{���q�X~��Y�l:�?!Y6�bR�������%H/��I��!�>3�>����e�Ԭ���s�nu��%}���{ه����O{���}������~�T��^2t��6��J�玟2��VJ��~����?0�|�C�9��X�2���1 ����ɶ,��<�d��!��ue��A}a�1.�����;��t����Kj�;w����`z  ����z���ltI��s�B��u`g��HT��S��4��g�jӉ�ԅf�l5M |����+�,I�u�>?S�4����~�������﹜��{߿�z���{��|����c<LK�2)P��y��A}I���S}��7�oRz���ɉ�Ri4��R��l�B�~J�������8�N�z�=�ɈJ�����~��gh��/wW+�a@�q�(�3Q��\	v��N�ɤ���I�ns�M3���o��6�\@�>ͤ״1 ����=q1
�]�Oh��O�f i*A�7���Xz�1��y�w�;��3�5���~��>ֻ&�3i1�+�l1�Y������8����u��/�
�g>��6�����AH�i�;�z�YY+����i�At�;�&��4�M!�[ev��,�9to���?y����E�x�{��~ ��щb�r�C�.õW�7��	.6%3���gWE�`�
�wU�"�4d	����(����WIP�z�\	N�v㿚7��F^	������c�ˢX���ƛUe�:S�R�>Я\ys�<� <<j��wn��� �`L1�b�0�1��[��c=w�H/u��6�H�q+7�4�I��La���M�RW��='~�ěB��]o��� �Y�������!_Tz���p��k��ul��1v���>@2��vy���
�L��ɖ����Pw����,���z��La���H/���:���Ax����L�)*�0��eg��g;�i4������Y�}w��W��w�w�u���A=B����>��i�
�� z�1����2mI_Y�h~M?0*Ny�i��i��M� �FN�&&�gAgɉğ�N�I�(­�wʳ��m��Ὧ�%Rg�\AO�T���M�@�V|�Nw����@���~I��~C={�3c�Z�@�Vm�Z�?2b5LgY5��tÈbVJ��x�`z } aS2�������|7�P�x,�;���d��i �|9���:�M!�w�o�
��'3�J��|���֧P�Y�?&'7@ǌ1f'�x�������i*E�w���LW������%i����2��O7י�����%|�þ��M!PP��� �]��aS|�+4�RT'2��~ɧ������ki?!^0*{?fZ�g�Xw�ΰ���Ę�@$^^������^��.�������H/��7C��V՚M2~egܰ��@�T�!]��4Ȥ��}dƿ2x�<�� T��N��Xϙ*�C��R~O�*�F ����Á�7v$u\��;r�9�V���FM�ze�AgYMe����Aq�C�r�2y7f:@�)�/��i���a�a��x���1�:��?'��i��&=<�5 ����(���`/kv��������_~߽�9g������M3�&e�����T*VJ�73 ()�8�� ���ُ�O�M04ְ+�'ɤ���I��Avg0�6��|���s&���:��g>�}�&_{���wo������q��c;�<���Mw���T���1�aS2c��$SHT��lRbJ�AO-� ��\g�L�HT�7VL@�?e�Y�4�������e��w�����xE��X�U���'#V��T�B�ng�K�U��,���e>�cu޾��vh�@����'	��kZr�z>"rd�Re���:����ŵ)�$,ꀍ��v���y�����8:�v��7��ލ"�
���c�����<=ah�1ڭ9��8� �G��]jZ�g���L�xs�ju<H/�OMwZ6���1 �gu�E�CVl��i1�Y�Y塤
�'�R�JȤ�+�`/Ϭ�:CfkϝA��������$��=� ��>}��1��q�s+�����6}����LLz�e�Id��}�M�x��{��O�S����z�����<��CN�1ĜO-1IP?%�?q��߾��t^�c���ƶ�=I}�c��P{����gRc�� ����i��
�ԯ�S�MnͲb���Y�Lˤ��rm'P�Y7�oK�
�SS�~�1�� ����Co�N�da&~}������[�y���zHVO����&К2���!�&��ty�����lLf�'��q&�O{�̋'$�,�,�>�ے(��]��w�������o���\偌��ܚg�4��g9�g���̧�X|�?0+��g���$�vi��X,�.��!���S��m�&��/�bbOP��~�OR,�u%n�}�5��o^������}����޸��i�D�� �A5:>�1�#' ������6|@��y�~�&�cF�Fy�0�^�Z����|g��	U�0�=����J����a�R��;�,��ᖡ�w�ݨe�C�H����ьj��?|a�:�ٚ|f�X�C��]�-�%�c�e����]�ْ�R�c���+Ix��47�د�Ȥn�yMXt��v�;��U�������*��_���mD���Oڙ���������E�u�9l������	~��y��2<�W+��M6���^�ЗY��� �m�˼>�YA�guQ��u�t*@��Iۢ��z�V��i[z��L�x�<�j�L���a��qŲ�e�����2-���1~��=F{W�mPT{̽��\v�8�e� �����	�B.Դ&Y1�_}�}��T��$�׭��*N���?�O@�*�=����`��V(hн�\���*��dd�L�Q3��i�p�G�MW\}O
�ǊK��$�Q����x�/k쓽e���Oi�����NY�,��Hb�vù6�/Dq"*N�,wuq�?
��>ײ�iz:���J���bQ��ז�F�q������!Ps�|�	<)EyJ(�؉�f�ܯCl<��_]�oT�yQ�����;x��e����z�sl��V(�~nl��]�;[��d����ЂI��=�`���!��B+zV�vdL�Fsc�^�Z�qsS�_����;;'4��0sU�Ʊ��j�]�\*��W^�h��Gx�����C��=��r+=�}=g����Y�c���A���XU��]5�8'�j�?��\�3�20wz=S�=`��_�ܑ.��Ph#۬�7i�7buЛ���j=�l���ؖq�����)�&������r�kX�F�ͣVDD�V2X}�گ���/1W����aza���m]�W�M�Ӛ蚂+�D�={%e�3�F��:
Ӱ��w��a|��Ʊ�SK%�,L�=�~�/@��W�U>Wr���.�/H�L	h_Fe��:�r�]\�N�[٦�*��C�&�[��S�BF1�OW7�����`�;�nt��:P9�3�?{� kw/i*\�J˃�*7��qaUP��!��j[Ղ���Õ�t?/�\c���Z���r��㙧�5��O�T�	J:��o]��Ĭi���tf�31Ra)Xj��x��%�j9���k};;^�W��ϟyL��9�˒{��F�;vi7�o��<��]8ܩ��߰y�Jl�����O[�gw	jo��ǛӲ�VA�J�8�������@S����ZHQ�蜍��ޜ�r�/V$�+����scS��w�{:����C��T$���^��]���Y��x_��V�~.�%�llo���}F���M��1抭%�����y�"�}��E���=i���H1�،��	0`�K�4K����՜���G��jdr��H<�n:����{f0F�r���Գ��t��X�������ρ��>��S��M3%�Ŭ�<d����yP>F�/n:̯n��dcF���1*+��բ��'gy�~�
��YN���и��7�Jsݢ�!)�V�<�vM��s�bCK)���L���s_�L�ǲ S�F��0L�&�o:1��<��n:�J�  {�b�(��K^^uVI�Ô�B�-g��~`���o����3ǎ^� �ķ����=Tfo����E���X�Ć��y�8+��f8��'V�X���Ԫ˝�3���gv���}�;���l4�g�i�Ma2�}`D�v�ƚ6�����[V�SZ�����Y�^���×��SBCH�}d�gC�.�y3vz�o[���1�����39���^���~{>����r��W1�;���r�/dI��0���T.������u}G���gG������m�!8鼬ד2
�~gq���t=Ï�+[E����W��C���."g�KO'Un'�J��Φ̭��~��se�c�`�5姫v�]����f/We-�Bkf���l*mߜ�v��m��V�'�uA�I�8Cٺ�6�Kζ��r��zo�U�hZJ��䣯w8aڒrOb���/���<K�;J��1����s�MM�<��U�{S��5CJU���v�u��w��w��d1w�b+�c[%M';�o�1�P[@��e��Ty�a�Q�w^���-��u�=q�;E���X����O�b���4`i��7rU��H��6�������uӷ��sR}W�I}RZWG���t��S+cs���(6�d�2;'=70���狂�b���]!�BO'u]�=ڢ�4�m�7�R�)j<�L��ed���i��V��8�	�o:��hzݺ.�T9j����&��\��|�4p��?onժf�{N�+��7P8�
-������?hι����2��b���0�o����0�2��K��]*�1Q�7zra�s�Y�=]�E\��P��l5��nqŕl�=0����Q&���]}����p��+n������bfz�j{�����4n�Xi�ٸs�-sZ�I`�C᳀��X�n��YY6�ۮ��jk�$�.��H4/���g+K��ٮXL�mX���eʸ��6b}c���?.�_$Զ���m�܃<������i7-Ø�뚺�t��r��Y�.}m#���b�W�Fn�sS���7�.ѡ'S6��;3��΋(h=ܳ�Ƭ��]��x��%���7�!�soi5��Y|���Zaݦ5��C0��4�V��Z�*�^,ۊ�免�\8��P0\J��4��)����=�f��o^��)*��w/�>xKV����m���3��Fr��P?2��{'?H��>��\��Rȕ��ׁ;j�=�V���!Pg�7wk����W���wɓ�z%��z��&�Ռ|��ys6��nk5���N�]�b���)����;p|9�}�v�X]����$�)�MU,38�&����J��'����"	��^��Be�b�H���D��[��yW���Y+6��e
u�݄{1q�-(����C]A��ޙ���׃!`,b�\��ޤ�ݞ�2}O����cߒ�{��i��h�L5{y�9vv�U�RwA�n�v=�ov�n������C�o�ׄu��U]�Y�qF�RU��Ϻ�
����I��.m��BS�t��y����~��۞���A�*x�\ϧk�O��C�Ԛ�D�z�s����0.�C��P�S�>Ӻ��R��vD�B:r�u�.j����'em�k�-���5��.p(�S�ͧd���'u�@mJ��{6ݵ����-��ɗ��"Ж����q[�vGg6k����T�i�Y�ԁ��.#��K���k������u�qZ����Z�/��C�\�ք�0?A=ˁX�^.ø�ת��1X���'V�t���5ne��:z9Ѻ��*��Es��y�Se�A��-!��د�L�o�7dمSȋ��C�9�Sgw����R��k�|�Ӄgf)���^ӘV����qx��fs�%�>y��zɏ���C�'O����S	�ٛ�[��OwUK�rm��r�ÌGwT��	�C [����V>T����c�1��f��uc�ͦ�&䕭a��#Y+�j���V'��{�j�����,sq#�C���էU\-��:�>�C��\��.ns.zrk ^���;�̨���ni�v�%��n )�ʀ��S-%�S�Y{Fam����@ձY�Bۆ�I�&�g^!����C����>�n�[�Fm��n��2�J=d��N�@E`<��M�<fW?)rp�2B�N]ӽ�c��&�82")w|zJq;�
�� � U�[�Xp8����J���K�s�����*���>�����7��6j.��kjV�0{�%���
5���kT=���������NC�.[x��	}����7b���e��6�Pu�2�(��{X���Ը2[�#u����v��a�9$�bm�"�T�[ΔV�w!�'L�j�v8�jߡܷ���y�fp��ޚ�f�}[��~O��d��S��t4��n�R��NL�/+t�Ư��h-ηGH�c�I�&T� ��B�μ2��l��+��w�PٗS%v����7�P��7I�t���Ivj�"1�\�/�R=I�Yk7�6�Y�dik-v
��[�&��"�\�d�.�,�>U��=6�<j�ÁZI=
�3����c�3�
�f���}2�R�'ـ���ҋtk���OF�@�����ًq"]o�]���]�*�%�lx�,���L'���ׅ[������N�j,p�Ï��g_0�L̜��zE�`GF�C�`.��oT;�˵:�V��X�+{�aU�b�WAxѻ,(�����6�����L���0�i-*����]\��wtFC��GF�ƍ@��ɼ��p�kB�P��a{֮8�<��چ,l2���2�]F~��f�73^T!�\߰{�5������p��s/�ޡtQ���1p˵�|�J����z�Pv>vU��u=ر8K�LOk��.s*>��w�ԫ�*UN��)9H:�b�e��ڌޛ΃�H��(�Z��Y��V�ѕ҆�����{�r�4}~(<��w]Y(�2u$
]�\ZGu]_ݧ�M.���ކh���g\}I'�s\F=�'�x�΢1WB��9�K.b����1����]�i���%&�����І��8P�:r�=E�������)�{@Ae�{w�d����T�Y�\�@���t�Y�=�[Ԇ+VU�����d�|�������rR{�^�h9]��i��̧n���f��Z;�bf���iݼ��f�`�U�Zr�{���nh��wZ�Vd��N^-�oI7�':�ր�������'aUxz�y��M�x�J��Tk^v���07�$�Աk5-��iQ�R�E��͏��2v��W��7Tm���O��g��7u��N�9U�ݟlJԘ���.ܐn5mT�*ʮ�IS%�íb1tWI�9b�(w0ryj�V��\��2��wx���;���I����)�n��ɨ���K����(�np\S���::���obb��K<<�p�4�h�����Sn�4������_n]m�N-�~{�mS��Aj��S�H����z^O�m�Ⱥ��7)ə3yF�����5�	j��e%��Y� �a��VA��'�PF�/c����\�v�'�v+\��v�w�[g�X��PT���2�Ʋ�6�`�"�f5R
Ԩ���V,�UE����Ң�#m+%Jũ
�D*Q�kB�Ab�F�UUb�H*�E@#*Ub��Dm*��E�Q""�,��0������еJ�(�Q�*(��PU�VQ��c�"�¤��*#���mX� �Y1�LJ�E�1@�*���1�-�j	CchQTH�*D%eai`�F"�Ƥ�,��1���*,X(�%B��)-��9j���Tj�l,Pc�B�D%K�c��e��QdQJ$���V���������EU��D��(�UR"B�AKh����`,DU�TJ��P�UY+
�-(
���EX��F*�F
(�ֱ�Z��UV(�Qm��,`��X���T+QDTQKj��$TDQ���� ��  ���t��yq�w@�=#�R�߁җ�/u���a��\-WQNevV���e'z1�43�=g�Y��b$]p���/燀�6]��_ccct�[��R����ó/��O�w�}N񌎫^H]e�[�yRxJ|��n�(0d�d��R;�� �{��$�M�G�Ȫӫ�V����>=�.������	�jt$r��Q�uz�X<���82���yv�R�����*�7`@�!i�yk�P}7����o�P�7,Gq��'2�Qgr)�2� �l�
�(�	_�vai��t���Ii�<uT�f��Q;��i���\n�rpW���~j�Dx��7d�;��ok^�����W�c���a�&Ć���lg�XL�p��q��Of�s�����f���[�Ւ2io9�����M��}���/��W-Yϖ"y�͜�̐�˕q�s��]����_����g%�g'-=�󧗩�����a!;���=�����.�@[�]3�t+�q�f!��l���xS�/x��o�dx�4#���oo[���څ���k3P�V�H.ݒ"섦7�;�|�ج|� Z���p�$�8��.���k��U��c4�ԗws��n7yj��ݝ�qqBҘP�]黵;:��b^�����rW�*pޥ�.�s���jK�F���  �k�Ե�����4�X�癇-���x��T&�jP}^�
�w�U\ŵݼ����S�l)��2��{��;j�Wt �%�bsbQo^-�J�c�|��V�s��/�3ʛl�|���Y����s���]���O}r�I}�㴅�)�}�ۼ����M��ΨfW[ex�K�S��[=�7}w�Jʾ�pznI��G�Ι=E�͍���'vq�3�(J�����mC��y�4�r{ꮅ�Y������3�Ku�Ԣ�V�[�-��i�VҰ��uo�@�`��R9m�x_��/���n�4/��>�=��mr���[�h��p�B�ߛ�D,2V5s�0�V6�9�탏��Nz�ܐ��	�0�t��sn�Xf��J�l/pGK�o$NN�U�j�H�λ����x�o��ޚe� s�\��=Q,m��e{M��jbe7I�A�_<�����-*05��n'y+ ^��ÛBdL��연;ᴚ9]�|Uӻ��G���l�9%���,�FNŷu���d̩B�&Al��q܇�ns�ٕ�ʔ�U�z��r�|�r���}���J�wW}�| ��ە�;�����"7rJw�-e{*����דa�aޅ�%�|߱?l}�X�eƣjK��U�k0���[ڃ�I��fZ�ӓ7��Um�.����>�g��j�U��?d�%��I�νmf̭�:jq����b����\�y�|��6�"�3���NP��&�o�����SpQ� ������yuyL�ޗ�>��=w^y۳-�f��mYp�o�myf�\Jg����;�������V:ek��|�-�Ӷ�!H�x���m_4�hB�;(��F o��\�*m�sYC_g"sj:.oz��v����`e�D®�:�I}^��.o�es�����]` sV�;|=��N�z���c
�İ��n"aw����_t����=7���Z�g���/�x����w�{1q�-(�,E�H��	=�^zׯ��m�3��7Sc�C�k���p(ҳ�&���0pv�ҡ�x(�u>|�ZRhn�^�_A}��u�M�n2PM�.�΃�p�)'�3{!ɜ�:���n�rm�7�w�����sjj�[��I�X {�KU�ڴ>穻Æs���1@��y�����]ϳ����֞����O��}N�1��ߒ���X!QָH���ջ�hdo?HiU�����v=��{�-�4�V��������V�^�-�UksR�F��S���ٻ���L32�T�
;�ly�yc=|�X�ɞm������X�L��ܐ�\.��<�C^�n*�q~C˾��{���~��
�h�=��~`���7(��<�R7@�(+S͝��w�cH�܉`^!!$n��8(5��L>��r�w�-e�
�]�s�/��s��Ȥ��{SAci6H>�C�}��j��/�6�-��Н\�vF�ʗպҪ2���2��Ҷ�XsO)M �����NS6xS��q�A�a�m�ь潰%\eNruP镗��|�����МǸ���t��\[J�'����m��1�LYط��-�;����Q����^
a�]Aਫ਼Q�.��Vmgd�a[�KN���Of���ޞ�M���X�J��|C��� ��y�9�d�� m����=KSܫE���l]2�[��z�K�Y��yr�맍�e7��'p�5J+�F� "���՗�HA�fpifi�W};T�7SIy%���UW��'�'������I�E��OXsggjP}�`�BF��*8�l�����7�q�,տ{о� �q��;���I}^�;��-�����fvڞ\t�;����w�*ݣ��oK�n s�oS[�{ý�-���;�z�AiU�	́�)M&���bۈ|��Q��ow|}k�}2�;u`ov��It�Ɛ��+��{���)]�:������rG�m����Z��.�t}os����O��9�s�OK���^󥷫�#��.�}��	������U�^�#�=~��@0��"*y~$��gO�+k��B��C~���-{�A��B� �Y�g�̊s���j��s�'&�6Ѕa���D�Zd��Mӽs8�i�[���ݮb��ѭ���Zi�঱��=0��N���J3h{;E_QΦq��)�52wyE�L^r[X�T[�_l���P]�#V���t�.rnɶ:����ڤu�g�q.�S��$y�������Wu��j�Wl(櫾X��p47#��v_&��Rr��bbM�V��&�I�����4��ֵ���ה2�(b���;؃��lKHľӂ�XL�^��5Ư������Ev�V�,��.�ߵfW��lv���КμW4z aP�uu�>��_�0��l�̐]��*�3��'Uw�����O���t���5�V`�y"M_绘��K0�N,��f*s��Bޭ��n�y��{ˋ����9�CS�����Ö�����nv���n�3:�`�P�.m.�/Aއ�+]��Rx���[�É^B�
�ꊒ-��i�vz�2��_e��m�Փ��e��l*m���=�a��o��@���Y��s���7,:�N�(%^����U|��1�-��7��)z��|��K:�߭�ʾspI���uhy���Iu9��#����t������9���c����%G�}!�^��ت�+��@絥SM$V1��{�,a`�E�v
����(D6UZK�\Iܫ��T�ܑ�
��\��9QM�Xz��y��n��$�����plR��K�� |�j��d_u276�ei��9C��o��h�F {�|��Q�lS��xvH�B��F#߇��Ļbr��n2z�~xd��h��ظ|-�* �0�Lo1N.��1���Z��ay�a�~mVi�{��'�V�/i؅b��@�p���T�*0u~�vny��J��쥵q�>��'����PN�Ysl*�S	:�y�w�������5��j����;�^v�f��׹>�p�k�cs�+u�����j��2�kV�,�}q:��Z��<T;���������(�O����F��7ڻp��࡫�P�l�/s
�t���j��AoR��Lͬs{g^�2ld���B_q�O��[A%T<��gh�n�7�!v�����#��s��B���c[¥��>mf}r�����Y�8�.wim6��Q��m뮙y{����j���y�n̷�����/K���C�xf���x��<;Xݺ���;/U�t�׉�W��rޭ;�޽'���,�=�u�рw�P�nCIpv��yE�f�/��v{ED5��z��Um,s�	�����5�^W�s�{��[���T�	�^)�)����O�g5�����S̫��'��s��S���2�gc�`cdv�6ay�U�� ��7Ui]�_x{�͵�Ě������vz�(>�b�	�\ͪmߜ�R�[�Q5`@���;5��Ԟ�Ӷ��u:�>�A,���	��T*e?/d^1�\���ɽ�j�{%�e��D'��j�?�Á�="��g��o	ʹ�IS��{�ܓ����cri;G�߱���� x���[�|�x�iI�9ς��i�/�n�	�����R�}�[�w�d:��Ǆ�a�F�
���My��tY�v��M�m�������@��݈mkڎ�����9.�sV�ܘ����c^Ԏʸ�\��B�l;�	����uf�6so[����P��0��,/ǖ���S��y>�6{h��򳆖k�&3��Z;~s�������v}\З�^�Y���j��N�\5�foW.��F�(��F�����31�A|�'��x��#۪�ò�#g�7�9��(S�4k����#^sw9��w��i�ݜ��ۇ�� 2�`5ڈ�����U��ڼ�8SVkg$�d;��
��	,�u��H��s��xd��N
J�rG�m�7B�g�QJ�KA���I.{���E\E���8����������ܶ��u_yꩯv0�6��%�a2վ�ݗѓ�Q�t��jkֱ;{�5d�ҭ�{}�9����C��/��
W���d�h��$5�u�����t���z�}.i��X$��5�[�k����IZ��f�v �mC���Q<ȼ���@_"��0��،��o�ICgֻ���3(�9��4��m'� 墮��|�Ҭ�s�3���qB޷*�v�S~��Y)��2��	��q1�l���&��h����v�[�{:�oK�n"aWTF3T�C�u[�����w��w�&[ۣ�|��|�9��)�i;G�������	�.�Jf�t\����zf�����:�^�K�OVpT������dԎ�1��"��޷�������ᬫ��U��պ-�z�8�b���StQ*	T���l+b.f���
���.�ǣ�8�<g؋Ii)S�5��|3A�r̤H� �Jd�Ua�AI�����6�k55;�ى�5�U�Bm�Q��Wg2�},	A�X��\���U��_,�ջ2S3Q뮮=*�#&Tځ��B�=��ڹ����s[Y'�o�X	��@[�TG���@���C�ɫ7p>��J �e�d>|����%�
�*�u؁������/�N�����Ab�K9�����ؕ�&�f_P)]	K�EKY�_��=섚��2�泸{d��qM�|U���R�oC, bv���BvE@-fm�U
1�BlK�k�y=s�@�_�nP�yX�׻���؃�M���}�5G���)l�[�<����n/Zܠ�"o���$dүo:��a�<�:�5�N���o�E>�g��<���NP���.2�s��Uߧ�߾�4`+���ޅ=�*�jWj�u8?f˚Y�M��a���p�&o՝�q�ɔ��ש��^9��v�E���Q=�L�y�姮��a�ockȱ�e��;�w/�T��J��QA��<���̅�a��bF��`t�O<�Zoq� ���M������f�c76�����;���R�)SFd���,�R[���5ދ�U���5�u�,���i}n�������d�&��6�Hi����0��w�ֳM�F�����)u�ĺ�O)�W�	ro��M��\�D0��B�] �>��u��s)��|�z��
˨�RZ��R�e	�`ϛ�&g��a�n�	J$;��{��.��3��CE�'>�ER��������C����`ZMM�tu�C��5Fo^��5vOJ�#;J
o��NT�(�ɍ�<i��ޗ��V��)��G��iW���C;��ͷ�:��W����7O`՜n�.G��љ��L�bf[�	�qwa���@����8m�T���]�uYK����A��&��D̙�T��Ҋ&�<CkF�5_6+Z$Ԅ�ɹ��i�K�,�����2kb[�t���vt�;_6����V\�Zz��5��,mv�������u����G�j=�Ӽ�M,��z�:*��2�&��}@mD)S�j�L��X<Q�I�HhF���X�-vP�����C��|*�kn۩H�D��>夜T�Qܷ5�pR#�i���bE��e%�� $3]5uą��}ñ�/�U`t�M=��.{���T�@��Z[���*�U<�X���h����w�ev3"92:y��˰��PҬڹ�x+�����qإ^he�1h��dS����>0�.�7ZHVkC�'77�Ds*��Ę���#/V�7b����7tI$�F��3(�.�n,`�3rf�6 ��R�A�ŉ�bج�ϲ�9�luҝD������sz��m���WUw�M��+�L;w2�d��5^3o����a���[�Cui��P������X��9�����M���@��ob��<�唹�Z�+�0EԈ��Ӥ�[Sv�V���C����5XyrR�-�NX����M�c�\�͹��ċu�zF��rO�E֓Xu������;F,f&�g\|F\��b�Kn�Nv	{�]ջU�_9 #2Һ�f8Ru�;���u�Z��.�v��&{[/Pl��!��t|�CYo!�ZL�d+FnG��u��\�z�s|�9k�uVn�D��Hu��]+���p�p�$�5��Ne���F��9�6��,���s�x�BwP�[$�6���*7�Ca�v0�Js����ں�`n��n�Ya�\�<�V��f�J��a߹��&573��6��Cq�2*;b⾝�
{��|�[0�4U�\u���|�lAV�v����WS��<*eBo�9(�&�\�90�#+eQf�i��η��f���;WW9%:
����-��bC��=���\��93
��"�����'l��>f��V��f�g�5-]�G9�|�:z;ڸjS=c��t�Ʋj-��9����}��\��V���1=NΖ�*�'�D+nryԷ-Q�E
s�s���ۜ%����N�*��y.�A>����ct�Cv�4�j��p�Y�������%=��QU��X"��Pek6�,EU����T��������b�5�-eER��
(�X����bƍ��DX�V�����+b�֥KlUUEXѱ��Q�����PTQF1@VV�b��b��DF**��eV"#[DR-�ڌQ@Kj���(��,T��[TEQTVV��64eJ��Z�("6�e�TDEjQ��[PEjb�!mAAR�hU#���"�B�ʕ��Q* ���
#dD+jZR�Ue)m������(�Ue�j�"���e�E(��e5
�����Q[J)ib����h�+V*�ւŋ��J��*aX�х�*"(�+(�AX��Dm�TKk-�F�-��*
J�"�aP� �U��DQH�JȊ�kmTX�����*U��c ƵZ�"�[H*1��T��`,U���PTU��QQ-��U)Im*(���DE��������V��u��$���_g\+��%;�t�r�Yˇ>�>�
e��S�!���Z�M�ؾ��)ђcX�����K�����Ew��t'B��K�C��mSn��9nl�8OLyl캞����~����8#��Ri9�v�˃zI����{�9������rR�/F��{�!�J��h�4}��;\��0�ob�<�k�����fX�+Sj:�cV��޾��4�O'u\3���S�b��Ml�*Lco�5��z�3@��m��V���꫆����iu����5��j�JN�����y�Ov��0�^�V!W��~��&75��غk�k����=�UÐ��_�	�0�hN�Ysn�Xg8�<�<@�t�,N�mG& 3�U�N��
}���}lHk��{n[;3��姥��K�u�;|k��%q;>��5+�OC��m6�6���n�گ�Ü����{����1X��Ӂ�f:a�� �þ�Uλ/��^ތ?Zl,�]�b���{䮥�4�U���^�����^���
��ee�+h	�N&�tM��&nݗ�
>󬆁�u�k����Z��m��B�0Ԕ��A1� W'Lų(��T�>3��u�<Vo1�m�M��ER��|i�i��s�p�]:~��,-ZeV�}����)���A�}d�V��vA}�sOH(%B"s3;&-q\��I��+�a�y*Sᡵ�o�^#U	8p��O�ty���d��k�4�����ֵW�ee��|���W��ٛ��TG���Ro:RK1�jr�\m{8[�����X�;j�=̦"��A|hL�u.��W���Q��#h=�#��ل篁��	ϝ�m��YΌ҆w/�v�"|���~��<�9��
z��0�=(uÝ�8��VJp��ӝ�/��p'�\���N�z�*��"�W���ZG�êX��#��J����&����)��#�Bи�(�@�<|���7�V�Xuq�g��^���;�H+�ޥ�ct��{-�c"E/w=���p�[�N�k�n�J��=-��ݺ:�cv��5����X*�;-�;��z�4����^|�/�WFK�D���9���C�%�-}�!���M4����v(��y�6�)�<I8f^��8q��'ۻ�U�ޔ��;H��s�q wa?�y���v�����|����bs�]oe�1'��>}	�Z|�j���H�&3�zGcz���=~�%���M��<�ݬ������o%�ν��*n������~����S��g-TA���+r��j(�E?FZ�����
٣�	�!k��]�v�;��g���G-�1�6��[�_4�bC\n�ܜ�h�|���P���N�ڑ�o����I��3�W�ckɱ!�i��k	�5o�,+Ι����bw��{��8�wr�����Mf���ÚyJkɡ<��\;1�uö���{ϖ"yٳ�#26��.�|�'^��<y??yc�DU��Lj^7|�N���^K3���=�&�?^WJ�5f&����m{�W�v'��(��T��<�9a����]�T'ghJ���hK�b��78��-1��ƦZy�f����Y�t�z�,�<��t�U��1V/1����f*���Uث4�/��
l֩:u�7{��-�[�m&�N�ܝ�&�`aq�Dn��wy��k����9���`\L��t�WuF�5ˤ�f���	�h�[��M`��o��|�)�pb��΢:a<��P�����=����u��
�����qC�m�O�=��§�uh�Ҷ:�9Lӷڹ��~��	�u�=7Ψs�=�G�>���P2��6��жr/H�7���n!��DWe	-P���`��X��S66BɆ��<���{#����U�~J;�,C�;�ꈎܡ��u:�=�9K#3�Cv�kܱoիMx��a��Bߒ��!`�� ��v��(��q����h�ko����#�;o19fKB96� pXh��[Υ�T��đМ�t�O�B}��'WA��a\1KNnZ��qb���։,w��s`��f���b����ճJ�.�Ch��X�K>3�!��C�?~m_�V��}�����g�Sc|�1wWi[����y��E/r'�B덨{���n���ٴW�5+ٞ'!*��ս�_t״������l�b7�mp�_,�KOren�z�	Щ�U;r��6���m�Mս�G2�\�1B�u�@�8ηFĜ�ӇzN�q��mdy�w2��寑�mnA�1	��g��ٽs�(��ٮ�Z�z{\����]7I2>�3� Ƽ��>9�hh��_�9�7���Y�rRN�O��v.��Ҧ�oS���w��~�y���a��!�<30����.�L��@�op����V]הˡ�+^ ��a뷝�:��PgM�f�H`�,KGԽL����+g�d�Э�N��c�S��.�&�-�ӷ�y�m�7�f�g<�V�ý�z�;Y�{R���E�7�3j�l��}��[*\˚�-d�Wyo]_�-�M����r�NI�x�YQ��<�����gx��b���;�BGoս�ִ��>�{+]�1i!���>�������||UL������2:���]!�^��7/��*{��m6��P1L��޴��k4�$��b���%@N�D'���^f�Iի��27��ҡj��ݻq���{�n����X�@7�߆B�2:7#.��}»���٥D�Q�I 7[��	
%�Ne�$�*ݓ�zq݊ls��x@���/��O02^���o����)��nM����P�ѡ�n���M��9�^���e��L��̔1UϊU֔ޠ�H�.��
�U���зjGd����u��å�N�C4��2g� ��U�w�����>�3�~��Zd�,Rsy
}ݬ��C���=g�ʹ��Y�x�s�l�ŀU�Ak:X;����}�N�y��w��v'�k�sV��ѓ��x�H��c��% ���>����+/������S{&�l��v=]�R�v��cS@�h>��2zw�U�~g��=g�j�}����{���sXsf���eHC�N:ʏ�>�&��E��ر��+�_ ���H[�٩tk9�oҮ2����]2�����>�OR}�2�sa��bn�%�Z���S�S�%(��[݇��X�v���]����u�f��{�/$l�8nz�q���˕宕ru�������yܷz��7X�k({_gXz���XAO_�Fd��9[܌I���8'kAOFv9���O��YʞXWo��f������tG��]rOiݨ/
;�p�IR�{@�έݫ&\cil�����Ei�PGf<̽���)�'p�o��U����,Ҭ��E�������4U�݃:Q�8��T��	X����nܧA��ZU�;q�\/�I�ÉR��} ;���y}Ʌ7�⩩=q�lb4�{-
�֔B�V]H��~�Ƚ5U�WjQ��3�j�J�w�{��9�)�}A�NG��.��cw�ar9��PC�~X���M�m�����S�n!���VNwd���KoV?�����~�x$5����kJ;̙�q���mM\�=��3:��uB�w�V!8̟xY���t:;�Ŧ��X>�4N��V9�WZ�pU�'F��cЭ��	+ŗ�qr�e�]�|3W����s�h׷���kM ܜ�3^��|fiI�]�8���-iA��O�fU]���]M{�4lKHK�6�yN�;��uY�����e-��b��Y�VHɬ���res�����Ks͚��~��7��{��Pkd�Yޡud����Q����Qd,ĚǱ�V�-�6cxV�K��
��]oG�޽�]Σ��o�Y�����qǔz,9։���sP���Z��V����},<�&w	�ot����[n��̄#;��r�H���NP�{hM���Gי�ԟ���x��Ծykb@s��m��*f���[�-q�E�Ss�<�E�Ex�O+����/��2_���G1%��A�3[[A���g*vv���Iq����רN�'�Ե�L�ٕ����Ň\pꮃ�q@�B���j���lKՓ�|��'�M�U4}~�$�����ݕvA:���ʍ����=�K�f7�RU�������5!4��{:yM�L��	�b�\�ԱpV}���Z�z����y�����K�OR�U��RiW�����q�'�Y�|}YV�����D>�w�����Z�����)�V�kQ�׺��ɥ��/iXo!׭�*#��B5���m�;��.��w�:��+�]��A:f�{N�X�A��@�v�u�iE��aZ��8o����]/\jgÌ�ઝ��^�b0��ə�(P�0= _v�ʵ�<�N��ր-��ʘ�㚰�W#�$���JY�vB:�2�ew��i�!:�n��E[f��0�v	�[כ���Q���v.!��;'�B�uH�W
}����j���76�h0��u�W��ifv%p��ۧi�̓{���p��ؖ�� �����ωit[���'��QL�,�>��e� �t.�V<U���ny62�$��:\� ����w8��D_��5��M�>��<�}�td�{Vo:+L�|��q����������MĶ�����zb�|K���V{�3[�1�����3�=�&9ߞ��^:Ck0�}r��#2M=<��MVt�XA���5<��Ҫ�޼2�����W����6��PgM�5l�2�a�F�����sӔ'{�c�Ɨ��M�:]a7�a�Ӵ1Ҧ^�E�,�Y�9[j�=�X��ň:�_�$o.f�6�ʺ�3O`������Y�5S�Ԟ�Ӷ�DL*ꂤ���uas|��B1�J���Q���7L�_(�=�DX�!�2�
X�2��������9�3Ϋbs]A���^����&6	[b�����Vjd�������1� �aD���Dd{8�ŷ�|Q}�P�t��#��2�=}�������̖�<���-ysuQ�'1vL����W���nnu��!#�Y��v����Y�J{\���Y�tN#����+�cs������c��A.<_@i��ID,4i߭m���� ߎzV{c��.^�oiX��V��x��T���.kv�^=�D+�l�r�[��m%o��Ov�n��^�x5b��#=�]�l�JS��+Y�L@�'ѯjGd���\���Їi9wf{��*��5��u^򥷪ߣlD�s\0��krS�����r}i��V�1Y�N��qP�Ng1��s��U�^�:��Gc���)^{K{,��d#����o.��R�i���֑��p5l���g]Оoi�î�0yl�l�N9M��sn��]�9O�a4$>�o��[��}uiy�T�Um�7��Z�5�X�FM*ޗ�;XtJ�	�;1X��c���x�<q��e۵[:�e�j�#��h�]Ԭ��m����݇\�{�<f�QA��ĩ�N�9����j�����Wq.w��v�G�EMfh�4SX�vg.���7�ԁ�6�&��J8�&�a�s7���y�zv,9�5�ʞ_T�;%ҡ����M�ע<�6�^P�&a�c���]:��3I<�A�+9vHÖ򾽌F`�(�uf��-�vb\�]e�hU��^�\��l����חc^F�6^!V�
��������A�+Ix[B1#�W;ޭ^f�v0�t�;��\cxuL�
�Y��z�M�VU���{��_=Z�m;6�\\�W3�0�}�
�e*�p t2���e�Y�X������Bs0Y]��/{��Y
2S|��W�1��J���n��J��F����{�	97D�������,ؖ��Y�g	�Ue���26�ަeu�R���f\��]���f���̥NoY�R˛�w#U�KN-9���oS�)JeN%=����y�;�^�\���z�Ҝ��q;�]κ��Q�e�sZ��[Љ��a��Fs���h��`�u��
�T!���Kyu��;M	3pYu���<�-�$�s��"kj�oB��c	����Z�}.l�ֹ�5}f^e`��f*B�G����n�sz�51[����)\B6�[�8�����WMU��k��V�v&�ĩE=�>W�8��峪���rv1ӹ��U�w��#����&mt���Z�[���	����t��E>YE%�U�uو�t��TƝ�V'�򣌎�a��S��wj��ێM��i'��+��KXZ;��8b����6Qb�ءxx=ԩ����n14�e���	:r�xJ�3�MN�����1������]e�[ ������SWU��a�꘶�c��ܵ$��$z@WoJu���N�����DR]����TCp�d�V���|����.���Ǜw֝r��$���X�+#1`��;�f;,��6�+|ݬ��gf�}nܚ��P*�������W��S6�Ԟ);��	�2��>�ިn��&^�����9N�Q�ʍ�z+�4+D�����7Rkj<��e�jC�0�kz�Spa�Y���V�ޠ��dL `W4�R�v��B�f�tR��`��Q��2�gIE�3shoǾI�Z��*�J&��r�n�$z�[���R���ff;M�R���,PhANk}�:���y�(KW����p�7�k6��1�A�t⭑o*�:�8G�7�5�:����B��]MRd����u�V)�۽j��X7EIF�ӥ��frGs�a�\v�&����`��6*��q���^�6j�^|�5�����|H��<�[�c��l�����'�ugf��5�3�1���X�W/���H)�i�sxu�U�ں��egt���XM�?GP P�*"TU�T����D�Q��m���)ib$F����m!Zŕ
�U��6µ��U"ʔb�XT�F�Ȩ�e��TQ��K)-���(�,X�ȫP��ւ��
�Q���b�mcTR�������b�ШVJ�,���c1#J�*��#"�`��R,QT��X*���D�DV��RF"�E���k�-�j[Q�X���d(Ȫ%B�(
*��E ��A(E�H�R,�T+@��,R�eAH�(�
)QR,
H��E�����*E�
�����ګV�`�j�PX֊J��¡T`��X%mJ�DP��YY[h
(�TAdmPQUb�UFVJ���xG�mn��'�\�Ժ#�iu��������=���Иpf�%�5;�iۗfKm+��L�YM�38Z:��[���L�m2G}�[ ��=Qv��]2���O���x���RBG&��_=�޾K�f`���1�/�59By�׆p��{�V����NZ��c��*.��~3�����ṵ���r�;3�ھ^�0��S��V�/�vƬ���7���ӯ̸��N�SXSk����%^��[�����V��:��3��m����֕n�D���Ȼ�n7]�I��_����z�C�s"������MG^�҈P���2@�O<��]��u���/�Mן�שn� �q��wKMb��VG ���dߗ��GR���-W}l���-��T�=����k�}3�mȴ��糧�2�Ϲ�G�;a��@1;�/9��7l��͙�!}�@�N�@C/�h��}��޳�P�������<6�jDf�:���Nz�m��j��Y�g2�
r�)�4�m7�Eة��}�.,�
���78_3�(VoV	;��7���H5]��Yk��Se��Lm�f����r��7�YNpwQڳk\�S)�+3h$ε��6`�ۗ��x�ַ��N�6����;�{_���y��3����\�oR�`ŉ�mu���\�g&*�Vt9��5��6Ƶ��8)�f8>J�#�ۛ�=1W4]v-���z��]ȵj���A�ؖ���M���Q����rը�]p��H�ۻ�ou]������+�)JP�Ϝ�qF�.��{��3��]�������T����|��;�L�+k"�s�Ș&/%�3S����b�¥��t�ݙ��������<��7�[��-���-*w2�񦹇���a�kcj6��s��Nʦ�um$�ɐ��x/�{5j�t�M�[�M� �a�
�:�����S@��M�˻O{��gS:o�\�! _'96��U�G��ͽ2��ᬾ/]�먪�O����W[�I]R��="�U^���v������%��oc�ɪ��zw�8�\���@�n�n��N�s�9�YG�N^,�um8b���t�%h����]��}�v�d��WJt�X5�<$s��L���c��]Gg����m��S��=����f��B��3�R���e�	N*N|��]�޻Uk�O�{�?v��N�����t�5Ru.l�bկrűZ�s�x��u�%@/Ϻĝ�uN��DG
��qRx��]wvbB�j,����V���B�1�2d"N�	5�r���S�R����GV&̯'L�/i؅ba�z���wV�t]c���q/�9���W5>�	�;�;T���ݣaε|A�x�m
��>Ԣ2lgm�_�ZC*�˥i���f��p�CbC\n(qԨ= ��QK�yR�\/+K�%~�з/�ޑ������m���ܹ">��Q�O{]m�b���N
�Y�X��/s,J�Cȹ��^X����{�v���ګ�$�GBh>�G }��3}Q�%k�K���<��6,���L߱��f�T��������a��4t��a}Z����s�ړ̽�]k�|O1�ܬ�2��7������V�?m�������(�� ��/��[\�2[8�LNc�<yݝ|�Et�2�=Ʌw(�gc�U�Ѱm��G�2�(Sꋝ
yXz��ݘ��;�]9���֕�ܩ"Р��]	#�oN♆��o4�U�*��/^y9j�z�v��o`���z�����pzD}�HA�߾�Ź�̣]�,��'��'=�^e�P"I�����c染;�Ǎ���Ϭ�>~��md��c����$hk/G�תgjs���r�U�	�:�Dl*��$�Pz7kw���v�8�^N�~�7�.�E�x�=����ő�qp��T$<����ޫ�]�6�zsjP���ƭ�yh6�s�3������OR��� �=ۯ�˔�`��ǁ�ܜ���O��K{J�c!з�m\Y{��8ͭ��bǚ��#k�i�w1ݺ:��Ov��0�t�<Ҭ&\T�ŗ���Bg���Lj�;*�Ϻ�-n��k�{nq�Y}��m��f��;ф�D-2[�)9��>���vm��![��b��������e��K�I���[9&A�tͬ�vM��-�J���vb�:��@���L����f�u�,9�R�Z�#�e�|��y4�ά���f"���WTSf;e������ ��,�##�aF����%M�n[d��3{�;a�_/����+����:���;��镗��*��=�B�o��J���k���+����I�-#!���h�f��0��"&W��{#���M�Tu;��ɵCu�xv0�@���4��S�j���� 0�f,��ޝ�g\�P��d��/4v��<�5��Hmft����5����^N8`�,��`]�&�g�3�z��Y{���.f��\�k��cu�Ґ�G�|�c�ʯ;j���w�n6��-�/V��;��!5׷O��{I�?�^����Ӿ���y:Ṿ���ِP{W�3�+oh��ڲ���KWX
[v沇>�Z���u:�I}�n�y�ڔ�7S���-�HM�hrm۔������0�:xff��"��["� �����N߱� �4��{*и�HI��N5�H������Xl%fL����{��C6x�� ��v�6	�ٌ9t0�$�+u>� <Oa�%v�g!�n��]�b�ܫ����<�/�q�9��9�����19ك�쥱�R�w.�Ӏf��(��rx�'��u�*�e慳���a��SFKѧ�)�9�����{k�L�F;��t���RݼA�>�~���Ln�:�%+�V=�>��@�\�\[�I��[1*������'�yl
զ�[J����O�i:��s�!�����rhN���
�nbھsڲ��.p�('N����B�	������'{�sp�h��gf]3z���lt���	�;�Rtm�l*�za+'t'8��y�ۭ�j�gu�p-yo��s9�>��5���؆Ć�����2�܅�h�)�<jRڊ��给~��)^{:�S؃�M�#���SQf�o2d���r g�u�K�Ȟ�'yu(p�-�9���*^���I��h�b��]u2���Q�>�z�6z������:_��k���}�M�Ӿ��Fk�ѩ��4󭵙3���q��ј����p|` ������L��K
p��P��	^vF�9%%�jo��.���mM���nnAƟ�U�V4���联FM-��	Ա|Q��v6T��GO��sD�ϢNY��=_Iy���` v�{��������e��=��wբr֓r�&�Y;�K�l�̌L�n<*zzsjQt\N'�Z�'-[�o.��{Q��Fr�݌Pvz����g_<'��1�p6�'�/U��I�9ϭ��i��	�GI>Telt�߻6j�
����S �BE��l*m�U�G���6U�n{"�MU��kV�)����GWTt$��(%��s��9s�}�a��b�[ɷ�=�np��$%�����5�MN륷����g��-uU�Vf��;b�/���V�c�ai*�2|�#�I��k��#b��w�QT6Z{���s��Ʈ�_Q��IM�#c�n!�K�2������rP�0r�Z���g�%�Ԁ	)`c��E*�0��xx';��۱7/�Ȱz�+�H2͎���}i��^O{�D@bQJӬ�W6L.N�%��!�w��K�=��YNn�v��4v��i��帐�0���cx������Y�G��Dπޕ�L1��{Y�ջ9 �S�+��X�@F��)��@��0��'i,��&�R�hM�Z�u���qL�V��1I���ywm^>}�1�Bj�>�G����R>r@�G�*V#|1��9����:�)��U���C��z���խg_�E��59U�a����D�.�I�����d�S���(�{�;왠T��Ћk/pO�:�����m�h����!�X�2v,�b�E���7@�y���S��Zl�k�1X��L��IB;f�@���[�R�5�{w�zQ2�P�J�d�AR5�OavgA㽬��k�n�O3����rV�tTv����?i�;g�Ň�_E_��A����M����6�.�A���*���K���zK�'7d-�}SKH�Q�Y5�B���0��A�j�v�7D��ks�Z��O
�9q;Й��7NY;~|K�<C���s�Wl~3�<o�j�o:�g,�K�uGCӰt�# 'T1T�N�~lS\��ʷ�*��@�#�9��;��u2��yަ��]�ck�#���vXz��9\����Wv��E�WK��e���o/�3�M<�I�bn��h�&Ԑ=�[���;7 H���]©	����L�V��Y�D�"�yY(�B�������3Ɣ�����wX���4d
������>����ʎ�$�ϳ[��L�&��"rs`q*éBwU'P�q�Q6-���|a��m�ιC���C���O?k�I��{=�1�9	�Pe����2�K�FFQ�,mNr��[�g�}��{��*Wd�*$��ĺ��e���sAjÑ���۝´W���O�o���]��3ewV}����bM���>H��3���KS��b�n�6�X1L�{��_lT~�^������ě�tc�.�A����sI,�׭R��ZC墏,�� $�~+�Kψ��V~ٮyx����wS�z��o�3fv^5�ޟ�s���r��R/%�z��]�u��B��b˟�3;��כƈ�^ʅp���#����J���)����VK]���Z"�j�c_k#'�om���ؐ���Ѹ�M#BG	5��U��eb3�������8�����mH��Z�������׫g����7������؇@�'uSv�#F0���ίT�Y�[�|�Kn�����Ñ���=�Fw��W��="��b�{6�CDFЩ��A��,}{o�%����\�f[H��t�h�υE�r�:��p�۬7�bl|nC��D�/s[��˳U/:��ٍ�>�:��A�*��:q�1��!��!��D)�fƅ�F�D}�L�Ȩ�\�;Q�iֻ@�:�$1Y�Z4 {�;���J�-�z-�w�H��r��pAQD)O��nH
�KC��D���Uy@�n��t6sP��N�t3'��4��5���T��(�XFR�Sy��G���j��%�J�ڪ���ϊ�緰�v�7�Q��y��hbt�!�9ܜ�+���"�癹�J���� *��6U8q�s5ls[�Z�$�,����9e�#�sz�����ɕ��)j 9ʾ�Z�f�@c�!T�C"�)��-�ՂG53b[�yg2/�(Χw/{w�&�%��HV��wr�(�S}*K�EK�����Ұ����5��Kz9�k{\N������,s���H�3�s>�*9��PU��5T3}1W��T���8�@��m�tٺ��^׮��R�g2u����C	&.�Szx��ςm�Ë:��K�7����1ڽ=�O���ek�}#��_\d�	����m�z�[���>�d��F��:���_r�j���t�lۛw	4I#��q"u��Uۉ��^�_�J��̯n�z�_Kd���5Z�5(#�A�����"��Dƭ�~����NλW�M��O�v|B8�:��{����0$gm�)��x�b)�he��j�5_saVN�<gS�r��h%�fj�<����7�$l�f�䜔ݾ|���ᗂL�#}V�N���j��2.}G8ڛ|��E���̶lC���H���!w�ڝ��ܭ�pS��h���h�m٩Z�����S�C���A*�C�κ��9�!��m�ZsQ����t��&�m:E��f��]G���B�;(FS:>���I2��~:�P�wm���BÕ'��U��ep؍��kT��ߨz�.���]�ۢ�Gp%���ov��	f�5ި��x��Ju.��O7��2�4pÈt�n�u�w{��}˶:��-� �1���Pl���pܵ��d(���y�����wb��R��Ej��w�4C���L)9�Z<1���v6�7i׻n�ň�m�p�v&�TnJ�&����lM�N�E�"L��c�x���~}}�����w5�wS�Z�+F��WP�v�66�_�^:�>��:I��p�
���:��N�̱B���4]��	����3+mM�J;)P���y>�a����I!��/� W[J�,�4�(�ᦸ��5<�יݒZ��w���)�]�F`�ؘ��wr�
z�|��4bi��f�c�z�ǅu�T�.^�X�d�
;�X�y���͕gw%D.�5�D,aEn�]��gI�T��S�u�0���T��&9L+�|n�wr�h�C��u�mXU��2��s16��%gQ��K%fY���Y��=i���
sw�F%����SMΝB�M���ֳt1�Tc7ݠ�L̛8�f���[kf}��D��*@8�};{[�jݓV�<Gq5��2���=a�<5��fKкLym�����Ŵ��f�	�Ӭ��KZ���܎ЉU��o�}�m|�iq�Y��oF�L���y�c��g��Pcs��u�(�"aa@�+�Y�N�y�X�F�Z	xZ*�jʂ=�$Zlv�gl@V#��N�(Į�z!�}
Zԭϒ�/�CGTKB_c8����u��ib.������z�v�=�\2M]�$J�u��[W�4�J�͖�8��˜^��s~��R��w\��uyE-���>��V�%|�^#�ZkHl������l0ǧU�J̣a)��{�e�q�:l��g�EZ$⋨�]<�C3},�����wtJ��vu��k���8L���7P������V�vͳ7��>3���}L*��Vq��D�V�7�|�t�γ��aR���9�;�U3�x1�T�Dŏl�V��8����V���`����8�Q�w0�z�`)j��׼�%��J�ߣ�1�Jէ+���X�t`,��[}\Өn��<�>�ܔZ���iه��R&P�����6�ɠ��E�\��7�&oV�՛�qx��q�ɠ�l&�rW���T�෰��.�*:�k[-W5��/V_,添�۷�=�m?|j��"���Qd���EEdU�$Z��R��
� RE�`�`��`"��F�d�����U�`)�Kd��KJ�V
(UP����k��B�E�YR�V, ��AJ�k
YP�`Q� V)XVQR��[B�T)l�T����+e���Q`�lQF2��(%)X�b��
Ȩ�6�T(V"��TY%B�AAUTPZѨV	��Q�eh�-1*H�U+-�U[k2�q�����LfZbbJ�V��⸂�"�*�3)J���� �&2��eLjeːX)�+��`�kT\-(�£\őLc���0�Xc�B������
��FB��+���5{��5��׺�p�L�k�Mu�����Ҕww��1K�B�(%�S�նl.�xƉ�;׽�qVf�hof)#2�'��VҊ��0��L/r}~���Q�����Y����&�� ����jjvN�wv�Ļp�/5��
�1�����*��veS=g�	��<'پ�Cf��%=a{	��6�gOlm�[�\���8�s�;$������#����9�����%���N��n�I
����`ru��Lz]�y6���5$�pv'�;;��l$`��#湺[�i%���E���h8�35��Ug����s#�^\��nQ̞�轌I�U�����u=GlT��k>��N��D8��B��݌���ZgH����%\�c�֚ս��..�eX����d��G{���0����t� ]_d������Q��{���,��EėC�M����7O��� Y�}^�QI���W�V���r�of3V����˫Ǐ��4�$�!��^��R��v廣��%��'��Ԥf7�����0-�,�x�!��У��ی�'IX|�� �P!����Fy��Q*�^*�v�OVl����4��8nnZ��~o<_�/[��F3O	6�D��`��s���;�W���*�^�!����W�-��rE&Z�x6c��r�`<�]%2��_jX[�7q�fά�{sU��Ox�
[�E�㺏�M�{�v�;��%&/r.����2��^�(�ȷ|6X>TΠ��\���R��D�:�r����TH�w7��kю��Xk�բ�ǝGӐ(�]�=� =8���n�ߥ�����@�kD[ͺ�D��,����Hk��q1 ��$��9`�5�&�څ�Ƒ	��{���C44�Û��]~��/��5�ȉ#;�O���!F庈q��yi�L�ޕ�I�a�3׃��7O%y��F��)�dV\j�:Hu�ύ�z�(�W��졕�V7�D1T!�39��_j�����Bju~s|���:���ʜ�>k��ʦxW�����+b���w/b�>.Д�]����\%$�Ӭ��k
Щ�{�9jצbJ��/��r*zM��{���z��*ó�]���~ã�~_��}~s�>mV@6��75�7\�mmȭ��+;q)K��)�,�=¥F����W�4���u9�p�L�]\��1U[���Χ�y��^�Ɛ�f,'4j�2��\L���v,�xr��,�)��2/cW�@H����wF*'��k�Y;���6�Wq�#WQ��hM�Z� HX�F�k:�Sm�ʻ��D�����YS���,󞞉f��V��M����ğ���j�x;�+*�juͼzJ��Ӏ�']���h��u����ciM��ɀ��s�:�d�1ӊk�7/9����ڰ3�X�cI*�Xkc�b���[�����|�Y�k`�ٷ��K��QղW^3�==6���	"�W�v��Q���E���XU4�Ovm�̬]j�\����C\ړ�>�_Lg����/5�&T)Q|@`ޡ�l�w�<<�N��nok�:f%��fQ�aqQWʊ"of��VUl�19�><R\�j]�}xY��\��osD��B���P��x-Y�}�`�BՃ\�
}�%��f��*���%֭�{ۧ�"}|;,'�����+튁�yz��E�Z�N3���ȧI:N���v��˹�ٺ񐣽��:`j.��"N��v"h��W�!�N����SV�
�B�eqz�����Q����޿�(�!.�K���)3�����E����um
�����Z��	�I����So,�6xx���*g�V(��*� �~K�r�%�c��1�Ӟ���}Njʻuut�$p����8����wF�q葑BO�r�6"eb3��x-��[֔�����S�ЧN8v�[y8#l�@bu:m��f��������wb�u{�R�d�I��nȸ��2̷�x�
>V�$�/@Kh��Ons��ʊ��ל q�T��痽�l�-�%�	��ӌ�����9󢲜#��h�t�\y�k\n;��Z��Xg%�O�x��0�;>���+�>R�g�۽�{�]���.^ſe�F8�b�ճ���ַ��<d;0�2�Z�UW��!�;X�F��m:"�EG]�e���xD:�c Ł�*d���z�ٿ��>)r�ܫ|<���sn�Pwi�b��=���Dn��n�P�C.l���{�U{���] �Uٮ8ޛ�̘�*"�K_L�U���x��������W��	ߚ6=��۵1��Ή�l%�u���{~B^Q;컬yJ��ܲzD,~�#!DE��\�yUS��j�Y~媶N�+`�`����˝�̲����F\$&}�j*������UoT2,��c��jϤ^҅3�Jm��y��o^g{���A�,g�\64�h#]ܥ
#f�Ӛ��qL�(�Ұ�E�b�Og�#ko���Ԧk8�+��H�ZH7��}M�&����IQ��X�tugn��w�Y颯V�{����P�W���1�x�$�	���$ҏ�4���G�M�{����b���v$^ݰ�fV.�p�*�;	�Uj���uY���|jVc���M��3%顮�h��8ɾ�4sz��w�iy[ǮNs�I]!��k�n�ctT�:�J�R�q|����-��S5k)m����֝��`��2Q�6��>�!��}����拝p�5�\nG�2u����P4>:�8ϻ�k�D����'G�tw�P�:����.y�0��].[6��ß%d��$����H��7�[�^����L��&���-�4���{X��s����Rdn���c^J��\��Jr�<NRʏrq>r#gx���qؽ�L��`O�������K0�ͣC駗Q+](W,h��Su���DtC�mX�e/6G���عz̫��%g�J�}�}�L���J��V׳s��Nt`�EAW�M����bu�3s�X���p�3�|%a�nӇ��6�$��Ե����T�=j��y^SA5�"���`5[3*�1p:�0��v|����� ���w�!X�Lڐ��O���\��lo:����zk�:�M���X�Nךz_+�y��g=dg�{��]�L�,i���e���W����ӡ�Ʀa�X:UC��(��1�"±L|�]�v�}tKU�ye�-%�1��wS�zH��aB$B��;�p��C��(�M��E JN�(�ږn�>����0L���m�{�_�N�R�����	s{�)#w�E�����k���ۋjd����DD4姸�t��YM/i�k�D�Op�%6�7s��\&K��}Y���n֙F�mZ7�h��9K���)W�s�)&����;�vYd,�����H�]A�G��W_m�Bw۞���s$mc�?�z����0�8LUƅ��6�'6�;�Y�8�1��q���8et\Iu��S`HW�����hR�|~XD��q��61�g�}"ॗ꣐ٯ:T��EVF@��kФp�9�ѐ��e�H�h&﫝��޾�U�5h3.3������]�O���*����#�I��gu��.�F��yϳ�u��ht^�~�,�%FxJ�7�3�΄aV��zilN��� 
�3ۜ�����*�����&Mw��un�s�'�t~��/����\"�(z��SŨ�]蘎V"b XDF���W�ao�;P�����V���������Y�}ou����箳P�
�I��� W�n[��(�#Դ�&s�l�����Q�nIŭ�%p0��B�G^�t�瑋�&�|
�t��{���]C-k�2�}�7��ϓS�d�W�WF�*3@'N"��c��NX�j����eN�kM�|r��&
��zhԳ�9$֌A]���%Эl�S�1n�����w+�[�Y�c��O<�JǹY�(R��ZE㢁�����~�G����%K�,�.T]�(#K���하f;x�W��p�m�Yp�fNڏ6lvZ4�J����[[|�� 2>j��oqm
��l>�(k�ٞ�T��0eF8��Ӭ�XV��m=�U�r�U&��k��0�I8m+�a{�G���f75!w��O�l{�~X{U�S=�����#��L��K-%�#��=ٔ-o�p���5�,���C�������ڏb�5�A؅g���B��L�{fl�c�|3!7���t�W�`�t����;+ �V
X���`�M�^��8�M��ǔ�n?}^~.՚��a	u»*�PKl~lQ��.��b�V�/T���<�2���,u9�)^Gg�GaE���c�,��xٝ�������5�K9=��z8�V��Ҩ��s� �x)��z�.9'��pH* �2�D��蚎I<_]��>ߜq���f�(֔�Y�k���%=��E_t�3躼E�
ѹI�lh��]�ܓ���IT��K(x���0S{��;A�\9�ewV��Tݰ�WN6w݇ �����.ً����0�Nz�Э��i��s r;���"9*P���o�����o���.��x��[,*��BMT6��r�j��X���1�XY&Ґ� �Q��Y2�W{fަG����)_l� W$H��t�&�B[Αeb�K'd�ȍwB�����"'J�o���gC��+I����Uٽڊ�O��ɺ�ɓ���<TQ��~!.�W!�<)E�&�Q:��D��ψ�����pQ8���lU�������p�e&^�^N�Ǭ��E�M�|���&���^(����b��0߼�\v���glX,WSĆϹ��(oJҦXdL�G$��\�7o]&m�:vǝ�UGJ�Zy�}%�Ơ�9Yt<E�į�޻�4�H��L�NϢeb3��oC���^mҘ䞛�z�����~x2��-U�Uf�*�wtlv��؇��Q�V+ؾ��1��ۆ��t��5�[�\�����Q���!���=/+>����2!�ٺ7�\�er�B������P����5��^�|}eSl�s��3�q�~�\���j�����p��ڏ*�����*�ֺ�
`�^{���A�*w��X��
�G��Us8�����ߚV&�_�	��Ξ8�xD�6����]�aednEY5�/-[X`�b�����}��[�U8#tG�����s�^�����+o�;Y8O#���ћ�`T�f0�*D���0���� �c�����F4�x�{2�TKv8��ء���ͩy��Nͨ�q1y5g��N�Ι�+1�X����P]n7�إ�n�˕����7�u� ���og>����
�����LӒE���w��v�����@wV}��}���V�C"ϥ;"q�z��>��z�εŭy�޾�|P���icl%��H�(���B:���/5��A����_��y�8����s�!��^$�4
OiwO��o�7ŉ%{r*�vM�^�~���V�k����pvȠ$��� �Z�g2u��|FiF����P�e8���#Jx֦�����'�ם�`3���s�o�K���*��=֘:�y�s(��T�fb����s/w��4�;��P�:��{��P�0��ҥ2������GP��27�A{ܼ�wȧ�	q�7c���oْ<�l���:����as���e�#B���K�o�9��:���断[R^���ϖU�^ۑ�}T�O��_Qj��ޔ�fb�Q�T-��H��n��.��q�s��e-l�)����Y3�u��/j�I�F��w�lz[q*�jd׶K��"�$huΑbΦ��(���W�.��q��g�}r�����9��w�ZGQ�=<�ܫ<y�&�����1��۩%J��x��JL������w,Sg����h+�'E���_j=N�^��z��ը�e^q���k�{�Z�6a�����v �꘴�n͎g�b�l��}ٙ
w5�G���qJ%+r%�M���!��+�uӰ_l�獾$�ҳ��������y�/�z�WV�\�HTN�t��ԇ����Ds��Q�<�� ���5�5D��g�䈌x�+p��_Uk�����{H�J��a"l���oh.�!F�35�	�C�A��1���3�`�|���rN��L~�rϜ2�<��)�5P�;ʌ��n��Ƽ/Ŏ�<�_�(W2���W��T�d�F�q:�W_mU�K�S��خd����������C=׬���b���[��u��1z��R���V$p����*<���h6���%{S :K.o��9ms���G���s5��f�*P�"�aFi���;
G��AX�!C��� Fײ����ݯu�����CC��Sjj�H;�w)C��*�O�T��{;�k�0��U��ƷG`#N"����U=+�\Xҙ��v#M� ���H��i��"��\���ib�)�8,��;�lQ���`c��^)Wq§ =8��/�ҕ�S�4��Dy���q��۱�͎r�j!���yX�Xs��R����+n�	��{.�4�7��a'Ɲ8j޻"��+�囻�[�:���}�i0�k!`
Ό��O�-�����l�mɡN�YTA�̺��֧u���HI�k�X6�wPZ�w4��l�Rl��ig[HN��&X�b�⺸�>�[R�۬�Q=��׭�hԽ�:��q��ҕfbZ���=zq�=��f�:_q���7H���<�x��z�&���Bܢ��I��8A�C8
і�ux��5��fmfa{
ھF�c�|���X(���wF�2Dr l��q�1�u[�vgG-���LV&���y�KiYr�>������ٗa�@݌v�Jh��a�!7�^N�e�ǗtzP���m�3k�=���B���;.13{)J�N�Lx�{���~��n�.�X'�.����d�BL�;-n�.�U�Z{��]*av܌d�V��f����k�!eA�^<�˶m��d[B��`<�u��)��i�P���zr_`C�_a�ĝ:���(CqӬRm�j�j�R�N�9n��ب�m<��;y�ٲ�u"�Wh��[v����{"��7h�V�47It��J۔�=�Kk]�׌�,��=��}(<\U��b�̭�,�Z�,�zzX\�5�c�����q<�1��c:�1'd���1��J����Y���3@k�Ot�Z��J`ˮ�*����;���];M�]�i<��s�ި�ob΂�gi��݅@�݌��	z��-\��9J��ܗ�'Cf�pMiH���sCk��jڲz�p�5�>�k�U�ݡ8S�Dx~���Ae�1����υCgQ:v�<T*g8�V�}�j�a���'�3x�\d� s�\���aiN�e�W���t'��
��˛��%Vcw� "��2�8�NG�m=�U�N_	8�����ܻK`�2Tv�_
Z��{enB��
S�C�D��Q&���p���]نNfoUZ�#Eʲ�q^�U+S��;��<��]�p���<wV���:�TQ-XyH��}�c�Į�������F��+��hʂ�T�%eLɭU���GEe�C�S1oW'3���q����Q)��Xd���r�0�J]=�.M��w��1-��Lc}y�	H��w��X��q���wӈ��4U�4T}�2�,�A�d�d���*�è+��^^q|�g1��ރNk8��]�c�#"�uJnk5�fA�T�Z�<����y����"Gol��G�7�"��ڄ0��8\��z�^�O 2�v���z��o0&C��A��`�j��Wi��V�w[0�Ioz�m����e���C��#S0�ղ$���}w��yל:��4���:����#����[�jb��Kl��ts-�d�5J�^o��`��5�_J�qF��}���i�`l<��,kgIx�&\x�Lb�*�e�b��P1�s1J�*b+Lb��7�1U`�X,1�+P�qPQ`�&F�IZ���	�m+��AIEE���"�e���`��F"2��E%s.V�e`�""��%AeEQ�R�UA@X�f*#*��1�IZ�C�)+YD�)0A��Д@F�,��q�cJ��Q���hj��J�+V#V̴�ieG)�Z��*�W��Ac��%T�lR�(�*���+K
��#R�b���%J���X�ª,QQ�PUU�J�E�`�V�ł���b(��e(,��Z+""�T-KdQ@1�T��iX�F(���"��Ƞ�1�fUV
1X[�U�,���H�
�����5���~}��dԫͭٶ�{K�B�5JvfV�� �mi��=��f�o3].tM4���)�y7Z�mۢ��8�'6m�(�Q�8~��7b& �uf�.7��@rv�G@q7WrmK쭩�Kٙ��/+m^W�d��`�h�H�_��|�\B,�n�{=H�d#��_j;G�^�����枤��TK���5ƅ�g�+-�(�!l��+hIG���a�j��^��(�y���/x��xG7j�_ڸĝt�M	���7�%	^�JR��R����eD�o����Z�+K��6�]��l�^�wp/�Q2�P�Jc�Y55�hP�񧤅��ɽe�ܾ��Ii��0�Ö�cpT������U�V�~�~ퟄf~���-n���6 ��{}5���/dIκ��%n���q�[��K�<�B綣����{�9�<�l�'�c���*3S51龜��HOya9᪔��W?����W8����_�ǈ����w!���un5�X�d=���;.|�c#���:xT�1T�%��?6)�����;�m5~ܭ���)�ho1��r)U�hS���m��;(<Ej���	�=5u���ݫ���ZWt_�_y�ts�7�7e?
mu�Y��:2�[�Ws����z��nP�C���\���+�;�ڽy�U<��m��s�K�F�6��R���r$��9Y9�L��0�W^M�4[ۋb2�VtH}���/�6�R�Zͺ��!�WH��2�]�w�e�9��'�ܩ����S�f���K�Q�w^s�Dy���/�{� O��
�Fw��4�G,�40���RQ�e4�4ʭ���Z0�u]cֳ�.+ zt����P�����c�Y����n39�q�u������:��(v�*�o�,��y�\X�1���bb�g�'�V��g#܎ۛ��<��Qɩ�[�.>2@C�����W�z�*�.�C�����%��Wb&����p�:�!��m���Br=�WV"��2��9].����7��;JL��yH'`��PJdKZ��l���5�d*� ����HC�P��+J�ea�2�UE��;���Ew?&V9K���Z��'t����9�U���^��\�s.�=;#���ʰ�L�F����յ�S̵�j��,�z��l�P��������X����K�W�|�`��{�֡����l9'oOv����VD�0��7��{�W<�s�|}@z�ȯk�7X���T�ev탛�S�c�g�6�=#y�!LE�<�t��O\����v��B��^�#q� �D?]��v���:vd-]-���S��-�b^v���Z�En��0֘G���K.�M۹q9�v�vT�j#3�:���*v�=�J��܂ �e%ܮg��6�BDF�����І�[���5ء�ef>2;F�L�=��JVΗ��;�F�̯?f5ѕb{�a�*�zu}Qmh��U�iq��DE���V+�䖚VL1g"'�=�E�Ur8���������y��Co��	��U�+GtZ�{dx��Ҏ;ۥCkB�o�ת�w��[8U8q�f�m�ksֵV��盌�g�
��!���:�f�{�Y^QsÖ[�";V8ՅŃ7���U�E���1fiM�X�@�{�n�ޥ}]��3S7-����H�(����u��b�f�.p־���c��v�<��I�_Q��,L��j��q-W�$�:M�|T_�e#~��s��H�=����{}��q� �Ӹ=�b��i�(I�!�e2����(��@Հ��=/[|^u�1�ڗ�Շh񔨇��`jb�9θYG�q�|b�� �Z`�Low��yY���vl�ZX��Zg��dJ{/ub皡�5��6�+$�LZ�{=1���zR�o2�e�(e��w��Dy_��ٜ�z��ג�7�q��׻�.��9����9=��s�S���z�'p[w��|�LP_N���]�	f�SJ�k&�c�ķ.�2��&>=X�`�.�hd��O�ͻp].�����nD�[ǹ�ݾ���"y���o���[$i�(v�A��,9�tE����;�23S�:�_^�Kmr��eD)7�3j�O�@�:�]J�crS7��0';h��L�f�[�I��5/����z�o(C��42�\��g;1��H��]�.R�p�O�ߕE�����>�3n>h�w��K9b(4�A���"�cWD{l*b�a�1���(�׹��k�b)5��Ν�b欸���Fys��/'�uN�M�rð'W�}i#k�����i�����z>yZǮ� v��cv�(�3�:�珮��^y���koh�}:�^^m�znS�3rs�ׅ�.zE;cƀkbX��s랡�c��0ȷ�S�����K%vS��o�iL���V�r� �`�W��D�Ϯ!C;�zL�1SX�Y1�'�jqc�ֲ�3�:X�<�ţ��.�����~]b��� ����:�:����_�W���޶�U���u�璥atޭ�����$�{uA!\�/i�>@wyਖ਼��*��sv�vh��/�}Kcj�v����n��Nѡ<�	���E�Y�V�-� +u|V5%.^]�Q��ˢ+!9G��ʙ���Ǯa�B��9I��ƫ��rD�d�{�H6P�9\�P��11��A�,�����y�`�;%���%;��1�(w]z�>��z��� \6hJ�<EV�2E�hr�����>�:d�3^Wj�ے<��>cn�.��@g1F�Y�b�Y=@�=
,9�5��U���l;5��������=�� K�1�WI�!�T���(�WE�M���A<�/FH��e���Z]8�j���)⨈���G���
��b�;��#�(.��X<5�ObB��q��}��'�4��5��TD��D�U d�"�#��/EUq�E`���\3�[�0�`���8���(ϖ;��R�hq�D"��#�G��,�2��_�n[��{�a�'z���V���}�_��Y�L��+R�c��B�G^�%�Q�ɤ4p��Pg�]�:)�c�.����zNXV��șC+���v���\bO������o��3�y.���ٜ[yi�c�z��{y3:D�t;���=�vEﺉ�r�WN�rk
аR�;ڛw^Oz�y�f~�4ߘ���U�[��F��~U�W�����l� 8�=��(%ޭ� ��O0s
!ygi�q׺x��Y��r�,�'sW�>D/@�CR�t`�67�4�[��i.�St.��#F�5F7|9OD"Ek85��i�\p�m�`���*Gq�%�itom7*C��[Ӌa�U��N������1p�K�tu����pGOg���
��!_��	[��xW,�Z�igRʡ]��Wk?w\��nH���'�P{]D'���b�X�O�[A�^5ؔ|�N�\ S+�_7��f�{3��CJ���{�0ٝ6_�_�� �����p���͊�}����e�Vu�����췄��DM�6!c�ȦJ�ø�/6'��;�vP$3�V�����a&�nn�j��T1�2��G�@�Y�sn����k�RuL}����;7 X'�z2��;;��;J�4l
�'�T��(.=�a\]U��g�+��&��spK��WaN�9���P�+�<R]��,��2's)�����4��g��q�^�.q�T������V���"W�Xw�ͻ��H��=�zK���>�@�v��:���+2VƩ��m�X���팇�q����lP��5/n��W��D���]���y�w{\D׷���V��l~o@���էR��^�##('v��\�"���J6seI��yT���{j��l�f���cVU�4��=rFD�$�Tq�����rE� &2�R �݋pwz��c��~(:�
V��ܥ[�_��JE/�i�������,��yb��̱P\WY������ru=����TW���o%:�����r�j&4�&17:ȱ@�U�$*=���砵�ˎ�6dlB=��q�Σ듼`]�WN����.�`��Q�J*H��ˡ�P�X��z=5#��ܝ�n���F��0^o�o�l�x�k�>>;(b���x2�k�pO�-U���+�g�fn)W��D�W6��s<bkܺ򮳞���B�"N�G��
=Ň>�y�Q�6��Y���8%4g�6�;�!���:6ٴj�DD�����І�[���Mv(E�vVm��c�h�Ét�}/��x���xܪ��ǵ���3�Ճ"�ڨ��T"6�=Bb�0�7F^!���77��5c��������茹z\_UW#�UU�x���a����>݈m�Nj4Ox
[�==��G�aĳ��SIf��d�@�N��!v���NI~�[uUCF�_�;���XĤ���z������u� �אw\������|D+y�"�[8-A"y�9�rC���t}�����|%�QTy�� ���DiƄ�vB:����{ޝ�8���42��������{/!�6�rWu��\��T�쭡n��q^7�.��!���i�ᨣو���9���c�7j��ʒ;|=[2�����%�到8u�SL�|�Z�.ff�\X���yc/�T�l��[��Ѿ�dNof#s�Ll�D�Ұ���)�'��,�� f���Q?o�G��g����Vr��`ǥ�j/�ōa�Gj�ez�F�&�܃)j���=�(a$�n��gS[ǻ&o��>������}�m��$d�:�f��.7#��B����*�{4�ZUY[�7�ЂYۡc�{�B��{/uW��3��f�۸}�u���yBg���g{�#����p$N���{��}l�����P�Q�5)�P�[�UXH�eҬz�5���&���w鶴ҁ�C�~��2���}���<\��N	���}���U{����.��.{;�(��I���b+ͣC/�40��j�{T�6e.�?�>sYQ�!^Ubn�9����\�|�r���9�u�j-��ɯ',E��i������M�G�3�1OW����~k��;��L��D�֜:%Vo��}�`S���:��	���?N�6��F��^���93� �W3Um���8C��؀�,���y�� ���~�D��6���f���[�]Uc�=N�9��EŎ�T^V4�wF���N����y�^X���#`P����U��wx�����fh����B�Pۙ���:֑j;lF�5�8	���,��퓦e����r	b���]�G�5aŶ\���uq]|�8��4�$��i5#� �d��(��N�U���e�����]U��Bt���[�J����f�펦ｳ6�8dJ��j�p�Zкã��gcU^�nU��P�[�P9^�G�C&�5v���O���;�l1��GZn�E���ΜY:�X(Y�W�5ӵ̑������Y�����'RG���0`\}�ñ�RG�J��X�5H�R�x��dq�ߘ�-Ӑ�_�j����izn�����	`�)3Xp٠�R��"�aF�di�#�*<ƃ�ƫyzcW`�b��7y���5���^%�z�CE���+����aܾ�5޵�	��JF��dѬU{�r���"/d���
2�quS�R����zS=��FmP1�OS���i?+}���0��f��vy p�u�6I���<"�un��Ș��=j��?��ο�M��%)T�$"�;h�X��2{��Bn �Ӝ��\p[�	Dw右s6��ym��ƤW�b��w��K�=��Yτx(3@i�,�2��X#r�z���A�=���m���V�\́wq����NCLyo/5NsL�Ie��Ps�ƳJ�����Y�����P�8~DU��� ��t+���B�A#����V�ݬ��Af�4�Ξ�e��)��]�%%,�����.\��圸��ؔ� ������MS�%[s��E��47�jS>1���T.Ď�Y���d��X�zcH��s�Ο����,he�f�˃+���v���\bN��P�^�D}���<�O+���ށ�5�ɝǷ67���p]�υs���
�I{�뚛w��T��<���>KE��yF�ە�mj�d��F�9�C��x2ڨ*ó�.��](�G����x;>x����-����������� ��!_�m��l#�q���[��'0�]Oc��9�;�&N�[x���يq�k��|e����ŀ�F�����㮕��]�%�/��WlV�mk��9]��flC�
%k��uUv�!�7�ٚ|p}5��+�0��|�݁:GD�Gh��$��>̵mٹ��q��c+Ix��5�����R>�>���Qo_\�g�P���)a��|v���}���E�}BX����@GW�ن��`?�y�E�o:��g�'-���S��Yڽɧ�������uYW�W:en����7P�.σy4�*2��+�t�5/�8lᘞGM�z�W.��DTG�x����j��5ə��k��Ic��d���rcޣ��}:�_e񭽮�"����G���t��J��n�Wg�K�`����)�F�h�{%mc�+S�ՇB�O�N�tx�j�^��z�HS�7�!�P����]��<޹o��.1Ș�j�S��
�\��p�z"�6�0G%ܗ�oV�˝bmsӄ]�����ft��HR[dp�& �B�u�`z�*��t�F5 �(Z�����ᱥ �S��A�Lu��1�Db�f�����k{�8������֎4l�곚��͗y܌���}��������s��t] i��B-���y{�f���f�đ%��33)v��l�2����%��GyHҭǪ�C�T�ngS5)-��� �Z��yKWG��G�`E��ۭ�9{kjQ��2�(�Da�,O9v���I�b��n��jeZ�|���[ެ����5p�3fBZ(�ʣ��)2_׶���8{EmНN�	k=Ea�O�=A�e�s�豫1jo��s-��W7�&F�B�����SM ��m�J����Փ���Pu9k�F�p�SRߊ�΢�cT� �.��b{�����L�aû��N������1�F�b�>49+���]N�{*uH)����VQY�N5�����>��W.��ϊ�����m�j�8��p�,z�ċuǮ�,��P�j������,B��B�6f_9�alj誽Q�f� .�:ʉ�Ԣξ�+7y1�#5�=`���c�mj�7�Hj��ӣ�4u�v�#�(���]�䙘r�f���
-�$b��Y�����b p�*B2��3�'�T����gsح��.�-��t�%��:t��f�R�X�܏eHw+���lT&
�*-6`�͒�����C��������#��y���.��N��pŇ�-�5-6��p)�;��U�@���Pu�0^�U6^�M���,*�m�5�����(���|�^��E���ҩ��w*ԝ�C����۠�K97�P�J��Z��lM����T��� 4����=�9������H�C,��,�J/pG�+���**����d�%+��me��w3E�1SY+%D�x]��5�T�7�X -
'+z��|�+�3rj]nN����=z���л(:�x�&Rl�l�}�v��݈�i�N�r.�p:���J �l�����7%�eD�oG!�s�`�(���Ք��G�K�7#SL9����2����.�d�����Fl�'E;9��I�W�-��=o�r�Tb�8$�K9�w[/��p�+T��gvq��*p������)}��׬G�.b�C���2��G����]nY��[gi�a{d�s�+���
���@�D��v�b�_j�J���Gui.O��v����\�ZY72ʹ�%b*�����jB��PPkJ�+Em��Q�����AR����TX��TQr�jŊ*�QJ��*�ܴ��J��c-�QE�0fQJZ-eEDP�X��B�
"0PY��#����P[f5(ܷ)b,A��e����)+��@��*T.W,-"��`Q*"9H������%̸8ثR
,2ط3�Y*-���D1%VT+,,LkV�B�V(T3,EmfX���q16�"�ҋ�cj���P��q��Z ���n$,\,����k((�Um**���A��"�Q��WV(��1�b�ډc�X����2��2����b*��=����)s��҄LA���G}��s"��A��g�eE���Y�x�{�s$��zN�<!*�[�Q��;������q�;�'�eԄ�t}C�1-����
CN�[��՝�uÀ��~�����
��:�(y<����b�6�/Dq"7끓�i�,�F�_lT��Ɵ��d�U�ıW�m���@뙟ͷ
4�gcq:�r���������
��5|Y ކ��e�^�k_ve΂Ϩ��T~��SV���(�pt���
;�_;�\�Ғ�j�g���՝�K3��B	`��%�i '�X��|���S��2㢍�U~��Ld�b�a{����Z��L�36}�,k���j�[��;�U��̑�COD�	$�l�ԧ���t�2��v��,�a@�9��ꎿ��φ(�x3�6��f��#��Қ%�;%������VR���C�D��n��lF0�'S|}_���y����ɗ������;�6�]ݺ���[����K��y�*�� gu(�ܦЯ���y����j�E��U��s��d��:�T;^���U6=�M�&�2�{�a�;�U~j�F�g�Ll��]n�r60~}���B���mm��Ѝ��>r�����U��JN7��ڛ�D^���������^�颇'�\��7��ɱ;�K��vļ��$��:�$�%���eqj���N+e����Ye2��B�+oev�n��a�q��f�w5-�s�*�7E"c!�`/K�j�yso�����̬:&��;����~��@���{��2w�
�V!>���\�1���\I{el\ۆ�#/��ǐd�q�h�lz���%�X����`��M��B���Y~.��5���p�7�L%�����I�k�7����]�߄�jf���EQ�gBZ{#M4's��Gv���bДK)�#�!��5���C�nzN��(�ǙĵX�đ���U��b��S���ӎ��1����{%af�*���Q�p�ӹ���UkN�&�܃)j�D�Lp��'�뜥*�;��������E� �偼V�7QBڷ'h����ͩ��kd��t��ի��>Qw�X��Z{ה,����V�4��q��A;w1\���
7��;��R��fVI���N�=����2�#K�,um	���5)��Yէ�+����&L�CihQ��Y.�&4�?wx���?EMv�>��_��$Q���&��j]�u�z��dXU�<t�LZ�4Υ��Uy\��NM9���P��u$U`�Q��p��xlm�FA{A����P��d�s��2Ա˜'��7�|%6��㒳~;y�8�-(���._{�ʮ�h�Z���r�Ꮊ<ѹ���n��ޠ�j�KTQ�jNT0ą��ua�-m|e.�?��b|�d�~cH��(j6�=�@�u�����+5�|�ד�"�F����H�a�:��X�.��V��Fw�j��'N�E����8L�N	�f�M�@R�^�a5�"���a�ٙORe� ���=���Ild�C�,7Y9YC��=Lq��31_��D�L��L����
!WU$�ɦc-�Yw�����F�uv�3�q�
(��o����ګ�Zu�S~�Ⴏt���)+��fO��wX�}��]j�*�^��p�Ԅ��GO��v5U�6:�u�#^\fV�=}���R�ץ���!�3P��7c"��XV�XO@j	@�림Ή_>@V�Y�$>o�
p9yo3�ԟ����J��!6��s��d�gn\�QD��)�"f�=d�Ә�f|~ﾕ���MN���C�,�>����p�^t�C�Ul#�,�;�ē���G+y�͹���0b�P���p�e�:h�(��;�f�8v;�rxs�~��N��CtZ������E[����A�*����t��Ig����|3ȁ�lh&��l�Zot]�e^�R��r����gG�+4֓�˨O�oeW	|ev�ީ&S��{�pa'�,m1��O�qRL���%4z���m;���h��6�i�C��)�N�*�=��<���W���v��Vj���JL�Y֣�kS`��n�F���~�c`�:��IC���@�^��R'y�a��&�l�q�g�z����V����1L��6��ԉ\�$�,�B ��^����Gxj�z��:��Wb]����/��,�#�8����R�(�� �h�H�X���\B�Қ��i��lw��K9{}C=H���3[ҵ)�0�v�r:�Ac�ՇΒ�����M��[��잹׬� Sh3MMYjș���n�]⡓5��8�j��K�9bJ�5�O���yȢɹ��y�<�����*���d*�뻁~�U���$�������C^�Ӿ�֗e��7XV�o<i�a��-zk�:�}�S"��������~��k$�/2�7�*�[�=7�����5=$����͠���GE�8��[��K�����Qy����w`��>�w��kB���?,��!	�VaӘ�>?%�u�~��Bfⴇ�ΝNQ���Z���]�(�]�~�"Yp���	t���s�����-�M��2d���w�A�lm^olR��N'љ}��Y�8�P�5��r���5êl��3���}R;V{)Fq�nwo)}NG(�i�c&~�����k�h�Oj���A	A%��5>l���_�+�����L��v?b����p�3O�M~+ˈ�;�1vG������{Ѧ䃅?V�ۭŗq��]���r�̅%��t�#��v[��1��ˎ�N����E�������:X2�m��L���\��o0׼Ȣ��wNO��/�dӓ���h�a^�z�����K*���7�uR{��T]�->T1CF���;�x;p�3�5�����v"���;U�1�p{�B�J�ޒ�(���}M�ǂ՝�����&xs��d��Ok�m��!F�c\�	�M��۸�Ĉ�.Ou�����������ѕ��oEKVz�:�J)�VE _+P�I�v59-ˀhK۴Fx7��V22�Q;\j�UVi�u�[����Rb#O@"�Q���|z0��e�0��p�j;�_;�C
o�]c�)�[j�i�y#����ZE�!:�ć�oG�Xe�l����{�LQ��������dO���j&T�*<K��
�є2�(8���n�ߣ�0-��o��D�k��\����"���J��#I����/���D�*���g����ga&��^X�R�(0p����gm��ܔ����蓝
�TQ��s�Od݁,�j��,y$��MN>�u�a9��Z�(VS�mt=�H�wv�u�qԏ'H��ti�˱�=S8���~���:�;>�=��]�!�.��]$�6xN�I��5�2���;U��R�:68b��DP����F0��t&�����G������?�β���r��`��N�߾�ށ\�=#��tSٴj�DD��d��)#O�
:»=푯\�q���-�d��ξ�`�z��׍���*��5W���2�{�a�g{�F�N�O�e'~/MkZ�ɝϻ�0��6�꼬Rؑ��*"n^��Uȩ��>N��|�y>�瓲�~3y�>�����+@'cH�N�ڼ_�R�f���8��/�l��fg���~|�i_�0���O�=�/��b�����
�J�¢7���b��J������~��u�'ו�ܳ�NȖ9mf���Lؖ�EQ�gBZ{��h4's���Y�j�^\��j\[��x�.+=��	�BqB��9�KU�I	i,������J/a6&h���3�J�cۙ��n�.[f�=�*���P��G@���G��˫��x����G�]vіpde�J�����'��q��k.H�B6Ν ����w{=�Qw�U�8���^���'���7����C��O�p���0^Ɔ^볜��rL�K�\?	��Q}�t��2���$���z��S�W�wRVb���\�7�p��)˟J���׼���~j8���J��X��rիЋ�'~Dq����CA���yB��{/u`\�T9�,����];�jx�"�oNL�V���l��?��'_ǽA�{��}l���xXU�A���ę�qm���S�֔Q�Ү���=HY�*�,���[L��e����/��¾G'��Ո�Q;1zk�>�Q;���1��%�"�F�Z�&������l�W�{�'�N�E��s�������5A��ZS���Y����&��"�H�5��H�a�{�#�s*��E�,��V:I����D|��|�Y���B�Ṿ�E���I��)���C���7��uYچ�%��{�ٽ��{6F��?11X#�,��6*�1Ɔ�f+�D�ɷG�rx<�cطb�^��?{��-i� /Xw�Y�U���6��@�=��V��&�$�	<�-d�k�1w����٭�u�]CC�1�r?�|���>zy�k}�0&�����h���}gum �VLCe�k-Ž�P�=0��'0�"�!]h���v1M��y�� IV,�X��K[=Y�	�+���E�$/�["�3Z�Y�C)�w'�����(�:����O��#�bRيu^*q�T�Zdk}��dn�8��:�`��y�1�7]��SL��Qɺ�V�Ӌ'I��5`�=>k�����0���^��՛��vR�EKc���la�9#���c��gˀt�(���_I�sg��;�抻կ�� �ȱ[1�j`M�g�/�Rf��l�t�C�����# t5�+_HBZ����Mj儗C^8�m�LC@6���.��C9�5��;�^<��B0�]�ҖM�v`����c��ܮ�Ka��N��'�*28D��P!���L�5�Z�u��]�Fi;Xn�J�$�t��kջr"���b�i�m�:���Q$����eE{c�D�k�����x��ٷ#�v��\���G�+�r÷6���P�2d��$/�XD�uf �ӕY��jc\5S9L޾GA�]��Tv�g�9ŗ6��nǰ8�"
��'��Uw{�\ܱ��q=֠�0�w5�l*�mT�D��Z��v�bG^�,��\`�YJ���y[�q^��ȳ�d�4
TQ���3MtYaY��w�uK~��������CZ@`¶���3VRG��'a�����X�O�۶��(̤��3z�G�\ZRr£��X�=cwP����[NP�Q�JB�k���+�`�ԫ�Y*[[Y�P���)aQ~׫�@�p���-U����X{��N;թ���
5�t6��)LNl}u��3���^��F���^uq�Y��u�zASs�pK|�ٴ�@u2����{) ��@r
С5�On*�9`Z��ux�)�#<����b�S���ց��:����3H��x@�-�W�V�DO�U���b~J��-Xk����������㬀=���U�Si��s|�{1�d�Q�zU�t� Ϥ~K����~#�h���c����6��E�
��<��1����3j��?lο����_�C�����;KG��HPf�ٝzs��eB�!�6F8ɛ�����﷘؅��l���v��sb��P��tr�{fo�[=��!�"�PO�%�Nj�]B��C�o &�"�V��k�;z�=S���u��w�ȳ�[BGd�)� ��!m�7�4�F������yے83�NZ�[��*�Xp�c6�#I�a����X�����%�ޒ��c���iѡ/vq�%߫�v��,F㼽9�ewV}��Tݰ�M�� �g�B�d�XOI`��?}Kw,��G5�<Y����z��^�9����mLc����!W��Z��9�Y\tv��%�)�Z�.��gV
��)�0�b�F�ovjӒ����0nӥ�}3��,΀Șw?,{��}�i$�������E���AhW	C�ze��Rj�y��D����rr�����?��M�rt�k� �ln'Cb�p�۴Fy�Y��`@l�i�k���W;=;̔�?@0��;?l�5i=o�t(aΕP��w�R�FX�\�ť��<ćJ/�)�H��K���C�Չ;�ޏ�pSp��t��h��ک�ǫ��A��mP���mjew=*:;\5�cNPt8��ޡ*����z��L��k�54r�=x��Cg*�q2��_EKk��Y׹�X'���9F�5X~ٽ@�3���{�v����:(C� HiTv�#����Bn|}_0��Xwʦd���RmT��|�I�G�\mmU��7�-"�k��ٴj�DD��d�>�dB�[���ث��t��L�MKg��bT����ڮ��UC#x��P}�~�)����-���z��R�.e��M{����] �]���xc=ćg�W/K���G�U{^�� 9�Ҕ����������%�j����o�V���q��~ט~7+�{��}{H@��	!I�0	!I�$�	%�$ I?�	!I�@IO��$ I?�	!I��$�	'� IO��$ I?���$�	!I`IO B����$����$��$�	'�@�$����$��$�	'�$�	'��PVI��P�8@�7��X���y�d���g����p0 ]���
���� �)�Ҫ���AAP�P��     �<M2�J����     S�IU)=L  4   `sFLL LFi�#ɀFS��)U@ 4   h  ѓ �`A��2`�$�h�i0��i0����Le?S)�wt� #�_�a�Ԩ��?���*�#���Y_��؟ؔ�:�d�n�  ~b� G0ZHH��� :@��iο�0�'���<�� P`_R��k��A��薪���kAAE����n|��{_Z��u�j�Gh�p��+ w(-NY�J��5Ţ�ER�(%٣y�U�y������X�]lm���+Q�U�����U>LT�v�J�Y�hխ;�7f�k.fQi��gM|�*{�H��H�՗�rt���?�3r��7l���`�+k)���6�5Y[�����c�u�������1,�$�P�#
�F�P#+F�\���Y$V�cC-lӛުV���2�
�������ܬ�Y�Wu�K3t�CI�b̵�Qe�x�E���rm�6���c
������U�k2e�L�ٹZ�"w
����V���'E�"wf��@���%�w3sN	�ؽ٘x�U�:�np������*�`�gWJ�ذ��6�x���������`%�p��2�#'J��Lm�kcc;�ղ㪱s�w��tJ�9[x��zYʝ�5oq�mK²u'J$۪�l�h8/�
T����7-Rǘ���V��hm�R�.�&��ڳطY�v��A�cJ�Jm��o`���˗F'$�r�I8]jmW�71*��e�⣬��)V����\��%�G-�[�)N]y���uز��5Y��̺��d�ح�;b}
�C�k�+��̾�����T�������	Y�yŚ�mf)���n0O)�ea�]:z�[٫^�T2]��	ގ��:H��Q���w:�S��ĪѪ�A�R�EUM��gv�����p�,�N1COm��y�ˑJ�㙈Qx*½$�|F�V7K��6Rۣ+	o����MN;�m�q��-����A��2��Ŕ�jq�!ʣU�U��4a�|�ppQ	�H�U	�W�SCNO�%bNإ%*?A�!�(�&ݛ����um�ؓ�hП8�˱i�@�K��ITm��,!�M�)@�t�Q�jD���%�"���(B!e��+�KiZ
�`���7I"�j�.�l�dAEO��dYFY�H��$
(��I[)�A��8.;��}dB�D��B4%��w�-AQ#T���f���D�dYT��,*h�(�$Q�B0X-!-RDQ�Ԩ�e�J㒭P4ݘ�_�&���f)&
_Q-Y�B[*�dȅ6m@�,��"A-P�BER����ʭ1�a�TA�$Y>hg�_}�;돟���_�y��r�!���d��[h���t�7%�*��fi��n�V�7D�P�V�oi�����1凂�aFE9tFD8AS)���|�>'�E�l�=A%靻����Lb �z����b=c���G�Q��o{m݉���{C��7y����^�FP��Ln
���Θ�ƞ�b��}�jh�R�|�6�\D`5���zx��΀:�����Fz^ ��ý��%�iICP�n�ś�#�x��+gv����)Y�~>�{��S�Rm��Mn"�� �t�t^.��,��[׋Q�E�%��z5tY߸8�YT�
�{�gv�\%�BZJ�E4*DV�*����:۬[�\eT��]�[�*�wnmc�f��/�>1��w��8oX�$RK��׫-�DN��*���Բ�qN�u���q�}�����\�𻙩����;�"TϦ��I��e[�Nw���À̮y��u ����q�[թ��ۜ��X����Z��q��$}d�]Fl��ÍDw��*vg���k�bx:�Ӝ�����fδŁ7����4R&zEt,_��e���	�X��Vy����he(`�nXa�W�5�{>ܟ;�ѯ�҅�鹷^�˛��]u�ƺ�(�F��k�G�~�=�ގ�ܡ����.��q�j�,�Ǉ)�}�=�fi��4�_!�9�LG[o���:N���k�S�9�/�`�7<�9_�/6����d��l�Õ�NȺ\��d�'r�Kh�}ú����)퉴�;�i��85-dd�vK�Cf��SQq{OL����״���ߩ�����iw}���m�_�)��\(���"��:�Y�h����E�:H��B��
�Na���w�v��l6�^Ѱ��|�$��L>�L��cv8s��������cA�܏|�D����0z�D��yz�L��Q{8����z�?y_��u���v�f�M�K�S�*ޫ��ڳ�XR�Ҡ�-�K��=.�x����;�y���upݙ;"��;ݯ�Q����&��!ۓ�5��4�Pb���G 'y�2f図�3L�*��U���@& (e,�faۉk�6@�SЊ��o\��3�s[��f�sF�����
��
�#t.*���M�6��O�{G'y>-��/uE��nR��I���-��=BZ�)�ON�s���#�6��������o2�h5Y��������b�B�w���`N�+�Hم�7���ǔ��2#1㤟F��o��w7�MCZ���F8W�Z:��)!bd���	6T6�f
kR�C0qJ�w�����*i�gȿUgx�c�3��t�@�Yۄ���]FE��{/�r� H�"��?X"@��.�q�i�B�͢�w�A�-��3 :�3
Θ�4ܙ��m���uv�hU� m��J�oJ��7��x����1H��b�)�3H	}�6�Z��-�:ժ_kk���2sA�\Ev��w�b�����F��(�*`��B�j5�@s��v��Y��@	U����\[}��3�ج���5ރh�E7��	�CH�`�*f:DL�8�K��Ve��W/3A���#�4��G/�U�V���1|�΍����� <E	���N�:�M�W��SީTF��u�kX9R�co]�D��JD�KV�e7��v��KH#��GT�^��#菶��U���G(���k�8W��Ew]�`B���ސ��Q˔�\�@v�]��+��U�3<�hV����ZBc]+ry�������UW��v4v��ol��cO��ֺ�O�;ɘ]9K(z��gJݥ��N����<L3ђ�-L��̬��"gb�6igN��w{wa���'������QAa���"���WҹWg1d1�m_[���w�����^�A�����x�9���7�������^�T:U>�O��Ǌ�jvX��	���1�=ګޜ[hP����!Rf��5hd̛B��b��%�Q6քsc[%Uыg���<�Z.f�lC��
P��\8i��rQJ�%�M�M��8_��5�pN�����'ł����߾���:w򜤏L��*3~�?G�&臫�l���Dvg�R�������D�����虻���Z��i�C5�:�;�B��ܻÍ{�>��)����.O�<c��e�P���H����k�2�u��g��|�|��?�����5ű�yG�%A,�����Lr���}�D}�ǈ��u�?�����I���b�/�c��+k�Y�s��kR\���G�z��������Mdq����I�m�n������3.�H407�:�B0G΋Κ�|%���R�{L�;`Vr��fnf��G9�C܉�/r4Y�8�Z|It�)�"�gA�,�Ld
W��#L��Z�zD�4k�d�y���%ǾQ��X�.�\���hFǸ�{���D�I�q��5�-n�m�r���iN#yO��ڝ��]��t�:N���T �����|t�P�5ꪲ:���n_J����A��v2Ɖ�y��8I@�Z=���b�ƒ��3��V�ZXs�����U�rU����3ğ_?��Z�Z�-7I%��ѳ�6�����]w�|t��Bo�&���
\�ÉC��fϗ`h�8I�5��� ���ٵuGP�P�옭��:�\6���"�(	�i}0[>�j���P"�7�(�Gyq���B
��Mە3���0M4�7�lw�{d�l�L�=�Α�xuG�츮I��i<��q<��dѕ�����)Q��׹�/o�ZT~�PrCKԜ�8wlB���9H!��wQ-�P�S�lD�S���55�,@
�����" �{��!碲�z��/,����6S�Y$C3�ZHy�B#v5.�K�l�dS��(��"n���o,�f����HQy�Jٓg)�^_b��l�:xaH�_Q�<w��d!-���w��{��2ч����a�N䫖��>�4�򔶐��n����ӽ�<p�v���y�Z��y*�c)
#A`�.�͎��Y>>	Q�,#�zc�rg�R֟���z|��K^���~����'�����wSua���XQF�W��ҫ

�]�0_FU;qA���T�J6i&鋑�K_z�ҩܤ;�+;=]��4�>e"ߝ�{��&,��˚T
8�$3R,�utf�ԫô"]�/������4�u��Ijec��=땘V$�8Uy�!n�<z�B�U0�
�2��Q�(Fs��qK&a"�WQ9����z�ࣜ��6���V���a��f-^�5o�T�4ДiL�Շb��l����y/\N�u�U�k2v܌�����YY�����y���⹈��Lx̎;Q�2��Ɓ�Tcܐ���Ay#����9w�����S�������j1
,��!�HPC�ő�}¯��(<�K$C�f`IE���Me���b) j\�
�~ǹ�51h#Լ���G���pr@�A���l�GԂ�]������|�oW��Y䏆&	�i$n�<u��굵:�ē����I������n���=���Hh(����Ov^0�����
����P�C=�M����z��Ŷ5�����#�A��Y��/&6�����8�3\���S���E��8�9au�� ̢��j9����i����[�6����I�.�`����˙���v��ʜ-�j42����)������wYB�qn�e��F�'{��
���f�qE]:{�~�"����_xඅc!CC_�W9w�1)5y��+�.���)*�j�k��u#|�P����
��r�|rk�o;4�̮=j[3x�I���}.zny�D8;������8��k��f�Y޺yy��[}�Ӌ�zy˜WL�5�v�A���y�[��LR��}}v����9�}�/5�S;P�W7�~��?/	���^��:�).�w�H�&��<�B��m�"�1�z	�j+�\w��q�=WS� ���3����^	�M=e�1��7�����<������G�������慎m*I!$�U*�6�{��
�ڴ� ��}�&��+[�SS����|nX�g4fRި>�h뭬H���&� 5��A�s�\)kj��e�$�f�v���8㏯޼�[<7�X�1����b/6]\��:�~9m�M�A�6�uƥ��A�����ۏo{����E�vODU�vH��Ks�q�e�JvPv�C�[��������<Lo �P��� ����}l�|	 06�ȀX��@гF?�=��̯��- ?��
�=�Xuu����	!��s���į��� ���m��r��gNۇ�j ��"&�/$�큢�c�k�[�\�����?;�@���t�WCO�z�q~b�=}!#�l���upSc�������px~�(�~������ (>v9�p�ܜt���!ʌ���NF���_.�9��=��]��!������|M=}��xju
�4�	�gh��iüs��f���=:,! ��'px�(?���Ň\��������+���0�#���NV tt:�$�f�Y� u}�)��#���� :�3�`���a�T�S\�Cm�]4����=��1|�}l����`��<}{�y��TA��y��:�`vA���t��lu���kaG�����������;8~�Ǆ�O OaԖ�:��O��MD�Ŀ>j2{�|�=
�j�w�Ա����mρ�r<Ws�6��W aYbǾ����]wx�=hw�k��z����t���h����c���*�=�B��S��D��]�`��x��9lB|w�!z�n+�Cuh=����R"(?�������{�3_7o$E�z���D�/�@���1�h� �[S��x��_RC���m����w$S�	�}P