BZh91AY&SY�,�݂߀@q����� ����bD��           ���+��d�[S@�eM�ֲ$��lȤH6Ԥ��V���mkҕkJ	@m��"�ٴ,Њ
IHѤ�TTkbU�9j�eV��-I�ʹ�e��*[6͵%$�m��b��5f�h��d�YUmeY��1P��Bֳj���CV � ��Z�Ff�nX����p�lU��֎�sVƲ͙N�B�Z��ə�h�%��d�5���Sf�Y�m���m����mRաtnT��S��@  w�/�km@n����Z��N�В�vWm�kWf�wz�lS�`s�[%fSm�TwhՃvC��j�+]7me���{3U�l�6&��i3K��%( ;��N�T\���R�VgOo�A��v{n
h ��{�uc�iC{��(t^��/P�6��U��{]����x�ѡ����@Sw��leam��դ���ō;�T� o�G� (��8t���={�� ���,�*J�ne�h= �W�4Q�ѯn���=:v��(���F�k�� om����kl��m����f�CkE3d_=U(�U�@V�����
�v{��+� �g��Gi^���+���r���@8��:h,�� ��U��x�P����z�^� ��ɤM���*JX��IJ�}��_��ӳ���( ���=zd�A{���A�ݶ�������C��ܞ��У^in� R�oo]�J��:u�vࡡA]� Ui3U�mj�F��[愈�}�P�էk���4�e���47���@ b�]�5��ŇG&ڨm�NC�4��ƺ�����[�������i�4�l����6�L��T���>������u�w ���� =��  w{n :���k�Ű 6:�� ����k�� �rD�Z٬�5��U��a��U( sݾP ������� �77 :��p ��V  qܽ�:h޺� �E� ��  QWi�k6�f)��6j2����RP 7�� �a� �}�z ���(wV� �\ ]�n4Pt3�� ;�������{7( zw]i�m��Uej���-��h�>��� 7{��K��� ;Zܸ�G� :�����N����w�^��Oob� �w �� S�� 
�((M@ L�)R��� �h5O41JU4�oR4�ф`i����?#!)TP 4   h S�MR�4c d�F  $�II�P@�  �  �&�4�R4d	��2	�~�Ѡƚh����X?�����uZ���'� �K�ݪ٩�>�����g��:�ajהP[������ _�*�*�D>�P_��?��@W�A!���У������?�( *���I$����W����EJ���/������>����`[ؖ���4�KL`��6��%�-�l-�Ķ%�m�l[`����K`�ض��lK`�m`��6Ķ-�-�lKe�cضŶ�m�l[f��Ŧ-�-�l`ŶS�6���6Ķ%�-�lKt�[�Ķ�-�lKb[�[��%�-�lcLm�l0,b[���%�-�lK`[0��-�lKb[�6����[ؚb[ؖĶ�m�M�6��ؖĶ�-�lKc�Ħ%�-�lK`����m%1-�lb[ؖĶ%��1�lKb[���%�-�l�m�lK`�ؖĶ-�-�l��-��%�-�l`[��0-�Lb[ؖĶ%�-��[�6���m�l`��lH���-�lb[�6����m�l[`Ķ%�ؑ���`��6Ķ�m�la�Ķ-�m�l[`Sح�4Ķ�-�lb[e�-��%�-�l`[���[0-�lb[�Ķ%�-�l)��-��%�-�lb[��1-�LKb[����-�la��Ķ%�m�l`[ؖ�L�%0-�lK`[ؖ�ؖ��m���-�lb[ؖ��[Ķ6�Ķ�-�lKb[�!�:`�6�F� �b�lm�i���"6�ؠ�`�lPm���A�%�T�Tm�-�A�(��؈�b�l@m�`�lm���A�*6�F؂�`�lm��`�lPt�؈� ؀�`	��Q� 6��
[[`lDm�%�Q��F؊�0�"���
[[`�lE-��m�`�lm�-��
����b�l�m���� 6�؈�`#lAm�$`�� �"��F��b�lTm����6��`L@m��� 6��(� b��l i���(6���b�l@4�bLPm���Q�6�V؈�[b���[Z`�lb�[R�
���(�-��lAt��"�[b�[ [`�lDi���":`�[b�lm�lQm��0� �@�B؀�@� ��Vء([[b�lm��lm�����$�m�-��� -��� -�-�A��� [b�lm��lAm�lDm���F1 -�lTm�lAm�lAm�m�1�lb��-�#-�l`���m�ld`�ضŶ%�m�l[e�#�-�`� �%�-��[�6Ķ%�-�lb[ؖ���%�-�lKb[�����[�b[ؖ��%�-�l4��Ķ�-�lb[���F�-�lK`[ؖĶ%�-�l�bS����-�l`��Ķ�-�lK`[��-�0-�l1m�lb[ؖ��b[ؖ���-�l�����m�lKb[ؖ���%�-�l`��6����-�[�6Ķ%�-�lK`F��-�-�l`��6�0�%�m�lK`����%��Ķ�����m�lKbSm-�4�-�l`��Ƙ��`�����_d��&b�~_��yA,O%[3EKf%n]1N�Tݨ^��è[n���Z�70X�� m:ͥCt�V�N�O;�|N��j��V��k�B�M�N�&d����:���!�ڤ����0Kǚ5އ��FXN����md�p�*��ob�m���Ÿ㙓i�4ke�xj��6��.90�X;yiс6}���c0�+�]��j�m�)����i�r��8I�,�IH�zb"�Z3NG�\.�FM��fl	�T��	�:������V'SK$j�4����n����Sq�.Vc�y���6,��}hE�j�d,<O/�W�d�kJ��Bn�HRC#d��/u�;g)�.�7&���݋f��֌w�ҳ�]�s��q��|5<Ճ+E���))2=�6�EW[Okl�pL$L+�6Y�_Z�\gd�p�����e^ࡈٗ�Dd��i��4�ڧ���xXe�Kn�B)d�TIXZ�������V"��*��(�� �C�ƚ���V�-�ģ���tNʡRib��n�7��S��,��Q�7�Wokie�[F�b�SP�28
�J�
sb�dy���n�عeǓ���u�.t�мk%z�֨��
AR��3Y�GX*���h�w��	y#��ø��Sx�MZ�v��{P֗/)����73۩9�M$�56p%�V�sf�M�����n*�G(lw�]����#�)�Q�Nmm��8�E���J�Ad���"�`�3�T���'����X���,�;�w��U�.\��.2s%X�EE+�u���h���l�N&Z��1P��M��Vc�ܐܣ[��\��6��g�U[L�0қ,�=Z�Pݘ`o8��Ǘ�o+m<:�k��b���,[U�C�;L�wW�����홻����p8�_1٨���UYv�S$�,-up1q[��T+naL|��h݂��v|	����Y�Bo[���;������c�b��[t\͚�
�+�j��z	Q�ηyW6���פTY�y�u����W�b�#�8�c��P�T�H���K�D����.�[�T�ۻ�Ƃ䍡�WE����2�����.�����or���)iaMm���.��?D��	'rei��.�.;Fd�&Ud��%�V��n�D+R"��3�͕&^���xPbVY�z�;X�ۭw[�wPX\��ia{�C4!��ɧt%b�J�����N�]k�x�;LjKh�*�5�bhm��W��bR(�^�&���3I%<m-=��^�;��a;��Ӯ%m�6n^P��p�'2k�M���fcxH�]��Z�Y��L$�r�z�2�+rm+'THt/N��dT;!�^����ػ9,�a=����;x7vLЫe��Ynԣ���R��R��'M20V�T2�����Fź/=
�Vn��v��t�PG3
6lc�U.�0Ln�^�Y�F-�ػZ[D���k����7�{�>�	�Եnnm��]j8��Yw�gAv7wAm��ф���3w	��[��l�sN��ʦ����a7#��mb�A�t7���t�g��әbƼ7����׶fna�usSJ�[�+	rl�qI��ʃ0����
�U�Bv�QKV�������4�P끝�����'�4!���F���e�ڄ���/�pvs�'��V�x,�+��e�w�4�Zk���vϖ�ٛaҒ�4:̷�:�T��݄B�%�X�by�3Y��*�ӷ)�(Ɔ
�:#��U��7"ZS��q=F�!�r�K��n���U����9214^��Y7�"�L��Ά08�t(�#n��M[��<�e��2J�%k'F�EV�n�-9a8�Vޅ ˇI*�L8k�iкsU��͂b���0��g^�Hf��*��\�WpLՍ7�ZDlV�V3v�Љ��X�1	\Ӥ�0����ĺ�v#z!O���w���o,6/P���y[dS�j�ta��&@l�Md�M�KZ���V2��v�����PI�/d�MT�Vf��P��+37,c�&60��LTI�Gs6��*V��Z�͆f
ii�5oDQ+�c��频P�t"�k؎Y�<s�C��Ya�AƍN�Cq���S,U�d�p��r;
J%���3v�7����u������Pa��J�����"�ܤ���c�=��="����J�Z/5��5�A�P���M�����Y[x]	x��i�Z���6=رTAѪF�{�L�6n$�vQ��Ă����ń-F0�.ʣw��ʫ�6��5�]x�c�N��]��J����tmi�L�-�ٍ��.3T�_Vlj�Q�Y�U^�t^b�x��7h�[i�ծ;w�2�,
6��̈́
�q��(�e����4�
�H`܍��0a�����K�9�Třf�N�Դ.��k�4SNc��$=������6��m`r���]fbS3wo$�f��k��1���YP�Rʺ$۸�����^ӥZ��ɮE�R�7�
�,ִ�'*и�5�ݷ3&�J��.��A6�R�Y�J�J�:)��F���	��OAbe�&n�ڱ"��i*�M�"U%]�FYǶ�bˀ�s	�kw7Jț�U�He�U�Ӛ���\]���SN��i�J�{�<�\Z��Cm��+jmV����6)�Mdz���칯v�Ȧ�����������Hږ+�MLb:[�f�D�q�l�w� �șq� �*��%�
�5:�zQ�n쥺�p��n�ƭO4ۏ͋��*T�uҬ���Gv�KqCUj�V�h�_U%��t�8tX����(V��+6�ͭ �`�ڨ�p�
Ó5@I;�\�U^L��"�wk��L���yYU����/)�ۦ�n�sn[٦����&�Xy���d���R�m3a���L�(�藅{S.F�Ĭ+�����h,�Z���ld�j�,���u��E�{&1�X��7�j篺�쑊1<��gl�ʼ��K�Z����b��K��B7,9��h���4ƪ���a�eb�5�2&w
����1�&�ꤜw�QSa�eP�,�azS7�J͙�N�dV�۵�|@l0�o�e �p��V�,��x�����2kU�8mE�m���p*�̂ؿbZŉ�[���r�؛X�[��k�-Ƣx�[ʒj��l��Zwq⯬��SU����X�ad�kc:��UN;8c��t�b���\;$v�W	�N�Bxq��)%Ag��Qѣ��nڨ]d0% So��^��Z������z����-V>�X$RwCb(hV��-�
�X��]�ң�˧���]��:6�n�p���#��I�(S�t��.6�y���,=�kΪ�D����yKh�%�n�R��{,��aqJxJ�!��-Tܭ0��,�3^迮΃S4�ok�T�V���)�!�[�Ѓj���CM��^1�Tm�����I7֑y��B������6z]�����I���|B�y�g�x�4	%k����pz��m���L�t�nS�v=v����4��N���/�3u5�U*��oi`�%<7W@��;zf�=�2M�;$ySC,IQ^8CRo�E��ʕd�4�ʙ�-�33R��՝z����j���ηK����A�����P(��S^՚0�D�Rd�+K�t� B�ƞ꫶urdu*�V�S�1D�� UU�Kj9Zi�e�֧��Aj]��0���+P��b��\�3��<���x�4�_��0�z��cT� ����t��&z�Z�o(e�-�����^�k�Z{�N��[���w�shz]�Zrʱ�����M����ȫH�7X�t��>�g	��:u�UY�{R���6���^�l�L��,�q��l���T������c]�b�Jrf�(L�e��J'<���Je^\̎�uNb�FB���l�A��n�	F��-�N����#1[�8�f�C)UP[6�
Ť���z�ui1I��s
�����[��m�V_$��\��P�˱$���Վ�1KUJ�3ԎnK�t;ut�:9�,�1�*R˓�2a� ̊q�����YM�k�e�e���^L{�l��ܲ�XDm�l��UV5#��E��]mA����4�UF�b:�*�;����nA31�,�]�REݺ9t&a�X{Q�^8�!�Tu�gCl���c1�q���4-��7%�U�]�R	�!��2���-�v�+��[	�U[�bH1�N�bh�К�KP���[H�K	�p'4Ķ�X�/�e�RG�0D]:%A.a�lje챹��
2��T�W�Է Am�^p&Ӣ�Ĳ[F��-k����V��m�]���$,+��b�h��䡔jS;H��I��&��L�qH!ݻ�-��/\���J�W�=�6&eJn��ڐ�a��M-7I�ud�Zl��Q�LA��AkODƖD�*�d�G��#1c��q��Hy�HZg�.�UMfU�[)����jNc�#F���'a1UfҚ��(�ٺp$dz�u�q�`�2�XpaO�	�gs�m�!�Np�nJ��̵xU��n�9���㐲�D`���4��V��V�iRU�	#0�A�bb���v�:r��'4�l�b�fHD�y4�u�9{X���:�t��Q�y�
�L�ŉ3�n�\�-��.ևhjr$V��.�eǊ�)P�<CV�뫬��2*V)��F�(�;D�k���ڂ���]Yv���j�����ǖ���TJ,4��Cv�UUa�`����.����F���Y%�1G$�����ˬR�n6�ʞӻ�ݼr��l�n^MǸ$ӻ��Biܭ�ג�2B�N�V��/\C%R����p�.Ĩ�NZR��FLF�u���+�nd��و�T��"͢��,!��a�����˅jn����m�P�Ѫ�ܨkȾU�-	��F�V�nU2��yz�Ra;���0��G)!�z�U��e��e����f�po��>)-cR�ƫ!��ͤ]êl�xU���H'�
05��FKW��23F�V���y����©9��\�9��g2�&���v%�o����m5��8�M�7/q,�+3X�������8�d�*�A̹�e10ƦV�
���ӛ`���#Ea�n]�7�d�Դo&�q��"J��kh�u��X�n7S7	�����rسV��9G�T�n
Oc�2��U�̩��87*۩fF��� ���"�hԤ�2�I��SZz���"���nV�
L�PB�s��u����A���`�b���l�x�'r�˷�9�[j�vaE���UDn��I	���7pcR���L��u��V����ʽ��0��2s*]k6$z6�kt�.��� M)���G_��F�\�jdٖd�Z��c$�a4�teeK{H(2�G0fY��j�zJ�D�x�V�{���z�ӫ3&c(�����7*�R�׀�A��L�Bl����ݦot�n��h�+E���l���9�b�M[0<���@�,m�ʁfǛq�xn7��6�&�TWo��Ir�8�l*'-�!���b�t�d�-�3�pԼt��B,u�����X�-{j0�꫸.���ؐFպ�,L�c\U�[f(�Ǔ5`c$8�_�Yn�7bd��RQ,+���'�U�%�+�S1�`�6�^}(aq��-jM7�r��E�Te��r1��] I�n�i��6���l90֩t�Qɻ��D�V7��T�K<'%�*���+�u�Oզ,h��K��W=���ס�9xvvP��"�H؛�&cá6/��)��0����N�9�f&�U���63.�\��,�;+fn��m�L5�2�Z.���Zٸ��4�t2��|�7G�H��9Ω#w�}�V�"�Zt\����]��b�@�:/%��T��1E�д���-�5`TV����Iʄh� ��#eȶЫ�N�=R&%���[�P��6�SY�[.d~�m���p(��w���b:i�75��������L�V�HK!>�m9�7l��P��±Z/�3B���Ŭ�,"?Tq��N�%y4�F��P4���J�MmĮ��X�����=���.�(�fr�tis��x,iE���H	�D\"Ș�0H)Q��H�
���%JpI���!����{r"~!2�)j�-��B@bD���-+o[�
\����Ȓ��:��W�SB"��]N~���ƹ!�r�!�.�ޜ�:�7m�q��pĝ�L�nK`��v;�kD���B�H�Z�A��m� ��j�3HW.�ٯ̤�&��6	��W
YkqD�b�!��gj�G�
z�֩s`g#�#.Ќ;�:�@��VȒ!����j�W7ڭ�s�D��������ʭ-I!Ei��w�p<�"�@�9]��5- H��E���`��Z�v��b�:�x��0�u�L�U�]�Q���x�/W���V��m�̒ ��I2�B P�iLN��#�M�9/96�j�u�9}z����3�2Y��c�D"�w-u�E��
L��iXX�f����"B̴�c�-Z����(7|���4R��٘�u�ݸ��]��Q$bԆ��f!dV�(6��x�,Yo�֫"�.N9������G���vVSP�_��W'HY���u pEu�D4MȲ.�+X���5��N�+��;�3C�۰P�V�)����]B��X�s:����-�e(��ӈ�f`�p;حn=Y�r�;Hv��7�h�6��?;@�'J�c�5�m�7e]eK�Ő�h5�Y,k�$��M0��h�����.-��'"Ĝ]���U*h���VR@��T2Wm�~J;�G|���V�g�ȵ{���\E��{�r��ѥx�VEb��**��,�N&jֻ�m 뒬�x`.Ru��sM.�Px�)���0�ؤb�+�"I$C(M�rU��/�$!���p.Ř��TԋS�E��-�VscÈ�Ӂ�TH#H�mgGX��J��Ȼ�J���nj2��Mږ�Ej��Ȧ�1�VWM��	w�C�d�2N\��BgRi{G2c����[��f4�J��M�a��(f���Ҏ��0��%�L�3=K����h���}��c{?@����������Bb�g�����S�]֬�_d��zkՊM���T�ĥ��.�Ғ��*�z�9RPyMGvJ�±���
(�qn�jh��,=njRo
���b��+�k�p��n�<qĪ�:�;��Vɵ�g;U�N�n��U�
�4�uu������Z��9	�Sv�m�A`3�m�xs&�i�w�:V�z�~�=<��w����]k�|��e�*Q�['NWp��je
V1��4�x��ѷֻ�<���F2��yqM�(�Z�Y�<�c1�������;zj
UU�݋f[���4��x�.9Ь���R�U��anKQ����q(��K���Wa��4�����Q3������4O�S�f��:�l�\�0���wBof����Td��|ڳZ�OR:(;W��v�B;�j����.ה)έ�g'vN48�Ԃ䴺!U�_�`G
���Â՚4�H�r�cmb�@d��i,y����UX0],�=��e�e�j��xgJ2v�={�ٚ�N�����0�V�}5��[���Q�Y[�X"�/[�p��\���^Vn��V�O
<�t�]�m�jU�똣�+̮�w�[y,�蹾�o����m_{i!��6�0S7̓��'�:E�vv��7�1i��N'�鸋��M5{���z�>�gm�;�:d��v�4M�n���Q��u򡙱q#�u�R���+�,��̗��LK�$�.��O�Qz4�YdVzK[O+yeގ{�O'mu��W.�S��E۷x�c��O�}6�Y��՚xӡN�&�9ݻ)�o�+י���ے$�]pm6渁����o��z�*��Ӌ*Hk1nQ��C�,.��3�g�>Ǚ	����f].�4vcݔ,��::��N�.��[�*r��*�N*"���+o�<HV��,��񪈞��:ks��Ȩ����-R��V�Z���Y���۪�����>��s�F�v�vl��U�t�FJ�!��5��Rۚ,�s���:��Zr`k�D%:�gE�*�-��7@��7Z��e³zl���I�4m퉬�8㱊q-']/��h����9ل�+փi�ʕ�u�w\�wp��W��J4b6R��mA�I}b��b^�+��[MF~�8R[�8�I�9�Y�=�z�%�fU���d]F�t3
�ek�&������b*��r�����g-��G]��;[0�]�[ErrS�Iu���a��>U�;:��Ju�L�\z��x�m��U���3W��jn
�;6��Z,٬�V��{����D�N�6��Φ��&қ�&<I��# �x�ͥ�b�s��(f��w%Y���2CGD�Z+���r+�kA����.�Z�0�6�U3T��ŉ������nv�zT�玲I���G����[av]W�3o�E��q����Qmb8�9��WT�f���T�;6��-wR]3
I�f�;�A�vrLW�Ӏ�.�}�v�&m�9TԳj�ӕ�=i�u��L8�C��,ZC{�f�g6�j���Y�,���8��uu	R2��������0)/�:V����=�U���-LPt�xV7��r�e)m$Jgl�v�:ɉ⣋&�[�q���}�<z��E��*K�&`���#�����!G�ȱ�����MYm�m)�_*�38�r����*r2v.�-t����V���x���ȁ5�ݘh�l�f֣�������ʙؗv��k��zx�Z��ͅ��+L�R��8u���ޥ8F,�����ެ��/^Ÿ�q��0�VF�Yc��o|�bI�^ә��]��gyNZ���[�m�ר%�B�_��/�λP:�sM���j]5�<Ӳ�,�����XY�%�*�<z�g��r7��@4e��6�@������R��f�dt�
k�Oi;�IA���,Z��I�/�%=6�BFP�����Ý0i�.X�7�XұhJ�$��0⪴n�K6BT�RĻ��a���/t�j�n����[[���2v�Z���!��+۳�=���X+�oP`��\��s���p�͟+����|5��{{�OlJPW�J��(�ۅAw�-yD�5�r�Lk#�/��A�Z-T%b�ڡ��9���ɧw�mr3��Իo����4_EJJf�t������+��c �h��g��v;�����}��&�k	bZ�T�*;*���j=2����{��w����r��f:��!�F��y�3�x0t�	���zf��-Ĉl�2�7v�)�;���[i�o.:�Ԣ6�L�	�]N�-GyI�3Ea,���fYj��M��o��!�p[��Z=,qOs+��))~f<V4��l�Nq=��&�O>Y޿c����#�윪anF�2��\�O��	%�O�k�P�2�옫Z6Ʈ�#��Ͷl�s6��$ȻzΓ6�IWХFh�Ql(l0W���i��L�}n��S~qP˜Xw2K�QkV3k	S.�t=β0�VR�$��3n���0�-V�o[�.M���vb{���[����3�]��^H�!�Px9�]�3W�ϲJ��Ŵ��R�[gO>�z�5:�/ҨlV����L
�6b�뺾�v�nC�pБ�p��q��}��F�ιGI�#��>ڣu����1ʢ)b[�d�뺻��1�ʣz��l^�����$�����sb����Z?e��)}�2R(�w�F�1������9��W̎(���3e��+3
ż��w\��M㣿e��g�\s��Os�:��"���%��g.)��N����M,[���kכ�GZخ��O�O'%���.ĆIx�7��'uKC���/�!Xՙ,J�DIY[���Ak	��=:
i�Ә����O_=�t1�;�f"�Af�n���w㽳ڥ��֕��S7��`Tӛ�Iʪ�'2���-�ųT�'@����I\3{ꓵ�Q�1Hj9�t�2�.Gp�wNMc��0oY��q�7�\-�h�v^��z:M�0���eQ;��^S�y�W��3,V_dN���h���&��B�:��-ՃP�Lbˇ�8�a�QITn��N%z�ȍ3kf.l��Jz�e����,͈��լ����q��q�W}H��*���p<Ur]�!�$d�UO���{�2����:��g;�/ɁI����#�T�e�-����By�e�N��� ���V����ڮ��8U���z�;���7��^]���an>���d�r�;y{N�$��X�z�;���sK7J�Yt!�ᳱ=�rZ��f��Ҵ��)����Y��yn^�{w�,��0���7���bv{S7�]V����l���ۘ�`"B�AC.��f�\kRaZF���D4e�Um+�#[ײ�gE w+yXx2��[ke�#7n���j���æ�\�P�:��.[Ǥ��ME"�m����e�U�c��5e2ޖ��P��i���r�d~-��m�.ב5y�-z6cߥe�gtE�9-���b]5Grƺ;o�7���C[��T���7�m�˖Z̶�nN#��5�p��E!ovS�S}��*��Z�P��/���r!����r����C��1�T����1�w��gN'��5,�p�XÑ��5�k��ְ��.rW�	��z$�ng�=.�\�0��k���Y�Ѱy�[M�����Bu����M:n�J�f��'<��-g4�ˇ1��3b�皲�i�=|�Ԛ�V�ꮧ�D���J��K��^)QPv�nu�n�r�Bc��:(U��`��cUȢ㪩r��o�&�q��V�h�]�YV���bN<�U�������,�:#_Y����6��db���DV�.'���{�YV��*�ں��}v$�N4��w\&PI�;v�gS��)�Yzk��c.AK7�=�u#�UL����}�5n���Ml�&ə�0���qm�T�Ɋ�%|�v1U�5u$�Wq�f�[�\�.�Z_Vu8c��02�?$A=��d�N�)�	vł�d����{H�ק�7�m���{u��,s�$d���(�,r3��l9l$�C;{h)�<t�ޫ���x�M�bF��X�����ۇ]mϩ-�4��Yܮ���cz�d��)h�8�Cˎ�w�ww.5nx�R��P���J�U�ڂh]X�D�h��J���u�\��93�So���=60v��ߒ�o���2���S�U|����ov��u���H �-�%m^c��o/��ur��`�c�D;ӄ#w2|;���#��CX����1�MC�2�Nȷ.30_!hes/'c��aZ��n��S˼���3�]�4�e���f��T���6�n��̓��,4��)^��F�A��Ӈ�;�
nd�T�^]bsnt��8Z�j̖�6:����Hku�Ӛ�Bv�&��ƷJ9O��6�ML��/����ѦD�b��:�N���o/��ia��Y�s[���F����[.W�U|��ʦ�u�*�{�ա�A��\���$V_M�M��ʞ�Tub�V��d�m��+%�ڛL\b �	���X%��q�a�QiΓ��<�г�w�oT�`޴WP�`/�4H])i���V��w��gOU�s�
�|��`�+�E�|��aEn�ʅb%V0�nH����MvS�t��-GA͌�M�IV��xY�y�*=�����ʬI�X�]�*�f54h�tރ��ԻS
QH#����AbU�*�����]R���Ի���%�xz+y�$v]py���{�P�ңR'�8,���Ht&��Zj�I�0c�Fi@�ڳx�Cj���n.6;o�������,�t�{��/j8s;eEW�������yW:�]��Ѽ����x5�Z'u��i2���rY��Iq��N�23yI%F�r�u�}K��2�#cz5���ؒv���wg[��
�볅��3k(̺ʭ�h@i"�bb��!��L�Uh㪸~��iNT�)��D�g��ix��UA#K�/y֘Y}[6�+����82�]�J��Q;��� �ڵ*z^C�t}t������:9�aUxE)�6H\f���'&�<��Vk�|.��)��X�(�'�WN���˽�R��d^uf��Хjڱ�'rW��ݔ�H����Cu74���!y��L���X�m�Ki]i��U-5���FM�$��eAtF�ڙ)�麎�n�nj
�E[�!=Yr�b�c�ŵ�IS���[yL��83N�	��ʷr�9�K��e��O=�W`pE��m�{�u�!�{ӽ��|���W��Vː�nJkjQ:��\Z˕��˶���o+�C�0�)u��R���Nk��vEM�����Q`�]L��:�XB*V�N���]�셔r�%��7��ڴ�^���n�qd��w;/��z[�͝y.���uQ�5�8�+��u+���ܹ2:q9����M9�Ј�o\�=w*e7Zӭyl��,�X��[�̹�:dޚl�ʓ
��$0B���i�cWvҧr0�h�T��ҝ��ka3 ������Q��[Dm˥MdݷN�l��",�L��n%,'Z.���r��T���:�-X�|Dv�O��Vr3K��7ibG���rr!J�R�^]��u*�S���i��C�y��B:�g�Vv�!Z�]���5��`!\���ϳp�{W:J���5م%Y���|o��넍��=�[�m4��L>��#6y[U��gaw:�k�m�soyo{t�y��t�6�\Ӗ%Wڷ����W��7�R�o�b5%f��;���'E�D���.;�)l��$3���zT��;z�֪%4�<�9RI�gj�W5���}|9Nx��oxX��,Ƣ36��́h�����\�J��gS�;�vk%�Ď��,�����Y�Y'�.�=�B9T�3v���[p?t���,$m�9����.�\��V��4�D�U3$rv���L���ͤ��6GZ��1NJA/�W8*brM��WNՋ�2oF3�ή�qӗ>�]U��ܿ�ڃ!ӗ{��.Ugl���oNNI$�7���f�f�*��6Q)�H �!�y�g�ҀȈd@�Xʦ�P�
jZtڴQISEșO'���¨���d^�Ex$i���#�2�P�yU�l���,B5��ZM��-(��Y�	]Lܢ�	2L�H�#r�a4ZK�/0���I��*�[��ua��"c���_����b��j�.��o�7	�ݲw�I�zd�����"T)XiBQH���'%��Ն6�@�6�$��ށ��M܎$R!1�F�����(Yp��*�w2�k���$I��Bط�MF�G.���ܧ�����5$�J�C����d�TE*�WTX��!���BT&B�T��qt��:©Oі��99%Sn��b�<�&�a�p���2�	�����e	$it���"���K`��a��P1��$�1���`$��h	(a"HR�҄�QS�7�)����m����eWIw#7B���mF�AD3�A�C�g~˗��Q'�h����
�ف4ZK�/0���G d�\^�U��	2YDvV,�h �"�Je�S�]�)$�%HF��S�dĊA�b9��J5Tk�u^��C�Zw��J�E%�"e9���A�q����LV�b��6Lад�H�".�0����eU�X]P2���d�k����?����b"(��;�	�?G��?��?p��/�������?��O��g�W�r���J���ۨ�X��YOr�#FL����%�ax%K��Τ��W��t�g,Ǉ��a�)�S�����@R�*��Z�ܬD���\n��F�<�u�k�N�]�[Y�ә�2���E�R�C2���smd��y.7q^^^���׏�Z�nۮ��r>��*3�[�:�d�S�S~�W,?`å�S[Ͱ�O�۷K��[�y�u(5��/c�7f�!�/�UCs�e��n���C�B�WtC�p0p�	_-�R�*c[�Mّ���Y젷,�Ǉ�Ϛ̱�4��g\�+)�0������[��t�/:	�w��/ZL�wV�OY�����r�N�ΰ�@7�꙳i�W���0<r�Cdm�4p�����#�x�c��X<["�7���ٽ�7h*�nҋ&nl/Z����Y	'Wm��y��]���G)��S�*�^.*w��&��\���T�4k����@M��na����t����Td���(����ܡ�M*�ҹ���E|6��.ҁU���V�����ȩ�P�3IK{jv3g�ݩ۱Y��5�w�Ϋ"s+:@�ou�֣��X'��*v�.�
��Jc9���*K&�l�Ra�{�)<W|r��\N$�B̾W���SO�:v�8ێ8㏎8�N8��q�n8�q�qǎ8�8�<q�8�8��8��q�q�q�q��v�۶�����;q�8�8�<pq�q�q�q�q��q��q�8�8�냎8�8�88�8�8ノ8�8�c�8�<����Q���/��ˉ]gZ/��с�nB]�3l����D��F��L�l�X狡��xiR[/����8�)��fR��u��˩|�u�0-�ׇ;I�وۙ{�WR��ޢ��+w��%H ��K�8�fU	b��
A�2��Ν�;�F,�pD�{�`��L]���'F*��J�*nK&���+���K��*�́�7�� ���δe�&����F7uy�uj��VI�t���<N���=��k���2̎aR�,'h��YlN�cj���r�g������(�Ɯ~|�B�m����Ɍ�֯�PU�����%�����	�|Xx�����U۫��l�*�;��L�&2d7�lv-[uBY9+1�&��� ��ڢ�����q��ino��W27y(F[�w$�Fv�;O��ag%�k�Γzq-��4�����I-[�P�8�ڄ���z��v����iZ��A�%�UQ&b{��r�[6Ӣ/���ɪ��Lp�}qL�	Nh��^RM��c��������gU����9�B�J����Ჲ���5ͪ��h����Ӱ�^UI9u�<��u�fr��v��oc�q�}q�8�8��8�n8㎜q�q��i�q�v�q�q�q��8�8���8�8�۷nݻmێ8��8�q�}q�q�q��8�8�8��8�8��8�n8㎜q�q��qӎ8�>��q�q�88�7�߷=�f�_�k̩f�.Z��3�����D9GE��Ӧ,��#��jX(�8)n��h+�r��;ʡǦ��Z��֎%e��=kf��hH=�;�O^�l�75�x��n�{�b�����j"�m�T�dT��9��-���.�2�3+z�%1�������c1Ҕ��8���U�T� �Ci�R!ۡ�=����݅�E܇F	����6�9X�^3�*�a_�]2z�+6�t�ټ�ذ�o��*7��h��d��=�W^T�P�X�Q�He���b�����("Ω�[f@m��=/{$Hu�r���H�U@�x'E�4[�<�W��9\)�R2�A�w�����rSJ�tm�oL�����mR��逆f�O/_�	7���^U7�v�.k˖���v|�q�muSQS�8җ��F�{u_F�־���$��ɣ�=eff%Л�=���:�8͍�V����Q��9s��&];�Iؖ}�pf�L.�ĩ�zƋ,�ntSڅ9�q�'��e����G��s��j����8A�ڽ2����.�FR�u�3��r�8�6�Jݽ�Q�2��gU"���Gʐ�t-�L��k�{�r��}��N�_�q�q�8�q�q�n8ӎ8�>8�6�8�n8�>8�8�8��q�q�q��q�N8�ݻv�۷v�8�8㏮8�q�q�q��i�q�v��8�>�㎜q�q��q�q�|q�m�q��q�|q�s��tvc���r$8렶,Г��h�:�(.��+����]ë��h�����ކ�p�;/U��'�38㾶�h^���@��L�Ӝu����/*�}��ޭ �9iI\���v_^=vkx̦v��m��̻Ǖ}�V�����S.��7�{]}\��3]�L�e�3��/r^��$�7Cx�"f]u��:�P����^�r�ܖ�t�[37,J�}�����S�������I�'��9p���75L��k�!->UC)<s!�OE��Y3+%ƻ���%�y(����TQ�ѥ6��g6<��S:]3�UO_`�RP���s�n]s��o��C��ر5�
UۖW-�%#�EY[��S��kJ{�n$�avҧv[7Yk{��}>��etM�ڰ{�e$zұU3�+4L�&��ڷ*�ՆqXm�Bpj�Й�2�ia��N���X���_=�K��n����EuVu۷�aM5m��PD�Z�֌'i�p��FQ<��z�cko8��D-�/%V,X9,�CZ͝{)��X��g�YM��Ʋ?��]塓i�:�#�%�4�M�F�_����j��5�=̈�/Բ�ed� �����q��=��3�6[�	���r�f
zN�`��$td��$�So{"���M�m4�3�բ��n�V9{�z��M����뷍8�8��q�q�q��q�qێ4�8�>�㎜q�m�q��q�N8�8��8��qǏ�ݻv��q��q�qǎ1�q�}q�8�8ێ8㏎8�q�q�c�8�8�i�q�qێ4�8�>�㎜q�m��+|-�K�U�c�:�I�["L�rf�P�����U�eT+|���	��� F�űu!��r��XL�ڂuW��3	�R��ot�Q>��h������8\��&����9�D9,�٪7��0g���<�Jr�
�������yi�s�����N��ز�Uy HV��m�����Z���_0m����]-F�`�4P����&S�lv���of�Q�0MiŜ��*Ӱ�#��J����rz*�[���]�� Iz���Ȟ�u[{��ylD�S�g���A��9�w[�0�ʢ��>P���}B�S����z;t�8�R�+K)bFӭO�V��K�*ϭ������#r�D��\VV�\z+#hw�cS�Z%���kvJE ��a�����B)�x'�и����O����ikrZ�^��|-�8ƞ�v��z�c5�qD�7\�T4�/m�2~(*2�F��ȵ�����lռ�h��C�:�=xܙ3jDj��$y��k?ђ>�n�����ʓ�!(bB׭rX�'�$��})�4��'jp"3�����M�c��|�l������D�-cZa�E�*��-�!�1]���5�e��5�E�2���|wv�|U̪��t�n`�F��=݀��a�V�\!�;cB��;��XZEC��:�CU�p@Փ�1*8|�lJ�ra�.|9�l���哫X���!��}S^8������'J=��"���]��rª�(�[�q�Ǥ��H� ���:L��^�������5�架j��ܽ��ΌoC�a	��dLH��@�Q�+�b^W+zZ>˳::���G�~@3T0�z�a��lI�X�Y�&[E�Tv4�H���Ss	�;����.�<fv�]>/�%;�Kl�y7�:��<\�л��%o��g5]��հ�|�-�����#>m�AA����x�����]]V���k�nsҵ�䶚�[B+�4�u�6`�n�_����G�:5�:�UD�mWb	���Zܧ�HC���\�;+*�����tzZ�sHMp�Usz/i})J�����,Ҡvzz��;���]��ML�]6����#c�m��Җ�^�\Lr�� ;r�M-��'k��p��y�a5'v_�}V�1y�7ZPq��c�'���P��U�z!�Bv�8��5�i��Ea�stXC{�:�NJ��uwc�9<��gQ�g���ݵ��x�RK�:ٙ��|�f#������"l+�HU��4����l�nCv9&P��rAݫ$g
3gj2�a21�<��A���Xu�Bv�ԭ�ͭ9����ܥ�(��8Qyi�K�"��R���7;��d`��W/%�{C��J���,��-;Te 6R���F��"�fV�sc��$���`��%��Mp�����Ä�:��6�k������W��+��K����5Z���;}�q�XV6�|SZ�\H�.���yHK��ޭ��1��9�wI�y2U�ב��\��we�ݫ�Ӵ�L�sz�H*9uB
��o�zhoIrU���΍�u���v_��ka���

��R��.Ⱥ��i�x ��Tq�E��v�7��r�qeC�����(�%;���uF���=ОmMD�K�^�t��Sڞ%ml���,��V�oW-=��%�8Ѝ���g$�ӳw�p=�9���]Cap#΢õ)r��s'>�$T��
�1ͺ��K�&�t�8K�i���շۙ!�s���Z�j�_n�il�!�B�e��N�K�,���6맨d�-�4!w�S%X�hk�­W*(�D��U�����S��:�$�Қ�doN׵��	��IH��'e&�RI���
�#m]'9�n����1����w�^ ��8��ZN�Y��c8,���S����2  �j�U�����%T+�u힂=f]�aX]�L[(�����	�,�C�+W���Z\���G}%�,��٤-J��*nX@�UT"C��z������0!F�d5��Y�e��B/�@�Y���U'>��x�g��s\"u�[�݊�ͱ�<��:)e����F���S"���;j��9)��;h�T=w=0t{�}Z��V)r��:4%Ws��ԕE�&eiJS���X\�'O�V+}J�Z�<�QA���Pd���Kvo/�^�M8*R/՘�i�N�7��Q2cV/GT�����9���]w4#l8%>���ۛ[zbWP�����M���1�n^�=qu�7#�.�җ��$s�
���]��ʃ��}ɶ�'O���휚i3F�r�j�U���:�F2h��=;����Mf����/i���l��c�o�M&Q��*��}*Xx��(�{+5�#+(�Uc����tpi�Ӑ�'} �QM�8$��!˹����^���5�O��ɀŇtֱ]I��� 7h�Cy;��s��p糰jݲA4Qǜ��A�'B[{�R�wm�(�Hv�����eSyαC��y���in'M���ֶ��M!���Ҹr�˪rRM�s�ToF�n9q����<�		ǥ=�q#�ݗ�v'nK�t̀�ž�9�9x���=��w]�=,^�#5�1s�XԮG�a��/'<7���K�9���s3��S���o���3��n�eb��Eu�!�Iv|��V�[�n�o�]96^-y�=԰Jh]j�%�R�W�q�rvt�;4���%�T��Q�\y� ���iR��Ce/���r����x72#��D����ب��ҞC> S��ww&��-m[��#!�L��N����<x������w��@�SvX�(�}�;*C�RNl!h�b��v��72�H`̣��V9�Y����$�����ӧb[�kkk�q�E��M�G�%�"��| �R�y�,ւR��R�q����8�̕,�S,�;'��N4(�/����$I�����b�����<!���Wl���U��vЅ�][]Т-N���սW��P���X�� �HYR�\�[��K�zh[̹�j�`,�x��H^�`J��[J��CӕlƎ..�Z�梬�5�4Dd�A*���'Y��iR�T����>��!��)�nv�F0Sz
5�R	�QǕ_��mi�vS�r���cAY�/yl��2E�yB�u'ʇ9�����W�nvӻֹ?����[�:����%���f�\[�h��a��tT7�U���s
��4�Z�f�R�vc�ԄDS��$Ef$�Sj�W�����Ջ�e_+�{nR��XY�1�ξ�l�]�-%v�uKLcl��D�z����YݳVޮǶ��U),Z}u�N��`Ȩ�`�5v!Ym�<�c��+u-\���q�n�cVMg2�kˑ�Ņqg�Z��AYU��ڡ;�����3+V��R#]&�n�6⼩���4ּ�u�́��'Zi\�T���ޥ�n\�q��N�~4.��"%F��;�P{�b��j�^�1��R���Y�����+dN��<�ST8aC n�m�5��T���:��|��%�m��\�n��Ժtw����!Ҝ�V�D���}�n��)^,U����}��{}[���ٺl�JF�庝���a��*a�!ݍ��UoX�� �pn�n����BѶ�^��բ�m-�G>���*�WE!zY��6z�4�G���˝0i�a���;�e�rE�+���ػu�v�Y��9w}�+��h)4�;K��>|%����dm�Vx��ߟI�%]Ku�R�;Hծ�6^r�z�]���*��$���8]g0�XY�.�R�������V�haq�޶-�E1�hj�ґյZ/�#�r�V`E���[�uk���zVꡭ��P�*n�FU2S��އ2�$+�p�k��B�Q;�J�E���Myj��@��Źf�w�3X~��}����=��������:ַ���U U�L��������������������V���@��=�-�� �!� B"�r%=�
W��Ed�5�LQ/)	(�ʑ@���4��Hj���xO���9���W�;�Y}ԓ�f�r�l�7�����62N�o_�tF5��k�D���BV�f�k�F-�S��������ʴ���t�{e: ���V.t���\h��u��}x�e��#)�Es<w�-&������*vQ��ڙ���ty�U<�[%־C�f�eǝ�Wq�ʪ<��]�5�m�7��uG�i� ��r�R���N�X僪f�X!�l������le�{R�᧡�ޫ}n�SmK��ñ㡄��
o1+L
�`����p�uRT�ʕc�h�:%��+�.>��̟l�ٛ
ү���/�6�}}εKJ�*�-9�˺���9�:Q睛̮F�X��}/����!3&'nf;UM���Z���5H��<���bK�,Ч\d�(����t;;��a��YE+�4P,	Y�2j�득5���n�Ge-3���d��Z)m�q�F�q�˸�	��d��+u1t�ncAc 9�uT����^�ҡ��31,N�]��֒2b%#d^�)7S`6N*�����`Ü(r�)dA`�\���(��s�`�����Ш�d[rv�H���Y[sW
�%�8���-'#��4{,���#�8*�=�QD�"�Ex�V�H,آL@S�J�1����E	��hHۈ����CD��NeDQ�"Op(�BE��b��j$�`��!	�2�B�D���ND��X��fŤ����jD�D���wv�n�r�Ӽ���et;�s�����˛�E��%��3��u�]��o)Z��A��6���nݻv�ێ1�ƱQ�X�IE{�㨴 PTo.'�4k⯏A����q�nݻv�۷Ȧ�
��r�4�69o���*j6�$IDdcN6�;v�۷nݸ��4A����{�cd��]�
/�˕�_�9u�\�Q�����.�wt�n�;�I�tn�7��߻�]�v�۷n�z=�Hǲ��G���s����V�:��wV���wQUw]���=u�.)+�U�ݹ��W��4b�DQr�h��u��R��tڹ�rܤ5��s����D��iwv����t�Ļ��Q6��w��7d�Gv�]ʝ�z/7.]k��뤩��>|��]�ޮ�s�n��,n��u����z^Y�ܲ�]�uit��c�������{���u�߷���]<�r���9�s\�w��\���.����ޟK\�����wϚ�[�����b�
��,�ݮi��ܷ�s^|�ܯ7��<���wo6��mr�����j3S!��j-;��_O)�h�Q�h����0p�_��0y[��5�r�7#E��.r*�r�^sb��j�|�\��}}|�:��
"�:�?[{��H�]�'��m�Pq�œ��d<��ฯUG�#2H�VP�(��tX7l��J!���`��`�UÅ���@�K���/���}�t�H�
(l�c��;�&M�$���ӗ����6��?Ge��7�a��{�6��������� �b�z{=s/��S�S��<�崥^�B9��E����N��=�,(4q��o�e�	���=dU7L��������\l����L�U����Ò�{��k�'�=��X:��mu�C�\�h4'Xi�������8l�a�I.{���ɾ�)�{��yG���M���� ��ɉ�͡�ni��O^o�l�5YUo��Ϸڞ�I�y�y�b.��z(y=�k�c�X�_��n�T�bs����7����uWޕ�2��85k��fߐ�ʲ�k���B'���|m&�������3���1�ңŊ�tG�����%���.����(>6"�n?}�_[Ŕ׻C����̋n�WS��F��g��skm��n�dhʆwX/r�*�'����x��6Ȍ��[��%�[~�{��ꥶz�R����b���δ��Wa�<�&^ݍ���7�Y��fÑF��WR�ƴ�>�����qe�]��	V �ϭtDy���J^��]�y���W������O�m݃	�xl�<��'i�FY�����	Í#*m�w�oa���,������R? ���<�W;�x�;�:���q��xɰg�:.>�����O�{q�I��FM;��S�+�ݪ�]��L#�#$���#���U�}]�IF��򗗼�l�t�Mp�}�CzK�7|�_{���g��B�g��9��Y�I�	��S���� 3��Ia����OJ����R�JGS�Mv�~��!\H���;O�Kq�ٱ�z(p��4��ʹ�cL�9��z���n��%v^��LdK�M�2�x;\�ٞ��Ol��r�y�T&`6U����:n�n��q h�=��=���7l�_�+rR^=��6������ai:GL������8ŭ8k}u%}�&�㺫�����eǼd�ytj�1�A�t��.�|�R��?Y�i��&r�.QN�厃3͹'�WߨW=#��Ri�d�ӭ�a4&�_� �6�NZ�%��Ow^�>�^���p��QXw�0��W|���s|�z����2�,��W�Y�;���2M�L3�4�#�+ݲ�5��u�������އ=���}^�Z�=��cL���#-��� hf��zD@d}������%j��Z/�۝�l=s�9�����ھ��a_�}�'���~w�/1#�:.�(��8k����
�[�Tk�Fd(��B�H���ǝw��Z_�y�#ׄ{���pG糼җ�ڏs�*v}#��h�WV�:wk86l�=)��
0�S�a�Ӟ9�g=��r��=����"0Vew��>�l�|�;�݊ߺKw�s;��{�}�>�2I�R���{ދ/�̼�����"���ӧ{k������V�eg����"�w+Y�ځ�^���(1ɏz�M�}�*��u��h�`���J�j�M�ɞ�U~]��.è���1�B	��HD��ZG+�}{,���&<�)Xu*��Vٷ�E�}�'K����W[�S���Z�L��r� �È^�]�۝�r�aj`� V2��PY��qMU\�}T~ Ks"z�=�F=�����V��9s��:�a��xb��R��5�/Ϗ��z��A�����1�OG��D�O��{��W��hP�V^`�6���f*Á&᯷u���x�2j��*\��uwZ��ud����v3��
�Ǵ�־�x�$����y�W�=���.I=�ei�� f ��8o�[�tG��<�:ۼ�2��#o~�}�����==!��|�t�T���x��j�sޥA%:;�dxm�����3ŋ�{}S
�겙�+�t/�e�/j��O��߽�ވ�v($@F�P��f���<|"�z�����΅��P�7g�3�'�}��QyW�P���AL�k�揮Vl����.��^�5�9�a�p��m}�מ�=�_ڻ9u�=�v�����ro�"������ud��������6�e����m�Uβ�F&�CZ
�O��1�N�U}z�c�3�wHU�-PW��n�Ze�u\��-��~P�{�[[5$I>����R$�@���uV�U/I= ����䂬=Xkr�
6�ݫB�a-g�#DZ���L*��D&�3}�>v��������q_+��AR�!9= �J{��Uu��W�&l��gON��r�F����~|թ2���/uWӔ�ѻ���y�ڷ��	^�Eg��λ^�E}��=�Q6^'=�����-F܈�˾'OTٞ؃�����:X�l�/�'�W�i��x_�p�|��S�)��ypT�}&�tD~�������yC�C5cDC�'/ނ����۝��?mx�3;��������ru`��f欯1)�`�y'�٠���{��O$�&��}���}�?Dǧ"�.��x͎�[�nO_PsP��Pk���]����
n-�l��&�ęw�gy&3�H�q�{�������ٵ`�'�g�Ͻ��#e���7K	�{�uwW� �: *���;�n;>���ٱ6��Ol�t����s8�\�>����lV_L����ӡY���J󘓇�P����8� (!�����-�"a�xf���f}(>��㷎�Ks���L��6���������p��x_,f��j	׾����1���L]e��Ҝ%p�-�JV��u�{�voq�i�e���i���y̕C�wC1�QU������]J2���1�L��%;U��0���[���ƽ�|p7�zI�v!����ML������O*�>�]DO]��Z#W��s=B[}�7��x�㪍Ka��9����=�}�s�2�`>fϳI��$ԑ7oy�7{�k��e��� xo��R�6F��@��&y�.۽*\�̐�/o͖��Xȧ�W�,W��vzP�A�����i��vͷ����/
�~�H�������p����o�W7Z���@}-���^^��0f��4yͯh��O�Fw����ī՛o����讇�s�a�)z�Ӟ�G��,9����7!�P�J���0���&�>�흜ƒnX���{���W�	���de�$�5��,�BX�o;6'��W� �����xޒ=�`C�T3�7;1�F��w<Km���Զɖ�����c>��q]_�`Z�M+i�)�^o�3�f[3���D���Π����(�b�2 ��s��Sj��q�\%�*����o��oX��[�N�W|omH�.`�Y5��-� 9(1����������~���=�/v����x����ݟ'�������A�la�q2h�?�穀�Lc�m������gN�#'����jx_y�a�?��k�g�ƛ*�ۧ;��������Kf�Y�P����/�`�{t;�`�}>YX׶�ALG�n:�����J��p�u�3�y�C/LN�6_c�5������V�cz�'��
?_��F�f��(�t�j�gٯڻ=�+[�w�Uӧ;t�޷p�QQ�܈��o�a=���ϝ���u|oޤ�r���Hl��ofݵ|�����m��Z�"�@���bzZ�P�5�:�c�gޘis��x+��\y-t�?,��|�c���LR]x�p��x�=���-�w˽碣�*jq02M��h�U��|L�E�vK�Gwg\ �f�x¼����<<	�زoh��t4*�v]z��l;��C��R�΃
��ܚ�
t�g�]N����X�R��Ǵ����v������r2�؅��,�:�t�q�> #.
N!u�GX����=�z�u�����3 �8c�f���+ǻ<љ�%g��G�|E����}7���w�5��	!����[��*��>I#��.��};�]�h�U}��oܭU;���kn�A�rD�3���h|�A�I8��}6��B"���y}T۴��
��w0�j��r�e��F߳<<�����������G��X��}g-��u����"��0���<k�q3�=�6�<dE�i�7����s�޾~az��_X�$س����&��/�c���2��ۢ����Ln׆k����Ǳ1�_+��s��;�L��=T��ו��������[2�l�Zڡ(߼� o�4q:+����o��d�����������;]��e0�_�|�}���e�=��&&9>�`g{n�wUC��\t�����f�[R�&h��!��#�JAv�Խc�{Ьr��$�ь9�-��i�{U������
����os���Dx� :��ܵk��ovY��ua�u\��2�/�U���M�D�Q��kw�UK���ݖ����U'�C~l�Y��#�۹�Umr���I=�����ͧ@e��=�����mp����6P�vzR�����������q��란g�����<��}S���o�fG*��5����b~A{��gPo��ݎ?s�ޓtc>z��?�fm���Y:�My������_�~�rn�v��^��C��7����B!{<�ǰC@�i����EG����=�3k�pxj�^��ކ�y���Ѡ}��B����:��D_���d��k+*u;��rމ����{��;��H��(N�y~�\7L���D�,o]��gnQf�Ʋ�����H�'Iql0�rdlS��l���R;�!k����#�ؿ%]��R�a��ɧٗ�/��>k�ɮI:�r��ӗ9r�黌�}ܯ��
�p6A�M���Olɠgq��3\1���ޕ�����MN��J�*����]X6ߪ�#�Y��4�t{hɒ;�k�E.b�7�U���V��;,��$��D=}�� ����Wy���ݹ�-�Y��d]X�7� z�l���}N"��)ҡӆ+�n;���V
?|�ݝ6u�Tw��ʷ�'�>��<�^r{�Mq�\g޾��o��l�����xb�<6��t	I �,�Y�A�{�׽��\'�3��1����vJ���
Xɽ�+b�����$�nz���NsX8�Q�,����rHsfq��잓�ϵ��h�'��L��;�g�yL��ȗC���`�)�R�_�]���{/�3}�y�^�=�E��hs}7��<�\�~���Zi*.�B~U��xP�/�,�.<ndoއ���x=ϕԾl�7_[���D�UJW�����~�c�2]� �%Jb~�V��I����6�����yj����3��|�.���׿V�1�����H�����o���އ�y��S(R���k�p���]��i#�/�f����2��P��K�d��Q͚o����+ڕ��:=;��)���#�~ �3��&��'��wj����ɉ�\'Y����c} �6#1c�;��X�<��.�Y��T�!DpKy�iPPWYm2whR"@��=J����s��޾�';;��E�g��v�$���j
{
軚r������C%]�F���eD�l7��	����(t�[�;W\U���這�!.��8.�/f�(S���״�e�θ+4M!���Gr�o0]�Ӂg����bS\�<�@�b���+v�~������l�!s�L"�MN�+c�;v�=�t�Z�5ՠ��EK���t�v�K�!'�":Y�w���#�Mk1�F�t�wy�z�P��q[��f���ō����cP�d���9G8GF�j7�mQu#P�.&u��߱�����.�f��\��7�ӕ[��u���UYn9vh��{0�[��|�AC��Ƕ_^ޚ�Z�M[SvӸļ�2���S���dM�Q��[���5����n��cT𦮻(���0���94�[��:��j����,$W>�e��wv�4��=�C�(��o5��:4"�k
bkcz�w����u9:Nˆ��i��5��˾=�@ܚ�fk��÷Rg�ٗɒq�1���x@ZBٿl��b�zs���j�q|�n�zblZy��4�H)�xB���t]P�;qW-m7O��f&����g�q����B�D/��*T�sso��hx�2��T�bS)�.h撫���|�Ig�z��u+�v%64Av�뭶��p?���j�Y�z��/��(n�;�ܾ����T�;W6�#nY�[F��o�$����Av0T��#�y�]#>4M&����R���wkg8�mb#�����(�5�n����ȋ��T�R8i]Mj�51h��ڑ��we�/�5[��]�պ�1��r�Ū��1�/#��^�d2��LZ*if`u{[�Sg0��hU5�P�����D/k7i��� ;�:KV\O���۫q��jض�����#��zj"�|��t-�ꊛ��f\ۏt5dt�V��F�[�SH��puL]_K�g�Z[��e�,�X*�f4d��p�������,V���Vͣ�"Z�����ʲ�L籭�������i*���Ӯ��\Gxn���-���G��GY'v��k��L�؃�Z�q�䤋��sΓ��x-e��P�H,�ru���
��/�F���ݷ��	R�s4N�ɮ9R�c��y��S��§e���Ҿ�;	(8�zh���*����wyOW��ɝ)Q��t�P��Y��q��5�+���7�஦N_$��3y�g1[�������y��8�gŚ��m��.H�^��G1%�=\��c���bUAJ^��khَ���|�����ߩ� �ѵ����qA��e���y��,`�wlk�����[���<v�۷n޽d`�	"�JF�^�\�_)r+�4Fō|]��5���|�\�s�5J��J�M@*$t�o^�z��Ǐ�v���dd	!BE�ȕT�K��&Nk�����,;��w]��y<��� �7�6�=x��Ǐ<z�sܦ@���׺��\�Q��nX��}<�ҖJI1��1-)�{�B��cO_��v��Ǐo���7��ر��(�5�%�ncG.��]���>�6O*-t��_r�k�:o�\�����v�h�EOt]�s�ݢ�;S�������E�lX���΄Ȫ4Tmw���lT����`�B�4��lV��X6��n-W9��&�h��P��M�ʮj
�M���-{�h�sQ+�;�Z�gNM�1�r�����j털pۮ�:c�j�jEx�b�)[�63g/����i	n���O|@���c��}�榻��&�_W_;
Ϝ��7[���'�qh�ǡض
q��|t��ʺ���?�;r��[V�VF���ᡄ2�Q��t��1-X��:2<⮶�&�l���-桦y�^8\1���+�a�~rM�����*?���D�-(G�D��\����
h��
�C*	N0LӍ۷0#�|���/�{�9�ؤ�����ߴ//��".�=�F��h\D����Gl�
T����Ig;��+��#�x����?v���}�1��xǶf�Ʌ͈�>�B�
�1a.7�&Wa��Fn��[7΀x���)�1,R�B��=���!�ƴ�k�	
 �4���̴�D�uj���J( %����bEFc���"�:"K�O�w�ړHµ}�ʔ�>��~���_��$E����l#��q�|�7����2�����ҥ'b鹼W��R���71o)悴���O�b|<$��	�9�x���u�>�8k�~S~h�?D�g���9�Į\�����-��T�������x3��RP��;�W�B@�~�k=�P��>�o~�r�S>�|3�\?T�m�-��42�^V;���m���'��������u9�����Ŭ8�5
-��A3��ߪ^]�-��hc��	F��"^�26=����&ᣯ�ɷ�Ȟ���q��S����ސ{Um��tG��{�g����y���G�U�>�i��oAO@�%����~���#�B�~���͇��PυS��*�Kd;�4�-����1��\]���^�>�S>��كp`-�����u6���4j�$l$M�2�|`�Cr�V�Bok��X�ǧ�j����Yy���{9�P�$~z���tZb!�69� �3����%�K���6de�I�(�`s�gfio��	/��ע�8�SS�#*�vj	�e%{��[;yHzgm���~���$v�kὟ�%����	�`���u�v�i��=����*���	����B�s��ht��進��*��k6I|�;z��ʦK2�b���@C!�b3ߖ/��r�����N��8>σV�ܿ��2*)�bYٷ��2fQd ��~��n���v&�O@ey [.qM����!�mL0��������#�ڥ�%=+1���G���l��׶�a�9>7k���L#�X�]Z�@�7����*���fpP.��2��yn�L˂�=��	��r�'�aľ>'�+�{��{=IW�+U\�_�����p7E3�/e��wֻ�����Iay�Zp��r�����K�)����7��}1��\5!o�eVԒ,���Z�/��GJ�^Մ.ר�Hz���Ȭ�H�#=�<����p��(&ލ3���9=ًR�vW	���k�p�6�Y�+G�3�a�����Ҟo��y����֪�Z���ԕUVS�1�0(�����3ރw%�W~����P/0���5�I󳁌8K��<�	����.��⌄�
qMXx��[����^O�t[BQ|o@���@�)Ĉ��=*3\�OwIǛ�����); ��>�7�{ݸ���1�[�\%~�ל&� ȱzX�r���u�o7=�vV+z���F�o[�Gt��r��@x
�nu巜�<ҷ�F���W=$�J��!d��A_r�Ǐ�ٽU�[�ힹP�����usxUZ��G.Qp,�.U�>O^��2;%�����7"�/�Y���)c,��$� 1��]K�p2�; �G��E��<Ɵ֮5�kmo{=�N���bLAn�}�rW��Ex@�M{=g�E=��y}l�k��ׅ�s'W�����K�b��J7:�8�2��W��(�`1�P���x�?
|`a���D�r�w�o'����c�Տ|`NY��������ϧ�p�(�� � �~~Ϙ�`��A��Lh��9k�'��m Z�V�,�eO�#y}���O�=��ˡ����â/������<�Ǘ��s~���Ml6*-���㪄5�� R�!�R����m^�Tз�d�5�t����0��%\�R7U{���'Ǝ^ާ2�����.T�fpY�˪�9&\�z�G��c�"ļڦ�ϨZ�t�>��7�7�l�ʷ5��A��Ȁ|����/�;��+���||||||G�g������ c �TkD�ς.��x�� ��e�-��:��!���5eS��Df��tW��R�)zOM|��=���)嫲9:Wo�4<�q��d�P���;�����2�  �G�*�/a1�L�/�T�3����vF�6n|�b��Q�cjq�b�p:}U������R�sW�����[�qm��;.��+���%5ޙ�L�)�ܸ�%�05��䐇�w�?OT��N (�P�@OqD��'�����G���O�h� cc�f�1d��=�Z�X�r�i������rqL�2��´��y����mJ@ZN,�@��20�ȷ�0"�k�5��&�:�v�q=�@�xi�� a�y�3 ���?�ȹ�
eI*M�A�/�W��a8����!��3�r����M�B<���^���/�����酄jQpx�Uk\�z1���1>{��nx�ܕ���Y#���t�x���Bm���f�|$�Jwf �r���8�]&���I���f�-A�|.SR(J���R����v��(@���lLp����Z�2Q�w�W�a�>����u�Qj�*�%��㱭�%#$��l&a/?����N�����)Ï�����\Ö�ԥB ӽ#���˲w��Ǔl{	�(R���wY0�\��j:NM�t9k�}چج�����,�a���>�/p����9�&����|t�1���K�y��E����C	���psഁ<Y��_���G}BA���4�[�X�Gԓ�2���K%�f��u��:����l�S�+�i���n�#��(�1� ~�����hrԮ��9ݱ�.�y��~[�I㮽�v�xb��c����s�V=φK?h�Q�«��t\����8��mvV*4H7�yO|�U;~DUv��`1/�Q�!��ܽ������
7���.>�Y�9XhU]��yY_�?��l\r4�G� |CD3�|�@;��߻ '����p�O_�˼Q�����J,o���b�"���ʹ1�k������[d�<-��	�xC@࠴��rp!��y7�W]Bkٲa(��Zg��D��0�&2��),�>��:?#�-39B����{���c,�~��y��m#R���-�e{O<�f�Z옞7��g���׽����������e|@�"T,!E�a}��C��4.|�o���֢��b�H ;xD�"d���$� �N���(�Ǡ-ϯ"e�[����X�o��y� �����_�:���LK+� � 3�c���6,<Y_�!R��1�������#4�C�C�+�8i:�.7	9�C�ڙ�7�U1��OF����v�%5�^�ʂ���p�;�RO3F��uW/2Y��4C�]Z�<�^�of)Β��ѯ�V�Y[��f+�Tp��9̼��s���D��BSM!M4	" :�1r#��|qP��0|*8a�&I��zi8T	k� k������L�V�a����V�T.^���Aw�J����Z�)���^�HA�S���� ���IyIoe�r�����rU]��>�V�I����ʈ�<��;!��ǟ���j0;�����~`#������M�oCr��aִMd)ힳ�ν�e����@��(>d4cxE��G���;N��@�z�L\�Ȅf�!��1�r�/�c.,21��Qf�ʽ�ć�JVk�>^�6/���H�M��UY�pt�.:2sҮ���knY8����%8�t�x�])�*��0�n���p9��~�LuXU.�o> c3��pd�R�j����n�z��w����� X�Ⱦ�� ;l�0c�X2i�j��:��x{Cx2�����!�M��%�>7��o�hFJO���s�,+�ŤY~m/�倭�,-O��W۱(!���>ih`z�s; _#m�3���#�^,�{o���K�p��u%,�,`��|��PCޝv`�Ǚ�0�_�+��!��!/�1���x5FӀqǲ����{I�L2�h�lȼT����(����ߍ�j��q֜T"�@�S�w\�A+��5�M��f�+�a�G��8��� W=��T4��Ea�	���7hX	R����+�2��j���M����Ww�c��8��6ϭ�m�%�q�����Ŕ�a�{z����#��D��D8�K`p�Q�BU��Q/ʩ.jkZ��>��O�4$ ƚ��)��J��"�����M����;ڴ-��Nl�d@|n����kjOÞ[��kd38�>2��W�!�v~>�]/?��f��]6�)�f���^����B�3n84��l����S��6��"��8�:NoB��\��l�1��|P��{o���r�.��3Ϟ�O@Z�,[�t[>�����A���͙O=��Rڮ>�%
�K\
�ŭ�Ƽ��o��|�� X��B��)~a-�nq����8_b����R���a�?e�f�&�G7�(�𺉔��ޖK�� |���c�%��d-��J��1k#$���Z��E�K>�;/���)��I��9�T�CM� @͓I���1+���+Gm���c�=��!�W��Qz�}� ���D"�`VD�_
��
)8��s�x;'����Z���t�k"���t�W���伷����4����ʐ@�iQ��Y���?ry�|���r��A����;���o[7T�B���ᙚb[o�E+4X/^ya�-�2Qr��+�C		��G�!��;�7�7������ku�� =a���L�З�uBLכ�:x���E��q��l�u�$'�>稯�wq?z�=��?��+] �L��hJ��9nwij�(�^G�fU��C��˫U�F��v%��W.+�K�Z=��u�Y�A�驼m�A/��C2�dwcudK��9˕�-�-lucT��Z:��B�یr�;ً�=����ԂSM*4�@�#M*ҤTE��Q	_��s����~|�B}�	����[��m����Y�I�8��=+^҂^��E{�5v�|(���8�2W�65����� �f�DT�T��;2�<�4ޣ^lzcՐU������bN�P�q\��U�,u�m/A�'����	��=��.��S?�W���+��=9�;�g)�7n�I�8��q^F���L�@�r�5��ↇ9�C�{aRы��%W-��@�-�m|n���B�-��B�/G{�j32�<����횛�"����[�;��,5N�/���Z�e{S�N�LEF���^Z����	m���.z�[佷_Y���=f���~o|�M��%H����`tC�����SY}AE�R-�nG4,�V	��>h���M;%��k��b�;���N�}S���L��aK0eN��q���%����"��9H�Cc�'!K<Sx��´N�@{�`N/���w'qQ��(ׇ�~����8�_�������L��!�W����i�֭�|��͚"�5��.z�0Wϥ���֟���E�I�,�<~@e	����d����z+U�7v�{���FQ���+dj�B%�+n�S���(p�ދ���N��z�N1w���u���_�����c��{v'X5Ί���Ą!�:��ʩ�¬k��*�$��[�g_CQ�������V?M4�*SM(4Ѐ�)���~|�Ou��9���^h���M����>��\��b��=��y�.A��e���DFt烝��M����2�A�����N�� ����`�B/���L�����o��0lv�n�y���f�v��E�mj�Px�@{mS �ȡlP>��n�Ĝ��z�Z~kAcK�צ9���E����vos=l/O@|����3�}k����ka�J��a�V��1�ڡ�I[k�dN=^f�~�����1���:~���ļIW�|G��??4j�����ݮ!}��������6���ex�I��to�\���w A���<y�H��n�9���D�m�;*�cWI��m�W#�ߧS�3�ף��v`X��ݮ�s��g��^��c�s66:W=mt�K�|8��D�wk8��0o6�����A#���깵)j�Q��eΆ�P���^8>C�J������}6�5�sŠ����p��)��[w��a�53��Ф����~�h��4!��ز/��n���8��y��?y|���W����E�D��?[�ɤ�1��u;7�e����Eb�T�i^�B��g)�Z5:��y�Xb;����K��y{Аyb&���B��3�b�P���u�M<��p̐��ȱ�m��*��3�>�;�씷z�@L�p����5/9���J��G�@�M4�4Ј�@ A{^|��>x�@zy�ݼ�Q��-����6#�X������Lz9���ؒ���w%C�U3g1tgU��<u�4����v�׳g�Ƕu="���[G�:/".j� c�����[W[�zg'�����p��x����J�1j3�E���f`�7�-��2/�^K2	�ͺX?�S3���:'����{��pF��I��)�V(UL'm���Ξk=ކ|����M���]R����C�%�7�k��`���j<��Ľ����ʐ�n�J4���nH��c'�k:j�^�(O?5��L��� ���G��-^C�����"�����s�[{S&r#j㬭�����$�5s�����ߔ<y�bלI��Bm���ٹ^}��CP�e.A��5�m��]s����k�n�_����mi�+�?KD&`ג$'��G8���\i�r��z�7/n��i9�a�>�ӧ�@��^���{��F�*���Lr҈�C���(���)�ᡞ��9���,i	��&���E��7�':8�J�%S#(l[��`�t�\���L=����;�o����=�ɖv�+x�U�S���H%&��J��s�M�����YMi*�:�P�cs��mل�e�gE����we���ε��w-��X�6�]j��y�� �k)b{��p��l��J'�ѻ�wz�u8#��&�:�c��M�]r�=9��;���y�����ƨnd��x�c��L�lد;���5�\Es���b�3roN��׵ �t�*NW�J������ܭ��4�ZZ��C����x�u6B�_7����r��t|fr������J�Z��v8��',)ƴ�Y���ތ��6e�]�k�T�	t��x˭
�'\BCF�﹪x!`*�ݱӍd�h�t�u��gjװֳ��5�%����ѣ�˖���-��8��r.��]`�r���њ6�r�����YCv�n��W7��74�I�UK82�5crq�:��[ޢ2�fs6	�[v(�s;��Y��F\7Z*&�0K�Ow���#�]wF,�[�mI���ikrd�L�a���WW�����#)N�ӝ���L�9�]�I׉f<�p��4���.�Y�4��\����ź��H�tev��/lqѐ�ӕ�fH-���;]�FI,v����vݍ{H%��*����n��U������R
^P˝{���WsEA�LлgP�y-珘�F��q���DR�ل��̤<ύ�TX2�l��ꎠ��P�-,����m��>� �YX���r&�Bd��HQ@����#n��#�w&�\j�X��BK��\s-��n���ݙ���
+/�jwL뎠��ګ�VJ�'�]X�y{s�Ab^`4i9�ۗW��uR�s�r�p-]�m�r��LI]X��Ù�(�vj�2��]rpیg�*�4h��jEΏcvƎ�2dI�剥v�EٮzLŢu�u*|j�h5��˗C@$N�05���d��+�';�˾�e'׹�|�g���F��Z8T͍u޾����Y�Jni�ԓ2���q�;ɺw[����\���X1���(��N�Y����,��&�<�vM"œۯdCIΛ�v[š,�J��%��=�8���k*K�W6j=���Yx�,<ji7�V�z��̘�ʐR3vNՑS��.�tĄ����y"�3n�b�/-6�u�rm&��i[��e�)D�k���&M�4h�����n��kk<Sp�u_3�::��s2����W2���o�{�0lfS�Ե�y�ʶ����v��|q�b4���Y��CS��5��m���ŷD(�p�Y�lĲ��z�By(���[o7�SNsj޵���X�]ҝ�q��V9.v2B�Ks0���â���4k�-l`O�ُy	������
a�K��[)�q�ٙ��ê���2q��������$�����>^�*��R)�!rf!e\���\ ��3
Q�1#�roV�a�r�T�p���=k�	���R�V�~��D(�
��A��K��,8'�%��=���9w{�ʹS>=��H�)��&ѱ�������t��^�q�Ǐ?{�~����FK*�F�[E��UrB�i{v�N8�;z��Ǐ<z��ѐ�$th4l}\�AV2D���MIA�m�M��<z��Ǐ<z��d	FBe5,�\�/��⼴QcTlT��! HH���q�=x��Ǐ7��߻�ߊ,F�d������v�&��D����-E6�بƍ��Ʊ�-��(�MI�$�"�r�b��\����y�+�]��6(�6/��E�����Dgu�Dh��IR$��Q���nh�(��h,k�-�c.j#E� O� ��@{j
vAl����?�>��4����3Mh.�>]�� �8�4��z2���j�U,@�U�f��'Dt34�D��e�q��k3kH����(i�%�!(4�*�4��jQDԕ/T�IZ��֯�*1�hDiH!h
����@��T��+�������^�v����2�w�C���sG}�ڨ����]8���k{�OU�b�O���ȼ@z����Ku���B��q�G�)��2�~�V~�' bf�P�ɚE�nv�ёX�4�$�Z��{[Y\z,C��~x�!���x�nn`&��_F��_".4��s�	}��r�ȗ�Z�j��7������s��AF�� �����5O���}>�ZD&*��k�g=o_>gI�u=� �N�pj��5��y��@l�g�3��N0��ȹQ�jŔ�Ns�:���Z�,�j���7!MId�ԑ�בL�:F3��zw>���n9�ӗL��Mig��a9u�z��T\7�y��R}j�@���,R�}1������zV�9���-�d38.5p��ω�_>2i�ѱ����X��B����wKQ6�*E��Y��6��EF@i����~�x�����~��P��|��)������W=�D�Q&��E�b�{3m��wR�\]�ɶ�[A��o@��Н'C*}n�|�k�}�3)��%�eCs� �n�e��Ϭ���R��I74~�K��u^*��¼��c��R���r檏k�x�9�&f��n(��4$���_[����O��Yfw^�������W��H��1W���[����ˎK��j��F&�f=�*�o�D�O�JSM)QDcME�4�� F$Q��#ѝS��+l�1��W4	/�B��_=y������-��� L�9��sƞk����Ŋ�����ۆ�N*J~Ep}.���[J�u�ape��79,�"����߉�V���Tje�g�;�K�'vh���v�
�,�熠r�)�,V��'�q vC��e\��ڨ�B����L�;�ٯ����?��_w����*�ts*�XH	�����&6Ί�U�ۻ�;�p��Xr��XR�f�Le"̊T�3��ҹ�t�kkS�v��2���ڛ7��5[*��)�R]��"Ǹ??��|�'�S��|���Xk4|�5��^��T}۽*������8��EP��9�Hg=��ށ�_i�~���2t��i��to�gyWt8L�u������u����1|�	�_A��t%ϛ"4w00��P�W5sO�;����
*9�X��,���z1�}�A.��x��M���ݹ��ɼ�8R���pr�B,��,2kܢZ����*��܏BN�@! ��/��-~;���-2�j���z��9�.N>�DV���s\�M�_=�H���)pǤ�������1����M}s!�b
�od���z�����f�:mJ�8ԮF=�����n!���(�W�N<�����.��}>�Buۉ�K{�ᙫ��,�T��B�T#M(Mnە�U��v�k�M�k�<�#�e�Gm�Z+�|��q1w4^��t��M��l�q���C�a����l�9x/u >���4^�7�Ɋk�����/�>�h>_?��ѓ|C��)�O��$�+eU1]���2��5�{b�=�~�E"�!�� �Q���^�X�XH�\��
+	~������0�7�3Xze�]q��	�q�Kѓ���ί�����Н�L���N~V>|��㎦}&��]`�i �K���n.�=�K�׆���E2IJaϱ|��Eܴ0Q�!��P`��UP+��͇C�E0Ƙ|���_Iw�y.�"�R��x�T���1����T�]W7#���](3�P�9��m��05��3�&�S�>9������ʂ�f���T��ǚ;Y�Q���!n%��P�~hP>6����{���j�dQU{�gC3�K���Sn�4�ޠS� s�}�����Xu>3�p躇��ɑ,bj�M�Ǽ�ѷ��3Q`�S�+����b�V|��ט�5B7u���F ������j���E\�Fe������'�(Q�Y;\v�wU��o��:�ǝ�d�Tw=Rv�ٍ�d��c���R/]Y_��ڪ���Ux��:�����.M�
uْ��y�K��W$�Eg>���"��w*�T�6�i�!-t#�(>�E��@M4�4�B�M4 �QY��+�~y��$�W�����4v����t������_�9�%`�z��ztr�n(��F��V����������#�e{�MKD���<�o �:��t=�[��}��8��)�ǌ3r�����A�_�/��iX_�	;�/���5��[i�l�Y��=N���U���-7�n�4�L�/\E���ʿ����;�#�~�P�ic���>qW�q1�6��8������B�v���z~H@/����i�,���ƽJ�0�ǟ/��)J�_�����9�ey��3Ť^m ����V�Mr�Pz6q=c�:��)�=aų�,B/?C��[�����vM���~ߨ�����S]�2�&��%�.�aG�1���oN��J�G�e���m�jv�yZ�-1��	�J�{ t�3����@���%�r�/xS��B�(�|�(-���dO?gD����A[w_y}�82�)�\fL�a"D�#����������ʑLh�&�i܇����wַwL��WEê1�:zބ�"a�2��l�*�L��)?9�r�xC'0���j�}�"cmo����;Ӥ	j�[z+FL�α�CX:1I���[�m�$*�E.^\���9�Q2���B��)��P�Cb�I�c��qz��t��79º�ƌ��*�+1���N�\�EIص�yN�޴���;��&�U`�i�K��m$I�����&�sG�v�*�4�SM�4Э@�IBAVO{�"������r�����D���j��|�<�-� ���Bm������Z��dZ�����دnQ9f8W(j�:���'��+y�mx�a=��`�ь���C���l�gNrT��D�uɎ��+��]�r���^���6;��K˼|ga -��n�*�oOL*j����i�u	�)�/�%�F���I�Yӿ*��y��A���lg��@����u��7.��4i`,-`�>k�;�z���0%c��xm��X�z=&#�D0 �C����2s�����vđ�����ÆpDsuy᱉}�d�fg�%~c�L(qh�1˼��E��'�z�t��JƖ�|?��HiߩS �H�~(��Wʫ�^��/9g��O�c�Y�kuK�3�T�Gx��Oj�K:�b�f��z�a�Ӳ%�q���)����
���Y4�t��e[7��{^�H� ;����epz���'>f�t�O��f(��8��48�0l	�"�j�+[:eEa�\�ݸ���zn=3QM���֎��K%�3�g��6ʇ@�t���ٶp��F�q�9v{��\͟��y��}uv�VѨ��Vwp*�9E�%�ΙQL��nQ!�6U�/s�u��=��C�'��Q'�������'�c�vfvE(u�bJ��U���2���J�"��+��5�o0�foz�"�G饨# !h)��B�F�E���7��V9G����wv�y`��E6�Г�_l �MV�K�]X�����":e*B"�#*�WJ�O�F\���8��P��L<s�/l���#C{΂��i�
R1WO=���X���_p��Fӥ�~u)Xol�8Bo'0.*p-�8oc34�v[ly�QK4�h7M׼���#/Hr4�)�ldzm�{r1�P���H{h�t\O�x�o|�7G��nt\���[���wgeF�{��mٹ����	��%�"hS�_;5��>���i���U?w�p5�u�����[���P��vܘ)��b����S����I��S��#W��>x�t�N�6j���!���2/��Қ;h��=Y�¯�s��tã*e�"�H/��1*���l�/M}���L7�C��C���ߑ�F�/�~��1"���TXPY>޷cx筘m��(ؗ]��ESE�����=;�B��m�Sp��95��`J������NTjMvlL1���\���}��EGb�>���iwF�<��Cc��j{�fW5<��m��b�H�J���Ɣ>�r���1�����{�������6[���y�1�wg	�'z��:[�nK��ܚ��V`�D�}����g�<�x�U��\ws9�I��'�����v�%�����+�<�����~4-AR4�PR4�E4ЀTI$�$@�D�AF@~fw��ϟ8���3��`NW�\-!��Hb��Q*��H/�*��ٺ�!w���+�s��6�vl�Q��7�KϨq�n�%�3k�&�ߺ3��yw@�3C�2��7P�a�v�	��K�:f�W��ۿ#T�;G���X��f��@�c��j(	s�Dg�w��9��F��;!"�L��,p���%�ޚ�퀁W�Z� ���B��7GgP�/E�n����qS�n�ɋ��^Y���bU�ĂD(q1�5�b\F�H�ĠSm��y�J�imT���?fς��Ԃ��.:k���&���a�L��q鱒ܟB���D�ۣm
��
[�ds*
O~U�B��u�P4�a�Q�<��E�Cޭ�]w���pq:���Ya�����r�� 7����ۢ�0L댎�����������w�)��N^&��;�H�5M���w�v�c�
��;fQs��,SߵE2��"*�3�����W}�T��۴���T�XsH���|zB�����]7����t�)�q����m���,�n^�����ls���Q�P���"�ܙ�Z��Q��-{*��w,�����h�MoNϘ�f������:�R�,�nXb�}5v2�m�b����ս��tv3��풟{��K3�?M���.���dD�Ƃ�)e(�i ��V�(E��2 �v������E�<�^퐷���a�m�y"M�N�{��1i���m�E�஗��Wɹ򕵡fL?5�?kB�Q�y�`i�?Qs����0�z��X�D!C�5Vl^پv.��6�7.�)4sW�g֖שL6F� ^��^0��=#�#��?j���e���H�g�t���B۔^W0�&V�{=�*4�Ot��L��l[��G@!��I�*�v[�z�[X�r������
t(������/ֻ����2����U���f�u�����*����<�t!zl*�K`�~���y� ޯ(5׷��=�"[���q�Ű�U�}�vd�Л��^�&��A>q��0xN&$��ܾ2U�����Q��{I�)~4~>�s���v,�@��I�S�o�芇T2%�!��\s"2OB^���O��u�'$���"��Uפ홳�Xn�GO;�ǯ�r���)�|a��>a�w�������=I���5����B�a�ڲ�B��*�S�$g�B76u=c�:�,'¡��z4����|��iK�Lr[%�.���_V׫�z3�zoDI����G���=t�(�Y®g�����&���N]狽�~}��;iPk%aʃZ
�C!��n�ؽ����&nӧ
�J��5��-Q�L����w�;pS�i(��`�R!��E?�����i��)��i��(H������ S�5����~{�l���|��<4�3�ÚD�y��O���y	��Ʃ!�PY].�a��f=���|�ݳ1j.���i�ۯ7�Q��L�����е�܏[kH؂�
�D����(�ҩP�Q���Ad֯n���߯\t�~ҭ_���:��o�1���!��@���tވ���R)�ús�1�Dh��X9��<�WW�Z��A�ˏ���Oz�̕xh� �SPXd��.�{���g���b.����ȅ|a�W<��1E�5�/O�獋aAG�Ȅ�YL'�<�.볮8�QmY����:��[qv\c[e蘵��S�-"��Fׁ٦��� [W�B
5��q�1�
��n��>RӠ<s�Z���U��\�G$&2�䣹�֣]ĳ��Ƕvo��-z�u�h'�P��TȝuS=/�#v���b@��<^�G�T���طp��_I�"��$W"4��ww��;�P<�Bo-�T�E�_�f�E*���n���I��Q��4j2<��`�����2h�Q��+lL1���C�,�N4K2|�2+�����������Kr ���nٯM[��=/ϒQg���������T�GW��"��;�\Z=�[G�c:��ٛ`eY`g�k�����CHZ�A�u���͒�sUJ�"��[T`�O<NԾ���n�w���_�������$�u��o{�t|}~�U)�i�j��
i�Z�"��=�0 {N�|YCR�d+� &�H�� ��?��XQP`|Qc�4�ֺ��M^I�6>�����槍�Q���މO\�w.Œv`�<��{g2ȗx!�4`��?a�g�S�����G[9�l?�WJ���zU�N�h�]���.4�{��;�(ޏ�Xn*�yq�*�~F�v����q�QL}~��)8�r7�Pj�FCO���.qL��K�oF���)Z��B��"X4-y�;���ws�bH sBP��v�	��E2�Z��{��7��*�smm!j9�.���?B�Xs��U��1>�4����,7qv����Y�7
���E>DJ��+�Q9�f~��|�3�^��+�&}�C�>����`�8R��x6��]cSP����R�}w�o9%�d1`�y)�ߣ&�N�[A�(��^��4�Ӥ�a�e:�_`����6�N�������}��&��K�&��q���A�-ᄍ�l�BcET6-y�2�z�o�>�C�5з�Ei�mɎ/��2.�eh�-��՜��/̯
�����x�P�ʋ�����qSǲ�J"��w��rV�Uتb[��;�N�;މ�_7p��0c/���WB�Y���4Tw���ĞV* n���=7\� z!؎dBc�)��Y�k�,:39�T�m��r����{(D.�F-��Aӻ~�E�:�or��Qj����Q3��L��x1ی��t����MEֶ�m��&���	6
�.�w$��r��!��9�����n<o���I�-9�[�U�\�X�+q���[�|,<���B�g&�1��v�Xrj�;S�����G:����e�Q���D�Ւ�tL�b���M�;��r�6ݗK�I]���rVl-��%헣��L.�s{�W"�����r"�8T�CGK����k�s��KU���Y�+�X�m�ۑ�θ{��hz���g-���0Vt�%�X�^�мt�fWr�L�Ӯ���7��q���x��=.J��qn���E,%��-n������Op]���U�ml����»`ٚ�=��+(�3����HK��.�1l!��1ʜVv��{\��3;r��,�Ά�Y/���G&^�To�my�wy��g������o������<��{�D�-���}{)&ˮ�kaˮ����}H>���-�|��]�蚹���0�<����r�LSe#�^�3��L�t��x��uj���C�*q~���E��v�:��D�!V�esu��������,+z|H�㏟h� cn��h�0�8��-��0Ec=�J5û�c����4��b�������wU/��X���^Cll�Z��4ɳ;��{��76l��v�S���p��=棒��U�*���r�Q[��M�H������lf!y]�뇓V�A.iz�ԥP����zW�'msW^�[V�!V�L-Rh8�������3ؚ�����2�d��p|�c,h]�"����q����_g�� �W����s5rf�,�*Q�u�k��x��)%������U-�o���\e�UiO�9[�j�³NA�$�n��յ�y��]��Úo\�yD�)�a�aL�1�\��a��\��y8���Zb��6qz٥���ܧ�2�x�+���o���=l����[�++Y��W0E�51� �+��$�mC�����;����J������ݶ�yմ�V`x=J\2v�1e��K3�B����{��/�-f&)[U�D��V�W�O���v-6zQyU �Ln �qvb̍{' ������u4�B�D;��ǵsk`�i}Ӛ�a�h�!�^��9�u�ni;ܒw��;!�MP�5�_~��j�c�sE��H��E(�D%�lX�۷���ߛ�u�<x��ǯ^�bH2$��'(�ch* �Y1F�d$CM8ێ8��o^<x��ǯ_�[��1�QF���!! SN8�8��׏<x��ׯ�~�EI�lb��vM���-�ߊ�1�ɍ�����7��q�ǯ<x��ׯ{ TIG{��hn�#Q�ߋ�#F����ۘ���W+�j6�j(��%}�h�Y��r6$�Ѣ�)#h�ӛb�cX����}-�E�J�� �x��a���4.ʟ����ڏ��A��P;]�IQ7z��:ra���S�,�N�<�h96v�7�>�_��
i�Zi�*$����*"H��!"|��>s�\��i~t|���.��̉��_BaU}'��˔_Jq��r�a=K'���Q���H�Ǚ9�Lk�w�[�� ��K�u^��8"�]8\]�TXPY��j.�dTܽ�풛zgU0B�YW��ۼc����|x��^6�=Q�?K�}^];�
A��O�qe��|���n�����i�����9�8/�|P9�D�s�Әoe탺�ǣΝ��o�˭��!SGy�8߶��}��"��x:ǒ���C�c�Dʥ3qK�6{�T�)�_�&S�?��_���H�'�׼�����ƜS9~�<��J�d�tuw����A�=c�yOl**-�&�K0�zh��ݾ�9D�^�e�o[m\�n�Ȕr�a��R��f�q�N'�p�Խ[�U��[�yl�K�Y!�k�15��r1|���ϙ�ɷ�1p��=�y�I��܁E�KǙ�h	f��1+��9G%���������=�~`��c�8��b�e�n\��xB�XP��.O������]7/��vf���j��Xm�-��C�����wԺ1���{����̉�t�	|�f�1��
��5t�Z{�Ә���s.�QYyPq�\�P[�V&��zq�?q�J�گ�I�Ө�a����uo���u��3R��}��G�j"F��i�������q�\��O/~�mw�!2X��.�g��=�3߻�7��U��=��(�=����[V��z5m��+��x��5�2}��_Z��m�는�5B*�dlf-�
���W;���ǰ�"�9����=��Eb@���)_�׏r���߼hc�v�$�[�X��QL�R�s�l�:�Ey�]:ՅT��e�5ոx
<.DG0ƟC�e>=!U�0�/%����ybh��\�_\<E�5� W�7Z�HO�J�>azyA8?�ף��O�ҝ�Y���n�k{1P�Zn��B�Y=�C��i���{n	Ĵx������`�Ꮓ���|F����O����s��z���]��"	�1kc�N���V�O�ʒ~�&>H��2�(���A>_�H�~�O�W���H��������N��?�Z��R��J��T6-�����]�n�mP���\�	�ϐ��MB]����Y��cK��eO��W���ۑ�!����4Z	�V��M O���z~\|��=�drx��dE���^��]>yv7��Z��N�Vk���fĒː�Z�r)�gZ<�e�eaF���B�n����r��Ǜv��זy+�� �S��
_�u�)���:�-[�1G]nWf
Ŋ�Iϫ4���¨c˕ßtu]i=RQecNMH�F���ɳ�$So��l]:�P�	TQZ�*�j�������{v۔Dݻ[�7n���ZjA@$]���$�+�9������I%���! �H>���x/�i1��?��ht�LM͗�}��W�`Y�a���\���!b�g��)�d�2��i/�צ�O�]X�L~����y���*U�62}Y�+��M^�>m���"Pޝa$܏�rCfT�|�*8h�9����~^��S�8�Q��<��ꗺzh���\�O��_��`��Kh=f�'����N�[<F�u��Y˶�ic��Be�O��P�k'�y	Mv4���D���N��ã1����ښ�N�nM/��)n6���\"�d�O=���V�� �>���/`�4�£B�v��<FfZ���\�����ȧ�x�����5)��ꅏ��}�DIu' t���Z�^����6��7 +ȸuC���j}N�����`����8�<8`��rI�e���]���9d�s�_<�T��F��xض'�a	��86�!�ކ�_2s6���,�C�%�|r9��1i�by�y�iȖ�推��tk_��p�N��4��w7�9������/\��Um���[��f\�l�4�a;���\�t�/]�d�gbַu��A��Z��}U����r<���^
{��Ʈ\��'p�[��-V���Bi��
�^|��k�[�o�w0����sy�D�P��e*F� ���,i����H��H���{���=�N5����ާ"X��Wй�H�|���w'�bB��b�\,�,Žyv7/S*:#Nb���*%�1�&�"�p�a"�o�����QN,-2S��g���Ű��e��Ze�:�G�wHծ�K�g��C����z��ɳ"�ts�78�c,~��O��M�Ϻ�0 �E8wv-��������#C`@�¸�H{��A����Ǟ#���6��o�o돯s���*|}���;k�QX�h��|���X�|~�}�룪������׺Α���v�z3�>����E~͂$�*0��>7��$>��j�U�?�o�V�����i	Ze4��{[�!���uǶ�#+;=D�N(7-�b_�׹��"b���)�^I���c���ɱ�R��<�؞��z<�I�\>��Ÿ%��P\gY�ͺӌ��P�3r��"��2��Y��y�3ЀqP"��y�=ہL*.��=�Г�_�a��P+��dS2T���\�:�}����n>t�������~B4�O|��`�ƌ�����jt�*Wu���[��3��7�ݽ-W2U�M(�u�л� E�s�n�^]�e�T��]���E�t���
׈O�'��^sD碶���G��a�w�%�8�nfͱ��p���#�uk�xѥĩ�$�5S��c{Hv�����������@"����M۷57n�ZŬU��4����[.�3}�+���y����������[>x ��EH����/ptiD�"寲*���L�E���Dkf���$��)°��d�b6m��E�wF7�H{hN���,:�u�p�V��l�偊����d��:h�y:��p�H[�Z��ϳ����K۾���Qv/cf�-���)���̄����eb���rc���˜��4�iyv'�]K88�)C�\r�o���H>���\]4��pn�Λ�Y�=WԘUz̖�45�)�`�,u'	�l����u�rx��P�z�H>ֱ@��;A���U �:�����}<\_%��35�����Z�3no3�����_(t�&���X�Z]�B�M�01��d���n�OOа�Lxӗ���'_1qqǣq��s�}`�\�WW�����fr:L��8�s5�/��{�ʓ6�)�4����Xs�v�\E��v`$�rɘ�34�k�?sdC��S�/�
K����I� �ޟ6ю͐+U�$�0����h��^�^W'�_��×���(��!�WzJ'�)�X�Φ�?EQ˺���8��gs��L`�B��Qou+�L��jC���D|$��[B�3sX{�S	��nA���*^�M� ��3����xЗ<!���]3~�{�,���g7S��5��=~�
�ijF�I�T�(�W�O�/y�|��|�����G��+���:u�A�Y!��12Gs�1~b�ó�bf��j[G���[�Ń�y���
3��`L�"ˉ9)=˼L���yYؿ~Z�8X����~�?�N��'̒9}�!�!�^iN���>�3�~a�:N$E��x���-��g��/��2�f~��=�ٌNz����*��	0m��l�	��T9�*��i.�V� I�c���/��+u>3S�ĝ]}����Vƶ<�Z\O�l�yGw�HMո�R{U�B�E�з�xjkgd�%���+u��豄wY҄A�-���kH'���S� �LP�U��f*�e|�%����o�_ג����.wTcG��8S ��u�CF)�wL�s��%�~��)���I�\N�|�(�nv.��v������f�S�zæ�!�1����K"���5��]u�v(.!�R�O����k��¨rsn[g�|���4 ���F�צm��k�ԝ�ngc.��.��g5e���r�t�_>������L?5'��C��/?��
��VW���>��]Xy2�7§Z�Ѣnt���"$�nТ�ٓ6��ND�r�7b�����[�cr��G�iMuo�\��X�~gϯ-m"�4-~�wN��jT{��!��{34�X/�Uw:V�LS�̹��r�z^ᩝ��y��!.�ꆵ�ej����Wzz���z߅5W<5L��5D���,����h�ƚ�I$i�*��{]���o�݋Q;���6�E�7�I�v�Q��,��{XՄ�����^��N����'Xt�y��q%�� їYM9v�5XO��bgβ`C��,+yN��J{��6��̪ e�[����m)u,���ҳY��žd(>�ȇc>�j��;���O�|7Cti|��}8�	�b��{�~q�2�-#۝<9`�< ԅ�Hv�������PRӞLZ?�X�	�+���=_KN�@ۮ���6jZ�9������o��8!��;�����%M����J��C����;�Μ�e�l�Νʩ׉h
B]N�_E���a��Ȗx�!����ȗL���OO:@��d�3=�	;�:����M�)��r��6���@r����N��3����i(�G�dQ;�i�Lz1�S�n�S���2��&���@f�'�1�OH�sY5��7 �k�dޟ߶���y�@Q�E��h~/^���OD{.�S���%5ޙ>A����I}	\�xP�1���rr� �R쭕K9�36�qD�Z*�l� Qu�7=�00@_7;��41,��)M21]�ݑ\���H0kjpM�fڢϞ���Q,N����q\������V��^;*��op��Sc��j3v���"��jK���sfQ��b�L���e0�QV����{��ݾ|��d��OC-ٕ�;�|��	�uϮ՜n˾s2��%�1�j�$i�����h�� 0e@�T�CjP�}����c�y��x��4S	�c�Pq�Ҟ�q��-��sbb��ɞ�F^�rqA�RS�ɭ�ܑ�����= ���JC�I�
�a���F��d4M�ٝ�����Mmn{�\�j\мԡO0� �av����(��Bn�|e�T�G'.3��\G����Wl�n:e/��>��G4���F�;�[�l�\¨^��u�Y!���Β3a�2���H����=�B�P�����e�&2����� � �k���IUީ��2w�*Y��*���C�q��:ꥠKl��{Э@Y1��)��_^����O�E��5{?p�s�l����oN���k	 ������vt�_�x��� F�<���DsF�J�IG$��?f���<�϶�ǚ�؇m��h@����qa��t��e�������yṑu������q���4&����\ׁc��j��~���AM�Bh���ݬj��򬍱W���l���Y!���do<<aۚA0� \�5ퟧ�-�t;~��W��Z$ۙ��dř�7i9$��.�qE�p^�
���yN�m�}:��v32t6f
#��dnN�s
j���\�'�T��W��~S��� ��T�Ir���x��'
��rX1B/h�%��S����ٕ�y.�3533���c��1�ʑ�����vA%a�7�&,�r���v2<���C}V6$�I� �˥�Ͼ� ��S�'���8�2�s�]^Eb�fPS��V�Vw�[��v_����^�k��U5�BF��OJ7ǎ���,{�d�g/>,��0�]�1�F@F��t$�c_l ��K��&��.睃z�6+�S� @	*\���T>W@fМ]X�/���3��4�|m(h3�\4����xl$N�i�����M��Y�%��NV)�*��8���6��"���!�
�]KE&
;X���kP#S��˞���Њ��2S����kP�hT�z="}��OavaO4��uB8��(rf� n>��͕)�����%�"hP}�Ks�w�xo�Q�z�8�9�9�0���������}�K+�l�<�Ɋ�E���M!iyF��<v�Kb�����osT�.��!;�@���?t|b�1��xY��=w��6�Nq�s�c{\�P���Uo����O,~�~{�O�~V��/��ߨ�	3���D�\��u5��}<\_�Y�!���������M;�狋�j����O�4��秳��O�巄얓�j]�dܵ����x����ipMU�4�)�"@>��Zݚ6��l��c���J�����U֌׳sjwzi+huZ��������f9{1�?_���a׼����}�~ڦ�Ɗ
ebH2:uA�e��S�t�̩T����K	����+���G�������������˺�U�e�|��9�8ǺV?�������i�Q)�>�G(���W�z�����=aK6
��!���W�K�ԉq��8����[�;�/z�4��Iz�GHf{=p�j�Z��/CBD[x�n��3$���u��
�Bϗy#�o��>+�'��ď�&��.��̡�I�F�S�<c�|�[�JVEO0�������]�yE��;��0ist`��F�/�H�^�vB��m�=OL�`38AA����De8��I�Zq2↜�s�c���'�����Uu��ڍª��H#��6�e:j鋀Z�X�aI�ܰ^׫O�K�����]�9�\��i�ڃ��C+ܟm�Q�u֮��d��.6q���C��@^��[��Ş�����pZ^�[5d�7�&��^��-R'�?��(.x��[ռ4��<>j�7�Rk��ű�장A�5��
i�D��^!��kk��z3ԡ�1�N
��;��<��{�x�-')I��^��?���d4�q��{5K[�`u�i')�f^0V^�/g\��o`�W@��Tym[�k��c����t�]Aa��:�R�t$�t*��y*�rt�:XZ%�1��3kh}�f�2>�5|Ϊ�u���/2�^�S
Ư\ɸ���\��U.&':y�e�s��o-�����>���f2(WN��������n����R�4<j�ϥ��z1��fME8�s���(T�
�q�f��u$�7�o��?N'�7���J�/o�)=��W�t&���7F��{�㝕U5gL�;�(v�wIk(��ܫ����Gn��p�D-!'�s�i���)��[}.d�]vt�KùF��=*^��!�d����I�-�����^�Fl����P�4��`��k
�jT�n�F*a5��cfM�����8���c�����L��e6�����歃=Eh�Z�͠�i3���cc)�$؂=��Q�1b�;��ҭ�9H���L�'�o�2Z�
�&��M �M
�N*�kʥ3m�)�Q,[Z߬��ˮgn�lO���.�v*enq&��gTk20v�����fڬhQ�rA���)i�Tw��_WN{�uH�4c;�4P�pv�ӂ�}[��t�t���dT^�6:���ŧ��%7��D��hJ�U��,:[7]�F��[:؃��oa'���c��Ւ��t�yF�аv
�E�J9h�2[:Yj�'ځ�#oyT9����0��z���`�ixf!+7`ԯaÇO�����G�T��#ΕZ�V˩�� yz�|�ڑ�7|�n��_IV��\/J�{�oa2��x��~��Y�充��[:��6d��|���/2�/�F�X�>3^ݲ&б�g��vKy-�����k9���n�Ep�B�a���L�2�9,�:�^��jG��wv����%��ū)YD�h��ە�����`��FW^ް�����($�0`V�q{2UH��<n�ͭ�L2(*�G�\;�Y��<y���j�b�g�u=�rEl�s5
����&ɒ^.����Wl�5*���a�㶑�I���]�*B̡s�nU٬�ڒdLn���Zgb�,�j�w��-���Xrd.�S5am
=J�nB0X�3w#�4�3F��ri�z��ƫ�U��n����z����mt���b5��z���!���Ջ�1��drX��%
;˖VU�ӄ�+KN��F����N�=n���z�\�fS�T��I�̋�J�Mۭ��#�ղ(�o�.!�	c���F�9��&q�+׍s1�^�1I��	��U]kK65}+�V�X��VRH�f�����4;|�+���6�oJ��)���
/����TF+�B���zi��o���f�Tr���/2����{t�I^��s����81�R�ᒕ��jK�풹lh=��fon�,x��|�G����SE�G5.6�W��;����'ou�H�$�l�}<�&3ܻK�J�R��7�5Z�ZqE��­�5o2�۞�0�R�k�?Q����)Ba�CQ�ڢ�$رuTS,騊�H�o�^�J> �Jd��"J��Q]%q��T"��^r�wt�T(��2�~�@J&�>޾U��"�W-�b-�W��B1������<v�<x��ǯ^�vH�eD	EI$c�N8�<x��Ǐ<z�Ό"20XH��"�BQ�N���8�㷯<x��קbH�N�
� j�Z����UJTJ� I��N8�<x��Ǐ<z��A�$!�I
��kr�.tߋr�cr-�E}/?��*��;�r�ۗ#I���[�2a6��ȱX�|��(�k�kү;z1��ѯ5�*"��*�Wa���2џ}W����j�����dI�p��IH4���oH9�na���U�����#��ܴ��MA3�k��)$��q`�#\�c��e�V���t��;@�E ���J�w�U$5�M}�?����h�����> �	'u��~ϳ�:U�K;Y����C�h	�|�0y���b��v!:�X��U,����eA�W8�O;JX'�ˊ{���E��F���|�PY ���s�%�	ὖ�,��[T��#��M>��ʁ�C���1�^hL�� �p��ǽՎ	��Df�Se'�E��w���zK�N'��g�,it�~�8�`�z���ό0t��a�^��G?�EB��QO�X�4������C�l:dU�*�=��f�����4�����!Çm���,�bc�1w�?� ߗ�/�C�R��zg�4]���I{��PD�c���֦�����>e4Y���`��:N��^9�1�&ھ���g��X/��{>�{�z^n�;�2��+���� �=v9P�t�D,Qz�֋1�d�n��Y(��n�K)Uͭ��%N�D;=��nl4Y��}"N% ��	��~�����]a���sG��
0�K>2S����9���Z�s�c1�z1 �L|+�{ǚ7�����î�+y�@�
~���k��K�c����3����:�}Ien��U9��e	x�'�kK�8�.?����ux��ǛW��ݜ�Ϸ{�ǭ��֔�ׅ����%勍�$����v_m�O�p,���:�X�w$Ȳg<�h�p����,f�:cl�C����Uܹngi/��� �j�����iZ��$�;���I��xZ�s�tǘ@s�&�e0�M�#LrW�iW�ܥ�f%~����}v{���*�fl,��l2	�5?X�����g%B� ���%8�5y#����G�(�~3�|�j1�7e��	�R8�;�D�;��+��B�ˈ��zY�L��[�o��=����j�o��[�j��B�(|;�`P���?~S�c�����a�.0i�d��!�T�0Ǫ��C^N\�c����6o�I�桯l��i�rf�V)��O�Ũ�XƊ_�8�&������s���j�]:�ʑLh$i3��6�v�\���<�@0"�����.ۘ.�p�0 �ѭ���c��"!�g0*i�Rg�Ăh�/��&*��Q�%E���G���督��<��)�c�v0X�:����&n���[�����2�,ŧ�T8��>�S��L;�_��pKZ�̲	FS�=��Ō���!�q���eOS��{F�@����t���'�q[�Q�ӫ������D��/�;+�HT:�C�;S7�o:�D	m��Ͱ:��߬~P�^��Y0����%��}O�g��!�ڪ����3�+����7׻���Ê�齇��ޑk�������u����̭����1̫�r�T���ǰ�q�C�R<�<�?����N�WD.�[2�N��N����s^s9�.����i�
j�h*2��g:���/}F���;z��xk��"t=0�C�<ñt^���Y�+���X�0Y�l�ڃ\�h�@�>�
gZG嶽6�Gf�
Ё^�_ǀ^L%��ɳ'�n�[6�_��s�ot��*���?u ~�;���Bx�\׏�
P:����v�
.O#؛�2���\�K�B��7,��>=ٵY��yO�9��	�e�<>��{��\���t,����~5��O���]��om��Ix����5�M.{���N���j��5`ޓo^IzC����-��6b��ye�1�ȝ7�<���^�	CF�;�=�d0��N����<ۻ�m�,�Ark5���qE�L�!�PN��m�g��|�̽�!>�D�c�oc��h=	>2���j�F���CI�3ڤK��%�I�$���K?؅�����|��O��t�ɻ/��r�� ��mꎝ�+��hk�u��
W�U�#��u�m����Op��4�Nb���	�-��b�ʅ:`�O�)�>C�T��]YJ��{ɔ�N.�6���{ǔc[������Yi�X%��V���f�Se�a;�Z]A�8C|�g(*0Ut�ԙ������~]�^�^�;�U؍�ue�UbFĸx�����U��z���Bj�"D|�oh^jr<���k׷�Q�Ā��bv+egg�׎��<||||��<<��f�Kk��+���\}��@�a,ȳ��ͽ9I���^�E��M�ؾ{��-�eC�;�����c��	osB�gb_�`�6�V��`ܩ��	�d]sl3Zv��ه��ޅиa��B�%�?����/�:G�~��\sץ�u��ҘMoI�YbD��y�;[�זf��,�.U%<;�숌�w���y���M�����uxE��pED�T{�u��z�K�A#E�,��5?G�~0��ɥX�ׅa�&E!��z�s��k�1KB��Qօ�Y�6�%Æ�_'�&W_��r�^�K�(�s�s���g����^�$������k!�`��K�͵짒�4��T:��Ǳ��������j{xC��A�������	��F��������2ΔG����V�,�ħ)�9ǀ����*�N�͋��Xz��p��\gǞ�E5>�>�	���5>XE:v~�`d$8��ioK�Oy�~����/OV��o(����{�|e��zk�x�?X��A�2�^9h�R���^=��������ˬ5�����c����'*w}�wt����SP��"�S+U�#��"�zT�J�Q����gz��!�W��lA�R{{�n�C2�t%SB%�Q]͙sporʮ���2�Sٹ%����=)�e�҇M|�q�����#���v^`���M)��,��#�^H��!Z�ʍkD������Ti�B�+��Yޘ*���q���Ǐ��Py�r�"gHV����=�GB(S��Ͷ*D�\�ym�/���o;�^�2E@���wd[P܂ٹA2s=,D�kD<��6%�~li�V��0��6!�a�e#@����Be8L��b�)�nH'�1�[ռ6q���@�ڼ�;���b�� r56;���|��S	֭�����4���LP�USZ��ȥ��:km^lT����g������f;ﷆ���m�5��,�K�����/J�t��Y�կ-sZ¨��ؾzf���*S��o��`!�2�o��ﭥ��d�RS�e�󟩌���Z~�9���uL,��,��ó�y�!�~�h	����1{NC\��ub�C�U��'�]�������'没2�I���X����`鱘ч-/-��0`ƌ2�e �-e	�ư->��B��1���5��U���|Ɲ�N���#���c�C�o4��C�0�u���&gqϺޘM6џ;H�R;���7��R��0K�<���+�`m��EfSl��WN|����yf$u�x���W[�<]lm�9�ei���OLù�t�ow��U�{vֹ�aLy"�C�K�d�9'S�-{�м��V(�q������X"�g���.5���ҁa�N��Ww�vL�뢻&{�������ٖQ��9c	�T�!�x:�1�p��r���P�O=�g{ ?���@�ƻ^���{M�d�j�B�ȑe�E��٨�f}��z�5��3'���VJ/���e,e�v�͛����m�qԉ�@�)��u�v�wyBc�NE���,)V�g�G~n繢¥F^i�ƒV]ki�	=g Ѯ�icD(A���.���瓟�b����>��!��I�����!��w�TZ{��`��Bhf�`ME���\�+;�e�E�7k�>��:Ѫ���oR��SH�	�/�c�Ңښ���
�dʂS�$rC�E�o$�k}c<���1�1��dĂ@�A��{�a�_!�PT��Ǫ�1������cL�ɫ�&X���k���g�f�9y���	��Z�=��^9j��J�b%��̰���@Sjv_a�.9�h����Ɍ"�+z�v"�N|�FXV��y��m�5{gO"���x	���*$��K��8pG�����vV�li8�tF�k��j 5\:�r)�$i5����u�����[?�)�K�M�u�4�g���{�t���l�=rw�Web&��O�lۚCm�8n9*3��'=�˫�^)%��""�-��M
єRإ�f�-��p�/wa�ز�(k�ՈV�xe�o��p�Z�]nñ(ܯ��O3$��o*�~��J�|c�1�o��j:t���\k���q��f���\9o;�R��"�RXsw�F��d�$lLqa�;.祶�������bȸ^}Z��oc�C�zOȄ�9�f�^;4�����-t]m�I�M
��E�8~�k��'�g�	�7
��;��'G$g��t��yGp�T���sw���!�&�t�+1׎��,~?"7��W��c��ݍ���n3_�9�&˕]�����n�@Z�����^�i�{���9�m�v.��y�l^j�B�{��2h�����f�jcۏ;�?UMK�bN�H��P+�~<�2/3ܶ���7:'�kg,6�_��?��Ig��L�,�ށƹ���<�j�5� ��GmC�WZ�8��"��io��+f|Ϗ�e�.�GO����C�)�cT+�)�øm����W��eR�3;�od��OBj;���9�dy��Mf�/B�q!�].�)qaR�4���U6a'*)Cqt-��2��	X>b@>�0 �����N��VB]��w!�K�Хɪg1,�|�j���^�<{^����qH�9�e�r)�s�9	U����QA����I��1/v�g;F��A�)x RD�01Ggm��\v�l�wmo�M����IyO9J�Y��)�:�&�=����_vU�˾���3�L�o�x���7����{�5�ab'l,��2m��2���W峒&���X���JD�踆=6��N�7�VD^��]/���	��	c^	ufy�f�l��s��Ϩ`��>/t�/��V����f���]��t�(��?}���5��W��	�,T))�a��c��.C�S>y0�L��X#�Ћ�Tm[c���Ȥ%�s����n[[6�s
$����aL�P.#f�H>��ƅf��y�]Cc�.^�Ɗ���Xb�����Bڀ��S�`l���R���%�K�&����Ml�.k���j�����.ѧA���	�,6$2�!�~��G=�vW��ꆁ�S��L["�x�-φ��T�eu��w����YU�(7���B@�iT�C�hG�C-{����[!���0��^h���}���i iᖫ�/~*�Y>M ��G�X!|v6>;ʢ��Y�d���U�[W�:uM��@���������Ǫ�=��sӼp���>6�!��
��w�V˦�î��e��`&�Ԋ4�<�P�ҫa�PKջ��8���Nr�w&P�'�w���qѿѺKzev�@��������a��͂;�VMX��.*��yڽ�͘C�y�\�"�Uԍʒh�@I�`ͭ{�6�ه7f�^���2��v����;�UwO��b��{[W.QʠM��e`����vJ���*4 ���q����������@�s����0n��>vB��i�C��S�M�UM��o�c+����=CZKl� n\4�%�7FM��׮�3ʫ�:�Ƽ����ԉ��lDǿ�����%��a۱�P<ӣ{��78Ǹ(�h���@��t�5��
�Þ���a�a��F)��y�W���\�Q�]M�U6g�	�C��K�f�c��ָrv����6����������Uj�{���)C�+n~�﷫f���-�(U�$��c)^�=��M^鋇�yg�b: Δ��C��KOL��ͪ�ې��K�$T�h�ж��г��g��L�a�~�v��N�^9�<��뻖�]�F��%�]z\Q�O���O�xBj�2%�g�)�Jܐ@9���p}�$�ZC������3�-? ����ˇE�&%��2�|�!�G�cFA��oD�VT�	�6�#���Dr�����>���b~P�L�T����E�
�	<��M��n̢䊼*��W;���g"�N�T�*IRaO��Wq���P�A�B�������A�F�%Ե�ς[)��pw�V%���v��+y��X��g57�2+��@����+,^{��B���k���ߟǊ �	���
�ޛ��G��[�8T�;]ǨQ�ug5G�N���]%N���}y|vC�U`�Ƞ�[����|��z<�y��o7��?��Ú�V'�E�y�}ƥX��n0q�;�mx�Ђ�@~�|�u��*�9�Ff�(Uy�`Ȝ�6\w����5쨾1���r�lGLk XC#�g�-���B,�;�b�h��/ԫ�qR���|�$�TgFc�)�w=A�0��>/OQ*F���c�p:�(:#�n��Ç�u^�	|��τ��ݮa��b��	u�u�z�{����ON�"_.��N�ψi�&���;Ɍ�W�ߖ�/��I,���/�F�|Ox܌�fX�~y�Տ�wRaE��-'nD��3�N�fq��<!v���̞���ȧ|b���(j�ͧ�v;Y�6����C!e�m���С�~�;��|�+��
|����b.u�YZ����c�d��3V�Z3a�-|i�S���GWD\;x�ٖ}��͸�4Ryq�Jػ<0:�P�˞��o[���iy�#r��y�H��/O�6��%4S�:ѡ�'h��iF�3��0n�>��)}q����v82J-�b[ݒ�#�����*/c8����³��1�[*��T��ΜfP��!�b��i��kx��:���${7�}�����]��n��"w�+ڕwG����辴\�r�����g���������͗��U̇>�Z�_[qS�+F�`�4����/%��Ɏy��V��Ǭ[�C���RWI��wA�Oo^�W����j}�sc�x�i�J�of���nQ�zsn�Y��t�HF�F�Y�e�r�]mȌ��;��q��V���®�<�'��#r�%ɂ�J��[�Cڙ�+�8uv(�z����{��"�ua���0#�s�n�|*�7�g�T�46�f��ZپR�/�Y���F�]����ԶÜ�|pQaoX�G�S#(�Y����%����Ot�B�6�5;���h�Ӳ��徫Z�6̚�Kr��rur�[M��Z�*�K�Z3d��kP��eA��,/r�D˪
��̋��ZK����s���a�kAԦ��Ӧ|�<&�0ª����͌|�0�Y�ΗIPӚ�E7-Ĭǉ�s��1�����(l"ւ{�<qtՌ�w�cUa��m
V���+�]�93�����l���m�'o.Dȭ�˫"f�ku+���6�O����澍=[M����۹Bei�OtVN�b��6��,�h(/�u�o<��Vv�Q~�ͷ���V[�^Z:�P��S-�eFQb%�!m
5T��>��{V/I�����k��Y`��e�H�+����\�m9G'|�#	뻒.�\�^1��s2
虪��u��V�	3U`�t�ū���%[��P��7z�&�+Z����R��ʤ��7��ؒ��4,Ĝ��
��f58GX5�JT!W\רpzof��Wڢd����f�vw3ve�*����}y���\p)Q,�T�I 5���Ǽp�Z��G��P���g)Un_#p�L}r�I^@Mdy���)j���g���j�4�_C��
�N�/8�o�\�!`�*L�0#`��ƽPw��kb�7Gk1-�jg��v����э���Y�<M��]�4�f�q1Z��=]on;\�U�K�s�N��t���bf3Z�F��KZ��{��e�y0��X$��fb�b�U�uϼ�SN�K��ؖW[k5et8��>��mE��Xٳ���0�]]�*�{/S5r�'u��t�l��/]�������i푴T����;������!��׷��n*�g1���OBx�jU��m/C�l�7z�A���Џ5w�.���ŗ��1�ڝ�j����4;��|1A���
���n�E>zi��'imf���wu�%1�8�z�Xr�N�찶l��:7�Q�h\vQ�}}}s�?��j*(���h��n���O��z���<x��ׯ{�ߺ��W69D�߻�����<v��Ǐ�z$�ص��nU���rו��I�A��8�<v��Ǐ�zH��حE(���D�%
z��8�Ǐ�x��ǯ^��FC�$ss��m�h׻�}W�����t��o(�<�u��u\��������I],[��F�7K�z����{�m��s]-���Rk�ۖ�{���I�U��<����<�k��Z�۞�W8si�E��z�C��D2,� #��`%Q���Gs6��Dk4Uf�u]�9ۃn��"`녥��<ڙ1먶��$�K��|�"ۻ�������y��7���x�NPOʐ��Xi@D.�[�e}p~�#��ǘ.�)�h��.��:��Eѵ�v;s�b��;�FC�"���&" ?�$�,.}<���S�签�̔�Ŭ��n�DwZ�.���{)M2�b�b���@��L��
���P����}u��L�O��<��eo;_m�F�s�tAd^�DIu��O"�F�[_�rxy��#'!��@.-�ږ��"�&jj{c)I���0q��9s�a�{%�N�*I��a1V9�Q�����/O������\Mn��8������	Dsl=�p\O5�]��`G2/��9%<�e��5J��yY�\s{��(�U�e�� _Z�����OD����^D.x�~��ϓ:��x�Q�N��³�����
Lb��x���_Z�5���$fj��.����|d��]s���~)�7������@q��Qq4�W�eл�5�3�H��S�E�d�??�&p�I��4
���igOt�!|��+X8����V��߮z���`��נh���D��?��/v��%yln����X������,�ܕ6B�]L���R���,�\m��_L]N�j#��Tk��n��s�[�9��Y��v����F���to�RwiYr�a�&�8r(��z���;[�~�jS��œ~�!������1�|�ə�|�~y�M���vO2qP�ΐ18�"��0��6��-����� @��K­�͛9W6U>��'�(g��� <A�� �VHl{�23��%���6�a�A��RN�Y� ;x�6��L��"�
�K�XTa�5�Mw�Z�/כ��y}[�[�y�p�D�ǖJ���ܫ�뼩���#i;!NZ����y_��6�q�[xC���M��EE4y\�6Y��X{����CK-��2�)��l�Ϩ��4Ɂ~�@
�jEQv�hW������Pru�#1�F��ըƒ5��v8�y�7��Ђ��0D�5�z\���b��Eվן���T����Naj�Y`*�i 53��ơ|��r�m�M$� �KF�Th(o)�!�~P]���3�����c����t��8����n\:Ǘ�~�5������W<މm9.'�XB������)M�7@,��s�y��պy䋈��%p��(3�Yz���	�4���/)���#=ь�_e �1���f:1�v�ۦ܊�OZ�^���b�E��p��ۆ����R	�q-k�͈�M�~7n�?�u���T�Ϭ_L�
�I19�T���}��}w��xq�%�$!���2=*�ij6�n���ᒻia��=6a�o�L�N�-ب��.��)�p�I
���%"PD�p���Z5z�5���f���c��}h�-��+�ն��_�6�E6��9K���������W*�@�iQ`|����~�^���̉�X-�SOyW�F�ݢ�;�wD����/`�5�ʡ��<;����wf�7H�	��F���c����|*���22l��U�2<9�ʺ�/��<m, �<�3N��~�lZ�]u��K�+�3��heH�^~�.�j�.��ς��֪K2G+��{�Dl�����7\1��Uu�4�<��o�������M7��|�Ec��Ml��x�K��ѕ\zc*z��@J�ØOE�~"(宱 ��-qZ���ފ/3mn�
ۻ7]��a�{q;_<�2��]���\�������{jh��F��;�@�m-,ٳ����f�x΁e�v�hd����i׊xn����(E�>��j��G�k�����5[���w�%� |uC�e����N䞥Ob�HA>^~��{j鋇�k�<b:ffQ�2K�ox
}Gp;�`�B,��	qި�3�Ʌ�fG5���l0m��͜a"�*�ô��2@ď��u������u�K茢�إ�o�;.�N�*!T���T��o\T8]��5���)�^�v�f��܆涙�)�᳹qs�T��X%�ǟ+���JsY��1�B���H��O��G�̭fo3/�%?�co9�ﳷl�:� ��࠴È����W�|��%5ޙ	��"y02�R=A�n9�^�¨�Y���T�n/�D�a��*7��F�Dx*|C@���'�y�:�e�z-�Ylӝ��y�L1�{�R���֦r�On�!Ŵ'E�O|��`�k�m�ɉ��K��wy��(���ޗ��=��-�y%I�>��os%���Ba�����A̋�t�g�/���d�Ӯ�LQt�ѩE�y�)�yi��r��k�w������Y�iJ}��9��I8�kt_�Օ"U_Qw�7i���q�OͅAi+���PN%����=�Ҧ�����K^�8pw���Z�Cc=��vt��cu�4�k�Ð�9��U�nwX����2NB9�a���(�vn��;�!Ъ�H��`���@�  A/5�lT]�@g���KzV�����ˇ��.�_16���Azzd&���g`0b9Đ�^a�oК�٦�k��ףU���7D�5�����4��z-�Q�>nF���(ɬ���&?��Zr�����~���x��ZZv��Otu����r�pMQru�.�b�q�T�F�����_���_ygL���t�˝�T�߹1;��0Ӛ��3E�|O�I"�ٞ>0޷��v���5��ݹ�}H4F����O�[���7��ymS���=���a]Q^�up?����ш�1���Ͼg�|����L�緿��֛��P���^}��~�v1o�k���aziw�M�9CB&�۩~m5�ru�(��^�}�C��揎���1U6�)�^E�'���J�����/dC�!Л�ܺ�l\�7��=qF�׳e0�nA�y�O� .F5pz�3�f{6k��o���YZ/��)��_.Z���*; �T���Eww�%��G�.����f���9P�et����08�a{.=2��q����|R�w�np���=��]����52����z1��7+�L@W�$��"5���Yb�y
���ý!��Nf�r���}���1�&%�=��4���ЧQ����l����H1�<'-7���J�%�����`��3���ܵ���.��H�-�	Ml�p0��d���u����f���1��d"���O�5��{<�'z�$���~�F�t���9��as���6���y1�^u1���B��r �W��l��	�L;e�5���19�O#���ʑ�.�&��0ܷ����v�VwGc�v�h���V���J�p�c���(��{\��h�\�L�u�����Y��?�n�#H��iSV�Q06sR����2�ר�}�*"���ec�]B&4�6�F!RX�9���Iz���ߏ��y��o7�*s	BBv]�4������Q����˞�Ķ��U��\�[+�&([FL�콫~�" i�[�S�|w���葏�� e�.X:������M_P�C���=���K���	���设v�p��8��O���Պ[����mt[��v����C�y�kt\��|�\�ӒpV��Ҵ��xb��������-���lz��}Ȣ��#��:3YŖ�-��j�Ά�^]�?;k;Sw:�`f^�O���K��;8�6��rŨ0x@'�x?���+��OJ�XXA�"o+��1�����>ͫ弑Ӡr��ۡe���q�Y����p��{gɿH�yA�6�~k���I����N*&v	���ʿQd���5Z����;gb�;q���O��Yw���U�`�0z��
�yAr����:��Eҹ�Y92�f �8�|X�������V+�Ξu���
ä�v���&��1���~q�A��چ����l/����ӌ��y�T[����`�����c��ƨ����>�M!�q���u��.���Ǘ|�7{��#Xk�ȳ/ޠ�Y�p*��͘�`��sX������8�uR�N���c[��8���_r������i5YUlӒ#�M�.U��Tsjk%L��7K���oN}��(3a0 
�"@�B!MJ�������|�5]6<N��f�	VP�fww��>V\}��1klkȄ��t&5劅+
��SQ׹Ɓ�/;�y�
Ķ��6�M�g����ѐ-L q��-��!1/��O�J�Q8����mq{���켬��QW�\��oF4_����zC�qu.3��;�/��3eJc�`_���dTt	�N�~��'4Ge�� K�#B��|�%V�}�|?+:���Õ��Vt�\΂��C�՚�':�vI�^��]s8M�Z^kͧb��������0ƭL!�����t؛�E�c��*��]%�P���\­A��(�NX�3d�B�e(��!~ϖ�`�➙E�×�փ��g�����9�N8�Ҩ��Zot���	?)�-/�Q*�?�Am���V���,T|�.�p-hA��pchLn�2)W�����ҵ�%�����\�R�2�����lL֣�D8�`��,���O\~�? ~K�s�M>�J�_���=��`?�3:	u��4 ����P�����J��1���3�A<1�������4Oܨ�S~�FI�Ƙ]�ay�/kUq��J�F177+���vBu�7-ΛE�/}-0�K�}��hJT�hM�9n(&6,Ku�ʠ�9WU�"O;ǆ.�)�lWbGk|J;��M�4>���kV�pP�֎�p���y�Ȯ�t51�ǁ�+4s4�{�����w������^�;�e�۰���x��H<"ڨv�F4�з�z8K�{aQQl��B9�E�Ο�� Hv���x���/D8�*ݫC���)�\�i�`JV`Jd<H�8�Y��oY�Q}����5m^��)�nBN��CQ5��u^��1�5B������/��0�Ӭ}�����
&��q
�|�ؔ
m�����2u��Ŵy���L����Uzz�_V#i�{�k�e�	�-���y�o4צdV*�L�a�=���ݮ�q���~uf(m�05
5������)�aH�16��i%�ϘPv��]���G�u���w��/�7����U|���k�:y��!��d^��No�<�Ee^t�E��d�<�:����7�wp�I�j�eA%I�k�8ˆ͕)����&���a�ݒwn��dɼ�2���3dl�Ψw��]0��J.�7E2oPZdp�8噃kϝݢT��Pa�b��\fá~g��Lc"�D����;$�������{�zK��%�'g���8��X��G�sђQ��n�d�Iax2������4}.�t���w��FC|���5�g���u�=m\(�S��[^�Y+A��׮����ى�A���@M^em����;�ܖ%-��֎��5���;���?������yy���b�jH!�a��G�`嵦4F��xN��5%�5g%B�Ra�Ǡ�\ؒ�F���a����ES����[KJ@f ��=#����j�� ���cv���H���a�oel��f-Ӌ϶�����1� ���#oHa|9������H��Φ|�t�>3�<֋����u���4s�=�G��c�	�ۑ^��^��p�σA��������]ҷ6c'�$�6����";{��٭ݙF� ��z˖�C�V ��$��(Aڕ4[��^���H~`���C��tFki���0U�ǹ|b�f�[�j͂^���E��_?����.`\��S�|9�O_?�_��|<�g�B�ߕ�q?e�}�0�ۭ���%�q"��BW��-�ҙ�N#����닫y����<�Ϧ�ϓ�\X{�Na���Tz*޽�*v424�Һa5*��Jݼ��{U0�^����ͼ��P��"å��s��b.=3��zq�62}�cq^�BvsϽw���Х���0�dIz	t�
���v"qW����~����L�H{�Y���i��4Q��I�{�6l���4g����g��x�7��Ff�j��L�f�V����n��o��R*�m57�-0oЋ3��>�~$�wmu_S�D=�9�\{p�o�˴<��zU��֞@�!U�:��U"��Y�s
�d:�˙�\��y�&���4�SM�@��� ��=̅��B�1���\GⳢYA0Q,�ThR~���s׭�=[�H-���I5:�*�['@�O��jB!0�q���8���L�و��eH�@W�4����G����F{[�ȿ*���Y%k����9��t?��T���^�w7��O�9��X�E),9��*[5�^��8{_�҉t�x [@Ǡ9�h	�v`�'H�y�R�m̋����6�Us@eq�nG���͞�Z�
e6���Hİ�0�4[A�'#�H��^��D���P���*iuu��(�W��i�1��<a����JN3����S;�{U�C���`2���7���Xڊ5� ��F�ޜQ��>gUĩW��F�w�]l���X0�R�;�u�0���R�4�Y��z�n7ge�V����Ux�v�l�����uL�i0�PoK�u��2/W��/U@�G�&�����\S_�׊����L��׺��kښ�ݯ$vP�CX�L�]Q�,����i�����
ފR�'�%}���g���U���^KH�Ǘ&�;b�^��9n�.���Q��l�h�*w��э]L��#�4Q�2(aګ�']�V�|�ǂ�:��%wE=�K]�]��~�g(���-2o;��t�JP���3c'�@b\q���xy^2-�hH��x�+�3iڛ�%���d�`w3G���/6[կSzL�.��0���p�_'pQ�#��qj7�$�4R�s�vqT����T�<��֦n�c��A��Svs�˽�ă:��j��{�\��%���K�p�!N�Ujk�go�<����oad�=w��>�/�ʔ^���j��ݽ8SЩT�ъή���Ve�3o2���uk�5mv�D]�T�u����NV��Kj�IR�5F��&J�[H��n�*C���9�g�Yu��1t�%eQË�gB�#m�;��Ɓ�Z��'�xY�{F�ʼuR�K���g�)���[q��ۑR���S�;3:����w�b�7�f������ͣ�N�RΚ�H<����Ў�"ك��)K��}��u�:_+�"�|U�M���=A�>!��U���F���z"�/�M���%�/�b�|�ʡ0$���A�M{7T��U��j˶�$�=��:����C9j���L0e)�I5:�%CNt::�k3�d����4n�N�JB�`�E/D�kX��D�P�UqUJ�5��!Cs+����gah��Z�*�\��VE^&�@\jS��I9R�ʈzь
�[���rJ����n��H��J�WAV�ȳ�j�\q�n�㗃ꗼ6Y檱�9���eqS&���"��^[̼���aU!��ӨDl�����jR�f�Z���]0`��u��O+b�\��!��8�ͥE �2��Ø$��@�f�=g�/�J\M�%�Y����ʳ�)
e3��h7ul���������1ں�\yS��Hb����,\f�ڧyCz�%Z'ӈ^h��wP}�@Õ�|Gn��:��,�Q�	�����G"2���Nu���u ��E��r29=�k��aS�¥�T�;1��/�!�$�_��6w*]	L��ٝ0�P_et|��2��x������룦���:Ğ�.a�1��\qK��������Ԋ�)����˷U�88N�rG�J�5�T��3�]-i���u=�i��{�»���8���{�q�����d3:��&
�������63D�S������N�ʻ�ҩz�;��A��϶�m��Z�l3�e*�-�L�-�Q��3��<���2�̸M�;/�vj+��!XyٚL��ï��8۴b�wK�.�tin
��Ry4�f��s�*��iq]Ϥ{���&ڤ�K��A��e�eBZ����2�%����K�EA���)F��#EĠQ��$KL��d9O�8bd��E!��!�f&�&�T@��`��,!9	��"I �^�aF���єY>��[V
it yH%���y�������͹\�D�O��}q�Ǐ?<x����$��/��o�����P�mN�eT�c�����x��ǯ<�{�~~~��Qh�.�HJ��$��I#z��qǏ<z��Ǐ\쑑!$!	!	�(��D~wy�!��Es����I$��Hƞ�ێ8�Ǐ;z�}���?X�m~����cK�%���'[�Kk�]��G��_&�|_���Iݮ$V!�!�4�`Kwt+��D$����$E7�Aݺ@�Ɲ�9�Y
]�����
�R^Wۘ��]��ur�>}}��u��(�$`�6�������;���� Gl��V�����O8[�:��˭t-��s��R�ֹ�(���/�5u��b��{�ƞN'd������P$��UUwmy^xY_`$~4�MSMSM%6���P���0�[=�37��},ld �>|���摡|}|< ��T���ܾCwn�U��n��ֿr�\��F���:�p=�Uq6[$ʶ�䦹�.j�n��뜫�@n �+"B\"���WޅF��[�	�����{QY�d�E'�����\nr��{-��'�ߏ|:����7�T�=�3��[�J�祈�9>���O�Tf6�5~��U�;�g�P;x2�e������o{�T�^9�g5'7~����ī�[��xJ�KZ���Y�6fK��}��6��_eH9o��B��2@T�D�U{��+��Ӱ���%��g���x�_&�N��$	�:��N�n����C��e�*�o�%��u����y\Lr���čt�6��g��1�]q��wP�i������t���c�a=@l�����t� S��\�EW�3��@mkfg��>d>��t��.૝+�o�[}ԑ�����7�����R�nc��Z���5QMu7�vs�ɡ�`MǊ����I��Jc4	!1�SN�aͬ���i)�&��7F�v{�J��,��n�J�ξ'�:C�K۵W+=P�]��3=�}����KM4�L~f��ɾ�Pk��*�]�w����h*�W�:Z�fnycd=N���S`�0�;�����\�fff�:qY�R���/M���� �l>j���U��}HK��V8U�Wkf�]�zl\�,���nA�㻞��Wn�����㫧ƃ�g`˩�-���r�j��Q�������6
E�����{Z�Ύ�p�h��xUS\or^�:3�,\�^�������.	$?��6�M��yz�k@Ǻ�S>LW�zߟ�.�@$@�%��}�R���Z1��.�ۥ�ۉ�oSY`�
ɾm�2��N�N��0%h[>�'2�?DΌN7;H��2OcK���z����r�w���E>��g�S���論�>-���U�R^�ͽQ�y�w1`�Ầy~��cD��qc}v
�u"���q�rǉ�$Rǆ��~��Lv�ϲ����ƼR�]����"�zč�ge��):Z�[+w�k��<���Ε���[����̺+J�T�}����6�*V_V�BkGOf�S=cWFkiM�or+��$�T=��Dm���cn�f&��$�E?���1�g{�����Y�<�׻h���~����`]z��l�:=r90E�p�+ar�s}�6'+oV�����	�L�l�*�)2I*�}���N�����f�K�F�?����Gs�����M���QH�BW+�A�v���+���d�B=��:sIn�~XXE��)��ؑ�GQD�����}mu��M���[����M��\�7מ8ú���S�z����I��tV<K��c>�vF�s3�R��Q�q�ζ����.�|W�y�gOT�c�bK����U����/q&怛s1w�)>�8�4�L���SVzg^m21�g���j��'���7[�l�9=��:��~�`D��3�x��朝6�$@/t�k��k�a���W�W7������L��ޔ���^7K��^^?cv�����m\?�*��TF�Fi;ŧ�t����a*лd6Ke�d	|j���|	��)�̇�DeZ�
�d�����r-��Y�j�,M��j�}:�s��1��=y{	K�8���)��g��}2�a��B=���R8��3iu�{�ɠ}�<���>�';q4Ow/%e�����c��}�}=�o5���{��Q�Bc%\H�2��d�9�T��|��W�:Dm�z��]^Oy�C��A���"��$��gSg=m���(���ٽ/�/EY1������gbU��O�mM�(��P7�'ȳ�pW�����'_�;uk�����U�AJ���ǳ9k8m��.QB6�VE��I<�3Ʋ��<E+ڞ�j�JR����^�uz�[�f��A	ܧ0�����X�軏35���x@��ˏk?.*k�$U7PxĘ�g]gu�f�n�����|>�����o�N���m�IKs��G:�^mdK�C&�ߔ�;H��C1��*���6�0jx0jg�ZI��x'�o�U�?���@�:J,��9^n�XK�qw�~�O^���&q;d,�j�/w�Gv���H�]�m��騅���zu�v�=�`�=#_E;�C���o7�����bOu���U\�vN�u��%���uou'ě=w���͉6zî�*��? ��v,�?���[���ve�X��(�+m�t'7���(=��Ҭ����ow��,.A�f��v�w7�}��d��Q�$�QW+�5\O�c�6�w�xg�w�}��#U��s��꡼����%*��fl�m�0#{H��L�3�m��/x���5�≘ˁ\�J��V�v����ð�Oh[[#�7~��Z�>���n�4q��a�z�ޯl��g"�v�v�����=��zj�p��v��<��d2��K��?�pk�V`̮��Pޢ<<	�j�;U�a������w���%l�X�g#���>�,�׉`��x���S���j��ף��3�/o�� iր9e��E��I�GCzv]	}����c̪�!��z����VF����R��O���>����I�6��D��%Ň����/��w��F�M��{O\TK��]3yWR�כz��[3��:*�p�oC:oGR5����{8���	F��c�C���M�p����[��-�RW"za©L[���pǸsNhKcJ�0���>�{=\���4�4RJ<�er@����[]�W)B�ywN<�1G0P�eF�{���S�ի:y��9h����Hh���cZ�q�M,��a�Qe��OMp�j�mu���T:�nIY�S,�||�o7���v���w��1�
w,&`Ш�ċ|J�!@��"�-�r�[àn��e�:3c�?l�X�L7���I!���}̰��[O>��{kr�ُ3�E�[�T�;u���u��)�$t�r}��{(��ԗv��OB�w��i���c5��8��F���W� %K?c]*����ڻ��� �y�],ڈFD���4�o.K;���oh,�v*i�Q��}�����_1��q C��2��?�z:��ՔOt�Ѫ�r�-D�ٮU5X'��+QT�������|�������(p�{�z���.��ת�¢������n/{H�D�c~�-�᜴��x��
4����ԪNwOt�˛ԹJ�-^�/�#�M��C?����"T3V4E�P�޷���) �ʱ�y����H��Ǜ�Q�/�p��51}��)�/ܛ�Q\�"�;MRi��	ʱ�z��5�i,��$�a�5��
�(���h�[6fҭ�[T�7(B6��,���QW�H�����|�K��Dj�����'���^�h���ߒ�y�����OX�1�s������̔$W@Y�蚖�]��=�WO���ƃ��{u��l������9Шm�h���P�e������k�.n��㫋@|��\���o���z�&^�
�}�j�}����\�o�ŵ�R%�K<��׎�ɭ�v�JzMA�;Uu4�E[?�6�#�b	��<5sj��>���3�[ׅ.) Fo� U���48�����SeV�(��i���2��ܖSu�k�����zr��m�
���F�����]9��<����x5\�t��<�	04�4�&�=G��I�܏n�\3	K$Y�z�)�6��0Gl�9q��zG&��oJĀ(���V�+�3�;/\E�6o�@t08p�w*c�go8dn��m�ڼ���i��޹�����d����^�_ox���1���ﾩ>�p���jV�.���}XmS:�V��Se�7��+	;E�{��䧵A:�
̼h�UY�0 ^���*�K��g6�3�>�Ñ)�Wȭw��F��0A^��A�E�վ9�֩��][�Ps]��h�����+^f���(;���7����y��f�~������һ��(��W�Ń�3NP�]=���G5e�g��+�k���9_�Y��S^��b��{�� ġ�޷�~���w,��,���.� ��AxC�\�q�P=ތ�z��:9������'�CjG79���F��)5L`J�h�f����/k��Ō{H�~�T���[��iq�TS���^w��|ؒ�rn&:*�B�<�U 0����W:�scv��h�[2���oKX/(j�k��C�vkɬ��S[���W5���	4��v��3qNS(��<���1k���aO9Ggϔ�&�7S���}��o8����Z{2�\�cx���v4�sz����M�R�dΊ��.�i�)(\�����WNX,��K�V��oX�:�ު}P+#�&�D�ׂ��\*�v*�K1K�bXo3���}3�䇺=|&B/O+U�hy9y��l<��w�"�2�힂��A{���7�C�U׊nE����7Ȅh;����P�P�
�:�J2�ku$�*���)�b7�5��`�4��}(�-Ŷ���K|O�BH���>�gv���K��
6)��Bp�#-�RP(H����1�c��d���3�9ϗe�H��}����}� �l��-����{�ޒ��.1z�]�'&���?]��w{�~�t6ӰA��#=���c�gETe�<]�n��F�����5׶�کPK�,Z���!T�r.�/z���&;������vnx�֑��]˱�6�������$;�8�oY鯫Y�u�a�7>����[�H
�zhҏ*�2w}o�=��YD�?lOYgӃ���m�F���ڲ���;99Co2!@NeWwn����+�8n�d0v%¹5թw�6���w�M-m ���˧�m�<�2��lt�P64���r�%J��V��,��w�:�R�T�<T��7s�I�$wJ������`>ca笯��0_4�}`(l��_���JT����{K�[q#uH�ӭ��y��J��z�~�C0a�)0��{��z��U�xֆ��g!��3��,�������k����WjȂ�}�\}ܓ���q�t0^�^\&�!!�!<���8��6���}r�l�ܴ�d[�$c(f��t֣332�]�5x夳H���J7��*�������y��o7�vv;L�9�R��j�++@��+"@K�
�S��Ou9����g�!]�uD	�[���Fr�]:�R2��fz�Ok�#%6���NVɫ��)3�qbzb:<��x�A��y"	��~�_�Իٻ���Q�&r����!}y �<	�~�L$㩿z��)e�r��,o^�^��݇�6u��5;zd��&8���Fϭ�m�H�I\�Q[ñ�ݞ#9��6�2��{�Ǫ�RJۛ�e"FN��9���m�¶D��m��˶{���Xk4<0ka�L� �ɠ��*=K�2<���<��(�k3���K�|�Mm�'8��6*���%�q7Ǟf�3h�d���;Xs���M�i����3��A�ok��fze*@4{���AgrL*���|�\�����.a��`����ߘO���R,ʗ<�JA��'z����揺&�L]n=�����P+nu��+C�f�d�hd��nd�U�)Psk�펗��X�PP�&�]�uN����wba���0��K0M������Z���Q�Xs�m
��lSv���sM�ئ�A<��Y3�)�n��.��:"��V*x��3D�wR�����o�集L�q,я�}�U>_"^������^~���%,�E̻�j��s�:f�+��yqd}�ѹ�q��Q�����U%�QD��#קzA7�t��5�
2꺨t���v���+zB��%��Z�	1��<�E9~�%���6���
�\)���0���C�.s;�U�s��4�䩬嗐6�%�1�:�g!{�C����5f\�h����d�����1����"���H(!�B�r)țX��K9��bVo&^[�ͧc8c����E�L�F�ͼ�'n��+1�]�vqz�k�9X�;KK�A��ڞ��)j�&x�+������I;k�z[������X�K}[���4,������c�t(��K-S<��VS�����f��u_5��*D�:b;�ݛ��f�+y��I���gY�(���;2�U���L��W^h�~�ZfS��ZK�nѪܽ�[ܥj�L\[Kk;n��lY�B���m�G9��2�*��	��S��i}��u�l.Ri]��+__VKn%�j	���� w!Jy�<'����3�$"���w^UA-{�#@bx,j��Kd[���=~�GW4���hma�"�5r�}���g�]��˾�R��\����l��n�ˤ�ك�֛����+���yl�wm>��9'Ǿ�zK�ƶ@�����F�<�T�[�w���.�ǩ�[�uWF�PV*��|8dwQ5ՠ��f�E�3(�,=&�f�����oUKd�Sl��,VT4���J�c9#%�%��˺��r���R�%]Gދ�6ޝ�����,#-�}˩��V2&�0���5�3�\Y�J�oR4�ً����"��ڇ%ħ�f�����X��� �E4�偘	syֺ�x"�i�[q�.ծ�$;9���kk�y[Re�Un��*n�Ɇ��w#3�W
�d�|�Kl]���o�1��0�ڽ��s���|L�j��yM[QJ���T%���sN85��a��w{�'j7��	��d�WZU�Y��p^N��a묎���}4�8��w�Z7��2�2J4��p_f��R�t�g��8�h)~�o
�	ɹ{��A"��//U���P_Y��X.�9�82;��h.e�V*g&�p[���q�ں���o��Op�E=�6ze��M���!�����uL��H��Q�j��MC}xh�̙"U�IWx��h��9-XV�}���IƑ��4��r)˥�nT$$$$!�ۍ�z�Ǐ<w�7���{�}���̌���N�q���.`J��M7��8�Ǐ<z��Ǯ{*���o;wr`/wDf&i� ��BH@�:z���x��Ǐ^o���w����z�s��R&�/��7��|߻�~o�����Ǐ^<x��d!$$��C�D�X�?7�\�{ܔPH3c�:����LTbO�"��^�cs���ĝ6�3f�2l^\���$ڻ�H���o����ė�J�����E{��k�1H�PDd��LQ��K�pb���H&��ݮb%�ٔ�"r�A�,Ħ�5Ο#A��R��*��T���#xZ�_Q��:R�z@e3]m���.}�Qv�[��5��}-ڻޛa����[3ͦ�_u�c�w�������Y�cd�9d�C���c�s��B�a����G?87���h�Z�Q��ر�{�����8h1�:`\ϑ���f��/���P�[�7(�������G��gҫ�uT�ƅ�5���ʹQ��y�]X�l3��)��o�z�x��HY����Z�������!�]�l��>Q<�O0�~�&qg��1G�h�E\���{f�FwV�$gjd4u��b����{~�QO@� ��������bWV78z�އ�Z������6o{o-M�:��΅8�?GJ��q�;1�z���1|;sD^��l�P��	���˨�n¹�rf
�܊�L�ۓ�1���B�с���gB\JGЊ�|Y�:ڧ=o~��G��i�sϕ���c��/�V#V{:L���%�I%>������ކ�w����j��*rC�G7;1���yZH��$aLO�&qujʯwT�t(U��Z��FZ�'�&8���es�Gg2h�Gpk��2���k�ͷL:ii0%J�5�n^AYl:�gQ�nrdlB�sꮾ��/}�����������9�^�w��� ���;g���"�Bг���8v3vs>��9ݯ��&�(9��Lj����Mg�L���r���{��O�;�;ǔ�"�H�HB7��1[��t��{�?#����L�j5�: #���ח�Y������N�08�*g�g�a�n�E8[���RY�V��i���'c+Hz�\J������/-y+po��pGcb�Ue'�9|M�Ą�H5������Ca���9\�x��Hm�g�c:d����1�~8�'3�#��9b�y�}x����]{��\���
8��tϣ���f��#�1�↨�f�bR,[�WV��#�w��Ms��M�#d������+�;����*����uP(����8{�^��ٳ���D�;�l��X�ǹ�K=���	��Hף��% ��q����~�p��{�de��1�Y弑F����mŒ�>�/���C���V�`ۛ<D���$��̐�Fр������f)��C\���&\�gu���-�r�͔�v�أ���U3�e�q�R�>z��9O/����+��3K�%4e6%"¨|�e�U��*��;;�'#�zs3�C�/f��n@26��c��6���l��@�z�7Y)�;�1��V0ȇ����X��r6�Sy�=���)W Gvf�Y�ɹ�3Q�\�F���ٯm7Y���x>�&3�a��~��O$�PS�L��>�;�w+���;"�6㧽K[�p<�^ϡ[�k��zQ��v�`�ʇK.�)��fcw���y	ي >\�}�Pם&�sQ���:L��*eop��J	�[���מ��ˏYo�m�7^�%0��b��8v�Gb"rj��Yz�mՙ�t��c����;*Ic�
�1�#�UTj��eؼT�a���]�i��֑�+�Wc�.�6�T�~;���Ek)w��mu�I!5-��3�2!N��Nxo!^�I�*��m4�;+`)������O�r@���qR#NMħ5ݙ�{�pck�%�T�9Y����_[o����`��̻ъ��n��i���Lv�tDj'3���E�*�,�ewcz]��=���(�ƞ�+լ�V疥Y�0iȳ�b2;��ٹE=ꛙ���[��������"��w�f룝�Ԉ�}������i���4C�T��7�Et�F�^ɳ�/R�c�ncu�O_&ɕ{��L5���Ĉ�����:F�VЫ�G�g�a�������ܴ�÷nI���9�d�j$a�=^�׾}�P�Sǧ�_Hy)1����g8p�eY{DfyG�-D�$Qq�Yk���ha`���hi��Of�9&�:�/E��>�r��Ygfe��arVD%�/)N+tO|T���k�4�\�����5zj�r�dt��Zz�}�I�PY��-��r����k�3E/��ED�jk�ȱ);4R��moObM]�=`ܽ�fY��v�,�����駡4�A��Kϡ(�S�Ƞ��E،�k��:���ź���W<j��
|��P{��N�vd����<�P0�%����T�ܐ��$-��ލ]m���jD�ǫ�M�_�+�����:2�$~�����`݆�Oy��I��ھ��m2\���	�J<3e��.�E�����l-��_j������A�'ǌ�P����^ۄ�0�"
��&���lV�����#�s{ѥ�K$o�a{ef�t�3���0e�ϲ���I;#��w���y��o7�U�a�u�mNF�uu��nx��\lk�+K��g��rz�]����Y@�4��~��z�W�o?�M�yI����;��n�����3���W5_�Ȟl��a�˷����&l�����V���p�̭�SV��]�ft�zԡ�-��!��0���R,ʐ��z��5L95��j�={pl�`f��>;�Jh];#��|�9���(UL��at"��f���W�j���Uyi���>:�1����;���E�=L�Lݖ�9�O��0@l�Vw.0w�N������m�G��Ug��;�t���b�ؖ�[����WO�Q$Oh8*��z�o&���6����`ןZ���DԚ���މfW3��-tڣ:z����Q�}@��l �$�E&
c2K���%�-%q��[���2��P\^y�;�m�o{��W`���㾬���r�{���S���̏k�9���}E��+�eu�#�Ё���y���n�l����T��6�.
Lx����N��X+�+M���'�6z���(�R�kǌ��Lh������o7��v���f{ B;��Ɵ^S���U��l�A*tr��1H�a,˵� ����3���x*�$�S���ۺ�s4�7Y6)=�D�U�X���*q�u0ư�~��ԴEvc)f/�Е� �-u[�n�U�Q2Σ���\=vm4w�Z/���'��M�AU�I$����7���[۹O{yb�k��|��VHФQ�����)Z4���*�KCd�5R�Р��Ǧn,�f>o�ނ,�ճ}Erh����]�:mn�ڪ�Ϲ�q)o+����:�j�,�Tp� f�C)���F6�������z�k��	;�C�ti;�q8U3�q�-�w�����h�KN�D���̪){�)����䶄���M8b�m-��ҳ������InqԵ��9<4>8��7���5�TN�^+�7�y}x��k�s����t��������j����qS�;�3�1xh�UhJ}�ͤ��0��w�Jk_nd4�/=����Ӯ�U\ē���knd}C��,t�X�7z˗�+r���7{AԻ���f�0�i�,k�1�a����vbR��G�R8�Z��*U7wuE�]�eu)��1�y���	��'	�;��� �S8��~倊�q�W�~�)l8�<;��^R�;��*�8�gr�`&�Z�.1��\O����jr���b�'��c�p�K#&�qۃXB��U`I�O4�s�5��e���ϙ�ٸ��q��/�<�Y޲w�qX6[<��5Q1Q[��V�ێ���ק$�q�.)t���W���m,��y�z��6�4�ݢn�of\=�ϯ��q*duϸ�˞A]{J
B��'qQ�ˉrۃ���NN����w�@���C�#Ϙ�>��V�p�΂y%)GEC�jo3����{}Zb׫�][��[<�T�����d�V�r0M�S�Y�4����{�َ�U�U�����+ɺ��9�4�l�vy���@H��l=]�X)T��1�_vz�noc@��]^=�f=��_���'�k:#�)m�E9�)3����;���gK<�!Zk��=~J��]��VZ=#��u�S+c1��b��p�Q�{~�(�M�[�_HnZ�9mfn�I�m<�S�N�7O�{j���]x2\���dW/���N��}�{rp�?�����}~��e��v]˰A�r�	���~���}�����-�a�Y���ϲ�:7m��"�øl��Q��k��(�]�c�imwc]�=2i�JdoDwf:aF�P�� EN{]��<7��{�;� �fRe/s44]}ۺ���ED�pR�ۊR��N�ڲ�=�p�r"�kx�L��<����,=$���|�!q�I�^Ѹ�kVs�S8x����STgs�#̲A]L��6?�}�g��u��>J���g6>����N��;:(�U��吅���:?O��0f�3h\W[��	r��l����W����U�9(��1>�����@Ӎ�<��5ᙙɆ�ٹ���4�Ќ�oI�Q���^ر7SSF����wԖH��E\��yy��7\6Mv�m\�a��6ŎP�I�ёt�T��ut���,���L�UQ�ߗQj]���*�̂�LB�Ԉߝ���I�k~���Vv��&��-f�#3����Q]U�s��c�]������h7uϻ|�İ�5��uȦ�u�J�̶E!{M�=sk`ǝ�\��K;>���#��8����y��o7�
=�Zz��:Ӕ�Q/�1<h�̟�M�|}��ؠ�d��,v��?uz+ {�ɿL��|���&�����	W��0"n�{�z3Xz`��Y]no3�B%�q�|��N�ݙ-�W�4��Dn��F�1C�b�xM�f�F�o惩-���U9̺G5VST�p��uܒg�_�iy�|S��ѷ<��R���-/^����ؚ���G�ye��m��8�3������Q���p��;}eG����_p�cH�wh{�����]K���K0c���t��������=�,��l�c�B���Yw��n`^dԑ��&�3���w����Vap`ͥؽ֗��k�o;�^�I��]�z{[�3�9���v�����eI����&���ժ��~M"��W��ޗ���ǻ	�AyԂ8&���{|U[~I,��b�R�⾂��3�*)��C�6�L�p����b�e5��^�Jw��_G�y�t�!B#�\�>��P@"�d�5���|��*Y�z�L�[��I�y��w�,ذ2��ۨ����v�*��6�{�wut�0���y��`��9��b��.�j��BqCzL��u�㞁�'���0�|BCwe�4���Rj=OO�x�U���oF�]<z�zB�"x�i��0��*�n.ޡ�����(3<<a�6��6��`=�Ҩ�����&6��~��������_-}&mX>���/,Ϻ)�l3�� �=ܚ�~��Q{��ܽ3;��73ů5Z�)WwL��1��6���0c�3�T>�x+��휺�7�p�g���]���wm0m$�����ޓ�bni����O���#�d����8��m<���$vp�g`c��iЕ%*��|��m2�)���:^�3ߎ�`���'չ�9�����ށJQ6���b�$��D<3��$ba�q�؝���&���!�ϳ�@댆��A��W��;������E,9ۈ�p�ξ��n��{:�����N] ;��#V�9������.��*�"/�>ٹ���E�*�F��3��X�X�X���ܤU]�i2�j�)UI��:������U���A���U��%�0b\31XѺ0D%i5���]T|�x8�:�R]��W�
�����u�m����x�d�[��c�k���u��.�p�n��V�)�z�a�F;��8Y��9ᬦ�˶�
� ���=��u�Xf��Ɂ���	�m)�뙪�ԭ[�[s.t�&�ʄ�\j�ض�d����:i�S�2%������K;��Ŕ����<���Ow:���1�EL�.>�����b��t���[
f#pJ�`�\��u���|��<4��R,Oά����l��b�ɮI�b������Nl=jɬݔ��%���t�%.�i�&�(�єmಆ�"��t0���.�H�=�u̹}{ym�.Itd�{���W#7�UB�|�EI
C7�@�{1o�3��e�4�����܇�E(�̹؍�h�%X���s�Nr�'*�Hxd|H�dޖEm6ޑ�&E`��Nm;�"t^��k&H�"��xV�wgT�u<��'{%vN���D\a��OR8q+�.���pt�@��Sn���k�6�i ~��ns�+U�����lENYBs�b�o+is/��uof;��TdS�y�}�8����Z����&���Q$�oPǜ5V�I����5,I*G�ꭃ
�(�P���F��``"�IR�i�^�e����)�T�eQH��S�8(��lUX��}-�\�(�5u/ɩ��Mw�4=�7�w��/7ԣ
�Ce�J�Z��ղڍ��koH��$J��b�ϭ9��h�*'�;��b)����j6�/���܄�;y����{�$�e�(�kU��{�k�o4��Jǒ�\e��OH\��xm`�,>4L�vd�s��G�vL���UkkYn��X�gsUEt��Q�����j	,>����O{�vK��n��WəN����*���|�8�mI��~�9����٢�SQ�S���#U����WaMm啼�\��K��6���U�7���C�������3,ԚE��X�ȓ.��J��#u�k���#9na.�jEFԾ���Y�	�y Jc0�{��3�'{�����ƍ�M�Dj P��x��gu]9��<��]Y���CDw{��O;o֕1'W�E�*��^j��l�}��Lb�J�k�Oj�	�����c!gI)�DA6�{��I��\�o�Xl�Pv���.���r*PՕ!{���&����&f�w���0#qb<���v]���+oE=����x%8gS��'>ֶѳa�A�US];b�}����]�2��ⷩ�2_�U��\���N���Q�����F^��/xO��!C�v�Bc �rr�D���&�q"b	B��H	�&���inQ�U"�_��N�f��q;>I��,$R��5(�� �U��۽����S�A\B%m�C��r�Z�b������&�Z+3���n�&`/�ۓsvA0����>?;v�۷������:BD)-��QBQ9�P����o���o���w�nݻ}z�ǯCs��P�IJ�*t*$�BM)$Rm$�!!! �H�T���޽}q۷nݻz���:�v�D�jNUFBcE&MPX�R%��d�c7�������nݻv�뷯\�$�����v��~8Ɛ�����ysXĠW�d�\�z�gӃ��
���W(�dI���f��$�1�/>/^tY�u�v(6����]I��4$���c1Xc4�E!A��Hѯw���^�2#%wt>v�h�=�W��K}5��bQ�H&
!i$H�&���fM&S?W[�ܮk���2����7�\��H�� �| >���>M�'�j	]����.>�����yS��34�w�-wmqZ��}rv̕jc�Ժ��d&��]��G�����VflV���H����!/ �R7�M!w�x����~?FJ�޾�����BPT�iD����եZ$�\_����γ��0[�k1XN��S*ab,��&,�rK�L�)�y�>'vA��T;;��{���}�ն��U
JAh֦�E�q�ن ܈��3�{y-������ޅR2z���-�#x��]^n�Hv|�y9�ЌdN0�N2��eK�e�Y^�3�O���53�\٦u���v$���z�o�h-B�>�А�*����'��ͷ\������t���8�JRD���3ҵ�1�<,4v0F��/�����ze�kuT�OlFci���e�n6]��D�?�*䩘���v0�ogv��ʌ�Hdi��W_�ղ�k5� ���?+���m	�O�^�����s;7>a���*�4����ƒ�䎶m*�[��#ϥ��3�ݳƌ�
!y�d���|�^:��A*}N�s2�.(FM,��ۡ�76+��C��HCO<����uNt�{+���Qt}r�GL�������*���;�*���;e��"�|�-�e�w�bj�btpZ.���_��v��9�%.r��Ӯ�-=L���΅� c�����q~^o7��<�oc�7�+�՟t�:�>U����[�~՛$�JU]�U�s�u�0xmM�[W#��M[@R�ԈF��9d� �£Z������ow��2{���uTQUA�����@=��P��!���/o�3�[�'�s.�oh���׫��F�����A[�[{����o!�9GzF�}�ɩ֊��7���f O�5�;%w7
�h~GZC�	=m���{��#����F��կ#��4
��'��]��붅�Odm�2�Cjܖfwv�eD�0�[f�-���5Cy%{�<#�f�f�/Z,�A�-z��o��F�����q���z�F�����n�f`�[�*�xq�Ƚ9͵Ht��Y;A�k�4[2�=�.`��f
7zC�ط�����]��͌�K�o�q�:z�g'���
�
�k���շ��I1�ظM�G^V�P�z�.���.al�m&076�Őv֞�留Z3�<����^b��\%�%(\b[����.7��d2̮�_��eS��k�se��Q�u:���v؅��z(/q\<��mH���wa��$T_�W���s~�L%x�c�1��y����پ�0c�Q�s�ͦIum7E��D�@��Kd�l�����7e;h�l3��F^kZz�19��H����Ro1WE�Rӕ2tl�ڥ�����8���C�W2*�+Gkr���dn.���xi�d�9Oo�E(��:��AP��Q�a2.�o�m�jD<��*f�dE*UIw�[9�AR�ճ��m|*%��dб� *Fo:��j����ǎ���4��&�3��ް�މ{��< }̝]ƫM������<��6�[��'�r�gK�JLq��X7-�fd�ѓs5��U�޽A�iK�Gu���/y	p�R֎^H�l�.@p����g.z!vb�
�d�#a�g'W[ͷ�x��׿%K��������]����:�=�CI
�.�]�l���}����96o��;�����6Uxu'z���a�s�8h�'�]kh��O�6��<��ź���"��-�Ȱ;�uƊ�f��JJ>�qj��<�D{�<NFtl�R/�״�*Ֆw��P�4;P����6���`���R]�qf����y��o7�6L��_*�z�{�˵v6Ck�Y�z�
s�\�M[��5��z�M���t�;�R��M���n0�Fכ���.~������LZ��Flvn*�v��T��(��<�Q�bWB�������pF�ר��g5v�����pj$�8�?d�J�a��j�M֎a�;WI��4igz�~]�Ev½���	P�g֠%�5�~�_9��=S�yP�DF�[����ݝ$r/��rԅ�D33�,����J�^l�������_�u�l��%�I����$ys bg@�z�����S��u�x�z��sZ�D��
~Ɜ�S}�y:��5�.y}�g9���=\���*r�#f�D��}��;g^&�ʖ�	]'��(��<���g��A� ݸP�;�z����޲��l�^����%*B��P=�74�"���=w�~������"��u�[o�Q��c-є,c��/4ɵ����,���ȶ:�:]h0;�
5�s�v�>�P�1��B\x��%
!��!%�g�:0s�^���J���
S�pY�6���c3�M%�ٺ�2��ɋ E���s,�]�bv+g�#�َ��A�,"�G@2���A`m{�YT_��y�mr.ݤQrA�?<�g?��~���r;}CzR)r"U^|�^J�Ӿ������}&����x
�u7D��D4��;����b�ۓ��@j�ŸfI�'j��t�������tv}�>\�W��%,�mW��}�����r_G�_��v/Q�;lugO�1�?@x}����-=]a�Sa�i��|ٷpGuVD�;��S'[D��V�%�B����w�;۔3u��UN�#�ȲMW^U�D�wg��m�Žg&{2�D�0��V5���8���X��|��(䶂D�ԣ/u쥲(tĤ�V&�!��8��1�z�T���6��[p���{'l�auz[H��ΩY�XF�]���y��2 �O�+�+��ޭ�cj�V�lYk;�����Zt�(����!����vx"Ψ�ґb�x�ތ`��Ս���zu�\v�>��;�'i�D��y}�X�n��w��Iݨ��_�W�ߟwj��F?!qo�"�>���m�to������7O/yV��uL4V_AOvE��.�n�:�rh��䑛DV��;�OY{���o7����k��1����)6�|iP�$-�qOӐϡ��W@~)��4pd���m�U����I���RM�>��tu�����x�ѱ��[�gg�s;03�+Z1ym���T��H�!L��RGZ|��c��(����ߩ�����/����s]��j�˧�'���Ph�"��5���<��{���l*i�iy��,E܈=X��߆��u����۫�ohד�1dl��e^�s�m �Nj@�b�D
8�	��g��V͛YJ#w55����^dK�8�F�@R�QT� _]:��� �:P�i���	�ޥd�c;"t�S�Z��q��<O&�0��4ׯn�h�k[t�m�"��v���!{����G�n�2�܊}���{j=��D��ĺ^��Ɵ0�!o����`F��Ft��"�̊կ=e����tD����VS�^ݤ �ܷ���m�Cb��*�O�綰�kn5u���$n0�m���;iΈ�R���j��>�e�W؅�����Gu�v)�_I�n_HL�w�eZrr�s��ڪ7$�o�:GK���f�V�s쮋��������v�o�G7"-�u�w~y��yuy��BbT�����N�)�zk��4�~�}=��fuF�J���`�l�pQ�r.����߀h�=6��+wšn.�����\|8ڪS�v������!���{�?b4 ,��gf!]��"�'_t�;g�U��1�UŸ�Ǡ1���#�<�)�|��h遼?Vcr:����UX�J��CWR��27�L����n�F0�.ڡ���4n9�x�P��{x[/4M竮�|��R@�e�r}k$�f��/S#S��fg��יo�A�>�j*榕�����*�/5G�n���m�q�AN���?es�(`�~�(&�=����J5s����HN���7���^����B�[I맇5�,�p,A��p�����tr�$Ni���ջ�:rz��L��#fMxΪ���:i���z|��T����}y`����վ�W.�mJd�b��s����ՖAl4��s'E���:�GPS�)���+;��#�][�w�_�ZƪcBH������ܩaIu��]n�����vv��t����j�� �EdJ��8v�9N���K������y��i���$��Ȋ�n���@��&��u#�*59��c&�+[[]C^8���P�\��WXm$%|�"d6V�DKãƉ���y�,o]����7/D�n��<x��aMqh۞G�q=��$�*'�-�ב�:��ip9WI���+��t�@4Q��Fz�{e;:���ss;�r߲K˙^[�./�ڽ��l��`�V�Nz��������ӷ�[|�}��N{���&���΍vZ2�8f�vX.��G�0v[i�\�����6�G)ӫ(�J�r�ޞ��X9�������1��mXˋ����\룗��=6�1ʧx�z|q�_A�غv�l�����c&��@���ϕ�#�b�N��w�R��X8��-sՑl�ƪ��Q�'������:�/��<*/6����2+�6r�b�}�d?�U�[k�	�'�/�cg,U�W�����fACdxm����U��\�˺�ƞYr���\�VT�j�v#5�e3�vY[W�,Ai��tiQ	}v��ǨV�[շ�We����V���V聾�k�ù��Ѯ�R�eDyv(sYB��5y�RSZ�`p���H�K��W,�\��J/Rz�c�1�����}�R�|� ��A=�t?��=4����a�)��u����u�2���mǿ�)�ɢ>�`���Pϸ���X�HO៨)/��qJ\���s�c��:�s��M�>�tb	]'����3�s;-^����˒�Ut��l��a��Q���}{��:�┛7�7'�|��EM?_��~�ɡ��+���غ��[�f>�w�]�*����GH΄�g=EUB��v�7��TT�̶������:�ᓽ�}�{�K����5�۪5���S��ɺ��t� (�M�;q@�*+�m;�^r��=1�wf��3g�/i�*�<����}!�l58A_��+�ũ������E��,���̇�������'�WZ�|�te|���O9s������0��&f�ڨ���:���5l.�d�2<'��x�Gݓh���.�wd���N/�76�H�.�>��j!����ӎ�L��\��S�D+(,�qfuV�i7V�ba�������˙�y~x�p5�	R���/>�֥b5��o��=�r:xw�]Ƴ�Z2�g��t<�/'@�X��C��1�i��k��u����������w~9��)�͐"3�!@��^�Kk�S�Ϩ���ľ���I9�wwxu�'���twn���C~��˂~��}Y!��Y-�xgx�}��"��v�GO8�F��m�M�0�0�e»Z�Ո�;h����u՝�=;.�V����GX�1����#���f�Ҙ;R.+��'r�mkH��Q�-���.G`�;�#!�h"��k��(�lĶo3�Z���&����D����l�<�&�����dd��aqK�3N��68�M��B�5���w�+�����#�>ʹ`mMl��&�ve43��KhWc�C����#��O�����P�"�%�s��k������dN֤ĳ�ͷ�EA�w��_���;G"s&"�]�l�#�.F�@�J�ڼ�SG���p���0+4=��nY�Z���p&qVCVn�m������G��9��(��"hus�|��tV�v36�9��2��Ɲ���{��D�������y���o��:e,�N�_(�m]�GHk"5'0�Gu���4�uR���:r�k���V9y�,"^�8�f�TeE\f�J�z��(I�$^:�m�s��'���nZ$����t�f�W@�FiT(�+6��u���䨇B�h�
�J�S����\ëF���'D�jP���Sy�/���P�VE�nWF�+m��R]�9�s1ɜeيݙ��ͩI�u�e�cKcӷ���t�:��t�5%d�ȫ/h��-�˖j5Nue��;�a�*�ln�^�Oj^�CKy:ۦ�a
f;��y:v���X�d�㦚�_t�}�	Y̛�w�`}]�������GCA���;�E�*���(�ٖ;�(�˻W8�|�$�`ޒ�nL�kJ���"�4��aRCv���J�2�l^W=��j��Q:��]�

]U���0���q�������H��s�0З�����yw�,���wcG�"��7tڵK7�i�bC!Y\��<�X&�����ݍc�����P��д���'#�mDv$�U��t�]s�r^�OJ�Uf6�q%�n��T�U��Z�m���A�cKx�[me�f�i=G����B���(G=��>i7��W�E�Ty<���5#gQ*�@^v�9X�9+8i���|��P�e߽��iV��M7N/�������z[��-Ŷ2�GA����V��a#f�r�$��@�}z`$�	��Vm{*����/��v�YG�:|��w���u:ۉ�.�0��)�v 5���}Y��w�vNU�kY~>���eA������|�`�t��'ТL,c�:b���ȳ�,������'�W徦1[��j��_����u%�$4���ؗ���:�������z�.�I^ˡ�x×m��{YM����a�nC)a�L�$�ė&���R�^'k���i��ͳȰ�W>�3���p_=�\i�D�NW���ĭI�qb��{�
��S.dӽ0��a��Q��dqL�	3C��\��'�����N5���kd�/���ۘ5��z3.c�0��/[}��/Dߪ<�6�T_S^�	�7r\<A�	�MoK���غ�3"����j�-7/�,�l���i���U�=������1�ҪӐ���!��&Xm�[V5F�k	��uxԆ�G8tT�Ĭf����]�;PU�J��L���i�nE�c
��N0�y<;`[�H*��z(nQ��!��n�Z[w2tE^��N<w��*Y;��s�A�,U-��A8u��CuΥ�t�He���h����ѧ9J�"��gkh6�RU[�:�A��R����jX3�����z��4�ޑ��u�=z_U�7/^5�m��
���љ�\���t���d��`�P]oD#���7��j��s�35My"PBfsBC��u\���m�j9w�h��y�xR[o��r�[��Ly�$�H$ M��]c)A��L�ƒQ ��bHBBE�:x����nݻv�������7ӄiJ�\�b��`FW롊,���I"HF4���_]�v�۷o�^����2Qb�X�-��]�4��$���n�!�$�"FHʔ�z���^�v�۷nݽz��^�BE	@��T#Je��#P��		@�%˄�H2H�޶���nݻv�۷�=z�2H0��S$�XL�Dd�M4j1�
J(��R{��E	͹��b4c+��T������.W�#Q�������̔j+��dR��:�o7ou׻���mݗ9���X�$Y�����Ǖ�^����׮�o:TF���^b掗-��l[����(7�r��s�u���k��co�^k�L�:�n�b�ݳ��W��v(^���*s�+��\���s�Ҟ䧺���¹S�����wb��Put	��;��&��u݄�K�	(��9�7;e�=ً�x.)�8\��m4�Msm�X�R�;"�s�k���w� ��ߵ^���t�y_�}�����y����:�����c.��}]*�������>�{��N�%������g�(�L]tP�SUWPd�P�h^�{zRV�ˍ�y�'�P=�[1���~6���L�6lb�!�I�7��t�k�������;��\۫5�{%ugA�(8��ʆ9��)�q�,��]�ᕊ�>������rמ���h��mE���!�_e�vO!�D���S��L���l��|z�猈�Sv|�����߷��ğ�_�LՑL��~��3*g% 6�$m6z �ւ7�`_�rg�C%�k]��[񛜽���j��Ƿ+�{�Ɯ�ѴwӾ๻�bd�p���L	�'.�r��f�7o���=*��9^�r���ۮ׃���#cCF�Gz#9������XU`Ǯ�#:�6��$`���E޻=�U��$�ǯ�g�P_~0Ϥ)�Z;�gp�e���w�$ �
�:v��Mc0aZ��g[��FE��z^�BĽ��iN�ofn��F�5!u�V����+lTQ�n.�_�����8�l;ۻw�2�T�}��
�n'�'^�p�j�l�^�:UǛ��үF��{���G�o�_��������&	bOY��W�-�|�q�"`֛2����P����R%=�.�T�u7��6�sک�]��I����G����{��D*���tک��	�%T33�8�5�;ƞ��{X�X��8YT���")�.pD�tNwu˭�Hi�঳�V`���T���6�M�@����g������	��h�mr}`V����%���"��c�P{�#r�Oc]r*�$޵ƜԄ�p0]�Dح�ϙ	u�����H��j�ɍ�W��U}xs�&��0�u#q�w��F��h������J���'L���׷��g��T��};��;K���Q}��j�X�:�����Ź}�՝Q�7����./7]j��6��C�oTA[s���j�·^�g�1��#s:����ʝ�W��T��x'�`��W}��_�����WQ�ۺ�к��*��F�v��H��s��&�+Ps�NC	��ڵ�n��q.Z�Z<>NP� ���m�e��>T�<��8��q�%���K�2��ᮬ�AA���6^�/E5�%90�;ڨf�d��WH!�>o�2
�u�){����n��{r������[w'��������q�ǖW���t�O^����YZ��4;�V����@����85y���.�;7��7��=��+��񷔚��f�ӯ<:�A�7<��Ϥ��\#�*u��x�.������kM�Q��$G� ��vu�W��$�2��U�Y-�N�m])d5=ܝ�U8g� ���y��q�Lu�@ǢP��?��Ǣ ;ǹ���+��s#�����]�ϛ�	f��T�3���B��}gGtx��ʭ����griș"�e����s��vd�הp\ӝ����Lk��H�|i:����5/H�������g���rX�p��'n�5��52fhf�6�yt�R�Y"�Uj����_zχ���MםXD
Y�:Ft%\JUS6���ȵ`�gL���Tz�k�N��27��S�pv1Žxa"?X0��h�e_1s���K��d�g�еv9e�

ڼӗUc���ǾĚDn
ɺD<w�<�!Y�wa���:�4��n�*s�f/�X5J��r��G���7�\)^]���Ox��S�n���=�sk�5P$���/�G�ȃ��?7�$�M���ԍo85�H����N��6�˪�����Czs��X�+;gݷ�Ŷ jA7���c4�ڹ�z��уzwʹ{*2h�GZؑ�KQD���B3[`5uu�m�˗ݪɇ4[uM���^S�}{z��\�+Ή�mv���C�[�D���m���0�@`c�L��j���䶒&����͖��-"�9��|�$px�7IH^n_���=�n�}�[���k��vEϦ9ڦ�){�3^녔���v���g9�G3��m�
�������_������pbZ���#���n�����:�:Q��;�ߴaىXj�a9��LC�>?(.tn�!�(��y��=�"�N��y{����~K��q����O>;r6ϝZ�����;m�g�����}��Ў#�j�7�~1�0f^G�*ur#�w�7�ś>����0ސUV�Ta��:�IwkT||2�Q6 �tg��6R^[ޗU8�
��MN�kr������G��Vf���U]I��[X�;S9^�[̎<�q�B�T3I�7u��:�$��a6��X�]�o����k�zv�1�c�w�ߒ�y_H�4[�V����$��Z丰H�y��V�6�3���U����v�3����Pٱ�V?���TE ����WCJ��,6XnF��-;F3���ݻW4�GSV�d���}���q׏��;~uo��tfѻ���������)B০NUϵ[��ǐw��s
ԖآFԷ5����:c�S6�6	9��<i�Mٞ����EUyC� �� �����1�;��;���\R�g�zRV�h�4;�Q�<���~����n��T�s:rq�{0��EgP��.m�<'F_r��K���Y���1�]��뺪����S�z�l�d��Hޑ��Sϣ/ӵ��3\��(Ȱ��B�<dq�W���UHRׁ��6��m����&`ɺ���NAZm���z�Y�f�����=�h�Ъ�z���Fl7��Fco|�O3>=4s%ST,f�E�Y�Ӭ������V��s�g[R�6��m�{��Mr�"�
!�u�/c����}��r��ە�q�2���&���]�TEn4�&W=u��X��q«J5�F����vT��^yu�o̧��1����9�����O>����Ɩ�<����`o��� Ȫڱ,�5CKF�(�B��+�Z��v���{�Ǡ鎐�]�JZ�sMc����wu��=߫z[~I��!�ņ�4!"hV_�$ga�� ͦI����bH7c�X]}���$L�w3�P����Hy�h_8����&BDcf�xv�݊�O��#)��lыu>�`�zP����S0ި�U:�v����Cm��G�f�n@�m�y�	���U�0�����U/I�F:v��5��r�B��9w��{ ɵ=@�֐z�����΂�� ��Q�����R`��+63���5��z�5���2hΪ�v�}�O��=��e� d�K4d���=F��B�u�آ&��W�\�#@�'��ߊJTj��ˠ�5��N3g�y�M�c^�T����[����s�+�����_��Ī�3����uS�o�US�/���V��D�;���Kzm��v_]���EU��b�=�����wC����g�!�<f��~��Q(�y�A!MB��t�s�.wR��z�8REq�NTn�e�nN���믋�1-�FZ��!ԆJ3�Y0,Nn�fouSV�b&� �I����.HM]¡��c���_����v7$�ƞ��wxy������u#H�9�w���
w��g���ˡ�S��޿\u����>M 6=����3Ѹj��8gf\1���%�ۢ�뻛f���=u���v$�F�]���B��cd�`��"!m�Xx��bN+�����ξ�|�vfm���<�,��6B���=�}�����������V����1,���P��ސ3��w�����soN��ށx]��-��9Ì�p���պݪ�צs�n����)�U=���N�t�C��k8��<�=~
��5EZ=C�g܉nΚ�'g;y�>�l�"1�T�͈s��xThE�6.��ޮ�_��1#n����ꔗJ�iD��u���N�j�Q�.dYg���L�-i=F(r*Cw0l�ӽ��ͺƲ�-^k�q?�{�(��|�:��X�tR?ߨx��;���r��ކZ`��o��YX���4��vRs5v^����|�{�n�ȳE�w]��x��9O۪B�W���Z�~�}��Ng����B/�%n�g-7�PY�1�T�z�-j���ب{{�����^>>o7����3ƴ�}&����~���7�m�2M��}yfE�!����E�l��~�0-�[�:�~��L��o4qIc��]��qZ�qvZ7�F[e�y�Tuu�ǵZ�K#1��1[P����,ϯ�+o���y9r�z8̜���9�l�i�O�9��R�-�.��<��C�/�Ӥk�uq��x�a�1Ȱ)�`�CMŴ1��{��7|g������7twx�O��{�T�vA��[i�[⌼��Bc�f��c:{�S�~��"D73����J�t����5����z;���M_]���h��l��%�L�/X�S1�ޘ��p�(�0�N�bv�f�^K���Y�E�,��`0)����S�'���Ԑ���km����u��O�b������@"����P��e��[�2�����,����us�A"m0Qﵫ�/C�6M򘭂%����1�;4���f�>,#|[}-0gN���G�.�#�4��Ӆ��=.��-�m�I�pJ�/&�X�Ec�m�ϑy\k!��c���۫�ϗ�S��{|�zk	�箢�}<�����ڌ^��#y��o&�h�w�$@Unϗ8\N�^q&_���Po�w��׽���9z�ߧa���o_�	�bRl�jV����3��*��Λ��V�9����2���9-���[q:�p!E�dn'��.���[�뚞���#=�Z ��I�ca�� ����7�'���w��_�% �h����D��L��L��2���1C3�֤e5�d��M�6Y����8a�6e&�q\7�������2N�鍐|#3$}�~�DX\既
�?XsЭ[6��g7oLoM�U��Kw���Իخ�|W��c��8�k��Ymx͔[6&�Y�鍜5$Ĥ+�bfG�,�ׂ��S⊪�5�35�*޼X��
bf[����Mlc=E��5Υ6\f�$iD�Q�H��=��k��2;���P�苣:���t�X�Ǔ���c���[�h�a����]m+b�$hs6���2H"�@�N$I$��N2W�%$Q@��( �	FЕ �)��,�;-�j�\.�@m��+�K;���4�Ȥ<F���FWU��aӅ�w������+6�r�0�پٙ���uo����7����;N�Ic^|����dX�"�����d�0�*:�����V��H����I����n�F�j��jכ���e�b���Ed�a�j�0a��@M!�T�i~����K�cd��v�7��H��raP#�OS����r����b'���OJ��l����5����<Ьol��]j��X�ٛ�r��3��N�n�F��d�<T�y��6�ʗ�xfxܢ�1f�}�ǯP[�Rh2�����'9{Z3&+�uuB�&fh��>�P�]"�Σc��o8}4<���n5�c��G:�8�5~�}v�����H�KL���%O){*��cL�d������@�.�{q�xx�B�y������z����j�xx�;��ϙ��g�V�5���ԙﵮ:�ץ�GN�U痟����V��*��x�(#�/�?�k�Tg��hh�T����>��B��H�R!em5&j�SL�MF[iY��em+5���iYm��Ե�SSZ���kJ�m+-�ƥ�3SSm��-�j2��Ͷ���b��X�mY�&Z�Ym�em�,fզ1�ڳ,�R��3V���5�Ͷ�c[Lfc6֘�f�Lfٌ��ɕ�,fem2jkl�f�MFkjV1���2Yke�-i�3mSQ�ibͫ+5idɖ�VZҳV��F[R���Le�1�����m����L�ҳm��5iY��Y�Jʬ����6���jVZ�����x�J �b,�0�j���V��YY[+5eel�������+5��VVV��l����ef�VZ�ͬ�5ef�Vj��XA��Q��X�G�z6j �� �b�R��T���J�کY� ��P �A�PY[U+5�R�V�V[j�fڪVmj�f�U+-j ִ�PQ ��کY�����R�kU+-j�emT��U+6�Wr
 @b( �@`�R�V�V[j�eZ�Y����j�f���z��Ԭեe�VU�f�+5iYj��iY�Jͭwjݵ�f֕���f�J�ZV[iLA 1T��Mk@:Q��ZVkR�kJ�ZVV��ZVmiYV�ԫ]�n�ҳkJ�ZVVҳV����Օ����eZ`���y���Q����PAEPR1DH��|
������~�����p�A�OL?��?����
��?�� 8#�Y���;������_�ߴ *�������?����
�
��`�a���䟲/���O��!�ʀ��3��������$��ܛ���?�',
��p~a�%~���0�A!�j�J��V�U�*�J�Զ�͵���-*ҳj�M�&ږ��V�Z[-i-��mi�[M�iVmiVV���j��+e�E�$U"�"	��iiV�ҭ+SkM�����٫M�mii�KSkL�Ml��5�SkL�R�kJkR���jjm�ҭ3kMem3kM5h��U�@D�AIIdA��6�V���*�kUj6���ͭ�V�[m��ʴ��U�kEZR��V�a#0D��BP�_���~)������) � ���~�5����? �>�,���_Ђ����P~����~��|��K?����[a��q<?J}� 
��C������M�W� ��?I����iATE���uЊ � ��_�(?���F�:P@��W߉g��Q���@X g����?R����� _�1?����s���Y�����C���"����ƕ _3���P U� �г����ק��h�`J'��~���à� ���D���P U�=�1�ݟ�R���wA���_������������
�-TE����ߏ��`R��b��L�������� � ���fO� �y��|� �-�BIQQTPJ�
�D�D��*�-��R�TE(���B%D�Q!
�T�P�B���J�$�UQ�$HR���������� ���R
�$�U(��HH���'A��U(IQ	 (�%T� �A)*)U���RDTR�J%!R�
��TH"JHR�GM)D�*��Q�*JUR��ER�
��J��J���E�IQJQR�  qW�h/n�V��B�VԖ@����it҆����J������R���U��i���0�i[�尚�A�JR��m��m�aэQQER�� B� 5�CСB�C����<{����hhoz�
�
(Q��=Κ��l��N��4�4�i��emN�u5)X[avw!ەC��f�p�魲�UR�%�B��%R�^  ���k�	l�m��S��ۦ�9sX�!��%*Sh;��@	X��mN�YCi�J��kn��jtі]��uݵ5e,U�3m�I	Kl(�
	*��� ����uL�4샹N�A���l衲��@�Y�@�lR���
��8� )��M�4�J��U� �'���2�-��w ��E�Y[�쎍@�������-��Q@c,��+��V��-j�E"U	ve%B��  Z�Q� ��F�Q�u���1����٫ij�U-q����(kRۥQ#C(m�wD�T	!	*�%P*�  ,�I))*[���2���c*��9�r���*[�wJJ�AgE�n(�8u��I��M��P$���n�"�I;�wJ�5���I$�I*T�%��  l{�ZB����R�*���H@�+�I*����MĨ�QXu�]��)Lq�RHJ69��El��)�%"�d�$��PnI%($�QD�J���  �<U"IV��UI
[v�RM�&$)(����t�RR���JWmn�qP��j;��H)7��Elu�۶uJ�%T��R�  ��u�K�c���DQ�ے�;0;��IIN��kr�5TΧt��I�-s@�gGpR�J�[
��ZmҷIu�D��O��*�d���a%%J2 &�CFM0"��	IT& C@�=���T���  ��H����@'��G��?�@�����_����L�e�f/z�)�1&�d�������M�2'� }��|>��˪���U��m�j�Um��*�ֶ���j���ʶ�����mk[f�UV�����P�������Y`�a�Ɍ�$E
�>U�\Jm�v.f�B�9j�+/v�����C*m �_��)��*Me�%î��eRK�w5��0,e�V�;�MB�m��֪PaԚ3m���)�[�e
� T�l -�7��fA*[bh9̿�����s.�-I
���l0��F�����T��5���1�S$�˷*��KM���m���A�.<J��5J�DA�v�X0�6��E|�n0���7y��m��w,H0K*X�x��r�	kC���R��A����v��Q��C��v�!�,Qw�Y6����di�27�m��vT۫%m��Z$z��[%����ika7����I���J�_�c���P��WV�I7n�S�m$����
��@k2�@�ܭ�[�U���
c9P� �ϞBJ���y�J��L]� ���L��Gڴ�hi�dn��n�qivȗ.T�F�nJ�/��]���C�;�,����J��jȂ��A]��&3U�\��xlmBy�	7UP��v�M���f%JJ�:��+M^��# I3A02�:a�q�֩��tJ���쇑�7t��t��F���[O0K�G�ؠ�b:�Kbуb�m˦~V)m���/wS�V��ī>Oi�9x@ű�n�a��P+mf1&.�jd=G����`9C~�2S��H>����,%YB�3+!+���3 �ض���ol\)}��U��G*h�=%�NSk^�I+�l�-��Ņ����NEj���Y�Q�9b[�M& ��E�kP�.�H6u�%�Ҷ�=���ij���m��%��m�-��'BL�hEu�-�v���jl�cpVniLk�B��5r�ze	�piGac+�3D�1�h�,�l���$�:9��-D؃V�j�%U�L��eiVk>*��S�Ab�����J�n��[���+"I
*��/�)�^�\�����0"��*h�t^w�#��`�b�f�Y�[F��N
{v���jr��v���V���f7RfXw6�)6�J�#�!�{ ��jz���3Rߕ	Y2�D3�8"�ӎ���q�W�V���s#����c��.�tn J0m���ӔpXŔ�ld��B�ҭJwR�Ɇ�
���8��yS�{V����T�N��r�k��h�(r����L7�ylU�Y�U줒�/N�D�G�=*�ٙ!Ӹ]�r�N���k�^ƫkr�=�[E�`��֤F�p�'2���1t6�&��J�۵.,����b�j�ˉ(HB-�ۚ�R�x�^%��w[���ճY"�n���V�Ϸ(^ n^��r��r�=ņ��(��⡢��N��p��3�q�4e�X�2��0�8�BHP���MJ��bc"��5TZ֛�/)��{%���5����գ�pF�[̼�A�F�9nV�����B�n��ݕYc��z���ؤ���n�8�h�kD}�����И��6�mՏ�nVbUa��8+M�IT�q	��vl���Wy/w].\��^�$ʊ��f�v����2�V�I�,�*�2�!��w7)[�w)��mˬZ-���7�^�z �Y��o4Q
%��(fl�aaPqͻi���v��JcW`�S]#�	� �n1B�j:�k�+p�-���D�ҕ�.T�-+ktk�������`7�[Y�O�]V����RT��j�JD�ͤ��b�������S.�6����ҕd�f�2��):cJz��wp��ۧ `&'ی%��읙0��eТ
��`7�M*�9��4���o,�9k+`�&e���(���P,Q��]�kBVt'��!,�#J�ˎ[ f�����1Wx�/F��� ���Wb;��	����f�fb�ᒲ-�P���w�ڄM��ku�Z�ƶJ�wT^PZ��4�M�����("�1|�Ȣ�F(X�ehTr�������7-Ӫt�
�7L@��J�<���4Iz����j)�2���Lɠ�L�nb����z$�odT�ܗBy�Ґ�Rv/p�:E��2�˽8^1u�j��fR2ejV3խ\��Z72��Ԅn�՛�.��V�Mܙ[�kh��<2i�6r����Y	Le��N��5#� �&�,BSR�4n� �
�X�h�G�F�)������8�#��a�/m-uljDf�@1M�	��E�ʹ���m���v@�=y��5J�mP�i�,���}�3Z���[Ejd���	��쳯4�L�1Qe84��n�B��b�V�ʘZV����RLD��7��D�Y�����<T������ �&7-�+�=3]y-7{�0ch�Od�XPѮin�V���qe<�*,2j�t0�5�/3�+%�N����ݲhݴ��ವ�,��1nDA��eKTm��X
�ώY�l�`���ɨ�t��uE#z���!���-L#I!�i&���KLV��Z���*��c�(���'�4�F�Oq���W)�����`�����9�pXڼk3Jp�e䤆�qP_2�_]��1����aPʺj�KSpn�����@��i� ^k˻ܡ@��RF��n��m$\R��t�d��WvB���dm)�Qf�eʍ`@T���kb���nܖ�ʤ�p�-��@�ɧ��4�#���v��+ 6��y�i1╩Q�wI��c��1�d[5x�ǘ�,z��t r��0��`����<X���6J�V�[��m�7n�Uaa��s4n�2[�05)��X��J,bEu�d��ر��QU�
n�"���Ǚ����YmT�ə�T���xތ8�V
�$�sv�in�V)�W@1&֣�2i�d�P��.�,&�FfA��Q��� b�jP4�;?�5���m�(�@�{��eLV(iǖB�Ch9�Cx�1����V30 ��@eh��ʎ�U��F��p�.^��w�>�.̫�$��W����a;+e��i��/^&En��ͩ�\�Z��i�n�b05���a�`:5�-Z��N�`bӪ�5l�STQ��M㗱�ne1��÷v�Xq����&H�A[��9�lM��H=
8���ï7n�]�<R���\�ʽ��jЧz�+T�G�V��θ�l�>�C�%����� cU��9Na� h]l�����&��T@E��=���k�i�����m\ǉ�!)೿h��-�a+�
1e&���:Z1�F��c�٢�,Yn�P�`�E�m�QVep�ګ/u
K,�Ҥ.����X��qg�)U����0�iP��Y�+!%�iÍ�&h^��F˕�N��A��6�f5��F��P�(VRĘ�B�|Cr�3oef��)�������&ݡ�Yb��m�+L����,eXN���Y�R���F��MMo0�ӕS0�SK%m�[�7xh �����T� �;�2��z���L�9��lf3��"��p�BR��*�W�����3�x�Y#�[�j��,�x�L����S�t�"��Լ�U�����s&�t�*��Ds0���2<u���nX9��@�v������+YA+W�,����MZy6���v���reT"V�d-�z4����ۥ�1$�-sf��	X	�K��P�m1jAUcV��ke�V��8�x
���Zs	j��yiЄ�4��*�)�yTA��(f�Ҧ�h�Q��6�fkK2� ��j���W�� �	ԑY�ʷ�-�;�:��.Z�+F��'��4�L9+��2�F��2K:��y&G�ɘ�j۾f�U�n܉�[J����@�;�V޺��aZ�/q]^k/��!<F�M�DdQVZ�P�̬���[�zr�A�i[���ww[۴Jh���D�+4K$��!cĜ�����I�Ca*�C.#q�L���U⛙��.��:��/�0
�F�h�D�Qb��.�νb8�d����wN�!��eCoh)x�yr�۫�i�"jH�Ś�2�tӬ����
{�]�^�D��0 S�
�Y��C8�?Zl&mK�ҒJ��aĭ*6T�)jH���o�#EڡJѫK)�q�tk�jQ���sh�SU��)�p�`�v.�T�4����n�
Wh�B*�8X�R�v^I��f�8 $&1+wb8p�M���q=��N��t���֘M���m��سt�+��Qꭽ�md�fŗ,��
���F[T%�[��/H�xS3`�6*Qª*���(#g�7�Z+P��^�Ӊ��jv���^b����&J��J�fB_��坠ј�47�OcwpbU��Gn|P��-v(��îSqcd*���0�LH0t[����6�#R�:��#0۸���0<i-�,DoR��f�¢�S��jt I͍�XԭJ���$����fsf��)����,1���R�`ԟ�֫��!=82�k��Q�Li��D�ZH��PZcI��@1IЩ�<4�������6���WS$U�uw��!͕{_שe�μJ����q�5`��.-�1`�4�J��v@�eO�W{Z)HA�	j�m&��A=b�h���$���ivhc%[z�pk�eb7�ۏE�Z� =�bV.��)�{�{�駢�n��+2V�ز��PU
�X�v�]h0<��.�d�ZLL$˔�t�h�U�.E�*z����7uWqJ �@+�h^L��c��x6%�kfL@��.��LhܢS�ĭ���Oa:F,�,#H�h1#�r��{NS��[5�bT���gM��l��N&v)0Pq��-[�kC.+z�ytځ�۸�D�gnb���^���B	�� JK�)M�c@�["ܭ��B.���Y͘�:��:)n��Rĳ2M��S��`�wM�a2�8��G2n̘�`��4�n)%��� 1Wd��K��{eJ��e�+t��Q�o0�$v�5�u"kb�W�@2�0�ڴ�<
�V������H��w�n�h�u�� �����3A)U�ɮ�;jhE����f7#����Q�Z,��qJT�4,b�(:����	s(��;��&�ǲ@c��n:��os`�\�0��b���{)�2�����RK\��V�(6���a�����č��f<n��Dd��Xzh����L�ׂ�U�rmَ���`qкB����2Qʛ�,$�6�M��@`:��m�s�su�6dKE���U�V��6%�I�6X{�Z�2][�wk2���,L�&֋5����T,���ۼ&��T+FZ�!�ܦ�K��I�"��p!���Z4�]�0���p4���R�j�n�VU�%9��٫5u2��(�e���&)�>M���W�XM#Zl�cBY��ǘ�]53i�ޭ��U�A�m�Q�Y�ʂdX$[���#9-�T����;f촱�.TG>Ķ��?Cb���{�-ՠ�\�Mي�������-ꬬz���)�KoJB�Խ*�d�/#a@0��2��=�F\�P�P��;�`g �핆".�]%�D��R�t&Z�ݗ��U���呪���K�+ ,lG,�t��n���.d�Ɋ�V�ۂV��M�1zI�R�U�EPM�9�a1�dcs+e��i�Nn]�*��*]������6�K��ih������M����u�Ť����%��v͌j�Æ@��aH�˦�T2^�6ͩF,�[��oC��ϱ��,�x��w*��#n��f�5�JdBd�<eͫ��W`4�F��6��r�:�c,I[�jpj�Cnb�պ����p����ˣ���8���t���iU����N�i ���<��kwtct�Y�Ӏ�(*��ɠ�6���ó�o)�G)Ů�@��ON�J�-be-�t�*�^T#Bo�����`Z�V
r±w��b�BB��%���)&K��N�Z4wf�b��dL�.�d�bF�[coc
��h��)��[�P����fA�%S�pX�,X�跑l�Y�]弭0��UWV�Z�DR�ۛJ�e�1�1�a��P�ZӨ��BkFY�	�'I���D�S[Oj�)��!a,�ۚ��ܧh���Hdz P�f ��ɻ5�.n �dI��6��Jɤ��bX~����h�KU��8� ����xЍ��Q=��oULM��)��zI�͚u�٤b0�6�����t#�&IU������%XZr����t�pZ�� �QSa�-�$W���Z:�i�Ը�%<�M��"���S��Kr�{���n�ԖQUm\�"���(8�rmҽzl�H;Ҧ.0���gʔ2�TN�,Y�bB�F븅 �.�U,N�\{�mʲX J�+m��4X�5��#i(h+�
���E�D�	�ø�¥����+e����lXG� ���TuD9��ʳiQv��.�R$��@(˧QL�i�t��ӛ���mޫ֚{)��ɽL�o��j��L1��N�x�����F�պ��ю��C݇��B�2#�fX: ��*j��×���q�M�"@!-ADv��u��U��F��=nݵ�,!z�NU՚�-�y���"\�ZO�!�����w���j)�%;q+�AI�sNd׋�%h�1cu�����)��	�Wyx������(��b�ƪVեv�]ڑj.��ct�A�hTܵ��YV4��v^
���.A�Snc�q�gh�]�83	�Ɂ���/R�2���L�J��Ƶe���͌ףa�2�m��a8F8$¥�B�)aR��.��)�Bo��`"��(J+4,c0nmn��N�T�S2�Q���m<ˉ�j_̧{Q���8�],P���"�c�Զ��m�[�hi�1�ab�j��Kc04������˜걚T�9 `�ή�;�^�腖���j*�f� =H�j�F���ͳju	���YY����̀'����og(��S�0MiV�[cj�[�"�hLy!���	�tZ�'@k����N��rA]����<�P��c��UV����95�n;EXۦ���Z]+�$�z ;����j��`̷�N���{J����XoM:�O��v.�w3c�2��t8)���.�^�`�eXm�����&�4�P���&a�{�.��:���_���Y�5�g\ģL� ��p��X�Ƭ"-�Πײ�ͷ�����٣-%oS���c�mZ*R�}YO�]�(�w�[�/�G���fkUK��b�bm���P�6���t�}y�b����*�I�z���=���[�;��n�d��Ž\ӳ]&�e �:\[՚ݛ�tu�����@p7V�w]��b޼��S�o�s-mJ��.au���M��Wk�Z�9�lw����E��A:zq��ԳU�כ��|�8�7�c���8�&]����]Io��i�����2�N8�ζL����Q8@ʹ�8���ԫKn��v�H��	3��l�p���&�����-�vv+���2⸓7�WZ(�1;X����h�<��1�P�m�dnl>���`�9�3e�\G��z�;/M�Eh�1��
!��Y�_�7lsͭcwa��owbT���.�qm���%�f��V,����L�C%qzq�N�\�wCT��p����V����s�',�˸�� Z�����Y�q�j�#a��=�u�NuN�΍�q���{����a�˴�|f��=�ɀwS;����n$�0��p��wH\>��o��H�vlR���b=osS�m�=t�c��5�v���뱣���RkWj\��[`��x-lLXdܝ�0�E����-�ղ��_"D_d��e��-���h!Fo-u˂������A��7����+�5;wn�.ub�Yy�")�FegH'�J(�
ܥ)e�&�<Mʊ��`��30`gV��W9v���{�u����.�F�2*^�q��`�.CyYu��u��8k��!��y�:��v8%K����o-W,Ԫ����ײ[�f6������|FU���7��e���һ�պ�L�
-��oPZ&E�v���:n���3Ao��Nq7�ܧXƞ/h�i1�ޓl���f�7{���7χ.6R,v�q�架�ǳ�ŰU� ��ښ;%�۹�V#wݴ�V�㻙4�m6w�(q�L��%F۴��U�"q�X�jh�e�R�L�2��/�X+����8�; �ZD�ZF!W{\�nY\؇��S�.E:��YU�R�\���u۷��෌E�u�)��<:��3H|i9G]���[m���r���$ҕr�<R/7.gb/XK�Ҷ�V(e�n׺�̇.4N�pw9k�c�P��!X��s��C�:�bև<�*)txjP�f雧)<��t洖���弑:5��3tşr��������]���}�\'9��б��`��bp�G�^:��Fu[�>�,bǂ�@�
E�ʮ�=
�8�Vd�#b�]v��ʁ�)s�U���[Ű+�x�q�]d����>Q�d�әw�Ik�;�Y����L`�k]@YY"�ʯt�2uK\L�G�{ۊ��bR=j�c���'���ǯ��y>!<��ґ��L^��[�lJ{���y�($q�/����� YS��c�#�lJ;�|�aˑ�=��\�G�\_I��tE�$����l=��%T�ºFu��;Ph��pӌ曝ٻ��x��J�).JFD\��q\�
�b�6񞾭Z4Y�v�t�Oy<��گ�'����{�+���������(݌�j�W]wwCZ������gM]�H��J����I���8��5�F.��-Gʨ�<��𺰞���5�b�bw|݅���ص��U\� +���uugZc-�f��[-�K8i�gAsu����n�W$�a��3�����+>��,�r��ʓw��Yx��Ԟ���J"K���V�����ӥj�Y���/�ut8U��@��~�eZ�ʍ���<=ӭXYIHc�3�v��oHه���M'Wr;�[؏�k�i����P1X�V�a������N�l8�WE��v�`�,��#�y��7`�M��C)�h�ˊU��,�\j�Fi:G泅늠˱�Pum��(�D�3)f��wYN��>��Go1̑4�/��^�����=1V����i���cc��۽�wČ�u��vЈM�V��:�W��ȫMN�xGۯu��������rUڣ�k�K=X�:��Yh�GһO!:9�6�s��}GOȸ���Y����òDv$����������2,��Y\����ۋvf�9V��-��-}��BU�}�Zo(闺���J$�+M�QʼBl�u��vp� ��vT�����5��E�S�qD�q�=}C-�5W)�i]��3��hݾ{,W(:�	0�A�gn��ohmN4'6��m�_�m�v�ک��;�����H�I��v�N�m�����x6��.V�ޮy���M�k�=�h���5�Fʧ+Y��u�Y3\=o��v�Τ������S�u�d��Ɠ�c�\Q��F���xʲ�=�mⰝ]�m��u��L3�\�(fl��V�kȑ=��b�:z-�;��a�@fӰ{Rw�����;�/��3o)��V�6��\�1�7����s��)����
�d嚞�Uh��ڷ3��Ռ5��nu����E��l�#@f�r�l-LiT���S��q�X2v
����WQ�Va�mb�t�m+����-�%��:w�QV������ܱ��f]c���:4Au�8�2u��8��Mڧ��.���{z�qJu�dɕ��7���[����rWe���(!��f&�݈���Gl�{fs�k�eE�,&�c(� E����B-�����ή�

��y?��{���g���8��r^b.�N�Q�n�'yڈS�3��7[�8�զ�|3�Tz^�csx^�j��s�]ʒ�oz�g%r;6j��
�
�II���:��/[ĺe��J)�nm◼��+���6Z�O��K��%�v��@�Ť�L��4��y& �f�����[�F�i���U�eM啣0�E�Οbhau'Vٹ�1Ѳ�@n꺵�1��r}|Q�P���Nҫ��ǔ5:��O���(:��1)���T����N��'^\�2,�k��'x�#�^8Cb��x�d�M�ۃ%G�q�,��]X�����uq�01������ѫ�R5yy f&�܉�81��6�v �\��͗yV��a�	X'�q	7�mccF�rܗ]:���&d�8��Y0��	�؈�8�T#�LK�v���yZP��B�:��z~��[���e���u�4� �m��N��H�U��]�Bz��.N��3��|z�s�1\}��`�A�۬��VC�Kh��5�B�N�Ҟ�T��D�9z&^A,j�л4k8��^h���ocm�EbH���D�d*��P���@��
���o.���;D%��-�!�v�&�K��|o^����� U�*w:V'g%��v��4�3d��U�[[�����J� ��>�/�.�m-���P��w[�V���W"̮�V�����1|�nG�!B�Ү	�[>���u:ΨF��5��!.��껮hu���S`CO�v�5� ��o;��nct�o�Z�/�\N��~��a�6U�q�D��͇��u�jNtz�)�O�X�v[�^:�u�w*K���>�Xj�5�x��)/<u�A��{�yjTm̛�1W4� �����^/ï0�,�K���^����O�a�Qx1�W��O緈��D��1v)�)ػ��Շ/��B��W^j�:�u���MX����투�t=�0�����Q��-mvd=a����15��ɏ;f�s��I��u3t���+��X��NaE6�Pf�(5�9t�D�b��w����z�qtS\�t0s�����Z�X�:P���Ak���X�[�t�U�`�@h�Nc=���֫&Ӻ�z���g�m��
�J�U��ڌfg��G���NuE���ͬ�� SZEICx;�����ȥ�݂rK�ًWE}��Z���/n����{n��
�b��,��Gzx`�zHzƈn���>�؂��x�r�qN��I��2��x�/BUӛ8-�u�]��
9�J�����C\ӭ�����ї]ZB�_��Ô6���y�K���{Vՠ����[;B��Xp1�ZEV��y��޲޼Tٽ�
TZm�:���/FxH�3P�h�Q���.S��7B�ż	JN�-���9���wL�������(b�|��Ֆ�k���$�'�)VsiU�xn��d3Oj�k#1\הCV�:�;�U����Y28Hֳ�A���q�u �v�@,��\U���u٪��b-�>�P���!L[`�`��cA$I�������U�s�R����Y����³z��:1�$��^e^rC;�9��*b�(I��T4:V@Ү�t���T½w8�v(���a�	�yM�1rgB�<kIdj,p.�jj2����Źj�v���)���U-�ʊ6{�yv
�L�=�PR�uj��&I��(e�nt�
�N�|nS1�K����Ӣ%tf�W�v�qT6Q�����yV��-����p�m�yE�_EMg+`lӄ<�9�N�e.H[x��O�<EA�d��i������S�d[���\5f	���o^��٠�=i����e_<71���/��w�띚 v�ޒ��Di���VdC�S���I�ѩ�PiW����f�ͷ`�:��݂��2��Wf.�`�|9b謽D�;��aL2~�52�w��)cO�=O���\��D6���vo�1���A RŔrp[���Gk��<EZu��
�nm$�D2P�%�Y�&;�:<|f�ׇ9�r �^vհk��C��яGAE��nI+���:xor�����{��$}�#y��rY@�����;;�$�^�V��M��w�zT�$�۩gw]:�=�wt2����ڃ�u>���HS���'}�軶�`�ec);z�)GKMt<�K�u�����H�u����%D�㾙Z�2�M3K��2�F�����>�Î1f�N�0[/��TDT�4ܠ���ww��euE�s_tmg<\�n�h�hoXJ�^ &n�p�3�lq�c3(�yKm��Z����&�4�Le��bV�AY�)�NU����w)0�`[q˧n]�B�9���
��.�\M�IWcw�+j[����I�l�)E�H\}Gj�������v'�yj���o)�]��h��Ë��x�m�jzyE�u^W�ݤ0�|ˊ�vs�se&��E�U'DX�f���*l�sW=�KFVf�K�y���z�1��J4Gq��'8���e��{zkfRǭA�diԚ�}ZD��ԧ�WӀ�6�;����2�#KOܫ�.h,p������a��C5(�x8.c�C*P^���C*��pT#���e�3�oCi�#�n�ѵ9B]����"�v��ג.G���xXpEG��ؤw�.�_���Z����3�+]M�{D,OS��:�kʧQ33yc���>Ȧ f�:�Ѹ@�"�G`�fB�ڬ�T�y�]jar�Y�PR�sP�;9κ�)�j�҆֊�%�7 ˧����;a�2��/r��8!�ɮ��*.�О�QQ�nrKt_Wd�,��Lͬų /@|�T�U��}��Yy8٦��BuL7���9G����}[X][�B��b:7�N�L��R��=��B���!p&�[smZ����3�5��o3gg-�N��%*�Ra����%;+NPR̹�������+�y�#�W�șe�OH���ʝ�C�\O@T�a�)jN+�"+��;�ɚwOe8����m���;�'�t�������[��ćE��-V�p]p�|U4�����˨�ڇN!כ+ e�7;�e��	�� ��e�fc�VbM��<2�W�IW�v�c(���ו��2xm+�FZޖ_P#���P�O)�X����,�{��s11t��k[�8���P���/v���%oh
��Pl�piY��pl8BpC;���d"��d$j�x��$�b���u��V���GmC3M�I�;�k�T��K
�ٽ��L��0>�7/// ���YM(�I"4m�n�y��{�|\����}F���w^��V���LWK�,������ڼ7�VP�]��\�\�u2�����Q����t��Y�z�[ʀŬ��2�tN�E�R�wط��+�}J��d�[Y����n�4���~��d�f��s���Sl�˭&�b�^�!oo7�1��]�]�Z�˯�;�=x'[����� e��v���-�C)`�z����%�ع���A�X�J�n>ԇu^T�u�u\*�#7s;[��J;bj	�؍��]ɖ��gh�w�D�iY>�Gҹ�-ج��8h��}�u%X@}E�@����#���wMb�r��X��97�?�G�*�l��w����>�;�_���2���(VWZW��@6��ō����
`U�n��A���\�,KwH�̣��4s�.���L���W�=St�U���T��E�v)u��u�B�oo�������.�i��F��㩃xn;&����lB��ٷ6r�Ĥˮ`���DT��B��d�C���#��r��eu;C���=�)���V]64\�Q�������˅��R��%�0T�b�U�k���$wf����4���o�����ilh$c1N�B9v�@��!t�C+[��;&F2'gM��e�#3'c7�QN��]XQ.��_�ꪪ�����km���������������~y�ꊆ�.٧�Ⱥ���/�Rr��&��u������YyK�+DӔ��49�:F9��7������v�]�#���t:�c�9n�Lz;R�j(/{
���ͭ)�wB7�sf�FP���wr􍏳3u�1r�kHx��:���Or�̎��®��@$�iA��䇳��7]����%p�];5����g�,@+��r�t���t��g#uH;7P<o��oYZ]v��]5��%�^����TpVK�kE�e��[�ܩd�J���>W��B����kWuؤ�Z���0QR�u��T�d��[)(b�y�i�b�H�ǘ�n˦�t���(��8������3Ilp9�=F�y��z¾s@!�^�k�LÕ0>{N�'NMŶ�jdUv",R�Q�w������U6y�Et�p6��Lu�K�nʅ&Z���.�Z��pu�uެh��9�d�o]�6��Z�1���ڧ\��ˊ����K�f��e�)���f�! f<�v��nZ�·������x���B�S�� F�`����j�_R�hL�$�,�XJ,��xqf�-|v�u7����S6�!M�q���ƅ�]��}��T�n=�� o�j`���ݻl�O��]6���``;(Է��CJ,��V�w?�n���j7�~�o���x7h��H�3Q�N��ɉ�����KU�>�n5���٢L�s�EVAs9���8��\���T4�:�s��*��Z�b��Y�. �����ܹ�F��SJ����"\Js�kąt2@��2�ZZ%�[17�71@�J�E輒�i%�w*p]`���C�����\��`D��Ƥ]ל�m�Eˬ�����+\j��v��۬��RXX���f1�y[ν���\<�ve���]����1%kt;gP�l3�G1ЫU6�<ޑZU�:���#F��}�z������ FJ�6�]��Ѹ�t+����f�opg4��,s��FYN
�rա0����gz!����M���WtL]�
�O5�u��˕�u���h�=1�t�r�-��B��Cj'$��� ���u�+Y�N������껮�QV��ԺPھ�E� Kz�u���*/qu�Kf:�Q�b��_gh���%S&<�=��5�@��E7�=�C�M�6��5Q��}`�of��s�֭�ٱ��������:��S�S��&ew�^�E�+�)���&Ū� ��hYg��Go��
�$�^�=)�
�k@XK�u�}�)F�E�y}�F��[K>���h��'`�ڽS�]A�ݮO�����)r�d͎�IV!�h���{ğ`/�.��T����&��&�)/���aE$No=�r_E��%VWT!@b�3���2�wH����x�^�:������re�u��T8�h��xM���.�\��YpU�e��W>K���3/��	F]
	N���w;�I���KFo�8����|;b�e*1_G��or����*��x�n\�
O]��}ـ���uOi���r>�j�
���\J��.�#�p��ؘ�rJ���H��1ǝm�V���Φ�4����v�-��a��=\i�/Y9ҵ���24��Mn㙝�FC���V�ѹ�v&�3�K��Һ�+ �|�%˳:8����m��4 h������ږd\��m���]ECƌl����ʒz�H����{�r�py���oS�ZN�����@&�Õ���.�f��j��A�>x�K&�����K��_d���-jۈ;�RS�n�JĨ:Κ���8h������x�_@��*� w�2��Ԩ"�徭��EID���sM��5�Rͳ%E�T��έ�]�/l�ZW�wL�'V�ʢ2�cC�t�;�m�@L����J���/o+!�ؚ��k��<-֊#��ɷ�a��:tN�ъ7��6��ɚy�b���Nm�v���
r��ɀ�ķWr��`��l>y>��:��FIt��w%��Q`��Ԑ<���J���̾���l[�2�x���r�FeL�+ �9�1�Ê�<=b���4/p�CR�o��]�[j�4V�4�}nP���zR�PX�L`��v�
j��2l��4*�wt�]���z4�6LX�u\���|�uŊ���BEj���I�}T-p��C�l�Z�,��u��Ҷ�0C*��;��W�cu�y`
���C˙�-=�B��U����凭���4,GH�Kvd�ru��bl�ս���b��"�Ҿ�|eY�l��.��!Y�]�#{	��b7��d��h$����b駚��f%D�d�`��5�P���R�X,��O��kKr)l��]�g;�-J+��v�L��{N3m��DQ"�Q0m6�t�����
r����r�C*\܁��k�s����,��-'x�b���S2jiǰ��w�iiQ�{K�˓�L����ԣ2ގ�Bd����R�].G�5V�`�B��XkkU]Zj�DT�E{[6:��U�(Kh�n��Ch^*e8)���l�<I�j�vx[{�u����}�#:V�P[�J�qa���놞�� �V�o�K6f�v����%��C���U�@1�ˉ�%;��k�a�aē7X-ڡh�v*}�s����ep��6e�z�� 2HhF�W�v
/,��j��dL����?��g����|�a�Ѣ��ڳ��;K)	wvmR�6>i�|v���upQ��X�Qf�r�[A�^V�d&5M5\�=�����X��K0���0�ɹ\��v���u{���[6�J\��oi��yD0���oJ���]K�w��T��s���F9�,D���B^��Yٳs��}t�h�ϝ$;9B�hR�	�4N�����1���c��ieƒ�np�n�n�!���X=Һ�e��N��*rQ�8�C:����i]���<��j'�����I����S]()������s�}���� �f�}�a��s�PPQΛ=c*D2��,�p1PP#,��ʽ��p���1SV����+r�S�K��'v�\�3Fa���T2�K�q�r��Y�:G�
�x���-�V���#S��{wJYO':�
�Ђ]�J�����m�\&fև��v���4J
��fn��vr�0�+>W����9�\�j�
�,��v��\J٧i��n�TD90�gF�G<��sQ-z��J�{�Žp�X�����$�3��mw]�h$/P�y���.�<a�^c����Y�� NH9��G-�D�Ci=�9���"\� gl�A�%+m�w(,U��N�3�fh�fQx4x�Q�9`���t��)��@r�H���)�EH-���*�#��M`{{P�����v]i�Ա,]ɪq���������n����,L��-����c�)������M@][�	Df5)`U3�γAĭ�KDy�MՔ��;�1��[t�CUY&O�4��I��"/w%��
��+)����B睋v�.L`}-��n�,4
Ķ��/@)ZU�fwRZ��ͬi���G;w����u�MEu=��ސz#�m1u]ܫ���耴T����.�Yx�Gi;�i���U0�i�oX�t
�����k�d��������qL�{2	O����g��pH-"��8n���(��͠���;t��ڣ�n�Z�}�p�D2I�0]։��t���v�AX��6�Tk�}Y����7*6~�%���2�Z�,�Q��V�ۺg�e_U�t�K���!�.�H�%�:�Ѣ1� �V}@�}�7�	���1��yb��!kI0Y�6���{�N���:��V�@L���-S�J՞��a�ُ�N/'2�Z�W�JF���\P�Y[vk���;�� ��\�[�S�ކ��_X6�(-�\&!c�R�-:m[�c�g+�������t��p��0]�܋���]x�2��8wgF%�T���\�ױAt�R�r]�Ow�[\��o%�a\l�ɤ;�]L�W��l�b,�V�	�|���o]k��?硄^}dn��+�kX�Ȼ���
�y��t;d��Me���6�Ae�z��څ�%� B4�Yy��\!vЗ�#�n�U}@����Y�n1��c�_R�+Յ�e�ϭ��7�1��ܩ���e��6�����\�.�cp��^է;�����R�|�^ӊ��1�S��zhYH�k�Xl�uGD��Y�S6h���]����T$P=q^�E^
R��������� ̧�GvN�D��˂��ѽ`���Pf��l< 7�:Ї+Xa���J�#9��	7Gb�
��%i��1�,��l�{�GQ���Ȍ�;4)h��=;�bn���*\"����ߖr��dt�v����=;�wP�X���R��W|xC��hAF�ps���>B�i�.�6]��S�2"2�%�j�%$� �o��]wz�_Am Ϸ��h�J@���Mb\�P�3 $oi��+9d9�"NwM�F�Ʀ�����r��5��E�.�i\��YQL��S��_wn��e��/�k5mZ���sji�Nc3�ч�s5RY9
}QM�#Ъ҅>̒��5%�xƶ4��h�f�H��I`�˭��{�cS������<��QB���*���vjfb�D�oJ�C%u �n����Q���E9o+�,��䙽/&�{�n�	��B�B�@pÊ>ŖF�@�<\pVX��H��WS�h��jc������WH��Yʖ9`x���B���������,��k���֮'���'r�ѱ��^���"�u�#dQ�u6o s)�sv��i�o�V�~�H�#6�*:����)��w��ؒ�(	%�^<у�+���ݍ��q��ԫ8ٰ���eW1�"�^���I9�憞��X+mȝK�lf3����X�뜆�}�ַa������ƶY�{+e�-`:7uk���<�/�]7�G��t+���ٺ�S�*k��Ĉ�U9B����n�n�Hm�'�V�X�YJ�vU����.��,|�m�\C����5��
o�����8^�r�s�}�w����TU�bʒ���lԝ�=�FV��N�!E��Z��&�=��T_c&:"ѫ2��+�&����G>�r�<�.��l��"��c��a�oK1���t{U�tc6)v]�t�l[�T:Mҫ*��]΁��;9ξ�՚f��v����r4c��G1�,�U�� 4f��1oe����,�eee�/A�N��r�����$ŋo���D�f.g�c~�k�B�7��͈�7��ˊ�=�â���i%�05Q#P�Ⱥݠ�)V$U����e')���n�0��ñ��7���^5�Ué�'Y��L�E�z֛t	u.u�a�fb�p5I
T��L<��I�֌U��/,[
�+�@�������R��oU��-������C�H�Vs�������8��
l{oEՇ(w4��%���4"ݭ[C�j���0v�W�gt\_׳{�
�������Ӿ`��G^GinQ��N�m)��	���HK����cbO@u� �q[mtC̭�����>�r�;T�Ur��>8VLG�R��'|��c��ZVvN��V�ᚳ9���|4>V��@o��Bk�v3�P�yM�u���Z~f�,p�rԶݮ��HW
O�����Wj�h��[9}]S���n>�H�# �wg�����#Q���1�Nt���;q��QaDT��b���@u	�����2�1���_=A�Zzu��ںP���e_E�9Y�MU�ZR��]0�a��m������t��/�-9�;�P��-�E���
F�kyu 2�KKN�������KY��Ǹ�ή�U�n Gl�M��xw\Vu�R�T�ڝ�]�W7���'«T�jܗ�/�\�����sOR�y���)�:����X�����J�$���B�i����%vMښ.+���V|zE����Hm�.�r�ڐ:��\�>S�3zՇ�N1|M�Yت��#שf��ު[ 5w�괯���S{���h��;[2ɢ2��t�i����.�0�{\�
Ղ �M�"]�+!�W4[�-�Y(��9�K���ʚ�^X��U�D�`�O���ܷ[3M��淧HI�tsxJo.��]Ӎť�eַ�21ßG�F]�B�̺H�cB�n��v����R/h�(�2��\��irZ(\��d�*s�]����MiN&���ӣ�ݺ��������qe����]`�i�r�Pf��;����jjAk2�[�[��r���Ԟ�K_*��#|�w$��R�]��!�����3��urS!��X�X-��Z�6��@�+6uL:Uʲ��p!]K�ٵ��6=��]�0p�D�щvA��s3fu$���#�z�Ӳ�	_m�����k��e���WCM��ëlR�v�nT��a���n��k V��R��HJ�I�٬��!�sϖ��h��jfTw2�5����6�'���d�:��du��QE��
ą�de�d��w�5ݧF^�|�XZ�J�k���8�k�s
� �|�J�n����Q2�n첷k���{g2��_I�l���W}@d����z`��첑�����`�@� w9t�:���Z�u�6o*>HI�*��Z�ʵ�%��u�9��K�i��k^,���X�L�L�ƱBj,,\�)WG+ImXIO���b��9�����,��s��λ��o+I�#ʷ��' �o{��
�׏�!�;�U��b�82�MwaxQA	�'s�S��A��j���e�����DVp�M��o��)��"duЩ]�c�2�cF����ֵ�TO�z��8��s����Fs���S�����SC��G���>}`���Ɔ�B�K%�nTE��@ùx�4=��]��e�eqUW�fV$zs��P������$۳Y�[��,�����I�d'Ã���Jk�2�
N,5M��Z,k��=ZW8�>§8�t\6�T�RϘ�Z<��6���h?D�j���G%<��ͨD�{N��a[�;9fU�����N	{D���]<�z�.0:U9XW�E*�u(�#�j�R7���b��n��ݾ:kNfuZ���0
�è;�l������[F���r�6yu.ܝtV:��qZ��H2�8qo"Ke8��l?X��3za�"a#}]nu=E]��
V�m�����Ѳ1�ڕ�,ݞۏv]Hl�7�/�t&(�ļ|�l0����o*�e,U8�06eն���JC%N�C{���}JR��Nk�)X2Sw�軺� 9���݌ʎ��ھ=��J�NW<Q֑wnZ�k,6�L���>��T��ͻ\��+�RYǍ���Uu�6�}�&ۉ�:1�����1$�y�\(ˎcH���NsP�4���w/��"R�nJ6[XdC�4�p֧e'f�£�ʗ\�;&V�W�{�>Yg�u&/8[Een�T�=���7�t}�c��VE��O<x����.<�j���W��ޕ!]m�ʰX�b��B2橩����k�>w�]�Y:K9�5r\wy�Z�����W�1�J�2��)K��>bM!��Nk�g��]��Y�jf���^��ݨ+21�)�.��:7u�P�0��{����~���k��kEݣ��MDU��m	r�6���[ss���5��cb J(�2�Nd��Z���&M�w4b�k��L���bܮ�D�h����e�\�"��b�AGv�ccY�3Ad���)4Q#1��t1����E`���M���a�a��.sE�hơwW+�ni���[h�$j�����*7+�1�܈������E��6*ĚM�c�ch�$���b��TZ1m�h�lS*1�T	�Ԙ�cP���QAX�lTX�lV"+Q�#F����Q���5%��5ͮh�*
�B�︻(��;]3S��j[�ɽJ�N3%�(g9�mj��qK���k���Sy��uo��V�*oے�vXz���2���\�!�.!�-F��#0�8��l�f�Zv�E*��*�u��M<�9WqE���z<8�W7}<�˸������:�=��]Q��טc=���R���v,�����֧8��r��뫺�K��������#&k`ׅhTb�Z��/;)��p�t�|��z�/�u�;���L>1p��p�Z��ډ�ŉF�\�c+�t�2p#�����{No7�s[4~q*x���`M#�W�Wn뿌�l�U����x�(�Q�(@|�9�/d@u9����1���xM�ÕҁX��q����Q����G<�	�tlU�;{�i��+*�p�ۃ?X�'D ��R�h� ����75���Q1Q��vz�5ӕ�9پ�s?j�gn*9 P��P3��$v��#/WF�Q�z���� uw��Ԯ?!���b�����zݼ��CA'r��k��!�c�i�湻��|n�붙�T:/�*X\r��ӑ��6�W\)�e�6
<��D��L�c)X�зձ��]V�JS��vnS�3����t(��C�J�L&�����\��;"�z	�Ή{sjͮ�%j+5!���j��g2�Kr�V5�������Mj�f�@�;��ow��G�(� -wL�o�S-�8bHY���|*�V���I�X�`*�M�Ê����s���/��H�s���q�*!��!�i�,�Р��t訠�c�����������@@� 2�y�`(E�6R��·<7��m븝2%�׼�t����Q㙇�+�0t�"m@�4LAJ�05wm�rj�P^W3�,���h�ލY��%����la�Dp�~�����0���F{��g���ˠ��U���N�^&B����J�9�^.���kZ1�L7'����5��p��|{��{N3+a^v�Zi-�0D2^{t��loޫ�8�IJdѶ������yՇ]8nX����ʞ���3k�����p�E�g��E=���������p'7��ێt4���:,��Ne�;�>��[$���*���^����X|-զ B�ާ��"�L!;7qZn͹â���_��EZ��큞��*��7��.5�2Pcw.�~�O��dD���*hMm�'�r�Jv:W��եO���6����r���:�����S
fa�!�63�L��c�l��b��a{�}yCۃ���r�-Z�ie��&�4���QѮ��U���PPY�	�z�-�c��=���9,��4P3+{vVo7�Uz!���W#�E�$޻N��@��q5a	�Ds�Ř�Xk��V[���E�����4��!��2�@ö��>a7-:�<;�c��X[����T�r�eyk�G�Z5��XyQUo�X5�!�*ZͥGMsסF:͍Hv"���22!U|��)b7m��+窶O���+�P�:�L��mA��\�9r��8��K�v3m��T
�ȖU�岝*�z>(_NP�f뤃�e�qx��9��������<q�Lz�ע6�T�2!tit������ڄ����Mb?\i�'^+�{uЦo��8�$�@�g��L���,�B�K-�/�O��q��Z��ߣP��\����k�g�-��,����f6 J@�.R2O�{Η|��h����P��`�dF�(���J�Z\Bق2�M%9�s�" O��
U�)�����K{����9�*2/�Wj���W6m܍�ub)�%�WN��3�ZX����å�O
J�N�Y�b�1��K���\�b˛D�f�
�n���t�Ԉ�1��w̋�&�[��.���\�	`�1Q�3_guHh�1˝x�/�(P@o(���r1��"6(.������W�²V2(,u�+�/s�f���"^%Gx`��x9�1t݄ �<���n�cA�XJ��t����k����
��V�Ҝv�'�uJ��wQo2=r튀���n�G����qm�q:�i��rO�w�}GOl���3�/�pX'����+�V�f�!���b����g�� wg��Anj
 ������X���Vuu�(�Wm��\�̦xW�2�vP���X��C4�I4q�C<���c������Z�ؘ���g�'r���Fb�Qz�|�X������s'���X�ܩ�7/9 �u��.#��!�,Vsy~��hL]kQ��Q��+K�c6gNF�z�w�-�b@��Q�On*��@��#НW�q��*�h�Y'\�?t�T�Ń�����L�'�4�<C�h`n*��t��`d*v�[�������s�x���b���3�#���8%>LS�\��S���=(|��¯�6y��z��_�9b�*b�lR���)m��J5b�����~?w��RK��U�ڠ�ϴ�x2#\L1��:a�a�0Ot\>�G��b�r��1G���r������'3�";���_)���t"?/������3tg�;~G0麷Vc薔�F1��[ԇ9���4JQ
@���<�<"H�♽v�\LO�)|zA2��6 �l�J�U:j�7B��P��Ҿ�G]-�h��SM����]R�v���:�����y������t5��m)0P�\�S�;�'2�2�ҹ����y�t�&gG+xǫv=���[:c͗Nn���s�Ǯ���v���x�F\S�EdC3��u����w:
�h�{�qf��GsZ�*����F���C��ޗ�3#�:�����2-UT�jƒ��|v�U�Q���[�]���&#�^C�:t|���ϋj�8LZ&�w�N�_�.śl��ԏ*|�Kܞ�."�#vP@V�F}L�N�p��8Wg���n����5���9끔�)�����mr�X�����(��҉�2��O���Lׅ�U¯3�8]ws����77 �s��u�Z����4�Fhe�q��:�=C�i�8��z�g���Xj�+@��z���J�Gp�K,Bo]ޜ�s�<����X���3�bR|| ���eZϻsڭt��U��6�Оg�_d�I��F�//���.��e����AWyT���պ5��fު=�C.w���Nu8���J�'.2P��!38>��Qo��K�n_i�3���._۵|����p�=�UaW·T�kӖ�(	��|�i��Q��ۤ56��iX�(�iޞ��ʬd-��u�8���kJF� B�po?�c���V���8^r��y_f-�E24H橇�-�7���k����˖�U<�o��&��i��ꄗθ2~�6z�Ώ�Kֈ���X�h���U�À��:�{r��A�1XP$y��Ӟ.����_n����l��W�*'k�ഷ�m���*"�*M�W*;w�WɌ��[��T�K��{�nک�������G �����|D>8!@�V̰�n��:
�q�6�7�����54�1r�1�eh�����Hh$�RX{Uu�����Z�7�Q��ڧ)�Ct�����v��9�9~C[Ur��^i��i:�C*���ͥ3��xِP7ܪ|��3RU�c�s�i�#OY�?eCuC���T���*1���
4	� @� ս���|�!vϧ�[��']���]�鎣+]�s��=�5��v~��GK�({�@`T{�L`j��ڎۀ�MZ�s1bsY��	�!p��N�'��N�XD�Yՠ\*ǑVdHC� ��#HNz�E�v�,*�hZ0�b!<���k�y��M�h�0���U[���D.4q|;�����g� YvcPs5����f�'Wq<b�K�$lr�ɢې5�6�W������^�/��ɴ��:��#Q�����r����s.�	E�Cns�t�,$��k���4d�"�D��2���u�6��r�^�s��^��{Iޔ��33!O�9ԏs��(c��w^�+�?[��̄�uJ�' ]����8�ì_u���D{p͋S�]���z��U饑����I�Q����ɯ��v���r0��~��;S�"��&���ͮa4+�Ğ���3]f�~W�R���� �>�~܌�΀�_<�Bv�n��|����;Ǖ��="��C�-���uq�_m�^ƫ�k���(1�n]B
8)z����1�8�mضI�	�'���ŭ�����.�V�t#־,�����*�ߵ�+�s%�v�������8��[{]t~�[,����� ��9*/�۬H�|L�L9ʣ�^.�y��]fN@�K LB�\�ϕW�m�)b7n�����-4��K�w�v��,y5m�O[���Mdå h�a�،*�Q�K*��-��;W�\/�Br�K7�A�U�R��g��'��i��E0dC;Z&K�<�hB�叻:c0��O�z*��\>O��°��9�V�����a�O�� wOҮ%�}ӥ�
,X4%��G,N涹»w���92�e�=�.0�U���T���.���F�~�S��IJ��7ᘵ�$���d'⇶�����'�0B%b9�#&�I�=��N2Si	��v���ǭ�z��af����Qۊ��r�e6-7�Nu�&lL��>ڕ|����ʆ�=7\�95j���݇hlv.���N����r��!�{���s�Ѡ݆��Z{՛}�[�>�g^�}��	;.���e9���uR�  C~h	Lҙ�/+��x��d�e�c�n%��	��8\������Cn�mӫiLI(TuI] �3�5��A	��[5kT�����:�D�a�ܺ�!��k���.�~�'�t�Ԉ�^i�yny���KPˋ��t�	�Y���Y�R&*9'e��E�&*'C��#���@���{�z�u�괾�CM{X���Va���1i+���}� {M!C=qBv��}�)��/���*HBˣ'#����Tq�ޡ�p�#H�.{M��\9��c�&=�+��j����?p��g�'r���a�u�謧�D`���\�L$���ѯ���V��L�����b�{T�n{ݚ-�*���0��Q�c����u�������AMyEs/�m��U�f�����ځ,�6�W�x�����N%�of�Wv��;�G(B�9���Q��J��>�u���N�+~5f7n���	�ռ�f���a�gA,��jk��I�L�5�A��msw{�.J�*��+9�����W�R��bӉ���k�t��>f򹛭g�;��NSѡ�F����%6�d�Kc��}Ш����1VsD,�u˖:;�3,������Ϗ_"���[��_Q��h��g]4 ���4hU v)L��l�����W5���ݩ}ј퍋�^���h
�~�(�|#K�gϐ�mPAhn�c�X'�[�f�SF�z9�-]KBN)_�M�++�ρ�Q�G�<�_����X�b��Y_U]\��(Y���e��m���Zm�R���w���U)���@��|H�9�3ԫ�s���z�����{3�3��\r5����sH�fp�8��d;@��9�̔Nlr��@p6P��Oc����ޗ�>NcD<j���<P�͵�[4ww�`��O���lo:7� K�^��t���:�t|��N�C>-�,�1h�m����g�qF���l�G{.������ejD{�@Q�8�LNd��!�s��sľ���Jc�,c;jR��7�DX����So��$�N���׌�^][��=s�vf���!���ڶJU��XH�E7,-"��.0���P��Ƣ͇<��g̬���a�#�=���d/C��4�}gV�/����\��u)�}u�Ѫ'.�j,܍�DJ鍂ݤ�y��'k�V+�b���)n[6X��gQ�q\#p��Q弇@6�]�M�Eo3p,���0��u�7���Y�R�(��q����9s{�Fνȹ('����͈�����N.t�xP5�^�b�y�JC�hF.V~��S�����":���!m��C�O�h��}0�����s9���϶�D�1bQ���������:kWӨ:w�������D��9��F[�2!UV��9�T>��w�:��FU�#k!-9����q#>=�i�.��n�N'f|�x���4}M<���5�O
�s6�>��Ӎt{����Zؠ=���أd����8+G�t���}��L_6Sy�q����-��=�oR�k)�U�F����R���p��'t�8�BH�*��L<�̒���b΍yr�;��8�z�TF�NӸlÕ,g}+/���]F.(�$�}3�L�
i�!ю��ڷ���2,C��3q�%���;zr9�e����ڨc�L�/>�8
7	IF횃�b����;o�oz����`��/Ꙏf⒯��/��H�9z�����!̌�=]0OVmu�W��G:�/`���� i��P��8*ď~�U��K}�l������A��{R;71��ɉR���PQ{��퀩WY��ɸ��Y
��+-H�p���}
7�SuY�y��T5ݻ�L0�8��ҟ-��0lx��vXUni��k%,t��d�r���Z��[xT"�u���Ѭߴ:�Ѣd�$�O���f�Ʒ�}Q�l�Q���
�ht�WH��+s�4�ۼL�yA'�6��օ��I �
u�]X+
�Ӌ���#�+�p�fk�w;��#�9��{�%p���9�rr]]`���z�$�v\r�,�����wv?m�.������{lL�	�`P}x{t�8� ���}���F�p�g��2n
�j�k���n�88��ν�
�Nk�[��� �k�q������v!�[��#�O&f�ރ��t���e�s��t�rqSfb3��nRa8�Y��/��sD�^��x$U�)+P����4:�pV���G��f΍�5�XJ�T�Yr�-�[Ϟp3)�c'�$|s����y�>rb�m���L�V��Cʿ�� ҪgM�@��^'}FS�C��M
[�IO���.�� �G8*��h�V�Ō�-�)Me*t��ދ�����`��tʵՆ�h3K+4m7��iV�s�h,]����	��@(iJ�Jw �vXr�1؛���a��k�ku�۳���y�1L$lg@�ݙ�)1�)'�(`��ǒ�a\��D�����p[X��A$Ov�-sT�zr���<jP����g%_��)��:��T,.��y�	ok���M�Ԕ���\l���9R�i�X&.Mp�ܡ��W��]s��0/h��Xo;,D�s缬�Z����J�p+��v_l�Y�s\I����f�o�^^�ǌn6�MZ�}Mf�'�R�H S����0`�ܓ+_h�E�Rpe����È�b+57������-������ں�S���n������p�`*���K�S��5�K�@ǔ�O~}�oZu%ٜ/J录ϸ��n�mu�n�.
77���`6Os���1���w�33@Dm^5�\�W��-=6Nm�Z��z�u�᜙dU�T��5%�zƺ�zƊQ]f�u�Ч���p-��͋(�;�`}L*FI\Ml0#��wuѝ|w�ήiʹ�cz�!�e���o@Wf[{˖m�:��ӪܘQ�M�j�t���}f�����iVz��XrE���Q.�Ǌ�����v��6�9��ǵ*d�ou�s8�p�g3m�j�(m�+N����X�ד4_l���}(71t�p�2|�4�U� �����Wtu�F�%�r�]����nu"��iΛh��S����mK�0�����K����v�m��T���'���ez/��`'��$��j�Z��`��7l��yt}�7i�>\��z�	��v- �_,�x\�52p^�\�U��W�.�ܱ�}j�]���O��ņ��V��`����M2T�Ee�+m���,���⫫�{�Ãy{* >���
�@P��R��5��ԕ�(6�i5Z
,ZBأTQ�X�Ѫ�*�X��N��6�S��m�5�c,j-F�6��-�nTX�[Ʈ��kAQb6��p+���I��#[�㚃V�W5��U�\�$	���F�F�W�sy�3ch�Qk���,Z1cX��r�V�m���lE%�-�h���h�o�66LTkF���[h�F�\����K���br�N��8�s�ڷx:9�ݙ��K�Җ�h8��wƈ�)s焪�!���]���� �ӕK���;�?�;�����g�潷��h/w���zEx��ž+��77����Ү\������m�W.W��[�~��o������_������snU�r�|��o���ە��}{�~���vp��.�Z���}b,1��"@���rߪ��o���}�����ݿ7�~W���Z7��y��w�۟*���s�����ߝ���_��Ϟ_Z�����[��W��5��-�~�ޖ�}[�����`x��6�6�7�p��[��|#�^X��6�ϝ�zo�n�ž�|�گ����y���y�E�U˛�߾W���Z��_=v������i�v��u�{��^��^�����}[��^��~^|���bjBt�]L�D��d��`�=�o�j��o�����\����?�W��+����<���^/�x���|����5����}��{U��\����0��\�7����j�[��������*� ��H8=�>�ɛV�^Dc����>���}�����m�o��o�=-������o׍_�ߞ���Z7ƿo�>���okţ���׭���ҼowϾm��lnoO�����_���m�_���=��or�E
��iF�'++TUa�wln��u��KO��/�mʿ�K�����m���[���m�x+��-�\�m���~���\�w��������V��|���o}�s���|�B��[��������2K�-��]ٽs�c����|��_���W����yoM�Ƽ_�{���zZ�׻���_��i���^�>���+�wW���ۼ���{���_7��������Qo���y���q����A�����Þ����ky����ߏ�_o��/M�������k��o�{{_�ڽ�ߝo��^����������Ѿ+��{�:���{Z��W�~�������[�^?���@1�1�0�LfU͆"Yu��a������o�_+��ז�|�\�>�=y�����o�������6���t�?������͹�����{�v�����μ[��x����=v�M�o׍�ν7�{Z7�~W��"��c�#�i덢Ⱥ�4���n������~����W���j��lno���Ͼ��\�����鿾��*���ߞւ�ۿ�|��i�����|���6����>/k�����m߿�U��<m�� T���t b������Xl�P���sTx;��F;�k����S�����c���{����E�-���>���p�B�	�w^��^����K�YoTÊj�6�X�#�n�>5�т�GF����P�A�1Ϲ�����W��{k��%s��<p[��}��;���}}���f*��y�zZ?=��������|�j�忿��|�^֝ڽ�?�z�_Z�|[���}��M�}k��~￞W���W�~o>y����j�_>���W,z_[x���ׯ`O�=���j�5ǫ}H���>�O�B�[�wo_�z�|����ך�-�-�����_����^���4_���~o�h��߫�|����|W�y�������ϸ�7	�Ii~�Nc;�>��p�+��W�<��r�U�����[�x�}W��ޕ�5�z�<���x����x���\���+ҿ���������W��r�k���m���s���5�����x�����'��GW��pavw��0>1�D�� >R!����߯���+�ţ}wW��׍�x���EDW��޷��i���ם��oj�r������m�o��ޗ��~��u���ݾ��i�������y����}�??>���������ۚ���7��������}����?Ϳ������^��\�^��潯>u�oM���������*��׍ͻ�n|\�ݨ��r��:��	��	�����D!X4��-��\�ļ�%��X��#���L��C�qh��>}�oo�|W��o>��~�r��񷟷�}U����n����>��U�s������ֹo��z^�x��Z��������B��'�|G�Я�}�L���Vf|�p���q���D�£�c������[�{��W��_������\�Z7�{��zߍ���Ʈ��-��[�|�}�_�o��x��~�潪�\�/~������*������{[��W7�_����y�6�y���X�0@��p����*��דo���?{������o��-�[���W�:�7ſ/���s^���h���ƾ�mx�W��oFc�g��?|dk������oǿ_ߟ�����*������oM���x������h���]���[�^-=����6�7�no��k�����x����h����o���/kE���>y����Z��|�שּ?|�@P>�P�	N_EE\{]x5��߿k��ͻ�n{}�y祣W���i���i�_�{_�m��׋���w���o������^-�u�oOֿU�_���ήX���~������m��;߯�}�b���|z��cb�{� u8;���2���M>)���o]��^u3�-3���P��8����=��7[��lR�2�O�Q��/%+͆�k����!9>Z{uDRk��޷+ku����W#�$��!�ے��]�
SK�V50*;ϖ��N�4�M��}se|��Z�)����W߾�Q#�#�о}�^�6���U������/�z�����5zom�o~y]�׶�5�^���+�ܼ^+��u���Z�����~^u�W�{Z7��߭��^6���x5��_h�2Ǆ����U����Q
{�}�>b�_w���_�ߊ��k��ׯZ�}~��W��Ͼ�j��ڻ�}�z��{Wջ������~7�n[�����{�znoֿ/�^�r�;o���皼[�<W�:�W�޵��>�����9&�*׸5�1�X�������x׍�^/���_��y��i���{��{o�żU˿sכ}o���~o�|���h/����������_��˿:�m������^/~<}} ��(ٚ51o�}��� ��ƾ�_���[��޻����Z�羾6�ݷ�������[wv����߯��AW����^�����Ӻ���;���׋��=���F�/�����~/���Ť�њD���	������s���@�+����~ur��}^�;^�.oƽ���]�ͼU�s�{��o^�����o����ǟ�o���6��o���z�Z76���<��޼k�\7�������xc�w晡�_N\f+�;�����1��_�+�_W�E���>+�ߍ���_��k��W-����Z|�+����oJ�.oKƼ__ͼk�{��zW-������KzW+����Ͼ�����>�*�^���(F$���.w�D��no����^�.��/���?��[������u�o����~��������k��^7�-�^����^->v����7�żU�{������������n��x�Ve?q���`}���z�����_�W���o�5�~�����/��������oj�.7�]_���[������m���j��wm���/s�wun���r�_6/pb�F�~{����0>� L�����W׍�_�x��}�߫�ѽ/<����^*�|��7չ��y����׮����}���o�^�7�~o|���6�DC�������pB."��yu���	Ne@�aqb.-=�t>���7����4S�Q9qN�l�Ż6W��	�Jhu,�k^�St:�u���Gs��A�L�ݜ���m%��[�C�i;9���8�P���-,Wi�����\7w.��'��*8k��kZ]��L��ʯ��'�yd�t�S����$,�;�Ǒ�n�4xh�&I��u�2��� +���<�f�M���R١t��v���W'h!�[VY�b�2��U4p�����k��1�~�K���r�"=����<��{'�����\�~6��Z�T�mZh����ݷ��io��(��'�鏩M�F�'���);���Ȏ����4؝`s9�Z�R�Y6������X"�������.0��uJ����h<���ҮY5�s����k@^��h�4�	�v�r���B�P� �ߛ�q�1)��|b���Iʕ�v[������Ջe�������E��+���[�+��0�ŉFҞ����BϷ��	��ce5|~t�����f[�3�UZ>�N��}4�U���S���ZS�-<��u�8Շ
��'���2�k�)`��(	�W������U�o���Aޮ{�(g\� �}�H'���L�l|o�l��W�*8�Y�Z]>�_�i�>D�W9��Gn�oB�mqŧI�����s��7�ko�ƽJ2���N$��_!$v+�䍨�Q��̺�-0n���^�W��Ffc�����α��+"��|�[W����e�ʙ�&�cQ��n3��w�8�co�{] H�h���-A� �,,=YsE%�x9����\��{�o�J}˹�����G�K�`���H���">�-�y7R�\��YT�dqt�O��lÕ,gB���<f��I��,������I����ݺ�魋u28EI���1(�}��Ӝ�2�������e��gF��}�5e@�v�;8�`�QA��023�+U���"��z�#��F���#hd2=��66��}]�;Sb����t� 7��p[�N�
������wl���KMd��Vg���g�ӣ�n��{��t�Q�~L�gb��)P��{* B�����Ch��B��v\�a�c_6�@�u�"�!�� \@Bs�d-9��7�+
��7m%��튎��*�%7<_3X"ь��*�u1q �\h���r��s��4ط�x8�﩯q�fi��+ꄺ�W)L�6۠9�5�WO�9���+w�ޮ��;�ճ܅j�� K��R�;U���v\���H�O���"���J�F04lǗ��˓ff��1@�����5{�]fç��jV�2�&��7���.t�����;�ڊU��x�Z욡�V��c(�t��׉�P�ޒ!�W۝��>;N��ie-��c<Q��ړ.Ώm���Ohw��篞s��ik����p�c?f�X�+������1)���Z]É*���.W(0u��{S3)u�`W�gf��^����>��ga���z��'��kX?NL�
{,���V���L!`��n]BïodG7W+"Cqy9��8���zV����N��{_Rw����a9���.��ΩEa�;�wWl�mu�ض�����i�
���)�5t���5��Q�+h��8N#�_{Rw��K.�@����t�� kK���ap:�	D�<��U_!���ݶ�����O��$�|�
�ֽ�0v��	���-�K�3괫�daU�"YTm�l��j��(_;,u��p'��Q�T؉��d���� Ȅ	��R�N|�hB�.������,]g�Sr��F���/t�G2��<�g�؄x���.|P�a�fxs�X�E�R�	�L*��p&n�v{��"�-1��8�����p���Q�G)��(*���t|��i}c�K��2��U�Z��w;]�;�.
�|wa:x�ق09(N'U.m BG�S��ź�h��5͸�N,*���k���NR(���l�H���SJ�%j�C�Ɯ^,����,m�	X��kBǩm�kB����zR�{�X�,0��{�z���z�ۙz��]�J.=i	�n�ڝ�U���uBl�(Y��T�.)�3���t��}ES�ٴ�Vc�7�{kQ����d�4umZ��b�+�:�0[$*���W+G���$:���1nmer��d�gT�Ō��*����5������fFu9۹!J�Ô��q�s�������c��U����lӫ=㹨��Z4�vY��#��֦�[��O�+ZsS�ee{�[@y������CN�c����i�WZ�����w�k=�������ݾՙI�q�( ���Tk�����D`���PD|�=�����޵e��Sxw�7�۬���e�-)�k��Yb���nhED42�EF��@6 ��l����1�4N��
s�}1�<,Hqe�Qy{|0L���:��LV���P�TH��@1D�8���r6:)˃�,�뺯��\�իu����0X�w��gT�"	gQ�N��U��b�ƌQQW�h���������a&N�b�O��6%>Cڦ_=:��4.��6V����]S�L\�:�j���c&��U���υA[��G@�<�t�;,�=������>`�;q�f��Շއ��z����2����*�UQ�����4��|�\��lp���}�=�`�eIӷV.�7܆WnQXʆ�j�9Z��?��0�V	̫�P;w9Q��~����r��&���~c-v�D\1�M�M�R�0�s������зһp�:ϖ<t3J���i�WOOn����u��zv�\��P.ϧ��ꪯ�J�T>��\/�����x�����]pY�8
4�z�3>0�(�F�ӛa4kl��'3�����u�����b/U&r5�f6� ��ޤ;!����͒��9I�	-͘5�r�F�f��@�Ѩ�<S4�TO}(v�����g<w#.)բ��g#���C�ʽ4��cc�s \��r<"�B�1��Cϥ�l�A7���NcC�17TDY}��z�v��[�}�����+h�Z�T�&#�2�:>U��gŵe��tj��U����T�k��{�?V�>5��=�>Ԉ�O���.��4�Z�����8RQ���3�sz�Kp�S�%(�Ö��"����>F���Izx��TJ��7Q�2h\�������k����!÷��DrUtoሰEBr�����]Y��|�������P{*嬧7֢�F��Uy����z,��{��q9�Ck���\�F� #���ٛ����!�Zr��r�jΕ4�.B��O�;��A���֊?s+�Q�����{x��qR�»M>�"y*�zv+�{a�:-j�Bv�B�iݺ��B����7��7�Y鯜����t��T���u�kd���#��;-��sm��%YN�{�D&�(t�Q��ռ)A�w��T�g�+T��ͨ���d�Ȭ0i����-�yl���^BB���&��ѨZ��o��\���Z��o��UZ>���\�}���S�X=�c�#9�9�	_i��xg
�0�����q;2���!��ޚ�!9;�ǹ�)�9��8uQ��Cu�q�y\.3ݱ���E} �[(�-.� =��+�W��]p�Ԧ���°������)��u\4n5��c[t;"�<HH��z��ĊTz�'Uى��_mS#��*0��i�6a:TƬ;/�Ţ�D���+��R%|C/��e�JaI#8��#hģ5��<�e�z~Ci�p�&�k)ؾ�r%T^�b��x�� �'@�<|
JbI�g~V�鯊E��]�w��=17j\��WK/��Q�~ǝ\#�M�f�9�P� ][�N��*��<O�vϲ/	lt
+h��ͤ�s�T�F�u�M��q:dJ?&`������_A1���L-�72�����V_��8��\8�����n����K��h��P �28��4�N������Zwx�:�b��iEcsv��U���F�
x�]�����rʬZ�yk4m����*�=Q��:���%���{��!:���J�W��)i�{�z�;i������%;�f�_5����Sn�G;��pt��,��L�Nb���޳���+���b'��*�r�ri7\�k\B1�L7v��Un�,��v��:��րMINqd���֊���t,;��}IuH��JdѶ������MQ��r�����%��:Zb8�:+�
����R����������bN�_�g�&��uf�:��7��Wm�����4���;"L=��xpTR�f/JY4,!{�� �uw��_FN���攍�$V��8�#Z��rg��>r�$+�nW���b�Pc�m\6��V�����w�`(�.#�>s�M�7�=����.�dt�9���#ؾ�QX��,jGy�����~��U�'\L �}hgʪ���1�fWy�3�e�Z)��k3�ozx�^AAuk�0�u�C�u�y�xc5]����Qw�s#>U_!����pP�V��{d�"!C�\�h�<h�'�Й����U)�C�J�6Y�A��|y��Ked;W�\2��Q阑M��§Q�}S�^1� �+��P���m�o,Y4!\it���8t�?���ۧ��i4Z�3��xg.�\{%�Jf�1�o#�GAΨ�T�Ayf�VD�_�Nm��o0>���]�Q��-���Ŏ^&���:��8퉛�:Y�&�:��;{�E��e(j!�pe�V!����|��tM�5�yy@;g&<)��9���vmv��6�ӽ�]9 ���+��o���R��`���][�>�|��F���^Q�we��]`�֦<��o��U�=\$�.�ɉ�.t�ѷ����b�3�4l�c	�9WlX0��+��-c����"�k)�ZF�����2���h�r��\޴a������4�X��]>�z�sW=�T�u@�+b�%j�,:Ŏý���6h��"SIՀ2n�r����Uv'����s�(�ȹ�4��en$sj'���]u�A��}�}$�{�y��������S�Xim(��LˋKË�U�д�(:N�y|����:���p�BE���WWT��vp;8��
��rXm`�-��]S3n�O�1g���M��H�k��A���=���*ů]0��:%j��u��Q�Üb_e�U�oe���{�{&Q�0��)�s�ޫ�{�'b��,����Ucl��k+1��F�"�Q2�.�;U�y�`�d��]\�mJx`�nw^�G鮓i��Y��%����!ӗ���ʮ�_�*T8�ع��7.�]m1��P�{�TdʏuX�م�.����`�Z�LԊ���q�w-�i��1l���u\k[J�����;>�u*�
n�f��;n.������y���Ԯ�b�u�lL����U�>�=��9�ל�o(�<�]��/0�4೺c]8�h�]vյK(]>����V��	��}կ�b���囫��ɽ2�>���C�X��@��4�x�8Zp�5u�n�G2��D!�fϭM:w7���q�VS���<������`��#���ua�Ü��G��Ŷ47{M%M�/Fr�(����7g4�bK������wp0i��r��fM��� �����Q�����<���`;�uʡԴ�F�s���Y�GŽ�]�k�!�2Z"�v�Wk���{�w9��%�ӚΫ��m��q�ӓ�ea�U5]ӵ���}\��T��$!�� ����#�:��[�|M"� �n�I5N�����K|�`�x՞B�_8���J�VY�د"��6�Øc�ؒ���m��9�����7,	}�2�'Y�2���B_F;�j2i���	�r6���B�r�n�|��y����ܓ�IoV�P�a�Ƕ��}���y��Mb�s��	�ɘ4p��HmM'x�z@�_u���K�a��wd�{m����T����q��7���͵��NԨ%����X���:�v�[��(0�g�i8�fP�]������t���w[��m��Z&�"u�$�35;�J�:1����+�\�1n` �=]S>��)a�N�EJ^�K@�Zt3������������~�n������Q&�b�Eb64lj4E�&F"�%����K HA�(dlh�4X���JX�cEId�5�hōa6-�5K�t�l�ѱhƋTm�Ռ.�b��6LFɍ����m��(ƃlXэcDj�cEX��-���V#X�h��nW75X�#Ah6�F�c4QQclTj��5�mō�(�E��I���Dn\�������޿����(ۜU>�c<��qa���ugWh�'���8δ�t2i���!�:o<͈Ԯۋ*�ANk��O��}��_W���Bq|��,w��SZ��(B�I<�+ _�<#J�:Ih�_�}x��-E�|E�<p��j�-���r�sn����Q��r����	M�����83]�=��d�����\M���e]>;�������Bi:�sh�!VM	v���Fl��A٘ \�=Yaq[�_qN�!����p۹t���SJ3݊MwS�̽��X'j\���W�%�c0Ơf��SED1��.m���-P�"3Oz=.�D}�r�C�ۤ+�!����bF;V�v���)#7y+&zW:E�9{��v� ��R�v�d�o���'��rk�Ո�^�0�Lv�����f`�V��sBUo+q���u�m� ;F~��.`s�2v(��'p�_K��qE{�7��SIe64�������4t4�X��C4�,1��y1N����<�:���g�1��w�^�Qz���<a�ϙ�a��o+i���rt1oj�������;Bb��A�;�.���U��P��UX0�RvR1�a��(9���F֞�us���V�@/�����7y�v)���`�3��h�phz�W0k�WG���-�o�V����츸�9w�76u
��`�����{;K�s���/��HE<�-u_U�<�r,��� >��Y����r�Q���i�|g�j�G��Z�� ]�ew��%_;e� �]�eR t݌h��(UA�I�s�[�j���FlG�{Vr��,f�T�
���mWL�d�Tk+���B�oT��� �n�t3����
��q�VS��ty���ٷ�:W��澵=�u!�\�=�;����i���Kh���Z�Ji{L|��-�c�|���ǏM-��c|S��a�����!����J���x����#tl��y�����o�虣���r \�����k��m��{ԇc�����l�j@��}�S���#�K��)�� 8����Q�S9im�����L0��6��.i]�NF�3�����%�D������ �T
�c��!i��ZKvٌ�oG�U��wK�Oޞ�p٩>��P*���aBV�׌� V�;�LGʼ.P(uDt��T}��<�Z��anW%��W�7�h�$V����G.Blj���L���$<t95V���A��n�Tr7i�mI.�8�h�Ɠĝ�9������흳��@�ђT���ܬ��]ϸ�F-X����vԻ����d�j	mc�a��H�����Y.�Ie,V�P��F���t.�f�]��̋�����ywFK&Ƴ��᜴M�}��}����'ǥ�nQ#R��6�y�^Q`LBt�Ԧ�ѿ��/����)��80,��軪�ރӘ(l��*4D���C!%WF��W��K�f�\`O:�%@��}x����'�;ox��!�(����Z�ab��gH%V�09���Z��ë�-.^��*y+[c���� ���?u}3U�[�`0~bxm4Q����(�?V�L�^�{p���y�M�+zw(ڳL+>��	�᪨Z�ѫ���VMŝw�����ۺ���ʕܺTVJ�yl�m_���R�w�b�M���U�a	��6gE)`��S#ae<�3׻�dH�7cS��!�4�C��G���� 5<�Y��x/�@s#>7�;����:+s'�9z�5LӾ���CR���� Td	�T��ה�u��h܆��Ʋ�u$�蒑ʮ��]���2�F��_?��F�B�̭�ahr�? ��pً�Ҧ5M�JrLt��-�E�=���*JA'I����qS#�T�9 �;�'oNDs������]p�@�8c�pI�nwy�`�c��yD���@�ub�缸ŕ�>Qb��3z�˼q�P����׬���W�vW'�L���B�v����E�ǋ�d!Vv������kK�^:+[29�
Ž��[ݚL�,�kv4���]�mbc���������|m��D��]Ȃ8�j�_���TiV�����=Ō�=v�̻�ETn(j�^�9K#���ބy��~�N��wn�* �� � L�}5�@(D�c�6W6��F˕}�y���G6-�U��;r��u�M�w��#�'0Y�D�� h��Q���ñ�F�)/.�3���f�� !I5hs��&�u�\KǑ6dHB�� ��4�^�}��t�R��#�*迨�;�~bc�EB�UM&�y�%q�}�I�y'櫍��xZs�J�[��]�����g�Q��o��5�q������b�K�$o)L�7��C5�>�R�R���N��~�⟯~@{#� Ίφ�����Z�;�:������R-���J��б�BW|�R�+���N�0�������X�^��58�^�2�hXB�㳹ݶ�0���n�ԭ��+�ۇ�'@H��N�Cw��^Ef�������ٮϚ�it8X6��B��±B��cOU�D9�q�����t�O���M�7�������:Cf�W!��j��[�����]3v%��\��}!X�6�N_�6��I�.��
s�-�lsxG{N2���5#���FPG~�h��x=z�X[~�i�}����om�����[��5{`�6q��(����.�bp�̕��I�<����vJY������&O�_|>�|��ث7���#�ĝ�}@H�5���`#gl�Ok�s����_��6-������;��a�p��QZ�c�7��ư�PJ N�db���,Sf��]f�b7�z����G�	~�Z:i�N��X:SKڪU>@hZU���ߏ"YTo�岕�=R��S�δ�r�Z:�g��e"�K=]$����B�:��������<�>k|Va3��\Õ�`����ɫ�����1\3��y�X�x"k��KG8u�s�[�·{kV4;�T���	h�㐎��c��Pݻ���(�c��&c`L�q��Hqҧ����Zn츩��TN�q7)\p����N��6�`���4�T�@ ��w�!j:&ksD/�3wP!�⫾�|�����t�؆�/+���ۧV ��\�ڪ���
��[�$���Ol��HBG�T�����h0�u4T1��.m��wl��9�w�Z=��u�d)�H_ڑ�1��*�A��i������\�4k;�A2�3���]����:���WU�8[�R�S�֢��GD�+i��B.5�N�)6u��^o���jY�䕻�X_H��\b�#]6�U��j��Q��.��Ѷѵ�����d��es�v����7�,����8~�興��Z��z�j�'7ƌa��҅7�Y�_gZ�kf~���Pb��.|k����t�G��&�3��������h��Cr��4���-C:������>���vmE�8�E���xk�X���&P��Ub/它5e�
vm���C*DVyu��Z�ܳ�ն�h�yܾ�P��q[KL��3f򶐀��������܏���o�Q#.n���(���b��Y?bN�h�|CB�|un�~������{p�L� !,�7	�}��z���}�7O��>��L�1xc��I×2ű��?�(͈�j�x|�|���4%�=�4��}�S���"�3�����i����+���^(U��8�3A�'�>Πn��ڂ�`�f�� ��e��w)��u��1\ca5�\s�0j���QZ�Ji{IO6��T�]�ׇ<�ꦯ@�k*��[��a��t��U��UN�P�#Ğ��1�vN[���/UE�NE��3���3��S�2ђxs=��7�M��\�cn1�M���^�~�t��
ɜ>[�<��t^p�b�t��v��5�K������K�v��ds	�+�+2�W}�8���a��	��𵏆ǔUd��8k��@b�\�{��|� [���6;3��m��}�]W���H����E���J����B�dV���2)XK%�3���ﾋ�̕�d- 8�# T���|P:{�'vJQ.gx�J�rm<w#�ɽ�`E![�.�OU�gjˆX0^�h�<�ùСZ�߄-3�c�"[��g�ޗ��$ni����2�½׮��}'��\s��Z�T���z�}ۑ�r�F�Y�>δ,�E"���n����wj�����ȶ{.~�����l��;�討�?T&�y�^}DE����W݇}��P`�����ط*���sr�����9r���d��P�n��5%WF�"�	���,�Ϲ�9(�y����nF�5���M�R��!�t{�1�{f�+����ȅ΀tn0�g�����KZ��3�_^k�0$����;�:ⵟ{~�j�ks�;��(�kza��k��n����ڨ�uL�kQ��v�=�s�w*�q�g�&�ѯ_V�g�8Na@n[�#4_@&�xr��j{�����c������b��E��\�+�x:��>|��&�7�*�t"�L�KW��[q�' �Z|j>F��*�X�
��6�����}��⛎dy��{�N�k0SP�Hᩴ�,.�p�1�A(��}���eº�P��XoE*ϐ�4�S/V�X�v���d�J�MՊ��79"�7r�+R��7���
��\�Ź�:�ӯA��z�_ܐ������4u���nR�!���f�wS�>-�k�.����t���@{zi�"�"���yLT>ݖ��������@D�{��c7K�)�m�;��;?�_�j�Y��>A>��0�Kʲ�p4&l�&�G)۠�s[yra��Iu3�L�u28ED�9�bQ�N��!��"4�����@̭㭦Q���x�ZXj����RA h����ZSLs:�W�E"���xB4(V>�]��R�é%4�t�#��~�n��wn�7
�΀�����jt8WP���t��Nכ]�J����w��nxn']���q:n(�?T'0Y��D�H&
T�0osw��H��R�շ�ה������� ���f01�	�mցr��M��!
� .33�Nm8G���uWBT3Eeu��gw���h�Wʡɤ�p/v<�j�^����4�KI��ں�]�mW�Y��_#������a�/y��.���r�ɣm��y��4�����an��`���\��}���>z+߳6�7Yݽ��e��`&ˎ5��$wp�d�Ϗn�!:Q��{���(4hO�Q�3�!�qm�t�3+���G�d��WaO)oNC��Tɤ@�OG&;��}��nSک\��gN�����W�=Vb�O�K���-�p�\�̫����#g2nz�1���[�n�Z+�%�J�;i]�#~�L-���Pa��QJq������4�;f���mtr�V�*}���<�Bv۸�6�m�� ����P9��U�;j	�[̮^�_!�p@S\4?�.����Q�yK�*�:o�{_T'xvҘ�l��A�BZ_A�/}�O���߽�:Gx����o�x]W6��NU��ɱ��+:�E_Z�#%%:+`�+�c]��.�%��%�]��rXr�����*WĢ�:�F}
��5#0��0��973uW/>��/�Mx%�
`p��X:SKکqD&�3l�����L�̠�y��9v��]<0�FΟl<&���K�^��+�_��\%��d�R�Ȏ��d�y֡��N7�Y���1ä00������ˍ6.Ht>�N��=���W�������~�y4y��p��F8[O8�7M�i��ܷ��Qɣ{�k=�kyVe�u)�'5wY�g�R�K/om'�׬�p�Jx�
�,t��t;b�d]jr;˸���.NS�L�.w[s*�q[7�R��������.;c�Q�\�u��5�ED6p��`�wq�8nƩ���:�8�g7�q5� ��F~�����*)���OԸ�g9AK�·ۉ�m<g*%�5	�j1���8���-�؉ؘ�M�����)�a޵��
m��ΑtKȯ2������w=̝ ~�d>�n.��Z��>���4�|��u�w��*i��6� �˵{�,���伝i��U�'K�����sBȷU�;�v%��O3V�r�m0�7��n���v渾��%ne�)�t��n1�/�����R�|�M,p桷��g*5�G:�Vo�-v�y�K�;G����+7F�VM<�u��Ú�t��q�fq��p*��,���+#byCD�a�s��S٫_<�w���^y�ߑ*Ck����i��L���`���ꎅۣ���:Q[[�n��~Οj[�>���3Cc,��&'�Y}{;dM��:R9i�k�qX�+Khqʫ��Ëj���iu���[����)�T8%���kN٤��w �Q�d�F�s�|�������K72����>��&'p����;��J�W����z�O_yKө�b�RK �F��ߘyiت�B�D�{8������\�@�{kk���Yp��ʸ�S���*�����'��ڏw���;���@l��D���:Տ3�Y��1oayt�h�l��� vu6P6��9���l$�f�n�_h��X�ʹ���crVLRr���ϯc[�5��*>/�rnQ�"������8���gT.wJ�}˝�*f�a��e�GYX5̇� J�%�.H�-���*���dD	G!��ע�H�Ӭ�G�fp��I[�5�Z���7i�e��Z�j�x{U���OK�ϓ|N����`ݝ�]��ڼHR�5>��_r�Ir��q��<��mwmL�1��!�v��t�R�&�U������[Pkp��e����s%�t�:��
hJQ��ᦪ��|^e�]���Ω��a���vkwޅ\�r��eY�z�%`���D�'�p+R����
�A��$q	�d���f����vյۇ�Z2,��J�v���68�D�#�H��oػVe������d{u�noQ`��|�#{���'G;*�b;u�d�q�t�]��w5�4�ǻ�6F'g)}[���#��.��G�7�4��{�lt���:�A� �����w#-ŕ�x�btf�[J�y#[��k_m���w�������b;�k��*��̏a)�ơ������3s�tM�̓G\�.�y1P]q	�sn�ԍ�{�����"�0*��]�]y*n�p��{r���e��nX�j�����b2T��t:noKT%���rЇ��]tT;��<�}�[k�����JS-e��p	� CJʝr�vh�	�=/(tm�H�yYR#��,Q�·Ӥ�B� �N�8p���{�쉝��T���g���4<���-��K��_d�@i�@X�>�:1���������jR���``Bz��]5U��//0�-��kX�2%�ͬ�z�*��JWC��{�%���/�������ok�K"�oj�w�Әx�{�Akt��X�
a��歷���,�3�39__��gio��w�x����J63��޾��T�p7|h3�ne����nmpǒ��5�5>�:7�w�q�n�.,�2�欜.�޵N:lh#��v���̼�{vv.�U�X�R����q�\o"{�w��ޗ�g#�E�`\)Pn�C�������,��D)�8��V�Fr�8��X���jQ�Nl��@��O��v_a�XRV����*N�	�gms��f��4ǃ���c1�6��	��us�X�>�8�m��">8V�>�TN�n>9��Jw����0k�+�o�h1�fovӢ�u!��ub���.4@f��!;U�m���ߟ����K�����_���I�b�!�ܴ&��ݮ�ܬb�6wZ6ܤ�ح���t��F���W6أ\�����6'w*��#h�6��sG#h�`��d�wq��b�\�]��n�EE6�5��h��r�э5�b*�j���r����"�P4	��k�{�^ܳ�os�V��֎ʄ�w�%X���M�*�cᰚ������g!'m.�֓�Q	2nq�i����꯾��ts�/G�l'�����}�-�yM��y���M�۝8����ԪɚΛ�U=���a�7{��&���>v�9�_T&�z�+���ZN0m�L����]Uٚr�Gl�z[��7����=
�p�)p�`��BB}ZÆŘ
N�JD>z�M�7�c�i�-�8��
�̦{�hRܑ��'��#�L���Xh��|����h���(��^��k�c�㞮ۈ�a�����?�F�鿾{��t-z)UL!��]��j�T�_��B�oe�5
d��O�4��Q+^B�,M_;9*���*�pc�m�o���
�m�Qv�|�\���ծTk@y���O[J�U��\f���-.r�М@n1�7	�����LҦ)�E�]��F�K����y��J��&&�q�����WBe�Ox��nn�����L	}�8!ũ���X.��Ǳ��=干�/�U�bl�z�+B�}�N֭�[A>8����y�+8!���j̧P�%�ތ�9�/2���Y6pHnϺ=�J���W�v1Xw���iK`-�$#�I�r	�#V��K�2��3]���>����r�9�k��ꈞ�+?�,�=<d��\�^ͣ�h�yj�Eᵩ�t�N��j�\Y����o�1o����V��GOs==��
������wF{�3��]��Ӝ�VK��Ir���g+[K��q`6J�W��T����S�꧙�f�zx�^����m/��+����8�FEN;�����w���.��~��:z�Wg�E]�$�{�K��Z��x�^��9�5�x9�eC�����(�I�P�>��]�mb�kg�'/�>�龔��Tq֐��)��9�_Wң�B�j�K��	4���=���f�Q#����>�W�2��R�:N���Kԡ\����^�k)�eF�K�Wg��q*��i�ڛoE����(4�Os�V�h��&����q��B��o7���ޛM�wl:�_r��`%7�LhZ@TK�+*�Ufn�Tl'C�x�;=,t(�94����U�2�`�z�C�ء��ʻ�QnU�1���Xn��y��u�$<���|�2����-P�G�Oo �z	�g�׿c�����V	�y�C�:'�X�j�ΕѾAݔ�V�c��壔��菣�Yի���֟<��+}���x͗(����|Ԉ�ȝ�sjz3�d�!l��Aن1w_�l�١riC�I�y��y]�P�Jn��٬]��13T�v���XNY�k蕹�9�Ы�9�M�vͰи8��7����T��o3(;�٭!�@ژ/\��9�wXU�76�w�:�$�ϔ�b>Q�绖���4'pP��]8'��=Rܻ�;�(^��mZ����]>��)+헉�M&��G9ʍq�:�t�[�e�TD�z1�m�n�fk�0�	X�('�bqJ��/z�r�T�gW��5�����F�Y}���ݛ{�Fy���r�_�o�;�����c+�mw��b��y�-ݳ1�Z�jm?��W�s�xv����jg�"�jw���o4�Q����ɴ�c9sk��.�Ⱦ9��n�W��V�=K7��~��o�0�%`�ާ[��ő����duLr�����u�ݝ��1Kb���������%�;�[w��Zj�P&��[`�4�!9 �(�]gA�wǣq������Hjk�y��f'����va	.�-�OQ]!�v�eT�^��kh�wʬ�b� >��=��n�Y���|��㒣25`UD��*Ta��@�d�$�۝)�W����<���}n���}_&�]�p �HsT��{4�+D�&A����vwSK�����Ɩ��1Cyx�ki�)�Wl*\��`>G��zXwQ0K�[]:�EcE����&����3��Y\X;	RWl%�&�<<�#	���$OMoCH�����u}'��g~)wB����mC�r�]"وoW!Qіz����q:�������LO��f;q���R�0����e����w~QިD��]a�N����<�����2��nv�ٱ5�u��xk����ħ��HTcv�|�\�����?�j%vM}��.����v�ۮ��]�/'ps��i$ø�;F�S��t��sneTܙ��u��Њ=ײ�rw^+�%R�Þ��k��qo�ԫ>�6%g?.'ٳ�(�������Gg'�S��I!��=Xܷ� ���Z�J��ٻ�bZ--a�ᰑ4o���Da��	}-��O#��w��WZ�Y/�]Fe :[;�Щ�*�q�!��c2�Y��&,� )�>�c:��ۗ$�o{����>x���X���ﾢ�h��~�m��[X�3O��ido:���sV��nv�iB9u+��� �����w���V�Op���Y�b��q.�8��˝���ŧ�۾�;��W�W?mzn���_�"�T���-^�K��2g4�Z���.s��o[�p[=��Qv��V3\�-r�;p�
n(�Q[��F�!��NlkB�!er���c�ݶ��kg��wP5l�㓶U��!"f��V�=�7�evO����Mˤ�:�_Wɭ���ڽ�����^�9��8j�����_-��7]����\:OB�\7
�"�!�OS�e�+�<�����g�픎��>ޝU7����[q��厬g:{������'=�WMU=6G}�lT�0U'�����K����UMf�",����r5��Z�g�T��a�/�ڀ�L��p�=k0M��jo\���3Q}��b����&�:��w�ӕ 7V-�Q�!�����z��y�nmם�D����G����S�)^ݜ�q��
>��M�:�Oq�8���ڑ�'aDv��\�.`św.DOLå��"z��7tk<A�ξ�*ke��~�舅WaB�=�U��܄�E<g*]2�+�[�t{%k�����8�7]�b�*��Pq�^8�c�i �p�_6�*�Q.s�]P#�}Ocm���ԛۗ��qZ�9��|7��N��6�#s�]Fֱۨ:w�KB�QR/.N��œ��_�*�����k�f��Ӧ�����@���}���VW�/d��g�Y��^��r�7�w:ծ��
�C5�=��Ot	�IDb��G���k<��r�����z��T�^��t:K���'��9��w�]�� �h��J{�N�8Wz`<)*�s%ur�m븅2�rz�>�ݑ�r����U��(�L��]:}V��sFu���/��|��{����Tc[=uc�A����@�ա�;Ql�����4�ܨ�:T.��01D����!�}p�o�8���,��}sF ����%]=%�C���˃��P�DW%��h'ʅsa;}�����،�)w�q"�en0!��-�� �7��&QK%Ȏ�|�e¹3��G��\YG'.���V�6[��}]��;K�(i�w��!ƞU�������ޭ�5ں��x�L��������W\LE�I�6�e^ޥYsm־�X�q�k����^e��� ���$� &{6�ڕ5�&�x����[7��s�p��OmM�zl*\;�4�Os�� w_ZQOf�8����-�F����P-��M�P��6(%T��B0�ڮ*w�Q��M�K��b/�����o�!=�OʗH�K��@P�,�93�H�s��a�
&*���j��J94����wa�p˶I��.Vu��9���e�ITFc�5�_J�ˀ��vhU˜��6)y��Zc�Q��G�v�3�r�O���u�>����K욌Y1�¤��n)>xz���T��-[���!.ҍW�LF���v�>��0Wf�v1al���Vk�N%{��Y]|�\,p桷k��F���ֹ�۞I�1a�ўl��ض_�@�X��гi���_g.^<���r���q�^���Gs��:Q���s��� b�/�>�{vv	3�,�۠�C������z�ݩ��\p�Q�n��웧i!���ec�������k[l���c9C�Hr�ka�Y���_T��3����2��/,�t��t5��鯞R��nv��7z�d���"���t�
�8��`ʈ��2�U���|�;}.v��T'y8�Z�3	�5��N:���#�T��lv��_>v�yũo���߅��?Os��1Ҏ���*r���|ԁ؄����}z2�E{;:�:�[��Ѕ0��x���<���zy�֛�j������]7�3��N�V��2a�]a�={-0Զާ\�*��v/G�h��y��p{��#z,��Z7s����1]�w>���޻�p�_��mCi��Wl*\��U[�3bc-=��H66spj�q%";��Y5��_8kq��y�*���6�`�u��B�QMU��8_M	��$w"dN�h��p�܈N3i�9���b������$��O=��龬������r�~	D���ny|G{�ߋ�W���]$����[�.����/�E(��d�O/ri�Y�kw0(1 	��r��S��]�?:L������o�M�����c�У�����8��\�t�gt_s]�ro��g�d:�2jvN��tݙ�#yǎ�F{�ݞo�
od����,�'(NG����,��YhzqʕL��d�!v��#�MD�yq�f�g^�#aOƻ�7Iwnw�]\��L(t���S.k�!tl�Z�vO"%dl�F��ˍ�m����ƛK�R����a���q0�\O;sQ���{�1�gZ�`[V'�C��\�8��q�v�w	*��X��6�]��游�vp����aiU�'Kd�s�_i����Ks����)do:�Z�͹G5��:)��K�OQ��o�V�EV�̛V���_g+Z�O�׷	���ᜎhY��,�Gl����W������b*�ɋ�SSjq�ڊ��4Pt"��D��9j�C;���p���ر�c����2�
�|�&�*T>3��Jfcs����t�گ|{���z8�R��������W���\EXA�Z��733�
n[�[�q�����Q\��n��u�l���5��\h�|�w6o�Q�z�@�mkg�]���D��R+��Iuc�R����:�k��"�<7N���Tﶃ�\`�#��Z����Ԏ�L�u9�VL�K�� �,�U<z4�-7Ws���b���c��w6�H̭5���{{:��w+��-�ޮ̅�3����]�F/�����Bo���0��wk�q�iK�KwxἿ�}n�ۈ*�+9����b^em��Vt�q����ʤ�Q%�rg��n��[x�m�/cg9��Qgr�]�'�1�݆�^�
�ܧ�w
��#��KAK��h�73�-�LW4�������t������/��N�Z�(x�X[�u�Z��s{X��nkΏ����t�|�J������9��3�z�XE���]j�n�����M(o�Q�6�o#K�j˚�h�У{M�P�j����j�ÊW�R�MF79�U|�9��|�n1�#q0����Eލ�=�]��7<��7/�!�l���MKy5�cu⸄�M|�15�n5�-쉝Q�7��(�QҤx<!^�*U�gVz:�}�ڬ���\�=<jOk[�:+$��/��oy0��R�@ڄ�+�q��\����ű/�eR��}K%���Ґ�;���	��gt� �Y��tnUu ���wQ��Y�ќ��$&S�t�ڐW���|�ZPU�}�b$�^7wa��r����7�!��_[�͔rc�psr�F(_f�,�+��%��#���v�
�t�f�Z�g3�(�k���1wV��i��F��L�ŝ K	a�ᆛ�J|��
�Xdn]\��u�%�}�V����cDZ2��CW���[�X�]x��N@3&`��}������h��ǋ;����j%*�؆f����ĩ�Rr�ݾ�࿞��׭6��β��L��N�e������eQd��9vP�Ֆ\��HQ����.�H^v-��X�n�B�U�q��L�9�[��@��CD,������OK��g�/���8�*�=��/lu�)+]e`�c&��7)ә�I;r�ĕ�GZ�5	�����ԮM�T�)��X�:�h��A84b|7l��ۅ;o�-8����hrdn�y�4r��ܯ/�8mi�*Ɖіn&�
C{�o����kX�z��	�sMu()=��e	JrUՑ�̹S����'G����z�R�='5�e5�n>�ݙb�Cfb�G�UY'��W=���vh(t�|�)��6ѭLհ��U����#ԶZ�:n������r�v��ꂔ�&W-J�>П�/�Zѥ����n<jh�8+�_F�\�]5]���C{�`�ѕ�f�io@�����U��3 AS#��f�Ltw�"�xsz�P9P�w��:�f�Ջ)�i[Z9`,���<q�U�aX�-��7N�,y}�AcJP΍R�/n�-{W�)�ڥOqֱSL��ܦd��u��3�..�O�z�����o$�O_a�N�[���_��Aۮ���=C(ܦ�\h�k���5�֋�V����`�bY畝Z�:u�Q�.:��d�����!�tu���>�0��9��E���w��؍��c���
��2��+vp�5;.����0�i����@`]��굘�����B1�+����g�[ Wi��@�)1��`˘{/"+G
t/�b���^P�قcf��P��X�I�,�,�S5�qF��dx��yq����c��ϵ��ݽ%7���X���b���p�m���&V�ڇ���Z�I���K�w�����f'Vr�Ӊ���]Y��QV2��覯y=�=Өd6�8���Y�V��o4��Y���7��%I�L�E����V������oMZ��rʺ}]�Nw�d�S{8'�;�j���A�J������x�����'�6��q�\�R]�ސ�Pu)���>G���k��Ȏg��Z`�"2�8���b��OS��I�=�	ɵ����y8��� m��"��=� 'U�����`� �Y#n�7�6�H��ov�V�*��>ú���;�Z�]Ο��=�������?������f9rܮt�5�*�b�X*6��5s\��˕͋n���t�5�S�nTh�͝���C���v�]�܍���l�F�r����,h��r�\�h��gw6���.a�(�ݵ�*��-E4�;���h��p�0[�:��b���r�JH�&���Fb��;���(�]�L�']���,E�ԑn���c���9`�R4E]6����ҀuWwU�b`�&���"�#]��LR�h!/wi�A穵�p^w=69��o^݄mK0^�qoQM���dKw�{xog��ꪥ57[+ހy^^�����9�.s���'W*�\ʂ�Fb��{�q�5U͵V�n�vZ�w�BY�>;�L�w;��c��S�[K�b<�-�ǁ��Z���wo���~w��Ë~�z.�r���_l��/z�3�0_o�- �:�����;���/X1���kg���`����[�@r�x��a`0�1����Җ?V˹�C�U�ۅ�J�Ue��.&�$�U��	�[I��ޝ��Mu�W��J��:N��I�%���r��f���׬-�hU:S͍�j�ᬼp��OmM�ql*�Z�7B�EBW��S�%7ɽ�l�z�[ɨ����ƻ\^tC�9P�7����)��]��Z���Ӓ�e�6��p-�6���MAK��
�n}	�ˤi9-��@�l>�/�����)p"�ߞ';�B��Ұ�[��D6�4�xgJ��o�h���u�ٙ�!M2m�:ֻ2e���-g��X|t`~��1eIB��Ջ���W##�����ŵۼ���x\�4��j��g�!˹�&�Sհ��8]wer���AR�'�n�yk�KR��Jň�W՗=˹�&���������ܭ̄��B�\�7�Ȫ&dh�Ϭ�ꏵ{�>�Z���l�j��P���.M��־�[0@�T�wa)W)[LKn1���Lk���ml��EG������/<�h�w�י�'%vk�uj�y���jp7��qq�k����jS�����d9�N�wp̸���׿F]Z��}k\9����[9����'�SV�]�|'��]nb��]Q�f'u8�:eh�������yfd��t����fs3s'�+J暸�ѻ���"�����6{۔Q�7��z߸L��}Q�ߗ����*�9�g�nuzo˪e!�(�2Z���w�G�;#	� ��ݾl׼�~��!�78*�UD����\�ͣ´gdq[m;W֕s��9������m��uϯ⯩>��O@���Pΐj�G��iv�xa��xRz#kF�ك)s������=bpT}�Q�U(r���a�랂{sS��v�kn�-��z��p�T�Y�I���|����8oTԮ���m�&s�vr�uw5��KE�(���y�$�e��Rc��ޕ��c��2m�N��Q�e��V���������1�چ�Я�F�
� �3����Yun�6~�O�)TD���Zɢ�ˎp��8[O8�7M�� [ڎ���q����#s�N�D�D,ϧ[5�K�>�N3y�$l�3եbɾO&:M���;Ľ�_r�bQ?O��-����H�n�'��^��s��֍j�T���L�ĺf�L�Q�P�#�M}+^C��w��� 9��gpW{�/RP�����7�4�\�}�.�Sk�;;g9�z�Uپ��N�.
�W��T��T�T�L5��h�O����;s��^�{r�ƽ	����5K={�;�8���I*���6������=�躹�+dL��u�(��ȽhͪȖ�/2�f�<\���?W�O���Xt��
��\3'���\^>�5�\ug�%���r����|jfy^K�)R�]��|����]��*�))�mz.Y���ms̒]'P�H�2�s��{�9�A�8�����D���p�!ٯdw�t"P�%f���;;�{yp��<W��,ZUЭkmv�iP�g����U����f'՘�6�{�N���ޮ8��]�SS��r�)��K��V�K6R7�:T���O���]�t��_M�T��b��s��[��jr#��ok7����3�j�����z!��J+�����t���Ľ5��UZ���:W8�R������7��d���
�+f�&OH�wU3��\�s��u��a�����79��u�n
����w,0gsi�03���v#] c+&]Q%�K�KJX�����\KOaJ���s4�gDꞾ��+��RR���ݠ#'�_���r]��SYv5)}�*��mn��T��0w��-����RXvt	]j����.�Wj�׮3^3{.�b�_j_�����w8"���0����{���~�S<�Γ�U��<��EC�r�]3Jd��w��8�r�̺�-a�]	�o������x�$+����P]�P�\��l�*˘2�h�۹�"79ݚ�Y����J6��6P�����*�Pw�d{<�3;���̽�ߡ��(ot��œ��J����^�����>�����laj���ۮ��_c��M��D� �yfp� �s�,�ۍ���C�X9�a��b�W<{bx
�v����o�*fyE�i����_%�j|�n1�#qS�}zv+p%�~ƞl�e��`fU��Mw�;��v��J�č���]�*�)�imtm���]�W�P�u��eJ�'Wַ�dm��'�Դ�Vܿ?W.����)�j�o\Y�p5D]P3D�-�V������٫��Ϫ�f{f�=1�T]O���ٟvh���-��"�!빌}�湾�
�3�W�^����g;3�<j�3�*~kW��yZ^կɖ��\�97w����(�����/r0�p϶{ݖ7�2�ח'�y2`G=�G�X�+*S���6��R����d�蟽���c�{��R���(F���-��{iw<�.��tʰ�jK��Tr�Z��)�[׸l��)v�]��=�;9��}n�૶1v�W�b�>[�M�3Ӝ[���&K��c��Ì�M@래*T��1���9�9J�hć�OS)CO'K�Iڬ��j�w.�U���ɗ'��l}�x%O��v�P�������̓n��q$���x�5]��;\��u�]+{$u�Ir��Է34#Sj�m�m���ˈ�SO9M�i��.����y)\g����~�D��LӒҸ�y!'{�<k�\f��9P�7q�è_r����m���rdl���H{�l-��%�
���=��s*aD���3ڷYG;�w�N�ۏ�B_,k~g�B��ҿ��o <���"zl<ɔ��_��-�;U��'��v���j%ne��4.Z�1œ�x��U�םx�q
#|��4清ѳpV�/�s��E�� �Q\e�i.�*�ps�N��I15��q�k��t�xS�ڲ�2y����X��!�B�9�s[Wr��5N�=�Q�r����01h�c��yj%�ܯm��E����g���T��P�8�������VhR��� V!��u�F�z�[V����k<�j�g���v	������,!��T@n;����)Z�g/��V��P��:�aHm�(㳂Ү�@�/��]vm�����:��S�unȽ͘-�<��r��2V��j�ۉ�̥H���	��K�I����!]�1�ӷr��k��|�"7���|CS(=�b�����.��Y�ݎ�w�+��-r���O\]J��v�y���Ԏ�ˇ�LШM�;݃Z���|�3�ڥⱚ�V��C�U�6�؇S���)�V��ClY��*+i�ևb��qjR�T�[���i�ݿp5\��������뎕J���{q����M�m�{�_Rke���t�_v�8G��?+����n�6[�;��Kw�t]��-�����������W�N�3�>��ӷ�Z�R?���ψ�{��s��_8kq��zmR���+!ԩ�|;����Ao����E@iTIY_N�h�!���8Ձn�����S��v��Y�*%R)��ڗ�6���M�l�n�d��y(5
/4c���8�P�ƶ�,��d���ہϤ�v�`Y�>�AH�8�8�w5�ur���q�
ٸ��횅2�]�6��wצ�-*E�W�:��'�q�u��)՜`@.sk/7d��v��/-��ۦ$��a�9��g^փSѸ"�p�{ 5�+�|�	%:�|�Յ\�x��������C;�8Њ�Ax��TQ7�g\�WƖr�Lw`7p*�}N��ugwK���K�a�ʬqAÂ9��Qf���;x:�.��h7���N.&9ۚ����ו�R]��ε��'i�r�]�����X��j1p72�Q��#�+gVG�$ �J��Bl*��֏�"����74�y���Z�Kv&�S�M�c��BYX�q�8��0�}�H��3D�ʕ�o�{)}p���yz��5���]�q��+{.w���~�8��`������*'�2����B�ڋ�����+�?�=v�yũz���V�1�N�,�U�|���[\ǉKK�f�~�\���t��|�ޯ�^�X��_�c�s����E�uL
�1�`�TD�ҡv�}p1D�|�s�;O��\�ʾ�����!+8#O�U���Z�=�*�K��l�z[��p�\co���0�Z�q�y�k8��q���.�p6(>UR�/���L�sh'8�@�Н���6j-����u�i�a��Oh�f�N�W.��^g��^�џ4Ւ+1�:L��ʘM�lZ��d#p"���\h��\�Gۆk7|����X1��;\Υ��HtJɇÕg2�{�$�p�f%�fd�7s�t�o%=r�(����q���q���L�;�4�O'��5��;M���礫��.7��X�dk��x�W�.���l5�-1�P>���\���;�"v�K5k�au�륍]�Xo�b��{���ڞ\Pٓ�>�^�"+,�͡F���dK�w�S������I�;f�m�iv�-�����sӝ'n�u2�'&�����\��9��gqU	s��M�w�s�D�a�p���]u*waU`z���#��1��i��֝��zvWw4e�����Eyr�]#|��'^xΧ�cU?VG:r�>���=��+⴫��!�^��Xp��:It����V�r�ځ����
)p��`Eޡ=v�o�O�D�R�I�=��LGL4�z~����j�̧W*�5�̢��h�#GK�7/V��`�q8����+���eh�O���_vU?5��b{�7��Y�*���
��i�^�=SΝ��ȩS��2kv�Y�I��j�R��)����ܐΦ����:^��^�ɹw8���1�:޺p�1_�0����LY�c���˺n�E:�J�_-�b;R@��»�A{u��(�d���9vCr1������b��;UM�T�;dv._8�R��|�t��tS���=lW�13_s�o{��*2��0}�ON)��|0V����I^�tp+�y({���Y�T����<��Y�w$>�'����=���£�`]��c�ƴ:��\���{�_WػJ��8lP|�$�Jj��J�Lt����)![�\���o.#\5��8[P�{jm����v"z����EΣצ]�$�A�-*����>V�k��v֭q�O8�D7M��l=4mI��&�A�v���|7�6�\u�'L�o�<����F���<g%A�
[�S�˫�su-V�K��=Q�5?�(���َ��I@w���M�6����-�ZvEAV�|�<��;]
�C���It;�o��Bw�^[�@.�R��0�!�a�q������6l�sR�%��3�v�YV������u�h�wFsκ鲞�9B�u�i�t3��1Jɝ'R���*m!wk���1�WHU,O6�oT 4t+��+�fg7��mr����C(��sV;ĝ%zv;�V�z58�ٜ@�
7;��T�dn��e�|9�cln��jz&aF���eր�Э��Rj��;9�	�ۡV��5�=���LT���b�ajt	�Qd�.^���٪�k�̺��xPtU`X�x�Yﱇ��u-mX��7���x�-�0���ځ�o2\�ۭ0�]�R-����a��Oq�.�%���*��}#��qh���ܟ>|�ӹdwe�ar���[����ܦTX�tv]`;:�Y��v��ace*јv1l��n�<*�ws��w}Hn�jJ�:fv ��j��������Qۢ)L�vݮ��
[��z��3V�\�t4H*�)-
���ԗU�i�+x�k4�J���rjԓ.�.ʋT�y�,�Ub��T7٤p�OnP����&�����J̠� !��q�&��;��S��#��7q��۱d����,���t�%rۈ^dw�NУ'`ۢLqXƓm���˻U�R��Si�ხ�r���M^ؾC����}t�<no���7�o�2F̮����8����-T�S��Ů�LM�����@�w4(�in�C s��C��k'4�vX��c�F�U3���Z�����Ϸ���d��aWx����q�w-�����u�hm]�!�k&�^n��t��7��iA�&!V���
���>��e���Q�ݟZ���Y��5e�wX
���xX8�E�:od������u��ܠ�mD��F�����:Sy�}:�r���V-�¹i�Q[�]�]M;&,���P�|���F��|�V�ѱ�m9��u}��x���mk�"�C],4�&�P	���� �/i0t=5��HH��s�O�u�{3����V"��e�)�3�fl��ə#VV\�^�H$�����[�Y���coP��z��$p��oi� ͞�f��u�����0��XƦ��9j�O���j�<���[�.w��wC9�סu�~is�f�p�k�]'�3���^^B�n�w}�9���X8�����)�ռ�2�Xb�a�3��ou�U�#v܉��H����4�I�[�|�g�<�n�u,�}���|u����Um�̽�QR|9�;�.V�R���bL޽�yڣw%�l �0r|��7G��G����t���o)mځ���m>Yv�믌�o8�ʹ*�:f�inh}�[�R=��=*�,#�Ë_ɗmWs�s�8Z̳���bm������Ԭy��|3+����f�V
����27A�kZu��	�5���ŋ��������u�v���m�v����F�i���wW���9:�����+�� WL^����6�ƻ�~y�������������e뢸BS776.��ݹ�Ld�n��&��*1�.c�+�K��r�$d����7.DX���\�X�B��ndԆӻn\�E��Q�,lX*I;�f��a(�r�(�Bwv*���s�FK��lb)0I$+����d�8.r�\��M&)��PRG7dmnu")�'5�d�r�4���ݘ�:D���&.�w.�����\�Q4��	ݺ(��鈜�fa������2��R!%�4L`�l&�LRH����q��I%�Ƒ��!]��X���jw]DS�*Ul,d)}IoR�
�l�.�	r�A�tz]�m�1f4B5��+6so���n.�n)Źrl�L�J�,'w?����I���k�n5�G:s�)�@����sٌsr�l46�ľɯ���igs��X��ns6��F�EMըCO;�r�h��-�.{�gi�g����/2�e#������ᚈyJu����ˬ�\=�gvL��n�Y�o�Z^��鵜�.�G_\GL���R[܉�o�O(�O%92{�mwi¢����y�����u
3�»��bU�q��4���V-J�_<�~��������)y[�]^߆�n��Q,�;݅V�G<.%k���^c��T�a���tz*;5����y�]�ms�6��a�ׅD�_ ��6�9�U�&�]�puu[j�iR'w>di� �_Iݨ�|�\����p�\c���z�ꆙ��:�*�q�Z�)y<�7w���*���U������9�[���e;�7��"5��e�u��"�oe5w~�#ݞη�sW���:�D�Լ��We���78෦։��	�%�����0�i��kzA����Jћ����kHte��1o��B��b@�)����/�q��,���#9)Z�]��7,݉[z�)'����2���!�M�_/�Iߒ�*���[4R�{��[������+�*����m,g�q��}�~1�Q#S�^�6��N�������SyX5$�;֡ݍ��ʗL�B�*��.�ls�z�V����ss�;�D�V�n7�vht�5a�0��_7lҙsQB��1mᅛ3DKy�'�"��={%���nc�������a����q�Jqq6̤�3��i�ۚ�s�Ay�r��ځ�%�e�-��b��x�S=��i7���g����6����Y̷R�p؛��գ�Y����_,է���w��`�q���;٥����e#��S���U�E�φb���TD�Q���4-�#Z�����Yx���{�Ƶ��s��[�9��0{�f*���{+a�Oqq̊Z�ﲄ���{�N�_)z������^+%)xo.�P4ZV%��0j4�$NN������|EkY.t%�fujq�@����<�+��<q`�2�r�ÃĶ�C^^ \�T8����+��pQ�AӖ����3rm#�Բ�9�\���eW_=�p�S)bc�G/$�N�����N��Y��Г��ʕ��\8�c�we�z�u���}82�F]R�Д3Rk23��1;����98�F����ъ'�䛜��}n��� _Wأv��͋��6���l���:J��}�J�Ue-�>��vW�یY�՚��yý��3��kn
�Q�R�4dp|�$�Q%����RF��.+gcqCan�x���c6��6/�L�;��i5���تt��#ez$3��}��7�����F��x��K����}�bi��6v&��ju� ��Ám���{�-�p��Ot<f�%�5
d�j�b�SyܨnL��ѪY����Q\ԽypLvh\�J|�6�|��V��l��U%=̢�gf�H}�F�sR�&�����)����^��9�Bנ������i���[�)�5��6l��)��bɍ׊lց)wx�t����ܹ��������sM��n���C��O��@V#}��;�r)=U�"����՘%:UP� �a(񡠮�읾�Sbt+�#+gɪ�JY���YY�T}4���z��e��[Yv�E�8ż���F�.L��KѨ���ǹr��j\[|�wl��I��mƻ�f���s�*%���Q=�_J�$�s�n�l�Н$���n�������jځ��ϵŚ�����3�)�r���ލ>0�n���\s�j���V�}�^Y/�w�]+=B�M9��`3�� k���﬙�c܊֮�wϠ���O�3�*~k.$`6|�.ȟ�=����V��jNU��\k�T]/~���Խ|.MM=���[��z��^��T��CZn-��,8?�ίM^��Uk��2�R��~�$ᝑ�����k������w2�J�ưzo��:S[���1���{�V���q�D�}	;���)�|U�F.Ү���`>Y��î�j���:�3�iYfi�/��\����\k�����M=F���K�]%k�t��'@����ra��D>z�d���<k��p�!׆�˻;,�^����eX�I\ގxW�{�-�O�M�L��m��
�a�+��of�6�Mrt��a�"jU���ɥ`��ɼ��mn���kSVvay�|�9k쨥���]����㔨˿�9��H���L�[�X$i^+���޼tĘ�l��f����#}�1�P�y����M|R�
�n'�!'O�ޞ6ɼ�ܫ+��8�q�]5�%����%cW�[1١W&����#���W���SKq��+����S%WH]P#L�jV�_��x%uEfvlb�;�e�q���o�b�|�D�lR�s\Bꁵ?�M��#�]�`��)D���;�$�gy&&��Шϵ��:s�)�
��jD�!2z���{��}��<!h�5yeG���d��sQ�\�+\dpk0=�h�V�S�L˕<�X�Z�U�7"[���唎�p����yJv�.�vrB���˛���uT'k�w��=���-�y\yҵ.w���Hk������ry��)���k{�b5���U�p!	�quK��N�n�̧#6[x�X��uC��]��u��V>6J��,9��B�U�.��A��@�ݞm���L��f��c�+� �j�h&7n�_��=��u�(a�ԫ�a7op,�|��5�\.��<S ���Wbk%�]��;3��I�[�PYW������gU�����XO,��^f�:�bS.�+pC�%ED�P�J���x�f0��\�J[j��kϘ�Mɴ8œ����P>�:����N$�Q��a�ׅD�|�Sp�|瞅Z�5��j__` ���
����+ .!����j�-�c��������n�7��)�{�fu��_S�,.�pb��	��+Y!'{���w]LƂ\�ѱ��n;_��R�F�
�ܧ�%=���,�������h*���7)Jډ�iM����������;*|�U
U'�t�i͟:N�0|�w;a^��8�SJ��k��{.����U�W�7.#[x�;��A�r�o���.ˀ�{4*�.j��l&*2!�f�˚������!��]nz�]���Poٵ�TF'?gqIt��L;�;F�gM޳ی��Y��-���y:��%��1%=49�S��{��wL�X��	2U��CIҼ@J7}Ż��F�m�F�����yVf��j%��gV��L=�7�p�y��vsO[��y{p�v�CI�^��}FgCarf2��ܳ.����Rb-��{y�ݾ[:�m뀮����BQ=��*$-J�\�`�M�z���ܝ�F�kF%��X11�i}�,HΨ8�s�G��Y���z���u3o���[�Ws��Э+����H�;M5_k��o�ᘪm�X-�͌5+��$���B��N#c�S/o��we�߽�P�nr��o��U��ĭ��+���(<!<�7X*hΞ�n#�����yE�z���t�^^Ӎ�r��h�=F�zQ�g�2N��]����S�q�Ef�/�{8i��l:��o;N����[���*5Jʔ�k�=r��s�B�2��(��䛜v�eg��Xހ�k�Or��S�}��$�I]�ė���җ}��sm��/�^ס�廮'���+�.|�NW��������T��K�M�VK�}���z�{�����M��T5��-�����z(%��v@�*Mc	�{>�Ž���T��xj
]�����񜨗I\3a�/�@�AS�:���Uޞ�_�qZv��e֋��!��W��l��s�2��Y �1�-ʹ˟r�:��흝��Y��v̇z�!��^���"�U/7�)*^h�uhd޺�*3x��-I*/i�ל�\������W���?=~�����t��+;]��q�M��Ύ�GD��w��s�l���e�� ;չ�{��3�.�!R��u���%�]��i6����Di	l������I|���z���Oj�N�H��^�i��Ue�˞�ر��V��؜�w_%�r�ͷ/T���Kg^>�B�B=���N�F����m�9)�⸽똫�3�7Q�uK%8��ibbi7��qc9t���G���v+�X0P���MC��`69�O��;�k�Nt-p歨���~�7~~��zM�����!T�g���w)оq9�^���.�^���Z���s���ٕ�ӝE���y=EIGք��j��K*қXy�+'����+N����\=��j������jk����O��}담P��Sk�ތ_^���{8$,^���VǼ;����([��6���6Y��K�Z����V�x1��uJŉ��AV]�%��x��O4�r�fr�Ю���c:�P#����vT}'���=�:mM�ɫ@����0=�����*��
��w.��7Ml*�R�MNb�z�Ӿ�~��A����7�h�%a+x2����q�Z�r7�֚nr���n�X��]p0WL@:�K�"�vn���7�}�:�+�Ʋ_\iq?Z����\:O���m|�1�e���R�þ��H��Hd^��Κ�7\�r�r��yk����i4�o��ah��{]�Χ�}�S��
��L�Gs�k&�O/�5ٮ3k�-���?z�%��R���7w�H���?��j������<����F�p8c&������J���n!U)�NK��R#O�(��\�[1��p�U�dk����P�ur���<�M��}<]rG�j��V���v]߳jD}�v8w7{��KZ�:�K��o�b�|�D�v�|���G�6v�Ca�(��n	�Z8��5.%��Ǔ�������by����qq<��d�1�"t����	޽|M�q#Y�Y��eG���gWg��{�og�pz�'+,FID�!jJRЩ*�ׄ���&�����y
�dW�Ty�s��Sˤe� �E�,f+�9���'u�hDxv6Ub@����Ȗ�|��U����Mn���z3��.;C��Ƃs�`���w!̤����� m�ͱ�A"�����res,A���,3�P����.�z�6��{���䶳������9T���G$�eI�����4��1s��"	�#|�V���R\7�Vr���}V<,�S&*u�1O>`,J�t8��>.s��W��NlY臯�7t��XC���5��-��+k8����g�Z���<�y��'n�*� �w���[�μ�m����{Q��
��|��Ko��f�x��� �$� �ո�Ox\V����DJ���}�F� Զ޹�����#_��t�X�Ȇ����֗�$�#tٝ]�S;����:�GGX[��b_����~�N�ޕ�{P��i=+�9����.s���g��C��z�^�Ԍ�%���U�w�7��+w�9��O��Ӿ�P��U#o޻��G�]� '5x	���l�Q�_u����f0}eR��夻���O����9\���4�Ƿ�#n�V�߽T��d���7������}c�}�wU����"�<�\�Z&4�!6^ʅӱ��Y/-pԪS����,��pޚw�X5�Z�k&:��W[��5)��%�ج`yP��{�z��?Xl��a����.���\��,|�Y՝����V�m�X`���DF;7�`s���!��)�+�ڜWʠ��g�՗���n��i�
��=��4I[��Tg$�.�G*s���[*�5:��R�dӹ)m����p��b�}�u (Ѩ9�-Z"�{�+�U��3���8���"�e!�x�X����Q�y�|�U�L��@��E�c�ݭ�.��F�Z)�:L_f7��*\�=����m��U���Ve4'/`�4L�̢%�{��G��3rڈ��]��`��b�v,p�vk&W��
�e�{��+�"�:�(;��0�#�j5�>�9\5pɖi2ٻ�wHv�/�iP ��$L�8�b⧧N�	M;Z�����M�;͔��})�FX�e��^�93�6�/2<��6�Y׉Ձʔ���]��7�5���=wa�����Ч)���oF����2ʺ�$�oa9�(^�[��@�.�HV�i��Ks>{5o=6{�Z�EoS���nr2�s(P�r�o�b}y�L�"�M^�ЩSF�GS�z�f\Ӳi�`�� l�A��ΩY�m����	�$6̺���)�q�=z��L1�����ᴬwfwR����x+AKw�K��jy������Q�c��y��:�"]�l���"��ҷ���P���|���a|��F��8%j��ՙ����]{��vY��m��e5���:����_�bK��m	R�@���Vl��۽\l^eJ��k�[�{T�8ϝ�Q��ײ���:�_,��5b���.�}O!�z�m2��o#�B�}0�;�ϻok
}�+�;6�af[�8�{]X+��ݙ���㰍��:} 9�� ����iC$wu��y� YI�X��]Ef>�/�K��N���T�$<�j�ʼ�yНS�Kٙ��>�si����-�S7-��ˮorA:Qv���Q�iL���v�]�KJ��R�V��#[�YR��r�0s�C&���N�ޕ$��ฤ��ĵ�=a�ge�,fWBo>�5���r�GM]&����!1\�x�"�,�Lɂ�'M]>�ۣ��C@�|'kk7��ŭ��^���x�Q��'V�5�]l��(Pe�>�mm�e�}h�Jj�w�G�9TG�� �g2W;��t4�/��mBQa<�qnɽ(o*滯n���B�T���7�<0�� ��\��w$���:]��
p�9�00���]n*Dj��D 5I|w�ȇ`8�$��w]�b/�pо����S�w�FN�x�U,&;)l:b雔��F�ϺGD�������ٷDl�y���%ǫg�wF�����=փsA_e����+׋�Xc]-��Mq'c�*����ć;�N�^�5O����PX�_��x��U��z
�n��_P P�BR%����%�iIN�ds�h\�ƙ$@rw&�$�Fɴ�D�1H"PX"�M�0����j�$4�2!$��Ɂ��4�A��ˎ�	(TEwt(�JE�1���1b7wh����);�¤���"!�����n4(��S�4"f"!)���K#��	�M�fPPlٛ"Pa	�JS&��)s�QCD�E)���	d�Q9�\�e4�Ƅŀ�SDj]ۑ&�	�.���ut���@|��{Z�z��������eޜ^��@�a�ou l�����;#�l��cޜA�RjN��(����q5h��Γz�@�[�^K���b�g��"yv��vK�B}I�31N���$��83ums'0vU�p����s6h]9^;� �*[�C���1�}�͂����P��BU��~�s����ś��缋2c2�NQ�Z>G��W�Ǫ5+��j��&���>��=��?P�m%�bf����;��=쌸�Md���\�/x�s6�y�Cq��m�Q[w�o�Ƽ�O���̵�x^�V����f�w�*�V�`�|n�p����x���&�=}x�%�Z���-���c��/�LG"��蜶�FP|����ޠ
4r|��������bU:^�s`�oo&ǶJ/�/���YCoT��7��g���N_�՞/�U��`��L��g���z�x��W�j��
M��<Q9�X~�2!U'�����,�k������dn^G��|ɱ/�尽/t�rMw���|%qb�&��S�<�i���{S�b,rM�֦��-*8,�����מ�ص����Zn���uq��ii���^�����1:~��0-oc���V^�j�Nm{��4
�P�갓����[u��$���n��A��}ShvP�`��|s��[��%1�U����r�u��R��$��T�^�A��*Ҹ鴠#눾��'d�O�#ۇ1]bM�V�M�G[�!�Dy��`�mc��3V�do{�Y�{�^��a�yh[�렲�Q���j��E�2�k�a�>NDϋ�B�����!׾v}��G���\{�g�|4��	�:vK���IU�L�ʡ�EL�1�6���7Q.��n���]�_\�U{]?�H�|s�%��j�}���p6. ٞ�\�����.n�cXfϬ@9�1qS)�rۭ[�0r{�h�zF���o�'o���0�<r��������3V�htx	�|d�W(�MM@c�z�x�!�����&���ӹ��}�/X��L{���c���ﭦ��?v�������r�T�����ޤO�X�&siwşXә��m���:��MI544�=���2{F�=�ʼ�2��J�Ց�/��5^��mVα��i��Ƽ �d3Z?e��U���I��~:�k��9�^�q�:�'�x�;�u���H���i��)�E���3T2�CH^��"��/�NJ�\6���\�=-`ѝ�'�ax�nU���uXE�0�4-�9C�(�}�E��X�	�N\����՗3�@q��^�VfLcx�[��g�~���r�C-\i{5+���mbA�<��{>��\H�S�^˔o4o�:��TA�8��Q�"��t��}���vS���}���f�`F�bK7(]MN�;C��ڷ֩��t��%�Q<����;�K7]LO��^��f{ᵡIzplS�'oenUXcyW������6Jee��Xa��G�����#��������X��Wv�6+�տ���:������T�N}ޟh��+�^���v1!�#�T����כt5�'3~3||��Ν�/ī�i��D_p6�j��:�����پ�0�$�σ~[��Ə>X�������=F�3�m|�H���Pm���BQ����_W�"9ǚ��s������̿�z�+ϖ"�}jI*�e��p�����%ϕM�o��r�Cl���ے��Z|�e���O�VG��yg��#��2��ԐW���\^2}�P�� x����j���D<��{���^0�G��G�Ϩ<��l�>0E�Y�tMNG;��������K@�?� 2�ڙA{!��.[����q�s|6T�J�T���Ƣ|X���,�9G��0c�_ź q^*��0��z�О�����'h_�)�,�jO��ֲ0����ǩ�WB�iK�b!��cwH�����4sDI��P��Y�����Ȕ}���C���;��5��`��lwe�Yc9�A�ܧI+bb�T��e�����ǼWc%��}�T�')���/�}����
P蠋ٝ_S��vd���Y\�����z�b�Q�,GǌIb��M�ʪ�;y�N���c������-���}Y�6�K�KR ҅`�|b�"�b���IU���5|��G���F���Yd�%��W�j�1\�4n!L�֑����ӗ�%zQg�=���*(,��U���cF;�RDokEܰ;�L\w�YG�V�[^�k�s;�U˴i���"��������z�]�c����z������&�M�rl�4���Z�ޜ�m�{cjr�2U�����x�����c�_M��ߚ(��EU�u���p�f&K�f��3>�mXs�c�Te|��sc�|��=1�H��Zh�����g�<����7If������w��6f^����x�L�V��f�뜣��8p�eA��s�:mCM��s�7��x����;�p�"����V����s����^,�~S��M�'����F�y1\�Q����T��57����P���Yrt��WC2�u�#ϼ���h�}
��q7ux5#I�4�e�gO��#,�V#ܣK��1�b�ަ��t��9��.��U�Q�9[HF���T�	Fӭxv�q#z�`E�Mfoe
�Chmi�.�htb�s-�/�N� łVf��[�f
�����x��nY��3J�4��J���n4��F���+�P��U��)�t:���,s7��p�5��&9�ƹ��uz�{9u׎}eUD��*Xȩ�������Q�ׅ����g2{��gx��ý�W�]�����D��@�e�I|f:�*�te�u2��Ǐn+��	3>��;O�����s=�e�9��<���鑎=�g��p�n@	�704z[>�diWbي���[w�م�9��V��.u��4���9�~jb�&���m(,�y}3��3Nv�.ıv	7r=�j5�og�= �B�ơoW�D��,��||\�ĶЛ��fb�$��
�=���[}�yQ��W�H>�*)9�|!�����N6Ž���\���#M�H<�y	���;N����17&v��C�;F�t}��j�e�TjW!��UM׉�]FLф:*XK$��>���_��TX��ˁ_/e������h��/x�s6�y�_��q�UoD?Y�w���q���U�Y�;��Qw�D5\��avQxš֬��}���>���>�����6����SW�o�z�Ŏ������Ƣ6��O�7J2�y�ٛ�� Q���N�6��ߟ���2�/To�+��%�Ơ��ZNf^��>��%[۵�{�
�aJH^V�߭P
�'�l�I�=����A�c^�Y�	�S��}*k�璳T��V����xټ깪0�SG{Xƴ0b&�m�e�Or@z��έw}.����*0��wɩ��V��y����?�v��C�^��cT��X�-f�Ĝ,����c��?��+��a�g���.�s��=�2��^��s������pO��'%b�
��X�Kz�_'YǙ�s7g����c<#�X2*s[�����UW��#��٘YP%"��Mi�� y\m0'��^^���J�#�E\���N_4}գ�/Ne����,,
6N�#��8�Rii���\i� k�=Yy���UR]k;݊{������C��Hxj����>�"�Q�-2���7\�Ƭ����������h^���s\�������yׇg�/m��d�r�%T�#ʡ�u��01*W�������w1�*R�rJ�U��~61�3�m�9A�hvXW��G�Yp MR����oht���Fz��<���]L��r-��7-�1=�v�}�c�(?:�	�q�s�>*L�{��u�x�6�2H>d
=+�k>���z�xg��;c>>ζ9�wI<����0�Z����t�,M��YYBk�f��ʄ��`�WQ�/��>-�!�O��1�}��g�ۑ�����3��������pT�s�ݚ�Vm�>�R���f��&�]fd�Ug�;������feݏ���)ubp��u��v�W67;2vԻ���U�8��}���3�_Vu���G�Ň4[`=W��u�T�J�`4;z��u-S�w<W��Ny�~���?Ws��D���N�$����� �&� �a��f�P�i�^72{-�{^�j�ǵ�F�k`�e8��+�s�pk���i%��96*_V����������c���,=G�{Mo����+�7��~&����f�e��i�c��ς����\%5=���\ǘSx}��ax��nU���u�a��hչ�9_s��j,����KbHۜ����g�6a���
JӃb�:N��;��:75=�`v5��W�d�S���%s��:�lc���Vs�w��5BwL;�����΃�����1U;�L|ڃ|'=7b�sq����^^�;u^�'8���ɻ�]d{UvS��ϙ�ڌ� ��&��ܓ~�O���;�n�hv-f�kY���{<�r3F�V�}��ۊ��/YUr���K.��y�:���T�X�E�~=�y����Yk����^�Q��y�1q�:�������do���;3����ع%)�DS���d�z�!�E��e���=���׺w��b�Nb�*"����R����}��vomD����IN��'IZ�D�`ͤ��(4'-�&�����ID��
��xw�ې��>K�i2�#��uiht�t\�����b�μ9�6��l�Juz�A]����W�^P�Ġ7z�����3[o�G(T��;�8�e��!2|��<���~��z=LnF��=ϐ~�����3U>YՕ�K�"�*K>�I`�
D�>�̒��<y����^�w/�/K�75�6������8������N����,���� ����u\H�*��	��b����b=l1�~�P˴��}�da5�~jc�Ut*җ5�"J�=�B���֬�NA��B��~�����p�Ws��`7���_���mע(	jٚ䔞�T�و���I�J�n�Y5|9������:������d!�ښ<�a<_���%��W���g����y������E��W�!�6��ʰt�����5q���zH|ڻ�7��F��#�B��,Nu�{�NW�g)�����K�Q�yv����"r�_K[z2"��M^�P��	z���P�OK��������n���� 
��r+M��!c�2v�T��}�; M{Ƒ��[�����x�(��/��<�,3��ջX��j8�j��&ە_>�\�����#pwj�ey���t���@L���g���f'�ٙ�9��q���Lpˌɚ1W�T�J����5���:�fd/	�w���*З�$
[��Ӯ��-�ߗ����v��u�gMg������wJ������,�ύ����{�Gl\v��1noM��hq�d1%,[�Փ�zB5}����Ͼ�u��9�vN��Y��',y��(v���l�:v�e����"�f�U�/��M]Z]�-a`#�N,D���w�)Z�GK�g�?m�Y���*xs�:wk}��4&VlM@�_���"��%I��r��>����#5�dF�t��:���{�I��d#D�u���מ���[i�,Q�s��2��EL����Uƙ���щ�[��W�S��X�׷̴���j�Y�����ǑK�L�m)q�c��tvCj�������N��bK)���<��r�|�l{�D��|;jY�e]D��?A�wF[7S(/��T�'����o�˕i�s�YwL>��:������]�{8�����<�Љǖ��F���Q��z�����lV�n&�[��As�+��uG��#n�V�߽T��{xr��4O@�^�ԈL
��v�(/v\+{
�b���w���||\�ĶЛ�Ꙙ�Q;�u���>����[��>�*H]p$�ښ�w>�R޲j�yY�6�b�mC7w^o�A�{��xO��x	��n��d���������[����칊���w�=޷����~Sh�ͣ���Np%��oF�7����oc�5����V�0Հ�t�7�e������_M�OD2�Q���n־TцR���2� ��XH���Z�'���c����֩MS$yA�1���F赳W�Ǫ5+���ڪQYHD(��N,����N>&�����X�B�9�B/]�F��d��1H=�vz��ڿ�j���^1���h�ś�yj[s���#]��t�0��*.�1�KՆe@�����[�V�Q�c޳�� �o�c��vϣO��^�\<����c����t�'-�Q���}3U�5t�A��K�gޕ�Uћ�z�Q��ӓ�R�O����P��T��o18�|�'/���g�?�l��d{��S/;3׋�̳�ߕ��Z��`�CF����~'%b�O(tf��b/�N����S;��#FL����W=s���c��6�GI�=x'ȱu�Zo�r��~��-W������z���T�pz5����#��+�+�����+�>�Zn���FGY@�!��ii�rWj���n$���5���	�_�+1�1|�7+�k��U��.z�b��R��*t��	=�|gP�F^�
̫f������s��k����N6��9����#}q�)�9��/m�:vKeJ'@Q7�Ũ���I<"͞�HD��ۓR��$�_0Y�ҘZ=�s
�2f�`�1M�&�z���t�*:�uuJ��K6����jQ��ӈ��Abl����b.O��z]����Y}�c��0�\`�㭫��ƞ9u|W ��Gu�4�
���Eɣ�&�Ɉ��nfˁ�]Om�mn]Ś��0a,��_�����с�N�h�n�Ma��g����{�Ǽ���Ֆ�,ܴ��fu�MŖ8TZ����5�V3P����9�7��Gib��[M�n��b۩��&�xxs���vP�j���agM�wt{�<�)��ڰ�gd-�X*)rǜ�+hsKju�(y��g��qˆ����Zw�J:'y,���on4�1�Iט���;f�KO[�V�6{Y��oQ��$j���������4��z�L*�Ҵ�|k�Ü0�R�k�;��xк�yu��˗1�[r� ��w8�aZ"uw�����ϒ��B�o����]]��ŪzU&7R��B�P��2��b�����[y9�J����r"�L�wי���3��f�L��e��e��L�+�Ͱ�j�j<r4�u9��z������9x��V&�kzT��u6Ye��t%J��̐Ta��nv��q/�p�b��;ΡI�obН��N�e���b�.�vmrN�@�f��J��oD���5]�۔����J�
\PU�E��9wuu�K���,Ȱ���hi��r�˻f��݋�����5���sf	eBn^��ho[���/4r|6(����J�W�Tfƨ�V]
��:���E{�E7]⭏6���"�]9�S���Q��҉@�ρ���w3��e���0�y��w˙l��rF��y�z�ed�{�:[�G�����e�s:�s80�Ġ�AӚ���$u����Zi��<D`�f:��Y�H(��7�)�­��Q��1/7������U
q�"�5��Z�ЗWM�2��B��;?2��3f��=���@Q�x�v�S��.�>�1grC�R��+�]e����S���X 3q��A)N1,6�pnfٻ"���˺�iȫ����Q����qW0ȵ�T�պ'#�sU�4�w$Ήa[�����+��,d[�v����R�m�\V�;벇G�>���UAtg5��Q%���p���/Ju3[������4��W:Q�=W�s�rj��M�TK)W#Sw� �}hY�q}�;�;Y�Q��Ǜ PQ�nuj�
`Ϟ]�:K"��A{
)���N�ɋn+�R]����|�.��)��67v)��D�x:�Y�����\�x@�r%�(�Um5�]s�'��t���vٴ�\��iҖ���AoWwj̴�sU�i��y�+=��dm��G�G��ғ���ZOu/�Z�1�ץ��I�g �]9;>�I�����UzNKS��-���Ͱ���4��p��|k{v��;GD˨�a��yg$�;u�kYu�t89��������ߨf$���!��H�,b������Di�&wW�Ʌ�$I��0J(�5DID�R6�IL�wr29̒&��QΚ".�Ƒ�E�qH�wB���۬,�fiM+��`ܤ�L)FH���A�cB��4Nv�l�!�d���  (�c&���$��2�w[�$�	��DF�2$���@"-2J�\����H��2&00ƒ$��swn�ai�Sgu���H�I@IJ3*##���w@I�0���ܙ�JiP�`3Iw��i���r��#���"�Q�������l[�aF7U�o���6�%#����U�$r|�P����������ދM��z�\�	�(�,�FT����Q�����)N�f���W����9�{�9�8����x�q�����/錘����
�D�&�_��.�S��s�z%�CFB{�h���z�����\����{ۏ�u~ǝ���6��@�2��@�@W��|X�|<2'�v���1�������^�k�x���/��ПN�q6�jY�D���J�u�(�>�TB��J2�h�c�U~�.�҅�7�;ɓ���&�m���.݉��&���=���2bh��+���I[qu3+�<�S���c��������h���-ĸ�����B�t��%mH�K��=63�7&e��}O�l�-s��>�O�/�����Vgz���F��̔k�~�;�����!zlz������N��:�rE��]�Z��=����/N�mxU�Ox�*C��갎�%��[�r�ҏm!~ր�����k5H�^�I�|�A=C&���i�t�I��enUXcyW�C�H�OM��?V5vnL��׵�f��XXk��J��'ޯ���D��ui��o� ��u�FMz�i�	�r(v�l��~P�5?Z����y�ZN�`S>J��S>����eVȥ{��~;^XK��I�2d�U����3K�q�V�-u�C�'�%<�zOmԣ��v9�,;T~Rj
�s���W��΅:�X��m����tw�r:H���7}��:�s�SC�N�w��\o�n����x��+����/G�;���F'B�NS�hS��p���d_ʽK�c���)ߟ��Y�����]EQ�P�]�vah���/Qȍyj��2��a���i��Q�Q}��Yi��s���>��W�WQC>�$��~�x)�����s��LS����3�"x������0�"���G[���u��<�JSQدq���N�j���e��辒��1 �X��HXJ^��\��@{���X������i�Le���'=w�W{ٓQ,f<�zF��h��$�3�H)* �[72��x(t��Ыϫ6�䙟)�KJkϏz!yG�WylO���w��f����d`���(����u_�#���Z���u��o���Ĺ����ONxsYM?51���WB���� 9 q��u2i�e��6o��E���Ɉ���$<�u�l��-�>��n=�^�O�<e�̖6Iju
��t�t���[�LGZ�T���z���"Gf��G�zK=�K蛈�ͫd�vs�lN:WH�N���/+��g�Mz��+����kh[N����
��ܭM�}��kW��c�^�x,�Q#~ț�5u۳Na(�Ԋ\��l�B�gYr��v���w� I�f�9��ܰ;C}�������ZD��gif���5r�Ρ�g砀-�����eE�|Uz{�f4c��$G&�f�����~�����ҁ�&{������1��b�C�M�܉�!K[z2"��M^�K��1�z��5�EH�=���[��W���-��O"��sB�ѓ�#�������&��H�������9�3�$۠�cݐw*��'���5�[U9-��c���]�PO�������V����Y|dt�e��X�	�a����CU='!:�^>S>�7ݚ-�+h�)�t������2�kk��p=����E�F�K�?F/+�{��N���~ۄ�z�������g�H��6���J=\u�X|h�</�	���TtK#�{���Z@���^01ׯ�+}WC3AW�nw	��ʿ9Kr/��n��/��HвR�,eD<X���|��]����]���1^�h6��d���$2-�c)tn�Miϲ�6(�'W�C�FU1u2��>	�<�3��R<e��~;
1p[�kC�W�{}�w} =_{���b{�c�FyO��y|�?�u}e��4-�q3�XOk���2�D� ��:έ��`���oq����WQ{,��g���5U��i�Lj�I��އ���inG����,Wk-5M�{�m3��#�`�tWew�;|V9�^gZ\e>�s��{�I�]���A�F�u�+qZ�o.+7E�����[�_N�~65�>���;?j���<�8K������E{��{.A�8^OV`Άk%�b.[4��xlV�P�Oun����>�<q���ϓU�i��������;��=�1��'=��?���
�_�<�_�����t�wI���P�(:��#]�gT�W�&jw|���?�%:hRa��b2`�l��8��
����5~dyY��lc'��&DkZ�ѕ����ȑB=��K�4hlɎW�	�1R��F赳W�ǵ*����_/v]Yf��uv哺�Z�m�K�\G��q�!�4r	/�d�ς<ϒT��u�z7>�S�^ޣs���n߫���*F��D5C�8�.�ʋ��z�?��Ji`�|6�r�F�L����,���x珣,��]n��=�b<-�q8ژ���f��j �8�ww���N�{y���20�^���Cn��:n4�(z�(u�R���op��~�����P	=�9����{fz2��m_�%�F�b*r���>'n6X~�9U'�����{(�M
Qq�K�w7�F�[�#!��;a_*���b�m��s�m]�foo�@�f� 'S��6�	�]�i"-Ԉ��B�#�����rr�0G�խR���庈��OP�}g�c^�7�_`*ap6-���Y�ͫ����A���;k->��߽�1F��;��`6heyP��ׄb�r���c�����h���;ncݟY�k�$���:W���ء��KM�6N�#��g��4��˦#�j��u�q
�V�Xz���z9�Ƣ/\�r�N�ޏ]����!�Ϯ�˔IF��k�*��&��V<g�ثם��]�V}G�4=�8�Ń�0�{��x'���A�Ӳ]�9@����:^�;�]3b��8����{�W�Z�o�\U}��~61�3�ly�q��C��W�gP�﫰���NU�"��B��Pp�#3�N�pnb�e?N}m։�n�џ'���xşm�:�*Hǫ8�c���!���j��B��� s����^SY �Ջ���'�vÍ�QX	�g�"����Z���ǭf_w�	��К�O�;TH$�WQ�/�� L4!�����Y~����{��v�z�����[ZK���q-��At�O|9$�֙'��1�Obh��=���]i�B���Ơ��q1�3��B���6��_�(8� 7��h���o�Jڑ[2^�c��N/�v��+�~�KjE�,K����$v�[{(�7Uj��\Z�ލӺ˭����:l�T�(�Բ*��H򞭻{�O	��;}0������2�<U�<%U�1�B�g��
a��ca�̐g�ܻY�W��w�&� �/�1����.�w���QG`��E�?�md*�Ni�5��x���c���p�_��oޠ;�L���P���P�X�:g*����0��E��OFTd�m;�蠻����;�HvcK�o��E�s��_{'Nߦ�qm�WOE��m*[���j�t�c����8'��	�X��*��f��/2����,r��=�~;��^��\V{�������	���z�N�u��7�A��`/�v�vs����W�}u�lo'�o粡��?N��P��Iݳ0��)���ZDy��@�������>��a=��`	��-S��φ��|�����/|먬��Pۙxnw��w����r�{�m���&k�xC�Cň�{�FoN��;���Z�������:�(G6=:\zn3z�4��#JY'},m	�$�Lm9	��>��y����Z6���κ��>�UU���N����O-�S��|�W�ȵ$Fx	���R���'9�ɠ���<4gz=LmPn7*h�U�)�Gh�8�y�ܱ�[��9E�%��$�}-����<�@N���&�I�}5e��Ƶ#���M
��e�9�n�홅��Q�.�]��NᾹ�{��a+�A����J�q��P#��z�p�
�; Q�5u_lc,ws̹�}��h��t���{�9�y|�Y�ek���j[\�e��M=v�&g*�f�������WW<����ɳ�ƣ�(?-����w�G���1�'�� 8�S�<�Ô���y�g�1xk{�:��,֞���q7��H��ݱO�3�`�.	L�ȼ�3�n��Q7/ö�K(ޜLD�þȑ�7�w��l���-�q-[2�fK{�#�㦪�/���V<z��H#����|tn|�[¡�&��o��zK6�m���G�>���n�u+T��u�'�����j�#C&L=���UON2�ץi��zw�2Cj�_ɿY�O�oq�"gW2���SY^P7����� /\���sV'��K[z2)ϴ������wmGy�U��7��=�%}���sQ�h7. �k��k�c�B����O�GPM{Ƃ=��}������>[\
&�6��}�z-�_�yUy~��=mTt�f=�>�\��Ơ�/��=4��OU@���B�S]r�y�N�æ�-,{I�e
�e8ٙ�'�q���Rp����ٯ~Z�5]��w��e���J��bwtrP7�g�'�ʭ7G�(ޟ@��Q����S�2���,�z�����	�적�F5\a��0.FY�~��(B��X�-_+wd1�6B�n��f���Ą��u�9ׁ.��2��S�U�hc�Zĵö *�L��T.���l��ډm��,��T�G����ڼ��rz��jK�E�Q)+����V�y�O�=:[��O�4+���eV�v�0�.�#^dٿ�h�A-�י�,�)ﴰ}��
��^02z��j��ڸ�z���6����Z�W�1z�]#�p���P�b�g��9��4<�K�b�bAwR9�~U������&�gm��{5�g>�L���d=(T��S)���(4F��q�/m��O�g�h~�/׃\x�z@[����qϥ� �e��Q%ј��aӹ��v�:�j�T{~�g�E�,)���ߨ*�n��x�9����|}�dg�U��%{� ��;�\Ƕ�?Mb��Fz�������џ�"���I\���#OS�Wɪ�3����ѭ�}�o-�<n �� ty���
Ȁ_[���λ���)��.}�f�c鈹�T���oVyV��X��({[h=H��'�{�ED��n 1ݛD.]L!r�=��y�Z��7}��u��S���f���f� &�О�-lɎ�qb{F�=�����8�{�|}����t�ͬ�=��t-��.�ˈ�ƅ�.b�B�tѡ�Izc�����]�k����8��NĝB���)�g&��	@}��&hy���|5(/Nv�e�Wp�(�;��Y8�.��d�:�NȎ\�����k�f��7:�Lv�&s#������sv���7.r �V�&�0�;Џpܗ&\|�k� �:ǝܬ�!�������C�ƛ\�oR�y0;�7x[����X��w����]��=I��0d^��ہKՆe\a��읮0�9w~@p�c�Z��a�0���W��u7��CF��I���FP|��jQ��{�|D�,uv��v������ј�tzK�6n5���YC�j����-f�$�c�k�S�	��S�����;��U��'?D��l�wS�t])�N�`o�~�2RyC'`��H��*�_��KG=|}�i������V�0��fT@�"��;�9��i�w~�T����C�о^`�����:�{ҽSct��<���H�'v�����C���9�A���;��'�S��`x�b<�B������)�,��hxvDK�B����Y(��Ih��o<"(7C-L״k�6S�FwM|���4=�tu���f��g�y�of�}^�/mrKĸ�
o�چz�r]�J/H$�g ��B��^����ԙve����}�/�F�C=~�p��۝�$��M�VeV?O]c�hh1��DLl�`y��%?M%8%ķhhϓ�[D��y�dB��;-���rf��@��y댅�d�v9�X�qz�ХjZ]K�Ϸdj
�?�B�v��6fm>��"� ܂'0b��B*K�[ЁĢ�&�R����Ǳr��Zw����wLW�nw|�j$��n.w��vZ�����kb��h�ٹ��[rlZ3��[X4O�n�q�;�q;qN�y�|\ � t��=�bF!z�!�m(��W��0oE��ޯk�eۧ��f�Л8�Bhr�,�" 5P$�^��!��ilW��yU��^oFK�q��[�!���}�D�<f㉦�Ȋ�n��ܒjkL��h}^���3}dӏlq��H���/Hl�\�C�m_��zP>q�^ o��_�����LvϗX�`M��[��!H3�>96+���RS9G����y��7�=��F����f(-��x:L�N)zzz�|S������m�ת���V?F��K����_nU���uXE�;M�s^���o�D*���W�e�����BT0͛��U�j�mhw>Ӣ�Γ�P�n]�b��{��C��L��r��+��G�?(ޛ��Vy�>8�T��`���P�a�VW��9�t?>�
!��UВ��D��� [{L)�Z��/NG���S���ͺ�t��a�S�~�o��Y�ں��4}\}Z'�� 'd\*�/��ü��'�%�/�󮢲�	C]U���������\�=y���&RW�v�Щu��Q�uӝ��<�Ȯv���n`�+�VΊ�h����Mu�9BZP��o)?�Q��5Ю�MX��`�:�����:���Vxh�|��[��0�|B�F�bC6M�iH�(u�q��q�ǨIw9e��xE^��+8M��(��f�q �Kӝ�A���@�K.�o4q8���Qړj\�gdu�+��<�ǘ;9}��8�3���* �&�-����S����	ӊ��ʰn�P��݋��9��*a�ޏ�A@�q+|8�&�m��+p9���2r���Fc�M��ئ^����p��|VB`��h��ѥpD�ѕy�wR���|TW�!RvS�-��DQ����2��Vj�#|��։�-�R ���(�yg5�*�	Ko\�u|�=��W7N�����rΦ�x����̈́_WH�2�4*eѓ�a=dq�0�ۥm����5,�*�aMfc�;Tb�SAos��C��p,�b��e>[5���,[�b4v��1L��nj�z�κ$�7ǹ�`PkG�_>��k��M;U�"[��(�J���ʼ�9s���Ob���ك��Hj�\�M=�j��,ߋ�tux>x��lbS��y`Ӿ��WA};�-+
Ӣ������8��W.,���grc���*�AKq[\i֋�kU����n�d!f�s}E��fcΝ�)!Ҕt�:�Ӑ��7L�P޼�yF�,�������8M��.�-�T�����v��ӲT������\�X��Ci���n%��̱���ۅu����pu�˼��"��t=R���g��l"t=wH��mZ�S��퇢�m���0k����՛���h�J4��Z �;�f@��ӷ)Mj�7��זjjI �Y�*��ef떇S�#Fp�ě�qS�l�/���������^(��g���J�k_PIDi���7dL����S�oo"�'}ڀ+>��K]�kqPA4n�Yb����r1�6���l�<�Kǅ�������fgK�(�
Z�������ø��*EvN�owS`e\�ph�-{��	ky�M{f���*���v�)��|��#shSz�G���> r��M������ܡOUܭCcB{�N;n�;���ZUH�&Ρ�4�ai�Ǯ����՘N�S]B���#R�X��s+�5[�w>�+��ҳ��k;�^V�7es1,���N�:�&}�^T�[S[8��h�X��`��/��.C�%�C�[v]D)���Ԯ��ub�b�Y� �y�:ղGa�jB��N�Gab���K�84����oVH�?�`���=:.�C�K�1�5uԚ��Nk1}���f��Z�F�X<ð�Mcs�ʋ�ULh����`)"ݮ�Z��.�s��� +�kG:��]�Yl�ʆ�x:�Ϭ]>͓y������t��(}T*�
���JI�BN��Ac&4!1$)��M�D����@��#��a�PF��6f�$��F��ݡ6��(A4�����A�W,PH�(�!Rd�\�]�ጛ��nl	�۝E��)����.������*�0(���̉�4b,X��]۠��Z�˔�k�4F�M�EQIh�D9�]ݷwwu�q0�H�bQf�r�c&1�hđ��h�#!$\�(�ZScF5\�ݒQ�����ww-\�F�i��ݺ��"�!�f	�"�;�r���(L�s��I���Di"5ˮ�t��+�rfR	���LA�%IF5wv,d+� ����o1���jıw�[R8ۘթ��` ��6��ɄV���9\�vu�|t���^s5t���z�p�&���͡3���3�Ek�^KN�p7��� g'K�վˏx��Z�����cpz���|������Z�Y�5VӤrՒIhL�h'#�)��(��_{�3ׅ��y�q��Kɾ��o���1���^��2��Ƀ�r "�}*����'8�h:���<4JJ^�蕯=WkU^ll�����ơ������(�YaX:@)(�[7S;�=;[E���h庅N�^�����}�G�?N�����w��f���3`�@M�K����vwu(�U��PcQ�{Q>�mb^W���Ѥ�o�F�޻�)�f}<��N�$�Uz�T��3�`�1�`ݡGN���9��C�y�q�kg���mע*Z�e,��v�;.K���Qb����[��,{*Ot�`�*�_��[¡�&��m�|���L�r/�#F�=�ԑU3^�ಜ�ȇM_���U&��a�F*�'�Q,��Ox�=2|ڻ���R�W{w�oO&h��xFwD��(�n�M���NYOnމg�k��c\K��R������va�& u�%��C��[gH&��ۃ���b�;Űi�it�6s.�z8��N�=��l���v�U�.]�I�G-��r�c�M��S[�̎�%�үL�nގ<�FxF�u^r�h�T�͓�Q��".7Y�6%SNk7�oV����.�+�:��F��T���5Ke�f�ƀ�<�!���Ј��O�GRu�[ϋ��)��ʩ����������[���)���3>�=V���F��nH��P'hG%�6�5�u]c(�����(�1��a��x�Ų�Օ�`jK�M�7��f�Ԝ,��\`�k���������xn^WM�NtY��u+K���(�ap1y�{����ϧY���	q�V���ۣ��*��{q[��['N���	�
�}GEӑ�7���K��k"+�v1P�v�`%��c�ޢ��+ˎ��Y��>�G,�)��3ŉ'����2�4�,S�z�>�A�=��\Pʏz�3NW��_8uЯ��go�Ka����)3Q�N���:�(EL�}�h�m9�R�v�T���7�7���������������D��s}@>���i/'�q���e]A��4v�>�4g�#�#����f����|���\�S��>���; ��c��p��3����v����ъw�w2�s�6�9T
�)L�E�ȵ���#��x�>�1��L\��P�-ℝ9���>.'P�Jǚ�-�x�"R2;���RM��}��c���g�M��z�`�"5��c��#���e;0��d�^�+d\�����;�.��Ǜn��lم	���n�c��.���:ƒh�$tmo|�Ҙn������ebcW<r���o�F~���(!Q2Cs?J�kz�<��l�A�u����/l�4^���Wz���YΕ��~��BW�k�sD{�@j�rb?Ox��oY��r"���Q���G��7�����A�t&�Jh�̘����Ѡ�o�>���j�a�ݮ�6����\�/�]�Mω���c���)���Zd���R�x�S[��w���u.��_*�?7߃nj����=O��4�342�ѷzl̩��{�F���wc�h��o��>����.^�~/��B�WC�u�a���h���8������zx���G7;��w���sܟ�K���6�t�~�;�F�����ܾ�jL�L'�f�u���U����q�е��Y�]�l���LN���·'$�إ?���`O�~����,��33w��yΪC;�ν|�C�׊]��0�}�u��wA�y|��d֛�r��`\>^��'�{�1jw}�z�A���c�m��Ҹ�-��[�%�E��e|���'!����/�T	�)�q�����2C����;��Ǔ��ȋ��e��3}��	+H#8v�n��	r�@���;3%�r8���<���T����}w$U��7gq{��G\n����,K8�p�iw%���Ϋ�	��ek��*sg(oo�����'V��fI�]\��;?�P�al~c]X�?zk�,{�U�����з��Ad\�'I�خ���k����E�e��g0�E��5�K��aiٿ���y���>R��^����6r�_��ׯlo��/T�Ӡ����0�wS-�]O�3�;��{�;>f��1�/�����9�T��]gfH�����^Ӷ�<xDF����`y����S��[u�n[�4b�l*�=QF�ϒ���J�{��#���v��l��>. ��@�[ Q�^SX^P��o�6{1/=����U�y�z�t�˼�����a4��O�|�:p�jY�D����T�����o�8M��Ukv^xLw�oa	���x��&�m����۱5�&���$���}����zoӁ��F6�Ȱ||�!�ː�vڿQ���Hg�x��k@�����FធL�s�!ݵ�!��y4MB�z�ͣ���x���C���F��O2Q�mDc�5���v���}��:s�/{hiʰz���c���86�ׂ�����]�7]VM,���55�o�@Kb�p7�Ż�:��-�g�����;S��乜k��iʄ*�;^��w������eT�B�ܥu�mp����F��YB�&0�5Z{_0�oG2�[V��ub��YG���a��{SK9��}\{9��.�^'e���Z�Ӆznd���wN�ȱ{<"r�u(�g�i�q��0Ս���tK:Nll�;�S�^���UǞ����[��c�=�}�F��Jee��Xh7~��x�	���z�O�GR����ي:�׎�N���
�=��� =��˭9�9����R�~����&v��0?�!j�����Ӏ^����^�謪�qEx�q���֬�U�^#W�yN����н󮢍��7Xij�R��ʷ$��r�3�:�Z�����K�*9:^2�a���Q��Є��7��,Z�א�٪�����g�A9aL��At�����L��hB΋<�us�֊����n��:�s'}ȯ|��	6�3�e�����<���W�ulL��9�*9f7P���L�X��q���P��]�棎P��_J��q�,�2�,D���,{p঺V�g�:�kѲ�z�w�{4P��{ף>����59_?-��m4���f�����t	KF��B�w��v�lr�O��|r|���__?\M�k�/+�����u���S���\җ9���mJ��ˋsU������W�}�haT$"Zw��Hds��wFF��E�T��W]mN9�Ж�}��֞Y�}��v�z�v��+�wg�3Es��{lNk�\�����Bj���1���i5���vN֝d.u̮6g-��2�ahH_�
�G��@���}X&�$v�[��\�ϋ��mע)�1�(���OZ�8�n������K��LFO�[
��G�A�P�d!ս�ѡ�^��n�3��օ8�����_�~F����ʓF�d�m���*)9�_z{�}�jc��	#޸'!5�_��z����Ί4�#�B�Ƣ�F����ڐ��NY����t�����nJ4\�n���7/������uJ+��54ܸ��5�^41�!�;��"}�:z����3��@M�ҭ���Td==��C��T�<jOM���fܨ���r�(>�\����}y�83l.�������y�y���ڇu������7���^�[	%�&��q��z���<���#��9k�Dt�sԻӳ=���u���'_�;e vt9ɝ:�F�0������ix����15/|�L�������9;��cr��Vy^5��؎�%�o����5���yOF������~7�������N���"'[�|]�׸�>�Zv�����2��ē�v"��U{���ώ/��HOn����ц�VVɜʊkP<�m`N;4�ym�S�Γx-�/,��{??���00|�g!-��"��w7�~�s�ȩ ��]��wݢ.�Ȍ�9b�D���}�w^��k��B�v%|��Y�A����w��pޙ�޾Uʲ��F�B.�^�����������"��Rf�$�CҌ��a+������y��n�*,%.7��Î�-�ǘ-���;)��xn%� �mK,"K��x���ݕ�b��� �#=Ƃ�q��]�'u6s}#�{} =*=��mǽw��\L,\�ݷKRb�ߨ��GH�5'���P#ų ���^ۉ�n�9\��?H��;�ؗɤ�y)�>Ɏ�H�R�Fm*�|m����:Cu���
��[���K��`Dϟ{�Gձӊ{��F�j�^�>>��m?\N�z��Eê�eI!�H+�hK=� �/x�C�x�+����-��+����W��� ��ώN2z�B�7M	�2�ݙ1�_�Fv&���D�����}X�Akϯ%?NG!�ڐ��6��Zn�O���o��n0
��ˈ�I���/K����/��v�K���`�O��{��;�n?S���H���ΜFc���Ǩ@r�ޙ�{å��vC��=�f������WJ�M���s�=�z��X�uXo�Ƣ4-�q9U��\�:��Uu��Z�Xlw���'�����G82]�S��� ��m^�3���t���$P�H=�|TϺ��m�����A��,���v��I<�Jz<�^�E���<^&۱�'k�<0��.%0V��.��Nm
ST���� @P�Xȧe�a�W��/�a5=�F����++�n*^���J�ܾ�x�k�b^T���n�����q|5-�H�;Gڪ���޼�kƼz!��vt��hՃѫg���'%b�S_}鄏��ڛ�:U�8t?�%��_'Y��9L��c����������^[y�����5�G�������:���w��3�P���B��p���+}u���{�Ho��"��):�I�^�W�YS=&���q�l�����i�>�
����^�c��v��d�����8C���cl�ѯƻ�I�bOx���_#/L��s�r]cU}1�_�����q���PZ�M�����#Wۊ'T��.8��(UD�1��u2���S�L�ɦj�5����H�|s�3Ѣ�D��1ގī���}p�!�o���3��p���A�B���.�S��s�w�7�&��'v����Pq���y�\??:z}�c�(?:��:�!�Q��� t�d
���)��E��Q�w������/ZdD�;c������a4��O�|�:\�O�;P��Ȱ�.��3꺳fX�o�C�>x�ˍ~�|]�v�꒍3wQ���ϒ��ۻWB�wl[�ƾH��q]�bŷn�0_)u�s�sb"94��(j*�Lv�6�m�P_�2���|���P���t~�v���4�N=�X%�\���v��/�4�xeN�3?�����9`�j��ŧ�la����ɸ��]]:��&��e�Â.eͰ���-���t*d��ɋ2sF�蹹�vD�ﷶ����.�e8���z!%:��������}���6�ƫ	;�����^�Jy�#^=�c���R�C�<�D�9�Mno��f�I���3ϲ��vxL�Y1f��]6j\mɸBNY���8T==�*�p>:�ٷ���7�0�^��gv��3�Z�s�')�Q��x�f	Z6a������t]�҂{78{��/c�ݏ��WU\8�����5�Ҹ�Xn��Mߪl�9��C�MY���`fn���s^ѧJ-i.���Hq��ኩ��'^^����וC7�>'޸�]�� ��@�9�#�,r5M%f�9��y8����\�1�rN1��s���v�e>�4��T�������_�=��t�qW?�6#�<,(���
�t��S�MZ�~ya+�{�*�=��[��u2�ET�
�<�ϔ�Ӑ�F)����y*)g~j�ff9QQ�Nf��q�N��}g�.�ɛ����9��r'k�wtv�m�׌d��Q�NF����t�c�7+�T�\�4.�7���M��a��k��R������E����7Փ�V�������W��}ڠn����1dcou`��7yum�.�+�~,�?��x��]G��
��/J�L� �c�"ĕ(o�S���78	�8}�ݹ�>Gܖ�n�o�n7LX�k�W��o�3���=�k;�7E�x���,#@I������[{����]Y�XKг٢��-��b������q��؛8�A�F6 FnxZ�`�EU����C7j!�4�Do���BOv���z�Ӟ������4�B�)�H���\T�d�wv�� i�-T
����`�|ioT;���G��|a���ɶ��7rnV~��F�����$������(�5|?���k��t�*j����m9v��}x�}��,��z���M�dqR���2c��Bӌ���Y�γ���J=�a:�ؽǘg���Ʊ�uH��h�g�_1�sQf!}��F�������W�}���ɯU��ѣp�$�����S��E��R��5M��ek��k�c�F�FN�Gz�nL����\۪y�S0<��Yf�9���.�G�R�i��9�g���:rsޚ~{d_G�񎧷I�_`��;:���y�����|��	�d���#�;�+m��]>N�9YN���+*� �޷Mji�*��ǯ���[����:�N��t�ve\Jen����X���{���k{m�d�s�c���<�N|��yl�;�U�㎺0h�>�\�� ᬻ���[����R��pb��Ҁ�)�{6�����nL�nLt����g
h&�,��b%�-��s���Cybܜ��o�PU�؆-��a]�E��W�鑒��QP��F�3-�ҫ�����ú�\E�kC��Cu�����W�sg�&V�]pY�T�)a�!��C�-��quCb����J�C���-�<���]Btw��E@��ּ+f�Ev����O %�f�G#zʬ��g��G(��fpFX���8��\5t�����(����ۺO�������!\����V�>G*����*F(O�g�ݹ��(1L,���u�K��VWn������m�5gc(�i�&p$���AS�\ov��a:�˰�;
�+�[�^�;4�X	]�`�'.���Q�L��N�d�D��lOk�8�Z�E�u��#�U�.�*�)�ܳ+�:�.K鈇�ofmjU�+���%=�jVR�Yz�i�,dx��b�	�am�:�L�b���4e����񅵟S3�)7������\:��7ٺ2,�F�0�Tb��K]�x-)�����T���N���GsX���!�؋K�qyX#�6m��Y>��������7��}��s��r�^���SDQ�`��q���vӃoC��a0!�]ȵv:��m�A�M+�E6��w�r|Rٝ��ж��7������6��v=�p
��D���N|&k���Ŗ:/v���Nunj����A�inE;�ib��蒬4�LZ��0�w�VS�9u^������E=F�TǷj���E�n7h�Q�d�`9��.J�۱<�k;l�W/N�-���X���bb�����Q��
����L�V����D�v�y�f�H� ���:�neλT��U��Z�,�ڽ�e >��2Woƕqo������{���&q���{;�ߌ�Ecc&uj�*=��B�94�X��Z���ե���s���x�p5a�,X��Y\��5yȶ/��{	�&��AvE��'�6�9��mܢ[����u���+}�����x�U��d|i�wz�{)�Z�T�MvѹWϪ��Ν�^���J"��.,��M�o�YT`�̜"�&�|���U��X{�y�3+�|��e�s�RU��6哓k���w{�j����Cy�P�f��8m�~���u�kx�I��@H�m9kH'_4{Q	J�\�y�n�|�u�ע�8�I.�COU3Q.f�3v�9U����x ��&��m^��ѦF�o����3��Ý��}d3�8��k�X�3`��/gmc��nHV�%��g+�f�m
S6r:=���r݆ �3WE�����w�������(ыQ���+���\�Nn3F19�S6"I5MI�I\���������F1FLl�4E��4wn�m��]ѹ�Wuus��[�1�$Tch۝	�wsF6Lb4c!���$ƍ�5���ۖ*5s��ķwDE���HF�H�lli-ː�h�5t���h���j(ɫ�,\��-w]���WwQh�b�s���F�l��.nr��6���DjMAr�`N:���kr����LDI���Q��2X1�nc\�Δ�A�"�F
La4��(ѷvLW.�Q���ɱ��(���E\�0S#��b�\ԙ1����]�F4�E�S,�c^�z���������y~��^��]����[w�Slˬ�X�=�M5�ý� &�ۣ6
63���wI�af��$o�����L�\����?�ô���LY�x? 5Hw�^���I?�z\k6$�b��k&(I�F��=V2{��myc�l��<}j��H�+�1}�y����'
�6�3
�tn]i�Xu)�Z>�1�j�f��M�Z.�Ò���壥S_���G�[�3��z1�&�xY��cR��=���DX�鳾��cj�`�԰��s3�;�����3[n�������;�d��qg��<]��k�ti���l<��+�+�e(�p����)��V9��=T�g/c��^�詔��}Rj#�uq~b[>��ck�����ތ�$�O������{/8Z�%�"�O�ZH�3Jg�Y�� ���f��0�r��Ga��Q�q�̱\��;�{9Z����^�~�3�������L0'��H�<W�Z��M�Kv�f�V��̉�H��t桊F�]x3�z�F�:�o�zp "�d��@�{Ǆ���v��;�\j�s�'
$y��^����C.�8��}�k��	�|�S3�$��i��#(:�TP]8ϟ������͟�ft�6qMʠs7,��EU� �-V���g:�w`I#��@n)I���݅q����}�4f����S�&N{��aujr�!D�0�3��_;�J�J��醫{N������9�v8Uj<;M��q�v�ꛏGb9��)�&�5>��1�m�1����E�[�,�5��͡b�ۡ5�SF�̘�O��b�t�ht߇x#w>�>��f��jU"5.��M�%��.#��ΐ��1I>ԥm�zt_�s�	^$������q%3j��;�1��ϻ�R5ޗP�N#�3��A�*�N)��yޓ[x'�eMI� �\F��9�����q�ᯖ�\4�U�}�@z��W��pg+�5]j�h��#>�g�0mV�j�G��)��t��W�F��7��Ƚ1�fs�2�����gn��sK��N_߿P��S)��~�vv�������t\R���B���Ma"�����V��i��u^�	���~��K{��b�ٷB��s,�<�>⇝�1�ѱr|o�WfAr�XX�vW���ޭ�����_$��j�0�~[��쥦�l�U����w�7\_gDcE�g�6\�� 5�c�t@�@W'Oޚ�ˇ�����]l_�W+[�b�(g�f:�\���K*N�@̎Re᠎��4=�8�Z_Lq�s���	nlp�|��ҙ�N�X�*c���x������S�����{1��,b���������ǖV����"�ډ�Y����"q\32f��1n�-a9�OXΫ�h����N��/i�<g��8S���G���	D$83v���Jm�t�2�O
B��ksm̉NPV���k}o����C�`��L�D�P�
gHBe�ӟ,�F�5z����T'���o}�>]>��o�3���}����q��d��v/�E)�gi��,�)>˛�x�_o��s�Q.uӏGu��xc����C޻f����p@N��H-�5@�c�Nc�"�=��<�]��9�묁G�kb�[�����a4�>4�
�\�f���C۟�|Gma�m�G)��胙PGτ��[�C������>�5N6�DN��ǧr�ڜ����2�mIb���ǌ�ښ3�����d!�ڜ����w�ez����=6�-���s������O5_�#�i�r����~;F��5��ڪ�"�x뜯_R^ջ���2h��9�C5X�Y��\5�`Ը��pc,�_�kNOx��T���T�4nIkm1���Wy�ѯ�����G��Y��zGe}^��/��⩦�x�la�|9j��vq�G�_޺���5vؿ��i�W��Xh7~��x�	��{���U*�S&��A���#5�#:���]Ӎ_<���`SY�If%�meŌ����n�o����d�aę��_=�Mb�u��*d)�k���%�v�!�����:LF��Z9YArI����㿕�P�s�u��IPݭe��r�X�cɵfi^dF��l�/.�<}�GF]<��UN����~SC�w�6�*�g�U	��{rDӯa���d��#�cH�J�['(ylDN��
e�f:eǞO;�����u�O��<v�ӌ]y�F)�*�Sd�z�]��I�I�}g�b�P�+�]���.��ʋ�Umy�q��5��7}�'�����QC"�ETL��"&r:�S/dW˦8��L��8��(��v1���术1��g��島���¼V�f��y��|�R�
����%1Wt��Ys}�]��2X���Ӌ�0����Q�+�Pyc�\�GN�w�ޛ�@X�V<��`��6cӒْP^�4P���^��^�3پ��\G����A�*L{.�:�!�/e�����p�`�@�AJ���3"����&���!�Ay^G�!��x�{}R5m�xݻ�.ڭ�{�/��_��׍�R���$a_U�l�V	�Ɩ�C��m��||�0���%ٜ�J�jN<'m�ܮ�Aw�������y���揹B@����&�a�2����3mצ"�T����<���g�up�d5,���or��y�2)��[:�Q��	yi)|VX��R�uzw(׳Ҧg�k)Q�����r�7&f��j:��yԖ
�ٛB:�|��=�Q�S��t�,]n��J5�8��_Y=ג���ǱKd���z�W�V�⥣�&;h�P���*+�r̘_[�f���m]��k��ndw�m]ы�7�"�ޟ@�d3B��Y�C]��!��#�]����7�d�ph͏T�PӞ�U�?g��:/u�(�9��[��5�^41�!�����9A�r����бC}�}����'��6��y`b��/]]
�4�߹�fjڨ��l�z�rz
3,gye��]�|B�ж�=Q �H��v���exT��ٯ��(W�+bƤ����.5��W	�L��N5Mn�f��<���R�ϻ47s�o\�f�����u|��cY1�<"Ec��w�{�fCSAf,^�t�y"�׫����^�hy��NF�6o�dT�s����诂釳"����LU �$����7����+ycqֲ"�:l�]�נ[�K}F�̃�Wp���9�#��*��5x��Y0�z���ǨD+�u�69��ۥ����zEs�I�k`i��pv��1��%��I�37���tu�����1-�X�C��:�xlOZ���DW�o. w���n�S<�b�/%Q��'�)Z�j*@���X�E�FӅh�a`K뗗�K �t
b�����p���uS�Rf��e�S]��pS��'�z���G'm�I�v34&m���"m
�f�>�K��(�<�ZO�D!ZB���L��Թ<��;`�U�t'��P�(�FIax�CɃ8���x�9�����&�2��&"�gquj{�#%�~�G�[ ��)�#ґ�3�x�m���ݠ���DW[r�����^��Y٩����x�y����ql�pp!H��{Ǆ���/?	��7QY5���}k��z���<��Ȳ�)��x���:�f(rJx֘���^J����l��eU�'�n
:�z���s�_�á���E���f�.o���B�&�К�4kfLv�_nH�:�nJ�޿\従�0�����ޕC���W").�иM׉�|=>|�E�����n����+���A�Ϩy,��~����^�Kf���>�1��/��T�x�z���>�h�(歒��:���:�o�����d�`��;8�^��!��ﴻ;�Hw���mv����a��+~)���{�:>�������d�lw����6t;�V���zN��+���E�����Ԙ���n�WLm��cY��',~�J�4�g77�?�Tz}JW�q}��ں�rU��D�fm�#�/T�?�T����U���F��dR;)2��v��N�L��J�2�kuxآ��eq:JEy�X��N��:3��ְ�G�Ӵ������Y'8�������	R�,"^��k��F�Z!��E�u}��tݱ�Æ�Jkb跫8����띈�t����]���Z͇����:�(�?ɝax0#+ɶ���Sß�{l{q�8|YcՓZn��{LN�#Uy{ d:�s��ա"����>�G�CՌ��Q'4�=�V9%c26�3�:�Z�7�9�D� ���:~�׮X�?]�ó�oQ�<���O1����!���A��$�_Ih��(ϑ���	��>G��2��:89�A���aj��rS<����-��I]3�H�w�L�1Uz�.̳N�e�b\�q�Z2��������<^��}!����w�s[���e� ��B���2|)�� 㡮>`ڙ�|���՝>�~�N�q��mv3|߶����p�,��b7���)ˏ1���3��4��O���|:�����mZ^z��~��k��B|e�B|9ʖx^�ai�*�fs�}�}(߄^���@�'�_�L>[�C	�R>��h���o��h&�M��j�:�bG��i��%;4K�D�nu�x���!�ݴ�����s��9���jW�zr�ς��t,�D�UfV�1ԯ��)f�����f�=%����qY���}��f��W��h��W�u7�mq��Ar��8$�l}s'A��̕�������e�uٝq36��J�� %u+�&Z��+j+,���+���2�V*���]Y��8��_���U��+�=�@��'�8T���4<{��r�V�(���Z�u�ڱ�,��J4j#��\B�Y���p�͚�0�\��5�Z3..TW1�2�^a9;��,ut:��uH����r�NkS�ޡ�
�H%Pه�kCO�2�H�7�KɌ��}(�a9�9y;_z�:3e���-�k����>�Tٿ�����������Ob��=��Ⲛ7Nt��c¾ܾ�2S�"�/N}�4=];�3��ܾ2^���L�����:N홅��ڇu�Zo�+ī�`	���qc�Z�_$��eT���T�����F~�����;��B�5���:N���^V����o��P��}X}C�05��Cwk�Ħdw�ݬ��<��947z#��b�κ�d��e��<�L�H�����,�C!L
�,��e꺳��"�tY�l7-���h=��ӟs�ƼrԐU�P
,wg�N�/�j�(�[��=te�4���nT>�.�\y�>����q��5����Y�Q%���/Eu�aT�d�~��d�*�Lw��Gxy''��w:��3c�P�E��3xfp�S��m<%֯oA&�&�LT|�!��j�WIG���߯�<d%���$�Y�2]��.�[ˎ8�LI�9O7T|fa����W��#��M��8�{���>Q<]µ��#~�<��u2ٸ���n�P�oױ���<�q��b|i�t�F�>���&�=�.s#o�Y���#I|�.{�2;�q�'�m�_ǭ=9�b/�{_������gZ���{fFK���U���T�o�@	�Ifu�K�U�	��{1�<��U�f�e�V�z�^�jt�i�mh7	��mת�f�UIb�Ijl�:�
���bȶ;�K�%{�63pna�\1��tٰ\�%�f���U�74�ǀ�F�d�mF*�=8ʎ�Cl����Tcwy������^��f�*��;����x�b<���Y�C]��l�{�~u��^�+pҥ/b3�9�ӷ��;e`��{q��;��E|;�CR����V��F�����K�W�ٝs�6<�-�5�s��[J�M�z}��S(z��5�ÿv5��ڨ��Uc��3h�Xo��#��^�6�]�΁*�A��[���0t�~�fZ����V^0�շ6�97��ٲѿh�L�[��h���+h�/PN�"0�}YU��d�׏���og�Sҝ�e���zm�8�=�d,�tq�$�%���cZV�Y����p�.�Y�Z�{�Z���x�'Wr�_q�yծw=��,��p�7�7%ms��	#�����.���'=t:uv�(^-�����0m��C�؍���%m�{8p�k(ɿF�N�~�9�R�X��q�2=��[�7�<:!�;L��=(;��:z�.�a{�曩C��Ѿ�����X���l���9:l�T��ڼ"��,.���c7,p5�_o����Sװ��X�2Ͼ�#�h2<�K��~�
��&��Ζ��<�H�ϲ���a�g@��8
}��?=�$�5���4�qL�ogݔ���an�/�Kg�<Ӈ�.��^����b������:��_�ڟeu"@=�ug�}=.7���%^�?��#�{�zhM�9o�|�0|���c��dq�%� Nz"O?�D9�5�3�����	����{�km�`Y�vmEq�F�{}r6���[/<g����� 7P(^�)O��wj�}�z�������{�^�_�����+�s�K�BnZL�p���v��b1]+��{��Px��Ѧ���/Oi��XKz�|���2����d��덁s�t&��8C��~�d�S;l_�/�-1^�9��5{0�;�B�N�Rn�����������u[Z���[kZ����mkZ�ƭ�km�kZ����kZ����kZ���[kZ����kZ���{kZ����km������j�ֶ�6ֵ��m�k[o�mkZ�ҭ�km�j�����j�ֶ���Zֶ���kZ��mkZ�~�k[o��PVI��R4�8
�w��@���y�d���^���{�G� �$��T�A"�f�4��B��Lm+Z��6�UHl��k�ݻR�e���M��[$mk}��5���(-�i�[m�%6�[`�l(�4ȭt�u�Ly�]mkAceA)l�T�+l�V�4�L$$!R(U36h�J-Q���Դ�g��-6�' �(���� 7p�:6� q�@ �t.�+Y���H���:ֶ�l���I��6�D��ʁ�Պ�ygA@��y@(( ^{��A@绀(((�7(�g�F!��� ܌M�k[���� x x:�ـ�/@��P���� ��s�� ��S���]�U�Jm���Q�o^�u�N�!k�mպ�c������3c��ڜm��v�U*j�]�i��+s��m�I��34�n;l�nݻ*JkU6Y6Z`x��L&�n�uwU
�]f�6q�:�Er����e�-˷v����5jѭ��\�K�ɃU���m٪��Y��fV�h��ʹ;�<��v�Y���v��띻tj��mۮ��U5f��n�λ�ֶ�vӹq�����ܶ�ۺs]�a�]�5�ӻ;MBe5�f��2��ok��WZ�Jղ�WwnZ]�v�݉Zη]v�N�sWZ��6�ue�f���wm�f�*��J�;���hV�6Ͱց��  �<��n��7(�kn.�f��Zk�]n�c �v��.�:`)�s����ie�l�kIZ� R� � �/&�]�J(w]�JMۀ�CL��Bwn4�2AV� ��ZԪ��1�x m���.� l0��fUU:����j��U�`6�V���  �  ���JEP� �  S�R�Tڏ�MCFa h����d%J)�14�C 2� �E?�*�M4� &F   F&�*H�M �j1F#M43D� �"R�MF 40 ���\ytۧ�>����,1�=-�����yV+i��sH�I�����<"Hr~T�A�I$D�		B�a�S�R��IR+ؿ_Ο����Y��6C��qQ)BE8APT$��O1EP�D�H�7"�*�~��e�m��0)����ww��"HI��m�r��^��G�6Q[l��gOT�T��H�Hk�`�_�����?;z��ݨ����C.�}R�\X!�ك�`��:��ٵi�1 6�\w���p�h� �b< ð(�K0��Vk�͆-�Ă�ú��$�&TvUQ�E����M:��K��˵z4c[��͡M����چl����`1P��Z%�P�����u4R��Ű1�$͖B�ǹ�m��(n�ǵ,�I96c�ҋt2�Qс+��5��Lf}�Qq[�P��D�N�OJ�:E�Ք����#����C3n�i�T�*�3���a�����НȎr����4SeYՀF:�k�<��\K���=ڶ	����4��-�s��Ql��H�Kn�!U��\�|~��B:p���c�䥳V����Ţ6m�{���r��A�ɡe�h0�H�f�͢�1�t�`��ֽw)�iPW�B��2�L�J֞�i�"i�5�r�E딒b�`�ܧjT�+҄7�V�'xF$����ӛq�A+YqHuV�/Us��J����ܳ ��9K)ƣ���Oi50���TS�v�*}D�l�'qPP�,Xb�w�������H ��H��W6��i�ۣh=�Y���Uy���4'r&�#�h�n�;�N����Br���OD-�̹�e�q�䬒�H�JÍkIRYr�-�Ru��Lo�qк�P�g6��ID��e���<���N�nG��dO(��d�n�K���hF6:Cq�y<f���ժ�������� ��N�n�q�N#�)˭7E��4ҳC,Be�ɠk�nk;E�\5�P�6�k;Y�h*1��sD�^�<�KofU�Ϟ�XI)�lwz�Q�:�Ә��ͽ�u�X�!f��3U櫗6��Hshլ�DIp��SB����v��Y�J�>��.�+ߵ$�-�[[H�ТL��QgeJd]�3%.-;��JnI��$��(��
18#Zc0ݐ��B�ӭ(�9��B�ʊ��ͽorSA1�m�Y��Vm�w�6�3f�.��5q�&�ƳJ;�e�ݨ^��@�����z��jjZj4&�X)q#�L݌I��M��z�]��V��a�"���t��q�ш�����n�8�D-���E�1aW�+,L�o[6��\�{u�7M%��� اx7a�0%[B�nV�dX�>Xf5
n��2cV��@Pre*�����CZ*�oڎ�Q�a!�X(�c�b��Y6ٙRT����'+r��\�y�Al��n�b�:�fML����#_Yd;��ܨs\:�2��7E�X�t��I�,`����Wb�$D��ܩc`(��Q��nءCwve�7�)ꚥK��Ks/.��]%J�fU�wW6,��X,�U��hjJ��S%Z������u�2>xf�ޜ���M4�;Q݆���������F�\iB'yD�b�h�Y% 	5�(�юE��F�HXB�T)�j&\�w,�21M�Z�յ�YC1T%{
��M� �yE�5��j��r^&Q�(ؽ�LIdL���Hf��K�R?n�g6����R����m����Que��ճ���/hL���f�݈d3�N`�t��k+s䖂�,�ͼ�Ke3hc���mK�Rw%�BK[���(l�S*^D��L=(��J��G���`�mM)e��ʼ��J�L����U@j&3�����H7`UխU�a���o^�LF�mV�rax�,�7(�E�MhsjZN��s۬/z���|�7���d�;�m2P�y�<�Z�ٗt�"vl f�ɴ�jd�Q�qS�d�����O �VTD�@�f�oq^؉aU�EG
��'BV~۳,�ڐ�fZ;R[B�Z�ҧ�m���S͔�
�k3g�S2C\U��4u�mB.7f�@y��'k���X�����k�m݅G@D�B����Jh�K7N��{O*�[��kݹ�͑�[1)��Jb�P`�m⨅C.��si��!-`�F
{{I� ���<tV����b�M�Xd�m[�N�L��6����Q��(ݳ!�c�ܬ��mFN\P��Y����W�u�Ar�2�bnnS5JN�\���� FvV�ݫ)
k"��g��z�ݝ������ZC��Ēn��M�!�Yx�!*��%k��A����&-JXJ;ܗ,B�8���t���b��Y��bx�7u��k�6ޛ��e渐��R�8�$�m̂�#�H�{���	��<Ya@�t�Vi���k6m�v��KwNT�o�ᅄ��MfUźq�^�2��IJx+eh���ք�w9Gf����*�zeh��L�K+l!O6������TԴ����K�XpA���eL��м�N���j�ݷd:
sE������m�EtQ��I@�ڵt���H�v���ol�
�nǈ6�"y-���+T%����Ȱ�.�l�N�n��(�&�m�	�¬�tV�k�%h�Y�@�	��n�ɲ�#!p%��^�����J�[*T*\m�tFV�o�Z9XmS��\��h6�Ӏ `�S�5���4���r�0&h��%���[zٱPx/6��l�<��X˻�E;[v���L��7n��Z��!����K7�A�ٔ.8�lkBd'/r�؍ɬ���L��[{���R�5�7�ɸ�2�F����v��Z�N���Ǵ��sH��ە.��w^�q�I�w7d��5�����m����Y�v�V�b�õ���e��+D�;v�҉�����($M��BFS	N�X�i�GZ��E���=Д%��e�i�:���j��6�wf�+:�-��X��v���ua�m7V�m'tN$��y!��Y�݇IT9�t��˓wB����Y[H�	sn붎��wm$ �;P��5��e֪z�\�@]f
����rn�Tl���R)5D��adpE��1"wbnzԮf�EP�nR|��=�gqi�[zf�E�����C��U-ƵFs4
��9�k.���"�%ފQ�f�-��ɬ���>��w6����Vl�����K�v-��5Щ�/�G
qI�+��H	��Z�C���B0ј���V3X��aIKH�f�66��;���:r�bn6�-|#�c�D��t��h�π�ah!���l�a��E�U�z7M�u+J˥o�з�ǵ,q��&���l+��b���F��3n������J�3F���Ż/>��Պ7�1`-=K���1=�kYx]=ZoJ�D�3>,*J�Թp��C�*���@�7��* 5Z��:w����6I::ʧ4jX��U�f���1�v@�R[#����ݚm��2��̽u{l�Ğ�9"�[�L��Igc�$J��y[�M�T�p,�؇Fn��a|D7��]26�ʹ�Gҕ�JgN0��d���&�ӭUe]]4&`0�g^�u6�SىK`ʘ�I�����R�,e
tkd�k`,�ͬ�J֕��j	6�ѷF�r"1͵HZT�K����MMÐE[[��V�fj(��7Y�Ѷ�ۦ,`��r۪X팀:Ut��`C���*ɑ��z:�t<�0L��ּӬ�%�١��Dai��kV��-�#�
En"������ Un��Z�lQ5�-��ׇ���Sg�=]ݝ��C7i������+`1�Z��Ht[�J�N���jS����-i�7�"�	6)�w6��t�5vu9{���&�i�Jg!�N#� �Rڼ@��Kr��7[q%N�n����R���/V����a�x���v��M�鳠�/@u!k2a�`�[��u�f�(	@3��F�{��%<Ͷ �e�m�	����F�w3�Y��.�aS��+to��1

������͔d�8��cU�6K�1���P۫�Z��[�[��~�q�¯6����oVM�4��i[ae̬a��q�t�ܫ���Y�a����!*S!�]u�en͊%����N+>�Bf��)�'�0-#V1�[t艴��������Ӡ�h�.ӫ�&�u0��u�yW��Ȭ4��h�Um�[�5i�iG@�!|�7qb�S���L��p@���[�����V����K
��Z��&�ͷmH�Q{��CE0k!7R5�!v�k�ˌS���l�l�b�v}��۶�
�XAd���f�f
�.F�,ac�퐭d�T;��ĝ��L��e*���nk��݈l����MX8��)h`�{��r��?:X6����q��^Q�W�Tw���p`j��&�j�SN-nݧ��Ǔn޽�q�����YN��ķ/R��-X7cwe��Z�����!�[�V=��:�R*�D�T*�k2�*�"�����
�ަh�z�J�]髶0bۨ0�{5�������N�A�ben�h�z�2*&���&Z�h�a�7�CEFw`�7H�x�8���Su�P�i-���}EN�Zr�YL9���^Y�RT��k��ﯮ����|[�W�Mu~��W�@i�%*�6��r���7n�T�&t��XSd�ਟ��n�e��L��V�m���JX����۹W,rvd��At;"�5b��e��y���$��9����l��;��ۑ��s�XSs)R�+��|n��	Q�!��Χ��DZ�Y����g}MZ]��L�<n�;��po�l��7Ob�e��-:Ee�[N��NYV�t�z�̓�Yܶ>�}9��f�u��.m�l:%!df��mA� ˝��D,[�����k�2k<�R��338wrP�n<�N���[�N39簨\-����L�K٩��y��g:[{�ɩh9iֻ2�\#��yW>��f�̭�Z�H�-`��k_<k%is+�Shg�*#�`�\Vѝu�����Ԩ�@�C�<��}��/o� �q09wZ�j���/X��!��b��N�p�&`�f>�|v�R�}�b=3rI�M���C�c� ��ѱ^���\�j����;�K�;�(�IWn��\�=;
߆�n�Sso�xC[���ũ��#wK޻}@m��v@��}�8�j����tGi`\
�>�r��,���F.���U���6��'���(E��J9���E�Ҏ۾�
=�[LJ��-�	��7Q�Y��G�z��^���C�4I�������R�¶]�<=����G�
#FE��5Q��2�*T�lH��6G�"��Q!��w�T�8��q���[�tcm݌Ê�.j�������ͤ(:@jQM7z�+�;s�)VY�G[�g�-n�ĕ�x��5�wWop��c+�r��%V�].��ۢL>���4f�#N�@���V@�����"�`_	��nF�s�����k���C,��N��:8-�;�w �N������Ck5���BX�%�3�֧��f6�v��)�c���ȳ���_K@�6hԼ�����"]9�]7��ݻX3�OY���X��&�)�k�d�]V&��#�g$��t��Ä�_]��H�r����-!f�$�O)"�^+K6����6�8C;���w��7!����B��"ӳI[l&��֮A�+��{
r�A����%=�w��\�0D�^Pnh���ron��ujҚ��g�w,���9ۼ\,$��70�������%2>�w�VP������_���f��8�gWI����QH�i���7Ov,7b����F���\�v�c��p�uˠ�f�aFE�z�,pL�ev%��
L�U��v�"s��af9!���Y�xv*�r�����ټ�h8dTD�n��������ފx�g^�=X�����K%v�����0tyM8+ODļ�]����u�Bibcs���2�!�er3~�lҀK5���R��{n�f��w�Ա�i�=�Λ�K�W]����O�\5�Ҏ��k���j�Yt�RM�d�� l�s2k����J�"YW[�Fr�)���c#m���Q��8���i��W]�&�Nͩ�a"��ҙ��C�
��tk �J�'q��$ϟv���Y-�H*T�c�X�a��-��Vn�}�t�f��Qi/,�|A1�Cr+����[G�r�Rܠ�ӑ@��}\q��N����@�xP�r�c152�Yï���&�ms9&-w0�Jz�>�L��4".�{Vq]l
�l�[6�ۧ�Zb�oU[�k���	Ǒ>tQ�n��࣑�M�
�)�u��O�e��N?�sf�vi���.[�2�s���z�<gj0b������o�3��Nqz*�ٲ�j�ָ�1z^4T�����6p�zn�e�e�����]�@�5օ�����k�dX�NGOY��;���+���c�Ҥ6�f�W�z��9ك
ǂj��.�C�}:��Gʛo0�6J.2��(��V�����xGHa5��R�b�6�xo#;Ή�Α�B���A�.��\��rЗB�����]7S�wN���tY���,]ïk��
�-ӡ5�mgWU� B��g�l��ڕ�R�o\⧻H�e�\�oms����z(z�׼�]���9����u�eXV@����`��$藹��wى�|�dtW��s����t�i2�:���dj�Gk��v�]�Z^R/�j紗\��gm�Ӊ��"�6{�%YYeZ˕���c׃�Ɓ{�&:V��+�5j��ժ�q�rD�9��/tZm�.�X}�:�1���X:5�����I�	L���ץ����b�m�DE4�\UΞf�.J�7�V˭���b`A]j�pp+��Z5��vo���rT�7��(J��(b9r���R�;�R�=pk���q��l;��w���Y�Q_fX�j^}�It�cP}������]+sL�@x��U�&Vԫ��9z�f��H[ݵ�G)e��\2��a��CeJ�m�+4A;�R��=r�|�9�
IS}�K�vwqX0�:���"�L��0����2�T`A��WU��Y<�q����s�+[[����-���[{͝)�;2�麼�Z��v�7O+v������F��F����i�����80`�m�(_�͌7��w��$(Xk"���莡ܰ3*��r����TN=ZX������!�/�6�o:)�X�k`
.`�������T�yNE�v�s��U�1'Q��E���J2���UŨ���6>Z_,+��� �أٓ~��/���-�\��r8B�"��Z]�hU"Om��*; vo�\��(��<"3g82�K�j_W�J9M�����Sw�ܣi����ǠhFVf�,��zw%؍�9�P��
Zz�1>�����UN:v�b�~]z���Uᘡ&{����H��~-����{���� �r�C*K�����-Tޭ��n�T�-����h�-��r���h1)t�;FBrT�����i�Y���`%Tz_M��2�X��o1���hG��s)%���~���<�`v�8�8��	��yڐjY����e!Ι�+�����-Z��C]w+��ur�ml��3�E�ɚ��R�(N�oM�
�;J���9h�Vm�Wobx�.�x�l�2�{2�g)"b�w53@�ud�e��[gX�E���4�s&\�;�g1l��c����U�ow��(����	��sy�ô����\���Y��񓫗��8\u�;���8q�إ2�Ҙ풕h�����C���ږ2��5s�l2��=.�NCZ��gϹ�zm�S��Ls�x(N����4�2��*�b"�]��ajQ�����xd���A���R6̮�0����VK&(p��nW㑶Xw�ۗա/�ԝ�Z�ҵ}e��X1����ц#�|���֘{�a���^ ��Hu�\:<��k{��\��͓nB4l�7�P���we�+%�n��s:�\���:�תs���j��H��m���D�ݺVn:� }��&�낻p�x�Q���i��a��lQ�X�����V���oxn���{I�M��fN4��&c��cf�}�c,�lK}Bv+ø�K<������І���[+bg�ݸ�7	���w��gP����l/�ӊ�o�8A[���e�7"C�[�ᝂ�v=��f�*b��v�Z��i1���"qN�
��U���&�+�qk���gGe�e�
�G�ӥ��uQ��(�jF:r��(��&l[>�	+��JL�n�W2f�����U^��{����tGT�S(��5H�Ϧ��¤(�.*���'wVX�����3E578�����'h�Ӓmstn���Y9����`
�8�O���dv��3/���>�;�4�����:4
���?uҵg;_�^f7Y�*�6�Za��Γ�5PΛX�l��[��M����MF��dȖ�tFI��٪1���h�u�H'w�����\��Z�od��!RQ��Ff@�1(��6)�(��'&�RfP��I$�I$�$�I$�I$�I$�I$�H��H�'�1ō&�R�-:N����*s�}�g!W#)V��gWe��T�Ty�u�*��(�h1#b�>�y:�l��)u��m��u�q�FE��P���q^�s���vb�xѝ�PCSu�^i7�	������O!�6s6�4�j��E]�͂������5O��'��s��\�z�^�����ZwF�vW	E��F����]��1F;!����V�Xx���N����
�A�����S�[� �t�qe�,����a�A��l���î�ᵜ��7w�QT�4i"��GJ��u{Bst�i�O��7S��*�p�e0e4�nK֫P6�:��lN���db��]X�+e�O0k�䆋=�������&M[u�6RG(�A1b�M�Po�޸����J͹��m(5�ݹg�m:�)���<�5��{������T��L�{eA�[=�����ho��K�_X��;�������ԗ9k7c+�?����w��p�w����������Ē$���t�:��f�Z��Er��C���?�`��c��$QԐ��O�`w�բ�!��Pw=���h���݊2����+mP��R�)o�n��@p*x����eZ2�U�l7�{(������{.z�k��@��T��e����[+܉
N5%��^$3&i�M}*!���$�I�����s]*gMV��=m��L��GWepL�����|��֯�H*Γd�(&�Z�[��P7Ux�i-#+�J� jA2�V0��ʊ��$]p��gӴ�L��ɪ���Ww���6.�Qhⶹ�CwF�n�O�T	y�٨彼W�,S8��!u�TmWKaE�)��iS��#�R�[��H`�ҋX-��������u1:e�/��(í�Ǽ1G��T����37:1�Q}��T����r�@��`=y�T4�]t��cťc��.�i����TKe�	d�qb�(�ufRS�gx��ݩ*��]�s83i�kj��!.�P�F���ܶqƚ �����N��Qj�Ϥ��pS�N�Kh�r�#�*5AZ8��	��qdU����̻drțY2$�~:k#��m2��"�ywD�U��^��4�AT�KG;�^>z��Ux@���ܝ:��&��ה�,��j

���>%�a�+�m�{�E]FJ7���ml�PR�*e:��(:H�	AĢ�i.�l�7K,�0�����vؔZT��$s��Z�%���M@�\f��K&�{�S5i�����e[t��XHlu��E]b-7)e�]%�QT�A���#��ᙪ�5�O%��ϧd��m' �)�L���?&��-�t����v��vc���Jn`�ԕxV7��LT�����s+$p:�Y*T*�RWh��P��FWƣ��K�Nᶶ�X�����L:�;��ы���ud�w�}zU9R2��@r�3�1\�� o_%V�(|��[�Ɛ�q#rW3�X�e�;�����ՋU���,&1���vR��GNC#ԁqڳf�k����"�՛����e �c���kI�4���m�w�/Ԟ ��_t8�:#V�;�2f�Y�W�c#KR�X�-qNv�uaŞղk����c[�[P�_bۭmQ��k��*��;w0^C�ګ���S:�k�	S���U�G���y)�X���V� N�ૢ�FCh�eHC�]r���r���XA^��P�*�Ӵ��72	6�#$l�H/�Qԃ�E���w�Wa[�񵱢�7R�3�(^}���v�rb�Uǲ����:[{ʗ,���%d��r�ԉW)|�C�]�&�*�Yf̨R4�Z��َ
VMJ�^@мJ`�Bh�ʔ�I%�L�:�8c.�+���z^rS��:*���-EY������_ϴ"MD�/#��3��ltug�T� G�����A��&�.�#ؐ�CE#nnc�+v�Jj���Gy�MoMԐ 1Th`���Wҥ��܁��۹� w;\�swtӒ.2��Pvٰ�����.��yۛeƙy Ǻ�Mj�G���0q ����ۮ]KiGP��v�#.����s�8S��)�`�+x� 
��݂��iw醆���O�g س��7 ���X_n�D5�1N����U�ӾhSy��kbEj��n>��X�QK�A-�'�h�m�^�U�d�3B�F�f?�v*�5���WW���1
є ▪:̵F��D�16��5n�8CȪ��=J�z�m*���ԩ��[s,L/R�j;n��?L�d�wkc�N��.͢��'窱ʱt�
Ok�\�HA��,j�AXmQ{�A\���/O2ނ><N�����?L#f��ҩ�|d7L3��5�k2�Nd)y��{m^^�A�4���Ԋ���]&���u{V����I��T(� I�{�*�=!d��'h�o���}C���mk�@�s�\�Y/�J�l�Vd����	I�V0���e�*ȼ��N��De�A�Y��\�*��)������)�-5+,:���2�y�ՅMUGJb6���-`�9!`b��8��%;Z��X���ẵ������v���E\a�]S���gU�U]�8�-д�m�M�.�t��e�j��65��N�:��X�2a`mVB[��1�X�[p: /�EŅѴ����Lw���C�.��284�)ۚo�蝆��L��m�%��� �1 L�c��4�,�KIK�e+��M����
m�J�Й9�FƋF�%�*;�6�N�+���(\Z6u�(��q��Ĩ���T�y�Ө�Q4J&����;��v�e�Ӯ���PН�Ƿ:��+n����H�is���m Lb�J�#[�4kn����wd[j��ŁW����,��Oaf��J���*;X�v�uU�KL��W���i
ǽ{��l@�@�֜����c��N��(K�(&&.�����iE�-�m�]�s3sŲA�9���Ղ��iU�DVr�[��;�AaPf��J5����@|l���F[��U�W��n��%����st�M�W�ʳ���&.�$&���+���� R�k@V����&8���QJ|���y��k�0`�:���3@�X��e^]%��t��������J�\=��F��6>Qm����о!غ}9Ӥ$�84�c4�g����gZm͸����w*��������X�E|�aKO�9L>���n�N[���;f�׮��zk��|5iҐ��h��Ũ�Ū��*i@�&;���X��b�0�Ҩ¯��qYC���c�-�*{ls
 <�&0�
�"�ts�,+t�9���<�Ӵ�Q�	Tzk�vM cLq(��d�77V��:���5��w�ː�-�\�iʓ\`���m�+o>CP�m����R;y��|���(�z��W��(��mm����ۥ�y����ͬC`�J8�c�P�h>5TR��̓��.Dp �o��%J$m
��-�W�֬m�X�"��m���j� n0:���������"F����s�DZ�WM�Wp�.\*vE(���t�ҩh+^-j�h�2�8f8*�\,�8`���e��� ~�`Yь�vIH�F�9��d�X/��7���M�Sn�%1=�cWз|#h��uʪ탕�Kz�ص�����V�	:XM�l-���m�8�WE*Gi̡b��rf�%�#x�*k��*�t�҅-K���Q����
�%l�p�z�Z�������=�FZW���5���OqIm��)(%HO�>Z�X��^8p����]/���t�EV;R����*�3�e 0��G�΢|��J����t�Z���wY\������5��F����y��i:[�4 "��ᒱû����X���ބƘ�8��-}�)���*p�p*�����h�Ls�G��2m^�� �J-�=j�wD�N7��͊f�[F��Caщo%M�Tޕy�D�ɳ]VPm���*�IȚ�m!�)�vD/=z�uŗxFr�ǖ��D���{���tU,�oL�p�u�(Y�z �m*�O�n�5b�n	}˱@�DeA�1����*�0����(B@�]�k�s��eB*�}B�F��t�f@�4j����7x�ͷ@՜�:��b�@�u�9>�IP�5�25�k	U�9|n�O�M�e�o�xf���A:z�t��r��h�8\4P���s��lNi��V<�,�*k��IDVLo3ڀIg9�orc��5��ѣf�e�z� SP���{Y>#��8l����N��2�8I��Xk���V�آ�z)Ҭ��,6��v� řj���*?i�fVvS�Q'N�ǔZ���VJ�u{ih��h&�4�/�u��n���oj��
��/���H���j4,�j<G;J=�j$�5ʨ��I| �N]�[�2�'���G�h�A0�Y�P��o%A�i2ѡF���JQ��ܴ�\�Su;R0q_*4e�=���*@R1]�f̗Ǵ�6�r���JL��?��R�x�]�+6�ى�PWqUrd�P�Ah6� ���Z1B(4������H�khMt�RhKJ�,.
;ىQͬlK�ۨ�Kkq���q�כ�h96���]����"�D�����s,�$`v69��A�.�r�w�M�̷}�%�aȺ\�d���e�*.nؕ&�tЮ��g��7���e@�
,.�D˝l�Ub�ڵy�^�@,͋j��"�k�Ξ;���o26UZ��>�s��ٝ̚wuDٙ*�6���陔s*Rj��F�#�-�5�"˗��(q�;{M���7��"l�pa0��ku�M������޿�T"���C`�B$�����$(�,���$��u��Qv�r:�aGp��46ڟ,�b�9x�f�8�㷂�� IW�;�U�N���%m�h�h;lU��f���l���!��EP���[7�AyZLscVH+NB�>��m�����2 oo*ww6zU�W���Q�[�c׏���a6���ט����t�미k��P�)�t5�AX��-��8<4��WqQ�R������)�v1���Ņ����5�w����}@�|W	�Fglb ��=���@��o�uZ<�t�cw��ɫ/.���E[�Q�N���5���Ψ�7��e��'F�'ڄ��M�E�K�}��vR�Z�����Va��1ym.r>n���6\��u�ĳ�qK+P�.b��Pێ��c�x����K�ҝ�!�[턶���mq���f�J	;�; Q�궃��ۤb�!ӻ��i��fK՝Hme�G9_�; �$���P�&T4��@P R�������N�2�(���i�ih(ii �rR���)hN,���
p�	C��NA�8 �ER��!�w�IT�Х47���!��)R�܎j��� �W&������)CB6��p��
A���J �N�������h�ϯ3�:���f�#�Y�cf��S�GjYS��Wӹ��bJ4�j�I�}@tg����W�T&�m�/n�X��E���١�})�|�	d7`\����8
]�V�G��k ��xﻤ0�<"p�SPmՙOx���1������\���Fѳ	@���匜��Ҩܑ�:9]�Ee��<3"+a�7q=���L�z ����%�]�f�Z��K��Y,4�g�PUA�A*�	�{�]�]`X��q0�m���z�3��*�}���Du�n��6�ߩd����N����˹$&r�]N��#dvj�)�8[;�5��QQ�zsRL�����VR�t��ٽC𽉧���7(A8g�.�=p;���R�s�z�U�3��q�������jB�mm�vz�N"O�����$o��q�eI�Ӕ�V9����/+$f��1l0��}�� �̾X4�����H,��HܽW�Ĵ�_��k &��������]�CM��iO/���v�r���=�j���B�,�a�cx�M��h�6����1'_&R�J�P�}���Z���gz��O�Q��,Lg��=e�����T����(�qI�e��Bq�x�d^��=����[�p����P�A��25�J35T\��$�x4�Vˍ4bq��*c�&�t�P[��0���g�(����]J��:3�5�K��!iu�Cv���ZR4׭X����&L��ͣd���q"�X��������t�v$�;D��rQ8�r>�-977��]���0��V�Ǒ�~T6�fӭI��V�@1FՌ]J��̊u�Aj7�T���𨽵��4���3b@�*S��.c]���}O4T�������Ɯ�ʆ��T�9�����c*��B|��Ow�˳��k�GhTp-�|_#8g%'!�H��D?GdU���d��.i���d*w�F��[H�\���S�	�t�k����--��wj�S�q�.;�yY�|����^��H�R��s�i\qdd��3\�H_7���%�K�ŵ;��[f�9H��M@>4��V��7�� C{�m���z��umXe�qa����=P������Td9S%;R���#m̖J�������eƜ4̓���&9ڙ�'�:�z�M\�O�s�^��'->Rt
����T���b
|8gf��싍N�tM�H"ebޱ8�cE��y�����5݉�h�P�ױ�V��T���q����43�<Q�Τ�g-Q�p����%^T��n��Ozr�pU7؀-����v���U�9m[C�5��}�x� Gs�`� �������	���k���˳�J�2��;�V���Ɩ+�zOk �uɾ�)��F۰���C����=�ݴ���ti,=����7�	մ�;y��AW�5���5���f�},�G�5�2�6	�Voڦ��<j9\�F��jocp8��<�s���8q�d���9I�,��F�m�^'�/y�Y�c�x��%r&��\J*�Ř���F>�r���]��[��Pٍ��;�D�h7j�ŵZ�<��|��\�b5d�S��1���&Y����
�������m=��p�6�2l��F9�J��o�ѱJ�`V�R��w��w�Bk&0e;}~�5nwK���4m�%���}�(�!���u�/F�yH����ӄ&�Qp]�G.�#�����w�g�|+��K�iC��8���N�	i�R�nڶ]��̂<���ς���yRp�`ä����~,>&��H��;U�8�0�(��=�]�
�Y	�b��;u-������Uh�ۻx�b#�MF'��(ܲRFH�,>r��d��pcw�B3`�"�8���J2MoK�3��8@��:�zz��-�	�Њ�#I�\��j���܆��� vF�It#7��n�3�EFq��I_r�b�X��9��.օ����U��l�3�����
m���gr��Z1�t�{�� ,����d���;� _*q�֚��{K� M{ad�΀���]�"�a���//��u��G)�7�q��$v�K`x�5RR����mߟYQܣ�G
 �j }�M��tě�}��(�%`YQ82�T3옺:�l�K�wP�Y���m���ӽx��5��㭺BfihZ�+�;�y[%+�74Iï{��}(I�e,M���R�G��p���(�֌��g-�,
#N�}��cLb=�7d�M/ ��9ǝ�{��OA��ځQe��U��iP�1��F�EC���6��y�8�rLdn����}I�=��{t������[�#�����{*}T��1
-s-�M��� a���D���*�w\���w�Y��aUOG-�j��0������\�[��/+�jy"ʍ+�-V���y�N��֡�������k�^�$��Oo�i��˹^BLU2�n����y����Y���3�ue_r�z�SȄ�d�KZ#�זm=Գ�܀��-��5����z:�-	6'� J�˯q��n�c�e��r̺Y�L�/MG�8�+�����<*�0d�!I�UK8��f�轨��s�m���1I�����o*���F8�q�g�(EBMi6�/�BM��&����4����=��^�m{���qk\�9o�V���_�n�,���<�j����>\[��/0���.�VR��z
��	6���Ӝ�ا�i���4p���t�u�t޵�6Ҿ^�/��^S�2������Ʀ�sΏx&sk��9��CU�n!2�WD��E(�c�}��G��y/k��H��1��7�lTd%�B~0*Q�ۭc`m�f�f	���������:Q��M"��*e6�X���;�<>+=^���Aʂ��"Q��l*�W&�R"��k�]�}�K��C������7�U������g8��M"q�I���,��(�������4��T���gz�M���M�.5�<&ʼ����,�TN��v+/���Ka-�6���'dN\��� �;�_Ѧ3�oG$�D�O{�e_=D�zr���mlZ��~��<���G7'a,w��dݐI.zk�A.���YJ�D�J���sE_ov�ޙ]��i�o݈�^�� �j/yS湭UF���{�^	��,N5ɞW�pa7�3U���l�/�0��G7�W@l
��-��}��A5�u-�;΋1�QHF��B�D�|�v��ӰP^4I�F�{�@:AB�(jhL��*��Pcd4u���1�wY,͋$�̵�I���jrEjGI%\֠�P�f�T;Ӝ���Hrr;��fe� An�6C��t�۬4˸�u�7��b���e{"��&3GC��۾u�n�uD��3,D�L�jP!-0a݋SP�4�-���7�:��;�<s���J�&v�f�k�zp�kId��^��]�U���y�n�i�{����c,i����MEѸz��W�c�%x����ݻ��PR{�dg��*�u�K�c�����y<����������4�<G������E��Ÿ���5Ul�%�8�����"3ӝ0��>���#銟G�'��{9yr����y�\��oW".��헼�Ł5�w)5�.���cbW�^=�.c�}н�K:k
���Ͳ�NM��n݄�8�b��A{Yjp��<�,�F�'i+�i
�n���WJ^ѧ"�q�H �pJD���<'u�ҷ@!��k�=R�pV;n���#��-ʾ5��n�V&����q�m�f��-G����.�oW��@��K�wR�Ӵj;����ֈ���I������JT�uQ�K��`�gpW�����S�gl��ʑgM�{}��G����2���Q�\0�GF) �f&�7.�X��3x�}-:�ހ��/���ܺ�.M���XCMCz]l��[C�*kw���Hv8�u&�GS�}��l�[�:���.R\f|���z��Y�������S��(�v�Vq\��G�]��-1��M��l+f�E�7Szi���	����o�5�*�84&�ic�^�-�5�F�g
��1����J0iF���v�w��~P��q�Ĺ�k����Jr�̊����7]`l�C*��f�����D�B�AK�j��y�B9:1�n��c9�+W"����5[�2�Gy�k�Ch�Z�l%c6��[i�[k�C�DM;�w�U,h�(��t\������n��«~gu�����hͪ��BN�t�K����*WV�+��q+��nҙ�o1b�j�wS����l�������73��IH<�]������.;gr�{�%RЍf�,�ʣM�ȷs�I@����h���]����YQP�ΙڗK^˜��vκM3�1N_U6�����Imtr��<��9�V�'=;��c8u�o�� n�e�+���#%�����ʁ����3\r�s�M��?bZ��r�������Η-�2F������NlD\I�WP�&�spg�N1��(�����O%#�HW���_WF�����"���0r)rrQ)��(�ZJZ��ƚ(iiB�(�hi�I�Q�\��F�P&�hC"��B���2L��]IICB�!��d�HSLCLEd5��#����A��v��QJ�T%
�@�E+��o�[��L�̿�%�-�5�OǠ��CŹ*P?�1C:)}0��'"���ԯ9�[��a~AlK�eD�����
�qƘK0L�\�z��y������V��Z;>��rml�o8Q?B���?���%���c�9ը ���X���}��(�%�
�<x+��g���L�[/��o����k�kݛ"ro�<�pЁ�.��>�Ƹ�[N��Fݰ+gI=��Q�{���Q�.D���#�W�3����֧4��9��Ʉ �u^$�(�˗M���tO��܃'��~�@�<*z4��ؗ��u���>��k"Of+n����{\T�\~R��{^��ȪQ2���+�7q�pۅ�aZL귥���
2v~9s�F�s���;tor�K$�z����0kەu�h�n9J�dJH��$G;�y���e:͍{����9�={sru��[�%�Mu�s4�]}��ځ���O�rVkXo���/"��Du�1���qȀgFe����	5��Ј�ٝ�>oA<J�r�r/�FD_+��m��Q�OF�oE�fN�m���\��,Ut��I��n1�/���7�Xo��.�=�z8)�\�$��ۣ��n]XK�Y�?�b�Pǡɔ+5w���9��^sN烊b�;�	T��JϤ�IE�;h_ih��Mk�kF���+n�邂�x�-�ё+א_�5�� ����.��=�8'�i��]cF��,,�Hj�
];zyy��A�>���A�u�V��=bv�)��]�۴�U$�u��9��+�uj)5��������&�%`��PDh�"�/�j8�,r��U��#V���hم��ֱ�nD�%߷$?H��Q�s��ven�6Rvlp-*�&E��f>0��2��(���V��m��{tx�iM"1�Fxڋ
�
�&U�ͿJw��Թ1���Zj�8$��k*8�KN�=���3�X�R�G�t�y;�cM��wς[��� l�ܢc���Бh��Pa�w�a�����]����R*��R1>iŔӦ�.��(1|#	�G�ҽ�����^��^q�}���#�y���y/�� w���M�'Q�P��ԅy+�G��N���B��S�g���s��Z��qth��X�yP�L�:JXwq?K���e:v��5'G��0�F;+�*W�˽ㅧ.�¡��aڑ�Nx�Y�g-L�DL���] daE�$�
i9+��ԛ��w�xwu}C�܏|璿K�p}��w��r��S�(N���F�{���	��O��?Á���N�Oa���_%�����qs#�oa�����{9��@�ƴ��=G�d�RP��]��^���=��?{�G��'S�x	�nO���S���_%�N�=��#���X���>Ƥz}s3�D)�:�ޅ1����M�����;��$>�;����_c�1:��M���C�ܙ!�s�����nf� ��x��|��w���߇�į�u�*|}�Ò�;�y��F��9���������9s)��+��`��m�5��y�������>�|��5)����K�brh�t���9 q�r�/���'Q����NNp<�/�7� Q�ƭ�hEܦ�š�D9��f*}�S菼k�A짓�� �]}��|�y�=�֖��q��{����䇱��.a볬�z����|�ϸ�cR��J��Ȕn=��C�N�(>���_� M�旻�_y�KK䆳�1힟��#ᚫ{�	�GO�B�F�C�;<�8����>��|���>�<�����eי�.@k��9{+���ɑ�~��~��_-�$>�Ney��`���xs;���2S�p���;>�N']a܅���>H��������.d����6�t���Z��ǯ=t��4i����ޣ�j��v�-9S����˛�#�{E?tv�d�7[�DWQ�} �P��S��=��V�F�������i�����}q�7(�{�C��sO/X'�;�%<���y��On:� �L���C�G�lu�G+{�����'������Dt���}��C|���Ԯ��y��)�W���T�5փ�O%���B� z��5��������u��}���܏�w/��/���}7w�z�ߘ�kx��� w����]���!���y�q߽}��>é
>:���|��N��|�����n���_%{�����r�7�#��E�T��f!�P���t�a��C���_u�ą!�?C�<b��ܛ�o����=]��ϚC�z������G�OLť9���ιߟw�[������(�P�>u��_���C�p<��~���Oe�M�a�/��C�܉u��}��W�Ͻ�>����c'7�џ
q<A���B�!�/0�K���{)�`y/r��	��yuw캐��9�Yg=�zwk:ߝ{�����z�e��P�qބ����;���;�>��оN���e)O���	�f���ۿ9��|�^�H��=Πz�w��Ox����'xy&HR��z��b>K�l<���[������ϗ�o�|o���~���܆���O�`��{#�X��=���y��5��縅�� u�/��/�Í�>K�����Fn�~}�+��\%�:�`T��40*��T�?e4|��r�}WEQP��UY0�9�����ߕ�sC� �d������4UԖڝ:S�������"�sֹ�޽����?�s]�s Q��K��	ܔJw=@���/P��i
�iy���-�Y�I�/��X���	����Q0N�ǋ�_���N��er2My���c�'��<Ġ�]��>C���	���Z�߾y�<����^.e����X/p�s��S�xH�'��Jpq�����\�c���7'��h��:���ǢP�/�X�.���/�x;š��Cf`}!�<��&�S5�1��)��tq�x��7��<�j����}�]w��R���;���C�|�}���Իy�K��ǒ���C��c���]����ؼ�짜o��������7d.���=��:��_o��C�|�Ͼм�l��V�~�a{��1�_t�LgW���Dr;L��Ϻbǣ&">=�� y����MB�`=����~����x���C�i���N'r��:��=�}ߞ�ϒ<�n��{l��>��|`=C�}�������b���{]{�}�Ǆ����G�GrJ���x���2G��$>3a{��������B�Ѽ��g�R����_d��e�|��>���xθ��s���מ��"dw���`u9+�'�u!G���ޱuՒw!Hp}�{/װs)�I���x�|���A�9��U���� W�K>���g2��w
Mܣ����;\����k�'�\��>�|-㾧swH��:�B:��!.5�&�w:�D�Wi +���/9��׾��������z �]��Q�w�Mw��d'P�1 �Ca��P�ː	��{	A�P�{���vk7�ǜ�ߞ��D9��˨^�ԇ�>_{��;�~by q��p<u��d�rw!��p�@�η�ֳ�:�z���;�W�f�<^A��}']�W�&K�}#�Ѽ Ժ��_`ߞ�O`vy�HR���Ho����&w&ݞ��?G�����z:���=��N������u��j��d6u���Gz�{��r%��)��u�u�z���\q��{�qHR�#ܼZ����/Q̞B�GC�P;�`�����Dd��1(=���G��9����|�w�z":c�ސ�~�����`:��q����\��'8��:�<���4��{+�d���y��<�8�q�|�����PjG�JOe��J���
{�-/W��;��Jw!�xq���!�茘�b=Ѵ��3�}7:����͵����x{)�'�HRs�	I��� )s���縯�/�4��R{!�;��w���c���޽;��|��{�޽C�ԧǘ/w&�0}�4������p�!I��_e�~k�]K�<��/��0hx���� �;����q�s���^�ߢd����n����yq��I����|��:���v`@w��Ч\����/ѭ��w�)fwdo����3�uܾ���j���԰�]�٭��,uś�Ӈ϶��&A�ߔ�i�c�~eb��F����d�.oVgV�րSTl���<�'�y+�*� ��{ޏG��N��c���DL��r?!�	䎍�jS�v��sқ��N������>@�>ë�3�9ss�=�����+�n\��ZQߨ�!�_h{� o�S��fc�F��=�Ѿ�J{�8��h��Od�X!Ԛz��}�����n��Z���k�z��0�6Ԛ���*�2�Z�t��y���w!@A���=���'�����(�!�׆n���q�������>��}`L?������:ylՊ��}�D�ħ��ă�:U��q�B��#�K���W�G7^y�|��r���Չe��K�i��bnT8�7ߌ�*נ���7���@;��D�nN�s��
U��.�����I;��Cm�2̍���Nޗ|��nb�VL�L���1�to,P�x�yդ�]�5.�/��������Z�Of��Z��]��� š��k6��?���W��>F��}ȁ�r�&��s�@�S<z���M׶��qh<���8�Q���舵���� ~�1�Q�ĥq������(P��hM%�������Q�\߃Rs�嬌BQ����~�1��`߳�T�E�EM��bi�y$D�E�+��p|B�ݙ�R�l�p'oޤ�>�Du��L,`y��,�n����[���|S:�����7�F͹�G<�QJ"DVa!��4� ZO�c*/.�+�h-#����5a�84��lc��#]���B�~s7��� =�|�����W86�w
�w̖�[��t]W]4Sc����m�˴oU�{~�M�-�iu��K(5NYe��>b�UQ��Ř���/N��7-jLZ!��Ȩ��ɗ��X�!��Cy�l�U���
�5*ۗ�CiƯ�W%Ȝ!���"#��Ym8��P��o������'g��g���9�uhk�Ƚ�}���!΂<��k%�n���;���/�	���T��P��'�ӛ��5({̄��4��;]�RtR����Gv�`�mU%��V\=Wg��؛M�N�:��J��te%q��5�1���T ����sS%�8�)�m���q�8�jU�'#oCev�8�u
$'g\��b�Yn�GLY�������Z�E@�-l�L�����z���S2|dcGKoj���D�������������'ez�+�{�}����0��R��9��+LWKxo-DþN��T�)��:.�d�^��J��{{Dk���Ƶ�O�ٝC�f��.�7S���Y�
���+�Z6Y���J5|��@WW{SN��N�˦U-�M�Ty�7ڏ�mN�2떩�6�K5
�\l8�η�-�YՖYť�ֵ=��
��(��k=�e��w�0-d���,��)��n�ӫ�Lb4�އI���Lp,�s<{�V�ܳ �������v�A`'�,n�L�o&6�Rp�&]x)�N�q�b���j=;�_D/(�\��ګ�X��t��d`g
.��Ļ	���<�
YXپR�B����ꇮ�.��>V�n,�_K�yr9F#�A{�Z�΍;�?���f���s�hl@��Ԛ���VT��<pL-讃��އ�US@���39���4
��ښ�	:Y�l�[԰e&oCY�'��G�:�t@!�v��d�D�='Y�A��%9 ڂ�*l��"�cL��Q\���Q�q������<Te}����fR��};?Y�y鼏M�*��W��Lp��Z�A;3�$�d�;z��Xu{V�f��P��b������
^��J���,�bfYr+��������нÄKƑ�eIY�� ���je��䇲co�ķ4Nz)��dę�r�눰E�U4�X�Ёb����.��iH.�8����7KZ_v�c&VH C�Dཙ,�5����:�=��Ͷ�̄��u��	�>��KS7+(��M��O��%)7/OLCeoMA�*�[+�V1�%�`�r�qCu�Z�Uw��v:�q���ڸ�d���*�O�>��$Ƭ�D�RR�������v�VgK��7����إ�;cP7�̂`)�yt;�	W7WJ�}
�P�0�{�F�\���'����H����])W��:�����q���7!��<��Ն�םty�w���׾`Q��+E�MR�5I1L@PeWZ4Uj�(�$�?��`���R���h(7�NkN��#�&�)�',p�"b����

�2Ɗ0��,
()����y���,(1���s2����0����2rJ
����̒���s2*�3"&���0�
��)�¨"0����0��"2&��2��f�`�2C1��
bh�rL��#
�0,��«3�*�h���2�7�&�ّ30A���fHeM�e�.fQ��g]���Xk���?J��3��W�2���q�:�jI��Z0Fm�('T���il�7�K����'���%�K����TF��� ��m�Qw�����u��pоW�����,kB/u7����Q��b`�Eي�W��M�P��Ba^N�H$�7`&�u�Ö� p*zo6�@��W�_�-���琛�}n�9�=�<�]�(�Cy��ȘOь�7$�uScB���"`���3�¾�χ;��]T��p}7��C�qU��J�����9=�-_u�P7q9��!>�-��Fl��N�i=�s���>�0��<WM�m7Q�!Ĉ��U���ܽ:��47��¡y�� i�]u1�v_ 2�2�wI�	��\�k���W�A�Z1�=�6e�7�2P:&��މ��/�5
*��,Vk��)A�G��Dy�v��*�Q��rM�q�Wf�=�-�c	:��e&Ɇ��
�0�X!-0*%ڧ;�W"�'�����c��*Q�T���F/@��Fܮ��Ky"�KF�ot��nq��8q+��;X[�@տs�����\=w�.f���$�MUycs��pS/Zy�a��pE�ݧk7��9�6���&�x�g.��MR��F{2��S.�,C��Z��OS�MlOO.�I.��j6L�Z�������֬\LmD���躜��U�bD5�?
�xo�f�z��ګ(����_B{�f�ո��+I�T1T�����{|��=i�^�5��yC|�[Ci�e�R�u��S���s�l��y��h3�4�7a���y�����{���UZU���{��{�746���?Lp��7҈����m:���D2����Ǽr �7��<�Q�8�&̺sΏ��%N��B�ϓ]��,Vv�]�j�Z�,�c �hء`�cD�w�՗���	��e�q�5�oYP�g�7)_G+�9vvoѥI��L֧6�9����%���@c\N����/b^[�#ܪ!ڋ	�D�f��O0
��R��Z������p����*�=M�z���Q�h��W:�Eѷ�g��^ʄx�I�$�ȴ�=�?CnVX�;f�[V{]H��tY M5��VYD�ӳ�B{�:�݂�*��X��/�����յ��V��� ȡV���!I>WY�AL��ǉ�x�R��{��D������3���`����pc/*��%H,ܚ:���1����z2��M�� �K�p�^땻�f��pm�@<3K� ��6����1�*�ې����)��ǰ"�d�
�鳁���oq~ۮ3Ѿ��UR�!�rs��d6'-��y�Qi��GB�F�%/ZK*6��u<%4́f�$
�f���5F���V%��zO=�ꔮ#�X*QQ��^j ��uz����<�.ޘ��:wX*n��t7�N�L�������E��-����|�����.reS�E14Tv4��!H����B6�|��w�36�m���޾�m:d&:{�ɈR&�!X�qf�a��3Ǳ��>۝QЕ���`ڋ�TX�`N��j1�+$�8�����Ie���]��"�lգo.�q��x��;�Q|���\84"@�_tI�kY�D�
�F=a����
yNN,��d����	K�M���J�8$|����$���_S�3u�^�Z�s�(2yN{R�|OT�lMU2�IB~ݻ�������I�s�F�w[ˊJ,'	�S�rZyj�e��M�hM�QW^��	-,�9�A3*9u�3="7�4�
3z��Q+�������A����
RY�v����\m,�ǡ�1��}E/^/r�������O3�cQ7sH����{�*�;P�����K���x����WhrMj���]G��۱��a�i��w,uJD2)���q./��z7���fq��9#:J��.�$R��s\�|d6��(d9grz�"��	�M�IxJ*�ñ�+|UT>���Wc��S�S��'9�	lt��{�FzO�u�5s<��on����#U�re���!x�\I7���]�@ݶ3'f-
5����O�:�j* �PH��ir�Ue	nK+x�]�k�:PU�2��TK�[,�H���9���u_�W���N̪�����q��Q�{7��t��+4�P�v�v/x����X���+7��J��1��A0��W����>v9;I�ӸC�mV��w!��<�[o}�0��3���'2p^nț���J�����9VNaRr}6M�]�vV�	}EE�m�����%#�QVP<BK��G�6�e�_Gk#�=#����q%_��m�n�5��n�0.D�U�4x���j�zyv�-���k`��xs�l�</��a��ҵw+ڙ���Ǜ\�����:h7ƳM=o�;�L'�'#2�]��q��)�T�+�j�p���+g��� ��&v���7�{�ѱHJ��Lޒ[��T�I �f�P�j��z��ڀD����I���t�t9X�}�}�j��/u3aoQ	gpzM�=Y��Hi�^.L4g$��/�p�v{ջۏ�ݪ����u�IW�Oi�)��/ڋ���� Ǽ^�>q�u^�Q}f�v��yÚНm��]J�)�x6
�8��hf.ތ�LC�W�Vc�� ,�7X��vE{��Ln��2HR�Ҭ�}��DD�M7��D����ykx�'J%wp��p\v��;C��kpLo��������9��cEC��k�N�OR1��u�q�8��u�{v���x�o&�U�����}]�g[�kp�U�ŕ�����K\�i<q�����!�6Ɔ��=�����|�5��#��fm�x)	O��t����-��`������3��$�K	{rN�=$C)�H�RVP�u�ץ�h`ыr�N�ډ��9%��5�f �+�/@%a� ?[o�}��U8�
��S��ڭ
�T^�����ܮ�oOA�a�a��Cnt`/4��p�^�Z3����e���J�M��-�ޜ��Y![J�.6� �_G��{�g[�[���\�z.�ZP3 ���ң�Mae�|�͙����uzZ�@�J�����{a�;_�w�ۋb��9��z�f���y�"�Q[Ƌ�\�(��՚��x��={ˆg%e�يf�Ed
E��Ͳ�1G*7�c�&��pP!l I��F:��F���N�I	�pYTQ�p1��c6�:�rX�H��H�ƃ��֘�:[����댅�s�����iWK��(MB�nrc�?Ca,/��*�{�}Z��`��tyP\�p�����/�TC};	�W�3��W���.�:N޹St<Z0���W�h֑r>/��NR��m ���O&��LT2�b���ۊ�
��# �첑 *������G�[��M��W�+~K}p��ϦeT&#1La���m	AnJ�34�۾�����v���Z��pT`U
�$�Z�����,.I��g5ە1W9x`�Z�[�FP����u=�ܚ�{'���/�_�,D�8�>
�_>�ʥ��T�ҁ��E9���|��_zo@ŏQ����Q�#G�g��;��t�|��Mn�)�OZiA�.:�f[�3&S����ӿi�V
5�S�b�K*N�-F?*v+�U.�g���7�<\8;1=Z�EC���%�9M�.�0�R���Β����<0l>s����.>��p�n���b���>�r"L�č��TBj"�Ćk�);��u�J�����P
�|����\�@p\@�J53���G��\�:(���`SxB콘��' C�WƄb������s�)<��x#����,lts�]ڶHz�l�h�N�jEK�n&��J���C˥�I�d�wb
���!b�F:�6�#E�Z5�qZ��s+8:l��`0�)�8��:,�E�����.��Ȏ!�X�X'k�>�`s����;�w��e��"6��{h���D�y���U/T�-���ka�B
�z�|�k_gD�����v�K�
�?CQ������JT/y���[F�[l�>Rwtj�&Ź�^��WR�|�7�рkHB#ld���5��m &�4�8{�Bh�Ѧ-3}���<�dy��\V���8*��6&�&=;c�ζ�h�8s�r�J"��
�Lm�{sX)������(T�ν�Lt��Y�m�{�3�s6�L\{#��1'|�B��-�z��7�����y^1��ފ�ۡ��EA�y�Y��;�K
�lW6Qu�͡���<�-�^w���(q�3��Q�/����;�k��W3�⼝}�"��M{�g�]�Q� �v��Sttc��V8�FU�0-�ՙM����.�q�A����/k�ࢫ:檿��������������v����́K뙉��J�"	˖lW�/\ٖ�gnwp�Q����[|��nvέsk����Uۼ�������%��p��n�v �k.��j,:�ُS�kT��-:�K�כl
���͝ �bgS�ԁ�\Q�F��E�ڲK���k=��\�N�=7$�f��P��oD���SH6����e:�/��c�
��$����/�V)�!z.yn�'fG����P��cy�I�Z�@��n��XӴ���!�WSx���#Nf%�L�&�H����)�V��`߮[��G�����G�۰R���I�3���~�R�W�DQAfa&a�UueR�2�*)J�(��)
5&C1TK�5h�rP�TRSH5JU:�*�(�����Q�DіT�U6�$�*
��Py���7�<泓w�h���vZv���Z��y���d�/�$����IZ���DG�ad&�;W�Vh��\�T�WL�K�R���\@�����e��N���BK��U���0p�X�򧇨S�|�N�o������z�<4Up�6� Dg�ٴ���h��)���r:����x��u��6��Bૺ�C����i]���o�*��>�2�C�bԝV��9䦣X�
�^�펧:���9=����!{�CV��s�������L����x[�i���l��yj'�T�P�\.���W����N�Q+x�M�e��ȕ*fzC�w&�#!+�O��d�a�o�T�)Ӿ[���U�Bpp�px�����\e��2���R�p�i՚��W�>��Y�R���j�VPf|h֯�x��/<���߯5��J+Y���D�S���(��=�ϓ�|(z���=e����3�x�Z
�n��Ջi����_Ъ#���I���P��@Gu%kP
_{��D��Ql==*(`A#����k8�$�3����j%�,��u]t����:*��:�YPe\E�	�S0'�"u��	s�T��Ҩ^�;����hx��T�U�q�U��/��V��rgL�l����î��g¯I%��`���4�[�z��#���]xxL:� �٭^j��0�Y��u���Wk�o���/��Kj����|�k{:���m��N�,�E!�2�_�nV����n+�)�5�q�MxJ�f�v�z蒙���,\򥇅u�cG�X�=�� h�u�e�.7b�q�J �0�\�q>�]F�Ǹ�p��U51�p�o�'ϳds;};��i��w�����-�
���;��,H(}� 咳=O���;^��Q֋5b07��3z�����eki�|�TYvaNN{�6L�bMvH�`ڒ�u�L�-�h��M"�,�є-��!]��f�V�A��ޏx]�)��Us�����t �/�S89�޺���W�A��O�+0[U�s33�����˻�9j��9��d�zf�ף)�t�gsΫ�����u��p�,"i˭�(ij�+'��ṡw����sl��R��P6j���D!PO�h��j��f�L�y���q��� �qݦ��\�P 7��ǟk�����ޡPZ��h$���<���Ԇ^R�TMz��{/swո��")}ら0`�)���G�ܲj�2��ӿ
6"�R9
I�ԃ�֪��(�'�ľ@���W��u5n�]�kc
�*rX�2�e)5�~H�x���g�U�x���[b�}پ�=�Xt��+E ���xFN�~������\��y������Ƈ��pگ�v[t�L�W��jp�����,i�A���C���}/�����3�;��n�MJ�0��Ū*�Wwr}�z ��6�䉩�K��
3�p�\&�*�Dv�q*S���ow��ѣB����\�h�K"����J�u��n�ub(�RE��SF0��p����<7��pm�T�*B���A�)��i�#%j��u��c����1r&{/�cY�۩7�HI!�����\7���T�Lta��*sf�}ݬo�㶣$KJ��+|m�e
Ћ
��N�
�EE>��\������C�1������N�uW]E�!\�����|�玷<�mK^�.��Q���Ns����1���ʮ�.�!�cO�z�k��f���0&�&�"�6oh�	�T�N^U��{�QhK��a���q��:� S���4��`�c��+F���dB��z9�O`{)9��%�ߔ��eN�C&���1�k&��Y�g��F|S�|C��Y#����>I)��R�w��������F�vs�DWiR��_DG�no6��f���b�5}�.M��/
b�j�C�S�c-�K2��t����ZQ��Q��a󿛮
�= P�\��{�Ou���qp� [G���čD��!5R� �ߗ�/3��͍�s����ߕ �M�|>�bB��5À�i���{�� ��5ąE���ѫ��f�UAu��r&��sN��|Z���q#�(��U�^Z<L`���Uj-�Z��i�w~y���9L(|3Ɵ��^��;�3yW"r[��=ϝYB�2Ki]If�(���T&n2v��\*t�f�נhk�76�{}	����:�%��j��0�����.�VUA��P�=��>E�S�)���9��)ҭ�O�3����	�"��-�p�ir��^��9m5�Ȣ��a2΅z�vW�D�]�W��=t6߸���p�R�yed�T�\���Z���U�(e��L��
(H��Mk@+�DDEVE��?(�#]*��B�Q���߽�W[�]NUJ��F�/z;�����X �0@5U ]�#I��W���,�;�����r�0��U&�A��	�0u�8WL��Z�wV��'*��4^�8�pr3jj�R�4~�!+^����Q��;��x���GF�r��x�UQ&t�T�h*����j̨|��?O��֝�f�rK���4lW{��L<r�eG_��ҧb:�]s�޻�2�t�75"g�Sl*7�_M�LZ=�у�^uw�Nυ/��J5^ہ7���D��M�������^�g���t�B ��������'תO?F%׎�ځ�Sa��
m����V������=�/���9��E�
E7c��<���<,-p�*",�S
���W���¦?j=,���żëK֭�t�����6��bg>㓰��8�3M��������	υ���������(����J_<�����t�v���
q��U"5�ԃ9R�xWicG�lnzN�]��U�rl���TT�Sf�ɗ=�%}����]{W?*�U���e�c���t����|.�\�`���C�ob4�ΚӍ�7x��J,�U�4*�aAPm�Hh�/�8;��W~��2*W(H�����f��\^�Z��� +�)�-_}�++��P�rV��\��,p�����u^��|�
�,�r���l�i��C�T�8�nV����e�
���Y��B��W���7��e��dt�PqZ4*��S|:�Q���j���Dn�)	�q����*�3�^�X�D<�B����on��u4�td>�Ňz��g{yA�y��%J>S��|�Ǵ?]!1
鶇&S�^j�����Ե-NwW�Z����W9��H�T�+z<m�?>���*����Ok!�^��P࢒��T�U�����Tu@|/��ފn���`�>*X�,�zN�=)/�)����j����h�֒h�8�N\��&f[��k���".��]������q�w9�#G�Z���/Hzh&p&E
�'_^�,W.M"�y��'`���4�k�]d@*�\ �Zx�H�.6�S��������h��*��O5\<*���u)J�ˬ�I�y��NvjE@Q��3A�����>~PxA�r��S�/2�Vlh�!>,�t�8�Μ���)�b��@��Lh�~�gl��J�`��b�^�pe���Md�����+)�52����X�`��\��*�"r��.p���� ��v�$|��zzV��r��7�����/MIWz�}�o��n�ʏ�i��^k�#�y�&ol[��3��7G��D�j6^>P�j���j��s�r;�����/�ދ��ި_xnLڣ-�v)SuOʴS�Vꮺ��F� �4�\�w����e
���ʸl=����u�Q��	�-6�t:P�%���K�n@���1j��6�U���=���ɅӋ-�Kwe�Tm��rL���&��P��p��E4#�{��3rw-U4�k��C�M?\9kz#��K�4��=��{����m+�tu��´3ԩJ4a�}o��S����%�;�'�*%�S5&LJ��
������z�z
�@dٝ�:����.��L_��@-4>�h�@h�J"�|���z�i�P�;^f��Z�j�u��qp�L�̔��j���8%�<��z�Q
�R�<k��ZU�b���Ls��2;R�1����܋u��^�L����2�ξcQ�����^<{�zCt�����KU3�Y[7F��]��"
��uض�]'�`\4�"�J���ш�\V�H ���7�lʉ���-/K�J��#�E|�֍e�xWL�A���<�w��^�L�$)�ULg#g��Q���Dq���]�|�J��&e�lK�U
^Жh��3��*1V�d�?'O��{w�j
�5J�
(�͸3p��%S����X&,�3��44��ڗ�s~��*�щ�1u�M���B�Fz�ޡP���X�������
�ETF3i��O�_d���D^On���j��}<�4�C�`BI�.T4%��]�l�í��L|<+�vt�R�j�(SǞY�9��7&��C�~q�P,<8T]#[�R���⮢l�H����f+q4�1���Ϧ�����Z<�F�rK��j�D��>ې�z}ktL�J�tq4���=&���f�x��jv�Ji�h���Y�Xkl�;������J��1O�H�����
;7a<%�Oi� ��< `��0�_'6��u9r�iko+7��aԫ ���o�o'�q������ժwl�6F�?ZOp#52��pZ���=DJQ]�)yӬKYЎ�f8����k-*�{��(wu���D���4}���,.2���d\�����K�.��-��4B/�(�Zl��Sx���WB�($Eʀ�N�����@�-���]��w|�|�X��;;S9�u���F|�17tM(����K�N��P.�ņb<M���29�y�Dr�kdMŜ�w���Ҍ��Շq��[���O3��c�tm J��oe�BvQ�C�!�fd�ؖ�CVm]��|��EN�y��f�z���[پK%(�����xa%XGr�p�[Gr���C��S�t�|n�B��y��/�݈_��M����wO|�O��r������i�)�s6ф��,U��%uٖ6�4�N;D��y;1����:[��pɤ���,&��Nv�V2t��O�5�u��}�٬�c!�{���2�Y�hG�8�ۦcw�8y=�2Ŝiq}6��C��ʺ2�M�X��\�Z�X�Ҩ0i�+q��&�o4ZO���<�� ��o��A󤷨�j�9zec;��N���샺�����o��Z�.�{	[�ёӚqj#�2
�kn�����)O60��]�wC6�\�8R��S['����i�{g��C�A��*t���$E^�]�r��]n�V��2��].Ր?U�W�*3u�,�Am�]LN�Uŗ9<�ۅ���U��(^.m	�B7(�U���0#R��$njg-H��
�[EwV﹉Xv�5W�P*k���Sx�ew0�r��x:ּ�?�^�CCT��A2EMw�PA^�Y�f���N���TN���$l3#3*J21Ĭ�� �*�5h��'	7�u�ŨYƴk�p����3,,�mf���9A�~���X�M�;�x�+�3cw�ḓ���)�i�Dk��A|�l*O�{�/e��힑�w1����T�%�w�(�hz}��a�ٳ���ouǎ�_x�X��-�]Jg�$���f�=#����l��E08���4M=z�Љ�3Z.������t���>��vy��i�S�ęr�$�'iT�*�&4S��{k[#��Ƽ��Otd?b�4�uS�Z����f�]9�ɬ���f�n{��Ez�*��#U�䅉�X8WujcE����t|���M�پ������QW�>�UD���>���򪺊����f��`� 5i�D�.Z������X�i\Ĩ>G��w�
O�����%a�F��a�S88���gJj�z�u��Pm<s�@Q��/�#Ƹ�4m/*����Z�����z*��~�y[��D1Mޤ�����=S�V|so\���^][������:BT�'x栲��f���(]O ��a@ ��J%_���o���V��鮴W������C�`���	�x,�c6���������l�z.��ι@�S�Z��$0�}����A�)V���^���<*��Tn��a�S��aN�o��<Pfԁ���A���t��!�tt�b^�Lg@��wj;���w�œs6���t W�R�;+���%���H��ߓ��i�<8h�Z@���ժ�K�go�\��=�d��F��E�)۹~t8- r�T�����)Ĉe7��4`����sg��"�udK�S�ݱwZ����a�l�=2o�#;|�Ɩs�zPL���
5� ��+�}���BU�0����ݱ����4];n�`��p� ƍ�n�Ue� ҩ���*��;��<��>'i�T�����k"=����&�׊�,Ħ��%�GܟcV[R�*��o�Ζ�tKԷ@V�"�$N���y����}ꗃ4����'��V��8k�(<3�I3Q�^��e��&�kaӞʯk��}D&Y���P8xVY�=Mc��9w�z�n��mB�;M�l:F�`���?�A��Q���������nf�v��E�5�5�Fi�z|�p��`�aR�t|$��k�#�ޞ��A�j����݋����q�T"Z���$�Gl�'��� ���5� )��K��������l�U��<�	h�j��n�lT	��1���&�U�:��!�3�o{�xg������f�q�-������k�r�5U�<,p��4�K�cz��ە�{�#Q��U��U0 0A�*�@��se��%��&�M@uz��+��s��sJ��O(ѳ0��nxThE�0<nf��q��b����Vp�y鏁%A�6[�H����2:�G��K%�fi(��a�9�rw���Gn�.��]C~J޺.;�'C�&¤��RÚ�m\)�����teD�X�.jL��"c|H��]/n$�5L���H�H��uH��o�[/��*i��pb� h�8��[ÊJ.��	.�DI��g*-��Q��ً�n9Tn9�V]��S2�}���u�U&Q�^u�S���JN�JypWB���[�1e\Y���J��#�֟�����F�򷳬���ҹ}P.��F�E����Y��Ȅ�dl�5/�{a��� ��C9�gM	��/�����K�2ʵ/��(��qE�kLx�{��}D���R(�0�j�[v�AV�:���L<�Ǚ�1��q����M���T��e��1>S;�ڸE�5���0Qe���$�L��ĉٙ�!��Wi�yg��_S���rWH)5����T��T�1ga�o�Vok�1���]o�)��9��oF���is�`�+HZh����>md`,��1���$VI
�"��7�!}�d;�%��*_4�&F�ƚ<+���,~ׯ~���Q�_D;�^W
�۸X���
y�N�U������~PSˌrL��.��p,`A#Z��p�5>ق˭]��������Gb����_���q*̹�]UW��ui�x�Lj����Nک���
�f��w�X<��;}��4���T��\+FĴu�tǅO��J�C�M�۹��b��Qs�&�4j�d*F̙��f*�Q���(-���	�1w��oS�j�W/
Z�U������x����_h��	�x�����Y.j{(���@72n��ՒYY��n+�72�dp���Rm��v��!OOY���a�*��vV���cO����3���P����Zyc�LZ�D�`�
-Y���1AY!Ւn�q�Rj�!荎����+��b2+`��cc�s/o���G��c��$%��|m�+��O�T�j�Ez����UM.%I��>�������b�w���ڮ�y�u^ Zj� T�����f���C��� �������s�ϴ�N/ܫGצb�F�: �?1��d(��\����]D+5�>�^�w���@���]U�䐁l�,�`�x�.�F�LnP����I`�C�Ju]�p� ���5���.7=�t��hR��n�>Z=qUKţ�ϔ���y6Ʊ�ְ�R�0e\�A�
���T˜Jc�ǫ�ˋ�����m�i�&b���1h�P��
�Y�����+����(EN�#r��)�mc�p]��@��VtW���+h�]�j]���-w<�� T
��j���Ū���螉�@��(gO��=�I-��6�	*�:�T��#�<ɨtԼe�{�Ի���Uف��t��"��7��n�e�W�Nnv=��Yn�S�O\j�@�Ѽ_{׃�����u5f��A�8ei���[��JS�F��Y4�&+��opb�P�x�kK�֠+E ����u���5n���C X�~O嚼3J	�~,p��#�!����+}3�N=<����qY5�Э�FB��p��^Q���ug]!�v�a�xw�3L�a�K"���(<2:��u�+����jv���4s~�Ə��f*
�@��A���d��]L��1pj;��p�
Q0e�@{�&og"b��U\�D�c[i�Ba���:�;�&A�#��7�u�0fvj����]ӽ���F�|�����ҧ#]��ޮ&�gZ�8gӏ���'�����81�X8L�W��;P�<��b��u���y˺����NT��}*ߎD������̃X��˱�Q��&�@4�_S�Vj����.L� ��<7��<�%q]�g.b
@�.:�FΔW���h��_q�N^r!a��
�Z+��Fz����x�֒Iw�C�J��U͚�~+ᩙLMwQ��K��s{&�"�4kyV��3M4Ӛ�Y}'M�v�Ƅ�d��0�TH��p��U�p���&��WB�T�x�#	Gsw��~n�+x�0}���χ�h�2���w&k i��R�IA���j��;���������P|�} ��z��M%7�fL�QD�9&�@��'z�c���{�[1l�\j�w��4Q��52�4���D}E�uW�����j��r͜y�/G����]&+�j��;���̞���`"�қ�U��ꆀ��U��%�~{]s�e/��@�8L��U�n]�pyo�]1��>�� ��z�
/]|���$���gB���Vj��G�m��w�I��퓈E���G���� 97����sI�[�DM�tS�����ʡN��2��}����{��q�2�&6��:��LT��Sm�RU9���aWfe�-��d�N��Q��7��ܸf&�aL\�V��2(�Tj��p�B<g�n��L��X ʠpAd�i#	��f�w�yk�� K�k���h;�U�7<�4�}���&B�X=�K�sM�H��BNЕ;��U�_ed
�~�U���X&t:X�\�o�o����Y>��T?<ehU�Å@A�<8uV��"�㋃��M%�Q/���>����?#��/�a��P�׊+GmZ��8J��Mޮ�պ�UA��<'�;5�X�ӱ����\u�d�x����)���U�`TyRd
І=ih��g�IsžY�{�6T˴�fҒ�;Z�Y]�f�U�IB	}�"��P�1NmhA�!4���|	oy��x�}T�򧖟~�~�{��d)�Y���g� �=c54�Q?�.�seӣZ4N=z�Љ�3Z-=�7��^�M��[�f���Kz��%Z�%�a�Ԫ4�h��~n;���g?�|D}0��pU��Y?t}~�r_��Y%���5
Z��q��@U�훽Mz���^�M*B������O*�*a
��Wj{�/XmT�==����
��'­b�<<*�L�qz�*�J}T�W�0�(Y�L\FY���@�Ն5�U�Bqpv`���.��L��4�S��+`Ҟ5�\�A���ڵF��͏�~��o�8��X�Mld�i�0
x�ff3��e+���{[��߹u�+�;���]��D9^�S��!Ll�#��Q����a'���,7Sԭ��FY�7��e)J��Q��[(�²�h� ����:�.٥�<s&��p]$jٹx�Gظp9w�m>Ȣ�!8)+:��]�1�'����Z���J���K�T�� ��ǳ苦�gXٲܣu�>vF�;uIB���4)T��q��X �EY�:W¶N~ktᕢ��_^��ٷ��9�xj2�����Y�36�TPkFe%��+�t�+*4��Փ����3"��ԁT8���ˎì�p^
�e:�f�5�4n��	��q-��}�on�4��D��Vd&�;������[��ps��u�W
��*)c���ض�}o�+xg�9sF3�Z/F��+��)���u��FvW��8ɋ��<Gݭ�.Jiy�n��_��&Ƶ��������RQ��Y��҈{��f�����;�PS�D��^�վy��2�v�kc7Q
�WTz�*�t��ŎmԾj�	�:���.'nN��3h	r�p�����+r�������`cU�$mo粈���78M���e:�v�����=y���Vv�cn�y��C��|"(�l�A�!N�(b����= �p�z��..�eAu����y�g	�*������:@5ڮ���n�/v���2ދ���i����Ź��4� ���Xv]e¨��A�z���7�sf-7y0;Qo��Bj�'�6+Oug+ī6ZW����GG�mU֪�Z8����� ξ�hm�ϝ����d�T��$��Է�.�tzk��c~� F_mp ��J}���ҺT�ݤ��:e��]NBU��G���T�@���R�M�n���,�;p͸^���wt�6%9T�1`�@��9@���q^�}�y̴BRf��\2�U`���ۇ��I�L\ع��FC%�3�y#��Q�6�lmj�5��X�K�\�k�C�p�Խc�g=q�y���Up�FXn0�-`e�5ed�f9�kX�2ˌt�0��0�,��5�&"2N4kIG0�UU�IEa[�i�Xe�2�a���XFYfDCF��q:��
�ɠ�00)��3*
�� ��� ��Z��,-���*���Y�e��q�:��(�&'V��ME�U��v,_����3�~zJ�O`������t��dw��U#M�VGl	GY���������n3�U?���"�(ׂ�T���B�R�~8s��`�6)<�d��mh�MXj��T�����+��E�{&A�e��G�MM'�_����E*�`��׆��⦀U7��+��x��<9�� ���G
�5R���i}��U���SE�A�.`�F;��Q�����x�����p}*�o|Fpz�߻���z)3��ƸP�ZU|�x�
�P�3#����l��&l�L�qFN��/�F�Ǩp�����=��^=��WV�i��]���A�d��iS��P�è��|on�j6T̾�/3�>�*b�>�����T�u��.lqӯ�%�����6&7�:�4�:��}D&Y����7�	�ٶ�/8���߉�{Ѕs�n=Q�k3�W�>�-xOy��]�P��.�>��I���S;��e���I�y�;̃�⼛�Pߚ͛���s�NF9'�g�-�*c�:S9]1�*;��p�
Q^���7�靡r�{����/f+���nsj�rdr�[�|��`��,Fp��`
}�I	P����L)������7
����T滋�Q�XM����Z��{ݽR=�W�`��`�
gU*�ަ��9��U�+��I�/+�1{M+��ҁ�NDAP]0R�Ƶ�y:&�st(�I��'�Gc.��75:jV�� ��]\�P��[��;��+�8��g�z����J���<���u�O�<�l��^��ᚲ�ԳSS��ee����,�p�5����W�N�p�ֆ>B�o�� F�[EM��0g76���oXmA��qU��x�M6e#�n��/�>T��@��;�l]���g�&�Ŧv�ө3%OC�^�}���{/U������Î�:���#��\]��#k��H���0Fl����8�:w$��H'pI~zv�sm�����2��g�/`�Ȱxk�
>5��5b�pg�-ޞ�u���J��\�h:�D}E�uW�tg�*Eu=}|�e����ط�u1�S��L8%���ƹ����"�P\�]Fva�T���C�IZ�I����\b�h�fi�gp$�z�m��DO�N9Rfr�Y�~��W
sϬ�T��F���wT߽�i�V�&�){U!�E�:�U��jDnv���r�� ؿPc��աш�P��GcU�+�s��K���;��`Xu��"��pV	ʢ@� �u�Ҫ�&�zg{�⚼>�T��a�yW�|k�*P��,���_;g�%�+&�WX��j\�t[�X���T�3"��n�:f�i�#=��ViK��2,��L޺�9#��,����<�#�
Q5�QpǓ�epɪ_^��U�P�7k��2���`jT��ft����,�*ֆ��vki�sk�n�t;���~x�у� Ek�. ��"����o�r�S�� ����I�����c�X�f�D���
*{>��~�@�y�m?��qVY����Hm�w!<���&C�4���UT���u���˩L�V����Z���|EU	�p��3d�Wqq&B���L�W�*�q'P�l�8�i�RǾ֬1^��<)׭u�<wY�\�r�b�j"��m͵�A_X��od��52n�z�K+=[l{X�GI�l���/��MgE±�T��5<HC~�p%L,7f��	ǸIEEt�e_NGl.�Y���|h�U��U�bT����Kc�V>M����JJ��p;6D��a�D֮Z<2�BW�����փ�=��*���0�]r�P@��	A!Q��@���U�'�2�wm7�\!��md�g,�������޻���Y��)�-�&�Sr9�To����5���S�5�\Y�ꫜ깿P�+r��܁N�L�����x[�b�z}~^7�� �z�/0x�^R��U;.-\	s(�;nT�D9T�䪄��γrx�����)�4x�)`��=��eP\u�\�����ܕ\�^6�k����wSsG������L��"�L\
�@lU����A�\X_v/�p�� j���X7|!��\�S(��C�m(�mɚ�	�Z�p]�Ѿ���f���S��¼��P�^�t,>�T��hP�U�R��O죦�ЖjB�L]�a��UyB|&�s�1��� r�Ky}�{б۽�����|���|*�����A	��-@R������w&�Ǝ��P[�K~@�-��3Y`��PƝH�|��e��î���%��\mT{.v�\��.���M4[L9�vݰ��S��.%����
���9��TL���ll*�W����J�4��C҂�WƸS���u�]���{��.��x�Qz��s�df�_�t��
V�wc6$�� 6�kC A�8�8=���3L�^*����T��ȃ6���v�$���SƘ���n����x+�D�_�*;����}���5�+��
�AJ�ԇ�ʳǴحp=��7�c��Vy�"�.TUE�هq ���t�o�L<7O<\*��kd��S��\,W�+�#Q������*u���e'%o.��5͉R��Z@���2�D��a���9��𣋎����K�h�A\�b�vb���X8+�h�����,S����y:0��ns�#�>L���ypߴ�O�/@:���v{�dT���2�}ET�ף�"�xn�ٯ�ͳAp��h�"��I����@�*�a�hE��X���*�Klΐ޹qKB  IOގiw��L�Y*~�+E��r�먣4F�������{;j�Y]��n��Lj�7a�T��ʸW�
_x���fVE�/�9�5ze�1P�**d;iV��^��?4;ˇ�h�G����ާ;=�WM�0z��(��hԆ�����2�m��hj~>�;7}`J�V����� Ad5�}Z��x���M���N�!�0��u�k)�]LlI�V\�u>�ʓP�ٗy�Q�6A�LᢰOZ��ʭT[B�o*Z\.���	}L|��9CӜ%��Y/�2��6g:�߅��m�R�IZ�E����F�l�E\l�5�Q�̹39]+�Ǖ�e�SZc���A�nJ+<�Ta��ڨ3���e�
�ۅ-�R�|�A��}Gܔ������V�0:S���q����\�[���"�I�0k�ӭ嵆%x�ףO6l\�Pi�pv-/�Tt�Ùu��ى HYe 	+�E�����?�缠��-�D(k:�u�Q<uyu.�+�U�b>s���T���Uh���  e�QjBV@iR7���R��@u��;냾��R]k�[w.�LVc����)p��Ti
�g��\<&�/*�1��5Z*�6�(���QP򊩉�)U)Χ=>�UfzP�#Z8�����ޤƏT�J�����ka��W�a|~ʇ��=G����y��Ђ�w�/��}c��)�.��>LP�[+9��=�\�wٮ�Z�`vj����_2h_z����t��_����R9�ψ�MD�Z�4p���W�K��M@hD���{�p���M����~;y9�ř���+��Zx/��;���zcޤ�r����$�__5����3��i�jM0�/u�7=�Z���|14w|O�y�!�,�,�
�9�����ZF��f.�rfٓ-�� %�xP��"k+�������Nr:�FF���~�s�/�ՒJ=�����Q�{<o�eY�VSJ�
|uڨ��NN{��GVΚ<�Ql����\�[=���p���R�U��|*�������rwhږz��q�^�c� ڰ����\�/��ɥ+׎�Ow�pT0AT�����4���J
���ϣ�}@a�����.�L�u팮���T^|���9Ȫ�����/��d���!��Hx5ʗ
�V�k���}5֊�c��(�X�O.^��M�1\ c�M_=hP��9G��CU�/�8v��5�������o�5B�\j!P�'¼8V�^�����2] wv<���� �P�T�¸U� 0|�A���Ҧs�ۧ�6�q����DI; �<:�{�x�4�gJ� ��cX����[�9�%�#�o�Ө�àӔb�}1�Lso��Z5ܱ�c�l�Ź��N��}��G���R_z%��Y7����r�
V�<j}��_MDT(�%{Ng�y/\���Z���T���:2�� V�XtxVV�*J/I�M���	��/\��vC��@��b��AUʋ<4m�52�ή9opъ%q�]Ũ=�~m�R8K¥Y����!�E��K����Z=�7Π�4��=uu�ᯢ���Ѡ�)q�¢ǎZj�J�w�3ݽ �Z�uƸh�!��#���^hun��+#�)�˺f{�*ǡ�G�`�gF׼�3L�^*�4�\U�;���h2���v?9�/v����SXfR�N��O	�LJP%Y���^���T���®��
�A\*C�ʻ��b�����su�a1���qK������� ��k�yW������9{5?�z������їe\z�K/�:Ko	x:՛p:Zn�cH�Sm��Xk��s�5�%��P�V4���{�ڃ�=-��Dr�R�m
{1��%c�@(]�'�H5�ݮ	
6.��'k�t,,�������wk���ږK�}f
�V�,}�6���'@ef3f�nv����7�G`Juҕ��*L��ok��g�h
p�x��68�+R�Ox,��V���[��_׷J��˩L�yJ���Ӑ����	Wt���+:d�iح�ea����5ZWyl�k����t��YC7-m��8l����x2�tK��2�J
`�6a]�t��/1�ΥXgn��4y(��q�ZtUPv2��[�8�tW]C��k��4���.[���;&�J�xj��zٴ2��sh�Uh��{~;��/��T�쌊3�s7�(���4J�FuV�Sn�t�xѩE�I*�5N��ݻ� z�ާ��i<,Q6��f+��D����#��]ߐ.�3�kƑ>��X�̎N`�vP�5��(�]+�fr8V+�m�[�=\!H�1�l�f�A�ֱk�]��tZ�˗�[�m=�'j��Fd�!D�剴���;��X����U��r�t��*�m�������1�����K^�Q��MlTiv[����@C�K���q��n�Vb݅�r��[��
=Ck�o/��
*�47��6�U>�
J�ޤ5�2x�lv��V�7jv�0�kX]f��LI��_
�J�j����w�#-���	!u%`�/�X��M� T�^��z$Hێ�V4��J��x�Z��ZÕ���y�'R�<2�E[�a=�#��͉Ν�1�>�8_r^e�4eW�}sGH�;pR�g�˗%G��<�j���&h�H�Q���"\����u& �s����U�OnT����f�j!n�\�����,�[��z~� >�(0W������UFI�Rڔ��Sbc���fa��Y�fd��q�UPU����#VTVF1a�d�fa��*�*��&%�s3&�,�%'�����I���XDDFf9!fZ���&LMdӐdqM�wQ�\��j5��i�j�b����ټ�ƧPVI�jw��i�q�j�ȋ3)�
�q�B�x�VcI���hԦg��ݸ��+T|��֮1 u1��'UK�5�:ی�9��%i��Q�֪���}��e~��pT`T��J�
оF����7�t����*r5�V��oI��7���9R�沙��鋳V��Ѵ��Q��tz������sZ�/K��W�M_[����j!CP#F
𭸱rHV����꣍g�����E�t��_S1͗�]݊O�(�]�wG�ɮ+G�DU��uE���GUM?'�o����ow1�V��o�<\)S4,������E/�xt::��¼����f�]0%�ޣLt>��F;������V���u,��n��!픫�$ �=Y�5!�pk�]F_��@q.�*�3F�s�m\K�x��gb̹�QP�z��@��|kV��[����=���v�@�M5��*^/��p57�u�R�4׉��w��n\���ͅ=(:-�*N�`}Q�N̾vE;�ݻ�!Om��kG4��xj��
�3 �����nә����q�稷����P�3e-Ų��)/���I�U?.LAPl�V=�N����-.�4��*j�n�qq62��m��6gc*�N.�9Pn���C�IZU;@k-@���]X�a��~z.�tjq}��J�ڌ���?C�,d�FV����Te֧fɭ�کP��3���ZW�FhD�n���&����_LBg���6Qգ���Z��m�K�ɽ�@W��ٿ��ӭ�s�T�V���1 *�2�Ћ��.�PJ�m�"�w
���;�۸���U�zOU=�
�'����4x_�G�pgT����?%�\�K8+Q��2��VV
��^��5�^^'��� �`:&�2���w��YR{�R��4�5����_����_,?_��7:�F��m�0=%tې�,}0��i�>u4{��E��߅��3~C��W8�cv�n���ͺQr�S��k��e��mG�(�W����@��=�G�޽���z4 �~����`���K5�Y}�{(��<��~�*�hS�H[��A4������KG%<wW]<S=;��P`�S�$�4,�8VT#J��}�p��n���<����b���K��e�
�X�Qp�#�iસЁ�D��$~��SDh�Q��A�������k���~�p����f�wp��Ky5�k�:���CՄ�y�G��J���jO+���vD2,�������s<�eK�,�UK0*'E��Ɗ�P?�|*�>����oy�Y�J�r�]���yUZ�l:�MX`
ۯ�hw1��=����򇇸��-�
�t��O����k�����(.ԅ{d�q]���/�w��C�"�et����D��6��C�)ۛF��n{9�a�lұ�k�o	�o�p�̍M�n�wn��뤐�q�m3��޽'��LV[��Q���!}LLo��&�)P�ZF�Om���������Cm��������w"r�×0�����NA`�C��i�d
`��!6.��Lt�V�D��4)^�8���Q��A��qт\������*�T�`�H��kC�;��T˜q]6���Y���Uμ��<6�
0�0��A���:>����ow��b>�>5RP�����kx�+�˴��W�@R����,����
c�銤>
����
а��cP{�|�lwd�ɾ�Yg�-���)�+�� ��g�����mf̣��N�^�r���N-/�Y�?�X�@�E��O�C}ᦨ��lr�=���d
�� jM���a_�_���)��괠��|\ܚ��1������l@Dx]C\4p!��#�Pq_�ׄ����g�x.�s�E՝+&�Չ��~�lp�-@�p�vدq�X)����>����gijPT,[�s���h�f]���B��sd-<�9�qPu}N�z��lounrD��+�-�����n٨h� ~�ø�b��b�>�EP#�c5,��v�n�!�X���תyR�L��}�o���X�`eė��E��rЪ�p��tj
U�QE�ʟ�i�Z��V�!ӌޚ�q1SUP�<SW�W���ʼ4f��]�����m����
�h��A^V?�`p��;�!�u�[�J�!���Y�.� r5�C�L@4Q�>�{'{��4��:E����.�U+J5�T	�����v��΄�1�ʨ]Y����]4w��4WJ�|4 ��KUۧ���Ev ��k�8z�"�ƻf-�ձF�d�Y�r���U�A��Z2T\*�]U�
�(SǇe;��TE)���J��h���zkѨ��Wn��Iٝ��|��Gwf��_m��m���X��Q��XlI�}�.�����,NSmY//	���^�l�	}����B��3���ͣ�ss!M��a��\İ�L�fB���B����g=�թ }���h��ˡ'q�d��$@�Г%�Q2�D�~V�k��\9�(pۊY���+�I:w�u_��lՆ*�<�4��|@���惭�B�U&e������׽��:���<L`��Z��4�-�[ƴ(kx�l���s�E��]d��ϱm�������"�s#n"�ZJԊ��o4�"zs��V2��A�|�_�:�P,�~RH����Me�ˀ���j_#�u�-Mh�i�C3vwXV=��y�E�GK���)S���셂b�U���B��:;>j�{�S3�yk}��'�<*
Cx���u�3N�r�Vj�o8 0p@��l�h�:�T<-���P/Nk���Vi�.�E�;s�������ڡ{��|�ׂ�m��]�E*ܔ��f<BU/w��T��T�C"�M�)}�c���x`��w=�q��b|j��[�q����q�Q]j+2�D���e��(`���4�
�4��E��a�R��p}���(f����(���WY^�@�K�F�j�<\^�:+B�Åy�3Ѧ�:�{�r�u͉rUGug�}U����w]Y���t��:��B3�q�P��}�@���0OZB�j���o+W�zM]�Q&�����_�K���
�T��+B ���8	s���[�wt����lS�W��Ur_h�k�&W��:{��Q?&�W���Z��zb�T\)z�P�<�^�>�$y��҃��Ѩq8(Q�Y��tg��ed��L�5n��j�(��%1��Ւ2=�:�U�B�_�z)4���U	ᾊX;c^:�Q�a�ݑ�I�H �'��J�:�)��z�ۮv�N���;��Y�����ܮ���_�[��zF���6Dd}�mJ�̫������c3��ޏDG�;��%�U"N�})L3Y&{�POaUb'C'��d��ԓ�՘@ivT�wQ���˭fԽw�;6D���Ն5�yþmnI���͏Y��ς�}��|<��]����M�/���d���2kg\e�ə��/וҲ{�*/�w��]8[�Jn��$��� �Uq�,�i!��J�|+�Z�r6ܩ���Mwy���k=��t�����h�,"i˭�(i�#��v*��lc�|���6��R���NdTD�̀�5�A
5��m���.��;�K�=M�.�H.*�ź�uq��qr�)�J�8@,!X4�Crsӳ��Xz��88u�j5+���AC[���Ky �j"�K�M�>�vk}�X�kG������ V�4O��C��<gרPY����Q�@E�r�C�n�˴�Y�������sXmzO=��:v���u��L��tG
1�wq�6����l�͂�ǳ�QZ�� ����D��!��WC��0o��|���Ю���N����̶��1�,��h]��e4>EV(]#��z)����
tS�.�+ո�6og:�a��a�fA�Pe�_JW�Sס�@��Wz�n�����| ��ָ8k�����Gi��b]	��gD�mz��t���ym���"\���{^�W]p+)_Zݭ�	.'�6�����T�86�J�9R��:8\�k��h��ۓ���W�e��X�*�Z*��,�O�EQwr���z�k�jn#�%된'��jog&*f`���1��w�ل������q��YK+%��5J�F��hTXT���
����ǃS����i-�
L�P�F�a7:ԉVk@P:%�Pe�H�Â�h�r�0�a���x��g^�	�(:|oz�uA[\��[�A�P�!&r�]|���Fn
f��*B�pS*u�C^����[�8�E/�r��bJ9��)U�}Ǵ�>"���M_[��������|U꾑ǃlF��*�F��P:��Gl�H���\�y�7���-D�O};� à
�h�X<�눊��p�Xʌ�3�Y 7��e��ytԏ�ވ�xRf��OUyѮ�B���\_������`�%ZQ�B�9��\[Ǣ�ƙ��[鞞�>G������D��!5RH��~�����	���oD���@-4���@x�Ыƍf��ε�⡑xl%m�8�<�n
�ۦ�t���j�X*�t��uE۝r8����n4О����a�uj�?*�v�_�ʗ�\=�&�V
��5*�غ2�=lnɩ���
ى����by��#�꼨	�˱/��XY U��-�w� -5*a���wt�.;cY����fN�j#6�?%8kt����o��}dQ��5���T\�#v�ջ�,�!@�^3��/�B �Gi�ҭ��w�{�����rkno"/-�e�}��}��о9k3N�����S��v�f�Q%չ>��� p
�xk{�E�|�+��4�3�o��3N^g ���ν��Ć��٭�;u���´�;��$[�L`�]�JR=�R�����r�n��
f�ᇡ�d�+0���1lm��Ӿ�u��Q)�N�(>&�)�ف����Z����;���9ɬD����Aιmꊗ}���ү#L�.���0}���ސY3�B�k��Q|�ý!���t�(X��fL�r���M9�G";�x̳�RM�	�������]=hUÈ��GC�/�V$�J�R�]Cͽ��pvB���GvMpӬ�\���O�q9;�lDu$��p�P��sގv�I��/���qaXOvH!8Kb���@�[�ؖtr])+k\x���� ��[[֕�+���u����e���ei�gFR�>E����Q�b��z������xp���Ĺ�ЂUƾ����M�Wn>#Xd��qy����Vn���U��''ũ�v7RJ��S�W܂$�Iq�F�J��y���W�����鋕��8���BWa�5d�֪"�gњ�u/L�70lJ�׻�U:v�΁�-���A���K�@�����8̣4�5>���֣�������r��g^t����wl�����u����]I�:r-7���3mJ��.��^��!����nR�!STbXu����yң�L�n�gJ��3t�3D�g�6���;3��u������a�D�Dd��2H�]E7�c	o����
�i��Ɠ�WZ^#����v���c��&��c�ѣB��HR�P��`�q��F��c�C[�P�kVAY��9N�RV���IA��fdV�rj�݆NAM:�)���$30ik.-�D��lPad�f%�9	EU:����7	�!�e�r�P�`������X�Z����bVC��VA��f5�N����ރ|f����TV�$Զce�f`VXQSn�YQ�*�5e6c�LUQӬ�(��֭js32,j5��Vf��+#$�ʩ���0�R
#,�&H�,"*I�(�dFF1k3v�%�)���0�Q�dS:�'�(�Pq��2�)�eDA�(��&���8�1��REIIDQ314Q1h�*��rJr�-YMQ�F�)�ud�Y�ITZ���.#URAe�D�2�j�+v�(�-iʪb��)7�C�4F�y�Z2����j����ʓY���xek2�N޴SS�fbQ��E�i���/=<�~��jfǣ9#�9䫈�$��y�+"J�z�'���I1�����I�~V���1�«�F��
/�C�37bTf9�Χh@4W��9�J�j_j;�QQ�or�*��\3qr�����ۢ�2o�]K�i�S�[����(+7���`Tuh�&�q��'��V���
�TQ�/w�=�o9U+5���.���kg�s����7�+��{w�6�O�E�AøRj�W&�nǳ�ަk̲| ��0u������q�~��=�	�P�A����X`�5��(Ѫ�!�F��W��x�0|�:���s��SD��+/�����;30v�sq���w#oeY-�V~���0{�(s�Z8���*����peэ������<!�W�fQ�H�ת�*`i�+D��$.�]��ۑn�az���(����V�s7�E
q魡�sDbW5[�rf�Ԇeq�-u+w�jܖӜv�-�5�YG�;��*rA���$��8oyB��1��K�n:�gE+�IU��5��ǅ*�4�%OJ��<e��}գQ~���W���1b�"�p�#�#H�0� \I��A�Q�+Ee;���T�:3�W#6�V;��w �����,e�W6w���Ы�r�
�dz)4�
|J��*��JF��#u��P$�1Y"Sw��U��Л��;T�ݵ<c��&���j��
����\u�^�j��-�E�٢ �a��+�����w�Um�:=g�[<�8�O����k�-7�.������a<=P��Z5�j��a�U�o LQ�������Q��n�*.+�� �;���Z�B�R��ukF�NT�ō���:1��RXF�/)N��� ]N]m�H��Tyh�S��bo�6��tij�Y�]����E�^����/v���w�� _K��	N��6R�� u�a����+,�G	�+Sv����e(���:(㒎�;���b��|9��*��i#A>g!�X\u�S�S]2�ie�7���ҴT<9�Q�/ܸ1Ѐb�����-��<)���p�Vu	|ﮠ\�s�*��AUJ���i+����e%tEy�I���V�b��| �%�V�+B�A����/'����W��F�k��K�H�t]
�/QW�<4.U= �`��©�f�,;��aUL�H}>�]�<��Ͻ��zr�ZxZ��U��̃]@0��?r�U��4.b�	R��xsJ)��)ġFy �ׅ���-<U����@W�rD�
�.8�绽��Wkt��Z��x*�Tt jǙў�)��36���k��B����+�@oֈV݊�ʕ
p���u��ׄ`�.N��x���:��42���U��ܕ����i��=��i���}�Q��k�:.��ƚ�I	�%;�����$`���y�M�6L���C�i��q��IOP��(�4=��\)�Z��TuQwr���}Q6����hm��&o UIv�Y���x��N�x�\����� ;��l9�f�vk�z�B��]���!>1�_�ʟE�#��ƨ9�;�Qo��M����;M���s�iD�g����Ϋ"�9����]:��Ϩ5�uP�wJ�!� 8�7Л�}��<�9�:õ9؏4��ݐѨ�1�klu�;�_.�(� ����#�mB�>GQ���Ԃy�z_m��'�4]�H�@��l�f��N�oC��q�z+Q��YMO�N�X�2t`���sf�H�?���so�F�������0�Ws�.9�o���ڙ4-ۛ`P��['J��!J9	�\bX�q�(D�	�F(A�K�
�N�9�|�~�1�,I�sq�b��X���&��f���V�I�/b����;1_�WN�j졼q���.4�,&1i�~z��:j� E+���M����n��/��z�EC�E���MgZ0�mek�i�\ZO.�e܅~e���ж�6U����4rz���k����m̞M2�4��Q�E�Zj�ᑥn��X���vo |Jj.�}]/!����0�jf�k]�'�T7;s�1�nh��C�N�xA���*d���*�4r���RO)Bs��0���c쭔��v�`U��}'Vn]2�ZZ��S
�J�K�Do�I/�^cq껥/a��c���l��fd���I-��;m;d����7��p�n/vZ�6+b�4�`�����	7!t_,/�+֠��:V
���b�Mh�sQvnQ�@6�V^7��]FЂvr2Iy)�×Es-��I^f��3"/��-�&f��h���D����c|��o����c�Ů�@N�θ���3�b���^=�ۏk����qVU}좲�Ǟӷ3����J��)?����^�T���:��q=�0�2���s�g=�֖0^D'��q�t�{�W������A���釘���C|�Z}��ܙy�?^c�v�Z+�U�U|�4����ꐹ
��#�oI���|��+��-sXy��:���M��NJJ#�rB�ӈe��hC��[�0�F۹�3G2�j�S�):��^r�� v���. �n��t����Uu�I�$�]g���3�0�SG��gA�e����.`�����i����Ȩ[�-%�zȾ3^�.`���w%f�S/����qQ�����zL�/���
�F7����4�_>���c~���֑b�=�\({�P������q�z�]jۚK�SB$qI�k�^������F�7~��s��waS�g��Ja��4Y�w���良�S�a����b���v�����;���oAڭ�5N��@�ȶ�H���X��{dQTף,������%���/��O��� ���ك�̝�������I+�mF�q�:��VJ����Y���5P��xiz+���]��EyZ�
�
��e\A��>��ڸ{�QO�5�~�+#M+���,�Zm��z�S�7/M�[�p�sf)�����9�����և$����ȫˑ�E�zV����zl[Yv�2�Έ�L嚂���1|����Q@���̬�ݧw���)��ӽ!]��K����Km׫��MlS�nf�U�6�kx)@qy���oP�r�����Q{�"�VNH�pD�	{������T����z�^�rxg��M�GP�����f�(�o���Uu�h�WҶ���K���7M[=�;��y��z^��#j>�r;����c�\.�0R����M��P�6�K�E:J�6ԖN�$��@��;�k�\�����خh�%C�z���n(�@���T;c]������e�ؗ��(TI����{g+@Qq�5�.O�Q¸'S�੾4]���WC�-ak6��.1���fف!-{��Ll�KH(Ƹ�9�A�e�b�k�C�Gz�pp[+���z��ʊ̉���ޡy��{���g����k+Y�u"b��xޅ*�7Vo����9��0����NkQA�E���m��w5:��Ť���#._6x���z7�#Q�:�50Bgb��0���[O;����y���tP ���fˣ.k�5��ǝ멌t�����������E��[s�4�qU��u��x�Ax�W((���ġ5��6�\��4`��-��i[���ʬ�y��U�����L���y�!�1{�Y-�q����9�;^��d����dbɀ��ӹ�� ��28e?XH��s�7��r���S�SL�wF�WP3rF��z]�E���9*�>ݒmR�M�%r�ު2��)�y�����]Ω��p
�O��-U&쓲{[D�!���)���Fd��%8n˘��l����Bd0+2,��".�S��]ᛖp=���t�?T������ۃoaigb�2^��Ta���"�k�{�^��McN'`�F�^,�y�*��͜�R\��̧�s����oTi�����̹�����.�QÚqP:�7ڕ���' %+��^�ݡ��J�2��Z	՛e�"�����v��q.ۏ{�.h��R^k|$��M�m���Ov�t#C����Φ�w1���]c������g����R��jGZ��v�4�����V�u�չV+EM�{6����e�'e�+��'WL)�Xk�4ڲQD�LEә6��ź��q�|2N�˭ۄu+�x�3��۝J���[�*��=L�wb�e�ό�nb���1��_y�ޤ0�DŹ���6rmʖ�9���keG����ղ���φJ|:m���
ffF�G�c6��P���sww��� I���-���H'�gDN�����!�F�^� ӄ�Mͥ��}�{�װ��t��3�
�OH�.��r�]e2��Y/[3.�|�،��hk/Xv�-)�iʖ�&Zy����x�ΦE<{3k��A�.u���b�c��SaQ��O�~F����81J'S���Em���T��u��12ݩ�3�VK� ��!F@�'���xܻ�i1�}����tJ �{7��]e]���x����Y�P�:�G��L����Yc��b��������
�Wi�l��d�c9�q�#�Ic�,9��6�������ցw�5w��p-C\U�%�2��3�n���5]�$\�l��w�>'������Ԙ��b݉�0�vCzL�;*�˝`֋`���5dtԷ�K<.�]H�p2�NȈ�}˳hkW%��/�����ªhS/���@s���V�l�R,L���L�9):���N���P�U��>ɝ�n�2��7E<�WL�y����� � W�XIM�D5ő�+1r�" ���"�u���0�ʊ�0r�J��u��bɬ��RP�i��k3�d�&����Mq:�p��ʭb��PU4�Y&J��nN%5qA@LR�J�@��\��������������)(�5�����ըx�%�����*��5	��4��:�
!�u9	C!B�TY44���IJ%T%%��J1Υ).�p�
�+�(Z%h��.H![�}�ɍ�GGP~���G��R�tژ�Ma�7��b����f���6����Hg_��%q*�N27�H�)�1|]Vv�l�~TT=g|��i�b�λ��O-(� �@p����j��A��c�������*Z.�κ�Y�z�ڒ�`��yc�b\�UD^��Z��v�$s�=�0���G�%F�����^9'�[���.��uW��YB)��\�*h����Gq�zP	��չ$]WIĚ��r�q9���s 6T���S�Yʾ�;Lg:�C{ºr]�v&��c���>���u�av(��+�ّ�[,�?q�D;�&9�#�UL��9t�)V�(��y��ԥ�2��sԷ��`�.F5����b��S�gڦ���KL��u(д3�+�~װ_�����n���b)���M�O+�[�}�$��%�7۱�kf�U	���,ߤ����U�\Ǿ���t����?>l�UF��w��rs�*%EF���Ԫ.����3�F,,���Xn�B�v:8�^�X����Rx�Ɠ�w��L:%[�Ti�qE�L�Ψ��H�z�U��C\#!ڰ�U�L�$�U��X��8FD^]�c=�֘�Id-5�ۢU�%(���/ge���xp�.r�*3Wv>L�.�sֽ-V�M�	],�(�̻�K�/؂B�Gk�k�?#6MT�q�Ы�W�wj���2��q+m�Z!�s"��^J7�L�ľ�!���Z[���\`g�\G7�%�8���`��!("�ӽ�Y��1C싒��Ť��	r���4{�
����٨����&k���"���n1׃��U�C�0R��z+�c��T�� ��G:��KN��0M�l�,$�C���Ѝ���;K��5n15ڹ��9i�⛸]g���ʒc9�'�ic5����3�?{hz�Y��0UУ�f#���K�'�KmN��ue�%
�\P�1�y��x��v�I��9��ѳ
�r2$��9�;�r��_r���,���0 �<���=VI�&��u$濑숻�^�;ǩi��Ap�K3�-�`�n{���xd�^�t~^)��i��o�Zo5Rj�X[H����b��V5o�sA=Lнr�R��T�x����H�"uĕ�Uۈ$TR2"�a^��P��q.�\�D YP�*8�]K ��zv.��uo3��M�ƙF���U�H1��^oH���|�E����y��cKO�>I�.����Hw�O~�²
�>��b{�#^v!E�ٳw��]��B^��G/�Fy*��mX|3Kw0�w��.%�s.��m��ǜ���_1F�g���vs%Z84=uU�v7"cE��-dI�,I�[)���@F⛵�`�";���?[���-�f�s��Q:� dĳ>zG�K�N5���í�{x�j�]2}cx`
��.��J���*��y��bs�D�:�_Cv�㝐���SY�qqr��Υi�.;ȧC���$�h�"��gf���lt4z�����Z6X�=ݚ�K%�ב}^��x��è�[B	�HD���XW@.`��q"�Ɖ\��ͼu�34#:Py�=%�"�l#.9��j-�u���&���YK%�J0< ��#:�Hs����P�]���"}|�8����*�ʸ�.u�X���YsoN��2�WgnhF�It-�=��;Y��2�%���lM��ӽ;'RY��c�ܬ寒Nf�f�H�a��V}�T<c�X���,�E$8S��qm�Z���eEMs�"�tv06v^���8��^*�����wKA�3*��zXH�eh=`��;�\������ˤ�ф��TA��ux/���k18���/��ZX�1I�^��"g��5je���	��y�$_���Sћ;ۑ�^]�n{6�5�t��Ća�v^�/z6P���=^�'%gep@d]PK�'��Mv�ps�c��6���ޕ�b�����rwg�{�W���#������=~�Z��b:�ɭ�E�Dڢ*Lm=�3�E���<yV7��)�����LArP'����X*jj[2����&/��)(Lw	=w^��쌰���1�/��j1���{&(������o�he�De]�ȫ��sk�fZ��6�����pW6�DO=��_y��7TTA�6�,+k���q�|b���,YnE��s5�%�Ȕ����T�srtK��`�@��Dȵ��6f�%ki��;K ;94��׼8P���r,��AA��asW�`�|�d;�Fa�� �u�KM��{�3xj����O`�-���K%Z�4c ��OC��l��F1��M�Qo٫�;%H����;MΆ�S���V>a�	F�U)k]f���s����8���f���ꉎ�o�Gic]ڱ}S�h��e�U	׃6=<:	rDg>O(#N���]K4ǫ�ЋqPi�txz�Ջ��Y xv#;D��.��/��~�f,t�u���.QC<�N|�1;l��r�߆N�Z>���ЛX�����=�2�l}�Y|;F�b�	�vLF��
���	,N9��>�M�
����r/:ͭ	��w�#I�v�H�@ӡrM���2m�e�c����#���{P��&ف�U�u��5�(ռ�Q$���S�w��p�)�����m�:��U\5/ �f�{w��.3X~��m�w����|�Xr9���g�1�>갫H=��Y�]�:��$�_U���P����2�����"�?��:u������=�[I�	�RV}��;�_�}�iPE���ם�k1�z��n3�J�I���W���W�q�+��4*�W����1�/�	Vh�7�6�EW�z�Pb��ǃe��j�KIOU,w!%	���m�:��t'[R��� �҅K;IVz�k����j9��%$�4	nzN�d*�5�S{��5p�����k�G�}�Y�Ђ�Y7�nw���pb���;��I�?yq�ނ���v���px�#�0�{9gxC'RX��4��f��5ѹ���H^Gc�f��n5>{��k�l�Wmv²�$��Ζ8�Y���C>շ5B	�WZ놵�8��n$Fƭ��(��Ց��ֲy!�-��t½�`84H�����6�W�V2�y3��ߑ�n3j��IQ6��6͢#����7e��1B����i���w1��؞��֬^9�UZeo���\���*n��0��)g
W���M��D����S/d<eN��ط�f��9��F�N#�3���[�e*�%��!ɼ���E906��giY��U�i��Ia�~��6�ૼ�
H��Pr\l֠��Nj!��T�1��/S�(�Qn��D1\�8E�/��=Z5F�G�me�N"��fɪ��E����+ԣ�Ae�A��8�s�	������n��jk$��n�8�;4��h�	7���=��S�\��%rT2!���E�Imr�;:Oof�Z���l����FvQw���.�hA˕[ӭ��q��m�B�)9Grx'D�P"�;��ބ�e�PWB��1����^�x��5?GЉ�Bb�
���/�<*��v�������WS[XΆ�b�Eq�����G��Q�a��-���Ѻ��$S�XOF͡�t�5]kC���]\oyި)䫦�j�͢�gP��jrm��$�#���6�`7����zʎ�K��Go4̶� u��t��|��}����+��}�M��P0iy�H�"�1v:�h�q�8�Z����U�@j�1`D;�;�r -���n�Ի�Š����Wi<LJ+����qkW�տ��/��Yܰlu�Ӫk�t�̭v��\���B��Ȳ/*��ۣ���nVf���=�n���,I� `^s!���8�0mj���0�h���ϐR����m�lk��� ��ɼ,�C}���u�p��D�W,U7zD%bB 6u^����quH&�P���u�Ƴ�W�yt�G)6�
  7����ײ��l��|QT�ָN[��
yR��f�A��wQ̭}�)�.���nP�� ���+�Mt�C����s�L Ʃ�p�7}�t��b��(����0���9fv깤�7O��j1T�+u�n�u�
�km^Eq�}�.�&�e�gS�v7)���#�oG`�ʺ�閶k�)a�m�k�5,G����q�AAQ:�	�t�D>s����X�L�r�m�-t�寞�wGm�s�����}�M�W�/s{��q���c�/Co���Э���O{N@�7����n��XR�(Em�VmǚVm<��BD�]������lIV2�g�����y�J�/��:�Ss���T���쭦+2�.� M��NĜ%�k�,u��	��-�)��t����b�����M��Ţ]B�wъF�Ǘ,f��"ډ�P���46(�h�͢d�H�n�1˸o���(����Hb��g��]l𻃸��9e���o�:�;�uS�9(S܁�k�)JT�B�"B����S!O �h
���]CJд	T-(P�P$T&��E�-�T� 
�������
(R���MȦTM4n����i)B���4�T� �R-;�& 2pjB��JA�
@�WR��Ҕ���� �e%QB�P(ҍ4nL��������,CW/�A�,�k�����9q��z�1�R�^P�r���L�� �SzO�?�� /����29�!��k.��K�z&j��paP��d���v��ou`	�����61�@3Q�\5aR�e,�����S3/��=ykZ��_���ϛ`���ɸQ�����Cq;aY�J��f�c[C�0L-�����o^����$�f���4i�lm�b�{�&�h��"��P�7�8��̼aI�L���)�K�}�Sl��v�\ci�ާ�Y�&�'����l��,%����#�T����[\�t:�`��m\��kswW�3m��4Z�%����32w��k�D�S�n��rX��zΔ1�)eJP����x��A`�{��r�ћ֏�r��8�r��J��\JQ��zwnuM ��W��@E���X3�)2��CG��j��ڍz�p�����ͬ:�%� VW�O��4\���]Ûs�;{̪����&��\���@�vm�Ϸx\�Iٓr\jwǢJ��H��w����Bhw�q��4ʸ�U�I��T����k�ަJ��6��;"��͸�xfva,��**q����Y����Θ0��.�le�b��+J��KV2�}f/��N��y�[U�vE��b�C	5�������<Ț�w�`*�km�W����;6��'sv!��D�]3�����خ�p���h�N҉�s]ͷ�tD�n��N�n��Iʰ&7%ı<Ӑ^жtH�N�!�Y9䎗v����L���	�/�����#7���io��2O	��`3��g�Ic��خ*ܾ�%�Ov�I����b�W�d��y}'$�X":m��;}b1��t6ݎ*��,�8k!�� ��D��ܒ.���)�ђ�H��eb� �7�z������Lo_�Jʚ'\R`Z�Z�%ŝ�M-�l�H"�<�Kbuk\�F;�K�{"^vQ�怣�U敔_t9��S-d�Ԯ_5ӝ�sخ����HnS(�m=�e��yE�Sݰ�y��T���;��e�v�Ķ�Q�%���|;
�VS��-5��m�:��*Z��>���R��fjc�#��tg}%�m��MD��|�>���З�_Y���ӻ$e(2A��:#���%Eli���Ռb��9ǵ�&	|�Jn�!΂�n�nY��kN�9f%��i���eMk�f.1 	8#:�{�c�%~p?oX��3mX؜������*?*G|�����.���$�2�[��PI@���!��b��|�A�.D�s�A�L$.�a���1yyw��_+�y��]Pcvs�A�������Fr��D��-Y�����h-s+�?v�i(�xSӬ�0�<�� ��x�zv�P��Y��bW�I����y7 -"i^��G^���p��mT��+��w�e],{����x�ʽ�U��h�d��|���Z���L؟=v�0[��^�B�c��m�3bRar�rT��>~�jq��n�L�q�r�_���|R���9���U�y��X�!��j{����:^�������=�(����W�Y�x4ߜ��`����b�UP��qOd��	ՖR�W0!n�V���r���sڙ�6=�d���4�A;��UOu.V����n���('b�OJ�uJ�	ٛ[��SP�t(��ǫP���v��V���2(���H���c��x�����3u\<����|y�QP�1��_����'	����e����v��
��ؐ
����u�ʼ����Ga]2�ei�}�8L,x&�2Lk|lN6�S(��

9;�6��w'j��W]�$�L]$�ʅ)y�r1��	���,U����kU�R����V�F+9�uG�E��&r����1�uvr	֞����a���]Ƨ�����X��ZZ�=/�U�%�b�&��~��Ҷg-2T^L)�c�p)�w鍩;s��Ik�|ox�ug{G&�,�}�ϯ�YE�c��F��3P��w�\X9�F�7��`�~�p���ݎ���2�u���2C}Ԩ�K`�b��n�Kz+t��;6'wB���n�+��I�e�S;�����=y���Ѫ^Cģh�H�@�u]�N�����'�����c|��g�}Ǆb=�5.�(�h;*�mZ�n�F�p��5�.�k�j�����jt흍��;d/ctL�>�����pX&'$�޸��^#�V^�c�3".0�j:�O�t��Q�{�Z~uN���xCY�fCl��a�k�,�P���L�͸���3��zmn�ͱ7���8��+�F4����o�PZ�qHɓ��WMb}�%�3���`�K�R}��|u�N�U��5�z�%��=V�FL�ǭ%l[���n���E�s����&�O9^#=�ӻ���Г�Z�k�9�o��J�{�=o��	�d,�"�U�^\�k�����a6W�T��轕��`�,�_
��Տ�O�F_��%l΃4I.q��մ��u�v\��܅r���͸������k\�T	��'d��[
Ĩ^=��Ǆk��R�Bʔ�\��()�D 
[(+�6NOɃ�e�o��D@S+�z�����/\�T5kK�sN�fD���Nujy�+�IE�LS}�)��µ���j�s�l��v��y�ԙ[�ї�a��ke������u��@�ڣB�LTli�����Z�u�:��$�̈%1�TH��3h��t�:V�c��,c.��r�8�ň& z/r$zN��	�]֤%ݢ�@1Pm_�+R�W�be�D���w��b�t���#6�[w3_"��+t�!��N��j�ʮj�g@����I�]fW���Mv�ن1N��'��^��P�������U1�W8.��&�}-��͍7��Z�o����}��*N"o�lU��n��"���@ T�^�Yv�7���f��B��#��@N�i�I��~��mg ��h�᪔�Z������V�s�&[Y��k	��ռ��&��
� ��&qҎia6�{�w���35$f_0	-l��A3���{ƒ�ד�+l�����Lp�E�p/���&s�OT�@����.�e+>��U�*�w'�������5����2-��:*��s��n���t]���h�Mi�D�k�~�Q&60��yI��=��e����ne<��¡[�+u�9^o���VV$�Y!%��{֯ҲIA�ܾ���Δ:}���wtn���X�5�M���!|�X4�Ƿ\�$�ͱ/���8���,�9㙬�	�Ik7�Vb�{�(�ԭ�0�`�{,�](�l%��B���ݹ�`elf����щAy��e{�pe7q�wU�e3�;P�Kcw\�U�v-�ŒJ@�q�m�~��GXW����E�~����}rhV�pI,m�+7�$��b:���:�i��l=\�7j5��%'�E9��$�\u�wPس|"�l�/S�Yn�Ev�f��f9sK�}b�d6F���>H΁���'_�V�\��H۝�BJA��"/�+j^E�;���1�b��Za��<tō��;��ٳ��:$y�*���,�������PT5a�pEAP����C��'�2D�{���/vW��ڰ��
��gv	�&�#��0�@"E�Q@��(�d
�J ��~��;5�F���811�3�C��&~0^�dX�T�)j�ic���h��j��I	!�RUo��+�q����z7C�����|�R��I��
/9�ౣf~�3���^_U�Y2�7U[93�u��c<s��I$$�ڍ�~���ɲ�I%$�:$�BH~�I�!C�(����vG/�Xx#U�G�'�=������x�~��bu��J���BHh=��.t�JR��d\��*E�F.�u0R3�%�~��m#V�y��zH��kv����y��s�gZ�w��ȦRץw�?VD����>���G�����Ca���m��|uBp8���?Hf�A��|�͂8�����0j�D����FJ�URY���c���Rpz^�1�^�+��ؘ�:�y�F;��|��nb���Y��ޛ�~F_�����I	!�zZJ�W�9���;<!���&�
p2�e�l-"�dy�-���ˣ��X�1'�v4�y}d�/Q��y����C��T�V��})EG��)�CB�S�,6��eKZF�H�!E.w"HI���E6��wեU�θ�cږ5�&��1�7�r2o� "��r�� ��@Ӣ���D�*�I"$����i1L�$s�W�7����	9�Y�`���a4�<��d!�9�x�;t��`}L�I	!�\�t;ޖ�R:!$$�`W�ړ��Q�w��I�}z��j�Ū>��9���.H��9�Յ���M(����Ӹ�|*=��D��9�a�s�FWִ$���xN8�8��^H��A���#H��脐��ۑ�q[%߹��l9�Oy��ڜ�������ڌ�(�
��{<l�R�\�����z��ձ��dmQ��z*���4�f�N,w��o�BH_����a���s}���Q����)��o�N�����5Y�VV�ъ0�ǵ1H���J�I	!����r��\z�Ѳ��=>n3gK���HI�:��)2LL���ɑ�2�,�IP�;�/�R7�T�GdS�Y#�sTM�fs���"�(H>�f��